BZh91AY&SY�ku��_�py����߰����  `���    z      }�4  :

P
`= �xjm�a�q�  ,��  �@�P�
  �8 �>�Ĝ=�V�v���g����>�zn/�մ��׻-��f�k����������� !{�`��}wji�����t��:�N��{bO���������M���:�Y^�ڰ�B7� ϯ�=-�v���8�{U+ݻwu�{ǝM��G3��U���y�*�V��7FW��l`�o��JF�f�]-t���òsOP�G=��-���eֵ��n�ɦ��j���  ��M�,�v�>���]�r����Gt.�n�k-f��wkkl��� (P    �      �?I�Ԫ�M4`L&�  L�C i�)��`      �L4�(UH L  � 	�F&��*R�&L�41 L�LM�	�@&�2�3*mOF��6�4��&�*�40  #FMw�Ȟ4�R@,�b���DB��C��{�D4
�����x���W�_���ar��DD�"""n��1TUI	A ˀ���<[I$�H	��*��C�����O�������$�y�����Uu�91�������K���Yh�g�7�>�x@�5��r��5�3��G�����*�X�V->�Q��>
-X�X+�UZ�5�R,E�U�+��R�R�ɣ�X��TK�?"G���VѺ ���nکUJ%E(uW��U�`�.���3�7k[=�u�i��e��^b~�qR�\Ux�O����M���y�Wї��Dx�#C\�
4[{=�9�-ᶲw5�g��oaD�Z�s�zŸ,�X����?��M\҉P�yB,�Xn �B�j����G�C4��J�+B�+�{�-�WKJXZŖ�ҡz�2�B�E{o�\��ED���L�A�)��,u~��B��]�1���~��:��:�8���rC��y�ҁ1xo!��_�L��`nE��q�؜i̸�ni�9.�,�qC�XT�e�Ż�:�R�R�j�w�<�7�녉���%��:߆��ٰ͇��ek�f�<�)v:U:�yO�7.�����-���c�kM�)�[��m����C5�:��蚘�dۊb�x�cD�M��cˈ��<�l����[��M��W���X��z�1ݻ�Se�jE7�b����l�!�[��M����X�y��߮�n�e��7���p޷��-��y������"0��F��9���2��Ǽ�޷�:i�Lm����`�G���n���2���D0��,�<�7b�[�1k�hmkk��C��K��[��HҘ��67y�e<-�!��J�l�������,�\2ۡ�U:��.7&3\M�z^=X�<ʼb��I�kHZB��v���Z���6����ι�Tꜩ�rC���F�kuL�~~�Wر��5��w[��ɗ��v�ٙY�.��d`�i��*aӔ:25ޑ�2�al���o\F?[�7n�f<�g����f�G�1�a�G�8!��E��:�S�NK`����{��dKx�)n�1k��d7��o�Hf=�c����LU�M�m�1S)�llmc[ˈ����6Jczߛ��66�f�t;���s[�z[-��m���#\c�1L�S5�`�C��n�N<��L��X�y��߽�v�91�����1�o��-ىߖ�^A����fDal�y���їN&��i�N�cl�k���Gz��ݻ����1����" �����n-��S��k[Z��鱸�w���@Ҟ����<lo6�{�tK<�dk#[3�/́��,�\2ۡ��7.��*6kć�V7��v��^T�"� zxqP?k�uE�{�g��Ů�"��Y��E8BBBk[�Bg�D�z/�hZ���0�"��e[Ec"�E}����g�
P��!��68�3j�j�lX���3[��z�ރ[�n��l�������*#��S:w;�V*�����x"�7_H�ʙ��J����&�4M�BT�����1��؂�P�[>�cb�,�]R�z�R�?R��8R��הlB����ʊ5���bǻL&kbѰoU��ݢ��c#��#��!��1
��+�[�pS�o���u��!�kx"���7ji��4AX�8^��|b׫&!T�Ezt"�N�{`���x[��E�#�S�
�v�U�F8BZ�����D'$� ���Ϗ�C��ϋq+�DK!J�<������򊈁�"ܘ�b�"|���^�n�ť�(����q
��?y崉�$�ʾ����MT�}bo�X(kp�Z���&�hW,Gۍ<�^�o�4!i�oۘ�`흻;�U�c�gf#ٻi��0Nt^VJ�ɫ>�>�t"E2��)���ߢm��lDk>��4y�Y1.)0S�q~-����V�Aon��E�!�y�)�,��,�K�$!�6�W�<؂�p�l��<��E��^�DE2�������}#R5��"�t ���6/��^���b5�O�h��W�~�y�����d*�������?
�xC�
�Cq��Z��nD�HU�Dz�m(5�Z)=;Ӱ�Kg���ֶ]��Z	tm���e.&�͘�S�K	"u�U�."b��,ģ��ʔ~x��)�\Yz?51'�Z3:��� m��H��4�(����7��Kv�e���U��I(P�#���nwb[kt�35ʹW�^s��fq��;L�����y�{��p�<�~i/m��
j��a���Ё��M�����oA��μ�#O}Ԧ���Y�a���C�o�)�j�<���j}u���,5�v�i�:g
+۩ӿ�k�M�������S������n��N��~�ߋ\i)M�/�����q7�Iߏ�s��x'ƺwd�އ�,��3ǃ��TO�|.�'�}�ף��u�];��=����K>���}��a����4�������'
��LZu���|�񭗦�u2�w�վﰾ7�[5���s��y�X1g�;�T�s�)�kf�wA���A/���IЧ_.-��h�@��ւ�ۻ��׼	�O.�m98>��{S���놓z�ovy;��:���r��\������Ϗ���ɐ���x�~�!���l8rNx�Ŋ���*zzMv��2������$�[��c/(WF|��u�c��|��wݞqtn�|�y�l������5ӏ]�֝�v�>E�[y4�N[�q��\������~;+�G�+����6�w=<���ó�sr;�/O_9=��b�vH��<��q��m�X<����.��J�N8m���������S7����ܭ���n�w�o�ܺ��{f�ͼ�%�*ҭ�S����{��߻:�n�VI��#O��'l�ܞ/L���������ޤ����7�_�F{S��R�~����c},����G����y^��(�y�^��_����jR�w�~g��+1�?M'��#l��?MO63}-1f������}�#�7w�x_�/sj�ʪj��_�#SH�	S���sZ��A���r���r>�RFHs�K�oVY!=<F^뷳����=7==�б6�z��v|�Xw����ɩ�w`�d$sU@�p[k�:�=�|7:���%}��~����#���ju;�a�#7���I_/�O����7��㷱��i�����ś�i����׹�[�z�dpG^槟x�=ws�u�s���Mx�J_~���8󟝿q�3�����=k����xK6���<�H��v��<�{:m񁾙汒{T�w���2�˗*�ۦ8v�[̙�R��m^�m�O9m�׮�+��5�EEx��nUӗ{��Æ�<z�Ƥ�EeӖ=t��{x����r�OX�r�+y�e�j�˧l\j�귭﹏j^���ۧ�m�uyr�Çlm�d�qt�˖ܽm��=�n�t�u�]������ae=d]=t��r�U����oU^��XW�a��m�z��v�+��:��'�mX�]�v��n����m�%�u������t�Çn�ۇM���۽�ͼt�޼u��z����ҧ��^nG�㭾8v�X��׮,��=m¹52���^��73s��6���z�ӷ�]��㧯$�'J�|�L��oX�ܪ���9p޹�gw(�:Ǌ��o�+�ܹx�����n��n���Q���Wy��n^1�n^:z��%ܶ�^�W����oN:v�]��=�54�e1;q\/3}v᎜*�=q�	]CJ���<os#�Mp�y��O[t���ghq�	�z��ǯ��Ak�wWq��p�֮א+�t�ӷN����C?n���Ǯ�=�#�����n�om+�&Zj7����Φ�J�`o3o�m[��.j6ܖ5�i�F��f�<S�|6��h���+�m��}�
�шW^jD��m����-{ZBS�U�ao��&;�c(VY��0��s��9�G�;7!Q����n�-�=�o���U9�b%Z�y0����oB��t�u�͡Zg0��tܩ�!�@����~p��y!}����Ǔ�!�e<(O�e��yN�A �G�G������ծ�C���=�@��T� ��*���x5�c0A\껪�3��!�3g,�	o���b$�F_6�jV���V�E�Y(a�[�6$!�<Ì�V�� Pͺu~��$�ƃX�r��� ��e�CGfZ
�FPV�Ql�2��Hf!���(7��31��":�e�i	�ё�>w�5T��`i�,�	��_XM��~4`�֬B�`���D3:��+f2U�.��YA%ZIR�ү���$�,U�sTé+tL�ʻ�$���[�
�Ls9%�l!j;% S�P�ޘM�@�T&��03ژBQ���[I�5r�Ԟ3*��h� F��+!D�*Ң��J�)����7���yǊ�<�h��6�`d0�ƪL0;�n��9�'m�ۙ�S����3կ"7�dT���؇i��?�h���=�?�<�����PO6�����<�yzq��s�s����<��  X $ �    �` / �  �   �с�  X � X��� �����w@�aW��&!	 �$�������y��9�7޽ D �  X $ �@
  � P��� h0  �@HHH@�  'wvw^�}������/�o���|PV;UTm�     �$ (@<  �	 $ � �  `�  @@HP P�  `�����ƀW��R�_%ɯ��wu{�����2@<  )  р `@ ��$ �� �	 $ � �  `� �<�� �b 7ov7w| ���|������}�K%W8S3�� 
 � �  ��   �  ����  �� ,  P�� � 6 	GB 7w5�� O�/�����T +2���@� �� �	 � X0  0@ �   L  �� �	  5� � (@����\9�s��{���Ha,L��~#�}DD BHF'��OO���/��Sg�>D�<��}OS�قmӷ��i۷��QS>��Z��*�B���ڏ��)�N�����U)�T-B�^X!j1R<�>>>B����+>�E�zP!X��E��j1Z)I�Ȅ�����*^�Z�R)y@�����+'�`���hϷwf}q��A��Э6�YT�vK6�X��L�a-nc�ˌ����YPns(m���WE4*�)42m��m����m�[ڴ��h��Ԭ��It��X�:�2�X8�^b��E�³;�޲�`v,���-R�hh�
��`3T��4?	��|�ʖ۞�XۂL6�d@��a?~~����貄�m�[��74Δh�`��@�	W����7�L3C�0���G����.]�mIe�5�"�i.똲�m5�#���m@�3q�ם��[t�ƶ�<8��[��[ga���.u���R��T��Dv��d����Ÿe�@�6���ն��ȥ@B���E#D]lECE�j�Ki`�0cQ8US����\R�높�&�E3�],e��K�ml2����r�&VгgXRmT1r&�����`&�͒�F���}��]^lU*�m�f����"4��ll��/�n����E �R�F!�!�D���4��^7�1�8�fp�B!�l[���aJT#N����\XV�n���$�1��ff0��I��3qmpˬí��qV`���eWcVkM�ف.�7�u�i��ś��[Jj��+�IS0�(YB��+T��)P:�AW��ٖl�&f�L%�5�Wk�m��F�W[F�,��h���J�ܒV[�X͛jT��LO2`�[��"n!s~���f�9[4�#M5$6]�c��^8#��Y���^[r��;s���[e�5�tWB�i��c�v��,,�&�}�[`��X��(d��|���.�#�te
�1��A�{3KE�mMG����Sm���]�ntͮe�˥nM��Q�2&Ȫ�V� +,E��!��]0�-����nF�YlͶ��Mkv�X��[��Cm�0�F�(��V��:�P�sk�c�4�]Wiuك[I[a�3���s�P�������Zbi)�a�ʞ�'����eBvf�fL��\��E�	�S.A��	d��'"1�Mv�������8�[��|�r[�h�Þ{B]�E�5[*do·[�8�е�fl�kn�$u`::YM��xW�c�M���!eѲ���6�]��>����ML���7��������ak�ia�s�2�f�mv�&�m$؎e��M.GYKX�K���1�\�;��������Z��l�����>��\��h\�5%���麤6n��SB����k����������K �vQ���S4��1�ڍ�n[�243��Ku1�J���a/n�l�
���`4a�7���g��mF[e�[�Zi[5NĶ<���6�P,%��ґ\�n�e�I���q)����d��A���-���%�@SIL1��QK׮���;;Sb�:�d�d�ի�ջKf��Fݪت��m�>��i}���m�v���	�ǽ�{�1����$&]��33<���K��˗wwL��,�o�@���{����>9�/a$-|{�����9��yv�$5�3��J�`Q�jS�F�ZЗ�ɚcfb�@�8�E����10�u%
����96;m�uW���n�%�@�mm�eY��-۬�٫V���u�k1��m��[u���0{B�E�gVT����L7K�Z�鱔8�t�kƒ��"�JSg;E�CF�L��C.>�>��y
]�6���m�n0sC�F:R�-����W�U��]��k�XDh,��18�hDW #�i��]�	ev�R�.�����/k)��e^t�A%�[�c�+����k.rB5z�����Z�X�j�A`���T��(ǭ�6�-�j�t�$��������w�U+�!�	S�@pNg�u9	s5I��܆�U>ud��@��h8֌%�.�.T���Z(�	A�nt5�M�^%J��=&Hz�̗E���%��M�g:^L[�:��y��D��K7�y�$jx���+1s֤��1���pY��a`c];����J,Qђ�kI�9�<�� �C����؅�fkH�'1���g�}>�F�"#	�����_%봾�Ki����n8���5�����{:Mqc�;l�
_��&J�(�G�K�����j��ATx�ꋩY<O�A���/X�fBa�|�����7�Nq*�X`���	[�	��+�ujJ��x�t8���[��B��.�,�Y.���2u��	-�p�VQ�tQG��Ƃ0�@JH�h��n�f�]�Ha�M/b��v�x.c�X��'���	�ڈ�*�'�V~������������:IN�'x�+*�m��le�����\��Bb�sS8���������*�j���b^��ܫ��L�xU�L�*Qb�̗	�����Y��9ˈt*��;\oI�h,A���s�+2�x�5�K7^�Qi�s!z�6a���h	ͼ��u�O�O�d��	aSy� ����mSz̲kS�z��zz7��ë��)�a��/@� a��(3��g�aF��l4������f츷uj���T��������YR�I���8͉"�0s[01+U�T�X:2]�����ƥ�-U����Ku^�hiث��1?=����.�Ӄ[�C�pT�2F�c��%T�d�o��r��.&��3[���kd�P�xd��n����տJ�T���m#C$���3�
jԭVkc�5j��
�Ņ��..ePl�tti�dM�$���0�?w�J�cP��^ Hp����"���|~��+	�i�� C!ЇÃ��o\��jv��Q2�N�
�r�R{���4ߦ�5f���%b�J�[�K�3�Uڨ���`�L˭M^�:���y�vI ���b�:hI��όCn"�#Q!�����ED�8̈́׵��~A�b8�c�_G���~!��+�W'�<�)�Z�>t��G�'��px��G�6���'�pt9O��O	����ׇ��� �D�6�W¾�[�~
؋��.�bO�Y��&��������G��>�>D}I�G¾/�i���̞3�O9G99!r��#UE�|��X(�Q�'_�ã�܋��C�3����A�>Q�'����7��ɷ�6?:���#O��(�I����ys������Tʷ�n�Ե�4��4��5#���'y;�j������n�z��'�ǡ���O~�w��of{�����b��тb�XW���ך���-�N٤y��l֜��K��^��5�bM}{��������y��,E�L�U~�?��y�]��339�{����wwt�����n%�>�ꙙ���y����S3<���o��wT��,���Z����We����.���(�``�0�0/p�h�Pt2�PȚ��/)�'� 6�#�]�K���kX���@�c�l\�~L��xB��O�U(:p(d;�d8	�!a��ӬP3on
E��1!�	�p3@��\��Ke��\�Eݟf�{QE�����	a�A�bv��Dh���3�A��@��F���Z{4��� pGY�6�cP�=D�W�*@� D���n�T��x���zFL�bEaln.�=�)��0��M$����
+AL:F�����e�٢��xb<װaL֬u�*��7��6��8�Т�(�b�e�a��j���v2�,�YF��H�������a��8kdl2�f]km�f%�4>N����&�&�L���22\JJ�7�EK&�5��A�|��Sŭ��D��L��@D(1�2�i�J$E�����vB�����hvf4�����cX�j+��)��B�8= 6��)�)�5���u�m��x��u�#e�٢�̙Έ�:�	��(��Bd�0��Q
5)t�	n��ED�5U*���X�R%�`]��]d�rf]]�'w���!��8	:gx3E���K\K..*LQ�O��(8 0CI�4,y�b:�Y�Z����.2]"��r����WX82��c��4]��G�^;��(��(@��\�0�l��U�ɝ�
M�� �y�BZڕvt�*̆	ћCQ�����(PL���M�`L���x�C�mF$��7�z��ٹS����&RE'���j�wy�Vc��Ҙԅ<Er@�j�Ђ��J���������V��䒬�d�N�.�j �)mY%����U�/`/���3QE&A�Kr���f��� ��HtJ�K���e�Z��w$V��;j%��`��|B�m ��;`��3�7��a�(\���RlJJ�T��ʰ��=D��
<�6Q��=�\��v��gA��-Q��g<��n���6L��wfO[�������L�o���mf�La��JIJ�r@�[���uD49��؄� *�v�P�%�5 ȭ@20��A���N����~Q_�����g�ש�ކ�K/�"�����f��s�d�T�k���\�e��˛�&���^��4UN��[�wL$��6Ԙk��=�1`�!��FMJ�`�ʲ�:h����\�G8�:bO5AͿPp�4|�|&a���>��(��v�W����HI--Qj��j� YA���ݞ���(䉩�m�鿳�DvЁ/Jݻ �����œǋf5��X�� �0Ɖ���/�W����!�-�	aћӡ��}�lnv|c��kd59g���ɞT�L~��~Y��Ӻ|N��(����7.c�50L�9Чs�|&J���E!�����dd!}�R�Rj�d$�w}U�P8i��n�&M�K(l�	�D����q�f��Dʋ�����~Ȣ;����&7�ݢ�N��)��6L���b�.��2d�����9%��f��8Q7������if�%�,��(�˙�wD�)P�	� ���N���8�>�k�a��#����ť���n"DG�'�O�_�#�~%x����pr9|5�sá�;<'�I�2>�>Q�5�\x��	�һ�.�v@�&��x���;~��؟	��/�:'�	��A��N��d��ڧ�'�SƧ�׉�����ǈc�tg������s����������8��948=0>�W����'�}O�<;.hq�i}4r�YYvX�Ğ��=�s��pJ�����_�f��X�S��z�$疫^{ž�Ao�����t��vU�������v��i�X��cM(7z◡�<槅V�ܝm�\&�UM��yd���������u�d�f}]4\��j�Cm�&�C��Yl].Xhߪ}��Ym�8��������O��wT��.އ�s��\t>�}��33ˎ��o����w3<��}���:���g����}��*�6L�Aϫ��p�-�	�ݒQ(d�-lQ�̊�f2�l�,-Jӛ��3���W6���rҬ�5.6�M5ɮ�V:B�a�]K7�s[�v�d;v0�H���R�R[���Z	���\KB*GXjCE�a��aFPDZ�ųF��Mն��`�[*�F�f�3}-ˆ�[�RY�֕���[-����!�R�+
˗XK6�[5�8-�˲�Ur���-n�ؘ��R��+lv� �:�E�f+�h@�@�M4�h<*0�QUZ��̶�x%��t5HF����:M��z-�i`�ڶ��lĻ:᪅�dݥ�z[��bki�B�qy�Kj���Ǘ��$B������i�Շ��a��g%rJ�{�O]�7��y�>n���L@+ʝ,�g����1R�k��vQE��9>�'0��}+��0^zj���}T��2&�ڙ��W�ỶT,���m�����/�-�sk�fD(�R�4HN&;e�$�oZ�(� �4B���C]+A���11���؝�Hb�8��n�Z6o���Q��NA�C��4�3��W3zZY��'\t"c��+���_��m��
���>�Bp�@K�x2L$�bt�rW�ڹ��10xj%�I���$P�Qh����3%�!��c�_��l�d�C�xD���ʪ� ��[LT��(� g�ܝ��/n�+�$VE5��]^X����d��2!r�l�����=ˮ��I�Ћ�ѐ�e�`((�}4Wh"U�EF�9�3������f���cQD)�����D%���>���WUiiK޼���g���_}�n�c!%ӏ*'(���X{�x�!�0=�F��T�G��ġ&�;�����q����&.J,��'�K.}�v
�r�Ɂ�� )�ۘ�>�e�X᢬�P&:[Pie������1�S���罙���@�b65ԑ��M�%f��2�YP�-���Č�v���u��Ű^�lMHĹ���ai)aY,j������`�3S=�c�2oA��LMj{چ&����Sٚ.�u���l�9b��UU �$p�W5]n�yE�x��(�Xe�;�d\�5�C�)����jI�
(v-S�hF��im��]h��K,�|��٦���14���Sնd1���e�����o����53�>O�Z&+J�M�$h�}���e$�9����Ľ���DT�5P���#��##;OYÁ��ϒh�$7�F�3)d�}9ކÓuD�
5�X�=271<|2��$�_�>K�2P}�S]�f��d&�C�K@�p��rtL[�M�5K*K�]�����%��Ÿ�)(V�\aZ��$'�ƻ�i#Je1�ά\X��Z��&k_@�|?e�>Iϸ�j����uR��M�$��~�əFj\����Y&���ӷ˝5�-��~�Uz�Wx�����ϻ<�|������+�ȁ5e��#i��ɲ�h5���Q<Y�}S4�5:�x�b�� F���,:#��""/�d���d�@��7����vd7�Q>ٝ2K�����ᨖYU���x�MQ�X�R��s(&5��.�[���#5fY���M���F�2��К����m�X/6�0�.�g]e�\X�WXK$j����D�L��D�y!g�fD�a�qD囁a�y�PL�+3y�U5NB�7<\���a��GD�!��ٵt����;�0{a�t�nď���ZX��M������;+N��M�a�z���Bê�T����ᨖYU���byI�Z��I(��ق/�W[�jvɀC2�t����sF	/eY%�+��n,��2��n��g������V��HWg�l��p0Ϭ��w�M���Rw$��(5�q�k	�����G�d٠�v�`�9�f�>!���?	~>/�
�E��$<4��p��|�yG��/�.��?�$>?]�/�xv�O	㳧�xm��F��>Q�'�_
�t�	�`����1؞>^x��xO�G���v8�~Q�3��
�]O�|93��:�w<>7������Nۨ���c��&>L|���TT������������sꇩ�>e͎4M�M�͌�.��a���?�?�����5w�S�ܿT߫uM��ި��"~����0~����i�[��i��!��JmM��5I�U!�ى����=_M����4��pu�<��PjȜ/;��>��+ط����ZN-�SP�Y1���K��9�OW��������8wGwe�Ur����;�.꫗����wU\��p>��˺�������������ǽ�2o���ᔐl��������]���i�4�<�
�We�d�䩭˹>=e���V,$d�,#\�7T@�����\<5cD�p�7ߕ,��}18J&����`3!�i&�/��[�n��#��.bl��J0)}�<�%*USb2�@ٹ�;�p��!�|�a׿?`K#:�����T1��n��G�n�t/_f���5�ʢ�։`�&��V����ē'�����bc��/C��`%�s�PF�w�`��.%�|_�b�Z42����=�^q�I=#3*[?;��[V��;a#�& k�S�!Q��Kp�7@9W2�a�!��24�S%f�M�a[\�e�f�mHڵٚ�DR�G�;�'��߿�=&�b����;�C�2��N��;
'��^�b���͹����N{�N�X�l���Ƅ�%}�`j캲��de�]�}+���&��,L�>��񑨔6`R�)���% p#9&%�4���rXj��#>�\��(�M{�3�wR�%\���3).���n�WW������ζ��B׶�!33D����>��Zm-��֧�12pj%���|eY4���U>P����C�*W�o���]J�J�I��w�c���e#�ԒBx;\���ju��+U�^I*1�0� H�$��t�`�W%L���EG���N�d���j{D30ِ~٨ɝ�|3.d��J2)z��s��tHny��;/$��ԛN͇�4N�ߥ��]Sr��υ�rh=(��g�URVΤ������NM�{����������'b� ��U��j�i��:�d�쪍�D6bTɑ��6tR��WK��'U�
�RJ]��!��t͛R,T,�WZ˦i4Bݵ�f�m�#,�h�Fh��j�ͭ�6�k�0��q�#�na�ٿ�g���H��D��`Pf]\��L���U�Ś�f!�;QC0s|�]�1�4.�<���������,[��ҋиh9�O�L�8J���) ����Q������uĉAn�G�<*W�+�ɐ�fw�N�ګ�KݵEQR�ԨpAԘ���5�esj5D�J
�R���xN�j���굉����|/`jx1������Ӂٴ���ԢM��VT��2�`��H=0#|��3 �J��$�n}4x���d��'������*����V+���Ut4Q�����D�2�6��0a��s��j�!�Xaz1��1������wp�:�͇B��6\����J�'ᵹ�Ë�bEK	�L[��Õ\�~9��bW���WO/1���£1m���%%d�\���HpM���$���\�D̰�\��O�۱�i�S5�!��app��|7���N�!X���x_��;<Ul�	��~���< �N��'Tm�Q:�|�_�(��SĞ����良�|<���|C����"A�|+�S¾񸉱Sj�l�����������RxO|C�Hl|�>Q�6"�W�^>!��g�|np�;��'�Ã����ى�|�|o����a�N��=:>�6zi_S����c<�>Q�:}O���p�89�6>�{48=��A�w����9�:΍�l﷿���s��y���E�Z�VZ�ܑ5YQ��k%���N�2��ڬݯc��Z��7T��wu{hw�m>z��=uS�Gu���z��ow�\֢�r���Cv���fkK{��ֵ��7$���5o8���w��w�z��q��5Nj��Nc�5UCC���՗u\�������˺�]�����YwU˻�#_ww��.�wtDk���ue�W.}������sCX�I���%�ܒCK#�6�ۓQ�v%Xn�K6�®��ݟ��e�E�*&M�c��ƥ%�e[۰���a�8���Γj3G9�Zk���r�Ku����袹�2�`{D��Q�q]i�������3���E� �خ�aH�Ej��˴E�(B[�Vj�%��Z�XEٮ��3G��kqn���mIt�)֮�[w7Y�Q7��ڭJ���du���M��q��������i[6��)`�٩\�ۗ6�F�6���h-����c5���	5���Zm���+6ƛu����8Ռ�?s��{���J��&�K��u؛)[lqH�V��5[��D٘�S^�؆�Fn���N֙��䗀�q�r>;8&������d�9���I��o>�Ji+A�\�(�OA�� l.��1�A�+����ff&�EpLx(7�r���v�Wv�X!ԡc X'p���%6���Ap5���E�5!��g��P�/�U������9����<�I��h���P��C~ރv}��v�|�џpT�� �>đbX}�s]�+շRvz�q� �n�ӄ�T]�*�rvo��8Y�&C�o<��fr�	����{���kQ֙�p����T �0^�!���$s@oa�M'�9�bg2���L�\qLr�x����[n�7�(�_?7�R,v:��VЎDX��ء�~�>�U�V�((�(�p��>��V-A����#�fB�.Po{�\��j�x�>�Hg?JO59(�a0��8eѭ�l�_q%�׏-`�D��&B�7
 L��r�&o�X|���d����$*���a;B�p�#�A��;4��;<dt1��b���f���0<Q�ۀ�}���d��nM��v�]�Ð��qA��+}�B�k*�0BzJ�����V���CO��q$�%������p0�M�FA�ҘY`5�� �%hQo
\\/S�{@��٘I����R�����*��K�I��iE�|��}�����ݘ�yd���&�VHh,5����ZԵXF["^0��.%^~_-~�g���V��B<��<�ou���k�[�^=�.�O�|�]���%��Y�p[f	v`��pW�Qk5|��C2B��Y�(��M���%B�&�CY9��I�{|�MJ�ܬ}������h1�!�N�M`����jfv\�ٍϻ��KY�5땍��n�
=�����R�bĢk0MC2���>�G3Ɲ;�Xw�d2�5��0SE$�pku�<�<�
2Ly��4,7iM��2�zCچe\����+ �?H��F�;��?j�Z/��v"d!DY
�DQ�xo}I8��:����`��Ã�����M�����>��3��UU2�^+�d����"��jA�L�zfQ�ΞE��d̰�b��rq�|��'��sBmB��[��w��l�I�E{���d06jЏ�a�+W3UfA&�d>2��2��[-�d�Wy^p�o�7���|k5Dmt��>.��`�?
N�{>������RK�4j"1\�5-,���ʮ	c�h��nr3�3ZғZ6�;D�8-����Ԍ���.ijj�]�����sY�k����L�@3h�*���C>�C��a��;�`8B:�
��~XI��5���
9��<`6Nx�M̜���?K	�A�c"�DU�- \"r�6���\�!f	W]4J��&�ԅ�*e�F@�=�m%���I=$��>th�$�G/�	e�����qK��ՇZu#��Z������ð�ɠ�P[�j$$����?Kd$E�6L��5��(���3���T�7.���S&C6g�P�-f�ÓE��^'�x����'�8�xAz"�����N��D�D�E���ñ�s�xkG�gķÿ�ׇ�!�6=rB}	�#�¿
�*|5�Щ�C:D�|8~	���į	<N��D���Ж>Q�t*xW�^�f<Cï(Ά(�ȊMr#�D��*�O�\�w���g��<�>>��M��'ڊ`��'�Y!��|+�t:.sd����dޢ����lg�DqO�aĻ����n���/� ����o�y��s\���u�Ɠ�&ְ���O^SOpWFG��E���t*�����#��F�(���ݶm�6�ފ���qqמy:r�o̜�Y~��}�{���׷+����S[���*��aκ�˒���]ϡ=}��=U�u˹�<}��=U�u˹�<}��=U�u˹�dwwt�V]�.�ё����g;ֳ��}�CR�x�>��?L��rH��@2��y�~6�:�jJ�R���h2d5(C�ͦEA88:���'��	�K��pbL�\s�Uoʶr3�J�1�D���h��fC��͇����f��Mg����՘7��Lg��h8&���(�fXԬ�%BE'�3\�w{��o[���c�jj|�f�^ʹSY��ٞ�ݗY��$��X�5�k�(�Ю�5)QŅ�«ax&�!���|U1�z��!G ��Q������A�fx2SEb�b��o\ˌM��91y�M4���N�����eM4��sVi�����h�2o�����X@~!/����hS[�ф�˟!5E�$ӥ�Z�kq.|%ٞ���m��Y왷Ŭ��)��@�}������f��b}8q�>���>�.ìy4n0���5JXc}�0�Vܓ6cV]\t�s�����U����r�b�`�*|):)��DNд5`b�Hp������䯾�'�>�փ��&���/�I.�Yu���|@�v��}0��p��q���e�uP5F�4��V�!��$�W46)�+!��n�$>ѱ��8T�����L�(�3�6��r`8�/7e�\�����E���T|�]�֋�rk��C��r���PDR���T��Er���4���.k4��ye���Q��VqےOk���3��������߂��B��nhbtz)Z�5�����1*���W���@�mwzZH��I{/I��j'��u���ځ��lߤ&3U��2]x��o!�&}�r���J�k9��k�A��I��`���62��'G"�b��P�mU-";�7����O]a�=�b��QwX`�:马8&�u���]�4���饄�a��^�T�&kjJYl��7Lbx�F��	7`��kO�@J�<Z*�VC�!A~�5�pA�5
�|�g|8a-��[����}Q�� QJJXT�Y��l�3��
�g|}�rL������)\��r@��4� oa�o��<����a�Xn��>Le��=�"��Q ��=��%�qW�����`>�5��^7,7,<L���5,b|<��V��1] D!��Y>�dśl>LU���c.6�jZ��Psd3[.� b0��`~�>H'"���2�۝�}Յ����2�AscApS�}\��/��Ke}��Tj�24��N�n�m��iV�|���b���ӘD"Z�٣�ka�����(�Z3X�垃�#-��`�'�Ǥ��k�5fg��ۭ��a�gJg�w�Y��I|	y�YQ̰23��p�ə�yT�{æ!�|.!g�0}9�^9�*�����'�_
�GqtǢ)�Zꉕ; ��O�O�_
�i|'��~×"xL���~&�	�;���"A�$�>�|@ҟCb��]��,�˟	��>�3��C�^��GN�Ά��v+�_��������|rp�ۃ���ٙ����v���>;<'|C��G�&��'����e��D�GԞ�:�f&ǟt���ɭE����ؐ�ODx{C���Ɍ7.��6�'���}��Bq�%#�.��R4|�|7�=�&��F�;l+�Q����m6��*���ۙ��Byj�x4΁���7��ۥǿ����n	ݑ�]A���zskQ����(���f�ǡ�v�q�)��i!D'�n���϶IU�u˹�dwwwUUe�.��q���UU�|��E�wwL��w.���q���37[˼���{��1�g�=�9zxbx|)^S��8���)ɫdI�Ǫ��ƫ�e���t��h�+ �5D �v��kv�b����Kdq,a����u[����jݤl�ҷZ�2�����0�}
��Əݡ���qn6Ye�b���
HY�P��������)�i��CԶ�Y�Iy
c5�/�\�3�o���%���Knt��him�ڷcm�iI�����4)Ѩ�5�>����È^�'� kh�#+$Q1`Țn*��e���!�o�ڒ�c�сv�{[16:�2��� ��ߩ$���4���>��������	�Sں�+��-��,�=�����V���"��������"1�g�ipE0ʴ������Cǒ��׼���ye�pl,��\9��L�<c�W)��-���,T�܄�c�4 t�}a��!Z�&b����Gv[�����L�T��B��St�{�&PF{��������sI�$:����9�B&xoqS� _��z�Ƌ(�01:;��{�:1�J.�lhTV��dNf"�4��y��fOL� �n���c�(&�p�Y֢ZͷVӼMd�#)4c�gJ��߳2x�v�뵒K���p<B�X�l|)4)|���'�oeU�b7��^8�m(D̍���e�m��c���Bs�X�ŉD�]�'oNj���8�����Mt����3҆�z��2V+I�>'�H}ӟ7%��}�f{zw5,O-U��i���tY�]�ik�S]����.�� V��l�i.[v��f-໶!d�Գ�SM)x	c�+D�V���_u&ֿ��z�ˬl.�Aa�	���Y��*�4���UFfo�� %�Mg��'��%�RQmu�0\J,�_u�Y���r���l�U�Z��LJ[K5塊k=;�~{�M=݌\�+����~���uD���tv�pQ�u3_"�����׹l�	ce����9ݝ�|��UUU,�<�h��5�UUV�gy�plI����6O���1#«����azxR�e`�P;���}��ݥi�ݤ)��^�QMk��VE�������U���59c��>C����kGC!��c��(��El�T��ȟ#h@�0Q���f�+�b*y�iG�0�l1�)Se6QF1�c,�u.�,����C��+�A�9=쇡��a�;&�=�R��E^
f7GL���hMD$'2/`D>�\�蔣��Hy���\�1����{�;�g��O�{�� ��]+{Ͻ�jk7W�u�@\�,lj9%]TxYJݠ�!l��R�-}��0%�k�]���[����? \�ϖ$����᱊����7�Ϟ�2s��R��u��U>o���%��$�͆O��@m3ej����ʤ��Ye�� V̍���.��Ot�DD�f^{?���	�R���	;,btO��ETЩmh��e͍�ۻ��U[��ᩔ�cg�G�o��X������-iW2������a���H�*t�:[g����>�u�å`<p��ɣ/&��O��[�}����Bb�)�)���t�M�;������O:��4Y^<c�)�-X!�J�Mj>����P!]
�,����R� B�`��-�Q���)yD&�&������^�Z�E�R�<�M��=j�SѳWJz����B㋚�^�<����Ƣ�l��\^���{=�[��매��J�y�n/D�Q�n�+���5Zz���z����qol�B7���/k�j_����z����W�)W��ɮٙ���s}o���fn��s}o���ff��s}O���ff��s}O���ff��s}O���ff��yɒ�^O	�x����+��9U3�2�Y�P9�ʰɋ�z�b��ၩW\�ۿ}��>���Y/CaӅ��j���MK���zwVJ��<d��ƓB�ɢT��<I�g� �KN��V(����X��Kg�>�������Z/�O��wwRɕD��D�PL�O�ag��o!�ѹ���v�M6k��ё�ŋU��V�A�*V��	��������&����
�i�5B����H�h�"�mB��ю�Yi�Z�F�4��*��٦p��KVRcv� �@XY�m�՛U�G��q��L��R9A�V��ͬ���gUKIwI��N]����8;Z:���YZ7�jT�g	������6\�J54r;�5�"'���'E�����Btԯ4/��*��A/��o��0���!'���)��i�h1M-���難�c
���=������0}�&�w4�\��𣢼QU�xVk�%]n����z�w���\���`�*�}�qX:����(����U�u(���[ꍆ!�-0�
�Ӫ�x&��S����y$��2q.��\Ρa�<gED$9���>��_�k��/�J%�L�m��J�2�b���2A0Cz511�M%C�|k����UT�����YE��h�C�צ���M�<+eA\���^�[Ҭ��J$8��j�=UTDv�e��i�N1�tn�q.��]��x��d3	w)��7D����v���ml��g�a�P�!óSSE�kRN��g��sux�g�A4'C}^V�U��Ыh�-�5(�"�OFi-�'Rk^;/"kD,���vV�*���am�m�l���fC!��ǁE�yW&(�_C!�u.Yz;\�|9��&m1x��b�V5�0�(<֫�&%Kgjc4���5≙���G�l��׽~2���}��������u���b�0�_�b��s$Pj!�㪨$�Q��]f�1�d��p3;%�Q%0��̂:J��I���х^�ī�&���$����w{
��ǩ�)�2���I":���)�4��{7�'�f���ܷaA�r�]��6y����+�~�	D��c͞1fΝ,�S�S��M˜���~���Bb)hR!!�Oɣ描��'WԹ�ԭ>\�O.U˕��j�yd#��O��	�^�YbJ�E�R�@���B�l�Q�Ջ)��"G��ԏ��Z���m:^G�	��g5�r���s�Q(�z.�vF��\�!D�Lq�9Nk�B}W��*n���v/.޽8����5���w��K�|�r=���D��d��wM�~hu���/l�\��{�+ "=%\�;Q���j��^������u5
�%	���W���r�o��[�� П����{�v�n�|�|�S��陙����S��陙����S��陙����K��陙����K��陙���90��xQ�<BC�{ϑ�.Ԥ�̥+��@��M,���'����)��4�Yu��&��fn���rU)e��a5�gBn�p�4�͋4�ͿO��/�;������Փؑ,q�A6)�� ׶n�B�Y�WB�v�7:����B-�54��J;��,`��6�飒���f[���C�Xf����.p�%��I�pIn��+�mâkhauͰ�f��&��a-�H�m���J�1 u�"��iFCӶqI�؇�Կ�5�֧�/�g�qk3�p��f	�B��fz�&ţ3yn�l���G���e�N��d�9K?$�i���ش|�cC@r]2ZZ��0�jhmi�l1nMIts�m�`���T��a/0�4ۢ�m�b*�6G���?s��=Y�r����0�	�����	�ka�wRH|�����7Y]�$�{�L�5ו���&��c��1y+f~4GcI�G��	˴��9J��j7"5f��AX��Wwr�ɒV�#E����[����_����~H�D��T��;d�D��UD{OUlI�ϒ�~�%��w{�S��=ߏ�p2#����8BJ��|7Э��3q�>�i�!��p��=Ua�w�g ��(�6��v��d��m�D~���$��|%��nA!7��$�;U=�'����;����1B�
�荍'��$.�Hm�\��:=R����߾}8���r��m�;��6���d35,6;�W�ρvsj�2C�@��N)i�2��k �Ȇ�li8(�!!��i�A�Z���Q��gB^1�%���e,��n�w�fĠۈ���z�#��旯$}{��yZK6�K�j����_�Ąġ �O֠l�br�Ys^�S��n�"���&Q����
�����x7��9D��4���9�)���p�M�'�����W3����"��5X<JN���u��p�nj�K.��%����gC&���t���2V��t�f���'"i���_�1�\���v{Uv{iE�-��L]٠��5�fkB���xQ�6B������va�����V��W��Wv����D���t}c^�q���~Ԝ�"�SΥ�y��m͛:$�Cc,�f]��Uc��MI8x��<&�T��(�GE�$9�d��V�8*�BBb2$��H��!������s����~`kK�䴍y��ON�G��Ҕ$r�z����d���������ʊ��Iԩ�Vp�d3�Z�J�Ed$%�ԑD|�� :�;5#�����5�����s��!2fV����JՈة�sn`Y]*�^-"��Y�F^&���n6[G(����X�XS����!�`��F��Ag��NL�a&yA����!���yH�G�h>��XY�����x������3Z�``%BViؒ��G��	�e+U����
0�0�0">�g�4�zB��fq�Á��܄����U;;�Y	QR$�#�]�����{>����h���_L��MJ08=�t��g�&����99(��﫾�r|�jZ�ʄ,�b�/&��GggN���ffh�/��5��t�1R<������LB��"�h�Z(�KҁbeE��j1Z"���Bh����X�թ�b�R�K��!4||F��^\O�+"�u;S���^M6�z�^K'�n8����}���������Z��Up�Oz��+7�L~���{;�K����V.n;[Ӂd��{��5��,���T�U�6ױ,�2��E���&�h��o��*v)�x��{Z��v��V�޹^�]o�k{R�����3�fgs�������33���t���陙��|�ywwt���t>]<���ff{:.�]��33=�����Q�}M�)�*�
j��k��e`3t��)�rvH�(�+�wͣ�Q[�^"�&!���`���*�ժ��*!@���]ъ�l�*zM����Y���~0p;��|���b1K��$g���>�}X�4N�F2������2�: L@Ng��Ȑ��s6�0ZM��m�F�Q_�3�'z�]c̊k�:��0%��.����k)�+n�3CJ�R�kf��m4�rv@�+�Q��[MDƸ�[K��o�'f>Ǉѣ���A�������9�	���X`�s��a�e`��o34��ˏ�@.�+S���0~K��w�;�VϜ��j�J�
:&�N��&�62���G�JMsKH��ٰ�o��|��d�a`���}��]>{Ӯ�u2
�V���h�|��e���涱7s&�J���Tx��#\���C�	���d�2ᰯ���EHh7ޓ~�:���IR¦fy�ӕ�1�*��bZ���1�'�o5��`ж��}Ĝ'"��Ĳg%ϻ.fe��k���d�K|��{��ku�T�`Q�2C�>�±��m�Đ�} sFr�s}��m��#mBB$Q�.u-�I�8$�,�32Xjs"���C��x'U��iɚ�2H����w3���U�T�`Q�2A�����쟕W���/�o�C�y��ͮ�fĴь�M�j�cT�f�ff�A�Ic�tbY �NHH��%M��h�~�/�LF���	`��,�Od�XXn�\՘�f�E4w�&�cd�n(TZ����A����6�[F{8��
>&H[�J��tu��7Xd5��&K�,(>���B�\_^��|���0���m��p\,'���5����w�e�S�V��K�+u�*T0(�� ���u\ς�^�DKy=���|��w�ۿ�ջ��ܷ{T���L�W�U.˼�=��<�k�58Y�,=���_}��H���&C�a;+%!�.�X%J�$!#�B*)lJb�
�hu�$ h��4E�VJ��YN�,rdC i#}���8���zt1�2'�G��HF��zWr��+��M��H���?��$�	�y�$�I$"��QG�}��>��͘?�	>ӱ���HC�(��h(�) L�/���.&t\o2JQD1C�+h�;�P� � �T �@ �T �U�@��`�  0 ��B`1V	`�X0F�`�A
P � �B�`�X0V�7t!h�``
`� �b�`��%b!(`	b*��$A�$ �"b�(A��(�$
�%!DB��	.�q"�����$bD�%$%E�#1#)]�%�A#1"$A"$@H�JA( �?��`�`���D�W�ES	0�,1"	�$R ��##%!
���H�E"	H���PH�"	�F$A"	IB@��B1"D�$bF$bD# ����HĈ	H��# ��Hĉ1#1 ��HĈ$A"	$A#"D�$A# �"E"D�$bR1#1# ��"	HȁHĈ$bF$A"	�`E�B����c���@�$bF$bD1#�H�"u(�$bF$bD2$A#11"	�H�"	$A#"	�1�`Ń`�2$bF! ��bH(2 ���1AA$��H�# ���� D ��Hȑ�H�F$bA"	H�F$bF$@H��% D1"	���H�D ����1"$F0A�0c1�0A �d�0A� �AA� � �A� �`��1$�A �Ȃ��A$PPA Đ`����A�B(( �A� � � �� ��$IB��
AAH� �DI�	A�1 �A� �	Pb	A�1� � � �1A"B �D ��$@H�	 �	A�DA$"$@P`�" �H1Pb$""  � � �A� �� �b� ��A� ��	 � ��@AA$ �$E"(� ���"�H ��"�� ���b1F#F�`�DDDRAD���H� � �1�""�2!"�H�A �D � � � ��HP �E��P �  � �E�F@!! !�!B@B $!"$����B�B(�1C����{f���zhJE	��>ƑQ�$	HE3;RWzO�_����ï���'��S�`y��_��ϙ�������w���,�$1|2������MwHw�v/;��zＳ{=��?���S�;�|=9���Gp������}��>ϴ�A�`}���~a��0DDC�B�Y@��}�w��0~�������J��������tG��B���!� >3���O�}4�ㄐ2�����>%��f�����M�����jq��i�k٭q�G=��̭O%�S�,�C���ފb���P��& 

�iB"yE."*\TC��Q*(��a�#kL㺷����=�nS��N���>`�`
,�,�(��*�)PaIAI~g�=���`�&������֏h��`v�r�0 �f>��?O����>>i(��Rz�K^��/ϯ�<?x�����>�i���8!�J��?w������C�D���@�'xC����<k��W_$�����DDC�}�X�r�~���O�瓃���G�^�� �'���h�_I����>J*�[��;��Fg`�H	F@�G�hTP�Z����%�8�%�DQ
 �����y�d\�C�62������&����T|Ll���k��K�n.����DB��<��$��Ȍ��\���{��(}�R|����w�y��?��A��O�i<��:��+���=�I�>������"'�Q����?�}<�0�"!�R����C�~��DDD8��{�^���������y����;�n��J�$e�g�p`�$�0Yb�·�n�X�����pA{���K=�Mw.�8�@Ȉ�����|�ф��OD�<����v���v���p�;	��C�@��4`2�@���'����O8! �)��<��}�'�ѱA@<�0���_.�o��g��e?���q�*�- 1���������"�(HD����