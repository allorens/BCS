BZh91AY&SYV�G���߀`qc���"� ����bB��    ��m)�i��4� U4V��#CmmI�5��F��B�f�h�J�TSa�IEP�(f�cJ�f�MeSfm�[|u{����5�DZm2%�[cRԍUM��6kEQCT�(fm�h*5��[U���-m�`�"�6U�m�d��3Y4�M�ֶQ�Gs�R��V�m�ٶPյ(�%5i�T�-mZeY�j��٣k[֚i���Kml�E�R�ZQQf̃E�J[5m���Yd�-"�����uY*՘   ]�s���me:��4��*����r:�T�cU��浫ZUw;��kE:�N�����n���iU���z��Z.�f��9��*̶�U�R�F�i��   �
�S���=�7�����nz�(h<p�R�������xzz��Ct�[�2�-�Ǜ�h�4��C�����:��{UR��"y�U#mXM[j�k*U|   ��|��v�Kr�]�+{
v�O8Uy2�z�Ǯ�Y]	y���ץ:j�n�<��PS���i;miiA��}��z�3��{�>��{i�i�97�)S֟}��e�f��j��0��jp  ;��Mi���U����m5���n����/�S ����j�k�>��)�T�z0w��n�Jwzmw�Me{5�Y������ܭ4��z�v��ͽ��/u{T�Z1�m[$Bə��  ;��|)T_d�|�������U�*����W��N��ֽ��ޟB�4S�|ϼ��im�f�|��_m��[�u}�_{�P���;��K��9S����>F���U��Z��0TU�6��  wm�����ϗ)��kJi�[זƖۻ�79��b�i[��W�i�M�q׫�����^��T�Rܣ�^�l�ҩ/J��p���S=��f�բ(U*-��M�  �o��W�����{p�zeU�U��5�:��7z�(������-m�����w{T�Y"o��i�����  L�� :�  ̮����Z���ZԬ�L�   }��J���NPz�FC@F�w������t
]g���twu�@�G�̸ (LX�:s��נ����ةj%���e�KkY�� n��v���u�  ���S@�{� 9��@�^��7m�tq@��\��� �޶p ��ӭM�6b��K�EV��  v<_C����op4�����i΀�/^��4 ���� ޯ+�B��q��]8 �      � ʔ�C &�� d�"���* �    �~LBR��d      j��@��� 4ɀM2 ��@
�CC   d   BJP55<��4L���M=OQ��Sȏ�?�C�f�C�?�O�����3�0�YH�3X�w�������1�����xx ��>L�π
�¨*~�TW� @��?������?� *��x����PW��%O�T_o��?��{?������?FQ�6�a}�_v݁�d}��d~X_����f�+����dL�����c�)2>�L����=2����)����+����e}0���/�����a}2��/��za}0�>�������d~L���#�����za}0��L��Gݑ���e}2��|`=2�W� zaL!�> �ʀ{2>� OL��Q�(��@�`=0��QL"�OA=2��QL*�A����e=0(��T̂��L���L
��L���L��L���� =2*�a���ze =0��U}0��d =0 �@=0 L(�QC�����z`T=0��OL�ʨzeTL��0���G� ��D���zaD}0>�_L*��T�aU�Ȉ��L*������ �� �d@}2>�L*�TG�(���z`E}0�<�dD=2'��L)�=0'�����S���3
zaOL	�=0��a>�S�>�S�=�S�>�0}0��*z`_L�=2�'��Ȟ��T�Ȟ���� �{�W������@���q	a���p���"eȼ�o/�hw�Un\��w�[x�`�m�������y0a�zkq�k�WP٠�'�]��4M�Q�4��B�xD[q������Re�t�fñ����巩�觪�=�[}����������e�)e!�^�j�3IH7i���ݳ���=`b":6�f0�oj�$�Nj���P��Ȗ,{��FT3 �XY�P�%�����2-��Ö;x�HЊ.��̘6\�� ͣ��3�f���R�Zl����m�9�cY�e���N�^吓�-m�ϥ�J�H1��ժ�o,�ǚ��r.�6fɵt	28��n�ͬ�b���f�%f��2�����m�Պ�+�Xuul���׮�N�ӌ7Ne&��;Q	��v�/-��_:p����n�Va��ۼ@�Y�[Y|�ob�k��\�:5ȱ�����:���^��;�H�8){z2"�8���A�Ӓ*RTK0õ[�e�X.ُi�,ִ&)z�n�0����p��7���˚�Y1˪ �(��ȋ��Уw� ��Ƿ3m=�[�r􅂤�+�[���I�Li�W�����ܬy�3@���Ä[�fL��i��k//�5-mا����q`���^���a)�O)�{B��[��/�:.����iJr<�T�Lo5d�"�bVp0S/>�ͳ��go�Ո1Lު�owf^����e�:nkg��$�E��|�=��@ր,�X�I`�y��ʗ��+v��j�CJВ�j��Z�X�~J���T�6QW#���A2�`�-��5���A�j���j3YsYJb���i�2@��b[�6h��ae�D�E롓6�]��5[yF\�tn|�UC��U3,���ɩM0��6���서�.�V����4��p�κʸ�Pd��Dcn�
���g����6�܊�
N,���w��Vr��/]�Y,��t�6���}����Aެ���aw�OwHx^S��a��/m�F|иf���GX����2�k3vm�qޕl�f-�5p���׮�j�Y�&���|e�;)�v(���mo��rԩY	�ǀ�J8Ҵ�h����X���-�]�m�R6�,n�C�Ѡ��L��o����]�;�]`I]�i�9&eTyt�y6��*�/T0;hh[fU!3{��+���!�.��Q���)D439@��p�SyN���7�27!����%2�����.��^�sK��I"��n�f�m���ʂ �{�61�6���
{diʒ,E�b �dʒ�X�7aܡO���[�5e�eڲhl��hT��/u[�Ң�7W�P���6�X Y0�نޔ4K�S-��]쬨���P�(-�{�b&Q�5b�N�隯]�;*r�â�%
�fܢ�=��kA�����(H�SVe�-5��.��r�)��e�<����;T��8~Z
�U��cm�x�8�54��8���K�R��`ckJ�����ʋHͤC+6�n�9�9�����:�݈�DVnƈ����0�vf�Q�Or�*�#�L±�Z����+n?i�̬���姑�.5�Y��k&̩��jHJY��h|Y�Y�\�`sn��\f˘e���&�ת����`��JJ�H�1v�sZ9mSgׇK�Of)q��Z㕑��M�ՑM6tk�x����mik�)����gM�s�Hݼ9.�x�f:����"�.�2��M;1^\y���mm^���Q�� ��ne���I���Σh]] ��t�H�[�C }F�1;�]k�њ��>��)^�h4�a��Vr�{�d�W4 ��46�;����	�[��3sPw.��2�ƒ��"�L��4�%i7zD�Ն�2n[Ɇ��n�:�;��:i�M�%��8���]K�r�JWK/��#�,�#� 3��&:�d�Ö�nS��Ffj�!�Ԃ�Zբ���:�V!&@��/	ٟI�GJe�a�ʏkr��^�_G�Ⱥg-�z��`⧏R�i2�<ƴ�F��m�.���V�꾅�܁�nP�0�a=��l$ܯ׍Ҽ�1��n����D�R-1��(֊��1�)�-�7n8X`GJ�XIiv���
��w��w�f�/i�Z^b8�k�R�
�i%���Mώ�X�IZh _y����`���Fe����W5���PT�H��I$楅�)f�,��4�>��j�of�z��8�jv��ȀuHQ���ϝDĂPP�;��b��
��ُ��,;aޡOQ2��.h�L]2B�0�7�6������H�Է)�l�T��[{Q�)+���%��w�~��(f
�WQ`�k]e�:o��ʶ�梘�ղ�j�M�kbiv=��6����Wu�u`�����05nn�M���ݛ܇0nmJ��Fi����-~�ᖃ��)k��^�d٢�016E�/v��� ��tŸU��dcn�&憻:�~�w��8Y���촴=k\Mf�"��M�b�UX�[պ����ٖ�f�6d�v�����ӍO�AY�rb�j5���J7� ��Ue����ݤ7��*�K ��֋���q�σ�ź:�l���e���=o�7dJ�O�^�}�b���P�Z�i�V� o5���P|��KM�0E����/oeq���	De�/(��;T,�!Pĺ�!Wa����N �v`��[B�T�Cy0��К�6����A�&�]0Xn�mX�������E�O.MQ�v%L{o4���� �����c���,V��Å,y��c¯�vхPK]�Sn,6�4fc
�JiV���n9B�h�;R��eh	TU�u�|S�[-m��'�W<�2e�z3.��y�ђ�i*��Ad�,V��Ll��j�-Vb�r1�(�T)S@�Bc��Ll��VЊz��x>��@!Y1T/6�L1���zPe�b�6Ӣ���8�c��+p�לx�4݀!Ew-	�����.���Ŕ��oJE]v�i��ym�.g����v��$�E^�`5R�w��ݐ���X��n*ե��=ФJéq=J\�7iޤ����[O��22-����0[�y�Yf�o
]O��w�(�Z�6���.&�ʻנ��gm��,�.���{�VX�P�ϩ�z���
^�L�X��_4��M��u6��1�Ɋ%�.�7���:o5�
�R(Ki�Znf��:a��ȶHͫg*�j �7494��tP5�c/5*v���%$��6v�4��Ӯ�8����e�91f!�x0��Owe�\(8,rQ*J:�;I֩�n�,�n&[G�̻2�Ī^���R^�zP�K��
�{@�^���;C�i��$mk����i�ҍ*�`� �&��\!�]�tuσ8�ug&�O�3UJ4����A��A�O]�H�����Hw"�o>X��S��F*	�쵄nB�T�h6H�m�I�U���J���U�]�;x�J:����ަ���w]ǚ�0��*�V��0L��wkCn�Uh�Sn�Bj���YY ;`�֞�:p+�z��uX�z��F'�ҳ5�vӲ��j4�$�O�%�M�K&S4
��E�﷋����E�.xn�,�渐v�[��"���V��R�{���
PD�vM
u�`�Ԋ�� �=u�YCb��,eK����;�d���ՠ33���6(��\����2D)���{JQ��j�Q���+E�n��3��a�6�ű�1�;9gn]��5d�� ���˟Kv�n�B�KX���	�t�-L����X���{��-T��8lK!n���Yj��h?���
P�ҷNdM	��l蝼;���73%���hV�e�Kd���4m�(��[v@f,ٺ���b�SoV�J(.�C3lh�6��2�Pz�&�g�z�%jw)�T�+���Y��ݨDlf�Qwj��˧��0�.k�.�y�cMZ˴"-�B!	�Q�ndzS!&�^9�͑��U�CWeQt0kK- ��N=�S �ص�7O��@s$8ւq���ݹ��j�L�u#��)�4C�<�z!���!�t�����s뗩:0M����w�1�D��GK7M5E�lx�u����I�XS[he�/Mѭ��Ze�w����n�l����ҜB�LG�)�"Fe`��a��j���.�Ný��ܩ�	I˛@��ݭ�jX[�A� ��Q���FQ�E�em1���d[Fɢ^�܍8Q2�4��n�4�{X��F^���Z�����ꎶ�.�bwv�j��;b9f2�ťeɣF�6ŭ�K(�a��&�OF�U��-gV�H=��h�0d�ܘ �-#Om�b���eM���j�I�%iL��h5��oWZ��Ӓ���2���T��v�E����ۻS�!�Y�`:j^�Y�m�q�JZ��m�1��r�J����=�՝�x�n�T��!ց�r��' �W��o.?����j̉H4 p�«6�n����h��wA����p���s.Ku���,c^�6��M!D/h#��ft�z�]�Q��~z�#�٪��(�MXl�E�6\6�+րe�aEQ�c�-;�6	��,�Y����B�o�!�%�^���k��A�W".��f�	X6��\ 1ݺ��	û��z� %㱖0:�VllV�����e�lE�rY1�[��#3e`J,�i`х5z�U%�ŏLT���b��5�m���mQW�\�����6�F�SA���Ҕ�Z����к���'��y�e��S�h-�W��V��&����� V��R�4EJm�r+�ы:x X1lA�˽�E䲴�V*��/"ǥ�mJݶ�2,�F �[�T�E��x4`�J
����G���e^P�Za�d���HL�V�iR���=��LfQ�[��i\.�c֛���f<�Pa[�t8��7LY;T�jiٻe�����q��޳�A���Lt�$���$�jْ�Yr�R�S��MB��
`�����RJ��m�-�N�N
���K�x�^ ���XDK��fCEV	��2�a�NL���Z.:t,T�S�2buR)��8�8Ҕ�Rق�j陠�;D��C�0gr�W���8K!�XBA�[��[�%�,�0*��W��Em�#�nVKb���z#������U|�*g�C���7˹�R�WB�)m)��"܉����b$������bL����_c�쌉�Of]�R��7�V��Uj�sZt�(LE��q"��N1[-͈	U�n�`����uM6E6�M�Zȩm�G B�L7J���Y��D4d��Q�n�N�g�]O{�����	�tn홡�u����ȭ�vi���ԧ2=�&#@Q�g]��WU��u��}��k1����x�\Ȧ��`>�n�7z#�EkA6�˱�FxL�C&a�ö�����E�nQ&c:7E:6��NE*ޫ�j'in
�*L����ek�u<zм�{n�1f���e��+5�/#@���ـ�ۨ�������'2��p�XCb%ͩn�J��i��x���`Wr�NQ�+��TcUn\�`�2^d��-�ˁ�C�X��S&O�z!k"�P:3)~�qX�*[��7�Y�L���jL��v6����h�Su�Jb	Ү�ё+ܐ[�Ha����`(T7t�N��emn:mRT��r<f�WÞ>�u��3�He�n���HVA�!1<ë7nT��L��M����l�t�h���%є�hgF�#
��=J�V�D�]e����d�����욖��J35ӎ5X��J��I40��R�Z�o%�ƷV�-�.����0��+vˑ��#��yvuևUkA���t�D�줝�!nήW[�I���81h:�sj(0����2�a81�6[��.eaosMׯ!zym�ɥ=�ջ{��4c�3hf:0.��*���i�o���r*��(jg[t�ɢ�#�aaE�ɩ��"tTe3%p����{;���R�8��u��鷵���ѣkbCpi�Vz��l1E֜Ѷ	�T�6KT� d�-LQ�^^^�o/"7`׻�n��CN�^��VUhr�ŀ��w�r�4���_��x�V��9v��,��op��wNL�7XEU�T�v%��=�{�*ʭ��aTr�	k�P�ĕ��ѡ1�F���0��h�˙�,`��^��$m��Eܺ�Ck2�J�	�Y�ۯŰꞡF��ҷE{H�x�xx�д/.n��kIw$�m�E1�UL.�mcojm�/T����S(j[Mmn�T(37wB�H1�ݺ�����3���aBղ��OoQ���PX�]���Z�W����j��P1��G�i�+h�W0����婝a!�3P�����[���$��Rc��T+p��6ua) h��޻4�Y�y:���nKi�3����Q�/��Q涻iQ��kibޝK�sK��sT�+���e�\[��H��f8S*�MR�j�����q��&�]b/d�z,�ؖ+ �C��|�����U��-��)�WM���;��4XY�D�r�\9JBK�wm��YvƗ����b7W)�te2Sv%i��˸p�&ۻ� w�yB��˂��u�X���N����"�v
Ě{��MX	Z��,�wM&�u8�(�����bVd|��h})�t�1�r�d]!�`E�2M��k06 (Lb��I	��cj*�
�X�-ł�*�k�y���] �7
aR!X�t{ذy-6-7R�ƣhdX�c,� �%�a�i	 W�r\�  �ٚ\3�k-f��$�ÖB"��굣 �<��	.\*��^�� �
����\�-�h�{	�l��ۘ�Qn�`���DEϽ�s�Ǣ[8-��#��~{�c��o?���X>�
���_��u����D�����`���VA�(���U:�;6�j�o�7-2��j5T���q��h[�N��e��JXC^0�,m����A��;�GΨF8A�H��}'����[z���?i����Z��+�ة&!?a6]C�Ǥۿ�8n`�d72k"��	w�ɯj\ui��f��Q�Y�<XK�f��Z��Y\��Q���
"���U`щ���]�����K.�͢��SrF���������f�v[�V�ۮ�E+�ފ|���a+r��?�P�y:��)C��ѹ�c�;����`�bn�
�yB��%-7��}��Y�\�R�4�t�÷Kih�x�x��͘����L�$�մ^ɏ�y����Rp����M�WĜ<��c^�h�t��eD̄����*;|���'��aK{����NYG���6����5�G�����"��:h���-� <��RW��%r�ٔe���H=�r�=�2%^+d��O~�8m�R��T��Z�{7�xC�@�#.����9,K� ���d��
����&�.+Ia�\0�t��L

RrT�q���@�,�uM`"�w_W_w4�V�G6�8&�.��5���Z�k��fj8u>ӻt�^oIt�Ea� ���s4h�����T���-�|PW��f+O
�]�KI���Ťp�1�����bܧrh�1�5c��ܥ:��/:%)JV�\x�ގ��e�s/�U���Jf�.����_"fK1v���v��+R�w�)�ih��C7�b�>�l�WX��0Z�9�C��<Bw.&�_e+�[�t�R7�o�'�;V�n��q=:	�ұ�OHrݛ{s�2�k���<9C�48\j�#�N�3}H����]�x���<�rb�6PoG=��Ʌ��¼��N�h�l%:��9l�tg~"��*�1�_eɋ����&:�t�t1d��A�;��n��jz7����қ9��ܲd���f�vPy�ᠲ��c��vP�)� �J��m5es��.��!Ӕ�������P�c_P1>�88�_)�^��w�S+iaK��a��j �騥Z�F-��EJ�un������(K���Pf>oJ��h���b`�,N��I
�K�ɟ��{�?�u�{�>�s8�AӢ��.��-�k.�5�����ß^X�w��a".m,k�Gw���r�vh:T�[�I��S�:(�R|��TI�,@�ҙq�=�WN�I���F�Zn���e!���W	�8v��F�8����
4�M̋�[�T�E�V���4c�>��V}}2��t3��_`�jw��y�$7ᖝa�Ԝ����J[�=��ioSh���(���)Qj�B�9����@n�m�X����T)��:j�Zޥ6�n�(V�[7�\y�oU�ǩ�Јm�l]�)+�N�lY1��o5��O��S*dw(7+$�{�H\C��r��ƺ'R�&�]/0Zy�&٨h.��Đpj؞\fƜ��/�c�a������NOn�5�o��&�k�un�e�b?�����e�ZU��8��	����ջ�ҥլHW�N��3d61���>C�VS5ܯD���#�I��Z�ϕ���M�A�'�T/)�M[[�3�^�D�q7��Ul�,+&�I�¨�[��c@�\֦I�:��\�(���Ȍ��+;�t�3�Q���y����N�%eou�S~4��36�v�>��vΆT��\�4.�˫_+<���B�[�&t�nA����!�Dk#�ES�cG$BV*���2p2����L��{��"���=JD�!-�<� %R'���n 1t�\kr�WVo	P�Eǝ���=��lJ}z��b[��qF�U<�DG�}�y���h
d���*��Zٹ|�U��Z�"Тm�径n{{5��J�O!_u�pI0�X�Ʀ��ugp�c�)�=�DT�Ul��g��2^�"S���ϒ{Y;�������[��C(���N�I�&�e�L�lna�etgi��;p��u1rZQ����}4��FVԤ�iӭrE
8n���r��em��]ݜŧ���莁�i�9]CUou{:�O�!���ovX��C�iby�?��r���ͮKބK+�7Y��vI�E���?=f:�x�����P�Cz�[�/PF��_�C5nTcǼ��1�ź�Ď�HT9՝إމ|*}J�q�Ŋ"y�ꖇ��n+Jg��SGP��U����{���-�BV�[�N��]�96a]�a����T�2hc���r�2=����3C�dd�=Z�]8MQ��s};h��Լ��N�8T��'0E�|��k	�S[�J�\�oo #�-�:���ޛC&]<��>���'%�P32v$S,�!qܢ�������Go���4#��ФT�x��N�"�|�:Y�l<�(���7Ի���;Jǯ��Rxb��N��u�k9`ג��R��
�~"���Li��A5�#�F��6B�7W�j�jG�>�hC��_4wY�IgMU{�!���k��i(���N=+e�qa��b�ult�1��؈U�Q�ji1a�;�o+�C��F��Ѝh�y���ݹ�.a�a΍obeۼ�F��c�uh��U�֓n�)���6��f���z��������]��A��V2	KNՒ� NGӲn �?{�p�`���3:p�IKλ:d�O>ʾ�v��G��%�Ǹn��b�2R�S��wv!Q}�����l��s(�.8�j�:r�˸��&b�OY�D��H��ܮ������)�!,��	����3����׼����Wo���mn�)5J|��"w�ayX]h8�]�t�f��Kй�x����h��5����C�3���@�gme(�9_�t})q*M�g7)1z��+�Ά��_u2����Y�j�y@e᡻�1�;��V��Y �*/��v�����U%b�`V<ޕ���O-��w/-Q�@�s�
>�Ŝ�%�2��5ޙ�v8�s*u�0��[����s��Oɷ�`9,4;��U%\���urD���y(^�͜r)�õ�7���rל�١q"����L·6Q���ڝÏ��λ^Z}���b����`R|6=J;����j= |�<W^����\����^��
��SQ�dt�������jn�"��Y�V,�w]旔\b�$�[�e+���\)����Ri��j��ކ^nl��q����&��T���ѫ/�YU���%(0��t@Ȱ �H��e��u���r6 nR�/�i.�_0��#Ris��˅�����(���s�Rƻ,��fǗ"�i�T�0��]d}IQ}��������W�fW)v_i�Dj!Jy��th\<x�ۼ�V�����i�I���y{tɥh/"S0�xn�mk]S�q�s��]+d�[��d�"Ý�X�*
��F]�KFJ4�o�e�c�'+UַZ���;z7��4C�n�2� i��u�*����՛�F����2�^g�u*��Y[�lW>��V���B
O�<����I.�ܜ���r��vo2���[ף�������no=�юٙ�4�G9��w�l�:�αI8��YJ�6�9:��Kɦ��yg>�Y)�s�l�|����E=�:�P�#|M��M*wLjP� !YCA�qAH�����S*ΨH�W�1k�Id�n���K�(�Y�vQ�>�J�x�l���p��.���fkV�J�qU˃/�Y�t��U65Κ3�,ƆD'c��T��2Ŋ�S9�X�RIٌ��n�jʽ�ȥ�Z�y�HU
㎷"û3��*�fq������[�h>Nty�c;(����'�ck7AU�Z�J��j��h氭I<ٔ��H��f�ˠ\��捼�57�^���.�*�N��$tu�>2@5	�6��J�̘�e+���R�KL��ޱ��n\�Eᾼ�X����*s���[��5���=��+� 	[�j�Uuj��}�*�صR�eC���=����[�a������N�`{Qv��ם�'6�ӐV��mw6T���Ğ{Z�v�
ɤ9�%1W1U��ki��rh�]�V��i�Q��ڭz;��u�$^h}Z�u���ǻ]��U�qq�=�tqp�M1��N;���)Zɕ�f)���fRN�����]FH#6��1�O.��(����u(��]m�A�{�N]<�'!����c�<�/�"\�,\ӳ�=+H�qaT�f+ީA�Q�^��u{�N(s��$���	�H_\��Ι���?����/Dn��y���A�[�x���ݝRw���-��YTJ&v�n
u���v���[��%G�Q�8���:e�߯2�_I�j�rA�o�Q
cE]�>��o��Zoz"�6mӪ;5b���K�݆��O��
r����A�k:���h�だ�ktwݑ��ݡf�V@֍����[̗\co���}4B�Λ�k����8��2�����\���!�0n9|���ᙆ�No�N�ɴ1���6��h�c��Ơ�b�ό1RU�Ck��'1c���Ĭծ�>)��g�H���:�-۾7c��t���Ի3�|�%W@>��ya�ػ���1A��f�{�,n*�+��J?���k#2uD�$�x/jnq�D���Yr��=ܕ��mu���+�4UV�J��h{�³�{�n>���[aU��F&���'�D�r�
�}�v�Z8f#��Њ�|��\�Ɲ��VIsD9R��+�
�evm��V�yw'�+�E����1��i�˳���-��5��Ā��g�@�IE�wuܺ��6X�&61]lJ���uy. �7;Z���}��xi�v�FB˻��=�6�F�X&�K�P��aA�{��+{�^P�r���2�f��z��щˬ�����{bq];�s��vʞuC\V.�l3F�Q�o)4WQ�:C)�dY����y 7��s�(޾�gr ���ܟ)ػ+��+��$F�?�l�
���Qs�p�%�U��m�äJE_C}X6�3}�f�%�Zp��J�z���^D���w,�y�@*�����9xyX�� 馻78�ʕ�������ݤwj�K�V�pm�LW���_u�@ Uj�ɷV�.���f�b���U��E�7��M层�*��	�xb����t�A`ˮ�¶ED"t$"�e����	����R���g3&�R�������`�|�#�)o�73F�mM�8�_bQv��Ǎ�h�[BM��V�z�tn�wۥ�2S���c��ӻ=
�E������֔B��+
�cd:��i,%>��u��k�U�`�Jp���;X
����T�T1�P۹|�tR�3A�Y��2���hۉLv�ZQ���NK×͸!�D�u�Cr�.Q�|oK7�A��MC����v@F�sT�T�W���w�vZ�j�;V��2��VM;\��(r╣�wj�@�-m*��k �Ɍg�ƹ�Y젻&;�X@D��s��Qo��ǘ�lNȩ�w���VNu������{l����7!Ֆ⫼bi}#�}�N)H���iu���v������4������w�2;a��ۗ�VoS� 2��ʲ�m��3~�m��O�Щ]j�����Yʲ�T�η�E��t#k�j��l�N�=fs�α�@�G.^�vzS�蹃a�햖l.��ӳźۜ�ވy��%��W�\�.���P5����L��Ů�f�5�yw�:>��b�A�:��O��M��w�:(p�%Y�Y������7%��1�.t��[A�I}�ș�9b��&_g�a�$A�ެ���Rem�u��]�Jи����Aer��V8�|���i�K�٧������]��w*Qu1{����В��s-��Ys&c#~�`+(�zJ�V�锠FE�kZ����r��y���v�:r܉ho��Qf�T�Z��E26�Ǖ ���gi7�΍��P�va�o_;!j"��k�ӱw�^N�ׯ�-]�hTn�̊���)�{H<�qA��V.�=��67�-JC�E���3��Q�ܽ��YS�eo1|2�-���Ѧ�*C�y���"{D��c��b�nAW�=���F���\(I���cXֶ;�O(n��>��u���=��c�D���ν�$��-�B� ;����٘jvm^9͵0�حEHwfj��� X�r�֝�s!��iZ/0I��kKF����y�/��p�1��S�������-���c<��ݾ���)3�R�����r���@��m��f�Dٝ��HլX���$�tU�J�a�Z[�6Ÿ4W<b��Y�x#�Yec�5�I�8�ou�뱁���<Jż�s!��t=O����t@y{�����I���IP��5�^��jV�o�]e�K���/L̷V����I�9P
���l�������=��$��YVYu1�ʔ�U�((�ݤ��Ҷ�r��X��)�k�{8c�9}���\s�����c�D� �E�N�����u`��������QY�:ˡ;�w �����9;� ����ո�bh��wSF]��ï��j둕�^Q�{Wh"^%���z��ݬ�[�S�C�.p |3O\9PUAv�:6�+��Cz�y�!�x�M@�� v��C-r+��JuI2
�Ö0:��-���7�&۝��4z����������C��M*�S�2�r67��2�p�-Ȥu6F�WE$��MYm�gaqϻ�T�	Nu�{6E#EsJAU뭿��ﾗ�]��'�!�{A�U����o��7��G��������X��=��i|�O6N��8��T������Ŷ����=�Jk�D��� z�����>�{�|��!��
���_�����P ��}�������>�_����={��?�������u���Uɾ�	(Aۚ��7+@�}�ъj=�o$~����8���ïZ����;��!0��� w��ןc������Q����0^�8����.����ͨK��N֞T�Q��wU�Ŕ��+v����s}mi� @�]	�V���(VsF�\��vڎ������.I�,�P^��� ����f��&�.m�q���tƖ]�C$
b����� �.*@"�=������kq�BE�Gz�����V(���9�n�&�lȊY�s�^peއ}���)4�b��)����t�d��.=65{,�5�ty���@���kכ@BoY��6�굇7�<�B�
*%抾���*Dg=s�����5+�s�sV�>&�ܒp�f��ee�AL�9��E���oN��:!�0}�0;��@�x1R�� 9Ќ�ˣ��6ʫ�7m��X�e&/�6u��*ou�Ҙ����.Y]1�lt�lt%r�ؖE�
�n��	���ܡs��s�?��1��4y)4�d�:J!�����uۀ��rr�I�dp��݂�{!��X�� �꥕tN6+j�����@�Zܧ�+�v3j�%\K�D��%E-���H��Ϥ|��
7�q]��7E��ŕ����v�V�s�
���䯏p3�m8�JP���Q��Vc����ѻ@�Z��3j��
�f�ǖ(t�6\n%ݭW-p|\]7�:-�i� ��b�Y��F�[�בq�#�F�4�ͻk�n��f�����mګ����R�6v�CtS���ՠ��h롟:��:�ﰹi�v�X��O|�v*=���Nͱϱaׇ%5)k7I�@x���Wkg[p��c��jM�ç�U[Hu*�Rj�F��H����F�Gfڻw�yY��CZ�L��Ba����ꇅӽ��7b�uty�Ej���v%V�e��n���[�b�'Z���;�V+1'Y����q�:�]��mp3m2X%�Q2�	uY ����Hg-MtwDn�(n��n\5(u����J��	g���W�U��ڷVFL�[N��V^�����md��Y�$��1]�^T���ǹ�����z.��m��-���*q۬�	m��@��z&�"O��{;-T�1���5�CCR4^�y4^i�;kr)�A�o�FT�X��kf8�_ִ,��t��WK��:����Q�����+��"C�~��cX�K��;��d4��w: ��(Ѐ3�:�(m�P���=/Uu��-?��̈́���R6����r�8�J�&X�lV����vio�@��p�m�[[�T3e����8��,M�#��r���ݔ�%#��q0�մw.7O�c�ޜ��X~}M�J�T'�y-eG�֢���v	x8���s��ek��j�G3��εtyQqm6��X�����F��#�VH�$��2�1.�a)�BJ�ĕkK��*��zW`ku����Ɍ��r}C�����f�`d�r�i�u:���I\uٴC�\��d&��u��u�I��E+�����Js[-�4�=hr���|�df�����%=���\����M�|��&\�6�3�q,�ʣ[�N�717m�?8�6V��vճ���&cޭ�ΡW�X�Qm��B��d�k-�ځh�HդY{X�n���ߪ�]�/��O�`�=���P\����ֺ[*��K���In�%��n�Di�$�R�����k�6��[��-v���A�'�2<Z��/�ƝڰO.�2c/V�'(�П><M�BҊZ�h���7^�֓��t��d�\�4��v�R��}�v�o盲�/`� �b<�nw\���/�q�(�/_^�v��=\P��@%��x�awr�ղ�bu�Pv���(�PE�%�r������Ք�1��C`Txm:t�oN
8�P��#@����Cr���(]�k�p,�q����%BIg��fI&lK���d��>g9҃*Q���b���|ˠ���2���T���k̴,cw��&t��񖲎c��wK%Y,fU`�h�꾷H�Z��>Y��P���&�����3�TзR,�B�U�����6k�pL�s�'l��@�_�%t�}������<&�����kw|�e>M	����fv��M�=6[�_ �.+H��Sw4C���h�]�9Ep�z���̆��Al�r��4[B���X	�-i[2^9�"Ќy����&
-���K77�GL�4��rjI��l��k ���mR��)���crȰ�M�2��:6+�峝R\�v7��s�F�Q;ʐ�k '�P���2�V�ը�因�RI�ݓT`7��8,���iX=NocB$��ouu��Ӥx�T���[[j�N�/h�Ǝ��
���m\����L�T��(��֧�xZ��[��nlL^��N�E	OH�Cb۾��m�)�̮��	���N�-�ݑ+$J�:�oX��P�������s�7z����U�mV���&���N�͹�l!���r@䬲4��-Zs5Z���ͮ�V6�����P�#]��-i�rn�%�R,A�WΩ����y) ]t}G���>�����.�Y.��4ӥ�&XRe��y9�i6~uk(輫5���\#3�7Qmʼ���%��pH*��'Y�._HT�N:/;�W<*=#6���̰j
�f�Ly���j��C��:y����*K��Z�N�&a��hw-#��mӆ��ף�U��wV+VW91�d��؛=t�}%�z�u^��Vp饀�Λ`k�њ��W��|��(����rB.o_���}.l�rn:J�p`���c��}|��D#�^:�T���TzD�k��S�0mf���3qs��u�áC��wA|�۳5d��b�a��C.���ԡ5�A��h8un��jJ2�8��C��WnQ�����ӶB�eb�P^)W�|Up|{1Ծ9��hyM�S�*��)����A,q[�J�[ڵh+N�v��3!C��S��K�+:�[�v��Z�n�˺�:T�uӖY��|�A�]J�p�L��f����)�Xn��qvr�RMO1�d�������|��_T���}�Pގ�n���B{hZ"�T/q�8�
w7V�)�$�j��;}�ә.c��^��.�C�כQ"�I�>zlA���X�G'�C�(�����zv����y���ϋ�^�w���y�7����x��|��1wϟp��wP5x�{G�ٗ�vCnV�E^���đ��8�Q��Uy׸+*LA�ё$�'!��8޼T����_\2���ЃˆA*k��O,�`w0�8���)H��SS@37v;t�><)�t��u�CN�}L�F[t�#��1<߇!���ͳ�s�U�6�����3�79���vN<�Q���z3N�mDRMb�em�`�{���74d��O�z��b�AÕ):�J�3�R ��x��!z�=Y�l�MZm��.�ώ�3�s�s/b꫾ٮ��Ǧ� �ZU��f�3�N�n�Ⴏ.�Lzj:AT7\���;pp�Ӏ��9R��Gk U��r�K
��K�s�7Z{� ����̮ *c��5;P�'t��k:Λ������]M9��f����68�£�h5��\n1�9�gjjs�kE���LJ��*��\Y�F���u�y|�V���z��������X�F͍"J��[L.����'��|��.�X������qB7�bqw3)F6qIu�Y)�D�r��� ,<=[�]*%�~����<��ò
�|NS���^��uë����<�7sf��� 㥬^�ua[�LV��.�ۮ��-�%�VF���u��NT��_ZÕz&5E����o���}�����GyG}�V��H�b��&�kZ���2��!Np1O��f�K��og�ZZ3���(�5ΉٺﺲM��mmݴ:�t��1��`$����b��$������4[��\z�����:�$�:��#�E_nXx٠_��_0[������jq�̄�2��z3��F�7ӯd��,��t*�a�5U�2���yR>�4Y7k�bc�I�3����j��J�)��2U�;y�9/Y�M���:9	f8����}�x�F�����V����k;�Uj��L�m�?Y�)�<�;�2�Ϋ�&QŢ�p`;ӑf�nk.u��w3p�8uZi�VM]�����}g|�f!w�]0�ĥt���S;�- V
������r&�WX^	M�}���V��Łt�w3�J�C��r�]���a���ov��i�t�ڤ^k�w*u���"�J�n�/35��T�k5������&#i�����d�v��r�D�d�849��mK���.���՞]��i�e?���:b�W8b�]�f��ʯoNL.��RЍ�Aޝ�+{�%�ƈB_$���U�K3X�T/,����nf*��,oq��Z���z�L"C�n�0,����t�m�T�_Vp|��N�g"k��t2Y	̮���(�ߟ.�tu��1�o��M+�s�sq��OR�f�r����\U�m�x��\L��]�;2�啭�������$����1$[�u���\��)k���
8:��C9̳��m v�ec�n��J���	�j̘��Ӹ���)F�Ո�-��\�XY�(�Y��Fi�3%���s�K㱵r�.�GR���&�{��v(Y4���D��v�aYYOmF�Nxq�ݻ�5����b��s���QÉSW�@�b)6�9�q�x�%k`^��PɨBD�\;$�"�(���kc�"2U�pb��.	�����u�}[W��4�称e��*θAp�U����n)p<�G8�5�ô��ATWջ�Q�a.��(��^��&��Aiu�ƣа��)��;�7b�Kp&��VS�3��;�If����fRIX��TFv59�I�;Vy�W�L!��8�_�ʃӼ.�ڑ)n�m���v���EL���p"S����z�yg)��j�
�(��t����:���鼑Ť@�+ȋ���[En��Q�K,�B��/g
e�M-�[]�8/fn>�I<���e>i �����͛v�Ke���C��Jp[]R��p�*>�)"淜v�h�U�V�twZ���#�2��u i��S8�4�����Y����T�\��.�A�@���+�,u�J,1yI6�M�6����ya\�i��3�+pw.S�����\bͨ7]/}Z�� ��;�u���59���C�a�u��}��������)�Xwb���"0�̠
�'v�#������v�8�t�aY�Jǂ���%7��ֽ�/a�e��\��R������C����JS��$=��a��\�5qkS
�u�=;c��-����o5���u'2�ͷ�WS��7s����C��b[΍'��_�;��l���9&U
���aX{Z_0r7����W_�\�dĂ׵*Tw�X��� q�Q��K��v�G���,��@ʼ,Ѻ�9�������*Q1�on����UgeY��y����:�)k.݇I%Ki	�yR��{��%l�E�����н/�n�2��.��HQ��?)��X�BF̭i��-9�d�tw0%�X梋a$�nvGx�aُ[��א5X��ӝ.�&rŎ~ Zd�C�˔6Ļ�ɛ�$���t[�����v��R��:�t�#ܾJ�y3N��g�IE����y�<�,Y���';+pUa�g]ѡ̆�� ��-�C��q=��n�ZƖ�����2��h�Y��_]�mM�)�;�f�;��_2/Ck�f��Ml�Vn�݂W��Zt_4DƺZ1q�)#K1}|Ƥf&j�ǱcWN;�V+<�Sw����:���1x�/�r�,��z�׶vqW��4[�t�7�i�՗v�3��ۼk���_җe��yc�u�̪��j�sX;Zd��1y,wt:�;�v��� �ũ5��P��r3��%��u�[�F�n�A� ��6�WN�����[�ˡ(�ƑV-�����X�c�)"����D��2�)B��
�+E)Z]׌g��^�VvrZ���g�u����Ԇ�tj	K�vW-<w/�A2�8�$_M��%N����K�;���%n��AdD�9	|�p ��ޱREJ��5u���A` ^{Q�{B)�v��j�f�Ge�jI�2��N�cp|��I��W֑�w�-��D�v�f��3����#j��Wǎ&.ghz����Q$�݁K(�*�\�׋���-�����5���YI<׎6�J.u�̜�Gxjĝmͦ%�Чʌ@B�v4-�q�+N��\�G#�'���I)V�[Pnb�</ji��M;1��+�Z�-�5�S�ͮ)���WbO_%P%9�%��I�S+$��	��;6��j7��'8�b�A�V�v:!6$�lʘ��Hr��
��"1�:K]��ؑ��BY���47c%7C*���'����Ѩf�oc��e`^a6e��iW��c9�Q2Y�QX�f>R,lz���I{�+f��ΩS���k�Eȋ���nn���R�0뿭�ȏL����#��O#�3��/����X��B_хT��/1�|�ሇp�κ�Oc�ya�F���;]ۆ�yU��\j�}rk��� f'��,���.���6s���t& ���șAh���+~���nY�8P�$��A����3z- U��+5���G'X�Q��؊���:2�_L�h�x�4���ݹ�GtlBx旼�bl����4��8�$�ݠ�
|���+-$�7��nk��B�c�� Z��yo6󨘬BU���-�yc_,.�a
qz��/K����˃_3�KW��Nv�1]���z�皧[YVq=�H�H⹭���6!1�]��'F��sc��H]سC��_���� *�Tÿ������_��������G�G�|||||`�?�����=�ؕ�=����X�q(�IP��%���ҍH�3�	���Fc.���q�A�b��P-~Q��?�R�H�T_�b��W�����C���_FbU�e�R��0+�E!�úZx�::�� �4�]�z�#y��-%�+�JӫYX���	}"���|#�!����qtvq̫���9u0���j��2�i�����i��l�i�N�6.}"�����{X�[4�=RU�]V�Oyk5R�Xsn��yB,Jpv=J�1 ��t�wY�wv���X�<c.Z�7�Z�6^2ݙ�������ذ�ݛ��c܇:��h�d-���2A!��>k.V�7�[Ac�&I9���_P}]�epSU\t9@Ǆ�9j�rܵ��A:��F��v��(U�K�G����obҵ�!��4�d^vC���e(T�J��c���@��җrZ�v�]xmN�[��v�47'l͢�Ԧ�!W����e��`������pbF�X�=#��[����p�q�9t�FVҡ�lle��*u(Ӽ��;�]4��8�:ܻ��ta�a���(��u�\�u��"{�:��5�/���oV4W�r��:c��"�h��oH���jrA�|���QF���4H[�C�N�TTs���iT�{��1�\��շ�6Ff=q&t��<��s�+�xpg�'t�H,:�c��m���!{�5�6��(fV�]Y1Қ���[�����{5P܋�[�,$��A��@�i6`(A�@�)��E&���"B� 
��R!"�4�� �����hR)�ɤ���e"��r�L�E:� � DbE"1�"%��O�6`��@�	�H�8�h�'�B��W��j����n�y�^O�GUA�e��A�c�t�
�U�F���KLl�:4�n�t�"6�v�:��(��.���i�(-��N�Pm�M�m�ƥ����v:z1mIM��Aӣv+���t�GIF�"'HQ������O���T��E;lm��n�
�(q��qS�@R��ƚ�ulh1=k��
��Z+E�TD����5A�tf��M1�F�]gMn�������j�Z���������,DUv��E��I�vn�f7mWI6�ڠ��j�m�#�:�D�m��EDh��1�Z��5���QIAZ�F�LM=��=]��g]m`����V�46ΓM�Q]�-;lc8����l�h������������X���F.���s��Em�-M���nƚn�qA������*�ꈨ��,E�h*�) A�	��`�tZDSA��!&�)Wժ+�$��a�]7�h4��7�Y���3��ڸ'���7̺�����3%"㮊��a7�aTמ� K�up򢸩%4$"�4	B �1��f�$���O��G[�{Ewiw������؜�ˡ�4��=^N�����_G����sf�5sR���>��k݇j�7�����M���[I�hz<�x����c��bk�z�@̓t0��7���5����:���Igvt�}8{���ѷ0K\��b�H��w,�=Ǳޟ�m�Ƴ��\]�<��\8�]�z����w�Mg��>��C�q��m������X�w��k�>��g�=���s�B�M$l��=k~�^{Ix4W��yC�z�d����>�zL<^{h���ٮ��Em����{JX��5ޏ��]Wv�at}P`Q֊��~㧁~���^6��ŗ[��c;׋<���O[�"��z�K�8wW%!+�[Sɏux�r�t q���Yȋqq�O���;MP�4���г/*�����������Ϝ��Z|�Ѳv�����&&%%Y
�q����+�Z��Av�� �]*Md�w��r2ڸ���ځ�ypfl�`�ƅ�G�v!GI"[U�x�]�F��4��;F"m� ��[/��ol"�Ɖ�@�N�㛫�����ٓ�2+�*����nYM̧�v7re�����no��0!n^U�M��a[�;��SV�c�DZ�H�w�s^��o>��[�|������]*��f�W�ߍzo��4��#�����OU���t��v���,&�е������x��
��f�&|P�*�����nZm�W�˷���~Ws��?'2-�f�}���{�����sX�r�����������>�Fx{�z��ޓ�:S/�/��z�h��=��i�Kً����>3S��+6:��Q��.p����=<@ŷ��M9�sݓ��w�c���{���C4�k��g7���^�Y�qg�a��1��ÔUF�����������3s��F���u�ߪ��>3g���I{0y�������1.7N8;ܮ^��a�S���C�J�D�{�����;w�cUѦ����� �JX���57:Bd�����p۞Ж]�Ky�w���"����:�(9�azn'�{��!���H�_�s�	0=��W�<�+��/�!��g띭/���m��f�rL��O�/���o�p��=1a��l�[ց
��T��H��$x���r�q4��74�f_���kt�ۧ��;>Y�ci��k/|
��5�\6�/9�N�
OOzߕ��Ǖ����~y2=���^l�~|J�xgX��jk�����J�⫣��8}��:w]�OB���,V,ߗ^_{�n��w�f?N�yA���y������Tˉ�wt]���ߤ���'f��T�*W�38m�F���sf��"�k��C\��zv����A���6k�FL$���UE����G�Ix�u'&�<F�5�3f����S���ik��k����R>G��;G֮���vT�b�ٴ`���N�uOo��2br�8X�2�<r�ы,�edV9�����Ĝ����I���N֎zj�i��w9��^��K��O���t�-U���~����|;6��iO��*�d>��x�е|���K����m�:4%Y�Ykq�x���^\��ӻ��.�A93:��:��o n��^<g�w��w���5�g�}*S��'�v�_~�s�������7��*$�m�A�p�MafҚ:�ܲp�ګ��mm��v�f;:ڶ��է]���T��9{n���֡9Qf�y�Ů���"ds8O�{|'QP�9^���Z���� i���%��qaM{$狷'�b:���^���E�E�4�<[����3<����u�wO���o�PwV��������"��3*�v�v��','���Q��n'B�ކ���=�"�P�g��Aپ��=�OPn�M��ۭA�1�w��3 o;|����[��x����o��8'����ߩ-�ц�<��FS�Pb�_�����-�Z~��c�6����y�t1E@�_Y������՗�l\����oǛwE����>��޹?�2� ���H�|n�z�Z2֏T�ӂO}KǼ�'��%���{�6g�:�>qPU��M��k���ӆdk� �o�no�C�|=0�y��O}� ����n�������Q��{ԅ?o�ȋ;vw�9�G�&�p��֓t;�˳C�̥ef�[u�tcH.Cy��C�p��Jzd�>. �bV���w��Z��.'�vZh���vC��c�]�PJ��ޭ���rJ����Խ&�CYa�z�F�s���MG�q���й�#b#����E��9�2�~��6{fvF�N+�6��]�Y������O�=s���){�H;�h��?v_=�^�׊�%\l���y��O+���?��\ڿ��Q�g�3Ǝg�*��g$e୪06v������ru�@&�{M9��پ4"v. {�CA1u;�[Pt�=@K�T�bO�:�ެ��g����z��cui�û�[�%�,Ժ8Go�֪�����{7��O�Ǒ|w~�6:�f�{��!�}Ǫ�pg���	S}Bc_A� q��6�w�rN՜�q�c_#��oϻ5��&�f[~��7U����~U}=g�wݾs�d�3��{�/�c�(�={�oP`fc�WzAX�f/�ސ�p-@�:������;m���'��]�����4*z�?aL��3�v�b���/��]y��i�k5;-�����ݝ�C�7�)����ĶKU!�x9��'v�*�Xv��޷��*Vס��-�x�ݱj�U�É̓y:�9Sfgn+��hcƕ����_c�҂ܪ��(P�R���m�4��7b����7�ꑚ�� �*��-�;i)�;�fg]������k�/5=�n��+-ꫛ\J/��E��բw����>�=9T򫟯9��~��'���^d8�� �|�����*������#�۞�,`1ޟLlVoU_����{�o�}�<���m�~��t>[{{�ReB��.9�����V��8>~S�<��`�
��׏����A����},����U�^[�Lͣ��x�=�Qiy�oF�p��+�����}�%{:�(�RW�ﺶ�����®���gy�r ����=��]��� bL��c5�
��<�[C�Pz�Ug��S�)?\(¤X��/q�V6�?gsP�^��3�0�+ŕz�R�B3���sL��d�/W�G=./m�T߻�Wz���.�T�y�'`X'��Z1e\W�ܪְ������x�{�|7P�t�ǲV�m���l8�d�bL�h���z����ۓL��(�"�{�h۫hf��Nh��=5����>�5�cO�R���z`�<Ôd�d��}ȫ�0GS�ם1�� ����팣�j)��y0�޾����t�Mr�'1��}w~���N�^��F/����l�	�ݺ�_��t�ƆD�����+�U<WuW����n|M&�������N�S�qL����'���j������#}��S��3�m�Zz��^5
����x�6|�׫>;�sҠ���{�!�{�{���F�E���;o]v�7�{��2X� ���Z��4C�/]����\��W�ď�����GS�1ʷkk�M�*�z��VwW�լy�>E'��_h���ׂ��ˠ˻ֈ3۶�"���z��e:U��\Sp7�fy�u�{�c���3�D�,0�͕q;M�j���/��������s~�K�M٫���|,<�G{ʵ�`�S������+�=�g��e����sK=��+��*yyy.�J51zn��S����W�[�B�������J}`�_|$����~Y���x�3F^�a͹�-�U�<�M$�̯z����k*�=�xrDM�i�{ӱD}���זt�-%�eo,�z��#A���'0��]Lc}.6�Du�c�(�^�O�	�NE�.=����i0�_Ȣ�Rr��3���#Cd�k�X���KU�;�78���3n�y�k+�o��k�`�3��iƶ�l�:���Q���[Nɞ�j�ㅴ9��@3�_0�~l�}��V�g�ҏj����H����8:zM.�A����@ԩ�7�����S���.���޴<Q<��?q��ٴK��K�h�4��߽M̊6Nm�������t�7f�#��2'���Xe��z���-|�(���4�љ�)q��9ݙKm�Q��E��O˱�ދV�%SН��$�/ޅK��.�מõ�1g���d<߽;���3�T�|���ӷ�]%ٹ�h��^��]����϶x^�{��S�H�d�s=�g�'yq�DY��Pz�t~H�y! ^4�k�rZ��vFg�4����]�ݽ��u:s���\W���4��
�`�>���M��es�����t�{�:K�$��"pnM�x��F��I{�"ד�F��g;]���hy�}���3�_�0A�����u��Ť��k�߉�?�V7,v�a�(G3N}���s%8�3L��`���*���rν���_7����"�3Dlz���XR]e7PC��c�ڦF��6Eq�6�q6�]�6M��� y�y��0��x�+N��7�s�߇w�;�<۔��{g�J4*��l��Ț�n��.;�/�õ;[�ox�T�����<fם�����k�ox�����:�{��h-��iɈ�ђp>�{$�U�yު��G/�L��=�~�e^�~�Q;���1x��hel��l���"n�r��nΑW��h�s������ތ�,y�F_89b�l^a�$cFQk�[������]�W�W'Q��KuWJ��H��t�Y���84�j�P��;1;�Xr7MČ�#�x�><� q�M9�l6|���A��P���0�ff�v�n��Vg2&��#3��6K�Q���</(��媧�A�����M6�_��zbw�����bE��St3�!��^�DV�10�wu<�x��w�5|'�ۗOq�߳����95�VV�,.�����u.W:vZFVhȘ�f�s�.V9����jTT�N�W���EM�){-JCA������aîض(� I�BQ�������B�`z�&�`���Ķ��L��z���t,�����mC��M���D2�c<� �wx]NO5zg����E��9lCg�>9w��^���a���P������2�ݽ���R�Z�*���q�:}����N���&.›5-n�;���+zQ=pT8=�}�e8�W��~����^�5�sڮ�O��6vϬFW� H�w�&�.}�U�w�N������y�0�kti�f�֫�^V�剌3B���T���{U�������ϫ��O?mW�~dF�̆]mX����e^U��J�����7	��qr������+�<���$����s���o�o�?^ߊ���Ν���7����y�i�R~?/�k+=Ⱦ��r׷�l��!qi�s�/W�j��*﷮��Y�tm��.{-�2}8>�b���.�\ҽ^�Uum���CoV�B�t��@�/������W����z}>�O��{<���oa ��Z�m����;�C��D��Z��r�;�D���[l�9'u�+l������mh�n��0e}L�]�������I�X#"�U֭vR�y��H9����ِ�rrͅ���3����`�f��%�ad���-y��̛A��u�T4w)u����ۏU&��ƴj��l��af�u����\T9�3��%3b�S�_\�)�2.��	!b�B�/F	�۝�s.<��1�7U˩H��=�P����vɂ����u.m�a��e�td�����O��妄-�}��H���N�mPǯ�����<�/1s�F�V-�6n�t�W�"�M;=�Ɖݏb�P�(�rD�"gtk�oR�:��.�б���A��7���J�$:V �k���2�	Y���s������[�1og#.�����r�3'%��MQ���.��V]M��ϕ����s�a��:<�U�ƈ�l��k�-7LV��qE�t+]aꋜ��q�I�U�uʆqe�S/z�ў��5tW�/���ƈ�;�����Dԍ�������],�&�U՘��:��;t�#b3l<./��ICs�d�v:�S�㸉уu���t��A��j��U�5�I�����WJ棕' q<���:鑀�_@�9���\��9�nǢ�y.��F��g���bڼ��H^;��7�R���'fr���,gYƧ��3�����_���w�E4ڏ5V3t&�*X�'����\8Ǖx1�-R9�p<�(�\�׷/��Чfb����5D�ឞ�5��l�����:�V��%;z�L9���9h���c@9�;�ݔu�؈"Ṭ��Z�p�i�k�9�Upn�G��lM9y5�P��4E�\E!Aa��	����{�Hn������np��Zm+gjm����-��4>{K�a��)}Y��!���v_v�O ynh�I@.t9Ltӹ ]th�`�_e��'t:�Єjx���2�d�����PuŠȣ�{`�#G���^صχiȇ^�.��p��^|qk�=!�N�w�5��.��9�:��t�t���&\ YaX���F5�83�r����LЧ9��r몇[vDu�/9M���q=*ʱ�I��=�J�πޣ����NKZ����躲��`&d#,_SY��#]}�]݃$F�p��,�@�S��oD`Φw2�p�g�o`��ݦ�̜T�W�J�#�"��6�<�Z��0�`E*�X9;%ӛƳZf����
����v~1刬����s���m��xP�SR�`�����}�I�"9ז,��мa:K��IQ��{W�i0������U�3DŷA�ʝ�!�W��?�7�������Y��SxpS�q,H#MVjy�C��ӿ_���=�W�'�s�R��xz)Q9ʲ
�K��j�|�f.G�E���:k����6���+j�'�q���Y�|���Cl��9 Z���}�<zڂ�4���hю1�h�#�!K5G`�8#O��j�j��N//{cI�n��Ūf��Py�yxh۷c=���u���͟;>y�1�qn�M���`飯#�rv�]��j�ֱ�<�u����uض�D�7��m�QL�S�7�Fe����lwc��y���n��\v���gf��F*6�;�����l�<�qyݮ�;>c��h7wk�5��t`׉��8z��v��.����]h�yo0o'=��5�O�bZ+�kl�ۍ��6���1�5��A��W:����TUl���1��9+��3�=kʺuC�"����(�رk`�f��[0E$��Ƃ�|�t�(4mμ�=�D���V؃cN-�y��ƃ6ص��� �:�G�n���^[�@\jF%��[�lm�Q��wn��[9|���bh()8��;V��kK��ma�Y�� /3��^Z(<�;y$mQ�f���۫�M���kSM�����wb���<.�y��F؍ۘ���^otb�'M��i�p���b4�[X� �>�_O� ���{�(��yp߭v�G��5y}>��4"��JaoC���P�ŀ���r�f,ri�2T�����.��Y6���Lg	���Ⱦ(�.�Q��D�b�A���b��ـ�P��M:Ǣ���g4"��n=��1to�ٰ��bw�ӷX/ �Q-#QI���N<�)���W4Db����:Ĭ��}ɯG
�{�	���O�o2Ho�ov�JPm�e�����[;�J�����.4���j�^C�:a��Y{#��S%4��'�5�\M0�j'�|e�ɡ�և��7y�/hr6r:{ͽ &f�AdM�¥V��3�:C��ΓO
��*[�S�ɩ����wu�]s�x��^0�]����1j��bۀ+�m���O�xM�����C�V?��� ���/8��z�;o+�cT�s��㗲,n��<���R)��S��YQ��ۛʃ�1=
��iU��k�a�e̻�A�v����G��
�J.-̪\��Zrs��^֦�kq�91�8ܝ��N1v����[۝0���<[E�z� �'�2y�:)��y*��� _=ϺL���xl�k@�Mjʓ3Lw�,V��U��N+�4F?��K�osP�75��k��i���i� $�� q�I��=X�;�t"w3	Ɠ��Y����w�ץy[� 8��8z��hK~W~��j�^�(s��RF�M�N1��hket3�6F6�23���v[^^H	�V�s��&���6N�y��V	f��0��x6�RÀn��wPKD�^���U;;i�3�F*Ӷ�ʏ��L�Y�\LG���1�)Q�}��㿷��S�憤+ �$�q����Wre��O�D��j�LG�ޒu<!�ә��r��\���.�����{��+�ӏ���eĮ��H����w�N"�8���/30��F�PYݏ7L���gɩף��v���V�0\����b�������فJ��-�E��O3�Z<1��՘��B݋��#�)�;|��n�k�:�U\�
����70Q�h��%�'��\ �{�v��Jj�����%@�i�y~��mށ3�6�fh��;��y�/g�{��1:_@D�r`� ���`��.�z�V�^���z��6�
�"�����5���RƋ�{/J-vW*��%�W���?,�O��`Y��ʿ�	��Lr��r��4�w�f�W�m������m{7 c1U.��*wG�TL<뵘s�OB�[(��T�<��?�PZ���T�=ΒC�S�i�_��|����qEyw�U竈g�Is^N�Ku����G�K�=�aY�u��A�=Y�/�VP��ʱ�)�tD8���=.I��z��t�0�e���=�MSz���uUE�Os�Y�t<��aT�g������75��#�ݏ�l����<JߢCfm z��ȍ��us�������u$��(=�\�šY�#k���޼��5��cGd�s��7�fk�Q(W.�����f�|(�`�+kA�'�>�4��S�Lkuʚ-���2/K"��;B�ڔf8�n/D�vK�t&o{L��Ff�?^Bvq�dh4[zw��%�I�M�f�ݕ�[�d�nx�_��O�{���*��S�5��x�˵����L�l���^��7�}K.j/d%:hc�5�yJ/Sxܮ���W�e����Wk�y(�n����P��6���"���H�Q�^��\�=C�ޞ}�x�U�>fn�[Wc%�~�<�L���EIe�O�w��b�|ZF����X@�����[H�d��X-mU��U��5c�yo&�g�E_0��)�����J����=�ib��JUN�< ���Y�i]H˴�R�Z��.s/��/�ػ�C�m�y�zy����L�Xr�w�Kճ���2�2uQ��f�jR����9�[�j��Lv�a�����Rb���TWzX]�V�u�̉y��^*1��f������d8�L,@}k�4ɍ�\�W���@�ۇU]J2���T\j��1����-A͉v�6�vf��>J��F��դX6~�~c��<���1]��4��1�����bw����M�dm�Q�j1΁9�{<��o%�i��p�voG�j5�-� �謧�g5b��ū-kt���� p1���-=�ү�J#Z�����d�S���qu��>�^��Y�Td���C�X��Sy����O���l0��ͅU&����TK;k���l2"}*p��mN���)T�o�N���r���*�VK��'��Ci-�����r�hOC�]P�����q���K�:��MWW74"�~����qmmۛ�M-B�z*moR-sT۸|�+�`ӵC����{�tJv������'8��/��\i1������ޡ�B�)ʊ��}/W����Z��/=c�u�����_@T��J����M�{N
o�cŧzO��g��d�g�SQp��#{�s��իi�xU�=ֲ�Rˉ��-�#���
8׼���xu�:Z��'rH�޼�WB�0C��0�
�d\��������aA(̈��]��p�&e�;�v~m�,�z��������\u~s�LXXJ��rSM�������k	���1p]������ ��櫖�Ԫa;s)�	�n�摊������qf����K�p��T+p9���g�[�B7/���mZ����"7�)��]���"YH�T��%�A*y9
 ��T#]��ۇmR���))���� ��|�7.�j9us~kP|d��;2�N�X��zx
� ��m&Ä孇:�e8���9�w���g�>W��)�f�U��`j�b�Ք���ѱ��I�w��t��u1(G6�Y7��&�J:U��2� x��/�v��h<ޮ���������4�Wځ�/ k	�z�S-{��[g��\ю6��pȮ�&ι۬�ږ�[�����cGpy�w�cAaw@���o����Κ�����V�Iˣrj��Nl��]X�6ْ��O=�]Ji����f�F�~���y�x�Ɩ��(������υ��Z��\e�p�7�f�ԖV]xʑ�^��ϥ�r�ρ�5��r�x�uz��~~#��Z�O�ܔ/'�js�1����c�?_A21��޹�=Ǩh�Up�P/a��^̻Gc���l�|�N�qWx+`�zҡ�y�-��J��Fw�q�����~Tx	�4�{�$6�=ڣ��㕘}��{bٜ���IV
^Z)<{̮����G��v�d���g{2� �2��B���L�͚�ϧ�јo����v�m!�j`�g\&�:�L���v~������PV�ڦ����kz�m�b^jV�f.�Ss��cڭ����Y/J�\��τ�Hb�s�ʣ�T�j�G(oVp�*�{��򑦐I��~�6z�M1m������֙�{WK�E�g�T�VJo	�ب�ڧ#�m�@�ϻ\����sM׫Gx	����Si�Û)�z��Gk/z���v4r	��h�5{��t��~��n]�1uu�;�;�II<ݽ	\6�3Z_C:nZ��Xs3�*U܁��e��2��GQ�o8�s_B��|��}|p�c�P����;��"o�3Us�k���)�9]���"�(�1��*u�^�l=:�!?�6E33��X��A����s��j]��B�O53t)EŹ�K��NNT/�U�����;�R���\�^ɚ;����*�ڪz���o��;:�������*,(�.�d��[&{zy\k��Hf:+v�3r�0��[��y��,�x�K�_��#79T�uȆ�~{9p_Ԗ�c����ߓ?������{���I?�iO�ǰ���V�6=��6)�fn.'\]fS��uΕ(c"T�:��Bh/�,�Ϡ,h�|�x�;z��G��,��5����hS��27y�S�t(ŧ�dU���m����?j��^�|����#O+�7y#�2����-ᶰԨgL�o�B\,Q�6��x���18�H�Ƶ�4�V�q���ó�viIM���D�Lٙ�S=�K���%P`�1�o��;ܰ�<� ��~���<F�İ��]4z���Sl�됎}�2w������.d[D��|���Ր�>��C��;�5.#��H���J���Tr���оH�fX׉�M�o�us.�I ��vr�{.��\�,ZmL��<�+���7�W�<@+Y�ĄҺ���0�Q�4��d�J�k^λ4�|����U��ܖ�;umˉ��
�y-��Z�b%66��?~��J��Y��k�<�@Z��HTF�p�g8�������ZT�sK�2>���"'ҧXLL[r{m��زj=�7ȋ�����JsYń�=�H�g��t�y�;t�˜���l���ŶtW試�%sM_J�bL�X�&�!����f#�B��-u�m��#6�>��5�X6�+���]gR�gf9�P��p2�O��Й�`�T�}�A�='�tUȜ�6�YbɈxT���﷉��n�v�^�p�\�ָ�\�tCY�#�xzv��12�@�Ƚ��I��-�z�{q�Şs������Gi�^;�v��o@�p��3�jfͼV�Z��2Y�)M�Qm�o;ʡ��kV/��(m�v��:�#�{�P�����P9���;#w���}�i�>�����"�ݨ���v
	�����4�X�59�9��ރ�� k��*x䅵�{�i����rmL�5�8`��-��Qe���b��M�uy0l[���<��
���Q5G��Vu	�f���7��3��7/Le�@c�<��P�0a� n�k�F�$����+�����V/XT{�fj^$�d�h��U$���SY��Ά9)���1ڝ��Y5�]
̡{p�\�w�����Ɲ/�mWe��K�}�t���{u��"�"i!�vY�(t�V]��T����ޛ��qbJI�D��1�U����sY�d�3*<IN5�;cq濼 �V��;��aϭ�LB}j1���{��8�� )P�(,ڂ��Q��a���"u)D��nl�U�W��R��*.댖��*05�b�ۆ��F��-�ڡX�OFErI��2T�-�U��_:&Z�g�U1c�m	�i��}�%ߋ���L$�4;_P��Lk�W1�8n�t���W��۲b��s�Q�o\k����O��b#��;��A}��y�'�KcD^���-�+,�fߋ���@?@��x�,��3IUI���C��t�<9�6<�0d#>�}�L.+{!�����t�������[�5N�vg�g�Ih,6��Sm	�]oU��\�&�@KЫWϰ��B�����+�}��]C6����z�PCm"�'5M��,x�E��	B�#/��B4��0^ɇ=�*�ϼ�xkT�C�)R�O�꣍�D&��iiՕ[Lͽ��&{��#'�X��4���O>��\<4��mm .�YDt*��؟�����է��� þE̵�x���I�^݆u���Ve�Ϻ�J�V��HfU�sT�Q}��ܾ�߅�(#����w㸇3�qQT���d�S��u�f�������9�|DU ��m��9%�xG�G�p���8ˀ��H��l!�x���g������k��8���m)��MJ�j�䱣M v��*�ѹl1��/�s�c�wdƲm����y�q�dd����'XRS)�`*��s�J�n�3&�O���W����ܻc�y�nd��nP��ǂݎ�a���GI��=��酥�E��)���)8����.&ޏ$�L�]B����̠��sW���4v��7�"��sJ�|
�l�s:~l*��]`���i�W&gD�8��3����[2Ls�r��z���	U�ӹ/�CV��n�ksM��\����^s���'²�%#�E��
Y���M}u2�7��[XCj��f+Z�+��r"^��%5p�F�>=���?�Ǝ��	މ���.�Z6��jη~��� %׳�c�h��X�|�2K�0X�Z�3@�V��l�]�eE��fKU�d!۴+z���ۉ���\Э5{Z�MDq��k�.b6��V	�f3�L��55�5ކ-������m�4ȴsl�	Tv* �gD�`�5��_���7��l`ks~�}z��	&W����2_���G>�7|pvf��54�OW���O�d��~,��O��*,k�i���!���7p�� �����n��>����/��ƚ�{�g�
�@�[C"	n�]�y�� �!
&�m���w$�Y�K���)*q��"�T��^i��D\[�T��ܮa��ī�ո'n����pֱ�|�Dy�;���Q������Z�;Z�`��+�c�� y0�=�{�n7��#t�D%����O�'FWD��}��ʷ�v��28����޴`�}������xl����.R�H޶��8�BUʒߨ&&���0;y8�t��z�'��v�%�G�� ^� Q�׊�S����p��q��v���+�b������Ma�p�&�'O�z2�Y�\j���~d1��ȫ�l*�ۮ�w���<�N�Z�<�v���eFJ��%�Z�N�'
l���m�F��l��)M�����m��9��CD�k="�)�u�z˔S��J2�284vb�`��q�eU#	=�'�����&	S��;#�m��5�і��2K'!�l{,3��M>�0�����h�ιgj�J�[�\cKÂv���f��s���Rڲ�1T=]m��ژAo&щ]��u^\�w�CJ�L.�kx����}�׎T���:T�e�yږ�3wݔ��h�*b�~�������inj���c.�fe=Q��ܣ�^<�SW�Q��P��+���]ou(�R�N�-�[*)�b���������~�o����z�^�p��yy���׶-�/x�/9�y�9B�7[���Ev{�ӷ�.]L��}��u�w�,��T�p�EPU�6�Y/��T9Q4����B�֒$�op�O��|�oo>d��^/,u������-kx/MLW����ؘ��YO.����~�U�ٮ�36r��@_bZ2��F��*�[�P�a�Yr���\*U�Φ;1�t5G�o:7�Z�^���h�0ԙ�����ܬ�p�"�2��N�3��5z�-!��h�IQ��A���t=�-�M	��xFZ�/�/�ќ�fN�s���SK'����va�1<�ə�U�]�,�3a���`��J�o�0k�IX����5:��m���� +����%l�MZo2��{��%.M�.֬bovn}U<�P��sF�jU�ź�v��v��ma������4/�y�Y9Zl1�=���8,Ⱦ���L����Y[٩6�[vE�k�<$"��d��z_*yz.贀��a���î<1Wm5@GUg�LN��P�(�x��.^�vE�1m^"P%���t��y�l['�k��fqV��B�r9:�˂���Jm����NM�+�[ާT=�,)-��.���M���u��(��h��cJ�aS��<�*�۸d��5SuSw���xgc�hڒ�u��AK[��n��yȋP���}�8�n#t�h��ׂ}&��32�����]bn��x�ɫ�}6����;��Uc탘r>#���n�{�Jtg\�qB��S7���&�����@�zl{�j������=���tQ��)}+kX�4lK������������u���-�+��/M}e�y��W;��Lx�mg6�y�D*47��(��:[�̐>��[�&_�=f���#ƍ��dVp������M4�4a�5.^v�4M�V���UfKYi��c�|���S�K�!�Qv���%�wQAM��N�i��3~SX������V9��']c2���2���{ꇆKM�}�6�ʅ�-��Qb�';맒͢��t����d�Z�vNt�͕���L`�-�#y�U�>=&�Jq�P�uɣn����;���wl�:����Lg*����Q���h9ү6Բ�\�s��R���n�su�A�L�W2�oM,K;b��h\NQu���7��>�l�o�� �'q�B8+#(w�hWt�/4i2�8󗶩��F��Z���I�ŝV3?vjen�czN����A��$w���MfEą[�;.�:��Y�;2����*��x;E4C�x�8�;�%RFK@e�B�^oCm-Lʹ]w�U�G�j�խ��S��5�f����r���tL^,�����u�ԅC�a��u��wt���u;Nb�{��e	���W�B��oq<򧕁dՙyq�������gע9[����e�`�{�T@0t���90Ѽe]賙��Lva��
<��I���{ �כ��ے� &|�����T���x^E%&�>^F�'l�M�"#�'ATyJ8�1u�����4�۶tii�v6wq�6<�)�#��h.ؐ�[th��Tu��ww]����֚�8�:*���j��Jv�m�Q�IS�h�E�v����s�w)���b

֨��kUѶ]u��lm��-�M5��Q�`�N�n˧�<�&gAZ&�th�A�#��j
&)*�j"��u�Q5F-TEUL�5��V؜y���j�&��@�X�#cUU�j"���C�Eyk�l�tWlƭ���a��:�T^j��1kDu���/#����DP�EU�ĄUAmI������PkT5KQQR�g�G]��U��ci
u�[Z���kh�Ί�ct���+N�5�6�%AV�S%l��h�*h61LlbѪ�bb*�(�ŋi4������|��+��J�VW�OI=����	�vy/Z�:�{�@�q�6j��7�R�f�%G9IS�����o.a�+���"��QQ��s{MX)6CJ&�m$����m�BF%��0��q���	��,U��g��X0�������������S�y�л�L6�Z���O[���xń�b����E�;��ܥ��}v�2g��Y���n�T��7�X�8cS�Oe��q�41�U���Cͽ**=�K�B��+��>��h�X���Lʧ��I���uޭ|��\Q5��S+�5�#K�2�D���úWY�h���c��*P`������h���!�C%��v׬�f�Ŋ�j{f���uI���qiz��kJ�P��PLMPc>�Ϟ��v�����I��	���/���`�늚���(8�nU��IU�oL
g41��o-�?�{��v_{j^3������:SJ8�^��k�^�j�C(zH��k����w��C㘔n�a�U�\H��ji��L�R��w�P/A��\�0��+^�P�U��/��Fh�X��Mɾ��f��ݻ6+�w92by��KN���9�"=ͼ�n����r��^7/a�?x��e����MfEgPH��S���7	��+��w!�Ȭ���@�?����B/|P��&��G���>�����x6��o�C�v�03N'��%��loa�S���l�����{/s۶��z������|w	�M:���*�;�R��;�wE\�U���n�<��c�K�=�h�(!v��_c?	:��`��mE���v��0��ۑz')�����xx|�xxl�eQ!�]��%>$�[i4G���.S��؊,ЖFJ�r�GOջ ��:�rjZ�*�sV���ǁ���3+��ژI�g�<��)��"�3�Գ%�<�`W�����.��m �0v��O�G��Xk�^���K@|�4�Q4���{�W��}[����ՂP��*�9��v�����}9��\3�j��M��c�<��OB�a��R�a�,���	R���2� ��Ĵg�[���N��!�ULF�h�	��{�����qT��h����??��drv㈯���֦	E�̏�|j/�������aP_=�}Nv�m��-��ĕ���}5�6svrqE?Hv�݈IAg�UT���1��`�e�6�?�ym���k_`��IѼ�Tٴ��O&���E��U�A(ַ�k��C�SƂ����w�C��j��@���Va�0m��y�m�[��I�����v�s3��K�%�������b��=��]y�|��t�I׽�iS��m������
�}�bZ�ڣ����=��!���*��O�M�'�y���G;յz
���&��U8��H���1mJm���WN��̆��=��e��Өԙ���R�,;C���u����]�.�Aº��:��/0��
%=�oS��6�W�-wV�u�M�n�:�E��[���$4� v*���ͱj�U��}�U�uōg��W�������5��L�����,��&��������ݙ��/6K{	�mE�Aw�j���`L��l$�	�[���+�a#&��hb�x����F�5O�pzVo��0�M�鼆�N���qh�y��CQ㧆m��3�'��Y���2*�O���sL�:v#Ļ�e�]q+ț̺dzY�*q�}]�0��w%aC�UьЛdR���~g��A˜vvl���R6F�RaJ!1Ԧ[��Ʃ�����y)���~|�S��H��]��J���w�d�����Z��;P~�/�c��%:a~K=u�ӈ��=2������rP����ݫSݮ�e<�4en���F]��H��Y4��F�\1�%<(���@j�m���=���%����\�e�=�F㘼��)G2C���ū��%�u�s�_En�B+��OS�\҉�:T�t^7IkQ/؝A���><���}�z�|C6�z�L�ϯU���-(͝�������ܹ�PtP*9�l`S��ö�@U���Ȇ&:�h��󡹇Bǽ�4-(��yBn̻�YR��]�W
�.��cP�� �'H�kS���oR�0M��9�������R{ܶ�䋓�Į�$y+ˡ�N�$�4�4p_v�6�+*�Us��{"��%:��2!h�U��_�U}��W��f���7�=��}�j&l&T��)U��EW7`]%��O���֮-��h`��b���uG���'z�u3��@�k��'8�v��F�����c֕�7�T�z�jk�j�v�=�Gw�t>(��]�|^ā���:�D����T���1�*�C�01����w큀�3Eۖ����0T{˚�@h`�D;�&N3���'�x��{�Y�?�Cvw��[p/��ls��λ���x�y)��3�c��K�=�^\ZZp,��@�&Zr���zY�X��4y�R�Uae�ج�m^N�hIN���2�-�U���WP��ʒߨ&&��c`v�����i*���e���J�r��M0�U_��a�ĕ<̜�����@��m#3�	���46�^�S����_�p��C�����\ԃ^=
���d�j%�e���\cN✇���/�����8�Σ�D���H5y~��vk��^&�k��q�):⓱����HZ�i�24m�%�6Gɇ1_�#/&���Xs�X^�ʾ�ƀ���qn����p�0�Х�2�����P��e���r�(7KX�䜭��<)��MX���c�}���9^%W����Ӗ�7��CZud���t�t��i�dų-��r�w����i��*��(M<�ު̨�u8Tܾ&ɼcުgu�x)]�b�Ҁ7+�2�(J�������_W�Cm����fnGݹ��)Z���������5�dX���eQO����~[C2q3:\���ﾪ-mا[M�:'E�V�Z�P��ADV:�F��Khu�����/��1��/���!��xd̓_���gL�9�Mٳr��(Ե{���Z<{���tke߽����q% G�*֍�A��X�3ݗ�T�X/��˛B�J{[�)�խ�mCr������tk��G
�@[
*��;���{V�xEƗ�%�?�z�ƫ���*�����U��>Zn�j儩�5"G��c���^�]��s����>��eŪ\v�zO>��C����4�#"�il�	V©b���wC<��Uޥ�􋼬���D$�����0>)-Rc��#�Vj���f��H��eq{�m$��)�XM�C�6�QX86�y��c�,�%��ފuZ��eV@p�Q�ע��*�]G����C�rh\{F��Qw��t֕8�/i7��G<����+~��K=�d������.���!��'3*�k���ͪ�G��W�RS9厊���d����S���~,��«7W�ڞF`��D����w��]���b$���A*���e�W���|�/@�Wj~(m<%��њ9�9_��xM�u�kr����!͂��2��s;���u���j��SOc����j���h�7���7����<=��YU��zro^�/X�ڽw���^�c�zJm�dK]_<��� ʈ�n��O��mI@]�]Ͷ�f���dUxD_\�*:�E��i�yj��~��(z�_l��Z��K�g_~�*s���z�1������DG'Fo�a9�Jv��a�ei/���f�/�Bi�M��S��Rڶ��m�g1�o�m;	��mL���M���͔���
�l��{���@ޮ��u�Y �g��
�>dJ�oJ�F.��s���榔B�ӹB�E�^˼���\��T�i���[�Eԛ�A�/�3HG����e'X��w�oVGmJ\���M��.P�J��7D^�.!9Q'{����V�]z]���%�Y-!�_L(R������8�<�@+\:~hw��s4��O�dT��ɵ��<G1�Zs�_m�E�idɇZ�a�d�Y,s<¨)6���̳��y/�)�h� %*���f-��I��Ϻs�
�C��Q>Pb���#�=�N�|۳}�tТ�ZFK	����~DȘ��\A-|���@����*)�����p��Pb3�w��u/*R\��1c����X�芞�b.�Kζ@뉅�A\�a���m}�e�ů4��׋x̵��u���YY���dT��N}��s�K<�m4��2���ա��	Y��YJ0�H�|{�jڳ�/���wP��L�r�c:ow^O�U}_ 7���m�e�j�T�ȯZ�g��UTt�y�~U���~/ғS]��!|E�Z�oʊ����U6n����ilZmYf;�|L���5Ͱ�bc��kà�Q�����-|����E���wL���G�K
��έ41���<��4IU��]!���gR��\�G%qj��hU���y��D?�$��O'�KU$���KQ<�{�=��uklU���ѱ�(nF�9�Q�a�=n�.I�Ï�'��}�%;�;�7j��z�zB�;$��*��J�����ݟ�g��� ��2,th�Ԝ9 +�+4���D8��RQ�)��]�+9s��
�en��-��Х�y)ʀ�!����+����+�JʮsB�	���
���a���{=w�Q�+ŗ)��<a��[4˯k{h�b��>�|w\�*��,�}mM���D�����,�kj����HA��ZA��	��L�Z��TS"�TSgZ���2 U�E'n�|�H@�Ư�,8;�,k·m^�	����h��={�R/a�Jt�ҩ-݁*�~�Rv}�;��/�`�)�˵l���m��[���[Y��>ߘ�S�5�i���(�|���/�n�V#�j��P��?Ke��IȲaܢ.���ڵ�V"'�5�7�c� ��0������Z�e�#���c%@]f&m=��x\�у�Q�,�ݮ���BrB��X(w�������U
DR��Q��r�_o���z����q�a��nK��	�!.�Y7ax[ƕ8>4��N�_��o1���R�ʜ�#���6"�q�_��!��m �2"!>���!���%�����z�� �v�N\>���ȁg/��K�F_t�2��֓u��JFS�M�G�O�!6���k�U\K+�U^2ͣx�Jۙ��H
�d(�c��<���]��@��Lh,����T)�l_��_/�����nm�K�CC&Poz�Χ�
��/�S�7�׼1�[�(�[t��x�ʢ.$UT���\��+�a��\B%�62Z��\U"n�����t.6=#��C�չ�̚�v�n�;!�����Cs��s	�X`@O���ީX���a�OM�>�CS�s�m~m��K�e�Hɦ�R]x�$Z�v�^ɖx�	��d�.,��vl20�m���J���܍�'`�i^)�`�oM�Pn�=s�Z����Ȥ�����ʈ�R�R=G�
�n٪^2�[�V"/`�PȬ�v�	Iq��%^���Ѝ�s��Иΐ��qMߓ��r�.Xs.�Et�ʹ�Nּj�M���H+��V�_=d���aQܸ����1�r���Qڐ�ԎV4e^��3z'Dk��>�\��]��i�y-���M�7��Y���ۂ��v�j\M���i)mf�����)N�����<�����y�~�}�_u�D)P�{����xx � ����\����wu�j�`�30*������rމ�_d�j/���}.*Zu��3�a:CB�ᗦ�����ٸ����"��� �ȹ��蕯��2jY���V�7_��ֽML2��l��35�")gf2�Ԯ~E{n@�Җ(���i��cŋ����{�:N��\Rsc�m�Və�d&I���q���9�]�v]�=;�����-Ƿg�O�G7���+�7B��e[s�*�s3��zkb��?g���)�f�c`ӓ����VRO���3�����|K�L����cs����T{�i��լ����Q}�R<�YCl��@����.z���bnm��#:���Q���
Z���}{Ӎ]�(�L��P��nBGh�����������m��w�wP�sy�^����
�<�/��j��bj_�������_�ԭXPS]�K�LP[����٘��d��\�/%�y׮}8Ȫ�U��c����خ|�L������fz�/	L57p���J�Ý�)�M3R�/7(�o��ekG�����t:˙��q#C�3���iG��~�<j�JӜ����9`0��d�����g0�S��F%�O�sݾ��/,�g�T�����]��=�܇RI�er;X��Z�~6oqQ�7�?����۱��-[�U��-�jZӴ����I����/㕒�$�ɑ f�`��]2Í7?�����몪���7��<0� �����*b���M�U�B�3�~D$����Y���ײ=�}��m����z��V��Z�H�������q��B(搘8^�21̂�N�r�]��ѝ��R+d:v�"3s�3CZ%W��n,��猻`i ��,x֕8�`����c��~W���g]��h��٣0��A�[�aOgU3����Rg���p6�����*`mP�����WA��]
���Ⱥ�����z��N	�ژy���=���`C]_<�̵|�w.���d؞pe�\1eG��I<�Α�;,�0�!#�A��~[.�(y�(�t��k踫�:�2���mh�x�ψl+U�)��rbA�u�B��M�Ά3�Bso5k��rʭڀ�MKlP1y7U��c+{r'*�|\�Β3e�=�"��U����ۆ1�W�E��������J�E��^3������ʼ甙7�
~j�Ru�O�6���	=5	s�ۋb��t%�����"K�����f�$u� �A�Π�|a <BN�<�c�J}������؇o�{�9�������~ϳ���ϳ������#��Tes<xo��ܘ�m����f���M<�ތ�x�OD�ɡY����>����<����� ��`-��:ޥ��#����h&��N�ɽ���24��8�3'�bͩ�b�_a�Ib����ɝܻCi�q�3�W�f��РRhb�s���֌3S���vv-�a���s�6e97տ��&�$�'�vr� �s�VG^�r��]t���ᗨ.�����6p^*��a�Vx���e���SK�k1(܄��i���tv�a�Y�u�l\�6�IK������c{��|�I����ǲ���&"��n�̼�z��c��A�dK��,̺�6�6�d�/=8���ŮL��U�s�f��*ͤu�*Ĉ���ih�9�jo�ew�ԙT�&�fq�çD�X	\E}Cn��U�,������T���M^M��u��%,ܼ��o��Ʈ����J��R���OL�a�t"+B����7X�Y�[ȋ��z"�:�����osx`u���*��Q�;��;��X��]��8�xF�r�C��G��L`�$�:����MN������aӥ&�AQ�Yr�̧�e�4�5�����c��w�۾�8��h*1�.�{�JK�Ӹ$k[

�ͳob3Vn�yy-�85�p2�����֤�x��6��=���C�m����-̜e�uG!T�sٷ��o�u��nߵK">� 9ιm�UI7��������\����'�t��.W/��5/�a�"8��1�<�����9|�+km���z��ͼI�݀��^Yo;�V\�M�l�&�t2`����W(���[�M;.f�]Y�Ne�`BD��ީ��Eg�"A�rDv�rGW��\����ct�P�\H���9��iM�Cl:��o�.�	)(V�'Mf���V��d��sM�ߓ�tD9+]x���Z�`�!X�W��g����Fv��=�e��k�&�y��;C�JZf$��9�R�6q��֙S��ZS�Ŕ�/d�3�M{���
� =�����]�[�[GA�"2�Y�.��Ζ�A;3��6�^��B����S'�凕jlz�_M7���t�<K5�zGhx��v����ame.��͢�����Ebf�YbR�6��+2>���Ĳ�F�=ߔ��en=�Q(�]ƥet1q���`_]%
�f���\��AՑ�B�y��KkxVjdU��iӈC����GZ�̜�J�7o��	}%��{e�[�=aއ���:����-�α'���)�\;�^o5��+�w�R
n�5szf�� <���e���x���c�	h��5ckENvMKŀ%z�jU���^A���˥�+.�u��[��
�z�
8i�`��׸����$����������"u��v�ؘ����V�Ỡ�j��*'ͻi�h�")(�i���$��Z�4t���+[h�Y���(��
�M:���AA:�:�51�EA��Z�f(��)��"{fh��!(��E�mF�ZcF"A�$����*�4h4kK�TִQ/[���d�*��f���b����clE[j�&���UZ��CQM%QVح�̚�%RD�EQDPm�c:ݵT�j���b֢X��h(+I��kl[Jbd�Zb��(�Jf(�*�Z�Vb&gF�AZ*�	�V�h�*��*���&�
����hm��j�+�TQ�kl�x�^�|�}__^���q;ɤ^���G�'�����=��a�O�{���t AJ�^@�;Xi!1V�H7LCu�s-c��̇����Q>�-B)�J- ��R-(�H- ҃��'����Mi����*��}����i��0��������ʹ��qw%���F$W5�jz�SCǡ�O̫����0qz�<���im�L8����
�]<ܸ���J]8��D��[k�?0�*�|ĩ�	���%��dy^�#�f+�fub��ܬ]�*�8�j�y*�1�e6F�5F�	Gs������4�`w�1����X_=?�ԏ~^�t~}���Uv��F�^�~��gƪ����KR5�֗�Z���h���2(F&��F�X%��rS9��EVC�9n��L�jœL�R�\��q`�ַ�5����j���`�	�(��´�+޸_��{�6Yxt"%Iזd���=�N�f�Z}���0��ͪe6-�e��iM�U�i����j���X�����|����[xԱlF��e�7E�CkSu]0nnaB����tU�wu�Җ�M�c�R֯Sp�8�Dg�bB������o����F�\��{�^��/��Ӈ��m%��}�[���X�S�z�:4s���ʍ���P�2RQ����f��|T����n��&�,۷�_��,"�(��Ψ�aJ�7j�k�sx��+?ndQ�X|��6����%2�g=���8hn�l�C9h�:�7����5��uNZ�׷(K�"S���˚g�`�j,��s|y�;�㾻�-�"�y
hA
ZD(P���V��f 3{� 6��i��fY���DkG����A-V��
Ϯ6�ʒ�Vl�˾�?��0f}1��X�X�7�gE����:���4�ە�ң�ڇq�O��L��V��z�Re:�$�� *��yYٵ�O��c7��Ϻ�����S��6����tĖ�2�rS,���n�YX�'����}6l��̴}r�M� Z�t���j�}݂@|ԭ7��ÞS�	L��ۡLT�n��
����׻[/�ʧ�!f�-ف��4��=C��y0���p\Ң�;��<Z�ER���Զ���r�V�5�-{��(�l�{]�����m~��,g�ڮ�[`ٸ����v�g[��;��P�=:](�]u#��tcsP��Q�0Q_j��3�o�8�9^��n	e92�n9�4�qRkk�UC,q���Q�أ<Ae�0��ͽ!�hh~�A:���X�$�u�KLa�6̌���=46�F����*)��9@Z��j�j��������\�j�׭I�C�~�9[{{�+�㠚v�.��Q\d:Z��Ǟ7gی�z�S^���)�Z������)��1�lA��~�#�ꅊ���p�[���sK��{S:�ݠތ֪���k�U��M�b������B`��ԕ�+�Zp���4���4iB�^g5w�A�s�*;�H+���"To%��v6&$9bye�Z���_g<��6�#���P�\G�� ���@� )PH����{�f ���Ft��&�T{���<��_�,?��G� ������<�A��*� ���`��[��sD"�)����|��|,|=*��T"��s�&N3��̟d��|�"s�h�0��`5��x���VZ�+S�KbAm�r)7�8B�{�,�`�y�ai� j��%AOSQ��Mi3S�=c
��漱���ڦi�ۇ�V3L����x�V���0�b�_X��?�d��盵��z�p^4�.�mG]MG���k���Lת�2{��}U�7���aR��靡H��.�(;�P��:���VJtQ�L.�0y��H�zis� ɍ(���72١,�7���@OP��}�Ko��rt�F��?|�J��Ǯ������z�9�c��{;*h��<�E�lQ~��صW[̛T�wuCA��5��Y�m+�b���-��x���AP��|��`
Qq|���n����*�3i,'V��Ͻ�h^�d�i�ra��c�a�9Mr��e:ʪӭ���Š�fkJ�v�=:�:������JGk�Z[C�S{(;O�􌚈�X:�m-���l^�r�I;�H�~<yż�*���5��-�%���vo��Vcq�Y0
w^a�ch�g���K��q_[��Up�<s�ڗn�-[���	��VT�+�R���|妟lu�M}�q�ʁB
P�*� ��]y����R�xd��e��w	�jܢ�<�=�ň���H�b`s�C�}a�4��Fᗋ
��eӠ�l�heD�{��2s�R'�E�M|tI���M%�����_���R�B\�IK٧X���/b6�)wv������ �^CG:/B���Gi�w�U&kg�е����jx]z�swx�o�s���h'�%d�q�P�ˍ��׎�1�.��4\%�ֹ���5�mU|Өk/.��>UU�_5#�����@�M�/]
H�F���k�ħ�L���q��m�-�� ��驔]�(%5�R�5�4HC%øqwܘ<��"��|���2���'�|*sՔ����u���z���Ar�ՠ�荃=�ύ �쯕���[�	�h�r�7���Y����~ñ���Y4�bb�k���1��"�8����{f�Uӳ��7�6�6�J�%7�(��Y�h�;�+�2w*��5v�Gy��V5p>jJ�+έ�ܙ���lԯ/fYs���'k�2�o��Ǆf��k#��2MC"u���)��R��gB���F�����Ci�Oh��&�a��1���@�y{�5&| �훜�dJ�V%�]O1Jn�C?� ����Of���y5$�7G1��k&��X[�)�V򳤊����w�w|���V��Kv�kG/�6���^�g��N$�hd]���l˕�:
ݡw�n�i<�~�磌�Q�dI�0ju��{�j��)�5*����Ν�R����MP���=dWn�:�2]Ebs���%ss�ۮ�v)>�-�{`��B���DA`cG�]��o��5�(oΞ4��iB*2�Q�����#\�� �f1�HH���ͻ�^��Cm�׬}HC�9�������·����R�>�][�84��4z��*~�I�Oǟ��O�@�r�٩̈����V��׬��+a}ֵ�xf�v5{G90�n+Ӛ��"��o
�5)�|������h׎��4a���&j�qLQ�7F�)t�^����P�K��j�#�r�����	v0��Z�auܰ9A�LA̻r�Cݾ-�����lJ����0%*�/1�9�~r���������gq�|�v�k�.f+zt6Nj��CKd�)rU�_ݤ�G����� ���_�����cCS[�5��|o`z�X�\s��;d��Nt�e�J9R�?�Ϩ���qV���T��1��0n;�V5��Hx� u�]�᢮ٖp�9:��լ�>2�mnޭ6�D�k� �Ʒ�ƹ�^�j���Ļ�����iH�We�nD�b:�1�"wk:�;&M�x�Xߌ�F�S����vMz�5$}�F�m�ZZ�j��?v�R]���n
F̹��$K�����	�=���o��Ԝ�f�c�uj�k�a�s����pΎ��S���#wrF0�����<�7�<=�/ԙ�����'���.���Ǚ�:v�4��Y�s>x��M�}�x@z=Ul�T�khu��\&�+bY��D{`6)0��b�(����vq�̧XK3CE���T�4��x��+$9�b���`�}0�>�e��:�kխ�y~D��I��\�89f�a���l\�Bȃ�E)Ð���Cm"�'5KH,��"th�8r�TC�����5 �m��9Ϸ��|�_�{�ֱ��%4R�����z��U{TC��,��*+{�ZV��to:Gt�?P�J��H�g��1gC	�l��X�ܥ���(�J����T��ӌ\��Odֺ4�O\ww:�vnke���-l�ߺ�K
 �����d\槛n�YX����J���,h+˽�S�\Йo���lu�lF��4;d���ې�p�^�T�ߜħL/�T��������/XNGt�Y���6v��4IW@�7�[V�9o}쀛����i7B�:��J�b�mD`��|�(���j�m�+���vx1[@�z~-���'Wo�`C�?!�
Ԭj�~�9�m�$����!E`�3Kܤ����童�x~��D�Y1��܏HS�9�:��h�J9�X����b����}���T���i_1�Y<�J2ƫT���W��9Ω�;4L*�|ɀ���M��d���o&\u�yUSט^����� ��$x .l�sW�T�m;{�I�E�g��mӶ��,公,��&#�������U]���ѯ�v��vYhRو�S*Β���)T5 r	G/9}�S�kT�o8f���42�drin�#~�*�;�*��m�E>\YgM�ޫ67��p; ]%�*�y���j[%��0�T�%��-�"�I�����5��e��%�$e\+KJ#��\d&,���L�g�Y���8�B]�T3KnU�G|�^CܮZ5�D3l �m�=!F�v�2��������i�s�i����/�K�oc:����L�z��D�9�d��x�_��<h�{�Y�����x'��vn��#�d-ne�vV_u]5y�!f#W�2Ӣ��+����*�o |�I)�z��\m��7,��ײ}�y�2׻Ɲ��R�me�R����B7��Oa}#��fp�o��k�&~_��������v����ы����U��d�%O3'��M���`���2�E	��v+5m:/����:���;�^�Ly��a�3GIxt��g�{�l ɨZ�b�eeSk`�d�E)lۯ]��Jz�v��q���h-ǹ&L[��np�bյ1Ʃ�y��+��%�	p��V\��{�4���g�W �7�&vc���h;��f@�/�s���a4�Ȧ����m\���Z���DX���L�W;����x&�� �f���RܧT��)�xi����ް��el�K2�	���y�����h�ۂ�Q0q��zׁ"+�naֺ���o:B�v�Q+>޷�!*�h8<藭+���=��XH|��ۼF-�ٶ]�6�XK��u&��
�NNT/hZ�a�\rr���]x�ɚ}>a��ʍh�d����ٞ�b��,*�����t��T'y/���פrF��)�q]��1��1��4��\g^���4�:�5��6Ԙ�m�%�2�kW����ǹt}k��X�z�gݙ����%M��#��]�u7Y��)����BJ��l������^5�:�9�/�u�E_I=@��Okh�͈�sb��sf�����L��;8��� (�r�%��]�i��K>V���y��MsP[����!��@�IC_�_|�h��~�_(:w�v
�eKW���v����g�b�J�5Z��j�@U�x��D-"q����,�xА��4�Y����Z��/E�ܬ%5��r�^Ѯ��R���E�F0�ƀm�F	� ����B�!W������^j�"���ƭ��Z4��hZůy�vӺ*��˄�]�zr9Ow
�_w7��fאּ[L�)�<��+��'ك736(��(�]G��Tr\r7fgWmp,�BV;ڗRm[|��{��������=�{� l��͉B�,G?�궂��eڶ�Q��'�`C�=���z_�t�8�`����Ά9���$�o�p���n�OO���v{���t�NӛY���c��c4��\3�s��Uul��5,1��]@�@C�C#͙=5,���_|�E����c�窢����zB��,TZr(�-��;t�R��� ^�,�1GB3z[�~ބ�f��L��|1L%j����hYʬ'/�e<�\��Q\�UȜ�ʱ�5bɈyM��ÐR~k��U>~�^P���6���̬��z-���,��[�o�WX�Q��V\���di��Ѧ��%LQG�b6����L�/gX��U��
Sok�,��4�hm������,*����'UR�7��M�9���~z�7u{$ �;�i�R���I�O�lK�Q�(݌�Aۅ�K[�/u�+�w���RG�jWc�0�s�s����<��Zi0��.���y���
w�X���¾E�K�������D�S�����8M�����>�M"��ƌ8�p{��|����{�ߚ��W���4O���2!}�4n�ʯ��\����t�:����}̰L8�qWQ<��QA�f�bg��ꥮ݅�{p�Ʀ�(�eL��B9��>�HJ!�.�[�b쭸:�4F�u�}P����6�>Ǫf��;�� ��ws{����x{������h�|�w��O����{�ƾ*u�)kZX�x�X�z:�_m�Ưߏ����;x�؛��d:���x���1gr�;��z���杻��5�ȃ�P�Ǌ�Q����P���˩��h^E��;.���}U�@�ԛ�#���JLdP��tU=�e�o��V�,Ή���}���\��8��@t�j昱��VZ����nߟV�}�<-��ڴl���=;Is {n�K���U�{��	��h�ao@��>yʄG�K
�A{�i��g��L_\`c2�ƎM���]K7�om>�"˚]X�KgR�\�ֺ3��։x��. b�X/��� 8��Y�ٸ��j?��l��3b�2f������U�Sl��,�(4�f�q񫳶�B��i~���k��`���F�Ô�6j-"r�5V$ﮙ������|�����ע��Eu&x��ܵR-n��k�5Mm��&�W#�QYB��jƑX���_K۾���+*3nP���\4��s�����t3�l��ɯ&�Ч�r�N�i�dp�ol��ػ�[[q.���7�����=�^�G����{S������d:��,܏wM�W	���GB�:�nq�vOu��1�p�6C�.��8m������A,8J�x~h���NŻ7LZ�ח9�
Z2	ڸB�Ƶ�kh�;�h��An=ŵ:�������J��J ٬A�{�'�ffӋ*�c_m�Ñ]�4�c�m�8����m^0�9�s�������Mz� �0	]�Z�7o(*����ӫ� �fl�>��t<)fu������� wۖ���)h�T�A�|���"*Wd�y�n��WV͓Z��t�����K�{k��af"���b�f�9�/�Gyv�dЫ8"��AL`��Q�@��/0�o�#}�gKnZ�ؠ_P̻��3��È�{�њ���C����.U�kXx\��7f}���խ�����]�_�(1�����-(�z��+��鸗VW�Xp]C�7Jﴼ��4�T�}�b\��e�˔��A�yQ54��S��;���%F�:AGr�Y�`��Ý���<���`x�b�a�Q5D)f����a���eRL�T�4�pAfԮ�G��v�T)��L����C�k���ľ�1�]�I���_ە*I����ܤP_d�O+�`@��c��.���V.'��#��`S������)��EV����@ѐ�R6���O*a�n��22�k3p�z�Zh�$�Uʚ���8��[2�v���|�)}7k]��R�z%�tz\�� �����φx��2�b//�k����:ڳ����>��۷��Y��-�ʂ�CEoR7���D7r"R!����9���R5,��u��N4:k��;��0Ifm���)cd���jT' ��r��ƚ囁��Vf[ޙG::��p�{}�<�J)[J�#��@:�GN��(Q������q��&�R�<�i�Uj�P탵�-��[�bHq��^s=5/�}�On:[Y�z> O��R2Q?C�Wysq��\0���F-i۵')6+��C�[W4���0�WƖP��F�k�ɹ���Vv鸒z޲�CDn�rM@��#�C�_U��޾���e��N�IN��{N_[��6��,蔍󡩐`����P��i*��#ti��L{�RٽD�!���檑��'m|�DF]w��	]�Ԫ�A��8��R��sYe��1�j��}�q�F�z4���Y��Qm��a����i���_9sC�	�!dGR�ܚ!���,��y(�87�Er��̕�m�z!��D��Cq��S�u�k���]����f����19{K/��.����b9B��l���N���T�m:ͭ���7�.����e�����������$��kY[�.9)�n�Ȏ�f뙮ڥ���Mf�^j���ʏk0E{�5�����f��/��zrݡ.[	�y�\nX�Fk[�O�f�f��uo��jI��1fi�:���m�^�ڽ���
��گ6�b�`��#��u6؍��C�s11j��lUE!���F�����)��b��
I-:"j������Av�TQ�D�փU��l�DTL���F.��Q1EQGU����*���������Tu���U34QD�v4]��k����"�ֶ5$�Km�"��1SDP�MPSEQ�TTM53D����Qb
5TѪ �;�
�тji4{nê�� ���ѶtI4ED�$Q$Q]����:�D�5v0AA0i�$��Q���hv�EU@Ul隦�袩��I���*�����*��b""b�n+�b*)&J� �h��;���h�$L���ہ��g�Í�s�78�"�ss$=�JFJw�hr�8t��r6�jMթ�B]m
t�|cˬ�o�2�e�]ֺ���R�~`������Y-��%�Jo���������6�m��޿P"o<�^{�)NL�F6�`�B��ԋ����*6Q��v����*��C����;�%�J��s�T�p�Q�f�:f�AR�6���f:���d@�w�wƁ���(	��s�8����j�v���
Rr�9`]<�-�/!?e&��zTר���'_�w���H��J�~�#����=C��v��v��L�!m��P�����G�4liu�f��g(-����j�g��+h����o��:�{�!nw�Ó�s2���e�_*x��E��"ʒ];�>.�v�s�Ƈ������:���uލ�5k�n�iy�`�+`�D�y�TCV�E���
UK l(I��d�HZ�.�S���f�H�[2��)�N���C��&_�Ŗt���w���ߵ�rz4��lE�$����q��n����S��������!����!�y�c�y=2����0gی�wl_I6�:h��*�4�d�L�i�g��V9g[5ٕm8�H�Z��դP�k�t&SI��Uwq���5��Yz�H��+ʇ��Y���qD发~.�*��eכTG�f�#�����_���D�v�1�8��x�G�J��� <�b�)�@~Ŷ�8�g�X�o�]��c�T$��C:v�S ���N`��/�gd���:�N�������ֹ��3��QS�,S��i4w��;_�6.�tb�9\���韕���`�����Uw_}�� f��i�C�]ᩚs�І���7Yx��-#������n�?4;�`I��|���NYEzV��]�ӓW�>=>��Lr�O�^d̶�R��HmF1�+��U�|���}�>7>��=���U:��
g�E�j<����W<���'�R���k"[(j�vxt%԰[:q�c7"�j_by�jW
���P�̑-O䅘xY���u'�Jױ92j�ɲ����5=�X�ߞ���ܪkIek]���xi"�3�&G��J�f���NV��M�vs������M��LaUsx��;1���5ג�.q@����=�[x�ʰ�8�l���F����
��}s��ߧv>�c���wu��WN,�+��Qi������n.��{.����h���7�t�˜�;{�[���ɽkMo�!3G��P���䨵�0Qj"���IXE�c�1G����T��w�q�J7�W���%�k�B^'Ǣ�N�sH��M=y�N�=���7(��ǹ��I�q_Go6iި�I-2��yE%RUЬt�q���?���MB�ɇ��)��F�a����bKčk=��4C�r��ʿh�Ye�3^��N���ʷ%Y�����J�0��:-Ĺ�^ը8sl��r��u�<��袔�1�짧3��r�]��Fs�R�h�����o�F�>���v�>��%f}g(gT�Ĵ�.%���)�{FM/	����ͧ����<<>`<��0{;�~��}�=�������*�g>���|D��U�E�ձ|��<'=��L:��c8#Wc��T��<�t�q��]>{���v�<��7��\P>�z�-�o���2�7�b����>t��5J�c5�q�5�������]瀿/�'�H�|RZ{�/X��m#3NK�1�O�9���x6��9�i��⃛��ܽ��~#*��?n�@{��䞥m%�_�*(�f����#��R�Ӹ��~�6f��������oK�ǍiS��{�-��D�1Z�ԗN19E�=!5G��즏vc�5f�!�N���l�e̪�;��ܛ1|���	��)�|����겴�<�:X���^��s����J��Ǟ�0ˁi9\Ѽ;�'��m��tu�ƀ)7^A��r\ccǤ]�I�i�c.�R��:#�h]
��|�qn��9���A:Kը��`�+o�z��5b�f1A{)�i׼�G�g	�%[���;n��o	��˺�F7Hjk�9�.z�Ȣ�cнJsV�um�
݋e�OU�Ur��� �o٥x�Ū&�j���b�D�)r�W %~�~ܞ/6$1����@R�Oo�G�����T�����G2����;�x<ַ�[Q\���ޅܮ/&ɹ%�3W&�N�/4BKKn�F���z�k:&�w�:��8N�b�b3������#�)R�)hO���j���m}�y������8�[�4m��M�KpfR~§ț�%�5�3$mr�<�N��X%������2��F�}�1�2�o)E���N�<���J}������?j���{���f�Le�9r�t�z�@N̹��Cw<�[�y�i6M&�jSa`��ZJ�nCN(=k���)SfR[a)X����j�
\��N\�U�od�,���Bډ��h����Ϲ��p�*�p
0Y�0������g�;�$|�����}:��o1N�[��u��Q��B�+c��8��ި/V����|�G�i�Y�Aށ1����U�������*�PԸ�W4~�;��|k��M�	�C��cq:�9	��t*�lm-�~r�M��v�3�\��6q���=�"	�-}W4�:�s�&�8�g��3�骒�3����%7<`]�t��A�N�SG��pN��d�ix^��i�1�iK�5Ne�0��V�o�q�0�l7�~���\��\�Z�M��z?J�.*k$��v�y���a�z8���Ë9_Ig�L�ֺ�f3=�YЄ�*�q��� �n�[t�V��:gC��-�P��[F�oJy���g8hk��dF%ay[>���m>pB�7�ڮ��(�r���_&+\�u�ykF>���{w��|�����P�w�_?]���.|�7�=L���r�����c�菱
]���T: ֯��v��@�y@����������U$c�eaCr/�KB�o+�Z��(y*e^E�NV��t:�Rꑎ���:۩�J�w#	Lo08!������t%ŵML��e����Ђ����+G^H���y��mn<�i��z)k�j�С���2���8KFl׋W��w(d����.�����UУ�'TU6��e���pƥ��28�|�I28�S��~a�}2�s�Ʃ���Ê��j0�Rv�ڎ���h��a[�ŌP�k�d���r�c��*�7_��Hy��+T���k�E��M�^rh��7կd�B�{`����&i����uf�!��ŵKD[O�J�mk�yθL�a�")��v����{�U&�sP��$��)Ӽ���j�m�
���aT��ꎑz�n"��fK��b�9on�;�1,�����z��r�Q*�=�D�2e|Ը��"�%�u!}�AK��p�1�Zj)h�]�,�/�DD&�b�[gqQkkR�jS�
)(�ӱ�3�hh���z7a�CvH��d׿f�3A�'�2{�cs�#�2c�����t�S]�*�v	2�Rt..�+���i���*~����ԣz�q�nV�I���x�'ncKrG^��r?��`�]�����j��ԛ��򓔝��n�Y��X�(�A�������ߌ,J�^{'w����%}|��/���8��>xK�:hhmk�ޫk�o%e������^�u�.c�!�4��<v0e���y7��]��8�������%����´�~+�Q����������f4V��5xؐ���9;�иM��f�+��(n��ɋ	��zB�/���bۉd��2ݎwg6�`[J"�޼�P�@�וy���#��2q���f	�O]^�VoC��ڭ{���]�)���-�X\��w1])��<!���,�)D��S��P9�gk;��pA��I�C2�e�MF2���4z�*��x˴w��i)^����S�+7tt�����t�bo#�uoFG������X���'��q6è-S^��,�(�,��VK����|d�	\�h��p괤s�NN֑�(�~X�I�����1F��w�*����-���Y=N)�}u�sTu�,�K����ei���L���Y��c079t�&�Z�kt�_�z����Mv7NPz]΁QE�|]��-z�ǻ*u�ȫaza,3�+�J���F���V��[k8��yǐ�w�*�'ik?M8���*�m�R�����ޔ;����My��<�4g��[���&s�O�[�6��
�HU��i��������*Oe䑥w���\BG�Q��r���h,���XULYA�x#$�E��?$�����l�?�����%4�K7�ן_��}������&y��Ip�r�N��ӓ��^еX�Z��=x�{*�� c�AȳUb!��l<+�.�U�2��l2~�\k6�gk��TZØ��E�q*����:�H����1��ﺋ�������o��!����ɲ��ۇg*��M�.�?�t��-�jA;٤Tχw"�"1��H�;&����Ƃ�`�+�2�]�mЮY���0��4���MǛ�40ev��z3�d^�d#��ڻ���Vp�4��5��بi�S��i)`���)H�=�Be�`�fh[����"�2�a��4�[>�A����4=�a_������u�P?��y��ƈY��";k�����e�+��~	ujzF�U:��04��A��'[�0-
�t7����YZ.�s�)d$>'4o���:lsQ��i��5�G�]/Y�D�e�0p��<ik�����M=��ؗ�_��k~��l�b�G��[�f��Nf�R�����ከL����ϓLTۺ��9jYˬQ-�A��}��H��g�X��32ju���*6��f�-�jZ)���5�L�o�wUbv�e�n=֋�}i�OuE1�W�J7���SjE�s�KD�铷 ��{�w,1�[t��*�6:�"������l�|^��q"���'E�B!�}Q_Y�e_�#DӶlWa��	���wE!���yݚΘi��h�;}z%i�Xm8X	���X�,H���C��?o�^�׷�������3|Uӳ���9��6��:���d]	��!ȡ%f�i��sk"k�s�N��-�2�'^��E�/IE�N�GZ��ݯ!��pDz�P%��@�nS2?FWt��E�
k�^<�`)[7��=�C�y/�\��9V0��1d�<�C���hŧSd��-�s�kM�^M�ۊt��:�fԻus�lj�t&\��)?^-�{`��qvm;�vԭt��q�(���s�h~�Cx�e�Z��\H��f��U�[=�&�_�̤�Tyw�ٯ�-fP��$�V�S��&j �K� �Od^h��N�^�@�_��e� ��v�{ʕ=�0��	���m������Qh��,���/��W"u��&S�φ.A�E��+�k"�����W��!�~Y�_n��{Zơ��&2�sg:
��x��O�
�}iMU��e|{c��U�s�=��Ge�Uqn�V7i��T�p����d�Y�3�$��ϭE��ن3O�F�T�k�T9d��R2���&�6��G�v���T�q�a��ԣu�X�%�֘}|��`0a圱
�}YWSlm�=s��Z�(��g���Q��6����O�5�ڂ-�ߜ�2�H����ek�ڽ������&K��v�&�6�Zq�`Wlx(3��v�bjz����{��/��b�+1Tȡ��`޺�\2*5���T�Y��:��{�x7��<�o 	j�s�ցq8�>'�	���
���	���N���W������	I����S���e��1��)�r�<�����^x��9怗���2�?oW�$�~){f��ziG�c؈۽��v��e�5*(K���c�v!�f��W�ΟZ�`L������
R�����g����xO�;�*���FR�=�D[:�c4��8�-f2ZP1,��B��!�gkԧK����F�k�f[WL����"�k�Jv@r��r�G�Z�)V0j-�<��]tD�^W�K	l*/_ga����S��nl�,|n�ٖ��2�P�m"�D3~�H,��"lh��ʿo��]����?7��S��k�Z��RSu����8�M �+(V=�X�*�e6����d�#��|����Z|`�כon�^T�O�HeV5��K'61M2�����ৱ��.zg&1�i��BU����p0�Pf��m"���5,�{�1%��˔�Ǩ��8��k�;���Tv��~/-���aIFd@�ƊO^���p�0.z�5�M�u�j�nS�����V���/�����a�u�I-v�]�ƽ-Oeվ�s{mۤ.��e���s���%ZPscN9�oS�uk�s�;|�5
�9��Jn���`P��2�s��Z
�o����x]QZ��9J���V���]��n��ނ.�0Wwϵ����y������,BEJR M��`6��q�1U����:���
���>�v~��-����?�e�0?}֎��*��Y�xZ�՛�S0y�v��us
%�RS��(�5��ʹT�~k
�1!�my�<d�u���j��M����^t�^2)�q�:�����ތ�t��9�,��=.,�N]�5��0���c��ӱHh@3�x�,�&	��.���)-MC0�p�1�ꄟ��AS��J:�T����󵧯S�s�{�1����Gϼ�|�,��C�과��]%���
�B�zț���o�%�y����!��.ʁ��f k7^m�^�𾁏I綺�7h �mV�J�xc�X
�ϥw���JB$�:t͗V<h��l�k�� ks�W�>y�n�7��]�!ue���ۣ���4=�w*�=��1��zFf��1O�!�9��,2����V�j����!����K�_Efö����}����a- ����A�t��שׂ�Sv�g�9���FD���<�v��T�MF1��O��o���wN�K�}�e�cj�����|�O������^�W����^>o?��S�|+x��o��ܰ9�w:��zR��3(��Z�uq�w�Hl�Zx�J��ՠ�"z5J�;��,��'XB�R��g��su�˂��/��麩�C�˩3�Pֲ����"y��K�=]p,I��fn[Ns��#�QEw�*�"o]c��G��f�����}�޳{�!-����+�֕@��g(��%���N����3^S
�L�}\/qe��o�\h���T��̉�᪛7[�&�J��s��:f�YI	���*z2����w��LHE)QF�gj>��R��wC�Y�G8ե#?9��v4��X��.�Kbk�:ƭ��,�
f�718��"��ƍYk0�$&�<�����Iije�s7^Y&����"��<��܄�67�L��w��2��j��6(Um��I���dzr����p�cI����a�z��@ �Y/i����S��E�;,op�7��r������Ź���CS�w2m���W1��/7��0��'L,|֮�՜��`�Z�Zsd6qt��h2��/e�//3D��k�Ds���M��9�Y��Y��vjUp���#xT������E3In�_��5/���7*%gfe$7�ILj�R�ղ.71���`k3.5�a��k�1{ݚ�Af���'>�Z͹D�vd����-P��#�Q|�>��2G�[��غ���7�E��k+j{\C��8#��������BqkNA���^Z�V.u��Fuc�Ni"X�t�m���ռp�B�!mJ��x���ۙ���kGU����xخ��x$X����yP��{�=�e߹]�c�I;��e�Q�ښ���Qf��%���T��p�uEf�Zs�֖�<��-1R��-徝݃^�}���v���9�p51���E�D�v�]�ePb�����58.�
�Z�K쵫�����	���kdCw Z�;'
d]�Ƅ��M��׏'j�|6�/�*V!��nWws�N��T�vXW��tw�+io������d[�e;3�B�[I��=�,'(�ڝ�L��3��Wf�^9m���:�҈�E��cýԈ۸5���CfI�,KR���3,�r�rB$�C�7��$v�A�f��V��T�mdyc �0ͭ�:�����U�ԟ}��;��./-[֞��]�Ub�ŇPt&@��̾m^޲�%Z9�TiPw���b���Sy��q	(s�BMh�d�G�Κ@T�S(��j�YX:�<��mQ��(HәنocZ��7��ݵחr�˖���g`|�@��E�+�H���0����Xt��]�NM�F62��vG!�;&�[}�:��1yx�ܮH�v�M>�/ ؇y�E���a�gWR�G�}�辎�B���oD:Ma3c���S����	�qn��,D��ݤ	�=�v8:5} �ݠ���sM4�*Y��m����t�A9Y�#�F ������XuLVH����MU�cS8ء�"�&ۻ�DD����"Ѣ��h�-�f�1T�`����;�Dݴ֨�4[gN�6Ά���`�����5���QLD�&ؙյ3��EkUEtwkX*���2�P]b�ю��Ӣ��4uct�h5�i*�bh��IѠ�`�KDm�h���"(��&m#���"��M�wsq��5Fb
j���)(����D�1LEE�,Em���(�c3m��4∆jX"�4�h ���U&��g�*�uEUDT�X*���f��������h��f�gAU6��T�T5E4��P��EEUh14�MCD�m���14�Q::3TGK�
�k�?^����p�q���<B�wyj�qN��dn�U��:t��vh��бN�#��p=��=��MM,�K$>�|�c\�ꧯ��%�����(�o��BS�[W�m�H�U���<JS���c�sH�w5Fi��y��r��q[n跇��X�b�{�.��(�C��������i��YM6#bc/�<+|<�x��nmW٠���z�z����]�mr��c�K�U�3ƶ�rڻ��4�d�5b���.��]��)�^IV��yE���L/L+xLր��Z&Y׭M�i9�X��z�]�4bvŰ�G�gQay
QpΡ)�JUڵX�Z�q��{�ly�]8*h�D�˲~�m����h���p��nuC;obTX��@N�Jj/�)�������設����Ucmue��׬^�-�TO�T_�Zg�?V���*��ju~O�1�(lD������4cRt`>lX�Գ�ݗ)����j��xk�\S�ތ=X/���_zy�f�on1=D �N;�ej�K�*v�Y����tk����*1���XC��͚B8�v�a)=R��q{ٓ8��wYH���y����֭�O[���|[M�)O> �fD;5�9��w�;{�[%�Iu�A���r[JM��g�b�*����q9��޾g�!����k��,`���u\���~!�xo��7�������w/İк5��u�:��*��&��
ܘ�4��*��U��[�_��t��%.����aɝC���z6�C3�o���a�<��`�������%!5q�='�gz�X��q����V�C���=��yO�ex�/�$���r�E�3f+��j���jc��G����`���ϔ��^5�3E�y͉} ��|���*��$[�0S��� ;@Oe��1U�lc'v�#�3u�5hFk�H�u[��t�����I}�����QV���PLMP,�O����|���̔�n��C��,�����
��P�k���~�KcY��g�3pv[��Bu�a�;�W�fe�v�/Wd���g^�n��������u�/S���7�i(>�i3=Mb��[ ��)��@�H1�)�_7�O�n�ې�;����[྅���E'�+*Z���	kϲ6�M��xp|x���߅ֵ��<e)��D��dy�Lk*�-�}Й��)?X��풯��`�a�[kSv<�@B�ꪺ#*1v�'l��or��l�E�f9f�S�Z�uQ�k�L$�Ty>�)4+J)��[D�q+[=�TN�v�Ź�!F ����g��C �,�@N�]�B�,=tMwpy���j,�3*󟚸�yO�b4D��i(9^���!��{e�.	���2���/�����ݞ�R�I�老��0|	�%��r�|�u�=������e�fM��v�(<�����j���R�PuzV9��Nw
/vv�w~���~$~� ��^EM�ĭ�������ֵ�;���W��b;��.5ʛxc_�3�{�q�<�����"�B5S�)_f��<:r�`�*�mO�*S#��m��c��ť���i�>����c�yu�½�d�r��n�Xe2p�$�+�N�q���Q��g��0���>�m��2�n���M�Rڝ��������N��|s���gjvoO'���,��>�M���;ו��#r1޼��3��"8/3�h}���c����S��ޯq8�jFbޓ�=/*�mjP����S>d���Qqw"�	�����(���M�K���^ON��F�-7[VFRa�ݬv)��̧��X�5��ѐ�5S�A�Ļ*�;��~�ه����H���7�w����?Q��W�_�_���z�jw�JU�w�iuc��Υ��DZ�Fq*p������~Ru�����Z����l\c��z�cH�3�ػ1zKH"ASl���U��Z���;_�?�Swq^1�`D�
gy�-���\.ȱ�ʯv����-~*m��"r��X�}��N;
�'�I���|���8�Fg5��:^A�B�J��d�q��?�/֛�j�O2v�D�d\7^��e���i�G˹G�w�p6jl�[����^n�`P��$�{-v��Vub�g�ज़��g�Ib\1��v�˙ ˂��ŵmGN�M��6�5�ov�z��305(v����4�%�RZ��i���F������4�M��G6�	e
ǽX�*❷����o�����ͯ��Ii�+6`[���p���4�'ţսJ�2~�SLo.�[�����.���arH�_N�L$u�m���ո��HCG�%u���=�?n�#��[�gG�����G.}�5���9�V1��8�R��B�\3cX�r�這s��[j�͞�T�_{tu�AѕD���NXX*��v%V�^����^�j?1��v}��R:w	��爮{��J��HRօ@M9�<���"O����8K\�l[���1y��E�*�N�f��!�5
�C�Ï�z"�T�6�PȖ3��Nޑ|KЂT�rA.�:����Q��AA��g2{�#���ó��ر�.C�.!�����T�7>�4w<�CPYaE Tsv(�X#��1Rc&����{2���W�6�x��=2�)���(t�ޔs{��.~~�������龕��]��F�#�ЂUXښ�ۋ�k]�d�c5�}1��}/�D�0�O���G�=]�}�?=H�u9nCl`yt�Z�k�|�)�>�f>�����M�r?���o�(y�b�B�lq\��u���'Z�Y���X�Ho�b�yB�'[�j�P9+9��]�[l��r�
x�q�%���p�ҳ�眺��ʅnKT�a��±�U�ww�]��OL$�W�Ao�Ц���N�݌���J�?o��ׂ:��;@��D��0�p��Ӣ&��U�\�t��:����t�y����}eހ��4Q����a���C�u<3gKv��욃[;I���u���>/�]c��C>焜��M"�5���Y�l%�X>*m8z�t���7��z٭13��N��U9Lѕߛt�<5.�7�wsv�Z��f�*HeAv�ɲ��~�k�λf��]��v�������r�!I3�G��LK<�du�ǣ���^w`)v�\�-n��'C5:J���vu�nr��ʀk1|�[�D[C���Pi� ���\6��ٺ_0J�u�JHnk �2k��������Ʃ�x��2�0D=c��d�4VG�}���x�殕��{�b��q��������*T�l���=ߊ��֡�ʩ��"��P^���S�/�R�����?5�����xH��J�X�R����u����C����A�f�=�oԾ�F��+����:E��>׮9��T3��R[����'����]��>V�7,���W�n�WDXy��V��W�O(�F�����u/�1�SX0����͛�m��!jk��%�x+U\YcaK���6�k70�����"˶;���9ִK��t:��H�&���P|�F��5R����p�W6�I�)s���ܠv�҃0L3�}��4�Z������VPv?<y����	xX��rG���Mnsӵg)�&�Br�-�5��8�ͱ��P�}=��Bl$������4�[�D��E>]���_}y�6�D$���o�8fF�KO=�d��}u(�XHv�֊�sb��sf��>]uJ:P�)�7����G2�u���vyS*�4��Kn��i��)�LAl�W}c�r��������V#�Ћ�W�?|e�q��{�粹X�&u8�H�ƫ]!����^��r��0������F�*������;Ϗ�^�Տ�z~�a;�%ǰi��kT�fuNz��껇�H����szd惽c�b��r���m8C�˽괺����FkXd{F�I5��荄�q�{��L��Bv��ܮq�ޚ糢�~��`���~bOҦv{�x�w�*X�m7d+2N�i�s8EG3kב��Vz�Q�9���a�li�F�V�TN�OR��-�	��۪ME��m�,�BUT�Z�C�*d\����wF)����Û5��-����'.�F�@w�-�k�z�(L�fFꗢҳ}w*>��w���8" W��Ŕ{�jn��JFf�������D��8�S�����d��D���5G��z/kR�R�u�B\Y��W���]v�o��-Ц���<n�i���H�v;�%lY��{w.h�!��<�ݴ��+��c���	��_{�o"�)�����c�e/B�Q}��+yM���q�:���N���L4+�� ��P���,�^�)�d����Ħ��t˜��O׋h^�9�*�N���a^F��	~̈́�3�ؔ5���ύ��?�1;�Y\Ũ�4Y�B/�G�u	��	K?<*����t�m�F�F�Ɍ_bԄ3��}*���Րx/�2�����_�u������&��]���A<Sw?%�]t0��Ȋ�?6[��߭�^B��T_ɪ\��=��ck��-��itx�E�r�LS��,��4[�|��#��iS���e|zC�u#�vV���m�[ak�@�R|�8/�q@��Q�Ƞ��!d=3�.��-�M�z��}/|��8���7�Ƅ��s~��E�`qT���[���w8��U:�زHՎ7p|R\:�#U�f#����:��LƗ7QL�GoYoY+i*{�Z=<ز��3]\��b����Ygk���J��*.j��A��%��>F�4kGW�i��U�@��� 5m�6� vU�g߅:��c"�7n��֢�ֈ�ڇ�����A��k*�o�R�:&��2弤4Gڕ<�1^�����>�r���lN傀��Ԩ��qU|b���z��TN` �3�Fi�ݑ^L]�$�������{"�eCӖXw+jcjܹ�*��,ë};�Qq�o��Y���,Ƅ;�@f���p^�"&vp�3'�xь��c�-I�]Sq���/�;,�F��g�gY��AUI��hu^�}s@D{a�ȉ�9�)s]��!�7ܑy2W<�b��7c��9w!�A-#���7(������l8sY0������t�E���n�����F5�h�f��K^�c%A���9^�X�G+�a/�����ι��U�����О5F]�"��楟=��M��i�v��ֱ�D��C$�e
w�ċ����E#�߿~�vt"p[���#�=:�T��x��8��μ`�,���n�S�6��l&��/K�٩I��������b�p��v	v�
A��*��E3���
��ss!��0C��7v��:��z�V0��2 W�!��65�v��}���zl�6[e�k'Pz�a��?��x��;������{OO5��u�P$.�~�T.7Y��L��\�v�S��ي(=2��sJ�>x�͗�M�|
����z]O{m��B�`Z�j�E�"��pdµҷ��jL<��F;t�?{"`�}��u�9�ٍj���ݾ�o��N��,}�ʣ �'�B\�u]̨�bA0��Jv��ً0���ͣ�Zy��]����$7u�w��U�I�|�t霆I��_|�2"!>5	�muC"YH��p��^i*�=��]Ԏ������ՏYOT^id�w�7@�2�=/���og�e�}�J�c1Ja�q����M��^���f��ầ�-[p���~����g�%v�A����UԚ���֑��V��uc,�y�k;P�}*��r�Kԫ�Ժg[-��h��34�ށC��*Y�_a��j���^�+!\�m�KC;y�[����'_3�Ϻʡ~�5��S�ӽp��Y���5����l�u��F0��n+u-�����^�;c��LL�nk �_;��4�/^n�dMmؖ�i�׭�ܾ&��`�#�W��<$���XG����smZF	��p��9�W�{G�]E�ْq�$�����έ"��#���|cw��̪���4�<T��wv��wjg�l���p���2*�C�����@_@��?�d�4�p�{"e�U2:�׹�EɄC��ԅ�V6jky@��m~�gY��1:�FgL 'HdB��H���nT����^���_�V�vZ�K��)	�X9��2�j��1�J��l��r�L1"y��ͭ�m::��V찛Y��Bq�#q�E����^v���.'	���R*k��x�S�Zpe���3nS���v��ʋ˨s����a�T9�ɽN`�(\�E�@8�į�}�d��q�=�����ć�y�ɩdK�)O�ݻN�P�9lf��j�Z��O��ݥmC2�	u8�ںh�d�X���\b��qh$��
S����N�V,`�>V8b/���!ynE;�T��m�2n��B�\[�T��1i�]"�iU�ƍR��`ܠ�Ͷ�nGeB�tt{.����4z�C'���3F���;W%%��\���}�۴ĭ�J�T�d�c�ѯ3�G{z�lVR"{����C̯�����i�2��]�nr�`
��z]/	�/r�Yn�Ȭ�=��<{��:5���	���g���n��f��70��?-.���>�t�.l����ܨ��lO��%��^���]%�<I�7�����"˼�V��.���w۫K��"��	à�ил�L5lsAr-l�옞m��|g�m~Ȍf"'	��U��V�U��r�ܵ.Ɣ���\@�q�jq����=!��Uk���_U���+�J�I�Z0��}X�
��T������u�G����7s�3�@�=˾2Xn�����x��>�O����y7������Q��V�T�k6�ݗx��n�pJH,���0�E�O���)��Q
��T���l�jvXO�M�f�w]w�O>����gy��7�Yr�:����W�p��+�]r�+{���a[ԉ����b�W���
�S��f�m�C�2�3���A����U	hB�u���lL+).��H#����}���Ӟ��uB;__�ۺ-����K�-cXO'SjWN�	H��9���C�2�w�Ү���Mf�L��[�t��'�y�B�u�&S�j�s�l�9�@�+;ZD�S�����X)X������P���sxkdn������[yk��S�r���v��P�����Y�O[�Yo�ڔ������M.�7iC�b+0;&�%v@�}c��~�ދ1`-�`j��{0��p��v,��h�\����L53`����ūtOu�a���ԫ�V�L���6�6� �����B�/��Ml�-�ǈ����y-l����ݙ�&�C(�kSء^��lm��r˧���Dl�ш;Ly�;}ϳu%�/��C1]�7
2���k{q��C�V��f.�}L�����ϖ�UՁ�ٴj劢V��b�v����Zο�Fd1i��aM��jڜ�24�Ճhk�!��i���S!������s/ɵ�P�e��Cۙ�c�uJ�21�eCeW"ROv�;�/�
w����VKR�t�㽷�3�N쌺��:(����)]�߆w-�KE^wG���clFZVl��<�Z&M�Wh���p����ˁ�!9�qt��n
u��(0t&G�V����C�BY��}������STs/Z	���N�{�1��"�} �pՊАJ�y�"K�%Ӿ	w��o1b�g7с7tÔ�Lʻ�g5�m�Ų��|��et�+�Xu�/]
��X��=Ǖ����cm�c�hM�`��c�����0�5�ձ*t�U�f�Emçm�Й��AԝI��bs�CR�����{X�<���pம��6fk��������A^-��-�޿�����V�hGkk�Zr�%l���6W]ɛ�ƞ1�UD�D�����rU���mV�34��c1��P5�MI�ՆX�t �b�6ʥa�����ײH�J���pK1v �7l�8}�vD^�u[���*oXч5	Ln��M@��S�CAǥY�R�f؝�c�^h�ޥH�̱��s7���5��r�$zR4qv��e�_���YOk����nC��'9�f[�v3n���XC�-H4�2�ͽ�hٻ�3�z�c�^���5���+��Y��42�+#���X��lo����/��b�Pa�R�;Vʪ�k�s;�n���-T�m��]��%���L�Go0��nV*��p'�
4m���b�v]�G���x��܆ʥ��	��� �AFͶ;��S�b����6L�U�*�� ���
�P�D�u����b�$�
*J
*6��4�5PSQ�AT�%D�Wl]uѪb]��V�!T�Ɖ֢�����ڴ�MRR@ECUDl��#�/oc�PL��%�Ŷ������bJ
)�th�5�f�ى�"��:6�hh�4o,'E%�JZ�R�V6�LU�6�*��ڪ�����Pht풊Jb|�*b�)+N&&%j�����TA^F�.�PL�1S0QE�h����j!�&b"^���X��(��Z

�6�1��5�)��*��tQ���*���&$)�'N�mӫ�M%�������U44�T���C�*j��f��4U,OE�����:��TTN���_q��|���J!�\�mo�z���w���S�;sP'3b-�+����)��wi�p�f��5S�s��A�;�ox�+�g1��yn��y4c�#Gm�棂~@��K���h0G�і��rϞ�3�d[d��p�t9w�*�[_u7�a������~�}����A&����}ф���*1�{�]�i�u�j񈶄��(���Q�0��H���X��N ���zޫ��x�����3�
�ͪ��/	��]"�掠����MP+��/~9����>v�/���|ƭ�s55�}ql��l��۹p,k��|T˵��k���B������Q������s��^d�/����f��J�m��*��P�_��e/צl�`
�N��X�-����'I,5dS���|��2�������o�%A�C��FUM<�����L��yO��h^���d��;9�������#n�T���+J��{*���o(�������ڗ��?������y&1��ZWN�v(���B��B���e�㷲���Z=�X�E�~�c����'0��Cu4m�4�F>C�	#�w:�4.ٴ���x�K��z�h��$Ԣ���/�q��#G-��~c�89�.z{��)�^<�	6s���f���������B���M �v�,<G�U:���e?��9�,�3p3�,Z��ؙUm���T��V�f[���|�Z��{m١N�=�w��sxK5�u��lD���=���}��Mh�>8�:h�3b�_vnj�v���5{v�,�]\bysl������x̓�3y�E�Q�˗��
7x����Îc��<�ȾM"�_0�Z�ae,�e�߈��^8AM��<�3G\��֩�t�:w�d�1���D9NMG���
�C�^[��Z��`�,"�r������S�d���E�13�!�v`� ��y���^YX��-��ņ�*\f�e�#iĵ����~����	����y�>4��*��A�@�:��@���@�ۚdǥO6�*����e�:�,�ݾ=q�x���i|jt	�gףU%�Їc��y�N���@����>XG1���9]n��f�`���E�9��?_�������4�/����^w_W8V�S��2#[��å���꣹�Ϯ� *��}c�h���_��+}<z1c��A�o*Ƅ��~}�e8�ïyp۾��٧u�5 ��D?#������WW�jZw ����J�H��5V;���}����mM[~�<2>��ܤ��V����m��\sS�][u�[�/��вlxOТ�]��ԝ��'�X��4���)�9RX@�+6`]��A��U��}1��������P�?Y�����q��JU���OB%�o�s�%��]a�F�*x�W��V�C�#iN��rXA_j�����)��4E�>�O1�u�i!��	'1��С\�շ�+,�=���éV�PiDh�Zw�gv[3f������+��sٶ��y�\"ou]%]1%�J�*�XYYF6k<R�CBk|��J��=��o8�> W��Ae��]��8�m��]c
J3"�uqA���l�ۋȲ�YZ�\}7���8��nՄ1�c��,�P~�(�9�NXX*��r*���I�71la��TM��Έ��S?h��o��=莚�ǫ�7f���as���r|1���G6�J��|��5ª���;[���&��MB�"�os�3ak̶e�S����/B+��W�Q�D~M�25/�:����������C��,cD{P���Hxa�iM�c.����KSP�C���SӔgq��Y��݄�n[!Ae�P���x���}e=	y.Z[s����_*�nݳc�V��%N����eZ�3T��j��.Ļ�.���ra7�L������tj��Z��ֽ'���9���ւg����S^�8����P�=�f]����M�{�O��,���1%K�{|/�*׹H�L:w����`�=%yP�v L�����+�d�J�`���I�l�=�N���Yi�j�a'�q�)�v���I]6���\���y�J$�,�U��xr��}�z�L�6Ɉo���Y�U�V��/'�̖���򡩷3#y�蘑��u�+J�H��DU���E[��穷\+	�ʻ��Ϯ1��ř>��S�H0j���T��Wm0gv�f8�l�ZA9j���Z��\�q��r:\�h�y�`�=����-"Ό���)��Q�s&}͠VeU��x˷@!f��ע}�+M��.N�ҩ�����TDi�f��{��q����o�	�#��ȽMG����i���Q�WH�_n�������6�y+�l�YN�VżD��	�����t��bU:Ym�~�޴���׶4ϲ㐵�]���2iW��`qڦ�K+Z�j��yj��E5���ی�U���Z�c��s.�n�C5����}�0~;�h�f�a%o���7���T��-��sV�]����k��C�S��J2�G�v)�ХaJ��ӓ�u�)6��c�3$�Ѹ��17�-�dӈ�f�AvO�*9��9����b����㩙����%I�~�mYOx�Bv��p�=.��*&ۍ�C���L�eo�ܯl�2��?,���>e��^�s��3��Aѭ���7�0�)k�t9-�aP�[��<n��u`=WU������Q�>�x��2�oJ�(8��ɢ���x���KR�����wS3�5��V��_4X9	^�k�Ehy���i�vN��	k[j�:;2�؜w�:���2�a�[��2����u�u���L���zDV�_5H�D�嶗E�}WWb�b'��m��X"�RE"I���A���u1�����r�Kߊ2q�/�cE;���f��F��Q�7ȷ7K�ck2��2S�R�+1Լ�{��y;���0�[<�_�8��Nz5�=��)�E[2緺�^-��{�$���UI1Nю1aSkY�1�a2Q��N7<�˜=�Uc�3p<�u,�{��lrx��Vs�b��*�)�
���H�u	v����LW�ݹL�* �֮R�e�z�kf|mɮ}�@�kE����C��X9D������X]��:b�+��k�{^�x�(r|���V7MM3��V���+���,{Y�[�L"[�����y��zF�q��+���fx��x6m&�;�j[[�p��̝z��8=�R+�t�����8��W�/���z���&8tY�m��CJ:�K�qmWp��j�C(r���2%��M���[&�"a���_ˋ+�'��3�=,��S"��]/�
�}ySl(q��^��A�=���@�(��X�voI/@�D�ݜ�����vC�
Դ�d��с�[x(��D�g啜���'���T��sҰY>#�۫3H"��JS��Y}(R�V���u(sG1߭w*�Ɨ^![4��������.O�֨ŏ<^^�56�R2�r#����h ��m�n#ݰvշu'CD�۔�p8�έ�J�L����ś[�T����۹�����J|2��]�3�ˁQ�]�򴯯eX�����L� ���h�{��1���m��Og�S�]���K�B�|A�#x�^=���'%�	
�%o1%���dS&��Y�:ּϗXHU��ad8�%�D"�3�v�����;jR��T�	�-H�|�r���<�2�ح�V���
�V=4@映����I���q�>)��l�c�nlV����X�h�d����bsj���x-�逛��G>ƴ��]�8ч��U�/�,�y��	[l��F�C��7�}�p1�|�_~Hx�m��Q�r�&T�2����c8�P�zx�Q�R�J���tI����l,T�°�
������|���-�b��׃1|m�E2��e�dڡ�ݙ���`�[��+s�vWE�Xu����{�UM�\�״�"�!dz��ٰ�a��Cv^�����ﶍ���z��5����|�Bw�Wlb�B&�>�r����W8��3\l��y�����.͌k���L�ŉ���Lj�T���@��~.-�
�L^�k�ΔS^�����v�w�y�=�g�O�]!%W��~�5�Y<E����L��Vz����g���W+���a�[I�x[x����<Ͱ؇)�A�SN�^\��Kp�c���|�n�\J��:8�θY���2%�Y��]&K\Z�#g�f&�Yˌo�?f�&��'�{��\�B���r����#3u���~o��x���ASl|9M�'眏5�+%;�Ƣ����f��{r�D�����5r/�f�SM;nAc/EB�iL�4�\��J�v��V�Wer�t�*W�ʈ�VJ)��,8}I��F�����:lg)�j�Z�T?N%�ȭl�3<���{�a#�M�WH��f)0��t	YW~Sl�#����"|Z�^�΋��aU�0��*i��d
R�Ռ�]~[X��^X��"j�����5?
D�`�����v���+'�����g�'�Wt�e�UL���ۨWX��|�x�	�@��V�O|�K3�����xF2�R�(Ǵǳ�13|%���%�v�3��:-��#s���uy��C�Δ-�4E4�t�]��dݷ4v���.-�*)�(�/�k��rS�͕"���m��e�w��N�NF�H�Q��qj�-�pݞA�d,S��RzA\���;��y���F�f.��Π�<�mj^I3�h�}�zD�����F�����n�������X{���Y�9�;%����4���m�2������r�ϱq��25�-���q|��"���T� ʽ����2�T��m>U(�.�B�l�EǙ�W�,��D��PȮ�Hgts�,ԁ���y*a�@�۸�9�v�6wVE�[.Cx�!=��������,WF�rб�]��1�q������}��Eq�;)�5z{�=��p�SS!�^11�;�_=H���1��'���`7}y��c�`��g8�]W&�j�wن����65m��r��ƫ<� ��s��%mC㮝4ƶoku�_�&����� �/ݦ�7�y��t�1=a��֙�G^�i��w�\:^0ٲ���D�8f/
�`_c�i����n�6��2�ڸ��������jٲ[l��ς��%LM���y� � ֓�՗}����w��5��O2��l�9S��ŀ<d5���	����E��,ʵ�4nM�L��2���#$Sx����x-e��Re�wY��g6�B���X��vn;��tQ������m�
�ad�rhyX���3��˪aE<��5]��tN^�y!�l�`���9�7C�R�d�zʬ��+���ɃLm\S��֦����:Ȼ��S�s-�/m�t�}`��ڪ�AK�>���Tnzn�؃h�:fF�P��a0֋����s_\�a�Og�g�l��[�.f�i�(�٩��_�$�\�Qշm7��p�#�7���5�к�3eLK���v�\e���=�m��Ļ7ov��A7I��n��cS���k�AM�|f�Δ���v�T{��m��Ƀ\�yG�.��$ܠ�nS\��/ �Y��U�N���:�ŋݻ����K��O����F��'�},�dFzנ���m9LaJLKA�87�ov�����GM�E�o}�u<��rC-2!��C�{�d�X��5�i�.���Fu]����e9庯�~P���|;��=��E�L���[9��n,��|�s�5 ���r+�1�%f=��m�/\��kTUFɦh��}������<��{&��t��l�O*6�]�>�ʙ��T�m0�Q��3��P2ƎlF�+2�2;W5�ou�7��x�{�r��N.W�����p�<��`I�6�`"���a=���t.�q#��v�/j�cE�c�[�X8��Q�Cb^0���,�nE�&8c2^>�sDw*���9�	i�����x�oQ]jTU�)Y�Ӝ�yr��*<��gN�V�iy�q�3|�3\����!S,(˛7�+��@yvܭ	x�f��+�meᴎ�oc&�MIFq�nZ�y�:��q��{WX�:.n$��J���&�o�~�R��nz�U{��r�X�U3@�N�Sj��"����:h]J��^(N�L/V�^a�؋��_��<�+U�B4�E�^��j�n�Q}�z%��t�}z�}W3��vB䷵J{(w���� ����e��^�*\��!��k�e]!�Z�Tq�;��JG*�f���؜��ȍR��V�NI'��eVر�:B�Y���J+j#/gXm�-�;7m�H��,cwl=~I-�NĪ�	̉�cB�aM� ���ڣ�kr�8vr�;Kuol;��zv�W�>c�畻`��)��c��|�v�q���b$B����Mz�z4%7�Nռ�2�����u�cryU���2����'�T\�o3��9������s"��=\�TWqV繏�t>6���{YE��ZZxw3; ��z�����	=��U�+��mo9^�������=ޟO�����=���������f[�W��`����W
��bb!�d�j�����CJ�,�Ĩs��B��ܘ�E+�ƪ��,�jq��]r���3r�V֎rc�^C��(&1m��Q�����9r��W=i��c1�w#S���ޜ��X:� ����,:��אX��u�Oa��$�E��.W.6a�B$�Ζ�7{��cnV�*LYm��τ�lTI��{/��/�Ʋ-���;v�	��C7�����n��e_!]&���cu�a �v:�V:���OE��G+ �N�b__!{��|YGl�5|%�8�<�y�l��g��x���lHe�J�s]�a���6���|�r���3�4��ؖ7B��_R�&��$UӮ1"�QWR�u��g\O_+�|%�&��vS�K��4/�n��=`�M�T�P���7������7�]V'�.��{�M���V�j<Š.9�W%tgyxX�Q�׏��8K�Z�|�_b9�ݍ���sr�V6wAme��m ���Ԣ����[���b�@�Б.��WyWg%�[H8{[�\��o�:��@�{m�j��e�٠e�H��%�()�^J{��(K�h]��
�zoJ��ʳ�)EN*[H���@�]l�}Vf�V���.��n�R!����S�{��\ìMd8�mVX/�e·粉�#OK�]����b��1��OY;X�ub\�e^��_rHC���H�؉�3�0���H�\O���q��KO)\`m����9w�U��{�o�f�eP�bVb���X�7/��ͩ����|j�
!�4����!}��X�Q�r��l��qˊb=I��tNR�gT��8v��]�ÆL��̬��z���+�g+�ƹ�_D��K��K��Z4=�����#F�T=M�*ݎZ��d|{{��]�8�9�s8;������D�4����̦�ŕ��o^���<`�<ܩ0lU�U3��t�ҫ���cZy5�Ѽ[)��rT:�'t�u�1Il��v,����P�5��00�gl��Jѣ7P	�>�M�S1R岹��h��Z�N7�E*���5��n��5ҷv�b����R	�X)�p9�K�m?+��_�f]��i�po�a���b�j��/`1ힾU@����'|y*�.�ڻ�)�ʋo����ԸxV<`��Ìw�k6�t�L���� >��|[��I�{�+=Vu.
�X��u�[*T�����E�it�h�����F���n��N_f�-���$m0�M�U\�E*���yX�4AD�l.I�=�N�*��a��G�jZ�$�X.��Vw5��m��s5�i`C�*��z��K�j8�yΘ��}Ҏ]�#ml ���#����1u����becm���)7�e#�i��Xs��ꅎz6K.S��upk� G��:�2����������&�¢̈́�O��}�*���:��f�y�1d��[j^��)�"��z�V�dNd�-�G3Y���k��M����Σ�VP� 
���퓦�&
""j��W��UO�tI�S^I�$ֱ34%QAX٢��6]!n�<�UMU�1�j��iib(8�V���(��R�6
�Ѩ�b����M�F�Zq�1SLU\mF�%A^c�w8�LAZ��1Rdִ�")	�
{��J��EUV6JJh*(���(b)������k[�N��ص�(*'AX�-�K�낍��r�[C��t�ZCF ���$�&hh��t>G���MEAT�$��QT�)����7gAW`��4[['m೼�1'ZX���*R�i�j(�"�v1��%��mW�Z6�I֟'�h�O�Gy���iJJ"(�K��"�&��֭�`����Ѫh��:6�MQ^N����E���0��m�Z#^mMA�ĵMl:�֨ʞuf<����<�x^O95}���#2�	WTF��w����Y� �Cq���O�V`�2�<헱��/E����gBɯ��>q���vˎ���~�im��cρ�o42ޘ�G�����;�֘�sFX���vnJ�R���.�����~�Y���q���Z�|��������H�틝��F��������=�a�|��z��%�v�o2��UdC�V�E�/��,���f��mܵ��Qh�o?V�����ZՈ�jٴ9�v�K1���`�t!Z���^���/w�v�2A��5�P�2�a�B�v� �;[�����%��v[yH}�"&�׮��2b��&'��ѣT[�#g�gO\?������v�t6,b��͈��6hj�S�s���o�m�XѢ_�V�#5SE�Ŏ�e���R����<�wgf�v/x�U�^�̜�G�ﷁ*ԝ����ef����h��7U�s��ɷ:�9�[�Xl�ci�Mfu�*�T����Ϩժ�S��N�y�,L�&w�T�Ï@{��)�Хh���Z�s:=�R�l]�uV�Mɏzo&����8�?h��c�[�(�;�˺�">R�{S{�oW�g��Yu�tl���AP��/E`U3����"@���;���ע1�����"�
¶����>C��.R3�)��ۣ�_oJN�Ʉ��G[��.��J���ߒ��]�����ô��P�GK<ʫ�r����Ԇ{lM�!�|�݅�z�<�y�M1��E_=�3����kh�8�u�L�gZ"�@����/9����Jn�n����R�:����k�=r���fp�������I��~�=�Yq|�+Yu��f���8GqדiA�0���N����ٲ=���C��T!��o5E�]����I34�*�ڡ�V��ST�����SG�k��%���z'���]R�1��}2�!z�zV+�Ͻ��j�����6�k��&l��L\�Ơ-<,!d�\/O��i�sЬݜ�Z;��x����]�n2�dն�+L��������e�h�\��U�ȭ�ڧ͇gǖG�E�i���r��T^pꍌYKʰF�e��Z������\��g�{9=�X]��]͘��u��M��/�N`;��SȠ�=ǋ�ղq��e�&���w�����T �JNX�l<��;R��O0v��I���-�\Em�|�����.�n�m�l�ݙ��&�rŔ.l|�����/	��j�:���ټg�M,���F�N�D*��}2� �ʵ���
��a��"��t��>�$oJ����S���#�F�E�8���܋�g̸��`��W�z;�R ���*e(�<{���z܂�S�qtpn�����!�Uԝ��Z�P�@��oAY8J�і�{Ë�!;[&�w&>�U��9��*�j|��}�2�R��*�B�	;�Ë�����UD�q⭗��4>�kr��pq����bSl1��'��v"T����Ļ^͓�d]-�M��;�>l���0k��2�*S���#'%EzJ3�c$1[��y[���J�����ϐ��i����K��w�j���ٞ����f����<x�\��rAG%�h��6q�=�9���V͝���c¦]�3�i�I�ܝ�|�E��=r���x��%���E���D����ӭ{�<s3۩���U�k��-�4�kI������G=��(��7C�l�0�?A���,�&M�ܻ�,��s�JҶG� &���ivIS����oL�8먒!���T�H(�/�����.�`s�D�1�y�ϐ�G[^�GEl:5�[W�\�`	�Z��q��..+�mRc���u}��V�n������n=1ڍ{%v�س�O,qH><C��^�-x���|��nz���o��S�WO���M��K9w@�I?V�A��Aܼq���j�ZbM����a�`I�ї��)8�D��Y�2�ɫ�l'1�����\�8��r�#�\*�m-�_�����7�A� |��W�Ӑ��g�����vr�&���=c����|�����-�p��A$����H��U����&$Y9#��yNj�n;c�����}�-��HE��@���Jj�:Z=3�V�����@�s8����P�q>yv�c���O�w��뷴���c�o���|����uR���!��m�{��۸fk!u�J{��ݠ]U�W��UnҧDm姝ES��Q�|껓�jկ00��'oÊD��&��*���lc1k5�W�g�{�4�?hJ�㊏&�J���m8�7˜֝
g�����>�.�{��#��jǩI0�ڰ�������;�]���N^};�UKY
�"h鑐fe�};�#f�ve��pĖ��G�Kfۄ]Є5��o��+	F��/x�Ҡ�ל�/7��9rp;#�6�7Sh$��Ӽ�5�0�r�ݰO\v�ߵ�L+x�h�h@OC̺c�Vm�Y��n�]eڳy*�*�y;�oy[k�9�歗�h�E��sz��ص��80�3<�F��4Q<�=�KU��+GHz�̹*���n����흙w��+u ��|�އ���?G�����ޓ88����k�e�a�ޝ曁m�23��Z+[�j�z�t� ��ʷ���;�l5/3�]!����+�|��2�+;lF.����g,��}�<�8�ĭ.��vg�ڎ;��K��EoV}{FC�d�aT	�i��['�f<z�v���+]UT�Δգ\�ۻ.C�l��>�f�n7v-\�v�W�yPWjM�{s��r%�q�Ȕ:���ax��]���y�H�QĖ��I-*����W5���zu�}gs���~!1n�=�j]0J��7^�����I��C�����������t`��o��ol�N*ci��NS9���UqxWKt�0w�Ş Ȯ�`�okd|R��X�ߋ=�ݶ���ͿzA�k�Lf���R�)�:D����<��!�o1�ɺ�,-Rt��̲l������s�<=��̔�5�k2[�k�z���5#�zj�*�#�8�����<y����s�d��Mj�c�+w�:Z��B3!�T��7���fi�q�����:Z��z:��\)GgY���[l�Al5Tfe
ٵ/4��Vk�5f��SI�5�أ��#��������/ &�RY������������a�Z�йnp�[���7A*�U�	V��W�e�&�@�|m*򉂶7*��zR[�W+�O͹������~�^�g��n���k�-�6�%��Υ%��m�Y��Dp}~��������~�N�k��Ub�t�}:ݕ���@�3��X]���j��[5gkd�u;�m)x>�3"﷞�����E��[K\�l���j;��1⯵���lY+z=HNw;�7ӝћ4c�F�����4]�����?AA�k���?nϞ��Q*�e�b�w���g�%���򶛣Indi�OM'�N�5�#o��m���M�}P�)H"��g9sJ�s�q�݇▦�٢�h:�ά��㧚9�v���x0#W��lD�捑�òaff���l��
m����#P�*��O�]�cKFl�:�E��r��R� ���Y��o�k�X[�_y����sn�Ya��}�����K�f��n(��Z�2jn|��֙�س5�"ƍK!�e2���:�c�U�_c2��í������3�/"u��[��`*U�4�Fץ�Px�k�!&z�%�[39��y?
�&cw�����LB�(H��w��f�H_Y"��5Z�H�w����\��{R��̝3��C�2D^>�L�g�k/����ŘγTfA��﫸�?L?kz|ϗ��n U,��VNQ5�:����f�i��ɂ����ju��i�y,��kD*���w����Q�-��N)%2�p��\-Ė�o[�[-��\�Y���mn�=.\�L@�[Jwy��w0�=�G+&�-��c����5�:v셴A��Ѵǿ/��K���m����ϧtI��,d�(儍kLu8�:kwp��OX���Z��.�C�\!�"�^����K���wX#U�!��]unL*(N+��_�ְN���[�;�\��5�[ֲ�(���Dc�-K�oPB��ǜ�U�;��2�5�C90�}O�r���w����u)%a<��G"u��l�yo�3�KR�r0�b�����v^h�ɾ��).�R/������\l�Q���Q���a�oV�u`�W'��|�o�u����H��o�+J��_�㔶�ew�i	k�}ɵm#V�S��T����:��`,=��u��i3�+sM�"�f���U�����a�F���^\ELp���}�����+��G!gG){[�d�vr�<��D�]C�ZD%��fvG~����;o0�A®�W�-�������_714v�`�=nM�\�v�U�4d�<0�	;��y{��Rw�c�]i^؞$Ŀe'����N����=����nլ�I˴\Sʫ��\��s�}kpe�ٌ��J!J-b
��]M�gF82L�,d󦲞4����鉮��ؼS�������yN?��i�T]]�/0��h�?/'^o3-����m�k´L}���_{VSq^�]��0qp��<o(�v�����pe�jQ�\�
C�,8�i��*�={��A�X�4�8� ��O#�{U��>��}�����vEY5G����<.��ןQ�3~�#4�jc�j'm%�τ)ymD�c9��=�9��e���^�T�<xt�ǚ�r�x�R��q�*�y�����e��8GFPz�<Q&��]V�
�*o�1���K]�,�AM� h�9ݶ�]d�i��7>q�wm�Dvs���(�x��J�=G���x�Wr�nG���'5�fi����/��]e5H�c֭���/�7��狀|�o��.G��}���ںȔ_��p��:���E��0������`���[�<�/3��q��>ġU���	�Jv�3����rcV�d���W~���k>gj��OX����� �fp/8[�!����l�z�S�[	�k��XV�o�7c��� �ŗ��Za������g��{��b��<�Ln_1�;<�>����H�H�-�'yd|�4p,G��n`0��i{P���c�H3��Kqh�mlt�+�^-�i�w�3� ۔��+��8	[��[��{\��αY����8��6{����>�������%(Y������HwlQ��r�)�K�5�� �Oh����9��p�0>� r2.r��'A;m q��30z�t�-���Zl3�x�櫚���j��\u-Mgd��{֐O`�	V^�G>ɪ֍X�2��.ˉ,̂�~���vΝ���A��Vؾ�Ǳ�ź��S�~�GL�g�Ȗ�#�s|$0:�y�
�m��6�=�j�EJ�Ŗ0��Fԕ��qo���oh���+���Y�q�Y�J����ag��v��O�"ou���9�r�DA�3]�cA(�qY[�X-S�l�{�w�Q("�Ce]��
�6k�o:��®0��,�AvZ��*��,Wcq��&��;;]Wr��z��p�ͩ�����Z.@����F�q��K��U#y�(<�pY�GoEv��N��,�{1vV��S�mg9�5.�����.�UeK.��oc�Ϡ��_��ʷ���D�t}�_��^��`ns�o$`��y{||}��O����}�m}�~�|>]�|�&�]�$.ɓ���
{�2��%��Sy�l*Λ���lt�z�ۅ�d%=�𹚨��,D�iΝXrq��b-vqN� #p�6���r+/�b�,�嫸�+ ޽X�(�*�"�ӻ�u�>��+o��6�0�"�fҵ��wb����8v��oS�m @����Mc��m�̧4b�ѵ��άјd�-���,R�������keɵk �⣽LM,��p7w��X����g>�.囩���V��.�����u�޸�m�����e���\���c�u�or�:�N�6�����t�)ΧR���ҷ6��
b#ژk��ejq��eټ�,#a�ж+��r�]�9�I�k��1Ӕ~uֺ��/]]`{܁��1T%,e9cjk��d�mљ4F2�^�+U聲o�ʀ�zc����L�����\��l��:c��t�^\�#��OT�OLn����֭�ed���/&�%>r��[���s9�|��ج�@����v�)�)���´T��{�M�R?x�(�iՠ�{ԅX\�g�ړ���w1%,�����IZ�N�[��ܴ4.0�Nޞ���$.z�u޷�'T�⯍�8��\���c���N&�٠3��hK-ُJ)�t�(��<n#<N�}X�3�ITPX0�͙���ζ(d�!O�SZ�v;��W�Gz!��I���d8�x)^Q<gʗ%Ի,+���P=��S��S)\�l\���Z�=4m�8�2r\����g+���+379�,R:5t�Wda���W�T�d��{��7g�|��1<y�"����D����k�ҧ�.;B����}�<f�x���.�1�F��#���%�4tG2Au�u˳(qdr�)��䝡�@��K%=6�:�ĭ�Fm7G��"�(�߈9ҩ>643�n~�hUT��S��C��,df�(�!P������Xyjl�λ��l�i�}��kT�7X]嬑[ɡ^MN`��'7iN�e*ʓ��5�;*F��Ż[x����d|�䃱*�T���'+'�'�4RV�v!cC�G�v7VTZ%l�
�׸�)O �9�N�u �%�r��avv2$p���1Ѳkt��[z��d�'p'yZ��Q��fO�Ԍ�D�2��2�%݅s��B��v^��ӔFT|+����*���gQ΀�k6�YKa����еoc���ԗ��+�S�qd�p-����zL;�?��	��{��U���s�m�m��ڌv�֙r��Od��+`��[
h�\�����E�̖%�uhį��ꊘ�*�WM���[�$��2��㳙�Cs��]�[�{R�	�ƥL��|����Vp,�хZ�6�;�o=�b�Y0���mhq^����z
W�G#@c�Y�xYR�������'/�c�Ш���F�;��$#����EU%,EUD�SZ4A^F֊%(�������iS�a)�;w����mI�@VKHS2�Zeհ須�M��J"���T֍!IDy�y�:���ѣMQ�qP�ҔWF���(�ي"cFZN�UIM1U5H�q9��!AQ�Hi��<��;j|���A]�v�Q>A�����#TUU�B�<�� �'IT�yq��� /2�GLS���D�Eh�E�-i���U!KLOiݸ��d�4��B�)������8�����y���tQ��4U-w���G�鉻:Kn�n�t�c�����2��dE��0�}�|�b��j�ra�(֊���Av�*�r}W��(L�N�sz�1�)9�e%]�����*cX���&*�+�,��\�z�@&Q��E��)$)�e�i�`!�mD�P
��;����?wl��uyIc>w���g�k�o�9lV-�"�i�U�#���j����.R�~ːJΣ��vYa�C��">m�.�b����w����DV��vd
��=iA�Wr��+ik�M�>}���������蒖ӭ_���0"���^�&���za�����yj�:�m�=٧n�לʽ]t6k@e�Du��ʏli�nY{�z���lAyi�h̆��!�1�ފF^&�P^�-ۻ�F# @Xd^aŹ�36�Yl�9�;v��}�����g���a��ey�8u]"9Y^l��z&߆�F��fӥ���tQ�v�^�[�$�
�.Yc��{�x�$�OV�����ȣk�7f3x�\	�VAV��]p���~�ϥTԮ�W�x�tݗ����"�\Ф��~���8F�Op1S)ck���_���ֲ����.���efE���k��n"z�Q�m�o9Q� wt� �z�)���n�Vu.dGx�֮�{�HH�2��z�29�ۂo7gh��T�Fz�B.�w���8, ����E��lu&��<?��í��{�K5rˀ׳/J�7�\��W>״
�`����M����ə�����f�h�
z#M�����vT�i��U��u� 4pv��:�tSU�M���4}�VR9�NV<��u>	8���b��K8��g^&o_/�Ь�X�t;/��}�'����im�̃;8ٌS]�-�fzm��W��i���#�]��$�<�K#Һ�Xʽ�o,�"�ؿjG���cM�f�G�\dz�3G�x�B���(�=��#lq��==���KL�g���`�0pp��"��A� \tW#U|KɺF��%�L�ύ�S��8���w�"ZwY�����7�:FD��a�ȭ���˦v鷴)��)�ʻ���Y؛��|>�2;Z�{��큛C�]>��k%@��bzy�5L�i����6���#l�%e�l�3��ߧ��f�sH��Ϋ�{�ۚj��ޫao�m�b���z�{-m�qFh�m�[��&3��_Ug��x���=�Py;t�lջW�1�����l�
��TCGx�"�]��n�R(���X��EL�x�'ucY�S:F�W{��o��M�g�9���C֚;)ݵz��7R����C	^Mū�n��g��I�z�����v��1$��=����I�(S�prqF3܃w(=�3w�0Ь��S���햠l?)3ήx(m&�(Y$4�;�s�9�۽Z��4���9{�����]�[�9)
��
�]��1fԚ퓮e5���?'��W����[�<�	y�ƽ�Ƀ�77�5������fV3@���֥�@b�C٭�OTTOHĻd�˯�w)#�s�ђ3��,��7��p�Jq�Kl��ߥ�B)��5R���y��Z��̜כgڊ�$��$���e7��Z�6�Mַu��n��|)Kk���HJ��=Ў��8�gzn�*ؚ��sr�&�д�����k����vυ�[����cꅘJ�)Ё�^��T6\i�R�l��N��u�ӑu0�<�nס�i�˴f�U�M"�<�#�z����uLUiv���	�K����V���f���.��8:`�+��p����=���[�i��9��9�V�e�V���ù �0�]�5Iy����e�ج](F^��Y/����)�l&�ٷeǻWHʌ�Xh�R�gwV����]}��e�U���5:5��]������]�B�;�Bhl��9�:)�%�J�]Ҷ�N�Xl�����r�����9S5��g�[���ss;(;ˊ�#����㺲�0���H�ly���'8���z���>�0�y��YIs�z��j;>������/h�CM�{ܪ�s:e؆�S�
ԋ�$}�o��cQ��3+��l7��\<�O��t[*��Y�ha�1�6k��\�r�dolx[�a�촃ZF��,�\g�[�1V(V�gC�q�<v��:�n;�Zgј�\����2}�[��fS�l7d]uWj�� qk�޴�m�gOy�C��L$�D٪��9��&f�V����m� �ݠQ>E��V�u#e��x��^�_f��V�6��{{��#L�2��U��Gv���T�-m�MM9�V�<�Z�n_傸/�'{g�99;��
�Џɻy�۩`n�o���H�.���M��m�۫�Ÿ �#�Ӹ��W���!(Gv�u�����ڲP��$4��:A�_}�o���&�����x�p�06��'�
g3�7s�v^�J'��
U�D:uY�mWo ����5�Hm���7��������_^{�I����U� ,�u�4�t��&]��m��(��
���\����v#��K��u,�%�F6��N���Lc4{�1� f<��tNo�K5�[���֌����%<sqU�X��q��I�-C��l\dUz�dg<�Kʸ�O)|]s��C��UםQ#U�j���,{z��bK��Y�PRX�n���,�m��u64[�t!R�1J���8�5���<]�\�'�5��%g����LC�w��Q���=q/��i�]Bc`V�֮}eA+�Y�m-s��C��t7A�/;,�m�8�]X-��c���fv }Ϊ�rXk�M��w>�6=[��tmFo5�h٦��v��I�1F|#��e)�gΩ��N4sW9�e*�u��5/;�� ��$�ߕ�������2���}a�;k�m��O£va0����L퓍y蹉G�r}�^J�v{�d��l�v��SE�20^�� ��u��RܺG�f]�}�~X�[Gۺ��m�:��WlJ؍�M��؅�-���Tiй����甹Wr[f=���s)lg��s�y0$�6{o�g ^��� ��zdl6t��8|򾨔W1��[Y���h|�L��ޞ�aE��M��!�2���!��jM��RZ������|F%�1��h(��̲J�h�N���^[LUp66/�2t�R|تDr/*U�i�=݄)���J:F*hUKb�C��i��5���-�!�a�zUu:Z=R�*�@��{U�����������Ȩ����T/m��<.��n��Q�}ko�lL���@�0J4T_���7ދ��g�]�{�ʠV=[-�:i�ম����g�4m잦;��ѩ�2���=�VQ���9� �Զc�0Y���Q�]�\�̊��6�D?^h���<ܒV^V��]y�I�wvF�+bVq�ˎ�~���3zCۄ>�Ϡ�V������^�L��"����(����7Dd
�V�]V��̣�OL#�` �;�*&��/;�٧�[
�#pe,�:G_�\���"��B�M��f��%��H.��Xgp����x���W;}vH8�l�G�Yk��1�&Z�[9�jY���MG�u$0Ĵ_P@�x~�.�{�a�5��m�!L^��7�U�%��d��r�e��I��o�����?.��5�m͟B�wH��p+oM�"�Wj�᦯�v��'ul���d�飪�}'Z�d�7F�k�+�;�����:��u;l�v�F�^s�i���ʳͳ�3��ߧ��1����xbf"�ރ�Ϸڛ{}�Br�����$�o3��߾�/ ��=tӽ�k�h�zo���mO���FU�f73:T�z�m�і��x�u�63P�b9i��n��0�1��"5Q&zL[\���jDM���I�r:�)�Z�C��Q�UgE抝�؛�F�{�/9���,���U��M��O=�X�Ԅ��/Π��6��w܀�^�h�s��c��j���񚭦�Z��Z�]p����IM��St0ڪ��g��ؗ��[������B��7����Q׺����l��GpuO��z�Ӛʮ<��Hۙ��r':}���nK��)Tz���V[H\���8)}w\M���3�ӛ̜��>��;{��]�������i�Ɇ�n��JXV���=W|�\y�	'�oOe���=��Cu$ml��Y�U�i�e٬���V��U�CV��3��ꈣ�<�}z6�VtA��Gx��qVM+����H]\�������_�����l]Ԫ�]jl}����D�ѥ"������+�忔DfWF8�{Qc/q��5D��0�<��x#>�o(��4�@�ED?+�����W�����}�����a�mP���6�O����սn{�ɨ��l�)7{���S�B��%�@�%,~�*Q7UO-R2"��j��4���f>v���Be(�J앓�x�>�ݏ~y��L;�s`@�ë����5�U��{�6ѽ�b0�FG�0��X����B,��WO��(	'�[�{SlݽX^O�q�ͥL�"�z�W�/_ur�N�A��nHR�u���c����
xjm�q��\o�z�l��غ��1�u�88�=����; �Xtw��V��0
�l���Y�_��S:�:-�K���4�O��x �yy�̿��36���N�"�*�|ʽ��!]9[R�6����KC�[��U�_�--�xk�Y����j8)���j]u[��csi���BZ�R��U�+��*��kο�HCge��!�K*�u^daQR��}3���jz1�{^����q�ܩ�{��=�Wt�B*bl�A=1�c���}��k��f!��E�*IHl�Z�b�h�N�e���@�G�a����8�ض���O�X,��������[�GNhi� R�Z��ʞ��i��\mC��ꗔ�������V�w�_o �R��4�J��c��)�C2���'a���;v����2�`z��ϊQ�x`^��Ж�JJ��N֍=�v�T��2�I�U�$^2�C�0�g���䌍��v���s�v�No\eL�5uǙ��qq����J����e��g����ɭX^����7���.��F"#���wf׵�Պ�=���8�c���5��P_"����I~7G:Ê"w�f�q��'~Xc��m��+:��������ݑ�� �[UN��1��_�W�:�I��|���kbf�1��x��70�V8�}}�0#��R�<�&]�f��Z�V�eq�Ym��
ÿ��I,c7���m���1���>���		��9~�9�:u��H�ɑP�#ն�2�t�K��Բ��n;汽lC�K~L�J�Q���oW�6+T�>�zS�+ue�V��km�wY�v��FP19��&�l�{9EH��Qa�z��Ж_��@���]�]�U�Ƣ�i�"��^y�-3��r��7_Nw?b��膮S73�P.{����r���gg�l9�{��[�]���g��v��n��/�d���ˮ�q�m��gY{��_���j�A��a��d ��]GXL68�잋���\C��[������gs���`��O�e#a�H��BU�9�0*�oh`�ƚ4��^P��y�7x��FO�2�[4T�4�u�?�ʋ���f]=C=�_���'z���-S��B�H����(LVf+���IY�-X��ߠ7���E����M<JԳq�P��r��9:;�f�)�����u�mq�T���G��L��-ox��X��|}~^�O�����y�����1���W�Qg�89�hQs⯞M.O�(���uͷp��L���^ZD�C��g2�(��\�8h*�7z�
`�J���Q�,�y��n�9���E��=\9O�n�v�����רc�ab�u���z����ǽ]v�/n�����0��3_��0Uv���t6�w�E��.Ev�5]lK�p��$��P�DFŚ�T��oFP�ήJ�u-�;w��pc��2�2�)�B/7�᭫ݬ^�t��EF(#�7���$\�%�^	�>��yUe1�m<5�o4��nV: ���@S��oR���|�p�s��|��r�CB���u0�wk��/��e,��(Q�qh�VhG�ifb��ec�Z������yP|^mL{t5:[��w��CyWQyu�Q�����ړ�,��3�Vq�T�|V�uu�7Z��F=y���B�Ӳ�k�e1��]Yn�)V.g^��]��l��v���!�4�oZ#�9�H;��H��I�j��� �37��ȸ��05�1���腲ΠgN�O/':B�����N�<tp���Q�Q���,G��z7��㷐;dlA�#�}P^%��T2�xQ�8b�-,��bq�w(j��m#T�S�ro)��h�Oq?�F􋋫Wuæ�f�|�n�D��jm�zr�p0���F<�KA���R�GS���'��)Dp�
Y�]�A;9}�mQ|\��V�=-��e,��]9�vow]Ww��jf����s��`�I�ɦ��ŋ�b�ɍ+o,��NKUGS�z%!Lo��V��4.�W��s�)�ᢅ�h�lD%�7��vLj�]��CI���P�rAƱ�ߑt�6P�%�˺
cc�;w
���gJU�qR�x��ru	�iP�.��E���ΰ6j6��wY[,6kV-G_h���.*௩���ū�&��l2]!�ќ{U��V�+�&��Ʉk��%:�.�U������S�U޳W���YP�ըų�9Y�����\5Z4T�8�7��o�
�����pBT8�X$ں��>� 	k	�̾�n͞{s��|:���->}* 6_\˨1��oj��#n�<	�� �ٻa+V�
Qk�U�z�B�0�
S���nǛ֘w
��T�|�f��y����z�X\�}��jbIL�s��pU���z@�"s"(� Фd��9���$��F<}�Y+\Rቑ{6�mFc��G1'��6�a|��V��^�F-�V$�_A���r����p�!����QM��Y���B'n�ۭ��Ek��'|� &�pL��
�h8�:#�*eϛ���?�cM����ES�/Y�X�c��6Yo(�%ku�*���J���1�_n���R��P��$̬�P��s�[ŏI��).�G
*����k��<X,��݈���W2��9+5euN����{ysRA>���%��B�p<q�b@򂭠f(e��\[�N[4�,Jn����-�뾍��@kM%:�7con�:J�z�m݀��!��{���bJ)4h��AAA�ݬwu��w!I��+Z���w`�Tm��TI��b�5�����q����y/�@�ǘ�ly�t�bǘ{w����V��Oh��x� �(̍�ϗEmE��Ӡ��q��v@�]%�v�w���y�I�������;�͆�+v.�H�h�͈��1��qb�w�n �$�ۤݍwGpk��)��Gc<]h�'��mōݮ�h)z��ZcG��9�*��>^c=%��m�4�tu�i�m��tͶ�N�$=�룻=!� �qk:i��h��Fϑ���ڨ�����Ӧ���VۧX�KA1U��OI��6���xc�<��V�=qt:4P�ݷc�,�y'G����̛v:&�j����[_��~�ُ��뽰��Hu:l�{��"��F�aCt��ʱ�p�6��Ā��0/��
�0�5���鉝ΝƲ]:9���<��j$o��IL��s���Ӓ
����U��_M5����\��`�h�l�F�aǻD&$�]u��F��8�>;�>l͏X�\����F��;�����Gf�?��Fj\9$�y;������,]1Ra��ٞ����}E�j�������Z:ˊ'�%ko�_μr��?����1����.��3�a�u� 񛍁Z�U�/ �-��$��:!}56E����T.w'SSd�3xX��4	���Q������wp�D;D�Tm�NFr�
/�Gv�{N�6��o6{E1]1ڍ�.n&��[y��Fj��\�K�q�3	uJ�������O���*ܲ=��^/?�wV<�k�-�8��굽^�Ѧ	��[{	�f����G3#��K��V��_KѪ&�iܢ�Тgp����/\�	���<��ct�k�����+ػ�w����q
�q52��y�V
.^hޡ�<U�NF�k��+���=\M�ALл��Z�v�j��v|��_:q�\�K�m�3]��j��B���.=˩��y�/9^����G������1���m�q��뿦�a��뵧�A�"&�P|���Ż�D,u��S�f�����n8�sq���y����-�7�:�O	����⛞(!Oegߍ��+��$��H�M��W�mw�����c�Ǚ�@���rvn��Z�辬���)�f;���Rz�r��4�B�g�t��UCr�+����C�������m�|E�����Ԓ�Iڳ�)]�ȷY����0���1�����K�Z2o��5�2k���X��UX������Ӷ�6e��2�t3Sd�[dX���|��#;����yׯ�_��3f���9�7F���Y�]Ս��w�qY1�t�pl�@���)���r����e��k	y��=�	�0��-�����ս�d����6��Yۭ�+�s�y߉��J6�V�샬��8���y����ʅn�Ry�_�����ooV�lQ3���k���I	����4k�Į5�D�ʓlV�fS������=�{���I(β�9�&�����a:sLZ�Vᾠ�e�DgP|�.c�|�1��fc�A��;9X���$�2����1�0[� �Jx&j�>4h
��l��W�ʫ�N���+^^L`-im���Xx��y��~���[ǻ�����MVdD-�͙ݼ�b	�B,��Wb���כ.z*��~�@��i}{v�#U�6�}r�l,�������Ǳ��`n:�'h.����e�oat�[����\+�����h��ޞU�	�
7v�(>B�bV�%�>�}/���,/e`.z��Ÿ>�=����
��L��n�~����I���)�Cl3�5wH�V-YR�f�z�b����dQ[�/3E7��E�*f�.�l��� �h�1�[�)��f�t�Π�L�ZBy%�U�P�m�;���ڛd;M���_���0{I����� �]�g׽+lr
%F��[}m�Y%�C�!�o�e�k��ȡ�>���ʮ|���-L�� ��#b8���d��췃Zá�TuЉ�o�m^���Ԕ{kf�j�g>�$��H54���#���rw{��6�����P���m�]Up:�,['�ngvLo1���Wj�y$Y���ku��^ˎ�'�ɡ��N����Q᭫u��ț��R�{7/��I�!+�ƕ/�Z���mgz�=�Ԯ�l���d��,c1XF�u�[>�y�ٝ��2ϿqE~������X����{�ѯu+�:<��ğ_��$��Nm��d��AIc-ա��2-��*"h3�����q�(���0�
�)�?e�%gQ�a�,���U���mN��{���U�mV7o;b �W�6+TϫW<�����]�-�j9��de^�-��>����ɉ���e���jT&v<���|��%	]����'���Dc[�`��~���o#�鋈ۖ���!�;�?:~�\��*�9�ĳi��Gd�Lm��U����S��6dh�6O�OH���,9�S����A�l��gn�ڍ���N bL�����.̛�I�p�&z�a���|����{ϯ>���}m��{(il�O`�+�g^�r᠜3�7f56Б8S-�	�[nq#hP�n��B�<�r4��}E��=�7��.�p
��%0��}�3�I]w�t>������Z�e�sL�m�Yx{
N�EuJ9��u"�M��8�/6��tɸ5�O�/&����Y��p��Wt�a��v=OH��y�,V��u�JV����Z��{���Rm�zjL��ѩ�:	ӀD�}�����|���]5&'��juEY��O��ۿw��?oYUЯ�u�g*�����o@~ԱCS�n=�G�����5`�z2�%��_*w�o&�6d2�]�}��,�:j�!!���7/tE�z��ǫ�$�YU�]����eo�Y�a��z�,�rN������^�(�Q4{���F��v��m
�䚞&�����a_קϼ�aپ|+4��D'����׃)�N\m���2,d��<Ֆ�^ކA�0B��i�\;�q�]V���cT8���(F�2��̗M�ȱ���}���kR��%�q���J�R7����cqy�J��ycSd����XvY����9FD׻����Ł��ٌ2Cu����oA�K�^��9+���z��{�ҭW�N >�e�kݖ5�ߗ�:�J���{޲��V�-�r/�
�z�كC�Z>�|<[�'>�هu�]c��M����Q1g'p*@q��%�GZ�v�:��:��T@�1�>>�!�@JVbw �L+�W�2*"�w���s4�n�+�Z�d��y�8m��sv�n���p��$���7�K�ݫ,�YV���m�6�=�1��]�o��YW^N{c�d�b���`�[�}]�����-��Ӧ$�!�S<Y~z�Mq��+q6%�ajO�lP���F�a%�i����.H�s����qN�}��eQk��C��
̈��^��Wf7x�:�֦����]�����`7EL@���"��̍M�CƋ4Ҙ�깣Ǯ��ɷ����9ע���9g1�o<���l���k,o�����CS&qo*'�f���,rR��~�!A�/�s���e��6w��ߩl�8Ш�u��s�ܦ0Ұ���'/J]Ad�j�Wtr�D^U��v}i�����uo���u5��Y"l�d?�V���볊=�ث0{M���qWm�qoF~�!P�h�GoZ"�S>	�	�ԙ�u�́\�ڃ�{��z��5vb�V�r�7=��	��ᗔ�å{i�Qf�c7����݄�벙�1K��Q�`�CMIU�0�0�6�3[��P�8�R�n_����-Ckx�noX�$��5 ����U���m��'�%ub�Sq\X�%�5���������n��j��E�Fn�z*��ڎ����m����F����Ʈ�R��X	������u��b���;��޼���X�'Z���cm�ؽVI��w��Q]��r�8`A�2�eO|cbv��LL��|��J�׸MߊOUo�4�Z���ڒ^)��æ,U�O���ra�.#T��ә�ƕ���E'i]��R�类$Ledj޾�U���>�$�ؓ��˕�	�۶��rٔIk�t�M��.}o3i�G<��Q�ܐ���N�F�8E���fE�~o^�����㍼��\�</8�;
{p�
��i'�qUz�����X^ʱqMo&o��gb�Ʀ�rx�����&����gK<\3�������qm�u�+!��)���:�?�?w��|���:��&�펯�O�\{�fI{v�V&eS�e5�^�X�^y�j�T�׾ĘR��@4進o5s�bY�k�Y]���4K��E�;#=t�/����E�I��v�wx^*D�@�r����d4��.8� �Jܹ��(v��������
�w7�{���"�qSC��ө�l*>�Ù�Χ>i�V��ߺzj�t�}:�D����
��%vג���lXg�n�5�Z�ڼ�.��ܶ*{{\�\��Jk�~�
��q^�e|�����m)z���Գ���f���U����h�����R��]��N�G��.���lɝ�>&{���V��Ȑ/T�`�]�y-��/y�\E�M��|"�i���Ǘ�ԥvT{�U�]�z�w�X*�^���x�|F�XT�����P��F��;�&�Ǝ�v�]�*�y��"Dp��k\�	�gd{�	:8sj�!κ6�q7^�(y%r����ʂU�r��.ƾc+޷f^j��^���!oP�Z��*9�i`������W��{������K$����!��F�Bgcϻ�C�,C˛1�,ǿQ�X(JX��;�~�m���}�zֆԩB'$K)H3�"���/4e�'>�i�A��zD�b��ή7�8���*q�����$�ۼ��U�J�	W�d����ojq�e��G6���ti��j��iv��'[�w�͜�q�=�*�^ωMR��Mm�Ͱ��y��3��3�ʀ��pf��޼m�;�^7�.^s�ul�GX�3; q��{��-3{��b,�r5.Ƥ����U�Qޝ�m߳~��'��9��Η�є�x��u�M���6v��l�K�a�}�ޡ�[�����
����w'��Θ#�3M+K�w�[R9=F�<W��y���ADY�V�G$3�(�Ʋ����������V�E��������(<,u�|�j6�Fe���M�����Țg����b�^�n�M�t�e<-�5��9�|˝�ĎT��0j/@���U�ڷ}L� k�cP�6.�Z���4���t�����΁�fz�-�sƅ�Y@��`���ǁV����{�\T����]�wO�f.������_� 1���D�ɨ��YA��{G��t��i0�6u���=5S��#��m����:c���gj��8��L[ ��a�d��س5aK6�f���E�t$L��z��̓6e�<pm����o-|�:cw�<�#+���蕝��3����[k2�;��P��
5����ꆭF�;����������r�� l_	�CrI_��ݴ�s[�NfMsE���ۄ6��F����c>C�� �6��[<�;|�t-<#'����a��ɓ����E� ɷS����ݣՔ�tC��B�g�ժ�G���f��g1=�Җ�L������,jl����a��6aoH�(�W�V�Wt1y�`��s��ΓT\�[�s��u��|���s�ݞ�<,�\Ȝ|.WX|�m��,��ha]1��Y~�ym�-��vy[�{I8�c�0�kk�Uά�5�@n0���I&�{�����M"u���V��C�LŬF��n���=�2��ᜅ쮁(�]�Fw���šȉ����a��6N�ɸ=ޗ1}��z�;�_���r�P1�]�#��j�&a����ʛ�	{���jƄ�1���ȡ�\b*�����������R?�� ������s����  � "*;��8��x=�����U�E�U��U�U�U� &@$!Y�fU�ae!�!�T!��X�0�2��� � ��������� � �>B"� !� 69P� a�T ì��{� 0�{��U � C(�C �C C( C C C C( @ʧ���P@DDD @� � �  �Q �UV�U\2 2��ʪ�ª�( C*����0 2���,0���"��*�
�"̋2�0,�����0,������ ����x1�~?֪��
(L�+0_�oO��_o��~��������g������������o�oG��ڝ���>~����@_���o�O�E��@X��7���؁�?�?t�������� ��������������������>�O��~�� ��  �� �  B B H����  ��
 BH ȀH  R�  A*�2 ��� ª�H?�$Ar�����,��!*�#*� @ 0�������@��@Ň�_��$�aE��hUQ��W��W�_�������}�@^݃����g���'�x������v?��'��~� ��~("~�O~I�"�
�� U��~,?�� ��~c��
�
��@g������!�<���{'�x��O��x� ��!�߫���W���=�g�������y����������� �����P@_���~^�x���~i���>�?/�~���I��|~�dW�=�f~>�2� �p���~���QW�0}�oD]��O�����2��b��L��En�@�3� � ���fO� Ą3��h�5��Fڨ@$D�J�l�TT%)��R�TBQE"U$���ҢV����(�!QU �P�(HQ%�T��,�k){�ګV�M*meH�kN�"�l��ai�Km�
6�R���f�M�4"���)�F��mV�*�eM�77.��ml�ff�Օ3YgwO{��1��HLʒhf�bԭ+mkT�M��ٵ��+Y*�U�[4٣cM���SmS5L�[V��+�M%M[bm�R�Lͱ���B$U���*��  -����g\��	fuv�t�Um4a��*�!�Ӡ4�LjZlh��m�R�v�a�㦃6hm���+b�7i��73l�݋F՛mZ���UVi�Zm���  �(P��>��B��|pB��� P���(P��t ��P�C
(Vʀ��T�V��K�l��6>���҃��Á�@ C�E�-+�v��+kV�ki�6EY�  �x�Z��v��-����<�jvV�F��ͯv;`X��M���:�1�&�;n��[۝OOTz�M9�
�4Y���f���5, ��^��)J�Q^���*�%���  n�M >����8fZ��[ms���M�C�N�t)I�9݆�R���s�AB�v*��¡ �n���Z�ŤP�:��L2���3IjڱT�̐>  s��րL� 0[:�45Ep�}��U�"*M��Q]jP�E�� eJ���tK�ۛ5U�7k5�.*��KZ-�V��|  x�p�j:w�6�e��U���m��݇m�TA��(%��9��C�2�t�N( w]��U��Ѷ��wl�b��PD�� 5�PQ�Z�}h�3��UQK�5��j��*�N�4���.D���ҢR�G��]��hV��(P%�wJz�[n���F$֦ɬԛ�  ��蠒����5���4�{�	S�zn���b��U绠R)Y�.�R���'u���5���ys� nz��= g�JIJ��j�j-�kbɶ��_   v��%J�t�碥����˝(�x].�QJS�pT+=��T�TWw���RAn�R�E�9�D��ָ���
��z����mTc5���Y��m�  ]>�����E�<���p�E$��{\�2�P]�U[���=(�(w5���I���ꔥig�� x�J���x ��1���R�  E=�	))S@�T�SѕT�)�0O��* �TހeUSM�ɐ�M$D�U"  b~���~��_���g��{����/��uy�2���^>z���X��y}���}��|$��r���IO	!	$$?�	 BI��$�	'�!$I$!$�����?1��E�~g�y;�� 0a�}�Zy���[Mf��dI�-�p8�Kv��C��Lc�������w�*�̨Q�^��I�.�|�C9Gɕ����	�5��-<7qfnf�cE]ʓRR��p�_Af�5� �4�fc�skl�-�Ua�u+6m��`��rk��e�F2kL/"b�ce[���i�*ZZ�j�l�� d[gS��s.

�l��f�5Q=��q�1����r�M����69�Z�&@�����ELTpSb�
��9�~�re���ƍң�7F�kyf���H�]�<�E���)KYr�i�5-g#fC��E����,����o׍-����v(���e(�0="��"��;���.�Q·-�y�~i�&2ދt2��q��*��ҵP�9��.���4��nm�C*���<�
�м�k0:�ct�z�J+�A\�1n�%�欆��5f�dS9y������`�e�z�X:�i�`W�n�UДq�XQ8Ad��n�K_2���nۀZ:Vŀvj�t2Ki�m[0��T�p\�������VŹ�7i��]��L;KV�V�T.��uyw2��h9��IL�D�w	rQj9ejU�^+b&iz�X���Pq���Y�9h340,b�@oa���;=���-j�34�Yi��Ұa�*ƽyQ^ӵ[kN��y�B�ƽ�J;����Ucv��Ӥɂ�*զ3M������*�2&�����P�C��7s}��x����ӥc��u�sYL��y�Iފ{�E�J�O�V� ���ԅ������K(�wVf<�4�e#,D�����$��b@��4�V�ْ�KF�Zj�QC^��(B.=�s%(o~�dv�^�" *�K�BB�4=�ӫ6a�,�[Qn�YLoKLK�wEGJ��s7Q���U�n�ی<{@�W�'C*G�m]޴]lϬ���Ri$�ߎ$��óq��T���㷖4ތj����O/mą�m	�L�/-aP��;�-���m5�5�-�)*�wd���5X-on��BW	{�sZ��S�Ff���FA�@�Z�e�JL
�v���c]����rA��&�y$�	�/aڃsj��/��nkإcw����u������Jr"��a&Θ�� N$oqY�.�ূ�����ͨ�Ƴt�P)���T��p���I�u-)���[V
�+m�{�ۆ��K4]�UU�Tl��+@�q��l���R�^�j�|hLZ��QI�Z��A7x��՛NLZ2e��(X+y��JFi�l�zn�wJ��Uj!�����j��5a��nYV����f�E�!?��Aֳ��oS�f坄=Z�$22��!i�5�o��5�ɔ�ծy�ݠ��F̆Y&bۍ�z#h�R��e^�ф�u�Z�V��6�Y�Z�FVԫs]�2��Ot0�*�M�&�7��j��Z��(f�n�e\�˥)�8�iKm���*y�Z���ڤ��jd�iff\��Zr؊�� �Y�w,�b�QoL刯i�LM��.�H��Ø��$����Mq�3�B�-�^kfYSi�#��:�k�b�HN��U��NL�5�ݻ�����`�VK�>U�RJ
�h�ɺwXB9����5.*NYm�����o\�x��xk��0k�B���g2�t����9-��eH�U�eB+M�y�)�bj%����r���2H�a%��m ��U�V�)�#�>�Tf�@k�\�#[�z����t�\��w��f�Mc�q�Qj"*��ӌ�����j�`W���)f,v����GwS�Z�:��Yw��@�'5zbK5.�|2���wf�[�gD�/K3%�p�o%���5\DLźl���"���;B�
��Tvţ&jȀ�7�Gbn����/A6�sj]���&�ǈ�JV�F�eJ$P+��Y�C%��5�n��n�@HH:C^m"�X�͠�Z72�R������u��CQ*V�H{���P&�i$3v/XYZt[�hQ�!�YF��Bݽ�ݚ�v>1:���۔�p3	y�8�Pj���2�m�EGa�q�Xc�"�v�"��Je���lC	��]Y��P����V3b%����h�C
2*xn�jJ
�Gu}�ƗG)�ѷ2�����KB��V"�&.��w5�N�W�*V�l����Ge(6J��z^�Ȁ��,�\��Auk�[,�8���\�2�N���sk����ћ�2V�D	ҥg���t��q�5ɜ�]ga�[��w&Z*�,����Ck�&�����eCp�y�Vjˣ�#b�n�����5�I�p�%l�]�G��Isop}%dR��Hj�x��Eh�1;�m�n�Y3c)�f�'T�;����"�X��ayZ4l	�Sy��i����,�io�]���p�9��;�*4qG��Il�4s(j��5;c����HD���[�X�ҫ�X17���)`��앺`����k�.��9H<0��T.�'!P'0�L�V�[�0���Fܡ6�R�[B�!�Vb��GVS.�nV,:&�7�(1�i�V*7���é�<F��!*d2dO1�4����i��?dH����s���6mVVt2T �uh�饭��V�^.�;�!jt3g�Ԭ���E�{Y]sC9�uͦ��SZ���b
�w%��1[]�E��^�+�	��;�*]=n������i���zj-��:u��˅�3t��Z��1�8�V��۵7l��NZ�M�]0i kb͵�n�xݻ�I�� ��T%D=%���t�]f���@MeUhͥ�5��+64#p���,j�u���,ۤ�謕�%X��FiLk�xo,<<�\�ih����1P�Ȼ͢�T��d\���7o
�H��[m����i��D�'�`�r��n�����i���AȨ��,��3߶�5��bN�������H%\9&-$���v�k��m	ň-9�5u��� P��R��)Mi�Μ��7�Lh�;��Q��IE��&6�m�Z.�(�4�˻��-�Jѽ�&ݼ�.�/*����U+i[��Ѱ��݊�,-���@�A��C(�6�Viܭ���6��k풱YU-��D���˺D[�^��[�s(��NƍȠtN�9H�u��;t�6]e��s�*�۷���$���hYBHD��Brn���A7v�I�kJ9c+v�I�� V׸%�qc ��U�f��E8,�a��4!Ji��l�J��5fK/d[w�n'c	���.����O1��Z�߭n��0��[ܳA3	�eͫ�[Q�I�0�aT�Fh�=
�uf�����o詔�[��mT�L}�FV$���=J�ޱ��k�kj���w��,J2���ϓ����͹�VOZP�d� �C]L3vi�+��d��lı+�\��1A���yN��	�0�(�m�35YB��y�ٳ;��SiF�D�x{�U���V�oIԿ�fAGk��m!�����A�Z��Eo2�����e�v�X�7�H�ZY�l�d�n�T�����jk,�C+p=��Ű
��m�ٛ�쟄rՄk>�.,��@ԖRW1���I4�em���[Y�����03{ �\[�daqbWy��@�B��+i�oX[���H���ed�ñ=��V�#ǧ]n�*���,�l�v��n�k囹��4�����٪f:t�^ %���2�t�Y�,��[;R˅�*�'��h1���6iv�5a�w��mTӹ���P�'������e�V�*�(���=j�V��3��.��aoKL,N��wV�M^�kT�V/�{hD�0 �Ƀ.�WYRRR�^c�b��XF���54(*Sq<�;�а�S�7v��͒����)Z��$�Q��5п&?1b�(�Q�F��0n��R]�j�U!ՍIZ �>F�ĖLE���-L���j����l�c\��J���4�c���OJU�8�_-��!"o�Ӭ8Db�U��m���_6�WM*i��ٷ���7.�Չ�*��-"&���jYLH��S,�v2�
iiA]lݻK�t����5K�#xЫj1�[P�X��4h�4	L��,�JJ��Z���i��.�-����A�si�D��	L]�P�X���N�P�ܬ$�ŧC���������m�!@�CKQf��-T(���%ފ8��\3 G:���z9;ND��Jg���x�z�ՙ�5&�4�ԩ�b;��B=���[t�YeT��Z��Syl��[�k "hAE,h%�
�ա�v���Z��F�M�c �,m�)֔����o ���1�I0�-����,�L��t�D���qQՂ�QK2�ɁMJ�\V*�f��*˼ڵX6���n�l�d��Bc�ևeC�n�ԉR�-�n �XV��Uz���T�U��r;��!�����f7H�M䄥d��V��Wu��\��n�%i� 2T
6۫5�_[@��ÒK��ԧsQ-A�)��G����Gk%2�휿�Գ��Ilb�ٵE�� ��J��*��&!��j�Ǆ���wo$v��b��Y�XS� ���`�Sm����0⛶cE������Q������cq�+EmeB�CY���]+��AZ��YP�P�;�v�,����R�+K����\���(��c~�-AO*�ٙF�2�ˁ�(��ͽ˰���X�
�!��e%$��L���N��
���b�P/U���ɱ�Pt�X��itK��������ܹh�
1���E"Y��hj�,�����,)bĶ�X!9O6�h���-"2��%\��5��ͼ�ݔ(���u��=#M"�^G[�-T�
rZ�X�'A�Ә%,�(^��u�.����֘�X�m����� �pR��X���oNP)�t�B̔�1d���w*Hݜ0��gf[��,��	��w��ľ�֧o�|��ʸ��w3Pb�6)���M��FV��S�s]�7WA�2�9Oo/*ŀ����\�P�q�v&k�r��/2�T
U�VU�QYp�Hz��cU�駔�鉋2SŴ�\]�P����2m�BK$d ����X���C��{.,�N^�h+$_bJ=��i�F )7N�ٚ�E Ohn�9F�,/sg���2!-!�,��x�Tb��h��R-[�����<;Z@Ah�YJ"z1��c���I9i�vҍ�NZ��)�6����Qd�M�A+n����B��2ore<�4�ѭGi�ӥ���0 2Xql�л����S�V���vi�Q�p1�e0NHq9FƵ�J��]^�Ū��FR!�2fa5`)o6��L���2�����(Լyx��o���.��QKI-�*<�'O�*�eq)��P���r����㵆�l�؛V��iW��I�����
��vP	n+��\ج
#"`c����6�,��m�yv��[�2��۱x�el�'b��R4�Z\3rk�12u���"";mm^v�9Gz0c�
:8A.Y���*�S����9s+Z��7�V�+�BP�up^�@��"o��p�p�6�aS�8ݵL7��ڶU+v,���OIKiV�m�p�gu��j
i�"�k6$ifenG6�6�-ܢ�m	��Ni�Q:*me��aF��0"�+.�kŕ5�ݙ���W��(��V��i+BȒ�I���h�V�{[��T�ޙ�ch��u>�ŸN��P&jU��h7 �vTu��B��ǃJ9x.��XjaT-S�v$Nm�V �q���L6&^�Op�F؍�k,�;��w2�a��.�@X`�`I��Q��b��0��eȎZJe�]�n�׉[�]�e=�k7ƪ��f�;r㧹B�΍9���J&�"�%,rV`W[yw>M!�O0˘�ƥ)t\R4���
֜� ��ٵ{0�(AG0R��;C��EHV:@M�ϲܧa�SX�-}r��S��^0g�.��x[����WX�XU-�&髷��������R���Ae�ާY�J�3�G��6�Z�e�������R�	��f�Q�0M��e-��m�f��Q3SciP[�<���mOl|6��S%�X*%���sۦ�n�e�"�Gw72cVF^�N�&���unW����KkMC��b���i:�L�m:�V�E����v�7Ȥjei�+$��2���PM&bnt�A����(=m�{�d��	��f�e^f˩���ŗvI�YiQZI�d��Ǉl�d�V��i�A#�hhǉ�ݑK~ǫ\t�G��:��+м?�#f���҉�-*Z�i���#h͋^��k��:��U{��IPb�1�4kg%��Wo�^'�s
���p+.VS��n�^�P^Sm$�;��/-f&�-�L`��iѭ���IS�'K
�jr��Lq֣���驣��ikw�K���cՓ`ii:{W6֥`n�/&���X��o%�w@C��@�� �kr^�e�X�8mf�m��v)f=�c)-�E(��U��	ޫ�IBJʄ|" ]+�=ײ�$b����D僉���7�A��H�1��S�{5�w��bu%A�dӱ��TB�V
K����x.��#x¡Y���MJ�B4v��a=ӱM#DB�:9r�/(Jwen�. ��YlWzbNށxb1e$Y�x)��A�E�c-�xЀ�u�	�4U,��ʕ���k���ᒄq��t51X��"7�if��\�����՗�oW�fodr�"wi<���Sis]{n��oo2�:xN�o�}�G�Fnܱ��ԛ p�Rs@������;��� �S��mf�c١���+{���H0�Y���_L��]��&��Z#���r�����յ�Ճ��Ø��;ݵZ��r�^WӟzX����<%e��X��ɰ�m뺊"�� �b]�N%���'��k�-Q���Q��������b�$� �	�G��8`᫴=6�n��#����GoDng�E_v�=�D�d�f�g\/Q����%��M�{��9,Ӯ�Ubc4�����4�T=��%k��5A4�����0_:1=�z�
���ؾ��V�`t��|O�ؼ�����2s������c�<�8P���ӹ��}�gY�(���v�Zt2�̗ɣO0NO�7jӐ���*�li+7���(]wA\�o[���3ҥֆ9!�m�޾-*�3�]X�խpwbKw��P��|[L-��wVe������D��8��y<=r��t���eq�1:�;�(���+aSZG����^2^����ǐ\���ڂ�5.��#Cw��<Anuq����k����*ۑ�㬮�YY�h����5���݃\�;�bQ�wU9~�	e��4��!)w�7�*<#PE�z�E��>��(���\M�`u����ffK�x���1�W�w�^bfB����ep�#�Z��%�m����>�b�>�\�f����95ȃ��A�75��u�sY�ʠ\��Pǽ��N}7���:��u>jIN{t�YX��g����-Z���r]�k�+���nwP�D,�Ʉ{�������S���)\�)/7A
_a�z�니L�q��t�5��Qj�[��r�i�\��or��P���9��YLs}``�,5ϖb��lf/Eg���z�ށ�o��BQ��Y����,�ǻ�� �T�c������@�����,S`�j�|�^"���=.����ո/�m&�7ޫ-�ru���b|��������<B�R�W��`��OH��}�`]Ւ�b����2��Bdē��4-��V�Fss�%gMO�>qǀ�����k{���#�"�E���K88t�J�u�g�Դ��cJ[K�Z�f�"�>K�V�i���Ze*����঄ͻƘ �2[ި�F"�4��w���G �8��w��b�P�kc���(h\�tzw~Q�� ���WKL�eA
����t������(΢fHl)�)����W[�V��,��2��f��]���Bq����,�=t��ܫ����b҆�ic$9�f��쾝�3k;r�T�;i��u�$��'���w.�9�.�W8���sK%��SֆsL߫� �I;�X��OB�Ԝ��[��[W�S�F|�A�C�A��*�!��c�Y쉈�Ϸ{��Ny�(o�/�:Ҳ�K��'t�C��V��la�1��Vx:�=�p�8N>�@�%��i̎�0��Z��D�n���xl�K�RN��y�Vn+nqݍ ����b7��d?a�;1�p:�>�9��k�Rv7[���FܶK���(]]������[`�c�nP.�	W&cf��<Q�*8m9�W7��x)��ڮoeED��i��Y�'�U�XM��V�0N/�v Ba<t�ҷ��1^�RZ�)�r���"D� H�(����,�f��&2.p-��U��!0�ױP�c��8��XZu�;�ۮ�p�5�;lE�
�Q���3G$y�~�<VdNUG��w=���������L6z��.Mo���5D�_'۲�*U�������.��P��T`Id?]��6�f��cLt5��7�q�%��9c�SE���}���n����Qg���M��\}�Kd+�P����Wދݽ�5T��`o�E(X�M�O��Е��ޫ:�qd8���ͺ���:���Ҵ����]��`�����h�sow��n��%�hg0}m�-2��(���(��W�+��j�5�K9lY�V�\���$�;�%�a^W���_���,17>���vio�+z�����h�R���z�R�3�rl޺��3Hv=��-܏�h�H�m�C�Eq�j'���lg�Z%ɠ[������cKL� L���s3��N�sF���n����x�i�i��N�c/�^�x!�=����r��c��sc��ۢ.��	��J,�5#9���$�:�R�%��fm=p[�.M����`�����Ox��GxR�iT�r���t����ծ�G:=[Y�Zv5Gq�/�����܏�7g*Efফ Բ,�]��I��n ��R��z��D�\F3٨J�vx��X���Μ:����f��V�}��L
4ebu������8&�3��w^���=��diV����ܨ�f��w��=�x�ܱ�FZ�Elm�f�e V�2eg+�h�ª���O(�y��:�:�pm<wS����73bͽ�����8�SHZ�S	Z���Z�q��Ǆ��a�+&<�f�6��(�{=�I���i�)^$-�{}ڪo�u�)>��޳������Գ�v�z8	m:��w��w, ǚ�f��L�Y�����X�rn�$�?6mw�#���4Q�^����켑�\n�h}B��қc���i�H�뵂f�D��iÔ��m�Ϣ��#tH���3�3�hB�{�U��Q8n�'7�0�0O�𣏕�����*gEKg����Sr]��T0!��:��;�_ CJ��:��k�2�S:�q��f�4K�Ft��Հ�|m�n���]��d��`y����YQ�V��U{i$���(�-7�x�κ�����}�E˛��6�ocZ��k/�=�Μ]#�oM�U�U�=����Ei�@��K��e�mNd�歚��W��stv����!��� ���V�畳u@�I�b��;�ϙ����o��~N1{�Wz��l�x�<c��������{:v��J%K>�`�R����d��n�������w�+�=ɉ��j�c���rD&�[�5׆��Su��ݢ;y�9��N⯯��5�->;}�P�=��;V�{|B����Q��s_V�z���*	1#b�yit�+k�=�(���9����Q���4֊�}�IԤ?$���H�]��ŏ�htz֝>��V�#7͓�^�|Jq����N�~d�
4�qK��t�e���B�ڏss����_]�1 ����| -ب�4���MUǬT�ѽo*��u�(]�鵩	2$K�ȹ�ilV-"ӱ(�m���
�Y�=�H��[��V@�VEA�2�h\�]�f�sQ3ކr�{�]LL���>��b6�@BS������N��k�Y�-��\��������J��Ʉ������;�CN����į��ܶ�:D:�ꡗW�����gK�j���EuϠe�����ͅ%��.N1s��F.���3�i����l�mL�M(֫ظ��Z��/�o�e�8�y��sz�Kl ��쿈�Q\�����e�ңt�YTl&X�ܬsm^�B��[V�ܙ�W�|�5��5�֦��Z�2�_$;^:];�dP$��0owEgB<�,�G�����9�@ړj��A�q�4�e,�oVAb\���G�2���K�=S����&��W��dWM�;�JR��(���9�9��r�#m=}+���k�Q Ψ��A�nZ�4�j
���2��t�۹��=��Qm�T�0W@5�#�2���E���H�ҏP��n�*y����wy��C��^>�dEdKq;�<����2��}���z��}�^u+d)b���/�y�.�h��-��ꍻ�;n�����S�2��s˨�nQ��P���%�ǧ�+9�QZ$� F�'Pޟg8�R����*��$7�r���M,5�("���8�\��]+��cv������O�qx�mb4m��xtgv���{ӱ�27Y]�c[�Z�b#8>xp�5ռK���������P�/N��xs��C��GW��t���Xv�m[ۚΣ��C�0���G.fMk���h¸����ڂs:ͳK1]Ǘ;&�Y�E���K��]�0���z�.�,�;z��9�yZEŧ"R�sM\�9�	�L��\�k,[T��پk�^]��{.F�s3�t��k�j����I���wcIm�f�Z�s:�� ;L��Z�n�YY����t�2�V^���Ch}��)�m���� ty�h0h�WW��;���������5hşn��nP�i��C�"uϔ۶�k붚R:|Q<5��W=g5���,(�C%'���Lf�)<W��ai�{Nb�ʲd�#l��P�����е���z��^4�`]�҃��Xa����ӣ�\�#>CZ���}�_�7�Zs4�5�]��B���W�._N�Kx�B����������C6�s8����[�[|8?�!�17�39Y��X�]B]��l��OUՉ�78�b���;�{�ky!`N«K��:�D��"Ii���:���i�N,g^�^}fb�r>�ekI��_j���n���y#�؎;�ؒzn�To{��>���7r����4Q,W�}�o*�=D�y�O*�;H�e��l�-�|��{u0Ztr㨱����J�����t�Z�N����g6�z�u�����)f�rzua P�ւ���b�]CJ��\V�s3\�y"�����Ƴ��s�nY��V���A1
��42��ijmv�hk�m]j�u�uc�L(���K+vj8�.�	�9b%�S~�y_^�Z�=hFwgY�s��=`+�M�B�7�B~��|�s����ޡ���J��t��P��n���IIw]Y5�=�#�q:E��T鎓���\d�!��7���z���'�O�(w��o�R�
�7s�Zww���NZv�o0뮏,��z�N��n����d/��K�5���|n��L}L���=��0��C����FhQ��^ׇ4+�i	
��	�>��{�z��NR�F���i�	��T�����6�S�������p�>���4�k�bW�������/e���d�e�����\����*MV6�&�����io^�ݖ{�[���C���Ϲ��X�t���;�Uv���V�3���{{ױ
����_n�=�2f�=��sAC-m-S���=�˥1<�����Fnڜ$hiќ��2�7����t���VK`��+�i�*7w�}����^�Oi���8�PL�ߺ�5�kV��q�aO�Չ�\���px4u�[�!|�|/���:ø�΁��8k2�	F�����
�͛�|��rT7G�R��)vn�"�9�w<�>�������錻�X���&��x7��{e��Q�#3��R�ze�x�:e�әCg����U*}͵��f�;4�M*��mj����z�4u��8����hƅ�adb{ӵ1�[�Z9[=AX�r& �=5xqT/��%���vL�����=Zf��9��W�e�*�y����礙7n��x����Mx�Wu�:���e���kY3���9|q-���8dٛ�q����&���9��%X ��\3j�����Z)n�6M �JG~IXQJE�y��.��
e�!�t�ڞ�}s����s`�{�����z��B�[�t�1���iq���Yܒ����1>T1p�|��ؗgo+�����r
7s�K��p�M�0�`Yaj�/P���c/z�C�	{7���h�eռ�c���� �ٸ�{h���i��S�bZ���Mۢ
f�J�(�նX��'��{�h��zo�&����[�S=��W`O���%oN-��)]	�lk��8��b�����q�Q=޺���ƣ���*�9�F����]��m񵏘����t������{�\�W>��+�S8��x�Jӑ���Iq9����{�m������Q�g�q�	���_W�@u�,�N�z.�A�<�&h�:ݎXTͥY������+Lw�A��m�P@ٽVE�,�BT�~>���Ӌ�����]��s���X�i(�P���!Y׭�e �[���vQ͸�v�f9�'Wܺv]P^j2>�+�޳-^a��f�V�atܪiar�ɶ�e��f��X��P�����[]�}t(�MU����k���f�.v����V,�;N��e@��p���b#�9�0�̬Ǹơ��]nh�I�fX �ȍ�W��m�=�b�-e�8�:�u���+f���װ�b{V��oFFq �J�.\�S�� ���L��x�Q숎�t�S-o��t0�w)<څ@}��J����`u<g��3��Ӆ�����]�^S�F�1/���MY�;D%�*4�����v�ɬ�w�{7UE�mයVt�Q�-�W4�ۼ�Ò�%�"�yk���ߖ�`�
��}��-uM	�F���O�'!��z�iI]��A�;}��W֩��ɹ����Y��'v�7��b���_Dz�F�}����n𱜋LXk�]���gmg
8�&��*:bK��C�{���B�21�-��xN[�y���>��\�AF�J��1b����/EJ�<+~��I�@��ӏ^f�y|ڧ�nM�V7DooT'r)K-[y��G�GIЁ6�Evb�"s=�W&29�d�̼������G~V��5�(��K���9ڰ��J�e�����5��yXlяNؔ��l47k�f �-^�� �����*�tޮ��O*�^��Iӛ�s��FΗ%���U�����|�2���[��i͊K���u��K�"wU��o
`�"x�N�;��:x�v�]�É�P10'}���i�ُ��Zv��yj����^{���^Ў��bM��v��@��}�����$�o��ޚsU��o���o|ֽ;������/�Ifh淹D(��.��4�#[�kᇶ��+]-�Ȫ2��w�%:Z��{vx�F�F�ޅ16JD�3��(��Bw1wg����=LRzMm��;�Ϟ-�\�hs2V�����\k~:e�
Z�{(5|�i��Mi�u���z_	)��.Z���\ۍ`�#@ܸ��c�[�*��M���E��8����z����ܢ��Qem�Ov�'�u�ʥt�����	�m�瓳����E�Hv�E�h�"Q�&D3��!��J�;�=�{��+ȝuҦ�,�,��!T���Q׃Y�#:{o����$N�i�J�E��F��I�.��$�>�K���GoZ
N��|��k5�G*�����N����֢YT%� ��ǉ׎�Oev�Հ�	mF�Cؑb��c�������wҝ/���gl�!��%wf�T�K')scku[�����쌙 X{��Z�I��c"�y����n�����Ҏ=W!����5YY*V�e��͹�sZ�-jP�ayˬ7�d���@�S���f�H|�Dz�"U1�س)�mb�=�Zd�;$y��0̼G5.F�����J�v͠��3��b��]��u�k�Le�Z��-ヶ��n��|�]�;}2N���aJ��֐x��w݃CYt���ŉr���y��S��Yg�0�+V�����n�m"�ܗ��M)ն-�"U��opvlzte�
�,)!�������}+�)j�Ѭ��Cmc�#֥��:ˠ8&���}g���Ma�2�����GaV����mӳ����� �Y�)�kY�_ ݎ��Ǐ�Ws�})��.��S�|�����V�r�>���d��*�]����&-՝01�YK1� 摭�U�u�fϣ���X�y�B)�Fg
�S��X����+7l0���F��q:�F)��Ż��:T�[Ժ�]c�J�.��ݰ�Q�@]�����PV]$Ȃ�v���N�H������/u�DTI�B���M�\��;�<5�;h�A,>�}w��ƸAJ�T�4�ꊹ��fM�V�f�j�{�opY�g;�:�����a�A��99+����a��_>��s޻9�1�cU���v��sx��hMǽ��){�}��03i9'��'ϦjX4%XC��hW���*P1��dT��#Iv�����U���
�͗(�yk3��JU!�^��Uk�S1�4讵���;A�|"^�5a���Gf��7ǢwZ��,�9�;Vj}��)|�+��V�3��{^�un�X�Ҧ�����rM�q� ���������A�&קRor�d�j����՘� �X��og'ٷ�2jوG6��QQ��T��|��#�0�!��%wW}te�����7��tƗJ�,���c��l1b؂�s���+�+ {B����5���T��!,w`�~���ۗ�R@����T1����Co���D\��1����lgfT��9������Š�m��PR3�{�.���.���,k�m�.�����8P�7��n��f>A_�Z��0�iW��%��
l�(���0�FV�;��Ǎfrۃ�4pT����0^��g	3s;�t�Vn����k/(�= A�d���^�9�5���e2�-������F�YB�n����c�m��5ݧf�;�<�fW �v�쾧>ĝ�<T��6�kS������m�]aR����}p͝���&�P��*Ӯ�q�$kvˍ����Ifb�G/2�A��:5��x��sF�N��w)9Ɩu�(wm˱z�ƚ[޾^�<�_�w�nU]��x��b�T摵���m~����}��q2�e�ćh^�Q`��i�Օ���͵�ԑ��ڤ���"��}.�=ˀ�X��q�0�`�T)G����
	P��핫��Rbz&~1=�I~/~۷{p[�[�q�?;�gl�v�4Q���t���2���ݝ��V4;x�,�^z��V�0t^K��N��5��qGGzZ_�h�[N�X8�ڴu_'��5��n[�G��Źt0���I�[�n\.�r�����!�m�*-W���,�S����;u�V�'p���#J���Y�:8�i��@��[z���Qg�����:�]�B�6�@��!��ї�K��Í�10�%e��{+���{q6���҉���#%�	�
\�
;��K4�A�34:{��J���/��M �]�PN��u�Ҭ�݊b�ȶ�;*+
�Kݵq��)�a<����g����қ��-Z�z<y��ͭz]�o��7���7J*l����&�jZ��ow���)�`MjD�gKp�ʸ�<+`t0ud��1�$�7��q�������Sړ���e�⠋�:����V�Շ�k�K���7�Gpm8�imVW@�Y(�{�P>{�郯iXDo�pC%���Y�J7m(wh#��3f�ko�ƛ��'t{+:������D�t��-)S�i�f0��3og��k��6�Ns��Ĥ���nѧ-��E8�xڼ7��F��0dK�a�7ʮKU*u�l��[��])9���ky�\�C�X-b�Q���T����JO<�!øU�ɸKL>V��uɑ�e���MhXO��^������k R�!j��o�$��X]Yպ��,v�7�X½�'��f�c��#�w����T�`}�mg\X �_�hz��^@��2r���T�Ǐ	ˈ>c�M���%J���ݾ��Uvq����}fk��2�\��G���C�����L����s�Y����ޜ$Ҽb����+��(9tdd��xA��"o6���v��
����}!̅	�ڎ�)X�b}�ذ��� �oN%z�=�Ε�Y�^"�u�G˜�ޖD}�'���j�B#Ո�SΆ�Y�������S��@��<a]�iJ�żK�n��Fw!1:��s���M[�CƷ��Tq��]�e�k~�r�M����*���]�e�y���v�����ӦZ����1�{���kAr����>0��������۷�rm����jB�ޝpeӽ(Z�뫌O�pB���C=�*�DL�R	�g1
�2�%��w�}$|�C���y�:����A$��B���@�@l[�)s��/0���V��$��+Z��er��Ec%���jd��E���)d��`U��r�y�{%&�a�*��^Ѭ�k+Z��oa.�lS��_-�c��G\���� ���@hx���#I���Յe�Y�΂آ����W���#�(�Yr�:#�F�Z���u�[|Y����2̽�މy͂�Zv��n�ŕ�����f}��1�y���l#�O8�P�f	�i���c:��T�P嘨�5s ���c�NI�_U��VJց�� ���Q�Ջ�71�y�Xí]�����
e�C[�c���'���K�U%ujN&��Z�]p	�b��%P%��v45��|%��\Um-{59�ڽ��ߚ��fFV���Mv*3Kʺ;����ʺ�R[NݵOF��G3���Y��a&�/�ὃ�KL�c�V����n �΄�o�\�X���Pj]3�ț�*ŗk����a�͝s�;"�ԝf��^���MifS�(x�+2	L�5��T��eW��\�DPz2���&!��%! �ڷ{�l%�ve�E8$�w�0�թKr�4�����.�pWG�^�� i���lF�.-4�b�4(�}w�	�RY�F�k&�Hv�)�Ğ���]��϶��D����z�A��t�4=61��XOx��y-��뫬U�`�^��x-��.�{��٨�ՇH{�w�Z���E>��:r��F��������5�]����]�Y7��h����4����,�$�ه�m9mS��μ*ħu�� ���z���pk��y���2�Fs��/�A�S�����!̘0Ej:�ʺ�7^��i�au>�0%����Q`�oMxo-����t�����8��n��hѻ��ג��v/N�Z��5N4h䏎?��p�&|F�C����h~�F����W�u���WZ:�T{H����A��z8�d�����އ����O5�vk���4sW��C{�7�V�I�v�M9��K��r��9�Xp���ct%;'D�	�Շ)!�n��Ç���_$KVV�j�s8������#��k�œ���1�m�=P!/,f��V�b��@Ԡ,�"�ɬ���7�|�h�ܳ԰��l�H�I�_cRG�]�y������s�����q��AhoHmȩNβP|�i׈k��h�ӎ���PWK�ӎ��M�ɐO�4Ԛ�Z2 ��;�%A�=t�Md#��H����8+"鏩�C��BUrF�&4�����B��&f��)ɄN��.���
d�^�?mh���o��}�b[�Ҭ�:�wϗP�lYo�E�Y�f	_<��~�B�z텎��^P�^��r�V��Շ���Ǘ�Y��̺P�E�&�����h�'��I��{�Z�Hh�c�{�-�e�����Y{Smv�_ι/�znt�vDh֫�+��ğ$ҭ�[��m�0&f�{h�7+Z��r�dn��Xe)���Y�T��L7â/{��vm����u%oXb�͸f�˶\����/���+��ᳫUo�n�!�v�G5�r��]O`��������yL5�!�o�v�7P�B)�v?<�˭$_
�9v�����&��o}��=������N��(m^>��"<�c��d+f��o��V�n�a��#������p��i弣��0�K@���D���{e���GM�L�`��[ۏoa���Z�'�ź��YBvU΀n���w����SSXv5��Z�e����W�B,�L|�"�۷���K��a͹έ�6�������E��4��[&\ T+�(��Yc��ɺ����R�R�R�9Yr��Y����=�~�>�bVz`ZrdL.;;���WQ�S�p�o�w{]ru�����T��j�j�۰�o]�X����M$�T���O����
��X�2�Sr�	Ղ���Jt��6��%�_# �J�K�Nr�4�%�u������p�up;&�*j�X�]�b�)��������)6�v�����`=��V�Wz"P�}t�b�fц���mU�y����̩�Z�0A�Sj̼���A˝ ��mQG�+f�ة�/��뺅�	-i�x�xB�p��h����J�Fj�l��W����f�ϖ�Vq�������'R�A&S�c�_������`�͚GE��{�1���m�\�{H�n�s7M�����YW������	T��9�x��YMu�*�|���iVk���_m��{��"��k|��`���AL�XC�򹔕4���/��+:�j"^ГN��"�:���)��]�V\f������90wD3ե��79���`���u�7�X�j�S�!�x.���K�Y;�e��V�i��wY�b>�nx�y#����%sM�٫6��Ҽ�\�c�6i�yX��a�)��:���+pj�]�S�i���w �K[��V��=}�[���l���)Y�c-¬�u�D�}ү8RSKʹ�I�s�]˺W\vZTV�W
���si�tpk��v��fҸ��V�G���+��v+F49��~S�Cb���I�X*pӡ���	Yd��5�2�lt�l_�=]����}6+I{w�V蓸��.���������=�XR��1n��OPsz	����t��n����8g}:F��Y�q���l��:�������ͱB�B_Y74jOk_D^�����l�;[�
���H�x2ƷH�n��'QT��p!$ȭl]v#���C&մ��Q���(��ç T��CY���w˒����˹x�ٔ�R'y��a�.�ßn}��Xo[��cAV����c2�7[��&-�ۚ��%bx�_"w �K�U.�"Ow��B3u�Ӭؕ^&0�x*����Qӆ=RdMt08r	I7�a(����ח�JP�Q7�(�X���ˠ�$�|�T����m	me��2�{�N7o���M�V���:3 ��:����Di��4�е��I���WN�I���]d��\�ugEGHj`�J�r���fn��Pi�F��c�Hul7p4�:3����V2v\ax[����ͧ����P��&�|���b�O�qh���h�WC��+��雷��J�Y|��\�)ܩ"��0!�o*v]��I3�F̜<���
�6me^}2�a����$p_t�+�y��`�Sw��Kg�O?>��Ƹ������8��4�Ь7�p��dK�m�Ja1l�ή�o����8�� �@Z�ѧ�U����ط(%���04[�BEt�?n�L���k�*�ic���m�%���_��ns���c���eXж��L{K�$/���O�xu��d�u����k��s�b�`���n�TO8f��`=��GI4b�4�*
���l�q�DM*��3-E�V��nFw5�k'A�����9]Ñ�����Ic�H�-:Bi�j�m�;L�.M5��H�N;&ou����˜q��nk�[
�����Y�lw`���4Q�2��T���K޻j��v�d��^�ͣ[-]k�ܠ�h�u*;-:f�J4�Q(0b�y��E;$D���;i��8(�>bQTỷn�)�n[�Zxf��2�]\Q�J�jv��vl��ʜl;�Y9��+wu�p�m�'��t'`�}������\���j
�{��b��
b���5<�[6��b;]o6U�G����n���C�%�m}_}�W���*��d�zn	��{�7�u��&I:�:)�|��(���`��.���rv?��R�w�����9/uu�F�5�K�{6���]co�,wWj5�5o��T�E�{�U�*��ӛ���w�vʾ�c_9�X�[�;�j�s�/T%5�68N3��mJ�ڎ�d��j���<��J���)U�g��d�HT�f�՝څxfOo����"�Oh��K�-]i��֧�mLG�jj�zjQtF�r�^R���*H�j��!f]����gx�����v�����٬�֫W3KH0u饝V���o����]�g���%[�s�P�P��Lb������.��N[�j���]H��d���jVİ�W�aC\u��r�=\��q���6>�-t��õV�w��]9��4�u��X���u�tj8����;����䐉�����*A��t�_'s�.�qp(w5��0S��ڇl���VMwi�j`cɦv��`����sw[r�tv���F,h=��Irj쳜h�^�����"M��$�5�Ϯu��wL'�	��ݏ"cx�٘;�JEy���
��m�c�Q���%K�\x��h�Se�����7e蝜�2���5��8����]Y��;�[~�����F�U51�wAX�K�sݛ�=����ػ18�P�c%�(����Fe��Q�Q_Q/M���5}M�JY��~�@��Em�,�
��j���E!R����A҃l�H�i(��Z�H��,
��*��Jŋ
%�%m���Z�-��`���E�E�idT�[Q��QIY*�YX%b�)[����X�Z�*�kjQ�l��*6�����Q�D��`�b���YIYU��Aj
)Z"�X�,���D�Ւ�+�\�İ��b�֥j����jR��V��E-�m�k*T%b�d�"�%����ҫUeh�,b�ee�-��Z�V���"����������8ʣTU�Z�EYm%d��%[m�j�B�V�����+
��UE�"B�m���j¥e�,Z�	`�H� UI'wl���VIr�qǸ��:�N�v�5a�(3�C�Y�-F�����7��A��K<W�ڪv(Ƿ $�E�:�`��	^�H��+q�6+��Yu���T�P�yH�!n5Ag"+ڥ���������D��(#^����?��5����1����w���?B�b��E���̔_��@$r%����VI2ԲV��`߅:����}8��CL���ڜ/�j���%�sJ]�4�1Q�8,w�(�� u�������3
B�%StX��bi�]͌|w�|��m�588�Wls���I�P��mY���[�|�h����P.�.7��ִ(���A��8k��i]1I��R9��׽_`�[��`����� �ub��ͷ<��J��3��8!U��7�	DW�X���M�b����Ma�ѥs����g*�Wv��6O�8����W�}_�R�~A�j�rv����W�4l����q­����ew�������/����o�S=p��a��9��X�]:����\�;B�(c�Y�-��q_<��QWLeƪ���@--b���SY�D{@sg�bt�:���~���=��%��N�#�ܦ_l�w#O�9`�6�'�6����p�u��ڱ��fĳ1v�ky���L��h����aU�Z���7��	
˗�6lϦ-�:��74$��^"����k�Z�ʓy�7YBG}����ɫADڔ��Y�,Cͪ��Sy�_�-�!�m��q����&������n�&��3�n此�M|�!�*[�ns�Q*�h�q5[�=�p�Kv����o�P��ov��^�_u��kvh���/�
���hIU�Լ���;H��@�� !��¦`��S7z��r���s%��p��Q�H�tШ+i��%#����6��_Ϊ1#l N-Y�q��j�t�8�z ��]H�J���2���|x}(��S;� VZ��1y��Iw�2V>C0W�9�!e�o#����{�%�*K*�M�
u<��Tkl��T
�~��G�Kɼ��^aL2��0�*f�.���6��%��y�#Z1���؞�K)�z(3o�{xN�s(� ��:M@C	����W%�B�mH��շ�ȁS`��|���h苁�eB}M^�R(���\�W�Mk�j�� ;�r����{ΘAH#�H,�߀^�􄯽��<d�/i�Ku���_��j�:��8����e)d���!��k2���(N�u^	ŀn˼��İ`�:���n�c�E��QIM�;��R2ҵ{(_�s=d���,bM[d|�b�D]c8�v��s���T1V�H�e��NZ]۬��`>{�5mai2��-ౕ3.cL.���y�ۍ�MNQ{���"�l�))B[��~�]Y�IT��r'`�q�2)�Q8c	bx�k�ʷ��}k��U~.�W�J��L_[�Q7��^9ڊ��%�1�{\����)�>�X<���`�4z����ig�j$P��O^
����|���a���n�7��+�P�)�W�^����w��(&��K	4��0WPIm�uR����g�$-���#���/ez��i�#��J�K&!k��	�����m�.�J��uZ��M�ʨO����:�\b���鸕uÂV]������T���j�܇4F���q89��%q�
�����X)���wP��t]rŹX��jy��!*�A��<\ �v	@#����+O���x��_]2���5\��LE��u�QFsOq7��N
yj�\CuPB��݊*<9�T�������m�tœ���Q��}��u8^������1�8?y�g��>'���uJ�o��G��ĭ%[h�k��@��w.�dW]u���;!�+s�n%�GRwq5j�<��\���}�XrW��N@;cxV�T����祼]O<�����N�ѓ&�U��R*)���f��wO����	7��Eтnv���q⛒�-0Ը/��U���ו�l�<nsu��-�hf�V���Q2_Q�}�lv�oT����
+�����EF9cw����(F
�.w��BT��4�A�`�[�`��8Y'��
�\���7P��+t�V�d��P�5���q��1hȄ+�m0=�x$Һ�[��x���h�4x�(	lI� 1�g�v�\f��pzcDɄ�r̶*�;vf-'��V	��m�'��,�~�M��M����ޘC.&XXn$���A�U�Sړ�;����m�IC��޴-D^OTcn�N7'���{��3�>&�:-����i��K���U�8���r�u�5(j.;dk���@r�b:)͢�Ȇ�x�v�$P�1�q0�IBE���4� ������	���0�c [ߗ<�ڥ�[T��B����7�ò>�(��d�@g';�{4<�E1S�%^�Ƴ��W�����q���ZSse��fk1VV1m���������Y�gRѳZ�>�RR�0��"��p�Ȕ��e᪘��@��J�����G����NC����z��׳��,dVO� ���g�g�|�®��=*�SL�k�zFD�I��Rm�uf!��ISD�x�W�ľ�g���g����R�j�K5�T��𻖥��^o�;�Eu�u7b�M����#4XA�u_Rn�Y��l�؏�5�Ltb6�	�ҕv���Ϣ�K�ܞ>�0v�jv����.粚���(�v�o:29JE�\a��B�:CGN��z� 3e?F\(^S�y~�:M:5�z���U����s�D�N�1�I��O�)�!l3t䡑
B�ϸ.&��y���u���WA�y�L!ke���pX�x_��qS�X]��q�)D�<�yQ�oRv���D��s	U�&&(�xl��2���y�\�/��B+ରz۽T.M�ݫ���<��=ب�����T�� -;lLM.��za���P�RL֋o���K�p�}�NOqW��[������d:��E��E}��F��x���|�F0u�9���)��(s�H�4f����ٶ���˿�u�L�,���^��8k�����~DyfPmV]�X���s��3|t$���F=�7��8w&��������bW���l���͎2SU�q�"t�f��	���[�Ӻ��b)�h���=b!�E��Ks,��Ѯ9��4����b�	Ì�~��GLRrE���j�m��'�e'�ȷ��5�� �.S-y`���ƙ]��y/0\��DaV0������N���1 ��_Ⱥ���Vd��U�3a�b���6VZ�}��w;)�^=�p�y���-	�|.�6έ�f�k��:��B�OQ`ə�E-6xt\F���%g-m�+�0k�����UPخs�!�\���~g�U;ω�(c=Ð���#"ͫō��k瑅
���Y�|����\,�CG�7��W��E�mf��3ށ�vU$�')�G�f9��-�W������ٯG���D���H	��p��a�b��Ko6���5�����.:���[/M��\q�Tp��Ƌ�㈬ ;; C�K���%�k;mK�+��3b>�X8SyU!�4��q��d#�m�|nU���B6�Q*�X��< �>�;]��3�\5y�����B�M����dYߢ�ǐ�ѥ��&��K}[J\��!�������"���A�KA1������ʎ7�N��7ԁ=U�;9�w�3ۘ޼# ��p�m�7
 f3`�$f+��[.���_	��o�⫦z1<� ��U�y	��,��@�f���=&�e @A�l��90��k�3S�^�}�Z�=���O��6��Ҳ����E[��|Uv��(�S��G��~�̫U��ۑ��:�.��eX�F`&_Z;jEܜ���\�Cz��&v���{�>����/N��a�3\_J�q˺���q����V�ƻ���́�rHܒ��`��t��@o9M������/G�sl��Ũi$�����5�O�CRNx�vs �\�rcj1��̜���+�����v������Sa�u��ȲV�1þb�����E|�]u��n������&�Fv����Ň!L6�I��~|*dH澆���6�yw�G�{�5�~�9f�L=:΃;u;}L1��J�6� ���o+����^�TP��r��k���{\���o�e+�C�����o��)zR���h�3y�����u���B5�=!t{��l�'�^u���j�ㅊ����Wv�1�ʞ��&����n#�c�؇_h_{{e9T}f�=���)r�C�ty��w�H9}�Mj��W��2�W��3]}����{J3Jv���5�Z`�+t�\�8.z_���ޅ����RŋM�3�:9��Ec%��j_�<\
�P�Yg�c��
8"o5�|ۍǃ�������Up�N���.X� �N�b��0=�nX�]Rwdq['<S���h�#�yPS�RMA1�~@ĥ\Neb���	�on@N��Ǻ�j�z�*��Ll��p,���(�^D����/���;��m���y;z�?U�-K�fOa�1��Y�u RV�C����f}�ΙČ�_��Z�XW���X:xu!|]�gp!JQ��W�����ɆFM��(́Oj[�u����fE�2�!����ɩ�+��ޠ4W��\P���Y�!)�F?o�#��\^t.�(��76�X�����ٲ�v(J&ok�u�G5n&��͌J�7Du ;�b�ÝTT�<��%��uM>���5�M��\����*��L�cDp��aV�.EZ�RQ$G*{8^��Z��J���gn�=\�eJ��Ĺ��t���yNfX����j�2Q=Ws���d�e�o�򪞸,.��|�牊]1#1K�Ɛۅ4>���g�T��1`0�;s猷�Ý����ɂ>q��`�L��������刼�¼���,=��qB�2������?�1{��@���$
ͻ���~��0��5I��4��#D��L���:�0Z��Q�7��v��t��'��������e7�L!q/�)���΢���
W�Z�fc��S�*�\e*�����|�QD�(5������a�ɋƋ��C"L���w/%7�k���E��Ea�R7��3���ረ�8������n�:cj��.�&�q�x_��f���G]�BU�hd�oi���רj��V�����X����,��T���E�f��*���ʵ�9�y,�e�9��y����GV�;F��]�>�p���s��XH�޴Ң�=��]������B��D)���t��s|���u��e;9G5��a�@����ȍSL@�SF$P���8:��Kw�7Y�J�,�e��A�(���^��ϑ�+U�,k<D���k'�!�h�~���/�������jR��^<�X���n'���7��v}Iih��Q?���j��J��e.������jك
N��g6���.s\kn��Ä���NVȭ��Z�X� �W�]C�{�5f\t{�yS����[��8N[,h�;M�"��9��[z����6|��m��Kwk��N�Juo#1K��<w8Q��M��xhڄ��c
�9�~�Q%�v6\�.�,�u���5o����Z��~N�'��!b��¸z��,j<-��;?e��A�v��Fp�^����)x� �YSĈ�NyY�{H�c�����X�SB(>(D���t䧜mf�VGP	�7�*>�<c�\����M[K�h�i�7o�B_$�hz��y���d�y���1��wP�=f����B�2(3^`��.��5�<E��itC���>�q��P��!�5w2�1z+��3ԮcV��5Om�#��3|u���v�כ5S����>2�C�d��,�6Ք��i���9��9$1#I���"�[U�;
5�غ\&(��/X
��=&V���H1a�1�����V�}��\�f�(��9�{F;���Y/r�(��5�o���jP\�@�p��8q��Kwq
�#!�d�ό�*:��J�a ��Ԕ&��
���x��2�}(;��3��0�����y�^U~Z0U�#~��W�_Lȵ�ʧc7�{W`�;ƶ�8�1N�xՎVl�׆�c��ia�Za?���R+U<k����r+,��1�*r�
���Ō�b�!�l�'�)9"��b�׻U��e��#����U�yL� �C����a��Y�[@���ʁ(���������'���ӷeT�]��zt�r��p�=�7����<l��ϙ��W�|��R��x�7��^�*^�����F1����0�ˇ_-4ԡ�W�Ѹ@ �S|��\
��^k��v�9�q�&(=s	��ua���i�e#�&8T]1��=q���d����[�S�]�Z�T�qovM䠄,���)��<
[81�G��"��N��ӂ8F��A��3�s�7݃o;��,���7����0�Qg�Z���V�Ei���=�8�����d�Y����/��x��V,�yeo[���z�����f��<2�U�5��V���w�u=�,�yݧޡӾ�y�z����B����t����Ϲ����<����f�I�~fWVA�"N�G,c#��֎�I[�x�
X�{�k���\��A1y��)O,���nC����h�_NIXX�e�=�6N��`���<�ý���W��/1��|2$��9ٸ���D�[��a�X:��P�B�U��#'�A�W=�K�s�nн�6��|���Br��iu&o��v��=Z����=\�8 ݋9���&3{����' "�Ӑ��������R6%l�Nn6��,�t�=��X3F�c�'r����:��=����*!���Ӈ���ں���Ք�f��Y*=H�I;3�' c.��8tݸY����5��N��%qȸ�u��F����=ue%���:�_m�#y�<��R;]��o����n�W�gf�"��7&.xZ�8pH^��&
}�D�f�4�
4�:{����K��kpe��nέH�J��3��
��y�ZM'�k��c��l=�@���Va�.�X�&�A�L�˫��{-��� ,Ŵ�VZ[u��jݔ/5�/4����x3��m���et����"�AU�2��ُnX����S����c;�nNy�~Ŋ��	y�v#�5�`�-���HQ,��ϫ5��]��Q�����^cڼZ3�}#w�CU7t.�q�I�Y���lc��2P
��O��ۗ���v�fwT���.�i�.1��<�v���5�Ls��+���� �۷�WhQv���dIn55.�t���GF�;�c����� �]��a罵ظ�'jK��PZV*У���O����	�[;�\�2���GS���i�ΫY�KkE�]���x��^�R
����²�E]�7���S|ۋPu�J�÷ڐ�:��s�kj���^�j����p����;O�B�]�n�tw���{wΨ�yw�9��}��=R�DD��z`�Ֆx�|��8��ֿ��������u̇���V��ԊS��[õ猔z�Q9Q�hO��q�
@cV������row2�s0=�P�X����ŭ²�s��
�+�hu�}Á�L�;�a¯��C�Y�9���ף���ou������Ww[�vI�^���u�|�>/����O�o�<��I�lGCm��)�݉ C]�3]�D���gH�h�D�M��=�5�����4�<˰+q�*V�� v���N�y�r�pT�_���%[�S�zE���ӛ\���tsu��Y�afp�q�ʅ�yP�{�tЕ6u����1yd}��)�ϗA-�]Q��m�S�έ�ۻ�,kU����o6�s�pS{0Em���A��ăVY�<m/&o�r�-kR�Y���e�.8�;ٸU�TnLu�l�Ŗ���Ʉ�7�MJϊ�ؖP{��K����ռ����vYඔ<�쎬Y����P\������Ɇ�v�:�^�{���)���Y[�3***��8��$�dF�Z�k%B�¶�FЫ[+X"��D+�*���[�K`���l���T�`�#%dP�YX(-`�mmB����[J��V�B�TQKV��[Z��Ք[ZEYkdĕ�"�E"�R%�hU[`�YF�6��%�DY3("�T�j"ʊ�e�Z�Q��ʕ��Ra�PX���j�ʕ�m�TV�V�PQm�&
�TU�cj�J�H���P6ԩEk*H�����iU�j"VT�$��J؉Q�T1!DR*���)R�B�f8�,1��T"¥J�U��²�b�(T�e,ea�em
+�T��+U+��Ki2�
 ��02�e)J�kAd�L��7vp�Ԯ!=,[}��*��V��|���]Z�(V�)R\W�%�C`�4@r�}\�u���˼�{��za�^Ĭ��@�ķ�N��SE�} |��b3���N5�H*�"$��bOr�>�*N'�t�>a�Ă���CI�<C��XM*0��=�?`m �����<V|��i*s\é6�8ɉշ��}wv�������E�"���Iә�I���^�:��4�Y�;��q� �����'��QV����St>a�l
�̼C�m�Y�bOr�3�q�����y��� G��q&=>5��}]~����"�$����6��<I��C;���~B�?$�n�z�ed��w�4�i
�w��1欟&��c1�_�*?�"ɉ8��>aU���W�k����>�g.q��ߩ�/u��^�}$D�8���@�|��ӿd�P�AV;Oɤ�B�7�����i�~���%eg^��m��!��v�VT����t�^'�L��j�ɴ%D}7�g�F�Xz����B}#��ا̟�V��'��!�����4�W��5�Ă�zs�o����$���P'_���\�4���u<��A�cL`n}��:�!��?!�[8�����sE/ {�}�>���m��u<�ٵg�*g���J�M2bn��R\�~�i'�Y<�4g�LC�/���W���w�&�����6�l<V�B�lj�����\5����S!��c����S|���&3�8�C�g�H*����<C��hi��d�6�u4��1��y�B��.��kOP*N�S���������x^[ه�r�b���/��
��N��ޅ�d�4��<ԕ�V�Y���c�P�a�?'���m ��=q��ÿP�AVx���<B����P�?:C�{�<@b��>",�EP��V���n���y�$��C��sDڳ��L}�'���ɛ~���=J��d������Ld��dٔĜB�2u1�^�!ĕ�<=���x�Y�<=����0}C��|avC�g;޹jo��`I��c��0*��tu����f��1=C�~��x�U�T�y��<H.н�!���+'���4�$���&y�'���joVLI��K!5�����<��{���������ov~����!�6L�k��oc7���^m[ov1M<�s�mf����ZΎ��wj���/��ڷ��V����8�VAV7N�s���
�o�]�m�0��R��:����#J}}1\Id��P��O_|��������ɍ���=t��6�C�kT�t�_5��:��T4�Vx~��i ���é�a\@����8�S�>L��3�3�|èm �|~�&���`n���Ag��1	�����{�߽��ٯ���xO�4��N��=`(d݇�'��1'��q�{t�~g�}��0�&��d�$���|�>g���~d�cG�}b>��|Cn~Ԅ�!􏐈Ă��LI�
���/>Lgɤ�ݛ@�VJ�oY??$Ǭ1O�!ė��������o�8�<K����g����ʆ'̟�c���V�-)�R�����~��#�`�w\�=�!P�J�Y3��Ag���
i'�l2�$'穽U �`T�S��6Ϙbb����C9I��~�R�^y�P�����?~�5O���!w���s�} ��|G��O%M!�J���{?wT*�]��l��u
�!��ԛ�aC��YXq��)����C��vjèi ����q1��+�7�3�>La�����{��H��1�kz����}���P�H(t���<C��1��l���<I�{� ��z�N���&�m
ʝ톒�T�'-1�a^r��i�V)1�^&�E�d�>1Ӣ�vv�����J\�V�#���>���I��'�����C�:���:�O6��k�$�hc��i�T�!S��cY<LC��{�x�������8�$�/���!�K��o\0�y��s����>��v(bA|O�Ӷ�Cb�|�H�u�����P�����}�"��W��0�x�Y�O{���O;M$���?2k��t�!��& (���;����o��.�l���w�{s|<�˝�S�z��Tg�������Aa�=��v�ă�o8��6��J���C��:��'���i'�z��]�'��9�Y7��{x�L�:��&�~��?���ɬ�zks59�D��"�C�t* ���SL>a\f$�:����ھ&�8���T?'�bAM��1SHc�l1�
���Cg>���I�����Y6��Vk]�};^����sp~g��ʞ�RZ��.����p�&��)��)Y<�3E{:Vy2h�_�Z���\>�J�'�EV�r��� ��7֣�XWO�{SXB���Z��Ɇ�.�]���}�$l����X�Nmd���9�]�$} �D{���
¼�ə�4i��J�3̓H��T;�T3,�3��Cq���y�O�
��:�x{C�~M�q���I;��2|}f+'�1����=uw4��/�.b��@>�"$G��}a�����4�^�Ǭ1=��
�U��]w�l�!�Az��{�T���<�b,�5�0�j�I�*|��[I�+�{���X#����[�w{N���vC�a_�cﵘ��q��%�I��4����iX���᷌� �I�{�h|�C���{�f3�16_�h?!���o��P�b��S;a�b��K��u*1�#�)�ھ��w9�+!yR�Z=��	�'�Z�R|·�L��������u�V���<=�	�q��C��}�*N�U�w4��u1��+���!�La���u>O4���L��<>Z����I�}n��.��5���%eC���d��Tz��Ղ�ԩ<MSI��LI�+�4�J����!�+
��ӟwA�$�?�t�����^��q���1��֫�+�GO�5�i��_�[�纳��������?0*0���׉4�LH)���%t����1�VM�I��Vi ��͍���%f�}�l6�<I�P�?]�������^RmH/�?}�����2c3�o���_���j���}����|�§a�Vx�yCI8�O̝5�mX
OP���u%M������Y5�4ɽY��%�''���
�2j���Ax��C���1�a���h� ����=�<�����ߦQϺ�F�6���������=�18��bO��4��b��5�i�P����>d�'�{�~�Tڰ����Y.��ˤ?$��?=t�n���%J�N3J��UI�V7��f��ӿ|�|�`�F����@�i&'��N��� ���Y�8�C<.{�'YP����y��XTk}��%I韰4��ɉ:����U���a�4°����p�~؟1X�Q�jZ�D1"��N�N&��*,�7<�I��0�|9� �LB�C|�O�_�
���s�$�q1 �w��'��hb{?f �'�Xk}�!���xi�a�U�Z��+�!f�}i��~Nfr�Vk�2�^�å@�+��5���e f��#nzxQ�h�9eVܦ�<�Vݐ4Ʋ��^^�U}{��lS��̤r�6�f4q�݈6�%8კWA���F��$O��r��Y�[ʧ%.'��ص�:�Z�q}���W�xϟRc�;�4�U�M���6� o)���L���1�2���,�k<|9�	��B�y����U���<��~d�c�O;N���&r�a�{믢��>��^y]��#�����U;���T���=���i�xZE�8�C�<5b�H,��M�M��1 ����*uP�y2ɏ��+=O�HJ�Xxw����LI�+���5�X
��3�3Y�{{�\�k&d*�ýt��0DH��,GގS����>|��u�Af�*l�5��1Y�%T+
���cS���X!�3~d:ʚH,����6�����
�:ʇ��}i���A}�>�}��r��!���m��4H��DE�#�Dku��'�Y1'���*�2nr�'�P+�����*x�$�y�M8�QeB�I�/�'��]+I�/�x���R�ǔ:�'��c&�_�����]�z띕y������	�Y���!���V}�1 �0��q6�M�����6�YY׉1��}�<CĂ��/<�3)1I������L��+�J�'�OŻd�8�O�������9�Ҧ�!�����c�� ��?i�,ĺ�?~�W�L�4�P1��%�,7;�����d�~�W�ă���|@_�|�3�����x�Y�xw�LC�1S
§�x�=�ϝ��>�kwor�s�"4} �ُ�@|���A}OP��}q=����ǋ�NʿZ����K݂��i�hdfjJ�U�\0���I�S�U��'"=��
��NH������]�h���aOf'�p/\�~��y-C��C��}U���"�m��(���[#�N���XE���'��ҵ�Y���u�<v[���td,u�_��q?�໸f�^�ueSm��8��{ye���b��n�jΪv��Mԧ \m����Uv�J;OC��FR�8j�sٱ���o�I�Kz��{]K{;i�G��z:��M;�c�)�q���)uu������u�	�y�&����ҵ���uZ�7�F�syd�O%��Itc-�v����1���E��}�x�l�"`�8���x��+_
W�3�e����o�3��{0���ua�����r�H�<��
zb�5T{��$)F���}�.Ձ�g@���&����,����;������{Je騔���v++���֦z.��#Ds�D�4v@�qN�q7g�Z���J>�{g��?K�Tr�N/A���ۼZ����]@N5^d!�9�o��D�ܾݚ+D��
���hI�#R���]�}����v�M��n�&=�7�Y�n��p%�7���!#?WM
+i�#�W�2Y:h�*�f�qR��X�_`|٨ۈs	��pߡ��S˩�(#�jeF
��.�u;p\bU�cv�.)�-�Ӑxi&+�o��.q'%e��j���k虅�+�'B���}��I��y#G���H���Ŕ���e��Vm�nb៛%��t ���qı\��R�dG�p�&�3�*0*��6M@C����#���N������j���K�=J�1�uD cY���oq��U��N�xa�_eb��pC�.��v��R�[[����9��:����R�6��+��S5��xx�.=�U��,]�+6"�uNn�QO �]�}@�;
�yP������ƞ���^F`�A��NOWL;��hi;�9	�����ٮ�^��倧pfk��S����o�̮�a+U�J�/��Ds0E��W���%%�r|��Y��:��;=��
��-�T����i�]he���S��sq���f��H�c:���M�.+u�-w���|�{�1�r���H�R��TV��<|1G���~w�3k��`U�F͉T�X ��t���^�y&��L�N���gT����1g]}�	;`�:L�;�S�_l>�<e��Sp]&��|�p���f�ˊ�na�,�Ng*t$�\X��T���ѵ�ʇ��MK͞]�Ɵ �YsQ��j?VAШW��m��O��k�:뒻�Ty�XΙc��A`�Kh]'ä6lN3^�Z0��6��ʲr������U���Bxs_c����],��>�^�w5�|�^dc���n��r���˄3�Rx��B鯉@#.~���X�M
����
�G3��K�/��=���B����K��7 G#x�pS�WA��!p wb48s�C���{�5�S��� h�`�:�n�U�3�S}E��(��[W91�J��2�����b���E,7gUn����
SvX��g�;�:��w�E��u%�*�b�(���}�y��r����
�Z�<)Y��Vv;4�%�a ef��u|;�GcxU�%v3*(x�����͖�<J�Ζ͞u�s9�d;�&)U)(���A��oI���F{H#5
�&'�/_��l��:��:C��+s�n\�tˑ�;�fg����z���.�J$�q����EB$@}��_/���T�Ti
����w"�h'�6Ar����.׾\����.��������v�y��S��¼��1�gPw�k=�6Mr
���k��8ȍ	���a�`���1PJ�0��5I��)���jz}���(Ă�G3x��1�d���G�7UP��K u�`��C���4��S����)I^��*�7P}3gLD��N����r(�������Q�|Y1�D�8;v� Xȵ�k�C���\dЅQr�a�r5�q@oB�"��#���s�kJ�J�����8��]/���F�4a�ᯤ��1Y5���a�� b��,vj� 
���p�r��ޜ�;8���+�t?Uf�ѷ[��aw�A����t:�s8��m����TcCn4=4���sBB®�������cK���4U�c��'3}Nf�[G� �h�Si��๛�%�j��s椽��9�B��f+ف�����5��z�1<�=�]&Ɂ�kd�Sh�+z�o�X�'%��'�
�o+��ю�jU�>�#���US&�l�7�B�'q���a��hz6�Z�#ùJO�?,u
��Ȯ���c!�a]]Qss<����]�����Yxn�3����	|���YVyO��4�d�ZH��n�@������9��BO�'-�4C�B9ʷ�3�i��q�2N��U��&{�]�����T< T\�ы�l���p��F2!�Kf�0���L4[�k^N���.{�7G"���9�:�ЁtN��A:�ٰz!�[,$�_�E�G�y<T�\Y�ӔM`y���h��bS�Lu�+�����GC���exݪ(f#��ţV�c(�w�!�Xx�t�T�2$TY�a�q͉���ؘ��մoL1�SL�t<��T�[�I��P���h���r �@G_� uCx,�NH����7/(�J�)̨�O�nfrG�$�nWG��aTw'�C�@4r$��I'"!9eN��`�u�	��бv)�r�k�fp�&N�J�o3>��0���EN��|Q��:QG'�/�͍�����_P�bDDɰ���CD�OdV�P�d�&�*sc�<�����u6g��l�4!2���9���;z����yt��ޡe�l*�9�'r%i���pȊ��}`7���n��d���O.��Z�9�9���y^ⶮ��ɀ:O��ي��¸80:��B1�ݧpÅ;P�_ͪ�8T�9E��v�[{KGX5��n�����#���B^�#���@�{(��(�՚�hsY8F�>�.��c쿤R����B����U-W9������I�N'(�O5:���?b(q.1�3ݮ�D�xe��w�l���A��/ڸ���;�� �sp{il��P����	����_'o�k�c�"}�i�CE�����bIC�ޜB9w$m����s<�e�øݪf��	���uad��p��e"ю��c5LU�Oc�506�5k:��Eĩ:�x
:ܝ��EBʩ�;������{M�/�;/���Ws��%���8SF�8�F�9 o_�N�A0�Vy��	,�Ό5^��h湭��1����w:��3��)6�ݼ�23Q���%3�c:Xs�c��[p{~����TX�u����\h��)R�'ԁ�@�P�#!�f�@�#���Em<.��A"�*��+ӛ��%���E �7���5&�&wQo�!��(��U>ۀ�ӫ5Tu�ڦJz]MY��)���ڷ1w{��#t%X��ŮOg�����h��%㼎,��b���Q�>z��-wgr�qz���n��� �OyT��&��q���I��y3	�����;u�L S���#�Q�Ip�L�A��!Β姗��X��U�����9��wN|xRb~�o����rJ���$�s q��v]�P�/9mO^�J��G�Nj#΍m��_+��һ�����Ɍ����*�e�7b�k�5�N$���9���fdeFW,l�`#������2�����[���f����A��A�׶���Whl�G�䥏�:���J�^��<�����nw$�nÕ:滘�r{B5��|x�^T�݁���#�JK��X���������#��cy)	j�oK�� O���&�)�8�5pt�ZdbR�V��|V,�E���x�C{��7vN��K��|A�b�p�鞫fO P�Gw>n��WTS���$f��d�h"��+����|rp#�#cN�J���\렌_O;�W:`��E��;MBx��ڹ� }K��3���<l�B;�z`9�
*���%}�<�G]R�Lt�r��5/�w�[Z@t���ꁽ��ns��l��\^�\m{�5����I[+���nē�m��ޒ�O��(]�� 닩Y�Z��Y�֩P��B�5���V�Rq�����P���+�|�����O"d󢲥-6�bpm����S�����1�d1f�W��[}���z�gtK�ª�K�x_K�y��Vn[t<��c�c�����V[�i��ۭ�)D��Jj�t"Y�ܯV����E�Fb�j����z���k��{=m�r��x����yF�~��s(u�5;�{M댈VZX��睘Ȍw�]��G��ys�[�T�-,�x3ܝи�E`���I�r�ᬰ;"��c8	v��0��`��.�#�yn(��6��'w[j:��&�+�	��[Z��R�9��[���,�#m�S�J�I{th�5���K��J�Hݠ���Wj;a���O��ױ�m=�l�ت|�W.룇^:���\�e.s�;qnܙ�BwZ
��\r�M�F{�zr*�`[�܇/�a6�"����}�G���z���H�8!���i��+(p�4��UQ����99��o�ƚ�G��.K���	�qr0X�����7]'}g��e_Sn��[�ށ�'se�\,������yt����C�WAՉ՘�}���ª���9dj�������4+U.O]�7���hŭ����5�u�a0�=��l�f���t^l2�U��a�BD��CfW]�ۧ��S;{Zcku�iҒf�]�L�gK��D���fNT�ՀZ�cWr���{֞��jt7�Sv�{�Sב :�E,��C�~�
ퟱ':^�W�6uQ<��kNN]�wU�����k1��i�K�\~�Xx�vwZ{K-����0]�Y��nX����KVP+4�9�HDw�����|�����墷F�P�<��ժ�*�2��;L�Z�p ��R�n>Ѡ�ӟ[�iḿ�e�{�:Wp�8T�M�aU�2.��>ԭ2+�����Ae�l��z�!�^}���\�}'b�$�������|�L����=�Ə91l ��8��j�ar��A��4��<v�>�Z����(3J^��U����
���Dz�C0��%�-����o�O+h�(�X,w��,Ѳ:�-M�=��V�K��=N�+��F	~�,@�/ΠB����;�,�»t�G�wK�f�yv��1Dv9`@h�����Թ�-�j_i�뵴[��w}r��˦�٥K�G�����y\�ж��,�ظn���vJ��֣�����!�xr��꽽�F��'��]�n�S����-�ܴ�M�2�j�_M�7����5:�h��9�����i��-+H��	r0sGf��g�1�tl&ݘ�Y�(Ր�;��Ģ�ކg��l����U!���=
�S�JB��͵j�l;�l��Q9��Ɗ�A���;Ԏ��C�\����۶�F��8/yV1�b�s�Ss6�������=�U���lOĕY+m���-YR�e��-+ic���R�b*("�²4��Z7.*������b�Eb�E�e�"ōJ��A-�1h�X��"��IUP�R(ԭ��1�s."��("�ъ����-�j�*�E���US�Y��QDGm��#-�*
�EQ��UKj�k��3(փZV�lPAX��,�U�c+�&.R�Z��1Y�X��cKm�X�KA�6�[��\R1[B���bU�m�EJ-�TPkEU��Q�F �1UEV�,�Ek(�(�k(��2+iQ*�"���Z�"���
[Vڭ��iQQQU-*�Z*�H�F�QVe��DV����?�
T3o4.X{urt廓2rz��
�[]d�e!���<�8.р�t�G#K$C���:Q[o �\@`e��1��oeo�UU}����>	=�����H�5r����tkB��:�|kx�pBG�]BxU4X��P�賡���{����с�yK�dC,eDJ�����ͅ!T��>��)Wxy����:h�U;�8�&��6s���Hq�����BD�۟k�4T7uM�UT ��:1R��c�N����ە�y��`��SE��Tr5����Jv��nH�������L�N�W�uL6r��&�_-�WQ69��T�1p!�w�I���wҙ�.cDp�nF��FfI`�R���%:��8`}����b�NTa~�0� �Y��gk�5���\#8]f�[�j�=[\s�@e*��eWS�O��&U#�z|��!�5t�] j�du�ҳp�'�'O��7E��RS�-,�A��1`:�� �~i��ne����孏�����f�}0UץE�Si���O��Ȇ*����
,@	�xŒ�������B��W)z*zL��̦eN�]�3�p�R�C+V�G��1��x�LFۻ��Q��0�\L���
���ǊH"��h�	�9���;3^�Ko{k|>y<)���+�hpSͺ�]���cǬB�uW>tꑨW'���W!���z�gKs3�mv�����������ۺ�h��3��7�Ma�7�g^S�f�o�p%5�v�,��������T*��Њ�>��Nƞg����=��;u|�'�f8�~n�ِ���YM��W�)��*W�LX2�)�������ٗ�g����l��O��|p�y�l�܌�]+gg��7Ԇ�l׸�vH�^ܪU�/�vxKJ�a� g^�����t�IC���{���ʳ�S�d�������Adr��U�)�1b4�L���}s8��ۿ�=��p�o��㜓��4�pRF�I��U�q)���>]'�%{�������>�����:�0�e������:��v�U�j���/���˔4?�����f�m��	��΁�y�����>�A�"��_�J���F����#�I����6s��8��i�9E��N��nKͯmX��3V�,������ŭ�:�S�D���a��I��?`���c�um�#k&��<4u��1���C�3Y��l�g��S]�-���_�_5Y�˭�xq^e��u���r*�.�ǉ��������D'<��'���+���um%#�R�ݮ����(�˓�=9N��n��{�yn{�& ���U�ӫ-�� �Ҝje�Q+n��&5�#q������(�o;�vv˘��%��o��7Φ�:Lw�yؐG+$���!�S����%	B\ܨtf"{Nݞ�i��G��W?/�}�DB䲏h�����:=<��\�(��@UD��2�p��W��i�*ޛ��i�j������ہ�.�����4D��1m�[9�:� ���E_{E��z��Z�|:���8�LL:�B��G��`GU&�ۂ۷��n���'�0i�v
>�7'_%K8jyF�.uq��H�
�+�g��cL�wm&rܿ��b�����UC]�Q3%���o�{{��}Zh���i�mpw3
��Ddb���w>u�#o�]��7�Z�l��0z�-7����+x+Mh�j�\>��
���^s�F�On��7O�[V�sQ2Wt�ᾤ _M�P�/��`V�ؒ�����Cb�yc2ǐYB�,C��ѷu��"HN;^X��J�ų���s��c_��7�L��fG����E�����W����
5e��l)1���Gx��a�5��:��y�F.���\��G������*��]W7�p��a��l�f�XpVy9L��w1��ul�78'�b�{uc���ܔ�����[ۮD�AӮY��Z(�{�wN�Hsݽ΄����;z�w�v*Iy\F�j�])ZoX9�]IR�!n�*�R�Cy�p����{�i\y��Jh�J�K.7�1hz�b�Z8�\�W{�w�R�%�Z���t�n��%v���j��L���U_W�DjKu��#��08�� N���`/���2֎�$c�T���J�`�o �q�|�p�90�n+u�Z��'��@����}����&T����$Ov5]4]gk�����׋����m������Oq܂�)��c>��n>H����0�<�aω����#(�mJ�j���p���ܠE[�C�h����G�[��w���݆ʱͦy��gb�W��#�8^��k��qV�3���u��R*�����(p��Lnw��ٿ�%�J�BA8:>�=�����,4��>j�.u����yd���8r�sA��=�� ��3	���"����a��sc���U��S�ω�K[�U��)�io9ۘ	�tI���%i"8a����T`Ur�ɯ����}�P�\�!���L����:�Wd)��X���vQ*����G��X��7t5�;�X
Drʕ%�*����|�G �cE�uEl��*{ΘA׺���y2R]�%,u��V�R�+}H��7mfW��rg����S� 2��OWV�\wmY����C
�֩�Z����#R��V�28����Q��m1d����){ռ�n�{W}s:�������9N�[Ovr�M4a5rgok�.Av�d��JŨ�Q���i(�mnQ�F���G��}�Nҝ������E�ټ�� X�Y4��ϫ�(�u�W��Au�4��<o��f��:*<o�]��O�J��J���c+�����/b;���¡��#�S�\G���{�ji�x�*�rS�IϪ��:GÜN�O�,򨳘�]}���`���+�c8ػ���+=�A�d��}���t�PV�t��9�U��į��5��k�:^���+�{����צ�����B�[�����J���`���bf{ޏ�3J&��K*�;�ʸS4&[�6�X�w�R�8�e���
xk蔫�1��@�ב?(��1|���<�o���W\�f�u�����	� �7:5�)��b��(���������A���E=��R�%�x��V�낍|/�~�.��|���'��2�`�ꠅ� 6bO!n���^�s�{����W1 "��C����֙\�Ư���4���������]���!y�e{�`�����*�Q11�牔a�\���0�TBN��2��Og�*(�bŌF�V����9.S��{W!���_"p�R��>�巋���v��;������ˣݏ��9y��vi��6/�as�FVp����)�:��J<��ou�]� �CPm���8+zԼ-Nwu���Ut*��V���b�5~���ﾈ�|�R��Ɓf�_���}�)9��&��;)G�:��ҧ��U|�3/�/�P��X�㛳$���/7��A�:�7��̤j�_:�����2���-WlWg����6Z{<޽BR��y��5��T��Z/��S�2!
��@>²�1��4$�%ˈ3c�|�(���I$���]���};���k�����s:Ȳ��'檡\�8o�C=j���檳��^֨��Ʉ.�k����҃�Θ��p�E����d����{W
X�Q�X�go���.D�
pÒ��FM�,M��⡮x 3�m�ا�Q�\xO9B|v�=3�~��,yZ�/$�4��fQ�^ث�_D��ZU����]��6�^�r�Ǯ�(q���K�UX� �yWAJ���l��ˋ��s��;���F�	��(tE��1o�Zn.�G9�q[�k��͈�����Se��c�^_�F�N����G唟ԥ�j�ܿ��ig���Jb���UG"�SW��=���c���h�.��/�2+8�v�g�<�-�c����3Py�k7Vk��S��d71�\��|�ގ�Kk��L��+�J��~7��w��͠����>����x���f��@�H�T��ր5o]eZ҃�9��I�6�0?�ޘ z����^wq9�6O�بW��!��ʄ?�W�}���Eԯ٫��}�e����=]P�TE�e\B��x�O�D,6s�v��P��V�
�R\i�H�rw0��� Wu�>~�:<�Pqphŭ�:���):H����2�y����o��h�r��>�ڜ��rP�0R4`���7�=�#eT1���y��ֶ(�[� �u}��S2+��O��;�;�F<�#��C���5H��DI�, .1y HV��]
[J�j�d���2%���@��w�+{�}r�L�u��/��&��82����u7'vs�h���7n���86ڶBroA�p ���,��9" �7�H�.فi?{3Ґ��G�}z�`WTZS+��Z��7��\�B�I畕���΀e8|���5���fX��^Oʍ�6P�2��Pw�c{��|�b^lT����b�t�آ�i����RiG0�@f�K���Aٌ���1N���MX�l�ׇ�T�lފ5±�t�>�T`��O��V*�=��S|�֋+u���<*��ꯐᏺ+��I�
�
L�K��Q}ɾ�f.��+��	�36ɘ$�te�3���}��q�
.�lku�FP;����:���jt���[N�!
VI����!'��̙�%���� ��s�N}�����	�S)n�2w5w>�@�oj�k�ڱ���J�X-����t��Sp�oD���#��Z5��c�*�,R�!��BC�_=��ED-�X/�Na�#�}��7��lW?6uA[z�]��R��]Z�4imH��O�Z;��{Z�c��_ΤE�K��^ݩ�)�]�Nzbw����Z�A+��Ř�k�p9������a������4SޣǗ$͞0P:��e�:�,p6���&��;�&Q�-j��2��i�e#�&8b�u���ԸN:B��h�#Nz� ��� +Β���9kG
,���u�/����%���.�V�ЙcJg՚�L^S�鶫�gQ�p�6S��1�I�g�[���}r�j��=݇�f.�7X(>���Y����;Wf��JwD��޳L�Y�B���l�
��cf��	��j
o.8H�N��7ԁ�@�L�2+�雅��ch�$2�˓���G��q����M� '�p���zѸ�}P����:@�wR+���:�k�o/q]��o���ĩ�93�x���1_TC}P�f�rfr۹-�^�>`p�ķ2��+l���5s4:���3�&�W*�TƏ��#�5fR��1F�y��U�:��eP3��cK�0"v�3$uePq���Q��MWg���T��}ڲ�z�P��
�ٵ�9 �bO���� >�q�{�f�����.&鈨�$u�C��]��?�u���b�zq�YRj������zq���t�������g�P>�I���{�Z1�n�e��Ϊ/F����vw%�U�e�9�RPc�l�jD�ֲ�hT�#=��J�g�h$WJY^c�@*G
�~�#�I<�6%��� T>�D�R[�#_Ѯ��W?*��Y�5�k����n�3������.�n��x��S�J���=뻣��/֡8�:xR���fnz4t�L��1��Е`�.rte�V�,-T�i��jK���.�9�1����MgdR;t�W$�9��VPq�$,7��TN�KK<�,�8�9�����������:V��h�o��غxm�
Nz��ΙB����r����}xpwm��ƴtZ��=��۾;�)�:�y؍"f���#I�0�=���~�F�!^ө��*k4����_܎��3�OJ�/�
ٍ�ʐA�L���z%i��Ү�+9�F6�HU5LF����w�+���*�|��U�����w�kw�n����}������>J����G���#���Ի�>3�ۛ�ROr��TT��c;��9�����N*΅����B��c��k�Q{�v�=�nhJ>ٕ(�.�>��hcb���Mܽo��D������ꪲ���#a�<���#�^�?!of@N����K�Ց���CvJ* ]2�k��LeC���y�ޠ�����,+�ŵ��_t����М���c��O-]�a�\�K5�7��d�#X sٹ��T\ĉ*_�:�oݴ��g[����L�1�8u-zk�
�I������)�Yr*�S��6�&9��9���1��ʄ���)�rM憖M�
�^�T����6w��ʫ_��):���&��;c��Ҫ}��_/˾�M,�E�d����w�G����t�=�R5�y�:�U��zK�r(�[l}�˼�����$�C�`�	uٿ>�4\r�L\#"�� � ��@� 4	�J��͘حNqB���rS�Bx�}�
���|o�h�1YP���Y��s����_��ݻ\n=lN6AL��w��U��ƣEz&t<7a���V\d�lQ��=����*���G�ϒ��oA��']$�V�tA����(�E�(p�f�	Zb��!�R�p+�W��x^mKY��\+T���z����7�X�:�bffu% �wV�
��k0�*���]��{�mH�a��-�vb5c��8^�{����p1�?���`n��]a� �6�@:�]����E,� oCGgPk\%������6i�U�Vj��H�n9I���Sem��{�Ԏ��!���=D!�������[v�vL=�K6-h{��a}�j�:�9��oi��Ym:�o_fG����3��ʼ�CI���8<�6F_L	Ӧ�;G�l� ]�t��wb���#�+�Z�]M��t���*�g
��!���Q�G�X�r(�87���QҀ�k�v,�\�#痯�K*��[�(�cӛ�Ԃ�9d+a����5���R7KZ��RX��$6�ss�6D�yV�O��J<���u�g#goČ����n���;v���5�{M�Q��n=�$W1UbC�3a��S����
�h�Z��J\���Ыǣ�\��KFP��e�HY1en��,@�Tn�\�qa�w5�	�r��J�
�����vp���V7�W�fQ诟���C��{�fV�U2�}�h$���c�ĝ����萢�<w��I=j!�K���9I8>2�xv���"���ֶ��S=O12��5��q%�)�T�H¬Y��u��<���\��V��ˏ��z-۔<!�g�)}��G�g%��Z1p�ND��yۉ����$�'4;r�&h�=j��ӫ�M͂���Ժ�e�c P�һ��e�HV��#��;Y\rͱW�2?���`��w^9>����]�=��h6c�g��ǝY���v��VB�;W��9�����I.+YCoT���:�ɔ;�v�gM��P��G@�u聫�E;��.�����Ss3ȏy�Uͷ<::�nᶳ�`�	"Q@��`�jv2a��J��=�)k�]��<Zآ�2�8�Z�,�Md6�}��nvm^��˖�o��v���7iN��:�ٚթ+qӗ��:;���K�5�U�uq�귦捉t�Ӹ �뺏&[���������ٻn@]�m�2����vuإ�Li��E��
��v��^����+]��亇_��ΙC��w��Պd���1,����{E��W�+�G�b�3�h���R0��&����AZEn��1s��T��=��U��1б�-p���O��ї�)�|j۔�{wk�k:r�K	���R���p�t�rZ�k�nL8�t�ڊP�&�[��(�+���R���bj�4r����CN�T�<j�ԩD��a����v/�#�'2�p�>�ne[�7/�A�'�ϟNO)�X�j��}�� �Ĳ�͵�������w�Wa��d�oT0f 33���A���������Z؂�E������J�QU��b��b1�TUU*�Qb"�i�YcZ��"���*#J�)����+-��UU���1Q�EF2�F1Il�*�(Ԡ�jF�cU-����*�ň��Z�*��iZ�EUX����Z����H�
�+V�F�Rڈ1Q*6�*���V��1AF�c-,b"��(�PR"+Th�P��TEc+J��,U�J�ZQ�AE�m�1E��1��j��E-B�
ʨ�X�HQe�PDT�j��ŋb�%j"-���`��b�Tb�
���TUc㛩D�-zΞ�2�N�vg1��n����y�փ=�wh�	C��Md���ˆJ&R1�9_8nͤ��q�r�f_Wﾏ��>�(�u�m��D�8�U�m�\���1[�Av��u�+�U�:�RɆ*"*۷Gij�d���ѥv1�T�Wҙ��s�m����nxԻ��LVZU�5������(H̃]�a�rej��U|�>8ˎ�k�Dkun;�:�]���ö	��IA)��7����CU;����8U�d�EZ۸L�Jj������})��,1үo��#2� 7��ۏ�ݥs2��7E4����"��ƾI��ςt��!�ӌ�T:�=y��<��=\�HS�Tw���S��(@��)�di��������F/�V����(+�ևo`�}WQ���b�g|:Q�P{�;�~ ��:6L�u������9�^�f�;���^����ok���#��9f"iJ&:�A\v����r����R��ø�Gd,��Q��k��t��q��TqXX+!;�eTXρf�%i�@Z`H�=q0�\�<�f2�ng�%�^W�.l��҂a�QɊ�p�U���8!@�o�;Ȋ�ڨ��ZI�4e��sHw��Cˏ�Ɉ���Ot�m��q���hKb��0uqWx��o�z�1��Y��t�����\�s���D�⓰�R�ڰP�����>X�-y�V
�w�����"�G����K)����MoF,J��}GC��)�����jKu�.�Ƒ:]m��_W���q#��������~Az�U�d�Z]�JcEv*6�;6m��r]�%����|uT�v�]ڰ!���^�#E
u^W��36P�3�Pm�����b�w$�M`�=Ro��t�>��+��mY�E��{M:�k���<���N�_]�1�z��w\�2dGS�`�k����R����᫳m�3�Q�����P[�n�A�<*�@<�ʺЯ�]�e�RS��L ķ$k{H@����>���(.���1�����v����edU[��M�DE����@��uH�~�� 5r�<js2�����_9y�l�������Տ�up�����!ЎK����뿫�1��MˁȐ���rv��0�g��Z��H���Ȫ�ΐ��ׂ�ƸR�'��L	��p�&Q��L���.!9L�n�#o�b��
�2�;)3<p�ߪ��k�K�!v c˺d�$�9=��Y3!�4��|�36;��|���0+�ApF{��o��Pخ��s#�M���ф�o�\�s㷹X��
���Np����b`vc
�'@`��!Q��x.�9����-U7�blg�
�C!�1;s�Y~�ۆ�;�R���4z�e�ie�V��e�O��X2��W�PIh�k��q��-{Z9x�z�K</Q�Q_{־��b}��}��Ѻ�a��XD{�n��q	��쎹�;�X%;y�}��}P>H�n�t���m�ث�׏�KC��Ou��]9�������,��"�S���"b�����dT7L�,3�Soa��e������-��W1��١Em<9JGu	�����)��dk��yC������nx�`�,�ɧ/��0������$�?���,Փ�G0�=��b������.q'�ք"b�I��wc���2�ﻮ ���2�GO"9��?/�����\2`տ4��d�-o�I�;�e{�3��?j���%��y�h֌uI����C����c��C�m�C�Ź�}^urP�mLSN�����w�H"�=��@�=��"+�_mn��j|��]8�Z6�Qq�t��� O�҃Ψ�����E	X��\�6J㇛��+k��]��X.'��]��^L`����ʹ b�s}������K�3
��&_N��� ���f�r��� �X\䱗[p�%���1���gk�K����u����[1P�<I1��l[�=��%X�F$�1��S{�@����y�u6]�S$�P�u�j��A7v��l��W�Q����2W�זb���k���uG�Z+k��[t�b���v�f+�WrT�̕�h�'��W|�s�o~�����W	I݉`�����>�5�)�EI��氫�v�\Ƣ�:�쿗s��3�@�7	u`��YO�_�������~�:�[X~b�N.P�7�(�Ã�_y,kG_R�r��-���=�-�6_�5MߞSF��\c.�,�q�c����@Q� ��9z�Ê�׆H.��&���:�fu��r��<w;��p%�Ж�q���|��/O*�Y���
��e���p�V���N��������L �n�*�:R��=F/V^f��-{�t4֯�����mA����䜤m�!�nDأ�ղ`V͹F���ǺԅrJ�@��&�

�bD�/�\C���m&m�w�����۷fmŧͬ3��}�P*0F�{����e���8V��J�Ϊ=%�Xϋ���ǵ{��Z�jzB�^���t�T��U2ᘎ�	���"���i���u��ک�>NxOt�W;���j��-8F����B0RN�����"LX�_�1\̾:jauvEpd*��x�n�<�P3yS;V���޵|+LǷ6��.�\���Jg(#��cg���NL)��zzqK�۫��P�l���aw�6���랸*��:ҥ�}݃�{]�Nnt�f\Wo��y�=v�:��K��^T��a��������.U��f�-s'����:I��}}���V�-ʬ�~��OI��e�s�ō�b��2!���VA�P��E k��A��Z�������Vz��C��ۃɽ�?'����|���g$}j��Qd\`n��^wSs\�w9�ͽ�KyՑ�?q�/�>	�g����읭��({�rzb7��;��M8қ���B���_j'��K};��q���E�o�ʴ�k���W�g���2VPʗ�I]�,Ե��\��t&9	��k�Y�'Lp,��P��E��ZU��J
;=퇙��X�{c'cPd�5�]�e�R�ū�i��ۭ��ƥ]��eR5cJ������Hm\����'���[p����j��[�Ꭵq*��ފ��A阡��aߴ�������\֎����|�j�H�U�۸L�Қ��k/k(hq+��.�H���yNMi�Z�ӱք��sR�:��`tR�b3"��$g�T5:l��is{�Ҫ��<l͸��V��eVZ󝢊� ,�{���`q�B���5+���h��35�:�ix��	�4*�\�:].A�I��us�n�L�/
�Y�v]����j+�w�ы���0.ql�VR��A7�TƭQ�D�j�h��M;�%H�9b+������mZ�y ۥŻ���;�آ"��wܐ��hm
Q�������}���7y��v���R�1�L*L��X���K��@�+��=&A:�ٰz���V
،�uE�{o*賔9���Σá=�*u�5��~�����
=�'ʕo�|MO/^��_;�m����{ì�xb�2������X���z�n�qs"EE�f8@�T�������c����=������q���0�n�b�gɪ�7H�
 ��Q-ĘS=�aO`�BnȀ�1��+���l��X�Ua�>fw*��y_F�f�j@|K4&�v��%M�b�w����|�
�&a�D���X�(!�y_+�bw�4��wJ����	ضz$���}IE�FJ(񶪡���N�@s8�i�mp𫇲���:�^b>v>Ӡ���o#F|�u���#��-��{"�S|ᔍh��\ ��Pd��^x˙��_����V-|t>�"Vwl��13ݓ�^`9gbJ�՝�]�����|����F*ϐqxB����-��]�/�"l!|US���q�n����u<��AK��8""����f1Jm�߁V��![�<��f�ٲ������#��G_#�`��R��[Z�x*���v�th�7dj��V	{5���T������AX�Y��f�1������\�M7l�0/�UU}�9]Z�x�oH�d)��XU�����.���Y�����L0�ΈZl��G9[;ui,��:��� H�X�v��@^����(��a3q<��Ϡ7t����"r��3��p�c�9��U��'��2��y��Id�z��m��[���+����p97����~��[Y�eC�2oT�;�E[�J��S�� �#�Ϡ>"�8����4����LD'M�e|��6+�7�S/|�ޚ=˺�{�rT��2e)}�ޠ�e�(�Y[}U�t�2�9�4�
�����F��]�]��>������֎���9\0`�$���x�I&/�pevQ��+���[�p��+;���{NF��t��{��Ykz5Ye�RU+�J��r�'�c���*\��A�b��k2�;����S9�\g1T���^�˳S���:*)v�1���d^��N{g�[Bf�`�,�e(�D��.�|A��C�S%ˤ0IZ����t��{��t6���?(�a[�_67{�0�0�G��:�WJ�U׸�e���O�ޓ\���U�u��4�h���;H��;oW'�V��꯾����{S�� �:���������hQ��osA�ˊ($����":Bj�'�֭~�q;���[����5�+X�:.���{�1Tݣ��-��~ߊĻ�j��[�}�+�3�y��]V�����wZ#k��%��K;��Lk�{~����G�^�.o˖�ˮ?K��"�O3�8fm/ ��m-��{��Gi�AuN?P~Ԩ���ØO�z���T�U9�5^<��紽߉�ꂬmD�1Z�E�N��U:6{�-�鎱���ө���e��ks�o�
�ʿ��Րx=�Te�̒��]+F�`���P�sC��p[�z[ˇ�n�&�%h���+n!B�]F�I�ču�O��t������
�k��只Դ�>ʷ0�'�ṉ�zM���=WKy�X3��7_�9H��R��k�\-?+���=!��\���kѵ�z���qݩ��\�k��P
�v�V�n�+��2���y���P�:�7L��:��Ȣ�y��7��4/yb���nE����ɝ0Y��5�gv���������^;58����yX�V(�s��U��mL�˩�$ﰅ���gu��[�����+y�M�f��"|��i�e\KD%�3/�	�����G�0���D��Jc;����.s�B9Ü$ꊮ�0�f��?W+^\@}���M��y9W�̞q��_�z��8��/#��I�WeD[Ql_oU&��̓�X�b���ݐ��QU�;��ꆬ��/@0��,et�v�l�����sA���g���z�n��Ŏis��A�9	�z
�v�����S{��쮜�j&�ǭ	e�Z���:���_^=�Z�z���i��1�>%7.j۵�ֱWu��{��n�������\Υ�����
��S"�5a={��AŁ���{{4���7(�ʃ���lb�ԼӮ֪�ΈŷO3�8��y��J�����ڞ}�7cep̢��ģ�ƲQ�	ݽ���r�����Kޝ�R�z��������ߐ���hq��u��a�C����ސ7�W��St��c����={�G1#zd'�$Λ�%y���h��[{���am[����W;���58�vE��K�{&5�!�]e;xg��¶^����xV2o����Z���V���`� mζL�P��|����J,-��G�f7e���F��um%���hST}ˣ��5U���"����w}.k�Ǉ�\I�[:�^�O�Av��N�c��[I�|�|5�{˵S}J���-�x����2k��l�m|���r5Ԩ2��T%�)>k᯺��Xmg{<�1å�G�e���/xհ�]!F�}.d%��W�G+�{rb����:�jd����r�q��:JٶU�J~��阁ϬP�J��)��.�v��V�t����o[���|8��>�"2�{8Cu���J�x��`�kQ�%������ՙ�������x�\7���yfiK<!+�gz��M�c�l�%�\S�B�ٲ�g5�K�ܾ.�w����P�%��qj�������X�H��&׆��}x:~��~Ŏk�厷���u����V�w���u�=.��&c���K�/1^3����Nk�ɹd�'����-�Y	�gE��k�8�9���wr�)7�Gô�#&9uf�vKc��U�,rkGf͇���Pֻ��m��.y
��6���CI`ŵ��L��ZPY�*í˅.fZ����,�E[Ou/B�o^^y�ލ��@�x	���	ǂbHXrX��& ��犳uT��H.ӻū�N�&��-��n�>5l*S%��t'x�=�oӣ��i(�����H�sȓ��l{G�H�ҾH�gq��j&t�]g+Nmws�9�tܫ��p�f�%
U/���!���&��,����冗-�9��ż�a8��	N����2�Fv���`.�x�&�-[9�M 
��.M���`�X�i���2d7H�fE�v�o�z@և�V���L�^iu)I��t�j�q(Fn䵴J���6�ԄC��Ŷ�;�i�����c�����x�8F]�p�v��W z��Ci�1S��+'���M,���	]׊%�EU���1�^��[,=p����f3��إ���!�h6�ʋ�(Cx�w�u�ބ������>ú1�T/͖����ȏ�M��>zox����¥��h�k�����Jl��V�Dm�n����Co��O>^��Vu~սg|E0�QM��z��vq|��	�7�)�o!�y85.8ݗһ�V}ˤĆ#x�T��J���}H��X�lٺ�"��!������kXf���Nіt��ڃ
B1�1_e�f��{���'��fZ՜s�v��N���%��` q��c���;2��iOa�*g7��A}��#�m�ݺ�乪˙Zsv�-�93C����)|��eG4M�!&������MO���<��N�u��'5�:ev�z�]��^f� e��_XkuM���,o:��#��[Yx�-lR;�dAs�	��ʒbv�RDr	�D�<zo�C�z�|1�W��K�\dJMzo���e������m ������|��q#e��6/rF`"��b�%Mٗ2B��-��0��IZ�E3XW�R��{)�V>�-���^�Ц�X�ҏ?�]0k![���z��ޱ�������Uvk�׆���'�؛�\��[ws@yȽӇHvQ�f�h�Z<e�꘽��X�:0�ʰ3z���u6����B����Wb,�I�ј�����z`������)S�`ϩ3Z�:ح���N=㏬�y�*&\����n��uf�4�-=.F��ۧ��\���;]ɥHmZUm|�|e�㢷���OB�vk����r��l��\\Mk��B���X��u!�T��-�$cYX�%���6�f���0��+j�D\����=8�M��2����%�D�t]Lk�o7Vr�����G3i9�`r��n%L7���s�/8q�'B�b.>��4�s�f���:'+��]w����Z�Gc�}�6��Ȝ,���,Β�x�q�X*���go�n:���!�R�"�R;��o�y�:��@m)��L�{%�]v� �;[X$/F���a�'-u��*�d��|���q�4��9V�������Ͻ�H"�WV�+U�R�YT��ET�"�UF"�"�X��+UTX���",U����,2�TR(��(� ""
E�ZT�D�*��
��`�"���`����ʬX�J��U���"�b ���
��*"*�k
�Ec*��b�U-��B�lQň,b�DAEDej��"��U ��F-h���U*VE+���"�
�@Ub*��J��X���"�X*��EEE��Q�TD�TR(*���b�E�b#�QTb*��YQVE��`�
�°U��,PX, bE�(��	hJ�EV*"�X*�Q����Pb*��-�Eb��� P�Q5Yٙ2�Tv^nk�]ؕ,�z������nn�S���<�*��R~���Y&�{3G��b���P��+4]*�)���Y�7m�z��Do�D���]#���EvTN���Qy9kbX][�gR�{�W"���i�j��q��K۩���F��^V����vs��M�ZA֐{{~�>O`�Eꕯ'_q���O�6k��%6�cE;��%��橶�.Ô��Ψ��Q�����Ԃ����.�j�P2�=ˌ*��Yب��U�u���c]�������V�9���7��5��}p#"�b�MN&3w�H{�p��W��	}-����v��~����S{4�p1d��R!�S���i���70UjՁod�;��Q;�W$n��e�����M'���=ܒc�ǡnt6��
���amB�1��D��{{Re)�4�\�G�?��{��?B��MSK>l%��7�)�e\�˫�}p��Oi�W��7G.���l�����.v�wD+�_wC{�^8���)�����wWn3O�$�c���Bs��w#G��p�wj���+�k�R�U��`�U�.���B��އqei]j�w2�`,��c���t�qR��UȰ�L�/��QH{���/��n��CKw�����:���E��t��{I�}�# ��� �����7��9ǔ�])�꯾����o�]�g�9�	�Y�t�Z�]���q����'�������϶����tl�w_2� ��'1\%n^|��RcTqW E�q��nˬ�H�jp;9��:�n�~��
���+i���g=1�u���GU<���S<�o;&�S�l7pr:�?6�e��Piu嫻�pc4���le�X��X\BZ��IQ|�Zڃ�e4(��|]A[���8'��V<�w��=���/�k�koKz�O`m�����0�P��6��Zn�]�e�U�h��h�Z��mՕ�w��K{�Ԍ^o�OC�iV��G� Yꜭv�(q��\v�(}1���jz�E�_fZc�]^���@wЯw\b�#��N����RZZ8�����uN&�P靖d��J�%Ng.�i���N��:�A��A��<�_V�T�w��'`x�#T[�������W�l�ՖU%�K0�;�^\�q��my�E�^��hh���\�A5����4����V�֌�MV�+��d��]�t��;U�+E��|��W^;f��ű8��U�},�E�_Mǚ��+�֮���G�G�y���Ӟ��eO/Dt󺸌k)4�����V�!� ���t� ��֊�V`��nn�N]\�'��es�-󿴷��-�M�|�8�[U6x�U�-��O��� (�=<�U�X�wG�޸I��m����;�B<�_uec�Vis�+����(�K�̄�_O\�q�vzG��5b��ϻ�����z ԟДd�;�-�WKh�U��'t:�>����k�V��/o<�P+d��8���*�yfb���6s�k��6�ƸX��_f�n\dk���y�����9�lZg����;3JY�pWn��g]���i^įU���n_�I��\�x+JM�9NP��,�E���"U�QU#� {ƚ��u��,sK9��TZ�!��
�4��e�K/��r�$=@+��*>4�}����k��v���\���T)#7
2�$�F����$G�����	���>���wxf_w#�d��Dg:W�/ּ��[�]8\f}�A.�ފS]�gJx�VU�{;l�j��yZ��k�Ddr��V�X��!qѩ޷�v�-�@��;ժ���p������[WX�$}�t�;_G�\A�ʃ������F/i��� �$TRQ����v.�uM�M��Gj���P��cr���.s���WTu�)�ʚU�������k婊��-�k��ߡn���PU��V���L��-붣rR�>r(<���f����w���{�^!�nG>Ue��t��y�Ҥ���gՉ����p�5���{��W���;b���w�>�ᗈlY��>�@p9wL�F.�<���a�>t5��k�i`ɚ�\�z�Wm]�N�K]|�����u*JL_%�(�$����7��F��n��&��k�c�q��.��a/�!��Y��
��X���֤Q���,o>�X�KrҸq�T[���X�9LJ{��U����y�PM��]��g+z�x�����Ծ+��j������tf�΃A���Feo<�{%=t�[:�3z;�mpз��S�<M�^��s~IV��we-;��jv����u�v����k�p�����'/��m�ۊ183��*}϶=�X���F�!��x��'}�mK(����+i��F�N9ՑBZ6�xi��;�>��\[�V��=蕯!u���K��V���
C�+��k׸{|J�O�;,�~��]sȦ����7����P�S��>�r�h�2JKxRJ�ȭ���2��^�w��Q����/��O�T��)[׼�;ؙU�Q��5/f�a��ήB�]�r'��c���K��^3���L���7i�O��d�;/��Wr�0w��;C��ʫI�h���Q=:�T�^���7��n�W�)���膻.��V��Ev)�v�{�a��r.�ִ�s����qob�E��5�\.ͨ}}5p)/"�
=-fG�q�T�7�!l�|qv���YԸ�����~�<ќ�y˒���n�n�y����NBi7��Q<���Uqѷ���M`��6 ��s<����3�b����O�����
��W�PkZ��<����P�}�7�2�T�&��=G%JgWr��.2,��#\.���u=v�
����ʖae��̼H� ��W�řf��\k�Y��9g�੫ɛkݎ�U澦�k�#��	�gt�)��"��ٹT����k��8NT.5ۻxmt�u�U\l����{G�|:7T=u�ks~	�\je���~+�/V���A郱��T��`��\�67}ݦ�T���o���e��.ۈm�AT��mB���č��e�� �yYN v����h�of����۝��i�uu���[LWkx�U3�Z����DOLs�����\;Z��WzM���4�K�P���l�UݻL'X�yL�0��5yJb�d-wave��:m)��5cRo$���rS��f֯G@�ڲ:��fiJ<,��	�p1Y�#}���׼����=����$��W�{CGk���ɐ�;"��}ᡞ���xr�{f����+ƽ�k�u�o,G-������I���>�*���P���h���.D����5k�qIsC�p�XDv�_jVZ㋛py"��%�
��K�YU�K��Ѩ�m*��W�k�zb��z��r���[��y�֞�3�N1,��u��A3������^v�&/rv����%K���f��%K��R���L�gzqV�-��:�rΊ��N�	Y��{����F�ͷ��jC������j�s�*l+����E9B�]�T��4������[�n����A��ffp+8؋�55������sG)�wDO��
�ʃ��b��A���}�j���������k"�pbԸ�Y�_.=�2��1V\�T[ꯣc\�0Is5�QZ��Vj�q��m_�D�����3W�{P�W�mVG1s��5dT�������z]�51��[�|�w���+k��[p�6��u|U���P.�c0�c����Z��N�r��T�cY&�܇o����>��E�z�X�z�K�=q�s��:�~�O.�������C�}��EJ��2F�z��	�N+q�J��p�L�65)p���h�o]�Jއ�گyݭ��e�g5Ft�j�f'�o����%06��2���O6��&�Eoq�p�!ӳpξ��'R���ɔ�}�1�q�e}�4�S]2밻.�m���4�9��1%.�w掶��1)���_�5��B������K�(�Y�d�)wa܄�̺W��Ɏ�۩H%�:Gu�8����ǁ�-�
��'��u�_+��'1���PϷ�GN�]��	.��G���ϳ��h-��Uن����Β�����wK8�w�_})�b�B�Uw�;9��ܩA*��{�� ��V�_N���v�������W�v���6n=�a��"�
���㶕�Q/:U��M�
opl�:����{�VW�Q�IӸC�9f2K��0��}{�ΰ��6,?�쯍-��UoL��4��}ج;���!��n�nT�oE8�Z�{Y��I�p��0�t^��ykb��m5��ɬI� �wQ`�^�E�}d�7�KwJ�X�����Y_wW�w��1{L74�fu%�d��V�w1]�-�N�pߜqx�i�_s�_`�Y��q���v����f�H�t�5ю���k�1V�;>�{�fo5oa�����ɼ^�8�IΒ7��O#߈]��^��]=��.�m>�K7��k�!�	�	@��2Z��rx3kk=�f�~�m�CJbߦ���[��U��&�a�w�ST���͔&��������Q���V9.����OO�~�R��tf��gx���k6�⫠�ݴ1̹�A8��u�*Ec"��MBz�zN�2������.�v������UQ��:�[���3�����=2Q�;�qv͓�L��񘞭�+~ݭ4;�֫�_c벫����*���(FtO|`�.�̓]�lh�TƵ��9γyfi���k��o?��W�r�FW���ڱ��O.�G.�p:~�Pe&*/���zt�"f�䎮�Xj�gJ�P�ݵ��w�	X����D��	p��ǌIq���x��d�'��r��i&���ܮ1�LS���W�l@����ee����\��\�f��Jִ�j3O�+��B�p��7]<T��P�Ю��S��ƅ\i��ݜ��)��ek�]w�qN�K��;�<C����	3c�&⃦�Ź�+�H��w�ݹ�1+rj�݅J90�#�WWugyC�R�^�Jqv�5�Lp��X%nE�駆c9��\8;�6��@��ƙ��9��MC�*]|-1�pWm�.s�(���٪��}�a@ɹݭ�mW>p{]���
����e(�ᗆ�[�-*՝��g0kf�7G9��!��n�;7��nK*�*�����6w�n���#��x`凱N�7�59+�C�X�)$�q�ddvɾ��3x,7(�+�طQf�&�hby�v�f�<+��s��5!9��;<�����VR2y��䎳�8�	��t��Lù�r��
��v��.'gHM	[������m�ힷ�lb�DWW�����qooTLE�Zc"ևRkoj�"nm�|3]W9sˠ��1�s�<���{����v�s;�띘��X��|���O$_O1}�p��D��W�md�U��`���N��R��*�k� �b�SkY���p���z�O�ے�	}-���ݤN�x�ȑY�rۚ��j+s_�:v1,��]���S�Y�d�%E�r�Ex���݄S��_P��]�)�'Πk쿖��pۍ��m�в�B���ʭ��ޚ�O���w�|�I��b��Z9S�\��>�F8�N��B�R�&`��yt�gJ�9��G\@�r6969�����K�/��/���pN�W�ZTc�O����MY��rʿ�5�a)������f\qM�����jm�B�������g`�=Up˜�C�3JQ�qv����V�Bwo� 
���̚	u}��5vnE����g����;ox�W�����҇X�0�}��T�ufoAI�oq�x�C��3�������N�dKdq�g���{U��FƬl�Ս�-ɷ�	��-����)s�*��,�rpt�W��f�F�/@�@s=��l�,���Fj��Q��U����wS��v���Gze�#N����	�'g:ԥ��S�qu�<W�w��E�tŭY�S���s�M�땾�K*�9l�gD�{�\(xw	���eM��y�.���q�Ώg=���\�4�L�l���h�KR�;��o��pP�d-�EJ�8��9��ӕ�� �"*���`�3KM_L�:�"�)�1\�M�t��õPQed2��~u/Y;W�w��2��*��C�f0((f�.�[���TAN)���r�Z޼z���b�`Dkq{(��Ϣ"t�y�E�=��}��p�=�m���Y�@�}�sY/t�\�͙ ��,ҕ0�`&NMw;WE>��i�O^3��jVE�`uֳg6�G�q�q1@t�]6�Z��=X;uԁD�*5�;�i���׉��C�	��j��E���_uY��"��jM����i)��nt�}���Q��]N�+Z� 7�l4�A�9*���k�[3�^��;����r��-���Cj}��{Jv'Nz��C0�X:n��Ud���()���v������B"஫�"�����/{�fgc���'Gن[�I
,k���j�+���k���Xz�v�x:V��p�)�Soy�뀨3)Z��F:-�kR��`�oi/"t*�,����l���Q �D��X(����e��ݹ[yKW����o]q���z,�;]�ɳ����~�G���M�:>/����NԞk5\�C�!n\�Q#ɵ�+�[���f��� �EO8շ}���_�|��Ov���K'd)N��
�l<)���-��ݝW�s����6ʻ��E�;����Q���oJ	�k7*�4���/+B.]�U���)GA����5t�bȦ�=�F;a�s��*�ټ�ESW
xd�;��k8�ŋ+�s`�]���]ܗǭZ��N�vA�0��l̐��&�k��w�և��[LG�i�:oRӍH�o.Z�\S���u���^V�6)� �p����7'v���N
��/N�B��˷�4$h	&v����1徰��nA#콊�Tq3����k٤!�ځ�QC�U��z��k�w.�ۤ�w���蘛4>{��ܝ��9����{o�f;=�1�W7xѳbn����1ϡ[j���Գ��G��i�[̨͜�����K��8]���m�ZʘB�pU���,��B�2�.D�/�E���DfCvI�!���6zav/S�d����x���}ٯ�
Ts�s?��DP-��DQ�b�����b��X1V#PDP��PX���X,��R+�Q"�,����E���$QB,Q ���X(PF��b0TD@X,��"DVIR��TQd"�R�"�,��"�(BV
VD`�(*�b��REP
�����l��"�"E�(�E��E���EdR��lkDX�X
�����B���Dc+RĂ ,P*+ ����X(E"��F����`�,DQ@P� �Q�-*J�$Q�(,�D`((,��@���0`�UAm��2,Ud��`�X�"�m�R������k��LY
��Z���]�ͷ*�U�Z�{���b�KD[?%�x>�1ͽ��ͺ%��ѳk�}p�u��a��vo*o�S&w�jcj5o>��)GW��LRc�[xim[	�p���Z���S�t���V��b9PĘ���>
���_o�vǶ�G�]@�A���7�셔�
IZ����3ڝBT]}�B������x�z��n3qro���Kb�}x����Aަ�5Hz.[���P}��&�6=s=�n(l�zپ�|>}�b�]�4���z�4����{�z��_�[�H���R�m+�����5Լ]����fy�y�g%�+C2c��ɡt��k���ǇkȞs8��=�2�dlJr�4���-��vuV_�6*-�ۊ�i;[�t]��z�̓qW�a>���u{�s�q����gU+����kM��V���>����(�'99I��҅���P\�D�N��������io.!�[�	�2v�����j4��f�ǬPv��|��O����o��j]�[�0^����&�;��w���_.����k�+h^���`��P}��X}�Ot^W�_��J�CW�ɋ��h��W��{K$��Tn'��tÈ�1(���u��Y/��Rr�Hh��c�Y�9]b�����P��'�:&��l�j�pdk����kn����ZB�/vz��S��.QB��<{���#���J��%;KGwB��ICj�N'6\d����W�%�)��p!-��%5�?����W����+v>�4��O��z�B/4,��:WÌb[��n�1�,�B�Q�랦���~��ڮ�]A�ɮ���;�g7^GW�٤Y��&����Y�&=�.Vz۞�������tSQ�����Y���i�7P[�0jo��A�n�Jƍ�� �0�A�ʃKo/�ޜX�b=�TG9	���2�nl�v3c�cy'Q��=�x�w��챓ȥ�W��>v3W{|�O'����L��U��]����ϥT��+��[Ax�������M7�c��Y�'��*�Qq���o[�\1����٦�eG;j�
�h���V��|3Z�Sn�%8s���`uu�7l�V��_U+�I�fT�ۜ!�n�nM��=��
�hb�i�3Vz-�-S�<��cy@���1�/J������B���S��=k#��)(��Ϟ�����鱡�ׄ_0!�]�*��a�}"��9�x�ZCI8�}F:\�:��қ�v�B�1uUz��/;?{�3������Ik!�#82I�[j�q�fR��?\㨳��8��u���Qm>�W�P���k�^.�I�s�=�I�;A�_Jss{h��@ㆩ�����}����g!�պ�V����g�o{ه|:j�܅P邻�Qs�TY�m'g�8y�+��fv����8Y����IvD;}EW+��W���&O�Y�*���gs]9�c����\�+N?��۾)��m�یkh���̮���-S����&�'ٻ4�.qia�o,����Τ�|;R�q�N��m�b��&� d�GZb�s_\�㪌兎�w�\�kN����֓�nj��f���ʷFY㗹=��J)���G,��"V��»wm�>�=N��:b��N'h����"a8���9����0�b�2�&�=�
�1�'�|xTv9�ɚ5��܁�˗g�g6��S��3oY�������x���95�Nw�yX
mm����S:��;R�ۡ�W�*;�;�l���D��!rܠ�]�]n^u���f�c�GSUر�4N�����t"yWubi1�Kj�t��8��^���wEf����N=4��,p�������w�w����GG�CziK�ʄ�/�7]f/+I���뾇	v���/ZJ��yu��8�޷�\a���{nGf���A��[�wt�9��m.���]Z�М��ڦ�M'�$'P�K!=J�s��F\~"��8�.'�Ҩ�[��^�:�b/�17���Y�;�v��f�"�T��ε�-�3>�<N�eAw�*��ؿm;�}���3���k<�,��:ߴr�}��:=^A�qh�ok'����!{~�9W]dreB�zhI��������~ƚ���mCV�^�� ���j"Tք�FH�z��;�n1�cy\Q�q���.1��M6��q�J�.:.��j�,t��T
���}NԨn�}i*YE�O���ޅ�m�����8�5�� ��%������oplr����WC��A\3W�q�6�f��sмX����2e`/�Z��j$(�&Y�a�+�B�Ԛy�нm�R�󝝕˭n@�$w��btnH�q�E`�Ι����5�"!��Ӷ	���峝:C�i�����j�x�1��9�$�z*5���ܱ��)i\8ו��pⲱ=��g�(���ٝ��j�c������ܙS�U��<�g3k�� �� �Դ�}۸���8��˖�<�CZ!,�+��ς�ˎ)���m������``�H�W[ݒ�Z���i$��
څ!ݚ�x�PV�Nb����e\�h��!VP|�F���lf��S��3e\u|��&8o�nT[|	��w�=BЩM�g)o�ь���U|r�vڨI����ayb�c�=�Vn�T5�Ge_(��w����]�|�򰪣�\�:�r6��CYOM�_Yηeor�yq�١t
yΰ���]|V�A���}x��^�[�7�뜄��łdV��w9���]�������-�����ڨ���X�w�ڢ���Z��C���j�}2K����n�Ky�2�~�V�Khq��ą7�̥�j�5��w�����c�Uu�n<z%��X���zt׽��x.��N��y-"+v�v�
��u��s]��M�����qž�}n��<��Ҍ������Q�MTV^�cm�ð�͵zA�Og2���N�={�Ԣ���WR�7�t�sZ�����H�M{[����a����s�;��G�c0*��.���ݨs�� �RT�4_Q���������r��'kK�~&��&��W�Lu�]O��d�&<s�a؛���w9\��V1���2����I]��Xs�W\Nu�c�a�x���{�Ը1;�7{݇�o9�iO��I�-+g�Y�x�r�z�̧��LXx�c]J���¢���Z:U�g�Հ)Լd���0�}r5�j���r}ʤ��ʑ�2r���;�wr����C\�Q܎���Ln��1�LSl*�BX�w'��b|��bP�ƫ��랹���K9+�u;�4sqk�Y�Q�[�"�T�F��}�������,>��W&�|Z�O�5�rtU��E)ʻ�4�l��;�{ś6<w��_c�v�u}�ۈ�)7�:w�}4z4�Teƌs��-&�Qjf���������xIy�{%�6i��|İ;�m��9R���ϋL�k�&�S�
��Iq�ci�S���n\�!tL-�s�k�ь�j��_	a����'}�tկ槟���R�oq�7���',����`�6��)͇;,3��D�9Z�f�àr�IB���xr�۩VLS
��o�
/���ڋ�귧9��k�����٧l!.2Y�&�`��'	(=MK���&������:���x�uh2#�V�-��u�#;�]�!C�y�+�X���,��TA�u~�?H����ĵ��+	�X�;X���ӽ�I�F�\�S���t���e|Z�۪ E���T�{��Z�i��|n�[�Q�����E�7�Pᙵ�5mv/v��˘8�u?4qN.sé��ۗs8��:�8����67�;����2��S����LcǦz�o��=&�h�;�3��.�4�j��yġ��20EF�.���t�'[�g��l^��3��Ρ�?v����y*7!�"˱��+34��s{��ɽ|���ԫ��;*��Ѭ���&	�\�$(�3�U��������M��Ҹ����5��wp%�Q���g@�]c��O�^��t�O��5�e��&E�b������
��{��[3x��������)�=x����*N�U�b��m�qf�l�y������=�n��<�vD��v]r�]�����ܙ�-jX����plK�o};��E�⭵+d�Μyw~����sjN1�sIBh$�N�9J��PURP���o]��넾��;��Ϯ��kZP�)�;��y���]�F���I�;��)�v`�šT@��Q9�p2���]�}қKz!��kf�}w�[�{{z�t��.{�G��[�s�B�����m.�fJ�����g�����)��W�B8Ԩn��Lp���Kj/O���su���]�+���=��\k[M�Φ�����
�����~4��q3�����'�bu����z�ϻ}�J����'�5�����u�XǮ�e��!m�Y����o�ү�1���F&�b��o�Nv��t�Tw-�Y<y��s�&\n��+�c��ު���QooTM�&-�\2-UR͢|�O�pל��CimFh5��9:�X��-�����S+Eѓ���M�%�u��4���!�u7���J���XԊ�UeWQ�4%&���i�`n�˜���rI3�	�qGmG��r�:���:�i�	Or�yz��IsF\|�3^w?B�)�ҵ��Hcj��!��~^��P�ok'���!z��J=�}�jV�U{���6�=s��6��kq�m5ku���W���S��ΎtM���ܵn�r�{I�r��ZM5���AJ��F�*����8=�-V�r��=F^�\�E�K$��i���Z���m�|z��1�B�ձ�y>޼%�S�wԦ��p�f65d�;�S��h�og~i�p�wmV�:�dWO�����z�\K���p�2�BS6�����kGt-�3����C��[g���af��p�J���E؆���S�t���.��F'e�ڙ��Ý<�[s_�í��*�Y��Hp�B}\.t�9y�
x�a�����ow�I�P�W7��L�y
�A��
���$ؗˣ
�ze�%�4Rq�Mvŏo�++����mC�*��@T>�2�]�u/l��x�P��¯��\#9��铈=�b�R��`��1Q�����XXЙ2�*�����Lf;��W΂�R1,��\���o
%�}{��<�Oz��̥랷B�in�e�E�c�e����S^��޶�P���y]�*<A�`���!oV���+�^�ݽ)�ȏ�h;��R�>b~ŀ�u�|�>�O��ޛxY��F�.:V55�Y��I�a�!V�Ps�^b�Ǻ���M�`p�6f	��#���}��W�HVo�������]��\t���X��w���2����f'ir��v�����s���V.c�fQG�Aqߎ)�����W�K��<F���,��wF:���lU�[��W��;�6��6�F��ɕ��>AN�(T�p綳$����\�Q���Ȅ��Y���;����\���yA���xw�nzV�Qg���5J��\Bi��OnbK<�X4Dľ�g�����I�oT.�q�Pgz&�����&������u]�d��.UoV.���;_[�WB�P�kȉPbR�W�e�V���<w�K����z帴�7|l%b��l%R�B\|C�5]O'O^�vdW-[ʱ���[��d��#o&)�Y��:��p�w)�D��`sUfgZ;W�4Nz9Ke՗Vn�k�������GVH�����Yq8����H�,��q�8�XѸ;���
���2��%z8�J9j�(YJ�1�Fރ޽�C��x�w�lf��C�d9W1\x�G
ѽ�'���n���wo/Y'{��5�х��i��c�=yP]�Ι4�5on}
�8y��(��l2t y�̌.޽<�h�سtSLO�-m�sL;�wD�F�w���v�-y���%\R��#ڦi��-`��Y�V�f��f�d���N��*��;��,j)���I��f4��0�9��2���V�h��u�#qDU]╂���w'7D�3/���<;jp�xL�r-y��N�8�Ѡ��
uɣD�Ai�7A��.�hQ���En�br�����éo]n� �e�Z��".��/��aՖ�3SM��_d)�a���Sz$[���OLgB��'q�+�.�G}u�f#� r��kU��};7�9�%����lŘ�����%٣M�_MzMܴK�pinst���P���ʤxPv�R�SyP"���b34���Q��Y�<�|��M�1�}p<B�4i��U�p���-V�9��mrǚ%*�V�9Z�(�:;I��1:����գ]�1������L�υi��X�w"n���pd˄`�=<7�K��Gv��E+�d,�w���ߚIlk�ѿ^d�W����3wC�.�-�F�>Mj�5,�����N��2�[H[
�V�ean��d�J�MԐ�YZ���˒h{��B-�9[c\��u�6JФ�uH3Pڼs^���/x71L<�*�fD�Pu!���^mX�1ݖ*x�(�C]��5|�M����F�#+@��A�Ҋ���i��
������H��ly�E۫B�}��I����w#�^�{�{�"j�7�)�����͓Nӑyll�b�#~���E�p��M�Ļ�-���^	>yx��.�s`T�St+u�E���`x���TѲطg#���,ݥ��9@j���q�u�����(�x���HWųGv���H!v���7v%�_s.���/ye��gb�Mm��r�[�o-u;r��k�AP}
J3,�u}�n�tX��]v�#��(_WS@kG���2���+�]t���u���RkR�s�2��0憨ܱ|��)��+�\iY��kȍ�\r�c�v;�����P:H����]�:{����>����Ve��?M��}ɎD[Kk3疸�J�t�:�%�}��łzl�{hU��O�hݮu/-��E��5/�qr�h���
�1ުJ����3l��=�*�p�0�K�����>�o�ұ(�Z�#����I��%ڎ�b,d�����HH[��ej;�V��6k�i-�i���dJL��]�����3H�B�f��S��o_PN19��v��(�UI"
�**� X��X��
���P�()+DU!Y+��,F(���(�m
�[,�AEU��`,+T`T-���H�IR(1" �
(* �`��E ��-�
��X
T�*��2*����QE�� �
�U��b�����b°Y
RVVAb��(�#�b�
��ŀ����"�`�ȲDEQH
(��mA`��b��TX���*�TYJ�E�U����#*UX� ���b�E�Ƞ�P
�b��R�QX��(���E�B����FL�dQb0DƱ��Q���`��������
��i$�ޞ��Q ����f�D���ɑo_0�s\.�1H�j}�HB��e=\�q�Q�ƹ�������v.w{�B��wC��K��-�.�T�}�9�x��}Ԙ֯�q�Y]+���x�ɔ�;y���ֽӷ�&�ƫ��n��RΧ�掿��O(�(â��b�J�.��;��8%|��	O�\%k��>̿�������J�Rg��r�k�T���ܜ�� �����Z7�~>Wd�'�q�eBTq'.���
V ���j�C//c�	��g�@t��
����h�6�����������;;��L�$kz�mBz���r�!�:���5ί1U��q1�m�9ø�UR�����wSn��!�Cђ�Ҏ�Y�Ye��2�v�୓��<��Q�\�W?��9���^���n۝\2-vu_��+�a���]�W���ʽ�G;���߭�TF8�W:�o���]�*[O��Bm��wۻ[Ƥl_#DVPV˵��}8��8�(���_4E��X��2r{z��<�9�����j�Tt���Id�q�)YL	9Ϫ��=���/y+�eĕ��U�ʈ^*C+�_�����r�՞�k-��]ε
ɾ�!��,���d�ee���=$N�����873��˒Q�x�-�E��zԗ_�Jy�GsI�/���O��6��)M^��T�g��O�s/��j��i���Z�������_J�:�Y䚌�.���$)���shV��w[�{�v;|�#���v�S
0$O�Vгf��� ڣ��7��>��-Ǎ�A������y�����F��rr&Q���Zj�h�}�I4��ù\F8�r�;�%�8�檜��d��s��at�}ws�K���v���	慉 �캆�����>Y�"TtӆY����5��חve��Ke�wӸw*��$�:�;J�&������y	�����.�0�b�2�&�ݚ9�A���'=�NL�\�Zj��Cu[�W�Jc�Ak��9co���"�ȝ'^0zp���a��_˵MC崕���Sj\)���Y������Ǌ�.S�V �Y�F*-rP���T�*4�bG����t���1h.�R-��k5��n;s9�a�Fszѳ%�G@�U��a2b�ϥ�3rV�c���4:��/��^I����r�Hg^ݢ�o����.��\�:i*��fT�.�wp8�ߊ��^V&��]��wE_ͨ<�z���Lf�պ}5��4��3�yh]�:+�Xz�&7���:�44��Fa�ͻ��c�n���sam�T�꨼���ƨ1]I�(nV�r0uͦ��b���Y�����h����v�=�Y)u./|�����-z�B���bN^����[��z���i�	��[C���죝L��M��O�^4R�����N���{����'��5o'U��ѩ/��> �&��V�{��ءMۋ-�ݕ�����Кj���=[�օ�]%�k��ř�
t��sN�����ld_%P��O�f��]����l)�h��޽=��.����S��3#]I��o�˅���ok�O"�v*K��n�:�H��)�w�T�ʵRmg�.z��Vд>�rg��uԜ�6��u��R��i/a
������Hn"�Pg/��4�����U���}��ס8�9�|�yofuɈ=֖��:�[�Z�񧙫��k�b���3ݓ9nN}S���;w4�N}��e���+�[�U����f1�Wu���N������^�xq��(T���ʹ�o��傛�+Qbp��g�A��*�������nh�oC�3JQ�}ח��u]��İ�O��r�Eȍ\�ˎ/*!'��S�i����+�єƄ�G�g����9�����3��{v���sa9���=��	C1�=[N�q�e�}��mGf��"�\���e��Pi�^gTE�3���juʃ�rξ{w3W\���`��[fn'6�B�А�o�T'����+�����sكΑ�۶��))�DޥȎ��:[���]k�o��{�.z<����n�8{��I�񸟞S��,�.��q,_te��k��⺲�����zf�C��ʔۅ�5G�ͨ����Y�G�׽��Z���]�/�p�m]E��ߞ��ؙ����o�]e�M��i���N����Cp+U��.V��p˝���b�L����Əڶ�ή|[���xv��r����,���w��bO3�g5h��xc�uh��E�L|r��==�=��wW�u=��M(�G�|;��:���8�������i�������!��9��53G�r�Y��IgH�������XږkZ����Om�z�acYbi��2Y4��6����g3i��-��?zZ͠��F�X���M�g�O`gb^=1[NgX��܅V[�]���*�_T�dc����b����J6�J��[-��j�i8[n�ڄ���t���j�f�|<�>�r�\N}�:U�I�&7y㌟�Ҧ��Y���ɽo��g���=甽��?���Ӟ�i�n��J�R�m��۷��!��Ȅ\j|#�W	Z�6�t�I���=N��du	�� ���9ۆ�7�Y	����sǅ�]�V�S"V��^'݂�w2�Æ�mw���ܞ�뵚S5]���s���zi���4���X�N�R*��� �c���Rk�?Bh*���
�hQG]DkF�m���z�h��<@��5f�G)v{����3u>�[���%}�e&�;�v��EOʗ�ϻi�"*BӸ��4&F#�]\��ؚD����ڜ^R�Ye���І	|��ɺi�'��E9�^6����x�k�7���`�u��}:S�����{�_ʩ�!<бe��w��A�v|�M�����^��t��>�xn�����M�s��D4:b٘n���l���U�(�����(��!o�6ٶ�o�v��^����żX�U�N�y=SP��L�n�rOK�,�]��[��z�(������ϧ���������>����K/RG@��vm'}���_]��
�k��^`���3.r�ue��w�,�ݱM����S[p����k�.��q�x.T�|+7�h`��M�.����f�N[�)�֨bwp�%��=��-P;NƱN�[ˌ�6:����r�x=^��;(���;��C��-�N��:��~3NYr'8���JG�)ͬ�S������#Z���v��{��:���QnL�/f�dK�f��)�� BS)��c��U}<O9�W3��]|��N��2��@b���倧x��{q�׷)��u<녝�B#rb��z��Z�6�}��hoa���J�v���qr�d��sQ�}���u���Ē.a�|�fe��SY�RA���J0vPW�C3�̡Wwֲ2�_
qW���l=��)S�6S^-	��k�-w�.�1�b���p��v[��m��6���*;��Ҕ��9;��0�#Fܨ1�~�D�Ɏ�!I�1�nt�s䍧�T4έ+~��*㩻i1¾;rg�"�]��ev_���Y�\.�1�r����o��n�7�32�+�\E�]c����#L?Q����ޘ��������N��Q�*����ܶ�E]ĥ}�<�`Wg:�o ��ܣ��^d�U���8�>ަ�#�S�1���7�m���f{R,�{��广R��Ԛ���	���)��e듸�0���}�J\F�����٤�eGX̯��aL��y26�O@���}�Ѩ�{/)>��dF���#�گi[P�[\m�d�2d�R�^�q͚��*p���ۍC\ޤݴ������ۍzz��p�U�r�.
�깧{���,�����і-�]�t	ڮZ3��ҫ��wK�sJ]�Y_A� 6���N�>է{V|��~��C+{�]��^l/y�L����xA�t,١��~D�4jN�`m;(����:�NVr�/�k�v�ў[����t��Oi�-����/u�\���?Vj���]��ΪW��kr5��"[����������d��m�;T���A�;����O�<����k�q��<���d��FG�KG����O(0.�}�����V^����b�8��(�F��9��_��������Tr5�<�\u����釙Le���s^�<��{��_�O�)�!@�I����M
�+ԅ�����-�l��b%�ޅ��x�mК
Uw���s9���Q�tǽ^%��Q0PU�B�>`l
�~�	k5���.{k|��;}ҙ�ґ��=�͗��۝󿽗X-̹RE�|QW-;��oۂ&+�+̇^P��	�Q������^�	:A��p,��Af��~	���;�rLٓ&�Q��ށ����vM���P��}y^&'���5��܄����������z}��k�5�[Wn�%R��T|}#��Q/����aV�`���M.�<.�^l���=�zwݝ<���gܕ��v<2�Dy�Q�X��`s5ugג�֕���v��Rڧ����]������	,J��|�>�B�^���M�ڴ�#�Iڔ�5�#�q��J���ә��]O�>���H���Q]q#����.��;Kf"bh�G3w��X�C�n7Ճ�n������V�䔍��,�V�����9(��X��l.B}=�Z<��rΜG��j�5^������	½[ꇬ���X�_�Eډ�5��-�c<�ϑ�Δ-����t�jO��u�\7�t�"4ਉs�ңaN����vuo�Z�|=��M"�#s�3�k��˝��8��۹�6숛[Q�z�0�$ˉ���������G������5�YY�𿺹�>�U�n���ב퇕����w�%ݍF;��1��,��jʎ"��t�Y;)��U7��x���Wz�:ݘ�������m�&�������s���S
�{1��댑=5X�@Mw�*�"��Be�7��Lh���ΰ^Xԕ�n�+�*��9,-����U���;E�Ϝ�3 �鐀Ȥ���w��}7�ݫ#66�x�F�� �!7��9H�{�q��������r�/�G���9�|p<Q�*z��3��M���x�>��W�׭���u�;�#���\y�9>~��]P=>�w��j�����r�ң$�m�Y��^n�{�Ù�E7�����X�j���퓠�4�z�_)�4,`���os����m�ZB':�7�C�鴱���C�з+c�.[AS&q�k`���O31��s�h����^J]�z�V�6yar[��T�"��
�J4k�pk�U�.�VY���%�jI�UN7k/Q�:��1����]���\r�@�"��+e��w�z=�0�y���y$z�����Fa��*��8n��ޭ_�WS�@��g��ƼtS��7_�v#Q��I�M��i]v	��WT���4����Ϭ7�z@n���(���[pf�y�
��['-�o��ݸ"���3o�{<��wz�9�f��zq���\Ts۸�z�	�dte��q7({�6����E�u�j%��0���½�"{!y��wa��2T
`�n�Cв���zd��o�w��b���o�<��n�w=�ד���k�Q{L�~��P�]�@����ym�Nd�)Ǟ���^+�u��xɎ�V9�ڋ���iB�=5�����`-��G{�O�֮�E�7\��U�{R�w~'������P���:/6du���v��Q�b].H���x�4U���Y �)̺<1������:Aw�X7�xh{�W�Q�9=�=W�WJ���]�c�:�W�R��[�7�o�C�����t��8l����֫�=y�U�*��D�����NA�]59_��.��2�RN�uM�*�,Τ���ҹ��j��� :��v���һʟb�����H"7Oi�xj�6��}b̊��֚XJ�z5�B��	�*��HDg�{�ӚAκ��MR�X%{M�A6z��sV���ܮ�� ��(���}ʁɨ;�X���Tнa�����4�V}�D�y�k�rFc�n�^s�����Ŏ���z*=���������G��GOp�}3�{Em�C/n �1�Cu��a愫���b�%�V{N���9D�o]�#���!$V���r����}N������%�d�3(h¦m������˯���NjDA��spK�j[8�}�M�ش����̷�fv��c3i��\Ma�g��~ۙ5�CUգ�v!GdB����A�l�5&�RD��z��R������Jt���%y�B����k�����{Ѻ ��e;ъ�ر�[�����}�����0�w�s�d�㋹E}�Ze��A`��W!e�PB��6���P	� �BsK���9c� �>g��Q�����Yp�삯��m�裊�YP;{W��rW���\���D��ta���.���%v�i��rP���Ն�T�]TL�;����!�1}�j�ZC����Dfw#�}�F����{�3�j��_O)��i~�gL�:3�̫��OK��`�|�µ;x�ԧWr.³}s)��'@P�j�s��kXS�3� �9dǋ�Y`�\jL�D�F�g=�)N��}Ԭ"�t��\S�ظ�.�F�7�}���9.���^������d$2U�*�7,Ry���;ҰQ�p��i'a�t�F􊳴�N��ԓ���j�w�{CLRr�T��ėj�.�
�)��p�3��|D�J��t&���{pz�"]��4�L
Uq���,Q)�u� �P#Ӏ���M�9�5�3|fṼw����xʮ���nT���7am4��h)�Y��\�� ��>\�r\�[2]P��<�[�3��ٮ���S6O��:K���+t�O(��,:p�Z�[�`���aa��㜏ID1hC�۲O�.���6��f�>N��+8�K}�M6n��o
�LN��������	�1��=��i���ө鞜�<�3\�}%kyȋ�Y���4VE3�DmL��.�P���@N��v���iu��ޕ�U�P��[��a��i��Co;3v����M�v��Z�EG�k|��xT�O	�k�jhR�0kor��W��h�q���S�S�6�W�3�i32%t���0�KC�!�A�K������ք�:��h�9$���nJ5�j��jM�;d�����V�5�Ⱥ!df��)�R`[y��$m���i	z*\v��I�6�&u��u�*:�c1�$�f�`�1* <�ܱ���Ed�1PQ����Ă����P�ӕ1i��+U�n��J�t*��N�'s4R#�g
�˩�� �����I���*J��Y-lPX��c�4E�,��"
,�*J�b�ҫE��1��!�P+1����QdR5��
ʊ����De`�*E�Pb�X�SF,X�2�9k3)�D()"���#�AJ��8�E�L�H��EPPPĪ�J�m��e�#K*�TFJ$R��m��r�2B�U
��Ŵ�S� �ŁQed[m��V�F�TaQ���1ADd*T�*�,U��aY��*Z�L@ơ"��f%AE��%E�[H��T*@SQ��`*�0*-E ��P�[����"�)Z��%VTUE�DYd(�,
�j���AAV(
*���P���QUf2�T��l��"��m
�
1�J���)G(V(��j��qmc.#lb8��AT$QFڅABUV���Q`,��CT\�
�"ԕ �X��W��߿~���~|�,�#�N�4�B���u��Ȏd,�͑��᧲��	Κ�=IN�cW�ɼ���}�qodޞ�E$��V��Km�,g�k.|r!zc�}O?J�h�d�w���v���w�o_a����z;������W1S̚�燑��R=m���#>f=��a���}N��ҝ|z�7�;����'���#%�!�<�A���^�Kex|Z�#�#�������Ox��߽�D{	�OEb��]�����{��9���f�&�t��s����.��:@W=�|xi�Eǐe�=y���Do�U{x��`��X=�2<嚎�N��@^5���}>���w{��]t�g�c�[WY��VC���~�ǊT�\�
��������MD���`����Dd��u_�^[�<�{7�{䏣
G0ۈxhrfF�}T̀\/>6!\��@7tI�J�5�@�^`�ViAXՙ�[��ͦ�Ϙ~���W+L�{>	Kmٸ�n�nb�����1�h�| J�&��Ļ�Ur�z�\��T��W7�y,zMw:�f��c��X�t=qq�*Ӛ�ɕJ�ހ|wzV�W�A�u��I������߼zN/NP��ήs�.�c�5{l\����yc��˹����g(湑vQ�;��V�B��;-�mb�K3d�\�2�o4-�N�!e����%�)��t� �ғ~[�=^����R�ħ�M��G��z'�84��/"IЖ+���]�Ԕ���AFøA��'y��!�:�{���.G�9]3\�*��Tdt����=�U�z���絓�I\l�G���/*���|7�(뙊�tz��w����_��㬳~W+�u�п��V�Y'N�L��7X���.Jv6߫���:�ݟB(��yLnw��юq��9;U�o�r��{������Ѕӿ.�>���z�2g\���������ϩ��S+N
7�Bw��{Q���;��2�nJ�u�W�X���Ȏ���Y~�q�TEm�'��x6|Ό��^g��ey�V!��k)��3�&gЯUc�(��^��+ޓ�Y83#�W�L��zW��?f��Ls�"ꪷg�4p5F���T�����YC���l�1M�'p����t��n��<�[��w���z29�G��>�}`h����b��ˀ��x�|dd��~���{�ڪZ�����iqF��V!���#S��Ź��g_�tW��^��2���sq0Xi����'��.��^C��� �zsl�i�T&��&l��'�g�W|��="y�#č�kO+g��]�4��*I���Y�q9����u����dI���|� oy���s�R��a+ٚ�}ݶ�DM�Va�oH˶h}��)L�"w����+�=;�eN��M�֕�X@>ȏY�u�od���xrd��g��.#ś��?HyXvM<���e�NN�Q��v��x�;�4�*5����6�x[O���2���LܿV��v����=��n���z���Y,�Z8f��+���5[F��>؍1��Y:.�_�VV���}������c�帤�߆d�l�!?@��>Gnn���V酞�����6�Á��N�n�mՎ����Gq#X�z�Q�� M�>��"��G	c�L�^7�P�3k�V���ͱ{���q$��b�̷U/��d���P:d7uAߕɳZ��W�ɲ�F7������/d":�^�Jg��t�q�+���g��/��Bit�28�s&,�f#ƮӾ���0���/&����
�q������`u��灿�լ�9�k��?.5��^&�������q̺v�QD?��.��~���+�.#��a�]�g̑O�3�׾�z�A[�r������C�Σ0JD�d��C�k�*�,��t�:�]~����.���+B�ʭ��up�o�5�ü�#�����4g�Y�%M}%������z����3��U�O^�S�N�#�ֹ���4��Y;-V'�6�+�5�*⦄����c-�_���v1j��$�pN@ ��Ox��z�m㥓��c7��Rژ���v+�� 3Ry@ qzv�����C�>w�s�NV��nԩ=ۻE�����g�y��"��R漲\�c4�M�v=������[b�??T+�B�Pg��*�΁ޛ�,E-z����H��Ǫ���v�Z�~v?T��~zo8�I�~�)���{�p��sN��������W���`��>]�z�m���W�O2o�<���>�|�_
����c>��v�w��e���m��o^�f��^�E�9��Q��r+�}$�=g6]/ޟQ�V�\��2=�\�`��Fc��7E�w.��y�"��^6:Ǌ���T�" ����+�2����ަ��l;Qcy�UԤ�T��
o��y���s�H�h����}~�v��~=�φu1�".��U~�����GS3��|_�vX W�,���(�|A���!z���G}�*kj&t=��g^A#�T��i�>�y���Ѧ��ύ�WT����eE�C�i��dzx�퉬��=�r}!z#�Z�N���2;ayд�0<Nd�>͌F�{�wσ�8U��.iy�U�]�U}���#�����ǿ���'���w�:~���Y`r�\xw���;�E�"���MCG{��@=�36�R��q�X(<��;49��[�e�����	ۯ�4�bT�p���$�u����]7��-���y!�:��z4�mzWn�ۄ���Y�����`�P.L7y��^s���nB�D�4�FS��7{_z�Fk�ɍ�At%]��&��EJW��������Θ_�D&pa�x������X5O�v���������߲Ϡ�;�1Ӵ�z��;�|Jsýʐ�~���X't��^)�vnra�g���r;��|#֯�Z�q%S҄�F;��l��ޅ��{-Z%�%%�=;Eb����p+��J�
[�*z[[>�:@��w��m?_��wz��]��7�c����z�$	�2���(?��V��e ���v��YQ�ɕ�c>}t�r%z�{>�zs��~-�\>%OH�մQ��HA�ļb���ջ(��� r�@eO{�p��On�z�ܝ�M��-�������ȉ��:��Kx����zuN�b%��Du1
L�r=�WU�5�-�M���Y
�篅?:c�m�=]I�^1�۷ݻ�O�To�P^��#�>S�7 ܁���Tb��R�`��ݭ�zH���$9s5���u��Kt����H�z�c�����,�z�R��6�������L��`o�9�q���%r�Mkdj4J��s������VG�z wܹ�\�=2��q0X�~�3�"��6n����I�qp�a+�)����N;ݞ�Õn��Eݺ6��=1C�-j��,^�n,f��NQ�J�7�|������[7�B�/j6ys]�{��/���C"�7:a����Y�<�-�N�K�E�N���{����&���
8�+B7�*��{��r�H��293!�o�����\�=�[�*<v��{ú��sSw]�cѼW���\b�=W+L��\�dB2��vj6ۯ����)ȉs��9ީh=�h���=b��L�IcT2^����CY;��O�I��΃4���c�'¡z���~��(AY��bjs�j�B�<|��f��(FH�q�B��zhk���`�;�
}��욞��j;T��ǻ�'���}��wU��xg=��5��Wђ�{p���b�ݫ̻q+359��]h�?����/:ݲ_�<P(�{���x'�,��ne�񸝖2�%�p<�{òb���2N���1�6]���QAt?m}��_[�Gw��h��M���r�m��cqy�^4��nn��z,�<��9훉��p���Q�k�b������,f�~n�y�}��F��}���{�Oap��v����Tk+۳2�9'�s��<���������d�mC�^���ʹ��,��X�7>�{��:�Dq� �=ޱ1�Y5��J(�!;*_�~���.�;�y����$V!�$;�oCt��뷲�d=

�rXwm�"y�\Ѧ_z�٤k,V�M���n-�Y|w#
�f��ce��d�]�p���
�8�է��下՞�ֻG��3���1:��+��ZN;nojgRj�chv��ʵ��6�STy����=�Xn�-Oq�C��x��C�"o
�{��h� X�V�3�3�U�X\�~q�Vx�foب�z�/�U]�!��t��4+]��R9��=�Ƶ�����~:oO[���a�Wn�i��"���N�e:��{�^�� �ͬB��v�'MF=6���خc�ّ����]/��۸�O��M��'���Sʘ�!�<۴��Q�qu��m�ޣ�8K���9WI�#�߼�ٶ�����Y����c���{W��\��(`��{������򻉧<O��ۉ����W����h�>Ӽ��������n�j�%�Νd��\m9�[����'e�{��A�2��#�u�+t��s�g
���d={�:�p��U��-����N�}�E�����c� �E}�$�����f��ݨ{^�$��0��W�{Y����L��6j̿�UE�8���L�ϖɳ#\7Q݄ߔ��bz�h��ޟt����Z�N��<���{ޞ�v���<M����:���E���p(].���3'H���L�}=���
=ʞ�(�S�� �c�{�v6:q&�^�%���Z��id5�H�F���#��vw���ޛXm^���:���`y5 9S�ϼ��&�J/bw6R�l>�9����sCvyziR��t����`���D;و''Y�:�e`���=�
q��m�D���;^q�Z^	ÿk������d$���d�,{��9W�������OW��N1}QxC
��������W��ic~ɝ��@k�k�c�ϼH{���4��l_�벳}�t�YZ:��;";�r�_قR7%��0�w�3��>���ވ��pW��W�����Wf��!^�1������^������>�b�(u�騒�Rf�w����Z��W���KV�\|p߾�w	��}�q�����Je��_�/��v�<�q��5����ZQw�����X��^`z#�W���{�ב>�5�O�;���Z�V��zj��,��W�p���5G�x�8���t*
�"o�<���!W��_
����c�)�_��~�ܬF��Sa�]z��ގ��\K`�]]F��fŕ<��]L<�(is��.<����~��'�.#����Ufc���*�ba~��D��O��p���ǪN�٫��;�9o!�x��W�����0W�Z^�ȑQn�m�2���dƢ�&&�V�w�?l��k��/�NYԳ�W:Y�9�[�l;r��{_i�:��ؐC�|0��p�ᙇ����8���(����WF��ot��N<�x��/�A���|�?!���Sl�WcS7��z�$�f.��e]\5[rm��j;Oy����׍�*�l �����QD��L�c�iWx�qc	�.�[��P����B�j����ty)|S�1��F��y��b��Q�C%eh��\�V��+��r3����l�};�5>fjK�n���U*a�I�^�)k��U������Ֆh��L�NI�:v|?vN���c\�oi�ʽq��u_;��0ݸ�٥60璸��Z|O��rʱV��:ju�����=�"���� ߲��5J[f4��A׏�nnP�f����cp�Ғ=˩"r<��w�P��xV���wM�x|�a�߲��秨��������W.K�[;]H��{��o�v�_�t���.��d�v�e�=7�=�A���u�e�Ȧ��]/Fy��79>�>�wq��~�q��O�Wo��x�]�����V}���?A�{p���ex>Lvʯ ��Up{�
�&S���O�?^�����<_�����j�w=�m�����V;���'�}= r��G���J�{u#�~�<��:2=��q�z��ځ�z�rh���пnI^ivw�����쩝~'R�M��/,&\�w�=<w:���̽�%����Q��虇�r c��I���z����κG<��bM�ͱ�(@\��s2ޘ(�Ҡ�6����w���]bM�����<&H��pU��՟m�J��~%���ĺ5����U�5�Q7��;���O�؅�8l�؝1/�:�~CN��|^Wq���~�c��Q��pO�*���p���4l?lŚ0f�����=o<(z\�S�R�o��u@{�	�#�v�@l�2+ۼ���?e�+�k{����7��!3���Mr��F�=��V�`�IN�ʓ�,>7���ف�/
�w�zØ�	�,��>��9
e�o�k}T͗��p�}�n���O��n�Nf�}�w���;&�G���$z��i�����;�q���s�~�Jx�t�1��'s6�?l�fn'����XMt�f��=B*B��0����`��A��ǻ����Ob~��QY]UT2h���<�����OM�mX�D�A��'�M�d�t.sW�����|b=� �ΠcM	&�f�����W��y��!��G�'��G��0Xv����9D�gN�;;��tM��B@~��U^y���/k>g���Fu�B�w�sޞe�<j=��B��Z/�t�̱�3�}�ޭ��~@�x��K���_oJp���k;����֨k^>���J�\����;�8����>Pq޶m�8�Kt&�1��:��ъW[�õۙ[��9%�ؤQp%��h�_T��7d�0o8}�:����г�񪆆�/7[;u�d�s�ъu����"�〧|�_;�1"O\
����op��k��5�T��ip�����KN���i��U���R[��m�W֟+�����q�L��b��e���g��ԭ�U�>�O��}���a$X�z�n�˴�w����If�;|;�#��ٍ%�p�O�����ٞ�$�^J��2-wC�-���������$�lE�V���4�&޺P��r�C��T��JZ3��E:�d���*��d-RRj�D�����䗮�<�yUxŲU���6���֡������8�"	B���a˵F�@cg}��Ly�gM4�-�J�KW�����>��3��L�� \�<��Qx���)P��F���}�&�'wy�+�jJ�(b'V��'mh���6��i��7e<�VtI���N�{*�j�7�8'G68�ǵ��k�1�}�o����UMg�b�/�+�}�2Ш�ƻk���7f�.�=���9�7}ŽΝ�$�;��hkc���ܞ�oK�p�Μf{|]�r�q^�;n�	���o\<��WpI����7L��ND-T�h.��&b�����%c����fk�ܸ���6F�#LT^D7lG��Ƶ�w�����+ ����u�f�tZs�on}����0�6_$��O^k[�Μ�J�c;1�D/*-���;Dv,������R�{�#S.���/3r��^�e��{���%:�a�%2ҷ��*PB�ƹҸ��ѣK0`��a���7�;R�Ʊ�r��U��ꇛ�L{�{��y����*X�h�ʬ�L���t�{������Y���v��w0����7Ci�R�慨�
��v�㮰A+r�<��,�j�Uʝ�oy�Sm�y6�������+�;�
"e�ҷ���A�:����| A�{��b��J�#���6j�!�f�2��4��i��7}���]�o�I����-��ڹ-�[�	��a� ��։���ێ�+2���
Os��-���0M��X��w�V�ic��G�8VzgFiò]G��u�7���\6;��\u�ᓱX�+i��8s�wrG/��N7y�\o.w��D�9�"�7�k�)�$��'���q.��3�V{�x��zSp<������F�e�T_x����ά�����x�/#}�Vm��V;ʼV
�Q2����}m��pt��������jU����kSvY�-c�Z��
Ѓ�3���OB��b����kC[���>����.������Ͼ�6�(���"�ȳV�Œ�����AE[J"
��*Q�b,1���1@EV���e��ETV���p�Q��LAB�J�AED�VJ�RUbʕ�Պ)R�dc
1
,1*AjV
����т1�̡���r�ɖ�@Z��Ɗ�S
*aUYrȵ��aPiTm
�r��1�)`(��� X6����R" ��f+Pmr�`ZP�QE��J�QB��d���R��,Y1
��aEb�T�%E��TX�-H��X�kI�ł�2�-�Ē�\�1 �(�U��X[`�LHU�bV��QAT�XT-���cK
��C����@�
UT����"��X�ĩ�(�)�Ccf2X���*�G�Y�a�J�c\���X"DF�}����-��po�u��iJ�ӗޥ:���F�s�G�r��Ja�(k��]i�pm�$k*�Aj��αC�w5b�=�J,-��k�J]�����\;�J��O�o��S�����o�լ����#i�������^^]L�3�<�Gfr<�V}����x:ɭ.�g}0u�NN�hco��n3��W���Gm�K��z��*�_�9r�����$��a�R7��z��`M�x�y3��+��5�:��ϙ�W`��=0e��{W9����\�i⡶�K#j�F��G��W�'x�k܋YUȫ�㊭���
y���;џ{��{ޟiQ.���7��R�0�R�&Ad��W��if�'��f~���N(=�?v�z���^�pQ^75��y�k�2���oz3xu����<�y<��}pQ�x��P縶}�x�b3��L��pQ���!������mg%�}��UB�������w�l�k�P���i� ��x�n<��!/{rfD����5:J&�v���^��L�9��a�FX��K��6\��慦&�\<�ݻ�3�m�L�T�oّ6�ĢH|qM�>�����s�܄��	���8W�,\����ΧϤ�|���+N=�}Ͽu�Y7;�s��4U]��>1X�b�@�5����
]�3o�ww)T�i����J����T��<�Ҁ-J�C�n�C�
�]�L=xSA�brtw_H��93%
/��5AS��/�Ի2��8&�{J�gb� �׫u-��I6=��g���,xmH!/x��#�u�2�H�q�]��9�yz]ǳrz�E5''�Hh��W��s�>7��� �xw��<�(��2�m���`�� $�s�=����?CT��q|L�����/�zd���} �z�1&�����D�[��^Z:������9,e��գ��N�Ά=�7v�:�b(��2�Й����G�{�,��q��d�%��V�z���m�iW>��\����w�}��g����ͭԏ�5o��k�'��t3k??�暟u��e#���o�ݧ��ZY�Ş`k�k�c��;���bu�,��o,��j${���������>��ܣ�R7^���LȾ�^�q����Dx�?�3�gFwp�C5�u^aꥧ��B����[�ð���,r�0��{>��p�ǫ�N����[S�_������/�p�u;���In{�>�^�(�� ��q�񦣽[���b3�n��W�)��ex��U�^�)>�Ƹ�,=��i������^��1�9_C��T�=�,D�J�W���)�#�0P�C��+�k���x[���j{��oc�ݣ��׸|������h��]��<I⮕������y�N��}�QB�1w��P��JGRϺ�Ҽ�>وJ�uޢ˛#�kR�t+3��	��	�= s��Т�o%�3�ڹ�Z��}ï��M!���z^Hc��K7��Xj��\��P�)����+�a�P��ǵ�t�{D��Vy�z�7A�3������.s} k����"~�(����6r*x�V��d�9���CCz�k��������N�C�>uro�X*�}z���&)�Z�&[;q2�W�1���3w���Pݜ��XE#�`3!᠓3����l��}X W�"���$����%?�k�fyF�o�~����;����J_�;}��p�z@�)�����%=��]�|_�}Kw�λ�S�'k�|�nXY���}��3[,i���Ǯ���|�T\�ǹT�s����p��W�^�oU��ۋ�rl�?ߋ�G�s�k�����}q�����_���`Oܯ����]83������_�s�x�WQƛɯM|�M�#_�0�$sgj^W���g�7�����c�P�u�RC!^`z=�o���{��r<�G\ye�B����,�Hv|�����|�j�豫�gN��C�+�K��qj��SordL9F�1.̊_ԔX���X�<�N8�5b�<@�T��˜�{��T6(�N�-rgT�x'���<tC��bch+���$�J��XhyjZz:��ծ(��;x���&,U�5R���-P��os�����}�գ�}w�C�u!q�%���0��=��^�C�����y����ߢ&��%b���ll�����������^��U���QE)Ӻ��ᘓy��r��>��}T���\z�e9�}R�\J�X��[ご��nᲺPO���q�&�n�2�^��N�늦�S��n2Pl��n�z��h{!�:'ފ��a����YWeG���>�4_�z���w�����D�4z@�3�8KeF��Yْ�Y^�!m�V��s�}���lg��6W������!Nx�8�Cn*�'����V=Z����Տj�ٴ�F��ZF���ԑϟ��/}@h��[��W���y�d;�Ns
��w�ﵤ{����>��w�q�٠�T&�s����x�����ܬn�ʓ>����0dط^���ZCQ�D��v�������_�a��2��f�{2�|T[.�\���Y�uy�ؾ����h���>'��Ǒۛ���Q����Ek���FXۆ����?�*�X��y���?Ev��.�`3S�+q���y�LJg�M]�Z�#A�z�\��ݔ�v�(䞞�Pn���<&�㛼E�w���g�vOnp7�n1}�G&��U���^h��T3!�d�:�"�=ev�ջ A��ZVN�Ƙ��� u�7�.9�6z�K��K�Q]b��f�2������M7>%iϤ����j�K����5�t]Ly^���Dǩ�����_Z��%�B�qq�#\ߞՏd�A��$>9���[��m{�$oB��Ճ{�u"��}��
�;��d/U�r<������P^�8;��2�ۉڇ�|�?j��Z]���Yc�ga�v/e{��͵l�'�n�����P瞜�Q8l=��05~Bey�V��=��蜝emÿ�|�oO��E.���L����ϛ��k���	(�F�a[u���]WV����>��Y$=%�X����FL�/��b\�w���~�q��~-U^�1�4z���V_Y�y뇜��QQ)�8]Sn{ŋɝ~�������=��4���}��x˒�M���)�r��]"���"8�Ǣ�W�cx�k�<��5��w�:T�F�&ʬ��n�	�7_����z�/����u�,�}���R�|�:�'@�\MCn؍�xW��f����6Z��u�,q�+�<y[�Ǔ����;����~�_�B����7$���FA��K�P20���O4�������῰w����T�U3=7\m<�W]��SSf��a7jb;��	)Yu�v7sZn�Y��d�H/vx�]��w=\���dh��hY�D"�79�-�t�֠�Go�y���p<�y��s�1��������J�k�\�O�]�������7-kꂊ��\Uå�l�G�~��c���XV����=s=�p�n�s�`��dy��@ /)��
��UB���9���n�e3_<J��=�ϙ�'��yg�M�I�7��`��ҏ.��ں��U9(���49�OTk9��s�w �^��Hz6&��C��n�������1�>�~��7�U�}@�ҥ����W�R��&&���z�ù���h	�@�S^�;�^�9� ��VN��~u~9·���� t5Q��?OxЈ|r�������#��-�����n77�h�+�'����ڭ�	П
^�,��@�/�=�ٶE����g�3 P��������\(f��)��]��<:4�&+$&yUK��2Q����d<�6v��q&0q�Cץ�k�3�i���3=8=�;[7��t�y{�Y��n5&��(����������(�����ǉ�=�Cn'i���kJ��
Ӭ���gK�<�5L��|n�:����T!�G������+���m���s�Y}bez��p�Y8ɵ����\�ף��2K��&�fgX��ŧ�)e���I:
��� �]Og]�N�\����m�Ő�Vz��roK��k�+*�W<�����˾��/쩷�7,��|�haOt���"��o˃���7t���)AЋ�z{�ùNϨw�uy�-o�y�s���y����.5*�.�)Y;)���|ׄ��Zj9����廜�ο�d'_����}���|����+�\��4d{�)�J=%����^���^���+q���0=��
��"�mPL�ПPc\;/��A[�\<T�����ٹ�#Q�-�=���>;�`r��(	���7�Je�7ׂ���Q�ґ�����9�}ǰuhx5vt����\]�2��Ey��:�ϯ�@l�����ar�7�Kgq���p߭�
��}51'k/ݻ�o�锈�l�+�)��*zL����*�>�����T����FNN;��z�D�����=M�=⋗�U�r�EE���V<W�9��D	[/F�r3���͸e�iS�7�q��r��[��e��
^�����"�-׍�r&Z<H������qMYq9��y�WQ�-����imzk��u~9�����@O�,�~��:1+���:̼|rW^�)�HK�lx{6H}���MF���m)|n�Q��F�|S�>6!]Pq�5Dz��D����&їr����`(���[��t�o>��@ƾ���_;�-�-�l�������k�\�eu�ep�K��k:�7���E\)���qI���bm-O�@$$��t�U�{[τN�z��Kk2p�iffe�!eU�C�}�,���>'ۆX\n>��q�Z�d��u1�g�n��ގN��`�6���V��쫬���7�����ߕ?��xH�8�k����^N��k����0/|�zɭ�P��쩼Ѹ�ƹ޾�Ƥ�{Q>�	�FC_�p��*2B���{��8`��d���*���p�\�k�U�:}~��~�������xrUv����֋X't�Ix|��4q��z6/���^r�v2:��<X�ˣQ�}�V�tF�؝2j�[������^�C���A}�%�wЏB0j�~v�f1g^�}���7ѝw�gT/܏��ZP����/s�h��߃>���þ�5�[���{��� OTA��W����ø��N|2>}t�n9�y�\�)������~��x�˭SX�O,�#�Cƚ�ߡ�/�]�ɀw�������A��py�\�>"���
�ٶ�䵆�ƦUw��B�й,��q.��9]W���D�^/3_Q��w1^��v5�����j�����o�����K�nj	��ʓ����eȬ�,�:��~v��y��SU禶�;�T�T���;1��uo��i�8P�;�wF7�֫�Ŝ �����v�/zK*�j��z،�Xp�)���uym�}��rZq%�"���B��]1��d�����1u>�N����E�7Z_j�"��o�N��>�Y�R:9ש#�l�[}���oվ��
�|���lk�gZ�N���mL?z�`=���ã����L��|�:Nv�6^N��s~��wG�ߙ=v�� �b�ۓ�-˓�c�n`����@��,x�s��.O�:�}2�2���]�}��Mc����Z��g�/}�I���Q�0�ۉ�c�=D:�Zdk;㼌��ݛ�(�f��x���J��ŭ�_����O�EË󯼪I2�2{�|v�T���aT.�#�0�y��l��}��ŉ��J�O~V^FDy�=5��ǰ<�� �$1{��2�L9��{n�\����p�]I�>���f��� ��N��s%l��g����vb���黉���֩�3�蓹���%�Ƴ�%Q��8sɜ����z{)S&�q������uH�Э��9y������9ղ���Y�鞤�aj׃���C�i�.Ɔ��R���tZ9iH�>3�aC�ּ�Z���_�9����dZg��b�����FMiw�d��`된���ĽL�
��zTf�{(��|�3�>�k��ֽ�ǓDM}�N���߮��Q�5ҋ{;}��7*}�ۜ��v[�~)e���:�8�i�'kA�J���ի����~w���Eo�%6G��^<;J�^E΋6�!����L[m�>q��8��&s��
���������Ԇ���8_�L	��X�ɝ~����SPf^� όI�����>�&��-)h��j9S�����e��Yx"8�>=4������l�{�W����6��٫鑼˗����ߞx��@7/�P���d)��;K�޹>�b���,9���^yj���k�I�6]������N}�2��C�0O�������(��ߍ{`u�G�7�(�Y>% ���JhT�@�KG�����%qV�֑ȏzB)��7�:)�ֳ�>���[�d�P^�O����`��L��.|�h,-8�_�D{����zH���0E�3Y[����o���x�}��+#��N�ʒ2$�z�$s��&Q�o��×����g���������ٗJc���~�ϧӰ��R�O�W���-�r�%t�o$^�Ey�ߣ7;ebr)�C}Urx_��^6���t����n�o�X5>�n���]]P=�>�����I�Je&a�='�}���xh��;�k�E�������ϋ�DW���l}�=1�k
��
�!�*��������|���kFek����ۮ���焨{X�Y�4v+f<ӑF�b�p��Fޚ��e̵�Q�bِ����K��+f�՞ʘr5�7E09���o�IͪT��m�6�&冧�/�Fг��߲��nk�_S�W��^,�j
�G+ֶYW��	D�gZ{i̫3nwl���6�A9�4ƫ;�ofL����)V�A��e��OM.�ڃ���n*�l��<>F�ٿ��h@�NGO,�����sQiǩ�zv��Y㚸q�#��,��e��⡵Q��"��7��v�����{��
0�(^fF1S�����U�a\'&�f<tusw#U*�dHR
M��┵���/���=�EB�nt{���3��D�!�}e�/�V�b�6�K������m��7�2�qC {�]�.A��֥���E��B�5����g�9{���V��l��l���3.��v���\����ZI�{��\�R���+�`������9��9R��6�!��mq����ƚ��Ŵ��l�>z{��H�njNĻ疴g-\c/rtn���Cu�ʣv`�'p;5�/C:O�q
ν:�G�U����<�Cד�z�1{V� �nlnaq(� ��N�K������ׁ���3�"_H021\��gp�1���:�Ƨs�u-[��>9�+�cc�Y=�Si�]�k�4.����MY�{aXX2_.�sz���6,���`P�jeM�2[7Z��z�=��uɦ�SK�-e����8l{���W�m�"�7�m,͇;����k��{ˏf7B��ʼ�*�7�Ǜj�T-}�����aA�t 
9��=y,X��eG��2�u�@;m��vr�)�+�n��gh�ǥ��GSoRb��f6��If5��C=�v
�>�pLj��À���k�[M�4��ΐ���e�yo˅��}��,��@���1P�m���զ�t�q˴M`�9���.�L��:��Ǝ1C�ޖ��k(��J��SՇ.\�׻��NgF݉��i�Px���6.]�� �[r����V�baN��L���-�z�z��ж�B���Y�g�)�Z<��~ߐ���}��kJ��2�Ybw\�Ʉ�+5=�p5�j�gĒ��,�,��=�x;�׵��-U␶ٷ�>��P��+���.�q'귷7�{L��´%ٯ��P����a�f�a��
v�o�k��xp;�Mo'�ɖ�mƽ��y��?q��4)��VA�h+V6��Gw7���k
e�yb��y �u�"&�;t�G8�P;*Sf��h;�����B�j]�b�.�9e�q�F��ܧ���*�y��Dʠ�.��� #�ggX����6��+�{�[��DkS/'خ�p#%su�Jz��ik�o	,,�z��w�+μ(�W2!����ǯC[m!�7�5��Y0Ћ�\�
�,��:�����+�'�ɊȌ�̭K�L�����Rc\I�Q����"��,P�Z�*4����,��*V�cZTm��KlY(���Y�����-E���B��VҊ-b��Kl��QTP(��RZV(
��V
(,���6�VՅB�E�EjV��6��VJ�hbQ��R6aYb$X媍�#
�J���Ak@�U�Ɍ3(,�"��,X�U��f �T&Q�S3-�Q"�!��$�"��-�J�*��Qq1cR��,��b��+1X�j[d+�XV
b(J6�E���Dj����Y��J��WY"��X�����(�"H�D,��k*�Ԣ�[J�Ub��-iXVb\}�ay9��")�n^��:�0a3(�Es=`/n��g��㒄O{��Y8����v]s\�F���[�Um����_S�����o�Y^���5�����PLоY���Ag@�/���{�K� ��*Us��=�`zG���\L�{I���zp:����K雌�`-�\{���Q;;�u�6���w��ғ9�M�`���M�5ŝ��q�ʌ��i��V��Vy��O���T�c5~�����$y>��|�~��Q��*���{s�.	�7%��Ϫ��ɭ,_�d���OXQ�wYuA�X�f!��(2�����e���W�H��#������e���{nQ��R$;'UT?���(���k�͡�ӿ?�CE���v!�ʒ2��Zq�|s������ P�"zv��)q~W\;�����씀��V�{>���&+z��d�>�����=��{O��W;��!q�[����9�f���9~���Ŵ��������⏀�����Je��jģp��Ȭ��lߺO���?���z���W���m�D7y�C�e� ���+��Т�p��q|��Op��3�yE��NL�h�sʪ��Ǔ
�9�����[�~>�����10�]* /d2�o#��$η��~����ԙ���[a߳G6���f�F�F����f�\n��sUZsPf��}�8�Ey|�ܔ�T�;���/07�3�^�j�#$��/�][W26nh���5��Ƹm5zٱ{���q���s��RJ��]��U�'u��0��C}_[� z�{���&X~�E����q06-�P��Z;q10�QH�����]��'?t���+>%q��c��Se�R����`����w)ύp*e�ױF����mݿw��$}��[F�4�ǹ	�����{ʯ���{p ��B�ڝ�џ]�.�k��ݍ����o�	�ς���c�d����5�/�����w�S�%��y�n7^�T�k*��LcZ70L����?v�*��������cL��ǻ��2=.BnG��к��ضיּ.cܕO�۸�s�̼$ys������>��tV��?�����GT�D�s��mtc�&�����!�N�`�4��4ʌ"����'ˍ������ҽ�����40T��mi΍�'�����Z�տI�u4NDy֎�B���|�N鸒��XrxC�R���+�R�s�9�};F�K�{�rF�ء�&�8�{v=Zw��1�\)lc�9�����2���F�3����U�+�w�;���H�S"�9XX�	�������1���lו>K9_9e��5���#��-��G,h6�B[Z��ft��j#}������X�:S?C����aZ����-Z��UF����Ɵ��hZ���w3z]E;CU�v-��=1�c�[��&ha�9q�v��`=�\J�+Veʹ�:g�T��v��<����r<w��U|g��T����ýڤ��c�_��Mѥ;������u�8���ݼ��,g�5����JS�s�,��6@�j'���0&����J��2<�.>�{_?�2�oz)�|W�{�;��n���{�$�6���;��K���JG�7���r#���m��j��f��ݾ��ڕ� ���ϓ��.�����yq�Xn��Tv��lf\b�,m��Ǖ, s.�Ϯ
�yi�RG��@�����wB���sN��F��w�U����q>��WD�A[.͂W��!3A����z���ǜ�*�� <��='o�>�N���:{T�1N�'�2��s�TZ���p��f����I�F�}T�Ln��e(:�Ø�����C;��������{,�V��I&9�7Lu�z�u���"�^ׇ Xˑ��m-�h�}�����7�(�s��^^{���$�2U�TM�5y���O�I5���ˡp��܊���}Eό1��΃sP_�ǔ���l5�C��H!G��ܗ�n'j��`	�O4M�X��M����
f�[�����t�çu4r�C���1�\,uB6�.�Kl-�ٮU���M�fs��D��Ruƺ�ff�����Yۢʸ�[]���@�}|��Z1���[�֋�0��
n���fU�ޛyz��62�@RT��~�*|l�o� '���3�uG�'<��W�݊����:rz�v�*�ގ�$Y'ɬ�������א*l�W�8h)�������R���Q�a�K�ٟe��v��/NS�'�G��O��L�c7��[p�'����7�p�W�d/W���N2��7g��+$���Me^����X��ĺ�ӽpp�6L���d֗q�;鋝t�ޚ�-��W��н8}�J~@�J��}��o��;��(�Ä�K6mSn{ŋɝ~�#_�M��)���7�%ς��]�`ަ����_��P��eXn���"8ȃ�*o��b�wB��8��,�[8O�iU�ʠ��/���u��[�B���.�9N�q��:���~���o�عߐ�5&�S'�x�\i�����>�g�s�Ѣ����7�#�x��7�RV�d�ǼNh�9��Ш-��v�>���9��\UïZG#ސ�d��Us�Y���s����n7�#�=���и�z��\ �0n�P����@,-9����=�L��^�N{����L;�*
m��;�ʺ���E����j˝W�,��ˑi-�U���-��ϓ�gƦ�X�]*�wnRV�R\�����.��=oI�q�;>q�T|���ǫG�� ŷ[�9������7�����z����A�H@���[�$%W��/8��|O'>��eM�iL�<M�qځ���&%F�������^LI���d�ɭ��,�:Ӽ�=��ˁAE�q�8�{��*:O+�P��������}��5������->s�g;�G�7(wdx�p�Y:-�U����9���=x��"��)s>Gzb֮�Q~��u���͟C~�S���]'C��}^������~r�p^]�+�_��`Yqy�.�1֬����bG�5���W�4/2B�y/M+I��4�e�d/Ux���s��w8�_�::I�-�+�g�<h���2��q~SyU�����`R��l{'&�x.���g�9����Q�_���9�#�6pq�=���Jq;Le��ZU���Zu������52VL��/�C^��;������3��Xi����+��������2�kKs�L��@bJuUuv�����Kݧʛ�;��#-ϑ#�n�~eS�����I��BR7%�<�ˮ����O�'�ޙX=x��Z>�g�{.�^L�9[u	��F3�����9�:�=��%ݡ�=���A��Vx��Ms�Ə$�B���&9oe�P��5��і�5VZ�
�BX�ȺћX*�X5~ͦwA'�A�VM�6��]}$s��[�EÆ�ղ�P���a�0�]��Lc)W6����R�e����3���6�5\�|��틥�ڸZ�i9�Κ����>�:M�� &����˷�p�r?<�ί_��x�_d_�<�od�Ql^-E�힚�<o�+��H�@(�2��y)�ojģpߕǲ�6r6���:v����;̳�l��Zi�;�F��dq��z�Qr�7�Ǚ�}D%�<� W�P�fv�$q�k~�x���G>�
�����P����Я�^+}EgG��\n˭P<������ΐ��]�W����=�\�����ndH���7h��L/y��X�s*����ӛ�.$0�gp�Dj�����{ԑ�����]l�x� ������x�x�I���}�{l�x]��&Q��%{ˊ��f�И�}[F���F���k�Ǽ��r���x^k�]n�/5���m�#�{�����am���ٲGh�9p�.OgBң�Z�S�Fln\n���Md�~��׀VO,����g��_�>	�nXY���N��l�&J�Ǻ�ٯ]�Χ�3��r���t{��Ψ���*�7�m�{>(���/NI�;};^�W��V�<?ǲ��y���6��e��حDQ�iȎ�������?f\�7�ϋͧ�V�-Q�����+5;0��޵�% V��(4ɅKy����,�M�X8�}�b���b]L�Jp u���9!I�L�3�B���c��2�0�����w�G�>�oU5�p�$����>�W�*�����|yQf�ݕb���L_xOi�-;0�]�G^��͎S]����r�Ӭ�����Kjߤ����'�po}喅}��_��[�б�s�1S~��}�e��m�emC��WY����>j�fk���[���!֎�����sۨ�����ʼ�H��bO�y��'�Gc$�9��
�d�8�e��:�E�����S;��юO/x�;��̮�{�ԟB��j�z<��+>�UL������1}�y2��d>�~9�V<j���`(���N�����K�>��-����R��UsVYY��x�ޙ`tT����A�f3G����޵#�te�s���ߋ�~��s�m�zJ�!֎��#g�y����3?q��[�Sjo/iz�c�=(�>gx��u��瞾<���%#�1Ͻ�t�?_E�AX���F�,�91�F�Ys�\�w�3VT��Ng$����	h�1��T��f�K�6r=�@��=`h�R�-B�d7�yF�ݼmFfg*�Ōx�8�}�FxǴ��f�+�e�24�T&��&l�wǷ�q��uwӛ�k�9u�cc]t���V]��<X��B����]ت�����ŧG����t�v�%������X�o��L�{�-ʒ7��Է\8�����:JԶ��>VN/�Ǐ�!+8r�a�Q�]On�-V��C+`��7Gya�Ҏ���Hb7�����]`z@+��ˎ�qݤ�/<���Gp�x�s�C�6�n�bun"v+��}�[y�	��YQ�b>�{�'tI�Y(����*���=D:�ZdV�������-g.���\���>s>L�Fc�jc�{·��lx)�O���lA|v�����,��6"iL��y����l�}�z�3}H:n�O�N����J}���D�+�|s+2`ۛOkF�=�qG_��Q�B`^׸�zx��� �W��ϗ���9�����
���v�6#i�O��{h�j�Κ��@Ti���g}�3�_\m/{�[��x�,��^Ȟ9��+�E�LO��t'u���w�=�ͭ$��X���c2v�_����K}6��u������q�^Ufx�Dׯ��g���?&{{���x�*��3��X-�sجLοΖk4��S��r}~��h��׾�U)��G9��s}I���)<V�<dQ�{�Q~;QT����`6C'�F'1{��x���.�什vi�8?:�=�_���K�q���du���0_�[��]��ϲ;������Wd��.�Jك��`��!{��B�*^֜AV'Y�Q��E�},�q�n,�;*s���M�=�����
�Iu�V�����+�3}s��D+���~vEC��]t�zD�1_u��٪�Uӥ\�HK��Mb�d���j�S5ؕ+R��ޝ&�ݖ��~E׸��y��dy#M��yW�(0��Qǡ�������A˼^#���e��φ���#0�R�"o�+��>�(��uǰ?Sg#�'�vo����g��stT
Ʀ��]ߒ�+�Z��@!��t���B�-��%���mdK7�G[�ZD/\`�y�,�Ϯ��Fxq�}�z+���^��L�K����a�Z�\����|����H��#�f/�� VJ7��r���vĸ�I./I�a��A��z~�T&�:A��]G����s�U��_�3�3����w�,���;���Q.*_�TO�@W��Qn�J&�v���}���<Vl��\�������1��T��j�ǳ�e�����m����),��G���1ʲ'��T��7W��V[�֭Ɲ3&.sV�`���|S���+�k��Yϼ� �P�^y�]�M�׷^�=;z�ϙ���l��+ɚ��
�J�bk(&hr���q1x�b.7-�~}Sx�'�d�9e�{����6K�Y��A��O¢�c<��;�� &>���Wy�	��рR��gMAV�mdj@�)���<����B�����A�o7٦!�S��4�ܓ����g\��ׂoecH��юjH��7�OgI�_�%���PLT�g�m���t�7�Ƅ�Ƀ�70ۗP��Ft�(*����9s�o��>��G���2fNc�#=����i��dD��Q��d흇2U,~*�������xE��b6����]����K&ؼ�x��o�����|x��x�{��F�����eS�H�4�\q9Qח�mJJ��c�9�#s��׍{,vF����^G��h��}��;c�\�^`��/v����Ez/��q(�d碪7�g]1dγ쭻��╼1��OΆ�:��=3��xNp�k��E�K��v��${"ϢJ	M�G����p�%_-w�%�\{z��#�)��y���*�U5�35Z�X�ұ[��><�t�;�qX�Sw�p�Z��bQ�o�#�X]�o��i���ؿZ�ݖ�����ޝ���έ߆GNQG� �ٯ�H��#>��n#%�3����FϦ�1��o-�%���{��?z�0����F�F��[�u�>%���ba���Qf{�1Ϯ�YN��tuʮ9���L����<V�\Kv�X��}:N]�"k�����q�g��Z���Cs���G�|�u��-��IH��#P���#�"M3nr�<޽_Ӟof?�	 BI�R@���!	 BI��$�	%��$��BH�R@���d$�	'���$��BH�䄐!$�r@�����$���$�BH�yIO�BH�b@����$�Ԅ�!$��$�	'�$��	!	�	�b��L�����n B8� � ���{ϻ �����>z���D�(���7qѭ �%-d5�f�:�%��%"�Mf��,wZ��Ef�[5mV�R��5g�ܴ��ٙkS�:�Z�Zح["UC���R�mh�3���΋`]ͩ�I$��v���eWl����t��p�'Vٶ��5Ymkk7u��͠+XِfKi�p۬5���VV�m�	�M����J��M��6ͣj��i�.�scU)��D"�    Lh�JR��C@�4b  h@E=�	)T�       s �	������`���`E?��4ɀ	���F	�4hs �	������`���`$�I��& �#D���G��э56Ԟ���~F_���	$�?�>����撐���H |АC$?�l�BH���������h:�g�F0' BHA*�jBI!L&APa��Im������Q���|x��B������c2t�}_};�s��Q����ڿw�U�Y��t�����雘�:wy����3&7��5����y�eLb�	Sne�?=�-������V3J�ז��35`� T��� N;�1Ӑ�N4@�巍L�b����FM�3"��T�ز��Q�-��f�)��	zӑ�
z+"ޛtb�"�Z�K]�� H//u�;���qL�su
�Z�nV%��@
�&��w�Qv�2�t"��++*��khU���
����3H��n��`Y[z3U	w��z�g��&��i6��WXY�t�&6n�+t�Z���U��)�F�ictn��+X7Sfs�/�grf�=�)�d�-��nV-����(�2Ey������^v�o
��E%J;uj�6-���FQC2�VV�1�P��֨X5'���aR�<zj�ҍasi��4G�c�]�R�r��ujp�ٖ���Ј���o���U(����%��gt�~���k�]k�cB�͙Rǩ^䛕�buj�lvI�%�����:4�6�w�[�s�ԣifi3@�����U���8�3o.$F�ڽ�rJe�49"H�x�|R2�&[��<���q�0k=��6�u��6葩Q�ڸ�j����+F$�Lӌc�,b�DΌɁ�U'v��VJ%���Ib3)mfزd��mBS��E[;CU�]�d"�"њ�P�	s쭭)T�0��OX�ڈ0aB"�ҕe'`�yYz�A��a������MJ*f$;ӆݣzC�oY�ե�e�+�q��kN�����J1L�H�
;j�3s�G���+�]�r˱f�e�E3E:�/1\	�Y��v�-6`uxLn��z��W�q��Zsl6� `vui����L�V
��!'2U��1ma��<כ�elt��%м7�a�ȕG3���>7!��MV�ը@Tf���[��!S-���]
�q�.���+E튺�X�t�`ԩ�̤3X*Z����6"�;��0��F��b9X�J
:VC�8�n]�Z�@�,X��b7.�'�n��/[�q&�-�F�i2^XF�
�u�u�$n��H�w+l�1U��:�6��Y&�*�HFb��y*�C2�;��&8�X0�6��t�=M�;���m��em�W)�1�{��+7����N��x#����E�ĭ�Zj�l��)J�-!$��i���N`1�#�^-ƫ�[ٔ+"�f����)�Ӵ�9,�Vl�
*țb��~��ϰ>�O�֍����*�է�qB�?C���~���)�V�pF�l͆6X�2Hma��-�s��0��R[����v;q�f�;3��v5��ƨ�tq7Ql��'��,к��ˤkl�àT�G��񃃩���6���m�๻@�c���H�����wW�gt1A� �.W�#OjY;�1e�Ԗ�t�8
��}/&m0}�R�dXŇj�����#%d���(A�o*�K�J���s��!�93w�z^ִ@���Tw�]�=�wJ���4&���Ak"PfYw�b�P�(���p�r�X�j���+}W`�XK�f�q�[{O;L��O.Ɗ�8�,flS���)�e��r�_\n\Y��O��^(��P��o;J�=n��(*8.whk��n��)^ܜu%j-�"����iX�_^�]�۷"s(�2��q8��7��)�Wy�"��Q�Yt 9�A���fD/��'!]�_*]\�B݋[�M�9�k_]�r)oڗϟ�kxŻ�3��X�֭h
�w`�����]��C@�q�S�U]��FG���,H�٦ok�w;�)汘��u�h=�_##�z�L��������8���K�X�y�O{�x��qp��q#Mh(��h"sN���|XΕ:��Ԭν�ս�&"��j����Wtl�e�݁����&��[]$�1�2�4ŕ*Pėh��.��Qw���o�u�&�V`i#�$t��_0��w����N�t��`^7Е�^<Y�ײ�YMu컇M$�M-�c���q�6ܓ����b
�=�o�<��Oj��;��Q�<�����)N����R.VZ�e�5}v�KZ���hvm��A4d��)���z�����N�ؽ��8ar�.N϶}0b��m���x���Ə�d+M	�,��ɻ`F����Ws�]R/M.'Qxj�L��2��K���o)�ۛlZk$-��k�^ �|�]�%�hJ�CL�վ2�S��}]M�b ��;�%�Q�r^5������E�Ý�e���tu�	�{꽵zq�nk���;NY�/_lln�+i"E��+q���t$��D��wu;��%6��
��FVs��;�w�����u�X�**�R�yL7�l��~M�BZ��EIZ��(՝����0���]�)awU�M���W���D�[�d�а�w��k�꠫���>����Fk�6.��GMv�O2����ob��0����8�Z6�93'5�cժ�6��?��O�������~������B�	�� @�����O��$!$!�g'�wϏ�G����{����Z�8�e�x���^N��.�;�2�)�m�����ε�A�\x�wpEK��u�s�Ee�t�|X�kWJ�F�;���S3ڲ���p�!�1WIy�Lvޯ��w]p�%�.�
@a�F+�3b�YHU�a�j��N�I��g�B��ι%��1�͔�>.�S������)���^sm|W<�Z����቗��S-��k�Fh�"�oc��$��N:�WS_L�'f���;��R����\U�^��L�3Ҩ��[T�gQͬ��|��ǭz�G��]ϏZ�\1^�;;�v���G�]K�`�v�0�R1Wk�[,��G鎦9�b�
�[7f!ä������x�0˶(���|�����2�hV|v�~�xN
f����������i5�LgKˑ�u7-�����[��m3,mê�ID��˧Ku3}�d�4(e)ʆ'�̺�Vř�����i�! ߷	�C�(:�<�/>U���ֳ'�uԗ4�vQ��cy����t68!K5���1"�qś�Gs�wE�w��dx�=ZV�q�
0Ꮖ��xT\�ݭ�I쨢;����T�E�hֻG0"�u5fmI�BK�;C��!|�`��8�ψ�Mে�_D���T�7�3�L\E҃���N�w�7��e��(�w��Ol���c���WŊ�kn���;����"�A�Ps���n�.ӧZ*��ݘ�;Ep�7ǹҔ;w�7\+�u\e$j�mr�*Cf� �\��K�=����-�(dC5%{��6���*�cୈ�r�ЗV�
� �f��`�a\���l�\�t
���N��r_�ܪ��P梒���N�\[kxPUm�v�K���sD��P�C��\y�J��ZgP/VEIcs-�8D�C���UU�fi�e�
��㩸KՃohWH�(�3^�o�w%ֵ�`�t�I58��f�j�m�_un]��T���ș�qvU��7 ��(SwCRx��@�]$�s�g^�ͫc�Eh��(u4.Z�B��k�Z�.ۺ|�j�:!���eފH���N5���n�%D�o��f�h�VWD2���˥HW@��gk54-6��� �ҝCS�@+���J(��p��O�O]�12M����>X��ѧBqa����"�&Ʃ�hܘm��&�N���k��fq�y
�5�E֨�ݔ;��o)R0�C/reX���A��.�إ3OZW�+�+�NY�*WK/+�[5M�~������r6Ņ��Cת�9�ۧ۞��~I��9ev��@�o�0r��ζ����2���y���Y��L#�l�+�N�%S�i�9��e[ې��++���,\]u�TG(%w��6�i�
�Q���Ί}�620@�l����kF���@�;)�r�Rl��:tV�M��B��аEA\[R�l�1��#ZT`ŹL[sU�ث������(єQe�QcD̕�T��R��12�Ke��Pպ�L��n3PjfS�"+U��pr--��ˆ%(����"[�e�2�jb6������̤����Y϶/G��Vj�^��m�����ȉ.�/��䱢�=��d�7e�vf~��ofjSGr��>�K�� D��:�m/ (]�����V�$yy1Qu�#�?~?�ᬎ͡n��<�
Se�.)��o3%�ڱW��k�jӶWuDwJ�<<ǅ����6���*PD��>ׄ+k�d���G�!0�T�ϭz�Q˶�z<��ƍ�1��X��}�厛��B
u�2�'�#��K�cY~��M�»1mDex/k2�3(��S뺨7�*0Iϯ��;:(a{�'fĖk�w���m�+ۑ�4��l�|��wߢ6"�n��s�oZ}��xjz��"�4DF�K��s�gg�7�'Z��×a����˦7f�����$��|�߳����g{S�rV�j���Ȓ��vR����X��'Yd7�U�:E�Bf�<�4��G:ՆK<GZ���Jf�3vƠW���\��/�,%��7k��\;�&�_�K����e�XvQ`��}]�lv�[r���OV��{��л��Sw:�Ѓj;�9zvW�Kj��q�x����Օ�Y�@��+��v<ʮV��mƕ�Ry��3�V�<(���T��Y* ��(��M�2�P��.��bq���˚;�<�#6�s�/��ϽBw4o�́��t�b���~~Ī�.���Ȝ�[ ������0,U�G� 5��}������U8���v�FH�*�*
�h5o�}u�y�����F����si����F�� V�J7.!Ųg;��κ�/��w�H�׷D-�gp��6��TrѾR����F��i`폏+14���[{:~�Ġ+��չ��Wn����t��
F/Yj�2N���M+�F�f��}O�"�&R��pކ�P��O�Ҏm����1(��Ǜ��|�����������Ll��[���3J��Sysb���>�Y���\v����2�zKm��A��e���Pe�i�u��=W�R�F�g�
t��nzz�lG�>�6���X��7v�h��O�Oq��1��*��|M�S�;_=� RCS��s���V2��z��vY�He@NK�@J���"�-�K�u��+A2ԛ1[Z��9C0�}^�������z�<���S�6B��**�`��Iwy��Y���᫢�;a��5�Bc9aEϱ�6��	������D%���x�d%�r)w��&�!��
�fe��<YQ��7��%�	�Hݐɕ��]+������Z���[�a�� ��iW3-�&[k�j�����c&:q1��M&���E�C2·V�5ea�u��B*�%�Z�VL�-V�����	͹���dړl4�z�@��i�k�sd��1��3Mq��@�����]�� ��?���s�;�%���jah|ldqR3�gg�[�U�v�>��;�3n���p!!�k�4"��.Sz�룷�Yp�+/���OQ�W�k6�WXsV���dlX�;�^�>aOTЯn{���l-�^���37y�\n#Ŭ�k\�r�ߪՓ8�[�E��d�W����8�{$�����������2ҐsklZ�ny�����Ҫ�XJ����������7�!�c�X�YI�E�kUf���q�8�<yz�f5����z���'�桚$wMx+>��V��9���[C�}h�u���+�ö�Y�i2L��.BC�Hr�m���C���C�mr�A�oz���!'YCĒi�Ch�!9�|;�$P!�$H)%d���L���L;�}N�^|�Z��+�WYf�-�/+u�kծ��<�$��HVr�āθ7y�rd�i ��AI�l�m�}w���x�11�<I�$H,�2O[�Z$�"��&�!���%d���*M��	'l$儜$� s͒2C5I
0��qй	C���@�$�$�Ht���� ��C�w��M�C�4��$7��>z�'lRB)$��Hm��Bc	��󳫹!��!!� t�
�>kεט<~�q�,�~��}�?c�^�����b���v1�[�j(��=G6;Eӯ�	;��3� �b��o�H��]Ϋtl��0? ��X�K�G~He8g�]�Su��2�-v��[y+��h���S�e��ʵ)�6N�:�zʆ2�l*]6���OY�>�CL?`6Ue�w����/�h�Y	�x�:̙5�3j�$��nf+{�uI�% �|�mV�U�4���k�yؠ�f-�̈�E���,輸�
��w�e��t�\5�s�ݬa�a�����h(i�r�=[2�;S�OmG:�3����C�NY��l�Y����1��n����أY���ȜI ���x�O����ا�LL��&vdF�l`�"��.�׽�3S�F�`I$b����^��C�'�ދ��Nw٣��O7��ismL���w~�j�T�q)���~�Jw��|0+qA���9볩����d��숌��\��@BW'��'�w���L��
��p���M5��f�o�a��-gW�[�=�G+T�|����!T(�*@�7Q:���]R�|����n�	9)5欣(���^��h���qŌciKP�jP.fa�F����.�K�It�g-em!��nE�F�v�Zb��*
��Ö�������G�]D�Y5����ۘ;Ww"���KW[f���RWt@DX�&��d4i*�N��ʌ��Yyt/1�L�d8�BiS,��8ءMdM�n�a�N��RL�F�L��fФ�F��"���_��p���}����ULJ��\ef.e`��*i����P�J����Z� ��Em&!X�Q���h�#hTKH�<�={��G�9ٺ�B�m7��i�E�M~�O�N�;�ox��-��z�FT����۷��C�c�_y�f��_������a\��/C7ޕ~H^������-���r�Cjn�8�X�� ��	ujk�^���$V�f�f��޽~?&�y�~YW�z%~a{���q<����G����)�P�k>�k.���[��Od�s�č��Sn�;��kx������+���I�������Hꔮ��h���U<��%n�-�y��C�oa�~�*+\�<��M�y �ҟ��Ү]�����[�U藫�]x]��'�jx{����2r%͡pG�	���Y�բ�Ank�qM��h�}�l���{�|Moî��M�^���gV�|��3�V\EO��8��ݫ;j�c�_��EN_r�\�.e��������_�b�¡��g�����x��I���{��Hb����}�Q\2a������ǐ�]�S�C��E>��gկ=���R���C���n��Òִ��{��WO�ҋUM����љ�n�YC���X5�f�U̩��ΙB2�A�"�M���}���-�5�BO_]M�}Ns_����
���Gٸ��Q.���=)���< ��;�N��zLa��h!4���)i�4!H�;����9�c�g�-���A
��6��hyQ��W��iT�{�#{A&���ȌQ��G�����>�]Ik�n򃫔��އp��x�}KHY7T�FG�Ыë�(����ip�޿��0��M+޵�*��i޳�0XvǊ�:�35�ӊ�V. �y��"1O��_|�D�i�z�?D�۔���  5c��=<�̩��Gv�?�Iw�W�J{�m0�g7�1�%�U�e^8��۠��믗��6i����n��o�"�yR����³1�:��g#MdŬ=�;gU')ƽo���j�NDwk���P���ɕ���ˊ�`���p���]眧�(�ȫ��O�V'�|e�w�"r�f2lD,uBoNYJ���bD��ڢ~�j.ͻ�R[5C[�J�@�VQ� LNќQ{�Mŝ���L]\��8r��֣��t����8�m�F�z[r����KE;֭t�n����o5��f33��^�"����%����ֹD�i�K+��w�3��m,�k�.Yq����*N��,�aE�	M˙����em>נ�M�6�U2&�� �t¦aec��Y ��Z՗&\����i<yO>Ħ]�y��$5mB��[
�¥j4�Q�2�"86�*0J�"��m�����XTZV�mZ�X��b��(��E�������F������D@ ���_vUrYQ�u5z�~�9T��6��ȡ�D���D���ԫ�~ٺ������{����-Z�^
�ޤ�I�g��^
ɢ�:xU/`4��w��1{�ޖ"<�V���o�D�׽&V�Ⱦ�%g�,ԫa��V��3�<<<6�17$~Drª��V�<��Cj�_���=��7����údv���ަo5 滆��&$�bԼw���@=�a�Ũ����ǣFH�3�|c]���x{�3�*9����W9Jd���N����̕ڕ��"~k�<��wK{:��4�W3�%4�}�\���O5xb�;n��z݃�'W��A�/�f���\
M��p�e&�7�x <����C�����ډJ�Y5q��O�.x�S��!x�'D��|
�43ʕ��~ǝ�c�bĶڨ�4<�Bw�糲��u��;u�� {v7^f�������%���Z������;S�����	m�}h')��/+�-�z�I���
~݂J�K>U�J3��َ�+ٯ�R��t�"�Y�^�W�oj��5~��,*V�l��L��8���ʇ��P�FwE�a#�/������W��j�{:�P!S�i��
u�F�ᖕ?A���=[��L��wK�f��%+`\���I$��k�u�ǽ�=`s��{������WY}*B"��ز(C6�rϏH�5�q�yǤF�Q�c�γ�7�8d̳�ǚ'��IS��l��l��MH��w##�q����=�-f8�����8f:N��Ξ�:�,W��!��X�_�W�۷R�����c'uTn�u8��oo_�����V>2>����	�kέ����)�T�A^�����w՘��4�ͳ���2�T�_Nq���=p��`i(����{���<�����p�ҧ��5�Y�m��Rr�ok�:���|zb�
��8J��W5{MU�����Z�LG�>�H1c�wU���N�R���m>�9��:ӽ��m'm/����#�����OI�*g>��63�6�=�3���2w�R������6���$�:�����Z>B����+� #깦���^!�w�xp��'Lu�T���o��պ�:혂�eN˴�ۼ��oGp�EN:�O)yÍ�=:k�j���s�[���rQ��iC��sJ�׉��޷פ@���2>���7�W{�R�����`�%f󃜺8q8v���	�m|o}q6ʚzN������]ܒ����9M�������pM��|�oVi3���s7�2�bO��*7�u6�S�VT��8u�w�]���Ņe�}x���f&Ӗ&wK�����M������&dX�kt�f���{AcXq)P^��W�Ro�RþT�x�1u*��i�&���]Ի���w6�;1G�,�E'�*lS����D�R���:]uUm����k��J�j���yM�-^f����R���<����OU��]-T.&j=�^m^���)��[�|m9���1�$���]wp��Y'�R�Ѝ�k/�p�����^j&:sN�4g+l��{j�]�n���ͤ��O��)����{z99�wb'4E��QE�1�U�j-��*c�bE�b�h%1+�ŶQ������,���,k[Jڅ��qpVTh�УmU(�%[*���������n���;��5�O�����\��=��wN��׮ӏ9�\��1;b�v��=����G�o.ӄ� �Q7�X=_���@r&<3��y���|�%>���1��0zC�Q��
B��{#mL����Xt�<���0�3�<x�'6ɶVW�Mf�z��K�-}"�P�O���Ý��oыw:�5���W�z�1��c/u1�Ã�5��(����9g�ᓎ�z�zH��s����v�y�:㉧�'��3��it2��^�PT{�z�{�j6�j�<wf�hi�.�y֞�ۮ�ZmAP��� �̃q�r#q�^��۴�8�d����N:��SY։�b�n��"�q���T�Kz�o�@瞹:I+*f���4�L6�PӚ��_[�Ӕ���w���]3�r���!��:�g<�wM3��S��;w��5lp��t�:�.�k�;�i6�5<�a{x�w��ӄ�4��wJ����vô�,�br>'d��4F ������
��������2y=��b�m�v��� �� �Ȩ������9=k}^Fl:N^��Ӝvq�i+�"�9zz�z;������x�Y3�5���t'��=�(m���n���I������S�YI��3�)�m6�8̇%��3i��q͜�<��N���e:M��;��o�T�6��X��vz���'��б��St)5�^��	7ߛ;g9LOI6����{u��:��m1�br����ðH���Xj�r�wsz�s�zf'i���z����N��p��4�t8�q�:� XL��3��Ǥ�6����m�;xyO:��p<�d�D�(,�\�^�V-Խ=b�Ѥ7�<<����1�Uh!��^�z��Ku֚� 5�P}8q�ܾw�9t��`�']���{٧�j�;eCl;N8�z�2�k')�k��>�״x�˷o%�G������Ӯ�7��'8L|e%M�,��.�q��2�<.*
U�!3^��r�3�]%N8��I��m�w�8eh��=V|�|�V}��`�i y�u�b
{��������1�1�OF���;f�Gw�1*�/O,��\q��M���zJ����Îy��Y��R��F�`h���yǪ��6ޱ���ӗv�l���!���p�sa]>�S>p8�G���� �C#�@�mxC��v�Ni���u�K�*t���>��4�ei�����N�{�l�u�Rπ���^����� ڽ�ۉ�1��OL;����m6��z����4޵�8�2c9C}Y�8q�\��4�Öb)�Vy�s��T��I���u�m^Y�T�h�¥x9��8z|M�z{H,87��+ȝ�yO6Q#� �}�2L� dvK� Q��%<��N��S�����,*�������s�tI^�μ��t��7}wW����8M������)��9�x�:NZ�&e��0�9ɱ��NҰޯ5��48M�������]4���ᕕ;�^\�5�2X�^%{y�����M�k�DjO�BZz�Jń��ޭ���F$�)�����j�����WQU�.��Hɜ+�����N��O�
J������x��ĊP��Nl�]�åi�Q�&ʑTH�}z�lӱh^��g+Я'�9(��:{A@��u�^�3pJ��:�_o�o@���^<�
�,���S�x'odB�/�J|�:ŝ���[����wOz����W�ѻ�v[Z]U��)�4p:�S%�v�٧�]n+/�,�u�w_��y�o,
����O���zϜ�8�)��!�9�.^`�ݹ�tݲ�Zf�S�<^+H�ܧǏD�o+�۫6�f��b8:::G�H���إ�q�%H!�W�o�nl�6�o'�SL �����	9���4��i�S4rƽ�;n�����gt�v5��NJ�����K��DhfS��(�V�5-kP���9�$��5��UkVc(��V
��UD�
�%�[r��>�P��j����,�/��-9�of�����v*�d~���_ˎ�J����d�Vs�ٳ��������z�����V��_�NY�ߍ?����rr�Ъn�h�037f��{.t�ަ�/��{&w��lT�#�I/��kN����\t]?�e�)�a�ɥw`��Gv��/L����K�YC�x�c�N�z' �:��h��TGS���YJ{՚
����`�iuՔ�S~�Ԓڸ?	�3�t��ք��,��-�G�o"�;�!������	n7�~�9�͜��2=���F�k���o�D/Ai=�X�N�8�63��S&+��u}�O��
$�^��>ͬt|�+�:��=o/�.�ʼQ��K�"��h!����B;��=LY��0�v��������QQ\�ź�=��^৫b3(�75��������_�{ON��Ɔ]z[�J4�0�q�6�VE:�<�,��Ǽ��-�km ע~S�=��B�,Jb����^l����7��cp\�]�t���ȺerB���+u�����xf���H3#�O��!�΢�@�p�u�je�Mi,��NNyf���5ܶ���D�=��5{�&�.p�����]�9p"+�R�@������,�I�W'|�L��Gm�q[٘�ڟ����|+�$�wE�߁�%��Zz�V��>����1u��Z;�ˮ�Xn��Ч;s�eˌ)����e͚�`C�'�@���n
��Ոj����\��@/.b&��I����6'��y���,ף"i�șܥ>쭦r(=u��݂����O����x�[=�t����%��\Z�r��2D�ޜ3��E�1�m��{x�-�Ӊ�o�=�~�Y�����"�o�����":��jO>U�\���A-�2���e���w���t��8�|u\�C�|N����k�U���E�K�Ǝ�0�W	��0w5e7��� <�����=Y��5ٔBC*ڳ����Y Q^\�XO{fu^�IZ{����#H��)]�2PL�s��F�Wt�5Ed��*�q|��fq��9VU��f�6*�2�pR7҇,zN(Q��;����	&�к�q��v�CUK}� ��v�����4Ey����c<Q뾸j�+��#t���*ɃZ�i�*I��S�/�@w-�ֲ*��YyR�,�wE%����*��}��̇$x��@fl_�L�����K4���98���W%�S�%P)�e�f�3!7�EF嫀e�i8\��s2�����W*�'��1���\���e�m)�L�0�\�ȦYT��**\�db
�D���T���"�m+D�M|G�
&�]��tի���d������=ặ���ջ�{K�Gq}կ�d���Þ~�<J�~��Dh#	�IS�\��Q�DMMy�nA�*�p���/�8�����$�(9�:-#�]O���-T�ϯH����_��:�͌�����ˡqѵy����.q٪ޢI��U�z;»��1���S������=����L�
����MХm�z��;;�V�F�n?k�D��my*�6Oݥ��XD��3�ԭ�K�=��
I�}�Vř&������w��v�N^��l��9����"jh�䬔�Zsn�,ҭ�F����{nr���T#��zLY^�h]�B�po��<�/n������U��Bba�'{��m0M]h��2����t���6�y��y@��Ʈ�W�Z��d���alteM>�M����t|k�V���x�f�K����"yE+TW�8��Ip�XB��w��Ы����l����z-:씣��a�o��Sᒏv�ُa�b�����tۃp�2�����i(�us=Z��¹��^���'���y�)[�u�Y�4�<ۋ8q0�͐a��LЁ̔�1PX�z!�9�D��hAc���5s�v���M<��9�G�=��/	�V��aV�]y�����Ώ��6k�μ�)�k��b�[�N�|�l�w%�
�Oz��_��3�o�^���
Ow�}�5{3��	���*d��Lw-��:>y:wq>�=���"8�4	�]�#�-L�9����n�S��!G5�r�|M��x�~e�c���'����IE���� ��dӴ� r�/P�¥�Vg�x+'�h��e�N���''6��,�K����FO��I�yG�P#��%�Nyj�#�X{K��;��c_�)�����:^f��^��`�=�I�>[��be,0^k*�G9����l�
�n7sS��M=I��j�}�4���3F�K��S��3�OZ��i�>��SL!����Z���)�C��lr� ����Xp��,(�.��v�P�"n����\D)�|kX�����NH�d���&�Na�6�Jm��Y���#���֜�Z�n�Z���0݄�*x-��;���\�;qY/#)�����-'Kg�E��0�+Cre^��p�x���͡�͵��x�[���ܘ��Gp1լ��gL��:�J���kM���Mҥv+(^U��%��4*�̼�j��N�;�1�H5D�Y��Ry�|��j��S�m&-A�M�4�[aªʷ����vk32&A��d�Hˈ"�s������-�5p�"�P��j�;q1b�Ջ�������q���h[kke�1�(�TU31�T�[Kl�#�lQJ�feT]g[�$�}:�I�"s޳��ͼ�� ��P�7S0�������ǳ�r��q�6�h�ŕg���[!#5}�P`m�#O���1��d�1���d���q��OY�:��MËy�ع�ɻ�qg�]m,�t)�)�2�L����	]p�#�ҏP�v�ıVv	���1S���K�������_u#��-�T��6A�vL�j��8ÊG�����	wˑ��ȏ/�m��B�rt#<U[�ĥ�y�^���J�a��MR�t��ee�Q�*o\�̯la�x�hT^�����|X�p�d�Щ�S����X;ט��+�,��NRsL��C$�^�:�o}���]�,w$C�U�ג�ɫ8�����7pb����k}�r��J[���)�d��Ig\��8I1ם��wuY�CO�@����[�.�f��O����c1��eM2�k75��#pu^�Qm���1�&*B)s+��BfMq���|z�W\1.1NR��"�R�Eئ+���!��8�&y,�d�S����xI�o'���)VL؂v�[���m�!����x��6�eL:ms�U����r�e�7����4;Vn-�-����^)�ŷM��6S���0��$ݺ�j7wQy2( g�g���qgט9Qh��;���S�v������ޜS{Z�ܥ1^�S��XA�D�d�t���u�'��bіTx�u��a6T��˫:*�^���Ď�}	y,s�4��6�؅���{��8`&5�Rlh��;�_�q�
��7cJˈ�Jjgc\1%ȍ��*�hk[l2v�L|$50G�\u�ِ&8�������c{�@�����S40Ǜڅ�e�Ԧ[c�[�\fd5�	��5�=tr����$��.�>�+^x��s�*D�#�IQi�5S"��(}Һ��m��#��0n��*8B�fb��&=1t;�w_Ws�0������2�j[\�O.U���'���S���8����/[��q���N�,J�`�9%��u�ZB�e�.aee��t�+����Vy�1t�ŕV�/o�M_��#6,p�v�v����î���3au. �4;ݖi��_���'2k}�������A��ˢ��&�j�q�l�4�U��ov���kW���g���{=�CJ��Y���1�b��x]��sW-0�F�9��hH��B�DWJ���U�e�t��З�U��B+�gyvr�Ç��'(��]}X��(�+�HXA�e#���̤��Qb�l��Y˙y�hD3>F��y��2��-`t,��5,�WIjTN�4Ң�u�h����q��y���\�k!����_T 4@EQ�G�[J��h�唊�eY�QWI��TƵ��0e�U1�km\�s2�(U�Qqb53%E��2��3aG,m�LЁS�{7%��*��m,l뷢�t�@Q���N�fޑ-�Խ�b��]���2t��2<[ov�.�x3�Ц𩏻9.gn�8}�8s�֥!�zύN��T莂�.��4Θ�tup����M㝥t�WbE��o�Om��gʛ}���F}*9O�n�S��J����(eĽ��jf��[�VѺS�OWӟ9Mرw�mK�W5
#S9K�lC}vF3m�מ��Y��p[i�����*�FM�J���PFi���*��`���vپ߲%=��ڂX�ڦ��]D�,�v`�<��������l��v6i�����zj~rފ��lj�&w.{�c�4�M!�|�T���O(�)^�<y>�����G=�x�V=GU�]�oDۨ�54�����QW��7ѷ�q�B�7�M�+�84P��l27W�4��X�x9ݕ���'Q��.s|�~����Mfe=�;m��)�bq���wRȕ�#��?HRя��^Im=�'sTo��;�c��̍� ����˭K�{N�0`���5eZ��C;Q�&뵱a��$��9���{�1������sxk���ZQ��;7Ԣ�̌�E�~���qT�����rlЍ�|j��X�)�����*��m��-��;��ƅ�Ɖ�/R����K�����!�fB�6#xn������BI�fn�>S���.l�_[�~6�՜�#N��s@��EԵ����nf�d�o���\r�F���=�d����S���ܽ��h��a�S�>��-c��{���h�+�n�vT�wx��N�ƾ�X�:�߳�Z4 �X�}�e�\@����ӅK�^�/���u�9R�*��I��kr�z�p���fW���dh_i��E'��G���Z�J��ypV=��zX��x:�/Ζ�žs{�z�>��K��aY������Y�K@���i?	�ȳ<�˓c�g'g�ײ��=����ۓ�w�f��gN<�Bͼ��g����J]\H	���R�e،�Y	�د�1�x*������ZC����5D�Z�08j�	}�I�b���2�x��q�nۘ������+�'�ƻ.�MM�/���ٸ�Z���<���j��T����uC�=.�d�8lYS:
��4i%v+���g4���l�E��-���)�4'.�$�9q��,�Ĉ�u��J�E+��qX��\�.=���/�_djn��~y
�wk�@��H�o(I��K�9�)��u��k�Z��)����Xu�72��[c*U�BZ�W4Sm���:v����.!�܍�g�㊍�(���ɖb1�-ekS��JcT��شr�X����մ�6�ܷƢ�5*".�.8
���eWe��s-jŸ�bVԢ0W,��"=&����8r�L]�)����~3ʀB��Ȩ<a>Wp:17r�8)m�����98=�<Oa��oe�9�]��iզ��]��ź���k5RzVq=���SXsVT"8�m�=9c��e-���׺�R�Fckj�8'ާu�@��^�W�)xSS�Ҟ;l��ڪϒ�{��]Q���3�{pE^����~���
�V>�������LfwV���:����]��;8]=T�B��WZ�M\/8d�v<crZ]j�I�<rlgǮ89+� mJ3���71�� c���a�(�װ�mg����f��_W/8*���:6=ΰ�*�4@�M���d�����şf�`r"�
~OUb�j��8(.�%ׅd�|��L{��NǢ�W�Փy���|���C�9vG;�����S|T��V���y�<����h�a���k�*ߍ�:��:��)L�ѯ.��*�e�n��;��
yq��̭���YRgQW�H֖n�m���9;сgv��{.ڽz�J�L�j�Ap<�`�#V{8�����ɦ�/��}���[d[�.��Z�^�#y�)aV���u�����o.��-��e�ɋfkre�}�N��s��0/RGM��d� {�2�u~�(`�S�}��'�� �M�næ��7m�f�A���F�����c"�\|4�H#��ٔ�AI��1�W��]s8�L��rM7\���sVkʅ�5��Rrc�Ҝ���Z:�v����砞7:���z�BXI��k
駄��?-���e��+S��,]\Zu�6�fQtf�j���56�d����;_o>��	�m%�Y"]�^*���'�;s���cZ��=��;�B��T�箷�0g�~�3R7\�i�Cxⴇ[�u�W��^�]a�H�&^p�M�����y�z��ޡ�� ����gzk�]�&��2�����)c%˯3��&�+��y�{�p���d�peOkv��f�ɯ_���+���������ҵUU[B���@BHC��ag`BHC��?D]��[tYy�����ߣ����x�LIk�}oG��4t��<!����g�5ǻ!8%����	�eB�H���v����{߿~��=�g3�s���㏖����Y֡��o}9����}�^���Y^Nx�k���������~]�k����@rO�B�	6@�B�(E������_|>T>A��?�a?~��ol��p>��}���O� �������_���L�?��I�g�:&8��n}���w��Hq�~��%�h-�3p���>�?/���O�_vO�q7s�g�l�!$ ����/ͣ���xB������xU��d�~��%��_�!�8���=��I{M���o��q�>&���XMB���l�w�!膻=�	'��5�ϼ��S����?���S��X���yc�|�Cݿ��}_h{��5O�O~�'�P,�'���������}B����������g������#�NO�������}"z�~_A?�{q��N�S������3���HC���@�����:u��}�����C��:98
�pO�l��I	$!����Q�?q2`���tOs̒I!d���I>'�6_��<��,�y q<�@���1��u�C�����s��i�vI��I:�Ϭ��}��>L?C������>������=��Cw��mX��D0~�'���o���� ~�����k���BHC�>����>�_��I�~��A�@BHB��p�#���?H~�G�'��|����p~��o�r3d�
~Ͼ��1����I��O����q���~�����������ǻ�� ������#���~_(9�V�á?B���{� y>t��{S��w���h����g���$$�?�$���>/�?W�{�?/��		!����6��}E&�Gr������}ٜ��E	��}���=|'3���H�
�p�`