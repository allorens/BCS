BZh91AY&SY�]�Z�'߀pq���"� ����b._                �                            EJH�IP�) {p �w�N�x���W�<�� h  =���)�H�lp�: W `  0  S @        � �� ��@PQ�$��E(���*�%TEQ$����$��QU"��P�  H-؀�TV`�(�����E@	o������s��ʣ�.�A�|���ν͜��]�8zh�k���Ͼ���J���E3g��Z��   ;n�JW�Kb��;}���}j>������� vg���A��¾��� y� |�	. ��ϰ��������}
�  : ����+f[P+�E
R�QIQ@�}��;�wn=o��`y��O}����}�F�����V� -a�|p4���k�ăǌ>� <���|�)�:��6��aw�  _/Z�R�� G�����>{˼�J����7a���!�X�}g�M�<�J���)����y���� {Ϲz��  G�R�[X |APH�RR+����U9�^`;����`����o���w�
S| ��>|�=�/ �}Ǡ>�����ϥUg�T͏��u{�|   �W>��TR�x9 ��k�w}�o .���{�>��>�ܪM� }�P�#xP-c������{�}�p��{ t�T  =s_e(�P�E��
(lb%| Z��҂�.C�>��` ��Ϫ�>�fύ�l�poXx���y���4
|o�+à���`�6   3=��vԡ�p_X��� 9����(���)�vS��<�������� �R���y�u��   �m���)@�R�D��J��	u�R��wpz�`|��aG-^�(�W< �����<ڎ!�{��� 9��J�x ͞@�.  �o})V�d������0 ���UF�
fǐh����Gs ��� xuUrǐ5sT��y >           i�L)R� ɠ    O��IU Ѡ �� �b'�R����� 1  O"����4�M@  a��Bh���� ��  �Hz��(�)��6A�i��6��ɤ�O��W���*)��
N�������o���~��{�����U\�LP����O�qEO� *�� U��������1S�����r���t��*�`���dEP��O��<����ك��̀t��لq�q�q�q�<d1�x�8�2�0�2��
c*Ȍ�&2!��c���.2)�8��7�Pq��1�e�1�q�d�C@��E�q�`1�c�1��1�g�;lc:`�q���g�`�q��<ld�3��3�c�g�g�q�1�g1��blg1�`�L`ƙq�1��1���g�q�`�g�c8�3�x�����v�3������3��363����3��8�1�c8�3����=63��=����3��8��`�Lg1�<cxɌ�3ӏg�g�`�ǎ3�8�3��1�cLɌ�3��0c8�3��0c���q��q�g�:q��lc1��όc<c�gx̘���0c8����1�1��8�3��3�c=1�c0v�0c&3��c3�8��c8�3���c1�`�1�1���Ld�{d�g�c.0�&3�18��g�q�1�`Ƿ�0c=3��8�0c3�c3���g�q��q�1ǌɌc8�3���3����1���q��q�`�1�c�1��{`�1�1�g�q�n��q�g�q�g1�`�q��c&1��ǌc0c�7�c<g�g�1�`�g�g�q���2c8�������0c3��q�1�1��i�c1�d�`��d�La�`�d��&0c&2c��ˌ2��1�g�g�c��Lc8�3�c8�163���1�c1�t��1���q�g�xc�8�1���1�c8�3��cc1�c�c�xc8�3�c8�1��v���t�3��3��83��0c2c8����1�`�q�g�;q�t��c8�0c�c8�1�c�������cc�q�c�q�x��1�g��q�c��L�8�0c8��cg�q�g�1�n3�c�2x�3��=61���0c&=<1�g�g�q���zc1�g�1�blg�1�g�1�g��3���1��3�ct�3�c=��c�1���8�0c0c8�18��1�����3����1���q�g�1��1�c�1�`�1�8��c�c�1��cg�1�`�1�g�ǆ1���1��c8�1�cǆ3�cόc�1���1�8�1��8�1�61���1����c���:g�q�c�q�c��1���1�c8�1�cLc8�1��3��c�7�x�3�8�3��8�63�q�c�1�g�xc�3�c�3�c���:`�1�c�q�c�n��:c�1�c��&1�c1�`�q�ǎ3�c8�1�c8�7lc8��8�3���1�3�c�3�����8���g�1�`�q���	�c�n��c�c��W�U�Q�A�T���G��2.2�0.0�������� c!�c
�"��2.2��c"�ό�c
�a\`\a`\a\a<dd^2�0�2�22�2�2.2�#�#���������)�����20�L�������#�)����L`a`aOWGGG<dLeN2�20.2�22��c �q�LaCC�Q�Q�A�A�S� ���q�1�1�1�1�q�d\dLd:`dd`^�WCGGRgSGSS�`W��D�P�Q1�q�1�Y�1�q�1�q�1�1�1�q�q���D��A�q�1�q�q�1�1�dGCGSGGG{eq�q�z`dLaLd``a`c�	�)������
cc
c c� c*� ���8�8�8�8Ș�L�0�0�0�0�2&0�2�2�2����8�8�=20.2.0�0.2!�0�ȸ�8�8�8�8�8�8ʝ8�GS�Q�T�����ƙSS^�q�q�q�;aLeaLaLdLd\dLi�1�1�1�1�q�1�q�q�q�q���A�@:dad\eLed�1�xʘ�8��2��+���$���8ʘ�8�8�8ʘ�8�8�2c �"ʇl�#���]������^������s���C7?ׯ7�(��jBg0��<��S�ovWpӛ2�[ ovh�í�NTK����WY�3�{'F����7�lz��U�:�5T���I ���_r��[������%ݹ�$yFQv�X��t�;�j�j�`�s��M��-6�s�zc�Ί�MQ�݁ly(O���ծ�n�ð�7z!�����c��ν�������`p�J��³�ϛ��BĸpY�v����@������#�7�+��ν_j�	ؓ�r�V���v�5��7��6N��;�^�we�oo=<s�5�� ����'Ewa{�^2����Q9r�7-0Ɋ)�c(�+�����;ȸ&��.�-�2o�����p�{M9�N�܎�t�*��u����"�U��d/�V{/F�4��X͙&�f�;��b�kA�j�A�ݿt�´��wGf�����S=+�j镁�ۯw���4.ʏ����H�׽�P�E�[�F7�0?���殥7���wC�i=��3od��΄���U�3t�q�&4��BQ%#h=��lR��P����@�u}�t�!��ӌ�p%�뽤�-kӰ��W\{hg9�v�ou]��%E���J�}�:W�9v�"Vwał��Z�(�Ђ�,����ak;�'�.+$���uo>�z�Fn��ݖ��J��`ww5��*�0��o�7���&�f��2�,�FY�����F �js��5r7���Õ�~U�^�zH� #�������os���Vm}���3,wI�/`�����6�&��L�+ûX]��-�&��0��wJˡN�Z���ɫCO�NK����B��a�������e��b&L��4�х�۵������} y�6h�t�eW&�p6�ެ����O[��G1�`������$��vl��*P�����#��d�m @f�r��
�C\y���X�7@�Q�P�.!��s�}� "���ܕ��5�oaޙ�vI.L�h�����F��cwH�X�1w`絖-%E$[��A�W���2vP���Q���KWk�"�(T��;�F����e�a��i�|:���2�;����Z���d�u�⢝xʹgE��{�f�r\���T|Blt�p=��k�X��\�w����c�Q�+�(�v��һ
禇�w��t��[�r�$��	��N-�I�Z�;;"��y��`���vɋ��Y`+��7��I�<q�`H�K7�u�A���^X:�׆`RE����v�¾6kim�h�nNGgזJ2l�o��ݮwl&$��d��ǠۃT{�5�1�{cG4B����N�k^/��\k6[��-�xެ�8�M�1��r�-҅qNĞ�����*F��;`���,Fo!�ItsV�E�su�EEtgv��8#ӎ*�s{ƌ^�^������V��3]�oK{��pa2!��qiOu�&e������b�P�Q
�����P"�.�;���-��٫5m�:�P��u]���R��.{��>|���hk4���ē��q�2m<�֋ )ؖ=��7�ɝ�̏���\t	��oN#wm�TS`yb��cg/��_�FP/I�C�1�]Ρ��,�)K�q���wt�\,<��
>K�3�/:w��AF��Ổ��곺�4����}V��x<)���T�1;�S3��ue8�y�G�7ri�d�(�h�u���"1��{����:�)���y�X�a�PpCO� sc�����+�!�PG����vڻ�m�-T�u�r�{�p�sD.�~q-�n�B�f��vRy,cc'!m(c�q�KJ$;u��G�s��/%u�ږM�.4M��7kһs���wT�\�0V���w]�{��4�Jܭ>Zy@F-�����ѓ�w^4�Ի!A-U;V#.^"૭4NOF�	�� �]�@W�1-�qkՍ;z�M�A*̄��C떹�t����0�g����.F{L�bC�����w�����0�D�ϻ �#q���,�A���1�ۮDS81f�{Wws;�!R$Oo`�7��YG��g$S��ob×�c��t�!�ts	Bn�ޥ֡�^�j�w�7D]�VJ�OL3$��x�&PQ{b=��M�λ{X�74�H���)Y�t��G>�o^aq�{�S��n���U��,f�ע� a�q����)�z:�͝T��&������ug6FM�6��up�%"��H�{:U�p��)w{����e9F��
'�f��7�ε<����J����u�0�;;y"��r]�N媨zxt�Zv\SQY:�S�5N���wu��yy
ţs���P6.���N�0'���F�.?����JNAS.ă���A��!ïbq9Na����]����b�ԕs�,�����ۂ�GfT
x���=y֮�ȋ_#6r�P<CFN;ڄ�ǣ�l�˸N�9݂�k��f�M��p����K]����
�w�o=�n��M��+�䳓TvR�B"�0��f��)���<D`�H�p:v�v���8�EY�:m�͑T�5N�n*ds{@�]]ٕ`<w4��ʭڻk���_f�Ϧ�ʆ�!0�o=.���a�֋!�9s`����hO�Z;
h��{��ỳ9i���#'�߸s���qԢ���W�`J� ��[	�P]k&^�m�ڨK�3��*�Q�0P|��O�ˍv=��.�D3�+u��IP;V��p�Q�+�c糆&#�eN��>�f�6���v��f��:�9��q�y�'��1s��%5��6���l��N�ں��vc��e�:af��L�#F� Ӡe��ٷ�F�\��y��Ҝa˺���R���8ݑ��9��Nj<]
���� ��t��c�¶J���+�;H.��t����$���a4���Y�摚W`lAۏ{b}qt�F*��#�sYК �tn\�afi}Z�ЪUч����Q��W��V�B��n	�s�&u`h�>v��Sv�vT��x�mݡ���}�.�f���y,�d�\q���˹��m�Sb��V��.R-Z�n��:�=��͝�b��Yۊ�Ck��l�p.�w�6q�m�ZT�Y��� �qǱ�jg@9䥕���Ѳ&Vv��9��|O6>��[Ő��� Sx9�1Q�`&�r;��v��dzQ����K��F$X�w\�=ް��M�:�]G	��V9s�e��<����#YR1 ���,�f7T�`�</��V�^܋bN�C�>�W��^��]nuͻ��X�|��6����#������IY�����IVr�~���%�b�x��`-�F�賵Ǣ���d�f��|��� ��L���n�kTzء�dcIiq@�o#x�z&��j����H|އ���{�Ǧ Yt�V){S���L�EG�ȘJ����{W`�����
*c��9��<����3�+�,�ۡs�S��-H��e���wAQD�x����RD.�a�G���>��Z�Ѵ����c�����wovy2�Ӽ�)L&�j���']� 9Dz±蓜�i�z�盍���p[h٣����Ѻ�'��_�Nr��/Q�d������,A-�O�"Mo[�^��|��$k���О���'���*=3B�r�A��ԇ�u���7Wf�������CLywD���)l�qvu�i��XG8R�.�Y��8>Crm��o.�yir���`��V���B�X�ƫ�bo_��IX0��S5��{CÝ�_Dn2�ä�Rf�a�๠���%��Q�#ŉ;���ӷC�e����۪�"JFm�.����ltӃz����7B��[׹kU.ܔ����2��̑²���F��4gG��Wbf(���_IhG
�� �4�E���̌!M�c�H�;�7��^wb�6Q����[�;P��<�]rv�����\�yB8��Gb�%Z�. #�ȯ�wm{�i;:d�w����1v�u���!����|ޚ{�g�v��b$p�t�q�رY�wH4!�u��N��f����*5�VYW,SG	��ͯ��/hz�s��Ϊk�2Z�M���b�O�G��G5��s�tɖV�t�
)P��z�݅j���OMkh��ȴ^��s�HJ1�
�i����ظ�K>��^EǨ�}ׯm� �1����r��]�Β*���@������`�3i�s]�Z�\,.���`�Z�]�f����b���w�M|UN�1�y6q;�4����w-OE��i��k�7C�_a��~�f�?����W�GwEM�{��)��SC֘��fn�Y�g�9�h܈���q"��Q}�C�Ӄ3��ub�7~n���G�DG�WU�g���[�P���A�t�5=��!O���q-y�yu�Ǡq�#��;�}�����Yb�͸a�')�R�œ4ΙY�lA<;%�'d��������{u;���-��G�����^���Yi�n�u���@�u��R������Ğiw)��	�z��xa�np�5p�y�!Sg�OS�t�:��DP�&qF;Oa�õM�C�fuqv.��6qljV�N�H����ӭЭ�0����(+�e�Wq��i5�2����Ĵ��ƭ�5^��(Nv��A��4 0�\,݅Nuk�6����Χ�x;�|'v���%���9v��8�;�sf�O�VN
%S{u2՜`च6��z�۹j��t'�s��{���a]؂q��N�M�&�p�3y�X�>3v�:;Yj^��9qn�o<zzC5�S4��bo���(:�;V��{�6�{���=�aŌf鼹���A��a�Z.vwWgf�W.��a=�)L���EPS)#x-��À�]�V�aj��u�Fv�� �v<=�bL��%�(� ��%�n�P��98�7e6�*�۷�7�h�]<�9b�:u�<t��8��r�����D2<D�,��Բ�V1�C.�]����ˏ���%���s{&������� ߭ܛ�j���ɇt��ԏ����O�t�c�շ�o�m�`F�G���w��.���l�l� N�&#��C_�di�_oO�U	xV��>�|���1N�R�|͙$'O1w;>���T6"+V���n�d)���;K��D�N
��a���|F����;K�g��%������1�a�o@UӬ�H�n�F��*KD#�$����U���j�JB��FC���uQ��N>����#�Q3M�l�OVl�[^��?�圎��m��R�Zx[�DW
��Wڟ�|� �)IҎ3�y
f��R|S;�$���^�q�Z���*"�8?�����u�y%�4k>x�ꜙ����LG��f(TBꩃ_��S2������8��_~���Ghq����o�^x�V��ײ/0ײ��s�����$�=���(�^&�}�3._�G�,`̮�U@^�x5�����3j.��U�2M'����s+j�O����<{��=�?-��f��0���5�xrbv����
bC���t#�b������F�ۿX܇ww/;t��ksJ�>���?��~s�C1D��i�V�i�wy㛷�8��]��a��<G�ʹ��8��*��6���Z�0-����5�d�m�}��F�9������/����
�x��=:�o�O�X����[��V���[
((��F��EOK����*e������
?�ƀ����M1~��������gi'���A�F��.���~�����H�~+i�ъH�A�NW�4�eڿ_d�Ȩ����/f_�����_د�4A{��R���On�����vj���ʙ��(�F���u�D����5�����;.)�Fc�B���d���N�#�w�z{Xȇ�=�Y~-�E��7^�$�;�F�x��/�a�ў��駒OwՎ���N{V��S��$P<|�,J���q=�?[d��~�$��7��<^�\{͖x]#��!ZwIBq�'a�wX������*�jO�[��73�:!�V�zW�<��^��dv���Gzm_�u<K�^�7�#g֢+ C���W��޹�������О�R:�y�%i�k��ou���nW�z�Ӊ�`��t��'�m[#މI�I��E�K2�6"&sg}��Ң�n*�A㯮k�~�����9����f�Pm����ź9�F/+z{���H�^��ճs2�y�!�o��_x5���-���˱���o��%��h�����&��^:���?����ښ��?�zCu�������_tM��=���M�?g�������C�r�f���p��wJ���yi*f�&*W����u~|��/�}S2� ��N��C	�/�e��6N�������\|�߁�7gbQg��z���ug!�8�����}���茞�=%���E}]>�'_+��~���q��c��x�Q^�
��J~��c���(�2���U�ZP7Y���}����X<�_�r��J�{���KV��|�)��!����<ZX�q�f���b�o����UX����;m�D���c���}�C?#s��c��g���r_t�{�3�đ�x���m�֥ۥ�_�Nqk�O����_�O�y]i���j@��r�]~���}�̰�d�D��0��Y$�s�h��l��;�;�n��i�ɓ ޛx�����y$�4�k�o<����l�I&��OvJm3��l������h���Y�wC����ǹ��>�D�Y��I�n^�:k��}.sQt�VI��Y*���ϼW,"�ZO�il+�175�$��A���Q�\FZ@�'�Q�N��t�+�1Vj9�D�_�~&ny�=�3��ߦ�x�|I'��e��X����૜�Mkq�2�����!��Ua�[�[���q)ֺ�D���Q�:\�)�<�u ��e��������a����?5��<4�H��*�"	�aT�!H�S@JJ "�(	B� �B��yJ�J ��C���/ A�(% �R(4�� %���"% ���H"������䠉@��AH� �*�H	@�P RR�� +@�@/ �B+�y  rC� 4�r �%%�J�(�H	B*Ѝ  � �����B4��hEZE���ZR����Fe�w/�>Is�S'�#�x�T7���\۠�5ǣҕ#�Ē�I�l����߆,��^xF��N
\K�5b�i348�m�soBč�P@���t��fb\a	��ly���D��ދ�ej�@IIv�n�W]�<&����F����+�;�;���!���A:�%3Nk��7_z;��2.h�W��'��r��w�kCLl��|n��5g[*a���*��Ė��Щ�-da#��Ś�x]��<Qw�_��f�p���J/}=׺����cD�����L�.�c�˚�������i5|NV��M��UD��y�.6����7V-�~N�
�4/L��؈��_�A�j�at|a�A	ʜ�=N|�μ���w;����b~��l��ViF�^��ً�҉:4�0�Q
#�()������I� ����ze���������gO	�׼2��Ru�a�"Lu'�d �y�:dgZ�[Tn�|t�f�KFE�Y�=8,��k�y�_9��T�w�t��.�L�	x�*+\������s�z��x(�~����T}�M���1z)�bųDnW���*�'$hNn9�n%��wka�LׇL�[3[ܐ��3|�n,��}��G�LY���,��ᙊ�����H��f;7�'8y���R� 03��z)�1ٌ�K�3j�{8��jIu��utך�sC�a�W ����O6/����T,��q[���N-h��R��������i�7F�����mֹ���(��[�p\�:��:+��`4N��&�,! B`��8��/=~����fmȃ�:]iI�I�#D�N�%�0�jn({������C����I>M�Y��A%&���[N���+��L�@EO����ӰE �?���?��
����������o���!�y~��xs�u�����~�|�Ч����@��ע���g#;��㝋F�v������К��ϼ�J����J��^�r*hfE Ve�cѯ�&�g�rch5N*z��YZ�mK�g7׼�3ݚ���*~]�u~�8=���q��o.`ܧ�<>��Ǻ4t^��Q*���v���9������ )�۬A�TP}wǍ#���N>ʗ��=c|��.>i�`o9	S���,�������g'_ �]���_u������ܖ{	���RS���nի���{��^ܙ��O�&��N�*2oSz<��m����U��p�A[�v����,V��N�	\���V�����|����Lp�\���g�^�^�{<W<|��;��-�}�eb}�)B��_�V��#�p�[�wnh���E�Z�K�ش��c��9�����W�1�%5��/,��1�ќ�z��9�_�'���f)]�m'&y��B�9w�����6��/��6���7�<���Os@�t=���>�wNg���f�����[�ׇ[˘x����u��~��:�C����]u�]~::뮺�:�N�뮽��~�^�?_������_��㮺��]u�]u��������뮺뮺�tu�]u�]u��:뮺�:�N�뮺�뮺�뮺믎��n��N�뮺㮽:����]u�룮�뮺뮺:뮺뮺�u�u�]u�uק]u�]|u��;��,�Ϩ���^�*��:�|�+9w�ݷ��/o�a
E��A�>�8�P�x2U\���|G��^zk�n�Y87	~X�]����P
�Ot�R<l�wɍY����B���g���m�x�5S4��G�/�xA��V����;;݅2N�t����x^���y�/;=|l�,���i�!^��^�V�=#>� �<�x��v.x�_��hm���i�oe�jVC����MW:{��s���n��{d�J���5�t�>*�3<>�f��^�����w��l)�bߟ���k5�O=;�W8�A���ͫ��b�QK۽�J徿NӜǩ��K&Q���	��2{�=�'	��w�}ō�W�y�K����BC���N�w�w���pk^��+>L\<׎�\{���2K��a]��v��w=��^����ǥ{Of*&B�V�~����|��/��<]�H��g�X��,��tF@�w��7�^u�v���2_}��ȿ��R������e7�팏-��d�� ����o�� ���s����1h�g����g�����ݘ�@��W：�Ӷ�;���*�os�������7+ØN/�4X��ϕ����,��LZ�]u�]u�u�]{u�]u���]u�]u��u�]u���~�?_������]u׷]u�]|u��]|u�������]u��]u�\u�u�]u�]~�:뮺뮺�u�u�]u�_����]u�]q�]zu�]u��]u׷]u�Ƿ�]u�\u�u�]u�]~�:뮺뮺룮�뮺��Y�]u�]w��*�[�v.��xnw�}��8��E�jљ��b�=ffaw����Jz'L �U6�,�r!���O�2g���e�>�{2Ͼk���:�{����W���9���2B����&*nY��Y��1(��b.d�d�	3k�w/�c�Wfhؒ�(�����32,K6%���Y�={�����o��y��wG�fg>��oa����5�~qMjM.
�l�4��M}��↿t�R$��3�f}��ٶ�� ���U�}�u����@���42n�H*�f��`�N+�=�/�o���f42H5��,gG}��>O���x��b:ܞ>��yq Iui���qxu�����N28ڻ9��Yw&Fܖ�^rǯ7�-I);Kfc��~��(q��ł�%�̨��'������R���}z���i����L�4]�Ā 0�� ���j���iM�����|���TT^y����f.Ɩ������sSʴɼ�r�~�>�����;�@��7����+�.eA���k�]�dp"�m,�3a(/W`�fh!�s�8A�}0|�^a�Ȥ�{0\G� �iN� =�4g#眔;�^�q���O$���[���"��z�4v�����>����>���Fڻ33�_b·�s��Z�O�f���C��w��s��c�;�n���0��c��A�w��}C����s��#��\�>����cW�{}q�������PWۿgv�;�'7��b��I�e��(�7q���<� �#1���>"=eX���t�<�m{Ni�K�����:�u��3�>x��������_��뮿C]u�]|u�]{u�u�]u�]~�:뮺���������~�]u�㮼u�]u��]u׷�_�u�^��u�]|u�]zu�]u�u�]u�]u��]u�]u��뮺뮺�u׎�뮺뎺�Ӯ���Ƿ]u�_u׎�뮺���Y�]u�]u��뮺뮺�tu�������j-䈇w�^,�y� xҾ�4�3>/q�צղq �{�D(�o�.,�o�[���7+�W�f�}��F�[�t.�]�$�ݿ|s�d�̞ۘ�G�F�ᑤ��4�z½��'���������f٘�2�������ۅM���y�>��]w/nN�*������}���o+���\���+�x��{	�9���ǳww�ڔҳZsZ�q57�Xyd�L�[��X$n������f�_{|��6uJ�Ժ�ږkR����fd�2�ξ�]��**߱y�Eu�Vx}��V�d����{�M��kWn��~��
�����T4���2�M�Ę}���oq�#Փ�P��-���wgg�ֿ1g�Ǚ.t��
޼��r��w��g{_��o�%�
zr�	�ν�{P�FY������}�n�p�?�C�zo-,vs�׈��l`�lgO� v�y�3Ŀ�dҾ��/���｛�#av/=[L;����ޢ�Ocf,�����3�3��#�\��r��,�g7&�P<��p	���x{�<����h��e��7ܽ5�n
r{z{����NI�z-"/Qj(���Q�N8�S�MyĀ�3������u���-ȟ��a������Y��l:��D�q�^9!�2<œt�:��ק]u�]q�5�]u�\u�^�u׎�뮺����]u�_����������뮺룮�뮺㮺��������]u�]u�]u��]tu��]u��]u㮺뮺�tu�]u�]u�G]u�]u�]tu�]u�]~:��]fu��]u׷]u�^�u�]|u�]zu�]u�u׎�뮺���Y�]u������.��:�^u�"��:G_�����:^�urF��7�v���5<���~%����(7I@��An3���4}{��`zF����_���2=��s�b��b|��G�=�n���Gjl�dç�wg��17�B�7V�����v#@|��{|�sf�r�!�>!d��>���|��O��n]=����]�;��d��x��ʽ��+��4p�½��jc�7����i|ޣM({�R{5 6�|������~ᯧ��gb۞w�֡��<U�TT���|Z�6��<���=��Z�u��͉�d�-���yo&�(�dw�dü-�ȀZ7�[1w,O뗸�ҵ��w~�9���'w�Z�Ǟ��w=!������˃���B���Ywr�{�����{Q��w�� ������){D�w���	��x�E�{�o1����g���D�*o'�-�e�`�zãG�'?s��c�;�zL��@�j�8Jby��k���͞���O��{C��u'���@
.�[��K��m^�����zfm�w��-!�_V��T��<�b���o�[�#'������tOg3'���~�e��dZ�sѨ�o��������׷]u�_C]u�^�uק]x뮺�ۮ�믎�κ뮿_����~�_��]u�]u�]u�_��������뮺뮺�u׎�뮺�뮺�뮺�뮺���x뮺뮿u�u�]u�_���뮺뮺��κ뎺�Ӯ�뮾:뮽�뮺�뮺�㮺�Ӯ�뮸���ɱ���	�E���A_�Tث�'�)�3'o[b�V�3ׁe�E��	{˂��X�78����כ�n�-܈nNZw�x��4�/a�F�!�t� �e����h��zU+�`�_E�pN�{b�>�-�,Hf��=�Bϼ(�3z>kz���S���
�֛})ݼGݶ{�X��+���`�;��nx�����6 g�X<<�Ү��aO��_�M�;TY���zݜ|@�=��7� ���{�7m��}Vw~�n�Ԩ6v�c������8~O�����op��*!��i�՞�,NF�zp�ϻ�&�j[ra��g5jj�s�{#��x~۾;���~/�F^�V}���>̐Lw ��92�:��/��s=��y�U��/G�S��4]M%���FyU���ff/{6�`�IW=	WG{y�"~������P��G}-��<��W�ؓ�=��=��io|氅ַ��Vϼ3��{�||�����Z����\�ت�5{=F�_�F����0������3��{�9�7C�մ�]s	у'
��<fbb"��U�g6E�����8{�����Ϧ���������Y�vK�p����Y����w��{�]��ӣ���뮾:뮽�:κ뮺뮺κ뮺���Y��]u��]~�_��~�_��]u�뮳��뮺뮾>>>=�::뮺뮺�u�u�]u�_����]u�_u�^�u�^�u�]u�]uק]u��]zu�^:뮺��G]fu�]u��:뮺뮿u㮺뮺㮺�뮺믎��n��{�����Nڽ=��r�v�<6���{tݞ�=	�<Y=�ٳ{iն�#��&�Ix;���#�tg������Ӆ��8{�#{ ��-�3Z}_@�K����sh=�d'.����w�;roy�HL���H�kﺬ��:��gͬ^�_]p��ڻ��g}��vx��3V����w��e���O=WJ����=�s�s��m��K��p=홷��~���`�}�k��=853��,�t��+gx�÷���6f�c���v7��g�bOsǉ���t�����y��=nr���C���ܝ��Q��h��c�4��q�k^�t��Zν9�}��w���}���wo�sɷ��V���"cp{��,��n=]�V����G�v����	��͏R�(�<��[fw�E���}���R����Ovt9�����z5��町��2�����[�<�]�=z�4f�p<����P�y�65�اk���a^j9���ޥZ��k3�_�<�}�p:���������M�Oz�Y7g<���z�������/�/a���l���q��w�t� ���9�C��{ˈΞ��w;R��ܦ�a�g�&�Ɵx��Gyj���D�Dlד���t�a�~|7�~Qս
v�p�+\o��v��e���x��ٟ�7=�w��ݻ}�����v�{�`�05l:������r{�<��B���=����o�8�1|��x��N;��fz��;g.y왵l;���峻�{���{���w���� ���Ek���ސ�+f�߸t�Ҩ>ܾO��(��/8y����{S}�^���_���H�
�mr!����@�%�\�/������lM������Z�?Oy�=γQ�D���)l��4M¢��'�7&/g1僵Y���N�%��ǵh׺E����zu\�7�ypk]s�}{�o���[�1�gԇ�e��n�Y�
bs�0g�Rc��<@م���}�b�\���Ht���3�H�L�t�5��u��Ϩ+���i�g��{��B�����x?u�w�-a��=jk$�(����[Ƀ�=�����ŤѼ=;�g3����|.Q}��T��<Q]81�˻�_ɂ�}��Ӱ�=J���Ԝ��^H�e�F+�G�/B����5�����i]ӷ7nP)��q��/7�q�ٙᘛ�t�i!��ݼ6'�v}��"$�=�+��O�`��Hߕ�2C4L�75�8.�E��F�3�����ʷۜ����_�}���طV'@E�Ӄ�)�6ߴ%���en���׸�s�����O�Ý��R�5�Z�����r��ҳ���s��$?s�m3��礣�Q��o`i�=�/wC�Q�`�;��^~��i��~��oF�c)14�&���^A�_c�Z�l�=�q��R�����OO�/s��ҿ_�b��ٖe�<;�Ǽ<^���C�\y0Y��S_{���s��sϊ��B����C�qϰ���7�w��{@� ��w�쇻���/w۱���[���Op�����o�O}�K�=ݽ�}���8�����&�t{>^�\����7��>�37}}�C^C{���ފW��O�xCٸ1���e@v��ؽujYgn�T=^y�d槴�M�N�I�u=�3W�D��z*+�0�.+�`�C��^�Q����ʯ��.��`�L#,�>�jѳp߰�Sw;ͪ1O:T�v�x�'LZ~����Un);::s=3��������v �;�Ov����Ӹɐocѝ�b�b��}�<�Ev%�4D`������;ǃ��M&x����F�nzZKl��h_����b;�E��gvWV��{��uv�$�ꋱ�R�Mw�f��=	W�vU���&������-�Z��:��6y@Z�n�ӛ�9Ò��>q,�{�{�v�����58���7a>�{�3:���Uc����:	�q�g�N�j��@�/wn��/nx6���DgJ�׼�_{�.?)� �bg�g3Ѭ���r8y.��}:�<k��nӚo����|����wL�����~GzQ�W��(D/{Uщ(7u����˒qj�᩠�w}����{q7�S�;N�[����ͭ��oQs����O���p�=�U�搏N�;�}��1���*�)�x����|=���{���12���	e�w�$1�������Gwjr͘��ދ��{[M�>,��&�L�}�����C�<���V|�dt�G;(�x_��V�.�9ᄯ4�x3��z���g��M�ǎ���9��x�ym����[PX�����+�=/����W�?�*�B����?��/����R�EQ�'�����ÿ���1ɭ�����*�y�jn�/�7PJp����6�vR�\���`/iv��)yg������h����Jh��=��&؈���ǋ�¥a,H�j�BJ���u�ɞ�7��O��'��@��>3�+�M/����.��F:���1Eu�b�J4س���4,�i����	��*�o^b^�k1o/R����X�x���[*]njj�.���=f��+�X���Җr:�ֹ�P������1B%�6,e��l�:4ݰ/P���y�χx��m������O��駵��k����6����F݌�&��G��4l�*޽�<n�fMC�㶬�hͻeݮq:�\^���m��<��\���ja�z�۱���4���;'1�g��g�ը �Z4��K:�s�ݍ�%����gCmۘ7;v�0�/�L�73�%��֍���6Y�p�Qu��0-�#z�,ݶ(%*����6T�(��8�[��x��;uAob��k�s�lz+�9�:r�]m\^���xW��NMش�X���v
UZ��]��P��p
4W=���k ��\듛`8�s7\nW����$v����9�KdڤZA3+.su�7 �m@�k���c��n㓠�>�����;F�%���l�N����؞��^{t:� (vL*��#������>���y4�m{V�Îڝ٣�ݲ7���j[dXz���vѱѲ�+��C�c�,K
�b��s���z�]��c��ݴڽ����%�F��p�Ӗ�Ve#��=nMT��\����L�*�jx�� �VkV��.Ʋ�M�T���Im��'ź�'�xDr�9���2s�k���g0c�	}�7v^ia��Q�ecKS����hV۫�E�f �HY��b׳)�L�`�ЭU�ܥ��nv*;Zx�'��wg��.����BȆ�˪���K
���1�K�.��Վ�xC�L�^�[Q�Z.��)�%on�'7G=`�gr���W����R��X#�-�m��c13.���hn�(v�m(rc`�p�p ��p�Ե�ƥ�Z.�g�xk6(���`����ʰm�6�Z��!+���kat�!Y��H�P��,�n�5��޻�+m�u���<�Շ��6�yǏk@$�;�Z�n�XM!M�56��u�|+3�m9:��3���e�Tt*�#V�&��f޼n�t�r7��ׅKG�݋˺n���b
�岖�.�g�3�lE�����x�{N�X0�<N�`��*�+V}u��V��m�Ps�v�K��n+h���d�\ot6���#���΃HG7e�j���n!�=vNݚ�c^���:����d�Z�d�#�Q�YL��N`�S&�l�2R'Eq��E�N�p���<s�%R��i�fH���F9ƛ�4flYu�xݴR�u���86�� ��rdJ�9֍�Ae�hM�噶�ˠ0H�ë+^�5�P�뭍�]h��9�c!{H�n�Jj�Tv�[;���̤A�Uv-���EM�J{t�퉊"�=��UqΧ;�@��}���.t@Z�n��usXndt��Y����eu��3͉m�2"�6�s�s�z�x�5�=(>�kA����^��[j;r&*{Jn{uY�ZpO5�'fkl�6�.���˔�[�z�t�Vn^!8;�f�s=������7&��E��zz���2�tzr8��N��r1g�4O\ܛ�mP/]\ݧ��J�q��t���u�/D�r=�vC��dC;��6��m�qA�K�����X3��-��fkk����m�Y�`�ڡ�:ٖ۷d��W	���sFj6�`W;�`Z\6��	����	��������N� �TOm\�mY��Y�U�й�$t��6m1��]l��zM��V�^ܠ��u�2�G=��3)d�XK�4cQ���m��;�UmcB�Z��e�f8�l�<-�JQ�-c�8'\���Y�׮G(WF�m�w;:�i�F�:z�=�I;8خ^�;{��z�8�]zR�ݱ��YE�u�� f1ڶ2��f�#4��eZ.ɱ�.�����k��UNG{���v���Ek��9u�vf\n��Ś�Y2�I�ҽ9���p5��y�<2�tИ��j�.��6���;���Nv=z����X.\m���ګ1�Y�:;`���f(�(��H��v���s&2�R;CM
a�ە� ;��Cv�{k0fs�ˣ��Y��ڷ�6�s��4>Sn��n����wfSMFdԲR۵�ev��Ɯ{�n�uy�T�8�N�3+���u�E��X�6�&��6a$0��^q��^\GGM�^l���jڃ]ldSrm��*�������m���e��S��T�l�@��]V�E�kX���R�m�k/[�/gg��0U�$ܧ�����ת����Nx��/F�
��W�m++-,R:ZkY1՚�f.u��Î�f�F:m�ڄ;��"�gx��9�[g��`��Q��CQ�ݻs�H�n��ر��kC��֫�q�V���׶�v^�o�����y�d�\�}n�s\�ͻe��W ��uA�*j�L�aX�[��Q�,3+syY�^��k��f�CFz��%�҉6���j���;�-��ܜ]�uHD��kv����4�2�f�j�s5�U�
J�ym�p,�c<��;0��x.��3��u!W$���ܥ�Ü�-᭱�.��h�Dܰn�Y���r�V���+ps��Q�������[p�n�)��â+�[cv1��
��`�fVr��mN��p���F��:��z�Y�hm�ڮ��������1�4�a\l��r�a���Y�p�l4�L��L�k(�h�0ͮ��9�46�c��\3űb��q�Fx#�+@n��6��Q��{G95�d�hًH�DH��1)JJۛ���UtcS���v;cs��&�����s�0�K.F1��ie���.�%4Ѭr˓�j:7�"z^�Iy�U�ݛ���\c��΋��4��l�J�V2�-v	��㬳5X���[��'6����s ��maRVhC�+,�]IG�r�y�c=t\7`�\H��05u�%����@v�&�Ҹ�yE�Qqږԉxq���[��*�`dq�RMղ��V�.�m���Y�ci���[*GQ��;$ȑ��lX�<&1�ú#��.%T�R���	��O��sT@����l� �a����ز����S�c/\�����p-�mѮ1��Ņ��M�D��B�g:m.��^�:c�����̔E��:ܼ<�[��K��U8]7g�iK�t�TRb�ݮN�6x�P9�ջj�P<���	tэm׈�i������#Ť�39H�����Vh�ZV�p��M�Yn�x��#k��(P����X�V�ع�Y�Ba&6v�a�tՇZ��l��Z.6�����lue]�76�h�[3f�@�¬-����� j����7la�
``�e��=�'j��O\����rq+�͠A7�K{UJ4m�vB�
M%�#UF��V�&��c��p�8�^6�k=�)�\�뱣B��Zi�Ε�%�y㸵kh�3s��I󷎷��AG^��#c�Z��6d�b�X�j���df����KY]�v�9P+�<������gF�ywi9"�ru�=���Y�ջ�D�WL�R,����T��-�k��<-�z��&ۮ�kfgm<������\7'>[y6�^�P{Dr�n5�F�FݹZg]�8�t��x��{k��4�®�'f��ѷ�i79��;@���te2��UcNe�n.Njp��/���km��l��� d��!ـ����N����0�EҬ[p�-�Q�k�>r>ۭ^��M����7]�bw5vG�ʩ$jnwnLڃ���q��ݳ=��W��i�d������X8�e��x���=f����Få윷����g��'D�l4�:�rn����7k6R�%��bI�x�9A���\9�b凮-�J9v=�,�Lםڮ^���0�@�M2kK�·l��Y�.��W�H�VѪp����uY[2';߭W��Шf{��Wk�]�jG���xФ[n�ZD��;b˦y�+(���R?M�Ou�ѐ���x���
P� ���۫4 �ś�F��k��ߟ>{�SB�6 ��f�)ce�fر�[����ee׳���&�u҃V��o����B�ɰ<�%�tŇ��M�R?�e9 �g@�[��ӛ��n�"�r=ך��|��|1���f\�+���\�n� �i���X��3bz����]��uSJkz
�s�6q�Y:]���ظ��2v�����r�f�R֢6�ġ�/k�6��A8.m��� L�bb�����}T��+
�U��7��J�-R4�����,<��A刘���|�A��ղ��T�[�t��16�X�s�cT���Q�ԯ����|a-��f�˵�6b:	BV���;�4� ?]�Z�G���Y�:=r%�+(����ʼjôc]��ɲ�\g���Y�a��ݶ�u��4���e�]�m���D�[�D��$'��x�(�O��1��r�RD�]fx?_����Ƿv��Ba;�:yg�V$�|b������DG�JE8��nY2q��ĒE�ʽ	ȥ^z?}fx:���믯�oooo�ERys��/ H�9!�qR�A�p�9$9 9A��d��D)Jw<�NO9���#�H��r�R%+�\�(�EuD�#�����q@��W��@s�	�8
�9� $	8N�#��!u�.q/�N��/G���3�����]}|{{{{}N��s�FF@�a w/�� ���+8�㹋	��2So�$k$N��z�"HJ�N(��Ӈ	�̆XHC��>�.S��	r�b�:�zĖ�Hأ��z�g��w���p�u��������������8G	�QҤDĥ�%��T'U蒔��k>�,�j|4���F!���>��4�{�}�z��������������wÇ �y%upc�"!����8��wÊ��T�r���wݑ�U�돏���\~<~����������:��N��p�9��q�& ��5s��N|��1��RR�~���8Yǒ�}Ύ	1E! �X���<B���/4�0�'�L��4x��|MB	���#)&� ��tNd�@���0�N��I��!�aQd����~8(��2ЂZp+L��cc74�}��{�e����y���]H�3��k}1�u�R7Yv*I�]����zݴq�KX�� ۮ�ֹ܈��<��9��pF`�vk �'������{0�0�e��c����Go=$v.:{[#<bo3ŭ�On�8WqۛWi-W�Y�,n9C�U]���� �3]�k�S
v.3���#�-I�����n]�#ˊY�@t��qɞk۪��r�s�2`��z�ƭ�m��Cw�6jz[$�l;f��!U�.3۩���v�oi��v�����8��8�-=/1����c���=�y%���|���Gu6�R��)�TU��Y��
1vȖ�.7sS���V;IrGf�7!t>��TX/�����r��u��=����k����AK�t�!ƃdt���e��ni�T��[���+`
�;)0#�J0)5�-��A[WC���eR�]2̙��u�vF��#C]�q�&����+��qi�i�!�Y�g��i��qTs�Iӎݰ[�WIH��N�|@�pN�vt���չ�^�"�]����x��[�)���s������i
���4l����Yl��v���j�9�Ǘ��D�dg�Y0�6���33����4��`�#�8M�d�[\�`Y����L`Ҡ�̱�͡�[��a����r�ݮ6�6�2��fʖ��I.HR�[�ŉ�ҳA���+i8�eY�[�0Pr:�Nֳ�<�w�ݫ҂�S؏��Ŗ]l-b+u�+�����U�N���4��ݭ�-�B��Ӈ��0�\f�+�\�\��:ɞ��p[��X���Ycn6s�gE�j�-�-��n��\�=7:z;͢�v�r�������b�n�h�jŢь��Eķ�r�-�9�Vm���������A��B�Jޤ,^y�U����,�-�KJ�(U���(ƕ,m���Ie-����Ie�%X�-+`�� ��▴�`�me���u��Q�����R��JF�Q��%)oB��m
ԅ����� �]��y�r.�A�p���y|e/+��c�+eN���KX�+XR��`��-l���*���s�y�6��6�mJ�"��ڵQ5��܆m8����-ǯ=��%��k/��T��|��Q�<�*�`�$o�׍c���]��fuQ��B	���+f���:�"D��1��D	�j������A7�C�D^��w}"�҄!<"�Ll�l�`��S$oށYܒ��h��Pc�[w;z��?�!�q�6�q���
�a�՘�g�Q������@{=�$k��5�դy@��	�u��&<e�K8a�Ġ:7W����bi�l���їb^0�nť�o�ﾾ�i�O,3Nz!�2�t���G��pN^����6V�Na�"y���=�Zﳋ�j����Wo���{���5�5��y����V�̚t�V��ע/rn�g�|��U{"^�eE�*O�`]@Ǳ�C��ʙ�wm����v�����C�_0�)%�Y�`<<���y�p0���@�K��s�7��|��`��v�B)��7 ���K���$@�K�>�/�͍�ֱ��n�e� ?�cnT�Ƃl�M[��uD(��U��7�+f�rKQ�Z�{b	;�"�O�(��ơ ���N�5�q�S�3}�erc��X?n����]���&;.�s"�W���@�}����|kZ8!h@ ��R9-Eb	q�����::���v�t �:<�kUR�߿��?~|�
(復	�p�|Sf�k;*�<>ÿ�7�a�M�k�	�g��?���'R=�Y{"w*��}�����H�0 �7|�ϙ�Vj��޴%܊lAuO"=��00?j~'/�omE{^���CD�`�ʹ�1n.|��龳���A;�ؠ��t�����ǟ�X��0��4IG�O\�1����u����8�N�`�(}���}9Q�����_?F���~�$�%�.�Ig�!5F}�,�q�	;�bI����CV��w��kh;�.j�sۿg���v�gq���k!gn_+n��,�h��)�ڑ���0�~�
��g�5do#�[�r\��Y�����^�f�ti�㴜.R���m���lKk���M{�^�5J�OK���D�����ȲDZ�B<U���z2��K_ A�H�z���[6�ڥnC{BQ���r.��o���0Þ�-�8sT��t?���-�o;���n�",7�y���(9�@��uV�ͭ���[�@ؖ  HśL�M6z�
��Ӿ�q�y�!e{_&Kue��݁��,�\�lL����=���C���wP���Y�'ä��K��Zߒ�{�bW6����'��B��5g�k��� 0 Xxۀ,�Y��k�����O(u-k�R����n �}k�wpZCE�E�	,�a��c}��>�'��4o��<L�J��C��kK�5��Ϛ�S��	���#U��T-�v�#��D��93��Y��c&�v`cRou�<��T���`�����v��y��S�ISށfk�EB�f��^������o5@A�����QS�O6�]�:��	�Э���'s4L4&�Rn��(2
.�F�Ǎ��2h�T�݁ ���8�%ɇ"A�������DBb�z<��k�4�����F�a+o5�V��H:�PJ�A��U�
��ʘ�
��|1�����J��:(0��yF�� [8��[YS[C����	�s�e���Ã��ۛ3���UΉ�?��Fv����`��v�-^>�V��,G#�4���-�"A"��U���%!Y�κ\\��?�gw��zK饤m��ց�:VՌ�K����.��$�m�t�Z�[�m�X7&�Z�MU&Q#5���ue�m�����k��1�n���vpr��=v����;x��K���Ifa��l�%=�鍈u-�(�e�j�&�H��`��g:�GUJ�z1��.�c��.T�d��eno�Ƚ�4�P��+�a��o;M��9�G�Bx��jhgT��n����C���߱A�$:��M�}L�Ě��M!�؉7;ū�<Sy\�bI�n�HʋȈt�2�L'�O�>H��w��u�o^ӯ�N�n;@"sb%�L��,�h�va�>�9�\eB��z]ÉjZ�3^� �Xɱ��F,Nҫ۟)�*�	9�MV9!Xsa�d'kPc�B+���6�mk� I6���S��׮�,���2��Ö���2d��{�F=�rC�s ]�7d���\�-5��qZ�Y���#.�p֣��7չY��}}?�k���O0���oܪ�U�D�`"���b��
Z�v���J˒KY��"��#�wM2k5@1s댳7cn,r� ��{�	�C�u�)���A�樽,��ߟl��L�9ۤ?L<'1ژ������8�K��y��0��j�T#^"�z3$C#K�0
:<�ޥ�'}�9�$G<�s��T�����'Rz��~��ٷ}���x�w��V A�I���Z�e<�DK��̝�5V�K�?��ź��̡A@A�DTl@����Vml#�[� ��I����p<�՛��mƺ%�M�S&���C�*�&�����;�ߒ$_bv+Uj�I��l�(^L^�ziD89��� {Z�1�4m��@�j�B8wm������(;�r������u���u�ʜ�!	���Tc�Ӟ?9Ȯ5�ǃ�*o���<����!4�g�x�ڶ����=O��ծ��p�Щ�$kЭ}��d��̺	$�D���� ����vI2ֆX�u�9r�7�Y|g}0h����C�C߶�a:��.�u7��\exo���o�5��6\�k������]b��R��T8E��R���f�.#D$H���Nn��d�c��<AxY.�q��W^g2Ozy�.O���{�ғ ������Y~�l[*	�,K*�3	P�A��f6���I&kci�Eh�,��1��m�MI ������<��_w�m�0�&��BvQ�']Iwn�;�������̖�&�[A	e�}O�/`�,4�F�C�I��v0ı ��(^l�9�jo^��m�W9��0^�u��`�B\�&;���C=���0_����������۹���:��w��uξ{�b�kָ�B��,%4�R�0L2p�1���Kce�\$�%V���'e;c26�-�F���@��`D�� �S��({l9���A#ZUړ��wd������쬋CL����G�σ��i�@�o������M.Jη$��;gE�y��Rw�<��{�����>~��֖qb^btK(-rT�����}�WP���\��1r�׬��{�,Pc�i�Ig�@%�f�J�K�֔�c֟��o������%W��:,�@u�T�[�\NTH����X��s�7$��۶�ăgu	�l҈Q�^;�1�����`�ʫ�z��Qa��C��Gݒ�����{i�|n����P|�(��VĴ�*.U�'{���$�=�W|��mzv��ʃ[|���6�$���J�Π&@~{[���=.�K��c�&8rj�1��]���Y%���ekx�y)C�g�V�{m{�Y���u�������9�=��P���Q���|ͺ��%44o�K;�Hs�Ϭ�����8��(�|d^B@i�=BN*��=F�a��������a:��.�zn��}�%�|�@����M�ĵZp����H:k��c(�O
dF�P`FS�,��l��@�?g����x�iLl�������⒙�tn	���&vw��m4�ۊ�v푱uq�$�0P�T�\q�96�,50M�Qy�����i�;\�닷)��̛W'<ê �3�[l3�!e�Ld�U��/[ %d�n���@��`T��+���cDѦ1MA�x�\�ve��q��Zvse��t�;��;c.Mu��
w1�3��[�C�Վ�̭kV���u����b�:�5�y�KYc�]l��	�p ���v�wHU�FG���<z�g6�{�|�y�H0h��q���aA�,rǨ(�>�mˀ��	�&m��`j�e$���ҕB��e+}��u7��5Q`x�6����]�X�������+1l�yi��ؿADB���z���ʴ�KI%�R�Dt��o2�r7Y���:�&jj��6���X�}��o��X���/���I�����{ʟlhJ4�]ŝ2,��,�$;�	�F��z��8��<D.�Y�cYf�3-��3D�h����(Ǵl����8I������Ql�\�q��k<㊉b}��|[}�˙��s��[-~|0KYp!���2I%nU���]:���5��Õ��%:��6�C�ػ�&j�m�.-��������K���������>���<;Ӝ�n�}ֹ���:�q�1!�%��Je�I>���ov�dx����{��9&A#F�=�a�N AyZ饯m�C1���/BI"'*�Hx>V�R	.�E)g݈��	P���![yF��R]����S$��؁l�%��]�+g6��z^�mQ�'���:ڪoh;�o���#��~V���ޙ�$B%�`�+��1�}1l�*ǯ{��b ���We*��E	XG��m����\[��:l�<�B�ajn���/:���)���N��C@6�/\CJ͍0g�쿢[Y*|8�糉r�ޠ-E^��it�Ou���0���5�*��!����e$Un`�/O�� ���1�ח�9Z�u��4� 0���h=���wN���P��C��%�>��G��H3�]�tܹ<��m��fȻ_b���r���xM=���/C��Ǐ�Q>�U�E��R�'���-K�Uf�&n��t����]���q����Z�f�8�Ҏ��;�H��9\>?n�=�1�gYâZ���yC��x�X�����=N<��ae��W��yur�GO��Y�y&/���ph�����j��]fn_�HA�=�F�q���c��j�����;&�n��C��ﺴ>�h���t�.�x���Q����\uŃvm׭k���|�{Н�1$Y{ ��l
�uē�Ǌ\�iFG�+���*n$�g��A���yĢX�Z�����x����>ߖw��̗�}k�w	.9fk��I�������ұ@@nw���n.���w%�ɾ �-.��r���>��شw.��2'e�\��	����XN��۾������w��z7�w��w���93�u\�﷼W������۽{���r��Z��^�X�S���^Lp��}���{ܴ��&�[�4Y�>{�.����x�v����,�gv���e�[��Ş��z�y����`;��8S{��f����d�ܻ���~p]4剌@�?��w���X�!��T�E4]�DX�mD�;�cz[z����d:R��t��*��É
��71t�P� ���t�SDS8�Z'�g�v6�L2Z8sD`��}�>��IM�^��g"���u��8w/� �D=����ǧ��q�������������ˑ5V�!�|ݸ����$��� �^GS�2G���G�����^���?:���������)Pvp�Fwγ��zo�.{�IH�^J�����w�QPur��l_^3�ѝq�������������W9����&̘� �D�LR�my�\9�w�p�r�>�_^3��~�q�<˝�sY��\�T��c �@O2��{�{��0��?/>*B"H�!���#@�1?��^3��~8��~�������������I�Q[a�jr+�A�P��&��ד��u:B�#���z>��^3��~?��>>������ʼ1���B�h�S��f����C260-� $�a1�r��G��ܜ|z�������gP�vQf)��&�i��Mķ��SŖAR6�̱����5�^Ę�:c��~ί�I~W�%��BH���Iak9$Ņ 5�R�>N��ϋ� �"Ǡ$x
�T���b����%,[�"��Hk{��O�����3��<����3�󈇞u�؟��>2t]G�G\>��Bx���������9@�8�7r�
r��/��p�,î.l[^��T�~��'�����~gBw�'$����N�=���䇜x�<��;�p�6ۭ:_�ܰ �KŜ����� ICZ�8+t��)��X�� 3��ǐ���8������N\��u��뾸_z��B`�!�s��o~|�O#���)�?=��ǐ�����&,���ZBJa_Y����+�~���K�`P���D��bw:y�J8a������ZJ&Uh�|/���|�uׇ���NG�~t�0K�zn����?7��rz��8G!8o��r>� Qr���F��TW����0vHz}�O<���w���#�C��������Ge��׆?P�>�|e�<��8@r��rϝ�|�ތQ>G�y�=���N�>3��!h������{�'�I�G��>����>���P��ҙBs�����;컮��݄�yԜ��<��a�8/pO��{�)F`.n_۽s�M�7N��o�E�bЃ��z`97Do�~v<��NA�y ����XI���	�$�����'#��Γ��矞�ܻ$鎠�L�{|!������N}���'��\������0�����;�[�Q8g�����1y�����0����։�{���f��=5�ɿ�e��e�=����!��Y1�0��	C����]y�ȉ 2!2j��Iӧ�\��,����μ��h<y�~��!�y�ߟ}����@{d������ސ=e|����p>��{�g��;6)������C$�i)�Y�m��n��Q��T�RWb�<�֤ to�����P;0�(�'^�O.�9�)ÜG��޻���G7�If����X�nfE�s�D	yA�s}��8�w���=��;�l�ͬೈK�C���b��ص�(L"�Y���.�W�0�������� �DY�j�Hy����a�
4���骷��f|�����߄��D����<�}�e �����@J�5S}��/6=U�ȀI���a��̙$Yf�c�gq��3��0�(&!U]���
)zm�kJ/��́���E�@R%ˑ%��M��+��[���l�$z� H�G����Â�BJ}1&KO-h�E���&����C��G�L�^g�3�CF�H��%c]�P
�I�A�~�[�#�p�d-_�X�p���^ǲ���׋���_K��#��1>���K|�ŭ�z-K���=�-;kwb؆���Ѥ1"ح���9�ʬt@���x,0X`��a�g�o[j�1�H���z�Z!)E}��'�����7fz���Ogkx����:ŬV�s���i��r>�[&�3��[��'X�C�^9e��G��X��*�c�&�,��]^4��q5$$S��)�6�Ò�E���m�X��Ax�XMW	k���щ�%C��lM-�Ұ���[=굠7w����J�Mn��f�(��T�5Kt!�R.⅗�4����l�Z�#�5��߫d��	��e����JB-��H^��+�I� ���R�@'�sԹ��R�����d�^ۑ"@Z$�$��n�n����-m���j�Fg�:�l�ٸ) In��j��"c�B-�V7��<w�k��[�Ӳ��͓�2w�A�h��zz[�R�o�A�,�X��I󢇻�T��54�$�:XA��.�Ф%�{�q"	��M1%�5)ף[�31�H�	z�l�ۘÄ�= �I�X� )	ZY���>��׭����% A'k���P�� �Цe�3��8
u�i}����h��51�Y��d�:���K$J]��%��)e�5�Z�\�&0 ���J�i9���v�r�F"ʉ��*�A��Hɿ;�I%�d����s�\T�_I��m��q�	�����o{ U�"eKN�&�}��ҿw{����)���N�.,������i/�<�t��š2Dw���mM���H�_zx������4{J�8�zA���6z�����X����)�.u�~�f��0��x�G3�K�_��y�Q(�o�Ȕo�3>gD��a�,��4J>Ф���.^�A����F�2E\�|SI�Ď�}S�M���1��K�]��U3�t�#�4�\�:A��;à���s�P��}Su�.y��7��3]�`��>/����d�Lq�P�����"�c�ܲ;\�@+�P�$��]�;��W�Xb�<d	$��șd�6�
���KMlt�Irŝ�nƙ�@I$oH�(�ӷ�s"vB��$-��[k/��[�e���K5M×z�V۰�.�Ct�t����q�o߻� �Z���v���� �f2D]�,&T3ͧ(O�I���$s�l����R<��Uҥ2vt��������M���Y��FB�&��(����k^�_N}LiiNĸ�������H��`���x��b�I%������æ�Ny��z7ŎuZ{�z����|g�h����D�غ�<J�}��^���z���Q����8}�b#����'�3���z����̐w���0�T�w�R�2 �5;�h��
�w�)D<�/���K���߈�����- $� ���,�de���L��<��w�c5��u��D� ���4:Q�z�wtS;��E���w���F�6�,��3�;�	 �$�޹�I '{�L�
{��&��i�э8ڵZ*��&\��{7Z{qf�Vy,B���!�Hc9����ʪ��h6@�a/Q qaw	�$X�ޘ���g�ޣ,`}A'�� �DO���A0�G�:'fA�Ycm��/���Ɓs� C[S�@6�1 [3Nol�P'�f���7���u�;��T��]ORa��L��0�v��>�F�Z`� �݉"I���A��[��t�	w�Ml7�ם�L�C ���{�$	 ��2�z�;���ܒy��B<O��O_�v[���Ŧw���k&���|2vnz�/�n���������'�^|��E��і�gb�X��p�X�1N�1�@(��&[��/$^"G��Ԗ�A �]�3lCl�f��͵��&�݄����]��{�f�x��wz��#���nEB�-UJ�P$̜��Yh�b:n�ԍ��-p���9�����ړ[@�zaݡ A�@����Gu�0��|=2�
f�8:}3�XH�$�]�ל	8U^	Kn���c1C��Ma�a�>b��}8Ņ�a'0i�6N���~�:-B:��d�C,{vbA ��D+��CPF/7_<����&SK"�gw�c�POH�=N��V䦰0@�N��&��U KW:b�w.�L�l���� �r�I����`�ѵ"H �[�,c^������ �l�5-,�ǒ=��� Q]n �Y��ڪ�]AR�y�-N��\��>^��N2e���Zo��0	���@��䂋ǻ�	���KG�?���F���s#eX(�wGpᘐ��li���ߖ����pN;�,|7B��lbY���³dֳ�X�N��ڰ�vG���v�Oc�wD��)����ΛSe�:��չ��V��4綠���SmGG�c�-��]4�j�&V�]i�0�q&ٻQ�&���ke ���As�ld�.0ᆻE�fpqv맷Ot��'=�nzN���<�Ʈ�`�n��b�Q��0Y�e��z�_K��MC�l؉vu͊�����\�[=��v��V�)/݁jN�"x��e����c�T	,.�cR,9��!ǆ���ƽn�Q�@�1��@'h����<$�c]�:Ţ'� �r��-�ޚ,'�nY��"��_����f9�wD��7�j��r\)��1��@ �1���F5�h*���nG@��nn5��bC�Cv@'�A�
�yP�Ç�T(fk��!Ґ��-LQ|�� d�|� �����9���ɓ�l GL��u�;��W��mK٘,��co�v����b����wT�-蘁�"^����lrA���Cm��^�&6������o��2릘��rJ����+����<]ŷ5��ջn�m���ږ����rIP;�����ؑ,	�ۆ-Sv��<ԧ��{��7���4�"�H���XE�EP>��쪐@#�����:G�g��U##�"㱰�xܩX��e�ew�s7�$���U�\/zK�΋5��d:��e���s)��f^K�+����9�~� ����{��*	㟝�X��'d����A ���[Ԅ��0ˋ�v�N��*�Np��<$�� G)�:� ��$�����'�;�D�Y`@�>��[�A�����$�H�t�ޭ�01a֕ "�ev�2I �bݵǷ{u�0E��bF��Mlt̐5�=��$&��ީ�}K�i {;'
=ީ~�g���0O�H?�xM�f��lS����h��=���\ĵ�����ڜ��$��>���1�=��ޓp"ڐob� �H���v� O����>��Y�:���H��͠wr�N��	Q�`|
�M2v�B�
�M����@N��SR;�,5�ࢡ��S���G����#D�\�H��,�t�ޝ�I$��B���K��\���S��"���ŅNK���]@{b7�Hz%�2=����{����K���BR���� ���iI�u���Ί,A"#��$�wQ;�ä�w������u�!��bq���4HɂY��H��_�o�R�5�1��5챘�;<�H�/=��D��p��ɥ�Ѿ��L�%1ޙ�L�X�˺ZA	 �sل����4�ޭ ��pQ$�~|�m�ѕ�%�a���KI[�e�W&K���#��[��
1��t�0a�S@�u2�� �=[���=�&H���g�\Y��qB���CK��'r�N�H��S�f�k;��~�:ld�$[ ڌM2m �{_�4D2�1�'y�ea���͕��0:r�����X@ȟL��.7�M 'Sމ�\��\�\@���CI�)�s�2�/c�Z%��""k��=1��K�=2>a�n���z|$�d�62��0�d��(�������5x{/]ezl�_+��P֞�	㦧/��ՠ���ۛ}v����R"��T<��"�pj �0�`b�֘d��O�~[D����
:�$��$�����E��m� ���`�� ��C[�[=�2�V�\���/< �CG�$��H��Z�K���@֔޸:
ǆ�4� d�
+�]���J�����OL� �d=���"s;�Af�e�>�����'��$K�C#]��I7x�
 ���v�Kc�Ô�,��0���i#7�D�$y�j�k}qZ܇f��������'c+�����^�z1� e�vE6��f�j+�^�ި�t�3�i�_=��>1�����?;�
?�;^	�'������kc|`8=���C搽�wb���2Pd�l�{�ffE�>e$	�q�=�Qt��\�����L�$�S�2�e�.�-S�1m%���gg�o:z�G����������f�*�Ȯ�U��J�c��q�^�\u~e"��{ٷ��CM&n{}vb�4�w��^(�ʙ�����'�s�>��ʅ����"���/\o�h}��]G�>���p��[���ٱo6/5�m��91s]�_z,�"u���'�E��y�HI]θ�M�W(\��������d=�g����#��Qֶ���>�� �8<��V���ڷ�B��a��);�8Mt<��iʞw��zvq~{�/�K�J�y�Fu~��<q��~Ѹ@�W{�ݙ;��A��N�c��n���?^�za7����^�=��~�{;���mڛ�P���#�1m}��)y={�
�Z}�k�3�����q�;%ͼ4�M���v��5/�� �h�7�Z��q�Y4�n��c~� r2����:7Ja�UzoQ��+�w�+���f�{
��S^W�����7�+�=y�qcw��iBN]�����`�}q�'ŏ`=�Hno7�H��eG����Sv�k�y����t]w�wcriM��k�w�QG���HZ��|e�=�;&�(ۂ��U団�1�oz�f�1�|�3���w�g�����vWE9�S���v��fI����Fw�� \Iw�b4��F?bz�e�d�,o2ZR�Y0��P|� ('d�׵z������3���x�8���-�ѣE9I����icS���c�|�^���4���/~?���`Wv�~��(����>]6����P �0DP�2]J��1�����fW���gB�~_��_^�u�=e%r�c�I믽��ƢE���@�a�^��������Lk�hü�'��~j|Q����ٝj���I�'� �U%��~,���
E�!$�cmB
փ �J�Ě�Y�w=ǃ��|~?zu���>>=���w��}��:��� v%,1�fUd�<bˋ""�eϷzY�v�����g��㮺����q�w�8��]ē�i#��1��e05ԫa¦W�c�ܶ�	�HB\�
��G����<}g��������q��{��S@�H:�åaot+����D���=rg���f4&5�Z5��� 1:�'���9;��׏>��?]zu���>>=w�By��mi	���W�"I��dEBA%�f�w�4%k��/.Gw9�ιgwG�s��׏>��:������q����Ys��κ(�כּ'��b���`�K�|��^%E�ql�0+��R�3�йz>�]x���8�������q��U�CFd�l�9wRf*8��9#�)1ѱ�ŕ���\!��ف�h3fy�48���Bu�Xy�5���|8x��U��@�~	L�C��4�à_{�ٝ|��cǟ6��gb���h�*�E�1��Wy �hW�0������#��f'�=yR��倾S(�M�`cm&e��.-�6��m%�qS,q-��r�r�l�Hl�<t�=�G=1Vٺ^�8�7f�+��Q6�[9x���ڜ�^���m�����Ln�=�zNnlr.L�5��Q���	wh�(�*8X�Ȃ�띜��X��M�f��3��D��d�\�tW�t���xYl�
��7Y�[�a��;W6<ܐ�/d��t���l�c�N����9�î:�\�P�Θ|����;��y�a��W�z6W\r���w��ظ�t%��Ժ55���偵�]�zy+���N'#Wa[�4�t�wV�0+�m�f�����p��\#�n��'*��u� �n�L���:�pP����tuj��WAeBi�������<���Y5E%"��r�K{i�JU�Jx��Ҩ����s�-������h��W��lq�mPg���)���<��x��6�r%�Yi�"ws�����k�h�Y�x�9H�.���;Yۓ�u+�g�gC����7�0��U�#/�KnLx1{K��tu�z���W4��VU 1F��7$e�2u����a�k�.2�����fɁ9��R�=���xKe��b݄f��k���1��<]���3Yt6v��{m"�H�p�۞VoG+�7�k6:�.u����V.��{-lZ��b����uӻ;��j�Ҝ�-\;>5=\>�n��z.�\��n�+�@�����S�#;��H&�Vm;�XG��bg����z.��ۙ�3�R�j�mp*�u���]&-�gCԒ��<m&=�n��nN��������(��t;��Qdqu�����ML�tMQ�@��]FՂ-[�`�ѲS2�Iu�����Ǧͬ��a,�3M4�K��u��N-�Nwk,�5�ZrƤ���VO��c�Kg!����ǋ�h�8�()��<Z��X�<=���ntt�"��qn�H����'X�Y��FWY��\L��d��i]�oU�jA�ٷz0���X�xNga�rJ`ەr�M��ۓ�#b2����˺���h�#��Ōb6�Nm�٥�yn�c��gs%�g�⥛��ϋ�ݱ�K�����[W�\��H�P:�۪�M��^����1M��Ľ�t��NT�'bsvCpX�nz�DtC�Hv�����߿!����{��'����ˋX����kU[ <.	�^Yb&-�� C5���O�u� �3t�!�H���y���MUםJN�H 	m��q�"�߫��b�.��mg�яz&'a�
HH�A P;f�
!�G�6���"@Ɔv�#��4f ���Vv��7��
$���3��W����D�u^E�$��xxt�,��lci��,��LH`	,=ux�@�(�`n��!��}l<Oz}2��R�=x�Q��W������E̻ � ��xgeu�{��l�	���-#LZ����;J$�����\����[7]��1�Ծ]^���)��)pV�&�lK��Ŧe���A�˖v|��!}:z�#�S-��/2o���+����$����v=���������3�x�A�L� R>ɉ-#����AA���d~{ S�Tk:��LI�r��O���{�a�(�e��o�S^,�)����etxT��	VG�E�PGM��ZL]�J!`�����g�>y��@��{!���R�C	��a���v�NO�vH�}���%�7�>u>4w��I�_ZNC�0J�2�ޢ�ɉԏf;1��(��Q�b�:%2@��O1C��K.�Ã��
�sTO�k��ee�ܢ�l-�hbt��K d���$����vߧ�83t0�I=�"@������;�y��Rfb������Xv��x+��1�'�(�EX$1@���,H������g�s̆ H�̼7�A:�m��X�W�h�e���vh�6�-;-K���m [�x}�ȝ�%��C�`��٤�9�b�!L�0w�L�}��{b^�;�1�=TX`9�������@#�^�I�;�w���v��@P%�z�Q�Yֶ�ȉk� �������@B��ޕ^�����)�}�r	AA��A$݂ 4�D�"ƶ�%�p4ǳ-�rP�����QR9�y�k��Y�|&Og��˺���{��:Xǜ�����/u��|U�N�	�DѬ�a�`q�Xp��D�ф!�+��a��;��ac��y���E?���`@6�>��L�jH���I�x��S@�rc�5FĮ�N�aL�藂��L����A �w��n|��.���	=�A \��j0ˤ��t�\h"l?5G�w2���25�@�`r��A��zd�Y�H���nRfr���N�k�晛��ʷ8�Ϡ����c<P��5K]�����������z|���	b�)b�Э�b܉)��;�y���ι�Ϲ��O�'a�;N�
J��a�i��wpb����s Ej��xQ�� ���@c�Ic{ksϣs�k 25ñz�$�K�w֫�6g�/2DL�LS�WH��C�	�q �lP��$�@-�Pޙ`�Kdu�܂`;��fr�����N��U�!� �@��D�d��,H��$�b����I��J�eڎ��Y榠�㐚��hN��w����(X�?=�g���<t�V,�B^�x8���V4�$K��+�Pʂs��r��@?FA������<��$82��� �@� ���t~�� �4�Ǽ��w��R+�<���|�	�z��է-lB ��L�1D2`���I ��v���.@�X���S?f�4l.)F����ѣ��^�T'n�<\:�]J
�mho�<��֭��#;浭	��Ȓ���,%��Q稃�T�E���,I�hf`#��d` ����^N���@���&�ر9@<gT� �#̐���	%� ��$�D�*�����3�G��Pt��1@��w��'�$�+��{�j�zg=3ӑ�2&�z��b� q����K�F��=��Ł��EwK�;�)�跻f���4�^:@�c	w�e@a��y��xl���,�\<�Gud4��u�ۀ`:@y�'p.a�b���h�&3��Yp�@=��2K@�;1i�����ן���c�:�yXt�5eO�(���_od{~�V�O�ʤW;�P��5�X������-z�1�D	��w��^;Vn��13�j���;u����G����G��9^�-���f%�X,X`px���C/p�9+ł� K!��)��c�M��!�_���ǝ���a��ġ��b���;�Ք�lbk<<�qt���]���sò��X]s
B��EV4�2��pW&<�)��4q���;��������r�7��=sF��v6�N
��<s���VX�{;-�����8�ݯI�Zۜ��Û���JəX�vԵ�\����fBiR�ӹ�[���f.4��mZ�}����u��֦�J���[��՝�ʏu.Sť��k��}�>�8)*i�/?�s^\�1 �"ŉ�DC[-g� @LB �~��e�N��ž��� �F�H�1%�u�&A�Z�9P�C��c�f@�A�إNf�������e�%�2@�gvt����oL�HO/>�
 0a�X�7&���wED�njl��E�>Kg�"G� �2Lnq���m��sU I�DAi�v-��bZ�li�{0:����Y����D	�r��3��,@&-~�ng<O�:<4�3� G�A6�}�����X�D�#�S ,�|�'bT�R3�\�\+��Sfa3�!�	�ɒ���� �׻`��s_y�<1��6	�R��4 �۟U�-����zN|m�]�[Z��E�z�t�,o߾~����"���9��8���H�I��'Z �L���C�]-h�0M<� �A>�t���x��w��R)�LE�[LUm��[��x�f��*G������?Bzg�)���>�%���=��n·���S�rƠ�%9��Wh��:��iAH��u�Q ����4��|���:ξs���r� �80�0�/�82(��L��W�|�J��~�~�4_�~�w� @�3��*��W�a��{��d����C�"�x-�3�L���܉�A��a��d{���h"<�	,Ia����zd�	̳|J�I�y3G[�t/x�/y�Lͬ�,��uİb -��2BH���楚.4�}y�	?9�K[�������J�o6�=̶��ҙ&�(��a�@�*�:�^�1���H �wCws��s,��ۯ��?v24�S���k66}�Z��stY��K����(��
I8u�'�'@�擕3� Gy��@>��a H��g�;bEEf;�2�y��{g�'[Պ���%���< ��@p��K7}��t\HT�q�7=��q�q�#{��7~<y{��n�J�[7�z8�M[��!�	U @����@ �[�7�� t<xY�.���5+��!woFU!T$��s��Խ�I������y�C�@�q�~����y�@���R���I���7�#�0����aB�)����"'R��|����4����R������@�[����WZ�9�ly����>wl�e����v�$&@ �YǮ�u�J��i�7C@p-�Y��$!���
�	�0�,����IbL5�uQڮA�l��x�mϻ��x��_��i��.E��~D�e=g��i�H3ј�PA0]ʎڃf7P[Mu���B�69��Ԭt�F����{�����:��$	;��C��F� ��^���n�Ƿ��H���R�A2ٹxR)�{bT��Y��$�@���� [	ngɫR� ���\�5���#<����bB�D��L13� �����]s���g;  M��H�}�x�@u��d�� ��lm���	�2΁�2pE������-@"�@ @-��,%���U�g.�JG�������U<�y�+ d7��»���n��X�_r�S�+_�������N�?j�ܳ�NHq�n���5aO��Jl��l���{O�I��[p�Ow�]8��)�A����u\;=�?E�B�FA��¿��t2�܏�����HPI! �����-~�u�in�;�s
xu�x�-��D� �  o'���{�'uy�0
3|�K�-d�t�I�Z�� �T�S_�v��0�턮v�aa�=[�.ݷ���8\�szejW#v�����)daf��{�޿@>e��@$H9�y�[  "��� ���	j�㗅Ј��g�
>��i`��y��7��yS����&�j���؏s�4�w1�.f����	YCP)8{bT�� ~��� K��nb[���,ښ6�5^8�@��vp=��֦D	]=,�@;��{-f�P�E�*����k3k3@4�%���$ X]; C%�y�I�M츓	跀��y,*r�+�� �0혹`A�j�� ����^�����뫐$��I\�0���av�v�_h@o���K������n�=ڵ`m���z3�`�{�.��(Ŝ%�ɼ�@�/R~_�N����������fq9κ�w��u��~������B�x0�%�<��	��I���O��ffmLK2���.��U����qb��z3��ݺ��i3�s�-!�vyxNY�i�fk�2�Yz�`�T�ΰ��gV�֮xFwY��q�\�I<n��ٷ;��꺻3��#�=���7M�0Wn�6�q��^i�f2靦{-�i��re�v��c�vݸ�Ͷ�M�L��Q ��^�9~Iv�΅p���m�jsY�gFY��ARh��K��4מ{��@��@�y�v�� @ ��XSv�0���e��g/�/Õ�a���j$d�V\�5�O��J[Y�����e1>ק���<�H	�m�L�!�cm�E�V];�;7�U{U�QÇx��|�T^̖��N=��@$s^�~�V�+�k�&bI����|�v<2�[���)8��LǦ�D�3�����"!  ��D��+;�[HM�-�=,�e���|���f��,X��]��������ج%���B<�x�"U�<�l� 5��`wI7v��{`$��̐	9���6���镆<���x�z�S���s�[ֺۋYl]�X���Yx��$9��E�>��\w��R4 ^z�Xc&�/�.�	m�t&�)4q�)}��4���Gy�U������������ 25��8�%����K��FpԦPo�/)�^�+��rv^������Ƽ�����e'q;n|
~Ćv8��Ċ����9�����Y�a��Ix2���*�80+�x<RT����?<�����"��z�RaR��!(�V�W�@G�i���k�3�I����>��X^����Z���׽��0�1"Y ��`AvA F�tλ�M��VQ]ü{���#!���;�k\bi��q3 52>�ِ@��AOD5@�~������D�;�cS%p
$��C;�bA ;y�qtL���^�B�� {�@ k ���'��톣/�[�x���<J��«ilUYvB����l;�9wnJ��u΢r���J5hH�����Y������x��@���`@6z|@�lwz},T�@aj��ka��/�x%4Nac��' g���'�5�2I � v�L��S=�g��z�l��ED�}o�y"���9�<����I�;��x��* �;6���y�9��C�o��;sU˩D������LIZx�}���T��}�0?z˾��z�����+f��/?r���6ǳ�69�x;S|=��z|L����s޽��]�`r���l�qS�{l9�M�G��Z�/+��%N�x�y��0�~՞�j�v�����<��N� J�SpL;�qMk=v��~��c�>��������^��t!b�O��gz�`	t�Sd��}��y553������(��'��-Q{o��1�pv����N��"�F�9�ƳW��/�d�%���{W����]�����w�97��4�x��m)RD�y05����g�6y���Ӈ�y�I{W���܄׫�sۼ���ۧł��鯲)����C^��:�*��cs�V�g���H��O��9w��	V�� -Cf��>q����Gy�o�D�������>�=��7ڄ�A�W���v9�&�n���7�Oǉ��Λ1w�����o�{��я��$7��~��\\7������mNr�vɞ1'b�}�ؙ��L��ټ]��;}5���ٽ�}�MuwVmh.oO�����9 ,��d��ݩ�~򦅟�c)5���/���7vHaXa�A<�5�m�b�ꮚ�}֑����������B�Z�������n?i6�����6�݉�1]�y�@jΊ�~V�d��WkWL������/f�C�z���f������ck}
���O+ā���-�р 2	"\Ä�K?�[@�1D
 ��r�6���#q�q�|���_f߳0rC�E��a	ʟ�Z,�mN�'yU���pRX'��!�Y��{�q��q��o��q�Ǯ̚��G$�x��$���V���T�
���܌)�;����y���q��u�����>9�D�u�����9Cli*s�ČP�q�K	�8:$&eOY��������:�~?]{}|~8㏏<˜�뜹Q����	��~.���RAyH@Q�9S�}�����q���~�}}{}|~8�g#�+�,H�N!9"�$` �DHC��6X(BS)V|ﳾ��;�q�Y��~������q����:�9˾@�||�r)��6���`O=�GE$��~�
C����ޏ��~�g�u�믯����q���R �B�e�	�������"�$@����	219��g�)%rp$�Џ@�\\�[����Y%#�K>��'N�z�dy��ހt�T���S�X�H�b�"����J���)�Ó���t�	98!�pB��H@b�� t�e�����a ����E�r��G�+�2�܈pa �9%(S����P<Ex	*	�����?^zݳ�^�kx 	,@_O�--yʼ���`w��ޝ���*<�2�M��$�XU��Đ&�wz��v��9��@`�ޒ��$5�
�� ���$��e����$�Y�v�Ͻn�FQW�G �K�t��H=���!;�2�.�M�! Ͼ$�-�68eP��an���.f��I[t�(u�8�d�7Ui���s;%Q��ŝ��4Ă<��	�$L@~�1g�Ew�� B�� H {��B'y��%$�@sK��_��Ů}w�M}�6=>� �u� �1.�cϗ2@2�wCbÝ�o:��ۤ���/�:x���$el�kS-�?�@Y�4~f���G51G2e�$gt7��q�LA��������#���[E�H,(���$	-��`,Ev�Tz|LK�vL���}P���s�8m���U��{غ��c�=�{=��]>����:���L���b;�5�wu�k����� ��C��� ���<�Z�e3>�v��$��f'xx�D����󰂙��X�K��p{��q3 �@%����X�%���h#C�U1զhz�!����~�mJd��b���7K0���od�q71�-v	m�A��b<���U���K�����c�L%2
��2��J���}F���A_e�I�)�l �\@�@P�챨aw���������e�d�#�����T��jH|��-';�%��	M�w}~����"u���z9+��1>}1x{�4���]\f�c��j6%s�7�X�n���	��bĐ��������e;���b�b$��^�%��	���y<3 [y�
Y!���@3�v�1Ɉ!�Ԏk��i��$��d��"0 q= �Lb�D�^Lsg����i���_˿�y�Kڏ����������{؅���g�|wO�-�<x�g��ǵ~k��ֲ,�i�b�L,x}i���S���𐗡�#��'�&�mW�l(L��:������2��"0*C*$0�C �����R$�ޱ��`���if��ݫ	��qf��bE�1\=Hks�Y3�r��8n��U#��V��{�n=x�+�wk4�*5�;I�l�:���3�q�uE�)�j�k��P�a3%�E�s���E Y����u�hvH�"Is�Cu�fXEY�Vݽ��3ˌq��m,��U���ѭ���X��)�[���m<VCn� o`���J���5�2�A�S�}���~rYlesK�Z嘿�׉%3�ͨ���X�B �NK͞��=2�@�4�ȋ�I�Ṃ!�D9O^$�E��=T��g��r�s'E�yShx��A����6��3�V2`���횇�����D1���^��x�Ub�����%�'��֋�-I��b����e����p<�ı��:��H,��-^ S���;m��77���3����q��&����ı$
�\ �(��Eڻ���y������A2W��������1 �)��r��:����H:��\�j@c��j��l�H-z��2�y�'�c��B~�ϑpYc�N���N�2tq�r�1u��H�w@�^�Ny��!C��x�]T��9��C8Z�����9�=����ʉ�LQ�܅��y'�P�z�}f�Qh���g���;����J;������x���;3os=��>����<2oY���*��T��S���P�<+%�J�!
E����C�B?���0+�T82��p�{D!�PȔ��ʏ@��`Z�Apv3��jD�����-{��Ɋ�w���}o�}b!�D:O���3�!�J Z���T�c�ax��i$	���H�,����Ke���0�!]��D@1p��ahP(�!fYGMBbŊ�d�4�-戨v�Ń�u#;f.EyM$^C�c�U63B��3�\9N��:�A���_G:j�Gho7�l�n`�Y �WcHr �C��^d�j�*�e��111P�yϼ3�
 �I�W��i�d�ɉϠ�oM�H,H���.�[��R�w{m���`��~<�������4�u9,v*��X�e4U�em�K��JW$u�XшZW�>�(U���y�#�X7�d�Y�ΟD`9m ;��}0�u�Z����ׁZ٭��I�:�Z��)�͊OF5���q��A�$w�&A����ܜC �F���(�,>j�I��D91"��4S�-b�vdH ��ؾ)��`��^��*�C޿���w����%�?v�p���}�;gu˝�ɚ3|���_K�þ\?c��ߧG}u˟�!�0�r+��]��"�2�C��0fjl���A7��I�s�5h��̳�"'�W�!X1��h���/y�{H�neJ]NײD��K�9�H�Gd���V�`�x����v~��0'�1���U��V�a��)nd��$�����́��f�~� g�nj�QW�c�ݪ3��ުܼ�n؞��\�����NV��q_����er�.���;��^���{o`K�t�L1[5.{�5���l��:$��կ�bd)��>�;���f���!e�dێ�$�-��6��+^�̆/C)��r���j�ĀAv|�\a����fZ�������A�!��Uo��x��h>�ؓL� �GL�3y{x1LU� E)�ͷ���z��@�SA��8�2C�2I�Vv����4�+��߱�!@vbE�I�*��]�#����'��_Wqa��Y˼A��\mO7�c�e|�{yߐ�$�,g�����I~X$��EdF?eG� rx0��R��������?~|��λ觊�|^�dIaM�|��h��S@�{�I.�.���b���~0^�_�������q�~��&Bƞ���tv��,zW�s����[e^n�+�D�U}�}����ޗ8��ǽ[1]���G}��S�~��"��7��.�2(`�����o����r�	��o�#��4��?q{�$y��OQ-�U�2 {z�d��>�_W|���!����d*��oa�p+�������Pz�V��꙼c��o2	��L���q!��(��j#<�Y�
�fH%���Q6ٝң�{����C$�zCI֧�8��N ��\���M�oM���3��k>�Ȗb�#�d|��=��Bu1���:�\xV}�oN��y{���w��r^�0��0Wx��k��hAwo5�N['Lњ�~S?�{�o�<*jWe�I�ɹ����Bԡ%���d��s�����P?FU����A80)��R�NB'D9
��X�@�Sz[|s� ,c^��G7x��{��mD��01Z0�Ҳ��uKYzˍB��N�0��cغ�iV&���/2�;jF�4�����eĭu#��as��\���c����v��ζ��p��eLy�ݘ�OmWO^.b�Pu��x��iJ�"m�vh*�ц�Z�V5����c�l���6���-�-e���d�sX�ā�!����B��\@ 7�w�Ĳ�Tr��x�NvjD�	�۷��}�'r� V��"+u{��a��}�I�U��j
YH�n=��]\C�ށf@:�����o�q޽"OtZWũ����k��}�Y�l�Ԏp7�$������my����$�����!B������>�����"�E6Ų��q�g{'ȂAڎ/���;��6�%^@��uN��� �<:7}�3-M�b&Z!l�*"��f���P�AV��v�
�v��֣��p�A	 h��������iՖ�;/;�&��<���������%�HA��]�8�xNH�*\@${��Y�,N�s��K݄��WC��"=W�&<H5�31�<"����8{=Fd�D����g��d�7n^L�Nϧ��z�%?E߽7� ��F9�,�
sR��F��}󾯿3w��.s�yE������+�(pdB>�'�(�(Y�%����S 'o�D�d��}"����ʚ�M�v�>d+�<P�HD���ْG�7WŢ���j�3:�c͈�ll�%���L�uͥ�F"r��z�G8��g-��aa�r����bA$��ْIl�WU�����ښ�Zdw7���w�b
��y�=0-�췃Kr�C�Mec�H��$�vr�A��絛Z�}������z� ��%��{lɮW����g��s=/��q�ݠ:�s�S�׾���p�a���{5H$���D��$��� �F��+��ؙ7�z%�����o[ۤ�D$P0��%�����OӢ��$	��Ζ!*�Z�/�tQh�vo�Y����xEw�};2!���淞�LA����v�w�"�ߞ��>?N{}�x���/��Π/��w��#!A�gbS�^X}�
e8X+LJ.vg��%B��A!�?`�C �ʈv����Ϗ��[;��$M�}p ����"		H��5*�}t�-��� lF���H.=� d�ێ��!=�:o��%{�gYw}�lAO4�YY/ &{������� ���JiC�W� &2ҁ��,W�����_D�
�����<�Ͷ�m%ni�e#M����n���h*N���kB�����-�gkDM�F���"1��X��tuw�,���̂H��%�]�!g�����vf�2	=׉�]{��;ĉ$U㰃>�AH1�=ı���i�T�s-�k�� � �^|��SA���,S\�Eĭ�}��}�����,���!{���&;�
��7T1��	��$h�����B���(���� <A��C�����n��>�Ȳ�9�*.��{P)c�&}���W7D��{v|�1�;�����|�>|��}�u�s�-+�T!�@�d���xA����x2�Y�1E����W�~�f�)X��)�F;;��eș��윌��`� F�SUԉ[��92 <;��w�y�穏�1 hB�-,�T�T��fX�klj�����5b%RT��c� C���?jvԄ'��#��܈$n�q$�*w�d��f����6�wK���v�m�H5�_gcBw���{�-�2��T����Au�O����<��@�*g[�3�i�2d�Q>�A�z�%{ޕ-���1ѹd+�!0�U{ffH��L� Y&�S��;�� ��h�&�u��S"H3���)nnpB���y�]�����f��<pՐu���!�@��wZ�$���\i�E�j�8F�ݽT	k�z7,<A0!�.�A*�O�D�(up�8a��w��5"a��@�(����Ru30`g�)oL:횛��%�.(�I�0=�7�&��Dڥ����������+�ԍ��}$ �3����x��%ٺ�6��}��<�1s�pB�\�{7H{n�ӏ�{��'��]q�{�:a��X���÷�{�G}�$�ɠzc�^0���?wp'��Np0gP�ݙ�g7	�9��L�B��@q���z-�G�̣��ՕN�\��ԍU�q!�X��k�n,6+}�y�����=gR�����"k��nS�;�3�UG�u���|��Y2�G)�?q�,�/�08��3W�B���͎�3Qw�$:�D;`�q�o������ ����1����>+�ۯ[Ch��8�}����/cX��zoyz��'	�^>��J���f�ѝ��Lq�ۍ����F{}I�K�'�o�={*�9w����'�_>��d��Q���h;�w��ݹ{�[�w����w�G}�ߏ�E,����qe��T6]!`/�W�sqOx���Sc;8��\Z��:wj����ӗg��]3{�o�������:��;�h�b�㞾]�=�M���}�oy*�pz��3^z$G�]R;�y��+|�������5�jG����{=��gI�{�����xF]= ���_����N�E��'�^��L�s�����_����:֡��F���'7��L���@�"S�H^׊�����-.c��0^)��� � ��^�lI��sE`<��q��|�k�]�mJՙF�( x�ht�S!P��<���Y�Xf�Hԝ��cz�ɷ�҅�sd�˕�+b��&��ڗs��湧�o ��^9t����yx��<������1}/I��F%/W��jb؟�
"�a�T�9)IcyĽ4�F1�^�����x�BPW����g^3������������v����rH�^��#`>%%$W�t���L'<����s����}xϬ�~�____w�|w�Hד���^B#;�$�11"�8:��HW�
�	��: J������?_Y��Y��~�������qǿz��R����Lbo2�$���B1���C�˒r>>�>���}g���������o7�.��� IPG#0���K��q
H�c��8������>����}}}|||~9�;��F�����HT^H�O�Ȝ�����i�a���*`%��Gs��;�口�Ώ��~:���k5��f�y2���CR:�ThC�@�s��P�%8��$S��$�Yt�IBV?-��,�G�Ax' "����>$$�c� U�(Q���<���{��b{��IX�� ?���2��%�|�8Y�%��W�Hg1�c5B�%$a*��[[)'D�&$��'"�>~����=���]�Ef�P\P	~]���e�R	}�� k�C	,�0��K]��V�"��Fn�5IC:2�7J��9z=[v�����Ӑ�t;�+��7��s�<a
7c�n_=P맙��Q����ye�lٍuI��,Ýb� #ͱ����a}=l�K��"�%B�L�2�f��B�=1����|����WUe�5B�\��c��$����,�[v��Y،��vuk���[]���휝��|�rC[g���voo��ыqF�Vu�S=��)�-��8�,��{lք2l9
tFU 0�����v�J�x�ؗ�Mq�r�H/�7��-��Te!���Z���c�{	�p(�q��v�7��1\����:c�/=:��^2�oP�����ݹ3�8�v��6�)_^�㴣��-*h.�nn��j�m7]�ܫAvXnlPe�0���'�ڬ���5��%X;<<Fp4�����O�����]ՊE�صY�U�UL�ݨ�ns<��:wu�b�^wa��e�6�U��ke��X�A!���cmB��!�ݴ&���ܜ�˹8����Vպ���ֳW�]�Iv4q����H�^�k&E;3�e�+���Թ(��D�,lŔ&їJݥ:�2�Ƒuv��:yz�?8>i��v�)�M�ݚ��2]n��6��z՗��*
M��hf]�ͪ{I\�'=[A����F%��Vf�#��g�1��̩
\d]��-�&��$�z�N�
�ێ7HX�N{m�Ͷ��]&aT�������@Ү��.��\��[��[1�02�Q�x��70�L\�-z���me]6[���<�Y�OV���K+F�2Lî�/n�
�k���"mc�h�@%�c�;T�~_8�Y_�Y�AN����)nsQ����=Z�L<�vwο���FE�U�!�Hd>������:�w�L�g�5_k4��n�1J���nҘ��8�����U�i�ՙ�b3�`��7sW�ܓ��Y1l�x��F�����pi�	nIv�u�֏M��c0�\%ta�9�F����+��l�hMu���z���u�}��U�a�rٷ0�s�df���W]�f��v���x�bm."�X�\dЮ�э9��w�ts���!���-�\��j+r�!��J)�'/����1	 ���>�e1c׶$�H�~"pv�ɾ��Clg�� �H�e{R쮳ىd9�����',֮�lw%��0�x|���{Ʋ�%�j���������w��-�g;��+r�c'8I��4���>�a�m9��N�#
�m>߂!�1�N���+Y��������Yťϵ-�E5:��o�%��<ԙd�yYL�m��^O`�����i�SW^�� �0�7�qu=Kgb��}���+��N9���N^"��4A-Ӱ��e��vj��=W�z�Vz����6��k��#�v�Ye�YveI{ �J�-r�!�E����KB��� �̚�&m����c*bX�vD���VB�ٕ��Tjh�1��LW��x����s[���|������]\=���kVaÑ����\�����~������=�
"�;����T��۴!B��=>��p:��l���b��Y� ��@���N��;���ʚw��3�{������~G^���^;�FxI���Բ@p��Sf�x�N����x���uT��)�4�9�IY�'+�0�I�<8O"�^c��w��/g�B��� 7w�$���}D��l접]�%��a��q\�qU��"Ar�\D��<Bq��́v�3�#�w2I.��[{*J��|�謂�_�zl96�WT���)�v.�Q�=ڑwn��u�����7�<=Q[SX���Z�����'��d�v{2\zb+/C�HT+f��A'3�$�]�s�DCǨɨ��g���캟xg�X���� יÐOT�UM��f9���4{rYQ1��*�z���W]2$P$�L}�)�����N��o�7/U�r�ȩSr���d�;���iy	��t];�eͿ�Ǽy���f���{wKJ��j�~ݏ9Qם�o��g!'�D�G�82/��l�J@�6pG}�L�-b��L�in�^�� :x�.f}���nטvND���w(r�o���]�������G���BO��yխ�rv$ݯ�q+�����"�.@�� �~q ��ʣW\�O�>��,_����ͦ�pYf���u���.*ڣ�p\�PUV�+#���������lV�&w���A;sq!2D�ށ�әO���p�k�A�w �tȞ����C�^EC�>d�ޞP\>I�򅵐����$Q� s��oLK���={19�P�A�l���~
"
J*��,I#�����������t�L|��,���a�I �ߚܗ���@]��rvpJ�݌́���Q>�R�$��ց���U�#`��������c��{�dL�F��}����Cݜ���9����=&���ך����*�_�AT%���\j��/�F�������:�:������~gy�?|���� :z�~k�1�C�����<����o��)g6�4��WwL��;}������8P$�|�֞�5�*Y��{K^��h̬��H\�,2W$��^w�
ԪX�����u�wL�wlH~gv� �gL���>�y0M���c��3�P~  ~��c �i����!DBM�mN�3(�@��-yO�@�X{� �΋c�t��ո�ל۰�"@,�pzÒ�ÒT�x�x��R����$�ڼ�Nl�� ���r��
�҄���=�LR��D�(���Mj�2!%>�_|�L�1w>D��Ds����9�cWt44I ���[����k* a�1���)�G]�4�7ьdd˙��<�D.���#��Jb;��mS�H^�zd2l�Y�����v�X3��\)�^2�}�r�.�w��΋4���dK3	*�! �����	�00���$I�bf,H1%�o��?�ʘݭ;6��#��>��[,y��K�� iaa�]�m�t#�	ss�ݛZx7e��ͥ[�ܺ�l;
r=�[#ػxN:8���^�<d��v��6v������ջ,���f�Q�91�e�v�I��]�8�g��5�;������<�l�ƠW]�`��<��:�`�Ƿ��?5��ׇh#��v-����+t��
�D������̑܍�/��ÿGi*�9�����y���۲�h��~��Q��e�o@�d��������y�_� eh��y�?C�X��ɐK{z )�y������=O�����.]�P��� ��E���t���Ou��K��ك.�x"Ò�ÒW��;ǽ}׾��Su���
�%�gD1$�t���xð�`(e�܉�=ADA)B�nO�7�ݒ��蔡�H�"�>����M�$�{d��&(�T�\�wLG�>�����i���e���#]f��M6�����;5ùy�Ũ�G
����D�o�>�ev'"o�2��j�K� �{��1��l��v���ԡ�,΁�Q$�����Q�@t���X*k"pT#�����ꨟDWY�c��~������~ͨ�w���.:Ɯ�=0(V����X;��]s�g����<�����gG�������0��eC�!��ߵ�u�;�C;���-	`�JJ�IUUX�i��"`����b�P�n��dA'�v-�C��mO�f� ��r�@�~0׏�è�@Â�C��r���Q�`@�C��zZ�� �q��F!)y�m{�䞻�>n���N����(6҇��$x��(�n��,;�c ���mA\�Wd�����;�'!ʑɄU��[���ea3ѷe8îYZ������o�Wz���QÏ<Dr�E�Y ���@��(_����7����@bqv($Sve7�:.�בe�ф�'��Z/à��0��-!B^�gƆ�t�;RE@����[�����=��!:����`����ȲG�6 �K�끘N�����]C]۵�{���O���X���vO������.�l������K�+f��ge�C�s|ў�`k�p�����?0��X�-�����NJpd`8�'A�+J�}��G����wA�K?w}R��8�vf�`�B�x��0�X5�2p���H����A-�2a����KVY��O�ݏ:�1�U�m����qT�=2%��=v����K�6��$�pH��P]���P �I���_H��Tn�$�Lܲ���Gk��3�Hr��R��c�������I��m�b����O�e�v0�n\fa�>�ؒI��'%s�;��u�n%L�<�Gtt�m�7<@!����x��V���Z�y���i�SX�Ͻ|y��o��%����� s�C�����)�Z��V�r�	��jx�r]çj��2<���F����W453�}� ��������dcD��y��$_U��u]�:y{��VَB�VP"Z��,O�����U��l���=�gV��������4=ԣ�M+7Q�'�4l9w�"�}��WCW�V����vv��w����)�٣��f}��x!p	Y��C<���~�`b dC3BL�~��?7G�����������$�$��ygk���ok �K�4����s�g�i��	|���?����#��tծ-c�D�&p�{g��'u�T[ǯv��'Q�/�D(�@É�[S$�]�;*g�.�L1��{��.�"A'�7�gD��	 �v��(����}d�3G�a_\���wL2D�����y@����n�l#{X��§�����i|�\� �ߝ&<O[�D�8�tܒG^=52�d���8;�<G�!ܗw*G��fg�V��ݷ���	 �k��{c�������O{-��Ӷ]Dx��.�r��9�=�U��.Fܗ,@�D7����jD$׶7�^O�}��~XEH���?��avo��0{A�=�I&]��~^[#w��
REzo���i|zn@�_��,��4l5�p�ٛSH��M� �ZQ�@�#	n����G���!�2?�B��f/2�7IXdQP���E�pVݯm=�<.[)�t�.<P�x:�UV���V6�Ffҥۖ<�k��AC����/�Ky�^��;q��s�`�:8�t�շjqUԲ�^+2Z7mp�U�k�vCgx�<Ez�ڕ�n��RnГ
i���c,�uYޱݺp�띧���y4���e���v������41aMon�k'Y�F9�t2
��]��D
kTМ�����+B�OH�Q�?.��Ok��z��~��9��Ǚ.��&�m���e��1�8L���1�]���xY�+k �{a��?B,I#{zd�k;�U\{e5߹�Y��^�Ȼ���d�u�c k"���=B�|2d��1�D���j�J�\�%�,.�>�]��xo�ǿW_s�'�	`I-^���"w�FoD�1�7��O��/�k�r[ G�\�'��}@�O��EnV_����z����E1�	$>��
$�c��s'e�)m!(�z�^n�:��_<�nn�*�m�x,������8�E';�Yd_y��H�$�9����eG|��&�S��\r�B�]İ�2d��qmH���W��0�)Hv�c=��F��;����u�f<�&z������Jm�-_��z�ܼ�j!�؟f���6�o蘼����cā{?�T�+�>ߣ+,2p���������`�@����~�<�n�x�_��a���#��A� ��]|sL<<C�$]�D̒ ��
iD�w��/�M�{y�+��"� Go;@.��4^����O��M>�iyWr��q���@� ��<�ʎ�8�J'l�P����On���|��%�v�GN�K�L��}�:��p�<�qdkݒ$�v�y���6����Wg�/{ �M��Yj�-=޼��y�����]U�Λ��WAͱ����?��K�yz�e�V�SM52a��<�ʛ�h���ї�ud�$�r���x`�1�����s��f�1u?�<.�2$�vA�bI����ѽ77l|Ő��9�[���z\�,��Rs#>��Oa��f`�0���˔��~w��R��U/M#���Μ�O{=�Y���/�x�����E��#����|L��~��n v?o�;����7Fq+G�� �y�ݾ��Ҡ�߻7�2��n�b���پ�-����y���命"��'�LK�mܹE�c��.�,8}�a?Ip&��nj��bOr��HP�\w�{0D�i����x�ck;��ݶ?>��s۝o���M��D���B�}0�ǻ$��� w��| ]���'\��.�gr�_�w�:}.��&}�_kΧ�6��7<H#�G)��#C�Ȏy�"�\��.�K$��Ǽ}���E%������n _I�o��66z�M���l�#Oj	{=����������r�#�~r�,�/E�ygz�w�.h7t�!y��g���̽x*�����(Lg��;c��J�|������F���q���pap�n�F����=R,[���k�Q��a5>գ�Sώ�%�}W*�����S�4h��^ʞ�����B��+�lfq��2���?M�K����`�xԆ	��p �W� j��t������`<���mC�F���{�����0Q��u����uԋ��z�_Oa8�� _L[��X�@�i� ���}��۠^�䱠�`�/���� 0jS�w`���i"����P��l��gW��H�7�@�����]|� f2���#u�������G-V`LT�&�%;��9���E*3���T̤�)���o��2~
�8IrD�H�!�z��~y�2�RX�����@%�N���w��g�����?��~?____;�����<.&��ɗ���ez#±�0��4��u��]r�]�.c�����>���������k9���r�-
�=�0�Zb�$	<R�RqX�'+8$�J�X��+���A������}g�����������q��>^wم�s�rﳇ&5W�����*Õ�x��sι]�s�9�������Y��~�������w�|�o0i/@@�Yy$F(�GĭF��@R^c����B�kj��XE�ޏ��ϯ��~?____�=��]s��D�AH@��b�D���II D�����Ĕ`<'
�-S��ˮ�G����g��u��}}}||||����ƅ�C�����UB @��C����b9NF��V0���*V�F�\@ O�����R��q8��Y�a�D�$^"p��TC�� ,�T��Y^���1y�l+�l����	���0�c��D�T�!ؗ�"��tF����	 *$8I9�3����HY��X,Lx0��)�����ڏ���#�8{����6��xx�H�K�V_5b1��h��cݯ-�� ��<��������Ǜ����Lv@֝�A���zO�h�e��j.$�U����|��@�eܴ� ����>�;R��'pT`�Kkg�h5ͅ2aX���Y+b��^��ɬ.�;����gC���9��� Ad�j��D�{}�;iuB>�܆7�L^�v��"�D:t�>����d����I�o����h�	';`y�H�� ������q��������DBt���c; �={�D�d��<%�hCu� ݽb{޸u<9������iQ�!v�q��Y'otē!J��)�.��b�0�h7���v��x��;��7n�����f�:s�qw�*���,�n�u>15�1��+B(xߎ�����N���COB�R!�ƿ7��Ť���s�祶YB�f��^T�$����H��"�?�Ēv�tI�K܋��Q���@�"⡎�����ٕ��jw4[�nS��t1Cv�¶��{����!���z�Wʧ,�M-g�"]J� y�V��Q;���;}9�\ؓ�~ِH�������_�
�=5	���ӎ����:��`D_�fA$w�[<��$])�9S�SDAwN�ϴ�$��覔	=��w��R=s��e���R %����T��WX�p]�D;����=M�?ne�O��-�9"�;��%��� ���t�;���]~�7Wװ�\�A���y�OD;�<s�������&���$�$A縈jd��v/���07�n�|�`]	jA����޽�N�^V�5{�R�q:� �(���S�N5�jC����}��:���F���G���	c|�9�4��w�GW?r��<^8�\a���ࡑa��A�6��ȹ^6W)����-t,I�"���܌�L�;f-�t���EJ��E�yNu��S1��^�\��{DqhH9^��u�C�5v�����,�n^�r�����PM����:Dъ�[�4�o`vz���f�9q��l�RW.ъ%.�����5��4�B2ض�t���N�/�<K��L!]k]��>�ut�����R8�'ln�Kkv.vؐ"9F�����6�5�������BŠ>��TȆH�{�H��HM S��Lϖ�o�<�<%�7�3����A��"�=���9w� �X��ƖH�P���5w�bI�^@�{z5��~�NW;������L� �軄��xF<��1������^��彀wm�1gtSbo	���kDAwN�Q�$����I��Dy���c>K��>w��AeZ�@�xv�Xz	�DC��1�� �ۻr|�D����g�I,H��ē5��kA����u�*v�5jq�K-�s�V�sm\���Jܕ4�ſ���Q9i�̙�x���I�ށ=� K�fL�@0JL����>��k�A��aďt���"���l�s��<D�D֘�Pb��B�����z�}�z���ڻK�bqX��\��[��z����W�=4� ���y��qpz���W!�+(�!�g���>�;��!�� �}^�$E��s�`����� �u��ǯ�������M8�"�:k/�A�xވ����${����G͝]U�����~��xF=,|z'�B�����<jd�,��>g�S��r�����M�9��g�E���{�������۳�E�BJ	���2,I���Ň~Q�#2�N���搉�[� ���`D�;��ሪ����nr�؋k͎γ���Q����z��/���`*��W�?'*��4����7ת�#k.%�ie���	c��fX��V!���ݪ���ݘ��C�AE)ِO�����ޓ��L\��ِ�1 �[�uḍ١&��j�v~���rx�x�aǫ�-��~��1G�"��q������}32�Ǟ��f~���*���ܨ���KP�wA�n��l�x���ҋq�:�	��I�"��5�����pT���`��i����
�.Q���d�������~_�\�4S.w��D�
w��(�N:���󐣼��H�݆�ׯ�ǛWBd�綝��2K����C���=� ����	2@�ys����3��O�ɕ���1D�?(�P�����c7�c���Tk��Mt�h�-<i�=A�r��v�םv�rJIm��y�z׹QU4��O��#�� ;1o(>��c�ղ�R Kj��~׽j��<�t�ư��D5hJ�u;�T�j-�Ｚ@#>�m�PDq�-+��A8�3y�ܗ��cA5i��EeU���xkϭ#Z;Ǥ.N����l���X��J�v��Z���5tݮO�8��U�2������v���^�M���"-�;�ϋ޻W	K�4�SD�B��P�/i�0����!�F�C��7���dUd�V�W%��Ǡ�\���т�Hf�n<�m��ہxhP���t�C�I�>�U��OV/^��|�$��P9��̸�����G��x�*�	�UOA��F��e�=�ԕM:�0=�7�����>�Uf�7�$��c�T�$x�@pX�w@Ǧ�q�o9��غ���UڲE6Ǳ4	���Jc�i
a���R~TY	n���s߻��_���(�xt�$�Vh�C8'r�E2gcէ$���P`ވ�c$��P	 ����k/c_{L/K�/}<k�t��"9Yh$Zj�D�{�)W�Q��_��@w�>̴WDDD*���ْ@֖��H�׷zӓޠ��g���N�t8�zs�z�{}]h>�UW1�ss<��*��9����7:"��C��tg���^a9�=��ĺz{�N�2`An5�Z&�xbP������Ff9V{��c��g�%��Ω"��BZ�4�lpJkR�
���h��#+�W[E��C����#f����Q�b��EՖs��bH���s���k)��e�^����b�C6�<E&�ݺS�MOX|�nxڃ���l.ݪx�b�;:�+L-z�']K.��\�f��n]Ε�:YC7ic�X5�'��S����+tѭ��u��13\&�]yݮ�s�ca��jN������	�Ih���z���.���A�+��I�sx�@�@l>tA��7�S�+d���L�.�A��:DBxJ<ʝ�gVo�w��MN7;��ʙ��H�Q]��W3]|q��}7KĈ�����߯5�<3�a�>��>�r/٧Y��Z I˾����"��>s:y�ϋ۱c�ɵ�C��8`.ۗsD�	*��� �ށW[c<�A<�[ȰQ�u@�
���D$R�@�X9R�`���e�D��9��S.��gDv�@�4���=2XS$�"!�';�@�����^��9m"�Z��eEu�QD���u�]���$={��N:�G��}���j,_wS�|�k�s��@>��^雞�Đ��L���y��u"�g��%��y�J�ۼ��0t���w�)�Lva栜3�%�''p��9�5r뗊�2-_���]����O�ٚ$G�
���?H���>]�~���J:r��x0C�5�L�1�79�5_�D���p�~�qfL�m�,/T�ލa���Q	�'���ف��v�G���~��Ou�<	��搎7��ua"	�$4�`v�ۣ^��RF��|m�<#��$wti$Su�����Lp�\4]�5���u�G�����v��)��u7v$�t�)۽2�n�z�/����R�"�W]��(�Y-���E���H�e�6p�.�lpW(�}��T�����|vjA'/� �$J��+��[�<$X�'Hy�qZ��p1���� q]/�,Z}�<b�^�%I�)����iD������~�	��]����L'R.����$c��ؠ}�{u�\񿦾����t��(��y�b�^y�ݥ�G&��Ӿ���-x��p���]��w�/�6)˧�T؏ˈ_��Ɛ�!�\p87�^�^x�yQ���Ӳ/�����=����TC�s	�@�ќ�oM�oM�`"qiA&CﺢI �����sy�����ة]L�A�}�TIvL�&N��K�xq�����	H=��%�� ��g�\�}�O���I��֚V�h�j���W���ƙ<�K��Ubu�T�4!5�W�>�M��T2nTpr�\��#Rd�w�!2��AE	]��y�mS�9x��ULz��]l��]��� �]� �(�t�b2��O'�>(���%��~ғ�H��u�'͌Y��ᥒ�ў>`��r�e��,���A2@�N��W�3B��`�	Ԋ$��0���P��.�8�6�^��lH{� �A�ܲ�����߽\����i���,)Zr}�܇ީ�O���Ơoׂ*-h��1P����K�w8n�d�͗E��m�/�_J�`�*/��`����ƳM���Y'����w�h;����\+��8I`LE�du��q�c�G|���]�2I ��E�D�]�YyT?B��!���A�~��ŕc�:�\�+\����n�ֳ�j��5� �㜈�
%���R&�y�,׀�sƹI�|�u�ӣ���u\ɆK̯c�H#7�IA��xSB���,�vaC���Y�U���D�f���A>[�;ysv{����e����>��O��x��R(:ۏ1G��Km�Aw��7WO�~��$�ݱ � .��q�)?9��bP7L�p��i�[df�͘�
dm^�gH[�+��w�>,�GE9�1��}�}�N�Qɥ��/�!�w"A�Q�e��@ ����C@�ܥ��goE�L������6��	�:�����龣Ьyn���ޢ��.=���k�lO ��{	�'�=-Ъ[�ooD�ś�r��
��bx����[��c(�yҾ��=�I����t>�^��<�5X�w�܍��<�݂I�|w4gN�=�E=���F%����nⲠ�Îf���m�Ѵ,�g�o �kg�+�����@f{��Ǩ�vSӵ�U�Z:�v/���%}
��O���%�$x���m�y��Q�_T�j��6�}��wY��
�)�U����р��Ĝ-��}e-x�^p���]7�ؙ�����e]ߜ�����95���|v�#iz8y�z��g���x���x�����[L��icn���^�!�9�^���s�ܞ#��ĵ,*=E܋�zo���ۈ� �
!�E:c�&�X�ky�η��ݫ����h�:�6��.�	�bY�D�����"��J��x�y�Z�����T�s٭va����/��!�ٯ;��P�!8<s��&ո���y�5��D�������ڳw�l��<�����J���X��5��B`���F��5�F�U��$����	�p�wK]��<��Ɉ}�ׄߚ�Xǅ=��(�ݞ�7����!�"ϩ��w*'���l>yⰻ�3̼�o�p�.I�u��>+�ڀ�<=���n�{�|�)]��n)@��7�GK<bI��8�dK=��_zO?L9�0Γ�~<ʡ�H"��`�C��=�#���ᒜ���^Ia��	`b"��T�ĠOuIvY�iu��߾���Q����Hdz���S� ���$ �e䶹@Ŧ�SVD�|���AIbBz�T���D's����ey:��� $�!��# q�*j6 @� �
�y���u���3���}}}||||~8��LW�HE��'��?;}������҅ D �9��rC����=���������g_Y��~����>�w��I�OG�p$���		�z�-�,�`,|�s�냏�Ϯ���____��<��`��1)(1��f~� VYX���X�(��J˹3ч?;����;�z�������������<191rZ�|-�_�X(�,�@������s˅�9�������8�~���۷n����#������ ��5�	 ;��)�e<^�
������G��g���������n��Opx|P�N��x �R4�T�0��htX�F p �� ��)V �K# �I�׬��v�BZ�������A�Fږ~N����"+� �!�B�Vz C�/�t����G��\X���c7��c��W�"���X�X-�B��ó5l��K��/��x�ur�Lv��n�w]��Yf�9��r�N�����^}[����M�֊��:�W)�&�Vs���lu�7\$g���Uy��0�#Y��ػ�8�C�)2��o<Nx;J��3��(e8�:ўf�z&}��l����8��k��{7b��m]��F�L<��"�㎋WM̷�f��8�N1;P�Z���%��M�}	F�b��!4Yn����v�A{d��=8q�-'^��b�B��[�ٞ�2��Q�������]�q�����qsOQ2A֎���V����Q�X�k>S����j��gv�2�i��lU�ƶ� ��m�#���Jی"v^�n�Lr�Z����]�g;;Z�h��Y�k�3��zw]d��&խ=s�,Ofzv#�K4^�%�TqZ�s^ ���Wv`�Jj��m�gt��A�۞�i�z�qo=���	x��M��X��VD�i��KSi@Y`5j��n��h��;��7m���ǃn+�=.˭���@�6u.N�fv�;���3�;�۴�ys�x�z�q&і��6[��Mm̙�m��W��N��^{x[�+nMn/#;��N�����{9Y@����	y�a�d�y��E��vqp��u]�Dc���H�,-��n��B���������^)�l�==]hw[�Y��R:�|o^�ͺ	��W����z]�k��(:)D�YV�E].KJ���6H��ƒK���s>���nc�^���o=�)��n�n�J4���k�� ��M:+r�$xs;��.j�ڲU�~>#s���h��N�Y��!��Ya{F:����[a�s4E�r����#
`e��#u"^�K�l&�X�;̹8/�Ҭ�v�y{���z���шfa�8<a�t���^A���[hƺ��x�jR���!��)l̶�K)Bh���q�Ji`Ö�&�ЁjR]��:y�K�	�a#�wHp���گ��%�㇭v�Z]㸋OdO>	1���v�eZի���l ���^K������l�H�^MGL:���ƕ�͵t/ �2Uag�{^$ؓ����Z��`A�#�r��'{�ɗh5���w�1��mq��[�ݵ<K�P�Q8#�o|�D(Na?���K�HA7��b��r�y�jo<�\�C��+�q#*W�Cm�	�Ӗ�
%H�l�N���5�.ߛz2a$$�(c����=���Wzr�/�1-����A�QwzaN��;sK�{�IY,e9K���Ѡs/�,It[7���o^�9�!"��Y��z=ރ�~���@(Rk%�$��H=��*������NL��dV���NT
�~��޸���x*�<�l�5w�1�8��ȐE6�L�Y����������w�+s݊�DIJ�Ŵ���v�jL��mr�=SK�����^��e��
n����Ls ���	���<�s�����OJ�'��h
'ͽ���D(Na=ЦV��q����ņo{�)��^�Eߪ`,g|F�ՠ�g���j��7ۥ{�Bl�w�b�G������юq�X���m����s[��n�X�B�~XA��X$ ��͌�`B��A ��&)������/��ô��J��V���KO>Ȕ9��� H�c��=�����3��AC!���'Y#}�Et�$P�	w��u�.�}R��X�z��@jG�y!P�%�w�����ίBk��s.fI����@x��R9�̿@-d�MZ�U����;��t�$�\LQ#�O��^n{7���'����4�n����ԂvsWm4�q��Ɨ5ף��8d��^�����F��s32	vJYo���!��`�Fm\�;s�/ڙVL�%42�ʃ�$��Dp�S��6Q�T[S$]���q��u�&6jF��C̺�Ă���S8�7鉾51s]ۄ��o]���'��(tˆ�.�k����T����US&֕�8��M�^C}�}��zy�/�)���d숿w�C�������
|���b
��o�5�wHb��CX��$x�������1�;�e���|�
m>�<�����ڽ�>�E��)���aڸ�$�!��SӴLsw��Us0y���	;��v'��#��0�M��&߃�����2D�}0�uwD��~��}��r	&$�y�;�����؆��
LJǜ"6%f��-�1>��A�/u�h�K8���(���K$Nttɇ�t���}�@���N���O��c�^Ei/	4����>����������h�F���Q$_wJiD��>�<cԏ@�9�^|��W�	�<TB��,}��@�n���ܯU�!|�ɖ+��d����w��w�e`�Βr�v�%�7�	$Wu�c(���}�кj�0�D�'49��1;����p��{��B�'�\�����ӝ�w�*DfK����_8~������!���9�|i���$�M��q�D<#�Mx�Y�g�21G��ў��{hӏB� ���Ă�Dk�_0�Q�H$�3I'�m���a�p7�+a��u�\�YL��5h��"wR2���[[�x;���1˝���q�xZ1=� ����ᾝ�Z`�� "�OO�=�z�,�YD"��>,��OA ���Yu�C��tD�E2G{��v%���Q}�><�k�!��w"�������a�*d���v8�k��6)�h�a��sr$H�%�"
j�B����P�@�a����W�x����w�bH;!^Ǒ��2[ƻ1]RpToSU[}n��!�^� ���C@ �,>����U�@����u�'d�G�#M��d�[\��B��<�ݾyu>��+j2�ˏ^W��&vÌ�t�z#alp��O�}{����oyxg��쇙����6{ڛpT�<�ڳV�#���f�O�w���a���Ć9<�t{�>��{�/�N�3F��-r�rKk\h6&9+�����m�i|��q�(�n�e��F�L�A�A�����م���-ԕ�u���y���e�r�a��@5å�`�ތ��v����-��۠9y��W���1�q��� ��M��n�:���:�����M28�x���C�L�YN�;���c!�v�N�3�8���a�ִ���t�m�f��������>�g�.����yܟ�e�i��WزsŲ��z:D�ǳ�T���b	N�T��t!9�}����E47;�E-؋d����`d�j�!�׽[$������bv���0�]��HG||�L5��=�����H5yb{_�e��$�8�8w����a��̼�͙l���T���`�*�v�L[�����x�O��Q���?yG�vs�� "���k�{��ky?y���[�BY&'���'w�K��ʑ>ʧ�D M�?_}rX݁��g��@Ţdݻ1��Y�di���$���/��}��YK'���%@7�����K1�cձ)�ÖaL9�����C�NK��;�A�KPQ�7]��s�￱#W.���K��K^�ľ�|<���RS{��o��g��^�5ag�k�+��X0=ʖK�pBc�4uب�f!���`��"Ƙ�,�� �2 "3�_��3����� �ݿH�T����GLSU��6���.���l���j�{�H�I�z�V���=톍+L1�['^��F�{W9��(FqO�ֻZ�{�����]*7���$�w�s���Lxu7Hb�O�v<e�+l��r�r�95@��3*��ؒ�3G��� �+�I �ٖ4���m9��w �uQ��/q �%����^��u]�����Y:��2�������\sO5��{�S�u8���ǵҁ���Ў2;��g������>�`:Y���^ݙ f���B�!���D�}�z��1>��[&;�tɆH�ވ�<HZDȩ��pq�<�z��]ܗ�Q�2�b�� A&�p&�ē��S�D�eOz��^x�N�������|UGo�M!5�/��u�۫㒷?'�{yv�r+��ū	_;�f11j��������P�::�������c�ﾔ�$�2A�-�`&9wR3rۢARVlՁD��a�>�yi`�vY��K�ca>z��w��ڇq �]s� ��Ƚ��A$�[����N�6[판:��IwэA	���ڱ�ьCm���,����&�;)�`U���
�ȕL¡8�B�� W}���,��2w7DL�$S��W0�P���{�b��[u)s&�|��<�;�� �ZP=�>���w�c�@7ݾ5b��by�c��,�1k$�m{�s�25`-d4��[��Hw�n�pH��"2�у^@��<�����qۦiX�-ZqѦ�S�DV:M�Q��?��rf�o�Aq'hjq��쇝�O��"�ˢ�!(�-e���I-{@�+hRU�-�u)"J�L2��9\��z�v���ߎ��=�yk�j;��gK7�7��x��B���޶�v��ݮcD�����J �m�D�u�=왋Le����*���w�m�ʁ�+���k�L�)b��-�v@E��vH�ށ�F��������l�HDn��?��o���"��fh\�y��|P��.�]�x�o��<=�;�ߝr��@d��_#����|��ד�NO��H<��BRĝ$��Rt��'!�u�[o���x<!��y��ӓg������ ��K���t���T!i/_W5wzSEx&]N�D��^�D�=�^ٹp9����������4q���p��9��v�]λ�w�`<�tAJ�y��P^	tf��9��
Ք�;��D2�Dz6�Rx�z� �15mcA��'�Ǡ^b��w�rڜf{ÞfD�>�|Xভ=�$쐾}#ZB]��1����M��x�֚�Do����Ru�[xc���н}�[*=^�w�{��}�����!;C'�ޙ&[������!��;+/��bK��� �,��g��"	�u��vH��$V���/d�;��^�j�Z�'} �mgH�M��=룱!�#���\�-���f�ƤX�v'x��f�tH뫘��d�2k�K-��fl'�ix�����S������V�`9����o�����AMP��*cа~��2�8�%�!��X�w-r��k��ĸ�r������l��γ^Dֆ�An,�I����V��їV�����]r��LDku��W��U-�^�h��n���m�w)�E/*.���=q#�/�^�˺N�o�g�p�^ŧ')];��xݲ�m��^^�B��y�vR3��1�����Ƽ��B6��{\�{K�*�pl�tn�!���=����e	�YVe\��+Z��9��;��!؋y1��@��o����/ w��,��j�Ȇ%�{�L�g5Ѣ9���	���dj�f�|0���FG���'w�ܿ<��t��LP�g|���H$��{�[�^=.�`�5���r؜g����O4�Gّ-(�oR���Kǅ�n��#_���?ow�]���]��O�_��טX����G��rw:�dK%)
��v:}$z�Y�4�� ��u�h�#D'�s��2�}b��w�F��˹�C��v�F׿}U:����������m�X����n#b�ȏV��Z�.��F�S15��`�'���u!9H�r��i��ngv91��6���u��}9�}�S �J�+�z�kK�I ����2 �g�O��{�`i�配�n��#���`�=@�����xLi�lX�r�����J�۷La�p�:���L��tʌ\��޾Y�BK?$K�_/p<˒�~��{\�Ig�3��CǄ=��I"�����b��L	�sD@�I��=��c>���H�4���F+d�p5������\��)�'G�tuO�[�����F4�2D۾ �{�<}�o���Ǎ���[2�k΢1JW��=W�����o�����LA&�Y�A#��]2V?�N`Ì~�}ܥb5p6{k���Y܎��+���ykb�m��["�ج��4���q�Z*��E1�K�,oˡ�$v�D�'��C���Ո�q,H�{0)����sµZ���H�P%��Et��=A��j69I�l��p�	�=`u�IL���^�O�J2zJis�o�Y>& 't^G�,h��D�$�A�+�������n:���	��z�
�F&N��BH�q���]zG!����{���}�������
��n�wzgb5Q<��yT��x����I�^�����^ҽz�3��1I8?%��d|���d�=��-��LX��4�y&�1s�4�9>����	p\M���!>����.��v����y�شa��l�׷ӽ���O��x{�2��cfI��fˉ{�ն���.t{�	��[܌�}u�{:��|f�u?wbl�C�X�_Y��/zv�{�!��z��spǔHn2DX��o}���	�	�ٯ��Rx�w�|�9;� ){ ����V��#Cp���_��+�_{��M�{ݷF�g�7|ݾγ_i����y�"���߮]�\�9��㟷���w�K.�^Еw��x��ڐ��e5��eҠ;\���4^��ot�q���������>㥯�|����V/o�~�%o}������k��vu}��	�b�o��=s�z��L̺ǋ���Oe�{����nq���ɽ��}�w���r�3�O�>�y��?i�}���s>�B�{݉"�s�����]&[x�	�{��W�~���ɾJ��j�g�ߖ��&���oD�b��-��Ӧ����\�*KB���h	M!p��Dx�E&YY�ܠ.<DE�O.b��C��m��R�TE�#�0DjMVT�-LKd'�p�ҩ5�ǌ��[�ci�0B6�lZ��(f�$F��b�^��~��A�8%���J��M��P���\�ᗝ�ə�J+�2�	�9���5S3�O�w�����BLB@�
(��q�@	 �!9<��?]f~:8�~�����������*��;�3�a)9$�N��
�b�l E`R�	�q"F����}}f{}��믯oooom���:*��P	�|�#� �u��p@$0�R�BC�}}_Y����믯ooooo}ԅ	����沊�!F^�I��1:
��3��e�0�+��~?]}{{{{{z�����AL|���$x1VBNH�Y@ڝLA1�\z�:�>>����=��?��ｻv�ۿ���@'�APD� �q���\��;/��ys�˜���~���O������ۻv��@����  �b�B��X@`�V
���Rt��˫8�@�!�ІC��pB HTc"DD���XAG�@T���u*��bBtX��I� BU^���8�Z�Q��#��'q�VR���'�� �`���%�'�S�tae%�C3@�RY�k��T���w���(wG� �1��u�D:1 �.���	��/�V��KoOD�$����$�~�ۚ�{1>��]���-Q �mm�p�øN�����2y� ���W�c�{?�{�!����>b�9��>�&����m�8��D��WJ9��"H���q������c:�i�����5\JG���'��V���Ǘ�$9�$�K��&����2i����l���%۫�}���П=�m��|cW�>Q��/�	5��%Õ��c� 'y��:ȗ�e����F�\��j��"��#bg6���c�����-���3fL�gLO�'�P2ɐ�Y�x#t�A���)��<��>Ϡy���vJ��?nCD�wH��/���^+8����o��9�'w���l9J�=��c��r��<Ɔ���0�N���тYާ�^�ԙ�HD�+�?�b!�o��9�x2'$8{�>���soL@&�6��i�d������Eϫ�&��"�=s3$�M�&)��u���-g�U�AB]ptke۔�k�D�Q�;U����W�U�G�e�3�;��I�����e��&�qϒސ ��{"������^7���A �J� A��5�.�P8:���j��D���骉%���Ϯ^�Qp�k��*����\4��@�m�gZu�4C�g�^��D���T�g��<�3���]+��kGP�X�(.Ru"��ж��y����s"	'�\��I�%{�⬓��j��(9NZ�����Cb2_�rx�fi��e�8�vR�3�LX�wD�c��KZ.k���(�>0�S�h4��s@��[�!��l��q)t�x�-�䆐ya���	����moQ�W���·�w�8�*L2���0q�!�%Ͻeܺ�fF ;[K��u��Ǽ��<Me��Y��R���n,��'�i,�;(���v�]{(=�'bSF�[�+�6�n�v��ִ<��.9:�g�(:NS�#n�ջ�&��^�5��<�Ue�lu�:��qs.s���Bj�	Xt��U�Fh��ٰ��]�_���k��K�m�_k�OQ[����B5��e��0T�Up$�5Ѧy��Q�M�ߧ�++��iz��QZ�� 3;�X�ǖ4���1=φ	v����'�t\/g<@,�n�vM\�@�I#��0I=��$������2�'���8��;�N��V�����LH�&U��I�S
��c��fA#���'3z$���wP�CD=y��L�/:�J�����5
aOW�)��7�=ӕ�'K�t�Ѧ@'rr�9B$�G��3 s�$��MuO�뺦���L ��@;��Xc#�2	ws��s1K��#�$7������μ�ٛ�0+]Sڷ���G^?�����q_{��� :.���7��R�s ��#���}��Z}���Pb���q�� �Ιc�H;w���%�	ׁ2��{*��v�N�az�6�9�y��FT����
B�� ��t���[�+�ގ!�څxw�h!���C׋�����#s���؏��,�)"K b��z��mL�7��IbA߯�D��ӵC]yA��@��:��ú.��o�Q�	 ��p#�B���蛷�0{����ɽ�ͻ��w�D�k��FAP�@�(A���>v$���.�FC��IIkal}�~c$�vD�}(u1*�y�fj��w��ײK��oh��R*	݊��̬��zs���=d�&�[�&��$���V�o[>�[:N[���"=s�=��\�Z��M1�lT�������x��Ӣ�мN1�S���2H�I���A�!�~0����ݦxyY��n^̱ �%�]��5�d�Q ��^G�_WB%U���w���-��2@k$-\;��$Ok�H�WF��/Jc�;+C;��ץ��0*������_3�/p��9�d�^�!��eK_��y���7T�� lM���S��|Y�y�S�S5�
�A�b���������N=�G�3 �x;�7�ﲥs����c���@�t��hk��n{�4"}���#��S.��,	�wO��s�����~仠�wϾ��'U��K��a��y�i�o�,�sݩ� H��"S;�E,��*}�aY�˺g��iqw�0��`�`���bζ�79�8��­�>}~O��D(r"�q�㾀�E�.�ӤV{�$��%� @$�,��5��|3���a�}���������'2ڵ&Ȼ^��%圄z��;J����YՄ��S��Ex��,���\H%63���F,��;�xj�� ���BA#�:dq�������c���=PG&0��L�̖2dv�fI"����ǈ������l�?�Y�^I^�5��P/,pO���w��eef�]�{�	��t�ѧ7�F<���E�,�{.�y�&-%`��}�&m��,�p�,&�w�Z��S9a�҂\�}k��X�;26{˞߆9#��0�5�tH$�w�#<׽�y�޻"p#��Ser��(��Z����uk�vkn��q��;�K�A��������J9N�:�s�bk�$s ����/��j�r�����{�(['i�B�"!�<���b��6�)���2N�s$�������{jr�v�$Cd��r��N���mt��L���=f�w�4@>K�V̒e�����)��p�|�L;'�+��w��������=id���d����ˍ�$=^�1�;)$V��C�:r��`~�h#&*��}�r*(_��o6��۽�-4y�,U�0@��H3�r��P���;U��V�t�]ڈĻǛ���^~���
��<K�}pw�u攠�a}xˌ����1�1��CG�i��8���OI��F��sZqZ��d�,�Øqӣ��ϑn#e�M��f���I�yn��J�)&/$�"��ƙf#F���V\A�X��	��43��^��s���v#î^˞�W�ԳB�f���U�\��Q:Ex�����-^���\�� ��ۚx���/b�\V��0�[aW���g�(�^f�`�n[EN[��VlF��s�!����2���=�P@�L��N�x�A�yG;��3l t:PK�#{cjdK.bYŻ㸃�� ��1T��B#�d���%45�Y�B�S��`_27OR�	��v���{֢�,I� v�4��UY���F���1
���`��2��}���,�����j=4�w���]��ݾ�ވo�f�&P�W��c��"�c@�2X�5�A���`@6��˺ ����5��]�����|��7��'���Q^���8D������c�]�;s�'�q- "�^ف ���~֗o��w�;�0�R6;�l����S��4�q�X�S��ȶ{j{��u�$��i��5C�N�'�x�n���	$���2�v�H~��1��b�F1�lg�C��2�;&�A�L��:x�>�Ж��4��J���y�Y^����E�X���?���O�4����m"lt�<<���s�A��`�X?��sY���9��C����D�ЕO��n��ݿ�y����q
N��A �oD�-�m@{�R���-�Rů�D�w��A-@f��#�ȈP#�6���������y����2@�AݓR���O{A����e��Ó�*�~��$WlB�~詎S�͞1V��A6���d�$J�y�"n�>9��&��/*�ƨ�Ȉݳ+�XcT�hc5�[Zd��	��:������s	��_"^<;���1�$��c`gB��6������xv��7l"�t[�v�wh�N��w>{bْ$�k�#������7th�vͭ����A.�ް;Zִ�[HO���6�nߓ��;A:eF~���t�ѧ8�P�dxY�u���<�3�,cx�6D/v��Ї�j�=��x�)�E^Q�[Y�k:`
`&M��9��dI ���!sv��!�è�zϪ)�lUm5LR��8��}h��I�dA��Y��>�P�黗35ªʈP�D?��x�I��<��v�x��Z�^H�ف �6�OG\Leyy6�H��d�T�p�tZ��+vR��3�e�Fu�f�5�4L�Q�Ϣ�Qu�&!�]����7Κ!�;�3z�>���-}���>$��A���l����͘�^\z@]������[ׯ� ��#�3ޗ$������y0�A5�l��R�Lmy�p0xs��9ߗ��G>�hd���l� ;�� t:P]#Ǟ#}���Eϓ�x�$w��ع�׆vRg�����o N쾼��g���Tg���q/jX{u��y��fѾu:_��A��:���F��໇��Drk���hbV�#���<����إ-$�{���g�"���H����+����Ui6�%�"%�����h�g�����}~W���]��lv>5eL��V	��n2�B���¹ىP��cVأ����}什R�`��qz�J�i���C��g��$B]���}磾RTB��n�B����ñٓz�Z.H��3�$�ݣ�0����@�Ȳ@�&��s;�H�_�s^����T	&Eﬃe�r�E�}}#*�ȒA ��_w����|"2M�}2K���(B��ϥ V�/�����88{�G A&�q�H7^ؓ�F���Nm���@�<�c�����
D�v˦�X[$�����R��a�X@�	$]gL�2@�{�"/n/����b pO�n���-�Z9�������0nx����1�.xC�e+�}���[��[�!Kw9xi|�Ź콺���Ţ��;�����W��n�G��@H�޻|��k�i^і<������������*����u�|�w��^^��w=,	�����czU�%���s��go�0�w��^�ͦ9q����ni�W�����$�༽��R���\��;ݧ���������b��Y�N�o=�o��{�g��0������g���̡���"P�W�K��������B��M(���婈��{F
J�IV�����, xn��8�0���/#4N®��ҽ��0F��m��>`q�;�c�q~����G�����~�}�k;٣Vm�9u^�ϥe)������o�������r�=.�F�� ~�r���К���f����xǾ����ơ,�-<;���m~ʼƖ��=<Ş���4b���3���n���<�q�`��}c��V1���<�{cɅ�{u�B�^D��C2=��@��Z+������w���'���ל�����^��w�C��/E���w\Hd����=��<��Ɍ�����q������H�^�i,Y�Y��x�S��n%�/������2/�C���/�����6{���Lg����D��Y���, n7��c��F+c`(�ߋ�[����l�L�=oz�C���4ݾ9����Q�=Bc�l�lcR��a�=���i+=�uO|���8;x\��`n804��ln����Dm��$�w�$iĈp�ڡ�s�[`D�����黸r8�s�����������{���nݻv�4&界V	B D'���19:V�Er�����o�������q�����nݻv��!	����3{���u'�a X��X�� �^��.q���������8�~������۶2�@	��+���	�BF�8�&ճKѹ=~>����O����u����������6Z�L0�x�z��*��ր� E��I������g����~������������r	� 	������#�'%y�$	�IO�	Pg�����fz}~?]}{{{{{z���ȇ+ #�9Y!�E�R
����&�� "$��!�2YK#�Va'=x`R$ G���	�����FtYl��2$`ߪq �Vyzo��ƄAb+�a�d$?�r�8�ebrF�����f��{��@��eoV-��4�����	줡���%8u��~��r�uEmӷX檹ss��R�u�U�g,�i�r�ܓg��f�g�6�#��:�s�r�\��{p���m���K�<�ي�ǃDM��9�;sP���:Z@5�E�6XÜZ����!�׆�^��t��&j1�ҷ!Z���2�):��.aIsv�ף��N.^V9�����[�Z�s��2�kt�&��"�R=DZ:��1�g��ArN$H��ҋ���9���Ɖ�h�&{uOU"�x�v��Ы��h�-�,ayP�C���q��<�v�[�&�=0���DǞ�i�͚q�aphJ0Q�����	b2�GL��wnu��tq/6��21cb�\��Pa=EM:�F]zkbX�
3{K{,뀚���j�"�ˬ�L�o0B��c�`��n'�)�����#d�v���Na �u�D�%���AP��uq��6�מpB`Z�`	k�T�mm��s��˻u=�\��Cd0%���mf����T)��G��`��h��gk��9��D�[h(����3@��0ckLa�����;�7�g���S�'��Ɖ�́��eu�;Nnznz������H3m,�R��]���X���r���	k�M��P�ei�lq�0��}����A<y�uv�tٸ�ʖ�Q5�K��������W[��l���۝Y)e
�f����G�U�{i�c.ok��&{�C/=u�:�VW�W�y�^��R�vQ��� M&[��mx|�hͷf^�W���7C�U�ƺ�Pu^s�uۍ6��WszR�;����'`���'�F��a�na�k�z�"5���Z��t��4ݴp�Ĩ���Y�>��߆����t)�b4W�dsq�
�ub@�������93j�<vC2�kہ�V�s�eKaֽ��(�.��;bkKF���	ѻ��qP��).�<�c#�^p��W��6׌�ν��6i%�u��EɷhxiV���5�LZ;
���y�\ě$�Y<4j�MfC1�y���G=�۞C��uc�qr(jo���}�Q4���]R6E+V][��0UE�VE�"�fݻ=�B.^�;���Ѫ�U;[x�QN���� [G#����I��{�I���20GGw�V�S��4�W��PS�h�:�"!��~��	~˼V�� R����F�]w�$�;�/)�k��l�OE��$y;�Kkc�D��!2���G5����[�L�A;�g�Y>xt\9/T
��+�R5�Ĩ�#�3��{U��gD]�n�w�����eG�,'Z�e�̓P ��	�)���V��YmfÜ|��vO����im��f��v������/���[ڣ����V-�˹����b�]��5�&K%n!	��x�A�GF�{~_kU#ƭ��Ə1�d���1���yyY��b=��<I ��f�NTD�f� ��^:� u����_�eⱇ'����26�FK�ڱg޻�|q��H������D�Y���2g��H�M��w��Eρ���׬��������1�"��4~0���L���b�L���^������%�m�CI$���E��[P(��V�KR֧x<�#0S�\�<.�`�4������NO�"1Ҙ���f|�`�Fgt�x���6���׏K	����â��y3����6��Ȑf���&ρj��{��-+3�%��)�:񛪡�����zU�mM̰�JƲ��)ś�]�`�\2�nz̛��1��z!@�f�8و$����;��%��֚ɘ�������MR�@��ll'�	T5�fI%�v�����m^�h$ǳ �@�]��'�!���Q�p�5�^�N]�wW�v��'��$�v�q����D
&k�Ѥ��Ǟ�6�����^�˼
ܨc� �/�f{FT�yA�������Z�c=
�Ǆ�~��Y�����Փ��2n�aƔ@&�:g�5z}��T;Ñ�^'���mH�O�y�'��Xկ@�MglsĐ9w�6s&AB�����aqh�P7`OT̒	c�y�`������g�X�D;$+�dK�Λuvv�w���^'��@P�0�N�0�v�-ɮsYz�!8�Ep�\Ԕ�0pe��O����I�@���Y "m-~Ȓ	9�M#��}ߍ���7�^�g��Aλq1	�-^+�7�<��7v�|d�,m��$�T� >��c}x{p����g7��+,D7�_�� �疘
㰺=��ס���D1 �9�.�%��CD���N]�wU@�w��dvv�������I�ˆ�k9�Pd�j�e��:��u�ڗ��{rk�:x��	q=���)�u�n�β�*#�q�x�(]����)y�OV�w.B0J���\	-7|����*��{B$��6?�չ�x��X�펑$U�@,�s��u�Ok�t�ρ����U:W(BT���ű�J�K�ٌi$�"�B!�s�Qu�E���s=�{���@���C�"uq��:�d��<�U^�oZ�LI�J���^����SQ@���|]�O{cW'���D�Kr�/ו4�<Θ���n̪9=��'�oX�x�E���8��{�K��h�5�~V�r�==��x�=$�}��"s�C &p���p��s���U�jD��D�th�C=lt�m��X������tk� ��y�,rZ܏K�>/.L�0��}u��_m=�x3�F#y�Y"�˵H:��g��Ι�g�=z�*x�[*�M�����d�����������-E���rv���:�U&�\�ᢒ���f���x�E�Լ�`�
d(ou�e]��c�NX�Z����g�z�'�:�����B�����طu���q���l�ș���Υ��\-�U��۞�Cn��h!1ӳ�cQ-�\�W6�����%�cZQ�\���!!��Ir/R��;�mi�.�+R0�8��{&�t�W��U�)�]���IR�6�V�e]�.������dݧmR��\[�4fSiL��Q��׮/W3	�#��b�зKev�U���-j/C�9Ƭ߿�����[�/߼
��J�4��|z��pw�W�c�yR���Ɏ����?��|�۶XP��!H���k�{�D<=��p\D�[+gD��PH��GUI*��	����[�/9.K��;��b5�5���g�{�&�l�ɹ���:�P2Gz.D��;pj|p��MP$]�pH��e�0k!�D����6���9f���!^������(.�ȯg=3��cx+�|{μO�^�t=�т�a�(�u��ă�p���7�GKQ�L��\E����ֵ=��r��m�3��c[s+�=���Is?����aӼBN�GCpXg��̑7w�$�u��·�Y�N|OB�q�3��ьkn9��vJ�rsh�,����߻��}����VS9�$߈ �u�
��Ois��e��H� ���&��vy��wG-|s^��lA�СOJT?��E�,�31�ێ!�]�P.�,c�� *�WW�R�^V� �m��SÒ�=��d�n��4�u7���˘�,ޑLh�`�R,�x%"伂{�Eu՛��M������2LHy�i�[�СQ�<�>9��Ǽ�D��ƧB�J#�=} A �5�YT�)��P�7�m.oz�f�1po&ZdH�ܠ؁��׫$���?��Mk�3,��#e�K�-�Ѱ�m��W�8�S ����9Ϗs��8��9-ύ��P�3�49G�A�EM�;����x�g��<bIz�߾���I,�^|��u�����Wo"�$�$e;�m��$��[<�2/}���Nn��O]���	�<(P xxv���Yݩ��q��c�Y��1#=ۀ�����������и������P�T�����էٺ#�}�x��ۆ���Փ'^n�ŧ:>��11!�$R�8ɑ�o�d�~B)�{�@)��Bh������9g�$a>b{!�@�2wT�l�R�U��&�b�6�Y,죲D���yओ��9�B{`�}��#�}F�/��x�i�4��hG�zd�� �;�G�:O�a�ց�L8l���#��WF�����UםM#�X7(�߾��k�]$}�9}���q���|����O��HG)V�d��/E<�d�x� 5�`q�`Q�T�V:6�A �pU���<�b�G��3�Τ �bؗL��>{ϻ���G����^gL���<:Nj��y��@F��$��~�;�W���b8�>d�7�A#���Q	�(�Ǝ<��|.9�0f`,I#�� ���������3�;ޅ]�ix�W��`���]w�C6g=�И�)Q
w�^_<���{|˲J��uSw�@H�� 8ȏ�fU�g0��ߝo�-�r�j�,Y`ހ!li���օ2N�J�U�t�Rq�������^ ��)(���7ln�n1�����%�,�t�)�	$����$�����b�:�"X���ވ��Dj��C���3�7s��9��m��A5@�t@�1f=]lE�A�>�\����ۄ�f�|9���˪� ���bg	�n���ꉻ銑.�؁�s��xs�{α��J��l�$�s�@n�X0����G���R�//�Dz*s�@���[��ޣ8Ox��w��L���6���s�}���_6���^u�j�s�9!o>ů;�� ��8	�qo!A�iBW@���X�WP"E<`IЇ��,L�X=&��ӪOG���������>�]�k�aw[�W� �G�m���n]f�ۖ��m1���� �G�)c��ԜM�(�D��Ʊy����]���L�x��pQ�Q×f�n�,�Lh�k@�K����\=����Qf���̕����lV뙬Aݝ�e�V��q���X�[��
υC܁vw�kʷV�?���V���˞XR�N^�:�[�5�9�'mGC��4�-mkIf��Ôv��Gn6��(;�L��l��m���a��<�.��jH9&�z�YM�*��,h�6 }�~_Pr�j�/�b�����A�{z�c����m6�z�e�2
�s��t1:�RNK�-��b ,k��f�Y�ױ,s̖y��[鑌�=�	GT:4{��>���6PP�	�B������搓$3��زlz��M=�m�/&N��$����P�ux�d����G��*oޑ���.���$�yݠ,c��H�Lt\�P'bޞ��۱��׹��û��
R=�\}I��#Nm��=Br	����L�mh�M,40���^yJ���I']Ө]E��\m���vZ)[�y��m�셹��T��d���86��xz92���~�J-6��Ơ�v��E
��^�7rEN�p걼:g�H�y0�;����zP�5��/>�L��s�,u�G4N�5����a {{�~��?~���A%{{��V�\�O�oF�-dZ�,�A#�X�$6�V�ķ2��w���0#]~��2�=c4���'q�����Y�dˡ�m��'K@<yu(�^2LO�r�����6��`�H�xpdzZ�{�����}a�S!et�����ı:��;��Uv	��`�k<��{�7AxwBȯ ��$	d���]yZ㵏E��G,� �%�s	���d����w����Ғ���OZ�2X�GNot���w;�.K[��lu����<���9A�O>��� ��^ı҉]p��.Cϣ�ɚ|�� I9y� �Y�O	;�t���:�����9��r�8�4��7�hI'z���~2b���vP�;Qz[�u�����w��z H~�߆	�j��~��X������H-��=�ޫ�E*���*nx�=�����Acs�ջb�����n�Q6�U�ϧ]�W�!)�􊻡��{R��� M�R�N�rǣN�[��j�?n��^��m{#�aw�^8;؋�=���Rr�Ƚ�+z3�:��j�����M�Gs�o���}��o�k$��lɍ������]�����Ӻzhe�k|D�K����3h�Ù�w{P�ޫY]��I��|-�4W��|¾s?��f�R�[����a��/b��_L]�#sl*�O��n{P�uG�nC�{�{�A5��wź��F��-��k�]`af�$��3F_߬�������zB^�ٻ}���|¼��od��{r��{�1��<3� �
�0<����O���	{;{<��{�d����H^p���ʗ`���r�z�����1��;}�Q�:zO���V/�姀�߇a׽���䋢�k8�8- _�yZ�dC��O�1e����B�냽=��M�&�w]î��ޫ;��=z=ru[�˝��-R�O���5ڪ�Q��I�r���
��t����Gޙ�Æ�ܹ�y^:�Y�5Ǒ�];��Kݴ��F�K,G�!�t��<2��Ӟ���`�<;=����6�fn�ߺ�(����>�����v�sO�b"W(�%2ow��J�zl���B�-��i��0A� B:m
�~-�G������!<rw� �<g����������������U�0���D9c	D��`+/�f/���e#V���;�q�G׷���~����������nJD ,���e��<��?W(rǎ$�H�hM�{��yg��{}q�������������k���+���%V�V0�!���;���QEu<�b��׌��{}q���w=�e˗.[^&�&�'�bc�AZY�@Hȉ��K�֟�) ��Ðz��Ǐ�����?u��������z�\���G'� ��&$� �9�C��:��zJ4 (�Fs7�y�=Y�L�y�s;��sYr�˖[`��	H�:�BQ����A@���
�^`p HO�@� ��w��P:���a�~=��la	`�� o�R	2�2:|0BJ/$ u# 8�!	N���9���N)#< wQ: DH ��!q)Ї�O�g�`$2�L�	bFw�p5"q�]�e^�2N|�;�#��%�Os�������6yt뷲0�+���쉟��8w�A"�w��{(�xpy���xkd���H������^a�EȐ	=�����m�d��{N��`${`'p\����	Ӛ�Y���܏�&�d�i%̖g�������s��_Oo5��b���̐<}
�Y�ƿ�^�4I�d�3��;��"r�4��k����ʀ����[iW�I� �dA"�Y�]ɽ����Qa���h���؄�S���\��h9�mP7� Cd�N��ʟ.�]0$��q�]�#w(P�u!UM�>W2b��L���Io2C�qbD�����:�H��Utc�Y��O�Np{��8r:�\Ր{����}J�^#k.�wGw���[ �_o�u�v䴟�d~��2��֧%?CD��2N|�;�N�N{a��ȓOw��/�^˺1-�y@6�?D�6Q�ޝ�_Qy��&Ԝ�܌�R�7[���(��6��x�`�b�SB�hF�n��7�X��n�� ����}|���2�D���BdYTz��3�|��1�0 �,� ,[�84wq	���0��~��/�0�y�H�.�g�L�l���`G-J�8o#��&/3�'t�8��� z��>�%���EKyV>���W@w� �b��^Pa���$sF���	�x%�d���߇������y���;:c&�A$�fL�u�ށؠU�� �(i�@��ue��E����芖�3�bZ�#z^	c}}4���	�٦�*�>��N�!�ړ~eu�=H�yN��D^�Q�2��o��y?8�k��=�G��f�ҋ]�{z�w��k��g�ھ����g
&�q�5�֔$=K9�!%���h�u�M���0e��0�sJª��\�[X�ɫ�宔��赜�nahw=��֎��w	r��t��ak��ZVST�:�l�ei��t���9�g�ǳ��`��Sdk�,�4�Rg:R�X���qٶ��$���H޽cat,��f��),�1�8 ݩ1S���u�1l��{���1�f�X�<l��	�UǬ;f3�V��!���";�q0V����Gr9#��7|1�T�&����:�SH����(�嗍��x�"=��@-=��Oi�Rw���T��rƯ��"����A��v�Te�b�o�]x�����mY�3H�
�(��~�H�F]����P=*��u˰֐��\��%l���>�r�~��	�N #��zbq�c_u���%11'�G+ti�t{y�]׊_�Ɛ)��X��j�v���ɵ�z""�S:-�ܺ:����� ����A5{��컥Ġ�s�#0�pS��{vu�8��FG��g�r�C�y������&읞^�y���%�>�z��UT���^��i ����I�DL{y��d�����frgVEX����B+/��ͳ�N�_�}�b[[��z8s�yާRDە��W ����Ό��{=2�3|�-��;V�g�N#�2�z�t�l������ܝx�vaŷEI �<��bw�Ѥ��3��׆$��qNVy�E\��,���;fI�@2��뜂G�3�ү�n�w���Ngy��x�[<�d�A^�"�HB�}s�ӛ���,�\����`�n������~u��~��Ҩj�gGb"woX.�;�$�� �c�B��:츐w��qC�Eڗ�%{� �|z�C�wqj�bz��%|uhw|�r�m"��u���m1�t��۞�^�n�H�s��:mH��O��O�U�G>��9eNd74#̑e��&�߬=M��M �-��y�M��x�R=걂��@N$fFNL�2�������ggֽ� Z�rȐI�y] �Wu�G���9�:t�h��3�PD�9F� ��oL݄�+�3�uh�B���|����4�3���Rwo�M<7��yy�Ӕ�@2n��ޖ�ܽ$�E��>,���r�����fC���{��X��t�$w]���N"��"�uLzn�㝷18c��m�Lߜ$o_L��-w�g���۠�
qf��X�"D!EQ9��1�ȑ���;������t�[#[�ju�	�ޙ.��v������D�A����u��ۆ�ZY��i�%�pE�A���(�{^N�:� ���y�����(��9b'obq����E7�sSYg��(bO_dI<�������)��Y��=�}�r�A$��L�S ��[�� y�y���H�dҦvW�$���Ѣ��B.*��ՕU@�G���f=��*z�QX�Y3�Z@v]�1�7��$�+��t�����VkhTc�ɘ�O�05�	$k/s���y���lFI>�cɻ��a��rs�8x������=��6����n�����q��=��ӣ�0�+�xq�<�e�E�������b�L�*�:��'n����Ek٦<nח�s�{r�ꉙ`y��ǯa�4��|�,��˿w�4&��K*�;���:��ˣ�0��5�ʩ@����%�� ��o�ƌ� <@"p&�e�$� ��@�C��w{���vE�����v�E�!"��Bڽ}{{��{��H$�q�!�yC�^x&$-n3�,K[�:�a�z<9b����r72K��{�m�Y�)�!�	:���Wv�X�xx��nTth�WoF���LLcK*4ڷT�$	y�7Yyꎧ��y�:Y2�l�U4Cq{a�spBt�h�ֱ:�XvvF���;�z��.A���	t���jA ���!{w}�.����z�g�ou+��iv�������H��B�{�)����[UՌ�R=����[��Ä<ٌd�1C�z��_�:��Ob�
h�N]j���Y��{a��"m�R�j��N˸��i����lW��̤VaR:�"˶�O+D�ۦ�urMbru��/kqW�S�v���^ŊVR��AQ���uљ{�����.L�D�%<��.Zۥ*�۱�5;\cg�`w0k����`5u#bE�����n�i*�1�� 1ډ���mlV	����&y�eT���q��k�ٍ��K�֤f�a����]hLGF\����=���������P���>�� �ӗ,����@e�YRe�����$�q �>�C$%z�ٔ=d@x�D(�k����3�Į�b������O���v힙$�g��u5��>��)!b�is�Mi�4��Gϯ��X���V���A2��Q ��8��~�
Y���w�\�>6��a�g>���.�Y ��DvԂ��uG^�>@��sN�_%�ݮR[j*�K�R}l>��b9P�Y>��Í�I�ތm�1��۪�w�r��|�C��ѩQ��\�Ӗ���o<;s��îݞѷ��p螚Se�h.����ҵ��Ɓ?�4O���2U�q �2��|�st���e֏�H6�s:�͐�����;�*
U@�x۲�ފ��(�"�)��ߝ'��y>�=v�_oAgmd¹�,�.9r�?�~+}�znl���>=�![}�}����q���`Je�+��2@왒L�]�斐X��md�:�B?���F@!��v����Ld�\�7���Yw�=���[n�dކ�3w,��a� �TǌȄag>HG�NNtscM��ͨ�A�\���P��*ݵL�D��諏�aaK8�{,ʃ.6�vÞ{��^f�NΖ�b����k�
b��r�w)���޻��pRR���ISUʨێB�c��<q�2������Z�7�qd�[�������� �Tp�o�B��C'� �}�@�����	���S[y��z6��{��/n!)H���3���em��竍�ۼ�̐$��X�踑�&�'�k|	~8�a� ��H;�?�6 ö} {��N�ɏ$���,�[��M]������<	���}�-3�������Q����Zm�f�Jm�l�X i�n��k�i�B�� �#��3��Q��Ht�^y��{f<=��ݺ�s�1lQ!*�Iƶq�Q�R��>T���_��V��a(;����P7`>�r�]ğ.�:0{���@#"��(o2��;���;�Xqz�3]�>�@  0eDP�d���B���#���#TѶ�ZTeе���K",�,i�w�y�����Q�0I��$���w���i_���c�q����cw����<@O ���H3��!��|��o2���/1�0|�ښd�����ꊸ����>D=8��T@G��%���<	h�t��G��L��~Q��;��Iki��:�à��h�z�mE��911�$��t����cw�jUwg���_�������y����/r���y{d�=�b�م��v-�}�P���\��.�ɫoP�K���V��Y��,��	c3�W�"�I �X�H@x$:yk<^� �Yq���ݗ��z�	a˵A ���.�!�y��tH��S�ʯ(�P,B�����r!/g��Q�5$n1x��R���p���`�m]�wm�(;�Q		a����M{ze����]�I���P��y�/t[y�iɫu�Ø*=@���2���fdk�g�,�s�ȓQ�����t�;^r��r�x����ldQ��S�2H#�����x��������sXydy� �v<gzϑ���x"�:u�{4���H>��F2G�n y����>t��#D��S ��J)�$��p�!��AAy	�]c���5�Λ&���s����|/��}��������������#�U^�DT�s����"?�N����PBy�d�� C;�b�! �!*�H���� @�*���V�VV�Ua B@	�@�S��(�J
��"�@�!  @�
�H���;D�	B!E�E BDT�$QH� BT�	A� �T B�Q � $G� �	@� � � �BX��C�� J @��J @��B @��P����! !�J @��J @� B�@� ;�:%  BP$  BD!  B!  P% 9��!@2�!
 !
� B���B u�@!�  !"�!
�!*��� 8�%  BP   BT U�	P� �@�� ��q�t|��_�����0��-" ����s��������|�����?���������_���~���Ⱥ��?ʜ���������/��_��?������/���� ����~2��K�4���!��" �������S�oi�A�C���O�������}�o����\�oTT@
Q
V�V��bU)�)F%J�a�J�A��T�R �iRe�D�FI�"@��&�T�A�D��bD��FeJ�RfD�`�I%I%RBQ�H���b@��)R	R``HF`T��!%H�b��H%HH I%� `�iXFRT��a H�&E��&T��$��"T� IHBQ�f�$	$IXB� �bT�dY�`�dIF�E�`�`F�f�F�a	RXRQ�T� Q�Q�Q�FE!edY�E�e�$ee!V�� �"Q��`YFe�dQ��%%HB�Q�Q�dX$F$Z��XBf��`�h�� �hT`	VQ�X�bE�iF�%P�V�hVB��h�d�I!�FIT)I�
bVI@�bD��JDi�Q�P�PB�DF� ?�! 9" R�:�����w�?����UDR�B��EJ����_��?������`������T@z��_����`u�����q����W��g�E]��'�z���"�*�DW��6���E@^~���%W �����8����t�ß��?G����:�;@o�������� ����P�ٿ�?����;�����$������Q U����8� �� ��?�!�RE��S���|O��?�O�h=����$��|@|L����������_ �?��}}_�*�A탁������?������������d�Mg���v�f�A@��̟\��>0�@   
   �

 @ 4B��h  CF� � ҉P  � �5@Pip���P�  �S�$D���

 m� AZ�@�Q@(� �J� V� �               =      P           @          @wϯ�����&�m��8�۝����gF��� �s��m��Ջ��95�˭R �Z��r��8���K���iWzW�nګ�u�/< ��9�w���=ou΀�g�`��t/0С@������zs����+�y�)��B��҃O9�y� �x� 
�| �K         #�)_@�s�:��^`޳�
o,�F�M���(� /.� <7e�M�5y�h���4�/{���5�6��M]�)��Δ�8ƨtԹ�	Q!Z�  /{��T�X��, T�L�NƔ���F�K�������(N� Ҫ����Q��;i.A���tԮچ� R�*�  �z   P  P �D����J]5N�5\�J�[9�JT@hT�m\mQNZ�mY��Wc5ks��\7 �BK����3I�(45@	x  �:�1��Ma�R�B� ��T�͝�\��MT��Ɣ��p ,��-NƑr�;�����ԩP��
���{�  ;�     P  G�&mO���^Z�����9���.� q���kU��ٛ���Z�Z� �P͎@��:� � )/|  ���wU��\�p͘�������k��k����*�Թ�媆� wS����M�����esw(F�']h`
� (^  �        �zZ���ֶ��p[5���jms9�Z� ��.���6��Nv��6��B�Ӏڪ�n�p)�ʸ iAH�x  >��;6�4��hj7 �V�\�E�;:���\
�g6�� �%�v��U��9��i�7Xu6���JR��  E?#)U4��D�2�S	%  !��?h����   ��JJ�    �Q5)H0�~߿��g�3�A��xo�m�j���i@(�E IN��o�`ILHB!!� IO��$ I?�B�!������/�5��<��3��8��)�af��x�n���S��ܺZ���W#��2"F�Z�BH�m�ջ�ꛃj��d��K��M�g+)�L���@еL�X�92��t��0�`�"�o7~̮شЊ��-��1��l��[U�'���9� N���Q��me���R�[�JWj˹@r���ҫ:�-���웪���]��D�,0e�1B���
�(�B�[5%��V��^�I�:�j����aF���vR���wu]��`u��z�jT�t%	��0��v+h^�4P����ݬ�y������ ͖q��c���J˰B�[����m���D�#[SQ�CR�H^��5�E{�[y����2�Y��x�%�a�=z�S��u3%��oj����5��o]�*�;�t�WI������P�x�?GV���B�5�͖q�lk� �l:'6l���on�kh�5���M�*��K%�P��b:���&��J��Ê��S-b�-*u�Պ�Ѭ���������%��AV�@C�j�%��K�ǩf������5�y����*`��((e��B�ı�ڔu�t 
:�ۖ�����7R��Wwy6�`�/2�YV���b�ݬQ���:�5mn���n���][w��Wn�Yփы>X��.�wmßv8���̫Б�5ؓ��%��Ȅ�E�h3�j��!���m��/,�
�0!����]��W����vR���,�
"�Ң�7���z��Jq�� $(��m-��,�Z�7++R�ijH�)j��@�W����N��-��S��/$wj��5�ov��x&nQ�.���%�ll-KU�ce��9H��f�dML6��Y���Ǒ�'�2�\bM��!����@K͒�ކ�k�(Z�m��Qܕ��;�(�C.���l���wmn�ƭ�KNA��m��t�Y%L�È���F�+o,��͑g0�<�l��M�ڑ���\��l�97C��Z�[��4��F�b��Z����ݨ)�ׯr+voẒ�lx-��XU�b�`�zFS��P��M��#p�%�ݟ �%<ޚ:��C�+s:&]�ԤMFҨ1����]��K�Я��Zwv�+�{.��C6�����v�3�P��9h癄͛�u�̄�	�oWG���X�e��␝A�j���"��eJÁͰ�F�J�%D�.���eKj��2G��
hȅ�jZ\h�y���⦴�����ia%x��جlz�ʵ*s&o\"�r�{�ȁ�lf��b�L�#mWm�G�N�VEʀފ�V�v3k�1�a��
�ƫ:u��kC�N�U�kV�n��5L^T��SxJ�FՓ9�wu۰����`�>܎�����"���4�:�P�+]8�̳I���?�n-\�vP7�ȼ�te�C4�
*Q�J)q��PL�҂�j-��wQպ8�˰om�������z-2�C��l���F41��
sjn+�Ӧ��Vk\mD텆8���;�n��ץ���l����Z�:H��@�ЎL�	��(^5�H��Ţ�ޙ�c	�7SEܤ�65^튥�n�Ղ�o\��n�^�H��9��f�Gv���B-b�2�f��&f\"�,�y4^�Vl\�fU�y��XT�%6U�z�ӂ��X��N�L�������&�n�d­
*��ܖ���&�J���%�i�Bш���i|V-`-�Yq|�ᩚ7@�oE��{G)Ce��86<�2�30�ݣbk*��%��#n]�MB��s1A�e�0:�ߦ�8J��fێ�o.
M͸�&h3@5��2?�;Kr�f�N؂�^�FE����%W�%wV1ڤ��eJ�l�T�+2��w��z�ݧ��ci��Ql(�n��35V�؋�2�jy���u{h�r�t���3opcSK�m-ܵ�ݤ�d�x�oS���њ�AZ�0�vmԗ�\#��d38�7j��"���o1�5B�����^�Uޔi����*\t�*5�S5�h���n��K�$�rt�oon
��3�P��b�٪�S!��[ZE�up��̅f^�j��h�����Y�xpV(���!س� 7Glc��J��k{�@R$pŗ�,WQP�a}�m'��i��EY�L��Xj"�V�o1Bhڊ�Sw���Օ�h0V�����+4K�9��t��k;B�]Yzcɴ�]�.��ѐ֥k5��F٥��,���U�)�FQbޕ4t!���+��!��x�3��sX�7.+�%�)A���s�Z{L�V[u�v ��x!�i��ht.Yܩe%6�!�5ڧp��j���fգy�oV�u��t|��?�

�f�w沝�8t�i^Q�)��{gov�-�[N��ʺ�ઓa��U�O��^:���}PY����9�{%.{��cx����nf�z.]0�&��(DF/m�26��×Y�滗n����v�x>N܆\���ې3x����J�߄�S!�¬��^�V��n�Iω���ubC*�y{`h�UxԽ ^fܵL�we�
��9�Щ%�Q;�,�ax���f]�#I8���R�U�v�]��V�v�5�� uem엱ǭL�̷�+7�X�ڮ�ڗ�.��KqO�fi����i��k�Ӵ��+";Zi�m�[�#��Ȳk;N[ǥh�¨V��,����������f+T34��nf�YW5,t�`��-8 ZK��.̓f��Z�D��P$V�ª�X���XU�^�;5 ͚�pۤ6ʡa=�񱒜����ܼW%]������8m\ݶ%�5sF!.#&�Ov��mY�d=��S%���q�Ѡ���=�yFCj�Qܒ�ayZa-<~t��
�T�m�-�vp�r���<b�Ch2S�Bm�&��l����N���a����'�]Y��8�r��;0U�n+-n
�.l5b� �Z̚ۍ"ҁ�𠬁�kr�З��C��f$�Ison�ˁZݫ�z����TJk��]l����H�����r�6�C�5��d3gs���̳��F�f����$���,Z�z�%/J�Ĭ� 
�E�)DMDm1�hT��E6��F����Z1�ZN� k���s��ڼ��ݸ�����Ȯ'b(���ذĲr��ʏ4�M\ى�1�EBt���1�jz��œ
�D;jC�:�{��ŧ�	a�k7̺�d"�&��{�a|������ȱ�-���O/nfL&�]��nB�ܫw�Zd�Wim��
��t�$�y6j��dm��p���rl�g�FT�~�i�vwo2^���oNn��[c���̓ڂ��KVr�зl̢����RG(-b��k��.�>���mM�xX��{�����n�3rmM�jbܔs.�"�U\1���2Y���i*��)7K���%<�vv����.#{����tĪ
"�@Y�{{�U�����_�LF���s��M�5tt,�����������v�U��NS�fnLn��Vi�_Z���Ui�x��0�Zo3S��nub�weQԭ�S6��nҬn #Yʲ��{��p)#�"��s��UIUV���!d�ɥ�m�Ym[�-:��������@��T�����v(uy�h��fmرWvΚ�AS�AL�74�tj�y����GnfEP+ �[Z8����B�N$�
7*DF٢5���NԼ[p�0��5�8^�zLޠ�ɵ�����&9n'fPVuɄ4R��ܩ��-ԭؐ"�YG6�)3�zB)0�L��+m�͵V�|h�a-���Em#Cɻ3]��l�*���I�|j�mZ���	�5���6�M=��wE�G�f�в���vl�M*���Y[����ʺ:ܲ����<��yL�yJ���ݖ��	�u�ƣ��F�tfѫ"��{�U�gukñP9L{�E�ʱx��
6���lh��i��}�Xwup�sm@��lz�ŅH�Dc!��Uެ�6�ke�����a8�"�kvٌl 
ƞ�̙5d�n`ω�Ttf]J�x^��f����F�m�:�bK��D��*�l�oY�݌V�n���&ɘ���I�S���kk����v Q1t�n�i�4;5���caB�R���7kw`��k)c�+��faSIOs�D���h6*j��6ԖL�A�r��q<�;�,f�1����ù�Jɍ���7v�u��3vo) Qq��0��n^αv�9�G%�2:&�v���V[f�]X�1�/ƝK�v�����7Q��*n=! �N��fKeZ� �b��Lt,�L5�V7 $�Yvcτx��ݡ��s.CW�lR#2�ډ[�=3F�*)*6��Ɍ�1̓.���cZ;��V鷀�Ǹ5<�X���2��m@r���B��� 3���J��â�p0+6��f�n�.���Wyy���=�JY��L���Y$�X��w,f�TTs6�5%ފB()���{[�,@4��x^���M�d'�M�a*�n�A�L^MGM(~Q��g��M#,�w�5=F�5z��ܩ�v�T�ٻ$$��ܘ�4%P!LA���y��E0�N��R� ���Ż�����Iw"
�O����m�r�[�/r�=�����Y�ͽ���ə��\>q��f�-�rո��8���cX�aJ�M�ݳR�*� �o�cQ�Т�4lg����ĭIm^J���YP`R��wz��� lÕooo$����ñ�e<Y�U�#Ƭc�O�׻�krͱke�p]��vri0������]�e�T0�S��:ӈd�Z�gk:��Sr�+j��2/&�[[�*��M���$�v��J�f+�6�Z��vL��<Dl߶YOMK��2�`2�}gEޔ��kX�٧D���Hg&Pж�x,6��Y@e�HTF���0mH�a:*ֈ���1���۽�gu��63E�7qῥ8�,Fe����eR�^�b��A�z��.��ȼ���j��(�9/]��IkI*eLNޙ&��$䧬V���m][���Ԕ��<�Mۼ�xb9r�C�f�a�p��Z����� Wz��NY�0m�ӛ�/re�5EiT�5j�Q�1E�GĲ�ә���`�S)еLf��ģ�i�n�0if�X�Ϭ��l��7�nP� ��+��>������r��L�(V�A�n&�4��r� F:�Mܓ����ɫm)�&b�w�9�\����Ĳ�N\t+%[?����7�5A�E^бt�e��ԭ;�at��>�p��-ۼ4N�R��a٫"g=+lݜ�r����kc��B���6�����ɷ*����Z�9�d4��� ���oh�)�6 �T1&���� wc7PKV+1�J�b'���#Ro|�Ʒ�rfr�����E�vaY�Pv1ѭu��آU�=f�^�����*&Y��t��u�]m������dG5�d؋@��Uw�v�ʵT�ӥۛoG3�87�m�u��Qw1Շ��rT⩲����[O$%[��Ā�L��Nmfi�.�۽+�+Zr#�FVYt����qrLB�2���d7l`p<�]^�R0�.���:�f���[flWd��j�uwZi5f�ph�A;upA,9DK�J$�J�t���q�F��;ݭ�C4-��?-��=i,�*��:+^��fM��B�;���0�����hڙ�!�w����P�Mm�ր�)�9,21K�(���^krS ��&�*5�/4^����]�K�p;�F��X���7*�$��UFh�*�T�x3fiU`�	�$7���a�LѪ�D�rk��n�]������6����S"�i���w��h���[�Jɥ�AX�`NV`����<JH� ��.�CNV^<�orl��	��[�wi�����ڼ��!1�o2dCԮ�5�6�
GFaݬ��`̔0݁����l�y��So^V�u>]���RK�ޔ-ǗF�o4R�`�I��LQ�d�ךhۗ�Z����������(��K6�kO\�X��lm�'�a��s]#�r*Y�U�O2�ǘ]�m�.����"��L��-e�Aݜʰ�9�f��V�a�Zy�e ���R���EK�m��e��@-���2�M�����n��&m(&�Mj��L)���`�M�+eŊ�8"ƒ�a��-ww�:�in�ȀwX�7YQR�$GE]u�eƳ������#ϰ�"�5�@[Wxմ��n��U�1aYq�)�wf�W�{V U5�muj�f�\W�mi��z㬺Ʀ�-4�v�k(@�.V�K>kf-vva:�!q�5j:�t��غ7',m"��$RE]2O���C+k5XB,{6�Gu��#Y�Y1J�I�����]���6�Ǡ��
�u���f�J��ѩV��t3�$�K[��yW��q����y,:ݷp�, ,bN��B�P�GqYyHŎe�m�4+qǷY�{��j�6�U�rd|�kU�r��9b��|9I×/Q���NV]�^RК��]6L�f��\����z15����1Xe�ԸI{eY�� ˵N�����o�ff8��m-�f�m�'�n�v�dзBۈ�Ř�n��������/l豕w���:G)�o>BR�N���ޛt��ut����ص���p�U���2�ķ#M�74S%��0�%�����sK�K]ԬMO����SY��eW**��Vkv뗜�w�R])����<�2��;zr/�`��bk
C6T��X�i�1j.팧y70�Nj*�G���Ug�vV�57c/7@��I0�h��ҍ
 �U�ɟ�ֽ�o-���q����s>�C�A=1�ْ�j�Z���dmO�t@5u��"J�H�z��Z2�vS�uůH���,�xj�m��R.$*��.*E��s;�q��mM��wp���+�<=����z@��HH)$	I$$I   (@�$ (I"�R� ,�$��d ��(d��I E ��Ad�E! Y!��HI����BI!!	d��	$R�a	I!HJI$) @Y� XBX@�%2I�RQ��e��Q�VuvwWՐRHa SSBS� ��
d�B(B ��PXHS$!L �!BAd���H(B,�!,���X�BB��@! Y  QIAd%0��I"�d�� �Jd�)I�Y	 Y!�
HJd
`H
H
P�R�)���$YS!	L)  SO��BC�H@�s�g�?~3�E~L��z�j��S�;{�H ��)
�f�K��f��/�����uln��l�e9�oo&#L�<R��xt�vڎ��S%&C��N.�����V�$�0���Wr�7j�5/.��؈��[�1���ɨ�`ķ�N�@�v*MΎ���4��}v��	���+��ʷh���5�qM�<��(�x����JO6�
���m%Y�;��t�\c���'��)E쥪2m�Xf��f��Q���U$l���|�	��MX�#�Αu��L\n�M��⬖����`CZ�E�䍫}y�I���bs&�v����#+���ʹ�޲'M�P�j���٫ԭ���LY`��'�8e��Δ�k��(�5��0v%�ZV��
��
�ԯ.�%z����,�ul��H������Tt&�2���Y��Ƞhj���˗Y4�h�w2�G@	j�.1�ډZ�#7*�F%�B��5ݴ��H@,`��/�n�\�\����&�{cf�%��/u��:c�.��)�"i1	��G�Gk~{eN33���tV���k��I���‽�&Ya���n��SW����q���t�*1��팤��9�M�
w$�R�%����f��1�[Gg�j���`R2��bo� ���g�p�J��"�[�6�۫�W��p4��ONm��c=���N�\9n+;�ۓ���c�,V�>;M��#�G�]e��CM�97D=��o&@4�1�xۍC^�䡘���.���ɐ����/!��7NÜy3;�C^>l1m�E��ݺ�d��T����P��6�rg3i�V���Q괵������<�G{���Y�	��ëOJ<Sћ��������yukL+�m�q��v!"]��\��X2� �/,kV�O� r��ZuԧȻc^-�Ϻ����F���3C���f!��]�����Nࡻ�o�0��vEґK{�OLozc��vJ��,�9�f@���}ɪ�\�L�6kq����n��Z��s��ݳ7M���\�r�S���m�>W��Ǽ�gd��Q��0�웜��Wk��s�D9xܢ�ؾ�K/q�g�j��\sN�ْ��]�A]j�ɖ�5�ŧ��^\�wH>������DجfB�>y7�ߵ��v*t�7�00���r*#��S��c��(Kk7]�U��ߞ�[)mwm�st�((�8�0����ϖ9�Y�D��̻�ea4�;�*�}�;��/�o좝�F�H�P)EcY[���N�V��X�c	Q#/�Z{����Dkl�c:���5��<�K�Sqɹ���A7v5���X�ʵD�Y.H�F�g������sX4�c�^���G,'��j�y�#gF4p�
1�F7_f��x���Z^��Zz����!qCr�eK��'�9�i|��{�Q�@�/!͟�^��
d��9�o;�1{ׂ��s��%�&FJE�[P"�ښ�iQ��~ͺ�R��eqʼ�=��yqg;����WE��iMqtZ�ɋu�U�O3�l�����xqamL��h-�{e���c��a��}����g���՝�7����0���`�M�ㅤfi'%U�kY�S�l��kVZ�S��cs!z�`���`�/�Z��L=�E�pV�G���z(ܮ��3au{}d���Ŗ��f��vc��V"��K�7��F˩�2�(ǊT��2��n'&jL΃8�i��z�jQ2������Z-��4F�ջt�RP�[�ܳh��K��jE�|�0�q`���aagxP�уdX*E�8.+%�샭j��wn̰��E��STTF1a85.,�Ҥ��1&ec
6B�ͥ��E39�d�!Qy��A�����+�A�P���)H��N ��I�i7;5vFfwݲ�v�hY�^ ��e���mN'o{���������S)Q�;�L*Wi������J�$�c�S��U��3���oQ8(��	�A�"��(�[��3��:5j�{��M��v�^����ގ����L�++�s�ͬ��/wX5���K�:�Cbƍ�Of����a�@�H�!���qu������(<͗�$���^%��⊚��R�[���vLO���r�dܙ��<I͉I�1�]����f9S;k�YApem�'�5j�,����N�6�,P�o�T�����U��b�ׂ�a#�H�"�#6(������p�xY3U�5eLk`�U�p]��w$[SVge��ժr��!���j���܍��q�tP������p;�����Ç%*ɔ;����QAӒ���Z����7F���{��]�h���VI�ZmmJU�0\�[�m���z��d��_�3����9f��nV�!��9�.���K�3f�ϛJ���ՍJ�1r��z@
���=]337`5٘fƫf���f�!N�L�b��2�%�I��͑P��8~&��X�w]�7C3�<$�7/�oZ����>j��z0c�Föc��M7}��v	 �7��i�)�aV�"�[Z��F�%���V�Ln�kFr ����*��#	�Ǻ�d}�j���vՍ�h�2w�հ������a��.�2f��N�ww}O1呼ꏎm�-��`Tkˣެ#faYי��ޮ]�i7{��VZd��|3�}�]�}�E͠K�����v�^9
�W��I������Qu;T�(;���]9�����m�����efЗ\۠�'�\�[/���s�z����f�K����m���/E��k��Y����,�AR�SP��B#t8ֹ�R��.i�����W��!^>}fw]G���j�����Q�8��,���Z��]JQ�]��/8������*b���.�Z�u�Cښٺ0�SzD�^�؞v��;-]*ʻke�L���.ڮ����g��U��[]\�w+ �w�f�%�y/���v�w����˻�4x�c�����O8d�-�����V��B�wXM6�Ӌd"
��S����ʪr�JU0�÷k���	V�M,�[+�܁���[�t�neH����ea�ˑ�f��4�k(LTiS0�F�a�c���-��S�-���lr��nWK���d ���6�lAw�&f�\y��`���r���'��+��kS�ɝ��
�	�!���'�F��P���̉���ݏK��Ψh�D�p��@���B����)v���/�r��pS%+V���.Gf�M!B�l�rGSf�oh��aLw��W��V�48��ݬ��o.<���;�f�����^0% y��9�{(�ByF�.�XB%&k,���c��m��{�(`�C�	��Һ�Ib���=�s1(���;0��Y:�!1ɕj2��mԥ{R�ke��%R�vp�5�qf�w:��P� -Xiʜ�CRpfL��^�w��5��^>8Ji�����v��{:������a��S)�c)�o\Q"�y>���N���Ν�yf��=3qY47�<�f�(����	�ÑXN��:jV_1����;bN��[o�<��zk��n}�#��{�*T�T�g�5͘2a�Is�/K��t=� ]�ݮ�d�ʙC\��j&3E��+e�fb�nR'/�t�m�f�_Y�y
vf���<��,
��רmI�ު�$簋���eW\�5qX��a��;��z���Xl�~�jN���P���M���;IJ9���鼱gE�YBt<��d�7h�/�e�ዦС���Z�e���v��¾��Vi�	��.o��.:�4��۟���t�WvAu�m�L�v��d��AީmX��CFU�C@ʣm�"��2!U&�����GZ2�m�1�ڻ��((3x�u�Xwxb]��z�Xw*��D�TMN(�)֜V��1Nm���hH�q�t!\M9��nUEκ3�*j� ��[u�9����[9r�р�S[�:v����9��k��Y&�I�*�	���l|%BTᰳ�f�k��I�� ��,�-�o�)��%�xef�|;o%<(u_^wVΚi�i��!��y��)\V]хK�q���8���3���
��Cr���v��,�=�e�>�a���oz�r�+��W��y+�x���ޛ����ب��g�7"V�#���(��91qiHnN���*�506%hPm�C,��]��	Bۺ9�"�^��S�7-\��fy�P�qrldީw���f�X����As�ce�bo;[�?�g*���Mе3r)X�������dg4�Z�>�Ė�Hf^���7�o.b$�"�U&eg�'F'��+9���ZgdU�qS7t6�
�J�PK�^	n���ۜ�3M�%D����jS�'R�rL!UnjwVkNڬ�%M�--����k��e��{(�+�N��x����+3fUD��˷G;R7J\��&g%;�Sf��!��rP��*�`�mI
kX15���F�pS��T�ڊ5ur,ALt��Y����eց�X�a�N�Y׸��fV�IY�)�1)b��e�Q�5�y@�_�a�f^�ʼܶ�1Z�ngā��jG\�:S���������K�,�wڰ��W���}�ǉn�m�ז��s���/_�^�Xu��#|�]Lջ������.��f`�1r��<�l�VvZ��^�:	�U���ɨLN^��˪��RMbrh���D*���U��_阨Wx�_B0.3)U�|*��R�z-X)8on�}���A�&��rVeG�� K!@��ج8t��.��Vqy䦳�H��|��̙�[�\�f�J��F2��âR���<����[��Cse~'"aJ�A='�"M�N��{X��u$�w�&P��G(��/�v�m\����E;�i5k��[0=���} w�v�!w�m�#[ۗ�y��x,qF]GS�Z�WI[0ʊ�!����G;������V�8��pZIT綫6#������wG+q���{U��R&�ֈ����s���\ʓP�h�6�15MN��8崪����1TS�F��ôo��0��t�����+���ȳ���z��޷��Y���;�΄V�V)(Y'����®���:�T���N�D:u
�5k�72�c����:��c/�s�+x�Ơ=�d��+hV�ܴ��j]�t7�$�cܻmd9�7+Oob���P^H��^޾���8����R�ڎv�O�Y4o :2�P�:t�|��i�3�,�4�Ńȷ(b+6�w+������-�&ͭ���[�-��2�[Wn;�+v�)�ݜ6ݙV����75���S�"R��iS2���y�S�Ӯ�ʝi�jln�c�5� �S����kD��{fă�(,⒋!e�����;���I���92��8n^[�L�ʂ7qЉsl�*�,C�Ɋ�SN��ɘoYnt<
��ܴ[���N��ԧ�R�̭��Fe[H7��Q���NQQ=�V��֮���	f��Jt��R�)Ւv�T�^�wo,�G^t��8-7m՝��]ǻI��D�^I*�	�/u	�J�Bʲȭ�V!�6 ���t.��N��eu���ѳ���lq�3�8+��̻S[�u��QerX�nA[p��o(]y[c(����g�����*��A���]��J��;8c���br�jR<�ee#���w[�5d'*-wjlܻ/B�G�q��+	��VXlڣ�A�<bR����Vಜɮ���*UTh�p���MIX�.�M'�լ�m��Or�nG���Y�nM#q���ŝ�]v�-;QB�`v�e�3�m���ٷV��]�Zb�+{6�~�|�;t'N��Wk�F]�Q��\�c�KreB�	y���8b:��+����oE�E��{e�h�)�+��h�Y��7����R��9+j��u�p�[���AW[�03�qZ�2��n�A4��	�&���H�v���d,�TㇹW	�uF�y��/^X��6�*��
K��#N3`;Z��
�:pu���k�!��օ���F��Gm8θw������õ�^�l��V�*_(�kkR���+\�S�AO�̜ڬw+�H�����Y���A��nRV�j�y��_�Y���c4��y�ٚ]b`��δ�e�̩��*!n�ժ֠�#�Y�`��h�5�M�^�	����٥{���s9n�[8�0Rg�ث
��F�F@D��ػ����I
S��D��s��(�0s^���NA-����Q��MAgfkO-��ܜ�L;Z|��-�\柎��}Dp;�L�� A[ޮƊ�p��с����g[K�����{,T���:�"p�3��z.�V�ə�Mx㻫��]��'��������Qt�5s�ң��Mn+穬��K�|�`S�+0)Y��nKVF
PL�r��ŏ2��݂�X�m��KU��X �v5�#T�lwF-�����֍�7�@�d���qaw�v{��+�%�	��
��87�,�f̠�w��Q<u��VX�[,Y���z��lj#�Hgk"�pa�5���gi�	'3��tBS3^,�`{���vM�v�Nw5��@M$��Xra���#ܻ!�����{��쥲F�j2��Yy"��vm]�Y�P:(ɐ��z�b��WA���������8���Q�R��ެ�crP���\I����Pl�P��,f����w4�5G]Y��>=w��R��X�*w�f�.�0�`�+��K�eXC��b�B���+�mD�J*��<1Sם�.�uEN��HJu���/%8�Н�/�\�d�}Kz1�G6�,�ڔ��
�I�7E�=�ו����%W�X-��F��-�{lV�-V�,�]x�n�՗�-��/��f�#�@�+�j�CM����<�On�g�V�����kn�*z�m�K3���4Zgz��A�ق�/���r�R�G��9N[WFJ���������.�:���w���b��H@�`�I��}>$U�k�9mvz��n%ݹL]����zNx�[\�{m͗P)��� ܷX����^8zX�Lh�����0�1�w쩣�6A.�ۣQ�N�kv��/nH���$�q�q�M�6�ӣv�.p�t��4a�)��v���Yź�����$%��k�u`�6�2vOO2����vO��(s�lge�S����^�%�ۅ����e����x;u�j˻AsgC��v7/��i5��^��m�ġ���cb�y����X�;]]b���=nm�����y6����Ò��=���_#am��6x���;w[qc[A/7c,�ك�>�������c&1����f*^ϴInݻ�;gs˽���9�b<��.'�S��6�Hgֶ�.;<\����Gõ�]�Q�ڎ��[T��f�m�rur��8<7*�<W��=�}l<�Dr{��s�:Gu� �3VGV7��i;;ָ;U���Z۶�y���	���^�ݛ@P�]��6��۰N�v�m�����C�sl\x�2�G�I�Sۋ���B<Ǜ]��p����w�b��*u���6�˳g������8��t%1q�͇	y7C]�����!��Kx��1�s���ͥlc�a�X��۷/]�v5�#���C�� �_Vv����v}��km��ۅ��pb�]]���pݐ��s�$c���r絹��&����ORn,��NPq�����n��Uv)"����N��ݍŜ:����؇=+�s˧<<x,������$d����kZ��֎E�0�M���˶�.1dۗ�Z�qP"�s�c�:3�뭜�۫�ӆ�&�;�xh��Y���aw����>Aq�ݸ�|e<e�ǵ�|ma�@t��$���#��[�r�8��%�}�v�ݻg��RV9�9::u��N�%F�v��"�;��2�]��:y�r�5�˛�������6�[����������9�L�˭�$��7��6g��m9̍�ӛ�@�4C��yٝ���W\��I��5X�tFx����\Z^װv��#�zg�zp�9aO&ϴ��;�y �k�6�\����CV���p<����Z�l���>8֮�N����c�[�#���\<�:�8$���\3f{9����+��9p��:k�؄p��
�d�7`ݐ�n^90k��]7����joF���ax���͎�iu��8�Z�r]���]��91��痎�9��k�N��6�A��w���i�M���7#���8{�`'���.ݷ�X�
,�؇�����]�i�ZKDݧR!�D��pr�]��ey�Յ�n^����6�.�5��m�<l-��p�<���ݕy��<X5�5d�>n��l�["lU9�'��\v���۱�PE���=�sնݮ�pb�ǳy�������뉪�Հ�f�(��c������U��ϑ0ov��)Խgl=<���m�3-�u>Cד;�i�vN7	۠,٘�w$����qc�zC3e�D�}�͑��H�=�\�,�حuoe���K�wG�ض=^@�d�,f���7x�Qɷ]z�㔷�`���w�5�k(�iv�S�U���hw�nFη5�s��9�`ش�saW-�g��c���%�g��pc��b^նu��#q���q��6���c���.�<=g�u�G���
8�A���]s�u�fBxћ\���e��q��K�v�{;��t�y����f�9�YpYp^�]�wOF�'\����dC{{�<7m�β�n���y�r���8���3lGj��<\�l�{f�A�:��W�ͼx��\�<��l�wGxAۆ�۝�.ṙ�Mm��O=Mk��n=ӂ�'n���y3�cW������Ƌv\�H�V)��n�m�f��<.y3���'Ob�6k�.q#T�o\���E��Z�px�v�<s;��UK0������tl��uΠwgƇO02 ��8��pd2�V�
�T�ݸ�Rd�v��p�G�ۗ��˧��y��������#LU��:Зs���l�{;�e�N���nG�M�c�ГV7�<+��k.�p���;v�7"�#�7>`ۖ�\�y��i�ޮ�7��/i�/Y����q.�1�w"�zV�]��8��N�����ۏ#�ȱjt$��kůvSm���L�k�o>��ۙᛎ{�ۍ��'61���ت݌Z��v�w�0-�Iѷ<�d���-덏h6��A�Gbݢk�����p͹�v͹�q��-4)/t9��dr%��]zQ��	:�3�M��mڡ�������m�[�����Ԗ9.s�R,kZ]��,�f�v��-ch[WX���\��6:b���d�W=���GG4��'OOg�\���.��bլr�k�,k�;bw��75z����vW���r���C�5�Z�H/0��F�ܳ:	h���cA�Ss�_Fkvˌz��6�s˽�v1�=�m��uk��<�8-�cڮ;v{���W�В�u�i���'�M��{��I����<qON-O\1�<�:����禮�GO!��y���L[���x�VH���97e9釶���w3�z]h�Zs��slk�l�v�L��|Ƕ6��+����p�����whL79.������unxw�;p���Ks�t8�z�X�t1��¦R�8��l�M׃.�����X��q��8�Z%8:����h�K��9O2�욍̾�R �c����t���x<�������\=��Q��6���h��Om���&�	���X�'p��b��i%��v��t=\�����\�58�J��=WY�;qv��8��^��|c\�kt����bDBH�T�e*����H��77g��R���1��7l :m��<1��g s��g��zsō��@�k]�E\�y�lwA�c�=����49q���r���c;�V]6�\��ز�7������=�ٶ���z:6�e���{m��7I�u���۱����{<���3θ��PD��ۛH��^�7n���뫎�75�t$p�9L��s��Խ���(�n౪���h��.��ݎ�<�5����/<�ʧ
h���=(l�\k�u��^�m:֋����	�z��Ü��Y�9�5�E�%���*�|��r�\v��8H�ێ�w��fnp��t�]Af%�F��ݴ���I��g=��,yH�|6ϻv��=(=6����6��<��]J47:�v�Jsv��J�f����Ѷ��l�֞��qơ̲F����&sj�<1�6y��:�Ц���d�긘�d�z#Gl%ӡ{xQ���#ۀ=��f�<t��&�(8���v�0s��m��v셱�ul��:x'Q���%ڼ�k��5G"���=�1�&�[e��e�8��ym;s� ��ؚ��E��q��[sq�C��g����v5r�v��h�[n�R�`H��'n9��n���ܙ�z�.�rum�����R�0X7/s�,O[�r���ݝ�&5T+�VN|f�3Ɯ��m�x`,�9� �/C[t��8M��v.��R��js��:�Dnw����k-��phr�q-�l���s����v���70�ۛ<��vF��Я���eN݂���å�uG�7���NP����OBQqۋ�h:T^GNK[QN1�����v,ܧH��ǜ����k�	����э�1��SCӫ�u��^ۜ/�c�9�v�h��:�熡������A"�{���x3��ykY���]ᢌ�J��<���c�Z�y�M�&�6���[�qǝ���=[/82lwKע���]�^���;r����uͺ�nW<2y�)��ms�����iw]�zƕַ=����:���=����:2u�`C��(�{&�e'��sv�/�����f��͸����\�n�l�n؇�
�ѵ��,�:�lm�%=x�3�9���w�����F�z8�M��b�Ln�K�`Y����.���X�53��ѩ6���y��Rv����'�%�mw3���8�u5 v�Ξ�}�� V�7;ul��:���v#q����y�[v��wI�� s�:���{t���&9fH��������֞܍�V�]��$��Gbs�f�O%���[r�V���v�����/3®��^���o[2p�3\�<��f#Ϲƶ���w�-��v�#O�#�;][�w^^9�y,���6|��.�l��v���ɭ���rmi�3غ��I��n�tri0�G����n��K�%W\l�XU����V(�lv�5ʞ���׃�����m�<�\��t��GXǈ��:6��]��ܾ��6�k��Ѷ�����:ݸ��mnzz�k4�x\���"r�4�\y
�gx.B���a]�qe�kka�)��q��uO]�)�v	go}�͙�3yi�f|�[I��*�썔ȁ�ĩ���(�3�"P��p!�w]v��U9}�rYSd�|u�(����z��{ݓ�*�:ɞue;Wl�Ų��w�D^�1c`�ݒH�v^�Y��x��9��}2s`�v�c�v�ڗv����)��Y�����\
�;b^�=l��g�c-��%�qk���;-�7jBN�܂�h+�:T�{B;��Ӄ]0ӐZ�O^\�������^��uO��eN�V�v!n<n^�;��^Ә�:����>mX-w[�8��G]�(ͼ{m�v1�N��\�<��.��q��[���� M��:]Z�K�h�eT��Gv���IwW��<x��w]Ɖ���p$N5[�){��Z���.��x�[��F��+�@ڋj��[��<�;!6�f��HtїBKl�L�{\�'�b�Y#>�o=a��խcz��i.�k��Bѻa-.�X�0��4r�wY��U*o�V�c{� �m����*����gwgU�]~S�.�n$N̺��N+��˳���E�[ۮ�>Vq����
�2ˬ��:�,�:��׷^u��y�wm�*����]�+�|��}���+���n�yt�]�:�;����eY�+�â�:����VQ���Ȣ�{�w�O��n��mn�:�#��ڻ;�vuf>�u^]�y�d�vwY��{u�����j�;��:��˰�;�y�G|��(�m�]��#���t�f�HC۳���ge�U������Tukg���3�ˬ�+4�3.���:�o��Z���:�o���3mXu�N����:x��嗝�����gy6�l]yw��[�{����?�nm7	�om�\uց���t71�ݡ�ݻ�gx9u��������μ㫖v���vC38綠���E��b�l�ۗ�_XQ!'����(�6�J���W;�*�m�̏'kx��Y�C��8na�|��v"ܵ�׆iN+�wXr]v�ݳ�Pv뛤��9=�u�v���]�Ȭ��9��`�۴x춱'l=�z�p����c�I�{���軱����ձ�M�m9���݄+�*�K�:n�;C�	�`����}��,��jqu�tuN�c�p�;���W�+q/on���qaɝ�o;��9=�0K]n��i���u�l�A�:���a�����;�kn)]��sv,k����c;pt�Ks��n0�7l���a4�''n�Ͷ�ts�db�n��u�&�,:؜9n�;����]y|f�.xZy4�z�LMۣnŮ63�S�l�)��k*��}z穻�w9;��هgPX�z9�	�J��-V4؄:���AG	p���6�^ �[��Z�������s��w���ѳ�����؎~h�����!�+���̼�����[��v��qخ^Ns���t�k>�vT��t�\�7k�#��<�:Wa9=���vƸݸ��NM�a$�n��nuۥ$�o�A�������6�K�o,e�[�ȍѧVÏb��:���C	�On��qXu�N\���6��\�+�ƪ9�k\�=Crb]a���x,�%뭭��t�<t�'k1���3V�Z0e��n�VZOv��v�;��y.���
\r����D��`��P�M��n5�X�Z���q�9t���t��mp|����9�{�>�ľ��#�p��������v�q��Z�����7Y�I���!�P������v�6��K�»�� �=�����<&0�r��R��.{vy��H��IǑ���q>JN8�m��>u�>q����=oo7]�����������9�n��۶�d˞�.����/!�eL=ǰc9yAyW�v1��{//�o[�ד�L�����/<�&��&� �
vɜ����p���w�Sr���x_o9�]��{n��`�9A�7}��ݰ���8G�w;p㱓'd{�`6_�pm���U����ɗۃ8�L�\m��nNy6϶��D��X�F��6���<}r�jH1&LO��on�#�6	��sJ,���@�N������B�V$�TEI�G(`��|i�����
F�Ϙ�H%��"�H+�����!��̇�\��9�q���O��Q�%Fb���M�{b�X�r\¾��|H�Z��$��J?��7��E,P���Y�9��s�N<�v�v
=~���Q`��^;YX�^�͌^�"�GlU�����{��;�f�*��w�$�O��쳀s��9�j���9�t(�ͺ�9�y=��U�˝}@��:4:�	�\�p.1`�ɡ��ݽ�>(�Ӯ6Z�r^sg|��Ee�O�m�@P'�yX�B�'�c�D����m����+\�X�bL��Ér����ݳ����mM흚qi��f��f���jA������#.�X�w]䝛��r�)ջ"�η�5�'B�%�92���Y���)@�4�Y=�٘	:J�P�X��zvu�٩�;BƁʠ�������,a�
'�L�O_^��IS�d���fx��R,Б5"fhʎ�3��j�(q^WCZb�����ȿ.�[3[�x׍w�g����E�I�Y����A�̓�)�J��0efx�������
��֨/y��d-V��k�x	c&&J[���D���:�WX���X#t��Hڄ�B����s�X���m7��M�]9�L
��Z�����p{NEM�w=����<�u;�Qkx�ب�J�Y��I��5(
��`�h zpW��aݼ�c9��J��e���4.Ńm���0 ��րV�	��X��,ǌ�#�0�y��bĂ�9m�Z���v�lNX�)�V,��4�eum�yv�ɜQcy���F�g��ÁN56�;55�@$j���H%�'6�z��(�9T����9���y�9B�n:b�P�޴(��}@a=�CBms��sk�D���\EIky��vM�|H=�����wq���{�xH:=�j��[��,ز����z���Q�ۣk���lQ�ke��a������W��+�}.�C�^���jE��<�w3;�g�|�Z 
}z�3$=�4����� +KNl;z.JjA�$�UFaf�lQ<����#r�;	u{݀`$�%�`O����_�V�bf�X����q�hE	��@�Ui��U@�=�`�03���km�OG.�t�8K̈�T�H��&'0��W�OM^�X�V� �׳~$��oĜ|��1���{b+f"kgڱ;\�����ٗu��k)uGS4I�W���2��NhwcT�kǻ,�]�Q�;ŷ�����X��Y35�{�vmL�Ln)\H
)�}Hޛ����" �	�$���KpfCY�9Q�
�Ѡ�+�$�Q�s��>[�s7GB�+\{��Un=f�GS���ij�|KS��ݎ���:һ��mۜm_��'P"ѻnm>u���"b���P�͂A>,�ɲI��s<2��Pi�U/Ă8�ɰ�m�&D��3.�ضU0 �5<�����<�$�v���A�=4��kܑڎ�9�s�`��&��U�����s'�U_q8� B���RˠK�[x^�Vi8���TJ���H.������ �:tvܞ��f�>9�|�&����[,P�Bf<�;�X�M�=�6#ܱ3Q%B�6	� 5�0+�Ӯ�/��<�V��x�jlh��e]��Y��\ݹ�o+���6�,��6���+�	q�	�0R��܈O3D�1�w��q,M�TɊ2E��;"eU���mo7f��s�GkK��ɞ�݇�\0��N��&n�6YЛw\��[Ut��tox��N���Hm<ʹ�C��ly��>3Z^�5�A�YK��{0u�N����r�n#�m���s�wXMU���6҇��unK$�[×����.]{s�;1�:�OD�=盵�)���ۮ�yyۈ7�����n����2ۧ���v�sGj���n��`���sg��q�<k��'x�z���)�_=�V�y�o4���x�u�tQA��lR�/��Sӣa�7��}��-o2��M6��nm�V�.xz���q���	��0�|�͂.��mLf�5I��� �DϦ
��z�a#�'"� ���ي��Uj|�9�a ���ȾދQ��Pd�5����l*k�m��
[xH$l_9	(�'�&ŧw�ۈ�bA"����w^Y�T啲V\=w5�i��߳�)�+:2�l:�
���z9�� �{9�sWe�f�x�o=��>�����O�1��1���\��F�r���Ѧ�kdkb[����~���$�MH��&%�Ĺ�A��f���M�8�f��T��Ж��x�N��~�U�qS0k������
��w2էP��Ҷ������ce���שVE��}�����Nwe�K�u�̵����V���(Lʹu�Н:���p�������	
9�߉��b�@���z*鬽��O8�x�;�=$��gS�8Z�b��f�i?=�&�]��ă{��MF����=��@� ��4*&���ܔN����M4(�� 񏮐K�����2m�����M7���Y-!-s1>�f�W���I��r0Ǹ��I�G�ؠI��n���j�L[&�\;��f��Bq���1�q�7Z	�fYzޡ��mۚ�zXu��
�/���(2�-��������Oo��V�W�٘k$qуq��܆G�t|:�Ò:�B5	���{���4�����5�%d�g�I$y�d�ٽ��TP�oi�'<]k����iN=�=A߂�H��Rj���ķ �	jF@�]]��@f%��VK&s��K`�?EN�mu�ga���#���ɋoK9]O�{܉��+�HωY�Q�NgGu�l��M�9��|ߣ���P-o2����V3�:�>"'r����[��г��:��>����6�]�bD��$4*$;�Z0���%J͒�VO������ә�o~淪�zB8.+!a4ݭU������w���Ť���f��T85�R	߃�x{��%vF���������s��m���Z�0�r�Уl�>Pg.��	>�繉����J��jd�5��iׄ����UB� ���3���O��Q�;��nt墳�M�ݼ���T��MbO5��Am��$���W�$6���A=�oĩ���5�S&�\4P�Ȝ�:H=x��#���X'���U=F��K��ٓ�Q�G}�37z��u�(^�:j�MW��1#��v�ة���z58,K��"�',)��Y�LUP���ٱ���X09(@P��n�<ϴs^�M�l��ږ����7��x��ӛ���\��v���矾��z���Z����/W<3�kdNsv-����:������1�-#__���燇ڋ_�^f<A%nl�Y6	���#���_j��4-�@zx� aY�A9��<���_�ye�2,���~b��+�{ց$�zԋ�'X�v�UmZ���*rZ�V]3��m�����&��}9����Y�j��1���Nl�IG�X��s3f^U��Ͷ�r%[Iͮ����H�9�"�O�Q��� �;fn�3��2|<V��u��˻�ρ�v(��Q�ĳ<2�L�	���C�lh&�76H!j�x�.��EW`[��/�����:�C������NX�xt�b�08�Vi�!q@{�{!�c���:�2�Qx��к6����I+��	St�ӖJ����ֻ[����+=�L�!���!n.pvy�ez��zqLW!�v�:�^��\g���	��P�=�������9mp�!�v5������ۚ���x��ہ���.�zW[x- u��ų���y,v�g#�����r��I�O����1M�dX<��84�MnN����Ɉ��ם�Ү���,��7.�z�-<��Ob7<QzS�,��[n��r�c;ksv��b���V+j:N�7��0�#�8J5ɵnݜ���K]	ݾ�w��:6��}���g���ڿQ� ��vf�I��)k��BNl�	�ö�Q��W�	񊨈��8鏂��`1��k��� �˯��v`�f�2א���[U���B�-M��H��.��ڿfwًm<f�X�},I���v�ʶ2��(�b�Tz��L]��v��}�6���آI#3V�x�OE��]�;<�s'����ֱo0`�����m�=��t(@�֨=CQL+���T{��^+}4߹���KK���$�e����D��K�^�^��n��'7-���$�MU�(K�uy�d�b���VoQ��Kpa�$��`�^��׬1eZ�@���y�c�D4A��e&W��ϛL�V�w�U������E"6�]�u-^6�Ss��"���|���Z��6 4�R�p��Xi�h$��(��#����+��A#��M�qD��3uQ̓5�g��_�	�h�HwV�$�6�߉$�b;���y�ٻX��J��3Ă޹����n�B���k�L�5ބ߻Ts�	9�s0��v/�l�sY[�����%����5le���MH��Pl(�s~$�9<�jÖ/�we�E�Y�	/�oē�9��X��ӌiv��Q�L��W����[��5=���zպ���K�j�X���ߗ8�mu�]'И�����'M��> �Y^ո����X0��,%C��TA��3&�D�W�a0ULP֣5�΍W��H$8�sdQ�,�d2��f:���d�&��S�P���H��՗�>'����Pmp���G^�G(��l�����I-�7�w�]��{6_]j{,�f�B�21R�9EWXz�d64�lq��s0���c��7�zkle��Ճ4`�f�܇u3xS����6:*mlnd�]N032P�� ��V�C��|;�4��.)G���P� Y�U1�q�ȨX"��6/�����A��3�Y�UV8o-c�P�e����UE*��%�j�DRg�eOa.�n�eeF��uq���V���V�mL�2�u�eK��Z�h*����#A���%ǡ/tY�T'1�ڌ�ĕ.�B����e.*����M��۵�l��{'LvӰ7��W��Q��k��=ts2��ʥp5u�^7��>�_/�0��ohޞ�6�Af%�����Ϥ�r��7C�
�N����ӻnƏ����A���<έ!L'��/V}�B]�UϬu�p��M�Y �	�����j+�(��Ò�8�k8�w/v_3����E,��i�0��ۻ����8lf�`�!ӕ �{˗ˬщ:Ӊ̝O�]�}�)�E즹"���۬�k5&���r*�ع�[�֜�t�죁�H�;�L��,vY�ع�$����'e�}�Ú�f����q�i�JKɯ+���Sq��j$9ٳl͝JP�*���uJى�y�}/ݽu΅�+f�4��[�+ۑ�e���y-홣�wpM=m67���womn��ݛy
}@��梅�j]�V�o^S��(=�fa��ٜ�F���j��)�>���� '"fw|Ƴ�mˊ���܆(��)���{��Rٰ�Y�t�Yz��(������nҼ��myGGGe�XȬ���6�gu��ۼ������t�0�[�;���N�gy=͍����������;���+'ۻ��۾[j�my�eq�u��Sxą&a%�m!m�N��x�]�JW�ee�h��u��t]^_>�ya%�a���ڎ�2�+2�˼�μ�,�{q�q�]���=�9:��}om�e���U�n����y��T_>_N�����Vt[{�w��w˲�h�:����\{[�����N�D�6�N��=��;ʽyׇe������Y�=��ojχ|��ｯ����|��(��=��������g�v�{�[�e�����Y�{�GE�1�Ǽ�y�'[v��tw��=�=�@#�t���O�-9	sYV5����0��k���t �"��2u;2)b㆗H�H$�~��v��תe��p搶	��ٰRp�Ɓ��Rd�YLX�`�Mw�d���Y[�>�����`�t��(�v��#����2�I��>�U�4ԑF��T�e½c�:�[q�+���T����\���޸��*EGã6��$��v]=k�3��a��=2ٕvD���smU�
�uڣ��/-���O���7�w7��w�GM����$��6	'�v�T�!]^��ם�#�jʅ-vG���y4�O��7�`'������T%��>���,�e׈k���7�[��2���Ms�g[�N�q��GFﮈ$�����\,�:��F8��/�θ*
3�֘�	O�e���}۩fx�k�k1d'iV��w3�7\�+8o�+8�ǝ)Fq&2�{Ă�nآ<��_��b�TM��ŀa$�x�́Y'Z`��Ǎ,�(T]Ѻ]t ��0�4��`�\�����b�g�4�����[u2���lk�;&�4���{=ߝNH�q���w���k��$���6uI���j&fG���ٯ{x�뮪�uIedTz~�j�6��ʼ�zo9޸a�s]�5��S
aI)+�߲e �Kޱ�v�G�n��������Zi#�<��n�)k��I��6��|��fH)�@=�~ɝQ
�!M0)��w|ݮ��3���@�h@��
eD���ff�JH(P�{�����5��B]`ժ�X��40�՟��ѝw����n�ݕ�e �����ɱ�d�RA)�{��FR
A`i���y��zw���-p�҈UJ���s0۸�����͟7J�qN+���Jƾ�L��2�%2�)�y��d���1��6��A��m�Cl60�P��s�2�HS%�����s&�e�k��=Z~7���k^+���2���r�ww)N�n���>�nm]�L}�95�m/yޙ^d��T�yL�w�<*����ƩX�B3,��b�zŎWq�}v�`��
�<��������uzM�p�z���v=�,鳺���p���������/�v�q�k�68��8^�]xF�	���&��V��{j�v�3ӫ��,�RZ����Ӻ:�7����u�m۲N֌f�;�n�ޯr��q�`�v�m�!!�w��'p�+��N=+�q�cdlj�\a��v��U�Mܸލ���2Ϋ�p�pĥ�4DIU�@���X�T5վ�}R�0�����Aa�k]�4�R�@>��dΊ!UD)�4z��u	�@F�j���3M�����s���<ld�(�}ϲe	)�竽���[n�Cl7S��������$ǯ�_4½�o'm��S��
��y�@Д������}�$B��s��7�{�ǳ�0)�{nJwK���6b��BJ���&SH�JH/��s00��JB��Ú�S��yí{|�n0�0��%{��L���Rﯼ̚_��u�b�aj|fpi i|7��`E��ujO��$*��߲e �Q
h`SG=����)* S)>����l��{�ɿ{f�sV�E�)
B��}�(hIL(�t<S�TR�dϐ�X��������	 ����d�6Ɍob��o>�ǽ<�iH_c�h�����������(�TB�{]�3;�
~�}���}o����M���H�y��C{f��g�1th�@���*����7m�\\s�Pj���c�@o<�L���]v���0�	) ���w��6�q�0�O���v_�z����$�+<�e&�)��L�2����ɤ�t�V��Ļ�XфSo;�a��I�:��g�wX����I���|Y����%m7�w"��{�)ٮ�ة�����ЯaS�`����ŀ�y��!�
�n����Bwy�o��k�3�D*�D)�`S\�=�@��% S*'��s0�6�ʌ��wS��5����g�2�Xk}��b֮�Sn��L;S����i�P�$�
a���d�6�P))�|�׾}��}|�%0)�4���f�Q
���߹�m��5�ܔ�Z���!�k����Zk�Շ�7�<��S=�ᒒ�o�d�&�%$}���i��
H))+��e%��&�Y�V�5S%�y��2i0�R�s�[�.���ލ�lJa���06�B�����D+���p�n{��0)�k�Zh@���~�y�i�JH(R���2��Sc;7�ޯ�n�۱]��)�qR�n�hۣ���N̼�c�=�`��]���^/���~a��7�/�<��솣$�!L9��̛f�)��BRJ�{�H,w5ǭ^�Q���}��s�
A�C�߹�m�?����c��)u�X������2�@�Td�VNV6�}�^3�)�_w���TRS
������laL)�$�J���L���C)������+�݂>�������"�;�٘��U/�ƌ j	L/���`SI
���}�q�_!���C���t�SR��?�O�)�eN�NP�Q���_W j��̹��,����MX�;y��+��wfLG�S"����\�K{U����% S(����6͌��)
C��}�hIL+��o���T�d3��������ƳG#���񤜈RJ��{y��
Ґ*v��aQ)�M0(i���fLg˺�u~��u���UB���m���~ۂ�����1����N߷��M�R����C�ηU�����6��¹�{���laL)� }_w�0�B�C)��S���̚L��_^g7W�������=�r�p���'�"l���]��
�A��s-sظl�r��[!/1{��Ж���'��B�o|���<�%��Ih]�-��ɍQ4�ܢZ�ah[s�c��6�� Aˮ�������P@��ֻ��3�����hZ%�|��ibMcJ?��p�s::K�6ҍJB�f��!�v�R]�ZN������t�������;~q%�I),KIiu|��I��ZKe�i-�6���3 h��LIr����F�e����k�.����O��Ae�ϐ��b���d�hCH[,e�l��B���̛f��%�hX�����9��}�}�9ڭ��!��h[mIr�o��L$�j��Spe��)���fM����|g���5��[��H���_-�G���IQ��}�(J�A��F�ZD�k�Lh�i�%�m�-ns��5��؅�i)
e�?���'X��-���dIT�V�k���b���"V�l��i��Ah̢R�S�����D��ON�}t�W:�Xn���vz(e�e�hZZ3^�icXҏ�����j"�+!���m�-���d6Ghe%���)��绝���Kq���?{[�I��%���U����L�I)����X��_��6��D�*�%�w*�=��$�)�B#Y�����EvB�48�dF�x�DcOh��i���[Q����ں�W<(����>���*�cc��������O!�-�2ж\e�o{s0�CbZ���l,���q%!L>/?q��s�m��t7��&h����ZKl��ܝ�[iV��W��l�9l~rb�L&Ķ��<g�-��KC�'���K�K��'Q�wy1��i�%�m�B�r��a�0�Bд�B�bs�s��IHS82д�層�:��y��ҭ/&���.w�㘀��]�h[������Cq�IwAi)
a��s�6�����$��5����}ϻ�]wI��ZKe��[-�ݿs0���Zeл�}�s��IM!��^����*��!����J1�k�0���c���qU��g �B�q������KB�R��}��hm�жB�]�߾�L$淟M#񝅤�L���-����C	)6s�x]|SX�%�/)&�il=�}��x��ci-�%�_}ܘ�H_4�����xc0�-o�c��6�`��ihZ�N��w<C��-e�д.%�}�ra	�-�=�;�|Լr�X�׋�Ϯ�]�=�/��l�[���D�ٛ�֞5{VWj9�5lN����P�<��٨�S��Ţ1B�����4��8e]r����5wj�A�X3�)=r��;j�vV�n4.�*����m�"rn+V�ۭ�;�p�Ӷ��n.�m�;�nkjvk�؞�����;p�ڷ���{;g�@$&�㎨x8��ݧ����F�j�CG�ָ�$��q;�=q�1�/��["����<:0{�(O��=e��n�t�q 2�C�����ȫM������j5B���d�9{U�E�CN���3j瓱�]��yvY8�c_+��{�N!Ĝ�	߃;�OV�'c���4���6���1̆ݡ��.��]�[w��v��Km�����Z\�ﻣ	2�$�7����wo��}��ϛ~����hl�Ф��YP����<ah[f��%<���0����6��дo��&@���X�Bٺ�w��g����W=:��X�O��0��Z���l,�}��q%!L8��ˡ���0�Z����-%�ÌW���x��ͷ���É�tw��ﯷ�W.c��w�ގ������<g�Ke��в薍}���L�Z�Z��ж�^�5�oz��jϫZ�!i���i)
e��{���8�B�l�-Ѿ��0��H[9׳h�)$�ٛiG��q������b����P�K�IwAl5���;x�$��-%�������wFe4���q���m�{��C�n�w�p��W�u��'�Vh]�>�\�x�-l�d< ��dw_!��m4�Nk����(RJB�R�c����>���W}�Eֺ�Đ �A�	�}����ж6�����}̘I�PZJm��Ч��;�i6	�����[�=��������B��̐���j�ԧ-�.�$�*����i�TcMYlr��[�P�d�_ʒi<���k�g���%�I)
IH��s&5D�����Z��w=�6���$�$d�}��t�O�$>�����)��-%#_{�0��H[_���w��	������m8Ҏ�ךCN�(�O��G�ec���k�4^=79.�NU�f����7�vո#n��S�[��#�w�e���B9@fp�Y&�mR��V"h�g��F�ч���u�v�3�-
IIbZKK*���a&SQ-%���[,m�;��CsKB��h^����k��Cx泟!䔅<ϸ�Q��5x,��P�������N!�-�h[,e�o��ɰf�����ih[��n���\ν��z�Xu�-���i,�﷓	5�IHRJm����s�i)6c�9|�`�cw5���=di|����O�<9fR���)�IhYtKF��d�L�Z�Z��з|�;�iM�Z�Z} ���v���j�y��;�߾� |�2д��s�Ʉ5H[>�ml�L%��fm��n4��}���Ҭ�.��Yt�>����3�-z��f���w��I��-%�Y��a&SQ-%��i-�6��c���ي%�WD�.����v���$	7�컺����o9�⁝<v�E�\s�tN���v�27:�3��m���o��c�c#�I��^g�BѼ��0�CH[,��-%!N��;�iCbZ���l/?{��q�B�';�ܪ�?o�ZJF��d�O�-%6���=����HZJO�ce��5�Ŧ-�d��O�[�{�<g�>�$zH��5�75�qǸ���>�i�%�i)
o��{�mIHRJB�g��3�6ϙhZJB��tЃ������� ��b�� I��{��bۡŎ�4�q�-ǹ�d6;C	)
IwAl5�{���q%��IiqQ��_�/x&��-��q��({�ӁuB�kns���Gݰ���@�����{Y���%~��v��d>����馎��ا����7%s�Q�"H��[i-�߾�;�m�hU�-a�{�������m���fT���E�z�д��}���oW_g���;��Rf�h[,e�n��o&�m!q-BĴ-��w�w\C�86���д�t7�{&d�uϱY�s�p2��e���[��^k嶷�U��R�^M��e��n�6�)����<Ci)�Ih]�-�^ɍB��,�����=���Ihq�����>�6���)6��l�5����gZ�hZ%�}ײakQ���-�g<I�Fi��欕�8�\�77N�u������N�w'U��#��V���ɛX���&�䨳�iF�C��{��0���$��[{�w;Ci)
IIĴ��W�{Fe4%��W�ɼo��wy�q�Il�����6��Q-
��h]�5�}��<Z�>�ҩ��n��j��`��y�a4!�-%!L�/������hGz���>���B���-���q�-���-%#]ײa&�PZJle����5�Kl�B�N}}�=S�~C �#�D������X��xƅ&�il7�o���-�6�л�Z5��ɍJ&��(���0�-�o���1�g���c�C�a8��ihZ�]���q���-��Bд�o��L!�4��������N�uZX��Hs������v_�>R$�)&������v��S��Iiq-%��~��0�)�-%���X��?~���AU����oR�H[E��������Z�u�r��次�,=K�;ckv7�"��toq��vf%%����eY��qp��Y���߼߃�@�=+�P���{<C�Z���fT�/]�B�R5�YɄ����\e�o�IO��v4�H@��ߜ����a��Z���{�q0�h[mIH���&jj��Sc-%��}�㹆�i���+;ˣ5����}�*]4��H��m�94�vU�vx�V�d�z�t�5D���q;�^��m����I�m�����/s��x�G�-�Ih]�-�^ɍM!vQ-n0�-�{�-6!hZr�����!�b'���<C�)
ghZ���^Ʉ4&��t��U�U�qy��`��]�9����.��|_7��c;���go�Ė�e������ʿ��I��ZKe���)����Cf(��$�+��u�k>�5���v�_��v�φ���=(��ؗ�.��aHi%#X�a:�����2�-w�c�6͡�--B�ж��{�`���]�a�ж6�������0�ST���-%��}�c���i���|c���8��8[�2)4��l��h���\h���!(#�}�H��&`KF���1�&��(����)�s��P��Bд�-e��~�3�8�}���>q�^|�<�Yᖅ�ih�{�CPM!l,�9�f-�\X�1�!�mq��̆ݡ��]��tÛ����������cU���uy�Ғa--%�\�y0�)�-%��IhS����!��%�W(���P�~�3�8����\��(Y��W�6:u�O��n�	�N�r�f�(��Mђ[R�8�m�f�9��К|޻Y���w{P�],њ�ٜ܄�!#F�I�#g�̌R��6ã�-��9��W��9k�`u��IC;3n���{f�&� e�C.�R6I԰1\b;�em�l:/9K����X��f�^�q��5�*�*��� j���j���wf�oM�9��@}9eF�|�Z��F��8�{�g�z��Iw0��#.L��U��fT�C5k��Ҳ��播���x���6B)J0��.��&I#6�w�NGWW��ZoD�d�kɓN;U�wڝ�u����{��|�Ẍ́��kr:��X(]�&�j��-f��I��utӣY�u��6�d�l^V�UK3Y�sr�8���]u�aC��mX��%�Bj���5V����ް�]�G�ۗ�(ԛ�2�X�c�����df��O���v��bjm�80��:QrY�A����D�|�g��ګ�S�q�EV������	�����Z�%�� �5v���7�66�N���{Pv���/$�n�Ѧ�r�&�m
�GIK �v�1�.��	���4�qFu��W�غ ��7vnܱυ�4�m΁���\Q�n��U�L�����{\ԙ�N`Kb�Äz�fE���K�O)�ˀ?;�^��є�g	I)��7r^��Ö0Һc��F���*�Et�כ���4-,6�M{�%ݮۧ�\���v�W�/���ꭣtt�}���n�H��Ɋ�bt١,�� ��F;� Þ��@.�n�U��
��lM��j�H�/,����Qz\q�|��w��^y�Z]Gg���w�L��w��W�yck�>^_�ϙ���l�:��﷝��Wy��\W��m���gNӏ����$i�W��8��ʏ|��Z����{�e�u����+#:��o���^fݹ����{s>@��Oy;�^v�ٝ�vW�YE|���>ގ����_�<�"����;ˎ��vwE{[��e�E��ǖ�������E���{Q�u����Ȭ��ʗ�0n�[0�Pa��Jd-�Ɇ�n�e�yէAgaGgv^^�ֹ��vfw̯;[HR"[H��a�Z#L��U��6�glϩ{%�O�{1��ݏ]F�-�rz�y]���n�=�Zۭv��Y;��PT݃p��M�6��T�n7OI� �ۄ]wnat�=���wN�g��8���^��A�ڑ|�7Gm۪u�q۳�K�a����Jnh�	+^
��Y��KLێ�C��^l�'n99{��ؚp�7E�=7�x�݈���;v�E��n]=eӷ4��	����&ήK6=T�wY���k K� �v0���=���n��Dr���Eٹ�z��N)L�M�q|/I�]1�v��&�6��+y�1�	�㗵�kRv㱸���[9r�Qƒ��ܽQ4�*��y�rl��w]<Y��-��!۳I��jl'>L؀:A����ޒ�5̩�'d�y8�gn��d�=ۛ�m>�. �s)���[�$�]�:��8�O:NMnݞ.s�ݲt�6�vb�{Ilm��L�Y�9��G;<�ѝ�U��ˌ@-�t��:���v}wҶ��3����q��v�؊���fް=g��+��D,��.fu���r�����4�#��ǁ1��m��<m�탅�[���:��<���ɇ�:�a��L�>��6����w6;�;mi}s�����>���v���ױq.�<���k��N���[ڞrvC��2��g	��5n��;q�-÷y�H�v+{a�n�s�9^1��-��=d�ut�qa��6˽�,��nw��ў=��n�m��x���v=n����u�����E<��]�����уa���9ʡ��3�n�#���o7WHz�q+�l^�G\��:�8�B�w]���$��<���r���N�=�{=i�7�o[w\sl]OQ�6�& z�1����^����v�#��7�8v�oC��n���I�S�lzy93�!�k�O&;x�4u�v9M�p莵ֲF�nL�U�	�]��=����x�>6<����ms��v�v4�ۈ05���Q۝Z�k�'�4���{�����&sX��5�s�-˗�(�ל��M��g`L��X�;�����E�� s��.�A��m���k�w۶�u���u�g�����ˮ|�8{���۱S!��\6�s�ż=g=τK�ꦕ�z雭�m�O���c�͎�G�	�h�z6#'G^]ɬ�n��3��c\m��鹫r�S�Ge�IݏeԦන�I���e��^�bM�d�կ��5�jɰk�x�bE��M��{�ຍ�Mڦ�ǹ�}*yL[�,��C�-%#[�ra?�ie��-%!O��{&�m!bZ����=����h[���Ӕ/d#�0�+G� 	#���Im����;�m6&Zg���X�1X�a�c^M$�ؖ�~ﻞ3�Ė��4i����g#I�q3��1�@�(����ж��3�ChZJB�Rͧ��s<C�)
gZ�5�f��&����e+@DaO���rI��[��������>�|;C	,�IwAl=�}�����-%�I))JKo&Ֆ�U�
#�B�G��L��e���1��hl�Ы�Zr��s��\|(Ҏ_{~+E�|���b��Ʉ�/W�y�kf��������9�1����B�д,KB�_=�s\C�8���д�.���d�OY���+5��������9���a�)%&��<.��ԼZb��
M�Ķ�9��x�Ф���ѯ��Lh {��w�l�r�����$	3�{5�I�B�д-���=��3�-e�Z�����-D��}u~����g��(����I~��ٍnuq��c 9��a:�n����0���_}��H�p���6�����Cq�Ir�-%�Al;�}���8�Ф������״ZL�I)�ݹ����u��IL�ۏ}�fCsKB�(���C�������������K.�!i�G�oY-4!�-%!L�1�޹^�V�ԩO�͡P��abX�q:�ٸ�7ZT��+��Ip+bl�7R�������h��ż<��嬳Cu�_�u���~�C�3�{'�0���i)
a~��q�-���i)޿d��B�S�e���1\���i�yַ���2�_-�֫_F��97e�I*��M-$�ؖüﻞ3�[-����D�~�{%�i�D�-%!O�u[6��3]޹�i)
ND-a�s��hm�h[-���q-�^�hi4��(��Y`���ݹ��-�ҏ��z���1y�ˊ�t@�=��G�`	0�w��oq%�I),KIiu�5��I�Ж��q���m���s��^sZ���{��1�@���2#��ﾴ@E|4��}��|+E�|����iZ9�=��e
f�Z�e�n��w&�m!��5{��{u�C�)
a���u�8�����$�]q�d������ZKle��q��i�0�Ѭ`�>�C�˫z����|^��l�����<BӢ�=��9�"'r+���:����}��Wv���^<)>O	l7����9$�X�KBˢZ?^��z
&��(���-o��{�mM�Z�Ǹk{�}��g\�Za���3�6�2д��!bZ>ƽ���iag�ޝ�1m���Ía��mq�c����K�I{ƫ�y�U^va�g����Km����ZKG���ZL��ZKB�S,}�㹆�ي%�I)
�g}��ս����;C�)
{��Y���Yw�mIH�����CH[.2жX�B�w�w&�m!ihZж5�_}��D�9z��.��F�ߖgDI�V&;f�+�'���M�M �bt^%Q�
ʊ��P��E��*������w����		�o����~B�[hZK.��5�%�ѪIM����e���ߖ��km}���&첲J�T�-��#H��?���Bv.W�_щ4G��񔖅�����KI�+TKB�R�>���m�д-%!L=�{��b�k>(�����Je S+��Ô�w�:.��,�[Θa�}��H��D��xt �i���鄝L�i-.��u��e
IL��KB�}��Cf薅YD�-��绝�m�����~�/����9�?>�e$�6�Ld,0⮛v1����Y���)p`�j�tv}��.���(�V"�_�!��~M(���ZhCH[-����Z����m�bZ��h[��w\C�86@�ࢩ�ņ���_eAﬁyz`����kT��i-�[�{���i����}�筒5cT�k������۝x��m��6}�5�_�Ʉs|�Kܢi��h[cB����a�6�Bд��2��绞!�q����Z���QZ�s��G��Ç�>�0���qc1�a��6���7�۴6���\.��s��s��8��i-,KIi��ɧ�}i���	2��[,���\m�>�!�6�Zeл�{��s�8�ah[�n�P���rk�(��Q�{y�����zo����P��e�l�Z�Z�!�4��Z���l/����q�ж���`L<�ő��n�����U6.v;��"���v(�-��U��R1e�{�n#�tu{�Z�0��eL�+4�J�a��R�%� D��l��������"S�e���[���ن��JO���X�^����k&�Zr%�߻���8�%��Ih]�-*���Ԣi�}���Z{�>�{�u�ah[x���Che6!hZJB�i߹�s�8��-�2д,D�0��@�F$�V���E8[��ݷfq�n��c���u���AB���h����5��5[t�;��|^�pR��N��iF�)�k�v��Yt���{������$��i---%�Wu�I��KIl�>��s�S��2�m�k��6��Q-
�%�wP��}��<�-l�������P���im���P�?ii�M,B�l�-�;k���=O96���fC(z%�i)
aw��\C�8���B�]�u��&Re
IN�ZKn����f����"��#~��3�T����ƅ&�il=�s����)%!ˢZU}��gEH]�ж�B��8��8��x�w�v!��Bд��0�}��hm%!L��Bд�o��L$����<�qm��1��0������ѝ:��<�$��ZJB�{z�����������ѯ��L$�i-%��i-����{�m�����HV�h]�{_s<C�Z���Y(^G�p�z�д��}���L�I)
g#-}]��63his��]wy��e������g�渇pmaq�-%��~Ʉ�PZJB�S'�~���i�F�!����FV�nX���zgOX4Vt�z���F����*�|']�Û;�M}{�6���q��Jm�lL��F�ǃ�̾���#����]�-�]����E,vh۴��g���8��lm�o���+l���avù�����Mv�Nl��r$���#�����y���qO�-x�Aml�s��[���웛��vz7�s6�c���Q6���n4�,���K]���2�0q[DvQP�8�8�u�Yɓ�l�Cu�ٞ�;	��\�^��n�C�y.G%�y����C��7���=#�Qۮ�ٱ�9냵�ŋ�٫EƳ}}����2�j�~>Ii�Ka�w���Ė�Ih]�-�~ɍM!w(����)�w��4�Sb����=�c8��2�CL1�s��g̴-%!H\KF��d�V4��E�,��Unm��i�������H�NU�����gO�Y����goq%�2�ZX�������0�)����m��X���{�m��� D���+9�<����>߻oH~O�Q��~2#�E�|������Ʉ�B�l�-%!N���0�CihZ%�l1g4r���k׏���Rà����߲a&�PZJm��Ч���0�m4���������0�,�ƅ&Ц���v����;G��'m��,�%�X�a&P�KB�ah[}�{����n!hZZ����{���3���ߛ7�ru$�)��x��a	�-��{0�W��gi%!M׷�����.��]�|>7z@�=����;�r5Ow�i�ZKK�ξф�B�S4�Ke����s��tKB��ZeC�{�����F����/�e������']�tg�x�vGpn/6�M� e��pi4����5u#8\c�q�B�8/an�!i�-���	�!i)
IHR��w0�IHRж�{���JB�w����y���N��~Ʉ�B�R����?s_,k�m��Q/iӛ�U ���ŶKMĶ���x�[.6�Ьk\�wf�<~�!�w:)��U��f�C�ވ���<i����e�f�7h��3�K׌�8���7�O��v�=�q��s��u����#Z��c��iIHSpah[r����CI�B�R�O~�{�!Ĕ�3�-B�����wߟ��g��H���L!����t���,��Ÿ��c[B�lB׻�����JB�]�[w��;x�$��i---%�k���<s����L�bZKe���m�=��CstKB�Q-�����\iq�?�iG;��� ��W>C�дo=�L'~>��cW^�W�q�h[.2е�f�����ih[9�w��a��-������e��(�G7���x�Y�w\#�_���ی����0�n&�ZY�{�u�[���*�I��Ka�o�g��$�[i,�3�A�αY������-�v��IHS���桴4�Bд�B�s����gZˌ�-KF��X�x� I��?tuJƖ\�扑�B׵u{vW�G.���n�qΖ9�=rm�Gv"QĪ����8�wt�	�{u��hZ��Cq�Ie�ZK�a�s��oĖ�$��-%�ʾ��0�)������6*q�>#�}fIw�߆�4lI&�h]�9�{��x0�-�>㒣�X/an��i�-�zɄ����@����0�W9��&�+��!�--IHS����q�ж6����o��L$֨-%62�[�ރ���Y=��Èdi�'�Y��*(�b��Z6��`�Û���ǉ-�IhYtKF�ײcEH]h['�H~���r��\Ο�Mf�eb��FnN���T�{�0���-^з	�ݘ��Z�X.;.-�=����g�񚌘�L���n���<ƴ_�	$V����O!hZ\BжZk��w<C���B�pe�hX���_�a	�-���ӽ2�!%V7-ʹ��mƔo���%��׿o�}Ϊ�k�B�R��Al5�}���8��i-
IIu}��0�)����m%���W���ho��k�s�e>&��%�vT>���<Z�?U5���Ma��!�؅�z�a&P�j��'���'c���@ě�ϲ��Ǻ��aĴ-�����\C�8���B�\��_d�MMQur��y�{�'�<k��gV�VsO#vU��US��Î�'��myM,���t��;�]8�:i������{]������$
��&�$��x��z��j�����g��V��$$�I4s]���~��H::��kG����vx�v��{���BI �˯L:��8F���t)A�����N�WeA�r��&#^����y��Ś ]L�׽n�����E�o_ �o3A��N�U]VTbF��s~7������m�@���[z@/���	�$���#��f�y']yW�����xl�~1.SN#&��n�e%��=a�Y;�v�4ƷcT����Ǐu�jޚ���Ass�*����=� ��� �f�5��s�{ӂ�I-�Kpo��$���ؗ���k��h�$� ݉�	'�y�d�����8U��5�8�gЇ�'m!�'�Z:�P��烞����e�Uk�"4�$��o��k�����W�!�J��=�x�h@�g���z�`I�´�#�H�D�>��&�k�����*�=��w��A��C�~ġT�q��ۈ�I�=2@5�~�4D����r��F�S�q�oD�31�T+fb󹫈�~�s6��Y܍�W4F��痷�wēᾍ��$>�������Tn4U*+ra�5�MfŻ�Y�0�'�|<��I�O���$$�$����jht ��1�I6�h���j/֫ck��7����'{�8x�o��(�㍼d�$�l���"��Z���op�?zz�Iu�i���e�ΓN��ԗ���/VFm����v~��JPg��է�pR�K��+1�BYinUB췻$������x ]X���]G=%h��g��1��ࣹ����K^����]�m�ױ���v��/WF^6sָ<]����'�d��q�n\�.#��Y�㚷�[�w���u��=�F]���ni���M�;o�䏕V�Hm�s�<���k�[�8�q�n����9��K�y8�� ���!ˌ�c��U��q������)��A���^8��N0���Ӷ�7���б`�NΑ���;��r������!%�<��8XI,�Kz7׼���;�f�	bL�=.�/����=�o���������$���!�,��E^`�禴�Į����6rc��f��@/s����G3�_hb������ц�{�Nڭ��.�V)�>Rt�`���ց �o��%�<F����������{��zi-�߹�h�v1[3>���|y��R	�o���� ��e� y�ȹ}�d��8a���}��s"�*���4b��H�I5��m�S�B�:��b�MfM�% ��ֆ k��5�)�|���߽}?}��Q*(�m���z��s�ky�9�k�n�➶Z���6G���c������"���ĢI49��'�@�Mԙ>�;pxy�����m�ID�M>}i5�Y�7vr�7��&�ӒtJՕ�SqȎy'V�gU���-�C=ժ�FLU.�N��B���C���*X�f¡2����MC�qHZ'H�!Yq�/�_�K��\�5��8� ؙ��� ��s��� �i�����"�۬���o�Mv���W�=sӚmg;�k @�~ޞ�켞�%h�Cϭ"	$׷u�|t���!+PA���y��_fr��q���$������D�'kN�$����#\���毮���P3ݚ�-���IQc�٘�L�g�0� �=�f;���<�2ؐ3�������b���{����w�[� ���0�;J���q;mgv֬�L��9��etTvAAȥ�FY� ��V�7'O!�M}�׽�gق@}���2Q˧ �u�
�Ɗ�j�[繭<�s#ڕʫ����{;���:��י��ȒMhn��$�I���d���~~[> �yY闁V����	f��;������oa�"+φ�(W:9�M
OE^eҧ�c5�{Y���a�ɤ�k�˦�5�"�;��e޼�2S�-�pܻ.N�]�k��vzZ��y��w��s{��@�fC]m�I�[޷�կ�`�.;�����,WT�o���,�*���U�u��]�y���r�O�w�^k�;:
z]G�nH����3�����ᚒz�S�(oo�-����������on�GzՆ�������;ru��ީ��5mw�>�r���ٙ�ݘ�O�m���iVd�L��3+��3ۇpw�do!�+a�b7]w�^k��Q�4R�"m�M�Ekt�6���L6J�A�˗;*Eޤh(�9���R�S��V�{R�FF���^=�-NcH5�[�r$mR4�-�0�ٖ��e�Wuf�� d]�����F:j:l}���Ո����$�e!,�+; �p�h��C�a̱�A�6�r��On�����h8���S��v|��E8H�*�h���X]�j���LȔ�\�\���i���(�U�l���z�W@���C��A��\7oo]�)>�K#���
mu,�k�GPX�x�92>] �mf8�M�/��>�Nt�j�'\�4�SܫRN�9*�ZK�2����Ά��iE�mJOVh��]\ҳ���d6��s�35��f�4T2�l�Mѫ=��5+�sn�9���*�Dk����y���(��3�l���]�+*_V�CY++(��q{u�K�ۥ��SNd&5���̡{ef���{[���-�jHa�V3#sQ�
�b�\��� T�&��M!ˢ�a�)��Z[I1U�<�+�(�o����{iG|�;y�}���N���{�e�{fp��7�l���Y�w��z]��m�{޼�*{Yvݺ��Y�/;���^���e����̹�V'e�v6�׶���8�3�����|㼟l+�mY����:�"�:���$����W����������[m�����Dq�\t6��*�->�{�yyQv]�{���]��֭��;K0�l|�'�iM�;<��I�$uŗbug�����∶՞vw�Sk���^�]�L��u�y��#��׷^w�U����m�V膶y�<��u}��xٵYݝ��j/���[c�+�7v����Ⱥ����;����̝�w�g�I�ƛI�so0�<�^VW�Y��,[T͛h�,�.�
�֔g$e��K�Xt]�����͢��y{۾�咥0�\ b�a��	 C����⪈ ���3|�{���ן>���A�����n
Ǿ�i� ]�i���-��A1����S�OlOO#z���H��r��{(ټ,t���N�I����#ga���2��I����N��nQ �^�T��/	7��zN�ӥ6����l�3�i�:Y�q�����8(m����qYio9�tE��Ud"�s��m�D�w_k��$�I�^�TO�������ƶn�� �϶HI�<������Ɇ!�M-{y��|�l�h�5��(�I4uz�"	4y�L�sE\]����Oۮd{�%Q�ma�徏����T��F���6Kc.��ּH��D����[��$�;�5�[�<�ct�,!+�s��M��x�F��kV*�I:�s��$�h� ����i������Z�;u�h���X�ȃ���%��H�T����&�i��^9o);`zf��X��n��)��B\ۦ�.�6�^��xx{�_�������������B(*�zϐ��o�MQ5���u���*7�I���@ �G5�[�Y�s1a;�����>�x=vu7)��p�x*���U��Åk�'�p'fۻz�9
'+���˪?TBVۃ��޻�� hvu�D�$I�h=I��nWY>Z�R�쒉4H��֑�۬ˡwyYvn�-?����d���޲�}{g�3��� ��s3 ֽ��o�߳e��o��ȁq�l,dnM#٩�D�h���t�$�NM�ڴ`syN�t�;٤�6�߹�i��sP�I*��Rgǳ����vOf�{�'��*D�H��&I�O���I�~�z�2��F��_f�X��Y!+Ѱ\�{��Q$��<�4f�'�<�D�b���F�}��h��9�%%�D�Emz���v�D�Y�����þ��
�D���
��{�Pl<6is�n���ū䦍$�
+�ê���ײ�1>��|�IN�z패��Z�c��cʘz�Gb"���=;OO;p�*��r�n�ٔ̍j�;Z����ݸ��[�r�v:8��j���"�hiX3�Y�ݩ0WN盲�p������u���6�+�8����䴦�5�����Wc��C{^8�a�q����GJl�^�d|tOce��s�z� �,�8���(�����˸npq 3�$�r�Ve���z�����I���p����*'m�?��B�칿�5�HEQ#�_���ihs�ϳ$���zHK�����U-�h�/ D�w��X�]N����qE��\�7����~T=C�h՝��D�h��{��H ��~���trF���8��~�,A%V��F�����>�7��BI4L���z
M�z&p Q������f�����T��:[ �ɆS�����Gu�V����[uM��?�9���I5w�>���)�z�{�Mv-x��f9�K*��Y�s����	 MY�H�Z\�/m���d�3�ӢOę�=$$Tj�|U#v0���w��|u�F�m��v�;y�����힎9�2�#�%�g����ꝱ�y���8� �r9^�g��� �3~���@|rs�m�m���L�vma^�S_4���礄���Vu�(*�z�noƖ����v��єZ�9v���w|����y',~����@�z��-���5�LNn,�z��u�_^;Z0`1\�n��	���χ���|��Z���w7��bB���h`+�<���gn�`zk��Ϊ�M5Y��w����(w����+�g^����Ȓ{��5��H$ѫ��U�^�~�J�*��홈���/�������[m�w��` lNM�����]�6V;~��UD��9$�D��<�S�����k@����x���@.�;�����5��/M��y[M\��z��3|`�`�f#'o9���@�x�'[s���M�xm��v��c�slk7��|��R(쥐�����x��@��	I$�M�2o̣�{����s�
Nt��n�oQ��+�J�ls�v�:p!�+��O5t�c؏Do�qQ$�F���A%i������kY���>W�w�ATH����k@�&���6I4K���ǔ>?d��^����[�;�f7K,�����-��^/�bec���y�g��Gk��e�6�,�����=9)������w�|_P��+z�~�s4�/L�gEU�F��t�Q�=���f��9���Q5�q_"h��z��]��%pi�:�t�|k@��w��%V��l��(� ���T8���Az�4+[�M	x�"@5�l�I�����m�����YEO�q��&����(6K��{h�؎G�lq\�aCe������lY�y�W�R &�_:lD����IF	�݆�f�fp�3N/�A��A�=TnRȣ��$�=�߷��qj�j�����w�h	���� ��������|,��フ	�R'�iX��j��a����f߷����sfi�נ�+����	���`πK��{{��Ϻ��0�
�G^5�^"�F�y����4M?H�Ğ��M��Vs��=JA�{:�L���pҧev]��Ĵ�u��0�u�e�Sz�
{=��s�5]ӗN�V%���m��\m+W����<I�@���Ł�g��
�J�q��	�7��a�6������$�k}�r��D���Q!��繽� ����Æ�7s�E�Fnq����qdo"�}n���c���?UC�+�۔�Y�3�W�޴��*�DZs�-��%� ���y��| �x�G�c�4߯�l�uQ��n��?Ool��>O(V�(Z��	�>�tV��������Ÿ�l =��ܢM~5��)�r��j��z�2�$j�d�G������j����8s�f5�{����K�D�f�ITI�I���T��c�ڱAڜR�0���w��. 7�wy������H����ְ/��3O����n���@%=���T�$Tr:��xց�.�Řqzk;c�t6���|H�_qT�4I�׷c@ߛ�ꕘ#A���>���K�xo���:IU�<o���fP�9���h]!�iV��o�Zn������R�G�����}����<yn�Wl�����+&:q��*���υL�n���<۵�l�jxmN b�1��f����c��/p����O�JG����ܰ�g�cf1<�v6#�:I���K��35ő�n�.�9:N�e��1=�v����IӉ��M.P����s����Nz�!�r���Q�:��/6"���@�x���2����H:y�&��a�^N\۵��e���k���b�f�V�F#�P6�6��㦑�����_��*��NsY���@��u��9d��FGg��$�h�Y��W�v�B�Ic�VW�
wy�,��^�W����Woϻ����b;��t ]���������|�w��na�Ua2b�t����{��f��\v����z�&�s�DOƻ�n����j�d�F�=��S3�~��S���	'ự�D������kk�k����/^��w=��T�F���d�>�M�MQ3މ��������c$�TkgF��{� 
�J���Q�1�S�+gԍB�ɫd��˭����Z�d�WV��r��}~{����/j8W�!{/�m�w�Ř| {�޵�9��!Ii��kx/��jwF�d��W:(�*�,s��sZ�W��8�iE�t�h����!�&q;���m��*�+�'je�Ԕa$���얯0McQ�
f��+ap޳c.%�����<<�៊� ����b@���f�]�=����<�mw��4��o^�\�Ui��|�y�f6߹��0	5���(��Q&�{v4$�ލ�}�tks���0��S�|����4��$�q�� {z$�?Me�A�u垏��s9�fܯN�!��$��^�i��
��_�\�߻�9���������g� j��YV���ӏ y��m��,���,�j�Ml���#��ֽ6ۺ���p�$���}R�H;������w>���� ��.�b飙罡Mwy�`π����1 ��pk+j��,�lԿB�$��=�7�#����  =��3 
�p���	Bsw�f/M^i�v#r�8�E�}�֟���)I���2���t�����o�^*�����r��D͛���b#���f�������[��TC�0�4ᅗ�FTKI�� xzƯ���{��1�����\�(W$�[%e�l��F�x���ڽ��A�I=���/}.� ��sx��n��w���y�k��f�e\���Q�x��^V�D�I��Bj^���ͥ ~]��$�F��ZD$�k��Г���{W޿T��T�$�b�D:s��s#k�Л��֔-��`|d�_�����M;'5I&z�k� 	�]��  ~�9��2^b�Y�>Is30=��KA۫�BX�ce�6���k�*���vk\'��Ł� 3��[���sY�>
{�_�׵u����'kL���L��j��&��N�M�����7�f�����u��6!�Mhb�{��bX{��#r�Q1Ŭ����yOj�=�Z| ��KA� ��sZ� ���É�!b�d�N.T���&t��D^���;�߱���2��,��X��=���l]�׏p�ʌd�S���g\4:�{�"WN��1������1ʇ���</�"!'vih7���e$���]�3�S���٪$�� /}���ŝ���8��$��]ݭ� �'��F����ZWw�:�����ӕ:�j�����#���b���N5��a�ETN
�A����=�ح�ڥ���o��.�| /s�ֱ ���,����ѭ��R �H�{u:d�קv��#RZ�?k��, ÙKβ���l��oN�&� �}��$�k�ѷD�%:�i�s{:P�f"bX:��
��[��w��o~����w��Gs���9�H�Rn�L��>�D�2�E��P���j�Ёs�!vv�q�� W7��0����g�| �=�鳰��GA�I�'����rύЫ�9Q1ŬG�}��@��5���o�����k�Q��	��CzF�&�5Sލ���H�|���#9XQ�S٩�/�i�LS����w��N}Y�>髐]��WGU�-����Ls�G�v���f�Sw1�^V��	
��ɹ�oq4�o��V�l�S9��� zZ�i��Cϯ�<��z����Z��v���
��h�S�����B�Lz�z�e�Yj�F�GC��P���h���y{�R�*ݗ98]�S��dT���ik��X���Y�5I��=����Tgk%v43fT���w	��3s'm�yn�w����0��Eu��!)�ՉL�&���(mn��v[C�x+6���o]��ԡTV�.�<^�u�;������Ze�뼛��{�K��sT������^�o78Bs�K�o��%n+}͆�~T0q�|�Թ�1�yN����X��0L:�{�.E^����*R�q�Cp��u\xҾ��M��j�X�`�6,g�᷂�{�z��'�0�p��l�l�V$D�D��n�Rɝ�+b�KMA�ȝ^�gpڙu̗��W�68	O"� e�(��껭�u��@�� M
���0�l��>�䍮�+>(�MNޖ�Ιt���w;��07y�X�]��T�s��V��!]�/�.���)W.͎������ݝ}7L4���ܤ�M��Ŕ2���i��B���s���76��u�E�Ĕz5�v�A�� �V>�vd%��,�|i[�8��l٥��N�/e�J��F�b��{���OE7���vY%CtF�|��ni��ʝ�E86r���{��I�$���߆��ݶ[l��W�uh^gu�ڷ�u�ffm�K2���W�����v�{E�z���N�+2s��mY�mk��γ�˳-�=���+mQ�|�^��+��o��חE��ayݽ�������^U���i���\y��wyǧyys۲�.���[rŶ�M���k]�^em�흜wokoo^�v6�������,=����k7Z�oM���z�[��GG{k�wY�[kBK>���{纽m6��_/^Փk�+�v�K���vebte���qy�^��5�w�,��ci�קxE���<�^U�y�[U�ݶ݇o{�|����_+Ώ��}�Hu���8m֜e�8G�25Y����ٺ����vﶏmܖM����>��,"�m���IryM�i�Z���6^��ݎn��a۳�<�li(h����xq�qhB��m��<�"��A:��J�6����GѤ�'mu��S���t��I��ɗ�^�d��c���d+���]���i��Lb���xݣrs�#�-ڶ�v�%���j1M�D��r���%Tu,����4��v��v����t�p������6�����t��WFc��/�t�rwg:ο�=K���hw��V�zA�`��bʜF��e:�N:��7cu�r�#½�[1��8m��.CrƧ�h�mT9����������1q�zt�v�h��f;S`y#�b���z��;n�Dx��^������R�v81`@������^x-{6}��m]�ig�s���R���k�t�K��oY�-ۮz�N�<L�-��Od����d��OU�M������χ)˼��ˮ�n�f�kם�ۣy;	Gk���ŝ�y���i���p��)�
��B5�m��\m��n#-���䭵�{u@�qg���ly�v�S=�g��:�ks![��-vTr]�Z����śs�\c�:�tj�1��n��gծ]ַO[g�	<MN�1ܵ���")�j�@I�ҰH��l��>��gkm��z'X�n7<py��!����F׼�ݞ9�]�v�a�.1q�6�K)�܇�n}�z맮d��Y��-u�sɶq��nw
�a=ͺ�ڍ<q���n.���o%��qmq��ٱ�Ո�������z����;���θ�J��vˉ�u�[���(Gg�\�wh6z�'�a�=\w-�ݓ7\�ְl��cvm��Q]��y�Ъ�q4�����av��׶B�Gmۍ:����8w��<8bݷp�=.���sx��n|p����;u\&]����Ft��`lU����Jzz�m��wg��nێ<uF^6�n�۷vn����[�\�k�F�P�OT�*c���U#��'���^l�A��jy@�8���V�Gfa����ε��w��>|��4tA�z�v�ϯhz��]�{Y�9�sm�<��-�+�Y�vm&x�k��e{p� x������� R���� lr�p�n봻�k�����7mn�z�v:B��]w]��j]�N��ܔ��v؜Kk��z4�[A��6n��^�^�%���J�$�����۹�nr=��E�p�x���b9M����r��	=����I�d�����<�n(��n�^��t��n���4U�,���󇦵~��O����X[%v�@��}�>@����ǻ�8��c�8�^�<���o��h�S���@/{*�V��R��W+]&��.�x��x��C�����Osm�I�I�~g D�{��l�k�G{�^A��dh���a�wy�  O�ɯ�6|��e�/�ɼ5�^ �	{�����M-��_\����[�|~�W��Zi+�Y�$�~��  h�TH�My��A�[Ͻ��$�sm�=����	�D�υ���@��}�֏mzw�iM��;�� �9����3ڳ=q��s�!�&���l��D�N5g���L�ı�W��� .Ë+���� ��b�3oއ���B�㋾9��f@ ]:�D 8zj�D������ݗw��KI �^��K@��z�p��[a]�0<�72�q5��RW9�6�U.ɔL��ؙyLgVX}�_j\��0y���vb�M����%SV"��ZP&f����f��"zs~ \���� g��� G��|����u浳�=�{ �zU[T�Y�Z�4JD�I�ӟ�$�>|Z��`�WB�-���5�����k4{OO���-��t~]�Y�;#~�$�VvH�$�x�׎� �{�w��w���o��Y3h��䰌��2�3��4~$�O��?�`�"�8#l�j�%�O6�$��6�>���-�x?/Vo]Z�$-�T�AeT��!
_K�z�F��z�xϮ�Fڶy>��-��ˮl��-m�����zih :���Y� ���kX��!��Lc��k��I?y�MWh��5j�M�;�湁��߯xgb�^2�$�i����&�?{��ݱ[�������:W�3�]��U�[
�Y��sz� {��f -ǜ���".MZ�nh�S(�K\];�����[6�Sw�L���(Jٍjܡ�H��h�����%���n�6��W�{;������{���N)�#O��=pK?~�f7�kuTJKR"���v\��b�[��>>�س@�w31dԿ3�vmk�S�||<��"ujPZa�滼�o'�d����V�����C<�L��;�i �$�h�d��W�]2��Oi�h����L�rg��Ō�3�3�[��8�Ĳ;7;��_����ߍ����[�j���m�����@ O~Ɉ�K��н��I�O]52st� �off 7p��6(B�d��rih��\���ھK�$�$���l��%߲kCm�췑uGV��w�oϖ"jT�G��^�3>�}�M- 3���U����y�~�I'{�` �Ԟ�K@��z奕IB�g����il,�V��I�}5�� M_3��$�ڲukUs���r�@6%�v�����#G���E�H=�������7f,G���/�Ք��ܙw2�w]ܝ:3NJ8F��Q�ۭ���ǉ:+{�f ?{7�Q),U�\���\5�$
��$����R	-GI-H���4I�[~�|� ����L˱[��{li���Ƌ\a3��Dw���kl�Z������Jc�pV�KP�K�{��(�'g���m�H��R$�I�ր�T�r��w���� �g8ih>�Ӭ�P��E�2g���5D��3fK����@ >Op���o��`���[�]+��[�{�������t�X�g�k@��IͰ��T��v����? �|���� >���`.��P���X�qf�s9�<����m[�ր�l� MP��h�3�����_�=�Y$]�ѭ�o]�-P��m�0���`I�'u�6J�v��<�k2��َ�� ��k{��2Ě���%���׵��w�n ��ue���;0��ξb��ZZ���ϑ���]3���X]�Z9d�:v�6��f]�����k�{����|~���4z.y0ݭ��W�Z#�� qTQ�X	���`��zɞ�V;n����0U�yk�!���՞�ы�I��}1�^nAv���,�nkI.L�nQ��m�Mۍ��hc�%-ݍ���޷6kq��s	���z�{1��4M\�F�kOtskQ�b\���`۴�;c�Jy=mg��%6�^/;6XÍ�O;���-�Ͱ��8IN�m�+�}`[<zx�8^�f��wA�s��o߯���3jUR:���/K�Z o�浈 >߳�L�ɝ˷EC�v��F�w[�O`X=J��Ylɇ5�ŉ` ��M�\ޓA�4�� �O��3X�6o��Y� ��N��N+��A�N�v���p�]�s1����,�1#͵�kDg��$�+�D��?r�IQ�ku�rJ�f`����Nd���'��� ��&I�{�*N�4I��Of�V�1ǃ/�hTI�5�ͶMF3{�U�Gg�{�Ř �'��e���gl3\��B|�d�$����I$��h�9{�W�"b���//6�d����ӑz�{ch��76�gpct�zE���ߙ�uw���HZ��� W{�f ���  hOf�D��NN�ǻ����0b�{;�3�=�f�d���#�;�lJD�J?X��"���FE����39�;գz�Rd�J��V����6d�uAJں�̲p�8��.�n��!h�Rג5�N�<=� 6պ��� �s�Zo B��ǭ���f��hvM�N�P�x��2�1�=�o` ��u� ��b<��ى�s�&�tOo���I�^�с}��g+���po�]��z�'=�us`�����|���[������.���L��f� 5�Řݹʥ����N[�0/�?O�7�y��X�c�׽Ř ��-���0�Ꞻ�k����q�6����E��u�\h-�6��n�zU
]��Y��4�|�����т��b��gw���` -�ᥠ$�h{�tJ�Aև�4b?^y0�o>�rk��qk��jv�B�g���$�ej�A'���z{�G��h�h�������A�m��I�N����K)j�W.!z\+oH����%��t߲@�^��J�af�h���rvF�x��9��$EU�w��=onZ\��ʆ�Px�EW���a��L<6��6�hTL��^Da <=�{O���'�KC>��s3W�����-�kO�����C��Wn�{��g�$�}�H�I&�9����I��P<&�'�{�����eZ���r��;n�/g{��� �v��5�I��4d�9 	�ڗ@| ���1`��޳��گk[������c����S7Y�]�(�wa5���v,��&��L�����~����@�����E練� Y��>��w��jXԶ=�x �[�kA��G�!Qڜg�{z��W;ɘ�^���	6�Ȁh�'�ZtH��(���1M�=����v�B�������]���1���}�|�y� ���o�[;٣��@؅�{��� ��m���z�%��9UˈGnL݂[�{'Q V/D�ğ�?V�(���$ў�'n�=m�<.�pp�,vj���ʼ�-�.f![�!`s1R�ƺag
���d�v����YͽoAC��4�MUbD�3�2�j���((� ���$��N�� j���,׭��	��T�^G_֍��$�6e>|�.��$�I��d�E	�H��յ�ŚF{�N���N�١s�֮Tu�|㲞��p�!���Ki$��k�G����;oO�s��{�o@ �r] W�f�^���,������v��*�������/�5����ͮ��yb���5D�f�@� 4g��D����)k;��.sa��$%!h�<z�^�, '�rk@ G��X�M{~���;��o3�> F�ɭ��̨��ZZo0��&�z_���J���I%n�L���rV�o��\�{,D|+�%=�c����Z�X�WW�ܘğ��wkn��B]LZ���/����pc�w%x2�*��N���[�sdK�I]n�Vvd�b�	���66.E:	����5��#z86�S�s�+R2��c+�Ƞ���!�d��_37���$��d۞��W�e�,�'��+�3�:�g����j�9�+c��2N���k�'S�9Ŭ����i���n x5n�3��]t�RM��:�u8x���l��,ۂ-�s���Ko^��Ge�r�r�H�:�}�����kj���)��p�9�'��#�oS��x^�k�n��Ý�6{vK3�Ϝ�U�9۝����	����;b��=N���,���-�������&�`6�2�O��5A�93����J"�@v���C$���O�"j;e�4�yv��	��L _%�N�9��kC���o=�<��z{���M#���v�S1�+����%x�jS�F�
�a	�'���@ ��s4�Z����x������c���������+�6���3��94��3��|������{��,=��$	HJ�XL�����e*j�*$�\u
��D��{��TI����@�ɺ�;�8�RgM}�����-����{3y�|{��O���w��z] Oƽݭ� S�Z���h�~�+o���=�(A]C�g��\�16뷲m�8qjp�@�{}ꃕYj��U���K�U" ;��$�O�;�C%�ƺ�}����iۅR �$��kAװ6A�b��0��O�kC��D�o��ѕmF��S�FPBX�׍�{&I)�5�uS:��EMN�:mEe�X98�:)I���fa�t�k(�Эb�/�|�ή���Cg�>��3M�~��Ǭ���_L�-닛���-�4?+G--��ု���0@��ǋ >7�TȴE�OTV�9%�ND@v��n]N[UW���j���p�|���4�{=Q$��kt���I���Cd�Oƥ�_�/u��Y��$���k�w��R,�����z�ŀD�gKʹ��9w��(�=;Z�'�塀�4`�2��Pͨ��Y~���^������	��E�a�	�]�s�&۲��m�^}r�VZ[�mw�2&[IQ`��W]�,� �o, m��h;{�OUVznjk�� �jo(���z���&�RWk�p�}A ��&�dн�wZ�� ��m�| ۞�_Q�4������]��-)L��B�t~83,��<�� 'A�*��I+���L=��F�Cd\�u��[�n�a<�8�&|_v�ߊi]q�W��p�P�,�]׏�_(q��1��]{���[�7gN��ngf,[Гw&�P\JhRT��\�w��]נ.�ƮS�sK*n��-MҹI�B�B�Tw��_M5wN���-^���_!�oS/��r��Һo\�X��8�׊C3�K���f���	�-�C3Z��x^	��aZ�]�W�/XYf��n����`A
$g�;S(ڹK�޷Y[�VKf��rNP�޳b�Y�����f�d}ko�_��n�9�K�;1�� ��K.Z[ɼ1��<�ճ��E�U�u�&���gfm�U���V�S���u
ٺv�1δpt��ɗ��a�eŞ���.R��"\��yqz��݉}�,�*�|e�ZwK0�J�Ԑu����BM�W�[Fu�S�T m�3S��Z4r^3���M�K�C���i���\���D4�ҷ[�}�{{�P\lgn��A�b����Ik�R����Z�+G�5+k.��6���{)�ɫ��݋��#Yɦ�/xn�H�$�z#��3��C�Nb�����e#�d�b�*�

���{y|�Xg����αw�NB�)��u��gv4�|�u��m��b�u�X��N�S��n��H^��nX�O�b��A	g�JE7K�`+����]k(6�U��st��I m��ѿ�X�G�Hy`�D
���u���h�z܈�!2nH�M�T�d�f��A{6��-�[b��q�h���R��4SK��O�o���2�r�����n�F�m�����0��gq��՜@tE�D@Q�7VQ�e�jγ�<������fS-ie�6��m��2��U���.Ҳ��Gagp����$��cq�����"$���n���K;q-�9�����C�-��d���k2��9%#�HN��״FٴI�;k2đCkt�8��i�X�t9��$D�+#��:G@�k[g"R9;l��9K,C,�i�%E�m���٢8��'#�����#���#km�&��9f\-�$�-n��7.٫J6:ƚp�&Nr�ɶ�wu�bƬ8�fqA8��f	D����[`�ٖ��eknȣiB�X�iMz�ϱ�g�UU�}��]��J�j�U���aIpρ{]�2��}�WX��A�r����˷&�&����n��8�D��J�;.�J�S�T+e�����Ҡ@���T��~$\y�՟v�]j-Z$�I��r�5��h
;����:d���$!5<��&S�L�P���ne����\�s���h���5�;F�I�I�5�����M�* ���� �������eJ{Z�� ��]�*��2�FKm�P�!�W��͒A�[�xy������v�  <r��| ��3M�N���cm99�eݔ�ݪ��P�fh��ώ�qǤ����`�	�<�ޤ.4��Oē]� ��k���{�T�O�통��\s���nOg%o����D��t�h ���9˩qK���=pWX�I�6C9��m�ɹ[��c��ڤ֡UHeTL���]��NNHD��x�-߽4sά~���Z�3Qܣ��=���%���\u�X�U���aIp�^��Ř؃���-5�RH^٭�d��>������y�1������e�8�z)�ݵ�[u�Uz��z�ػz��&{1����[ڨ[fg�Խ�u��U>�(��^B�^�- oGM�I&{��%d
��Ћ02+�i�� k������D��K&bE�s��&�|o׽��V
R�$@$��Ѡ}��M�j���z��ۙyJ���&�#�[
���|
�ϳ��:dOeE�]�S���I�I����w��,��w�8:�UrWk�pW����ڜq{vI��[d������@|�^���Vw�أ����O�͌�RE>+��G��b����0S����A5� �5��t� S��G����V�Q�Pݥ�&�����ַ�@\{�;Y�XSw%��^�������$R�|�8b�|~Co[/Z��!���_,S��>�D9얪�ɃP;m��b煻m���y����&׷�m�����=�;���bnh�����E��up���g;����m�9a�ۑz�zs��'��7���nN1V��(�U�nH;+��0Fv�su���l94��U���:��6D[3<����h�{%ه����&�q��l��9�s��2Xxݎ��	p�ib��a.��^v5{��y2t�k��K��lC����\M�u��w;�yu?+JKm�%���뿖a��wU:d�5���뱆��!�5푿�bs��,���S��|�n�,�_)�q!i���J�ԭ�c0������M(O;T�$����l���5����QQ�T%�&?\�2i	>�q��Lbsע�1�:�5���l ��&��%��r`�p��2��5��;�Ӛ�9��v�$����ɢOğ��y��I�^���C�n(C�Hf�!������s7�[*�J�w.}�>��H���ӛt��?i��k`TI�=Λ�OĒD犑�k��uL�E���T��ے�Za���Q�Usq��ս����M�ur�gh�D/Z^�9�~�������ص'P��R�I o�*D���y�=��{��Yκ�y�b��>s-z�V���-��������o�眾ߵ��w�Z�r�	��b�f ����l6�c��u���@P��&]r��q�_�vHw_+ɞ�Wqת�2���U��H���` > =ܷH �7�1}�>jBQ�xw8����^��'J���l��s �o|�I�&�ir�kz7�Q�h�k�� �hל�tɮ��^r��"ۣ�5���Y����z >�^�Z  ��s��@��y���g����Y[�� Z��Zsk�#����#�������|��ŅҠ��S��$���_h�F��[d���� ����}͵�7mm�9�p�cr������l���c����A���r*߿�]��U]����z�ր \��>� s�oX�~��vY���|�k;4�1[�sY���6�iYC���ay�q����̻����M��|��X	���;\��M�57��<q %Wk��hK�k��w�� �n�`ؑ7w�-�m����P��jN:�1L^�y�"�Q�4��!�W����轥lCŷJg��9ev(l���Z�ő�;sF��D�sk-�U��w�&~���}���'�Ey���d o���ٔq:U\-��5�̺��7�^q�Πn��6h�I�w�� �;�~���Z��N���-_s1`o�z�����K1�>�h2~$�4;e��n<^Mk�P���3Y���[y� >{r��\Wf����r)mr�R����[�9K���۵�o�|w�8��c�P"�B'g�ژ�{���F�8�#��
�o3 o��y���'�w��3$�^J�5_���y���2ϐ������͔eLV�m��\�v�D

�{��-��F��|٢M�{ @2I��w�"k\�k���f�Y�>i�J�����ֺ^w\x�l��Z;g�9t��Ź7y� ߻��m��G=�KA���]�����g��;�=�e���i��ھy���w�.�6!w7쉾e�=N�j�8 �S�n^]q��Pv7F����7ӻ��*D/������9j��!ά�q���3 *"��I̓�=㤟�f�ט��[}��n�Wn�׻5H��MQ4��HԺ��H��&�|L�c	�&�?'�$A$W9�Й��e{?��z��c+��'�s[cϮm^���>z�J�p�����_'KA�e��;�#��u�}���{7�k.���vQ��Y�m� �wk�s�DrBƎ]��X��d�xq�|%Ӭ�^��1� >�v��B���Ń�צ���&���>� ��[�c�%��k�[-� �^�T��xOw�vԀ��% ��ֆ$����İ=��A4� *[�"����緾W�]g��=> �v$O�I#�֟Ē}��R�]��oH}˭˦�v�����{�� A�z����ҜO�����*'q� ���'��A$��塲F�9׻O�x5U8��<��Й��h�)�@��6�r�\�j�0�eɘ���]�)���b�zط����"9{�+*ԭ'zWy�S���Y��#��Em���.t�k���0[G8�Z�:�����mkg�Ӌaºu�׎5���=GO��-��6^N���[�ݞx�K��U��vBۤ�b�ӗk��n��I���g��
�n�<L�[j��4��룶���c�۪�������֟�O&C���;Hv�����v��&��0g	&�^n8��ǧ qۭ=����>�U���;i��gf�ٶ�C[�4�Muo\ڏ0{[�6�/#�y��+�&��<&׋������B�U�����o�@�����j�ݮ�&��[��[8��bD ~�Sg7T�����a#2�+3���|s&����	��rH���- *t�$�{�Rd�b̜��g�g�1�3����)dy�����lA���&"#j����t]����� 5��5�|ﻮ<o=�+��T%��*�pnU9M>��5��k�~ϳI=ݚ���~�lw���MQ���L�A�%`�w@��-:9��?�$��|�|�������	i�h�S�P7D��@犩�fоR��#5Λ=�:���6�nQK	�;�Ohҽ�sܻ^�-y���T�V�����E3�7�a{�浈������ ��f�oRS�^�k�F�2	&����[� �]��US��ăr��	U�'����������2�MS3)tq��.�M��w��k���x��A��Z������ZL�w���T���[g������y���cb@{�������~˯���K�h��^U���������,n�*����#�޺�`�o�2�P�|^<UĻM %~�塲@$����a>}�fJ)ly���[�m�o[��������	 �[�������oV-?a�� L�o���|��P��yW���U�;`TI�k�9�ڟ;y�]�洁���I���x��פ�l��w�k�{k�霜�����h�UQ�8�hE�'����a;<�K�5�4c-���q|�?>�o+I-�k����|�ܺ���y&Nq�%O=Kz�Vy��5 �˭�ⴲ�K\�@���M�~W�j�f�(���!���$���t ]����b�w�g}ɣ1-�|�� ��o��6�UN[5��˭��",��a0"��+3S�������50�X�.�+sM+��m��Zͭ���N]�:��M/���)aλ:T�t�a=��) %n���k]�m�4?U|��|��  ~�]-@���f�枣��2�0fY�l�E�T��ԽW�w.�����@$��Y�]7,9�6L��vׯ��zDb�IBE-�I>m�~&{�Sgٔ���{��H>�.� /{9�� ���qf|�}=��;�^�]����H��N�-B��vc�$�[^ۡ�q�j�>��m���w�^^N�/֪J�o�M�ց ���X����qcg\O�<�Ѣ�^ 5#�C�7D�c�N+-�����Ř��>g9����M��@ }�{5� ��{�1 ��w�R#y�Ĵ	z���K\�׽����绥�� /<�e�ܧ�!�sW興����d���� *�o������~�No|*��M���π����� �w�� ��rvo�4�C�5>���G���x�ɴD�Q��]�j)jy�ҽx;�s� ��7��~��|=�u�Gm�k���
b���<�i�gz��B��U(��j���u���K(�a�7�Y��6���KG��^I�W�� N�T����;��Uq�f����CpX�a82��1�s[��1r�ר'�[�ɗ������vU�gW���"�qIj$E������,��;�,��  ���'}ق��XC���DS��6��Ř��VӲ5HJ�V��\�O��}5��Y]�٢@5;��I$��;�9�.D��XZ5sY>Bmh�vT�-��s��.`��'��kCf������-��Ā}��M�$�E��z�G���J���w�z�9�w��|��K� ��j]b4�<��1!�׉d8)�Lk�'D�X�]	�%n;Lτg�4�6���K0Moվ����I8��0 f�y^  ����LK=X���(�}%�Yu*�6!�k/c�q�0��a����~���/��Q���MgszT7�l��*{���E�yV���]�%\���S�.C�A �@t�2�㦱��5��ǘ0Q۵.��B��{e�:(9'�5M�!�ݣ���:�Z�j�mU:��H�
Bܱش�+�O��_!�% S� wv���;D���$��qr��^��̚�q��7�ovh�H�ͼ�l��e�{мVٹ�S������KI�w�eV;x�����C�W0��I	[��q{7^�ɩ��U�i5ۦ<V��pZ6�	}G�˹�L���Ի��>��3��]��еY��`��x���c�]����lwU��K��ǩB�O�!�h�v�ŦMQ�T�	j݃��gǷ$�f5]�7Zs�����-����h�u�eˣS�"�l	��&TN]�`2����yD�H�V6�wZ	1bAK9^}v�ͧRu�i����.��%�.�S�2�����B�뫔!�H��xH���N[B]M��!�ʪ���O2�%P\�����9/�,f}ö�Ӡ1KsP1f����N���y�Sq"�ٕ0cj�6�f�+ڲ��-��{3��ύ��`9��k}H}�ޮ��&�թ�H��)9����4;x�Ӧ�f�9� '�4Vq)���x*l��h��S9H��16����MQ4]:}u��E^�hG�w��WAN7ӈ��S0��refTz3e+6��d�Ȼ��-x�N��r�����q6��;������k��y�"�L2\m�V5EET�,\���kn��ͫm���Jav؝i�Yaf�af6�ӌ�-�:�޴��\�l�m��Ir�jt�����d ^�����Fn)F���mvvۙ��B"��A�a�3m�q�����%I��ێ�"���Y�f�,�tDP�8&���#
5�{�y&�D�˓��N�n��TB#���m�v��'$H�n �r8��m���8BI;��&w��(I6��8�����9	[ZRw"9��M5��{Y��mh�t[on���a�a8ڵ8 ��dC�N%3q�mɶ$ᛙX)8�,��n���˥0������E�zTд0b����4f㲄C��=nŎ��J���.qY�QƦ����؃���u�m��\p-�[�v|�P�֢8�{`�	(]�J�c��E�����������=��m��W+�#��x��Gt`��mo��|7���w#����S�j��J�Ս�7�^d�sţ���.�a�tc��7n���Fm�6��a�MV������.��3���6:�����Pv�K�)��9w>^�7nh��l/���J���=�n{�v8�6{'Cu����x��t��P�#�H{u/n��e3�b���D�Zm���8��m��z���[�G��wS��]���+�ݻ{m%��
�d�HK�x�o\������mar�<u:.��7NsI���[O	Ҏ���a�ً���62.���{s�b�l*=k��R�b�p�lk1�m�7k���[�۳����d��u�us�������<�݁��c��{nc�v�+��S����f�筙��m�<��&�T�:�<�S���B�:NG�3�M\#�,v�y�gZ�l��\����v��\�e
�9mz9�ɲ�@���[n]O[<���)�����D�c;�y��Xf0��A�/l��nM�'<���x-�*� �=�z��BT�|�@ڞ�燧���q��y��m'����:���g�u>rv�t�ӽ���ۺ�Rn^�q������v��<�/X�mH��3�^[� ��.���nƤ~ώ��7)��hM�ֲR�>M;*r�'`'��7�	�|��B�]�Qj"�[mD۵����z�;Ki�,�b�M=��j@���e赭��d��]�����z�[�&�z.��k���j��n�i�mmOm�W^�i�� p�I�΀q�v�n�#��n���gۖ^viF��{h�2������PDTun����=���ϥ�٫FU��T&�:۷7�.�e6�0�m�O+��WD��:�]V�uz9��̝mY����M������|J^��ח��{1�m��v�q=<SB�\)�rv�^��������=)<1�Cl:�F�i�7��=����C����K'n5&�\Ep�z:������ W�u���Ѵ����q��筶�v�N}�����^�8G�+6�B��y d#���]���cκ���ՙ��f�݃��ݬ��g��u���i���Ocb�ͳau�Ä�w@���u*�����[\�#�����c��=1p�������Z��bv�{�>9�k�O �y���@��y��5�#��"�����������H�RZ�lz�Z�b�on�RmX���_�F�$�r�D�)��l��<�$�^��4GTI��e\!H�Ԅ�ei��ހ \�wa� ��j�W��^��� ��SKC w=����mZ���%�ְ�޺�KSYf�~����zW�>>�\�`6{��^C��jM��^�}�K���+��J���=��X��r�������ٳ���&�}x�4I5ܼ���z.�*lN�����O��e�X*�nb�fx�t����{6����8��Ǳ�D�D��\|�T'Ԋ��5��&��|)���$�I��������F�=���6υ��ً���s��E,P�ct}9@�D��37�~���!�|�\��y���|莰>+TA�,��r�]Qquqsc�Y)�C,���6�����A��_ϼ6�44"j����k/=$��u߯���UUT���:
�*�{�^�$�5z���
���Ț�dۺx-Ih���|
�w3��g�� *��ۗ�'N�ڢ@&�f�� K޹�0��Q͍H���U2b�jm>���|ހ�k��a�}3�� l��J޵5�+~׾7 ^�3�����Ken�Z�k>/��i����c�h><�b�4�I����D�#O�ҽ\�w��L�	��G���),���ɮ�S=W�۱ٸ5�7J'Bh�m���o\3��o����ҫ%��{��cm��<P�׈��e�od�jy�����s�b��U�"��M`�ߢ��^�{���h��sS`MT����;}5��^m�u]�s��|�����N�=j$N�K���N���Cٶ��MQ$����Yu�ާ��sU,)��ڠS��ڌ��������t�/'�L�[�i`y.��K��h�]n�%և��&'L@X�ӼC-ZR>��N�޿|����6���4�{7�=X9ed���j�y��y�W����ro�/�> z�]$�����C�p���e�}��ܱWc(��s��.h�~sX3&��Z��|����$͵�?�$�G�֩I�ڛ5u����2殓�[���!?�#NN����X�V�;� �����jE�>�v�XXK��ꔥ������}w�� ���� ��q��8��B����^�B�h��m�^�3NWU��J������قto�[���ŀ�r�]�5�s�Ń/t[v)���{��5��W�oS�
�#��L�#7�^��w���:�Y��Yu޿y>v���#��Z}�f`w�zD��I/�0�^����/P �禾�k��5��=�3���z�ꪖl���22��P&xC��9�Mm�Ӆ:eXKB̥{��X�=��ul(���۳z�v�t4'����j6-�y���L��œkA���L�%+$-bf�f�����dS���I���u�46u�$����f�I��I��=�ޖ�34��lM��H N*�Xinzփ���3��6��@���d������n4�e��@$�wk��D�}���7��\*��2h�־D�&�}��&��v���U�f�#^��*|L}�����5;��  {������񘁵�l��Y�U�,��k��Zݖ�L�7��5��t��m��0'�H&m���?^mh��l ;�<Pl1��
����Mw7���'��|��Ns2�	};�d�����J.�����Ў��2&����\�E��N�`,���9d��J��	����9�r�^P�kدȡ��4[і�a��ݘu�dWB���QC�#������b�E߱U�&�b���t�|�%mn�n�n�s|����.�6iIHA�~��ᤷ 'f�睅���Ϙ��|�JkAu� 9M���h��N8k/F�e\�m��Р�t�#v��9z��\��6㚣�z�I�,��X9�:x|�x�<��<��0� )�OG��
�5/�\x�l�N�ѳ۱�ێ�(80��[��:5���x�!y�������8��]!��c����N��FS�3p=/�ml��l/3shsa㊹������{�����'�O>7[jS)��5�7m�{��";@���'����cm���i��=��ROE9=R��pa-θ�}ʺL��
����S˱bV⚜i=� WF�Y ��X�J=�ޜ���Fgt�������U�]+�4��6�r�ł
���j�=u�A�s��Iw�Y�{U5��j��D�`�&Y�&VE�;��M�>4�	$��U�O�O� �OD��o��r�B�b靖�r��`8P��ؾ����w�w��96G}��/�T�POމ�=�{�dl_�������6�4q�Y�`z��.j�'�u^�W/#�S�6�l�[[�;mR)]rֵ��|ʡ@V�n!I��:An��5�V�-&�[�施w�KDGh�z|�{z�V��q�~�Ve��jW���z�G�[u*�}�7/2��f��
����ab`kr|��7뚗53QT!��L���)%ඨ,����P��ˎ��,-�n��`V��G H�^Ʀ�j�:�Q�K=v�z�{��6�W�y`�+����P����^mZ�%u�U%T������٭��i	���� �j���蕴$�jݎ0	"����5�ݲ�%%�T�3�{�w1�����t	��n���:	��3	�'�s��_G7v��&՞b �EQ �ۆ�o]�c;x���p3�ی��8�Cfh�۵�|�>����Q4$�G����	�<�$NtY�y�M�9����	"�VfCbЇU�.���fo���c-m��|��|׬�I�͵���d�����DǪg�W�K�Y���0w�EK�P'�:,�NxJ�b��6����@[v[�P�GiӷD�Ӊ�gY͢;�C9�۹��ר�"n�.��T�`��^�D�W�Fk۝ґ	�T�f�CuK����+:�bm��xZ^��ب���GQ�K;����9�b`� :���<_@}@P��uXp�\9g|iՁTwco�+�F�|n��f�E_�Nt�S�
���M]��&�_fH��,�|����=���a�xET�L��>�JA$wj����x�]�X3���*�>��_ّmEt��֛� �Q��|O�s�)�1���^�<���*��A��ʲj&����C�V,��w�D���e/Y �:z�X��e����8��^U4u���bDT�U@���Qd��Y~�6��ٙ|�i��I�ޗ�~$j����o�v�J�Z='9��l���i�M�@��ؿA }�d�:�{(��xk9�^^��fnuOn�3��od[�$�j�;���R=xּS2���ɞ�h�a��	Т.�:f�8R�NR/ڴ�'x^���k�c�V�+F}�5�	���ԉ�a��>��Q`|C}��B���<�n��k�Z����9�gn-/<�EŬu�7d�7$��r	����Gk��3�]uۍ ����9B�U�����٦�m5�<�`�f�`*UC���J��UQ�m��^�sK]�ɖ�IK]��u����04�Ip��,_l�F\���V%�O�*���DWi���3���P��ꩡ*&�1Sd_5~�e��'��3���q4'�� ��.���� 40uF'�5SUT3:��i˵ԫ����W�1 9�����r��;F��[��w�+Z%t	-���c���Ѥ����E�x0
�E�
��`P��hd�2�	AD�t抪f:af�܊�vNH��-d�t�jY7�n��<qN�k�fb!�Jj�UX�7b6�jPSj3Dc{���]Y����(�o��q�(TXRw.�;X�la���.u�{<nf4�{e�.�s�/"+p{vθx[�;+����%ʻp
v��V��e�Z�۶�E��:��k���W=���a��Cl��v�s�6vd�ɯn������q�m���Ϗ|���q�Ӯj-�]���{j�9v8��xq=��7#��h��n��Y��n��0'������e��p�8ї6͜��i�.���Z��綍�n�{IӬm?
S��p!������MD	�B���ʲ|{n{�:�f�6�E���@��v��|�=��#�rk�,�YiK�}۷���w���f�==v	![��$������wםw��r���T������UF�T�f��	��B�$��|xNIj��u A�չ����斛�xW��R*K�,�k��r.���y[�Q��H7M�� ���b� �k)�Xk'B��טlP/j�Ϣf��h^�W�'�cyw}/5�˛�.(R��O����A#�*�5K.M�������g�u&�8�vY���qs�m�Û��>�.@P�����b��U@���9{��2�n��I�t�b����=p����0�O���ܥN���h̉�1h2�y;UT�aa��{$"6�RGt�S�L���������E-�`�N��%x����^�q��W��G֑�;(X��y�s��.���@޷b� �G:V,k0�åG.[���~�EE
�����ؿO��NŒ.��;W��M�JW����KV,�j7*�Dɚ���3Y���]V��o.��]2 ��I�}V	��eed� �a1ۖ,6���n�T���K>��KI���gٽ���x�Q�&� >����_�-�Gg�O��{��l�R�F���A�j�bc#��wk��\�M[���9�@.'�ꋇ�뾻�Q��S4y_e�'ĀF:w�g��z�f�skH��ؘ�젉��:w�*�L�ύ�a&�0�7�#�]{5��ط˨g�$���Y!�,�!	�q��!f��D;%y��w�Tnu�+2�.���qJ|�=�����~����VK[� ϷZ=z_r}�gV	yg��K|�¦�<��E�*��8�f�[\e��L���]8]+ri�`̱�Vc-��
{]��vs'2� �CN���i�qk��M�(��!V�ʆ����n�x�Ty���9����B�k����^=N�1��|,��mf_J�˒�]��d*��aK�r�:Wn��z��t�S��)�)��]�}XTelY��)W����0a���\l��Z�N���k�V��]ʮԩG �����Mδ��	�v�����
��*̜;Q��W,-b�j�ab�=2���7{�[)�(b	��f}�1SN�nDD�s+���fn��la_GßV;U���Z
t�3U���M�����}i��޹yY���.��X�A;޳��4�_��	Ëw>�y&l�ԧb�(헗$0�J�mhV�h;/,@��:8¹�7�)뼗��\[�\��3S�]�a���eh\欨˻�����2���u�ti;���n9*��R��F堁�Ȃ3�o����K٫�︤|�3���Y�6��r�2�z��l���մۮ�5�:�2�b
o���3�襤��n�b�f2rv��p�R�c�q���f��Ôr��pGo{QYIU�n�*^�]LQ���5Ї8�q�+��7d:�������a�B�n�f1]Q�፝sU��F���6�$KL�Z��5�	�J�a��X�V�ݾ�%8�4��eβ�u��;��ٌ�,U�EVG?܅��m�'�n��ٓ�A�F8Hu��
#�k2)�j'8Skmnr��%%-�"NN��f'��k8���6`3��ܸ�6���;���Ël3��)8�:H�9�q�RG'u�i�RC��Ad�P�f�n�'9�ok�)�۰�$JE�.F�c��9�V�n��m��om;���S@�$q�VZ����2�P�V�Yם�9u�{���s�Ci�m�Ί���NA擑��w�M����ٖ�f�H㓔�Ӝp��<ӌ�e�,��9�%j�2�Mےq�&8Js�J9���K��gv:f8����J�A$%jł	{٘	��zJ�bv�K�}۶��>Y�����(�k.ŐH$m����@|�Mv�/�"OtK��L˺��r�]�ޓ�t���2/'�MY� �!B���f	}/b˝T�K1ڊ=2b�EW:V�Ivy�d{.�um��H;B�C�� En=��6��	/}��v;T�e��y5��4��o�l �}
��k�є��J�z�*_k��X�x�閲��\���}5�I?�P�j��혀�˹�({�С�Q�h�:�g5����/b��U@���˯oX߁��ϲ��&!�m��O�[��M��}3���/9B;uȥ��Ϻח>0��y����� ��/��B�٥�^���:�2igf�nkg�FAhR�b���-��Q�W+��xՈ��3�hi-	�%��]�	1�\&PƗP=��N������p^$%ݹ�'�cl	� ��USQJ��4�G*ww��]K�Oeb�� ��<i|>�f����+�����%
��4�O��>�f�m�l��ݻ��q�g�R��',�������Y\�<��s���<g����W�����W�~�d�3t��������Z冢�v����}��y�
n/B�݄�"i�_Z�\�� �ҕ��q��؉��t�a:�3S&M����/"�Ad�B�t�%�;�Ltwv�A)N�$���Y���r&��7y�!k�"}K��}���Q!�(� K���zy���w��F�'ͣ&�i7�^n�tq�E,f|�u�6�y��˪�d7\.�h�sYA�=�,�f`!����Q�Fz�adDN���3fխ̬9�����J��(]r�̽�X@�C惌fr%�U�b{I�y�Pdf�¢�Im�Q����t*�^�u���N�Wk���u��w%������s�דg������$,��4hav�˺֩8W>_:8W�+�P9v�	tm��d1n�}��cX.�]�<�x4GH7���[n�kn^+r�����6n^�E���9c�n}�׼���6�h�K�o��v�GpF���{i�]���UF0mJ��6���;nӊ����͍�c��ф�P7(FG��x�� �e�on �>.N {Z�����z���uKe'��l�I�Nz�6�]ߵ��ˇ.���Q���ϲ{�õ;S`^�ʻ�ǺNt�nb��y�+�ghA �ޫ�v��/�34V�v���Z�4�Xd]�� [Z�M$׷�k�6�o^X�΅$�b����p���X#�ɧTm.e��4o��7^W̭�v�I�Dw *O%H|�{SN�{Ǵ�e���^��-?]��kD�����;�H�OҾ�4����;A}V"��@�}�^fx�_KQg�[a�fM�O���7oi��<g��.#����-�8b�u�z�f28EɷV�	.f��$N��"*��Ѯ�Ii��n�=�ĀO�����r��ӵx�B����|�u���%JJ�2�JM�};�**��5�y��W6��7�0M��e��:"�ֱ��3bFգ�g�$^P�vU�%��$����cD1
�HIpoWW<���!� >��0;��W�/��F�ȱB�T�ױs�0&љ��}�����=�P۸u�f�6��fkO����ې3�%q�YR&b���Z�7'p
�yxA� GR\��w�V	�[��9
���dѼw���V��T�.]H��>E�u���$�-E�H�J���q�8{Y��*)S�؄�"�`�"%n�$�ՌғJ�(�("��ddqZ��eN��?{�Z�%C,��ǘA��Y>$z���r\W_.\xmon�%�j,�Y�3$В*(E	��.]ؿ��a�ҡ��rĳ�I�:��X	�X&WF�ka��sОn撲�2�a	��g�-'��;�6������.��k���{ٖx�AQ�p3jV���1�B�NV��Y+�^�>f�k��ϓ��#Y[�,|�x��+^U'W��f�9.F�Ϋ��	%��P ��jC���"�̢m����°IOY�r@$�q~$�H3�ՐW)�����C-q���zl�d]�]+�M�� S��P�S�{T�u�>�����D�u�X ������k����Zѫ��j8�+%+P{s4c���/�V�E�3n�I�4}F�-�����gl� ��34/��mŒ	"^��|H���l��C��:��_�>$'yز�8DD����;u��,�\��{��m&�`��#�{/	1':��Q�;S��=�ݒ7Tj�C>��kI�k��ω�v��)P�tuF@>�]v	>����ٻ4���e$���٩��/sb���<�d���ω��/<O�/��7��1�i��)�����)�s8sb��_UAz�Va����~�x����ze��٣c�&Ӗ�LA��ˮ��HM+*"������1y��1wx
ع!�
y��м�y�M������i�(\��˜+���t8�0��{`F2p�ݾp%��7C�z��I��Q�������	��|\��Z�M%�������$��9-���]��Zde��A$���Ś<2�z]V����ͮ�}�ϟz�Y�Y�%Z�/6�
�Z�ۄ��l*�9!���ۡB���W�P~���k�1m�8]*�q�q���(�e��wZ���=��6�g1��\���d�uT�8�f`$��<��+��n�*8�(�>���ڥXx����Wna ���$���7[x��U��&�K�緘����J��
2�M^N�@$<����!��x* �w�3����D�V.���2f%��1��D���"8�t^�5^�u�Oi�ޮ�LOz�Q�����׎�h��UU�3,���VE�m;�r�Z8,�k5����׷����ϰ�<���m�Nѳs=�htu���.0�';��d<�`:�xq�$�H/9ڴ��8��=�Mm�;�l�&�죰
��ۏvNex.[y�	E�ܢV�m��v�N�ntA{s�r��ϋ��k�[�7f:;q�`�\��t��l���;�;����ϫ�Mͫ��:�q̝F���[��ȶ����c�y}�:^+4�[76�V�`�v;�a�{�L6뒮T���n^��sͤV��NI/=�V�NY$��~���co�<��ę��r��Y�n�#{�he�[ō��N��{�;�H�#�؈k���v��W�s7Qn�N��A"y+��Ga@V�[��%:%��T�o]�7�k� 
o�!@o��,�ǡwQf�� 	��*� U�u!U��
�~,�zw^���٣~|��|�f�Ҁ(o�@W��h�=g�׵�Ô͚ms���"��R��3kS���OǛ̾���ޓ�X*�Y$�#{�Y v�faل�2dGR�y�B��hA����a:�RSeA9�rQ�l�0j��Ǩ3k7\�'w��Օ(Q��M����m4s��b����l-��N�&����*�
 Q�u� r��5Q0ԙ�������|{���h���kg�
zn��;^*7���Wk��jhص�i	�k/&��r\�n��]8+�3�qֺJ3������2�!SwQ8���	������ �Ƅ\���}[��N��͒EI��B�S���B��m�����y��'�]>��G�ڴ��fkk���ݥ�	]��Ͻ���{̯�[�m5-��m6��`$��k�M>U�_^1�������sD�
�~,�j_k{Ɠo~���ɉ.@�5�ﶫ��Zud���xI >��Osj{����/f���BTEd�����GGA�WB�vԉ�UB	U�#©;�s�ج>�5���7*�Y'ǛY�I$wmq�8Y#j۳�)�ذI�kY��f�fG��U�N��i�~�����8����vI��3 �;��߉ �,W��!�J��D>�˧�vhf�̻�]�Ә���dO73{��p5�]V��:�Ko�P�f������g��a��Y��Xٙ�����F����u��4E�^��)�mx8�39�������	�3� =9���6���|��kvvI$r["�Y�/��_n�� ��טHke�g�<�CY�۶J�$b���O*$��NJY*�^�>6�i���KWy�o�Ƙ3|��'����Y$l�|b�7A������T����kv�%v�w.�f�Ip�*�������_�P�Z?'u��}LP&��J���Oec��̊EL��L߉��MH�>���`<��'Eם�1-�յ��>$�;��B�]w�o�<�\�nZ+-mtL�/,�&�����yL��>#euY'U���W�Eg�ZH'�=�}~!N��e��U���UT�a��C���=��1�<��(�
��`�o{r�p���е�gj$3΅��YJ*�N�^���{(�W�&�ܞR"��s2��u��P�Oq�Duim�t%N�K�gj�)*Ot�o�zsf��p��"�RK"!�ֳ��� ��n>�"�1X�x�����M�����Ge�N�RfD�Lll�ya+��n,(X��(���ϟZ��k��ꋌ�D��j"I������d ��]�of`#7}4jBiVu�lIyս�Y������G����ƛ�9�ng&A��a$���W��vfAը�Lzh��������YWf���U�b��HP ����k�k��b���w��$Y9ڴ��Y�fbo��vӖ�XI<_Ce�X�g��>�J�,�|	�י���7�bȞ�zdr��e��F���B������Q�*�Y��$�Sn1��"�H6���ׯ�0_N���k�8�̞���
ە���-��h%ݫ$�|��t���\au�"�[�y�b�mXU�ywY�:*.[Gv8�w����lc��&8�>�}���V��(��f�B�������Sn�0��|mݛ���u@M�sm1qև�B���bJ�W,@^S����+v��s2��
�����V�n�J�WX�K�����acO7q�x�X���*ՌQ,[o���^�'E��Ͳtŭ:��!�o/�[�A��7������֖BZ�e�yI��c'�vH�ܲ��������r�k��mc��[��um��~כe��=5AcP����,޵6)'Z�Hu��^����ۭ�.��6�x���Wg�p�YpV�jl����(���n��ڱ��\)��hُ���퇹JJjK�B��י�����7�Qʔ�:q\\5�L6�B�H6��4��E�{g�]�{i�؟2�zƱJ��S���e��q{졲�ڐŹ�l^e��x&�fHIB����	8̶F�A�U��8���Y��\����R�a���0c���U��#ECyN$�Wdi9���wu�����v7Q���\���p_Q�K���[ٕ�]�V�e�]�)\�����.�|�y��;�]م��]q��� +J�u�20�8 J��+��[puf��H�),�Sk)�oD@��ً�]tj
��8�4B1M��W6Y�7	�Z��;�{��21a��U��T�k*��o��e��%�poh�`]|+)gVr��9j�#�s���^��S��4��'q�ZM]iv	�����H �L�� ���h$f$�"-�mg8;�Y[m�Q�q rG%e��ۈ��������VwE!�9	�m���[���,��(�kM�"��+)��q96�)����s�yY�W�viqYM�K0����n�:��B�B ��,[�a�/nȤ�(���9$+��s�3mkm�dG%YM���:m�Q�Y�wOb����YŧY�mh���gt\ts�EE�vtY�n��fv�Ӓ[M���RfE�pY��QYv]6�clq���]��t���gV-���۷{5�m�uA�G%�GFw�ywG'Tq�qw��^� ��%GGRハ �x�w|���&p�C�Fۡ{qTs�G.c�Tl�Η��}�=�ͯ�7mǣq�{tp�5����oP'k�[P����zDͳ�j�+u�tOpD�f�3��Wg\s��<�m���:�6��q�A��S.�^��I�n:����윔�]�ۡ��=;{�e�tR!��5�Xtv�6x4��)��1���۸M��Ƶ�;��u��V�d�1O7Py{U��s�M�x{�-r���s��n���nٷF�E�x�v���\1��(9<lu�"\�9�lq۶���@Y��T�5Ŗ�x�ugK�mў3�&�嫷V�^l��b���:cy�!��󋃁�m
v�l��&����;;;��Pv��k��bB��M��n�$x���ɀݕ��٭����G�os���'nMGx��ݞ��cp�3��d�9@��H��X�H�nݼu��ݵ׀�NwR<Y�쇟`��G��!�[�V��7k�]s����Vݰ�f��:'\������TnƮ��3�mخɉ��C�f��6�sg�G��wdw������7`v�;P�67NLl���{c7\�ۇ/G3�i��Mvj�;�vsON�Bu{g�84�8��̻q[QnB��zn�z��u��,��$2��vyٺ�>Pz�pv��Í�ێݺqx�O��ly�s���Jv1�@x��{v�)\��^�^�;z m�n�Y���v�����v��jGu�yrj�;�6{9�"v�]Þ��M�ÖB8�*^֌p�r�b�nl�f�o3��G7*��˩�mƭ��u����Yó�yւ�9�
�a4�/�v^�wg���[z�������y���2*tn;88ۜ`45�1&�4y�wa�gY�ۓ��sm�	i79M��"O
Y#m�ua���7��������gT���ݩ���
۝ob�3��o\w㗱<-۩S-��q�^����Mס;�n�� ���=`sr�ٝ���q�!6��9jK�v���ˬ�mA����:tn��k��=�nS;�]��8�1� v�Ed����7:�Wk����JŽU�I�y��rcb�e3�u�n��vCc۶�f��6M��^Lp��g���m��s�Ÿ�j��l/S>.���<G;vSqγ��bz����*;%W��w!�\�b�n��l���<n�b�u6yx�.}��Лk��nv�htf�k�U�q�z��g�^.5g��[�<tWn;�%R�@�1��K"�D�����o�L ��|�z��m5�L(���:_)�Ӫ݀x(e�7���7�|�/�T�=;�hȾv	 []���H};�t>�ȷ<��jj�_$�����ß�����1�'��@B]=�ve!�ﺍonV�|mr�_F�_��j��b����T���.���s���<�ؖa'�z1œ�H|�hX�S��)�sy��b�aVۈ�r�XI�y3��ͱ�����lq�gA"6��AJ1ŀ(|+}�+���%�]�u:���
�6�&S��9�nζ������[����vWl�Ti�	��gWk���T�۞|�����gE�I!r��gZm��x�0H�;�O���Y+���_w��M�����Ѫy5Qŕ4Y�ˋ<@L��Z3��J�-�_-_�e���!u{�ǚ���w���e�7+ޢ��%[�(n1�/F����w.Ճ1�U+o�O�#��ԯ�	�v����®�
eVq>ަ�r�䌔,�1k��i��k۽����e�W���H]��hZ����R��SE�u�>'3,/���9>�E7vS��|I��Ȳ|I%u*�A#1�g$���;�}>�{���v*�+]*�]�W[J�
��so���������l�@!�v/ٝ}x���[t 0�EO����oj-˸*���0O��C��'��B�c�n�7;����ЮK�x��n*�*	;MaĂA��~�����tf�\t�U4�X'�oS���F��hT���K�1��P�]�����DAݮ��$��/:���mѝ����x	Yb3�x	����$�K��!B��Ɂ��7e�p_��2F��E(�lF��1�\���.�TYZ+w���+����Q=�V���Z-�����_�'9J��nlp�A��Y fu�a<���3#%*�ק��ϳ}9��k}�4��i����z��@����;#`
��!Sjh���a����,o͊ {N�To+�����d��{VH9�n�Ot�����O_�z�{XCwx,�h ����eۯ#�q����ݺ��(�K�^w.C�ft߿����TB�aQ7��e�-?��w;����}{ƣ�etT��)��������9P7�uIa&��3��i��3�[���}���$Z��^��@�b�͒,�[�2M	4(�����|���	;к,�2�S��qދ�ӏ)�J[k1�׽9�M�X��mP�++Mk��ܶ�r�푧;�^N�]	$����?d���I�ˍ�5}Z��34
&:��a�V`+0�ڞ�Cə.	@��5����®����S�śbK�Y�X<,>�Q�H�O����&n�C�Zr(JU���=��ww�[{�Hs�=Y���	���A��u��E�r�XZ��2W>�T����8�?ݭ�����J�0i(r�1�7m�����>��Y��'��˷��P�X��O��u`ֳ��nv�u��w��yB�ڮ�jT�Q��u�����zLѫϹWU�{�
��J�H*�v߳ٮ���9[m9Zn�,$׵3��M��^�M�֌}6��7���]O�.�b�t�H�fa8.�o�fZ��}��P�)�I ��ՂA9�قh�7���ּ�0OӓZ5�~V>�KQ"�Z��{��Ϟ����r�r�+�D�;��*��,	#uR��bǇt���"efd,Q����2�Sj �^�9;��'ڥS@�N#q_0���폻U?�����(��ɹqn� �q��<���:Ӂry����� ���]�s��0��جur��u��-B�=�wZ��@+�]��v뷹�a␷�n��YЎ��G98S�Ɗ�q��ln�q�>�XFy��{0�ǎݮ׋lu�Ү��SJ�����ݶ������ɝ���{:��Nݩ&�]�9���{[�ݧ�;�Ӑ6���l��3�Q�6ݮ�s]]&�aK�s�Wk��ڷ[m��۶�.;f�k������8PZZ�ʅq� �C�ud�Nv�f�*���&+g�,�H!�wgݡ!>��1>3UTl���a:�A�x󈀦a(�H$�T�� �f>��.ok��:� f�Gp]e�Ã2�+����~��b�y;��du�[�	�PD�>���J�ڥCUY\���Mk�ɭw�ϓm<�� �Fcy�	�8zj����Ǐ����t`�15�*�"�N�k��J�]F��(�U�da�˫ ��<�`��_<�繳{���1�����������qp��[�.�6�s��&���Ie����o˞	M	�2*���->�$Ƴ0�H$wJqg�-�������lP �%������N��v���h�M��:����R�D<s�)�wҶ�d��E���
^��D�ԭռvw$�YW��4��_�6���O���NaB̛*ʳ�(�{3	����Is�fꝋ=m
�9	�L�ĈU4EK�� �)9�G:V E�����?��3$��s�I�o�\�ʥ+�Q����d�����ǉ1�� �R�A(�"�&�oL{73R^�?s����l�T�j��I��+:li�w�Z�_rtu���<�@$wJ�I�+�0����n�����Z�^���w=���r��K]�+�pm�}sn�Fu��-���K�����[N���=��}�6�ޅ�dB��6Bu5��N�t�N7~���WIH�R+\�OO��ӕ��ɍ�fTe�}k�'�S��R�+�+R/���L֦H]D�����2j����u��8�+�My^�9�b�2J�
�⽯&oU�/�Ґӯӆ8/��SEP��`^Scu8��]�2L����!LBbf�@Ú��`�j��$�������BB}&�L���"��l��e�����LlUł|A�]N�9�zS�0�c�ⴠ=�p�r��4'0�����\����*uL�$��^ŒH#]:�q�fz$q.��۽۾�޴�K�;F5z5�;gq�=����=QB��$��2�J���	�͞]n��TZI7v8�|F�t,�����Ԟ��[��ߕK�i������FE~vЮL\�{z���]�f��]^Qf� nn*�~�m�#��yNEC+�v6.��R��Bzko���0��Q��~���Y$���w`�Fv�fyQ%�"�ȑ3QPst�D�&��Ro��>m�_�-Y�I>�t�����0,��b�RwC���B�o��� �u���=Ð����k���\EZd����U{'V��<D�[�>�ԁuQ�$�WFM=-w�}�Ep�E)(�n���6��s��lг���"�\������i��S��͎�GoN���]*C�"b�Ꞙ�,t�q�wY��ll�컙&t�:ӟ[�jۇ/����h2�J�R��&�5��i�9����S�aM-�wn�[�:wlX's~�,�ٲ�n��TZI4�ft�ms��u�6V^�L��<��IX�g�>����Sw�N�\J�|z�E8��>�Q�$̚�TD���y.X0��.�$����,����d�@�O3$��N,\s#�8���|o�w�|����f ��+�X$��[z��MW�^gf7���mWGTRR�'�hK�M�Nik��J	!�b� ���$��)X�����g�3�2pӝJ�!e1)P�mi�X����f��++Φf!�,�ʞw=�A�1�x�d�S����/1S.��j�,$�W�1a��B`M	�L&��v��3�]qtf�I\�{x�/V��u�ˁn�JJ=u�8�ק�W���Ͷ������r�{v���Ɏ�EՎע�u��s���g�!筸n����h��]=i���{5�'oma&Mln�\v�]&K����'8�S�9;3L���րO؜��-��qm��7:��u���13I������7	lܛ��z#gV *�m�vU�ns��k<[��ԭ6c�X�Ŗ2��w��:�d�RS���;��M�p�M?�}/:��Ȣ�ԗemze[�$�+��>���q��W���]o��o.>�x��u����,E+�FÚ���U94�ћ���6���cu�J�RK�gE�A'z)ܐI�,�u,K���CoӞ5�i�t��kצ�8���1�����n39U���P ��*���ɝ�`�^���>�FAO& ԙ2(UƵ ��Y���B��f�>u5q~ ��+�A';;3^�7o��N���#E���DҲ���J���ۈ�\�bϰuZt��H��J�D����j Lqs�_"�
 h��X� Ky�'�V���7�@P��c�M���,�^�8�t�n��}����`�h]H�w�8Z;G��.ѤP�dz<0���`o���y��$EW��'Y���Q�VAWp0���S��6�QWO�'��@���٘	����
�^\#����*b���V:"�D�J�ٞ�F=�z�Ƣfz:���A��|}�ݙ�lP�h��(L�LM����fSo���O\V܂-� ;�x���� =Yb
Lƾ�3�L���(U19�$��<l#�GZ;�;
�� �����*f�SL�qg�=MHr�*�v�C���<E���Ѹݺ�S�E�t="+C�m6Z���.����rdP�'��J䑯Vf�Gr�o�T��~�=8��1�$��3<O�P.B���_z��ڙE��x���U������ �T̀I��n���&�qj��cx�H(ZE�+ۭ�6���פ�M��L/f[�<i�؆H�����~�:�^X�W��/�Z��h�z�jW�Du��
9��AKp�!R�N��Ԯ�U���}:7�;([�{ϵ���x�}0�[-��J�9\��&�ݘ����F�J��%7���7.�pT64O�h�%���x'd�f����T�4��Os{"\�y� >��[\:�7,.X�m��V��QZ��w*�@���8y�o];r�H;c�[9��� �w]e���"���\�9zȍ`�Y�+,����ӕձ�e3ha�sQ�!����h�WD�sT3�L�N[���^vݬ�3t�'��D�h�ã��ޚ���^��UQ(���QKM�S���-���H���ssR��YƬg*��By^њ����p�{9n����݂�7�4VӖ��dxK����/�:8�#[�5�DiL���3��4��e�f��u��V6���'ץm�/�`T��2,�"3E�(Xq�`sV�D9��]���s͵�՗��C�y/o$؎��oL͂Q=]���JW�e^��N��O�0���'����j��M��v=�3"�D<�X%�B�b�3�6��ò0�d��H�����5>p�B8�Ks�Z��I����Φ��@|�p�`�f�%�v`����qi�r�]'rE����������is�̺��.�h��j�Y��̷o�\���,����+:�+��;�.��vz(ee��'�xo��T�]��.����K��偃��6�F���ݮ�tN��[��'Gf��;��3�V��ئa��� �����/����\e�H$�\^X�Oh��fe�DV]yޝE)�PA^wg�9��)ʎ���g��;��K��gq�I�w9I���8	;�(㊎��6�q�ggT�gQ�yv�yXtrr%I�w6m^]�t���eD�Zy�u�Vsb���mm���뽫E�Y�{b"������*���Iv]��qu�]�\ǑubQwq��s��A�f���:s��)"��ʳ�n����K��B+����[k�ȯ���;���X�]y�q�Snθ�\�(��DE �B�).�����cy���k�sX�'�ru�mx�d��qZ�.��N<}���Āk�m�'Ò�E�t�)W�棭oҟ�ڝ��F��&����L�ڬ�6	�=N�]An�8a�r~�����S7�A'OR��Z�
��G�!ٓm'e0nT���,�{<�O=q���J��4��=ë�;�V�ɵ�Ox` �)�~$O�:��K��]���l >���PYҁˡ����zr�P����aW�=���P7����mҡ�Qp�)yط�f��m3��r�]!-o^ק��M7׻�%[lua�¬�oo` ���E�H:z�������j
Y��?ff�,;^���߀��P P�mҠ:{[�ط^�K�mk�r��ϟ�x,C׼��o���\�o&�:Qn'a6��s�	�u
�*��
E�CM��n�B=pj��������{���;9�I��/�l�Ў+]�O�o,Q� ����j�AȪ�S�
����/�#��k�Bʣb<@����p#q��S��.�0!���:�;G=�Qoϯ��߉�)T�޳6-5���*�m7��ُ��j���{��T �r�]ȺydXϲ��n��N�(J[v�b�{�;��$�O�9�����A�Pڑ1=(�<�~t�A؝�(UczN�o��W�^ĳN9�Lɮ|+�I *���&��fx�t�Y��&��TN`����n�U������+��|A�f`#�1�N�������zI��$4b�0&�ᙙG�I�1�=��T�2�� :�l�H�י��qŃ{��x;��E�IDmP�l��h�C���a��c���`_>]�.^<�z�C�j�o'��X.�)z^ق�UӜ�����;��s������q�;����Q��q�/V� q��I�l���.qj�v���6�rmڼ۸� ٷH�3�y���0#;�d�� c��S���>K��=�]1Dw逺<s�ڸ5�Vm�a��ձ]ՠy�m�=7xꈞ�jcq�xk��w�nS��F8�*t���E]=�3v7e�:n����#)v:�4\��Q�ɵpzq�u�#�sA�۟FZ����%��ؠNPlC���ع��Eb�AFӒ�^�t�RB�����_�
S���� �[�\:|�-I�Y�]v(/_f`'�v(`5JU�^�:k��s|S����y9DIƲ��&�y���N������vd��xc��U~ތYb��U+�����5�О3����*�<f�� �y�@^��E���dr�k�Xڏ��u����|i����uŒ	,�"1��/b�)��9��G�t�iUU�K[�קp�$�;J�k�M
��{����z��H����_�!���d���me�2X}'ڻҢn{X����=�nA�������C+3��j5�{���E�
Y���9���6�~ᾟi����~;c{.��#';s	�#����#�8�M]�',�1��z�HC׵ۊ�R�ز�}�}��F�� ����70�����^
�޽��[d��]oL�Z����Ŋ�B��jb]En�|It��b�$�)Œ|���`��U����\��/k��AR�B�=�3��O���A&���r��ٷ�'��t�H$���<�0dQ���	�&'0�\�0����ʉ ���X$��ʺ�N=�ͮ��Kښ]E��_6�]uX�nX8Ucz����=5�vq+�>�T���� ������>�mr�b�P�z�:M�7i�W<f��Q�!o2cR��t�kqs(;n�߹�~��cRT��vw|�h���� ����Q��Z'U����	$Ν�=�+��5>5UV�f�qzB4io�o��q�T  C3����g� ŋu1���qv��0H�X^��,c��}���lP|t���e����(�-��Y�l�e�meE(F�W*�V{7f#��A��:V-XI�
.�G9՜�o)�2�UݗR.%�-|}M���{����{٘�]͕b�,j�IH�^�|W[�ȥ=@��*�(S{���޽��%g�,��)�Ek�Ⱥg,ɡD�19��,�|�.�)opmB�nS�@�<۠(
��x��q���o��~�#jF�6Il	l+�ӆ��]nV�n-���s�����Ud�
4�;��z�
9Sb�I<h��D�w��H'�S����5.�p�s�;�0���H2*H��r�:���8�_U�-�Y	I
��x�fI�8�L����h$yҭa���5>3UB��w#�Nl�yeμR���Y�����Vwfg���͂���K�IQ�c���k9��\�^`V^<H*�,�*�n�З� �ZN�]XH�]��M���.\4sI����j�dl�1�f>ϕ���Y��Y�Ǹ+�8���r�����n�:/6�f{1���*�PQ�FJ3�o�I����[���H�3�Ud������'�3ԬVeU��Č��Ǫ7o;d;���w[b3wD��!6<sX��X֦�2Is8yt)~r��՛�w�O���d�|	qԦ�r宪̧��-t�P��5�`�`���ʰP���<vҞ���/F	�'�9t�$�z�� �	��e����'�"h�"������6}�iX�	�"��B|�$�ᮛ�R�z��BLɚ �UX7ٚ���h\6nk�L�͂A$��iȰO���3�'1s�(�d�wGE��&(�jj3��D���eW`��g�&�ҹ͂,��c���o�p�q;7:�1k3
:oQ=�T��ʺ.�S�F��J\�i�,�Y��#��^�sA�F�*���9�l�@�vw����zz�K�q�=D�֓u6ݜoZ�r��l�;<�
�[с�4�m\qס�3�����[l(���m��t;{�q�ۦ3���VŴq��)�m���l��Ƒέ��ZZ���v�:�{mss�� ��m4k[�Ǝ���{R�k�:�l�m#Ov�sQҘ�O�WG<�3��'t�������������5�]Y˸�dMZz(��uǱ��o4��78��Ɨ�GU\�M���Z��w����Q`*�%|Vt� ��S�`�۽��i��f��y�\�f�=�i����W����/�Q����c��:�nx�)~$��ӛ$۽�����H���S]�)�NN ��m�0�������~�k�maq,�/��N4�{~��M���l�-�j	(A��r�u����X2�tp�+,�uq�wD�޼�'Ď�Nq8{�뙨���O��_����ݍ9�.e_%%1B�7z��Qy��3�(l�i�<=�hG�}ɫ���,��ʲያ֢� �gI��Wt��F�"�U;ok��m��F81Fd��I��|t����%.Y��������1˺A�yC��[t;!�E����f��s�I��;�r4���՚�){�1&��ba9�9L8�Y"i��d�[�R�0]^��cuY#o՘^v2�`玶�P"�"a8�)I�.٪��O��f`#�'"�R��bg�)L��l�饦!�~r�ɭ�o����O�T �\�+��ܶ sۚ��~�Κ��G18K ��Ǥ���F���,IQ����e�#T�� �=HܽW{T�k��c��a"8���A"V�J�e��=|�>��Iv��m�o�M�|*�^aj��>#OR�U�!�V\o��-if��V�l��Q�\�(R��y�Tq�%OE{y�Z�7�'I�r�k����k�U��x�` ���� �v:��8��4�:C9��$��q�{z"įT�4I55�8$�sV'Y��$�Z����Ru3~$�t�)�6���Hv����Zf���u���٫צ�Oo׺�7��^��A̋%�R��ܹt	X#Y�|%��_��<qM�d�;�Z�&*A�fG���kQ��zB���:�#�U���X�u�$�w���@'�OR�Ds��"=SPA�2bs�k�TUص[2+"�g�����"��>Y���qq:{�[J{��oڜ�Z���~4^��|w���#.�8)\���2�l�|�R��ܳ0�8]��jNRI�3�m��'l�������5��������!�K]	�'�y��A	Q�^z���?�\�X ����;����	��3� |/5�k�S�l/Ď��;�f�o���T���j�>�Qdgr��b�z��	�;�>��V7�4.�ᗅ��Vߤ�J\�0�	C����ֽYҮ�K���}M�}��I��ʝE����e�e����Z��,�|߉50�� ��Y� ���(�\;
�t��T�&�#%%4^��e1b�mz��<qoV?,�=dU+
�;{y���O�*���\�u���2V�"������6N;]�������ķ��Hi/A�z��&oLRk�(ɉ����	'O.�%���3PM�Ӂd�\�z99�c0վsڼ�ܜ�K]�X�(�*��2E��n6,qZ��B��TeH�i�V�P�|ﺣ%VADTh��%`I#ZYxI���Vnr���+���5���t���B�dM����L�+躙���KMfa>%��	=��ܡB�a�J�:~���<�'>7c.���9' P��� �/��Z�rۉ���axO�yf`'ľ�qK�Ovw�4.�ᗅ�����Oy�m�
��́S�x�>�9�w)�7��Gؽ�wy���+u;�Q*�m�7���cf��Z"Ύ�t� �F8�V;�c��@�$��H@��H@����$�B���$ I?�B���IO�H@��B���IO��$ I?�B��B��IM@� �HHB�	!I��IO�H@�`$�	'�H@�HB��IO�b��L����¾�n� � ���{ϻ ����;�      �        @   r�
$
 (P% H(P�P�
 (P�Ig��"������	R	JR�(J��(**�@ �(-�T%@����Y�IV�N��v{�Wq�;�[���r�ؓM.{�.�wp��qR_|DH.7�/���Ux罸��i��ܳ��%g�ON����4�ۭ2��D%�)HJ󆆽���;�&��\<Y�m����W>�������{�>��wf�=��@����z	���<.נ�Õ��u�_+���������h�c��3�
Q!�� �**U(�EP�S��4�k�-��C@���=�g/v������8��i����]аWж��xR��T��)("�
Px(=��@P}3�s����4ժݍQ��ܕ�4ٞ
���=��}����򧸦����:{jfw�^�]��:�Ӫ-j�UU_>*U}�R)A*(Q����4iY�⻨v�Pwn�݀Q�L�8=���W ��U���������O*wZ���WwyQ�V���^w7m�Z��(    ���4�)M `�4 &�4h`F��4ԥR��      S̪F)%A�44���@ j~)R���   h �@ T�D���U=@       I�5 �42M4�F��=G����56ԟw�� O�Z}��ow���4��� I�Nu��|�I=����&IBC�!I�?�I �a#}�����?�O�`r��Ќ`M���%C�����	$��2"��	 �M���������������o@I8��㩭��jr�>����YJ"���=���|��vv�\7Ỳ�����ӳ���v@gG��J���4��O-%�ܓa"�0��Ox�n��%v�1�58S�ZS�+Nka�J��2�-6�1^b#�w9G�nJ�8%X�,/WasK�f�NL�/(]hb��ǝYؓ��{-���oX�$f�ͬ��Σ��'r>��܈􊧆t����ȗ�wK�㉮��� :�ю+��vmq��(pVv�&Vn�t]#^	+�p��ǠP+�����U�$��hdn�%�ۮȺ�8T�+A�p�xޝX��M@K��:�ܾ��}�Fk��Aj>��np;�.�z�ı�1��A�t�_ �#�ػy��,;�ٹ�&��_o-�d����lS���n��9۷d�p�ݹm��Čjp�gEkU>F`��T=������،�X�����]s�p��sl;.O�`��)�C/li�ht+o�=8v�TA;D���ò��Ȣި�������pЋ�;D�F�� ��7���kc���	�=��8�l\�b�0��9 �W1q3Y�wq�gZ�g^s�֞����!f��"Ž��~�np<X�^�	���
��z��(��:V %v��x�\�5�����+��kg1ΰgc��X���M�S5*���&�=grݸb��<,�/5䳂��^�7��'�b�΃S�Ӯ��#k�Lq�1�r�h�t�ނ��so4݆c㫏*�`:SGeY�yd(�7�jLλf�m��z��E��6��ۣl�^G��	M��GC|�MΈvuHY�Ҩ����oaܓ.Ny��g��G;tB�AB{��%�C�������/���=З.��ǋ�]�m�+~[p�r;�����������N�ˏ]�8�ڭ���	�D��ZB߈ ��5M�B����nw�{u�7Y�:�:!�s�hoQ�[�*;�*s{��("Kr�!��9�� ���3�hU+�h���M����5;�.P�6f�K�Ƿ@;�ٯ�� ��Q{�|�$�$�rq���ըU&��I�u*ŗW�!&]��ţz�޷WSy�g��єb�i�V	�;�4���I��8+��&�Ԕ�FnȾsi�e�E�I���ٓ�z;{ई]�����C�I�F� v����؉�Oe��W3��E�Q�v܅���J,\���݃H����VqV4�GZ	��V}��<����n�5amX2r�G�B�}	���Tꡒ��U���z���&D��֢п9н��;YH;�9�Qڰ�d�w7	H�6e<�x"�;N]����w>��i�^Lo  v��f���v�0g3Fi�9��\/����a������ĕ��cׂ�v�bC9+S����wV���֖�9�<��4n��;��퇉5��]}F.�l��Oc�������s!JgnE����
����L�&�(���+bngGo���"��M�Ԟ��%i����G�x��`=\{jJJ�5V�v��{/vu�5����('t��1 �D�x�Q{n��0�Zw�����+����b8�U�6bB�*�wn1�8��t' �X	Zmu�;���'��\��ߡ=Ż��:�Dx��7`ݎ�ptAd��O,;��D�I:zn�R&�(��IN��X�G����sZ�}0�/cx��c��.�#v�,f�Q��/A�'`_vʈ�IM�투�tr#���������@\
���ҋ�oi�F�Ls:X��Át'E����!��\���s�m�*o�rk����(���pT�,��o�����7b��W��;i�SsA݃���s��Q`)Q!��Y�rkmX:ٚ���c�8��ESk�B��41U�UB���f����[Xn]|G ��\��h�D��n��;v
�P��L��Դ�L?���v��
��W�8\xSO���a��ɻ��8oO;6cї����P�C
�m��;\2��F�!ac1j�r�<}T�O#NՂܐm�>])x�z��ED�I>�HR�4��#�����St\��Z��pY�S��d�
O�+�_0x]C��Y-�/t^���n�g-�����W?��l��P��Fwk+n���G�I@����
���w�K�oh������\�;.�Ө�m`%�#�|Tq].�P�Q�rGӵ�I�^���=�;.�	�{`Z'rg:gP#qp��s�˷�s�X3�W�s"Cu�w�;��F���*9>oF��b������/��{��|C�5�1�O6���t�ۻ��f���i'��SuWKZ-_i!�N7��qV<�{��wH�:z�5Y�5���x	���7���}7�EاQ�T����4Q����.�^�Ł	9�K{76сn��E�e����rX1Zx��z]YcYE{�Y�p]sGD�i�0�4#O:��� ���9��7�W��仂�]�}�P���1Q������ԍ�l���\*y|w5�T�N��ءK���2�w �U��{��'��	-;���w���cOL�����Qw$�2P�[N�R�d[����u<���;�\�ڥ,�,m��_#�ڌŸ�^�ďc��i��q�To-���⢘ ��7$��� ���E� <(��h�\�	ju����[sm��w.3�\g
ѽ7L��	��n�u��t.k�m�>�P�g��7��qTG�7�N�V���k��m\|�,��q�d�ތ"� �>2���9����:M<z��P	�d艸��y�N|�o>ji
�Ŝ��Ϸh��O��F,\�j��K�Y��e.�Ϩ��w�a�p|���䣰�vv�<�+ފJ��z�2�}T�fO��7� �ko�OR���0�;�c�S���+w��w�"{5iR�z�(g7j�c#��wO>Bp�*����޻�[QH�`\�gp�K���tb��@`���צU����C�r���"��Q[������ڃ)��^���mꋶ��1�/[9����e�M=!��4V�Ĝ��!��� ��(����n93W_���W�ܐ��3����q�[b.�V�/�!�;t����N��#nI�w�����d�s�US��e����V�E|�yqb!�;�*��r�eHP�c.VtA�ޱ��)�LW�>WwFD:����P��{)z!�zwvN��.�N�qr�	%Y��c��,�{��w�"rnw1�^L#!\���y����Z�����PF F��'�:�[E�Dӓrm<���\]ӫyHŝ�;�nM�B��N��� %�M|Z|N�_B���d�(�N��>]rn�".w��N��p��Ȿ3���$����b��7�&��[¹,{(�hݣ�K#�.��jR-�qg�]�!����?�������\?��NSq"S��H姷�h�Ǩh	s a!�� VI �  �!+	%BAa"� (@RI+� �d�P� P�(B,Y!"�BTH �!`@�@P!��$"�$
��*@�� J�E�)H�
H,$P�!*BI+	 ,�H,�YI	,�("�
"����%`R@%Bd		>�g��|�;��>�h�|?p I#���IBI<�mB�C�����I�?P�M��>'��=�p�����݉)�g��z��K��˄_Q4.�����ѹ.��v��XzY��@�/�"M��ª�b�
�{S�ܫ~u�S������BH^�+��Jr�[�*]J��L�JC0n�9�H�n�]�۷H���
��u�;�h��=9�9$�`���`�\���f�V��D��|�G�ԿqK�{{�~ݻ.S�*�-
���Ve�d��;L�B��f%��Ս=����������`�f��b��s�vjqE:�y��I�y"6]ί����o��a^d�'�R����g����@��/i�$|���|�b��2j�ȹ
K�X�^*j��jdE��ҫx@���=��FW���;3^-��:"��b���~26�5��)v>���j3a�[BCAb�X�7�����Y�q3�;���� �MB׾r�R�L��>�$��.�<��2�,�,��5��3�U�}���p,�� �D ���ȡ�òD
J޸�y��	lgM�Oc�������)��s>��,xh�i4�<���t՛k������1*ʘ0�V^�_0X}���P�s\��=����7�k�}�Rٿ{D�-����2�w���i�ݎ�|4��_��>����F�FζY���mF`4�Q>X����_��#� �
�	;����zT� ��z�}��P7�V�W�}Ӽ;	��^;�շ�-[R7AH7b\���k'*�͇�/D\�QrЩu��̗ie:�5�;�ٻ���C�ܺ�y�w�7��w�H�g�ݠ�pM��y=e^�VK��|Ƿ��\Ƚ�;�Á
^�ya������������|I)c�Xa"u)��%Zw|d�z������Rq<➒HŊ[~�\&���Y�qB�H4����1��)�wcJ�0o��=�a�E�Oi���1�������Q�vz�N@�h�Aj���NS�Qr\�p-�=�q�*��wg��y��
�r�m�R���*�i�ȁ�0�4�qW��.2m���">��s�='ܑ�Ҵ7����Cy�}��H��\BGɠ+��]�}b�{��wW���II��
�d���jXL~�����j�,�A�����j^�(�Nb��A �w����O��;i��3��*?4�'qGP營��f��=��z�|�&����ý��9�aV�U(���#&���2-�I��Q[�Vyn��3��9I�R�7�\���q+7�[���&E�����7��	>"}��P�\�P���f^�Ff��rj�Onvw�I���A\p6T11Q*��,[*����LUT�7��N���=�t�)��\�d1^fp���1��{A��ww��}��g{q��<��x����g6`0�HN�%�>�uY]���B�^q��}j��rp&1�k��Iٚ�5P�+vT�j�6���$i/|*{���j��f��~&K�%L��*{sg}ܷ���w��UG�-b��q�F��I���kޖM?]z{���~�ڦ��l�{s�n������W����m�9}��yos�}�拸�����|�_���4��#D�AH�4� -�Rw&]֭�b
�%�)U��sR�\�4rΧSmʹ"����q7���(vy���RG�=b�YJ�n�@���ܗ��x�El�2��;͌TH�qf�V�hn���t�=�:�}��燝�/v?���rd�����o��}��3���L�r��c�wo3\vz���%k_�%����}�7�v�{�uM�4�����>�a�;v}c5�h�C��[�������7�u�c����&r�l���m��[�2�#.E�7fXa5�J�rV=w6o,�f$�F	�&���t$C�5�����5�;o=�l{�7�ݜ{�9ޜ,�_�˴g���v��vt�ܟ�6;����z��?�ΙǼ��j�
�y �A�$d�2��k����j}޹�=�bXni���hKl��i7۞nd�5���L[��س|��c�����*�؏[�������M���g�ص�������=��ė�8�w3��ܾf��=0����i�j]��G�X����:�����(5�B�'�4�j)����[�����V5��}�V����M�q��'e �x)	�*C��~%m�8)�wۋ%=�^z�;	g:�OOc��ou�㫺0�nE��O���wh�5�CL�QE�c]hOv�2��Y7qg,H�/�����tN��O��n��S7��AD%n�	���F�˸�ՃVNQf�z"��n����Y�j��?k
��+讀��߽μ~[���;��^�ӧWM:U0�<�\���2&es�����4�����Nb�L��)�c��&���i;�lM��b[?o��\4�㽌�}	>�W�Z��\�'�~x�R��]��F��Y�/h�q�����ϴ���#+p][�6�xvsod��{�p�(��Wӟm	�w%U0��7Oq����Ќ=uYp�޿u�_H����7/�����Nr�2��b׹㸅�6޺���|l>˛�U������Y-�zp��Ȃ�g���_p�{	�r��i���������l	��=�����J��9q� ��.�i.->�r��or|"�<���k�Ü$�bӕ�W�C�5=��eg��������B�Ɨ�m֡WI�q(E�~���
�䧧�7�;�:u9���/u�'u�{��)�|��r�w�d���j�����2�v��w�ۆo�WW�����p&%�n�R��E�7�n_�VK��<�7e�F��Ͱ�-�bV�K�O|����[{�����{���r��І�<�d[��Ox����9�7f,���������=|�]�v^Ow���bb�i�8���{5	ڐ����]�;��	}�?�p�ǌƏ�L��Ga�u��(ʇ2�����4s�d7�<K�������x�`&���}�P՛����s��'�6���/�5r�ȿ2S�;�;�s����)��Q���;|��=��;���L�v/ ��4��Z����|I��MZ:�˭inUe����ܩ��Q���z�N�=�ù� ���uym�"��%+�h����f�tͧ;��|�?M��$a�$�;�:�tzik"#�b}���8��͵wi��2XA<�>�zJ(���֯5�_>���v>�C�{�=�i�P�'�S��~m�T����tG�}�MMw���Fx��^u�|���鷓Зm�F��|��}wX �����.]ө�ڜP]\Nܰ�Xrn�=�gL��E�g>=*8�Ŵ7F��2�T�q�#�W/{�0�*���G7K��Y������潂 �u`�P�ެ���@cݣ�u��S�	�#W�ꢼ�ົoh6���I�ٷ���<�{�L^^;�m��{�������b��L[���	K��E�4�錺��A(���`���QI7�*�-�M{
��/]Uڴ�.?�d��p�/($u����.\���-�z�����t��u�.��aJ�����f���;�n�m�^�� H�,�@���������F��n�Z�p˦�ґY����fJ��m�Ɩ�l�hFl�E\�l،]�ԆA+�ax�T�`��*g����<�����L�nf��b�e�%�Vn�Q��.
d����d뀎�� n�>���r�-��,�ql�Um��H����[F�)���Y�¥3��ƻ��󞎷u�n��(ػ��w���V�xx�S��pZK�Rͳ���1��%�.Pݹ���g�!����Oa΅ДIK/3s�$��-n�,3���٦�-n�i�".D��\%�V4�I�6�:��m�	cF��cM�$]��k�qZ��-�ű���)KMv��#q�GӒ�>fk��ny7�۹�.<��rZ*ŗ]�ڰtr��j�lɔ��cX���i����)`4�ux����أJ܊��\�(�R����l�����[Vm˂g�k�م��y�A�.J͍Y���̵���V�a�[��-��ħ$2��Y`٢�5��X-�;�,u��tJA�,W�+���dY�:�4�Z��M.	�p���<c�s�\krI��n���U"g��
2�du�X�VX�^WJ�<��YM��^�X�	M�k-d훬��Qp��iN��X�z^u�Җ�F��*��\�lD�� 9��cL�ь'���@K�<���twf�d�xO 9|�r;��$L�Nŭ�c4u�l�mQ�F���m���ŵ���2�v�ۊ�B�!t���ffSdͲ��Q�\j���U����<�d�6�6�(#.��$<�Y�F:B�X,�;��h�j�y�rF�p�0��"f30�K�f�bb-���nYm&v�kk���3I�f���Ҥv�&�%�կqk�u��½��N��y��n�al�R�]B��-�J�%�n��խ��h3!P�=��9�s�,�֬+��*YJ�FZ<�hl�V��%�y�Ӝ<E�ݹ����ٲ��"���Q5&��ah3
���lFme <iH
1�P�e4���L,�9�]f��Z���:�8�:�����-ew6���F�<�ճi�^���E��2n��vy����J��ss˖V'��KH��x)���%f[0��X{��-2��\�:;%�-�Z���Ť�G38l���F��h���_&熞pt��YR�e=Ѹ�
��V���8�w�5	%��.z�w]�x�u=i��\�.Cփ�T�hLW�͕�*����\k����̨����2�9�n,�k��.�!v��&�x�����ҽ�zZ�|v�����׉�9y��f*9�c5�*Rۛ7�YR�(�֚�4_';������O�G��t!��
Dkf�h���L�E�s�)61�V!�6�KŜ��q�J�՛���G3�1�A�Z[�Ё�+�G�,Kll�XG[0���؎E�P�p�E��z��HR.b
���mll�뵼c�*�h�rg��qkfZ��Vי�j�B��	t@�#�(���5����s�æ���t�6��qytqʈ�[b�;��:�i�K�@Ņ�ZV%�[��h &<�e��]���G]�܁�V�l�`�E��j��Llp6�J�[�s�^ ༶٬��(��!�Y�^��l�ue�3-�$%����C�{���^�
zw/g��^z�<>��������[�����k�n*Y���R�6퓋h�"�<�[��+֨妹BۊL츍�sF�c�� ����6���9�iFfQ�c��:�p�-�u��b���m��w&h}r��{�ӯ��%n�y�w&�{`��nn.��&7qm.�z�ѳ�"�]Z�ݬ`Ɩ�֢�h���KB�K��L��ɞ(ů-�Ɨ(�ɀ��u������:�R���̫)�t�3�0CK@�,�hDP���]���ғ&�u��i
�E]�1�D�ҩȋ�<$���0�=�ѓSQҡTC�"X<�٥leu�b�j(�B�b&��r��:k�c�xB����mk�3EƎ�Q����je��.��.�n-�b�`w
F�mvbLgsJ�64�Z���ͩ�鮶�Ü7S��-��k��p�X��A���\b8_/hR�m]�ڽ��Ff�Ck�
���\YZ5�s2�kWL�]����IL�]�MN�3�y�L/{�]�fH�[�ř�9F�cX$��n�n�4c:����3\>3g�&<wa�N^*:j�k�q�Qwn��u2�s���j��)ƅs	]��5�u�z#A�N��v�/�<Q�(k��4eZٷ�E��r�,�04O]8�sݣ��0�j�Տ^��<>g#g��c��t�c4� �{qۛttc��f-f��g"4[e���%e�[*͚50��s��Tg�f�l�u�C��vfAb�:ˁ*�.���5�+����F��d�+�TUUUUQv�eWl*�Q�L�j�DU�ю�.ڵ,#X0Z��J���͚�F&�Ͷ#�kH�Hlc26�6�2��Kv�#�K	r�dn��4rk5B��c�]Arm*���ˌa���c���4[X�m�,A�����Eâ�e��hM6��g)6��s��\���2��Ҁ��K��9N0�"֩3A�]��o?;�ug?Z�B��m��F�d�-��V��P���GL+P�������H*!RUf0��`���KmEmk�\`�7�ڲN���ن=�&'d���6W�M�pG���XQ��
�����(��v5W��!=�l �ċ�D{&W+�S������M�p���6Lϓ�6�� ɲ�����`W�=��p$d �7�%�&�/�����Mj�0D�u �n��nk#�lб6qt�����r{֬`+/�۱�p���8(u9ݧ����d�mE]c@tM�&Z�x�H0�<\����t/ ���n�]�u�몸\4��B���k�}�;Ӝ�0]��%��%�%���d�g6(b|4�'���]��%2��L���\���6]�2\�5��7ͫk�ۓd�5 ��X�jhM��iLF[)�p�+�l)<v�;���rr�5�py��]a�B=%��B�{w:��U�]-e���nc��
�(����2��ӻ�wZ�6*��C��Y�nŘ �\�X�s(��,Na��o��Ь+-5u���U]uѳ)�\BaH�֕�6Y,�st-��*,��Y�r�T���Që��W#�̍e��x����oG�q1�sg\ܤֱ�!�d�ڵ�i������ص�k�Y���Һ$)��m�ڨVٮ��*�"mT��jڥ͖&�X�Z����m�+(W���+���s�{m�n�u�F�,��,i.���V��TW���k8��>����L�ưz���o> �l�`�_6�ӯM��eĥbe-��BV�-�9�I�������
���޸}Ɵ�6)'���w�F�S�Wq�IL�Z���(���2b�x�I�AmKΙ�Y��[44�ĳ� ��0�eL��1��>��&l:���m���Q��.�P���tT.��0G�z��D�dP\�P%:Mc�v��%���߉��j�br��f�Ս�X9*�+޵�h$�f���o�*������L�F�4a�>M�������2sU�=}tɑ^���T� Z�������}��8/��� �j%�"�۸����聄u%�z�2<B'�IOt]�I�����W�*v�x�g�HF<Rl��f9�.��b"3a�"E���(OF��	7�/�)#�~�����{��:���*� �As�!mW�{���(u���׀A �� c�\�@�An.�i�)V�(�С�S��A�k�!���f�ι�$���$��6Q*��J����ۧ��8�A��L]P��DP6uu`�:(�[Y@�7��3n"UƉ��f���Oyn���J�3Wc�2E��h+G#������O��N���O�x�tp��c
�*͢3\s�����I_�ν,����摣��n� ��P$ZV҉�Rq`��eV3�*�t��������cCV�)P���]�@�蠩4'�Α .�Q��:�G��M��ެ(�A�@=�=p�����c�W.p�=Y��h��w����`�=��<!�Ũ;�x�IL�cxq�*��t:�g$B�S�/{}'`�ۤ5�O!�Gu�+=�3�w7go�.,�3�Ƃ�1w�*�b��V�5M/Q\[Ƭ��7���iT�Z���^o�#�D�d���,�p�:H'�"H�@#�CS�R�=V��	�> ��"8��R�n�ޏ��%�����|��>�<��%܊Q�vb��N�@6r�U�
rM}�����}#IwOjq8�X����<��'Y��s�yi@�.�E��m�����^,�����tع8�ϙ���Ɗ�+4f������n֕6��x�܁��U1ݎC�V��9J�x��J[0�F�p�m�l0����K6�l5Z�^}�y����oo�[g��,_L�C���)BTYE����v���ǂ��9/�OK��4��"�Ӟ�F(~�PWơe�[�H��Q� Z� `@`�𝏜o���Rw�r���^���s=	�r��"�t#��fqR�g�����Ŷ��8J�-T��l��o��%�� ,�L��#��P�B�1���(����x�FR�~�?@�?���Bk�K��b~��� }"q�g|Ԛ����4b�@��{fIإ��[H���:s@l=d hD^�\�P3v]���h�N�>�o�=\_1�&jV$[����O�(W;���e;!A�ALLX���Q�P�Zj�E���lR9��0�3͈�$�|Q�N �$KZt�"�Ha��d���#��8�>���.�G�.�4�:
��[��]<����>G�b�H�Vj���ϟ@��U������7w���~��;�a���=��7�C�˱�����Jf�w~=}{B�L޸\��N0Bj�[���;�:�]Od>�����׷˼�z,���4c�6٦9)l�7-U����0�t�l����wd��;��� ��r#:I�bdJ[w�\��q��[��o���2Q��� a�$p�QW",U�[�:erߡo��݃mQ�k��p\(�@�t�8g:�'d�;�h�;<n�9�bwGU������:��m�7�}+��:q������,�*�� j6)I�j]��7J�������w�į���� 8a z'��r_|b+����M��#�i�u���I�o� ���>�k��n`�	7eQ �@@�E��d`�+�8���J��`;\�Av�{=J�B��#�Wz�ϡ���Xh��n�J(��8�F�M�Nհ<�9����7�D��A�'^zE���y������q#���`���'q��\^/R�4�CWM�
,ǆG(]�iV�xw@�/&�{�u��X	c�km��+V0��en��>9���y�������ZA{�wI=鎮$l�w��se�f�K(A-��+-ɮ�I��0�/���P#6=<��,��8Z�^A�W:{�t����c 9��=�>��Rf�y�IA.�@\���3�d!�E��+��$Dݔ_\������rځ��j��_��Af!�������G}91:	�@m�߀�hA��e�B�e���$inh�5lq��{���ίz�@9 �+zC�i�Y�@9�L�t��	1b	�p�	%ԚL�]gs���3Z��T.�DZ�n�ᨕ�g��$8��}W�G���0������ ���n����{^��%���BB��1�g���|>��(�9�`��GO��U'\�������3s,�j ����y�����m�4�
�8��|���߷a���lf�d"]�;X0��@Q�!7����]��]{n��ע��H��R��K��*��'>0��Ơ�?������	J
���o�r�lU�WkԎ(?����,Άt�V�-�V\9�j����!��|+$���{H�]�;'gQܰba5�n��s�~�Q��.{7(��ޯKjO֮3��ˌ\l�u"d�$�CV��:���W�S�BS6�+�cz��W)��o+���ڜsw{:{V~o8"a�A����%u7Y	BV����y��4�������98���<�}�ߣ�z5�5w���}��ޮ;�t�����圪����2��Saž{�̷=�7�,�%k��vc׀�EȻW{�nS�gj�leN׮ҕ(���^��6��x���6?�,\�ؽ#z�5n<`�!5s`[ވsO�J��u��<h���W��6	<��7فڅ�m�z��aŷ<9�m��4Ŋ, l<�yP��%�����&pO�|�_>809�6&=��7�h�c�,x5m*�ʲ�R��R��P�ŋ��k��ؤ�*
��6�b�J�:L�J����\C��-X��t�X����t��uxSk+�H���u����Fе�F*��eGN�)&SZ��-��LTD�aT�V[֍X�Z�g"y�ő��p{
��d� �� !�s��0Ns�q���f2�=�g9o�˃���pt�wNr��M��o>�7-�-R�E��ꕖ��}�?E�?� �_l����ǱǙ5It:�}]V=���&wHH]00�]	���D@�Ax�n�ܬp]��4�=���ww��M�s�.���'X�4�[���\��5HER@�v�GQ�RAv�r�g��-Ǒm OkM�)����`�lrD�Tzl2��H!�E�B�l��	�r�Z�"�"	�Xп�Ɇ���Bq��@�����UYݒ����K����i�"=_	�E�D����@����#_Bݭ�蟚]�Tآ'��g�~��RU0C,�,�Lm���L�_�wߡ�5Tq�Hwc��1�w�rd-
�hPf�p�����zA���$�ڠ�L�JcA������P>� �[��yg�<*&������OjDZ[N!��tEfP33
�yG��T#�D�1c0'h"� ��T��ߨ*5!���? &~�.������o%����WH�*w�Ց�ș@�t�nx]��si뉱	�jA�-#]���%Ȗ:�+�	bk��.�F��հ�i�c���ܓ}�v��Io�,�N�^#�n"�CEs-��T���9�1�śN�k�gv{�q�1�.lb\���X%�s�=󾂐3a��@�]I�C�a�X]Oty�,P������ɺ�v=>�Ax����&�)M�Pf������Y���<���"@U���r�f��K��#q�}��������}��#)=< �j^{Ƚ��t����#�m�|TG톞�������n�aI)�r���mT�=G�S�E�~B5�ܶM@�<.�����9#dp2�%R�09\�&F�X�J
��s��9tT���ttc����s���<�.���x�ْ����G�����?5aCi	:ב.F��̈́⡋�<0A��A� �z���<�jޠv��`�ʈRl�B���vl]��#4�G��z(^����e�H���A`Kŭ�R�4�y���~�=�l��}���8��5�H�H"����R��د)�A���
##�N0Mn=�Rk�K�� B=G^��a�����n��?�7 �v]K�^����u~E���Q�P��)�����V��@�q�	mki|�Lk�ȶ�er�Z��5��j�^e�x�$_��N���F�C*������4̬�H��*=w��M���>2ڀm�x�WW>��>r}[��PdMd4�;N�ʠ2Kp�����k�f��(�'3�� �!����N4�]�j�Ή*�7p�>��|��7�:(L|��n�n�&��B�%�q�R���UD9��t!H��x�ڡ�Ju{�@9��\��E_$Gݽ����Ϡm5.�KsR�s���7av^��O}������[z���v��.a�j�+���yT9B20�we@���@�3�I�/mɜS�ڶ4�;
�"j�W�=IAv`2^	g�M3t� J��f��H�£�4��$�I����Gp�<:���/!x�p�+1���K��!�y^ ��V���z2���H���gqu,�p�p�x�����:xt��u�s:�u%io�f�ʖ�L@Z�i���=$i5�����n�#q/��n//f8Ɖ�k��ÎC�t�%	�]k�6���q���Y��E4�FK��(J�C�Wvi�v��)�_s2�ʃQʾyߞ7����r����d_*$�"��;i��=	��x�m�ڳ�,�	����kq���|��:;p� Sig��cXh/gpv���i4�6z�&1"FT ��GV�	m#��b��I@؋��� f��S�h�X����$g$|���&k)m���41���_�D������y+aAm��8�Ch/�ْ����gj6���q��9ӧ�.�C�4�P��Z���㈫�S�K�1Ād���H�Y5�v�!�(M_��Q�D�6q��A<y"���(Fs��w��B(�tH-����S��WF�d�"i�h$�8	j<Q$���pMs�m�(�k*�"�-W�:mj�^���I��0��䁻��k�ɽ�`C� >�7�% �{O����f�G�֑ ����[�,�"��JFB�K�i2N�7�M��	l�8�����Th:�~���֜�@@T�F�����1r7�Bh"�eei �3�DYb�8ۀK��l{�����u{;��w� g_�<'�ǯ�7�����*X��΋e8��	LuW�Z���Y�܉ �� �l�T������I$M<螬��H!�	q�jyM��1_Cp+��x�����W�_�����R���w(�E@�x�䢛���17e�Z��F�1��U�r���lucc���=������jwWjL9��5fN��\�e;�3��B%���s�;�qpDx�0A$)Y��
̷\�;�~z�6� ��du�k���4�Z��]g41�	W�]蹜��$�2�����u,�-�H�2N!�o��gD�;�1k:"3A�cTO�i�ob�˛���<"��HR�N �5���tknqd"�=A|��'�~S�d���n�aS���otZ�N,�5����~��o��w��3�tu{j����l���o2�����ƫe�;nP��}4&.cPɻ�E+x�Xo<�P�N8����U&�l��tp�]�����0곽��֊�k'6����yz�؉�tAG:���݉:A��qd�#si}��}+�2�M\�@��-��6�Oy�{/�����ak��Oh��	��ر�y����j�Q�v(D�Mo�q�?<g����^<դ�>�az.�]W���<{�7�\�ٛt��h3D�;��5ٔ�;�1:�vh�4t02wp6|%�53ی���&�9z"�1��R䰭�yn�kI��qD��T�b����&�cY9�L�����3�glE4zdܔ;�/ ME�mZœ ݩȪP�}���$�A"�A?����Im��l����¸�D��4T\pF\��G�z]a"�/#�o�7�ˀ���e��G�lkVqb`B������7Q��#x�-�Ű�YY�nn��K��1Ǔ�.��ǃJN�s�;�1�s�K(w�78��=�p׍>��h8�z#dG�^�]�Fg�V���k�g*茑�h��:\���F�d���h��}�+�M���ܒؓr�k��3����-��s��0m�����<���h�E�v��	Lf��N�Ѹ�$!��+5kб��+6�#l�i-��ά��'Vu����W�o�m��0�a7K�ƹ�Fa�T�ZgcXb��Ta���M��p�gF�Wh�"֭{�*�d%�m�Ð�*���N�rnb��5�Y���6��ا�!7c$����]��J����`�/�rV{�ܮu�asKQ�,y���Y�K\�4��K��m�X�-��2��X`��1�mqMM���+�\�iY5Ov����x.�Euu'=��V�.u��˩ev�X6��-��ѳE�'U&h�Йs�
1����rB�����έud�W���c��FyΪ������.Ū���f�1�-3��f]��.{�'��ݸN:��Z�]�8(/+�k�L�33́��J4\�]'y�P�(Sm��sl��W"�2���%�a�s
܄HJIG�6:h��a2%F�\]�٣s^#ޖwi:���c���ٚ�ʈ�6��(f!x�ٌ����1u�[l�5�+2܀�ꭔ�F:��g�.��E�]�3,b��-�ڵ��	JM-G5,�7Q
��p��DW�����<h�F�S���p�ҁ=�ްvVݍĬ���s�<s7y�㻄�Y	�3�s�ܲ��n�^GeD����V�k�&�ܤ`�]n-���%m��G��2��C���ӄ���n3����vP����~֑��+{���u���A�W�Z��Qlw�nP���rs��>�y������BFI��1�I3n a�ǚȋYtqwl��@�n�L))(a]��Bp�Qt�@�.P��"}C'r(3a�/S��3<
�
q�{�]8�N��c���8�]e�m���M�33{��HȞh
t� �������I&�G����&��@G�%����Y;�#)�j���eV�]6T�wV�J֦~��7��u">�c��a�c�M�9����| Erx�u.u�#6=?`bf�DE��dN�$P�33�Pǩ��iL$�Rf��3��^����.(nB���^��'�4�e�u��&��R�.�#��n�0������A;Ё��LU���z}���
U��H��C�ȑ1 F�Ӕf�bk�`�5fz<�t I'@5���59�"��v���xi�]������9�y��[���ž���|���}�ܝ��j|kS���Q(X�>/��=MD ��!��Ø��EÖ���~]QN����XD���1��Z
���g��lC��"�To��@f41`����=�@���9PؠgO!���r�(3Y��3����#���m�M�{���}�*B�b�H {� 7�*k��� �-ӂ��qS�.��N[�́��I��P ��h�VP��+:�bmIf�h��v0&+b�Jˡ�����|��.�:9�{��3�~-+�� �O���}*����[$��h�@cT��ha9�*=���{���3�"g ��*�OEm�$����L))(,�!Wv�$����Af`H��
�qg�L���Vs�@�[��n`|��/z(=䲒d:��_�5����e= .H�&�&�˄I��� ����
|��oM��6�<e��'�9��5��2"�4"�Q�mة;�3!Qh�ßrNs���5M1�!��۳ʷL�`��洅Ium���u�����l��s-%�3q��-��8�`1l�&vVU��ٵ�*]C@�y; j�n�Lb�K=��;Y�kZ����e��-�/)� �O2��х�T~�皇�ŗ��m�� ��ȩ��UG����c�f�@�ɞq�"�<�myP����j���q��Ε'@��D��C3n˼�=Z�da}.� =���:�����Or�T���\Q�6N*��R��5���ǖ��^�����ʋ�X­��.��DL��p�,+�6�qsC"_q��Ĕ���_0$�Cƶ��-�uC��B�"�n�fи'[.[Bj1N������. ��Gڐ>5�>���9Xp`RL��{��3����|���@��ޮID���o��<i^G�^����9l(؂�2/	�f���8B�Qt�T ���y���B��7e��g�H��T)��7q�ҫ-�Q���QvN��[��=��*�#)(DT�*�,!7f\!�y`�D��<|0e�ŀ`��<��m\�N�7y��p��QU�{���C������T`�k(IJD�����c��o�T=��5������sc˚��~�6�#�؛n�_�Z���Y���k;�\��#X�@���={�j��.�?<	A� ��B�2�kɷ�~��x�e֑��5Ȥ\�2؍n��}�������9އ��Y(��~��R
A@�i��`]m�y���u�2�RP��5�Ӛ̷`6@Ω���J�Mi�}�����%H,/�Aa�*A@�i �F/~�Vn�n �8.px!4,�0|6�Z��RZ|SI�H)t�q��p8M�*T
ʛu���*%B��TĂ�9�:.��[��XoT�T;�͹뇬v�:H)���F̬���@��4bA`djB���@/��������[��ˏ|4a_
�Q.L	D,$ݭ&&&�7"�:�� =�ῄJB�ۭj�
���<9..nj�ND
�YFJ���4��m��&$kZ��T���4�Ad��g%��zq��O�����������W�p�j8��͋6�G��?'��׆���AH);���`T����& T�;���֠�*AB�w�1�0�9�j������ �{�4�Y;���JÜ֍�Y+*J�{�F01�!KNy�e5��|�s�'W}���ϐ_��19�9�]f[���ۚbd@�����S��IXX°���뾲�����
��u�1�Y++%S�i1$� A����<	�H���n"<)�i���_7��
�YD��;o����l�P�C����q�xq�����a�
��!�* ��h����M����{�t��*���R
CM��fR
A`�K���Hy=!����y���q5`�#���u ��<��;�x&�����Ns�����:l-�R5��M����5�E�t!���\�ⲵGc��E�!w��:;]�L]x*a��46���%8�H���F͔Ť��][^[�mjl��/+�vr1�îYqn6F�F.�Z�1��WE��sJ:������ͯ䓤�9�bAf2VVJ�oLI�Q>b��?I���{����lļ$�MA|�|������PI]�W$�I��Xw�j
C�Hg������q�4�R
ANw�@bAL@�8�Z��d�q�:�7�<�b����xp�S��sĕ
�Xo޵ �bR j�gn���]��<	�� L��+<֠�5�m�f7`1:���:���n���:*f�Ę�V�az�2aR
J��Ldθ�m�w�E�vVJʝ�I�b�θ�&��� �����jB����;��B�|5��<��S
ʝu��̌� �P�bA`�޷|���m����%�6��-(�^���z�1�ɯ'����G�bAd��;�Z�Ƀ*�S�4c#X�r���AN��i �HV�s�j
ALۃΎK����qy�P�A�|϶�,�w��f��#��?{.n�ͫ�M�L���OZ�/)�Ȳx�Z۸��O��H)��fAa��IP�*u�Ld�T���u�����i($����I8��X3�"T4�-!mn鬤+X �����o��m�t	��R�V�AH)C�i�20�,��FQ���*w��ߍǎx
�a
�YXk�j
AH(�M07k� �=�9�n���A␭C}�PR
a�s��s1����M��$`�R
o�Hlf�ݵ�\t°�� ��*J��Ld�T��S��11����cѭ�GtXN�v�L�3���=�vxy�u�ў0<k�֠�0�������
�S�(H)�:���nü֠�1%@�i�0�)����k]o
�S�P�H,�v��fw�AH(%@��i��R
AOߚJ�����2�Og�n�����bޏ;9..l��N�Y�����`�
°d��3��6�:��y��̰XӇn/Q�F}F��n2t��t�W&��������p�\(�5_#%��0�ļ���KEk�m��[��ԆM�}����3b�tl����ǌ�����ra1+g�a�� 7������,s���o�ނ�w�徻��/��x�]�R�V��-��cܔz�Ꞓk����#��<s����z�)�xao
{ݜ|���_+����3*�ː���w����{�;����܅���o�dUX֟=aL�#c\w�D�h8*<�މΚ���!j�O�Zy�}>�Up<4j>9���y��:OC��==m�E���lT�T�/�u1�V�u�%��a8��ܵ�K�O����ï-k98GC�}�zf��y7���������݇���)r;A
{z�f6��k��Z*�iyd���i-.��-��ӻf󖗇[Y�]�% =��ݹIs���>1�GIl#�Ku�ί5��Yt���9B^\�(�Z��*�vMR�͚�#
�,]�.�]"g�tǷ/�v���L�P�d�d�ȧ�F�ǄO ��1w��x2y8��c�YjPv��x��ɍ��D2�cA���6��cI�&1��ް�B2&t�������v���*�ڙ�e��:@Kt��)XQ-�J��Vk�@8�4
AI�ID��bAd�ʐS�J�0㍼wֱֵ���a�kA��o�6m��Hsi
Z^SI�k����1��=栳9�s$��T*sLa�+�ؽ�em�p¦���1%����wdT|Ͼ�7�^���W����jB�q�I
B��j
AN������YpӃu�ء��%�+I�@�r����V�d���s��6`�YFJ��S�(CV�a{�2aRu�۠ě'}�&2�VTۺL<6ߚ�h͍��Z��䴅��^��@�)���^/|hH)��:�5 ��)��˝�'@��a����=�td�	_�0݅O2����Xuƴn��YR
���뎺�'L��R���
Aa�Z�vM�;�丹��N�y��H)8�$�(���Aa�*AIS������y'T�鹺�(�}Am1�^��ͱ��q�ӳ�ۈ�5�V�CiT��9�� � ��OA� �|�4����n��j�[��Xy�j
C�H[@��i ��z<��
��@�bH,�m�j
AH(b�LH,=5����:�j���Wn+�hma��v�"��<���#��AM����R�֠�`2�;���{uy��AMw@�AH,6�Z�����o��s1����o)�� �����'	��!�J�X]�̂�T�
��S�}���~D[� �pXBla�p5��kA�H)-�)��+X&3䘽�9rb��IxX$��A��I���w�1 �Í�Ì���|�z4����D.;H��>[$VJ�R
�}�Xԅ����n��~)���Ap`T߳��K������9d���6�9��t�M$� ����;ed����8�7�n6ߏ3+|�OZ;�ȝ5�l�"�U�[���d5nz�?:g'gl�������1l[� �$Q	�ܺK��GSZ��wjê�PT���f���Oa%���滖��`��٫\�������1X*8�\����s�����d�m�j؅�VK����"9��:鎰Ȼ����GL7at�6�q�g~j段ى�փѩ!K@ۚi � ���8㝸vvi3|���P7�a�°��ly����xp�S��I���_6�0��j'1� �y�4�X5 �}P2e ���:�`�\j����w��s1���4�Y�%H)���|���L���;�l)����Ϗ�IP�uM2c+%ed���4�&	���BhY�O$Wc��՚G�HqhښH.0+FJm��Ă� V��Af�Vs涓d8IP6�a�
o��f�ַ�0݅MuCĔB��Ad�w�����n�bA`cRӾ�H9HV��u>@�@�������#�"�I
��2�֕WX��߽���ͯ��z���
��YY*u�H`���+ϙ�Xc
�k�l�q;�Ɍ��������bb��w��]ks��AHpZA����Y���7pl��-bj�����q���,ev�®�VDΎab��������� +`"<	 ���Z
Af'}XbAH(k��p��;�i�`�A��tbP*�0�;ށ���R��1���T���k�Y��	��R
u�2�RP�p`T��:�Nf7`17I�T�d7ל_8��o�:H,�$<�!� �ߛ\���gsy��Y+*k�LL@��<�WFln�Xg�9�$)i�m��[R��3&��o�~3�����_%0۝� ���3vJ�IP/���~��]~�C"�����m	�F+�60�J�^���#�F�x¦��i&T�î)�Ă�P8�`cX��7�t��y@��A��a�H)�����������=��Y"�zn��+
°���caRX�IS�i��O��%�1�礉P=�I <���T%BH�ýP�ą�������������[��ڇLl~ܚ7:�v���kٍ�v������K�X���u��?���{��������r9h�%U�{ك4�����D�;�5\��jM�2��YȭI�ӡ~$r^D����g	����e};��O<�;����%J���q��P��K�{�V����95N�NDy�VF&���}�>�P�w;Q�8��k��+�~@:�A$]]w'��q"Hz���N8��(f����pBl��j�-Q��
O��У�v#�|�m��5rJ��!`991����v�o]O����>�H	�ʼY%I�Я����d�x�z��^���G�\N��Uȇ�Ss�ĸ��r�ڷ"��w��
�ǳ�R!-�@�"��̜�*O��ܸ�A8kzw���z��H[^E��*��
��H�uF}�i�X$���^S��0)&l��Ўm�X�ă���$�p�����QY��Vq%{�^C^7��"��$cK�rI��D�[1�r��X�n�p��8��ٽ� }�s����[�#v���JK�3�+f�bE�)-ժʓ,È�s]0���J�����
�݉3R�,Yj�b�%e�՗R0j9]���3���a%�-	[�Z�ѮԒ��fQ���x3�9�ݝn��u��\**���<����u>�����'ZEf5.�wRv$O/\vJ�*{W����u���"�0e��ۥ�98�ڬ��]�^q�y��-�7�Y���_�
���)98CnlKCl I&n$�k�B��y>؋H�=}�s,.w���dy�'�վ���{��S�\��+2�c�H�5�Y�MV�^���3�O6��%z<�q� �唵ԉ�M!ֆ��T*��̐u;;�K̜�j8(��]P6��[��+*���jA����� n>$E쀀�����?~�\*{j)9�X�$�]�I51|�xY���2�D�޹�7H�2&�ˋ髒B�I2D�3P�$��H�@�n�jD$r����^�I[�}j�����~9�ʂ��r�-R��]�wt���\�2�z!�$N�$�$mڒI�A�:�s�"����//�"��TZ���#:,�Z�r�5���9��t�
���<���4ݙ�T��#����շ���Z\udi.��+,�=t�����9��$�����^_,t�����|�$��[[1B�I�2\�PrdMٗ@��EoNЎ�$� �}wj0}��l�|�.3�=9���+�S*&w��D$>�	�GlM\�CK���a�HU��"2a�R�J� ��I8�E=�������JLB,�]@S)���Cp$�C.G�T*(2�$��N���͉�j��f"�ώv!�\a�2VX�j���6iܬ��q0���x?�OO����T���E�ڬs)���WPmE�\>��S��-{р�D۩�A�[���y�4�߽�ֱ��9�i�^#��4/m�N}x�&Z�4�D�w�V��"ۍ>̀��d�c�����#�r@�:�dvV��B�q��ެ��!)18��C�d"%�̂I��ѻ騨�1n��T+�Mt!{]�q2l�v����/�1��_z�j;t>Ve���=੼E���^����w�sT���XN�sN!<5�yT\���;s�}�h��J��o���jT�v!�<�^�f0���oT����:gd�B���|۹��ػ�5��&dV\Mcp"�¬�]��xj/�J����7�2����}`pw�%�h�K�����R75�;^N��M0T�^qWP�i�	{�U�P�}���n����z��1wd��A��ɯ�'s��x������FP~�:�F�,CW��i�}��[�iw�iŌY�r�P�^,�0����*CX2�+vD�w.���e��V��c�'���F�<��3�(��������zr�q,��,9���@��x#�W���e<
���=t
�j�K;��.u�ȓ+���6��?��s�ZwJQ��,ut鎋VV��y|��1���\�D��d}��\�rw(���;#����9v4�c���Y��/�`�����1�C�+L8p`Kǫjϥ�����t�1*쁁PeL���¼�D3���ǌl�C*�F_X���aE�R^P�.<1�ǌc gυ� `D<��S�4
��s��5�Ɍ#�����ww��� �>�ĸ<FL��G�L��f�0ͧ8.�>N�#���n���34��'3������G�L��v3v,��1�%,c��RZy[!��h�)Ic1������f�k�r�8�>/<�v�qAY�[���B���WS�9���suY��q:�}�S���ƒG�=�qz��͏]
� �txz�+Wm���7V�j�JܙՆ��۵�7pa�89i;.��`��-���h�¼#]]SQf�& ;.�،��,�ؗ��V����wu,+��f�W[f�ˉ"KD.�0vh��8�h���"ǚ��K�-��8M\�tu&�4u�e���sY�k��b<�hn`�ګ�D˟JG;�oOt�hit�N���Wc��j�q�nng�k[�q��^jZ����ܘ��W��^[q\E�F���su�n�y���R����Pn�xlM�J�>����E��[�y]�U���-j��˥�j�Y4�yn��]��6������]�:z뫶��b��Gp��z^l	^��eq<q[�����h��R��㴬��K
[�I�q�`Ơ��Il�im���ےrr^�����ѣ���q���)JJ�(�YFjW�EMI@���xY��O��E�%���XM.�Lf[>t�(�[�n՚�0��]iJ�X[V�e���6�Fe���:Ri��+7-P�][XU�J��;������?��9�6��g���{"��"io!	܆��U�Ʈ��΃jDD����m�l�Բo;ۑ���T^��C�+-ch�;�NՖ�^��r����=9�7�v�.ϯ��}l4�a�V�v&��K�B�S1+o��]Ҕ���,kr���Y�TL�=����<:�L
oyߎ���x��_����n;��aث,�̫�� ���õ�7�{�ΪŒ2��2&��C�&f�sϫu��\�)`�yGy�R���s�M�;jz�#tGU(�6�ghSʮ=�mA�-~M}%ƻF-L��L��A��FLD�o�
dDQ���g4N+�a���;CBZ�*';�⮋����h�rqΗ:%L�U���.����)G�ǔu朩j޽w(F�j1Tm�Z-X���{�/���}���L���a��~p%��j8��K���a�R"$7����4+n=��srl*�:�J�[A��� ��R-8e�S������!|��uw1 _ru���8͉܍�W�bx��;��̥��h����;�>���gtb�T�6�v���yur�7�/W����l҇�l1�N���b���}������5�0J�QI���=�����&D��|��rv�bq	�C;P棹��S���k]� m4�b�as[a�L����Ԉ��Z�]�m�%�+�D`BB�{N%�Zx��.�6���m7hM�236� �cu5��.�J4B�+���6 ��	�|��;]�b��T�.�Orcr�2�6�y����{�L\�G��&�a8-�h[]3&q.����ԭYt�V���<إ���v��q����<cg].7w>3p����nx���)H&y͍v�1�;c<k��Km"h��q^��\j�J���e��,�����[�6�K���qj�79ᮉ_AN{q��������LDL�o(�2'�|�N<9������7Mƞ��fQ=�s;�ת������y�	m�4����Ȉ���9Q��*��3 �3�k%9�hcu��^HU�
4%�.u�7�m$�nȠ�����ƻ,R��J:1ȷ�LJ�R���*Du�N5ͨ�a���p�:�rdM-�b�A�܋��JU1��.'+�6_ƾ���z$o���{�xM�Z���ɟ��g�r��J`Ďx:�z3xj��u��Sy�	
�"�uow.�f�>�зj�@{�U������*X�w�*i:ť2&Q����.�+�����u��K�|�	�^��9�k���!�%��!:�t��$��wf:u��	��2&�j�����z�@��A��	�s�U"f-P��!�k�(����<�{��5Y�F$7����>��ي庽}�28�4Ξ���	��`_a�u����j�]�e��%��U*��	E9Y��UJ�*֯=3��hzR�oO��ļ�|����NB!Y'��hh)��l�2�*�l	ր�w �whp;yy¥L��&���Gnu@�hos���Ɲ�p�>Fy�ʮTI��j:�v�I���*kA�Y�Z)|=���Q뿡ڔ�M���[	S6@:k�����4��
�,����Z�(�&�f�ĩ�:�����%a�/�'עr����C�V'U����f�c��W��75z_Guyl�0���E�Or�L�����l��![�j�_��=7�6�XƮ��&�z���Zvmq�z����hR���4/�04�T/TBC1��/M�sn2�!<
�Fۿ� ���Ղe�Wv7vŌ2b�TAXf�U���9�,XN`�~��:�GK�cTՋm�Y����r�Y�)�v��1�н�\<�XŸ=qi��{RU�Z���W/wcv^1c�4�i�MJ&��xRfTʉ���}����v�;cy�uB��{�����\��{���~9^#��n���.�;N����,�b�ӝ��R�Q7����p��?Ms:�eǪu4��!m\���<z�r�m����]q�j�qG�i�D���#��a�6\��_~��c�����V���;�so��7���JF&�|�r��"�N����0��Ӎ4N+�u�̈K,��*�����<  
��=���>U~37��pF!�R#J;����m��_3��]Z�(�U�kk�oE�@]�p�2�lR܁�ژ�r�Ӏ��z��BZ��[Z�ximx$�SV����3)H]w��m�����yx��\BbDRmWǫ��Z��ȈO�Z{t��yvzNq���Śd�� cud͠���H�h�		�b"�=����	c����0*��ܦ���ݹ�J�?PG��eR�]��Y�qpb�˛�Ƿ/��a�jUW�U�����e�S;��[�Kf��qd���[SMD���Z�C�8�z��S��^��S}��rd�8Y|'�J����ݚ��{gp����Gf�����g��o4����]Մ爏U�/�+�"��˷(�k^���yA�uo9��V�O���a^���f��1�QI'�3-f��ۖ̙VyͲ�Ξ3�[w�Z�D�C��׺������ϗ�ӉIG)��Z���zZk/�m9/�L�=����	���v,^٢o�� j���gK^��p��	՚�c:|�q��D�f��j �u2�����˄op�!��{+��`Pɐǟ;�f��=�p7bA�|��)8D {&��}�>a�y\�s��Beq�`S�cwN��_8�z޽����#&%b�px�TC�6���*�ú#�fɁ�%Z�Yim,Dr�14S>�jDv]�)��q�{ $EA+Kh���������QDX+�Q[J�Z6�X�JʓIE�V����$=;�=;�S�׼�Έ�d&Tf���0���,ec���A�1��K��w y��sP�;Gv���ί�>�������`�e�j!1
!L�M��0��]�K�� ޘ}}1tg��^y.��3˻�ꉎ	R���T�M��q����������hp6j�bh�k3�pԽ.�a8���L׬��Q�[��}"���L�s]��g�r֗$�|=�
������:�U+���;;���6�z�уWy�߿a��(m�[�2�`2P`�����Jh����{��r���0л���aɔ���[@k��@E5A+m�*S
$N����J�8U'/ {�9\�NI�M���U.�Z��oK����H�λ�S��w@T�/9HN�H��<�Y�U�P�"(��.��(�p����EtT���J���x�b؅���ݓʽ��>�/gX�;u0u��W ���.Ѯ�-��gD�uSZ�f!vL�աs�U��c
�"K�ͨUv��[i�����3�vܶ�����H��u�ͧ�ԝ�wpO\�C��2Vm(2�s�%KT�N%32�~g�|��z6i�(�:���t��ȈR�7���ޚ�����A�Y�-o�����)W�$%�*'���1��T�&�>�7wQ�h��ɛ:���)0b��w��j�7�{~팚����{>u��s�RҚK#��2eO^�򔒞6ӻC:=׽��tJ˵��,F!P�#�Ou�qIY��ɉ�����;��W�m���<=U�z����=jj�V�鄥(flK�L�Qj�\1������2�:SOr$��.mUQCwP��T�H�˖��m�ʹ8L��!��(�)J�&F��)��h���/�=�z|��\{����}�S|��t�e�I)�8��^ޏ6о�w�^��ݳ�0M�9�G���p���p��S���a(+��_�r���W�3�<9V��ze�GuEU�)�����k�=���L%)C3_fRC:�!��e�3�`n�2L�N��h^���y�mx<p*�nv3;2�B�Q2H˝��
�+܊#�}=H��\N5͡�.��Zh���(��-6�oqFɠ旛hl��.Ԥ��mv��rQ��7��S\4F!S��$Q��}����B�)�qa]��4cS=n�^��-��	��t�;fJ4��o���{S^���	JQN)	��n��U_b-xc������F�30���C[2����c�{��ap��ؤ'u �Wn+�q��Y�J"Dש�zL`*C��c���]%P��F����²�ˡm�ݪ������+��9��vR�Ͳv�X�����F!S��x�]8�����A9��}|r�~׵vvq�vl����=b��`Td� ��w1���FJM�=X4������6��*mFC�,���Yp��4���"��`�5,�AtWtPt�r=� ����u@�F7
z�S9�wG�\���.�p���̵�u����\7-��pҲ�!m�FkIT����|!)J��= n��8o*8[%&WL&̘�7��)�����}*"D�`��&�M�Ww1u�Td51�"��3�L-���mUk��,܋�����Ꜽ^�������Z/M!�,`�Xڔ��$x�Q�&n�p����eR�x$�����;RJq��,��.�����T&��"��􄧊�j�q�q�r/����V��O���'��{8'%.P���Nf5n��f��beDH�v���T��&����Sڵa��b"�D��U��V�>��7�¸�X�ƣL�(��*A�A*����|��� �~zI��C�"	�!<��1w�	��c����yY��(fr���®"�wht�JJaEtR�Jpb8����(�&z��Vc&���rK�9�P�Q��n�Na��W_|�;��s�0�JT�V�B�#����Nx�v���R��5�w��J@m���xڻ�3"�(��.���70ܮ�q��_{�{��ە�=[ ssѬ��:���)D�mG��P��͝���T�vWs��0
�������K��e;ҡIQ@8��zT�)^��jн��%�9��R�i�*��=bpDgYLf��VvDK�L9�+n�9�U}���v��	0���'�}�Ow^@��񍝯z��{V�(RN�HV]3Z*���Ӕu㝚ʞ���j�Ӛ۲���aw/dY��b"����w�<��IywQ��0�L�;6���p9ם���5��0Ux��r.=��Ԡ+�xk�]w����ʷXT)*3��u!����[�.:4J]��12��[ێbn�!�5)xnvGa�͋yR�a���3r��xx�x�˞��i��{�4��W��-�9��|�R5I��8�(~S�K���^t��n�	(�)cՔd��}쐏,�o����{�0Ipw�c%������w�A�� ��Ź���`�9���x������;yy��s���6�5�k~����<9`͞��>]���<7��ʜ�.��7��j�(EJ��h"S^W�)��
����zB�y ;/b�(���P��ک��[i���4Sɫ-���I�]]ۯ��Kӆڹ�*f^�p��ZD�r#����mwZԄ�N�Q6ޝ[N�t$�kB0,P>Dx�nt��J�=�3�o�i1z\|��� 5�b{k��T,�h����6����5�y/��� � *=:M[+J���V���UEUU5�V��ə��1��c+����xщr��U-,K[Qm
�Ep��0�h�F�/�eb,@�V((�%�R�Z��j��q�ꈊ%�R
��+\���O+�* �'��,Um��-��q�T��R�*YQ���(Ք��XЮZ��#�1߬�:���\ f�ܰ;�1Yy�ڨE��6�jf]cuҔ�i��x��d�ۙ��MqU�1Q]�&3��2�̍"[,��[(�v���;�h�r�ņ�I�&"x���8R��Ҷ��B�X[��XCA��#����#�,盫b;��/�wg3�y�M��I�λi�[�{Z�*E�&]f̗m0�pEy��C��\����S�s��G�<6e��i�ܓFF֤��nT�փwm-�{f���^������^[��3y����k��:��4[��Fi��Ĩ������u���a\ķk	c�5�k�
h�s�&�!̺h�8-,nn�����q�C9�:t4x�k�;��r]��M3�E��q�Ý�s��#����:�̳�͸2��u�;����=µ����<㮺�Bn�W�&vņe\V�m��Yt(�f/*�+�٭��K�f#J��뭖mE[t��mk�m�3���*��#��9��Q�]۹�M�'�ܛ�8�],v�A������N�m�۝���������具<j�Pqv��uƼ)��W�t����v�.������s����6�R`B1vH�[�`�m3M�Kv��pᑺ[���bM�/-�Fc
�!�\,���ѡX0ZWT�Jl.����K�$����C`�Alϳu{�`��4�sq>ջO}7h=�*��U�fx�Q�WF�Y�6���6�'��Q!�������P#eMoh���:�)��X�h7x��9��s��$n	��i�U��6]��`��߾�b�n�ʏgt����ʚ�ˮ�a&��WD�Ч�Z�s�W!D_�<�LZ+��ʸeJ��c25e�rg犙߇�|��&���T"��n�[^$���nǳu|��*!�nw�V�\�C[2�okwJ��h<��o��Ҽ�ev[2w�c�>��Y�3����ڴQ�IR�S3*i��`��ѵH��B�zV�PЦDF�^��'�� �^�/#3�����%	|�sN��{6bDb�����_��;�iS�W d�����Z.���M��	f������Bb!S�1M˶�?���㞎�)>�
f"�5]qtn��m����Cv&3\�vz����7���ZKal�1�顅�����FF�v�;b��_��y�)�`��C�����Jj�7�g@C�/n�=�C�̃ⓨh��*����%Z&\�9�r���y�TiY�b�w�7��Y�
B��"uE��@�!���܆<M��ۙ�qq$0�>�P��Dј�U�������K��͵��y�s���ىqm*6�V���fQ$�LDL���3�S���9�T� :�]%J3E��P�۠k���F����T�R��d3K"fP�^� K��;&d������$%� ޮݰ���)�aH���Ձ[�����n��l��Pv��l��MdUA�"l�1�R�y9�,֩f��b-
�ӐETM�fO����+>�lg]�t*�kZ,��Eb�\�Z嘱�Hmu���^��ڞ���֮H���mud�<�ci9.��ny�����W!�nU���Z��v0v�Gj�k��7Z��uuE�̖鸞ø��	9s���GϾ�Osv>~K����X窎�.3�؊�P.‶w_�nr�j��;��hƔﲨ�o Q-�9�K��Fl�:� �&4�*dQ
�%����8p~�t����"H|ԐO58��Q( NWX�3 �qH`!�R���$kAA"�&O�R�R����{P�����BK�8��n(uBs�s��I����j����Vd��ZDR�E�� ��ٓ��nT�
��n���h���ֺ�dt�SND�3&�����f�1T�E�i��;�� �w�@�����{�ͨ����J�	g!��m"ID=��ihD�-�E�e�W�A������caC�nN�K��|���x��B=��uC{���)$m�$n�F7JN��`YE�^1��9���:L�*�R�H�A׊U;���+W���j!P���,���#;�cP`��q|��C;-��=n��d��r � }z��[ɝ���dtO+C��3�w����ٳ��e\�B������&~�����D�5>7�e'T��{��>���j v�O�'s�N��o��T�0x� H��p,i`�N!������-\��C�I�U@7B��5�qS������z�p��O��Aw�I2n$����u���*���#G����o����r�U�o)�>�\�Q
��d-�$�����%� ��x�u�ZL�&t�W���� ޳ �㌗p�N!�hn�z���ʩ��`Y�h�=��h������w�o���
��N3�rH=�:y�.�.�\�@��R�������5�:ﳸ}�h��c<A�*V
����Q3��b`��2 wh�AZ}荱�H#k�I�c"eF��m�f3��!$��^}G{��Ar�	���P�� .�Ey�q\̥H݋�������-�s�=pG^�$��F<1Y�ՔwHv�o���JeV w^���M����$����G�s�`���l4P�-m�!�Y��B&�Lc.�d�� !��j<��!K�9$*r�]��c\��K^�2�9l���h��7\vmk��vxEY�F˩I���Fl:�H�u��^ݻM�n�驚��糃ܖ��B�iX#�.��\�fT��ʒ$v�
�,��rҥwwƧE8��~B�HZ�Dh��uP�ȐE�N�E]��pi��/k�P�I݄O�:B5]�b�8��Dv�Ț��7��^8O��G1zWA�j��ꘪ�sϑ�\�#�B1��,�,��XIt�\,�DE)@>3��n�UW����x��^U�/�~V���HV[������J��c�0���2��Y�1 |h�6Ԃ�l�VR������$^H�Lk���[��Qz���&}��R�lK��LT���X����NQ��ֆ|<.���,�O�~�$������&%va�� k6<���F�CƄ��(� ��ِ�i�.�� �u[���+�j�6ځ����U����yb�dˋ-@D�Eۑ$6�Tp�u�-�SbT%Im�ͱM���Qv}���P�m����o� zC;2v��H�P���n�Ҝ��^��6���µ�WqP$��E
�lE���@ɘTs$�n5���o���]M�����*.��v�Љ���6W�����bƍ��)��xh=�3�a(��_29��%Ρv6$��瘘9:�a]j����V������4�l����2�5�j�lJ�z! ��UY����^�>{�v�]������H����?k��������>��I��86jN�:�k�W15��@bw0���o�@�	�-���s�o��%6�K�Z��kqvt��}��d��R�e�Kn�jC̛��'BMy��<�u�'D�ۓT8#>)�\���P�.�pvA���:�m��z�ܩo��oRG>ڷ��wճ�0��s�^�Q�F�x�3�^Ǿ�ၞ��j;��}Ϡ�7�M�Ŭ�_K�����}[5b@��� $	��1�� ��Hqeǅ��;�L�&��}g�(y"�Z5��Z��A[k�L�qE	�Å9�7� �1�輬f��=�Ǔr��8��hg��O`�ݍV�[R��(�J؈"��Ӑ<Ӏ4(���V�iaR �h�X�ul��d� b3�/��'��#�a��Y,�3�x6mε�Gt�K���?<<=� >��I'��ڹD�P�8f�Om���}�u�A��WqL|��Tw<��A�ߠ�ԫT�kk��T!���E>4k���_!�"��*	�0�#-�����|��!�c�n��7D7�к4�U53�-�E�,q6כ�#��|\9�>�=� -����Zz�����/�7����t'VOP`��;��hd�&aCk�˔���Ֆ������'��VQ�r�1�7t��W1Œ�W���?  +՟#�u�)%`�	.�c+u��b�NZN72\�pԍ�}�:3s%E��F�ڇ0�;y��RD��q�	�d�a��@�A���Ȑ�����s��ȁ&��ْc,Rx���`�B"(� ���T���=j$�@���s��&(:�<�ʏ�$��S�H{�`�*����ygH�L倂o��(fA�^!�R|�	��� ^�� �q����fz�iTd㋰&��a���b��w�U����%�Iz"
.�eK1�L��Ʈ�ۘrn��:J��ǻ[�U��u�v</*��0��+6F����4�fi�]0��Z��֞��+X�����`��k�L�"�%�Қ�-��6,5�т���n����5k��N"����T���e\��y�i��RD\ìn�v�0I�>��^�{e�P�h.���L��ڹ�A=��E�N��$��R>=Ѕ�Q9Co�����T��J	����-���c9%'vT��v�&*˸^"�3�oR1҄�Av�%��JT�/����Z$X�u�ٷU�2T13w��2f+�I&�^��}o�n�R 3d+;��U$������u(Nݯ�6�`3̯>���+�r'�z�l�1򶻮���*;�}���?E���{)��۝�����oZ�d��[�k�H&�yx�זS�$+qK*�d�\�F\ �D�rJ��^��w�1��'<NL ?�O�[+>?Z~�/}�����>ވ�jZD�.����J�H���\���~ڍ���^�Yi�D�y��-���#(3
�t�h��7�3h A��'�i&]U��)���e$��`=v�o��芢���W��(�95�Mּ0lQ{1X{)�ѳy�(�zv��[A	��E���RuB=9{��U��� ܟP9����}- �3|�LH���\�$���T\���F�̒F�K=��s1�\��//n���v����C���_�ԩX����ȨFzDx�D��D�%��4�$���R���̧b>�z� ��`�7{:���,�2fw, �|��c��^�K�"I:�D	���2�+ǟC>Y��tHm�.��v�Z����p�*���쾬�D)מ��q���;aѭ3ڤ��dL��:����(k�>>x��ޅ�{�w��׭��]�F-r��6�l$
0&�_|��#�ӯd�����p=)̥eP!e��S�U:�OF�����̭���pF�Qw�3��f�w��	RL]��"�y_^eኡ@��x�k���L���HƑ!�Iz�uUDCZ'�S\rfT%Xc`v�>�"	)�7 Pm̕ޗ'F�7-P�3����3)���b���^4<8Sލ�s���4��'�.]EP�2�q6P��j6NgnY����n��z]��l9�s486摰���ƚ
��*-��KM��!LApZֹ;ԥwuE�7D��p����x�*��3��p�u�B��\�w^��sIr=��fx�U���!wv���ݴr@�ւ9N٘�%WE!�
�=�*�E�	'ϐ@��RuTcu�f��6��h� �^�1�D�w ���$�CD�&.�v��wc"��q�	�"H�ʷQ�	�K�uHt&��7�:�\'��Vv*1��
:{���.��M.3�+�� ��(���F���'�2 ��R	$�i�x��\Po*��l�UC�Qgʳ�X����h�N�%��A	�{�4��c��~G�^n�A<�>Ie" 2�R��/�:���u�)7�H`#�"].
u�&{�H9г:M�*%�;�r)byzI|�'��f�xr6oD��2{f��RLPځ��SS��"�H7� O8�C��(��E0���!�ƹ��6#����D~}�{�p�\�����/�s�'d����Im(*���8<;O=r��5/��錺�{3=��wA�3d�0�z��L���k���)����8�E1@J�ٽ��M����mO�m�w�I%���t{)֙��U8�Y��Ef�|{aw�7���*�QNoI��Q2GDz��Ћ��zc�� -}>�Tv8�5��!Ynj���lp.�K+�0����$�q�H[�HmȻ
���qŖj��� o$d��0��z-�����=�������o9��Y�MBWf:$���7Gz(My�EG1��L�����>~�}CuF:y���	��/�X"&��Ν���1��D��j�!Jژ�K�c�|��i�3$�lR�A!dN�N�TI�E]���7Ui�7=AuMIPi�C6QM���̰KvS?=�癧P���o��_�j���wk0]�@H$n9�TtJ�bè���b>n�3��Q��� C��ض�5N;��o�D�
�z�v�I;�d�j
jC�e�`>&���<�zD����w����mlf���2,�0g���;�.�@��kA�4p�{�@��}�v��"놝�`/�s4��}��b�R�mHu�ST�S���:�+kŋ`��Sk�5�K�p�Z�Y���(g�k��������-����eMfn<��㠽��f痥������8ܮ���������ٽ�<,�b��C��Lfh=�"��H����x����$��������F�w��g�{5x_6�#�@nL����=<�Z~���x���p9��hä���0��Ͷ����ؽ�O`���Mi����n�EZx��cJe��z�ok"�1���[��CӚ+�_2�����rz3���^*t1��P��وjq�Vс�k�����&�-����a ���F9�9D��TTV;�q	⍪��c�;��?�q{�;�[=G��]��:6Y�"�PQVUb�X+J�����K��(�'��S��&�P]��F��qcdɈ�	4d����X΄%���\���Tb���i�X��B�g	�PM�1�p9굈�*Z�+U�EkQTQ\j"��X�GV�x��\���eS�C�EVZ(���ՅV�Q�0�b�0��y!�����˦�JŴ�˷\mV���nH*WVֲ͍H#���wNu�ݵz�碜;�s��,����u>	�+@��� ��E��:�R�Wr�����࢒������[��(cB�pn0��=sN,��;�Qy���<uC6���u�ӂ�,�Fi�L�����`Л�ţ�sNWJ�z��[�K]�7v:Se��[]�A��XW��rlf��`ƥt	SFf��k���R���x]ŖНcOr�v0� ����LF��ܥ�ghC:�ꗛ7B�ԱWZ���l(���.��7Fg�ݺ�_A�]X䕫v��ܣJe�GIV�R��M5�(�9�ke�/��35����9�cN�]�W�b��ؙ.y��4��h���ͱK�nŠ�͵�{��><k�)[9���'jw�(7�)�b��9�.̹�yv,�6����\1��`��j;=�5�y�[A���kmЦ����[N%\Wci]��	X���]������,J����+��%���Ss�;�r�c�Ye+���2k�uDlaG+,i�� ��9�Q-n�CRɢGk��im��V4р�n��B���lm��%�u����I��Ku���P�5X�!v��";14 ��V�53�CX��.&�v��h"j�\���ڴ����ڡ���Bk���v���E�y��	Fd�j$r���$��-ǐ";�k��/;=Q�T�e�"A��쐻�H�Kq�5��nFP�
\K��|�$]�D�GwK���X��$��১��������whn�r4u���A��l=�l��}�k7٬Q���J¨���d�A6�x��E�n�Q�=��v�=[|L̃a��%�1m�Μ�<Hܣ�u��k���{��'&����f��V2nŭ��N�H���,S���R���:yG�3�� �W�y�m���	��D�&.˵AÚ���Y> ��d�sGc�7��.�r�IBR���H6Ҫ���0������r\��ߧǖ#�[.4�JA�V7�)����;���_�@�E;@s���d��۹��`̐\��LZ�	2�I$n�	�T�ڈ�ޡbfA���=" `;ߥ�B��R,���n\E��V��A�v�۳ϠEn̫Bwر�N�A9�"2�nT���E�۬���yU@� //�w�SwQ��W��g��LPuI��;ѻKt��̒H5���,���~Wu�-��*�\�捘�e%#���}��wƑ�	:��ZA�qy�Y�s �s�	��RJ.����IK%!0�c��-� �A=Zc;:����0fM�$��GͷQ�y��X��"�>����UH}�~�]�̥`�j(�6��H��ۅ��l���Vd���V�4�F/ �%���s�9���ܩQ$q��K��`Ǚ7��&c
��48���+��挄��ʑ"�Κ�$[2)�����+n�%��E��hL�,r���qF�nba	J���&�e�l�Ƒ�H@�� ��8����sj>�CyJIEك�=]k�v��q�=܄�9�ܓ2h��l�!9���o�p���\L�!�^v�sd�<���P��f�-�]��u;��&w�\vr��N[�s���ԪEQ�,���B	�>	��*�q
�k�CK�#�)��T�mBM��[��� �;�F�����ZG�u�j�"�97wa�9�!s�9��Zg����ܹ㎆� ���ʨ����h��yh���zS����(�E(O�Uț��~��*7T,o��s"Y榺C�z� �$��2��bfI���"m�}ir�=�:� /v����6c2eR��m9ډ�%*.d�o�$��7��5ڤH=�M�mD�V8��=�H�jA�X�`:�;�D�<ɹ&dц�$���bƐ�5�IQ�<��{>y��:��;/�PZl�QEI7)�!P�]��	T��>D�� |��+�sNf��cb�/~q��lh�I���f��B"�.����Bō��סͼ������`�{;݇�n��˲.2���B$��\�.���3$��.�+�#�ͭoo;(��^΀�#��D��6�)ڭ$p�� F�T��
 �-s$c*TD]��D������ܗ#�=��/M�O��]z8��+�jk�iD��Wa�/߷���
�z�> 6���تdB�3�l�2]�s$���i@����L������w�hd��4Y��}��IE��̂\��:S�ޅ@.�<�������q����&�1g�`q�	꜍"D]��Q]Ы�0g.>��[k[���F-t���êA�OAƤ�'�("A4�D���w��[��r��n&��:�nW�B�&��c�����g�Q6�{.��4��/�r��	;���9�܃2h�H���5'Pw'�㺗��@�b��YU���b�C�C��A
�_X�ؠ�^$��ȐF8�j�A�2l��-o/0#[�A�d"3`:�=u�w!�7Q�l%|���unjq<�':0����-��*�<6-Sq�dH�Q�W@�mӈ�`�ˑ$�}C��Ƚ���u�1)̦��.аՌ�b�S3����%*�\	"��#�Pڿ6�3r1�*"�p0�yF��VI�=��!9��K�q"&H.,���)�z2����0	����w��&�=��҄�_G�%�}�M��T�HYh��:9@��eN���P>�����q���m�Q����ە���f��C���tp��{�)ikVO��K&��j�I���=NL&p �0V"���fj���2�8��9��̗��8�#Q6�1.B%s�e�:��c���l�cW!�V���T�#M1��沖�xDq�˴j5�ۖ75c��J��%Y�"B��1��hpŢ٭c����~ob���"� �r?M�1�����@���̕0����Y�+���@���1Ϛ���[r7��1A� ��RA59K�;��OE�s^���H����E�}�ȳE�Ԓ�Awd 3��޾XJ�>[�j��F�(�����#wF��N뾯^��7�-�(R�j�:	�	���MvS>��@��VQ�@iHNQ�Cp�D�s'*r��b�V"\��U{�DD:��qw[���7�=on�r2���pe�X�t?�j��%:s��̟g%�31<d?r�%IJ�t� ���I��pi��$����&�s3(�[�|3���!o) �r}�����`���_��N����ڇ���;=�oP~$�	����N<~�����NP�f�)]���mJc��^hJ�<��Hơ���CmY����(�2f0p��G]Cκ^�}Z���$�ى���R�R�����Ϛ?{?{������/���VS�A9*��70�N�t!�;"�0�aY{{�
��yKW�(7�|܇ݯ�M>��&!�wέ��L����j��Tl��&~��{�����u]��L]P`VzK���^:;鍓��y[��]�ó��Y���(Y����;��_�nֳ����}�����m�4U7G�\�/�Vs볞2���v�f�ׅ���<7x�+{%f�
�������7�5���^��1�.�x�B�����hՋ˗��;�h�US���"4o��̰���L����=��Gxrn��:gf�򮣇qy���ysD���6�VX�U�.�p�ڧQ�yL���ƒ��_�É.����� �,���x��B�h���w�������-�T^�mUvq�*�u�� >c��x1Ⱦ�><R�:c���,a�SIQX��UeacEclQV(1cF0F+mJ�9p�0l ��D"��5��[eR�X�(&��N�h�G��q�< �6�
�hi�VQ��«r�"�* �:De"%��+-��j�h�XekUkQeb�"=A�2`D���7���܄>$���}���D�0�ӘW�k�:�$tQ洣Y�
輑�fQ��Ls{(�٫NDH���z��;������-���,�tE
�s
�ח�o��o�����Yy�9�x`���1P��T���2Yt�`�sl�%���g���7�?���O��^b�P�3(�i�Y����V'
�{�D���L�"�n���r빓���\�Y��D���(��3�����"{q^��ϗ��[,�����t�(q*W�;bD�0���=��|w/Ot�\J����vOwN�U*l�e	�	���ڱ��n�+��~N��]�+sݔ 6C�u�/��k ̺�p�-�uGIt=Q��!_�(����E&k�& ����)㫰��5v������C�!�P&J�-Gt�N��2'y	"�/�Qל��+�H52{$�APuH5�)��K��L�$�<~���F\�5�>��������ݡ�<'��y[^<4��y�@��ϝ=}ӭ[.���ĺ\[�sXi��q01�-YB�Z\q�'1��׍k���::��!Ǭq��֎�a�5�%�2��[JM���Z�in����mnF�c�B�*A�͖7[�j���<�6\6�uYmt�ƭ��@���|�ȍǯ�V�o�R�6� �1����Kh)���1Vg��ێ��W@@��;:���\�x�xdDɠcc�⏮�_R�j�4�� A-���Q �8�xЃ�3%�!փ�r�_Tj��y��[R�(��<�kȐ3ɒ�<3G�\.�+P�ڹa)�����L���AMt#��nC�&.0����x�LɄ��TU���4Գwݼun�`�}��֩��.?v�s���I�q�:��8��gL�yY]7,J��6Pޓ(�a��^x2�w<w&��_h��2c��2�](����|H��	�f3�\�1&�$m;�2��!����Q��1^��7{!nI��s5����TCf�H&l�2ږ�z!�����Ҩ��=fD�ϡ��7\��Dn��92qɐ��=p�p. "hH#vi����h|��UT93%�]�P���\k�#Q���<����ӊ��8%���yS�n�(��7w��3�2	#ZFjF��E]�p&(��旤�1�9�jt�z}g�N��?���{�'��x:�uX��������5�(�6�cJj=>|�&A��W>��Dk����V�������BP�*4�D��RiZכ�4�]sN� �d�����ӏ"�b��n�I��Q��	�0�[��輩��v6;�k�$��[s�A�`��R�T=[�`6��O�m�S��X�bv)���+���Vk���|�*ǖ��R`��zD���OE���+̈����7L#M���ԭ]e���v��w����l�n|�s�~sB�Vq��yN��RL�E!�4ԿUL,�	.,��W���rⱩ�Ѷ�ġ2TQ��&�]MO��O�x�I��B+�����4P8l�Z��>�V���Q���̘KZ�����́4MB(�V���v���DP{ש�:��q����Ff�b�\������}:7����}R2�WE���r��ľ��Nǅ���wj;YŹ��t�\7i�[�ε������,[,.�cA^-�����,�Z�vB��Ж[�l�n,SS8.m�8��!�E��뮩щ�#�ԣ��f7EY��˲����Ly�2p�]������� �QE{�	�`k""d��g��#�e���I�z�Ӹ��\�)&k���:�����xTGm�=�>��1͉AHP<=�:�c݊��@x]Ij��*�Hr&3B�v����8��7�H�J�͊!i�nz�2���>�T-���.Kn�n�����fbI��qdg+�MQ�.d�p��b�%+�Z�k��Ɏ�nČ�.n%F7�D����Hc�|�'T��H���+`�˘jϋix��Q'5T-���A� �^fϺ����O�t{�y�qR�g��.�����A>ݗBH5>n6yH��x��gy�SuHOr�8|ޡ�pV#U
�La���Z��ٱh�iX�U���a
��qu@ ��Ɏ��!��\2�̙R!&֒h�aGJ˗h�� �l�#3������3T�%+�Q�Ğ�R&��4l�Nu+��1��:�ʝ8�m�/zE!�d;�|�@Ԩ���;v�U���ܪƭl-�Gӗ��1"	e9�Iw�b�d����%A ����0�J�.�g�i��$��R?�g���{4�V&A!� ���3V�[`��}�ߞD+��#>�bY��y���k��������Uż����ۭ[W��e�}_�!��w��L��i�K�@Ұa�c�t�p���IJ���]�<p>͊ ���A׬=�ʽu�r_el�3�?b�=�離}��vXn♸&�ۮ�y��_XU�h��^1�@�x�T�@3$Af�]����↾��23<K�U�)��)���}�HR��zY�>�I�ɉQ� I�H��є�������or��nD#]��Dn��均^'�TF I��K��v_�&��e�_fSuH���Q�	 ��
 ��i�J��mr�b�%+Y������\�M�D�}���A��}������B� $�i���@I?g�:� I��~���ȶ2�B�}9)������3�9t��[�8)$		4Ő p� 6&��t=�vz36��&ᴲ^�~�{]$��}�E�C�������o�������y��.���`��H�e����D���-�N���{Ƃ����Ԑ �O��y���O�?� ��@	$�`�xI?�>�&�����|������w	���lS��k���}_���O��|�>?�� �N���ڟG��I����rM6��o>�M���jA���i$�����6��Ϛ����/�|�>��ou���Ԑ �G������/�c��:6$�!#��H ��qVC��Mo[�%־��c���C����x~� $��p7I~�8{����g��g�	����m����!����I?�ٟ����%?/�����M�ʞ�P2� $�o�Yݎ���]�0��|~��m�Oޞ���S�(p��w��|����|E��6����C�������������� 	$�ψ�����g��O]��3i΅?�
w�>�Od	 �M��� I����'.~�*V���3��A��N��<6'����! �M�s١�?i54>��9'��$�I"2lRlp$�������Ѯ����R�?�Ӹj���i���m��AC� I'SA�|���$���H I#�����bA�O�����B��~���v{����{��������X�#�D4>��'���>�������k�{�?��� �O���v�����E�!id�/���0~� $�O�`��3G�������>_�p�C�{�h������7$�)�>xhI��~^�6�	��^to���������s���a�6��'��@I>��>�u���zߎÑ?WD�u=}�w>�����V��ɰa%�}�� ��I�$������S���d���z��I��|a��znO�I��h�,�����S�loQ'�	��I���	�q?�.�p�!N��