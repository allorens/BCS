BZh91AY&SYC�F��/߀`qc���f� ����b�       (    ( 
            �              -� ��f           �                �       P�� U��	�E IIP�%@��@T�J�(I �
AR��*J�E%*�T��R(  $�| ��B�*��D��
�܈����I�* ͨHp�Apr\�)&R��D�ͪ*�9 ����)V���   | �0�1 [�D� �a� rt"���� 4x�B� 	{ 7���X�����J   }J��a@�D��E)H��AJ�@7X�������4��w� �x>���@u����{�/�=�pW�Ǒ�PG��}
| 	'���< 
�� �7������x��� ���j��ҫɧzïFl��R��x����q�*��8�Y�����=k  P{�  bA@�(R�� )�W��)�Ω>�;�ތ5���(r
�ޥH��
n��zҞv4�A޸�]Ƞ�T.�9l.m`   �  6�{� r�ܰ(!�J)pz�.[��U�iـs���zSW�@���ffq���p:$]���  Р�>  ��@��%�	U*�>�h��*R�3H;4w��wp*� ��[�g^@01P{���U�%+:�*��N&���9�   j�  ���E�pz�(��b�����ww �:w H��$��!wwE$��׀@ ��  ��IJBU*�AP(P�{ԕsH[�Q@���ww@CqT%wTw8�.c*�d4R�B�
�Y�*S���  4�  F�1�'��Jw �`G �DEf�D���UIns1QNF���dh>>  �  ���*U      '�h��R &     D�2�J���P      �%Jd�J�4Ɉhb&M � �OT��2M�       H��4�L?�1�O!=&����M�'����|(�����_;���B��MvvL��g\龺�(����~��*���U }�� ��+����C��#���ҧ�UE`�I$��UTW��*~�����|>߻���+�`/���)�1�`���i�v���;b.أ�
퀻b�؁�)�(�v��Gl�6�M�SlLb&ة�*m��0l�v�]���"퀻`�بm�;b�0ClH�M�SlT�6�M�SlD�6��^ػb�0Sl�6�M�lT�v��il�m��`�)�*m�;`�1Cl�v��G� 킻b�؍�]�l@6�Sl� 6��L�X�M�Sl�6�M�l�6��^؛`%0ClP�6��Cl�v��`cQ��@�"��Q�ؠ��(.� �ؠm� ��(+�
+� �� �� �� ����"���`�"���PlGlQGlEGlPll�"퀠`��؂��  r��QlPP�� 
�`�ؠ���� m�`���
��(v�
��b
�m��b.أ��6�l v�M�C�m��`&ؗ!�6��lP�6��L �6�M�Cl������*<��;�h�i_q��5�JP��ON�^��̚���q�uu��Т��r���B�5�y�xi�&�0·!�l�����L�����F$�s���]���`yKh��hT�6�CI;кx�6�˽���̰y���d:4		h�j���4�7V+t%�(f[�p嬴��Uw�Q�~��\��h�u�:R¤��]�7i���o�r��pؒSjS�ٓh��ٔ�ڊd��~V���t'@�2�&��(nj�[�3h�F��GJi�T�S�B+3V8Њ�ڽ�HnV��ʚdۢ�.Q�1K�*򶆡�v��6�/`Xv���^bqn�����ѫ�G�����B;u��k��x�N� �5`a���/*�96J*�J��5���]�JY{����Xw�Ō���V��@/2�X��b֭=s �8h໼t-%�%<m蹵���p��{%*Wq�t�^<�z��DŇ/2�T�Ǘ�*L���q�7�&�W~6X���E�&SB����Z�����.�	y��B���6�k�GCz�
U��u;͔,Z�M�*M�Jdm�l�������~�S�A��L!Ot�<6���CurἘ����5�	�x	�H����`���#hi�7{V����5:z���gN\�޴��m��KW�I�RS���G�+�t���)(c�ְ-����Z���m/Z�K}sN�-�WkAWDV]M��I��57��Y��ջ)]���G��bv�L�E���3+�T4ҭ8sL��[

�
��E�O>-���4]n9Dݷ��+s��-C���ƞ�7kF�wY��݃�V.��JQ������(��Yن�����[���C1�Z��ա��l�^݁�S	uyt�勱v��75�a[/,mQ�Z�a�����r{1�y��oH3��Ddb�+ұ���'�r�-�(Z��)�[��(b4S2�fVeh�Y(����Ħ��7i���k1ś�7���ܤ�d2���3[Ѹ��Y�#����j�b�ML���	[����:v65o(�"��������"yr(d�l�17������n��U�E@������0��62�{�i׌��f]���Zw1�t��2 Y ���P&tP�x�#/|7y(����p���Veir�v�א��2��Cq���A�7����1FJX�V�;�7Hێcӡ�ʹ�1̨լ#_��S[;�lY0�������:��٪ic�Ǻ6d��\����Q05T,@���R�\t����U$(:�1���,�Xq����cV�j��'<(\S�i��t72��(�j�	9�����Z�vC�R��v�����utY�D���M�H�rZ]��+wԴ�{,�H�5^��Y�,�m�"Q��3Fa;�K	m��`Jb����Jc#/d�7+0Y{�Y7BC-����$�*�/���bWB�^�<�J�7U�w��R���	ID^����]���R��.�F�h �Qk74�W��z�[��K��vEC2{Q��������i{�����7�EnG[�r�,�(��+�H�T�Y�Q݁�XH�kf^�j�լ*Xd�]�dJ�)��Hi��������]�gy�i(e:8�1C]�"��,5�1a&\�c���ʙ�-U��kXw���X�rGy��2��7�$���塧,ۡw��jǮ�X�H��#F�d*o4��@#$k4hwx�x��jR�,�`�z�ӯd��&��ڗF(Z*ln�kaڑQ�ͳ��D�4�U��,��m^����ی�n�9��51'��b��b�ܼ�jHv��fV��xJ��Vڠ���ۙ�4.[�Xн�5���oj��ɦ]
�n��7ts�ov���� 4\of*�.�=l�ܰ8E-Ŋc��X���^�9E-�0��.%w��e�x��j*Y�MP�nY�Ui�yRfu�T�Y�dJd$�L�aOMI�!b�#,4�nc�w6�dݽ���^C����*�N��bb�ȑt4U��fQ���:dZQ�T��9f��[C6������U��;		n�P��݁�Z�]�l�zUm�R�c8(���t��Uy�Ϭ�0m��B�ͭ�m�m�F��]���3.D[fȶE=���qj�S]e���X,^&�VX�2OC����Y�i�v�fWkkf�af��Q���Kn�*��X�*�,m]K��/HRn��R�Z�6����/RF�8nݳH�%��m&v�G���.��nV�˙�Б�CD"~���œ��5����.8��xS�E5��c�m\&C���)��C6���)�ɫwC��De�F�=�0��,���x)h�7M��<D&S�����v���j�ڲw2��u�.������n�RU	�[5Vʸ�2M\�O"8�5�5�,����Ň%f�[�yۊ�]�kw	�V������e��Ƴ-P��@�.�.���nؙ��u�{[f�k)R��ӱR	�ځ֡g1=�H�R�;(Qˬ1<+1L2�ǡ^f��b�1��^I��6��R��(��R`�+K&��c�CrVwy�
ӊ��v�/,�%�(�xY˫���TM;��%��^'q뛶7H�`f�ѡ����r�[�׺��V�43L�יF%�n�E��TF,�Ut��بt@b�	^0�����Q�ա'�����q7�a�GdP�0�irŶ��Պ�Tc֙ŗ��cڵyulͭ�˵�[�K-�tT�:f�[5U��r�+*0k\L�2)��u����[e�V�Mb7y3@Q!1DF=�!�U�#R���M�lfl��w#Z��h�fV���CM�VƳY���ux6�애V
�y~�r��H3E��M֠�@�t^��řl�"o�`ޢP�#Py��5��i���I�GsHz����3q<���u2��єl٫%]@�Qu]K�e��g�upa-{v�yx�-	����+[�V�C#�er9�/hT"�ۘe�7^z���{S�j�9�jxm�@�Sv�<�r�÷Qiu��
A劷��/lMZ6/�+.�X�{�:*��w���3&�n`�wNٸ�U�26o0�z�݋��.��ZP�V�����+ׅ��%XydM��52Z)�Zj����w�����lU���tM$�n���=qL�W��!i��Xe#F-�oI[����W-��+*�h;5E���N���Vf&1����X!�C7�8���*��xd�97n�)�Qn�7��K3�n�R�N�!�w��ܳ�m�.�����&X^=�~2�Ы���;W��N�E�j`�W�]�� �f#z�x��ł�[����sR˸���Jɥb�̲���Q�ʒ[�C�$e��i��wL�.b�a1J�k�y��or����kr�]p���ţ��a��u��������Ď�
g){&V�EiY7Hё�i�N�0�0n�医�����N�Yckl`�ӋL&-hp���*�#�e���1Xp�x���V���j^+43=�*z�gD��S���։��VQw{��xf��3!����!�L�j�����]]`Xa���0b�b-9w�Q&P�n�l�zr�P�#Y���>�����X��7n�a�y�C
�r�@iU��8�ItF�))X�^/nj�������KE�G2nݼ�"�;����$��6Hh3-�ZW����6�,��xѰS�#1�y�A�T�c�vo	U���0e%z&���7���z6E�Q�ťff��{rP��ד}uw)�*ML���O
�[�)�%�@�*�1�f*��	��X��l��R�+77�J�`���J4Sӈ6ۤ�Q@^*�'Ӓ��J�6fa�ø.�V��p���e�[X3fbۅ�[K2�V�t��j+B2�) �V���sc��j�<�F)�n���t�3a�Owb����m=�˖�+%�ܖ���͛yN�K��sh-��&��Ucv�;N����V�6��*ȱ�uڇuŻW�fmdݕ{N��9�D��͕(��k6niH!n�>Zٔ�ڽ��nj8'.֨/h�[��m�&�f�9��7<�̃DU��L�W(l��m�

����Zl3kl��Y9D���OE�x�m�2�Q�T��,֓'l�I�F�]Cn.�Q���T�bj�{��^�h�$�rfP۬�뫴���TB�)�W,�Z�aP� �b��^Zq�p�ā�yX�m3D��
͌R�휢%��j���]U�P�Y+6e��r�9�LY�]V�/ �͸4�<0A=O��2QR%�*�+��-ڄ�V�[f���8i^f��9K�n�4Z9�P^
���J�N�^����V�WvC��YJ��b�%�B�n��u4�n�)m�(�G*����q�N�	��&�K.�r�0ރ#��[KJm8�0��+3؆������u�B�Z'�ʆ��lص�73t��X�s]5���Ǫ��UwWW�]#W�����(�u�M�ʭ�Ehut��a�l��P�)��5*�^2#���F�1�LJ����ZڣeLӍ������p+��ꞼB#V"D��}�d�ĥy�r��`a	X4q�d��1�^n��o�D��n-���\����Ŵ-xl���&^cw��42��q��YB��Ygn�(W��P�3�%��v��z�n�Q壗��i�,�֪�r�bW��e�N��;p�K8c	ٽO"6�1�eǑJ�$�ڑ�^:G�DkqeY�*L{H�{/�S �aPUe��/�2�ɧ2�sn���z/�h�xlF�u�%��-�Y�����*C��^m�ik٢г�F�u�v'�˽[j��(�sv#���(���DƓ�t����gn�FŮ��+rC�~:#�m�n�k�)�0����J:[ܣgD��Y�P��e���Q��h����ݓ[��r�e�n�sv��q�@�9%���C���ʶ�Ȏ÷!�x��řN ��-�6�etF��щ��F��ĥ�S�cY�^ݚ��M��`�	��4]/]7�d�DsڞL�F��cV*�^X6�xȆ��$.�'O/��i r@��YZ�L�{�(���m�w�h����t��0��±�YR��ݍ���z�t�j�۳�p�+1�Mf�^��(᥸KڽֵK�����znd[Q�fkos6�YN��xn*
�F��<� b!�*۰N!�����p���B�Q�x�v���P�ei�Y���]f����e�Ȯ�ڧw�x���H�g%,j� �X���
��u�$��R^��un%�ɗM�SFǱ���2�+2�U��W�F���g*R�h���l�khŃfnAa�K!�۹��q�*��$�d���2�	���ܻ����Yf�����l�Wz�T�M�Z�'�a��[M�YN�5m�OUQ(�Pm3%1��k72�.��E	w�MK"V�)�K�5`d�� /{�}2d�\oK������T��K�@n� �0N1V��ÕuV���HX���@�9��ч-z�ɳv-;A�[��n��M7�V�U���N��~�Xu����-�q�o'kq�������v��]`v�n�T
�V3Y�+76�X�9�D5D�,%osud(fHkd `�b��a�1:b�s�X4�@�h��o6�K�"�L�8p{Z\҂#*n�Z��ҭ'w�O)m�d7�,[�, H��7]���0)��bRcoq�X]��im۱*�<������m�����B)�W��V*�@G�LE@ū�E��nn��c]�n?���!+Gi�b3�\@�ʐ�l���V�u�v�b��Fl�o=�f�k#M�	<9A�a���e׌^q�v(Y��la�i	U*+j�F�ԑ�$h������R��V�r:�k���yd4�dK/Sݿ"le๳i��c����V^����;vU=�NXԯI��,�,ɥe=�q	o�3��d,Y��jf�vf*CZh�N5�Z�w���"�d�z��]����0)16��Wy�ӛdwc��@S\X�3eӲm��v8e�5P��c	x���CX�2�M��M֤��[x�M�c�X$Vdݻ�!�S�D��s(a�0��Q5gr�i�z�^���h\qޫ�MA� +�b���}�&��f���G{���sH���k1nc`k�h���L'q���q� Be�[��s`���6A�	��HnYeBjj[W�r��%�v�e'J����uvMvYi cX:��wV�P��%X�-�3sj�j�0\��[�3m���SjU�X�T4�ݠr�K&7mk���)Z�F
��镶�h�qL�0���fPj*���wl�k6X����kjfT ��Y�8�ժ�������h8�^�
؈O_��a:!4���N�f���Pj�+*Y[X��ͣa�OA:Y&��f���v���$.m �.^��P�nP;���u,Ŵ���N=B�L��uk�ɫ������uf�n��������Wx��EA�z�6���i��ve���*��>ݣ����NV����@�;�a��@vd4��JɵxsnQ���@z<z.���.C"�֥�aW��	��h)�zM����
��q��b�b$V�ʅ��Y����R<̍U�j�ŷ����pm-���<�2��e-r�Sf�]�W{ec����$6�q�Z�g@�6�+�1GSjس2%$
d��H���[������{st��5u2���d1��<ܻ�ސQr�ޜ�'+od�{J��V@󋫲���������q�&#��̛Z��]L��wl�l�[Zls���^�K�C(ۛ�`	fѸc��n�΂d�͛C�m�L��6��=���s0���ۻZ���)�_X��yn7��6�l�A
��0]��7�+*�%<wy�����䀛:mݝ(�L��CQ�ܼ�D#
��;:���O�PD����9f�r�g��i�Zwf�JJoC�,��4kcy@n�or�7)�<Y���%rq���Ca�y	���W
��n������9���<y��I�a[�yh���AD$��m��m�V-m�b�m�m�Z���U�T[kj�UV*����kc[[�Em�UlVű��F�E�c[X��c[b�m��m�-��Z�m�mQ���kX�kkF�Z��֋m���ZūE�cmc[m�Tj�ƶ��U�-��U�km��[�*�UF�X��֪*ضִm���V��j*��ƶ�M���X��cjѶ�M[b���m��bڨ�Z���mV5��Z���U���,UZ��E����j�m��ժ6-jŵ�Z֑DA$A@G|W��UʜpK��^s���&�mqn�:)���#��1aE]�yyW��`a�I�r��g�U�.��-�_6�t(*e*�Ԩ[U[����l����K\д�\
�� ߎL��e��[,�
�(�-m�
2�C-U��.˥�d�����(�<IJ\��ߎ���Ԯb~�EE�{O����� �g���|�S����ǤA�D���z��{�|�������R�yW���{]���U�j�r嫱.�U�;��{om��kJ�Ի��Y�0\}���X�u����n��ۊ�c�q��1�0�
b�[{N �n�pqy�4� .��&��S���\%jݺ6:�&��IE��ZCD8m
[�� �f����o�����n'�) -u��i�X��[�ޥ�fT�c����>�����m��]��&s��Xo�u_0�R{�*�Wu�)�X�Ycs�3�7�����%���;�X�V�k� uG�V���3��w+���ئ�f��sE̠��.� �s�)�+��:˳�d�y���,��������Yyd�6��J�+�nRj�i�.ś��N��X��[��u��gj��:�uk��U���;�A�Q
�2km�4���a�2.>ہ��u��t�e\��
ޅd�mv�sSz��)�V�<n�bӡXl*W!yx��)X���{}�oU�ź�W=����:����v6U���Z3x�kM��ܰsÉ|��Ɩz���{/,v�5�ي�ҽ�D�+�-�Ă�y-9F�Z����ʚ�e�%�����vU�-��e���d�2�ۡ��Y���v��h�%�r$����xD���L�+E˸�8�-;��kNi'�ĝ"�'��$�u1����.�w1U��iWcs8hw��n���K1�@�yV�q��o�Vd�q�d�8_	b���&�ɰ\
��p�/�r�U����cc�{]�0��׏'P�R殶%�&�Q�H�ܴץWm�]^�iSi�6e�����Q[6[�f�K�-s��\��&i8	V�5�/8c�'b��[�n�Y��3K��:��Y�(���a�Y�"g�u^X=@��u}pW�H����t90�ȝ
Gw��K�2��˜����
Y�������_`u};r�;	��Ƕ��-=әN��U�vê��rjOL��6'uԢGV`�8��R�Z2f��w,���.�̽W�5�|�X�0Fᶠj�x��P<���{j]v{V��g�PkZx����t�����u�eM��N�iU���a�6�2�U�g�r�WF�9��أ�,�x�D�����k�m�g<k�V�޼��1��+��X���Bb�HV�o����t��ס>���� �Wq*��^����}��K�`�X׷idB�%L��a4M�b�S��.W!ۼ۾˅���WP֊���q�c0ַWʕ���qu��s(=�}Z�:���P�������9�9q�]��]�����QC+8�'k�/���1��H��l�3����tmJd�4m
�k+oלصniƥ;Y�̢�x���y�}f�;�fx���u�B+�b���'c��J$x�InuX�3*4bSd�ݍ���o�w,76�ޮ֍&+7+���s�ě���)�.�sὉ�yk��˅�|B�ft�.�C�z]�t�]�x��6���,�{�/��X\P�H潼��mMx���g`d n%
yY�������a7H�qnjR�����V+e
B$�CYt7tU�ՙ�䛹׷���ǝ����e*h-Yg�ob��E�{�F�$V���CTB�L��=���nŎX7Qz�CZ9LwJM��Q+7�S/��Jt�R�n�u��U���8�v��x���m&ifs���J�Y.�v����#�śn��CS�o+���ųi��7�}o���s�c���<��1��üz6����T�5��.�L��^�X���&��N�2�\��W�g.���L33u��g���<��eo^��V�Z�<AEV`������:��%���F�r��$c���h���7hs��F�7�th5ƳD�̗ov�᎚K�sAS�'zB�m��;�¥[�瘹KEV�5�:+ܖM��^��v�曵���n�@���)R�ɓ����_X�lJ�����SH\�� \%L�����wW[�L�����"�F���WΛ�c����dT�K)VV'W���w����А��k�w�)wQ�(>���gTK�i��9���m�B�E��Ik����6�0��%0�:
���8]��v�JqV�5���EbV������;שf��[�V��K{�%;���'�(D5r/	2��|�:+��8�^w1�r�;L��[�&7�E�c�0�P�ʥ~F�U5}8�"ؑ���� D�z�b.^̹�X֨���V&l/���%����de�9�۳#�z��kÊxC�w�Yt�^��;�R�Rˌ�,Tk��ry�:]��u�bH93=��;��ܫ��_㛆���-viy|���!�PGEUJݮ��7���Z�[8�%I[9*x��Uҿ�Z��v_q��/�#�P��(Z�5�/2��M�Q7h۲ف�"�Nuz�q�;��BoU��ے�)4���b�.����г2κ��h+k0a�H��|�rf�������ζz�]���g3�6w3�eؕi7m�:����)·T;x���V�ۯ/rҡ�N�]�խ:����e��v�k !w�	]�iZ���&[���$U�u����(;�o_|�d�kۍ�Ť����$єU�ܽ�` �ئ��^�;'�f%u�+2�Q\�����gnL�5�P��xK�Z<C/v���U�.�_��0+F�Bniuw�\O. ���Bk����j�v���]]��ٗơHgh����Xj���2�P�9�=�t���+ȣ\��4^bA�{�v��r!֭��pd�nޫ�Y���������i�{��a��E�l_�⹙��u:���E��Y��u�]����WR����Z5��c*c5��sn�.���w�P��Eٱj��,�N�p�/o�W\�Vێͨ;-S�6��vOM��8��`��!B%t숺��Pd���5���X��nҧ�fٌ�]��Owi�fW�zx����(-���E�1+`�WL�G����-����k2p��wk�F�&�ԡ�A:U�Z�ŀ!�x*��E|{�{)����PFnT=9�Kw��mWd.����ٽz�P����W~tըn���3/�v�����{ۭ]s�=�E�
㧶�ڮ��1�ʶX�m��]y�}r�!D�5���<���p w{o��kI	Л�\�ݒ�O�8u��/R!ь\r��%��V_!X������\������݌��u�V('X�wL�h�����,,�0�Pi�=����Z�DF_P�OZ3����`��7k����KP�Q�-I*Y�۞:�EڴM��
�4�z��u2�e�kh:j�
�ǡP�����%��k&	b����| V�reWyz,��z{�y7[��V��i��{K��֚��Y\��Y�*v�u��6�n�Mˉ���j�}A�f�E�g�U�h�ϳj��ٶ6nd����[�i�1�C���f�&�w	[��E\��Q�ųUD�#�:�f�un��ެ� �p��ۡ�8��MR���%:��A�}{�e��hU�n���t&�T6)w�d0쭚n�b����ۥ�\}�E��ut��GPm1����2	uG��w�j����+bnn�5��SNI��JTkԲu�E��]��3����E��ݧ+7��S�}�jv���e����)�h�9c<�!r����N�@̕������PY:w:��l7z�Jy/�)c�ԗ4��pq�\��pЇb�Gxq�Mp������[A]V�lλ12�gv�G�gL�I�7����2����X�꺘�k<:�� �S)t��-���w���cX���ۮ�Ah���S�oe`�pl��8]� U�i�^mbΧZFؗ�},et�'m�IYե=�4E�R��h��wV�B�#J���h	���n�q
7.��y�ke�w`;7Ҹ��H�q����}f�d��ۨ���M�M���T�/n��]�$P�qK���hlVu�e�k��g�4p��n�	� g7{w�k#��Hxp����X�;|��j�ח[7t��^�rғ�I7vJ�vcR���hz��[ph�.�`�tvv%Q5����c%#���-��ל���@5K$�p��yq�jy�l���9���҂�}W��6�P&P�t�e����67,�e�o��̻{��*[N�kr^��k��J\�(�o�]��92��,�����:]��ӝ%�]�.����J�;Uy��R��Ӛ��-�|�p�,G����V�����Azvj\�5 �\f�yőSei�����*S8�,��w]�Z.�$1漙���j�:}7�m�Vǭ�;�\�,0K۠�jۀi��{����HT�s�F�w�{:M�%9��kn7�}�_2��s�<��m^W���A۵��M�qn��+���`��o/2��8�y��T:fD�{*Q��{�����狭FA�ԉt2�
11���8�:�b�鲶J�Õ�h��}�Z�T�s,�x{)��׻vW{��d��s��R��$�ۗ���p��OJ��k�Ě�[\��맣�NJ��8����sw@�OU���mr��n�W�W�J���1�1Z�o��L�-	m�d�6�t�(sHi���Vk���Y���YL@������Y�ܟ[���͚^�����w����P�Y�����:�bj��I��4���<s2�J�:u��6EjY�nX��{�0L�6��I�F)�]/fZc���6���)-�,[u\G�4/r��ə�3�֊v<v�$�R
wԗ:�k�물��m	�P�c0S�Lf�I�������z�mi�O,�5�3�	\�9յ�}b9%���	�����������X$I[U�8�B�ݪ(-��ӊ�Uy(��S�/K����z��������3ft+.��^���]q>]CnS�ػ>��1YU�x�r���ۅ	qʹ�n]��@R�����(�a�2"�	�����6zŞ���bHg*��f�M� �ucU�:.:�U�S�Ms[ǜ�A�&�cse��j�L�K,-}w���v��Җ���dE��+M���K�.�Ε��v�]��J�]ɂq��㣖w�e��[���Y:�K��:m��"^d�#_f4x��t1���[V;6S�]%)=;���ä�U*�icb�.�B�ͩ����w<�wc��
�[�]r������~5����^�E,�j�.��Y�9�/�-�6�Y���N�(�*PBfZ/�dJNО��C�u�hZw�� �v�n�Ւ<ީj��s�/&	���-ů/�; �wFf���#6�s�w^��z��#ט����P�[e����< �y{6��x�3B[����ңh�<���V��i�۫�omF��=S��f��R�*k"�S\����(.#Bc�Ƹ^6���'8`���|8���,^��SOw k*�������^Y��Q56�It�8���\gi�K1v 3�S�ݵݽI�@��N��I�4���e��l�K�`h�+o��r�M%1��8��S��Xق����{K+cĵmy�*�����&��P���)T��kSH�-Px�"�m��[�.��j��]J����:��j��\h7�ՙ��>HX��fdÓ�N��w��]�h��%�������T��u8�{�ed�}��r�Y!��YO�fY�Ɩ��͇��MK.���y�`��nFk2��y97s�u���+���T×H��B���5ĕݨKɽLo���_��݊Z�n`SGr���ڕיP�ݦ(�6��sAV�f[:o��x^�;&�g)�� M�J��[�0�t�1�3�[����)(66�/N�@;b�A��X��+HK(�<��W������1��X 7Õ�]�:j���2���KE��3�k2������u::*���ޚ���r�1q��7��)n��R�۶�ۢ�ڷx��9>X����d�l_l���um��E�Ȼڗ[��ۺ: u��ظ^�n��f�ֵX(��w1�%_Eu��Y��i��+���w�~��Wu���`n=휺켘�h�a8kmd�
���{�Wci{53bc2�(Z��7��h΀�uݮ��t���q��\��ؐ=*\�Vp%]NA�����]�oQ���2�ͬ85�T��Y�1Wm3YF��V:E1����m�z�8!�m�u�l���+����dO7)G�2��$�����o��F���u�52�x%�����
H.|'gJ���}+_U�G\���ݛ�A�cA�$ތ����>V4e�ul������r����-�]jd�9���ٹ��(n�p^Yw�R��ܙ}Zs�����5z/����C��K3,�t��<;R���CH#�uM�<��&�!x��m���/��~��6��(�,�8��Y��ջ/�gA�BnND {&]iU���J,�;ˏ�i!|s��Y����WNˣg�
��v�N��U�9�n�]5Vp�#9W!���У�{P���wX�ʽ�5��cg�^ۡE#Q��S%Y��`��:���c˫��-��6�,+Υ��f�>�_��&Ggv�b�5�!k8��^�2V�q���]�]�G.��Y�r���$\�/���:7���L��(����	����]�����an掮
�ls� �w�sMZ*d��h,��'u.�fh�"X�iĩ8�[���Cy<;����$���r��;X��:�t�XJ�)�l�:�v6R����CO�\9�rS����נC�U��e[�졷���m�]-��E�!�n���_����7�x�j�����4���-�����e����Գtn�\�.�]��s�7EL��y�4�NT:G�TT*f�P����li�;:�$%\TT5�_@t�D7�U��5=�%g^�k4��Z;	��Z�kp�wg&�<ŭd$k�Z�R����875�o.ر�`��6���W��y��������?Ծ� >#�~/��?�����8�=?�����*]�d��*q/�y��LD�5X%���y�t.���f�ڣbM{V���{,5%U۩�ny�q�pO\l&l׳�6n����t�n4t몶��Qc�k�[x��4H��3�����b��:M��>���n�p����Vw��ŝ�(�s{Y��pq.��Zw'��pש+��n:-,#��p4���ˎn���+c��Dx��A�!-�f���w��q�[?`�r<�c9A��jn�m�&��4ЄVR�Qە6i�il��U������,��NWs�M�|�m��%�Gq�a�\%�(\om=cpzhz�t��/��(�7��E���ۨ���6�-��o<:���ƉT���7���9M�(�Z�6�
��]��j��Е��]�.2i]�pk��N��uU������U�ƻj�^��Z;pVS��7L	����n�ւZ����T�E������pq��g:�bxΧ�7<rs�� X4a0*e�����.L:h��fx�^���+�k�1䶉mظa��5�l1�MGir^֮�(�FT���a
���%�Pu�Q��SJ�v^- Ƈ�<٧�Wi��F��� �8�^%q�lG7e�Q�1���M�Gi���x,�hyc`j]�oQ�hn�l�=�>nٽ��r;���u�	@��E�U��#�EV:�tszu���y�S�l�st�L`��&l��g��݉r�/l,䒋ٲ3��m�rn�IY%��a}mm�ZL�
J�V���e�[,�����[�C���3s��]��:�cM�o��Nc��BN��ƙc��Yc��W&�d�s���|�<�a�\S�%�ШF�ԡlc�j��#�F`B9�p{�,g�%�Y���y۫��F�&Ë��8;(�	�p���Yf����d������mn
��÷���6�v9m��a��a,ZM;�N����mx�:��� �1	�l�Vi�W��-��������x��\�xjf�.ޘԙv��me�5� ��s�ݛ�E��ٺ�[�GT=���p��]�����2�=����:��y�&�m��+��,zu��6�A�0�r���r�6�g`S<q�֢q�n�����.p���ȒL!����Q����óHU��Mq��&s���Z.���t��{/c`�����6)��<w7����
݃B�f��ۍu��Hb9��k�r>��x��v�=P�z��g�m�l3�B��M6.v�XR c0��,
��3]MP��O��pr����ø`pC��[Mq��[<���ջ.��豮��nt�H���k�k�&[���m�6�<A��a^T/�<�6�gvuWY��k�7bѴ��,��\:SkW,��'�����B��S$-1@(d��sո�\=�wXv�����AU������c�Ǭ�sl� �=7[��2%�t����Jf.�����B;g��n-�]H[1珚R4�ai��v&��TN�<]��t�ØSVU1)*b�[0������[CpN�ToÛN�H�n3�z�Ɣ�yܭ��y�֏	6ta��k=��t�n��II�Y�mMv�s��oX�&��j�F�i�8�:X7AV���9�;d�8xũb� L�L١c����6�:����nL�R1sV��|'[���z�'MKRK��;�M��РR(Z�ec�iP��lN(6�6�����t��-�������\JĆs,IePk�{6�mM�E��77d���q�UE=���z:,m^��ɵ����tnuص��l��M�϶��D/2z�b��g	�nJ�/�K�;���ݵ�.�vV�A�w3��,�g%��!�W*�HB=G������4�3�쫒LSP�gT�~3���1��[f*cA����jԒ�a�5f��5P⮌��':y{Zgd�f;ʚ��9}̡�ÆM��7vO\�{�W)�^�\�D�0nݻ�x3q&��ԃ �ώ��<p���8��m�8ٚ��pvV�ܤVܾ�qmι�{rZ]��v�|�`�qX�&ږ�s��.���=i9[�]n6b��6wP�ڙH��	��Sk�%�{n�ħljBc�5�77�ڶ�`�Br=� �̡�X
+=��o�cZ��ZF�٘�7B��1|~��{�<�nې#�\�LF�h���s�ڋ�dݴڈ�-��`�\���6�]���c���73KFFXKvGk-�����@9��3�n{T������+v�����k�0���X�=kW<v��-AJ�<��:9�`��]I�q�����k�yӐy�$H�Y+z�}��:��t�`A�	t-�mxy5˴BYb;Z"Z�f�԰�]
�<�x��1��zr�&�`ձs�l�@�I��jV#Bu�V�y1�f�)���5�Z����r����2�&1���gXx�#p�����s���7��͎��y�,x5���4lƭ2�,�+���mX�,.�H,Q�n�<�ҹ�:���cc<8(��q��l�uqc��5뎩��-��`��'Z��<�U�1�B:�{j�b���f�
#���F���l��cC��\��ug8��6,�^�n������W*�=u�8Q�mN�q@ڂ�����;�li��%a�fV2��������>{Us��Җc1۪2ϜE��9����ugq���ֳ�tu�Nݞ�lv��q����ri�i<S��z�CgpX0]B�(�k5)6r��˺��'S����x����+hKL:����K��n]n�ݶ���B7���t	�����[�ժ�\�9�KǨCc�=��N��5�b����ʹ�������wEٻ8��۱ղ\nz�I�K�:�M�5:6�t׮.8q�9���W���Q��b����R�t#mq&��#2�+����&�ClTM��.�&�׈���ݎX�-��V�u�M�$֜^z�;r����eظ�j��u��C6���]B���^6�3�J�jݲr;o�ys�XM*��g1�,� HnР��bUR>���ٸ$�3�pv���M�I�q�fhVm��d4������ۇ�<Oq��q���	�G�a�� v�R����M���Ij���<��d�ܮ:9w%؈Nwc�]ړ"�����꼽E�Hݵ�색�̋���#�͕Z�ʘO)�R4�>�9���l!�-]tR�G]Wch_����2�����9�Eۃ��1�\��7i$˶���r��jB+v=�M�J�n�l�q�m��b;ׇb���[���+�H��{nҺX��J��T-n��v)�m�� n;��B������
�B̙�b+�Ji��H�����؅�\zv˺��u�\x'v6�����9�g�����k�[V#XA�(F\Q=���h���]���F:�TwQ=F`pU7i���絚�SG�.���Gm����u�3XL�B\�n%-¬1X����\,f�a�om=��һ������f��� X��CB�ispk�۠atH���&�Yx�=[���3P��L#0�"F]s��tb7U���S��f)�%6�湒���8�pۢQ3,��]4��P�]	��ĝ��;b��s�h27cN�{���� �Xծ�4��ZZ릁- ]\Aݐ�k\��=�����9J�R�%�Y*K�Ϛ����;^ї�.t������X�69�ͺ�8L�c�r0��CĆ+3mʹ;v��A(<�S
)-O7nM��gN�z3�U�k��A=��ݱ踆���r�F_���͵���Q��5��Z�B�^�-J�N�RV��Қ*h�:`�����r[��gW��u�b���0v�h�CH�C��ޭ�U6��n\n=v.��0�����l�Rg��)�+
�봖k�D3J���$Vɫ[f�md�]��#�:�qC���:�6y+S��v�aaʽnAW��q��4���-9�[���F͕0Z5�]��kE�U�	cj���==�p�
˴��ܼ�{,Y��m���b�8�q��Ԟv˺㋋�o0��D�Ɲ{dMm�ciG[)p��{Cf9��s�L�X�s�ouu�Fe68vu�a��1L(ʛB��8BjklъB۹���7�3��5�\lV8�/ж��D�ҔYL�ݱ� �v�9^z{I_+����Q�A�	�p`���^k��d4wSe������\Gv�������x�s��2���8�����u�[��s���̮s���N���Nnx�eS�h򫦍٘��@�xA��֯S�$�ܫ���7t�=�x��je��+���"n�n�kj�{0h��h�:y�]�����qO��9絑혹`����í�������On7R]�ͮ�X�W d�.x������!.붬ûa{��C��ăv�apBnxm`�A�4k�d�c�nn}�g�n{C�����#m�"=]ۃ����6S�ϗ��ϧ2N�M՘�ۜhe������!���{a�Iy]�E�m�� �۩ǰ�[k�t�=^����n���t��kEc��ֳ���y��:�gr���NX���`�[����wǤ���]\�.x-X=w/��n�7ܺO7H����Q�eg�Yce�mXyw��GŲ�ЖR�ǈ���3��-F��gۯiX���>{�=7p�Q�cu�v���ݒ���h�1��qv�Tl�k�NJNJ�Mk!=v�u�z۪�`[�m]p�u��ݖ$�;ժ5#t;v�n���*B��e�\]�b���`[Ha�enյ��8zkt(D�;F�&14�M�2�v\��g�s�W;A���0�7m�gY;0ns�nB맒�#܍���#C�ܺ\ˡv�ą��k��D�I�Hz�RYn%D�d+.�A��|��ynGmF��&�y�5��PEr��EE��sTcDQ� j&M*�7^륐��-��E����F"�Ҽ��]�%��uy�k����b7�Q��s^sl�\�!-�vQF��So��EA�ѳ��-��1�llj5�]�&5��Uͨ�髕w]$��Ǜ����ͼ+���m<�˖ŗ�w��M�7+��[�hК1�$�y�州�d,��wsշ��_���Npn��m3�tް�M����km�;G�5�N���8.�iMmW��V(�T,���"��&�@د7Lr!�x�Ѭ��7c��'V������&5(�1ka��0�I��n���0q�0�]	�wϐz���f��i�%��U�$��싗�Y���hx�K�m�;sl�p�����r��u��8'��١�q�@��;<A��U��f�1�1��n�%G�{q�;���A-6�+4�`����,�"D�Vņ�GeL\]Y�P�c�{/nz�:�Z�[V�U#@T�.e7&�xw`jz;���L���b�xs��5��gOK^G�d��ەሚ�W�&'�q��í�Mg�P����c@���#��VO5Ԏ�c]���#�]��V+v������o+�x�4�+.��΂p�v^.�leqͅZ��j:cm,l�"���2����a	KQ[Nh]�hB���LQ�4�B%R��͸-IIR���g�6fkД����A3]�r�X�Å�\�X���-�)�v5��N|m�����I#y�l5KƮ�:���V�^ϫ��.cMe���H�;��ôU���yx��[Zخ�n-ݠ�]����%�����J�޳���.9���Q��v8�]�L`���d6�[^:k4f*�-��0�b�c��4���r��]���+jq6v����� ��]���6��K^6����J�hr�un�Lwl���6ݔ�xfjk�e�5�D��VR�F��I-e���W��!�����4�c��rO�O\�6�����.���	����ꛓ�b�]E�e�;۴�j�P�.4,1*���q�"�4����[:�������۩��Y7gn���qɲ��v0ٽhs6!,A��^������)㵤N"��UZ����7	�s���͛���ࣣNٺ.��5/m\6�upQ��z��ޝ���~�<���2�F���lyJ��J�
4�z���BR6J6R5KE�G��-��ca^�4�+y����^�	b�������XT����F{!,m���6�N6yx�8G�����`�[+%%`�����[Պ�H�� ��Q���m��Z�i#*,��ZQ��M�jI5��r�O�u�����κ��8�L���s3�n�!����X�'�I�e��q�(�Vu�q�2���ͪ�k4��"�Hh~��m���/w�+3��<���+�ͅXs:�]0��]����$�K,��~X|���UR>����z���K�����>��J��~�����~���ؤ>�$�U��3ओGV�ϫ�T�o퓾�~v�]{�?��^�~�ۿ'��[�/g���H�k�жgd��(�35��#Ui��jue^Ǳ/.�/�9�̵����tw*}B��"�%�1 �YӞ�$�gky����qs�p���vy�|cS�l��]ۊiӻ�U�ņ1\�F���?V�lv�<U�j�C$^�{4_���J)�q����υÊ���G(�n��E0sf�ə#�2VSN���Ҧ�ݵOGn�F�K&x�6Л.�v1����8�kl�Ŭv%��%,���x)Ć���vVW�d��a;_���ᮇ�ER��f��]<�H�e}��qn:;>��v/N;����u<�����]���n�+�1�b�Z&�k���;���/b�L7�٬�RO����***δY�k7�%���e��,���7�z�C��O���d.F��yI4�S�.j�R�{b,��ܽ=`�Y�`Xe�v���Mm�G�1m�J����$핛Cr2����ܙ�y�{~��uU����2�"��(A&ݽp���VT������J�h��NZ������=�}�ڽ�j�#�I�ܮ�����v������Ƿ@�}anY��Y�He�h��#wi8��-#�ڟ.'M��Eoɤ�j�튳A].JP����(5&N��J�y�^^�qR����T��>�/zC_Gv.�ۣ�o�z��L.̭AJ��9����^�b`c��tZ.�1��|���p�]������g]���ӥ�����=�w���a�Ϸv䲯��ͮ�G��4Ke&B�E��W�҃�X�4��M��t�m�´�5����H�����`�ZY�����T��-����(�����R��_|j����/F���}�G���n��>�|;;X��}˳���:}�Q�@�*hF�3�9j1E[�𚊪IT����������G~��rw'�2�]7���8�`3]ٔIP)��	�ؙ-ᙏ���N�KvE�Z��a;ֆ�<U���U�-H�F�Ӫj2��A�����ɯf�l�+u����\��*i:�&w�N����H<��6#�P�UvE!����U�:+�_x��_�>��w[oݦ����z�R���V�����,J��%��c.�(����s��YD�M�n�)��]�۝+��޼�׳�����+��܈[���m&Z3f�4�,��j��*�2"� Y�O3�/��K��p��٬ķ]�N+Id���E�������~;{��v�__GRI.@7mMWr.���S����pv�[�ܣ��Q��H}t*X×�ox��.�����E酪���l�w7N�0��r݃�[[�&�$��&�MwmHi�V���+/V�>ԉ�I,���]��wg�ՈJ��������W��qL7�u��Q�Vu�&����-f��3`�ra��.ɻ�.�W8Ucw1V⭜gp����\[a٭�s~B��P|��H��25sch��8���#�l����d�9p���ط��<�1��:EhM�����"f�z	N���+����2��i��ۙ��-�sl$5�uv�1�h[H�jͼ��#u�M����e��gV��4�blc��a�t`t���uvS]��P��T�M�XL�{F��C�u�Œyn׵��e���xv.,���~~}��Β��4��ّś��m]n���3	,Xh;SG��v.n����F�5��ֵ)	0O��'Ƚ��YL�-�4�����@F�K^���צER�˥�VO�^]\�k���W�I2����j�p��M�m8�
Iǫ�lݸ����Z�m>w���u�dFe*Y&/j�����T�?H�����!A�5�*�>������O�oa]����}��u���x�Z�s�T�E&l=uy&	[&�c,9�f�N��X����^d�$�}!��U!��1�]p��F�N�Ea&�WL�uŮ׃`6���;�s[�[nf���Sa��w4��E���b����+1n���foX���Q�΢0g�����*�T����IL�>A�Ux��Q�4�UAWIb�8��_�&U���%<��u�O80�1N�]��f��r��ƛ��>v�1����__'���W�d㴔,����YMG��[]�	M��Rp-�k�}�*�C�#�!;�6������~��;��iߪCU}/�g�1$����MD��9��`��O�NV���2b�Y&ob-�Ɲ���b�p]0�׻o"��"�sC1��ɁYu@36��m��^��oa}��{�TȤU/q�|�x�Y�r�h6�-q�� m6����l5�4s�B�ź��D��)���ު��Hj��>�|e��tN��R-}Օ�f}�U�Ԓ�nٌ�)�3\ֲj������[�pFl�O�id������������u�)j�C^����_�ʭF{tkm�{�ƾ����l�fg�ݩԩQ0�H�KN���*pd�>�H4���"�nY<q���V���ȹi�J����+V�t:���;ϥ�����_`���Q�C$�I��z����
y�K�ݜ������k�t��w���R��Z��e����ZMH}�"��C�'=���
[r�����w��j�{�����U��CU$C���~����<�!�ÑIp:���PD�۞0ϠBϤ��=�٤�n���D�C"�!ݯ��%
���2���mfY���E���0��>�5�*���>�)����S+�n�zs��c5�ܬ�ɕx�}v�wX��[�]��8�Uk�].��!�*�8U�����Y��{-�!=�F&��O�[��}�AJUx��b��kP
���x]��S+Y1�m�e��8���z&o}���>�!+�8�N���G�b��{�:��|��wv��-}��M��_]'�A:*�3j4�Z��aEi0/v,i4o�锳2ˏ�o��|d�/z��2a�����ړ�b�f���̩W��z��_ERT�1����(�%� �9���{�4/)���i�{y�;EùXm�q�dy��ñ�����X�]��퀕[�����f^�y���ڷrH�Ӿ�����\�w�W�S9Q'ej{{m��of6��+̝���bj�;G��C�dGoM�s��鎳Mv��.�x��Ami��x��mLՔj�ƅ���R�o��N[��l�Db���H�M4�z��n�fF�PP�bS�Z")�{�����u�}}��[�ۧۺ�5ȅ��'�R�k,ݛ[)bk�8�{,��2E�d����w@��@�yt~*X���?�S�Ms�shDXhU��`��̼z2�8��-�c�'��=�?U�׵��U�h>���5z�vPu\|���_C�yp�����Q� V_�7ʮ�Ǭm��特��١�Il�\:��l���5�1�{D�1���� �1�m5-6n E4,]��,�����q��9ֻ͇K��fP�κ;p��\�+�lܓy6�.�녶��YW��w`.��l�Yļs7b����c���ݍF%�5�k���!ۄ���v���ظ��@[0r9uu�:<h8�����g��m�Ͽ>�O�@Ԧ�]��3�	��,P4�SM��s�DLY�@Zb�e�7��-_���T�R��<��՚ж�s*U�-�ݚ��ٺU#1f8���*�N�>=�����{4�f��ܾnmK���>W��!�;f���؎�3UOh5�}$U!�ϞG�'�~��|�;��7�w�ΐ����z� ����r�X���̷����/.���[��N��{;�Jǻ��|�wT���q��)�2C�}����}��ﻺw?�=�{ݳ]�Ԟ/d2�$�kg�3�-�?c�������MS['6���s۪41����nm-K�l\�`Z9��O�<�:z��`�`.�y�Z��l��]b9�̲��`yvo��Xϳ>U�H}$G���}2��m�FK��5�x�-ۓU*<����;����n�G�!�9��O%;���zk���E����b:���w�L�x���6V�ʅx�B�>"r��H3����
�&qi��`.EU%s3�/�}�O�Ο;�����&�ωx��k���p�1-y�^�2@�o6��e��j���G3@ܣV"(Tc��U.׳O�C�"���Ib ���i�L$�H��:�����k1��}^�tX��:]�B��J�j�B���1M��̥��0�lah3b�5�W5��َ�.��߭�����RE�Uϧ}��T�S�w�U��%t�[�,U��:�mwo>�p���,�2
�ST�X�l��5*����ʒ9���޻��#Y�2b�Y~���&�A��v���ˎ�v����ӧ^�o�ҪX�Uq))�0��mJ�%]詛N%���aʱ��J�c�꾻�ݾש	c���m�p����v�V:"�+%�VU���ɦ]�k'w#����[z�Q=�л����ͽՃ�7�U	Ʀ�P�eWL��A�F�Nޭ#��L������z��5��k���*Y
f�������k'��gV&�y����W{�[]1\⼢tKy���s��/�=�o+��$�a�SI;�evPݻ9*2Wn����V����2�ċ������v�n_v^I�&e>�7����j���n�R�:n��Z9if��ۣ}���LT��R��V#\�G���iT���Y�+F��k�OC��VS�=�ڱ�����_Zۭ{��ģ�����W@�����l�L���4v�w���oqvN���:R�}Yݨ���:GD�s=�����t�e����u �u7+u�r巉�ض������M�Z��c˵�f��A���ʅKj���v,�T�qKB�W���P��V�|F��	Hn�#,��)�ywǮ����7B3�ֈ�n�֩�ۢ��x/�.E�a�z����io2	V�t�0�.��{V�9E�$�LWm�*���8e;ѩ�3[��wB�4{7r�7hse�E��~�8�)����Ω�#^l�sA�,
u�:���Nг�@�V���f�6�Ko9��D���W�tn����;{��ۚ��YE�*V)J�ou�1��C��"��v�l�@�����i�F�QU�d��dSINgɷ�0 �V�Z7��b��kr�k�mi*(�����[s���9�����Th�|�6�^V�m�Ù�+�^���_-���y���k޺��ݶ�E�lsr1�;ΣN�\�"�>��{��r۽�(ѾUҹ_�w�:Ѣ�k������k��;\������ߋ�m����疸g���ݘQ�o{�Ϸ��wEr���\�^nn�<�;��w�W���ݷM�]6��w��FVI��9汴l�t\;���$��r����m	im��ɮ��oD$H��Y�k��!<�K���J��``ⴳe��p�\�^n����ח?��ۧӇ����oW��ޱ��}����C�||8�r+S�&I������j�ef4�D&E���'�\�of�3ܕ8��:�biǭ�j=�t:v���I�o9�ׂg���)(Ro�Nӣ� 
�"'X[;˧&�.�����A���Q)8��ȼ��"c@o�_>���@p<�II*��l.c4��d
�f�a�4� ;��{=�o�~�����K�3�|�I���X�=]�k-��:<c����U �\ѝ�0w@�u0p@'�u�(�8>ʴk�����9t����,B����ܦ��x����������89�I�˝puܓ��n��'���x8 ��G�*|�BM�WSŅf�ƨ���E�ޭ���T��s�<t�����(�K�#���&p|8>r�Z�;�`��d9I��RN�{c�t�e������p`N[�<|}m��k�G��s-ݖ�0�G.�aO]s7�R�����W��S��?e��w�>*��:��f��b�c��)�eܗ�ykqQvیV�R�|���z�ǋ����$�\�|`�y��T+r��Ix`��g��}cW-R���m ��r	�o]��]��y]7��<��I�3���祫e��
Ȼ%����.�r@#��-5c���k�L��G����8��Y�����{�6P��ذpgN��d�2��;�#ª��r���hV��oz�_��)3��I����j�ӑ�n#�]��ճ�	�ǻ��~��YMwkG�88 �V�&c��N`8�����*�x��AI��� $��C�}�$��]����l��qb~�oq����AI���8>I?��?��C�>K
�`��32 �j$�����;���x�.����L��:.�Y<�,������j�R��D9I�����[f��|,�S�!����{-e5]�9���oe8����Qr�!'��}��3 ����μ��B�Q���P��&�Q6!!*.bFG�)���ݮ�]����PG-&�G��ִ��#v،�fp�&f��� }����q_V�0��B5�Zg�B�u�F�[�Mv�r2�9�S(vv��p%4	0�0ƓL��[�f��p��9��(�N8N��v��8۵gۖ#In{a$�����v�nm0�8-�ChKL�L/i�	�e�%�s+]MB��4�lc���c�����f���4��='�f���[��:�`���������F��}��D�l5��\s�uX�E�RT8xY.9�f�Fգ��֡F|�B>���_����pT#�2!���]Ǯ1�*o2۳��Ir;�0��y���md9�RO�U �������9����d����`�����ɬd�x�tx�8���V��k�{%����'w�E�&p�N5�Q����"l�j�̣WY��s{)�����(��)8~�̟G���Z�����<"������=	�����z�&"�,��e�x�M�	��S�K���Fi�~`˹������-��%
(���.h��B�q�ݬ��x�*��t����p�����:=P���J.�l�@P�b�.�۫��83��h�0<�1\G�ح�Z77���ʩ����C�M�)'��rf��ِeNhc��	L����ҩ���D�k T�����áA��![��
4 �/��I~�f��g�-��/�2Sm',���5ٗǶ�Y�ܒX��b����eT�(��Z?��r��N�{���5���x��:�gg:��E�;�P��|p�+�[��+|k�%�),�M�7O�����u�k���~g�@�:C����P ���R	�d�ȱ�g��G�d�e�I_�	ӆ}�'�*P#��C���7���|�r'kSv>��}M�;��1�Bf],�ur�2�hc�p3�
z��lk�7=��6P �!%�"��a ���b�������y��C<����K,��l��Kp�� �x�2#�4�`������=��¦��] �.!�%��٭<��g[5뇰v���K�"�DC�3�(�y�=L渢�.A	8}�sul�e�I_������CϚ<��
��R�ܟ��i���Q)'W�5���a���`�qT�sV���n�8���J����`NS ��� {M��c�,�	Õ㷯�&N:N�jx�DG����e���e���2�Ӥ������mG��+�R=�\��)9��ƃp*�w4�F����0��[/�ĝm̫�r��b�/#�g�� ����S#27���D�Z�Z�� �fi����)3�	I<N��D�n�,� �!�#���V\����BL��`�9�sٗ�Z����@ ��<p�5t7\gQ������x��?�1���'�A6�9��h�-�)��x�|�n�il�	��fU+|��?��8U��	3��p������@������/a�A.����q�d6���Tj���h0g�kg�2sh���H���a$$�Cx�&�	���r����Sq�k�I�5:x���r�T�����֯��<g}��uL�%r�4��)ɋ=wd�����[|A�p�:lcf�Ib©.�[ހA��6�I?�2�tg��$����o4sA���R`��A$�oi��[�C^ښ�+>!��0¹\<���-��<A���3�1���j L�R��1.x�<AI��Z5�������S{�f���?����G�4kj��O��-�f{��[+2�d�b�V���XIGCQPum,���}�����!���Jܼ�If��>��{���*� w���x�;�
L�$�A�I�}���<�@G8y��-�w��ņ��x�t�g �pO�Ĥ�
{0��z���m�{e����Ԯ�6�[`�nJt�0�.i�jĲ�hF������>K�������8)7���{�֜����
�p�o��!���`�X��Hm`��9	(�HI����S���A	'��:�d��32���r�Sq�S�>�&
L�s�O�[ݵ��x>�`�S ����&r�
�Y����)ּvZ���Y�;�!�X��pA�8!Zy&Rg>]��vy�# �0W�9�BOz�:�f���/uK��y��9m�\��C�Ui�{�p^#9�����	(�O�L�pO�8�����n<�S|�)��fe��r��A��  ����I�AI;x�^�Tc�ar�Q�D~��U� ��������s��7�L�nU5�4��+31�3���S��{c�!�lM	A�3b풧�������FS`Op8{����>�LU�+�3��]9�; oK��z��x�^��:uۭ_�K۱��`N�<[�4˽���т��s�#�^2�	�c@^7s���W��m�j��lT�=ի�u�W,<2ݢ�gP ]۵�wL�p�����[��㫍y��#5����J�nY��.�3N���:B买�9�u��^�Y�e��N[�nK{$4��n»����
<�������:^�⣟;m�c�����I��G!w�w�~�z�8+ǵ�G�I��'3fֶ��Zċ�gx�w��]d�ٿ%��"值��R`��A$�A���a�Dk��Z�疲�XZ��q��cs�V"�6�ͭ�Lz�G�����s<�o�X�p�";�d���9��#3� I�˫V�M�S��e��S��X�LU���M�]ۈ�l!��g �㙏!�&�^3H�����#X@ �(E ��?�t�ú��ԱYz����,x�ȑ�%�dc^�ٵ����x��|ٍ������3Y��k��xllvn�Ob-5k���[��� ���BO����Ⱥ!�����v���KD��u�V�te�-�1�[D6�B��������p�r{K���G�y:�0���s�����|���Xh.��ɪ�P�g�)��6���I��!�)8r/���
g�<����r���B�nK��9�NTԐ�,��W�{5����F��,Յޔ��eǁY�������s�ޭfC�u�|�u�Z���2O`�/�P������h�#y��mfn����^[=�w�gz���N3�fc��cUP ֺ��q^�:��A������A�3�3F��1_GZ1t�"�"�	pc�ür��q\�AE���	*���+YDc&O�&�h�L�u؛����j�*�e���x��gM�����e�gX�8#���������I8�Q<�R��z,jq2�w��tN������p�x�pF�I@�ӣ�r��{f�I��r �I�J��E�<ɛ�ƅ�8:�� ���7h��2gGn�����yU?�&���y�I��b�4gk���^a.w��vmńᙹ�s)��*�:QpBL�$�ȣG�&��%;E���#�`G�6�.��Nn��j��������S� O�&D8Kѫ:'�LU��'�~aǠ7��8 �́ ����'�@`sҍk�h��΋�TQ��ꧬ�u����+������ݩj^}����B�J��!�tq[�����-3P�����U��g���� 야�0~���{���� ��Lc����Q�8>��\n�v�4�O�<}����)��{��w[_�L�	pc����\���+Z	:l�^����Qr�p�����)u���!F
���=n�U��U��x����&pA$���C��ϛ�|���I�Be�ݗ\��uk�ε=��s���
��Fk��O���~�[R���_ty4AI��v^��3]s�9�+|@�ͮ���S�yn w�і��=�"��� ���+�ﻫ���LX��0����/3s[[��<�\�y�)���(
(�vR�Q�B���J :|�8rQ)� ,�X��3e�FʎYG\�T^#����34��L�pRg#�'�B)�»`S�����ކ>�\[�@�vv^���j���+�����r'�ѓ��9�0�.�7j;���4�ܰPE�U|�pq�\�_ƺ�M��Nq������5�r���ÔA��}K(����\[+b+"i����d���{������w��ᇪ�,��6MkW�@�dC���,���[�� X��Θ�ѽ6-���y���=r��2(ǈ)?�N��!-����{�����4A�"T7��j8qD����n��"f�����o����_��PA���%<S"V�p�ttU���x�d�hǊn�Y������AI?�DP)0s���[�&m��7
{税Q��ώ���,�uUW[c]�w�g@�.G&I?��������g��D9��A�72>I���g��َ^{��*Х��7fż2�k~Y�T�޼�j��Yn4j�C���|E*� }��<I���zA�`�/-�YÜ���Xܭ��&� >�#ns���C �`���|�y�&RP �\l����w͊�M����-�uLUqQw��l��;�rp�#Z��F�x��˧��v�ӧN���mXŴ��"�6o��b`j�*�y��Sq�n�2�.Xz��Y6���[@�*��X��4�(��Wx�)b����aP�v�"�*�}�&��P�E��v�S��h������,:hv��(*nI) G`����d�>˃���eC��A�v}�"fiT��>���n�6�����tPF^̌@�!���n�u"Yv.�u�ymW �%V~�t�_}Do��V��^6^�����O0���7�NS\�t:�ɭ��r�Q��u�i���a�y���Z/Kv�e�������Tdؽ�s�+u���O�;o�\BݓI]n������@*&�e*%��j�u�d��&u��тc����S�s��G��X�݅Pj_�El��y��|K�]n�P�ٖs��;;��^�ʃ]���G�'y�Y�]2۶)P�ˢ�o^t�=!�z�UvIϏkv�����m�DIpV�H�ݎ�0+:��e�*��W�l�Z��e�����2�J�"�35fShu�R�K�`���ݙ��E`��ZP9�!oqy������p���u�}��L
닡����B�]�*.�\�N��z\1e{N��gj��쾗[b���S�[������S����Z�(����zWu�
d�f�_rX���g����/���f��Ew^��J/M���v��H�Wx�^�yC���Ι�n��\��si�ݔV�;�K���8���Md�oE��r)κ�w�����̫]�s�r���F<���Z=�2�خ@DP�p�+TN��6wL�n����ꚘY��4��%we�Z����XEY  (+-,-b'�(r{��3n�0�K-)e���U5��RwWw+��:A�;v�X��lB�V���c),!�$��{�}�^�4�-���4_g���7�tpﻑ�����\߉�Ɔyi()8�DG[�m����_sn>us�'���v��\��@wA"��#[or���Il��� 펶6pWi���e��u��k��#�xI吥��,P���lyy����@�ptG'Ds۝��S�[m�
^��R�:��^���+D�^l�;��vF�+]A�ܲ����Dk���m��y�\ؓk�;y�۝(���-�/7�\,���-�&�u��|������vNW��ㄑ_��0�s�Ȉ����r�u����A.n�Ƹp���~>_V_�f�]-�.��mՙF'u�;t�j��+���ݘ��3��(=��/d;�s�nY� �7��F.K"�J�6$�55���K�ѴSpK�%M`Bl@ 'Y��[v�lj���Tc��Co[]h2�\MX�����뵪��Z�\�WCƜ�:�:6���r�3qպ�VN/k q�n�qn�Ѷ�*�q��'i�&ea	L��m���>y�:���4�X�ka �4�39��D�x[��c�H��ts�n�`�)ëY��A�=q`m��)��s�SF�Ɋ[�fnL�\k[gOv���t�8U��&*��9���Omz#K)
�ֻf�����2XkQ\��WH��6g����6��%�ۯU�#����^�d2jzxLq�.�u�����U�ZK�h07e�Bb�),�[��������l��Ҙ]ID.t�1X���qC����mu�h���8��������'k�v	�a2��Wnj�2�fh^si8�y�䈣n�����Xv��r=�\��ۢ뮘�҇m���C��=3nxf�1���%-g9^�9��i�,2�LRM��X���}���m���\�q��'S�6q��$�olz7v���Bs͏l��r �t-�h���:�$+�^�� Q�-����&#�v:���u�nO#Ѳqۧ���F骷T�n�	S�J0a�����u�;md2�k��ǡ�wƸv�P��I��O9���A�6�-���˞lґ�ƱfQ%tF�3d����G���;K�m8H+��&olku꣦��0��c�3w3i
�s��bF#+�d+�vkv�ƫ��2Y{$��x�U�X�Z��Ɲk<�P y��5�7d��M.᎝�-u�|vv�n���\u�ke�,v�>ԯf&k0:��
XJn4�Z�T&�m�QHRa٤i.��Ц�c�	�Gi�V���X+��6���@�6�v�aK�8wlݵ��7��e�I��<�<��7'��r" Ȁ��'3&YG4=T�֪����!m[a	��:NgN:L���ݴg.]۞���-h���4�lY�,	�J��6&���hV��e���e� �iӵ8p�[7;%uXݙz���#�v��%]���WG7���
w]s���T��^Cb��T�7!&�KipL=�͚1�ífAP��;`�z��}�>7Z�n�ͱu�R�#\���G����6��[6����rY�I��M�8�m�3�n�Ƃ������^�o��~�#�߱ ��xh��v�b�/�����jf�m�����oc��Q$�$�C���	3���̓��![p#��5���nVh�*&+7$��OM�œ����6�?v����Bi�B�J< g�j�˶�|٧�y+-{�&��M^Wy�:#�����}P#�L��Bj�׸RZ�p��p-7�9��
I��Gc!�F�q�1��m���2�Đ���$�o�%3�A��$�@ �9$��K1���mȮm�	���ZMM��r�b�1�&�A&�)��M$�z3N�p�[P�SS������}��=A�3�ٴl)h����f<���!۱��u���E+�M�~��}�a}��H�v�G��c�3>f���OD�Xɻ��6gzm¸�2-˗r`5mG�L��i5�޶M ����۰�=h4��)Kv�A�Y�Er�sO7.�.f��)�WЬ�	��R�`�Z�ͻ�C;2�s���	��:p��'�ʂ�$���9�@��
H�$"
��5Y�峂�ݯ�G�!�ӱ_c|����W(BMx{Y��(�U����x�]p#��Fc�!$��Ra-W�c�>�LU
8��9���7��bi��R`��A)'*��6�m�&���w�f�蚀3��8{���������ɻ��6c�v3�/�Rc������	���Ey�%�)3En�Go,�n�ä����֊�lg/����-��+��(���p��K<Qb����˨t���ZW�4�Wr���l�N� �˦��hb���$����.#9����� > &DnRLjo8s�����ԛ�"��u���k�
��u����j ���� ��ꝉ؍����
(�s�����Kt�k�]�o�3��O>q��I&]��W�)�`fr�N�Dy&�A)'��y��8v�e4u�`J��v����6T�V�=�K-L��6+5!1��e�2Nd���; ��^q����r�4�m=aM#�{�|}�{h�U&��������!��֪�����c��r�P QRq���q�R���"��=4�;���|����Umo	oQ��y�֛�kŁ���+���['Ÿ��V >����PG�C�
�RGO�K�UX�a!��*m^��^:i�*�'��2�O�0�BI�	��u���W]�bSߞ��]���mֆ�4�14ԁ�"=LfQ��n�l�h����a�A1�� ��O�	��&�I�H�@�YO\���c�m�����m(
:\��W�I�P(��L�Î�R���gP�t+/]?<)t�n̪��5��y�֛�A1T�!2!�M����`4�s�I�	���AI@�QE� ����{F��Q�]bL>K�e+��5�@'���?�I8^2��d��V߲���P���G��+]�%$�$y�u�jk�؜�w�`|r����k����җ1�gby�)���D�)1��C�����e�^M��=>�~��SZ!�0)��E��-�|��-�j�\�ץ�U $A�Q��mlU�U�U��{���@�<\V�	*�@(��	8rQ�d�o������i�kv��V[��~��&*�E��A$��5p�?W�GunP s�H2$��E�z�*��&�6�on�Wt�QXƒ0j=�f�������㎽�
(�����[��,�+������׏]f.eq�R�ӮX� �E���)�
M�$��29�gV7N�d��87��w5�Za�_6��͊���H���A�_@�Q6::��w��;\:�	�����	0pB��&D;�SE1�h��uZ�M���GZn� ��x&D9I���RO �S�\�X�85�����v �:\�p��ZVi�i��U��lN8���H�݈���� �#o_�a��)3�|RO ���)4#q�n���p��'����gK���vB��1�	�`+��(��$��}�j_v��n�1;٧a�`��v����W/�!���}k��h�:`l�u�3w��q���ۮ9����V.B���M7�j���5Q��+ERH(��"$�|s}��BUQ�.��I�ⷉ�#�u��5FZA��vL��qF�VM�(H�wk��S�4�;Z�͸�����0<Ů�YC�z� B]vs�n�:��qD��bR��ĔɓF�<n.��j�u�<g�P��՞2���vn�e�ϝe9���@8d5M*�C���%͌U.���	B���{7�z䭌C�e��V忞L�,����}�$.���힗$M�6�W ��\'O6���[kg�H������_'����v0�C̀#�p�5��{���������
���1��o�
㢕�r)'�N�����nX�f!�2h����whn��3��jr{̓��?�'���%�`cX�vi��u�M�x� �Ro$�A)'1�u|ӳ��}7�Rwv�3�Y}���A�x���$���O��9�9�74�����Q���I���»��;*_|�=i���f���z\�Vˌ+*XI�g �ik�>I��0x�8|́e��5*u-����H�p�z�p�:��ݖ�'�n�@$v3����	(� ����a.zUe[Yd��o��z��͛�����M��c��V07 �wC�6�����_��e��Ϯ�/_���8 ����w6���΂��60�G�D;wGN�, Ff��/Y�'���0	�����w:(\��{x��%v,�E�,3����b�u������=F����U� M\���z��\�<�/6h�R_R��ι��'�簏�_�m��FŴU�mm�"�!$���fY�!�w��'�ê�����ٌ|I�*v�q��� ��4�7K���=;l������?d^T<s?�V�G�I��8Ys��,��1�ѯ��P�-�evZ|��$�jnN��G�&Rg"�Z���3�/u�oX4}�����v����Jˠ��1�om�T��k�2�ǘ��<\k�!%(���0`p����߷&W3��w��;9�pޞ�n�lģ2��7A���L�r�8 ���.1�:<qQoPb�Mf�)Xe���Ѻ���x w����7T]�Ö�!)0#|Ƙ9/i�>!k��>n��&D�e���2]!4��,��E��`*��x�G�4�)'�F*�&۝�����"�g �X�礚�m��SA�,�p��;l��EY�9��7%Â�@'� �'Z��	���F8PD�&��[gl7	�*�=Z��ԻY8N�$�M��ё��w��km�ӻM��7d3�:�ˆ4��s֜�J0�� =���5b�QTE�cEX����������!�1FeN�o�A3t�!2!�)3�A)'�p�92�p�Z�4���:\|���T79�ѵՖ��O�:t�#d[Y.�����m�F��=~�b�� ���� �k�.�v��<g�Cǟ.����\Ћ/���pE�q ����$�`̵8�Ǐ���KSb��Y1a�\�&���u��N�fx.4�X� �(�nx�����T���![���&D8U�F��Ŋ1T���Bo�d��A��;�9�I���W��?�{��w����� ����q�V69�s�=�ӛ����K��G'�,�՝[j��o��� ݳ��^<Ao'G�5)'�|63y�5_o=N��9m;�4"����;��"�@�QE�I����5<����`��c�˟ȢU�!�;z��#OZn �fm�>2w���b�B�N�����N��������ӹ4H�!��m����WZ
�x�;�,Q��w|3U�6��3u�S&fCD�S>��������V(�ب�F��f��w]C�7�d$�}�-���,��� ���?�v�j0�AV���s#��i�b{-�;�˄xt�pA��$��""�g�a��5bY�s��;�D/jLt7a��q�=S��s����e��\�:�� ���;O �a
M��I<S	B����c2�67x��׽)�[�Z�&L3�w[���`�����@ �j�vIC�?�o:��5�w�ʾ���ûyݲ��*���A3)�}�ψpRj��5r[I�g��_֚�Ey�e��%<R`�����s�h���A�Y߶�3�j��;���Ð���*�W���T*ӛ�S
q��Z�*'���r	I<5B���=UBlf_����9�ovnM܌����^=��f�rQI��Rp���T?F��gi��W7�^�n1Y�e��*�����f��F6��3���w����͎�Ȭ��%ܰ8�(�}���u��[Zr�኷s}f�mX���̚�d����f;��~zuOuq�{�YgqZ�,��3���w�m�5�Z5Qlm�"HH��H���"�}�γ��(ݡ�v�O<nڒF�=	���ڢx0�mwa�t�>F�q�$��{�Z��c��7�۶9nW��n:B.��s�(�/V�����p�Ğm+�N�q�ӏd�HS@hV�Zh���`��1f��2eaD�aݴv�\Eڍn7M�5��Iq[�!ƣ�7`��{&r��=�k��E4ٳ�\�i+e�.��ƛr~P�>}�=���,\Mq��� +a;q�қ���ݕ�W�X�3D;g����0&S ����QE�)8p���Z_L��T�Fw��� =��o�3��nr�|A�Ñ��E��"�>)'�: ���.�d��I���z���R��n�OUP�×���i��֟ȣT���C2N�c��/^�N\��8!Z�G�L��2�;��%Fì
%�gjӬ^3*1L��w� ������&�AI<�p�3�aR�IKa��j��t�r	8m�tP��1ѵ91�8ۨ�|t�zwQK/�#�_��l!�Rg��<z���#�L���`�-�yw;\w6F�t��	�9z�y�9L��@��.AI�n�y�����բÿ�C;	�IcكjܸB�i�]����m4g�zG�n9u���?:��p�"�BK'��1��>�ޚ�ts�ʌȞ�n(���M��*���1���� ����L$���i��	ޓ�د�ukn��U�!~��[��0�fu�,x����V`ӔY5��ۭ�@yԫL�--��+��B��9O�걪Y+0L��1J��� 	�'F��S,h֍�����F�I�U%�/��� |h�r|��o�5�a�y��|�U?@'�?'�X�G��V������A�ׂD9I��b�:ll+���	�5�T%=Bo_9�l�b���í@�Qs�BN���(#\q�zl�<�(�D�5�`s�<S"����wCp�YP�'���ǁ�)�9��E��pA�<�8&AI@�ky׬�͛y��8w���%�g�^zr�;��ހH�g �����J6|�1�鹼�Ws�� �@�2	Hx0�*tK%&����nm6��]���"hِ��71�]߯���ϬN�y&�A$��J���
���͝���lYQKa��A.i��$��IDI����S���9-'x�Ji������n��0�b�'���2� �o$���кx �xݶY'����5�8��VBkVr�{ycn��=�>:qۧN�:t����㪧9��̙�WB����.��2��щY�vl�kU�CC!���!��we�F%�/�j.Q=���qOK�V�՝Xd�:��(��6��)o{3z����՘�.ys#���u�t��V��>�v�0�x�ǖ�,J�%����.��	b/g^	u*��}a�q��m�n6�MVi�]���v�yL`QZ[�r��[O]	��D�[��)k#.��t$ap;QkY�;�|%n,:9\���ͬլ /on���wJ`��7��fr7�Aֆ�����w��C��n�q��굽7r�U�i���˼/;�	�C����6�cH�"�pXm`W�s�a����B��q���^λv�~n��{�ά�`���q9�F��D��`1	��wC%�+d�����bͤ��@T8aZ�w���d������DoG��͖�M���*R�B##
@�lL�f=4���5���y�����`܎ z n�nWH��5}���{{0�Y�%f�_�ՙV4�Ԁ�����[�ǰ��uԼ�oi�k��"�U��[O خH�N�-��5��U�e���Ov�/�z�;W����<��vIkl'B���醸�¤�.��B�W�A�)E*7aV>\��`���ڼI����ڀ�2;]�
���Z+1����%Ń������5⏨��{B͹��ek�U��h:"���@I]</6�JA�Vhs���pM�w,��\�Yk"��ľ�k{��)
�֏�У-��GP���;�̪^���|������;��s2Dn\��r�r�\ט��ҹ�|�o���2Ļ�ܢwD������$Q=�vQ����˗�t���F.�FG]wuӜ̈���!�˜܎�r�RNrWu�m�"^�gs�B�Ŷ��3�i��^���;�\0ד���y]�1=׏nK��`������w_�2Ƚ�#r�)��t���nn��p�ss����� C�[֡՗�ix���owQ�1�p`S%�+�v���y�w�C�%	.�����л�L\�ܹ�s�"iӒ��DB�B.�)!s�B&�d�����q��v�ߵ�%m)�6�61[������|=ރY}$��ODC�[gz���H�g ����	(���I����-���w8�A�`��3�$�*)Xܮ�����/���RÁ��k6m�)�E&pA����9	0pBK���UQ���b7�sY�4VV��&-�v���aDP)3�䓷֧�Άʆ2��E����]�y�Y]��n�Nk\q۱e�n4c�ꤹ3�w��<��1�4���QE�A'�z��w���v�M��p�M��|�ǼA�p�+��QRgROj���L��׺|��A9|���l��6��U����w�S�AÎ|�a��,s46XG��؀Aӥ�!'�Q>L�x�]*���DE�d���C�,������	���2!�)3�	I<�p�Z�
�$�I��E$���|�xwg�'�6w���
<_�W����8�-1�אhի�??�5]���sM������0DAǡ��ˋ��	�U��(�\=]s���Mp&Xj�w��'���W�
$dA�A;������z��&s���ɑo)7��*����v~����I��1�`A�`�}�@�QE�!'�R\i�O%�!�\7�&]�cs���4��-�hֲ��;v
�^ݙ�ӹz��ûg$^��:h�5�I?�2!��s\7E�S���p>
�M��X���k!��9�I�N
LW�<�3X�b^�`/8}�]������gz��<8x��jp�$���Kħy��&s�h��5�B�z[^2!�L�RO�;��Sv�V�3��t�6E+�/C����rP QrIÐ����݅LkH�m:�ģ��[S�Z�<E���&����:������e����F�wD&�Y�o9�O$� ��8I@���������>�t��GWo�b��qFw������A��$�G�O�����t)��sc<v�(�.�H��yi�C���4�@�ޢwâ��p�^�O�)r�k=q��*P�����%�Apꝝ��]�����יC)��xi�Yθ��|prz=AdA�T��V��?<���L�khW$#��:͖�GKh� ��Fĥ�і�s�i��]�����j��Kz7���9�n��1�u{h��$�ؒ#���ut��s�+�
ZY���p1�/liT�.q���w�Т���b}	e�է�-�ϥ{'D�y�띓��n�!:���ml���2�`n�i��Uf6۞�����Ŏθ��sE�μ4�ٜV�C��f�\Ϟ�����.�W��u�yy�[��m��v��1�I�v�v`),�d����(]�c�Ǝ��~�x�o1�VU�wWG7E+�/�;p"��M,�T�c�v�
q��)8�q���x��M�ף�� G��D?�nz���ac�xμn ��[� �q7�z&"������>�D�b���i����3�fd#1���3'ҥ�q�%[�h-,�{-��zi�q�� �p�$�<AI��P	.�H!�d�64wY�|� �;���$��y�9��ʒ�/�#��`:���y�\��O��>w8y���(��8rT��6��'IH�r�|Bn!�w*�b��	X��3���x �=��pRo8)'�L��ۂ]�c}�,z�9pᡡ�>�q��[H�23�/��ŻBƸè��
^@�g��x0&S ��(��$�_o�<�ld�̭��t�P��64;�[>�m8r+u�:)o <]P�;�{�O��A�K��>T���>p��e�.\������y�$3}��s�KM��]�~`�ӠT���u4�ᒌ ��ĝ^�ந�U/�:���H0���GƓ8>����*�����!J��1�`N� �Ãf̽%S-��������]�����T�L��ed5[�SG�����?^ҹA�J�I�6�p �=U���t�V]�2�a�-(������&E�c�_��`�HL#����܈�)+�K���y�aWwPt�6ӴX����R��P��C!!�[�C���-=�������n��)^_9��A�U �V��?�z��Ǫ&I-P*�d1y���î��R�v�Vi�]40C�^ViT�߳}%������Ȼp�[Y#���*�?X��s�7�<X>4D�oN�!��g���W�AQ�BCK§L'��2�>����n�����i��̾��8 ��}��.፻s�r7����),P���BCHK(P��]c��.�B���Ӷ���jf^f.����V׷�r��H�6�����+k�v���Vf��p�2�@Wr��5�L�S\�eZR�2d��J�� "�ߚ��}ou�fh�gy�]�#7�By�Y�l̰����Zq��E�pgś\9���#v��*�tX��9֛�&i��n�l���o3WT3
�@M5R_�
�T�b�j+�ᡡ�������b��̾�����O�n���
)S����~�����]aΦ���i5��H`����\�舫s�M�Z�]��w��Ù}�#}z(7l�b��2����J�����㐕�j,�͕��ARp�W3�n�9nE�8"��'�k>�w���-��ʮ����6�q�r�ci�����חYGì�w]R�3M!BEJ�/��LAS�1J��n�jk�V+����7�n���ya�O.VB�eY��J�������dC���p��4T^?l��M�	^._�v�9��#SV�ƨ'n$ć�=pR�=;#*-�d>C�v5�#~��;2q�j��(��j�=UtM��m��s5iu�)�'(dRԝ�ʋ���=/�$�H �vza���o�,���E�y�v�Ȼpy
�=7ڛ���V���U�up�-9o�Y֛��4�A5m�СBC�
�\�bN�P��������E�SX��lf���q�ڎ�\����Ga������?��X
��Ϯ�@�stv�X���3�/�+�p���A�d��7lݳ�=v�ב��*�bۙ���I��U��Z}��H+X�͜��`~��LT�&���U�]�L��
�P� Eۇ�笞O�y�����|zδ��P�@�T(C�7C�*�ԟ�<ve�V�0��h�r�p�v��glOY̬�K�\x�Uǚ��)���<)U	
��
*=!��;ە�T�W�k?�2�3��,\w�W�E�#�[�'0�e��c��w�π�����\yc8�}d������epV/F7������ͭ]+g���Ev��<,m�3o��gx��@ve�,��m�[����,����eCj�<��/�w���Խ�ۣ�wJ�;.�ؽ��s)�nHj�v;�mv�jۙK��&�B�X�4�huc�IuVe�9e$%��\,��`�\0 �����hy.ת�uZ�y�B�y��&�d��cN1�k��h-�>n9�#�ݷ1̈́X��C��6�d���q�ׇDtv�ݱ�t�j���ݿ_�?�r���{\�A�VK�v�C�d�c�ԭ�1L0n��&m}����̲2\��Ñv��md8�뷵���NRȊδ��'��	�=�b��q���d85��n��"͸`M�o�^8���L�1-��h0x��dm�kta�=g2s�/��<QpAm��	F�e�t]Q�[�p�u�YM�6ed,��dI3+3�7�L�F�^ʩ{�@��Յ+8Gx�0z��l�l��&����=l�#������R�R�ކM�����;�eu��|jY�]��;p�E˿;#<�}���a���9����͛�4�owu�*�v:x8�p��1e��P�ɳ#;��^<.An��mdy��/�������/�1�鵕[f���	fjF���e��I��k]�-ҳMCm[��Ǫu�};Og��9��-l�8�����9�`z`�&Ò�w8&6i��)��L�n�8�06�	�u�Ex�w�G8��&\w�����$���,�bw�,�v���}r�
�ii8�u�OC�|%_u�Sv��Z��`&�e��* `^�q��8�����&���}�����q��z��M�jY�5��ݳ�f�_W=����
�j�4���*A�"�����$�ڶf��jVs1�}/��(�l;��=md9�o��]�)2?���u��ճ��ϙ��c��d,\��0pC��/7	��Vz��|�8w�� T(H�P�/W������Y���j���s�M�Օ���Գ��붟B����C��|�~r�vJ�����Κ͝XpL��h�ZԆ�MNϞƃ�7c�%k-�9ٽ�^4i�zu��c�6l���p���5��f��M��~%��)�P��snzk&gp�^#��W��E��|n�|}v�w�ڼ�î�\m�m3�:�êZ�:���U�u���sSu�plن�2;��P���8 ����Ñv����^>�|��J!bS��g�m�9}�i姻k�F���*�ڬ#�؀pç��z�l���{�X{c��0 ЦlК�]G*��
�O��B]�*�/]u�!� ��붛���f��m���S1<�]������|A�ۇ#u���*ݮ�gP!C��%��F9~�Fc����ݳ���P���چ������;�|R�{���6:�c��s�r�nٲ�$Ue��W����b���&, *nc�Nz�W�B��/�SڎE(y��/���ڿ?�j2x��c�"퇞��}�X�28Uv,|3���Q�y�>��z��C*��UHP�"4<$4�rʱo�>D�};A��hYG����,5�qWw؛;�����w;x^�����s"ܷ��7��n�Ϯ��1v�&Ʃ���˨eV1�_;�����u�6\�v���ԍW/���J�����B�4�@Լ#Y�ՙ��k�c��]i��o��z m�;B��a�sE+.��sQ��"�0�jaS��������q�2G;t_{Y�E��eA}��'��!d�Y۰��f��{=BD7\�3�+�YL�Y�aD ݰp�`�rP ���U�՟����4kۆ��%�.�Rn�f�?���oJ�H�xz*N��x}x\���#8Ѻlݼ�W�H���`�� G7X3X&��3��@K��i�
�(�����)U_����-�[��b�:�c�_;�a#+A�uH�D6��`3�Ã�˂ہw>pA�e���(�Y{��\�I's���޳dHRk�3#��b�Ê����Ʃ����C���zc���V��rI��t�Ylɐ�2�k���5��ٳ!e)�{�M���8���E�y&DQI�P��wD�6շ���g �ݳmR܎k��c��1����`��o9Lr�~������GN"~5R] *�R*B�Ʌ���?o���Y��l��=���7 Ae����&eYʉ;m鎞\t���ӎ;W������^�-�KCM�b��Y��J�r���r����y�Hm��@�tQ���eu���IαϠ���]�Jv���x������8އ|��Vm��+�sYk$2�J��yq铚�#ji�W����xq��V_1r��Z�d�s,ԝg��,�]C2aoL�A�oj˕3�s�wgk1�я��RG�2���*��@�׏p�c�R�_v��R���[���G4=��e�8�u�`��и�X�z��0wO_���6�M��9I�qy����ۦ�����5�ᕴ�}�w;���˷�Vu2�>f��f	�A��sw9�yY�A�X��w-r�!0�D���J�A�E��D����4���6�o7��9f[�9�SYk���K�Ν������X�r�2��KFE�X4\t�."�q�B�z<�\��E�+�.�ג��{E�ُD��� �2�u���=�.K给b��e��t	����}N����@%�:�v��7�=�e�J�4�����u>��W�Y�J��F�Ym�)�t����,�8IȌx�bZ�*�8�5H�o\�yY֦b^���,u��;Ρ˵���N�mv}v�wŎ���߲��gG�fu�?er����s��Ӝ�'׹ޒ�v��#�N˃EN�����w�.S�ẹG����R�5�n�%�β#m�t�M��+.PJ���Q;D�L�(N��Ք5<�v��r���y��ȝ�15�٨6l�
T�ꔫٕx�,�]�M|���a����u``{(��a�(�LG��Z��J������Y���v�mM%J8�X����W�<}?�͒8s|b�����u��~�R�Ww����fI�t�>]�ӗYspĄ��r��w������s��;�{�{��B����t��1"X�%�!�z�.�2���;���7���!;���:��v\��w.����H6
Owc;����]w\�9قFw\��^W0=�Y�����ur��s��7*�F��ٱ��{���Y�Mss$F4=����%�����%H��b��Й5s�����wWE9FB;�^���<�-25�u�MF���hK.n!	���DQg�2r�/9�̙�B�q<�^딇���)��j�]$S��b^[�I�s�o*�"H�o���~w��y�^�q�'g��׬q�Rka+�^�R���u�=�7@�^��v��rl%�6�y�sշ��v��m��-N�XA��2�7T�˥Д�P�V�!
�������vMy��5�u w�7�籗�i+���6��[��z��ls�Ů���]�[krmk��Ip�ؑ��hP\=����&\b���x}&��+	Hd�i����A��� �5��8������Q�[����vO(��mĹ�"����wk�V�u$�n9l���"�bF<�fq*�܅K6�y6t���7s�"۰٣ 9�k�%	D���K�S`�6FL{���6�3�z�oTp@a����v1μv-G��Y��L����[^���c�D�]�LAv{sZ�Z;q&ܽ�����9;O�P�>y���0�Kqz��T�� ��9�;Xb���xI�������v0�.�m�+<�E�v���K����@��;9�n��%D�����K��琂iP륣���ˏX�l�l�n�هE���Tu���ɻR^�CX8cx%J��:X��#�n��+�nE��:�)'+�ϗ>�u����,�hy��rn�F�q�v�5�l�;]6Ф��]f&5"D�l��̠Ŷ�lՍ"��DT�%.#�b>��8���6*��Ms]]KBY�[+T����thAe刖�`uHvVp�q�՗hz���s�']����k0v�m�� T]�5���c��4ˮ�K�2�2������N����l�7m�;�P`Tۛ�iћx!�G9���j��0���q{P��N�M�s½=Z�r�9.�*��"dt>�xD��:zHRx��1��Rz�ݻd���z��rq�ʥ͖���n�g����B�Ñ��N�̽^���`�Y���6�˃�u ��^�K	5�C��hMku��])R�ohb11k���df�z�82�4@�	sذ��F2�q!>�]�I6�������$�	�I���!|��ZB��M�`��9GmLT�c��wLÓ�Iz�r��l�	v^�v8��\YN�6�#LH@�1�����F�̰����r�7l��K�1*0��$	H]*lA�eK4�HKʻiH�0��f�<�b��C��r��h�P(:L�����n'&���'S�ÇǞ�̩��"+�����\���Y�� Md%eslٚ.�G:S��?����ϳ��=�h순ּ�����T��M���#����A-Û6\�.�7Ucf�.�Wo}xپO��9�muʹ��x߅
�T�g�ʡ���}!����Y��g�H���A�f餷a�-���=b��{�9L�Y�[2�nfѼ3�@�A�.!'�p�"�Ș|ax ssP�ӝX�Y�s=���M���^=�Hn�P��#�_�G]�g\T�X�ܥif�`mÃ�K��v��*�6";b���6w���n8`�Ca��M�b�����|~���
�J��f��(��ڗ��ާn��n�91���0 ���/�ۃ�:��v��Jy}�<����	��MX�ƾ^�'aM΃�� ��;����lk������F[��V�8pEۇ��C��dۇ3Dvf=���M�!�vCV�w݉k�4���g ���j�����ݿŐ^Zҫ	T++���A��f,�ՙn�A�X~O5&�G�w}ch�n���-ؠ���S~��%�rNeMݴv�{��>4x�&�T�������j�
�'f�Q�ۇU�r��rw���G�q�
4�
��7B�	�2�v��g���o��S~I�PY���L�C2��e�J�g��� ���G��ɑ�X��p�Ŏ.��f[�1�	�Ď���:��|�o�
��@Hj���������X9���Î��ݞf�۸������8���9�f�ݿ��\�52!L��~7�Sq�� c\�f��aZSf���;��O��ӓb^�M����tz�(Uo��BB�P�)-~}��P������5_s;KE��εUA����tr��Y�rd�S�&����In�]?��Z�d�O�Vp��N*�p �2�A��svێRa
/���i�w�i�`|o�9��؁xw��U��\?Q���뒬P�I��͕x�mݧ�d�'[ڸe��׽��a�ٜ��n�;��k�هgU��W��v+f���+ԗL�������o'���S��oye�̶�ed-��s��s�5-��O�wB�0U�ќU
�<b�͛ht�Ɍ�w���[un!����8Qk�!'pG��.A�p�"�[�7}����D<U�}��v$��3���P�vP��
BC�T$;a��~������{�+�st���	Mrn�2�!�
�5��V�C\�&���WK�>��;��=e���͛.7nr�W3<��S_e7y78d�����z�n'dɏ@�p�W7��Ϯ�H&���f�(MgOJ�2�Ȁr�� ��F��	�-?3^L�k���8�`�7�8sfJ�cC���"택9,!�E�̶ٕ�ٽ�s}J��.����9R�����	��N?�(U���a��>�g�n<�Fi�sÍ�{<� "���<\�v��V����U�_e7y7y�<Q���oLk�v���XYP��L��L�	�Xtт��,P���AJǄ��ʇ<O1��&�~�읷��O�?���vF�8�_i��G���*�#�?��9ݷ���sv��]��P�a���?�r�x���y3��#<_��w�3n�Ѳ� ݸ�˨1��a�ϡOb����mb�6M-�l�n�3rJ�ЎvҢ$ь�<�h�6��s�>}��|�6�GR�ђucr9m5�����ڷX���D�'׭'�m�6}v�����yx�FfDug�ْ󇞥�3�5֫�~�n�npO.F[ T�r�y� ʵ'���¡���
���DYR��붿U_�k�a������Vŧ�jS8�1�8l�޳fH>�p�]�!��A�jE��@����Z��E���JV�0Of�#��Y]x��e����#S�Twl^5L�H"͐����"�����{}��*�*_�7�����j���-���� ��H�xC?U��f�D�_D���3U�,#�M4+��LPV�}�V��!Gn������Ͼ���p�}��X��!�˸}fі	z[���cl�3�4�����'�Ϟ����M`�d�RSikS�#pv2r�]�z¶C���������.����Is5�Y��!�=���=m�Ws�k����V� �c����\-1���O\ ��m{nB
�S��qW۶��E4���G��"�F��[jk(^�mg�Q����f:ۍ��s \����(���MW�٣n����*���9�z���Q���6h�e;0�Yv����-�%�#Y�ntҨ2�&����VY~����c�צpA�<_na�}�C�T�p'y�W)&�q|}n���,����e��r̙��*�m���_��w���'���Y��e=e��7A�g"͐�ݴA&h�Ǟ��=�#�����r��͟Mۊ��Ӄ��:ީ~�b���n����ㆋ�U�pE0oSQS?�7
q�������>MG�ZH>7l�+�;�)'�K�w��t�Ȯ���ͦF�N�$��Kv�L��,���MKa�E�39�仲����]�����Z��e=eW^7x��j[�-���]���]|��g��e�'�T�ͳ�+:ʳsuؐ��;�I��΂�p�֩�f�?a}~�^�<'���.q~8p� ���KtF������~�oʇÚ�m� Ѣ���/
�K���J�HU
BB�/x�֝��cE@g��1�W{)>�r��r������;��|��ǧ휴���u/�Hy_<����I��KX�x�:�|^fMܥHx�t^Ƥ����O%���T�Қ��1��S �sf���t>�7f�g�x�ө��G2�!�W,8��o�/-���V�s�'_4,��������>P�J��P�BB�T3���s���`�{u��Cy��.�a�K6
qWYwϔ���8��f&�k�}C����HP�$*�
�
^��n᭴a@��3��僦b�X�&��w�U0p#mÃfːn�b�m��!��fhq#^�%+a�#6���c�P�'=�ܑ�(�n�pB����,���YwE�̴�ܙ��[/�cw��yʫ�,o6ɍ��8-q�DQ��3���n��m�v�u��S�N_>�a;T��`멛�I�g���i���(DY�ݒ�6���ܚ�!d�@��Yed,��q̪b֑�KH�ߐ�A��&�wAf�銫7�˞^�wH'�v���f�p۶ ?�n<Z`�`X����kp�O�fJhy�����<Z|�K��|ګ�����6fl@͂�'��~	T��n�<l�v��"�5�ގ&n�5Fȿ����͞#T�VN���ಞrk�� ��,<����g����*o��jj�u�/����.d�f=����9��z8pX�������}t�&Ⱦ��8'L�N�zE��r�_O#�=7�����I���<�,0V��Q��R04q6���0.��n���Y�</�P��!!������鉱z
��w����N-�.�����a>��=ۇ]�Y��sd�g\���D�z��>��읓3��f+}���</�R��{*o˿qv�+�=Í&�/0�����0	7�ٲ�q{S�������^���u�<g{[��L��-����6�}v�D������� �&pF!��g�v���M�1b�w;]d�c��$�����>��Z>t�-x ��䱶}'�v�-��۠�;q��[�坧�,q4�e�Y����g�m >�RnN��t+��9��¯�*�v��>4\{�8"��6\׫��Q���ÜS?x�#z�Nщ��j�g���P�/
!T(	�;�����K��e�Ͻ�Fֱt1z鵂&�ඞqd�kuݩ .i�;,v�w��|�Kd����386l�������J[5��������=[*�^��F��=0Z�EC<��Z%&pC��\���/��4�;L� �L�"���T��k��w�U3�H;n�͝Na���!�p�#u�p�pE��m網&ɘ�NUꭥT�6�,������&i��������A~�s��\�ټ��&*B.�a#in�~�p��c�o���	�%�1�u�j4a��l��"	I��"���9��>/��=g[f�=����u����U0l$6\�qT��j��h����ଓ(�f�D�o����p�2�3Q �ef_s�{�oH�[�� 	X/8r��[���trO��6�D�0O	�Ce����".��A��ř��O�^��t�n�؛��`�����ȴf�
`s��`XLJGhF��l��s/�(e8�vۆ���tw,p n�bα�%�TV����1�m����=����mn�`�] ��ICɠT���M��J9���<�.��/�]n�k�� ���EϞh8n�G6� �S���(��zv��5���ݢ�h��]윅˙�:�~�m������41-5ݗW�;�1v�y�1���N�]4�Q�1����ߤ����l�|�c�z��mf|c̗vm���^c+�[���z�Ar��ئ��Hsv�}v޳r]�pDa=���1���2�4����$*Y�_�\%�X�=�~pN.F[�M��z�3v�<�}�O4x�~��
�`��zC��d��"�eo���f.����w�S���
�A�p�ٲ�P�*!��.��ލ(\T�/[Y%-��U3��d�®�n�8#&v��mG ������f�ݰ$=ۇ"�m����q��*�Bqnk�u�K������8 ����-Ñv����?�ύ��*?�e$AI&L4�.;t�&B�=(�Ӝĭؚ��uq\�$��N�}�<A��`���ݳ�Wf�5��+�v�����"vE�:�l�#S�jg����g3�|||�)�'[�ߝ��ZQV]7���+������ڽ?W[f��B�x��J�VCj ��D��^Z�:l�����2^[G��O|,���0q?-���S��9-75׭�5M�)0��f���-�i ��V��"��G�͘�,:�d۬����+U�ϖY-��}����s,�;�.�l���W/���ˡ���*)a�]P��[U����kB�:��`�����NEF7Blx�pA�p�]��f���v�]���*\��Q2��\�N�#��u]x�&����}v��A�MH���Z�P���+��C�R4��E6Yh@ګY�Lp[lB��E�(g.��;a��������ü�#(9��6d�8��f�tS2��O����1������T�t>P���P3�_���8��x���U��[8}�7��ւ��*��c�pS#m��fδGE\��@�q�aj�.An�̶�ed嘞;x{q���N��:q�o����CfF�2E��VHy���S�"��^�9�n����)NWS����*&�1}5��3�gs���0v\3��ka���Mu�m���٥��e۳����4����"�#����{�Oup��q��kR//[��I�r;���m��ٙf��w5í9���A%n�zN̺�`#.B�9�=t�o����	�s#
b/�wu��d'z���C�L�:R]YBM�z��ތﷶ�*k�A�٘�����$�u��1t��%lخ�ճ ���_b[�:�K�j]�O`K-쓳A�Y��	�9eѠ+�)c�a�9�uMt��(��9I�hp�;s,guwF���]x(������uB���RW�,�X�wS���m�[v���^�+7x���
�/EGS�u�m���,[z6e�$�E�[˕�q�)��d�:��W\�z�k"� (_j�9�.��x���O����v�����{�b��0�]F��������e#3���Nb�.��s'��j�n��s�.�����qJ�NVK@;��h�4;�*�yBi�n�[�Lt뷉;⌾CI�{�%��.�Ե�wuYt��u
�un�i��)��L9u��י�&`:3e�z��1ڝR�2���W����R ���/��y�]�0-�L��0�R��+fޒ��h-c\�j��;]o��2��iȲ�oe{k@������@B��tB��u�N��z���UeX��uk)�P�b��5�7V��H��I��Y[.\��N��yG���-�9XwbX�s(�۶�7���e^<R��~�9�}�ށI�|wb�&c�L�������ؐ���$h�d�\+&��N�w2���#r���r�F؂ɬ�F	�]2E�-�"-wW0�TQ���H;�BL�b��A�d��'u��݉1b��b$2�N��5r���`�+��ag8�]9\ ����F�nnws,F�sr��ۛp��5%%w[�����t��F���4h�pخk�Q�E�4m����E͹s�:�J7"�QbHFm3�\�#F.m͝���� ��Z9�&��	C ���cR%������&�˗$L�bѫ���av㚩��p���bo�A3,� ��HH|�I�N��P^ۺTV��Z�1�}]�,8��o3�@I�	���ڬS�5���k���E�O����_����d^^;M!!��7B��ҡ!��[S��5�ջ���֑��i)�6����(W�R�
$T���7�4���
͘��%6�sc�Lb2ٜ7<k|���eL֞u�s�F;#%����`.�O��4ݮ�&f�7bص;�u-��g$�����w!��I�x���b(��U���v�ꑵ��tdr���~	,�5�� �!�P5Cvu��F��k�5k@ ���A)0sv��	�n�������i��&�]�%��Q�ma�S �nv�A�p��������-
�^�mܒ!8��z�hm����"�n�p>�o7����P�Trfw����ОSӦ�^_c�<�^V �����!� �cc�|����Yge���Ö��ʁf�3����� W�V���_]Ռs:x8r�,̲�����N�Ez�'D߰5C�>���Ω�29Z|���y��Y^3�!R%�BCKPqAj����#���i	���b�q��f0����u�[i$ɧ�E\�-�<��(P�����K�B�z���/����Mr�c�W��ƺ_�a���^,)�q��N��8 ��r+F4���1�z������v�k�n�7uڛ��e���sv��P���{��G�7�X8 ����2>�p�[a||�O�p"���۪���I�;�����K�Fr�*E�^�
�@�߾�a~g�:�C���&�>���隞A��W� ޔ��C��E��0Q�c	�����fˑv�ȻD�]�uM���P�C�j�mw��\0���jn��̳�i���g �nټ}�^�r�h���������Z[ ��[�#}k���Q�u��_�¨��j2"��}W�t t�Y���"�o�g [�GQ�)���j��R%��{��v��T�Y�3���Ge�#9�[�n$7�[�]F�8����{36�f[&�]�^F�K�&������)���VM��j��x�� �f2�mս3�`ܜd�a��l&����D�Jh��m�;���Z�qqq$�^qɂ�	�\�(��.�x�ݝ-���Dt����i����JfYW l�3cfNz8T�\Y�ڞ������������qgj����c�aJ��l[���b����|z�9n8sfϮ�Mm�ΏuX���c���&57t���2K��o�G����Qn��n������L�mL���$�9���������O!/�+�t�q�����l��X��9�h�,���3sr�fPfr[+!�3�kXӬOT٦M]�pa�����Ae����/	
���K����e���n�4�
�p��Ӆ� ����K���X�ҕ���#��x�r*��tOE�Fˇ���]�md[Y���#��ګ���?�z�v��G!/�+�w�/7����7M*��B�BEW�����IY��Ӧ���@:�ٲ�Z�.�p��T؁(�Pņ��f
��&�W]W�%�h`�]��~T�dT�!�NZ�Z���殷m�.��{GU��u�L�rg4D��XC�h��e�M���ᛟ�	j�U���3R��O[6�d�5��{Q�\Vm��!g�yo!$�B73��A\���ԟ��u�����&a�Y]U����/�f�x����jKYw�&�:̙�l�.>�p�]����1U�o=G��g����q�f�pj���R��~r*�U4䠠��uG���c�����n6\��v��A�7{��F����CD��5�~1n�Z<�>L��XwN�^)�e��mk{��9�vҖQ�>�e�A��UА�$T��?1���R����3g���'X�{�<��x�r�p��R�T3s��9��qm�A6�s�s���8�v]�D$lu��}zr`.�Y�ʜ�c&���pA�6�ݷ��eb����(�wJ�|\�7��D���>3��Ds�6`B�4�'���Έ"B��l��^�ڟi����	V�p;��w���L˹�md9�n�$�5m��y���jƉ7�.̷&Na2�c�a:��3����W����`m�k�ݽ n>�r���VQ�&���x��qT���E��s4�J��.K5�W��a�݈w��)\�T�n�G{k����K�[� ������ݳ�(S��u=5�n�AM�9�gn��~�;��G�u;�w|�7��9
�hnࣅ�4I���)8~��8>(����wqZ6�7�.�9��+Bnğ�����a��,���%&�جݪm;�~�F��Y�~�:�(�m���J:{<�[���5;7A���i�4q�S�i�-��E̙-!�5�֍��!;v�1\o��^�[����=�Q�Es�f����sv��	�g!�ս�u���%� ��Ǜý|�j�⫽t�u��2�9�f)5�)��J�^�
��%�|>���
ȩxCfSj����)�p�P��.�Sp���lՉ
�B���AO��:.}���P�����"�Í�����:�2�W�pA�'��^or
;�ۧ�k�e�j(;qlw��Xo��o����Ŋu������ʽ�{�W�v�O�w 31u���j��@�7�}\F!��m7V�*8i��<�C���@��붼];q�I'��N�F�[[|�j�⫽w���`�e�6\n�-���O&��C������'h{�8��F��M�4�	��7,r݄G7"�[\߾Y���Y������Eۿ��'mn�Y�bn�=׭������X[m��r��M�8"ͻ�v�F�I�v��KF����8�H%�ԇE"�2㽵�pN.F[v�q�)�e}>�V�)��W�8),A5M�uw����u��ev(�/�n���
#7�B�2d�L�-�eٛ���-LX���j�x�E8�@`���f�yĳ���G�1*�[�ƥ��uM��k�w�]B���-(�3(,̲�a�x����X�`�1�z��Vedw����%��"���l����w]�oCeZ&�@?�t{"��f������Y�p�* ��1��x��x���f�Ƙkj��TV�1��%�o:v�LЯ�w�J����.��;t�*��^BRsζ��ݹ�X�7n���Q��:����v`]��\���i�2p���ZHm2=�#�mu��gu�������gzq����V�*܏E�L;�&�ǐ�&�\.��Qt�@�!Xn�g����v\M��.�t�E��Fz�1�e���A�{A\ݸv���P�6��&�JۀՆ�$��kz�^�-�����[�;I��/mU<�K�'h�r�c�������F�Nn���@����|�5��^`�����%&yV2��g�⨾)���'y�a~�{���N�;�QE��ݰ�D[���6\R,e
�7X؀��?�6;h�h�Z���7������@����h�Y�'�O���>��v�$T�A��U8Dpc�g�ʅ�,�2`��X��⌔(Wj���R*�
C!����~i7���A�~"&&��ݕ��1t_��c������G]�8�d:v���x�rۇ]��l�&��̈�]����i!�{4F#9}��R����7L�Y��	
��������~�(��Z��6��k�=�������\�R;fx�;]Z���R����b��)��0a����g�v� �s���1V>�k����p���y��;�f��O��~�/Ab�	T��������8�f���{_���'�7��K7Z�vn��v�8{���Q��5f�Y��ѱ����q}�6�,�W�������̦�l�����g����[=�+!M�;��)���x�EW�2n7pm�#e��]���v޳d`�ygK�~��v�I*�uk{��gk!�7`3�	�gY�&&P��'�sY���(p�M�8n�v������V?{k�Q����l�f����71�4H"u�Ə���P��Hn���j�R�v��{ʺ:6��J��w������*�!
�
�R����XE<�Gn�)��7j񣱣�ZF�ϣ]fz�Ӹ��j�p�w��pA���F��0kojdE{�n��k/x���WV��*CS\䡙I�4������8"�	�`:eA�^R�B�����:N+���[��/����8 LF���K����ўk��k7\B3{��e62�9�Lz�꼂�>��o�ɥ�����X���Gf��g[��;����R�+zƣ�uص��{��2�K�x=�3s1���w�k�|m>z��J���=�Im
��#lF\���V���]Qp�Qd̢�2�!�vs�V�;�����n� ���_���������eJ���t�C�U�]���tB���2��e�Yd̢���<�6˺L;D ���b�ݮ���������q�O��v��o��+�1��}��Y'�ht@j�-��f�&�#��^M��v���ݺ�:3ź1eu`4����e��e�����y��<����{��2�S��:ށ�kn$K�!u�e�U�x��`���?�I�n�9�6�u����a%	��?�\�~��nl����dJ���}v����i�I�7�����nl�p�X�'��p.�87lݸ��U$�7[���3�2o�6��{����j���U%�	��g<.G]?[��?^v�������m.=�^�/q��=^�f�AT��^>Uܵ�DP���\����-	�r�h\ں�&y�읊�%)R��m�ޖ�Wf_�>�պ�^>�u�o��2��h����Hw��LG�q�`0�3�3!�i��Rp���W��=1ɘX�<����%�eEn��/WV���o]��v���~�_��ؾ��lAX�h�IL�*�[��3y���:�-��Ć��(�.��16��r���C��PNK ����A�p��1�9���ZG7ʸ8��/���
��/[�m��k�l�!�Bu��lA�@m��u6Rһq���[��:�AS� ���	�}#���#��E�p�+p������T�H�xH�3��
�v�|��-_q�w���W�}�Pp�*E�$(zB�E�9��(�3�,}��c �����|�Y�p-����L8�`�s_Ru�s�"��
Ȫ��O�����R*��7��"�B��>]q��zj��t���n����!�.u�\&e���]=���o�n�:qۧN�7��y�T�[�q��n�E*�c���l�y}�;��B���8��^;�5<{Ig�>ر_��Y�޼����W/�ە�ծ٬��ģ�w�Ϻ�m�]�|��<��Z��V�3�k�X7FR�I����:��:5v�٧9�Ǫw��q�݁f�V���O"��\�7�u�J#�k��J�YY2�B`�:a�9wjR��ܩAx�Tr�+z��/O!y�Y=�%�E�zI���Xf��0��ykc6�����`�d��NTӨ᭿N��7!�a�Wi�u�	�@�Ə%�f�5�f[�6�oM�.��,�ٽ�Eaz��v�_����`�=el�eG�O�����M��f`$����x��Ϟ�y[��l��L�$їN�j�V�kz�!wE���& ����;Go ���	�fBQ�(�`��U����˙�cu`oP�Y�X�n\��S���mu�y�e;ûnS��VG:v�։�Vi4�A�Kc�.�Wθ3�/���m�C�
x��Ȼ;D7��6��0���J����(�h�@PkK\iU�R�1y��`��.�'/Q�.a<�7\*�HA����j��u����m�������[Y٩v^�\hr	����*���^_udv}d��*�:B��]��3Z8�v뷱�ini����2�T���TT�T��$E�4�P\�Z &�^rR �����xe:ͧ�r��Ia�����\�*�X3�׬lkO��Y�J�S�X��{3/a���L�R��K��K��G�F��{"�p�u�;W6r�����ź�P��6���c�7N b��H]h,�l�H�-`a��+�P@z�iLDmh�m�5�M$��جiݷ�1 X�b+E@k1"*,i,�;(ܮ��1)(I�1��HĚB#G��*!
ɰU��a(�F$�Ęň����)(��,[��T���n[��r�X�(�6�,Rl;�5�U� �F[���(�@&1�t����ؓ.\��J��
�� �0j)6��V4[�2AL��cQb�7(0QcI�,X�nk�(�EEd���4�($9nr�$���(�m9tX�ưlE�̢�QPY(�\�h+���Kb(����O�ulM�B]6T�,��!�R$J:df��5�Mt;:Đ�3P�����'33`�֘��A�I(���iy�h2c�x�ӷZhq�ꛬ�o]=���=;�u�He}��X��a�#8I��0J��RpG�1r��������r`�|?0�ex;�Z��P
۶����Y��:�9	7��<Oo��ҏm�v�6z	��vh:t����;�0	��iط l.�f�,��2ٵp����m�q������ �\�D�դ+��+.�d��	
Q+JͲ3B3vB�J�]�f��UYXG3kw�R��(fW�6k�;aD�n�ģ���J����4�ř��.��N<�f9�Ò�t&��m�����N����G�u�3\�R��v�<]N���]5˸ãip�i5�)�]�u�[���K�;(l��qn�^�0p<
'��uq�؜��6�
�06�J��t�3Y�n%���zD5nG�݋=]�u\�������V9I�d&��Nձ�B���8؝�J�����-em�D1l�\K���e�Uư�(�	K�X�!׉<��ys՜�;�f��[�f7h���v^���Ѕ6l��%��1�myѶ;=#�=r/\����KTAUWE��ݭ�j�U�X���ۭ�GG^ˢ�K7#����Xff�i��z�W<]��sNH�l�⹋��4�#kN�^�҇HN�n6�ԍ!��CF�e�ܕ���@�U )5Q���!t6�ٍ��[��8��/,
�g���M���:)F�����b.ۭC�ݮ/Pu�&�x��m^q��tb��c�Sp:S�7M�]�]]�L��۞)�;<���p��ӔM]��[�3��l��o*�uᵲ��6@se��%�Xi���"�V��ܢb�.��玒��	��j�ru �0�t��c@���*ڄS)�u�7Uvx,r���$�`v�.Й�f#��x�\��=z���.X9�HM��z�f�nk7�E��LE�1�M@i�u���-״����t]��w��ܓ��u��Y�0� hԆt�����X�	��OuJ�E��(��%p��+��`���U��r]dK�qvͳ(�3��d1I�5���æ7�hv��P�<���d�b눶����<�خ#l�����ԛP��um/�=˛�-6��v��v{f��G��pQ1Y[q߿���~�﮵�n�ڮ��uvf���+���B��f���E;�=,����w��'���&TV�y���oro5�y�c�!�Vh�	3�K&���fer�2�!q�Y|��e�%]�����O�ok߿E�N�no����l�/\8+�-mİ��l�k�s�M]��:�ٙV[E��3*�մ��ȹ݉��}\��i��[�p:��sV0�7�a> ��l9�������ʜ
M����{ۢYD���<��n ��r1G�T�ɖ�t�x���'�8��*x����$��7l*�9��2��'y=��޷���n����*�9�E�y���y�\�u���Vz*e�Ȧe�D6�)�G��Z����b�V�^��ap�.�v�L��/�����d�g?��r	�n�Nw������*x�[��Q��ihqL1���A���A���fYd	�E���^d����T]����m1�fa21�]m��gT4�Əu3+~G^J#�>��'�[ޣo.b�ЋX�����K�}��/D��uߩ����X�qם�%���ر�v�w�&�E��!�;T�|��@~*�o�P�T3�A�.�#R�/�rS��Ay�w%S�d.�y-YV���	�`��Z�
�/H|�$*��~�!��;�}��x��w ��>]kwkmݹ޹T�<���`���7O=C@�`� ���!�*Bxi
���1�`u�䏳�UݢS��-��s���j��l�H4�m�Ǫ~��ٿ��<�i�E&�x��7[��S�^�Aˤ�(C�ݙ-����Q��;����U0���� �����dn��j|����_ �&Oz ɒ��˶B�K»�/	���B�H}���#z/��-6Rn����l��	I���mn��[�l`D�1"\:��ј�Я�4�wB�H����R/_���:pa�VW�=,l�n-��m�X�j�oU�jq�V�R�1Y�5SX.��A����3*�R`�N*���H�/	��5|f�z?�έV����=}�>?�=e7�m�2�!�W�!,֫�u�jz�ci���{9�`��.�e�9�:i�*/3}����i��*���v�?�=ޣ_�^���d>~B�>UBB�{�Zt6��;>zo�u�-��I��u�	郐Eۇ7lEۈZ2ۊs\��H�x/�w�#�3����\t�{�[WWn�Wj�D(�VU�%v��o�Q�]�Fϸ�]ϜE[�Ǝ��8��C�l�����3ّ����^k2 ���L�v�E�9�탑���%��@�0q�`׮�u��9�xͳ��fw��q�`���8r�k^>�l7>�����A|���>p����s붋�Qi�:v[�p�խ�M�חT�e�ne���!x�a6c��9�����t�����z_c��_�W@��v�|����k{α�s�[�>5l������ъ��_T3[%u4溬=�������r�t��,@WgW_:���0W/��{ ������WޒЧgʮ-�k&f&��ł����gY� �����pA7l�	7l!�Xum!N��p����<v���=(���W ��v��An����H�/)ދ���DVd;X�4 ��n�
�My'��Y��.
kf�Кgb������C�1�g�s��I��8K.���깄&�k7Ss�0��Xh �F�sX�8n܇��<@�5\��,n��#�������m��cd�V�xA�o8�87m�s��Xti磴_��q>a<ޏ�L$�A�q��)fps(��;YzQY��]�Fۇ]�	�
t7J��Lqҙޗ�x�
o�8��n���R~��n\�p�&�k7+��l�k�i���zw=8X������P�!�B���
�gO���w�K^V6֋�3=�J��άnV|��o=	
<2���b�߅��[7�(A�b���N�_u��}��ٳy}Y��)wG�;�,R��W�H[�a[k4fp)����\i���Ǎ����
�T���X��g�$i^��ޅ�V�M���]n|��s�v8�o���p�=�OE��p�fx��D닯�]���;���|P�yۍ��W[/bnn�ֺ�6�sۑ`0�^�u�\u���Ÿ�y{��gf8N��K(R�V+-G!ͱ�.�KK(M�ٙz�oSz�령3v�	����W��r!�w�AE�ۮ�i�'� \�++__����;jNh��<x�םU���8�����Qļ���T�Y�'����8�!ye��s,*�W<v����QY��qq����f*T*C���HU
$(S�g)�[��������A;��ؒ}��M��;��U�����	
���Aj\*�J����-�\�Y�R�G����Y����4�Z!���+��ٓ�X�M� F&D@&$�af��*2��I��=4��8QpA�q+�V���P�bfo�y�Fϱv��s� �r����ȇmI�$�AL�pnڑ��w%�M�ghc��[����͉3��N���l�.�9�e�7n[Gn���������c�g&��#��hWh�8��{E�V2u�I�Z!�v��B{ ����]�k!�%9�4ToI	�Nv[p!G��9h+�pB��syW�rg4I�E�Lu޶N;>�n��E�|W�k�CalۻT��X���K�J���N$�D��c5lZ�f�rw:d�g!Hj�������u��������+�H�W�Φ�;�L86W�����	�W0#�nzΑ~8���5���B�2L��Vc,͈~�=oO*�n1H�����[���v��l�pE�]���w�xlO4�>���oY�'�-M���Bl̮�nҙȭ+���E]m��޳����R`��9�fB��wƱ��q$���u�%�Vf��6\k����ȹ��Q��aU�����iL��%2�HcC%��Wu��.�1�7�Q��m>�5������}��?2p�O��Aݳ�$�6���$^�e�c��^=E�9
/�8�ga����.A�p����6l���Ŧ���"'[�)��B�^�[D[fe�cp �)����v�-q^7=v�pI�o+oI�`� ����	]����{���mA��,Y)q3F�=�!t+��t�?�Xۄ���,n�<X����	r֎[Y��.��$�7�i���]�oQ׮�V��@��RJa�qNgz烂j�8#-���%�F�E�BB�W�s3��v����輁�o?��g��f�gp)�|��`�!J\��T��X��f8v�]�r��9sڒ����_C���c��[dZ|����Lմ��
L��3M�:p6$���a^wۙ�عg.�Ҍ6Iu�l��n(w"O��i(�p߮����X9َݰp���q���60#�U�f��UBg�K��L�.N��./*C��Y^��:N�-�P�(P���r�Q����t�nX<��`戮�v���҆y;�o0ۇ�q��`�n����]��{����n��Ց���>�U
�B�٫΃�P�
���1��3�R�AV���`]�q=[��w˜��gz�׈["|}�'C��ºq����EQYvP����.k,ցu��Aں�0�i�1VmC6�L�� �ml�,i�t�Z U�}Țf^f%��c�0�>jie��m��8�	T(	
$^U~2���v=��7��L����w+G�����AT���*BCJ�
�Q��$��W�_@!�~���̍[�kwkd&�S7B��%�Xܳ`N�چѕT��J����� ��>�J�H��$?�Y���5���׍����]x��An�H ���m�|n�j��fy��6��kE���}V���^�H|�a��q�~��Ԩ���
�
��rRߟ�;�ؗ��|�;��R��P���Ž0�o3�<0]��1pln �L�lO�I])�Dۇ���[��ڜ
����Vv���Mi�2�����½B�o�TE����P�B�T�ʄ���R*T$5-����UmM�K;/���N��v�����8&������]�/H�~��暬`M���T�Y���)������������y8n�[���m�K�6IY���DS̝��*�O�dZ&e�ٻ�t�hQ���H������F:a���l�Y�D�k�Cً�]L�&�f[��Ux����痭����E�b��pjSV�1��P���F��,]�m�2&��`zv���k��N�X��뫵�/f�pi��s�2��љ2�ݞ1�n���`ڰf�]��T��4a�>�d��Sץ�8x���=������<���4�Z\4���.2��l��~���A7]0J�p�9^n��WvS0&�a{�hM���b�с1̛��[��dC�v�v���f^>et��vP���80d��j��k����0�Ys&����Y�FgFq0��eb�E�x�����?Y�]�-�9M��լM3�i���(���7�f�hc��G�m��nנAE ���;��ִ�{�y����cF#�x��u
���P�B=��B�>P�����=�f�E�c���	j!��y��gKo�tu�(fpc�p*�U��2z�����P^�ʪCWCP�K-zI�:����:D��wh��m6d�V�x�^cM���r	�gi���w}��˼�vq1V154�f�8�D��%��b��0uȓR�X���K%�����l�pA�p�J��w��q�_3�s�:Խ�3�ל��&L����C��md87
�C�B�/J�jsߣ���)���gƖo2i�e_�u���#�l5�����F��`�%�����/4��7��>���4�^]���a��n�`'���3�Am��MY[X+��36|\� ��l�E[�͙�[��#P5��J�6Y��<�F�,��e9�걬�}�z)���A(��i�':����L�V?����ݳ��$��:��M#U���91���Ey�w;��n�;��ܾgz�j�9�;��dl���a:����r���@HP�	T��g�?0/�J��U~����ݳ<)̡����]0pA
���`�
*^b���r�wٹ³����PhR���;�pM��:V�m�6����L��F��W��$��?������fȼ��[�5GM��feukq
��*5?3���h��5�z<nY�^�8E���L�9��]������ޑyH�5?.:NB�ž���� ��E�����҄ޓ�>Z�y\���ul!���fPfWg��\v㧇n��:t��n�7�U\q;�;���{��Y������M��:*�n�?k����Bn�(k����[f���5'+�Vj��oD=�DY=���(�鍼�Y}�pU��p�x�uwB�6_.�4Wh�cz��jr v�cQ�����rWk��i�3ygWcemش' ��ԍ���h���}���cα{���:XKU:�VQ�T�/m	�A�
�Pc�5��v �F`���vR��Ε�����ܴ��P��Ҧ��{��0h:��l�ma�� swa�w�xj�
|�����\����EP�?�*Y<�"��b������;�S�аn��a�����OL9J��}�]�v
3�	��ޔEhܝ�/��w���,�2�Ɔ�\��7�肦듎q)Re]��}�v���W<%���n;���Q8`-]�Ih��Ĭ�T���i����H�t����E�9˺���I��nJ���N�ܨ�ɀ���o}y�wW:e�]��3Ҹ���>7�����`=��8h's��s3�h����ڎ��j�fuǛ��Uu��֨�o��;L�N���S5��WR��&ٽ�g��hU�����4-cL�ihv3l^Ö�m� �-�L:��T{C�b�Ɖ�/�PY�,]�mf�s��>��>���'\L
�N��0���;9��d�u�\��믯�>��(j�Z�zE)/x�_���x�=�QnU�6���0m��̏K�*���[	f�f[	�M�Ô�$��K���"S���]=l���ɹ5E�&���w�|S9���S��B��V��	���� �+�!�lL�Ũű`�Z"4�0�X�H���39]*��mA��Eh����lh���b���ѣh�Y0�@1hюW"ɢ�`��F�*��c��\��cLoӮجѶ,h���EFH�"�D[�%6ō�lj��6�[%�XŬY��E�6E����
�%�T�ȶJ6��E��6��X�m��i5�kXţh�X�\�Q�Qb��*"Űch��͓E�M6�ŀ�L�`��X�����,N�+y�Ni�p�7L����6|��Â*�V"]M1�@�)Ð����!��]v���7q�3+�[�}R��:"��ve�1�EI��iY���v�Ȼ`�6l�	�3j���hp��p��l�m�}����
����/A2>�|>���e�"��Æ�MM���ٓ������֣+���[���3�ub�����������bݳ�)4-�W��xKC3E��8���s����d�"ӇJ>{�n�l�}��UR�,wc�-�Lp^"e��sa��K9�tͽ�feukqԻ�m�8*�b�77�p���"�+�4CHP��z,P���-�!�a���j�V1Um8��Y	��p�yic�m�VB�z���LW����s��{}���G�P�&��<n�We+ٽ��Ɛ����n�����|s쉔�nE{�fR=]L|s������էJ=��uZk#��9�r������˙:�xޣ���hP�-D��������w��.<An���^8�ʾ���v5��ݗ���e���2�����R���6]��t�˺~��������GаJc�<V���Ȅ��5��7M��$�l��D��}�/��LV86\v��h�n{\�evӋ����^��_vA��=}��x�T��I�fȐn���`�ݳ��M�g.������B ���N�p���U�|�!���p`�̭��@�p�6l�VH����O�Y7e�w7s,�fZ[�!��}���M,ѭ�5κ��dfR�[7MK9
l!�7l�kfr,ۀ�"oDj��a���h�pA�p��"�Z��Z����(���f˂$N�=�BT��d87l��l�Y����CL�����EkMB]��x�chfhc��AV��fAES����.?~�݋�Z�����N���oh�k���Ƨ_ґYNo��E�V����AxZ�v \f�����,�M]�e�ݗŻF�xb >F�Xh�4ZA�Z��&���Mr)�0��6ZِpG]3qUA�l��l4�V��
a	��	ͻ�5Vc�Et[��y^;X���#-�h��V�,l�s�Xz��ɝ,z��3Mh��B)��Ԧ͒05�˼[�۱��X�穼6�Ë2���g)X�N��iZ{nc[���{)�i�$M+csք��2�0�����MHXհ�1^�|����s���*��V0�SLCg.�:�GC�ɬX�#�,�:6��`|�'��y�_/�eݮ��k!�L���t)���̭��^�;��&�c'Y�����(O@¨������"_s�ߤ��l�<}����-�nj{j�]�E�8e�r.�6�sٺ��2xL'Ʃ���3[9ݷ���n��q	ƙڛڊEp.-��cz���Ñv�7n�UEE
̡Z��2�9.�O��]�ԙ*ގ}Sy����ٸ�Sy�VCU�
R���*��W����PEG�B����g�T�D��L��@�p��!rL�ssS�T��(���ٲ���.�?�'Dwp�'F������PI
m��U��E˦5�5��@N����y��.5�<�tu����ߣ�,�s"ݳ�]����OӶc(fpc���y�>�Z����FS��2A�p�����e���V�}�'�������s-�@�1+�i�K5ߘ��J��s���hG,>�������P2f��;^�*�<p��ݗ��%�1o|U+�B١l^�O$��@��V"��zg�M^dd�V�A�ÐA��붕R���)��.��M�7��v���0�u�QE� ��B��z�Kѳ3-Xy��CW=��\xBd�p�jˆe�̬��2��T35�oAZ�(�gv�>�s7-�v���e�����܎:�z\r�޷�k��IHjO���Om��Y�}��|��܅*�2�X�l�ۈ�"nO��3�����}�,Z�Yw�A����ۙyA!�H���y�
�$�F�;��}Wƽ�Io�M�|%�r�m�P�8�GyV-x�z�ئ�����j��ݾy'HT�U[�5YmS-���b�}�Hpw3c3�8�
�����0���3�u�|�5!�_��������e�bj[��I&S�X�sI�H�!xM��Ø�#�';W���}�
Z+]o]ֶfm�̔2Rؗ_P���W+5u�m��J����}���'ꫳ����!����K.�̶��jU��H}�¢����)�g(�V�[�K	�9,�f;�w��m/$�H��O뷹����%������m�Hhw3c3�8��O䓥���ϯ�>�?|����	��0�9�{���q�v�v-�t�O\�"�-�:��ߞ��Uߌ����Kg���F,{�����4�H}}ݡ�]7ww"�ݝ��=R#�SD���۬�57�2OL���\���x�[\��Uf�ҢsH�wwww�;�%����Oia,�,f�0
��}v�m^�
��w��-�+E&�ݽ�K+7�]F,zUW�a��씮��\<N\�mL_�Ed͋MZ�&�P��ɑ���ͫ�ƽR��Tn<E��R��EFL�{��T���ńd�}Ʌt�{��8�y������$�j�es��f�q
�`�'i<L��[�+��T��~��~B���*L��iQ�{W6 	��t	ĳ�4R&16�fW#�4��������E�6��[��.%�ܜ�l�Ȥ�b���`9���aܜ]��x������r�b�Ġ��U���+�w+z�XԪ��gߺ*�Z5`�ό�Z=֫�פ5R[��=���~2E�b�uB��\��z���ݽ��gS������˻m�Uoy�9�9���L���C���]ôT�{n^�{<��i8	0�w�ҩ�i.��֏�ә\ٷ�����U(}�ǻo]�W���؍�jT�t�Gi0��޶�����H��ƺ^���ݮ�N�>1��ek�G��t��J�WwLd��2+t/�*e�a����چ���5��w��;b
Հ��ki���ؖd�aѕY]
�,6��fv!ؤm�u�Pۿ��l�|����w1�
��;pnJ�hÊ*�1� ��	�v���/��j/F�v������]m��WOt��Pm���Y���>���nmlx,vI]��y�v�\��h���cZ�BfR�q���e��A�GAI�Kt9�r�rJJ�������m߁�#��6�����8t��^��Fd����詅��;��F|;]ہv�7�����K\'���;���N��F]e��ʥ5>p�y������j3`�;tD����T��f��Mq[�����͝�t��מ������m�x��of%"���/�&��"U�*��J�h�n�]����{ov�ؙ���LZ���f����{�'����^���l7;�q��^s���oXwu��p׏2��;"D[ȫ4��w�3'��0��$^�=r���<+?I�OЛ�C(7�7n7�j����Nbn��n�bIx
{/�7 ��S`���S���2�/M����g��Fsd����>4���p��.��@�a�z�ȋ��lh�"i�=�̉u���hqi	i�W��+,�Է��VaY��JX���]	�pͭ*���x!�X,��s2�;�Y4q9������`����6���/��ڍB��\��Bq����>�;>�`6�s��5��}Ƥ�CR~8��zW�չb��ۻ{�A�9g����[z����C���Y�Gwry�ɮ��=�ו���y�*�p�o����Glv!z޴��6������X�g�4����V�5/�W{�	�
���v�̹�ᭃ�g��!�8vZ�4bvΠ��ږHQ���h�pchX)�#.�n��5�����I0�͕�Y%{�ƄP����]g2��h`n�5�]g�ڽ!��]����6(m6Gr�esu�^cʹߪ���ʤ��u�a�m�O�{8�CY"��{<�\E���B�����u^3��}O4o{��a��)ͧ�!R�.��<"��ݽ���ɹ	�̼y�.Ғ�x��(�ʺ�i��+���ө����}����]�ݽ�M�ɭ��]�;S�ϵ��no]�l�L�.]�lE	���V����\�Z~��o�|�l.��v��l�uS21�+;��kZ��,yW	{j[�z��r�n��\��ϷL��gY&�*)2��b�α(�9��vM��+���Z륍���Fo��2X,k�qv���#W*�se�r]鴾�h��8{MT�z�2���Q��<��[���Y��It5��9z��V����YPA�.��K ��Q�p�����n�1֥��ekN��*�l��qv}!�"�ol�܅� =��}�T����^��z}v_%���}��WaF�.��r���n􉛫�5�2�4������
6;�W�)<�W`$,�i���#�����qk�Sy��Gݽ�iI��Xvs�]��awow�v�'�P�����Br�7gb`17�������L��'O�l73X@4!H&w���{	k]�;Z��n��rCm,Q�-p�,��]�T�mv���lK+e�:��V��%�6�z�3�ز@�awo�v����:��v��ë����oQ�*��r\2�޻��5�{s.^���Ӏ3X$��퀻�4��_k9��"�����X�3�WpV���<��`oq��c��\�0����Ww#�\2�gOuq����F��v2ʆ)�]­����<�y&����j���Ѻ�=굛�Z*l=�Z�	k333h5�N�{v�����qǧn{|ԉ$����.v��(ˆiv��l����v/ja؛�`x�U�{7���n�h����7W2� ��.�� ރFk����j�e�]��XzM�LeH6j�W�:��O s(��L�2�ߊ9d����#PG�r�P5�d}DГ8-2�ThP��%X�R�u�F
�x��-�ԣ�DN	�*�t[#�Y�@�50摻��^#Lѕ�-���/�|���k9u�ONނkt���W�iۧ%�;�n�(N]����1[j�7QAd�,c|6n���ያ�WՇu�u�B�es��{;.��s����1�{�y7:��4;�:�f7P����
\h&s;7��+I��aU,�2&Pl��SA$Y���J�'1X3h������Yv��#9W$���w���`!��En]�Κ�C��ӫ�ޛ�Fr~{ܟ-),$���I�ޡ}a`�5ԫ�ڵN��X���W-�z���<���r��_Q���G��ɝ�r�+�X0��ǺPnm:�j����C��d����ء�������Q���K�s��>��n�Ӊr��z�����Z����ݚ�3o$���cl�����m�L:u@��_-����Cf�-��QF��/��jo^�t��]�ݣsUhެ�QWP1uv��*�уn� ��t�7�p�8�������\�Y���em�퀣Y�i��3�j욑tw�zҌ̡}��^_^����ռ����,��2$Q�G�w��j�]>���"o�^=Qz�Xf��j	ey4�4�$�x��ͷ�;`��@�V�2Ƌ�U�Bk�7��;E6��L��e�w[��!n�30A8?�����pt�i6D�ARQDX֊��ۑRD���[rű���nJ+�(��lIE�����F���ƋbRkܹ�D���3E�[$���E`؊+IE���Y�˚D+��&���c4Tk�ՄԔ{�����f��2`5H���(���E�ѱ��4i5"��.U��ų����i65�2Q��&�{�CPk�F6�낡���E͸V6ɬb1Z,kٕ5snV
4BE����u��l��-&�4QRI�0Te�bw���=���ޱZl�2�mtF`푄.�X�B�Bm�ͷ��X�)5��Q�*mY�n�nn��p=n�����b�G<R�Ҭ4�u첅�Of�q�]���8�1\s�Zz����C�D�mNn����{�7M���\�6��]M�9�v���.�̰�5�sLin��f\p����c������Й�w�h��+Zɡڻza�;�z�uZ�k3ċ� �3J�����n�׋�۲>e�����dW<�lEK4��z��
P�.	XIM��W&��˷=l�s�M<u�O:YщݍTN�
-4%,Q8��;A,����A&(d,nh0̰�SX�u�6kc�ӑу-�)EK��UʳG&rb#a@���w8zC&n;�7���=��Cxvϸ�N��s�9lL�(�Y��(b���)���v�S�x.7�O&����yL2�,ЗYh��D�i��s�ۋ�r���N8#��64���]!ز{�ڑlŌt6f��)���j�n��ĸ�7\v��&0Qؐ��T���5�����w|���T���ېW���x����:�#^Nr]q�����$dr6�.Ψ�]v���s�l������F���v�-ə�{i^-#��ڴ��XHa�.&5��;+<�o �,�%�b*5�v��i�g�t����
����۩D�MQ��>��5��W9D�sa0۠�&�����;WH��n�wl �.z�pp��O=I�:]�S��c+^�^��b��u6�r&��y�l˅W��H����E���KZYy�F���t=��uz�^�Ap�-�g��unvӤE�c6��K�qrҝQ��3�O����v�P�U�d��|���A�E��ʴn�6�� �mK3(MM�Y��T�,n�u�l��Y�U7k�q������8��n�sˌ�\���YE��y��s�Nf��we;�-��\f�[&�ӧ�ۥ��CO7�������/mc^�ub�-�4�	٬�ݜOM,J�8�:�'q�&6��"������ێrt盉�611k�U֤�x;,�����u��Y�2�=�E�H�:��Ek ]e:�aŽ��e���CA��Ƈ<5�ΛΘp@��V�؈�v�zѠlӗ֞�p%�;�m�]�K�ֻ6{ ��A�ɡɎ�\FXXƔ���v�^u[.�-W�v�h�'U�f�\y��~@�ye�\遃b�p�ּ��tN2�GG����Š��][��߳�<�¾�m붷�	�غ5F��eǔ�*\{�z�2)&V�述���I����f�:�;��J�p�a��{�C�iȲ�W�����k.Q���G�s�Ѽ�ɂ>�;��U�:�/H~�O�<0e�{S���z��ċvWl\�������:ʪ9��5�����IHjK�sକ���
}k׃�
e��]C⫸Z�OXr+��%��`�n^i��,o*�J�A��N�T@�X�SWJ�l�v[e��LgQ�Y����y�￧�^��l2�Q��썚iTn3�84��UQ�b�ڿV��z���l��j��7]�g��O҅٢�N5;���gX��[�`]Qի���Y�+j�R;����d�i�ͣ`��׋+D�ݼ��㺣AڌěhȪ1ѷ�s[��og����߽]�%k���\g�w�����gj�F|*HEg~ζk��ȇ�A6.�,��U�-�a=n.��<E��φ��gnj��:����`�Ef>��ٶ�B�:�Ql�'��o n?D\	�𾷟]����ww�u���cR�2���Uie���������t>�d��&��ߩ����]�~���O���-�)]+
v.ϛ�G%�cB�8����aW�%6
�������CO�H��jx2��,��r�e4�f�}/0�T�������$�g�Ue�>����n�n�W��}W3\g^o���Z�__�1!Vg�h���c{�m��{���}��0gU,d�&�*�w2�"#&�"�VTb�+�F�%��S�&�{�)k��Y��t�];�[��Ԃ^]\�aVf���ʁ$TfQlYo�&-�(��켸�ݸm�v�tTS��=�v�o]�E#:/��2��Wq�Q[1T�-Ô�k�ޙ݋�{�wv���v7����.d��������.s�8
��l.��d�{t����eU��ŕژ춒��lL�X!.�J�[�拑F�� S��:|�2��]K���bⲊ�oD���#���R�www~͕�Y��y�_s��+F�����w����?���25�77h�`��y�����l���-zʱT��=� �:��W./n��V��I�n<m���q�qp޵o��:��L\VQ���O�M�f�e�	�]��|�^gfL�íU-kg5|oj	
\]9�#Wr�����-̾��鿳��Oe�Ģ�Qכ��n��:n�룅[x]���wxTz넰��\fP��~���9*�'@�a�]�}�uI���}0�@��s�	x�N��A6���n��^%q�R��S�8�t�*"��S�#5���od��I�ק��n$лeU�ANs
�z����j�������"��}��:/h�k�J�֥V}Φ{�
k(�����k���;��67�����k�w�4��h�T��`<�Η����%]dǷީ�?�u8�o_�����ƛ��Ƭ�̟]�j�W��7ή�9՝�Qn#�(M�{i����	5�=�1����r��&�*������5��2��+�±�2�]��]ߣΫ�s�n~Nozpb���y+x
��S�]uܶ�I"D�ۤR,���kAuY=�V�Y�/�wVh�8�E	�jQ+A��e.��z�e�μ��#�}�����<�yq��K����+�p���b��ӹ$}�1����n-��k��&�㑹r{�v6箜f뗴,�Hd��	i3���f��.�vz6`�ԑػl8�<���^�sHD�7R��B��ڼt�n�f�,����N�s�Nv��կi��'c���C��:�,=��0n��hKten݋��]�,f���Dΰh�xY�lU��J/��W�P#���7��z�ڊ��x��2i�
ֆ���$���ޟ���d��v����`C2�cr;�3J�uc)�����ᳲ�~���*���%�I������Jg�7u�%[�5Ԛ�*s�8
�q�� ��Z�.��˽ګ�O�H�5!z�����R��w�������J������	'&l#�f;�b����mun5q�Κ|�cJ��J�����<<me�n8�7n.�y'	+�۽�;y;zYI����m2V�s�x�.S�n% ]ǟ}�+�����VAu�	��6� 4��ay���T�pͫ�07ZK��3\F���7�ߟ~���^M����V5�NI�����7�q:빆u���X޻������g=gR���YI~���Vb�V�����c����8(b����<�ɱ�ӕض���1����&~˝{m��Ȧ[�_&�&�g/�YޙpjZ_3f������U� /�Y�*�̞Zk��ˮ�!�*����/̸��s�:�y���i�[BΝ�&-�X]��������R�-�k�n[�����e��k��=�Ƶ����[n���m�*�Os���v޻��n!�kA4)�n,8����Ԅr٦��.*�d�Y�*�H���Av`�ӅL���
��E�.un3�Y�y/3�ޔ�X�{F�Xq��E���w^7��G���$��e��gqku��]�u�[�[ �eL^:��`.�����5�}�wQц+[=�͗j�_x)/]m�79'����U�̉�ڦ�����<5��^���?���kk.~&ν��J������Un�e���4(|�B�*cSP�0��TkOY+SC�͎eb�h�5����f�&�͈{B��PJt���wF������?}�*ə���3��$�9"�Y�`�F�[N@�N.��/ص���,�u�:�z����b�^�5��C!���*��i��iDSTVYx���Z2MEs���I]޼a�wsv8���n*�,]t��!��]�I��ݶu��1.V�7''2���nm(���Zȩ�3E��߹�Z�퀻��'7f���8��U�Ws0��jJ�N��������m�`ُo�P+�z��Ɂ�R��O][�d��x	���}q7&�W�ol_���0r�Io��"�t��֍��f<��d}�{�x�-����]�o�t�u�s���swn3�Nv�76�qSr�#w��-��{��;=
��`����*eX��2�e)��h�x���<��:�1�T���o���+R�ǥ��s�w��'}Q�,fn�n�Op�lL+�m�.�]���v>�D����9;9��K��w�_߽r�}�:����O��?~���� ]F�)[��ԋ�ºjmY�6	n�t��,R%6�F�T� )��Fj���T�ޗw;&�CM)�������lp���d"�9���?/HjC�+�<�I׷+Y�_�l^�wh��d����ʬ��oUs���Qvr;���]�k�p.ٻ���74Ś��?K햢����������2I>��.�i�ȿgc�k���k�c)M���b=�=yc{wr�SS��p95�]���n�
�LU)�:B<'M77qsp��@�oW\�.���o_�=o3�qN�#���f�u�&]���`�-�z0�:m����o�zy�~��םR����yc����)0�$���Õ�2�_���Se"��ul&�
�4Pz����F27K�󧞭i�ywமg�0�n���92�*0Yr�R6��'�]���{0���W1onBz��+tv�'%�$KX�s�KŎ|�D_l��.^�V������kk{&q��7+��\	�s`x�n�o:��;�m<)�v��Zx�(���!�	���qls�]���%ﯿ�6���}W"A[t�ֹ�z�)53��7Ba�-4v�b�Jt�$y�;��}�{݇��/Hh�=�q�z�)K�%�;�[ő�~�y������Q�L�xL��P�B_3e7�	��k�iǊ짺�G�{e���x�֖g��k<g�Bj�p.���w++R�spe\�Şa�&�1m77
�6����B�	/8)>6;TC�,KW��齖���l�b�n�ĥ�Ν��wwH���z��H]�T�K�z?������<�K釿|o�ϻ��<�boe�ݸ/<�m���������������V�z�D6ITB���F� �Vڕ|^�U3N���_��������1o�Z�b�cl-[ os�z�l.��w~�_q?p����Z��]NⲸ��.uj��2��ysoQ����brպӹ�l��m?9[�\!3EK�퍅������&qˡ?a��	m���W�>=��vN�FJS3�xD[ǖ��Wd	�3:�q��RER�?�RQ������|gkf+&�-7_M�wr.��,���������=p�iq}�]�[m��S��F�|�ƫ�է�~:��5$U!�$�Y�$�dv���	�ɫ��ͨ�J��ft�z"��Z�ݱ{��}j��a@r]��:^5��$�����c���qF]���]gA4D�9�v�����R���WDeͶZ�?_ kqx��ɛ}踦�۳��$��}�5��x�E3����n6��g�����qI�}Rޮ�b��9T)i�z�;�|=�fQ������oo/oN�]�zzzzz{=������gW���kiE�sY��!泧C&RC�5�i�v�^>��s6�\��1���`�us}�u�#�%�|�N���lw�̒�-�t`�J���%��+Ű�}��ݦ9�Wuv�����l�3��;���A�U�#wׯ6�"��vЖ�y��,�-�L�)��Q����ƛ6i����{J}K�d�Y�iU�=ie*o���{&��g\�7�|JѶ�31�[���y�)r۠�,K��j�$����(jڐ^PY9�Ny�_5�vV-q��U��F �<�o���eTz��v��P7ٕ�x_�^�:P���0��c0V����t�d���uũ��V΢��%�$u(.��2�nbd#��oS�Yy4C��_e�ɻ��m�yD�F��8���̍�oS�$�R�ᓮ�V��V��%͙wĳf�/ ��՝�3eu�U��R��v��J�emfg���S(f�cXU�� ;,��j��9Њ�q���H�.�T���Y�Wn�LM�,�t�*9�b���+}!f�\���*��+���g�'*��z�\�AR�_ƺ]�`��T�9��9�R��q�Z�T�푓h$$��p_L;&tv���cD��v;T���U�7�m���Z�NTմ�;���2�.�<�Jto�ފWRk�QT��e�cRB�M��[O̦��h�6��,%z#1�k;J��3�t�c�K2�4)+���5\yw��:�f7�Y���8�n�|��(p`y#"�ج�/5�p��w:-��g^����z�ab�hyZd���F=Y�blP>> <A���\�cĖ0��؄�X�������E�p�E��r5�"��*�aI�-�d���梹h�%��Hjw\�L����4`��s�9Q�<���lmݝ������ט؊�k�5ͮh6���_������ۛIEE�\�6����U淒Z7<�<�P��#E�9b*��wnݷ��b�uQ�F�F�c��nm	D��VcY�/.2,[h�-\����Q�Ou�ͣj���I�m;�h���y������F�����W�\ż�;�c�y��0 �1���]�n��\b�Q�67��ʇ�M܁7ov�͵3�T��Z�!�G�#��o]ҥ/c��tFT�e�봺*wY'�$y�{xԆ�I%�����g`���������ƚ�%����>o�XW[ݰ�G:��5�a��=�}A� ����@4{6��S�%�q���%��(qq�u[]Cwo���Ǐ���ƻ��eOV��\d����:7�4��c�^��]���ݸm��{m�I�ϵ-��7/\v�tF\�e���bol6���2{�4�=}~[Uׄ�CRKDq�٧��/��9X�j��z���3���l=v޻��Bݧ�͡3
9�w��;7l%�N���(�E5Z��#{�	�y�8���q(�<��z�IL&�)��TA'���,aXgob˾���V�IX����؁���aKF_
.M������݌CO��UW���8�LOw� C<�lv`%R�#r�v+.��u��e����Ό$�??}��߂|��jB��ln�rk��vq�է��B��9��F �E$���a3t��*��!��,�0��kG	~z�����@��ʹX�_�^�T�H�CU�Zv)��5<���{o�jZ23���v�:7}ޙ���d�q���u��v�v��w�� ʦ��r��K鹯�ΗM?�����c�H�-�\�-�x�F�zy�Qkg@�?�,`.X�W��ڶ�.v��>pLl�:��B��P;��ofǮ�[]����G_O3
ǟ.o�_!��Wk3�x�}ƻoI/����_�v:ʟ�\���a�~��j���%%t]0��n�%o��~Y���F�Cj�}Df�G:��7fMsכݿ5k����va��#���`d0�Ŀ�@2��3�@-�Sli��0�ͫ���nM
�Z��b������
�G@2ە9bn3�Mn�yy.Y�#<p���ͪeǵ�Y	�^��C��VnmJ�]p�+�k�|��U�tJ&������Q��7
���d2�g��u!����Fiy,5��4�:�b��l��������P��ع�i��Dv%�����Mc�Ku�ڕJ�GDƚKr$E�X��7n�+s��G�j��������z�UC'�<�����Zn��4�V�,��m�C{��(z���wn"y�3�͝P��z�\+lۿ=W.�&wº���nɦ9͒��ӏ-k���]����|G� *��r� !���.��Dc�q�ڼ}mo�]��C��0�^�������xU��S&�=�5�F�Zn���c9m+hSy�"�F%wv��\�������b��8��=J]>o���'�V��Y�W�H*��a4a�A�l���֙��V١0��6Fm*���/bTA��)`7]ہv�1�Y��Љ�7+wS
Q� [��	�usB��Z�"�Zo��%A&>�oof���t��W+�yh�����:�=y�
K�̩ik�ޱ��I��gf������3�0m���9j�w7
�)I`��%� �ݝ����,���{!W]e	�w�
˻�۷$B�� ������v���N(�]�c�*G�N�f;J]w�{޻oo��I�awoةх�7����1�Ky����nV.��"��So>U������W'���IL��/t4Ֆ!�մ���y)��6Α��f6[]��]�&G��f%��$�a��]�"�\�����\u�Fz�i��ޤ�ў�U8X�퀻�Ve�ҡ��m�]�&�����o��~�����E�	�.����m��=7��V�_((�X�5��Mv{`LՑ��������K�Szn�]�g��ށ�7I��<�DZ�A�"m�G�qɼ�������k���X���Ge�狭�����E[�����]o�O��S]��a!��^-5!��EPf�	0�B�M]%9wf�=�3e�v�]���什R�����w�`��2�m�t�ު`<��LlT�V"[���RUHd�Ϸ������o2w	��6QR�v����w�Ԝy���XE�wu�}~�gi�z�\���.i����=p�m���؂�6h4�h���u�~���C�d5k,�����uf�qq�����6����m�wr.�z��,[��������طĆ��2�u�:l�
���t���F\��>TөƦ�o]۟v�_s��/����r�R�ѽ��S�v�me"6T�|�9�O��	~
��Vue՛jK[��d{=�ݡ��u���P�f�Ӆ�A���J͵J�=���3��4Y��iW�nfe �#�hP��hQz;���0���3]�!�eL�y��7�tzս������ki��۳�P�*󊧐����8U0\�]�݃bz�O�?
5�}���Im�C�I3C%�u�0=اT��(5�`�ufI�[�F��W������޻��a5]���pfR�Ѽ�������{�8õ�wwm�Ժ������f����e�|��1Yܬ�˫6ԑ��f0mwr#Jݾ����\��O�]�ÍE�|�,?�J������}�x��~��4}$�+:�V�������}��UR����=3 ��KF��� Pv�����uJ�wr�􊼡�@$^��i}Y���[�����y��f�˻ԑ��f0$�U#����ʗ�!�!�7X�[�s��Fr��hѳ8���;�E�x�cS.�ز�&+s��д4b��>�)[�:�9��л�M�w(T�| �m;�Fe�Jj�x@�.�e��Ue�4zXx�$���:���B�0;�踎�'[q�xwq�%p�&��Ql2e��`4*׳g���۶�MC��l�d�����f�_9tU�A��\�Ul�ǣ��xι��js�ט沤��P�4���A��s1V�u��۞؃�nv�	��pq�9�a٨�Llc :%ҝ�H���+�K�����5%�4�f�F]�E�a��sm�r����5�S�=Sl	T��!7����}�����[��u�=
��N�TK�CZ��u�m�]���^>�	�g���u��ޥyǡ�3)b����8����D�#w]Sxm�z���.�=����ΒG�v�Y���ĵ�yved]ہv��[tHf���v�[��������7r�{����})���za�6�fSxf����`.���i~�!f�6V�R��^CZƵ��x�~M뻻����~Y�0�${?d�L�(��tcŨP��b2�6k�h	Mm����9M��QYwX�_#���Ͼ٢L�Sp��|�U�v%�#˟u2`��U^�&@R^�׬��o]۷��]�c�����,w�X�[!�Z5ʠjfaܼ�@4.�tn��ǖ+�z�u&�\��g,y�:ؖ��]t?+��w}Jn\��ܽ�u�+�n�j�3zf1O>��V0�%,U����*y�|MoEU�Ԇ����,�c��I|�c��Z�kXֱv��n9]��ո�)�]avDT:�rgYxt\\�`����]�۲�����ڿo���Q~TN�N2�"�L)4�59b��U�l��vИ˦���?�`#�j�j=�Z]1$��`���ю�V�s��c3!�N�c�;.=va!�m�eh��'���d�\���I����]���۲|���K�t��B�m�F]x-a������ܰ��c)zS���Z��x��������H�/o���,�C�P����v���ͷ�܁F��K����k��hFa���UC�4�O,{�vki89c��ӛ7Kٛ��s#����N��l*�y���j�.�Y�=(̃�v�hv�����7�P�L=�������wo;l�ty��RvN[Z�lOV�gi�fX�.��2}�kS=r���K���.�]���#���.��e�͝��*�.eؘ{.���z���F��oϿ�����
��n��ij46��3k�k����M9���`���G�Cס=N<�|�I�I�b��ySp�Rc.�4T��^1؊z��=�\V7�n+�,��/s[�r��T�3ܜ
���۾�,�NS�X�7�x��on0K�����)��zz��n!$�I��h��'�!�Z���VD�5��e�b`2������źib�+/�.�o�^%�x¨�F]2�C�+`4�]l�,�+�v$/���n(���s!XYL�`�6�،\eQ�.�&!�k7@9�Ceu�v�_/�{�␤���u��awn.I2p�[�\O෍=��N��,���.�g��$� ]��ݲ�g��5�o�C�<������9�ͦF��Yv�$*�.7(�c`���ċ��c��.��rݖ�{e�>NC[���M��ω�6�ʭ��aV�V�Z���øv�lDبa���|w���m.���\5_��bR�,�ڬ&������y'I8J�
��c�9�F�!�NVJX�g�콫�v�����
vD�Q��?��mM�L�����rZ�^��&e��b��wq���m�wo�v���Lٷ��;2�ɚ���6|�̼�:����O��_�Gࢪ�ժ������" �����(��`u��QZ##����L쵙����k,ՙk2��Y�Y��+fmfm�Z�6�-fZ̵�k3[3k3k3Ve��Z��L�̵��3[3k3m3k2�c-�mfZ��̵�k2�e��l�Yf�f�f��l�Y��6�-fj̵�mfZ̶̵�m3k2�e�ͬ�Y���k3[2�f�f�f��Y��6������2�eY��*���ՙ���l�Y��-fZ̴���
5O<�
 [Q�*���*�0QX�c� �LQV0X�cU� ��cU�V0X�c �0X�QcE��:��E���-1DX�cE�Q1DX�cE�Q7�E�1DX�cE�A1X�cE�<]6�,b���"��
,`���"� ��,`����,b���"��`�b�`�`�b�`��q�H��H�mfkfj����̵����-fj̶̵�k2�eA#����drO���� ��"��b~�m�����C=p~���?��
���?ǃ�z���pO�P}�U����Ǯ���*���>�������A����������'���S���k�C�UE���w���KH��u�&��a�	�@���}����Q'����,T@duU֫�QmU�ST ��E`�DX$ E`�DX�E��`�*Eb�Qb�`�bE`AbEdQXAcE�P~iEPx��J�寂����"��� �H 3�=�_����}� w�����{�k������}���G��~���	��N���:��C��p{�`��+����'�o���j*����TWꇼ����APEk�1��*��� ������Q���T?�+��=�g1��, �EU��?O����*���1$��_���?��O��{�{���?���4�����a������`����''�l�g���9>`J6���G��t����&�`��+�PIX}�>���a�\]�'{_j"�+��xPEz.�����<���!�M��1AY&SY2i"k[ـpP��3'� b�>�         >�                           �  ��   �          �                      7�  �T �$�P�(�*��JRUR�R�TU�IADE(�(*�D�	HTR�Q*R�� 6�E ��P�R Wx�{�t=�� s�Ҁ��a� ��*�A���@���{�B������J�@\� ��=�    7�  �G��@

�����(BK�<P'��z ��������Pv����W��#@z)ΡGu��;� =���{��@    o� �"�A
���E* !Q_{��w�x{f�� �{�@���P.u
70:
7s���6�4w��"���O[gz�*Oy�� 
.�  .t}��:�gZhy%	���l9��
�ޱ���;׸*��
�c��/]�"l�w�Z <ڀW-.��   �  ��T� �%J����QOy_M+�4�^l �se
sol+@��
X����ѶW;
u���H��M(����{ t��    �  	��h� 'U�:v ��@@�� `�*�� ��: 4 ]P       ��U(��P�QB� �=7w Q݀�gEv ����@24
w`���*�� m�      ����΀�U�
������ �� g*�. �� � 7`!� `P�  }� {�$��@
�) )Q> �} 1��r wR�:�s�����Ξ�)�[�
�rzI.zE'�ȥo-ԥ�]�    � �r�}wBQ��w
�� ���5y��
��W�Yj(�oRR�u{
�Y�^a��2iT��4����Ɗ�H��4i��?M���   ��eT�M"�!��M��	JQ�  I꒕O��  ��MD��%Ji'��d=������?���I?Đ�|?���Xd�q�r�]LM��	&j����H$��խ���jڭm�u[U���V�BH�	!!�����=�ow������h��p����MmK{�負�]��ۏMP�{[A�eh�n�R���e<��B{+M������%-����5GF�Q�`�E��[��jB;{R���y8@G&�;+/Y����11Oef�իI��¨e��#{���&:&���qF����y���i�&�����mTpU��M]ȥ�%A�����W�LF�|��5a��2���4���h�D���Ei�w`������]n��"�J�a°aõ+T4���S��Jɥ,6i�ٯX�/#V�	Co4�7b�l-�d���5���n̳w��ΡI[�ѡZK��S��Բ���$��^��.U���.�&�2��qitD�q���[YxX���&���Iռ��̈́���ګ��6�Pi��{���&�)�4�Kc:2�L������F�:�ޥF����"�B�яm��ޖ���Ƴ��K�V�X�����=�`��rU�I���o寉�v�,�Õ�j���^T�j7Z��chl��z�)�x���lD�	-,ryn��S+p4^7�V�ӧhĝk����k.wd2F�TV톎UB��ٶ҆URx��NT�G^֤�����^���׆��:�ڳ�j��ս��aŁU�;ͦ�&L���{7C\9v���R�V�:�S�����x����R�c�{�p��K�iDD���s�kva�ӽ�B�!�q\�vV�����PL���o#��$�e�B�8�W����.�nn�h���� xt�S2�W��Zi
љ{�V��*�S*#Ye��I���{��t�t�e�OFTN��ǍE��pس����iB��\5 ���J֪׭���0���Y�K6�ˣf�;�7��vBx+v�,�T���U�1�{s-^8��G
#&\6�RV�+E�^�!����31Xq��749L��1�ߒ��qҪ�뽉ӻÑ+%���5LRh74�ɖ�WB��ڡ^c�vɣ�U�S)f-��ʽ���g���[c*�vj��MM��8�%BDx&7m�lP��#T���ݣ6���*jĠ���*}xf����b�Ίp����U����(	������̈����Eb�����˴Ҵl� ��b#SO%�������p��HF�t�ȉ��$���+m(!ͺc*��6/>�`�����	��˦U��ZU$u5V�EX�E���uU��î�ݴR�v�����xw3�'"V��܅&�U�����nU0qܶf�k�*�ы+TA�x3E�L�J6Ha�7v��������Zt)W������pԴw+d�we
Ұ���ɇ�GE�8���ŔQm=�cSq��mK�H�r_�2'4���OT�2��:�ՅT��/sw(��>����]�_]	�X�Y�qø��٣6��u׊�i�*���e�F7GPP�z�-���r��ү��.�R�x�(ҒC��X�a�GwfV�JL�ԕK��{�����յB`�Ņ'b��QUgmn�E�5�3�5�ކUl)��ň�/)�9y�Aj�5�.�*�_Ee^����E�I����e�j��pn��jIR�r�U�hҞ�Q�H��;�V�R��(��kD?`����.��]�b�U�*�U�,c�u�~�2�R�g�����/���H�@U[vQ�;��R�r��E�E+�7���&��A����ǔ3o*��dBJ�m��0��R���:fk�t$^U��&bckcJ�x�D7H��<�vmR�yg
�WBU;�� ���B����ɭ�&Sw�m [���3����{ׅ�ɥe�	5�jG�$v�P5���2�"��e�Ĳ�U�j�m9ҭ;�K�4B�`�
��5�^Y��!&Ԇn�z`w��X����G�����c+&F��8Sl-��p'�Իi궘:��6��ژ�	��H�c�����xض�j��2��m��]��w1��{1Z,���NX�s)^�T4�T�2*gv��,a����ɓ5J�5Z���C� �U�ct�ӭa�zc����V�4/���I�SC7Ah��	je��Ռ���R�ͭ�KmQf��ܺ�jv�^�dZ���͔f�F�<;��ۣ����Wy��ŬU�3�[�f��KlV6jM��W�TF���`�۪V�ŷ�rL<8Q"^cwo5Vf�Ң]�i�I��٫�Zl��	Tq�V��9):�{�ԡ��TvmE�Y��Ĳ��*�e�Q�U ڹw��y��f��]K�,���7�ͬ�����#-XM	���ej�'m�3��OL���j����W�-"\VN�S6�,���w!4.l�����{�����Y�]ɪ�츨,��*1�Fj��w�osn�l��x��.�he!0Ir����"�PeK�+(���J�ei�8���ܸə�Ua���1�ˆ�^�m��ͷ��m�&�Q^+�g 3wr�ٹ��z�mk7A� KP:*RP��3nmH�.#�Z3�WVj�B�33Y��fG����tŵUJ��]�YDuy[��Z��IA�M�,sF
��[����K]=�J4J'qTU�\�'kNdL��v��]�˪����]���VS���&�Vv����tU�����K`��v�e<�g,7u�J�b���u��tP�<���S��j��Z����b�ږ6��/��ݧ�Ty$`�^K�l�0$�jR����:�l�T!�K�3JL�J�㫩q��z]+%�7Y)*{W����,J¶�ø+^p����(��f��sD����c w&�F=�m����A�[�'(�Or��e�	w[f+sh�6�Q�t�ڭ�I�^�A��Z,M�����Kn�WZ�c���TՉ�N�$�[���!e䠪���^tu�5x�Nf��>Ŵ1�Tf�O�Z�^m\�ڏw�#�
E��QC�ɴ1��3*�7+�yf��,d�4}[%��g6M��r�Y��Ii�L.^��eji
�:-��W���36�Z��KoV�rƨ�	y{q����\���xKaV�ݘ�k��[���sK���BZKz���xL�f�7T9F�ݗ��镚�5CN�*�0ٚ�U�Qɸ���4Ч��nݔjn�{qܫZrN9!��MZݣb4&e�m��fh�crD++5�f[x,�l0�I%Rë&�l���.�4	���v~b�ݔun���6�9�c�i�V-Ct�s�;�)�mm�o%eK���n��_;F-�K�A\f�x��7���[�ە�x�Z�H.��,��h-�Z�{:*��û�ٷ2����]�;V]ÖF��;�r�ˤA:�[ۺ�RG�w2�ѽ�tҦl7F��V�ڔwpʛ/n��ڡ3b���DKtFd�V��+n�Uk"��YZA��t�r����z/6�ɹ��4��,,+V�^HM=��4UUUL�ώjz���7p��x��P2Pv�d�a��ܸ��-}xb)�:,��w���ǂ푪��ʪ�&�͘M�(�w,:�K�4�m�
Lz��-f3U�p朳Wn9.���E�<w0��ȫ�Sm�E�u�iKTB�fX]jm����ͺ3(3�iP�	k�s
�7^��M���"4��Ȁ���lI�đ�Yޭ{�b�D�ǗUv���iM�ܻ�`���0�*��=�V����O.��)�ڰ��ѧu�dQ���R+2�ug%Ѩ���*���)<M%����v�f��i�UH�LxP�ZeVc���Qd�wY��,ӆ�;#j��w.�=�N+�L[�wma#���p@T4�$A�H#��hь��j�c$5dn�Ķ�X2��4�S%ҽY�/.n�հΓ/Yx�9�X�Lk�-��kl�G뤩<��ڪe�w-����۫Y�A���f�L �U�*����[JP϶�Ӳ�_�RY7��Bd�.���۽�cmB
���*�t�'a#ٷ�7ê�^$3�u),�(5E%�؉'*��v�p�Y{�c�ړ'2<�*�{H����R��cek���w`��>�{�'�E��������0ދ#H��G�U��ǐ�T��JɊ��^=cA����Vnf����P���XdB�f%+sv����b���d�F�c�����)��owtPe����s	�5_�H��(8˚*K6q�Us3��Ԯ�d��v���f���}0�m�X�vm����*�?]fc�w��Z{e�s�����T�ԫ%<Yq��f��V���T�ʗ�+*bd��)�ˬ��c&�Zq�W0���-p�4�Q��kv�J�1,?Y�
m|T{�0`r�JWu�墬:�`԰�w
I8Q�6*!�lf��#4�ʽ�B�����H�[B-˴sv�`�(���5X2�AL�Y��#^忙۱mp�;���N��p�
.Ʃ�4��֫p�Mc��W���ܨ�w�gJ�M�+Rx):u����
��ͼ%�Y���3 ��]J��M{R�.��gBN[���ģ"2���O�	��-�I�쬩��ꞿ��:Y����4��34Ҡ�æ�y3m����٥�`ז^��y���d�>���2�7Qں�H
�(�XA�����,�n4�
���ͫ�BUm˶�΅جvX*�ȉ�Pl-=�-�uC	N�8Wΰ��m�j0m�[{U�]FY'B��2�G�U�p�:;��U���Z��Ut�.m��-[bΨ�A���Jg�[��-,	gd-M��f�a��yz�z�����KT�^�.�}sk6�WgP�_��������aj�T�PY�T���hi�j�7�Tx]U�w����[q:��7-=�7hT��De�bu�e1*ie�Y�Q��SQ�305w)��J���5��)�gV(m����gBXB�l�3���p�ܕ����bXA�GQˤ����j��]�������K��te�8o�Yu�j�C���֐�&^R��]R�y,����X�6��CܼkpLa]�h7�ddC69uE�"Y���WM��ӡ짴*hܓkl���Yc4TC^�b���s��nB70ѷ�����<6Ȑ#{��ujdr*#75��ԭyf�ۚ�w�G.E�0L��o&������F�Eq�Պ�L�F�A�Xl���D�`�&⻀���հq�=t��Uz�Y�TK�k���י�������*�M%J�]�C����
������ݬ��yf��r�1�6�eT�������5�݌�����]�d�iLV�#��8I��+^-�,��
�YoUIU�Z,T��锋�k6CY�D�ʠ�U�ջ��M����������JQ�c�k甮��X�ļ�p�4J�Icڴ4��퉽��UUq�aLQ�hk���)��n���@�B�h�R�)�U�E��&h�cUoC��UM^[�r��P�2��Rͱ���Iz��X�Ҏ��w3)���|~R՗�KA֜�-�4��ى7�z�i�YXN�M�4`�j�%�2l�D���4�J�,ё]�ygk*(\.P���OV�tA�J��Y�2����vrT�����͝C7&e�m����&^`��l��f��ţ�R�h��vdmވ�`/q�`��.�=��5�XQG%���ٵ��f�N�f�]3�nVڬ�Ph�k1oN�$9������� ���QFQ���f��U�_ْ-B�2#�n^Vc�����F�#M����D��d�D�m�'fɰ֬үn���M�od��Y�*���1�O��Ũ�.���]�+�BGs.�Pa�{zwbAQUor+Aji��ʡ�mò�͂��o2�V챹t2����c[u� ʢ�&bÛ�&��;�*�]Xs�K

��7�է����ff�+R�D�ncwS�r�I%h�5Y*[ɺ���V��Da��d�ʻ�E��h�*�h+���u�$��6�qGH�a�Ҷ��n��,�K�W�B=��D@��j�N���˺8��x(ϘXX�I��[hA��XZ�c.Y�P�M��P;����l���/дl��C.�ݲ�7V��9s1�6�f�4�I�f�D0�2��cYv��{�I%nݼ��c4�R��Kq@��5�w�P��K�P��)0���Si��1�����p��VR��`�UJcj�݊�ʠ�ʧEVEJd�G5c��\̭��x����R�U74C̳f�m�&ռQYI�8�9��s�2�g7!D��L���8�ެ�ۖ32��\���n��+4�<�mYպn?��	-M`��k�3 y�j�2�卽�!6kr���\���l˨��ݘX�(�S6%�F+W��cJZ��B;[��W�ùz������b����ڢ�f^���u����ݵZ�B.�l�f��쨛@��9E�f̻ÏN0hiy����uGN显��e�S�ܼ��V�GZ�r\mlQ��Ŗ����Yq%y�s�7t�<�v��B�4�d;�dں��L0�[i�n,�l^�MK����tc%]S��R�jrf�ܨ,����a�r^��KJ�Sn�f�֙DZ��ȆQU)�F��ɗTL�ZkK�*��q桐<U��-�qT?W�Z��Q�i�WT٘����1�ڼ���,��o%)�4�ee=��=8eJ�T-uj�.��d9��ի���h���[���Ó0$��͗z�R���b��#ܩhl
z���t�gf������ѧ0M�Ԑ��wJ��+v���b��^�Q�Х�Nh�!KI^R.^�wM���-�z�b�{���O�uCf��+�f2�2���v�#�{j�a�j�tf��b�w�%*����$N�J[�jUb��nźvn�sj�[C/e�cjmi��Y2�?j��:�A�Wk,���ӊ�j4�����Xk�"P���Y���U&h����b��,���׸���t�Fʘ-T[�D&h�MmbY���J�����&L�%�� D�W�*�4��[�"hR3k.�ࣹ�oN��r���5v���][��7���6f8�Ch�	8�2��2,����J�f��\}6�tE�W�U5��D7FeQ���6��k2�Ix�yf�a(������(�-Kx��-��m[up�b��UX4M�4̗��������T^[�|�am]QYyN�C̀��F�Q�֍kh��mE�l[X���E�F�ت�-��km���+[b�mh�QF�b֨���cmF�-��V�Z��Q�֊�ŵ��llmV5��Z�b�Q��[j6��kX���V�֣mj���Z��FՊ��+Z-E��-j*ڍj�m���5�m�5[kE�V�����j��ح�Ŷ�U��j-�F����5Z�m���Ej�ձZ�k��+[Q�E��ֶ5���TZ������j6��ѭX�b��6�kZ6�FѶ-k֍mQV�O�I ����B	#����?�畯�?2QU��!d7��u�E�&�9̖�*��ޫ3{y�9��/e\���Xj���S���K��Em���{�Sfҡ[}1���
	�ڔ[ݵSosM;�_���WSk4-O�x��\�ݫ������L]���t��a5:,̧��9q��MZu+�Ʋy��&n^��wԼF��*x1�x��S�q�3i�]RV9��gou�B�.*�褍�ɻ}u%v��k�3)=��6��~��Q���ڵ�s��y��m*��B�ԯ����_vN�nT7MY̏r�c�:�L��o����Z�r��hf����G�ۺ�m�u��������L`	���pf�����$Ҩv4���y�����u5����P��]$����4:�NY�e�9۲E�+L���E�mP
��sⱍNU1���M'@�R�`�Hẹ�\k ���t�^p���X���|�ѷ�%�Kfy�4�_�W������̫�䏵U��ڭ��`X�;���Yy��0ӻ�G'G!,�:�ݝSmI�*�����V��u�˨q4�T�����>z�c�IfX�ئ5p���WD�9.����5[iV;7.TBtC�B��B�j,��:����璚�z���̃k�}Օ�Y�n����ѩɚj���D�ӑ�ù��7-֍�3z����,�+;�N�=}sV��'��wY��Ū�y���mѦhv��9��Қt��e����k6���R�[r�^���tJ���ӷA�囐����Cr��Ynb�{���,���C��eoA�iV˽:�y���W��so^1��o�Z;��7���Z��,�c��U��ye���]��)=�2X�N��9aK�r�����9�2Eۦ��h$f�[W3�YfoV����fdU�cj&"
��p����{I��j�ƺ�U7+��w������M����ܼ�D�X5��:��wB��k�o�S�D��Τ�_9���3�,�NU3�ޮ�p��)e>n�pI.�hVsRZ���yǸU�Ω��b��\�_^��n�<����	<���gF'�WYU�Mmf��8,�R9�(Ƴc�D�u}�5���Cm9!ݼ��E�K�ط3�����v�	}fT��\B��ԮՊ
�M]#�2�=��y�����cA�����﷞��(�a�»7r�Y��F�|��0wv��z�}�0�᯹5pǸ���F�et�!+h��ˁ��걵C�V5-����f�7
ܪ�����K�3ۆ�*�qR�{%I�+}���RʆQ�F�y�r�t��A�5wUS-�ܼ�wiV�U���T��z�� vmN���N�oJ�1�n���j����R�m5��p�֔ l���h1�
"�k���8�\,I��N\7t>'��(���}�f��w�vt�W�oeb���ܫ�R��Q��9D���)i��T���q���y��tf^`��]�����_V�VӻOR�T�V���\J�y�k��B�Yc���oqp�aV���f�y�WrU�?C�q�������%`31]'f���s�6��(��Tp$�ۦ!i�X�:NZi}�Ȝ^ޮ�l�K��W��]��lz;�7�&qbw׏3Z��N��mn釞>PZ*�}��$z�g��2�b���Zu=g����Nw���|�H����Ut�An�U��B�%�%ORe�7R�6Ƀ��}���Z�J��r�r�r)[-�M��3U��+�Cv�]g2�'V��J9I޵�`�v�j�����˝��L���t�\�wl*])�s^n֌�bj��\�٫�/k-����tq^S��G8V����V�jJ�ov�p�nB��&�w�˘`�Hˮsu!Sw��[;f�ǵ��rm�uknR<5b�w�.��[�7v3s\�F�ԳH/�����|�mҼ�k�Sz���h�ޜӳx�8��]�n�7��Ori�_M��[�5�6�:��B�w51NXuW�s��f�ҳf�{}55�oJ୦p���U�4����y��,�g ��Q���o���Z�>�f6y�R�n<y�:���ܧ������;�ig�oW�|s&q��tڴA;�০�J� ����I.�4Iڔ��unr��nZ
��1���V�,}���5.����G��K�I)�9K�W;�{���!81R8F�&!����sF�m�R"�eaD�݋�mvޫĈ��64f�*�7mDu����{{��r��I�^T���w�pB��Q�q"{�-�W�U��ݻ�й�Y3/r��%�m��]
��
�F�H�|�ͽ�Բk��;�K�ͥ�,v�ݏj_��#��T������UŬ�ӆ�
�4`���p#��mn��F���f:�2-�1X��5�dn��zc�w��uw�=����wejP��Y҆�&��CvmT��L�%�΂���7��c�iN��X��mйVk�Pӟ6�up�ށiM�7Fi��wz3v���_^^�:!ݽ���ۙ��C�Z��9�{��W�Gz���qXy�"Yj0�S=q>��EkV^u�
�wWw4:��u!��̒l�W{�Sşa�ݿ����n5H��eO�]��óy�:eƙ=A�<�;���RH��.��h`�7WH�j��Y�\�q�rb�u�4�)}2�k�n��Jk_�d�ݵAo}��;\�"�[��}u��f	�Пe��N����Z�t�*|���л�������qkk|��׫�әaiou�7��6��n���=�[Ϊmc7�4m}]z�u���F0ur�_p+Ъ"�u���]ֲ�u�w*m�̛�0��j�UySGn���8���3oEUb[YG;�>/{>8,�$���gX�n%tV"��
.K�uc3+�,�a缆&:��A�c�e�Q��6�^��d�q�S��6fulG8W`�%�MMG&�{Q~u����������|�ES�JY+��]X��m�V�s�Y�et��eڂ6�9�ɞ�xI7wh+����s
`����a���Gk5�%!2�X�KْN뽆�e.��;���J�%���*���TR1��9�U�:�y���c8;7O����OjKg$9M��R�)�M^
I�fE�1�����#��Ά�]���+�X���+�����/�
����(onr��<��gcۍ�c��{v�ܲ�/V뮦fS�Y-���z�r2�d�T���#X5f[�1#3GPٻʎ&5����k��{��9�p⫯r˳_Y�!����˻!�>��Z�关U���t�^h<��]q�s%<��]vnͿ�՚{_T]�of���v﮺%US{N�(��m5w�����6o��;D���9�Ck��As��L!Gk����ǚ6�fQ�ʬݏH{�y��6���mՎ�8�݇+yk��m�s����\����V�/u�Sѱ��u��WH�Q�[Uk7PA�u���Mu��s.��y9ڼ��;L ^֬�\{ 3�I���S�"����Id{���ג}���y��La�;��ˬw�<��ef������=�]��;�D����\ή�Y:�n���4��VU^7�R��Y����[řy���;{o�8@nH�u�'"u��݆*�>`����Nܾ����`��uG6R�hd��Vr�t�K{���4�ڀ�kØ�-�ܜ�����,�zڡ�!X(�⨗��Y���yr��Zn�pSn�5�E[�t�UuN���3�j�Wݡ_���͇��on�b�7yg*�Ue���zM-�3G����Z�J�U��wU��}��.R��ks��o6P�,�W��5��]zM��y��u�����	�G6���7�gm�8T�x$�����]�v:����jg)TC�#����b�5��2ش�i��B�رEJq�l�]���S{�W��4Y�o�#yYc��Wq�D���+E[AVV5�)֖ƣ2�.w��7������o-�����fZ��o32��l`�UH����y���[s���w�Ì����L�A��^h�d������*��+
f��mN;�w�B+�+���#��X���ʳ�ҥ�"�]JuԱuk1���������u���SolBO�C�ڷ�b��O����6z�f��)�B�҅�9�ar�$��7�x�L���p\��j��nbJ���#�s���[��㛂Ь���y���S�R�dX���P����\:�ΐX)AkL]x�!�l�}�w�6�y�G�8pYҲ򌺼}��6�N��V���9˰o]�ib��1f����4ܜ��yѮ��Qd�Y�ކ��;����"V��۔�fnU�������Ӄ3r������h���f��G�F�F����C�ar<�9c�Y�QwB�6�żʕHFv�����H\ى%B����Yú���č<+b�(��PބQ��k��+.��ls��C���a�4(M��}�uue��[��o�퇓v��:��mޢs�����uU�Z��i�dL9H!+��YǴ$Z��i՗[�����UH΢�X9���U��)�Y�#\��0�r�gf��A�Tb��'m��W©+}zhE�w�,=)����ry��H��7o.�P��{����NK/;[�Dm���n�o|է�
#�n㼜eΪ��8Ֆ���n�]��ۀ�:�`� �����	ʖ����u�n�nJt�d�u��q�Cum�W�rʊw`��aՒr�������V����
��{dW�����гE,*��&�}� ��\��*iC���������Yf�f�����l��ꢕ%�Z��k�]��w=o[�5��u'�(�E!{Y�{���z�{�dk>����u6L�u��em�j��r�E4.�n�bV͘�b=9�iTU�����l���.�E���YM�ZM��6�7"�6p�͊�����55��4����V��U�U��rv��UH̻�ՇF|�ZU���u��{-���#2-z/9�,���SX�Pז2wmR��ޫ�{�l��nf��Ux3o_`8
μ��!v�ot�/�W��ly�ٷ�yr��7/^�V�[�)O��yÎ���wyQ.�X�n�/��]�a:����r��m�W�Wy`٬��s(,r��d�mZ� õV:�]���e���^.��:���y}���+Y,���K��]�k7w��e���5�Fd��O���T�\tG��q^�Kܪ����뺹BvBWn��C
q=[u�Ӻ�l���fGw�_Kv�%R�WmIJ���!��*�f$/p����[��悮�f��L��^�;�.��ڻy3�-[�M�[�go�|�fe���L
��yrGW�S���m�vf���y�a�W��v����딹]s�Ev��{6��kP��w�b���Yo1Ota5�r�Lq��o�\�X`���uW��ýT/9]�!H��[a!�ZʜЪEmv�tQ�:Z�2v��rP�v�\2���#痚-XJ�F��X��&�:)L�Z�>�:T�˿�l�b�$��ղ�'I��y����,�7�5K��I�������-���42�*�ݤ�r�Ǻ���K5ǺwL&�յ3�թ�Q'n��V��bn��#cL9R��n��_*����˧J[�޽z�V��������Ub�AO�rU6L�WJu�w(3��)�l�����Q��>�9x��E݃B�7O;m�wR���r�˽n �K��R��A7��B�v��6�.����'n}y���;l�*����יΞZ�٫2���֊YI$�˼��o]���#ug�(3jQ�{�#��=�=�T4�d�8�<����`�X��>�5�Z�·P�#�V��Ջ���0���좮�t�k^'�4��E�i]��wTT��}�E�����GE�׳Mr�A�U�0�I�Ֆ2��^j�ȍ��B��d�b+�Y��f����4�uY"n��iGd�K�z���8i�vQ��]؞��1<˽=���b�2��)�Q�k��� �t2�\�'��1o	}UEf�J�uB8V1w�Zd�J.^A��u8(*:-��)�Y򴵎�M���`�g^10p���.��i��Z�t;��x�^m�1]�����+;w�;�u쮬ʬܽ�u��]�e͹(o����<z
�[�����b�w���:n�)u�J�1�E�u��{r����%���6�ػ��U�b��I�ە{B�Dp�A札��CѴkX�,�ܝ[�tVwF�bޡ��M��u����x:���b�I��\�h�D*�U%�dP�ύ��csn�wJR뛁ic����2��͓ZۤU����֎W�#�2B�F�m+Z�co�e+o�Jg�Y!y�ݤ�]��]KqV�\gv`F�Kcj^��2�z���1w4{����f�Bc!�4��6u�����7��cc2TǛ������!�k�E�s�p�ʼC���,�!�wQ۪�5�]�Bէz�C����Yݖ��eلouTY�{�;�e:xz�M�f��Qm�Lɫ��$�Y�r��wwg�E}J�&Qw�GS�}�4+��f����r�EN��EUN=���������j�M�fK�o5@n��-�w��r
�����[�QMa�TE)���u�u���ۭ�8t���l㛌��p#��M�-��j��W;�&�2�+&�xS��
7]���m�GV���x�%W���VFe��6��Wb�媚/�����;,,�חj��T�����6͛��*��2=�m�IP�#oyU�#Q�U���zt�y�tʡ���Xh<�Y�6���١+�a�ɽ3�U.��V��5vi�OC��;�\��s�c�:�
w�����S{\�ѩUf�we�0�-�Ψ�F��bvɧEL�Cb�3zE���w�7l��mq��Bj����~�`���h^����C���A�ڧ�QC*��k.u��6���Oq����s,�0KS��'jw,��U[D��k�	�J:�%�p�,�����jb��x�ڻZv��FL�	�v����K�T���.9c{gm���Wy�bq�l;��u����y�ږ���.��5Zc��c=��2���^LG8��䫷�x6wi[vɛq̮��.ZF���j"�g1�U�6��f��u�����BI@ V�c���:2�;�n.�ee�\�FSܸ�(B��i�Rd����m�2��^�/s^bػ�.�h.��*��Kc����Z�����Z;c���s�rk� 8�7�c<u�>&*=��^^;<6�u5�+�]��|�8���/\tt���=�=�M�LU��"��]��l��5�EƊ+j擉��7@���uv�n���8�ءL(%Ug��!�Z�}�d|�::�����pW�Y�c]<�[E����,&���k�Ywhb�O.�wd꺟p����v�N�s��o$uɵ\v+���,k�CG7cRj)�i��b�v!M���ƪK.����p�Ƹ��ר���8M�/h9�6�m֢7db���Í�"�LEm�`�2�m�fUH���oyPvb̛��촗0�KO�w�L���!�+vٙ�i�{\"[�'�mm�R�K��>9��c��Y�����l\[�yq����e��3�K����Ӂ��q��kA�ɷo�a3�cG�te"��&��]	Dѣ�5a���,c���ၽvx!��n��w	�N��y�waEu�89����Ж�5�J�����A�!�����x�F�),�u��[��=���ąn�n��q�.M�tT�Į��V��4�Lq+`��c��㫹�/m�"u��JR�������hn��v�0g�A��\\�r]����te��K�k(s۔.q��.�tAQu�j7�L�[�����ݎ
q�:z���6:ݎ5]�7-z.�v�nب�>�ݶ�Pno:��<�-v���ۅ��tN�	�ݶif`M�K�V�-P]6l��s��@�Mˎ�ш��Gy�˺;A�w��z:a���gf�5ckn���LqɷU:Z8�r��/�zүI�Q9�<�;O�<f��V�n7n�Wq���V�ŭd�J���'����Q���A�Tl�[���d5�f��C��Ee�e���f:�v�'<K�÷��������N|H�q"�۰���kȇ�H7V�BK���j��c���%����e�!��l�-e��n���j�q7cK�S;��9�h�q��6aGil�i`��j)@q��'�$�k6�F40M�n1bA��ק����ocG�)�//o�|왇�RG8��L5��e��.{%�S�kgfNλvO\X��y��\Ѕ��*6��@E�����K�Q�^!Gn�S��n���k�3
{:��d�v���qa�=&��K��mX�˦!���8eH�9�=��)e��k0�LáX�rs�g>�۞��N���n2��Ū@6cl�O<�Y~HU�K�TǶ��y8��)݋��������nЕ۴�Ӑ� e�v��K�Pњ�K[�֖�R�4��uv3ڜ%K��GI��Ȼ�皖��K������Onڹu�xM���)�꒻�^�.Iytv*M0Y���X�eca�k. �$#CRnطl��ҍN���L��pfP.�r��b�Bf[(n��C3m.�L��Ȱ\�;��Ιu��uպ�9LM9�'$��D�=��x�s�`�#��]�����(�MX�*v�5�`�!.�N�:�;\5�U�Л�m� ޡj���hR�����nSaZ�9����L\��:1��\�Zl����j�(lj-�l-��B�1Yt%�3����5�IJ6�Ӈ�䷋FV���oux��0��^�a��v�g3@qe�/mv���vq��I�+Wfi\��-�(�ƫ�� ��v8�����1r��;X�vy��z����V|�t��q�In.�N�U�)�EƸ��y��tp0 ;6����,Mo�V4��e�Д ��ظ����L��{>��(�A�9�[+h�	hZFč�3B�	��,[���Qt�j�x�r�:2q�"��n)�Z��%�)ӊ���k!��5Ѣ�F��ہiK�OK�khJ�b�-���9hn:�ѽpٶ�ݞ�6-r]"1a3(1�iXihr�ϔW�������o��Y1\uWjCd��k������v]��]�6-˚���(\Y�<4��O!���ܰ��.7m�|�ȯNyN�`x۬F�����C�F�c=k4Ŋ.��m%�,���8 �#�v����J�iQH�KC6
1Ų뛋�6�5k���y���ʮ�����G�-&�8���\�\��rn���`�H��՚�:� �R��^�+K�Zf���.ll"�ǩ�ď6l�N}k�gF��+v$�g���0��l�VYB�=y�������n{�	�{\�.�зD�� �h�p�op�;��pv.p��i��ܳ�:��U�v�ݍ�rWZgu��k����q���΄�F����u���a(�Mp�
�t�ZZ˩|e&�T�z�A�k�؍�2k3�l�m5�q+̈́cl��;M��]ugpUc�\��;Tv�.7Wy�i8���]sv^W\t4e1��Y�^�n��`�����\����M/����0�;X�<�:Muzz�@N��V��[�ù�h�z���C�nѻĵ�]�t�k����qu`D�y(����{nIt��CaЂ
1�h�](�|�lkg�Zd^�� �9҆�f��e&�k���,��>ة(�71k:�m�v�ړ]Jf޷�3���L�1L�p�V���Ү��4��:gg0#������Mb"����4G,ƸH�JX MpL��fR�`���1�ʗ:훎���X�^����L�G=��:�������] �`�y�Y�We��64���+6��%Љ��V�j�Vc8�a��P�����󎪐��<��Ղ��BkI����x�)eB2�P4MB%%Ktȼ�']`Χ�­�.��Z�Ӹ�\=i�a�⣇2\���(�iB����U�Mu�Z�2�e
7B5�c�h
u��Q*n��;۠��[���+�qӹ�[�����s����ͱù���1Է��--���v�֐�KSsl"�ˀ�f��2���2��.q�R2�)`�=A���&��k���&.t��&ۮ����5�_ ��U�����F�q�=�Fa7*'6.�G������Ӛ��Dy��Iy���N�ע-��϶��a�<�.9's�%[`쁺x�ez:��X!Z�XB�&͍hv9	��3�H�i��4����������8��G.�I�h�*X�����hڼ��6J2�k�fԴ��@�k)KKm�k41bV��x1X��H5�ƭt�Iqq��]���sc"��`�M]u]�y�$���3��8h�z�6��s:�0v5vӔ&Mk.����J����{�ӷ��Ŵԃ����D��[ڶ;1�&�W=b��:�X�����h[�r�b׽ gtd�a��=�����c@w/����n�(,m�i�k[�ܶ^�C&u
�m�XX�e*a5�9������NȺu���V�������s��T��mef�Q EZ�)��Ʉ[�����!J��f+7z'�YIo�񅮔 �R��m��9�]�]ʘm`gv�������r���g��iv��[�d'�kud"ƚ���#�of�܉O6��ka�`=]v�B�2C��g��G
����h�dG2��7n��7'A���-6&|]f
�6�x��=���X�:�^ay�S<m֡.:�n+t��3�Xwi��
�����){v��\lj�����)�1(�P��i-b٫�<:�F�$�v\[����3f��4j�2:\Ҍ��6��o-��6&nqБ�6Q�e\Fn&0L�ł)�f���9lDa�5��:�a�
��0�ˑ���N/&ݻ���V�U������@m�;Q����p1��X+��q���*s`�K���e[���˲��I�Gy�yY�9��[��]��ML�
�9�VRu�.,�$��&�a�l�9�eb���gb	��Rl��9�l�&�6��v�F.�m�󬥆�Pu���j޻	�$
<�i��(��n��m��s�r�%F66���4s�V��pe��e��.N^��7:$��v�b8�k�̆��9���;tC�ئ��4�׮Һ$��R&I����Wc1e��.�vs�`lf� ���p�hK�Q.i������/[ȗY\(�i4jA����`T�<l���ݡ�y��� pH�:�'Z�:�bw������F�a8�Pv��$�'��k�##ġ��SX���C6
-�ԣ�2�&��<�8�AJ C.��m�����-ke5�J�e�]�-Ֆ�[n�Mx�W�KL�i���f!�y����f��\�z�U���f@�4	��RapSE�C�Y�Elt�uњ��W-��k�۞i녤���[��������D�z����7o!f1]��&k�fsʘ�Xcgb�SD�G�$�$��e;>��ۍ�B��[p��6�9�7Fz�7�ͭl���^�1v�#���`���ïmy���+In�M��G=�<��m��ˋ�|&ֵf�X�=Essj�u�Έ;s6D��@������!�\TZ[�ۍ�`��Ex�-)��h3J��k� 0q��0��"��<���o�<lBl�X]Y�X�ɶ��s��M����v(O3ЌpV{��Ꮭ����<m�ilᲡ�*��`���N��\��sa��R�K��(�I��4r&�����#U�:w�����I�{]�l�m��Ϟθk������n��y���a#�l-6�uqd-� jέ��pNz��o<��)Y�ٮ��;�"�U�3j���Rn6ɍ,��Ƴ��ۣ�nރ�pc4N�=�8��W[>�'u���hK�q�X���&nmL��i���G��0�u�n�v��㧳l[ѷROl@�7GK��i�mWn�[me��L�	��=v�\VMڻ@�if�CtM�We���)��Lp�TK�f{�G����_f(�Q�~�nh���5&9sj0W6�nWD�Ѩ��F�U���"�j��F�`�E�LPE�P�;�$J0Q��8���&�Zt��z�r�h1�w![��ەû�Ri((�ԕr鹳��Q�*4 h�F64��Ou�`�ѧ�Q�ۢg���"��刍%'7v�+��*(�Δ�wW]�w\�¢�v��b�!6�E^W"�/s������^��"4Y6���I^zM��d�XM2���z�p:����KK�n9�a&.՘�.bSd�D��J��.
�j尤�-&OGnNwhx����e=�������4F�{i�ۦ��UUt
t� &"ݞЌ�1oq]�KMV43ݵ�Jl�b�&�l�Ѵ���S��$q�j������	�plT�j10�1S9�lvX%��(n�W��:S<�F�-�됫̘! p�<gRp9rlq�tv��y۵�`,�kqm��k���ʷ@��n2n�����<�Ǎ�$� v茊-��N'f7���Fg�i��Nwg�n�Mu�=[qlգ{q�Ja*���z2iNGO��A��݀���p��]���n���=��58���/���Ɨ<m�\D�n�j��)x4	B�ift1e�R�YK�>�rz�Zx�.J�,�9渗V��.KI���Phq�{Y���	;��:�c�v�'&��<=�8݂�]>�
�,����H��!3Q.x��[م.]M���@e.f�t�>܌Z8:Ѕ�Wo> �����۠���<qx���y5 =�\7�g�}Aֵ�qv��j�OltnHN�I��>��{�7Ig��^ � 4uUEm�VF$K����nha�o𧜝qx�zk��ٍ4��]�7uNh5$�nH
�K��ťřL�m��{����>p�MHl�z%�1vm`6�Da�4s�4�.LU�Rk)ZB5��n$T��KKE�Q���1YF�&��j9�w\JPj���Nwv���Wm�GpQs"�0��--8P��헧����X��wCm�\��f�oa:�8���{�M��o@i������qz!�Æ,�h�tm�6���<�ˎњ R�u�O
l�K5�sش�������%"q�ݯ,�R=��ۆ���4�Ж�til%u#׉�mכ�<n��4v�<���:� ]a穰�����i�J:��I$��@�ٚ4�8e������h�^�*�a
YJ���Dmm������'+�T HA�,HqIE(Kb"�Q��JYkaG�QU�QE��JX�-�sV���a,)�Rն5��A�Yg
R��"�[,���
VQ��[�Q�k(���YK)K}��C�=��������T�Cڦ��r��!aI�+��z�kIUZ7�g���E��X��f�e��u�o�9f��ܼYgm�� �"�B�n��,��!����}y��Ӿ�A��OOJ��ݼ�f��9_oP�7� �*�u��=���n <^P'}_7C���:��Z��y��Ϯa�w�1u��u�A<t����� �Ye Ciڽ�1{�Bo�o�3F� A�A
�~Q�ݨg�gc̱G4@ ���V���������_��Ae��h [���,���4�ߌ<P�cq��Ϟ�TK��@�.��8~����{�5ƒ%mU}E
�Mڪ"��M���'<�b�ˮN҉��&����@�WKs�k�P?�v �!����
����~���"�4�׾#	�;��TQ`Gjԁ����@��#�������vߌ�S�E��Ă����N;�˖ls8d;�F��ԕU%ǟ��~�$�T*���_}�S:��J?^����k���o��p�,��L�����C/V���i_�g�"ߩ A<|W��E�DYd���+�v������&^)۷���w=,]v�G+�r�#9�-8�ϨC�%�h��_f�2|+��
�=���n��vT�)f׾?qҾ#Od�r�5;�_==�@�|Y@��@���|韛�?w��M�ւW�T�o��oq�L��JD�A�U�m�@�eY�������ҝu{U�񺐴�^��:����Y�m��4��j,�`���>t�������h#w��Y���������e�G�4 f��%�r���{�r�o��B�:@���T��H(���;
�S0�u���-_�gt������'�Rͯ<t��־n��g��8�^��a_q/��� �鐁n� ��jmW[~n�B�YCǅU`��.n�]���[N3�{S��Cf��snr�:�m�ug�7�՗Jn�giڡv�̬ROfǕ���su�GՍ���6�C���%"�!���A�}g�C�Ү ��,��� �.RYew{��^]��S,z>w�e�Dx�
�sP�Q�̤A��Y���A��e�z�*��ޣ'��1�9+���.���k�:QZ�	e���Y��m;�Ș&;b���jQԆ.$��=�P[=��N�k����(��fWK��.#�İyʱ�Ck�؝�׺�n��f{���2�u��_nj��W���@�K�,���m��9U60�"6Y@c��})��{w�+�u�<?J�"�J�w�=6�Y����"��u"���_�����ٍp��n֧�or�l�ʷ���0���Z�_/�,�Ct"��J�I�|f�����Bh-P[3�m{Պ��a%"�4g�۫�[)���+[�9�]��W
髹�N�u�M��e���w:������S���j|�d�n�>���vp���6��[w>�!�B�n���Y_Ch!���!��;ꄘe(	�b�gҟ�����jw�,`��L�Kr����9nЧ�P�]݊$"Eo8��)�Gf����x�a��D�J���y�5a�OW�N~��z �!�~n�}�9�~����{#�8�k��^U����> ��n��	e���%��]����^׻���6�^�޳l����ؕ��_d��� E���պ����͏�ƎAm|�aYr��J߯��l]@���s���������PD�Bn� ��_�B�+��3�6��T ���1W���g�W�~��#�:�hp�������u"<Y_�@�[��B-�y%����}1���}�k�����`F{�㒑( C-W��u��U~"�=�W����=>4��QK���	q��ù+��F�+���d6zmf�}�.�d�;�_�2׵粳����3����_���e+Fń�ݥD+�P��umn��`p�:s��&�h�7c��q��A�\�C�iN��8�k�\�Cpq�����2;*s�}(Ok�n�`��u�9ڛ�Mk��0bj�H�2��]���Y�����ˮN���RE�q�=�8x�:��v�/��+����&ku�y�l��m�z������t���P�x���wc�]B�C߯����4��Lj��q����d3�������4�ԅ�o[��X~,��[�%�W���~�ʾ��yw�k�~_��xg���T^!J@����	n��j��O�s����kA|Mk�5����ܟ)�߈%�?*�-�Kr��مg�h�}?���?7Y���vﱟr7�̽��{���p���9+��e�����D^Fa���t�����H�Ye	������̻�_s��A�a���q>:��y�b3ݰ���B<�X�9���Z;�o��N\��Ҟ��\��8�k���O�k_7_ae���V�&T�=k3��n d��D�f���u=��c%���Ƹ8���ZZ�C�Z�9b�tz��<�K�嗰]��y�>��z-����>��ڕd��Y��@�H�,�D~>��q^�	�ѽ�C��T�s���l��IQ�.�f��?m�\ɏ-Z5d��z�s'Y'.�-�OI�uZ��	�H�����:Vk�y��<�kҘ��� AΠ� �*��B���iE�I��n�4����!����͡4z��v�rN����q^ׁ�Ҁ ��-�Ȳ����C"��n��̪�+��Մ�������x�їa��x�^��xA��,�����n���,��h"�ub��54�`�EwC��f\�7��7�x��@�:���@�i���4�m�
MPUD�Jҡd5��Է=`'��N1u��[�t�p�Lv6.�~���w�΂��Z��m������عH�-��+ξ�G_��� vW���(���@{�'����YK��f�/�;�3��^��}が�`�=@�f�;���{U�Z�Z������j�x�_��g�fq������.E�!Yҳڳ�(��ְ�~*������ꔺ�l�m�[�^>;˯�\c���5�)<w=�yչo;�`�C���D+�@�H���@PM�e@�䄭D_����}w7�.����ڤ}��xO+��1Tj�#�|�h:�~:|Q�E�Ι�o�_]p���ϭ4=������8��3�	�K�A�����-���e�ק�T���e",+�+��՛(Q<��9շŧ��N�1�QՒ�ڔ�Mh��u�z�^��ҁ|��"�͕���cv�K5�X�N��~�qYt��"���	�??V�C-P �_z�|m������|E�����K�y��f[��^�����E�^���9��F G���P�A��!��f��a�fg��.���Q�����4�
�m"���Z����t��~�^])��=�f�>�;�_��_c�6'wŧ��KS��P�2K���̬�H<�Z2���s]+�R�;4[���;&Wr�z��ol˭�8M��%U1W�A�>�ԉ���^m��j�׼���~r�D�C-
�H������jίe�ݖ�݇z���l��{N-����J ����#�,���>}n�ߡ����/�%I.����[�l��)��́L��!4�qR�����O�o�ߞ'��"B-���C��?h�b�|j� �=����{�U����!_����f��[4p��{���1��l��4ܝ��{e�A�h.�"G��Y�ˊ ��������c��me�_���E���y3�9��9��{N-���������H�,�H!6
�.�R���.�)|Am��1�f�c���i�	�H�A^�UH�4�G���|�a�+�͠�n��8���h����]�,4�{�Y�!ބ�� �2����������~ͣTA�'��-+�7m�5R���$D��Ң�ۨ{7���h���]�vF��[\9�ۆ3�:��=o_=����/ϳEu�`��L�uVWt�wM�pwN��5
�ܵ#=�c	]��͵�<�q.T��C�[bs:�;^�[��	ũ��xc۲:�1�N��tvb�pÊz���up���`:f��E�&�n-tm�m�q3��Ʈ�wC��яf�"�-Ȋ'd:�m�C�δ-�[d�)9�#e��6ԂhH$&�hJ��"���������5���2�%��gWq�B��b�^|�#V�L�y㼙���}���-����A�B�!���������K}��mx�y�f���m�s�J6 v/�V|A�W�6��@e�9u�90�w)|A�����W�R6o�$`�� ��Ds�m�Au�<��ܢ��}�����u��,㪤#�޿��JY�UT9� Om �q�H�C,�ܫ�8�Ū`�ڂC���C;�gy�?d���qn��>:P"�s���ؗ{�0�G�0�Ctn�韛��b��� �2.�A���{�X�L�}���f��q�E9��fv�i@R"H�b�E���D�μ9�U�@���=�vS�n38�����e|A�A|[��,���x�=|q�֢ ;�"u��`�;@�����͠y@�[��~T&����vk}yd�E��FL�z]����Uf���wu�J���A�ͪ�#������,ͣ��ɗ,����*�/h��c��/����2w��O7��k�;+��?-h/�uf���%���(�;k��C,�t�-�{���Z�^h��*j��;����U�4�<vR���m|�}�V,C��p逍�)|~�eޕz_��������P'� �:�e�A�$�DA,�ۥ�#]e�N{⧺�o�|�D~`�{�?zo_ga��^ �(�5��t��9<��x��r�����V����V gXCg��h�v���n� `��Rl[�����P����}A8��t�!�G�{ޞuq`�=�f3�<y3]�n�]Y�#~���g9eǜ�G��y�ߵM���7���6�E�ǚ���.�B? A� ��!��Db�#i�TyP%�"mC-_�}�:��<�>=�;{��F�A^�E��e�gc�嫞ۖ�]19���e_V��csPU�tov�X:1M�\�c�uⳡ�6�۪�LY�2�J��W^URVn��{��ʦ.��ռ�5S���Uȩ��j^d�����)��Bk�5�Z����Q���wF�U�u�놵�H���U+%���Eй;��,�Ol�cJ˸�!�W���T�Vꘔw��y���y���j�[�;&�o���U1A�IA���ý�S��ݳg-��̺��a/���\�k_.�e*���p��V�
�d�]F�I6t.?#�j�
c^<<9��ฤt{��յJ�ͬ���T��*�O.��{tv�m��I�,�4`Ν(7�b4½"�N��5�;����j�=6�ze1o��&��d{|\�	edW�J[�{s{�ʛy�h_�E�sIok:+ �결�A�&�]�P�u0"�y�C�f�m��F���ӵ��K+5�}ۋ2CƺV��pG�ݢz��S�;)K�.ڒ���[�_P5Pn�[Tf]e;!m�m��mQoa�x!�U����P6��{�{��e�y�\�R�Q�Q�!Ẕ]��7�V���v�:�n�Euyt����Gw:Κ�\�9ׄgLVu��ח�OK�]�3R�=[ڷp�� �K���q���.������n�kY���ZB4e����\��-�1��X�J��hu�O�xs�Ȫs�h���:�bK��Pg
�@˝UO��=�*�s:��+�B]��=OggZ)nW$3彋34ud7{ӟ���OM:��.%% �EH��c��l�b�8�i���<�7-r�r�bMAt�I5;�9c���3�IΛ����o{qW��]�ʺ�����t ûs./wLG�ۥr�����u�0���ӥ��b�\wnm�˕ӗ1�;�J1\�o5׻��\ې��s�zF<*9q��u��ۋ�����!�;��s���G�j�ǆ6�.r(�]�snF����L�ܹw'd����^ys��s;�T�ܯN봽ۯv���9�����܈������+y�nt��׹�/u͹�i��=�s���sr��N��Ou���QI�u�p�.�(�njw\�r"�Ξ���*��-2*�RJW��C�Ώw�s�=��u������i�����I�2S�r�R�) ���p�Aa���E��!I��NV\
@Д�XfPh$����\� ��ZA�D) �_5�
j S��l��I
�fQ���Sٜ�}��ޫ/���֟�Ԃ�a�ai%D)�;P�MFRA@��}��ʯ��=8�X�H/kwAtAH5*}P�At0)2�MD
H)�ˁHhII�C2ᤂ�L)�E��2��~{[���pG���%C_ ���yl�-��?����I!AT�E���_W�$؁L3*�2RAB�3(�Aa�����}�~�ߎSk�݈@X�^q3���5���0�+��8����>�ڬ��Ѧ�����AuZ��R�l�I��4�Xi �Yp4]Rʅ�~����7�{7�??߀� ��Dp #�O���N}�<o�[�v�R�) ��T- ��
@�h�����C)�ˁH�I�e�$���E���]�ُ������U�) �ꅳ�%$(C�F����߾�o.�o���k�bAy۰�aI%SeB�42�
L��H,4�\˸�g7�׍w�zAH?��$���Qi�
H,����� �̸i ��3(���R��� ��;[]�f���R`�8:<G���h>��
B���(����RAh���
AM�2�l�d���D3(�Aa��$2�4
O}�y���0:�YP�OFRA@��I����������h�fT4�&k�w�Χ._���I ]@Dp 
H)��p��X$&��ߵo�Ğ5�����4o���h�|�9oAjH�� ���&a�&}�Y��إ�4�ʌ�<��7�{��g�ix�Ry��~��_���l�k0ߊs���9��R
A@�(���) ��T@�JH,3(4�
B���- ���TH)�eBؐ���s����~�95R�;��{�?q�Z��MxyA�o� ,;�\Bs����
ܧ�D�knU	FIQ!��$&aS���uͽD�ڧ���aNݦm	�2�Y�����i��(d�����Y높)2�I�) �Te<ʀ����t�L��M#�O����AHU�{��^�9����ZA��RAk;p4�SB0�T-����P�3(�Aa��$2�ZAI�)�eB�
A@ᚯ��g�c�g��M$���D�R��jH.��~��W}Չ���	 ��|)���P-$��³.H)2�I^����W�s�{����S������~�Ӥ����v�H:��\ʁi4�L3*�̔�P��eH,9���WZ�tw����_s;�s�������Ă�*��Sʅ����v�$���P5� ��H)2�H)��~{�U7����P- ��ˆ�)�E��B�%�s#� O��j7ݱR&tty���|	�{A󤂐���H:(�$�f�9��i:�L=ꅳ@�I
�h�Aa��$�A�H)(B�fT- �fY���Rs#�.7O����n�?B�]w�#�O�6>��>��|����ۗ��@�- �|2S�*��%$̸i ��3(�����C(�G�" �Z���?2��/a�+��Nƥ��U.ыnj���4L�٣���\-��׽O��v�81��V���d�Ϟ�݁�N�.1�����K�Ɨ���\*���bFQJ�V;��pX M���t�65�<�۱��K]n��v'\�X�hͩ:�!<st��q!$��!2=Wkv���B5v�Bj����y�҃<��1����qfeǇKcsź5��6ᵽL�3x#��^x���-��٧=hg:�(d��d<�N�e�Se��ȗ=Yʥ��{Zz|�H�v}�R�p�n~�����F��mB��Al7d �h!��mm�Yv�س�kF��)��6�XsUH)�U��iR�RAje�RAMD
a�P�i��
�eH,5��^�ﾬ�����_�Ă�a���
J������e?��z�['�RA@�9f�M$�ہ�肐jT3*H)2�M�RAe��e����X~�t��s߻����aH�-&����C)�z�R��}���ޭ�x��vߏ��{A󤂐�TyE�J!I�_��
i�fT-��UP�u���A@����ñ�$���RAI�B�g�H)RfY�����Ar��RAH'�%|w��s��C�Zc��<&�������� RAe%?W.!���eB�0��-&����C)�ˁH�ʅ������e���ٮ~��=�- �RAh��RAM Sv�l�%$�$��?	y�W����|���+�H.��
O�)�2�l�e$���g��[hϹө���AWn�� ��j�]
@̢�B$P�NV\
CI) �̨ZAa���E�u������7�����Ad����p)S{�ו�z�����ݷ�i�{A�� �*��H:�B�^�j$�0̨[4�I
3(�Aa��_U'��������\������0��v�]��+��b�݃�8��9��t�˹oд���aᅤ��}�ZAH(���H) �Yp7.�)�eB����>��s��Ͼ2�����6����
Af{)���|v����8��\
H)��ˆ�
A@��-&Ф��L�+. i) �̨ZAH(�ZAܢ�]W3���׸��G��ݝy��E��x#��awsr�P��VK��SQ��2p��~��>��×�3�l�p%\^R\�j��@��޿�) ��@��f�JH(#��$|	�H������z�G��|�|0�]�l>ai%!L7�d��H(=�4�XH.V\��.���AH?��v����P;�Zm�*2S�ˁHj$���2�i �fQi6�$��e����\��W�R��ȿ'����D|	�7 |�
B���H:��Z���$��2�l��I
3(�Aa����H)>����������a��H)a�Y�����Ar�p5.�)�eB��O��{{��2�L��Q e�Dw�Ae2S�r�RRA`㿽��yݘ���1 ��E��!I��NWn h�I�2�N�
B��̢�
AH.���
H)��fT-��޽���~��'R
C?Q������qw:��z�� ��aj�H)>)�n�l�I���I�����e��� �P̨i>�v�����*mh��(�P`�7nn��\��:���=x&�5>;A��ou��w�7E�� RAe2S�wCI) ��j�R
e�R&�Nb_ H@�팎}��F�������|� �+{�+<�~�@���H) ���Z���@��B٨�I
C2�$aI̻0���XfT- �׮��|��i �7w�Q �C�H.��������p8� �|\G�%;����RAaFe�I �fQi=����=���_����S߮�(�ݨZAH(�- �RAh�֠) �̨ZAH(lC2�$����_��Ο���v����j��::���prI�^�L̊�"4���TjP��I�D�oeL�8���C�6��TR��A��{���>���o����P�[D��|/yv��$��0��-�L���S��I�����]��TAH5*�$C�3(��@���_r����ݓ��	) ��rᤂ�C
@��ZM!I ��p��J��dm�K��G���8�">����H:��]}��Y��^_�}n����0�T-�) �B�4�Xi�$�v�
H)*!L3*ɡ��P(3,�A`j4�\˸���?a�W��3�AH9*��>���9���U�p8� �|]�R>d��]�P�II�eB�0��-&�) �P�s-| �����5;<*$8qQi(BT�/T&%�[!M]Tģ�}��	1wX�>�V�i�uxR�I �s�ZAH)��֠)4 Sʅ�L��P��4�Xjw5�k;�~����H��bAw۸
AI��6j�su�ka�T-��RA@���$��_e��Q �T3*H.���E��) ��Js.�) ��?s�u����ۿ��}H,<;�-&�) O�G��9�| 	}ۋ�΋�K���Xgh>��
B��;�- �B����R
i�fT-���*��>���?$6D?v�$��_z�6
Aa�T- ��i ���]�R
A�P̨i ���!�{��7�l�w���� ����
H,����wH)Fe̕��d��!���^�@��1���$_ })[A})�Zr�ײ��'��^ ���3��ΰ�v0G����{ͻ7Z�|���Q55n'���k����Pu���TFڱ�`���qW�_�؉9������b��}?��>��v���������v��������#�|+�n��1j��osK/�k�����n�M��c���J6Q
s�-݄w٧
�W���=��v��b�\l]
�6�R�A�쯐�����h_p���kr���o7k�o�0(Z���B1�G]"ź�[�� ��3Ʊ*��c� �(�p4���f��}I.��x��yH�("��v��N�~. ��e ��@���-�sό����{C�ɏM�:Y}�Z�@�6�>�����n��VmgJ��ξs+�t ":6���S���p�	Ry�^ �s��V�B�9�z�ŃΗ�{� Cit�uc�L���Щ ��RCt�'~���{Gex�R"J���ֆ@��5��zfƉ�B��aÛ����w�Z�w��n�Sn���9;|��U��:QڛU|��o�i�fok?3J����ͷG}���2O��Ok��{��g)�X'�hA飂)��e�0�c��:�Sy�#���n���u��M���y�$��L*��`���9�MO5íGܷ=�D�uЙ��3ӹܷ%�,�w
�3W���AY�I�B�cr颅�9ͻA�ĝ�L�=`�,Mq�9٦��۱�M�]���F�'�P�	]�ͧ���cF�\F�5Nmni�j����~�#��+��6y=pУ{e���u�-۶�'�4��B		5�� V�F�>@��O^�W�v��
��E�A�m���T�B���_ A|Ct�%�@��^�m�]�lap�N�w��tgFF0o7k�~;�k_7Hw��������A[@7XA��<�5��r{���;t���{Ge{��� A�D���@�H�*���ܐ�.�A����i*ѻS����^��~��#���n>/���Rhh Cu���|���f�>z���x�w�w�^��v��tt3�� �r������c?G[fT��e5(�rv�����'Z��0�3��t�L�M�b�z���w�d�g�g=}�"�h!�W��c�����It�~"��^�4˚��P���"!�Dw
��W��O|Z����*<�.�˼;'"�����S�
��R��5�m,�9���:{t�,=�T�se�e��f���W�/W��4� ��?����I$�����O}V{��.�g��~�Y�vÞ� �("�g_��.����_��|����@��_�C�:�2j�{}�x��#�5xJ�����:�6�n��Ct�!�V��2��{������ 㠋��6���*�Nܥ��s��� L�������܏~	���ź@�Ct�!��wu�a��S�A�7�g���3�ב�ö��^W��t����|�[�0п�7�P�8��������[Gn��su�;��T�$�6���׿{���C%���7��9�~�B�WL�g��F
���c!ç����"D������ An��r��!_��������w���)��Ur^p^�^Oh㞠A�HD� C.�0 �9��G��|�|A�(���H�n�3|��ݮ�ej��P�Uo,𥉉�YL!h�C0Ž����Wv�f��J�\��3{�,J�C��t.�^�^�%f��>wx��>���vg�'^��p9��/(�r���_ A�h!�7���fWב|ϗŴ���s�j���n�^������у70��+Q@�_wW|A!� Ctn��[��D�n��P�!�;*��g���y���3+�� ~m/�m5~��}�~���\3ٙ{��S���)�7mk���8��c[�,��Kd�7�u����z��-�����t��Y���=�[�� �z�p\�{���C�N�}�X?6�?;K�@��y�7+v�0~�A|~�A	��������V=���Wɵ�uA�M�5��w�,c��h�9E�9V"o�/Z�Jk�Ǿ�Uy38vb<,�v�fR Ⱦ�_7A� A��O2a0fT �_k��N���3ށ?�u�����9e|s���ʭ���{�/�n��^h4�[��ۺ�۠�Hi�����Դx�۰�M5&
v]�U�+ͣ�JW'k�����r�Ǫ���&�>Wh#���C�����X��u[�њ|+t�+�7Ԉ?6�n����UZ��V<L�RUOOC�t���[�\�֫����$�/f�ǡ�U�B����~��器�,����U)38{+�������o����>h ��|Ch u�!�ʗ=i���9���y�;'^���aѩ�<��( [��{���Y��-��vW�6�?6�Ŵޫ�2���b�łߟ����Vd���R���"�7_7�i����Q�0�����v��QS��4�K��o�fPyomW�шz����/�� [�A7H���f�<WЊ�_[�(��Ʒ��i�x N�~r���H���J�`��=�Z��Yڪ�>���V��ڼ�s�㹪�Mt0�����vpY��*���R��1-�j�7}x��&����N8*�v�I�-wr�咮��z
c����	����8���D�یn�s�ݸ�(s2�k���X�WzT���;8�Smb=9����M7���U���;܆��j��F�ڸ��f�5"�����|Q�L۝�֮ٻ�?w1I�f'cyɽ\�Ց�Ɗyy����YC�Y��2�#����W��D��NDaܹ��G-����2�=\=$�^h̵�7�ROM�R�|��48�9}�ܨ�]d���ԗ�DVq�(�����iM.�x&�k<$�_����T��~����^V��in���W�)6Q�4�7���o�1�,YN�2�]!���׋r̬7��>������Ѫ��$���Z�Y��h��	.K�b�1|��y��+���/�!�-�[YG���}*�{79uV���зUÅ�wG�-S��vK=��� ������F�闗שY��޸(�f�NF
��Ya{��Wl���o��ҡ�V�v�':Q"^�	�����7�l;ػ��a��s��R��_EGq^�v���t��[[�8ʾܓE���_��D(��]�����3S��(���o�5���Z$���#�㲣w����(��ӫ��MQ���[�֮�엝ѓ4$~''=�+M8�d����V�Ž�p��J��i��\졨�u�N����M���Fs���s�u,�9��Y�X�m����c:�d����Q}CO5t�S7wݷwi�u���9�>0gE����R�iӼ�����:M ,j���R��H�]�c\�E��ngs���S��sr�h��KB\������5��w.����99�۪�9�]��h�� �+��	1�4fwwwQL뻕���wun�͒0Xs���+��(5ˋ�r�θ�3L�ʺr�v���4:���ˁ����rH�nnE˛���˚��쓜f��;�J�dш�'t+��J-uf��s�s\����1��r#����#��c��\���ܳ� !u�H��&B�!E���۹s E��wN�����fu۔��Ȉ��pۤ%��L������ZH�RƎE����\u���^��>��a��ٸ"�^�R� -��^v��M^݋��ga��;e4�zz�c��]���ʤ��r����Ͱ&�@�.�ᬰ2�<��Y��G��C�]\z��E֫4s��H�b_'`�.Y5��Ѯvmn9ڮQ
�Vͩ�%�s
`j�8�̘�7b �-���d�]��i2X�*rk��BE�@�C���]vob��a�u)-��:3�cUI�N3n�Y6�$/@�ƺ[�au�g	��4q�6YWa�m�k��Ԅ�Y�� ���u���Q���ւ�j��6{)1�ff(^vì����i{f�ha�V����J¥FXMt6if��x��f\�(���] K��,㝭���ţ����XC2�;u��.}WeG�s�J#�i���xV�Iϋ�˶1�
&8���'v��l��;D&�N���]h�,,@s�.&4-�su�f�q�hCJM^�@<<g�+b�K� gx��g�e�>V�4
���[.�[�l�k��۝�b8��g2��yx5� �α�7�uy\��v����]���Z]��wY�qԔ��ppCv
����Ž&5���
1-�����XU����1V�����:l���=3'`:��\s�qɹ�#��h{i2q���7DyM)X|��8r��q�lt��N�v'�Of6�α˵� %e�Y��6�,��$�!�3�
�����-[��(�El�Ei<��|s��P�q��\���Q�2�2C�p�C�\�^:������XA�Q`�K��(qv��b�8���0�-v}-ڬ�mÑ���x)�,u�へv'��Y��U=qS�f�a�uĮ�Q�ay���/"�f���G1����u�����ͼ��������H--v36�c$g�ѱ��,��#qc8���,����!Hk��k]Nc�+H�R\��/@H�����kG@ka���M�Y-5IZ�fÎP,ˉ�˜C��Qe�3mIE�8��".��6���a��iK�j:��v���:wN��0�l��ٙ05�e�pV�5�����c��MJH�SCf`ևALJ�Df��,!�]��7J̈́&-¹��#f�=��uUn	���ݵ�VB��l!��x��u��S)i�7m����8��nu�7#���as�+.lU����R�BdU�tj^1s,��sSUS�qu�unCq�J��J��֏��|)���ےa:)q��5ie�����I|�>�~��/��)����r�s	���9x5���;�V��Ŋ\]v������6~�F��g=�����ac�Qʪ{�4�n��X3��<��r�9ʜ���<��C����T=+������ML���^O?�}�̥����{r���=W.��v���/�ܤ�D�E���w��z6��w�L��"�����s:����A������6��*�eyڼ�젏������Ɩ޺�N��8߈�@���'=��+>�W�?�H�_7AKt-ՙV	�+�I�Y�]��;����=c?U��2ˌ�.�9El�y����Ѧn��f�9�t[��ݚT�v�VK-�74`�lׂ��Wj��_G�d��e�~�D.�
����'zgd������$5��;T;�Y@p7���_ch#�h ~-�Pڸ�/]k���j��c��yH�xgF�&�v�jo��+7Ws7r�+FAh`w��}>3im3UV��X2��ѷ���YZ�Ӿ������I$��³���
�#�}��\��O�o�
���[��9(xU
�`��7i҂�Π����@m����^�ڰ=k^��u飼����fY`�yaS�� �K�</[�Q��/73(@A��� �n�/�wcwю���!��B�B�����X4T�ǔ�A���t�n�n��݇:�'�*��>Aw8��V뭗)z�S��?V�D��F��E_h�Ư�P�o�B�*�n��ω(û]=ۢ�,�C+WQFW���������J��|�t�!��_��W��#k�`�9���U���3Bζ��#�:�~-��-���-�+=����}@3����N>)u�h9�ܠ� ���-֧��/� ��!@�\��6���Y��}W��jW���\��Ա�\��)r�k{�OJ�H��H��Oem��}�-[8�M��y��ڵ�ٝ�[�j������|�j���y�]�`�������n��G�Y_�rfs�Ȓ�e�^!�H[A�~�1_�}��}����+锈`Bv�q�b+�f�|E�4`~4h��ݠ��^�z\ڊ�q��(t��wܻ��%�<�[A� M� ��B �H������[�� B��&���s��q�5�8�<Y.����jY[��x�1��N��g�} �z�݈7��v������u-c/��C�����4~�����@��!��n�?j���������?lBa���;Z,�?��o`~�A� C-T��P�]x�W_^Ѐ�)0��mt� �Ye?b�T���J>ȳ;6z�--����!� A�x(u���i�}2KT�=�{>��m9øg�s��yŝ^�����!~�Ó3FԪ���nZ9�^tܭ�ewf��2E0�1\�oM9ż�(�&%�9�j�ot4�S�{��g�J3��F/[W�U����}N��|�~����t��[�N�e�7���W	v��S��_o�5��s���_H�?6�Ŵ;�}�3OyP�f���Q�-}w[��tsq��8���u�*��Y`ʺh����S ���F�t���l�����>�|���Pr����^~�'6���6�?7A [��-_Ǧ���6��r���l|�PT�0����22}��K����@�.��pԗr�3��r�*"�|�z�[��n����՝P��Ռ����F�����`��O��@���7����_xU��p��X믘�A|u���u�{˦�C�G�Z��t���5Q}�0�}%?6��͠���;���L^�& ������6&de}�9������!����a���{�Ǒ�bk�b��E`5KZ���d�u����M�k�5�w�Uuu|��8,���a�Qvy�=���0���>���np_�0e���HJ�ce#qeM��Wd���cM%�M2�jwf��H�ͳ1-��!c�T�pB\��c�����͗[�nm;�4��p�����j�Q��7e��Fť�<�1�{Y`�e"e�#���������<>��gä[���<2L;l�����N���:�۱b˸��ua��r�'��b��}.�]�v;a��pA�'��}�~.0�h�'Uۖ
ш-���zN.�3G�]"U��Ci��n~��	ۀ�����"�
S�х�[�߼��=M靑.�"� אG�i|[A�|�.�[��%t_;���N8וR����>�y��Ar�-�z5�/U�M����V����	�HJ"��|~���ͯi�|2Ϸ/h���X��W��$oR���H�_7�	R�1䱿XS�4�{�ޯ��A	�N��ւmo����o��<E6���`�+�����n� ��� ��E���]�=����!z�zz�����G�r(9��/( A2W��~�����>���|��\┣M�B�1m>XX:�"�&���g����lb�f~��^x�A�A���h!�2�p>���1������17yNUx���ޯ�����t�v^e���A��;�����e&,�N��x;���x�}R�Z�FNfW/�n���T�i��0�E�s��\VT�+{T��� >}���B����%�Ղ:|��������yH��D?7����D����/�u A!�/���_�S��rϽ�.Ϋ�~�j=��;A� Ay@ \��t�!��_!�.��	J-��dA�K�Ca�'���j�V0s3��)�ņ��C�V����5�"�	�A	n�-ӻ�G�����{� &��Y���Qg�C���� ��"j�n�g��TwW�xZ���WF�лZ�Us��H,O[�¥�b.��4H�YL��$��@��P!�n�|A6l��N�Fm%�@��,OCg�h1�<ڍʁ����_��6�2�@�H���ݳiI��,⯏�_s��}��]����ί:x�Amuz�V���s�Q�{ ���B-�ɴ5��^�n���4l-}�)�l�Vw{�\�l��0=v��]��w�"���AS�y���x_E�? >�I�ᙙ�VP��O1�P%�":P��mt��������t�A�A A,����o����W�����r�a��̽�������C��Z���-��!��I��%��;�I=�y{���껻���ίA����t,��-+�}UG��۷��5�	�G�l��[Y%8�7Oi僦Zn��E��i,�/
�X�2���c�G�]�;�t_�峩��3[�Z�G��Ĭ�ڰA�r�x��:�K,��n��U�`�����<w���z5쮬�����}�AC�B�o��f���e��۔1�U��Qq8�s�s�6{���֟�"�j�X�M{�4A���6����?7C��;�d>���4@�g�q���u������HhY��|�yH���bKtk�z��v���;�U�!]W�	mUG[�W\���jT��5���T��//�ƞ���ؕ��4���ѥ���Y5T��5����!$�w����ˏr�yʴ8�|Ctn�~�U�����0�H^8��s^��#����x�PD�[����M+>s:gߏJ! E�@�M�[�k5�u;G*���]�����c_�x�4.5�`,k���(=P� ����v���ˬ����VZ�f�3��w����+����A�/�?�|�|�F�U���w*�2>b�:�tD���:y�@�~��؂?7��s�&e��d_<�6R��_7X$7U^�c�>录�Jf�]�֖��yw("���H�p�� ~�QC)��b���5�G�h/������zu\��f���N"*��*�=y�Ԙ�>������-�_-���;z�#���c���,rA�d���^����v� AyK�Ѡ�͠�6��>{x���{��A���v�g2a���Kؼj������4 MV]4��Л�gP��ė]ԑ�'u�漗��f�𻷪ѝ�8�T�phv���}�����)Y�K=B	wP����[JR*F�;EHh��
�!�$�䵯
u���e����6�R��Y�a�4A�]R��t!�pq�Vs;�g�]/.�M�ٶAu����9 4�V�XX�R��Z�W��V�r%%�*��g6�WJYL�K��v�P[�9���؜��S��TUY�;<�(�:���ǰ%�xS�(�T4���l�~���W�[mi�u��qk�lݍ�䳮n�A�:�f�5�N�nq�B�o���*��+PF� �E�*�ҫ{EN쩩d�znŖ#h�f3u��_gͯ�x���^�^��\,����qYX��iꍌ��L׼�H$S�?6�n��/y0�#�|�>� �t-���u��:��>�n3[��|+7O�*��w'w��y��"g,��r��r�n���;�z��:���� @n��5W�g�eMy�P-�_W� ~�;xv��_�S߫�����\,^r����7q���,;^��S}��!��{=�޺�u����ί|A#z����� A���>�?>O~����X1�a��8��r��1�<cA�H�ur3o5��Bf�qsނ|�����[�����]���S�#�(n�t,���2��z�zh�S���������G]/�?� D�={�}㘫Ү��Q[U��'1ݪ�_K�����l��h��Ij'	�֨_�f�����7�՗M9Cl�w*�������|s9��n�_���t� [���oEw5U��}��V������D��n��O#6Ÿ(8����n��u�t'������Sw�7��Qp��I��Q�+a[A��m"�ʁ�[]��� ��݄E���tG����ZAy��}~�������*�n�����"	��@��y��C�[^��e׻�[��L�V���'r�@���/�b'9s�w[��;w���F��Q��'\l�
F6j\��/b��4��v�P��mj؟�e�ޤ?F�����f�Ϧw��W��\��y��6g�좦TPeՀA�/�����+�H��"ۨo����6�ƫt/{ꀴNAx���"J�^��Ǝ0��Z���h wԈ?�E�@��:C��M��ر��\�CjZ�0l=L�p7���R���]ưjf��F�d�H:�����a�|�#��Z�{rm*ʫYUCn��TuLA�Wl�*��pP[���p�s��ZZj��5Զ�ݫ��q';:E:��OY�\6R�9���a-ZU؇+�^����i{[��XݽT��{�&o܇��,�N����&���e��u�tQ%�9V�(�F8Y59⮭�����[��Ē앷�P�v91R�sc���wWou"�_ۍ���.��cn�84�)]3r�_WZ�[8���ʱ7p*V�ܫ��>�C/��2��=�ۗ�n;+�;�y�$��Yv6����=v�f9V����0Q2ҥ�V�����s���Wm�5����Cm��5�,����زZ�]w�ڬΪ�er���Zp�wH���PWJ�R5X�*�7P�3{���t�NF����z��P����⪴���jŬw���w{U��ԛ.��e�@��j�����e�=��zE�,[O7jr���A\�tq�&�&�U���v,�Ś�{G������&��D8�8�X��u���qBae�]���a�����wX����X$xGv4�:u���X��u0n��D4X[&��A���?��*�w#���"l�S>۝�Y��ǔpoHk������m�M{�|!j���*qG��65�Jm�yT	�>^UϴJ���9VD������[���6�w*����������Q���i�j|m�=es��VS���c��P���3V&y���7>��P��,ծ�����	�6�/���j=�ec���Ú?/a�)�P��*�I�w:L�uی�C�tܹ�E-wrhwZ�r���1nn�4&��ܵ�4fTJ��1Uîu&ɇv�dL)��X1����1&Ɛ���A`�C&���0�s�a;��s��p���%��9� ��d)#A&1�PPĈh\��HL%Ί��@R��"]�RCBB!E$@͌�K��H&14J��	���Ewq�nn��	D�2��˙�a��4�9�d�]�ܙ�s�5Β�Ƒd\�J4v�s�v�D�FF"�U+�I}���w~�뿼��~�v����@/�q�H�AdWexn_3��Ӟ���A�A4�
��g���qF��9&�>q�GJ��B�kC2�`;ԁ���	n� �L��n��F�N��j�W��2yP^(�_�^R Ȃ?6�_7C���	w�}(����cfniL]����8ӵC�Q�
7NK�a�F֨j�,Z$��ެ��z�?|c[�$7K}���6�<V<�v��!GsD�\���?^PG����n�����G$��O��R���-�o�����]:坻ί�F��kA [���z���]lx�X<�K�=� A��?7A�/�!�b�o�l�$!�������Σ��~@��$A�i|�|�`#6��E�]��R����/��Ct����m�O`�ǜNP}��r�rS%�F:R�AQ��r�wնall��S�eg�g<z�&��	�1������nF���^�q��x4;�zl)^�k�¯]c���j]g� �]t?��|�����[���?7I��O�J]u5�<A��N=���k$�Ϝi��Dk��n�@��e�a.�_��Ŵ��c���~/�3sb��:��l�-�,>��im�z)�t�ދF��,�/�Ζ/��E�(���m�-��fOZ�3�����Ǟ�y��|�U�G��y������� C�ʺ���s�x� ��A#r=w.m�O`�ǜNP}��;��ź���6;�-S9�Yl׮�;�K�,����Ŵ<*<�g�^��cO��]�],����o��t0�Hn��%L��qqW���Q��q���������iس/�:����|�k1�th?MK�A|[�A!��6�-�M�}LZb�x2�F����L�囜NP}��;��_W��[BE���m֋�����^hWu��N���X�zc�g�f%;�zZ�d�<S�m��{�aV3-�בn�Md<��;v_�\F��pM�VɄ��['�<b�5g�As���$4F[s"�6��*��s�[I1Ҧ�XkSlH8��ո6�Z&l�3U�{m���V�ػq��.�Ҥ��3.̭GH3�q�^��5k4�����^OO{A"���"R�S!�!�A#R�ذ,і�2��a 7L�3�\b�k����D�:��n��Ŷfiv��lp��>~?B��c��:��n��sn�����oc��C������	Ѧ>�S���� � �?]���X���s�w�#J|�Hm+#)��#]� \���� ��|� ���@z�Jй��k�E�C@/Ԉ?z �W{Ь����u��_mׁD����]A�G^�o�+����H������7Aì:�1���9^m�L��78���'r� �_P_��_�������˶��]H��A|[A�����~�}�]�>q��El"5�>�3ndYw�#2>o �A|A-�E�V�A��W?�*�D��/'U[^�m�3�P%�/�?H���Z�����#k�v�N����[cI�����qkL�i30Yt����5���VY�t֊S_��L�m7�9���,���v�{O`���s�/������,�x�\���D2���|E���Ƿ��{D�d�d
�������{ކϐ[�S8p:vZK����{�~�����&����gbK�3�T��|>oů��B���Ϳ-�R�����_6D/�%mCؾ�M>ߵ��Ǐ��o�h�Ǿ��L�Ks2�ȃ��F������×�	T�8gQ��=*o޽Av��TL�ѡ̫@�OiD@2d��_V�l�7Y�xZ��
!� N�-�@�j̸��8���u�*�$W�D�OP�z�7��-����[��~�e+ί���D�Ń%/� �)�{��{�=T�v}%�n�k�%�]tKB&���)qP퍃T*��,��5W�R�\��a�w�."�fe�L�>{�&}�6)G�y����@���LW��j� ��A���$�,�_	+> ��a=�Y��~�JD���M���v�^��Qg����=�2E�[S�vT{«� ~�@ ~/Z��#1|$�����K�z�`��)�ٝzĲ�+��l�����ygz�*�8��գ�o����Z�4������:7��ov�e+��5��F��y�G�ר�I2����������㬝��ӏ���/� k�����%"$�`�q��+���	���m��f ����٣b�{G���@�{JA*fnb>s
�����{�_�J@�D��"Ib̕���tߡ��2SN��nSyr�X�z��!���	{_��+��$A�x��z7�����BZ11+�#%"9����\�7q��(�m(8v���l>p�ԗ�߯}�OR�"_$�a��L�[��}L�W�^{ΈY�����)��b�z� �$�D��%A��3}(^��(Y�j� �<�;[��7LTG�œW��@�{JH#Z�f�7U�73���Q���L�Z9��@�HH���>��;�y]�Yr�.��]�\NP��@#�_I�A ��P�[^��UY��X> ����+�"�m����S.��W� ������j߹����q]3Z�'R��r��C���ߴH~W�	����յ[�q:<�譵8<=��Nb�mn��؀na8���UV�w�s�HI���=R���Zff�.e+�"����y���=�;���M���^̮'_�< �j���#���XI�������=y���rpݛ��92#�����3T�����5�	.��).���M}�Y���AmȐd @̅���~�؉�;'	�	���c�w�P� ��@����/� "�e����-��r��;���q�D�{|O9R��W���7,Y���Y�,�#���)H�v,}��2E`���Ʒ����b�U[�4���d�����ܥ �p?H��D,)N�=����đ�[��"N�|�̍��zkN�o��F@�f�&m�Y���my/J��� �����}bD�G}�%����;>ϒ�7��^��9R��W�$g��ܿ�� �D���
�
�}aV]���-�De�If_-�N=����4]��{��U�c��9�Y��%����=Oof^��v��/�%E�&�`v��\�r���t�����с��$�l0ڍ�z� ���1����$a�OR�68p�!z�%ԏ�Wʙ�x��]nֶ1/3fw��ņok.����Ul�[:�q�]/�Td�Z,��öJ��2<]tk[�mَ����Ƃ�K��;�d��d��ݱ��Z�:��m�,�,
"���Gq8ʋĺ��8���9�V�f��N��C�����u��͖g�؜�lV��S�:R�6㵫�:j��n�K}Ϗ��/_�H����"��2 ���x7�S,z�:���O/wU��f�^�x�<���/��ř)	W���ۿqq;�����-�R�N�N�0z�o��TA/� �*M�}���i~�A}���(i�D��!�[v"��W+��>�R����$OޫD�3F�2�DLʱ32��ss� A/(/�>VA �>��7�Y/Ư;���<}5}�7��Ctt�a�5ۗ�����DLʱ�ѧ2���}�0y��RcэO��V+�"�r{�͠� �P@��"�� B��>ױ����fm��\�%к��֋�s��ʦ�1p��=n��Ua��n��m4֮��w�b?f\������3$H|�c�ڋձ�Y36�~"�#��Ż�����D(�%�?( Eo���}~���~��}d���BeA��V`g���]��wR���ʮ��+.�
�~����n�p�UU�DT��teePf�2 K�KS����H��T�A�#�zr2�W�t�����6����Ch"0��ƓAW�b��݄A��−!)|Af�5��p-�{����^���U�Й=���AǈFH���� D0���n�qR��t3�5d����fd��ӌ�ڵ�cԲf&iƂ���_OP&s�|=�����|����M�E����eꫜ�T�`�}�k2���e^p���5�(_�X� ���K��7�y�����#u��kq��j��k��+5���66T8��E��k���#�lFo�ѡ̫Bp�L^譜��z'Q*{4H;��]u�Pψ#Մ#�yX"J�a�H���Ѹ}����D�?k�(ni�[ڸձ�R����NF���+��=�E�ކ�����=�ք{�-�ı���G�b$�_Z��n��B��DW4�W�j]9��,.<�I�d��Ϫ꛾���j^��1]oc��t�̄i�����6�x�ο:�K�)��MEw:Ҩ���7�v���?��X����U�D�C�D4)|��q��}�=���b�����(p~��qw����	�'�����{����y�ȳ���C����X Ȁ�]e˜n��q����{Ӫ��k�][�]���}��u����0�w�4Z�{(�QY8;=q�ʛz�pq�n.|zV�pc�2�q������\�w�C���Ա�˚��[�z	S}��/8`�!~��h�]>���R��M��N�eD��s*ю8�#p��m�a�c�*�Ϗ:@�a������6iu�NЙ=���@!�� d��ds��Be��N' �?lA�����%��5Q�iK�;<��J����_V�wuw�^Fz� �����D��"Iv<������𞡦tVA �w���޼c�3��M��j���VS�U��V��ub�F��k�w��g,��12��Φ֛�C��Y��o=�t�Jc��U;Ye^V��ӥ޴�-�7W7^�MY	l��$0~�_/�����I_!��ř)��|/��q������0�NP3ٿH �@@���+I@�.�?z㴽/����l�y����q�>��h�H��M��"�g]g���'�/ A�������D�D,zzWR����^��Jf�h!F�� c*4�r#��g�HAR"H��d��(Erī�Y6f���D� {�����>W�$U��о�� � �ٔ��$Dm}U��z"��K��ʴbfV���\=���)��F��;Bd�~3h A��PFH��$_	(_�Q�ng+����K��]J{��+ٱU�������"-�@:dz���^����_AԾ"Ib�?(���i�6�=��^	�i}[Xӭ��Ի2+>����)���J�I,`�{��Ev�n��=\v�:��9�t�c7�hVJ��꒓l�Qɘ����ݩL^<T��O��T�1�Ţ�*�/\o{m�a�v{���c)����� �����]2�U|p�+�[[{�X�]�Q@�}���j�YV��+iFj�!�L�ɮ����zo3T���Ī��'XLR�í��X�� �ܴlWsx9�㻂�V���㣅�q_vNU��S\«�22��}kj����n��!r�t3"�B2�R�;]�K��W뵤粛�<�]�TY�J&wNڵ�)�Pjd��4A�{jH:�gNe�Ɇ���]v�ÑU�����Mo
��5R��� ٺ�ַͤ�M�}�9*��h��իe���lO)ْݠtN�f���.ѻ�T	�2��������������1�=��oY]kf��ׯ�.�w��=I�Z��n��XUV���ݣq[Ӷ�)�������^l��q]�5�R���7[���7
���]�n�����ʸ��m*�J"U-�%e_[ɚgU��y�3�ۨ��pY�r��]��n\?�ɧD���09�X���mE}��^J��u�K6�I����R諾Yw)��{�+�2���S!�Ug�v������º�GJ]D8�**�/)�9�6���
���*曫M�h���v�x'�F�fjS�e��Nc�c�õ�v���M���b������.���[��XyV���m�ެ�j�-�&?�������l��x6�]�~G`1�:ui�k�./t��Sta���"���mZ��<�:K3���Ρ�ܹ	˻�&��D�#0��1����DCG6�H�;��h��I4�#�5�Ԛ��Y��"��� S���)�cwW"2�۹Ќ'.0� st���Ӻ$�10JLd��#(D�SW����e7Mhɡ�Q@II��gw�� �.\��"Dȇ8�F�����e	΀�Fd��iG:#K4\�F4X���!�t��Jh���ݢ4A�E&���wb�p��+�v4��f�����M2�&nnH�	@�)�.ErL�n!P���sr�:㣺�T!I	$dU�w9�&l�Ȏ�c$$D�F�#��ADS�_��_����M�)�e髜���ε�q�ą�+���L����J��;����Zla+6B���-����E����n�pC�sͮr�U���������v�������)m��3.rk��ӱ�P����=��YXu�"Vj��%a�.�VnR0�\�4&�M6�o	]��A�iݝ��k��`kf�䎱�Se6�E��!Hk���ֱ̦C[�����$Jg1�����{Z5�v��c�.|�٩���廇s��{\l�R�:.���M�]�q�ўQ��V�wm��,i:i��6�Wb�:����6s�&��Y�	���lI��a�-�7l�F�%���y��t��x\����E�yXw"7��-�8֒T��<b�\0��v��{n���w�]�o��B4�7@�t���ؼ��[�NKF�����QFˈ��s�����ƭƅ8�A5�[�KТW[:����M5�h±��r�_Z��N���:�.n[nؼ��k���N�c�Z���{t��޹�a��:��6�՚�x��D�hk�K�k��"=���S��k]�!�b��&�ogW<�5��c�Z�c���VXG\] 2�M8�vdl�K�֎]0�iK���&K���{�8J���{q��+óJn��v��e���g�;�t�I�v�մ��jYV˞6gHe��,&��:�,�u#mVێ��&
yۙ�2q��y2i����dct�	6�;f1s�V*����9�mӸ���J�˶	8;jx�xSruģ�^�������k�ɲ �n�њ��R�6ja�t�e�7>�LIF��&;]�8�<��ׁ
�a��{g�0ӌ�XݧU�,�Wg�Z�⬼���b�S�V.�V*�rc֌��A���1��;V{q�]�0��ؙ�r��72 -窙�KjU���L::�Y*�� 2ʃEi.�4��VWs�q��!��i�Z�E�uh�:�v�me�;�y��;Z�@��C�:.���&͌b��Q���wm�ֆ�I��<ZN�u�X5�L/�0pnQ�݃l2�`�2���c��y�H5���G�w �U�-���9WZ7��h�L\�I7pk��wJ����^�1���\���;J�[�,Ԅep�by{u�c��#R��e�6�Ǚ䝮MX�6�Gcż���7�}b��X]x�����H�mX��e�_����C�d]st�]u6��Nr�P�t��k��Tc���S;��� nB#[BĀ@̅�^�����;B\��ǃk�gg��r��wh#��`%|$ϐ&H���;ܽtjn�������������z���j<�i��@���d�`)�^
^WcҰ�b����Z{۳Q���2������e������zA�c5�[��|͍�\��_�_�t����I,Y��!�u���U_m���>`��A�zVh{�F���9�3h/��%d��%�P�����G�_I�� ~��:stx������=�JJ��[�j#�~����"۟�"� �%n!a����X���qUvAH�T�x5�۵mf�S[&3A�:jێ���7B��gx:
�@,҂ ���X"J�����m�]��l�e
��X�s��ZA� �?{���,Y�� �%|�گ.�')P�#{K"��t��f���5J΢a]VP�m%d'����Zm�rЩd�CM��f�ݕ��vn����'������/� �Ѕs=4f����jNl�m'��2D=���X�묎��P�A|~~H_����&|� I,=���!�8iE�^r��B����"�>X܉2R���K��Tw�K�m �:� ��?H�ݾ�o�����ucg�<��U�r��w���m���X2R$��!`�^�K/j�a|Gu)�0����QSh����|~n��� �"�U^ּo���(�Ճ�� H�d�m5z��l��ř�J���(#f�I��/�-}7�#�b㙒:�E<��oURם+�w��-�y�֐fz��})|A��)$���!�Lۋ�u�,�j�=�/�v���zϯ���L���欂��Ow/�jz��꽱JD'��$�`�HAT���r8.�XUz2�y_�wLx�p�����:��8&ɷ�P�Wn}�d��B�/&Ɉ���W�*;uУ���]������Un�<������=���iW��CqWGFϝa�[�Ig��'�G��٘��W�ŷ�.gi�B��8߈ ���{v����ԴYͤA!�DI.�H�d��ą:�HsH��^�>���g��]�)����V+�%}$An`�=����Y�M�Ww+?]�.����u��t�ӫ]�E�nϠ�h�\1΍�+�����8��@�)���2�75��t�p�	��a���]�7~S�������~�� "�~卉�φt=��;��:�D��h�ot+��b_�G� �=+�'X���٦vˎ�9� Ct��w`�( AJ"��kw~<�^��W��͜wC�ͧ�'�������tA�K�$�`�K�;_��O#ȍ"f>�-܉ �G�3"���ͳ��AJ�Н���9(��Z�F-z�}��Y�ef�0>�X�~Ei�O��b����q{}�2��C;µ+�}��45��9�՞1Ku�W�*e[��w�$]�C�Z�ڡ�{W�' ��D ��dA���Gk�6GCe�c��ׂ)k�
���B�����_َE�+�����}����4l])i�X[4�T,\��׫-�KBg6%�3��Km�m1�W�d����9����b�V�{s�4?vm<�>�B������\̮.u߯PG����]���2��fU��=���dE�����7cq��η1F���;=c��?�";�`��) �݈/��_�"�%|��Ξ���s�W��M�����������d��� �%"$�?q���f��T@�;P;�}?f ��k�����ݧ�;�(x��4�[�G6f�g���~����h��U��fU���ř)�e]f�I�chh#e/d&��ޮ��5w�v���@/k�:��(��w��[�~3�s2R;���8.�������=����1u7m׶,��'����*�_�����1��.]I��xVZʡq��#T�.�Ձr�Ũfi7�,]-bq�Tۮ ��d(M#So(� O�����@��-ӄx�GX�����l�m��hFb���Ę�v�uts��hV�!I,L��wM�F\�T4����:٥�ie���XF;�kv�E�K��Bj�2��F-��i�&�A&��6X�KA��Y+l1b��t*�k&����,uo�p6E��O��f�����_>����01�ؘ9�e��F YtU֛jۺ� �1�.κ]�m��� ~V���?I_/��,g<�Ww����o]�^#~�}��kc���
T ���Y�R 9H$�( B�̬q�3�����`���m=>�z�=��7��7��#��ӭ�>w[s����C��q�,��s*�h�m���x���D�vr������a[k�����:S�X�6nڄN��8��3$N��8+v�%7���U���[<$B�x`)�H,�K��{ԁK��2P�%d��Շ���+V���t��	�wn�f�]7��=@��_%���I�����0l*�WwH���\
�=.�/WZ��fN2��N`$���߮F'r�"w;�Q̫�fU�έs��=�UU�a��������W<0��>�.yX �"�I��"�Go�LX~��:k�Ƨ�]��z��^���t���i�M��5�K-�B��k�!eɆ�Ζֽ�4n���ow<�ns�V�N餾;�"C��pV��JoK�4�#A����,)���r~=K�ǁԾ#_�X'�A~2PFH�~�W�^�'@�9R�ٳ��;;������+"e�w�Ѩ�T׮���͝�n#5�hIn�Fd-�]n�s�"&}�P��`���O����߲�*<���~�|��/��@�&�z�t�Z;�[Cד��ݰ��.Ҭ�������,XJ@H��9o}޲�.����F,�o>5ь���I��Wq�-m��\Fɮ���&�p�礪�(�^e̹�2�z���[��*vw�;�1�p�nvޞNn+ �5�?w%�_�V�@"JG�C]���_"�=8������������� �:� ��s��%d~B�s�,G;��fe��R���|�k^������Õ�/.��l����Z��\g��-7(�}�_[ƽ��˚���ī���fb�c��SG,�º�m^�.ۂձ�M��^� A��J�̩��W�f��׋ю�UG�ݢ�~��(m��w�=�v'���	��3|���̿e��G����l3�b���X�d��%}$CL�wuV�3��"-�SoC�1>���7���� �{� d��"J���|$B�H�}T'�#ӑS;�lh�B`�L�KTN;��n݃�&�л���b����}e�3.\��'�]�d��h�V5�^U����{�{��U?f�o��E3*�ff�1̢��a�!����(^5$h/�Uk��zV����>��o��%|$5��v
;ݹ��$�e��:� �$�mL� �9i���}N�/H0�6�]DA�̭�ݞ������$�����ӽ���ih7���!����~bR��5�Yip���]����4MGVj�^s+e�9�1�n�X��L]����j����rl���uK�`�}�
;�lV������RI�����( d�z����~�Ӧ�#ڐ�T��7�n��9�	�@�7��(i�_$�8�y�������Wh����U�(�6bLl�Zm
��N�={��\=m�X9+=����G�����5ʱ�;�+w��{����̭��=��3E��l���CA��@��`�"�b	�+$1�N�Nm��hG�n�ڝlz7}�%cY;�]}�|Y@���b���x*oި�T����=��S��љX��e�"��G�M����'���sfdܡ0��V"D�>��������Tf�e�;�l�$��.D��� �p��b<�q��y��:g�^�����c�4��C�"B ��@C���}��<�;�{�s����hIX�My]Ƃ,��}�X���a���pwj�AR��Ƞ�s�K+{yA���̧WaV!��P�ۻH+�;��f_=7Gk�_�^Z�4�6�F!w�K����uA^�� ��G]j�F�b�R�0#���<���s�D�=s����R]�����2����s��X����$�ɓ�}<����CG��s�{U��;U�G��`lܑڱ�7[l��l���яF��ژȸ�۪�Ž\�uۜ�u����|�ǌ�N�͝������>��d��l���cۍu�;��Y�qפ"��X"P�����-���IB���6��u�h[�ŉ20�q.�m+�!3Η�`�G!"��"D�~�G�ٻ/ �e!���9VQ����b`�s�X�z�33F�ʴc�6	�ޗ���;�n����>E�V�I�������+ht�<��� d�V�Z�MTq
�$W���@C0}$�×~v�Ry��½��$Ǹ��~�_k�I_I$�{���eo�5����%/M�O2߷b�=�BI�;|��MU�h�R������L�H��)=�t���k�{����^��:4/7+zg�yC� $�h�M4����~���2�v�z��Hc�7)��Iڕ����4tͻKF�&���5���ܞ�}{��|��H��Oe)��T�����$��4p_f�o9RD$��>��������7.�h��_:� X��в��z�]Ǫ��j��Cr�n�[��}K/�Gy��3��6��;�F	v+�U�����R��>�m�#Y��{���%I؎�<Efu���휾�/�����.��ݯW�2=:�j^���BP�ܭ������"J� ho�]l�*�x-Ͻ��τ��d�B���jj�:��!M�^k��n�	"J�I6�Ӱ��	�������d�GI��}%IOR::U�n���������VQ0A�X�[�-�2m2:�Ea���H��&
�J�
����d|31��';��L���S��"" @�7�٬����d_{��$�$��j�>뒮���� 'w�$�R~�*��z��=_l�C��U��^��@>�`�/��uJ�9�Ґ�ax��iR�ٛ���F.5ٵ���&���fm\�v˝־�Ou��6�Rӥ�Y��wYM��n��E�f�"gF��V�ۼ���=�L2N�ج��ל6��Nd�OAy�BF�B��w��B�i:sW#��%�L�{o�-�ە�ދ�kz�e�.(/!������)���eJG�Uk��-���lh�r�g}G]-ū:�����]]K}���d��^9�{�-֝N��+ڤ.]���ҷ�������PIu��}�B��]���e�x"��5���[�$%u&-s쫺w�W*'��q���B\���o��)��+4�úg�n�oYȝ��y[4ʄGֵ��sH�ct Ӈ�3~8����Ղ*Y4^�	'c�Pm*��TBL�wa�7p�f`8�UmZD�]R���|M^��f�9{��[�'��5n�,Ac*n�]�c����	S[��ҥ�/���-�:�'yYe��N�ީ��7�K���;h�ٵ4����3/��+�kD�b��Վ�΅UgA��n���F��g/Q��3�U�K�&e������:I�u�>OJ�y��[�T�oC�F�+����&II\�r����Y�t�n՝YlZ4i�}����L\�n�wu�q��L�ݦ�S����������ý��yJ�r���Chr�K;�<9�n��z�Yٵ��t���S���0n�ב�L�z�ԛ}}����%�򖳥�ߌ��p>��'q���H�+a��/h��w|��>�˜��û�e�ݷ-(a� ���:b��FM��n��0�22Q�Ō��r�F��0cIr�.r�ݻFM1\��9%��S%,��m�!Rb9E\�M	��DQt�1��$�'7hA�!$Ě�*-BM	�%0��'w\��Ih�AWwcwr��pB�Q�A"�6�	�9r�,��&!$�E��ܮ$bdQL��A����	,hƠH,r囮���-���9wv���3��ccKF�F]�ሬTV@��!�Ph�C��b�Z���I�Fdm�%d�r��I64;�Nr�Eѹ�����&�sr.��1??I�2�d_M��Wi'�y�+�"H�����i䆟�Ɯ�"؇s��vɑ5^�s�>�E�s�jeǄ<w���zW�D�|$�&��,�k$[!i����ݜJ��X3G�k7�t���%	'�˱����'��G��]�ش-&��#��a�<��J�������c]	�[��F�x��m|��D��۽�j���d��"I�)^z�M5��6W�7�O)$�$�u�r\������;a��ͽтEMyS�߯���H��e�FR՞�][�	�_	$���|Mdۧ*���K}~��fu����ݓd�$RE������]����BJ;w��[�=E�t$��w��F^[)��Z�?mr^�Xj���7�\٫��Kq[�r�s��;V9P��+�����8x�����a^m=�N,����ٝ��3��_OE%}$BI �Bu3�z����+f���w�6����>}�MI�kz�����hYEQ�u��j��Y�y�,%��]�\�	i0�*\��e?�n�x����?~���������6Y���5R������h��o�wr�u}$BH������w_?#��=�&{w���מ�b�:��k����i�C�1PK�e}��	"���Yˣ��;�?`�cn^��vK�ռ��+�9	"JE�Õ�2��|��r��#�D=��ϲy�,�Y���9]w����L�vb�ve���� $�I���&�xh��������eE�k��z/�I2I�?F�ª�I�����n����0�R��}�m�D�F�[mf�x��ՙn��\�Δ���lew|�~|��ߞ�m����ծɐ���5`S/���v"�B	��0���:�e�N����k�&PW7VKB4��H��/N=�����>S��u!�q���aͻ���s�t:���,m��ױb-�nl��5,��>A�x���2�
{/���4�(����kn9��c�M]Y�;�y�M�X���]r1IslZ]wv�����U��_�ظ��HF��ʪVGE���ٞބrMʶ�m�F7Ś�j��O���g)+�"�r�d�޷d��[�{���Y;�Xx����%I@���eBso�D��o��N�j{#d�����I7��Q�:5���_>���I�I۔����o|1��y7ڶ���T��瀞��$@I�l;�n�����f��BI�»َ�z�˫���<�����f7=�=�I$W�O\�/�v�~�[�>{�&J�������@l�I@I<k����|=D��Z���e��@�iX�[)rA���a��A�&���-ۓ�4���@l�/��;��<����]���=�6F{��>��ݡ!$RW�IO�ڍ,��'��o!��
�U�B�h�/b�JYk�fUU��nyj;3�.y�]�v�(!@�s&����nBp�i��㴅OL�~\�yy�S��f%{{�x����$|�̛=X2��x<��_I�J�)'�q��=W5R�:�"`�k�u{=��6E%$�h=YK���bP[�wP�3kj�c|gr�V�0*�~�	DZ����q7#t�0I�I&�_�k�w�ź�
�=h�^��ͳ\�V�y~�w $�}%{_�ek��TƄ�n�	���:�`'�䳢v�۷\��{b��C�	!t��%=v����I�I��v�7Ȗ3*4)�ǧe��Y����;I��ž�$@IPt|�)��[�z��Og����b����(k�o�}ң�ؐ��FٟwS�I0	%�y�W�%ưY��z�]z=�8�-5S�Z��hX=U���֗��c�����9��,{.�5���X�bݾwt(�fb7��Nͳ\��d^ nW�I�MT�S֥�Ɂ}\��H���z�o��i�Wq�n�./n�������$��%}$RI�yY���ͧ퇅o��y�������=�}Q�������������j�����ti��>`�x��i}�խ��&�ɦ1Ԧ�UL����ޜ�$C��G�j��۪�u�"�ɂo����61 x�A���JE��M~�����з���L~w�o}��&�w���q} fX���w ;��$RD$���u3�1���*�7�/�Z�{�$_}$���79?�:yt�$C����;ֲ�]���6��/5�vx/��9BQ�[��u�Y�nߟ/mӼ󒬡�42�MM�W*���uI���o���j���=���T��]��$C�"���y������Z���Փ|4p�O���﷚�k�I@I������~�v5�h,���:���T�m�ۤJb4����uU
	],��~���@�I�J���x6��D��כ?%(�7;��I� �c����e&���_{��k}��e˭��������gi)]�'���t/�7�	$���K9�ڊV����
��X�� �Ow��o4����RDqe�!�;ݗ�n'"�I]3���z�y�����������W�Z�{��PD>�)+�˼�Nu�,��{�W��M������u�"���};��! ���E��Q���h,�yr��˴2��S.m�t�-����/���e���C��㙥��.�!�n�P�댊�F�3|(w5;0n�A:��%T��H��ӑ�u]�V�;h ����cn�*� �n�8[��6)���Ba�*w�E�Ml������^��t��kXl����b�������� j؅���e���ut]�ûZs�q�5uxCm��xPF��/�}u��$�Cm�v^��Q4r8<�fu�yF�f붗n8��q��&�[��{^�a�KYn4i������S�g��� �ZŰv��\�#���C~	*��D.�CR��{b��� $��ޛY<�$��������_�?��t�}$_IBۯ��%�¯�3���'P����9��Og��|�}BH��j1��d Z�L�_I��A��_��­�����ثvE��hT�����\�mY�v:zI5����s�8I��]���ڽ�^�O�y_o�$�%I�׈��	��³�F�g��\"{=�{�:P� $�+�G����OR�)�ݛ�"6���qq��WnǕ�kێA���B
TB�2~���\h��>��̌�O\h��ӻ �:QU��-m�\��|a׽��*��I0I���&�4�!L���e��6�Z��/�L��*�L�_1��(�3��m�{t�5J!�s0.7j<��G\E�oW<��ݮ���\�B����t���k=Θ�&�w�Û_k�#
��J9�_�_>���	"O8f��5ԙu��<�.���{=p�rx�@�$�}$BJY�/#���o���ukrf/��{��=ҍ��y_x���C{�~����$_I����WRh�m�޺ʷ�<s=���<>
�g�6���$�����z���%j3D�B����.��a]���<��[r],�`C�"�"�k�k�<�$�$��}g��]vz*���l^>\�j�~��/��	*H��W�����i�ږ�%���' ƞ�xS��{�2�j��+�<���N�s0�3�M��_}��%	"I{����w7��+>2V�Q��.V���3�fl���}L���Nܞ��-���\.^\��L��;*n
�B��]�����]}�\oGc�Lp�w�n���	"^]��pg�.��X5}:u���\�w\���g���'�{�(��Y������q� �RW�D>�Hf�{�\ݾ|2v?Wnx��7�ҳd�|��}$BO�!��W�'�����
�YTJ�����%v'���t@4�N�]�@�iB�AH�]V/���LD����c�x|��}�e�D�v�4�����H����7��=��|+��uҖ���^�<�e��)\%�O=���$���g��Q��f��^W�k��$RT���o^}%�W��6gX���%{���II0o�ުʣ׾���	#|�/=���>
�g��wۨ�<i:��*��T��/�v�篬 2Z�g�}h�Uj������康w� �L��3�S�شu�}6�{�;�V��^N���bh��jj��w�.��)"W�I$��o�S�=|0u�I9���Ş�\%�O�C�}$@I)e�0}���&(�L�9eۮ��,q211�Cuq��h݀n�V*�{��^����� =�;�ݑ��̍����{�͸�����oݠI@I�I�jX�_��M�{���&��ڨp�T�
f�@wk�W�fhձ���_۩��ýRD$�I�_��[�sU���n�����+����_t�$C�$��5(����~ �4=���D:y�}��\0!��%xnP�*7�W-�E~�_OW�I&�%}$K5f�ǃ���ϼ��}���k���>
�g���)(}�(O�=�� qE/�Xe)C&��g��;a�i=���K;:7a��hh�]�˽['�ML��U�Y�#Z[�wX��x ��
e7N��Wn*3wՔ���v�"�r�R����у�
�T�p�ٶ8s.�fek�]h�YZ.���"(�A,�<Evqu�9r��n���Q�Cmp�8�v]KH�Ss��c�o���t4wTAV=s��.�=3秭V*��Q5��;O�3�]�:����q�򓑵y�B��Ⳍ0U���Wx;��EQ"���ۼ��^*�uO6�����P��A+Dٗ���˻:��sDU`�B}�1�pf1�g=;��r�Wu%U�G
�ѣ}��D5kX�жz�}<R��`�x�˽�/&*/�9�ä:�a�Vh��ecQf���ú����^aN̏/l���V�2<��7i���N�X�<�U-cګw������9B�.;�ǫ4�@�y��͆�ŷT�VU�ac8sQѰ�J�u���G6kN�l���iC�*6��Y��noZ���O�^2����+��H3M��kj�[~7�39�-1g��ٮm�8���n0K�����u���t��}�D:�Pgo��8�������X��^/��v�3w�sM��u�d��]|���׷�h�Pܹ���ن��ɫ&���V�x�S���	��L�Ӌ��w����4[���ѳ��[d�_w>�	��틆��9��^S�������yW�Ýg�T7N�̼����M���2S|:ƫ=��ٹ�h���?7grfwn]ӺX�m�!�(c�bƍAF"�F�fh5�-s��wrh��D.�ƒ��(�ssD�ܨ�5��ݹQ�%��A�F�8%���I.R�ؤ�V*(�d�2�,Z5&��E����DѢ(�c�ԓ4E���Eh�*��QQ�MQc`�H�b#DPDPdɬd�"����AԖg7IX�$�ŌQ�6#Fɱ�h����b�RmX���:h�J4ȴ����т�ɨ��E��d���"�4h�CQ�lT2�6@�X�\�5�
��Dh�#cT�=o�U?�y5�(����h��,�քa�Fbа�thbk�Yv�`��lK4MnS�9���A�0���'�y<������!����df�i�����*2��S�'l�+'99����	\jḺ6}T��DĪͮ�H�\!��U��v��u$c�9�,^mvy�p]����R�O#c��X��[,wNe�.nu@[M�2��;G�b�n�Ma9�P�C�72�b�g��=��2Okq\;��v8����ع�|룊֮��:*��cn6���m����g�i��C����u��Kl�9;Q9�\�f�9�wm�d'����m�Bʦ4�8Ѫ�s�5��m1�1�E���h�v����QJ���e�D\T�<Mnk�8���-��e��&��1��gPd�q�l�Xk�`�8.��v�-���=��kd��\������ے8�;r��g�-Y+�������A�zm��� Kp�㛀��u�V. d����u�m]>ؔ��]�ݡIC�9.�u �Z8/%K�mʸ��nNc\��;<�d�Q�v6�c�W7�b9��b:ˏs�ٝ��h7���e|JFĭ՚S1]�ٵ�#��x[c3����t���&��1H.���my�&^<v͓����xx�4h�rSg^ҋ<f�ISz򛖓h��K�a��׉[��������:-T]7/b^���Z�^NdJ��S`,�i�������>_�S�,UV6�;+m���if��טFi��6���u�E�g�X�"qw!sm��ӻruq;�w����G��V���v0�v݀�vۤg�4�MDG$���KXK.y�H�����N�"�"R�R�ݶ!A�j�;��sƒb�f���\չ1s^�эٛw)X%v�5��i{,�e����'P�&؋yu�W�\Le+dz�v���Է�gG<������ɫrݨ��%^�]x%1GmfE�ћ��][=zk�G�ly��	A�9�����x5u�u�2gc�������LC�w7b��,��e�ˡ�T��:Ν�Lm����X�L���5�{/ehݗ��L��]*k�0˸n��vy0��5�0��	a�v�b��J6����M�b��!��n3k\Lhv�/&���W!&��J��k�ш�rݎ�ԹPѦ��SlVj�І��������$�i�����KZ�\Tmzݺ���KIj�̜8�
�FłE�j������褊J�G��I�[Y�����Z�=�矟��tC�$�$�䶼<�]W�ǫ�c�m �3�3����;݆{���NBHk�'���T7<�{�P�/�����5���ؼ����m�w��9��I@I�b�u��~y�=������o:����k!���߅֪��85��7W��f@�H��)�Ni�y�U�[����z{==^� A����Βl��u<��xЪ�fz�ps�؞m%� s3�ƪd�t��Y�l?�k{ŏU�b
�" &:���B�3<f+��^���l�]^����SE�3�+�#�D�%}�x�w-��畮9�I=bnOj8�|s�a��x���pz+�a�י��}9�֦Q������M�����ܠ���L/�~R��C���؇u{��u+2{.��+����|�JOWB�ú���\�=���E����ݯ{�Y���ܲ}�w6uy�*���/�n��NRD��|sM�xm������+��&����'T��h�0�w+q'�����{�� $���I.����t{��U�;n��{7�=�$�I^�A���ue�j��
ՂM*60�G/h���j���u�����;'\���޼�����0	"&w�_���⪫{�c#׾Yy���	�\�	(I�D1.dk���@�=��y���Y.�z��}�v 5�$�_�������9�_zP�)"�9VM�����T~Y�f��<��|�jݭ76�^k���]/y���vQ�L�ͱ�5�θ�cF�W�wv�N�.��p@�{ܫ-UJ�VC���ͷl�G�-�ڗ<�����=��I�I�G|ș����)����I���]��^j�Su���w��TE8��-��BH���(I3$:��H-��^ɛ��Q+d������"��D����K}ݫ��uX7f�����R�S7a�Vˍ�1Z����۶�;5�k�n��tRD$��y�}ڗ�"��f�.�kw�g���'��'`E$�A��jUASX�Ɔ�u�gu괲�)��������q��ȫ=���+T{�s�	*H�J���[;�=J����jU���G��\A��I$ГH��&l�j*���#��k��U���d\��=��򷏡�AUxIg�a�ޚݍn�iK0о����y��\��*j�f��.2ì��R`N�����mKo[�`.��:���g���!$��	��9�^�������߽��T��7\��n��r�H��dW�&o����XG���C��9�1���J�L[w7�*!�L��hP����T�7����$���~�Z�'���������G'WA��Bu��H�����Q�ת��}�k�W���y1y�R�d\�w�|�T����x���ٴ_�ف�_I���@OPW<py�z�|{�R�T�rxڝ�H��$����=Y�+z�ѱ�_w��1��U��ԫ�wK�{�z�}���u{u]̞���I�I@I�m��SzVz��o-���W���s���t�$_}$��H����~�g�g�z�=�ew����{������[_Zb���;����3�y=ʄ�Gz�r����܈�y7+p�$���QB��^th�y�x�,νX ۟Xa1��ZA+U�۴u��GC����)���\��[�żF;o�v�x#nh����2�(�CE4\mB�#v�g��D�춝p%�:�kr�nr�^bɕ;��2��Ԋs�Wn�,q��py�s�c��F����J�Ukj��ͳ��q�����7=QS�5�i��Èݒ�v%�}O~�7�:�aQѮ�7�u��T�A֭oYܕ��&Ci.��=~����O�̏�1h�Z��[d�Y���4;�g4o���~��D�|��O��k��U3��7�1��o���������޽C\R{�wz��`�+���;?W�H��|$�΂�p�锄�5�!�*����
�Ƞy��|�P� $�JC1`uvѮ;��}��$C��W����`���L�}>��9~Ǿ�}z��/��	+�'ge>�á_�ح��EU8�;�^�����}%	!	]��M�m���d�mq���Mn��`멵�f6��5��n)YU@��~��m|��E��7=Y����f�x�7;�1X{պ��������I���Eֹ���Y,����P��@�9b���uN��e�+LWca����>���kY{c.�_W�CQOY���V2���������ӟY9S'f�}����g��{�y*��s�n��t�#�V�3|�[���BJ�H��N���m+��|Ex�z��R���.��[$�$�I�"<6B�o���/�Z�fG�l�_�],>�!y���?5������TY�}�!%$BH���V��MK�v�����yF-��{_N�&���r�*�g�d�z}U�O[�$0b��=���`�C\p�y�����4w�X8_���|~$WL�~�$BH�a���]G6{�w�|G��N[���^���I�P|�_�/U�l��7�OP���w���&vNY�S��.���f$������t�}$@IC�'���3�;7Zݭ�m�,��pj�D�x��U7����<<��1jj�~�{VW��j��^ov����U����Rb�����_mN\k���v��s#(ź����;��}%	%Uq�ܾ��U�y�~� �&����ͻ��my	~��l��7���+>�@�BH�����$�����;�{�q߽}�Z�����������	& ra�{CW�y~���ۂͭ�Y�M`�#��{5���w����\WT��EZ�u����������޿{l�J�ku��܇���7�����I2H��p^�&��<v����~���s�r�*�y8�Cd����,<��l���I�C�����?0d~��%�]wSK�����I$�P����gq����cBu|$����v�K���x��ݮO-�Q���;\5�r��w꫔�m"�s���.�"'_Z����Պ�L��r�*oWM��3s6w<�����}$BH��$��w��w��{q3��	�q�Z�G/{�ͯ�I3�&Iw���~k<�y����٪v�Q���-����`'��쐼��F2�6.�53�w�d�?|{�Ⱦ��dazx���4������i�Ҫ���mG��	+�$_�5���}�S�\w(��Я��V<n{v���N]���^']Ջ��_}_IBH���رX�7��t�мO�f^S^����h�IBH���3���y�|��O $��7�{�:VZ�f�g����o�ߐ��%$BH������������u�g�[�4^�s�f�ӹ	"�O5hgR��.�!�+��+ڡ�(L�X�s�W�v1�K�SW�m'�A3CV
��+�_f������Q�t&#�ZI��Rugp?X��)}v,]���v�s�ױ,,1���1�� �9��nή1�bݮ^:����Jk�$���[D�%�,��+.�9��	�.�Y5�;�k�3��͚v�=�6�A��׆�Z�$�,��.��-$n�Q��׷aؚi��ԫe��Ȑ������E+�!i��G�ݪ��\�l�_��ҕ��"@k;gJR3����_�[<�����}�b������%����@{
�f�&�9"ܣ)�hAK����O_<��(	"� ��]�1Aה׆+���[����W�E��'�f�+k+|�n��k�q��;u�O�r������_t�$�Ƽ�nL�5�}=_?y}$RP�Ij�&�c�'ǧ\�ƭ��ks�^�w/���*I&���wY���j҃辒7��~gq�yN�1^���4��������9�I$�$��w�{7�ԟ@�xb����<�I0I&���{�o=z�����5�!��Mi8�g�'d��f�Nܽ�V(�R�n�7JȺ${���!%$�7ˣ��ZL.�=r{��Bo��.����o�t�IBH��H�7\�U�^|�:c�X�+G��y�`';�
�\}}�1�b�V�x�}7��i�0��ҽۙD>��llU��+s�g�s���+q���� ߫������:��o���I�>���b�I��	�E$_Hz��ٗv�����W%��0p˹�&���<�*H��}%;f��3o۫�|;9	��H���]yz��-��^P��wX��w�1�|=��I$�$����>�t��f�K˕��{�c_l�JK�*9���!�f�v��`,!�N45��]c-���a�#!%vʺ��UEN}��|��'�%y/zx��n��M�C/}���9_s���LE����*�+ Ģ�ݏ�n/��1M�Do�]{췭�|/(>�'S�۞���_!��P�/��W�.Ow؅fҾʏi(��Ke������8��ں�\�]�B���MV�Bu��Mf�U�Ü3�y����!��o#��@ڣ�G���91QDAwm,<7�Z`���V
R���`�A]6�ޛ}fɚ��ۼ=Q�=��m�Y���W3�K��=a��;Ũ��7J��n�UD��'^w�Gu������>��VWM*��6���ל���`��}I_N�rV}�e�l}*�+��1��5H��		%�ۖ��:X�o�&U*�l���[�2�%d*��Ci�f�������l;��:-�7s	Ѝ�v$�a=�Qf൛-�Ȯe��;�U���K3a�.ڥ]��h�MpܵV�)=W�Y��5�л˹�I�=º��z9����T�2�%(9�N�aٗBe�w��5��I�L5�,Х�X�n#*��P��y����qk���N��a��s���M\z�V����wQ9u`!T���B:]�*�C�3q�^���ivVߞn�������
��fm���&d�^�-���y�ܓ�8e�aC^�.A���,:5���m�הR�xEݸ�c�l]�w�h4�zX��-�B�y�/��Y�zGK�y[��Cd�3+��l�ih �sj�n䊶X�73\K�Ly�팋��;�Y�I��ժ��tZ��Ϟ�ٵH��md9;s9b
�RʫiN���N�́�2���oa��s���0Vl2�ޛ��f5�]-��W����[4��]}��m��y)�n𛽮�+��Q'e�4՜���;]��kaTyX�j�w��? I#�~��Q�2 V1��(�#E��$��b���L��j1XؙHI�@jK$�cI�e�"Z5�Ě(���4�I��j0hђ��wY
,�ƍc$Z1X ��3`�,ccc͋sW#fh���d�!�#I�Hl��0�b���A1��)��m�c&�&�d�0���ű��0F�+�ʮj�$T�`ٔ͐Gw"�I��L��#F��E�
a�a�Q�"XѤ��"��膢���g:��+��}�~hl�JI$����l�|�����ƽu��tL��dy淋bܼ\z�곕��n�$�I�?{Ft�Gǯ�Ư�������b��o[��fW��I$N+���r�>t{�gƠ�uƴqq�+-���H�i%�m�.�oY+��t|5��Q��_�_���C����f+���an�L�^v��+}��y3�����PE$_}%}7�lM�7�3Wϫ�8׺{}K��v�����;��%{�[����u���q$BJ�H�����Ro�~嶑ɭ��+z)"�JE���]ټ�!�8�}�� �ܺ�sUq��˷���u���E���>�7�C�l�T��o�O+~�.�ۂ�)�)�,�vR�:Z���.��S�R�^5R�h���=�1=��D�s�K7[�}�rI�I$����OƧ=W��t=�Fͭ��%T�Y&{�=���&I�_�f
ͭ�N靥_�Wj4�^m��1��4q�5�k�XK&�ma��%a�UZ�W�<��)+�$C��]�Q�{ԵVT׽�������|����I��W�����/������u�'��jn߆]�x_��l�}!��o����N���I�M�yz�z��'x��+�M��T�| ��;�8��!%#�5������n�В����r��cT��y-7�k���n<�]�z�5����}$BH�����_m���WS=��'IMON�;jn߆]�x^�l�I_	%g]u�//�%�x�V�c6:�a��/���ۼ��TZ�o�Ͻ*���/��#�<W�j�S���6��-�M֛/,b���wL�|f�Xhv�2��;�.�>�Il�=��R��A-[]����k�5u���m�zsT�rDj��X���4��HJ�#q��t�h���<�Ņ=ngs3)u����*6��sB�/M�H�ۍ�z맄�B��ڎ}����t��]�2xxWj�noB.ᙸp�ŉ�Ѵa�����6������krvƹ�2��lI��e�K�a�Ќ�@�d�q&a8��]�R|���>�۱�q��DV�ue�yd#j�݁xN�t��n���f��k���������:�9ݣ�쥗����"�Gh�E����>�@{�C�$�$^q�t�����=Y��\�������w���x^Po��J��ya��;��*^�;�@I_I��Pp���箵cޡ�u7o�]�z��}�!%	"E����+�v}]�:�.}��WN@fC���;�w\d9����o��Uir���;��}�g�H��/�^����&r����#N�ƾ�nFR�3-�B�;�u�U��RE��#�J�!5���V��UQw1a��v{�vq�����D�X�mvW���l+I�G��{�J� �<>��}C��߰��x\Է���c=)�3������I��t��Q�]c+/�����m���\v^hQ��{ڱm�Z]9�vF����Sꏭ����O=����۶�5,˭��;+*4R�����9����l|���N���ss��߇g��&�<�.�Zi}쯜�)+�'����Nc~��%�r��u|wo��k�$��%I�X�]��v}��o��PG�� ��S�wV�l�>�]���{�}������ťdd�VL�� -�۹��r'�~��1�1B&u���h/��ݑ/��1ͨ��Mp ��_N�����-������ī�+�"@����`�d�;z㧎���H�]���&�8l�Z��`L��;���5����nD�o6��'��2C�pʹ2�}6C	�F�6;��r$�z��������Rڟ�s��������@ �Ƨv��i���].��xf��r��	��G;�'$��Ǆ� �w"A9Ј-�Cn~�mcydy��엏���@����/^[�0pY�� gnT#v������JZZ��Rc���������i)CD^,��zi0ʪ��q��bp��n�:k��\����Ԃ	m�6��3�q�v��H�r$�&܍o6]zSq^ћ\$�ܽ�#f�_�ml���|�T ���-��mkq�8b�E,O�[[�y�[�}�Ϯ����;�����"An ��V��s3�_���S�`��J���4̈́���[��z�3�����L���13�	TG��=p��ȐCn~��h!��r'��x0�و��k���-��o�L@�A|^��~-�$6�@��Uҽk��%p�T E�#�ͅ~�(qÊe׸f���}�� �͑$6�T�
�b����j�~-ꟈ-��m� �ګ��K�n�
�)�Ǐ	��o��7�@��BAۑ?�n@m��;T��atA�꬙��r�;���6��v�r:}�y�߰�g:k� ��ԑW�;s�E��R�T���|u��nُ$�.��'�^{��eG;��&;����/���}킌sT�]��n��p��
������!����)xԂA|�BA�$�U��z^���Ew"z�M�Z%���{�y���B��y�$������PqڡA;�_`LL�svK�Vت�n+	��U����+�6���x]M�7�
9�S ��Ԑs����A-�#=���tM��{�<3`u�(B�bdc6����ٱ_�@6������U"�r�C����!�W����Ç�b/]�������k=�2:VB~x,^RE\su!�"~-� �ۑ=��R{�<}�1
�5%X������A��!E��������ԑ����w��}��/9I��ৱ}�Hh����xf��U�I��Cg&V�Xߍ� A�Cnd�|�m��� �7������n!���9\;�L�^޵��_Z�@z�-� Am��SVW�ly�{
!����<���f���wS��P\�y݅����!�l�5@�ԋy3o�6�vq�5K��U�-d���ϛ���d�RfʻB��ЋE��@�D&B7e�i���5����npv[=�8�6�G	�l�i�]=���ZVU13IZ8I@�ek�bK�E�^=��ئ=����7e�RݴG".K1T� r��V�ɓ�� W��{r;=J�g�Aס0d�y絋�V4L�R�`4{������y]��b���� �	իN<�%��Fɱ���g�ǐ蟯���9�5�Q7��7z��jmF��nq���-��5�Ato3����9��٬��"An�"F�Ţ��|H����������r%�G�=�E���Ck�گ�%����5[��NV��b~;����mH��3v�4M��{�<3x/�\���6܉-�m���C�[;k4z�����r'�s?@�G��W.�[�~��lC�b/�Z�/�I��m��Rm!UB|�p�@Sn~݊ �ۑ��h�좹���4�4�O�q���J#2Y���=w3��"�@6Ղmmo���w���ҝ��;j���P�z'�o ~5\��@��H-� ��w8�b��t�"�	���kG:�� �'��4�7Y��E�k13-���rA��Bٲ'�Cn~��h-ۻ���Y�b3}��|G5{���ҳ�K��y��mY�_�����5��^~��8c��L��+�Q���7A��}�w��/}m�����z0Uvg�V;��l�ΦQJ�*/2�$-W]f_���@�y�'q��%�B�&:���O�"��$�����'���}k�<�@ڐ*7��E�_OŶ�{�ҧ��q|&��-�&n߽ћ���r~��H-� �r$�B�;s�M7W/zD���?7��[�u���"�85׭w���RG��6��Fo�BwQ���������@��[s�q���#$(/�;"@�ٸ9^��	a������?[���m	��י������g6�,s�rr`��M�l��E�q����#"J�`�(�R���RAւ-� Am�7s�7j�ɛ��>��!�n⮆����l�BA�r�B���BH̀�̄F�u��:U�V���1�ϲ+;=�g���ѭ�k�ϭI��-�����}<g1H"� ~;���k��-��x�L�+�m+y���8�1�ZӢ��PW���(D����m�f�����	�$r���A�Mx�{'��������!����;�ܷFnE�	a�����$���{"A�����m��2����ְ��־�Ƴ��Tk�q17aw��f��}\��Dl�z#f.A����~Ύ ��Cm	-��ro�������e�s�w��a��k��)�-�$[k�oُ����N�#"��d�0J���<�p�x�;Y�֕�(�hq�s�n�ܖ���>�>�K/=�%��|ۑ#������˾�oc��7�*�	n��[_6�-���+��K��D���@�R��&���޴��aJ���>�������_�$���;�C̙�{aCnD�s?A�bb�޽uw؍�ߡ��rZ>��]�־�7W͵G�ڒAf�Fѳz���us��P ��Oۛ���Q�Ӈ�Æ��d/��ڡ�5:/g��Fq_�.�����֒�+�ۻ�x��\n�RK4��L\�[U�{�����3)����B�Y5B=��ag�W�p"�f~#u[j~?6Ԃ��mE���a���b>>�R/ǎv�ay]��p���>�BA�Ȓ� Am�!�,n��l߽�	�1��3�a�h.�f)��Zh�Y���b3��h;�c�F�v�p���b~n�xo9�w1w�h��j�+W���A�8���R��Z��|�/yH �ڒH�m	yz\N�ɜ�Jk� ���"~����`��+����H'�+{ 6ۂ�uCۼw즂���N�)�@�ԐKmddV�
3�{lA��o�Y�;��� Mu� xВ�"͹mȑ�k��\���c�$>r'��y��}�|�ߡ��y��/�H#�#~����u5�V�3����E���r$���AW6����U�1�����>������~>��ݑ ���Ŵ,|>�t4�=������5��5�V�͡�9=�δR:�ıf���6BT�/o���uЅ��8JS��7�����k�]k/d�:�hNӼl������s����L{�8�9�Y�n��{XS�{ҷ��޺2�jK��l�E�We^U���Q���UN��1&�[UQ4gD�
����p����w�̲����e]7�ٝ�/��ep�L����CbF��ʔ����ۗ���+�W˱,������_��Y�yߍ�`��n�t��㎤K.�I�q�9$�*���i<j�$:��K�t7٦;���תuN�����ܒ��F�Xmn�g��$��l�t���w=���j�loX;"���Iu��ǖ�.Oj�,�|0�e��M�0%�mZuoz�n���=T7K]��vň��
���⓻�9V겣���N�|���u���*�v��C���感|n�KރEʯ����n�%�Vn����Tja�{3����w*;��n	x�/�$�����Y��5�ʯ�j=��)��<�P���tgL�z�T�Չ�q�%� �u㣗.��ć2��:�����4gi��Emu�	U'3i��T�ño9���[̪�B�t㻵�Wת�H�H��x�9X�F��9i9�eUevous\G8�*�1n�ܣ�PX�ir��rb�Oc=�p�}�aL.�徥�C{n�Mͭ���>�=3ز���q������7m���_�	!��9{{k�vFD�����Xw���E׹�܉��Q0���'}��g���T��ʢ���;��~�w�ֹ��E��Q`�F�b��Xѡh��E2$��1	ED��Ɍ��"�K&4h1PX�F4j@�1�b�BH�d��\��Z1��ō���!�40�5��̨؃j+2�F
������EIFɨ�P`����4P�2Q ��XML��(��b1����;��1�6H���
4H��D���lE���Q���Q��Q&�F��h-%��`���AD@=��)���UU:*�ck�u�(�@5��P����q����sE0���Z.

�4ic��13.ЄN�V7ۍy�gp���噤GZK�P�)n��.jz��[�g���]ηHK�-�7/)�׳AwY�9.λ�ݒ9g���<y�Ƴjx�rH���oK�4%���p�M]����e\���v.�,��P흺�v`��K�U�M�Z�AtT�ƕ�]6��kE���e�qc����[��l��h��)�1t����3IԖ��k����g��,�ŷeMu�!�4�:{8�M>M;^�.�ks{ ��O���3ؕ��Vx�ɻ`k>��na�"昈�A"ì6V�A�3���c[9;@}��ۮ��ы��zwP��,MӛY�ȵs����qgU��f�B���%kf����uڛK��G�@���؛�R.�F�7;K2MiD�X.4���n�����<�Ύ�01v]��wn���TwH�.U�T)�rݚ�#��vl��1�;uN�vT���ƃNw�,�ň�n���}���]`�%c�\v�uy���tz�A���KW8}׫][l<��8�ɣ�Qu�{;�*p�Z���M�q�"�����ɷ\6��{��i�:�VZ��c�J7W�j�>e�*���A[p��^3�]�����s�xd���c7V.{ph��b#l�P�&��ꗓ���hly#q��հ��Rn�	���K��H�Ym��n�\q���nU�:㞵�8���t����f�hF͙m�0���YY�jL"�l!�v�i���-lXqn�zI�FƐ��h�$�m,�d4Y�*�a������m�ŭY��pd|�I�d����V�"�լ-!n׍R1-�7kĐ7n�f�xx.{[��q��J�w=P���v3fu&�0�	�.��kٖ�ym��:P���d/b�\�+�r�y^�<.�xp8���y�h�4�A�Vxn�ܭ���ӣrݹ��u�n|n�^`"�zq�!ٺ�f�����ֽ�Od��66��5�SY�[YCS�9��D,[l��X�he$z�c�Wjͱ�.��%��q��-�4�luŝ˩]�ph��e!16�5ءv����p��ܽc[oq�Mv�.�^+��y�`%��B�X!
n��e�f�X�f�Bʑ�M��[6��KY��úyMP�ͫ�[�����up��������nJ�T��>$O���ߛ_H�� [k����~�޼����\�DD�Fo!c��oaD�V����d��-��!�"A-�{�ۼ�T��J��{�1��~�Awn�g�Ŋ��J'����Ԃۨ mR^������?X��+�@�{�A�����99�Qܡ��k9~>���q5���O� ��������j�ʟs6u�+�.�+ ��7���[j~������G�{D�����8���R���g�C��� �;:D�1�A-���ۑ ��X�$��C{:�;�V]4�sָ����$�Ŷ��mE{r+�Y�^ve�u��}($�12f���A͹豴:Xd�%y��%�Mvi�͋L�����P{-	�"An �܉�xv�}�����R���,�`��$�k�;q��*�@�w��~mm����ʞ�<�P�{%�YrL�Cy^��\(��^v�!���8�&�Z�Mß6w�!}�����
̀���%��o�v���7ܧ�ۍ�{5{��O`�����BH"ۑ%��3~���\��; U����A��"A����u���0Ui����1WTҕ�Z�A/�}#umO��ڒA�&��z�gCC�u��;Ј 6�nn�X�|���=:5�H?d"*�D����,u�?��͵@��m���h [j�쳍׶&!{�1X�^yUlo�mzߢ�{B������A��ȟ�p� �܊G&�����l��~Y�꺠�]"�v�]ػe*�Sv�/iI�F)I��� k13-�����%��/��D��_O͡�Z+���8=uN�z�|��m�]^�7�w����_֤�jHm�6��Σ���a_���cAބרs�q^9]��sG�ѮxH'�!��$��ٴ�9��]+�3P@ϭI�S��"�@6�ښ垙�;��~��^�]w�ݞ334Y�bf���W�r�ei9��Vw��gu.9)�]��tY�q;W�ix�ٷ�[��0P�z�1V[�AT/�n�{�n��@R��|�5\��A�r$�~m��F��Etu���܄�1�����¸7�y��eJ�ָ��w��S�M��m���6���@KnD�q>����=�"Fn�v<��;�<�\5�	�����m��6�_oF^wN�+߃�#�j�Kj㲂yN,k��m���&,mGImewm-��\'��=����]e���4-Ғ-��z�ٵO(�w��Fl��3�ąE=� ���D�s�p�K}<sF�-��r�����Fr��+^j�~w��+��YwD8��r��.U�v��q�A�p�6�X��^�F\Fһγ�շ����5�_�A>�_{�I���E����&=u���A����k�-�#76���o�Uw�)O��}րqR{����Opc��ʨeY�Ƌ���N��^�Ǫ����Y�-�7�*�k�������d�kW�nb��/6)�Ns.�{�����6�A-�~x�H6œ~���{��+�Q��ۙ19T�S�Z�.�}#ڐA ���q����L�'2-I�b#�q��20Xɛ������t��x��u�dxڳ��� M���G=�?�nD�z͌���u/�k��!^����>�~ʨ��]Ȓ;�D�[Aڒ��RG���{u��r/G�R �59�����;�ݒ��<3x O��-�[�g޾����}��$n����A�m���	��E�ڏW�(W7�19T�S�Z�A/�}#��_H-� ��C��|t�W������OǶ>xС��E��t��_��A>�@�Gz�E��nvH�n���$>��~/�G2�b�A��Ȫ�T��=���j�@>ƥ��έ�[���
x^�@�"�BĀ?f ~횇mT��bx�N K�NO���l�ù�DD۱���Cr��+�;o|�hV��kӕ9�&&�o˰b���ܞ��hxy���{���m/\�ct�\��T9뫮D�X���f�h�4jVk�\�k�rnKF��p��<�n!�K:un�i�0�5պ��Rlu�*�i8�D���2m.��6�j �An.�W]t6k��bCK��k�����׸�1�0���;�W��;�e	D�Ա��Y�0!-�u�n�!���B蒵��q:�g)ֲ������l�����b�P�(�,&ơ�cMwLMa�h���k���1���G��\"4#3&~9�!��k��vd�ʦ
�<�"a��9�w��y\���A�G�"�$_ A���`����o��_��d A�n���:�b��^o����g �t�?? �G%PM{��O���my���d�_IX&H�z{ނ���b1����-���/��"�BNd|��D�Q����T�������n�Z���3>�`ǹ�p �si|��r�=_wG@5ܤ���@@���H9��l��g�.�G��*��v�7�׽`��C�8��A$���{>U�����}�?���@�5y���֚�lq3at"ἷ��M�:���o��߯�e���̏�f)�����Ϭoy�&x^�zߥ���P�{ޱ�H�D�łd���E��:��;�k�F�2�z�Y���X/z�Ja�ۏv�$�Kĸ:��]��xE������荒��#貫5�z�"�uyS~�7�G_L�wP@>���{��f}���u��	ͩ�"�s �I�g��U�
6�Y����?I/�+~������.&��'�ӷY_����s�����=@�%��D���/��kg8fߩh ���} �s1[׽�>������{� ~���S��M/c���V�e�&fjhG2��-33�+;to��h{�`<}['V������m���m/����dx���ĺ���g���3�(m�N�r��y,���S�:��z��C��DH�S��>��]�$�B �x�w�7�\q�ch����H�>�����7N��Fw�X�}�˙�?G3/@���s���v�=���^�l���X��xL������ "�ȓ��۱��Qxf�\"�;~�L��"DK�!<j#8����T�◨MTM!oyɦ��{t/�����Q�M��d�;t�w���T�O]��n�1�P�P�S}v��z�e�Z0VKn���ޗk2p7��W���Ȓ��+��Y$2���Hɹp09hI���bm����w��>�k8O��@����.�/j�)���x2=���(i�� �$V"E��¶�VP�j�����)��y�l���1��{��@@�O$H9���{��������=OM�;`�i�gm�����pSӗ�ٲ��v�Z#�L[Lbf[���������e���"32~���Auw_#��}3�0g��;�+��]���'��>� ~�+����@����Q";7��,�&8h>�@����y݆�i��	�ѵ���B ��"IO�������/�'}�`���9�� �s1ƳF��_)�4�,-�O�}��H�s!Fb��$$�+<���j��Ԁ����Ck����L{)��k��%�)?\�0�����iR��2h��G�B�uc'��J
E�2��7�WN����	+Q���AB���+=���r�Vvh�/)#}�\8�B ���~#2>́�31	2.��{�Z��B�#i;k�s7��uuއ�{'����>"Iw��Mچ���%�@��2eJ�PR����p�1n�z�A�ܵ�6q2�����X��Lp �mI��2>G3��������ǧ��!�g�JiT$��qP��4h}�fe�foB9�i�;�û�����N��������[�;��}1�"}�#�%�)��dnf����w)!�_s��3'�Ƞ#1�u&X�r��Y�n/3*��ΐO� A�	"��)��^���컇-o�{��x����YN;��9�C�cӣs���*�{�4���+ӆ=H��K2W�DH6�����SA�߶�꾩��a/s��'v��b�2>�3���ވ���v���xY~�$?C{*�c$�_q�uU�^7W�`�g8z�M[XENХ�HP��Wm���G�[��0��ᨠd)�(JH1L:��eI�헇�N6�[xc[���S�x�W�x��˸�U&��4�Uqtt�{P�h�;�g��Gu#M�z)����hヱ@�܀[`�s�J�B<�o�xou�E����ƴt�J�J0��m���u)@0q��3�v'஺7%��x�B�����76BW�9��E6B
�a���~�1�V;nBm��[i�;d�v����F�=�n^��kE�ѧN�MS�9_��y�#��d"bٯ��Gm�x�
����	Ճ-��kAŝ��>#҂"H��"% A���Js����OVA~�M�wv�l��l���h/��"�! �D?Y׽j%�'Cp+�'�dq�#2#3'�?��*38s�ܥ�����YS���N���j�!����-H���{��O����A��t A�1ۗ���wRǒ�P�y�	��K�׽�7�?\_{܂2R$VA���7�ˤT���"�F>ȥ�C����k��,_ޢ�w����U�32Ą�|����~���߻h<[X%Z�+J�Qam%jC���1R�e>/9��yV#�(��Nr������N=k<|���E>�����%����XA���|��}%��@U���y�=w'�Uq���yi�����ר�5��v�5XCeUNe̚�M�J}aݜՊx�~�Qr�3��"h����� n��ۛ��5=�X���ᷜ/���I3��⟨����Zԁ��`�")�����h�G��,��:�*����*x^�@�lA��H�2���\L��h��>���Oe�'�f~9�!��|��u�*��)����H|Q�n�d�D�Ⱦ�B�JH�|s ӭ�}c��c~�ٹ��MOLvt9��3��	�H��@$_X!�z����������<�F{�ٝ(�g �i��X�|��I�_�;@���v���M���-��b��?_�̄A��b�f��uӴ6�4iKё7��R^mƮ��{"A�!��#3$H'2!��kX�NޫkѠ)���A/z�wT��*n�z'�#�/qI�2S��ל7�}�堎�����$��� �"��<�������c��3�h��RY�Z��h>՗����(��ܨq�w('�0uO��^^�&��\�J�.���2�v��k����YRXý�0\��w�e�Φ�������v�J����o����ע�:d35m]	���ྕ�w�JG���Ɯ#�OkF[*�����ޖ�,��Mv���ej�[c;�v&��f��Ǒ���m��̽{r���۱��U�ǣ�I��L]c��"�oc��簳�uC��KB�^���ś�h��L"�ʾ��<�;V���W�aG6�;C�k�hL˼xv��v���>Z(^���D�F4��D��KЕ�V�U^�y����
�}����T8�q���ֽ��̻��]�K���n��X��ĩƶ87m��-v��e!�M׌iJ�r|�2�^;��n�J�7��17^����R��rg
W�3W;FK��Sy
v{9ڪ��;���4��u-�q�T䪕u�yu�y'�N�<�:�ܶ:fl�c��a�D�eY��Q�Ρ���;[u8�ޱ��]�r��וe�U����jUK*�Ki�sytL�꾕�ݎ�S���CF�vK�b��tٕ�oG+�kB����ٝr��{M}K�r,�
��u��o��t6��M�����j=��G�}��}J�Yq�ܱ�����~V��{��^��lf۞+1ܿ�̻��J��n"48���L��uc�1�꺂ӝ���U�U��k�]�����UP�:w��Koy��bl٦bwU.���X�]0i�u*:��.�3�G�lD5�|��e�{��~�֙��D&2Tb��4_��Em!I��E���ՒŋEE2��%Tc%��ƍLѢ��DlY5�S�p߱�"c&H�M�dѹ�m�BF��ڌ�0�)Qsk�4llX�Z(�)$�MDh �Z���Qy����r�.F1ZѶ�kG9���&
.c�&
���(�����+���F46L���,"�HRs\�������s���Y����࿲R����I��"D��k�fX�}�����-�G��S���}ǩCF���5�#E]bz�!5�������%�)� D���	ǬWtzw�������mKu�1;%~ �z+ ��%|��)�}k��������ƞkn�[],��4����=�F��5�]@[w=�\[5M�)�s����2���#=~�"A̅�f �n�_.��o�I���,f��9�m\�� ���J�Df)��|�)?��� �]��Ϲet�N҈b��8�}O$H9�ׇH�C�E��A݈H�>_f ����������3K��Sr�����m�v+��+� �y�}H����(D�?;0�w;�:�� ����_)_>����������Hp9P���g�Oټ3/�K��v�o/3K+���[:Mc&�y�������YC޽���g���M����u���-�īZC����fߏ���=�9�h�3/H�Yc�N��Y�5��������,��q�QR����"��'2�=if}>�쿣-�8��GSL�2]��ò�T�7tJ�x����5CU�&�]_�^��~ʹ9�-31}#1=�ֻ��~���0�2>�`��ׯj� Gt{��f)f$	9�/��];��ݞ��o!�A}��Gx�g<.�Mpܮ�AʄA�A��'�������Me{M~�oQ3t\s*�̿pk�Ϧ����φ�A�*%�9��l ���%h"J�%�c%�����WS׃ӫ��!�_H�A	���_W��S�#���T�F�m���`[��'����fd�2��]3�+�v�]���컙>ѹHqʄA���'����VϷx�F/��Q�U
�,z��%��M\�fG�
�T�qdWI�c���G.{c{5:��6ns㖜%W*�����3 -�Ƙxj5��\��E�u�!�=oW��>|�h�]����Ӌt��|q�õQ�X��1���Q��W9W�شN�q�j|��b3��6�h��`�3Beԕ�ҖWdф6�4źk�,�Ќ��&8��l�Y�ՙ]u�Y������5�Xme�vd,���0�q9�+�;L��0� U���ܓK�YKWtH�>�/Wms��8��Wb/M<��at�z��[+������ը�u�l�� ��"���Q̳9�L�m�iMQ����Ye��������2>�����ܲ�xn�c�/A�C��ҩ��P���gޤA �K�L��s"��'�E�L�E�<������^�'%�Z�8�^��@�_fF�oni��65�ޓ�(���,3,�s*�!�b"Cd�^�q�=ʢ-���H���p��n�9�-33F��e�eZ5���=+�םK��=� _B �s1H���/5�ނ��K�s�հםQcA��;�/��]�d�2 �N���~�

��9���3s��˾��%�\�8K�R./�����d����/�h�u�ʓ�S�3ͅe��G0�!��ri��|F��2����:);Tu�P\��ѡ̫G1*���r�Z�ԏp�h8vo���"x��Η �V�#�f~#1s!	��;A�ߧ��(�4:{X�鱟�L��3�eb�V#b��LɫUh�*�$ާ� ֟)�VR�w���ܼ3V1��q�����~���@��S�ܼԎ���ľ8 @5��	2�g���ƹ���&�	9���1��"~9�:�T���z����uI�rW<� ���׈#� f)��(J�[�8p���*Ao�XJ�JM��w�.;�5><6�H'."k^m�.��9o
#7��z�9��?�_Nb�a�۩~t��JC�۫�dww��f%�9��<�?�@�3�7�g�r��\�I�"$�LHP�$�
���&a�.��A�ʕ�ԣ��T����G�������@��FfH��� <�����ʹ�PÒ��q�p���<�^/�����S���9�"���;��7'/1g� �hU7�<&�m`���F���.��/P@�̉����"et���p��r�3 /�d A9����}ѣs���}0@v�8�q�J�Mv�=���������n}�zU�u^fn~�U���	,\��3�1�Wry3j޽I����N���_~��;�#��9�q�,L̑"z�1�|��>�Ⱦ韏�1�������Z������/o��2�|�?�� ����P�%2Kd����;ѵ=}�S2N�� �m�ݝg��SS��{{��t� ��"Iw�D2>i������g��H!J���b%0\�K���α��l{v��_)G�m�;���o�����c��A�_Nf.����&G=�p�a=;�6�#��ځ����آ�Ay�$��Rn����?��ow_o_�/�4W7'w�~�Aȟ�(�K�gh8�j�� �3�"H��)�w���~���=6�<��1]�<7���-�?PDI/���FJ_N���yR�����+�Հ�d�矗�}�{�8�L.�;�]"ƈ��cw?]\�1�.�3tp'��{q�g:��y����]��(�Z�=��y����<b�($�S&#ʤ*�ᦺ>@tA��]�d��PK���]�lި߼�v��ޯ,�ta�\�q��Ë�+&H����������?˩�/פ��0F��pnZ����NX�M۰�:;84�[��"�]�~�@��AG?�����UO_OY�蹱�p�}#4[sg�t{��^��8�{���J% A2E�y���/~n<A7����寽�O��8�z����s"���p���p� ���W��d�������u���6e�>�Q_���A�E�4%#�f)#1'ל����z5l��D��D���wW	�4�o���5p�0��?zi�u;�"�g������HA�+��"�K^����Y���|(�ҟe��O�Xq�>\79z�"<��"� �3~��;�j��E��Qg��-��(�F�h�0�[t����#��9y�l�ԑ�su���ː��^`��z��P��3�ev�5��O��g�l��}���Yf \�:1�].)0B��|�HRCӭ�:�8;h06l.�bUĭIC,��Ӊ�n�\�q!cD��v��3�Z�a����9wQZ�ُewQm�@��;V��;KCL��X���a/�Ʋ
�՞#pqg�D���A�Ť���lq���l�u.arg��
�Eɴhe���j�g����f�v���s);��nu��q���9�����Pc�G2	��\���2n 32��3�u��ub�x�����06�'�nnl��V����ޥ�"�J�J�3NLx�{�/�Y�1�U��WWժjO�����D�"H�7�G�,Y��Ӱ��,wڱﾹ�F�ʴ\̷�v�c��J�d���=ˆ�	�@_���d"b�̑"�|���x鉞��}O�/�����1[]ݛ�QT}̸pW^G�<_?l\_G��~�6:;��߆}�oBf\�s(�34j9���=�c����A
޳�{ZW)��:+_} �������m�D�-��J��ٸ.��b�qF�͜C��^�d�ɐ ��a��my����2�)�A���d<����$V��f��s�=*���v"��I��O�|�b�̙�2>�{�w�^��O���x*�hlmV�x[	��,��/V^��W�S۷X����*���d(�G��7�L��O��Èg����_�~=� )�of�Tz����u�p��y|s �̓aGw�
���'�P@�$�/�% A!����]�_~�Z��wZ��R����z�H&�>B��K���d�Eu�虃���O?����:�G�>@�b��|�fx9�O'ˆ�}����z�^���<t"@Dfd�'2�f@@�̦4X�Ԝz3k~�J{ٽ}ݕ++�N
���A<�I��dxL�W��č��(ݥD i�A�O�(�k\ؐr1��.�1��[c^!3<<��}C�o  ?c��2>́�U����G�)^��</_HU�8�g��$��A��'���B�����$J�iVg���v0ǹ���{��S�Z�T-��>���_�S�醪��DI����K��	&�����ݓ��nL�O�KGz��yyzu�uOp��f����厬eR��/��>�ki�~����z����*��L�eP�ܱu����Oyۏ�w^�*��>
�+�.�feD�e0ӂ��>��j� ��V��ȑ|��8�n��t�Ǳ�4��R$ۏ��1�8=7Ǹ��W�|��� ��/�����A�v�����~�@(	"�A�d������[����R6�=�ҟr����p��?lA��OّD��#���UT]��h,]f�.����#6Z��`u�����5Ȓ<�(�$LW�|���p��� Aր���~́[~����H�V��������f٣"~��g ��RR��M�("=�S�C�%��cA]Ӄ�c���>����y� �r��m��c�փ���6������E`�"�J��^?�e�;���J}޺��r�ɏ-�'�~o'���$���X��o�0F������s@t�����2��K��;�=MH#>��Ȝ��הM����b�ݛ�d��Yxo���l�@뷾��5�zN�ǲ��c��*�ɗv"��j�\�̃YQQ��XxFI���A���S�� À������Шt?��{�_ն�|�w���8�y�p9p�$�mFf/�1��{������}�ri�ݮd��v֒����F�͎����_��=�Z#��O��A7mI��dx�s1H�܌��ڙ�t�s�������$��~�G���t"b32g��_"���]p��ܾ�_.����z$]W~0��>��ԀA�#��k"�+����H=@!$�����"�w��Ճ9��̞��'+7��N\ A�@��'㘾̏�_��t�{F;f|���� �|�f)���'�ک��Ը�z8^���q����eD���F�����2�fg�j��gɎ3�>�^�y�>�|ʂ�������
 �_ [k� �굶�[m�m��m�����Z�Z��[n�Z�m��kU���V�km�v֫[o���km��ڭm�䐀BI��$O�@!$���km�kU����Z�m���[o�[U���V�km�U�Z�}�ڬI?�! ���B	'�����)���$�]��9,����������0��,UT!�EHP	  �� U@ P�"E   PP ( �PPHUJ$T�H%E

P
 *�*HR�
��(P�T"H( ��}B�R�
�E�(��Q�*�J��E$��������U$�AIR�*��IUHP �"�{����5A�C� .�I���2 � G  ]J*� 2 ݺ>�IEUy�ȼo�`.�L�l)vuT[�U�U͠u�U�<��ޔ���W��w���6��t���ͥ*�B� �GѲ�	
U%UT���H���S->l0�aꩻ�����U�IUΤ�I*��R��	�B�uK,)NM%JH�H=�=���f��*��R�� �Ψ6w)"��kR�ݝD9 ӻR��	� }��URP�RBT%/��d�R֥w ���*N�;�Y���ʆ�'6P�������� �� 4��<�����J�� d�w`�w u.�P�$�4Qf̀��@�	G�  �*����� �B�O�%j@�&Q(�΁J�R)XU�(9BL�R��$�lUU;�C:D��Na� �x   `w�z��**[�Ac�U��QMۡ@f9i@L�I\�&+�ʊww�;�R�
TA_| |))I��QB�� $} ]�R�� M� �ΊS@�� ���4O���z#��+��P��DU� @� td �U�8�;�8��F��(Yҩ8 dt d��v |      S�A��� � �ɦ` j�ш��$L  �i�a=�L%%4i�&	���i��Ll�!5%5@�  d@$�IHSJ@      $=F�4�Sh#M#5<�M4fA�'����~���~����"=(pu��q�Z��뗩�*�ۜi?�	G�@UA���� "��� lS_�Е	-DUA�kӃ������?Ə�h;S�bl �� �
*���b�Ъ����i40RA@UC�UT�	���U�_��o���}�QT� w�iD�j����( h��yT6�=X~:��k�N4RE�����k�c������"�☷����!&Ks%F,�b�-�wc%/�Kc�ʘ�F#�[�J�Q,� s�,J�W�JR�SSRM�D����V�\Q��LA��ŷX0�D^nb��S[/t�0�	�0NӲY��6Zl�]S����%M�QLL$l\�SE34\��m�Q�taS���ż�S
ܧ!H5&f1J����J�����B�JH�2�[���v�S���G1��k����0̉V*7T�P��J���Z�[�۬bh݇f�e[�g��a�*�] \����"���BgR$̤�lH�tK�Z7N!x�UF=^��B�5��9y���z��.��7J�	soI+],�Xi� ڿ����6_�z��Q9%a	�G1H�Z�qэB�rqһɘ^�t�*^G!�f��*2(3I"ޫ������3'ų���u,U���QG�
A{z����<�j�q�ܩZM\֋�OQ��@��]2��m9B�i���.��c+��2.��dsq䁳��;�;ʗ�QɚU��s��̬��	,�F�I�̧qM@��e�Rt$���]�eD��\�a$�Wn����J�C�nrq�`y)Q�$<�f�L�
=�f&ȩW�N[y�_j��AK��[�y���m2jT¶UL�1�b"������AnՍYF�NJ�&	�u̩X��j��*�q�mf�����c�YA��F�LX�nfL�1ⶅ���0k�T���̄�U�Fp賹h����k$<�a9�Kr��%<�`��I�bD��-d�Sl5S�T7-KY��qm��y)��,E��7f9+�-P�r�(#Sv]�yC���b^t�-B�f�Xyg!����*��c�0Y�735Pk
��ܧzMfE���U��0ڵE�u�xf��9v��۬+wE+��	TeN�eaA��]Ǧ�ǭ�&����Y+�suHܢ��j��P�5��MP�F����4��d�D+�2�����ط7vV�ʚ��Z4Æ��Kb�+G[Y�*����lX+��6VG�"�)F\D���!}Y��f˲��W�f���E�b�"7f�P]�+ܔ�f�rl)��^�������۴�}t��nM{�O��*��k-�G*��62�`'%�%{v2���um�iZ�f�+7`�zj��ӥ�N݅�
M�f�a��\��O�2��ᬪ�2�:�#Am��Ҳw�B�V�r9{(�]]��Q�!�2elҥn-v����3T)չa`�r�YQ㔣N`N�J��-mI��v�9�?�][�����fa��(Ҷ�[Z��M�7l���sj�ڬ�Ɖ��ǺA	���jU��FӼo(�����*����=Ef�&�ʖ�R�y�IL�2�W�N(U�J��.�$�l��ՂG��+[�j��9^���cͣR5I��J�h*�2���E�HnS��{�����4L���=�m̹{p�l�w��%���t˕��w�ULOTtA�{of0F h���XT�hI3R�5{R:h껦��"��7��GNy�Ժp�E��8�r1B�np����B� ���X���5��N[�Ȫ^���i�y�2�bq�wX��$*�LH��w$<M�&���2懸N�c�SYur�b�cF���Z���J/	P��T�yG.��Im�X*;e�Efl9�A�4F�%S�w3�,e(�`��n�I���F%Z)e���bUq�#+F�vd���cE�Tux���Ab��Bn66�m˽����n�J�r�&b�^Z�,ٰFh�V�j����0���n�5��������Z�Oӆ����I���%��5��6�)����Wrz�m�W��'.,�A��61Z��U��)."�Ör�+hē(��~X���O�"P���b�UȐm`H�j�e�'�Xf\����&�Р��y��2mef�̥��Zw�C�NfKO4᠌{�������\aⷀ�XuJ6Dϥ�P��-�xn���M�n���2�g�Ĕ( �E`EM4J �f��ک`���5�zI��Va�Q"�#"ؒ�<DD2!f-�EU����1,*h-M#n�V�6�kIi*�V�v�S[ͻ�ǩe^A���Υ���/H�b(]ѡ��q���0��*�S����r4l �F�D=���U^�̩Q�M2�{M�&(���Dj4�ډb�c	���]�w�EK���� �nԖ&%�6 �&&�T���2 �Ļ���x�C�e:�w�3��,��r��%�i��u��Z0M���V���K��W��mQV�ŕU4"f��8�7�7/D�y`���]Y"*UB!��u��
�ݬ���B{5���˲	dԶ�]5Wu�*	���#7��*:L� �wsuly�g�9G0V3�RX� �j��L�f��iXǗ������h۵�ܽ71
��v6�#�ݛ',n���BL��S]U8�:�؆�\���2Q"��l$Ҹ����$L]����p��f�^��q��f4�'3��I�L�l�Túyd�	8d(`�ץe��&l�e��,ߜ7.�C��c%�(]e�Ɍ�rˆi���V	��$3u\nMŮd�q¢�ڼڥ0��8ۂ\X[��h���n�K5V�췦R$hw-;̳z�(�X^͕kfn͏H�͢���ѥ�\�ɥ&E�1��n�ە0��9�^�I����ə�dNd�#	�-fR!d��9t���fp0� �n�в��M�jE!S\��̷��B%i��2:�-�چS�ll�\����Srr��Hr�]#<�*�Â�D��Q2�IfeL��#�66#���&Ua�������'6�a�t);�Ϥ;VQw��7vM��}����Ʌ+��wVl&��QAD���P�s.���`�U�p���Ź�ysCx��rA����X�-#_���a�	����\�������TH]g�S��ei
�^
�/n��4�(��-B�GT2T�h�f SE��NL�ɒ����j�S����z�:��B��vU�e��N�eڧr^��Mykn隷2;&U75���h��U��j��d�-	��ݜ��Ln#D=�3˕b�r;9,ajZ����"-��흧l[FQ�	���b(�"�ևZXY��mfN���h��&��d���R�̕m�-�5��'e|�m,32ş�U�.E�<F�B��*�-��{��oEcwW�2OfՍ2�*\�Y&�J�Q�4�@.=)T�7[���˙ɔj�ݽ��hkB��*a��D%�j)5M(JQ�!��eoKZ���N��YX^\�I�cB�4�a���"�,�dc~6oJ[.Sv�/7���C[&<J�&c�Ղ���0�����A���j� ��U5N�Ct������ҙ%�F^�n���
�j��)[&�)�&)�5�n��X��$���r�U��pF�-^�.�p�x��u����zotEV�lh/���EXv�wUN-�H*�yQ`��8�X�d��]^ʵd�5��R[˧T�ZXvBV3A6�^�&<��,�#3X�I%��rl��L۠��*?]UD/J0�P#jmū�Ob�5�2:w�]�R��son+M��')�u����`��s�{�"˗z����9hQ
Q�U5x^4��b�%e�3��
�mv���G]��1�PTv`�5���vա�����M
F*!�\�F֛; t��Z0ʾ�uH��x��i���i �Auw��paŅ�{ �z��xbv��a��P�U����T]fZnN��t�ԇ � Ў�7BU��g1�XB�-��mC&�ؗ�ѱ���$�Ŵ4$p��P{wv�R�����	�c���7 �����$�3*+���VMf�������D��d��{�i��.ԩq7~�)\	�ᨔ��{��{z�Q�-L
���V�ö�X�@U*.��L�ld�"�N��1�]@5i\��IXʩH�c�*Û& 0JV�h��&�%��,�*,����T^�	�F�Z�Sr[xٹ`Z�3t�T���Ai^�i�0PyT5I��Zl_:F��z�B6c�iǸVQ��f�]V�AZ�2㺢�-E�+N��n���e��%��R9�r��h۱T wrBܴI�5vɇ)
���AU�]��;��&G��Z	#��gn-�qӻsm��dJ�d�K6ƭ��Z˰����a�b�4i��#3�1�ۖY���	č�WT�JP�a�(͵EB�m:���UA\2���UՆ�q�w-��.Z�����7Z��F����B�n9�3w�VEm�X��7aQըJj���g ��vF��^�[o1C�/��5C��8P�e]��4j���J���U�,V�m��X�[zZ��!�A:)D�[�2ʵ����Z���*��E'�*�SJ�U�q�YilKU�h���3%�U��e����W�-��h�$ć���2༄�U��XL6kp�l����WC*�/T�R��!4p�d^�ʶ*���UI�f���k0ݝ��Z42]-Q��j��n֧MR#Xf�raȑq�YTISd���F��(A
WpBr�Z6��UF�b/j�P��J9n-(;*���P��Ǵ�E�[�䵕f��5V�n��3r i�N�*eP�!؍+w{�*��G�e�m��nf�`eZV��1+az��
����8Aݻu��]óvV�Uڍ^�{�q̶��:9��խT�h=K[���%�)UM�ے�Zѧ3,��B1dTn��Uf�)�駣"�T�M����:�˹�J�t2��)S��ߖ �uzTw��lP�en^��������he5Sr�QT,��k�	�n��wvE^�;a�y��)˸�S%A�:��aR�I�t�a�4�1�ǥ뽩V:�H����j�T�x�����k3N&����\�n�CB�faՀ�v��4��/N��a^��:�@�6[�F-ݢ����w,�4(m�]Qk,ݫp��P�0����w+eaP{�U�Z����n]��ӷY�o2=�\u0ȁ�4d?V�wm�-�������SHՃJo[���y���m�j^iަ�]Ew��J��$�e��.�EV���cǖ���ʤcrSP��A�
�J�ᄅ)!�Q�8�ZB/Z���W1��3A׀�w.�v���RY��¾�ҩ�#e�ѕ�Kvl��k(��6V�b��sMe�tm�(h���e�F�*���"��͋B���	�T#KY�����օV��$��J��e^]D�A��[�6K��-u2��nѐ8Rww�em�n�&V�X�V+�o1>�U��K����,еL�f]�j���kcpI�8�VmH���Q��har/�e=F�;ћ�a2enޣ˘PB1[0f�9����A2XV�+ڽNR
������Z�Y���O7zuf��Y�"n1��XC�z*+0m�J�l�2a�Kau0ChAUKv�5V�����jQ�����l"�+a8�U��ҏ��p��n,��W�T�t<��4Js);-L���oS[��"�ÈKV��rSr��f�ϴn��㤞AcU��(6��{���b�^��?+.�2��n;�6贆���
���z.�z;���<#��w`�*VR�d�O}]xzb4�c��֌4��g�,�uZB��ݯ�B�Ғ�&�-�E���ӧj3
	����'�]�u��YVطX�]��n+��)���v�+gF-[m�(us��a5W�rU��yi���-T���ʶ�3����X޶t
ՂƇ3&%W|3��w�ZuY�s�ȳ��o3p=hjߦf�@�\�YyI�ۑ[Ԏ�an���C��wB�w��^B��U�rdIm
�����Me�(�wh���9��X,�K	�{�+%��H���,�{w�a�Vh���\�v�[LZ���R����Z���Q�3F��$�s{ڟ����5���C^��yaGI����w��=U'�룞Y��VrY�:��
��(2*2V�mm�m���6�(�V�j�Tmk�Q�%Z-�ѵ�j�F�jŵ�mm��Ѵm���ֱV�mh�b�X���*��+Q��ض��-Tkm�Vѵ��h�b���mV��lj�������U�T[lj���Q��[U�ƬUTkmE�E��m�����+j�Z�m�F�Q����+m�mk��[cUc[lm�kU�Zѵ�Fѭlm�FՊ�j�b��6�����"��Ȉ$��(����>�G���������	�ނ
�5��<_|* �>�{�E�A�ʢ�?x:@P~���o�?���u7~�,�?������]S�NgqǛR�M^���J&5[�*���}w���$����ϱ=��j�*��P�О�����H�/�P�����J�����4�V���ݮ����U0eu1U��e�#/g���C�8�+=ti"Ůw�a��b�by�G	�v.K��o]�lJ�M��Y29lP�ӷ��)1�v��a�hE�{�]�M�.��!��QQ��P(�Dz���
�WIRU��o\�%Dd�0�yT�"�fcwT�/(��T�s֞卭�e\\^"�j�Ҥ2+e��n��j�+����jH�j�U��y��ȶY��+�f�����ыT�(T�������iYEY��C tr�"��9U�1F��Yf��sH��%q����5�R�t���*�B�;�jjg5a��Wm�%��ӓe�Em̖D&Wˮ�WU�;%�ۚ�A��ݎ��{YԮ�Z�P�m@��K*NR�Q��FMsHe�G6$*�%W/ ��\H�B�)���C��+:�Q�X�(�Q���� ͺz�������V�qt�d���UWO�(�݋��iɊ�<F��G,�����m�<:��+5>���\���XiuS{����3�����y0+Qut���շ�.�iK;�5�*���*rq�C���������I8}ј�����D<r̈���ذ*j8��3Zr� F��yjhA�ԩ2�T@(P�,Vq�c��A
 ��4��(�n,�9;���꘩�s3�J�GTݰ��9^i��J��*�.��F�;͐��ʦb J͈�&i�T����Th_28A�0Q���bX��uf�I��;�R���V�������/�Q	쫶�Bw�̌AD����C�{�)L��|#�WҙY6:�ZϷ.<X�UЁ��Z�.���d\��'m]%}'e���\R9�v=����.�Q��ҵun:���K��ʥw0���{�Vn�f�����p؆�`�l�+U.�^���u��N
��*be20ы�T�$�f�C,�����YG#��T-��s0������.XhԠUf�Z8����0 EV�wM8��&b�P��΍��E���.�IՅ�9V(f�t�<Ub�M���Ѽ#�A��U؏���Mr%0YR1�R����e�0P���(�f���.�G��(�P��j����6,��0S���ka݈��)�S�װЕ���4��	���Un�!amF�"��l*Z�����3�eڜaeP��[�^M��|�ؘ�
?�pY�
��U���
{P�tK�t:@�!£*�ҫ˛�&]͡vATj��j�����i���ҍx�T`�B�Ke�V�rr���n���=�ٗ+h���l2���.]ִ�%Q���\�{�S$y�vee�	�ʙ�3��bȃe4&.c�v�Cj��toQ̢��V�齍a��Va�3rK�`?6j��(��5�m^y�#�GUB^�ܶ�x"{oJ�Y7z��z�,�h�$D���)L��Mͺ�/EЙ�4�ayT�2���;s4��UJ��z�Rv"ٚ~��J,�ۚ��*��|��d�<�12ý�Fb؉�}$�N"�Q��mV��9ѭ�,��V�[��\�6��6Yq�%ݓj�u�{�y@������ќ���ʲ;�o	��0�;Gln	XC���5�2]�-�|jʼ�y�sK�r1�XG)`�1�J��XR̓
ʙ���bb�
foQ)V�c
JʣTJةj&L�\�7}�r�Ф[g���#YB��%�fm	Kv�u����Y�ɜ�lU*݋J�#+,���CH�ni{x�ewmUw1[Y;
EʹYJ�cW�CT��V��@��z��U@�GU��P�o��K��&2Tɻ�3�
�U�=Ez�D)�g"h_\yr���i��θ�q�Z�w���"6\ˆ������C�Yˢ����;��f>�[{ƚ��r�2��Wc�R�Q/�^�&^��i�G5��r%��H�L�3��F�0j�w���82J���3�m(��X�L�񳎲�]���US��	�))yd�3��{[��ٰju�dFt�qk?wnХS�`�]�1�bth���k�}��H��/%�3%,/0egfEK2�lzީ��'���L;؅�K5����6�^�����Qu�q�ʻUN๗���Q6��M���wFPP�K�Հ康���X�´���\���׼��*B��9��u�X��b�j��L&���-I1���gK.h7���F�u�7<KRʱ��6���f���]
5Q�jC	&]���q���S�"�w|kz�:�cK�.�RK �r�ds80��9VM^�w��lc˃J���n��<Ѭk"�t��g�2��eZX�ͫf؟e1u�!�:��q�kK.��ᕕ�h`�p�@����P=R<Zܴo�1�jlP;P����6e<G推$!]��uup�Z̫V�
ˉ�',���2�^��>�79�[�Ҳ|~���5�X��#3�_b��D����餆r+%jF*��$����p�#�b�yB�m�,.�j�%��xUv�CF�edZeY��#v�7eSM�k]@���t���jɺ�T㪴�L]}چ��q�c��s�M���cv�n,�]G��J�&�X�3�A�*�5�+MLA�!�y�}Hs�J�`|]*��K�Bm�x�p��'+FȳPL�)`vP*��7_Gq˸%<O4�s��e��/�iQ��X�.�Ъ�e�jd��N�8K��8P!F�M��R��<��.��5W�uX6T�Tl;%R�w���uU1�\ov5Q�0;��C�����/hl��9
m���:������aH;��J,���;-K�*�L[j�]��EJ��׶��y�,���������T���tɁ��ڹ���@���|�ͼ�ܱ�;U�Ym�n�eV�
/�ɹ��%Lk�u����76�oV�u�WST�eE�����e,ʼr�JX�I2�Q2�S�
ɡ)�=f��t҄�t]m� ��Һ�AU�ύ���|� �PŴ��7�!!�i��S��%\��r��|�l�D(iY%�̼���t�$7*�6�R��:aX���F%YW��AUm�1��D����B���G)�{���i��1IϻK��E���t�w;J�c7/)kWetwi����g$��ڭ"VYrd�-Y��l��ue֕�������k2�T�x����B,�n��ͺ��v��nmаҾ��%Uz�Ij��ma�y�ή�ى����U,�]}������H�t��ub]c�lv�<.�v���f.�C%}�LfUSט!T	�v���8p=D#J�S��8�!e��a�;ϩ+�Q�:6�aU)0 �n���u�h���hͻ8ʄN�0��T�N�|���^�Se�=D�%0�6�6E�SD*-�вuf�`�0,Դ/,�˥�sMs�&��9'��Q��qݾ�1#]��`����UCF���I�D�J���hQ�:�>�墁�f�f�/Fާ1�����]ۉ�V�s*��i���gv|�,"ŕVo��e�Y9O&��L�5]"�bJ�Ʉ�@���̠�yo��Qv����7��-n�˓'2�7K=�c��V
�6��(�N��$՗H�q��v���f�4ʔ��M�"ٵk*�9_Z<N�tW�,�}�XWM��ԡJٖ��a�6�M-���ph�j.O��fl�8W���x!��[��a�\�ɓKLѕ�o��	�+(�����y��;�b5_}c���}Fk�R�sj�wC~�E�ˢ���ӂ�I�#�sT��6��Q:��B�L����i�g9�����ъ���$�@�e��g)]��P�Tj��Uc����8��k�5z9�Q����R�3N]R��Q�R��u��Y�Ѝ=t��!�w:d[�eȗs�S���W��F(i��d��LU��e<��P�ZX��v(]��7du���Il�"�Z^P�h1��t���J����oT�2�]dC���{]N)��*TRfڴ�]a�n2�����VM)��I��+1AF�ڦn���&#�<8WF�ͬ�)���6���e����ϻ�6�i��s��OU�J�p$V�g91Om4�q��5[��K �Y4�[�+"o,�VK1F�pʀ��j��=n��2�I��O�z8vqҁ��_pr�������Dg+��2�\��W0�������r�V�6�¼��p���P�2;���٧����G&x�a��WF�ӗzv�{�c>g�	��dF�L(���:Kvy;�����F֮�Nм�V�������"�x*qǠ�͜�MЇUua	K��b�S*WJ\;l(r�X`�����J˽����n�`+�Z�!N�]ΫLmK�'^X�J�+�6�b����S�sO�j�ѹ�����ܤ�y�gmu��q6�Y�XV:����44�˻6��
�	�[jU�YF��)�E�X���aȳOhFM�2�I�T�*&=w��"�u�t��9������
�3��l�E�#j�7t�����	2�Wjj-��l&�S�Lʫ�Ќ��wi^*�с�MbZ���qQ}��f��*�ل;Hٓ#YUܷ-9s�d�����ԫ`lU�Q�52Qb�pbŞ'"W���Tw���ḙڅiˇ��6{rd��.�;S5�x
���7->���u�:go#����!��{Î�sHl���
�t�1W2��2]�͌]ryB�gY�A��������4kb�n��8��p�c��M�s��#���l6�5D�O+���!�λ�2���S��Sx�"Gm�]�$6g�(�,n�5#��e��Ҭ�:Ne۾u��B�x t>�x�ۍZ������w1i�������[�1,�ySr����hl��:UT��
U�rUĽ�=ψ�v����-q�����)-�W�+��0j��y����f·����fo\��l'^�W��SO���_-<�Yj`!�&%쀧�8L�Z�i���\A�.<��W݃c�+tc�$��U�-�2ӣ���Rx`w�i�"Յ����v�J�pŗ�T��+eu�_H���TY�DXbԆػU-���v7�VseT�-|m^vf��N�k�f`(nM��0+�З�v��X+2<	u�OY��v��L&�3gƝ��V�[�)�R�F�����$u]��s�2�Q���Yd�T�ǈC�l9W���[(�p�,�i)�ܳC�fi�ո1q���U�ߩ#D����:{.��;�ٽ4�m$Vdյ��vJ��cw���o��&e'W�gA��/�VY�"ymT����_f�U@����`�����i�W�I�B�J	USu��L9,���Q�U:$�a�m��a0�!�j_��ن�KR,e�YP���0\���˅�ߖ]rK�r�`S�_]����AAcH�T�0nd�B�N)Q�	���i��o*����R�B�z�P�2u��X��I���{�Y����*/&J�^<`��e-C���공��\�0)K.镕R�Ъ�mWi�����x�,s�Ɇ�p�.�63&C{/��v��9kֱ�s%i��%ƶ���c+����5� '�����\��g��+��!���k*�V6�7��o]����[V��L�KeZ��Ѫ۶6fJ[Es��9�v��f��/�
�V���R�)]�.4�l��b.����T5Z�M�/�;e$��P[*�KJ����(e売�^7��:�Pc�B�����'ض�V�"ɺ��Ǣ�Ղ���	��E�`|��r�F�ƭ�k@�G	�T���ע�f��w3.Ŋ1���5�qe�VN����YUƾ�W �Z�N�Õ�8rX�Gj���e���5u�[�v\I�9����b����2��,�\d-�z.�$��t:���uN�mkWi���bdL�4G����(�H����.I�$R��'��|��f��������c�fuB#��cHV0�]������ۛ�er�1-&�cK��l� ��rMN�hmi'b&*� �k���8��-4ki](6�&4n�\��i���n,�c�l-�fCd�6p`�T�&���2��gJ̀(�,-�)�7o0�tfTi�\a�rh�+�1+\��.4#tql�h�.4Q֭��RY�f�*��S�����,V��%�6˷Ja��T�k���������pu2!e���2��6[֐�C���Ֆ$yYlSmL��
�ys�Ě�6u�X#����7fVX�lѽj��c�ku-�M��gPq�jB���J�7��*��t4�6M%;8�j[�k+�$-pV��4A`�2]A��m����̬Vh5���c+�v�f��fP�(]j���0��׵�X[p�)Xv��f��)q6(��M��]buR�˘�m,�f2��9�Z�pe��u�H�J�L��@�h�.�l������EM�PD�5��;U�Z�͐Ie"�5�ÖQX3h�K�m1�d��@֑
&�X�v�����X�C�G����u5wV��g�u�l3v�j�ы@���Rj�eS
 Wml�mB�t��iX�����n6�%U�g�Wy,<��aJ�.WWl�$���sh:c�
-�Rb@,@NCB�-M�̥�GK��%���,��F�K{r��3��ܓ���,J�ڮ
<@�F�le�St%qA1��[-D�m�-����W�ךCJ��B��"M��X�Sr8�͗�A�(Śi��u�m���#<�;^�1��[L.LTIM�J���ɘ�6�K�M�V�WM4�a��{B,�D5��.� %3��a�M�[��`�nڶ��X�\7�#L�c�Ihq6[�1ī��0��Q��WkY�n���J�&Օ5��I�&��V��h�4ԗLr�4��c�Ԍh�`�s��aCe�Q�{;Ul�ڴk[���;
F�sU�[,.v��؃��������q��+J�@�66�ԨWYi�n+��i�\�B��P�ְZlmp�0��4-��Z�9�aG����&ֻ%�š�mΡE2���0���+H�-���,� �����`���:�ƺ��0`�qF�VY��cr+��2dCDƭ��5��B�JA�h3j���tx��i�^�hZ\0J<�ub3%�X7T��S��e�yO+ڮ�Ќ�)`D��;0��Z*@���6�������&��hHCF[),B�LT��$��g8f� �S[�,c����Jf�cX�A�-�M�\ҶԺ��	��ۅ&14z���РlF2��X:,v���M)h�֕�%���	k�kڅ�,FԨ����ͼ���G6��;+ճSj����U�����j�V�ۓh�P��F�KB0�o[4��mͽ����cX��#@5�ms� ܲ�6ȁ6��+4@�T�teC0����ѥ��!��c�Ս�s��dc����Xn�6(-qH�/]���Z�Ũ��8��kT6q]NEq��͠�KA��j0�A�,����zõN��-E�й\`ņ!)l\�MCg�G$�61s�<1ǆ�.���1[[����Ķ���R�f[j��%�M�M�vQ��jh�"�a�ְ�5�P�1a�3K���fQ���^������ g��m��b�6�ع��66
��\�ؼM2���݈V�0�`	Ju���[J;`v�q�H�Qؕ�t�j�hڵb$�t��
�+�H��e�og8��jDC3jhV8Yq�a����d٢Xi�v��+���A�$��uنu�1Z��SK+.y�wr1�uc -�f@�v����]EI�iN�H[�`�f�e�s(�kve��y�f��xgc3[U�5�通��2˅T׋+v�ye�n&��D��suj(�ۉIu� ��
�r\V�t�7a�
��Էh�KŴ�����a%Mֲ��ۂ8�P��YD�Lݷ	Nd���^xn�	-�v
&�C�v��<��S87-��nʲҍ�T�^-���f5��f�2jI����%�*ke�h��U�5]�$K��a0%44q.  �\[l�CQ.��QՖZ2�VתL,3-�T�"��%ʅ�f�Z���]hgAΎ)	���A̺:Yvև��YL�3MmB��X�Ga6"l�ћm��.̱�]]5��4If���6�RWL,�.�JAuԴ����dBYn��] Ѷ�gb�LZ��+6��E	�H9ĺ]i���e��*�a��m)*�k Zq�#b�SfW8�▙���.�t������iz�-5nL�m���Ĵ�֨��؛n2�[��k��F��ۮ��2�v��f`�����%tcv4m��D!x.S5��b���n����a�A�	��,+ĕ���t"5�f�hٺ��-K�V�ZmDۨ�0������s�M3Xh�xFT���7*��u&����ƈ�Re�.�Z�� �"Yea[��q�eH)K�"[.�1t���j�
�j��YiA,��ض[�Bh�)Mj;Z�O1��֣�����ѓf�����9U��9Q̹�X���:j�J���P�)-c��ְ����)Qt(!-�Z�0��Y
��#ť�Z[(Z�ŋ[v5Bƈ:�(#�hX��FC�Yb�h��ՎL����M[�����&�Y��ѻi
۪�1�-r�����*�H��KvĬYFR�n�mkL�0�38����0�62fЪ�b#�K�;jlS;h�&H��XYh(�7T X�E�*�D`l|\_�X��S8��*�ͮy.�%���!ͤ�C<R��6`�Kt�1j��1�Ǆ�H���]��%S����B�h�mŘ�Ք�-Í�95�u��q����9��0����iRb�ìn�l������Е�8f
u*Dx���#6Й[����e3e	������Z��.0��	�P�w)d3����
�3:)S9m�]c�I6��)y\�kj´�-`Ж�,�m��7I��9�JU��RǮ�n#��B嶌F��c,���;b��֦�.�ĳQ�5��ռQ(��ͩ�#F(ع�M͸�z5�*1֭���j~j��)n�:..e�����m;��5��@(�v���LĉV+W\j������Ѝ�
A����0�V��-Mu�Q)y�YP�f�n,H�"�$�ؤ�c�4-t֢��:�����C�H�VlA����ZG)J�W$t5���kR�֐��^�U�X(F���ڎ�`\YZ������S�6Q��t�b���J�"W%��[Ye�j�:T�tQK��Mlf��B�B����WZ������0�	�x���HJ���@���[3Ly6��7GJc�� 
�f�^h[��n7^���"@i��#���KC&&�5�:��ցÛu�
�J�`gR]��-�-�XͤeBR�ILJX�d��ʶYQ�B�5��	�
7ʻ#�r�RT�bK+	0h;]���F@@�к��x�T1s��rX;Tk�5p�#)s�Ko\��Z�jAKlK5�k�1�:!�.�*Q���,�3nL�78��B�O"D��]��i���X��t�i��3s�e� �5�%1�����S�Ͱ�%���2k7bU�h+��b�g	��R�)3v���ZĻ��f&2����L�v��v�-+2]v��,Ch8��3���[-�H�{ ��t��p*�һ�hAs/l6����уm\G0�`�KA�ˆ�G%�H�e�<�A�;������j�m�ݎy)�]2�n�8Gj�S1u�+�a6Jm͹��Dm����X)|i�M�>x�Ri�V���bYsW]ܲ���`���"ZXW��
W��4��0=�b�v��ʥ���-�4���a*-���Xo<f-�3� �-ejV�Eh��M3f�=��=Y�0�KF�]kq�5��˦�hE���ʢ�c��ƛT�]��cT�)r�mp�b�l\X:fꂏ1��9�Ƭ��fC�hh��̶����V�n�"��1U�t���L��Aͅη*���,Ius`���W[��b�UJ��pf
�2��ʪ��j��U�UUUUUUUUUUUUUUUUUUUUUUA-<�#[���6�A�8�f��Jء���aݡժg ��F�.nC=�uL���e�#Ԇ��U��6�m��fp�xr��a��`Sמy|�*�rh�b�2LBl@��ꮦ�a�\CL@�v�֠����.B����w��B��C���~<�ni�m�����w62%�*6����5�5�wu��>.�+���ᯊ�)d,���C�$&�)��7�~{ו���oF����w�
,{�	�۴y��mr���5��o�_�u^y^7�O,h����ۛ�:��W�pT�[�����n�y\\�u�_=�X��v�wv]�^ncϦ�ב8�vA��ӻװ��>{=ϼ�f��3l�L���rWhZ�l5u�\L�Z۫�[J�)IKN�FZ�	]h°�hffZkfլ#(J�\"�ut���2F��-6�.��"��ŗ$h�U-����We.�uAT���˝�j, ��#���p���dͮ�-6�LB�a��6Jf�a�	d�T�����,6"X�l҂R��4���q,�ZP���%fy�my����X��VZ6LF���S)f��Kh����Q�ݠX�؊vչ,�f�c�0��jV���䕊�0�
Y��T����0d��E��1]p��5WL�	��j�!qa�4ҋ�]�v��$ť6�2S�V��n!�qU&�L��13i(Re�iR� L��R�M��,f1�Ii3Z���M˶�Ҋ�Kr�30z����j�Wk�75�M��	V�f�F7ZZ�w�F�- �i෭�F4C+t���u��-�����h��k�k�n��[	^JT�)�6�*��Tݩe�;�m�a3M�nZ�t�[-]���F3[-��
$��\�]��`�[)Z���혱)hT5I��QA���].ѥf��� �bib�C �i�e�ceVQI��h����U��(J��e�f���9 Ls-5K�`ɨ��ur0�i� ˣo�N��얰�-��Śp�ne�èE������)����P�[\�&f��9*�i�D��G+Z�����l؍����i-�G1��o��%e�,,�!*��&Cf�W:[�F�@4�������X�%����1[�cьlh�2��ѥ5���ҮQQ�]U��UUUWM�2�^n��+ݶ�Ҫ�٠,�����@�j��֤�#x���HQ��#,(Pyk�e�u�m������T��se"�l��%�[T�h���Um ��b�@h�mZ���D��ŤUh�mc�62�%D$[KJ�(5K,�RTF�m%xDh��S7ϐ��5�o��8-֭��]uM �3Z�aK)Y�
fe_�ZK���nj���@�f)I;W;�\��`�"���W�
�|G
x����A��m̂[��Eq`�utϻ`���y/:��A=ܤs�@��o1+��J�R|��9��"An<��r�Fg��g�^�ֹ��^�(p<�}�m�7�p���#z��A�5x��h t A�m�7�&m�tc�7#ys #�˅��Z��=p��"r�p�!�6�8N��0����ʓ��n��.���4-� ��L����"�vcr�U-e�Ԓ���r������lS*�=[=z�7P�p�n�2w�>��1U+ҧ�L-����r҆A�4\�>!��� ڒ>\���\��
��7��g�<7)�?53F�{R��8�����}�^���G>�������_��C7���2$�B �Ƨ'/;���3qb	���A�s�%������輀ȧs �q���ȟ7�okt�Z�z��M�]�mG/�zy��p��Ԃ@ uX#:2,p�Bb{�(���q�m(!=�ޮɊ�^���y��Č<�m����	���p�ڟ"rnX3�JX��T2��&oN���7!Ǫ�qyȒ�yx6���ׯ�&}E�]�7M��ȱ�*�1+�5ѵJ���n�&HS&&eL�=9>��9�"s>!���z�N��-��9�%���9�OZ^���t"	m�7ap���9�9��q��'�	{��1U+�3�A��@�A��]��/<���Ǒ�ק��-�m\�Z�E8��Y�����N�s�.��ێ��/:�h�*s1�oJ�*˱�j%�k-��؝��%�&g��탾��S�]��z�mm��T�J�qu�;����6����ӹ4�.j8��T�s;YhI�� �l#�Ƥ��/� Cmy��ggV��p��8��{��ez&{�9�圂 ���|[B^�>��O_ig܌��!fq�m��Y�:6:8�qF1��Bi��*fGx�SRFl[�|�R�YuOg���Ն�`����[qZT �wdI�nۙ�q�v�]X�k��#���w �j��k�ܚw�K�A7ڤ�����n��-�������%�Cn|�z�m����vv���L�D�{aG4�m�7�p���t+o�z�]�>�i���/��xv��X���x�����T��Sͭ5:Bc�73=Ӕ5��,2e����Kb-��6v,�J�9u.��(9���ө���n�q�;PD6В�"1�D6�3c$��2�Cާ�N��mG7ڤ�-�>m��1"�j1?M�BaLD�31�h͠ZbW2�U�Bg^�M����|��l�~�ǻ"Kq��(H����d�L�D�H�v��tn�ST�@"r��"||��q���:-��[/����vꕆ�/�nxs-���dF�B|[�26am��@��2	݄-��mȟ72u����n��;�%Ïq�� �9��p�Ŷ�݄:p�u�P�T��"���[�Am
V�"�ML�J��|{ax�]q��P�Bj������mI�E�ԏw���0����7;#�����'2�"|[�A�$��9�Fvs`��M�؉/�J�ӞU�XhJ�\R��D���-&�رJ=����2�T��u�)IT%*)@�ĊL�\V��1z��3dK|V�ڡ��D&0�]�R�2�kT���1���a4�ˑ"�6�jMM	D+���֔2 K2[1�:��u��ٺUj�ɦ���C[MH-R]\n�ꕀ���\`1���if��a����r&��B�`�B��f3���r�]���r�)��V��5L:�f��-c��*CT���ggf_=3�~�Az�!�3���B�.�uU��%Î غrȕ˓ �܂��"�Rm Kp�q��1Y1�q˄A��
��|��SS+ҧ����m��Ť^?]G�!�A����_�p��m\�w��p+gNg����|,P���>n,��ۙ*�cZ��Q�pc��mwy�Gz��j���s���ܫTd��%�yx�r�H� A�nD��xͨ�m�#�����֪�cҧ���/G4���4�_��zߍ �)�o��cv�B1���&���4�ib :��B�
feS��	�jA`"�"	�ԡY�ok�yd6�|�1�yۗ0�� �B@6�A-Ǳ�t:TzE��+}b-6ں�)R��d&|�^�p'r�1ժ���:��n�0c�\���M=�5�yv�~�bP�L�>�!U�ɾ���w�K�}��H<�^-�z^Ҏ�_)�����$��ǔ�f�*�85]�[jjf=+�� A�!�>�A��Fҝ��{���A�Z�6�Ԅ+5��t��M�� À�>5��yw҄�����	n ���/sv�}#z��p(;���rkx���>9ܤ���� A-��Fލ[�c��b%�2"`Bj�Ҩ-
��S[��8���"�ʪ��g���,��=���m�1}�z.jTz&zExn����+���6� ����^ع�z*�a�܅�/5HB��r�
ܷ!�^̀�yȟ�[ِDw ���;��A۟O��g��[�I��F!;А蘨3�5D��F�Qj��a�lIk�T�\Q+P�ڀ�=��Yʷ���;�P�?,��Κ.@���'b��v�O4nD6��!9�1x2������� �l��,[AUP����[��J�D�	��z��#�nI�C|C̙��E�D[jH-�7d��3���kÎ�Lv��n0C� NdA|�H-� ����,,���h���W�eb�[JMGk�ec(���\`ѕ���u�J���rW�c��CngŴ��ϲ/*��;�$vAʮ��ҰA�s�	m�6���Y����b��.��Az��G�Ӽ�T��L�� G8ۧ�"NnU�S���z�[Ax�����KF�F��#I�z:֦�>^yC�"Kq���~�V��H��7�#��X��Qy;�u�����H�L���Wd�o;4Ă	p�54���x��u�f+�u�{r�R�S3�;9�>�ᯥ���/\ӗ�������X�O-��p,��r'ŸQ�1�vL]pcZ�1��;���G�g�^���"r'�6�8���(�PsD!A�52v����@v��;� �
�m�[X=qv���=K	����A�"�mJ��wL�ũ���5�ʤ&D���A��ly���[�E�Ņ���XmT�-m�e��������H#9[��	�����|GZ^퀼Amȟ�ɴ6yap��MQ��/4��71�<$���mϧ�6��DE�ed�ت[��)��l A-�}�k��V�q���ӳn��ݍ/! A���m������m��b��'�O{ ���m�^ff�; ����[�k��!v�!Zn�b%��u�L��WcDi����dͷ�M��2ĻF�6%t+1�.�T��a���^�8����;��jȍ�u6v��S���Cu��2���@u������+��ЄW:��0llt���1�\a�j�2졍M-r$]�M�sm���jf�ڵ#�k����3a(�a6J�h`����;���ݳcr�P��#cc�a#7kyK&�FW)��R�a2iR�"�ܤ66L�;rZ�{7�翟Ann]���4+BǮ� ѳ9ib��#kj�&fT�;�z�"��q���SD�����	��x`3�9����>?O�H C�3���KmH s�wvГ[ ^�~T�k�]���� N�A�������:nH�\�#�מŐCh��||��Qʆ�]B��쬻��v{��Rh/�	m�!��"���m!�Z܍T�QȐsax�ATш�g8w
���B�;��sk)��{��arD���n ������y���0s�O�n9�7ݑ�c\`���C愖�[C��O�67^&p�g
�M3)�[�iR�QMm5f) �ə�2�Gt��@���k�A���쬻��`�8�C����2��M%^ ��ޏ [k���"7C�T�+���������X6\ž�����Yؔhޖ&5�%��g2nz/549�v䝹zt]����X�GW]�V��VB �B�K��/�FT@�(p;��<�@��}T�>���k�o^=����7����AS55���}n:65�}��� ��`���ۑ#>���>�A��'�Ǫ��e�=e�� ���>#b��vS��3��R�E�6����ħ���'��
���
zA=���h݉�m�bk�����<�:�s=��ǴE�f�3��r��]tw0���\�S3)��A��>�`�E����C�>~><z|,i���QIáB�w"Ot"hn�[�DC�����H�T�����#uW�q�Y������yO���nK�6h���^��	������l3(�������:��z�~��_�&l�'p<��:A�2��T����B��G�vN�������
�ㆲ�v�s�z�u�*�sfi�n➝�v��jӊ���9z��ő����NF(�v��<�HYa=אP��G���Q�����9�J�	������9%^p\ݝ����8j��z�-\��jH�����U�鐍�R pL(UO;=�FVl��ӷ�e��s&�nc7q��nk��y#�Lv����w�ۺ�@�8�Bc5wrhy�-��>��0����u�C%���FU���c��<�2���\a^�%X3�V�5\�3�U�K��C;r�9���d5�ni�S�U����R�G����x"hhF�9���d�8��=��ڼ��ON���z%"(�jN㜛w�m��QWp�Ֆ
�B��[��_l����X�c���ͮ������`+�O Fuλx噝�ofsq�b��k����]�e�*�󅻍�����@U)�������BC�mf��e����"�(�1;B���'	zw.���I�ۅ��5�􎫺�痘Gn�	�d�v�W�f�+k0�OVQ/O��^]ɒ���#�E����p��W�p�Kvl��ۭ�K��-�U�c3�e�>��������֊���v�'���U��95_8�Uف�w|���fN��֓*攌PdT�/��� ؀�S>��&A���Y.¡dj�@��Kg7����-�qC��lא��p�#jK){�͜�c)-��Fǽ��v���t��9]��5��5��R N�bpD�n$�)N5�}l'�����+d����s�	�;�
�9'7A������_��h��`�w���/;��W�8:`k/MlN�v:XJ��S�C o���>���w�Q���@���s>n-�\�U��W������9���wuQ�Ε�~������A퀈�fs�����7���>7v�۰�um����
]^�n���.68�wyH �A�x���9�{|:��S&DH&T!L.t
�8��U��q�"�ʪ�v�G�l�翬O~�!=�)3ü;����*�������� F����q�mzm���.��(Ј ��R�����7Tk���:�"5��R�S�8U,��@DgZ�����D6�O�h""�{SYF�M۽aR��ɣ��� ��R#Z�|[k�ߐ2]��;�!��	#]�%�"��MD�h�£* B���^H����v٨#��f�A����u&��L��CRł]��{��}]����'sy}y>�M9�^�LZ<����=�g�O�~�7|�R�@qcӒB�6�G��ƶ��`�i�@��_�!��Ǟa�5L�{��6s.��B�rR��ke,`���[�h�m�{kU*��/���a6�9� Cn}>!��x�+�p�Nŵ�-�c����F6�`"�<�P �ڐCq�����7����;�!H�N-�x\eDS�=����b�)������Ϲ� |�) ���n m�!b];�w�]}�57��z�>�$���s��˄��%�i�D^�v�ŵ�m�W��蝋�'w������Dnډ�PG.<���� An m�e��6�ݙ���v%�ø�NA��ݰ�g ����7��Gt�]>EuY	-��͡Z�W@�tt�ܹ�Wgv���4��X�G<�3}2�(������xl�q������=�|���B\Vm�WB�J5+6���T��rj��a���K�
R �m�oT���ye5�`3M��Qej��-<s�u�"�](��&4�t�u�
�!m�Q��01��K���[Xv��H��r��f&�i�L^Z��v�K���J�λB^��m�À4fK��-#ĺir��s��Q�_ߟ���R�	snk��l�2�nYCL�v��<�!x��S0n?����ւ�������;][��#{6��ˬ\�P�c�I$_I1oL]���[���=5)M1=���[8k�癆ι|���eX�#��>�\�IBz�͏y:�n׸���R��o��?	%���dH�_{;���.s�%�H�7�|�ñ�[ﵫ�Q�7Ve�y3��2>������!�<;/�j�����u��I��몟���HD��՟p����=�Rk�� �1�l���5î��!]�%D�3*df �y��d�c������2�</nY��{��F]�CӬ	��%�埼x����h�����h��_M5��u}
�u�WXg,�e���X�wRsn�W\B�����Y�SE�+a<y�����{��&���!�Qx}пN�vː��v�����Wq$�$��:�NU��f��&���&�ټ��3#3̏c|v&����Kʵ=̟$f5���\&�%)�>�f��5�B]/<̜�^̌�ͭ�M�r1��u����9Hv�#v\�	9��.�-��,�}��Ұf�୬3qr�ޮ�kLRM�-�#�gg`sV���I`H�L���駹��~�,��'o� �nI.C�?t�׾>_G��5���u���} vff-�J3�Ҵɶ�Hd�Ϸ����*�_���JjѴr�}T�"�����;I��8��zm����y��]9�BGݚ����&��q~�<<�%�����?2�l;�l��`HD�Iuu/�Ů���������[z;�m����y��{PR��^�g��$R��_�V=��n��n6���NVJS������=����y��N�������P��I�L$��.7-��U����R
��\o���$fg*�t��ѯka;Ԍ��:<9�>�^�!KI[�F��\č�^�R�7G��ۍ&�ټ��d����-�����վ2K�}0OG)Q���£-owDp�����@���[��LD�3)�e�D�8�&����z�{���3� P>��^ };����z�[��ڠ�#�ȉ���K��Uަ������?;���KR�{�+�F�(�8Gv��[71�C0��3ݗ11;羭Q���7�\w���9��?��x�*ׂy�B�	"f��fXh"$e#lD̠K"9�`sϝe:�R����|@���qo�h��mv�i� WT���g������eq6׀�i���pd@����f	�3)�a������j紮���jK�"�ʫ�IVO��!�t���h���RD� )�Mr}��%�'� &i���Y�/讀ީ��y�K"=���"@��Be0̴�9�2��]�H�z�."B}wh�����7���8���A��"u@�D�w�@3)*y���+��N��:��y wH�D�e�Y��DA̯�͝�KF���дm��/ܫ���s��@��p�v��;�3("< 6׀��|<:���;^r
vx���tDI�Α5�)	"c� B�����{�e�O� L��|<	�)"'�3�7}dG}��t@�t�d@̤ �`�"C2�� ,"n:Du�t��z�y;ߏN7;�����ꁸ�3��&�9������� �c�����a��յ�A�v��O*�N:�%���
dv�.����ǟc��M�Ɂ�E�������'wN�����:�����2���5�v+�kR�J	���2f�:\��:ط��f�s��n�yBZ,lZ�Pl���-�^V���f%�l܊����K[J1װ�N�ņ�J�v���)�.�ٙ�=��q6������%��eՀQ!l�n�յA2�B�m��Wլ��@%͖��>��K��,v��`�뱘�!]�f1�4m�-�mV�ޒzߚO�9�Fȉ��̴^`fR<^y�tzg�Ѷ������xm�ë-` ��b$3,@�@32�1���I̠n"L���8��D��Ax�f� !"]�C���2�+� &ix g���$�X%�̰7�����ɻ�8�p8�@����p7���C�q��Q�� WP/��ؘ�������3]�[ �T���s�lD��iP�B�$��@D̰�+|��w~y��#�#�v�sߖ~>� ��7v�]�|vV�� ˤ��v�J�:�&��%`��@v�H9̴@�A��elD�fiD2��w3�8΁!�(�&��7�5��5�,6DH��H�D�t	dG3,DH@̤3�_�߿�����K徲c3Sà��)��%v"�պ9�HKu-�Tֵz׈� �k��DI��K"9��H32�5�w�w��7���{�� ُ�쁢��?
< ԑ2�t��2�,��a�"� |<&���~_����M�q�A�A�ER�T�&_���ك7Ef����V��,i�u3nY�
��ߛ��u]�=V]V���{��{�| �x 3i�玸�}�.�:���_sh]ȉy�Q��؎e]��ߛ��W��4��Z�{��+��7!��D�̤.H���w՛�ι�W��oµ}�ǈ�,7! �t��I���#�����BeD����GHK{����]��� ck��m��__խ;�� 5 ||<>��"f��g^ux��=�{�. fe���H�3(�#��*`������<�����T%w���[@��6DI ��:"$�D�>n< ���y�B��gTCɃ"erl�.r�k��t0bg;E��&b��Bjj��?d��Y;b$�kt�H���&�e"�Cp �Y�����'� ���>�����u������ȉ:��7�$D�3)�e�I ��DDu��ZT��X;�</���� G�z� 5���,͗z� 1@��A�� �<�-D2�羸�!<ާE`',M�. g��h����@����fX"e f=a5����
�tR�j��͸��KfD֪�p-W���v�e�0��h�����P�[a��5��r9B�eE�K��}�xxx����wϛٕ}��:�F"@�y��DI�v�a̠-������� fP\D�$��Ϋp����"L�:D��� $��@k��gy{7����mZ��dD��Ё�}W|�k��N7�'��E���be � m� ����G����b4�go1(=���)��Gٿs��}�Vl��� Z��9� y�iD��,"e ���5LevDFQ`�1!}&�"&h7\��&r,���K[i�mCUJXGd���zI�{zI?^���<�.#���� fR�q�9��~�������WKy����`o��t�uh�Dw�ȃ�����AqD3(��5���R��{q�k� tx@� �f� *�7;�78�����[@ָ��D�}�7'[�3,�$��|�D�Ω�}�\D���DI�h�̠�xk�����GtWФ���՜�~ W4���<� ��$A̠"fXj"y�<u�y���D��X%�|��t�̤8�|���w�{2��x���m����`舜k=O��P����юt̎�2������]���*����&��s��9�t�k��Yȋ��2r�}�x{�(@�ґ}��@3(9���fP6�Hff�5̤7�T�q�z�5�'Q7� �<�S����w���^�5|Xn"B��"$�v	q̰4@̏ ^]��B>�����$�(J����S�׶q��ˆ�et�fWy�C��:t!$�߽DD��3(��h7�y�����֝j� "��������Nx�ȉw�D���E�&e Y32�DD� ̡�淝w�g��a�'�  �@{ !Uw��j������7A�"F�~X:"$;�D�#�@s���<�'��sh <�ȉ!�t�I��D�̤- x� &�d��H��Tgۂ9^��/h�m �Gqu��#����e \@̠��\�\rg��N��� �Z�t�[��$ fe�i�;ý��M��w{ �(7o�� C��8�����]� �� ���;�"fZ�H�&e�XD[h�3GV���	 eǀM���g�wǛ'z�����n"�ߖ�$�-�9��H@��Pη�w�YǝnUs��u�|$I��n�)����7g����M�Y�e_L�{RSwQiP�T���a'�Z�߬��ʷ��s#і�V]Zs��{�:���d��LD�#�+p������,*�gay�ː!
�j�m͚�;2��F]�5r�V���S�%� ;�RբP��ˍ
��5,�<�Qb��J�-��Ԏ�&0QT�N쪙�̊�:b)��"���d�y��|h��X���N�f��ol'��4.(r�����2�6�u��	�%�3ʒ�O��#�p+�^@�j���۹\�"/)�Rf�V���,���uGT��BJ�ʾX��>�`�u�Jx�t�[Բ��>+a�2�l�\�#|y&�5%�6�+EQ��6~0.C3�A&��$>T9�Ee^^*/9�`���գv�v%RQk/�rs6�q�zYvue��k{�h�2�0�+n�m��R���g_1^V��2�Q��9R#�۩]k쾩�ۏjqoq�Gq�IȂY.��ꡣjX�A(qN��X{a�C���t�sX�z���ݶ	�X�:�h��$WXg_=|P霞,z�B�U�D���;⨭������\兂�Y��)�d>� ��1�v���Ҿ��{�ez���oA�N��CP�̅9�3v�oU���O�����P�A��%�-�?��ݹ9����2I;���ݢw|W�%{ޮ��w)2O}]﮺�%��Jp6lZ�	m�	iI	@'R�gn��Y/��(�s��v�]�wk��^������9̑�}�/]�w2��������V�����"��K-�˩	}+��L��n�����<��4��}���ݯ��s���y�	9�v$����`O�����F��!5b88����m�B'�2���nt��ٱAGuLFin����GbāEq�Y{\]a��\8�dΛ2隥#X�-����C1���Hk]��j,4��mW��)�F�s]G]ZgUxv�(icS���6� M���P�YMP����)q�IGr���D�]�2۬3f�*9 �Y��2Ű��,�XA�3��I�hh@ѱ�j$�v�b�gq������ �2���fa�O�_/��#��D�x>[G���4И�VG�)%�����mF2��LM��^%�%��-]H��:$�3rJ$ع.�2�04�iG��3K��:��W+��q,H-P"�a�QҖ;Z���ܐ�GH�L��h^�mF1�f--�큀�ళ��[%tRJ�d�6�ɦ�	j�@õ�5�+�fX]H�tY�+��tEԮv���YA�4�G8]7Z���)j��G5��y
�!�F�������G:�pPŅ��M��ܑ5ñd�S3Ae�4�Me ���n�.C#�l��jڴ�!�閆,�,�s,���t#.��$c�:��e��'�o$��R�l�T��2����ciG��- ��5����u��&3�J�mf�G"�BŅ��R�Y+4����ܣaa��2��k���6qr��"�`NSM,#��5��%���+�U��ntR�3�&�v�vu��%�K{�6��%�sO<ڀ�B��4<&�B�Tc��j�JDI�FjVU�ꑱ�L�m70�2��b�6�Y������9�U!G;k��G�a��+2��Zʼ㵄����,�s�j3^nhm�i��)�И+�)ʺf)�g)���UnWeUUUv���y+w�%b��ڜ�^S4�wN�Fo<�\�[v�-n�x�"�l�u��WB��3B�.�L^LA�.u#n,�,��KbB5��:f�3�ۢ�\-&˙��6�-X���L�s�Z��k]Uΐ2�f�eй�X��i(P�q��53H�Km�h�u��X�ЗIJB�k�#c���)5i�)C8
�bֲ��(#*S�ϳ���b[��V7I�9�-��; ƻW�٢��i���]j��p�P{`���oy�5̡.
H��|�>^��U�vWY{@���'E]W^wTw���/(@�@<�,�e�DI ��Q�����,��h�Dw�dD�:�Z��u߇gg{��]��
�qw@�<�-D2��a;�]ֺ���vDˠ"}sa��}�7:�@� �|<�ǀ7��L���������sA�� y��,@̠8"$`fe�h��:��������@3|f�5��`$"fP�k�{�[��W��u��_V����l��jy5��t	�#�<�4�I�(@̠�"�e�̱2���y�g�S��;��H�� $_�w�8wۗ���j�qw@�#癤M@s)"e h��<�u�eT��c��FQ�,��gl����])��K5tq\3*��$>:DH�8�#lD�y`���LG������;M�f��6�w���|%^�;�]t��l"$8��<�^ u� uA�D�C��"&��{�ڞYfe~�n���&a����mR8�5g4k��N�VcA\�wo*�9�]]��vr���x�N�������W���;�m����/�|�ߧ3w�vk���j�7# �T [��ȏ]P��|^����i� q��̠m���D�#�T�D����:�y\y��7����ܹ� �����D����c���������>�Y�k�<������^[.t&d/�ų�l�l'��u��d?h=������ɷg�����Cs�׻矞켞9ղ1VZ�H��d"�������K	R�331��l!��`�N�tOzn��;�W��FN2��/Ke�d֏u������n,٥.��wZ>�o�bqz���F��e������`�2�����
��52,�=:��ÿ8���s�\	{��U�ݫ	�|�s���Q؈�Gn�T����8��� �\�~s?�v���`l�!�:��^Ю_gVT^�q�vͽ�)Z+�]eE�q>�n��g͐!���5P"B3��|�?����L���~��~'����]��a�WDF�](2\�6��g%�ə��55AXS�1�qwo>}k8N4�Z[O�s�Y�v��g��l�a�&�׽�=�=���A���u���uǵ����կg1Tm}x��l��mp\���'�7x��Q�=8�t��[-��M/��
��.�t�w��o�[IpΏl�1�ő<dG��+���I�ֻS6o�W��Le1�x�t�g��E�%���r�6xو��#D��2��S���� ��?����6[!��N~j��_(m����yyv}�{Hl��,�T��PO@�P�u��(Q�\�p8Hv�"�mC�4Ф�.�j�+�P�9�n�_JZ�6x�t��TnUţ0�f���l�����i�c������;ӣ7M[Iw��m���b�7!�3�q�q�w���CS��Rl�}̎���g�E\��[��`�B�������;��{�1�~=�a�[?6[!�y�ۮ�#��������>�n]��|9���*�m��/�h�=kc;d�"�p���sP��TK�N�H�F��g^<�+�;��̳7�G����]��(a"��SFmQ�-n6��F�rЉe��6Qd��%D�/:%!V�#lF��e�n�ب�յ����e����Ixsn�8�� �RMZ̘ܠB,
��t+��Ɣ�e6q?s��Jo���:��XT�2�n�M2�Z�\��L��W\���j�II����������e�ՁJ��K=���q��ݢ��,ƶbT���r�fhƢ�I+`�M�e]��������l�q�W��}�0ᕯ��U����V�!�dx���*���|@�~�+��;o_[H�{Ϫ���sS8iE�P$1�����nي�[��Rg����uė}�܋��/cU3��G�y!�Ǯ�vɸ��|��L̕�;̚���я�ql�?6[�+<�����b���]/o��-���w}�3!Uj�6nƘ&�BP	s0�f�`���)�1h�Zb!.r��O�;�������|����w��6L���u�>�n}뻹��a�|�p�����Z� �uw�a��թ�-{�C��k3UG�ܸ��ڼv3�������u�vU̷���P��� ���}�����6'��tT�+�w��;�0�Ӏ�d4��x�b�^����М|��1gY^x������w��ﳩn%��� ]����O�d캴�_G���SS�{�|~��d�sy��~�^�cɾ=*Tp�Üz� �����G.�~R�K��0� ��݅����\щL%fBk�CA��/3�@�Cd�s�	�s��k6���o�N�`��?6[?���W�*��!��;�6�;˖�w~�Ѕ���I����N!2�������UQڮ��s�;���,��n���<���[w���zO��u��VŜk���ڈ.�l� �������kc#����t%yg��[!�٭�=�c����{���[??k����|��b�|'��s��sQ0.��������e�}{��,,�n����;����]߾~ -!���!�qW�<�ev��WEm�AūԺ�;D�B�L����7V��ᱵ�����s�U.;�Q먕���[��p�O�l��ڋ������i^����|���^�y6����!L��eϞ�o>o<c��z��[�վ\����~?koͷ��"��a� w��w�)\���F����2�^���X=��ѹ%s9��n��!Z�uy�Շ3v5֝�{y�ꓶ��sw��9�U*M�3$h��¤DE����������x>l����d����{�H�������e.YJo�m�ͻѣ1�>�D�(d�8̻`��.�����e!C�ea4�[uA[���O�܋����3��^���P�Ӝ'�M�Fg���g���n��籤=��������1y����=��uw�g��㬆�l��z���J^��z>��\����)�����g�Y�[;l�~��=4��}�o�os��yu��2 6[nŜ̐�g��<A�-a�T�ήπP��o o��1yV�h�>ݰt:���8%�t�N��#8�\��G] fd�K)�;H���θ8#`��Uޝ�Z�򢨋�����@ ��6 �f�[JҰ]+��ڶ��U͉�R.�����Z#�V\V��]��.���F,�ef��VWC4���aB�E�-t��^4T�6Ҋm
���;kA�RZ�M�n�i5���n-�G/溥�sU!��e���W��[���d��`�a`�7b�E��llX[�@����KO���Ja��k�k�0�L�3X�i)a�/�#�-?v��͗�< �������L�Ǌ�{{���y�͑An�P*�@�[9�b7;n\�\�����[P㴛|�6[ 7�έs�;��������)GY s�]���]�W}�����!��q��/=�*�k��S��wOr�!�����l��of��9K~L��Ӝ�w:�u0��
wr.�T|��G�_y������QZJ��t�+u���,�cA�fz�%��p���{��9]e(玭�zc�ۓ�l�[���S��33�0�>9~dac��A&���ٷJ�glU���ט!���׭`�(�c��]i�u���k�W�N� >
��H<?^��9��w*j;�<+#�bi=��O[�|Gx�d|���{D���}�;���梳~qO͖�d:��z��q�pj��=��9���p�7���k�������!��2��W�����I޺阏����l�݊�2�݈b7}M�ٯ]ֆ�^�$9��3IJŨ��e��#b�+<�#��[#������_8�߽�������-�#��gA]|�˫��],s��)G^G8�//�՛�����d�!��o�}�uP��
�M���L�����u��Z�oB���D�p�����,��q�����D40N�-�{xl��Sxj�˓
�����=����]��J[Sj���y���iT3J�	z�����\���u���u�o7c]�ucO�F�8bB�W�c~堎�܍ӝt��ݶ��/z^mUX��-A{2T�ْ.�Y��˙u�i�d*�x�<�gz��|4��0�5�ΉlYB�Ǯ�}�[J���N��/Y��Rle�2���dNC���J�N� �K('��f7�-5eU0TK�vm�l�73h>�1ϻ8;����q,x�P;R���u[+1e��IS��Nﮆ��Z��k�4��dQsJ���"g�UP�$<;�m�e���j��8���+�d���wݺ�.n�_6�=Xe8���X#��7�:�Nm��ݕ�&�J!#[��R�m��-�u�e��-<U�ٌѾ�/P*cki�L��7���oB�,l��r�,�-ݒe@�ӵ��2tɘ�V��nf��+Ty2�*u��u/H��kj�L}�s_S���ti �gaʧ�x���k3��jMt������W�~�b/dr,(9Q)�W�N𽽪X�ڒ��X�}jn��Ci4�hћ֬��:�����=�	'T��r@�9s߮���#�zU��Y��_���rJ���;\�\�F��{֋�W7I�;�wr�v�(��s������Qh�y�2[�wr�w�뻴SΨ�g;u�h�{O�N��$�t�ӵ��S�C�	��-׀-��c,�����.x�Y�nj���r�L���Mï���r�;G+�S��R�#r��	�tش0!$�sr������j-vۤZ��,o�վwX�������t�~w#Xϥ՟� >_��-���L��������M�?o�M����q������>����~��i�VN������!�^�r��q���/���R�zU��8~��˹v��"�Gr���FDD�$̈2�s��f��qB���ܑ�=��8M���^^f	ۄŲ>n��>>3�oϬ�w.S_n���g��/��v�j�x��<���X�����\��x����Oz5�m�8����~d8@����m���0}g�C�a�NFGp�}���͖�Q�駳���V����[��z��:^R����>k�)2�3��f����۞�Z��꼙)v?.�y���#ט���+[ᕏZ�}�3l[�S��d<5y�����}��ߋd|��6Co��=�ф#8�Vl�^3۽�a��~w�<.�Q2�A�ڂ*2 �aK1���,ѹ�6Un��ef���T,_�fffᨎ��d�ck'�#GaEp�(NVJ�F\�6~l��Ja��	�3U�{�uK�]��l�v�
[�o��Cm�l�_}=5r��3�{�a�zd6~l�ʺ_>�w{��]�b����NF����+*>�/�8{<�X���!��v���,��}I���F��Sq�v���w�z]�,�[XQ��կ-��j����bD�j�7N��;}M�\��d��8�I0�bFz�hX�݁��f��߼�M���!t���S��0�c�G���IRd 	��{��gT�.�ma���ssa]��k�SQ�]2�t0�	��Q� ��uP�jVZg�Nn��K��",�q������a.ΰI5iH�q��-�����Ɋ[L14	]�i��;�7a�F����R�{L@��\�Q��1�퍡f����~�[m�
�i�[�kp/\�����RhuR��eZ�7���|@�!��|�c���{w�,7��q�檨�-}�6�|#�Q���N���8�O^^���(xyU���O��ِ���v�Nu�{�g��x9E.zO��&sܔ��g�{��-��#ճO��|�q�2�y�\g�{��~�����^�I��yL��}wq�壖ЃY�=�v��</ʍ��{[����=�4�ǆ`@�"�t�
B�JL6&�:�9{VV�u��T@��g/(�v@�f����q��Y�!��2��w]/WQ����p�=wo>mh��F�S��W}�<v�7��V~|��Z�6��K��b�'&���ߦZ�w
�t�{�t<�Mi��u�  ܿߏf&�����wE���~?}̆�Y�Y{������!��uFr�rD�y���S��Q��=���6[?p��έ���C@s!���B�����g�~��M@z����g����f�<;Б������a�zs��o��f~{�H���=:�S�� ���k�k-+�jK�3R%#v�y����f��7��.�]��˶��6|�\ڳ�-�l�����J/gU�@����q霉yЮ^���q�m���o�+_I����e�\/�}mmI�-d�<�P�K1����H�����߇^�~n��v�Mۏs��ke&n��+fU�g��d��� )�������r����̶[-��!���zz_Ug�?=-�������4M����W����G��?�Ͷ76ZnJ�ǝ�>���ިm�!x������U}�J����-ʵMJ�,,s6�e�3l�jUl�*�-.�<,vvfc�d|�.����N�uw����f+����2���d6o��߉�h%�ƣ��=w�w���ܞTj�{�io���C���lw����g�٤�9�Տ8$=�$�Z��T7K�{O�l����+3n��=>=�!�Cdgcx��S�t�۫���3n��ΡӮ۱�"ݕz�N̩E��٪��1ɅUtsU6�M�'���n��=T�&gf�W*�ќ__�m��7���~��oW��oCsT��$�W�2���i�$��B�, wi2�,ڪn3�)���Ա�59�8�&��ffvY��}ב븻��l�Lw�i��[�f�y�l�[?t��l��p�oH[���n�Omt�۫������k�F0!ǎ!��|\��Ά���k���3�i��!����_��Z��8."����W�7K�{���#���቞�?�m��4sF^i���'���=�=�Ϸn��{O3�g���+9�>�-%wy�RT�ez�ܔh����-".s;|�NIFa��꨽*L��)Y7K'#�??]�}z���M��5G�Z&f���Ihi�;	J�,@Mr�a��G�h�`Ժ���I^�,]�U΁��s����2.�6�X���:�M*j$�1k[��t4�2��N�Ԗ:��R�@%�h�ڑ�)R�����u�[e�5����[\ో!Zm�hb���a١t�lW2�j���8��o�m���l�Qr��P��j���-�,����Y�y��vB?7�S������:T��\�<�!_��K���l��y��އ������n�*{�V{G�7��{��͵��#��C����~l��R��N���)���s�[���s�[w>�����%���V��@lx�g7��ro�:^����龲# (����5&���Om̬�P9��;��!LpݏuǮ��a�:��! �iD�H�����"2�	Mp�T����X)�	%$��S�f �s��W9�Fv��MT��#�s���N�{��@m���7������N�&ff'FŹ[��MݜکL��U��Wک�bL�B�%v�H���w��� <�����,X�͛�;5��!n�
K���i���79�}��xI�������u�u����[!��f�Ѫ�n�������oC�u���p[b�+D!l�Ce�U\��V{}�b5v�vw\3|�������l1�<}��Vuv=����Z~PV(�U�ӳ4��y�7Q�A15�,%.jg!�y���-�%"��ٗ����{����׎�{_|�|@��-�ٽ���R!\���\��NpyӸ�����=w�kJ�(���gѐ������c+��s&�� ��m���ѐTR#\�̉Y9R��8ڳb3��Մ�'G���f1�t`b��JE�]������2�:��mt����O����Cg��d/�o��o?���<���Y~�=0��@~��w�|�p���?�͖��w
��Q����s��gr����n����>����%���Ł۠����ۡY�L��TMcu��xff`�����Jbuw��Hw�˧�/On��Q���6v6[ 6Cw��Q�VU�38�im�9/)������@nΆ{�e#����e��g�Z~��2cO�����O}��[-��6�;�śy7p�-I�<��}\]?|'��3���`��=N���*l�zov쐭���3��v�X���Vm|�t��L��s�:�&n����L�������|�~��C�l���6C�������v�y���_�����qe��~�k��~}��=�5�c,�t%F��U],��i�6�� ���˼�̕7l��Êe�O|+|�eOS�نǜ� ���?6~l�j^���Ў��:��V�����~�t��Csb��<�O��Be�t��;�Z;����/�;KT��F�=�G�l����l���+���u{�z|.�J�r�y�~U2����-�{���Y��6�}�e�F/�wS6����ӂ����b��q�.�]��Bq�vt�eJ�j�ӭ�S��5�:�3%�	�Ղ\�L��0j�[�jtT��	����F�?K��ЩۇgM�{��P���K������i"bހ�(���C�`���a��ne��1A�,�:�:e��@��ݭ/h!L�uai��f�2NmP�}{y�4��5���*')�/Gm7I��$י����"::F�n�)+�i����Q�|�i;��D�gWƦ�{sZ����;Qo6���8����w�1�5J���nB�5v�n��ڼ����М~�p��o-��5�Qڶ����+C���<��W�S)�⭑X�����+��Hf�޼�h������Rq��>�n�Jg\�eC��\��"b�}��m��:�9��N�*��)�Y��(=G�܅:��JVD\��[.�t�_r��ȶ�M�u*�D7^Һ;ڴ��4�Պ��5̧k�dk��{��N��B|]�c�*VЅ��}�kU��'](��ݗgoT\��#),2�34�*��a�Ĕ�m�(�ГW ��XU'e����x��0'ZH��Ț/+j���;ի2��!=�ű��ޑ�B��f��+c�6�Ӷ�@ɩm*�^u抋��+׌����+���k9�Ō���y4��6ɩ�����&l�Qml�B5l(�s��.�+��C�O ���d��%�M�QQ�\��j+�r�\�~�����QU���չ6(5���-�sksb,W"���5�Qh��nh��m��-�4�棚(���~����wV4Y�[�m�ݢ��n`��(�|�ͷB�-s�+�nsm%�cQ���؍���$�6�cQ���ܶM�X4`ƃk}6���c�k˔��Q�mͺUF�b��\���Qm�-y�6-o���t�2�	
�A$�	
�VvoY���K5�a�k ���c*Ak�fk
��5���C�H!�9�L��.���M��퉄&��V5J�e��˄�?��4<.��&�La��s�6�Rd�aX�q���q*�nWh[���F&K�5����$��f;Ԗ`�6��-������_��ˡ��1�6�Msl{��6#��m�v��d2��I��,a7:�ƶl���.�ZFf�5i�b�LE�hf;cLKmc&�n�h3�h](B�GD���J�it ù1L`"�yٻg��ɬuV�ױP�#m38cMP��խ��6����f�9 X��1[&D��v��lõ,���j��2 V��eM�ma!ՔXK�k�Whh�0n�e�eV��W=�UI+y��q)��%Ѧ�٠1��͚�f���Kut�BT5͎�h2�9䔘�q��']��Z� �@D�Yi�%��٢YNek�pDƍ��Ƃ!K;ji�&��h1��aHX@��b�usL��RB#�k�`�b҃��+� ��a�V��H1
j�cb[ �t��N"KHۙ.�Ōq���c�bY��e6�C\�sC`7V�������v\��,Ը��j��a��h�5ؗ�`�b[0�n��rCUH2�MKZb �,�\U�\�n+]��^��M@�t[t5���a���g8#�J�Л�]�aD�RBfk�fG:�ZB�Dy�7Q�V�e��hun�,�Z�%ë�]yy�5qi�*ɵ
l����I�`$�-��KeHQw	6=v�z�+�[pf�`��HCSBZk�T�E����o1�g��*��nF�U��r�ʹUUU[H��[���#��X��2j˕���I<o��1�@����sn*@�&1����d��p�]�m�F�-U�י!Ǌy����2�1��fb��PЎt�.u�pj���Q�k\n�r����@���²�Ś؆XW]sc� �6���v/9��#����سM։iQ���v�2�R��[\�+r�s-����g��?��J!n�7$Aqa)f�n�q5�� y@��y��7���#����͕|��^,����u��t(eo�c��ql�~l����˾sz8�⾻���_�;��=��[�����,�խ����=vs-�7;6���K��a��p5���o+�ai�oZ}|�O>��6U�;�f,����u��9�(Ι=��C�Cd�d6(P�sU����S�b��V���w��{��|.�t�멊Մ��1p�k2U�6\�X:�39�2���lc�.��y��=���ף�{�r�D�|v��* �����r.���@fn��7v�`S�$D�F	a�x�է2<�J�Rɼ���^�t�}�Z��S�ԅ�O�n9m�ѵ�Go��e��oՐ�GU��_c��{wv�e����/��{�������ţr
��g��^����������ϩ��v��q֏�v|.�!�n�tL7��3ݤ�h3쫿xq��x��l�[���T ��/��^�=�n�o�� 6]�=�=�_(B	�LəFI�$B�H��v�9�-�����R&
II*f&c3�u܋�
d�LGm��~�&U���{��������ۿK��csc�\k�c��&9�i��f������r��&#�~l��z���_��z��%�Ӆ#n��n���h'4d�4��ϫt�VƝU��g-�V�Gd��N���MC��z��k}�o��W���U�~��^-��l��1D�@��-�̥¶s�|�h�����s������?6[?6��B7�Q�x=������5����z�gs�)����)|�����:%C3@��qu��M6����t���ȶv|�l�J'��Ezp�ʺ�W���Z;��w/���-��p��vy�o����p~��?&{�<y��yr_��61YH�����p�\��Ʊ��>/}�w��rϾ�?�-��@�qq�][��y�l�Z�{3��p�Uu�zG�8QA�c�R����K;F�We8&�����#�&[�,<Y�����n��Ғ��O,�P�lb�ʯ����G��l�����u]XWO����Y釟��'���d7oj1��8�U�`��͠�CзX�ڛ3q�d�&��L̪����dz�.���m�;�Mt��T��X��X�����ͷ����3��u����!�i�S��G�yU���=+�68�d���6߶���v=�D1�J��zx�/���d6[-��f7�w�^��}��y�q��\��y8���uQ���j��ų�e��z<u��y����E]�u���z/��]�pt�x.��"�\L�8<��DnT�M�afq1&Kx�!Z���ǃ������Zq�M	y�V�UA�4a��#�F�2�A4�Cb�"hC#�^��.��Uҩ�R!a�j�.�������M�ƅ�M7i��#kZB��&l�����p�-0�G$&+��ikC�؄T� G0��%�ͣE#�QWl۩e@�̲�ڹV�1���R�-0B�+�خ�^8*�GdcV�aي��Wc0�3�ϿA����W*:,3,K���2ݡZ���f���eL�%��q����]ǥH���ڜ[�"�����*fd6[-���v�o��ͫ���k��9��;���]��JPR������Cd��u�c����h�k�Mj�
�������UX񳵺�úCg����:x�/�x�c��<{���?�-��!�����y\k.���|�]Js+p͏wwq3j�.	D�0it^���������Y�4uW1�ڃnh̹g��ז~|����Οq�o�y�Fx@�;���ϛ &k\������P��7�]�gT�s�c�("3�G�{r��l)�YjrHٳ�aG�F���>|2m��KP2ȮuҊ�����ݱ��_uG)���Er�̷wPb�.�t^��d6~l���A�H�V�T|�8{�.E,�}�D���6[�8��ů{�f�:o||�s�:4��
ͷ�h��C���l�C~�S˒��z2O:�ʞ�4J�����Cm�男C��޲A�R0"�"d�}"�X36-�مL@ؖk�/ㆳ2�����l��UN���;&A��P��l�8�Cm�>#Ď�������n�:��O������p�<1�wr.�_���+n�3�屳['ZǤÞ6�����v'�����H�Iϻ���Z�Bw���V/w��g��[yx��`���]��i��΃_{��ͼ�6�Ib�^z��9����g�;�o�ǧz�ȝ�i��:�9�I�y�l�~l��*�N��|h{��{���*����[nM��U>���%�cT����tu���ڭ�-�M�]�v�|�$�?M-���Ϟ�~ʝ�4J�pc>(�k����"9�o l�N!u�T�^�����}�o�ǧz̑;>��7K}�kL��^�N�?Ҹ��l����ܪ�gU,���K�8n��zW�͟�og_�w�0ɻ��JwΗo�~�����y;�6��D����r4����UE,��ɅzT�T�LFRNB�H�|n<���=v-�ܪ.�¢�ܱ���*����~�?n����d7���r��х��vw���������-�e�)�$L��
i�XMv��ԫ�i̱��)�3JZ�
��>��;��`ݼ�<+G^B7ƥ�LL�۸-���Dyc�vd�>?yS�wΗo�~�}̆���7K̋Oɐ�p.霩x�U��-R\��s����K���[?6Co��x]vK��-���ȭ�N���rzj�+��I�TS>�_�C�7*����M,��VT�*���}tM���d�nRROQ�R|WY:�H��[���U�q��d�f"@�b���������Y��~��E)�gn�����ǝ8���@�vѸ��e����X��^�iYn��1)1Z�MA�V�7XKIL�#]a5%X�Tc��SQ����LK��ˁ�Dɴ.�`lMū��֎�)JV�"�F�F#�%aB�+�V j.���ͳl9��U��йi`�W��h#L�,t�{f�̫r˲�����>��(k���Dte�ݥ��B:����&�`�R괮
ffgO���ܻ�]��5ӵ�V����݄���Y4.6q��=w��U��{il%��V��0up��M#|-���]���zW��r�.!���!
�;�t�0f�y�P�zD(������x�Bِ��!�7\{n�TA�0���=��̀�K�l�d�o8{7^K�������R�͊�6u��p̄�#�1{2;�$����$ʅ.�h�F{�4�Z�8�/oP@�G�bbkNk�Z��a(�2`L�]�tˈv�<��`14q0�������޽ɡ��. �A3#�1䦏dƎ��|&"w�����Wa�GD���[A��A9�����ͬ}�d;�5�I;.���W>/EXm�=�{��^���񹷄��	�;�%�Xacz�}�xȯ����0v��W_��� ��AO:�����U�/_Bh Fa&��;�^ &�2��ly�9���!ݛ۽w����E֊�T-w�' �P@�6(W�X+j0�2���E����K/1�xy����M�
)��G9j�3������'2 ����܇�t�B��)�WF{sC٪�]�7Ј#Z�f ��v�^W'(ȱ 	HDj1!����o$�q����B�M.)�3.P�{ԇ�/~|��̄A2��,s�݆�UP/�<��HV�w�3H/q�3Df//fG�d+�Н�7�^%���9dw�OFl�����Hm���)3���t!��3�"�>�^�~�]�쮭�=(��9?F�17P6ڈa�ҡ�b�)�qjt�此q��\��9fQ��Z���W��Wq�$F���Lw)b���w���]fÙ¢5X閡���!P�ꖲ�4����gps�qn��V�:y���ٽ���m��/��Gs�,�����u
�gl��yYC7&:]YG:���Ex�of] �$;��vЙ�sp�8��5sQ��:Ϩ�~ﳤ�o,1�Yڞw�#-
ݸ��)B�v��.��\4r��m�"����V��3�r$�`s��v-=ܺڅ'��C����PDε*��ll��UR.IO���j���n���J�^Ih��1XF�DXvs-�̋�ץ�`�#�1$�{e�ҹ[���蹳Mec��x5;�.��!UKd�	��徙s�_կ���Y�Ĝ�&�c������>��3]�����	y���Ut�ɮ�ު����h�\���Gu>Zom�K]�U��#&���"�N�\�y�u�
'��Oz3�i���^S�f㳳B����F�N���8�3�t�;�������l��6���l�;���囌E5b��+��o+v���VLfeX�1�uaޭ�6����x�<�HV�c��g��V����2�@㉑+sel��ݸP���]i�;g��n��ŋ�\8�8���۰s"��-5?;U���5-y��TPQs��XŢƬj2[DQ�`�*+Fƈ�U��Q�lmc%b{���t5�[��1d�j1��6��E����X��Dl[A�h�Q��[�T-�ڹQb���W�r(�EQlmI��4Pm��m��ci5�>��(ך�k�ڋ%�l�U�F�E�آ�6���Z)6�nX��(�T����Z^�p�j4X�����my�-�i�4��6�	���ǽ�,�N��g�������7ЁkA���b��ܓk��iđ�p�A9�^�9c��n�T-p@��@P�����a�F�P�b�Ib���3Df#�J����-N+��wLS�Q��A9��/�G2�'2+�4���Bb�5��h�k�պ�n�T�����7V�����}b�j"�N"���%�=��k1w��ג�;"&h��`���"�/�̄A9��cH�w�"�� z���Af�r�<=�Q�-@� �����;�gq�����
�~��BK�Ibo|:k����r���q��A��+�̄A2#1��+N�ځ��6�E�y{1�7�w�3Oz3fkл�o�ƶr��}���l������<;����hHl���QP雜�ﳋJ�QP��;g9��^S���	
tKK��'`>�P�X��ءB�7�	�IE~�?;_q&�N�U�W�4���#B.�?\�=8��U,%��H���pe�Nu�Ť����B��3r&�H�Z�����2�>��Y��#1/f �I��=ꨗ��!G7c3t���H<�=��o!x�ā2"i�O2��������h)Λ���.�vl*�\&� ��#3�S�Q�3��y� ���3@�B�9�ِ7n�G7�/eP���^��d/Fb� ��8�
��� nG�f ��
��/z�'8\D(���^#�Æj*��f��Ÿ^#22�d�b�&ߟyi��!/v7���:�g_Z�7����x� �F,j��uO��R��Is%"ImM�ئUn����a���uiMU>���8�L�Ƕ�&ʣj�hr�麄�̳�,��2?�}��_x��9L�i�F��J��7R�?u��X��Vͣ
\�T&Ãh鬶�!�"�Y�p��3ئ�uT���р��°�����M���b�2��r:�/J��F` s̯)n��[�z˚75[J��lR\�"� M�5��ں�� ��Yq�n��tk�j�a��\?~|�{�X~�l�n �:VLF�H�X�T�0��0̙�˨��;F��dQ�Dc��fZʡjfT�r�V@N��l/s������\z�av��В;�^=�(���i�UJ|."&8�v � �dXY�tC��R�>:�Ϩ Kd]	��C��,>	��+�T�9��:z	�m�K�1{2+�N����r�ˎ�Ah#�Nd��O^Y�p��A߅���b�f��>��X� ��e Nd A�@f��zuJ�:E+f�d�+x2K N>)��Ԇ��z�gi�"$($ �l̢�1*ii�$e�Յ��Ҫ:��mK�32����@�嘄��MǯW� S�5|.Ի=Ӱ��@ �yA�AAx� �d A2���ɞ���`����i��5����1��U<;O�[�g��΢�t�n+2+-9����%��'w7B�s�o����� q¥�s'�tzxnʡ�/^�^ ��9�QE���0D���A��������b�`��%҅�9��n".;�Ё���2#1 ��b��`�My��f ���l�uq˴��\�B"�����P�
��4�����B ��Df �̍&�˩�Q�L�]��t�+g�u+|�7��{2=^�!����>��5����f(\�:�Kɐ�lZ�mcf�@2�S0��؁�ysA�Y�U	��<&�M�Eǐ�s��p�A�Ds! Fb@��@@�Uv�w�b"3��u:���sV��LW��/[�A��Fa��졗br߷eg�vG�b�dP"�Ba�5�ު�ꖡ]-b�#�΂{���=�%_^t��k�7t�c��\�������z&a�ǘs;�m+|����k�/z��Uº�n±k��7�q�̀3 LK=J$t���wP@�i{2����;��]금��	���]0gs����]@��#2�̀�B�Hv��}=��->���e>�Q���	����^#1�3j3u�7~��8�Hۛ��)\���!t6�h�`�M5�c2�&�q����dW�'2O^��L-��J�k��z���.�V@@����=��{2=���t+k`�����SP��tw����� �����d^I��uQ�h��aB#�/s��̀�̄A�^�#��.*3E��]n�����.q�A3��#�հ`R���;�'��M�*T���f4c�3b�/> �����r���[��jS�5YR/Bx�AטiE�ZJ��lv����H�����]���P��z��Ľ�����d�a@2�����5��KsĖ@�~���!_W��p����o�K
�%���\	����*aK1R����\�@����D��SU9{����/%:��[O2b�;H"ǳ#ِ�`#���F�ҍBθD�*���<�Ʋ�J�k��6 ޯfFy�
ٽ#�������v�������'aɚ{.Χ*)�Qq��_B ��̄A�̄FbB�fy�[Эw:/g* w���7A�A�7���ocٕ� A��F��\LJW�Յ㺂2 ��n�	,]HKTX��+����ev�ץ���� |s�"/` s!b���0;I��_�BFns�z1�M[\N�/3�UK.��&,˹Ӧ��[N�箜��"�l����!q�t�~��.�о��8u�"B�MX�.Ҳ�Y�J�KF[����&��x��dYo-.ؚ`�(:����Ķ�6M�������	�����LY�(��R��Kh�١$�GC.qu���76!s�0��5R�%y�h�(s�iR�%tvcF9K�[x!Jlsie�M+1Q[\�/k�s��￿-%�R�E0I\��`\b]��Ԩ� ��FlX[�Pʮ����?oz�g������"�Ѿ��N�/�8Y�ْ��`+e�!�(UHo��!
sZ�߷6�n]G��A�U�W<#Ocڕ�u.6(Wm��!�����x�������6�Fb�@�2)��y�6ܧ�L>ҰR� A} +��d/b�ąoץ�}Q��ր��㘂����{���� N>�ۛ=��m�6(W»��]�!�u!�=�]��K%����U,d�_=�����@��e/�N�ɛ�d@az�R"%th��#ԓ-΁�ʷ@oh\j�	A�E~���!����9�� �B����0�J�K��iu���A�q���̄�g�E=3y=���-�E�(�
���!�w�����.���fS팔�Dcw�ਖ਼2:,���
�IÝ�Q�b���f�����? ��?3���b7߻��)^�D�ǸЁ�s"�t��i뫁g�=��s "�A�}����+���z{���O^����yka����,]Hl
�1����~�gݱD�
���js���U�\�� C�^B��u6``n^��̀�̅�b��
��=�EZURY���E�~��??�Cb�T��J�����|��.��1��։�Y���t6�b�"�hb��ړ1L���;�Րp+�2f ����5�I���K�@�ΐ�x�;��q�V�D=@/�̏/�@�4����j��[��U=���㸚�1b�/w@@���d+�~�VdЉ���%� #1��!W��|�w2e�y�Pn{�h���\*�;ӄ�Y�X*j��G|���,�+�+��d_\��r�Y�ݧ�W���t�����?�����	/��~�w�@P�+�~�$�c�fŕ�I��ԗ�� |i�#,+�qUn%0)�^#1{2(�s!��#]�Y���Qw����K��\E�\�=� ޯfEx�3���Ol�UD��LĒ�&�l;ie0�[Ga#Y23`�!�r��7��@������	.��,Xt���z�=��ke��p�'�\X ����Fb@��Ä
E��g�r)r�Ugk{u%� M8�����w5=���r�G�݄̀�dyx�Ea��ֲe�=\��lt_l��t ���dz�@��<���nǬf��Fjx���T�{�qp�� ���ӳ�M�9���\<h�\�*A����ޖ��v�"�-w.�X8Ɉأ{g�UN�n��u]҇����{�N��eys /�ȍ�\I�ot�{�Vi&��a/%�i�h/�Y����t��?=}w��z��R��5;%Ϊ��.@թc�KS,��dHS*d�� �r�oW�"��ms�6�z��ݎ��aoA��z@���b�̀3 Q̄�¡T�X����Ax�O��y��Q�/���9�����0P�Im�D��d/s���7r�l[������ӏ/kA/#ِ(�@(�����c�bw��P�E�OM�_Hl.}f��f{��a����
�ߜ\�B���!b�C��,	d�y�}f���0��f��5�3
?z�����E���
��4Eꤽ�-U��?:Ar��w�8��KL�ᾪ�т#��{W�Ԉ3�����}\�v��N��ΒV����4U��<���E8K���6����zz�^k��������'7�K��J�稗cwq�k�JX���WJSӫf��3N	44�36�]�N�����K5��W�,eڱy�\h��u�ʸ�N�zcL³
���-I��*&��էE,�H|��o�s5�@H�bX�;D���V���(l�j���'+p��vh���r�r>�.?uov�˄W+JB��29E�l܇�]h�5�7:�o��4��{�j�E�o���T��CV|Ep����nԠ�4֒ސ��V�.wgrDI.Ke�^���E�oy�d�xEϭ���J�o�P5G��6j���|v@�my�Q0�C�u>N+�rP�40tU������m]ޟ`�AM�[�^̙xh��6� W��a�8�C"�bcU���%F�
�*��̤Y6�&"�$;5��nf��#T-���3$��[���u�g`������j#c�^��J�Xn�q]{U۟+���;�A݉�Cq�!t����mNF���mܦ�R'C��D���tz=8��RL-���Vz7K٫�+��:8,הocނ����m]y�2f��T/r�ʏ*K��m�}E�����d�It患 H2!"��^nr��m�5�鹹�����ۛ���˦�:Z��v-9oٷ��6�QEp���Q�����=ѵʹ�U~��6-��V��[}�j�m�ű����W"��u�\֋���F*6/�sT�m�_�}��}����KF򫕹r���ƍcW-�Z*�o���Q���QOv�*��k��K�\�)��nTU}6����[�KWMk�͠�5������I�W6�r��W��t��sr�s��m�t=�������{49.�Nl̳Y�i\C���3[b���ȶ�R�Eí�Z�����l/8)�ݮ,���G�0�Xip0��j���t&Z��Q��ۘ�܍�Y�ɖ�Y�؍A&%t�7�( ��8i�ૹZ�&�@ױ\cY�)U��k�Fm�
�X╠m2�	R޶�\�ٵ�c@3dMK,#R	s�F�������"�6�jWhM]H���j��Q�k �`�b,���iGV7i�Z��N��`�*��X �;$1P6�LĮ��0�%75�[��;���+X���K	CZ����u�HQ�#^i6�mB�9q�gL�k��hܽkR!�#�)ac�m1m�.��i*���EƴB8iBq��y��k81��In-��v�m&��X��hW Ɛ��J1����&���A�K�%�e����mbG��k�;�4t!��͊g1�1�V�E��#�-Q=�K���%�J:%
bRٮ��;J#kY�. �c2�F]�`ޯ&�v�
�f�����<��CK[�ae�c4y�1�(muMJ$q	�SDU.;l8R� �s�+
�����,5X�kiʅi �s���m1�nlb�&�l��C�,�����!m�����XîGL�қ.)u:3Wl�%��%�˛�`0��m
]l��%A�]*�Ya�5̊�E��%:�ej���ZT�G.s�X��u�sC�2�Q43��[ Ybf0v��I�i��)�R�[`����K��Z�A�M�#n� aW
G�ff-e�
�D��b��y�[\���bFj䠲�4m��8a3ن���asņ,*�^�8VZ�m���2�*������q�f��-�P�YYK��ZՍv�,�o0�2r�t+\[j�f�����!��x��A�Xia���0f1[��CD�av�a�\����sd�|p<5<n2ZkWp������a�4��ΌZ�V��(㴦j ���7K4k ��œYu�����nU30��7l]���.@Jif[CK�6 4Aj�U�{Xy��y������H~��ö-
nd�&���K�XKDmc�.����~ї������s!b<�V�"��a/B���QdC���!��㘂9�dP����3ͳ���|�~u8�~��R��=�]0������A�*B��2���B�̀3(/f ����]�&UNE���.�2&8K���#��2��Ht��a���H	��H~�%��{-s�����/%��X��Q9Cj������dQ�2<��#{��R��b5�|ӛ����f��J=� ���d 9�+9>=7��R�(8����S-]-�l(�t�$��W`oh����m�����5Fb�12f�67�o�\ه�.��stV���J����k�!x�ā�̀���O�t�{H�MU�xύ����YB;������������u��X�lu�#��f����ٲf&�\-UU��/���#�D��*����i��i� �A�}�r�$j�^���9p�}{����'2N⽼�/����C��Hإ�{` A���dz���#1!-��؞�L�ycAx����JQR��wNJ۸Ș�':!��G���Pmc >?I,P��%�26dȾ��F�~�B�;�x����+�rӏk�@����A��kX��>���~	�0\AsGd&�XR�����-�,���V`(9!3&fk�=��B ��̄A9��m����7��4)r&(�U+��=�����%�R�͚�ܼeg8�����X����;�lÇ�*����b�B�Ѵp��da����A�Ay�G,�g��^U�b��冶���0�8&t�.�OWZ�D�F�y{�0��u�sC7\�$��c��/p>�6�t��ky�U�tKz2pVm�#Ư���_y]��#\Fb^9�#���;p/`�f<���~�!\�f$���՗H�U{��A�Jp0�� �A3^̄f ��p�h�щ�w�X�Dٽ{�im�dLq�l"b�B ��b��]SY�e�LG0�n��M{0fqRƚ+n/؉�"�UY���lA��̄Fdc�v����4��!��.j0�{Y�ّ@�R=��q�ݡS�b��6�gf8����(Х�����̃s�D.���������A����+���Z��b4Ko�jm��� �����B ��B#1yz���ܳjmG�� �1��-�@��7>JN�W�nc\� ��

ͣUZ�nA���XK�ۺyG{������k*��n�)S/Ӻ��v/��Z�U����!���G2�D��9�7wQ5�6��Z����rDN�xv] ��
�"��]Hn�Ic{U���:<��fO�)�0!DJ%v�lZ����a-{f�$Tɕ3
XOW���Z2�^#13 �]���\�|(>�Zk	EB��.��СR�!T�=[ܔ��o@�l?'�J׮f�9�n|� Aw�9�2u�.�#{w�t��b���!R+�����A��#����MW)�9]0k���݀�"�s#�1́{]N��������ԼFb
fL�Ow�M*�9��6$(y-u�^3Q�oaP����"�T�.�46��`��¾؜������%�]� ���́W!n�K�sg6�V\�G1��A�˰�n&�'>Za�aRF[���Kո{�fTvɽVp��)�"�fGX��n�����濚��R!p��J.55��Ź����MV�iLA�$&v':bV��c)Zv&%bV�:[4&��j���E�--���Tn[� #5�h�Y����U2V�M��c�m�G]�bM��K��jv�8`:ٛm��]�Kjh��� �R5JsjP6��7�B�֊찄ۚL�>�}!LQ 
�f����dtѢ�n��ݥ=�лE
�S$�}��ڄA@�B�{��n�^w�lE@�.GU A�B�q����*�ءl�[�g���1H���%%
)���*v�E�^�؂2���{bn���݀�9�.�7B�����\����+X�t�_i��\�.�����f/fE�����6��/Nd!w;��%��qv����p8�R]A!.���"�P� �Bf ��qf{r�a��\��J2���\�g"��kab�B �ȿ}|��>>��0�	}f1h�k��$ٸ�b8&8& )(^SfR�������FdS۩�[�`�ley.C��΋��	����A�D[�,��ȣ��^#��5�@�G.�W�bi[��/��(G�����J����q�9�+�b�r�b"5��/eVAɬ��זQ�	�(��X?^1�˄A������p��^�i���wt�:����t�� d#�n��KA��Ib�>]q˞��K&�'W���م��\��=,_�!��Ct$!vC���M.��@����U;��u�fc��B��n"f&���^u�ߗ���dW�>9��	��B��_/P@W�ݽ{]�4���f�/��qC��H~�,+"�8�/Ϛ��l��h�v�����B�
f6�q*���ԩ��@�P�̀��Kِ�F"��޿��?M�Vs����9b��x� ��Bf/ NdD�5Yb��B t����̌�B������	̚w~�#~��Я��`T�9��؊5�T��g�P����EN��㧽�ޥ���r�׍�q��wV�D�z��.�D��{��l���v旵=��s�6"�|w`"�A�s�����v{W���0n#���/T�}�<"k.2.8��o本�|��A����ۏfW���(S�.�02h{��^�8b�T����H�E����s7B����������7�^C��~>�R��Q�2�Zh-1.2H��D����-ƯhPrJ�����B�f��o_��Hl�E��!�6"�%.�Ȕ���,u��/a�3�D!妥��4�Pr����k:�o.	dy<(P���q��j]("��ڐ>:�"3 _�!�BB/;�
Ⳕ���s�^���߬P��iC�X���Ws}�  � �/ax�s!��Օ]����|�`")Tm�s��3��135gK�Tz.`����re��Z�%�V�{���~);`�8��W`ۏ_az]��̱7�.	���c��=���Hs!x��'�'�7�6����A{d(��sz�]N\�\pkax�؂9�� ���p�������K	FbfQa J&�T�֦��Y�K�$�"&�2����,�	�ݘ����Vy�>�/ޛ�>��5�߅��3�8p柳�`P{Y�#��d F(��Q���nFn��z��[���plE�۰"�s!�تn/3l�¥E4 �������l���4i�ܞ7p��{�G2�>9��� *h�EiA���������!q%��}Y�n���rǮG>���^K^^���}!�%�!���0��ը��vm}�	݀�E��dQ1Hv�)�3c8�^`g����lߒ�^X�t�=�[�CNF⼛��Li���4�	ED�u�PKc	�Na� g�Z�p6�LK����ٍ�R�C����q�k���)��Tܜ#���Qe:�`Ebn��],N���ubm��C0�.1X��ah��%�Q�f�n�1��mҚ�+6�B\Q��̥�[��K��"9�ŷ*�D��s.+��5�[ ��a&2�n��)�J[G`����W,!̱�߿o܃��e kC:�[����ȇ&�&����	*d�38G���k�3)x� �B�����7Yw�;��f���A�Aq�d7�	/�Rb����*����(`���רR舾����f��r�����ʮȔMcMZ^Bq������Hl
R���K��r�W�����wLG���ol]Hn�	,]	,����g
رBm�HE��g��yw�˺Y'6!�b�@�z�ˠ�����2 C1s"W �*^H�몷�!�$ę��&������P�m�f%㘅�;���8�="!"�
H�0��Rcr9&�0fd-��HZb�˴�2�W��=�q~��!���/>W��^�ۦ��Q��=X��/��HEВ�P��zCzG+��v�ʣH��+^�������ljŌ���f�GO���f�Q�DNw��u�Wg�:߂���/�!(jS}?-Ό˕�Q�^�;^9�-�ܵ����]ǯ�Q̀�G2I`�ǆ��#�z�3S|��K�=^���Fdy�̄Ei�uVθ�U�@�BN��v�b��h����wr�Ff�w#��Dhf�"�3(!U!�B��������}���jn���˅P�[����b�7B�HB_K>�}z�;�4J��V�4tL��6���YF�����#$��SB7P>;P#6=�9�/T�ZWgGoS�5^J=#g�tQ�ؿGr��嘂9�dQ�������"	ͅ���'�v�E��@��v/�R�גs�Wwb�i�$?),g�����
��O�7?e��Z��VYa�-��cT7*:����g"���cbqC��ɼ��In��Uy%"u���v����ٝ϶%3���R#��Ym_%�#�ܽ��4�e���,joK�Ϝb��WZ6gl���`�L���mc��t�}��C�94�}���Yt�]��l�>UݗÃ�N�-Wi݀����V�;�r�,}�9��ͅ���I�ׯ�F�|n�x�܁�׃{�����u3.O��teazgQ�(��W�8�l�K�<��c]��i�ӑ2�mG��x���i.C�{Uբ�\�L+����pgĿ�����_\�39f�tvIڵ{ǂ2�r�ͅ孧\$�u�DvH��F��4��k�j��]6ϐu*ɱa��av�YG�b�J���f0	��hޕw"{4��I�j2�%cr��J�l�ۻ�Q�0Ф�q]�zs3N�����ѷ{�$&C�>�D��
;�]ޜM.p-��f��ظ�:�S���7Z��~��m��j7��`�=.��5<�l��J�#�n�����z��l�>{�6�qښ�f���Ѯ�c&k�3��e�[�gǻ*�U]	�AX�8����m�4+��P�k�I�s�F+�G6h'�fC����o�זl��9e\{B7��K��j��3�v����ƣd�l�P�n�f�Ɖ�d�����ۚ_�t���X�R�'<��ĉ��[�]Σ%~��������@��I$Ow1*����I�Ş�]����^_��jM��C\�ĉ H�Q$�5""N�dgK��{�Bb۠h��e.��Q��B{�#{�);�bu�f�1)d��� /�p����;���G;#%nt�7-ԅM�s(��]$���΄��dD׻�n݀
�s�H��d�T�.t,�����y��șo9���e�6�\�^W�{��ۼ�K�snN���Ӻ�+���s��3�V����^_�k��^\�_���ۛcp����Xۚ�o{��v�/�͍\�lV���汱��Zj�,T��X�,h�j�-���Uy��;\֋F7��[�nQd�~wU}76���Ս�k�U��nsX�Q^Z�屯�^k�h��^�O���4����Ό��qQ����#�=�����L1P�p�u�@�b����ū��{z����\�7Ё
����``���/�9��A9���9�V�}2�l@+aCǖ�'�s֋�/=��A�A s!��TȨŖ=���Pe�1u�qM���QGZ�,R-͖���V���A��8�DfG�b�%r��/s�/%\Tz��<�ն�v�@��>9�e�8��������ty܂;w;�;z���z7Ј#�3r�IUi���H oax��"3 *��
���^�y����]��>ޗZ1w���^ ���d"b�&&�7���_T�U�q� ���x� h�ڬ㹜�ܫ���S���]N�7�J#� �����:��
iȈ�u/qE�0f�8=uע�f驙)T��&��9;��P��}��������	�RP�%��E",���/Ha�%L�~��_��(S�����K�f �$��UI���*<(�a:`���Ķ�-1�������¬�S/��,���|���ِ�m����29�"�.�swYqAt��m�!T$"�HEԇ엻u/	�(j?l!���?Mߞ�E�+v ��s loiq����H�/��.�6(HB7=�ԖjD�9�3�ՕUU�\ �B��Kِ̄D�6nX.�Κ�3"�v����9ިы���*��E1|�e{v(+��Eb�Hn��	,�i=��>�A@}7�O�����Tp �q�|�9�R�Ok�G�y��O�����*�W��g���z�֦���s�B��Q�r�Rɶ��+���Lĕ�л,/[��D�gLTQ�$hda+�%&�	B ��S1K�Ի��e�!h���4�j�6��7j����P�cttܻ&��X��hC��.�mʎ��ZZ2��é|��ж��t��lr8eʰ5�v�h�3\bf�Ƽ�1�����(؜�X���giiC]�ϖ~�~��a��ҙ���ō�t��9�Mѩǔ�2�d��;j�dQ�1	s�xZz�*�kй9�tfl�OE]����B��G�хmu̎����}�����>��xK#�V�(H~��������H�����f!=�7�t>}Z�M�*���'\ A�/��А�@�i��T(Eb�a�@� �����;]5*����Q����L�CU�S��C�Щ/����h͍<��n�,�.9֨ы�������%�	�����,�+���l�&�HD�i�m�v�Xе�c�. �9j�����p�Z����@�Qs|ʸ��<���8�l����̈́A��n���B�ڊoB��+�n3G�i�`)��th��F�q���aS[1ۏ��d�*��Z��>���;�o�c:v̹�s��.]~�|���Azv�����|jx�^��<�DfQ�p."k0�b�$n���	�����f�;-��^�� ���b�B ��e&��\�d�z�h Fb�1no�^�w7�UEǻ�\"Y�v���M*���Iw�]
�K*BUw8������u���
�Wyo����@����CeM��কG�Д$	R�6�"4])6��7[X��hM���l_�ν�����y�y
�uC�մ�5&1w���3�fe��a�B�%�b�Ct-�yf��J�fŐ�/h!U�qz��iU �Ǖ�ȍڝ��N�.d ^BsH� ,�̄A�Cl؁F)qf��:!0`R\|ҩ'۵Q7Q*�X�Ӝ�
ڼgV����*��x���Z9=�&����]ln�B�W�|��y��̏/f �̄Qq�!t���3� sa A2*)�Z�����I�\��}�z���@�B �Ax���B�f ��=�ě��aG'�;�6iw3����Ҧ28�oc���#��db]G���KDu�FIG&$Ĩ�1�P[���n�A(�5r֤�21���z���ߞ�,�����c<�;8n�{��}d��LY�tj�ې8������G�̄E;���^�s`Ș�-oM;wӚ���_@@���@��Ee[yӤM��k���@�b����bux��wN�;�G^>�0�P�|~~!
��u!��HA<��X�@����9Ј́;1�b=�-)�@�}�eS�64O	�����q��:c̆���,\d�������̫K���J�]yk�h8eէ��9Ǘ�{2(�2=�̅�VO����N~��j�����.�E����C���|,���w��`�t32���e-�R�ዋ)n.k3Q-%�R�WOw<�;��2���A���!���2a����	��3������P��?H���)����k}U���j!���=�1)�^��kA3,u���1�I�`-!
�~�N�!T���B�>�dQV�w'R���jLb��:^@@�B � ��HJ�W:��<frE�F�;�^̀�-3x[�-]�������@s8��4���j��f ���^̊����JnV[-�ˎ%>Q�A�@�^�^�١�+��wvLqD��UJz��^�\tPJ嵁�w����N�ٜ�ˏ_]��"��cWҥV��6��76[d~7��'��hU����Bܵ�@{ih���aeV`it�CR�.-��Eb��1R̸�Ҹ��P�.�1\gi��tڹ]�]�'"ޚ�d���mc���3����	]X���L����iqm���3l���T4
ۜ��uԙ��dJ�� �i�F���*Չ�ll^&�+��߿�lY1�fh�ݙ��K�ũ.�u��7-4�*d����|g�˵dy�
����R�_CԘ����r9�c �y�z�b���dQP5y���Gr^;�!ˌ�23*�L���A;��|��̄ޕ]~^3Ј�Hp�̀�̏f@��8����i�F�%>+� ��h	�	,X�и`�Qņz��B�m��n�dR����QM�=K.��t�۷���
Qt��o! F��3@���d
#2�^����q�x͠�39�#�ī�2�Ǹ�B �/fG��2&���y����=K�y[	�c�sb`k{Rggi��8rcMjJ��<�fT̂��=3�ّ@�3�&29���
|W �t����^w@DoX�}%��B�]�Fz��'^ik[O�����&�(y�J;��q��>��w*}g9�l�)K]� ��,n�>9�zY���s�C�O��PE~��'�<�|�\�:#2�̍��OrA({<��Y���1.���YgFf�7��ʇ}����Gِ�FbL�e��a�Sװ4-�@�� ���Q���F7�B��oa71ʠ�76Mt�!��͏ ;PG2T��P��ԇ�F1|kQu�u�1�V�X1p@��s^9��A�C�N�<	�'�ׯ�k�	u��4�؂AK�#�[�Ba�,2Q�U2bfT͌�@��@�9����ِ��k1v�]�(q�o��YI^�2A�A�@��x���7p���E��W��e{j �z��c<��NDϊ��Ⱥ�_�$췬vm,�q���S��*��!7c7�W�>��m�H��^��K�c7 �;.�6��)�&�E	J+Mn+��ϭX]y�B�_�O�ל/��9j:No��LE�': � �̄#1�A���Lnr
�.<��;c�16sZY��Uv���;������Ⱦ��8~��Rb�}%��4�n��lXi���Ll�NEO����B�Z���d4ƹ���f*�c҈غ&ڥf�G8�2�r��";P��Xk]���QB�O�����!���z��N^;�z
!�����ʘ}�=A�D�#29��Gܖ҈萈�Kǹ��ۮ�]�(q���ؽ���U=�}ei�"��
�"�
����B���@���R�:�.|Tr�����<s#���l:�R��Mu� ��TR�{�̜�w��~|G�nzo�Fr'�L&��tA^"TtI�k�]�Q2`�4m-x\c����;�u��o9ֺ�j}�U�����g��~!�=A���9��A�ύHσM|���+�t���Uv���k�쀼s#ˡ��~_^���^���5*��ګ���U��6
���v)(db��l;�~{�xFY>1�߱�� �z��z�_E�ϊ���W�'���G��2;���/�Gّ�6�n6��F�<�ͅQ�z�o*v�7Rb+��;�1dj�|��&�T�{Y�"3#��;��hܛ��j{;��Ҕ8�A:�x�/�@�Dd/���&
r���A����f@AN�Օ��f�\����^!�:EF�7cِ8T��W�!�BHW���T�������t�*���I�P8�@D��ȯ� ���z�
"�d1�kl�cO�C���g2C�V��Fo%�I�'ep�v�H��r�<�W�&��NA���Q�E����w6��)�C���f��٫�*���e}��W��hiֺ��q}Z��/SRS*�4��ҩ���CUVb��b�DKͽ����u�]����v��c�^m�q��^����G���y�;��uϞ(�/1& �A��naʼʵ8��U�����;�}S+{�P��bǘ�݃�`��U��P�o1Y���:]m�����	(�ʪ̏���,K�&f�=�ںb^_r�G��d���q�Y1V��ĩ�TÍ;1.BS�,�����54��qC;	�����_R62e
�p�&k��F�,A�(<Λ��T$���]��I�9���,Պ�iz��n�F�whoݹx��\ՔFX4�*�YB�7:�iB�*P�[�J.]ѯQ�C��f���u�v��"�*,+��H�H)S�2Jp�Mi1O�*�ݧ���g�
9S��"����wY�v=����흑���rˡ���-��{�w���q�{�A�\7y�[7V�#l�*��Z4r��nk�=�U����jL�xw�+�cSK�[W�Z �匎�Y)A˜�8�#�vY92�����f퓂�%#�����r��*�����xi���
䲹¹��i�� �$��NTU��"�X�h�%slTr��msE�cѬW��cU�6�%��Ouʹj5���6��lh��MW��*����5o����X�QWҹ
1_}o1��6*�|Z�6���W���|�i��
*�o��1h�m�Z��D��6��Z�nmE��+�w�m|k�nj�.Y(�����v�[�܍cݱ�+sc[���.I�kzH@'@���>�_��k6��&ƕ�Sb(䖠Xja��,Y�BQ�T�P�f�P��;%���5Z;����ѽ�	q,)[G�.���kZB���h�Z���4�|���C.Pi�z��sf��eα���̦��ش�dl�AV��2(��.5��f��T��!E� ݜ����Գ5t�@�H�)��u��b!u�� PɊ�D�;X�W���cM���T�Yv�)3cUf��m����v�*��ԃr)l"��m�6��C.�������It��6C'(r�Uu��X��VUa�ф��A�4p��-��7F�h�j�ۨ�1M��ki�uz��PXkԆ�yw9�A��rViX�e�Y���-��aZ�a�-Rݩ�v�����En�kn�QeE-{5c df���r8k�TZ6���F��̱�j���6t]n����\���P6�\DW15 MsL]�2�fuэЃr�(���h���]�N#霖�\��&.�yJ��K3����IP�K0J��۵j��a5��ᮚ�Q�ٳ�	�Y���u��k�SYcR�R����J��*�k�a���Z4��e&�aVS/�拜ef�A�bi���bW&�328�\����@��VXҫG]ݕ��9k$���5�k���Q���Z��� ���A����mkk+]�kD*��3M�=�*�&�s��RW5�/,%����$nD%�c.su�j]�4��ca23*q�v(MvQ�֔����4Ճ�Z�P\���)��(JZ�%%u����m(ٚl4����:8�Ze6aX͜���.V�vUUU[@\iq.F��/[���k2i�vR��CoھoOz����k\�J��[)��ՈB@���[.�c�,\�l��3Y�7+d00�)�R鑶W�R6�R�9�ڴ����V���!x�.�
a5,�p��Yv]Xܚ0G3;�D#5��m��m��GZ������R�bp�Ps�k���6+Jh̚ш�1�퍋Ʃ�������A��&bk�]�;GYu,E�䥚��mMFusvUP;ɏ�f�Df%㘂��6_m㚮e(q����/fƭ��1dԂ�<�̏fP@��=��gMD{n0}��S'r�����Q�� �k�@��͚��ѻ��A�D�����̏/�.Έ�J�w�U���n��*����D�e!qE'H�	�����嘂������%��)C�p/aNx�\B7��/k��Hs /@�AxȓC�r��5�]��r�u����y�#\�K�1
��6ϟo��xy^��^I��E0Qt��,]���������,��32��FOG�� �d#��B���U���ݔ�W!�}�0M���L��<^�#2 ̤	̄��<��.ʃ��^�@�R�0�ܻ*�Q���U4�+����²�Jr�buẳ7S.\j��WOu�)yvf��%_��#�܂��A�����t�
P���/v �s"��� ��h K��������d�'0�{y�J��Td�G A����@/��9��8�S��n໏[��m���B�k�eZ���LEr�tF�P̥�/��ǖ�ex/fG�b3c+FS���������[YZ�9����zX�R$-�ض͔�N�]P7�&2WXB�W2jk�`6Δ�Q�W<$�ǔ��g��4�>ms!sU..;1��m����C�c�x��Va[�*�(���㘂9�� �B#jnND-��E7����B���U��Ż)���E��d-y�i���a�����"���^^>�C�OV�S{4*�*����^���畛�tk�9�F���{�a�.ŝ��b��ʦM�F$e��6�ﶥ�A9T4�M�uf_Q�)C����@��/ꐁ!T$!�hb��

_�BB�g���s�Y��Y�?o/q"�5=�w5��s!x�s!x���̌rC/���mO���.�/��+�Q����D3D͇(%3Y��X�A��Lhf楱/*93���Ŗ8��yM�����}`�������%��c�:��G�����P፲%�Oi���w$?7�� 'O:j�oq��bA�C��)u��em����\��}��y�k��Nn��ms�M�"�A� fAQS}f�۝����r�v�� Ol��_HP�RX+w�4w�����WӬ��Ł�P�[쑮�CvaiW:�r��k���M�����:��s���^�Q�R$���]�˶ig�3����f�kT{�5�䑸O»����$��HE�BB.�>��9/r�	h /6./�ie�e���s�����Fb���u�Tpʁ�H���)fɜed
��Z�Í6��2�6˃�ߒ�c%��� s!xNd*w{7�}�q�I�\Ȥ��}K�#uq���A�s#܅���� ����Bk�k����|n�� ��_ �̄�-�=Ȱ��^#� Aހ�^̊#2���h�����{��O���9Ё�^#1/��2�y���t{f�^=Ј �B���q�λ��LR�	퀼FFl���Z��qV�����"r$�"�uK���/M �v��S�ś��T\p ��T���@�ȶӓ݋.X!��a�zgݯwfE׊���j=��L�Xq�^:��%�̋+q��r��Q5s�힩��'B��t�_��m>�P*D�ql���h0�%ΆK��50���c�\SX�ha��jG���XJ��Xk�����1�b�Yy��������U�4���Ѻh�1	2�Q�;6R�氰�ѵc��k�*LMf�B�u !t�7\���a��%3aj�J0i`ñT��6Zk�9�Q��3�퍸�:��={���Ϻ
4\�����b��+[kc�ܭ�;0ҕ�M�b�?����x��dO�p��SG�����Q���RxefW �E3���Ax��'ŵ��%�S�2;Z�#5{��7�^�_e��w�1K��lFsBKq<uYUQ\��ݹ�A{Mغ���n�h7ƙ�����I��z�%E���O�9p�%����A�̭ȫ��S�F�^{A�h)��q�ge�TZ����@	غ����dn�Ϗ���p��mH!��q�5��[^��U����}W�b�/v�D�>n/�6�W�r�莓NI0����(�H�M�Kmn�pE(�J�7�.�������y���ϗ���7u�ۤ^[~�K}��3�Q����xQ����jH#�q� ���;��f=~+ޛR�/d̥�\9,�b����)�)�f�>�	��]Bݞ��#�IU.�SnAJ����b�u�Q�H����U#���
���j�^�E���;ǜ"h"uSo������O��E�"�)כ������=�S����.���{W���{` A�r$�^mCm
���{F��DV�f�D<r'Ŵ"n���g\c�Q**=�^�lS�G��Ջɬ��G� ��@�p͹[��S�`�
b��D-��診�= �q�p+�6ץ�*Q��O>|�����6�Ѯ�c�{4b����%ԑ���fY]���5��fT�dp ��S��n �ګ5�[��b���@���;��ӧ��r$�&�D6�H ���'i�ެ]X���
�sj�쵛��U(��Ú�p�)��B+�4����`"nD������ ����&��]8��y�'�#"�,X�[z�+�(��a�^%�`�{{(v�0񙼃������� ��J���7��C��΋���S�8D�@��}>-��[�P��̅�p��[jn���}��[j�d=��LJu�
��nF���m�7A�h"wf+����܂��|�)�Z��q** �k��h [�AVk��g���@��(Z���$�T�1 H�,Ѝ��\B��R�mf$�d��S2@~3����%����T��tMV�˙��#�RU�7\Aڎh �����q�mI�d2�R�Nf��;���=��mP�� OlE�^n3au���";�	=���n�T�ꮇ�f�DW�fw2p�Gk�>#�q�m�!�{�=9T��A�>΋�^*y�#U����L�8�vƨq�qkz���d�	�Gb�_��>R��T��\M��	��T�B)��n&�T٣��-[�n�j٭mQS���έѝ�s2�ff[�2��g�n��q�aDZŘvm�/�ڸ�j�d� ��Ȓ� A�������ߟ�����q��3��Y���s�)�&M������2:H��3��^�� �Aۙ�m������=s
"����i�2-a��B͵���� �Bl��3��H!�(R��ºo�K��LO	ǜyc@6�̈�`��"�� s5H7 [��-���s{�*^�C}W��Fr���#�� ��Ak��F�P���;���g��^�7s��ρ�REL���y�����Hn���Ȓ�T���c��K�� ��W����.f|fW�#�-��m����>�i����^�&�Ne�p�­[B�\��j۳v����9���(��o-��F�z�#������WMCޘ�#β�4�6�T.���Q�i)m��T��b�I�u+_�^�a'����$f��,��+mظN�.Ȣ5��n��ذ�u�FUل��ºP)u{K���ؖ�XZ�j͎�<�lt�eZ��%��&h̔v�!�h�łj$+iթt%9̸�7a+��̪�R.K����~��ii�������Km�v�P-&�Q�[�[54#�O��9��w�p,���V�\���͛�z�C���w��׸��@�����-�w ���X�{��p�pq��%���B.��獮������H<�@�`�F�`�Ԃ�w@�n<��fvnwfen�O���g�3�H#Ƕ�n!�3���q@�rK템���@�G�m�/3�;�Y�P��ݰ�!��N�H�k�}܂���7���D6��i��6Ї��b��k�aDl{����p/ŸD[j��r�98z�bA�h�kB
@R��kD` �, �_���̽~Y�>n���t&�����e�n�z&C��3��1�F��g��A� |�RF��Ǚ\�Ҭ%�)�9,��R�QVB�XA����-ź3(��*��Lּ�R�%�
g2�x�1�����~�>�U�Ӭcn�nb^��;Ƕ��In�]Ɂ;b�khI��m�����
*�`ՋA�fVu\�t����Q n����n ��RCip��Y�~ysH>w"An<�h!B���S��^ݎ57FwGUu��&4	����E�D�RCp-��!�yȽ2'��[v��zx�{��7����FsBAn�靬�4��J��WG��ڬ�:iB��d)��ͨ֨)k �s\��}��H ��#v mߧ�͠������o��Qj8�UU�&�{"yҲ�P@�� ��Ԃ��p"7��jWL��j���P.��=�b\Ϧe=Ј#��Q����1<i/^�[� �A�y�Y��,��|��a*֤�X� �˱������d�&�Xq�jgP!��D�[1�:� ��N���b70���k�U��*c�Ks��,��~�.�<G���EB���ү=��Fr�GJ��x��)�N����N�Dxk�捘�lT�G�]�3:$kv"qA8��)㺘�Y3��7v�b��7��:�]\r��䋤�);W�pX��B$6d�*I��(�sM�����#P��#Q�5�A���1!I��E^����*H�p7F���rΚW��週G-�t���LL#;N�E�������t�m�l�f�jE3�y��Xx)�w�vBc�:�@�\�b�
ش���P���d��j��c���vl��!��Ù�k�U&M�W���=8D�5�ʧ��}x-պ��օzfĆ	�*���gc�w'Cuoe䏹-�i��u�b�zsd�:Q�k-��1L/�'V+H��]DbaVۊ�(�&2UF[�z�!ջ'"�O���qQȺ�F�r�缹���LK���.D�.�6q��B�H��#H׻K+�c��v���C�C�[x��L��u��7a��2�;�����}K	��Yʹ8ѱ���U�q�*����ݬ��k�6jdUha	gn��	+y�v��Թצ���U��OMF5�r6�V��/
�J�/!
!��G�o�b���cgu�����wW6�ܫ�lm������+|ksk�F�|]ݺk���͒�X��F�W�s\�/��|[so�tmF�ђ�����ccQwv���w������6�Em�sA��&��э����F�9�nkP[��H�P��-|[��yr0QO��h�}�,X��b��5�n\�w\��(�N뙟]�	��H'Ē.̎��u�1��Dl{�/������D6�D�W�Ah/zפ6�
��oM���]%��'�T��[�j{����k���5$6�� m�7���]g�FG8��]�<;���s>���A�,h݉��ޛ�䞏��{��EɆ�2���	��Xͮ��Va�`@�2aL̦z4�m� �� [� [jENoj�W\æ�F��8n��@d^jq�6�6��A��=U�c;�^��d���g�n��������o��Qj �k�A�-�D��B��`�}�4t�����^!����|C2ÖTv�꥓7B�衁�_	Ng�3�}�X�@��ϛ��n=}���7̞�\E�{�(KmH�y��y�WR�T��� :Ҳ(�Vd�����1:n}kb�o�	��F�3�ʹ3��yg.�b��z���\!��=�.����G3u�����8�B^� ��m���@�1��� ��X���XN�3vmn��t�E�Ov�s��n���G�;X��^OX1i�J�$ƴ�+�+ �:�m-GZ���!���3�#7P�q��P����z�Rs>����E�W�A�j�fl��my�������1��B[�'^���9��g��Ω� 뀼A�ϛ��4U�>�����Dv9A=����D6�|��6k��뎫�m��T�##���H9��p�%���Bʦ51�y\�M��D7P��Z����� �����鱞#�L����� �ץ�n^�=j�Х��Z�g=�k7���R#x |[�|�O�p�-��U�˚̙��VՌlT]wT�Ad�ШM�d�'���w��]6���B�Ns˱z&�ݛүo*��1��E��$�R
�aAbl�Alie���6j�Km���1����ț��qW����4��:���{j8����j[�&�%��*�ru2��Km����K
�n,-��0��6԰Ȯ��l������Y��g\�ь� ��4tZ����Ը���m7"�A�)��	�vQ�݊�9[�mՔ2�����k*�ΏUź��mHC�+eb�.�R���I��2�\�OU����F���m��3z6�_7�1㈰N�`&f4M����l/Am�!���:��JԆ������WV��ï��3�3���@�5����l/5kձ�sT���n���]�*v�T��k^�K�R#x An�"Kq�@6�F�D�Ql�[�z�D<���X
��4��o�^LD8�	�� �����V���3ƶ|��� [��6�H-�mP7B��Q�0N ������ע���C�tysAۑ>-��+����U��H��f"$��%�u��j]]� ʻ �

H��3 �L��q�mM������ܺ�"7���ͺ����a(ky����IHtP�M��:�E�w��F���h�b�]�L���oj=�Q��M�\��a�K�'�8-܍"ޯO��W+r���̓��j�A�E�v4�"�P�3+��@���ۑ%�@���fm2A�%N,��;4Rs>S<${�9�@������D[�&���V*�f��ݏ [i�w�8�kv�j�������"��0��D��6�O���mCm��[3S�$��(%Z�7Z�<��0��w�H �A�����7�=��}�>o^ѿ����],����B�3��ivX�feH��A"fR�#u�� '�"Kp�СJ�l8�٢���B)�n"c�#���O���n�m{O;3Qd.��y�x�=t�g<�Z�F�@�[��#��7c!�wUR����}�6�m�����t�PS�ew*ح�Գ�fC
	o\�J�FE\�L���¯+�T5�g��ގ:�����v�Н�{�k�JA���lO+��{�Is^n(�mI�y1[K`O�7�"A{Ch*7h���)9�L�t"������;�y��^>m�7�p��6���Y����V�9�:�"�� C愖�|�
�ō��
�S��Tvt�b�6�B�R�K2�n�Wb���333(� ���� ۹�p"�����vU�0㈺��뮕T�*v��|�RCk���@��ofA�ѽݸ/�.�9�!B��.�ó�'3��H>=���h��q�������/Kh"�#���'�idc��:mns�u�D>�A���n ���܉�;��Ss�(�-}�>-���������.јq�A�� ���fvjY����,���x��Y*]`5NŻ��R8�=}�tKf���燣h��v������βc�P:�x��)��E�����������r)N��tv�I��fzA=��<�D6�O�h0�h��7�"����4%�]enD�����)��Y�]`���K��n# ��$>��p�A-�!�x�;�G�Z��"�3'}��Ώt)����G�mCnD�[�EH�(�f����n|u���y��M��F��	����-��v�g��r�Gj@�p�[� �mC�}JhD��4�N3���Ϧe=��pmϛ��p���y[kd���r�G�m�����]��]j�~����:G�Cϓ_=>�S�.����An6�m��������1�6��]Y����q����9�E�^>m������3V�5on(��dɤE۸}:+1�LA���PȉZ2L0T�#����wrZ7�4+�y6K�׋��WKHc.3�;����4�\!W2��6�����FcK�ءm�l�E��c+e�P���6�5�w2�f�Q��Va�V)������*�TE�n��uڕ���6�\��r�l�&��U3f��WD�4�Q��4F��j݄%���c�3VՁv5�vb�rڹ4Z��׻�}��R��Д�-Pل�*�S9m2��9L2T̩�9z\ �vȒ� Am
"b�Oq�573��"9�����{9��FwH��@��m�#��s\F%�����i��M�6�.:�l��"���-��s� ���@Wu�A9Ј 6������bt��2k��7R�;r�9=��r�k�Ǩ�כ�F�����쮀�#7gݱd�
�P����{*&�zfzA�����B�GK�7�>��Am�Hmp76B��P�����Mw+�=wZ�lH�́��9n<�	��EnUdS��J�"f1oV��G[Fjf�iYMtԱ�kel�2�]�s�t�V� �Aۑ>-���q��U՛Β9=��V��y�Ҭ���� ��^n�� B��"৅3{bˈ�
����%�e�2j��@�����U�}�r��j�BƝS1 �,��
ݬ����,i�X���ݖ13YHq��#�
�M��]�&�zfP��}�� ���W�i�o5ɠ,��Ƞ}���Apm#�f�o�����{�j�4VĈ| �_9�qd7x�����ͽ��@������kr'�6�
�Nfʮ�|�Qp��{�z�t��s��9p������/[r'Ÿ�����Yƃ�/`������΢nW�g��Ol G8���|[^Û]¯9��*",�3�J��0�%uh��BmZ�u�BM��W-?/�������ڑ����ӕ�+bD8.;�Ulw@X��{������y��Bt(�v�-�����eu־w(���\A�E�<���;���#q�����?[B�b��	ڠ��;��b;�t��� �ף-�w"�+���'�R\�i�^;3:q[��0��9�u�js��nW�g�{a3�/ۙ�q��ӂz�k�Oz)zE��Ǒm�ɦ�����8VĈ|&�F+q�5�e;��>����[�-���{��W]z� ��'������"ڎ�^�h"�y��rE<����$��(�ʉRI�$ � ��KV竬k�S�J2L̥,F�"��p�-��)47�oO:��^��;��}���@��@������&]���ڟf]���vU>�" �7�Ϝ�-�mD�6�Z��du� ��^!��>m{�t\��*+���[�o]�-��	��>#�[�"�S�AZ�̈����|�H-��!�47�oN���^���Ol/��T齫ϫ�0Ї��Du)�6�(��U�B�eJ�yt�7e��cSƽ��%B�J7�x��jr^��]ݘ8��D��^n(�mz@mq����,���8��<����7��#yȐ[����<�����O�}�nt]1�]�e�D�u"\��g0�˗W*�|����q>|�߿k�� �X|�v�<�-�����c��ZZ��@-�$6�����M��~�n���<�&�zf{�	�9�"gqe���ٛ�-^ʊ �sZ�k��Am��y�YypV��V�NE�o "7�[�Cp!�"G+G��5�";�z[A*V�]�O:�j ���%�TF3���GϵI�E��nD��
e�ݖ-@`HRr�����T�J���O�n ��"|N��O����~�H|(�RI		��U��7(���U�~�i{EPv���0�!�%:
��o��t��5����ix�ׄ<#�)�(Aj� �"��(" �� #sDut��N��"��
18�u9-)'4'�èzR���Pz1�-Oer�%-n��S�. ��?yOd�������^v����a�~e��������A���?�κ��:�,/e�P���+��ܔ��~'	�:�UEP�>a��7��@w_�V+ЇԪ���0�����b|	$J[>���k��A���������Q��,3������|À���>�YG��DQT������&a ��O�DlA��ϲ �6�����;������֒��7ʰ8�|���d���_;���-\'̃�pP�*�=N|b��՜F���$>4p� "pQ	��P;	�$P����i�!V|��:4'��f��wG�����>�9�H���C�C���נ>��~�N�'��S����"{�ا_k�8 �������h��������� #H��1�#�b|�)�����P~_j����M�P��M��R�
~ߓ_w��9�?@}A'�^����!���/�_�9�!��'��i� ��>�|H�&|?�`@�A���8���@y�'��5H��*������EP�~���Hv���_�S%	�lv~�(=4�~A8J }��<��Py@��$���[d�Ұ?���d�  ���K���� �x_�g��!��Qh��_9j��A�)����pi��O��9QEP|l?C�a���)� ��3A?#�� ��� �X?������y�=�K���!�>�l����������,�����}o�8��~ ��'�M/y蘚����������q�=����A�(�>��}�(�/��s�	�������6?�>�����Q��'����=��� ZC�|��@�n}Tc�`~�C���z@�:~jx@���$��?y��o��8�k��PQT��A����N��������>z�a��#��DF��<׿��< ����UEP������� ��~��=�K���QT�~��>��@�>�����r�C���>۾T�$� AO�!�J���Q߹�����)�ރP