BZh91AY&SY6���ݔ_�`q���"� ����bBπ           u��%H R����J����
�dh$R�%�T�R�A"���
 �d[�UP�$��Tm���Դ�R٥C{��E
���P�Q R��	H��h�4!B�HP"UJ��E�j�h(fµ�J���  s�J0z�mS[`�mp�)RWT ��j��l��A��HIhm��QTl�����-Q��Ԣ�DՌ�A�)� uT%`  �JP ;�=g��*{n��m{lwj�M���j⨭Qj �3Pf����*���pvOv���מ���U��
U^�IH 7wƷ�%l5^�z"P�%ޕ�a����n�iT�p�� �Ǟ�R�U"���{���*
��z�ZoU�xT���OR��(m�(UHS[l�P��<�  9<��()S���(zOW{ڞ��+�Wt��U +�Wz�� U�O<�*
�K�^p��(1��(;e���ݠ<������TT������	h,�'�%( gϧZ[R��=�JU�AU�O{^U=�����hj�ާ��������=�*n���R�j����
u��ܽ�T�U���CF�@f�	$�	%�@-��I @�Ԫ�������=�곥@*�;��y*� շ����:��@�ܮ�S�Q�]�@���:�]¤t-��:J���PJ�L]n��/�R���P�>����J�
�9��B��u�*����T�4=˳�[f�*n�U*�)s�꒢�<���*��n��= Ǖі�`ф�HDk�(� K� �� (�  ��� �p Q��à�'� �vV+�P�XW@5���)B�X۳�C�@u�|�T���[�8 ��8*���� ` � 1��x �j{� ���op ���;�Z$[QVL��� �נ�>� ��� �`= �À  �� ��: ���(�X jV�`�����m��JE��W��@���: ]w�= ������ ��/x �y^�� <��pPWE�"�\^� ��l|  �JP����  ��2R� ڑ��F  LɈ�C����     5OɐJU @    ��L��R@h@    ��)*P 4     D�a�$�	��24�h�4�#L�����?��O�O�n#��yg�w����� s��m5�7y�ɾ���k���3S+�g�T U�O�m@EO̠ *����~��M�?���?�����>�?�* *���I$���� ��``D��?� 
����������[b~�-�-�lKb�ؖŶF%�m�lR؅�m�l[`��l[`[Ŷ�K`�Ŷ-�m�[���[`� �lR؍�d`�-�[�lB��cb�-�b� �!l�%���
b��-�[�!lB�hJb��	lB�%�Kb[0`��-�[� [b��[�	lBإ�m�)�[�!lإ�m�#�-�`ŶlB�m��!lض�-�[ض�-�[�� �lض�-�[ضŶ-�b�[ضĶ1�l��`�-�b[�lض�-�[ش�@S�-�b�-�lB����
`�Ŷ!l��)�l���-�[ �!l��0`��-���-�a��`�-�[�l�[`�-�l[`�-�lZalZ`���m�[��m�Lb�Ŷlb��S`Ŷ�m�[ �-�m�li�l`Ƙ���-�`���lb� �-�m�lH�b���m�[ؖŶ�m�0-�L[b[�6���m�l`�#ض�-�[ض�-�l[b[0m�[ض�-�[�6��[ �lB�6��-�m�l[b�mLض�-�l`��-�)��i�lKb[�6���,b[ؖ����%�-�l`��6Ķ�m�l�%�i�lK`��6Ķ�-�lb��6�1�-�m�l[b[�6��-�m�lKd`Ŷ�`Ŷ-�m�l[`���Ŷ)l��m�l���m�l[`��6�-�[ �-1�-0`�-�[�-�m�b[��b�-�[ �1-�S�[�b�1b6�m����%�b��-���1�l�%�K`��-��#�)l؍�HĶ [ -�[�0-�S�	lB�%�KaLB�%0Bض���m�0-�Lb�ض��l؊�[b S� �� ���F�
� Bب�[`�lm��1 -��lD`�[�*�����@�*�H�؂���"���
�U�
����� )��lEb�[�"�V�"�B� �-��LP`�[B� 6��*%�-��iP-�l@`�[ت[ [b�lm�-�E� 6�c`lm���E�*6�F�"�`�lPm�-�� �6�V� �؂�[blQm�-�U�
6�F�(�`!L����
�[`+lm�-�@-�-��"�H� � ��V�(� �%�-��lTb�lc-��lEm���-�lA`+l b�lT`�1P��1E�*��P-���U��-��l`��1m�l[`�-�lر��؅��1�lض��	lcŶ!l[`��-�[ض��$e�m�l[`� ��-�l[`Ŷ�m�L-�S�l��`� �-�-�l�b�ضŶ�m�l[b[ ��`�ض���m�l[b�)�lZ`��)l�6��%��K`�-�l��m�lb�6�� �!l[`���m�l[alŶFl`�-�l[b�ض���lK`��6Ķ�-�lK`[ؖ��-�lKb��Ŷ�m�lKb�m%1m�lb�ؖĶ%�m�lKb�-��P?�s��|���y��ݿs�����kz��b(�����dysj	`F�ٺo]�²k;V��wDPc��������t�PIД����fC��̊y3M�u�d�U��+r�iI��m�a����vi�+�*�m��XR��^�����n�ʵ�$nt��Oft��ܵ�O�
�F���֌vu��[
9�ӷz��3N�i��M�
wV�Lʔe9��V]GZ� �J4-����,V5�o6މMс���S����aVj֗m�Ɍ-n�����T#+i�W��m�o]�H��B��*�f
�Ʋ�i4E��E㧬�l���4Tت�L�����,sl���(�u(2m+��m]u	��ubmfa-��%A�D��#��VѫƯqJ7�è4rٺں���;r<o.��a�2X�1 p"�Y���1�g-�8�D���>V,i.��J�e�P�5*S�c۰�65drA�e�@���6r� �A�V]��$95|V�Sq�F�$](E�OV/6wS�V�=�sD��3f �n�H-���*��C`#�EL7J��D\�+n�WR�"m��R�!j���M 04k�Q� Z��ґ�)!pE��iܽ�Qj�f�S˦��Ȗ�-RH�����D2 �Q1B�޴��j��ҫf��{&c�z�� [�RХv����4��S.׭m�q^�HR7W�H�x���U[*C��V�x�J��ua��C�OJ�b��2�z�4�D�� hг�x�c|ՠ�NWm�'�h�-�Z��֙*
��f�T�c�D�mJ����2j�5���7]�ĕ���&��B�t[�E2igׂ̊34�De�L��4,;.aa7��~���+t�@��˕v��r�{F��/f(67
�5�iU��]�-SNV��X­�t(n^ ,���	�f�$:"*����.V[��W#Z�����v^��.�瞺��t����j����DB��\�IfXA����uaK���4���C^�ф\X�f������h�4�ҙb�)�i�f��N9r��J��V�6f+j��T�]��qm��{oj�?�7��F�yy�Y��Q˹X������W ݰ]
�ȷ2l�J��YB�*��%ϰ4�alGn�	�eml�o1[Y�]�,K����4��cK���O3�e�m�܁��f�AV�B�ab
5�%�f�ZT��U[en&�m�L��*M ࠦޒ�˭Ԍ8�ä�m��5Xb(>FV�CX�#�!rgb��jZ5��=�2�,�C3f)�R�7w��K�(�Y[R���!��z�B e=f��i�q�2�m���B��U�",Q��$ou�p�yS���i�=�6YX�6��j���Uf����9B�����H
�@j���N5�%�k^%M*Y�|�3�t�hvgcS9M���L�Js^��5'�_��R;9kέ�]梲��S#
28�:�i;#̕o��ٷgEҒ )���%�;�(H�SI�4^�'�������Yw/F�X��EY
�;���k9b��7������f:a�u䛇XX��K[�ũ�StC�&U�L�4&��L�܉U�5�6��P��x� �{���1�Rf#B���LN�l�5u�YHЩ�I���n�f"�ͼn�OG�B�g04$0]�d�u�R�uwr�Խ����P�.�Kr��:A���UAC	�;�ͺ0Lt�	��5�(^TXv��۽�j���)R9&�7JR���S��V�	YbK�-�+^V1����F���P�M�X�5��B�J�*N�h������Ҹ%J�������0L���$&l�Mm���x%��)��T(F�b�v�Tmm
��#�Nf�-0�Ի��RT�ǭթ������*��ʹSi�W����+T�*�^9�8��sfVP�������ҵ[��p�7wO,+��]�"30��!�V& �zP�פ%�G�� l��ZfM��ni���jM)�^��EY50YɦI�m�R�N�2֫4^ܱ!f�8w#�z�D0�㥢�f;m�p8cěLu�X+;u\=h�oD��c��u�i�г%<	�3o(�f����*�����dӧ"��f��0O���Q��T�M�y6;���+HT/Hf)-e�28L[z7/5*�u�7Q.Â�%鹗z�JV
�W����挬�5)���,ʎ����Rf���(��GC*�g34�3Yˬۦ=���m�J��T��F�;Ej�����:�/r��y���Ro4��JJ�ovi�7o(A�YF(v�7h��r������4S8�Ӕ�&�^رq�b�����q��o'Jۉ�Ek2�ְ�i�V�&�ɢ,&���X��N�Ŷ [O/h��r��q�b�h=�.�IQ�x#˸�RH�,�ҁ� �2��{Rܫ�]�4�) ��%�6�xo�g`����b��$C�6�!�y��O]�;��-7o[
�2��@S6�[��[Z�)9�fU���R�;�n��Z�h��yN�5L�źYv�������Z�Xv�=6� �X�/6Ԃ5�����
��HS�:�Ea�W,] :�V�7Cs�n��+B2�e�E%2�H7Ch���=�9�B�ǭY�B�5����t�E,T��ݐ�voY�6�L���wK6��m^n���]!I��Tb�T0�OSX�n1��hc���0�6ÕX�W5CGH��%C37,�ܫhhm�m^ʽ4o4�Rg��0��KF��m;T���NrPAb�X�Eh�U+e3���c�!Vc����q�/Z5m�Y4+`�N�;��gP�i�v��v�wm�ۉq�&�Y	�9#�a�MN4Y�SU����Z�C��C��w!�śjGuY�h8	��ma�� �Y��M����l͖��EX���������+���	W[nD��vd��.	W�:����.�A5A����9[n��[� 32�R�����Y&*�ҀT�^��5,"R��F5],{��u&:F\�t�1A�,�d�H�K]1�:�R�j�2��hdȥQ�
�n�Xy�x�#�E4�����36�ͣ�4t��wcr���,��Q�D\�
���q]��1�xp�<�6ؓ2],�k%�`bX�)�;�z��ն��eZ&�k>�Y�;�l$���R��[���12�̵���%�b���Ck&V��yIbR,:��5[�+.�hr��6�\mUJHL:�[Tu�wbYZ ֦�y�-t�\:�Y�6Qb��wv�ˀ��Ї�u[���sP]%��UJV��.Q+��E�Zmm����&#P�N�m*�2�{#RKͰљ�&I{[���S��2 �u���eL���ԭ����r��I�fJӒ���'�}id�E%�&��5Vց�J��)��Ѱ&�d�1'fXl*7���Mt� w����+V��	d?�)22j�6��n��;����D����]�)��!���Fl������̔�y���ăYu~gV�1�E%L-�.B��n�����=��,�/w�2�Ͷ�3���l9�%��A���P!Ǉ.#���q�>hm`��ɣowL(z���◡�Bf�@�%���6믻�#���F�i��+�ow�=*ݳ�b�25)�wHe\O$i���a�:yb����&�m�hI���\Z��X�_S�5�J����E��J5h�] n�Ű�,x5�6�Z�h�f�1�]�)��mԠT3.���lҪ�v����u!-�_7��#2�BST�O�0u�r/*T�ͥ{[R�A�	�;�v�ٷl�L�����ǅ��Rb��v=E'�t
�x���J�lӥ 1��<��ۧ+VR�-�hz�,�yWs ���/5���/FM�pT����͎��֬5���bnb��7TY�h�k2ᬩA�x�V�Ѧ��ZQU�u�1�f� ��sCt �'tv�-��s[)�f�5c*��ݽ��N�9o����ok�l� �ج2*6V��VR���[XXf��%�E#�ի����2��=G]�S7��K�ڙn'����6��H&����һ(�꥗��t�tCwE0�r��f�]��V��қSj{H����V����ӕ�,��=ĲH\d��;�DAxF������n��������T0z[���F*JD��4m0#�Zș�A���M��ә�����ٍ!216���[�vch��mf���m�nώ�S��{@��6�`��q�DH�m��,�y��Zڶ٘~�e��F*�c���֩P�)�`YDz	��U�����{�`�ş<m��R��iO*���Ԉ�f�䷦2�^PS>��!3r�x�f�-Jh�`���,y�yS���2��g�zJ�&��ۘ�����ik5xv�^ݍ��V0L�pƀS��Q�Y�J�-Q�r�9��V:Z~��\nU�7c!�t�Z𫩖(�2��*�j�y`:�.��gU��j�Fs�*�X��ݑ{i^G{�6�8��ژL���-�JM۫��F�ٻ h�v�Eaq1zq�ҋ6�PiBX���ՏA��S�GH%i!U��b��m[6�'�7���-Cl�,-T� ��ۚT;-ۡ`�4	�)�raU)mX�GZ��k��n������-4��B6��	w�ζ��7�*���J8	�����l���y������Ud `�A����`"ʲ�,]B�d0�un�J�{u��ٺ�-IP٦5nڗWv��з�fؖh��;��Un��cD^��"i!@�"1�^m��j;cn�<��x^nX�˱a��*�S�p���U����w�hܽW���KQf��Y�^�1"K��ue�-)v�Uc0�NY�F�r�Z��cٓ��5njBY$ŵ�/Z��;.[���UGy-GX�8Km�Yf�bPfZH���f�V�]���L����Rwj0�jZ���o@錊J��1���n��]�lZ�����e�u{{�ǯ\�]kF[�n���9��SbFw�u�`�j�Ib�*
��LE�S�W[CX� s�oQ��ܬ/ط]�Ck�V����l�Z���"`�)���醞$A��m��GX���ΊKn3���N�R�Q�\�YX�^��]���udS)���g�kZ�%�P۩5 �,a�+jO;a=�����å+wZh�c+7Q�c1�v�8�®�V�1�A��΂���ɹ��K�u.7����z�� ���VA��r;N���"�#Cq�1走�UM��/���v*mU��黨(��#2�{d�����^�v2S�ۛ�.�m]�%����;v �bh)S��]Ki��u�5�1mк��KWOVʱb�
:uc���5�c���w�b�cW0D��oRU�X�-��`�E��T"O6T7>U/f6R���6l�6t*�X�J�uǵ��b��Ac��Xi��
�+q�/،&�tq�Z9�s���u6()�I��V�J����vo.�m�6����f�4ջwDQ�Z��sVd$p�B����(�)�Q���մ#�V�'A�mR�My���I��hi;*�6�n0�9��l��mbw�i+:lX�h�I]�॑��Z#��IP�C�4f��gv#Tf �3�S��u�q��#��M�m�i(��Ͱ���ut�U�sh�Ձ��ۥsv ��(�[6{i�)�٧�dcY@R��dU�;[�nٻZ��r�B�Ja"V���nX l�oN��ybj��9kƳP�r�n��t%:'ʶ��rS1]́Q��ҶQr!���N�_m;��.���(�3h\�!+�$�N�b��#ј������
���ۄ��tH�H�l�ÚE��0��=�n�$\�%�$P0�HFYVJ&�:�éJ�	\T$��q��Nt6��Қ��n��5��]j$�6��e�Q Z���bƝ���+�ڤ�1 u���6r����ʺ��BٲS�:y��>J)��Z~WR��W%5sN�h��RD��1 j%I%�:M�՗�A1e'ˁ-D�e��p7J#z�&*�U�%�Ř�T�5M:[����l)�H������`�Uʚ�'�Y8I��YqG�p��jF��\]�q0X-��ge�I��ꔷR]"���:�;�����f��!����ē��sð�B6�qP���7Y�^�{��O�ڴ�J���Yk0�Z�R/o�LJ�cD
�V�L�JҸ�E)h�)��M*Nҥ�����$�l}Kq.E��bi4j�%QdQ��%��\���Gv'�#	*�=2�dY7a�7�޽#���q�'I�rm_$�&���ih(z^<+N����b9{[l�'I�8�3	�ɐ�:*I��Yt-�C�!�(�R֩��u�VD�k9(��j&	�M$�1��ݫE���+�g=Q��)o`�nwv%j����܊���WJ�M�_r�](�j"W]��f#u�㳸nrk���ú��ar�o���c#'C��ORX�),�T���R����~Q��bU:�We�h�w:��X�;i�mkI%JQ�9f(B��5��6��l�F��㺚[Ut��@�W�qe(
��6�OSG��N���+7faT-�f�v��h�M�'�;&��U�z��+�\�G`�Z���%�q4��û]khP��A�R���'qlqwQJ�[J�Ð�,���[d�YxZ3� B��zl���'��բ9RJmh��$C��ХX�ORI�"T����i8��Fመw���;B�S8����Ĉ�p�+��T(�<]ݡ(Hr�ٜw侕��V�V�#ˢ�����<'I���v��NcF��l����QU)k-+I*��ȶ�O�u@�j��%ȋx�0�T��ٱZX����O�D�V����U�}қJ#���j�cK��
���i.J'��yKN�꼸H+�uC����{�o�����������������๬ۛ$����-�պ�[ݼ�^O0����/:��s犲G��Tw�,�MM�ʬ���?�𸰢�X2��.��7��ɗ��L���#{NZ�Z�U����6!7N�{o�����V�_^fhт|�V���TN�I�F40S|����.\n2��,\���J�c����1��&�S�����.�"�i�\���kՌ>4��Ύ
�f�.;�B�&�#4v��RXӐ�4���P�iJ�+r���������_|��RŔ��&�eܼ΂�#}�r��N�Z_e�Wٗ�I���������^���S;k�\O:�k��tx9agK�F�)Rr���fv����]�P�)Nn���n숱������[K���%�)́L�e0��Yi���}�P{�1̈��Q�/���ٷ�w�F��q�l�Ԍ0u��4�y��Df�9���������q�TW���fTO�ި���%���`ꃝH�e2���]�E���2e�Xk��ȧI�tQն���6��w�rƊ�7i�Ii�3$�|�ִtWmc���"+�+A��2�uv���{y�qI�s�>�Ō��t��k�XT�㥳��`RnBU��Hv�AT@�S8a�֔s+qÅ��|���c���]� #+c�Q�������V��5�O3��	6�w�K$S�����V�6Z�p+���Z�dּU�+��K�ػ3�\Ǽfe+Eic�Q�|Ļ�R�
�(��W�_[)��xE_mEoo��@���k;&v�D9��W;"ӕ.�m�#��=uxcJb���κ����j T�G�ȣch��=��)����W�p���F��q�T�f_j�9���%�����բ�������ߺ�r��;t�ꗅ��(=�����hf�*<F�ջwwǹ[N���Q�G�MsDy״.�K��A&+�a���5�-j�mU�]Gr�B�'�sgehٻm�n�9�-�T�n�mv�����vU�nR��X�����ܰ�^��BR<�L�|�0�!�_R0���X�9���e��E�>˃b��v�O��C�L�i�x�Zj�ݾ�x�J�	�,g�,�y�0.;\]NΦ�t�wv��w"���&��腐PX���M��9���YŅΊ��]w,cCYG���������t�c�����㸱8#�G�2�ٵ�b�պƔY]9@�O�9���Nh试�W �ެ=m]K�v��"���1sz�`�R��G�
x۴�� �3���(��Ts���;S�_��t�!v�����c�Ƒv)����\$v��z�1���q+�V��J.��5uAEt'n��v�N����5W>�|�3Ag;:Q70��K)35<[����~L���U���*���Ͱ�A�sI��ŋ|l���ɯ��lwb��b��f�(v�-1|.��c�53�q,����vB	�ɉ�K��`�*�<�P��I/��w�
�KE����`�ɸ��������oA<Gox겨J�y�o�N��)������R�ss�.����$�Y�ѻ�+8&ᱽ��>��{�Wc�^��n�es��ź��+��GfD���x���=1�b-i/�&]C��u�}:�t��ΐWv+�A��v��}�a�#'L34�Z��۰������(Q7�%�
���&���`�[;}u�e�N�.43�$0K|����s;��Vڱx~o�3\�\�]3/E�'s�ԥ^)��Z�s�'LK��a��y��+q;͘y�R��C�]\6���ؽ1���l�U�æ�Q�v,4:�nM3M@�m]Y���)�!�/)�]�����1P΃SbƗ�y_���\���d�Ʒ�^����_�������u�P1K�G��oi|�������(=���嵁�md������Z�כYڻuJˢ�K��Vn�'��c�<)v��ȩyۗ��3��9�*��vxT��w6�D.K�S�B�
��W#t{���u�\0"F�s%vK����r6�C��ڮB�s,s��tz�v����D�v��撂�{4^N��lr� �2��4�;S!�ѻ}ջg�h�صmک}p͋����R�M_Q���e��4*ǂ�Z��SGvY�
[��5}��ol,����[�9`-����;qP��x!A,x�Go����1�ob2!%�Vm��f݄�]n=G�җ+`��L�ygus�VĮس�!޻��g?uo	�¢�pU� ���PjI.��ײ��h]��G5��9��r�y�dn�̥�ʼV�H�`3����خ�^d달�Wr�Y��aw5Y�LD�.�O��Z�𑬔�M��UjS���
Mn�T��L�sН�;�>���.+=
��0��L;��8v��AwdF��B����>P5��̪��9qfR�����k	~�h_N���I�`��q�j�=Xn��vL�uA��ol�Lj����6�a�Rm�w`�8
K�GF�����F%evVv���]����Q[�F��2�T�W���泡ۨ�����T�J7�{�u�f������:Ȝt�kp��PA.,��8VR^q��+[��h
��Jꄔ���+ir����c��u���|��a�c욗R���`���a,rHB��B��&���d�mit�n]�l�l��>�gl�B���n]����]j�������&��o��Ń���V/(qT\Eވ;;so�d��mo@���zzΗ�]4\��ܱ݂��&�'��|�\����!����a)�i�捗���X;��!˕�̱����J����G�q��w��e��+��^���r�Q���r�5�gz�)�K��8m6*�� ����fi(��4V��VKo4��� �}Z�����;k6.Vl�n&��󋁫;�������W�ռ�/�R��G\�O;:a��� l� 3bnfQԹ���gP[R,u=y*)Ҋ֭���=��tt�q4v�(.EA+}c�Z�w>����̎�Yr�3�B{>�+"��]f1d��ֵ�>.Pk���S*�n�ÖSg�S<N8���ۭ��i�=xM̳c���O98��E�͋����z�l�u$�uw�,�Vܠ��C��v����{�]��ס���JS2A��w�бgK:�+8`���{o�޻N�j�>F���I�Af�-��8+�e�a/mUjv�쩩��n�9���.�i�|�'f�e���Ͳl�U�k5����m"�]�t����FY�C���Wg��;�(c��Ng|�;{z[7���BtQ�,21ű��5E]a�U�*P��W���}��y�{v���Z5L�c���01�q,�9}=Z�ڪ����>��Z�����x,�|_w%3h\��*zG ;���́^�>b��[;Wۍ�uf6��6��=-�%�{tj���]w4���^��ͼ�����UwAmU��gyqt2��b��ô��s�z��{�����#�8�躕D�"����ǎȫ��È��>�j)���y���c|�ؔ�Zz�S�R���}�����P�^�w�=�/�^�!�e���c2��%K�����bŭޝ.�f��T���K�9o��ͥ6�X9�.i}�*��J�TT+7j]���-ʰ��0M&�WLU��Dj����sx0�n�������+S��npɼ��!�[�2�6RSzK�3�^UA��.��eX���N�5<�~Щ�aW�q�b�`Tu++�qǀ:�1Z�y�%��@�0hb��5y���B�IE
\�Г1kU�tQЀ�n2Joy�U�ƻ��V�L�{�-�;��q�I�xo�Ĝzv25�ls;Z�X2.k��I]fۭ�uk!���n�T;�p�Z����Ĺ�`R�i-i�mY�v� #WM㸯�dΩ��d��evkVμ�D�-�<���Uq�b��X�M���,s��ּ_JM�ov��;Wr�f�%��w^�����5=�J~�������%Nf�l:T��}­�Uj��{����z�⋄;r�i�o�c�Gxr���$z\/��i��H;�K�^Ѿ���֗�fj��#⫪vm���[�1|꩙��"靴�S��4,�}�9���gN��IچS�M�RԻ��ɺ�v�vP�؄՗�8_4Ol�"<:���-m_)����;�	��X+����WR�Vݠ1WNh���}��gs7C�u-W�Y��#�SPa����湜&P��ˬ����� �y]DA���	m��I*}Rܬ���7�t��(J��vmq����fw-�{��(Gz�Q:A��J�5�1:�l|{�Pq�;�ݐ��o������H;���m�u�u&u��m�@��h}/�ލa1:�:砝��sk�6=�V�n��v�0�Woe����ݭV96,udfg���&՝��Uzlk�pl�1nc�s�Z��F��~��*��M�����k�m�j��]�VoB,D�]��y�B�<�x��6f8�wF��Vs ;[�~ɺv!��,�^��{�CO���Tk:�yWg��}��j��U(;�����G8徖�:�e���XR�gq�i��b�V���
\{�v�T�SN3h7��
��&d]�W����^�js��\-�\�huY��I�P{w�+��+���Z��'Z7��bQ	l�]]w
��H:�Gm�V�-}�B�*�SW��u��u�K�64���C_[�C���v."���.�o	zG�����+;ff�����.�S��,���]ձ�t��}����{Z�T���|���7cs"e�t��#:�D�j�b(A9�id�����+sik]Zs���}g;��fծ(#C���z&7����`mT[�����h��w³v�.QP�u
�y# ���ޔL,tb���N��l\�,B���O���m,?t:Xy��fVS�Ԅ0��U"�f�Ә.�Z}Kԣ�HK������4�����M�XE9t;l�j��|�1;]��"60q��t���R��ͮ�\�ɵG��}�]+���a=	�7MV�=M�;�V��+W:���Z;�.ڡ�6�r�Z�qMf��[��x�}�4�̆L�6���p̬�T� ������)�"k]ntywZ�ݺ39����r�n�/��#1[ڈ���Cjٔ���6�_8,��'q�K�9��{��mv�O����+���k&����=���МE��F�Xe�n�C��䊭��t��]ϡ���
y�_�Wn��4�Ԥ�gF(�&�i�͐K	�k%�B�mc�.���b��s%��ځU��A�M�[��/g�cZ��t��Z�j�Z����8Rc(���)w·��B���&�_vvN�XX�}yF-�U�J�&�qr�^����t7��=F�/���쾮�l9��wm��UF	0[��y/��ZÖ]�7w�k'?fCX���E��w�&�-�C��Ņ���yB�u�u���Na[�jj�d��g��T�ꓺ�`IG�2��cg��l�oj������ᬰ����^)y
ZōJ=g�֙�>����H��nwY��_�eM�X+rb��+%�ض��X�bA�uԨr���vx%i��/���t\�F�%)ْc�1n��v�[�pp�Y�s��,:��ԗ;Xm��֫��L�2����s�z�+寙�6�w��A�]O%�8c��WSii+������kiX�r�oP�쾼�j*B�w�6��䝙��)-<��7{0��	u:���6��9���x�A��ى�����0�M���9�����ںW]�9�������tX�OQ�� %b�ޣ4W��ge].���Z���ޭ�%���������;��.Mwhb��x�5��8���=��X����y�H����_S�ۋK]ԁ�aZt��ͮ�{35a�I������k�:p�|;�q�N�f���0A�$�>��x��v�@� v��.@�DԸ����9��t�=�n�9�v+�u�y�yUp�T߅y��{���.���P���9T#�҇ �r]
n\@ު���{��PC =*y�sT��y �t�����O7⛋Qd޻b���7�77#�|�<�M����	��*I'����ȡuEO=��)��+���^tߖ��.�R���<݈ku�|�$�)��<�lOw~� �lכ�y;�	�A79 9 ��P�Q�	P�b�A��<׋QC9Hs�%̋+v��v�A|���{dW��J�+�ئ��[�����_!�@���������������<~�	����	��� (�����|�����oϷ��7��ﻙ�O9�à�ʃ7+K�8�Y�	Jݬ�u8�2���-�����W0�3�T���9�=��	ڝat�p�����H�t_���Xjɬ�s�uUK���ʎ:{=�8[�ڰGI@fYkv��W�寑	��$�s�{���z�ϰ��wIrmrV�aJZ��K{O�����s�v��ut˹7aQ�C���<�����+��|�(��1:
p>���V>�Z��z�����;�c���]�k�G8�Y��a�J��۫��|���e��W��� ��Mݴe����H#3��m����7Wu�
���y޻Wufb�ޛ[4췗;��*�X�A��f«�0Nڼ��^�ʕ�P�}2����r�Q۹�g��$��*A�kx*r���>�W��S��nm1o��!��mp��j�K\0���a��\��y��a��޾;Ӝ�qݱ�UX�gO��������p�f��&�,��^O�Gy��f�;{u����6<	j�ӎ�f3Z�)�3c��ԫG�nݕn�,�P�#д�e*2]�]e���R6�w�T"�0K�Un?�	r���]{nh��=VƊ�m �8��R[�`y{z&S/�,��q�q�q�q�N8㏎8�q�q�c�8�8���8㎜q�q�8�8�\q�q�8�N8�8�q�q�t�8��8�8���8�8���8�;pq��q�8�;q�|q�1�q�q�q�8�q�q���6�8㏏����<c�8�q�8�N8��q���q�qێ8ێ8�8��i�q�qǯ|�{��:�Dh�;�J�RM�͡'ҐsQD<F�a�ْtk;��u�tp���ck}en� ,2F�����yEn�nR�F*O`Ls������C6z���KF("���kr.7�\�X�-��6��o]�$m�,*R�4�A�t���I�jD;]���+I�O&�R�M���k5"��hЍ̗�Ý�	t��ʴ�­+���V�A�s7v؜.VT�e���X�e��B�\ B�em	EX}4�ۭ�TT�3Pjj����:�4*��bp�'I|��mu��y���7����Z{���}��8�`�8K��5�Bɤ�l��r'"�l��X��6^�َ�*n�!ib��op^�0Ʀ`�j������7Y�����H���j�`z��[w�u	� %�@��
uo�\Dm��� ��Z5��o&��^Eb�]/�I���i�d�g#�I�KW��'gC���x�⺮d�2˾u.��͓Sgnۣ�OL4q�=(���
�qX��z�,���J�.�c����޸tvKL�IF�{Ā��RlG��1�݊�ȶw�Lz�D3WX2���l������N	�k��zx�/fNL߉R��b�f-��_���ز���Lr�[H�M���Y^O�F�>�������88�8�<qƜq�q�q�n8�q�qǮ8�8�q�q�q�t�4�N8�8���8�8�8�8�8��8�8�8�q�qǮ8�q�q�4�4�8�\zӎ1�N8ێ8�:q�|q�q�N8㏎8�8�qӧ���N8�q�qǮ8�8�8�q�q�z��4�8�<q�8�8�5�r��[s]&v�ܻ�BX�Q�=���;�Ņ��{^�{����eM��{t$��sB�3!��ΩM�H��R=0�e��Q�����+Y�e��Y��ުa렼=��
{�Թ �`F�YV�OG������Vç#��ҝt+{�ɬ>����lsU��j�-�W9w�6��S%5��,d`ےŢ]#"��2����s�uɕ�@�_P��۔s'kuAA�i��(��˩��"Yݷ��=��}���1��]d`׫{��N9���]��D�S3tIc�S�L�֒��[w��Aq��r&�����C�ӌ������]zh�c����fMiK�*!�9j���e��O��z��jر���]r�[Z	��z&w)�-��*ö�7�79�z5�����)Ъ9���f�x�Rku���k	�[YxːT=&�r���B�J�hk�S���-�g`�/5{���Id�TۗI��]P[xDS+��Ý��Խ��8��8*@غ���MAAkʻ����ٽQq3��9��`���#zKPZ���:����9�ʐ��+��vf��+Ec�rfF:���sc���{�ە9JYW�fv��m����n�8㏎8㍸��m�n8�8��q��q�8�>8�6�8��q�q�8�N8�8��q��q�q�v�4�8��c�8�n8�8��q�8�>8�8��8�q�q�t��c�88�8�8��8�8�8ノ8�8�>8�ӧO�8�>8�8��q��q�8�8��8�q�q�t�8��8�ރnl���{�p/oaM�2ԾnGS2�+1���̻�ރ�%a���Ykve)�.��'l������Ӻ��2���0�׉w=C��W#n��h󾼬�N��3n:�s�˨WDSX��a's��n��ZŹ�:Pd��/v��N��� x5�DZ=K��EE�m>Am{���\�Fޔ�L�UKt���gj�Re��ʜ��2���nKjt�cP����f�N��.�Ot�Cj�� Ma��e̩5���C';j��=�RE{[�[kt�Yj�	c�xs��r�1*�8�WӞٷ-�򏱧E��͸w�٩�	Vw��֪���B
�_{�=��ԧ:�b�kw�F��(��}͝`m�{iS�Mf����v7�utO&p�6�
���ɛyV��w-��Pb���Mel��d�D���G:y����P��/;Y3`
{W�,�B�S�=�Us*�LMPt  ��պ�k�T���]���N�{�Zqc\`�S�)Y�i]d�؋2��T��ٌ�����]NGv��m��(ͼ�\r+����w��1-��zA���D-w�d�Z���,�z<"�n���HZ�}�qNgz�����ڻ�]����.����.��,C�3��޼�0v&��f�gY�XO��G��B��WQrY�`�E˻V�l�@Lbek��"��������u�=�f�." |��d8�-i��dj��i���C���nۋ/�Y�A�v�Q���.�}LP��vu>����0wp�CF����ӫ�T��X2I�#���5�\U���u�+;�rGA�����YE�&��;D��r��gXv�&.ۭwko�ޔ����oy�b�Hxl�Q)F�{N���շF�I+�j�W|6�hiH�yx�����"�x9)Rn�/�J��ga���QvCn��r��v��R�2�c���u2�o	�5��Fo��Hl�{[ٴu�*�m� ����[,��g�X7Zj��(U=I�c��C6�����K$�xVۨ ]�ZyI%{g� ��o�E)�
�K[���������o�0a|eL�L����Jì�AU��Up�B�A�wQH��r`���X���X�n�Y�u*��a��{�:S`�꒸�dyD,W4�ݩK�a�g2�X���q����;0Ȥ��Mw[�n�fS���Q�:�%rx�����<'s���u�6y��߀�m������y��Gh:ܰ�ޘa�V��[�� ��Qǡ��墵���X�Ġ^&J�{d��ݟ����!v����WVN�\iK/�a�XG�)��������]��5�b��f���-�choHB?aʇ7	��V����]2��&ZH��P0&n]��e���'o�7�q����}(�a�wX�ޱ���&l�j���'B���y�Ou� }�r��Ӯ����ToHu;��&��%e�t(���Gd7�]�v| �uf���91�v:��W���d��6�px��v]�F��,�APowK"�\SL�i%yTE�q��۾���I�-}�+~����Y�-����l����%휡mzz��MKwN�ڽ)8�[^�T:.�Z����*i���Ռh���]������׈;O�:yOz�3�Z�P������ɲ��!!�C��S;qHgWtۼn��tn�h��H=ء]��Ow^���rW������D�q�V�W{����d�0�۠���e�F���oc跰˖�[1R�WM`��c��+=w�K�&�;g��40pc�弧ȱ��`{�k�����N���W����y����w�hw%C@����J���7���ڲMF��gc��]O��1��QZ�!;hQ���Hcs��p �"�w0<�2��<��LE�I���rM�2'.�ۜYڧ8��bl�n��Ge���5����Ԯ��[(��4�K�fLr�yx̌[6�u��r��C:�l0VN��0��i�ÖG�V��kFΚ��GP�|.�,n�{Do{T(nt)�;�EM��[���z��\F���� ���L�T�r��t�ZƆvn�wAro��/^��v��j�0����<Q@�Q���|#ރ�WE��%5yrY&ٵץ����Z���V��}�P�sO��.���'la�yܾ����FjV�A�rR�s�Kٱ8B�9s@ ����n"ӳ��/��6E��Ñ�ħ/���r����ܖP�P��,�ۺ���3x��}�|��t�{/��ꋩUǲ�-7�T�a��9Z'��>aWk,T��������ӳ&z�Of�ޱ�4�2�<�g�	=��y}�=��6�MO�D�H%滺���鉭�a���X�#" ��+�*`�j�MQ;n�^lvX�U�*�m�F-�z���:Df�;Y'X�%s4�{�B_u�n"/z�L��]X92�Ch�j[
E4�����W�veW��tZ�55�YG�p���M�Cx��_�m�ᑙsI��(駷�)��G^�7*�s�=�a�1�Uz���c"���  n��WQk	��Wӭ_$��]��12�檺�jI����Y�{���bٚ�m�+� ʺ>�ʯV�M,�&�Z{��H�QmVݑ� J=3�-�cE�4�ޤU��/y`�����4�At0�Y��Vn��"j�ݭ�p�5�zn�u�)��o�H=x7q��n�w'��v����X{��V:ΰ�jjZ%ۥx��E:�o*饱�Ձ�������( �Y��r�l=��κ�r�-;҃�oj��EW�{E�}Le��6���^qJo��Z�LY�P@^���eeI��(��z���~Lv�IIH�Nl��WLP�٫��*\��`e�O$6�b�����S(Jiӕm0dw:�p   ��I�c-�#��x�8>�X�z�S��9�}���<g�؞�������mL��
��ƹ�>�A�7�m�5��{���Ρ��)�4v��Uz�d�w3�i���$z�U��2\%XP<ڶ��kpU���+I��
��㓚R�l潪O^�o*���k�+�v�(��F�!s��rM��L�n�����
Ն��.͓��5�:�qǢWn�
�j�5[�������3d
�����T=���&�x�)���g��l��x��l4Jp>���lnab����&^��&wC���zܺKJ�І����u����I��zF�u�V��w�/�We�9�z+8^	"n��W0��{]v�n2���`��{��{����S�޶����h�k�vs���=<���� D��}�H�:�!˕Y��\��ZB�J}.�0M��-�\��ѫ|J�Y&'�� �\Mdz�mu�i��(��R�ю��8s�/pW8ق�|��1��opͳ���9Pi����w�`nA6<��]Bn��%r�Ǎ���ڜ(�/r�b8�����`�ʍu�k��*L�9���~Ie������p�j�pL�ٵ�������v�W[�n��_@�Sӊd���Ϲ�|;k&��_R|w��Y�$�onq����;e�p�I�Nl���y�����dk�� v�v��*ֵ�ƞ�׼��M�*T�&����&��[̯W���c��S��<*��e\W۫*�/r�M�pBcR��V��pOR���w(ڢӛoz��QGz-s:IW��;��]�uD�<�7ЪH�޺V�'٢�U�N��@�ѕOpM��g�y{_T�O~��1I�,�9Xh\+	X�=F;��IR�ۣ����=j\�&�j�b�w�������[���k��^�*m�X�p��Sa$'��m.�$���!ba�˵��#KT�mK]4����r=�t`A�4^!�V�oYF�����}%���W9�6�]Sfmt�:�����N9��2��6����)
�mHs&�&��"n���n��3�'�Ju]�)X���r�nek[�}�];D�Hrp�΍�WP����qmv z�����1\�
P�f�[yHkŇJ�; #h
�^k��!q�u�Ne ����v*�Ɇ��Wu�
��D9: p�:�}�����wY�6VGn�6U����&��]��ި{��c�w�[X����xs�˻��՘��N6��cyΜ�fh�U�p���h���fie�5	Ҙǀ�D|���a=j��Y�=������8Mh��7&�$��rļ�XJG1`�/�:�h��>M�BՉ�r�˳r�ńP,P���6}���q]��T�Pfyf��n���/��֋zq��+���P��_%�Ũ���BԳw~	��r�ìI���;u"��͜d8/��Z���=�wn.d���e� ٷ����FS-�y�^�n�>�r�,+�^��Y��M����$�0t�]hB�V����f�S#�V1B+2ble�1i��	ҹ��ɜ��W�[L��=y�{�e���u�t����wە��}l[{�2�r����;#��A�6[���xwC	J��cr�S��4��E�W^,r)���.������Ly���+#;��m�et��],*���J��ĵ�n2���1��� +�2���?���O��������%W�k�ʵ<�W��I<�L)�rA��MB�!6َ��?�#�#%�""�DFxn!$N2�F)#I�ᓑ�Il�<bh�E�UQ�0&�$)o��Ӎ�D��%�8Al�I#D����1)�J@HC�T�
-&�?�t2��l�<eP|��b&�%�M$�E$yD@g$b([-�ٍ㌠K�Im�F�d��P�2.3F�H"��B�P�,ēd�$*ʅ�ь�L��J&80���#��T�G!q��DA	��ۃp[H�K�>�Gs�VN�s;�nkF�:�jah�=`ż&ɢ��@fؾ��9���\Shh"�*	fe����Yw�*&�VtCA�o5���q�Lͳ:�v��p6�d<kU7[gP˾Z��8���nKU�vX�v�WN�j�L"	A\�B�{A�'Ke͹�����vx��HVIthGF�Ur#k��g2]�pE�ӓE��f��DʁL=w��\x[�MNq�Ou�F�A��w�3R���ݶ2?[�N�u}��=l-f콵R3�q��+S�:��pv9��dٛԷ�L��{�&�Q�`�\�9wu�x�9��:��Ś�U��.�5�4uQ釹�ڼO�+�����
��a2��u�I^`��AvܧѨ\��f�vd�O
��t�����kk��(/��,��у����+1�i����2���6�}�p5RY�t=k�F��u��[���vn���4n��zx��Pޏ.BZK����jh�K���x�0�Zŝ��ϰ�f���9����S��:� �����uS�[V�!x��\8�֘'<�
}ӦހA*�P*�5�����b����t-VΆ�6g3Y7v���L�[��>�v���7���LCoes���}ܰܺ�q��ub��yTP�8�E��
��[�D-�
b#PDBF�F���YRFCqȔ!�jIb4��,�l�X-�Si��$#ʢ�d.D���FF#)!	H!���e� -��1E'�rHJ�6�d��jD�)��(�QD��HH���.҉P$:��cMc�>3#q4�I�$1��A)�$E��biچDR<��k��Z	�ZA�K(�DD@�q�Za�b�IAa��m�� xd,�
b�%�"a�
�U!"�TI��L&\���I6�e�г �E�IJ�""Q��%�#B<a��`�L9$�����&�d7�E"I��!B�QA���@��SI�"�R II$�e�G��fJH"$$�e�!�(Q������P4x�r��)�-���DI!B)2�B2�M	8�!�\4�H��Y�ZN2�bA"fDTd��4���S����	Ear"�Q��e"��|h(�-(	DZ��@�ʀ�Q�D�@�-0�R$IL�� 7�!)��u�^��Y�"64z]�޼�c!�nk�����$������}q�qǯ^�|q���{����E$�`,L1QF�u�C�wu�7��v�q�q��z��M�t����]������D��s�so�]��I��$�������lx�8�8����:mӧZ�D���ђ����Q��

���i\��b)J��\\���.2����͸�72���U��s�"Q.��M�殗8mw~yy<�r�xyI��WS����k]jCs����Vw^�*�k������#T��ֺwww;��X�g6�wu�:��p9�Nv���r���o��yj��y���v���:5Io}��<��[]<^}�u�v�{�y�a$o;[��wr]�ܺ�v�����o.�8�����宪�B�Y	S%�
�MUCUݝǝ��ݼ�����;�u�����#3�y۶xn\���;���ݺn��޼�/;��[����wS;z���.�]�����7�\]r�.�'l��\�(�WQ���>v��М�W�_( x��8���m�$0�d)�h��,8I$���J3�e S�Q�P�ȋ0�a��6O ��;�����aʕ�cx�^�eG�%3�y��|��3W�}VnYTy�U�/.�F:\�ۑ;�|aO�Jkd�$��,3 S���I<e�Q��I)�`q����I"S���ā�A�i���q$�P��Qq��a�‑!	$# �"�3a�\15~���1�ch�����j(2����[��4R��`��*���w�Q7'��Z��g�H6xWv/.���<�F
�����+���%�D筳#��YԤ�*�;U~���)�]:F6j6�����\T9��WMdl��TQL���vgY���2B{�	����4;�r�H�P+H�Qq��m��Ja��T\D�L�V�8�P�طFΉ�9�d޺�`0�Q9Oq
�L-�td�sM�#I]�ʐ�t�8c�>�R4*�X��0��m3"�	���]��$��	^��<����w��`�`V�5S����r�!���zj�(ąx�(���~�n5�uj�C2)'��eF(>�R"�ݗk���ݹ#u-�ME*�O����WxSd�dM��>�ڛR�Y��inK�N׾���cJ�������ha0
]~~�u��쨳-cz�N��gh�[RzI��J`��nwG��}C��Eҩ�5)�ܿ�E��,�[bWWl}t�j��^q�r๷e����q׷�]��[.��i����˩V����;�G����cS���	��fm立y@�W�#S��R����dd�{�J+�����G����%�O["�g��L�m��6"��t+j2M^c�c�h� �����:����֏_�ᘬ/t+r/j�1Ȝ
mi7���T����+3��|q�UK����MQ�-���ERL��{D�=��d�^�`4�ޚBЕ_�%9^z��[������[��k<�Mb�^c�*G�O���+Ƴ�h�V/T<[һR%�F���R�X*���@b��qhJ��u?��Avµ�<�A[�R����U��p��7�v5	L���S�@3�P�jaM�40徇1��8�^�u���X�'(1���IG��|�ۧR\�S�{9��JI�ѧ׊$l�Vޑ
(����)ZPm�ǽ��;���+m���IVO���n������P���:W�^I����v註/�㮙��f�TB�'�H�u��!���}��?s�+'j��gE��{8抺t�o4Q��iA/�d<�CL�ĭ��b�m���>��2�	��
�:��W��xxW��_D�j.ѫd���#�3���k�Ǒ��"���󀰥���E�NN���msQF#4؃Ѧ�_�L��9jf�k�J5-�ۈ�#dF�zz��w�"�XӶ����6"1H��#6�R͆Z�&^��D�}[4U�#�w �򙼖�_��Iw�3��Wg}-���*J�6�ߪ��v�}��1=�B�A��p������5�������6y�������F�O5�Y����ٱ�&�ڰ���m��{hɠώ�5�fcS��Vf�)�i�'�l	Z�*G��r�*p��~\��-�h�iy���*_�_�y�`���a]��'/ �#����)o��!Ia�C-��u��u��:U�*%\^򬬟h����_=�
�N=0a%zBL�Zխ��[j1▣�a�
�����y���`�=�R7�K�]�χܝ��ӂ��0U�H䕎�B/{χ���fG�d�~ޥ�*��������q�svT?fU��᳹?%���zwr]*hs��oK��K<C��C�jK���f�1��[���7s�ݯ0�ڙz���k��Q��y��a�j���k$��"�)	g�t%5�<<�$.ߒ�6����V�Oc҈�9�k��}��Y�3iNЄs�F.�i��+ü���f�;�|�Y���T|�I�kv�aW��
S"ἕS��Өe0*i:K1U�&�!o{��(����!"4�2
"N�eU�
s1�e�1��t��s��r�jH6�s��@ '/gg��Y.oc�$��s��8��y�{W����M
Z�-�1�6���f*W.bҫ8E���1���!it͖�n�2 `�:�w*=�eJ�`��rF�g@f�TMy���� �h�~b/!�3f��h+����NJLB�HV6#ڴ�yn-�AN�+$m0Z"�c7������_��Rt�J��--��9���v����r�UN�C�4=��t�&�������7�˜^`�g���ʹq�]���\�č�I� �Wݵ�"��މ���@coM�H�2m���:��Ku�z�zm:�;�v�6��{���h��⥓#7vb�G XN77���^3�x�5���S��� �~R����%1*���ϝ��Ӻ���\'5�K���7f�ta�ĉ߸9��"Ύ<�({�H2{����0v��Z�zNibl��ȇX=��ŕa��t�W��u�B�`�Ϊ�i𙆽�;��m���x���W�-W��u��������	�{�N�,�?���^�-ո�V�*HCQ+)H�`���M�����wu��3�{����T���H|�2�﮽{!�3�Li���C����U{����IT��`:!�J�nf�7�3|E��Pū�+��&f���S#��W�q-����L�&�%d���f`Е�yXVf��ɿ�qt/���4�|V����Z�J[s�[�"̈\fB9�����$2�ڕlQ#[�}-����IH����`C���al�TDu�BY�k.��mV��J%B(dn�6�3�CI�h�����Rᵩ��.(�t�쥫�>�Hg��Y��,�.�Y̾zS�g�z��5 ���=ނ;��b�O��؅��?h}���l}�K��O�O:k��[��N���ou�,Qr^�ف��WqE&�ڕx[⃃����]��
��*����RF�;y��	0�/ m���4��&B������������\̊r���FS��Z3��
�BY��i�ʙ�&Y�Y�ږ�"��̽��c�Y��o�
Fl�u-�Q/�j���E�D�[�fD��^,F�_�*��0�3}:��.�v`��Y>mŏ(U!j�����srFV�m��֑���lȀ�
�H�F�C9��`L�NU�Q9�Y�-�~���;#h3�n�װ�<*$�q�v�wx~��N��w�뎁n:��h*<�Q/ �f+�uӸ�]��_�o�9�*�?]��<Σ�|3���j"��ک�!=�ȝF��IϜ���%�i�)I�JR7s��E�d��[�i�m2�i)��=FzUz�]�'+�(e�;bB�3������m�����0F��Vc��W�k�V.~1��F�jf�����:�<)��~eH73&T��Xy��m�����ͣ/���!�ه�G:�1m�bd塽��c&T�ޒ:��0^<�G��zPV�y����ofX[��������U\��f�|}�ZfHݻ��sB���"��Ǖ�ߞ>� ��Ͻ����@_NR����5��K׼�:�)�n�cL�yS	7o�"'0S�S�M�l�Q�٤�lT-	$�o��/�Z��s{v�I��yV�CC����O��T�"�AIhMkc
'^c�ͮ�5�K*��"�5��>��"�G��>�Z���fh��-�N����)mUjIVF����,�L `<���ݽ��B� �Qb�6��t@�������&� ��A�~����){��U�b�Ś�ߏ>�9F,Ҥ�Ḯ����L��c�Fl89�jw4��2�U�y�
sYX�$H����ePo����f��߃��}wC�T����kmJ�#���j�o&�I�f�}8t�S�weL玀j��!�<��ԍ��$��i%�ZEz�#\2�+�tk$vC�n�il,dt�k��]��f�olε���!T��D�^J���G��;/B}�W}kI�
ҝ�3yf�ˇ���pK�=�Q���N�Jo�&�b��Jt��<<<<=�7�X��-�>�V"`�-���G��û���.����T��hX�鼹�ô�0tV3��(箪u��Im��f��ִ�Y��1 Fk��d/-�&��0o���h�|�����JvS*�T�Fi���Z��S�/jlm2�5�'Ð�ޥ#3���*5Ò�1Y,�P�J��B�R����v����3�yM)��O�gaZ�e����IW�8k����/mp�z��{'U���2�o��'2���T���������~ݯ6�T
 &IN�m7n�Xv[7�xOl��{i*kn���{Ǉ�Š��H�iJ�l������[:a��[��b�����]�+E��J������ �c.O�p�C��qD	չ;M����A>{gm�^Nȗ�6Hhp���ζK�X�W���Qׅ��C��VD�`lT��t�lHl��;��쓕Ѽ�!��˷y��
<g<=-�e(
�P ����!��@�ҝl�#��,d<�;Ǝ6xtQ?2�^����u��K�q�ڙ{��d�Fy�t����i
�ѹ<�躕ʻ*�-�#Ľo��\�s���@���쥛����c�r�	�Wl�+��]�f�نN�"0]��w-�W�����^}/	�����y����ܸ65��q�0�W������x�%Y���XϽ@�|�z��4�+� f��n�)b|�טNό-�fT�gN����
vVO��\�Fao �h��eG���B�"��IP2��/�������ӭ��/�e��P٩���X,0m� �1���c$uW{(w��'���?Wt������q��[ax�X'gi�{!� \`���4�7a�lo	�2n���!��$@�Z /�8�����p�D#�g�	zLi�XE	Ut�dN⻸mM��Ω!j"+)N�<d3��U,o"|x=�nAՐ��,�2Ɨ�vK�
�m)�Y�ɺ^U䖴��
��/K#�R ���M+�ӗ����J��O�D���Л�u")NMks�_a>�I8�u.!w�VӲ�ob �<��՞��ӧ�썬p�E<�ݝ�~�B�a^�3Qh<L\�m�ٯ�\���f�.�Kټ�ܺf�Y!��&z�O:�6(����D1����R<FR�� ��xG9G:VV��ȟ�)J40m5ɀ�{zYM�d���,�aN��H�y�{�0��|��꫶�JK)���jn�(�E�<�|�i5/S����קS(�Kkԩ$��T�)��p�|�1R�_vJ�%�-3�:Jݔ�ժ�V%,�;ZYyy̵ЧP�<1����PK@oE�&+am��m�� �D�PL�O���2�FS�eE�'ܭ��NjaB��v}����x�-�Y���Eɽ1v�,�0�%E ��h���o�m��*�%k�Xݟ%�
�Qx*�`R�3�H:XX��n�j�y�����Ϣ�6d�������#��Ι�������R��d6��g����l����Mh�L����!�_'�췺�zk��w�&�R���>f������]���<�Pj���Ϩ�����SC�G�ͨ����[�������k�jd1�+����N���
��,	9�|�C����r& �#���w�+����5ݧ5�5���0Jc�������;"�=X��WoD��G^棐R���3RC���v���i���"y/�z�}[}t��tK<��D��+��2��p��?Wn%���(g��"�����g_|��qPHJ��v���'rhy��Q*^�W�ۤMz�k���H��ӎ
ZQ����63;Ub˺R�TP::�y>fe몔lݪ�x#ג�gg��&�7ٺ�ݽW�#��w�#qNڏ%k�5F����[�ju��ٻHV��K&�%���,Sf59��p��ٗ��%�fd�c]t;4��W��]�[���X�{,
6�����3�s�c��,����
�WL��̔P�Zz��A��ҷ��d��M�{�����[�n�o�t��S]0��NZsT`���Ú��&Q��wB3Gz�So�5*��jZM�b�Rb��`]wC�Ŋ��S焷�ғ|�8aduA��ӥh�]��bv��c{��+�'b�3��o)�[J�=�SU��u�SJ)ζj�]g?f�X�3�����^�jK��,�CZ��E�L̔���n�܃\n&�:�B�
�!J���Vx�6ī�էtmN�eU+DI�{��������SX����Π��R?w	嶣�	�N�(=�V��C��[����}�W��Rt�]�+�ut�Z��m��]�M��%vݢ�O�핋��S��e��umS��c��Qj���+M�M�@K.��@�Z���g��ǈlA]�J�\��h��6��ꇱ}`P��-��uS;8kf$���.�;�S>'�c�K��kj��U�0m�ou�Q��Ƃl�ZO������`�%�I�lL�b�����w�ݔ�qNˬ$S)�k��ڪ�
���wm��"+�R>�-���fm5�79M�v�3n�m��ەS*F,o�O*.W{z%?:�ĭ���,��j�ܖ+�x^�����z�f��:Pl)|*�h�Q�r�6��NY��j�r9��A@ފ˫ڴ�3	���j^N��/�`��g΢�G/�!����ENx9�w�	j��z]���7�u.;aJY�h^���.��h���k����Q۩N'�AbE.n9���mҬ~sוק���o+U��Z�& S�z��6k��,6#o�\8[ޫ'/L�#XW��@�ͻ����F�9�}�.�����=��S�2��Z����篸���\�e[������2<�]��v�}�a�DuXӈ���]�c/����G���]��w{��ַ��$�9-�J�j�THy
�;���޼�����9��]W1UIʢB�U�(�c�_^<xǯ�8�=x����]�|v���$$���_%�+��%;�L/}ǝ�D��LRO;�s�B2}}v����}q�q�׏__]�|v�:$;*B�6��$a���~n��:����3g�h�}t���ǯ\i����z������nݾ5�$fJ�$d<���(�$�	�]9�ho��}j�H�7��	��wFd4��P�DDK�铜zv�۽wH�I���3�vbQ3ӲB�=;���׎����ώ޺��Q�Z�y�$�2'����\B~�e�������# �D���\��䍐@}�4a��m��t"#`&��Y�rI}:��sIO^���~~�~�|8x�Dr𫤧q9���pJ�f�rR��˟c�O**���,
��]˜<���U�w�ͻ}i�����SU��l�G��k�����U�?�\nM� >g�V0vF�$���W�*�6�^�T8�D��8����egU�]�% �!�~�������ڼ@L�!w:
�� &ʤ!CT���s�Ou�t[a����j3�����+�6�m����K>���j��}b>����@���B�ק���8Ù�����w%�(�S�l� v�?���ֶu�E;�������"2=3ql�r<�y	�<��v�tv�|U��,��xo3�-��Jp(�8©�z��x���=�àdE�>�X�_�w5�����	�@<$�H$�I���o|}�;qu�k�徚e�u��3twH��-�lj�E�yY��A��~O�-���ѕ��9�/��y��f��<���������|��iY�i?`�Su-��{$�b���@���kۧ��!ot�'�Ap��ٲ:��t��n��&�w>yDs ��Ȯ��,RQ��퇣��{�q��1�w�=n�>;�#�)�5��r��p��^V+����~] \���5�7�]U�̋�;�m�����~_:h����*'���Ǥ����Ksx��Q,�,�Λţ���u?�Y�pc'n|.�=k�TTy���i�	F���8/|�۲�s<S�J�������^�c���J��e+:�3��[��9�t��ݼ֙�zWEwh�.�/��� �ټק2ќ�y���\��g5�<��0�ȹ0d�Ha���!�i�u礗�s�̐�����#�\`��5�T�(V/7��>W���sv릉<  ��d'�� ��C���x�O�4��v�>0�C������kۋ:5+�9Uu�Os�N�L�|�o��+��0����{���r�zM0ye�ɴ99����]_u+��On��.y����|՟j�+���Y�� �Bs4���?�%��ͺd��aUy�n����3^��7��_�?X��
^��#����;�g-W�����C�i�P�$d��]8Y���se�<�t�S:���C@˂�H���zk�V@��ѡ3e'��q�ul(/ʶ̵ƕ��;����vD@��M�R����	s��'��,+v}�s�98n�r���k�7-�r��J�C'����W�\�j�|���B����I0,.|E��+�n�B&#��S!�n�v��{�����6ж
|k�9��!���U��͸�>��ud�O���-���*���d����^��� �P�O��~6zl.���n?�
���OGI>qL�\[H/�\>kK��Ο�5�7˽�O�v���)ܒ�`�s�M3KPǀ.Ȫs�b�Y����BMy�{�;�uTV���`�����[r��[������WG�R�vۦ7������@�u�]F�0����iNΩ9����b���>a��y��pВ2*�q�c&��V�]�ދ���:�fa�����������"_L�:Np�2z ;\��Y,Tsc6?0��1<��H�#���-��q��
�!?-���r-���_Ӎ��[&�qp�7MF�e�7aO1A��ѭ��)�VU����zn�Y�-� Eƹ\���ģ���*M��\
�\�jd ^}n!�h���DO3}������d��+�ɻBxۤ�/�>R$�J�Y���UE��c4c)lU��6���=�s��-���]�o_x��
�,�^Z����ݾ����z��k�$3q�$:�B���Ͼ�y~���S,���}��G�j�j��ۍ.+��P	�_-�}u�$����E���%��3�����>vݞӜ�0˘=7�80�ÌcJ��iP�`g���I�	�Z����3���昖��Գ�<��z�0��f�:"�yEz]��h���5x�ex�s5�S���Gk&�~Fj�j;� jN���<9�^�_A���)���4�mm�O�P^q��龤µ�hX)<Wtӣ���A� ���_�ö��<�E2oQql�E�x��#�|����ϸo�{0�ԏ�gB��<�ٟ���ַ�_'Mau�,�X;�8��|qR�<߹�0+HR#��C�y&MI�������咁�}�1��&,x�De�cl=�;9�)-�^��
\ƍ��]dL�(�#U��X��˱�Շ�k�n�qw�g8�xG�y��էw^섗��f/c���������9��P�/᪢��eW�h�2�v8F��$��1h��Җr����w_��P�VhK��̽�?;�c�j5��y6x�\<��<t��#:���=W�կ� �H���!8������)�-[�|-��eK.�J?��l��b��c��]uyZ��x��=��;{��Yv=4�
��*>�vs3C��F7w�c���ifܺ��{
��4���I��u����i�f
VQ���!���<��1����MM�4�q)=�:���޶9��uK���+Dd�8���i>@��<���C�b>�}�9m�Z�5��x]ɍx��"���4�1�~�� Suwus
bˊq�h�5��P.b �s�fZ�O3�jhǨ���хp�֠�5 ����b��=S����]���(X陼^���f�G��=x������u�+��,5���"}�И��͏;<r��N)2�=s��?B`{��9j�Z��#�:����]�w����g��d���x, `�����)�J}̥�[����+��[ig׈]螷�DN~��9�t�X�'|zS�z��]�
&���+v�o�.����!��H�x���5���ck�#n��o�w��Tx��<��1�4�!r��ї}�EYY*wMw���7�x_�`�c�Z��_y�%�5wpΧ�7z���8w�{�`a�1����.o�� So_�D�I�V����Glz"ڃ���mg�D]�֫F�iB.8�˪�*�e�a��{�ւ>�9A?�^<���4s������yn�}�[��7�<�)�(�[���@��&�vc��k	����@
= �_(�Z<����n{;x/�/�վ��̡d�p6�x���h(n����tt�6�E�4��"���=�~��R�=���rwg��v�h�Y�����{�u��rm���v Iz���ԥ� /��M�w�} 1�矅�e\�Լ�3�����
1�7'�z�����awFD_�e7��j��5�^�*2�& ��x`\N?y8�:�����������М��#	<�j�'���b�Qmѧ':�Y]�-=7�7۴��������q�ž���^��'ρ���NG�B�`�=y^3Vn*0�,��|��.���E �}�Pb�}����|'���☫�� ~��,S"�����b�0��y%f�����0�}n|�N����Y'�Q-�{�Ut�65��~}��%˃�6���0.(P�Uˇ�N�������q��P<;+�t�l푑N�dAJƸ0l��CT*�t a��{�x��WJjRo�ar��J7��_f-Tb�ԪA�N�y ��곡;������mF����O_1��`���{�k��$ݡMa��DYh���ڬ-s��}��3��������+dOl\>��Z���h�W/��7�p�c�}�xo�xNR���\I5���b��]ldWWu�XhU�r<0���D@�@\?���ذc��p�/������W��'/������ǫ�!"f7�x=���kwn�=[�$��x>��
DK"t !~����۵�L,Np'��b���w;�3Ej��+���m��qQ�,�ώᏯ�4OJ"���9@��h����H�c�Ӥd��^XkOx�P�|���_�4=ps�v�A���DB���A�z�m�&���G^�2�����2�l��j�xD��~��Z摕�O�0�����xz5v� �Ph��c!�Ӛ�m◖��_-u� ���Kt>���� ����=�z���S@[IQf��M�%�������y�Vw�Y�
L�,=(�y�6�{�X�&���qP�v%= T;&�n��£��*�kjG�.��;�E�֫+u�x���������y�"�_-�}p����x��h����f[(���U[����ۃ��C����iJ�M�Y�~��1W�y����?7(�����-�1w�V����t͉n;�t��go[����Y
�$�-l�\{V�㬙V��
T��0��K�Ҋ�ε�ek[W]�r����HuS��6\���1��@�b���Uw��T峎�,6�Df���ّZ1#d�e����,��2��Pv�_�M�)��5~���w+�L��a����@W�> ���$�;<[����-�N��O�MU6��y?x���v�qVa��C�<���Xg7π_��h��������=5���}��)�M�%xco,::��k� &���A=z�	`y%X�J{ TW�^P��f/��{L�cv��z�+x_*s�D��D��$�K@t���Յ�c�@�V7=����}B�ǧ���N5>�q�.���!5#Գ"d{�*���N��>��(��~��pE?g����K�s��*>no@}ժn�\F�4�5r�s�mf��'H�:��CgO 6k�|G�>X��A��
�2�^?%d�1�G��]Yt�lu`� ��6��t�V�q����o�L����x|�l5��o�CuoCg?���V1]�.���F �=ܟ�8�>�3��8�
��/N����M��h�9���X�)<'���ح7�5��K}�"z�(����E'�_�@��ZUCgw�����o^+�"���/ݣ�� @���ŝ�TP�B78�]I�/���a��æ$�+|�>���Y5�F*�.�!��b{�<��w�u�߬�|�a����ݮ��_"/��|9������0��ޱ�pKR�/%c�C���\���I�֝�[m�e�a��B�[&���[Kl������+��K������)�4i��@$�%gw�k��p
�$�?��@B�?����p����P��Q:�P*<Z8��M���uBd�ӯ��;�f���#^�ѵ�d@���Nc >��xcҁ����M>	�۝��l'3Z���y�m�/X���Q�*.�� �p�*A`8M��Ԍ�{�4y��;!��y`h���z:��l�0#�9�_�=�y�d%�'�maǢK�}�\�P�^���k�gNXw�8(�by�3�I�������^�z5�3xv\S<�H��
�JR�=6�/w"<��8)��6f{!�>q�e�F�,��N;�8m�Nu�yC��b�R�<�dܯߣ�s��[��=C�k�&��≮^�b��{�wx��~=#A�ˁU9��҃�PQ��)��!�,m͗�:�dgS��-�Zn7*n�����}���o<0�~h����gAŰc��v_���ͺ�KRF|9�B��Xfέ=�Ж.��)^'.x3���*�2��~;>!���>������ ֋��r�]p�\^n��|�� ��M�z%:oX�Ú���[�[z�����[��>knnO�&<9��(T.��md��p�յ�G5�~5q��/����r*�%�iy׻i�vgr7f�2��y����Hk�;��#J Y��A"��}�xd[��^W�o��u�
j��-W��k��H�''SX����9R�z�P�]�ژ�ؾ��^�4O��߸x�m7f��ݶ���[X����b���PK��3��y��3']`bYs�� SwwO7y����O�1��.�-J�>��L�29W�c���M�NG����I�O����O'�^[�i�� ������t���{�Ywܳ�ם��q�!�gLm���+���\J/�����)��t�b��bl��|1�����c�aջ��5��zc�x@����Zg8p�|6����y�m}{���L�!䂼��ϳ��k<����!�&^fez§�Q�!=;�9<�����^��p�ϔ���OᯏK��3�ʄ7Z{�F2����r�:�� UR2�Ű��8@Ǆ|H�
�M(��L�B���u���N{#Z�ʠ���4����J!m�ᡪ�FL`Va>|�W\5���䛩�ss����L��i�?<[�k��Ҳ�1�`�,ohn�,rngM]��H	9�z0[�,�}�Ǽv`�ü��F��<te�	|>u~ZzC��d[bv
�����L5��;����y4C?p��}�7�7��+Эz)���n�ɤC�w=	z���	�5�I��8���0Ae��l^-��ǹS.�L��;�ۼ�<]v��|)��[P�#�{���;��<=�3n5���(����L͵z9s&�6��m>]qWs9�<�r��6��L�mc��R��6�GZ��0�i4�JEja���n�k�;��.A�����hi
���h�󼯆|���������z���'1B��ȧ��������* >�ޠ��K\8LU?oei^ ��cݳl5��[A�6s�� /@�I>XB��N;|�y�x%uJ�UKYř�S.�{�8J�>`ސ(75�z�@�>d�M���V惘��Kc�t.8x-ك�Dq�67�W�5w��o:��۟ ����\����U�q�L��On��ҝ���m=4��Zf�x=�
�* �:�4Nr�9��5��>X��>^�ϼ4|}ܽ��3��������]�f�R�4Օ�=� ؙ�3W<��~��Ե�;.	q ]@/s>(�e��3�\�S���6��]iw���n!����;,|� ����g�����|����a��?��H����\���ɞ�������5�gW�׆�4��_���!�k᫂��*��	�{�����<�le<�Y��Kg�	��$���s��e�(%�s�L��=������7��S�RIl�]�rv�n�׀��¤/[���e^v�#+�P�2[����*��9��T_j=&B!�QA����a;���񕫺�u�{�n&ҿ�x��2��OG3G�U�k����-�a�Ϲ$��ܟ/:�H3��E*��ֳZ�F���ǔ�qKtt���Z��9\�oJ�B�	q}y̡A�c�	���j{��0wI��288�{,�+j�w�Y7��tR�&>Uk���-�	���F�v��t�;-{Vj.�-�/-�m&��ȋ�C���j'�V��g�n�[3DRT�v�ƺ�^n
s5š���I���;$�;8hE1���y�
4WP�^�u���L�Y��}�ƍ���Y����ܤ;�y����I�^�hu���[�M.��<��ɰ��N��\{VU���wqú��T!�[Ĭػ����e=rDԬ�M�����l!�/y�pun=�X�b7�`P}-Iݕ��r:\`��8;݃.�<��;$z��늠�<��{{�j�ի�_���v,�Ol.��ʎ#u��a�8v�0pʻ�KW� �e=s2nRAG[8��R��s"�)��#�I)\l�{Kc:=����,����f�m��G�_by�T!���6��cqfmGY��r�FsĈcm<�X���^#�j�<xYƶ�Nc�w�+m�I�T}Q}��v3I���H��ؙ�+����=���o(d�8�Lo.ݭ�C## �4�U�4���F Aw;�3fZ�=`a����BwA+�c\�Ͳ}�,E�~��Q�t屮haB�$J:��,,��XM�{hf�>8�i��΅H>�����S�c��[ь.��g[A�g���y����zk���	�bm_Z���}����l���"�m9�6P���\�wj#*v��<�go`=�Kr���PߗۭG�/E�rռ/���0�:�yC����vm�t�p�h�3�a[��Ms�VoF�)��7��f�&]̨�!v,lA�q��R�n�G��>�ʌJ�V:�S���.˚b�N�50�wX�x�f����5�<���u*�X�����s��� Qk�R�0�N��
f�B���T��5
b��EAp�u�������/6�@��V�D��9��6�%K��9Gi���V;�gU�S��
=�f�ݼ#@��i%�9��둏��7<(��t���7��lA����ݏ��q����5>:�s�ď>�tUe�lޓ����Wq�����V��O_P4v��p��-���W��y�Wd���3�'w{9ݎYD�[zhu�Yb.6n�t�)���GOL}5��Gݷ�M��^5��F��ލ�Q�ǔ��φ>y�a��S8mB���W�db�Q�LVWb�*�`�Cm�۷��+��K���v������F�v��7�b�./�&���yQ��Չ���������7~L��	�/}x��e�v脝�y������$$�:x����׮4��������Ǐ���ݻ||&U�T$��ή��wv�wr�$2�$$!#���^>�;x��o������=x����nݷ�R��D.1��ۉ�I1�uV�Q�*H��H��v����m�������x���۷m�I	R���Pa$9W,��`���D��r��o/�t($14�d�"b$�c�졄CI�(����xL^� $$Cwr�0b�F`�{�v�m�%}.ѯֹ�A	JHD=}��(dd����7����#���Np%2Qw|��u���f on�?n��s.�ƐBs�`D(�1��BJ&,���ɒI��S�R-'���w�rm �����PL?�0���	Ę<��P�A���Bi"�ĉ�V�/~iwf�������7q<&�Мn\�_i�,w*!�]�m����#�C���ύ$�k��Tы��(�.�nD�\JG
WR��*(�*3�3���bI�	nxb�&�S�&��$H�q�i��ˌ8AP2bd 
P��J�.�X!�ՔZH&�"�I���9�[�4 SCJ�42��T�YVE�\�������{�O�ɻ����3]������ngq*�l0;�UR�$ŕ�&�ڼ��ЂIR� w��_��(q�S�]^1%��}n�AF}Tΰ_-��$wm�s����j������ �>�tp����U��俘<�����a9�)���	Qf���ܞb�7S-��Ͳ�k`p��#g��Qc��4���oDc��=\������t4�' 짻ӂ�ET�ORv��t�����}�H~�`�y��t����x._E�08��5F���:�]7�W�#��+[�̶�xS�3G��^�� v��O\����AJ�i�`ނ�.Z)���d�>|�I%�+v}�����@�)��#�{�f8���u%��MK�x5w)7ֶ���zx���2C��������6��}Ǧ"��\�F����\l �MV�K*�J����Io;	���C#Y)��i���3�xo}���C�!�sP0�{k��ׇ�����eWʘy��z�xS�N�]�q���:�w���f�	�z���ܪ�7.Z��������Q�����?..���w^Øy�{h��_��wt�w����|�3��de�(���:x�������?��rޛ^��}r�Y7���⬷��m��G��se�{����ٕ����z8��I:^t�x���&k��]D]�WY$�$i'��j�#�����л��<��Ϥ��P��lfu;�y�S�ou@�[en�{��9�uC�u��q�YӔw3(ߐ�Di���hh�����)��~g�}9�ψ{�$�Ri	�b�_1�\�ܕ/M���v��1�8'��p9�b�FL��W�7^њcT�����1�d����'¢�����Ǿ��`�%j��8��9<A|W�wh����Yu~����e�R��{Mz+7 ��O�u�ª�z�H�0����ʸ���C;����5�q�vC_����v���m�	��4s�JA��N.��{�0�0[�{�=`k
�>w�3�ڽ��&����:�C���
�,Li���@�1���IO�ar������͢���p���D�3a�O��빇���	~��� {h�\��7��sP;]@�Un���J�y�*tw��oú�
z��i��&#��?��o�i�)���0`v�ob'�+ä�捑s��ӵ�T��צ��#�^*�Z��	��-l�ǅ������8!�8b��kY�JyMgN:��ü"��팖`�p3���f.y��)K��Z�*�|�_���o.����;nC�chW!�zr\�oMl6��yj��S��^i��t���@�o���������w�w�;g,sŢ �R�n���m��h�焓�}���=�*���.��%x�p�3��@$�M
���=��۫{�0��G�3�ࡼ*�x����ے��Ʀ��4nj�k���4�r�p�݃%]b?���>~@D#CB�M"-AV|��� �Sdd.��`��.Z���<��o�k��!n
���z4>�q(3�Yt�l��F�Q�����{��/a��%�.`D��!]���w����Z��+>�vqfh�68.�1woe�d�_���HNv�*����ɪ\R9��,EE��d	ϐ��lo˚r�ݩJ����WQ��#X	ė䣷�8�'��.���U@Y^R��|}�ϕ����9g���:k4e4��k��G�n̮u��K.%��t_��G��s��nex���
Dg��ѩ��w��}׶�*�n����z#sL?��!H�I��LR~ag�y?��}�h
{5����F=��Ǹ9~墆ǡ�<�͵逛f̉�+�ĜR�3���p)��2Ɯ|ѳ��N��߽ͣpMf+ڞ֬�P�5����Mq�xcL�7C����T.��R��68aW�z�^���wvy*!%�4�z1ܽhi�iur��t��:�A�-��� ��3�Θh�����T�ġk��BN��\�	�;X�� P�k�c��8�}�4�4;���LLH���D��q�&������fM�&��ܩ�LE�0���	�+U��ډU���^�g�Q���f�wO	����/+v���|��MCĜ�zG�5�1�J��7 ��|nPBpb�� ��z6R�ULEW�����iP� F��ZhhTJ�"2��o3�w~��xs䁯+��]��Z�]�V`��#ӎ���-����2 ��ϙ���+ҧ	۞L=qx5��L��zm�@ޑ\�שe�|��}����ɟ`�)�F�;`<*�Q��y���ff?ow_�^��C�B�!��7���#'��<r����;���)�) �f�f�~�h�ѼYa=B��a�fz@��.qxc���E���qի�Gg�mpEn�`b��V�am�k��t�8h�Ԅ�w�CP�0uB���<<�
�����ً���
3��o����
t�t�n�� �s�{g�2)�����.=<�H��y�m9̖���O��H��cT�nk��O9�R��9Fc�M<s��ס�C���治%�5�D&W�f;݌+�ב�C3d�^� h�87����)������A�Ƣ����d!u<�=�TŤ:4��D?HP#�X@�2�&9�V�"EF�?2N��?%Yp�ss[4Y�������v�s�v�Ǖ���1f5ϼ��Z�a��E�.$���|Q s.�
x�Vu�-���v.d--UȎ\N׵�@���[]A��)�qpd��wH�1�Y����՗
;�k��z�DsB��~MQ0�wk����K������Q��	�X8+���֕s����l�w%6
u4e�uA��+2�N�fV������C@#M �QTHQA<����4�A62>������owG�e
�wS$x�$�Lh�U�Y%��Io���|��?������qb���>>/���ʋA<�p?��=+���˛���8dv�YC���`��W�j�ޣW�(�sW4�����}��������ɮ�|�'/Ω���=B��e�d�n�����{��� ']�^��Gd�qw�sx�-�:}�[٤Y�̒�&������퍔Հ=�/�y�r����w��3��{sC��5]��x!�7��w�=�1t_��M�5uXm ^v��gԢ5�	�}d����̱K���pNkOE!C�6Y����q�ǽP��Æp�uy�T���z�n|�]{i��=�7k��Ys4�hk55VK��WY9��{Iord�ɸk�w����= R�-�#z���ok��6���}��sU�&�V����� /�>�֪���8e�;2�^�îwij�Y�6����}�f�F���{�ڥP�P���O)v�'־r�O�f��'�[{5���w'�W���s��m�n=2(E5s�q��Cs������^k�a�j�`[ ��ӽ.}
O!�z�R��ׄ��bS�����i�j��R�+�9VH,�Ů�����(��EY��;v� ����@p_���>7��ЏR�`�����ݹ�_k���$�l,и�����e(�E��*'ՓeN}o���ٹ7��}��L�l�8}�_�� )��)��UG�7�/;��|)����\��.�n1�X�7�3��z9��1Þ��2ԕc=���q�E2�ט��ܝ�����ܯ��;�`���.j4�O+>2�:5Đݎ��wYT+�m��(Yɾ�y���a}���YNڔ����y�Џ�R��� �z`]~�-�vf�{bj��Z꛱-=6�# ��t�8���Ng]���Ξ8�<�� k�}K��s�0�Uw{�:c`�٢�#'�zzUX/Hf�+�\�;�P�1e�����}������ymr�4$�FSUM捹<F�N0v\)JmɎNS�qu��7��6��f��-���Y5�%��m�r�:[���ڬ�B/����m�x�9����\�=�Be^����
�Y��1;�mݏ}���"G|Xv6<sUD���3��)�+��s��e\:�X_f�c��M=���tՅa���-��x�+�t�!eq���Z}�A^�s|�Fx�A��1�Bƫsٗ5��ټ���z��Oe�=����)���@_i#b��4O�SH�����g�x�x}�h�y�oO��"9Ф��x.��gq%[d���Z�h�Q��o���׻�Xy���d�+��T�9Uw�"cF��ף6G�Z&SvOwst�'Xy��"�}�g��o:�u����q�ǹ����� ��"��
LPT�k���=��֯2�«��{���S?Ì	�J�i`&���:�~}	��~`|�nPi�Ϝ{ӹ�xq��f�{fc�7��(���T7�034�{J�3�6�E@�t���C�@�݋펙�d�vf��}�gяwjR�
+;�t��n��̐K��1J�-�b�O��a�C(a.� �vF^���k��`��q�g~O�5-C-Y�u�Lޯ�����f��`�w�5"}�X|��ST)����=TJx`�EH���t�[`b�#vށ]��}�`�ݖL1�z��*3?���l#��˪��-�K��7���Ѓ����U��q9S���Ҳ���M�����+�"yϧ�PQ�o���"��ۂ{k������PlDFW_5F�M�p���G�Q��U��(���Ѐa���
����cU��+I�������n�Rq٪�S0懮��V@B�z��g��c�u�c�Suwus/E�UDsɗP*4K��r���hpB�d��S���]]�z���۱I��.�)�=Φ�{L��^��B��}�w�ș��k�۠ҮܩY�tr�C&�:f�ףuGoF:�+=���/�Ѝ�	,�����XHr\Qv��T��i]���EJ�G��ٍr_hE_k�R���NR�r1���5·�6Ρ�t��lm�J7	��*M(�44��E�PL�y�'��~�3�k䁴Ң�y����C�r�	�s��C���O\���z�jI<c{N��Zw�s>z��Hg:��\�p�����4�^�Lۜ��ƽ����|����r^oe�xZ��鵔	z�d.�jw����lk��[|���VWٴ�z.o7_j�=\|㟣��9/Rꟙ�T���M���}�R	��t�.�gsfv�ǳ�|[�_���[��+���)�1����S��^��-��3�݀�f��X6]�z":v����wb�ϒ�ϖh������.�;}uүG�`������=�,�]���Z<�,���u��������uj|����D�*�;HݎO@���/:1Ef�������.�\��4k���z`k��&q��Ʃ-�t����l�o���,��aj`X�	���x�����<�����?� b������o/ֶ�}�l�[/�5=�n��+װCu��ܶ���9�X�����o
k;�����O2���b�	��3R]�Q����@���{��O��p�%�������+ymٶ��D��m�彐���/eS(sWa]��z�P/����i�V%е�v"Wr���o��_[L�o<\j�+D�o�q�B,�_����������i`�{r��'m�[��&�њ�9����6��Ă{�F��k�-Ӻ�y��]��B؉y�g���-y`�޹�xO5ީ��������ݺ��xO^�.�)��c=S7����</�!T�O+ )��oG� ��v%�{+�u[DwH�HՑ�ĸn�ϱa�����]�s���s��>��oc���>~�d���~�,�y�ey)e�"ŸF��p�^=�Y����}`S�=��&�z��$W�/Ao>�U����ܩ.ђy~�U׳h�,��v���cp��:͵"m��*��nՊK8�y��T����n�ls(z���=� ��-#Vĳ��2� �� uaQ��j�}��]�U�� OQ�Ȣm;<?J�n�shUz�x�W݃��W����ǖ$�4�gK#؅z;��|���S���X+��{b�s�u�;)������W\�����n��~+����wݙ�h�~`���.�=||���iK�
�sH��vC��
3�3���j_vf<����Om���z�=�� � ������ʄ�����f�{�m��Q������l�œr]�����-c���1��Ozq���"+��&&�(��ӭ�s���+�X�eYb��
[4�1ƭG5u�-��nڸ3�p�3n���Q�����$�ܘ��>�3~�����e.�L�
'_��T���R�E;�Y�r{�[���]I��ϝ2�=qcY�&�^0R���>�X=_\ά^C�)]�I��ÔIyI�C&ԡ�G��tJU����ұaX跦�]�#j�u�\(ȭ��Z��@w������m�����85���n���[�y��[!��(��[t�wR��>ZÞ��x��zl��/\�L����!�b���ş<s�f�q,�ԩ��y�W����=�>9ȮՐ��.Yy��f�|>UL�Krm�9������=$�W�l�P��Mz��N����ϐEb���������!��;	�m���awհ�;�����awm��Ӷ��_+�|��^�AU���[)����4�2EsKs3�N����7Ŗ??D�V;����{�5�N0�λ/�6t����W��������^h�)|�|U�w�A�����k���)�&G��Yzw�xa9>�eKW�V��L"�-��ܾ0B�\"y��&�KHܩ �)�?p�u��g�Q�O��6�{��=���[Ԗ7�9�7����b�����M�;�}u�^Qz2���zs�N�W���t�n�(�r^Gu�gge��.a�w,m���ֻV�!�;uR��41&�qU�Q��obwM��E�����E���l�vr�{���9���]�vS65��t����L�DA�-g;۶���wO�R�{��S���}��s&_RCn�y��\uaN�Y�Ԭ��P���*���DSW�n��;��9;�V�͹5	��ۦ�� �}�'��wҥ��jE������w���B�VfPy'��ݷ\�b�������kzֻC�V����W8	�_��n]������9��s22H�Ѻ^�s����]e
\/���H���$۫�,���[H}"�;�W�u�9�$��eF�F̖.r9�=h���ۛ�8����"� �b�[���{u7d���z,m��Ńf��[���ecꓭʡ͗�r�<�V�y�%����B�q�]3���ј*J����r�sX\7e����U����Y��7׆����9W�`Y++����uK����u,��v��O�S6Y ����o�k��E8�c�dY������u5�oiM�v�3I�,�|�Arړr�s�޲�SU	(��Օn�c��Ό��u�%��Q������~Ane�n��;��;R�6�;�[�.�R��J�3�ED^%��6��D��DK��޺zF��ʸ���=S�&~.��g.�9f읊L��P�y�^^�gPڏ�mV��H�ű��c�vʕ�"���xf�g��7(�곫n:6��Wm�Iě��uٳ�6��Q�pi'upe�R��U�.�^�gh"\����S��8Fl�e���8��{uVhot|�w'˺�*5�-�ܑ�}�
��D�gkduetX��Uw��Z�q���tK�L<Ф�T�ۦY��A7��%;h_-�d��f��q�R�i�D��̔���#8v�Y%����f>ɰLR�Y��n>X�ܣ}��(;�;v�����mo4.B��)��CJ
\���6ؙrd�$�4ڮ=Y�t#����"�2ie����6i���i��n�3��1���N�-1Q�`no�v�#��%k5����묩��(j�G:��\��+U�քܼ�3�'fL��+�8����C'���Q�j^w��N̫��:g�8�Av2A�����7��u0J5���`խ�{�K�NR&����|���Ч95R����wfl�S��%{f`E\v;ogX{99v���r��v���i����keη��w�t�3��fG-UQٹηX/������]���5YS�����
En$zֺ������%	��/ݪQ.B2HL|t����Ǐ_[q�}}q��}}v��.�	$���霺1b0#$��;�M�;���o�o����x���q�}q��>��w�n�����/2A씈����ק�JR(�߻�~�}m��q��q��q���۷mߏK���+��g�r�R�������}��E%�3F) �H!Y����F7����ݿ]0BE��gn�"�.J~j���y��E~u�;v���wםB��$��F#A`�!X�A�	-���#B(�ƽ�1���%�L}i��?�%W��7��/���ѥ�A���"hv��b�%Y��#_���o��֌��%%#I&I�\m>uߝ�w��g�Fa`ҫR��~9]wM6�Jn��4��B���XxKhD���7�Nw�Vy�e���r��]���}��=~���D
hhW����o�ϙϞO��F4[��^��P ��O0��R��R˞��L��T0��v�*Z'K�l\�̾O�CӭuD�2�$>9�k�J��\�y�6"�$��K�0��d�W59��}��c��#p�&��Ó����\0g�"��!ir�r�?��1?N��C�23���ڹ�ɖݦ�;�N���'�����=�0�5Y٬���~���Q�}bPKW?ag���nCH�l%�
�ә�{@���x��y��ԍ��;@��=zF���}�OoHM���r����ʜ�f�y�f���5�(bS����_{EC��,�-4��6e#��.��+&�w���c��{��g9�� ͨ�� �V}��]�)���r�.���R�zi�ǧg[�����r�Y��_xu�P��%�!�o�@TUj�rմ
�E��H�R}��I �f�3�Z3ۚ��w�Zm{������XYV�tx/yܾ_ϼ��\�"�c.��\Jw�uE��oN�hc��y�PS�ׄ?�ԥ��*�
>O���9�g�lt|3��ο�Q	�H/��ng��|��ySvF찶�_��5c���7ԫFd	3Uz���ڰx�F5z�}9��v,�Jmu�y�-�+���)��!��*��uZX���3�L����M^.�NQ���t����s�ȭ?a����j1�1���9c��M���󄦻� �_)�n������*�̥e������Ng�q�+n���7�8Mw���V���y����at���A{3ӵ��^����}��O�c=�3�ݫ��z�$�����[�`sV�"L{<3�y:�?k�$����6e�W\��ǹ��;�/� �c�\oǃ�5��9��ՂL��cm�~h�^��r~�]��g6s���^t=U�{kd<υ���Y�VS	Yc������u�0�-���Ϛ��*ۣ��P_6����.�ʣ�z�]4���L/4h�̲C��A��W���}�|rO<j��Z�L-Y�.�3�3���~�l�Wu��d��9��݀�Ѭ�1���s�g���5%�նo;'�D���E� J�.��z���*�e�a�6p��[չ9�j!�n��R�XCݴ���g?Z�tv���2�����ӎ��ж�o��gh\��>î�zּ����}��	��C�R>=�����7�_w����4��Mzs���C��xo�Xt�T�/��K�Q�n�ך����]DJEV^U3
s��̳��޴l}����	��{y������x���bN�vd�l���%��xE��q<$²�\�6�&����;��K�Z�滯's�ܮ��ԛ�8}(;~��Jh� .!� ����~�Z�����U�_�v)6��;d��d2�:�ee��}({O�gCE�4�0/����O�zm=�_��Hl8}X�	��c�woUEM��5ƕC!��Y���)�>Ȋk��
cC�z`|}�QU���p���v����z�f掠w�w�_��W�޸>�5!9o�.��#�ʱ3 �
|�i�����>>s���F]��V�>�NUgd�9}�O�O��|�T/�q�a�ܲB����¿{��U�,��������;�۝�}�]��ql��.}��sU��籝�W�@��f=[�dO95�ٶ�l}�ӳ��\�Â�S��4�� "���FF�>�33V�⼌Kw �3M����[��Qv�|:^l\j@�=P��^�z�Z�O�}J�<5����<�4A���'��!�9�=��J~��Wl;7�x̭�իD8���q���'���:�q@��=��a�n��^q�2q��"Ň��VFI�\iQ��̺���XE�����7y��G�F�>�XE9�5�(l��ܭm��9�����/a2�����g<��3�H�[4�L/l(p|�<�]���!��-��ZO�4����(6*��bې�CS�����s����Q��A֟�Y�uU+>#�;�����1�s:m����E�)AA��%5܎c����'X"��v�ζ;Uח)���E�W�p� '�i��B�j"$ ��}߹��:ĸ��'b[��B���x��G7K�9.}ώ�þ5������E_a�n�.��:nQ5�	�-�%�	��/��y�O���|6���b碦�K�a�����{w2�drE$���Œ�	���/|�, v_�W�"���=�`�>�y����u屝��gw��U?�|�[!x$A�A�
㥊Cܙ���BN|̓n�U�f\��ʔ7!�gC�(�m�NY4�����8�vz�v�#��{=Rw*���c�ѧ	�4F�A��g�4�������v�ϱ��:�X���I� �跦������h�⶝�'"W*~����}��+�3�,��*��x��#��V�9jU�fr�g�[g��6L�(OG������֎x��
yiN����pA��Ud�j�|E߶���vSs4���&Π����^������az3�>8�>����ن4'�Q�jd;����Uy�f\�+;���=ێ1P���8(a�8�"��-�Qc�Z�m��C*zSű�\ɣA�+����f�J���l���~�7��Q�Q�ϫo�J�(a�xo���ke��f�Bcͼ�D_�N���)�nGX]yB�o�L��mgZ%��xܹ�7�i���T���Y܁�ׁ4�]+4k��U�gg�F�eC9����~��
hhP�����O=�t����: �A!�/�=���٤C�[��S[�{g��]
E��>[�b3��Ɂ��[KR�͎�K������P���|}�"���g�gO
�^��hSA�(uW�]͕��COT[ ׮,�Úp��l	O��P��,�?z3XP���e�n"���_N��X7��᱗F�F��۰
R�NT��TSr~��9���6�{Z���v���M����`�H������Cɴ7>��5��Q;<�tS��^[\�~�L��&6��f7@����_�3̏�HwR감�/��㚪<�� ���V�Ԙ?'qZ�=�Nmm�����J�X&�������3������>~5B1����5�?|�T-��c��P����\p�/at$�_T�5v��P/lg��O���6s�^���v�%�f��Ypuðn���e0�v%@�s5�e@�,;��10'����6�A����F;c�1Y��j��)���K�OX��7��+���׊�e�A(C�+�l��n�m͓&�V�]����W��o
W�!�+ROy;V���MhV�&wћ�����4���G����hB5�ݬ���r�� ͑�D��d��H�����	R[�:n�E/�r6���ذ�D(0���]�=j+���Y�<�s6^ge�Úɲ�`__�ҥ44M
���������UWۥ? �jF��#��/{$+��?��P��'ΥC�R!�on�7gk�fs[���t���Y�'�9���#��*��j��\^���{^5��C���s�﷣0-o���G��k��R��lv��
v>���@�����W��eAG��cN������}��
n*b��$��C6t�j5�㢘�b�/��h=Y�+��!w"kr�Q��h\��:$Jk���n�||�_>M,�H�cս[�O�O�hn	�ZFi.��-�/,�1���ϰ4J1�8Ab^9���Ra�q��-U�l��t����7�9����s��4=#��A
,u}�ڌx�V1�r�q��O|��O��>�]=��!Wq�"1�EO�1�*�������#]�1�;\q�5�C�e��#��9& ����T�~Y�+j�hj�z�xo�[��p������C���c�/Xt\��+#��94�o2�G�'9K����ˡ2���Z|C6�#�`D���C�O��4����#`��K��Fu�G]��Y�� [�|K��2Y���nkefŕ߱�J{��=���MHX�r�v0��̶�����ղ�銄���J���c�٬H�W�7J�_GX;,�j$�U-�I�=�c�<���ď �(�CB��xV��|��{Z�����G�����R�#˲F<[CZ�^ӄ����>�v0LkL��WR������@��W� �'�x܀�9zK���8��A~�|7�'{ܯ�¢X�dKt��,(��W�е�^�\UR2�Ű��S�ם[�Ww�|�����ݘ�k��o4���l���7�l>�z�K=%���#����>f^sf�[^�'8z;����\��{�7���C^Y]`��kKig�+�;~�YqgJ!�Gwܮ{�tK?���ǼHd�о��->	|n��_��s<j�����Փ
�]X֨�g�)09�]q��S�h��Q�����-iG�� 6*�_��H�.pb�`�E�,�o{�T�h�R���� ��_���8h�,W>S���:\6H���C��Ŷ�x��){�#��*/(�_^s�=��}CݖG�r��ϸ�������.�9�7Q��:Ch��(�|Z���T>p�� [�G���k�S����'����/5��c1͛4X��~��������4�x|��S��D�@�&E�cuOu�N�yL�Lj7?'\�[�wn*	�"�bp`�a�[y���&�U���,Ö�7�+��Xx\�Ս����s��-9�Ru�f�
��wUԽ)v�Ĺ������<��2��<��Y���(8�b��APG��ZD`թ�ٽ�.#{I~��Ès����ҭAJ�xy��=�߿9�s����:�p�^]�'�4�">�^O�2��+`h�P�۟�'�է)44�ꍦ�=����]"���kk��$�p�@Ǟ�m1�"a�n�Q�;�������&���ihi��y��N|�_Wc�L���u�(���y��b�@����sl�;&wC�������=��{�.ӆt_��=�}��Al��7B٦�s�-��5�q����z���ۅr�9��(�\W����%DÚ�4*���Ad�n����s߲ &wvR\�]v9��Z�L��G����B�F�w�	��� ��M����<�:�Κ���+�󺚰����}��w�5�4�`����H^YH���5����u>#a���V�P���#���;njt�i��L���d	�c �����5��r#��/�]��������V��z��"�%�w4�TY�>PZ��5q~��K��F���O�{hc���V�S_�Լ�W
�����j�'�
�d��a8"�P�el�"^#�鈶��_V�l�/�VD;�:��pQ�k�����v��Hn
H�\5�zy/
�؍��a��0��mb�嚮��<>�9 �dݝ�[�&t�S�a�Q�4�ɇp�J��|ݼr�_������H�nu������jY��vv�C�t�JhhiC� �.��پ��lH��e��қ�wi��/�c�6�E-�O@.����^떹r�oE��N3�t�=}�����w���|5�2��"nϾV%�xd�����@�r2]���w)�93'c�y��g3�P���N#�5�)�b���b����v��v��n��=9<l�_�C�;/�d"fgC(V��q��9q�g���$���&�<��|�=^6|z-t㵑l\�V.�|;�fe�ӆX��2�|�
�ԘSPG'���y��~��Sz:��Lv��]��z��G��=o�$v�2i|�b_����+��]�u�8�g��e�����@��]�>�U[m�s����p�!���d}fn�W2�0wY�+ǋ���5��RWi�h>�tt����Y}�oT�u��n��<��Ct�2Zw;�J#�~*-�D��3=� ����i�P����a��� n�䥝�c_Ө�m�!e�_��W/̦�D�9\¨�R/Mam�k�Ss��ռ\��eii=~.xO*��=5(P�kHw��ՑO��y��ܝ���6d���{�ն�JJ���pK쥽w�ssn��g���;���l֨1y���������ާ� �r�0 �(�ڏj��_e.r�M�0��/;jw���q����^���N�:�vE����K�=8tn���$���q�7�y�<�����qi�w��F���"|���I>u
�.����4������,o���4����C'u���x)�[_���F_�=�ÍAmjbL�gd5��:�T�f�e��fd�ݙ��L9�n%@�s5�I���Aŏu/���	� ��}�i���_բ�?xp�am�����n�q��0%�=�J��:w�Z��<���N_ ����UN��Vj.d����߅��N���dXt����a!]�*w���Y�n�J�H��v��g��#{|����S��uo��$�B;~�ޚ��U�/,�+���y���̍�*����i���p�߹֎�ML!B���G���7�]�r�x)�:���%m\�vUMWׄ��c>~zF��!� ��*JV�z6q���:�cE3��X�L���f.쩊Ü��|~��r}�l���29���
�<��#�Bޭᦞ����>苓����R�GKt��^�	!O�h�i�$�;�~^��Ú�wu�9���A¶�v�3QE�w>]o�dw����Yl��u��U�Da�#�c����")l����(J�5�f�5���.�Tk���2&� �2���]��UH�Ҋ�3��LV\1-�q^Z����]��t�hZ"'�����ѻ�6�z�5gmK��6:��8�jE��{m�6f�E��t5��b�Q)e3����z����e�Ga_3�i侤h,R�iؤٽ�ʬ�ˠm���J�P�ܳ��[���J՝�K�,4��588V��+v�'.'r3��4e}T�N��#�w���a�y��и�'Hv�2U7B=�qI�
�\�U�|�/b�jB��K�N�5�{!�X�p��U��T��������G��J���*Ąf�4���j#�q�g�U�Hn(��H�^<�e�^[u���iAMZ1���vl0���*��[�/(�K�g��F]�Ί ȓ{OW^"�W�rМ�⚞=(7ݘ��e_Hyܡ��5s�Qኝd�E��[V3��v�c}e��B�|L��Kdѹ�דE�(c�]�,N�t���)^]y�3jE8���˴�<ۜӨ�n�̆�(����o�֣����;Zϕ_B6���Pl�ॻ5�H9:�e�����9a&�X��[�Ri��׷�r�#�VO^���s�/Enq�:�]��j�%��/�� u�#C@1۔�S���WH�QSu��ge���vAN�OL��O���dr}W�b+�˪�dqnT/$���TM|E_t�yP�%���G$@#��Gv�����n�F;�	=闼������5���͘`�&����;\�|�8n�g�|�Yj�<���ʎm�ܱj�M���ھ�om�z��}ǣ'N�*������r�}]Z��@f ��=��?q>=M"��摈F���yW�8���ۜ)���j���;�8��o��S8G}�^Ω�v!]�[�2���@��1`�N���,[�a_��K�a�_]�ϡ,��gʯnX�0��=���PN�s.�кXJ��[z���e�1sK�������U�*���x�;=�\!ʬ���DX�]�:5� ������w�vxu��O������:��60d܈�-Zz͖DwI���;X��'y�l[�em�s�Fj"R$����}CJޫ{���C/����ә��u[lڭ[:ƕ�bD�&vQ��d�P_J����,��kz���wlN�h�f�wKm�{��˯��>�m*c6����o�h�z�us���na�-�S@ ��Y��Z�gD/=�l&	��C.��[r�Zҝ��Ibnft��|��"y��hU�dd9}�v��J{z'q��<8�d*螙��k%�r�;��R��d�h�8�7tG]�V��X�y��҂��1=w>�J�&��(I	$��$d��qێ=m��q��q���6���۷��$F��*2Z���Db�4%��F������[v��8��z��6��n�/�k>�ζ���E�~v�B@�AB��D�$�=}z��oq�8�_\q��\v��e@Ka B!$�eTx��n�h�M͹b�����-�3�*���k� W�t^ת�����Εː�1�d�ɂ��"��\뻽v�I��k��RRkېj�/�ћ&�m���1�1� ��%IQ�cF��͍�T��sW��F���E,Zk������^1��F�
5+{n�>�Ww�梊4F���Q� /�B��,���F��h�RLL�Hi�\��2L>G���TP4� m�ҒC�{n�Ǚyn�[)2H3}��:ۺ,M�TK�(��Qաh��co&#�;��b����!����h8�h&ʊ2�Pq�aa̍G)8�&B�M�!HB1`"�H@ i�!�"�M8K!�dD�.�0�i8�,�Zhr$)��	�a)�$�� _<8��q�8�
��?��8�~K]7ur~v�`��֠�0��᧰��b������n�}�R�֤�B��WY�.��c�����%�=�"+<�'$��x.W~^��onw�h�W�Wq�a������ 9�`ul$���?0��x��;}*�9�;*��Nޗ��40��M��ƴ?�\��+��8s:E@��gs��5�{OK��E���L���-5�!{�0��d/��<?u���8U��dV��`��T=C�	��u�]_E^���^��	����@�Aa{�Y�w���5f��
�w�=T&%��e��y�	L�{vzR|��k�Uhc�/���gVRU�A}��y�}���(���Ɖ�+]W2z�á9�����z	Ak����y�N�����N#d���z퓐�.xG'�A��w���Ih�x����U���%�X�n��� ^U*ǫ��3\?|P{`�4�8~��h${����;���(7���=��wW�Hl�&����]�$i%S�~J|�z�T�[D��b*+'��E��ui��>�}�Լ��pe�g���xNK6���9d�v�'{˗x��q�9�A�+��Wq�֮=����nQ
 i��(
CG
��+j)���>���Z�okoUf����׬��!�����̢/�p��v�#R�"�Ơj�9����|YN�nI�����hh)�׾w����~R+� z͏|.�hEn�a!.�,��/^���=o-C;�M46MlS�������a��-9�^�K���@��B��A��t�n�oyY>�-l�v�n�iƞ�<f��m��^/@��0/�����g|��=��sW*�55�D��q�`p�>��"Z//����i馞��3���v]����d�ư�ĲO����6vZ��oOm
.m��~y�i8>a�'�\����ms��Z��/k�����ݕ��wޅ�l~�)����;���}�霐q��ǟ�b=��Vs�G�mC������#yߦ@�c�"Z`;�ra�Q|�B��\�ߙw1�]C����N��{����~i|w�u��k�ܾ~-����P�t��C{|(�i������ vxs�/�y��H�`��d9��ݕ����)�ޣ��s0�Z��D<2ׂ�۷�$���xY����})=���Ʃ�{�[��u,���t����g����@B��5����#�F!ɓ+M�ݞ��{�Io�2;�}��3q|!i����k���G�^�=��JrSuK�ͽ敁���+�o6=}�^۬�Y+�R^9{r��D6?���h�뵷}��T�t�{�Tհ�P%4��s��A�e�=�5���e�k�pS�q����ᕛ�_��߫��|G�� ���v��w�Vc�*���7S�9c���H���5"~^�3�G/�{����&�!�QQ��D�;-�i�7K���ʯ��Zk�Y��6�G`�A�@���~,5��]�GVa�^�6������qEp��9����M�X�%:�9d��A ��e>v�H�����^d�����Myw�E�9��ƲCcǎ_P%�>�ɥ(f��R�5��ȗ|]�'gs�4ti�̎�c�q83w�#�bcy������2<��݄���84��iO�|�ⅿ7I`&�Hi�X�s�՞�x\.C6q�l#c'����L�4���	��qCrne� pgE��Z/2���7g����s��F���o����:�@�ڢ+�c�F�y��>��k�꺞T�����`/��%��U���ޡ�M}�~b�>Bq��yY�|s{'��z3<oz��� ��\I?��ؐ�+�����"W=���������� �>1�F��^8A��^z��z�D�-�ܳ�i����o���9�N�ar��u��@����צ��gק,K�+N�:�ג�j}o�p��'�Cٍc�-JW۫��q��fH[����㮉d8lIFK�J�����̡\�6Q!0�����}��Mu�v�S�a`�&J��[�cUn���h�T]�v56�����u�{qwbL������L6},~444�л��r�{}j�����\H���N��`@ݞ�e�;� '޳�W�N��|lXZ嘆>��al��}�m��d{�a�u�2t��lh���b��ܘ<�<�\���i�k�P���:��Rz����9l�z��|J��_<�jd
|�����s�BJ/-i�����R��{���ǀ�DM �9�⤅2�N6<sUE>~�R^�̈��9Ws��w�2�|�G�kO���?}�gO��� ���}`�?1�6ڸ��s�Qs�n��{�4p�#�}`�w8��Q{]�F6�L$e�=�pŭ��a�"=c�XY�`�49��a�1�5�7@|��vn�%�i��~8��5e�b�9^	P-+c�4����)���%��9�����6����wT�ߥ�sױٲ2��^�P��p���sL�q�9.�1�9&�.��=�-���%��;�w��,:v}���B�ۢ�2s�Kɐ�.i���̆��ay��%���'I��u�}��x;���&]�a���N�s1��~w�)���[�]FѤ��$���	��y��zuzƎ�������@��s����8\)n�J�+������֑��7j����=����m��驷ǥܳ���t��z���y,:R,T.�K�{]�r�W#����n/xfe��~�41�O<����Ɇ�j�#i\�^3��'��mΣt�8�aS�W�*��(� �0����L>��=���P����^��X��~�w�y��#&WF�"��wa֬��H��*C���peAe�EB��ga ��c�>�L��)�[���\,''��p�w��źAy���#~�����с��_*f�{�YB��f=���>4LkB�cި��я�3,~��5ĶLG�>A��2������lW=��L9�GwP�����+>�6vz%ֽ�i��
P_����_E��A������T��1���hR�LI��!��9���9����4Yy�<��rc^��	��u�^�oj�7M�n��q��ۂ2�e����Iv�L8r�];u��/���P��u|i q4��������ݧ��NC�C}Iqڧ#�W{g������*/��s�HoJw-^��ׁ1��ϭ�Zx��Ut��w�z����a���a��nY�J�e.�/]���ރuh�^��gPC����iS��;^���77{`_[�.=>h<��ĵ��۰K�%����z{����w"�>�fyR�_��7�F��j�W�	�k����*o!٢�ua�86Ч�f=�J�ø�L�ܸ�w#�u���j��Ijfx���@(�d�2���[�oi<"�b����\���AE99zI���8�Q�.W_nw���<��fE��n����v�^���<�a�f a����wپdo�`�c�'�{�q��`h�ڭ@K,��L{�]��T�q�6j2����SG� �b'�pw"@Ǡ��F�fq��� ���ߗDG�%�|I1۞�bf[�c�^�i���&��%4ԧ��)�����w}0���8~��Z|��oa���Ɗ~�����4���,���碚*��D
n�T9�lK<!���n։�I�LPx��:h����	������{�[��� ]zS��z�`1X��)�i���=Ӕ��8:�ۻ��.{'��Ǡ�4��T(Y^���6Ú���X|ؾ~��n�J�����8"��?;LpR)�a�2���q��U�p�m�^{�<o>�'�����璠���o�c�u{�﨏�_�օ���U�|>B����jr��n��^��A8]�]�|b7q���ҭ��SL���B����Ǝz��;��5��q����`kD4'�����:m��c��d���$Su�kg�c��m{W�
 u��!��G�=�*�v�G���Z���7�v�
]�U���d�\!���oY�IE��� �A���S�}):j`ϕ����&w}�#���=|��:VǑt�֠]�[�n�<�jm=//�r��M��\�B�����.�1�_����y�����Y�&���r��	�W¢�)��ᰚW���s.��EuwR`Z��N��{­�LFu:U=s�g;��=�Kҽ0��Bz�-��t=ޜw=��[7�n��L5�I�lF�:f�s��0��̚a���^Fnu
�fx�,�H��u���4s��w/Rٓo���u��s˾2gaC�c !{R>;�g�B�6�9`d��`^��q�;p�X�s��p�A;3.���Q�b���w:H1��<G���y��?Sץ���	�I٢�z�b���%[�:�>��k���\�¾]�ɔ99������ū��ܟ��(���]����}��}��t܅+$�a9�aE0�%�+�q��0$/U_h��U/K��{�(�K�6�Rʃ�î%�7�r`soW�Cc��	�OEC�d��Y�&x��q��R����/Bn�+J������X����ڑ������.�h:�����H�ԥK�;�h��k�^&8O�_W���{��0jbv�G��S��r�w��Uy�>�7Ǿ�������j���c�}V�d���ˬ�ϫm��-�:��F�v�viǦ3ǀYg����Qa!t���h�]E�^n[`��k�;�.�]�9bfq���.����E7ۄ�"�Ws���j��,S�/u�Ɵa�����<�a�j�x��v�|���ϨkW�LJ���|�����?�߽�9^K㻲܎G�ت�G7��֖�/V��YPIR�{bpT{�4<ë3�#0<'Ξ�n�bk	O�V���]ӗ������l���_��}j�c�W��
���&55y�c/P�N}��M��R���r��6��з�]0��[�)�co��k�C�����������qw87�crm�,��FÛ��#.�W'�jݘ7;{����5�8�}���6Y���̱����m���\�sݳ��-��W�t�{�;���y.�dI�;<���������&��]�=������un��m0���)4>E��ӫg�~�,}��A��	�у���<�bg�暠ʗ:ٿ��9��a�H�ָ5�'�%�J�)��q���(ƺ�	d/���QO�c��灹��u8����Gi��iu&�u!��4��gK���P�Xu�����������6���������+γ}�.��O8���{]	=��֓0k�;�6	����m�����M�蘊�-�6�(�у��QIJ��vZa�� �LO�R03Y��h�ʂ�mk3j�Cl4�����8S�q�n�n�#��۬�;�VA�յ�^�՘�rat��[]��QM�W\�נF���]v�M�;�Q;�<�@N��xxW��{�ZڌMg�~�F^Э��mA�r9�8L���I�Ÿ��]F���J�oC��K�c#��q��V��DHp
�G������k�P'i*��`&���R����W��V�Ԇg2��������"��Cdnu&	/D��P���2rD��W�$�S,qV��~a��$Y獐���ټH1�ų�gY�8bp�O#�n鼢k���4%�����3�:�=���a�����&e�z���鴻��|)�m%��L��kNX����F��q���b����� _�~��{s��]6¦�]z��zm�\F��l�R1�(�Ƽ��*	g���S�^��e�+�f�?O��	~T�n.L8�����W�n�;�}S�W4��+�PE��f�St҆`��ɜR�����w�����Z�w	p� �){�Z��	L��~]�mQ��4^�>ߙ��mM��U���L�@�9��|�/�^�v�cƦ1��q��O|��k�D���[{S7mܰ��k�]ƻ��^"���@�7�`c��s���0�8O	�	�L��f��7{�>�����S�R4�;�Y��ϙ�p7ˈt�33vP�խ����a�7�[-�;������y���{�Z�w�sqD���>A���[w4�i�;��E��!���"olj'�[��η��Ÿ�gSD������y�����m�$�Sw[{���z+�0�.�I���<\+
[��;�׀�M���r#�y�3���1Euvp�zzR'���
zT:׮r�wBe[ҝ�sc�7���i�ބc}���9��_n���Uv��q��o�H��	P��]J^�dkt�u^��d;HOO0�Qq����l�ħ8?��8���Ǳ��9�2��7d�aA<^��I�� u�l���B��n��j�Üm��2s ��ǁߕ��7�D�ԭtU����1��4�&\�8���7�����g=9�C9c_AMEΖX5����;��a1��.��>�ׁ)����R���y�p�����kL��6L��5�{b��a���% Zt*�ς��ӿ*�]X�/8�/��[D�d7G�*�;H݈�D�>�o�"�tR�n����E�>��K��t#E�Ra��+w�8�C0��v�Z�%�ހ���݁w���	���!
�%(H�N�Z]�J2hI\�_w��7�����|�f�ψj��z���)Q�=�<+��Pn��m�7%�ǻmN?<,hZ._I�<�;�˻ٍ�
5{:��қ�>��32�X��F��3su&t��O7'����3E��eh������ ��*L�ms���G3�ݻ1V��t(W?-�/�J�����ک���h����������J�M�׸�m��_ta[\��:�u,�üD�r�T8�7�.��]ݫ}�!o^9Q1x��R��] .�����#ֹvd���u����mA9��[j�;f���f�3��A���&U����vWe���1m�2�gx���ĖR��J{1�i�lI
ڀ�s�v���"څ��Ά����R�i`�D]�QR2����0q����Di�(�����<a݉��L>̢��u���7Q���uqb`��V��.�YҺ@/I�v�C�.ɯbλ��BV��/��.U�d��Д59:������C-\v�k��,f�D����od�଺��YM6{pKᡉW:�*.�,�r���>�/��7k����AT���>9�	����T����í9(gl��@QϺҬs��>�~M.��+r���&�=s7N�i��7ΐ���o�[+y�xWoP ;;�nM��=��ݺ*U�ݿ*芞�.�V�E�%�5l����_f�����P�E�Jmhxkf��� �_bиR�ݼ��h-�OG[W3w�.��Ef'*�\uw�Y�*ms:�J 꾶�����̺�3Ʃ�#�3���t�'}\��i ���g�{dRE�K��	�|�ށS�s����^{{h��Z2�'���b�M۫_q�ý�זV�#�g��^BM-��(w�p��Ԗuw�R�����ߤ9�n[����ĺ�:�	�9}ΟV���#f3���%%}}c�[�3qۮ�Y�ؐ�C���f�`�������Cn��%'b�+;�ҩ9	�-,��n+:k�Gy�	�	7�;U� 3�OQ<���p��;e�7rz��#����� 彔v���$b�+#�r�K:%�a���w\�w`�
yn��q���(ILʩ�"U+�ЬXi�*�ͷ��K���JnhFoC�l=G#��k���7}Y�w\��p��ݟc�r��kP��C�n�u�%.�-��`��ZWG��`�%ó�N�ՙ���%;Q�_TݒH̳1�ި!���]%#��Vc|5�.�zre��8����k�*^�|3g�N)�1B��gs�#82�=�'��^��F����ζ��n��{%ښ��Zv^9��\�a�2j�Qab]m��돺Q��v��}�b�DV�ly���Z�V��
�#� �9r��-t��I���ZOM��&����K�7�Q�k
����nH��̂����V�\ŗ6Df�R�ٽ���6��F�Ww�#է]-�݂�j�ZhP5v�ws�s�ye�:�b�vwQ�h5��N��fGz� �^�1��,�����Do�督�mոj�2��E$I	޻}z�o\q�N8�ׯ�8��ݻll�H�/��hح�k�BH,��*2����}}z��N�8�8���}qƟ^�v�Ȅ�j1�6ME���nBP��R\*
H$�{�]><}}i��q���ׯ�8���nݵj�G�v1�V5`��5�-�=ݷ5{y�X��.Us��э`����k�i����X��Z��c^շ2lF���͹X��6����E���E�{�_]�st6�"ш6�ţ�Qk�~M�+�ʿ*�o��5�h�Bm�����Q�1��M{r�^wL��� F���D,�w*�ۭtڶzU�K���NΦs������@�lU�Va���|!���bX ��*J[t�Y��y�����6�X�ǳ��Z���dS���a������-�Ϝ�'��T��αa�[*,�[���|N7���.ڭaa�z��xOV�3?�j��j�Q��nGy�dk8(fY����|�6�N;z%�u�%�	��UvzN�S�xg��k�10x��r9����CĒ���D�޷��C�t(p��{rJ~��"��������7~���q�	�2��K���}����YmO�,�)�Aou%�����?Fˮ�2)G�����ק���i�|-�Z�[�������Y�l9
�2Ͱ�t\;Bx���Ź>����g<�~z�- ջ�����n��Y+z�G�#���}�@�!�+�x�y��j(}�O,���ޑ$v��~푭��`�=6��c����������&�$�(V; o�u��]#^���w�{[e�1�>9w*k�4-i-uTK�ݴ��T�3wl����^���mZB�|���;Ɂ@;'��/��s8`#�Z*���I�
���i0T��^�F}T�u�>[�}��ۨ�C�Or/:���Վ��Y�j%v:��b5ݼ�Ն����]ϥ���;q�)���S����׹wz��w9���M�	{��{Hn!DnT	��/��f<+m��C;7�s/vm���c�O"-CR���s�`]�|��S6�_a�f�[�߿}�8xG��#�9�4��]��� �~tD3y��}-b����f�P)�-�%E�',�4�q�������d-^,rg�&GGl��+$Hy���&25��T(����W.ɩ;7y��h�OSe�0,���L��-�^����Ave������<��r��α���7�+vRz]�2�������v:���n�ƾzכx5����Y�����H)�͙~<|�}���a�OOG!j}�[�vN�����גϫX���Ī��=�~��z���<�>>n���n��W��ɸi�kk�О��b�U��ͻ���0��Z63��>B>�W;�wF������]#�ׅ�ŭ���47[���M�R+�ORaMH俱�����sӬLr��������񍑴&y�EG64�G1.�㟗�����FN0����e5t�ճ��\�����Bî?���:r�̂�*��	���<��K��k�����iU�%v���Ϧq��G�M�P�ۮ�ŋN�I�T/��5��r�?fD�v�ש�m�
ޥ�j�����+=y��)L��4����2>��M.܌�=�֎��6T���"��^ʍ��BT��[m�c#�W�-���{8�6��b�r�L�����:���=��	�~���{����mx�cu�m�I;5Lq�s�#Φ3�P'�El�6�wp�9�!�ݍ�����؋@�Fh�|�>�5��΃qz�Lm@�΃2�"�6��j���c���a\0�s�P��~�L����<�Bn5�q!��㓍��s>�ኑ�6V.݊�y�<'�t��Jqv�� ���O�˫�~���9D�!���/Ly��t.j|U[��0��8a/�xL9�����c��_�����	����Qijc��a�YM[ֈ2�=����zc>P��੤x��C<q<U��*�a}�Bh��fo�F���'f/��|G���`3W�P4G0>���{��K���f�}I�bS�扖�����
�D�`��'�;Dž���A�q�^B�,򁩱�x����,�����"��Ʃپ�-�<y����E@A��.��-���Ok 38	�8E�o4���x3�pA��[��Nis;�v�>=L��.��f�x�>�1����\*}��ڃ��a��<�*��X�o�/NA�ip�Q k��T�h�w͍���/N]IJ�^͜a"�*b�l9���~�u�V<ƪt�yJ��|̙��!\�󤅚����,�ۂ�r�k�����}4܁�U�.�+g�p��B�e�i���T��6Z�"�m�{հ[β��n�1�=����`�x�p����G;����:�:U�S={����7�{����*]]l�p�M�i��z=�ד�������W6a���}^�ϓ�hk������l�Q�V��e����o�W�<�}0.�&����s��W��=��d+w4-�I���x�R��ט�¿,ZP�f���x�X�Ѕl�՞�#��z��;X�VM�O�<2O�q�n��aNb�
V�e�x�!�p}g�Q�}}����m�ȫf����tkp��>��tÏT�~�1�k���30mv�=6x8���<��ؕ��:[:`&R,Ȟ�I��Ra��Ӝ����L�ޔCX[�$�b�N7^�.�o7��X[	!�7��*��O���CĹ���a.�.c�n���ݐc�n9��_}��ߒN�^���.P��=qÞ�I�#gi0'���	=˸���ӛ7���BX��f
�z���1�"`0g�p;�|h��G�IW v1;7Y=C#��_k������Ǯ�#ӏI7�˰[c�ch��L
���-Y��G�2���t�]-�abx8d��i�j���L�CR��[�y�i����t�D�������7-�C��7M�D{9�]+�ͤ��m�x�_nw7(M�*�b��1K]�l�5bve����Ql��uWE���4��J��_GX1�T�з��;������y���c��<��ic{\ݮ=��顶,cüX`��8x�a���'���$���/�^�n;�NU�v����Jiޒ��O�U)�}��3;�}�|H�:�Sx�8[�-އ,�З�zX�G��4"���z���̸�1���g[�J��=���K�u=z�'��#0ջ����w�}��>��Έ�!gq*8�;8�e^��f��{&uP~��O�AG�����t/yG��!E��u��HO6��z���p�n�q�#�K��ް�oD����^��֪��]�
��\"�c�^�_`��'��cf'ͼ�U�O��8�%���)���E�3�z}���򿸤��k�1���O�#�����m����9F�:�E�y��Q����R������WH�����sp0�\?�;��]�ؽ��sk�5Z������3����|�k��c-��]�I4����s.���LRQ��U����;�:��0l�#�s1���]�[���Ts�zy�oz���v�
s�YB�a�l�J��0&1��;!.w�7��x��2�ua�+TLl�-���nKa�5�{���#	k�B<�l�9���s/���l)ӧ.�3����S�|=�."�0�,5F*��H����v҂�Ǿ��q"�GU��&�޿9�������-
ȡ�_<��جMp�v��z�q�i��2f����>:;��1�
�M{�'���R�|�LuYD?u��!����S"u�O���&��'9VI��.-�x5��qW�@��S�>�U#+��.�A��1�Y�58�~�I��fDY��*O+�'=��y�2)Q���v-�sdD<ޖ�Zd���6�:<��G�zҊ{��x�C�l��>�\�"3���R�;����s4��SC2�J�,�ۦp�����d�y�m�Qۜ���Fǐ��ֽHq�]i��cuW,yD1h/暺����ba^1׬�@��ԙ��v�����/�hA�:-�as�=5�B��8��B7a'~�Ǌ�ͿCo���x���b3��<kT���d�:>bOd>+v}�q�W�tj�Ƴ��6���� V�+`p�vJ���]t}�ŕ�Sk�>b����v��{+�Lr����
�#���Mm^�����$���_���1P�\3^��c&ѵ8��
�(��P���V�ϗ���q�� M�?�tw/�'��y}x^���Bm�oc���b�c/����_��pT���.��WY׷�n\~�RAe�7�T ����`k\�����F����Z*��j�_I.���r^d�}�p���XϾ��+�,Ǘ�=r��殎���.2�S9f���j��fԕxk����q#e9������V��o�|�[��L�������*�hQp�9��j�̧[)��[�j�Exx?�:�8.�~�KCE/_OS~;���?ʇP������i��~k�����8���g���̋��@����C�5�>�Y��2:@�(1�d��P�l`kYk��-9±�qoB�yN+�;f<0�������ъ ϥlئ�}�nչX_tw���d�,Y�_�<�Z�vqi__2�Q'��iQc�,{��W"�8��1�t��m�k���3�Ms
����P.{���2�ǪO<;�܇�|�2�g�%�g�=B}~�vo�����s{����߻�&;�꾺���ZAzw�gquvq[��Ҳ�ݎ�\=0n�(�X&��}"�S��(�>�.��Ʊ���۝c��Z©S	��(-Nw�Y��oH�:Q`��y�\\v�3��Dy��;7]A`�o�F�'3Z�
��6��P�s�GM�m9�ǂo�	ϗ���_[�0�0?�o���'�)�D���|C���
��aSS��Z�ٮ-��R��*6ƙ��Yݯ:�B���3%u�-JȉJ"��'�]ʨa��n��d]���D2.i�S أX��oIƓ�uv"���n�]�j�ye��4w�����<�r���u�����vfC���1�Ms�l��"k���ؗ�5@�DM�N)�(���P���Q)�dPt�����^S9�/�d�Y�s�{�L�)�<��4}�'9��}����㖔__0	\@�i���uљ3m3ׄ��~��zkjj��xm�oG/=wd�*�����SW��V�vL�ٙ]�צ\�*�޹��bz�,�Af�h?n��t��Jצ���U=D@�����t8�������^g�׾tS[V<��<L��Om�Y>}�'���Wʅs�ܴ�=����*��Yc[#���7^�����ۂznb�������5s�[��M���T=`[�~��}�8�-Q��e�A��u�Tcn�]B�6sZ���w��ڹ�>T��[ ����4$��7��Vu�.�;��S(��@D��1M�wW0�1e�G��@���
��d{c����S�s����*�)�d�W-�1\���]t?`c�^�4/�B�L���C���J��z�ʻ�2tow��[p�e��5+=n&ʓ@x�Z�t&[Н�q,�O[={o-�:��5�:V́�Yy{�̸����Bt�&IDv�w�HB��4r���v{�Mk=Ս����z���n�`�+E���L�9�=��d|����{*s0�O�p)�۸@����&�&�����su;�S�c0I��]����l�~��p�ҺO�i��eM#Mn{(Z]*]vF�Ot�]�/5hK:V��+�ݧ��Y�5�K�0�a�!���\� �Έ�{;G�%���ڬq7�zkg-�s����[z�CՎ���`��5�<��h��{jV�?]����Ct����m�k��0����ӏ@%�/�I�~��Ih���>?%a�=�{���g�cB|��,���p���6¹\�~S�|S4������nGMm��}M'��
;04�؊[�نp̅��D��{��]��0v��I�g|TK���-����\4���ty�nVt�=G�-D���^��6���OZe|�x��A�������P�	�w�Xv����r�����ޘ����K*��χ��n��k�Wi��
|��f A�5�,�z.�j�����cnv����z���H��o1�������w�wdx��|���tgJ�td�`kD�M]�(2k�}�S�)�PZ����&�������|]��=�>>�־N�c�3X\r�Ω7�g`Sop�2��,
w�.U�%N��8�l$�}���j��N�C]Η#�*�Ȼ��cñ�2�X"��wc�^�Lы��v\�|`�9��Oy�s&7�B����]SjH��ҝ�����,b���s��y���䶹}2�ؖI�.�*v��B�ͽ�jm����!?��	�t\�wCқ�m���#�T9aެ���G 2�6��uuwwU	����oiz��wRd��� �2wݻ�s~�G�8c�=�`˛��I�6�g��Ǌ�6ʔ�{��kd����̩̆�ƱڴapY�_<{,��)�v�u���D����M���ul����*k0=%�q:�궧��0{#��E�Gl�/�}7�]-�h�F::q!o'N��˜�3������͆�{�T0�[��^�5�z�bx\�����b!�&"dOD��vM7,�*9�94*t�wS������6�\�R]�f�;����%��Q��'c@��V�D�)VN^�m�����zVn5Mv��<�������$v���{��ꇪ��e-��zEA�Y��Ke����'�7p�g��G,�F���>l�f��xO��C��E�ь{�Q;��5E�c�J��������Mۗ�FoS[��i�9Z�4Y�I�5uS�T�q��]a%uN.yP�/"����s�nw=�:r�Ov�r������ˇ;k�]��v릸aS�2sFҧ�{qZ�m5�]����!�q�'[��B���u˅m������W�k�3לG+��IgqլSd�����KH�i��*>if���J�#
��WI���B!�\�����)yX��0Xqu�V�,�PY�,�ˍ	����S�t��W4˚Mv@�V�7��d��KΌ�(WY���Xz������U�*��A�%v���j��٫��Q[�������7��ʭ�&�CL��j�ֱy�/Y�^͆6�a�!����
��M皤�#��N��df6T�F�]ʧ�1	9��Q��_|2��0n�7��k)\��8�˝Õ����[;U���QN�LV���Vŭ�v��1�����rf�������ٵٍY��a��"U2+�㛕;��ڥܳPsi�2����;i�\ŧ����J�Z�t΅����9˰2��3�:w����㽩	����P��X��k�c�]]>˄�r�弄�5��1N��>�ˌ�G�0n�x���^��5n�,˽V:�Y�h�Ie��K�W�/1��N��*��V��C���Dr(�
f�5�����HըVr��"цݼ����/�1���(F��	��t�w!X����u�كO�}���R�g�^YTQiRuC�����Γ7�}כo����zͩY��Jܼ��U�pzm�'��4ճ5j��"�� �� �h5�7�_g�T�쁥�\��7Eᩛ�#�2��d'�U����[��Ty�`Y޸[6VV_(EI7P����������wӈmp���drN���w>�M�E}���2�������-\oy�Z�^��1Qc��Z�q�7�ewA8噙B�-�x��k`ju⬰�6�AP*���؏>�8S3�^%�9�����}c!ݗ��; 9�W0�|�8`�-`qq[�#��1d�C6�F�r7Z2�!�r�2d���=;K�x�#��&R۱{��p����}s^��m�y����+ ��R<u�o]�Q˜�9�v�wpI˫WUJ9��9�XHPj�aw����:�m��wQ�3*ZO��oX[�qoKX她HT#��:5{�R����}���g�.�O5�E-Z��f�d��U4fZ^��w[��������w��^���8�Y&��
��j�z���ŭ�ǭ�uF,l<���M��'C׹Wf:�l�� �kuE��Ԙ�u;�c��:Xν]�(]�"]kwu�G�mKyP�e�� �y��gRGVVRJ�yP��5���آ6ő���
� T�N8��i��q���ׯ_���N���B$��,� U�lZK-�Z�߻���{�;x�8�z�����ӧM7 E��\�"��b��`�=�]+�勎��N⧛���o�x��q�n8������N���z���x�6�En_��h���zk�sr��r���kw���`��m�m�h�xۖ������m�b6�_���j�o<�m\ڍE���\�r5|W��v�\�ŷ6�՚�נm`���6�sQW*6�ӕ>�����-F�X�sQ��l�Tk\�wu���j�r������J���¢�&�mH��˅"b@"Q�"�/���1�����d��PO	A*ì��w+z�c2��vXH���t�n��m��V���w�I���%��h��ݝ[�;��(�:��d@�܎(A��L��i���Z�QB��� �b"�I2�+� q�I ����hB�<J����2�D���8�f����i%m8d��M��C#D��|�p��9�������Y���8�dt��5*�qy�š2&h��yo[˗��Ce&yD;��c�ȟ4y���4��)�VO�f\�B��܎�9KBJ�ѫ�0�@��y<�Pؼ�*���
P�|��W0���ʂݒ_:�2������8GO�Z�M�n������;���7`:�oI,�kn9�mOjU"��&�$�1F�TK�L��q��R���i�k���p�H{�##�ܚ=��4)���^��}�kQ��KbQ/��4�ث�����:�0.�c���
!�Y�t1�Ar�q����C,�Yw�W�/�n[�́Y��0�V�u,��s��[�����sm������Ӳ;�����U:��pQ����F��5j��ț�}�3I8�_�eJ*�m��\�ϑ�,1٥����Q1sd�e3B7آ�^4F�F���9��wv���á�)���VUk˩����+J��'�U̮Y<3dn�ŧ
��Ќ�/�ga���/wc�-��Oeog*�m���3�n!G�F�=#�P�~T��}�%��M�=W�5[t���s�]ǯ:�}sY�ܲ�.�ǯFk�0�NlY����+����gG�o�� 7�E���J�����L"9H���`�){�gL���6U�n��(�9�����8��e�pÌ(Y�jzL�{4�h�������9���K�گ%������MҰ=����#���A���Q�%nr$'3��q�p�V�$NE��݄QY�,�� ��>1猳@@]B�f>:w�6�&����Y�>�K��Zex$�<H��y�n��;�Z-S�Rg��vQ��vf�<����U�R���l� �GpAw6�`���� ���F��hxU?}�vf{/��{�9�� m�a�.��st-�����Y��$a��yi� �8�
���Cvf�'����3�=��C��aP3�gz�pR;+�wc�\Q���������!�
��>js��op��(�ۊ�*ze�ӽ[/����7Y�HT���{pd�%}h@���Pi���[4�+:��"`�����k p.����B��s��B��^̣�X�^��	��C V�Y�����
j�ZQ��s��tu�XN�לRn����1��iuI�S�R���Wg��皝/NQ�Y7���0cY�^��2��^Zd�׫w��7�^�� � �X򏜢�qܲ},��<h	�����o�!�i��[�0��e$�9�-t�#@`�R���3|�YZ��a��yt����^IN��=\���vn���M-�ݗ<{�"M�����oN�LB�ݳf�%i��i���,���1��[�omG��!�`0�n^w�rw=�ʒ�u�M&/Y��%�k��͋t����{Ō�M�����a���[RZ8TGNVv^v�`�i�v�$UE*s3s��>� a�g2��y�8�WY9�zY!�+%d�C���:�I'V����Ag�~P)��\F������fɇ���31�Q�q\�\+Gh^U@�p Z�l �Q��6�<��S٥��zbz�.e-/.�z3Ot�n��v�K,�c@����ͱP3�v�[�T��$��q]^wC�Zr�} ��[Y�]�����݌�@��;�+��M�%���;�W)ʑf2��������:��eT��V������C���r��ڶ-\4�M���$�ʫ��i��~a��7�1����iY�s.�aȭ����Y*�q��C�b I�AFҁ}�-��A�G��aD�:�MҜ�~���������@Uʄ(R*�;�ر�"�����qܭ&`�̳<�ASYƁKZFm��G��m3���{��|��譮��@˳�K���+pY��ŅuZ����WB�����d�z�`�×�E���u2X�('ok�4�R��$���v�ʗ)�R��z���Ad�u-�5��>�����6�H��7b4`�x�����ۛ��0�Cm2��	�5��LҾxp���:kk��&z}�w;*�e�dk�vͭ�iT�Y��lǍ�୐�k�fd��	�Z�A�gxlO=M�e˾򚦲ڎ�������l�rzIc 5�~CL��'� �q�zͮ�2k_37 ��J�I�Ի�+���oS�P�vy<^"=�����z!�Pz���eI�Y����oْ���W�E|�cir�4]z�磬Q�J��٦Yta�^�u� Cz���ڷu���ro�~C᯻һ�Ie�s�w���2��*mw_%�v����a:=Q
�n��NC�:�AA��9�,q�z{���xxW����~q�[��+BL4�o�7�r�n��3u`�������J��ꎬI1��e\(�W��P[��Cw�Mv�T����oM���3q�l=MOx��*s�˞aR�wT+�FV�����we;ed��ڧ'�kO>�w֌yg�w�i㻫�;"��m�mx�ʠS-H�(�w:�ږ�VM�
Ct{7���y<h�g�����ͣ\]ѐt]n��fXӸ/����jN4��<o+��`�;L`�p8���:�w��+��`a��[3���2�v=�-�P\���������1n�E��8R�����s���W�'�]�l�n���\ޥ���>�����*Z�^�ʆ���~ڃ5\l���^�A,����5�@-�jRKQ���K�>�����&��͗ӓ�jH8�o��UXu^w]޶Y�^ѲX&Q�|�P�U���.�C\E�Zx��Y�^2%Й�<��:ߌ��zŞ����v���p��u]0�!����{�kZ�;�����*޻���J��'��%%���6�>5ӧv�y6�\��;_�%Ub�
�b��a�V)�(�M��2���A)�1e�Pmt+S)�e,�.Ҋ���h�s|�vc�cw��z�¼<+��ޑdna?}49%��m��I��s�-�t[z��T�M"Gi�1���b2x�Ӏ�o6Ww$6w�T-��_����fm�̨7Q�7N�<�=��Ej��'�O7��ٯ��ey��+uq����pa�F�o}���'8�>�9�0r�1W�@��P8�O�����4��v�q�Q��v�Zp�"X�K�?.N��г�G-p����'������C���Oe�>L��:�쀎aa�:?�K���������D�cۜ���1�D�ga۳����7z��ڙ�_��LQ��f���v�ӣ�(O!v6�^4�@��("�ӱ`�)TF�6�0o&�_��f .��\L�0멩��!ڹ�FzAM~L��ؓ�P�)�~	���joeo1��^�b���j8�c�Eq���b3� R^v�8��žx�:���*�O�3���~<<��gVbP᷎Ɣ>;˺��W�3E!訾*����U������c|�����5cze��&4cqm�;�wU���]�0ʣK��,��n�k%�I,X�WNʐN�n(_v�»;���\���I�ݤ޶1�K��~�3��͒���Ü�zg�U^�MOP������V��� a՞zȴja�a��)3�HQڭq�~3�x��d;����g��_�3���΄�N ����m.��V�O����4�F�p���y��_t���3/K��m]u!��F�P�kNoa��&�� Zګ4�@�g�Eۥֽݼ��N�P�:�2��www�^ Ѕ�JH�!s�~��9�[��L�����Um�)�1�c%x��	Ώf��lauvʔ�^��H.�n6��p��wΥu�x��j��9i�q�$�EX"�g�I�#R~�B�~�P �H���<�k��vLj�/������=�{�]ssJ�+���OY�i��b�=%2�5t0�9n�BGq�ܽ�W(���L#W77:���漏a�;{ʙ��~��,�n��|D@��f���yg~���{X���:o�
^:�Y�����G��ׅ��6��G;3���e��w�3I�va�fKiV�"I��_0�? y���O9�}x�Z�����Ze�:;K�D��«��Ĺ1�~S�n�u�w�uX�T6N��y��z��o7�������L�Ė��*�N���+o��6�N3���լlռq������e:��������|$YD���+�܂���8[A��g:�L��_b�{�5����I��J��>�+���9��>�F��4�`�ǳ�͠^S,7�#�|��T-�a�`]5�q��Ρ���G���N�|�H)�B�Ct���n�N���bL���� �{�!Y�3Z�>��Ul*�����z���]����˱�f\߱��|��8uy��P�ETy�����Fu���m�5�����Hl�]�ܵ�+��r�{,���f�=�zT���Vm�+j�mf���Q����G�Mt)	��p̟\ө�W_Ut�����`���}*sջ_�@�o��Ҫ9L����~}ۜ�РED��^����F�uR!O7�E�d7r�m��WQ�]4�\��iiǇ��]3�ݻ�dç�e���7z���ci����{�kﵺw�j	�=,��w��CeU�Y9DӔ��1]r���XSt+����:޾-ʾӫv��!�2{j�ܩ<-\)M�tXJ�Β�V�#���
Y+�� ��7f�?E�6*�t��dK�Ս���;�x+��w.��@�s���¹-�ZΌ*��������w�x}���z�L��w1x�PL�s335�<U�=;�����VY�;��^�{),S��x�qí���2��O�9�0+P�͝��%��ІB��Gq>���v�[#�WH%����}�ؗ�,8"��]y_���wzc�joMiדܣ���8�����a�s��C�p�8��BL����;q�I/ʪ|㤗�8L{��v�
�ܮ�����_����5�>0�im��,Xp��dF�(���ҜP�aeeD(3���4��vf�,.xO�W��~Ĝv`�p�v�/�5ֹ���݊2ݽ�v#�����z���!�sH������u��+q�Og��̺F���6$녴�oX�dm1��p1 `��w�t����.[�͛���0�+3x5R�����7�.BS��{{��b�N��� �K�/�߲�J�j�Yo��� xG5�*7�n�t�J��j�����ŢF�t�`�S[�ӏ*����(��&��`��{K���է���8u����B5bgJ�.���x2W�Y��a����U�µ&Y����55�'y��P����12�Z���s�+��5]zt�/�z�wqY]:[����3j��P�έ�R�){��������=��ͦfd�BВ�F�Ѭ�dA�ȯz�x�1�gkjM�o��\���;iKs�r���}Ц����+���%����l���j���Yv�|y~�g����-	��x!��{ы�[���;O�z4^�s�ej	�t����7-�À$[�u�o����W�*#�i���8ᬵf��B`��2u����䥶�|�N�Y������e|�u���lc~�J����Wsڧ��ٯ����}p��(KT[]g6���q�D"��7o��[�ϯ�牐�?H�h��^��U3p��,�]��i���l ��kў�΀X�������w��Fmt���GŻ��8��8Ck��`�;���*z|`����}K�0��2^s�c�*��6�㭷øc\�[���9��흷��ҵ P�f�L��J��R�t.��jU�`Q�9��z�,�ӓB9KB�]^�5U�uɴ㯏��ymȞ���zkd�0v2�'>�l`[��������\f]K��6�K�{p�yݳ��i��3��B��h����bKu���cd7�3��_1B��;�O}y~ćdɕ'U���m]�5��4����9ֳ��O�д��eܚ��p�o-��%�⸴>(Cs��ھ�e��_aN�iwV4�m]��+d{��a	�UMg�T98+N�D3��{�f���˗[s��K��8��6��n+�[�ξ�B����O,B�.}nCL�]��HI��O,;�B��5f�ͮun���b>Hg"C��9jd,	�1��6�k.t��7�{)]Ø��a ]�t��I0II>��W����Q��\�S��c}��n���۠���`=�/;QY��3��Xa?^��y~]�=�e&G3~
�Y]v�\N����7��:����&�T�s���v��P��o��v�A����tc*�G���bBPQk&���h�i��d�⧝巌!c_���d����G��7��i�q�E� �45�D��zQ�o�G0q�]m<&z+��x�$:D�R�+Q��y_I���0�d�y٨A��%� �d��Bei�V
	3]�cW�&n�R0������  �Q�{��@���G1�{�i�E�&z���������{bdFX}�|1%��m�'d��ݫF�c'd�4��Y���ݫ��j�'2�d-�~��D�N��ÊL�}yW0w&/��U��v�Z{tl�b����q���z��F��ނ��SƵ��W�6WJd՜v.����қX�F�JR[��$9W� ��Q�'}O�O�1��t�PW<Z�}���-X7ś�KB��>�&��}a��� �q:�3�ygL�<���fi���F�����M�+N�ȱM�r��ޱM��8��Ղ�Cx�f��I�b^��������ŝl��8�M��ن��:M�2���]�PsP7Ydu�70�Z���F�f�y�0�	FȨ��p��u���٫���jW��XB'�Q��.�γy�9x&;���m�GGb�§�m���p��r�<�8�g)�`��ug�7*��۫��s�*h9Y�����6֒�n��%ݗ��|7��6�}�$Q_;�9�ް�oT.Y�l�ݳa.7���o.]��(ݮ��Z �ce���l߳kh^nV
��	۠ʐ,�1֯���)�u���f�3��uj�׳xo^�+q�n�\6�vC\��g�S�]
���rwI.M��ͥ(��Jt;��z����6���V�m�.H�%�H��4FG��8���q��q�^�}]�t鱸�^=(ا�K�m�5������*��Tj!��������q�x�ׯ_G�n�:m�5 �	�/���;[����j��j�z������q�x�ׯ_G�o��{�k���"MzsmxѾ�j�)��.j��RG�rs�_�]5O��ʽ5�k�r�Μ�ʍ���kv�J�6��m�F���-�ܵs�,\���6�����n��sK��W�s����η��-{W��,�wk��soKm�x�5�Wwgv�����׊�-sF�AF�c��؊��ޛҽM��]���?���4��7#�n�Ý���������)O��&�6رo^h�l��g+�lN�5,�Ǿ���������J!�7dESD4�����[�o}��4ǜg@q�J\K2mȌ�����]�>�-ȚӬbג��RF�R��;ƍ	�x�1^"�)��F�Z��/xl0��\ޮ������pI�N�l3���;{4eY:�u[[�T��A�W<ݞ`ǻ�v� �~HRT�傷|���qh��;�p�M{û3�s�s�n�z�>����
9yv��i�Xé��<Eq�z�܈����޼���8���wO�2���fE�+��3�̽D�A�{��䕅mwob����_�f��?y
~7c���3��"�N�����+���M�3�H�vb�O<�6�*i�������S7')�ܼ;�r�Zzލ��@wq��4���������� 9�2�s~�� �4s��D���S�����B���<��P��l����uh�S��)��U�C��䰞��>��$1؜��ݽW���T-�b���o�W�*\�t�Z��c�U%yoF�9��%@i��P�ؒ\*�`�IE}��:��{u�{�y��<g�f{�@�t6����u�����%:�C�Vxxxxy�OKwobR�U�� ���Y㯣�z���=ǧ�s��ݍΘ��e8����'��K\5���� F�ϬW(V����m���3�sb��]�������->�+�=����r6�L���z�Ja�0޾6ة���.%���H�ҏn�oq�*g�g�<�L8�3�l�"̶0�n����vd�l W.� ^p%1�ff�ev����`a-͉�Kn�M\˓�G���]=;��ui[��� �m�0���Vv��Vvt��Ν-���xvx��
p�j}\W5ǲ���Q�w�rt�x��934�&`��f��7 �d%��K0�#�,�W�����0�{�̟a������wl�:Nh��.)���z����.=�W*���Ug�Ãw���rzs[n�5��gVK6YJv �2�X/(W@wʽc5�?��Γ��*7Z4��C�y����n��U�}�J�۳ �ݮ�%�}�.,�4�Ѻ΀�~}������	Tp�?C�+B���n��dkD���T�a ]�]�@��lVV�j
i�R�'���b��\��>�Y����R������nb����ޢ����_e��>�*8�m[�Yz���=ùql��3_v�4���U�O�pA`�wWr֑�} ]5��Z�,�c����e�݃#��	�D�tp��>�}Hu�Ï��ҩ#���`��R(Y�I�˱��c4Ӝ�Ld�P�U�Yh��˔��n���M��ٻ�&�S�?���]~>�����􈥐ܧ�߃l��㯅�<�3E5����P�at����]���魿FP�x�vp�2�����׾M�ʞ�{lܾ��:���'Ӕ�e��Y�2����ޯ%�Ce�V���[!�pF�"�m��#Z5o6A�3�ڪ����3ǹ��5���rX�k�3��.�H���a�3=�(��x�0��:�Y�wE�g�{|��gO_��]���nO\��,�m Q�)�1�F�ƀj�=�۪
����ؖ�:�D5־���NB3��,fǜ7$�t)Ok��c��'�uݹ)AuD�Z���2�S0n�A�fR��U-�WF�Ú�y��5Wn�R��ez�(�=���N�L��K�}��7lU��2��9Y��Nw���hn���(�����í�As�9廜�{I���i#L8�V*T�,x������>t�f}u�B��1>`�>C���.;2�^�v�}��[Y��*�n.��kl"�zG }��z4����=8c�����e�xe��O\��D��vw>0��q&�e�pu�N���e�rֹ�"5��4�mi����{��g�K|���~/ �g_���i���ń|ޒD`$�L�ʕ6r�	������Kk�W3��\��@��/՞ P�.yᦢ������Wm�6��sx{�$��6$�t�b�`�5�vz/��z��gՈ ڕA%�+�����+P���jA��b^�o�!�"���W)��6hUgR�60�����#iel1����(Y�F|sS�S��SӸ��H8�{��u�x�]�i�+9�����*��ۙ�x��ݏH��\���w9�M쏷5���ϱH��s�$�oɽ�lk��)`6�T�f��S����m�UA��w�M�g���z���N��;�lB���3Uy���]��@}�W};�}��3PA���]�$�=��%6�Nw+Mwo>_fu��\p���e-]ZC�wx����/�*�ju[+n>C,��ٙ}��xxxW�xV9�IY0��gwgw��AyHΉ�&6ꙃ1Z���Pc�> ^��ɟ0�׮��f�8kW�ukNd����f�J7o��D-^��Mߧx����O>����ˣ+f��m��ם�L��>�l���sΎ�)@���������S]�6�j(�˝:Nw���l/�3b]�h2�b���_��L���rҥ���u���)-U�:���AnQ�}�:`8�a�{&+3�\�7�-�8�tޜ�Ng+�Ta:m$�2�ha�6��Uc��x�8�OΤ�gT�
끶U�2�ex���*��u������{��g�k#��A9"$�TVa��.�fw�t�H�B�G/��9mM�+Jt�X��&Ms`O�ZS��ET�����H��̧��F���㹹̮=K� ��g��{�T!�3����ϋ��������	8�v��ߛ,#O��uv�!���L�{��H�Y�K�s7�2�AM���g�k�ڛ��ی؞���d�H=.����/p>�#XbM�9�S쵅g!�{rܨ2�ȳ�
��ɠVs����+f7�7�$�{cm�m/>"�l��
���j(۪oV��,���U���ө,��d��^Q����%��:{ᙖKt�U�j�q������0�&���mz������Yq9v�o�Z��y�R0�|zN��Ir~�}��n�m�3��͸�\�v���w�s��"t�t�V]]��$��͛�P���Bj��+a�qu��T�ق2;z%�W���r�`��ޗ��0x
��{J�����-�<wN�6����dH���ԘS�����S-��ef����Sxf��;���3�1����k٘�k2�'x�F>-����:���Kq�*�(��JY��z��J�=���}��v��&S�ݫ������(�#w����:l�܌���0@쌵g�T�1�[FN���¥z}�q�2�lvμҀ���-��9L���od����_�a��7�ӸO*Th�i����~�%M�>������xx�ۧ]��z;e͕��}{ϡբ&L��±w�G��東�=]��b��K5�;*i��V���7ڽ����rN�<��R������z��oz�:*]~�O`U���1��{�jys�=��M����p�}˻�up�x_i`_��02�Zʷt�^�JH�<�z
+�־��|>�B9��,c�9$�AeKh�6�뛴�����'�`��<�ӝӂ��u�|��F�b����
X[AՉ�ȧX�C��
0��SB��W��wY7ײ�ĝ~)r�CV��e)ا9VG�t��A��v�z�ax�۵��F���"�T���ˇu�P�Z����]7oz^�v��3p�/��B�����#3�j�y�5���h���Y�.k���������&�l�� ���~�Pq@�F�;).Q�}=���ՕJdtq�p�O�=k`dg1�P��^���]��{��#M�z����NR��\��f�a�Y��yv*�Vn_�S�
۸
r:=9�"�q}ك�b��Y�3kTRѤd��bt�/2EP��]]���X(�b�u�ϸ{��)��џ�YU�k'o�l������a�j	��o�Z��W=֕Z3�ѳ.����ղ�7�tn�L�v����;���N�U\ �y����j���4i�'?,F=}���b7]��7�E�k{�̪�����Pf�Aϴ_���8j�;��#�0[�;��߾��ýY^�GMhZ��자Ko�&ƻ��k�%��t*K$�� ��W�>���(��ܼ�-w�;���v���������3���$ǜ�>f:w_L�=�+��P��*�����9ʡ��:���^��#��cn�u�jom1��+4��/CD��Y����J����>s;��0�<�9T3v@��v��vJ�����&H$��-ۯ�0�@C(�a��#!����a��ݗ�|��տi3N����7���=]Φ�@:�mfk��� ���� 1��y,��Ψ��=M�{��\�=�k�#C��TL���D������)��dM$�m
����&��f�Z[��)�$wf���ycPYPib�aG}��|W��D��=T��59� /V dR���㹖��UEh�&�ر�n���^B��hF�lC�k}�V������hAg����Wr;��6UK�(i�a� �B6�7����ӷu7��7+�i��n3vlˋ�L��3�*�_UN�VhZ�#x�8��M^U[�zk.-]���'
4���!�}���QC�����h�8V��bz���r�.ۀ�[ӱ�]��N���s�=�sKĵp�#=$��YN������(���/��e�R��ΜZz���lS���2�w[E�-�M����eq���Jr"�1�8�˺��Ot�*�m���u��B`8)�~&����5��3��v�`cх��3�R)�m���ޫ�@��k���9t��i蛸j��ڤh���Ì��fl�� �1
�Wv�%��M,r	��8&��U5���m��ᥘvO�z�ǡvF<l��=�+"�-�5�צ}�I]��6|e�H�<�w���u�]	0[t��ƅ���3�������[^a7�(�5����Anu��{J�Y�1����`�Cu�ܨ)<k���{T�	��bO�
�(1���s�%�<�`�fQ2vf�h�R����*�	�/��qq�K�#|����`�|�/zy�<^�E�/t�'��gU���Z��O�C۽�n0���30��r*���e����K|�k��a�;\��"��X��2���jg�-�c�u�w�����Zg��|��b�ܒ0��2��q�-���6\cu�3yަ�̍�&��a�;��gTUϳ�`�c����d�#�����CW4�a�.��&b�C$��}|΁�-5w<L�]����1A�c��N�-7%	��p݅�9�e���	�/�{�N��2_�T0�ȃ�l�F��'zx�3Ƃ�R-^|۞ܠ�Ϲ`�U�����f32vv����T���V��f��|�y㍭��TөVzO9��g�:ߺue:>>��5Fs/-B��c�ˢ$�x6o�4�oGu${�8����I$]��M�SR/���窻��8N� �0�9�@Y��t�@��;eJIv!Uq�nSk�-�>/5��g�:�}
���A���ҰmD�ރwx��k��-�>ئ�0��%��v��m�Y\� D��|����f1��3��V�8V���p-�]��6Z�o��f���QJ���E�hV��1m>��eI6.��ֹ�Js����1Lu��E�!�7^Փ�,��h��B���Ե����=��c�@���D�v����j��#��7;��ú)�)���}�\T��b�ٰ�qI76��*���f���q��v��1Z޼(;|�\���Q�&n�%���$e<�{ҹ3�V+�Q��"�G[�1$	ӎ^�Ź}�C�Ev3Yl/_]j�v��3at_]�q%#O�X5�O9� 4���L�r���ɸf�:�=�<[t�pf��,+μ�����֐�s��E��\�7d�,��YC\��oZe���h+����`7�ewa�|llʚ�2�7s�Y�+��Tyf_^)���b���jBk�9R�����X53i����}�=}����WT���C�ag��
*��^Zl��є�neAzgV$k8QE�9�}gJ�2Su��w�� 㫃�{�[��n;����#��]8�ˍ��^RMUN�w�jO%��z�L���#A��*���6Ļb�wn
˻XE���.��{�Q��O�v�fڤs���[��ŏ����)�<+�:6�N�]���V��;ꇺ�i���d�m�r�V�	.������qT�jUR�����ʤ����C	E#�.�� �J�a�(lۏ�*5L�.���x��Jg�������&�|H�מa�tYv�12��m��4�C�o��:����&��']����__oZ:�����[K�d�M8�_^���崮A�W���t�Ҩ�t����n�C+� ,��{��f�i�*�y�P�Wuׂ�5ïYQo۲v��R�۬�G	�����xm�j�,dJ�kvNoFL�v��j�bD)'W\	�.�6��}Iq�Q!���Q(>D�h*[e�Q�0����[�a��fã{���2S�w+�ɼ�:j,.]��}6���˨���է4��H���#F0a�,�T�1������T�3�a�◛�f�,�\�����.��٢p��ufP޼{̈́�V���sl<�`Fg��j�u�.�E8U����5�N�$�B��ޚ0i#�Ǟ��b
�,YhZ峗ol9f��[���G)eҹlm�޲��V1�����dt�=�Y�X�5u��d�@�n�J�4R�+�7�4cL����Jq�YQ�D�0n�7��;m�n�u�yQQ�YYZ`ʵz�V񬕔��K.���7a�:(���C����Kv���՚e��W_3;UN�]՚OB�����AǯFm�B.`�ˋ:^�T�.���%�����m��e�7v�}ռt;�-bɋ��J[�ʉ�ݣ7�����r��v�R���o�Uj�ms~���cQn�����!! HhIQI�����㏮8�z���]�t黂y��V#_Kƃo]�0HH�b�0j�V~�}x����8�<q�ׯ��v�ӧ�	�HH��;�X���W7\��\�	C���o��oq�q�^�}}c�N�6j	!<���s�Ȗ�6�75��}��=-�-\�آ��v�b�����sE�A���W�e����6�i-��PPD[^ۖ�4Z
����Q��m���[=v��\�1��cF�h1����DT��]++���[r*g����\�&$ɽ�+���ll�أZ-E~J��7���a�4I���M�Qi�I
J@e�*�d�l2M�b"���B)U8�L��e���ˇ���ո�U���L���.i���W��jtc�w�F=VUQ�͒�
��wt��a8����2�DQ�0D������b��h�P�	�H$�-���A"Q(R���l��	I&Bl�J�`��"$Б�P�JC!���q"��' a�0�EdEQ�(�(h���C�1�wz�|�o�L���w3��A@�li�T�}4ȸu�ۺ}�ӻ�"���$��v��a5���z� 3Ϩ��WH��ɏ(���CZ�������a��=��p�uzLJIF;�J[��PV�6]۴�72Y�w]Bbe^d���y��da�(C��� ]��7DDVOf�c��@�c��7fMQKh�ąTz}.)L��g�[s��cJ�XVK�Ӕ�;mqe#*�ov�����wgvyP�g����mLo]&��g-,c4��0mݲ0v(ݩ:�$�+�e|�C���g�V"��]��n��%�p��z{���Fٱ�Il$q�=�/���8;�(Õ�@E/e9���!�+���Z��o	�xf���u]�ɴVWO�)ԁ��`��Β��}��ݫ�7��Lۮ��?��\{`��n!Ԧ���6��}7����t��+�c763�X:8{E���̛�oU����P�.I��G2:Z$�N����sgi�&c�v����[q���9��h��8�<�4g�o���+�-Gr��wȒQ�M�r:Z���R�,�E�w�pF����'�2yu{��a2��&k�$�Ӕ�{f���5K�����1�b���9����{ͷ{�a=�4��Bz�����;)P\��v"zC
�w�w���c'`ff�[��>�-�?8
���f��w#c��%j�Y{���jrY�4zkI����[��9o���+����o�}Z爋����um��9f�"�Ͳ�#ƒ�!�=���� :��ۣ��ƺ�8�"`��
�]
�=ͻ}�C�@����a�6

gD����g����F�`�#ʹ3�ѱ;}3[���EwGq$qǏ)�<��jh�2�)��8�iwP�\`W�䡝�sע�&�B^�Y��~���
{9.�-M7�*�{:�>x(+g��ΠF�p�H����cV��;^C67o7e��sP��׏���\�5�������C��q���XT�g�"n)��F�kJ���[ $aj�!�d3�,��;�K?8�������ƃU��鎾ˡ�/i��R�
oT��$��fq��`���9)�fݾ�=��g;Y�Uj�AULz4����A�uu��,{2�b�]7���w�_�lU��e.:0�&�!�'��l)Z�<�c�Nr��O
���T�����w������;����N�.�HH9�&v���a/���S��ߚ��gOi���y��V�������<���E�ǲ���uN^�M�tVꡣ`<�|�)�f���#��ք��1����N4ef��3p�{[����`��U&�\yn7���X���oR�z'롔m�����7i��OC�8�3�h���Z�^��d�νH-�V��6�P|Zo������G��9����g��>��a����m]�f��@X��|��M��;�r�t�S���?���\�p����w�tN�]$��I���jG���J�Hl����]�k1:��r��kNA|w��>����g�l��ޯj�*�ot����6�/]��M�E�w��ȫ��������f��k��~�~LP�"��;t��Y`�F��hXRa{���5v����Q��{�h:���j{:�P�B�ݝ9:�]l>�]h�KO�������;�rJڍv�5ۙ _U�Wo��]�.��;/�7��
ł�VD�S��-���|2�z��>�Ȧ�\J��ۑڋ��g�l�����ӑ�L��#@Fj�Oѫ7SN�A�גN�r���W�{*��ɦ�a![0��0\dAΚ�lp����.N�a9Ka$��x��]ߺ�����x���t0�{��ʋr����ɔÍ����O>5��6A݀q)
�(��)��ȋFt���e��d(��o��8��NRJ�2��6yjO�U���ԷZ���-�U��R�C90�ԟ���`ǻ��'��ǰ�잭̚ݍ���V��3B���|����}^����f]�xs1-/1���#x�N�8�͉��k�Xb��#e���ݯVy�\�*����{L��7�1�{Vj�zGO]$��]-��S���9m�Қ9sm-Rb�s��|��d^�5�+���G/,}���u"�|�/��a�y��.ƬZ5���勁�c�zo�b��&*��^�o���S�a��CUYwO��ݶ�p�}b���va<NZ��#q�qb�l�S�2ҌL��;�2U����$���:�>�I�^�Zޜ��;\��50�{*���1I�٬���v}�}y��󼓹�]2�i�s:��:�tevNQ�^�l<_=2��c�M3�8�Jꂪ�]vCb|v;���u�t{�Û���u�Ӥ�z����Kj�hGy�n�LDN��t�V�Wl�'0��MMiݲS-�+.p�����=�\ �k��q�E{vOw@�x\�2=���ĝ���2��,�&���h�Gv!��#i���t���aqj���
���Ռ�����,P��T����L�;ʠ���}�NFת���j�êf�-,آ�!�A�¨�Nz�D��>W�KG���0�٭u�199��&�a}�,��������k
�)�:Q���e��a$շQ�Gd��`��y�q�3���7:��T����5[�l3�}ؒU���"��hŶd;����>�r�/��s3�o��g�e[vSt1W'{5���+�q�.���vy
|p$^;$�/�1�A�53���LMC#�lU�x́���v�W�C7�XJ`洋W��3�����E�.�ݦz^�q�C9Di�5��/uD��F����!y'L�F�Sۘ3��r��S�c�o,mi*�N�s�Yg`�v���7��y�<��d��(�Oܖ��5>�/�c&�uڸw��������=p.��D�{�u�Mj�����8������Qh����X�U������r��g�$6 �GhGB���.�$V��H���#6�E�wKbl���%�V����v�w[���-����v)��Ww����1��~�*�'��4�o��[4�@�>rň�#�sg=X�4���S����;/yQ��Gw1zL�{s(O[�ճ�@]>t��Vh�Xd9��17w���ӎZ�(%.�#���>�t���G�}�.GNQ�ω�����x&x��;Fsz\x�, �Z���Wu��*�eHH�Jրُ�8ub7��
��Wz�t4�� ��w`VqQ@���ۢ�[$��K(k��3�*޴��^�rD.��}6v��M��$����=�W[E�DJ{�y��҆=�dKq"�bU[�Oj,�ʨ�"��ն@2��ϩa���j����[
Ó���S����U۷��8�wKz���wp�d�c����WϤ	Ty;Y�7r���6���ܙ�P4ohnn�c�H�핼B���*��������?�Cl0���G����žԢ3�썍5@����n��1�˓y���:Or�̖��� p��̹>�Ҟ��Zi]Qג��{-����۞I��O��}�v�d6�o��X�'n��v)����VLҗ$%���x�3;�l�aj�!��π����-����aRS*��=���I�T�q��}_�{�.���ט��JC}:*vX�Ž��a����/#���bg*�v�zi,�{��׷�\rp���A]5l���oƍ���/.7�����y�w�QW3Tm-�N�K�A�,:ח~��b"�ǰ���Yv�ocﲏz�4K��LTI�������h� �Ewk��������ܗMS��B�@�֟"}�.iԍ�p��S���V�p��S̓��n�^k@���R2��s$�<	�pG�\o'��yl�ϼ눻:�F'|{[��wM�S���`^��w���1t�Cx���f�4�sYp�6I�W�b[�F\x�Ļ��_j�\���+cζg:�w�9����ohO�g�����%Ω�����]���<Vw�T����>|��9�����ɧ�$}��s����Ɵn�r:�2o��l�s�����g�
U���PD�3#��mK;�4OO���6��l"���'X�K<3�z��;���>��'"{Tv�{��J��&U��k���zڋ�Їt�c�
]�4r�Vp�y�e��2ԩm�K�V�&V�����}�a��Ј]"�<��Hf��z����H�D���OM�L��|�[y�!>͖�%%�!����&���6"�L���0���㽵≮�/����&����[�4�es����OŅS	,��-��Bs���6�xxJ�?�l1�ԧʃ&Ζ󴧐=���}�`P-Cy�R�2�o���2��Y!*��Y}�m7�6�Ժ����p8s�Zh�W��X1�����ڂ[X��l�VN�cW���"&�)Y{���\4�T��%Z�[w׶�vM�?mE��a�Da�(r�"	���WU�P;�epl˔2\��W3�L�jT����S��[x2��9�P��ʎ,�u.̑��ȕ0ٮJ�'�������T��w��w֤���,f(]��n���|�:�h�=�;և��P�_�֙�Q�j
�u,��s�ê����_^�%����u�q�;����y}&)�D;�&�wH|ɥ�.v��Lv�69fw�w���;W{�O�Ҕ�5�,4�}��w�5٢`T
�c�o��!{5?F����m���
�}H)�L��n8����	��^�S���p$<�DO_Mˣ��W����~�H�u�{��swlk���1��qx[M�&��u��Ɏ�"�LgO%~at��1m�!�6Ԡ�Nx���OÏ��H�����rC? C�Ȁ�RX⦦����6c���2Q9���+��c=#�k�@�Y1�4��b;fn���|���(m�79���kN���҉�X�R���_��.6�)��2�":�7/��	�6ba�6waQ���^tJK�ע������ӽ�`B�y���ЮԻ��k����t]|-~�@�f��ݘu���j��:��e���գ��"�xu�c�6���2�!n�k�-w
��QH;�k�lҳ����X��xN��1u��gGV�$����y�N�\C����`���`�MVaën�����a�D.��I#�B䞛�&"��n5�U�"���[��«�/��مxks��!��qJL�c�[s���ʘ����\��R�ٸ}xL��wwDU�dw�H�q~�m@��t�|�:;T&wU��픁'���[2@$�&C`�g^�P�֫�}�wF�6�lg�Pi`H����qK���7��Y���8;�Gs��fC�(f��%jV���+�*��wZ�Y����W#��k����ٞg�����I�w����Y��S���F�2��rz��}�>OVψ�*��o��Nw��Iq���P���Z�(l��,v`ܬ=����5{�uZ<:@�|���C۹-�@��z�y;kq����Y�2i��Ъk��#��w�AΝ�wO]ж��hźsw׏ڌ�K|}E-�]o�*��8�ʪ9@��!������m���E�j��,���fՕop��f��D1c�=p�L{&��rl]JbX%��][���9��f���mv��DGm��)���u�(�R�O5$��o;;���R�2�oW
�W7�ŃUt(5}��V�]�,�Ծ�9(MCe�|6,W��v$�<{���=��I� ��i0�c=t�V�z��z�����G�^���Y�^�}�+n�(󺕗�@�e�jv��%N���q�8 ��/��g:�h��LR���w�Rw�^_Z� �Y;�B�����n��]�1Q�\���@��-;g�h����l�U���6�FkK�R��<�Q�g7P���b:�b˰�b��Ӡ22���ζ{c��k�:Mpc`�x-�(@:���v�K�X��1R�Ks���^$���ݫ�kX�9F���=�<��[�����xF]iү1k�qn���M|)��G�\���\�9V4��
�Ct��}�x.j	��`��ܾ�%ǌ�[u�u�cbƖ�m�ޱ�`	֯.����ֹ��Ya��yo��˦vn<M��][��鹉�qr���m�^���0��"֛�Du�&�P\�F�k���j�:�u��WQ��e9�X��c���6<9�uP��6�f�����f��c���[حꕜ�s��	B����C���5�U�|�1u@r����U��t�D�|�0�(�1R��h�v�u��d����r6��W�Α}��}�>�ұ��ڲ�[�wY+��.�g>{ij(�Wuv`��G:0)��vN���
�Y'b�]t�љY�!`G��وX���,��7�e��soOw�VU�q	�c�2V'���z���YS�Q��%��_h��8�:�kS�V膛��,ٰ��N��\{t]R}&�98G���-�Ɣ{ǿdǻ�Y�b�t�3�svݱ��r�;ܨMg]��r���f.��Ֆ	�+�"�$D�ȷwqHLu���:���y�ͥsU�{H�ث�_s�i�V�S1����ӧ,fjv����h�ã�'1�n������y�HM%�ِհ�'yb���M��e�>�Pν;̓�����}B��7z��\5�l��f���.�R��y���x�T'Y;�[��!0�m�N�ڻHUl�i��[v���,l�����,�U��^�XE�+:X�}��{��)4��F��]�!�"�kqR�{7�Ƞy)��r�+�h-���̡�(�ȋ&tk鋻\%*�[�k�,���#]�=գ������t���m��PX�������pkn��h��=����o�ٲl��%�h���^���st]�{�9FIA��	�I؝�d
��FA-��n;�z�8�^�z�}c�N�:��F@��κ
��)/[���}6��H�__<t;x�8�=z������{����m퍟}s�c5HD����C���^;��8�=z���릝:t��� 3���n◾��7�F�r�Q���U�b�/}pɢ�4X�ׂ�k��X��J�-3��&ƫ��/NXۛ_�v5��.����~�J�(�J�TVM�ܵ�k�y�D�(�\����^~n׌hz�X���_m�E��*��^��5�r��k����i҈�\��[�����r�^5��0�.��̪{b��/o�f��~r���k���s�f͡�L�{A���b��,�u�nB�t��wN�roX����xxxU
�����p������?0Ux�����m�7OѪ�,����n��ʬ�ڻ�Zs�Ȉ�=zI���!�.;q�^K�vͱ>9���f���牨��D�����"QN�375�Ѫx��ؾ�� ��"h˃o�i=�D��h>+�Y��`��^�}���5��>����q7%��f4�˻�l�=%�O���6I~��M���{Z����}�F]l�;��W�Lc�s+f�]�[�r��g�0�4�p�>�z�Wf��k}��F*�������.&�G�]H�����qc��:�_M���|/�`���l����0[!#Z��e�!�`-̟e��͉�bÕ�k;�v�Ɔ������үQ�SE����o���&Vk�vkr�-�:7�(vX: _3�1]t��j,���ԯ�! ��y�����ޭ�UZ��_jѧm7A&��,�����gY�Ӳ�W3+���r��4���ͮ�!6](L�1�R�:W��}Wy����ck3�X����u�x���gHyc2�7{�voF��ӝ�V��I��$bF .c^���UFw�-��^
Mk�ݱm�>�]����8*ڂ)@�Mʦ���b'j�Ղ+)H޷Re��z�ot ��u*���-��1����^�7/�s��)���y�6� o�RKY+�%��nub;�eV�ుY�	�34�v�96�k<���t:��UG�O���4�5[r�b�=���3��Y��h3G���N�dy���q%�{����I5Te��q�M�e^W0�����enC-0`����� Q|��6R�1�ĻF(}��^K�$F&�ŝ�0k�w��� �uǟ��P9ucvOP�<Q��&X����&��iӧ{qb�M�%�	�8'Gk�أ
F�#����l��~����a�pI�f�b��+���B>�{=Pa��nC�l�u^�͖��z���Jšւq�Ԫ�(�voD�nϕ��K׆�����*��G���O;����F�g�n���,�w_]�Jھ�ns�Q#.�+��SK1��	5n�^j���LF�I.�$Q���H���!�@{��_gv�8u\
�@���]��jU��-�g2G�5W�B�h�D�yJ�����f�����z6����y����KS�r�~�F���<�o��K�Y���ގe�������vp�R.�����\�����m&��S��������Y� ������X;�U@{�k��C+�H��=4������6-)��%�{u�N?IÃ�P��;��4_��:�ǽ��uE
qu��5��ϐ�/|���T�'��,�����Ǝ|	C�R��R,^�5�7"k5���a�t���9.��w������L���aC�µ�A��a��o��婄Dh��6�^�-����:/"an�1��m���w�,q�GEv��ɬ�~��{gLR��/�[չ�8����qy�ns�L��/9w�2n]_E�4�؝n}�]�8�#���W���mmVv��,�A,��/2eYs���U�;GTm��tc��=]����1�]Ǻ��Dp�S~� �3�YJY���Acz�}��uV�\qܭ����%ܑ~Yw]Wu-_��"o/]bwi�F��������]rF�F�$�e��ʬ�7s�
�td�<�`�R��´w[5�3�Ӯn�wDW��{d>��}t�G>d����C�Z�����"�#��^�c}*���u�gu/~]�3.�y�L����`FU��6ĭ1:Lg�I.�ۃt�>�0�}��=�ii��Jb��Si��1J=~]˫�f}�;������z'�߅;�ݙ����3��ٷT����,x	& �\�z����>FN{g��V�D>.��q�,e�Aܙ��;�3���(vR�	g��_B����⒨��m�4�6����O�f#:b:20�'�B�z+�]��Pc�����o�yWg�q�L8\v4�,ʓ���8ٶz��IF�j��fgv~������Cdf����96�|�fg��#cB���u�E��^�I��O�#��%���7R|^����]N����t���a���S�� 1�'tV}Ԡ❢��Y俢�vT��Q��7Aՙ9�\f'�ot�&�W���8���#Qh9K^\��b�z�y�r�Mn��a���iJth�WKZ����4�41n['�<T70����&�[���	��]gI�*�)���D�{�D�@�9o��j�r������&��/c�*��r�=Pl%�3���n�4��Iu}����L��[�;�6h�t��o7��ùR��X�2w�t��KkG�����f㚦/�+)�c�[%���ɖ(e���{��oD�a��RCK��������48/H�F�m�9V�Y{Ľ����:c� ã���u��M��G2�����|:oA�D��<�c۹��}�zE[?��^���\r��MWS
`�=o��Ǩ-S�My��+����>]�}�o�(��
Ox*�_��]�/:�&itF��{�Ym��CWl��=$ٯP{�������=���.����ƄHاS�~�'����s�8��i�߱��캵$����`�@>��������Mok�wR����k�Rܼ�~��1N�@�y�jz��,�������bL-�m駪}W"s���\X��d��I#qJ�VX�g�0B��>���G��W^���_CEX6P^JYк���[��_R J�j���n���&{M��kۥ]Po{��S~�k��S�aw�t�w�\O�̌3m�>Bt�� �7�k̾|.�u����X�d��=��hn�4�c{�R�;�0�U�Ϡ��1C��7�W����澜��IZ��&�)�YY~���v�#�9g˛�x���Y-�xev�XA}�R��F(2e��:�2�k"Q�ݛ�-��iM!@}�3{{A�ǟ@.�JeHa7�>�Uy#�R�ҥ��%��k�V]ܨ�z����t�<�*���|�H=�y�6y�3Y�[i���#f�z�ط5��(��hv�*(Uu��]���oyµ>���i���IYJF���P7ù���8�A�쨼�K^������~��Փ[�M�H� ����p��,_�s_<���]Or��(�R��`P���U��r��;^�S0aܮ��i曚�O�n�����Rn����a'�Y�D�Ou�.�IP����2����LO2��+Y�����{�`�_��V���H�E�dJa�j]�g���EC����tA����U�?-�Z�*���ҾU�-�a�n^]I�.�2��k�Ώ���Z_
���Q;&v���Kq�y�4ko�[�F��K᝛�_u�te�=���e���(j9*<��G�F��^p�����wj�n����e����ۅ�|�>�"�e�z��p�j4�,]�-��Ű^���l%�����`��pch\�h��=�����v�y�;5z�q�;N�Gc�x�H����n?njb0r;p����o>ۉ����ݽķ����m��mv��۝o�*K�Z�+�b��1*
W~�+F�p�FoA�n��}��}Ct��c��5��8�0d_OY�%�%��b�
71ܦ��p��Aq5���d���s\��cPq���*��>X:�m���1y.�e^���7��S�x�;���.B^��S��m�!�x��|��P��4*�� �sߦF?(���iu��K��ӕ�z�G�h�z�5ۂ���'��GR{�B����̺��������vAlI��|}��)����<'�
^/N�bn瑢��ǽTKC�㻻vEݓp��w��&}��'��� �86��b:��{ܶ/��?O\4���2�ݽ�(H�Q*�ڷ}����9�7Kh�i��r�sg[v_ZS���3�{��p>�}���aUk
[×�ڼ�(������nRʝa��ǭ.�yz�����H`7J��0��/P��k��uF&3�U�^�5�ŝ&��)k�fs�ی��6�ٹt�g�Vʊ�b!`�~��I�v���Uܯ������t��2}�ιm���x��쒵}3�AƄ�뫐���鬝�XUo=�s3����24��e�N�-����mU���&����G�,���"Qo3�����|�p��8r=��Pn�R�$�����~�k
����	:��j��F7�Ub�ӭ�g7)�7d��ܸ�۲M�dϴ�p쮀Ǩ�DV�㫭�rg`���DE��#���ĥ�:�Uƈ\s�j0|ņ�㝜���8����';�c·C�R ����<\|�,�]�Q�������H���?]��#~��?�g��� Q=Ҹ����9V#Mgi�j����Ж"[��\�t�p�4������|�̳*|c���-�ljtl������vWQ��0�\T��3S�]c��h��v"���\=J�S���zHģ���X��� ��5">>H~�g��T��3e?z^.\v������f�G7i��ʆ�J`s����Z��v�<9]��79<��ۙ��z��\ʥ�vHS���W�/���ŰTk�C��5�5� ������b�֤�˺�&c>]��}�=�Ͱ���{�A�2q����[�]c�� ���/��)#of5KdX��������*�plJ��>ð1d&��Y}��{xS#bPB�?/3�J��K׷��@�X�sO�N��=�m*t�ԥf�K�k��(�9ڀ��F�L��JEa
OWr/�&���tk�fl�2e��1��>z��E��{;�U���j*�U���u���v��[�6���o���o��P!��!7\�qծ����^�5(5��^�zW)��N�Vy{A}x�^~R�(����*6U�:�����׸G�I�2��x�����z���֘�ʽr)�ة��mZ�W�l:
'8ٿ��CW$�ޮ�U�7���}�㱏
�tg��+�1(�F�׬O�5?y��Y��4�����Y]�%�Т'�j0�X�e�������)�\��o���!XuE�&M�����q"ld���H�&
�OpP��rHw��¸�h�,���xU  x6�����(�_M���� [��K�SǬ�\�ra��o��!y��N�/��h�j~�G�s]��otϫ{]ڣ��D&�Z��N\��^������3�ޖ���x���a��S�n�B>#5�]��3q�܈��)���	a�j�[w�Ά���<a��W�?6m��*�ic����zt�m��N���m6ϳ�<C˹�7��\U2��>n�*�_%"��F���V�1��Hu����h8�rܰ���
<�����N)���k�˧,�C��Z�[�7h�9��c��}@*e��yC�`��t���B���0�=1GFt�V���w����V�B�ө��G
P�LM7�EQ���p*o.��nnǸ�3�ⰉDM¬�v���%���@|?w�_��5�����@Z�J���������(���� ��=��E�QѺ�Z�)e�����Tԭ��ͭ55l���b��Ե�R��,�Lc5����1��jV�R֚���֦��LYmMKm,f�*�UfK5SU�,�MM�5-�R�5-R�m���M�ڥ��T�ڦ��5-��j��ښ�������6�Z��5��*�Sj���ԵMMT��SR�5+Sk-SSj��i�j��T�֦��5-SSZ��l��jjV���55��Z����ڦ��5+SRڛYmMM�5-SSV����֦��55���MMjmejj[SSZ���Զ���jV���56�����Z���5*�SZ��ZjZ�SmMQ�E!�c�)����V��TԫMMjjZ���56��ڦ�kS* ���	B@�)"�!@ � �DE@! *�
 �P@m�BjkUKR֪Z�j��� A" �]�������Z��RԵ����U-JکjZ�K�!@ �Q �D(Tjm����j�X���Z��R�e�T�5�R�0DD�B��l�Z�d�kK�jZ��Z���6Բfښ���զ��wm\�����f��56��fkic6�Ե����
D"�wbF(�Mm1�*�R�������bͫ,f՚��c&Zۺ��ڳ&L��2��2�Lfٕ���٩���*ٌem1e������r��U@$QR0 �O��W��~?9�?�>�j?���Z��?������������������}��E I�O���G���"(��H(�*���D h�t�q�?�?3�!�Q@_�~�?`{��촋_�Ԝ����N�~_�? ��?�}��*0��"�B"Dm��l֦ԵKR�6Z���J�ڙZ�ij�m��j��j+R�j��Kf�KT�֦UM����f�fkR��R�e+T�T�j�j5QmFڤ�mkmV�*�Q�U&�Z��"�	�	j��T��QkU&�T��Rmj�U��֪�����MZf�5-jm6�Mjf�)mK5�SZ�kSY�M��ԫM�����5iR�5�ZZmSij�J���M��*���Z�SZ��֛Yj�f�5��,�J�V�R�+MZZʴ�Z�ҭ5KZ���JN�����g��䪈�(����)  $���_�������@�� �����J����ͣ��o�i�D�H~ ��h�=M�� p>�?R~��:y�ӰA U�� *��?�;��Eu��7�\O�����_�l|�����������>��`x������O���y�
�
��b}�P������~���O;�����"���U w�C�����PW������4'�_M2Y��(:��A����=΁�;ЉϻB���r<?BR� ����8����ŠDQ�N�hE����ϭ?��!����PVI��w���A=�V` ��������>}>�ŕ��JU%$T��[e�AZ�V�T��!k-+DUSlZ�!T^�%R]�RR�� d력$��R��ڔwn����������wnѳM2��e��a�)Z��[X�ҵ�iT*5���6gmѓ6�����l[m�mU6�i�i&QV�6���cZ��WCve&���w9�-mDQ�%/l�*k[��j���)Qm�kV�մ�h٤��m�&�i]��m���e�mY��Y+Z�%�����6�ZJ���\�֚՘F��嫻��)�w�  ��^��ڮʮܼy�ܗW�=z��^�ԥ�ݬ������n0��m�ۼ٦������v�-Uj�^7��7��N�{+ǽe{Ws�큻�wm�U#��w��˶v��.w���ʶ�d��3:ݖ�鋏�  ���}j�J�!$*Q/<�Ҫ��i�liT�����T
�a��Mi4����y�.����/�V�v��g�I<^��u���U��Z;Ý�{:�۶�:��z��J�f]��[m����l�^���b�m+��I:�f�i�   ���իn�j�9���F�6�n���U��7�ww�oM�ڥ�Ξ�K��m�l;�v��Ԯ�;��<vҕ͗z�kzm���J�w�mx�f��ݯs�w�m�8��m-�n����SRQ3Lʭ��   ���U�֊�Ի��P�vy[޴լݽֻ�tw7{j��z�P�����z�]�ݞ���֪���u��\�X���z��Wwu�p�����^٩mYZ�M���kX�A1>   Y�=��kf��'��S7{���+֞�����P��Y.��Y��j�<z��W=�����T�����Y&�p����Mz�{)�j�UOuW��&��ҥa��l�jɔ�  '>��n��ȯn�otx���Z�4ޤް�����z�UW�ۭ��u=�u���m�u�0�t�K�՗��T��]y���j�oJz[m�VE(��3mk#R�|  Y�PQO}���+�X���( u,*�@U�z{� %E�c��P��8�]纽�(P���` ���@ ;ʼ�mm�km[�slUJ�(�� �z�t�S��{Ҕ
 ���xJ� ��ǝ Zz���A����BU���/gRT*���@�X��AE=�� oaT��J^�R��V��T�k�ݚm�� ޽�:k>�k{�  �=��%sޗ=�I�:J(
{^�{�RE	���T){��<�h ��w�zP�F��k��Pp;���w$퍭)ݜ����]� �z��)�=�m�ҕ��gx� ���xw�hi@��8u*U4���� ��=��@
9n�Rj<��P$���8 {�S�	�T�@4@��a%%P��S�6U*(   �~%*(  S�	T��� �Iꔈ�@���~��G�'�Q����Ͷn�jƌe��y8�r#mTF��\}V��)+�P#���������������km�m���_�m��kkZ����kl�j��׿����J��?�����8���%SYL��A2�F����C�b$q�u�w�)t ����rbj	��s��1�MS#"�]�y�6���~�`㬕Zu���,*:r kD�ؖsBŤ;�/r�5�j���V� [.�V˗�@L��F`&�Z7л���z?a��g%s�F�0��.#+#�,��3T��9�ƚN��dy`SzJ��ĲT�u�Wt-;!�Ï>J�^���"��'��h�z�m 6��K���ڧ�!q](��]������	2i���T^���I���ZƌQ.Ý0�rg�70�cZ�4Z�I�Kߜ��������=x�.m��<*��Q�2<�Ţa�}�'�`�=��LN�f�\��6�{I���i�z���dX�X�lR�t56aLF�����=�L�5�6Sz��a��ҕ�h�3n��c��M�8c�":�Rgr:�tÃl�ȗtɆ�&�Q�Ze 6�m�&���]�<�q�s&X�=X�2�H�l�\�oư;�j�C)�^`��!!,��$��m�n������w,@����g���goh�͸�"si�Zy�J�٠�n���w�I��&M��[��`0��F���U5F�#2�n^��՛Y�,��`�1:7��z�^�)^V�l���6��Kx�@�Z��Dl��C���m-�t�)����#z������F��nS;��v�)�9b� ĉ��*ĪΙN�ٯ�ʛ��l�C_��-����Yy)m�i�KpKܫ_d�	�^0sˌQ1�ʈ�C�O+/\��R�p+ffgU�d����(l2K�vdH���b��a4�s��J�v�R�{,�]Ƭ]d�br,�N�Q��t�lv�&U2�-�ɺ�ttM�I�f��a2�()V�Wx�r��l*U��r�M�%2;m�$�rc�B�'���
h���J1��.n��w�c-m8fа����	h��v]s~ۤ6��N;��u(,���T�"����!LHV��MT�qo��2Kz�C��Vi�Fā`�zI�,�����i;R�&V���I��[b���+E �v^�cN�� aHcEе����Ϳ����2L�3)�$�z��0�����TUk@Z�E��!�Utm��3�ItChԍ֨۩�mb3 :�a���&�em7aI�X-���V���h6��*#m�ec�B�!����� UHt82W��j7.�r��VM�µ�qp:kxLzt�4��FXK�Y�n�5z4Ħ�Ě�e]ap:������F�է��6�7��骶k.�
5��w.`;jn�F))p(-����4oo�cf� ��v]h�+Dy�T�c�bf%{X���Zi"*��GlJos��x��0Ǩ����D��1d�03�t]��󴶞���W(�����ljq��`�^+��6�U����66$��f0Q�Z%٣�6EK2�"��ca
�E���P�ҕ�"m�WWv��=�8�5uF1m ��-nY��s7h�OG6 ����<����n5.�:�ֈ���Yr�+'AJ��b��U���kvƝ���Ŋ�@��R_lNm6��[�ɃyT�[�X�S*͔��Br��ro�����s{��2Z�"b���2٫XƸ��ViŹ0�ś�]#,��8�僷���&�@J�K��@M,�T��2�|!mǻ:f@�z���*ܭ��+�h�Y�am �m޲��������T���-�b��)Y�5���YF�$�F�p�������!Lj���H��ź�̂��z�7�.�ӵ�
ؓ�2�"�݉+�+5bc��)vКû{��hJj�V]Ek�o�RV]���# �xlKN�������ݲ��B-�3e(ֆ�f!��Z5m��{4\���R��tk>;Yn��
�\�4��n��^�ەnvi�ⶆ��(�73$�b��ތ�� ��^j�E��s5�E^�4� ���;�Z�n�� �c�Vj؊X��b�I�"*�Z��*�'����&-R`��!	*֚f�J�"ɹ�Ý�	�J]��,!�y�9�:9�4oRʖ�M�����V��h�wؗJ1>��CmM#cQ��T�s��W��B�xs"�ǹl�����N$F�+Aa��-����ڪ醪JOk@;��ֵEa,�а��-��C�.9r���kP�3Zn�7J�bp^b�oIc�YR�w��Ij�QG/mdz,�ML	Z�̊����/PB�f����	S/��&��3%�Ɖ��н�j	!���-5n��"l圵Z �4=�g���r����0mJs�Iu��{%Dv��!�� ˦��lx�¶wVq�Ù5ћ/
�G�5��PU�t�uAr�n������04��;��/���&��(mkG� U\wm,�7Tx*� �wb���&�+t0�]b����@)�>(�Q�ˍi�S[�:���ӽ,�p+["�L5���-��!y'�C�x�����\T��uu���tݡj� �D�X��	�Y��6�f�6���Se�{X�9����1u�^�J�B �n®nBm�Fd�4���� u�!L�%$������iU�RPf��NW���R��eG@i��$���md�@�9`%l�g��x��	�����.K(4^�-w�����N ��7Rf����K���`c	th<M�h��nJVUQǃh؋n�R�ɍ���2��®\���"�`f͂�!gX�������F�ɛ�0v� ����v�:Z���^��z^=Pm�'��q8�]*d�U-;f�{�i�\{�f�����0v�����2��a�v�T�ĩ:���xQ@�Cjh���E�,B�fdv3�#��z����)\ڱ5�i�kT�K4�ʰE��H��U����P�x�Q@JU.J�e'�Si�ӯVJ�!o �4ۡ&�K-l!���ӽkt֓q��Pdl�1V� ^�tdˡA8�'�d�[�-Q���eC�\�����V6+�Kiŵ{�MI)�����
 �Qn���2YZ��)�Ǉ5�ylh��B=U{���d�V��*�@T��kj�Z����>;����KxzZm�[��P��kN�XZ,�EU��[E����O1�-��0Qݹ" S��Ж�拖��xŬ����z�xl���[�Z��3�+&�8�Ԕ�@$��4�iu�j,����n;f�M�5�IE}o:.�0�ȳY�Ș��7�HY�k�;��.;-*K�p-�Y��zB�5���6	�N*h�-,�*D2{cg�3�{b5v�d&d3��4���ch<��Z���sD͗{I �(ʊ�nZ�T�kRv��r�#(��#M�OP[�4�0͇Vհ#�Xpj{��V�*؅��dѴ��6�'Z�I���Fm8`n�l�=A������;u��$���&ip�,�-�:��@WW�ڎ1L)2iNk�+lO��@:���t�\��a72^�#�_
�����Uyo5�+t�$D�zr�I�`&���ڼ��Y�l���\.��{O2^b1�v��/��dя5�5�CY����S���YW�`%G&�
��]�GP	���e����Ŵ��K�.-1b���4ۄ��/C)�F5���!�^3Q�q껼�v�\rF�ąY�4�ݺyo�owe[��؋�l��n8in��A}��%Xk�7V�b����.�T�@�/]��4�ǥ5Z��*���H$�k��f�fQ���F!Vs��ڻ��#T웢6Tz(w0�f�$�yV��̽��: 
d�R�\ǌ,�3u��I)B�M���)��V�dH�L��Kb"H6hRe4iX�%p��eZ(1�;V`"n�Y�ժU�rƃC$ev톭�b��őp�[U��ۏj�K:� %!� ;bhu�E,��3	d[�U�"k��4Hc�Z�Ayl��Pr�"���̼�On� k�6�K1�!����ke N���M۸�)q���n�r���෩�%uc��ݛ���ʙJT�[��P��B�t� �jX��*��� �n�"̗(��e@�����k��gڝ&4+r�"cMa��XC1$�t1=�t�'oJ��-:#�Z�}z�֩����:
7J�X�F���\(R4�(�Ѣ��Ǚ������R��7����Z�NJw*dg%�0��yF�*vjK8�we9X�o�84�/�{m0�)2��N�F�J�Z��nH���z��Q8�C�+t�����j]^�
t��6\ǲ=&�8�&�Z<��+m����Եh��DI�bg3e���I��<����ˌ�ؤ����P�0N"��o.��t@�Ԉ&��jeh��M0홶�2]J�����ް��n�,1�B#��Y�ch^Zb��٦�]�������2�<�[TwÉ�CU!EB��z>�k[Ąj��al��c�ɂQ��U"�b��Ƌ�� QЬ���]\m��3�G�h�)h�#��j�M��F񱠩��� N���,f�{k,P�C�7Iud+�V�{2�RJP�w�U��\�e�1��j啮M�/�W���a�I
�L��釛n4��41(г��-���.X4r�عD��PQAqY���*[6���{)8��н�����n�J�r�[my��Q2��	,h���@�'�K�F�/	�8F�[��Ą�Y��h3�2mk���4�VE-=��bh@Ę�ͻ	:�)ڥ4=��[<�>��N��)��+*������/DY�oL���Ś� �Z��p��;�ӖJ�1y�:XUۍ���mQX���4Jmr��Un�.:������^%�P̤��c�Q��@j\t��ҵV˱,�4�"|�v�!5M6�b��m^e<v�A��.XF�OZ��Z��E�6��3���&ŷ!'Φ5#|3Ҿ|�,~��/�s��e�[%�Bh��cS��͍%��6e^X������xk
��Dh�X��֚Gl�h�c*�q�'*`�SVA����Ԙ�,�.ٛwI����L�����w`�i��b(ɰ�d�����n�cՌ.�4�S�UfF1H�*w���ګ����b�5�̥�P��eB�hm5vCٚ�XbL�_�U�B�N�n�*��D�_e�H��M$i3m6S�Y��1�TF�6��SR��\9kvx\y��Km@�˨��r���=8��е2�\��u�*Ǜ��J�SM�]�W��KU�w�v��ƚ��Q֤�7A�&�CO�oA��!u�i���Z�n�lc��Y�0��%*.];^�R<4�b�GS ��-�p ����W�llC� ���=�S]"݋�r��ź�lw5�丯jbbi0����n��2�7Hb�*�l��]���^[�Y�H@g�'"�i�1Ռv)�	`�6V��I�&` �=#�B[��j�L�C,�����z��ǚ�v-JQ��]f�`�4Ҕ�0`e��;0fb�[��"��P�*f[�"׸l]cj��UҽDb�u�ވ��HKD=U`ۧ�7rQ؆k6cp���`jÒB�v����7&�j=��J����Y0����G"ךd��>�E�Nwq���a���{$�A�r��02�*q2I��6���[�	�ʻ�h`[uvj"�ʳ*I{����n�}�*2�@�����[p7DXe͡�Ij��2�}�De$�)Լ�	���[��2cJ��0��T@kn�UAFؑ�E�b�+H��<ˤlm(N�q�t�deL҇�^�.��Yt�Y�uRM���Tbm�J��[kE�h���VIv[���Y���v� �՚�n�ܬ*��i�5�o1�5{�M�[�:vjɣ
��l"��;O%�2���1�S �{!�����Y�v�
1[�Ժ8�/�
��$�7b�<�SC�\b��Z��75b�����Ż��+�����-S�A����p=�j��V6�{��
�$�9��O=Ѱ�f��"}�bc���ޱ(+�rTώe��c�lM�V�h���I.�<�
�  �5c�h�R1�`Z���@��K23z(YN*�m�?��8���,��Q�&��;�@�2Ek�(�4e��#��1�r8�"�Ϥ
]�Ֆ��6-�j�)�X��0� ��X����8�=���\v��2��P!��5+qT���l�t)�H6�2�2�ˤ�'�8�Y�q����8�3L�Xm@��47x���� Hkڙ�t���c"��	�A���ht^���,��m*
��!��6�#ed��Tc����(U�w���O�JT*�X�H�M0��+N3�KQ��U� [�c�)�4��Yk@���y�)�:&Y����Qkh�#�3,R�yT$����X�I�j�Z��bhh�u�{Fi�WyN1)-&n�,��l��jg(�s0M5tQ73X�-��R�gb 1{i[�kR�/�,�X"C73Q�lO+`�AN���*� 1JfP(� Ygi�6�Q,�.�Kh#���9l6]D,��"2�=�Ä��t�Im)zv����B����WCQ�+*Mۛ
�[t��6�70���ؔf�N�RI�3E����&L��i?dtf��Q!����UY��Q�����`{y��@C�`8`���=�hI�GQ���$'5�,L$�.��J��l�*��h\����tlJ��Ҧ	S1��O	���6����$N�Z����V�m��Wc�I9��	{��s%*�L�k��4
WT��jع�N�&��wPJ�����k��VW˸�/�Q����CR�=��G�^梦�*�W�ؐ�]�l�x���u<w��8qsPYJ+�%��<�s�u�ի�ˣ� �;oe��7��� w)�N�m���>�Hu�8g*�4��Ê�$���8�ȋ�+���-J;��@���&z�3v�m�2&���FǢ�#���h����V�gPTn��M��ٻeS�1�y�6f�V�P�1o��C��m�T�.@9��o���t��kT�����<	W�d[p��n�L°�6�Z�-bi����=Gp�tEdo.�(N٤V�Gv	d4�=̻�'TQ�t��:�+T�Ez���)B���9�jP[Kr�BB۲.VDxJ���n�+]�tV!�;�N��-�i�ԅoV��Y�����4�@ ��(Yu"�3z��D6�Ke32|ͦ�U�Y+Wg���"G�]�ީ� A��_#�-�h@L8-Ş _�a�>�����BZ�����+�=�w�jPKx`�H�K��0Y69<���z��_GK�SrG�|ET�vF�
���{�N�'�����)r��c�֑[�Dh�r�q�4s@�W�Ca��6r�KIc��z�g�U�#���Z绊Ժ�鮥�-����WǶ�iZ�#>.�w�TI�ۣ�k���pS�Md5�{l�MS6�=q��5�9��^�6�,�]ȝcƞ�-�C�^/j�m�L�k�k�{�p��*��\�v� �>S�C���TxK줔���h_Xyg�� y�K3�c݃_���m��%ձ���i׻x2��o����XJ�:vh�;!�]8����u���z�Af�����2孋<����N�-�;��Z�a�{�Y�WA����7v�0����*Zə�=\	�5;v��y�hCƌ�u�`λ:oo�#���}^g,yP�	PM����E�������Qy}�(H��v<��*A���1=�W&��u5����*�J��#t�Uvr]I�b�ZՇ����4�׬�&���6�'U�ቊ�+�m
��odTKK|�6ouҠ`!��Lu�Bz��0s��|���G��*�s蠶��Y���hWm�+hcU|z�~H�5x�/VVz˼��^�����lk�{v��O����Kϖ�F;�Wuq�&��A�b��S�����X�J�R�2����x@�3��e!��0(7:�N���M�k�p�Z��ۣ]s�4��]�b�4檨)+�!w�n��I%���Ң�1��8�]�w����*�LNӉ�9,��i��8�ev�8w��=�J�(�����2�b ZmJ��̈́q�̶���.���҂�JB<�RN�ug-�)� .٘`n̓E��T�v�6T�z��"�q�Rt6;��!v4o�p5Y�*��87u�Q���|�a���r�,�����3a{�=�� �.����j��<5<�/{lY6��6����Ol�gXY=����{A��}�.��K���#C�������$nU���Kp`t_m�o8��K�6�cF�'ʺ�S��N�2R\����뛷CGlڃ@\��T����j�ƌ�x'�j�L3g1��/}���[w_2��^�oV�{*�݌h9%4!�Wy�ӌʩ�.,���YM��V��Z�8Mi{�@�t�q'��,��
7�����ɷ��<_���S�<�4;��h�G]Ko�wT@`5x	�����#W�	��v�z���.{�����^��+0`T�ue3�/ :���;V��>촞���V��[=�^��.Vb�74pU4)���Y��=�Vz����*����[�m%ݔ���4'(��=��ы6h���X�������	�����p-z2�;aF���� ���y��Xq]:�''I2d\�N�j�[�]gS|7�.�ʥ��r���t�Y��sm�8�t���lX�:a��{�^Р��+_J�mM���B��
-��7�ٜ`:~���ԟ2��վ��]�|xP��֖P���+�_a�\��;���?AGk����'6�1z�e�79B���Մў��lv��Yc��9�e����DGAtIOA��GӋ3���#p�BX}���ug�
�wR�<=�x����s]!tD���s��Vp�5�S�{�z,��57M�Q�Na��ZX4����ա��f,��˭�g9bm.������9���o�;�f�g��mݵL{�Z=��}��-�ao��j��=k}�qu�U�-�*��մd5����-4 ��c��6��O�b�<}�o�"҇��}�x�7��h>����a�K�l����������<���ͫBf�-�'8�N�-ge�rޭ�i�`�ʂ�$��q�)������u���U��@9�c����H�m��VB�R�w68��ݫ��0_�奣�N�oM�{��A�'XV|5��:���3q�n�_.)���u�#ٚR���c��7U�P��j�;pU����M�ܧ��v�Mñ;�j��.�M�c�\'S�s���=H����5�%'�{L�J��XZ;�����=[:��o�v�ȵAOz@{���U!�<�\a�pN�j���Y��^%PƋ9O����ȅ���\�9�4��++8���x�G��C��{
	���?U{�[]{��G��Ѯ��
� �:D���ճ<�#�y��yN����P[�8>}���.�V������|̵St�{i"L�|Q.kѨ?^�6
ȳ�)�����w�pyN[u-��C�R��<e���{]r�f�����cE�ѻ������裙�ln��:@C	21`aĮ�
�Y����֦�E|&���^�~z�
fܱ���i՝�>b�rm
�7w
5�Z�y�:�]93`إ�ά��.HF:]궘�[1�Y�V�y��2C{V���b%��b��Ӆ6߸�+Z���i�^�Cu[uؤ����_����?�h4BN3������Y�x��z�M�װ:n���3�r9HK��9�c�6g�`�h�����;i:�}j�Ɂ&��̴9TS�7a�L����|��UM���i��e��S�|�I٤$S���j�J��Ǒ,ʊ���U��ؒW�`Ǔ�]�O�>ۅhd���ZJ��>=J~�yo^ԦF�D��K	5�X�gI����v֦kZ��N�I������
���v��A� �7�9jY���os]Ӧ����y�u����0qYX�ʻ���,��`�t��Qk�U��/I���N�=��{���d8-�]ׂc�4�\���B�h������c�}
b�������g(��R��Կ	��(�wʥ��_�xH�/"̡�s�F-��M�;�T�`�0���m��e9�<�kI�o`Fy�n��;$�ov(�� j�v�H��c��h�)�Aj$�#�j��@G)�st�6�:<PV�[@�e]$�Mk��˗pe�%j�z�'cs7�%N�[Vb�ԩ��TĲ[kk(*����]����&��g�����7�LG�׻C�7$�/���{Q=7z&�X���`r�SW�z�=�Z��i-���P�s�rm�%ʗ�w/F.�F'w�����)������%ug!�0c��ߙ�+��4R"�yꦑ��?V�gkt�6��hG����1��h�[:���s��S�2�(���.3�v�q�ݚ.��>��,�4l��VýYe���n �9(P�*���	H9v��ӏ-�e�, �yy�5ţBĴH�[�W�o8�gmͿ8��+�^XM�~�0���9s��?L�h��l�h.�B�*��R�A̵F�����V�����
˚�h�H��Z�;�ɻ�o��p��f�13�4��^W}΋�.gJ��½�u�<j��!4Ӧ��Yr_t:�,)Þ��Ű�8+��`G��TŘ���Je��l����Pf�������^���fN؊�oi�R=��R�er���K��f�h}}b;��z�"����=�D6�!X̜V���l�;6�;j�j��'�w���Ӫw����J�%X����R�z�@ު��/����"��I�Q51ZG��6��D�̓ԫ)�ݹ���Uنъ:�����t��ʇ���SM���[t���1�60����}�e�ݏ�\��R��K�5Jd�>d3��ZCuq�6`�w)��[`�P9��m�rV���0��@�)\�1��i+!��S���h�c���p>�ĵ�#�f�Ns2iJ�oQ�@Dt)���Ɋov� ��&�9*���+e>sD�0t�3�O��=瘲Ԝ���!Y�w/1���\��n�t��[�k�H�Wr/�GgcC{�X���=.��rw�;�=�l�S"�<������nf;2u����.�M٥�iտ��Y����g�k��3������]'�n�y!�3��}9�����P�QY�&˶�Hk�*�������}�|�e-�EXn�V	����8Ԗ���IEv�A#֧]��{���(.Trڻ�G[(���'z0�y{s^P�Z�����y�+� Ι���c���ȩ3�^�7�\>��f���u>�{�(�:86.
0���l���.:�O�*�����K���5�4c¤�=�`t�B.�#���˧`4�)������w�D+��:�;U���=�N��4S�Y�g�����ۼ�֬ő��������ǫ0�����pdfJub[Vi����\y��ޗI}��f�;<�</˄�v"�BDJߍ�+�2�ug��g׽��z�IL�yS��Y�a�g0$1�:@=����r���a�K^���f�a7fESV� Ҥ�ܴf�M	�q�z��^�؞�H�,y�2�4�5����.[��<��ضy�ܧL$����j��z�ڤ�թ�9�G�bS2^��v�	�+	��[���פm�̘p�PTwJ:���YЩ|�4m�P	&�*�˽�I�m^;�J����w	���In�^�]E*�8�벛d��WED�ސFݾt��rj�����6**9za����v���"��:��7s��3��,SjpbE���pZ�+���Ge5��8~�+hԑ-�-�î.��א�7q���٠�6�J=��}��T$���V0�+.}�\VN\�g�rdֆgn�	t�d��uZ�Qm��O�t�A�m9|�\Kȧ�݂�'R����|�E��`s��fn������Vx�<
������3d����x�e]4Qmp��sw�d�f�Yk 6�Z
�MIM��`�I�@��篽�³n;5w�~b9�+�R@�Ҙ����O�K�C�c�zT{��g�n.al�|�XcQt�~dm� $y+���p��3�Iu�Z��hĜ�<cl��9� �l�kcR7��Z1v+8RtJ����RS��]��3��嘀��i;��N��f`�e���q��]{Eb�ob4o��u�����,+�$׸��ݸJ�7�r�}��7�^s
�Q�ur�F���P�x^���R��g�]�vOp�O F��A�g����Zhe�����b[�؞�tf�h�H�V�g#
+�a/w]�$��G��Sn��\h;���o_�Z�N��c.�?&��`:���r�mY��	����7(B�!��>|�`>���,fc�,�@
z1e<yS&��5��X�D��F��6q���{$(������G�{v��]�t}�(5�
zU8}�iI�f(��_v[q^�D�&�n"w��ރ��ή�W���b�\�ĳ;+�=��ӭ��"�����a�N������u�y�X�-eM��ǌ�ԕ�Ʒ{�p��˚r�Jxw:\����)qTUu��J�ٗ�Z�{�P�� ��W\&���H1>��{Ë���W�4U��g�1��Rޞ�4G����*����N��#v����(!�*��Kݭ�fv�֬����3��e\k[�������Y!(��. �BC��E�R��{�%�4�}il�<r�Y�#�X\V��;��H"���$�ٵ;�}��:��s�M����x�`F����X���iY4U�CQ�g*�@��۴�RZ��Ep��oud�Uv�%:n���4��/��M���&����C��e�Ĕ�2�~:�d�}��BI�]'�|��:������ ���靺��e�s�E:\��řH>*��4%vf��d;�S�Q9Մ/�H��t}O��U��m#�1/�j������s�\PH��f��v2ў8��#)L�ou˖�LjT�
Ϋf'Tm��L��Ӱ�+�i�����#D���=�Y�3�!G�)�R֦x��)�|oz���vx�����]���F��(�g+ݖ���&ͼ/���C��������ӏ��D
F�3u���Ɩ� ��%�Zb6M.K���@,��%9[��3��ԳsY=�*z��e��e���g���ܻ`�0�g��ٛDR������]8����Pg��FH���
����s�T}���o���X�sEƠ��9�e��g@�d�WIi�V��+cw�ä�_�`�#Q`�O��Ͷ��*b��}��N����iG*xB�k�j�I���|�e #v�2�gKK�&i��c�{fs�m��X�{���j�嘽s�Z�$%ԫsU��:Q�Ïuu���P�\p��v���hMa�ى�͙�xJ8d>�\�;�.�PO��B��R��j����͇Tv3go.�S�1���9駏D�$(PF��y�,㶵�ax�N���^wg-~��!^����*��M�ur�{F��m7�>Ǜ8�D4m�OnYL �;׬k��=���uR���U���`v�ΎZ��dw%c�+��m�r��~���vڪ���ݭ�km��Ͼ��������-��
�Qv8���k8�v[X��y2�o&�i��*����X�w�9��N㗩����5ncTL%+q-�Yp�������8����N���Ȧ��i]����A�<p�gF
��{��Z"> ��lt	��vK�ٝj���/�"�X��yJz���1���簒�~��0_�{�r��>!������u�^���w��/ޣ&�Z��oI4��'��Hd�挕j��CgT���B�o,�wU�V������f'a��\�A`w�Ð�,�e��yv��	��q&�W26)���SQ� {kGm&�O3T8Տ������?	G�N�0��҇n���8�'v>u�`��̘ٗ��%?���[�׃'��O��}��fBR��b�\�-X��e����X9�m�h�d9��tܛ`d��JI``Nݗ�e{�OL��e�b�)��{-��}��}�ބ�hW|-�ml�!^����x�����O�ϴ�)�h1�:�.�c�=��eg\1���^["�Q�`1�t�9���6�!Y�k�[rgf�j�^���_S�����})��輐�!�I~�����i��C}�}�9�`]��;�Z�9O�<�ʁ����*Kf1�Gݫx�e�[�%�D�V1��k�y�_2�n8'xyaS���O,�n��Gk�	���#�� SKy;�9�n������3�Tɏ8e/�r�d?-ފ�|ޕ����"�6Iest�����7��lQe�͕kwmMRT�+���{'UԎ�.ҧN����.�d/0�N��4U���(���'tX.��+-8���b����o|�P�-h:��vus7B��y6��oB��n��ӜƋ�f3QMYEE�)|�=� /TY$te���:CxMA� |��`M�4�०�V4l���n-t��Uܭ^T�PR���M��<��P�D��?`j�:kl),-�g1`�*%�Ab~�X�	��iP�&#l�\�fI����e.ш ��)P��}��1��
�ѝ	;`	�� 3���J[��	�]�˳,��qf�Y�_X�����`[�c]�q��bg ��I�9�-s>�=n</r��w�w5����b��K�O��b�ï�:��,qo��ʕ��VIi�g�M�dn�.ѭЉ�ݫ�|i>pyї^��a�r�q�F5�M�4aJP,G�M>`n�������3U��z�9�6�T�)���qj`ӫ�����`
z��^uC��X�n�6q��P��(u>%ݥ�ң-���,�l�����T���h�ĩt��v7���
X1i�6�Ր<=�\����e�+}�Э�Ϳ=AuN�k��F�M�e>ݫ���r﫲�R�J7D��A$ֻ��;�a��ۭ�AP'�(�=}Zq�:G�:>�QIξUط��1nVu��Gv������}ye�������M*cVV�^��f+�];�ؗ�-���'��,]��;)���2��@�q�8:|��Vu6�e+����0�C/;s���z�%ۛ����8����g�e���m������Uf��3�6;+uZ�~ng�X�<ΰL��v��۸Xt�^G"�U�Q���|!�Ŵu���_O�g��W�ow���典�g�Ů׮��]VF�F8��9�1��#`\�����'��U�2�@սJ���)��f<X��u.�	��,���X�Gi@uL4�SQἮu�G;2��M�P� �x�0<�Y��qěɁA���e�M���]c6qI6,��e�O�B@6�����Y�ؔ��AR3f�V�0��W�JEb7mI�����F��ՠh�(nGB��&�u�4]ل.���c�m���K@(�m�~�9h���S���t�NKa#d*��n�;z�Yͻ�����GԆ+��t��[�|7��Cj��a"�U���k�L��t�|E�>�%ܟb::�w�X����K��+]A����U�F��_�%\O�ʒ�6�ӌ�<��&��R�"���qOpkWk�W�A�J'�
N�3,�-7�;�'��BQ�(�3���F�c�qu��dٮ��E�Q�����Y�un:�
���VȺ���"�����k��J���"1����o�P��;/G|`�rx�e��������L���_��g��}}Z��0-�W�KxecQ-V���V�z����ΚƱҺH��a���j�e��L"��zT���y"9ԇ�:U�5�m�0�
K�]�/�u��kYWZ/��g����e�FZ��Z��AW;�Lޠh�n�)�����`ݟW�����õ>�Ǻ�Q]��;�T:R ö;K].��ۼ�.�x�N�#�ɭ�#mևyE؂�u��+ǵE�ų+X�֏h�*��3F� 5����X���Z��Ӈ�t���1�V�/c�u��gj��-O��7��I��<Ty��|�L���a=PE�qT����Qoʛ�D�P&�m��⫨F���-��e�k�
���:�db��7s�CM��fJ�n`߫��C�Ep�v��Gm2�bZ�xrR�o_(�ۧ��î�s���#��?:	�7 WШ���4,��Η�������kճ�.�0�#gFsT��m��q��#��	7W`�ɱC�<

��̞��ܩ�#}V���;T$K�[��E֧�V��lRU��������q�l�J�tMv�>��5.`�tJz7	R>���=�s���j/�V���dq-��^�G�"a3�+2���1'����p�%m�	R����ufǲ�p�s����{\WW7c4�R������[�^q�Y�0�m���@���c��4��K(�:~]X��w��1���$X��x�����N���N`K��9�����̛{Ѱ���{���23�zy��;[��v��J�v�6�:�F�V&�ie3g�wyqG�2~��k��	x�o��Ͷ=�¸e�c}�X���N`��;�DSv��|�/�ʫ��|5�XB��ii
�;����>82Rjk/���T�|���՗8d�p�r@ԓ4��onv0���%|n�_`�Қ�j�ٯ�l�Ӝ�O;V����6PU�n�t-t�t�i��	���_W%�룲��e�ItO�ԭ���"�;4��of�r�1e��6��3֓��;�|����1�ͨ%��u�����řa��!c�M.�J��:��,�ϝge�¹�
�2掘;��/?C�Vk�i)ecҹ�kyګ#�;�q�NK�Բʕ�a�d�R���9O�F�f3<>�g��� ;��"r���P�Yp������/Ȥ��G#@�Bt߸���h�.o:����8b�ux'�y{�k��C�"��ܩrAs�g
��Eu��mw:Օ�V�t��c�dvmc��4��]>�o�\�������ށLSW�+k")GOL�E��LSrVj��,�*}�vJ����Cf��݋�5��/�#t�J��>��2��`}�I^�(��Ϣ�u�t*ѹsy����A�-�/sa�����Q�9�j!��iE����ر�h=*�[��X�{)�Q݊M>ߺ(1[��:#��w5"��j�+Z�bԾ�s:�D`����"���H�.�oc��U�dA��x��ʛ��YY,q����-�$9��o�y��luek��m�Վ��a��r�ʹ�:������a������v�æ���6$�8��
D<Gd��0������wo��O�{m0~�|q�@ʙ���\LB��B��HTr�<�"��IՆ�)�L%��v�O��S*���e��u�߶�rb*�~���8^b�7��9���1�@�0[�x�۝��յ�kY�t�Ӭ9�����=�X���Q�ee���3���O6�P�㕖�"L�`r�^�-ږ�B�4y�ȭ33!����k��vsU��Ii�9������{�/�k��I\	�F�ː��w��;|�-�lS9yc"0r�̗n>!B<�8U��tƣ�rD�v������΁�ywp�60�z���C+�.�u0�Z5��+ir��_gI������&A}Olu��\������ 	�nm�jP�S2��p��>�ec�H'*�����(M�vУ����ZW��D�n�����4�˹V��rRF��쭲4QǏ�f��p�l�<x�%�;O�P�U�Y"8t^L�ȃ�;At�U���t����]����k�Q�C�J3����6b}�r�EL�|)̃(����ɞ�2*��3�۔iZ3ՉN��R�t�m#�34_1.��k��	�,�eu����JH����k j�P�5,��4|�&PG���,�;�w۸�/��JJ�D%�W])&�:�*j�Z��p��N�x�coܗ�D�:���������KFƸŨ��ΙǞ���wO��i��S];:��pM�������W�q�|>n�,��T��j�nC��5Knc� ��c�FiFAJ���p[�u6U�ϩ��M5��O�+x�.:.�zj;�[C�ЍX@'�u;��`��v��v�_�yo)��i�^B�"x�U>�9����]*Ne��#��KmN+J��ّ+��_'��`����1�{(f\#9�;Gwf�n3���ԋ�$��J��$+����\z���C{w�S5z��� ,���7ۂƃ��%h�|�-<�����C�j�6��솫�o/��X�5f�;��p���f�b�����nu���Ҿ�C&(�U�E������~[_��_<�	w��y�;O�����Є�e�(LF�7�5�k�T�]���3�}�4\�؇�>0�V,.x1'ǹ�Ϟ���A~� ���`1*�^y��ͫ����T��U��M�{I$�5�D�8V /���X�3��J��sN�:k��X���/��(U[���eL� �p��p��/QF�HL���P����r��9I	B,�.�8��{��K��i,OG���0Op�{��;���-����v�5x9�a+f��Q����<���1�C�ɾI�A=H�9,��k��ɱ��j 9��Q=�.\Qͫu	��6��
��Q�<���m���þ~9T�v%�T���w։{�ˢ���x�Џ.��7����s����
b����zS�aةjz`�M�6��/���,(�������xF<'=�!ͫ"�캂s.�h�O �H�oq���a)�5|k�����Rѣǰ��eqٓK�jwrS7B� ��Y4�� ���ba=\�@�傐/a9�u��I����{�p��ڢ�@nU�����In���5r�.sPb�{�a��ďF�r�ۤ�t[&��<{T�g4Wuɶ�z�M��q����RVo<B��*L��u{)8G�8�".9F�1H�G�&���u��w��k}/drdm[���y7��\�ͺ���\ѡ�R:r�K��`�� ��70�*����k� ټ)�p꒖R4~�����tSu&c��U�z�'g�EΙ��V'�������Oʯ$�C�"x��雃C����_ ��N#���Z��]������ ��_@��́�á��-fC�^�PQ�j�s�sp��~O���^�_K����\z���MrKL�{�swf-;��oR*��LT��!I���twX�6��IyUk��W=�Q����9l}���:����S��' ��9�2���Q��ȥ+ɫk)	�ǎ����Z�t��:�*�����9�����ل�)b�!���+��|���v˜�-�j���v�@�t��1�8���KB�z�)#�6�3Tڝ Y)9��\Z휮v���so	!X*�d��t�P�~�p6\�W����ڣ�PoEv�3�m�(hyZ=�/7���W+�������.O!%�^�=�gxZ]NϢ�J�0���f�+>��=d��/on{]�I�ڒ����y�
YCv��(m��-�ᨡ�%�F���o��糷/nq�8�"�����:���U/]H*{0��9�F�e���-^|}ϵm� �M}MC;�m��,R�BL/�7z����AU��3�v�{���\����v{�uc�2)���I���v�k����*5��(��z��&��m>��/�F����<;ׄ��g1�2Iu����|���0��gjW, �N����-"e�D���GNa7�nw<}��r|�L��1+-�|8�ʳ(־�Etɐ�@dV�W�$5���˷��x��ufY���n\)(��þy8�߭~�f�v(;D휠��C/'�=�:���.������͏
B����zM<C�Bs՛�k6�]��ܙ9R�t��*&i�T�q�\��.<-�Y|R����Z�����p�u�nK���{�(�K��w��p�:t�'����m�.�.w�шۭ��<�ڨ_d���%��7.�eC������Wqx	'����sz<0���qX�P�۱��Ԉ]���<�V�I��w �K�τ�s�=�7V=�T5+c1����Be�xM܌��r�u՟�U�mk�|��b�7n�0-9���)�����}�&#���z�4�"��?�Sk[̕����������s(���b]�o��3���,y	(���,<�EO[��:y=��j����t���,����lc�P|{se��v눌ުkYiR ϵ&���x-Z�cp1�d��͏xvaε�
��ZPQ2c��E���ot௒���}u�ꬔ#l�3�1k�!�a�w��k,� �U��c�DX]���t���ZN���Ni�eX�n��1��*0j�&����ś�e��5k��c������ﾯ��sO7p�7��~��{b���R���-��Gk|e���C�<�����caV��^#��_Bv �	;�gI��PdfC�hwř"�J��eK#oF�D�[���)]�-Y�y\��*�RWM�
��3�f��Rp+X�������Xum�c�ĨW
ym�����@�U敆Yu)�}�������:���N��)e���V	�J����3j�	�N�]ɷʖ����33P��#���[����O/vq]i;T2=�ε���.u�S�i�v
�U LaQ����i�����ưe~�6GV_qˤ��)����.���.�{��3�P��#���TpWDH�"*��,α�8��ݘR�����2`z(j{�+"9g�x;�ò���Sj�Z| �9���〒�1Ƭ��e�wSi49�J�/v}�Z�y�n��7�T+��V׌d��_Bm4�W�ѻ�	�E��8������P���x�y��7FP�{$�aξ �
{GA��Mu*P��#r	|���<���vߘ	��[KFyT�$�4��]����h��	��o8��
z��r�`#�eܾ�/��f�	\�!�)0��դ_lat���5�ϕv��s;1�7�,X�\%�l�զI�.�:]Z��.��?`��r�����NW<׹0�7eN�Wq[�eBOL� ��'�h��"��$�u\1�����3E��)6���E�j9\�7u���w��(J�r�ns`78�sb�k$[��R]ۨ1&1�Y7wa2T2M��IˋsnF���F�]�i#���]	'.N��fi$���ۗH�Z,�f$̀�]ɍR��h�5��JI���#�9�v����s$BFK�Q���Ѻp�;��,&1��]1�w]�$M���˛;�	��M�wtF�cI��XNU͍.p�DR���wZ��F��t�$h1.əwX�E�\�4��b����g��̬�Lz��{��"{Us��P�=˳�-x^�[�4V����-�b�%��m�Fr��V�����SWӫg�{�Ӻ����Ôz̠Faڠ�<Zh������'�ԓ2�Yc�ǜ�}��&������v\���c(.���#�h?v'�qG�r[T%k]*V���T�w'�w����������wy���_��عY�-)xV�\�>��{U�U��,�G�Iu�]�x�"׉ܬ�-;��ṇ�/�N+E�u�6�3�
1��AH\�8�goME�[��,{�=��x��y��Y�@#K��!�38>�ju��=�e-u�0����{�Wm��u���D�Oz�Cn�1�fpΖ�,	�W����i�{��E�o����L�}�o������"���x}U��(��TN
�G�imH},}����r�{R���T���jiH�7bŸOo�k.��\�'K���4k�_º�����0B�6�d���u�_����3w�_��1�kF���jS:	:N>�\�*�E�FrJ���g�uOm{e�Z	&Zj��΃˚�7��hq��/�Yp�j���!�/��k�g't�� ���ǅ4�����'��7R���w�t�l����ݬ�O�ٻ�\�0J���Tg{�=~�}=K$���K���vQX}�l�r�$�ѳ���ڜ��}����>��a�k,�켉�G��r{�qLz�&�[�����[Lj.+U|j
E���;H�5���9�����rY��E�t^߯5,R5��x��k���p��o�%.�J�|%��6����3����Rޅ��L=��gDY(]��܃�v�2�`j�ٵ!�5h3s�ǆl:�ܱ0%y���s3�P����W@w��,BA7� O�JE�[Ӓ�V�n�}�+���l��N�\]"��G�����xp�`�E�C ���`��u1�Ev�G��?��gY��z#��y0:VӤ[��A�}���E7)�F�����x�_0o�z��^�m�~�s;�V�v��2��@w.z*��\{o.N��/���&��|�H�}���g�����3���O���1�γ+F�6���^�_5��\I�����>�݋>���O6u�p"�:<�Å0t��G�J�A��qH:l�uo�����Ҹ�3��~�+�&(�r�$A�YY�:�@*���u&�!��C��9�梫�w���W �l�mׁ���B��X(��0�Q�މnR���sͨa�E3#�IVQW\�����U�'5xV�����9��~-�GH��X����*�F0j'1ut/lq�m�Q����z�E�1��n�o�ܭ�#]�f�yiEo7���:KLΙ���z����[P�}(��<@����{.��K�����+N�T[��h��
��G3�gF�%��>��Z.޵Z��u��)��ZwcSttoגt����(�t����ˤ��_R�fZ�͗r�MP�4mFP(�%�F�n[<���ߏ��<)x��A�ExnAvI���i�ı�U��G�J��o-�4!\x�c������|ڨ~�*��VC\�=�+s��	:���V��F�pt�Ѿ��x�.^&���Ԭr�Ø�p�Է�0���vֵ��&e11�rr�������yn�1Y���ư�q�dq�@��?ۯ�e�=�Prl��Q'0V�&����� BG�ǹ�cx밫��n��jKZW3���w�;KW�]�K
��^�W]�������春|���G�B@�7�E:Ex��&%%n�3����������ŔPD�?����|\ƈb�.m�̀��4=�� �R#�pS��j�C.X�7�__��g,�4~G�??[㏸����&+RvY�s1��ȨN��)��%�߲�����52O����Qy:ٶ%1H�"�2�JN�ż������(1^k�ȳn�W'I��cFus�u�ݜ�]�������f���=�6i��L37%.���l/�^�U��*��֖[�-Xf/)�G�ұ���34:]J�}��jq�s]���g����{k�^�����}mH��,3M� ;
~�߽��T���d��V���B���w�!��%G�=������\&o�>��,i��o��4�t�}+s&g�p������:�TpD��
Y �=��s���Bȳ6����g�&��L��$�bO��8=e��B�S��s��LH�D.���a��������X��GQ!�<��W��D4��<u5���X�7	�}��3f�P<j�f�s�ӱ��mf�dn��N'����w(�&z\�gI^��#�9b7��l)"���x���b���3�c�b���ɺ�g8�A(�V�1jD9rی�o�p#��
)�gs�s���P/���������x����Z���h
�~���Z�%4��q�4f��yD��X~*к��k+�ޖeH��^R�Y�t��~��t��2�^��>Su��,_�n�{���ow
�N͠���'ב��s����%" �;t	�L5gJfє�*x�������z�e�/�Җ^�z�]�F9��d�(s��9I���%�yi���јN,�J︜�ضT+�
B�w�V,k�T�m9q�ۃ�O�3�G���'V��K��,E��,�̵���/f�e� ����ٷ=n����u�WE���l�ם���|B;Լ���/d�J����X����Z�.�삲�[�B9N�:�h�4"�/
͖z���]�_��q�X�=�F�ޒx�)sg�� V���w墶�&q��<zuFа5��zh])�2�Ch�ʵ;A-�,�1h����m�UAM��=�3u�h�c��"�D���QEx��J�7nB���u��fXy������5�O-��iG�A��Ӥ>z��f�Oi���j�q����p��A-��O��G��lE�h�-8J��VQ�����ė_.����t-���RqG�!�bV�Ҩ4,�&���θ��/&� �hG�6���C�@:5|@���b�y�J +F�mY����]�ȶ-c����S%�VӖ��a��/xC�}�3�37�Q�TAH\�8�ԙ3x��<oq̹�泬�iu+�Ꝝ'0�=�e��CUx}z�k*�3|;��Q`���!��'��$��*�������ϟ����vp��OoX6:d=Y}��bq�sFڧ��u�q�.=�C�L���Gw��v.�%>%����5��^�x�]:l�u/�R�Pt���~��m�.��|�'enC���]B���ݹ�'I��ޚ���r4��Ѕ��6V�Vd���/��շj��H���p~��)�	\u$�',nV�J
ؗ\<o+W�;O+�ik�Q�da�_ӰOe}X� ��� ,�{�&/`W��Vқ����C��g��[^�~ڥ�Gn#�G��+_Α�it+�oixlPhhV�ͺ�{z��R�?1�7pً�j��]�D����Q��i`{]tirO~N��ִߵ������f�*j��ƹ����p�F�{�O����`;�����aڍ����͈ܘT�j2��}"��_��u�����o{k�^4����7���'_'�v�~@e��?�� &�[5�
?E��yg;�����Kk�� j��h1��2yz������*��ק��sM|���@�<$�@W������͸!
�ա�r��>0�dqn�T2�#Ki׀*���J������0�=�ϙ�9�T޼��6�&����V/@��XN�R�9΂�@u��.uL3n��!x�>ϯ�z�V�zi1�B�D����x	ܛ��6k�oj$j)�G~M��:��_0����1x}��)����Y�v�r#�B�8���6���Y'�,�;�*eg^�����@����v7�Qz�����Cm{��װ]�&�YF�����4���(+o����R��&ž�����B�y{������NzD��S����&�Ŭ�w�K0Z��w��˱���q�s�[��˕��6�w�}Ⱥ����vԗ@gI�L�_���p���9�nֺ���U�
�0]?+񩇅�A���,X{�J3]J{�"��ʞ6�<�`Ůk77�$�-c�����Z�_�ݚ�C�3�ʻ�<[����(��ݎ}ֱ0()���������>�����q��ݰ	,W�a��kR��<�v��>��hf7�f�JxM��0��w~��]nLU�=�F���+�^�5ݏ��9S�-T�;I�v�j����ɻs���]這> O�:�FD��YMtu3}��a���b�!�����f��=;ܽQh�V1v��!]qZ�Q,�)��������"Y��A����x�f[}�]ۥb�
a���UJ�4��[.���:C1�|ڨ~ߊ�#���Idn�[8�3�	�M�q�X�xO�U���o��u�BR��bo�{�J�!�#k]p^j�/]Zm���ѳ�*�N�Y�1ʾ?��@`*=��.�)�����{�`qz�iAK�dS�����\����tx�X�rq��ƦVDp�=e�uuf	Ʀ��y_�h�odj�`�+����Fѷu���N{0gD�0�T���h�6��^.pQܨ:Y鍏���FN{z�Y�ns��ݓg��p��,v�VG�RЕ�Wo��q�liA���oM�)�&��.n "<* �P(zS;X&�*�kXǫ�MLځGk��j�9g$s��X
n��SB%)�%��{T�@�|tR˲}�cCNz^���	EҢ�����#7+�C��\OW�;�x�>�n�z������f
�����j�su�!�.c������_f�HW
tT���'e�s1��Ȥ؄������W�ϫp����}�����z��K���!y��a%UAn�� ��jh��b�Y��{w5|G�ꎆ�eϨE^��Yg漮̪g�{%CC���'~�0���gQ�wI��~�b8a~<ŊW����4�_՞@�`�=��r6�皂,�7���{x19"����p%8'V�d���_�ꘝ�۞��2�PP�#�R�c��X�
^$���^��z@#��T㡙
3�(�]�3���*<i
w�,'��]Y�aNk:v{�\�Rl�Y���%�؟>C�L<������|h_OWr�1D7[��
��bJU��]<�#׌}6�6�?��Y�ɗt�yr�u�{՗W�!��t�:�Y��s��$�{��Š�loU��嬏��Ќ�!�,���i
[Ř�
*�4v��u8�ٔ9q��o���[����#�6��]J��ǆ��O�+/�X��gD��b�.C�ʴǶ�U��Yb3�r�ܧZ������3��$�Hs��yX�	�iW	M/i���Hѹg�,gQ�	dnܛ�vV�P���܋�6�����yZ|�D#�����=0��2����\਌��[��Y�em��y��ґ�s5k�΃�:��u�y^�:����W
@��� ��C	�x;N�����z�b��#�y��Y��������}�]ҍ1�5�lr�Q4#�dD���=�uAy��f{V�iD�d�1���sQY��\wWrU8֯z"��uT���4���S��3}I�q2��E�(� �}jz�V���}�3z����,�A1�����DUO���>�ڥވZ���1=+G�0�ШJ^15���ڐ���~��i/��s.`7�*,��}��aTk�_`��MӣC%ةeH[��1(q��E��=;�6&we��t���{¢�,�\�ZQ���Z�;]9�:�W݊BqG�=y���W^��V{���>��xR핪	t�z�4�nV	7kn����'���)�S�e�+y:� vf�zTvh;$��`��$X:�V<XIT��\A;�g=��l��Dnem���t]������c���;���#�ad�]"ʺ��+�uwu���lӛ�I��ϖ�ѿ�"z�l\�<ť��\6P��sv�������syXMY��0w8Jh���̯D/xC���ۆ`���(ƪ��,�߯��(�-�kX6r��1sa�T�?Wӳ���2�� �g�#S�g�2��v�m�����y��kB�Qk�݀Ku�U��^���������}7��5{�p��#�>IR��ʖftw٬*]&����4���U�V��G�`�+�1O�v	��$Gִ��$Ԡr����#*ď���[�<�|}�ug�Z��^����۝$�!"�ޓM|!@�_��gsΎdwkpo�T�C���g��ޕ�����.�d�;y�5*��I֖1�BP���Oա����S�Tj�#�3��1�$ޮj�t\�di����e��JH!�6�3+N��m�ȕ��k
�tHg(ݏ���K5㥥�8|�i�):�!�"I5P���Z��!J'�p� ��0k;"YZEgC0_ѻ���х�Ci���e���1��^�k���Oi6'� nJ����/'R����ŷ��T�X1ʀ����`��|��WzY��!�<��YY��]{9��7l�`�9z�.�k�j��D�离�u�q�lryձ��.zyfY���l���D�����O��*j�nQ�\���Dpo��*q��o�Y��#���S�HQ�WΕ�Іa�><]�ƃ��sU�`$v�J��]��ol�+#OL*3�_���ǹ��RZ΢�ĥ��)Q'��%�Q��.�R��7/u0銷�%�Y�e����o��� W�x�m��]H�#�om��,&��t�ܴΞ��)k�vWo�Nܴ�M�B�<��,���z����Z�*w�Q�X��ҟ;M �e�ŒD��Gr�wCKpp��f���Y���M%��<�����J!�#�Ά�(���g�)��8V
��O�M����V#�^��m.�Ђ	 ��-�U�O�d�81�I.w����.�;�����e��gB��PթY�Xa����'Z�KWd���-J޻�fx����SPu������H<n;E�ۺu� DV�'������{f3=D�w�{-������e���������Ӓ6�9����e7Jfݽ(�u[��jQ���+=��Y�F���`Ć�}x�<��<�J��wG{�w٧���ge[Z�����I��Ԋ��ԳN�� _S)*̆͗y�0�&��],�nЅ^ۈ���r�	����zh�qx�/U9S�̑AQ�/���N�\���ܾ�&v*�Z�8V#Y@�}5�^kom=�7�ԣ�z:1ռ�3���g$]	�ݚ��;�Hd�bW��hzs��mK&-��8.��\��s.&��w��9aq���`�:�Ø�L�N3���u��9d9*��ZtlY���|��p��ñ���BB˔ \�b/t8I�J7Me�W2�:�!�$�[W����'��"�iz�����GN1�y��f0�D���;oe���u�W�^;���t�KV�`�׈9XI*�ɐ�&�w7Z�ѩ|�c���*:�fMB�i��_)�P��N��Xǹ�x���m�pr��Ç����O-�E�A�Xv�!�tǳh�(�O8!ۈȪ���fU��'f����u 1`�%b�@�� ���-�{�/��Sf',�	%iH��vpAb����>!ݝ��=0%�1Ƨ�0�]"�J/1�ᵠ�H%S�b���wrbn��J���������tj*�-S#'�H���r	� q��"�g:|�B��8k-2��e鱴|���d�+�f8�LΤ���{�(��P]������2lO��$t��mo}ᴝ�%��0a�EBŃ����r�V.T_�i=�ib�}ȡ����{맂������ktq�vyM{��[��������c%(���F4Q���4PHh0�D%Gu�JbM��\ܹ� ���(�Q���%�(ܺh�a,w\͓Aҹr�)u�XȘ)#s�u!b��I$���+��܁�1ΖL�����#$�BM�c%���QS9����J�l�3&$!I2Z�.�B��3;�	��D�ݻDi"��i(a\��E�����KG.;�b��I�!5ût`�wud2RT]݌����Ωh�@��h�S�� ��sQ�I&������2fA�fX���$� 4h����2$��]�nn�X�h�Ѕ��r�9���Ɯ�>O�WƂ��9�>Gk�N��.��%�%�'�1N��yhn��2��$"UΥט��h6��OHa$u�y`5��bpI7���i�Ϳџ�}�}�������׶�^���~���H�_��o�^wlno����so�������ڮ\�[��۾u��x�������䟠�� !C{���l����`�zCP�W���k�AY��"	#���G̀����#�o�C�G�?|���� g��Z7��o^���m��ʽ��૜���W�~v�;�~<n���^���׋}���o��׋�o��w�������o�Nj�3�����=�H��@����X��6񷿟<����n�ş;ү���?|�#�� ����~�ހ,ߐ�#�W�{�{_k|{zZ};xۆ�߽x�a�I'�	�Oи�"�#�H�wOjJ�I������$$�x|�G��">��x��ڼo�~7����������wl�D}$~yG!��D?}�����k����yoj�+��~��}�����y�_Kw����z\���_�Br�3�F8��Ǟ��F�����#���������ז�o׵����}_}���G�`�+6��E��'�?��~~�<Z>�~z����+����y������"�����a��?&��������;�i������> HG���_+���KO޿Z/�mʿ�_}�o�ܽ��|^�m�/}~v����?}A�HV�����U��:C#�O�;��ԗ�#">��$�GшEt�r|���U�׷z9T�^G���
0s�d3�(��� {��������0׻��^��~����_j�i����K�o�����ۼ���{ﷴ��?|�c����������a��G�#��ĩ�XU��O��z��������ү������ۆ�~����5�ס�ߟ�<�k�}+���������x��~w^-⾛�/��ץ��/j�o�r�+�:������\U���?E6������ʼ!T{O�2 �9_7�~�[��r���z��n���ߪX�O�~��H@���Y�O�~�����|Ȭ_}G�$����H��`����9_'}�����^��{Z7�}{���׶�P~-�l���Pﳟ�tr1�$�� �(�@��_�����MDt��������G���� \�QI~�b x�O���ίc6�߿<�^��oo��}�yW�����^�;o�W>��_Lv�pTR����[�
t��8wvt�&܊l�zE�����K��F�2눭X�!���i���>e���aò���aʓ�+*�ny�Q&��F���r��~��������8�t�9D dP��z@o�����Z��ր�-�=C����Nv�>��/
�������^�vߏ��h�����������x�>�k�
#�R�
�������ok�����^���׋�z������߷��n}�����w��\��|m�?|>��,�v�*9S�33'��?~�������k�o]��W�so��[����#�:G�[ 	?}��k�︀}}G~���[�����z���/���_������������h�vM�er���'�Ȃ4_;����W+�n��x�������W�湯Wy�����_˗��Kz5s^<W��[�{�o������ߍ�W��^�������m���^|�ſ=~�_�u.�/{\MȾ���#���ε���O��^��{Z7��~�_��^��x���EDW��o^w���ln^����[ڮ\�w��7����m�契#�O���=C�,���5�{��N�,xG*��J&�=]�� ��#�螟�E�����>�@� ����DX~��>DY�>B�>�'���
���|G�__�x�ۻ�����F��+���H���������}F{f��;N����F�h[7�G����?#�w�#�d|	�w�}G�È~��c�hG��~�� ȓ���P�yx���̎����Z�/���?z�?��/�h��I�����a׏fz�U�s�3��-��g���zT��A��4��?qO�@k "��7�>����H���D���x���� &����^?���kگ��r�_�<����oB��G�d�?�4o�)���i�<����"� ���@�_a~��Ȁ<��ɷ�szmϾ�.�����}��-��#���(|����a����#�~~�y5�}5�|^+��-�Q��]Q��+�yi���x�&�׻��Dz���A "�ޏ�?Q��}����ޗ��~��v���������񷱾�s}z�/K�o���sE_˟G��H�>��@F�����"��?_G��?|��T��*L󹼿h�K;X.mx?Y���#��/D��'�F�z>�G��oG��?A~F�����$}�~��޼��^-���>��W�}��^ur������׵_˛�{��>����>�_��.�W�aݭ,[��חjA��a�����Eb�ѳ� �7A��#y��^7�)�#����޵3�R��K�}Ql�r?�� I��>m��p�H�} ��Vw)0LD3j��ݷ�T2FQZ(�����S����֭�!�o�tte�N�ML�ض�^�V)w�O$~ ����t�D#��b������"8���w��%������]{k�\5����n^/�׾�>��7�~���ο�������|k�x���o���}���|�}T{1�<�����Iި���@����׭x�?x���痥r�|�]��IHG�V����,���">��G�����k�����W.��ou皼�~�
�d	h|��ь�����#'���7��?~� ��(?q�i~~� � I��A ;���#�|���L�G�<G�@��G�x�����QG��Fo��M�@� ��+A���O�~�X���Q~��^n9���oe������?=>m�����E���~��Rl���7Hx�����t� ^!��ۻ�������堫����׵�~ux��T}����G����}SY��?aGq��xG�D��f�"�_�缺�ɽ-�M}��6{�叵��^v�*������y��o.}o}|m��sQ�޻+����?z�_}^��n_�~w��֍͹���~|�ƾ5�|���ޖ�G����e��T�͠�/-�٪v%/}�����d(D�d"�=�� a�M���^��W-���;��o�y�������_˛����o��}�I�'��PhII4����|�X���ǆjޔ;#Ob�ts��#!��s}���W�_��{o��{����[����� V��G�-D|G��"�W�o���x߮x�{�/�x���{���7��o}^�yzm�?},dO"��>��^�z"< ��_?�z��η�[����z�6�o��I "~��>ha�� !?G�k��[����+�������ޛ�wv߯��x����wQ���h-�����������z�j��e���J��0~�8� �^􏰋#�O�E����#L}�#��84w���dc��V�>��ޫ�HEI�m�z2J%������5��,���8�q�^�dW���'�mr�+�OwnR!�>�r�-�	RO;{�[p��Ɋc�iH�Չ��Q�Av����DZ�
wG؅ ��I>������r�ѣ4W=4)�$z�R����Kev��6���)�k����*d@�W�"b����0���o#Jn�픬"�I��b�9��$��:"�R�w�!�D�v���`�7���N�A���ɌD�Y_��7&ߛu��I!������V3�H�t� 4"py;+��ίv!»|�͚�@�x'��tJ7sigr�%��g�&7��ϔ~fiD�L;:]���xZv�u�`h�j����
�۫���()�SC��qf��%x�����g�b�Ue]?Cm���������Ôz��z�8��F1#=�uB��D� +B1pض�..�=��ޒ��GO��&�F�9���=�֝��^`m�	�V�1�!�.F�1I�v�{Ok�c���.u厎�i��!��C�G�Ս�_��yY7g���+�}ͼM�=g<�IH5�QO-%[�4��n.�Vk�e�g�h�k���<�ٔ�x���U�"��i�
N7fb�x5�ȩ��]�,����ߤ���3�v>�Z����`��x���O\s;��®E�{���m[ {}�}��O?
ؽ�յS�������r  ߰w7�u�4��ڱ���귱sހ��r]�v<z���c���Н� ��t�,��w�R	�x�'B�;ɳbb�F�����g��㇑ͦ�ٖ�tH������U���b��=.OaXr�v�o�yOY�;�um#S N�X9�[�^�t�𻥱��*E\���xu����ٝ�r��9N��졎%z�v��i�԰0�|ƒ�k��(����2��}�f�����k�����z�W_�N2����l:�&Uugq��=��`�Q�G��|"�X/T��LƳRU�)0\k󴏡�>0����ר��N���w�zQ�t��X	/Jd�(i& N3�&�ZD
Μ�h�����-�M.�~~�n�v�2g	z���T���}�A�vI���\���F��8����jbߧ5�Mj=9��Sf2M6��_���M�dHB�� -5��)�ѐ��C��M�QF�J��pkr���6j=m�9)��\9��!`Jwl�U�1�#q4����v3�^淘�E�����i�ea�Y�/��v���̄���_l�@O�U�;>���c�!�V��ul�8h�ё����fh\kR���UJ�>�S��p0붤�A�����'7��7��}G� z��Dc�5Y�*��k�l?�+�Xx[��p�f�˱w���h�S�^.��+1�<h0�M�$��K|w��*ƶ�i�ט��}Yy�w:~�4�zB�Wrş>]��jܩ�vJ�p�}��Ő3�|�۽���}@+L��	O���)L4���t���.s0̾Uk�����9I�( YS�ɲ�̅���Tlk�A�[�z���t��`��6���CM�V.t�ԍ9��5�r��?���Ì����SٷB��߷���J�� �P���o~+U�rYƎ70�Z�=C[Xn^��U�I9��t̎&����#z����������x�������}ǲ��Jigk��Ӣ�kB�ǴUt�W6��w�{c#%S��vc=p���z��������NqS��0�;"�c,zI[1����n00�%�Fۖ�Ȧ��4:�my>����dSUa�7�o3���A�W��"�'�k�^�O������Ӧ��u<v��n#����eHq���?\ab��J�3�'�^�$�@��Z�K<$X�U��8�a)�~�lk~lU���x�NF�Z��p�v��J1��c � ��T��t`弒�-�̽�%{�(��=θk��RFx��s e}h!5�( 2�ݐa+�]�f��c.^^�&�Zt��f���pS��|�pBG"�`7	��i�Wʑ<5گwg�hO���x��6^$"m��[7��s
��sw���^�h�Ojթ%��;�e]� "��Cv^�pֱr���2�`{�,��k����L�ϥ#ۗP�]C��*��b��ɭS�o�|�@��x�<����V�Fo�iP;.^����p����|1���r�9'	7jȯ��,f���0���9\Ɔ/���+>�
�:�hG��9ѵx)�<�
�(�=��+�K�pA�f��{��"�f!�ҵp��c���9
�S�n�݈��*���!��o���Z��i��V'˗��F�Z����wt�o��m ��V�s�C6E�2���S���z����
;(E]���?5�vP�^�}�C�ȫP�V$��� rn|m�S�g��r���N�b�o�4)��@��b7p7 ��j/c���ӛ��i11B��������J�!���וc�!3��d�n<Wٸw�C���jĭphSΆ��&'5b�z#�w�t��A���Y/z/�T6I{�{���1��þK��_y�Q����0��G���=�|�=����_y��:��B���ҁ��f9W�Q��9@�<�.C��Cۿa�@:��e�R���(:����)�g��(n�3W���m��hT~�(�|%4��U>@W?�!�} ��߹ڙ���D/�qeD)���eT�����W.��}��ڨ��>�D�Yr�xlk�bVbwgX�#�ݍΟv�%It�0�<�[�VB��T\Ǔ�{J��s=����[�f=�a�%Y�d(�'e�^)5�E{	za�p��a����x
j���}�G�l�ݿ;o�����4_c��;��ܬ��Q�GI;Pg�!�Te"� ��ԩ����qi�`�>�����VA�_I:�s�Ӗs���j--��ɣ�y��Z����,�e��
���gmH����܈KK��8� ����"y��{�`"����V��Ȏ�q�+��}���A,v@4P�XE�G³����܅�N5�o@fk�B�"F*��j�5����V�uB��y#g�D�
%�+9Ě�8��%c_l�ޭ=j���<�SĬL��*)M��{j�'��O��)�i��Z��@�d��(vWk��u��Kq]5\�7<�$z.}?4��/��O�Bt��
m��ZQ>��Mv�fS5�k��󛄫1�����ZG��c�f�Q�\�nX/����	�]C����>�~�沶s�o�gn&���KI���U�B�^T��閳��OJ�z�F��s<ť����ׯ�C���xLqi�=V��nMV�ns�LO��?s+�U^���#�b����а�ɑ�j��\�׌� :}��{!b�G[���9٥������ӮpX�SJ	P�ˁe߈���/x���u����w�ܟ���v�˷�d�61�&s��C75S�|f�2%i�.��)J���B�W�FV��:0\����H�߁˛�)���Y��O�g{���*D��� ��n|2p98��&���[ܮ\������Z�Z.������E���g-U��_w@%�
"�i��ٔ�xc����A=��y~[^��Н�l��b��_��N�����{,�vG��{%��g�io�ҩXq�n���YK}+� q�-:��Y�����V��?o�܎�� L�J����L��҂+[�f��~��ʘ}�@L�ѓ,o��=�A��w��j�k��e��z*V�`	�1��J�ڐ��N�)N��_}1�"��4�P�z���r~1�c{P�*q�R����ݳ�Wwr���"��0F@��/ꙍf����_�/�~v�h�>��I`�m05^�Z��RE���u�2�W+�hD��Q���$���%�V�7��$��ܖ�NnI�o��@w�-�����"�E���׽A5@��}#��P�eP@`�	��X<��Wc>���*P�ߧ�ړj"CM;a��fa�JGwK&���E(0t��	�R�j���0@��cL���ux&aʷ���i�S���>�
K�(������OkVX�Vt��s�z�]]����V��"f��ޥǜE�MӮFh���䠶�o9��E�-ަ�1^�5B�r�E:�=����e����;�l�������^�� �	X�{���):T�}� �jGf��X7�p��``�X	ݰTͺ��"��7��(¼;ܼ�yr�<�^�p-�9���_T%�#QL�;��5Üѳ�?qe��j��fe͸��5#c�G%ټ�ȇ���zG!)r����W�|��'.���Z-տF�	��0}�z�Z'�ڨ�rA��vP�Vfv/�gLϪ�p�^�[=��-=���WShk���UU��v�e:����_g7Sj�r���@ݚ��{K�p�m���s�Ϫw۲1���NNǃfY�6�=s�kͺy����;i{�"^B�ϖW��nk��@�Z��F�4��I*�r��D'6�����4/�\�C{mf$>Њ~ý[!9/�糣��ΣqY���ٖ��@n+:��}�[(Beٌ��wW��z��Sv�67<a{����-:p� ~�%c�=�������1���:�eѶ岲���_w+�ɼc:89$�\C"1WӐ��Ep�
��Z�$}���&+��|�>�_�υ���CV�'����RK�rTU��w�3��|
���}�;p��c�McǍ�o$N�|ga���Y/�1�<q�G��.j�����Wt�ɔr�#2w�ι�R��5|��,��Wp�Ǒb��:5�;�����^6�4�+�e�R�%7)��։�.�M�����
�;݃��K&{�Ӑ��H�yp��Cp��yI��/Q����%��Ɠ���v(佖�����^�R�T�?���uCo�.��o'R����7+E��,�'$��CG�Jy���Qv�Gjp�����Ej�[�d8غ�tPm���R^�o�ǌ�ȗ�v���ge=��n��L|���w�*�W���|N��W`�p�✾Z�^�f_;'$�G�9FX�M̷a�.� ���nj�Q�}M��#x�{i������vf�P�Y4�]��A�]�тl��ۛ(��v�g�Htl��,(^޽���.v��U�a7ѱ9�h�]�9B�{6�J��q����4�c�g{��2�/�l�)[���g�I�
O�9k��J�XSVI��.��-�Ә��J2�Wkʋi-��NNr @���^�D���]�3&+���!L{�(�j���s��'�u��96c�cfF���;�5[�#Uu�|T3h����a·O`J#]�ya·��lK6.W={A:�e�T�g��*�0N.��r���܆���x�}���~�r�V7�eji�Y�����m�[A�@�>MYLT�1����c~w[�G�GhUt$ڕ�e��p�향N��Okg�^Q*'sh 5R!�F>��������!f��M�Z.
J�M\�;p:6Z�um�];e�$�é���	2p�����\��Gw��\.k���W�{����������r��mŒ��n�N��Ekd�_/��y^�,���/���1��]\�}v��.��.�`]�B����S73�'����M�7���xt�[�d��[qxhv����bpWz;�F�
�AۭqgD��,6�b�&7� y��D�jK|_+|B}�]�&�n���R��O�~��ta���D����f�0��?gh��v]����A��xUPw����k��F'`�{G�5�G���ekn��fi�&:�=�o0��(��j���r�q ����#poQ�d�X�t�����T:]��Jm�%�v&fH
.w�qx*U�*�:D�����l>�p�8���:�a�Dc�}c�Nvz��W��K��T7����E�����;��Y� Y�X�o.�*?��ȑ���$ھ��o�dK��t��hѨVLP�;�Ħ�Ǒd���x[#b۫#��%Ե�\��ح��VN�1�+U��j�4��o��GZ����m��� �j<��l���R`�v�c�ڕ}3m�6|T2�<"�p��SfIb��W{��L)��%H��\�ϴN����y��Z���eu��òv��믍��,�� � � {�A�6M��`ɣ�2�4 a�&!$���,�0Г1���H�&�H�%4B0���hFD# �D� ��#.����Nvjb�I�1!��%���J$�E3F,M�F�@�IE.� �%s�(�hf��0SK��&$e���tMH!18��ws	���&�B���4�s����#4i�`���w]N�q4�C����d�B����dQ�$�$�Rnn�%Κ�P��w]N�%7u��Q��K�hē���S�a�٣!) �C1I�\���"0�f"$�������&` >��䱴�ɼ���No�<�j��m2�N77s���z����/���m���kh6��+z8�->�t�Gv<��Z�������yWyw�@�3�ۍ���G���:IU|�/O	�J�to�w^&�R;td��{��n^�w
捞�;�����|�I�n���T�p>�Rf=`�@R3kW��v-�g����9�ȓ��t"��q�� �������Nh!5�3� «����X�\�랽��M�@p=>�U�	���n��S��C��	�P�z�i�Wʑ<&��.�U(�+*s��p�S���.!k�0Wi��>&F���As!����+��R\̦��r�)b)N��V<�ٙX0��&��\�+��ኌ)��ݩ	11��K�o���cq�]�^�<��l
�t�D�۷=RDc)�^Q���l�WZ�<~���%�j�
{�E����L�Ч��P5�;�r�Pd|�=����❠��>�&��h�@m״Hp\�\$��_м�3VX����I3�L���G�RnF�h>�ps2��������+"=��ҽ�A�̯R~5	:��T��C���o�Q#-u p�N���OF���n��U�H۵/`j���m�c=���^Cz�k�	�0���J��0�V�4�e9^��K {�p!k-J��,yϢy]B:����S�駸��Q��@ѻ���8vXK
7�������Px�ۻ��������lm���� �ⷻ��(��k�8��&�Z�%g$� X<�m������qz��8���ھ��ڔ�D��}ٯ��H4jwc8r��C�Ҍ�R���'h��eֳ>�N�+#k�	|�k�ǭ�J��U��L?9�:`�+u��P8x/+!�e�=�9����y'\������q�{g.;�<��{�����ݑ�h
�~�(�|#K�P��F���T4�f�G��LY���x2<�a��t��u�ÿ}++B�`��t��g�0�YJ�5gWª�U-{x��g�*�-zb�+��{��VA��'Z��'NXξ�U%�lsa�ENø�!�M��3�0t}?�������w�Cp�0���@�qm�n���0�������wC�V@���DZɈ%�ǺAg,!�5���g�;���f.��5b���w�#��_�q��iR���''˛>3��Z�2���R�c.Ch�ʾ���Q��n-�=!EC׻
���E"�%_B4�)�O��$wh@h_�ȶ{+<<�=�ql�̈��V�.s��̅%O�����ǐ��y�.r5��
3k��@[��>�2�/8СRd�/�����}2-��v��B���&�r�)Ψ�r���B���_y��9Φ[�ﶓ��o��n�F����!{�jd��}}�9��V*E�럪u���fXq?X�1�D)�tt=����ǆ1:��Zy�t�v,\����3�t�[5E@�,_7,gbK�1�#�h?v. )��}%+1{��:�F�2��X�:*5ee�usco�� U�����)�t�ꩡ�9���-�Ix)�9@�|��V��04��ߚ(��1Qw�g��~�ໞ=�y�o�E�~ZW*�o�XP�� M[�\6���j�~k��r�p
�{n�]so΄�k�*��f�yB2Ie�4�Z�p��8/�� ���
��/�x���o;��1��]�n\T��)�+��c4��u��k'F=���6O`?1(����#ݹ��	M�L�Fh�>~� D� ����[�"�l�mOC������r  �*C�Zy
S^z��%'��Gy���m]z�x$����dZ�4�V��(Gl�v#]`���w�y����{ ��`m�`��d�{#�LA�$B㚨1�/zz��<��6F���4�t�g����w[�̨���*����M+ܼ�xp��I�J-ԍ�4�c���'�]YF�DѾj��-.c![�qt�3XƳ�����
�(����{e�zꋍ��+H�?�6LM!�$�'F�ȁ�ũ&_(�w#O:w=扃%�z���J �i;� \�;JW����_}���s�YGV�6�A X�ՠ�ZSS1��%_)0^�;H��B[�5c��h��Z�O.�����8��m�]D��Z�k��}��<)U�w��N�~0)�����6S�>��!��m.�A5_����夃���g� �A�i �(r���'�o���ؘ���#�����9�X�6���J���:g'qHH���R��;�W.��س����� m}y�^Q�mq�vÓI��^@u��.�wl�U����u����qx�bw��0i���x<�(�>5�q�g+7�����yw�fw����,$��{콿j��Q_=�89j����m���;Z�/�ٗ	'UF���p�dX+o�{m��#��o�>�1dU�
#_���V;(׬�>W�R���� �H��}��^�7TNEʻ�	� ��s\.�-P�n�Ռ�)9��}�U�B`v!��h�;F��Uߵ��k*�$8N����+v9�ntIss�뺓}��l��Tߋu�x���<��#�]x�-��f20g�Ý���ܺ�{���}݀Q�a�ަ���kv��8��6/J)M���̽�����X�0ꃇI�7���}V�S�}+q�V�NX���G��ٳ��P�X9)���������헛�}f�*�(�I��P�[lgʪ��B�c�g�h�ו���z��7a�e��W-SsUշ�Q<��v��NF.
:GP��j������%�C�TJ�!��.�g����7�&�/X[I<==���;���Z:h>	`�'�1�R���S`�%�F�l�+�o]me`�����%}L��j5J,�V�]Q^�B�:K^�������t�����sS��dxʧ��ԫ����O{dsϖ���4��bKJd�ش��
�?�Z7ɟx�Ý�((��{7�x��D�$?�\��Ḗ�c!f<�	�P��>�
��9w�mP{��5�{pwe�>����%=딥.�Z'�]=>�7D{M�*�Bi���� 2�5�ji-ZTm�\�c't��MDbݿ��IM�H���`)�#<��q�\�����m��;��J�Q&Ʉ�PH��V@BָݕؤZi�[m�h�5��7�o��B���>�āHw��ĭm�R#�>�k�x �p�4��x��u�Ӗ��_A�Lvһ[f�2����L��ٍ��}\^;�V�ohɯ)&<�c���t1̔ڥ�^⿛��G{���d�W3��Nnm��-=n�8j��VM���3y\�D6Y����R����0��Y��$��LQ�>�mۆC���y�>����3�P�j��GO�s1�*���b{���$Ek��X�����a%�TW���^����Kj�?�`)�� =
~�_G�]@�yfNع����??���@M�	���v�}^��T~�z,TMp��pT��1��9b�+*z�����Xj��@����{!I>�|�����{cE+�z��5"�Z�~cy:��T��?۞�bE��&�FQ^����c�'B�%b.� +�=Bn���D��DT��[��֢b;�uL�����#9g�LU�>�Uȹk��ա�^�)�q7 ��f"�Y��=�Β�*��l��`6���+q��>��Uw�+�$]��S��Df�hi�����qܫL{i�a��=�7������36	z��#��w,�=8{J�o����Z�ݥ�����>�svX����^�n�x���S�*a#��ལ]�Ayӿ��W:�8
5#���?B�$�zT'�J����9�j�d����eG,�B*#��<�3��@/no\Y�~�@���>c'�肎��(��(���w�rg��]��L�=����@��]�u���L�\^2��Z�[(��1�IpQW|���4�y��������ZIR�{�x�)�ͨ�
����tN�N�-:}�B�Ud�Sr�u+
u�%0
���}�}
�7��� �"��t}!�F���L�YQ;(n�S-9rz��#�!�/�凩�*V����f|� i�"	pwdFr���ΖywOr�T�Z�Q�wEɂ!A��q�V��DvwHW�3�J؅�$=(�s�1�q�Q��t��8���A����s��VY�c4ۿ��۸�&]}�$%_'|g�H������O�z�tq�w34���p���u����`y�
� �N���G4�/Hژ^XL�&�i�{y�޹�r6ە�Pf�E��-�SIUѸ��)�`x�FF`o����6�.K�[~^N}��f���q9-�<�Jƅ��DngL���������;���
u��I�J	���wN�K���y�V��0w<#E��ez
4�ճ�ml�n�溽�A
#��}�t�1I�)
a8-Y�b�}Q*p�����[܄06�T�X�S^�X�ӓ7Yc��j��e-u�aG��T;���x���M����X��Ǌ:�����g���e ��գ!�����hY���ܩ[zGړ�Ʌg/,[`�oH��^��׆�e5+I�{a��"b�k4�F��A�7zu��zAa�'2y��Z��!�p��s�������p%wz���,��':At�!��P���_}��UH�7e=�^�@���#��O c��#��u������uX�ik���$�2���k��7w�v��e�פ�� �~�Z��9b<�]h��׷�DcYt"�9 u�]睒�^�J.�f`�\����� �5H��8��/�ZF���0^�����M���{6q�feA�٤ $��k�F��N���5��/z���:.j�#K���9�bs�Df&����M���t[Ye�1ʀ݄Q��$b¨۰!!���?)[�����m�����鴚���wBk(+���ޑ�u�W*�B'6Ta0CI1�y=3UX�S�S�}�����2x��z$9i��ͳ�؝n�q���J~��-$Љ���w: �d`����*��&{^m�Tjj�f�Y��c�	��x���ȐAdF�i���R�����oz/bb�.�s�*�w&�?1{�0���ɨMւ��p�#��+���Z�[�Y��!�(���_#��9M{N3�������] �ys&��ɺZN�Cwp.�q��Wo��u#35�h%�l+�/n��-Yi@�4O�G�����s���#.y`�1{# �W{���0CՌ�{�e蓗7tIW����UWɍ�]���=ݏ�׽�B�`�붬F4��nK�-��m�R�>���@�����"3v�;��&T�����Ս��}G�3n����|��ɬ�����i�(<�N�.��.�@�[WC��i��D#�������j�j�A�֛7	pA�wXr�WQyl��%\6xoOe�}�J3]Ju�BZ�3�������J�Es���k�O�z�7�#�!� �`�}X�hyq։ZW}����Mg7?oUL���8�e�q�䰬�����n�m�F�*�z2.Df������̞����}�RO��bL���#3^o2�A���T��V�s�F׮,������ۢ���	����"��7SG2WT�ţ^\vH��7����,6�/��]�I��P����e��k�����UIݨ�z���*ȸ��r}�j�q��=�abԽS���u�o^ ��h�n�:��l�w�^+`�\��z�I4L�{)�Xh����k�|5���s�=����߳K���w��Y�ǃ���n��is����P�	�;��M��B`xo�u�
�Z����u���c9�����߅
!�L��>f��5�ܑ ��#�:�SY�U��S A��Z	��l�oO^�;z^"��P�"�u�MaJK�Y�8�MV$Sbu�����&s�7�'�M�ٷ�S����o}���W�����)�nC�������ۡ;r���!��azb/}�Ҷo�C�M��=��d�ş-�{���T<�䍺�7X���Ȑ#_] {#�ƶ~����@s�͢��~��?P�#� ;��])�S.kH�c�=�Mvھ��<r�
�y���^Y�Ǩȹ����-���L[W�F#�#��>Z��F��x��Vo8�۹q	��mT�,p����]��+�2�9����u8�7�w��ӟc�qb:|\��~�go�	�Q��r��/�1ެ��\}�/NL������g+[�)�G_K�u]ާ���xC���;Au����,q+A��z�fTA[�Ѽ�c*1A�~W�:��~N1��d��=ˣ�χv��H�w�ߗ��}�m�㖧o�qmgW�����gKS�Y�u�z]�U��4�K�������C�������
��E��Y�
6G�ݥ�Qu��4O���.���ʾ�{�B�W���� '�VH=g��D�0�1ګ�^�]������2��.L� ��j�� zjr���WV�_���A�A����4��o�m���7���3+�-��3rɊ�(V>�1��K��-��ȕ�֩6�^���d+���7�����`���3�LF�s3��w1 4�묹�dZ3��H�p��ޢ t*/��(��0K��+��<��"_]��}�7Y�'2�`��i�X��L�2��x�:c�M����J"�T}���M��t��v�k�caen�6in���-S�$#�oe�l8M�r�Ӯ]��ccY��wK��TT��]@���M��s���=mƇ�jr�ë����y|~��4m�b/X�S
n���Zk��J�p�su��i�'W�^�{Y{k+-��@�L�1]�?�ױ63�j�
�lQ���ĺ��0ЂH#��Jt��h�c7�P9�B�+�H����.ne &���[*�3ud61�.ur�rR�B���6.0���Y��q^��Q�]�71��M��5>c^����μ2Y�GxA��\q⊟zߵ3~�tE{Ck�5�X�������W(r��7{ȓ07��;��ي�h��TNp��`�`йО�IM��8���ew_+�6g+�Լ+�i�l���m�u�H@� ��杷��2�����޽9q��AʥZ`s�"U-������������B�F�{�ٴ�w]���Mْ�5I���N�i%�NF��x��`=nn_`����pӦ����h>�h�D�[n\�q�Lʶ!�;��XK ͥ�D#舭^h��a��=hMᕭ�9�Qm߲N���]�?/n��Z��6����O�h|���k&Iv��c�� �U�Ž6$7yժ�%���v�L]1u��ͭqֽl��PbZ$�,ɡ=����K���jzh7�qv>>u%�=ug�O$Z=0��d�-������+��o��&��Uu�
|]���A Zأ7��0]@�h9��-�wʲ֊<�OP��g/�3�ܖZ�<)��1�z��j�+#C�w�ͺ��X�`eЭ��)� ����4���~e�kK�)��y}؆������N�B�=iY}
�~����Ⱦ C�uP]�ys�H�lIu���2J)���Q�Nn6��W�v�C9O%�lvu\.?{V��r'$�M~4� ]3%��L�9��q��[��J�������3݋;���Ѣ:��컭��~�K1u�,'��vIn��4��VD)p�F=�2��[�A�!֧vf�[J��zA�������vŞ�K!%;��>�q�A��e>{E��,�\UǂJk �->�jY�t���T����X�����;Y�_u�or����N{�������H&RE32�RM�[�A�G:��1� RwtBHA�ƄE�CK"�tNq��WdY��M��먍r�$"	��Rd�E�cDX�f2B�Ή6f@ ��D�P�S��4A�"d&��%4`D��� (�0h�&R�d��0i4�	0	&JbJb$�h���"h�X�h2S@X(�6S$��dRd�A"�M��"H�,�	�!0�(eH��D�C&��f����H�D(a2"����@&c$a0��P�I#I�LRA��T`L�f$#I1HSI2REb1�*B&�#� A�%d�ۍގ�J�n3m[qA�q��}RX����n��80ǝ�����V�y-������Z��_(���4Zy��&���|> NKf37��DenG���O<�Ʋv���U�>U.v�T-���_���tl/^���x��R���9Son%������N�h���;޹�m��--vG��]P�%���:���
W���������aUE�E��d~#{T�Y�����m���Z�D=r�7����z���C�^�/8lDf젤3=�na�0�F{>�0��0w�k��ChwDg/t~���]#�z9Y�|�R�`������ڤǌ�K���g>=ۡ��[�,lE1���.޸w'	���­1��:�5HU�-�N����o��<0r��'oʕ[|z��rm@�gW�l��m�{�6栩f�H[B<~�w"q��<E�B������u���M�vˌp���m�F��qT���]�O{�{ӵ8\G=�,\Tg�+�IT��5��mǝ��G�\-\��~��2Dd�+��p8:�j�N�(:�d�jӂZ�����(Z�7d�f�����������!.�ulm-��GW����>���^�<�]`4ڡ9b��:O�;&^ĥ�.�8"���Br'��ѳi�����]��o7��!ҒT���ϳ>���ޝ:�����ST={Q;�^9�,�ͫT3:s_��Пg8�v7���}�4��W<7�)�3����`��#���77�ϑ��4k,�}�kOIׇ5���y�뼖�]L�K��l�ՙ��LN�NN�-P�NN��8M�9r/H�y,F��6~9V�o�q%�瓶�V�ׯ�;/3m)Z�TΞ�]�}���)){�C��3�&V�T�=�{ڌRGc&�9�u.�c����=�[��m��.'<�R�,�^L4�|����nm;���`U���*5`{�*&���oKO%�b�=�6��_���6�z�7�2|���!j�;��^�(�bo/�ɧZ�^����n�W��&��m���n|2�>�9�7B�uH��|���WE���\[賽�/mi^�^�U�i�kz{��=#~͏�� ���9(�2w!��^�͇�zݠ�/gu<n��Co�o!��b��w��FG�ܕ,:��#Z}�5��.�=���%�1�s���u��ʲ�{��J�lJ=��Է]���]����������۳�pw!B��a�L隷X���i�׋���}�Ei���8�n���o}�'���0�G!�|׾�uz{=,l����s��QW��}������V������yc��Ȩ.٥2Q�������[Fof�s`�}�[�\����Q�\�&�;�v�nN�Ս�J������Pp���x���%�ٹ�irʤ�;�f9���`2���:(߰5X���Xf'�<��qQ)[;b��o�+;�5r�4������b�'P*�lwûF��pN{b�> �VI�rn�s�mVr�yZ[�3%)��z�-����vܽ��s�s�wsY���{�3�5I����ʴ�Ŭ�8��*3V\��dF�[��@>�Y����w]���Lh��zv�L'��{W�?��ڵ����޽v�u�/��O7o^h�x��/���&{����M)���FDk^V�Wd�z2�;8`[�ٟ�o*\��z�㫜�[������w��/�|�r�,�YRǬȯq^z��K��K$�j��w/] �[ l��e���D�/8���y���f$r�B��d����#����љNKӗ&�����|�����y� ��qZ9~����>���Y�7[2MUr�m}��lpn���P9Α���Wk�����K�t��֡*[K�79B�Zz���Я}	�K��4=�uTI�%���֥���nVP��>���w��~��~��q��oK�σ�W����w���`H���L���@߷˪3����r��q�S���ڰG�o�e��6a^)��qΚ9�y1�{կ�n��{�������|���+������z�F�d�]�^@4{���(�3ث�����(ycS��Y`8�"��J�����O^��~�T7ڝ.�\�7
�Z�S��^ϼ�b�5B�#3�X��K���ܗ��H�c=�N�v�_{����^;��7{X���	��MCi�l��pBq1m[:�����=�����-���-�g�Jg~X�Kl_aع|(G��VHu�x�2/���;hjq�rj.b#֝H!ҖF����G�Ҷ%�n:��\�~:e\�z�l!�
���z%gM�-�)�wz ϵt+ɋ�&��mj�v޵*��l�HMs�Km����1�Xe�^Nmg].�ˏ_*g.�+��ԲE��-�CX��=LM��mo�����w���uZ��ws�Fi�b:x������G����c��ok&'��^e]mwx4[�g�A���9Z�=����w�����E@����v�V��};F��_�~O��ih���V[�����>�������}	�Dq]C5���������~kW��k�e��>7�"*-h�w�%7��x�w*�̤�ʡUr��+\[�����޴����l����_������������T��"j+�=;�TO׫[�m�DK׷G�_{�l�z���̨�2�E�7��'���R���sP�=�S���j�����6����+5_��V���̶�x�n�5�}z��r^��(�bO.#���|5�^kH���&#�9yy:��t�'<���ߵ����ҩ:��g�-�V׮%���fۣwm[m�܋�K��̈�c����4� �/; kVs�Q��S�Z��m�7R���ܠL��[��:�1Z�ܻ�g,�9ɓ���.� ��f\;��I�1RKv��}�}�*r��uq�׭�)�p�VV�Ɏ�R����+�pVsn��O��n	�z�{7H����%k�8�ygX|�L��2My����U_|!N�{�����B�s���le:�4T�_o�g��~��^y�)����ŭ�ZRPkre�Ϛi&^�p!P��f��,�ik릭����G�ؽKj3���j���)-s�����%:as�\�6�q��>]'L��[�	����7NyⴕM|�X�mǝ�8B��M&w�g{��Ԩ׷Ӗ@�_�'�۷���t�b�x�I��~�`:R�\t�k���+bJ+��o��B�gP�T'm]�􇠝W�Uqλ@����t�$=~�;H��N{�������y,&��������Y��;Xk�%���V�����Qr:�C�7��s/�S�~+�^�q�2q����)Ү��><��*�R'<���Z�E����ԨΗ�����N��m/r����k`}Ft��i���G\����xǫ��ꘇS�=�����O(�Y޲�����/�l���d+���~Uՠ��w����AM���i��Wtq��'/�l�������{����ȝ��{����J88룠t7�׉J��R��L�ݕN�r�҂�I���Y+^��4N�v��{��Rj����[Z�܌b[��ٌ�������ۋ�@��wՀh{`�ԗ��Ua{�Ej	��obe�UM��ur=Mm�g�ET��������+@�>���;��^�R�&�M8��`��Vhe5�2��/1�c}I�낱��{
Z�A�CJ�N�b� ���
��{P��N��i���5��g�iʄ����}�`��*9�,O6VG:9�߫��'=V��Fs-ۄm��
���W����:��<!��im�s|���C�w��t3�>��U����~o ?`�M�3.u�ٚ��}W9հ�ƈ�R�� �?��w!k��w����\�oC�L?����;�I�Q�v��R7�N)ȱ��H.`����Mb��2�䶦$�ֽ�I��R�ݘﻘ}Gl>(v�,��Iur�z�E�+s���OYw��g����1#������9틐�P��QY αw�K�pn�=�f�J����N��6�TeJLv�r�����	�}��W������ Yr���rAZ���x�.82�k'ٵ:�m`
WXS�ɗ�.n�7�g8����X�p��A�Y�����h�l`�._y�=�!7�۝�iF�-�nh^�T
mm���}���i4,���v�N]^߶V�'�[�}Cz�븧����Щ��hT�ב��?K�O}����kW�������g���.O9��븲r�T�eʈ�Ï�B���T�c��np�7ъ��jg\"�f�z�N�|7ю0-g�k�D���.��i�UPS��rh쟯F@��>y��5�ms}v����۠�����3<�o݋c�u���#�t��]�j�"�=��7%4�/}ܹ�n-�T�_���K׶Vjk%�V����:��;�cUT��fr�6��u�G��<�R��p�[g\�o:[y�]��7	��1�"�(m*�Y�iEM�8��Q%j�K�\k��/W=�o{}�V��Q�N�^���g�����g".\��y�Ց'W�+^)n�;]��q�?Wq�N���m�e@��c�F�pU8�;���8�'tA{�[�oh-���r��J_�
�������w7LP$F�+84A��)[��9�c�|6�B�Tb���X��4����i�S��ؙ51��KV3tX���>Wq�������z�}���V��y��Ƙ�3Ty�;�LV�=�jͩ�沄�C���[�����F��m/l�2<���T���Ur@!�vD���G����b����S������E�k��l�
�<���}\���#��J=�Mvڍ_�|��s��]��ǵ8�s�6���Ra����Y�qQ?5l֐�=,��/o���j�<\�<K��������k��?W�[O�a�F��N��)�{"���b)K{�^N�,�t���l<�^ͣ���w��H%��+md^�+;�(�[�����}��r���8��'��cSy��-$nw����%Vl�o��]�ߗ@����U��B~��]@�K�i$gT��B��,��c�]�;�[������[��y�=^̨���/�-I�7�{�_[���9z��KoK�����k'n�n�W ��{qߦ������E���צ�ΛT^�nTE6��^���i5���5υ[�ʹ��(7(���%yΦ��W\r�;�V�"'Cp] -�.�ØwA{Ԋ906���^�ՔD�?*L����w�@��ԯl�ŕgU�M�i�bs'���\	WY'i54
�dp�0y�[��L�w|�.f�*s:}��}A�>�gz<���m~�ꜮG�-^(N�6��낳Q{6���묹{�ɕ �q����z�K�%꿩J5�ˏ8k��y�LY��/Uc���)U$b�����/�L}�+��#S�Ԗ�瞒g�W,�[�w����O�w�3�i��ݡ��o٬ ����d0u���q�f�f�e�O��N҃Gi�i�f���'�5�i���:��}� �3�]ъr-��}w�T�M+�w���H讉c��Gq�.�mV��c.��?y����5�y�Z�����*�K\�&�6[�"a:bE��q7�i��sZ��`���\��q";�/j��״7vbaf�5�n<�v����<��!%�f')�/Q���ί})�dHr�:\���Ƥ��xCO�$��@���Kd��,�ig���NGl[�1> ������#����74���U�m����JzjnzT�,uZ0������k5��(Y��k��%R(���3!<��ff�k:��ߦ3�ԋt{#���O],����
l�/���9Ǝw�&l��T��V�5���@�S�sd
ͥz�#f��@�cڱ�r����sj�Ԗp�}�8<ͮ7��JFZ�+(q��\SD�3U�swy�Ъ�:y�,�];�������+Bi@�vz�m9m�*\�Ւ�:�������f�J���=iB��nJY%�見�J�"t��BfeF[7�7��C�`��:���i�ٷ���;T��E<�0���Ń�0]�A�HnP�H�cNi:��w}l�_��%��}��]mw����f�JrݯCz���(�6�<ڴi���-�#��&�FdT�]
�Nٹ*dV�,K;���[��j�`�f���7QksPRQ�#!�uT��Z��s�8K�0�3���$����;M"�\��[f�F"��Iչ��c�f�&��j�r�|ͥn�'�Ha��B�2���wH��@���:�N�QT�=���w3�;�M&�Js�pZ|;rV���0�y1�|�SGy���Z��0��{�[��T�[;��i���.�C��\rI��\uX��L����W�����EC�_V�/P ;��c���i���{��ib��i�hĞ��Fb���7	�Nݚ����Èœ+�u����|��`�d��B�*ql��3�G�<���.��c�afvlhؼ$�の�Ȝ��4��c�C�opv��|�m��<Y�8�1Q̔6H0�����,8�Pz����Sa���xb,y��{���Os�f2)�o����z�O������g����ܰ�P�O�Y1�愗TA.�!M�6�VGN��v2�ǇZ�(��z����c*d������Q{Y���W��5��no]���)��2'�0^ˋ��=[��O��m�g%����ck�nIq�ų榇lܫ�ėP5go�Z:5Y7���ͼKim%���¶�љ��v�����G.Oyd�8�ܡ���3X�_���]����u`���u7�{�Z�e�T��r�D���J��X��_Sqn�2jD(^�B�e�샿6��m^��>ʁ��8m�h�c{t��ŕk��ؚ�����8L�Q�>�L��}�eV񈘪
LW���ye_`[��egc��Ĵ�\�E��H�*��B՜:�2����`�+k�Txrnbn�c���*:M�U���զ��	o(�7bqkG\ƀ��)f��7n���uc�}K��[�+��g�(3d��`ۚ���3�<�<<[c"|V''�hh'�)u��u�\��RK��}�s�YO�{�����#�N�LΘ�!��S�'�_�e�{��u��KN��)��">�'�ʪ��#=�-��"��R�h#���{��� �0h�&l���)	Jh�Ғ�L	%3���Ř���"4�e��e!�&1IM32Q"� $���3&CE(�2fRC6řd4�0�&i$� ��E�� ���FdѢ!$
2i��I
!R"b) SR2�M0c ��Y$��0b�b5$$�#&Q	13Q���H��&E"f��c���6LE�DR$1ѲcQ	$��L���"L��ldM-	bF)��f"�$������ �%i�2fL��^�~���������W�����zX���u�鰗�{��V��]�IJ���{$x���`K�C�:�ݛ��t�=w��|�g�}���~���`�������]�9go���'�7q�2�����~nr�'v�<׌S�D����c��g�������zE��[T��/yZN�����d��~��dŹ:�����/fzz�P�>���Ns��r*N�yW�\��T�Ǜ��:�{�%�I�Ԩ{X�g�*&=�Y�Iz�<������g���\��u	�r`/nKڕ���
����18�D��e��G���z�垚9��Sk�y�e���0�7r&^��(ª@l^޿y�yⶼ2g+1���౽X��� {
�ZN�	��d�)D"�c])�ܷ��L׳)�XBn��ǣ=_<ӕ�t��x+��Ӱ:�d���K)�����xlp��b^�;��5Wc��f�����?wA����Q��2���gV���hq!�9���*�4��o���M�z������ի�I�����['<"l������[�/�j�=�i/)nR&*��ܽ�d"���K�� �U�mCl�{�������,<����piֽ��;�J	�2%)ѨQ�����]U�-r���ZQ��sl�a���n��������|go���;?W��yrm]:�L9�#}���:t�w��C5���㢭]E���Z��R_��o��6��O~��=m.X��,-���y��s���9}.�&�q�clC�";k���Iun]��ql����
m��̗�%�@lߎ��Z�\,p��?P~�W��k*����^��K���0.�g<�u�������a�5�iň������ᚷH��9������e�CD�KvE��^�(��Շ��g+K����fs������xC��}���S�ae\'C\��M�S|;Yl�ٻ�J�qu�EggP،�Ao=��]����[���ڂ�gv��t7Zn�T�H�:.@��𽨯��L�a�Y��d1�{���[_I��?yq�X�Mɴ8�ۃ�~ή�-{ۀ����^Ef���=-0��6��K׷f�&�.����W�]��$ ��T�"�ʵ�9�a��eX�l��s֦5D-�틣�+;��: �:T�W��6ɨ ����~�N<�8=ǩ�c�f�Q��&�g���qx�}qa��Z-(S��gm	);
�u��[�V^^�Q� ��S�ev
ɔ.#Eէ�k�W��9;��q�F��3���-_�wq���/Sw�u����_�<7�A�$�3�7�h\8쯤�R^��V$�z�^8^�׊�z{��uR]�'�m�b�;f)K��4z* '�H�Y��Kw~
����B��sX�}�ÕSD��VM}����h��dQ������r�����^��廰�Ny��
�c)���#�P�b�����=u��G:�YX1d��3Ԉ�����a�ٴ�v#���Ժ,b;� ��=ވ����1턄������ћ�R[S_jL;�e�8W	�D�l�iMN	�j~��j��Px�<9�~�m|�e)���ۜ�]�ﻸ>�v.C�C�ф�;lJ��KGu'V,w��M�f���/2�g�����^p�[�}�!�Z����dz�=-��y��Ρ��л�=A2�����33ϧWb�:4�А��l�W@�.��#:��{A��9ܘ�շ�Wu���6�I�Cmỵ�ހ�y�UҬ8�vL�&֋Ϟ���U ����B�;�+w�.eBk��'-�쇴3�o{�Z�9s\��Ŭ�D*q��\��:����HOI�8��gCS�n!�?>�-t��߆b�����X��f/=L��8ץ��s�p�S�C�|j������c���ꇎZ�C4�w[�M?1��L�V?��ޭ���-�)w�\'�Ʋv���Ds�-BaW�|o*w��k���J�Nʩp������D�z���ߔ�{pVjk'S�ޔ��v�����ai��߾�h�Z�o;;��U{��on%��гLx'��T*TNlX��NIT��m��?�5��.�;��wx�~�s�jr�Zr.g�[���8ED�����K���Vvw��L s|}ݸ'{;��{�3��p�y5B���fګ��x����6-L�p5���%=�g�f���5��ϛaMx��{q�M+`�k��z���Ge�������� T85Oi�''��
t5~�F1���wSz��
��C4�>����#.ɩ�F)�S+ۚ�>b�������~w����9�)�o,�̃�:3��f�%X�i� :�v�w$bl�r٬
�� ���#'PE�)K�x)�4U�!��H�]��cV*�tU�tڝ"L�3����eIG(^�	Ib�!���`!\��{N�j��ub���TT�g���Nc7J���oC_2�+�=f
Y������X�QEmM}�7j�J�IN�#Lg�+��M,�$���ٟ;�����@�5W�B�v�3�?]1�s��+�ͫ[lU�4L�֢֜�E-��6$u�NF�\�¦C�r>/r~6�~�%�g+]�V̔����w��)�a�� ^3���vp����ц�U����͏AqU,[c/w�k�N^�]/8+s�<~��H���w�K���եw�Ə/^n��q��M�WӬmc��ꗵ3��~���)�s�/G�վ�|��,��>��_����2 sZ�ֺ������V9���ws��&�q��d�M�v�j�������6~+`y\���T=Ϫ�r'�=~a�O��{�s/݉\��i�������^�J�FG�Q��y�d�Y���d�ʷ��ʝ��pʈ�ม��{;��)����M�6F���U���9Gj�d��T�s}�z5ա�M�6���í��`�N)d�N������WG�:�\�NQ栧�k��pAb���p��8z�z�{�n�����n\��8�+Vv�Ua�8����V�z��/Zyy�Yp�������K@R}��:}��BԷ���Rpۓ��j�E'��ע�a术����VzF��ZR#sl!l�����)�𼉁�M@ܚ�f�����5��ß��W+vʭ�n6�ݰ+��3�(�?���� �}u��kdf��r��`�Z��'�clص��w�"lkf�d��dv��Oge{2�s{�V�i?6#�������ήl��J
�S��:��=Sy�Kܚ�YR�}m� ���ǎ�Pp�%�.LJn/��v���mr�2{$�>[�n���K��`c@����饟n�������r�P}%`����mP����g*�a>���t~���d\����<j��CK�^}������y,/�����g�r�0w����U�����E�%�X���}��%�����Fa���WVM�f+P^t�89�&VZz)��5�����`��>����	������J�x����s�}8汾�kf����Px�tR4].&n��iuǺ_-�r�o��0���g�:�kv޵{�:�
�-�����2Rp	�ݸ�ێ�ԅs�����#��T:*|�V��k��?M��}�o��A��x>TX�%�XU�=�ۡ���7��x�g��4	ʰ��{�uz.�=��ѫ�c��V�����Z����K�����E��ʚ9�f�{ B��p��uv���+�"j+��N�}�D�����z^�o�f�k��+@�/]k�
Q�*�,�ҫ[귁j7sx�N*�ej�R��n�5�z����y��q�hvτ��=�P��x�`���)��1:��������߾��W����v�f�
�����ٙ�+s<���_k��4�$��ּ!-݀��At&�$q���Jȸ�p�Ȏ��H߳c� ����\}[�%�=��n'�ld�m'��T&�S�sP�J���?{%yߔ��WS�i���Pkr��l��iD�;��AC��N���e΀��	��q{���,����V��&G��w
��wĠp}�e��Q����Z��}�������G�[Q�U����M�ϫohv�H��%ѺB��1V��]&yp<��/�����/��FW�F�]]_=V����)���b��Ӧ$��eB�K���q/Fn�ImMjL;e�;������)��ɩy���[���C�������u��������5��5�n<���.���pK���]f�U�(W�x�U��G۞Hr�o�U#���9\�^��zkh��e9ՇHHo�{���5P����Jz�ˬ[��Ŝb�X�Cٌ�8׻�f����8��xC���9~]0v��Q79S�21�Ņ��E��I�N/P�	�l�q�S���s�?-^+���G�}jq�w���8�1t^V�~�]7��>3��T�OQ���x�~O�X�N���a�1�����������p��z��Ȧ��K׷�����e�;��������~v�m Vt�]�#Fl�Y�k�~��W���2%�_�6��<�FT���x��au@�>�ꯤ�R^��(�$�G�M=9�U���86奖#�MKR��U���;�=�w�c�s��v�gT�}0q��%_Q��h"BN1�^7��9����ӖA˝���"&��qV�Cf�B�=W�۾����.������|��un(�p`��,���!ɍ�g_VL��f����Ө��~�\{�r���{�R�P�ۢK�:���V:��U#����DI���k��3��uI_��t��?�N�^�]�7�y�p�\���yO׫�ඕ�7���¾�le|��RF��?��c�+ɠ�B��a�;�B�E�Ұއa���e�/\��|�W��I�6�R��i�|#м��W�j19��*�K\�ɽ�b���Ԇ<Q|�K��S�)Ӧr+����c�_�{n~Ve������7U#�YF�[ѪQ�����b��=��H�Le��譨�:���k7�#i }5��ۇ�i��Nr�����H7z���&i�����O��6󛘎�\�CT��<W���ǽ�qTw!v#�IZU&�ɧ��Y��:��Y=L�������9?z4�N��0���~�3(:C��.��VoE^�>)mD�_z��1^;�(�P��L�N$�T���7���qu�\*�I;�n��d����R�0�W��x5�̤5�7u�n�p۔y�P�*odU�RYo\�)��B�] ��(���:�=���1����.׮>�-�R��2�w�燎Z�%����u���OQ�w�E�NR~T߮	��3�����]�|�:��k���yB:2Dh��-hy��Rh�lt��[�3ט:eRݧ-g�ſcY;:�
ـ|�$������g ���}P]��$�\������O �m����Jͨ^�J��6b�����(����Ȯc�{{��#���ᴧ����9}ݼ���E���'a1f3L��-��{J*n��y��J�t�);ή׿v}x���=��������Q=�^��,
�V=b>=����_r�)n�6�������t���*�ƞ�A��Mwt��n����u���Ou
ĥc��2\�:X�%�0�ﳺ��6'cR[c �H1����0���64Lo�A��@��%��;�w\',#Nv4��鸂��^上`�8�4�|���D�*���׋�M{/;�=�.���rfFX�E@�|�wA�.k�f��Vq�ڕok6ɚ9�5��]�x�.|�ŨX�qa9u1��q�,��]��'e3z�S�|�;���\��$z ϰ\�N�"_J��h�C���.N��sy�8�}2��
b��=G�xu�5"��Kvk��]�0�{����ߴB/��-dO;/=���"�pǑŗ�4��%a��t����sUBr����p�K�{��­Iڰ���L���چ�&��>s+��j��:���rx�/zF*[(o&;d�1���l�!�aCi��F>�)�3I��F}��K�=�Y�q��RU�./~(�V���x�(OL(��%�T��>E@�]a��Ճ���I��^�+=6H���}��� wKO�Y�����f�X�C�.��Q���_|�[ĕ`�˸�0��[Ac��}��.�I
�H�������y��Qa\Y�L��<�'�X��p�ɑ���4�y�P�N���o6C��=0g���v�E�^~��
��jM�Cs淁�w6Ц%�$��2�Y�a�9ۇW6��G��U7O�q̚#7G���c�[��%ɜ4��L�	pjP&Qڼi��;-1i�â�yf��v��v�pv��W�,�X�8	�с�{�5�fm�JnU6IU�78ӢΉ0!Wg�u�y�k��4/��97^���U��!N��.�e�g5{�����m��T�ۧk܆Ea�E97���á�0.��7b'�P=���)�xjsV�kz��!��Lf'��I�k�h
�r����{"�{�^[|L���(IF;���ECet��Ndy��JF��I�/$��f�G>�Pq[|�����t����;�4c���j�漧�*��oEڳ�}ƆRu�JQ�j���Ɖ�Fw��0��ڟ2�s$��K��).�X�f�eG����oA�[�,J�����i]��.jV29ݶ{���tv��B�)��|�(/��m��?W]��L��ǭ��D��%a�hbQ{YgT�k��<����c4�IQ/n�8�U�q"��[4���*}�ch�쮲^�u�}R�D�Z��[8E,t.��>:NXO0q�������#6�F��u{κ�f��닆�݀&PV��p�[�`���u����`���	���	 ��O�o��1{F��r�9���f8F`�$����G4��Դ=;%��^�ˋi����Y��!�$w�i�e�{�cލ��r.b��\�]�Z�r	A��R�@�i������9@镝q�v�E�[��s9��fn���0�q.�J,r�582ʥ��m�6.�3����E�,��{9����Σ��N1םx����Ÿ�%���>=X!1��|�Uɂ���h�*�=v�RT�c�=0lu$�ۺ9^f'�_YK/�˺�8�7�]V�1�+�4R � �����,�1L��h"&"$0h��Y�0�)6J1E$HD�L#3Tl�2�i��d�
A,�i ��I$��Q�4b�b�jM%�F�f �"�
���$����`�Q55	��SHb2%	P"(��$ER!H@�a��	M�S4cE��$&L�hآH�aM$CMb*�P�2DA�,��Q!�!+D� m0h�%-2�%2�bѓd��` �{�9t��6E��i�!�c
�������f�ǮAwA�A���"1t��,�Z9��Z�,r]�#�*�ȸ9\������y�w�&׽���bF��h>3��dv�7)����揲5�Ji��Onoܼ6$��틗�++z�v˼������oX�z����-�/7����.g�]��u<���,+�{��/�f���Qi/��{�^8�����w��FU۶�����h]�*���r����9�����b>�m߶��Xq	뎗P�==*yg'�ta޻�Uݜ��\�k��`=�m/��s�M[��ض���at��
��[)�8��_����;=qpSoUg�f��ڽ�!�7&�9����^�-�l�h�W7i,Q�F�\��d��¢��[on%�Я}&�.�@�>h�fW�Ԛ[iν�&m�����%j�ԥ/��z/W=�{���;|+�c�m�\Ko�zr�
S�,�&�����3�Nрgu}�;]_}xUl�|M�d �� ��L����
�Ȱ͕��8���P뛎<�&��Hm�����M�r�9K`kt�{{��h��H�ӐHD���kp^����5��`7x��������i]�)k��MwZ2EtѸ�j�{�_C��|�δbK��q�!q����لiG�y@�]�f��;�><�}'W��ᢖ���xC�`���n�7�����S�SM�u�B=P��y=�ދ�1��n<��[v�53���&��(ycɱ��sEHZB�@��)^��L{��4�lJ�^�K��1�z5kW�oC��mq�'.Q.v#HZr�{@ƴꏼ��v�j���q-d���n�䶦�&�2�+��`�h��j���>�+G\�\�]�}��5��J�c�;���a\�w�u��x�h��Q*xo
�m��n�c��/'O�|��.{au��1[��������7B�r-_vÑ�)L����7{"+��+Jy/f����^�o�_5��U���+͸�x�}^}nZ�~��#1W�j���� g����d=����e{���dFp�����������u��g�O�x�-˾ۻށ�6���n�U�����h㊽�I��"��*�h��G)oE�.�d��,Ǻ�"�)H�Ӗz�+pž�&����=�R��x�5�:4�0��a��v-7c�6r�
��[�/�����P.�ޡ��.Mwk�@��LC���uբ�6^�E���1�~ڌk'|R�9�q�[[��h-�~�%����]]�2^�z��Ȋm�Ľ{+nZê���7c��Up|�u}8NG˲Y��X����7�FT��e*F63����/��Z�5�<vc�כ@�[;�� �G��Iz���:� �w�Y��=mG�NU��;�g_^m�]}��Vv~߳Ks����0�����Un�For��5��)�\jƷ#�3��T��8|��4)�԰�t���U�|�+��g�����	�[c*S��Y��>���Z��ش�k�q2�3��o�����l�����a�h<B�����ܝ�8���<��z)lp]����>��w19�7J���|���E˽���"j�ڀ^�3�D��i�ic�e{&�<�\����S�{"'��ͱg�%Ku2f�qU���.L-��f�E��Ӌ�(wc��2�5��@-�5�tm@y���7&���tN��d\~��:��DQчk�6�T*��=�����f��-t��������֌�fɚ�1��M�]�T�M��Td4��v������9�E�E�-�Bi7v�:�����A�_�2y��k�����6urܽ���Z\|�_�'Z���x���9ʇ�:�W���ovn9�����7��w����'3�t��R�T���r���w��_��`����?s-G$�s�ײַma�k"����|��39�w���L�Ѯ.c���3f)���5�LE��e�]Po7p�����]B��{3��j�y�7貖(�V�^�\�����ث9d��R½�	����Gd���E�������Y��zs�6��{ɚ���Kܲd��tϊ{"dƌ��
�4�͉Z�O8�R���N؛L7)��-?_�Vm|���8N?���ʫ�N��Rﷺ�dʪng��)f�yy�Yp����ecw�aT��(l�L���Y�[m5�4Ѹc4Hƪ$�wIa���ˈ׍nCў��r���y`�t=y��/=rg\��TǼ�f�cp`@	ğ�Z�����Dig���+=O�n����ԜÄs���쿻�h�d�jf��H(/��pC�0����μ:��N�~Y�+�Yӈ�rD�y`��*e�<�\"#����{�8�w'�ݫiڏ��<5�(׳��ď���^r���}/�L�m{�����"v�Ԉ�{��օ*`-1�:mOِvw��������5�{�SK0zl�T:���k�?`��C2��ZB߳�٩^̰�z2�&jY�Le׎�b��Z�d��=sM���p�1:b�ۚ��T�^rזҒ\���3�WJ�Nz�����t�ؓ_&���,��8��j٨�{:�Q�/M���Ӻ_#��i?��)��I��X�M6�z����q�/S�A{�@�n�� w���6қ�K~�/2�e#���g��8f��#���sc�2��ڙl]Lo�y,&z�e��iv���s��]�G_�v��W�2����1߾�-;����#�v����Z]����ͪ]W7iC!B�>I�V;�r�n	��72��s�z���o����7Zn�P/+��C��|��bc"U#�f�O�wng��>��D�x.��z�w��m���6��w����b9$ĩ�;1lY*ܮc ���	�z]�F����Ri��%$�n�*���%ŵ��
�f�.����1[]��p��b� ]Ok(�{ON�nԤB�e:�W.=]��@ͭ^r�!Վt��z*�ϼ�i{�C���}�b���;K]���M.�B;�Ձ*�p��^�Q�^�ܶߔ�z�MzXܗ����\x��u�N����#�z�)JW��ㆭ}�����(����%��˪}=�zӢU>�d��z���;�U��q���2*��Jb8=Ǻ&����;�^twg����4���Q�o�δ��7HSL�\s���C*\�U��OM����}w���{��O�ڶ}=ǾR��ٕ��_Л{pSJ��o�g��&�T:�4T��-� �X�3�n"ۃ��o8�p�WQ���|wf"��Wڵ��v͠��d'Nk�2��y��������5����	1���^��'9�UB[SZ��e�;���ܒ���c7%&�=�n�Z���|����f�}�c5㴕J�
Eǡ�s�{���� �p��wP���`6�!S��9Z}o�u0���B�Q�����K���.�-�2��6�Y��䫽��N-��%���V��*��1Z/X��#k(��}��ߜ��@��Ͷk׾ydwy��wFn���#=ݚS�T!�U�
3h��g\�u�w?m��}�y�8Z���b����ѱ WN����
S!�8+��7{ M���`ŉk����QJ��Ƒ~���N�ۙ~��q���;o�b[�k����Z\[��J�Yj���{-a/՜�m.�w��̝Dw��y�O�o��c�v����ȇ����{�5e�ݙ�ʉp����h�������!?m�.>�76U�Z����R�83G��|��s�*�d���/V�9�6�նL����bp���/�%�3��ű��=�7����ޱ���%�D�-������a�E/W�:�w��r�L��v������{�#��gJ�/hJH�1{8w���NIBi���z�~�5z���,/B�VPt*䶱�������|�8h8}Xw�KoU��(�<g+�T���Q�Ǥ�U��-�O:��b�&�dO3��Go-���SYpk��L#]1|��R�̣ؐ�k(uрV�~ՙ�&&*M��iX轸�p�p�rU���+,��{N'X�g#�?Ey���yVx߬��Vo62�-A�m�M��0n}ŧr|�Â�K�;�FO�?��l^�0�LVn8O|-�~uNu]��
���	�q8��<~����g��Q��p����	!9�6$W<��z��RHr�/W�:������e����׺y�o�ߪ��F��x���]�SDf`�ϣ�Y	���֑�O|9�㊗$��y2m[�U���7�����-�����.'�v�X��=n�sڨ��o@·��n�zi�ꬡ�ã�B�7���¥�8�/r4D�nR��_���S���=����k~^�9���C��T���s���K	��yS3����3�]�n�~��?GY��T��"5��}��9���74��{���0or����}�~s�S�	gz���v�Z���\�ym_�^��n�sf�����>�6��d5��3@��g�nu{]U��л��>��V�o��Z'��۶���*��4����sʽ-� ���?�v0	�ٻ�����I�9��q�̯�%��K��t����jb���vl#Yِ������E��O��t[i�Τ$�w+�%�ǥ�γ�ˈ���t'��%^]�{tN�z���S�Z�o�ix�y�~U�d�z�=��9��R�W�o�=�_���&�[���0�����6����
�^�:l��>�V
�e3��Us���W�⨙Z��R�&�=��q�i��nǬ���
j��6��:�����@�����7_����I�Ƽks�C�8�#��/�����mGy������k�k͚)n����cA��嚓q�7�ݭ�M���ǫ��f���}���^��\X���n�_URr��fìm~���ͤ�?`��y��ܑ�����a�G�J�˟�����Z>jn\�M�W�뚄އa��
�8�lWF�˝Q�]p2]+���S��Y��w�5�'��.�-��I�M�<lGτ��v�!sQ�A�gz9��֩;���ß	9�Y��R�x�'�6�z�'��}����)Fb_JbP�-&s���-[sR(��ޮB�K�gqG|�ΖNm����tMDl���v%������as���M�0L�y��T�V��*.�"a�	1Ʒ�o�b�)Oxs��K�;�XtL#Ggq��dr]�:�P�rmvlgo�����Ox�����M����+��ګ���K��y!����#����+�^ �7��k¼����!=�s����)9Y��M�ꛟj�%?�~/�}콶6]	J�`ܯ]<�����y�0��ު�+#�s��}��g:� ��?!����1����2/�vL���Օ�ܫk���ܮ;>�\@ϥ�O��-��<_�_�OrZ�znA 6Wד�<��0�t�2�z�W�1b�Q��ã�d5>�G�����}}�O]F{{�Y��=�G,�)PoO�|h����:F�<|/�zn�C*�49_��\+�[;�ԇ ����c���N=o���T��=gėPf9�ʮ2����	ө5���dG�'��{���=;+�0327eH�������<vD�Fc`OǕC�[2J����+�"r�ĺ�A�Vo(��������Zm�T�\>���6}%��@	�}'@��
�t�d^�i�W�.v�h��d�މ�y�qo��O�x��u���f��Aヂ:�~��o�;#��W�W;���iFC�b�����׽]�kcx���l����i.�X���-� �Œ�эpa����C�LΔa����Xq���-����1�Cě�������֠�&�iP���{ζo���Y�.���6_������^{ݏh���+�ogD�/��"�U^#�>����F���H�W�z[k�w|H��	��,����."A]+r�6���9�hM"�/'e�WR�h�*ũ�<���=D&zTﻶ�t���Ȑ��n��<��4�"�ݕ�W|���le.{Q���nf��WW�T��{�p�`�j�}"-xH�c�C(�cD�{��z��h]�Cns�S��]�'(f��@�d]��noΚ��-dG�ڱwH��}����n�
M��|���0���t�Mqjwm!m�팂���;��Uhڀ�>�{��Μ�ΰS�2� x�]wwׯ$SI�o#��2�j��o4tf� S��!�4���7�m �5�Id$wq���Ls�'�����5��?7\���/v?{w�jQKc�C�m�c������'��6�؂�ƙ�xl�Mh��+�z���"��Ŷo��U�Z^��D����9�L�v�q.�I;%��`��3,�5��0g��9�G��Vp}�.�;}.�	~*��&�s��PF�R�i�*�t��Tk9�!��ȕ8:I@پ0X�o�\Cp}�����^tBLb�#y��8�^:Մ�f��wA_t��u&q�.6wlGLҋ�J��`K��6(A���}��'����b����"��ޜot<U�2gM���7/#��y���\�.��� �'�;2�,���y��O����4����0�Z%�;&��\=�ho٫/�i'���/�N��<�v"��n�u���O�^b�Kc���彳��EL:K��f�Wi����u3�%7��J��$��j�v��+܂�Re�TɕgX�ݪkw��B�j�����Ct�yɃ�l&�|��ƶՍ�����'1�=� ����:�6���cWS�S�N0��3*�=�	`�G����њ��0aWC�p&{�ўQ��,�#BKؓ�Y��t���Y2���zZvwD�T�u��廬!��2q0x��޻7_ud�Q���wm���z:���4�=!�j�'�W��ma�+���x@��x����j�!��σR�Β�$m̩F/i�wVk5�Q�/]�ٵ08ɣۆv�'B������]��ps���F[��SS��P*%z=ؕ*o{BP�jT�^���T��{�"�T���=��i�2�#*΀��Vo �� �;�oV�Srv���_u�|(��|.���ʸg6)h�c���]ҡVq2�/h���ܫ�f�&X���{���:���'���L�5�����LH���t�t:�Aj�"F���ʹv��.�~��0�Ǖ:�&f�B���n���ۤ���)��;����>�H'�$�H"MœPF*J1j(����@��K�~w#s��#S1� �s[���Q�Q�̱��gu��H�F����%�X��h�2Q�A��Rh���-c�e%$I�l�渑!F�,ZBJ*i��4�Y5˚�(�h1���"�F4C"���cdA �(؄Ě5���ܨ�wEE���	�`��F�BNv��F��i,h�wZ��.��"�A�"��3˾�^{����KfMh'e��龓��j�dpn�cqnq+�K���{­~Z!����U�{�eva�w-��p0�G#���wB~ԫaB���¿@)��[Z;>��ٌ���l�N����\_]��7�!����/2�k:�h0} �ޚNW@�z�7	���|{��9�8�yƣ�_TU��IW=~ˮ������n�Q�2F��&�k�t}��5q�c��Hc~m]п�7\Og�g��Gs�Y"�H��\s�
< �w�P2m� 5B]��������'4�i�|pwtԬ���kӞp��v��w�נi�懯��˃#}6�6�*�b-Q�>��k�f.j_�S][e�Zh�� �k�{��G���󮘝ϟ]�]C&n���A�� z|�Wn��E.UR�{��(�d�����e��Re���}��{��J��x+�Nq�8�H>�\D���q���r}y~͵��s4��צ6S59��Mײ�T�@/�̯�Mq�﷯|b�ݞ��a�w�C6M��8{ݸ�݁�N�a�	�<."�k�������N�"�r쁎���OM֏�{b#���?_�&��>�gk��I�����%-3��y�uR2�oު��=������#�s���:���WF��4xc�]i3u���Ov�A	�:w�A>�}xn�H�r�=���ET�"<��pq97��Sz6Wu��
�Vk;�N�ٺ��Mɜ�{|��cogq<Ć,�/9��7L���	'Nv<<��O��B�6y�r��^�.!���Yr�(Ԗ�A�P�(�#Qp7��z=��f8�c��/�z����ˤq]���uθnK���Ϥ�r�%W�:��P��nc:�G\�����i�jk�����i��>����^��Y��+���8�3�Y�������> z�%��ݷBs��u�b�e�M78'b[�<3�����oAk(y��:�Urc���ٯs�I���{��T��������G�55� ����G��v�GNm��}KI����3�2��ʇ��}R�4�*���讞�:m*� h�+�ED���5�F-�Z|�=(��XIً�U~�Q�Mxi�HΑD�>�:ǑE��������6��惑�R�T�q��NN��������S�@���pݐx
��]�2���j�ܑ��P:^ׁƽ��3�8�z��=���t9�w;(�>�\,��wtn�q4n;��އ23ѽC��V�9炍6:��i����)Z}��dw����km0����n��P���>�C�8ۇ�C׽C��	O��v�fE�6��Hѕ����V��7ː��t��'�
����fZ���_/z����5�B�4�<��Է����#kbq7�XQ�����.*rg&;���7�
��ū�x&leP@��9�j��n�f�D�N���0�2 �G�g��ۣ����S9>8�MZ���B����}_LkL��4�}.��<�2<���Ͻ�\egm�i������;��Z����jOV����f�����7�9�>��L��Lj�w��Cu˧т�� ��w�k�!v�̖�8;��R]�zq,�
�J{#�鹖�	]䶇��&15dv�<|�p������c���&r�i��1�O��աd.���s�)E���4���gj�U#qE��nn=2���U�{��W|`>�;@s�\f\�GҺ�=лq��:�2-I%t=�U�����:7(�f�ul���x����N�=E|�{���qې]y{+M3�Z�
�	���_z���h��puJ�%�;惛������ǳ��,��s��ϋ�q���l���e{J����Џ�:�`�$W��f�e��xH�o��vO3�9Q�܊��}}�0r�6��hr�H�E��F��Qf���1�&t��l~5{�q7��G=��.���2�C�>'��z;�&���]v��GuQ鸆@�$i��u4�=[k���~�/ۄ�x�`��pìc��x�o��x.�$Fo�������E1�:%�Ϝ��'ϲ�
wF��ky\׬����A����k�</C�x��^�'�=�w2�1-X���N�J�}�5�ET��){ʔ�oڑړj�!���9���mx}��/���[��,\*����}HR�_ �
>�����iPУۇ�:�-3���/�"x�ӜOg��O���p�+��)��
��ƣ��<��Ϲ�uҨ�A��F5&�#Z�9�y�!���Ʀ��}={>��[�,����X�Xy�(�*7�R]{�c-��˟G��8��U�67}U&��Pu7��Q��i9���W��L�@^K��r�J��P=����K`�����w�4Q��ۿ�[��&#����oI��|<g��X����k�졛�R�*ϵPM���n}����&��)͞��Ꭓ��z�m�@]@���U]��wW�7��J����z�G�δ;�=�����L���8�n�v1��V�"z��{K�8��x�iq%�k9��ۑ��q�ʝ�N�ɜz.g�h�,��=�]7�\�����!��`-�p+WZ�>u��W���w���(�=�Eh_&�n�=�򩎾��1#Ԗ? ���T5ƅL�e��߽49_�.�
�Lu���O�O�b֦4�O�;7��I�&Cu���Q'��l��hׅ����&�z�B�L(��mNwP���9�-�|�&TI���GV1:Ys{~����pJ]ӵ�q7h�j9΁F��Oh۞޲e��6�:�Wܮt�����$�R����P�]�YAs��-�E���>ίP8c��n���+~3T��S)���ޱ]Rx���ޫ6�#ܞ=��S�uq܃��~�[Ԡ܋�6���ZOd���2ˆQ%��<����L��ӹ�،����������̭��9]�=�wN��⾎���|; l�K�r NjN�0����z(�����5�r�vz��q7��8\���}}�Fw][5q�TpB.�d�ƶ��?c蚼���ܕbo:��b��Q�kCȗ�ٌ��6�>=;�o��p}q�wƅ˪,޼�j^/yj���kwL�G�p+zh\WN��|_bې�5|ʏzq��8�d
��
X��T]����8�b�+���q�$r��Љ���7Z���X�%r��Wt.u����z$Uz/9mGa��{��ͯI3��Pd��
�do]zV���`YR'��ڹ]����L=�	�׻qߕv�qs�g��t�}|�Y��<.��E(�G�PN,�|'�ں/Ǵ�^"��?m{�w
�~���06k����=�C}v�ސ:���'r!��ۈ]C&n�ޠ
5���z|:2��B��Wd^�7wh跁�w�=88�̕�|�lM��w�(N��Z��X5���j:�ԖK��&:#:���	�4�qƯ��jӛY�� 39����h^Y�)�3nN�sg[��gS�Z�.�^��V�Y8��|�o�9qs6>f��zMlti���]#o���+89 �G��쭨{�k��7�K�G������y{_��~�/e��M�bS��N)?�A�zxv�)�r<��㉁u��Ry ��2���^�z��=��P7&����t��A������;�c���.+&�n)��,F'hp��d3�Ӿ��m�EHOZ�8��UI=b��C���HвR�gj��H�S���P�<] �fY�j�n��$���\�W/l�9Al����:��o���˔IF��R�du	Q�T%p;ɬ��TI�7��ٕ�ޝ�%��!��UX�C/�ݷ�r+�pY/փ���.���S:��P�r:��r�+��q��G��&?T���ȷ5�n<�����^���,�����=^�����,�N�{pLA�_~�m��ȕ̑K
�}�b�y��^[�0o������ey��:��C������}�9�xC ���l<�� ���k`6�^���7�ǟN���݆z�o�]�>�֪f%t.�j(钏|��ʢ��J�R_�80կ\�|��D�̘��2�G���9�7��6��Mm�F��W�J�;8آw���2R�]l�s��w!���J����sɭ�I�������^Wq\�E\���P:���99ȍ�q������5�n���z�7no<�{x��}U��d6�.vʷ2�`�����QÝ�T3�����}qE���FIh�#H{=G(�>��C�ۃ�-)������W}ܯ��wR��5�t9�=���VuL_ЦO)�;6���839�ݙ��:�`�KA<��g||�a�Wtmz_G��t9����E.�NE	��0�LL���v-oAp�՟}8�L�q��t;w�8�?D�=ޖ'_T��oP�bk4ک~��籘�-��.�5t8g!z՝��u�C��w���\�<�F��t�R�j:�%f���o;Ѫ*��^��m^�
M��hM��MϱG&U��1u�7�=Z	� ]9�6v	��$���KFn9��LW����>�0T2�����k�C� sJ��NNK��2o����N��U�Z�>� �e!���uۯIcI� ����=ru垙j��p/ǣJ
������9�:���>���.�b��(R$��2®��Z���}�*���7��|�.�B���P1:,����++��hs���ei�RG��}�U�ϧ!^��mۀ��~���HE������H����g���=[�q�����݈� r&���m�UM�)|�h��l�N�2H�-'J������M�,��ی	�9�Rxf�|������N� ʨ*B:�.�X��ݔ�]mk��g^�32oȬ�
0�)����盛����4������7���dv�gl{�{/kz��r�=�\�>R��43�;�:mI�t"EA�l�L��-��q-��dB�W2��*��N�N�+�M͞(�wR�.���>�Ł=���$�#|��C����B��5b�����n���Q5��C�r�;�Ԇ���G�+�؛���C sD�2[�e����=*_V��9���Ί��3�}m����=����6���\uU�uU���	'<jnC�52=��}�u�}�+�������Zj�&���ϧ�<rNq=�`������E��r��<�����)7`q�6�T�u�NW�_��׷�C��Wtb�M��6�z�92�y��"(?G��=鸝��ꍅ���$�t��G��8�j�񸄺���Pu>TH�D��_P�J���9��%O��ĵ@g��9�*�P;m�Eڃּ��Od;��;�f{�<s.��-Í;"�<=΃3y�a��C顫�.��z�>�����z��er7��`Ŀ*6}�|��鶒��WQ�Nq�ٲ�D	���vfc�>��n�C��,Kٽޯ7�2�^�R�v��))�GZ�%�9`7�x�'5��p����qz��Vo��}���QS�M�gu>�f�^�y%Ϣ	�mEv�/x٬W��k+���֯�GUWi-���z������}��g:�t�}3�G���|sfU���t r��=�Q97٧���:n<\MTs�;����}�܍���T�o�>>]�3T�,���d���_�'z�Hށ2ø��>]!��x:��������v\n���z�8��_S�yW�w�+���������3���S<�Ӑʸ�MW�� ��1�»������꺟'�Tyw��SD�|z��Z�\r�$�3�T��L�n*��t�Ci���F����ˣ.�Gg���7����%���}R��2�,����2ٿ�e���Y��R�t��w���KZIރ���N}�#��G��zo��G�]�쁳�.܀��:�n�]����7α疩U��%C[�u��&�[��f����;q��G�j㺨6��_�����@b�Z��hp�3���K� �8�t5��1�9�ܘ^�iW{��UW����Gi�O"����p�*�7n��9���Nw���܇i����g��l�.���a���õp����ވ�q�F�z���ʏ�m]���W�nh|����x������d�Y����Y��yڊ��{�\���ՒLGdw�h�܅�����𷺦д�xݕ8��tQX�����,�o�fOD��}��Tңjd�PdEƽ��tZ����c��%r��� |����O��s�ĉǘ:%�io��a/�Pd��
�g}u�T5B^�r`_��-�Wy9�0�I���>�����X�;N���ή������_�����ˁ_.�3*�=��G��[O&W�:**���	���,�"�}�uڝ�/z@�7�(O���ۅ�2f�7��|rx)�n�s3}*���Z;��)��Ω~'��{�G����*��1��E.9������*����5Ƭ{"}�M�fG���z�tL�U���u����O�������c>UI��׬�3��a��0a6���cgמ�U�#�x��_��\s�'t�~�X�ɯd[�`N'h��\	���:Ty8ˬ�I��7vQ��s���n�~�{���ȋ8JVfva�EuR2�o���f�;++�誜��:\�}\9OR5|�օ����,��IF�$�k�*���w���u��̠0��>�\w���q��b��!���S�θ,��AƜ��!��S:�7������U��A,{�R�����^P̹�4*SOu�\I�'�)/9�7��{[�����qhZ�<�l2BT���=i�x-�J���R�j*����ծc�nư��ͫX��,<��0v�>A��m�X�W�E9ѷ[�K�-��	�/1<�o�-%zK�v�a�眾\����MD�Z�R��<��8��I�FP�+2�u�GV'�%��`�a����g{��OSMvEw��77���/��Bd�Ӄu�y}��fX ���7׎,:��`��cq��ՔL�8���iֆg��
�?;t�΢���%]Σf�+����2�YX��0,O��W����9�)��6]��5�V��Qp΂�3*w��dtl�][�R��]�l:��ۛR�L�WR����1U�TXY�e�s% ���a�! ����i{YI=�GB��:XW�Z<[�49�K9n��|:�a]�Z[��^mh�G:�OC;P�&�Z#\P}b�ީ�q׊:��g+~F�!d+)���d����J�wwn�"O�vyI�5���!P�˓��X�F��/k�̚:� �Ϋ�N�0��A, ��u\����2.��Qt�t-�p�E�g�޸t���ꬽ�U� �[��o|�w��<����#�/{U ���{rl��ĺ|a�9���.pYy���\+�*��F�6 	��-�c�^�RM���,�up�=��JD"2��&���q�.�~ۊdK_�o;R8A��r��qVo";��R|�J{����Jj������ڨ���I�Ņ��_.M�
K��D�m޼/��A���O.�s��`^�8i�U-*��mL�+s��t��f�B76��h\�A[�j�u>���&��il'��णN����G�Ul�ta�[�\�ZZe�+J=瓕�H��r�x�#/w�mX����ya�:�+)�[���t�o�K�Þ`�m[�K�l��-�j�s����D�QTM��W\�x;�z�u^ ��I�/Y�3"��fufT�xy_g�w�d5U<o.	坄��nɀ=��,'Q�}v3K@X���u����@�\���W���e*j�7�,*�f�U�|6�9-\o�X���:� ��"��#ez9Yj"l,z�pY�[^u��fWP��+�\��u%�;P��c��+F>�2�`��u�k!m�����o����o�I�%�uܓ0u�ھ_e7�Ѱ��sV��F]ftt�Pan�Ǔ:�t��v0wE:�pgvKʵ�8�1�뛘�S��Co0=�׮;O��pc�\a�W�B��iW��|��_N�!q����d)��V12���g�/aS7QTq�3R[����(Lc��^.Tx]Ô����4�w��˧��wX�m�=����SW��0��L��3_b2W�^���3��n�D�j�X����k��Cx������i��ơ��U�&�6t�Jg��{z$��ݻU�����4�H���
�3G.�&�ː��]w�˦Ĕm�*.���.�X�wj���r��6LjM]݌j6
�WwcsW#�˅F���uԗ(�-��̪�v���A�4YwQ��h�W9���mw\\��;�Q������'v�ȋ\�s�ܮ���G4EAd�mҮ��\��W(�E���jM���6�E;���2(��Gwkwv�J.E��خp،�t�\�QÕ�b��u��k���ͱwuF-F��]\��;����-�/�E�?|O�r�h��BwD=:-�`n���ٳ�^�i�Ü�	P��镙���3�:z�hWS;A''��Ɇ�ZxRa�f�K��n-����p���Ir�ط4���n��x�/���%���z:s�/�τ�/yЙ�fk�sX���p�d�j��/�O�"ۯ	���������{�'Ѧ�B��&#�+���NV�;�
	�{�J�4�ck^�=��Ȏ��csѯ�Y�����8Ft��]���Wn�%�m������y�j��)x���gO������Fz2s��L����ɾ�}Y�q.��o�d���#L�^�Q�/O�s�ML�����[w��A�Ό�ϸ�m�+�7��=�x��� ����Ω�I�;�ٰ߰���bY�����m�����r��5/9��wL�߹��h�wP��F{z�K�S���e���VF]��ûk9�Q�LkL���\*�=/Ƽ�.B]v�=螣�T	�|��z:@Z�v[�4�	��8:5�%T��@�g�&<�5='AƟHwUg�l��/>��s-����^9�:5U�=�Q^�����ڼ����{d�hu}7>�S��t�&>��WC��t�!ъ�����xE�Ҩ):����&�*�6����`�4��>>q�8\9�+��m�`m1�*�R�f�������;@�;�\�gM�2l�ǋ�`m��+�eu'3��t�ܫ6��������C�>��5.�J�t�N��k˂Q�55^�˟,Iiɛ��9Z�����S�Y,��u%��ޜK2�S�{#�M̵B��W���,s.n����/S ��VE�WR�1�p֧��Ԃ�޴=�}E(�N�".Ԩ�����н/#`회�ո��G3#���pG��+S��e�6|����޶G�ר��jI*�ާt��&}����nD/I~1.��v@�"���^`z#��Q���+"��r����gK[v�V�7W�+WY�PyQ�=~��:���T��O'9nh9�������u1����;��A(n䍪�v�)� gB��<cz����(���:�)+��ٸ��g�m焋�o�o�-��7w����R��GM�׭�����vߩ	�}]Q�4��d@N��l	�� 4�3�a�䍳{�T�"�z��Z�d�D����ӕ��t��+��6�퉾��2 �4H�%��� ����	��s~w�T8T/���j=�MGZ}m���sOq�Ƕ�����_�U|j�UIb�U%��91��#,���Z�l��@�W�]O3���b1i�w	��7��<p���`�����	�;3�|���J�g��3���!�x���)u�����=�e3�^]�4
8���;*He���q�.��j>-_��O�A�8��P��=��u
���r�|�L����j1vAQ�"+k�˻y�Q9�{
*�9Z=�2S���O4M7�K���
�����+�r����kU~��_G��CmUQ�M��7��o-�C߬M�m�	/I�.&:!� RYJM¹��Nኖ�~�a����*�y.���(��"/9�c�}�l�������wX���s�JѨ�a�:��گ�s^���ʁ!nc���Cx�4{W^I rk��zq��}�V��>�k�ܛ�������U܎��j6�;5E���YH	ud���5콴2U='�;�`g�|c}����9r����p�Y`Dz�Xd�̄�?u�,�2���dE�/R��\	���L�/�N��}�܈�~�~��T���*�L�E�=0��m%��t�dؾ�L�wS�|.)��7�x�����q�竸���.7c��SV'�ӊ2�����$t��ݺ�g	H�Ζ/��n��UǦ�+�w bc��h��&Y�y}�:l���u0��#����(���r �c*e#uS�<�wA�N�{���/V��oٶ�����G;�@=��;N}/ԃ�ɖvD�Fc`S���;|�~ǙB˄}���oF��p�&b�R��`���a����:� N7~5�U��4���J|)D}z��nP�r�z)خ�L��[8n�Q���2��wGע�ʄl�z�Kޯ��.�?ʰ�7���_OȼL�ѾC�"��gzxηǭ�f�����PjW[㐺G9���@=7�U#���v�Il���:t蘤��>v߲v�M�>9�J�^�V�Њݤr���H���;��\G][5}�@��ٺ�C��vg6}�n���0�L������B� �Ά���c#�6�>�Ӿ%�T�gU�ݡ�����Q},�螪:o�RBW�6b\���9�>��lbې�U���h��.��cء��[������Q�)v;�rg��L�Չ�����!����(�W!�j��aMT���魩����s`ߢ��C��Og�=�ǀ�}p+��}EO#�n���{�"���|�dH��EuUwm^��H	�q�{���C��Qy������oF\
]XfU�a�>��p����[ho�	s��HZ���_h�~�}1�k���ZTCޠ:���u���G�Pɛ�� ���?Q�}�*�܎�z�|i�FzN��ឺ�c��K�>>��/n|�k��|�E.9��+#�^��S��ե^Պ%xtk���뉖O���|%'0�_nC����y��v�T���*�h�C�8��K�iC	�_6��b��k�;7�)9&x"���Nǣ)�_�v���gz��Yb6����u��(vVSMR���)`�k���y���<P�n>;��v��M�nˎ��y��|�6:꺾�x��a�"D�n�A�m]��XР�n���F%�P�0gȱqY5�qN@�~��v�	<�|-G:~y�73���tGU6�z��n������hY)o�a�;P�"��� 5���]澌���վ�����8���Ի��}\9eu��d:��q���˔ID��U2}�L�NYQ����(ۣo4�����|]X��!�ێ�9�s�"_��6}%��P$�[�j%5�{'�.�};��z��_��{�W���-�3>n�
�zG�;d���WrW��pS2���Nc/�8g���������@�ۘ����r"ۯ	�n���O�moH��tN����e
��L�0�T��]w~1���������\��1���p=ΘYi{��8}�6�4���w�q*���T=U�B:h�h�P�4�"�x&��:o��5�k2=�7�(�:!���ǥ��%�8D�vDܺ���FIh�#H{=Fj=݃/^��Tr{p�r��k��mWQ|�A}k���:���}���U>��Y�耬m-����/Y>Ś|����,��&�6ʬ�N�����=�3��M�K�vD�"�GGJ��`k�mԶ��U�8t+:�m��2��j����̆��լP3�l���ȴ�WC5��U���Al�5:Ǿ���%s�:�m���K3Bc59T�<����tm�WF㻨��z��a���������nmˬ�n5plA��2��9v�e�>s�4㚗�t:�蝹���}+�p0�Q�k.k�������R}���� {C�{ǚf����=(uG����E��Ke�p)��Bn|o��Z3�w�n+M�����oII��@�Ɇ��s�Qɕl9�M��OZ�U�_o������Uנ�Oo��A��n�/�s&߽8�e��)쎪v�bUս~B�����Z����;����"�:\F:�������h{����>׃�bA�
\�/�~��Z�:~6��E�̳�z#q��G��+�N����Cgr�\{qv��u�(Qk�����@���7y�jbC�I�DY���3�1�*����g��sӢ�Q���+"��r���}��j��F���Ǩ�=�;��ȵ$Pg@����J�/���-�7}�<7����ے�8����Qپ�sG����p�t��7�,�(���/�R$Q�l�L��"��	
4M�.��b��U����[�[�I��ZJb*V�$4H�����p�`;\��iY�����Knv���]	��_Y%w �o#��Ս��������<��NS}�)*[&f�d_X<c��p�T��^&�c�o����*<�nJh�ڽ�q0�;ws��ܫ��>�|��ZǶSY^s��ޯP��僑zT�+���4=���=��x=��T)��:ۨ����9\�����o;����'�d�� sPHӧ:79}��{㴖��`�t;���iŦa�}m�&��{k����:f����T�'en�xt��K���0�����^O��Ǳ2��S�-5�5}F�}<�㇧8��� ��
�t�v�����=�Wz#��>��s�T2$�Q�C"zw�	�׽/ƽ�Rj��oɾ�G����홙ᾫK`/VP+|�1#}&�3�uϡPځ�c-	��OG����!�U�>�_z��srzu��IA����6�*��O w����o��9�D��6�P�Kj�s^�W��TT*�=z�mpu�H�}y|2#����>��o:�9�ϟM���P����D{��?W���O�j��ż��=�|n<S5콾���-���ު�+#�-��9r���
ł�Y��yT�L����ٳӤY��s8dy������ʣ�>����]�m�ߔ�6��^v,p8�+��$��4��O�eZ2���\"�z�$�D�A��mȮe�-"�M�M&Uժ8�o��X���U��=�K��jaHGk�@��ely�'0p
U���IV�U��� t�VE{|�u&��[X}4"�cܦsއ@osy��~�����iۤ�\�dT��r9O�o�.�Tj�\`9��;��k`Õ�rr�r��;J�RMt]�^��H�Y�R�,e:X���o�=�Ӊ>�u|)����}%;�w��r���s�l��C�D^F.=��e � �r4eSS)����9��\/������=��+���|9o�͇���>��u��K�A��nD�l<�p�<�a<r-_�s�0��צ!��YPjR��.��w� ?�U#���`���q@	�;�}N�}�w���~��=�:z�TO#tg�ӟ_eC���"�+��}�gu�뎺�k�,��W3ˌ��|�H�E8��=��*�d��P+�u��Y�/Mb���%��c��6G��1��-���s��6fD@��<UV�+bđ��`� ��Dl>TX��T��ԭ�1� ���G��t*�33�=�4�ϙ����*�MuIh�1�k��Qk�W�����pci�iVu��j-�;a���4tw;������_q�+��w�v_Q�FI�nԉ�-��0���멤�,��u]շ�֐�S�T_��mysO�G��:3i�E��^\��8^�A��ѹ+�t���U;�PYd�q��ؾ��ĭW�Wۓ/�x��`U�|��(cb�[\nwb���u�r cb-ʅ�Q��A���/1��^9����Ii	h'���Q�5�^�1�WE��J;�������]@���2�M=�n�v�dMN���J���-�8ֳ�{ƣ�yp�5u�8���q޺b��Hy��M�T��{��F�\����E�x����՗�7<]1�&�5�R_�1>�;�#<��c0I�&b��WM��3s������#�?���3�T|=>NI��ԧ�>�Kc/�!��T�@\3f|�\w6�_qؔ�z���D��g��s8���o���	����Z�=�i�ݧǄn�P�nS�s**�y�::���=�:����!���~�F�������s�(�؍�X������"i�{ѵA~.����wMz��r��C��^�.?]�(��Ih�g��1�;���ڽ͘���~��	\��4��4h^�G�;n;��W:��~�@���]P�����c�<��UC�	:O��S��WLI�L�2̸�7}��8�=����yX��	��TLeBs뗸gfX]g����p���@� nb�S���ۯ	-�5?u�s|�=~��~�=vML�S���/������{�qО����#���[��Pz��Ϩ�m�삓�Ƞr�m���3�u�n��.�+I��9[vwڭ*�i�m�X�/{��g�����2��-Ѷ�זMS��|\[a)s��Ͻ��e�^�wj�\4���MȾ�n�s�]�y��x��	ѐ6Al�4�SP��ף���b�+���깪�X���C�q���ZNwT;�}qW�(h�4LA]R+�/ǟy�c]����JQIA�Ί��ݒ4\s�lq�D���ɸ��q=��7.��n�Z7�*��"��!OCw��qPþ��Q�>��=P٨�F��6����g�� :���3}Sq�֣o�~��j.��w�:�t�^+滓�MsRy���U*�8�%*���'=��X�]e�G}�/��{j��z�\Ҋ�$t>�����6puԯ���W�����W��c!�Eus0B��qX^p�w��'�-�	�u#;��l^������=Si��Ҷ�>�uVx��n5.�9[���N�H�W�ϝ��g����8��s4�z
Mҁ�a�:���a�|V�+�]	ɚ��h^�� wϹ_ꮽ!��Ӽdw�W%^��޺��K2�E�Q�|\�ޛ���\3p��RŃ*q枊-�#����"�UԸ�u\5���Rz��9���zK_G݈�d����|;�}k���{b�;WJ*�D;�����sU��ToPhC�Z�k�K {4�äe��������+��\�̮���������7F�Wvtf��׽�[��6Y�Nr�.+q=1����w��zU��K�\;0;�r���}Iv��5��ĩӾד�Ɣ��%�+6�O�*�Tc��Y78[A�G�h�}�����;�q����{w)3:����,c.B�x��r�'\ۅ����Wvk�4R����0��;�OnNNsa�|kA�~�Z�Y�FpEbEv�Sv@C�(�������Ó޶Qf�_Mr���3�ԗ�6,1lU�;ܯ0�t
v%���̞Y�r.���J�I�O����5�"��JZ]Q��+��pt�J5e��L>�'�K�jY�,���>��*8���dN;dm���
��wԦ�;.ra�joDo�����/��'h7�K֘���=��9N��S(����\��	�xGtAa��g.�0�e�U#���g�f�����bUg(���:n�|��'W��7�Q��;�*4$�yԵ�ȁ}9tK�=o�
��X���b�Q���]͎6�����6C�r�9W$�]�+G92v�}՗��G�8ۓv�+��^��TU�^�̓�٧�S\2�Vo=�宻:��hN.�gote�үjNh��3z0�77�Y/N�{�?M+�0y�ۺ�*�؉ooMER�����Xm���^�Y:�`ܜ;��תP=��7t-�p��g/N���������K���k:,S��5Ei����Źu�bb��&���{���J�򱥵-&�;8򦻃pn%9��d.b�ďE���/���<��W����'��F��\+�M�-a�s�ִ�Hz��ꏕN�hQ�o�qу��s����Q�Tj=�z"�ӌL��C!�!�}�(��R쎠�tUɀ���h�
�j$ܔ�vmc��w�\�x�c
���v��� �s�F�̷H+,�J�,��%���1Š�Ճ��4�-	V��N��8����EֻӺǑ�iSm�m�`�F��x��Y��{�X��Z�[l�p�:�G���L���������س����A�u�X�V��ޚp�ۍ5t��l�(�`�D��i��t���}~ΆIb�Y<�zD^/M�پ�a=l�T+g>��Fv5 �1S��W`�47��~�J���8.���.�ܻ��U��3�[b#���c����n7��TZ�u}���U�'A��3��$�x����V�>Tf��P*�v��עދs�p����#���D�;�Ӧw7Y��~�E�8��boz�:����tVf=1J;�u�2[\W�O��^N��h=�V�"��f���U��Yt0�g� �J�L)Ѣ�ڕk��m��5h���n���D�vB�8���@ۋ����T=U�R3z}�| �¹��6����9�����m˺蹋�"�u���3&�5���%˔�nc��'.�s\�7.��,X�wTPS��r�b��5���\���+��i"�\�r�(�wup�nk�+\�[�4H본�X�5�C�#����ۥU��s���ܪ-\��N�a�h�.nr�٧w �-�sr�U��ksr�1]\u���#��[�5���24���A��"(Kr�6�\*wt�i������gu����p(��$Q@����DM�g5�fe�܅GHw���\5�iQ	����Y\�ٝ[�'&�0��g1g�I�b��NkCo����ڮ-�D>�:���A��T;���tzF�z�rjt��S�l�G���ڻ���6�\=Aoz�욽�q@w�g鈓Β�9��~�/ܪ|��9��<]@����{�q�^�"KK�(�Z���ʩ#:�8�|�V������.�X��T��UO'9惟>�8����v̙�_v�z��/�=���;>w�׸�d|7�,�̢K�:��"���d�^���)ӥ��'��'���<��3���s+ܨ���ޤ'��}~�����@r �H
{���N���흟iD�t������<o��n�n"[X�D9��w��Hi9�$zz��}�G��9g{2��uӘ{�4���n˅C��y0:�"�=;��;�>��Dt�����,��z�>��)]<Ǹ���U�[�rL�
����H!�B�ꗧ���Q�MC�����Ȟ8zs�ࢋ�-�K���r7Y��.@�}V�
b�s�H�����#�����]f���m]э��!�x���h���E��}�zC�2����*j��e�";]3s�楮7�s^��)��4eeF�<�x��$f��(\����;�8�}��i����:�����w���l�=�0�:2�
E{����$�|����'��;��!�b��b�w|ޑ��o��N�/$BTxݪ̭�P(Q�]6U��h|�vqGNA��:wP>/��U�uSq�<���Ex�oFP3��P�J�]����[P�{��I��,�(�n��p�×��}켴25U4s�C�\gU�;9���.���oH'6��Ʉ��۟Z�=Uouh�V�.�[���q��j=���|���8�p\w�xN����9G�uU���}��n҃X�Q]��a����ʯ�s%��Oы��c����|���KPe.�Yw��X6�!���GV���T��]�:w"gP�Яꞣ�qNG)��`/P25u�06o��*pw+�:v���a�w����ϗ^��{t�%-�,e@3��'��S�ʸ���Q��C��=�)�V�j����t˘�B�WqY]Hr���ž{u�,�J�1Ȃ��%#wt,	�OF��R*?W�ý�/�����X΃��{���lv��_��}R����l#|Ox��T��z���Qsu��=��e��D[ʃ_JW�rH�;������}wãNIkZ���;�S�vw��3�����	��P(t�n"����ֻ�Kv���9n&;�Z����c�ȹe��é'��ahs�WK~�Y���5~����Y�x�����˸(�ɺ��Q��l�Mp{����ry��]�tj�v�H7AS���҂��ű��[���D��p)ա��7�D+��%D�J��Uŵ�\x��ޮD��w<���H���T��ӗ{�(�Po��gOC�ꉐ6���+zkև���1�9��~��17/��r�y�p�s��u:ݳB�%�T�߄�� �SB�����Wض�5=���fN�/�"sђ�����A��K�1p<�:�MuS$5bhD���7E�Mu�G9u5���'�O�5�w;s�_r����'�8U|�.�.��({J;u�w�����V��j�R�P�����>��Tw����6��t��}�|����
�_����[#+T%7�*w����k�^����	^kد�\��_ں���@u��t�n|��l����YD�����|��](<&g:5��O���}Bn|]	�i5A��w9#�y�7�K���f*n�b��隣[���Vl��7���TB��Ƹ���ؙ�x�?T��?��ǥ���p�]����TK><s׾�WS����x��D�f��cB����W�:N�1��O�b�k��� r�MG:�ɺ��������d|�/�]�1�wt�WV��҂��?]#�p���<5k�^xv~�Ƞ�Gl�Һwb���H�K����@z�2pLy�/i�n�F}��w'��؆!H�B�C{4a�.<�+��p=Ǉ�����uo�n.mYr�j��x!�\Z�N����ţ�4����_�� ~���Q��ʀ�e�������-s�u5��\?�f��=TW.����wMz��r��C�s���C]�$�=#!����:�m��*/��=y��p/�J����X�4���G��=��r+�p��vײ�tn	�{��ՙ��MtB�K��t	�:�e������[�fo��x�oH���l�u�u����)� c�|z��`��7���|g@�
P471u2�N}o��ޜ0I3龭S�e
i*�>��]6�U�ý�����:��C�����I���
�D�#}�6W~����+޼3�ַ�k�d�:'�_7�Ǘϩi7����뾸�̖}�T	D�]R-S���?B7�z�u�����	��1nH�'��Ϻz�=����}�^���ț�U�6�������������L����\����9򗺤uCj����@�	�r�}���u�����?X�y{����}09%�<�(Ȏ�fa{��?�������Uq�&�wH�ۆ���=��#ܶL���}CNl:s�炍62$��xV�_�٩�愈S�fy�uǁ�b"U-ǣZP�2�솨�Щ;�g6	8ڍ���	إʠ�A^C�];�f���/�4w���\X�ܩv���d�1	����
kL�O=���D9{��B[��]{��yT˱t�j���L�G�v@��_��'oOoz�l�Xz1��T�{�5Z5C�W�р�{����B~�)l��vQr�Pi���Ӎ>���;i�����]�`�@��á�r���t�*�D��	�޻����AI�l�huMϱL�Ǣ-�/ד��N5o���g��Bc-m���ރ�7\�r7��#��XfU��(�1�\X�����5�W�>�6�VjY@9�L^�Р6=+�ϝWj}�H,]�C�rN��"�J���=7����@w'C艜�Fv��L���v���mG��*5u.9�����>�����݇]T�f�A�c6<��e���Y���·$��9���T
��g�Q�qB�x������5!76[F������f��9Zi��ԐU|f6b�X���R'��fC���[�s���78�=z�2g+�<9tup�}�E���qۅׄ;ʔm$�t�-��ػ��9Mi�4��������	/��1t�;���eyΘj��W�z����9��0f�\�&����x�&��+y�q�~7�������2�r;�1�o�H���'��g����{�mj������2֦٬	m����Y�����(3�D[!+z��Nw;}��� �#�:�]�y�:�e�pv#j5u�1�@��=qI�٠�R�݋��^%Q����I(�uu��=��8�8S�˜<��Q���*�����R6�� g���'��P��=Pa���O���3���^�eP�z��jy���)��9�E�ڋ�f�:���)%)�@�:&J�ក_Ŧ��j�_ϧ�<M��:��\�RU����C:h��6B�b��WQ�S$5cj�gx���8W{z�6��]U�9�A����c���-��vQ�~�H��B�=�e!?Gc�o�=jri� ;�漌s�'�'o�zu�џs���M�t�q�+���*.�2�J��#��d��R̎1ٙ����K�Jƽ�2t�?ut(�>���>S���9�ϟM��r/zA(�ܭ�Z�o'��)���u��	�aq��^�
f{ų�Y�2��v�x^P����6��6�%�S�~�ӡ�S�N�s-X\H�.����)�K��g|�����֏J�����׈���N��=�ӹ3t,����]9��X��
կE�5����y�%sO�s9\�`tO;l��o>������WJ�̥nAQ�H�G�G#�eχ�*�ٚb�f%bV������6`�k�B�=���`��(u"�ֿQ�����F��]��l�����X�ɭT�[�ruЮp �mSK�r��~�0��Z�a�ϓx�n� ��pŮ��9��3Z)�t�n��;�ov&w�灞��vdޫ;�ҳj�D�� ��\%}��VWR��F7��n���NјzA�A��;��;(ջ��to�O}GC���걝����P����9��R>�XD�F�/]�s��j����:2ڏH<Ͼ���3Ү�кG9��PM�w�G����]�x8}'��'[X<�X!��^���@@0Fꂱo�}k�q7ݠ��+�>���b�>ɕ���;�WG]_����. E�L����@��szt5��0�e�G<�߷w{�f�\Ͼ�F4�ސ�:��и�TY@���v��s�}5�du�]b�)E���#Z�A��0�+<rN2n#�� Wϳ�*��S]F��\	����3�.�kd;W�o��!G��5����H��-wB�u���g/�����|�/��2O"-j&6c'Z̙o��4�j��vK4!f����sO=t��n�����u�\� 懷���B`����d��q���%����}8�t���^kŞ���]�3}U���O�zօ�b
�a���#��^Ń�M>�Gp�����+��Sux���nF塙:��i�ȸ5.K�������״�؎T�*%ݯ�8k�M��=��篓��I��Ӯ���.ɜ��&U��CX&���m�۶���,n��׽�(��fP.[tm19��sr���^�����%j6�X7v���И�T��K��٪<���XIz�!\��J�o8���~=Ω	Y��c�M�8�H>�\���V���?�٭����T��"�t����j	��˨�׬���k��o^���K�ކ�v\����k,z�w#�߹��u&z������\*k�|깝ϻ��}�A{���Ϭ�*��g{۫�QX<=5�Ʒ�d��ٖ{����8-�@Tjt���}\9eu�k�h_ϟ���w����M�:��Tƴ�jj;I:z"Ni���:�/L�Q�xj�ꊈ�!���r+�p��������zv=���9t�J���IU3�O���qS(�=:����3~]}�GQ4�^�irF�k��w��|�M�(�Gr�[�z�ǰl�K6�	ѝb�����ɉݛ0��"pq��~�u���2��.�_#�F(�T��l��x� kfcg�[ T��kަwj[h>��
kzD��	�h��[�Դ��;��_~�����Es� 4_���E��$����K1)6�������ڦ�U�6�U&�5��S��>8�2e�qb��M����]��y{(�*�9�:��c̧
�!Y����k]Ӳi�u���{��ze!a�<�,�U�;{�a���KX�g�ƍ�I^�l�#=���^�o4O6���`�y^J)E�����<��rC�;c>������d�wux��Ȓ�I�q�:�.Z�K��^ǒX׾H��}*���r2a��P�W�_t�y�q�����_{�w&'�_Wvm�qy�$��۩��f"��s�jc���sO=��ɞU��\M@y�K=\n���z��P7׆X��3�u!9�ԧ~7<��'pช]\*�/ƣ����<�E�4/'��{j�ȳ�Gw8�F����}R3ѽCTg�����E�=�YJ�'���Ԗ̺��|�ܮBy��3�����8�Κfw"\V�}�]a� f�1ʠM�[�5��E�-952�ޣ]eW����N��T1���l*�z|�r��ޚ�Gn�}�]g�դ�>��+={��-�=�Y�麬7Gx���L1�����dC��O�z�X�և}V%�v�Q��Jy��[_�3�w�2%�8�_�͇H�U��v�����3��;��w�n���n
Wan��Jd�qwϷ�9�((�U,*�3���3�b��f����A�^��l!�y1��5�]`�E��+b�dOu>�(���XS�e7�H���:�|}'{i����ȹ*����)ӻ�p�r�FO���d��C/����G�,Z0x��*�YP뮖��:����L�9�PQp�u-�G}���լ�8}G��L����*�M��V�g-IQ�ـy/�HL�NG�X�=6�ۃ�wЯV�^�״Ŏ�GS��,����;C�����t���:�������݊���~��6��N���}I�	�_�B��w>�Pgn;Ԅ��ϯ�;4��@��ݛ�_�K���_F)^ ��2�F���_\M�kȇ9\��Lf��Dl�S� �P>�o��)D�NOi x�#�O:�_Jg���X���}m����0��ʽKq�]B0���E{��F��3�EwUZ5j���p�O�7� l��_T�ρ|qi�i�p�^`]��t����E/.�TFw�J<zsI��:�)�_�9]F��Xڱ_K��BFٜ�\}���N߳��(斂=a���7������E�����=���+���n�T'l�K�_���<�q��z߀OA;ن�Ld��W���'wBߺ���<��w�{ѕ�e�*��=��3^s��b�q��U��kr�|Y���j��H�W�V�2=���^�gZ��<{�n�Z�	��������i�J�YLsz�3rN/�gS�91�K���:��T���?$&���11{/yMҋ�����u��j�h�קx�v����m�7�X�I�C�R��o7u��G�\q�v��Jl�Xv�٘��W2�ڛ^Wn��(������S����]��io1�e�V�`>}�C����l���U�z	�����_��Q*�f����6�Jy�.�]�k�T3�m��)HM�m���L}��q���:��7���[ ɘ��pxT�[��a�n&��{R9���n�}�6��+��޾���x�t�,�!�cb��\�T�����wsg��"��!��/.�Z��WE�9鱗��;}�9�wR.-(Պ���^�2[PgQQ>ΥL�XWha�"�j��r�����v��Ogj�OsL#���U�,�	�I-� +���wŇ�s7.���4����p�yU!�Tu\�}g��zx���3���E>*�c�c�z���̺��ـGtT�%]3���b�(�jgV��0^�w;���A:V�n4��Fw�����}��,����x�S���C{(8凫f7q�.���}h�g{tWM�OR9r\��ݚ�d�B\X���!��i��^F��x&�t3���ᒆFj�v��LouBT�x{��M�\���.��È�:{�,���$�u�vӷ#��2� �ml�vYӗja���r�V	s�t�]nK�� i�
0����-�鯖'Â��L��d� ��,�=z�[7��V˨��cU��F��ťW�#�=X)s5�S�jZodx}�r��hs���\b��,�3| �ޭz��ܒ,�0�L�,��Cy��Zڜ�.
�����hs���BZ᫮�H^lL��NVkͅdID&�L5oM��>�8���6���Ikc!��V1���DS�M3��
G�n��M�g�lۭ�@Ƀc�kq=�"�u���m.E���G��`���;É�u`�Ӵ/��uG3�?}f���Q1so6A�a�﹞���y�0���v��"Z�B�0+�:��1YiN�a��'T:
p���G��v���c6�
�CKc����iz�u��g5ä�y�w�9픇�����E����|�G<�Ý���;~ې0�wnɽjHT�J��A��Dw\y���4 �S�v�_^�J� ��S)
3,ݽ
�-���i�>�΍G8v!.��:���!eD�+�:������fn^��f��|�xFd�ȷ�W9h!�M���TE��,z�n�D��{IPކ +HMV���w��<|�[X4n?�`�f]9��Z�������Ď�d1V�i�4gz*uN@�����{ٸ^�+h⫷�֑��~��@��Z4�3_a�黎w���g)�,���wE��8�ݴ���������r�]݊�s�;��b��wWB�
�k�n]�]ݢع�#��]+��]E�;��s]����*#p��[��.�\��tܷNY5,1]ݷ;�S���I�Y7!6�]�k��-\*.�բ-��.�占��풋��1��Z����F��Nu�+�r��S�\�(ւ�q�q�EN�˻����Q͹9�˔fcY��عwq;��H��\"+��h�jH�]u�	c��w#�cW2QBS�r�`���&6$˭ҨP�P��P�� �\3k�����{2�k�Z�9��>w���}۳�#��q��pܭ�L,���I�
ٌ�����=��GbIUc��3{��?T
O��Tm�S����¸����CUv������;�Z'n=��=�و�u�g��N��H-:.�8g��10%o�2-p5����9��_�o�vj�y�zeZ�S^�@x�5����]�:w&b�d�W=G�Y�cŀ�qy�N���ެ[v⪲�B�k����Z��A�z���u8�R��
�W�Q�<�Hd���]}�v�]J�5������]��������+"���ב��{�4@ѕ�5�2�w�+�׳��P57s}��Tϙ�,'y��걝���T=�;�K� � o�Y��*��5���C��L�w�0# tutgY��e��"���į����s�@=7�Qꌍ��x��OD̿D�xl3�}��{�:#8�}�Ҹ����Kv�����?p��^��*�'r/��M��+���p:��]}2�s�x�x�^zp���z7"��b/�F��q�P��_[�;�o��p}u��r�6�P�6b]�B��A��t��5c�v�94��K�7)Od�o�8���@y侑e՝�'�[�§�h�Z��r;���.����a����4|+0P��ל�`����Ľn�÷��4fu�Z/h�C��k�r�xP�F�V]��c�*�U�ȜÕ��Pks�zu��>�3ܬ�ȃӌ�鋀����:��6�Hj�kn����[�uk7�8�*�(��M_��^J�E%�t-7\Odq�ݐǀ��p)v_Q��N��E�|�5>IcE�y,�-�syP�j#�޶1�WF�����OC20�ç� ���^z�U(0\�uc�܂���dY�	�mP��zS=i��t:�K���{�Q��޴�������{�r��5��gF���rG~��±��u>�]	�i5Mo��k;z�T�:C2k�٭W�M�,1ϜRg�3�w�T�������Uw�Xx���v�ߍV������&O�.rk/���b�d}�#�uWnA������^޽�u�VwN���c��O�c��6'Y�F	A�^{�T�f���(q�`O؝�E�
�v@s=�;������vN���N��ik/���w�=��/�ȅ����T9ٝ>���W x��:]�^���+���lT��V�QK�U���5J����Q�<�;1�Fy��&|O�.���HG޾�{c7�PV�-�s�8˫��E� 0�n�Z-����K[*j���]��[�z��S�����۬<�:Yh����!�}^f�}�<�/��=��ͱj���G���,��s�Pk+.�g�ܵW�.��y��l7FK�����Ϗ��y\�73�Y{����_}޶/窶�e��Q3�OÕC���R�����[�foϯ�g5��>���V1�>iFd�p�����v�;��.�ǣN	gZ�@�
P471T�]*n��Usg���7)%�=<}���x�yTNlC�1�2O���.l��;0�sK�����]��X��ɮC�N�H��ա�C��C}�i7������U��4x� s��lQ�yQ=��C�B��h@WĤy��{Q�rC	�3�+x��t��7�^糲&�o}骏9�i�b�Q*' �9:$�x�<x�J���3�&Ŧ��&��������������-�fzқҧ�G� �Rfojc���#M�{\*⧑����5�WtM��!Q�����Pn�t#|��/��h�wm�p�B�ՃӰex��er֬�=�fi�4���4���7ӹ�tU�ڀ|o�[UTc���N���z����z�z�+����釶=^Ox��H��d-��W9ن�J��]�CT����ͳHϓ��y�V|�'8d�!#�S����'�ԅvX�{��o��Mӄte��c�&4�4#S^�۫+�o�;)�R�{�Zmu�l<�D�N^M�zʝ�ɪQ��G4�o˥�J�Kk�V��='TYFS�Vvo��D�碷���9j�F�&-ƍ�qy[����/g!����zN�s�� ;��66g�
�g���D�FǱŜ��IyY�*���'��;�����Ц��%��z�n��s-T�q+���k��UK��u\5��>� ��~��.����l�(�_��s�@��ѽ��=�.���I�8gj�Ux�Qp9k�����d�N��+W�U���oa�.7�\�=��q��s�QC"�J(�	a-���ʧ��{��/��Ou	0nQD�5;��Vw���t���GOqY\�9g�ב�}/Mqȵ$��ĕ(of���T|��%�V�9��=}4�=|0d{���v�g˹�v�8�5\�*�.��	�;Q�=\���;z籭�=�|$���S,'��xH-�`]��}���z������h�,���.���^es��M�(c��(^rL����a��ս�r��1�W#��<�wI���V
ꫳ�t��ػ���TT� �RF���@����ȁ0��-ۇ���9�9���釶:�Vk���at�DgC��j�UIaI-N��@]HU�K��� �5�MC���@����WAw6��.��ta��(.��ֵ������,�.��h��F�슘�0�9-�\Wq�]7cc��v+ȐoaW�s�>�r�"�r�/zZ�"#F��s[[}��Ok@�9���j�DK6A��V���Q���n�k��l\7��Vn�Jw��:9���?gx�A��K���>��B��WQD��zho��xи�+ƒI�� ��ޮ��0's��>ꐯ��wF-7�x�L�v@u��}B��zJ&;W�wz.mC��*.��>�;fF���	�Ʀ�x�{�ύ�uT����M�t���W��FT
�e�*(N��3�����&�=���5���Z��i�%y�e��fC����\���D��O>���I�����=�v�H��R�|U��[��s�W4������1���NG�� ����wZ� γ��9��՛>�}ݹ�'(�u |}py�=��+Z�c�e�bN����gn?aW���&r�i��j9�Q���ߟ����d�,��a�<�.S1��e,��&'Ҳm��^�O��e�=ۃ�GWZ� ��㮻.=��u�1�~�E��43֪�����:{�q4w	�)��7(�b3��2����5�½��VEu!�9�c_=�F�$������$��s=��n$S���x#K�ϩ�ޙRW���y�|qǺ�r��c����s�|UeA%n�'L`o�^E�
�W����?P�:�k�d�����?�{$��R�y�Ǒ�l��ڕ�0���	��1_s����+H�܄�Y�n_��F��,���#V/�kcSz8�.-�+�4��I����"`�ϡ�"�	x���-\_@��۽d��&W$�����<�:��f�g�g-�A�į���s������OJ�^����RFs�޽Ϥ�� '5'@��A���ِQ|v��Ė�a&:����]�tQi8sd����>����͎��^q�����g��@�ut�Y �8e�Z�V���K�m{��N�y��}�3�6ޟ>���w\uUq��uE�P@j�H0
�=�|!nI�[aG!Gݘw�A�ڑ��}l1�{��9�7�q�՝qW�����Hk����0=����Jj��z�F����W���Ty+�Ŷ��[�Og�g��`w���A�y�n��0�.�>�C�W�W���"c�\���惑�K�:���2��{>*}��-xG�"ǟ���=t�o���5�x]���GکdY�N�j��kҩ�j^�\<�.�G+r$G���j��K�k$e�Vs�a��R]������\pZ���Yt&9��;����q���׼{AW7���\�d{�)q��Up����W��s�q_�99�?��芜�tK�0=�M�ߞ2ӋmPoo�9��
����|,�A��IN���h��I�׃1[�&Ɲ��0��Y���l����7)|v�]�-Ӛ�ͨQ�<����n>�N��Ed��J��� h�C���މK���OF�0\F1#����[u2���^�a�;z�7��lj1���4�[�4���,.�Ny{rx�]���n��y4�(z�WL<��^�s;��_^z�u)��R�W����\*��>�U��wNҹ�!~��Uy���`�hﺪߵh5Q�N���fva�WU#,��c��Q��
�N�tע��rȮ�<6��p��.��z89zφ{I���H�Q'����C�yQp7�
�]Q�B=�Z�5��L�0l;Z�7"���T���A�g�[�@��"g@�ʡ��2���u&r-�3-Ƿ}��[�`_��د{�&r��:�e�����s���.�ǳ��,�RA`��hnaN���Į�,]5� f���jpOD�����F��*��}w�;4�� �΁�N5��3W���v]�����9��X��H-�A����}KI���>7�]�������꠆j�	k��w2�"4x��@�4O��D��a�\�'��Μ�����	����{��þ������>�`���Gf�M��$i�Q�/O��a�Ŧ��j����@�Շ�]`bT�����T�I����S����1���*��0�W6.�&�~�O���7��	�d��@����}{����Ce����=0���Sv(�E���ni��[�[Zf�Q͐�wP�g:^oy?q�Ӵ���'W�ו�%]u�����^�kc�_=C�{ca�ˮ�6곪b��jo�`�����*�\Լ�ӎ�fן��2f�^�y-Ql�&�|����DoP�*M�Nŀ�<v�E�ѭ3b{���1�e�r�T�wW�}�S���}Ϯ���?tS�p�z����@� �a�~�z���V�0S�w�o��v��F�}�l��eU�=��G�H闝6��|��qP�7Sj��Rk���z2$�^���.*s�w��hz����_}=�Nx����m��T�A��NF���S��^f�Z;Wb�w��+�����i;�c�����eW��\J��0��|̮!C��N���8�rzT�ӓ}��G�޶/���芽�%�	&WO��u������vZ�&|"�C#vo&��]VW[�����^#���H��Tg�z�q�u�(e�U�q�1z��{`P�{b�W0})��o��"��{�W�%�P+Y��{�q���^F�K�\r-I�@(�
~�th�f��-���7}�d�9�sC�F��=���8���w;��.��<���f�Iw�0����Tz����9�`$�G�%.]�ի��97\6��҈]-b��]DM�o:�j���<�g�Pky@A.y%g�YPߨ�b�m寑: X�>�,�����e�)�}�%\�:����4M�^�+^��+��YnAZ��&�owgY�>�|W����f������	�_�B�gs�A��J��uC�~�Ox�dRg;P��|�g�<��l �@��Kf�f��uD����3�9\�����5J�����ͪ�w,����aʩ��E:��[�%�2 Nj$�2[���|Ud@�zj1n�<��پ�*��@��(꣇���mx��Y��^��T�.Ijo�@��.�*��x�]���H�a]�ou��y>F�K»����A��O��.:l��зU]F��\�.w�	�h.˳�=S��~�f�����k�S�k�T�pڻ���<s����=���+�WI�3��-:�Fr���oiv,�����dV�����.�6wt.����<����*~��Χ��Gٮ�/�l��j�|a��i�+�{/'�3�c5uZ9z����gՐ���S� z������u���/�F\�] ����-�����W4�g|��eq��f}�*oaiB�5k����/ǣ�R��sƻ�\�c}$��/j-3�73��o�i��Y�r�n�z�NU�Q�59!P����1碥�Q
��s���{6�f�@r�SP��.d�-�7�+���w�=\�����x�Ƀ{�O[}@#y����.4燤[�x-��
���fXi��z�Y�բ����f ��WP'꟫����ޜ�c�2_ϩ�S�[���q4�hZ��&.S;չ���0�Ȍ��;��%*&k��{Kq5�n;\`g�����WeǷ���/sۤhY)i�3��z�6(n����v���g+��Ji����\zhr�pbk��z/�����9g�ב�|��=�a�\V�֯=�QO_�MGi'A����W	'��t��ǪB
�y���%��{��,��c�������wW�-���d���gOB(���l	-T9��<9n�}�_q�#����u�/�ȩ̞��y���\��Ώw�޾��Il����O�*�C�� ���yQ1~q��]^����ⶲ�<y���#���ی�=}ul��3�xۂu2����
�l����FEu���m�5�2zupY/��ӛoK�&��:�f�DK�,��T	c�'�;//� ��O��e[�j,��M	��9�@<F-��>�Ϗr��N2n;���.#�:��׌�ԿPd��.�*��Ļ�0HYx���>�NV*�݈p�]�hw���u��~����+[Z���V�����5��kl�;[Z�ٵ��m�ŭ�km�������v�����ժ��6�Z����mk[o�mmk[o���ֶ��kkZ�|��ֶݵ��m��[Z���-mk[o�kkZ����km����������m��kkZ�}��ֶ��1AY&SY�S���Y�`P��3'� bG����(	������T��[e�V�@J���U-�*	)UEU��R�QBE$��Q!D�Z�m��UR�(�фD͔m1��Y2�Z�2�6�3ejV��1b-�f�5Y��� ���l��E��b+`��Ŭ*��j��m�[4U��T�ij֚�Q�[I�b��e*�(��F�VѶ�Ś%mV������&�f͉T�e�ʓMK-&�T�m�A��b�h�[%Z0�Dm�emU[Q��;-�V4���  1���L=qWm�(�C��]EV�V������u��T����ٶխу���*�l�U�Dݳ�c��Sgk*Tڑ�m5�2ٴ�^  ׁ��ְ-�����ZQ���E(��z㢊(��(�CQG@�;�ǼQEh �����(��(��{ux
�(��E��ۼQEQGn�Ի�Ѫڍcm�%�+[kVǀ c� ,�&��T�W;M�F���pR���n��� �(��s�qA�����-���pP�P������ۭu��VE��%-V���1Bh�   �����)�l;�;���u���w�t-��k�mv��t]�v���ku�u]��u��۸��4uv�w]�қY��Uuոwf�i��n�ӱ@W+�V��X
kJ-�I(�f�   Y{{:�K���t�me:U.廪���Zݧ])�:����Ki�nٹ��kQӗ;�ݳn�kv�L���5m����.٥�;�hVtn�.�(kuIT��,�J�2�a�   /Q׻��[��ݠ�lh9��ml��s�wn��i��n�(��5ۥ�Mla�w5t���+����뮻��h\v��ݵ)�7vX��[`�6ɓlJVmmx   ��k{;[u( V㲻�aLvЫ�qZӥWj%;�Pw`�w
�T�]�w�-%���YGI�u-�[R��K.n:���ͫ�3a�M���V����  3�ٴ�n��T���u����:�5N�@m(�P[PwqR��]�j��ۚUi�wt8�]Qn���ݍ]��i��ʧM�u*��ٶȊ[-���^  z]��ZVk�;�ڮ�ڶ�Ӏ�������].�9��:kGn���]��J�Eݵ�49iwZv�wnwmim�+w�SF�6�7]��N��m4$�a�N��d�2�mo  �]=:���+wP���9�Aչ��m� w%�7wWM;��M�:g:�v���UڳSU�Peh�Q˭u�/ D�*RP Oh�JJ�HF�M�mP1  S�A*T   5Od4ԩI  RD�UJ  �&��[$dH�j�«��'�\�R8P�8{�u߿���Z��;��Wz�1WB��h��+��* ��Q`QE<?}��z�}u����u�3]���Pz�SB�*V�x�<򬬩�i):u(�Ӂ�����#��1D��ui"�U�2Rh4tP����)0����Ӗ�*�\�PȢ��/p�րf*x͋:h�k�2M	�A�u`���`�*�F�:���*�-rmYR���NI髵�~� ��KSN�K沛L�z��a���,S��zв��G�O5�Zȭ�]�X�*X�CSB�S	fVN�[y4���a�U[W��`!N�F����ݭ!�3��$`�D��I*@,;����E�ջׂ�2mZwbz���(+c7q#��k��{�����P�n���k;�b�Qb�TP$��hS��m����vU�� �*�k��DpT#.)�1�H�<�]�p۴	qJ��+jY�t�D���L���4�Ӧ�P������H�A���֜tt2���8�'Y�+��Nvӻku8S�U�HF�n���Ԏ��+D�V��a��K �����
!��z5�d��Y�q����-LN�˚[ueEc�`�v[	ͽ��J�t]�6���	�ۏB�q�kJ&9�Y�Y-�ǻ���o�I+D	0�6��Y���;I52��Y�$�ߘP]�Y�pڰ��հ�J��Z�I	��ŷ�C�����E�kQ&��˰��x�V�5�(ւ�ʱ�^Q������h�h�3k`�]��R�St�f�n�*�f��CN7��(�iU�&����*���5��p�7�
Uq^E3�*�IBH% �@���R�E`���	[��ժ�kWj��ie��d^)u5Vլ����i�sM��Gz�\�ۼ��U�c���U�S8��;ҶPhoҰ�)L�a��f�j]n,��p�D��V��Mf�.B�S��x1����~����ěl��i;�f{.��Y���K�1���f�WCi��67X�(����-�:��fL���UC��5vwi4�ҫF�8��m���Pe���B-��Z�lT�jV�^l�y��%K5-�Q�M��X�f<��7��8K5x^l��e�ՠ(�=ͻ�c�����ò���]�� �!@�S�4�2 �@*[�)�i�QS�բ��vѭ���(mчt�z&��@਱V�Z�͝&��d���n�t���wow
S̴�kB�v��j {5�<+awB��ީ�e�A �����{1����7,@Vj��Gf	I�G�:Y b��"�:�gQ��T1���Xv�^B��Si�t�MZՒ��f��ϥ+�Ɇ^D�6S;$�*�O&le��
%���f�V�5��n�¸4�P��tVv����եbVcP���hm��M[ۂQ�h�Vp�,�q��퍹���x�jV�u�&��o��Mb�
Y@�AĦ�]�ǆ&� �tpn�P��%�,,۬.]��
ĭ���nC-ei�j�+(��3CdBv��蛲��Ä-[VT�v���o�b�XҚm̨�#��h��Ale�ڼJ���0K�En\�B�dl�ne'�h����^Zۖ&��,�$	�!�%�DZ2<{�Vm`jh�� Y4h��Q�ź�'n�[,��H+zL�.夎��C��0��x�<�xC)Y�S�7�g]��n��d��Ʊ�fXY�`�5y�N�],������>l�l�V�y 5$��[[�`S����DUȀ�U�3FMJ�o/(�l6i͒�ʸwKU�T��#����(n ����D�J�CW�T�4Ӊ������-��M����Z��ɪ�%��\7q���3r�r!y��mY$�IWVj��BO���n�����e6���Ҳ��׳.��2�\��J�,V<R��`����.eԳ1Yse��SfR��䰙�>!jÍ�3.S2��Y��%G+V8���e@��T��k"y���/.V�%��0��l
�լ�M(N�è�¸�d�6]�+b�a�۬��y�+�<I�x�k2X�+4�lit�L�@��݊ѵf�-]�O�0�n�F�&�C�5@�
Kۼ,nԴ`��é�nPj��sqQ�*�B�Ll4}+]BƤB��^{��TXeˋ5��`�����̂���M��f�hqXܺ���y�XYb�B�N����Ѽ�)b���J��X��]��:�����9N��
�R#�h�D-���&S{�H��S��Q#IC$5��.�L�ST�L�i��iV��x��9u��,,ZJx����0��	v�7��!�a�y���P3$[H����J� �h�Y���^�
\�:)Ax2T4�8 FQ��P�I���h��{IY/d����!��dqSQC�$��(�v�.�hd�Ǻ�ƪ�b�CU�ZEyL��t�8E|��A;(1�r�`
7��	(�	KC;�7GඣET7�te�J��ޑ+r�!A��q@�T�+c[�����!�D�wwQ0]B�T��w-^TŐe��o ��Kb)X[��eD���
��]��Ȓ�GFc²��pQ�r�fH 	���Lܢr�l30$/��1�Y�Z�VB�4��[u�bE� 휧��P3Uַ�h�w$��X�E�"*�$��j�O,Iwd9&�+i���n�ݲŔ�]��-����n*K0�m0ڂ�+ZЛ�Fe[?'e��5kD��o9�!�^M�DL5�8];W��e9M�G��R���56�4o(f��2#�Ħ���=z���crjԊ��˸/u�-` %��Y�⧻MG"t��̗WM��W[F��
��W���)U޽��m]���kfՓoʥ�m�6�fQaʂ�/VK���\��cɪ�sN0��o&��)���L��A����
�ڏU��M��%L��kr�X�.E�0�
�����K@%r��QxC�Sp3YG�74Di�:�GC@x��Tڥz���"bE�ok^�����YN�K���T&���U�VV���6��Ҟ�lZMs0��I�r���(�.ֺ�q�Z�3\Վ�75�C] 5Q�-8��!|1VK
��U�U�K$y��ӧ�1l6+��wh5�4�Y*�1:�x����Z#j�0�N3���J�.�6�Gh��m&*V*@��:��<̛&#�ѻ{F��v��m�RzÛ����gM]-���)cm֚�Kŵ��=�����X4����fM�6,��h�Oq���֦���I�0���̓9,��ҡMS�a��X��te*�n�Z�h՝�j�jҁ�������f� �[�����U�l�I��Ovh׻%� I�F��<XZ.T�$lH��/�i�a���Ta�fɎ��ț[��X+,�[EOsW>�wBE�4��XX�m��k@��x�ͺ7ɪ�ܐS�ur��}���k��F�Yp|��%]�%�=R�V��0e�[���2������.#6�렌�W�Iۋ3J�r�̤�j�0��K�#*|�ZVHʃZ72���p�A]�7I1��*�Ĕ�Y,��@�hd"��U�V�)k�vڬ�Y�F�\l;��D�h��h��䁠5�s+���A�����"�.�WoD� >�:��$�N�J�bÔ�.#W�3]ܛ��"�N ��N���BP�*άN�]5%��-Q#FZD曡��܊Um-v�7S	�j�Y��mRʥf��x���5e�z�pMj�<NXթ��7EMB������Z ��(�S�Z�X��-C�c@�u`5[���1�n�J �t��j�F3��,��Ce-��8���4��ËfB��(+�q�ɢ1�nһ�H8D�:��ʗ
E5h�x���W{�٩Xjj�SX���`=Rh�Fk"�a�f]�B�V�,���(z��&hG0�, x�V�U�*b4+ej�+Uh�m5f��1I�D�2Fu�CSC��/
P��,�6��T��A�x+sp��l�N���DH�M`8�8ڽ��
��R pd̷N�;5 bQ��f�Fe!�qk�g^�k�ku\�����L�4�Y�uo��uz�:�q`�P� g )JVZ�vU��{J�`j؀e�+ƚ�)�y�6��j��`�,�c�%��[�`I*g]-Qi�mK,�+���5g/z ;�n+���DrM-�z���	�X6܋vKZo�H`RM���Zbq�冂&�4��`s=�Ι�}��eGW��n�	+ZT�x�˦r^��񛭁�[�F��Un���J��Y���BM��x(�"��N�˄Vاys�a*�W+v+�8(�G��n�S��y�-yv�@ xV���J�;����²#ZcW���#i]��!�#,�$������C���eG��7fRJz�'BE�B��)��M���L۰Eh�ݕ�"(iJͨ T	jKd���V�+U���(�r�� �f#f�R �J92�Dwr`Wb��j�v�Emm'q��q0�S:b��n�8EK���[� ȌyRCB���n�Ĭh��+��P�67.Pf|
�[���!ؠEC3�q��JD�4���M�j�=Xi<���ʵ4���l��8d�8�z%�t�}���41�:���j�X[%��ņ���D�E�$�+j�͈���N�Yqm���0����I
��� "�޻�O�T�����W7/mh,��j�ԛ/
r��v������A���@ek�A��
ܵx�16.M��eּ����抔�����Wq���X̸)%A�Z+ӷj�jSz�U��]��[�1Ӕ�&��0�76�4�*si�1CCd�!�扛NM��Dgrlk6Lz��,8.����#֚�.�7y�^j���L���Gh��i�4ݣ�$��e;7�u�`��v�4������깚\M�jһ7�M#i���Mm9�b� ��"��Z�w S-�tt3�pX�@T���+
���p��ͥ�{�=���bCz���ڹF�4]RrV]e�HJ�h���%+03Ch�x�U���ar� '�`Z�h�˨CaD�[�b��4��[z2��Ǥ7���ڊ���eZ��1Ivm0`slKͼE���P�r���(��RS��`5S �VfkA�(*Z�	��e[xXB:��'�����`�f@���]��U�S.��]K_*�E�PK�2fhC�V�0Vk���Z�,�d�#�f@��u5T��Y�ۺ�Gh�f�9f^�YtΫ�KT+];�IN��cn㫭���I̽QC�ѿX�M%[0��wwkt`X.����*4���=��a6���i�d� 9�Ck {����5���Y��3��|�j���;�C#���Z�ZU��m�Q�y����� mڴ>�-|�;oRV���+4ٽ��L���[A=[�� ��yu��˨�V�없*����нS�t�4��P�k2,���vr�Z���������(nm����էT�$�o��û)������B��^�ǲ�Ü��PI�Z�L�2ɨ�b�mn�y�����S�,<(�hw�n�smUc�2�`ڴ(���9V�xԠa��u7w6j��c�p-V�vh%��#����k%�������S��伡���Wh�NQ)[�SB��$]n�	�V��܇�y���i*����c�0,�V�)�[Z���@�"!ࡍ�r��N�c���ݷ�C��k-�wt�m�lj�ڽ����[4FD�ڸd�i
�c�68�yh���"��kv�n=�Ie��O�ay���մP��EFL�˴iV�G��zF����5]h ��a���jBܭv-@��C�?���dݦ���Q��TmF�Ua�Mu�`Ֆk@RZu�u0���El�D]�*���Z6#�oL�U�a��X5�+F:�ij*(A�&�թL j�)f�yqE�7\�h�Yp�Ms;M
���'�yD��Y#,,�񜻦ͨ���hk�䱘6��"�hGzr��IN�𯖋���RY�b�L����in���ӛ�8q���p���m�.�9K���Fu �j�[dm��+8�kWH�'�ݻ�M�JVF��Z&a#��۴�L֔�{/I3*��	��H� ~SC&��6��B�* �J}j�Ykm�U܂�Bt�e�J�m�������*��zZFd�m�{+q�P*Ȣa���ОR�Ys#�spk�N^��ѹ�d"����p�.3���|�v=�+��.�;�k�`-�
d���/Ch��*�����b��2���fޝ���V�X���p%W�uZ-��J����q0N"��fi�B��
dօ���&	{I�C$����W���f��5E�B��x��n�)���6�a�q���ǰI7X�[�p	��˱��P65w�IR��[����lf^
���#E��3a+:�(%\[�ޖ4�!������_��e�t�֠f��F��$rYu{ w�$�qLltyj6��3E�e�$�4*ɢ9���ԥ@���U�R��\��b��V�[��q`�( UIb�̭����qS����̢c̙F�L<�L.ft�r[�&���BՇa]d�U���Pn]2�՚ ץ��H�7[�S;3c  +<:(��l��;�@��ж
 ����c�6.�P��݌cu�h���X�ʶ&���U��(l.H�C2,Y6*��:�֤R�Rh���
5.��"se�M��8��fͶ��q�cE>���iжj�`%�׉PHUk��'B�B-j�����ğۋ
�Z�,�B���e�^l�3t��Y�Y�b���&'���3e��!���
;�Z�H��(q!X��;N�x*���U�VK0���R��đQC�3��g�e6\U����5"�T����!ƹ�n�IKy��gN�������Eu��кw�h6�T��]3LM�kT�cLo��ۏu۶-�;�j��Ŀ�^�8X\�%��K ΖV.��Hv��[]ӷdz@݈^B�����^��;��Z��������](2	�k�ɿn�%UL7���i���m��YsT{����e�L�f���
�1�nd�+�u���s���iǙ3T�	mK{fgS�����V�xܢ���WN9��2�Մ1ϣIeP����㤱�Zm�T��HO�^��9��|hs�U{3E�׻Vv|��L���b�;�n-�Z��oqId]��5�v�i�fN�jt��n�
�yB��f�{���������b�x�t��[�pgn|���Vo�BH��b͸y+줋y�P�*+�����v*��R�Ԯ�:d�����u����mrE�@өN˻x&�W!P�Y�a^�J��Z���E����;�ۺ\�b�lW�ʦ'b�4���Br��	�-%�x50���K�y�W��Q�Gog�q[���y�X��v�0�Dq��EM���]Z���(K5��|V�_Yc[bu�4��t̘��µ�D&e,�Sd�-:)".�,�d;���v�o2X�޽zwd����u��7.�������=��Qs��(�:��=�ХN��
�Z��-
���rd(r�,i�{�{đVe��hS�h.��r�L�`D����dD��=	P�'V���,j�OByD#�ɩ0�v�h����E�h�7�M{�,A;l�ċ��x�vf�PS�H��t^mW̢#Ӳ��d���n��2񘲻�Z5�]�l�omI�
ˊ�!��&�'���.wjm�����F��`�T�7�" F���e�$T؆�z:L�up �y@�[����=���B󹭈qVp5���h�c����Ղ�y��e��c�K���;�B(;;�Fq�����|�@�>�Fؗ 06ȩ���a�l�c�`��V�`Gۑ�}�+\��8���c���t���Q��7J'�:�
��tg��=r���bzU�T�YVH���'�L'riI|��ܺ��WN�g9��<`a�/䚥�t�(1�P�Z�Y6�V��@]n���9Ո
�xm%;���L�m�=W��pdZ��kod��V����1۝O��n��/o7��ͅIN�o�p�@�©A����)mhv3W w�T"#�3�YR'�H���Ո�Tj:���Qn
pTr�g92�Z�fLU[�;�`t��r/JÍNXX�LDu��/�+w�:��0)ۄؖj�(gswɝ�6�y!�W#�7ܪ.��qj� h�/>�hX��Fu�J�ٶs!����P�n����u/�Zx�u5X���ǣ�8��[������p]���j�Bnǲ^� ���0�FkqE
J�;�����[������Q�ˤn�'p�_K�|C�_���Ef�y��-$��r�6XǉE��5͌�&�ԇ�g>B��)3��E��n�m���5z�<�o�C[�Npx�_7G�I4��2�niT�μ+�
�f��k�@H,�N��S���7�ֺ��(�0{���f�3+��t�h���ff	�j�6F��,���T9<�ߚg�|4�fS%����C~'�v�#n*�T�-Zo��T)�ޏ-u������ӎ��b��t�F���9�SO���o�m>���gP$CÙ+k�ڑ#>�Y
�H���A��9���D�\�WQAG��d<tmV%;�Eð�z�y�o�)p~���)2���2���l��+�ˮ�YK R޴�Ŧr�87��l�E��.dY�W-�J�0v�{}7mG67���ۓ�;�[Gf��!.�ն6���a��	����Z��@���/oR�њ��SN2�{��P+/!�ڮ+o�V�$��.a㛉�qv�[ۻ��X�ۻ��N�0�O5n�#j�v�	WA�ɵEO���y��y��fib7a�<���n��,���צ,�GY�vԗ��9��xWj�j��v�a���m�����͐l�n.ous��8��k%���E9�5�%���5-T�j+i�D�H���Y*�6{��w$�GM�g�%��H���^`޷2��\]F[��,]�R�S:�6w\z�]�7rt2�S!���8�(�S�cH��Je�"U�B SY}���5k�35���N�Tzwb��vsf$�R�g9�c,s+�X�k�:�Z��-	x�X6�jwt��7qtaQ�T�v"gj�i͸Mo6�D��/8�%n�1WX|ľ\�ĥ�jI��ȑ�k��1�CO\J=O�H�)�<x� )�n�Fﳫ-�"�]Y39#�)[{{�jG/�T�m���x�މ��Έz!��!V���6,U۔r�y�[S
�pi?O���ԝX�bõ�V<���eNs#6���h^�=�t7&�u}K3D�K{���ǭ�@�
7n�PePy��Q�Q�ƟtS^3B�ﶍ����qG۹��f���J��Λ*�r�?�K���4!�e��������A��3~{�T����S0�U:}ͦ9G�ڨV르0i��T1vN�T�t�]֛�����T��2��{��Ҟݡ'Q�ehX%�Ԏ�Qts.ͥ��&WUw+Z*Åhu�<�ka�=Gk4��k��ؑ�yIp�QtK�^ָ����)wF��D[E5�3�vs�no9�-<`�1˛�k�y��vNTɛ��ԣ�W�J��ܚڪ�S�n�U�;�N��鏆UJe�{���~�k]T�o�$-ġ:�-ک���r���,���*�M���l��ڏw:��=����ZH6��p�}Iu�A�;Lɷ�_\Zjs��1D=�6�H{����%��""ATG�Z��'Q[��Q��@Y��]�]UG�m�7kX��(%Y�giQf�<y�0hp�s]��Y׊��-d�}
��PG�gRK�*Ǔn:�Ս�og��Zw*��H���D��^�
�5]ǇM#,WrGyݣ	r�ZƘ�fc�����v�6�b��V�EEf�S ����e��S�K��+l��n>R��P���u�r�V��o!��v�2:4("�Uق�{&r��i������x��3���Q�����\�z��ͥ6��vԘU���f��V��{6T	R��c+��M#羼��<�Û��,�zP�X������s/|��jx0_�u{q&>װo*A�G�֕�*�Wo�[r�t�L^L区��Zb�^��7�L�b�����N��$�N�cE6�\��z����������hȷ�G�f�i'S�ޏ�NovXAٜ]J8lF��6j�5�<.u���.�\�%$�g۝�f��:�H�bvb�k\�/��$�R�7�1J�%S{�B��^;�C2�[��sx�m+W"ѥ������Wy����I�Gh��jҖ���:Û�*��;����2��r����t����B�\rt	c����	�:]��WDRt�PT�O%Y��!!���^f�4�R�٠���Vv�8�9A׈�rqz9�v"�A7ze�9�p��^8��С�+g1�r\��V��g��s8e�5���/Tqή-�� �l�W��C^&Y�@ԅ=R���H��Wi���5��sT��/P�Ƭ�H���B�a7���.�j��n�+ۜ�r�Q�'	wE�����ض	h�&]����m9�>��	mgU\��U�Ǔ����L1_U�A8:c�7��k"�L�ıخ pJz�l���,M|�ƍ��{םf�9��@G^�y���q䵐֯����adN�׷"*6_fέ���1�LqYٗMXXG��r��R��/�d�*Ru1��	����:.u��rB�߮���.��/Ԥ7"M*���y][uw�)�JWu�d�3X$蕼��Py�yI"�]WN�%�a(�<�4�sZe��*���_[W�]B3�}�|������]1�%N��v.��l@v=�mmlit��W1��)�(Qo(޼;g-��a�ϯ�Yw�+`�Nڎ�M�eD�m%�B|�m� 5ȄhY�u�H"Bvc�_�~�j��>��(-~���+��U�M�<b���^wNO)F+\]�\��,�n�
w{ֺ7�gSuq��6�d��%�X�=��WU$%X�V�i
!�o&ɗ��V�Io�Wy��IǤ���ub�w{V-mtmIJZ;`���8���x�7�6��+P�x�98���Z�zP[b�(NN�<o���> ��]j;�:M�7o����A҉4t����u�,�Tt�u)]��x�[krud�α�E��˫�bZ�\�P̍ou^*3��	���MX�Nt=�0�����wU�*nc92e���Z�9Q�%|V+��y�km�����t5�T���_��a����'�F&j�����cw5I��o;�5���ܠ�\�ƥ�sp���H踧,�T�o �#��WoA��ʳ����J�B6�c�x ���t�s%�E=ٗO@�x��X�����2�v�\^�@���M���1�]ܲ��	�ᶂ��_"gg��O�s"�Zi����v��Śuc��:̶�"�"�v�w*ܘr�J��3�z��@m��Q��� �(�7�����oF�f[u"�$AtnJӻ���4��a��ㆉ�:�6s�&���ɒ�����-�֚ЇT��j�Z��o�ؼ��f�"���;��X��z��L�{K����X~�!t����ѫ����vCr�`��޳K�;�U&I=��A%�,=�^�5\�A�s����;Yi뮖^���:�ϗC���峥BTm飌P�yʚ��XW׊�Ħ�~��i�)Ѕ�o)C÷)��y�[��������7vWkJ�\
�X�ۑdp��|�:�Y��9��]��h,Ӭ]CeaV8����t�=\R]��7ͱ{�y��F�ȊF>�֡M�sM��1�t*IJ!�{2ݺ��"��ARKx���o�W��Zp�s��"��%����z30$m��.��	fC��/�w;����|KS#��e��������;e��h��f�vCnV�J�U�ԛ��-Q%�/�ܗ�^���6�;�̔��'Z�v�=w�
�N����㯞k�s	�f���])|�
�:��!J�<A����E�`B[�\e��'�����
�*��whV,
n���JZ#jU��. �e���f���.��Kr��y��&K]{����E�AE4QT�aя%�K1� �ɀfpv[N�������6�D�KUJH� b�*��c4�
W)件���u���Kk8�ظt
�E��]�����XA��YX*��  9�)�D���)���L:���
c��w]����Eʹxݙ�A!�{�7])n�=V6zq��D,Gڞh�����	6��= �3''��٘_7���pJ+ISktG]��#Z4[�y���Y�!�(Z���ac�j��;�t�j�P68!>��>Go9$����+V7�hޕ���S��8-ʮF�f��&IHb�xVL* 'L�R��r��bIh\���f��g5�l�}WM%d؝R6IW����N�P��z�m]����gA�r�0��n����t��j�:���*��:���.���v.[:ɹp�9�3iL����q�b�H������.z&ҽ�Z#�jtyWW����\�.Mr�:��[	�9��m��P�B��ə���G`�G���&�{��.WҍM�f�w�0u{G�&a���Fd�[Mgw�D��1\)3���<ܛ©��C'\�]նB0c�Wnd�6��R�9To��B}���$X�y�HN���\�j�?(�o�F땬�HUy�v����EH��-��k���^��#�g7�����2��D^@��������Ǹ��Xr�b�͚��b��:���3&�+��������Ŏ�������Qfv����7;( ���\mo&m�v)F�!��}��}��͖zU�)��Tl����,�c�jeݍ5m�wם�+-�W��M.��+�8k�#Bܭ�r��n�����q����"̚�Ί��ݕ���l#u��*���V�t	�0#�� }d���B��f�5�ۗk˴,T[��J.!�\���ӛ[��|p-쨄6�nd�X�&M�/En�wy>F4t�-���Z��F��F*�a�U�@����#َ�Cf��v3+�Z�t�Gެ�/��1v�V�`�0��J�;�\+loM��Ko	�ԧ%,ҘA%�h�\^9�X:)����pq9U�XͩN1�ږl�1=�xV=ؘ�8_b9$���%�ɯx�=���M\�"w7v�:�>�9YK��ȫ�5D�ܲ%̑��7\#BM%�V��䕗�o{L������Iۋ�{k���79�ȶ,��F���;r��vMOu���E��[1P��	�t�� ��r�pn-��e�O7bW��سѓ	�9MK[��h�2M2�eA����	���3��hU���x�l���pf�������2�>s����n�3����j�1�ƃ��ݱ��Q�'ơ!r��:QY�"T�̱�y ǡnTf�eK$r��z[�+qϖ�/��+�z�<�x(ic�Y��W��n�L��pP��w$�.�M=d�NV��D�|��]6Q�Ð�2C6�YY��D+���ʍN�˪T�i�^�"�{�Ds�v�����*ryq�rV��PH��u} ��+�|�5��jdP�c��_�CR��zFb������HV�$�9,w=j�ʳ��ܚ��eU�b�����L��U���?���|>�~����꯾���ę�|�{P��ݻ;+i[8s2�2*�t65i���- ���ܦ0#�kgN���s�N�So�[�gj�g_;����e�L���'���*ۋi4��d��Yt�됂���n�t���/�;}���y��U�7�Z�
 �_RL�M4��v;'�a�f2��݃7�&�S�Vq�c�J)�0C�{̠�a���&{N���:35����C6ŕ(
����Wb���Y��e�|"�Tb��h��d�W�4�)�	ޭ��"�m�Er�܏k�u��fD�Wz9�U�ң�hIɼ*N����]��%
��y��2@x�j�Oق�`�uٚ�Gܺ�JJ{o&�C�n�zқ�Me/�y�C��*�gwnӭ�x�8�(ݨ���.�WA��4K�6���X�����{��u�/��\����&��66����,��iTy�#�9�]��R�q���
�mHufr"���.,���[4�� Ne��'7�4
5�z�Ѭ\H��t7�q,� �r��J�!��	h#-l��n.��J�����,l�Z1�Ѽ�$�oWj�3�����nk�j�'i+&�wWԎ�u������éj-\�څ��pu^!�����g:O���9_j�V����Ǆ]�+C͋����;�Ӯcۛ�O]U�m�.c�����]�EUJ�dz���n�C��g@��q1�����;�t\�KY�駻9���6H!ig��8	i�'�7b�|( ���Q���*@�E�Y�֬�ê�9��[XezDBd�0�z���0`"b$��sM�r�4BE,��ai	�݆��˶�3��Պ*��E���5�Y�:��=��[5]��^�u*��;5|���(�=�}�X�Vof�Xm:MM�i��R�P<�GvBrf�8�So^�.s�� �:̀�����6pQQx/_Ho��tH��GHN�"]j��ƍCY!�W��T�/@T���vK�S4]�{l�K4ͼ�xf��9��!6v��L`����J1��n:�biV�2�Ïw*^���W��<���w�Ye��Y��*�R<�;'��턌�T	m�C�W%	6��6]�^�:�\ͬԚ� ��Ŗ�ύ�N��R���ZȾ�C�k��P�]�ˮ �XE���Z�gu0��AhFJ3��	f� Ƽ��9V��Kf.��@v������b�8`p��V�ʷU�]*A��:����y��G��u�ʶ��4�dӚv�e��I��0�f��՚����t)X��̐��J��e����R��dJ��[2�W|�=����i��r�h�Q�.`O:ɫ��	���dF�u���.�1C�Y����w4�q�Lo2*�@�JۨZ��8�-ۡկ V����G4�7y(a���\ֽ�Q>\�&;�i8 Q��I��q+����ʙV�&�}��+d�=M:�G���!K��_.}YD���:��AU땬�xbP��̌��Ʀ%����y���'lZ��}Z��kJ��@��l�0�WJ%#զ_(3W��Ǹ�<�vn�Q�8���S���{��aX�Ǯ��(b�����Z��D��g^>F�Q�5gt�n��1ZKDzJ�@+Z6�#N>�ϩ'b1�z��f`��~j�\V�T'um��Z�X�w>6�Q���E�Ȳ��!�����t��j`���olǥ[��Pf�nD��ӭ��f %ڦkWc��^����ll_<B�O�/O#.���vV�T-k�����5�0�AM�M�Y�����`����֎�	�e�_no1[J��C��k�+���Rr��<�Dl꼺f��.�6���5.�b�^t2�l[�gs���V�m��ffP&���!�G����,_e����i{E�8i�\\�ߵ���'""�es���nb̴;��U��#<�;�ҤJ��fг`A�w�+�Ni��ܝ�C�uZ�ғ�����+�b�8�D��';#ݻ=���O�|��ׄ�O9V1F�w\�!�h$5�w����{s8�{G���⮣��-1}59*Z�81��ۛ����Vlu|1���&ښ��ۈD9U��t6,���k�Z�`���"�7�f�Y�tu�9wu0��%	T�$�D~��û,>T���Wqd^�xr)"�������TQ�&K׶z��/z�6WU���E��K�0�)���)��n�0m�m;�����@���d�2V!C�����_#r���|N���U,.>�V�;�@7��;N�pgG�sjR���rE�u��gl�4����]����]�׀�ͣ��C˥p��K�b����Wح�Gk{�l��:�Y���@^�[&���V��W�Rt��f%.,���}%�bJ�NDXDOj�d�ԅ3�͖�r�YX+B�St����sO-Md�2�7���/��7��B�x��ѣ�y8�Q�f'�]�Q�X�\�u�� �ٹYsK=�l���pn�[Xڽ���8.��k �t������[�']*�G�Y<W[wyY�XKZu/q*VoF�z�'�3�6�][ޮS*Z������f��R\"��`����JU��+r3 ��<,� ��E1țW�T+7�{�\mK�r0�J<�̊V�ֈ��z6/�P٩�xR��y[YP���VZ=m�@��2�fӕ�P|��]X�YZ5�9jd�T�)�r��X]�Wee����� �
�p�l*��n+mU��Z��#@q�c�u�&Pb���K�Fr��a��t�;�n�C{��0��a���3"o��aJ�͏�*�[�~7ٱH�J���b�۾���aG�U\�
�s_mE��	w3,��2�[��T�*Թ:�ŝ'�栙Ot�w[4(�5�p眭P�nS4�Z6@�mplw:w̹lҁ ���ۧ/[[cu�9�)�=xK,J�!ǴNn��ǆ�y���[5���T8�1��XR�N@u�X��	;mk�jR�W�X�ʮ�U�,A��i��b�˙��5T7�B�ŝ �P}��Ճ$����"�5����2�f+����ˢC��n���z�Nr���{��� �a�kO�֒]��oW]�_^A�9oj`=����jѺ"��ځ��9#1�NmgE�Y��E��{���v�6*]�:�]_&��Tl��n�Hs3uf�����Y�h�v��O.�	T�"qu;�v[�9d��]Z�h�T0I�c����U'w�� �8��xvgwY����f�쿜w�X%�C],�s�Q�Z�nνmN_1���U�}�9��6	��a@ŴSȷ�%�c�6f񷝁�]>��]؇��tkH���ZD��8!2u�*ӗe�Ͳ4�yӘ2�T{�ѹip��P��wGY�ݬ�V㽔���᷏���U�z��Q���ٖ��P�j���%���:	�[F2���^oh��k#؊9	�N'BZ5:�9����F;����Uc=z�h����lV�n��$��g���F��n�fX�%���5aR�w�+�}��JV��p�Z�a'�m�@�u���p4Y�,b13-XΩ�v��]�P��!� ���S¨(�;�j�nK�{N�4xG�9v��)�F�����o"4�W]o`��øo����g!`GX�"�2�1<
���9e�W`��x:+V���{l`R��d�5���X�V�٢�`,݉G b\#��m:a��0i��Ú�l�T�����T�P0Ů��#��(��p����%Z]��k��wf�V^�p�]R���91⫁D�8�����}+�8�ֆ��[ad��U��Κ����+c���u�P�}gVC�N.|��M�5�u������@��/-��7Pe,�k�Q��|��˞�W�w�Ήi�m�QU	��RO�r�(k-��ZI�n޺-��C/q���t)bϐ��sYT~0�F�=v��j���!���Ǐ�P��Qio[� �
�̉t�Cl-���V�d<��w�v�O���S������v��YM�[QU�3��껨����]�>&GΫX�5Y�����[�t��9H��P��M���Xz6��3���Ĭ�v��_q�E�s4�;���6b�A���A�J��P� 8�tj�B�]УP��kowx�6�F�Nv�n.��Yn�h���uŜ���a���Z{�1�`�ޏ��*vp���Q��@T]�]&Ӎ��ݤF����U��6E��9JR��vg��N�f��	G�d�f�'1:���.�-�y��;����q=���\�l�w4kh����n'��t�J�6�-P����J�}�<�x8
�ks�x+�n�d=*[��ovr1�����G1��&�;vљ]դp|Z]{|�P��$�o#u�9��m�4n�t�ܶ���Yri	�g\+��	§v��M͝YÑ{�*����7]&�_R΂�
��3��$�;�ռR���eL��^ln���2L��-6i!�u�w�EǴX��W+���ڃ!��FWP�+�v���(�
�9�q��U����A�1����mr`�R �Vr�.���,�p޽��XC7dk�7h(�%��M؈mC��M* ��@R�ه6�4�o���\f>����ɭ.oV�@t��U!{l��hl$�����v3zY�+ox��tPÐ&�osx�/b�� .pQ��z0lU�͹}����L�{g)�>�[��T5�3v�P����q��/��treC�uх���j�)-)���Ղ��=NdC~ΩӒ�s����B���R�u����R�R�X䋭�4���_7mN7��.��c�gJ/��Xe �f�;Gxuk�gN�����k��P�r���fLK4 !�m��T�9�z����-�T�%_$Q)|c�����ꗏ-����븎�'�bGk��St���NӇf�ʖ�C8�Me�&Ŵ��b������'�k��`�.�4��nƑ[���n�\2�<f4`o����I��n�Z+7f�Z��4�x��\�7o%v,�YЖ�ɴe�}{VA��9���1W��L�5�,Sk�녝���8��R.'E4X��Z3Vm`(͂���/N�i�yƚ�4]MWLܬ%����h���i�o�v��q�UJ��$��P����R��M��Y�����^N��
�܊��g-�j��	J^5/�Ǻ�4Oo ��s���L�b�s�y��Q���>��K�6��Z��T+*��ڔ���e�H�1ٙ��rPEu� YQ����K�����!`;��^��#�&!R�jq�X�e��V�;�.v˽���
毠��RT�N��;췎�B�j=��}�R�#�
�碌f]A������ob�iMj�T�]u��gs�4��5�h�2���
yZ.=E�3g��U [2��z)�PjIWM�*���yga��I�1%v-���`ZS
M��܏uG�w�<ԟp�y��I���]X�[�X�#�t��UۇE*b�8:	DÍ�`h�8~8*,E�P�l@o2h�3D�X�87����%6>ǎ��aIҵ*f���V��ݼo�ւ��ݥ2�A�����,��Δ͟_v�����pV�N��	��3��t�)���)2�J/--X�G�B�d��I3�u�B�sd�0r%w��N�Q7}�8�����,�W%��gb�`s)Fy3G��j�̆���ˌ��:^r���v�+Z��7�	&�����-ݵ�DV���`ng�-|1��Z�ש^���S�^�Z&��N��ݎ�����6�qt�G���p0�,*s)����/N:q66G˴�g�+ї�EQ,��sQa&��V�x�y���Ǭ�s5xLݮ�"���Q�8�ĝp�h�ZѶː�]���vK�M��9�J��Dc�C��[�&��Iv�]WԞS���=��6�6bu]�vc)�7��叆зS6�B%�*��v�<�qu ��R��N������v�t�k� L_n�Q{�3V�mB����j�C��Lɷ7�K��P/_M�xQ�x���)b��&#�[�ۼ���,��x(�����]΀`Κ	6�p��Q{;g#,���������1G*!��p�^#�����/{�0ĠQ���Ӥ�\�q�G�f���]�f���Pφp
��֣��nV�p�#J��BY���1�"ήlm�ȁ1��+�>yl��$�M��Wl��֯��twm|�;{���D*�]��qe �v�TլWnc%[��
핸�3;�'�u�V���O������0jo�oǒ2��V�[��9��|�:E��S(A��-W&�[+B�t����2��D���ac3�=��`���r�璅���M�ZnF�;C���Y]����[բچ�s	�����:��Iʠ��`t5�M�٫�YA��ژr��6{N�qe������mH�4v#�S��0��l4�D����d��8KeJ|�Z��j���*�m
uF���;D#/f�rV�:Pl����IB�?!��u�#2�"���Ydu=���̳Ԇ�p6� o+���v��P�e(��^�n|�u�l�fЦ�eY��d�,P6IuCAKBD�1V�u;���ݦ�g�o��}�#�e���nf��o�n��uڈO*qf-���
b����@�H[P]hwH��[)��b�ѯ��G�b��)���i���psYX�h��:"V���A���s1���J�4(L&�Loء(>#j��u6��1>�t_Io=b�ޝ.Y���^gg'RO�"�@��J�2Ж��k8�o�EB)��m�+]�ǝ���T��.�`if�BI�wZ_V�l��WMQ�X0;��ByK��cN�!��ۃSWp��ǹ��o0,ɩk�*P�yA)�������������>���3l^��U��^�o� R��c�ZcQP��.R��V5���\��~�7�<��OĹ;��ʰl��G���������O|���Z�Ps{������\���o�����|�J�H��ݫ�ھ�����]g5z�3�]6������S}�d�vw4�(�\h��2��{N�i9V�Y.}�ַ��	%Օ9���SC;;o-��ڒ�}�wv�}��W^"�R��l��48%�T��(.{b����qɽh3|n�8S9)���_eB	��9�"G.)f�U�s�OV�KNCԉv��aE�>�V��c�0 �a�[�T�b?,�0*J=�xL��#�Ŝ8�A��;��\.����7�r���K����KhR�x�\�Us�L�+D�b�}�(s�7�.L� j�*�f�x�q]5���:�y����]����ֺ̢��e�K�@@���f�s7/����O��"�c�&S��Wkiq���t�D̂�\���@f.�2�0�M�ӖVJ�� g��\�N:��2�P�*�KP���'ʥ� B�)�ܕ�a��)�sM\�+(�ة�:%y/GS��K��1�Xw��uN�v8�9��Le$���3�Rfl�v��S�j������-˯>~�~��nT�#d�#/3%��v�p�Z�}�'bC{ԫ�/�1����e�w���~���43O����eSPC��LNT�c�$Y�TFf͙�Ae����aY�MfY��1��Vb��QQM�0Y��Y�a�F$T�6a�Q��deUMFYRFT�YcESQ4Y�Y�M�AVNFfFefffTFa��4�C�faFY��9e�FffeTdd��a��aU���ّVYf�VC��d�cfdd��Yc�S�e�fVU��T�YaUd4��Ee�Tff8Y5�D�e�fc�eNY5�f�TSAe�c�d���XfTT�1VFEQTљ�M�c��EQA1EMQQUR�Y�FD�F5RQFAMDNYU�aa�U�fTUEVFVf�gc�~�ν�~����n3�칭��vV�����4}� �}I �a�����^����5�d��e��A�U�j}}��:[_OI�GR��w�rht}�\[|&u�@��9Cf���&��9���B��h��Z��)ިE�4�c���5=
�1�CB}��k�f���k�d�������.��J���joj�:����{/��������rWd]b���3�٨N�Rp�6p�Y�X��ͬ˶�꜎~j�-6|_^_�9�U�L�^�ߪ�ނ��q���7�y)����}"�fu<��g�^5R���Q����,��.�g�S�Vv7ܼ��%6pMz��y��Ǖ��ߌ�8�L������n�\�o�{еd���X[��.u�Z��o�7S��{^��E��jZ�M�(�����=�
5u#ў�n+Ӝ�)����i�(����
aN��O<�ΰ���K��XҙX'Ԡ��QWɅ��N����4�l�P�=;z��a�o}�{�(���GI�V]���� ��Vk2()�Lœt��gљh;+��I�HS��nշ诙)o��EYzu�f�[�(�le6�f���Z��w([\��މ�g�F*�b�8I/2>���\�N�N�t���9y;f{�)ea�K��	�U��!P�9i�0�cWc�S]�U�H+��ۨ.˨7+��VK���}�gE�_�.��ǚ����ל)�j�I�ó�Y��t\1ѐ;]A<�"zxXѓ��5�N\�ɗW=��yMht����v�T��k�1<�D�Z�6_n9V��<�Τ�y�o�����v?j|�:n����r�u�aN\m�.�y������F�v�t���w�Y~k��]<��n��b�b}�M���/s�t[����8L�5+f�U�7cJm�^aK�к������Wt0.��ǴC��r�X?+�Nų~�S�ݕLh'���x3���o=�Ƙ<�h�d�wN�!�ud���b������q�cG7���!�ܷz߹p�'Г���Zu']�n:6���7\	E�1R-��:�����
,}rM\.�"5VZWP֢�d�
�,�Oȸ��v�ڏ.���{��k�P��;��,�ƥje񳹒<Q�m,�8�$S.�(f���	�0�D�L��=cT-�3+#ے�V��:<�"@ONcM�ȴ�����G����徧ݭ��;�s�%cB�Ţ��6qޚ�%n0�{�vk3}3�?;�,S�y
k�jsֹ�-htE�[����٩.�Q���}����Ι��ʯ�b��*2/���U�ή�&���u�4S}��Y����5���vϬf����B�)���圭''�8&���f��W�z�\�O�E7�r�)!7^7.��J'S�����'��YǞJ��$���7��↻�l���m\���3�߻W��(	�s9W�-���ڭ�
U�w��+zl�m�u�gΆ��m5�[��0�g��dZ��~'�E��k��BЩo�q	��l�y��������X�.0��(��G<���E���1w:���:n�/.8��ȾQZ��ot�s�<��b;!w�����+�[��M�=�_�7�z{��;1��TW7Q��8�{T������§tON��x�}gCy�3��Ν#(���C�&+�9�����e�YN��r��g��\nU�{V��WRd��BN�ܣ�|%�Mʙρ�Q�w&Khh��o�Ϲ�g4m4�P=���5�V隅����8LA[�Q+f-�1\1ɨ�v?5�l�����s=g"^�a�����[�Oj!�ï#dN��-s��s}�Ab��u5�8wk�6�!�������)QI�Ȥ޳R�!�tu�Uڦq�Su�������a죩��K���͖�F�p�W8��wN�^��ݔ�B���Vg�����7�B�q����{^���j)<Z�]pyk\Ci,*)��Lf��;�-�^��W�^��~�{j��*�®���6'�g�vÝ�7�t��~�s�9=��@��������tܕ�E�+ny��N�-Zв�y��:rj��|}�o8��Q�~s0���+�{h^��j�tP�u#��C�ic���I�=�;I��f���k}��g%�ōF��q���b���}u��xKN<��p��*��P�:R��@M�KT�����_��ީCw�.�S�@��V�w�I�8P�§; �� 5�ʘ�q׆hn��V��b�j��A'��g6��3�ޒu^G�r�܁Յ��YK_Ό��C	��N�/�(�#:��_,.������o���N�!,H�y8�]Ӂ�2T�z��.�rw�z]�D���&&�!K�I�+zt �`��iou�v�\�U����uTK��DZk-hR��f�r[��oB��Wײ-c�wn7��[gk�h�:&k�+����	;��w��R�
.{�O���������S�1��D��#�z�%�D\�B,���}^Jy�'�_v?ozr��b���<���g1�-�tA�].�^���y�|�j�Po��b}p��=%���Û�I����sלr�K7;��it�޹�����Ld��S�G�Bq9�ި|���l��;�ܪ��!�X�/\��u����kg��s��~1�*�ˠg7���TJ�趺��8m�GXZ��w�Sw:]�:���U��md�t�ջZ���g��(~K��1��׹��m<��,���⼰�g+8!M�_6&��+ϭ�4��V�M�"|����)�h+��SQV@^�=��ŭ���B�_�]v�ܦtN���_j]�=�p�_+��,����9gM47��ƴ��_VD�'u\]��y���Y4W:+
1s���*p���ܽ׵]�������W �e\���e{��pss��{�kr�X7�r���?ENZ���-kBݬ�^�6yFi���5��*exga1�䧍�␘��.3׍�D�*�ʭ&�cO���M� 2�{3���S�^z�X�~*��N�Z��LR���:v9�ټ,u��tiD���C;:5ﳒ�cP9�@k*�:�!P�0vgp4��λ�8֋��֪��UV�k˅�g&��v]@ѹG�U9�yu�gV]L)���|�,%�7+;�a����
��y���η�z�:.���� �I��FR�a6�!=X�-;N
��[�R�;�O{/UP�S�1<�Gt�\�õ��B��[�}i�cUiᮺ8���u�'ȹn�]�Tr�w��1��;(�
UiS�W�֘~L!0{]x�s�LV�TiO;<�z�YpҮ�����&2�q��7 ���d.AB��fM/{�7r���T1]5���]��ՒW��e�x	%�^��U�Tb���H�;"2�mu�1��3tfH�kTK�V���,�pzlmՁ���4�+��	��RԶ��K�6;��]*]6�<Ur���̜JGr}(�͸�q���sp��'��>+zJ܋aMp��[�!M��	SZ�V2�1���F��tE��y`��5�9O,���9��G��6oE(�>1?7�	�M߾M�?Z���dRq��ӿ#�:�����'�t+hfE����q[es�4��Vcc�OA<&S���pw��*�����S�J�|�؅V.�����8�Jƅ'�E�8ٌw���Ⱥ��1�k���Z���d�~B�zf���X\��;��nȻ��r;\���4���;�Ս�ip�U�~����[һٽ*	�y�̿y�K�������}vn����;g�3]ٛH\?A�=W��2�j�U\�Hu�g*۷v��k.!4�.��ۇ������T}��`�-�[6,1n���z�A�ך�'J_8M�C��֛ݹXUxp�U=�vp�f�:]��f�'nV)��	��,K��9�^47R��W�����a8Umi�]�#8q�˱&y}%��^9�/0�f_�z��Х�����}�ɱ�-��x�W��u�+�m�R�Mޠ��ԝ��qY�mn�%;���@��՘RRS��Y�S���{��w�\|�j��p�<�}����yW5�pp�����r�>���
y��`(���K���Z-㰩�Zau�"�xlT%|����;���mэC�"j���Ҫ ���;�]'�����������M��+���/�au�bc��%oT�1\�?-�=�\���,��a�W8�-·[N�뛅M��c��5��Kh���oh�^+�K�����=ϗ����=��طOj�:�6Dơ�J�0f&X��2�Wm��ִ���E�ٌ��}�(NBo5��B�r���F@zF��}����Fq��6{�p�'۴�]糛5��EBp�Ts�Ah���uA���\!qOiZ�����z~�9[�<k2]F��Q��M��>
���ǻT:�������~���(XڞAx���PSoW����|���{j���^AP���9���336�Us�MK⾱���^�6�&>��xc%�g��]���VB�~��o��gBR�ǡa�l�J�CE�J��q��LL1/X��iT�*�*)�֫w�d�dKV�ȹfG�ܛN�*p3b���f�=�s&9m��ھ�݋�������q�&����^��E�����,ٞ��V�iO�%F;,C�ⱺ����R܊.G�	���ڏ��+����RͨO;n5�L��PX*7U�|�(�$;�ߪ<��QO��3���z=������7nc7��<�;S�eꇚs�!G�9޺5�z�����{{;	��z���o�MD�86�T8�o1�}W�ܩq��r��7�\t�bo���8O��j�ĩ�v��$pW'�u�t4lHz�	�Q.x.��B�{[�����i<�oT��yڝ����[G�1�0;X�Y��_\�A$C@�O;���7='K�ɹ��OK���/�;!��
�����Y��7�3�K��79h	�=�e,�S��坞v�j��Ry�቎c�C]�*h�t���c��!�Z2w[��;��]e���}/��X'�r_^n�(V��-ג	KU��+6�qHxrKFϗ��-�������n�j<z����:��ڍ��ݗ��mu�;�m76�\�*���M��kӶ�j�n�tF�q�9���4�ѭI;T[������� ��1.kf���Ϻ��k���59s�LAz�/g׃�����.�Њ̈́�r2��{Cl%�Qu����9�ڎ�B/4lt{<��UQ�9c��w�*�l�7���wWEf�=��v�3�в)(YU�;�\>2��С�n�Ʃ,�7<�������$Q)�����_���fz���5<���QyWУYӱ��e�ٴ�J�vy�Oo�jb�{�}�HM��-�6��F,9=�Qt�Mq��[�<��H[���V?O:����kZ�x�q��睽}"��;p�+��m�8�(/�=�}�Pf�Ö�����&��k@�ꪬg*.bm6�o^�Z��S�y����Yg'����u��Lvse:w62/���\sI׭��Ok�S�'��/��)�s�e�R�~��Nz�9!��Ҁ�=ns�5MOn��ѝ�Bj��Y֛u�t4nT*��Q.yǧ�>�on��%r�U®]���{,��T*���s��5�ʯz]���	P���f(�sv��;@�L���sO��fإLm����~כBY&���|�s��i�^kt�=l�e�6����������"|�M�>�-U�1$7��N�΂���j�0Y#�ŧm��[����׌�T-J��oo;OK_Bb1b�ln��Y���Wml��]2�����ui_Db�t�;���*͖�?��8b�1�SKMȢ��ňVWX=�����<$�=���8�!b��4��P:���,d�Ŏ܉|k�w��h�BȊ[�u(݃/E�␫'��V;13�4����.��sHN�ɢY:��ΦEe&	ab��MX�X���΁e�(���=�K|v9�k�Ct�,��2l�ʆ�-FX��w�5��ZP��<M��*�*����#�D*��U|4�Z`�.�ٝŋg.��X��\Bbv��bYj��Q�9]ݣY�t�V�u�k�>�}��L3�^>�kn�#V�WwD󤛋N(T��[v���w�.%:gZ���3u�3o�Ցv�WX%�J74u]$'py[��e��:ո�F`�rթ|�v7�tuyO7U=X���K���AhQ�r��fA�}#ܬ�G$g�N\���bQ"�u2�4�_p��m3[�a�r�L�'�W�|������cr��|�a��[:�wU-iB@\�c}����[���*�<�W^�6�7��r��w1MҎ�F���^l<x�'��ěŶ�|�@�!<I�v�h5գ�]�+l�^!�*�b�����N0�N�]ҬN����9V)��)h9�i�aߖ�ؾ�*
X���5f�EJ�Xy�ݲ�oU�k&�I�{�el����5Hι���+����CN�
쳹8��8C��PI�i�-�l�c_j�A<���fcE����]El5�X5)����Xp��g)q�
�x��ճ����FڮYe��}'̝7�Sw ���n�Y�."���Τu����N���V/��o��`�_9�)�i�ƨ{g-���G��.�0>���)�E\ թ���A}�R�`��+��O�)�x�F���o7q��Ƚ��둜�Z��^�ZnV�b�%b�q)�[���0AW+$Ԁ|u����x���p��|��Ճ�Ќш�8L�c��`F�\��ķp����$�648�/�ۖ�'t�\Gƕ�8��1�Szd�����b�
���D�1����i@Z���u��Xv:T�W}wD /+5�������TݷS��vw��]�Z��Yg_ۊ0*<�z�-r���%Nw�#����_*��k��_e�^�I$*��h�]�Ξ�+3�
�N!Ұ�2�&�ofr�)dk׌���S��Ӄ���w�o\�t�w+t�s�W�Z�5|�ц���8-�h�<�ʾ��3�q������
�
  >���jd�l�1�������',"��3,�b�2��',��)�2��r+(��rɢ���&�����0��gp���*�0��*�0�s2���lr�*
*��(�p��lɪ��,��$��(f�0���b�2")����bBb�"����2����(�q �,+"�0�2��3
�""�*(s2*l��H�k1ɬ�+0��J�0�#3',2�h*�r�"�"�"�(����j�(
c*��p��l��,��(�0�*��3$(�����������*����J�"�0��2%��
���$()��&e�j&�`�0¨����f�)�Bh�ƒ����&�32j��)�Ȣ(�&���C�s���w��orp���27�8��LA41���X�lw*�H�"�fb���3(OV.�qh}�v�X��WժGf����-[�֟+�ó�a�N���D�׀i$�򃵫�c1��V�\��A󻅡M-��]��U^}��ɇc��ٳ����m��V��3�I�]\^wQR��S��>F�7un����Vh��~8Em.�;���E?7�'+�������m�����}{�AF�C�D����{�WJ��Z��B{M ;�Ԍ|��z��V��~��z��n�O�9�}�_:˭ce��(���3P�6F���k�����C��56o��{D7�ؐ��ZK���6��ʄ�\l/R���u�~u*�̩�ԇ�N�˾��n�[E��:�ڬ�c9@���T'Ds��N�׹�ǵ�����َ�wWΣu��W.s��vK�ףy�G��W��}��D��ٞ#Z��S��;�ܽ���ߦ��d�y���9n���T,���}��%�s�v��Ar_	;f���hb��J��n`'��F����xdu;b)���i�b� 5���UA�{8;��^4�'CS/l���t;�r�x8j]œA�ũ)_oD/:��z�[)Ny"��t��wl�-VFR������:��OY]�,p��WӾǛ3Q�yU�M55���x���NU��Z����7�7w�DR�<o�H.t�]��&����v���6��(c�k��.�c弯��4Oo��˄�[��iWy		��u��\OmQư�N���,0�;�E�b�bu�R��M���δ��VV��ض�!Y�b�M�i�un�ƗH��a�.|�ZЧ�޻	��[�=�x�,P�X2J�t�Y�9�p,o���yTK���M�y~�}����g!��D<<{X'g�kt[E�I��;!t�W?X#���K�uR��]��I�\�pM�/�#�^֫�W�\���1<�	+z��:�կPZ�,f�s�����f>��\�z�ڸ�n��¨oO��V�ԭ������S�b1���gj�!n!�[��P�Ĕ�)X��äl����f�}�h�H�`}�*6��&z
��9$��	w6�.�{���}�����1�Ԑr�R��� gE��͕��
������C����UA�\U����A(�)��(�:b�2���4ܷ�P�Uڪ�0��ۖN���2sE�������k
K��0�{=�:�����a�������d&�a���!e�>+�w�D��H��
�ɨ���X��n�ј����y�QP�-��h�[��iEò�.�S�^�����Գ�}������Z�WHzd��c�ɜڅﶽ�47����Ӿ���ٸ���t�un�v{���a���)��k�Jʎօ�X�^לj1f�׺/$,u�dS�*	�:�&�py��	^}ҷ�E��X�����ȥ�^O;o^��^�^�+�W�l_z�����<��s����kb�9ʢ:U]�kq�ة�ۉY�Z�Ұ/M�>���^�>�=CJep����D_$)jt��	��z��x��(֗��V��UiY�8�p�������#���pR?]w��y9!�O�ܻ��C~iL�rt�z9}+�5�e�s�̯���wn��R�`�P���"DD!��~�������Ԝ���Oc%�
N��ù�Y�_`�v����W�bn�$:���y.�'^o����\�Q+6��_�������Zi�`�Cݱ˔��(�wgÒs�m���R�u����`�p�k]�
�,�&��1����2�����o�1N��6�=[�ʻ~��>qV2���U�������b�.�*�7{�n�1vZ�w�K�V:�l�e��`y�3���]Um�()�H�/�a�}���ϵ�;�����u��޴���OLÐd�AI�`�A켎���nz;��:����s�{�;��������&���S���y/��y���Hr�����Kΰ�m��O��i�r���H�N{�K�(��pd�AIј��_��w���}��F戨ǟU�޵����==�#�#��Gr}/߱O���ײo}id9f���p��s���ܾ��s�G��M�΂����ΗPP<�o�W���z�;7�>�B<D{G��}b!��{�ތGr�==�}d�#��=�/%=��r/��}id~ݏ%�O�ޗqܿAO�}�A�9לﯵ�[��E<���U_8�=�`��ﶽ�D{��!�~���`�_e�������,��O;��9y)׾�܎G$�ژ��G��1C�c��"$���_�}<��������AԿAOh`�^����y'�z��d/G��r_�b��ܾ�˫���}�;��ܝ����/pv��+��y��=��վ����s�z����כ?C܎��{��y!�ozJ�����	C�����^I����ܯ>ť��C�X;��^F�w!�����C�~�ϻ�\�|�y����kn�w��z#�1�`�������}��R�}��pR���w��~����z<���u/g����?�Zײ&bn�^O�뗩v'�_,��k>��ǽ!!�P�h�h��R�
���A�ߴr
W#�����2��O��g �}�!���}��{�""��j=#G��"f��~ǲ6��y�=�ο}�\Z����G��x���z;���^I�y��K�+��4/�7~�O#�_'�tr]�@���|�r���7�=��z�|�����u�{2�/.�D�>�a��\���d�ksvT���
=����^�Sⷍ_���N�
��wDN��xV��Ռo�W�޹����Yr�\�:(]�B����	.�E������<�;�)K��xx �@_@Muˆ���q��"��9�T]/����$�/��hp���~���;b�������;��2z������������K�+��4������r��������b���l�G���,���H�Ї��w���K�>ߍ�΅�C���>ڇ�|�ΰ#�y;��r<�pR�{��w/����<�����v#�D�V��}��꯶z�Us��d���w~��9�r�m���4���mo���!��%�O�w�S�u.�XjW�9���)]{�ܿ#���o�p�|0˵��<��������>�2_d����/$�f���H�9�7����l5��.��'f`{9/�yHrK��Xh{���g�Z����>W[��g����+��`n]�Hu�p�/<���t�K�7�^���7���nG�ϭ!�>_K���t���7δ��������Rϱ˳��{�ڳ~_z!��=�#��R?C���qԯ.�`n_�ҝ���~���?�ҙ.���z��R�����|�����w��>����{�˄����}�f�����R��" ��wK�����0_��u�'�Ԏ�X����ف�w��>wք��v���.���y<���F�$���w_�x0��h��{?���.��~�R����|�u��<�%�2\��>���#�yI퐻����>^J{�nC����z�<�����O���6o��Z��P�!Bs�ܿIݾ�AԾ���AJ����Q�>?a�2_�%���u��X���:���$w]�}^J]��}zF�|�b��CP�B�=&,z����w��%��<7�)�=���AH���K��^��ܙ/�����}��a�u��_�_����믍z�^���o�w_���Lե��l�Z��$[��z�ڴ���Y	o~A��`[���=E.��P��u�<�*���ws諦��r��2���;�?]���]M��K�c���5�U��S����/{���̸�κ;�ڛG��������?����+����p��=����FI�}��I�]����w	�bPn_�S�hJ!�|���/!��^t�����4�]�ka��o�9',|�bo���X��G�ts���s��.���!�y/py�rW#$�����˯����
�|�Pn_#$�����z7��=��|>������������o���h��x~�@u�O�>���~:�w)�y��w'�؇�Լ���u�`�=�AJ�zo��q����7/��~ͯ�]w�,Z��'b�>��= G�����u�ޙ}���W����Zג��w#ǬN�܏q�j^C�}��:�pZ�B�$�7��AH�3���s}`�ʩ�k���R��0{� �z>Jb4z_oa��zC�~��oϻW�{�t>�B��b�������;��2;��nG���z�pP���K�,�U��3�SI~<�����y��+�_�Uh�A�h仌���4n^K��>�Hy/��o�h_ <��P���b�O����r�FGrn
�oy��~�����=�o5￷��d��(o�7.�'��4����R;��ϴr]�H��5�C��|;旒C����оHn�K�{���u/#��ߝg��k���y�ε����G�2y��tu��r�!�~��NK���~h��;7֞}��Oٽ���?��>���w�^Hy��[�ԛ���[͟s��0���Ϧcg/�V��}��!��#т"e�sXj�n{�pR?]w��~�����r]�A�ߺS%����⼓�oG!��/=�C��}�㟷�5�UVo\�v�w�G�{�B���z4{���NC��f	��������}`rz����&��2C����^^A�qL�ru���P�ל2ֳw쾷����O�"�hb�RɶZI9ノ��S�k�3�W�]�A�e���D���^>
��4�*�jB�j��o_#1���4i�u�:i+=�_ۛ��v��6��>�3ӄ7����1-)>t�*�\���a�z���,|B$�-��gwFl]����#�����=��{߿�MJ���.��~�A���bA켎����:;��z���k��~��>փp���;�y�6z}g�wO�g.�r�~���z#��槂�j�ޗ��C����#��/g��ԏ �������wK�d��<���F+�<����1]��k��}����M
w짶�nr��"�����L���!��s�!쇒w����|��~��;��{���:��u���wo9�K�P=g!�~�� 7'��uo���ߧ>������wN}����zD}�����=w��9y)��!�|���}h�%w�接��~�4<���
y��<���AH��_�NH��/��kS�鬊�����_P��p�=�ǰ{�<��;:�~����w��A��C��=>y�r9<�cܜ���ގ��'{撃p�=��{/��y׽~�$}g�a��v������������	�ť���X;��.���O�9?�;�����?G%�N��[���:<�O$䎣���ܻ���_o��sW��������5���w7�)I�}���^C�z���W�b��w�krC��?=b���w���I�y�yK�;��rG�2{�����������ov�����x����?K�(NozC�}����Д����?u쮥���t���h{����NH}���u��;��<�K�7\�޵����}~�]�����߼�N��
�}��I߿h�������w9)��i���d�������<��]K����}���;����NbnG��s]��w��l��k�y�^y�=��&I�>�qԻ����{ ���п�ܝ��G#�_'�t��Jv��r�_oa��z�a����p�FG}�B�{�#>�{[7��g�Ն�����F�j<"�\��yI�R�Jd�e�rƲp��^Z�
���o�8�_:"�-LP��$(�Tެ�[W��J�����[������e����Լ뽉��3T�#��v�Ή�s)б�J�]���Q�<����E��jY_ns��z,F�{D~��1�",&��G��5/ ����y��dv���M���h�w+��O%߸���9/%��=s���u���y���~��ܭ���K_��=�ɏp��X�h��N)�u.�c����NAB�N��r^A@v��>�r�2;ߺGrrN�}h���$�����b7���=�g�w�J�/f��N�B��{ߑO�Ǣ�p�u�y���w��FK��AޱO'�w=��J���bn
G��7'$?I�;�q��4�K�>������st;�:���*_E���z>�1�<��?����}/�}�܎�9ޗRr�1=���):��{�Y�_`�w�'#�_����~����o~��|�ɺ\hEg�]�k��V8�=�=�=���@Aß�}{#Խ�z9��y�d���~翺B�=���]I��fa�2_���0O��^Gf�W�7?o�>��X�̸2�J���Dp��c�>�=�§a�h7.���<�H}!�?s���_�w��}�/�~�7�#��^}�C���=��_a�2_���u��)�@߆��Q}����D��h���O����;��y��07.��{&�֐�C�vo�>�����yK���?i��{7�:
W�~�i�ћk}C~��~�v��zD@��C��=�=��~��b;���Y+����r�S�q�!��O�֐�G���y/ry�������
w��q\�'ٟTm_}����D{DB��~�)^A�����2����?NK��_e���:�w�t������C�����r9��h�!~���rq��Gp|����S�X��z�����R���oz�{/g:��ܯ$��^t�����9/���ܾ�˫���}�;��ܝ��<�.K�����k�ץ^��UwS�ȟ]�F�/�A�t���l�5�V�u ��I�3^�rۖ��oK��ƞ�%ΐ���A�q]��7������k�fWF�&��5�I�SY\��=Y]�j����k_��I�C:��.�7��%U+r��_��M��kV�O3����=�ޘ�c��i��]�Ho������4%����W�y�y���+���Z_�b�w/����@�C��<����3�������?o�������?C�<�!�u/�v��+��y������z9.�;7���g ��4%�������^��.�%y��KC��C�;�q�Fi���\�]B�A�[����A}Gލ�LVN��NC��Լ���оA�;}�G �r7��q�>��!�>�A�1��/���u���;�ܾ���oE���^���=ߟy���QØ�?�$:3�cs��p���<��䜇����Ի��z�B��pv��O#�_'�tr]�@���|�r���kʐ�>Q���}�/�X��W���DH���oν��C�����G���-��{��J�>x�p=y�K�){b�%��^h����Ӹ��{�}ξ=���5�!F���0{�[����^K�p|��<��}���_{��j��r�Լ�]c�_'#���J���%����#��S�>UB^Y�����5^���I�a�u#��ϴr]�H�w����n_�����~:ߝ�{��r^��f�O�Ի����}���=uW}�[��5��5���ɺ��>O�wR�!�x>C�?NG{�Jd����h��/$���<�w�<��>���;旒<��s�K�y	ۘ�K���r}����1�特���r���̯�������s�M�R�ݦ�>����`�%ߘ���2]���h��P����?[��ϭ!�>_K��y�jW�]{�#��'��$;�����oVwUk���=A��%!���p����R}���9/�r�f��^~��o�)��N�����]K����}��h�`����n�wL�NP�HG�X��f�l��~`5`�p*]�o(�*�tk9&����Q����[1 z�ꆖ6���s�v�xg3(	p�3c���o�q���	�p-�n<�]΍�˂Y�� �ވV�F���$��&ڝX�z�`��=���Ǩ��C-!���{ވR�X�N�'wߞ���������wK���ra����~�qܟF�w9���S��ܿC����B{�;�5��]z�.KѮg�w��^�+���X���]��/#�w��
W�{�|�u��;�%�2^��na�{ш�^G]�}d.��=���N�֍�r/���>��6*�uUmn}Fn���C�.4/P�����Or�'w���<��y�����|��d�_a�2_�%�X��_�þ���u��H�;漶jM9w���9v��E��{��{�������<y֏�rW��:�����4�K��o�S�{/|��AH��z���2��ܙ/���b�_e�T��j6�E���_}_F�7�z=#ޑ��=ۅ���>�/a�O<ϥr2O��rrW�\��;���|�Pn_ ���BP�[���y�z��d�%q�ߴ����ܕ��ǀ��p���O�c��\��X 7=���.���!�y/pw��FI���7+�_oO!�'{撃r�'g�Д>C�w�w*��k�ׯ9��ޱ��y��zF���>š��ӬNH}�����MXy��w'�'�y{�H�I���9+�����w�o:��_������<}���'�8��|O�R�-lfʊ����5{;ڧX���s�5�+�67�ϯ�yX�iX�vf��lVJ���P�r��r��=]�o-d9IsY�B��}��u<��ޗQy�E`|�f�L����c�,�ۛKiR0��Ěq+h���g�clM�j�v�IE]"ӧk8ǰ��+E�h�,n����lL�CI��H�o8�0=j�>�'UD�oҞ�YpM*�2WP9�WyIv�`���V�鲲���S[�h�g�H�#��R\��[�������k�c5F���:�ӽ}ն̩�-+d���D���w��#�]X3�����h=�woX*���+R���ي��E}��Qī��'obwWc]=yq�ov�(31�7I ��*#o����\v=�L'^9�U�=ܝ��d۫=�ƫ��(^��5��ä�k ��MKk&^��cT�G��e8;@g+�3��eߊK>3M�L��y'n�G�Q���*t;՚\�k����I�ֻ��&�Q�	���b����%�0���+Ripq�&N�OzL�*�+�P{�#�ku}'6��]2վ�n��RL�[l4���k��쾊�x6v�����4�v���M僸a���,.M�!� y�d]}"�����qӃ"�U�лqn}|ztBj6�'��ұ���E��w>
.�X�v���t��{�:�5ad�u��&�������R"���qV��9uC��|�c�ZK�R��+�:cY��J�[Q,4�lRJK4�{ύ�X��j5��|��N�^L��1U�P6���Z����ArZ���]`9)��`��<K9��s{���)���J���6B��2M�[r�IZ	�AƵ܎��<�j��M��Tz��6Ri WƲ�h��5���m���}hB���R[�I�:���,W1Q�t��o�H+f�T�3�:��
w�eg�T� 4e��?z&2�+��64���mEt�R��U�1��S�+�	0h�:u�(q��r�휂�;Of�F�L��f��9nɖ#�*�͝�m�AQ�31� ���\�S����Z��D&� p�A���֮���k�m�gIx�jB4*(�+r�K���z�u���PDΥ3N��G/���XE1Gq����I�wuq`(vݩ��bF�S�ǁsU�M5yJ=����)����������r3�~�6�G�<
'�D2��Q��,	�L3'h�����T<��u�u�E	���񕽻���-2Jz.l�������)y3�b��]#��-��#�8Sw�����ͧ��+���m%]����Nd��q�B,��ݩV�F�!6]5fj�b�`!Mv-��|~�z�K���0N�ޚL�C]������s��lۿ�N��.:/E�Fc7Y��WaT]')-�]�D׻c�+��T����΂��.6G_<�쪈��x!P���T>�Y�ayY��=�w�t'k�N�V��\���z��cS��n$N�j�f4N2�{��j�y2�w�#[�f�I��}�2�n�&�a��=��b��C۰�&�]T�ݡv�.��/4hN����"kR��]Sw�G�6��9Nt��2i*3#3
�'1�
Z"��
&��b� �i���j�������j�Ȉ��3h�f��j�X"�h�
 ��3(�ʢ"bI��"�Z��*"��*�)�*���H�����h���"�"��b��%�&�Ɗ�h�(����h��b"��B(������2Ɖ�"�
&���',�����
���3"
��J��j�"�"�f�ZZJ�(����)�b��Z&*J���
�
�,ji�� ʊj��",b�
j��"�)*��,�	��*�f�i"$����������0r�(�"H�JX�i���
hP��
> :�y�3ڌͥV��JA��=s��"|�Ee*�	���u�՛�)���#i�ݽRC؅-��틨4�(m��/�������rؐ�+����*'9W��p9��&�܊o���HM깶��6�jq�׸��YZ&=[w�����z�M��i���ݽ��R��c-fb����q��r�JQqҴ(�k��޻��'�P7l����)���bͩ�pRN����u�D�v�9g��Q\&�<�-
��.8��OS�Fޥ[E��'m�����-��D��Pc��J����i�Y�;x�1ie�K�E�E�uN�{�Qh��!�`���펕����vމKCנ.Wm����W.y���ջuP��7b29�]jU��$����d���"��ᙺ��4Ҁ��nr:=�7+�Gmb}pr���k��Hj�뜗��]gU���=]o���,�ǍVs�����h�e�%=U�:�/�*�y����Q�?��w|�a,�����\�-�;^��1.7�	�v���������s�X�-���6��*Pmy�k睎�c�? �E���4����� �ޚ�9��w�"F�{h��Bn�Y�P�:�j鋫���8h+u�p�����/t���C��c�xc}o�Xz�@>�^�s��{��ӸL��w����ٞ�[Ƕ\�tM�t����s7��>^;����¦O]���W��J��b9��9���^\��81v��gv{2��=�g!��[�1?J������x�5�|3x,ϕ`R�a�s����m?��o��.w�V���e^jyۚ��k�S��'�<���q�^����f��h�Pf�W ���:U]�s[��Ȯ���ͪ��w���:��x�?^ɞ
n�x��i���!?x^rB�jt��W���:�H�y�j����p�z��M��J«Çex�5�J��LL_$N�4Y�|�l�z�E�Ԕ'�=:��A�x4lHz��N��]��l�F�<]ꐳq��n��h�g5'�@=�:Ǟb;=u���s�]h+0pɥ��3��Z���qŧ����zn���j��Oh����p;�ew��NuY����eL�{�+Z�9�b��л���l{iZ3��9�޽�ij�ڌA�[G6��m���uo�-�j�K W=��&��d�8UꤘfdY����ʙ�Q����w]�r(9u\�A;�:��-��:��Jw�ruM������I��>##�э��W5�*#�Y�
u�w�(���������}#���F�k�չ���)��&5��+z�-�aMh����~�ͮ.���9�\S}�L�F��])��^���_M4�r��>V�ͮ��_�(�yk��S5�WS؎�C��.9,nn���jXV����u�*eƚ��9АT6��f�������|��IҊNEG8�N�ߑ�n㣮`��ͻ�k�:���*Z\��6��Bǧ�Ig��v�@���'k�wF��ǹto�Y��'{%�ʾU\�W��R��Q]��y����`�y-NکM�ٌ�9ٓ����zi�a����w���Z��ڨ��-kAN���UL�r�=��U��񥍭����{3��,�WJ��n*s��G⢎{����&��y��OG����n��3{�^���W�;1�QF�}F��윫.�Ak��I۸Y9�z��i49	�R�j�>C"�	������h�#��a�7�?<g�"1�SXZ���
n�ph��׀���ٍ�c}�:�[���\�Kc�vu9��q����8j{q�#'h�b*�K�R��lo�� > ;�~�ޝ˽�e~	��@�4���+˄�D�PN�3�F�U�VU^�zc/�8��R���a5�Gg&�tS�Ѹ3���+�c15Oo�%�ɷQ=.�W�ahS���=z��V���޹]��gg*H�(�]A<�zz�_]�օ�Kx�*{�czMObp�VN���}�S���4��N�R��hT�ٝoڠ�S���f�o��P�� ��H�Z������={�'܇ ��'��LV�D�<z�j2߸����&�j�v=�q��¨O�c�[Ӓ����q���6��l<ՀV�n�SmXr�Ḝ���ӛ�u�ֶ˭�K�K͙�I�D|�X~�Ϋ�Y���3С8Y�d�t��*5y�Mz�Ku��i��U�J�]���`g(���p�FjU�Ķ�
��Y�V��������:��z�Hz��O�j[��+A�)f�'"�fXS=��[�MA�SmURMO:r��u�!L7r���4�ʘ/u>��I��ש���1N�}pgd|Ko�U��[=�o:JUs3{Ͻ�G��D��vz*۬���]��8�JgB�p�^�1g�?;�=Wm㊍��:^S\��ûc���c=0�����Y����SΫ�/���AO�a�
/|䥱��~>\��9���L�^O3���6��Iݳ��Y�賕�ީ��d�=K��9Ώ:��M
��l����j#oK����Ch��!��o�N�۠��J]����PyR�j����ۉY���Z�	Yy�t)�[<�GP��҉��rC��R��M��٭d�m���?r����i�>�A��.-;h��_\����u�?=��F$���B�����x�]�����W���F@�TOK^]fu!���^�I�կO5����\Mrw���7������`�S�+.?h��Q��FCX�vl-���ĳ�T�~lI�8�I�����n����=:��"ݖ�5�If#��<�c�/_+���!����"��'=�v�{������t�^�)����nG�u9�í�m���5lz(5��8�� �ۙ�.���7̣��㰃F�䱭�/�j��Qm�������ܺ�>؆���dOn���<K��W�}�|��w����^�����E�w(������yۭ�v��¦�G]�%7s����*��>�y��ç�s����}����Ecm�×�p&��En �;�h�gj���͑8Ɖ/\ץm�vE�����������QS�wv��ʉQ�/Wa�_��T9C���'�㫎�$�<�<>�������Gn�Χ	B���2S�w�~�뒺��U�U;O���x9�OR�P��������	��Rv���k�Ax��W�Wmt�G-��yZ�d����nbx5���qQۊ��bօ;���^q�Y�7��ا=6_MvbG��5P5�_*��qx�tNZ�\�-kB����K5ޫB`�"ko'޾�W�Nޙ�ު+�)��/9�jgi5]=�Xu����o�D���	?l�x��VhW�Ϋ�>	���Β�9��{���*����"b@���݀32/�m�<� �֖�ԺW��>��L��z��t��jf���R�ݛ�me�)\��+�a����r�r�Z5oL��'��\���Np�\�*��#tA���tY�dz5ѕv�K���{����������K^��i�M�Ϡ-yq�jȦ�nVP8v+ �u*:i0�-K�|�������'�=C�'��|����$]�Q�b|�'V�O_���3�1.��}C��G��q�R|����ul���GT�����Ƽjw^�K���:�� ��	;{���\��S�+��"�I�Ǔ�ٖ��.0�0�|;X�S�w�^W��!N�O�s�9Z��;�yP�����6�zw���d:oH_t������Q[�A����?ka��)�7��ǧ\��xt�����,�����8O�ޚ�������; l��Wf�����(d�̥�)[p�NEBoY�x�:�]x�sQ���ծ�'&[j�|5��4����`v�yOCNEG8�N����P�E~�$�A�����=9�qLUe���u���(���x�\s��/����O�����n�WۓP���JN�J��SE���y���t�ף0��q�[4k�7�u��y�&��;�]*����v�kno�]���p���`u����X�ħ���h�fdseı�b;|�E�7o9� �W�I���ȥ�s�T���c��|����v��\�]Z�U�Q�8}��Ў�Q�8�o�cB�Ţ��+hF�:Ι;؎8��H�(�͔V}|��{5g�i<�߱�����2*~�ucSꛢ{���H��S�ڞQ�~s3hћ���V��+ޭP��͛�*�9�{��^��Ms[t���)?sz����V������T�]�t���֧PS�c��M=R��D����A�W�]��`�ŻtA��ܬ~��
�����~	�����n���^��1kOV�K�S��u�^�=Ep�j�hS�of���o�gt�q�q���Soc���`�����ʫ����.���e��fGQq�g���b�rv�f��R����N�Y�{F'܇D�-tc��t��:Y��hd�9�,��|�������^/vr�o�h�!�
��DW�o.���/J�ӫ��Mk�㚳{k}�Zb:�����~��n���p$k/��J��2�^�ͱ��6�J_J6�Qn�]j��IxS�gK�|/35��n@q�:V6��u�-)MB��{9�����|���6��|:���������<�[�{��DqkC��E�[J��[�jvG{��%oH�r�Ҏv^Otn�ZK���dǷV��Sm\@r�ۉȤ�ל�:F�u�{ݵ��wRJF�R�WL]b�[U�	�mC*58Y�g\n�t,���"���=����\ߥC��F�{7W]9�`lg(ɢʶ��K)��-ۮ���T+ w-��*�y�N}��K(^�S1����/�=�ju�<����]=� ���
�y�n����%9�j�=��u1��z�Nm�s������h�r��FiA�����&��!ݱƎ-�U
7q2��k�/9:�I�uy��x����âW�*9Ϊ-8�mS�mmh۪>Á�'͡��WZ9 �%�;{����'��P�27'C TNO~�Up�9xS0�Zrۮ'K͜2���Ե5��v�:]��`��E�G����*�L�x��m�1����
[ق�����^����;Z�u'�����nƆ�4O��Ng˚�u�t����+��V%Z��jWE��lw%8�N�)��֥u�C[]r`-�6�f1�V�n�=�j���Yĸ����,ե�8]JRq��P�u���y!6+�)�Nok���ޏA�j�V^�teꟙ�˛�������D?h�𮬆�Kr!���<�gU�����R�Jb��{U���K�-d�I���z uʀ��7}�P�l�E���ŎF��qx����*�+�n�7��bP���/ˬ���(8Q���v_��F?�i�����s-�Gqb�sC~�^�IY��/�{cTw��rb�tQ���R�S��ސ�g� z��1�5��,vl�S�n�9�K�-����U�ȵ��.��K����s|*�U�Dq-j��7�h�kI��f��@uLvAa��U�Z�+E��G��iü�xy`��!�D���\I����c�2oJ i�f*!�)��M6s�[�~&�!�y����F@�۴��(1�fD1�p��~��B�2�Y�� ��j{+`�7���^�L�	� �\d4h(	�XN�6��4�S&�;�i���Hp�5+n�~�(�ы��7����KX+��i�j��m��>�>!���}�:�_���v��Lq�,�ܭ�׀L��[G�WXi����)c����j�3Ih��OJG�e��2�;U��b�^X�q�:ӏW��B�]/b��}���T�&�d�P�CS�xm�j*��ͽ�,9�i���ou+��4h��;X�v�b����U�LZ��)��x��Ԓ��
[t�V�Zvt�
��/���=�xq�X�|J�F�t�+U-�/l�^�=0�|��v:�´��LN������}�E/m�UP�����C��P���Oo�me�vH�q5�ݝ�x�k�vV��u��B��_L�J
�]"�;zy���-\g9떾����v���m(��G��sλB��7�Ps2�#�v:��z�Е�;�|d|U�3D��������Λ�Zg3
��jYm��6xݠ�\r\fnr6wU˺�;�ݽ@Ď�����p�3Ku��,Ij+�m�0d�K�V��f�	�o�㰸\���)��j �d#2�֣Xzi�q����uŴ�>�Dq��IrZ���zn��ܜƦ��z�˴ �d��:h�!��2�w�3���R��T��ץ���mI��LV��<��ģd�k#�
�6����#�t�A�mՐ�h)[�'�i�,���5=���r�;��)�N]����;`�jR��ы
��u��q�^��2Zuԩش)��߮�	��z�R����}f�C �g���8����ƒ�J�}�a�D��[�۽�����d��Xdm`֬�tÜo�������F�Eu�gw���]��i�Ο��Y�����Z���<��<]޷9Q`�]w�C�M�GGc.�3p蠑������W)C	@�b�f;�܎c��f�:�C܃����t��w L��� ���Z��o<�.gZ�4Y����0^�,�9�F��Ę�uޘ�Wf�r���5�v�i�F9���D���tUemz�:�"����vy㦶��u�	!�:���Z�-,'(�B[�ɧ�9�S�[or;��N��?&�ew:sz흲e�5s��cU'�W4!M���B��ʶV���KvP�a�fjڵ�|��N�ׁ��hVmY;�S�(��K�XDf�����u�۝�A�3-�B���F^��ц3׽U��y����A�	쫗��T����SYjv$vu�Җ�|��%����F�/�M@���xP�5�n�ÄVF'`�<�^�����k�R�Y�nҮ�63����f.�i�<�`����"�Mݤ6�b��ѥ�˽�S�|��6=�\9�U��.�y�{�:W*�x��9�M_j�s�x{�N��s�ݣ�3�V��;xK�2�M��;`�>�݋9�6�u�bWָ���tLq�4+�i����Z���l�/I�1k����k�ښ4-�3�'ڹ�da��ZF�#Uqu�q��h�fg+�ǎl�m啜��� @ ��쨪,�Z�����"(i�j ���)���R*d�ȩ��f&j*
���	���f
����Ȳȉ31h��h���"��"
)h��������"��*��#�J����*�0�)����"�����H����2��ʢ ���,�
��ih���(���l�(����)��ZbZi�J(�j(*���*��f�(�*0H)�*b*f"�*��(�(�h�b��)��*��Jij���)�����#*�*���*(��(����
*��ʢ*H��c,&�����������j���((��J���������*#0�h�))*!��b&*�ʪ�j�*� ���h��1��)�����1�����$��"��r�2i̳"��"��
b�0�j$*&��l��	�"(�&�"�321�(h�"�E�Gl"ep,��=��^���zW��u:�(������IEub⪠�k�^�|��{nl`�3���drXO<K������.5=�|ĵ&}�:������l��N��o8��Z���:D�V�_�9i�����щ��-�>|�o��U,���̏�����k�D��ǧ�P��-���Ɲ�=a�蛄*^#�_�/jY��@�{4m�B]m��Z���:��]�c��ҹ�Ak{�9�a<��e���Fd��
�ӯӓ�Ꝣ��:�o�udY�q����O��Y�("���Ī���U^k�1�j�3�:�T�<�����c��(m�gh���,(�=���s��G��l���q�kl�('��Ny�O�������L_�I�*c��"q�F+�
ׂ�X�	C�=��]/fIc~��@��×Mۗ���K�뭪�#i�d�޴�P�7j�Ut���_>�#a���&D�4�a�)s�?���e�D�uW����-�Pd9��O�x��&�����+�Oq1(:�D���+�R��
���/����9�N���ء�]����n!e;7duj��'�!i퉉C��r�b�}'M{�׷�x�ۈxC��٬uE :Fұ�C��q�E���][�I���Ӳ@���F_n��Kup�ڈ�#ʖѫ6J��Pʧ��̓�������f�ɀ�{-�{DuCʎS��3�{�n.���Ū��QQ�t�N�ү��ծ�=w܉EFb},�������o����{L��#��n��B��LsGA#�u�]�o���D��a�v�r�VԞ.#zX"���1�U.8�M�a��:���)�DW��HC]Kk.�4w��^�l�D�-{]�L&��@JX��R��NB;���������S�{U�!�fbp�Qv���ӿ^ܲ^���#gh�}Ή5��A�N������UOe��.�Ѵn��L-�*�����p���3HgՆ��vP�2����`���[kT�Km�1e�����|s%}��,.~x���^��h��H�	l�{6h(���7���q�rŚ�Gd��lh����"U�f�S���j���M�^H�7r�4��!�APx�K����3ӵ�ѐ��˕.z����Zn1�b6\��;溸u��;EߦX�h>YqD�Բ�0��6v�t
�+�6�ɚ����<�i�5e�c�UՌ��h�F��v5�Iڑ�<^��Lͻ��ϩ%�Ҟ���P�H[%��Ä�a��P�a��m=�f�,��J�\�Kt������w�h�ι�Sv��,N�er��J����B�*���;:�f�w�`Rn���ׅR����T^GizJ��|��Ah��=z%�I��o�I\ɥ�]��+�y�*%=������b�3dO��� ��M���l?�����Wg��S����aa�[$*���)�|�-�ڹ7�!斥�vvmO#�it�oMC����K'�W��.�$�qR��r�a�����:��].��ߵ����M���c&�=�O4`aIP�*G\>��Q�J��V��=g���FOk�
�n���i���Z�7_��R|�C�.���W�S�*�+���CxA��b�|��D�����=�^��r��ܺcVÚ�
٘�7J�א�ذ��X�g	"x��Q���^�f�����rK�CbШVx��3�X�@uQ��r/��>7�Y��e�rXY��6�/>���:l�D�MF��^]AXK��
�坛�I<9��:��92��0��-�z�$q]uQ�!�%�PV�ٔ"D�B(9/َ�5��Y��&6S�ۖ�uL 8�@F�'�X\;�#��6��{w��P/�Z=��,͛>%����"�=d۰���]�Y�'���*$8�n*��i��iyVi���p�jK�G��m�s|��G.�Kz�e�Y��o����|RU�/@ƏWw�j��͍�2����"fT����n&�\9�S��˷��+ ��ov�("�"���s��l
�Ӧ���.��μ���<�-�2[;G(�hBC/����%���vjr*��  	ϼ�T~d����,𜘶Pp,%��8�P��4p�jxH��^F�B�L|Ê�@���yI��B��w��ip��B�t-w��0��[T�qص�ò �:**Q��nfZ|�v�/ݒ�=�E���u9������d�`
��
�yU��	���&{��)mv��z��Gt�o����o2�
�J�g��`T��_a�$:��������cy�/Q�����ظ��<:R�9�"V�.n�F z�ں����*��^E��j֘��z.pvZ�sJwVt�o:�}H/>�NC[R��C��OTH�F��Tu�K�J�;V�)춙��{�K�t"�z}8�tcx�[u#C�.�@T'%^����ǉ�c��k#!eɍ��U�o�Z+N���[�r"�|��l�-5�?zʽ�o�L�ɵM�g��@x%+|pP��=���W�z����:�)���]��n��mt�m�c��T�k*�1�����`>rB&��WT�Td�
jx��(=��YL,���yt���s�U��;rsn� �w�'�6*K�J�dHj\������qO����BH_���{��D�]Ր��N`m�o�q��N�XN�U��"���@.�wSxY8Nt�8g����0��KQ/���v�j���]���M�UJ`��S��Ͼ��r��B\;�B����>�7�&25	�j%OS,v�&��q`i�RCo{p��V	�����ۤ3�߾��,�Xck�dC
l��}�j$�;WH1^��b���+ �{Ɇ��66�����%�u�d\C4
�N%i7΀�.�P�dy�ʻQ�]�H���ƥʇtmd��^-�e/vL�t]�a�����T��,p¹�+��E��01:�����%ڇ�����o;�2j�C��^֝�
�9:���!8�6x�,`����=��b��[8�y��Ԏ�X��ƪYG�ǦG��O���{�Jx�z{�s������]\�'��ne���vHO1���<�?=�6��t�j[5�B�ћ)�q���y��ͽr�l�m޾���ʡ鋏ct�N�[�'h�=�{x�3�dX16����W,܅��Z�t�:A9a�@K�&giA��0\=T���t��{��%�v}�:��ZM�oײL�g�ZFĨ��	�<�+h�!=�N�����=}c�g�����;*���bl�^4��WI�۝���KGѩ�q'74< �5G�c���p��XB�!�K(�T��I�Ƨo\	K���7�f�gK��S!�G�]-:a𳝂>�^�_T-X���؆�1�k;��}q�Tg6f?������od����C��l)$B'��&V��Q����O�{�	C��Zp��B�����u��JgK.HQP
ɀ�صTġ�E�R�~#�מ�`�_tOJ۞�˥�^����Oj�Ǫ��.��s'(?��������R��Qq>u���W>��gC)XXp���+װ�u�v���ٝY1K<+���P�ޥ��1��%�\�X�����T�:%����ۥ�yݽ,\��t֎�e����r�cne������'�����]T.+�=�I[M���Y� Vrt��PB�L�tT��FC0�)���2CGY� ��Py�">k-=�hWڋ5Ա�7~�w�JX�Iݨ��#�p����,���TU�����p�s/^����֝p��0�9%�U�av��b��'S����@^Nq'��s�j$�p��!֞�Yp{�r'-ٰG�˴Ǝώ\���C;f�E������cF�[tZ��.�wI�8��ZG)�7�f��7X :�x���7CQ��}�]A�I�ঞ��ug��J�BDr����n΂ˈ�Ö�o��7\���A]2y��]�s'69m�V�V�q��<������3TucG�҃v���'�n�$\,��E��J�q��(E$t�<�ʳ���⪁ல�w���8t�a�6R�4$�}y~ >����NW"d�=��T�{j�~�,�=����gގh���q`��b�^��!+�.�2��U�;+��΀�!"��+���VpBea^Ʃ��sc0�]\.#��`<Ôt�z�>��Wc�=6@�S蘘�1�+�y�mW�%:�6:ZrE�T�gJ���;�k����&�m�̽����(S73,;�t��X��H��,׃}0�'KK�P�)���Qu��~|�'YKuգ�UA�^'��7�sAܙ஝PW-*1L,7�BX�ŪX�:Ì<�ȕ͊�C�R��ǒ�P��l��Oiw&x+�J��˕�2�V����j�٦�ͬ�y�Ev�h��[�3K
�D>ʑ���`E@B6�'��*U���Y��G6�����˜��^�I�;\5l9��'��\;t�˯[�%r����e��y�5Xŷ~:g��yb�S{�����^�5�~���[k�+�3��ԫ=x�رn�)߬�/�I=!���{�YI���>JP�6(Jk:�K���O|��{���܊9	�=6�@ٖ�w��'yСCw�1���5y�vvY��g[��\�swڪ+d
k_Yc�]�v���4�=�r9�U�d9Wy����w�M4�i�j���#�)[A�v�}�U�g�.մ�ej���S[�F�[�i=rwY�XV\���Ać}�����J�ܵ����|�'<H�qyh���ύ�2�9�\e�e@�f���W��{�{�R(B�k˲�y�%��(+K���R�e��>y��ߙ��xwz[W#�o5� ��Y��J s Zw5���L5��D�C6e��يG
y 8 (1�~�ܚ�6�(�s}V/y�������g��+��HM�9)��/����r״�f2��}�C�۴��z����E��K]"q䡻�Ǝ����U(���/���Y�n�����]�k|��NC)�w~��@q��IWg���>���{.)x�[��g����>�����d���D��:}]-�q:�9<�򫅞	�җ]��b	z�1en�=eiv�p�[z<�9&軗\z�@�����[&W��|�\S���<9y�'|����m�k
y��y�r�7n)fJ08��5h��F�CC������Q���;��<��[�d*yQ���O���^��v4:y0G���mN��D��:UY�x=�_I�'��݌��|Y�����{�o�ҡ��]$�"��=qȁ�f�w�nj�o4��Tf?}1R/�qz!�z7Z�g8�T���b���I��F����m�E+�U0@�!�l����r�vd�K"���캷�w^�Inqg�ޏ{��[،��a�����Q�Pz��a[�r-���ġ��.G�]f��NJ"y�]r\c譼�Z�Ҥ480c���aT��7�)�;K��Cw,T~n���+��o��v��ty�V�o\o6�;�9!^�yM���@�_RF������
y��%ي#��0_E^���������Y��	�K����r���V�T֓a��W�)��U�4/#^��o����Fr�2�Q�
��n*2Lf�<MzT�u{���f��c|�@�����%柛�"߶l!Ќ��8���H�P�^�m-��ӎ7���杵Ih<�e�=�_<�v#�*�1�X�"�
y8���3K�A�S&�>#�q�C���/<M8�՛9�&{���O�2�����A`�~�
��L��eS�~P����MHvClB��s���d�{3E���SNIp���Te�o� i{�n�b�i��SZ�|�P;e�/-c,U8|yX����L+���d*�����ș��s2/��=B&��G;�m1*��7�S�GP�A���;��xj�"�w������^-�>��Nm^�:i�h<��^�Jr����)m�z��ن�Z�Փ5mtt�܆Q7�A�2�N�f��}(t��4��45s� ͋9ocʝ�E�*Wō�db��ߟ �_q�A.�zv,�c�K��g4�zp(�{]F���PP�3M���
�l�M�݉y C���|�g*Ճuu�̆����鮝�k�9{pm?o�t"�16�)yXs2���_j���]����΄B�|XFz�i[n�]��$1pP�6�v���\K��Sq͇{Os"�9Q1��<8��:��B�},\���}�~}h!r����F����-f�U���<C�pc72º��2��	���l�ib�a3Ⱦ��{kw��t�x����n�NG8n�x�$(�d�A��ޙ��ҩ=��3[�7hX�X�^��]��~ž�7<����}R�f���
���
�(��PT�W�A��%��8�VuT\*z�(��C1ZjE��y��3�Ӄ��U��!�+7��7�w��MM,�����}V�[�O!�c~��v�Q��S�j�9�p��:Bt�V�2W��8A� R�#��G�u�T����T5��$fM3r��$}����]ʸH����S����f�uwa���F}�<{ь��7�R5t:+�5[
`o��Vi�Ņ5�O��D�!�ʐ�ڭ�L �ݼ�h����u���V�雬P�'�6�����㻗��z��l����]3�ZTjf���R ��KQ��7��>��۱�f�D*=}h�4�3����b���K.ۛ�a<�]�ȈJ��nP�E�F
*��XkL������Ω��/T?K=��쇚j�YÜ�G�jb��
��y[�E�NX��)���]����6���jP;q�'�'!��*��t��ѐ�!�nF��ثP��o��j��I�'��^c��b��]�2�]��z���X�6�bָ�KM�F�	��S��7N���@��i�-��a�y"˔�wMb"�<y��쨏0��*f@�v�dQ�(�ݺcu�ED�=Y�Hآ��s��b�tC]���p�;e�gvu[���i�oۼ���������\rk�!F�b.�)�]}��t��Z�]%\UۤK���-Yk���a���,}�p�u}�̷3r��Τz�	&����D�꛷�V�P�V�;U8[�Z$�h �ǯm ��Z=��e�.Q;/8<��ړy�e::�:���nص��l�q���Ce"����hTa`� �UlPk�.m@�t �U;n'�Š�d��7\��n�giV�g��Tbf�k��E���ײ^�vMҫ�j��ρ��hU��u�yNm��%�S���S��*�:�Dqfy7����5���>΍6R�hՔmKҧ#S&��T�yL�r��q-꛺Fu�X�ac�#��k�M�)ځ���YC�xuR�^�FOg�mZ�cYө%�2U��KN!u�ݦmw9�����V�2�ū�5�Z'���=�v�������Uǔ#I=è�Ş��wKvz��ք�ZbH໡�$H���J=��k{/JgeG��E�+�������6�������t`źy}ƺ���@�si�U�`���\��8#�%	q����8C�W8�7��ߥ:�#�|J���y��"��KNd��7I���wU%5o"%�X�@E�b߮�̻`pn���Hn)[a��yP�d�6�j�ba��ͽ�.ۢ�9�z�c��+���"B�)��"�I��%e �j�=�m�����jgVd��*=w��w.�Uw#�r�G�]m!ӱΏX:�s�m%�g��ΤȆ�+WTsnh��vH�74�	��S7&�F���.��j7e�*�APF�\�@�/8��}�U�4�!:�4��Gu�����u�����R�R��Q(c뤋��GvF%
Q։!7a��+03I�BoN��W.8�Q�f�z�A���Yw3N_�z���ĵ����Af���]�<or��ϳV<��V�����	�T��#�'Pn��I�)���JP�N��z�b*jrR"ծ�k7����>h٥^�.­c8�ީ�1r*u��aV�Ӗ_ז&I�NAe�1ILQfeM4Q3��ED�5D��L�fD�FDEDĄ�UMQT4P�QFfQL�QQfd�DQU$�eXKTQ�FD�$T���EfcA��EQ5MQC$UTEU3LMD�AQD��T�QUUQRDEFN$SEAUAQDUTUCe�TQD�TUP�TUKQD�%TE50A0�ERUA0T5DMPQQ�-T1DS4A1E5QDP��E,ITf`DUQ$�5EMLQQ�35TILQ$D�DL��U$�X�1CQUEUUPRD	SM4��dEAEQSdfc��d1�UUT��PdeALC5DS�`DDDT�CQ�D�1UMEIU%SMRTԕ�T�NPELDMP_���s6k�����mj������&<��w+��s4qSM�qL�Tz2{�<1el�.�*�@��NeE:���9A������+�=]�}�.���n��emBܝ.n�]�&���:�b����U�+�=p\�+���wmte���峃�J�1�6�p�%��X���Z�TN�@��5/��p7u=�-Μj�M�K�r8꺩�����S����r]�;�:�t��ɪ�]�mw���Ԁ.V�"��R�r;����s�牛�f�����n%�$�ˌ8HT��kV��ض���U�\t�C�jȼ{Q�Z87��Y2'�a�4��a9��i�zO,�C��4C�ڮ����nt%=J���Zn1�wMo�[c����(4�wɥ����\s�-7�	���A��
�<�6�ɚ����t��E���i�U��L%p�z����pf��+�Ih���O��,pH��,�o��t����wc�wչ����c�p:����혵1����͎�{���]fsF�}V���X�����ל����<���ޜ��� ���Y=�OiwgGJk��*��Y{�,-e�
�=�fbwE�e�1;}�F�:�h'��p�s9�~i(��|�wM�����"֭������(#H��{25�R��7a"+��1[��A���c(ĸ���g���4�嫥�[��J�5\]T�vj�9�W��X�v�/�UWԧ-4��w�Њ�*![��#�[�01����=�*�
�
��>��o8�'8S�1�ˀ&'z7�:P(��r�[k��!>W"����y+��)���e��y�X��/���f��*L��K²��ї�4�l����؇5�B�fb��7.�[�b�C��cC��j0>�9��v ��I#��%�Ί�X����qi��`��u��+�y�w��j��F���QQE���~NV����t�O��K�|��2���M.��vhln�$�e�1ܣm4NԷl��J��q.JFO.��#�$��:�����L+<,A�w˹�K@��9����O3w�����"y8� �rTByW�*p���j\���T���.�	��8�{+{��|;e�X�j7��"���"�<+I�s�"b1��H�Zv⸋فT�*���v+55Uuow�W��iS]�2�����¶�!k�M�=�;�%�*!�� \-2ũ/��9�o�ǎ���Z�`	Jd�E�ڧ��D(����O:��R�&��c����aGR�\��(�� �P����J�2��o<M�A�I[2�t�
�f�/����<J���
7���4�2�U`Ꮹ	p[�9W0��*��*���@Ώ/Tv0l�3;#O&��S�Oj���{�-N���v�tZ��+J�/3q�Gd��[��N��A���7��p��XR;�ƒ��s�l���\����"U� :V�t�o9]Fx��hu���Iuu�"юei��6�d�(A��6ϧ��A��[�̑q�['p�u�Y�}��^k���gV	�������qh���\�P� �!��#���1�e��hBڤKl���G�o9����u��Thb�S�C<�K�9mHV�Q�=��
V��j�8�P�ǌ��o0B��UG\J�&���<��b�o�ȸw1�S�}�#���4j�I�{�=�7ڶ�����?� �8q0�"]v锊Ӱ;�o����Ex����yyrX;O���{3�ʒ��<O��t82���%�F���L���Iќ���$�φ3�E)�wn��2<"��Ýz,L��S��$��T��2`G�����8�f��ȸ�ޛXɫ��y�c_�U1�' tC�b+�n*2Lf�<IG���7��zP�Cn{�5���z��sT��͆9D�q+H�,1��C�8EC�tOa���]�+���*�}��UK��qάkE��u��9��3v�8���xy�v�sZ.T�RW��_JO=�
?P;^�b�,�"�|2<��'|�Hk0efQ<��v�<��C�k,����UU�άa���#ܳ]����\T���
킷y�VW���	���1���&�	Ux�T����w��P�,u]�KI��@htd0�4a��ʹ�[�����8�o=�`W�h���x�k:o�L��򊂵Ӂ��CO:Ĝ��Ԛ\�]pХ�Nof���":�X��ghWkZ/��w�����
�''B���]�U��(��L�sUۈ�bU�6Q>�f��&{��ƪY_V=+#�^��Da��յ�����"K����{�zxF�J�/w�v"��/��c�X�ttSg�YT߼]MLu�ي�O6�Z�ͧ�+	���S��T-1~Ʃ���r���=��o8��ȓ�b����h��j����*u�ʵ�[*t �ʩ�c
u-ꥥo�����c�P�4s�'/3��+��wگ��N$�`����d��QQl�*},�Q��}�o�ъ=GS���9�کq\����@(s7�����\�*��l�ib�a3Țѝ�kf���~\��jC������b`�1C��jE�3s^�UA_�c��)��y������)C�5�/Ɨk�]�)ח�&7rȲ�6�����eh�iw����
�$.����Vfsv�8�摇��L���uUtvbwSa�I���J×�����pݩ�(Mg��f�	��X��ͤ������ҩtC���W1��%W_z=븧k��y�N����Z��aI^}$B{U08"v<�J�Q.����e
+rP ��]X�V�o-JӮWp_)��۪�})Y� ��g1<MD���bP��)��FZ3V��n�|�'�六g�������YB���t�۬����s�W�&���IY|/;�5ӊӶ���]$*-I��焎Jq�P�^��q46.�N��1^��(TK[����W�t�,EЕ��=N�7f�b�n`$�/�t�}q�!d�ͬ��
t)�&guc�l�����@�6���r�����i��wyvx Wݥ��7�_n�I�7,�+��ad���/�v�VQ�� K;����\-Z�</��O��Q���T�>��h`я{�^� ��m;���l��?<L�`f����ϑ�GOF�Lz��E��=�`��x�Ⲑw��Z�/���t�S���j���a�4��a~�k�ީ�y�D<�"zg`1ˊ���
�Y��2�߱�b�ߝ��u�ע��#UA�E[n'�W���06nɍ%���5|���&Q+&��=$��de�����b��+)�UĎ!�p��n�º�A6*w�����P�-�N�$$�n�B�M�x�<^^�l�:Jۃ�|$~�P�s��wq떅�}!.��镧��-�����&Us,i6��WL(9yW�5)ݱ��-0�c;/n��l�}��g�^�����f7��4d��>1%�ҟ�O�h���C��<�}wU���hIS�ޔ���32		cQ�·~�PY����B�3�����&�bJ�>Ӫ�7�C��h�+�o����y��D �R��}�0�����'p�"�tk���������$U�6Wq�;B����yԫ��4f���o������J�щ�kz��[nkf{E��D]yE4�^�5k����T�v�ἇ����p �y� `\�,d�}Z�w5�ф �!����F�{���7ҩ�LΌ	1z[/B2���ٱo���Ʈ_�j޵���8I�rx��B:O�܋b�W�x��І�U��C���X��z���n���z�]n����J�{�Fٔ��Rip��b�:��3�$�!���L<��Ɗ����١�mS�~J@���tOn`���v��di��V�r��ze��ߎ�-��+v����P�{��2��S�-�P� �ߌ����1�����M���Kuv��J
��{T>�޾${�iP���YNͺW�<U�]�q�qq���.�&���6������!��/"cY[�\:�u���6��t,��}�<�����|�WF��Ws�g�]D�� Rq(Q�U[b{o�m�#���^R��zD�^0���y�y~��X(-��XnS�EB֬���&��1���E�-;qF9�'c���[X� zY8;x+�#BVV�{c|r
ڿ���s|��GY�w-�@����i�狤���#�9�^)ᄺ�^����Z�.�`�z�*�cΓ�U��f�r.����v�t�2|�-��N�Z�+�dld�`��,mQʍl��y/��\�mF0����a2��s�z�ވ �N���������*z�Ą�z�p�׻��gY2����K뇞
[ٌ�Qž#������!�`P�e���f�#ܣcY����;W��`yv �!����F�/�S�C	z�!��
��#�h;A�ߎ˵�W7h��{�s�8E�#���U�Uq5�Pz��b��H~w1�S��r8K� �!^u�'�Uw�؝�j��rY(���I�\��锊ӾŊ��W"��1z6����7���q���W�e`�Z�զ`ᗶ�@�5nH(U�΄�� N��/nT����
��*J�t��j���`x"��41�Ӓ�L�B�\��O�օ�3���մoS��v:5�;I�<B���P�v�f��v��5�{�]��t��Y1<Wa�>��S����K�БR��}HK!�U�^��9j[ă�ɹ�SkΦz��l�!�p�]�7	��BrB&��WLu{ɭ&�o-�����w����J8�^�]�,\�̗Ք����,:;���D�Ȅr���Bx������Ls��������9~Sɼ
��
�2�TC�)��Z�D
N%i�6�Ub�؅�x�Jȅ��f��)k�;Jp���#����\ǢU��RUft�]^Ox���	�XN���]�8!);��i�/���Y�MW�G���en_�<v���4�p d~�
��)��5M�2΄1Wy�E�:��uȎ�gk��ٳ�r������\]:"��m-#ƭ統�K|5]�s��:a@����~3r�Ϟ�uZ��دŝ�^��D^N���&_�h�-p��N䴞e��{�E{�d���@��f����ǅYM���.�%�V��ι{J�W��BSR��{2�G����j���r��yq�ޙ�$d�9��]��$i+��i�u��ܦy�uBwg^�H�g�D�W�Xe�,'.=��QtaꝹ.�.�Jk����hK�nּZqr���#.jz����z���t�ibQ���7C{^>�PC�5C���@)�l욲�F�n �t�:��������ݪN���&:~JU�/:XF�B���2
u.�ZVźavSܐ�}N�hxf�<}�M���]��LpA���Ȣ��C��b�\�>���s^�Ը�k��S�Ur�+h��t����Ih���+Z]���=fUv!×Mە�ܗ���L�!�g���=O���\C�5p��Q�$(�P�o�W��u0$;�z\�ZF\\{�u�ĭ��hX���W�Y�B?<�����G����C��L{�v��V���l2�^�s.���-�G]�/Ƈ�f��𼇔�ø0��A��OQ%i��{�)3-:��oaH�(��N��w*��3���˳��'H�WLm�:��x@�̚�;r���:v_(��ݪ��oO�n�K����Gf9�uO�y8�����l�ֺ���2�iݾ�W�CC�:h�b:�zK�n�Y{p�'K��n��Mz� �T�eQ�F޳�	���X{DIP�u����NV՟]j�C��q�u&Kd�/��%s�l��ʳP�;n7[uf��-�"�[�ܖ�]�ї7�D�2��H�����]�V�e��5��)�lut�O3�U�^q����Yi��˴�ʡ]�E�Q��'rR��J����h�G�})�� �m��F��q����z�zYk7N��2��\T�����%8����G�yw"��p�H_K5���xn����Ae�q���nb��:�y��m0Ry��)�p�ư��8�ٮ���r���3_��������>�D?'����j�X���kVF<��-�ՑÞ)��8k�ꇙ�h׹�T���Ҫ���]T�X�e�VWsԬ��	���b�}���z�.�a{��%�ߦ3yORvf�2lg��A[���/�=)ݱ��-.�a��@�����{��t�������X�ڋ9)+����F�	�� �� yl�cv�飒��*�.���~i���P�p6t9s��x��t���"�t~lt��Ċ��@�특�QW�hf���'�踍RGT,}�L��0�͖֚�p]b�d�
�=�ܙ�\�u��eVl5�x�r�a���[D*���B���b���o��P�8P9�UM�w=��n<�e��AUu�P����,bNk��>W"�ۧ��oD� ���YJE��
��!��:�K�eT��<��B�)�r�-ʄ���� ���2��(����X�g�Vl��h�nդ�m��hfp���ܐ}��F8�N�5�;;v�ƸVuڦgu1�!u'3hKw��R*2�\�A��[���$��o�ܯ]Y�
��yOO ��ӄ�2�9����DtĖ��"�����Wɫ�9�Fb�ΕJ��(kga׀i�8_L�R�kr�c�	gzm\߰5g���Ŏ��b�*JR�2�+�v���n��q}��<��SdQ��pP�n��>;�����d�q�,R�W{�K�U�$�mE�
3�$�>{��3Nݵ'T��ʓ�QV�Ɍ�Ī���7��Ru.7��N���ݾ={@A����.��D��6�����V��������S|�gE�����R�j�4���Q�ڰ�WN�h3ݘ����5��S8�+���Յ��F���,pnJԵ���RV����y2^j�N�5x�Dv��I�MK%6k3p�0�(�N8�BV�)�����n���2�&���>7sn�;�`b�YЍ%�Ҙ�@B漢��H�f��,o�f��KuͨC�j�Цl����eѢqBe5$#M���Ws��.�#"���֫+����7C��f�~��T�!ɳfS����áL
�"�����Tt-����.We�8�:hX�3+���Y|��K�#�q�l�W��w��`�y^ʳ:DOm�#�$��*��uZ�%s�w/S��1�
Ŭj��3=�i�apr�w]�ip�qY�;ѶԪ4'� 0�o����˛c*�1�����OA*3�r��2B��y��te���B�DI����py2]u��	hә�ޅ�����x��z��x��8�p�� �e�3����nT�S!7���qI��(�9�|H*�o	��T��%�i�P�XU�ח`� n`��,��.�@��be� ���M8�,�t��}N�Ak_d���lZ���ܗ�C54
��6������k�9^2^t7L6v������SZ}A�������&N�
yK���d�"Q=#�iU��*���t%���T��"�&	a��˴U��pS˔-!��F-�I��f	ו]�N'�/:��l��hS��&�7��nq%l�s*R T��y�#�K�N�3�u-���Ŕ��Cʣf�hi-�jT[��W��ץS%�$�V^t��i���9���t�'��46ku]})��E�J��;��oG�޵<^��;��لVl�ݺm�R9�����(�C�pvk)���;�����-����RJ�N�`�r�B�;w�����Xe�=:�����yY���m�Ә��їt
�gI>�5C�vdd���NR�t=�uz^�ӍS���uUT̕�A%Q%STL�LMSEQMQ1UQCSQQD��QTADLDU14DPTAEMA%DTS��ETEDD�U1D��0T�TSADU$I5QMEIUQQ0QQ5ASPTUS,MCD4UDDQ��Q@faR@D�U%P�UU3Q4�U4TUQUD�L0�Y8��SLAMTI�STATTUQ3PM@UE�A1TQQDJAL�T�SU�QSAQAD�EUDAT�DL�QEEDQNfE%T�E�1QFYUUQS5DQ4DU%QPPSU�e�EHDEA1E-R�UQLUTIUQQEUQ4IMPEU5�M5D�D�QLU3,�STQQ$E�Y�LQT�EAES�TAM1D�k�3�~����Ȯ�ͅ�8O�liUx��t0��JmX季����f>�[fj�񄪐��s>Tj�dgq��ϟut���C�_+\p�9 	����&5|&_V龕Lj�s\4,b��7.��t.RN�ؕa%�u�j8ppSq(6p�'��$�C����,b��u)�Y�{�CZ8��ϸ��51��G!)��k���O���]o�d�襔�e��9����ή=��A-�qA8@�zP�S*� F@��a���#�$�p��5�s�7=T�4����5ѫ��:��Y�&�:�Fc�{[�A��'���+���O-�+ӫ"�c)���q��׽x;�V��)�Ô]���׷��"��dXxV�~�@D㽸�Wnyeս���hsk����}���͠%�ʳO�T^�B�h����vp0W���&��!&��N�Q~h�U�����P�۶9V����,��X�w�Y��B[c�۴[ui���x�al�=���������a����
އ��ƞ�&�["�'C W]��wi�w�ʷpc��P��)�L�9m��W���"�?V��=�Ɯ�(B#���?+	R�Lz�0��n��\�c��ūw/M�ǌkf�JO����hMU�J���������
�ǦU%��U�ssA������E"a�=����_cԮg�=z�m�=}�*�Y\&�X���+�E��f-��}>�n��fS��{.CX33o������54�O��"�����-��>�NC0���̔b������+�<��)ǩz�[�:��*-J&���Y�Thb�}hc�/T�5�![�1S��Q��ec���k����D�H�*��U��)A�y���E�W!э�ɉC���s7���y':�d�g;��vhD� !��#�W&���89)e��>�Ύ��k�g1��.�B�ծVV�j��^��W�5A���Z^�*<)SЫ�!�W��*x�ŕ���|�%s:f��4ޞ����]��u�P�!��2B$��R�c���iv���B�ݻ�Ovt��C�L����tX�jS�N6�4��].Z<��Z�޽)ÕG1F�7�"^͢����>�TB��u�)�@��V�~,1�fD1�p��
��ۺ����W�H�*���b����͝w���Ͷ̋���J�o���O=\F���h�j�Uxhhndخ3.,���GZ�'�x*a�o�L�V������۬����o�ЛNfﮅ[����Wc���a���� ڛ� ��B�ᮀ:f����r�Rݩe{=��8�P��k�!���LXʑR����V�^`ڗ�&�N��N����l��L�Ԝ���!��jp��I�>��l�F:�5.:>��%b�y���>���I�j��.�Eh�9��ٳ�W(U�S"6v��k�Dk�N�X�w{�o�K�_L�R��x�p`{�[���Y|�h�*�;��G��1>#y��O�C�>l�X���w;v�8�X�UB2�m4_��}�g�i�7��c�X�)	nW�\}4�%���PA˕~O'�5�z�~���g��Zb��S];nX]��#E��5zY�O��vԉifb�oV��La����Z�'R�)~���g�h��KJ���av`�xg�Sw�U�>T�U:�i:xvf"�P���Y��P�Уp��B�'��NyF�D9q��fcμǚs��^�۴�xi���<Ex9�O�S"8������kd�M�W7s#���T�T����ҙ��x!���P�1�T��h^ȕBGY��Ş�Vն�mwkܴc����{��N��£^}$B{U02#�'�Tx��&%t����1%E�6���/cq��Jp���^r�a�U��x�S��C�w��ʣ� �{0`G0t��Ku����淪�>� �9���3|�>�]Ѕ/��j	%��d���+���]���櫲�q�'+��%lt�5(�SrV:�۳{�4�S��oj:{C9�k\I�g�о�j򫄘lY��U��6@��hq�/|6537��c��r���Ђ:��9�u������֎@�85�+�U,f��X�U��
�x��,Z@��xN*���(U�:k��	��0�̽=	�������[0����3T�`��:���"�d:+at��S�g���+��>S3Ή<����>]���K�ׇ�oKR��!��*!������:@��Ж�_��YW����^7��fb>9�����q'��,��*��ad�s��]�H�#��w�i��&��<�����V�kgg���:C����v���P�R�y����\L�dXX�	��c�:��n�F���095Ƅd�f�6h(��c��-kVF5��u��p��*��	54�P�g���[�ǋ�Y����7�=B�(+ho����lOR��eiƥ�η0�P�������d/>�r��;�C�j��פ����g�eO�=)ݱU�r���/����3M�u�"�$XՖ�a���E�����$�z?0� ��_-s��)K�8x�$�]Z�%9�����s[�N�U��D��(�x��g��R �U&c/"W��5qٹ ��_���R�CW�.�82M\��nʷh5Ԍ�A]\]�502�⡏z�3n>�ί�ΖǷO�ԝvP�K!�:���;�OQ�{b�7K|a{Ầ��i�|%G<:Ө,������O�Z:?69��0���7[y���.��6�Hu史*���0�͞�Zj�F�Y=��,�@];���i�%�g�nv�g;9C��D��E��-[�3|XTjeH�}w0 F]��k3��8�ڝO����V]�L.�E�Q`�vuK�5l9���\�v��r^�YeV��p�������w��oQ�Hb!� �g=|&_V��TƦgF�a�止]M�X��s�!�=Ȯ�*�<�.!�E1p�B�#��R�#`P��Ԅ�\Z�u)�/���^��y�3�W�Fx��R�e+�	7�|m�E0�̓��H�7.xD�fu�j�S����$��ś3oӥj s,(s*� F@��a���#��z�uC~�d��}����_��ފ����b�Ѭ΢�� T'���O*�o���L9k+��d������P7K���ŕL`�ًf��(���4�p�ZՑ��w��ȑV�X���bN����|�֦rǔ{V��$�}ف
�4�û�SZWik'�w|�	�oE�J�@GpIV�[���=����Om6�Y��ts����k8�h��1sB%�X��f�8 Y��+7Y�����pv��;���,����S��k/���3-<�X�fi��ڨB��Qu������*7�:���5���e�����Q�0{yh!�~��9��x���ᄹ����]!б[/��
�Z�r�[����J�7����75:||˫�'΢���\������u�X���s61��՗a �J~�up�'OND3	��"ۮ�+HB&�zNQw�u�����r���9�۪��Y3,�)L�{LB/�@R��d>�K�gB��F�6�}�^.��םÙ^�%���X�\M��+cF�6��g�έ�7��mH�`��+�[�l�ǜ� F�g`8'�:$G#^�U
�WX������B}�4���"Ώ`V���ZY�V�m��B���P��Ex8T1�Q�0�%�a�锊ӣ�����j�cV��v*eR㋤>�����:��=4���:O%�gʏ
OB�f�քc�[�b�(,�_�=�󃬽��{�ܖ�O3�q�1B��]�7[�0*�/�壜o�jx���=�h]�\�e�)mJ"�1�:fژ:��Ëh;:���4>�wnם_��`�z,���|�e����7w�
i
�k7)*2Z�^[Σ����,�s;2V"N�c�*�:���=�Dv�W�G������ZY"u.k����g4gj� .(�aoNyVS=�1�Xtvùb)��CB�I��Bx���k٦d�6p���0���ڰ�,�&31���c�DN%iXc\̈b���.�(�i��;ռ�i�z˒��]SV^��:"�UA=�m�ق�x(Ɂ�6����3ެد��|z,O�#zji���V���xشk3<�	�f�:0�unض��I�Nn0������G*�7��``y�؄�V=*�q�᷊�\&%��gh�
fkOg3����{��.9����~���o�n[|�h�B��h�y�Ha���ܭ�YX�!�;/^��!��	;6S"--���i��Qnw���v_��eP�Z��V��#����c׶"��\m�J��A�Jwc2!���/��w���Or4:�2��\|�
c����襅�Tb���50�A���n'B�*�s:�-+(5�`��=��n����ST�T������$�� E�a@�X2�J��ÀG����K���LLײ���3.:v�ǫpm\��ʚ�۸�jW�i�;�}.�A|��?co�],(��
��D��k���ī;�zw��A���u��V9�*���b�z�Jg�x����N�ưq�f�I{�JsuX�����OTQZ�ڲ�q���zhvޕI���ⴉ,|\{._��o��[�����~��J�r&V��P�9��WU�s]�o;���XL�/���(}����n����
ɀ��2V8�jb�i;��S~�ةxMb�:�|�&��*5��U��E_O
�T��ؗ�<����$̎
~�d�c:],=���;��N���r�ø0�=�0#��D�Ty����|�-'��}�)]c'�c9{����"�]��au�xʾ5�L�Sc��R�vJnMET��*�Gm��W���#\��^���T.9����'Mw:�"ҜfDT��}nN��Ig#�wѫ�o��׹V|���C+ah��Z�2�m،jg�1�`$��OގrY��=����;�JJB;�����b��*p���"��C�����swR�uY�Yk�絨�|�j58�5��ͣ��#Jחr�l��H���^L#�^� ���X�ss�E�Yё�4�,-��B�`�O)h9�w��gJS��E��o�yID�7 I�↊^���^�l0T�����@��Y�aX�=B<�i_D�F�t��<s���?F�VS�f�Q�V�,7O{ik6fS{L�RĿ��s/R�֍�y�}6��Y'n�y4�Uv����	��+9`���x9Y� �����/\bs�ݵ��_Y��|���O6�'f�ޖ(`Z���j7N5:9��j�/��66M���'̣~���a�4��a>U�>��R���*�}N��)k�l]_xs�b���ҋS�$�t�a���{���=	;>'��g��� ��a�Y�^L��K���q]�gT�nJ�W���48)SӐ,j�L{:V^��4r�g#~��\�<X]苒�l��V(�yǞ	
�q�O	�ø	�Ӑ�J�·t�4O�n'����3�
�s2D���7�؎N�#�ʽfv"9����>Sτ���Zj�F��/v�u��[�{:(��C8�+���Xؗ+�r�]�-���=������Ć�P���ǎ9�szd��}��CB�>'t����Q]E��xn�cV��R|�E�ۧ���n�`T�4��׺q����� >r@!�9|&z��M��S��pЌ��� L��8�AK�#1<\r����-�n%��x	�rx���#�Є6m��^�㲣h�WG�a�ˎ�3� �Η�Q�OA�N�et!�S��+���FCW����[�������G��ǲM�d����Rޛ��[�*���J�Ĺ���m�"va�1�N�X&3a�g!0<�ѭu�؟�_T��|]��g
���.:Qj=!R9�f��Yﺱ�,�46D�����Y�Ü�%�f|��Rt����y��5v[�]�0n��b�u�&�s,+�uJ�rd
NFO.��;RK

�,�4ex��|m����w\G�������,:9�H9ʀ#��N% 9�/!<�
��m�=�Ĩ}�<�[~�\C���].\/-�b��U�gҵx`.�5�Z�8<+I��"N�����ZK�u�^�.����e��a��,�֗���Ln�J���+U<xz�}K����ԍ�P�\�骢\wm!ݱ(h�Q�Z_�#Uj�JK���^c~�~�:!z�:�0^�V����*�e���fyK��j��;�[\;Ӣ�ƒ�Ec!<p��~��.uﻷ'� ޲�w�f��!�����ߢyU���=8�&V��n�vy^ދ�V��]_v�ɕ�/���Rӏ��j
WD��-�oi��/�x)of��3�˛��=f�O!���Է2N�^%�I�je@ᶥ^�,=�}d:��	� ��5�Ei�	@�	n	x��'5�=�최Ë|B�	/�֣j��б3�Z����f�;ː]͏n�	��M��`ʵ6�nL�͊^����M�R#�6�c��p$]�-Ȝt1[��l��2���e�����[E҉�s�T^�7.�����e̓P�46�+i�e?�\6ސ]�Y�<���˾Lmn-�9L��b��;0�X�u˛!{ʴ�(n�q�pR�{G��&��������-Rvkފ��n�ä��snT;�We�D�"4�����\�m�[9g���ٷx!ŝ+E���-CGm+v-̼��"	��eMmU�8+6T���
�w���V��u%:�fNu�w�Ii������aB��/D�E�m��¥�uk�ʳE���tg��<v�p_9S+iT�2fj�W-]�/@�[�3�3v�Zo�L�+�Jj�9�|r<vN�sUf�Cw,�m],}F�_ri��� u�׵����v�evQ�4T-�4�A��Ÿ����Ea�^���.4�$��٬#:N��7AE�(�k���aߙ{6�d�%��
���#$r80oT=2��z����=��3^�-v9�Ԋ���]���y2T��J��u���a�@��^^�n�ƭۛGo�`�Kej[�q/M�+Q4��B����ßI���ާKBR3�%��;-e��:kG�v��el�;E>�(`1q��
��s5ǅ頨T�պEu�'s�>�VZ�K[`B�R�+�pDhqs,+=X��U��Ph�S;w!��+���E\YOo��E��]ܭ����u�rp��܆뾈s�<�,zY����Yg����]bj+J�z�����ڶ��T*�+_�8)�̬�J���n��3�29��E)����kh3vt+��6gZ�8*�Z�T'�*5v�s��T��mi�p�1�
�[Q5�
E�5�-y�+��\}V-�]�jPZ�n������&�4+u�AJz�,&h�ٽ0BQ.�[C']
\hù��a���!��;E�4�mf�w<�;x0˖F����\m��7{����aj��M�g6��L�(P�^�5X���T�.�j��6J�n����f�A��3�����)�:����9:���a�ݡ����KM����s�i�1kW���w�~7��3j�4N*r��ŊWe�'��9���U�T���h���7��(�����zEt���(�/u�gw���CӶ|=�(�����0�R=�}�Q����-$�fn�w�c�3)Y��E�=dun��3/x���<T�;[[q7�Wp�,��\A�ra�d��;**r��&HНA�ڲ�7n��8g\95��'�9�F���k����&�O&��'e� �pb��k�ڕ[Y��$�*Jk5ʬ��3�֨��|l���%��{�}޷����J��6U*૦�c
�����9ees�������A���׈:�Hczu]]�TTUUQTQEA�M�DAUEDLPE%APTAP�%EIE35:������"�*f(���j������� �(�*"��� �������*�� �fj$�0*jh����b���*"j����*&��X�)�)�
�"��(��&�h������*�%��*�"
&)#1ʨ)���Jh"("���if���"&�*���"%��(�(��J����h��)`������)��i�ʈ���������fI"����*"�Z�����b*������J�0Ȫ$����
	�()�!�*i���(���0*&b���������X��*"�"������(���*J!�)������)b�"I�"%��
(�� �Z�i���&�����������������(�j���b�"&���&��h"f$��bs2*�j�k>�{�<�W���w��ֳ[̮Oq;Jl�s�^и�#5<��y�4�.��;����œ�u�\���e\g���sk�wS�;��V��W�#��#@@�'�0r2�c�Uq5�P{���+��\��2P��v<޼W$%.�4H󗞸k�9r��۽�rQ�0c���aT��72�Zk�d���f1psO7�r'��;�GY�#/�u�OM ��`&O�2�#~�(D�p�J��
K)����w��v�{�{��L��N�O�S��eъ�ٸu�P��������s�P�ID��-�Z�j7i-�� �S�����J��9�5����sqP��&�bau^ESc+'֒��K�<]RY7�4��!M�:�)�@�N%i��"�F�c�g+�sݷί�FW���em-���8�7���/	f�Vk6�2. :*�9_f��WZp�wc**�/�PQ��b�ɳ�����*�k~�|W���������z�K�k�^3�d�k^�mm}>�<��+} ��ױ=f�zr��oӋ�h��_��̤{�]
3�#���ӈ��tEF󊌸Z�x�Y�X��~~��X㾳y�4�[^N��#:
oCex�� wwi�/��5��gfj��x�;ɳ��F��7(��M�m�!
ž�ܭ�et�Wd��w�a�f[�Uf 躻BN�۠vޖ�"��FW=5i��W��;q�u��j=���A��|K�������պ|W���k �{^�J�1�\F4��[������'h�԰�����g����[7z`ܡ�P����t�p3Jd�O�%;���B��S];nX]6l�[4��:s�9R݊�8ճ��"�w�<(�~�yJ��^1>,�,F+��;��:�n��m���{�8�R�k���$1q	Cngh�p�����(2f�"��!etM`�̇���UcR���ܞEh>�~}h!r����x��X�o�3��";=2�q��w�xY�x�VK�r�9E�)(�<]t.g��>����j9�T�#�x9�����a��Em�	Yn��,��0�ǧ�N#:��Yp�aIP�H���`pD��[1�8��ý�+��F�����U<#*�w�Upw��N���yJ��yT�0j6�������£鑂(u�d�"��+��K}'Mw:��yMh�e�ё�\C�Qi���J�]����"�v���� R�|���a��������|�!>�W�\-�y-�ꫬ�G)>���~�v3<�}��3�`��)
l��nX���=�,Q�N�*�����3͑����`Rwy,�{nI[�iR�g\Sq�9eV�K�z�mIsk	�f��G�q�*K���g{��7sk�⾵��]�.�\�4�kR��ԍUqp�M��SmC��g��(![G�y�8lv��(�<VU�l�睭Z�������\f�k�ځi�Gj}�``~1�	�ڳ��@�6�5��{]�S��-��Cf�䆻~������Q��A�N�@����s��5��E���w f�0�v[�!c� *�����֭��s��Ӓ����4ȳ���`����-#��x�&�����J�[7�\�1��PLh��Y��B2Kf�6h(��c��-kVE�=��/��@>�N�b�4��\��9�dp�圥9V�򒗝a��U����_���z:|��6)��ج�=�����a\wqp��?;����kҘ�K��/%��A}|�cC�(��x@��c��c��9^���ʮ �<,j�v��\�;Qf�%a�I-^@kt��Z�F�պ:@,f��J.}0��:Zr	CQ����)�@�z�zzh,�����ʾ�j�b�n)�%"E�
�[$*X�"��>S��{zs�i�V]���%J�xg�Э�yƊY�M�F�1"s��U-���y([����[^v�q~{4T���ja�Ya쫅K�V�kk���ΰ��&�����n���N*��;f�f�ڋ��TVk(�7fb�Sn���=E���:�Z]R@�7;����!	��:��;�w]����Un�T��Գ(��;�����B�[|$\+|�FiaQ9���\�@"����Į�dsn�`E#�O�z]�bc�E�QB�=/�tƭs\=B{�*C'_/5����9oCt�⚯�u��N ���h
�$"ި�	��/+�Ƅ����(꾷g���L�.W���aL^�����-��"��eZ;��$�����S���Zҧ(�=v��ݻvzX���8���U/�ȣ�p�C�n�)�s�$�$u��墕��{7��絙;�h ��g���I��
êP E�L�*<�]�C&IaS�݆�E����u��'t�E��t߅*e��(A�n��9U������J W92ˑg�������-�^�dXk���|tK��,9��f��cA���p��Yvn�p�ͦ��o&]שB�e���3-<��e'<jbU�G�]���6n!N��g�wy-]|�}�j��I� �{�#�o����0�څ⒒���c~����\���'E/���@͗˫�3�����A��wt���EF�t��CV�z���{��V�b9\aj&d�:,�Z�+@��T�PJ�K'm�V���^��7�֣�X�6_8�]Z�*�,ؒ����Z�Oa�A��.�(�o��[tV{��\�X�ॉ.�`݋�	�E�l�����X�Kع��nT�.��l��X�fK��a� ���tp�'���W<��!�L�4��ޅ{z."���JP�]��g;?:0y��Li�]cD�cC��2E�)l�{LEB��"��a�<�w�z���B(���(������c�*�&cU�S���D�KrY�Ɔ:
}h`���q4��]�nmSg�R��ԇp�T�*	��z�TqS��Jq����q"+��Vb��0�d��vq��V�Hq�0�l5�h`�a`>�<C��Th֎gQ�t���/���v�����Y��s=V��C�}LF[����	�T�NJ$�9c^4wЎ;;��Oln'�l&a�M9���:3�O3�r!�1B�˳n�*yFd�&�D������E%��$+S�a�d�G���X{Ӑ�)��Srr��8sqP�
�5���>p9�rŵ$���(��<\U1ՓzP�N�*!�)��\4�	ĭ !��t��!��Ɏ�uyp��1RǭW���q3�XXf��VԠح*4��
�tmi����WUX�&�됵{g^+�*�����Y�V�䗘8s�X��e�+KW�2Iۿ,��r�q�5ަ9e�س���2�<�3�n>�qmmtIP���MX��XG�q���;^x�T�ft�]^Ox�����b*��m��ڨ��������A�I��۞��;6r�Wn�Ӵau5�+l��;�nvgO3v��|�T���gn9�+^uȸ`w�"�P�ً>qp)�O������Y:ǽ�n-%!�N�����~Z�~�s��7^60g��2���.�e9��Iu��=z�ڧ��9��*/f�������������1�[���(^�ؕ��qU=1�%���Yf��P�P҅�񱜮��֧�MJ�)����#"�1�k�^�9�6-�ons�VR�nC��o߂.Ȱ|� ��'���y@�Ѓ*^��W��ܞՁ����94��\��+;t�짹!�(J~��>��B�u�^%a�a�Y��'c̎sR�^u���(YN��>��}h!r����49������Çkv�+�-�ϛǪ��?s��r�tXL�/���/>�Q���Q�*H^w���������=����eJgz�:�(e#>����� G{�OtͪU9�=h^Gtw%���F� >IÀ-�f������������6K�sU�T��BL��u���Uoe��*��|f9ݯ^c��$4�E��(k��Tgwr�3��B߹�Lu�.y��0÷�]V�N�Ѓ�O��U�s pjg\�x\��Kjw�\��S��LJ
�Q.��`�*z�纩p_)��;��C��h)��X���&ѧ�yѡK��.&ь� ���|O��"͎�_ϡ[]�˳�9
�v]��5)8�܊�H�tx2s�=d
U�GAh���u�]�\O#����>fw���I�轹�6��on�lt������~sm:���h3f�T��mO֕J�bi�!��B�:Ǜ�oy�%MomA%�,A�N�@�NB;	��,%9S��Hb�;>�/7�C�zJ�3D�٩���`�v3#�}d�D8U��x�tCLϱU	����mr��q���t�k�ҕxka�u��(��Y���L�R�r9��P�����̆�Z�>s���7��J	��r�`�"[;�4\V�~�b�ZՑ`E�6��fuV�sơamN����dp�z�&}hNRR�.:�OR�*�}N��x0��zM��ՠ�b��k+͢^�����6����0c��ąlJ�(Մ�hj�6{Q��S ���};!.W���}�~�0�V�r5ܔ��+�,:��n �s;����f�`b�m�Z�ܻ�s}ۮ��Wdj,u�.PN�:��i��u�~��`���릫}�3��^�[4�2�,g��K�	OR��t-" �#S������՛H�}^H���t��h��-�ۉYx-t�9%a���_[r�V�l�]��W�f �vP����[%�o��i��P�p6t;�PY�x�Â���ј2��[y�[��%�)�L�w�A��#qL,6#F�����C��u.|�FlJݫ����/��_t�<�I��K%@�%idjU*���"��
��	���[q�r��<,<J�?=�:m�g�M�O ��B���8R&3����}fVOK�j]1�|�z^���]����n�+�#��?u�<6�xW)��Ȑ���x��f�[պovkZz�j}��������Cu�Mpв��7˳��-�n%�#�<NL�&�!��5F6�n�A];�JΨ�� ȧ�vhhCuʛu	U-�r�zzdS��'|H�Q�	<�wz���=��R�^e��ӊ	Y��.���t��J�rd
�r0ד˸o���7aԞ"�A��皽hߡ��\䱕�k6fV9���fKr�q뷂�8%�rN�/���PC��푕�=)1׻��ؙ��;�l��˛��v��o��]������qr㚲Όm��P��q���6x>Ǆ�3
�ݝΡ�![S�o�Ƒ9^��'ǫ��P_Y�(X���9 ��AA�y8� ��%i�vG^X���s�w �}�)J�ș�i���k�w���E�Ɲ����A�oS�@�[��W֫`:{�%J�U)�i>.�-�<
�te�5�2e]��9�Ncu�Y�z��ju�Q�<�汙���F�Ѱ,8��H��=�;�%��h!�~��9��x��.L����Q����V;E��r�s��Ť�@q��ʎf��b,"i���]���^������5������7z���"`�#U>�)y:�9<�*�Y:zs��eiȶ�*��R(�`�U&kh���{-u��\D�Eܺ�j.T
�"�l����_T8E��o��R�@�`��[��Y���.U��]\ ��̝1g��
�UI��uN
��D�)a��!�-�~�])�A]N���y�y�^�'��&%��[RÚ1G��
'�*$GB���R���1�{�^�����*i���DPq�z�\+��6��:�e�ຌ��NJ"�
+�pUzL,���8}��B�f�n�������8����)O��ʽ�-ұ:w��CoU�=ס��f=��s��H°6�K5h�͛�*JF�!vet�c��r��j�t��5�Q��"��fA �h�bWN���bΏ�.�G�-�s��1�}�M�9%����##�������0���|�GC��#/�u��zi}u0*��%�F���A��"Vv�.�����s0F���2�ޕ'Fr���eъ�]�ע�ϧ�!Yt��J��b�ol�ݏd���S���!�� 9��'{Jzre0��c�����;�#����u��qUbw㹏]_EF�g*I�`�:��T�VM�B�0��9��h�c�Ó��
ZrŴ6{��̬����z@�b�ͱ^�Y�*���h��q��Zמ��'�蟛�@TطݎQ[�o���Y��2�.%��s�6�]���5�Z��h�KHh�I�~.�)M�o=1Cf��.]�gQ���8�<�8�p!���+���Ň}"��W�\;Mg�'dĹ�-NW��vˌ��N��o8����)�gI�g���C�i�ܼ��8ҕ�8����~er������W�u½�L����a�5T#-m4\F7[�<���]����׹L��9���v=e�t~H�W�����C�^l�o�[(;���cuL(�p�Խ�8C��U͒��3�E�PIng��k ܸ��7j#W#��싥������Q
�F���f-8q]d�-+�D�B�Y����о�t���EU觏�����V�\δ�r���K�ѷ[�{��Ԯ�_+ХwK�d��b�)D.�ٱI>���gu���-Uڜ0Ы�rv��}�=}M.�i��0B9*:벏M�H	Ǥ7�e|�Jc�ҮӼ�y�!�u�6�fVoRmj9��Q��H��4P�jR�;7�*Pڃ���z2�se>�8��m#6H��!����r�_D`�6gL�qɩ��;��s ���;m�b2j�gS�PY��*�=�P{2�uЄ��c���Ug��b�X��Mm�
UjR@۬;��I*<[nn�#)VU􇴰���5���Nd�`U���<ԼE�3�UF�Vj�9r��M���u����ҁ�jܤ(�W��4~OLk����f����F ,8&l��Qͪ�.z�Փ7(X���kY��������&�W�!�Ɯ��uQ]J"e-��(�$��� _�R��׊.s�o#�%ʴ�{�r��$3V!�I��m���]���2���2.'E��g�SE��sN��BJ+|9�W:���2�-]j�|�mI��ܠ �7OL&[G臉��6�j�s$i�ĩ��y���2/��cH��sI��0,:��-ijډ)��ʬ)�	ռ��4oi�Z�+X]J6\�z��y\�x{1�,���1�Tk5�(_�&����7�wi��3�[Q<��k�xᠶݸ���o�;|;/w ��f��ɇX�o���\�9/�c�h��Y�Ci�?��`j��>e�tT��Zl0��w$7jҺ �LL�.����ί�Es��'���2����m�9,�A�ޠ��j&�Se<��]��#F��aJ��:�6 �>�0RW3-tީ��ҁ�!Go[cf*�X
��ǴM��"���/k�\Fֺ��s;�b���sO/����]B�a�i��U_�Qp�N��xfB���ٵ��~w�{:ҫ�<�8k�#_���l^�v����1j�8��\z�%��O��)Ƣ������V�^��w2m�T3�"�5���2:���R�d޶�f�X�YeG9���jZ
�	>b������e�哚�~�Z�v����buUм�A��J��0_n�GKBv��ElPb��7l�[�u�`Z��J��/���*_�8�s�R�y���h�-Fe�>wU�DΔ{D�]`��Oo/ ���1�+���Ù��黁I�[+���-L�ӎE����#��Rț�[V1m���HR��r���yknG���/�i���(+��2��İ$gnh	[y�0���]���9��K���q���6��OKݔ�0�|e��L���K(�
��S���Lv�uB�Rtqwա��#3/�=5{u���IZ_ooP�
 �5DQ0DMTQMDQTPQ�3�DM5EQMELMRSE�$^FIQVa�D�DQFAfQ0��MS$RSTEM����VfU�PES4UL��SED��M?@a5ET�T�f1QZ�)��b����VQTSD�5QET4I%4RQDk��3
jh&b"��Ja���)���d���QQZ�jb��"�jb����X�PI11DF�2(�����"��Յ�U5M5EF�"(��H��*$�*!����*h
f(��"����j"�(��0�5eEU%�&��"��(����Q��ML��TSA�����
-a�U5fUDUDM�LE��ՁD�8�SYD�Aj5h�
	��Ĕ-�L�s3$�Xe~�� P�B�@�;豚��{1�.�(-����94Q�oZ�L/FWy7��{I�>�!�׷Fq���Z��L�O4�n�DG|3|�Qj}�H�M#�'��þ��`#�a@���J��N�X�P9]5*�^��cC/�,_��ZU9c�^\�\s;Eߤ�p���� ɚZ.d�m�g<��2��~�d!^��K9C�����v�/08�;�X�n&g����\Vɶ�g3X{:"��@Ѝ�vI�]����L�7�OS�5q	��7*HP��K����Ÿ���.$�uj�;���1EO<�G�b��Dں|�p�
J��"3_�=j�ww�-[T��E��<������c��g�Ά�؇۾��4�����7cqwylP��D��E�T��k+%�����R{~S�+�}k����ߩ*�C(b�v'���%�B<+�¹cn!�XXx@��rx��Ջ����c<�.�>w��D&���퍻��ٛ�Ō����l2��7Ca�c7ή�S���@B6�k��1��k쩌,�!r8�׺���N��PŘ��MBR�TBuJ�!�N��L�%r����H'�N����-�Q�ri�%wvU�Ȕ(ZK�wX��'O�X���lE�G6EXM����՜�n��8���k�uf[ĳU��I�m�Iv��E]��٫���-7�7�!���Do�XBu��\���X�m=�Ėdkv�]ӒRΎ�4����^e��tI���ד�P*!9C	�r4�yw"/���c���e��X�8܁�q����r]��٦lh�����4��+ОR�o���v����MU������뉸�:hZ��kŭ�d�lP�}j�k+ϗ�mAsc����0�އT宛�!���=�Gg��� ���^�b��`e�AZPU��W�`��s��&+uOT����:ޱ�'������1������__�pNid���h�s�9���*�^t��t�Ƞ�*�3Q<���t��h��)�ˉ��&�\�
fѬcUƌM�W��8:�Z$[�T���Y��6�X��a�N��|%G 6tTJ�(ܡ���uт)�t��I_�_�f��2×0��EF)��i!r��W��w�/f�xA�e�/K_E��x��38�=�����&��@��`�뤩(l�B��P���B�[|$C-�0(LSv�3;!ҥ����6���^���#�I8��뭣��\�6��E�0ɘ��_s	����'@���{4i^"���-�F��hZh
*� `�ktk�1v0@c�++�|_��~qs�6`v�E���;w��Nw(����񿎥*��ndWt4�d�eCA��5��37#PI��Z��� Gh_�_	u�m:���r�7���6���7�rɮ��]9g������W^�P��
��ү�*�5�,{�!��%���֡nrݓ�\t�CV��pЙ���tr�<�,\:Ȧ!�1��O�F�:9�6r͘H�J�-��{��0��Ɍ)�U��C���НC���Xf�IU����_e�0��7�ҔG��$�����gf���hs,+��N@��P������8�d3����/eN���W�{%��.��	B2���Ay��]Q�� luٱ��N��t��ʅ@	H�sCGy��=�)�ה�z.�[YACuh��ƃ�A��Fɾ
�kkwz�{.�]��XV��@�u�;�����/f�JyVi����늘��&iny�w诞�.��҃�ac�%c�C���Ek�b��&v�/5�e/�S���rI�L��-`:*���pra\��a�ڦ;����p#	g�m^��^����=43�R���Q\S#rt0D��WJ�-'ON3��=m�NX�(���r����G��$׈]?W� ym�+|{��ᕆ�p�ܗ�&���lz���l׸'G:��x�D�Um!Ã|�|��(�&����YE�A}�H:�dۣ�����.<�f�A]�k�Ek�T�b�XP]2�[����	7�Is`���O;���LP�٩7E�b����L���M��b*��p�y1P��IޒA�����kމ�8���7T#R_UL��R�hؾ�N"��=�E��Q{�w�����ꧪ��j�2	z�=mB��`�GB� h� W^n�Rׄ�{�"ձ�$��cڵ�^)C-�+!
��R*��6��:��\���&O�C���� �� }+�n��`q�?)���;��X�|�Eþ�]_���6��B���`RrQ���+���[��ˤ�M� ��
���?j��!�����O3�q�1B��y<�����̉k��s�V�FV�`8y$"jzx+��W0�T�8*4���M�w@N��ã�ٽr]�4oUCv����s�C�Q1=������<IG���U1�:�00��4�.2:0�8MW7E�4��8�ZE���\)�*+Ѱr�;��S|<\��x~Z���n�㤸��{���C��>��U�,�S���� 1��,xO�#zji�5��gG���wf�<� ₦m���G.UB5:��"����`-�³z�	��(��ڢ���2�=|��h<-G�8KJo鹡�u�p�No=�sx������L-s�C,���@�η�'Pچ�r�f\�}�l�s&�s�}8٬�oK-�S���W�����c�������v����!ъ*e��%�te�jS�j�ԙ�9Y��\F��p-t��qQ^X�p��<NC84V����ݬٛ=N�nw(	��z�H��VF�t�^�#qt6D��z�P�[-���s�0�U7ۅn:̔[9�Eƭ��C x�f}Tѫ١�/6[7[(2�P��M��k�MX�I�}]Q(Ïr�k�b-�v�{����,"� �) D[낰k]^0e#���7�U^j�0���5LPi�-1��;o�U��<	;>��B��m�;]��yz��y�b��E��0�KS�-�^�v�/1pzO�=s�����د`~SZv��M����=������x�c�q3��>����F�wr�*$Tu��m����W>�#a�:1����21�`#�燹��ț�|�p�aQy���'{r�v����x��EOs���DZ*U��Y�K��Tj��r��Z)C�� 3o5إ*�k�"S�PbM�������Zv��v�`T����I&1ɰW�����ݯy��dB�m(e��Ha;�3GtH�⮥ݴ�@��Q#/&�5Y���ye�/��ކ��_)��/zچ<}V����ж	t�U�g�w%��oXn�qM����,���=c���Y)�� ��x�G�L�r{>1��x�����ڽ4a�8��8�;gG'O+�6�e�����掂����u~�U�j�K,%������9歩<\o:���0�:�����na��Wp�4D!G=P�S�Qπ��Mz[��t��#C�a��:n�U�&�)b�P59�\'@h�3v}Y�[j�Sקh��5+|���:��H�)԰��{x0[,tw:$֧��B�I�O20��O�sV��yί+d8�8~�D�>���@�K��#�i�����`[L;��@��S,�T��;r_�G�.�s{��Zn�dxث%qt*#�2��1�;�D�w��V�X[{�z�`q��ȼ[Q�r�]�z9�`~�X/U�f/Xf�X����H�w�F뀖��WW?E�
���+��;83�2��,E�R��!��\3m�	��[�x�;\�f�KZC���1�Y��u{�<���t��E�����G"*��j�5*��H��Ꚅ�J[.l�`t!��Qۚ[]@��DݍhM�;��Z\�R��^>k&�%r��%[[������1PNY�f�̛WE�q�H�)&0.�K2�D�Ղ[��[=�a��u���ĝ��l���]������+&��Ϧ�@>���(c�t�sG���f���3�
�� o�e��o��N��|%G<:,8�3j��5���^f�t���t��)jc�ȭ�s��ć|����B���-�|�:n'���d�0���{�6�3�i)m�aɆ6	`O��(��r��<'�˅��]���ᖼ۵o� ��{�ѷ�V݉oS���>ʑ���*�
��j�f������ǫ�����s����iWW��r9vo��p��S���hD�0B�ba�5�Wq�	KKՠ\.S�_��cV��-9��q˳�β)��� 7���dܐ�������rK�!�hL\Qӓ^z�M���:��p�b�w�{O���uoPI$���粆=�X�$��B\���L��F˖vl_�d3^�
ʁ����6p$[TV	����Y/��M5\���9��d��R�e��| �/��Af�Q��atuIq�����ҁ��� �RW�ʸ�6a��J�YB�e�"Q�rψ �B7�kt^�H��G�6��k�rVp'���AD��ovq��B+8��:�\��4�芏[N���B0��Vh$���}|u�M�	n������.��gC]�v�Q��Q�L}C!����0��ӹq�kj�:.sϻ�EE�z����T�{���N@!�ԯ���y����H�zv�㈽���c�Dճ��\�3&���z���8�بYQ���Xծ�7���>0:�,:�����&&��hw|�kw9�����6�����
�ڮ�q�D(�ʄ:��R�&ږ7OZ��a�����Gh��GVƻ�ց�%���b���l����+ӓ�\uMGs����'�wv$�C��?\�`������y�����P��"��s���@����b-��1ؑ�rw�\9Ѻwr5�.!�Vt�n?R̔b�xL`�
��c��P4U��qY�\nZ�E�K�p��[�:HǝP�S�A�/:S[P���X=K�X'�KД���d-T8���t��׬B���B/�~3+;�������+�N��!|����o<i�����z.���J�Ϩ��x���;��o�H�;����wf���A�̫�n��E�f/ ��{9�{�eo� z���=A��C����:�=�x�h��W�mǦ,Jq3��W�I�2�}��\yt���>�14H�'B��-��!f�Y���z.�^/�NR�]�!�V�	���,��z��ܫ.$E����[d]e&l-�.i� �![��,�v��Uy��J}	}|pI]e6jIӖ��\�퇯Wu�-gtZS����-ʷ�\�炸��:�`>��phA�OB��뀝1ֻv�WA�ƚ���%܊G�?+X)�J���4M<ഗK��9M�k��	W�V��5�s^N�6������0ffs��Cc��{!��P�-NQ�6�D���e62���c�f��V�ո���Z;�������ّq�P*��eo��>��	�k�Fň�KRg�7�)n�䳻��X�����Nэޘs�TN�,p½���Z�F(=}�8��n��7���|��q ���8�|�_���c>�+�`���t�"m9�x��ph�3�Tº��z�kW���24;m �j�+�>V=+#�0��:"vl6�DZ��h���36���(ZJn�ݓw���fm��ѶU��¡M������/�g�P���ּ��ҩ�n�N<{+t��Ǚ�������C��7��h�b�"
-��L�9�'2�ۣ{��MY+O�H �U0��1Ca>��m�avDSܑ	Cn=3�Y8@׀�׆�Fɾټ:$U5(VM��!�H����;^:��(ΥY�~�@f(��d�c=��v�{5uh�蹯�>����`�	�q�}���3Wfb0�B#���,�r�W!M���پ|T*���h@y`������E2��T3:�����h-,�m��x'����H\=�ۄ��,o�I�QU�9��!���Om�T�Q$�N�D2W�&�@bE�v�_xN�%�>�#i�a��S�٪]՘�*JgHD��
�ĔD�0��"����WӾ��Bɗ����Z�zn:8.>{jt[E���v�<<NPgV�EK��E���/�\���Upf�ymvP�A��ً���t����Ї���^ye+7�u�O��Gl��R��Qx��Ձ�˫Q�O[��oWoJ=��5���gF2�q��O���Y���tH����5r�ʛ��y�7:쾇��a�rt��\"қf9����M�sk��c�����
|2z�]�?H"<�Z{�#�z�.:�'����pIH�	��dq�p�������]eQ{[|%*�X�� R�ٞ��txຳ~>��2Ks���B
s�V���ǲ��c]�����gb�*�\5�r.4�8]�H>�p*ס�{���,{7�����mR�f��<�3�qua��w�w�v����������ܼGV��VY��mv�"�$5������(���]���Z�V6d��k�0VR�Z�5�hw�w��
��&���"����هC˴����W��C�f'E���N��,I��P��vs�#����1�/���5K��mk�.��b�wΩ�m��v+h�TK��%�p�娕�	��UZTFֈ1�ֈ���[ق�HSMZ4槁A��V0�z{gƂj�>yƅ�[K���l�`<�aEYǚ j�u��f�`5�ROvXb?�1PcRtb�V�L�o�w�^o�N<Bϭu݇;��N�p�1�t!]fأ�5�F�j5�y��r`TaV���V��:in�Q�L�� ��l�l7e\��>Z`[%,=�Ϲ�YQ�+5_I*�T��A��Aj����FQ�q�t�!'gJ�mMu֍�P��#�m ���aA���c�K���&�[+�^�,6�fv��)�%/�g��~�^����V�[�`��\����W��w�=�7l��(���'q{&3�$��8&)��(�\�����-�Vh�6@�__46μc9B�;��*C��5��8bK�as��,�\�w���� �Xb/5f&�34,�ive]X�We��>֤��st{�$�u�f�zW�$�-�
�RF��V�V�ѱN��}F�n�N+�]'�&BF]ctyJ��0�B�� <�)K�7m�@*L�����S����4�̝��h��mj2Igzf�sxjG0b�uëM�ݴ����>�'�v��JC];칇x���*�hk����K�f��2�+v��.�� ���%�u�1 ��9�{Ő�E�Dʱ��Kuw�'���Ĝ;�怫���ީ�4ӛs�F����ȸ0,峪olO��\];5V��; ��lG��6��V]��jh�aj���r�\V/'
kz٬��6N.���%�MJ�V���^D*i�r�\����p�r�)e�hfIcs��z��o|��}|^���wTCOΕ|ʴv�c:ƅ���2�e����+�۲�]�X�6-�)x��]�:�\ܮƨ��P2;���3'wKu�������US��t���4�U�Z�8���,C7.�}f��{�fM�O]�r���Yǅ�}%"�����7��N����I�Z�����.�aC#7a@�WNM#hbhT\�^�z�d@�=�F��>�����N��qeKѯ�V$ۻS6�0��h-�X���+�+�R���+Y�;�9�R�n��=�t�J�57���p%�6SW� ���{u|ǫ�1�x{	��1a�6��Dv`W9}:�6�j�sAL:�Ne��s���v�)�o4���Y�n�ޭ��:p뫙�v��c��/{����Ұ�۵me��x2�`���h̤�)S�W,;ժ�ٷ��z��}P|(
��*��YUV�5��HT��"�l̢*��������kY��FfATQ�5�PT�5LSF��j�I�*"���+1�"�����2�&�0�*j�"l���""(��2*��J���,�e�2�����r2�"�J22�K��� �l���,�+'*���0�0Ț���',�L�0��0�"��̜�3
�,��1�,1�ȋ3")��'"�2!�2*��s��)���"�Ījs��ʲ+�̠��!0���r���+,J*�h2p��2��3	��
�p�")��#
J�J�,�����2�2����,�*�rs0�r��\�0����h��"��̤���(�+32�3
�#��"�Ȍ�,̣	#+�,��r,� �J��9�h,��e�f�s���C���X7S��V���
�ibF�Jkd��PSe�w'`��܇����P�ۼ��Mwu��E��*��۾���
i��&Q��-��ch�	���U�]7[����7��o�����/=�®�;���|i�L5���R/:����P��g�0�=�ܭv=�H�W�+C��vp`L�V�1����o��W��u��)��r��K���ڱd�A��Ŗ���#Q<��ȃΖ��S�=����GM��\㐹=�˺�q2�3~�ïE�c���8$yl����	���3��OO#�Sk�e-�V��,�'p�N�rg��S�U-*1L,6�HT���r�b��NzL�_lPfbr�|�Fjra��@��~�::��@���g]{p��A=��Mrp^����=o�h�$jeH�}w0"���s>��꜔���Kں�~�6iSW��t��S��5:=П+�n�<7�+�ߔ��*�+����yf��Y���.�7}aW�JA�ξg>�/���	�^�n]��ylXsq,hxqZ#�A4�f�C�y�������K��Bx�����#�7���lSc�q�1A�v�\������?G�jv�zi��;Otj�����4Ŵ��	ɽP0�ܱ�Ŭ�����>�I܆��u��ruAb"�z.(�'�l�A�ܬ�Ηݫf�����Cf�TLQӓP0pZ�M��f08��E�P���:�_�[Aɰzw�J?i�]�ؚ%�y��|�RuIp��bƺ��qA7d3P9��uJM�݂/)�q�a��}��*@��ӂ�e�<�v��R�ф�e��<��"�}b�X�Kn��fTe>��p������ŸO*�LهТV��C7*��^����_�y�nc�dIԚ�6�/vKvkz�)kW�ZM�s�"c�ĎxVӨ,�����+�΢�ɉ��z�znG�]�X4���C!p�VՈ�p��{HvAc��:�{T+)��S�\��{Ǟ�5T�8��F�J�ڧ�Q��W�;��R�&�ڦ;�ŭ�3T=t��4�Q������^!�/ӆ.X�t�z��%Z������|�J���ӽ��Ӑ�&��ܭ�磬�.v�S�)��2�����r��O�cqKd�>� �ÝՎ��4�k\������~y��{�qo��s�suB+�����EU�7�0:��M.�}u�eQ�2{v���S�V����V���-Z�G�	ق�T�E�` J�׮�KVm�������-�T��L:�GE�[����K��/#��Q��\�B���\��){��G�u��z;�dī���v�"Ζ�\yd�3�tB�7Q���)����/�c���!�<'�Q<!T!Y�\���38�<������9A��!�H�ncx�
ϲ�p��j%5�1Yӎr�^䞌t���Ʃ����v�����Gqb�*����up��Y���{7�)�v��}|�t�D�F�`p�\&xƼ����Ω��!O3�s�%يv��U�w�Swq����)���Ȩv������Ig�ٖ:�`GI���+ϖ�����]�ыp�k�=�u�V�����v�����O}mO8-'j��_������V��*������Z�O#��^k�SH��q+H1��M���UuYG!#p��7���o�ʙ{[T�OV�᫖a��O��1�]�ّ~��Q	ĭ7���2ɳ���V
����8�7|�b�fE�wj�Ӵb�]@�&��������;Ek�"�Lƪ�1§Vv�yb�5�9v��ٳ4bm�F��p/˧D9����O���'F�P9�5;6�a׷[���=8��tH�6��$�8M"dC����&>��� O�%����'��g&0>�� �}�\/����^��1 �|�JͲ��I�#�j��y/S
�X��.����k��U��,�[۰�� ����$��қ)�ص��^��Mx��j��@�3N�<7�{4�������5T#/�A2�N>��7��n6�s]k(i:�9	��g8�ד�hvA�"��4j&&6���^��T����<=mm߆�/�j��{��cULcR�ez��m��/�g�M4C1
@�(]WA`���]�x���v���׺t�PD�A�J��΢�}+(�L.ȧ�"*����v�_^�橊2��uC<�Rs�s"��p�f(�<n;l�+��b�
t���>����,$��(�-TK��U���GHN>���F��iv��xl/m5�����#o����f(�NĨ0kYi��Ɨ��OW��9��uc��p#+�2]�$u�P��A���,���<���t�$�|�x7�G����%��"|�`V�'`W�O~���~g%ѽ����No�������7�sӽY��3�ӂ/�۾�)Y��a�{��F��T�y�^'���kDa���[�hٮS�gc���GN�K)�st�'���%i��uN���JT�d+��^Jm��T��,x��K��U���v�8�����[�8��}x���V�d����=pe�\��/��������w3\�Ffrd��b�:�v�ɩ�G+"���ץ��"ۥ-�)��W`j�7:?�Od2��w�!]���nuFq�l�yY�ϯ={���5ܫ�S6�(s/O7Cb���uv���ed��ݩ�s�{	��πGk�k �+�݈�x��o�	4��
ʁ��Gb�����XM�; ����Y���c8=�m�Pp�n��j�ݝf����'S����(�Y�SVu��/gM�K��K�r4�uR2!ϥj,�\��)WJס�{���΂�2D�z's]ݺh+�]=H�8 �	e-9��Q�:�o��Κ���J;2KG�np\�����_=�Ca�R�py�0R֬�ǵ�3�_g\P^O6�+7��7-Pug�����8��)`����f�Y\�S�� &Q5mS������\u�e�Z��)r�jk�=7/}�ٿ%Éu:�'��B�"�ϵ<���Ζ���anE�c���2�Ox�s� ,���[m���o ��@պk��*,�H��L߄��v���
�1GD�˧O:�����r.GF�*��A<Oa�須<Ӡ\�M^�&�ɩ�o��ma�5�6����	]��r�����*�@�q(��=t�+���D�����˞ҿ��z��j_%>�H��\1�9EW���9g]��w�Gwl���>�DB���u�a�r��}�MT��}�qھ�+�{��]�.+c}���z%�ND5��Yta�8���OiW&x+�tP��(��[���UJq�һ��{j���V�V�����	�����$oݶ��ݘ�(p�O3�!�7���]�Ao���V8�{GJ\��9t���V��-���7�+��`�5������:�]�;���3��f���ԺcVÚ��5Q�r˳��-�n%�	^����Z���.L�ռ�� ?+�����k����P��<u]:���,��>�]�Y�/aa�q���*�'���'��N�������p�� �s�$�7"Q,�ؽ�E��
�wTR]:O���"9w�uOw7������yF��'�u��^Z1��R�C�ٿh�CǍ*<h���)��(X���,�H�P�J Ts�2�<���GjP�u"V{:�[��w%*ҝY�[;������0�ާ �ZՁ��Om�g�Ś�5<�5�U�jbQ.��C;޼�>���rԃ5����׬�GQ��o�����D��COK4k<�Y[�[ɑ������wD7J�dV����V�b�����#��ͳ�O�������a��3׬�+|.��f�R����4�v����g��v�Ʈ�:�[����å�&�v4[R�&.</F��9&�ntnA��(��M�@�#5n�\�V<b�������%�ꤴgqx9����8+��TZ+�TgF�������^ԓh
�"׭�J4#]�w_���f��i�p���<���D�X< t�h�Z�ʷ�s������K�M'�״��c�Zr-���}�`�fR6Ϣ砸��z��vWg�l�3���(�0�k�c�J�{�!��Yॽ��|��v�R��hK�W��`�~5��r�^���P���r6ֽ�x�'���C�n��S�C	z�����08�U�'F��`�M�ٹ�]�z�RebUg�b��>�����f9����.G]f��X��[yR�t��0t`#�d�R��)�@�,[�R:!�W�N�Q��e�w�;�����L�c��5t}] e/�	d?j�JT|���W�zd�@�Yǐs�����˳p��C�>ۘ��MD��bX��T3�ؼ<=���ի��k<�|�[�W��s�44pr\�r�TC���i��1QĢj%�W�;����/��K���E���Z8�r#,ė!�הV�6j�� AR���	��#�n�!�P;r�oI���g�������S:l,��-����h��EJ�[/��-C��<_N��\Sd�}J*��!��Y�eݩ�,tn�7w��d�RN��W�[��\<��\T���c�)�tdy8��f��P�%W+!��l�{O���rX�&��{Q��Sfsy~fo����v���ڐ�����	ĭ"��]�"Mh���R*{ޛ�Ms}�^�`��g�,Ǜ㡗dXo�	7�����\<��g�ۺ~ٍs9
'����#�qg���z�Y�>�!��>x�����8F��p-t���^X�w��ND@7p7n'9�Oq�j�&�%�84TF��*~Դ��P��+�5~>��U�^<7�;)d>���w�[�L�NL�~Ǯ���s��9�F���B�X���k���WPT0P\�K�\�\���;6�\�!Ҥħv3!���.1�k��Vܮ�U,�����!^S�f�L�s!��{�j�`C��W@��S���Ѓ��T챇�F��=*��ڢ)�H�k�y����]� @�|���A~��,&B�a�aϣ�^�=�üS��	�u�;a��{�5v2�z�;����=�Ǒӓ�?I-�SHV��\�V���]	�G=�S���e�Y��I==���Ň6�8a�ޛ�N��[��ὡܓ�uӛ�nS�0Co��準������ٺsd����4E����]��b�g]�i��ԫ�kV˜��-	���.�����w)��u+&C������w4��EV
�����������C�7���wr��rB�f�eqJ�+���T���`]{��h�f'�\VjI�ݖ���z���hu��!V8�z�<�x��쨹�JKEA�&��^������pBԭ:�O)�Ca�W��ʣ½�zǝ�( :R�MFy��{��ж��v��y��L�O&ό_gw�[�ϑ�gCN��,�.��,.�O9<Bn5N��\oz�}�N����ڄ�V��w:��ͳ
����1���bN�bp�ګU�{��<Xx�| ����jS>��J�V�uI�g�k�K��P.��Ĥo6�\��u�<s�:HV9��&��%�HbCg$�{{x�f�Gs�MF�Ps5�u�rh���K\�ܲ��q�}�S6yw"��p.�:@�5�S�ˉ��%��g����	����c�n�͉0Kg��s�ݍ�j�qج'�pm>P��WA�!U��r[N�̋���	;e�9��~���2
ZՑ~Ǵ:�u����.����y�����+�t��0#Qш$e�Z�Y&��7���.�\d�W�SF܄�7�]��p��55���:+��|�ֵ[_	���>����U!.�^�<�6��vwK��h�Aⵍ�۶��"]�X�x� U�2	|�K����;D6��N]���y�[���ǼԢ=�ڗY���Wp#Q^��
�'���	�J�����*�l*�zl���V��l�����X{c�̳�;�{L���=F������)��ʩ�<�i��ah;Sܲc�}�[X����+/�d���
D���[�&+��*,�H����	}0�G"��fv��O��E�ƣ�:6T�GI�{	�!lI�\���-*1L,&��ziKpkW�o���xo9�
���/zq�5
ˣ��'���3�]K��X�O+�	~�n�dn��=g[��C���B��x����>ʑ���hS�¶�'p�ȳt�Q=q�I7ٛ��EB�N��R��)t���V������x�]�N��h�z�����t��g�����Y���poǄþ��aK�5l9�-5Q�qܻ;n��t�|��nF��rV��]��38v��x�OJ�pB6�B��g`hA�N*�p��Thp�s),�;139y�]4�5��EU��j�;���a��'��Ig�NL���CU�;6/۪�#��������U�[MJ��ޭ�c��N݇�XltMd�zY��o��� ú�o] �#��!���K�j�v�Ӻ��#��kl�L_p�(�#J��n�s/�f��*�+y�Y}s�v��!�� n�����y=����V]��ai��Uq�]@��n�7%�o�����o�{-d+*� ]�����yE
�;�㵺�[�~�ʷ'0�8�˻L�d�Xʙ�-�0�� xq�F��X1��*�oV�m��i��ac���T�B���a�D�ˬ���+	��;�n�T����rFc|x��-Hiژw�v�L6�|���=�Ŭ8����|�uI�`eF9;�h��kөƟN���v�l�5���h����'�̮��2qj�o�5��xj�k��P�m<���!�zr�YR�ʛ�x�*�v��b�L�(�o�c[�'oy࡝�YFIE*lMp������j��Z}Ƕ����&Q	��LlW^>b�ͫ�Y��%FTt/'�h�+�۔��G[*�t��|� n]����d�p����'�
]���a��O*<����W�ou�LXee)4�w:�K��:���y ŕ�`��v�-u=�
�����=�I�SsC�XWo��e���"�5�*m
��끆�g)�a`e[��}r�nڽ��L��yZ�P[���o.�ش#��7[Hn���:b2wf�e��[q�wE�m݅q��7qU�z~U����z=u��<wf8m��	�.,�T���X�������S�F���h�Iڍ�8r�	�[EwX�7���f���*.�'}tY�����C�����F|rs�,�+��u� ,����Mj�:����v&K�6�/��&v�jv���9EڥgL�y�(�m]X���{�k'	�;��wׁ̭�,�'�}cF=�WGx0�N�
Ժ�;�3N��F��0�ʇ.��U�2J�7dp�չ�wt�<��G
��\Yk�-Ԃ��bYлNl�(��8�"/@�Ί�C����FdY�ǙY��U��0z��[2��Y���ԛ�Ѭ׌<AT�-�'2e���ᣫ��.>v���bB�@��.��)��:�Rݍy7vHf-u�@�����28�g��)%7�q�1�ek�z�.�h*߲m��7|�'�'sf�Q ���i��bM�t�}Y�t�${j2VԖ�Vs�qZ���/~�����Qupgm˕�o����Pm����Z��m�-��v}�I��r���1��V���3p��S�.�de'�[wI�ϻd�"`4���(��gG��xe,ۼ6$+Y�2���J���o�pKW72[�$����_u\ꈼ�� qIϪ>��>�4�\:�ζ�WM�6:BY]r����4<멙���c1�5�(�N�����p��ּ�e����lV�,M=|�<�[�#y����pH�z����dv�Z����n�	�Kb��n����y��G���6a�dQC��fdQ��Ue��fe���U��TY�NFTfQ���Ra9fQ�FY�fXe1dXa����a�D�XQAeYUFee���9fX��FT��a���Y�Qfa��Y$Qdd�fY�MDdё�fX�a�E&f-4ffN��f.Y9.Y�d�FY�IT٘f%Y�9�TNQ9Ff9eSUPY�FfQfFF�Se�a�F`dSE�E�E�eFfY3�Y�Y�DfY�UVJeE�Q4�e�FA�ffՕ��IFVedd%��5e��FYY���aaDQE�NTU%PQNac��X�5d�U�PDYE��efE�ef�eT��D�	�>��@8w-��p�Ea�2#�HE�2��_3�MmH��=9Ӵ���k��Vh��U��wj�S��Wu���֫������K/3C�"��C~��N�Rd�����ɒXp 3M�.�yw(!���W)��^"k�����y�m�-��w�H9���X�@��P��Q	�\<�;S�(���.P��/����RO�֜��f@�3N"+��z�)kV��i7��w�/���Ó����`*^���*@��%\^�S/v��GQ�i���j��~�M�=�8�,`��/��޼���:[�3���Wۻ�dv�l?j�D�3�\^��߅f�B�\;;ف�k�	���Yگ&z�E�o��a�c�G��5|�����mE�a�.X��~r~"}k�Z��2fs�.D׼�.�s=����o�i��Ӗ�p�[z"���9�9EߥWe@�Et�@S�#��bg;{#;��,�VNt����������|���޾�\j|t*��Z<�U��a֦Ͻt��fU�p[u��<MF)A��{d:n��>�1�r!��L�!���z JaeA�&A�*��{�sݜ)x�S�j�eOإ����C狮��1Ⱦ����y�ϵ;��H���>��Luz�������[������72=�N���z^ثKZ7P�[�(��&𫏵8ȅټ\�9ˌ��$GaZ��Z8>vn�U|�����U����,���v�㇑C,�8�^�K���Hm�s�ubT����* 8T1���Q.���E���X�|�Eþ��:zp)i���Z��o�d��~kM1k��'%�D�B;��aW�kɮ�AoJ����=�Onz�}+��;���=B+l�+���D�{�0'$"j%�`��s�7
Ү^�-��z9�g.%��j����Xtv��k���i��1Q�J$��V�Sw8V,�SK��py�4�a�#�TC�Sa��
i	��#�my�P�-NQQ�Oa��O�G�Ϝ}�M��^��Y��]n�ƀ�w[fE�E@�'���t�vh1SF$�ߏ<�N����#}�U5XG��֊,;��gI��0I�Q0W'n�8ҟu�E�kS���Y�J�����r,n��:E��X�ٚ(o�]Xy;E��Sֹ��"�1Į���1�ҦC��4��1��u�V�~P域=�4Ъ(�����U��s���_I�ڲ�!~�g}u2v<�����1���y����P�qѯ'����8"��"��f��t�Vz���3�7ؔF���3� ��Xv�3c�;�G���ݨV��ی�d-�uVߩo֊���zō������]B-H�!�y�ۮ�E���Fٛ�Mp�¶]�R]�M.C�Y�tYn��I����,_G��}�;���nmk����U½�Hk���N�cs/cT�NŹ�݉�G��4XX�$���f�oR�������Z=�B�R��y��'B���`s���MSҶ�0�"���rŢ��:�L��}��[��Eܙ�"�TLLE�^�ȣkl�*},_�t���>�n�gٗ�inH���]Ք�U\����Z,��:K�$�z4�kK����3��x��[��՞6�U��r�ݜ�x`���u�"�$ue�|e$�zS��J��a���X���Oؼ2���{�E�uw���Y�~螑���F�_�b`q��1ux�+�b>�[f��}����ƷzDpqӕ�{UW)�A�Ub�<�d{��E�K���g�IW���� o:1/^%Ռ��ϹK�z��!�gF2�q���b�!�X\�kMK�,ٕ�û9���\IH���|q�ړ���p�fم�S��M�sngabaA�],�r]rgv֪��4#fHa��$1��b�Q��
�2Y��w����R�)���UGh�u�.�'�i�Z�(V=�x^4�@��NM����u'[��()BJ�J��W��l�:�����2ߕ<У�c؝�.��d^	�hԴ�kt�/�*磺�&]�B��X7�(�v��d��`�ޫ��5}�>�*���>��i=�k��r����)�2�5�Ρe_'��ܞ��NW\���������\��5���Wq�8O�yS7�yw"���7	GՆ�NK�����MEX9i��kst>�幋���[��5i�"��Zs�Ƣ5�\M��:h(�K�.4FW^sU��ǵ�_}�t��
JӚd}��\d��"��l6tO']��h�~�V-D�����/����}-Qk}�!��:��~�����uF_��	�	��~��Y[�pf���Br�k�X��َ�=��T�|sR�63�� ���ǅ��)w)���^�j�+j���z�x��y[�Oq��ڴ>Ⱥ�܋6M�㔼�<�OW����]�tV�z��1[�7k2�.q������XZ�(j9��n�AF��=��=4�� %-9EE齞pkk��я��<����T����C�a򘸇�^���a"��O�(�ү�g���M�C�6-����2�Uq��%�'B/am���	�o�h��$jf���NU��]J�'Uw�/h���R���bƧ?U��_����Uҙu�&�IS��*�S� �º4K��#�wEcL"Lx���B�X�<�ZQ�ڀ��=�d��0Ŧi����v�0U��������J�G	4ؾRS�5���U��S�;�u�= =����f�>�H��Bz�˖}G�a�.�Z�p���[�O�C��h�!�<WaȮ/u�Uٯnq_;\pD�@���&9��0�����.�հ�h��v҃�=�@��\�<�+�0�o�b8pp~u�LC�@�rx����|��P���=��X��;E��I^u��
C��ac@�c�|�/S�m�$i8��Rt�e�����
��A�o���r'�	�f�=��:᪾��	��*����.��#�$�p��5��oN�]]k*���\QlhI�n��^�tA�kv��))8� �r+lOm���K�Ҋ��(��9�:��(��x;�V�w1l߰�{,h;Ҡ�Z�.´�rlc���[]x��{�7m�\�T��3~��Y��T^�B�(��ڍf����P��&��!�q(g%��U<���o�VmN�^�F�B�Bxg��W��ߨJ�� ��2����q�t��
��u���"s-h�>��D�X%g�j)���Q�w��FY:��r���� 1��z�Z��J�C��z��E걐S����A�#W���l\��'�Q�Ӵ�N�EbE�t��%ܙ=]�,���u�(:tNR}w��
�/:3#�r�tl'V:��$g�+�$X�UϮ���*��� ��q�:<��,w���8�1�:T�l��T٦�����&+��>�ѫ�ئ,R��})s�\]B����t����a+׺����M�>�!��)of2:|�l��K2Q���c�*�;o>�՛�Ȁ�M½���Z�T�p��(��R�/h��Ƅ-��s�K�3`�*6%+�*��]E���}#��Um	�hHTHv�|M����YS��BṎE�(n`�r���l��[�����H��5��T�D8d5��F����3R�>Ãt�9��(;��G<$G"��R������Sr�vx%p��>�H[멁I�DT�"`!����k�P[�q願V�t8�bEs�ѹ�دe~S�s�yd�1B��z��=���*`jrB&��s�Y��/^�1����ʽ�n.�ݲx?qaj���М�����y\�n*��$�O^pU��}��Ց��0���g��/=(�*�3���jl1��:2��"�ƹ��yNQ#�$�ֈ[w��,��Q��+t���]\U0�e�1�H��U����"â�W��ZE����oEk�0i�>��a/Kvc�v��n�l�0"�jLZ'�Ԙ���5`��^e��ۂ[�;�R��t��Y�(M���a��Ja9[����n�֊���mk��Ӈ�̽��C���YU�g%�pW*�}�U��U����&\��mEO�v	Η(��}�/4�:��8D�Uڬev��e{-�x�j!��`�Y�*G'n\���±]��۝:�q~J�ѽuR2�G`!��!Z���S�\]:#��M6�j��.������GA~]��l�:Oz��]�C+;��S�g�L������㷵m������Q����`ZC�X���~�{�Ey������
f���f�"����Z��%:��'�
yǋ��A@���E���T/|�B��S];�܋��U,�0iawgA�s�MF��/�f��w�G�Bp�S��[�W�N�:�N�y�`�MSҶ�0�d]f�N�����7��R��ȷ霢�1�2\LLE�Qg�Em�x'���N��̱}<�7YN��kg:+ڟ����x_���:r%��bKG�SHV��A
��h��ʪ�0U=�^K^r⼺c��oτ���G\Bwr�d�����.�����=�//�#='��&ܴ`>���*���t��OW���\��dt���$��K�(]뼼�ݴ{S�5}�2��lG�"�n��m�0��[���dJq�2������em�Μ��Z�u����e!�Bz+5w	1vKa�Irf�'Sم�/�vVY�&�sS9|0݌��@g�"����6�rU�F�U��tM���r=�IW���6�t珞z���S�>G��wV�j��!�C�1<�
�>�N��ENr�N�K½��sZ*�o;!N�B.��]W
�S��[�۱`�-����\������Po�sG��kq�,�����x-�X��:��#�۞�ߖ�xy`�C��r�X?MD����Ulmf 6;�WM�F��}���%�<;��bA�{/����ñ���'�N,�uĔġ���n,Ξf��݁;�E'G8�N��oz6�ǡG8���8rp���/UE�k���p5cA;X7��q֜�&���$�=���nzQ��Of�A���[�#���Zзk3|��W�x�vT��:��8�/xf��m!}�/To����Duw�m>ۻm#�υ���w�/O[����2�]�>�_\���=ANt'ok{�4�W�C(0tl����Z�!.�l�Ȟ�O&�GooV 2����HγÒ:���59Cq>�!P��z����6NmWF���kZݘO��oc��%� a�]+�^��Ӱ�=S�R�첏oY��Jk0a���8��\:h,2�X6s�s����x��Wi!6,�/�҃:�����u��20:y�U^꾬q��_�o.�οB��9�v�r��3�ߕg�Em+�f�U�f�b*;u��óv�-[�	�7��[�=P�^;ݩ4��+k�����Fb���ĩ�g��<��R�;T���y�w��+BJ��1�k�9V�
�����t��}|��]έ�5���;ڽI�!�N�V���'wƛtbuV�|*{6_k�P{�U��ΞP�*=�f4EԻ��i%'��v��ee*~W�^Sp�����8L�%n[
�fF�{���=O�L��|�2����	:ظt�������{<��U��Ά�Ne�{�@��5���J��\o�{Qn����jT9�氜��k�y#��_�}m�[E�k�z�j�8	�L�t���-����?p@��Q���l^�ҩ�eqp��7�p+e��o`�mx�~���s��ZXUm�!�h[2�V�
Ŧ�c�J}6]��
A\0��#h�bC��reaݐ�\(n�;�%޶��X�\���A�ʛ]5A{��u���7�-؎���Eu�ͼ9ϒ�����fq*#%�:gm7�
9�7�,���VAK龂�:��ks���]r#���idz��.5(��B�Voed�y����{y�TBևn02/e+�M@׻ ޿}�=�K��ڔVU_/o����@r��֮��ŝ��<�7�$�X�O7�����y.�]�V	��TOl�"\v,v�-��ז�9K����.kn1��[��J�U�lYzWЧ��]N&����k!�1��E�b�s/U�K.��)�Ҭ���ݴ\-��_k�J�\j�aM&&�!^X����\=:��!�y�{Us�w�N�6�Y�ک#�p�v��uTK���LZkpGQL�OtݕW���g'��'�%a������}r���S�V̚=��^�ƪ�*�8������큙��-RnN3l��D���8�wno��}��
��
�+�

�+��* � ����
�+�DTA_�AQ�W��TA_�AQ�ED��* ��TA\AQ(* ��Q�W�����ED�DTA_�AQ|AQ��d�Mem��4�~�Ae�����v@��������/z>�f��I)��E$����RV�)�l�RDI����j�҅iKX+m�q�MaV0���ZG�uk�fմ��U4��4��c�-�-�[[4�6V�6�(�6�w|op�U��يB�MF�YU�֦��44�d��,M�
���[[,��[V����l�Jٕ����S�U��x ��V�C�]\����Ut�:�eZҭF�H�;��kmZ�wk�UJ�\.��m��jæ;]�c�+G�����[e�MI؍Z�  �tQT/;�L�\�j���GZ�u��֊�[��k�֘%6c�;S��f�U��6�j�
��V� 9^��EkI�+Z��p � P ��g��  �@({��  {�x�@( o^�� ����ڵ�j��s�Kt�:;u�cj�T��]�Z�i�n[36��M��f�K[� ��-�l^��*�u����4c]6��������m[a�k��n��\�ͷj۴��ֲcB��ͱʹu�S�Fm�  �^u�j�hR�wU.�B�̪�f�*�5mV���tnV�(F�۫�ӡ�9���3��ѵ��  �� �Y�.]����w ܸt�p7wL(�����e��@�ʶ��6R��mF�� ��
lb <��*�!@�m�M&��5 �q˶��
�� ��խV����X��� wj��c���U��;� gc�Qhv�F�k S;� ��P�խ��Z������z	ɺ�r�Gr�R��� 칎�;�
�]s�`�UA+M�mU#��< ��-� i�2u�Q�θ�b�np��ۦ9��	^j�c#e4էϪz@  �)(�� 0L���"��SM �     �{&M%U@       j��	R�0 40�C (�	�&�2b��O)�4�jxLPI��2�P�F�i茘 M4�9���r�8��˧c�YeF�cu�I�k�[�¸��Nޒ�zיZ�~�I$�!�i���a�dQ��`��@ 7� (�G�TD���/�~��	@�1�$r���
@��UDL`�HH���UDK�o�~�~ֳpN\:x�ۈ(�� �ؔ���ᮁ�&����W���)D_���/��-��Z�o _��T#�h���תS��7w�N��H`����Vʇ�N�uz�R4������h詳e�0FV�u�1V��Vp�S腴�+p�ad�>��ǶP� �O �.7�HC�Jo2X��z.��§�Y��a���q��jT�X��6k$��-��2��GJ��T��2c��Q�z��1L�X��%n�Q�ܷ���j�p���ٵ��j��������A𲙻mp�ͤ����3Z���z�u��f��>�Pa<"��L�]ݭ�f�Q�'
i2Ӭ��/N�e���y�`�#icbҚf$�r�8��ɷ%Q¶<5�245��,�en�Tۼq�G{�h�����ӍQ���JD�V��6��E�)�r�P$� I�)Q.[�-��3d�ٖrkQ(/��n=�R��.Z��ЇM�%%j�k2�`6w0�O+57)d�7TT���@ɺjl3*�-��*��n��t��oΈ���!3W�95e]H�������1�³B�=����a��
�a�,(�!�n�0�M��J#PGD�)�k����n�_�S�ȁ���n���aԏw!��2���d]1���|q7�gv�X2�nԼr�ƶF7V�v���/Y�X�,9d04c Չ�ݐInއ
�
I����#Y�n�℈^e��eY
�5�R��!�Ct�Ң!�%itŸt�ݪ;�R���vIm<�K)�`�4�9���w",���	�RƠjH�� �)�Z�#���Ɲ��#����[��MiHW�z�U��5��y�+���;Y�h��r�����*A�2j9R��n�)�T�ͣ�>�t7&$����:E1�Z�xvل��P֡�t�(�v�V\�V�Uqe�35]h���A53G�����@J���l*�=��6�f��KY� զ����V��	Bʳ�d�n�����v���$�ۆ���Q�vv�oma�Q
��±�W�h�.���[#�,��4ӄ���L�]Ea-nF�������u�����*����#y��MB�hn���9B��.5��ӻ�E	O.nQ�"�8�w�wlCJ�ҥZo4��R�/DB�f+����+	�[�M"�6���9��,�m���^F.�8`�BnC)W1�MX���kic��ѵ5�G0���+Vm����Z�2����n��)4f���&�˫ךY2��!UW�éT��ȭL"}�I	�CIӦ\�6��7aR�Jvl�m��?9Z��I3{Y3E�i�`�nR����)҉:l�r�؛�q��B����/r�cX۸��휚!����x��!�E�;zI	h'r�[I]�"�ʽ)���VkM�%��-.��!̘%�ͻ&��ևF�j�-1�v{la!��ne2P�ڙr��ҒL��h���E�U�f]L�^�XXr���X�(��pCO/(+E'3+[�*C�@�uik�v�%��p ��6(�*�<��k��зZ�+^�\����m��6��20��z�m��#�b�yPZR�9eX���>�w0NR�ԊKE�)}�i;�o! �������1d�=�$�h��uè�\��R�����d�hRƥ��h�Zܧ�6�A�^�JU�֪��ݐ$���(fi܆�:B[UM�b�28uˆ5����ۛ�br��lWJkKU
�7���D+sL���:�S)��C`�K�8tUd&�b7��D0�=��7v3b�q��Ż���*��Z�̇D�oE�Sj��]�H��tdu{�K�)�d������}��(Ce�v��4j��!��q�C��Ejv�����P�:�/���bϐ��{�-������Gs(X����9{�l�ShPr�%b�<�	P:�!Q��o2ܨ�Ge+/���(-�*���
�UL
�($t�50$���ճ��i�ڔôVJd˭�JcĲPn�V�5�Fe�Z���Kkh��٤��YFf��[m�*� �S�`��i�5*�\��/��|V��]��!�V��2��`�����]�D��έΡeB֐ ��A����2��
]���g;d�ȵOxe�,�{�Lm�ä���=�f`M��AC�p2u�zb�g�R�B�EU�0���$V9uz>&լ�lf�j��ZJ��m.�$��Ȱ�feN����t��bYXs!��R�si}�spIZ�����n���˭˭*IYvp�g--ݯ�%`DQMn�8�n�ǎ�5�"�l�R��)�[Xd���d�ʎ��� �X��R-��h+	���b[��U�P6�����A�w �qj"J�Ö��BʫāݗZ�p�<��j^�a�y�n��S4����f@�
&:�
�hc��YM�y5�����O(մ��L3.Q�n��2��æٿ�E������7���^���݄�j�rf�ut�q͊^mޚ��P���Y�,c(�YM��r��Ř]��eP�e<�P�`�=�A�^����b�D�E�]X�،��VV�����Wx5e(q܁���&�-Q�J��ͽ؝+A=s�5�ً�rV�#{N�Ueψ�{[���^�uX���Z��ܚ��zk�����'ۏE��b'��Q�'�i�b�m���b@«���e<�� n�YŶ��n�Ȗ��,�j��Tj�Z��nmM�$#V	0[)�y(���, l]�q�em�>t��xL�%�x,,�����F��4���U�he���E�{���+8�W�[��3��%�z�Z�ܰ�s���<hs�H�	ӷ�"-u����a[$���H�7Os��N�з)<Kc���yR��I���M�Uk9o`X�[�Q����HQ�Z�R`�n:�� �S&�v��t�J�X�l
&�u�m�N�M<5zoD��y�%X�Ø�ik(�6��3C:AÅEUZ�*�M�*hґ�ƃ�fL��h�j��7	�(���ͷ4-SM�C�	r�Ĥ��ت��1�Rhx//e�36B��2R�jJ�wp*�B�:Q���r!JhU�x��Z�Й&��M&so�B*�rQ'��Fp�+3d�֛;m^Cy��$��TjZAn��ٗ���Ѹ��7L�f%e%.�Ò!(j��M���-��3j}������4rۊ��0Q�Iڻ���[��e=-α�.�u��pCyf�\��޳���ڳt��@wβ��o2�V�(^\�m��v��ֈ6\ͤ�a�%K~��6���H����he��١���KL�M4͊ٻ�p�f��ɺ+\Ǳ��Fni���w��>�e�
�ef��"{w�� 2�h*V2���̎��7�D�-E�SX�4�<s���J�����y43^P9�VdYo1@��U��m��GL7V��)�U:�U]3�Y�*R�f�i��b���qMT�k2�Z�60�)�6$^�R��&�T&;�I�55���`PBb�㢁�5I%��%�ϱj%��`�xmme�7-�1�۶N5"��� �h���el����f�Y5dp\
��[r�m�����4M^Mn���8�6�%ؖu��SeֈK�hx������B�@��ԕ��қ������Z��/�xr�DT&]�\�U6�v��#�!Em�&�SÓ�����*+-|u!F�4T���Hb�l�1S�BK�墂)|�-��De�f9�*l�cyA����Y1l/v��蕖�ۓ
pn������٫�YKHں7}H��[���E[���B�kv����De�n��&�͆�me,$���x��@�F����n��)�b���IRβ��U��,G�!{&(,-	H&\²����Ȫŀu�W����V�8�&��iThL(����w��q^�_Jݔm0��E;�d[(3Y�m���/+)����7lK
�$Y����[��U�H�xT��k"��XEn�&!b^��{�h[�)�w�mL:-�u���:���_DQR���p��Q�lb`)٦*h$N��۬���V�@xV�Rk%WA(A��`ଈϖD��&�T�U��W㧵�J#-��Ƶ��x�S��b���;WbC���R�;�aj���]f��:�R�Ց���)�T�p�ٶEi+%��GS1=�e�E�e�L�D5&�ݠ����PGL�V�GXv�@��rꊂ���RܺN;i|����KR�mP�a��؅<�rZ%�W%�V��Sv�,ڸ++e��0эi�K70�z��vpb�l���F�"ZN�uV�JmA�(e�5��/��"�ThmL��<�p�l`�	)7�w&B�C0�7+�B�$�qm�1�9f[�2�J��GZ�f�)F�6��@�YY��w6��L��Z�z��v]tN���X1�Mc�TCT���aі�jcJ��R�kmk�9�D:Fƍ�ǘ������&�`��K;�e���Q>�����
n�/)~���f��������WF|^=0M�^�CU����v�zC�LJЃK�S,!Hf�@EI��i��ګ)8��z�̛yOr�,�<�&��E���S���6EZ�R�*�̺7rn���8o�-�^�D�� v�V��%�e
��Үڼq�[SRfUG!�]�$`���˗7[�I0-kt�z��ܳ!9�^+P��sEm�
�)6h�]Kw�hN�c���Vosw>y�h3��&����h�.�������CPU�yN�S��
�[7]��b�]ؠj�ytv��n9Bd��pZ���w.j���vQUI�	`哢��Eb:%��UO��0T���0-���.��4V�j���E��J�-�֠/�ۦRx`�4��j�*���s���{g\JZu����zOI��+H^A��T� %ԡ���/.5�A���������$�v���ܲ�&`κ�ݴ�T����!,,L����ٵ;H�/Mk&��j�\w'+w�3Qw�EΫއ��,�U�L�ԅ�;;(&�wϮ��L��Q)6#f���(E��{����Cd^Σ	�Y�Z6�愡j��Ԗн���Hv�k���f�O�AK:_"gG�t�cy�(f]��(��Ә�ǀ��1e�L�2�}�;#ŝ�:�{����9V���K����J�ա[�Y��3������ǅ�9.t��\Amo��iۧݧw�]QUϸ#m,XF_#�4�D���U��՘�->��b>������ϞI���jW\9?�6�guq]fœ�'���|���QP��l�BV�=CG���BKʴ��U{�1��ʒ��+�>3����k�N�h]��b�{�"��ݼ\u�ކ�oCpM�0�M5��gb;!Hy-�P.v�|�y2��\j.
��y��]g���1<���Yj��]����0����gWT5�K�\�2)Ճ������EfX�קbI$y�w3���⣬>�z �}�x�-��%#���v���ȵ�e���k�m�s%��y�첩Z��汊�7��-��6�}��;��.�\	&���&��f4%
f��9QU��C��2�7w�m�WjW�3q%�I� ��9��f#��8��d���c��ħ��LSWi# �q�.vu�	�f���i*t�|Z��݊�+<m0�r���N�6��+n�ʮ�7���^��Ќ�ؖl��+LR�J,Z��q�`��h��0�֦t\8�C1oP"R�Ɠ��;�*V�(U����W#�u�z.���^sKso%=I4r��W�P�]�J���C��%dS�h̋[4Fv]`�b巏�T����#�(��^�ʰ�؝���p [��6���~g���"��s.4޸ze����lgn.*�rD(�Lx�U�\M���sx.�ê.J��gw�ndaD��}G���+���;�[ڭ8��*�77����I����#4��b��-ȹd��GVS;a�M��:F�
K�ᷝ��*����9'Q���}0���R��#;�v"W�/o-X����%M�D�^�2�^��$ս��z�
�i.wRMR�U�V��N=4)�.�Ԝf���1���)��[����:j�Σ���6YW4�sl�i�^�INҍq�\�R�|���ǝ�d�k1�ַN*)�ǚ�e��Q@9�e��T�X�ݩ9�!ޙ���첂��"W�ۢ��W�q!E��_UǑ�[Y�Q��M���W6SPSNͽኡ�ܩ�Ϊr�cI��v-�\�	�z�a��2�o���A���-:.���W�U{0J�ټ�l�2�V��f���ְ���%��ER��!!�������f}�z�%��v�{�Ԅ
�A��,��$�-��rޡ}��\�U���������ۼTl%9�x�]�2"-B��]�XC�~N��3�9���n�����,AK�Hņ?�\J[B��W��]ݍog]i]QD6͹twd���; �x���|��3z�eJ���ֲ��繟4�֭1$���0�R�f4z��jr7�pwk��yXKyS^_N`�,��U��^�M�SOoۮ���x��2	���(l	�%��;]:;S����Z�2����u�U�rM*ɅlԻA�uԓm��OzoepX�	�t�.���VZ6�إ����A������`�t��J�kۙz��_�� O&N��Q8�׹�t����/ޒC�)6n��Z���Y��{�8�b8�8�ф�;KF"ºZQ��(�Վ��&��3/�p�/�	�/f�8���E�d�ݪĐ���b�wScb	���)Ε�\ je���Uβ����C��J4a۳(e�Ic��~g%chM�;*$1���΄�WRPc;L�ףjce4�q��ZBKi�-]�	�>���Ӎ]6t��L�ݮ��#�%�����gV�{˖ۋ��|�w�I2�o.��JTf֋� ���&��[+�Q�yʆ�����&8�x�E����£L�)Uћw{�f��x��԰� g�eI�B�D�۸rQ�'22�Vs��V�^k
��"fU8������N�H����P����­�Y[ysY�.��9'�r�W�6PЋGp������*�KX��!s(�;9v��]��;�h�ӣ��c%aܮQAڸ�؊�V�*�;ЃU��d;ԃd��Қ|YO:�lښg^�@6��涋��H.��opu���c��{[8�UyZk��0���%�bR^�ͽ�h��%�f��h���ݨ�5�HLvevc&�7W��@\�����i�vّq�%:��)`��d����s��;�n�AX(���z�t�'��y/��OJ���Y���ep1勾��l�.�����qVə�����xP�mBZkP�:�ɏc�o��R�s������I��.]۱qҘ�i�� J��w)�Ŋ�̗*aX��i�.}���ê4$]�cL���������z;V��;�&�<�}� �[�8�}-,�X��Gl9����y�mR�&��u�
�w�$���sdӤ:c8u����_q����]}� ���O:��
��Gb�;�G*�TC�.�b�A�txl��=W��fь�畵k���iU��T�R�� lcg�|)���hg��v(D���o0�tNs��L��RVwa�R��̹���o�NF���rn��BQ�8�=���፵�	1>D���Ҷm�o^���Xn\9EJ��=�&��45%/Z�pN���w��Sg@u��i�2Z�ڴ:`z�b���ިwd�yo�g�é��E�����b%ze�V�6	�����y"���X�b�4����\y6s{�"�[y�	��'���mtkP	���xAod��3�י��z��<�����$�"Ɠ�"�%^A��{Ī��A>Aٗ����-G�[�E`�`�ʜ{ ��Ë�i(ܳ�����C���.�����j(��ò,�Wt�7h㛱�3|����,]��H�-衙A��:�{]z�����bEC��J�ڢ
��\)����l��{s�X�$���éMΕ�n	X��*��Joi��PE;�nhM!cM��w��%h2s�.��\��ڸp�v�����z�M�L�r*(f-#Uo��ѵ&^"��`��<�ݦ�u_*���3���*�*���G�U�kOnT�������)5y�-��s4Vr%��K�
ͽT�Ʉ��oVEI�?3{���l��o�����x�?T�U-1��dݜ�x��F�qz恎jE�э;�ȼ�:��@�wm���3�B�&B_Qx�#����ٱ�2�����sX6znb�&������:\��tɺǔZh�
���K��c.�ڢ�rYE��r���J={��;��{��2�I�s��2�D��T�G'�sӾ#�)�V�������`n�Nf����9��e��0�ˮ�Q��)J��Q�WǩLh,A]�����ZRn��-\�qm����[;����r�j��)}��Z#[�..J���\��E5�ۤ���5˗s!!�Ԭd됪{\�3%Mva��e�y@ژ��#l#�������|�p՛���&[)j�8sE�������+�u�V�O�F�)֋G�����[��&`��Н�1r���L��d�<V�6��A�������ͣ�zN*�`���\�]�BQ�ssf��ٝ��N�t 騤�T�',V��\����1�╴�y�Θ�	C����ɲS�u,JR���bx��|a6u6=�ep糋 �*I
u��搘Qh��A��\�Ҿ(���n _^�W]����b�1g�@Jb��V�O1n%0��^�z��(a��p��24��8GQдu�kW֖�ȴ_#�%=�͕�[�\X�Q����uɫ3���>Ha��޽��U��4ޜA�ᮬZ�V��b9j��v�ۻ<إ�:�ٙC�R�C��$ӊ1��ꥮ�B��PS��+�i�Hq��e� ��vb�c8u9[v�F��R���Ji�z*e�t瑼U]�yX�[1u�O�,�r*<oN�+~gB;��+8�ᴎ�׹&qG/�� �F��+�!��:湆�r�3;�)��%�|B�~4d�ұ�0�cw`�V#;�5�H��iE�:��Av,[�&ݗʤ���d������.���q�ә6(��IS�n��ɓh7ٷp$���|Zҫ���6�mc����<�d*�M��*;��� 1�EE�)j��r�WYpѨqִ{�V�i�m#x90�^J:��R�]gi����Xm-r����T����.\�V^�'-����]tr�u�!��QY�]"��ŉe6������V���Ws��1/��QPqf�q��$�y�W�=5�T����]nP�j
|[��/;ge��J�s4X�M8��b�3�<�z)i[D}R�]Cr���F��+'1�+prm+�����\
��rN�]%�r�v�Dʄ��opB��le+��\�Jf�������nnv�=onKV�&�w"��nU�9�R�h���9:F�!��#�I7�NI�P����<����c�#1_׀PUwQn����U� ���'v���լ�{�_^���."���y:m,�j+�����@�M�dx(K˻�J�,�~!��]#ԑL��u1�r�Z���E�5ވ�N��1�CH{��A&�d�φAZ���+�c����j峛���]�]m^T�	ci ~6[::
?Y�N�0�&���k�H��Շ���I�7)��<��Lo����q�!$�8�f޽�%�e1�V��`���2Heup�("����7�'`dUTTD�L7_��iJJ:.���օd���+a�?��t*h�B�Pܬ�֖��[)wW��GhL�5VK�r݌��ů����2������R8��G8;Sr�2�5���d��`u�#�q;��7ʺ|z��l{�*&�6�<�6�2鮆�`hq�L!v���B�/#�����-�F����)B��X'!i!��\�y��ՖX��6�l�	�4���S����$0�3iٳVhrz.�+z�L�dE��nq�zb���=X5K2jWg/^"�l��7$��R�kN�s��{��u�-�S�yM�H���"5��Ӧ\�����eQ��/0�������&j���5�5q"ژ�u�OY�йb��t2��Rt�h pMj�Y+d
����ڝe�v���zI6d�l�����P�bDz�Gsi�3b����d�lpb�or��3U�ѵV�Y�vn�I4��,�8t��Nڸ���ł�y�l�Ys+� ��Y�H�ҷ�+��&���i�Mj�c��Σ���@�d�)�ƈ�[��%��.�H��pn+c��V��RS1^v�'f2���J���YS��,�{l�ω��T�j��N�z;��D��U޶I�L�VۺTsk�@,8ڵ�qG�d������,����gXݾ�o쵫����E8.�;�Q�xFT|����t�MPE-Z��Uu�$�΢)C�V��Ԕ�p\�7�d*:����g����ҵV����4,p�SY���.�^���6��V'z~Xe̲.u9�W[VV�P�	{�,9Z�^\�mt�%UM3jh�.;�퓹�����I�ar�B"���f�:U�6N�K��ܽ���8�GKE����;�uˮڃ�Ti	k�Õ4�YYu�v��Y[P��+6n�;�\�ޖX�cd"\�C��s,�Bnɠ��c�P�6 R�E�&��:jaO�q�[�)dn�+-iTn�T��wۻTŇ4Z:�%ZmjE�'����b/�i}|�Zµ����ER�d+߹��oQu�KV�38e�p�`�6�D�Q+��VS᫛�t�u�*�����+�1��!��	�/e��y2�'K7r�,s�Q����;B�L�������]�^�	���M�����v,I/�l�������jj]���������W6�5�ĮӴ�qD���%�&�G:�룬���M�2��1z�Z�KbU{]�5=��
X��fcsP�
r�
bbXS%���pI�ҋ̤��]1��:�c��[�$X�e޺��=ݛ9Xl!�휡 �.!�&�o��ۚ�$�5iνke$sU���B���3�:�9W��Ƥiow�4���u��<[,��n���Q
sE�z\Q���0��zFp�yϡ�\УL1m�kbJ�+Ek
S�W��`7���cj�oI���yљx�G4Vb5�k�2씐tX���{/E����d3j���#�\X�׼HU�����FM��V��%ּo�Ѧ�P��"�y�dd1�;�4��r�һz�3�Y5��XǮR�[���i]�	>��oz ���+/��g+R�����gDWZ�ʬ���^n1:}E,p��,�%oڗRzz���H����^����C
9�����ɡ���؍y��DV�*�yb��ì>�x�.�����u��Z��ܽ����a�!�:�=�mUwn�K�
*v9xY��>�)�(�c�,5d�}tn}�Nف<��.u���c�5s�K�Ոi'+��iK�u�;hI��gWl�pWs�+_mvf /�5�1w�/�:R6�{�^U�30���Cʇ��X�{�����}��t��h�)��mj�k��,m�7�2�2�qe�dձ�e�ٟV3��[U�K�T�oWn�o]�Mz��4Q��ba^˳˯M[Y�����V*�4�ʋ�H>mʊm3M��|}��|�,�nc���f�<KO �gQp��W�
&X�+Q���Sqo0sJ�1B٤��K�u��Ȯ�e���xr���!+^3&��5ݯ,��{xq�����XeO��{�[��˩�}6�҆�/8�1`�<=�S��d&�ΐ��vJu�%����2��ccJ�ۙ۩���<7����`�F�7yg���ߋ���,�/���N'���]=�H�U�2`[{2�6�2l��$[J��һ#9+��c[y�up;]Vf�/���s_E��뚱nI)�\F����[#��	kp,�,���r،wv*1d�꺰.��`)8c%]Dy�$\+vn�mt���ܙ��yw3���uwl���6��='�2^S�swK��67�jg]�9�Yy���Kc̛�'m����t���zI�+�}s�o_'��Nl�}glՎ`�O��pڹ*�w\�5b����\����<��R�W��nn�sH�*v-�ϭ��ȯ�)6��2Ԙ���꺼S����wr�����yU���\t�ܣ���>�.�ibء�]
�[$�E\/J��]��w�) {s�a�&[�y!҃�����P�����^����ѽ�18���z�i�m��:�8�\7�o/�.��bJ*�t�Ô�4��;_"[�a��Ϊ���gUT&K�7�r�Y��U�A��^�tf�<8ʽ�G�Q���\�4٬��
�lM��Q�59[2���n:]�![*o'FӼ�΃9%��vL"�)o%eKY�Q=�w��1��ٱ@��[F��k��x��K��Е`�9��q�Q�6��D̉�iJ�F����VPa\,q�'\U�p�kee�x"5�6�|��:q#�rrخuq�m����١T7U_f�D���;Y���V��+u�/7T����IXm@��Au-qC�-GO�(���[kBz��!
��Me�Q��u�].rv�AG4qy�y�v�7�޳������,R2�}��q���d�ZcW�D�y+/�n'W���;��m7c/F"���ذ�!�Ēƞ�C�hNM��\��)��q\� �����QO��è\��8�o����{US,���/�XE����D�KL]��$~��0�b��Fմ����Z����q��霏0��㡝@��ʮڒ���6�awP0v��ǑBs�ϡ�'3K̮D `�'�S�"�-a��B	XU���������(Z�kC�{�:N!ÐGR�+[����������TgC.�U��k9L��`G���RΚ'-�%ލcy|-.]�k
,�2��o���ڨ+��d�Gn�0N8uc��e���&Y�4��;����V�^e�뜎�+i�F i'pG��ʅ�.5�\��Ъ]�F.�L�(���@ԭ�������I�!tخ]N��0jУ`�5oj�*DjX�Y���r�$�%��]}�+��q�3F�Q�y+Fr����c�n���xeuGXʬ5����n��l�ܻ}S�؄ݚɬK��$��]-٣1�T'ŏ[�Xǝ.
W@�Y�֏f�B��c3���T��4��Q���Ec8�ˍGFO��kb ����)��l(q�E�f�X;!������1n�®(vd�n���`���kjQ͂�Rk/Y8S0�+\˴�ޭ�t@G��[�\�i����\&�pn���`�H"X�Ȋ+]�R���و��W4�એ_9�:�vo3(��hI�ʵe�}��n�a�ZRv)F�b�$��z3.���'7�]:Ve���5\4I�;sr<*��O���k����x6�e��#p��{�OQ�]T8�Vkn��ϒ2�je��[�[��vɆ���Vi5���+��{ U�Ӎ_mUNw��)�)���&�8O�,��dn����KnsO�.���f��u��W!�w��ڌ�:��yL�/�^�'�qE@b�wuչuN�����Ԓ��]F���i
z�#�Yy3�lȲ�J�T���B��p�)����U�nV�V�׬6^�{�,�w2�G�@��Q�X׷��u�P��V�|Bz3ĝc7�mqb�W[��N��Ҥ��cT�J��Ǌ�Z�F�nC	���W���5S�Q�CB[��3�b+,��8]�H��4y�ӫx̸0��W��Q�������[5��P��F�:�4��t4
ݨ.�)uxw�����Ӳ\"���lvV��v��N)���5�3EA:��>}}���A�#���Ҵ�qs������ɳ0-�{$�|,n�J��2�EK:����uw*+J���0wٺpdحP�G�u���I1��t4���������}�kYQ]�O�\�;|�No��:0&�
�C�v���&���yb]�Ù� l�����@����G��-A�$�;'E,���gRI;����E� RU�_3N��x����tku���0WE}�0�����8�7l�X8��'r����Z�2�Mb�y|Ѧ�3� �	n��P���^VN0İ^:s��{��;�T�-}��\����*PH�s����k���'�SUHM)	j��������F��'�ْ���v���0^�-�+5�g̮}KCcz���̸�Y��֮�B��-3�#W����4���(�l���WPnC���<$�h�j���'s��{E&���H /.ڹ��N-���o"m�c/�\�F�1r(�j�1�{AњoP��*�dst�Y9&�	��N��S.x�g*s{h�{І�bHrt��x��w$��͂�X�k�	LYb��;XU.�����UN��(�MQ.�,��۵��l'N���ڰ�������y�����q���yD��!Xlᩎo\<C��ϯ*��5n�TU���*�,*��ulyʜ�Q��������(U�Dt���u�Oj�c7��;.�\m`�Vڣ�왻2�rfʸ3/��u׺����'k��A��m��;Q�T�/�1Ң*"@�,�H`%Tхj9�O��������w���T��y�U���a��t\ݕ����5v;W'���"T۸^�E��kuخ��)�P��Y�e��[����Ba�;��Q!4�"E}���.����d��eL�g{h�ɚm#��mB
�"����4��[ gU��T����C(��
�_a�z�7�j�y�r�7�%û5����=�K�m=�9�K���¢r�`���\��H��@fA�x�@ۮ3AΏ�-����k{ں�}|�n_
����'
��ub"�rk�d�mcΑ��7�Gr�:�ު�2U`b4w���lԮثӹxkv��k7V�:�|��G:R�������;�$)*R6�a��A�&��og+f����P*�qP*m����_��v4 Є���j\A`�x�(iݤ�ۋQ�� ���n�GF���n�T��(���ܫ����*	N�Q�W�&	g�!.�C�m�˻f�d����'i�XRQ�N�<Rr<��4c��wd�"�b^��V��eLK��AR���0B�eEZ�h��,UJ��kh��m����G-��jT�DclXQQm�FѴ�DU�eedR�+Z�Zőb�e����6XUe�V��
]6��aR��aR�h��Y`�ceK-�(����H,Q@F
	�U�+�-d�b�DX(J�X����*���� �-�Ym�Q"
��ģ�D���DD(*�*�J� �,���H�,U���X�� ��TODD�<|�o�����C�k-vet�엜��P�e�������a��W-׶�Z�/f��U966�4��u��d�ViǨZ�_�4�[��.��p�^��T�F%8��hwJ���>*�ڻ�p����Pc���f��n��ܵ:�h�+m]K�@=�,�������p��,�}1,�m����n��W9�+��˗��?��@�j/�k�Q�cbEI��M��a�@JrQU�2�����~�
t����	�ʕ�/�kn��Emd��IГ��z��AHj��1Eެ7�C9>e.�l�b�e��B�� ����瘑��s�7$`�7��os^L_g��x~���пWA^o��nyA����D����{
��e��pM�t��S���U'g #>QT��2��h����9^��VC��\��*�6�
��sg��7#�j>���E����}�j��5���,� ��9���f�y':�*:,	�����S�Ƙ�z����o3Y�7�*<57�VeG5et��=�*�����=I�|u"Ʒ#R0ւ?�d{�6Qx��ҫj����z+��Y�-AݠV��@��"�����R�)k�ٳ哥��۟�bu�vv7�D�YE�ΎJ����T�Qc'�-���e���`O�Ջd�=�c�h3�&��=�A>��O�
�F�b�V��-WB����1��=���h�m�=ɨ3����� Щ�zeBb���}�2�bx���"��Y��3�,=H��@X�S!9�����J�6��7�����b�Ƶ^���6 :��S�Ӊ�� ���*�4(�[$��d���9R`��>�S����B��!ElLX�׸�lה[Y:+ ש��\#jF)��9�!@p��	LX��Z�k�c��n{��8��|D��DBS���.�G�n�H������6��,f�\Ϫן��w5����mC@�ЅW:�]=I��R8F)f�ɳ���غ�u/k�t�Ƶ.����L���9F�6"��OG%0(�
�Ĭ��$r������-Hx�?c�5x���J��S���'�^DfH	Ĩ�1�2+H�tNȈ�V.R�X�'�6������Q\�13�Ȝ<VqhX^�FA��h����]�CM���W�0W�\��C���,]���(k����'O�11����E&Ш%K*�\�;���#ɚZ�bTё�Ş��u�Eq���XOT\^��+��\���Ŋ��dt�ʧz+�Z:�.l���C��A��F�=� gh�7K�'������Ⓧ�ʉ���Va��r�|L�7�L�:��r�]}�˞9o�ky&��S�n�+�c�H1�(�D�"���ҩꐍ<�aI������zC��V!�oHr�1i�R8V�6��u_3��sҋ�u3�)Zţn)��z���|�h�7�%����4gmfU8���r�t��<���̙\gTD�GW�g&m�v0z�:H�7���gE�pf"B��r0s��K�����ϣOT�4��Br|�r�S��ez8:��e���`q�>XK�)߳�F�"�85�L��w���M���nߢ)zGDd�
�8��>:|h��㔙���{ʟwN�O77���bY�\�0t/��� y1�b9Q��*�r�Eq���ZGt�ʊb����|g�_40�;_D�&1�f�f�PFt�讖#�	���7�.U���j��ǫio�w�!D�OL<�G��XM[s�5@S7:��v�C���j�O^��w��a�ڸ�&k=�cb�~���vm�k�	Ϩ)jN�Ms�.���cGc�X�C�#"�zAΪq�o�^c���<p��.��:�J���ȧ6�s�SU;��1�݈)��[t�>~���b"�3ݥG}t���i��]�QNƘv�	}9c�#+�����j�Qdd�1�Th�ᝓ��Ӻ�jV{[�k�B�=u���*�d]7�nا>�еW�X+x��H�qB�Fߣ���[}p�ʯ�nj&d�#]]Sר�G0B��X�<Xp�hj�~���F�Ɛ�󹊎�Vy6�i�1"����%������L��t=�������������X�T��.�mX���d��W���;T��i����	ne��E����
����O�s��r���{���z�n�_)=����D���b/� �]�t8
z���=���bI,=z�=��^I���s=��f6EL��0&|y�y(r���'�*���a�Diw���x�y�!\�~\��9�g$�Yqe��ه�J��\��^K�x��^�܅2�bT�T
b~���U��Z�R���'(*�\Ô���t�~�||��,�:��T�F���%�����|��jӢ�Q�6`�u����[�*���Q�K׉T�$�U�lݷ������yS$4̭��Em�݄��M���-U��;W}�ʎi�Eetq!��S#6LLV]
�7"�b�B��(u��n�h���'��>��?h~,g�B�]�I�Z~X1Q����8:����w4O�����iP���#�r9^Q>j�c*��k2�[̕�p�>�c&�/�CJդ*��c�џ��>����)w�x�N>\+��Ub����Z�e��p�+P�nь�;*�T�Kx��m�0`WH�.�^�Lm�o>�z��������;aHN��q�yXn���#��i}��c"�ƃ�GfQQ��ZM5ş�"뗒�bq��+��:(7d1<��<��ϭ�PR����������i�y��r���1,5���CK�����)��i?C>7���z+�2a�+�WR�`R+DP�	�����.�Nβ�R��j�C$�VڔL�uG2*�_3���ǁM��/���=�����l�����fk�wTMʷ{�^n���m�m�YYN�����p�au�FWR�Y-�Q/���8���W=S>9Ն|�T#4�͸��9 �0����\�YK��~"�������g=vN)�nT	�)�QZ�����<�p�˒ާ���y��L���E?��o!B��%a̱��:���M��㩈T~<��� 9}��1)��"{���G9ȓ�1ӛ��b�ΈP
����Bbt�!�8��:sU}��M6t����tFt��h*pb!]"��*ЉB;�Ƴ��W���:������L�Ubg��hb�Z����ƌ���d�v	��r���k+z[�e_[R0D�Dx�b�����(k�+Y>2�5Y�خ����ݛ�g�D;��傽t��l��3Jku+e��!�=%1�{=�����X]�R쭵�T���9B�mS�4d�pg�C�ج��c\=�t-+�]�崦�f�!�7HNPp�_n+J[QGShmn{�)�9�ޤ*vy+�sMi]�jvu�]�gY��bo�,�-M��k���efb΅����I�%��tқ|�<�PM	�D#�;);2��Z��DK��k���r06\T[�J^ϭ�S* ���3�����
L_5y�$rg$�)�P��>du�j���~��a�����ԭ��E�:���p	����9I�V1�ZG�k5t[I)�n�5[F9ٽ\�j�@!��W��B���s~rVJ2/تԨ	fKv[���["����;��A��0+v,T�(]8
I�����^�<Dx��^�����&+σ/- q��e�9J�ٹ���v{YUw��d(۔��T ��P�@U��+��-m�:�L>I'�3�j�pl[\���u�����Z��`C�h��߻�oxEkډNI��
ݖ�Ź�G��]LA�����iAqA?z��-+�P�57�h����5m�v��֬�^�.���U�v�����L7�\�k/���U�j�� 0�)9p�����Jq�s��7���x��3Uzݨpa�K6r<T[nG|���D�XNۜ�B x:��@�shO��.�6f�r|ٍـ�s��+��Ǵ27�U���b����"�K�yَ��I����H�~v"1}#"�P{Ig[���Z�O���}f�k�Yvy'��0�`C�`I���r��ص�~���\��9=�"x�'���d1����E)��do� ��Y���b�&�nC~z���b���
+6�
w׬0㰇U�Ŗ�Wd���Ή�DUK�Z�P��{��R�R�}2ax�隅�t�zA����,��nFC��m���T����wA-<R�ϥO��v�d,��͘���Zv��g�xފ?

��QS��tb�T�9ߤ>��q�~��_s~{����u�����ݸ-��/��r��7�T�rT"��ssk���(m������_�д�ev��g),* �4��ͅ���� �5Ye-[�i�\��Y}�g*��T�ǅ��I�N"W��^ۗ9���|��_9S��{�;T�6��d�V�[�ch��n�͇�#dX���H��p8�uIkIA���ō��o+ˮ�v�չ1S�]*QhHTj:C˨���Skf�>�6�1 ��QK��UHnEx*�"Ҡ�T���5�3~�C{w-�D��_�ΰ+��\B��;]LG�C�"e�u�\�+ɽ�����YKS�eH��1^���L@ts�N�.���b�T� ���~"�P����^���X�T��i��t��$n󸥼�#���s	�}�A�͌+TG�}ž3�+���;ٗ��z�^�g��t�̬���pс.h������͐���6.W;�ĥJL�ݑWT��G�Y�5�/�x�����Go�7���y�캎���-�1�6��0�
)�Ǒ�~�UpaF���~�9��<*�5UB�����pHHPj3�����QČ�J٬�$vn򹣵VGY����rΝ%�\ki�����ܤ���Y���A���P�]�V�q�f�.^���Fs�*7��:dO�7\���]u�|��]2̛�{�U9��;(Ƭիl�RՖ.��X���z����[��c�f\5EK�E�����E�'v�'i�<�u�!]U���To-�t蒺*N_RA�ܪ%�;�êL�/U�4B���
�p�Z����I� AF���	5w7,�.����;o���6nҥ�}�ʲ�t����R�F�;]��m]�z�z͓,����ʊ�\�A�Vg@�<(;�����n����J_u)�A�)��F���5-��c[�)���f�u;��,����6����G6C�,��,�j����|N.g\�n�NJ3���s�&XT�D�������nHҁ���읷>e�Ug$s�kV��r-��o
�v6�[�z�]��V7$���5xB�2���d��}���l�i�_'���͠�\쳽�Y|��/��y�R��<�7|A�Ӊlp���e�<�(e�*���p�hқ�0�`ε���P���'h����Ac|/�t����T��m7�l�g[�G���RT$R��d�gH-��-�&�⨘'{:��+5��V��3�� Y��M��^�}���'�8c��1ٵy�OQ��4X}��Mާh-
��;el0Nc{-�]W%��r��hS&�de������ompڭ����+_S�vܽ
��)uX6��b�\����0�Ȁ܋�a����I:�0c��S�d]s���gU� [}#J�O��w�p��wyWR��-5Md�yt�R���]uG�*������Rk!�vU�؎)�c��j�F��p�AI%�$h�����]B{��\mqě����W[=p�[:"����okJ�p�]�H�+pWw���oJ��g����Em�&	\xu�Q�	������S�k�o���*\�a�Tm!�ӻ̙$��<�{7��VS�����~=���QGM��X�-h�b�0D�����+UYҐUQ��Z��DQ"��lm��¢ȱb#D�2�EV
�V���b�6�1T��������V,X(��1@F����(�YEb�0Y-X,DKeV*�aS-m�b+*�r��X����QDFD�R�@D�EDb�S�1Tb5�c�c1T`�f(��,D!mT�EU(�"��DAd3-��ł��A���0V,Q���E����TQT�"�*$EX���w�����\�L��6�HJ���K�YE���;� _�����w�;9%5�H(#�|�-��~�ێ�$!3q���S1ѧ)}���dn��� �"�����,��Q]����w`oEz��ȝɺ��&v}���rLKq�x�ڛ��ߛkE�������\����R��ޑ< D8`�5�;1Fkq~Iu�����
i~��tnM��JF ��$*�B�EL��lk�j�-�Һ�;B�T�b���:��V�Q�թ���ǂ��Y����R��+��h6y�Ǔ�5�vАs�\�s-�@�@Ⱥ�r�Ϥ�Sj5(Q����0ݗ��!����qo!��U���w�y��∌��C��Q���:P*�S�&!)�b�Ԣ^wrwb�9�B5Hj[�B6&䚠�G�VU��׼�[l;O	m\M���^(9�X���ڻPv4?�'b������Z�������Đ���d6�`8�oU���ѳn�,+��(����b��n��B�5:>u����?|���Kj�:1��m�3��rGk�.J�U�t��x���C�&r�̌�s��c�_�o<+�[�!�)��BX�qcBø�u����GM�q����iK���/�ΚD#A�q�B���M_�hR\�2y�[)mTCb:���d>�~�((z�3@v�au�J���4�jv^�'):C=�t����F�.!�k�[x�j�3�Pw ���9c�����UI���H�x6	�:H�{��*�R�ə�vk}{����=:g�񚁃���puKh<�r�(����ᵉ�������"��Ϛ�}eP�gG�V���G�ccY�L�6����C\��܄�*�;�#�,U��Π.X��k��"5+=S.�;Hw��s��S��1�������,�{����φ��~d������Ҿy@Żv&��T��
�����%���}N�}�P�a�~u�S8V4E���n^ڱ�l�YN���]h������M}�z]�y^�61(Uֻg%�խoB�֒0X��.W3Oo�0��U�+R]RD�p��v�b�K�M��'�a4����O������Z9�rK�|�
IlLn����W�**�9b3֨C��X�&�<����&�~2
�{/PQ�{b��rT��t� 4�E�|V�0�_Tvr�g̷Y�o���� Sa��*-N��vlUu1�B�#�<�����+��M�ڱY=�l	�����P�� 9L@�-ͭ��[���g_{�{�Ⱥ�v�W�NZ�4��w꽠�m�{GJء}��4T�ϼU�y��03�6��5q���q����޷̽���m��j�z�k�9#e�#Sނ��)s{Pkm#�;b9HP��y��jE��Z�b2�U�hW��<t�t]�?���'�fX��{t��+>���{|���e�
���o4f5�>[[�����+^(P�j��ػt7c�w,��D�6.�����\E�C��t�'�+w���F������ ������\;L�<�Z�fu�]Wʠx�����⛜JR>gW߁F0�3���Qw��wVA��&�����Y�F�1 ��E1z!�JH�^�ʀW^�W�2��_�ߛ�)��y��]Ĵ���}&-8�A����.69����=?�!�ny���Ҙ}s��ⳇ�ןN�+B����Bdbk�U���)f^�}����*�Q��£}�:���y&�n�ͿH�&�`$7&+Ң%�n�o���4��/b����Q��܋8�ҥ@S�����a��v{���x$i1��`�$�gr\Zu�܂SiPY.Y�'n�e���`tDd0�WUk�DMe�C��U�)K���#�|s�񻇘���!������yę
�P��Q1{t+7"�L@sї�]R[��ͷp"���7 4����QBª�\S�cR��J�8ͥ�T�V��}?���n���x]�N��5ъ|ݮV��]}EG���sBu>���[pQ>wiry�뭊��-�h=��R�'6P�5m/�T��e��Ce_�V�Z�!Q�;��^ܿ�9�k	������C����µD{h?��������ߦ�_z���8��W��t�C�k���؇o��룈Ga�L�� c�E+ۙ*�xz�^�O�e�/�x����6�ҷQW����2�hW�y�"y��x�w���n���b�Jor��x������}g�.��`n���#��i}�y����k�jV�ICҒ*�w,[��%�"�h���qP3�+"��<���,�7�ʯk7YK&����.�_���ht�F��	�E��ccg�Nt�x��o����|o���nЩ�r
�)�J��
�������H�IK��U�'���/���%���s���UxMi�����>Ko�X4�u�r��7���y�)R`#��*��>�T���?F|���դ��.jy owo�׌
��!�&c��]/^�Rb1�!�g>}���(���ֺPx�J�4j�xO�Ά5����r���)$��5�ټqG��w�slI�O��~wi����Q�՘o<]�u�#+�.J�b�b������S:Up�r1r��D����9P.�%�td�˦�e�C�d�Q�
X�
CSa��R$t�I�TW�G���B��N^kMI:e�*�gTE91�kY\t�گ��������yhń����讚�^�yo�x+)<�K��n�[@^{��� +���*S���g���jۑ�&�!�#JsP���t��N��c}l��PS�mnNT�U�ܠ�m�"��Ѱ/��fJ���+�Ԟ��=~�G�a>Q������^���|J��1�S��]f���^/����L_in��	ҁ�Ϻ�����l��>3#�F�;��/�k�çN��!��}~��q�+�gA�\�o
�Lr��bC��
BMx��;3�O�c.*�j��7�P(j�ha��<KM�p��U���.�}�dm|s��Sr^��w�ʦ����M����Y,�1����i-U�^)"������w�;?�VV����<��j�y�mh�gF��D�>�.➳Kw;�W�];�S��h�WX�<���wY�oPw0>_M�e�[�I�q1-�J� 4$(��¼7랯eM)ph(ϝ]��o3KiY��cPg:��<�:t��o���i���T��t�\���]Ȗ^Xޖ:}Նۛ(��t���|��,K���:���f�r��kmR�״����ÿR�u�.;���Ә:�b4�@�FV��t����\C{F.=�]yaܼ�\�C��sK�+o-�Z�~A&>�he95@�p��za�6*���!E'�ʈ��;�sf6v:�&o'c�*��Nۜ5X�K.�+�)�D�~���q@~���<X�Gcp�pY����hxص<�7R�n���c�}��0ޫS�8R�.�>���u��������Y}�Y��?_ń�L������;Շ[b*U2�J�d�7T/22�g���zML�ֳ҅h�%�3+� |1ö��4d��9.L	*�@�
Hȳ�aP̵��u�K�1X��)m�y����݀B��z�k�Ɇ�����.R�M#�+��q��q���Q�f�}�5�c��Ms�����t����9(�����I'V����>��J�Ho)x�x��a�Vo�����`x�yu��R�.��ʠ��r�&�z�9�[c��8m���{Y-Pi����F��}�ű�7���<F�tZx����N�?N��-/8/��\��x���j:D���7&=�����AoV�?|�ş?��u�c���~�KʻK��N�L��Mt uE��kVN��pÑѱ�e�nP�6���`(�7Nf��j6�ۘ�1T�T��o��o/������z�Э�k�<)t�_�	j]�܈K�����c%��`�Z��A�9��{q�fײCR��Й�n��X�7��Nk��n4��ڽr��/��f�Ն��f�r�e��.�WU�t�n_��ME�w~ =���i'���g�4���lc	#ڮ����!������.R�Õ�9z؉�Pd?"t��<��Z�N�`��'�vAN6��t��GK(F�D?9	�X�\y����E��Q1B�,S��whᝦHNM�Z�Ie�chGM$((Nv j��Y��g������o�y��:�w��]����G��Q9��V��_�͌ld^\n[�D���a�߲e�ȘBܠ�"�B�2`NVet�������\S]�|�gT�#膤W������񼎏Tt�N;rj�VĎ�hH�'�����rՐ��2|�x�s�>F��S����r�i(��ʎz�;�f��nyPk�/���0��6��ܭ�5j��e�.Ջ�Pb����Dҍ3�7d1<����6o?*��H������q�5�Uqc�8�"pJklV�$� �/�{Oy��{"�<�[W(g �]�7���v?�<o��ۑ�2b�U_dw.]}�~�����e3h\Uɏ���C���)H�ƇL߈4(H�*eB�4h7��MZ	�{[���7J��¹t�]O��6��A-Қ_��|����}��C.k���\�����V�s\gk�������u;wX��.|
���Q��#gܦ������:�<5��wOO)�Uе^�K>
b�s«b�������\�!��3��Zڸ��wX�j��R1
=I��� )t�^J�n5��ſ,���%Coe�f ���t
�@߄:b���B/��L���za��<���.�撽�d�
(s��4�������g:�d��aXVi�yN����S���iU ��5l�ڐ���
�l�1��$�AgI�}b�@Q@�������z��{Ͻxi;a�1 ��ud�Y�}��:H):����,���wq��T�(���L.�S�M0�+&{f;`VbM] (�`T�@�m�y��1/9�y����p�)
���,uH)7�<I�
,�,��2q�̂�{�u�i�9a���1+6�+4�b,�eN"�{CI���ݜd�aT$u�Z�����}w�j۾�'�\�sS	�>�WZ�.-t�Ye�\oY�qv�xn���W>}V3^���k���Y����&��&����;7��rZ:Ӓjă���P�X/6�&��[��6���5�w8#�r�ܵ�
[��uC{�y�@&��8����~�������%�2���˴���v��:���K^Fn�.ҭ�-sH�9��T<ڬ%�^��:	�ZWMV�9��7R�:n�M�5��ݱ�������UKWwh��Q1���T�N�a~�o�B����1٬�k�|6lmog_@�#A!����U��]R]A�YVF�kI#�����"^�T�H7^+o7��M��Q%�o���7�B�j�v(�:q��q�4��5��Z�3GQ�R/vgT��0�e���]�du�ƌ��܇����WwPb\x�{E�HG}�����R˫�=��nt�:����i�q���h�G�kv���o����;�ܳ�UB2LvD�]����MU.mG�:�8�\�sq�S��\W���TE���y�w����X��6�9�����"weͣ2p�d�B�8��u��z<��,:��&"�[2��k�x�3�VC�7�E
.���gR΀�'}�-d���2�Ʀd�MY�:ʥ�j��td ��{��վ�i7p����Kj��K��b�ϋ�T�v���v,���+���+&�9��Җϴ�\;��uv�#x�C��<!ͳ8���h��5�p������@�mv��������;�F󯫞҂�A�:�S�9u��)�|�_N������4Lz��&0Z�Ի3�=�)���mؔʈ@��_\��1��Z1���9�	_0ka+�Q���fY��R<e^����B��j+{��ng\���c9�R,c=̔Wv���fn֦��&�7uM��y�v���Im'��u��x�t�Ҁ�����Q];����<WՀ-��W��`�]�:���5ے$P�԰��m̽��Rs�����3�������)~��WB"Q�R�5ۆZV�X�"���PQ����U�)mX�Q[JȪ,D�"�Ŋ�����1�(
�EV"i�,kX�QV5�UU��(��Q���j,b���E��$`����Z1X�E
$ѵBҊD1�be��
+c�"9d��� �QF12�,X�����e�X��EEb*�*T��V"[q�-��b%m�\�D+X�D"
b ��RQ��
�Ub��em
�#Q�������������Է�դ!�e�/�]�/�m�ԇ%���S:7�F�[����/��J�a���<=�{Ҕ�����<"=1p& (��?8��t��R�f�HT׶x�O���0�Ն3�J퓩�:�R
x��ތ����:��ά6�T�
Af��w�|u��5u�m���=@QH/<�3�$:�&jÌ1����i ����2T��Lt��T��:��f0�f�<�h��Y*t�	�T��3�1�zx�o���{���>`v��7HVg��Y���iE'��14�l�m����|��*vä��ȡY�Y1&%E�0���4� �TxJ�F_f�W��v�+�}�G�Ǆ�rr���C�,�����=@��:�����Ն�P;��ͤ�����i6Ɏ3�y��H>H�*<O�G��i���L�-$K� �+6�+ɫ&"��*z��LH,��frϙ1��x�AH)����H
)�:��I�d�*x�}�<0���|d�1��$�=d�!���Y癯����|�tR
t��2m� �q�ެ=T+1��m��x (�5:��3��^��Ն�bw}a�����1�2T�P�%t����x��o�:��>�}��1�2u�d-��<aY�sv:�m��IUR
z��E�����!Xm�}M$���4���E��bi�ى8�H?Y*3��w�)�#�c xD|χ@4ιd�8�E�0���r٤�¡�a�
��W�g��1E�'2�|�R�0��!Y��ud������ދX���k>G��1�T���x��P�
A��|�0��1'�TJͫn�E���͔RbAC=��gl����՚H)[>d�
)��=�]�=�Z�z}뿼�����S�
�l*x�}�s�i��+�'i���1�2W��Շ:��S�8��e@�f�e�
�u�������(iE'�T��������������+������`Go��4��"����}�Ny�9c�[L�g��Q
��%RR���k�a���T�W�j�;:+b�pS�`#;��t�Nɠg5Q<���Q�����[�~o���_�$a���Y�$5׸M3�J�ժ(v��v�ީ�d�o cXVi>5aΩ�a�i�ĕU �xmL��k�[�+{��{r�O/[�{�݊bA@�+1�Ɉ
/�1+�����a�dY��`q�8�f�d���(��9�>a����g(�V0��]�+5��轺�s]s_o�NI���5݆�h�����!_��uH,���IӉ<J�AJ�湝0X)/8�a�Xb$���VV(
,�Ntg�{ǭ�ky�s���'���4�|��LaÅ�$L��4�d�
k� T��^Y1;@�Xca�퓰ߘt�Y�%z�y':��SOG�M�eI�z}�fsy����������՜�� �N3�b�NRbq�a��eH9a��XV �����%a�*(t��}a�Vt�Y�N���B��c��e�{��������5� ��mORUTyLN�+m}`^�
�~]��� ���Y�>L@^5 �0������t>�,�6�1�'�V[�{*��w������|�> D���@t�Xu޲�
��w�4�]�.�2zɤ����I�I��7�A�����o){�+6�@\�P"�@p��t_c�5��%v�/����La���@���|;�&�Y5��4�E%Hwi�8ɉ�z�I��l1��T�
|�S���C��w�w|�9~{���=��|��l�$��W]�J�Y������QH.�������tZG�Cya���I�����8� (�P�>a�<aRXm<�#�Ǆ��k�F�ҏ�o��(���i���=I]=���C����A�{�+XW�Qd�T��z�I��J��S(bz�X�ʐ}�+�P�6�$<IY�=LdBL��/y���|������4R��TQ��K��H �u ��U���
m��'��`�Ej�i�u�+��6�f��:�c[f��JQ���z�Y(�ݣǏs���ʅ(}9*�v�#�{{�{���1'E4�~'i:a�~/I �M��,�|�x}a�8�g_P�٤�°�)|�bAg�E�wE��d4�^2k��>d��\�O�+:��׼�~����}���I���9�0��`u���$���H)��0X,��Y��6��{���gI�M��Ă����RVMe��~�������c�7��6�.�� {��HmBI��n�|��jP�x��|��!�z�>a��HT6����Y��Z��������ef�ć30��g�1:��5~�i��T%C�+6�}<���+��٫"�Y�d��]oV��SL铙H/]�l�N2UC��z^o���=���>{�;O�*O�� �`s�L+=LH)��ea�b�&$�^d�AHk�rJśO�bv�Rm
�n�a����QNr���]"�u纼�y�w�|��h�Vs�q����|�P;���O�+�̤�y�M0�7����$T��󤂐Sѓn0X(w�&Z�ot���G�t�}�}�>�'����ꤩ�2��IXm�H<�l>����
�^�`,�%g̕<@��1H)�'~]n��1�uי'i�Af�{���>���7����p�:d�1��Y�P(��h��A���=�j��}a��8�2t2��6�\�z ����,4�l+�Cĕ�a�SI�W���E�S��G���������	�<<��t��X�gl�6�U���Ĩ=�ۤ��M}f�m�&0:>��Y�&'W���=E��Y9��\��{u���߼��'�d�Y��	'hVs���:H,:;�CI�(�ߔ�a~��^���$i��L풤���;`T�O�H}i)��@
�'����Y��g��]��=��O%���W�WǱsU��(���(�Y,�GJJh�Y �f��WY�"�v��-���^��GDnoI�+�b�_�N`�tq���a��?j��{�������;H,���.�Ro0��,�(���:�ޡ���3j��)�w�'Sh���<�bA��3��tö^�:d�g;�|ׯ�^�<�sw�t�v�S���S�>����+��Ʋi1 �|d��O���&'�d�\ɤ��!x�mP�<�8�>�� 8�+�8��9�JX���<�;a��Vq��ĕ�3��0:@QB���æ��bA}E�3�!P�W�gL��N�P�z�Si+ݪAOP*yՓ�������Ϸ�}����a�t���*Af0�7��AN�a�4�Xv��d�Y�xϾ�I%B��x_�� (��������1���'sWL<aR�y��_r��}s�|�|���4�*����0*m�^Y��큢��B���:����Mr��H
,�=�l�q��߳>�11��Q��I�b��D@��$����&fU�_"~�Sh��5`bA�ν�i��T�wC=I��S�
��$�:�G�B��59f�;L`u>��Y+�M��y�)�e�G�s��_f��=���,� ����XqP��Ag��΍Xb)8ν��A@�\��a�
�u`bIY�,������4�����Y�Mf��S�S�!(��\�R�q���=��hz��$��:2��8��z�5 �L@�gɌ1�H,�������L8�H,�VL��X�i����
M�~�ٽ��]��~��g��VL@QxwCL4�r��wi����:a����5�Y�J�E�O�bC�d�.�
�L>�ֈ)>T�������}^���k���>�p�4��bT����5���$m�&3����t�Y8ʜE�xT��m��,�a�
���Ăϙ���(��2r�6�R
}������n��r�^�}G�i֟�:f�­�n��Y��:��(Ϣtp�c�Y�׵��j�����Z����by��l�6)��1M��[&>r�a��3!CL\L,���0N�v�����M�-�? g��Cj¾2i1��wf2�W�M�:�a=@�Vf$�;�Շ
����f��g9�4�AJ��Ru=����0�����=k�y�o=��������-8�PP�^a4��������m���@���aY�Ne:�����8ϙ��>aݳjCA�8B��>Lg[�$�AgI׎����~����3�N�P=J���bAy�ud�Y�9�t�Ruw�Y��1z;��L*s�{���awE>I�+
��+�f$��l
�o�>�~�/�o�y8I����k)
ä�ݎ�!�Ğ8����SL��Ö�H=P5�i�9a��l���T�����q�8�y�$�}�5˾�ۯ0�wә����n�̳�La��R+�RiE8�~Y��
���²_��M{g�4���c�1�2W�N��Z�� uތ����<d�6�T�uξrz�VW-`D�Lx���d ��\ݳl:H(m%�0�s�(;�t~�	�F�/P�̕��yj:���_'�J4hR��'a���^�O������5����g��hro|���[Q#��Q~�q׵��ƃ=��|�#�1 PU�k.c��R=�L{��cC��&!�,�!X�َ�Vr cnN����
s	E�B|�� �Q����z|��B
O��c��"��r�iV���]�d�e� G�����cUz�fԳ^���)T;��K�q���{�7/��������!E'ʄ�^�TaQq�n[9F]�ޚw:BW��xz�m�ڄ����n^�����$#��i�l�Ǔ�W.ʞ�3�P�o)����M�#���x�گ �u(�:t����4�CL�����G(Rr`̡m��`���ϻ� ��s�����,�6
�bՓv�;�4��.0�#�h�d��r�ݮ���NX��B�F��=F/l�;��,L��fFz���E��c�.��J���0{�N�2��g��B��]�B�
�L�qJ@�m��+nSBef�AG��c�4��/fA����|�V��a���S���
��݁leh��W��kDa'Mj���5���~��쑱%��+�[Bጛs�O��(���s*�\�HW^�ʝ���:�~��G�6����-C�b�}�X!jȣ6��O�Ics�!�o�a�b�u�Yf�kT��V��b����~*sgyYN۸(�vM�*��vQ�^��-�<�uw��Ʒ���1J�;�P���M�8m�ES� s}͔�gB߽w��C}�HF��Q[��f�(5C,թ�B�p�<���������?`�L����C��^�t�_
~
Vm!N��O����?Kfߔ�**[�q|m?g�h�Ë�����e|������s�6a��Qu��ű��?0��>#��Գ-��h�W��=�ԡ�g�}�X������>/�Q� Fܪ��Ի|�q(�F1G;5��*!�|���0���Pm]�OO�8#Ei�/�ae#��5�.6��A�J6�m����_�L˙����2̧Qv����c��29M��T �><x�^���Y'�~C-�ok7�����Bkcβ�-	����`9�T::b3c%E�w�jz�x��K���ԏF��c�͎!�D��CR<��LR�>���N��!)c�ɇ55���c����Y�,��Z�6����W+�}�S4���EB�n#Hu���ݔD����t� �.�*yECY(�e8Ns/)Y�2��tD������ ޗ�5�;�u��HG�B�!@i�p�� �"X���Z�ф�?/91��@` �2�1B�����k=vE(�awgj���z�K7��cR��nlT|~��Y�&5��!j�p����m�{��O�c�bu�v��2��Lr���
&�h��f\m�����MrX�AXb�&sg��7 ��B��E��^LWZ��q�����~b���k���br�'�ȼxG���̙��(
�S�߂�o¦���=kYߋP�tU��ma�G�:�dB�l�<�U!LH�4�Q�u�#mر�`j�GZ�~�s������V�w��l���l�5!���b� �9�__���q��$t���xru|��c��ˎ0:���)b��/�ő�|�,Շ��neS�9��6�k��b�G��W��G��M�Р�w�'RTβX��n��+W/uU�G�x�*�e�%v։�]���	zIy�K�zc�#z�3&˜w�.�ʬ������
�{���Se&���/��I�>k�s �r�E�c�mua��ES|��Ղga�5}8�8��us�67ڣA�_O���GH�4i��u�w�S����s�>锧�#F�� l�V�9Qw�u�
H���e�B��%)R1M�v��R1bTz$�1] А��&N��ijL�V`0��Xbv��LCS`9��!��CS~n�b�pr��eйJu@�zzES��yz.�d�-$�����j'��J�b3��э#�b�!�l���~iX�|_!&}���\P��*���j�x���bTSu1v8P�ݟDR��T܇Ed�3�P{�/7��=ɘ<�X�Ƿ�N��QXj�ϫ��0�m��L�-M���G���	Ԭ�2
nM��M�p�p��%�{":�I�U���x�)�m�g=7�9{�<mT���Ӕm�.�_�i7�Rç���gY��|����MsO��[�؆��6͔���'2l�vʩ{9������]	�B�@u���%��磌���<S��>�6��(d�9t��қ����MA4'J�׊^�"����]=M�o�GN`���<:f�/�9��}�\��̣����q�8D�8�=DR�᩟����.�n���M��o��#t�������#)�p(��=>qn�2iM��A
5N
��8V�EMd.r,�5�8V�6���<��k��������M�ڼCЏJ�O
ޙ�q�o��d/U���憛4<�Z�MI#!�f�ԝ�0���⤧��D��߮�|(|��L<+k���3I)H�&���z� ���W��s�;
U{����9b2�6k-���ҖP^ja�L�k1
��g��/`�:.�����:�@ܔ�N���4�ԄvC��Č5������"}T�r����ߍ�c߆���{�i�(�n�3�Ň���S��5nٔ�z�cҸ�[�^���P��A�mmWX��Ռ����w}\9�F�}�ѡ��Ʒ+N��m�������Q�@M]5�陹LQjɆm�B�a����BU�WT����m����^:�%ъ�+��u����b�c' �R����U�޵�J4�c��y6x����oT,��:�Δ�.���;t�W�Ū�%#�}�2�,&���FWX;�����+yŎm:&�ɸ�$����Hl+�2�kjQ̓�J�n�<0)Vr<z�Yn˘N��뻪6�3��^�,'g&&q�șc;��t��P��<;	�����5b�I�l��A�JTm���&R��kN�ee�;%Ex���Iﮪ��5w^��i���28�FGt=Q��x{Bq��Oon��3��F4���ӛ�4,;ܐ|������1���m"FtQ���c��}
�f�h�Q��8��g���n�����4w�Q)���8	Z���,yٮ��΢�����K[�B�-M��R�ƶ��](}Zm�_�����~��(�Y��+�p˫Z7�:7K�������/��.s�)WC\`Ȋ8���Y�B'�<+�09J��|�*˂Qgme�D��e3�YI��Di�DS�ݑ֕��]͔����H#s%G�|�r�xU3�ٜ�m7m1k�g2g(�"e��[���A�If��ͺ�{q�J����G"ܩY��\�𩽃v:c��eE�O{6Z�K$ʤ���#�n�s�}�r��Y��J��y�U$/I\C1T�<3����{/�VZ�M���3�y��)k]$-�Fd�Mwa�V;�I�t3o`��������(���|�9
�5��^a%��%�1�H�
ɽ�V���ܱ���JV�Ret
���"{`k� ��>�Qreǁc�W��Q5�i�f��u*�QO����ya.�Y:r�p>c^i����-�N|*�V��f�����~�8����5H��kP��f����h�/$��Q�+�A��R/{�֦�rʾT{�p�@����Q@��U����[b�*�"�AF�6ʨ֨��EQDE���"EU#DjX��ZU-��1��""*�*�DTUIU�"��*��-��
j������1�qR�k �TQJR�)���U�`�ʥB�PTAH�((�*��F(�"�q�D+mQ�"�Ʋʐ�fUR�VXc�*�J��(�TE����Kl�,*,-,RT�lET�j�ҌkV[Q����\�6���҅�U%aZ����V֖գ[j�eA�ڲڡl����m�Ymem��YkIX�Jإ���|��}y{͏u1e)�9�.ݚ�������Ϛ�*�Em!kbX��F�����g���x{�4�i��� �1>lӍ"B�]C&o&�6}J���-<��5)e\p����9w���H���.�I��v��~<c�x�#ǻ�AR�F���-M�"��xJ���D]F[wڋY�����ͷc�u(��C����l]�b�t��~���TϤ)�~X����O�s�%�j�x��5�~�2��R�:����|�2�W��B�0.�r���I��Do�^?��g<��-6��QC��*6�ۉ�N�>ɶ<a˨��y}��P�X*�?)�';��޸&S����N�e���,@��B�#�/���W��o�;ga�D���M��ӛ>�~��d<f�j:EzD���������'�9l�ڳq溶/��{W���M��V;�R��/O�_��|���U~J9�h��w��!�,U��Lh�6��x���w̚����S�SA��%�]���ʑ��4=[N\�F��ⳁE�.c���yJ��D˩��@un==���_}U_W<��&�i��v\�������pe��[�BR�8�P3}�㮬�,b���#d\�]3nt(p��Fř�޻Q֬N�W5�o{5��zC�G���s�q�����1��ڠ��h����ǜ�����(�!�~����9hm��'�@�[y�$c|YMP��0g�+]HG��ሥ!�kx8�dl+�P�%Od^e�ͫۉ��B��#b s\�
2��5�g��|k��"l�T�^�H����_� �7�0[���G��5��aj�W�=W72�ɩ��]���gcڄ���W�Mۿ���`ܫ�h�f�f�WX�
Ox.������R+�3g��D7"��(��4F���RN�+;y>��/�!�1LnJ;��,,y�(5d9�2	p��2n�ێʊU�$M��l��-".O��'��Vz���e!Q�Buѣd���푸
)^.&��.�ý%��j�l���c�u�I�t��E_mp����PD�ff�����6�Mg^NG��ߧ�^A�r����Y+j��zM�;��t��m�g�di�HYl
zǭi��	��g�t�S�6�v���&����(
�.��HT�ϕ�)����nJY�H��"!���"�C�]����H�4�rLP���x{��m(����?<�;��yF��&A
�������+��u����Ώ�	q��N&��J��fQ��H���8�#� �pY��_5˚[�K���3�2��!k�܉���u+3ˌH)�O=��{��^��2&��ꘋ
C�!G��1ç�72ȓ�����-0�`U�tS�Ɉ*\�A0鈰�56�Gw����|�}��S�*����YV�<�ܮ��rb!�@�J�<�)������{j��E���<q���X˾���U�ւ���$���P����K%mN#+Y�t;�㔅+٦Qf�R\�BV��NZ��`�ua��{�������7�+�+��,L��┋5���f�4�y�?�_�sxS_a���ƌ�n�Ԕ�/�Ξr2&�ٵe"֡PF�a�sQaϢ@��54�ܳZ�AQ�����a唟O
�rH�	]`N�$���G�h�31�*�a\����+5�,ј-�3PK�;�~?>�O�>Pb�H�0�=v�ޝ<�{���|EqVe��K���7=4=�[>q-��f�B�L� ��6*j��
D���xU*�4�k7fK����xW[�=�h_a���ρ����ź���h̎ٛ��-l���0�b�L:�e+BZ�C��OUl�Ւ�秒�����ӯ�z�!��������`�'��;�������}b�c���S�������=q��j����������Vθqtu��?m���+3��%��ݮ���N�n��a����ܥV/��[u-*9�aAg ș���N~{��{Ò�e��\|�0���O���Λ 6.W�}w'AԲ�<ҩ�6�>s��aC����n{�;
�_�à�S�#'1d,(W5|�E��>a�d�ȇ4�r�}ȣya\�tb��]^�e�>��os���^ZU�aN�ĞXAH{V�x�T~G�YU�;�ni�eZ���(!>(ҍ��d�Uk�@��Wc��V���ҹ�R�j�� P2���f`uݻ$u��3o�0G@l$�=&�N�U�~�
+fܱ��N}jZ�H�aX��Th+j��KKj`t+wchf[���B�~?;P񘨿��B�<B�ںT(���������ڛVg�I�.wA3*�f�ޏ�¬��-yN��<�xjO����B�iם�^�����BȟS�#�Ascz�xWJ�e핮�]���I]s�ĝM�+~�Mp���Fw�	�۲DH�m�䟫Ϫ��c���7o��^]�n(p��1�d$]���)f���F�V�w������ZRuD�B��f�˚Q�E�6�4�#9t�[s��f1���<�^���t�~��隅�t;h xp�ű��?��WC��ۊ�ӭ���cf��O��O���\f�� �T���;�y��4��1}F,~*lӟ�=��+u�C�����a�����>Ur��Q�q����}G|������r�湢�sI)��!�����1�(L�����<�x�^������J37�{���1�fF)q�J-	�t������u!wQ���v�s���4�⤆+K�~�;P�w1ѱ�=D�ylll�cP!�/�^�i(<c��.c�V*���z���5�c�dl';� �Qh���	�q1B�,U�QR:"2!��(P2��5�k=i�:�IΫ�5jpB1�c6���C}-��ܑlRxz��(�g��w1���'�+��[�`�W��f�eه��5��7E�M�.a9�0)���Rv����~�_}�}�Ox��}C�>�������UJ/&��\8�D\�2��e��z,�<}�����
���q���M���:}t�LtE����t���[��с4�ܮ�ȟ9��R�S(@C%������KLڼ|�]]��-�<�^B�TY��hC(����x(�Ӿ�wG<k{3�F��C5��ъs�ll�+7�n�3�Tu��Ex��H�«"�m[��չe�)Edt7>QV�tg|�Q�ڱcd�=�5�"�A�;q4����%bx��Ɖ����E�ɍ���-}~�Ҕ�b�@B��ﷄ��x ����Ɔ�xn��K�}�v�+b����^�Ey�a[��r
BB�+DT�Nf<p_X��Sї*JE�����Y���l@U.-��/��h_\썁��A��������B+�H<�n�6���*��l]㙬v���f6�d�^�g�ǅI��6�,��6xZ�S�۷zQ�(\�eh��l��f��bv��T��p(F�^�{����_4�u\��T�v�s�2��!ը�)�P��U�t�X��7�ֲR��LFW���U�9R1�����X�R1r��D�麑Q3�ie�������^WE�'nr"�r:9:b-Hjb$���KMfq/cw�ؠ�:\����5WܽV2_��O�
����sI=�"��]��̔~��>�A�� ���L�uK7�Bk*����|)a^_x�����ѓ
���"��ezշ!W3E��NkV�-k0R8'0�w&g/��_ٶѫD��@��(��[�^��|��tO�����%M)��#�"T���ʻ���_)�.�]��c��X�guCϧ�S�1}�k67ԽL�̮FzB.:걣�+.{�k/�`��-�.����<�#F�ƥkrÞF�sͺ5���4�d�W����-н����/���oxܑG�i�O �Ij#�줇r���짲��l�N�N"�Ί��j�+����U_UP4��Rq����S? m+�lT�B�|�R��U3T����7�����{�}��b���7�xT��ƾ�1���
�ߨ\�#"qO8��D���^����E��]�p�n"@�x�-=f�7	�ݾ�i����O��<Pb_Խ�JUjT	��P��1�Gcmo؄��?)�~
���״/�Q���>9�d5^��磖N\"V������&�#V�ӥ�Q���9I�=���<Ǐw��0�;ǘ����!�^茘�Y���(��E�
�91J�3gBΞ;���⨀���|��PhaN�ĞXA�Ǵz�y�epQ�-y�H~�'���J����|wB^̂�)k�;;�8R�֓��VR�ؘ" ,u1�2���]��"t�j�׻r�|r�U�.��X������Ld)�� �k��R��B9b�4.��v�������;}�j_�|Z~uÑ���R;�n�tv�w
ڻ��=(�Z�y�mD�:ҴU]�n��_� ���\�Y{�����X�(lۖ0x�	ϔ5<�QT"S��!�{O�2���Qo.¬�Q���ou8��\�C�{[WA�����v.�?Q��㠬	�9���U^��[v,eQ�6��ޯ+5��6�]fݞE���"�!��$'�.[�sP���[�"�H.wj�v�-����
���m��boӂ�U��|W�n�xe�D(���i�^~Xv/���VB�vs��52��@�1�c'���{n<�MT����dY�v�-<T~^����;T��m}�|_��!S�2j)Ք�V5�#��G�ɏѐ�k�c��c��{�򔪺���Z"7�+�b!��>�'W�F���r:(
{ �}�:/�r��l��4�Yd�c��y�)�Z��H�H�G�9hY�~��˯��y���}����*K�|S�i5�5�0X���nԻm��i.7�����}[q�	�2��b֪t;�ı�o>��@�}�~��i��uv�j���0���ռ/Uu_dD]NwPm��X��ssh=�R��ivTL��{f=�T�;3�1M僥;�̨S��k\��P6;��u� 7-_c�j\x��1f�T�f��*�v9�(�-��p�����:�d�[9֚�!e��+��q�$�E�c+nn�b$H�2ܡ6v� ��Ň,gV���.v+$��G��5�KU���h@��.��1��
6Ú��VNJ��$/+�+G�\A��d8��ob��@t��z�ȩ��̗E����\6K�J_=I��q\�fqV���M_M�.�N���FZ�l���sVh�f�Å �׍i��((��l�w瓖�H�� s2�cU�:�n���.�H�ϗ5h�N��Sv���J�zFE��^�I5�'Q""�Is�YÂ4��DN�e������ڵu�-������e,�%�򆝬��#�f#���a����հ6�F*�G�l㷤�ʬe-��a�;d1T&�r���2s�m���n���k��{�1͔v���T52�m��{ĸ���3u15��ٓ��RA��PM0j�wenp�M��u�kG���l�{L�u1O��|3��40pERk�Γ/F��k��q�r��o���ۀ������魷�F�H�cnc�Y�YǤ�%�Q;&g:姺d���.S��Z;{}�qj�+zk����Q�fx�#f���,U2�>ܵ��Z�ə)t�Q�8��b]����n�6�s.�W
�Jib�b��"b#L�bރ����w��sk/��Y9�zr���u�-T�����+ow$;glA����Ib8�p��r�k{�wP�pUѩN��(*d��3V��7�,��Wdԯ9��_�,#Y��R���O2<{J��y��F�x��7[�۩&19G+����Cj�H�wn�*8�����ϺG�F�+�ƭ��A������ה��y����<~�}�2�QTJ�F�11�����+-�m�%���-���h��Z��V�����AE�Z���kZ��h�J[l�RƑmQ�m��+n7*�F�T��̃����D��U�YU+RV�[j
Q,�A�Z���[mm���4�D�"Xі��aF���Z���֖�b�\�帘c4�Y-R��mn6bJ�*6�X�U�T�j�B�Um��BԢ��[�jUm-h�6�R([hԨ6�5P�kQb��--#mh�e�U�J#Z��Dcl+R-b��AR�l�hƵ�ZU)s.V�[�m��Kne26���eZ��(Z#Km�m�ҍ��[kF��-�KU����Ee�[KmZ��[V�eKeV�j���-*Z[���Lʔh�[Z
�1+�fL�hQ���"5X�K�3,�+�G%�h�2�`�h��%Z�@�-�".���j_>���=z�-�����*kR�s!��*q�oY͆�Zl���>O��.o����jK��ﾬ��d�^�����j܋�N=*Tj���٧>��B��k-�j� fK�ɋ8��9����.�
�1� ����X�wx����t
|��9/ v*�S�E!��X�X�8��U�Z��1������ܱV���s�H�-��ce��'sF7��J�aԾg�����es�}����Q9�#��vyonM��QK1����)͈q��"��@�����*��٨"/r���š�m�&�:���	�j�����8���~���WB��}�Lv��!,�a�����f!�j[���-�������.R��Z����4��ʙ���Pu�G�\F�R�%Zm��QV��)���/�ߐ�l�C[�B��E�3mX�03Y����t,͡T����
��̆h#��5���ڝz����n=ÀӨ8��\��1�.)R�I�]����C�v�h���3cYw�
�S
V���*>k
�����S��ū]_ <Si�ڋ~�D���gDn�Mx|G��H��a~��*�В�^�ڋ���#fY�	�L���6���)}��ic���{��Z;D�g[�dcY�㡹H0+�HHN������}�k4d
��b@ض���6���9�;�
�B3J{�Ӊ�O�S�U#7R)����Z|Z�~a�t����65ۭ_y.�#��t�"x�~����0������;:|�Ϸ�-H�R1L�C]S�8c����D���GQO(9�T�̘yN��ܘ��܎�B]�n��u�̥��;f�}�P�����#�ʓ��滱�����:��ˎ����L`�LS����4,��D䍙��
�(�"��7'ϝV���U��Y�d�ZS�_�/B��2}��-6>�0/�u�Hj����<hO/z^RUi���"��gd헕�6����^�z/����	x`{K��YS1'Ε��yhܬd����r��M��;�K�SF&g��}��_4�4U��!�!B:����G����d]��G�,g�$nM���.B��M�L��X��5j��%y&�G��(J~F����4N��{���W�@̗���J�bT��1x�X�F
������7�a����ب6Mm�	h����m�b���u�m��nK�+֯W���\@�
�ߚgA�48���=�@X���m+���/ݒ��;`H�qNׅA���}db�������쩹Y�n3W&�U�$=�S�C�0v/��ku#�1��z�C�)�P�)�U'4���-�˯eM9pnO@�Y�3�2*	�6!L0eyN�T�I�J2g��#biPQa۱u+d]H*lt�hb��6j�i����,��o��51��}~\~g�O�����U���ٸw��G7H��[Sc2�p��.(�oL�r
d��#9ɹ��^�&�;����79mbZ�q
�V|t��y�����Y�zPn�����1�2�e\�<8^����J����%m�m��,���"}~1�^����t���^�Pt]�3٘[D�M�oM��AЮ w.6�*hc
��'�b��k��Wn�I���/����V+�;!9���hC�ِD�"����w�yy����])QR�j��S7:��@F��N�z{[�6����7�y�r\k��]�V͹c ��CS�Eث���\�ftD#`���b�<�Q���nˏ�x�����`KF
�W��~��%!]-*
�>Pcb�W�)�2����
7����;�5��T�F\�SJC�d)��^HO��9뚅~ɯP�HC��B������[Ð�ٳt�o�;���],��9^��PF9�X����N7�T�C�p�+!v;9���52������0
^5xUr~�/��J���2�H��t���^�$x��?Y�j��W�ҬK"�YR���޾4��u��31@�ZCǹ>��:<K��9J�J��,�ݸ̉;����;��_��}�g�2Q�DT} �j���鱓�W��A�讓��W��Y�^��s]����P�}"~�T���n�~���V�����^�:��7;�ɥ\��1�b!�=`���U��8��m}G|��w��ݗ4Ug��T�	�oH��ŷNe���2L����Å�q����m.�rFG9�HWxn��BW0�/B�2~����ǃ<sz����b�����	H�6��c�lq�D��C|�&��r��e>-m�D��A�P��):�� �0`5���z��k�;�l?
6�P�J&6�fIȱ�瘑�[��}_s��[��e1{��'�`l9�C�B���ek�P}����Q>��a�x�=ۼ��ީ��8~l`aTF��N�Jo�Ui���y����3�6��*9����� ��S;�SVb:��GK�Y�nݟz�\j��8#������I���ɂ
�Ϊ*�]f=���!K΢�;v.^�F�X-��j莱2/7w�@{��M6^��Y�<S�HO��>�c����V��W(��.ޛ��kO6d���Ccd7~2����CJk����@��/�Yc�E_��ϛNL����	�G�/�[7���i�����L�$t����3����5����<�_�n����P�C����X��Sk�(Y�A[�Ȇ,N�-�Y�20ҿrv�#�p�ζ�Pe���(� @����4��d�y�є�����Y��axumh�&X�0�O�U�V�����Ml�h�a�t�#J�n�-0��/m�ؤ��"[W���N��X�;gm�W��I+E�vH�l�V�H9�,׬���R��lm`�܄���E�
��ݸ��#�]��H��N�0z@� �̳d1j��y8��{���5vZM���,��W;"��q %�>㔦�"Mx��ļ���v�Y{�xl�A��%~{�'{ŶcG�>xjC��W�ʡa%a�P�ue��K�y�/JFc�<�Yf��+%�)3�[n���)2z[P}����><a��*�Y�zwE;ְ>���=�`��/~R�GH�s��?>簆�/�rr�`�������i�>�S�����q��(jf�Z�eMA�n�u��$��p��}���<|)9'�ooNZ��8��'��숝���۝�{Yʟ�9٣�-*9��c%B��m�gR����^�f�Nԝ��ɮ-����Eu&wcW���E`��Mmg�WOz�ܝyƔ��ogj�Jd�2���Fy��{��)=~��;[���OJz��(�TM���l{���&�cL�ʻH��'�Պ�ާ��˱̘;|wk3罅<h�`���d��Ƃ���tãHemQ��ow'����q��f���qȘz25���h�Ҟߧ���R��ӧ�+�wM�:Ȃm�6t�<Y���6(/pι�f�8*�-��K����qً���򺬶.� �� )fi�#(����RI��׮�R	�	(*Ⱦ�
Ge��f�D�mBյ���u�c�*��,�̓������i��\���y�H-�@�1U�H�W�KM��l�}w��U{N��rsI�>
�֣8��:롄�e��7k2^n�+mWX��FU�<%��R�K��ŀ�B+�ۦ��sY}{W���d���/
'�A�7�u���i�ʷ��܃l�6���ZV�Y���4�\8����}z�u����%�R��x�yN�o�����Mru�ɚt��`;J�*ۨ"�F+�7�"�e�k�-�����L��Br7[ʕq�ΏiƉ��>��y`�1����S��(�4���
iN�~SE��5��v���v�C"hv�⹉�fӶ�mX�r�A�}M��꾥�Cޯq��q�ً�u��B-�`4%H<jѯĲ^|���GF��}���I����H^$g��=[�Q"��q�U��^4���Յ;i[n)���=�!wL	a���!�"qa-*��k]����дؔ�D� gi;� v��Y�)*��$1{V魘H�b����u��-��t&R�U�!��d�,�m�do������Ĭx���d�tzV�NޤMF�O��`�p�axő��J�6��Ik��<�E#�u�(:`s�e�u�˺H�n���\m��]�����xS-���G�!���Xis��l&��ܸ�!sv��E�n���bsL]e�mw�K!�0oEۗ��r�f2^v�ے≧e[�W��m�.�*��U�z ������K/����73�L�k2[��ު7�g$���6Zڰ�X�� RX�k�mr�'��\��=BC�����nxe�"��j���f�I�64Ub����k�K7�ɖ,�lbw�ti��}�yZ}6K�k*f^o���:����'��V��흴�nf�Lɾ�ˈ�y�B��n#�f�{L�`i�*��6��;u;��g�wl]�i����kҐ�$����ҵ�ڡ]�|.+�|o�?��6�J�k�R�@�شNZ�+e��q�����(twАrdѮ�[��2��wc�,T5�ʅ�м�^ְ�J�"/��jU!b΃^ �{OtP�E�/Y%�)̆.����&������C�پ���[?$FZھ��K�^��!�ي��C�9)V�ñ-�ɢӕN���é��j�@�fE�)�LE�B���V4o]b�U�:�2���H1"��q�͛��1]��; %�Q�(�����Y 1��vGGԶ��n�6�
SHS�+Z�;Ƚ�J������pT�1�6�f7��qR�EQ���3P�ٛيԢsn��0p��*vT��[˼l��%j�m��]��KȷKu!5w@����u��,�/���8*q��Z�����]8Ef�2��qW�/���������n���<Wئ4����<��6��r�l�|�j�ʫ���F.�1be�E:4�Վ���C��>�f�)�肞�4���f�:3P�B�%:�U����N���+㶦�̬���}L^�z�dH�+�����OHA�Z��I�]vx�!tz���D�2���+���V��;�nK�e�s��{$�Q�k����˕��7���rx�J�$w:�i�=��ޗ�o���
�ɏ6���>�pI�u���5ub�����ѷc��|��t�<�B�b�.Y%�c�5Qa�����6Eo�:EY꼖 ��v��ǩ��W�]��6wH/��:�k��%��r��2��-�H�P�r9�'�-���Q v_gL�t��]�r�-���ZI�Sm쮻V��K�BӋ�=��L��ȵϳt֊x�)�7�6;��6!�ѻ0�a|�V�SUjGC:�J㢍�u�sw}yz�a:�k鰉l;��u�o#o�5d ��(��j�%-ͣ�������RS� �)קڽ���u2�Z�ḙ��$�����t�E"p�D���)ɡQ�%e�˓�{��"�1�-�V�VV�%2�Ej�B��D��[i�����q��q(ʕ��-���8�D�fE�̙2��K�b�
Tƨ�\��؊6����ō)F�2�2�kH��8�(Qkq(��Q���ֶ��Z!ZELA�E�"ah�UA�h�TFڬTTQ��Ȣ#iD1��[U� ��Tc�F�*��,T�,�V�Db2ĵ
�V&2�d��m�ԬT`�UA��ֱ-�H�
ZQDZ�EAF���"*��s3*#KJ��ʅYF�QEEE���e����AU�F�L�#���X��

̡b�EPEPDDE��b�eI�V"�EDU��1PPU���y��E��W����w9g��VO��Fl`9H��LA��Ѣ�
�72���'�2�՗}�1�[t䒃"0!	����d����0Tm�\�޳jJF��⟒ү!�r���Jk�s2.(5-��#��݈u{�1E�^x�{r�����f��F�B"�]X�,r�	�b��7�ܵ�a�	��`��55��ʡa%~}Oc�.2�-w46X|(4��F�r��8�-�x��k:w9��^�>H*�$#H�{��ۊ��#ݲ+�b��盬�'.�t�B�5ĎJ��=\#3:�B��
�"�Y��e_5���`�����H5�؉���N�t�ҟ`��Q|ŵ�/7Z5:�kT�C��Cf����	D��ci��73�*zz�늬X�IAL�2s�&�A���Nq��9���v?<�QOK���R��ea��"� N<������P�,H�Vk�x��+Q�(�_xx@)��b��}hR��79kj�z�4�0��:w��e��/�K���FP$#�s̭�Y�^]f�~Ũ���ݪ	���S$P�J����T��m�����7�EB���z(z�oBC:��A�(��)S�̵e��|��t=��
�fz(w�]��&+hON%��As��[��o��2p�&vv�
c"<����c�O:�\T�W����eֹ�TZ���GlԎ�>�U�(�q�t8�#�w��[��'��ui�(xpɀ�3"��f��ͬG�J�f1����J5�T�ܾ�F�]D/ޠma��Y�V�>[aŷN���, ����Y���¥U+�3�,��c�8$��؈���	���gt�nk�.��G:f��D��F�$o3�DF��nm<������?xұڱ����%��`�B<TB���)�CY�ь"ql:w)���B�G1 �AW�{:r6��"Jf65��⩫��m��yM�c���bʭ��55gX�T�p6;2�R�Wr�u�r�0Ձ�e�y��TR��w�}��O�ұYT-��#2�(��f87�ɖ�ݦ�<J��8�Z�Ln��(U�lc��2�7��p�c5���=g慆(�T�E��i��O��*^���Z�\^���r��Y�Y"�X��v"�ɋ�$=�'H�=G������Xu�Ls��ws9����i�IF�1��Ht��I������t��=p��!J¾Q*5�?\Ojl74q,��A=�5�e�jWU��r���)̰pWs�s�Q��y/+/m�K�V�ݮ=Ă�7���C���K.���<H���+�XdՊ)q_�UWծ��~sYW_���I$A�:w�:Gr��b�<�m������6���W6⟈ι=Bf�˘z.��U�S|RRq�8v�#ֺ�:��ĥ�"75a�׵Y1n֢���UF�k=f���	8a"�%@4�C��s+7x���{R���|XI8�846��d��"s��^�5��'TMe�6��D;�mS;ɌՅ����B�ڪj�-�J�Z���R�����RՄ085��=G��m�l������y's(ѫP��e=.h�G'6�N��ZғJ��{�^aA�9��æU���^��a�̣p]�6�ɣow4䠲���Yϧ�<�m�ƕ��&+P�t�\�r�3��,齋w�/�b�[ۂl��F;\�;t�.l��)��V;����g�-q������{��7�Ko�p�}�mP��e��9�=c�*)Xm:�c���w��!7*	��X}����n������;̥�t�ě\7"8F�E���;��z�B(_>�K7��?9�Λr��N�!BM>��V:����-�e��ri�Y��aHٞ�4L1��|��=�Z�'ft��D�h�lj�����ūV��LJN^	9�GoJ��=����q,f�!q�H|��U6�"���EÍ�ǘ�P�0{.f�M���Wty��<b[�*�e][�5�(R2�����r�T�5��m�!I�  b�݄2��?(%T�8j1b�w�yl�8�6�C���h(�TC8Ya���S_òm�T	ݩP��ǥ1�����ٔp���=���6��ڹ��O܁�RE��M�׎s.Q�T�d� ����t�DG�H����\47<+���j9�yx-���-��99����MY4f=�)N�t��w.i,�����R:�0�bԴ����_2�b�OS��3�Q�J�\��ȩ�g�׽��\_s�*���hɺ�X���I�=yh=%�N�Խ^K[��v�Q�K�L��Dn*��96٢�r�22Mƻ8��"A�3K��:�$^S}��C��p�Q��qS��z,��oZ/�pB��<�Z��L�gH�[.���l1;q&��\�c��[�Q-�4o�o��и�Ԓ8��-�Q��]f^�;�K��[��P��VV��}l�X-��)m"�wSut��ƔwY	o�%6�-�]��>~g,AU=5��Ev��1\8�
��E��W��6�W��p΍q����6p��xK)l�\��.�A� ��@L�莌ڊѺ�$�PXc������]$����B���tx����^�j�K�s<�
�Q�S۬�Ŕ���*��Q4nZka�k���F�SU2��+�I%�u����ꚺy4ګ�{M+j���l���;�^r�tO�ݣ��ݬ����Ȣ�EnT6��|K�v�m��F�\x�TګmW[�6{������囮�@���`��F��Z~c$^��L��֋����]�3}jȡ���X��V�������VO�Mz��:�F���x��-�Qw� �QM���4*f���nӠq��s���Z����_��9�/O���OFoP�k�k�p]ՙo\;fsI��O�pڞ\x楞��m]ڑ��P��Bw#f1��Z�Y�}J���l���Қ�,��+�{ؒ������R�+wj!�eW�j_axr�Vy��Ȍ�w=>�yXz�f�e��iTֺZ��춒2�m��������g/̌6��E�D_6����Z�.�	���MDڵ9�i5��UB�/�˵	8A�����8�a\��422C�R��\W�$��2���Tl���N�ik;E�H� t�s�QYV�W��v�	g�k7Ǯ�����@��(ni��]97b}��.�8��)';�|�cp��%�un�JéIJ�d�2a��o�8m�{]m��.홀�w��#����:���3D��g���g�DMRj�ҭGz�]��͒�ɻZB4�4{�Ep˾�&�Sm��v�Nx�$Խ佤J�l���&z�:��܊s�-O�x蝵ޔ_��E��sI�*�ۍ����}�9�Bgx:s��h�Y����V8��͍�4���(�H^��9F۝����3�-gLPt�5�$�7r�ݰH�c+�7*g�NȤ��fR��ܛ��{���c�պN�P����)=�c�r;k��4<i�'93�D#C9�EDd�e��a�Yʓ�����r������X����YG�'%�����Vy:#��uT�&^?m�2K�,�JՒ�N�=.��zc��JE,��t��E|�Sf���'kA�׷W������n����Ż�2��Rr�ĭ�K�<�7�:T$�]yM$`m��"%-D��m��!�ίNK5^�٫*�腃x����������-��$�=� )f��FV���u��DY-j)n��% �G�*(��r��mެ��Zp%��|�Ƅ���\��S�ufÉ�R93�$�QN��&��uO$G`&(��7����-���D���R����ށ�� ��v1���x���] �veܚJ��Ou�ںHY�6'%�ĚJg�I�nC*�j�;J�eP�>�F^,�s|*M2�Զ���@F���1������>�e��-���Yŕ�9�ە���t�9�ڨB�OpS����I��n���)�좁����&�<�Ġ��qGt�5��Y��gg]�O��jJ���򚄢V�G^�)�x�9�ٝ���
�����p�$�v7G}/�V�);."�`��][K	ËAw���8M�]�G%^ΊQ@�o6�Z���&n"I��3�r}7#�m�R�.�Z��̜m-РK�f����ԍ�.�ǱP�5e.��.9Hڏwav)��zC�ʆS.[�)[4��Ϯ�d�mA{�M��,唨n`�U+^9Lػ��3�����v��r�
ef�ZS���ڑ�kxrys���T�q�R��ӻ.�;F7�.A���
9Y��Z��MV�eg*Y�7�WD��Z�Xv^�[vm,<OJꏒ%�|E҆䛩
�"��M���+$2Bs}���T�Eʾ��N��G���[��+�˃��eY�����*^�iO�r;ΐ�Y.|E̾�af�@����,��g�2�We�}u'"DH)AZ��U�ex�J������ag=k�@�k���V�� ����Ȕ�ǰH݆�TVN#��g��*̶��A����}���h�X-�m�v��W�P��F8�����ݓ�ɳG6�j���W.β�t��9ݬt�-\�f�r�Ma��qiŐ3f�(���5vi�äW���we�Ôm�g!�pnF�B�R/L�Q�y8ozFݮ8��(w-�[<���HWR�3���R
� �F�v�xԨ��.�ՑN�4�;;�����ta�D��w�@o4�1ʺRkrU�9\E�Ư�=��M�\^mŌ�9Ǚ�OJQ\������[��:ٕu��R��<�2`r��LS"
��CnV����(c��+���0�(��-ܫ�'�+�;���]j_to�+wq*]YZ�fV攓�*cc���a62�ލ.�v�婟�'��^��	Z7Pn�-�V4�tӾ0�N��ؽT	�&��(��IGq��$攋q�w�zt��7y�_Q.�W�r�"+EdASTU-�,�E ���\��EPPDX�b�Q`���D���"�Ud�
(�m��X��F*�X�"#2,��EX��EX�dAT����1B�TX��T����1`�b
��U�
*�*��R
��@Ab#QTH�"�UV"*��b���""�*�
*+V(��H1AV"�Tb(�QEEX��U���PchQb(��DE�*�o�
�cA�`�ֵ���PJ؊��*T�cPQX1J�R ���TX(Ȃ(���Eb���e�Ecr�E�(�Qc��^��׾>|����+�s/vi��TxD�c������޻(�.�i)�+t�L��5���~W���]�[9x��C�dC�"��g_e������_XΜ�[�w�Æ�;'�lR�m2Ճ�K�Be�G�]�^�/&K]B�t�3���0�9�RS̓�ɞg��WӋ�}8����P���N�:U�V4�^=��f���[��A��/�7�fl�S����L��V1�]ҝ/�N�bW�f"��LQ!��%ܚ�o1�5����e��%�n�Y��)��s��G�Dz���*�JÞ`�� ���\�U�6�n����Se���y��O,�͒�7n����"끔�W���~�YZ$Ӯ�剰�,#��.��>)�%�Ӗ���R���q۔�R
51�Q�YTR���?_>�R�}��76�v�M���vM&��S�m�7�*]�1����&:z�G
v�z�ݬ��%�ĝ�k�[V^�7:Mx�rv��J�g0lGCV�:Y���t�[�C�ţ�P|��Z�~�u�q/W<�w9	S��b;�Z��y��s��]���I(�Ňu*�η����s�}� jF6!���m��N�n�(=r0�������M�u�MlSOJsn��n��;�6ĹFi��������:�k��Z��j���<�P<,�Yӝ'r^�%�Fۮe�]$R4����(�V �[�6"�o�2�]����j@�*Bs7ta{�c��^�b�^L��	/����Q�e�ں�졼`TBR�R����pw)��c�aʇ�� �9�*�u�DΝr=@
��v�g-H�\�超4�e���R�K�������gV*��0�Sv�����u1�ġۊqGB�����/��s4p�C%��t�C��>�Ee��0p�5O�4�^�֐��F�5^�g�ERhF����e�Kf��0:P�#\rXzOEPᙝ[Q�5v-�����wO�\���\	��X�=�(����%���pյB���B��F�ūbw��=�j[8U��S�o�ڶ�et9YV�m����}�b=>�IZQ\_'n0q^�7Br��5s�os�;����)֓��﮶�殬UahӢ���"�f���wz|.����LSX#�]���bNv�e���cH��ʳ�C{D���P�w6�����WX�b6��ĥ�E�)
��{c��t�b����Y�S��ie�>��LҺz�.W������ ���H#��D=�-4y�d�[�g����\L�Q;՜z�6Ұ��=�}t圡�╡V��W[�G^����6��`������{y�Di�D���q���HG�flB�;6U���toC�g���'���l] A��7Ms�hU:XkX�٩$�V_o�<ᰊ*	���]�t��Kj���N��[�G0hB��dp(v����kRF0����ͦ���F�Iɞ�M�8ie�(��[8;d�g$p\xj��³���x��^���I��\�\�@|�Z'+�w_��P:�\�=��{�Q�u�\a]����.I�]���i�E��؎��jr���ٳ�T�sN�em��u�ؾ��ͮ����ٽ* ��w�x�}�)��Eܐ�t�(�`kM޸˞��)g��Sb9�h�"eeP�4��[���[}̔�شմ��.�8�2#-��4ཬ2��Ě9��^��U��Ⱦ��f*f��8�
�A�eC,��Y<���FS=y����`��q���]y��L�rT�!�6��3T�~貼n���;u�,�<��,6��9n���Pgz�pʅ�La��������s
D�/����t�b�F�7�����If3z��kYZ�5�^���~��휂��a��y�x�,'2�%Σ��~[[Kk2@�֯����'-֕��:���Po���.���jPCz�Yx�Nod╻Σ�/�Ze�޷�ˤ�2�0V���дؿR��� ��뚩�.��_�g�7��>]�T�}��b�U%@ޭ�4u���X���YR��ٶ��$��0B�F(oFջ�X�`^��@�5����m������ھ��T��c�a��T�p	���)5V2�pXD�j����d>��"c�ƌ�}%z�d5�+,J�w���y���������2�U�I�Έށu݋�-Ts{�.X��^ϖ��x��Z����Szn�h�"�4�=e�]f�l��.k!/Q�۩o&.��#)�R�'�L���W�G��臅��l�W]���p����Sh���3�sE�Ky�)-m�E�eЋ;��-=��^[.���G���ջc��γ*2a�֕�<����t��wv("������[{�wJ\���*vi�/s������gn$��v�Q0�^�H]u�y��C^�z�_��'��H]��I"P2��ճO�	ie�����h5�;-%��m��4�ڪ1N񤕫b^�TA����k����s�5���Q��5�����������F���ȅ���$�`C�8v_@EDٮ
�$���\�q�q���9�
	�i�~��b\ꉬ������d��l�Ԃ�/�I���ڋX���'��q��q�1����{��`��|0�^�SL8eGԖ>qM9e�ȥy|��<�;)��WM��P%���g3X����G�b�6�`u�"��+2�s�%�v�N��,��p�v��S�<��d)(��9 ;�����$e-§��*"�(��M5;�_���=��\���,���/��Rf�O�xj�I�~5��vNy�:\1M�ҭk�������f[r:�W�8M�J�j2��\��B�S�ޝ��C�|ubd��ʎ�
����Tܼ��y3%��ct�כ�ֆz8 f�]1�*�(�ש&O!�r�3r_-�4�H���b�7R���|^�bDO/��u�JC9���J�o�#�8�:��.Ǻ'��AΡ%T��N��%	�S���[�,�w��4��'%��
]�vU�yֱ�UH��D`Z;�>��9�ْ���o݆^e�f�Gz/���A�zĭZ̖84�,�+���*�T%�q������i�,��7���ǋ����{�++;)l�f�
ZM���d��>g3ye��{�Py�|���g!�^FQQDF�wV��q�KSb�6�z%��`Ѕ$#A�z̳��Y]CY��y�`ǃ��T��F)�p���ӟT�KB=���5��(ml;���Υ�L�6��Fׄ���:��Ƭ��j�T���>t.�f��\=$�<28�Q�(NҺʫu���뵾�J4hso5���O"�i�@_o��� }�&����*�Yo{����^|b���c"-&��͎,L�r{�"���&���g�����涳n[����(e��/��$���ֲ[4)�Q�*Yu ړ�W:��8�F�ǔ`�@�3�ђ,H��sr��Y0v7V�H$��$��}��l�JD�{�\RB�'	�(L��M�Wʆ����y�x�jVt��aX|h[�Wuz�c�1�ϳ'96�i��Ux�'�^',Aq�+z�[���l�M*�r���C�kWᒚP�ÆuN���tf!T��TX�4�P÷t�R�/m6,R�	OY$�����y�>���>���&�:O�e�R�K���Ǯj��9s{����x96V�y�P��+��Rv�$��릍��s��+*[h��&j5(���U�y�Yd5�Q=ڢn��B�*Ǽj#9=���ɭ�yo��#�If��=�#s�Cߵ���f}��ڪj볫��5�K �n�"�b S7��8��<n��*d�Y���ё�q�R�mdGѳ��tƗfm���ӏ{�s�Ҋi��^s|��vVoQp�A2^�֛&a�y1x�o.��/�n��c�&*niJ��S�H(rsYs;t����s��T�gf�گ����6ʔu:�꨺�"���_]�0�Ok9�',ZU4�N����Ӱ�S5-�Ϯ�1���-=S:�3�j����8��Y[��[�)�ۥVu�Ok^N��7&��֑��.<�lV��0kVpݣ�co��wT�qb����US��d�u�cJ1�=,�������[X�U&Z0�<-��
�6 ׉�k\+l�Q���j|K�Q���6{Z�r���e���&�3����L��J�l��	9�UO���ֶl�"�լv�����pV�n_7I;S)i.d���
<*ػ؜1���-�p�n��c!���w�Mԅj7�Z���n{������|��mh��7�Ѥ1FV2��9K]&+�o|���)�m.�oD�4����%�U�n|T������+��Vkqø��.4cʴ6��e룢�ܸjt{z4�g4ɓ�U6�09�X1&Em�ǩ�����-]�[F�n[����\t6M�:E͊q貕c�M0Lz!��&$��1��r��u1�syh��w�5άj>�%p\��VU�wiι�k�-QXZ�h�YEtΩd^�*��d{�,���]����<��G3�q�Zյ��)�&�	X��M펫�I>�IGn)��F;7Ը*��ʻ���1;�ͤ.��z���sQ��޵�E.�M3�W�x�야0$��m$��1�T�\]v)3V�ש�@�6	��t��:ޅ|w�1��P���0ۻ�:8ù�O�y�)I����K�{���T1Q@+���놅�V�J�/P��|or���Ək�.�)�EΙ��3�e��쓎�1�k?
��E�٩0��jgw)����i4���gu� ��N9���=���ƹ��|�َAF*�h(��"�QTX�-J&[Fe�b�P�V(,F(�TIZ"$EQ�YlV�µ*�R(�����X�X�"*�"����bbUV
+���cQb�,Q`�����(����DUDE�"�"Ա�DQ�**��,����H�����"
**�X��1L�"VUED�Tm���AT����"��UH�F
��UDE����PH�ʌU�S),b�aTDJR�VV�F1T����Tb*�E����+F1�Z���1(��R�m&dD@��fg���N0�ΐ�T�����9�֕�q�@bX��F��tU�.�����k\�䤚�@g���Cnt����Z�-�rxt�&Z��֯�~�C�Ţ��Pa�"��<3[.�u$�U<"���V������=v�jݢ9�(��j4�������R5�0���5�k�!�	�0<�9���ܦ��BTv��3$T�=�Y"�WU+%6���t�䯏A�G8^�h�q$у���e'k>Ok䒃R���Q�n��v}���H��Y���JY�֤�i[n-��ʝ�E����O(���t�F�����/�\d��bk��fm d�5�֦�g=e\��;�G�w�$��p&o>H	g��Z%5�νC�e�/2�;��pPHl�E��k�@�uf�޻�;;�iV]�a�F%
�}L-�ݬ�U��Y{�`s�u���:��r&ԗ{,��$p�� �R+���h��9��Z7w�J�&Zӄ/�ˑ�0���Kݷܚ���h�%W��E�OV�����3�$�Ss�4��Sv:P"ƨ��=p������-�Ҝڠs-7��(P�B� Ҧ��9�'C	\Y�!�F[wOӆ�im�=և{S�|��l�҉�2L�c�a��p��ϷΎ�cizZ80�x�s���q�!��oe#(a�����c�娶�T�����tV��Q�t�>՘,��-f7�?M<��}KV�-c�NǙ�~�6Ɨ^�nPT���Ų��ȏ��+�Xr��]kJe.���������;=��~"�8kt���m�X�b-/r�O.�*u�X�;E�A���)̼/ f����m��{���6$��i�U*�<�Z9�vq{]��/j6 �ǲ2��v�L\���!�ԩEY���T���sS�y�diX�J��ƹ`r%x�Ω.�t�J���ȫr���\U�=���d�M*�3�NHf�5�vs_ws�V�Ԓ�ǉ]�*��çV�Hx^@SD�bιZ�����Leu�o�����J
�b�1�]��d��Mti05� M�ܮ�-ߌ��B��16����'u&cq��!։�ΊU6n�Jj�ȥ9ԁ.�3f�Z�N����A�X���=��1C^�&q˦�0�$�b�f�f.�����v�����O&F�����3�6�=SP6�F^[gH4��lQ����R�/rU��f�y3Wv�b\�`���|��¥�M�8杻&d5����o���ľ2�v��Q�s-�����r��jɥ���c��kx�g��1�wwU�=���}�h�ךM����#�9Z^���	�ԗ����zS��eh9Z�jy^+) �僻O#�6��m>,�-�y
Tsq�֤,q�)�ݵv����==������,����Y�ԥ���m�Y��SSY�O0g��遃a��V�Y;�'v*���Z��m1]�%x���)��M&[J�]��K��CW�4�q��FvWi]�^e�KJs3-Ƕiu-.���
K�۩�y;5�SYA0���� p�o+}U-��=]�2,��k-�q�ܦQ��{QoM쿲����J2��%\��K�{��m�ƋvJ�Ck���Չ���w
�v8�:P�蜤�d�J]�1K���`��;ƒ\V�"��p��p6k�U���<%ޡ$>�;��	M���&�Fj���m��ٽ�eb]ݼ�K�$0���T�b髠�K�4x��ݦs�F��7Oh����Q�g�D�ѹ���NJ7�[Mg,�c)��7�n����b]�����OqgI]�XU����^�c/�g*r���2��WS	@�y��%V�#0󭪵�-����F��G
��(�⸾[OW��p����=V�	�ȼ��>jW^o7���U�O$:���&H��S��(�b.��ټ��t�)�X�+�)13j���9�t�0'�џn������,mβ�s V�x�@-�t��uq�^5��`,��.�i�z3B�o�(�{��_�Z�V�`��NW����Ҧ$H��nV���\��k�RVN��|�e}^ghbU���Ra_N�㌤{[K��1�+�S4��jQ��Nl4$�ǥqC6��9 }ed�[��:��[<��-��ѩ\�xSj�RF�֧@�$Y��"u�ԝ�d��Y$���R�yp�&�C�}p�Kí�B��<WN�F���֜Rӆ�r�&������;%W+���uG��(
}\���#�~��dۗ[��Bb��Ps��E��rF65�0�7wM��+-
�ҧ��jr#mgM��Ud;�MD�ٕ��9Ou���Z׭
����s�b���%�I��bݍ�L�{���X��oo��QZU�bL�ּ�� ��Ǯl�ЭѦ��X��.������];c/����\:�c�.Պk�-���O=8��d#j�R�NҜ���l�띊��)���a�T����cG�D�NSX*M�0��V�=�2��j�{:�[��TPX6�섯����Ţy����[\�����5y�*Y�vǸ���Qі�!�i�o&�J��^�4����zEDeV#�
mF�?d� ��BT�U��Θ.�����QS��)�-"B�R]I����e��X���p�ާ����B�K�/�N37�F��{���o�aۜ;-u�v�HIxa�T�%���Z{5�FJ�1R���Y�IT��/R��p�����p�2U�t�G��$��R������}�����f�QF�'��������S���Kk\V�O�<dթw$2��q�7)����.u�(���H�]˒���	���F�n��0hB���[�4�xU6���̓�5�u�$S�m��B�ar���V��Q��Zi�������55tei����bDE���2����d0:sA�JM.�
�2�
Wjۥ�]曏8ܧ�ə5�P�~��ǔ��4_P�6��y�5�ii��G7�B匱�Fo;8�Y�qG+\����x�5�4O>u.�v��"��{�;������)KNs&�&y"��5ժ؊��X�k7]Ŭ-��8�m�^�lp��R3jQ=O�4�d�T��
�I=W̵�g1��ߋ�c�H遃j[�L��B�;���i�z%�>�5h&��ѧb�.�cSV�#�q=:a���1s彣Yu�K�/�c��d���[9��+G'�_EJ��(�H�ke��l��\��� X���-D��Fc�3���'��cR4�+�|pH���x�O6�)e���7~�-n��hbK��~���
ʊ��i4�+r��dATڬ[f�����զŊdڅ��Q���I�01��|-R�}T%�Z!V���Me-:��Y�a�!If�Ua$d��:�p�e]�0Y����Y��Qu�-ǫ�ՙ��W6^��!��H4��R;TM�;@ݡYJ�o"�Tm���4vJuԥ��x�j§ֳ�N�ϣm�1��l����cd��[W�I0��N����-�l�9f�[�-+�.���5��Mv���ڱe���3C�%�E"e�A�]�xJ9�k�%�8�o0��Ԯ��Em݉7f�Vm��ݚ��Y�r<?����nM�77`ٻ)3=ӎ����R%c;���sR^�H�*/'�!*Y��F�Y[T-��-3��B��dFQ�e�̻o:�u�<&�r�Σc'��]@�T�W��$�U�d�N�,��VKhУ�����Y�R;g����`�T�JL(ڤ���k�[��IE��W/�є�;i���Rb�D�"����{�Y�lJu}5+�R4��5���ז�E��-)]����9�F�f7�:u'�i,�&;3u�*�S,4�D4��U^�E�:]^+����hJ4��	!^�$p���R�*:�:���x��c��"�H�Ccj�q^C�{���U]�����������K2�j*yR�T)�n�e���r\�[M���R� uI2P��s���J�H��vf6"rw<<TMV��kf&����n3
��h�T$���ٗ�6�K{����)�zJ[�}��]3	��i�T0�E�Z����OGf��k�,oe*�����p�3�Q�M���%�>9������f2�D��<�mͅ�r�h�}xNR��:M�]���kVвx	f,+hWDSBՐ��[x��;KiE�@>ۗ��F�\�m�D�c�,�SAt:��C+;�]E�2�D���#<7 U�g^E��G
vC�R�6nI�4qc�}|����	Cm��d,�$�����.ū79nV�!�˨@�����_f
�_7q�ќ���66��$��@҃[Kf����Ш�TQ��0ޔk��5���n���f��b�mg;R���xzv�`$�����V��%h:E#�>y�t�����-�v�$�fIB���gaN���*š"��kT+����+w���XJ�N�3BZ�,�c���%Q(�[R,�泐�Fe�ؑ7�.�[t���{iMGv3�n���_;Ř:Y�YE�"��b��9�W�`���$[z��'0]�m�E������	�+4��Ҟ���{���(-=r�s��/K �Mޒ��s�*i%����������|jMYpD����Y5[��F����s��Jh�=�׷I_"s3���i�Jn��`�kI9���\��o�S����B�)fXn�&���x䱯�˝v_h���iU�|��U)ޮ��Ү�d��Z;�x�ӫ����{t������/8��t}�4g�"���ᧆyf>^�wnLE�2�6��n���6�*���{i��;à�Meq�(sjjɤKl�B����>mr��A����^,ވ�ɍ9�vu������{�I�z����֩#t����{��Sw����SN�T�h���u�t��䍘�r:=�%%��$��o*��Sԑ�~��U���*���ڨ��R��H���&��U�
Z
��"���mmik*���i*��҈T�QV�����Zʠ�KZe�5`�ԥF�Z��ZZУRԠ���U
�-Z��m����q1�UJ���KT����IlJʕ��[[j�f*�TX�Q����V%�-
�Q-B�(�2�9J�Dm��QF�m���Աljő޷��ߺ�~�Z�xv���Ok���{%i�;�V����H�Y���y���i��ׅ�o�o.Ij����7�h���`�d"��8���G�6��}C:KW�ҕG)��@�}f���ڲ�<���!ؕ�����w��R��76���$��K��N���=�X'����Zz�I�}���6�~�<21Q��Y0����r����w�%�"Y�C�y��t����E�"n�)�fD��ۊ�<���ʯ[�[���^+v�eE,j�r����Z)X���y�[O�:Fu�{���+�dL+�hJ�ܓP�	Б� �,���(����u,�o�j8���qY�S����y�}���l��ķ�ԷL���gf+�㦰��P��Z��L�_���b�'Dە����SJ`��H���9}4����]�R����[�wz(���7���vn����B�D����0V�f��Uኝ�I8��-�뎎����[Y���I�����ĥ�+�vmcJ�J-�3��C�X�/x�]��J���@<�÷u����^�M��7Ʀ���+�=�.��oϩ�2�9]��R�Ca%��Q�����!3�ą#�M�mҽݙ�gOm�Ē�̒y���h�!�W�0R���wҼV5'�e�\+㭫�2�w���M],�MS&�K�X�kj�)��<��R�)wk�$��/Ni1��9����ã��
�]Z�3AѤUp�\ev����6Z�Y=/����Y��C����q���T������_xp�Ө�y,�N��BTA�iY	Xr�X���P�n&��:��NIq=b[Y�+���D>{2�om��W�}�8���Zյ��w�NMrI6U1��б<�us�Fz�P{��:�G`��*mjN3����;F9�ɟR}��!�􃰮7,T�Jtr�oos��4;`f�S��Sϊ���x�K<�8N>�<��ޱ�������l��I�<�;�p���X��$�"B�p"q�U�e$�)��v�b��k{7F$������M��7��}Sʦd[Y^�>�u���-�x,�Gi��]�����6D��P����b�a�t)d���[{��ڨ��U%A��D��<�/�![p�6��Z3u����:�ep��Y�έ�!j�Wa��j��ǯ���n�km�`ͺ3�۴�p����fB^dr�`�;��F�w�<t�@n(����p�5^�Xe��د1�]�-�ܡ,�X�y5���)*9+>���-�ֆ����Q���g���t�RIf�;2�r����:�RÍ�j�׹7��y�c���P�V�����d�kkJ��FS�~��H�:߭����M�\��E�=y*�ԧ/%���A��VL����hV'�zr��P�\�=�V���
����;}[ʆ�Y�l�%ţ����yf	�Z�#���^�%���M��T���i�5����<�҂�V)55n�um�Rv�)XCc,S�ѕ�|v�*�u�%p,f��?���Z.WzQ�V���0���i������*E����mI�q��G�gs��qT�ݙv�����&��3��̎�B���Iز��щTǰ���݊�.����8᙭m�7)R�������b�P��[�����ۇ�MJ1�\E�'ә��:Kj��w�'��I�8�Ϛ����3vzњٴ�mP�x��b�It儐�$H��7:��e��i1=�nj)*-��UXeߟUK!��e�B�"LE�l��e>�%�3+,��t�h���0B!ڷ� q=�u��n���7m��J�)�(�/#c����ޔ�v�)D��fuͥ�I�6P�B21b#�O���cc޵ZuJu6�,��w'H��<a�r���)!ͭ�g6�����Y0�Y�K�k7v��K^���y*;E.d��=R��FPĎ?J�s��-�����G���Sm�|�<k��ׄ�N�y<�C#��gLzI�B�]�kٷ��YΜk���(n��Q��l\��1�������gҌ�a�~.S�>���k9��?ƅRَ��n�-�Z����XW���^������{�x�V����~�z�W��S�{����Mۥ�gCY�2�7w���}9l^YnOx�Ex�F����j;�٘)}�JL�֬y�X�b����r:�%C��W�\�����wMWf�K�������#75ݞi-J��i�o*mB:�:��ŁHM䚏d��N�yA4�s�E�rxb��vY�l^N)|v��ZЋsn(!��ă¦ٶ�^�l�Jۙ�TNR�Uy�P�/�e��2�h��r��蟽�h8jG�pq­�3�H�_�y9��Ԙz��yK��[��+/�Y���,Z�td�f���ؕopl�Gv9J�3ծ�f����	<=>��+��oV��E���BB�.��&*�#p���y���ؓ��E���R��B����k|���
{2�i�[�������{�yOoJ�ը��!ѡ�Te�묲ޛ�Sev��*���<.X��#7��j��v�Fge����̴.���r�7�T��u�}�x��^T��A2W��L���8��xu�ˍJ�Kׄ��u���ު�~S��ދ�:c�G�¸���,p�޻���4��t����'�g��WJ��<�5CK���݆F�O#��eq�G�&��&�`f^��,�t�3�C^��wr������0G.X��3��K\J�ȕ�.Cy�=�c��z���^u���/c�5�HT1S�o5m���J�ِR�V*e.�D�뜞�j#$WR<ר���IE�ܖ��º
��͆�C	]S!�j�WRAlMrx}I>$�r�&�'^�IS����Л��r7����zN�9i���ʒ[��:b�wSi��5�ç�^� yX�Rj���xڞ@��$�AD#:��34���y��J�.h6��������pA�Ǳj�U�֚�Q8�u[�Y+F�Bȏr���.�H��U��L�Ơ��J]S��Sw�FR�m�ҧb�*�{Ji�C�4��pی[m׮P��3��:���Zj&�����ݹs�4��F�S�m�z���)��Y�,�xZ�Ԫ�[]�(��Q���z%�ՙ�*��X)�j�f��װ5�s\�@�V�ݾ%c)��%t�Z�*8a7v8�����u[�eD�8�aw.ڝ�k;a�CL�]�;enN�4�{c��7�i�t�:�Ko�穹����_��[\N̢�]�B�[Z(��r����]��~��B)�����KK����eN9���G���V�@�k�[���;i}�`�h_D´�-�(屲a�w�(���'�\K#��$������nvؼ�lӿ6��Za�����;�e"y5��k�vz���(Pi ���V�u(���-(,1��|n�a����$O���:A�%T=,�ք���"�I�R�Cb�j�P��n�7*����yy��x�X�RL{F�U�K*�i)�*�KkK�O��Ht�h��Y�ɛ��j���t��XO�:�
�(�7i�U��j�W.����l`�#��0��+r�U�27��f��8�)�L�\5�n�^<��,��S8n�>��Nܳ���-���J��zk�5�7�33�l��������a�Qx{�Z�f<ۗ��a4�˱8h[[4�d�eaM�&��b��7�`2���4�J�;Jg3q�|>�o��P^�3�w|+2�݆8�n=4���ޒ#I�B����f8N펋"bj�\���A0�e	�+Ӧ�d_^t�Q�v�V�;|n��4�{�w�W�:k(QYBJ�3�\&P�z.�YT���Y��;Am��F�g����T<+Ӳf8(Q�)��q��gFԘ�j4�"B�BKuۗ5r�ӳȲ��:h:p��ٻ�+�B�J���N�̹��~U���c)M\rR6��r�5�{�J�;;B� �<T5�}��- )��mL�q����p���j1�pGe�+~4O^7�{T��;ڈ!V�Ŷ��2J�B��]�R�H���H�\!><%�W�n����:lr���#�d@s��Y�C�F?�ܰ�QA�v��H�3)}���gtO�ޫs���3�]�ՓU���U��(��EYl�X�Db�V��M�
��@�jUk̾�����&�܀q����#4tzr�\�/e]	��dF��[��jXꔊ��^�vl趻��s�k'j1w}��n��9�ͳ���d�:��5g]�-8g�7�%�l���Q�om\���R����tq�T�G��V\��ӎ��0��E�XB�-f]��i�W����Cc�9}ۤ$��A�ߣ՗]�T�=zѺr񊶚�������ˈ?B͈�����K췫s�10s�JO8���Sy��g/��Nq����
�#S9.��;sM�f�[;������˦�r3g%B�����9\�0m���(e����J��y"�ϖ��鞋j�Vw`������Ɔ[�S����ƀ.I�.���puB�������������gIWҷ{�+�����,*�	��:*��� ]��b�g:��(.h�]���Cv�j��7J5���A�W��k����@!�ٍ�{k�6�Mw�\�k���)e]vJF���p<2_V�t�z��v$�R����ZY+�Ri��� ��)�������5���i��DD�I�Z&���c��t/��3��`ۇR�:�N���Iͦ�Z�<2��se4�2�9۵��6M:��L[ԌnL�p�%�b(���M�����˸#h*츈����$��\���n1iuƟ\%n�ܪ�ٹ*[���&�OL�k��ꕜ�U�R�ښb`��#4N��λ�b����9E�A1��#Rd�0��[���bcg�`����1p×qBz�'�YQ�Pۡj�I۬W 3)�Nq���;nB�޽��*'0�'�Gf9ߔi���-���R�J�lQ�#h*���jZR�TZҵJ�[J�M[��Œ��QVPQVTmm�T��lj4��(�b��es()��Q�-)QJŊJ�Z*�)YF6��*4U�EJ�[s.�Z��4��D��3E��*)kDh2�j��)��e�b!FTX��T\�Ar�F��khɉ�V)+
��(Ȉ�dY
��F�iUV�(��+ej�ZS3V�ZUE�U��rᖨ����7=Ǉ$����;��ITj���&3��MIPf�ύe�N�ނv�+1��,�.7$ʛ�C��S���et:1h���:��y{GuEQ�{�ҍ-`@r܊j�F�R���Y���=Cb��'�����W��l�X���M�ܮ��m�vl�ӛ.�e]���:���y�d�oZI�t�?M��J�9C}�V�,�ځ�A�'P��H��|�J��j����y9MpRkˣ��х��j�r-Lr�+g�o2Nn����A�>a��^�������E�sÇVɚv�T�|+�k�[�iM����I����x�!S��J���f��������6��ܗ***���~
M��y��w
��,5��kՄs�X�w�]u�w�jzb�,ddv�����(=�O���Ȅ4QY3�r�.�I=.�W&i�w_/uޠ���m�(�9��DҖh��*c��8�rH���}�g�I>�Q��G(WDd��`,ǫ��`��d���xV��Q�g���6�P��Q��d�S|hYV���8ڮ�^p��m�Qos������������;6�$y�V\	��y�����S��$�Lȇ�ڬ[f�=���Tu"�e?euYl]$�#=z��#����&��琪�{�Kwu몔iK��*(��pHD��m̤yM�͎҃�9S���iB3��8k�����m�����Mm�"���瘒�jz��0�𓤾�|SWC�ժUyOi�GPQ���.���L��f�7�S�vx�Bݫ��L����;�(CS\VEr������|��S舼��'��t#	>An�JRǷP��C�}�J��wB2e� ���[b���k)H�YyM���U�׎��Ӂ�Z��:XbC�A�pRsn�[t.P�E˙�O�NG$�]�z���M1:"��p`��ݼGw��#F�z�f�s�݂���0p^p���}�C���S��o��&�v�Z�J�m<��=�g�=�/$�O���O.R��P��Rh姅^z���m�@��1(I3K�	є�;iX�����b�aE��RRy�'�yɊ$4\'Sƅ��)F+�x�ef�ic;f�n8?)Za#x3Z:�k��x��i�G�o[�-� |Ҡ�#Ll�Z�3�ө'�V�_dS,K2�vxU���f����C��ug��\��5r��%ǙGwFn�Vt<���l�S���z���,48*�®XN�tJg�`��A�S��sl�H�����/o�h��'bHT�Ò}�2����E���v1�a���W����&�T�\�����{�؅8�K��t'KD=�`Ј�9��)�HČ�/�hE]&�ʫ��Jtb#'3rf0�ZT���z'�fgE�̴�~$J٨�K�Kj���t�.玟��N��PS���,���vz-Z��kB��F�Z�SHϑ�z)L�*�+Y�'���m���4�+�U�b�-���%}�Ҍ	���T�èð�r�^O>h-�+�ϓ��:>ձ�Do1����6�>�7���3���W��^�=]�@�]�J�{�u�S��z��Y�.2�<�S��
���ՔKz]c��P���nγ�Y�!:�e��}�v��v����b�[y��#秬=+\��A&�Q|R�r2Ӛ�on��=BF�$!K����E�{uq�yɥ��4����fz(� ��e�|*��Wm�قÞ˪�;��)H�(9���0�Vu񧶑i�Td�3FUͯbK!�H��@_j<Ik+̇ЏH%�X��W�.�N� ���,��z5(���LR�����FQ�b�o�Y��T#=��2\^���@�ι
Gl�t��(إ�����f��L� �C�B(�!I�v3[(�h�3/_ie*9/�Y��(��$G�#���]�Z���!֝�o5�B������S��Pqt֮g���{\���/oͯ{*��RH6/����̡H����3\r۽=���&u������+L=AvQӓ�r�u!�h���9,L�Nr���s[D,[�����✜��.���ջ;{<O�#�*��0�كo�5����f�C�l��e[u_b��V3J3�D�ro{sj8���8�x�
��.;B��ފn�Y���֞�Zn�C�]��U-�s֤�J:�>�΁��=�����bkO۱��(ֵB�?���h�<�
e6��=�������t�6���J�wukMff��R���7���VMe:nq�]��+�1��7���J���_�Ʊ[�Q�Xh5�;6v^Ok�����c�u�⟈ι=^��]A�^Ŷok���:�G;%���7Y�^�غI�l���CW5.���Z�M�0��O9C ��9b���ۘ�w�˗�s+7���<)7ٹ
���$#��F)�&�'�͞��.�y��˷{n�6���-<�j��Q�5�Bdregw ���]$�/����ٝ�gN$ڰ�XA��y���M4�s%+�SE��i�M��\��YsI�|%�!��'Ŵ9�WN\�f�)�l?�W��s�u��9_V��Y9^��q<ڤr�nOMG�'�c�Y�g+�w-�t��]�q=��.y�t�����}��S�����<!�.��e�]oo{���/N.Z`��Tܘ�o�]�U��Ǥ�Η�1��I�Ԯ�[�����W����՘sR��DT���٥H|!�o98���{��h�і�N�Dd��z�ZV��{G���_)�q��͑����Ua��a ���p��� ����:>xGv�x%|�N;�tOvEG��>�6�Z�T%v��b'B��&M/�2�_T�Ga�Z�P��JC�jGcQ]t�ݹ#�I{!��2���D���T�V��'Ʋ���#j��'Ԕq�e�"��̛sǜ���x|S�>3��O�k=�0�W>�9OO]�FA�HF�{��[Y�{�㝀�TXF�Kr�O��HU���f�E-yĦ��ܶ}�'�@���<u��e��5J4)�QB=�s����L�4R�PÝ����>�jG
��lRV-�1�8bz$R��^�b��-��T7>��0/%��7	Jr:9!���K�5l�|� �l���!#�n^���(��ї�!�Nl�c�Q;UgYc �b�����^���3p)�b�x�B}I�yq���A񊽙����u�pz�+�ZS������3����/W��d��Y٤�E^Hb&�$(C��L�/���V�hZ'K�wI����ﳜ�׀��+4��(͆��!g��wet:��a���t��i����te�����7�P�Ѩ7D��R�	��1%gDJ�nR���$��(����)bI*��~{~ܐ�f� �F�b�Қ�@�W���:�*Ǉ�RIv��*U��u�v1��� f�8���d����SCKc�Gk�)��u�PA�:Q��mH�*��㖾���	��g���ɽgIEt�6tϭ�s<@���i�ǡB�[�-��d��4���Ƿ�㞼��6��K:#
��������ρDu�O�c�o���E�דra�+�d]�mw^�x�bh|��"�3d�
,���o���f����hߪ�߬
�r��d�"�U���T%�sb(*��)y�/;
ibQ����,��q�zzz�Do-����ܪ�<'�a<�����ts{w�_���i1'U�Tz���v�vNz�a]+�o����D�%�E�\�(E9���Dd�s���t��7AT��z+$n������[Z4P�ᮡw����(�#u��f�����R�̠0��)�B������g+��+J�Cj��ɥEO��=)FAi��*6y�]�b��u�V)aJ�Nk��r���껗���,N��#Ɍ@�ǵ1��Mo��7����sl�^���o1�������@PA��Y"�Xo��vf�U^����nʜ�B���2�ߐ_v�D�N���\�U�ﷸޘ�7���_���
+fܱ��0��CS�H�[V�niTm�g�FtD��PR2,��tv�7�f�����ܾC�>1�tT�l�n^>eH��p'����)�S�kߪ*۱c$���
+����3:a��4��r��銞s�CG�c9����E���D�ȟS�#n���KRiY���E�5��,/�CM6jǮiF�x�/���Dg	e2s�Y�w�(ߖ�^���_�TEdܘX��L��~�@��[c�h*���}����#ƈ��	i����
�S)s1��	V|�#��GgU)���I!$�IEQ���TD��Z9���8	�����/�3
�y)�>�U�K�WJ�%�>5Q+@�
��@��B�hXn��P�=�\�P=��(����J$�fr����e~���W4��<��J�����Tބ�c_{��A��m�@����< z, >c=���$QQ�]������P/C����� *���tH��E��g�K���t̵!��[��M�3��o�:�(p�1���O�C����5ü�T�T+�|���1_������)�[��7v߻$0������ҝd�̠(��1�e}����w���
%� T O�p2�*�{�)���v����Ώ����;���QQKx�������5���Ūv턎cWO������ܯӬ�xu������ghZx�h
*"u1ƌ�v=���~a�����5ZQ�h�|8��9;�)�\�� ���i^e���!���Q5����p��g�q�,ԞI5�@4� (�	�9�����K�,7Kz`�
.�vG�M7�dbY(#��%��
�"^�l��� �R@��1S@1mE�� 7�`.���akRRa�/P��-V��y�5"R��qk��}jв(����u�9�� �M�"�%߁ԧ� 3c�X���n���H�#r~Z�r�G��k��f�y�9!�>��s�<;��_~�&)�������e�����#�؝�"�'�.r	�S����^g��t��P5�;0[\����;�T.#����ڇ.�3���p2���m��0�{�A�����Q7�J�pM�v���p��La��Րlբ@��Sn��r�BX ��
�'݂���
�}���x�0��TD໎#��x]��Å�xQq �
���$$ΐ�� e�L����]��BB�O�,