BZh91AY&SY|��� Vߔpyc����������  `�~�     �( ��X        Ϲ�m5#�@ y�D�(EJ$�O��)�\}�)RO��}4x�W���{�q��
>gH���t�+n���;d%DC�cωϑ 5�I���4��2���e@�����R_��X�f{4"�����TI��X�Ss�{��_w׼z�C�;����*P�֎쪪��1��D*PWr�vd<w�`w������]���ތN�Ԑ�Gˎ��N�^�:��uy�^�Ls�����D�oy�"C�Ѐ P     @   J����UR�M=#!�� i��`&�i�R�iI�bi��2hM@  i�U*� �d � 4� ц�� �*P�2h�14�14�D�&�@	=L&�"i��mA�	�&�*U4d��	�LF���#�"{��C��D>�~P��_AT?���QTG�  !�@�����"��6(V~�������ȟ�DD��@
�nO�*��!($��QU$������I$�~�DQ�C���/�'���������}r�̚�~�g�ܺ3�9�_a=c�->1���J,�9P��w�8���:d�A�u��+
�U�MU�ʲ�끪9X��Q��O�JOp�t�tpu�840%*c@��Ӹ�\^�;���r�:�]��88���O�]��8
���hXU1��
uv������W���ݖ��}�v�1o�e����ø8������9�Q�(÷�\^�덎���N�{��k��)_�g�V��n�a����w�P��o��xr�j�w��qQ!ޓP* [c�;N�x�\Ήoy���̮c�Z��r��{�ܵ�h���}�zʵ�-�6�[:M]g.��Ipr��&5��^�z�q�+8Z����(
N�wtJ	��hX.S�6�o`E+]k�tl���e��'Mp�hv{�p����O'��or�gJ�S�`Z���MW��Dx���Z�]�7����p�V˲�]W�:��	���!�X�o���������[K��5</H�%<L"ʳ��m��K�U�<��7�Ͷ�[t�ܩI�����,[��5�ÃO4�(��v�΃�����-f*`�NU��
��եQTU�:��qi��1;
99"���w�8;D[(%k;Ӱ�a\͎�����cTw��-Lpޖ����}е�������L`Qރ��;�����.˳z�v�;Äpސ�'a�m���hXR�0��҃�]þ"�w�_0.�vOX��fv��0 840���/����{�:��bW�Kg+⸺�1p��\P:tO���J�'�S��x�"��m��1w����U{��r�vC]��o�ǳ����:@t�i�G����;u���KYE�P�I�o[}P�3C��ٍ� �6]%��Q�r�9T��I� �	�k�ƨ�;G�:\��նI~��}����ɣ`�����8j�h`yv��5J�+x|�W�ݫ�U���P�z�V.�\-�O �*�W*]����x�)�Z��]G-]�'��W�W�J�m��F�X��G�7砅�k��a�R�rŜj�%ds{6��o��@�`F���J���0�5�ӽƥ�z��Zu���pr�=����>���p8������.]��E)\�����n�������f��z��&��QDra+�N����OR{+��ޫRk���ƍT�	UE.SG(��V'�,%��B�j���s��J|ck�k�J�39��Y�z�K��|P��^�>�ѭ���}���I�\�j!v�>S��gVg7�8����9u�����k�'5´s�V�M	���������|5��t!�u��J=U��:pʫ�8YIg
G�j��L4�9����x~����۪J�5�9��J��\@�M�ʖW�#pﲫ����ӈ����U�p�/�5�&��y(����ֽUbZtOG�t�7����窓ٲ��
N'��JN�k�"�8p���JO&�
��xP�e�{����������9l+���u*�X�URr��M�5�r�B���k}�w�B3��:��ZV�ޭ����Gʃ}Z;WE�j9d��W�´�Է�[��y#�W�E������u�{ۭ�7�[�vB���W\�帲�/=�=��rP��|�UO#�9d�Z3V��K�����7 ��"�\�3��#�f��2Q	��O�����^J��:j�Yf�Iϓ��y66`�߳�5�(Ĵ�}<�;;�Ӗe^%m5�%#�á���uF}voF�^��L�cW<*\�F����h�*���R�eZ�:Σ}����3����3��4�����K��n�ɖ̐&����u��(�|[Y�J�*�t���U�Z��!gK���84�0i�Q+��3�|�84;[r�l;���T�.x;���z�m�_�A.i���r��ݞdJxR�H��LITw�v�×����_�,�m���v�C�J`�<��=�m���Y�ѧ��>$����G�����!A���ǨPQ��@��+�&l�p���g�Ef���j~�2q�qEQY@Yd��Q���P?�P�,�� ;,d�2���i{���1�Ē2�� �M,��$�Q��p͎����,
;b8�)x$a�2c&�:(�-[Ŏ�(,��]ׄ�A�0ќ\J��
��8��H��ID�A���w�N�d�=ȁ�Q�pĔ��zaƐQ�$geLM�E�F�z��&z4���1LG3o�M$�PY���8�i9�I�,}ћѥ3H4�8���:G	zm�&�nF�$����c8��0;��سM�@h��/iE�I%>��}q��e�AEYD�`�$g�H�A�ag���d=� �,��0� ��I$�AEq�ýZ�Q��qQ��
E2�d�P^�A%q�;4�N�6v΋������=��� �,�� 	 ��,F�Q�A$IF��P�c��1�f$��E�FA�c$�@iD ,��8�.�<�$�IfQd�z�c@g38��M ҋ 
0��O ��4�#�4�K'�,�4� �Fi�J�Ğ�K(��0�
4Ê4e��2I4�4xi����K.�	,р�,�� �,���  ��82e�{G��d�GQD}�+A�҉4ehAC>$c�OɁJ��v�>0�K4�(�0�(
M8����8��P]tq!�4��TA�|Y��5������q�ČË0�y9#��
���(À1�I���.,(�F�@�����ɐ8:�"z(���(Ɨ`q�p�3J0�V�	(eAŜtT*����lGƜQ�|h�((��i&�I�iBW#J	��I�2FQ��Y�Րiq�A�Aj�y(�bFMF�	��p���(��`�\8JfA��*~�4�Cf��Et�S�YU�4ݜ`�iR����	eW�YK��C$�B�q�� ��((Pb,(��fP�6`E�t�$�@��bc8٘��(3"����c4�N=����.j�bJ,��<��]7%�)�}u��|q$�XT�OE$��zU����2��ycxq�E��I�h�d܇�s�ctae�y{��D�a�S�%A��|� �g!�1��;�O��4�6쉭&r&�|%��Ϯ� �%���� ϶��9����<��\Da�t\����6�$#�I,�$�Q:׮� ʸ�N�+]�~�q�a��Ճ(�=���#������:"�(�����$�C�@���ʭ�ٵ�aE�&20|nѲ�8�0��P���GNE�5iԝ+�@�^g��R�&�J��F�Q��CNƞ���L�� �)�|I�3p�K��K����0��/a��u�P`��(J1�Lw]�Z�n�.$�M2��$�f�35ٺ: �
�Е���.r�&.d�1/]�����$�٧`���`Q��� 3L<v�)8t�&�m�Z�d�֞0��Vi<�v�ļղm��8ɗ�^���\=w�)�xۦN�W�,&<p�N�d�Zdy��i=���=�2���P04��e���U�zOh�>��ȋ$^��k�$�k�Q���I�s^�KT�@Q�2��{�Q.#ނ���z����N�}���%����?����z��6$=�S�J}m�'��z�1�	��>&L{�|q�굛.�0�g�o��1s4�v_Hc��'I�H�2�\�69��l��⑓tPe�Bc4cU%1T[B�A����� �	�fb9�T�R������y,P�t%���]�E��K�v�E�y�>���* c�k�RI�UQX�U@��+5a!�(o4��\Ai'�K���L�Iyl5�P�W�)��n8�ELC�)��pP����WWB���r�ppR�BaL0�M�Y"�(
/��q�Y�/p�(���D<��!(@<��Oz��H�/�Ȳj��&١��h[�	��PA.	�70]@E�Z� �X�詟������ _+("
%s��$�z��=��::!�_I2g���Y�C��ǭ�W� k��o�~��/�}�]6��W����W�����v��+�Uq]����UmW�J��J�[ZUUZU�+��+�Uq]����Uh*��������U^��V�x��W��fb��UU|Ҫ��Uz�UWڮ�WU\Wj�U\E]��*��UU��UW��T>>�ᯏ����TUU|Ҫ�WJ�kޝ�sTUUTUUTUUTUU|ҫ�V�UW��W����8s�UUUUW��zw��a�@RA`�Ԅ<0�I	"������Us3+3_-*��iUW�J��EUUEU�^-*��*���i]��*��UUV�U|��u���>���>W�Ҹ�UW�J��EUs337��+�Uz��U�t��UҪ�EUq]��Uz���Z^o��ۊ�U^��Uq]*||*�U�j�U\ZU^�ff6��U�^*���U�j�U\ZUW˥]��"��WJ���/[Ux�ڸ��[U�8 �yH����p� P BH�H���������`*�|}G����|������t,M� �� �B ���(DN�tN��<'Lg�t6"P����b`�:!��xO	��X%��؛E �� �<<Q��x<�O	���8~����I��׋�f�����c�ѕ�U�u�p�2����t=�m`XፄX��{)�˶[f �fՒ�%�K5���
ja�؆[[r\����[�Gv�Aw鲚��,z�nl�),&b59��6c9�bJUч��F�6nnҚK��[�ᶴ.�j���rkf���:YXjҐ�9FaػRAm�jkF������h�j�ֺ�[��h�2�qXJ��F���5�-�v�#i�(�>v���h�����9)d�f�����f�V׈&��mM+�1�י�ʷ���Q΍E�1ι��ycn��b<Ĳ��uvAr#��-%�n��#��КGl8�؎m#�JGf���k�H2h��ۥ�@G.񁆼E-��F"KI���i��s�2�
1�)������0��lB�*��ͨ5���ER�Z��ω]�Y�cR�F�0 ���6�
�Xݎ-�b�H2P�����%�m�fkm�ܘ�k�[b�>�������Vb��V�M��u��s4kwm�EH����:�M0�N��V�lH7:�Ύ��&��e�����^y]LGRh����̡q<�f
��pF�H��^i�s����g�ѭ���:�8ce�b�E����7]-�f�� �.��6�W�V�)KE/<gL���D�3Q�8 ������1�%���h��4�h��h����`�Sb꒷A��s����]a8���&��]��k7
*�[��6ٛI�J�i�ܶ��	���&��eb��v-`˴�"��`Fʒ`)f��xWt��P���2�e�Y*��6�0�l3%��eCAԤv��->�z>��q�L���1�R���9M6m;̧h1ee�"И�jK�i`��t�	���(kγ4Ѭ-�ң��lkSh���,M�qn�-"&�v���4#�N��{)B��p�Zil� �mYAK2vԠ�j�W6[mV+��ZVSF8����,���hr1����\!��5�h�vZ�Ѵ惭V]jbE
`�Rxc���S^U�tٚ\&�ƥ�6�v��,ee�R������lt�R�f���v�f\�ֈ&csu��XB�2 �Yf.��Y�cm([�h���b%�H�h4��50藓T�V�Q�eD{M��`%�副$����L��ml3��4uA�k��D�Y��v��*��G:�cfG3��n��YH�9[���=�!S�u�syWL�+lA�H��ܛ����3�����u�	�{.ﱟ+>����I��w$�+ ���&f]ܒ|�� $��wrI�����&f]ܒ�'>�&fg9���ϫޠ��L��3'�>�|��)5�Ch;�[A������E�љP�-�ir��C2�i���-�z'���}��X�F!	�����n�tp��ڭ��˺���bk�N���Y�Xh\��yM���[���il����suhؚZ�hK2��Y��"�m���5if�.���Ĳ���`��ө�N>�[����6n�E��(U���)�M 5���,����ؕr��A�����f�!ز��ij˭	
��m� �"�S���|`9_�V$A�D@J���ǭ�+a^F�JZ�x �V^aW%Qg�Iq���N��|r�'����(�z��UE�aa|9�5M`���s�d��^���Tu:u*bn��Ɔ����Ĵ�#n������*U;�.T�C�,((Ȝ(ѐ�w��*誨6鰶��iz2�'n�UKN%�PK=|�WsS8[�MʆC==q����H�`�JN�#��+��S[�*fm�dJ4�e�YwV�*1(((��2Y���Rں���Cm�xi2�8[]c�I��+eV%B���lL�����J�4�
%�C=�TLJڏ����Q�Z�;*b�:�Yuy�d�`���b`�fC܆*��*u���sR�aڕv =j�U����eD�'D��ӧ 'P�`����&�:Ӏ�ѬL�C	s�u�Hi��J
�
U(U�Wk\�q
�S���*M5XA,� Mk��&�4b� �l�%�c+����E�=�I��\���n%���Փ�G޶�u!!�M�v� �ďDN�E�s������7umUߡ� 3��UVB�*QCR��J�Q��z�

6'��d9yC/�8b�`�u&����vU=�$��Zt��6�fY�&��M�\�1
+u��V� Ű�qk����/X����*�U)�z�:z�a4�bdۇh5��ĝ9hL�,�9t��]SM�L���өrf��.��ܩӰ��{�6�L�srˢ�XQbjb!�P�J�UV�� �ܿ!ܫQ2&�$�M�*��ne�(((��6Y���U%0Fƽ˪���;r�/n��k�zI�pV}2��4��Ci���A���M�Ӻ!V�%C3�aE	ҍ,�g\���5��!�.!��*ZSN+��ษ���\'jn�˭�l�*�Rj�"2�X�e�*�UAB�&: ���4����Q���P��b;7�����\B,��� Rፌ�p�[�2bWTa.�j��g�O���B�fjb<b�z�-0V�y��#�uZ
(N�tvY��\�U[�t\�P�0�n��vw��͸��-VM��M�{���惾��3m;K��.�Mf;��}�N&d���!o���<³�W�G�6W����t|<E�J
>�����O�O"x��D~�(G���E�4|?G�<l���|>��epv��%>���QB��G�xh|���}NJ�Ҽp�9O����|=��TGDф5�B�p��6C�>��>+����%�|'�G�cF�Z��(�xQ���B'��
?G�'��>@���z����C����ߎj�cއhvi-���7�M`����.�\� �D�A�Ue���ӱ��֔�p�B�l�e�D��g���$���"n���8Z*P��%�\ד+�T}�}�>��������T��&�ff\��ܒs332I	Rl$�/33$�jM�&^ffI ԒI}���$���<Q�ř�ZEQE�dI*0�`p`ۜ�\�.�uS`�w �zK�dF�
T��HF#�!N�D�-D� �L��*��U�HN��Ӏ�	�LR��I��ܢ�%[t.�)�#�t��ye)�1�m"u�`d�$�I�$��8 '-�'X4�eL��b��C�%��:Q�ř�];�9EQE@�Ta��P,f�%F[bo4�lP샺w��\�%J�嘻�T�hGm%Ӷ�$P�P�	D\�pºb D��X@�!P�aeJ�Xt@�IYQ����8DN[N"�m�(CÁ$`���4$=
�?Le0���,K(�G��d4yS�j)
T4홺r��,YV(���:7��ic$}���D��������XB9�$�Nh��
f	�f�����m�l��Z�%�T^�א���6���ǡ�Zuh9��M��Z�&4��(l���<q�:p��zϏ�4b��[�F��bt(2�}��1�F��g@nUC@Pm5�9��.U5���S.S��؛�4xĿ{�^ʎ�N%�C	e(��̆�>�����EQE!�R�'�-� Ô�I&I��ɧ�Ҁ�Fw�ˇ��[�*Zu��dp$#g}�
����8ӕ1D��W:�bV.꤫�%d�;�ڑ(�X0���A�:`m�֓AL�7����f�τ�YBYF�<|Y��o�ո�q���c&��(���ϯ��� |�|�\�(�e rQp��f���@�&�w˅��"�}Hҥ(�������j�< �`.{����
�����P� zrsE��h�p��;|Me��x���6�$o�w�`���,���|l�����M`�[AS��Ԙՙ����,���wG�:5��R���8I��a�r��*C`�^r��z���}�t;�L[kF<&\��l��`��qԒk]����N��UUPi
p8b��*�5 ̅4dJ��(�fΖ`4��+��6�󉠅�ny�Q�e.ecV�v�4�YF�2ڜ�Ք@����k2����f�e��)\2V�@G���k6�Ͳ$K�f���@)4�v ���[o���������N���nN2���td��`a+�CƜ�7�ĉn/�H��X�a �� �V�=!�+j߫��!����lt��tb�B'oT�H�!��v�5�Y6C �YE,ɲ��8�&E루�Oc����<�U�Zs c;�n���j�j�5�Or��,�#��Њ�L�
��x��0�yG�T�XیH I�y�{�y���d��5�|�d\��(8��|:Y`fs]���Լ��d�(�%�<Y��:�j��)aL��g�몪�
�d*F�	I�i�6�M�O]Y�!���XU�8�j9&I�guUvT�\����&%����r���}�J7��4m�hF���]��J�;5�-�,��2Y���CEۙ!�+R5te;�})٪oe<u@g�*U^������c�Z�%6��/U�� �1�m6L����\ŭbUUIU���2i��d��ы�[�O �np瓼ԩU/�M�N4�C�>L�n�a���U�+��86D��^�|t��t|<#�`lO
>�J<(�C����O
'���D�S��2�,�~�|l�	�:W���xp�+�D}�'��xg���4�]���ڨj	�sUIP������⦏��>0Q�ʡ��M��|�,��|h����D�*>7J"hD��*"xQ��(�"'�'�O�+�f~7\�J�������"����]�K�U(-�<�%����4�����t�oaSn�"iГ�2iP����MT�t�ۓ��)�5Dj�wSQw5��+l��RbwއQ�ɺ�ҩ_u�6�z!AOO�/KiZp�r�~�FB��fd��$�����H5$�_s32I$ܒfffd�z�6I&fffI'��I.���$��M��F�4h��CsI�O�|��<eH�4[Kkf`���d�m���i�}<;ڍs�l���m��W� ������@�xB;�*����hKb�R튍�Hki)\�.n���&
�ۄ���p^���d,��ˍ�O�ۋ�٢�L�g,���fVe�2K�6�m�-4.���S-�L.�F�a�jb��Z1���IFZ�K��(54aq��/�޺�X�&.0#0[0s�R�˵:�Ϊ�-�ɑ����������p�:6aƮ3�Bk4�'Oy޷�Gi�V6%����kMLA؉f\5��F2�Ā9�kKU�Z�]�CE[V5�
$p�a�µV^O��.�͎�!� 5չ�ʝ(�G|gX<�Ud&�p�@uTM��mxEZS
pU�O�z%/�_���语����ED0���e�bx��0	e�Q��,�h>��}�KE��������9+Yrf�����N�M>a�;,�0G j':�f��#Hom�>�B�b�@�ئ��P���Wr�nʤ���v]�<DL�s
���T�p�_LM�Yb�n �Y��Gr)T�F��pf'Bp�&�6h����H�ŀ��C���%0�	��X�UQ��bh��K�8x�J�i���6yL[uM�Z��.e�J"O\����w����1���Z]�*z�UK�<�$*2ɑ�K8�S�ɦ�%�p��n+���hLP�>Ξ0`4XL�<d�VҦo|�&�;mM�:%� w�JwZ��(j��bh!�b 73��s2&��݂�����v�h�p�����S*��xJ�`N즹}\����<L�H�a�%��J̉f�0^u��[�}Y�ܱe4�L,�_t!��N#T���v5,$�H���L��������RP����+��a��X���2�dy�tg�* xL����{̇
eJ;(�HgR��^3�<���b�/� eL�oXti˅6:;�a)�w�u��"�&߁�C���@V�M�M��w�C�&x`�	Blؖt����}�<-q��(��@�:lm��>O:�kCni��Ó���G���,Zg$�;��g|�A�"T�v/�e4�T9��V���y���UC�9�\h�a�τ����lك��k%�)�N����řP�!=G����l¡����D������-�S�) �YL�TD��&���$�:��>j���	���ER���ɐ�Ϧ�F�pM��u2X�	B`�l��p�[��H�Q��uO�(�������#�]S*�m*�ոd�391.Ȱ��}5櫷vT�����Z���qjNP���F��<H��w.ʪ.�N;���e�<J��pL�P�x���0Xh>�O<d>����B�o��,�Ka�󘆡14�fRX��cp�CmL�I�ز����4E�1V���[�3IXͨ1MsJNߎ�O}��!d;V��l�NS���kǱ,zC���
Ci�[L���E �=wf�*���0x���
���O�y�[V[=�1%�m0:�&��Pi���L��J&�(���A�REM�B��4�pv�k�'TUe���`vv��'UU�懢1�/�Jn�ٞ���}�YW[1�V�V�eZQx�^.�UH«/po]gYM>~H�r�ԭJ&O	�>��և���tJ���Ӆ|'�|x��t~	���T�^xQ��E���xQ<(�b?'�O�+�|8���Z���Z�x�G���x9W�"z+�O
>(���jd4a5U���Z!�&�ID0�O��Ҹl�/�48<V�c�ʡ�D
 x�
��h��D*
!�:_D������b"x�|(�D|(�
'¯����S��WᚻB�
"@��I-4�Z��].��sJo�+�ۘ�Qq1>�p��D�S�WJߓy6����n���"!ۼ���w���q���DR:)����*����$r<��2;�	�;��*�o�{�}��fd�Q$�]�32I=D�Iw���$�I%��3$��I$�w�̒N�$�]�s2I;D�QF�(O,�G�����p㹞�E�#g��:r8>]v�2/O���$���6�wCuUwv�ފTst�8|;�ò�&��8e0�|V����5����,�OP�0Y�G���7�f8m��sJ�9�nޥ���4�_3]��Փ��p�U�Tf�b�7�[b�i:t��]8:�:���ux��|#�&4Z���P����X�����J�<Q���׬k_n���
5�~q�S�)�X�h$.W�8ûBޫ�LU�]�l�#t�M���IK�֭��,2Դ��+\Ѵלx�x�=z7�p�%�l�$0���C�liM<�m�P�;^�B�{��UEU{0ܯ��ޣp��N�K}�c�5u@�m�tXULoSNMo$؁���qu���D�%	㥝(т�AN�"x��i�;1����bbꪯ����&P�Ge�<i��}�;�zl�?;6�r���Y�̹:,i�9�"Kn�9dbk��Q�0	Bl�g�h='ܮ��(�D��Er@ɉY1�E�}\w��D�PL�ϯ�砓�?#r{>E��`�U]���j�c��xI�XU�p-�"N���p�Pքh�@>�칔�Y> �&J2l�C�����y6!�@rSE S��9�*���8Ywme��ᦓ�y�s�����ĭr�wWX�����;bg=���L<�P���Ki��,��F(�x��t��[�.3z|��Oh믯xJ[[�צ�X���,�	-�QM���e�f�l24f!m��o�wm]ܦt��\��.��M�h�eNO�l�G?01�<tQ�I��R#�]�ѕ��������$��Ϗw��k�D��d�ZFT��LY�W�a<�~�K@�'J2d��A��=4�u��o�5�����sT%_��'i����ɶ­����ʽ��sO�5�)����K�_(g�&��p~l�D]Ȼ�k��������"n��h�R�IG֪�s��2&�(K(���M��Q�BII{&����v����_SUW_K�����
z|���UT��N�y���C?IA}Q��qܞ��A�=nk2�&Z��JC-`*qJ����ʓ2���� �'
8l胠�O.��Ys x�r��B8���[8��a*��P�Dq��ۦ׭���v�B�QeZiA�H��4^Th��\��\�TskCc��x�|3��/�tO��⍌��\��G�J�=��|(�!����~�D�Q�TO����S���>��||p��x�>*tM��4�z�E�C��F�yY��x�>+G�O+��B���`��	B��7ㆲ����p>U)<��x���^	���GcC�舘gE:P�(G���Q>|�����ri��0s����ka��>�"���{�.yK#6f�J�m{a��4���Bc����Z\�8�v^9��0YQ&���N��q�Ki'�A�ˊה�8fv9kn���מ*kb|d��r�i�Y#wjs��uz�˗^9[��\�[s3<��$�K��fI'h�I.﹙$��I$���d�eJ�I�w��$ʕ$�.﹒I�*oE�%P�(��@h����V.���W�n�Lh�񽳥���祶�WjA��MZ�
�y��.�T�v冴�� ̫V).��-#��@���16#"��y=�@О�Z��d��Վ�t����sXMk�R�Z�2.j=e��%q�����!�аL��u�:R��[�_z�Y�fĽ�$n"b �L�&��m��F����1��\i��X4Ŕ�7-Jnu6���f�q�f6v�6���$�2zz���p꘠ݥuH@mlt����!���m���@*�JL1s�j-�(
:Ya3b��E[�����vf7��hW��|t�NW��Y�A]u*�H\����<I�yi*�0��e<7G��u}(���c�a��:a���C��̹p�g��J%6��}wM`�J�C�J�5�no*��>E�f3Sp�4�t�J|:N�5J�ă���u/���R]+M�X�b�w}�l1E2��4������wӻ黒�(�:���'�>4��C�ŜN b1�D��ON�� h�T����3J��}<Xbu�i������L��;|^1
G�ĳ�'��[���������m��1n�B�F

(Ox�4pU�����'�UT
h��-"h��'5���^�P�26�L��4�U*�f�)��o����:z�	b�>`z�)QnLM'����P����L@jn&Ed���
(K(�`h��y�+	3`�N�|'�V�m�5����;Y��kz�и@�Uђ�롄�a��(�R69B�&x���M�%�HY��R4K*jg��\ä8{�S��l7����>���ߖ`-un�P'��:����O�|z��J~�,٠Ѣ�4xà4u�k��*�e��S%`2����V�ml�U8p`�M8�K\U;|�>t�~�%��۷�ݜe[�����}(���o�eYUT7��b��������UUT��4p�AE	⏍E��	L�Sļ8�b3$����3ģbS��φ/
�[��⊪.�f0(���n�11�jrYg`��*��	��_�uU�_�����OK��ꪪ*��|��6h����FNEꜴ��$�?M�J}1pg�^���{���V�v��gKdJ�	i7FG�H��-�ĳ��JL08�x�\�Wt��"񳳢���<l��>�_y����zٟkL����r��-<��b�jb!=s��:�5���XƌmJ��vX�q���M�b�Q-��Gnz�J�!���}O�d<��-0�&N�a|;�	ـ2�FH}�yوz!��D�Lr�HjJ\�N*�Iexi�nʹvY�>�>��'3�kT^�Ѫ6u4�hP��r���T �J���nb/�㊪)�I��R��Q����k�Qq#	~%���3RK;"觶�Er�vJ���Q(i���g'����ɐC�&��js����L�
<&���OdM�����T|(��H�|(�C'J��H�
'��#�e,���p?�d~���H�'���:3c�4�z�E|(����,|3Â���aJ��ڨj	�RWHi�'
��Ex�.�<6>��<R>��^����O	���Dx3��,Q�z"t��&O�F|*�|">�����|�w(T\TUԄ��
O�v�X�y��ԵZ����O�!�qhT�V�pi	�B�0�6b��3��g>/���(��������ˣ�s�Z���s�nc�*I&]�s$�*T�L���I&T�$�wwܒK�5$��wܒrI�$̻�䓒M}�F��!�Ggf���.�[@���BQ��˓)]�4�?Z8���I� �A��pb}迎쫤�wmU�W|i���ͱ9\Ի�R��-��pu��b3��ó�(M��y>:PQBx�͆�*�_^� �b�si��5*�+kܥ�߱�L4�b�{�3gL��3�f!eT�s�N��U�1蝌צ󯒴�A��Ȇ��`"l�aE	�G������\�o_}Cz�œ��2z^��og��ʜʻ���R���*����� �]j���[n��0��+Ιݫ3�{�ͭ#T�EE�P���7F\�W�KUTQ*��p1�=
2Q��y�����#����}�jLz�yC�M�cS�toc��MĻ������"�鲻u�s$8n��gŅ'�<p�h�x�Q�(��+��������dŘbp��`��i��8F�)Eq�X�>i��Uk��K�Y�>�u�������3*v�B�J!G
(N�d�Ѭ��cnI7L�ّ.3&�F�qW2��kQKJB����/�����yI���a�x;��%�s�d�b�����^��Pɩ��edL�d��h�g�&I9�qF�36��ġ��r=�rݵh�*�]ܺK�G����|���*C�<rT=�Z����nj8��� ��Lu�����ggl���	bh�g��z�M�5�+u���E����N給Ҿchm\�4��̳.�Kx�c���71�P�X#ne.�6�Rb�ķ f���ֽ1s�$�����lYV�g`���f�+p��ӓD.�m�*�(����!�Oh��Ɏ�F�%C��`�!�C'�Ƶ�[YBXٖh���c�>�&���hO�2h�h��}WT���5eHZA^�:��ʼ�e����F�^�d�,UĈaÆ��˳���5pj�e3/���PZD��wR���ǌ
M��Q��4%�6h4wP�5S-�nI6}{��k�i�������Stc�)�:+h�9��D�C�1Yn��UJҗ0{�90Q�x��#X�X|JHx����1��J��i:���	�4��+�
t�� ��+0����;e.2م�E?�4#(�,��ae`d�÷�͖u�h��%/�/i�n
���嘌9�����̆#�|=��⎍�>.xO����&��dh�B>|(�v4>|!���D�Q�D����O�p~���>*|;>(������:&��Z<P���|">|V�D3UVCP�P���U�I^*�)�/�`�[<V�Ʃ�I�'�(�eQ��>|)�5��>�>z"r�G�'JFt�'J�>C>_
�(G©4�ȥ;��}�w��V�s�*�Us���<��P��I��v��i��T^_��}ϩ��7Pb��d��Wp��=[.s{ji[�[6�n1�lAx"����%���<E���ɖ��ZL���{���5�*e^Z�����(�˽�1˻����MI&e��$��jI3.�$�nK��2I9$�䙗�w�NI&仾rvI�&�f�46Q��W֏wdՖib��5��һ���a���{�iw��B$��(m�6P"f��ñ�5���c!������b8Z�ܕI���T����ȳlL�SS@�0ԸW����4A��4��6�ԗ���>���xX����Vj��]U�]����Di2��K�$a�pk65��% ����k���!��c+nFR�Z���B.�کB !36�,]�+6+i�]`���y���{g�k�#[��(�v!��G��>�/�*D� e���d�~{����zm�8tpbʦ� �M;�w����\}`���#�,O��F�.����l���Cc��X�Ɔ��7��{��跁�&h��O>t��K.����U�s��%K��7IF��9�4PCn#���)�ۢ�2,F��a�Ϛj��_�
�:s+JEY���Y>����aAE�ҏ4�>��u�1�L�U�F	�rRb��UK�a��InT+G<�|Y�t�QIU3�M٩�.\1c�4�4ʺ�tU���N`�u��Z��5i:i�fq��3!������4	]+��4�������^����H᧕���	�αR����P��ɊM	ʪ�(��l[�XN���(�C�����a���lf�c=�j����!�AAFD�FO�9�{h7�q���%Y���d��洫a�S�T�2t�J_U)wE�]�)�*fl��Y�s'��� �e졌9�����CUML&C���7(����%�2�p�e�%:h���ܨ�������o��>xF�16��C[m�$Il�p�L@#W^Y��U�{������1��Jb$�l��ϙT���2�Yl@�cV�^��x��]��^������*��jhy����á�^w��wJ�]����&f��K�9��I�X�Щ=�W9��Z\U�-��Bh� ��$e�;*���O�&I�Ж|�z~'�7�'���c/�|��D��ʛ�5wwx6$>�UW3���0T�����U^���m�1x&*˼U�7I���ǌ^2n@�rtvѓ�$�i��R�7ۀɐ��bl�F���F�/J�|��'eɄ�CHff!�+Ψ�L!�9)k��5_.+���nY��Ӂ�Ģ�xԜM̔b0�E3>����M��*sϹwh��g˰�5�E�


8&�2t�Ws��7EV��`��ߞ�=+�}~����v�s��qZ��0`bs?c[*2b����`���`�ײUo�P���"T�f3�äw��'�g��x����`kV�K�k�U̥0�����,n�L�v��4G/{|�,�M��r�	T4-5XŰ�;h������^�jKK�.و	.���z�8���h�LBh 5���f�o��w���ǣץ���U�Q��
�oM���ɢj<|\x���n�uj��d�M�כ�%$9�˂����mv�%�[�k-�1X-u�'�9��C�O\,6PPQ�(�A�r�=�-�|u�5M_��`�F<�FJ��K����9��CeJ��Z��w�U��{�f���
�:YsY�ӭYWv�9�`�_Y񳧍lpx�Ύ��B �&���A�Cd<B�C�!	'
C��	���&	�<'����t�,K6&�	��A�hD���а������@�'
��w�u�U����*%��I/��#q�Ƃ�y2N��VމY���>u@����ˋ������Ô�U̝��-=���n)��v����^�m�S����bS����;=&�r]�9;$ܒnK��'d��I�ww��&�r]��vI�$��w|��nOPQaAE��4���<}2pa�^�\�p�ԡ�ӴS��,lF�-Uv.}>��RuU6p�
����.�`�r᜼��q��tNp頭���"��̎U)J�Bse�(�{��2a��1*��5��2�� 0���5r��xj�����z)ƶ�Aѣ�Ȕ޹��U�>�
�,.}�cx�]��/m���U^d��!ۇ������F�V��_6ڈtJ���+�;��Cjm�EJU[2P��u�t���5��P#]���-4&��j,R٨]e��8��*�춮�4�M�M�ZxlÃ��X8�ǐ�P����=�(��j��i���O\O�����ƣ��f8ӁP���RR�z��tOp٠gyEg��38p�Tԭ�0T񈹪�'�������(�a��9�h���*�J�A:� ���>$��5�A��NA<XPQ�0Q�Ƃװ�}�]��#���j^���+=��0��A�>����3����՝8�������&�vN�rx\�5��AAF�G�S ��ZӀ��^��|���uM]]�	}��U�����UT4��U=>4J��QgIV�i��e��Bjl,���"d�&�s���I���gE��Ü4Ά�h��J̖�!�r^�e�2�FB�#�:�������6����V:ف��.��s
%�F!��X��Q�M�r��g��:��.z}���(�������i]Nt��.�3)-Qi.�n���რO2}��ڊ#�Wd�

>�4烦/+.�QE^1����c��lk�V&�+s���Q�7�w)���n�S�ړcc@�11�h�t��B�E���$�^ݧm�ލ>�I�աrj��KjGBb�69�'�|�7�������7�e�a����c={�|K=��~t�-�A-�$�Oi�R�
ш?t��p垘�5թ3=�u��4%V��a�hߢ������AAGD�G��e�x&�h�L������SL̩���Z�O{=�ǳ/�%�|8o�?��|��w�bx�{�4���0�	I|rc$���]U��+�����<t� ���ѳB �xM<�P��Cd!��<B�a�8Q(؉�0K�ӧDO	�<'��F	bp؛E	A�4""a���x<x<��r�.R���Kq�*fѻjU'5MY��[L��Q~��w�( i�y	����uQ*��gC�ӝ��\lR���Q�M���y:�\�fo�����ɍ�#��g
W�[ϦJ6������:j�4]�ɿ^��X��pLLT��U�y�vco�n�;�I�3��H�'���U��F�(�Kv�X��S�q�}�S������$任��rI9.��'�ԒNK��I�5$����zMI$�wwrzMI6l6PPQbx�Ǎ⧕�7Ku]�/�(�4Y�֊ U���3=u3MrĬZ65���%j��y��LÇ�k3bY���IFeNf���J硯R�v�6f�M[1j�L��[�b�6�[�ha@�F���-���ѥ-72��f����o]�!�,7��\m���f�V+�u�c����!,#XX��a+S�-�{��T-Qˮ��� �K1ihٸc�#.hD*��!{WX���Y� T7\��P��S^.�FƃC�T��;m���%\C��;Rj.��K8���10�e���Rh@�ΦY(X��,X���I�)���5�����V���>��0릓�2z���Y,@�F0&����<����q�j��;���K��b��X�1���}K���l�7�N�,((ț(��A�jC)5t�H�l���(����)`b'!�0�о8�=A���>�n�>��d��[�i��o�k-���^I���c8��]6�4PPR�+Mb�i8�mD��)|TR�kҶ@�0��4���9��r����t�t���NZ��J�u3�E�1p��W�s�u��iWV��C)�V��w�pѣ�(AF�FMr#Xm���%�4*�.����v�QwC�fg|t95.\=b@���s
�x��X��6bOJɃ�O}�7uwv]����h���D2Q��A�pyU'�rB �Җ�����}h�&s��jl�A��	4����C${\�MB�E��l�ev�%be����Lx����g;/���
/ن��vo�{��\ZN2�z)��TSX0�;�}�iil���uZ��>�|'�>:h*�2�����`�O���>�1�xx�4`u�e��9,��yj֋�Yxj��UUӗZzp� ����$�["AưF�?�%��i5HX��j�ܧ����*hp�SnDm4�Kۇ"k�nT���B��7�Խ`��Wl�T��KQ�U@<��\tm�"&�ˣ�&�5����Ís��XƧ�^`�\5/����֪�����p����`�&����`t �z' t�$�e.��C.LL��J�g3�<*j{�5m_�(D�lk>�Ym�·=�q���׮���}+�Pf6v3Mm}�t]�.Ya����+�Գa�`(���bhА����6]m���Sۯ^����s�}�����ڠA�Q�����4
b֩��%p+f���m���ke�̓��Q�j�j��[,yg��{�w����dSђ�WD���=8&[<#^{H�x���ty���r��U4��n�G��*r	C��j��J�4d((Ț(��A����\�*�ˬj���0��h���OO;��*T�`��k3u��!�;�t�(������C�:-�����-;x�6t�$ÿ�1�����~6l�铧J2t�:AD�B!���(C�Ql�8B	�!A0�� @�@D�8'K�5^:p��<�xOj��,Nbh�A<&�	�(�t6���</��H\�(B�[�ks��TdPȻ�&�R�����m�n���Q6��i~�ݷ�Ob��o�}���ݢ��>r�l����zr/��ު"a��2�q��D�.�Z��Z����E�z+ڧ������3~��{$ԒIwww'�ԒIwww'�ԒIwww'�ԒIwww'�ԒIwww$eI46(��4Тp�h�h]f��q^���߅Y1P����M�ߖ�Ŷ���n��(6�4u�S�d��;ׄ�U�G�T�1�tP�p�PQbh��C�	��Ed�
yg��a.�q6l�it��珿��f�O(��br�o��Tc�J���6����f�����;u����@��PQHV����)]+����Ey��/W�Gl����p��e�	��r�M��D�{m����.n��k��в%��{�ί��yɇ.�յL<{�x=9�nY���j�3D(r�C�?*F{�u��3z��=�F��Cn�>�=E4�OML��3��.�Jn�������0lLx�Ѿ
�CW�Lr�kV䐼b�7i�m����=��V�&����v��2Ǫ�����T�9�����V�0j^��7�3���&mG�e�,((��(ɐί>`��#�:x�f�&��θe⡍ɤ����L�x�+�Q�m8N�SU���֣�dW�G���,�3�pLh�k8�EpL�s��M�f�-i���k�5��y�+1x8t�2t��Q�l
8D�D��L��q�a�a&f�+ǉ�Ό ��Q��l����l�FA���z.�u;��n�ؽ*�J�әdF.#G��3�l�#sb�inM !�� ^���ڨʘ��V+at�@��ń!�7{�{�va��[2�F����<klo:zmﶕ>��N���/�K��±��zs����3�|����uwj�Qc]�<㴎E!���1�^�wZe��Z6j3�/&�^g~]�V1XѦ4��	Ii����
`�Mrc��j��]c�u�
�OOJ/G���.�1:b�n?Y��h�PQ�8Q��Β�U.Mz<0��nm���a�7���Ue�*ʶU\�L&��8�p��ŵE�2������p�]�y�0��]<�&���0�d���$4Q�!C�f��k̎�cc/FN�ۯz��ko� ��&5*�U��i�<z�XN�zr��HͻQ�	"�1	$��=&y�
� w���?����	�{��I$�P(�����?�����I��?B�d�8Dٚ(������7���q��QPC�I/Q*�X��`���X�A`��"��$ 0X(�b��0�@"� ������Š*�@1� 1".�!p@b@H���� ��i!H�� 1" 1�!P@D
�D "�,
 0@P ,�B� 1�
�.��!q�	� 1�	� �� �� 1��\0#DQ������@`��@`��)$(�A����(B (	��	�!
�D	 1��	!#H���$bF$bF	Č0H�F	$`����#H1� �H1�`��H1��`ă1 ���`� ăH0`ă#1�1�1 �H��)�1H1�`�`ă��`ă1 �1 � ��(c$��0bA���c0c���F$bB)1#��1 ăH#H1H�#0A�A�� � ��`�b	# � � ȃb@A��10A�0A���1 � �0A X��� �1 �  ��D� ��  �$H���dAb
`�����(���`�`�E(�dA�$AE$�#��0F	 ��$dF��$�"2"0FȌ�A� #"0FDDdF#H P�
�2#dA�#DdI�0FȌ`�� $�""0F��ȌI`���"�`���2 �F	 ��0#�$#dFD`�`�#dI#H Ȍ�2#`�#"0D`��Ȓ"2#`��2#�"�Ȍ�"0I��Q���@�F""0F�0F	 �"1#dF�$#@FDDdF�$�"0D�Ȉ��#(dF�$�$ ��0DIDH��0FDA�#�H#dD�2"�#�`��H����@��VDH	��H!`�@��H	1BЩ��X A`,*�`��� �X7 J"@�(X�Ab��$*XAb)��
=���Tu3^�]=�%	���p��("�*�!
 �0���RW�'����u��u�_w������m?�y��{��|�������ν:�}c`�$3�=�z��$����|�GG���8�Hz��>\��u��O����aO@�)�|9��'g���W��������J�pr����@�~� *�)�����'�,�����|�B�!�ġJ_��Q���tӇ��?܇�4|�d>��t~�T	�������HJ���Y�o僇��J�������?��q));N�V"�4T|u����	�䟗�j��>��S�,�C���ˏ��W�N:)��#- {�
b" ���(���D�"���?�B6��z��%]7�}'ۃa�t���z��x(@bBI"��@��" @D M R$ P  _��!���G�����������|���H0<hO�S�`@�~�d?�_���6��	 *�R}������n�p�����>o��_���}A�a2WH?D����I�>a��2�&Gb@���{_���^��>����6~#�?H��~��_��,�����>g8l����W�>� !�|O�U���b�����`}�*���P��zd�p�Ui %��� Q˕�d���$��0�K{��a�����e�CXID?�)�=�Н]ꏼ�����k�� �E�O�=
*�R���$'�������r߼U�����R}��}�������s��Ӈ�?e'�l����O��!�i=��������DO�Q����G�����0����)�=B��`A�_�U`�Ld>��g�0�C�>�bz����>�zN���ڻIA�>�|F�`�L,�hg���_L����|��� �/�!��D���k�p�A��;�~�Ui��{��>��j�����~���1���p����6��	�I�����=�*P:�'��?
q���=���EDi�~ !������:OY�Ҋ���&9K��_����ަ�O���!��i_2�*�- 1�D�������"�(H>J�r�