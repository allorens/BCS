BZh91AY&SY�*Y��_�@qc���"� ����b?�P � �A@H�
� �
 @� (R�� (� U P� (�	
�� �UB�����
�AJ��REU
(�� H�B�EB�QJ!% ��
��"T��T���UTP�EB*�A*EIQB�PUT)IE**��U�
"�����ET*�D$�H@IAB)%$$�UUUR�J%L�P(PJ�C�  ���҈� ���`����eL�(�lP4A)��m�m��mklEU���j���j��UV��k/]�TP��T�
*J�UW�  �� �PI�0�A@Q�(��c@ ƌ �0�  �� -&  0l  [<�
B�R$I)%*P�<   ����@3�  p�� .�������p ���� M��  j�{��z3'8 (sE�@ =*�P�QE�(G�  ��� z �G8  up  Ԯ��t,�� �Wp�t4e]à �0��3H�4 �� �T��B���RP!<  �x  f� Z�h� �  ����`ʣ@i�eY@i@6�h��`  � 
^�UR�TU* EUx <�tM# 4����L �`�m� & mm�` �	�� ,S�kA�K @�܀R�D�
T��^ T�( # � �L  �` �ZF 4(,� �,�h�
�ѠPb0 
�uT���"����R�D� �T��̬ hk0�h l� �` ��@+` � C@4�@�A@$���*�TDEx 2�(�� 6  Z� �F  Z �L
�H� +2�l�`@�*URRIJ�*$N  QT�1@ Ռ C
�����`�
aX�6&  mU�
<  
� j`�J���  M10 O�aJJT��12` #L�0F�昘 L L ` &O��P�      H!#*~D���M&���j�'��$�JQ�II�     8���ϵ-ۮi�S����ΫL��8
N��զ1��u]9�"�h0d��T�uª�+�@aUNJ�{�:��QUTW�0	�����U>B����@�5UV�{��M��%j������� �<XD�`���L0��6�����ek�6���V�*��[�ս�|���5or��m��V�-��k^�k��vm�k^��V�e^�k�ּ�kܶ��k�-�sL��5�r��5�sZ�-�sV�6׹�{�׹����k�ֽ�׹�{�׹Z�-�r��5��^��V��kܶ��[ܶ��[�����e{��sU�m^�k�5^��ڽͫ�ڽ�k���e^�ܭ{�W���ͫܵ{�^���j��W���-�ͷ�kV�d2� �� 4aRXVXE���m[�k[ܵ���m[ܫV�6�o��k{�moskj���ܶսͶ��-���U��[Z��[[�ڭ��[[�5[^�֙���-Z�嶭�Uk{�V��V��5���kU{�km�Vվ���U��+V��Z���kor���5���km��Z���m~smW��[{����j��͵��+[orֵ{�km�V�^�o��Z�-m��[j�ͭ�{�W�m~2��6�r����׹Z�6�sj�6�r��j����m^���vW��{�W�Z�6���{������k�-^��k�ֽ�׹m{���V�6���{���[�
�0�V6`Sf�?$�5�3F)�����?�6��w�v7f�9ZEly���+�
�"�
�d̠�V7�����l���f��D���n�śk�Y0n]�m�P��� ��m^AV��L��k�4a 
�0|ʼԢZ̹��tec�A�p;�w5�v�L:Yɔ>5�M���c:�:��	)�ۛ+] stn d*ڣ�B��F�Vۗe�W.�Ɗ�O%WEj�lf�M�/2�)���,��bWb��f�sW���\s��u�A��b��U{K>�����om��+m]'O����4*�n=��[�MU��fU�'eم�n���#HK�r�ǔ[�)��*����Y���2f�.ɡ�4\��ކ�e��qAm�@����:+P�@�O$MVh�kO>�c��eZ	���$��HT����7E�bGm���(����d��㊐`�h�3ER@�z&D�\sf��*[`hj�#(n�OI�"�����Dq�B�ĉ^dr���{����V쬠��a�W7~Q�;on�Ĉ���{�l��u�ۉ�%�t�Zs2�w^�u���(�;��,�PX�,F�Jf���Cr1� 1V���p^:"��X7�tRj���{uj%�;1c�pՋf2�3U�CmŖ	�$�˴��%4���H��'k�k��x�]i]g.��4�2��yu#��e;�� ����_%�Z�IX����Y�	�P
���x�X��"r��k�������cʖ��[�o]m0f^k�w�ܛ�����2��f���t46���7"��5�AYUl���P�Y_:�˱.G�W@u��u�:{:������B-[<��|�l#F,J���Hă%�W�=��{��v�#]4�f�V�HD���g���̓q ���,jGv��)!9t,�dEnRTf��n���{VԓS�쪝6��\8SR�e^9l[��b�Go�
J�);�5�H)��DƝm%��ɭR�(@�ā���v];�u�A��������Fy��T�Y��YL^E���Ic��:�8�*�:Ƶ�G� �����凁�Kf���LJ���#4ɤ�ݓ1�w�c	�;X��G1��v`ה�mqHfue�l��^ЫC�<��q�e�!%̣v~��s]$�Nԋi�a��k��2�*�p=[�N���Z��o*-���B�zk�L�RPJWn�Ԭ1�t�ּԫP�(�S쵙����P�y���\�/of��$�{t
�GN�Xaưݰ�4��t�fV��7t����TkvHd��1Z0h�ARͷ�F�^\��6H�Ff�Kh5�,\Zw��M�vݜ�KdXN�;�����nH��t��@�)��TiJSv*�k4`vw5A�Sq�.B��#(��1 ��x�ѳ��oU��&Z�ٮX�W����0	ö�f=�F�c���.�COpx(Վ��qC�n���b^jD넭�n�\;���۹�<�P�"��Hf#W�-em�{�*VNγ�۽�+8�V�2��N��7�%3-h��n*��f��ݥP�Sal:���㣁�5��:n��M�q;�{@�	SS,��m�D�̫Ԩ���)ӳ[kLͼHH�fVj�M]^�l�X��;`�]���RVtT�d�u-5��%�������7ݚ+I�yoK��Û���[J��h�)��|�܀orf�ooU��hܬi!ƴ��i���D�w̋��kZݦ����5�����7�Y�,Q�5� ��C�ZV�gtd��U.bbҠp�N�q�1��+5o���)@oo6���p���ġx��Faej�2�Y��xhX3� J�,i�y�$$T�^��N�;�����\�1K�X�cˤ��hEouj�-Rd�B��ַf��^�±�Me��m�y	w���t�Ņh�z����\���c�M����zlͭ�6��D4(�ܣÑ1v�Y#8C���lc1�ݗ�6�w�Ĭ՛��E{3dR��{����V`wU�%g�yC�լlr�Š��V�J����[Ƭ�h����������7�]��,�ۖ��sE���Ś{�"o/0D���DVCm]'b��x�	��ۙv�T��e�y�F�JqT����u�-T�(n�f��_<6IY���� ��r^P���n�SQ(c%ŗx�V�������,�e6]�w����{i���g"�5�M�"�o|;�!���r����2b�3��I���"�K��li�B��v�hm䵵���K�N=A�s1=��QT�H����N��:��S�,GQ���^�2艨�Ұ�ͨ��V�`�7Xɷ�`�Gii(�m)&�zu`j���!�V�ݤۯw������8y��n�yZS�:sC55ǔ3�J�d�&2(�M*�ցZ��cj��N���.���[�6��t��m��ZKM�Й��Vi��$�!����=W���'RňTj�k]�y�FX�̠´v;�aoD�8u�V�D�e�&ܸ������Ml��O��E��@_]#Þ<Z�N�J��|Ep�|^���z�>Y���E�k^B�@�stV��;N�{H͆2R�+Zn]���K[��hW���C��l���6�2��q��hRJ��	X/R�gm`N�R�Uq(D1�f�
�x"ǩ۰�a��fn�m)��f��� <��)�y�ia�{lU�SUau�C�d*�A
�^m�fF&R��ʘ�n�dZ�q��(n"5]	�
�����]��nT����3�j�6��b1�� Y�8G��̩/#�+/U�KƝ$�B�L�Mz��?�_j\��]YJ�X��\x���U��6
А�X
�	�n��֕��ea�O)�wH�Vh�;-�]պ"���8Է[Q}v��R�Z�+)�2���y�9ktꭚ2�>f��oKw�� �c�ެ�m�5����[HY����u-�/�+���U;�Aہ\*$�ZT5��P�c	<�m�Z�A<C�@�������a;�Z�6��H�{A����)YU�P�j����"Хʭc���m���u�-�hZ���"W���%�Lꦵ�;{��SHk�M,/
�U�PJU�(�d�1���:i���I����g�-���w��[�]�d+���,���F����@Y�E�sv���Y"���ؽJ���h5�*���:"���k-{�әB����c(�U�r�)U�z��5�s)��Xs�˖�R��z^f�WHY��� ���E��R���U-�������6��[}�e��v�0J�^3/M]͂�]^eѼbL�c�d�Wٻ�b��B)t�#-��h�n^V�J�fm��`xp��4�h�yO콈�aэ�Rz�tT�x�;+�±Y��껬��U��5JU4Ba��(K�A`�x��#���e�F��ڴ +2`˔��^����v��TV����d���3둚��"���ya�.�t���h��۽!�*ɖ�t��-��+�tSp�o1�y�C�-4"b�$���ڤշM���;em�ɭͤ�U��rP,�;�XvV��+P�"�nř�b%�CY��/H�E>�sq'�Si�T�ɪV�.����n��i�/����ɭ�������A)��S�۷��v�ոlP˕�([�гZti9Q�5�]���P�*Ui����[0Ƃi���YyZ"i���� �e�M�0�R��f�i��.��
�,�co�[X���.�C=ܱ=��4��7��%���[�Rz6�\0Yf#6���u%�����R�0��ǆ���+�	�MƵh�VY�ZM^_�R�n�]׏S�BK6]�R�݌�[d��ݷt���]Z��5�ЅAJ��7/4S�2�8�ܠ�r+d�>)L��:mYu�z�R|��4��^��_'ie�^U��(�ɓ0�ʸ�1n�e�ܗ��e���駚9᫲2�&����ȳA��ۋ3� fk�լb�F�R ���^�˦f�)+ݳ���jimm:��[u6�8�T9�l�GdY�Q��d�1���N۔�!��8+,j$��B٩j:*�5$�&`HrT�7�hF�bZ� �/6��c��J���Ҙm����흺3Z��;��D�Q,B#LfV�S�2W�F�3kk���FL��Χ�G@��Z��Ŗ�z�1h�,�dVM���*@�6ƒ��	�ʮ�vz.�RYz�'&��u��,���I&��
}���U;��(�Z/�J���ʳ Y�Vދ�dF�bf����M��DHY�J�ٕ�BKr�߳j�-�d1��mA�(�ZCY���6��+��o&|�]�DͱN��m�d�Wx��z�-��D�d�'eN��a�Q���L�(G�1�!�Q�zh��7ِp 1wVՀ��蒶��!t�b�0�O[�˸��1L�\�	&�$�@i����Yν�_�Z�etވ�]>�0���ڶ�˦n�M�N���+]�/&�Ǆm���R.+{�ƕq���2��R�3J�L�2�2+��{�%#����ܻ)�F�+<�o)h�]k.hǖ��� 8�%E�ACGۚO٠,_v��kT�J8�Ze��0��-2rd4rۙ��MtU�Un�\(�w>2�Vm���U��f�;�V�Wf��i��y�ubf�����qЕn�5YB��IJ���.��S[c)�Y����w��¦�bѦ�f'�]�pI�cjj�[
���ô�(巶*8�g�����i\x6���S.��$��l-|�b���� ���Әi�l]n˼&&Am���Yv���&���2˳��ú*:G�Q���R◉
��"�˽��૽�]��rìӗz/Am506�'�v�*��q�P�Ӱ��\`ѫV7M�WYv^S�kM<ͽbn��r�-'z��6��0f�YX,�5ԫycF��A��sv��jl�L��3�\�w~@=��P��[��F�r���R<�	v�^�A�w�����h�[��{Qf%U�B��2.�	�A�$���0�0![$��{@i��cFX���u�)���8��MwY5V@�cY��M�޺Q!n�u�c�����E���li�SY���Ç[d�FH�'�XJmSc�uù���;�z�SV9]�*��iP�b3hVH���su�Ex�#�`�3%�>WR�h$�����A޵�3a՞�`Қ7EX�����;H6W��1!����v�<ݒȭ2]<�4/p�/��J{YZ���\L0�veir�P5���c�@�Ti��U��rćWwm�VlT�owMYS,�3f�GV˦���@�x�L�9����A��i,w/-i�M�ha��։���\�3�ͳkףmf:�2�'�<wytLl3B�@MZ-�:�P��1��n��ݴ�Rj�H�@<�P���F+��e٬�J2M����$�
,ͳ��a�R�D[�68�D��{0���s�,ݺG]p\C�-0Uj��,����u�7�m$�����@�Ң�%f��? j���n�p�7,��;4���aX�s&�V�#��d��Z�Ys��e73i��:.ⳛ�%F��FČ�p�w+.뷉u������wo�T���pLj���;�NX���U�9dn��)5��>9��K(����G�ۡ���JSFK�reB�It�:K 'ƴ�{f�klc֗��{ƈ�Qd��T/2�
����wMt��^ZMwk�v�?��f�{dgeӫz�P�{l6���fX�.�[f�P(��[��qG(�sY"������n�ɷx��z�3B�xâ��E��S+6�M:�Ⱥr��C�F'^#kl�$��E[�Aj�8�KW��7n��5��7[(�'4!D��vca�
�]صLɭ^Wf[�ywv�"�(�&��v�嵊�x �i%c sn�n��u���mT�$Mt]Ś�-�� �  �n���%�	k�ܭ�w)ּ�)M�w54w,�[U�;5;N����+se����[�VR�IAQK�k5���o-��{����]�]c�wF������RYM���rɡ%4j�P�f�D��nU&Ve��yr��/� �Jâ��`�!ir���g6�5kϻ ��� �$gu6���SX$eL��lF����{NS�K��ifm9���j�Ǵ��-a�hXÝ�k$���Un�H)fj�r�"@J�V=�%O2yW`����Փ2ڙG+6�^�N����B]�6]X1�Y�#|5M5���[Ж-�WW�&;8`0n�0�p�N�܃vCythͩ�^X�Y��&5��,��,�DJW������r�	�c.��+��F*0� �n�����D��lw��v�io;���e"{lVo �{]�Lf�u���� �,$J�j��CV],���m] �l�/��覭�Z�c��xDŊ��P��6vm��vK�uZu�m�k��:�v�!$o�m�T�C�Z�4h�XF�*���������.	�^YEjܭ��3��n��٬�m����l�����kE�ƚw[�h�
�T�kF<Z�mb�AkiG*���	E�7q�J9�maWn��n�L�M����v�2wR�����{& �r�����b*��Qѻ��h�z��H�����/���-mi*Rj���ÄMY�0.�m�W��b��������b���]���6)ܺ�3C�,f�{����� P=��b�D��T���?86�\��^Wkh#N��@ӽb��=M"��q-s/=�Ed({U�ӌ�ն�zS;�\��Լ������<�������i�8IӰ�]h��Q��&�s3p+v{\�aP���oFr:p��r�;6{n\/Y�W���i+�e�(]��`�V4�=�PY؟Y;��%#	6I7ǯp�ͮ+a�r�G(i7�(V��m���N����J�B(�o�ͫ��;y�9�{h`C{oK��e��ڎ�k���p�t1֐��C�R�jJŗ��j���M"S;CS�=�(8*�e�u�d���7G�g �k�:,E�JD�1K�:��O���S{����z��-r�'������{�9�t⻲so[t���{"-�N�#�����q�W�Wd檆��)+�<�+�[�dޭ��91�W*�Y;j��LI+�
�Zi��	�^��S��f 8C{��'
7�#��ʔ��T&�t�����mL'4�6	bt4%е8*�kX�P�;ƖF���g��
d�]�Ŏ�ڼ͆��L��&X��A(Jq�k�-�40�%Y�×Np�4ME%�2���yV���js��Z2�=��9�ɶjHg�6�P��V��v�w.�e��!᝷���Y��d����x�s�0ly�k��l��7�s��&�E�̉�H���.���Ĥ���e�8	익�!��NV
��������Vg�R�����s����(-(jΤz��"j:^Lu=�I���;xT4qu�X��rn]�7��X���e�GΜ��jS���v��iĊ�P�kZʃe�ʻ`�(����chb[G���`8M��v�P�5̕�e��2	V����@]�0��5z�����4#���bs�5n+��w���|��+Y��.�QS�-��¹��n^Q䂄�����3gy>X�5�ə�JNu�n�ŋI>BZɔ�h��V��%b��]��ū2��zt&��t6�=�R�=}�[D�jb�t��ˠ����e�c�}��3��3
��Z��;��v��d��1#=��Ό���x���S,Q�B8�U`�9�6��ݪ 9G(�Y/w�74�5�������t���>�*�jc�i��]7:ulf��3�`�TB��upZ��*W��6�7�'E� {#�#�ثOx{2эu-�N�'z]ݫ��kV�iΨѭ�����»
�0��P����c
���|]qV�u��ycpTqiM̡���l��h2lч0H���*�E�Y���E�:�=�K~.�K�%����+&�+s�5���ۥb���U��h���y
]�����cY�|�I�nsmv���ZB��v�K�|��*�V)$kT�8�����'���2�PJ�ם3So������j�E�[��r��Z���VPۺgD�v����n��:���hUJ��Ξk}�����5eK}m�]��(���(n�p)2�}+b���Xk�کk*ۛM��g�[X�6�4_�3���\�:k�#l�P�]�m�w�w[p�d4Ղ���!��A9��pn#�˴�ڕw��(�H\Xpd��m-EU�+T��T-P]\�j-��P�[.qz��������؄�We�ϣ.��r�)�X�����}.��|ȭ�G�~E6��ɽ��%���a� �Ҩ�,Wu�ػ�Y�z�h5IW[r�u��5���/k7~_o{yZ'���F���%�ݓW�.�]���1���+�veG�}ط�⧠*s{v��Q��7'v�U��X���Qwk�i�;�η#��-�{��iY2a$�q0G͉��ET��&����M�2�u�i�fM�!蛍vb����g�nG�]��ʇL�:�$L
�N�wl�{�V;�::0�J)��H֢�%��EQ��U��td�:lc���\Հ��mg�8���/�jU�X��+�rV�ܰ��7Y���;W���}�f��
�/qæ�Y�ty��IĪ�h�V3 �>��S/O�叜���u+GiC�8��1SQֹ���*U����zi��Q�Rw2mӤ��i��������0�x�v#&�ZR9n<�h���R�ӣt%�J��vE��os�˩�|��r�u�b���<!���lO.��bX2�����(���@��u�W�V�uʹr�u��H+	�D���Wn�bbG$�k�� J�
U��Mt�;-�Q����z��SrV����M�~��l���]��V��[�v7[PYyM�G Po����3�h,���mp(v����is�:�h]�7�at����u7:�E+��im�%�#햸iV�+:��+G%�rGV�tAɷF�$P���b�<��.mӧ�+�{t�wSM�>ɬMtJ�X�9�#�d�t8;��'��nK$�{�o�����aX�v���RN�zs`5�.��|ҝ� ���!� �����j.-ٳ*ޜ�:��.�hF��ę .λY��,pPW���K��:�L|��j��OPn�PO���9&���8*\��W�o���NV���Q©��tȨ�GS7:�e��ԩ�APqSc#`gV�K��L9F�wNv�"kq��ߙuBN_�e��e�u���۰�*���#�2ɥJ^pV]J�K�2	8�����+�t5��_�E�c5�E$�t���sMwW6p��57����}���,g7���J��u���J[�^f�
x�{�j�Ƃ�E�h���u��Sl3��iu�k%��/7�=R�d��]�}sǍv�xi�}�La��;�;�Х�X�]>�6��a[+����ױ�ss칽�vV�o+��aa-U�.U�y��x���O��-��FQ��-���s��L�z�F�X�R��>��)eI�}b��htA]Om������i��캗�f�6gJY��)�>��·*X��{:���a]4��uԸ��b���qj|)>.����.��"mt=�䒷�ӣ��: "��ŕ�����a�yvU��f0	M�t%��Vd�n-�u�h���w�#�I7ݴ����M�r���t~c��I�d��ͬY�]$�a���-��5aV��RL2��Q��ĝ�n�s8B&i.��}��!cVQ�w�etܧ�ް��*m��
|��J��X��lM�f���G:�]��:�ٰ�6i�Q>�"��"��o#���9wzK���q�n�M��a�4L����:f�G��Yqt�zv�u��G-8�����K��bw�lN�M=�4��]j�՘�,�Tl�y�[��:������xTu��y3���@�A>�[C\�-(�LOh�/k�=�kK������ +6��J�21zLۢ �he8]��][dU�n;�̢E[���50�IF�2v�h�`�d��.quj���Lpۍu�ه���[̝[OX589��<R�Ʋ����c��D�u�N�%#��ѽ?^�Ƭ2e��ܼ�� ���އw ���;��J��8	u�|�&�O���V��6�c[/kc*�j�J�4����P�v���7 ٲ�W-2����sq�+,ԩO-��9�i���圳{�%��Ǆ9��l�4��	�F�:��Q �<�#c�.�Et^�����7P�[��\�T<wl�66���r@Z=]qf�N��WEջxĚ=S�gaX���5;Z�@���t��,�&r��]\⛏�DD�<Խ;�wI�p�F��qc�ծ;�.�Ř�]=В5v{�6]���e�ݢ+1sFe�G����R��[��@I� �#QoYذKqB:��Z����H�]+�ѳ-��	t��ⶱ�f��-��]��-���k3�pN��kW^-L�?3�>��%����h�b�ܲcWO�eO�\X.۲��.�������wK����cz�/���
���8GSuC� �7t����O���������;����,�9�F��ޮ|��S5p������¦�c���l�+^-���lt�����>��գ1���Y��C�MӋH�sn<��֡��#4�ܳ�iU���(#�.�v��T�4d�u�.�`��sh�ǌ Jw�_<�)R�*5\�u��5�*[��A0�Kc�2�/n޶�\-���p,paI��}�y{u(�f	��*��9�R۬�;tث6,��|������S/q^qܛYC�4#��y�ᑆ�P���İ��>(�Z/H�[:���w�G�^�Kj��R�`{U#˛�)X*�wo��dvpTL3�R��-�&a��\��y�`�;���=0��	���}g�ud�ד���#��c�����P�^���53� ���u}ӫ*m��&Ʀ�;9q�D��uqZ�nb�
�Z�i���8�{NX�ye�*6}��	pR��7����D�m�T)�� u�1�P���o�
Y���������o������ڿXG3��YE��Ex��(��2�,�I��|^���w��8����ea�R�W����-%��K������"�K��M��b���������],r�����I��x(�
W��B��	�,�����f�No���NJ��W;��/��p򑾠��Gk7ԅw^� j4�s*h!���� ����Sx�� ��p5nq�kL�.�z����&�Y���.w�H֌-�)wm��0��\�i;8�iZTOu�ky�d��i=؇*ɔ��:��R"c砷i����Ԇm��wyG ����[#�To�b�J�i�V�=�;P�/;z��:�����m\��e�N�2fN�vjĵg[&Vt��W�o:w{��� y,"�ך�@�R�+YkEu��rMۥY�u�32 g=�\�%�r��gH4��1��S3]�zK�yi]]���͑��{�-�N�s���a�8�:M)�诱��r�sn��޹)]6�V����]1rè�õ�{�i�%���m'G��'�s.w,~ujJ�=�%�(v����h�W.�kZ�ɋ5��v�x�fWf>��k��� K(���V��J�FT�9o�Ļ/���V�MG�%elO{o���5_���c��2&^��S���K��j��<�"�S����Ma}����*{¥�����'syl`mɁR��(M��P�]���dg�n^X1����gl�����\-
������ܶs�M�W2n-��R���"��/v��0��Kr�����i�b䢽D��mi�9���]XƂrVPfVR�i�4��b�:��j��\��>5\�p����3*���ѻ��r��q�6�'�@����f�g��_g*-j�~�����r� �,T�=�Xp��$O��엶	8C*������ʶSt-壹�r�����v�Y��U�Շ�D�t�T!�cu9��ty����|�T��L�"ݱ�@#S��yW	E��b�����N�6��CB�s;^�FW�cѨ0��1�f��9�ة�N����*d������
����褳���V���������S,�@�F%�39ĶgZfP�/�oSYt7-d��3)*���5�E�f��f���{J��y��c˛n�WB�v���&���ڜO�;�`f�����;2.N���-Ͷ���7m�w+�nZ�9$�����v�������VN]�z����Oӷ����5�<��B�"u�.�H^�K�oc���&Fs˨��;����nk��&|�v���Q���a����m2:UKn|�+���RS	���m�n�ک����-2[ݼ�];�L֓.P�|�yU��mp��<��cnĠ��F�����MdJ��͜N"jƳR�Ф�ú_E;z�R��7@�G)0�fWO�����kz���m�̻R�a}/K�fK�4�΍ff�
t��:mne��`di=�y�vƾ�-@�s����L�7�Jܬ�q����78��h�C�1����2ū���z��]����k_��rrw��ئ�O�1I�\���wVk#�X�{!��r��]��3n��-���ΝFF+��6�Do�G�6���怗Q�kt��(X�@	��ga����㋧NΦ��*�QjC�>�6�XYm�8Nu�]��wz�<�M,�pM��m�=kGgs]���:HP�78��ы.�*�ց<h\�����cw�qyɫ�2sA6���r-�^2��<�j�[jpOm
�P^��:��w{���M��9�y�-�:����|���"�G\�`���)��Д|*O��4
�7S{,�s�}Ɓ'4��'
B��F�����TY���ZS�¡�0nB�9�@���z�8���4P�����+�|6<}e�r42�}�^����13YH�2`T�u���rfW��,�E�ۼ�*�B��XI7Cc6��Y��՞�:���}4j��f�ɢ�k�X�����u�]:�M>�a�<6�t^ܤ7�ﺖ��֕K*�~D���E31���i�秩qLۛ,�V�5�SJω�����y���xt(-LW\��b�V֞��Eu�S^ʘ���Rdw`���r�fl�{۝�Tk�ia9�(�������k�:�I����p��[s�b�IA%v�Yp��Q�o��`Йޡeb�jۮ�}gT�J��7Bi�6����]�NK�-Z��/e�=k���w�(�C�xK�����ٕ�p�wn�w���}Qk�7���ةF�k�(�w�fQ�{dU��Z$������'�:w��_W6��u����^T|s�,�����2�Zq���k��O�E����G,�ז��n
8f�j�a��p�k4�3@*�O�pJ��tu�����mҵ��=�l	.�tҳׇ)��]Y�vT��Lh�+�홒jjK}�Nb����j��,و��>�#���Ɣ�Z��=R�/c�; ŵ���jy.v�XU
�����e+�G+V�F�OV&��ûd�5�ԧ5��WR(��0��N�I�6��o(������I�nα���ۄL�F�.\�;���4���۟u��4�ҥ�5�6��aK.��U��f��jq��2�����}�����;s4�*INIҤj@1l1�Ҥ�Z��ZۇS��8�:��B�Ɇ�RN?W�.v`��HfԡY.�X�B��|p7�S6�΂��Ղ��}f�WB�al1�!F�ȚB�8�S*���
�������M�����]D�_�1TF�T�\.��"�l�SM8j���*�Zc_/�Om��G
�j���K�(a�kZb)a-���4�� T^|����n;��o�?A���9"�����z/��S�>�Z
�iK��?�2?��B+�<��皇�#J�Y�:fWY5%�ٺ��B�`�F��@W>�&f.O����߰�g�㬬�B��t �<U�D}�2��I��Pts� �q<#�|,�Y�2�YƏuKp7�a3�<�h�����YQ#2n
34%|����yt��lV�(���^���wu�jd�Bq����:0{�W�I�*i�ҙG]շ���;A�X'����&�t�[�j��j|�uouKbK�c(V���YW�9jE��뵁�̓�W[�Ю�Ս�t+!� кQd�1���ئA�ΜֻV�X��2�aR�qO�c�p�[x���8n,t����4�p���F�-|ȸr�-PT�*9W��_.-�@D�S��#���w�uqoS�sq���Ct�gK�eӀ��_p�!��>��.����Ӛx�4�Q��j��M�[ڍ\t/�>Z�$����v�S���BxT
w.���Z�K�*�o9f��&+�ij5�JK�ƈ0�����݌�)��5ws�&2X����e&/tI-�z=W|�ɝX�V! u7[�0�̤�]�G�ҥ:�M��}p�7s%ʌ���aTg��Ӻ�p����o.�L����N73))�;#�N��8�ܰ�7@�/8�ʶ��nK�G�
�2�@���]�m��`9�#�&�&^mĬ_Xxn�VS�s�͍t�(9YX�YI	���yخPO\��^V�LwkŻ�vlcT	�d1�t�x���xj�W'85*�W�]�l�[��rr��?c�����R���C�"]]��[yt�
��;�5��5�bd�
1�e[��>*�M�����!�O���kbc�QE�����ν�5]�ͱYx��ċ��K�U\u�D7:�h�&���7�/3	L�w�H�je�났��02;&��ݺUΏ	|�P�;Yލ��K=Y���Y�]�`}������O%���=���=�(��Հ�|��HJ;2�G��-���!�84&���;�8��zi�6u�Zy���!'ٜ��T�Gm�Ē�xU��Pv{	ZB��Lx[t����.�8mY�S�>����t6pڽ�B�2�7�WT��_�#��3u۸�Ӣ���E�}��*E/�BkMiz�Û��n�wSc+�z�iD*xe:"�Gcvd���Y�AT��Ǩ�n��WיN�P#�HZ�Dh7Z"�s��&٪�j��^Зc���ۖoR��ك*�um�nE�h�^dD��C�T�\5�n�����ڨ1W�D��}����Q����2�,wtR�/d���e�����<�W[���NG�<�0l��܆�m�9n��N��!Zƭ˺���j�]�q>�J��piy�����CI⛰�]��.<�ה�Q����쀀3�\&�6mwr���l��vo^��,)6Sn�W�﫰���q�{N�*�z��Ukh=����i����K�lfU�T-�;�*�jbZ6�L'�ٲ��9V����U�o����8x�Y4+R7ى�h��2R��0�*�{^5�zp�����37^�55�t7�5]Ko�䫫Jq�Y=����Ɲ���3�4��g�t95�^� e�vwE�&��c����(ʺ|y'J3�Q<��ff.ӵ�حG�u�8��ɛ4;Y)�B(��d�[2)�	hh�#���)�xɺ��i�W� ;�:O	p�S]���r�q�l>��t`�,.�2�o¥κ9�M��g3���=���ܩʰ�#�*kV�*�R��[�Ѣ�Ԭ��o��t���k���|��E��V,�r��Ѓ�	Y��7���@n6����z){�M�S��V�D�#VH u:
4��[��|¼�6���Pm� 7%ʊ��O*�Ռa�� ��Me@����b���X�H�7!+�g�Qu�m���n�%�b�T��]Ӓ��/�����=k官�м�� �������*�gr]��T�ڸ�i�r[e)�l��I�{:^pz<I�u\n;�[�v��ɲVeI�%�k:��|ޓ8�+v�)�'�:�a�76�A �-�]]�hBޢL�Yp7�w��F�Q]Zл���K�}���&.�ۙRd%I�N8r0k�5Q����Q��}�O��=�B��� ��ؑ�y�Շx�(_����Aj!�J}A9���d۫U�(T�X��OE\�0Jd�j��A6��)����ꬋq�ުG��u2�����0��D�S�h�{C�ֵ�e�O��i`[{u��2��vb2T��jc7:^�ʛoCD=*�����_S{�R��C	Gr�Ҳ��b�*����tBB]
�΀���2��7��?�Y9R�����.��p��V)������S�[�40�["�R�j��m6����jurD� Vum�+jp�(Ч�u� U�B6.G���%\�ĺCy0�Ǎ�JX���3Z=F<�q]�UbcYW� �a&W>�)�ɕ+o�.�ԡ8����>�Zy��c�Y3M���d��7/.������ylC;�Α���NۡZo=�#Y�e���g��&	�d�3�T�o��yV�W��F�l̝n
9O&.Y]�}u�z�um=q+��z��b�n4�奈Tts���� ����qBo�ih�\{�n�{�Ew��]��Q*����	��ɮ�.#�5:��Sk-��﹧D�'��AvaM.�n_mt�en���g�+l��ةl�lzT���A]_[�ȅGk<u����-�y��t�`�d�"�u�&���	�en>ڻ��-٩�%ߍ��z��\�V����Ao�H�9{4�󈰸�]6�E�L�J���f�,쌣O�j�2�^+	A������{���S��	N8���\yt���j�if��dQ��	�W�^S%X�jU�p��q�̤��ے��s��B�&�cFᗔ�6�\�v^��ϻO>t�'���J�4�ue��ѫ��5��K�o��/Bk(���n묗3�����<�9�A� �Y{e�&���\P���o�GyŪ�r��Xn�{R�p`��Νu6jqsՃ
�o�:���WH��7�;L�i�rH5}���FY�"��7��H6�ն�0���Ύ������f�e���^˳G�ͱ݌��u�j�bѮ"��Xi�@u�c=�9��Vo>PB�Wh�|�h8q}f�Y�)]�(^1�(�}N���y-)�>���aszgG��H���D�b�4[�k���� v-iY�aj/jڗ�U��r��e��v6�jY�f��*�rK�Mpx��h�����ׂ����Ttq��E�[��P�G+X\��Q�&���. ��	g˲>�գ�fȹmmt��L�y;�oJ���}�z	�i�J��,�)�q�R[8A�q��O��]�
S��2"5ش�r���r��y�F�'�2��fm�6uY:����!�ǻ�̬��x�:��|�s���@D���X��~���:pO90�Q��i��G��}ib�����8u:	3�gQ�q����P3b[y�r�}R��Y<�5�t.���t�X�a�
`�1���;coH7] �t�T�٤Z�	W����9�^�Ts/�i�z� m���(+6�W���a�n��m��*<p�,�h��!0mYx;��=�R��P���r�h���P-"Ѿ���ut��vH3���Lk��	��wYAг���mGl�Z�mb�sn�Z�Tܷ�s��{�8�|��Z��~�e]-�!ba7%$�"����/�ѽ&�D-�o(�**�֚HKO�hn͝t���f��l�I��ۣ���7Ś��+N&u�ӯ���ʴ���n�.�q[a�,mG���w& ��k�!�wK��!�Y�Q5�T�u4�
B��S=5��u0o�]9���Ǵ������O���.�Օ�R�yx���mi+�*��)��.�jU��nql<O*"�yqmGh�$�l���|l�WL!mֽ�X���dV{�Z<n�Z�ER.����p���������z�D����&]Iٽ�oW�8������D�g)S�9��<8�N�pWK�t�������lO���u)�C��Ω��5�M!��б]����V����nU�B�5��Q���	o*�ٽ��5]�@z�7VA32���i�KKxq?*�8���T�Zp%@\*�C�m�Ë�L���n�5Z�/�GC/��ub�gcYw���f>��!A�l��޺��8Գh�@}�e���� 4�ޫp۵Cq��E�:l�)��L��qiy�8����c�`Cd��Iv�k��پ�\�6uѹO%8���x�&�(T����r�{e�yu�Ԯ����KaQ��<Ѳ+*��3:^;c��i�;` oin�w\�֊B%���o3{���}����O��I�o&�wJ��l�@��tQ.>���a*4n��o!)�.�vh 6��t�m����U:0Q����g����uF�Dt�y#�pu7%�� �\Ku�M"��nΤ�>)��a�|���73wx:�\�\��z�u���-Ul�ԁ�V��n��+��)�%�.S]w�I��0KDehzE 
5�2�j��`�s�%q.��5��l��'8��)@�����su4�Ơ�;s��샹�r�]�l��<��:"s��֍��7��a��:�K�J��΍���Y\�Rf��S[l[����)`Sz�My��T+������=�k��I�͔�r��u�W7WxU��v���Oj�[����_0�L=�"X|��'{/�:���)��G4th�C����.�F��9:��E�N�Gd�֐��w���o��l7�H䳐Bx����0v�xw�6��<��9%[a��ԃ嚳5<��U���ȘsO��!�n���H\�J�+9�W\L}ُi��s|8^6�"�+40*���9���
�K9C�NP��-I�h%+�Wn_e��)7]p7�n[)��n�չX]��f��
Ŝ��h�X��b��h�"%n����Ӯ	�X������]+��[�c>,hD�ܷ)����	�z�A���$�!�����k9�ϰ`�j
��1���_]�=ǥD�f�;��u� }7x�Z�4�6fP��Lך���� ����4viͨ�ug����I��k<�Mc^�F�Z�
«)$�b�鸅$����ڝu��c8� \�xh��[[����1Cɲk#K4��XF]c���[�@��(�ɺ���9�]\U0S���FT{-#�Du�۵,Ws�kC�A<G"NR�8�a�����N���,12�A��;kǲ"�[(��u��HQ�utJִyJ�뫣� EÖ�!�� ��a͔��и�rK�:RjR�36q
��%m�,\��H�o�j�p_
��Y���t<Bg8�S�켐3Q��J�sAB�P�X��s^j�waJO���]r�AY��q�B�)]S�4_)Ջe�}њ�a�Z�-��6/x,6�ΛbA#������F�u��YgH��儚N�&ڙI�(7���޳R]]��B��n�����j���ч K)�h3 ��+�KXW�;��Ķ�w3ݧ/���b���Y�voVb�[H���;.�s rwڠb��b�Ytu��"Vˮ�*��P��Xtf�NmȨV�5����v�4.���{�e:0�+�,���f��+������/���̃�ؕ=��egc�V�N�v.�[�᩠qB�:��Xvrm۝y�dY�.�h�h�9)@1b���%�م6k��͜O�q.|�^�3<ꛌ��}Ε�kh��y9�J�N)���^i˅z�]o2qj`�ko2�A�	FU��9F4�^Ǎc�E�����n,�a[�]�3�4��6�;�"q�ܓru\w�X��>�X��iɍm�n6yu�5��0[�]2�K2�o\��3r�<e�X��ٵ{ڛ��}�`��'#WvMr(���F��Uje�EM��o���i�ͯ�m�j��s�.�� ���ҍ]oq���C�tG��&nI�=�ƨ��3���V͡���1R��S=m�mI���ٕ�7@��]��7��r����wg>��uܪ��XD �c&����3Ƒ�(sR�W��0�\�[��\�k�����#��d��{X�dr��(�u[R6~	����KU՝�tj5GF�V�m�wW;rR0��k���;VnJ�N��{_B��M��;�ofD�#����Y�U�w��q�H��_.�����*2ڃ>q�;��x
�3�-.��"�.�p�+��;|����w�Hj��-�楸�/�W
������Hb���^�5T)5ZUe�8e�[v���i֒6��e���+���j�f�E���0���6�1��!4���a��֛����ǡ�4o�d���c�ozc��,� ���^Щ�u��C��ۃ�kr�����YEa�6��`�zQX��J�K�h��i
�q���k�V�i��X���7S.C���.Y�t�XtX0���S��]V�f��4s�;L��pmdˁ�uko����4��e�è�Z��U,K�Ѯ\�A7��O����E�G�'b�[�>}�;�_rT�t*9(Žp��9P���׶�p��Z��rكyY��Q�:UI:F�Y�B!��XQP�O�l2�G{�j�v�J������a��+S}R��{ya�jP�[��8��
ˑP�p����d�ĉ%��x�w!��!��S�߮�u$���1U�%���x��WY���T��C�}�㲓F�xb�����1_'q��i�,�F2;i��Г��K��ո���ͦ�pf3�u�dӔ�FPF��F�U���R*�����M$p���sƹ�TZs���erţcr�<���T�z�K%�q��[�UҦm-縤Y��m�wT{]Eq�܎�Ժ ��Mh�q��SJ�/Y�S4�kL_�r9����؃��o�����t��s�=��W��.\�r�������C�����~���t��D��t�$��4i�i�E�U���WE+��J5�%m{���|�`߯�����}��>���;���{���i�lt���4��wS8*pI��HwJ"W��ج�q_e �T&W��q���WL"*^������d��V)�����2Ҹ��G�A�v�Ժ�����j��k�(G7OuM�e�eȺ��t���:��5v[]��EZ��V��L,ܵw��V�:v�P����.DvqS�l��M��	�lu���ժd�,iVw9u�S7h����I���qy���7��p�xl��|9��vK̔��Ou���b� ��َ�u�}c�*r�N�c��4'ֺ������	@՛ʈ�>8�&�E�Gj$T���r�:�I��;���fma�:ѹ�f��.�ӻK;��f��Z4�ڜk��q�&q9҃��u>��)�w�e�<0�9�v`l�Zv�U�q�Tx�f��˖�S@�}�G��o:�j:`T,ד����j�J�rDK���v�'}�uF�_&nn6SK���U���Y�@[`�;��kt�]��ܔ�p&a����%K�ͮ�6��&��{����y�������9�e����~13��2��o�	=��-��vEu4ͪb�0g��bi�Nf5!f��4.���s�T�׵/���ɘ��t)c�#㒇2�E�:��K��G���d�JY\�mK�l
����q8��q4h̻��H� �G4�t@�&�E�dA$~I�	QT�
��i*5@�h��m>��ɚt�J��P���X��S�(��@*���Jwr$�3I*9�9�F
#I#���>:�	4 ��F������N]L��[��A$�ȴ�2%��F���bi��rJS`��P#h	����˜��L����dGu\�рȘ��@�32(�Q���D$�0QL���$D�g7#B�A�n��d$(� H�d��*yۙ�e!&����E(�L�D�%4�� ��R�f��0�h�,�F&�����F#cb(�V5�3b���6����\�Q���1Hd�L�P����*(79"h1L�D��9�s\ы"$���w�����u���>|�3�k|P���42!|�+�)eYS$�5�μ�Mr�gv�u�x!Ϛ��oA��&9=+��f��n{`6/`�к��! *d�  ��2������䫊�woV_92��u�t���g�0z`�K��ézo�R~����.��&6F�+�I�Dɨ;uC�2A޿u�9 �ԗ�����L{�<x���(�1�5� I2�ʣ��&\�y;���[�{�,^�{�m�M���e)���K�O^�Bj�iBy��>��vb��a�[��*_�1�N�o�+=�]</��iοx�t�������9�����/�+��9n���,G�ug2���0ٝ��aי�FN�'�N�{U�4
wB��ޫ�7���T^;�ǧ:�.�W��~�!�s���̞��Ľ�®��=�&v�=����D��<s�6s��z97#N���1�� ���1��E�TE�O� �0��ː2���g�ٺތ�@�o�ʄ<��e�&׊�YBܣ��O�K�3&^9��;xH�'}��`�+N4�A֮���Uu�k�ɢE˚fo�3n�9����5pS��`vJ���+m7 �w�M�7�l�X5�$��@-�,���JH�bnd9��}�q�3ϩM�=(:��zeU�3�=(,��N��z��#m�Nw{ь�)Ưkԥ#�&g�WG�!��T�Tf}y�z�^Y���災
H��Y���X������7����_;�(�--��o���M���-z���SeV/��}��~�/����Z�hB��X��Ks�{�⭛�|:�伿>Xc��CꞮ���ҏ�����]C�qrw�����Է
��>v}z��7+˾~�{k���%�����{��-�7�k*�%������bȂDV�	�;#O�½5)��~o��g��ob�����!��e�K_�u��wMh��oX��w�-�c�[��K���xg��)й{�z�ӎ�0��w��k�M������Aё�_:	:9��g�;�;���X���8<^�x��6���#G�i��tC��짏k{�U(4)j���~�\tS���gk��t�C�J��=�J�s�%,�%@�,u��%P�Ù����Uc���f;��PEæ�t2nl�ēٔ��p���� �va���2T9��8$&��ӕ�r�eu/��s���|ޘ��/C(�'O�Ӈ�_��St��Y��L���z�r���ly�;_f7</NU_}����a�sr}�������Fxૐ_ޥ0Syu�ǯ�2+��������C�^�jrj�����N���v��b�JwU��ۥ�FM���^�{���+���P����z�����e=��1r�2��rc��t�>�=��ώI+�����$��&��ݳ�Lt�����g������*�(a�l��tT��y��%=ɇ�ay�9��S�dU�i�\}�[���T�z}9!�=J���}����=+6����>���5y��+�%+�g��n��;�E?��u�uY�'�'ʼX�y{�����rB���/m�
L���m�+�]7@�g�\X%��Q;�1��m����w���	�]�9j�G��}���s`ɮ$	��ڥ��?&m��;$��|9㶪5~h`�_n��,S=O8��;�b�@�92�����z9I:�Ԑ'��f��=���Y^�J�!���q.��šQ��*2�N��z�᠋��p����>�N�`ݙY4�"�x�QB:��eM1�3'wk�f��õ������{<�}���&�Υ�J���Y��/�Q\Tܽ�u
"�ѱ{�*�dߝ�ޮx&�4ht�A���2�6��Wm
�3y�v[���1�٠�h����	�����S�Fu�����)��[���l1=,Ge����E�~gѼ:@���_t�4��,v澛��zs_u�Ǜ���a�r��7gѲz��vΣ=�ۗ���C-*�]M�zt�����<�6���/#��s�1��N�14�Ѱ�>���&&	����Ӿ��y�7W��Q����Vj��C�k�#��\��vpث�rE�NM�1Ӕ;��&��{:���2�ĸ٬Y�(�a��M_{(����ڶ����3ޜ<����>ړ^�c��{�����kҩ����n�Ϊ�<]!�9���N�>\\+�'dS4H���=�D�_OMz�0M{d�ˮ4o��t�ゆ>41����Z��,:�n���S3�]ʙz_.ٛ��K������*8�0�
�}�֒�D+���[7A}z�D>�qJ��#z�T;�p[�/�NŮvG��I�a�9���T9���{�w��m�=����)`��LʥFgמ;��>��\zVIk;ݮ�����,�^�r�-柇�*��w���H��WCd���[�Z1�j�M�·b���9$���D��MX!��YFF�9��qc���qVUIҰ�"�|Gx!�[�ӯ����y�^�mw������Eodu��mw[ER����]ű�>U��f����/s_��I�D�s�=�e�˰�o]2%��1{�k7\��pڏ�r V��;��C�	�H^�wrgX��7}D���eY��ܜ���X��n�.D?Z8eoo��4L��:��ͮ���'��/)0�	�jz{h=z;�ڕ�J9~�**2�քd�X���}�������99�8���ζ���Pa$u��v �}���˥�3 +,�uw���;���x���+���Hg#�x!�3���(E����d���v��F1��μ�WE`tk�,�Ƥ7l� ��:^�P�.8� ��)�/d]{���t5�x�H�i�:[{+t�5d�N4�&�9!^��yz�����~���-�U�Ae
w��7�1�������r���)t�}��������w��sEg�w�;3��Ȗ/b��^�ゥФ���W��s��_�u��OI�=̹��D�B<���q�"鯽$k?�q�.\�/h��=^/�m8Ò�������R_�w�w�W{�$�uүL�Fv!�X��P6�����ti���� h$uw?v
�A�6���|����۩P"�*Y���ֽfy��Ǹ������O'�y��P2���p_�eM�}��|B�&wsO��~To�o���M�FVk1�}[T� R瞉��_��ع=�J����߽2X�P����MxD�Ȭ���H����o��c ��ޚ��-M��%�\���z�0[��Q�L�5영���^{���I����Lv��k8q�n��a�:
v8Y����%���W��)�P�\��+�������}c�reB�{��+�ٵX*V���̀��)Vf':���0f[3	�F�u���6�*V��C5L�=G�����G%���nf;�w���RQk���0z������ �z�������l[Q�=츛��G����釫��A��Ύ&K���|��m1��q�<c�߲��ٖV#&a���:o�zJ�����I�x&����<j��{!���+����dI��B��}��\���g��vT>��M��j^��<h=����'M�%q�#stW�7SVDFz2�CC��[>�ѳ{Rh���_ =GIn��[x=���[Ԏ���� M�@a}9��a_��k���L���T���~��ׯ�u���|��s�+iz��M�Uלڬz�s3�CϢ�9|����U\a�"���$�uE3�Xfg�p��Ϯ���c]�Uk�y�]����-{�.(��X��휮��� l���0�b�~��X�k�i$!�a�m���Jλ� \���[o���}Żd ��=(/��G~�7q�l�O���2�q޻'�R��/4�v�Ǩ�؍]jo&�WU��jOkUԯ�X~�Y��E����WQ�s�Y@ɽ0u2:\��\W8<rql�k�k�I��J�ʐ+rݗIo\�JN�e�1��v�`'H�pb�jR�=����1[�-�V=YG����Sܘxay�Nl��q�QWMN�]b���W���x�n{�r/�;D�T�+��Ko'^l�������;��+I˫�[+���7�>���{KE��z�n�^n>6_���e���%F�k%:��{2U�����
�'Q�c׬]j���nߢw�R�uWKo����I�\��9�d��UG�^�w�/���C�K~;ֺ����g��n���$s�H5��_׹"�@��r��I��MzN�y�=������u���c��Rr2a��6�O��<�N�h�5O���sNb�ʒ��Z��Օ(��Ap7Z8El��Gl�Kwd�u�ѵ�0�Bz��I�Z���n�DJ�8�K�����rL;��-���{�������?KyF0����ݿz���Jo��VN��W,��^)[=	��{yZ��Fu�;t��f��u���}��G�li�s4���nR�W��o������r���JW��w2��f�;�S�dU��j��!����y/G5���L�t�b�k6@Q�DL�n흒����{��N��ˆ�t/⥢�fS�/x�%�}[�y��q��<��I��H�(���ѣ�\{��dH�8�l��/g�W��N�+m��ߏ�q�;�����͟9�q���G���dz8
q�����j��%���(olZ~�B<��8���x�����4��y���=�@�t����BY��$�w��d)o_�}�z�O
J,�_�Ǵg�:����~d�|(�'��{3�_.!�gI#�=�W���&�_��g&f�����̺fv^x7����ӕgޘ3ʹ�>)`��L�Fe����i1��z�R'��$�H̽�O϶ۢx��Z����?`�τW5�&SĶi.�a1�{�:H\�/Q^�³z���xg�(�ا3�{m�NXE������}gҺ㮞���٧gï@'k��F����mǪ%�m��0�\a��ݮ��~�\'�Ci�V@t�I屳������&��o=�q�Y�u�؋�#vY�K[�R� ��wO�@r���j�b� �r�!]'�P���^3������0��;y��X��H�^��Wt�x�u6��ne$UϷ%���hq�/0>�[���\���>��l�zҋ��}�ub����pi|�l�qc���pN��˪���M�U��t4�k�	C��dʛ6pE�q��܎ˮLC4�$o��_�P�_�Fįu+*��,v�7�{<Q��QC6�1i�X�����e�.��#xw���a��ns7
�����
2Mi�����u��v�b��f�^����I�5s;�}t'O��^�wYx�9��{����~�+��x�� ���=���so��W�^���'M2�=.�߻�����K�fq ���Z$>����K����� E�w�rC0���d�ѽFܛ��g��������S�-fw��j[]�&U?���^}Ҝۣ�ߑ����<G�����J���7ޘ��j#S~�BeJ��U闈Ϊ�<���W��ϡM�ŵن�Pc'�u����d7Y5��LjQ�g�M�:vwe�.\�r痈�^���^������x�����E�,p��d�y�9t��_��Z��]n�;u�aһ�������v��	�n�-Ӣ�����.&��a�u�fT�.�n��Ӻ�-�8P١��25(+����4���^�-"�)��)Q˽hlsiB��(�N�xJ�`��^����8�7b���
1c�Y�T�2(������P�~�Q�K�	��v���%	���ym":��rwkO0��t0�Н]�!�YV���v��U��v�]�n �P�BF�F��ީ&�fc�(�/h"Xwx�����u}{���-�Q��az���D�*�8�-�J;:I�t�e�t>[d]"���5� 5'!W1�ͮ�!K��SĀA���N��M��kt����Rd�����V�߻����B�J�]a��8�q�Nt3S��ۭ��L�{c����/Y�<�9�E+zVv�oh�[�fwM�΋������]h_��-�s�K!Tz�v�v2�,������a>4��h)5��]M�\:���V��$\;�GV����Y�eNP�B��շ�.�]EU<���na2V�	�;VV@l�M޳�[��y��Ff�x-U�	K���u{Sv�T�er��wfV�y�\�Yq�.���LǧmVTu�.�����ٛ�ҋ<颹C2RV/�MT�[���Q�ﳔ�V���S&�̲�W���2��6l�2.:��ĺ��P"�c�f���R6p6�.���z��{��̠��M.F��)ɢ^V�w�u�C6��o`K���w{�F����>o�E���?Vy׸�\�D���.�
7�[�Gv�G��V�+1LC!tn+��GkWd�k��-�Hn���
�5r�[f�w=N���b(ۺm_O0���SZ(�]t,<��{j�@ot�mc��Ӊ��I��]��˽'FPL��&�a6�_\R�����J�\R<�gWC�ݏ�7��x`�7�ʾV��v�8S*f�[��L�g�K��kw�0���s�:c�9tN3@��ے��}}3Q�� �fH�h��<�����)�Oi�-�)�<xzEb�m����Y���*e�Z��YWEf�ҹ��E�T�N�U��P�[Wu}CgecD�2�q��Y�֗ǃ\��S�YZ+	x��{�;n�l�6'+�Kj���P���v�H�)賖�Q�7y�#r�yO��b�K��(�h�Ǻ���&0dʙ�3�&��]v�5�!n�N�N�E��N"��[H�����7�_eE8n�}��O�1�OvV�����d�89(r|ttN���m�u�ʳ�*e�̙��a�c��u��a�Uǔ���d1�oW.n��� o�-kv�{j�NR�����0[�۽YZv1:��VE���Um��H�-�ڑsq%�j���lK����"�S�t_f�f��_?����w��%�
�0��Ѣ)27��2TiwWD�,�#";�����jf��X�u�EQ�2F�vja�lcY&�h���(ք�TB�b�h����4ͱaCwtc`��2L(�CdM��a�hL�&0�2E5$�H�"�(���Ii0����;��Θ�*O�b#�4RX�.���-E���.�ɂc0']�+��.��B��u�$��Q�˕��r��\��<�K�H7w.�Gv�wn����Z:����x��^tu����cN�F�s��)�u�+�u�]�]u��':ww �w;���F�v�N�;�wu1\�ܝK���wQ%��ts��"ws�#���x܉"��g��yN��.n�r]�aȂ���A;��$�~ϝ�;	l��3����F�J��]��%�ã[�v(�����L�PZ΂�c�#�7���m����Tʹ�2����g:���[�n9��gy��g���4�mc.�zB����F���_E��^�n����0G���Ŏ�+�%��>SK-l��i��^9���z���f���$��B�K���^M�.뺜4m"ς��c���ޥ���<��}hjC��No�S�罈���*f�;(2�Z�`XW�!�DҲz�V�����3����O=�)� ������
g%�Q^��D����x�oM6N�������LO:���60��ǫz���-��P2pD�M�L�Ⱦ�7��(F(�]�/9��7�2��QQ,���YB�-N�ol���ȧ�x�]��'H�3	P��:�6�j�Wv���G	%�:"S��l"S�]"��	Mm`Gd�P|��T:�wC��֮Q�5k�i5��72�R�F�:0�0RrT8���$�b)9Y��qO0��bˁ	c١�ٙn�;^;y���L#��_�=K��z��g(����пÑߩ���<�\";-�"��ic���Owu1�f�D�>�|`l
9���#c�N�䜚c~«Z�B/����7G��\�.�I��{b?�ur���j��P���ʸ��͇���uS�0�v�E���b�XtL<_�&'闃���%�B�d��1قN�,��bsz��ρ��4�A����ݣYշ��lWI�����F�W����C�[V�x�gp��QG4�j�D��������������ݙ?�Ό������mvG�浪�v�}�������_���\�[�W�``b���z��U�w�\�z��}4]�!�2�:2g8���gŅ�(L;��5�X��z}[f���u��:$wUrm}�eZ���Zw�,�1{���R�%����%�z����i��C$�ߓ����䢋W�r1�P/a�����z�3,��x�W�Y�<��ɹ�D�c��������aΡ4����hc��λ��g�أy-���Z��]z��YvP�g*d��i���^�]>x6ϳWƪ\���}��ƉU��
[-�	��s����k����\�O��?4S��l�S��)���ȹ�;�B�sY"��Oy�_�)*I}�ϖ�p����ԖI^H�0Y����3���N��NIݳX&�`�]���e�gv24R��@�
����M�O�ga�-@�4�V3��{k��s��3?�P-�����=�G8�;VZꈞ�����16�=���C&=tB��r�N�-T)\�,)�=0;���z|J{Q����:�V�<=)���_뾓�k��=�� {[�%=�K땶t��,��T�f��U��	�Ģ3��mqs��t�u�\�\�W�V���'gj6�b�ӆ�[�݀O�I��7����뒸�I����p+�dRC1I�.-���?ƶgGj���,0\��M�,�^���j���}�)�s�d��D��+IP�bU�͍���뙂��x�����'a<��z-��!�Pq1������_v�z�&X^b��2���=j~Bۧ�ڸwl����c��#��6^����);�@m�f��sH��ꧤ^���P8���SQâ�:��0l�G7��K���⾮�����T���y�W*X<�t����*�z/:���st6�wA��^]\«�%s�PT����!�a 'x�f�vC��p��l�����u���79OV�۾�)�^-�!=t,ߜ��`�E�z�O1�
�[�K���8٢��4(UB�,��
6#N�����	ڼ����r��͵��Bպ���l�V�����%��'�٦'�����-�e�Z�T0G��`��涥�m����ڰ�@��6�9C����_�ӼC�:�����Z��^�@d�����'��:��K�x��	�<F��d;$�6���-�7�gp���z�y����6��CL3v=f]��-��l��k˼ ��3�0���|aQ��l�~ߺ��/�R2v}�ʑ����$�9���k~+�{׃C�	��'�v���k�"j��K�p�x֯!�ڛ��N��� �2Q�7�v��&�|�N-Gp�2��(�nf�G�N��2��BǖnH"H�V���,+(�l��R��UNn���'<R��[qv�E�y��@���7˩ځ�ȼS�,�	A쿇�|<�fp��+5����zYO�^��<��Pyn!��P�hy��n��b��{����Ut�˽x)J�n�'����0^��N|љO���jY3l{�H\��A�z�P�a*:���Ӎ��oq�j�+�if�"�Wf��4�ϡ���C� �]���2[3ͣ��M�9HL�֕
N��y��S�r�-���1�/ԿS����z������-�!�&B�|Cg��7!	�y����� �c��Y�}�v^��)�`(T�c3�S���o	�[�Hp�ݒ�%�����C{�=��l��&�)c�'�m�kyx��f{]bx�t]H�Lh�I�s�8��s	���Aʠ�g�_��y$l��s�և�􍃺���+˧��ud�s�):a�aK�����Њ���|7�hi ���>�S���L�Źa[^\)3k! ���Ɔ�F�;JSz�qOK�zO̓�"�L?5��\8Sl�4��smd�ֈ���A�0�l0rŤhmcBvh��&m�l&�V�Ta��w9�
�w;y��ْ�a��z�RZ�Vo/3?q�\=�eAr�F W^�ٲ��|�oW* �|e��O״�0�\+;�+�f'�o٘	h�uV��6��}�):ǌ�	��6\\UG8���WE.��F�w��s�HC/s+%�M{3��Ϛ#$��������z�ۏ������[�(6*�3�p-��&�G0S���ֿP��mV'����J��] -p'�Rw&��g����Eݾ�c=���`���РG�t�#�ȇmt� ;n=��l��:x����g�w���c��=�m��x���~1��_%��1a��j����1\�^<ލ�q�����]��p����llK$���zHzZ��1�tE�j��4��D�ǐr����г1���p�|`�%�5+���f�\d99�0R�A���F���o�؊�����l�ޏu�D�U�YС��4?�s"ۓО�ǳ��9�73Od�K(!^�%�;z3�S�Zy��-(��ҳ���e�� �X7GB�W���,�ɯ�=lE�ԥ�P;0������쎛��/A�n�6i��XÙ�Pz����N��͍#��##�_�J�[�����i9���g��������$���h�'�J���Bޭ�|o;@A@�"X,�&BA�&���CK��sl�}�����r�PQ'9D�/`�4��(�k�Dn>09�<�Sۼm{)_�����������R������W�K�~�x�8np�����i��T�y�	�2�++��Otʕ���4��"n����"��s����jf*G����]�1}47��H�݉���r�����=Xw+fwM��˼ἥ��[ײ�W2�q�������_�?~;x�<�9n�p�X_עG	�d���	�r�	�(�B�R2���}�P����L�7�Vl�Bd��vme�[,�Bvx1�a�`�BoCiRO�"��
��kUs`M��QT(��-ð�u~�lA��:m�	���ugM�:����s�E���ո�q����Vf����Y܄����t���>h�a�Ϙ(�|�\`��`x4��c�gɹ����Me҃X��8Wa0�!׉�����G=7��������7s�;'�Bz�s��\귅�!�9�����x���+ѹV�`%)?5���o[M��B��l���p��?0!��Yϯ�]�+�d��`�u�S����BՇR�u1�e�h����b�%x�Q����T��E
�;g��9��f��Y�=�2�=mCs�v��e'�%9�`���z�J(�y?t��B��2�:坸�]f�V�p�ៃ�;Dt&�D��7;#Y+��}�:���4]���Lh�q̧�SUmf^?U�n�w�X增5l�wA���~l���\��m�o*��/��_~��R;��B����a�^�ë����d�FWNs�f���uz�]��X˺�@prt����-�UĞ�o��f�T[���k���gj�4����t��=����&�=����[)��KB���vh�����o�����z.����}�{�^�R+�u�����7�LK��[`o�&]����P�f���,�*o�,���m�N?Gv��]����.���{�^J8��b�\ ChH�3�͜eC [:y�x��8!'�ݳ9�W&ˮ�y6ԱF��*j}�4�S��m��X;'�Z�,R�o9����eE����fA2.l���V_�%h�/�8���nFy�v�g=tB���-��Z�J����2�^�v�Bڥ���<�񆮗�6<	���&Y�����{,�'ݒ��;�I��Jua%B����PVM3��16�;ݼ��b�t��$,�h5Ӎ�>5äH��U����� ;�)�{�b)��Uk��4�^p�!|6�<h�6^���H���B1�r�zzA�a�,��՞Boۼ���t��;5C!��qyo`�Ⱥ�^6.h���=;�?<�m8Z�[�����/>M���lf�֩�s���R'�I�P9+�Z���^o��,k��Cx&wvj�d><�|mo5 U�}��)�o�p{���Db��b���>�S�X���uk��ͅu�$��}��������~�<�D�����ՠWpa�7s8����uMee
<�3:#W��	O��-�u3��c���^�7�=�����0���CG�A"�'L6jC���:K��t��&*��u�T�o0�SX��`���m���L�*C �ܸ4oX���%�������a��Y�e-!�}a�X8�8��1�9���4-2�n;�˥k�Q���A/�1�d��췼/*'z,,e�a�'à0A��ls8lNpmK2��,9�
T]nl��p�\�C��Q�7V�s��^J��R���^��"]������m�_�'=���v-�}nP0٦*s6�i᝽��/.��j)f�z ��c��tg/�ދB L��ݡ>7�E3�Snon3�����c�vy���A!�%�����eC�m᎟@v�[͌&�l)5M[�3�a�4VJ/sQx�כ�5�-�!�<�HW��[�:l鋇M���y4�խ�gu�Tνb-�:��S��cW^UKcW�)��vej�IJ{<��w,���"��h7]������0��T?W�S<�sF>	���s����������"g(	�{�w	2��qw�ʷn{7�
�^��B�t�4��]=�� b�0�0L��P�5킨�H�3�� �)_���C�O��0,�"�]���z��	�|w�!��vH>`�Oo9n�%s�۳�s���2�sb��O��i�NX��M��t=���/��e��YbG����O'��ns��آo�T<�K�o@�zR�
���wH��D��ٙ�ť�6ۙ�%���u��QG(l����4x���NY�e�����]Sw�C�{��{�q9�Ś�w�G�,���2��/Ⱥ��4Q�~��sL&S�4zA�lo��-�SO�Dn'{V��s�N���9J@��0�r�E�{�=^�c�Ք��\��p��t��O�/P�u��=��:X�t���ƻK��pvT8���]/V���ZPX�]%z`���^��C���34u���-à&�>Ha>nmg��ݾ��N�L�Ԁ�KpQ[&��w9��z��� ���~孷[��Y�y
�<���	���l?07�`�_�ӳM�稵��!*��q9�P��X�:v�S��0��s���.���+�f�z`��!�?���Dqwf�L���n��/� �2�7l�$Q���(�B�1�'����>�rb9��f5���0����4B._b�٫q��vYm���u9 :~�f�v��K�/�!�Ĉ(x�"�t=1l�C���.���h��Us�Ow���`�>[����f�Yƃ���
_���8!r�v-����e���nQ	���h��;��ݎ|��\K?ֆ�FBi��==�gzF�{73M�,:�YA��s_(��P&��vR���������9��Y9����Ջ����)�h$i���꟠��R�Cgæf��U���Ջf:�\o��n��(�U�9J�;�_rKky^��d��jU��*f�����}:�d��++1�]J���T���ׇޏ�����< ��9��ڻ��6����ͼ4��<�Z|���ꜜ�6&���B�@�e�K6��/T�b�B�շ���׼�5-3�5�r��ŧ�z��]"�����â�����O�5Nݳ����m}Cw/ {�m��A�Z1)�J��z3����c� ���,np=m1�=f��:�v�8�׈a�����MsWD�W(�E���4��Mn�om��Ξ�����Y@Q�^���x����:%;7T�k	��HC�	~w��1�X]"��e57��9��q#Z#yu���[X�a��<���m�'g�*�,�H9*H=J�|"����)?��4�ܩ�quQ�lݣ6^w<%�-�1����a�<A�D&����
!��jO~[��Z������R�+n�h�gu4_v���@��_Rh˦�D���>a��`��}G8�ؖ\�����W�H���`u���h_���S�y�F{˸�Mv�2F�T�Z���� �̟��xrb�����V��nk'���r���P�[]�2��^#&�l+�F���3y�)H����lSPB���t˗N�]2�,��.�εmk�L�5�61��gmN�ūz��}�; ��K��B�%;�D崣�z$�M6~�0Ӑ�b��^_lm���,�!�N��٩)� �t�_l�6���ۭ�j�Vvs�#c��������p=ygmu�����@���C� qeम��I�^�b8�f�������΢MkE���:�yD�'%�L�G�J޻�;Ee7]���/U`7��fD�Ont��e jB�jm�Z3"�rM51j�Q���ɛ�뒬���yP4�cG��5�Xz��w����L�L]�C%ɩN'�����]��&�k8xS�zJW+�1����rõ�B�
���U��gZ߆��r���,�7]+ja�[���!��\�R:)Y�|3l�j���6>*� �`�z��_%��m˝:6٨��������JC[u1؂�_=n���}�>�rc��0yc�ACW��-���ݕY|kR�9Vڐ<���G.$`=��
B��N༣8�S,��4E4�b��ۓ�Hʄ�r�M�L�	9����ײ���y*��R�Q�(-9��wMz�o�T7�R�*�ظ�չP!�	Hݛ1�R�P�)f�[ؤ������fl[J�YB7k�-�{s9��m_u��o�������Ax1*��R�Z߭��I+�uqR1�;�hoi��iq�pEd�����J��ُ��
��E�c-����}s;�K��w��%��e;c�G�]1m�]s�f�qi��(-�k>�?3�L2nKA�[����G� m�~�hde�f̺&�\N8C��`�'S4z2d���Q��8ژ�����ViJ�-���iW��PS��u����W$Q��[����t̕�{:�r�%;�iR�6�a��V���]�C�	�T�ɦ�:���3g�K�&�rU�e��l�=�:�G!s7k�Wu�y���v�9�Ihue�ܝ�o��������=hq��6����s����,�!�ۗU[s>ɬ��a��4�r���W|ᩫsl��U�q8�t䫀��1�,fS޺����W�'8+dܼ7-�RgQ�3�3U�m�T#20�F��KI�<�*D�W[��k�d�L0�aV��son��HYKlX���0�Ė���T�M'����'����o[�y�@��|�G�w]M�)���w��<T)Wd�~�yŤU��Y��T���+Z\��-�eu��q�T Y��E�Z4�j�I��H2���a�o��/;B���e�3R��v�y���*fL5�=K���h��J���Μ�����'dhT�%��O�[�ݢ���r=//J�tJ(�Q�����f�h�2�y[������_u�f$���
#�uv�
�Ft���7�F��[.�$k^�o�����JrWx�q���08�Ԉ���w��nw!��f�HS.�"6���n	��%��y�\�q*�֨��/��;����������I+�nL��u�E�r��Ȗw�Q˩˔$��l'�<q/s�nw+��S$�Awrwt\��n��덺���\��w:��;�N�h6���;%��^+��U�t�5�X�F��]<t��ם�����y�L�5%���K�����Ñx���#&�-Ҋ@�L"22Ƥ�#i(�"H��]cb�I���\���R�	#�D��* �$��60T�EF-&��6&k�M�!a$C���KIj@��E�%F�C"ŠI ��&do�%C�#��nW6	 �TYLX4�"(�h�F��! �"�Ϊ��ٕ	$��J����s�"��5��L|��2ό�-]���@��f��˙����]YZ�����Z���.1T�
;�&������m�x�F�x��.�P���������/:�s���&�ک�~����8}:r�H{����x�g�ԦLcYc�=>�J�E��C�A����PT�0�$Z�7D�|�c�^��ρ�&����Vܱ}�wp�N	��e4���-I�Kmw�5�m��0C�Vr�ol��;�gg��&v�`PY��9���oH~~s�Mq�.Ϛ�������Nw'O��Jq,�%�|o�½>�t�_��VxZk���|���OoO��S�I��ʡa���\���̩�v���a�m�=�6�k�"���/�T�K��E�,��5�}��K^�v���O�y�8�C�㐃�I�Q�E`�k��}�����������BO�.���5vC06]���bvG��V6�X�]P%�]6Ϡ�c�W�T\98��}uR�����䶫���`l���c�v��&?;��yE'X��GҨ�S���� ���f�Sѻ|�.ֲڌ�T.0x�ޅ
Y���$�W���{%1j�'.�u��,,�Nw�u�bͧ;S؄�Z�[�[�d[B����b�	2�2͡��;O���Cݧ`[�#�Q�Ψ�b�_��ܳ�E�����S��n�uI����P��2�3j_����7ܭ�=�ƀ�ʻ�p"jQ�z���V�4��TΩ�tq*
ۺ$w�H{#���ftȯ�D�鱒;ܙQ]q�i���^�q�#��R���s:��9�s8��R!U<=ܻRv�nr�[�ޗ��U����2�W9�o'F@� �cLC� ��1[��K=���6��܆7!�jE��ROY�m�:�^6.h�;5�N���!��G��,�;3�gʈ��٥T�j�W:��O�=u+�kT�	�rW<�z��/6T�5�v��gwf��|xX��+u����m�:_�jL��34ܟD����*�_X�㋲U-t������^�>�$_3PS
)���ܫ�eOV�ץ�|�7�1d��==#�k�ƅ��X㭗JװT���U�U�qM��m>WQ��]nӂu�PwY�����ghLsH�����2�΢Ú��@��l�D�r�C`Y��уF.��t�i�J������ߡ�9�"]�Z!0��oѐ쓢���6�X��+�7���'l=s��Q%ځ2����;a�ƺ���k˼ `L���0�x���8�H�ɮ�����6��꠶nl��ȴk�d���O�t�I�˞)���}�m�l3�f"d�C�J���b;>dq}j/��as׳a ��J	�J�r3��t��#��8�/��1P�w����l�7�*��-gfVޜ�P�H�{�8��;�d�:zM�̾�>�z�9K�����97�w7fGJ��(S��Cw.��u�S�T݄���=�IX�TӲ�=�ro_^2RB��m�J�&�\�mjN��곂8A��ڭ���䣶�~�"9�X~.&.�ľ4����Ư.R=�>���P�.���D�zsX��9y��ʹì3�$��sCc=o� ���������d�mT�5{��M��}ӆ&Lu]��n����HO}�:ze>ܕw\��J����:-�����ح�pe��EZ��9�Ѻ:�x�'��3�s��`���B�F�c־��z��x��^��$"�)�4c2bɢG�o7e���`.���ʯN���xd]/
~�c`�I�y��qOw0^����+������
��kE&nQ�sН�k�(�z/)���]$��Lqt�wNZ;���l�`��_6e�8�z�jn��M ��b�C�ttČ7B���(qU�*���~n	Ac	���n]��r��Qۉ=��[XC�I@}�����֘��^��.�L��MȭUz��^Fl�Zhwu4Q�[/r�7As�Y9轸x�l�s�ǭ�οW�k�ͪ�2Z�I�;,$U8���&r��]��۪�[=�S��.���T3a�E�~�t�Ü<�^a�]6���^I����R؏�`��M��!s�:�bk��u7�_`�2m��t��Yu���3����(k-V_�?[8��FQ����PKr��!˕�"K57�uN�c�$ś�c�VVΓ��5��Jjw!��lȝ6q&��)�����R�b�4Vf#6���*�q
�������MV��Nٯ�6�p�&6�;�q��3�ǯ3�Gr@f4b�;0�p0#Elf��ba=�[^��n��K��??Tf�vިE���zHz$@9D�zA�ź��na;l]S<�-��'x��y��~���}�49���'c5��4�mc/C�$�hH���aQ��[�J�&�n�P����=��;� D�SI�,�߯��aV|�s��M{�س¡,x�)���lYl��|����CB*K�y��]T]�4 e������~b�}8�<�{3���8��LZ�4	�D�lؼ���L܀�k��8��$r��͜O�4��"��`qm���ǧ�R���rbB��������Kj�+�BSm�2�&�h�'��l4�ǡoQq%�[�=�\�0�����u<OX8�1zd,>��+$�5�A8�Q,���Y�����8'�Oۮ�~��=v<���#���u�a@R:'��*^9��|$#�Iz�N�ሔ���E1H��{g���u�]�I�ɝ���fY0â�Xp���D,�^���� �q2yūI˼�[^�e\�Ӗbc/ɯ���w�JK��r^��V�7�,I7���4�J�H��u
%#u�}�k>�d�Y�������O�9g�E�s�z}�9@yKۑ��u\�wxY�{WKϊ��"Ҩ�x���6�VpQL�����n���+;[&�VE.������?S�z�Z�k[Z65Q��������ؙ��5���	ϊ���.����<ǟe�[�G�9�hN�p~�鶢�uL3tSP�̹J�lf4�K5�u�/��'�K�M�t��zC���`d0Q��G8����$���v�i��Q��v7��sr�����(�P�#X�ג��'�q�b]��3���0��K���}�ι�<�Xb��kz�9B��="�Ђj����)?6#�J��yUK6Pطvm����ǽyΆWLv�;-�	�+�����	�~}��hZ�:�é�k,{G�ն��jv��5��(���t���]�z��~�8
��/����ev�Q醒pB1,x��v%pyv-n�)��u<�u^�i�C�~jOa�FtK<Ȏgl�\L,sbvF�[�������o3B�˥�wS�A�]��~w�,�4S���%�<��m��X���\��m�����DCSF��R�{��9��5��O;RS��P�e��X�؞�ͼf��{��`J�1t��f�֘���b�-}�}5s���lV��Pq@� ũ,��pg�c�l��;�7�:U��0^ ;���'W^�Ϧ+9PN| �㢍ޙ#��rT�7|I��j�6U�3�kMI���=u�Ƭ����/s��`+���q�����y	,վ�g�w<ó�98����E��Y�����n��-��U͇ۘ�!�5ӔAi��:�';[��s��:��W_�U}�����6��+m�kh��}{����߶y*�r��;]�1���P*������B~k;'�j�K����c�u�Q��ȵ��š7�Y������sb$����zu�P0���e\�(���*�=F�Z&�^�0(m���:��{7'�V���XR�K����y�r�_�*���=���tBd��_M������޾�TC��]*3��g=*�qo�l:ޚ�oH!�66e}�5�:�1��o�R�L��[�����X�b����2	f�Ӿ[�	F@AƿC����/�a�;g^J무xmޞ�0At	m��T2���͎Sl��/�qsH�;5�Wp\���"�p�k�����v� ��858�+]�v�k�?/I�o�i0���\���j�?�IPX�Ɇ��ݚ,D��s��kDu��ON�=��,f sqx�u�Mгnd㋿U�9��u�&�S?UOL"j��)f�a��xڜ:.3���C��������jéX�2�Z���.��+h�V���챼n"�r�{dF�=�y��̘�y�~j��f[�:�c���Jl�E����o����枆�7�C(�%uJ�7 ��I]}/6n����J�Y��O�]�0�Ut�;�A����}9��6�6�wwL�V���\zk0���Z��c������M(���nn���&�"m����!��������궓7��ʀ� 
�(#�cdֱZѪ��ƶ#^��]�C!����c�X�P�9^&��������d�\!�S�mܔ��0b{B���ߜ�c��ޛbn'�,#�bK�x�f�z&e�|tE��tg/���	��J�X�3�p*��Y�<ۦ#.q��oS��yC�2	@%�].��-�{�m�u��N4^���s�Ո3/H�:!k�����/X��3`��̈́��P!��7�r3�B����Ӫg�*�V9d.b�������\�)�z&���cW_��[�\�.{�҃-�B-㼫'ݴ��9��̝�����/�������	ѕ69�tS<!	��`�L�^h�k ��%cj��K��9&ʑ�&�0^�}~��e�%#���
O~��B�Fc�M<4�3��[HN$��/EQ�M,�W�ub	]ܼCV�s1"g�����U���z_q�=�;�`�ʝj���a����]ݬ��t>�K���W�|��4̤��"��4Q��W8���N��n޷_��OFu�0N�Ō�Ca��!0��=1�"D����Y�N�X�R��g�=ዩۀ��w��P�Ҳ�\�Ww���!W<7�F���LF$�������BRt�E�}��Ѿ���m���/���'<�L�u�+�|jRL�Ӯ�y-�l�Ŋlp����d9P���qS��ʌne��\��':+B�����kM1Jfu{ZL�ٛ��W�G+� �Cb֣V6֢��ժ�3x7�7���!�q�w������������&5��Q�v�8������Z~i��9��wg�Z���^ol&:�'��\>��}�:ni�#�Н��A�`[p��ei�s�S�O�!
��S��%�ں�K g=���ݰ ����@p�_�vi�]]�9;!���{�7�ʛ��Gmc
*�ԡ�%�^¸搮�k��=���0g�P����xըj26���ku��n���Y�vX�/T�+��1��:�/��qɈ��w%�ы�g�1-����SS	ӧ�8!BDf���|Obv�Vl�m�_�G$��.���߼��%��O��bi�jV׬��*�w�����D���z�4ϳj1§��)� y��M*�h.s=�y�j�ow�;!O���EC�<3�BiiC ��{d�9�������4�$�{gp���d�{�XR�vP�J�4v���+��������U��/��Ŕ�����uN�I�T��T>��E�Zi��l�ʅ���$r��l�z�o
�H�x[E�E�����vMʶr�����`IT+q�v*c��e�8.[��0��+��|b���;CM@Z&�.�c'C��M��)��T�9ԑip�J<�+���oFy��ď;��#fe5ʆC�B
�IKH,��tS���n�ݬ���-2qjj�W���]ߺ��Z�Z��Z-mՍ�[h����m��������h�Ǥ��z��a���z[��Bl��Pd��Fi=�]8��ݾzޭ�[�N;�tEK�t��f}|���!��"X^D����:ǢN+�K"���+Ti5��=�Y6�*���M����}�L_�b�|uo��#�d��͔%��X*���<���'.�-�-�-�m�.�;������{��[c>�kz���8����a)f����f�(p|z�$�֙-�z_�����9Y�󝜪^�1�]Xk�sQ1e�>@o3��PA�9�hN��覒�UT��p�"&����؃�z���a�J-?$�	s�4�]�3Ǥ?y�
9�C���E�qD?N�[
j��N�Vü�{��4�o�\P�#X��Q��|w �v��gaCc|�j�gNK�����Mx[�!�\��):�&E1�&��L$��،�yU��ݠ.���")L]��(��ǣ��w�2���<xB�vnr�D���~ҤVs�L:��M�k���5͕�[I	�'.�VwIr�C��;�/t0g:g�!1i������k��~�a�����|~O��)����-ݏ�8M����p�u����~�K#�98����u#tU�����������'u��3����j�V�ǫ� �(ŵ�z��r�Q��A�l�oc��苩1�0g�kj�h���I|�n�\��%����,��!���us(~C�#�onן���[�kZ4kF�TmI��6��V�[�}|��_~��Qv����<Ŵ[��/a�G��D�H����
I����O#���P~}�������햗�{@�%y�v�Y8�d�Tq!p�O\�o`C��q.=�i���Kg2}�Ƀ[J4F�w����g�/-S4��+��%ޭd�J]�:/L�.���d�W�>�Z6�`u+��*eg�9е�q�����Rѽ�u��̂Y$5$g�b�n@�t�������R���SK�;�X���>|Ǧ沂W��]�B~k;'�j��%�3�Z�A�� ��5��'sT�]_Y�̆�\9�\g:ϬD�^��v��u�W�as�D �^�E'Qx��sN��U��ǵ����=t3��*��2�lQp�1�$Ao@Pe��'l���}�)�d��d��<pٜD��y�tb'_�%B�ʢ���:q��ȶ�^8ށ �Ƙt���C+܊T%���3h��?3� �%�|�*L����)��q�l3e�;�0�h� ����y[r�֝E�Z�/�vB��z�Zۨi�R���d]g�xӁ0瑴�sӿ3���z|��g�ۺve˦Ye�YwvckՉ�fokSk�ukM�ºջV����齢ܫ�	�u�̏#�k�Ö�'fc���*�S>
�����<�]�]-�Z���6�ԥ��Ny�۲�`:��䷚c1�H�1k�y]h_���uYf���,
��+6q).˝I���Q	[:�fm�U;6LѮS$-�)*[������,e�g3�(�s�#�������DEٱG�h5Ե���wV�t+	��0�4{M2.ka͋
)����i��1>�"�83k�z��,���awO��E����w�.�9ջY�H�LG��B�o8]�n�#0�j��cws�kRF�d�,��[��M+ 9i���n����ї�7Q�h[/��B�-1��}�o0Id����n*D]�".雉�3z&),�K^Tzf#<c���]��E�V���� �sL��i��@�7wf���
�voܝ�V��d�g[��/xL�M�R�8�}cf�9]6�4�><of���r�Ӽ�Q��R�*��k��Վ��f����x���Տj8��Ѡ��b�-�f�1|�4xw-
�ޢMF�����k/t�ɸ6�e�6�5��L�a��+:nfB���6D�~O��Tn��)Bb���@���h3U�N)!}I�yQ�y��r�}]y\�ʘ#��zZ��;�-栃����<���J�ͧ�	[@w�I��aS�x��[��8Z��kz�i�8W&�"��ٻ��0h�Yi�v�����R���Ie�E]�_b3�{�Z���I���&Y���k�MI[/��ɚ�k3Z�2]-��[)_�)�c�IOb��wo33��R̴�c+l%�y�8dI_T�%K!�h���`�4m.sZ��ys����Wg^h�n��OX.]�t�JSvp&׈���]�nn0�\G�N�\�t���@��M�h]R`�����5���2Y �ȩ,�*��"%'�6�u��׺ї���A��p��B&L1��x 'f7}h�5�5q�Uxa��sV�R7��%n�� �r9<d䶇-��	�x��@�٘_2p;�.Xl�r��vPh<a=�wi�������,�R�q:��+���&�1�Vt� �ά�[e`Q]<H �Q
g9�U��,�JWl�C\��'8���/;8�Tl�v�,N۾8�����'M��C�W����2��컐^��W	�iJК���SO��Q�h*�]wr�����R�N�ڧW*+���'wb냼wZѲ�����<*#���40Tݷ��qC+(��f+������f5��9�Y���ck,^U��%�������7��YL:Lgi��G��\&N��͉��'��2���_�4��6֠�N���j%[�;��Vnv�s��s Υ�3�&gFN�j��(Q�6�
�(����Y��дf�3<N�N�k�o�/'-�����(�(���Q�ű%�ڏ�"ѱ�4i5�AYA2�66ɩ�mi667+�*CQ��lb؃��c&ш�ƨ�h�j-hѡ*#!��20�4kI.�,��HF��1�AI�F��#��Y
,RV)&TF�w\�LT�ţB��4F��E�b�hƌlX��b���	(�-9�b�!�1b�F�������Xѹ��H�LQ���wk��h�F�[b�Di$ƻ��5�E&����^��3s�����{oǏ9���xt�ȵ�u�/�%�{u���%+>i*��R&b�����mi�LWk�֯K[�9 B�� @��(�ţm�k�mQI�֋F��[__?��P�2P1�+o�5<à�^9��$�
7��
9�[����/6T�(�����؈��T�:�wG\��ݙ	�|yp锰r��q|��W:�&�Y��N8��,-tsk��=J�����k���I����c\0g>�K�� �cBzG6��:��9�ndw]X]8퐳����i��%픹/n�O5�θaC�y����4�@|Nva�i
�s���4d�u����Ƙs͑�̺k�(v��H-�@�/E�3��.���x�	���0�g&�\����\,��9.˜�ޗn�9E�{�Iv�L����	�v�tE�O�U��鸁���rZ����~��RpB�3pSz6*K��m=�N�=yCΘ�I��.�i8"���dڹVՊtF1�"�UGŚ��N�c�DE����Ľc�^���	����%r����yw�'l����^eq���b��tS>L+�'"�h��h�u���KkW�=!s�GwOMSѮ�ۂ!f�ԀӔ+lh뇭��.b��{b��!64��- C��ig ��7o$x���?A່��P�8��q�H�C� u�{�G$��tzp$t�'�D�u��5��)\)�A�N�N�ӔV��M��f��+�v�k�Q�ϩ�]�	�.�ӌL#N�Y3E��&bV']Y�3����{�]i]1W�Z>Kg�?�����6��V�5E�)U�-h�DV5��l�{��0oy�xxox�L��-O"�ߞ��<�~*Be@ZT)=��vzw^���i흡Ʉ���.��m9�5mw#Ys�����g���D�VħW䤰MP��w9����m��eC�k;�33<ʭ`�?;����/y��W�/�zF���`�YX���F��q�Ki�ׁl�L�,�V>(�C4���b!0<�'��5�H�^9J}f):a|�Qu��)����v���7JP��v{��;J��t����4��X3cLp��^������sǩC��iWC�i��\bD�R�-sU��"a1��a���\<{��:�G����ng!��	٤��Ͱ,�iyə��OD�}�#�{a=����w=��,���_>���x���ǘtz:�皸[ua�Ȅ�n��UY'ysq^�E�����P�ҵ����{\sJ��m�t[���à;ܳ"]å��5[c��1�f:��Z`÷c�雧/Rc~eO��S�Ǣfy��K1�����0��ʢ������� ̨L�Sϡ�_ƻ��6C���zQ~�1�IGD�^||�$r1{��R���j�h�wIn�]WKqhKq3)���ִ�͢~�z���n�n���+g*�#c�t^�gpLjd5t���O*�[m�Xl\��� ������9�Cf�.��!.9�"����%e�%/�1�k�=�N��������}>/�~��j5�6ƭ�cj#E�B�Eb�Q�[jM��1V-�x 
��枙������w�z`8"����LK�円���E�;��q��9���'H>�#��XI���ӫ��{{�r4�w�'�o���T9��,������n��X��Z���{�ޡͮ��}h�i댋���>��Bf��y�P+(!C��p��I�sͷ�u�=b9��	�FFS�#7b%���&��u3���.�ɜj�(����U���7!�g{�S߆�c dS�-���מh�uq�V�D� p���(-��oj+�܄��P�&>�f���^��U��LL�W.��B~�c7��6z[��t,(>�ò�G�}���\�:!��%�{�Ji��*4��^�����Be{���/u�ܮ�[�:zkw��,��;_M��`���ArIz)�|"S��n��=)��q�n�GlW�-�����O�pꑟ@���}��kӳ��f�(qt��SZ������#��r�tE�:���sW��/O���"�BG�Ȅ��x�JQR����s:��� 6��]0�-Bn�E�?"�%�I�r���a`�}������cY��둾����=2�5��V8N����F��RV����2ž�]e� �$�v/#������[���]|��/o� �2=-η9�|��m�Ա�\��Jd�^��7�&�]3��poD�S��#V�i8���ϔޥ7/���� ���Cꪈ�����b��lm[���f�s4�P�EĲǹۚn��kZ�a�^-@�0�>�'�q��ݵ�-��Z��Jܠ�e�-�u�X�)0|.���GH�tD��5�&����O�~�d�ʨ�yUK6b}��fr��vbv۪�|�l;5!p���0����ͮ���?>�q�j��S�N\N��DǶ�����۔�[{U�����`O�v�v����$Ini�9���}��s��"�/��&�4p�s����p��d��M@��q��?3Ӱ���T�ss�5��z܈,�u���9�'��wr��͡4T�"w����u�~2��+�]2U~�I��R�Q�h�4tL+��Off�a
��NN2��z}JY���<�[ �9v�|kOC�m����p*�^n�^��Մ����� <��ۋ�Y>Y��� ������!�1l��l�4�/�r�o>d�D�����}��r��������D䄻�QX��'�:�'>�K-����lg�ڻ6 �oR�u샏�C*.и΁�r,D�^��v]ɴd���	�̵���D�[�q��.�u/{��ɥbb�Q�[QV�2�M���n�ƏI����hV��5r�4����;���	��>5��w>&�^�Y+�S�p+��u�H�Zuh�HpU�Lr�:0Y'
DeY�{���Ǔ*']��_;<�4����G2�J�}��־�Ʋ������+3x����M����%B�ʢ��x'Eh���N��ʿ/0.2�~"�ީ:јFB۫���#�4��@�krt�	� ��j�QN-�-�vE�*�����������Lp�.�#�m`b�K7�*]�J�ˁx	���"��+�pf��w�xa:2;4R1���5X����3E̽�?_��p/�L	eKCM���oܦ�X��������h�lT�\�9N��S�Ӡ:h!�/>����S�É&�Q�0�aVas�u��^l%�ݲ�Rx����V���g���P�xwf��������H���OEs��t�رԭqv�,;��p��j�n�j�s�p�=-�R�(��B{������k��>�K��p]1�OH���4%c�o�;r��-�ū��m�WS�;#q��s�%PK��O1j�����3��i����]vT��`��bfY���;p{�6�y����jJ��6�9C��jXc�,���̙���b2�Ŏ-w��B�8�	�(�X��m.�z]�F�¸ėj�7c׉�v:��@�r���骲����!�X���8��{	��3�(s�Uc'h�@ܾf�8��*K��Xճ8�)�ʳ+�O\�4�,�°I��BT�T�E�P;���z�0�B��nt�ܝǠ�c����\���S��McV���FʬoN��v�;ȴ��N7���ث/��rq��>��}X�j�lVѴZ��������ϟ�z���
gD.y�ό+ѷ8����/�y�2	A(4��v�Չ�\]һ�oA�r6K���X܅���mx�fq��L�\H��I�j/��l.z6��>���
t	P�{���q7ku�$ w�C��5>S�C�.�E3�,"ä�j���^m�����!�&�~"7��`U5X۷8�{�r_Cr��*:��y�V�G�T���S^Q���b�^�-��0ER�Rƒ��L�M��BeV�
Or�(Y��{i����F44�c^Ľ�n��|��y�U�x`�{^��;�P�Jee�S��RX&�Eu�=J�f����c�l�^%�d�?�N�\�!��C��/�z�@"E�N���g�Ĳ.��)�FS�m��yk�t��gL�n�%�ss	�ց!C6;��'���$J9*E����E����7g]2��k�`ޛц��6"������,�^�<����#�&���ư�
6҇i��ƌu=]�2�f��]��a�=��~J��0����\?k��a�`鵟��vN�U��ؼ���o�і�X�]����j�[@`��k�vD6m*8\8�X� �>��(M����^���r�py[y�ԋ��&GH��7�r2"���;Tb��U�]��qk�܁��#�#s��]dkkl���SaW8�D1�����o�|�������V*��W߿��^��[5S�SC�gs������}��=f'��UH�un/_��9�B��0��uaa�T�BF�A���Ψ��]�Eı�=I���U�(]+^�T�.����l���s�A��F�ߍ���f�ީ��:��0쟙�ݷ"��Y\I������ӎLG6�w%��l��ΰ�Q������&��]p塝�
���@xA.��_<'a��{6C�����~c���T�eښ�_k��z^h����>`����T�3�� �, h|.$D���;��ƃ�ͬa��4�1{��Y�n����@� ��i/���6"���D��塐�-���=	�{)lcg1�������y�c��k͖`%�Xu%���K�y��O\�o#^Y�X�ii(Lb��V�Y��5�.�����q�c�Lz5� ��^��[1��(2�S�W�9A�ٳ����P"��x��Ƞ�9+��_S�vc-:��Ӣ���l��=�D���MBњO~�ӌ(��Yx��gRJK�q=t/纱t��K�S�x@��-�"B�Ed���t��Ƚ�R�d�6�v��"�=�tz;���7G*���Rd�q�4���
Jȶ�Y�uu&��F(kc2��Wl��;���5���+u^��'Ģ���\ �ن�k�2���՗���Qrr�pV��x��|8��K�cS��:?���:�I�����3y���UW�����=���D%v�b���G[��r�On�� ��Q%ٲ��0W�=�$���'��^�F����e6]kTC�o#/k�dw��#)����<͏P�G��ki��m	��ʆf����cnt���tGo<M.��QO��NV��ث�sP&,�>G�e�[����K�	�ƞ'�D��ƈk�{�n���)�����j�ia7CФ\N'�O!'���G.�`y��4[Y��xvV���A�D�d!�dK�=sM�3�k]�2�Ũ�{��2���~�y2C���C�:�B���;;
�%ݛ�����T�8�� ���L��׈ɷ�
��sl?L_���^�k��꿙��n��HP�����|�vn��	�~}��hZe����1����Ta+]M>;��h�W}���hҜ%x�Q��JDs��(�����A���-����?[��W#@%��b�����b�#e�ow#n
vi��;(�@�rŨ;��x#��0(->0������ف�l��+Y�/��Su��}t1gJs��"w��ˉ��~2��+ک����\��>��{ ��ٵ,�V��X��]��l�N����B'�jմo�qq�w�c�.�1�N�����XF�ؗi�p�<2��O��*���sA޻wۂ����L#�H��+D�i�ʖ�ܭe��*�Er�rsG5����]��������v����U~~Z:��`��LZss����=�>�yf����<�IN2\��H�ƴ��6�w�3f9�D��s_-c�eX�;Ч��qm��j����حj;	BZ��!�1l�1i"K���ԙ9�0�*��1�Ϯ�ӽ��,`��D>c�
���TV5{T����A<QvQ�7�V��|9{�Sr�c ����*.���r�?�8K�'�z?	�~�yP�436�nƓ�/)����v�3�1��%B��TXSR�jQp�1��-�Pe��^v �/�����޼�m�]ɘ�/�5(��9w�� �*U�ߢ�gd[B��o@�DcdD��g�%�^�C�Y���/a��h�]�ǩRe����)�ޑ��\�|��;4�J�:�Q11$�Z
#�D9怞�Az`K*CH�R���d]`%�Aj�H����\���R/0V�!��Nӧ}g�8{d-wd��g���:�O`4�U�\��-\���.��.�h����4��)kA#P�?��٨vC�ˇ���H�	��	�urn��0m���zqn�K��'��N�)mz?���ʝY�7�¶^�[�m���]�L&������×���9<���`������j{D�X%����+�JD͝{�-�G:�F5	Vzu�G��T㜂֗J��-�b>��Įt��.̷����z�x�*��[�{�u}w��?<>o2+9?!R��,>��%��WZ�G�֮݇{p��p��mn���"�Ƨ�sm���1�A�V֮����(�n9y�J׿���C��lN�5~�7�y���KYk<�;GSi�8�q�-��:��ua�Ú��ꁿ2�{�ӄ�71�\���s ��MP/���Qo����{���/��u`NK�V7�ۧQa\bK�,ݎLC�x�b�'a�p�Qi���ŭ7���Z?�d��T��<�gȿr,dse�p��!�LC����c]�7TS#�6���c�����N�W�)��lg	��Yq1�)<K�=6fƴ����� K�<��g���u}�E:�(�^k|�M���tS<XG�:N&.�ؚ�j庡�,��LΤ���C���E��;]yl ʼ-e
7��ދa��*�ئxBdy�Ahx�6a��,;imo`�ǣCr����j���t)���BeBҡI�J�vN��M<5�{gi�B�-�+f�ۑ����{E�e�%���}^A��O5?!)���N�֔	�[osk6�i�F�Z6p˻��Yt�,������>��9�'D>>���}0S_sXF;�/O>�T7HV�
h�+
��+�[��B*
2�3k�R�$x*}S$�=p.]�6x�Ӣ/X� �\Y��MӧiN�X�ma3����ZF�yڬ��z����y�"uq>((Ի�v�Y-���sp5c+'S�q��W.�I���Z�n�T���0ԉ}`C�|[���n����������],r�C�ʋ�n�:�b�:���YOd�>fح�zp���++���o��Dt�����]gZ�7iM�2	��`N���������0�ܶvf%"�p��x��t%+�겵[��Vcr���h�M9��h���D�^f8�,x�pB� �t�nkQ:xْ	�Ŏ�h+�G������ƛw�6<� r*��*������{CvAs�[ɽ`��q.e�f��]
�#��^���8[ɝ�!q��d����0B�q�f#B{�����@%���jAH����#бF���!�{u�2i��:��j�J-��h��:�ܜZ[�!,JR��n�5�dg}l��a�`���2��	�������̱K2C��5GV�8ۗW�|Ԏ�ոH9}ӭ
Ri&�W�Nњ���H�p��̽�Aַ�����2ݮ�3Ss2K����0?N�W��r7*Wi���Vj��gU�X�b%�݀�q�h刲����aێU�XZ��#Fu 	{dh��;�ai5�@Yf���q�H��&v�����[,��T�ĥg��˾��'%k;~�#�4�Z=z�04�]�_
�~e���ˬ
�E���T�{�V�N܌S�H�r�S���U8Wh�P���k�"�����r8v����-�I�b��tGue��S��{x�a�]ZU�"ר������o��;w����w@kYu��G���6�S����s��\-Y��WT���Y���|��ZU�h�W9p��ͼ㦌9�Ɍ�&	�p�طäU���c��u�g��ʃq�1޷63Z�̈́ty��ea�z;M�d�6Z*�&�L��Az�ܝ*��S�+�˧FL�V0��th�B�l��q���P[y�ګ�y��/J��V�
���!mlg��
��4��TgV¬Kחn|�:��sFM�Q��2=dc��+P����k���[�����J��[��r�@C��3l��jN7�(EJ��3lܑeMT�n�N�X��mE���FN�>Ӆ��tՔ��ki)x�q1}t11b7��ʽT�,�V�ru9��֚�f�3U��aҒ*¢�F�q�2��b0l	r�^*s�N�_w�Y��j�za:n�Q���\�T�&"�2-�ǸR���ų�%[J�WT78Җ��2�����I��:�g����.h��l��	���Z�k<�gd�9r��5,a��a��_�}շ`����z%�U0j���ټi�͝��X�N����i���YH;�w���8�s�B�Q�d��:��n,����o,�q�\ب��ǝ�{Ϟ�Z$�VƴZ�&���c��m��%��aDY(�h���F�b�h�6*,��lO�nD��X��ت

1��؍F6(�a66M�n[�р�ص��EsW1li5�5sW(�j"��j(�msk�Qj�F�X"���wv�j1�TmA�F�Q�1���I��k�5Z��k��F�b���؊ƋY �F��(�hѲj-رQ�����]�{�������be���W�x�[C
�:�����J�[h�־��C%�m�v���&�Spp�� �ƝqW7O�hK��ж�����A!l�)���?����.use����7[����?W%S�V k�(K�!=_H�5��2���x�t]KtS�F��K����8lowva~B6m8l��|��։
�b�S�CD�TR���0̐��>-�euo9�Ҧ߹�[W��;ux�r3׷M(fƘ�	����[�n�c�p�x~;O9��3���޵��;�za0�M��d���]*���p���|�=�d������n�J4u�7]��{}�N�)3l5��|U{O��J��K sIzp���aΫ�n�����3;��qU�^^���L��z�[+�c
�ҵ�%�^��9���Y��-��W:�'�3�4F^�W�`��� ��v��ۏB���\I�O���=����4�F!������=w��\�t�f�E�v���!�h�^a���:~��!�f�Q~������J/�R��C+�,�o8d3F+��-��sþ���ā����f�X8�s��xHm�a�iP��ǘC �w�S@#�K�l�<�"����,����2H��9�z*���ۆ�F�l��t���6��@�N�+���g�Иc���}ОY��MT����kS���V4��qŹ,,��tt��3��}$��|����[�/����p�/w�*���d	�`�CN�\�fl_{��3�ǋM�w��yf��T9�p�4�$���YA
�%�<�M���6�����~hjj��Y�\�V&sn��	s�e���sbj}%��g�)f�;(2�
q�jH������V�R9^��/2�UT��#а�Z�:�"��EU����Oq�oܥMh���+�Y�{��'ȼ˻�z�/_�O��,�3�8O��x"X[�D=�v�"�J�nwA8�Q,��9��6��ٵ��o+�;1[q��Ԁ��|njgO��� H02B�.͕/	��|$>�K���&]�#"��k:���Go/Z���6�E1H�jn���lz�X_�� �64�R��'��(Y{�l�jS[��*����)�p��I˼��n�J����5b���y�C���4W<��8��G%�fg����!�gM�:����t�Z~X�A/ZT���L8~δ)LUWD]�U�;n���� �`מ��C�O�b[��%�|3�k]�^*ԍcS�?��:1��:�gk��V�Sv��z�� �n��v0}�`�G�ؿ���Ĉ&���4�O�~�d��y���Xe5�
�j���*Gq-�����v�늜\7�����iK�8��p�4��tVgw!.X@6�k�*:�:�÷#��xu���Z7��2_��9�������ݓqV��hfM�F^EX�#pr���
$�B_0��X훙y����U�r��s?Ϫ����Q��폾�˪Y��b�ٌ�0g?0���$K��/^�����q�XŃ!U���{)X�k��st��Z4p�ڋM:�gժ^y��`Mt�G>B��<��h��b���^�L�l�w��KgoI��pm��a^$@�LW5�Z�^ø�v}��x���B�����Mِ�_P�����P<^{:S��s�J��#üx��m+�ࡃ�dK碴F�ᡆ�@�y}����y��W�O����vjߜϡG��g��Jq�nF���=vHޘ�cU��f�~�-��{�,׊W"����F0k{b_&��ޮ�حe��q�� Ũ%�CWY�m����f+��7��+�װ�2��l�����qx=�{�	���"nA7��Z����{����{"dPm��:#�yH�Z�Kmx��g���C*.��fp��0D�BbK��k&��;���4�3a�����G]tF��{E'V%B�),%�.�Ƣnrc�>�0iM�Y���7Afg1�3�a����Z]�C6�rS��	�{���J���E8�ӌ&,#?L@@|>~������\aTz�gUh���N����O�����t�Ve�]�O��y)���'�����Dƫ��h�;W�2��,��+Y/X�J���K8������lѦ��z�m�)�������QL��ۂ�]�GZ�5y��6k[7�\q����}_;�v�GLO`��gm!��641�_K2"�˴��I�����t�O@Ɓ�3e��M��V���4�Q����`C�_�	��0%��0�f�'���"�z��g�jR~��xMr���p�2[���z�	̉.��?<�{hX4�P�7cק����t(��{�es�IX�*q续��Y��]�Jm�{��5���0�'�vh��`��d8���Kq|�\���7�qQZ�b����Y���n�˥�!˨����d����k����nX0i!�������	�&��8|�Ϊ��5���k4/�:��:�eҵ�r^���a>[bu��ÿO@`��#�˶�˚J�J�n٨�����\׍K7m{:�jl�k���)%tů������:�r�3�	��x�j'����V�����[��v)�ޗn;�XhbK� L�z�3.��x�F��Z��=#�/�lW���s˼	��_=)�ۜds��� Ȳt�$=q�;]��w7��ifke�v��CC!K��V�T:&�W�3�`0&|�Yq"�2�x��zmѭ^������d=�;���l��hC�xm�P&��]W��vЫ�zL�j6�vMW��X���y+�˼�z���3o/Q�Rͽm���V��Dr�6�:����Z����:nm�rJ��PU�6#>���#'w�uK�,����F>on�=xU��M�7|�����)���b���B�#W�^n����tS<X@��8{���(!O�QO�Ϯ����r�6���ƠQ���� ʽk(Q��|�E�N����5�g���p�ٺ��b'��ִIx���;�l���[U-�C�	M��BeV�T�n���W~�gՆYC��w�U܌��e̺�<ɕ��8������أ��Ly����5t��k�U��͡в�u^�]V����snq�����i�������� 7ƽ#LΗ8ķ1��v��/�{'l����O3���?`s�K���]D'�}`"A�l��.z�CD�U㔡��>�lw[�-��U<���Ύ�����^&���xn�gi�P1���6�8zhAC64�8Bn��	�z:v�EU&[���u����7���qV��?Z�O�~J]&���p�����0t�Ǭ��n�MT���zqS���T�_��Մ���Q��Z��2�Gs���Ӈ�p�O��1s=9��<v���,)0��8u�hN�6�����Ҝa<�V��^��\sO�ܳly���^%(�M~KI��t�둆��y�˚kE�p�[o0�K(�b�����w����9�<�B9𰷳2�ێ	.�1�Pj4�Y<�B��z���pT���U�fM���1�=�%\3aV^��D��n�ٱ$�nc;�����yӼ�E��e�თ0z�p�h��a�]4�C����6�ʔĲ����ӎ��.���>�ލ�_��p������N
,3�.�����Cξ��t�@f�Xzf�����Y�R��=Ŧ��S�~��E@i7h�:"ص�!��ý���\X�Se�Nϧ5Ҽ�B�T�LCm���-����a �$={�@!����j�ε(�J��_~����X�6Ij>��T�����cy[d<S�z���73Od�K(!C��p�y6��)���ύ+���\��m�����=l0"��P��NnjG�=ٜj<�3u���*�8��{����8�̢��ؙ<�ζ"�t��x5]�8����.=<(�c�mE{x�M��,�iM'F��.���Ѭy$s�d��7����m]�0c#kDK��]��S��tB	����znU��Bo���۠��b���:�-��q�,�^5y�?22� ��H>�lHƨ�~�0,F�]gK�#�5u�:���D�K�K(�kk�<��������,��_�����t�E�������t�t�=��m��+��J�m�+Ī!���>����Lϝ�ӳ��Q����{I5�>X���S���oi�QC�`s��a��7��o{���#rhG�;V��ܝ��=@6��������97�uA���:{~���3��'ǩRO��Rr���ث�sQ1e롆��8V!R%���}��u�^��͂��}�*rx3{���K��0��0���#�� �A/�@�t��QK2�2f6�]���νb��L�
;p���"�&���kZ�a�^+��̡������T�o1�^�M��;Wz�cû!pY�B����v/ƀ��\�ęƠ�����I��-!x�Ps��)>N<p>w՝�۹�e�U��H��0�763�����v�E�z�hg�5��꠷��r��r�s�m�K�շ�	��G�tH�B������/���^�KNc�1����ۃܛ��C��I87�Fi�!�^�b���r����{��Ds;U�tI��Wg�ZW`��_�N��*��瑇:���~�.�aط���A�^�9��
n�e���֦��V*8���w���}d"c���N6ۜޟG�,�4״��j	N2\��,�7�E��	��K�d����t-��4��{��3dK�k{dkрU����3b�y��(���7��9k�#n-�1�2j������}���yp���{��?/L6eӒ��ӥ��3�I�]�]%cї�9^������Iv�2,ϯ1K��mݐIR�Fa��F7�')���{�&wmD�nr&�7��˶a�6u��tpt��[;�0�=y�9�ٛkC"��={6q���V��	_]yV<���t�a��c�u�]����+���+UOC�����\	(�^�j������v>5��sW��
�x.3&'���
.Ꙕ��iB��w*id����e�|����
W*�
�Պ��ҭ`.��ف`(����K��i�UݦlR�څ�p��%�WD&I��Juc%(,���]���d[g�������e�%�ݭZ?N_����0Age����W��CWv'�RdY�b����w�uz�Et�4��COKp�9.�؃�+�L2B<�Ð��OH �a�,��ijRy�r�d] �B�׽×�4hv�̃}�c QiAl�=;�?<�mA�טr��OE'0jD��I�nN��=A��f��GuxnڍהT�4��0L�����ȧ��d�^�鐛�Л��HCI�vh5tU5*�۲ٽ�w'��qe),���c7�k��(:�����f���
�Q��Q����B����J�3��$�b�m�B��Ԭq�˥k��1U�V؝j��G@a~+��Lv��O/�t_V;Ɂ��i�(\��J(oa��9������������OWV�b˸�8��z�������1ͬw��+o@�!Y�؇(�7�YRͨ%��9��]����:r�r�cH������ޭ�
���nZ����.U-�ٰjt���e�°�j��޿A�����38���@u��a��@΢Û
R	`�t�=�P�:L�sqe�J��ڳN�a�=�\4-�D����<Dsx����쓣����r����Iv&��`�I�ky�v'���y�ks{S��"�i@�~y����ߨh�/0�P�8��ާa�d<�YZ�«G�0������A��hbz���]�6��g��`0&P�.$Fd��/X����rlxT�S[y��O�c�s!F7��W����W#^i��[���NC�<�ߖ�e�f��8�}�R���W�*󞍵|YN���]yw-���Z����P�a*:���zq���9��gM��j�-wY=��c`��^���峌U������M�9HL�ZT)=�]�,�f?m��˴��b����ua�xd-�;AҜI��HH��݊9�?!)���)��),l��,،�մ�ob0O��Hj���M��_}o��[Rt��3�範$_����=s��D�>��'��o"ӎS�⌦7GEs�w0��XF���b�S�C�"Tz=�X����N�'m��A���]�n2%������֓e"_�8�{f�VAX�Yt�]�v��{�`3^��������+y���;��;�����ps\���)�r+�j��J=ae�JM=�{�����kP�j{5q���sH:�\��]j͎��Y�]NU�+"v�T��a׸�k���t����S].ܔu9e�p��=4�`���� ���eqP�v���;�m��rڀ&�V�\��UYU��j-?2NX����A8���!�{�tғI�!��^OE�CNM��DU;4���`[F�.��0�-Gs��+����9��8x�;�:-,��flOn�-1�oY�b`c����ڴ	�-l�)�9t�{A/WQW�e�I��N��}�����nw��5��l$�`�s���/0��ݷ�M�� �Ll2���Y3+����k��|�]��O����;�xņv2`3?�!������ח��|�Շ����g��yǅ��tj���9A�=< �A1^��-�W��;�t�y��Ĉ�9�����T���|[wX���2O�u��?^M���L����q�v-����0����Ain����xV-��pZ�v�<�v/�{z�4��4�=�Xw������^M��xc�#�g�d�&̽V��[Պ�Յa��+ˁÌ��q��e�x?w�07���eV����� ^�O����������]2�,��ڱH���8�1���Ԥ�&h�$F�,�v�RsW������|l k�����Cw��K�rl�f3���Iqy�ؑ�˦ҀHm��J�ڰ�����U�������M�[:�Pє�f��R��f�Xw�\�Mbv���i�3~�j�}��vΩU����s������T�c�{�bN0��;a�w����t�n>�՜C5��@w/^)p�
��8��Ok[�u�K�㇯��֜�GE�W./��V�!��s7"�S�$e���H,'�ΰe���Vw�0���A�6��rQ(����`G�B�M��r�bXi[<+�!VH�u>$zJ��H|wV��t1\^eE�D�g'k�(���|l��t�hi��SN�S��v�*��K+0�B1ʛ�eu5oŀ����XwoC:�9�v��9!�dh�ڝB��m�9�e�y�(�i�+s�i<�7pt��Mm<����,)��v;���@��v��p�	5�&�NI�[}���KZl>��"�M���&Cn�^�R�.ocCy��lgp��Xt��9.M���v�Sskg<y
���竵+Hn�S�7o�!6����T��-�u��ŗ[$!�|�os.�_'�QZ���9����c'ny<�k=��\j�n�~[�,t!���޳,�����7VW>��+��.�&�M�
0��I�72��c�L³�v�mҹ/u)����6.�Z��|� Kz��6[�8��ٜwx�zm��n�0�.�B�f5jS�0��ZÏ��֒�7����[u�k�ʣ�������ohu��T�t��,U��n �����6�I%�ZDQ���� �m���uʓWDx>�� Ik�vWwEbx[�6�V�a|��4ӎ'��a�숻c̛�X��e�B�}�+��ja�^�W9�E���W���Y��yb"���f���T9b�sKa�Ob\qi6���f:\����[x�M��B�g5�z��W6f��Ьe9}�Èf̆�2)JR�'~p�c}�Mc굧n��e�ZʅᑈeerC��9��`�w:��86�A%=�RB�֩3g�5�E:b(�e�im9]�ʵ�QT����ϻ3���je[8���y��ܳ!�F����M[�N�Y��a\��1Ym[��W^�9f���,Yg�M�v'F�Ω�ܽ�ص��X!ڲk�ف�R��;Y�9Nu�^��K�%��yN��3n�4�_El��ã.ӏ9�K�V��TÓ�2�p���y[��W\s�`�����i+%�_:�%ً���홄�oP7a���D0�ƹ�7Q�f���Bcw��"�j�(�k�J�{�'JJ����+K���(���T���I���H:�%�\OX��mފ��y�V\j�ηw���K|͠��]�*T8�ˡf��T�ޤt��:�Հ�>z�.z1Ԩ�5ǭB���);������(���ϖB��r���8PU׺+N�λz\dsx3�S�7W)��D��:�C����cFM&���h�[5����ZB(����U"$�Dk��+��&��(����EPF��7)-����E��F�Q��j(*1X��%k��DZ4h�`,�h��h���n��Ѫ6 MI��h�1��C��9QU�Qss���EAH��QsQmp�+-�nQ�W1b#h�E��sØ>��������ʭR�Ç{�0�D���lfC�к�F�ʀ@��g��\dJ�څ9��|���n��Բ��B�'No� �V��u��ܸ�����Q�/FE;��N������W���"So(A��M�UMɥm��,��W�����[�3��[�z��;��f�� v�"�N�]�ɉꮎ���+��\@Eᴽ��4��Mn�Om��t�On� ���.͕/	�Ƨ�f��g"oy�CU��
��z
"S��b%:�.�Lh�I��G\�6=C�o��֎�Y�=��Ο�_���������A�Ζ`d�q �*I��NV7H�X��sRJq;k��x�E�GfNTE^۳���
���"5��;<���mI�S [���'�hΆ��9�Y�ɠ��2�֓�2�u���8�
���-���ƴ�G8�ؖ\��ݹʵ���/���j���Ԗs��7��q�k��������q�?s�2~1�'�G@�����q����Y�٪x�Rڝ;M{��B�ɷ�
��T�f�;�n��~`Cqwf�E�z�]e��O�xu���	A��A�k,{�����6��`O�R#�*�Chp/Կ�}���'��B��v�M��?R��)^^P��?)��^�	� ��-G3՜�Q���X]�z��,%�{5|���Ϥ��On,��[Rk޾N�>@���6y[WN7c��ʺ\�f�&i]� G.��:��>v�Fm�5L��Ծ6��M�$M:�fV����3��^�?=�K������3v��e'�8�;(b���r�^ø�xg��y���lS���3�{eF��+6C�9�&���^�.ŧ�s��tE���yqQ:R�ѹ�q��[U��Tw\CA	�&
u~��m�9����f�0uإ8�5���j��k���~�W��i�~k/J��^���2�cql�߄�ϫ�ٱZԶ%�=�5�d۬��8�jd7�t5L�=xf�2��l�瞝�x!"��JN�{ʈ��bA���~=[��K�9��9踆7���z����z�8.3��%�_[4`v�S�.oh���l��������sϾ�k���^%B��UԻ'��S�>[a�g�ƻ��r�+o!���huD�;^t� �=�gt�?�N�$�Z�J��]����w�xh�z���EJ+����1��o@���C�J�q(3�C1��]��I�1!1Y�2+]���kr۹j�!��>���@�О�N}��; AF3�	���ʎ*��,Ԥ�>e�3��uc*/ݩ~v_N�M��:h��>�G�/�^�(�պS���.�(-�啥�n��f�^����������:�խi��A{����f��]֓6pyZ����o'L��b��Y����3Tl�����,U)�X�>b�s��1�5�tTgh�ng��\��lD*�����]���
�Q��_���q\e9�&�Q�{�yz0z�^A��k]�o���3��T"���,k��C	O�ݎ����|��t��_Y�~���;vT]m��uʓt/mԜqd�,�t���h�����٢�Рk�tw7_�}��c����W52Ad������h
�u��Z�⠗�R��B��\���<X����\��fu���0��f��Y�^?!�,�s����)P!tM�'v�$Է6��n]Bʪ�}����9�Mf��3{�&D���D&��br]�u{���w(�8�%��r��>��U�/�/�y3e��e��@�r���^@�n��x���
����Ϸ���T:z��¥g<�m;ˤ<�����N����D�+�ǆU��`P&|DYp����Ķ�ƛ�9�UT��k�V�ĳH����U��^J�!\�y�fKۦ�t�îo<�X���4L6g�4v�a��ap������|��3mڠ-t�A���lY�+��z-���sh�Y0�Y���9Z��
�_IS��إ��`���{�'0s{�i�S!q-3[�Z�ʺ9�dt܁�]��[�˒wl�5ޔ⩆�]b�%�{y�^�Ss���#�*�Vt��յ2
�L��*r���ǧq�567E�6�����7ܾ)C'Ki9.���d͜=⿐��5�J�`��i���Kfa���-�T�i�}�BeBҡI�J�v��v�/2�-W�J際�W��ǫxjkgkCb�K�!�Bo��4��O3r�qx��暡�9�!B��*�o �v-ā-T�k�FNc�m�'�o��[Qt��K�!=���g̗p�1Q͛��:r�pbh�:ѧ�^%���������Qq^{�����A�l��.z�����Nʯ7
�Ś͢�w3���y������J.��X�����u9fj����F����@���6nl����۝R$�iC��eWCը��֔4I���\<{���"�.�֨�o���{>ah0}d��ʀ���V���	��I�"�w9�
�w=.��vSGL`u�P��1Í�t�����u�6$բz�]��JU�+JװT�.E��%�2�{1}x����K�Y��b�9����g�f��#��6�k����M��*�ħ�M>�+���Aݨ���2���T�5�f4Xgc&3���x���ξ�mC'��yP�xdw��p\�˹y,/ʆ���Y�/V���`���/��랐'9ԥ�KB	}L��3Y�q�sޮɈj�AI%�!r>x�l	������'s�&aBK�m��Km9,�ٸF�Qr�h,� �RK �tco�8D��x�~�-�����	h��9�ọ�C���	��-�uv9�.�1aZ���V�=rJzM7fE��^��O� �Ǎ����$=Šǥ��Y�֥�U1�y<���^ˉ縝n~�����uLB�֫fg�Ψ6�5�{�K�%��r��o&�␘���y�=���=zPa���KA�r�kG11�筈���S7Y�A�jq�eyb;\۴&÷���no8�A��;�X�o�E;���%�Eǧ�U��y���3;EtFD�c�k'D��R�{R��I������
����;�
N��	~]�*���d�b�)�!֎��:ˢ4s��Q,��)�W�F�]�m�5s�:y�}>&J�.̀W����)i=�:m����-8O�J/C�%:O�1�X]"��Mm`G\�P|��\��l+T+@����Y��42�R��'�k�e�)%C�ҥ'�I�WU�9�z1���,Ŧw���������L#��DsmN��Λj/`�i.j{F-9I�� �?��1�JƆ�̧�)|�b��M1�15��@�t�f��Ȕ�z�V�D�۴/1��Ie(��2��8f2l/��1�+��v�dJ�;&T+����!ivW.��[l��+8��	�ĢGn��:j�}�=�e���jSa�m��Owu2���� �2�-���9#ϑ̹�O\�u�g*ּ0��^W�^^��y~���]pY¢�j�{�\a�'�qҢ]�:1�� ���7s�2~=�=B��ɑLH��"fo�W�E�؅����#<_��6�a\���l��n��;�!�����ͮ��d��pcf�U\�Y�ծ���4/�:��q��1L�������`��5�3�C�C�S�j���H[�0�T��x���:�G��Bؗ��Ͻ�C�4��l��
$@�b���rŨ0p]1�1�KR��yͭ�C�JL���<q��|뇦k���Ub���c��o�خJ<
����-=�o.�]ܮ��g��elT����AVծ�)��N6ۜ�ޟ^Y�i��O;bf�sٗ�������k���t'�X�Gz��m�Vȧ|� �����5s��͊֗��e	��s1��=wV��>dF�椲Pj�#8�Y��� [:y�x����y��L�F�vea���̎�]ց���e䠄��vi����]Z�F>6K�9ˀ��(|�9�ϸǕ~��d�fY�nQ���R�}��f-ʏFL�l�>6W�}�z�=�Ҳ�4˳�3ev_))�4�zf���tͱ���kY�J��Y']�m�k����F�Kȍ��c���+r�Pw��+��Ľ��V.���;��k\J0�aZ�l���̛'�����3�LN;wF�6��<�:!Z�9E'W�P�r�����8�:���	ᵫ��V�*c���:!7�ll�\3�v�{,�$�L[��$�b%:���j��e�U�ҨVd<estmS������8ޏHB1���Dlʽ},�4�v��I�g	�u:x՜g�Ǚ�Y�\;k8���G!�3e��-��{m�� ��\C#㊡�Y���x�I�T��𱳢�7��	�b]q�kZ�sӿ3��p���'ؑ37s؞�ND�:�S��؃1�y��ۧ��^]\¨Z��B��/6
�Ƒچû4̵b����_�
�=3��+��Ѽ�.�m�8�5k�'"��G,be
�W��]<�o��=�(�`~jǷ�7>��i��"�q��l��р�W�z�c@u4�m�2)s�X㭗Jײ���R��V؝i��{B��t������@`�Dy���z�6׶���zKר��v&�K�E�E�fȞ��Y7��扫��͍|��ׂ{�L�w�\=h����߬	�vI��;wx�Q`|���=�P~���jڳ~kz����Tdh��ɶ���395H�+��$��Wbж�v��z	�U�"RW�֬#����Xg�v��Jd�=�".�����8���Y�a�������t�3������\�ƍ�jgf�̎�Iv?;��A��-U�n�򻺰�p�s�)��L�n=f]�lhtg/#^]�."�	���/�/ѷ8��Fbv8œw�[;�;���C��C�J3˩��ze�lM�1��̀��B,�7IIM��u�+s_�Od)����Z׋�Qb_/W=�B#^k|�M��.WE3��K�M�ecR�ӽXa!���]����jS�R��;���`� ʭe
)I��¶=]&	���p������(\S?���[D8�v�vq���R��:��c��ʭ*����9J�a�{��ݽzFf�c�M<6�\c;@B��S�I�逖����6�uIj~"S-iǮS�^��G&�mw����`Z�"�]�Nc���xOB��Hqm	��/ ��| ��z%\B���j��th�����3\��,��n�c@i0ny��s	���� �6H�L<A��Z��mgZ;ݫC	�R��1I��Qu��c^�����\�0l}p�ϘF��%�9�ͽ�"�Qf�^��%�����'N҇Bʮ��j-?5�%�.��Iĸy�x�J,�.�~n������W}�:!ΦY��@ps-�5,��m�`0)1�AU�u(�{�f���l�eĻ��s�e�Xg���z��:5d���I�τ<������Ar�@�rN;��l3�(��/�uQ*YZLa-�n�ۃF��_K�\����TQ˼��LU�V�Y�شƈ�5;4]X�6��'(]�Ta���y�ʩ�CP�a�ouq��4,�%�����0@B5���8s����j��-l�BU�(r�Z���g�[2�t�{��ڶ^�׍�1��m΋`� t�@��ʊ�Ի�}>hi�����/y���MЦ�B"��e��h�ݦؠ�6�,����3<�n�����A������u𹦷Y�T�.q�iKT~=�p{ܚߑ��6�������"e�D[���z%�r��VN\�c�=K[,��C�"nO=��k��h9��X�F�$={�@"x�;O��􍈨~��v����U?T��l���ք,F4��B�,?Z��U�*s��׸�|*~�d!�������V/aC�n�i͉17|�g�
?x�U��ê�y~�,�ɯG=lE��J����A��_<���r�e�z�8�d
YA�b��=[���N�[P���ǧ�M��	XQ^3|�7�|i�t^��(��i�����ZSI�WN0�ј��z����;��e��as�H{����߿gg_���L�C3�@JF��#�]��gw�WU��&Ƨ�vjW��݅�ӧ�_����Xfq�͢9���px��]@�rrc*R86L5u�PKT�#]F%fq��2�Ê��&��ۉ��X����S�(�ɇt��,��w������韀�9���7�Q폁{�(��q^�Y�B`��̔�M\":���<�ۼH03S7�Hh�ev$՝�y�9��j^�z$p��$����>)Յ�)�xi5�����h�p�kK��1��#Z*�\�=����#a����c�vHeC�'%C���T��"���n�K�k�ɱ�(��bL�Œ�_ϫ�"�G�B=D&���ݣ:m���S>�M��zO�2��]=���p=�Xj���tQi���?c�|���;.,FĲ�O\���ʭk��ㅷ�n��h��L� H��z�Q����H1.���q����ٓ��'�W:����qtzT��Fi�C[�nU��R��X�d����*�#&��$z�P�O�{�[�rg����,ѹ8�5�cŻ�Ŝ�Ze	�s�X�.�VߍEsP/���!ۤt0g�_Z!Co\��N�t�RΨFg�Z��mOC���2��.923L	:���j/��]��c���;K��m�C�R��Dc;Κ�`�����#u\�־ԋ�kR6�)��ܵvn��ݖYr������z�wd��	{�u��m8w�B�۱}):����l��IY��_V/��ڈL�mģT�Ul�ǵb��46JX��g\W��_U�d�9�2���Z�o[,w3�޼���0��銮"��F�u�6o^�e΋�#N�l3���ݻ�;�{i�;���1:���uk�<]���b^T�i2*�p��f�����;6���Ϩ]���m�����ږ�}րn��S{���Sة�C��bwB�%�C���;n�-�5���q�!�wgQ�N�%I�~�\2�%��C,<p��.��Q��b�̫,%g��&Pu9t�:Y7ph	_sO3\���\������.�=j�-���LKH�q�o5ж-$k�}(��X^�q��)����(�(�;��й�kCN-*�v�
��X�o��h
�Ƣ:2]n�z��O1_7t� ��%SxJ��m."E����r�E��7��D�'���)o+�F����9�h��aO���5��L��:ٙ[#�_�0��JĹq�;�;8�x���O���a^���َ덐���X�f�7r�ps;��>�R�u��n��<.�ΝE�gv���x����>���5
*��.g��Ѥ�	H��3~r��2:�c/�M]��Q�9Mn�첩S��u�,�â�*��芥{[ut9:8�q�&�E�v03��J�9Y�Va�X,�cp�s�ٌ�rn=�9Ҹd������a2�:{��U�m�)WQ9����%Z:�U��6©�p�a���P��l%�#����&�$.�v��+�g��4��8v����t�|�8,&�`!�]������Q}��39$��Rɽ��Ӯ�922�j�Z�Ii�a1:�벁%W<gvLêRCV7JT�ZKpE���w��0W�W4�έ��[��j�u��B<�Pu�u�8��X�7v]l��k�NR.�W|H�+�}�,v�{��e�&՜���Ҵ�lk�㙅�K���0TF�s$Z��v�y[Ì��/��͛,�	n�nu�nr�bR��ޥ��K�y*&;��;�XU^1�j�8�|/�L"�za��	U�Д�B��ݘ�wk�: �D�.c��=�6^om��p�y���\�u��uJ��x��[1��갂U����Vx��S����I�*�eE�����mZPo[ щ���b/yf�4��r����{m(_j����nEv��>}��N�xD� �jR���M�
�Nge>�zf��4���\����NC��t�-���s�ޒz�-�̆�[ss��S�q�J�>���*�>�Y��1�m:���j�ϙz#�p�K��*b��� .��̄���HrtB�{.g,ߤԭ�'5)��O��j�
��({1\��Ы��w�v�" ��p���Oo�N/fs�E��G|7/s������]ϰ�y��^t8�062 �r����˘F�����ɭ��Z�
�rr�ebub�v�'�a<CsZ��7�6L�қ� �]S�Vɳ!C_|�G�@}c�������9%I�Z�ە�ܚ3,��⫕l_���\�������Z�m*1ch�\��6�W+����j5�v�ƹ�;���m\��Alk����s��k���9LI˚�5�����ۡb��1b��;��ɪ涹m�r�gv��:vۚ���V-���ʹ��rۥsF�r�nkct�r�6,ms��}@�Q'�߾yJP#Xd ߦU��m�:�m�ד���.C��1�Ł�C[�s��J�3�y����	v��q-���6�r��ڇ_NB��'j쥦�ƈ4
����5�ٙr�\�x�����X%1�k��Qќ���ک~�H 4\sLL$����m����zC�f�F�Bsu
���F���3N��Ӎ��0�MmI��m�����(>0���E��W>��ԕ���"����mK��q,��!�,��W6���=��T2���z�����{GI*�+;�zںF)���;#v�noZ��!?5�0�z�X�^��Y����V�9�>ڷ��Oi��Z,���N1LN�H�Y5�\���L�˜��tq*�Ҩ����'vFƥn:q�&�b����Y�����!����5d�$�B�Y�H�Ź�2O�1�w�(�i[BYw�:��WDp����m�/���-��N7�HB1�C�H�C*��b}|e�|R��4i�R!s��D�us�vr��7H�z�4�l� ���qń�i�9	���1C	e��H�p�.FggA:��vj���QO��Y��9�4�m�\���ρ�� �k؇!��H�����c����u�ܻ_��D�&^�+��B/$(���\�FQ *�G4pj��xW���뛖��_�=����J��`
�]ZI�"m�H�G.���o�<N��XE,^�Ejҭ�ɕ��t'~�PۣoE�U��� +��rÜ=.�ŧ�ͥ�٤ ��w�^��  �Ƹ��t�)���Iџ���{h'�e�T��YyCB�v�i%|Ts��nU�_�;�Bz���~�7B͹��.�TXU��c*�Xi{���=�v��w����i�y쥨0jMi��L�_����͵��B��Ԭq�t�{*	{e/��u�#�Vms��R�ދ�a�$�!��i���0��Գ-Β����*
���U��nv���VI�m���ܝ��J��W�@��3�2%�=¼dD��3����r]�u��/��wfԥ�}oɻo.�3O=ܭ�]��䥘��d:�ұ�5��,������x�FS���+I��.�Y���o|u�{{V;a�v
�-�d���H���p=2�xc��`0'gs��@����y~��<�t&���65���}s�P���7n��b���sϬ�ag�D��=X����09�軚O��ەR�ǔ��aUk(Q��뇍Αg&���vJͧs_W����y�߼zw����4�5����C��i�g+کnj�"Sm�)�$>��UU�U5����݋���+^\�K�u�cռ4����1m 'C�L��W�i�S̼�ͺƎ`��dY�0��*��*��J~������g���Y�J��VV	��#ڇZ�qܝ5�s��=�tn��Cc��aaa���=�7$�0d)�g�M��82���_��ວeӺ��׳�z�I�H5M�ܼ$ۻq,�`�.�wpR�1��Nd)(�B�S�����rW�����]�׿o�	�Њ�w�9�Z��	����C�h:A�z^�\��N������������x��θ�d]g���׊4�P�\ᮢ�ch�a�hu/8�X�ن�e��i��aY�+�4�"x�}b��ʥX9�ױu;uNY�6����qE�WpњFl��d�o��c ��R$����U�]B�Z~k(,h.���ӎ��q�rR�ᗃn�B�<S��<�<`0~mi�5��;4�X�6��'(]��Q��Q��BU�UK�y�����'��D�i��Bq��Ҟ�<� #Xt��8u�ѱ-�g����J��?V��X�w6�[��ݼf��Kܽ�q�>Wrʹ:-����:��]����6���!�K0��zY�:��+�v�������ӏ^&g������0�:!.��b��q�r`��3���.����7�K���=$= vQ1^>��"صu�v �D��2x7k��fg���t��K	4�D����f�X8�s�8� ���8�'�S�m��7�Uv:T.2�$�6e�Q�M�r��ʸ_F�	�2Vg����݌�Ś������X�<��x��{Q5}k^:N�͸�WTYh\��s���GMw��@�� x�f���;̖����wg3��B�'R���zħ�"N���h���iF�fҝz�n�̬�Z�?��)O��LԴ0�X�T��'�=�gzF�f�i�ø%��f��BvZ����uf�7y[�u��颞Ƽ��t��P���\���y�b-�.J��vFoU')��U�^^V�ל�5-3�5�Ĝ���i���W�E;�a6�,:/1q��@�	q��H!s�3D5ջ�7ܼ��ͷ�MV��{�ӌ+ǣ1��l;�x�_=�������Z��ۖ��[_z�!Ѿ���MsWD�P�Ƚ�R�eaQ��`Dm�5s�:y��v�AO-,���j��k����p�̝�.�N��%�Xuz�HB@�_�a�%:O�fi=Z�Ɗ4����Q�}7Q-�ZeZ���5�Sm�|���_�}�� ��=4�~���0D�pzT��b)9X�R��(�{g��Ϋ��k����XK 7b��|�>��pB=Ȅ�Sd^�5��a����&YK�c��[�{�Q��#��fs@<�RiK���d��a�����5�����N�M��Rꟼi*�-��MTj��N�s�Kb��P5�?x��zO���vosc;
l����!�?�}�o�*k��=��ۭ� x�"�i"���g�J]Vx�`T�p9Wp��o��f��6L�XR:�V�<�����k��m�5j��\���{L`#�𱋏��.=�s0�����i�f(xT��ǘ�xp�
�u���vmi�Ϋ���s&�'��&��Y��t��{�sY|�����*L�n�	U��Lkb�y530�kb�ٶv3���x��u;Xۊk��t!۞
���r}cMP�~u)�S�X�˧զ^y���B�)g�I�*�3?O������ `�ɝ���mo���_e�2��C#4;(��g�%�6�
�i����g��ø�����сAi���oӲ5���A��u	��h�4�qE�bb�mm�vVQ��3c��d�O\�o��P�x�� �q� D�N�zq����������yc\��|�[����f���;�6�F]���׹���	U��M�����c���Lvhx��q�Ӣ�wZ��kP[	㐃��!���=�8ʲ���zw�X00FPx�TP����u61!O��v�y`�P7�ʊ�zЂ~k��P%�$k�]�����x�����tU��e��گf�fq�-Š&'��wN˦|�\��,}��>%B�)��O5vg����j�f��Qp���Dkzf� $�"�Y�Od�殈L��1�Gz=wV�&�	��j�;^�X�iF�Q@�>��.�Œ��׹g�{��i�ܣ�{!C<M��*���ehz(��9�6��l
ƻN�	��[˻8��π<Ա�L�3qV��S]�R��v�gH���gR0�]�Nf��,��dWcK弐:�B�G�7��	�*�8��t�	�d[B�t�z$��q1�C*��CH�2�N��ss76��|x��|���Ʒ�$�+�����|��7  ��\9	�����e�V	lx��z�¯������i�R���d]axӋ�F�ٮz���.ڽ(@Z�����Ae1�[�]1=j�W:�O�=t(~�I�U�\�֪y䤱�v����vh܇��La�������w���ܢmOS�\�ě�e�q[�U�9��u�$���i�2_z��-�eI�á.3��S�Y4�0�О�ʹq�jéX��X��Tdf�Z|�������k�C����=�s#�0~�g�#c�D�潵,�k��XsV��N�4���b������SNyݢ�K�t��z�^�9��~CΈL!�6߬NK�N��(/�C���R���gw'mC�V��TIx��&��� L˴�tE���l��^]�dh�/�aGd膷����1�.���r�{z]�[�$i�Hz	@A��K��l�tM�1��͞��?�{���b�sf���q��-|�kU%ױa<���\r[���Xe(�2�kf�맳F���ʵ�T�������X��R:��t����S���M"������ݚ�'c��r��F��H�m������JۜdSt�3Y}$�ވ�˝Ap�:�%�fN霕��L�y�e�4�T���l�{����^=��ƴ��	-W�G=%roW��H��tս�1��t�x�=�Ο�gQ��P�\)U��+�<młu�le��8��Z�r����F�N���Y�ʹá�q���9��L�9lk�0Za�s��l�%�0�����M���+���9]s��o����&D�=�.�N��,k�<4�|gh���S�	���}^!��;,��7�r�P���̺4O2��)�P�&"T.�'1���������-;<�VEl���Z)v��4!eW��Ʃ[��YX�ƁF�
��W8�˘O���oxQ.�U=5:�?�m��[���ג�}�V׶��Z9�����s�)�{6F�F�7X�SQ[���*�Ψ�8��N��.
�H�#��zAc��I�v�8���]B�Z~k*lk,���.��05MS��x��%�q.�-@}�0�t�ZDp�n�N�W&m�jw�lfE_���Ȗ(�=�=�N�*+�N���H:��b����hA��[�G�:�����j�=E��y�4ܡª~h�J��{=�+5��ɋ[��&�Ӹm~�t��ʫl?r�����OI��q��hMK�v�U�E;q�yq;�(���Z�<�*�j�3L�c�'�)u�EJҵ3eAiV�!�fV�ث=�i��ۯ\�䣄ǽ��	s3�N��\��H��
�����{�PKܽ�Q�*�Y��E�~�����@x���C��f���N���"���U����5��)�BT��eO�)���3<�<w%�ы�d�l���4���l���n�G>0e��q�{چ�����~�Ǥ�$8��b�>:"صu�v/y��	Μ��-��T����L��~���}=6^�c5��3��;Ӭ#{��,F�l�,�ؑQ3��ƞn�E)y{�d�De���:�vU��|y-v�m˛*���;[�(ү�= �|��ο�����tfQ��&���eBe��7�eq����{;[�CO�h�m	i͵74�oi�`9��rAPw�{��^͗~�]qѢ�{_���))��H)��;KOfO�i̊�AZ�݇q�
z��{�v�$ص��+�$\v� V�JP��x�ʹ�n�{rl��gR�bp<n �f��Llho\�}J��Ga3�	�N�<
*��N�k���j�S&ClI�(c랡�m�+4���I�b7~<<W����h83��X@Иa��V�劂���UD��df:Ps�B�gwE(�
�t����ʜ�ʛԢ<ȴܓ2���l�޶Ա�U���Ҷ��/ag0&�g8>��[�5��d[��^���l�~��m��]V�)��_���=).h\ky�v9�}�úl�5����W��-��,-�B�9v[�`
ޓB�3��Ә������G5�7��ܱ92/g�W�R�[}j��<��9���U:V~©Tk�B�L	�ѺA�ʫ'�h�1Ew.��0�� !�����߷݂^u�w؋������-�&�Urn���-wTQ�
�d�m0��x�T!�zΟ[/e�%�9����z�k7�q����J��������[f��퍼9M���C���n�t����}>`pc@��B�U�I��6Q���D�˕
Y�E���;z�Z��{n�V���h��h�ά�H�7@�}Xvb�Q�����~3�q�P=ͪp�A�G�\��g�h������;)ڥ��!�j�c�gw%�DO�������������l����B�y��n��ld�E[uo=z͗��k��)iR��j��ۮ	u�d�&��B�o�U}��)���|��5����@I��ٹl����5��#�&*�#��u��.��r��ݫpd�|�o]8ų�D3�����լ��1��J�b�3���%��X�a���*�&J^�E|w՛ߺ���u��H�@�J�K���ԋ@[��Z�!�d*P��Rڴ<�V��Cr��x���ǈ[^� �&�]� ��F\f��d���i�"ok�u��g������5��y�Y\�L�̜���&���4��޵��{�f���x�  ��BB+G���\��,�n�k��s\�s�i5�=�P}�=��}ِ$�����<�����Țs��:�y���Y"�t�+�S�t�Ӛ��A���[!骦^�����ü6�{G5�'T����Q�U.7κF.m�=-��S=Ų��}V��+"����\j���&���_%U�+�C�q�H	g�Z��'t����yu\KD��i,+=�A�q�<�A�4箨w.Uk��yV��˩8�z��>^�ym[��0�>4{EzO�]G��r����3e��a�^�-Y�a�-�6r�˦Ye�.�˻�i�>n��y���I�WO���K�0����T���UZW�7�$w�q��:��n�;s�Mu�/%�Dy%�vǦѽ�R�S�o^���q�̩su�Wx��I�:�peنڻ;�k��[d�_:/Q�]�)�Cլܫ; ����Va���*��;�^ݸ<j�1�U씮�?W2�x��5���Jjx����<+;���n1x1�ߞ�*�k�z�ue�X��L�@�[�S6j�?�x@����b��;���2�S�4R����̆�E�Y|"����ס��6/hܕ��ѵ���BS�D����.w|�Yt���#y1�rΦᙛX�v��.��f�����9B��$d:k:��·mml�	U�Y����leu��U�K��-Ӎ�|�����T�b�{+Fzg>6������ʋ
q�K+8�t���(�odڕ>�sT�Tך���ô�� !ή�Cv��y���BsW�,�y��!�'k&��X��+mwWL��1&��VN磯W���}&���j휍��7YB�\�U�m|1K�p��AY�+Ab|��瓱�w�ɥ�;j��!�k�@�E4�vDx�b�DW���q��n�,=���OV��g�vJ��P[]w�76�<tV���Z��r"��ts��a�Ƽ`fA]�,Җ�>������1F����D�a�ݾ���nm���>8�Lo�s�ʕ�e�h�ǃծ�ht�TO,�R��y2\ܳ#;�:��L��J!'fU�/5epI�[D3,TB���w����V�w�V@����}�a�*1C�R^8��<�#�D��x�_��r����u�I��Ǽ�H3��[�*U����·j�	��v5]0�]���q�7��[Z��V��P�E�K�y�%�� ��Y�մ%.��e��X���U�e��.K���j� �غ��B�����<a	����Շ�{��2_9C2(b
���s)��L�w}�Kʗ�*zq���[/��:^�Ѧ��a��9q5�ĨK�mmf3��Z�ˬJ���ֱ�2��X1}m�vM�	Do(�}����Xj���45v���;*B*��]�Ṋu��ܗ�V#YG^%��ޢ�8#vy!5��]��s7*�8Y�.�s*��$=]��>}� 3�ѧc�;^�Y��j�!͓+��Ư�/k�s��\w���]Ջ1*ŕo�j�]�7�_��tF�wp?x����4+�j���#�{���چH+�jǦj�Ѱ`���ǰ��ԣZ��2���;�sww:-V֮�$�Ԯ�����WW*�G��e�E����ڊ�l�H⾓!ol^Q��ح���W	qD��e��?YYdWMPn���fgҳ"n�*}��[Y$�էM�O���sn�^Ԛ;��E�0��:�&�<�CyH�:z4��sLK�yO�]��]Qgݛ��B�;\Ge��]�\��׫4V�j���պ2'Fov5s���~zأ��[�k� +���F����]݌l:��Wwj��+�%b�7]ܝݔn9�����G8s6���s��vEѲQF�9\���H�;�s���9��Q�r��6���1���r9�뺤�Ě(2I�n�s�w%9�5�;���c$��ƍ&� ��Ʌ�f��$��A�ňI�\�u]�I%�w5ˑi��9���Er����.�
��~/�|�?>y��~~��O&;%��X����ǎ[�q�`#ݻ#`·�%Ak���N�Ou�v���)�#X��X�)�o��v�I�߁�����І�F�Bɽ&l�)=v6~�T�)zI��-=S��wF��:l1��g��y�o�'hrm��M���l�y�U��Q��g��%N���**����c�z�l������4U~�-�璌�*���זDi$jI	�8%s˛��8D����ߪoMbd$T@ж�U����nǯ5�l�h���MzDYiN�(�����Q=��|�E>ϺY�cU���z&��.V��Π�{5���Y��A�T\ܞW&m��쳄ǬA�?G�����jZ-Yf~:b�^Q}s��4��׭)Y��.��ˉ}��p��$��BB�e硚U�!d��EW8�D!����A<���%*�"��.��u>l�:ŷq'_�3�j��fM蕘LC�]УE�`���2���*�l�7)�{���)�3.��9�X�	�����EyY�*Y���˶A�'$6��P�S��G����J�t[���Gd-�*�f�f�åGʷ�c{8�F۽��X���#�\э�Y}��I��zz�Ћ�L���#���L�����C��Z�'g�נ`�W� Ȳ!O��J�r�U�y2-km�a��溅<���y�b;.&�)�A>��v}�p���O3EkυuU��Z�ŝ;��"�ӻ՝�h�~�. m�_8`��ޑ%?I;��t�����ڥٯ�#�-އ#������ ������LÏ��X+zDl�%�8z��[��ݙ��ؗ�=ռC�Z��≨�+M@��O��n�G�R��ϛUZ��NF�鍫�J���l2��峔	�^����1���s�{�-y�����{)�R��֫1z�>��<A	��g��6tT���)>�rk�=m�O�������_����yf$i$I,CD�)�I����՝��ƌ��~�d3���siW��w��Q�f�˱
����M�����!ݚ$��t����e��A({�/ޏ���T�~�<�婿�eX�\�/6�frF�Z׍L=�w t�|��ƥ��Yݮ͙��qX2�=W�ŉygd�ј�#tY�d���NE�4�U/�麴aٍ�;S�Y��.s�	���;��f�H��N����UEV�X�l��P63!��|{�9�u� H4�ԟ���G3FѤ�4�6���l5X7M�[-3�,�_E�sN�R�XB5�k&6}�B��R#&��=�74�E[(�[G#��(�l�����D`��#4@]�O�\��@�J4
R�)�T<�W�e�q�<F�a�;S�/�N�1����d��VJ��Ga:Ηk?wb��Q�[�m���}X�4>���/�e���j@B��1���Q��JJ�m�N�M�E�w�7YE�t�h�:��WQ6g��d0�E�!��Nȍ��/�Mݾ>8}������:��Vl"�r���6�ʐy�Y��<����#o�OA�]w}�u]i���=Q9d��~��
�]��a��6B�Sh$��{�ʻ�΋6b�	�h�v�kђz�r�NM��-�k���%R2���j�c-ɐ���G�g�tw�P��S�b9�/L�J�c�(rQ������z�o�>r���^\��S�(�׼{r�)nAf[ڌ�)S���i&0�z'�-����R7��w���YGV�v;�� h�*Ԥ��_{2R���� ��3�td��	��w<��v��ր��ܢ�]v�/罷̛�Ǔ�Vk6��'���fN�-,n��sf��Ί	]��7�LB,v��e�lvٲ���ΡQ��B����Z�u5}�.I1�=�΁4@�g�����<+4#'�R��;�]�1k{��_�˦w�鲶�����@: Ϻ)̌�th����[�qj�9�3j��WGi����>�VnX��xJVD�i�Yj�E��j�a��n��ٌ��j���hh�׆�&��͍�ԁ��+"R�i������ٮ�Ӓ���u����2�Y����r�D�42b����4T�K��o;f���ǳ6uۮ�F��4���&�բ�+�������<���%�Wv9���N��Om�ɽ�"��ٓ�y����PE�B�[�=���2������*�����4�gPOԒR�P��*=eHYa��B�ڣ&2\�c�k�Ak��r�q�M��V��+����T�s F~��؎�P��N�t�_��Q���cg�1�]����E 5�<��ǔ9��e�^f2xێ5-ʺ��EZ#�lT�o1����K�\�H��Q�/��f��]��g��<|^K��9�%�'ok-ԣ���eս�q�#��(g2��7���M4�������
;>��?k�Oe-P��tdb��g�0ǈ��3�Dh�����dcPZ�:d�l�v䪅��JQԻ��yԊ�:|Wa�W�n�)�p�rv�z6R���g��w.Uk���ʅ'<[Gxe�oWoBAu��#zvt�3�g\+;�K�4�T�1�s�s��ѝ�^��vRUˤm���7ͣ��އ����Ė��Ŝ+����rGx�.���/��,5j�,�&q��)ܵD�3FDp�|���e��^a�[�^;���"I���]#M���r��s���a�Fe�{QP�zՁy���tz��ΒF���Lય�3al�dUF��a�E�r:!3��RR#k+�gl^"k��$suQ'�Lq<-��iسW��)���!E<���J�K����yj+��γ -UC���L�1���UT�E����m���J���K(��˻~��I�w�SpW0y�?; ���/I;��*V8g�����%��F��M��jkΫ���\��݅�X�3K*�L�5u�s�f����H;�N�s:LؗM6��8�"s+K���r�����gt*�6�%n#E�2��ɷ�wn���f���{�u��⒫JUB�;U1.r��q咱��:�]&�NFV�N>�њ�x��A���-N��%*�US���+��9�ڶyط���;���N��{���5��gL��1oB8�x��?�[���`����+���>V�����]�˶�x+!O�:IV*EX瓞Y1���U�_l���>�g�Bk��v�}��:�Ք�(�y���e��X3�8�̱ǩ��f�������j2�u���.�=�!���K�&��M�k1�N�n�����۝�d�y������i��3��a�����N�S���&�N��>Ő�W���≨�Nf�W�o�T U�n��^׷?$BX�yQ�I�ۗ�'\���7@�%�A��g�����M�u���T�I	��k�a�p �����fVP�!�^�[:]-w4��C�G���80�!�����u�ځ� �턼�C��2��wf�*��R�4�#Ȟ
s������:p
�Q��ani��v� WB�N�d�+�h]&;���5w�N;\\z�[&�B���3s�ų�*� ��}��z�ǤՒ�h�u��j��u�y��U���w�αuR�P��y�Ҭ�n�@f���f$$���[8"pm�x�wq�$�s^v���JF�M��k��t+��$�Y&���e)�lx������;���BG"�WJF�9��X�APT�����0L5�-�f��ۓL廜#H�d�QU�t!��:8ӛjE�(e���+��V�ݰ�A~��G�Jn��q����o�$�R�'i���0��5�ObO�f}ޥ2e���;#+�#8Gv�g�����R���a�l�L��U���m��ԭ��\"�^��b85�5�x$�8%멨�-S��v�W8S�.ʠ�:�ԍ/�\y�3�𕽅��C�X��^�dJ۝9���6ɞ:��M�����pC��Ï�����j�d֧����w4��^cGd�|��fE�KTS�Sï��ͣƹ�ηי]�EI+N��	���r�nR�AI��t��tA�})b��NGMv��7�q.=%�ʖ)�����em��8��S�5�t;J+ӈ�#3����s�{�T�Mɂʏ���EI��<QIE)ZKfzζO�J���-�3U���zjLI������}�����k�H��>��`�mu���Զ�7o4�i�%��7:j9QbjsJR)n�W�(UC'l��v���G/q��*��`Dy��V�!��*�Ҡ䮯2Օ�]�i��������ݻ��7��z沁F���H~�v;;^���&���2lGݽ	�nHJ8��y�tt`fh�!�3��I&{��m"M^cNt�w{�}�V�ֽ<7�V�L��A�fz���0_/�8�D&�����]q]q|*z�⼲#=�� %�g������&z\da
6�Տ'{,�tI�DP����M͋Ųu h�BVD��+)@�.2���Դ���.�-r�Y�k���S�{rb�.Kk݄����:
�0��DL�.�E_Xr>��hY%�;G5<7儌�g �8I)]*eG�j��@���\"\�n�z��&T��S;e^��u^�a��H˛Nn�����_Ws��y9Q�k��cP0Ѿ%������A���m�p !Ռ��IM%��.�i���?r�_�5� n,A�~-i�4�X�9Bg�3X�v�{�������;Qڪ��Ήx�����.D$ V�}.�6껍�M��w��u��<%A$����jF废vdHY :Bꮚ�Nv��#��o��۱����3��̓x���\e��<ǁ~�˞��;_�n���o�{K�g�/�����a-P���F|1sl��N7�.j%��&��S��>��#/ú}L٩��U��+=K���-�lo6r����9�ֹ�ޗHt0t�!�?�m;�#d��Fl�����a`Ǟ���l�z;�<�����~���7�uz1�Vq�LoI���m�y7����v���7���W�\�Fߺ��}���b�P�M�V�;�m�6v㻅����$�2�OY� sa�l1�8�w�F���@��7I=�S�@�F�����]����U�ư�Q�V&+���-Z�h��[ۀ�����J�c�$�����e��̷<]� �dv�8͎:�8���HF\��[Z�r�#.m�'nl��v�����Ю���J��u�m��ST��9Gjq@�|"���F����k��$�nI����9���r�{V�4l�'x���ip�<m*��F���,Ɠ����r���<�r�ͩ��S�7m�$Y������:#�YjJ��ǡ�7�W�Y�t��
y\�����x����S����J���(�ٝyO�I���ܗ���c#8JuO�M/�9lM���\��iQĺ�|/-M�9��!N(#��Zc�Y�8�6a
�펞�>�A�)"-)U�|v�ji�ճ�mGt����y��Mr"Nq���Y����ð�2	{T#\JN��|���ɞ��⫍$f��c8�=1�<7��	Gg�C���"E���)"Ώb��q⚤�����oܙ�n����0pE7%�'x)�i��:IWʑO��{M�Օd��7�:���^���a�8A�pY1����v�6�2:��.�����r�˗.r�ه¯c&�Q�5Lt��P�#yZp����!]�:<�8[����י����W	�3��S�4)Z#������'v靷Kv����e�Rɻ��5kj�}tۛD�\�:�K��b����V 6]=�C�uM��0�Dޢ�L����R�@�M�RNȯ,���5}�>�Z���\��:�1�!84�e\PMҪ�Y�u�UF�^åZ�tz�P�E�M�K��xR0D�9ӮP�k3�
&'=��(G1��X���8 -�
Z%F�#X�9��]6�gë����̢(�J��Ƕ�Ƨ)U�xV��}q�M��:�f��G�C�-�����ݸ��*fZ���m��ֱ���i�Q��d�ί�RN�[PJ'o��n�9:�Cj�~���F�p�V�o��Wt����LEy�._G]i�O>��i
�h�������u}�Z�]`Lš�&jIg2F�L�9���F��ͥ�נ^�y6�k��̌_q�p��&���Z9�Տ�Ŋ�W�z���ZZB�����w �Η�٥Xi�I��i���R����Ӥ��C�hc$SB_7D�Ꭼ�)�z�C�ec&u�smT��p%@��r�J��2h��݅�q��
t�WV�.�]���+)��+O<�R����Aj��3}��3��>r��s��Pw���n��w��>��PY@hC�`7��&^��)G��V!��܇jcÒ:je)���:��5���+`����� P�����u�S�Z��G����j�(YtbŻ�l�2��Lڰ��n;Ӧ�V��M�9�6�<�oU�BTF�Vr�'ZP�z��r�e���7�5E�l��F��n�!�IJzVɔ3A���q�7Z�+�.�i������{Q��;{��s��t�Ӹ�16j�(otc#�O2Ь;�6��PЙ��'f���|_YX:j̈u����+4k&�(U�/S�+wR������Z��3q�����ʉ��3�٭�)��[X��xw2)+��英f�IQ��m]�]��[9ٺ��:[4�VVu:�5���=3wa��B޹��ǝr��r�Hi��ɋU۫���\�,�En��<���4Wr6r��S��8yMUΞ�ʻ��@|��*�,i��Et����� d���a@�l�S#/Q)P�4p�v���iRs'*W�c�� }k���+z񳵍��[�?��7_R�
�Ȟ6Fep�Z:�39v_Ky�*���
��f�>8gAL���s��t���j�9p�q+P����/���ڑ�\��M�g;m��=t�_t<����4mPa�	��WK-�=�B�_�U�6q�{�ԫF����ч3�]�4�N�ݱ �2��)v�4Ұ,M��o�7l|�q�v�z�;ԡ����c�V!���ͥ�0���R��<�������iU�/^���oĆ�t�)�TŶ����NY�0�t�머��,�&�w�я{I�R��|dN���Oks)]j���?�O��"����"��76�"�s�I T�p��˘,cD����s��r�DREs;�1 �\��t��I3���ݮ]z�*������<�3D���Fd��M�ٔ+30\�D��QL��y�a��ġ�(���P�BJ�2odx�A��4QF.�w"%$�Lr���`d!�.��Q�y۩�FLg�]����y��wr$�È�y�bD�$B� ����c#hE 
���W����Q�.��46Wѽ�$�Lܞ6C�l��G�%���u�S��/Nj��]��c�QR�J[�V�j�c����(g�>����bO��ˡO�]�>�KB�%$"��B�lv4𮱯�;����}]��&W�F\�>��C���|���+%s7�������ٽ�R�ʤ�y��|	ݓk���gCzo]a���	[,�Us���*}V��|���ZR�QBS��y)���0x=/J�i͗�]S���x���ܑ{ԩ��n�u��r�������`�ɟ�R)O�3�)U�~��!`�`>��+K��z��D�Ɖr�Xը[��5�W�ګ�b
�>�9р�uf��Vklz��!��!+\U�-%�L2�ί�y#�Uߵ���v�}�!e�%����DT����w]�M��A��ܻ�X���h�])ا9B�D ������+":&��״�\^0��>�Sw�x��=hu����l�Yt��(k捫�/C8��5�Z���q�aY��B��SJ:I�G�ϫ�sD\׺�?�;Zri�뾋e���ZJ�)�L��!5���(��[�L��8�$I�U�5]�5;]%z�͝O8�;%��{][������*P�҈ �摺6���=z�t�˵����r;PiVQ샷K�Z�λ|ʧۇ�mb��@_M���jT���&�~4>tꃫ�< ��g�����6Z�wjzZw������쪹����l���T�B�p�؎�F�y�9�W7P����=��:Uu$T�`�p:�֗S$8>�z��C�v��i��o�YgK�5�ϛ�K�#`���&̆�}���[�{�P�v���ѵz��q �a��a(C�.I�E�l셜|\σ통�2�^�X��v����D�������=|�k���H�]ܻ����פ&�֪���h�λ��x�)Pހ�|Y����G4��W��N)n�P4�C��>����S�-��<�}?�V.�����@C���wdޚT䮠�Vl:�MQ�+EUE΋�q�حx��6z�tw�o� ����[>�;a�R�b#��u��#OwWݒ�n��1�v̎��C>�g��W_�� ��ԧg�bC
��x�[���m�� ��L�_Q��6�e�Cl���P��2�Nش�J�hnq��}���`�wW�˻���SS�-p����Ѥ��vZ�2�H�N�%���+���ɨtf�Q2�9��2Wb�ֶ���SH��}Z�W&���a}.Z6�6��yWZ �u���$o6�'����gK�]5�z�ɾ���bFWh���g�}��63@QydF��R"4�@���u�;�wD3N�s�eR0B��}��=ު5uxsN��J��	w�e�2��$d�h96o�FU��Oq���X)�]�W�p�ɋ��mvDc<��ɝ[u�⎙�l���{��J�>�sO3��Wa�7�Yh�J���h]�ti���y�۲;i�X�`�$�Q0v��ٓ�O�dPPEϡ!��ݗ�ֺ�6KU�Em��J��I%�9�T-N庑����'��W��9n� Q�|CѺ��Ⱥ��
�:<��t� �#cl5S���'%�U�n�c��#ǃ�����R���e*�q����@����7�fvOb�WKp��K��n�9�S�;�+�T���ds碛��ڇ}�+um�h7[�KItb��.�n�]����aq�]�'�/��]b5��b��ٛ�f���S��.�f��KW"h�[+i�D��\+6��:��;RuCZ�ht�u��G�!KX���Uxޛ������_G.���ڣa�p�0�����b����`r<���F�T ћ=t�LEF6�r߸F��ބ�b�U�*�g�Ls<� ";�!�]1��k[[x��ufv��b����<t�{�u%=�[Cg�}�9�0�LF��U��Ecr���b���n���aH�e�z���6Ga�F�>�L�c)㢝>�i��DPµB1�ax��\�<d�� ���=�4�+k����F�z^��eC��B2��n�^Y�I	$2��r6�fT�}��ݭ��)�P^_-2	Т@zJ�N��ww{�f�K('-�G�tE�;$9�؜ɰGw&�yjGE<{a��t���Q1�^b�éP��g쾍;�ĜG��PSJ̄��o-H��;A
z���}v�z�m��ńu�rɈ�,�iIZP�B�v����������~"d��2�~g���z�R.��T�؈��n���,�J��Evv}H_�6��̥����Y1��Ǽ��[���u�s�N+{	������V�L~�t��R��̋Gs����uh�NM�e:x�e,���Pj����)�/�_h:)ȩ���\W�IiXD/[�y:���kgEWB���es�]�H���9�S��):�+ϗq�m���ފ̽��ņ�Xk������&��FV�RVxF�O5����۶N��1�cOoe%��L�/��	�%m	�
l��8��R�$����Y�Y�k���p�LV��;"�v{��2m�0�A�,���:��լxy"^thW��8�h9]�Gvk�:��eqw�O�4�㭐��<�l�D[��m��Q�Tq��oovi�u-�K*����Y� ���I������e�Em�i�V�;:��R�!���R��W��Q�)mMD+�9I���p��u�R��f3����=�,3U�ے/z����S�	��H�>5��GL�_�+;:S��gM*C�>�A1�}�9!d���ȾG��I�F�kfa���GWT]��r��)h�#�3�]�;�0��n%Y�6�|�q?��p`x3~�ذ��^q{���#G�.�^��[�� ���{�=�OGn��8j�(���Pa�u����WJ�7``ս�/�S���	�/$���;6V�[���Q8�L�}��S�}T)e3�ݡ���ifüҺ���;1��w�wD'�N�xq���_��$�04�@���S��d3�B���I�纼�[r�5����y�舟gr�	bȴU�ח7��x��l�C�e|�+^��~�f*�H�Rkױ�ܐ�ևH��^s���e2���n�S����7UZo=d��F���MxĲpo���"�t����)4\N����%�]^���f��A�ߡp��U���@��(���Wo5�b7�{�k;n��ِr�U:�V� �	ȩ���Gb6���������a�Gota��%Q����t�F�h�� ��[��3���|�٫,�*�p)Z�*RV9��g���l�f>����>U�n�^F��~��w��фl����/�%�r 'ص���+����md��P��v�t`��C:�S=�S�|�k���H�]ܻ���\i9\TG����?={�;��F�׫ݰp��I��O�tn���ې���c{��ҧ_aVX�\$xQ(�P���Bre=�5n�oX�'*��*;O�t�"�u�����*�ĝ�٦e\�P9�3���e㥺�:^��]_�:3=S��#�)���Ly��;�G,MN)M-�錛��*3볳H78Mv�K�Y�q��3c��8(�v`�'֙)��1)���ȵ5j���hч��{uI���6z�t������l�����*�!v�Ft��x������ ��a��C>��[���GY���ݤ�=�0�p�XV����tY��=�a;ͦA<��=,o���M�=���W���W����ݔx\X�5��i��#I�BDG��@喤�&gE�k�p_k{����2���)[ݓQ5u^�:� x�*"k������o�����ސD�ٯndg�P*�OP6z�L\�K\Pi{9c�|��rDvo@���I�c�/H�΂� ÿ���l����dA�Ȏ���5�nW��>�dׄUG�+�:�����!=
=W������~+���Vϰ�\S\�\���:K���{����Ot����Mo7@\��b޳���p� R٧��njȺRd4f�m<�
u�zĦdw�MҲ���i�y/�T�U�`��Z��p��\Э@r�R�M�A��Gi�%7����2�NU��l~���bRI&[�C�ܷRfL�-.Ųf�KȪ�u1+Ei�}!>�8/����Љ�ΑC���[gg��uFp���b�7e�s�e8�a9	N0 �ΏO�H��z��q<z��CT�7��	X�6�d�|��7g��̓���~�9�OW�� ��rQ��6'Cl�ܡ�i��i��ǎ�
8�l�{k��~\j:yP�EP��fΊ�h�Tϻv\�w{b���B�q�
�e]�K
O����
�l��0�X)�j��OUd(�p����έY^��J®����St{}��g�/�ίk:�~���4���f�^M�]��; ��;xF�|�^ۇ3C�^TTؕvٶ(��}"�o�B5�O�����n�&H�H8K��:����B�<\��Y5h�w�of����YgTlF^#~�n�yf$i$8���^�k�kD�Ỏ���c�ux��N��{y?.���q��mҼ��7Ż*�zK;PXE�0����W�e�nw���Zy�x�_'V�uԎ�o;�\Ӎ���R��o(���!bX�כֿ��GG�ڞ��g,��^�Cw/�R˓�������^���TR5g"�k3��r༏4��7����IH��쳛�����'�����^�{{ E�f��#O&���/��(wB	C�ɨ�wb�ŷ�Fu����:��#�.GK�AO�Y����z���:�&��r��mջ�/���#�vd��QHϨߌ�����n�g�~�ŕ=ٷ�~�#�ht 0��NW����v.�A`��)!K������I��{�#����0&�e�,�M�vJ�+_��2��^[o���1�-�U�������}-t�@���O�EmN��B6��1۩�n��;T4l���)\U�o��.�ѐ��8A{��������D4S���D�|T����9|�eOI�{x���^Ѫ�_}�鉣�^6P.�e��U]r%=A�������\�G�.7t���?��~��'9^�T%�"r��s��t�س����<Ũ�zQ�:}e�v�ӳ�v�i|Io23iP̲9W>W�Ԩ@X�6eco�<�+v����&v���ux��dd���H;U�g.����(0�W�ED�Cפ��~>�+��+�������0��y�i�>��p��Ɯ��/�F����D�T���S����/�A��#�<�^o`N�P�Fc[r��k����7@�����I���o��C�Dƽ�A��&}�Fl��'¯\{�xA�g'wu<�d`CNڊ^<ےLq�G:�8�����<+4#�ۉk���뙮���ܱ:���5�֢|Q"G1�Z=�(��?NC?�w�B��.�%�c �ל�羙�ѫ6�e�8v����<�ψ\�E�)��,ܳ�k�f0�yZ�O[�U�!���%J�{>\���8�GBGso�,d+Ya~Ne�TN��B{t[��(�滄f�'ɍ���Ap�U'�8�k�v�i����}��ޭK;2@����5"�u��av�u�(�O53�pr�6ufD�m�i��Ȣ�zd�܍V�E[?��UzB�p� w����yx�����g�����{��3��ͳt�A�g��h�l�4U���V
�rvS����(��`gk�Y�[M9B�����5bȔc5L5>�!]1'��T+�t|eھ��u���*�Ky���]u�pE{�b(aW)a�+���'X0��S����[EvBH�T�Y�tM1��W1ثQ��{���q�6k.�|Et�cu���_�tޙQ��k�$���l�����-B6�3Nef�efT�Y��c��+r��W60���[�K�ׯ��ݗ�k=j�.�^Tޖ�e�YF��]j��
n��JumŴeo�����ֳ�Nm=[Jv�֊#^�#�V9��/RV�dI���" �h����lp�|����o;����0��;�)�:�>�7$�0���50p饬������]0�.����.wyCsN�(♥YM��'.���:2*� ���&�5�z�ΌAj�A ݄��3^6�>ҨQ���-�eN��Y��ucwpl�!]ڌc�J��5;���ݺS�v�SY]��T�Y���T\DwLo���Xo:�{v�DA�雛�0�J�r+[t6�غ��B��w��rKp}2�t�7�i2si�LG/X�T��E[Ǧ�Ɗ�F�����sr�ɏMW����e�J�ޓ�9g}H����o9P��>��*�9�u��J�؋r�5�q�0��Q�`P��V��W<b�M�ޓ+�{��j[���$T��u�n&������eZ���}�Y0f�°cH�e�\�*F��gj�q�N���4�7N|ŗ��7���c�wZ��6��EfQ�^�B�S�s H+��V�<7ޮ����D)�BJ���ƻsB���T�u4>Y�m5k��6�:���S�v�$����H4k3(H�Q��9��\��F��'tW(�|ޤ�"���5U��t6pb9�� �˅>��2+%v'���b�hyS�ȁ�׳Fm.�e�m1rJ[fp�����:�v볞<G.>9{"�6�˅>�Vj�l�֒�YG�y+F�Ec���U��΅�Q�V�Z�3X����)��k�&�妱�f�M\8��4aI�`�etņ6K���͛f��SG��C�y3�,��k�dј���]�q�đV�b�+���͇ue�MC�z�6T��R�Y}�@���S��L��N��7�HҲ)U������R6�B�v�,q�k�˫��/m �<Mtæ��Ex�_�%o6����ӼMu��weiT� ��1�G��Ch_+�3���Z��S�׷}`Vs��7W�Q5�D���<�ż����).d+���Lr��������K�[�Z��$+mqs�}�oHm�
w�?��Z`jUݛL�������Nڽ��Eַ��QԸ��`�m�12�kU�dY+����ɒ�D$۸�:���F�����fi�o�G��0VפoK�˴���W��-6���@����"f�N����׵r��z2���L=�Ӎ0gwSj��	}v�!cEΆ/��XdɃI%���H�0(F$$��b�dbM!F(f.n�i!1�$�e	x��$gwL�@ � 0h"F�0��2"��B7]˝03 �u�̑��71H̆�)2�v��J.�@�L��(�	4у��r�IH�32��boƘ��rP"c2��d �4#(�u��&y�
I1�
H�K
$����&	��&fo;�̤4Ȕ��I/;�RdL��b##(�)��;Ɖ�v�#DB���"�(U~�f��L}�1O���%����v�������"��Rh��M~�����v�yp/Os���g5b+
$�n����m�S��Z~�����Q��UA�㮝H� ��Houz���;B�5��w��w`X�'=	-�\F���T���%x��Jb&�;�'��o����Ч3�H��>�O�(�9R�i��l��+��#3<>�@�u���j8nƻQ`\P%�j��=^��������>���{���� n��¡;A��;�6�Cy��<_cWG,MN�+ =w�K�8_y�����=�Ki��#6ޏ8(Ȏ�zw֬O�j���!���n{�׷�vP3�>;cgè7Gy��0!t?b4*�bIi:���w3�n;�^;{g�I��ʮM�>&:N��lt3�̟��=���1H����!���G��v�Q�J��� Y��i���d�h:+<k�l[鷔�5M�Ǚ�^��
4.����h߽�sӏdD�<%"4�g߾�4/�@OLom P����4{��r�S���!�<=�VϜ�:��w����ɻn�y�w{k�F��jʔ�1�e����8���)��x���K��RھC*�jqZ[H��ug�:�^FL�:��\��pӔ)op�p�ɩ�Y�.��<K��=%I�e�/�.�\[��X�(�{�hD��^�-H �K�V��{fl��:�+h�n`<H�YGi\��g�qA(z�ꉳ�옹:��;G聤Q�3�q}����O��I��d���Z
��w�WK��%mt�%��i��T{`��qJtW$dQ2hA���]�&����ݲ���\���i�z�Ř6#՚6�s_���/	$�9�}w��Q�~8�U-<�����7�J��\��S|�+�s�ts�P�:Wnv�b")�6��Ή#��S��A�K�Ѥu��h�.(��W7�6#XW3�e�탘���"�r���za�_���r6f;{���q��V���<(��F��{��< ��ڃ��{��s� ?-����#*��k��#/Oh��l��#�.�yP��b�n���a�q������Ϩ[F�L`u`۽����cr+�i����$�7S�%�&�`���p�3;G$[��+�vL��SS;��"5y���T:��{/4�e㹬��#)��b��N�*�%f���o�DK�����(É9ݘ����S���7fh����͌���},�a�p���ƱT�\�Z��Ǻ��U��E�n��Dn,a25�f�>V?B�	���p��ۚ��"@O�t5FH��6l�]iRlsđշ\;A��8r<��#)�l�m�4	�	�̿M���T�NVk�wU���+�d��~�j�f�W�ʢ��0�nR򜲬gc����;��kO��n,Ė���y~��tBZ��W\�\^��SW|�����;�DH��oDg��i���x��=�A-d��7Xəv�.V�����w&&6@�����Y��W �]myKU��t�nb���46Fg7f;���G�2��`�-²8�gJJ�)T!u�;wT�E�{��!��ٺ��V��=�c5�!e����s!!��'�t�:;ĥV���[ywM�B��~{�{$�۹'��i����0�H�V��	��#��󚗇dy�Es5�j��`8���:��!R�em��iS�����3���7�7Se]�͞��n��|������g���m�7%���9�q;+-�L�cJ����ܷ�I���D������T���6�Ft���LaV+h��	�aI��h�y:8��{�6�����fh=�b�o8"�Ί���vi�B����n�wNj���(�g����T��,��Z�s;R�[Z_1˾�6�Or�@#w��ĚϪV�oL�E�P2��
1+���:<8���G?~�j�_��]q�Q����W_�g<����I��M̱�k/�aa�f"�g�W�n��j��R�Q��-����Jn�j-��$f�h���cS�:�Y)>��p�#�Fᆋ������xѯ3�p�⋤�;ʩ Lt��#�6Ƿ�ƎgA�dd���}�[�13-{�Z4N���-�x���Lt�����gC� ��:�T�DLZr�p��ο���K��lZ��I#G1�[�I��O�1��0����B̠"6����g8-�Q�������K�q��Z*�Hا9��l��牡8�o@dG�
��@��/���Ov�s)��T�DΫ��q��H�H�VY�`��]y	�{kv	�:%*��w6���Z���x;w3��v�s�ͤ�����u�CI��X����u���Ĥ�z�?-
����۞��D���z�YB�	�/Gu�d�HO����48���9���L5sL3�u�3r�j��6ǺY�v95T
�,����k��]�UK`�Ԍ�=��g/zt�q�U�ْ.i��P`��#��0xG�l&{e������v_��b{�i����	gz�R��<r�@�n���@)���:+yql��s��y�؅Q��l�$�<J��H���p]:���[SǢ����ֹ���T�ȹ�t�=	-�\i�L�:��6d�s�v��
�k�l���
�1�:}}�<�J�R�i�քͼ��6�z��#���N��%Di��؀r7�6WP������)L(>�B.��iau{�}�����mp��`y�����8,X�����Ę���Z���q�Dp���C���x����=f�#zf;���r���
�����fݓ��ԧ�6��3It�^�nܜ��W%}��C�r�W�8�!"V������ܙ���0aTĬ*�UI�ދ�u	�FZ��O�>�S�!��9��곒���H� �3k6�V+IHj�Ôe�Vh嫛)M%.�.��4X��\S�I6O긿���������t�퍑����|B�"!�����0q���!l��m�x��7d�c�����CQ�V��K<TS��tp;�{�.(��Y��4�	�����y��3nE;�MT";�=����h3�@"�?}�F�L^Y#I�)KY�O�[��3����#��w�75Ъ4�`=�4"j��ԁ��Si�]����|S����x;�M�x��j���z���M�d�Θ��h����CN�v��p�"��A.Ɛz�\�k�N�e`�\̷7dK�-�c�W���_ט�d���B�H�d�UG�$t���L&��Yܑۅ��N�Ka|�:��ml�r�,�pI)��>Z았��;X�y��l��ǬaE�If�C�.cH�*��"/�H�%�lvz��6b�4�QNy�	K�C�zT>�O]jm5���Ve�3om���v]ƪ,X�%��C3l�*��aa�]�R�d�� 	ӧ`��;�%8��բU��C3�ǻS������QŔb�,#E|:''J�2�M_ܩ�\�+���X��"-f��^:�>���n��.���(6Q��N�nhC �+�H���)�Q�����y���βk���Θ��Z�m�vzXc���VX~�G#"�O�O�"��>����Ľ�x�R�ZV&V�2�7!���,�>������:Ņ��o��4�:�l���ʭw�[��Ϻ�?�8#y�T��h��5
������7��H��4�ҹի(=Ԕ���6z���3)E���P��k_ �[3���>�f׮\���"B~���bߤ��-��q��}y�=��o�}Ԯ�Xl�<��}B1��l�6ϑV��fj�YޘE+Z�d�졼2ɸ���U\��,�xThFg���ng��`^Eme]�����ف*or- ^_�[s��,�I[��YL2.n�a檪���K˶�م���y4����S��g�ݞo=źf�;s��mOa;����{z�	:��q�h��
%~�O���X%�j����%"�=�+�;�P�7�M��\�p|�Y}R���L��Pt�;C;ϻnX�4���N�T)j�R�(>-	���{j
��3����ɛ�,1�@�U�}W��SA���H�"q�뒔q{���d\�җ_���R�)u���R�90]������ު�]ylhc��:�$Ĩd��x���-)T.��s�;H^����s�^��D�B��6���	��$v.�s��P�6�D��9�E���vN��ugf.s�S�܍�Q4�:�ߑ�Q"�����m3!)�њ;:�qs����	�%�l�R7�%�ʶ�x(���)���A��I�;��*��q�od�~�H��f���W&M���!K���4�=����wM�����������*hYMV�飪�'QnЌ�m��ތ��ʦ`�/^���1�R�1�Ccϑ��k��rʡ��Y� �&�UR�v�y��F�ѓu0")��	���ޑ:��қ�Ni�%�U�������f �^I�r/�v�dT�';�#��[Q�G7l��I������ތ��x��B38{{J�����W�"�do�C��h�;����V)�<�e�F�A;^_cu�'���fց�s�!�}����[���p���o�˹G��cl�+r��q	�����Mܻ�K��Qx�W\�;��%mJ�2��fu��z�>��FwoD��NPJ8�����q���#�g$,��>����p�|�Rm<~n]y�'�5�-� ����̎����� L	s_Zh1�dSDT��&z��"��;٭�}j4�7�Ō�<�3�#!�Iiv���cг��쇓4pC���KK�d�Ϋ�#;��%�H�Z�Pz�fL&�L�jz�#+!R��^�TMD��z�2B�����m#�ky����Fo��w�X�Y�.��e�+��{�4�J�Ln�6X>pDoP������7�M����TfH4�}A�U#�D�Pev�#.�.�V����]�}��U�)Juч.�S��gt�T!���*B���;�;����wQKG��$���y&�*��EU��W�&�_ᛦDXc�eh���!�Mh@)�/�%|��3�WQ6P<�E7�Pw噵�WY��bΝ��T�p��-,_�l`;�@�Z�=!Q%]�`�d�����R�ɮ:5��XM귝K��4����=��xM��=����Wv�j]>�]����x����V�u��j]�۬�-�,󚰴��h�r�PZ�ӑ�1�:o��Zx�IG)\�a��[<�&/7��c�$�u4]�^E� an[ޘ#���O� ��kcwYځ}m���nH�4�\0k8d�+��]� ���B}�,C�3���@G$vwV�f�Ԟ|��{٧�wz�2/%��A�F�8(�Z��g1�5�6$ֿo_v��J��-Y˺x��������}Ϊ�L.�3q[�����3Wr2;o��]�����zLt��g�A�#)���N��7�8wY�'��1�,�?�����8&Q����t�)ɋ���U��L���꽎3� 7X� U6k����������4���"t�������L�a�{��Y络�������F��ba�Ѡ"j��� A��ۚmQl��okOl��D���M��ܙ�ng�C���j���1���=�W�(�EUTV�b����}��|�(����xP�L0�i{j��k2�f�f�3m�[2�el�lͬ��2�f�3[2�f�f�f�f�f�,�fkfm�+f[f[fV��̪���5�6�5�+fV̭�U2�3[2�Y�̭�[3[2�f�2�2�2�f�Y[3[2�f�3[2�eT�ٕ�6�f�e�eT�ٛY�S5�6ٛY�R�[�-�Vf��Y��*�j�ՙ�3[3VYVe��Y��-fj̫3[2�eY�ՙk3Vf��Y�f[fj�ڷ㷞|٭��j�f�����vmUL֪��U3V�f�TͶ�f�ݖַo�~;u��e��f��Ͷ�f֪fڪf�T�j��UL�U|v�o>m���m�*��m��ڪ���fV������m�6�l�+���[m�6�l�m�f�TͶVUVUVUVUVV�m�ٕUL�m�5UL�m�5�ٛm�f�Y�ٛlܮ�������fV��̪�����j���y��[2�el�ٕٚ�-S+fV��ճ5�+fV̭�U2�fFU� �1��������UA�EXa��!M��]����c���ö?���6��#��t�~>��_��t�,q��"���'�y��G�QA��*��� |}���<���O�~���C܊���/����z�N��y?�~�M���~��u��G��յV�km����m��T�m�6�l���5UK6�l���e��m�J�SYZ�ke��-eUSj��l�ڪ��m�j[m�Ͷ�&�T��l���Z�d�QQP�"�����>b�+lmkh�Qj�����Uw������!���<�p����<�jv��r�
�Ȟx[��:���8>���{�w
���D=)��Wt� y�����:?xw�"��;p� *��ObP>v_3`��4�������ݰT` V;�����UEzR xc�۰z�Ӡ����pdh����~��UU���P�E�'U؞�S�@�{hI���HP��K�AUTV鈀��N�DHP����p�2�;���u�PEz�
�,����>�����Ñ�C���e5�}=v 3&e� ?�s2}p#�=�Q)*�$����JD��UHD@�H@��IB �P�RU* R��RI$R�AT%*���J���	U=�*�lj��*�R*P�U
	_ZS��J�HUH$J�*� P��"*��R��e!*
D���R^�B��J(B�$�����T@UH��*�I(D�	(��U(�%
RP@IB�BPD�Q�R���URQR<    �+�{���kή�큵1��l{ܫڶ-o[z=��m���7]Rƻ��]�zV{�����mȻ��v�lճn��mk3�ۺ�wW]U�o������m�:l*Q��4H��   Z��{bCFMhhP�.�.�����U%��<���44(�dg<�CCCC[;ӭ#�}�n�u�vۮ�fͪ�۽Uޯw��G�]�wL˷m��]�FuVUۻ�ڧ��1	(�J�U*$�JR�  F��A��޼��{��[s�c��<m˧N����-z�#G]���
ۍU[m��:��z{��W��8�\{{��O^�wvݝ6t�qJ�kv�%.C�V���{���t�J	QIBP�٪�| ������v��^�]�]m5�{�����m�ަ�]�u�wS��mݳ`���k��3����f�Z�G\�g]@��';�(���n�UP��%%T*D���A��^�J��r�kkg7ln!�ov�z���V�.9λwb�u=oTZ�'Z�V����N����q�[P��x��ۭ.��J�٦�IB�(B-��	�ƭ�d���U�]6�9ֆ�T�'\t{�釧�v�TwVCU�m��M���݄N͎Jn��N��j�z�mJ�/f)IaUNڋ�ۯsj��L�K��OF�����PM�v��'nѷf�w!���3#[����*5��g)Wp���T+t�D�
)R�Q[j�|  ��%T*��Ф튆:X	:;��TZ��y{
A�K@�"��u
J�+t.�UH�gST�t�s�D�vh�Т�@P�R�
)%_   	�����wb�BJMʭ�ET@�-�J�J���l��U9��$�P�]�â��)qu�d*��Î�Md]۟x��ccSr֪
J�%
DJB%>    ��7�I�p64
���$�UA��qT�J���OzR���7%(
�ݦ܈�(U��J@��T�TU:WtP��> �~@e)T� ��F�Oh�JR�`  "mUT�U� �S�A)J�  ��6��   	=T���R@ ��O���_CD{�k���vr;7!�NR����2`Hή������=��p�?�Vڵ����m����[j���ڶխ����V�����[_?|��9�^BT0�G�� 5]4�-i��j;YWׯ��c474��	
L%L�����QVD,�;F�7dvް�ݫ̼�t��E�mB�論�2K�J�R�%��J1Pc���v%H�ޛuhf��ٔ-*�1���bu�ֱ���t *,�t^���]�X��54���fG(in�W`�S��8T�v
[R��Z62%Ʈn�h0K�؆�6�{�U)�6f�B�Ԩ	��R
�z�T��5�tZKj-���r��B�Sl;�	�Klb��!Z��OH�FU���u�WESY6�,���e���B��4]%�M<�A�r��ؤpF���&%�5U�5�t�,JN�wh��[P?�R�cw�yR]=_Ce̬N��QPYH\���skfe����%��[O-+Gs�tR��r��jȖ�HS_H]hJ�W�r��.��Y��2�٥�coe������F
;Y�I[�h�D@8u*��0yhk�+���m���.S�������Odt���C�qbܕ����4��lEZ �q�.�f��t�X̤����Lİ볶�5x{�����[��<2̉�`�u��r��i��J��I�h����H���R��yLLӵ5��3��m^.��ٻS�)ˀ��%"�����ҋwl��e٣W�\�	"�Wm %�&e1a�ub^��F�%D��e�TQ;�j�x��B��ܧ�f�k6����('MŚ�J�I�l;��,�Ƞ�Z���Yi]^����[�^nj�,7VXEv�H�\í'W7*�bl�N�~���Ve�� $ɀ�,��>J�6;�ڛpXa��XfR݁q�LSTy�t��Tv��o,�ڕiTUt�e[ ˥sFS��S��E���J���x��M�؉VE�f�z�nŲ�!M��97-��N�V��ӥ�a�h�^]DM9������ GH�����3^n�ݕtąkf�; ����̫��ZX�vK9{J�q���j��ʕ�5�\K��Ф�B^����`��q�j3�4Z���v7s�Uk-jhD�K{r���5�r6��-��e��e�l /6B�YH��T׮E@`� �Hč��p�o�$�@pe���"9md���6nI(�%KQ�e���?7/\����n��YB�Ѡ�(�-U�b%yF���>�W����am���E�&U����ZS(��mL�m��
�f&�c�+*i����{4�X�N�6j0sUif��7@eז�n�F=�ĨA�Ɗ�z�n�#f�ňaf^\����c��'Ld%.X�Y'�]^ZI����ZәiK������c�����h&����Pe]9[�"��)X�y�N�C]��մ/\�;F�13w--đ&i��B�ȨډS�@8�#t�ݠqݩ�nX��<T��sR�y�As� :���J�@��Oh�ڔ�Y��Y�[rV��v)�uҎ��_,ʄ���7v�$1<N���,�c
1j;4H���4Y�n�b:�lv�Z�2�2R�4le�A�O� �y�{w�0:wj�+r���tLtͦ�7m�	ϝ$P�r�(��-�'-��JC,q�n�mHKQۂ<;O^k2���R%@�t0ı�Ys5�q��F��XU�{
����-aV�n��

ǆ(�p^�Xs)���h6�ٵ�aX��]%iyg	$=2�ì(�kN��b�fc����Gf����V�arFΕVO�LRՋ�h|G	F��uYՐj	:��oN"�_�@��K1J4v��H��T���bZ�Jf��VӼD�)�;�f��/��r��'H������E�������'t����f����q�4tO�6��Ze�Q=��i&�n66�b�òY�e�\�j0]���z�ջ���pca��j�R�L�j�����ӻKHQ�
���[�7B]�4���wd���RsQb7A*�$�i�EC/" ���q�Uu 4<M�.`�Jӷ-�JU�oFV%{�t�!�c�	�u4^��u�1Y��ס�а������ �^b15����YĦ��r�z�Q��2��l#z�U�қ[�J%fL�.e�۪�w�Ym��28�-�e��\0К6���y�+v �K����)�������R�XƤ�A5n�0�I�\/�3\�z�tŌ�W�7 Wt�㡘�f��^cxjS��.��QB@�Fk�^�Mr�J:�v�0K��cʻ��S�~�d�	Ȱ0��N���ݹ��)���KB�j. ��Yl� 3�V��ڒ��@ ^`�r��a��x٩5����I(�jʋ+{x��Ë+�j,U�H��@������#t�R��] �|v�[l�&kV���X�LM�E�lF��y��@��X���q���-���z]�GEG�2�m�>J�;��Z5fҚMc�&c5��6Ģa{В�]�K@�5�xSn1h��H�)������e���$F��I�HT�j��]%Yܰ���溸	��.�ۥ"[�^�ʀYy*��m�3�i���EbUفTgS���e��i@��짘T�6�[E�kFk�X�^�CC�vN����Ëc&�ͨ!��1r��{b�B
iG@nӏ1�/(/��m*;���0��nl���
�6��D#���M?�Q۠h��2�
���J]n2%+ ��:7�Xկm�R�R!d�/k�j76�Ϥ�d[ѨKǊ{M�ZIɳp�e�6���{���8�$�Ö�r�I��6�C.����;�.`o4&��o]��+V��)����%A$�)���9����$�wh5Zq����&���N��KV�4ش���hKt��w.�OV|�)�1);��b�M��0pn�ŧ��R�(c�۵WD@rZ�Wv]�#\�)n�W�H#�(Zd�7nl LZ^;�fl�vL፾C���^ڦJ�*jǲ��`(�ڈ�IL�ѱ�E[I�����Ҹ�6�����e�*�ȗ&�af���SQaJ�љ�#�ikcsp�QVӱA�̬B���aVe�d�ʼ�]Ar-��Uѽ_%�V���t!�y�A= R��������*­� �$��:�季Z�� -�nCAH.<F̛ 9%�Y�^L���S�1���&����gj��N�S,�%:d��cM�X�P�����SE��^����Y�� ���lhݩA�]�-��J�CʇcEc�֚ͺg\�kVD*@-��l���l�܊��P͂4:{�*)�8��LĤX$f�YJ���u �-l��z�t[���cF'7f@�d�"���`d�,H#m2��Y�
�j�ޜ�yHd�@d���%�&miцH6�&����
$�b�nh�����/vT�x��-�R3���Cu��\�,8�;RG�JΖKŖ�[eZ�強W���q�����a̧Sn��
�-*�-Zݎ��u�P�F�"[yB��ۼi�V�i"�������MR��ddcZ�/S%�W��Sg�EJ��n��Ǆ�368���g]�6*ɧ�$O�X���6����� j�	�3\"dg5�Z$� � �jܻ���2чTʽ���=�v֓^���I�T�YR�n�m\��[$��N�k����VL��.��eڙ3FL��4�R�Pa<��f���mXo$ #t��`��,�Y��k�!?��f�z�ǘ�4�=��E�)0��K5ں(��a�K&�����[�Ќ��&����V����e�٤��4l^�L��g�ؖ�s*#�ͭ� :2������d���(��Ѳ*�[�f�Y�{�a��iK��(�44�Kݍl�ȵ�u(��o.�K��D��li�[6e+X�)fô���Jô+f�ۋa5�u�K�z.*�#'f`�t%ktfn}�45�n��t(��%��M�*L��wh�P�OV��fPZ�V7@%��@vƻ�O"[2����J%u ��#LFƻ�0 9�b�C��@��[��h"�ͺ�g�R��!F ��,�lk��2�T��Z�k
VP� �n"�������,x#���5- 1�Wn�\Oۂ���SL��K)�
Ôa����ߘ�0�/pe�݀,�� �lJ�R��)˵��Xx�ʏp�(ʒ�ץ�L6^5�^={,?�<�ItڡeT����M�J�kz@�DEX,)v��U��(C�e/�E+�R��6���Z��	�;3E���l��u���M*9�r�L�n�*��:��	ffT�6��fL����Ew2�u�Վ�i���"2��Iύ2���]F7EIV:��pbG1]�Ѵ5a���J�7#ۚMnm+d�҄��,\�n �aR��lf�7)PWtZ�4�r�jDT�/o�5��5co3 bN=q�cs6�m�14`H��ON�P-ޛ�Jd�[�5���1�WFމ�4�5ha
�V�[4e��]��W�-I�b��މ��ӬI�5�b%٣�h�U��~nwAb��[ _�ޣ��v��H���nK�EA���r��I�ni���B
��5fL-��t�8����	9��y���C^���٘�0;�*�O�&�tڈһ��S'1k�WR�8Q�FÐ���A��i2|�5� ���⹉���b�[ܬ�f"`N�M��9��z B��d��y�8s#���r]�n�J�]�1V�m�Ÿ�	�N9]�v،0^mr2p,m�ZCW,Y3v�[�
�E�b�OI^�W�l�i�A+P���4޼��A��6K%��5��-�h�e���D�	�*�%�G��Ԟ��J͆l62DDTu+71'1�ܰ�z�������b�g%�;�M�(V�ʢj���DHRi蛎�PY�q��DJY�����U��3tEsh�R�;4�c0��&�f3���+Ӕ��2)*�ϵn�4"���T�E���^�5N�ݔPʃo/iBU��Қ���OP+[Y��í�_­3�� ��-��A�-Z�ݦ��[�$��0�/*��bP�9(]���
b�;�
���Pc��LA&]աJ��mn����r���R��[�A�i|��1�ӵ�o+-���L��6�e+�� ݭ0+CC�m	��y�1�~P"�\��[Ȍ�)����ڐ�ԅ��2��m)"��R�TÒC�zS�j�Q4F�h`%�W���=%nE�$�j�V�ò��4�L�a� Ǳ*�K�̕sqV"�ӧD١�e��̙Sd����ݭ�Z\S�JvNHZë��Eh*��K��KI��a\8m&��'���6��I���QU�����3mA�
���ùZ�+����
�X-	u�.�ԩ��6M�����vf(,feL��i�˂Ea���(ag"��e�M]f� wZ0X�L=��kPq/�t�7J�q�5
ѕ2�b�»_$�EZ�ft�2ka��W	����^<��5�Q�R �Vsif�O�7���w�mV0����R
5���*��sY�Gc����q�馭�i�2*YgЍ"����K�
�����IHې+ɕ��BeK��l!tM���x0B����#Y�6�f�8�h��H+,�u���r۽#(~X]�K,
�m�QkM�,�53%�Ѧ*��`b��0��5�x�˻b#*�wY;W�v_$�������
h�u��J"�����*�V�u݂:5��&z��B��r@���*�1)%�R!y������l�UV���u�t�6��7�"�Z���E��)cYY��m��ahw-d�Fl���c��~�F��[�wc�qb1�5!Q빎�e��6�XQ]=����u(˧��D�z�:�@�`�����4�і�yt$��SU�[�M<�X���j�����)�`����S�W�cyqj�Gn���aϑ4�V�.��@�-��m�@^�*|��A�V��ͽ���2��(S��`C�eG���X�k1��m$�a�3@/5���Ǵ�"LԓE'M�n�_�]�ق���U$S����q&+PN��q"ico(�x,�!�b��d�E,U������VSwOв�o7V�iF�;�Ǻ��\KL(m)6*��e�$V�F�Yn)��t�l�[�������9����hzkb��n�u/pb��-5�J�&@al�D�ݩE���y��t��@n�J�ӎ�$�*B1��2�},����ՀUØ�M�N�Ѻ�6	R�E�n��+2�Rˉ�C;,��'r"M�
T���5�+R�E�eJ!N? .�R�.�4��Q^Gx�ĭt;�[��(�P�Nk7d�]�
J:6K��Pݔ^K�Z,�.��Q�eL��kr\��r��,15�Twnl���5G6��llI��-��- o#F�]�t,�b�x��n��(�oY��כ�5j�h�t�^��KJ-9���a7+!˳�A9E^�/y��*`DF�f�r�Csە�̺Naɒ1D��i�pZ�U�Xr5.�E`�-���ҳ�]�T�T�m��4ݍ4��#.SyODp:��� �51,Z�a41����n�%D���4����1j33 wm��'E�`���� �[I򉑔�����F��9gq�*Ь�t�h⦠�iV�F6Ҭ��t�-V�#Z�y���3i�D���b�*�ot� Ǭ\ H(4�VZT�חE�MHқ�F�{$���@)-Cr�
&���/a���� �U�lx�XfhVT#�,<Ԩ��';�]�4@�ŉXy�!��/iP�� �e���������y�J9�-��6�r�LE�)w�H��
�c�с�4�ǫk�,��ȗV�����V����p��o_po��yi@,{:�Vֹ�^_^m"!�;;o}�,@tӒ�N!w O�h�q�ʝ�W`f�����ӎ���{E;���l' �k�
���=Uvd3��v�N��[eV�Ѝ�r�wd����h�w.�Dd���V��X0�W�Ʃ=w{���I���3�1��zk�׃���	����&�M͉��P���,6�7}vp��W���J��4m\ڋH�4��o�%{��@��Y�~`	�RQ�;>d�o@k�U�Z�V�&Cy�ܹ����GfX�Ϫ�k;d*��hB��*N�����zc����p���� 똈�)��T��n��*�0��t/�vb$v1��CICkl�+ju�l�u�3o���>��5���I�G�t���ֆ��޷V��R�� hjF�Ma#cO�ao��N��sx��[�vp4� �/��B8��dFJ�Z�a���p�����I|�ףmްoM�Ch�{L�T�^�;��_)��6�i���& 3w��GZ�Vf�F.u��,o?��Z����N���d\p�+3*�C�ԭ��2�8�N�kT6�1}"�lK����t
������jVLA��kNl�PkSX(�u���U�4,�X���Z�3(�xsw,���Y���<����I=�9����ܬ��y�n�h�;�ˠ�a�l\ۭK��)�z���+��+5i-�ȿ�Е�:��s�ř��ݺ�[e#���J�G�n��$Wi�' �w�b�)\QM�FecHt��f��x���9P:�3w,�K��ގ<S�"E��ر�P��3n�N�Aԡ�權�Ŝ�C.���9�Gw��9զ���K�AQ��*�,�'jX�9��).��9�Uu�y�b�ѷI>��5y���D؉=�y.��N��y�]�����G���v���Ds���8QR�ב���#fPm����K��r}w�� )�ʳ)��]Jqn�Ի���L�w�C/-�狹��8A���z�*���ν1�-��y��yt���m���}W�"���u�K]�� �u�K����%k6��U��s �A�1�\V����n�K�˼�L�B��e�텡Ƭ�֝(�=�:45F;oqi�n�VZ���VZ�2���ߖ>�V;)�d(����W5����wC�����ʷ����bh1;�W<�T�V�/�7��N��f�x��՚��������k�����ч�_�\�Jr�3b�@��oh��6��C�Ų�=��}H�qWK���ۓ�/�\�nm�!�SDf��l�����ƅm��q��u����qp��릹K�G����j�Q2�>�8�
|����k-�v�`�������/I;v���z��E��k�.3a�vo�M>Z%�\���f=����F�n���\r25��-�b��M�Ν���}.�][	���ѧ�Rd	���RW�nnO�,ثF�.��(ܷ�NK$5��Z:���$S���9��Bt/k]|9cicC7d;�<Q��r��O�z;İ�.��r�!��fk㻼�_F�[avV�u���;k!�՜�☉���n���n�<�i{Z���׎�e�̩'%�IV��}����𱝂�Ӡ]�#ڄ���c�%�ւa�M�L�tD�)ռ� ,��Pn��w�+���vEȦ����I���_w�z�Wj}�%�����v�43U�U�8J�CU-.Z��W�/����Y?l�eQl�u:WU��i�N�9����(�Z3_�ql���7��Τ� `���YW������ .2rњ���+�w��:�r����L+Gp��· t��	6�(*�y���a+���˾8���+���]�V�v�2�[��"��G�&����V�;����;��nG[��ǐ�٫���et:��s�L��!�[q�鬮Is�Hs�+&�n����Fu�WI#��c�o�yw��b
b�Y�YRf�ɂJ'ɳ��+��{�5w:����]��	��*j�Q��-�ڡ�Ɠgz�k+J!a�YNmv*��M2u�9�c��N�_O�}n7w��A+'Ka�"D2Ƃ�wP���Ox�|��`��i�%$���Z8�a;���>o�>t����;Q��'#|�v�Y۲�}"f���d\A
��K���V]��!X�3��V
#�6���l�hA�6��wN��Zc�;GcG	2���$kUuj�V��v��X�j�R�V�p�6ڎ�Su�V֋J'i],����R�n�WSWji�ɤ��WA��J�o��Z̀V+�����:��2�b�Յ�o��6�Br鉎ӓ$�����5�IAnՕ�{���E&��{�wUw
�@疧c�wE�<͌t7�iu�x����}ʻ��E҅�	nYwE����\M[�Z�-�����wn�r!�u&�經째k'LN���A��ږ��Y�zkf0��Z�%��vĦ��
�n����Wn�U���K8��d�ΗV
�ʮ�|*@��<��ظ����|}�uJ��;B6���G�em=�l�J�96+�(>�����=YL��t�1�3�����[�6F�.��m��fi�w#�j��I��v'��뼾
���������š�ŀ�V�=�YI8�ۣ�`!À��c��T�]g��k�������z���橒! K��[[�2ʣr�8>�z�趱��U�6r����FK�{�����R��Cw���U�1��-K��pVR��X�כ�7���t;���[�y3�^-�H��Ǚ�
������ޕݥ�`<5��0��iU�<x�a�;4R�����!ZG��-�Yd�ӎ�U�+%W��SXX�8��R�oK����N-���,ܮ��E;Q��ģimN�a�9xD��շW(AǛ3�&&�E�̼�u$Dt�+����Vrb��v�k8'C[�XP���}�@H���Á�M����:�]��Ft*��EuC\avЃ(�Z+f�/,�o��ie%�>���W�A�V �H�̹�t���TyI�;2��GQ���'|u��p)+;��3��	Ȫ�P�w������L�a�Dw���na�A��v[˺�<��D��VW���Y7�����{��8ʒ�>���9����Zy�ss*bl�Q�:q�X��%�2>&��S$<4v��&aoo[�G��<z,
�+�9���}W�V�&�'|��\-�ag2�c�|�V!z�4q�ݭ��r�*ס�5C4���6�k�i�]$s:	��.��95���_>�ǰ�vY���� z�M�[���K܎��N1���Yl��9��]ˉ��IGnc��t��6�G�(mY�X��&��[VO'E�u�W.�V��YoD VD�jK.�b!�Vn�1y�.cU.�`�]3T��He��8P���E�E]M��خ<>.ks���lYv)݆���u{-&09zz#��Q.��6+z&J��m�q�B��wd��t�/�!����m�Ȏ۸�mr;"�/��]]�X�}G���є%u9[����"1-��rp5��Vr��G8W��(t���Zݬ�F��z�rNՠȷ�^R��YԸ�x�}O#�s�d"[N��I��t�X:�OwRoU�����mm�`&D�x���,����0�9�hi� f[��f���Ҋ��%K�U���V���fTu�n�:d�"��{�N/y��K��Q�.�]�|�ج�fI�T�lk�*���^�AO�mN��y&Iri�b>xgl�B�V�|�����,�]����|��jʭ����(^����cPL�}�F���U��RY��ޢ޷�w�0��fn�'Ej{vW'O@��TW6M��q,buy>w�g�*�إK�Qt�Nå����ںv��������0n`���v�8��?I��}S�,�޺Ol��w���Έ;��,vv7������`�kR���6�u��)c2��&�]+��f��5b_X-Qѷ�b�X�;(�'��m2��UkE+�EZ.�]Ԣ2�Ȥì�n.���e\E�{W�#��V׮����Ӯia.^a�9�V�:a�֋�:p6��W�쬷�
"��+�p��@_Uy�,nM¨��cw��XEK�]5�X9s�w�M�Yx�ytz�v���S�7�RXU;'�NН�V��^�ɼx�!뿺݉�9�k)nr芘�3���'o�JzɓY��m�8�BQ6��}��.�[��urʾ�_\i��o�u	�s�0��v������o���7�2��-b�ZGGm]�$����lu��j�rީʹ�}�e_���u�&�_T�0�b���
v��*]��&d�P�Y���Lι�.Њ���S҅����l�Q=��k���l����r���tO��*��w�mD��q��7�ogb�����Q㻙�ׁ��+���M�ͧ��T�2��]�U��^p���c�}�l+�tɳ�q�v�i�t�jT�X5��ϺJ��I#��ɻb�����Z,o�/3�5��@��kO��G^�Qa���V/b����d�ϏOn�%:��{�d��kf�Ы%b"T�WP/\a� \���ç-�T���ŝ��N�YC��N��-?�jU��5���[G�EX�����Y��u]��
lm$�a���*��L�f,��v�ލ��}�n=�m�׆�7�ܩc>�q&�����t3��YyAu#�_+��Y
F{Z��L`�z��N˂�Y⦹p�� 9��j!�ru�wdZ�h��wѰk&b����G�XM�LkN�L��T��O�����U��ބ`b�HQ�|k����8gH>�G�C�x��Ģ�v{�S��Kmж�u	��;��=H�Y�5��K�C`�&s䎈�]C�(�	nΪˢa�iW��\�h��aƥ]8���}����q�q1����b�)��<a K�Y��Z,��1]���S2wY�[���uvd2��)�Γ���b=³��m�h��]W�����d�#z��S�W�y��-��ã@���3�n������(�XH��$'�V}��F-rڍ&�7��n��}�j?�+�I]!�dΘn�Z���9��:�Y�S3����ADQ��"�0� ԴU��9d^'-- �ٸ���qo7������[U�XR�+Oo ^�7]A;��0�ɨgp�*a4~D	������=�͔��76vuݥ"�l�4p(���I�Vᘬ��x2�E�#�S�u}uۘJ�&��'.뚼�Hڰ�p�v��Ō�=9,��ѵ�5gy��;�f��r���y�-g ���Z��u�q�ng ju��o_Mo���9�n���Uʲ�ӏ����H�h��γyR(n�x�.�yy����N�v�v�
���V>��h�ʼ8MNW�m'�]
�6��ߺ��ri7��X//�#���Z��}|U��� ���d;�oG.���s�w��Adlp���Ae�gf��"T88؋T�㺳����)����v{
��V�q��+g��{�v��l�B��L�o�(r:�j��N�{�t>c,R|C_Ǭl8v�'� �6Nv:��x�,��h�r14{�Ŋ)��받�|���z5qs|8<+na���g%f����]�\�f61��Ƒ��Mu�9ƃ����D�=����.qY[��qS6�*V(���.qg^΍�gU=yCd u=�/�,U�5�v�xd��C�������Lv鎾����$�5W]]��0rN\ʅ���e���	W�k1J��[V��\��5���Í �	՘�OF��T��zU��P���l�2�����h+�`�=6�� �v�<��>_MJ��@��qѠ\2�@��g:s�2�	o�W^^�*`j��T� �ⰰ�ՉyΊ�v8
'$:��z���chK�O-hf�A��7	�;xЎ�0��DN��ν��f��ڔ:��YFNJR�!��V��|N����\)Zё�d�]��$i�b3�Xlo�$�DC�@Q�V��zn��sE\���I��]�#�U�#;-�N���"�M3{�5��y2��|Ŏ�w&_nV���Wc�ƪʣx�n�+e�k��Ľ�;f�:�\I���v�������&Sx��+gl�����,>OHM�85�b�]�(�!�E��9�oV+Ѓ��&9N@�F��(�������=�O������5[�:��u�!��.s��`������ov�'C��Zw���pO/�	i�n�:�\��\��+��{*�f����x�X@�v���AW�a��230>|Br�4��U�tJ�E;�k\�ŷj��9���C��3�!b7�]�f ����fK��R�����Z�u�*ĭ�6̓������TWf�A�V�[}}]9�U�~̜A�b6N�Z<��� ��f�9h��-�y��
�T��Kʔ��M̝/k��ݚ|�܄��p����t�����O�|�:s��BI��ڱ�oH�-s(��"����Y����Ć����2ElU']�����2�n��l��v�����B^t���U}3J��a�x�4ǯ�mŬr޷5��vV[e�� �
>Ҧ�о��K���rM�+H�����>�_B�7��`����X����1�k�n�]��N��n�R,28��n��<�)���D�iln>�X9}��0��f�8��X����GV����3P`�A����9��E���6��XyS��|��6�b��ug,�5PfĴqf�ΚM�r�a@7Y�>Ի�\�nQ{(.��i>�:�����/��Ռ � �E���oiT�KlW���~�]�︂�y��$��T'�F��+=E�
M[r��i�ɔ�N���tq$%������u�k��0RG��ќ�nc�_[s���c�L���Qe��Ȟ�,Mԇ>K{�
}��[�}ļK�=w��m�q�2_���sUJ鳤N˅fȺ��ww6V���ۧvG��[Z�kk���խ���^ߺ�8��_��.���
�[�(A?p��F=���b�P1vM�Pܔ��c��O)HFJKn���*,�y5]^-��-\짵9�\�ڀ��OHUq��+8��wU�;ҎT9�74d��㿞dg����Xi �:�.���:���I�j:a�|�b�8�r�����v����sCTv�&��[a]�ae�/����=��.�4O��'�D�iWZoK6/t�I&h�8�u*�z��5c�εϢ�&�b�cW�B����`��
�p�ʺ,�x�a��V�/U�Q��\��z�YF�X�a\��X�P���6��'Ie�m@%��f�1,di�u���ҕ�C�����*��>9k��p�`dZ�Z���fm��^�����۲�_��1�I���1|��G���L
�N0����O���)�B���j�]%]��HG�2�Q]0��J�ھ�y{E�ݥ����3o�ۚ�;:���.P�� ���d��ʈ�g��s�f���<,M���p�o��Hil��n
,�뢊
�E% Pԣ���n蛸�`!��YR�*����*��	�.N��.#����7�:K�b|MTă�6�ˠ�V{��Y�v���&��H��B����1)�L0�񅘪$tJ� +nA��9�s��N�gXgM	���76��F�ԂwԎ�f�lτɴ��CH�N�6)�i�������NhX�-nZ!�B4�y|�Ǘt�Y�#�]7������A��n��p]���HbY��Cl�z,SS�e^6"��Y�16/AOEX� ���J�i%S4'�cN��m�ʏ��F�K^�tC�ɗ��+���[�e����mF�SW��7O� ѣ���+�E5����C�vT���>����ˠ&��Į�eH�N������C�IVfн��;[��Α�pQ�$U��e�f�����5É��A�;t�����9^��.Z����+�{+&��5b��
c&l�ۤ3-��%j�kf�*���@:U�u�Х��C��ƚ9;��+�o���vrn|0h��v	�f� 4b���\�#�����	���/��,A<h*Wv�9$������,�����!"�ˑ�iL�A��G~F�S��8!ү=�-�X��̨�� �$�+ih�o 7Hkǃ��뤝���7wfrq�+�
wEط�ܮn˛,0B��F�ܣ�3��9-��{Xx�¥���k�ʾ�}�Duk-� ��`�̪8�E��ͼ�-�8Tr�Y��\L��!a#!b��`�*|���O2�tH�f���Wk0!����/�X�[��0��(n�JEl�u!���Rǁ�\��=����^JU�MGQD,m�~��bw��v��h����v|*R:"�Vq�r��t��Pq�v�4�we���g1+�ZW�������vF��]^Ss�T�`�:n���\@TT�P�2��-CK%m ��U���lɿ�Zt^�	<Ӝ������-jsg�^p�6:eS:j{�H
ySv`��w":o�TQ��t���YͲR��Fj��]Ѓh�s]i�@��ز��m
�̻2�����M��)W'@�p!!�l��Yql�2&���ka� �a�����|o9ɑ�EN��[��XUqgZ���gJC6e��i�zX]�N�4��\�񫡯Qmݥ�촊����iV�^P�m�i����isI�d���q���b ���6�!�����"D��ӝ�9�Y�b�?���%u�%��p��|/qʗe9dcF�O-�Yڅ�0q^�9VK�w���\��@N��of��9f�ݰ�
�I:�2��@u^Uދ�YZlFd���+e���;��L�X�+��-2���R�
m�&��Y����7;��Np���iZ%䊳K�ut7�[�(��EK�Fh��c*d���k"�A�.Q9IS�[��+��Z͑՜f��uJBhm�F7�I�B��\C�Q���)��r:CH����mb����h;.�P������&��V*uo��ט%�W�.*����Uܱ(�,�3NN�?&Ӵ�]����j�u��Ö�}��a��;��v;71�T��`6[�r����x����HM_3��Z��L��fU�/�m�:c��Xd��G{bt�ݤ�ʻ`����b!��^���Y6hϋ�����#V�[X3qk���n����Z�xh<�r��q�3�0n<Y%��+����1���3�@o	6is�:X[�p20���kv�D�5R���h�2A`�$�Y�T��#FUبOG� :�/�ka�B\5���#I�MelD�	p���颯i<�[�n���;����Kΐ�׹��"�Ż+��c'��$'�*¥|�鏲t��F�mc�����c�78>Wk�;2�ǯ/��r^F)ܮe֛5	=@�}t�
s���n2;��K���ĔZ��,�mtk
�o52�?.����,�ϻA���\�d�����חCʛ(�DE������JE@HJ�J-���_�_.v)P9�A��Q�v������Y,Jx�0Z;�i�$�qbUEGnI-:�,������33�>Y	�w0t	Q�����c[�k�&��OI���9"g�*�_ ���T�mJ�ʍf�,�Gst��I�	�u�Z��	8a��ڣu+j�v�;���4z��a%�:���Z,�t��>[����H�(�s9RB�v� ��`p��B���ͻ�5���Kc�CG�w00v�h���Oz�I`�\r��#�������9h���;�T�~6m�l)NV,���oF9:j��Q]+8:۔���v�4����J�)LwK
���;v�2���(���A����;0�(�2��C����>�V-�U��577~C��Ϻd�����k�!�XlG�O���V��Z!_"�hiv�\]�%$��v�:��x��&�!��+�nwnV����(U����gF�n��٣�KAZإB�0����E����4hR�̺�%>[]8��0�����Ռ꺱�K��sȒ���L�|j#+���]��ݜ����*|B[�B�
��J����a���{�Cz>C����DR�r0^�R��u�������ɕu%�D�Vb�e�T���*I���9�JPYU� UMH��֖+.b̧i�9j�p�eGr�����m
�	ڕ"�;WZ��f�h��T��j͔��]�4oLEՑ.���6��[v������-GF,єB���vC�tciZRj �Bc��V�oB��6��{���iǖ�:�p�ԥ�}|����}���4��d����gUw�R�Q�b�;�wE�h?�[D�7�:�1�T�:�Gnn�̨�� 4�0W�j��}}@D��k�GK:v́�x%$Z%��]H������)��Y}�ɯ����]
th�"���p�e,�00)k�iF[�(WY��օ�
�˺�2���ahV!�<����->Y������ �+vsU��
$ϲ�ԩ.Ф"m�$�4�*
�����Iӷ��;(���#w*���(��⽧P���Pk���������R�+�ضY��S�E��+�k"e+��n@������ѺB]��βs%HYQ�^ږj}9��"�)&j,J�zSoAUض��B�]�,'�њUH�Ȳ�D�V�c-EBKYb�E�V@��S����Eh��2 �4���4��J"��j�	Y�����+:��-�D�k ,l��M�]�B7r[*���&4ʔ�J+�t�c�q�.�×J*���n�,s��j����o.cWSJ-�hw�+�{4+��:݆5��4�*����q�z��r��ڔY@!�»d�~���]�[�t�ʂ�zM6�\V�5k� ې��]�b�����A���2s�=�Wh;��E�s,�p�.�S�=�@,��䥼����ƙ5U�c�b�]&{}��μ}}��C��P�J�02h�f�lڇ�.��u��r��/qh�xRN^Ʃ���h��.���v�C�6x� �wD֒敢铷H�=�F;P��y7�����c���8�+B��{v�-�5Mg���}[of!�NW���W-�޵�	��[7�zn�;�Z�
�(��\@��i�PG.�pu�e-��,;��U�v�Ƈ�Z�����.�\폛�rkW±r��اBu;�N[�3�Y�p�X��t���-�1��w2�˕0���`|h�����s��z��:_oL�J����k����t�/,�B�����7m���nԲ�:��9ֈʲY
��B�]���+�-�s
'�d%����,[LA�2��L2P豥mu�b
(87zn ��^_}�N؝T �ƭ��^�Vul��=�3��&�7K�4t=�՛/���9X�-
;�R��ۊ�����㛷Gj.so��o:�_#�u�9�H�Eb����S���eC���6+(Y�0�=�V��3����_[dV���v�ei�@Y��=1_.�����̭8��Sem���{i,Lm-_^PWq�Z�%��*#��ڤ�	H�P�K�=̗f���:�=H��*�y�'|̺��;��Dy�3M%I0�n"'d�e^Ȧѓ���Ys�%5{&��nov��:���
�I% ���+�����k%�����bF;�Z�7b�]�CD\���vV������\�r��j�[�5�c����;)�X��C�ؽ��L��cU�t"�Giܺ�"�@һX� ��V
�U�c:-p�E+i9��
�ۡ�����F�3;��/�#�ΕM�7����Z�d��2�&)�o�����n�;�	=��y��-�i�I�E�E�� k�fKWJÃD��(ڒ�+�X�Z�@�W����Pڙ[T4v+�ya�s�$���`�]��E[I*m��e���Ph�$Sj�L���Ğ���`�*t��f�d���4U�]b� E����کW!�]�t�J�~P�ZvJ�o�r��:O�ۻ4�Y���]`\r��xMkl��24�e���i㱉��m��ɊpU�I�G{�XL�����=��G`D8㎃���=�f�v��}��+Y�@��TeQò����|�M36�=���
S��wJà!T5���\�E�Ub�Q���CJ�\��v��x�
6U�M_��';����K��RY7݀:`<�������E��(�˄��D<3N*%a��ԬP�9�	
�X����:�*���6���g��V�5����Wu֡���c�a��i;��2�cJ�����S�ͭ�F����1���z̖�*ҥ��� ���C���Xƞjc�(�H��ոo�a%BP��eh�
%5k(�de�*��run3}W�C-SiTm*YHDd���;]AA�+BU��F��1��N�Q&����z��0�Q�.��s+�ʚ��y�Ö���_r�vD�K����-�1��x=gY�>�=���Z%Z��7�F2g2*8*�ZvD5�+��Hi�y�x=�X5W*���v�Xh@Wn��Pj�<%m<&P΅ݜ�I �a��4��  ����ӵ��fս�t���AR#g�N���D)�U�����n(_,4�8)ǃp����tn.�N��󔶻�v�%ݙ�΄9�6�Ԕ��
�̂֬�c�١H��x�R�z��JTh�cq�p�i�?]#�n�_.C��#�֒,&S$��∗����w��Eb7YM$�Eh��V������e��4a57tV-�F0(�*�SB\(q���xR'H���`�~�x�J�.�[F/��b�Ԏ���0]'y���f���Qx y��Լe�R�-v�*W��"�����o/>�z
�,�HݫӰWB!j�8����ks��tqv�82�y/n����tP��Q����.���݁��kQP��w���*�X]��O�#J�v��PH�x�S3A��!�y[{hC�5�껦 2�D4U�2�Z܏��7��G��`H��4�*&ʆ�Ta���������|{��/�G�hs����i��g�QV��ט-F��2U+�׊��*�u6��c�m*�3W\�,B��l
]];Vc�j���W�K����n'[PƳ��yQoV��d�����,T֫����#q,Y��/D.��Zt-XM�5`�\�u�u�T�FP��Mӹ�ut-�RsA�Nd�삶����4��,6E�b�T �q����`����
W7@�����oY�3�8%ɺ��Ca�Bʅ����(�4�����& J+����D����x�Vw��E"n(�y;�t��]lWSr������w݅VH}v���*zz�!���B�ƻF'y�y�iuuwzŊq��])�ټe�a�#�qAf���;Ҁy(v�<0�[�L�t;���d.�ʥ���l6�jУBP�[���$]��(U�D���dU�Y�c�v2^�k��D�v%��A��K�kh[	pY�*��	&�B�����3��X�s{i��|.\K�N���}g �t�)+�55h��KU�zk�xTʾ<�n�aonU�É�0��)u��/iZ ӧhU��k]'u�Ka�S��]4iZ�mR�$\�lt^�U�1kK��q�h���h6h)�2�+(��2��A%{׸�q��b6@�*�=&��;J�]:�㏯�K�W&�BŇ����4��8>���R#��TKGAt-|F�]���S`N���L��#N
�s����7z�����h��Sf0\y�eX��ȞY[�������9���:J1��gv�~�������>�8uU�t���r��g�s�rt�;F�ݲ& �F�Oab��hrX������G�vX��Z^�C�6�~(�7f\c�1n��\ϸd?ve������R�r����[ɛ˔��㗸�s�.�^>|�k�sDa"��^��w1fv����Y4��>sZ�	���9,1�Tj��x���O�����m7�-;�,�j�Q���̊���]Ok�؅����\ʳ"��;��:�����f;j�����c��} ����ȟ��dÆ�@*�f�S�4/��$�NH�o����*�d3b=�rZ�32���S�E:�Ѵ�ڧ����\š3����$����LZRMΩ��ٷ��y����25��\�)v�?2۫!TοoK��i��٫a���6�ˣD`[=4^Xx1�pSkvK�ҋ�aŴ�`5����$� �X�B�]�jR/�c���I9���M5�tX�ڗ�e��]:o ]-�B�K�r��$�й�v�o~y�Wlo4�R�؆���C�қ]�ҧw�݊qM�p��0�R��W���8��;��e�imDG��؎���5��-���ݞV�'cU�,X*^s L��?���`��bVRo��iD���iF�>=�g{��%	��;�b��eLw�㷮o\o lf�&ά���\'$����u���S�<��4��[�����J}i�����W�o_9��_���F,L,L��	�LH@�ƌL �"1F
Lj,,�#*J�!��q��c&�LFi4e �+1��RbI*�&BAl�E���h�¤�b�H�d�Y2Y��Q�X��IJF"H"#d�F�1�@ı�6�,K�"�DjMq����58�A�$F��S"ضP��d��MEF���6E���ش%*#EA�2h�	59ˀ(�QX�EdQQE���llE-�ŉ5�B���cEHb�@)�j(� ƓQ�$���(�dIb�J$ء$�b6M�Hch�M	h��cX���4�F2��	I��(����2X�AI&Q�%cQI���D���LTI%b,�5d6ō��̣�U
�}g�����v){�|������WTl�dm��B���R���14i��},'�q��gZ�3y#�΀�Ɛ߾A����%�.�������χ=H/�WZ�HԺ�9�*���9��޿��p"Ͻ�5����pO���j�u��aX�~y����uѹ��7S}��r�I�/L��{�]��]��}����yTv9��:�!�<;�G�w�5k�dO��U��gs��.:�8�<|a�C�����󥖥��g��5l�*�u�%�f��:�A����J?8�'����G���c�g���Q�`lޑ7�+`��9EJ��3�F�'�4hŇ-�sXn*����|̌V���c;Ѝ�tF�R��'�^ɜ���ܣl�/x8��dpυx���#Nn��TX9ݏ�crEZ�n{~yLGF[\����ݦ-�D\;JV�{���Z� 8w�<�A�_V�ÓZa;9T.�.��9�V�j=�uz�;3�_;�ԡ�{��Ȍ�	�sfP�B��ꑆ2�)ؼt��L�F�N�����Ȇ^�p�{Q��6����x�A�D�
���\��������w~���8
�̀*���>�6>S�`b�(��b�|*h�`��Wfv�Jm���K7��lXIXL��*+yQպWgS�_uΛs�}�ԑ�i��}�(q^��T([IjҒ;"�ܣPkJ�b��-Wf�cg�	N�g6T��v��}�{w�b.�W9'ܵ����N�9N~ʇ0�*�RQ��sPA�k*�}ܤ1�gy��F��Z^�,�pV�y���6�����:�n��ف��i�	K)�{VBOV��cy8����&'������wm@rj��&,"r�F�-�Y��޹Γr׎^U�1�M<c��~�#Il�=])���1P�
��J��=�Ũ��:��<���jTS���6�:`�X
�I�<O����G��r����f��"V*d� h�������?jW6��n��w�H'�j�+Uq�ͮǄ�����9"�+�Һ�^�IGbFm�CѮ��ԙ(F>�:])[:GK�Do��L����օ	�׺�[w�M-���C���
�U���l��ɠ�9{qڤq�q��YV(s��)� 8��O8�]�5�q�J�����5���atO��srpk�c��q��N��h��86���09�^��=�g>x�ՋI̔Um�yW��`ό�d�I|�܎W0�5Dl {@���1VW,�jq��αإ��W������V�9����~�TT$'���1�}��a\�t%g�b�[i�|���kj&�Q�o�¯_48`Sz�<�q��gYǀ�v�!o�H*�q�/ G�^�m�`�U�z��;^h|�M������z��F��z^Z!G��	z̕�7g�d� v����.�5.�r�7��� �V����^Z+2W�h_LQ�"M�҂X:do�Rmw1g��3}.��=]�r׫R�q��nD���6zg�`E�8(�t�q�\�ѣҶ�������q��	�/��{,0}j��_�2��p�8�m\>�8���&VJ�{yOT��Cn�yI����/��rBjP�[S���-T���9�4c>�#�Ϊ;�d��O-�]3E���-�0\�.}�¡M�@��a���M�k늸�n�u/�X`덄�py!�Ƿ�OCڵa�L�e��S%MG1!��J�qx�O�Ɩ��,�ѝNngF��i!,#��a1���	��2�����'���q��w��z�i���\���g/$�r��;a�yȌ�7��0��b���%�#Z4�dd#H&9���LVr�l��[}|�h�*���$4Xzb���7���1\��D�Q�C"������^�7�lYh��R���Ľ��P�����s��|����
s��99bV��),B�dM���H����^��?�C1K�Mp�{Ye6Î�o؂��>U蔴X�s׮�5��yVOu����N��m���z(�,V Cz{���[�k .�9wֶ����*K�lC��2r�<�eNߗ�&dܟ �]Sá��_�R�ܞ�$<R�؏�{cٖ=K ���c��HMu�)��v~��=fuS-t�d}l��j����X4>��H/�cB��&�0oG1�+^��+�eL����שza�*3Ų��(�tˎ��#|�箴w�K��cЪ?����2�[��>*5�	���kKH�vV�Y�0����l&�����{��`����u�A'�̘w�I��e��(�u=A)�;,cj��<��g� �ݵY�+���!��hV�D�Ě=��54$L��RX��tY��VF�__Z�LBe��-�K��T5<d����(�%��b��^�QZ�%VF��X���wH+�A�i����^۾|[��V�>����(&��x�6r, V+�=/�-�H.�\LS"m�z�V�V\�����-�Lnb廥���]���{5!{\����z�� �jJ`)�>Б]�ڱ�Y��>�C�ꒄk�ut�貺������S;h�q�ƚ�hb
�#�WJ�9�rX��5�	�|�^�޾Ra����F�YW9i�^��Ɉҩ��1Gi`VQC��qgSz֕��cS{(��H��t.�Z77��R���v(�]�L�˃N7y�L�1�Z|[�́30�i�nH����sH�)�DOAz�]?JU�,5To���2�M�6����6!�c���p�N�1���G>-U�~��+�^(g${�-}�Q1��yE�Gkw�4t�o:h\m��6a����*p6�c (a��T+W遶���WT�L�^e4j�![T6U�ip�1�jY��D�1��ܕ0ZX�MF^5����9]\�,A��p��Ga��-{g0��j�B�s�c!�WD�CV�oA��OWt��Wx@A����#�b����d����FxŻ��iphjU.��u��=]��Ř�yfƙ������pP�yv.8���G7(ta��.�������t��=��N@���ќQ�򪇂7|�j�+W��E�A��.�b��
7Mo,�1�!D��zO�K���@^�p���+�#�����nE5A[K�q���'�H��^p�#9��dD�P��p�X�Sf��PX����W��ȅi���Sgr�ۧ�ynv{2�u���i�Z�ɱ/᣺�u�+F�	�k���N����5Ժ՚�
c�l���t�b��v�B�p�;�.�����c`Xca�	h���hv��jV!�����������j��%<	=��.V+��ý��5
Y��%�R٥�+H��� »��&�h͹�]�KW����7B�J����̙��6Usu҇z�ѯ<r=׹�d��K_t���#B��x������ב��\P�
��ם��h�C�[֧mwY�=r��3�4չܬ��2Q�Hn*��K�}��ri<�Y(G�=�����4�4ӷ�#��_�?!���m�� @A;�*ld5����B��B���C�j��eߪ[$r�]�Qv�[sB�RQ힂_q�?�V�U�r�����#I�9
鋈Z裏=M���ӝ�n��1��3t�׃V�)���M�����ԅY
��చKy�3�ثG���;��r}\n�1�cV�զNu-��9�$q>��N�������"˱��ORG�9_�W��
��.�F<�6�w�|�$�I��@�� hB(2��GJ'�@��tu|;�mV��=Ԑw�͓P�hD��R%^�}�O�6�*nR`Ѹm���v�p�$�t�=5��B(1c��%h!i�����Pz2X�CO��#�}�J����ծ5(Kd�U�B"N���[�tk{۽��]����.�5�}spo]�M���u�
9��^�>�g/�hn���|�3GS�4WV0c��hn�@�'>�{g9�2�G5U�����(�,�%3y��\�F�-�ᅐ�%�>�:\�v۽�q��< ����#����v��Q�UGS���c+�i1�Pj�3�����u��4������V�a���2��a7Ox8�
�z8�+ʢF`�&�%/���]C����|�s?H �\�ܞ\��azR䤽C�}��	����QU�Y�?�(��)w�ۤG &�s�'4m��P�j�wi�ks*7����qM�=+m`T�h�O��K��
ێ<Y6_TC@˵Al�O]��]Y2(<K���_l<���<#v��0�l_ӑ&�Q:<�%��ٷQ�e��]bx�v�nZ��˹�����nAe���M��e�i����f�$�םݎ\�T��G5�f�s�@?H37�l����Qr5;s�����G9�p�>3����ORٸ�T����E��ՀS2L �;����w]���/:nJ�s�y�##]N07y�RJ��3���U�u�[@��.����P>��f��U��#�Y�W�)o�S�ޕ�-�.�ᅇX,�]~�WN�^S�t�{��*��J��7��3+tv�a�g�׿]�#�P���#M�	0={��:�v�q��H��_7״x��e�9�;�Vf9ŭ}�wcw�˺���b�]��fwQ�����NiYht|f,Z�[ۡ�ի{�ꥳw���&��0��'!L�5� �TK� ����=��׷�V�G=/Nn���ȯ�wRg!����A{X�&�@��͈(�W�R�����3�7�Z�����%bER���tkS7x�����s!��3l���h��̊F�)V�9c)���zkX�g�秊-D��	��L_t�+����2a��;4u�ME綞
�{٢U�*�6�����޽�W��k����UU[��2T�.'�O�dܔ˪�7Nd�l.�d������I�R>y�RGK'�>��<$m�0���s�}9f��r�s<z�'���I�7/��ɘ8��,/�4��=c������;~��c#:S$<��k�R�M���V��mhp&J�3����wPr�����_	���?b�Ř���)v�Eg�](���j�#����Wi�D��SG�f>��V�� �fu�6�GW^&Q�q��	
9��T���J�S�e���Er�a��f���7O��ɹ6��R�� 4��R�uc�V(���ƽ�"=�b˥�nn�l�V^��\�E�Jj�)ԋ������o�y���ן����wSm�a�IGT�Wһa��L�}Y�`Lx@�F��p+=�Ń�S[� -r�{o��W�)gJc{�������ǮbQ��#�m!G=�Z#Y�b��J�+>���.���:b.��g��K��7�]I�z_c5�(W��\X�+,��QZ�L��򿄇�k��������k��8�TwQ�쵷+���r��8qܭ�c�����"�!u�K7���� �	���y_�'p&.
\��|��9�l�n��$���@���$)�"�(��& �?2��zG{x�bC��N%�Gc��rDm[vF_�iD�"��#�TE;���a"�m�_������5���dJvٌ�oe���`��EwlT�*���-	ә֎#�4��s2+�q䉉+�п��C���z}���S��C1h�b�a��ޣB��J�
�}h]�.'f��Ⱥ.��4�E�,��"\�K�rT�x��Ur�s����/*�♲�L'�A����2���WV��0�O6k���������L��2���s �%��(���	�ЎՋ���&:Y=r<�N��w�����x��>�t�;Whh�eզ�c`�o1ǆ��u�Mt .�'Wu�v�}׷ۙ�(C\�J�v�R��Hyi\�ѹ)�sm&�KyΙҭ��l�D>�Y�WT��4�����q�|(�X��8��3LY�S�����r�Q���PU����J�����e�<WP�w�й�˾��϶��&8=��!�t�Hl��]��Л\�Z�6�7�u��z��`p����(��UC����Z&�w��0Y���5��AgE��+�����Pl����|�&����uׂ�n�]/n?��nE5AO]Hl�6�OG,6^����W3�V��v��N�/�X�ޛ���O���}t(]R��93{��Wz;�_).�~�,9�?��}'s�_�G ;�]P�al�[���ۢ!r��k�Vc���H���E�ug�_��[�{�i|s��G|Y\�x�y��x��ُ5gh^��W��g��f�#�B��=��^f1r�1�����c��ɔ��	���x���ڦ�L��4cC�s��X�:�==�2��i���p���@�����!�b0�^r�{w�w �[�Rc���˿U�6:rO�����r4��Kc0�(U�̌Xo��3JC�(��:*���I���S������vz)�|bY�s��p�f���4`>B��l-�>�L�U��t��cuH�cx$��ӷ������im�/�.�ת�d&�Ÿwb�
�����IѴۮ
�K��ޝ�VWU�>�Nww{7S�fT�;�a��)�Ml
&�L�9=N��(���(ix�˜�����V�����c:��#�SD���y���]a�Qut��d�y�3nY���t����f� /��Q���1$�9n��T����>������9c�����<aW�2���Ű\�`�:X�z�H��\�m`��,��	}	�y)j*rㆺ�v�!Enn��j<��/1N�fn��9���&32"3�m�WZ[�f��B���D �_5#���|kya<�ϭ;�.]i�f����[�-�\J��}w�2F�9�<�[C��!^Ӌ4n�Ze��2�7ն�N9���^�b�noB��n��P�Q�¥j���*]�9��Ճ'`��(*�b�@��-����o��Vp������=�q�
<��}+qad;�+S�¶!��� �Q]���/ni����k+�����k�V��g�D2arr:���܎�[�B��8���0N�$���ĭ7�m��g�=7ϛ̨-��c�et�c��#��.)WLK��M�x��`�A,��]�j�R|��uv�U�n�,���}ƺ�(��O$m�Br�����\�i���v�|aY�)�;��:Fm�c�1R:j�P���.�K���t�ǣd<̭�E���,�y��R�.w�u<�zn�D6�/��V�LC����:݆]^�Je��C�M�����G�e�h�u��.��Y@�*�{*8����t��ͤܢuS�@�,l��'sz��vt=yd3��[�kj�ק#$j�d�A^NP]	S���h���n<�Rh�z1�Q�z���h5p��@�l�j?}x�ko�m��x����!v�'��Z$��d
T��r�2a�QRc�����E�݉�/�ӷw��OY��Q��fm�So#���grp:�
:��VB0��aַ�d%)p�Rv.��� �s$�����kV�l�ٗ��S�;;O	�S�U:��Y�P�����;�c�2��������h�t�mg
�M�h�X�"��۝Z����5�V���QeD�����W)Ls�p=1��0nְɫ;]4K5)���ܩ���Ŝ�-V����m	�b딝�d�p9ػ+[)�N��	���7/A�7�{.��n\��"���c����;w��[c�ܼu���mUEX$�C�R�����sȠdX��ݼQ]�v�\�cCpW�j��W��xg#�\U�'&���ӏ�٣�ESN��7+i�R�o��`n婖�ŷ�>/5�[a���x��Y���߹+��A�Օ����Շ+����Hκҫ�Y�4�z���y��nV�S&iޓ���>�C�>�|��c1Ih��I,�$�4��AF�$cX��!�j4L2l6Z2�đ�QHd�X�1��ABc
���F�أDA�4M��&h�1d���I�(f����X"+��ARV+&� b	���`�5�lEmA(BJ(��I%���ZA+X���U%�KL�A�IHQ$h�ZLlh�HfcAh��%�54Z
�J� �#F4��I,RcQ�&�+*I� V,F�ōd�DQh�TQ���%�,`��#m�QX�h���X����E�(�̨ъ ѱ�J�VLj�ԛ@h1QEDTX�4X�Q�I�s�;���^��Q��5*�k��n2�k�Ѽ61 �żf���֙h�ӊ-|��E�ܝ/�f���ػ��� ��B�Wm� X7���]�����~����n����k���h.�s]"��+���y]s���?+��]�6�t�ww�����[ҺW�ﾭؾ�眷��+���/;���q�#����t\}��� }}�_k�"m^�w�}~�ߗ�z}m��[˟��[ڸ�ۥ׫�z��6�9�W���ѻ_:�r�:c}k��]E�~�t�u��n��7u�z^-�t���ޫ���5�B#��'8#� �#�����{��ͭ�j��'�0@�E���}�L}�^y׋�}mι�Y�;[�q�۟������-�\\n�r�=~�WMڽ_y�U�Ӧ�;��6�ߗ�����C�z�� |h�s�)ԶC�X*�k^g�Ӵ�G� t|��*���o���7���w�+��k����ץ�W�~��ܷ��t�ۧ�<�o���׏����oj�oy�?��K��n��v��Λ}]�[�6�W�ɮu�{�㶨�⩕�y��^��">C�g�\��t5=W����=��\����7�:k��������o�_�y��o��h���}�Ex�WM��m��Z�t�_)����\~*>z~�Id �v��̩��y芢�SPk�0D@1���/j�i�/��r�o��U�r_�:om���}�+��n�B��s]-�Dx}󞺉�Ax}��뿾�B4G��׻��9oΘߛ�|��5��_?����.�(�q��G-�9���|���0쎁�ץ��˥{�9n���]/���u�v��]�?��WKOܽ���ǋ�n��뮫��6�\�����[�ߕ��nz���צ��+��~�����-�nל�w�^�9�]ҡN���������Wm���.��u���߾o��]��|���+�����|W�r�hߕ�qxߕ��o�|�����ŽW]�]��WK�տ����ˍq�-��.9*��X���֊���#�#�W��}[��6��[��;�������ߟ�ߛzU�r^��5�ݷ��k����6�z�˥�7N��\�绾j�-��]r�/KF����}^/m{zWMG�X�ѧ-�z\��}Afט"(��^#�c톓��|�(���_K}�u�-��^u�h/s�/~w�}W�9|o~r���w�k�n�7�n{����v�K�w�6�o���sk}��N���,�Wګ.�i��R�^����x%Ὗ�'���]���Z:�{Iօ�#!�F�۲+��^��eI.Z��ʺ[r��#��ݤ�d�ڻ/*}�+�I/�=|���٘��aw���_ڷ���<.�����T�4N{*�|�'�pR�g��$[Y]������-q����.���^�kG�ﾯz�-ۦ7�����h��:����뚾����]/�]=��:��x�k��y��{Z+�{����t���u���!��>��
Oj�us�WWsj:��7�n7���j�ط[��U_U��﫶ߝ���=u����.��Wmn.����{~Uz���_������r�_[.������Gr�4���Ds�sw���{��m�|WKE��+Ҹ��q_��[�t�x�7J�\k�|�:�������\_z�]?6��k��=+��|��_�����U�s���]��q��q��|�lL��G�ʐ��y3Wzs�᝕L^��}t�����Ϝ���o�O_y^����o½.���]-��r�����v���\]���oO��]+�31�/��c��s��� ��7��!�>�f0��\1U�`3����;͇����}�;���oK����M�ן�����q��K��:���W�ƻ]��7m��ܮ���?.�z�˦�ns����r���_�r�7����󮫶�����}�8�=��OWHkYs��-�-��]/?�y�q^����~�z~k�m��}n��\X�xۯ��6�\���{[��^���~�k�t��˵�n�~徫�m�U���|�M��">�Vxm���ǻ��zeZ��	c���.�M~k�^W�]v����WŹ����~W�Ҽ������h���}����oJ���λ[긷���םU߾[�t�x���]kү�Ƹ�_��^ߖ�&� ��A���
>�NC������R�������@�E�����*>���ֻ�����q�mǭ﮵�\�;7M��P>��!@���%�1�@�����T}+���}������zWJ�y�V�R@��_T�Y�7��;��BZ��ML�tzُ�&�&>�@P� Q�G��h��s�����t��ί���n7���ֿ/K��7����u�-�}ޤ*� }���s��菁��r�}�'�(E��V��i�>�m��W�lָ�1�Ę�D��.�h��#���?�^������-�~]5��׫��]���׾w��_��z���ݿ��WM{���]��qc����yzU��6.�}��G�|=� hۺ��|<+4�.�-r�������VC�uw���b٦��u�sh�smgr�;hG-S����w�5���h���N<�����u��h���45�3���%%��2�T烺�ֻ�A�T6���t��h�P��8�����f+�4���Q.c=�� ������*��_�}u����ˍ�t�t���F������mpk����o˥ҿ��\�^�k��^7K��.֍�����ޛ����{��[���qo�s�������J�B�X�i*v��ep�w�@
�~���oj�\k�s���K��ߝ�����W���6���}�{W��\�^�^צ�mž/Sn��鯋��+�som�F��
�\(�D8p����>WV:-�ǚ���V��h������}z��Mt�]/���Uv6"������kO9����[�~x�Ot���7�9�_ܾ~���kA}^��5߾[�TO9zm��͹����]��:o�3ݱ=��~>��]`�r
���G�"���.�cQo����^�[{]|�9�/w�m��v��_:�m�ns��|�opU���[���뗞�Wm�x�K�~޻�}\Z7��{���+�Z{���E��[c�Ȫ~��1���:o9͟y\X��\k�_��Eι�6�oþ]6��q��~z�~W��ߝ~忹����{m�_��:�M7q���^/Mx��~�v���Ҿ��F@@d��[�m�:�}�c�#�/.�ڿ��t�^���U�ޛ��]5���t5�qo��\ŧ�[�u�]>��W�����W��/�Kx��������m�߻���\Z~��޼�o��ۍ��'�	Îk�Q��]���t�C�>����ޫ��W?so����5�>��{W9k��kӦ�o�����n��].����]s��؋�s���Z~���~�0�}!��_|�T`�����׼�d�	�*�=�:��� L�D@k}?}O��WKy��m�����������o���������W��W��j-���t�ۥ��j����s������wʺo͹�Q~t���z���_���^�F���O�����>��jG����_}~��W��z^n��q}W�t������n>��]^yݮ��qc��{��������o~r�����Kv�oܻj|d��@��D�#b(�BK�z�D��.��UU���|D}�1�E��4n-���]��}]5����]T[�}]+����v�����U��:ޕ�]-<u��W��o��mםU�����8�|!�@��"�T8�� 	�rs�N*���^�UꇻS�.@�8�K�.�D,�b��1��G���@ ��c�$3�U=&�]� c�9Or�ū�k���I�.� R����$Z� �Q��j��Z�W�1�M�����U������f	�oe���͘�;X�gǩK�C�p{e�뷅���;?}H}^�O�zv�n��+����z�r��[�qW}���x���6����[~^��7��s�V�o�9��}�pj-���ץ�W>��?s��^��.��9�zk�(�(�=��Lm9�FY��,���Z�羫��^���z���m���>(�.����5�s�yo�t�z���ny�v��߮m��_[t7m��ޫүˋ���>���tۋx�=�Ͻ��v5yX��>��<��Z�����E�>�E׾l���}m�so�痮��ѽ��9w��������k��u��+�9�ߗƺ�/��Z7���Wֽ/������=����n>5���|�������ۼi��psk\�˽�.�X�������w��|ޛt����;�����8���v����o����s_��6�s����F��}n��t�k꿹Ά�ߗ����/���\o�߮^7�|W����(C͕�]�Լ�:|�~���H����V��W�o:������{�������ۥ_���;�5Ƹ�z[����Z��-��y���-�\[�����|m����ɷ�����ݭ�\��-z�cvW�"�h��Q�DG�D��G�K}W?�k��ߖ�鮛��}����Ƽ]5�������{��}�x�����wk���n�W���Z������߾[�U�~�н��\��t�|��x��u�l*T��<bG�H��L|E�q+��o�m�ۋx���;6��(J@8 Ï�Pl�G��}aŇ4���u:�d'V;���9{�����VF����針�,� ]�l@��
���T_0<'�� ���|P��w���[OExaZ;
~�{�)�~�����N����Ҿ�U��E�d�u���#Kk��8�٫J�-�ud}ͽ$<7����i��z��nT��>$��w��W?�5^F�=Ǹ�1��P**癍�͘1���OJ9�v�U��M�g���
��+��ݶ)���l}�Y�����	A�p!�y�����\|�X�J���H��y�3t�֏���ےPȳH<��Ee�	�	��1r�`ܙ�T�FT�5\���u�c#V_u�٨�ށ�5G��j���8{U>Ԯ�9xTi����0_J�+GX6LO�߳:�R�=j��&�R�o�jq`����WAQ��|�&�R��#��_��������ôR�-e69oS Pd�3q�y������Xlt���k��u:;��wo����{#�^M�e��0����z���I���S��Z熎�[W�i�.q<��O[¶�X�7|�f�q��V�;�XM*[��ثG��m>5]]��^Y��)+e[�:;��3Զ��`qU2b�5�n�n�t�b:'���&�m�/�!�踼"��Zͱ]���TcsJjt���5 U��)�Z���|�GWў��Wx�R��pnt�\�m��66���|�z|[WS~YI�`��g����� �uBPj���'��g�B�É�2�����.oD,�G,��(F>�:ґ��X���]Y�+�th��F��g|�]�"�W���+�+ݝ�
L ��a���O�9c��������=�����f�g��Hz4.��c]�۩D��#{�-~N��!����8�٬��Ü��Yw6 i�v�쬹��e:���~��"��v�F)��8�+��Qs�!5n�N�M�Ov/�h�M���]wm];�{����ݚ���X��eB��#�t�!<�[+�������[� ���XHWܯatO������^3��m�>ăgu:y�^��O��0�\�ܯW��	>���B����?�VK�N��Ԓ})c�+-�ӶgR[`��kVH�f��:�-�Ҿ�=��~���"�������V�v�8m���� h��D$�(�����x|珝t���;����d�@�WoZ���d����m������5R�y�i�y���z��Ӗ�t��8y孙��p��J�uq�/�N0P�E��T@W�tÛ���lg�e�Z�����k�|,x7qf]b�����^�)w�)����^�|�_i�'Y\�w|���Wq��Q-Ӿ;�R��s#�*�9����5^���-r���ʞ�F�W�nJ1��3�I�G2�"��R|V��r���I{̗�9�m�u�Ò��u����9�6�R�*x ���� �N�p��s\�#yhפ�s��.��+�NR)�������n��6 �I\rJEutng;ʑ�gi���4㠼}>y!>��G��ξ&u�3�k(�􏥚�xop4�l.J]����Ե0vvV%y^eșS�|�ӸB��|���^ݾ@���8�b��ά�{8�l��|�;x�.`�z���T�3���/F� �ۮ���9�*�\e���>���nw��"Q���H�݁�ٿ��1��.�FӘ�ŇE�����EUT�4��ma�[�����VW�2� ���1�t�W>��m-˝�e�MЎiر��Dkgڨ���έp�]��oUͥ�l�^�']�mĆD\R댓���*v��)6أ�N����nZw��y�`r[�Oo+��:�A�\N�Z�sع]�iz��H}n��7�>�j���܉r��W��g�(Θ�;`.���@�!�R�O�p
���a��5�}��F��9�o��ngG5ц���f����c L��e9��{}j��yQ�b�l�'��A�ֈu��F(�6+�Z��|.�#�ۆ�]���4����Q�~�dՊ#�v5iY�ǭ"�{�[���xڳ�*N|vX
�mC\��`�;���5��0��i�R{�=�L��W
5���`Δ,T�#eHEp�V�a��:��+V.�� Q&�o��v�t���չ}�+8B�T��;P<���𕑽~WBC�5� �)zɆ�$�]�3j��+<���)��;�f���w�\�ڱӎX��Y7�L<�V�k̆�S�n�RB�v��̹�{JưpݙMo	GTg8=�T�l��J\�5�z�i�ed�W!>Ru!��s��X9_LK]��]���Ժ^��>�>�������j�T�!�Q0�^:m�|�5��$��|H�\��� �fw�iL�}�9���܉��s���OG9��:i���H�3��h���鯤�2��U�Q��y����EoB5oj���m\U���#vnH���쌿��3_)�G�;�^�����.����N9�"eu|+��B��з��b�m��6Z8\�
M��mL�$gT�>w�,�eGbF�P2�ٌFr顝j���
Xv��˩�ՖK�z��m�V��-�g{�j� }��d��i�9�*�J���4py"�4�������<4�ڧe=/ynX����d�e��Q`O��Q;@�Zn[[Y�[	��[��){>�C��Nc��#w��6�]�Sr���ڱa��OK'�����rI�\�}I�y��l�FB��o��U7�p�&N�\�eڬ�}��&8=��!�t�����l�t�3}�`�Xju�#��s�8��8dGu&qG�T<c��alCD�q��h����6)��c@��g�k��TrG=�N�w��}K�UΘ �dG�H9s�Jl��Vh�!NWJ���;��=2u���7B�S����-��������:����:�B�����*뿆��^�sxC�c�5�{��W_4�;iu7�!�������z��I䃍��8ɇ+=9Y(���"ON_m *���1�+�#N��`w�U[��ex��;�^�}5xV����>�@]�*�!^��Ӊم��U��;g�X��{�c��֒b��I��"W��U���3���-�,q>�~ch�u����'0;������o�2;��+�O���*�����si�O�_ԭ��#B�\I�F��\�����/0������mB�؇!�ZɅ�������/��l@j��5����
A9���8=;�"���g@=Bc�q�T�1�+�,�C,P�J��d2��>S��)> ��*t�K�ヮI7���Y�� `��<�Ɣ�ܶ��n����c�:�.9��ݷ���fs�Oh�����vpF1Rx� ;�� �ZH�y��D/����%�q�ѮP���Yܚ)Ӿ]:mm��)��� �&`p�ǲ�� ������c��
�S��Y֣՗�ޣz��A�r�r������u�\<w 3����Vˣ�P����xM6@�3���
� 8��lnq계����[+a�i��.�.0M�@0so���ʘt���y٨�;��:Ђe�-�۷�1��t�>�R��rK;�0�g���6�z��l�%��ɰbҷ���ϕN�����WwK�[ݜ�W����}�W�Q�Ge�
���#��w���������p/� �p�X
eI���D� ��w/ޠV�� ���}�	k�;��=�_�I��m��K%2h�6�leP؂��Y�G��������3/D�q*L��v^[���j��p��I��dC��ɨ�(�5�
0r�6�qUV �Q����{
�8��U�X�F�f����&:���7�?Oo��¡�ylۣo:�Y����
����u�v�,����n i��3�U�+�W�֬(���=����6{tէ7YG��Y�§08ܯuSg�H��P�Xj�~�J��95����>�Iw���=X%L�x��9�j ïb�0Ҿ�>쭽��`���z�EnXK_E˼�-^��c21��M���>��r���}�x|珝t��w5�hd�Wrj��lj�����IN��%q�2�zP�8��q]�hv�2��S���e�n�$�wQُ�j)j� �d�B�{Deh8W	X���uSm�+� n���s��ڜ~��}r�+.���7�H��/1an
Mo�ky9zw��G��[u4�q.R�:�ص�ST��W�s@��o"i��<�FZN�)��jՊ��:S�[���M��*PJ��h�i$H��Cj.S,墲<��{S��ꕱi�%i�tm��E(�������u\疕����Wx���U'G{�bD⺺���o�[j�r�>�:�Vh�D����_�hu�}u n�P��w��+@8�G&V�X�S��nmeJe�KVst�4����3xw���֢2�YaN��`Ħ���d���QV72���(�ZK,f=��T�][�D��n����z���IN�.����<���6��Cb|k�	�9��\�S��U9�[��O.�^���+;��G
s^ӸfT)�T���uc�o ]�WFgn�.o{ϯ��"`l1M�)�j�G;^�1LcL� nv���[�%ߔo(�7;�����>�	H�k�V��w�L��;f���╍�[��Vm�k(RI����l��o\�F'�}y����i���wa�K�Z��cT�P}��֍]�]	F�h�1�tU�+4P�9�$k3����&~F*̊Y�PCy�-Od�bɵ�}��F��a˭�qFm�q�����xLn���VP޺"�S�Rg����Ѻ }[�����S��f�$�ۖӾ���qrIH�v��wv�Y�J�����XS�B�R�<ޙ���^����FkGhM ���7(���vP�w{E@��V�%&��kI��������)p�^�6���:�`�X�L�<lN-�m��J��9��f���ء(��f�2'�&�yS{�wo��ܚ`�����u�i��/F�
:�Q�'3 5�(%!���+�7��/9�=	�v�j�)#��,6p�Iٻu�S;m����sI����F�������y�$�[�2�=���CS���@�ڜ�U�3qp�LE`J����)�����س+uTl�N�7�Eh͕2� us����&��źbT�.�W�Eo�c)�����u%�lm�σ���V��2R+P㏒��]��=X�t���k vyYu*a�3�Q�n��_Ċ���C$��yOq�:C���;�8���[���`�+w͋�^.R�Δ�]�<�6ORŦ�����v��J���^n�W)�p�>�;���꒟P�&J�(�J��Ӷ8vsx5�&��eb鈜��Oץ�sxF�@X^���^*�i�o�d�ɐ�F��w6�IQӱEn��h;+��V��2Y�Y�{�kj�!��Z����q1��s�ɛ ��w�r�A�z�'��P������iw9���$i�,r���z�l��촹g@�s꿲�p�#�Y�k�5�:����@��2����t�7X�� �OB{���J��kX��)�]�g,s6���K]k��.fR�2���Ư]�bJ�]�p�f9���Tyq�fV�n�ӷ���X��F�Dj���cDE����)���*����(�K�l[�T$b6ѱfcE��m T�h�6��*�Z(�(�i"���h��Q�- ��E�&LX�d��63M�clh�I�j*LcQ�ƓX�e���F#mdD��i,ȓE�F*(���Qd�4h�)6�(آ��ccF�(6Q�Q�R����kE�E�ѴX(*H�%��_�{���խO@���}2�VN�;*ݮ����J�+�
�ǫ4�����j��<��8Ft F{.���͜и�}��U�}�"|�����#5"�}��Z�|I�Ep
���BjU�{��?L�3��GW���
���{�
M�����j��4�>�P��� �U��62r{�����'���ŚL�I�����ю�gmݩ��T_	�B*"\��Cv��C �@�gQ{��з�}Q�$q����y6����sb%q����YQ��P����,�3O��|tn�:S67���������p�4�}� 5gL�]�N�^���ErBuN��z`i�(��*�A�<7L��go��Z4�ZdX�/�����:��|8�6UiQ|4ȩ��&t�:,�� �?/l���?aw���l�px�+M�r\���U�Zo.���S4��	������ו �π��������D(s��3
�Idz�k4qmvR��bڪb�֖.F�"����L_� 2��ݸEf�;{H�3ug��[<�8P�2Lb���ٷ��@!♴���;�9��Tw��Z���$�?o���a���$���+`���.R�,��8�P�(��hi�g���)�aż�glIaz9u-����=���\v�:�Vu&*X�w��:鴙Od`K�8��퐵����e;.��ѳ:���w;$�n�)\������}�U}�w����Ֆ�W�,8eo�� 6�\5U� ��SG�c���;]�i�{"�����WV�]~O�d�@}�T���4�59vX
��1��`�ޏ�u5\�ѭ��v带xy����ޚv`6]
�]������G>c����,�.�yܘX�.��;Y��P��*j]yL�"�l�D1A]g���w�}Ek�-~[BC�A�/@���d�ް��
���3���Nw2��g�A�5��M� �E�_U��T%K���s��_#�gӮ�^�]���
���)vw��co ��ީ*��	'ej {U�f�[؏g��a�8ngy���j:b�Ӓ�em���Z1f��p!T1�[$Fu�de��f���j�G:��e�m��pE�S�An~6S(FB1�ioWR�����`��P����j�j��g��T���o�L�Q#R=�Pj~Ud��$��}j���Xk�<>ʎ\\�gt�:�Y��0���D���Q>���\�R�j�q���lӤpy.]ԥ��lOZ��]+ٺ�(-̊Pb�J��ɥ}�i�Y&�]t����Z�4qMל��n�ڭ��l��9tgP���`�VL�R����|�h�)gS�E��/T��ߒ�~�9wE�S5�׼t�u���֘��ֆ.6�u�Di�"nj��Ղ�@�z�R��}Q�z1��=��1���;���l9�E@w�KO��P�3��t�v��\�{]-��wc�;��B.1�p���m���]�T7,/!���*�W��݇j�����^��YM70�/Փ"���Rmm�ۨ����`s�>�]͇��%�|d{�)�<�F�	ս*�������G�r���8gu&g||����n��^����)�87yMg��n,0S�V&�ѭ��*��~h��7+q�g�����}p�c�E�5�6��Iʇ=�4�f����_���q�$\�i��q;7� ��0 +�j�����N��Ilݜ�R��>��v�܄o۠�5��Õ�} +��$j�F���9���U�9d�+J�}��GZ�mnu�@��c��\��)E�/p��=PP��Y9ˆ��5*sg�p�c��S�\-D��pv�dh�����ί�k�W�Q��}k��˓�ĺ|{!�s8�u�ec�\�f�e�Q�[�s�΋�?pʅ�q�&�JGsK�+':�.��ؙ�O)�D��c�$*�o� w�eGĚ�8e�s�@��.L��*q��M%�F�n+P#�
��n�g��<Nme>��ƱN�,7���T��:	ԛ*WL�#��;�:u%3�,u�!d�tq�çGx@�
� %58�AQ5�ވ�G�)��8��9Jx���f����
<�����-��1�~�����1�YH6ȷpN+��L�����k��ѯI��1�B��%�prG}&�+��P:#�k�2�k�X�SJ^�ڣ��nP܄븜n���,�?#�T'I��z��r���7�ΐ��:��K��5cMR��a�b�&�mցo�т�t�8vH�$⠮�.�*	�[���v�G+����Te�%P��n��� `�L�o�N�W���+D��=^�*18TF�pn~�<�I��Q�+Os����M��Lw3�!�&@�Z�}V��{~�O=��H�i��t�W]��쵥��mB�z�X�%|<�6��t:�ot֔/�n:��"ߣ��3�>¬��@jWl
�s5�6=��iA��Ѱ�θ:�L����X�gka�r�B��᫚�f�����^u2�r5�8O�o�s�C��ҏ�K���H�*�-�g��뙆��ñ�?L_�BJ�\N`5Џr�v���E��TZQخ���pڽ�K)�3�{��Y�<�b��������yh����Rc>;���I�w'đKrC���B��V�}��˩��L�5��f��-g^�<u���ˋ���w�t�ݧ[O�vi.�������������/��3-��H`���r��ɷ?b�+��EO��1Z4��|.�t�����P�6`-���!Ts҉�o�! `m9G�0��s�a��>s�t��w;����h]�{���	��Ҫ
Y� E@<��L����T$�B�_+�K��N�
��h=)�i���j`�>�����: �_S�����b�ڮ�g/���EȽL���A�B�7����� ��&�l���p���<
 �Gs���P�1��NlNK�]�ޗ�;d��P�mm4c#\�;q�}ϝt���W����<&������v�KP�n��ѦyObۋqM��>���p�o��P�S%Mq #���.'���{u�{�4>��Ǡʫ+4�����zo��N�0ؗ�d8M��>PQͲ�+�s,�����"u��& #��%q��:S77�������u0�X��<)�qՅq�%搛to�܈Z�I��MwV�.�r�
{Dޥ���bY�]7BZ�VA��0;���w��
�i]�|'@�3�b�"���^����d7�&q��J���5{/b@ Ŧ��eA�h�J���F5�أ���g J<�qʴ1�|������gs�r�������4�F�&^pr�S���tY}-����h���R�=Gc.1���{�1�;�ӋvJ�]��^2*@��Q;'s��O�z����q��顡�9��؜�{jU�i��8Ԯ�\2�s4ܰ	����^T�[,�t-Wl0��y]�����⎙���=��Z�j�Ek�vƋY,r�b;它5���`�b��wR"�
' X�P���
��]h��[)�}�����gS`�i��="^*������ߘvo��Q�qΜ7s0�i��i�~�(Ќ��WBng]���$����2��1�����5��A�vD��mrxi,@�!č�6l�	�s��9��R4���EG)�X;�31Y cŐ�1�z['_�:�]�
��7�!�B�(d
��Tm*��4L�NZ[�Ui���=�ߢ'��ùw����m�zi��\X�+,��*��|'����w8��<�V>mu�}^�����v#Xn�c�-��_<=7::���\Q%�!��fM8��wh����sOv�D��S��%.�2�� v��F�*��	'����j(��.6Y�������kB�9]��2x��[����je-ކ�R�E4>mWj�m5}`��BRc}՝R��n�N�����&��kc����&^ZuہoA}M����w%E�HxjBnU�5�JܦS��T�κ]�w-�S{,�sڢ� ���t{b*����A��F�CUh����{�1zv�{�9�^�|za�ӐܑVݑ��]�E���n���|�Q<e��"'�eI)W�4�P���5�ޮ���f2͖���МX2M��ͥ�k��q��+�*mU�����"#����μ2�r�����=��\dY���rS缎�-]��8]��;�_Z�ä�	ꅶD�r9�.E2��1��A*bQ��ӫ+�m��/����䩒�5DX	���"V��yq��*.�/�iOy�9�B81hl�9�>�0�/˞�9�6���C&����8�yFWbr��m�o�	�����Q�b��>	*��ܬ�F92xg�;�v�"4��7��R�Ǚ�w9z<]��j�]�Z+B�)���;�ns������8�⪡�=�ހ�:��b֤ �K\�U���զ�0���5n�p��t��g�K�mLߎ��硂n*j�1Vi7d���gܖ�u��E^���}5A[K�S��0B�>(M�Æ� �p�a���Ƕ�'��Vt ��Ch�)v��;�b���Vf4P��#�Z`�5�r�:Ɂ
�eIaJuEkV(�r��C�U������O�߂��PC+=Ko4 ��cfY�R�ϢWVU���7�Ą;8-��ݼIVX	�P��whJ����D}�=�˯����=j�����lnz�n��l�f�փB�+�g�tB��hH�4����si�Y����	dwc���"�-O7=�)��燭L[�Fw-9�2�D4��O�q-�Uf�8�[~���B���-j&GoF{G��8�6 ���;����9.ښE��w�˾�h�^�	<�K�Cv�q�B�#P���Ƥ_�u,><�Em)
�X��Y�|
�f�Rn(� vo��|]m<<��A������eߪ�9:+u�Y�'1��+���N�#�[�S
��!} �Ḡ�vՉo�fqZ*ϣ������Ƌ�S�����t�>>�v��7}��uO@�~�F3��N�<먳9���h�R�5���*�Lbo� �ɪA|[�L\,"i�Z�Q;1�>Ht�C���&�����ݵ`��VG+��|�F\BUJnx�:`�1`J�Rg���$�B{��4fU��i>q"Q:�P�M�����1�K�I��mTHXS&�|۠9��2����ʥw#��S�}W2�P���8��:���L��vq�,�(�`f",�/�������뮰�3�����$"�MCUN�*�!�J�=�nՁ�����}[�����C�8�:��r�a�s��E�5�szе���s���8�g���WY1ܺ$|���z/��%N��3���J�U�S�k��u��~�������8ad$�B:��K��������
���gXfx�c�Wq�g+�
W�SÂ��i1f��� �}��3j�fv�R�b�$�v�p�ܡ]zs��f���@��6hg��	
��nW�c�0�޳Y��5Zt�y�S�-��S3pu�90�1�Vy;� �Us�3r�PY��}Ԁݿ��,3Mn,�����W(���ϜOL`�3)�B M��2�6�^Ŵa�}0}�['A�	_G[9n�\������`T��+n�(��!�0��2�|�}�<���s�7FL_m�����<[|kf��h9>;@�r�MV�1���A�sB.��>���?/Ge����z w�R��;ۜF��͟`���ӂ����8�+�@�WK[�ʛl�S�L��gy�S۹t�lo=̹��װ�pX�j��6�D�У�,��� w9��t�$y����w�#o�Y��u�b�éc��i��aۂ���R�W�C�}&a|��31�����
�v �h�2�0�X���0ͺ�f9�d�z1�]���	�O^,�9Ll�7� �Z]юނ�u5j�vV�0=��Չ�6�m�%\��	�-c�����g�^jg�>��M�hRG�a�osge�vmu��N�����W�Wի|�Dg�y10"��}¾Z��[��K�΍%�9�6�RJd�����OB�7�) ?P�����2�����𯫓��9���/kM�Z�}84����]������0�i�H�1�v��\tn�����2�u�7�s!��*M.�5l�ַk�ح��^L�j��=D�
��FB槈S� �R�|��_�>��$WA������s��k8��E��Dk(\�x(��뜯m�CO���Ů^�׾���[�}Juf�]�%�]���wt`9�� ��9��F���e�цh���4�b��os�uoV�c����CE���c������gmtT28�gT�,����s�'�ŀn��k�݀wh�+ے֗v��KG����yҙ�;�0�M����?0��(Ry������JëzL�uk4G{�X�d�TyX��6jy�������T�dࡌ�����&�7^D��<��������d�:.%��K�xߡ�!�Bπ�
�Q���
��9V�]�SF������U�Y�E�be&��ٮ�l]2f�K�v�㽼���PB��u�\P�X�S*˜L�N�b�g�>Lq�k��!7[������j�Xnd�̅e����
^��'r�2�ݛ,k�*v��	��­���o>�t����Ol�B��i�Xj��]ٳZ�k���4�7 [��d#u �����s3�h�_O��fY��c-a��+Ŗ�]�a����%����e.�H!(� ym����]�L�%v�v;��X�~�.��ü�*J��r�#Qc��ޭ�?�ԋdn؋����n�\c12�X�8�k�:P�Ц-���^ү��vӫ��|��;@��S�vͮ|��t��պ��uGN()�q� ��:Z�r�4Q�%�;$�!c����4���u�@�3b)�r<�)I�v�T.���-�W+�ٔdg~x8��14z��� uE�ѭ�zv!9�k7�/Q˭k�#	K�d7׹�;�,7�c*CI���Zhh�J��G>h¡��V���Xi�(h���׀q]���kY|��핋���-�Q�t���1�V�>L�銰x�����˸%ڲ�,]I��y���"f���B+�P�D��{����#�;A������C"��2ݹ�F�Pu�[���	B뻧o	QB �}º�ϬWp�ܞ�e�VsZ#MKǛ˞`1 �t1�g�z� �d���Я9���$�e���eEN�y�ۓV�BB�Y�pu�F����æpYY���P�a�U��<"�h����=&�p$�5㙸�;����Lݜ��Mo�Oo�>��=�i�>�<J��u��s���l=W�ǯ'+!�wu咕2�O��V��%o]GQ.�2mlg^Ќ�q�;�y���uj@jy���'@{<�+�m;}@]v����&����T�0�f��:�Ʈ�	��__k�B���Ҏ�<�v���K�P��-ə�b�𶑲��d}�����J&P㷚 \�ʂ����W��a����[��gp�8y;.k�6(*��5��3ՉbEZ=kX �R��ݗm��[䃱������r�ŁD:MK*�'B����a+d,���t���]N�3lid�o.�Xޙ�զ��F�v⁁>�ϧ[Ycҭ��=��b)����J���<���nL���3X���=��1R�+�u�m9p��t��wO0�S4a'�+Ҵa�}�p��O�Ԗ"�`�����f`$G\˝���=#�D)��:jPe��[O/H�v;��GJ�4:mf��Ic���� 6��s$4�Ԋ��qǏ�p��;h�~w.nu�]iued�'�6�ٸJ����Pؙ�*2/��E��WOt�u�`f��'w)_ZfӦ�Ձ[����ek�<#�2�hZо�����%e�p�VЍn���Ͽ=���6JH�cd��dY4DTQ��X��TX�4PJ(�h�$شm��X�E��`ѫ$Q�(�	�4kF��b�b���1�Rh�4��#Z6-��#�ƨ*5�(�hѵmPV*M`�#Bd���TlE$V(�%�h��F�*66łƴI��Ѭh��PP^��m�S��5�ލu�c��U���V��1�p�'"g�:{y2�X.�jtc���%VQ����$N=��ވ��G��'��x)#N��%�f��A[H}�^�gY��	A��O�|��E"�=�~��y�ǟ���;�͕���t��}/��v�\d4b��x�����h=�9��D��	9��\��Ē<��I�0��gg\RTc���>zQ��1hp���>��/"eh]�M�Y?��6EզB�b��{^����K�̭y!|�ڏ���9}��
䱑��ގ�M��l��x	a��)l��<�����;�F�-�#��䈙�I�ow]�[$��U^�+
�A��Ӳ�'�J�e2�d#Ɩ�p�N�1[�+Ç Z�7X�n[�;K
�&�2�ߊI�YE���D*G}��[9��,=�Xu��x����z�H��v�T�]a,_���\U� 6 ��V�w��z^b`"`^ba��|b\=��+!���~�J�/>X�(��&�"&8�v����$�ͩM�v��JE�U�a��=��}���Utn2�K�GjŇ���{�zXw+�,������h��5l�s�Z4,E"G����5�XY}^ $�<�m�8�ئ�U(E�]8e;��St0�RاemƉ�7��Ze>zE���-i�qPՌDYV�]�av�:y�uѷ�����X#�9�RdM�_A�')�T;��ntWt\�y7'�����Օ�TL�wR�S��Y�mTb��9��OxٿnVL#ɓ�s��}OA�n�7�Bn[zr�=5�J��h8��3����iO��+��np����pL��>̯!W��5��.���>�\ίkE�C����o4\!A���ק+�����}'�'/����s�bsJԾcO{�R��a��U�����7"���Ǖ:n�3(�!��U�a�,�d8��j��s�xs�
 p@O�����;�:��t#~�!ټܺ�r�k�xȦq�*�mm��HY��r�I��@5�z�>�g���+�{��랁�N�F_�����M��3�T2�A�A�t�N�C�X�~���B�D9\-D�������Tc0؃��΢�Í��3b��̛��i�Mz��$�K@_�]>۪F�W0Y�X�5�[��C/�[�}�FHT��j\rܿ�c��n8H���_t�%y��)�-��qۯ��w���<6�M���T�in`w�R��8o(õ�?\��z�'�DDn��0�5�י=��=vP�a���j�0B�́�������vF�v���.�ע�ܬ�N����wX��o��%@�d:ƣO���wY�� U��0��
9�geؗQ$��R�.��bV�Ǘ,�Wmw^�#x��,Ԭv�Otnк*?׽�{��u��m�xdG��T����a����q7��6%���`#��N���tm^\_wgr�!gT_��{��j�]pMR�-�&/�ńKnp���h�f8c���n�&OE�9���Q���rD���Q�-�U�xL[���M��� `�DTDNo�`�&�-N�ʼZ+���DL��������s`�R�Rz|[U+咙4TX�Trv����kR��\rA8ՒV���ͮ�s����2���0��j��X�m�!o����ż�4^-�����ґ���t�
�4��U���׬�[�	��9XQ;T����9%}hP�488j�dd.t���ᵕb�sʜ:9�~sa��uv|�D5��f��
����%�_�m�/\�mp�s1p���9��Sѡ&�'3�xM��
LGW�����%ղ'/�J*�襼N�R#�	���j5�aױm4�f4���W�g��+j�=����ق�� �C�5��D4;�6���`_��0�^9���H���]ڧ�Ꜯ>�46Ɂ^���uk�<1�q͚�,�R^�}�x����3v��¡�S���8���p�[���,�E��ݏ2[8�5��{8՜kqwUÊ�w
�c��w��b�ѣ)��j��Ի�j�r��ˋ���ʎp�P��"">����ti��AI���`SF��I�'G?�X:VF�u�U��Z���C�#���4t��o[▭tg4�،z��×���Эc!�GK|�8�+�U@�W��~76���+����s����t�Rr.}�)*�m\>�8��(G��Ps����c�bպ�������z���i��r�Q���뭦H����5�㋛�;;ͱL{�.0�%����OD-|b�Sf:HF��7}<M�c�\��+��ph��j�]q�[c�=$�� 104|���+�݁?o�?lrt��3�9�`;X{�tN�,v`}��FM�AVb�=�b�̒���#pL	��W�:S67���\]���@��/�pi����E�
��rH?��*�U��]�K�xe�q�4�s�K�	�{�W��᳤-<&L8i;4m���q�]l� UA�Jc�x��ΛJ���in�vV���f��]�T��*�8,1���Cbwt-�l�	�s��w2�NŘZ2��]��v5�FPʃ�S���fDW�kN��D�c�϶�ΖM�R���7n�"��ejԸ=u��9E<�T�ϝeG�p��]��s�ӻ�xF���]��6��]���c��4��/����Ô�:�d�·]���2T3����> ��RsGtN/���5�R؅���k����Z�3]�Ń������qhW�c�;�����)�FJ�;�F�#&2oѝI��x�ɪV'~h�n!�]��i�8����T���Db�"�� Th��M��ek'�� om�L��̗;Tމ�J4���������W����ٹ�\-�K�xߡ�e��e��o[5wKp�@W�K�����[�i���PR3�Ͷ;=u��^p����B�W���P8x]Ph�|w:=W]/��̏dw��1_0���c}X|�ΧLBe��)��s�T.ʔn"�'ɇF��o5l��!����w֫$����[;9�*��s+L6|�5��MOmQ@Ա�S&6��aU ~�^���!\i�ad.&)���퀕��X�1��V��u:4�e��=����%9G���4J��d�jKB�b*����cxⶮ(�;�ASv�="�x�o�$2&��F���~z`�>s�Z=��ҙD�Ǫ%�)�_�e2�g����2[�;�gWB$��f:�NS�R[\'3���:V�fKag�uf+�����%:wl��o`�&%�ݔ���VwM#��}�H
�fM.'��3��.��nm)���w����*c}����m�R�Q�ݯ,ƋY�CC��v��óo�_UUz��wV�m٥f=nS,����;n��rG�O�_s��H�1>�μ3֪^N(K27Hi8U��+J[k��0��c (}_��Z���@m�Ts>��0l8�^��%��V\�
K���#k�o����}S�}�S%�r�ןQ`JuGN���Nfأ=	(zrޏ���h:g+��l�]o�<ϭ}���2�K�v�W9H�S� 9��n��-1{�=/+@ۑ��p2��{�h�/�JcEnN\�V��΀t�͜F��}�ˤ�m�«t}O�.ƅ�6#���:ᵟv�����$��C�诽BC7HYZ;ݞ��E��Jc�z��Q��;��@a��Գ\<��)�g����߮�}�X/�h������<����d:�p�98��'V;�:��Tc��ϸ�l���{OS*��AS�u&�6C�K5�00&�_3#"�wm��W��ael暭B�����4�)D�.�� ��xT��tX9ٟd����n�^[���w��s�Y~հ�Ik��8����;�m�����})F�`G:��s�-�P�fd[�>��t!<;$&-����\ؓ���z� r{= _���΄�B?P�%H���f�m���Ϛ����{�V�B�a��+��w����::w1��;� &��6Zl���﷖�J&N��e�IG�%2
���ژrtB��9qt�f�9xc��I�&7*I3U��,ɔ٫Ղ��!���	;Q2����ea+�,�C,P�J��uK�)�qwZ�"��0e(]ok���9�Y��6����Dt��@Gfr�G��ux{����PL���p'�a�=Ak]�y��E���0�*%�p�\��y��eQ{R:�뼧�����C���ONSh�ĳ��s��p�ك�P^?*�C�mw=��t�Ff�nEXu;S5f�f�Gg5�9qɤ}-��,���E�Ĥow3bM�a�]�q�^��#2�{Uu��1����%έ7��n1� 	��9��F�u��12�q�;���Yy�w-\�o��v�ur.^���j2�{I�y�ު�~~B�\��}~<"*��������8���c�nȮq�_=p�Aj'n˽xƹ�+����&�=��<�6;޺�r�Y���������5Gu5ėc���=��Y2c��jef�	��<�w3)���S'���wS��.���Ut�m�u;���K��-T�n��\���jL�� L6�2}����ByA[7h�)p������4�菩or��V�i(g��_^ջ�r�k�|���W�CU�tw�:`놈�̕���G1�[���_	x2�TLV>h�l�'��wowŐwg"il���VCו[�te?�k����-��*&�s7
�rb��.���ZkVL��|72X:Z�g���jV\j$o\m���Pщ�%��fp�2���!���K��Q~�[��:F]���u#U�ӫ�ڀ��@V�ж��l��Wu��BX[o�'��{]�u)���z_+���g4��>��>��y�͓#��+8w����m=�����邠=���M�
;9�b���h<Z;��Pn^�)������6���+�)P��S1��"biP��*������o
�<�b;Ե��� +}��訶Ƙ�W�Vn��]�Ԛ�Ԋ_�E�ڳ��)h���y;�[�*94�0u�n�It���	�v =ލ��(&{JU�(����K�%*�Iz��o�F��]S�z')J���Ԗ,��3�2E�X��Z\��;�Ӵ�;5���f#���Cd	>�	W��Lī\�]+�NX@ʂ�{���P����J$�">{ٔ�:[Y9eg<�T��!u	J��S��]������̝������y顴N�N%�,�
���ox�G��EO�`�}�M��!}�>sk6_s_7�5�14ۍhTf�3\�j$���u�?U��D�z���c�E�Oh�7Vߗ^#����q;~畮��c�'3f*��s]�n��J�s��a��z�#�����yS��v;��h��	=�Nh�i�K�^]9%�j3��륓���A��e�t^�\�Vֳ/�ϩqNϾ�c��S���<k�Y79Q���¢o�9l�u�Qش���d�r�S_C^�Hag���>r�ި�u�T5e�KF���{X"�	M��ɇm鈥ۨ��#.-K�z*9�OGT^(��e�}�^Fҧ�5�t`nn
���|��;Q�g�)���?U�a61Q���4���U(-͗���;\7eE�S_4�*d�EoXy;P%��j�o�y5C2l׹C/���ܗ4xX�A����3j�\㶱�H�ׯ[��:�:	S��Cz�G�ͽ�zFԽ������y9Z�Rٜ�7
"��|��g8�&���dڌ�Q�t��G�Nh��eK�u�W�J����c��ㅷ�� �y{t�GFC�C��UN��;�0tP�u�I,Fø�oi���8{5j6��Efѻ�|%&,��[�7.��}A@�I�Τ���*�U����mYG#5��ڼ�yU�?����2���W�}�0X	h1�5�o������ln�:��\4��3z�a61�fQ�JU4}P�lYJ-F��i3ef�q/��ޜ�\Ն�;�LTb�g�;@�޻;����p.X�����o��sozR[T��9f[�g��ȓ�r��Q�2�3t:͐�#sƂ���������y�up�æ�cV��v��Da�!s�U�=��Fny%�����q�rwη��va���j�x�;Ӱ�Z�.x��)�������3��M�������#Ypy��&�v|C�t&��f���{�[�x,�%>{�Z��g\���]�zN˕�����.Wջ�9�.�#���T���zS�F��0(�2�;L�I�CW��M�N��k���6���pI�ɏ*X�hvu��6G�u�åk�:�pt-��_��ں��r��|�l=�)�mU��qL�e��詍�l�U�{�5շ";s��k��b؛p�x�n#�oe�G����]8�%s�u�"�b��T��2�*��p��#�m���R�U��BP�Re����,r��������|48���K�)k�@�}i�W�K�+�6�Wc�.|0������i1���;cb"��_,�1_[�|���i���B�L��M&/O6��$��k�����2��l�cC�!��b��yy�/r��+Nb�cA���R@FJ�Q�RľΩّj�}+hh���a+9��{y�yp=�F���!�P�$���[LV��j޾�;��<f�E��p�뗕�F���уz0�&���.
��n�T���˕A��n$C���飮�>�G(R�a�{,wX�-;d�5���+6�E[�z}�<�\5K�\�8'��Fm雫+�R��dŮ;�5�/{�6Y�J%|��q���]��T�.���鬹mbFfF�|����}��mBR��/)Tݳ�(���^:_*��gQ�	�C�+N�8�����l�Y�5@�<��ಢY]���|�;;%\v�eX�i�bi\q��ܱ���j
�ě�he��o���-���ohstX�N��8���:�l��ج&�]ZO�`6�r�V�2�ł%�Y�3� �2v�W�C��z��.'�f��=���E��9�l�].�8n��;����愮�uT����wfҖhC�K�ӆ[4����]�9�B�Vq��'݀��vg˟m'���^�D�kۘ0/:�r�(�
�в���w-����l�'Ȱ���T5{J�i�Վ�������A�w�ٕq���Z�B�V��S{�C̾��ړ	]j��a���" ����A�&l������C�v��X�;��CT��:���q�Z��3���1��feHz�n�rP���r���KF�^ K$��5ڎ�9b:����h��sbk��5l0汥�3�Ib��5Vo[w�VeC��D��]G3�V�5����c��F�m�tN5t��8g��x��Ao|ie*�7�A�\����:WV9!�B#]��4�gA��ܛ�v<�S{:\��]6�4wٴ�����ݪQ�#UV�,ouվ0���WW\�'W���&�u��;2�뫮Gl,e��]I��Kv.�w�`lF�V�Q}D�ՠk��֋<��f0Hx[�Ȱ@�ѻ�(	Mˮ+~j���[=�-\���+7K�ƅ�ɵw�^��ý�"
눈��#|�W6�/i^j�n�<�l�I{Bf$6�$����E)'�\��~} @DX��d�j5E�*V�Al�ch*-�_[�5�n-�r�F�"S��4�8�s�رA�V��q\m����F,U&��m�4h��"�5��Q���n4��ɱQL��5�m*��V-A��g����Ͻt���{����]6�wO�R��g:�S'\J�k���F'[2j�}�5�r榕ۜ(�[H�]7�+��|��75�[�{�#j�i�5��s��+���s.<�NbeX���xM'�q):���o�T^>eUss��_'Y��h�2��XGk(�#��������7g�s��<������m�ۨ�僕�*:�F��pP�t9Y �=r=�3�m(J�k����+��m�S�a��7��nz5�z�x�e�U�l�JA�QR��PUB�h�oc��o��h�uI�32�s�(�Zqk��� �EOs;^ϑ��I�6�C�uy��;O�鋆x�cS��C��͆�,�y�L@)\��y����@ԒU'6�T��^�Պ�hnfUd�>�V֯��m<g)�U��ﻦ���!��z��<Х��g�޵���-���y��cj�0�Xo7��q��s��E$+�NL��U�{�����ʎM+�7�ä7��F�#4L�j��������qW��N�)��`�����՞�s=j���2�Ӻ� �0(2zWy��]��6Z4��t2��`
ឬ2y�Y}��u�Z��Pj�Y)u�w(���鏋������;������t�xG'�R.�o�Fow��N�G1r�<}׬�8:�yF���GR��y:|�%�z!7��j}�0�+լD�b^S�.���5�/��;��	���Wy��[~��-����i�w9mǋn��5M?&�Y��_����y׷�dKio?e56i�2n*'c��Hl�T�8�N��k�Z}�ok�Z�F��VzR\~HjfE?���9~Lk���C/9z/j��\k��z�eOw�֗ƶ{L���}��L��ò�
����'�TT^>hX�w��׻[4��y�R�����; {Ī}*�f�����Q791ۅE��z���;ų.Z`�N2��5o1��L,
�ޭ�SS���Dal�U���V��yjy%�?S3��ll��Q�2�����R5\mӫ�P����Ӫ�*�҇.<��,�o&�;Oee�C�������n�>�>�;�k��S��sw�YL���䋎�|��o�e��U�6ʤF\f��nt��D�"Q ��
̄:8�ӆL���o����קU`kv�]L~�:�����;�v#���ؤi*������+A�j�<n%�HugL����W-N�\�[����v?V�߇{��Ƹk/-m<�6�
<�����]��F�m����Ĝ�~��>�r��ڿ*O=k��΂�r�$]�ڻ9��yj�98�p|z���oG5����-}5�o��+}����W�H�'@����Q�j���3�t�|�1PR�QW<�z����Ҋ*g��z�W5��/V0�CO!�9��R����j:�kUs���=pųD�'�����ngr�P�J~@�+@T{��H�q<k�k�b�`^c}bJ�9��]�G��;T����sNj�q��5ؓ�j$�=���x�����=���:p���+_<o�<<�u59���s��� !���-b�]�L��
g�����"�������{go�T��k�]��4V�F<;N���u�-��C1T��+_ќ���eU<C3�N& s��v��tЫ�Ϋޒ4���F� b��/��i1�a뻺o��)Y F�g�^�Ɲfsf��݊5���j��AJ�o��QYx+"͠Bo�����ַH=�/zS���R�j�ԩE��o.>v�dK�Niul᭚Yu�������Z>{��҅[�K7$[���w���c0:�Z4o`Oxv	��ۗ׽u���;��dΤ��ӽ��^���KG���c�`�ԻŶq�\q�F"1EtwF������yފ]�agW��v���Vs�Q��J�W7��г\�ONʆ�k����Cx|�|<�j#���]�x�\�]�'�+H�d��FԹw�]�R�#ÎÎߛO_=kro��7U�A�v�����9���|�JK���~v��L�s�����HPk��^,Avz��5h$�������޺RO|�W+}X}�'�J�VOO(|�r���Ks��mE�1�r���,�\iMe�Y-�u�l2�:�4����]�<H��ֱ���9���)T@�-Tb��1�����"9Py�K�X����Oxg.iz[�f%�(�+Э
�nz2 ����n��e����=������;Ux,X�=e���7!� ��ؠy{We>z��y�|t/J#��秲�S�oEb���f�|��4tɭR��c���;W��EN�N�-'����Ud�N���3qu��s_�Y0q�Fw�e^�s-xH���q�qO�����:����a��c�nn���%wD띭���i	ܒьl��@W?����ٍն��0ں��)v_��p�%O�Yg�ʽQGd��<P�T�����s�skNe�=
I7昚+���T*���f�9�7�J��]��O[�_`��\�,�Ax;mU�ps���b~����s]���YS�;O�-���js�+'���*v��}�K൉np�qx��*�n]c��1Ɲ�,���S�j�覛��r2;�&����5�4�q�㊃˘0���vޟR��w#/�l�b�O��ީ��Ո��ў��s��Vm�H�뵒��\��C-�0�3���+�E9vI,��2�}3��ĎWt����+J���L)y�U�j4�1F;����I�^���P.o�{s']���zs���<v��U��,�r���c��}c���yaJh�2=�t괫�aǬ6�ӛ�wu��Wm�O�i ·^�XzYS�DEf �7<����yKu�ٜ�ݚ�vY/_,Jc/'j2Be'
p��ct�,��A�oh����i�(������S�:��٣BD�T����1�m�<�����h�cw�S���ۛR-Xߴo.�n�{x�B��~����q�p�IX��;��#j���sQ�:��n�uUA�=7�<�[ֵ���bY׸���AlmC�d�jewh�C���m��x��� K''�cR���V����O�)(�UE�ڞ*�6n���çdA~�AZ�vN��t�K���ya�W
s��v��%t��c0���V��;�;�6��uXg��9�{�a�A3��}��mW=J���9�MƲ���x'��I[��ۑ'�e.��G5]y��}�����tV�'|ak�VZ��o/Y�v-ok�P�3sm�Q�J��$]b�sas�5��gs[��o�=>Z���s������`v���M,��`�a׻U�p�g{�%���Q5��x�z�CU��zȊ8�ݿ�����WR�gll;�-��8h��d�;��R�˻BD:�ē������w�yV]��v~�|s7�(sZ/Q�a��ܶ�N�epz��0=��晶�uv��Œ83{0r�>�i�=sc �����3�3vwZ!x��im0�e˚N{%F���V��$�{��Sy']�.�6��r�1ٴt��Z�����wWZ���
�Q������[�ܶ����Ks̷���z����w ;�zFJ�n�g$���Ǉb��=�㡹��M�0�=0/j;H�S;^��!���~��>T~�8�w��)_a*��:�8�m���Z�M�v��ְ���V꼇!��� [�p`cCg��W-���I��=k���/�
1ە}�IP	�c+k9'���y���`%�q���Cz־��E��'ƹ�� �J�7]��KCۺᚅ�R�w�J�X�w;�c����7�r�rr���[.t���]-$q~�Zy�&�y�X�";_�w?�G��Wm�<�g9M�nz�fl������r���@v�B�>T��C;�6�=�e6x����>���l��p�ͫյ�ʺQ��DgSk�P���p<.xw�H��GYc�]CNmX�V���a�r�F2�I$�3�t�*�ICtɾ�Gnn��w>���ݫt�����4�R��;��m�k�5������VFp�wC��Lv�Y��\��ok[΅�]�}u~朮��<hgI���rU��9����]]�{��*J�N�O0巴wV���|����_�q;�Մ���Ň��mb�n�[��_Wl�/�ۢ��������Ӟ�^�>E�-p�i���U�+,���dC�;�C�Jv��Fr�K����vN�N���5�P#3��}O��׏nv���J��������c2�����T�tw��UjU�|���K��.�vCJm����WMw{��dg9&U���*26�)�7Z��;+\	�J�8��ZԸvޚ]�}:�H���}\{R�2�S��Nje�;�R�i�V5Ҽ-͕�M�>��H:�U���2�p��aA�*�e?U9���ą~V���\c������k�]F��H��b��$�!W�N��
~�IP~��I*��:{(�p�4+��.��Ta�8�Vc��7�X[���*h��ɱ����pS��zb��␛�A�ǡ�����R�)Щ^	c(Yh�ޭ�k,b�]v�|��d���碳�O`��惔�ĤU�����О�wU�J6����#
'x�v<�s{g#yZ��g�)T@����*I���#��yۊ����SXx��f��i��N·ې�ͨ��2�"�}�0X%-�s\� ��TO(-Gs+�sj�ĳwYM+�oZ�gpSl�,�"T	Kg{
����l���Yڿe��i����C|�LTb�@q@OH�6�s��A��n�ED��M�Vmv���v�M�O4�_@n1�X��9�qKp<mb���DW��E�m}c�j�o�+�S�f7V�.z�6��6���s�9�R�]�������K��n�?!yS�2���m�y�쵯�;���;]�]J���e�V9f����������5�q��=�%u�b�eO%ʖ�����mv�%�n���0��sq�k�Ό9Q̃z�2A�P��r�+gN��Wú(��r�MNv���|�ܨw������k��tz�ީ�cPK��/,5�X�3���kZ�d�\]O!��'hQ��sL#�Ln�������z��aW{�R�/o�΂�`ݗ-��ap:7QT�4�Օ/��6c�t ��J�dB)�v��|j�3p k6�/��Z�+�gJ�G�OFPce���fHK:����u79C���s<���1K�AHˡte��ʢ�S��YFq��)]�����6��҄���������D�}��	������U�����y��\�)B�I�+0ܻ����*�<P�������qsʷ��{�oO����#Sz��#�t�oz��N6�����1��p��r� �;�}�D�������3�����Em�.�Uç�a-k���9�]%sr��:Y=������}%�D�[�qy,�z���-���7�*-���Wޤ��i��E�{��B�,�Ծs-ب<�kis�X��ʎM(o�Q)쌙ћ��z�:md�ݫ"��(�����V����7��D>C3ؕ���mvrܡ��9�2�c0���r��HN猭��-�/A�ƅ>Y�j��b�땴���w<B��w[Փ7u���Æcu'�S�>{���cD]�9p��p�,f�7�(�N�-� p*��Z�\x�,�>�f�lܩQ�Y�=���Sn'[n�t$v�>���b�T,��ޚ�Ԩ����1�u�EU�ʝv�,�T��j�9��K���d�z{(��3\���X�cz\Y5v]�grru��Yīܮ��$*$әd.�4�:�d�r,�V�FC[7�Q�t�Dno:� �eY�����Ѵk���{BV�}�"W��K;M�y�T�u�l\�r����8>cE�T ���zY|�
�셊�PMnХ�z��U�)$��u�z��\�7��]���z�˶]An�gj�Jm���-�a����2�'��=V����в@ I�z3n^�a���mR�b���Ù�{k6b�m1� +;9�c{EKs[�5B���q��Ec*�2^�d�����um�%tKr���*s�L��ܐ���	}Zq��2Wa@Nnb�8��-
lޱk��� f��������۷th�遃�wJ���μ��[ŢSi9�:��뢳1�ge�g+]q4�Tk�������Gq�D"��aS.�h%�7��Nӊ�uݢ��,���"mg>t�Z�}�����T�y�O\����>�ɷ��p��u3�Ih����)<N$*3���V����īc'�W�Z�q押�ǌt3�Y�j��h��s�M�M��V2 �ݜ��;�c�B]"�f���U�8Jg��r�R�V�;�϶�X���wo0> �Ž:�Q�
��+�1&� a��$[��:U������Ҳ���,�U2h't3�6�ϒ[3�v3��U�툫�<Ek��n�,k[�Ze���dwP]ᕱݚ�Q�Y�F4Eu����^%��nI��75�7%<��T!�s�p�&2�+HV��\6�!�N��C�
�)B�un�q�Nl՝o
�G����	��/���g2�œ�a�i�w����ɳJJ���\k�:��%o�0�v3H��t%+��˥Òb�Z<���)r��O]e����u,-��[(֤�n9��8��evmt���M���]A�a�Sr����1짐�����}�4�;�Ý�F�������0��\��Z�D�"+(�F�rք#��U��V_;�����:;`�Ă�Y���ܻ4���˫q��m6�>Cug:���#��ޜ�w:�p
yi�V㩀��蝖�H�.���E73�'�w0'r�lV���)a�}���
��A�$6�(D��;����5�m��=MRBgF�Iu��NU�����7}���x#�,�|;2����1�v�AW;�]j��l�S��U����·�v���a����A���wb� �������s�ڵX$9dL�µ�G��Z����ܷO��GS�-h�i!�WL`��Vn�{�
[�����V�[�z(���O�����O��������2^���z�he�b�nl��u@P�U����n8�QV5�.+�1V6�VlZ�q�#n5��\�,j6�Y*Tj�F��8ѴZ-�A�q�Q��."����ch��g���PRDXэc���\pNr�F�V7�.��q�0��R�)�ԅ��E�Zuezue�·�7WHz��e$-TeYR_m��p>n� �W�\dڅ��w�jUv�}�rζ�J���&�Y�*�5�5�S�{n%��b�h1}Gq�Z(3*ߡ�7F7V�j�E'|V�upZ��o.��7熅��;8��}[�WgL���nNv�'�ߨ�>>�OJ��k�ی5����9X�N4N�~��O|���=�i{j���^r���QX��)���|����1!OV�b��b��/J��<��K�tk '=�:�Ζ����x����L5����,���!��BοC�[�=�W�r��n��'t�Yn'[�����C-���,�x�qjghs�H�tu�1TTN��w����v�m*T�'�Z�\il[��M�r�t��=����e<��0���S�VmeK�=AoҕM�F�kF8[p�z`�br�sSq��j�ݺ�h�.���P;��a��v��ؼ}Հog{o8^rodi]*��a}�²ob޻7ҵv����!Xܤ�M��N���n	d; ��K�%���jK�|s�Vi��u����ގ���k{xd��_���C-��i7�����!N��/�	uB8�vw�6k����H�Κ��F���PS�.
(%���Y��TB��E�� �7���s���G)�֤�Le9FQ�K 0JZ+J��s+�����0�8����);Ƽ��{��y홄B�)d����������MvT�,�:{�+�9M�h;a�Q����Cf w�ˮ/H�"�خVNGb<��gU�մ}�oй˸o�j9�%����vE�n-��hq���E���dE�q(ׂ��m��Z��lBN��c�-�&��g.�qPaJӺ�=��Qʞ��|��)��o?ws��-��=[1��<ڧ��;
��A��UY�c��k�7�]��Ok������n�l%�-ď6�E�����U,�֮��Pʏ^sF�����TM�3��y�	C� 7�Νg��ҜpQG�3�T���z����G.�g9̕lo�*��P�4稵��5k�s�o=��;5O)�+��͉h�6�U�&+f����8����F�=�@jZ3�3��6�C���u��;c��ג=W���
�Z���{u��u�g��g!�ٜwiT]	�k��y�-�9(t�oº����/KY��\��]w��\�ި�̈́����P��㎼������ziv���;cn�,�P���&�#�:�×���;d�ݥ	\v�`nJ��y6�����3��y��q�+2{���|�uO �G���Ƶ?���17�7���͛��on{XQִ����� �\��s�ꀠz_+��$�ݽ��X�{iP[Y�(Ʒ0���z}���p�T�T��y��$�bu%'_R��w��Y/j��Lu�U=�r��e��79����g��Q��@sA�1�]cqY�Uډy��y��W�{��M#k<���o�1HJ���'U�GCYF�&dT���W)���=�	���2��5a� ���<{>���\^ ���SZxۑ�����W�l�o'O�u�MG4ø]u��͑=�4V$UaثqTG2&���D��셹�+9��[p����)ösaj�Õ�m|g8��^��6��,�Z�0ovb����ǁM݋�r8�m�{}l`��L��RD�9��M��*Y�t���PG�`7�g�T��{��;8%S6��o�dbtP��E�굙!�yd�llI� �\�d��
j!7�ʯ�^<�L[C/��9������^�j�xJ�NL�{�5C	;�\:��rᬻՀߵOW����V*R�����r�y(��nt��wm3�T��q�dk�ܼ�s ީ̌��nΞ���V���.�H}�������Q^���U��yޮ)��ӳ xP��j��|+��g2�#^���F��>�Q��0a_7%�{*��3]�����*�v����(܉qퟏ�A�biX{��m�7�{��ч�7�-˞����ָ��dk��[�����s�S��\m�
���ݹ�y���k��b����i�z�竔��P"_*&l��H�s��<guT�Ҧs�c�p�ㅜ�R��>�>��ڳP_Y�f�u`�����9��q6���v��|vֻ=���/����;�	�e�3M8u7,���%A,d�ƯlU�.��e�!��
[u��׃W9Q��fp�ys�n�(��xYox�[��b��w�i���X)�-[h��Y�VͩC*Ӿ_�ҍ�|�}�zT�z���i��u1��%W,r����Ɔ�ctFO��迭���V�k2 -�Z�Ci/��{���R��	��@���6&�a��e�)��j`h0y���K��Z��3�Jj%V���Ċ�|�q��7%].\7�q����K�; -u}k���sd���_qXʚW�Y�CdU���m�w�n1�7�O!�
t:�ܙ'�K"��r���Ue�b6����<fWV�9���k�g]|���ϱ؍�5��}Ne�<��t9�oe����[~�x�$t�Q;p�^�.��C��
�����#������Y�ֶt�pv�1����L-��wnQ��G��A����ʢs��I�v��^>eU<c'^(��r!�ix�gj���6w����,�F���ۣ�}C�ΔV���z��53�k��[7y/Ʊt�yڒ���Ӷ2��(q�q�W%n�u��x���U��r/d�0�e�b�̔�^S�Ug��t�;���y�q���ko/��Ε�Vk�8qk5��
���ϱ.��\h�����_k��(�Jz�z�Kkzj���k�{�XnH��d�ʓ^�tZ�V�MR���z��g1��Ju���힮[�ͥ�QՅ�\��tިwۦꃤeũ��tꃃ�z|Og^�N6�����m@v��>�ܗ��m�i�@;^�#�yf����)+r�e�v������r�+�*�J��7�5�Xq��m=�=չ�(�ԮYVY۾�oӁAN�~.�;�a����I��u̝ɺ�9����X�F�ˎ��2��J�1�>�*|�Q��̮s��U����*vcw��W�n��U���rW��ַ��2���%u�	�ܬ�`9�0,A��U�CSg�&^k�I}޷��
m�W�٘D.�)F���#H�����K�*Z�[�'OxeG.sP�����q0�	���'R�-�r*�,tX���±t�ī��1���0龩�i���k�o������wt�9�����Iݸ�5��0�-=����ubI��,p�rp,U��[\a�z�`X��Hə
$vc3����v���+4����31�NQ�φjA�E�B�<�|�I�����l�ؚ�u\{����kf,���
+*������K!w��M�\�7��e��-�n�][x��EdkٝҊe�k�� ��u��y����kg����Y綔��S9������V]�+uz�<vS�|���~�P��c3��W��n1NA瓘�*�T	X0E�M̮������P[k�K����v6#���T3ՙ�4o���.�{ǳ�m�](}uBn�g(3ۺ�O��M�1Q�̪���;��5�׶�sw�pe����7�E���52�}�Ӻ%�Wv��r����Sٛ���[:P7+�4�Y>�u��߶����n�_��$g]����*����"�j���|�0���Kkt�Jgr�U���&m=�6l�j�=�j��]�&%h���7��t-���ۃ{�(w ; (�m�#aġ��R24�m���Xp]��5i�c��8e¤��s��}%A��LA�hBjd⨩w�����q��V��7�e�ۍ�inK/!*��S7ʃ���݃��
���]�@�c�-��3T�I���2^�J�򳻽�RJ�]=]��̲��(��T=��׷&,z�؝<����-�{{gq�vM$_)
�K�*�ǚqes����ߎe����w66���I���y����I�p{�q�n�_�i��H9�y녽�Bi`�Np��6��:cb�;����-���|���`?{S�k��D���r�7��v�Q�1Yf�ltm��{�&��X4m�j�:ek���l�'p�K�o��#�i�o/(#QU�j�]7�S�@�BdO)��H[r̭�<�ŕ��0��;�:7j���O24�=J��<ۍv�Uk�'��kj_T���ŋ�J����.~u䣛��o���X�9�Z��E�_5�Z��}�tĕǶ�ë:ᥖfM�	N����\V��1��ǎ�gʩ�n9��s��9�ݧռp��[Z�m���?|9R^o�2�TLe�v�y���rs�8T��3�޽�ЍV�2��QO�̢�,��˚P��qA��w��r6W=��"�b�6%x��5�z�%��c��'�Ykz�7��>��^�q�Wt��=�7��l�n��>;������ &�=�ѧR4�]{�qx�[�:^�α�rc]�T�\U"��C��cZ�d-��ji.���(�Y�gmur�f��Գ�#��=�(70�r��"	���T������Zq��H��R=�x����㔹>�_/!��ɆRt����~1�5^>��O+�>��[[�n�X��{=�,�$$�D4�ж�@���������}q-=����
1���h��"���CM%C7�#aߡۺ�Ԟ�p��c����J�,�T�/�h1J������Z��p��ӗؖ5�\g[�0����U��2Q-�6:�ܚ��s��Il�F�k3ҷ�k�>�o��ӷ������:���>NK��6��(�1�%04{7���|���9�u�0sU]����!�$v9�r�K*i��NٔY���᠕�k�v����TlLr�vl���2��)�|�w\e*�ĭ��{Ά�x�a����f8���T鷶��B��j��'5~MƻFf5��� ��X��Gn��IS�*�e�twV�F�ē�X�S>귾����O/�{W���7)�D���d�
˼uyZ:�Ƕ��Kz)j��������w;s�\3k�����
ҫ��kr@���3�[{U�j��=C*��K�WX��ޢ��,ڗ݅�<6�2f���L��Ǻ�{���zgaH���N�A$�ngu�x;�)r���/ny-���O���,�*z|��5Q��j�6��]i�׵;>�qM�������>{W��j��|�mI]ZmRY��&��<�k�=������T�>Ѧ�Z[C�zr�5�4��j��rV�h�UXK�֑���;�Wj�k��5�,����}�nG�V��F���ڴ�T*q]Дk�e�|���e�>wۥ�;c2"�Ϋ�s.�U�PN�����)p��7+�����F47%�g�o�SOH;@��E��GulN�U�R`o�Q�u�j�{rUY�M��a�8Z���Ә���˦oP�����3<��j��F�UVwv}�ÿ;{Vy�z���WvB�]t������͸+�-RWr�����['G5�jlz7^+-�����Z|��ϢQ}�	��nK$%Wy*�r<������i�'E<�e��Nn�Z{|`�1�T�/��T����++i*D�d��S�ڎ�e�9��w!GEn}�whF����oǪș%�{@���s�F>�2<��'͘rpqҺe�;������%s��<�7��Ҷ�3gd�X�qܑQ�è�@#"qT�u`M�}�����)��Yt9qIN��nu`Wp�97�(�L��әT���y32۬齹&<c	|�-��U��6��|;s�ƑLn7���s
���ͽ�I��
҇gh�Q'B����5֬��=%oL�� �\�+hd�T�1�i@[�έ�cf��v����J��z@멨��ڲ�h�-���0
hs��
	s̖��Ak�_zt������� 5���*ɘ�����`�ZƗd���^���[tɰ�R�s���U��+���׶�d��'AB�a(�A]�A��i��u
-7�j���l�pn����d�[�m�v�[m^�u}������r�dx�Lщ�EX�Xj�I��'y�����vñ& ]F3(R=�A:�9�l�@��uoV�����mM%��rM����6���h.�ʝ�7:X�
�T	r[b[
�5{��Q(ks;��r��u�{y���u��$�u�]*�=�Q�� Zfl�ΰ�{��׋7��ֶ`�����]e����<��12�"��6���N����jLV*��8��z1u��H���Ay��S@ټXN�fry����6+�6�%հ���L�������QY.Hr�`�ޥ;$7o��ܱ�sk�P���IP$+b�:t	:����[�2�h8!��i^tk��v��w,��|-�^�+��Ӡ��q:�]X��cj�f�t�sا.�GXcX���Yf�kw�{9�j�_�w�G�U�h�v�@{/�8�ԧJ�:��N6,>�B�����ӓ��[6։�V�����H����d��IZ�h�d�w�
a���A}hjTI��V�|���ɎQk��;ج�ڬx�y\��K(0���Z}iV�[��r����� �i�i�������;�O�j<�=z�^���J�e�"�աe\ƥ�vgc/��7��KϠ<��]��P�f�yη�:��!}Hhi���
���皉�Y��{+���J8;bƐ�`�bl��V�h'V����]\[+�Ol�u���;wWU�"�Y��wP\��-��U*���ѝo��S����pR�c���v4Χ���p
[զ�M�d��A}�Ő��.����`Ϋ��j���s0.�G����i���d%Ϻ�J�� .�6�t�k���o4\�&�Z��9�fΙDc��"�n��55�S�7j��_M��hi:���@���B��C4r�n��n(9't�� a ��(Rܑ�o���c�v�wi�F�'�e4��F�bl-ch>�f)���2%�W4�%Ю�5d�Y�z�����Ͽ=}���+�4b�Qb�F�5����q�neq�h#�+����WKq����lF���8�n��HF�qC��.s��6)&1	�Ǝ6�6s��\k��h�1	(Ɛ��8��`65a�2P���pEAI�q�PR(���8��r�}��@_��� �P�L�mD���������7�iS���]�G�i����n}�W'����v�vn�����m�+"���Zz�~�ozr�H�u���7��E��*��4�j훎�=�E�$Y��٨�Kw>�D=᜹�|�����q0�+7
[@L�#�8�W�]�XGm��i��F7���.���4�͸�q�f�ez���^�O=�HW��mۭ�l������]x�N����̪�ߦo=�����U�T�ݪ~B���Y綔��%�Sy�I�pLq�h�x�};���Uc�gR�\:��fvᚨ�A�gZ�3���ۇ�s��]ZQ$�N�Hu������2�_=]z�g�3�7Q�fQw\}�t���Cٻ���8lQXx������>fRnqޮ0����v���J�u�-���C�X^�{��^u4gu�nn9sra�z}
�w_U�'(��{�@��hȳa8�S�~ԍW�.j6�%�v�Z��P䪊��7��@�f22���y��$�nf�t�E�y�X�t�oͫ{]�''I�4���v����Ti]�*��t���g�+I>rm�>6�}�\ܾz�mƪ��1�Z���c�q�D�R}�\�P�uz�����l�4�f�r����!���ev�"�^����G���x֧��u�^�a����xFK���|]�r;	�m���w�P��O�T�FԤ�� ��&u]eoO�.��ܜ+�N���t7�{/�_V�ܠP���Q�c��H�}Dȴ�.����9Ȫ�p��Xo��/�<��ߋs����
�� �#nLr��ȫh*�[��%o
�-��w��hO����Le����&c5�4d����u�ubz������pyt�u.{�uxeG.j�|����NwUL�Uͣ����q����3ŝ��"ܕ�M���Mo�����F5y�oZ�C+�N%��|���I�S�+L�^s�9��To�T9=��]���{6�{9�j��c�WۍjMdk�5�z
�7�M����?*���A�V��7��0���Z�k�V]�[�o:�y�n�4	����Bɗ�	�^�����9�"�.�ՙ�Vs<�t�4f�c��yu�]4h�9�Qe�d3x�E��߷��2��Ȟ!��+5aXCP��S+Hd���,ƀ�/�U�v�����f	�kӜ�fT�m�f�vI���WJjD�����uc�*�OӘ�(��swS�;i�B�y���:����*N�G=/�Z;ă�`'әa���tk s���+�|����z���tj��Khq.��Q�3h�*�#.#��XF��Q��M(|bqEx��4}1�����WIS��Əu��lR��]ۥf��2�-K��F�j�u[J8��AJ�ݾ}H�����c�͕�n2�?{g��Еo]�����.���Ft�:͡�sYt6�*P�Z�l�K���m��oD��@n�U�љ�Y�IC��P�=E��8�_eJo)Pu�N��\5���m��Z`�Mz�c�,}�h_U��;����[Xܾ�r�--k�5�u�;5�6,�K!Cuxn�c�P���D��V�k0-ꅯ��i��*���=Y�VSٽIv`v��r��!O��%#@�qK��� i�N�՜��h�x:�k�8k0H*E��n��e^����t�ޣs��Xg�0���Z2-��������*��&F3Oa�\�M�<It�+lCUu��#ִU�e:䫄9�s
6��=��ܖ���
t�Ġ��|`=Q������u�^n���ȧ���|��
�y��E��*	Z�#"0�j�[��:n�֪�K�Ο!�s���p�hTb�O!��K�A��l��qZ,��3:�(��=�ms�[WW��\Bn5�u�с��/��dc�R��.���xvOv��]x�N��p��Q:.X�{"�\VB6��:V7:E�s��P�U/2����M^վE㬗T�@;�I�[�p�p��u��a��A�S�c�z'1�2wX5:d�@⦩=S�y��T��7�5Y��kŐo��\j_+�Q�hS�r/ bsfgt���Wc龮JU�v�W�K���Q�3r�c�)sn2�a���R�~�P���~���s��o�C��,��B��h�f!�X�4�Bg��߄Ui��m@W]��ᲚZ駻�/f$�>WY��ؘ�M���9��G_7�	3�`��U'���l��ܡ��t���2];C&�����cj&�(�#�ݐ�Z^f<�йn��ǻ�5���-��Ԯ����8c|2�+S�N���U���P��ƺE6�;�nAFqWRW.B�O��Y�2o_E���������^�u3�U�Z��M���k0r����^��r��7���RH�ݢ�s��0;�����E�C�����Y���{jxy�]У��ɯz'�Oj��r�R�

{��T�Z+O5��w�J1
��M��+3�'=�C�!����{tT[c)�(q�%0�e�ViM�9C�\��&�y��7��-�ɥl޷��
�m�S�P�{xm���{aUŐ�[2*\���u>����=���&�;�w���-�>ǳ\Y�i����*q�G+�4����l�ym.a�7�<�P�Ȭ��ڹ�IMn�T�J����Ț�s�V�+��Z{Gum.�@c�ǔ"�9���m��y.7\)���yU��c����.����&c���p�@<�@K��~�\ޘZ��fv٪���=.<��ZPҧ֩����9���X�{F���ǈt9#!)w���:Lv	���bdM���5��a<;���3��|�w2o�Վ��b�{�`�S��$����y�̫P�.��z�]��;��"䨺������a�%��Vv�"/�o�8�p�;N�*uٺ]X��嵁>��\bN�k�%���Wb�~��捺ڑ~v}������k��R��T֩�<��>fRns��q�{�����Wd�9%{�A�f��l�TO<љF���T���X�͍�͋�M鼌R�HVV�\˷���D_��_��JsQ��+�\F�ц[0�)��k��y$�-���O3@���λX7ʁ�xז!�v�fz��A��C�w��oB����1�m���=�gB�� �5��f�M[G���=��t]G��W'��8kq�·��
ү����
�̬rv��Z�֕U߯e�M���U����_2�q�͸-�[��C0����$wG
fu��<���#����׼3o���No[xf�_������jf�S�@�g�1}=�݊�<��O*�ܝ���{��[a��۴^��%Հ�]�H+uy:Ns�[�v`�ŵƅHB;�o%l;��u��ȍs�.�٧)L�u���}m�N�,���l\ ��s��.�.��U�9^7��g瓵r(��_7+N�T�5��FtW:�t�9�����e+҇nXOR=�2U��l+B��OЩ�(�|:b~ͪ���s�lQ鳇,[hL���q&6C��5�I�a�ƅFB��Ɉ��N�sח�����'�����x��u���:���k(e޼]"o�b��bg0���~�d�crS|��ۈ�'|�å�SF�Ŋ����v����tq��M{�N߫�\Er��������n9��w;V`�P���,Q�yQi���F!�Pw��0ie@�c;Tv[�je���U���ZrB�;յ�bGb �z��є哴!ʾsp�ζT�$ia��}�~���ޙ�u0g;�t���ۅ�?^��A�U1 �VS�a	1���c�qj��b*N��am��F�����벾u�=�H��iD�=��n2��UӅ�� 6�t�U����M�P�=�[1�;'x��ԝv%�W�s�-l��)�r�^k���jkHT��L"*��-�*�go���ϑY���[�Ec�K�uTȕ`�xy��4F��w&3��b��bz1,�Q��uL�ԝ� �ޑS)���b�lA�M2��4�]�ok��0wJNq
��y%nM.�б`�C�mKw=A)S9�ޟk���Yp�-�3�R�o�4�m'i���9�s45%ki�C��_C��k���b{[���Ex��=��ާ̘�����(t���Hih��_|���9�"�N�T�o�w����1���{�ۋ�PF���}��d�a ��b��]�����r�s�?fLk�9v��c5Č�s�a���P>��^�zo�Y$��2�H����'Zg�}s쇖_D���8�X�\��B�����/ĳ��c�U���Q#ǎ����㇈�LR�`{��x&.l-�X���_C^���{��\w:2hsLF���N��=%ߕVUS�hV���8;�LwAV`�͋�/Ʒem]�c!�]Ž�T����}:B�˸��5�[��|�4X����Tqd�5�A�]7���q��>��j�(��Uߊ��R�7ݹ91f=3���tY����Β��\NL�d��=:��'�*W��	���+�#�G)j�/����a:1ޭ}��t:7��u�eм\�\XTqv���`Bo��P�mgov�V�v3�����*
|v%�R=N^��S<�NNӧB����Jy�W���J�������1�-wk}|�"7��`^c�u�%�(��<�/��-��Ɩs����ꑔ2�"u�F��.��).�%��{AüT��Uv��y���x�t�@�W��%��u�n�,U�k�6Nd��]�~4v�]\:�;�S�>�3ඥQ��{������.�9�.-�l펭��}7�3����*{�~�bл��E�r� 1��(:iqCjeɭ���]�j;!�=|��i���%x=/0��޻+ޏMp�eV�9�)��ĝ��/��@mL�Z���z��sqb���Q@�"S��W�z�+#܎�5P����f�����=Qa@��Q[R�K�Q>=�Ɨ�N�����|�_+�ע�<���9�=����j�n��p��(J|[����3(<�5�|{����W}�H���������nL[+��(<d�N*�s��g�e���v��T��W<��"��8��ʣn��c���˂��-���eF�/Q����oH�9��Q��	���T�����:�!�}j�������P�S�@s~�͂��=���^C�!��MԽ��w�;�b�"�sQ&�KA��7�O8�����a��䡞��RkY{�E��ohմ��,��%�o;����ŹJ��V6�s h��qE���i���?h��U��ʴ(�GSb#Oq�ů��kq�6�V��<�����,�g_p8�B�������r'����p�Ȑl�*�ٜ�7�qz���wC+<��}����f_���WkțE�
���rD)d�E���r�zka����T���*Gt��%m��oz�z�aO����4�1[���^ڱ�ɐv��P�i����"s�^�[�u��]����Z^��н���i���s�� s[˨��l���t5%d����n7����6;/�!��1˟D���N�<�5{^����[�g�������H�����.�y�Go*������p�/����T�}>'qK�ǂuO��w�\�����D�[��������:c�ٹS��,��b�����U��5k�V/_�	�_�=}��"�n�VV�ܪ{���n��AVT�5G�{EY��D�rkk�#��]T���$m�)3-�ʟ9��a�~]�,���+և����UI�QW�=0�����Y7d����yab��N�F�U�r��5��t;M�\i���d��,g�XC��q�4z|$�B�u��V��J�\�)p�//^�oZ���q�z~D.f����g]c7
)S��X ]r#�4ӭ{�s�����2s���V]Hz9�jbb~k:o�P���2��V�	y�J�s�B�j��ʎuHi'�MX�����<1����Փ�43RF�5��Z�N��<�ݬ�4���1�\�{�oRЋ��J�Xʸ�!�6Q�y�xdA�w�R�/l���}�HT��$���<s��H�,!�����9�7�,.P��nh�rΨ"����gxuf�^��\S��X���*����\��h��ml�YWc�u[��߃�O���)�� �c!��̙dܻ�n���ε�v]���pܫd��WO�R�[����WY[�u�:�(��2L�96Ř�jPꏲlů��Щ�����5�,ni�D�����Yy$�{��}�.����@��r�M�o��Wug��)�|V��qM�ܺ����l�\䌚�Τ#�ے�C��2w#뱍.����j*����`TvY��A�W��r��롤��T.�R
��O!ܧ#8��PRl�ƷV�3>˾���	�HKS#R[DFa��Qˢ�n�����r]�Op�ST�J�ym�uh�tyna�� �Ѝ��`�#�k�L̳����j��s���V��
Ggr�C��U�� ���O~{7[� }ꉫT%N��mK���v�uh���5T�䤥����N�,��[(:��� �Sq����3�[�G0�m]臲�u����f��������:��K\c�Kts,�c/Z�Ә��rzi�*v���;k#Ghќ�u_�����;��O��yD�X�­+(�hPp#�b�|��[ e��M��#U�mєM���׼z��<�������[he��N��>��Տ����1�����<[JC+�8�����r��*�P���y��^V�}XGT��z�oq�7���TlH�[9-�的�M���4v���y[	A7��۔(�1w{]jk&�ڤ�9񨮹����b�9�7���.�Lfw�����F��4#�}D=�
��Wm�9�Xã9ཻ�	h֨u����t�ś�G��B��kka�c.\��@u��lA���wo�*�ypͷ���h���V�WHJ��,�#c��Z�}��4�nK�F�ϝ�sR�n�ݼE�u��3�}.�wZ���v����j�8���E�t�4p-�/%���]�\�@g7���G8�H����f��X�^.BSԍ�U��
OjUΥ���X�B�oR��fu·v�=m�fLJ�wGI�P�[���ze#�vw�W1�Y�Kug�*�dǘ81��ʼ��9<��ŀ�Wt�.��	����ژgq�!�*�U��ޫ�e��`�@.�-N�u�I�w�&�W�fRk�;�Ak��ξ�è��8���j��og}�}��� 
� � ���n86�.Wrf�1Q�%qh�ɰRF..*(dq�$2cH�j���F(�Ab�qrh�9n49ˋ�pɉ1� �(��+\k�����1D�S��&
.8���3Ti �1�� ���5����&��Ą#)	d&�,I�Nr�4�!�d6D$PFIL�c�9�r�����#Lh�$h0L�9\"Bd�HƔh`d�����w���wլ���7�R��p�{�o6.���U��Am�L�����Z9\�[��͊v�s�:�Я�j}����Fj�V��wU�XחS�z�Q-:��<V�d3����f�p(s��8��m���x�� s��&�Zg�C#}S�zZ�Inv�t��l����q���sq����>�g�T�E�#��]C}$q>F��z�C%����:�%���ŏVh�����͞�v��'З�-5���G��wgд��^s�vOx�0�޲0"��Jt1f)>���t���g=,�p��٨�]AO�䶾��x�Ǧ$��Q��KG�5��T�Au�o��{�;ll��8� 7��ןK���r�#B��R`�^'"AK��-\B�7b�b�VN�{����M��x��C���o�d�v'M|ۘ�v����#?yҜb�u]�T�}�ٿX�+�W�l���OE|2�Ӌ�]���(u��W��;X�Q��L󫢡8E��E��kշVj�_xM����i:(�qj�Ԧ�E>��v�ݞ�W�A�y����<�J'ٻGpDQ�(0z���\1^{��B�:����iD���a:�N銛�i�J��� [�Wኂ	���h��=�[��0!=�e���K�ީ2!L�+ˡ�#�����7ATm=����o t��[S%�W#���W+�n&y�Q�g\$S�v�4$�Fgd��P�swz�}+;4�+]ui]̴.�e�#}��ϡy�U
�;fJGE�F+���g�ٜ����Ӽ}a���6�ؑn�D�&������Ui|<��+}��t;>���wv�5���C�����Ga��ӱ�;'b@�V�P�ĸ�z���=}�VΎ�['v�����%��xGq���="�O�;ǳ���Xu��l`��G"��$�{���ފؕ�[�Jk�+�!�s2�
NayP���톜zچ]��>s�xZnw�<���\X�諽�2���4}�A`�/�R>R�þ�tY�n�U�/_��G���Hgkz2:��P�©��-�|W����������5���fG�C���
�ҊWw+��r���?^��H�M�m��{VU{k+܋���U����r����Gʌ����W��S��_H�q��=�K�.���8������\�w��&��1� o�J�� �����^��G�e��"0j�ǵ��מ5lC���{葔=λ�3����z77�S*~�ؒ��rbmT>�y�u哪�B;;���f�ȗ9=�b�ɳA�Fy�\�i��l�c�P�I	��/ϫ�h���n���{دN���r�
�o��w}�Qv��W��u�w��n�W,	�@˛���hk�}@������K��S��F�#o8#*`鎬�ߺAH�ORd�|�S9�D������ٖ��;A��8��Ge��nlݬ�ď`��mK駥�w��ᔬh���I��H�U���¶���Oi����̑��td�,F7c<�v�Ukn]�'�a�Gh�gN��"��	�mTX���f��vz7�3qѽΨvz|�s����gv�����O�tA�w�QC^J��O��;k�Y�y5�pz�Cۍ�c�����\ϓ�B�vvѾ�93�g�{K֡�������;�����<�]��&����}�v&o�/2��Gm��<M�tMc�8����.hk�~�-�NF�H��t8OQ���Ё�۞�J�k�.3�J��q�Ȟ9�*-j���Q7
�ͺ��ң���t��_���c�}i�u����t6����������at�ל��&��V�ݍ���c�TҏVoe,e�.S4(�n��8�V��S.N�(���ǻ�(_.0miL����&�'���f���?��ɕ�*���r�i�,��
���K��������e?\�l�9֤=���:����l�㘎����zl+C����Ğ�0�L*��jR*m4#q5~�2q�^7+C���4X�΍�i���_��n7;���K'o���lb{� �;�j3�_L[[�R��	�t�������|\�E�)���U��uiOpLy[���״nZ9�D�v���j�[���6eb�,��V���+���-�`vԩ.���U�N���z7*�RX��4:x|�g\o�����m��
&�� �MI@.f3|��p��w��|�m�O^��Xeog�����W}�H�.s�q~86��#=�����̂�yW��"�o�$���Gt,^�y�iAvOA��.3r����3�縎j��g,���Cl/țE��q9f�{�r���H�(Do�6LL��EGZ����)c��VF�&��-���06�&z��m�������>&��b$z�"|Y;?Hy�вȐ�eɡt��� ��dxt�c�M��o��k�l��{2M���\Km8�w�<�\N����v�a���vb��B�o"z�*���h�]U�(n�ע��5'���z�y���{jAGĭ��
U��]��,jg:��v�X���\�|�yv���:ǹ�i��1|��;@7�b������R�zʚ�_��D��N��q�!Л�_z���7�����ȧd?7>g���-�U��~S����`�:�ɺ���ᮑ\_�|qa.;b���N�4���j�E�G�:���>��~<��;Wƚw�h߰6*�Q�w�df&��F��`��.�7t���!ɔ��ؒ�N󆨺��Qf����om�g�n�+;������R�������}����{I3�/~�1�G��{��oL��T�ib�����.��VH���v���o:���k���%�^�7�_RXsœ�uX��z+ՓZl�LC��W��*53$�}*tHj36K��j~Ik��?S;<"�w�@��%�q�D�|� �< ����U�ta��g=��sj�k����_/6�ˇ����l+��m%�R�N��3�uH��v�#�b������q>��'	��2;�K���5����~I�q��F�A�U|��Of���`��S��/;�+&5�L�N0uԦhNj&���zlkP�i����z�m�|{&�t�'G��z6�\jQ̃g��PJfo��X�w]����J"}�CF|������'O���V�FG���4���j�==�\c��F��.����I2��u��z�C'�v�H�@���(�~���춆�)��8��}�оt��>Q�#�#�D-$%�;&��x����%�g�h����w��Xͦb��}=�>%؆�8��9��\KK}Gq����\����jO�M����9W�7����Fwz\�|�0!ˈ�v8��OT�*G��%.g3��^u���9��m@HK&Z*�J�a{�4��gm�ʰ�\��:&
�5��K����/qԩQ�ۙĊNmswN�u��;R�:ڛP��.`�Bo��f�Na+\X�zV�+�Y�8��Ȉ��2���9�v&�
�W˅dd�:�VήZp�9gq)yv�%���;G|^���}U&�b�L����|r�+KĊ͡�=�g/h��e`�SRfӌj<���\���v{M�YC��Α��%ɫk���v k=�U�8��Y��p�#�U|2c��mhw�O�踤���=�U�â�ݑkr��}mN��ˬq|�����*�<�U��&�>(yȅ�GTܽ0�d����L]���{g]��j���3՜V �����Q�lm���[�Q~<M�|P�3�~��&�p�؉�FӞ�99Փ���mx�^���?;Q}K͢��Zu �O�:rN�\�|6��xp�!��t:{�����L[�T��� u8���M|=�̽u!����7]O�E�r;�oo_����c���!�Oz&P�'Gg�S.P���ar��5`ir����xo�i��u��N28��:�.=k��og�w�M�(֒��(	�Z,_�t��r�QeӚ�s��p�G���	5�_���F�z;ۗ�����v�a���D#�O��@�y�uwr��jBt����T�N}7X�>�����x��ɚ�Q-���̽~9TWGW�\�a�wY�5׃l���9\{�e0�G9^!�8FŮ��R��"��hk�u�;�����f�|�l�[�Ck鲭N���u��9�<��tG.$��+�	�ܩ�����Fή��va��1��x��;�4�l�8z!Өv"��#�?IC�;��z��쾫�s��6�c`.���efz*��9;����aw/�[YO����ә�R$yH1ܧ�щ�0��mU�a�U�����eg�F�����:�6Z�-�����")�eO$Ox���{����C��G�A� �J��������~�*6�y[�_sOĳe�d��78:#�ܥ31���̫��X�$��($o�zn$&��X�q���_5�#��+�1p���/ڄ�������Ě�;oY;~p+=�5?y;(��œ����Nȕ������Ϸ�������������ꍭ�x�ͬ���0���U�8���y��K'��Z�!f��0שv��p��$dU�(�o�ɜ�<��b�m]!�����x�c����jbuܨ����7f�d����W�X���T����ݥ�M���W3{>��x�憿.}RV]dk4�^���*|:g3�����'U����;E�k]eV�5<�G6e���W%x�]3����zsJ��+�]r[����7x��1e�ۙv�jl��1?.��m��תU�%��?;���؀܏��уe �.Rn�EmG*Or7nrwc�uwl����P
����ΰ�5����&���S�������r�[3�du�%M#���/�:�+M6��O��`�st�w������p��Ҷ?C��P�;>h�x�z�����׼{g�|���6�SJ���T��ɿ7�+Q�{�WE�V��S.M����Z��}��ǌ�~ܹ����繑�ΞG�^�=�g8�B�F�8~8eS�]R�N,ʉh�N���z�}G��O����_�E����c������zo�kc�"���Ĕ8|���.$'���R�=H�=�	��{Bk�u<>f,��=���҆�:�
%" ����~��lz���ޕ.��W>�XW2�v�F����C��{��+g�s��;V��W*��|$�c��N�m�\�$zx���X�u|�ȗ�l�}�ο2<t�!j�S|=z�VΞ����N��/?Dۍ�fb~Ԏ�)�ńw��^[�@����dm�rV�
��q���H�~�i`�Wk�p�m��d
�ۨ�Y=�@��돡m�!v˓B�w�N�t<��:B�6SY7�Ʈ�13}ɒ�=|�и��t����v`��0�ڮϜ�?3\o���>�_K<�U���5ͬ{,Ǵ�1s��١�O%y,F ?���V�Wj��N�5pb%0��I̲�s��hJ���o���;�|�o��ǯ���j�w"ꓨ7����"�f������D)q��A��_v>��}<^�ʝ�˫�ә㝜nX{C�hw�S�o����s�n�F��jc>ג���d�`�v�Wd\�H�nc�R[���j��/)w��R��g^�<��w�z��)�\��o.��^%j%�{W�-��y���=O�䱶6t+��U/�����s�T{åK�,y��=��Al�6��1Wk^�j�g��/����
fp�>;;s,z4�rnN�J����Q{��ꟳ���̨G�=���ön�q�7�Q�cf��VGw����z+ՓZar�|-0)�ms���\I���b��WU��#�m�WA�R��S��7ֶ&��a�G�~�P�2V��3&��lz`YOt���~q�;��u�-ъ�ͭ��\?[�8~uJގؐ̋ĝ-�q7쮋�xM���V3�Ɗc�:S�46�Bf�oU�.^�2���A�$�8�K#�6J���1=��@8�b�뾝S���i\@ևXڙ�N0uԦk���D�t�;�<V�o�3���\>���y��a�U�]�g+ҍ������_���[,-w]㞿Rq>���"��Ѭx6@��>������A8��> (
]��X��r����*�ͬ�j5|
���ق��ږlӚ�q�޳%&�ܟw������YE�;�Z�J�9�]�ګ�)i�a�{Y�λ	�S��S6%���p�SڰI퇩e�E;wWRK�4.�[�qf�ж���u=�a��|���Q7�G����>������ǔMU<�X��k�շEz��t�����&�΁��At�������[K�}�N>*�,��l��A^g��ѽ�#E���!��_CWM6�"+�n���4�PTw:�Oa0�%�{�l����=��/��'�qڿ��s4��#+����k�_C� o���K�9�O��ksP��+Ǳ�FT/8T}�|rp�ElVSg��)|ny�m�T��s&M ۘ�v8�Tfx{ɯc���d�;�i�*�>�f鯍��5�W��P]��l��;�r;�����%ɬ�bቨ�o��3��gӍ�~J���i�<+�0�l�}S�:/{� ���_�T�*�Y�`���ঢ়���p�M��c3�7��k����X�Vk�<Nd�a_M��@�NA�?,Bi6�=~���]�[� {q���z��2������Q�oml[���yq9�
fK�>�6�ETR��Y/۠���Y�����q7��j:O�G��gj��>	d�7':.Y>QZ◱�Ԃ+6�+�ě�)~��j�ĨB&�e6�N�hwSF�ڛX��\�f�u"�o�M�]��(�C���x�f	q떫U�K�ev �j�W�v����t�u��ŵ��ר �y��9Lb����W8P�۰�.�wo�n�s�!-��oo���J����>ř�l4����Y� �9V�S�p�	�*�D�k4�k1�-\�-�f�).��î����;d��������/�b	Ff��"���X�8J��������j�I�7�-He�!]g����W7N�бޮ��6� �Y�|�+:��7�98q��l�·¦+���}/��������%syv%ۜ�w�%ֻ��v���Z������;��ʧ�����Q"Y����*�"'��KJ�Ӷ�_uo�>*�Ѯi]���\3zb\����,��J��l�_(��ww�ޠ�t���At��w��j:N;�pg([b���Eq� �nB��1��Z����"����V�aԆ�ndn����(����b6�I�)�Q����ݡK��Y��^��q8N�1��rE�G�6ҧ�+�f����q�N�$&�����*��S��gf�hǘ��M�NK�6��g/s�����6���{RvB@
�|��SqiT�m��dt2������wx��f�����**tܻs@��n�Hp�6���(���\��j:�bv�HW:˻c�M̫�%���˖;U�LSrh���V���^��#�2�VZi�>��3_.qe8RҺ��a֬׀��t�eJ�@v����W>��d�Ud#P4i�v�pa���{��-9�]}�[�l	 ��{�(�mS�n�[5�,��<y%Gl`�n0�R?�Vvdє.�_�+�T��]M�/�����	��]#.���L�[Si�wH�hr��Kո^X1��gDWV���r��g�hǑ�U5�*Μ����x�0s��N7��� ���7-M��[��	g�����.*yF57!�����s�S+ObI�ņe3�t��D(��r��&��=�X��A��|yVi���w]βܡ��nݾYՠ���=�������"{хX���\�� ���ײQ����V���T9\��Ɂ������[�}CUf�x�Z�	Wח�f�2�_\f䳻y.����r]��=����,^�5�vh��/I�DV�B�ܓ�|7v�����j���8��a�֩���T0@�k�}�h孽U5�8�}x��	[ܱ�H��Q�c�9����]�z�$�wʖ�b������6WM�d�]�_1��S�4�U�1�h�
ŋ6�F�>�*u�Nh���g���l�C��9l�z���e�����;FX+.��Ɔ�:a����A`�λ�>x\��4νv=X���A�	K}�AJU��)�1�V��άgN���Rt>��O_/K�޿�}����IH�9ę!���p������
Ff1�	LD��Ȇ�Ɋ(F8�)�4m!0���1Tq�EH�4s�$&�DL���M1A���d@$�J �@�c&�LY�,�b�0(!���1	��M�@��4	���Y"0����Q�r2d�a�
H0P`��HY�"	4�$I�&�L �2KJ%$�H,Rl�)	�AbH��Q��b�$���7!BBM ��
B9r�D39�7&�\����+��sD�9srDhÜ�&f(�Abi)) ��(4#K2��. %0�hR�6  >�P�(S�wp���pS�8��4fV=̩���C \���'c�x����vn���ۢ�+�A�#P�,�I\�y�äk��<���Q^u�2�U&���l�q�0�d���^��[�P�u>���sz�'�3X"��<*ZGa��Ir���B[�ڙr�mt�����{K���0��|�g�\fms��17�i{x�cO��t��
h��tD��b�:�]xҹ,�V*�9��8j�6���W��LnϱX���3�w�Hx��xñrQ��|ITe�?��E��m��	��7>+�Yr���6��Î��FB�W�[ޡ�_���7�P��f|`C��:=Ӥ�f##d�m�:�VH�����X֝��9�v�P�M���4uG�\8������U1,�� 77yM�HL���ع��U5>#�yH�<�݀�o�v�$es��e���ϋ��5��DW�S*_*;'fH�}���c�Ɖ��jwM�T�2�!W�*h���)~7�B�o����柉f�-[%־�붞w���7J��b騇J�J24�ϊC���<wƆ�X�q���}�!�=�wF&���W���h����Mh�5^�d�|�F�����N�&|x���;hBvD���Y���̙�u������F><���Wq-<�t�]�����B#��йnsQꩥ��*��� k�3mܼ\��-�#+�h�y	6�H♈:�y�`�R���2���\���v�݅�N�X!�0�V\+����X�e쭬ݲ��i�1*�����[. ���EF�Jjd�b��Y�z���/��D�Ebv3w=��-W�C}��z#ʜlW׵t�Ǻe鿇k�f}x����H��T���N�8�My�'t>ڬ��e�ދ>c���hO	�y�١{^���3/9,�#ϓ�A]��h֭�^w<����PBr;.W��ޖ�����C���4Kd�ե�&������Y6�g���I�	/2G{�i�ia�t��;�>	�f�'"��}�.�ŉ]0�X��}�Ӄ^s�\6|b�_���r�pʧ�m�u���E�%�(�/�]?AZz(mL�5��Lq��j9Գ�f`��mQ�/(ۮuU��b�LnG�^�Y^�=�g8�B�F�$���~5U1}uJ����Y�e��O�cm�ڜaK�����n�,c	��1�Gks����kc�%�Y%Q�p7:��l�t3�yx�-���\}S�=}�A2��л������#��=*2�L�u4O�3Z����ցW�x r}��J#��^C���+���޴�f�V��#O\/߈�ʺ���臑�;i�5�ZM�\�qw} MU���p��<���
��G�_��ˢ5�yK00��'<7{S	�.���6� {wQ�z7i^�Z�u���_��n5��O�7]�����o$H\*>Ѽ����}�����[W!Ȝ��B#��Xy7y��Q��2�`�|\�q-�_��Y�_v�}k�wa��|[�1�f73��rܢ|���ꙑP�KSq��u2W�п��^=�>�r�6=u������:�Μ�^����l�|O[2,GO �ˉ�H�l��v˓r{ث��OD�l����@{�=����
��z�C�UT;��x�G���1Q`7���z����\�z��P�O�Y�nޭsy/��K�ټ�Oyܸo�d��Dt�ODahd�ד ���J��{�̻��ʹ^��GIgá>��@e'�����i�{YA�~��������*{�t+ؐJ����N,�	����1z�Yq��!Л�_z���67W3W���T�"Ǜ�3�4��U�K��3����0��M�?i�U�C79�Dχ�:�S�t\U���,
�uǂ���4}[�г�97�6MkY�[��W\��z�wgVq��eN�9�þ�O�b��_.@��wN=^�����FZ[[��V�#޵��>�������>y<3�gN�e��fa��QA`���Y���`|}m��jJ�ߟw9w��Q�G�u�+"���^�k��ݬʃ�}V��\���Y��,��@\t�����6��Ų#ςp�K�^m_Q�.�:�r{ʔ���7Ϲ��w:�����+��tK���~��zŞ�����@b�s62�����%?�N@K�ýv!�z�P�ͭ�r���ס��W;=�*2�q'J�>��5U��[�9��RԖ[#kᔥɯ���ƇoU�i����^^:�\��+��]ŧ�����2����ܣ:3|1�iڸ$���G�!�ܜ{��3_Nj&����֡��c�:��9Mr�����93�`�t*�*�W�DH>9
@�.��7e����_z�HU��ֆ���O��r��w7�sk.���;B��9Ng���)2<G�%�%��/�W�����S!�*�s+;ܭ^8���\5�u8��iƶ�	��5�z�Q4̖P�<L��3�]���g��Kӗ��o}��r�4Z~v����}���8��Ȋv�)�K� ��9q��+Z��`J����9���"�[;V��e����S�ͯA|!ˈ�w�n"GT�+/�w��V��h����ޒ�%Ylz%�h�����Y�R���{�=��UI��̙5�nb5�ù5#��>wsU^��rϐ��&�L"��Kp=8���Wm8���|7�(ws��6�J�+�U���/��M$�t��v^��sez���<N�.�yb^���{}u�� ��;5��Uq�-p�A��D�,R�~ǥmwb���K��RU���]��CNE\���&�����$ی.�A�z�H�����KP�p���Y�qU���4��,�{���k�v������yz��a�+��U�Ɇ�mhwS�9>��v�g���˜2�Ϯ��V��Ҷ���P^�ޚTm`�K�S�C&�C�D,�:������E�C}�Uuzo�'�4��DD�?S�2�Y�|ϕ~���(�Z�s,������&˒�nH^�Z�ȹ�	
8�g�p�)��M0F&���I~��}>nxr��³���]�֘w�g�Ǯ(p�zܒ�X	ẑ�C���Rhm.�Ɨ�.Y5�^e�����7e��P�3OM�lTñu�����:�h��+Q'Iq���ѵ2�
��ʻ\�u�4�pk�s�>����[��kZ���?	���]0u�e� �`H>E����׍+��E7V���\�׽����e]$�����_��8����*�_E#�>,��+�)zd\�܋\r(8%��VsCs1�/�[�����}����1��-Ϡᯝ:�b�H�Ua�w�
"N��-ή�͒��_�-e�hg�c��o��I��s����ܘ�g�Oܑ����~�2�����7�o�9a|e��QY�χ,w8�nK���y��_yx�XN��]I�U�����n�n�=�:��r>��>��{!J��1N]+��^�WZJ�/�N��j�<�M/D}SV�3�l
�<I�3Mu*�s�g�v�g7�,k1q����YaN�+�������3�}��u���
��O��Ϗ�8��`�kA��^�@��E�^���k{�8Ք�$M�eo�Fk�7��������D��w�ɮi��i�yjz��}yi$s���F�iL�ϑ��3�`,����K�bT��^�<�m�w&������Fm��O$���4�b5��d^�E~<N��hv��]����j&b���8@^}�v���w&n6�uS;ÕA��ם�T_�����*�0��N�	������U����?<?��g�y[/�����N��o��3>�5��%ظ��8<�T���d�l�vTz�����Y^F�K�p��.f��z�_L��K9���>�+.�4խ�%�"UU[/S���1l9A'fA��73��>d�ե�$_�Pw�<�&å�wq�eDQ�Ψ��yD�s��~�kY��gB�8p�-�&x+�����a�'����TMD���zǖ21<���@��ۮg�=j�!�q���T>'�O��
��67����0˷�-K����d�߰f������ZZa����8gp���|g]�)<�K�=&�.�:H�l��������R��+�!�����P+��ʽ6k-Iz���Ήhk=A-��:�K�]���2�2s=:��,�&`�2v
�w:uǲNٻ�G����[��O��&�ﶴ��x\�1B�9q�9�g���=�U��^5G�; ���zz,=Ň=��f�9OޟI��:�����u�ź��f��v�u��ڵ���)E�P�z.m8�򑔵9��\���<˿�j�f���&���P�m�s�i�Fr]�p<���ˁ~-o����4�DE�}�>��һ�\C�Ⱥ���֑Ȃ�<W��F��Q��Exy�ͦ+$��f-�S�N�ơA��]?Ku���~,n�:��T�g��m�8:��<V����K�7)N^���X�tW�e�${ʾ2�uFɅ�>~S�����|#���m⦻mE�rk�}�f��~�ԭ��*>#��)�#��\NȄ��B�"Wl�7��@�7yM{�{K�U~�Og�|��=�+�����z|�>f� �~ːk�,��Gi����H��R�O���^Nἥ�vo�A���q`7�Rhv9�rܸ|�ڱ}��j6<��pe�ގ�S��<%87W�e���>��5{YC�{�V�֢��w �`���@S��uTE�Ń�c��U�;�2oɵ����ZO���y��9v����p�mn�O\�)��)P�n�R����o�#ʮa������L�|gEÏ-�np��a�η_K�B��݅Q;N�Q�L���0���N�ݎ���4;�t��[sR��t��?���3�O�F�K
�ΎV�^z���7��\���ȧdu����n��V�0�<��Z/�🧉������38P��͙��CgC����J�����z!�Hr�=Y9sy�k�T���;��p:�g��j7uV�N���x��#��?'�j TËK]f{3�1a���S���^22�_���׼yԡ�y���;*t�Yd�_�a�[���%�6���*1G!f�c�UG�n���޻�{�B�)���p�`K�C�4�0{nTe�hT�Y�H���Eu�2I��+Mu
��Gd�\tުz\�7�5��t�/�ñ䩧0�3�+���琾>�^�%�j�$섽��ޑ����rq�)2婉ĩ��zG����`O�;jWa�����G}	u��m���(� ylA��R�f��-�T����B�:�=(��1}kx^�mf��r���f���M���@�3����( %P}D�I�+�v߆ǵU<����Y^)"�=B�޶ȗ�}�w��s��t���4��R8��G�z��W�ؽ2.������Џ� T�����C(��B�c�NۉڬLѡ��s��.���l���cF����V�|���k�t�yx ����V��[�\����!,��u�.��٘)��k��@�M��h�h�8�e`�Hh[��iW�7�l��zJ�8�tG�u�tzcZ|��	��E��Ļ��8�m�DPv�)�i{��ٞ��7�����娩/�h�Y����'5�C��ϢFwz\��Ϡ���F�!��1z�
B�jsy�L�r��&p�tx��7�S���Z*�)x��J_��ý2�v.d���g����{iM�&�3�QC��F@��E���j���g���Ro��յ�3Ȱs�Ŀ�t8�5��
��{D?�xOI�mt��u�hi����Ĩ���kC��i�t�q=:/ޱ_v���}|حګ{ν���]���*���ʳCFe<��:ߦ}d�g����'YѾ�}��r���qX�.<:e�2�s�3ϔ�aݵ�6�T]}���y�
*���Z��Ep�,r<�,9��'�0ˈ���:�6�z�5��y�Ad-�)]?m^~?��z���5�'Ḩ��xL,*��̦q|���U>�>�vNdB�I��|I�Z|���Sd� !>��Kc�je�����5�ӂ3`
��G�}��?�5]�8g"}��ή�p�gVF�o2<�Y/}�ۡ�Վ��,��#S���E��
�ђ�f58u��8�7P�Naș�ѸK�6-��c]�������U:�g�⫓yW�M���rU�YF�N|�z���IJГ�^���M񷘹p[�g4�\�ڥ2�=n�݆o�#�e�$�2��|�R��i\�wu ���b��⢕���*cF�r�z7����ǻ>3�0�\�iP,�R�Ȝ�\M�r��3<�9z��u?�ڐ��{����2��0��RMçP�\�k�D)��g#�N�Nl�w�������[ 8�e��3�ݯ�&�~�D:O�=�s����ܘ�g�O�u�F���a��}��r�{�Y>LQ��� �0�nvi]��r�!Q��~��Nq����փ¯�y]����ٳ�/?Xm��L�Ѹ5?��=$L�Rj�á���!Q�	���vd	q�W�T��]�����>�k e�$.�����A�å忋�iwޞ�[Q���d���̬���9WX��s�{����ѓA��k�2.F�e��w"��	���p�(�3����;ض�V��Q�熽������7�����v�󼊊�^J�:�>Gn梨��n���:F�(�
���W���+����8^u��d'U�8��<ig���x�߭0�[B�}`yg[O1琐���e���_eN�;�b�ξ��֒Y� ���B�k�4�m(L�q^�ugr�V��Ǌ�

���C6�/�;y����X"�Ee)J�$�&F"}�4ٖ:F��j"�܇	�л0ɕ�	��{r}�µ\Y�y���*����B��*��y�1�9t�=��m�B�������g
g2f�2��M� *xX&�=r��4�0��ܴ��Y�6��U!�:�]\�T9�Tӷ8d�n�a�C�U�fT���f���C�ì5y�`n�2�t��Ԯ�I6c�X��+U���ά��U�3��9Ra��<�Đ�/�[ �-w-���/x�A�� u��Sb�oOV$�q�n�)k;��n�2��z�Y��D�c�1�r�P�z��P��������Χ�I������u�m��[C�6�2�ɸ���@o3���F@εYO��U���l�,}pe���7���v�gfQP���h��r+��޼k7��w>M;�<�m�vmc���.b�zn7�{S*b�A֚�Ѕ]�#/f�vS�FT(T��ر�*�0�.��v�<n �䷕���fNj�e &5���׊�..�u�޼J�*~r֓��lib��
�{NL¼0VA����箆v�����Қ�bC��G���PVu`�J�@Z'U�6�8nK����+�Z�7�'��c僱.�nZ�Mo�Sy�@_p�b��9{��T��rDlQڽ�9��T�L�X��aC~�E0�v�Z��2�%�w�����Ê�6���S�1DAz���.��X.V
40�.�±nR�w\��bo3m^u�|�wS��;�Z;6��gI�AJ%ԓ��vn�M��k �H��k��HHp��=�y$�;*��x�J����-��a�,d}����U�hs
Ben�0UZ��V`p�X9���wd�QyX�;r:�l�3���x%H�lዥ@�|v�ZO}ҳV�f�qU�f�R*󜣰�5# u�r��{�v;[V��bd5���7�h��j�n.���e78�S:-�\I�k,, I��/�n� �}�`ͮV�T�Σ�Gh�:r�#m��]�J?�ό���H`���6Ʈ��Rou�&*�;��W�pc�z-G�~En���xrϋѴ��:�aXk5���K�؛RPJ�6�b�e����������k�'P��d�@@��9cMh#/�=��Ȯ�Vz�v��I8���y}�8ZT��\�
�K��p6�m_A6��T	4��W3iY���۽V�_;Ne����)b�I�iђ�\WZ�TO4`��F�\�/����������}�0&�[�u��`�R���yO ��0)c<2��WV:����[�˥�q����',���`���j���y�슢���o\�[\���u/[����.n@t�}yjR�YYOJ#�<ݏyN=�wm��sm	b\zi�����8ަ�c�@tM�gK}hS������>������wK�P&&4�DJHH�FI�63#&$A12) �"���
�03f$Bf�M��3(�F�cF%(�4�E�
4�2%PI0d����cDHI��(�2`�b$�dA���D�LA�&i��b-	JD�H�Z Q##R1�	bBe��cAI��4��F뜋!����)(Ŋ1���5�iI� ����1�@B"Eh�(�b)),`��� eL�#�H���i���RTQ@T11d6�&(��5DBIF���ƊE
,��E����#62`���F���3(�H �Re
Z"H̱����\뿞��{������(p�z��%G[������V=��-k�jVپ���� ���6�.Uro�mA�ι.]��%ԁtD���`g�¿0h7�j��/�?�g�JS�3/9,�y�:�r>�kv��:��(�כ�߭���ذ#�ΰ�5C�Ϩ���s:k�+̟ĸD����s,��beGl��wv�'��n�q��H�c�y��Y�i`��9)/a-+c��\�9Pv|b�Ю8��=��������b�e���!ڸ��X�VvT鸲��,e<X���Q���:�(�k��z1_�$��5c�+����sM��.}o�H��^8(�'g�P�iL��:y4{�����O)�7S>�W�	���cźȼa6r��1��t=&�Ƕ)���6�GD��r����M��!r;ey��mPLӧ�&�]��ߚ��lc���A�FX��6�Q�����g��I��^� /MI���7�l���j7����M&��6+g�U��>�Bg/N�O��n������/Y���$z ����2�p1�����qo�!�����|V�:�/o�6�zr���+u��9d�ͺ(9�TOÒ=�FP��B�{�&9�w㕗�k�
��	�e*�MV�c`n�쭫��8� ate����Q�t��h�ڔ'N��%ˣ�MKPd��L^��9cر��qT��9S��Y1��=m6C�{��>���6�m���_�x��C�bʝ]Y�y�}���r��%fA��Eo��-P�1�G/Y����V|s���'�3"�H��ǉ�ul�f�����{�t�l�I}K;T��OC��(7ꩊ�K�8�v8и��t����w/r(��ĕ��MF�`�ȕ�Ò{�O�hv����7�d���C���a~�QAE��ݽ�8f_V�榠�y �a\����k}����~����0�?]��}�ԧ�$5��Mz���[}�}[��~Kr�����_K���6t;���WO����s�T{G�ʲ��%���u{a��}����[������Y�����|vv�g����(�4��:����l)���3���[~�2�� �S����x�~��՜b��eN�9�fP�"�m?15�T���o�7�ƕ�>�;^22�_���׼yԡ�]�;*t��Y>@y�k�<ǜע���GVW���Ә��fxF7F(�����SY^�<;'+�s�C"_�kj]�X�-F1K	,�>� �H{%99������l4���^^:�u�Á�w��^�X��d?�)�r�5��Vo>�Pu-�6(��wp�˾�W��ѵ���d�V�JhWS^�wlL�,VȮXiu�G��wmG���u�����[��˳�`�C����D�����B� �U(ޛ.�����U+쓩
��7<6�
|	=S,	��:���rq���3AӚ������9�G������F׹N�C�l�S8�g}��p�>3����F�<��&��<q�알�T��e�U�׽��N�Nl�.}����õm�9Ng��G������-���]I�� '�1�;�૏r�W����G�������O�������a,[t��x�";��^�����쥷k����D���$��K�������Y�sĿNM�ޭ����
~؜�30��L����ԤA���=$���)h��~>�&3ͫ�~� ]�\Dc���"�W:S�v�n������T�3�'�'̄llD��qYKǬ���i��yA�}U'�+��渱�!�S��Uw扢�H��݋�>ٓQ
a������Gd�aȡ��N'uv��@��ٛN�ܝ��ALy����.M��s@n��ixU�Y>��z�'#�SÑ��{g���v6��u�Ov{	|M�.�ګ����v��5ٮj�ɸ��<��� ݊��~	�RL$��?��s�:Z�I�	^��5�8]���U:��,�Y��Mb:x��v�Z���7#כ�՝���iMv�����6�F���뷄��ʳ]3�k�k��w���o4�Y�kݜ���p�:���+�w���ʎ�&�`���^Wp�&c=�\o�^�r[ W׾W�:�^��������Q�omlH�r�Ύ�>���[86�дw��V��ٟ��C���5��>��z"&��v���6��R3�X}ԂYъC�Y���o���c�=�9'�k���	;0u^Ӫ�_N���:�u|4��M���u�(��1o���f�%�2�o`mu�u�4�F}MvB^�?B[Cje���L.U��sQ��n�����j|e�Ck��O�>�1Pe����y��ǻ��{�E� �,ȱqs�^B�؝��rN<��j�fK������G���/�sv��l�du�|g�I� ��\���r�X/<$�ey(`rY�V;jBt�{�β-����j,�5�l���$�>:=Q�6I\;t����b��_R&������}�QJ}�a�W���ޮM�{�G{����:�uU�3��R_�<Hڜ1����?Ku��h�v��_!1���>���-���{�-A��X����J��Ac��@�s��$����l��&_�
���G�hR�o�r���iD��D�r+`�5ܷ�U����o��FԴ��� 
����D�1�Է�8;r+�8��Pb�͉����+C�ۦ�m.�I#�>Xs�u*�@bh;�p�G���~�Ie��M݋8�W��7�Ձ��sWG��"�͖�[��ʋ��x6�d&�"C�d��*Ӱ�Y8-���BCx�,����D�ʹ%<xꟊCξ
�T����q�Y�G{���=�4����,{�Ly�L���4�b5�!Z]N���Z�!;#�s�⓺�sw�|}xS��[�q��c_U`A�߮�Wc�r�. ���y���K'ʶ�2�l��UMK��[����0����z���o+��}��ᐝW��}�4�}xv�-+��w�Nԗ�5%���� �>1��ߦ����Wa8o<����Lc��k����(���yn�o�Wj�wx��뮉�Ѻ�9@��g#�ngL#�O��\"E���Y��k�������kس=|Q>�g���$����}�:.!y9A.��Kc�6��ع]0�f�#�U�zV�x/kٶ�)���h>�2�۩�v�W�n��{Ia�<K��r��¼��9�8�/3Lu=��q>�ç0�X�sQ�0�pb��r�/�r���z��g�s�T.ʔn"�$�&@�iC54"o!�_%��v+*e�+������~-�E�	��j#��7]M�kc�����~~�V�LZݹ���s�p̴�Y��]l�C�����u���<K1��c���a��Z�
5�ʍ�wj�
����	V3LܟswT���Ж��7|�2R��;�x;�w.�)]���]V]l�Fr�p�2���'����)��pzl�p���:��QD��4Dn��+�>v�˗�'Bx�9�������{�=XC�5}������ )���&u�o�˸�j����%���x�tF�|^X�Җ�Z����bu������Όe5<T�R* El����끸/ō�qf��$A�p����Ӆ�[ޮd3[/��	����eD�G��݂6L$|��*pI�����,��y��Y�}҇��������ߨ�e��y�#:�B�<���<����h�4ٸ��^ߏ�!���5�^�Scޗ��Ï�U1���|!���ΥAQ���xfR�F�b�7����Tu��!.��7��;7���C���7�d���C�n�F�9+��72�ϟI�/�{iAcɓ郃�F�b�[�h�>�J_��ۇ���Ҭeڹ��w�^��VV8��O��u������g/���PrXQ�C��J��<r;������<��N�}ZjוN1�ᒧ�����������o��fp�>;:O�큳��T�X5� ������#�8�w���+S�h,RB�.�\n-?__F�j����O����:lv��R�WiU��MNg�©ka+����=�uI`p�S^e�|����Oe2�پ����K������w;+����q��qX��ç2����F�ț�z��W	�?g��N����F��6�����n�:�ۙ8#D���u튛�����Y��#��d��'k�F;^�����g���'�}��:k�{W_���:�J�AB�����0�ѝ�����=N@mD�؇�}�#^k8;���^��=Q�Ed�lv���[C��C�ZI�c���zGP�R�입�GoU����c�^^��1^�n���Koѯ��RT�dNW`�+��'I���u���� �Lӧ5��\�r1�ܼ�z���qy�zlg�3��P�e?��Q�*2��W��Wq�/J���ue�;��e��Q���-s�FE���]�Ŝ����.#��,��	Q�Ҩ����=5^��}'���c���l2�=C�ף�i����Ӎ��t���4��S�&�Mgh���
dn�9�����d����k��^����]��=ϫ��n|K�\q4nt��ascY1�`t��i�D�6e��G��:� �rj|��j��9��*6�W�7����B&|��{�����rc��tYnৎx�����/o�O�4gm�.K�þ�Ź�ɗN��]:`pკ��}X8t��)�=e�j�s��ǡ�'3z>�.�
"P��gf7�3�]N��c�x5�`U��:�T�`����0�t 0�8��A]��2���O� w�@5�E~��~'E��pT�/�Eme/����6׶��ϼ���u�$-��-&��l׶���M9���9U���C���]���W��W�]��{�+S�2��y����Iy����U�,v�.M[]k��,�i�7�Ī��_�6�;����0Ϧ����ixk�pz)z�OdoS�κ�q`y����<�g���}�q1#��Y��������ڪ>��8�������w��٥Z�˭�+��+��u.��������MF鱶�'�u٩؍�Ex��=su�ڸzKQ���_:̞�93�I~'�i� �M{$:/ޓ�Ų�ld��d&�=�m1���B�%��Ӓv��X͉����B���tg���Q��w���_�� ��מ�5����F/fg��u�:��G���7'FےO���q�U꘾�B\��?1�^���
{:_F�=.�^�>��u�Ui�{�qnH=_`H>E���w�F{0L�=�L��:];��}<�o9q��5��9�;M��V��),��������,X�����f�	]Δ.�ns��tYV�uz�����,�ʳ�jf�<�3n^.uˠ5>��Q{bAW��ַۊ0˝���:���)�e:r�FT���Sf�AmBx�lK��w�z����l1��p;8�m����,���U�v�}]Pńc���wVT̋'���Ԅؘܺޞu�a����j,�~�a����AJ������Q9������b��H�nt�Լ�f��C����M���w/�p7;Nwx�3��u���h�7W�#=��p�$�ϑ 74}$L�\�� �9��Tj~������C�)�=>��z�FZ�z{�r7YA�eOܑ=�FWq�&/��}p��<:~/+̏�к��]�W^v���1W�>��i��l�l�c��D�S"�g������X=�Ad^�J�c�O�ﯳr�Mxݾ�-��M}�ra�o�RE{�ѓ_6��w���D�8�ش;`;Y2����l�+���e�!�y����������j�C����Hu-��/f��(4�;�L�f�kp0���o	LdǶ�N�.w��q��W�ö��9:��}�a���upt��(E��v�V�u��xl>�/�T]}��� �{�|s$uM��+��7�\�}{^��L��K�Ͱ�-m��͝9�»�ԃ�S��kV���,;e�:EeW5+ģ��c�)��'�oKvY��ek�ice ��=Q�԰*tbՕ�˵|.k��x�zo Ϯ�}Ư�q�I�17@m�0A�i*�eɚ���_I�)����Z����y�����N��yBL�k�w�.�J��X��2�9u�-vXDJ��[�ziz�g�꟩���_��;|���~��"˴�(y��(%�s	hW�]z����ƶ��j�^n�b͕�JX<�#��>kY�,:�gz}#3zo�M���1ĿA�q՝B��;�ӺUc�ST}�Ϥ��{�5�GX�������?W�VW�v�0��Q'3��S�|z��va׷�'C�`�豵2��܅�=�P:��n�/O�^9��nz�w�0��+��U�ⴵ$��$����/�;et{}�A3N�К]��ߚ��us�4Ủ���-9�Ѿܿ ��l��D*����H�j$�&u�c�e���ÿ+��uO��>Yir��}�X6��Ӝ�õ��F2�S�O%��U���-�_��S��+�/'}C��v�̖3\�i�=�sW���9d��(9�Tq'����#d����&�;S-a�{�4=��~=�����+#m5n:,��,�5���fE�����ˣP�V�|eXN+A��g)�T�7f*s���\��X�C���b۪�_rT�p���ն�m���mZ��j�V���ն�m��mZ����km���խ��um�[o����m���mZ��Vڵ�����km���խ��[j�ۚ�խ���mZ����km���խ����V���mZ����km��[j����ڵ����
�2��]�� ��������>�����
.��� 
	*�!% A%"J�DPU  Eg r*��R�����)J��JJ��R�R��TIQ 8�J
JD�QR�" HRD�)	JR��J�� �71ҤM��J6[��+X�RhM����UY`�X� ֦�v�BQ�		��$ڍhɩ�4c+ wX   ̀  @  wp ���(].;�확�6$��6���Uf�Zͥb��f��Z��F�j� �H�&�6m5����"IV�U����fV�X�Fih�Y
�kM�J�5֨ ��0P�(�(*��7 Ω:̓A�
$�j�J43j�@T�@[h F̫�u���h2��,B�n�8��  PM�R�j�
$�%�Q���(( J��TVؒ��T��m	n��D�@�SmMiJ�@"��ca�Q  �P�hhB ���T��,�J�p�:"J�`V�����dS���(�l�֚Vl�1�e�c	4��e�S��:m�XQa�fْkY���[��Sdƶe��#VY��*�
h%[�s�af�(fj��H��R�6�$5l��l
R��     �J�*j�Hd�� dhi��A�B)�)JJ��!�� 4�24@sLL�4a0LM0	�C`F)�b4�%=T   2   �12dф�14�&�) 
HИL��Q=MG�=F�SF�6R}??��f}�n�_�����u����73[]�B�(����i0��TD���8 l�?`�(��M��?ز4�
 n)m����������l��z��H��
"�@v	�("�ȚIa�)h@����}Y����G��?������AD@���:�Z�|�`��3Oه1��O��;M�1#�?����ޚUd~��퓋�ƺ��-&�7�f����RSZ�TǵnػR�$l���щ �0��*�*i�,
or�B= ���K�[�
�kCM����hH��ˎm-0`+*�㉆��l�J�d\uA(4p�r�\x�'�]����v�n��� ���V�m]��(�J�����U5�-�8���n�Vj��[��e����	b�^2I&�n�X�+A��v4���Q+;7<�����Y{z��5-7@ްB{���(V`є����4l�r��g�f�e�E��T�5���Y��C��X��b	:Ҋ����m鳖�Cq�mm֬;	Q�R�$Cs!���ʹ�H5f�f$�B<? ��/)�dY�	�B�]�7whL��;�VY�v�޶���*��I.�r�An��q�L���X���ʹ�f��&� ��0l�([v2nQ�iLp;$f+�{���m�Q�8�;Ы��[$��<��꼱HS�^�F���V��m���;E��^�Ef�@�]\�<�Vo*�����X����x�g�eo"nÙe�H��w��D3NE�j͚1a��X%`�/P�����T��-}�H�)�74{�;H�J��ӝA0x��٤�-��צ��D�HR;�k�S�aY��%���3#F�TAJہ��Gp�o$QÔl�7{��ߤƉ̺ۧ����D�(mZ��g�t��(�f�V��V+	�+Yˣ�kz@f�0�Oi]�&�fi�4!,�6�d�{��ZoqKZ��K�,	��.��7q-`Qω?]�:�b�qK:r��H,���@Qk�*�mf�=���f?�G������V�f�'�n�+j��;i[&���F��Y��\)2�/ym����VA@mjtN��=�"���^c�e9D#7�l�f|����bV^���V�`@�X����z�w0�L�k*�v�%6U�f���U�-V�X�)�L*a{�r�¦��v���6��
eǨM�DйSk�/Vf�Gu�z��֬ǚ�`�9عs"�����V��$�M�'��ݧ��]�z�ݮ5�����ز�H�	���GP�a�NlU�M�s&�ol�Xm�������,J�x�Z�����H�[�t��u���r��U.�ׁY͙Or�2�]����2�<�ޥOPIRvt�7k(��4�i�y�<%��I�ub�G�i���Z'
h�Ց��O8��4�7d��{B�nĖ��������J������y)���Ê&����&����2�4����
e��l^օ+p� -I��2�5z0
Z�]���ͦvЩXa,���ͺ�3q��?I)2.���i��������##ۖsuV�YtE������$R���.駻�~�43,ē�D1�,kz�=(
�0�f-�z�n=���J	�'ܙ(P��;L<P�b����6��b��-C�6��X����2�]���8������a:~�'�J� ��X2kbwwq��!r�e�#@9���y�� ��2ɻ��j����ju�	yA8Ԇ6�.���%L�H��\�sLZrD����+��~WnfLiӺ4r�T��Z��&
 �f��`Vݨ�V\X��!����KA/����/{n�!�(:�0f*c.���^Sݳ�a-���"+��#�J��7,Jߎ`��ur��%mc��^r����㆑��ɲZ���"�sTG`q��}�e�X��{�Su���&�+.��A�7:vj�4ct�$����C�Դ�yø]�/�֠3�K�r�k�� 0� ͇4��R׏>C ��+���: gp������kCP��sDzr�9���Y�����ٻ$��f���/�]Ol���z��٭�{U%�1Yt�F<w���6pbNl�tn��Lډ��`�,��GkoHֳB����9�9��އtT�:jH�չ��/n"u�֖����YM�jĵ�̰l�ͳ��@��VSxO����׵��hӫ?F쑵��x�`�2c�N�k�!7�\��h*��N����t���wZ��D����`H��5��
�kX����˿�(n��ح��uzNh�	nJ��ZX�놎�;������
�c0Z�u�Y{�b���O�y�H"Qj�bF�u��|>?.pj���M�DX0�*Ξ�{�F��H�wŅ�WvY�X2*���Yf��hm#jS����L�5��X0�6$��YXނ1^���lӤ0�4�X�V�8Vb�u�7o6����!HlH�ɀ�MQ�k@�e�J/� O�im�Gu��,WD��S#>��(�B�t�^&5Қ����HK60٫ʲtAN���j/h-ժ�5"^�Vc���s݂���׈I�U�շu��}��1'������U�z��6�4���۴�'VK4��l!h�y��j�.�����/t.�L�yK��a<ջuÕ�]H�����]m�d��ѻ�`%N��˰���r��'�kK��iԆ@'�l�C5���+��w%1R�(й�z��Ǝ��Q)�����w[����)Y��V:5�Gת<��aL��P��c@�2Ӧ��V�a���u<�ʰ�(,�6ͼ47�:�,��-Z�����-IoR]a�Km��:�C0U�I�j�4E#1�2�������6��GTx/��6�4f��3q�s]"KɫHjP�����K� �*�:d��Ʒ.�8nΗ/v��kDZ4K9���w�Y���:�d�P�&:�m�hS�;WYr�*� h��N�Yr�KYͩ�S�J�w7W©�E[�`
%溳յ��қ[�PAR���Ie�* �[֝aᎈKV�z��<��֚��'iPհ�t�6�����u�L���ȝ��r=%]�k���{�Щ��w�9aђ��U�O �����6��*C7�f��W)0���+v��j����B�:{��P�u�S5+��-&��EՆP���=��n��XՆK�A�V�͢��Yc@cC�˟t���+�d������EX�۹��i�4��u6���YgP+.�YlJ��h[������qc��gu�v�/mӰ����
�a�@l��j@���2l@��ԓհ�[�0\t�T�QjJ�K�N�R�5��VQg5%XѬͥ��(ꕊ�T�hY�����)4U���,���˴�lct�U�wYg[�/^���lӺQ��Ve�Û���]c�3��י��m�8�
;d��-�JXm��,��/%�y�b��!�7q�.�F�4rQ��cWK.�sڈ!ۺ
K��q\ב�:E�؎Stf��
��R�{���ݕ�pљ�����9���$��P��!!�E�ú)��_x�j,:���MK:m��c�X��%^�F�D^�՜�J��n��f�m	)8 D�%��1"(@�
έ����j��IOu���@�%��J�x�}��8��#E�lea 2��Z�(���$f�b�w�������Y��w���i�JJ�Z�s.�I$Fؗ0�'�ɔi�jN�P�w	����5l�8�l\��yV�P�j������'wjLB;1ݷ�Ɩ�U0���@6��
�y� p�#��#SӋ �X�{r� R�z�՗d�F���i6��.����P�̵��;)W2pm%4^Xv�c�@T��A�{u��c\knw��]s�o�8���<AP=������d���m��n�Ӈ)��`��?��������q�ב��ؘ�z?�?����@                                                                                                                 `  `                                  ܐ�^��23�%��`E��\�%�'�38vwL���������bU�;0�\�y�B�+�(�V���<�b戨���.�Z3���4�Qo�Z�*�=��Kn�S�٢j(M;me`�+��S��`�Q���T�J�#1k)޹�b^�6:�r���̱��rBi=�X�Tޢu�uyyٖ�W	ڎ��7I��¯x|��M�
%���]�>V;x��zNt�F��o_L7oCE�d����FI^<[-0���}lC�	�5{x�%ݴ�%VVW;�H�pZٗXv��T�A���;�nY@=�}���v����*I�6���"�w�V&J�9Yʎ�OMt}�Gb��g^��Jt����%��;�{=2y ^����������A	j��%��{��9���G�b�~��O^�/��`�k@���U�7x�XS�|��ͨ�)�Sت\�ӱe6k�:�M"�:;ܯ/�I3I3r�����Wy�FĊ}e7�f��@Ȥ`bڝ`��mP's9��Y�m]r��nKhe[���Eip3a�o�U�u�v�N�ta��COt�t�D��niN�6���\]諧YNm�7v�5@]H;�����X�V`�X�w��-��"�Ms4��Iu"��$N�]����N���0����ݽ��#ֵc��ݢ���ΨoNV���wCu�IFΣ��o��8�yfL�;+V/6��֥LR�P�(n�};9�[���Z�|��/,Y�{ֵ7�;eu�V�0[��@�싖��<g1q��꾔���P]���g��yR�؋
�irT����4j�5�>�������\wsGy]�3�]VS��ѵWI�W�A^�x�����e΂P�6Q��b�c���خ����a�yh�7*v��7Y�us��s-�K���Dwښ��v�¹k��q!e(�G�IkZڅ�yb�u�7ȻS�2�n�	�i\��T.��(+-uk�9�m�i,O��������ud�6ј恕`ptq��Ƕ�KB���ڻ��A�]J������F�f�Z�C�\�\��w�yz�Ԁu���3��D9o��-��D�-�5Sb�6�4l
���y\
�!ҙn�`Mi{�n,J��p�q���ͧZ������@�F��#��Ql� v��=��$��,���y3���X�qL��֞T�'^���88oY�;��-�xH�b7`�w����9�p��&�����.u˫��-J�g4X��l-�'ZʫH4�u��7QE�����%O+���֝vq��s+���E�n-�H�մD�M&*���x-\�8�z������$�4�v+�����oi�d��v������f�}�Y\+[U���}F�ڽ=��uZ�{���#
L��,.���%��h��V�9�l���	�<VH�t,�@���77�/����zTR�z����Z@2�s��ﺧk����5�W]˵x�OB��1�X3Vr�1lyZ��HWv<�����2<2����C@VU�P�� (���r��3��C
� k���ެ�.�GC5U��X�4�
�WR�`��2�.Ŭ:ے�"����� �8�s;��Z-Z�x-�D�޺h��DPX4iΖ��o���qf�z�,�R$}�}�&f�hN��d�k�ʀjg6�ee�9�7�>IF��J�"��¸����1G/����(��������x�r���Qf�vI2�'��雜Ӣ�7qt�!�2�5a�]�i���`�=����X�M�U�G*�o�䫙�l\��^aqu��;�����u������nc�{�G=1^��N�A�ҔZ�Y�#S^m-���*�׶�Eֹ�bu���*��=w����.^.ԝ��R�Y�#�d�3O\x1��a�2�8l�Ica�u���2�s	��ܠyt+��\�tB�t+��O(�e�_9W ��[F�b��}�k>X*�'�.�r.���8�/V�dv�� 9�^��	�y�q�\�������w+_���&p{5�l�X�>����h�R��[FGB-�;��/����0֊���5J�n���8'�dea��@$�@�6��\;�igb!�KO/���L�}ؓ�9���,{���������B�+R+�Fk{��t�kZ�繁y�)��7c!�93-��@���&d�V�w%��(��W�80�J��t�ђ�Wv�d��C/��}ZJ��f&.���J� �X���yZ��x���GY2Ғe$�c�uuO3�a����|����\���mޫc�%-fj�bS	2��rfT������h]�wN&ˤ���g�
�+`de_Q�S2�Zֺ�|�x5}��b�j�w�{��xw��wƎ�.����t�^�
�(�g*򷔖b=�$̠!c/����t@˒LR�V�8�f���H�2�n.{��3PR����+Wq����p�Vwl:�zԓ�����K�w�e�Z-+.�fi��gNѬg����-v�j�jلk��[�W�8�M�nPTp�O:���{us\'b�{�Y�k��6Ӂ�
={M����VHQ��+:�Zn��Ε�q&L`�VO������^�h��v���rF֬�Ćʐ��_h�Nd߯5l�#
��0Uf�v�k���JSf�wwv\�KU@���B(�b�iCǻ3�Ѵ6+\$Q����ȯǝ��7b�EbT�94b��^��7��-�M̵�sK���ob�r�yl���,�[O��u�7�������SS���#J3Ð�B�g=���'8�l9�t���ay�{Z���a@\v=�n�2�`�ʦ�M#ܱR�}�D�7�&�ts���9�j�J���ˤw��I����M����.�d��H��	�8�8�F��y�n"fNV�q�v^!o��l��|E���u�o�N]Bd\�
oj��$m�Ԁ�P�O��h�SB��9�d�m���4���ؔy��f�溦g4��F�B��*�`U��SGU��݅vk9 �C-Z�r��P:�R���W]�K����hsUˢ[�Mm�p�<@
*�s�DZ��{Y+2N���^L���/͏I���1�����*�b��zV�!c�l�����Q��,�Y�T=��1@C�C\fN��=���ƛ�9 ��s�n���P�*7�0R��m��
���%|bq�O�$��/t��(�֧-�ᡩ=�����{<�*v�g99��<ϖ�2np�,�����f�+v����pj�F���r�>��b��`��,x�r��0/�uEW�Y.e�Z��z-k��F1f���Q���^�3$�g^�E��.=<�\�N�"�G�+x1��G�&�E����˳w4���roX�����=6�cV�[`�#�P���*�ĥ���PnF->�E�3P7ٙ�����Wk�IiԂB��(M�/� �\���7��0�x�r,��v].[7/GmkPXP�Ԭ���&��59+6��lJYE�QZ�q�uw��j�+Bӡ�3jT��9��-��'�$�7������n�                    9  r   �@ � �W#�g����^�-@!           @�     ;�����~ϙ�n����ߠ����7�DTDԍ�כ�"(.;Ш��y��?�M�D�~d�}?M�ӵ��s��8�>���Z۞z��u�h
Gf�����t�ݱY�;��#��9�",���&��M�Y�9�lh���Z9}{�Xn�ң.ʦ�6U
(���u�����5lyݝ��B����˺�c5r�m�9�w��\@��;��^�A��#��j[�L�X���HU#xl�Y�D�Z��2q��J��U��7�W�<f*w�jU�=��T��VWK��e�
%R�����{8��]�4��vܩڐ+,Ϡ�/��Y�1�Ю�v�K���g��Wj<�뵕��a���mw]�4C��*���G�\�en>'JMݢ{t�q.$i�0�4�9/�l��w�kPX�+Q�А����[���Y �{|�m�L�Z���Y�'<���(!�[�Y�p8L�*�Ma�X�\#��T���vv� �ޤi��pK� �>��;_*#�v@U�!���R��S�P�!�8�U�nZ�u��9��Y�H;$0�6*]��4B�\�A�@��������5�Aeug5��{���Em�MIM�-_��j�1I���a�������|�:�P����M	yն^�Ѻd�yi��`-S�`�F����J�i��4�b��g�*%Jf�]��q6q,�:aKUGr�6����-�`}���Z�B��7�iNv���&n���4F1A\�����������^KY��bTA���M�5�i0����l����;i�EE���6�u��{��P`���ʍ���F7��܏o�"�haA{I�{��BXyQ�W0��wr�cU���/��o17�XZ�d�Νw+M�]	,��Knc�Q�������Y�K!Z�����b����vl��Rw���P��/'<�W�Ҕ�����
{p���O���l\M�[5��o]MϮK�w_dk�V=�ʖ���Fj������c�Zm����unq�ήʲ0U�7�Hϰ��ń'��'^8v����3�+~TЗ+��w���<)w��F-��K6���`ڼ1Q�I��U��1O(�[ǫ&;��x�������ZUؒ�&��\l�
Yj�V��۳�4���d��0m�j�ݳ� ���f⽬��_��S2�RE�k��^J�؛5ӤT� jE��j�ɸm.}ͪ��[�:U@;�X�i��iֽ�C-�9V�"�𮚂9p�p]��{Hn�mk��T�%���[���J��!D�u��d3U�w�Ѳc���^����.�1.��ʛF��Rb���^��mh�i�F� 6P|���pu�{�|�<q�ۋ��y	�Z�=.^�-�e�<�������)rQ%t띹��u�Ũ^Ί0�.��Qw�~'����]��@��f�(��%�o\�ۚ���il�B�c�3v�I�:�1U�y\�b�1].O��|���k�̤�J�.ܣ�f�B��ֽKs���x�v���ǀͦ�����s��Ed ���9�v\�"��׉��X�p�\��8�:�t�Y=�b�ǀ�+����.8γ+1U������W	�������(�;��4�Շ��D\/*���25ݎh��:z��/�4��ܤQ��٭�G(Ms�]3�t^��)ޱ6����5�b��v�Xu�{X��f;ׇ�����\8���X�����T����B���7�s1#�;[m��[SZ��6�n�ȁL�K��;����'��d6�n�_B퍉�Sn��H��k8⦥���=���.��'�_��4��9Z����"�v�YY���&�Ρ�$2��q���A;�9��oJ�mA,�:�g�����.�rӳC� ����Z�ڒ��.��3�S!�6ܧ�����h1����Ɏ�1ҠBPe�]��� I��|s9�����L�f�.��WȾ|qW[VŎ�7s��!�� ��6f;S��M
�i���b�A�Û2��L��7��ШfJ�1�3�.�wm֤v�ܮ�eӤy�Ѳi���ZN֛��K�._]20i�zIk��s^�c�f�\H�q��1��b��Z����-ћR�X��&�rQ�$��V�3�.���\.����7�¨T��׷����XKqY�:3��c��FZ��l��*�B��E�|)&[�����`��·s]Րq�����GSu�,5Y�>:�re�/�P����
���F�6l5��t�0�d�A�G-�E�5 Z���@ãn��$���ӛ@-V�ӡ�ҷ�=�*]X���n���8�%�+�(b��]�1*��I�)5Zx�i�B��ɘ�ø�c�
��K�����w03)u�L³�5|t��t�۫\���}�EHn�_Fj=�w�����A���uŎ�ޥiwVD5��ee���X��X�(a0`F��������%�:��ɒ�l�;H��.��;�Wv�ب;���R)��7�Y��es����-�����ö�"�`�b�uޛ��:�M�97�#��N2QÌ9g*X2��'�AxS���*ւB]�$�9�ۭ�}}�/��Vn��@�"��YXE���nO)�s�*9�!�yS�I^��w3�XI1M���bFgN�%���1���4�n+��&�ax�Zjb�G_Q��e�kE��GF����TJ���|�q�Q�/�u���gu���'6���xı�+&�ܝi��e�R��øI]���Q5��!h�W¬�����Vr^Y�N���|�� �zH�∛�,�[F��� ��˖�P(-ɔ��4�E�!��"��Dw��l!e�Z4b(fn,���hb��^I&�T�C���|���sga����ڔ������;�&�y�6t�3����������6vm�Ǭ^j�7x���V�C\�U��Tf�JF�!�K���)D5]�; 5��۩R�������:2���M��3�(*`U�ǐ30��Ku�7�J�f��[��ݛk~L�����S��+��ms-s��+������*�k�i���=�O9�%,a��7���T�K�u/�ƴv��gqLTG489c��e�=���ʱ�NZ23�V_K����VMZ�q�P+v�젟5�[v�vr�͇�N�ywhq��9��n/4-��T��<ƶd���.``it�߉'ru'j���h��a݄m��\o+\�v��9�.�C"�K����c�(idvԾ�����ʕ��i\l-�����z���6(<��n#ۄ�U�c����v���v��*�h<�fwedgr�J@���<�I=��G��"^�ISջ�*�^�S�D�y�D��
�ǇI��{,�i��TJ[Z����Â�m��ٸ����wq�S�[�o�g2��Ǥ�hn�;��h��[V��h\lt@J���b����i�Xn�o+��fm8�>n�^������M��V��+K��0:���J��v`�
�S4�H�B�u��[u`���V��.[Ǖ�9�t��_2�P5s�4��U�DWW
;�YV\5�o(en�oM筐��j�D���Auv��7�t�.X�Cw�'������/�m�!�b"��
���,�M��u�F�qba{\u�Ms�-e&���Ia���s����+z�1���I�,J���y0���!v9/[�ե=�L��@�Q�lَ^�{�cƪ�����|�Dp�h%w�e*�܈uo��7(�9��V@�z��t�	x�q
��쭫3^���0�������
���hV���g~���?������R5���MD�v����>���T}1ﾏTV�%�            �(]h�ԺH����̢{en}xf�������q��7v+,���hmB��r�f�QۅXW5u�֪5��*3�Se�	Ɵk~e������+ua�/k�(�#��=���+U�Qڍ�,�bR�';�t<����(�ݳ�3a�zd5��+�=W�h%("r9Ԓ����۫\}y����n��K�Ħ�34��j{��O%�]�����o����U��1�)vD;fo*cw��
��T�nW>Xe�������GX�����I�[�,2��I3����\p{�����I�5�,��u��n�H���Ɛy���՚��ڏ���\p�#[n9�t�[���Ȳ���7�۵|]�JI"cR�e�g  � ;���l�m�� �hZT:�L�R�����^�8!����C��!u�d�@R��II@P44PPP&�2WVQ RHPUC�BR4'$9)�8'��'0�HdM&Ha%
��JR� қH�j9�ԩJP�H�T#JR�@Ц�*�� (i�Uy��_����+�w���e��Y���jt�7ط�L쮤�Y��(\s7���G�]�7��MW~)0�:��C>��B���x�]�oφM[�p��S�9�B1c��o/xOz]tť!����:L������y뫯}S{ap3rR� �_�o��$�/D�F��m�/R�[�7C{�m�+z�*��������KꍺO>����l|-ϟf�Q|��Q�?y�� ����6�'�o^r�ھ4����	y]��9ȍ�JΝ������,ߵc"�kq�ߜ�R��t��&{��������9e�]�s���wFi�;�h)U�<�#uY�эԌyy�u�i�;�mS%wG��y���b�u������1�i�V�L�\�h� �6�Q�@������m���f�ǝzؽ|[�d_��V�E�uҿ2�ÒOOo���R3�CaÒ��^s͗)z-�:��}-�j��GN��<�Y�	�4��EP��;{��{u�I�Ó������w����T�~����Om�,��C��+jߦ�����G�:��թ6�M�N�\g{s�ʔV�y��x֞�%-폽 �w��3ՙ�^��ӳ�U�����i�݁��Ъdbox�u����I�z;s=�"��vy.�{�=��<�26l
��,IK�wG�>��2v��=M��S)�r��{���jy:�*-�̩fL�36^���3+���\�S70�����~2�����U�w�һ"���}Qݷ����@>�{�S%��9�pS�x��t�F}�|�b
n�,��IB��'�{i�f�r�y[�˰�F���[�v�RG��=5�_)����Gpse6===<e[�����ùgg7�M
9��aw��I岨>�e�Sޘ��ڝH�w�'#+�$�7ڼFE����e�:�z�����9X�t~�&�/�[�x._9��<�۽�����Bt�-l�<��u�.V|�+޺�63�1��f+c�tR�Oe��&����n���3y�w!Ͱ���I[3x�F�Wln���*���Gi�m��k�����}Z\�� z+�����g��L��}\����o�l[[�M�]��w��M�'�ʍmz���Vv3ZI�w�&�^�,J�P���=���c����w�{�wF�a��*��v�+Ѥ�&����C���5)�[���X����E�3�2��vs ���>*ނXuoE��S+�8���1�}&�!�в���Wz�ê�2�Tlzi�9�*�l�e�X����9\��afo���x"�`�2$@e���5�g�Е�ee��푵Ϋ�7����(��&0��Q!���OQ�r�y�Ms�G��7WI�"V��`y~n�9M(�2�����^�\���{���c/�S��n"|���O>2�z֟���I��5x`�ms��k�v�f�K��u�{g��}�'����է�+[������g{>z��F���5��$�����Ή�cT��y+�S$�^��Y�ӿC�&]�OE�sf�ޖ������i,�2|�U�z���73�V{��b�����-�!��g#�߮g�8�;�=ɺ���ʞ��n{>���Hꭧ�Gr��4���L��hw|FP�yr���Z�9���u/z�[�Yا'N�=�7n�WD���d���H�sf�����
 �wG�u���k]��	q�۞4���ͭ�j$e���ɏ7��T�׺�yٳV��Yb��[M�5����#c`���[�	���n�k"^��D���sh�����ٞ��y,[��7I3�Q�*^�ƞ��ou�~�l4�g���CMq���-�OK�[�9څ�.�����.&k�F?C�b����Κ"X]-��֦>��§�{Q�S�s����}!1vCKf��LgGf�7�0��R��J�PSy��_j�x����"+)l�4Ve��d�	��6�>Z��2B�k�9YQ�}�g��Dv�G�^p�zz4}���Q���u��]ͤ�\l��w:�:��_׊�{N. �{ܼ�'t��$(���.��(��B���5�|S��W�3Ckk�.������}�PR�����6(W���34_k{�X^�r=�+.o�**�G��'��͚�ێ�n��F�Ի�������ާĞ��*[��Y�b
�U�������ޓX����ǁ�X��F��5h:Vnci��⭝ټ���o�ӗ�^&v����:2:�Z���]{@)�( �?V��YK�-9�莻��qm�r���5×�W,%�,�ju��'���f���-�_L/y�lQI:?U�WO��'�R�V���3ĥ�۾N{(#+�xhf-�k��c���!���8��A�;ܨO���(v�-�A�R�~x-𺙤T펖y�]z����d�f{���>��9~���u��E��Q>�wC��^l�S���pB��N��w���y_zz�Ѿ���Og�o�F�m��n}]m���ؔ
�1>���r���6�&����#���ü��v��\6��܆]v�/�G|�۷^�	p(=Y��Ӈ0�ճNmmu-�	�2vp�d<wo��d
�-�>vY�ܒ�ҮZ�O�"Uˮ=i7ʹ�f��o۔k���
;T�ݡ�Z�^^��'��jc؟�=��Y�Q��^1E�=�g����796#��sj3]t��{�ez-Nƙ��ԟ=��N�tM���-�h{q�ݚzg0O���7�_R��*�m�y즽(�6�Ä�/�q	�N�WCk:��J�W]��n�8H�Y1հ�>����u��$w�r�zV�וW��A�"�\�[��f�OG��ed��\�=YW�o����s�����íc[��<S;����-t��׬��{A{r�<+%7d����hfSk��iΏ�:d�lk�<�D�Gwh�oSо�[�h�J]�j�[�ce�4g�藤�R�}5�C6�,3Y�h��P<~���.�u�Ժ^س����%���z��YϓJ^F���1�us�T�}���F6Ҹ�3]7QR�5VuЅ*�oH,���a�KwٮJ"�p���+2�}ʭ�1YX���U��rS�|C�ɷ��:y��)?���t�]j�q��L���M9��oԫT�B��;��W'm�1�8}���F�1�`SD�oF��<�´}�m�sNb���s���:�瞷�p}y'��k������y]��pG�����ֳ���Ri��W�1\�4V��dv�&j�^a��Wt��s���&�VWR
�k��Y�.��j�ү�+��͜R�u����Y|D�AjJ�P���emǎ��@n��f��:�o)����V �B����ՖrS�r��/~���5�U��@��h�AT#ap��n�����7b�8c/��I��j�`�Pg��g�]r�)j��K�9*�D��mv�]�NҔ��L�Z�-f;��d;�W���1ήЭ.�A��!��|7����׿:(�B�$fq޳���G@��r_�ޒ�5����Ut콪���]��]�|/:v�����&sӹ(I�S�m�3���<�F/�㴉w�y�2r�c�6��8D�w���ñZju��k+v�y�d�)���NL��!�7�#�}����            	y@�Q]A~�y0�����i�w)��;$�̋���������s���qC�K����5p��9�4<F��fs���jƍ,[���j���}1�7&��9j �q���gv��J��V�&��k���䢻�u�!���0[�iVl8����W+��td�]	ǖ:�}і���	,k�#��`[��,�b$)���q�W)�*�=����2e�Ǚ<ݨ8mG0l�J�x��٨"i�"t�,�K�13�k;}���W.�=��5�GU���6��SZ�u�s$rs+��L��.���Z�f���g7esC.fj�V�\��Ro�BZ�E���F��Vɦ�#k�-;:�����Y;��垨�W�\�p    ��fs̩C�B̔3���Ւ�*����@1)@sE SAG1�;�a@<� UD
Q����.čQ���
oM�R�doT���
P�*y��	�R�K@f�Hv�gs���o���Ӽ�~{���2j��r�7�J���z5p{��s��YW5�E���ն��S�ַ��;��}���?'軓��r{w��q?�;�z���'Jy�_��B�9������ٯ|ҹ��,]�6�~�ߺ3_�#ʢ��bе�>Yv=�z?��:r���>�î��(^�W���4g�z�֡ԟ�U_2[�٩��ȹ�92�.Y��z����g�����k�QK��{����mJKD�K�
�����'�ts�mR��a���q4eK��G�����6�����q.�Y�o�d�t*�X�P�H�}��uZ9�Xj�%�5�SXCBV�t�o
�X�w_�Ιv����[�2��ҵ� ��v��hq-Sw������
�~�*��N1�tT��c���o�\~�Ǜ��-"���h�fމF����e�{����α�Hڗn���o)�o�y�u՟�䯔���|;��BN{���'���D�G�ߖ����v�s]�L���ߢ�(~jĖOY����:S�R�Y3C��?��g�w�x��s�<�f�އZ�n<�K�9��g{;�{�П*�ٳ׵�?V��3�I����C;�#<�|>�9�p������ꪌ~�s�����͛2Q�	��o�L����h]Ce��ZA������'_��TF�_�e�̞��6WgV¶��)<�$H�X����`���������_}�Df�����+�-~Q�`d{�-幇?(+2�`C�w��bf�6׼�,T���%Wƅ��^+ �M�ԉ{F�R�š�[���*.9���̀�ޠj�xv5��
C#�]
C+�;���;�k�����Q����b���,O��{̈5��i��s_�y����Ԋ��yÈ1הoN�}��׾��O�5�\����M
Q:m��{��r�{��hK֓jؿ[⼊���G���X���͇p	dq�3[7<�ꏹ#/�@��E�hvlu}[���f�?T��߁�mf�!��7d;.�����r�].�1�6o-/���~V,��o�w�+kf�؉���{�Gn/E��5m��w�eD{��?kg'�Ү,��z:mK������{�%N*��C���������'�������w�r���\hL��}<3#��yQ{9�z��W�O�>�u3����Q�q�����������U}��"!_W�z_w�65��ƹ�z�Ѷװ���s����uζ��}��5�uoPs"Q�y)䇾���Pu	Cܻ�ir�W�p_d);�մ��ǯw�<q�\{�>u৛bw�=�m����`��c���>HPy y.u�B��4����o����~z��2�'R�NǸ'P:6É�یS�N��v��8�7��ԅ��C�{�Լ�k�s�|�s���.���f��~=ͯ-R开m�@K9�/�����i�Y����Z���/8,�k��Ti5�� <M9ܯ �V��)��_}HSŒ=Ǿ`�Hk0Cx�v8�:�Ѷ&�:�o1x������L����r��o��׺��|�%Խ���Hs�J�h�B�a
9�5�r����܅��$�η�|���������S���]�$w�a{���iSyh`�Shԅ qq��ܮ�yl��{і�s���c�:��Ӽ�Nc��^��C�];�\B�+�u�x���� �{��0�W�;����{�^q�y㮺�S��|d)s��/�lo�u/Rm�\�Hqs#�Xܣ�q�#�'y�Ju%��t��[{���Ϟ��HR&�Թ+��:���0;��}��qSQ�/R���p�G�=B���s��w�u��{�>A���B�!�C�ry����}�����}�n0O$u�ys"d��=�w��5���|w�^���9�2�qh��z������!{��=���:��m`�H���]��w�~��~u�Ԏ�����#�� �S�^���:�$)|��^��b=��lo����+yO{���{�޹�2 �O8�N5ȁpHd��ԧpy
��!B�q�I��!KԽ���rm��<��񶏍m���W~�/Ƶ~�8n��I;��{2��=��V�0f�Tg��x%�?NW��`�-���yi4	�-��m0zoA�]o�_%�~�㞼����P|o�WR�w�
9�]b�+�1�	��J�;���(^a��*k�_�xv�9�3��u�����/Q��[B��)�ܮFI�X�Xo�p�Bm�!�/P�=�P'>��w�u��������x^�|�}��`&��c��Mm��Rl{�o;Joy'0�+��y{��B�6���μ߯6ߏ|��|��^���i_dv���� �=�;5���p�)��ro�w��=�.8�.��7�z��B��I̾�K侽�Mo�B����B�8�c�N�z�P��qw��N���~���y�z�C�=�P�A�up��y/���B�y����|� Ѷ솳ew��%My�5o����>{מ��&�Ju��0�2d!�{/��>�B�"�vm��!�0ig[b����n��k�׻{�^x	���/�g�ym�2y!N���q�=J�&��Ծ\H�+�̏�*k��;�ݸ�~;��}�${�}�u!G����
f�:��5�2y/Ro�)ԾA���u!�/F�i^�!�6��m�8۾���M��}�=Jm���`�A�J�K���'����K���u������69���f�绽��̷��p�㨤�T�_w�9|�c�/xV~���x��v��+?�+���bR���h�5;6rF��Np�]'\v��Jr!��۞z�ξ ��/�| ���Wxߝ����{�!:�c1�)^!�7�P��y	����$w�fq������^u⧜g6�C�؇�>�w��;H�u�d�@� �N�6�;�{�ԯs�;�޻�~��s׽z���'��\A��C�]a�	��^c����Jw���������ԞK�q����v����]x.K�y�'Y�Jo)���+���8Շ�=�m�!�`z��N�y�HR>w��Ͼ�u���������ӜG�x���Cs|N�{�n�J�xC�7� �W��5"u%p��Pr��ǚ랸���8��=���qix���{��x�3X�����=���' �T�|<��n}�\�|�~��޽J��lR��u"f�irW�1i|���V��x�R�6����!�{��y Pm��������{���\�8�yGX���R{.�`r��.m���<Hh�N�v����T�Xq����o�Y�y�]v�=;�v�y6��\��)��$_%��W�{:š{� |���1��c���n{�7�n�ﾽ�7���۬�9����=�G����=�R��y/����.w����!z�7��]�����lx����s�ٶ��#��y.=e�ˀ�s'�xg�kv1�l?�/��U����N�o��RB&�a5�6�l�@��6��s��gY���;�n�����ҡ�>m�~���!A�^�#��*f�9��_ 8��Nx�y��:�!'�z���e�_. ]]q���u�|sߝ{Ǩ�!�x���6��63$
5�!�.��A䡶��RklG�;�c�:�:�c�<��1s���{�ˮ8�z��}%�W{Z�B�x��2�6�Ԇ� 9����C�]m�܅!��9��M�$�����\��~�ׇR��̇2;]��q
���'���d�'Py!�gr����6��B���|�����~9�z�L��y�S�vù��$z���^�{��z�*m�)Ԛ��;��x���k������^{�^{ף���z����^����oq#Լm�wԧ��s�\f�g����ڿI7�
�]6��:��g\Y(j�7���Ø����,oʾ���X�ڢ���"�=��R�}u�3s�#p�%�CI�(ݍ�Ҳ�S{p1���(��z�r��u�Z�\E�[������=蹱c]a�Ib8�?��ߧ�QE�,�9�N�"m�Z������s�w���[�q��w�Y�}w��|��PJ��ޏ�"*�0b���?�<��9�킽Z���>��k��nZ�:.�Gj�q��C릣:�-j{9�mMQ����p�2c�䛇	�לVN�c����՛�]�s����!�VՕ6uj<myԇZ���4���lF�M[����8��w��z���\F�яE��]T{P���z��l雭�,"���q�l��{�/֕��f���!,i�ma��<���z�Xw���sҗ�z�3Ǭ������{�����zL������ﳎ(�z���
�jn���L�.�)�=���a������{��/��a�Oo-P�L�z�Sx=k��"�펟~���PB�V���)@��(B�hB��)
ZJj���j");�<߿�Dl������F�F\G��L�9]��	��y�h�����y�Z�T]C3<���^��r]��|�
^�����)Muu+��j�O�<r����:F��$�i�Wq�`y�n��M�I5�m�/]��nۚ^�EZ�OB��O3`�oyy���}1�j�:��W�	�(��������/0#�����T��<ny�Q_�V5�Ki�[��5$ʼo�x�	)��MV9�/�	=/=����y�w<��_���n��|%�3�w]�2�Hz,Z|�#�
���4���\|+�YY�S2�q�[u:�6���v%*�\�CI�c�x�x��l,��W)RSyWÔ�jd�Ǘp��YL�^nϲ�
�v#|�v�*�St�B^�"���|w,V��b��w��2˵��5��VE�r���{@�Q���b���[��V��._r�/9�e�@�P�`�p��Mwk�W�B�}��>�{1��*��{��C�*H�a�Jnn���5����;�/��:�Y^����H�e� �(��]��@����+E9�^0��T3k���1nɇ$�
s�I�a͈܋J�n��M� �,v�s{��ќQ��Z4�9:Y���/UN��S��G(
Q..ׯ&�e
�ݪ���u~�ܟ���            �x���D����7�Mx��1��ע�K�Ive���ݣliP���J�)i�n$Y��C��2f�@n�,�@��ꇇ��)^�a�gAu�P�s��t1|��n]�8^��ru�Ȼ��N�	�h��w6<qV^�+?���fyǖw3�y�3$�+z��wW.�W�I���ʉ�oM�է{Q�3�d��o6Y�XnJ�Ae���v��L�HdK;4�d�9k%����0g]���i_���2Y)��q��re���Wsw�=�>�W��J/&u�zH�c�j[SN�ܜ�/��7%�J�[�Z�y�Bi�!���9�%<K��]�]M��D��������=��@�0L�W_YtE�Ƥf7��-)9�T�-]�\�p    ����?���ޟ{�Y�&FQe@5�>I�MFJĆ@䔭��Q���9d|I�-X�N�jSR��IHPjG'$�*" ����JiG%7�6�.J��:�B9% �R����*2
��j�C%r}��CyʁiR���F[�B4)M/~���q�||f���w���Ci��)��7V�rGRsw�#r�^ՙ�%fh�_�舏���Y����giL^�+g?���ls�߳�[{��_����{�ov�z�v�!V�널��m���7=N�����>OК�i��]~��ǅS;�ጸ�^��Ldvx�Z�1k��9�W;S��Q����������}�ϒ�K���o������s��
�[��y�ٱ���S�Ϭ�o�|�]��m���q=ֽ�Wg9~��I��n\h2y�&�L[T�,eǺe��K�<��/�FB���&k��k�~]A~��ޠ���pa�ԣ1�ԩ��l��[V�Mծ���U��r�D��g��ճ���ڏ���{z�{)�NվmX����}���ҎHSq��Ρ�C�i�8����f����W��Ӛq˕Ư]nO��`ҿn�����M۷�\��@��LɼG5>U�3ڒ�SR��	�Q1�U��nUE�����"h�1_�e�$5��SU�������}Dt.�J�+>�rq�`$��{����놹���^����M�kk�5Zv�ߵl_����;/��lZ',[�*��wdoM�m��t����A{�;�1Q�v����z�і3�f #5=_����D9��K9�#�tl#��[��Y�j�fd��1��壘vs2i.��o|���_%��˝\�P<�S���r�J���4�o����W�|��{����#�;�����k�������g>�}�Y�����f���*}���CU;-�z2}E��;HK����}���� =B���w�쬬�A�����h��?6��`��
uר+��`�N��N��n���U{V��ߚ��S}�ņkÓ�SN�u�Mݱdh�	�t�|�߫hw�����d��G�^�g|�md^m�g��`��d��aL�Z��W���Y�M��]y���\���;�rC���c�p��g��}msګ>�����1��s��v����R^�=�+���c���Q�U��K8����+ߔ��޳�f�+������>��6��ܯ�?3��o#J��T�U��݋�DZ��b�W�̸��R�����4��v���]�+t׽��x�b�R�%j��d�r߈�~�S�&�;�^������o���}���wج������Z��\�hu�3H�<#��N��$�1��`�0���!Y"������g�{�hL�6��O�D�Ȩ�Q9�۝���5lFr�U�{)Tʙ!�%SwI��=Ǟ{y���;���U���鎋\ʄ����%�{�\�q�|e��&��yu�V�B����z�N҃l$�Q:���a���c]1(v9�S�X��2�{�8��#���}���ՙg&�(�����^��`�ge��{�̷V%��*��6����1ldW��I.ֵS1uc+2�7+}���ó(�<�o%p��J��@�&�S������^DHu��f���[�E���eܙ	��W�1Z^�m��>�2��Z�+��yi����yVU\貵K���\�+��5�Hy���h�
�g|[�{�u�9��A\ѵWq����s�_����S+��S��ja4�[�ٵ�Y�vf�v2�=��kKf��U�q��RQK��5������6e�Ŋ�vFL�wyħP��N�d;�p��=���x,�},���}_W�W.�=�S�X�_��/�V{�颟%��@ݤ�bM��k�>���ב�B;���sĝ{���I?"1ĵ�	�qm(̋%��*޴cÓt7'��^�˪+ց6�x�]���jf��q}�̇~�]���j�'��ԹOh���6��2�i1�s��e'/�&�)X���7�CN�籪/+VjN����M�ï���V�����<;�O	ʦ��ָ
��[�W�ӹg�]��4���+���^����o+>h�<���4U�N�V�m�h��;V��z�c�����	�%�t�%�'�r˕���޶�}�W��k��x�}�ۏ�~tts���ܞ��7>I�Y1���9�F�ѫb�g���i��ɷ�g��.s_\=5'����<�{K=�����������h�W�y�o[7ϏKُF�9[w�k�:&m>![,֒F�g�T�*��ݢvn,5z�yso���r�>B������U��؂۽ؼ�O����-9hRuՊ�犣D�X�������{t�_ӭ�.�L�:����yV��y�N����v�T�үjY+�(]y�i���zҚ��o�/�+����24؊T�'+D���XH⚱ou��ʊ��n�{�)�x�jn"U�$bԈ���yJyj�����}�}�U���=��p��D�[ut��D:>H�km\�,��$�8#]�y�MeVQvT;R���uc��:�s
�.���=���\)${�w�b���s�\�Q����׶$��[yf�<�Dޭ�lz�W��]0��k�S��g��2�W�"̨�{��̅���k���q���B6�H���v/�����\T뽴�f��.<�u��5���Ν�:UK���^Q��TH�M�u��u���}��_���f�����:�-b�0�Ғ<��]��7vN��7���`��L22Z�eGV33MYj9����iJ�ϲB��̳�ţ�gd쩪>ع^@��k�O��W�UF�s����7�+��y
?z)]�l��Ɨ���4���t=����E�zZmz_�{}���*����ו{ݎ�����ss3��Ոܛ�z�hқ�/,���t�����:}���f����c}��De��N)�{w�j���l�n���$��#:�;��4���ia�E"1�L�i[�|�]^��x�ǠRERU}��6'���V;Ց�8���G�n�6߽�:�yv6<�������SiU�/_�;�v\�L
y����4mg��)k�Ot��rX�s
� x�����r�4�S�0N�Qzx�GP+�p#ܻ����o7��}�#[��3IM��U:.�n?�-�==�Ϝ�u�;G5b��#�oޢ�{���Y�-�5�zs�@��@_*��Կt_ן�C�g�M׉[v��P�/0�?t��-��0�^�N_���wR*'���j�|ޞG[��]�~��
��c-{�|bMbo�i����W�B��'�c�n1��@�;ѯug����QڙeD[S�K�iXq�o���W���-�r6r�h#�!�������/[�Q�L��^v�������n�����ټ���Ѿ�Ӷ\j�U{���F(7��iBc�b��Ƭ` 4����/�IIo�q�t�	�m�������;�/yr�7��j�ls�ȍ>�d	[d��K�70�����m��D	ܑ�#8T��QГ6�w[��u���ݬf**akht�7�뀞���f�XX!�7�������͠Gm�w�U؀g&��L�v3SI����k�����s��ִ�v`�y)���H�V��G�|R|4fì��Q���}��o5v�ӗ$�3/��,��-Ec��L�]�0YBA�x�G�C��p����`��*�&�6r����.�Mct֢��kN��-�3�z���ۉ�D�q�S� r:wkwē(��L��J�,0���t#[�66��O*舍𛺠�"��Ȥ�o������3V���            ��c����#r�1&]ֵŨw�	�=@�t�Z1�VWf"I����lޮF��uz)m�;���Ly#�8�Ь��\�D�0�b�/�N��8z�:H����8h3�����Z�+1WrזpMз��ތXA���fn(�oѹz��ҙ:�(�+(��n�𙏃5����|-i;\p���Ŕ:�:��/Q�էF�|���C�lOPp��0i��đ;O��S�' lY�/����-GG4�A)i�.�*�xFmh��(�W�+���p#E�^� �a�ˁ�kW:��Ֆ����E��}u���"�X��r�1s��v��r	�i�u�t��*��ɮ�*�x������"ي��.�j�2��  H��iSh2@�)h�B��rJB��w�P��HR{d>���e�`LP�<ɒ����Z��!<�Z ��j�������lƔ�І�AIUHq.KT4�E D;��4[�KKAQ�[@dS:��}�\�_t�ev⻍���M�{������\�_,ؚ΋�Y�+�_���>���6V�T����&���ϔr���{��|��p?9®n���o��WN��^�{��hZ/KYSe��F��Yl�7����y4dzH����j���Z�rZ�iq�T	彝<�3�PL�PR���Np�SXU�ż���b�g=��)���z�I�����~YӳW�f$7��w��E��7�y�J{��`���gӽ��>�*Uc�̵���㵣]�I�O�VMR���.�ݏ�=�2_���ށj6��}{~�g���Q�l���4��`���l>�\y���xN���IH=DVe �P��3���Ña7���ڻV7%�������I�����q'��
)�v�{�yu�E���t���]d���B����.���=����ҍ�->������4��i��oY^���zY:k��V�|���е�{x]6�@���aMs��ut��0��/$גn�O)m7�A��5{e��K��琮��"&��ߵ$1ΰ��l�ɥ�C7��l������QI��d��V��i�1�E_�X�}���o#|��=;ϣ��i���z6��m^��7�	�F�yA��ϯM<IW��5�R��IE�p��7�qe����4�[ӽ�S�S�4����g;���*�U����S�,��}x6�kc�d-�����:��ͼ������u�ɦ3Wg¡��/�;�{=*�:����^}�xַֽѿ_#�2y�/}�g&��������(�ٿD,��d�&��Ε�D͎�,�ϐ�kA#���vI����˓�i��N:ÍX��s���|�ϝ]z*��Ϯ	f{�&�k۔��[$���O.����O*�1q���)"3eA}��#�,��:�'6½�{�&Br�z�i��Q:�>ʮ�xm�8y�M�z�����;M�]�q�Oɜ�¦Ĺ�r�p�'j-�k0q�G�t}�GX��#ھ�F��f�c(�j�rT�?�UU����|�#ט�Ti[Y�2��#M���)v�����R�u���MTa�V�L:7���1�~��9�F���Ds��S�;S��]W�s�uv#1%�Nc�ůzy�~Y��u	���V�+@�{Ϳ/v��V���СU���Քz��/M[3]����,��pK����L�z(ǇdC�[�nH�S�tOk���gw�{w�g��g���mKB��m^�r}���W<ixf�j��蘞��${-]Q��m���Wp-Mt4�2м�x=��1F���X�Uj���~u�~6�H�g!����R���kft`�<]!��?G�}��OxC^�]��#Toz㛚�mb������mz��vI�oFC�s�&fǛ��/��m���ދ�md;��d�bcA^܉y�=~��7�uԙ��1l~T����ُ�]�Nk�g�L27��
+=�وL3'a<��Nt�чX��

�n�����O�����vz��D�0�ޗl�ѫ�õ���S��+��kSqk��o6�w7����W~�&cڴ���ʴ�L�O7n`�shۈ��0?y��^�<�߭RIQ��E(7�/$���F�v���H�Գt���`��9c�P̓��S��9�]��K���}�,��꯾����Է�*~���Xx�Q,�/*�����N�5��9�m�����c�c�?o���k'��crn�Ww�<�8f��Z3��Ȅ��	�]���O= ���>:Sy\�
��K���,�}����;���ͨ��Q�����aX�<�Oo+$\�(r����jdvE�.�yĤ��X���s��ҡX�ץ2)l'�OJ�s�xv3~J�⅕8�Z�Eҁ3a�G1���9���Bڬ>#{�r���wز����ok[�\�B+X��k��/;yqZ7/d#X���
�O���%!�����W���9�'ns���_W��s�w�s���wc��#?j��=�i{So.tz�����U�z���l�\j[��Dޛxע�������n��C3�;��kyٙ��~uH�<�3�����k�:�������WVx��}9G\ML�Ⴔ�8_Ā�	�&��m�C��VT�w�׽y��*�����I��*Wz
k!��LU��w5v�|�5�?Es닊��)�d���pX��k|��=��t˯b�`�8i��a�nS0k��io{ܺ���ᆖ�EXwu�
�<�8n�+b��Mڐ_*�窌�x+F�}��ƸE����L�V�\¼ƀ��٫"o'��s]*<�5]۽���r�FF�D{����y�~w�zm�]����3�w��Ǎh�M&��~}�Ͱp�|,���P�U[��0v�X+�� �I�{���������*��dX4~�fz��
9났R��<�
�{���������X�\i���3�p�=I[��g��|d,AcU��y`z�4!+ �
�dg������jq�0���J�;�f+Ǡ�<�1�O1�Y�y�xk��z}�}~Ƽ�&R7W޿z��}�Öd�ҰA��8��B6GR��X��l?g��K7�|��y����4彺���cBb�Ml'�t��^�M���Wz72�f�h�#�p�\��F�`�
c���L�!���9q+�Z�mU��I�:�]:
W�a�@���¤��ݪ�Х"85PC{�s��:ً��d;�r{����iOy�^2�m�_��\ϑʆ�f
�g;!��F�x�7��t�k�a"��A�����ٮ��ɗ=~���#�#�>e?�xk��^���3[^*.Q^�s|��6����" �0y��b�`ax�����N�%¹��r�]���+�,�
?f�Gn).< �qw��N�/���7���o�(A�� �Σ4�=����t%�����F��h�c�&�y�0�A��LX�f����l�����WK��/,���J]��0:� Ū�M�u�l�g���o�Ozip�Uz/��d��W��D�A�8��N����^pO�������L�N��c��k��4�+��_��k5��~�4����x(E+Yu»iǲ>��|�9W+�D�WÔA�U���P�.���R�n<�����Q�D�:�+���U՟�x�B��(Ֆ���v�����.$y��k�|+�0�VU��®���I��:2�d畂�pr�
z�G�p���w�	4�Rw�vo���+�]] 6z�POz�L�^˯-�����/����k~���B��F�]Ҽ�B�A�r��y�'�Q�W�V��*;`a�\
�UăWu����a������+��n�"��B�$wMx0(!<P�o´eZ�;UϽ��cܞ�
j���*�n]J��*I~&�=���rn�\it�u��,]�c�+Q4"ǭ��w}7��7*ǩCF�a�Z~5/±hׯ�+�8V���ؼk�6h�(0Sqq�f�G%��QF��]K�Ț��w�q����yp#�>�v�1*}��m�yp���rn��-�e���`�W`D�ϧ�����X��/2�&�J��Ӭk����z��ʊ�^�ƼM��FH���Yz���@��t�VsbH6P߸c�X;O\�X��=���(sZB3,첝�b��n��R��r�a�(�^�}�����Ɠ��l}���+�bV���{n��+������u0.�+jml�an"�1��epT�6�Jc-8�mX �9
w�;�[�������YtI`�]ƥjJ�D�SF���.ɣ�Ú��f>�X�-7���Ζ�wT�+�e����1V���;7s�����2%���"gA�7���h�D'��tBy���E�x������gdI�            (P�����F/l��3� �����9s���5:���&�*��Y���s�S�"�駨Ek���Ps8Jz�Bͧ:��nft�t\ϴvu�t��͎Z�73c��ӷa���}�y���ٕ�h�85�yw,�e��)٫�R}����>�w�N��M]�D��i�"O^�m=�Mޮr�#�nvӤ3m���#�-�Hi
��8ustof�h�*�z
�@Ĭ�m��m� �s�a��ǘ��13���a�xs*Xs�ҎQN�nB���B>��)j��Xe�B=�N1lβK����auNT���I�3"��`���N(�S�GY�Ru�YH^�5��t^[�$��T�����2M�gVS{� � A3�c���PГ#̙-�4�Y��oeIH�P5�k
*�ix�))�(Jh�P�TPR�H�RQ���&�u�R�\Jq�F��b�"���"����MMXUEM10E5�D�I��m>�P������� ����#dr�-�
mC9��r��N��Ӛ+�ɗ?u\�g��{�?uv�h�FѬ�|��x��x�Pz�ǧj���V���X�R�щEK��~�T�

����&g�<�8� X>7�����e�i�I�C+��f�k�`��v��8�	Ŋ5����],
��r�����A7�yaC�����~��*�Lo�.�5@��~H]fC�
~~�j'SW>��8)]��;�u㄄��B�<)����/�;���:��zq����L@�o��4v\��ׂ�r�����u�@�tX�|�<,pt�񦏆���g��;�f#F��NWL�Bv]+�-�.B�
on��>����ϟT��3P�p �@��v>(eP�3}ԭg�;��bv�pw��K���������ȱ�&�~c@�\Q�w��+�{��T�3;�m��|>`�x�&r�b¬�6Й#��>���y��[��ѳ��r�4���SJF�k��&��μm��n�r%T��Ϯ.��C���;! +ٱ�Gމy����s0`��f
5�P��n�5.s%x?G�=.��l�x���1�EXvi������y�|�ZLb��+ޭU>��d�XH�ZD>o�T��G���j��@�<4��W�P�U[��N�Új�:����m���� �WC���l�(U�4| �k�,�4y���k��sRG�����X��q�;�]k;�^�k]Hz^L��B�i��0f�L��>������+��{׋�NsR��>�~��k�P����O�n��5b
�����w��`�ߕ��`9|U��++������X����5�^�0�7���a�����wT��<�<g.��u)I]�䶢w�!{��~�И7�?Vu��.�����޺�Є�f�=��Ş��0��Ǉ�K�|��f�8M&P�X�Z��Қ�ݑO6�};.�+�uqt%�ݠ�4U�{���ý���MS���o��q�?]p�8Z.+�'���Y��_x�w���Lz��Tb���=�xV�
_��u׍U�`�]����x���+��E�ǆq�}lua��;��ݥ�5�)���VBG��/�h�b�y���ztރ������^);�	�R������ �|#�xy�b�t �],��+ �ԋ���eײ�ثF
�k��H1.fAu��թO����}h��6)�a�LWI��P�v�=2���[�E2Fc��a��jNGA�zvf*�Y��j�Z�aX��##��Z�"nܮܚ�Tj�3˦���N���d-�V�;��8��꣘Ӟ�~�x���Ƴ��72���t`@��5�
�O`K}�&�S7'x����;U�K��^��h�y�T��(0i�gGj���"
�u�[C����W޺l�K
�5�r�+�@�z�y��Px끀=�~�@�iB�����كf-����H�ڨǕ�诹��=��F�%�
�+nU�2G�����O�Fz~�
��
5�3�s�I�@�j������6�[���]Ѻ�R�VVV�ex��4ǅ`c������w�_iYM��<�c=�������?l6��)~�k�_����%�$�hz��< `xם�iFP?
�� �^5��ãx�)�==*�\j+���P�ĄMp�2�����'}�a"��{y;ד�\�+�i����w;ynE��m�9����Մ>FJN��b������ѫ��'ɋ�*��j9�i�>�ӒO=�YB��P�����.�&zؙ�߅o��2��7�ߋ�����~�uS>��D�
� _�3���\�WC�ϒO���ז���+�VPxX���������3�Ox�Ww\%k�`iܗ�WQ5�0L4����7���y�=C�a"�)Sp�i�	g�����!��3u�~�vzGZ:��;�UZ@��]aЌ5�N9�S�/G���(y�7ky���{�l�n�Vaz������*��C���'��#|Ξ����Ӟ}+�E��?bu�G�i�2��c[ՠ�׼��7]!�T�Z��b�è�b^�w��~�ކ)�b��!�Ы��>t��fwU���:cU{Z�SxϦL}a��9�b�uĂ8tÄ��}Q��N�v�u���7��kQ0�}Q� �4w�<�z8f�}�ҕp��Ug��{���:�4o���������!���,��gI�)��z0a({��>t0x!�|��a�o���~9ƀ�NWU��.� ��f݌��]�;$qs��j���W���t�� �S8M(HB.���ħ��vX�+4׬�C9̪�x0i]�t� @�{Ucȅ�.�J5�ݟ�i��˯eu�U�,�<$:-|i��P3d·��p����.�m�]q���[\i���Xr��5���Z��z5�|j2@G�!����4�B
�B\��X������_�+x�r�
9D��]+5�B/��y�R�~#	�"p2� ��?:W��x ]׽ĭ[���!Q��]Tvk�{@E���e^�!�S���G;;��W�lZV��1֬�)�����`Ԥ�Ay3^��q�5�7��UQ�zG<�d����;���ZɆ�+��{�
��t���&�HR���y�����0�
��F�6�ϐG{�g�v�?��3Oևٶ�`�lAދ������G���#��x�œP`���x��`�������d=3MP��lW�G�}p?�ZP�V׆е�m���n�#��b�x��t*�9�	���ؠ�t|���]��wK��t�uCK���E��(��'�=X:?l�Q�K�y��`_KBqcνu­��:+���P���cK�;�ExAXĚ�uQ��v��'��/��=�Og������{�k�Y�Kj��	<}xh�\�@���� �}^���@����2���wN�%�c��՝G������я�RW�Ǡj[Wi��iw5�ec̹8k�
뛔����V�"r�:s�|s<�'�U��P��dr$k(1�h�j+��k�m�5�s�(�I�%��~�0X#�5-L��@��2`�٬�ҽ�M�^l�,���N�RS��K���X��du�F�{�^m��KM1��Th���uu�=��F�}�o��lQ����3�Y��&�|D:j ;�E&��b~~����{o,�i��~4���4_{*�0=���l�ػ���<�*Ǹ��,d;�F��M�+��CEI{5���o��hׄ���Wu�΃I��	��zG���;��]e��t��4j�%�
�+V��{}i(��mp�)K���B��Z�_m�
�e��j����=��;���g0�q�^ڬ�4BcOq���iӻ��m���7����^;��I/,�b*�=�hg�b��Y��n[`�����G�y4���D��&��<{�u�,���r�G�\4EV����c�~���^�v �+)z�� =��������]yYaP£ٳ����r�x+�^D֔e+��Ӹ
��N��p�f���o��j���Wu�������p��;^�ٶ���fl�&Mg|������WZM���W�����[���6"��n6�WTmٶ��]��qގ��Z��Ɗ7*��s=5u�/|כ�~�D�eiB��y\< c����|��f�!ڢ~��ۻ��Q�V��k�
��]���0���\���V��U�"�-V�~���ٓɽ��Q������%�?��c٤
@����R���t��ߥ&�W���	]�r����!��s��1v?rᩨ���^П���G�r}ci�K�P�^�*c��tUݢ�_r�n9��S���~����˭����D��ׄ2�4��s�!�y�~e����G¯�~�^ƣo���4�~��_��P�¥�C�����]hL��AVֵ�b�?:�һ'.}=� ��ELS���֜$ �:=/�!�.����{�>X7�4���>�xV�A3-9;}W���� s��ɍ����� h����~h��Ҟ{�{�]oR�C�_�D��d�5t�eҼ� ��Oj����a5.ʬ�^�le
�X�d��	�){�D�u/;���pd�o�:�.�a�8��)k;#`��iv���z��]M�IP�i�9��<$:.b���e~O��ء�t�7��H�Jh ����)B*��Y�+�'%fݾ7ڰGf��ń��KnE/�����i3٤����s&�n���<��JA��&33��\�"�	��H�]]����Z��m�z�{k2���fe�2��a$�y,U=e��u%u_���ܬ��k�u��'
r
WQ�N�N���h麟7�2[:�qK{J"u�eKƲ�6�.�nL��:<�rnq��S9�MZc�e��K��+��������#8u�*6dά8-�,��g�,E@����x�hm�Z)���;3ᦅ�Y{�c�Q�SN�@ܔ���&��<���X��ǩЮ�����8���6�5�w�pp�"�ט�8�QMn�[C�$���N�5J�*a�f���F��u&�`            
.�Y㦼+�����wR�
�"�T�*��M��v����Xv���V:�����uQ�W��9��\��f��d�+�=��Mmi9:TՖYP�Nr\�]�\;#%�O{�T��G���@/�2]�|��b�r�{�y�x)@"�^��pg�r�9����}mgY�,f+�,����|�L+9Je��aQu��knR|���7E�򺳵J5�ɕ�1e,�M�`�����.�0�M��0wS�W����ͩ]h����h(�jB$��*�:��ޠ�7�:�3jJ�8��r��9���wD��r抅S[�۝Zl�P�pu1�/���S���7�+rTb��=��޷3�2Y(���m�W�   ����{�D��fMSEQIUL��P�Q���URy9!AE QNӑAE44��+�Cy�7��X�Z��	��V�92Y������Y��QM�9ƳV����jM���FeE���;˯�qϾ����]���6
2g���Y;�T3/Z�˵;�M����Jc
?��k�����xg U��z�m��V`��Pxi��sqg��T^�[�F���5���B�¼a٧z8/]`@P��o��#����������\<(�j�Y��Li���Ò]ʹ4ϑB��@A�"��Mw+��L*�י�=��� y�z�ea�@�A��i� L�,4Ὰ�h�}ɜ�>S}�RB�r��7U8�FCN������H_���z����1���c���W��!��t>�Yl,�!؜��G���U�;L�
�}��
���փ�ix��y��A]�ޏq��HA�|N
�үAϽu|`~5�l�#�|�e������?&|>6`��K9�
Z�lC�/��0�t�*�`@�N��Q�=��G�ϭ��]ҫj�v�v[��VV�9y��E��殴�nBo^=�3q5Y�rz�N��?�F>^���E~^��Diq^ۯ���AC�:�-��i~~���.�0�����=�h�V���<�].>������z>�Lm��]mS0zu�W���JR);59nK��3��^R�Y�5���(�~����h��b��۪6>���>>޲:6>Ȯ�|k����i�`Q��k���uh��b
��R �y߃&a�(>�-�o{͵LW��f��i�K�H1Z�s W i=`+܉x��6���8J��
��VҢ��t�!��Ӹ���~�����x�~&���'��������O�z��^��D
��dU��B٨/�!�9�>�eGI���B�Y-�y�/7�{3�nfo^���,ƫ��J�����S`&s˵0���{l�&۰���NX���h�;)�Q�
~���9瀁�h~TC�h2箎x��H�����˫پk��{v��9�X<00L,���76�_j��C.9��b���V�V�_�k��Y,x}��d���*�}#U0�.�2���H�4�]{�N��1�+�&���{#~Da�)�;���<�/ S�0�u��p]`�3����0]/q �ׅx� 
��Z�u��n�b����H���[D���U��L�@̺�]���}����mo�����i�μ�#�%�[5��+�~2��q ��
�v���<������V����Hs,R�vE�d�������S�gg���w��
�m�)���t�eرH��@U���(���Fe�ِP�vۮޏ:��j���L7��&�2����&g^۽IX�I3;�N��1���w�b��A7��6�ɓ�	�}�|�)����朞���x�X��]E��h�b�{��z���z<i��mLz��]:�+޹�U���ؙ�rx2M��tsҘ��{8�U�]��D�6�fq�.�q��aN���wc@҅1	B��*�Qxt#�N�߮��g !���D����<< @3�q,�5 f�%��;u�4�����X���!2��G������vEw�i�hya{��y����&��py��Ƙ5��@��Z�x�~z����у��θ*�c��u�cV�C>�+]���/�_r^@G@j�C�P�7�Ld,�C�蟛�Ѷ��^�b����^�J=p^�(:���~�^�{F�	�Z��+��M�2�d��ʌ��B��'�ŞCu�Ͱ�a&U�PD�y0}��@�d�S{v�sX�,��UFrjO;�W������5�s�4h	��mۜm���Y����4nOk�)��Z`T)�0*�A��~�(b�o���~������
ݮ�6t!�]V��0U�ٓ� 0��8����<Lh�53��n�וa��V<;+���¬���<��>"�H� \=�1�t�_��k;�WƘ����x��n��5�~0�Ga�x��Ш0�Hhh�=;քSgy������F�f����,d�8������]��o���f�}�����
�D Sx~�ʾv��^�����o=�v���V�j�ж|4/_P�(Uֻ0������YO��J:=�5y��DWn�݆��;�������_q���щ�e�����Kxd�J:rY'&ĵʇU����[��B>�Xؼ	�ޘĽ��pW"h�$�Iw5�_.�6C�~�1�o.'߻�����i�Py^���kn�ƫ9X	�8zO]I��M��p��
5�[��w�m�i]x1Q��{Q���F�B�oüpV���*��Ѿ���SMc�w�}DDP�w��`�φP�5�ՁJ��mf�����{��ǩ႓� ���].*m׆qa�?v��}F:���J:�ʺ�~:@Z|0p�]Q㣂g�l�{��l�(�5��Mx!��]�u�p�y����tzԾ��j��i�k�ye��
�+� P�̀��p��	
�Ȼ.�l>���a�Q#���p��?Di��e��+�_zt��Q")uu
�p؂��\ y߃&W��х�Y�>�Lܡ�o���;s49�L�a��Mve�η�r>�|�ny���=8
��H�r�B�+h����noA�oy������}@X����H��.�$V�,S́Z��о��O)�Â����<8>7Zj
�t�?.�Jc��JnM��M���^M�K�l����CWg���p�ʾmޥt�{����Nm���k4�(c5�x����.����i�d�I#wPW �:� r���z�u���*��H��lCw2zE��kxי�~�\�2� ��+�^��z�|�漂�a��^�B����b�Y(AUy�� G��7��u*�q�j�h��듯�P�L1��4�.���B�����5C�)�R8"�0V���^?_5�h��vw�����^D��i
���=������Y�a��e�[�$��}���Xi
��yS��,6��ǫ��50��/x.;��i�����+:���S��!���Eeڒ����n~���I<��i�?es�IAt]�˺�*��bqr�o�F�ϟ]1�z;��9�]q_����"�cr��y�b��uCv�+���h�����j�b���S��w�����Ⴐa5�,S���Iӻ,�+jxI~�kҮ��|Mzղ`�>ƟZ a.�.��Xܜ�X�C¼���	�MM�OƊ��K��働9x�����]��Z<j�g*�y�]]&k�O�������U�Q�t�xY<9XA�}�z	�S��-����d(i�+�E�(V�,�W^M^<�{�1�s�?��0<60W�cG�O��(T��E
�T6�zv���!MA0,mNJwX���sX���B\Z��*Ķ��rfdCd5|������x껻^ ^�i��_��Ûm�^O�~��U�ֈ~����L�,7 ���s��{��Tj]KBɭ�hU�Ul��Xk�'�KTC���X�>�ތ��>  xѽ�C!����o�K�����h��4��n�3ń�C���èk���w�CE!]�Y�_��t�5l�tU��>�;�2����!+H��E*�l}�P�d�C{1�x�{��8�)�؃�:�~�4G��r�Ш)�¬�����w�W���ɭE}.Y*J�{_i�Ryw�t�1��=
�60 �1��]@k��z|���������
�=���)*�i� ��!;<2�h�~Q�ou`� �a�`�I"�����.�F�j���s2��w�Wu0K�<�M�P/�i'/8��l�Tz�������S���i�P�˝;7�Ugw���4V�?}�a
p�
�@��d I�q���)�V�j��;p&��{pY�~YW�j??<��]讔wF�ᬡL[$wZC|``	��by�5�5'�M"��_�q_�w�~���M�`���ד�+��澂��87+Ç��筎,5��z�cboپ��掏
��E`}s�xL�Ț�b��ފ'�$5��t��;׌�Yd�5��|i������xk���eR7W���\�,W�f)���B�o���Wq�I� Q���,=:��
਻��\i��<����@�j�{�R��Z+���+p���Ft�>�����a-�C/"��_��['D�Ա�գ���l�fd��NVlA݋�0�(���U� ��/�ugof9p��¹��\0�E,��+U˾.f�{l5BzZ�#�Z�pT��͗+u�m)U��2�f�^n���':nٻwc(w<�J̋�v/�<�b�$㈮2���H 
w�`4����3������x�Vd�*u�;�R��Y���E��绽*�7pٿ�����f-�Y빺ҹ�̡k 	�v�EO�k��l�6�	�q������z'X���eZ�d��3�an�*���q�-#}&A��*��3(I9Ö��B��Ǽqu�:PuA!t�q�{AV�2w��v�c_WJky
2�ͻb`׶,�n\IE�[��J}K>�%�W�jJ��             �M!�3�W��[IH�.-�F	�n>-��`X�=١䝽�V���9}sj��M�X�E#.B�}67���D���\��4�[��3u��]�>��S7�oePn.e*�@t'��Y����ݝO��Yb��Į����IR�k����`*��l��7�U��jܣv�&�����7ه�SA �=��b2�guĤY��;���е��"V���l-����%&�ƅ�%�M1���4Xi�x�e<�w.��{�P�Vܺ��B�Ι�0vF���7��]A.�XyvO�M�w��.����%I3��e�s�"��"���;��p��NR�����a5�:�fsר����S�\�9�ԩ|�����ܐ���T�:� �7n�P   ^���{��D�}똟DW���F7��9d���4Pjrm��m٘�N�v�8QS11�m��2�j֦�+,����j2��6��Y���ffFU�;Z6�}aF����X����ʨhi�Z֔�|�k1x�u����F����q����8��5[�h�.A�٠5PRw���.���^-�0;��ڤT���]E'�u�����9ta��������w���у��*+]dʿ=:��#����(ҳ�5���f��
��B� iv�nWK�!����|$Fm�y��ތs��F�"�Y^4Ś?�],��V�E�}���Mh����0X!
g�U� ����Wؤnl��3@L!�z�S�v)+Y��������w�b���X���Le+�ƕ[t����ʸo�׽G��Y�C|~�Bg��B�\��M����U׽v+ �c*��^�T�k���|h��N�t�:uneW��< �~B��^�P�v���K�`�)��<رQ�������~�� A��d׷}�,$�^WV��;헛�@Y������j�ǹE��5�Y{�­�F�Ȼ�YYz�ˮ�뱻}8�\����b��%[�uB�T뚟��㘣���1�����޺ˮ�B�K��+��(HvS�����ӫ�~�Q��Ge�1RV���F���
��(��3�:aТ/�]T6]@���JP��E�~��=�2�A~C��]x�$��Q��X�wMA�Yײg�������A������"�,��Mu�Br�N��zy�Fg�1�Z5N�g;� .2��;9�ԍv����O7bQ4�6S�C�v�qb��P�&�O�Q^[��π��̱�0V&��[A��$p�po��銥K�j=���8r�}�X���T���]LUf���BPOR���i����Zɡ�χ���o���#NK���}[�Jrle`�_\	�NY���㘺
J�)�U��<�3��RՐ,���fV˧ts������]���R�US�aW�
����;�6�c}~�Px�
��
� �9WI�c��fb����0��&���LùY�(�>��ѣ�X��ve�:I5���d AC�ۤ.) ��Z��ѯ�Rܻ� \�)�Կ����
���P��ǏO�aK���;(I���d�_��c5���O� 1\9���s�`����
����a�Z��RȮ�v0���y=i6�2�`���.�xm�Pѽ�Bo�-\��ޏ��u%�^v����`U^, ��0CEa�[ݽ<��A�K��xU�Uƍ��&�c�z�E�ޝ�?eՈ κ�U��]�uX)���hb!��H�k�\8��#��2��Z�Cwm�++���^��C��q�a;N�<�Q*����dʹ�s��:�\g'�v�Y���HC����{���{��:)�#�����_mՏ9˪��y�H�6���O�V�<0�ٕS>�}u�?mt�J�ۃ�6t�Ǽ΄>Y����>c��4�_��Y���Ф���lh����EA��I�Z ~����+�����y����Wu\�a
p�dD�:�b��+t��M�3UÙjV�����A���g̓t�fy��K����x�ټ5^j�>5��< ��p��v>O�+��"��P��ا�������/e�<�?i��8�@p�=�nVR8ވ�~���{dWK��t㞓�܉ �| �2��_C:��u�r�(��`��lV�����o�b6T�2`����D(�Ѫ.)AѥY�q������]�:��v�Q¦���"v��`u��.��	,1�2F��3}��b����^Q�(��	��Xd�^U�4�D݌���{�{S
����5���F��b���E���^�^D
�`�ح�����>��&�xpa�k�oD��I�����D\���j��}G��b�e�ϲ7o|�'�H�%��4�51^f��exA�K�(�����\3O��e�K.��
�vhYD�%��,P�F���,z{�}��k?j$j$(i�C�����n����n�ƣ�ω����P�`��ȫ  =b�sO����&�] ��Éژ�a9ꘟ/Gz�/��z�3�������̍7���j�E_��!�}g��z�34�)\�oڼn�Q�oX:��;���Y�fe�',� }�(�Ή�Z���罘�7��E���N�2�� �����DكCO|z7߹��Ң����]��{�o��	~�()㕍��͂2��)�$!|@��<��Z/�~��w��Ǟ���r<t�����4W�1�|���*+�W��s��F�=���Nأ[�F�ƍu��+���	C�8�6,�>�������Ӄ��EЧb6��*����?vyy�����}�7 ��a�ƚ$^Um�
�2m쨐޼�y�%�G������T1�
�`^��kT���~�f�v�����+�� W
�w��y��|�;�V������]\8[6 �4�bY��C�;O/���2��0L)~YX�#��׮�"@V
_��ueumL��#�t:�DN���e�@r���mؙ�ϯn-T����q�WV�ˣ�۳5��GrӤ�\[8ȑY�(^7���_��]����?�v8��Z���|>"��kp�4]�g��o.r~���C�L���> f��pT��w�qv�]��Ȝ����F���:h�fi�4�8A��3=z{W�d�^�+�Y��껦�o����Y�8u.���>�C/���5����J�v*�'�a��3�c��X��/]_]���c���5�
�HW���w�#���%^�yX�
��d��Cp���D֢B�j}��~Z��ҸF�u��=��i�"�޸+�e
�_]�v�ͯm��g{�x�W��U���H�hw���@�:'��]A��|Y�;~8Mw��VMu
�^�U���>W�7]]��"z��J�!����ks�_8F�FI/�;�"�Y�P�K��;��#�ٵ EήC�[�ɸ�u���8�'<ք7M~g���y�%'!��H9�=r�X��ގ�SWՄ����}x}揁��4��M�ι6����G�3J����\�q��P�>ߴ�<<���)�!�-�tl��t�UiC��ʭx�~�ͮ��߻�I��@���t���
����`*� ��F���2q��{g����vg�8SKD֬�b�>�C^w�� �=��8�����]��l�M
�����O��ؼz�~���z�­�=�����բ 2ؤ2�S��s����{zg�t?�W�%���1����8`�R�L�C��<ʄ�z6�}v��c��i��w��@�-.�w�q�B{� �/`�qv���뷜�m�m�0�:C��4�����9�E�J��v�4zWI����'���[�k�N��Q.��ce��}y�ޞ��]Ba0�F�U��Ɗ���h��B
�����y��8�
\�7��*�[���o�>P=l<�� 縜m��� ���5��\x �ͩ��c͍�~in>�덾��~�`[˃AP0���^�?V��-o���H1]��b�ŀq�C�h�5a�����~����}�f�3uб�+��v�a��/�I�_zNK����~�h:
��b8(��ݾ�k�c�t�k���p�/�.ႈ�eL���x��R��^Mi3�O<"d����t��k����%Y��ŀ_�0zV��½����3z��!8�k��
�pO��ʅ� �g��b�>z���B^=��� ������z�Ն�(���R�j	�s3:)�flP��f��t1s쑳�%[���ϑ��v�ﾣq�9��2��׽�X�
�xR�96`�;-%Q,���دj��<�&�hc���YP��l|�=�Yc��%<�� �Q5/�t�^�E-�O�Y��HK;O�3uz&�\?{�X �3 ��Z�ӌׅA��ޙZ��L�	f���7
A:5�E����s>ö�������L5���Q&�#�0N���{~$h9`V�#b���R��Ļڗ�z33θ�\ſ���:���ع��x�����T����8��/��/'=��0�D�(@\���u-��N}�|U���՝x3�@���W��B�01�����1�{ۦ�#���C�[�^N01RV��kJ��[��=Γ�~	2��e=ס*��˛׸u7���u(l�n��/l̳�@�+��Y��ct9Jǎ̺٧)��S5uf
@Y�!>.fE�MY�n2x���i:)�i�b��!9��MM;X�q �Ǯ�3ݵz��]Jk;��g�ڴl �,ގ���FP�/>5����_Veib���������r	��:��8�!�q�ƈ�]�5u�Q&�V��"��nkf�,
em����O���gV��x��*�8����ī:�x�����t�oB9b3.Of�E2�fȝ>ѐ���B(k�[�W��z�h<s8��"ߟU�q�-��4k@kvb��	W�1-��"��*fTf]��hb��X_R/Vp��"��Y@�oo,�3�h�|�Z�`��2�������%(��x��[��ԥ9���Gu����x��L�}��         �I$�/.�a gu.�7"���)�v�P��Y\�1.W%d�zá9��j��t��#� Ҝ��nqMJ90�J�8(��K;n>5�X9[�a�ʴo��zMB#iuC���dV�z���ģ�uofn�f�M`�u�ص�g�dF�n�Ю��k�`�T�d��a���oje%\���m�I�1����OBN�۫9��; 4 U}���p7Q�BU�^�t4gm:&&�Yh��:4���p3r]J�X2u�m3��a�N1�@�Sb�Wk��Xt��F]�����#8�qV�N�Ϭ�ӷt������ٕ|�[�`2�	�f�.�,�m�S�=m&&��$b1ܼc%���(��4��i6HL�A�U� ]��}��|�߾xTQ^Y$Mf9DM=�ym�5fPd�U5��e����­Ye��bjh!���Q��+'�0U��u9EN�YEA�ũ�ՕC�Vc���AQ�r��ɠ�!�a�,̈����1�����H��0�7�5SATT��D�U�M�}bDEFDQEUMoo�G1�o`TA5]����𒳳f��A��w;�t�Y���6a�����+㻯�y�ZW�
C�X��U�C]�а4�-�+r�YY��lS��\v�+��<��h҇l�HTg�(�c��ܻ=�ɽ�B5��� c�i�v_
4]�öD e�1ۯ���y$U�g��
��]ڪG����H����!�
�Hd֊h�m�|�,�p�
>�cWs��?Ou�L�P��߬�T]״��'�����"v�uy{s#S�m�*t�E�G��`�>)�c&='rI7�4@��*��VhA�&��~�����e�{$���ʝ�`�1,�9��p�P~˱B�~��2w/�z;�_��:(2��t��3P3z�`�;���������+��{�jB4#�`࢙6�'�,�Ff��x�G�f6�4Ak���;��I��Z|�Wi�Ky��}Z����^B�:.���*��&١����`�V%�K�Jb���'�����5�~���Ƽ,߆�+!
�0Y��¼o�aSHz�űy�%xԹ�:i�!���c�-����8;z�~��&Ոׂz3�K�o�
�r�+	��X�^Rm�o7�"E�F�3xX���.�x �_\�^c�����y�z#T��EF:d�5����0y����d킳������	CD�v��/Ƶ(��yos���Iy/Oz�0@@��^��C�J�YU���p�5�Z��|����!h�:e�$�5��S
<}3=��MF���\3;3�RKD֩dP�Јk�����A7��O{�\�)��V���t��>��&lIs��{�:���N�,�ѕ���Eh�üB�F����/6��!_Nw�t@4���BǄg����2E�>�Q�/��W���������¶���о���l���D�� i{�Vw�!�3����U����"��`�"#N+T�5�j����H�+�`�w~ �k����ul�L �O-��4���ϫ:��
�V��P՛*�b���Ǝ����~֗�",�[Ċ�Q�*�}�b�}���olX�ۜ��nB��i�c.�� ��>����xi�M͑�t��g�\�+�@� 8f�+�֑��6��&eeq�KMxuW�e� ���M1D2]�p�w���9p�(8xx.(<�n�>�f+J��u��Cv0���*�@Ϋ�ɩ��C���}SݦEco4,�U&0ɩ�z̾P̾�� ��@� �Ҋs˃'���?{��W�?��йlb0Wi`a�[��ru��/r���)c�8m��}}���A&�eL�����զ��L�j�ߟRy�6��I�@h5���՚���E����z�p�.�G~��p�V��&P5�����?�
���Fih��[>�kYB��;���ȳY~���u�P�w�9��Mh���}����$�z}�O�����d���xz��� �eׅ@��]���z�9~lH��H�xW���<<r��]�Q���5�u�p�����3Eum��.e`�WV��G�ՙ��<>��9�{�f�{���xeW��]#L � )i-U��|P;՜���-�ِ*�7���r��|ձ�U!�%�����[�}��of���}iP�L�R�@.V�j�f�����?��tM��m��=߭�[���c�����s\񇻜6|�����ZP�r�b��Z0Tf�K���!(@i˃�ӵrո�I�T�׆���+
+��e�^4ΙB�_t��5�����g�kէIa
��n!xl!���˨kI
��{���$�b������4i[���MuVჄC8t׶׺w��4~h��u����Ф�^����먞���FEJ�!j�l!Ⴆ���F��Gl�*��xꜻ�w����a�>�XR3�����}��D�J.*Y����?��R�]��w\*�n��|�,�p�
]��.�D�q5����
=�DxT��g�pT��e�h��Q:<]�WeѼb��ʶ��Y΢�q��;/7� ٩.+�ޜ�X�Yr���$#�W�X�qLGglيk'���t��=?|^b�߶��L��(�Q��"(Sߝ�`�>)�ۃ<̋&��4M� t �ۺ@�]�G7����Gw9v�y��G�>ʅCbebY�}����p�!����o����"8����@2��F˩�j�c^��N`V�)���*���d�f�ۤ.�`�%���s��
�/Y�����4�՟3�x4T�V��Jշ�z�^w�BP�4�;�������J�smo����ja�W�jfS.��]�ZDc��g�ƒ��ҝ�h�������]c�2":zroת%׮�g����D�n����ž�3�EF�[NF�g�au�z.wEYه0��mr�����e�5$}����N7�e;Z��JD��Y}�U��$y��fkb�2kz�z*����n���o��*��Moz�Bޗ=�����~QFg��r9!��G��Q�TL�H�n)ͥ�O؝�%������t%���8�u�v7}�ۏ�v�-G�uZ��@�;~��bc���M�mM^�Y�����Q���}�^j���o{��+��E:���y*���a�F�s��=&U4�i��6�6�����
�n7~�F��Q6�{�J`�R��m��T�bi�B���_��؁�;oPǗ�,������t��{tS�+�󽌼��I ��E��ۏz�	��)"|�����o^�FS,Q��G'l������F���V���RRx��2�i���"���Û���R�9ނC8].)e�uL�5u]��OF(��O����<��g�!s�C�,_i�������%㺯&�ML�ʁ�R����W��t���\��S��7�0�GA�w!�tj���֗k���^�O)��Ѕ��Nw��
�Ӽk�gc��j��I7��*��]f���?c���������Z�¼9���/B�_�������pt}VD��޿n����G�X�-B��hV{
WF�
�N���V{h/e����yLq�^^��`f,Sq�*,��e�bJ��~���n�_�/�3H-U�#�8-��e�i���D�_�λڷ���)�=5��+���^��������]�$_5w��.r6���'�u�z5׎�i�<�|��z/#4��f�i�䯼�]��pя�[����gK�*Sx�Lޜokd���94���븽��P�έ��/0���؋�s9�eM���8v�����7�V�k���N�i�ƞ�Jv31�O?J��נ�ʍ�Ǐw�u�ȟ�HkFzzǼ��a�2����=�k��=����Zۍ�GLJx^5�Փ:�N�� )��[��\�(𽴩�Q_\*É{�,��9�O�IΞ�?��t�.����2�t��ȗ��jZ��d��O������QoT���5���v�ҧj$�hy��Z�y�y[����twָ��2���+y��ד|�z\۵�u>K�M�=�mp���f�����=Q]�g���!FEe�W�e���B}��y_���bs]-C�տh�{����W�U.�Ht�T��&F��j-����)Ď���]i{���]L������ÎB���<��MW�M�9���)���/V,e֪���[�NrӜ��p�6)�d�tju�Ԡo37AC���ӛ�<����Q�YH����)�2�7�b�����tV�-8Rݕ�YS/{6��V��M>g��76+���xA����B"�G\�X'�(v\{Q3N��}`�N��0�=�X��X;��gK��}�]�#�d��5��Z������l$ Â�J���#X���R8��5�8>}��__L=�k��	YDu�B��*�yxV�e���T�������M�X�
�u�@uǉ��Ge�d�z�=kd�U(JP	|�P�z�L�6��۩񶫳�D��%��J��f�Z[3D�|U�omY�[+ �D������,z�������K�e���!�1�$�AE��+�̛�9�\����vf�             ^S�x�o*&{p�sz�<l�\�%-Ύ���M�e��K�*�a��!���T�@�w���	E�-�޸\ۚ9m �̨�����������o�Sƞ:{ғ64�2vm<�+�	n����cYHl�"�F�1����ԁ�}������j�#n���$ɜ2��o%XF�r��c
5tv��WY��ΖC������reg@je.-��Y�Vjn�J�̤l�ys u�V�uخ,pф��fVG�۱+��mط�������8M_G��f����͟ozud멩qʾ1>[�{�:w1$1�D�xH̛�N�:v���w������6��>�Ѿ�D
v]M�d���ؒc�T��d�=o$ܻ�$�G�}��}��]��S�d��Z�*�j��b(�lMN�(���Ʃ������1������
�&��
 ���f"�b
����Jb�M�`9Ō��DPDUI@UEE�QQ�8MT[X�m�H�U��1��JX��+|� �(���Ģ��$��	�7����\�**"����j ��*�̨�f(��*�lk*c|&�
��Q�1%	��U-E��w�3S�z߷c��dN^��}|NS���tì9P�&�ȭ�ᓓs��U���p���t�����]�7ļ�G\�:4�,Ƴ+)7+=ܬ;g-_�6�cĽ5Lha'������ח�[^^K\"b�V� ���}���Ίx��uNwZ���RͣT��n��y�,i�԰��5�ϳ�#fc��n'�ӷ8or�j��ۦ�%�������;���WYEI�s�'���]z���^���^�l�gao�ܛ0���ގ΂�2�g{V�Bq|��e���zq�21���^vkԦx�}�W�X�Q�
�W��b�E_L��U������^�G^�R���OS�5��2�Y�ȷYf]lA����:.ɕ�U<�q�)������o��-y�m�Uݮ~����/Q�z8��\��x�hO}J�Q{d�̯�+�e�T=hQ�ﴌ���{�L�X�׼���&\��©���8����W�Ư�9�ڳֺ)�\��y�uɥz�u����c}ϒ���ESoz���[�"�ɮ�F^�7�sp��nz1F��1ѣ<��Ot�~N�����£y!�k����%$|WJ������|��r%�w���M����?�Z�%�hW^&�K�6�2��� R�o9e,㛹ʺF��k�d�@�6,��j��i�8�|�u���[�C�kW�9:�]Y��f��6)ո��L����<4�?�OsW�ѻ����8� t�\[Yؗ7dn��SOL�]{9��(8z�W��O==��͛Εִ�;�۵��{�8�j��E���jq�{�*�K��nUs���(G�����sxe����0�s��S����^�t^c%wu	''-
N�WR�^�Ծݯ6}9�n��Yr��\:]���;�NW��&����d�0��:v��JC�Z�"r/y�p�g����*�Rv��-jtfSǵ	��u�W��&u5�[j�M)j��<�rEI�(�A՛��>��Y���{�Y̚�6�s�s6���s��)%�>T��P��fNB���hLm�iF��jnl�;�8�PK�՛�ҋ��ك����j!)�+n��N%���f�|f�������\O��)���朇�F��ב�]vv�jo�ʜQI���6eg��%�:�����m*��W�r��L�7懱gr��ﲔ������sظV"�N6��H#�=��}�����W�X�*̷,Y9ލ�N����O��T�a����֒��&1��Ko+��(�%� �SV�
䘵��@�+"�@됊��Q{��� Y����ۓ;��=ը�X��P���nw�;�ړB�wp�V��{�I����6��E�T]���2|�|��n�n��W�������M�^U���kJ��3|�4�Փ����z�	�%w��AM`�?9��8ת���	�t}�Ȯ�9=�p���y}..�n��^W��m���B�b�{:6ƫ�RޤZ��V��R�2���1���鞥w�O?_Y4ށ�yO����t�w�a��x�j��ꭜ_:3Z5K���E��`����Ux�\�U�щ�9��8��Y!)�
��b���j�����.�*5���+Ϣ�6i@�z��7`�����"6�Ǣ�)GY�WNɈ'%�V�m�Ӂsn��Y+
��sz��$��u��3WW�� ^�����ۢ�/{�,��ɪu���
�?Y�^���1��l�Sw�H~n=�#�OE�݂��q�2aw^�����OE�T�����$���ކi�lE�LE\��s�+�1O/x�&�7�+OO75Jm�F�昽{�Y{�[W���w��&�T�:����8���;{����`��{٢yc��OG�饵�	��V͎�륝�%�󞖷�Q�۹rT}r��7�����M��ka��5�Y�cU��n��֧ղ���t�%�fM�g^�v#Z�,�.;K���8Č.�u�F4�J(H]�y���{��ɺ�9�b*�x9���~;�����O
>f�����e��E��C-_��lŽ�;YQ������e����%�iqf=&Vg�	�j���5�Ft�Д�aW��m�jڏ_����ks���޶0�J<^�tԛz�v�vw�y�7��{�GL=�s�؉��حcK�-s�'ӽ�i�+��Z�b�m�֟�t�~�x?�:��!^��):9��י>���ʮ|�'	w��"�u�y�5����U�wvm���yL�-��"h�zn��=�,澎�]���K��!\����/FE�ĳSwgN�]�	_/Hg$(N�	�z��or�����Jս�m	'R���Ñ畨'�nw�<��bIsg8�����v�֪�ߝ*}���Zn�Noޮ�k�H��ܩ.�Y^=^�՜�j�|��N���������k����t\�o��ՙ����j6V vaL�o��͘����tRb���5y��c���.�4ܼS���[�`����Qk'�5ǷY��z)���fde�wk�+oMk�����덪>������}<�]���;M�naض��P��Y��)�Sҋ���w��g.m	a1�U��:K���5�݊��뼟c��H�r'�N~9�k�L_������s�&��7�s��]�Y����~|�w��u�����g�m�H���,���*_Wev��ao|����1Y�3�̉0Xuy%�7�/��(엣')E+�b�2�K�Q�x��:�R�KWy��:�>u7}]��,����+ݑේ�\��U�9L��/{��kiL�.���uq�/Y_J47��z�yy^Xu��V���b����;�K�>�v�r�Z��R-̡}=뮞��� �(���;Qp�T��5tb���Zj4^c2I��1����%9CP7x�.:��FFqN�WD�E���Rfi����8��u'���a�V�_Mx�mf�����p�E��l`�Y��jC����v��$K��#�f�����m�q�[m��An�M�
�tC�yw�yy�{�>�Nn�V(G.��&v	KZ�^f�S�;�MgH�g��
�3C���=Nx'��^�ڧ�jP\������:O��Jg{(߻�K�\T�<z�}����o���A����[����~�t̒�{G�+4b�7V��]nJ��b��c���Ǖ��4����W%a�\�A3!��,�E�uS��^�喞���0���<���]R��ƓK]��
��Nck�o�-p[9�Vf&�3�*%`�#]��oU�w?IR��B�[nz��P����;̱Gj��v�Z�0��x�RC�W�.���q@αW��+��������n����p�<�6�'��.�l�v�Ҋ����e��j^S�.��u��R�$jhc6N��iN���}��G/_A9��u
3����B5:4錢�s4�B�:[�v�
�	wu���v�lw^�2J���->��@����BA�V���eZ��폏|0�K���S��V��7�Eq�.�������5�.��2�<����:|�P���>&��r[5 ���շ�1|�2��U�G�}:�v�����+��Nr            �H�۩�jsg!|�� �R
ܣ�� 9(M_<-�c
�I��؃	װ����)�ܕ�Zp��/�~+�����Ouh8��^��_�u��+���ż�*2�B�Z�+�I���<��0�ײ��,:���	�5B�Yk;���6�#��MN�_"����f�u����EF��(m�s��_WU� ��kįS*�-/g-�=�-�����NP�;E<��M��Z�2WA����F*�9�ثuIf�uq�.���낓�C�-�9�l���;�UEqv�������q��hK��)(ȳ�e`[��@5�n��D�wН��+R{�nv��	\GO�b��pB�ʀ'�i�U���i��1Rrl=c�k�����   ��
{홈�z=��UAM�aMD8�VP4% Z�2M�rZZZH�x��)�C h����y�P�HeMRI�F@�X9ՙ��1UP�a!CHo�A��RSACHT�f�jֳR4�%H�&E;˨MK���������r6��2m�r]XZ��l]�¥�h��,����~�����:�t��\��_� :96��u\��]i�/�?��mI�/��~���\��{.���M�?u����{�m����^����PF�y��V*~�=�ދԦ�*^��?zR�{2	�Ɏ�n�;y�����ם3T�'��rY�^�eY.���OS�=�!�xfE��k����7����#9�����\�|��~����"{�H�x��*e��ɷG'{o/u|�_k�o�^�#w*7����cO*����jQey�N���"�Ml.s���l_�%�{=���<���t��ޙܷ呗7j�Gs��j��}�/0x���+ �/��,d�v@�kp�1Ĳ�7ٸ�����s���pmgWe<�p����Nq3�YwhHq��=�^�^�u�y���U#�=��<�s�w����w�O'���t| ^x��|�JeY4�߃�a�~��'�*Y�7#���1��N�f�
)�ݽ�;L{T�&���������-"�ܣcb�q��>F�Q�z*m�qpXNJPg(�>�3Xؙ��P��\�:-ڌ��ZMF�a���څ�<ֽ�Wp�/����4�z
���$�Ҋ9�Wy:��'�m�K}��k����_�U.�ZC'?��{�u(���B'�~*���`/K� c%�}T�������w;�wV*K���p��-l���t��+Osg+`Y}�ʷ[�'0�g5L�؝��rxI
�<S5Qf���d�귮p܆�UK4[	�m�/L�`_qsޞ=׏y�O�Q��N��,m��vgMG������y=~}^�c�w)�������Kw.-�]��,u~���tr�t�ډ5�۫զ۹�ӏJOӼ�:���~������i絏^�J�s|�a�mF2�'{5�"�ίf1��ƟNDJKVT���Q��;�j�/j��7Ρ��O�!y]!����[�e}�*f���t�s1n���\ļ+!0�c�RV")/GPV�븚�6�^�^���݊���]����̴Ƒ;6L�V$i^��1�ْ[�opeΐ�I��l)�_o �{g��.
�5�n�K������(��{/n��*�bwx�7qߓ�����N�u��[���J���ޝ�]B����eꕈ�5��yʹ5�]�U��Z�����������n����L��s�أBfo*�q�"^��W��dv,��;���=���,W}�8�ܾچ�H���Tf^�xVy�7$�[Տ�ekC ���磣{"2ZK�9�j;f+�y�j�Ts>�x���Sl�O>S5���N��7�%V�2��_���+��
�OV]�aN7�3��b��j�9�雜ݎ����q�ydh�l����ZXӹ+A@b�]� -���ǋb����2GI��׈��[Y��ჽyѿ!�C\z�>�y����]�nV,��&=s�.;"%:�~��\�q8fa+4Md����ޞDʦ�^��Mr^�W;���&�{�_�S,�Z]Y�v�rOF��Z[^u
�@�:���ݬ}^��i��'��3W��%��\�����{);�2�oC��'yn��9�G�뫪xu��^�Mw.�z�=�}�᪽�����cT�^�]�g���0d�[�6:��X`���t���[L����V��ݒ�!�6C���J�S�j�WP(��Z����ƥh���,�䄹���Kcc�4�b�����=i$�ƑXb���a�*s=�M�v3#��|$��ʇ�X6����*:��Q������^���ً�Ǧ��1*{+�mǩɼ|�O���l$N�^�UG5$'<�<q�Ǿ��p���F�������lW.��5Y��u�VU���v�{�o���m���Eo��o�!YI��Y��ks������P�ץ�!}�����Pm�KG=J����S�y{���+fب�f��W��WsغՒ�wUi9N�juw�n������Ui(��
��ڞ6�6/W>���vNU0|�\-w0�5c�4�pY���}==~�ýJ��%���C�nq=�{}�I��K������3��mMR�t���p����*��
Ȟ>��5�;Y�s�'�~�Ϋ�=W�^_]߷���.�ܶ�9�1m{��Ǿ������&4���ku_�%�sP�o^������4�-kN��.��2����]�zo�z��V%6l�=�ᬄ$����Y"ĭ=�홲H���,r��J����ϻ6�{I�o��zV�(�|~��B�hۡN{��+~�	�V��#��ݣr�.����W<�������A�"[[k�������,*sj^� �(bmQ �m�X���Pn���0qw9�7���k������T�~[��^�;�ih+ǫt���y]�J}7��D��i�藥Jڷꋮ=��˱F�
������GX�
K9w��dk:/����Ǟ���/�g+�Q�7�y�;}��ƽ�Ih���������:,��Exo�[���p�z��P2��.���9*̗9R-tZ��=��4��ǚc�|��3����c@ʌ�5']�x�M?LQ~��]ݟ,�,�l���k4�2l�=4�6a��	��O��gK
�9]���������({��)B�Gy���X�ʆ!���#��x�N+�����������,�[7CK7�D�-dō�nWv�����n)��r���-V�c{�\-�H{��5�����}=��x����H�ʒRe⦳�F+��#��=��?x�O�9�&����hר�ϯ1	�9����{�瘮�س�f���&��}�%2�KZ��^��~��п-��k|�f����\�p�~^���frQ��L4��@�m=ެ�l�co�]�s�!/>5�]g���S41���C���~�k��R͆�R+q�eꃛ�2� ��[$�v�]m������/)x}\�+]~�����R�5��-&|G�|Iuu�!��t��3\D��y�F��앿sa�I�r͠���4yxe�k���.
��o*�]��Y��e�@��s�������I����8Q�̢�=����^�����=!�mI��K��5�W9M��Q�`��~o�wE��V�:��W�8�nF�-���Q�:�>��ʁ ��S�Y��6��z�=�ysV���E���f�!����vx=��,e����Fg�����vq�ΦO�w��i��n�]ϩ�Ɨ��=of�xq��:�u�]����}g��_�Q��CEE�S0AD@Շ���D��������m��Y"x�0�4�Ɲs��bmq��A����6��#��E@h�(���*(  $����;ߓ����80q.01��a3��?�X�×�7M�=����H
"�C_+���g��G���>��r�a�L"4𻛇ױ��5��Ѱ���s��u飠���k9^~i�Z4���;���(� �'���~~��{�����Q?�%� @��Z%&.��>����!>�?��8���w0�_�_�'�������~ �w�Q:������!���u4��%4*n}�덈N]��}!�&�]�����3��l�������?(>�?��������í7�C�M�@Q#�������h�5�"6@Q6O�k�e^�ިC����2��o�׮M���!���l|�AD@�/
pMR�������6��?q��7L�M�/��p��$�����?K�ۀ�=7?�~G� a����ڹ��������qD@��Y��P~�|��O�����?������|����)��'�}�~Ϸ�8�? ���~k�?�x}���W�x�����'�~(
"��K���?P���|n=��h���0?h}�	��)��A@�4�AD@�����H�-���lk���g�������0��~�p|��
 p�� �� Ӣ�pX?��~Mr�� bK����)�Xp������׈IƲ�p�.D|�M+�?�u`������N���[��((�:�}��~��O�O�D@��?��7�� ?S�?���>>g���>�'����M����~�o�?TA���p?����?)?�~i����}_	�m���b�������>w���&a�����'I~���~t�����P;�z����?@��G�O����Nx�P'I���bb����O�����?/�����)����_��:�r=�����.D}�h�X�&�zs��ih>Y�q�'D~�C���|��=��$��~�3���M�0?��)�z�L(� �_����??�N�S�G�~�����QD@���?��<��'��`����!�:��C�k[�)�Jb�H�#?/O�~o/���H�
�W�@