BZh91AY&SYy����_�pq���#� ����b*                 �                             �(
!T�"Q>�B�,�Um��P  `h@��I)�1H��@ �0 ��!� �  �    R�  ���4(�$�$PT�� ��T��B���AR���%@(%%UIUJR�	!	"��$�C�i�kwrv0���@�P���RP; ���Y7Ѿ���D�77Ӣ�p�E/@��Ƈ{t��þc�D��6��:�X^��;�����  ������i[m�5Ow����K뜟}�zj |��/= �}������ >^�� �������0������P|�;���  ��JV��k@��H"(�)B����D�_: w`}��<���=>��}w|����G�7��T^ ����� ����=��ǈB\�A+��p��Xﳠ�  P{�)**F�p;� ��=� {�>����|��tA c�7��^�>� ����@>@ga�}�>@{��9w�� yA@ �Ғ^�V�����$
" Yj���۸���9����O˻ʊK�����9}}��;� y{�QB�G��;��  =��R����� |�r ��W�^�@u�{� ���0��� mc�`���� �d 0@ >�E��|P
� �
U%(��DW�G�s�7`�� nJ�� 'c̀{��� �}�ψ w��U$� H� d   ����JR�^����� w� �����Qް<� vw� ��T�`@ [�7` H � >�_l(4G_ 
��	
�@%> -c�`� �;�=g��[�!`!�}�}���=����=
/ w=j�;�(  �}��Q�}`�� :�H��b���{�# K΢�������C� ��`�   
@P � � R�ɔm4��2&�O�4��Q�  hd  �ʥSCRM @    O"��T�@di�@dFL	4�J�       T��?R��h�i=C 3(��~���~��v�~�P(V�hV��(N���/����������� U�~NAr�|�?�@U�A?Z(���TP_�?��$�����?�~O�0�����?�S��V�r���J(���p>�/���U~���G���M�� L����0�� �?��!� c"��2.0���L2.0�2�¸�8ʸ��8ʸ�=2�0� c"�l�(�L�+�+���������
�� �&0�l8�2/L c�
� �vʸ��=�0cL������q�`�1�x1��0�'��g1�g1�g1��1���x�0c8�63���l�&0ct�3��=�c8�1��3��c8�1��3����8������1�1��1��3�8�0ct�3��lɌ�1�g�`���3��>0c1�8��1��q�g1��0t�3��0cx�0q�g�Lg�0c���8ύ��`�g�<lg��0c8���c3���L��3���q�`�q�`��&1�`�q�`�0`�`�`�q��g1�`�q��c1��q�`��q��`�q�1����8��8���60c8�l�0c0v�����c8����&3���c8���1��3�c&4�3��3�c�0c8�2c8�c8���8���8�㌘�0c>0c3c&0c&3��163��0c8Ɍ�8���q�d�g�c8�������x�8��g�`�q��&3������`�`�bc1�g�g��q�`�`�1�1�c1���1�1���\d��8�������0cLɌ������8�Lc���;q���l��1��8��c�q�c��q�g��3��1���64�1�c8�1���7M�c8�lc�3�c8�4�3�c�3�c�1����1���c�3��M��0c8�0c�c�q�c�c�ǎ3��1��<q�cc>1�c�0c�1��8�1��1���3��q��c�<c�1�c��8�3���3�cLc8�3�c�3��t��1���c�3��c<c�q�d�1��1��1�g�q���q�c�1�`�1�c��1�c�1�c��c�;g�ǆ1��ώ<8�1�c8�1�c��q�`�g1���1���1�1�c1�g�1�c�1�c��1���1�`�1�li�g�q�g�1�8��q�c�1��1�lc�`�1�g��&q�lc�1���c8�3��3���1�q�3��1�c8�1�c�7�cc�c�1��q�lg�1�g�;q���3�c�1��8�=<1�c�c�1�c��g�c�1�g�ǆ1�1�c�1�g�1�n��q�g�q�lc�8��lg��1�c�1��1�c�161�c�1��3�8�1���3���8ǎ<8�3�c8�1���7Lc8�3��3�����x�3����2������0��	��*c � �8�8Ⱦ8�� c��&2�02�����#������������o q�q�:`dLea``geL`LdaddLdLe��1�q�1�1�1�1�q�1�q�q����(�
c"c*c(c(c(� ���c�����#�)����l�����
c*c*c�(��(c#0c
c �*c
c*c �
c*c"t��CG�T�A���T��a	�q�`\eLaaLadc�)�)�)�����"�c*c*cc(x��)�Q� 1�d`a``&��T��A�A�T�P�T���W�D�D�Q��T���&�T��T���D���W�CSC����D�D�P�P����D��D���A����S���	��)���#� c3*c
c*c"c �"c!� c � �(���c
c*tʘ�8Ș�8�8ʘÌ2�0�2�0�0�0�0�0����)���������#�)��!��0�2'GS�(c*c �"c �ʘ�8�8Ș���*c�¸�8�8ʘ�8�8�L�2�2�2.2�0���c"c)�GSS��A�T���A���WGSSx��� �� ��8���8��������+�(L2�0�2t�.0� c"�	��0&0)� c ʆ3۝�Q��4?U~�^��Θ�.���Qx�f�z�ϕ&.��d�q�H=���\�A��rI���b,������r&(uV��d�/�:�e��|%��dy,�po7q�]8qn@����}�c�r��R(�H��	�<��w��%�{��Ȼ��;��:X�H������(=K?Z;+��1��]&^%n����ǧQbp�n�n�P��&��Toh�jb�̘����3��զ53�kjM�'EY*4���q�7�ۃ��za�-�Z�Ӌ�u3f�dv����c�3�gD��Ύ�����#,O:Z�vu�gU������/t���;>5�y�2s�Mٷ^�V��u�#On;����ţ{a:�E
sW.����0u�����9�]��F�nn9)��u��I�r��y��cQ���f�ܢ��K{GvO��X�0��Ql��P� ��)��.?�[�/il���C�
��;�ͻ����X�;H��2bc�Q��$� K���(���E������hy3^N|dBp]"�׍�R[�ք������Վ�^�>mgP�ھ ��^87 ;z��Z��;9�]&n�5kks�/�n��a
T݊-����9�=N���*�E!&m�מ}=�g��P���q���W#�7F��r�gn�؇]�8�3���x�Zw�b�-뽺Ɣ R��k�+��q�ue���9n�޻�AZ�y3u��Xa�� W�ql� 4�
UQ����u@7O'y�⽐awp3��斀@ɋGN΢��,��8�
/d́��"{&)z$ ���a��N������!ܴ�{�,1�Z�<�'z4���{����u�lL�|�ᶫ�k�sxa�$ܻõ�v����ae�h����8��9�J�̦�]�k�5X�c��&������s���Q�X�d�V��3qҀk����h	�d���K8�^����`���|�nR�s��{ʺE�(���J�_o-?D���k:�ɱ=��
^����Qϵ��H.Lt��Z^�V����c����qvI�����6wM�;3c�[�sw#��\;v3nCK������ڡ�U��8@�E�W!�� ����9��o���ǒ���,�[�.��Μ8W>t��}�M��V0��6�+��{�L��#3-)����`�sSf�'�6��7{E��-��tɓ���f�u����2qJ#�Q�q+�_N��h�o{屭�3�9��m���D#; ��!�(�4�#�]���v��7e,�/|u]���ݢs��N�:��r�w�8o06>�ׯl{�&�Z�ss���T
琑۸S�˞����9x�56������$f!�hFLL��r�P]��yG�&^�;�T�D��q���ռ0#��e�0��=�s�!oua���`,�����!��\��t:����\՚ ��s���ޮ��g���L7en�����1*�� .OnY�sct�,80��xgs�wd9�!i�Fq�a��WV�~��$={w����ȣ,k+������7Gu�ŗ��I��&�ў�����]ԑ��Xm��(��	,*�8q/V��ź�kV\ۺPP9���x�ά(N���Ϻ��V��j��\8���$�f�7p����(��9�L7�80�d��Ƶ=厭4<L����l��:����)���;xp�P�]���Νvs&�~o�;���_s��v
[�l�����!�I��vr�a >�xos�Q�t�>�R2�YȰ8�^���vI0��ˑO�2��	s
�fM�`�).Ŕ�V��13���t�6�p[�1gH��q^"W�p��ST��S�s�GX�GY)��S�%P�IG{d�n����G|�o����\�vN���o�zq�#�+Ǔ��P���g
ZT⺫ua�����f��̡~{
b��R��w-=��Fw������p������׈+i��`��δ�J�l��4_�h��k�kL�Me�E�����,�=��I-�7W=���uӱ�ϷS{�+�gw]����ˈV�0�`;���!�:n�z-=S&��1}��I��ơ��I�3��],�)xP<�X�hA�N���R�ǐ���`�w6�s��f5�m@����+㽎v]���#�*���G,��D���+ۓ)\��oo58��#�/7ל�]�g�H���������gJM�l��-n�|5p��u��+5��^�/�v(�\���
Lx��[��F*�ز��&:��䯻��k�&r����6�)�6̈́28sF��b��ȋ�,�g}�(�o��8
Q>��_1r\���4�}�
i��7w�Pt\ս�rG�	��%�ۣ�/k�LJ���8� k3P���b�5�Ǭ���PL�si��.�wL"N����QZG��I�r���0r�,ҒD�y��q������x<X�"pD�sIv*��V\��;b�8��m1v+ò����
�y8��%����ǹ�t!����4(y^�"�Z�޸1C*���G�J���/Րr�黮gC�V�.3Mo�|�%y�0d���{ݛ�{��;��q6�Z �$!@�I�H��Y�a\o>=$��������]ם��{^H5g;��)�/�'�u�1(F9��hiM��48i����.�j�k{���!;M��$h�-�3i.&��!��7�r�LW^c���!p������w'V�x��J���� p� �4-�eǌ�J[�rpY-�J�ـb�W2�wIod8�D�;t�K�&�>����6�(<=�r~���ضvx�\J+)W7g-��DbIh�NoI��8n�U���sJ�4]?pd�g�G����ѥ�0׋6^M���K{����p�u<�TS��A웸-�_tW**c��i��n)�{�k9��z3��-��
��u��f-uv��t18������.С7�n�H�tê>}�G�RѬq����^ѽ������&��K��4mc��(��A�޺���4���V)���m`
,��Z|�ɮ�ib��n<����{\�c�h�������78�>��yh-�8�Z�.lm�^����#�᫉Sv�0
Wn�D�H{y�Ǭvn���2pgl�pg`]ܶ�k����5u>���B"����T�4��C�&qK[gGڟs�d��D��s[��l��&.�*),�ذ��e%vڇoh8b�J큇t�ʳޯ�����9c�w���� S;��u����4�;sRU��{t���I��1Sy�n�'���� �\d�Kn�kZ`\r��T��N<�����*;�յ�M��b�0�y`����|F\|���7m[�No�{\Z�����gw�o>����n�=���0�j��sv���K{���&L�ڠ�����n�`�ϊQ=9�٫�K�Bٚ�Z.��y�4�*]�s�Ʉ�:�+0���Ɩ�aX�<뻍S4v�3U,Q�v�t�8�#^NW.%�v���ިaٚ;C�;D؊\�!�ɶ�P��ʓ����&�66@�7R�l��x��P��!#�7�D�|��TCu��p�ُ�:�f��&ا<T���*�����A�hӃ����ÑM���os!s �q<|�u8���'�u�mn�H�2��Íc	�1�5��Cѳ��
�<�8�'��׌� }�ķ��^ك�p�$�Y"��:.Y݋ ���ɀloq[������ިg*i@�]�H�y���� l���UA�D�~a�;��MGP�
���7�!�
}v���@-q����}d�7B=��f��â�T#	��Ho'�JjmEӇ����^���t\2��|�0�<�q��\��I��2��"]�����& ����/�lI��l�F�n�:M��Gw��~��X�7"��(2c�茸��f�*�u<���"�4Ja�A��[��h�L�A��Co;�ׄn]g;��qb����r�>��+�m�ݽq^�	���4^�9ރ���9��8����]�{5e��Yԕ�f���s�z�H|�s�3����i��	֋���#x��83f9�ݨwΐ��Awbۓ�.���,��;^��L�C)�4�.���x	spHg$t,��C-�,��mH`����R{p�:%yh�Ex4�ٷk���/@�s��)F
^@���g^ΐ'�Ȼ��Σl���o`�5j�p�ɀu�w�5�N��Z��;tG���)�;6��NqԺ9�FQ3�]���$��{Q�ɜ+jBj�w"0�[Y0���-��m�xD��ާky3�*�f�zi�כX�&! �@��dC��};y=�D�g71=2�ӈb�.#���e9���1i�����;��;a��^6����6���Xd�Ҵ�wu� S�& y�K9MX@��0�p_��黿9I�G:z;9uٰZ1�M��*�-�2��qG{��w�����)�ѽ�%�79t�aW�N}�xv�������d�|�VN�~G��d�m�w �0ӡc���.Y�����
�]\ Y7��z�ĈD0�!�p���9�hķ�:Fn���v�㛉�Mé7�T"��	Ɉ�I�u����C{�@��4��8T�;�`��ώry1�^EX��.�@FqȢK{w�,X6����Wm�i�Õ�W9J���8j�\�d!)	�Û� cŤt�Go!s�b�ⷧqV���!q��n�-R|U��+ew�'h��)�Mnn'ۭ�C�젙�{R{��i���H�!1%�i�ݘ���s�����g�!S�ӻ�>!��
:�v��w[�%�)�Mm��JF2o�5|E4��,Ǒĸ�K�t�k�&�n�a��8b$���8f��N�8���n�8��İ�ր`��̓�3�k���u�zcO���6i��B��c�5��s4k祁��Ѕ��÷w)�Ѩ;�:������d;>��1�I�n�xp��q}�
��N�g�����*��s't��_g`��f~a�G;oG#|��NS�{�r�<���Z�.\n� <M��^^���1?g��}�ZV��s��>5�^�2�
�&ױHQ��K���Q�~[J9_%䁔���Q�5,KR�m>��|�T�ѭ^�S���=?#�q�?o�}c������҈��D$�j�UJ�E׈}W�: ����t���pDJ5�����JV�ID�Ȳw��(���#�d~-��!Z�[
<���Rp^�/S�)I��W��I4���I��Į�։h�5�5���Uu:��=�i��f���>��,�����1�o��Lո}����4M(e�[����nߒ�����4��T:H�s3t/���tb���-���3ix���
��=O��?�¡�G����9A����oN��xYڪ^՘�#}����P�=TN�yFP>KҞ���������`'
�<���M�B�������g�o�B�p�`�S)>"�������~������p$H�	>��ӥ2�(�6�%Q�[#�P�F�H\ì���l,�?��ѾE`��Ri(�T.������_�������C���I��<� ��QJ1NIȇ��.�1h9ġ^��e���(���%+�:W�����Բ,�ҤFt��r.�������bt�'KH�D)�ۥҢR�^��7�eg��ҩ,��Ӏ���S�!;�"<�n�������unB�y�گd�Qz��J����U�d+!�T����H&���A��yՏDD�t�px��J��Q&���4��F��*�a�;	Gį�;�f��g+?�7�z���B��.����{�w񌱑1���tg�G��x�`����0a�I��#��i�z�Fx`e�IZ|�d�<}C�'���*�"5L���{��+K�eE���Uj�/��=��zI�ad�^�0�=�B�P�1����j~0=!�l>$�0E/ߏS�MC'����_���oH��I�<��%d��S'S�����έ-��/yL%
I�pL��}�q��g��FiP��X7��4�].�l�~���k$N�B��^�_�Y<�#�����k�<J&�R-kmT)�{�s�������+�JP��0����R�����ʱ+Y
�(]�1V+弫���B�Q�$����D,�y@���t�fq��yc�뽜u��R�)/H�>'��,�1��x�ZZK��|�c<�iy*�D���u
HT��T��Ig���C)��L0g$���R�M*��Rt�$�$��}U	0�{�7IR�:�r�Jڪy�����)��Y���0� �&*i�f��x7Ʋ���ȯ,Ԉ$x�R�Q�P��{E.#uN>��N������#+�>)u�PD��Y��@�JR�V�Rt�H<�e^I���e�	:y����M*���89��z��_m-�1&L+O"F~�D������S�	OC����'��;��R�$U����*��t�Ty8��䁸��'��'��W���&R�KT$�6�ѵ^J�bQ�O��6�(KѺ#|��ҡ�O?S�͏�d��'O�T+ҡd��x�'�;s�ЦQ�QE#?�>PC��KV��X��D%���(���������}:�˽|��m&�|J)��~>7^?��N���� 2�e`d�u��t���ƒ�p�{N�ޑ)Ŗ�����/��JWZ~H���b��?'���^ժ)k�ͧĞjg�X��.���]{�t�.�iM�� ӥ*aH%%��ƵvTL$���D'H��"�RDb^��s!�d)�	"��a����cϴ����-�f"Q$�O�x�e	$�U$��~3�(�Wg�>O�� d��|��_�Ӭ�o'�
�e�R�뙔��T$���B��EƤ�;�uϱ_��p�o�����~�����'^����G?gÈ��@ZE�@(rNA� PP���!Q� �R�T	$ *� a!`�P
���N@����T) 
�A���E�A�"rQ
V���� J�
/!�E)A��A
������A)@JAX��	@�Y Y$Q9	�PR�
R����(AP�Q)AJA
�)������A���y(rD� P�!$
��)��?�������ޖ�+�=����t����;��@/� ���iY _�|�8�������Ϩ�����Td!'.����Hr��D�Y+��,"�`KܾF�i���`<=�����!e���u4��$�`�wL&�8��֘��u@5��y�g}�$P��'���r��S����9��M��@�u����vmt�]qM�����=����/}�
�ԇi=�¡�']�g)06�쏑�`=���rN�1����%gN���H�t�Hx��q~C��!��:��>@>���C�LӡrS!iN��>B�#�d����s� ��I�P���q� <N��<�y���|���1<�`>��=���7�s�}����{��|Ȧ��}����מ�����w9Jd�����ǉ��f��U�T��30�[�g�rzff'��!v���dn�/~��v�}��G<�҃A��;��C�!��~-��*��B��3��_���(� J��j �*~����آ�
~~l[���O����f��_�����N��?���'��撖Q�W�9;��y���.��a~:{*it�a>��m�]r�W���� a������6B=�F6\���֪�n�H�1n]:�\����U��7��㖞��W�P�*�ڪzb��7)��Q>Φ���ţ�f����*3]#��Ϣd�����T����\�8v-������.^�_0��q��;ӏ���)v�Cv�F����=�叞ŝ�x�]so��L���\��1�ݏ���k��� �z�|���'�gd4���:��Q�O�z-X�ru񉞅A���o����ǐ�o��ᶠ�C�-v�!��`�ƽcr߽��A�Ϣ/�omKO���DV�Z<|���ܹ����=�xI����w���*���%ҽ�_(��^�@��.��������o���G��Bs��\4a�������� �Wʕn�1��5^ �u��=S�O������+��Y�fL��O���V�v�9������i���FK*ޞC޹w��{�Q�|7ʹ���o�"�I�W�qɋ7��u4.��^.Bo��S2��
�>WF6,���[�[ͭ����f{u�]u��]u��Y�]u�]~���]u�^߯������~�~�뮺��u�]zu�]u���������]u㮺뮾:�u�{u�]u�_���뮺뮿]g]u�]u�]u��]u�]q�]zu�]u��]u׷G]u�]u��]u׷]u�_u׎�뮺���]x뮺뮿u�]u�]~���:�~s��7�~s��v�\X��9��{��L��g[@�{á���������phk^bR�[Ł��X���J
5#�{ė�d�2Af2���Sr{6n㔉R�*q�U�-[�'�wͅ�<T3z./���e�p<���yyA�rw�x�Y�5�a�y�TFԫ�	��h) e� �G����5�����5�y����S.��wi���FE-�&PuP�h�7���,b��oRɡ'^׽�u����=��u���!�(��[=�gk�b�]<�nwp{�p{�X�@{uC�^\�����ʗ�;�³Ȭ�g�87skj��0,�/Y4��3	�U�1l�|=�`Ǥ�^��vޜ���D担C2��XYtcF�E�^-p�+d�qr����z��39��������M�=�.���`�g�]]]MѶ���.�����n{x�.�=+O�9���3�n�!+���J$OOW&ٴעL���n�l~�����e;��:�]��o� ��'\�߾��L��Y�*�goq(ӛ�Q�4���abA�,Fe��v�ﰪE^ͧ[ߖ�����-I�k�
���BȸZv��I�����C�!Z0=��3֏D\F���fwwy��Z�u�{u�]u�tu�]u��Y�]zu�^:뮺뮿Y�]u������z~�_�ק]u�]q��]u׷]u�Ƿ������]u�^�u�]|u�^:뮺��G]u㮺뮺�u�]u�_����]u�]u��u�]u�uקG]u�㮼u�]u�\u�^�u�]{u�]u��]u��]u�\u�^:뮺��^����1�E�;�f�>z�[1.�l�,��٘�q�]!�?��s(D�s��z���]��AR#
%f�#t���6���Ԫӥ�Ľ�N�wq�"B�T��f�arw!�3���;�c���y�1�5�P!=C�Fg�d���|���I���}��i>he�|@af�6��(�\K�R��-�Z� ʔ�f�ͻA��r� �qE��9��|�=Hy�N�.��Xp�K��`}�|DO+c�oHF����k�O5�!&A���^BA0�&i!t�ӄiHƇ�L�IG�JS$�vV����,i�cƱ�$�g�0���#u�%����Z���� r*��t�-��7cZp����f���51�t�Z]܎�ԷS�tNBp�?}����\�D��y,�λ珨x�őAEdQD7{��#�B���Ӻ�˔��+�D�>�����ȭ2��t\ہ}�//��� ��_w�_i�F���?���q��_r�5��<9)aw�ᜳU��Ps3�Z.��;U������-��<�3k�G�o�0>���:��y	H��^�^�8���Y�N1�6I�!�Z҂���tJ����P�0&��-&V����Zve�̌VUD7m|�g�輋g}��6>x^ٍg������4��f
�8P��Ⰷ��V�m�s[H`o Ն'֭�&iG"r4=�˷�0L>��{��9��8�(N�1՟}ۚ�sy�X������}�}���1W=}�G�Vϻ6����~>?]u��]uױ�Y�]u�]~���]uק]u��㣮�����������u��]u��G]u�]|u�_�߯���u�]u��]u��]u׷]u�_u׎�뮺����]u�]u��::뮺뮺룮�뮺��Y��]u��뮺뮺�u׎�뮺�뮺�뮺�ۮ�믎��N�뮺�ݿA��7z|��WRa<��-;�2(�^��"az[�$�]$b+���>���w����~^��\��'���5��m�վ�������mc/^nՙ�;��A����.0zr=��{u�;Z�᷹v�>�׋.s��Xb�)�y��ϳ��zEx@�{8kk��ۀ��x���wX3�5���DH8E�'pCT��C��O��=���'��3��O��{ϧ���V�.��5W��ȏ,q�<�zJ;�+:lUS��������1��|qt��;���W�l��<&s��:�=U��y͛��}Y��Ͼ�w�{�X̝1�	�����]ֿ{bҾG��<D��a����m��z��>�U��C,�Q>�&�x�Y+�׍{��C�f�z=m��{<���t#/�e��E���﴾�z�ς�/�f�O�pg�����g�}�ظ��^�7�����w��{��j�H$�9���뚳{|�X0*(�� �Z}!���wb~ɻ��������4^8�|��W�6���Eܼ��z�z=e��k/}4P3u�E�;��ɟ9n��^���]��Q�=x=} o�:����$�T;�^6���G��u��w3��6�;|�g�i�DZY�rr��n���+�u��������㮺�:�u�]u�_�뮺�ۮ�믎�κ���������~�]u��뮽��:뮺���_��u�κ뮺뎺�Ӯ�뮾:뮽�뮽:뮺뎺��]u�]u��뮺뮺�u�zu�]u�~�:뮺뮎�뮺뮿]g]u�]u�㮼u�]u�\u�^�u�]{u�]u�;�yw\ם��:����|Ǚ��˖����C�Fv�h���=��&�b�8|��G`w�*9�rn�H��X%�"�CǗE��_�˥�E=�6^�uzz�]�7i�=�Kv���G����Ǳ����}r�}����btwa��Ϙ��XO�
,a�ٜ��tnwww��FG#�W�g���GC��_������v�5�5�\?� ��}��p������3��,^�pi�����w�}���}3f�wg?/\O|����SY�%��\�Ƹ��}9�y��{�4mJ�QvԦ�w��/N�$]��W>O	}:Ε�{����{��s�e������p��{�h�ٗ�yw���û���K!-眜��~3��}|�=��}z"�a��{�G<��$�Z=�&�ֳwHګ�-��S�u�o��bp!��Z�lK���5����'ܡ�����N�t�VF)rj��X�U@�m���}D<����yƭ�B��K��w����`ϧ.:@���g+��G2�u}wv2�9L��:#;��e�N�)�o��r}#���W�"�B�t�����_xs���_������]uק]u�]q��]u�_u�^�u׎�����q�?_��뮺㮺��뮼u�u��������㣮�뮺��Y�]u�]q�]zu�]u��]u׷]uק]u�]q�]x뮺뮿u׎�뮺�����]u�\u�u�]u�]~�:뮺뮺룮��u�u�㮼u�]u�\u�^��y��<�S*������3^ok��������q�#�#�t�=�7ܤg���~��|T�������Z��س�l}����ג�.�kf�:��/�KElh�z�72�u/T���[QU*A`�eF�Nju������v�fZ���l̃���{����	˱�>T�Zb�׍�U{u4�d��r�����òf��)1&x{}g�,<0�1(���Щi�w�cc�#�C�Y��0`��d��!��9ͽ����<ے�w�d�#d��A�v�������+�G����LsIYG py����zgt�]!�4&8�F]�ai}W(^V��O��w3�׫y<٩�����)��#{���{�&��Q7//{g�x8�`�9<KU����$4_�] y���rg�7浞�R<�W�>��D�4	;���߷۔�����|��5w=�=RC�0�Tf���y�x�j^雛ݤ��^4��o<z��s�򗯼���w��j�s�W|����]�H�;������K�P8wM9�W�9�1�۹�^������ږiز����t#�ּ{�ߦ�ً��S���'ʱ������뮺�a�]u׷]u�_u�]u�uק]uק]~�_�����~�]u�_����]u��]u�����������뮺뮺�tu�]u�]~:��]u�]u�]u��]u׷]u�_u�]{u�]u��]u׷]u�_{u�]u��]u��]u�\u�u�]u�]~�:뮺뮺룮�뮺���zw��Ͻ�r����S�އNG:R��Dgc3H�{\3[1�Z��Y�jr�.�C��Hk>ǧ;�pB�3�>�|C�e�=^��=�i]Ulf�'=H��y#ʾ�`�Њ*�&�'l�O-Mxߐ��_U�g�g}���[�rgOa}��4=3=� Ҽ{���9���M������0{�����{���p�Z�j!�ٵo���ܳ�s��^G�t�g���N�����zb��ogv%۾����L~¥B�'�x�f�fwٯ �鋲���珽���]�q�t�h��=�g�GyLf��}}�U�"f��zǧ�y{(Ͼ�=��M�;�P��dXJ��H��p���2��ݡW��Ouz8<��{KX��f�*Q���횲^�R~�xw�뭸��8mk��
D���Mn�1f��l� �{8)sJ�v��6�֟��{�xꢵO�z����y⏲sg�;�||�R���qo;40{(G^y���������W��ǖl�K�'��lA�/u>[=؏S���F�q�z��0_3h�|���w*�gdЫ��<��Cn��BU�������ٷ�3��9ݧ1o|_��,Ef�é\.֌�����ߵ���Q�4�W�R����އ�yxv��6�1����}���� <�X�b �"k7��.��&݈E����}�c|������[���~@{��S�ya�&��CD]�(/�V��Xtۡ���]�[<�>����_٣3�>�1u���]��Ułf��:�^�A(՝Ȏ��x�Ȍ�k'�{YH��q��٘���{�u�0���W��׈���ۡr��/w;��1��_z�rݛ}�Y�~�q���)�x�@x=f�Fl;��;��r�Az�|�"O���=�+�˻�&��B�{
78�MEz�n�#���~�{��w
Y�,A���e�������el枓���}&n�a?g[�<x�#�W� �F�4�{~ύ-A�6�Ik�B3����D�#���,��t����gkZ�m�&�;��A���C����B�p�ObY8�z�w���L㺼.u�������}�}��Y���-��o{�,�ٞ�Ȝ=�a���r�
og�|����pɅ�>�|DNJ�}��|w'v����%��,y�4��wy`���cG�hckx���1�w���>�	�����-m�F�;�^3o'��g��H��^^��;�#���W��`%���n��!jO63�u��z&%Ώ��/@�^>�aF���qվE�.����J���b��^utܴ]��".q�ӳ�3�ݸG�~zâ�'o#��a|Q�I���{����F�@�.FF�wR�s�<k���@b*P��/�3a�>y{D�a�h�%د�w��r����n�sUPP��>w�nB� �˻k��sݛ��V���3�jʷ\�\���G�[�Onfaވ.��٠M^���s��x�A��a��8ȶ�jG�a��������Ԋ;�Ǘ����G����4�X`�J�p:E�=�[�-���]�o;��ۡ��E`���yz�0� �����C=�ח��9��y��ly/��Uyތ�n�T��s�1Y��['�خ,���ܢ��cj��u���EF��#@�bo{���^�K��Շ�b�� �q��|Z�zZ��b	�۶�y�f�!W����>���p6ǽ�v�n��V���j��z��C��ۗa�*9fq#	�{���jFv��C�S�C��:��=<;�r>#���^@0az��<B[L5��r��w|j$ӾA�yA�{�
��U�Ɂ��Z�7bu��:�	�=Wo���Qgxn�QS|��g�����z�Eq����M`m 0J�W���wn� ?vo���J��/i��#x+���V{����p�����_*Q�����L�yW��M\��w�R��'-�f��~/c�낗Nz峮�����sA��Vt㷀V�����ؗ�m�.��^�o��<	]2m�`<Om<f�w�JnxJQ�Z�O5�����z�浻�^ھ����|��Z�5y���Ű.���7�Ky�Ay1q�7m92�8�p����1�|6e���⴬�h�y�x��N\�}`��w,�غ1#IK5zn4G����<�量:�����h��{B�r��e�`���}��,3g��Թ.{����V�[�O��_L�\4��s��7s�^��ќ�݌�Ǝ�c���g��Y��_J9�VsY6ޘ:{>�<=�w��xa�A]VYW��N���Ӯ5`�{���Ͽo�<�����Q U��_����~�����袷�~���?a��y�A���0D:$��n�QЭ�jy�<J� _%�9�j֑q�.�k�#��LU�p���� C��uE���Wz���Iu|-�/�,jkll�`]�Z�7X�O�x�	���B�|.�� �ز�L��h�����e-�,��s,���y���a٪  ����q�����xN�9�q����{U�5�!V�*���.�)
�hJ��5ԅpRYXX��dƆ��H44�k�-n�{lL͗/oo8;>]=-���V��[�V��y��]c�0������@=0B�ж��U�W7jQT��mb�r�ƙ�4К�֐�6���7˼eY��|��w[�9�.�m�YX�"�+�a4�-U*�Ҭ�jb�K�)��U������_V�=R@���c;Pf��1f��d��;u^�����w��w�+�j�uv��\�<pvH۫b�.�Ėm��r"���ۭnN�c��<g��kɮ��'NӰ�3���$Zv2d-��:۳v����G���W�6Xا��N[mC�tݻfIz���cH^� s�#X��/Z�,bm+Vj��k�a���ZF�Y�"�f;�����۬�v؉��޺z�HG�n+�MrH������&����F&��jVZ����mk��`��wG�c��e/N�:78��df8s�7+��8:�c3�Vw	�[8Gn��.[	�:�\QV�
Z��(#.+�B�W�
�&���m,rk=�Y�c��y����3�s�瞺T����2�S6�&ζ1`ʺP�&�n Uk�"F8Q��R�mu�qftr܍�.rL�Ia��������9��]p�r�],ti��ո#�z��㊗.���Rj�����&�d���<��ʹ�Y3��%�z��9�(���Q�{]��g������������;K*�7/U�Y5.��Y�:���i�V�:��aƻu��֬�5��k�:��u��Ȫl� ��yN]=�;a�p���d����a-�����m��yX�i���W��u�^�#kk�س۠��k�B�WWf%��̶��4�Sń4�.��Z�Q��f��qЦ^۹yÓan���o[�Tq��{rc��;��k�M;��R��=���l��wT�b�5XX6�n��tv��V�$f��R�Q�h�0��jY9!x�eHQ��]���%� .;uy��r�uOsᴚ��]sK��X�=���Q��g�v)sfb�KokKj�h�4獺�{e.���F��\JL0،F�)�q���Wa8Mq1Y�q͗��k�:떘#oD<�t/</\�,c�gt�U;����Rw.�����5�.�d7�d
�n#��>޵�gs�t�lk�y�=5+��z�vy���t���.&xj;�Yx�Ѽ���ױ����N�U�$�y�MY�T)b���hF�-�J;p�wa�K�;sRV*��f黌�[�\����W�Pceˇ�M��\�Yv�v�B{qq�6M�`�ь!2���Yaԣ�5�j��� �
nx�&Y��643��ε�0�)�l2��З^���Үs�m���`��Ў\3����e \\ʈU:U4
����\{GGN�]�o �l����e:�a7Z0�λ[,����f`� �M1e�Ŗ4���w]t�<���.�':س.&k��#�B�-�$3Yf�+˳��dV��i��gTn[͎�8������u6$y:�E���#a6���[�na���F�m���==��m�nJA��XL�`A��Y�v�
�� ���h6�c�A �Z@�JB��jM �m�����r�'v�ڝ��k��Ƹ�9�ą���D1C��Q9�	�Wk0�2ʕb�u�yuA�lth���Ŋ�⸖�Q冸.�J�]���aƯG=эՏ<^5vT�8�Xs��eݫR字��XP��g�;V�X5��5k`E�A��qH�];i2j� ��N�F�dΡ���se.��OauPr]�Nw]�k�NՈ5<�;vs�qk�[Y�:�Gd�v��U[
f8kZK�Ie�F��D�xB.�b����gA��ut
䘊�9�K9�4����u�b8:1m!��g$�mԈ�tc�.�c ڹ;z�x��]J���SB�#��ڼ;n�(����Q4�Y�ǅ��J�,9Κ7db�-:W]�su�v�T�3�N�N���T��.r�"����&,H���L�׀fl(�e45ֆья=YZ�n!5��»^4�8��]q��(3�^�Z�\�`��r�-�죹s`cA���Y�h��ك&�r۱ź 5�2��$�n4�i��Mܽ�V��[��5"u]oi|[�d��m)���k��0uˌwn����a�KFg:d��M�ycW ��cVhO��L;o	����j�W�T,�R�s�4"#�qZ&堗II�*�k@�X�+m�M�L��[�ٛ-G9Y���)��Υ�f�nN�p���uт���J*�[����B��C;�6��]r�T�]FY��Pf����U�RŦ�6��#��������L�vJ.��k4�Dj��ض�X� C�i}�O\n�Ϯ�nnE�a8}i��2�<��5���·���qb��T�[Zm��^�,��T���N��ۮ��8�\\�C2<n�k���n8�7��Ͳ�{'gZ۔�������n\E)��-5�&��Ԍ5+4.5��e����c�!�T��̇gw[=;im)n�K�ݮ9Î7B�G2C͹�̸"Z�u&�W6&c4&x#�l��"��睱��Ӛ�]!��Da��G&�:�q)U���n/\�tw4�J�K<�rx9��³��[C���=j���D�cMg��Ũ��r�u�1��
ʧ0`M`$�V�Y��j[s�s��UԽ�<O+�CjW��0��dv�.�x xWm״��	�f�uny:]�W�����s]lj�u��=�\痟k���iwxiݻ�;7ɳ��u�W����n��:��ɺ���Md��1Z6����z��u�7��S�V����e�$^�ʅm�k��=7��x7f�ݕn ��{VD�kX�"�M*b�8m��*�pƓ	��'��^�GRɱӷl�E�7.9ۭ�͸�z�^���%&��K���Gx���m�<l'aݎ�zUq��n��v{b��Ű�V��z6�\Z�r���5q�n�W<�mSg��v�}mn;�O:v���e[cEu��f�
6�dr�2E�V�!����e����>�XM�5�/X�ݩz��Y�kv^jE�b�A��jXT�����޸��r��ű�U�J�ʅػ����l����cqY�p���!+y���lik ��g���k�n��ov7��k$�t�;M5�����L���hѻQ���}��H�n�(=mϩf�A�$�Vl�%�%ٙzg�H6r@���,�oR���SGA��e!vx�; m��v�V"Gl�CXk�lu�8�[d�4�سpBm��m��͝�Vz����x�m�f�nli%���" ǜ@qp�qc��a��;	���NN�ڑqE��Q��bȉΝ�	����Lvگ�W��LR�ݢ������Sv�&��z���70��X��(<��k�[n�[T�itxc��sG)�CC���u.�Wa�cf���fu�Y�)^N����ș�d��Z�M��c*���q����d*ٝ��T��:a=�X� 2^n1z�=��|V��{�K7;��4� ���V�ѥrd�^��U�n�3T��r��\5K�f�sM,���V��nl�%��z�r�Yl�xK�ͬ�K�nnɩKdzqݥ���f�E�����,y6�.�[�YV��>�v�庻�F�^D���h�.�>]���:��n�r��f�td�nxt�#�I.���.�0��1es-��bg!P�i���Q�g�ck���=l�<^ͅ�M�Y���70��h�֝�GJ[��F4��]�x�&��u�Xh����6���Y��	L�6����H	L��BX�j���&�$�(J�';ҥ�o:�z���:�Kz��˻q<ڠ��qs�����E�&�u�f7<X�����g�q�I�4��CE��3\\���8),
�\Y�4�Kv���-ί!�:��m��鷋�#��x;Y^�{gi���,yF��n�'4c��
�f4n����FU�G�y���ʒ2�[�|��#Y���8���gB�ғk����a����(v*f%iw��)Y|�8���Kc�oyXY��acΪ����њU�����cf���vk��]liUNe���{���8=\j�s\\��\�X�y�$�]��g��mm��\ڼ�{�b�]��=�����Ni5�E �n��F�i���c��Gn�^'�/���ȍ���Z=t�U[2���:�:�,)tr�+V;�	di\���+�]� �7��m���tS�约����������;�I���Y"�����#�X{=-w?����qeNS�l.�9���j=
�[S�f���n����vx�1sB���`���R�����T�;����x��9P�&RlL�+i-R<滗�W�9��&{l]�!��>�m�hp���g�5�fi�V�K*r2��9s�Mf��ͷP�$_
*@�(M��s%��9�]���­�΂Z���O^o;YKk|V���-tm3ͥ�y��R�τz~��<�n�8��p!��,e&���[��a�_�,F7������V���B��U�;�[.�4�c�L�U�2���<��J���/�l�-ؙ%j�ݻ���V�,y�]���zxGle�7h�[�3
���=��r8kkS�붣Z����S���+�:�@��C���Fi�r보Mz<1\�K���cL�-��'ע@��JF� I)%
�$Tc���ruϝ���;~���=���]vlٳf�T�Q��[TQ�s�� ��~ީ�{c[��L�Ȼ�0/1 �)-	bm��c -k$��PV, ��������~?_��������C�XF)r� $u�*LH�(#�
�E+LJ��� �A Rb�`�'{a5$Rk1$*�ED�&1s,"5 ̢�K�5��W:�
���XE�^RL~I4N��w��(����2�m�7�lV �{~>�<����}}{{{{{{�ATYDzd8���X�*�*����dȬ4�-�2�`�EZ�k�ŋ䄷P��J5�C�������Ж�N�/ ���g4�Wn��
W3��N�����믯ooooo�y��Ä��^nGǃ������x;-,��^����DHZYa(��1�
���.	��}�;��;��'��f��'']���V���`N=jQHF*��ÉNI�e��SVO-�`�EAA$X���u���������������������t�Q���(���iO�Ɉ�LLE��j�#A+Xѩe�̱�V��D�RSc1YD$@b�})ENN�rF ���R"H�[�ބ^��B'�%\���JLǥ#T�j����-��S���eVE�E2�Vf�X���V+�ӻ��<ؗ%]���������E) 2c2aN$A��N(`em��7��Yq��XW�-/"dR
8�O�$�a�x^6�91��������g]E�)���J��;U:�<�\ny�)Mv�s=��ri��9�q)�Ķ�ۭ·,�-���e;&],]+�'P�%�L�����;n`x����}����Цb㙹띴�s=�$y��[gIX �(�n��-�.�^Ku=vݺ�x�WfD�j:x��1:vydN����B�G6ƏnӐ^7��0"x�b٭ЈՆ�Q����Y��v��*&)wr�H`"ȷqs�;@1�1(q���V����Uܦ����99��'=qWn✢�і����ŉ�����8tR(l���n,�=�x�ùǊ�pv�a�:ٹ,cU�3��|�����r�x�=L�爷��ι5������jD�,M�r�Ck�,1a��ʝn:�9܁�]۠�]+F���+�l-u�c,��j�v��G]�s�`x���|�+��q@����,+�UՈ�S�-g��۵�1A[�}:m�n��)�����D%#s+<�j��8�KS6퓱٬M���5R��4"Y�i��	�1 �X��;6�u�#����q�rPp����n9-�$㗮�]uɱt1ɧ������	��jmm�Y�F�rE����\��P뇎-6�un��9���g���eM-���J�bpU�x�>G��)�nש��N8������H�v���RG���6��8+<�ƝeEYr�р�c��o)�c.0�KM��K�@1��wj�y^3v��&Gk%Z��������
��%���.��z�c�ll�`�ѻh]�ulN��f�FJfCm�Q�=xŵI�qb뱫1��[Xl�б�Ѯ�H�/Z9�#�s�n	�-c )�e��Uj3<��S�c9f�u��w=�;>���zQ7��P;s�ݧ��8%�GRl�����Ǟ���ǹ-��<�b6��)���s|$�M��]�^5�S���"@4��J�"�YB^"���RYe��jB�����jRPZ��4JX��m��[��oV�-a�h����#ר���Ic�mD��,	F�+[�Z����	am�,���N���i�A�R�`Ճh��VX�Ԅ��k,�ekb�VTZ	(
ą!�iT����_�����Gy?���O�1
��$Nk�*�%��kt�J`g�qS%�qU߼u (tj��>Ű2en�����H��%1�$o�$|�"���-O4�|��-�@.���ˁg���|��t�{b_�!�bF��M2YSN�
w(C
��w/f��nKJ��ǵ�`�/��ͱ��w�}�៞�s�rM6P.f.aL��t΁$y��<��ԅ���C�� �^|"	c�y�e�9���w"�܄O]K�2��{��\�^���M�r�%xC��7kA�1ٟA�7���A �{���`�z>�D�X`�{�)�m�s�~�O'�i0���s��b��X��{0��Y���;�QU��G�^br�;*��p��~P�U�>����0�C�S��d%�Y=2
$ ĆĽQ�Aݏ;)���ǂX�V+��*�{pA7|q!w2�ֲ�\=��lC����>>ʣ�w{RA��|����<m�dlP���#�����^�%�	F��RŁ�e���9�	��*� �*^�1,2.K��8����?T�}U��_K��0cg��jv.zb/��5�9��q?;q����-�VO5�k����ѩ�nksu��N�N	�ES�#۫]�"@����*��b$����1�e@���췆+��@9�m3�>r��)����&����ƛ�{�qè��:t�{�ξ�χ������6���������ǀ'?,_�;ت���������3��*�}��W��wٳ��V�wdrM=�'qޞiS���s`CI�H�Q��HU��y���"}�5��1�����<E]�Es
��iy^Myd�#5%N�ϓ!�oj� �NףТ<�j�ڲI�S�H^��jF!��Ƌl^�yX����橓O��X�5�<I;쀨f�Й,^�p��)��c��[�����6�k�T�ٰ�7D�8kraݮ��z�v�\�F�%�;JM�ￅ�r��i��X�։$�o���1{�V�<?���p `�͆]3�)��������+zv4�H���1�YlD���A^�1�}�Mz7�<sb�x�yH��tY8��wpw
�6�0$4{� ?|-Ηߍ���;�*��؆��[j�*$=�/[��D��9�*��^}��I �e�2 ��10�H;�9Yi^ב5���Q�緻X���פ쌼�����_�q27��?��ۊ�	���ޏ��>���9\/��D)��;�/3��S��	�P8�b�� �$/!�������eeX��7� �����}>-�o�;���9���1D2�m�ch6d�#R+�u�n�l�k�cZ�!6���=�Ħswd�j� no�4�;��|}� �EW�]>^=s�/h��r4����ĒbRrXb�R�o6���"�8�4c�O//O��F�یœd�8�52p}�p߿1m�)����=�~�Sm#���4f-�/����$��k�͹�x&��YhD�<��i�91
E	^����OP���1P�&4�C�b<���|���n{��^��mM��"Lo�'�p �zc׆���Eb� c�"��)�Ƌ�1����W�)���ߴy��s�9������,q����r��ߖ��Љ����"����k�����t���i$葓�w�o�e�\$ Њ��j�Mn�[�xR\G(jYFTl��R.�e���'�,��#X�饼]\��$Hi��	Ycu��:2nR%�Z{iQ��d/]���netu�Y��~���|b5�%+���vҲ�:�3ժ}�cKOS�ช�v7st<���Y�]��t�Ů:�Wf�껉��J��LR\��T���K׌%ʝ���G�P��jm����Tp�����t,�&�Y��n \���<����Ϩ�L<C��������s]��I:��8��1����PP�`�}�x���:�E���XJZ��;���{E���ҕgM2�y��H�����@�������ס.`�x�����r���+���+kg^rG������QbA��>�ɽX֞!C����O�הN������=�?�2Am؈$��N��P���x&n��.��xV*�
u�z��$���)��I�Tӑ�c�1���v0K{�dzn�r�"}���qk��;�`��m�uc�P\Dv
�$�ں【Pg�~=�oX]�	���_��؂I���z978rTo�A����+_o�)&Zl	�?�|?#�`���-��/Е�Q`���^�0��v��OU����x{�['����?G�o=��{�w�u�|����sw,	�L�]�� ���$�e��<���i�<M6"�B.f��;W	����B��>u��G�|$��zc4���`��+�5���&\^��^K���1}�D�TK&MlP��0E%^��+>Y�q��		]�`�(�-��	C(��ո�
�<Sk;�P�- ���}��	�{� ��U��O�L�C�bRy���|Yb㵫Y;P�b�ś<j�5լ�c�]������-t/-�s"�[�%�^4H2���De�~�߆�ypxz��&S)���(�뷪=fU>y��H�=��dȟz��KZ���۟N��;B
q;�:��37W�H���w͢>K)��� �����O� �zy._1=R���;~Ig�*6��箒�ɨ��c�o}����މ{�d���pN���r��N.P=N:�������)��y����ϛߑ���<�?���.D"�h�3�;解hN����Y�C�WnA�3|n��j�� ���vn��q��TN4���R�i��d��q���_ѳ��h�5A �h�� ?o����x4�A<����g[c���\0��t2&-2<s]]��k[�����������������%�DcJ���~Y7v������A9~�D��%�CЌ܂�:������|�cը��f�>�A;`T�$�S?��Ab��vAw���m���5�s�Aܐi��y3G�mߖ7���l ����G�6�|�#��I�z;-B�p�wxP �ǍPͷ�s_i���C�,[2�%�C��7�<�#��U��Q���W���[-��0׼��7<w���bZ����\W��h��ˍ�y0m�ľEU��>� �06��RT�E"�K)��<�yϗ���q��\�Đ�����~w�G�喭�f��^A4S$^e��I�\l>�[Oк��o��*��Ŵq]��u���M���<Uۗ�N&��ZlfQ���_��d,y7~|�I ߲ �b�/y@���9�c�h�C�00 ���A��g�)�_�L;�@��ϓl�Vf�]�/MMq��$�Ff�&Ab�(����y��=����IN�%"@�;�b(�)b7QRH�t�{\� ���N-�jc6���s��È^s�u� ��mCZ��H�^� �I5�y�ד�LV1 ��G��
�w���	�V
5PX�{{.���,'�Y�!�I*�ǝ�ڣ�d�=O��g����6�?A�Oi|i�ETKY�T@�iG�����%�n'�vU�ǳ��ˌ�%/bÆb@isS߿�p�޹���\pl�p=UY��E�.;8�6��kǦ�أǉF��[�V�\k�֧ϵGc�IW4�g�:�|�[�h컗;V���gU�]�+jW%ĳ1Il�K��&�� S��.���8�h�%1e�*t�w]6�k4����ۣ�F'��U�:��x�p`�j7C�+=q�ABf�W`ō�\��L��(�N5r�m#'b��zJ�β��R&���b׆��ET�����sY' �s!���T��	.׀�̭���J��
�V\YxۡD�V�BF��T ��S�&=�Y��0~ǂC�9�A&X�|�D"7�vf�G�\k������x���� )��si�b=��	�ۼ���\ |V�8oTc��x&j�F�P�#w�;�=o���{�߳� ����"��;�C:#���ȃ
��/LnI�w0SD5�E ������ >��o1/�z�]��E�@$��<I7ş}q�*�J]�p�)��&J��[t�c���x��B%S�fr��f���r2���~�]m.���}��{�ri��q���7넦�b���� ��w�������' �s"���`�5�f&G����9q�ء���\����?x=�<#]�>�~e��o�Fy�{ߜ��g�dy��C����$�,�޻A�z V{�>�Y@S��o�s�KH����_��� i�~�F�!�b��s�nnW�-{0��{�	O���A���ݵ���}^���휲$ Dמ �Y�ŷ���ϫ�3��L=�4�/��}�	FC��p2�_�d���ߤ�b�~mf0
�����lo�V��=��I��v?L��$q8�u�9�u��_9�Лڷ��1�QyX[�}�f�o�>�����p��|�}�;�D���	�~�J�����=����M{"��bZ�C���n�ޥe��1�̭wU*�JX�HƉ ����=���Co�{'�{;�AAɀ�D4w�ty�=�^�J�('�>u�}�w�8މ#�/�!�sڟ]ќ�=����+�X�0���P��u�a7��f]���ǳ���.��o5�����A�0qv[��QقƔ����ˍq�����ݡy�]�����0���@�����w�,������*�Ʊ-�읒�;����>�O��w!%�A�9���6>�W��>99L��J�9}Nv�-�͇5w��j�gk��6A�3�������b#�{��3q�3�;Ow�{{Nz�~GH3�Fc�+�}�77:l��ǝw�ZT�6����3��|>g"ǼE)��M�:s�.�{�TuW�� 	8�0:������D�;5U�:wIy������S�Ȝ�w��A|�YNg�՞u�6nC=�qv6ز�y�O%�N��Zݡ�H���ܢ{|��(�vhRtcK�R������vFp�x�h�s޳a�x�\D�;ᦁX��K�����;4��rm��ֱ����3w޽���ӻ���g�ځ	o=>]��� ����L��������R��F����>'���@3�=���ٝ���F�;��%�)D��7�s�ὥ��=�J�p;�i7���G`�C��{�k�������.��,��;��Ex�ݞ��v���՞
����{�y�M���u�
1���j/=����<;k��+��a���s�|)�'v�'����}�����1g;�I�U�*O(hA
�1�?0�{o�Q�㿎hVj pL��҇�^_�>��1"��ptw[ԏש%8������D؈��O^u�u�q���θ���ퟃ��__^������)2yˋe��:4��o�E �y�(
�(w�x�ǣ���g�L�q������ٳf�r*r�/.[�\6QnRX[R�>�N�%&X�� 8���j:�p�_�>�g��|qg����rlٳf�G�����$Qd
�F��r�^�m���S���PQ`���<��F},�c9;��{>�NM�6l�7�Z�3��5��^��F��O������B�F�K6�ݷ6�O&O�������}}|{{{{|;��\h����;�h�-$cJJp�,��dX���(�ZR[T��Ogr��ќq�����Ƿ�����|/+�Yd�Z�R5� :����'���aPR1�̬b�[�0F�w��tQ0+G���$�)+&:�
��*��	>�[�䅵:�''"�# �$����YR5�Hy�� �2%cX��mS��e(��@ƃ�6�7��f�Čg$#,HČf ^������Y-<�� ���,��C���`T�`T�<�L�M�s+��z���C�C/~n��|�Y�ON�C�z3�@�0d��� w!�%aD��Oo�J�(��<�~>�ܾ���u��(���5*w����EP3�Nu��~������a�rz��>g_���u�qNs�^���������s����H�C���̈́� �����IY	
C���	acb�f�z�滇0`4I�ş%>=�XY���v�e���m軟>�yM0= ��#-�9��~~Z黗]�ֳ�'���ߝ��G�>���R}޷��1�X+����C�Hu��������"�u��1���-�������XS�|?{�&��9;���DtAi�" �����[|��O��	�k�1!RE������8��bL@�w_��u���I�^��9s�}f` ��p�a$0]��%�+s1����?w�hd-��e�z��׌�2
X���Γ�{��t{<��!�;`VT
����~����q��
A�������^��<��!�Pg,��.��'�8,�p��o�O̘!P��!�nw������2q1�}뛩a�@��B�;9�`�g�Ty�󝧗�&�p���{V���_O�;��:|Hó(
��;��(��1��k�Ti�)�K�?}|��7�|�0ﾋ����0�3��aBе� ��{G�K׼���s+�6X���vj�+(�R�O���5�s߾����㞠%'������g~�p;����N0'�A��tr�G�����޿O'I����YX݆���uuv �X�z:���R����n�(�$���/	��Q4��-��/ցӉ%ə �`{�ٯL%lHT�#����g�!>�'{�����{
T�����q��ﭣr!��0I�~�0�J�iߟ��t��]�vE%��ؼ@��`�Y�f�yێ�8�^g��=J��S��a{����b :�0@2�Np!}�ܪv{���?0mj��D��o��
w@��O]3 %)��[��@I(�%���~������-���Y�0H�&^�q�@ ��iyʇwuH��ֲWW�=�Ve����� 	&TΙ�_�N�qގ��P�d:;p��H^� ��\a�r
	 �(�Il=�ي"�t���!�nt+*�{h�Ml�Av�;)�2wHo��)�u�������i*�=�@����-��7<��QtxY�Sy`V{<��t���T7V� �O��y��{뷯_2��NШ~�1��1#�,e3�~;��r�mKpW]ݳm�mv������G��rs����c�6a��7��ڞ�ۡ���0� ��"���M����C���InS;�xXy��k�XB��5Ѷ�[aL���)]e���2>/oko[{��L7&�n��C�,.Ƹ(Y��R�3�.�q�4G�q�zvz� ]������풓������.���h׵�z�i�W����nV�n�u)he�f��[�����
�HǍg�g��*YݑwJ��T���;�YwD�:���3�7�[Nz�@&�R'�~\xL��n�=�0��G�AO���HƐ�A=�c��)��Ґ�w ǋe R�w^��R�k;��}��*�n��i���E���� Q����Uy�l?J�-�D�oV�N�S$H&+Ѹ)��3}��@<�-��ұ� �s��$Ϙ;(9P����-�{�<���nN8�����ę �:΋�יJE�l�[�qq�=�������dH��۩y�P�"�iq�@:%�5x�k`n��sM-�  �� .�I����~�L��w�H�x ���]^C�k���xyŢ�'#��^
P�.���'v���f.squһL.�jc$K�����A�#,�:ޡd#PA"s��蔐.�y'}���q7`k.��,% RKm�T�9�����4���<� "v�[��^fg��6#a�;3���yb���u�2��ft�ۙ��⅏D����i���������γ�3����0�#�_����C�_&s�����>J)k8
��f��^�JC6��'��tH7`��^�t�$�@�yi�3�@,�}q����U�gw+퇔I �	{��@C�^u��ESKZ��GD7�Ɛ��[��:h� 0 F	I ��̲HE�Ҙ�W���>vq���cf*�A��* ��`U���̫d2˽�S1���˷�4N�M��y�Y�$���(���ϙ~6%41]Ѿ��]s�A����vg���m�<�t�l(l�њA�[61-Ơ������@R<�x.7��$�Y��,�$�m�qe�����;���ܭ�SC�K�I ���{����^b�@H=Q6c%�`��g,�\rs{�ͪ���BL�	"^8! 3��tq����ϓ��ꬆ�7U@4^��8���1��h$�WD��&R�|1H���j/�*�XF��,o��_���^U�b�,���y�����/d؝1����h�Ҧ&����"H��Q`Bѱ�?�vx��0�3J���g[כ����c������-���-)K�S�	��:%��I���{G��X|�KaX��e"Ɍ3�t�̪����wK���ꗠ2R]�y�h��vJr�<��f��Ҥ���s�!����;.v��	 j-�@H�id���XM˸ˁ)	���;�O�����=��S�%��D����ۊ2����u��S�x�I	D�xf�9P��]��e�z��G̀G�t&b�;ݒ�U���E�9O2Ӭ���b[��"ٹ��\�(wJ��V��/$7��a�Ǜx�=g�r���,i���A ���.ŚI�����Q�q�+]׏,b�@H=0�;��X�5~�@ �s�{�=V����7}�6�gp+�ٸ�C�cM���A"�]z;�݁� X;��,@��2@ d�u�I�����)�@ׅ���~�w�}�f���Ե2ِ�R���z�/�BI�{�/b����ǟ��a��S鶹A1*�q���?&�,��;�Y���de)�����v��hʏ��� F$/�2����@ I��&@���ƻ�phe�n�z)���a�]3��l ���pbC�O�:���݂�چ������n�¸:8�t���{�(×�!�{��^I,=Y��-� Jy4�R,���v���Ku�jr��y�.b!�	Wj��0OC��[� ���w�e!��"`sL�հ��cVo�/9J�]�K@ޜ�j�H��̆�=�s��d�O�����L� � �w� �q�4{YC��T��(���QWs�:/>�m&d䂁lj���-K�b{]��#=54[�� K�;(.�Q���i%�7|�
3s{>��2���j ���A��ǜAi�[����<�N![��\b����#2�oV������?����|��\=k��[���!�\-�%�o&�8�ر�3/���'�i� 1g,�Y8�}?oҵ�ѥWIV�j��a)�b�-�6+��Zx�=n�]�Lv!�XlTܗj�i���Ɖ.	3(�K2��lH�6�i�{@+15�	�sj�W�<�V[�-Q���h�KpUF̹��Ԯ���m��[ Q���	҃3\�b-�Ŧx٘�O������]˰�Pr<�q�힎.���v���͵Ojy��.7+t��l�ֳ`}�M�p�6�o	��}��+��j��#>x]bbT�Rf�]2���H�f��0څ��g��_���v�F$	�I�
/c��D��p'_�X}��I󽴣=��-��G�Hh��D
��@�]�@��}Λ� H����r�,�$�I �y���C5�w*�U�n��3v$�oh�����y�IS`ܫ��	vL�דC�A$x�
�?�9�`
��;"X�M7tII����t�'F�͘��o5H�{�9�>3I��� �d��!�����gu����&=�jƹ�+0�B$"	g��e����P)*On����}�zh�����t4{�z���ޔ�� ���
HZ����ě��q����N��Ms�E=��u��tIss���ͦ��
�����~�/�vP](��=�Ȕ�3���� I��$��n)��z{�Hm�����Й��.� i�*:�	b+�\=-���e��g<�}7�3�.-;�9JQٸ��ѫdv����{���fy�0o;��3��?�~�Y0�JD1"@g�?�����3�7�-w� y�]�)�c�a� �����@��;�=P�9���B �@�݉$�L�w�;E��Ŧ�%�%�V.0H �zE�X'��P��� ���6M�t�"��T�"E�ݲ�E?w���a�`Kw� �n�>��t�'F� ����4��ҝ�*���Ud�lam��`o{d I��I":}>�]��o�b�i|֎�b���/;qN��ݝ�n�\rJ\���PX=�{����5��O���nS*�P&~ْO2d  �FL�|WF�獺�����Ȣc�Ng@>��e�w�$Bt�M��A�y2G�Zړ�>�$�a��H�j���d_����K�nƓ��m��;��V��gO�Ouh�Q��n�8� G�2�i� f�g���!T�t��V�.&�����Mμ�Q�+8�WYD��ZS��:��S�@N����U2�x���FZ�Q%|?"~F`!��F`{� �5���b﷦@!��} I�s��(�Cȶk7�\���Ձ�Đ%���2d�kb�{fdy� oǻ`uU6.�MX�8]CC��j;�HC$@�[o^u��v�0,R���L���,c2�� �o1���|��'bo1����5tc�-�ph�Z�fݎѮ�	�T\�c)5Ʋ$���_�˂pa:0݄���#��U6���%9���~CPӊo��f�5�wL�P@C%v�{,H7ۣ��� �"��Z�� (��q�0|��Z�7���:���c ,����ϙ�s<���F&�j˨�@#=~���H�	@��>��͙�,�Cmd�S%�fFf����I/��i>b�.��1�z:q�}�I���$A��i��f�#��:�;8��[7{�ׯ*5��b<?߽U&v�8>|��U���mIw�8���V
�n������b�86L�軂��=:��� B,`�_ḻ��?��$�Hc%%��R���	
N��w��C�߿}وT�!����TX�4�'��`w���[[���̐$�Al�	R[����o_]�]zR@��8:�<p�M�nm���1v�+��]�X��3Et���������[����L�'�
��I$��/�=���O��\0���]/U��O 3[Դ�[���80�
X&�m�&HK,�[d��77�N�	 �#m��,@�����l^ZP�>�9�E70i�Ȯs�<3�(q��@� ���b5��h�K@=;��EA�9S�O~�h_���r()��p9 u���8�� �c0��z�~ލ��������XV�0K�rd�c�-,�FK���c��?)0- �'צt�����ߣ��	��OSH�y����	�;7�,@���k��@�]�� ���t����kiQ��l���(������Ec���\��y����F�<Nj}��^����#t�-o�� �"]f�k�j��ǖ�>�NUVTY��pZO<I���;zG��=����O?y�w�ws�;�x����Q��=���3����۝�e�g��RgƢ}���z�]c<-�!�x�n��)��3ݡ�����vM�G�	���H'����HbӻR�6Eب�S�E��hû����;ݧ���3�r��n�7�o��1j٩>^���	ѯ:|�.E���2����b�j�l�J��v�y��<'��ͰN������[�>~y��㈺�8 ���<���d�se��y<���D[�o����\�݅ a��أ���j�X1�X�t���C!��w.Q��@淐&=:U֮��ۮ��Z��ڎTG>�^<���Aѽ!y���份�ˎ��������/nz��*�2}��o���r{V���v���bś���u�Sڼl�5�o���&(=�7�zk�EЪ����2�Oy�ݙ�O�nkc|F(�wK�6A=�ۤ�=�=� [����`_90�j��w��y����B>�V�[��lM`�Ϲ�Ĕ�\��?j@{����S����R�._��8p#�7�����+�xׂ/��y��0Y'�3@�T��cSϔV�������`�oߌœp�X ��@uk�=��Ӱ���Wm������ot�E�S�X^���خe���΋�^��^{�˺o�#K	(�����@ 0HW�)J	F��j��b�6��b��O'���x���q���������������2��Y�+�UO��kjW�9����XU�e-�	��},e�E��?��������y�9����r���.7�X;t�܊��H��(UZ�mA�h�o-��O'ǌ���~�{~�������ٗ�ɩD=���a��1���1���A���Jr-���C��㯯��?�Ǐ��\q���ï8yB���pX��r3�.������YZ�'����x����]}~8���㇔��^]R	�%J�V[c!a ����SY���&�33�.^���>�g���׎���q������E��Q�X[q9�]u1Uj(HrGӌv$
���m�b������?[�NP��E���թyK�9eL�f穐�'oκR�Q��c�U�-��0Q���-J�m�f#cb���1EX����R�Br�%UQi�==�<	 �0���bK	���l�@$��߃�/���J֗1]f�s��h6h��3nĂ�� ���vA�ܯ!���v��x4�hN�^��Ou�������֮
Z�=<ը���H)m�t���e.뮱mЕ�%���ʒ�a���sk�rs�6���Q���!�B`�غ�4m\�5ul��g%�eB�*m��2���z�e��(a9�)��tEyz�9c1Oc��!!W��kƜ(��f���Ɖڻ0填[��y��nq��s��s#rn]�SK/"]�]a��B9��Y4�[P�iaZ^�Q�A̭r�H���ʫ�2CJX\s�+#�j�q��te�j!.�Ӓ&7�\����m��=4�ڭs��"c;p3D1�����͗^��[e�w�l.\��i����6�ѵ ��/e��UOaj�����m]uΝr�wA&5�vw�:ghV��lƨ:��sKvۉ<�+vj�hbt���*�qͲ�Ji���CR�j�՚����m�&�KX36]6l`��OW��L[gk�lk=���[1(��R\ű�[.��h�ۮ��	�x��/n}u��U�d`̛��/]��K5�������B7����y���B�u�v�؍Gkn_$�u	<�����2mݮ�p��u�L�Ce�\�s\�+B��i�D���[��f�];J[m���5=Tv�5��p���E�n�z'L���E8��7�n�I­�f���a�nr�qZi[MYsx(��KŠ�o<Q�P.�uZ8�86�Z]B��懷i�4��$t��+P�C�aYr\u�[�C@ȕn���{hiɎ���4E�=s���ime.7=��,�&؝�n��ݰ��8u�lH���zk'!�y(6������8K^G�;����h�7K1��Yo�GO�B��V�zɃ��r������U��2���'��m�e�Й�{"� jیܼ𬓂�u��=q���6�q�����A	�F��@aXeXa��C��yR���&��m��'�(Q��I�@	k�=��;ۅ>�D�A�GEaĄj���ƅ�6^�ƛa����V*�;*��Mc�G;1ѩ��d��;�O��s�vpu��݌�����=�
�<�R�V�%�2i�jE�$H�!m�l��4z{T���9H��X�(��]]�$p�r�{��ȼXBv�t#]������y���a6�*��a��[t��u�f�'�Y��ؤ���)�u��q�����/���*�q��٥��~�_��A.���C��>�	,=Y�$K�G�k����qEcQ��GA���L� ��7?��/T�@�����Y~�p q�e��PD���L�����h�H>uw�g�|bH3}�^E��R]� *�Hc$g�e��.�	*�/5��fO�� ��ސ$b����J��8���(<�9������_�� s?:[3ɑ$�7�$�'}�¤f����c��,:z�	&=Հ��$��eX%��H`��$�x2�z���1��{ăMMVnL�XKOg;M@-��j����sSz��N�	�<  ��4#�n�l�'8�m��6^��; ŋoϞ�|&+f���s�t�"ڙ��y膲H�΁�&��/#1�WtL�,�u��CJ,D��b%�9ylo���N6�5\��9:���R!�D��纁*3� ��_�].��Q>��c&�w�<�nN^Z�&�;��"j�5�=lX�y Q���	�O���D�!$C	�P�82�P� 2����~�������G����a�(�^ɬ;ی�o۵E��lq��I�W�1��� �v3�b���A,iz/��^����P�q�,e�&Xk$}� �{�b�."��1��&�&v�j���a���I$�`KJ,@��D��v�񩰰  qSuP&Yzr�Ԋ� !D���q�Oɛ7�E��8�Ѡ E��d���H����A}����$��f"�RI�r��zF�m؂��g��'ge1v���ytj���0Ǹ�I����H1@��H;�r���@���A �f���K
�Y��7t/u�%�"	����l�]�Ò��X;�Ȗ�`#za�P��,ݱ,d>�t �tvY��k��w��ed��j��f"QP��2��\$�%��6�H�>��31'K蒰����~�x?M���
��m��ږ���"���S!���Zp��{4?���E��:�dI�Os:/�/�de�G�
ʄ2� �3׳2E�_k����G}K|�c��Q�OT�9]���B�GE��5��	,X�]y�$�	��f���J���T�{$����b^y瞭.Wxl�:s&I�ANAs`�������rC�DZ�vfN>�e�Gvy�s���4��z�s�Lmƹq��k*�9�/�q�ٴ�q^����v��a������)�ћׯ��[��,A�CY�g@	$��u�I	$�H��_k�o���$lz �AvI��e��R%�NV�~��1@��tԁ Q^~	��|gbͼ�	,A"�� I �Y���@'�����h6��]�u�AA�t��C�Ѭ@4T1�� ;覸/C�"#2��Cd}��$@ �t��P���D����n�y��yp�w�e%�3���_/>�pQo}���3�������;����n{�DU��z6ag�h�i]�4x�cʵb��y�;cO������=��5���R�g��ϛ�X!愈�
����@�m��1�ٚ�x�~��M*b ���Z�z]u�Q�����
�0�C
�W�f�|�~|/v���u
�� ���ZH-Q?k� )A僷�+ �A @隙H E^�I`e����Ѐ'�K���J�%�\�蘈)��i�����׻vyN��vwZ�v�z��ݩ�7QU��^�t�!'���&H �=� Jb�s�L�����u��OO���;��v��Y��7[��ϥ˾��#�l=+! X�����T�-w��ł
��$�X�7�� @&k�������	�O��BD��]LI:婢 �A�PZ���@l��ܯ@ڊ��eW����w�!��G�~�gz�?l%PO�������2�9�y����<�y�w�VX�|S���k�\@����E?{��^f���w�X�_�/*�(ú��H�1���2`X�ݛ�*3�z���Ō�A ݾ��� c �������#�����s̢�.�yp�3W��O�@0�f�g)4�/(��;���Gwd��OQ�񽖄)k�ϝ<�q��D# {(<@!�!�<�N�'!��x=X�dlO�8�Z@c1&�C`��/ݝ�W6 �!9�l�X̴v���Y�6�\�0\�W>8��]V9����t�u�Jv7UX�6ʖO	��u-��4R�!S;�X��2.؏^&޳�.8�m�1�ң��s��k�Q��J�K#;��n�oOe��j�&^\�K.k.�����9��xv�9j��=��cu���닮��]XaR���J���Ol�4k���Z�=��R�.�a�Ĳ�k�����p��:;��@@����s�@,}��
�.�^�TH$��9P��tD�Z>� ���ّB@$�~~,!�Uz�]8�I�T��^ ]7t�Sv���yW3�LGSKs�B ��v{�Xy���c��,0�ͱw2�d��Q������*��0���$bo;fH� 2ڑ����`�ȍ��.��(0���2L��5�H�����]ӿ���[k"@~V�	BA��Gvl�&�y�8+�da��~��� �v*�|����]�y�i��^����b�w�����F����x����X0��� �I	�09`�=��0Z���#����ѝm��ou��Z[͚�f��Z��Kc���~�>D�O	ʪby��N;�2� ���@�1�ɐ!�)��[y�ݱS��T< K${�� ������!�@ �U�J�Xe�h������@��{�\�ڞ�}�R�U������r�� �����9c`�'6�js1w*��P�l~�X/\܋ P�8�p��M{�}�}�0�u�ɹ��_���0�����y<y*�.�E,b��H�0L��,5��a��Yv�0M2�XS��gN"x%UxK?�#� ��$] "�n�^�Þ��٪̱ Vf@	 1��i����JJ��&��0���������s�0�̗{�œ ��w ?��@�Ko����Gt��� �Zv�$wV�~��1�e�)�Q0@�.�L��ou۶3\veg��Ō��"�\�@�,���z:s���ޫo���!��̘݋��Q�0��v6#�ff�s�����]�S����n� �&�	`C7z8�%�ۗ��H��#Y}@K��;]� X��RJ�D(*Y�X	W�Ihi���[���{Z|X	�l9@��Ė�."�@h�u�����KP��C��Iz����Ok�"�,���۰�:9�pz8ܪ�`���VmH�Gbh��8�B��f@w�f-�<IxϏ�(,o�DGy�_}SrRZ-�\n&&�2,G0�	�!�!�NJ�!�� �����{�΂�O��]�����*�~.��
�.�we����k�T��Y �ǡ�Z@<�����e�};y���$�5�K��4�~��G��PT4����K�,��f�ķ���cѲF!O� $��tH�rAwbī]�w�$	=c߼���w�N���Pi�Z6].څ��Msp<kiꝗ���a�i1u��}{��S:�>��0 {j�G2 bY A��p��t� ��oc&��1cɆ�:ƈ��D�i�g�<D'NK�U0-1���s����uX�{�k�����`�@#��@�@�`(	�3����8��4:�?�e�:�2�餡��<<Tƹq��ï�5�+d���l͂�o3��v�t'�}�L�H w��K{F�!@� ��`Y71��ǜ���O;���L"ՖIbս�mH�F���G�jmN�m�De�,�����/{�����J���ţ��w�����|:/�}��ϼ������q����q�7Mx���:���D �
F@}Y�"�0C$0'!�T�T�$�C�/��,9gm����<���`Y72 @��f{��LG�<=2]Q���S:�l�$�ϢX�A%�� �_��7�xz�:I��}�Zݭ�U1]&���vR�dIG9���T�u1n�BZ}���!�0����{�� O2@W�`	!�{��"�m���mY;���0$^����@E��nG��
�n����d�Ȑ@wyG�ո�{�H 7�S !� K��`��ۙj�pV3gs��@V����g����y�	�jy��2@ �<��5�ѰF�3
�q$��A]�Y��gZZH��`̴fU���=�' s�_�b�]LI �Ae�I �;�1�w=�󁵼3}%� u��B�/"�T?��̔1�=�<i��BY��wP�Y"�zI�K� �t �+���;�r���p�+��\�M����x�ˑ�y�X⃟���j�ݠ��*��G1���������B �����a��@!�O�/:�x2�䠅�+��E;�f�pi5^Ȕ;��y|��3�l����û�팖��n.Ԏя$"LR��u����.��sc����������\����y1�ȥh����3�1�Χm�(�q�/�h���f;s]�v��GS��"v�{Z��&YB����8�;4/&�nJ��{p��.1����WG4�����KSm,de���g�������	q�u70�.�G%���&ս=��n�k��R%$�C�����vf�AH�s���a�,@ ��tP�����b�����*�e� �B�� ٜ�>��D�Z��uc�,�Ip̯x��ĳ�dK�@U�$w@�d�$��r��@%��9�5�F;��I@` u�E�1�@��_�kͫgS���X���2 os��{km��A�.K��cCTs���=g��}s�<L���n@�d֝���,�<s;��0# � y���@
�r��" )ka-|�����މ ?��|3-ㆍb�v&��n�@�<A�wL��q�I�W���7�0Wl�VY�#L	��VxBۢfN���%�]r�i�70o�ޟ�馋���P��}�$ /2ĢBA$�� s�v���_\�H.��� ��e��<B ��se9��Aɬzźi���s�i���El��.�&�'�����=�ދ�O���Y������W�q)7�'6���A��A��ҘB�F�$�	<����	��¨ri�	s�:U����:�����$�@��:I�좧 �2@-����b0��bE� 'V`d���b���q��q���[�����W� g�"�q��`c ;������Z)��F�A�ɡ�6g{�
��u��X���fb1+�L��ȍ�J�!]&� �ײ��2Z�D�伊���P��� ��Ww�F �]�	��`�-�ސ$&H���@ʝ��q�=�a����
v���Ү�f�X�+w!Ўp#P�M�6sȆ\�Ӛ��"�@�p V�B&X�=q� �ř�wt1b �ڢ���L!�m;�0O~���'g}���M69�w�!u"IEG����>v�)��9�Oo�@�8�0{�X�=�<�uw���Z�Y��U���w�	�Xӝ2X@]�@�%��&f	���S=	ś�~��${�5�[pA���׽��7�4��!Ӗ� ��E�ۆ����S'�(���/Q�6M�����E��~��%H;�w�0��.̌����=��XRcy��g��ؽ�=�{�z�����h>n��M�­�nƇ�GbAi��z�2{�n�oe�Ϯ�g,�vx��>�"�Wf�+>�V�y���{wM��
;B�^�d�}��'$$����ۻ���)�����q�>~����ݒ��{����:7;�rvr������\�N������_���M�g��ž�
s���
3˰k�e��}�ε�S����^��F�SA��1n�d��[{�@�3Sq���`g=�ǒ�͙0)�]��������g���>^k*���/|�x#�k8ľ��;��IS����,�{=��Z̫on��-;�yh����2�3ƦA���e{L���߅����v���F�)W�p��g�{U�;��C��TmgN�9gN��w_L����{ˮ�#�f���l�7ӊoޔ���8pW7�g���݇vD�2)�B}Pt*�u+9�H�+F+ڀb��bݚsg-�>,v�.{�������/-l�[vY(���dm����`��p(�:�`2�>�0g��S�{��dl�#*�Dx�Db�<EI@P#.�H�)-HR��wj$� (@"�K�"�(�a$x�U86�!��5i��Ѣ�Q�׎���j�W���p��]&�v�B��z���@@2�N@r�ȁ�?���yK\H����1LE�����<}g�x����:�NNNN��Ef�Z"�Z���DD�Z���R��=�e���W9�t�p/��v8�}x�Y��^:�>�ΧS���N�l��rتΐ-�K112�ZBʃ�S��n�Ύ(�8Q����x�Y������|||z;Ă��;�sϱå��
�Ǝ��J[˓S�k1N\"H�(�}~8����~8�~�?O�'s�����\�Vq��\J��j���Ȃ�E\��1a�k�m����>�'��e�}���}z}}|~8���TKAwr�g\��rԨZ+P��zD��,]�(9rK��O\�㏯<}g~?^�__�8�������Q�<�s��xM)��U5XX��g��]�h�v�S��1�""փ�\Uwi�[�U*� ��k��ƒ0�u�jf5���X+�+��1�}h�&XQD�e��<ӬV�0E��TPyaFj����Ue����2�8#�O��! ȁ���4 �qW��>��� �}3 � �#=��b0��cd�l�LLߧk�q;�>���U0��I0�d�#��Sd�C����ɀ�	%��bI�׫��$a;���S����́̑ ;g<�G�4�v� �ul�f��.���? B� ��i?���:�X�n��K��nuR��psd����mɥ:l�\ �7�Π<BD��2Ž��b���g�D�,X.��d�p��L���~�����A�s$X�qhb ٻ݄��WCjZ@1�"$%�,X@�~,=��O�~��6�`c���.�"xn��
 �b�v
�5���55 A ���@$�+z8��y��`��@��W�5�2�P`=���;�.�<�7�9�*���eز�fe0����Z�f6��l���~3C�W�z�7Na)�/���c�߷wܳg��p��S�/�������ւ�v�o.����/=�<��8��������!�e�OPt2�� � 8��}����ο9��j���΋��p?J��$�w�ēF����se� E���r�@���`y��c��;(g�￧�)���n�T�.1�u�Pn�e^����ex�[]]�YܹrH@���A�Fx��|���d�1 w� �-=۵Lv0�[{ݬ1�C�L�y� �g�Fi���^PA@�P9�R �Kz�L�7u=խ�u2H�㰂A�� U���fjc=Q ]�&��"�"Ŗ�s�1�=��̘\?��&/J���P�7���	 �����D<#^@�1��R���L,)��qH gf̒ld�Yt�@nlKȢ}�eVyC�������KC*�*d9�<�fm)m
��e��2���ݙ|�.:`4�ٽݏT�W<ܽ�w���#����Nd�}�F�f$�]�Ł��߄��mx2�ؐh_g�H����Vb�� ?�O��,2�}�$�H� }����&���3m�iA������4�3��^�1�`)1ltVq������,��`��X���wE�X��Pg�f�7�T�/@RRݷ<pDl�-��'s��i�̘�	��+�`�����f�=���>�1Ύ�'!�g��e�65'"=��R�ݯ.fѻvK��=�.�h��۳����,v�h�s�RZЭ�]7t�ۜ7��/�<����Ɯ�����j�d��gK�e���zҹ�tR�+��Ҟ������Ч
*������1$e� Sc��M��+�����2,�4���6�^�aф� �Y8��VL��cG
����~ȢF2C%�Ojj�A'��&RΣݚ�Έ�S��p�篹�����]�p�^� z��bG� ��KI$��O�G%l�I6�}�L��z/L��K.(hA�Ɉ�M
�wlȻ�%��;���I%�3$I������rQ��M�d��6�x��J��.נ�z�M5&�l��^�O����k@d-k9��A��C9����?w:}�9'`���&������Pm`��G��d����^�
ڱ��u��3NX=VԺ(� f͂G￟�:����[�q�
��%2d��D��u�Y� ��V��uLKTf��D"�(�vǱL2 �C ��������Nl�ky}�{�>gv���#凳��>�`2w8*@�vb콣�H9vv�̜((��}������H!"D$�@828�(�dz���
�IE~w�ޕ��_�|������ �fV?�[���3�O��V�-l��v@'���< �t�8��;=�e1�~gu9"A������5���t�Ow`�nf�X �eE:�NF��C@b�d�Et���QJ��=�� ӧ��U�p���¸����D�9��<�7
f"+�o��`�+I�T�p��X�+�y�G��f02|�87D�+ޛra6jN*�5�{��YE�F]{Y��2%͗c�#sv}O�ox�"���U���	5}r&�,`A�Ɉ�@֯B]y�a���u�K�U�h�Ia�<ɑotd�%�ԫ���r`��b:k��5Qڔr��ehl���B�Ʀ_�y<�X����w�š�B���O�z�-!���X��HRъ�Tù��=�i�#V�{�;�t�EU�+g�$�-�s�h�sd;e7��B�,wˌb@�-�z�@+������k N�̉+�0�!�q���ڣ �vdJd��F�t����r��������UN����p;ې�
���~��?�>�����?�?ev�����]3��{ѿޠ���~P_���� p��C
���d���^y��??�����w������ރ�0"]�	 , �no��/{=k��X�ۇ$z��.ҝ�0�DΓ>|2A�mK2r�^�	��l��˙$s�'�f�������^k�V��bkٳ$���/޼U�2�	����ͪ���y#H7�|��v�wJ5�T�s�&�6LB.\�T�>~�c.�v�h�~�X{�� �<ɕ��H>�ɖ5Y�-�	�6�OJ��zй�"<(p�h�}������9��}c���}2l��K8%��"�^TK�V
Υ ��vv�P�Bt!EP;�A���w"@L�k��T���P��c���S[�@�w��[�)�)�SS':wØ��AN!ꁦ��M�!�rz�I$�L�$J]�b:uA�'�qPz�'��<D۲?3vn��y�Ü���^:9��;<=�O� � �A�r�ɲއQ�y��旰�(��O�f�T�Qa�:��A�BB�/b�����3����v⮙�P8^�&�6~�=�Oo���K��U��"��F4�O/r���-�
^�'��*��z\�t���8��[\�d�f�Vfi@H��
@�P�nx�!9D��>�\��"�rfd��H.<_���U��\���ں\f�n+�h� ;��{١��Ò�$&�G��9<�kR����Tlօə ��I�ܠ�ugT;�ݱ��K@��	D��CX�]��4�Ð	b�c�^F*�w/p,EU�	����Y&�̾g���Js
&�a%9koy��R�3�'#{�:�oc7}*Q ��qCG��s5.W���мʧ�->B<':�`��h�]�˛�<�_F���6����R��f��驔�Y�Goz$�����=�t;['SCs^�e���N �.7���S��&�Ɖ��C&��s���>�9�6�d߾�I�/� 	�Q�^(C(��2����tZ�gFM�s&���;�nM�y�3=ַLq�d�[2i������Ep�q���(�!�Z�=ڝ���f��6����Mk�o��q̥&�	%�M̓]˭�g����9�5��i3����ĥ���s��u�Nc=��c���\s�z�cUi��Tyd�.�=g�s�tg��mܦ�;����9�\��\��]v��pY�<ܷC��s;V��x�6�g�����٦��	C�:ߴ{���z��|}y(F5"p��$���a����ǯt��8��nD�	jW� �Jw'/t<Aw.K�f���p92���W���� ���C�s�'�nO�|���.��[����((Xk]��"7Fzh�����OS��%-� ���2N͌��;��
$KfΘoK�^s�;z���3��=�i�ou	#ݒn�tS��)���=�@6:�w��J&�)L���b"�$$6�\eE�g����jx� �o۳ �<���4�f�ԓ�^�NGB��sJvm�ݡ�ypu$���'�r{��v`�B��e��%e/�~�Bq�no����P9'�cqsd�d	�H���; ����OR&'P�CZB��{�d���xN�bՃ,�{"�Koon?ohFNd>
�P�\-�0-��vV�V��M�,f﯆
���?�P]A/v��z���\%\�6��~1{g��<�� �yX���!�?��	"F$N�D��<�����V<y��}�O}Ƞ_�#�L��P	�\���IÒ���詐Z��o�fH$jOWp�<{�A��H���2Fiݼ�s�@SE�a��}��{�"��$��ȖbvI�"Y(ɓ,$�<��e
�E=�b��fX��� üA0�E٧�D�d8��;��#Ȥk�bA��N{����'W����ݧMS\�Tx�NS��x��۝��O�m�VzB��&���W����ͮn���s�C���ln����$��e�$�N��g�Ý�؜��&�&+ޙ
KTgx�vw�yG�:el[y���j�c�"����2<�2L��2-�7�Ƙ�88�/Xt��ۚJ�Ӄ����p��dId�e|��A�KG�G��-�`)�KՇ�/P\t�,��ٝrNퟵE��D�ÏA����5��^f�]r<���{�}��ao[��? ?��!�!��B�`a�+
of��@!$�~�Ȟb���<dʪr@��'r�}]S���m^�s�x;:k�I.Wy�i�����/��#��^�,�B;,	����������``6�"	7W�
Lm���G�`w�2Al��)���!��·VH��4�a�іsur���qa�3�̽��ޥS���ٍ.P����� û�0b��\lL� j�D��w�O8���I���x�TH�I�|�R	��x�r��"�Lu�P%��Á�)mj�� �*��äK7wzd�$�Q�+�ѿV�ΙO�oF�����R(��ԯȒ�/�$ĝ].��"��@"����elhK��q���ǄF ]�+A�n��X�V�!��g@���Pɐ�9� �y��~Q�Z����T߲��!~�������5OpbR������z�|�ln��R/��F����~�}�^�M��;jD���B�۩�rW�7�1
C ���D �$%a�i�г�s]y�_݇��S@��E��2c��'y�^�Tuv��2M��D16��mQ��;T�R�=�<��XYE'���ƕeІ�kV¦�H��F�e��6t\Ar��ڽ�����X�̾�E��9L!�Yۜ�LI ��sĔ���Txm¢%��gGD�E���:sU
T���L3���݋^��Hݾ�$�=��b�;�ǽf{,����úPH�#Z�㣉b)�%��Cgd�<zu�����U�H��_�"�9��`���+J�W�\�.�$�
u=�M"��[3��$�sؤ��t�,��lgN��T� p�`�����O�=�p�K�{��i�oY#w�2��y�j�����=n���`ro}��v���EŊ� v̊���5.��� Q���c��=�A|Q�}�rvlU��mV���*���Zgw##|�K�q1��)�m���4����Ic�{=����.�{�K
�ý�.u�"K�lζp��_�wۼ��3�#�珗��t�_Oz�׷q���D�օ����}�W=�Y�D//3^����'B��%#QcӉ�;ǗR8>!�b^��̰���zٽ��ʔӌ����g|3��vl�;=�F����A��j�]�t]T�k��w<�\����f[�G5U\d��w�R���,v�ٲ�q���2��O�}�����~��
i:��>OH�&G}��e���<T�y�&n��{ �W�O�>�b��.xg1�r`���/�k�{�7�Ļc�8��;��,'��,Ƨ��iz
��w�1�|>����d~���[��^����VuHz�|�z�D��Ľ�U��.����4v�Y޷�~�bE~���^��Ept"��z�T�i`�-��ݞ��b7<�z,JBI�_�٭�7��o���@�$xD1{��羔RH�j��Qv��sE�Ν� P����Ol����.Ku�t�V��o���?%�u? @BS�� ��XsF�bI�g72|}�����wv�Lԩ��;JnFf�u���A✑��^�׌�嘕4���^��g~Q��a�*���1����9j1FL{�,PDb����Lh�6�OgS�e�~���|~�>��?q�����G/�����e�*�#�md�*N%�*�*(�ւ��'�z=��^<x�ώ?_�O����||�N�iQDW�\�V�"��5�TƱ>�ł�,W6�9�n��G�'���E�c>�����q��O����||p���<��2�V,���9h�#e������X�ffaS�}>�K,��>8�~����?q�����U���!%^�qe�9�B�.(�j���O���},�Y���׷����>=�w��9�:�!�"VSR��j,|$�A�T��S�b*�kVR�1>'ӹ?3�>?_��^�_�8���P�b��T�e����EQ���8��=��t
 "�o1j��r�#Y��Z����KR��(*�r���Q�cE�Lk�p�>rN�1�,��C�*�a��R��-qЪuJ"�1J5;ʂ� �b(�j��*��Q@D{�TE#�
�9I�o���0r��Y�w2�f.�T�̹��r�G;W&���g�\t�[��J�;sΞ��=�'u��D弻u�x�r�;�\��C�ob����	�MZKB��AytU���D��o* ��8qu�6�k"V�ٞAvnA�#��$O��7�A&nv�]սZ�C�֓2��:��#��)��B�\�,fGL�eqt�b;�jD�	I�&��.9'��.����oM֞w=�#�N����T�S��Ѧ׵�n��N|��#��a�F�d�%�V�,��=s�%�&�Ë���9�$@�ٝ�^���<k�Y�dni,[1ַ,��V��M��j��=&�^.�f��,�$�Y�k<�[(�n9l�q� ��g=�6�9u��]
n���l;Sn#�k�SCT&�aٛ&vQX�=]����2�zy�ђ[�\��*��ܰ��yͺ�b뵬�ۧ��v�r����"�3��t1׆�`b�t��5ͽvqX�dbW��W:�H���;9
��Z#�Md��=v�^1����^�JKZ�1����=���r��cZ+)�34"(�Lf����+���\e�N��v�g��Cp�չ���mn!t{{m��wg�uIv8�p뇂uZE-Ρ���0޹����י9ö�Dv'c��.݇�F�ݍ���rm]c��e6{B��d5-��Q"Qۃ���	̊�n_#�=�c 㨷8���N"8u�:�ɕ�ኻ>4��!� ��9�@�96�rQm|��>_5] �+��큚��������.��0T�a&�a��{q��!��]#r�i���a6
.�=�Y�n��-���y�/1k�n9��)�Mj1kv�8ضc���t����INo\�+��.�kt]q� H�q����;<����U�KR��N�K�c�,�wnu����6�َ��#c^w<+\�Sq6�V��9����51�U�dk6�֡0[-����+� ��$�FH��"����&ts��ڳ-[�6�Kv�	�̬B]�1�9:Z�qZ�b@�cF6k�1�[�1Lm
aRcpm��U�V����<����B��"��Y[��m�9S@����B���3Y��.53C`��҉�H�h�ywT����v����r�'iywm媴�S�/v�J ���I����&����c)l�ˈmiYqub��j�;q�c��Ǔs�:J�wnkz�4f���Y����":6ܚ�P�����E��<$K����;�J�ߏz�d�oѓ$��$���� ��z��S˿�6�r(�w�ɤI9�c$�1<�9��q�i�Q�1��}	$�];"I�? k �����}��:��	ѱ:A��"���t�LQ��>�
PD�F{.}U��a�"j�`K��� ����0�bH-w�:��?��l!�Fe3��y�G����7s���q/����
6�ɥ��}�b�PLD;�xx�(c�QJ+��Q~KՔ���r<@ ;�G�}O���{~��~�H	���q�M��5t�N��e���zL)�R3�IMY�i6_~�O�i�tl��S�ə:�>�X� �z�GQ�u���CWcyʌ�䂂����9���NRJj�%n��H�U�k��6g[5�q��
�w&n�?��`���G��L�1�{�ȟ�.��"���O���-ֺ;��yzd�lK�qG?wy��{�s]��($H�$a 	"D���$�y�s~������jϿ��i�Y� fN���l�����P�	0AZ��8��,��I:��k|]G��Ww��;'�ڠ4�;��HL�ʱ����9�o�퍅�����d�ޙ�I{�����y��B�/9u �qk��t�$j�a���h���ğ��KyA$���3JԱ�{�e~��V.�Kc��	�6��1��:����Y�䫌��p�np瞠�79��H����)x������+��Y���96�˞�KԐ��L�(��F`��+P�֑W���0�@O*ɷ�1���$ƿ*�;#�pc �@rE^�
j��t4�����1�'��	$�X��dB���铭�q��މ�
������7N���:k�����٨�̛�}�\X=�d�����Q5�9Ջ����.�>�;�x�R��L��@��a!��)-	H�$I$� c=٥�Amm�}B�,~��d�D�LDC�'��c���.gwL���]�1r[�왖Ar�S?v���nKy�ٓ4"�p%�<
EY�މ$>����0z��Ѧ~���$	cޙ�˱���L��joV1O��?���ٶ1��g���f����ƫo9���D�u���w.�"�j�۝�B�she��d�d�*=�M���ĸ��ZYm\� ��ɒO�,>d DC��f����W��F�h$;)b�=�)� �!��(`I�}�I^���G���7^�A
x4�\H"��!�Ab��
���D$������R	Y[a��Jh�A��ǘ(X���`��黖v��'�bĎ�d��͗73z?���D�|?�ܣ�p���Oi���p��Q�PM���i�O�6��?*�Z}L�@�)���P`I�z@��>!���C,3���t@%���̨��J��@/�&Ov�(���E��_\��$^�ΖLEZ�M]���_��O��|cx�_��V%ڻcZ1f��1�Y�uK�u�Z��0]��_�y31%8m��������*�}�3z$�h�a�v�w!{�2q�A�K�Y�s �U��5� 0�˩C��iw.��Ą�v��ZF3�����{�rI�[|$
�z������)�Q{�NQ�w��2ro�áDCȠ,3Z��{���v2�C�z;^w%��9�����%���]'	��� , t^*0�8���c�N� �f��j�,�\��\���09N�&��,?(&IU�^�y�1��wؿi�	�e�9( �ḟ�wbO�zf�B��ݳW]����CY���n����3�:�����m��}�!x4��Y��y,Pv�T�f�) ��tK�58ǘ�S���4����He!��P�N����_�푄f4��@ظP�̑Eڵ]m�^��oq��
z%�F��&���[�u�!+��%��Q��4�kH�3�4��6�s�@Y�0�]I���\Fen"]�+e�v-�"�Ѱ.�o�l��Ʌ���S%�N͸���f����
�����dzs;(��il�n1t	Fcq�[�[��e����kHV�GU��Jܜ�pn�}{&�����})]�������p��(�m5Z��C�Yy�5������1�?߀d�� ��z$̲xd���F�7�x0z��c�B�)�#�$����\��x݄��NtE1���n<&����A+��$�+��2R;�|��! me�w&15��ܿHH�CVF4�����"c֣��)m
��s�bX�z"Z�%GQ �Q��1�vD���,b��K	 ^�S)���7��!�o�S�Έ�A�ry�6߰%�D8O������{%�o�?��Z@7��Xe��hor����:��Ҩ>Q�g!b��qc�Zvwm�;���ڒ�sf�����(	F�sI���T	$��$���L�Mߢ-� ���-߯}��̻��3��,n�h��t�1�<�V@�.�&��c���wxL�3j�t����]3�����;V�<�����N�C�4�y?�����c�µS�X9
P�"����=q��C�2�$��nH��%��� ���0i�/ �]'���:�����U;*�L{�<� �M	1�<8�,��E�7� ��~2	���p����WOL�k(�5>�1�	�i�2�p�t�g+3�ň/M�ΌC��É�H_� y��Q�L��͉5pe�|h�EtR�L�r� wwH�٭V6�ДD��~�����g�f��G0�@P.݉���cbs$cd\/n1�'���z�۾I���,�R%�2��T�|�j�^i��.n�b{Ӷ=
���R`:�fI�#ޱ��"���U�&����A��2]�3��p_��� �
^���@/�.ؔ%�H�A�]���gLI.�R������?���Ǽ��;�p%�f����nv:�zk���M��M�W�}���py�^�K�͋����.�]M|�`�A)"a
Jn�P��λG�3�E8�}��B0L��.��(4(/N{���J� ��~�I���=�@� �>��|N���˿��yׅÇ�R�����G��7w�:�h>J��{�2@#̐�Α�H({9��[{L��O1]4�,{ j��Fǆ۵��p4eq���юe�lXXUJp��^|9�A���]�b�D�%9�F���	��Z�u����&d�8���܌����T��������=��_Wp����$�Fn�dւ��)3���QW��68��bhN��t(H�^8%?�e��l�9�	kb�Ў���(1\�Q��a${�.*W&"xg֢�w?u�wfT�<�wފ'�L��D@$7�OxS��'�o��~7�7w�^#|f��S�GI�ˡ,���Å?t>ٸ+kޓ9&(��u{���i��M�
��S���E"	��8FLU��Ͼ��h���]��<`���d�`{F!����d�ɒA�J� @,}����������*�3�3l�鹘��L�qA.�	�چ�VͶ����Kk_?|�Yf�Mw�ւ+��pÁ�Ɓ$�w(/2��C��|�C��d�A�~[�!_9��h�z� lS�CI qu�(���1 �{�r��X��k�wI�����P���`%
�sy�K�=�$�O`�xQ���z�mP]���U�Lh�n0�^���m� ��H��Sc��Uzף6�Y�<1 ��ր�N�td;����u.-�\���k+ؼ�0�xg�'EF� �^��s��nA+�=jw��!�z_~a�����R/��Z��@��č��=���T�tMR�Q�z���v�ɛ*j�`����5(ɭ�����R1'�(�Ii�dξ�|�BV݃-��+	�\�3�����0�M���A�F��+lY6��\]�]r8��q�K!���s(�4n�4;:�h`��I��c�ٲ�q���`�Ŏ �3�甓.UṺx�vV�g�v���!�:Ch�[��]2�Mcy�Ύ�Pt.Y��7�:�������d=w��E�3�f7M��*xlBڮ3Yxό��2��70���D���ü�'J�ڴ�1��i�ű���n�����N�
)���-x�y���!����.Ҽ��z���\߮g\o+n񻸙R����g�� �D�3ݓ$�eq>]e��g<ܳ��%s����'��I����P��!_9��E7�.�/غ$�igql���Ѿ����.�S$%�B�Q��M��P�wx0�t�T*����{��\�Sm^ֱMi�t��1�=J9�Q�fO��`uO�I&�r�)a���W���Id�������V��HH���\A��L�7�:R6le�j�v��m�Ie�����������ua/)��5]��9 �J:Ѭ�)0�e�<�MU���KG`����'w�
]�KB��'�!q��WZ�|�o�|�֕����χ{��Ӗ�4�\ї��H焞��ڦᑐZ!TEO�qĤH֑-%1%�L�y��@^{��Eﾁ� ��f%G2^�Ԃgٽ��8PR�T[��X�e���$u���~�̕�jؓw}i�:��;@$k�E�$9����R%{���t��!��K�L	$o�	bSs�-���8h�D�wvUs������*22�M:r"��%��b'�)���m�f��V�ޙ�I,v�����Р��mxFE'��������z��V����86�'7nl##�(�6JѢ�`n�G-�G?������P�&��$���� �܈" O.� ��p�yړX7"Cc�����^D�D�3��l�(�{�q��#�n�LIb3ވ$d��B�|ő�q9W���������=��\��
P7��fԁ����{$ C}���kOks�����f��f�͑J��O���p ���Oѧ��8�&(g%�������w��P���n5
�{���l�f���o`��(�9T��x��>���+q�~f�S^���K�>����w����>ޚi����V,_!w�+���u��O-��0-۞�x�׬�u��{o��pɖ�g`�Wѯz+��n�~��m�ϧ�'W���O׹�r����G���M����F�˞6��Y�0����|�u���>��=���寛^;�ybE��/vX���f�}��(-lnХ��������ɛ�.���}������ع��UK�$�!���m�Z�����	]ۏ<���L���)Mz^����g���㊩�[�2q��lNԪy�U	�*�9^�g�ңۭW�u�x��a���0��2U�y۬�yW��{*��5�=�w׺'k�Ǟ�ii���x�u��5s������.��.e>�{AN��N-��1���|y��ٍq�=��<[x7z�7�y�����m�(�a]�]o�������s��Yb�������M����ox���N� b-��`�>�N�=i��={x-�5���qai��	#��  ��}��ˉ�������i���Ir�=1s��p{Lf�8����v���n�����E}��c����A�W^` �g�=qf�3t~�Yу�{�&�������'��Kf\�6�=�og��p|0��� l�F�0UX��U�[AJ�z�����P�{�
�8��ǌ������l�rrw:�NNt��DR*�m�り�/��m���.���j(�y�:��������q��u�����㏏�W˝�릎KO!��DL�1���h�SR�(U�B��
��N�W�};��Y>�㮿_^�_�8�����ޏ#�/�a�r*VJ��4�+ib*&�ːņZ""�嘚�;'����>��?����>?q��ʙ}����%�ت(�U�����{��ڱb��>'S���^>8�~���>>?q�ߟ&���8C�(U�TR�����^m5b�iJR����QA�*�DL�����Ǐ��������������6(��������*(�r����Q��+2�> �2�"*�4U�W�2���TpB��Վd�=������3������OO��5���G��Ir��2#D����h�bBҋyqGF*��D|j�k�\h"��b'W2 �O�C)(Ԗ$R2�Y+;�n�b��s�O�Y�Ӟ(8x)x���M�+���w�k�H�۴	W���ϝ��(����)qK�Z=~"r
�Q"�� � ���%Q$4I#���,�<��3��gjn�F�����C7\p�z�n�d���+t�����:��}""�B'��)��0�tX�h�~$��B��Uot���vkէ�m�e�0��-�% ǣ+L�^"dU���H2:$U����K5w(�C�o���!w��o�����U��i�'ab��F ��2sa��'ݐ�@|������.���	�]�	g{�J�Q�;��(UD�1��{�h��Ǧ�H!��H�43�>�m,�R{���J0�5��c�=���;�Vl�wO��t˝���_q��zaLlF=�<�w�Z?��>������FV�
�0��� r1n������(��La`X�}3/�俱�1 �^iD���uP$�=��л�Ӂ�@����;�P`)�I�ְ޴�u!�B�F�j$���x2�����~��0T9��Gkj7�c$<��$�2BY.�}�b��'o �w��O��y��Эʿ��F.)���^�x��s�a� �#��	���t�(���<JqYɵ�S+S5����m�=<�ʵ�6�	��!�;:[cT�)��<ԉ���/*ms�@�Cȱ'���^��8��<-��J���x�!�ܜmwW��_7d��/�I�~wND(�U@�f�xHY�@P�/�,�'���̔2wL4s�Р�i���6�Ŧy��P��s�"�����툚�{���Ox19=���4$G�#����Q�:<��C0ܳ7oۻ�0��"	$f0�bKg�&	�h!�=��3���^�N)Ѩ9�q�r�/��>�_�1��&���S���h��<�f�N�ax������q�7�Vy(sm��4�l,�!ɹ��ccy8�]���J%���;e[ݪ3��Ytvy�;Z��:{e���^
�nf�v����t#��qHps��]����3�t����XðS��	]����6�	�RX�[���˲�N��fZ.�eֽ�ʥ���k�k��J�Q晘(7C��е�����m]
V������H �{�v^�·��3h.�U虦Hl@Z}dv`�0�U����ׅ��j�!�����a�5;�C�KAn7~y���VqN�`B1�V�=��q�eLa	�P=�>����I�~"N�߈�P"j�v�0?U�=��>��S(:`C�A���$���M>��ȂEx=^i��G��lB �P��9�o�|�7��$	�Z��U��^�c ����G��Vԇ�>;��ݝZi�LnnX�b
%����+��]6�db�ew$��{��Ә)��5��j�"@$�� �`�<A޼��yʩ���A��	gq]�ⓣ ��(�3��$����w�9�TaʡJ�>C���|Ew�8�L�Z_���0w{e���/�joB����2j\#��W�w7�����JD�Hĉ4"J�e*0A��\��y�S'��H]�k����r�_�� ��aC�v�i\"@,}Y�$E4��ӣ�j�^A �+-��dח������b��߰�>�,B�����7>N�UG�"vz�X�
�O�M���u�5�II<�T�V��8�uaB&��^_Ѥ��=����u��x��L���e�{� �H=�#��2��-����?'�}��]�4�rm���4a+�ҵ:�8�F0�O��wˢB���H}����"�:%�;L��� ��L���P�����o��)�Q9�l�x	Ҙ�G������řm�;+��~��3��s�(E��<�F�A�� ��{�f��(	�(�@�ك=u2H &5ސ �J�W��LG)s=��*�d����Dȓ�a�����rR�w����-=b61�*Ĉ2�Q@���AGR0Il�`�阋�����k=�:db���c=�p�`�0��;Yko3��{*8�lu��#�ƣ:$^��#�r������q��� [���Ӄэ��	s;H̟
�c��K������験���1ȇa ���PL��z���}jVY�lM�*�b�p9�^��[ ���kt�j� $�e�w�~��:��=��?tddɆ(s,[�Q/��*C�yɈ�Ѳ<�$Q��衬�}�޻��C�TD �@�h�A��汷ۓ3ZN�� Nvx���PH��Q�W�s��${k?(P`��<�l���u�b�A ��y=	����1@���q�Rz��
�`"�a�zzg8��^[���,����@�{��2Gy§��q�L�j��7:c(�)�W��z���m�L�?xjk�K��Ǻ6{s�2x���{�͵�E�"^��0�����KH'�c�f��<O��Wa屭q��y}�z�^w�dOc�"Z+� �m�_) e��~��lZ*z���w>���N�&���֭�l��#�-�cu�f]���VڳR�E�>~���)f���%�o�$�[L�<�<��G2�WSe��@��r�C=y5��'@��H7�S ���{�_���S���	d>���}��mp�����<�0o��J��D�I*#���d�G���b�]�� � �w�e�ۡ���A���-��{�W��Ϻ����X�$F�t�������!���%A7y��T�9��q�̎rcn��os6�����D�t�o59f+�<�]h�^��Eөw\���7_������[gBvA�n.�G����?w�I�+�ܓ����%i��w��GE� �gI̦x|��!�-"��N�#X'|<�p�܄�m	���#�6͊��bB�ڶ�p���,v�MH��д��1&��]�R���Þ�S�hy���3Z��z�˩LLfJ,"p\	�x.6�^txx�L�z�HA�x���};��8�`{;�����Ÿ�.��/�e�4a)�Y���c2Ҥ�0aݭfQc�r\�۵�'{)�ٮ�r=Vm�`�&��r���v���ōxqRog.#����s]X�#{�p�DA&!�Q�����/r$���&�t;C(�vA�ew&ƣތ}w�lݼ�r� ;�ؼ�e{=	�V;שj���C���H	��t@%����W�I�r�K<�"�f#	�H��A�H�뎟C?�^�(6�y�{ș �.�p%�&���!�v�Oqc/}Iz��Trx��~�b(dkJ$���O��W��;2�m������xw�VgCG��"ȳ��]n�x����d��yɦA�H,��T`B�(1ԭ�.N�ϟ��H��,й�.��E3�:N^���w�����zv��c��זĎ�	���ϰt4G��Sw.�� �d7�yoq ��i��fM���^b��ion���764A0���y+$o	���y���n�ؽ����7�Qǖ7���0���-���5�9N���=�!�<���{�7����+<gHx߹�O�����D� ��8�d�7��B|��rc�&�k��ђ	�����	w�Ql���;F�sg�I�׊���I��-�� ���L'=�^L� L��ªf蛝��;}>�H1}��Z�<���DvGOW��)׼�����r�"��ڿy��!��AEy���y�$n�bA����) ��=\��HM����[%��!�*�������ߧο����[tnх.��M`���F�'#�w.�ݏP�d�(Sh	\j������[�^/,bA߁�� ��6�����di
�dp�掟L��ډ����<����������d�\'�[uo$�.� �'��dd�Ȝ=ڗv��}m�ƈ0�)�H� x��ތ$w!���������mO�D1�dj(�_�+��d��}��p�Ρ�vk+xj˷���k�dVa�_r�A	$�*�(1DR6��R%=wO���}�Ã�o	���pr�C��v4���\�,p�Pra�5��l쨎�_��[��{X�/k�*�]�3��`92+'+�$�2@���c���";,��$CB�Q�0���fI%���;�=Q��\��/�0�D�!��9 k�4eϪ�ݜ*MŃvz	z���??����(�A��cE��g]w�G��YwC&1�R����sԴ1�ށ��6�p\���a!�:���9��~1.�����s��$[�L�	���f�6�ׄRս
咍��@0�"�r�2���P��~��{ Mf����E�g��戄���pq�����7�2Z׫"i �43����=��['�'�zP�J�L<>m��3oj�}[���3���Ue�.����>����x6��F6���9\@o&\ĽWL�>��.S�(�6� ,MGJ"�D����;����ҭ�3�LI&�� qM�����z��s����"��"pTAG3�^^��<���Lv{u�ˌ���ѧ�� ;;�/��y3�)93@�w^��1�2@�lA��+�,g�/�	�1}2��$�*�^i������
"yp��˖Ԥ�fo�����4��}cD�?()������Q/���2�p\����"	$5j��A
�п:�����^�A=�t`�˹�;�����,sumUc�W���K�� �<�j��8�Tu�Oq���8}��g�1s1� ���6��D$LM�`<r��X��ؒ�7�;v�Q�Fu��1{�	�3E30`u��W6��)���uBh�Ξ1^���s^���{�=md��Mk�20߼�Ǔ�F�E�Nξ���>Fr�$�[�j�ܼ*+�ϐL�:k�W��.�精�iߗ���폲�V���4�q��(�F�=Ҏ�Z�f�:K}�S�w��>½7�s=l�_ݛ�+����g��-���kv����ܷ.k�Y��U�؏�#�bk�Ὓ���Ş�?	q��L���u�|�3�$|)�;y���ͯ���w�}�K���%Aeo�䧻�f�7w�ŜG�[������4�Vj���n�bs6P�Á���	1��m�t��Jv�?yzQ ��Yݏ�//c����dǧs�o�po8��W�
߃�^;�a�����l�s�8nv����}��V��Ed�Ȭ�4Թ����ۖ�5Ot7Y<����������=�
��=�ͺ15��ѩ�n�S�"���u���x�p&���MOwô��^j�z�̚�����ˤ`�����s"��3����wr�W�.��xm��O�I�n��ݫ^\3F�������9�+���w�������l��\��{BB���r��3��o�~G&���;����7f�ޫ�/e>��O6�ਇ�=wnӇ)��{z�F��pGө��-�xh�r�@��������}�?��	0M�{Rƽ�����yg�ܓ�3����5�ۨ���l�]x��� ��e���wV����R��AAj�*��#P���#<�~�ru>?]}||||~8ツ�Q@\�p��*��L�p��"��E*��~I�G��|x�������������u:�PEQU��VwL �e��b���(�|J�DU]���>������������u::@x�*��TEb#�a�R�T��h�J����*����CQki��r1�O��q��}{{{{q��s
��#�RR�Ѐ��C������#����p���79e��}}fq��}~���������T1$y������S�1�Ƴ�xʈ�V/����E/WW����������ٳfΧ'ӝ(���b���ښ�z�-
��r9~lOhP^�k�UDƽ�AA���P@X""�J�)x�"jU">P(&0*�J ��-�J��D�P�XdޭN�`��P�)��p����G7�!�� �� �g����*/L����������b�&�s���EɟgB�񷟾-����O�Վ��:�7����օ�L�Zi2q�-Z�IbJ)S%��2꫌SC���k����@V�&�]X.q���n��n�N��H��l�����P��Ep3�cۙ{#ѵ�<�Q��N���=q��+�-�=w&{7��\�촠���:�д�f����%��mZ�+=���<۲��`��s�ݽ7�[U����byͲ��̓b�8ݺ-���s���DZ��eI�)a�mD.+nI�X7n/]�zR�hw?3��1˒\ i�m4�����'�jX$6��&
����;-��L��i��4�n-\��Z��`w�����5�R����SK�Uصs�ss�n�haNx���ݴ�Vy��'rk�G6Ŵ�8���>#a����c�fIwP��wAB۬�6������	PKn�u��Эe�]�U�V�5a7ֱ6$��3Sa�����k���Z�Y���cbLE���S�r[͒��9��t��o��c��8�sa+�G��2��6������7P�V��.��M�Xu�ͤ�`�w`�rC��+zƓi,`Ƶ�%�� ε�m���S����0nV�g>��y��}�^�M^]�(���m2+���u�:Z��ݴ@O@G�E+��˔j���.�!��&��[3�溺�{u�onS\��k�T�]G�#��m՛ay�.�{	"����g�ז��Q:���$�fk��f-������Uq�<ڊ̈́"3n�ڸ�.3�J���;P"F�Z��6��.��E�q��a�9/�/��wm��7=#6��Ws�%$]�i-�؆�.9@��-����h�2����0�&��<���nZ9�E�뵵[�H�)���x������v�r5(��y�=[����`RƷ��u�6�Ī]��b�J��1������A�p��]���x��|N<�[���m|£0��bR�it�bƥRm���d*�vP�[�����E <#$x�%:w�Jl��L��n=�x�e�h�݂w�b�u'![�v�;t j�.��Y4���k�rv󲙮����������>㨱I�@&}9�[��IIh�KIu+j4��9��1LՍV�V�ײ�v͊.��導�k��/�Wt�#n�Of�Y��^�}�ɻ$�[3f�*[5]LU��+g
���3�pV��Yc�Fa��f��?y.C)J��k�0�	Zަ�4]�l��r�n�ƶk	s`j`����B,~}��<�'����J�����tޠ-�c��z<�^�c��2	�|�P���g�0Jtdl�����0G<�!j����6_�,@B��\�c�/&��e2��N���!�c�m�7��I���#f9�h��w����վPI�wD��Q�cs�'��x�@û۱�y�i/�'�C��2D�'��SF7��Tjc�PM��������w�"i�������^:}���4,�m�G�fdA��O1;睴y��"b.C�8xq>�S���h�%�a�K��q�y��<#���v1���_�Ѥ��H��D9{� [>�<>��Wts��A7�t�i��ē��sH�~�i�����E$�ɻ��.t��4 �o�{��2K��#�����>�p��W=������tqԅh}��P�VL�Ƞx]��{��;�f�$_��E>�o}r�{��F2M�����A.�׽S����7G�{�)Y��=�mCJ#�=��*단)�"<� ���t��� ��o3�w�9�$%ܝH���ޱm1=�,s��_����x���X�dխuA��]G�gg�EX�z!51@y{�QI���,!���Ϲqy�[˖�/"ńK�Q=�r�g�l���&�٧��c�q�(#s���;��&/$=�p���$�� �l->�$�␦c;�A4�g;��YL�$ǚ��O��&۽��������ɒͦ�Y O.��}*ޯGGzX��^�xP���k>1p �K�E�B�ɮS���!��ڇ��|�Yr����Ml��6��´�����g:���x�3s���wJ�ؤ�;�l��`4�������4�(��(�Um��<%��se�4�b�Y9�L���I'Wrh�{���yj�H���P��1���\�A<4Mxl�� ����Mڲ�c^_@FDX��( c �wGL�3buS����!�I]&�Kg���6dyx�.�8��b�����aK�˻�l!ˢo�wK��4N��ti7���,�1\��͝;��sT��d���>��cgq0���%A�IxT��2ĕNg���P�SR�d��w!{:$H���r�@�xLH�>70�z�"y�1>���]A�R�VI-��2ĵe{^%�C�ڡ��:l�}5|��1�6#伵��2�zfI1�Ԏ���_��2�.-��"#JZ\�*���F_V,�ۜ�n;�g��i�7POh�ڟ;zo˗$ŗ���$C�`, �*iA5>vO	wF�}�T	�K�f;���#}��V�2ǳފbA�7���s_��?$��޿��i��5<<�m�2�:]���ޭb}\�a�}vM.a.��U�f��߿ߡr1؛����92���x�?Dz��f�6q�Pƙ5H,M�Y�b& �W�I2FW�"@�6�M���.'e��9zB��t9ioFU0�|\���m������s��
I���J0"�[0
��P��H�z�s�]eOvڕ]����!�����s��81B�٬x���_s�p��ȒX�E�DZYx�)����rH��bIm��!i/
���)�bOr��H��ڽ�d(��I ���rANH���O���ٕ�^4=�t73e`���>�E�xYd�iMV^鍻;�m*���a�ʙ}�*�'I����r�KҚ0GH�rs&�c,���άx%��T�&P�-�ݨ�Bc��N��v�\���;�t�HÍ�Q��f!Xg[[c�Ơ�:K���5�P뺞��X�;�K��v.P� \��֦�̶�`�̶�0�43��'�V�oN�&��K=����T= �Іq�ѻtՙݧ����:6n8]l,-�YY�F!�mN��!{�Rf�q�3mш z�:��]ډ���E�+44�Ԧj��N��{�ی��19�wi��vN���C^K���s��]�)n��K�k�����ؓ,r�`Ǫ��B�QQD�8(��q�;�7pg���M��$ϗ�c�"}ˢ_��߽��歱����������r�M��Zf"Ǝjh�D֡[>n����0$��r�[;3��".`D���
v�v۲9�� �U�$���{��ٽw1�^��$��� �&��x�w���e�s��dʳ�%'�l�	��վ ��1"|��y>do�d�Nrj�=c�& ���.�F��Au�7gۓh�F�ΓY�ܜ헎[�7��O�sm����{̚((~����I����Cn��}$���;0!؅kz^A2�k/]��1wFh�s[ܶe�����wBwo",�O���f���5^K�����x���������{�5ū�pg���=�x����Ķ'3�sx�j��}<{0f�=�8��������<Im  �zv�-�^�g�2����.����x�~��gTc�t�a���y�i���9�#}�$�d����)c�0��!����P��uq�2}D䍾A.��Q �x�&w3ޤ/&DO��=j�Ɛ��zD73�%�]o���L��U{w��".`EP.љM��%���wվ<��x�"	��6�{�Ax�U����(���ue�e�9�i-����s��81�P�]krW�*<￯�wL�y�_����6}2�כ�no3�2]��2%��腂2��À�wL�&����!oAY駂���X���Y��X�}|�1�9�����s�L����d�]њ3[�[E�"H9� $����HPM�����A�f]��<)��.ճO��0�1������t�
�N>V^����eu\��^�S�o�S�U���D�"�� 1>b��g;bA���������{:;�*�	f��5V3�k&�<�i�����"y�Yvj��޾��d�g�fN@��*	Na�Hk���Ω�I�ZT�J�o�>��P<��tȒA�ah�I�����<)�����(G���t�)#���'3\<X:���K��g�a�{��P� ��,X(Ȩ��2GϱR�^��X���[�T��8�����Eq�f�����P[|��Q� n;�
2�%�*:7Y'�Aw'_cX��,@�B�W��)�R%���]X � ��8
�X �y��ӊ�mC�ªe`�0��&�@��y�C�`��7&��x�ͅ���<z-(�G��"�pڦ=�ڷ�Q+�M��e�5v��xɹJW/7"��+y+�|e�G�r�<�
P��|�������3-�>�0!\P@S[-�q ���h�X���.��o��$|�G�r�%�l,��gw�)ё@���}3�K.�j΁Y�6������&;��=7�4_��wZN��+����7�M���f��ts����m��?�6l�~�S$����s���z�Va:Ld�0��'�BT!�5�1�@ҲT��X��*����O]�g��R|$��b���w�<��~B�bT���� �g@*�)}���,�s� ���i�n��c�5��wjz�^~���}�}�V�mR��],�ؗY`�UoZ��"D.�
Ms���IFė߹���p��>Hn`}��A�f�D3�p1��q��|~����[�3>qH�{0	���.`G3���ԁ<�d�t��r ��\a�#��d�el�̾�|g÷���L@xP�%�ڮZ\�M��bD�I9�j���`K)_($��9�m���qAYQ&�zd8�����L�!��/1C}ޙ�{3�]������%���i�w�˿ ��J	���2H]��ݝ���l��O	���}��$�y�9�pN�G���K��%0f�AǼ�^�2ল6�$�hĂ�`N��]�<rP�`�>�)����'k�f��|7��^e��>F��W\�~�y|%��!Z�KեT�u�:4����Ҝ�
�k��nl��洨{r��p��;T�	J��.�x�0j��i�a���=��x�eN`�����c33�bK��̢���h�=Y�gm��c��|��(F;�I�B=��Ļ\L�F��.竍X�����q9��'��㪥��z��m(�+,��T�DX�[3n0ם��	�n:�cU-�Sx���^;�Ds�r�lj.k]�g�L��=]�	�T���E�����׉t��y��>d��z$��=�̶���qݞ��m���Ѡݔ'y;èyf���:�фu��'�ޙ$��@&_��>>���k�iI"�w�����y�'��92$y�8�]�d�'��a�8�������L�	��"�׋������$ܲ����a<LĐa�w8r2x�-}�[�4����"�����A��z30h!�|nr@�Zs%����sޥ�ϛ3-��D���yv(2�4�>�ˊ�}�P�R;`b镺�ZgV�FF��1v�-���*��;4`"@p.�Ef�Pr�%����ˁ��×r��+���9��I��P �{���<4+k}��b'�����+5��]��<紘xS��Wױ�/�)��{�y�%M�&d��K��4M�ɣ.B�:4�@���fK�Uǘ�q�:D�%��A�w���<����`Nש���e�s�<C�{�h7!1k%���mY�j[�w�d���@$�?%�.�".aD���t�g�޵�*��{��	9�d�p�%>�L�X���g� ��f�����R��H��{�N�Ô�D���l���HC9a��"m��-O�D��X�?
�<�J��PblK��]t6��X���n�]c]���Xj@g�^�|NL�tP�q\ ��8뭐�,�������z���%��@��W�r�	ȫS=<����On�nc��A��Ac��$�B�}����Y�&1�!2xDC�X��=�H�y�������}���RsC:�~�M[��Y�-�8��O��N"A+MЖ@vT�g�Ok�\pj��<_U�VO-HVĳ���P4M�3g����c�W=��طc���N�+�ݧ�:o��b�gh�:�n� j�'�M���b
��F�����;w5|�Y�z�{Y��I�����]�OQ�A4O_W����g�{�gn�ڡ������d�}Ӓ)y��H��72�����4D�{8]��g���H+�4�oe�}�o^��9#R`�^ILU��;��9�s��z<L4������}ٶ����)d�i2g��X��J�@�_<v�g88�60 ��ާ.�=�>�5���U��,�/��{��6�{;�������n�p`�͒�9r�yoFd�76[�v�Y�&�3}o��뱡�K�N�3|/����ݞ!վ(�;��٨.Yrg������\5mԯP���p�C��nB��vd�3�<7R>���zq��h-{<N�܊��8�4�N��u{�xOU��sd�e���ē��v���{4{�j������[>BMbil��)q��B��2K�&��o;���e���O{{�׫��Q�$�NFX��:�5��^��N�vx�����&�̘Ǻ�1!	2�E��i��c��-)ȚZX> 凥h����v���@j!�MQ�X_���,�H��Q뙢kw�1:�/�ӷ}��+̺�
�?>��Q����O��u��E����ҡ���[Ω^9�,���R������=H�ϙ�Y͡�V�{�Lj�nQs)��L9�	$�fZ�t+(��"s�){VW���sp3�tr��x��2�l�_�e�~�D�;��_�? Sr��+naL�D�)3l "	� � ���QUTb1A��<�-��
�8�3��gu�׷����g���3c=acl���$
Tv�!��R��O��;�EU��c��~�Y�}g���^�����}s���pf�����#ʣTP�P����Q�BTPU�z>>3=�ώ?__^�����}q�ɾڣ���)>P�L�Vj�,�T���T�*�kO���Y���~�]{{{{{q��
�Op�ANڂ��v�,�%zID��}|f|u�~����������gp<JȖ�;��RZR����C�DU��}h��a�>�&q��~������ۏ�|��>�����*ʈ�E����  ��~1&:��88pp�[�U;��!�TR��("6�U���r�5�}!��Fj�Df\Ū��0"��Lj�B����VZ�m�q�k����XZ(�(��"�I�gIz�a�K�M@����$;�=��� �sx��û�w�$�`=}ٱ<qg��U.�@vߤkR���{�V�)��,�YcB��B�ك�dy�>}}S��P�����f	�� I�(����XβS[����q�:mZ-�X"1��n��帡��ë�#V�m������ϟ�k.�7����޷�/����D�b�DA�3w��40��~8���fNȑ]\��O����\$f(�^����\K0b�ڜ���w|݉bH��R����C� �,:���s�v�w�� ��Aw+9��=u �{�ί�}�,����ME�&x�٫~�A:�""���s�f�/Rq�+��O��P}�� �ܺ����t�o��䌂��2{/�׸��vP�[��_�9�w��':�ԄIՔ���y��5����^�n?����v��`��(S|��֜\����@d@�W	SZ�3�y�:x���`.�!��qǎ��Z��w�j�H^�%�n]�� ���y����S�E˄�J:H�gK\�נ�J�XR��'�Q�L�m��@�bz����B���vJ�F�;c�f���D���H6:'����~ɖ�}�m- �z�� �1T�rl{�l��w��f��]S^d�	8�@Q�L� r~PD;{L�"�8=�����!Q��y�'�A �G^myQ�d���H%�=�ld��݌�H���b ������w��)Y���+:#X�B^�2��t���o:9�$�tGLs�.��DkP�[�d���'F��>N�q1�����v>�l��9w�1�e���E���=j��Ι�xb�S󹍮)̂�߶|����;j����IG������-=��E��k5>��矪_rv����&�DH�M��瘴��v��vm�z�_៧w�r�n�� ��Wr��'XY�8]rIZ��򬆮М�����9h��<+��v��m� yu6�N.nSm�ջ\u+�7��h�n�ܮͭۋ���X�΋q���爻<t��s�`��re�<�b�9p÷���6n݇v�$'�:#���Ĝ�FZ�s��dV���9��^=�v�OS�"	7l��՝*FS���z���6�l)}^�`������������i��� T��&H9��AvC��cW;�j���j� u^��Y���C�b(P# ��	��fhwչ=N0��PKo�njU�����/�ݍ&#3��!���9���C�#�z � �ڵ��DT�@$ɾB��otɽ�V���!���QڇI�Q�8�,9��9'Y.�ɓ� J�[v�{W*�b]D� �����Ap��yU� �I��h>�|�%�`���� B�P|ΜWoKH>�{j7�����k:JX��$-�>�)�|�ty5ݨ��u����a2�����S�￟�έ��z���e������D�Ws���[w|o�b���\z7�''9� �������O~-;㚢Ю
?h"m]U����^;�X#׵�����d��~^�!��u����Y3_����������<g(��:H
ٓ5���x�s�((vCD�B�/w����6���w�<LhrC�]{�d�܀!��c����Pm"3ݲ$�<�t[J��:14N����E>L�>Tn�o���DD*�v�~ݞKW�ص>�97���D�Z��c�<��w��i���T4B�p;*>�{���C2Z��K��EL�Aw:�ARH��C�qQ�(�}��#+X��Dt���V]0��99-T��u�6�͎ �f"��
͟_�?|q�����.�ft�#7 v58�Ap��B�s�\�СM��pl8����b��
D�EP3�����A#lS�s޼�N�ML��C����%�������j��{�{he�"��	s@�271y��BM��ljJ�y;�؉�p>վ��u�:�INw��M��o��}�8I��a�ȳ_��7ϔ���*K�����^;�y'�K�5'hJ��Kjy��J�� �8�(cU}��A"EW���b���k΢��D��2�|�F��/G�m�3�w�LW@��<M�:�4��@>��=xl�T�K�D2��P�f�D�����#�"U�I�[%��Ɠw-�1�m�3�*��-+fڼ�e@w���b����s�t	�`��1N�k^�Kg{:��lL���'k��xl̴� ��(��n�r�80M݄�Y�皩�'�A,��e��0�<�T62���${3�/ۙʶ����/=u�D(xx��u�N�g$���4��>r�9�Y��=��ē^�P.G�t�Ñ[O�O޸@z����T9 ��铬@@��p^�5r%ù3�O���<���q�;i����/�÷����x�1���|4�����:���E�&�P�D���b���x90`!�v���$��ȇ]o��d���RH _{`I֖wtG9��Js�dz{~�!��#j^B9N'u��a��ZT�
K\ͦ��3�M��xcm���g�~Li��'�f�����̉$��s�1f��\*���i��`&��n��w��=sh)�S[%/�X/m�i?�F�Cr�uqH��b�8�O� =W �kn�A�&l�#ͽ9� K	5���>�J��
�PA �OwD{����0�	x1U`��
	`s1���sX�K�Ή�����ğr����uw�F�d�Q2{�e�:w�"$KP�FA8�e�l�D�ҍw>�O\U�
���"�}�-�)��]�1ל�z���,rE�����Y�A���@d�E��.�ɮk:���Ḃ���"V��Rxʯ;���nQ'�'�p������b�Ff+L&�vĻ��g�uR�ewk'��J�8��
-���v�e�k��2rmftWonk��3�(�6u˞�֋e�1YtK�fs�������^���㗨��eJ�hYe!��fi�c�&-��Z�#u�f �c�]l��d��㭷nm�}o:��[�kƲ�1�+�$Ж�]��ۛ3�Tq�؜�����e�b
�{Pz|v�8�u�)��7nt�����w&Y�w!�������]��Jݞ��bIy/��iB�/2P����s�J����b{�t��#:�T�n�ÿK��7�46Fg��$��w$>z"i݉��k���G��Ǯ�_��<��5`���D�8o���]X�My�$��� �?:�	kf��B��"�z�kT{e?�jؘԙ�y�A{��4�  }���j$wg���� �\C�W���%��P)������x�� 9hW����݊�bS;�����ybH-�/�W1�<x.�< ��\p��3O�"�mº�v%�v; ÷]���M�Ö�x�Ip������|�Aa�M2�wt�}�����ưm�Aeۈ�Hj�P ]�p��0��`Xݳ$@<Hν���Ԭ��k��ܕ�y[A���5���pQY���E��R��$������OpC�nֽ�Cמ�1А����igYx�-��D�@��)���2|��	n�#}��ջ���0!�*�)n�5��3�Y&%��?���{j+�|	*�m^� C$�W�@�z��|��L	���o|���O�xD�>2L0�@֤A�wM�t�������|-�iO(F�u^��!P0ف�=2K����aV�^��-�Ь�$�j�����$�k���վ��eM�Q鈇N!๜�<Q�V�^&�w8\���le�ҁ�&`�JO�~�M���J�ƙ^�ĀK	�t@6 ]Kz�3���5�3���	��I:!�U�cL�Aȯ/ltq�ٯ�ˉ:�����s�� �Ή�ki�{�`����%@�g�fI���v������E��2j�=E
�!�Qܬ]����H��9n�&9�s��HgA�Ё���[V�;��O�h��h,�!�!�Z��8��l�N�CE�5r�EB���3{UO�5*�7�Ďl30%�c��d�r�/���3}��m�d-��_;�x��j��3��=�!��O�����v��o�θ �0��i�ld�	��G��D�m<^�)�����]C&�a�5rj�2ڷ5���X��M�e����@�@��eL�@Go�$�^�-�g�؝|�s�"a���i{=���"Q*����g��;�����,�SGc�I���� ��(4������ץ^h'���\:r�� r��0 �A��H�6=ܻ0�r�#X��<(8�]�xy@J$e�fϽf�g<�3ad��`E+� �n���/����j&���Kn���d朜����D>��G��wr�0Ѷ��������z�&���	��d �d����l���<<���u��4���E�u^^d�=ı �/y;��,o�ۛ��R�h"Ar���F���x�q7n�9�8GU�k�66t<H�L��c�u���Q�@8{�h��r	��t�k�حT:�� Y�Ql�O�\<( �	��{��Y2��.U�N�$�m_($��L��M�������.���17`�a���C�E�lI ���73���o�2��z�"IWw\��Cr�`.��4A8�^NQi�q��	����fM��7��N��zc�� ?n{�a�P� �TNc`�6ƚ�����h���8��Rؖp$��C;�d�k� ��{B�<dҩ�J<7�b|{��wl�XʼFL������ܾܚk໶a��N޻��6i�ۣ��s�����>F����I��-����K��=�ri����^'�������|�x�R� `�O�݊�p\RΥ��KyN�P�{7�:�_v�E�ûLWw����fk����F�.�d�W��N�|�^w�����^�m���to=s3m���t�q���P�͈0��7��=��x�{�.��y�7���k�K-�a��v�3������G�hS}��^��OZ�\����9�
��6�S�����	|=0��3v��HC����[��O��ݾ�}J�h�ﻸko]��<Pҟg�	�=+}PgD����!9xj3w����z������m:�m.��Q�x@�N0vn��N���Gď7����V=���\�!ma�U���"�x��{E�f\���)���b)��_goH��xg��Ź��=���TΨ{�{�}���t_t>^[�7!��:S10nhߛ�|�^���+r�v�b��	&�nF�H����t�����;/�gux��<��1�g���ZZ�S|T�j�����c=�y!�gT����h��Wy���B�Ļ�m�6k\�#�Ji`Ɉb(�.=�|UA���,rrX"~��v!IE����(ЁedכDVDQZ㉌�1H��8���*��c�:���Y���������ۏ��ȣ�T
�wK`v��Ī��k��(���}}f~:�?u��ٳfΧ8�l��LeV?
Ǣ��N��Ld���#��wpr������������?u�������7�V%k#%���y��ԗ���>,8	bȿך�a���������8�}}}{{{{{{�Ig$��,�ED���eB�%D��(j�Ե,��E��|O����lgS���}6lٳfl�J�g��X�+U��T(�XVt�`!Q��.EM�_G��3��q�믯sf͛<�t�J"�|כq��[V)kb+S	75p��N�Y��Ɍ��E��ջp�Aq�H�FF ��P�3�jDb�K�53�ǧDF,Ċ1���/�\ȫ��Ue�q#ݕ�hQ�X�*�ҥ{J�0��G�QGį-G����m� m�G���C[r�ML�ڰ�\I����<)�<35��K
�:�\�k�͔#;;b�K%��<��Ƀ!&�y"�Y�m�`��n6�WJ��.��MGh�l`��ڇ�Q͸�^^�ۓl����ѕ���A���:x�E����2ںLe���*�b�s���E(YE��eke�QSD�	��(g)f�;���ݹ�غqv���^�ڞܼ��y������=)=�N�՗'����X+)P����b��EĦs���@�f��^փ)���匈�=j^dظ���`��p��G<�^a#�]u�{�H.@��x� ��ޝ��C'��"���aćX�Y��&��i�utՍ���e
�̝�f����`�sq#B\�n�W�y�Iɮ4ݣ�ul���RK�֢�=*���x3]��vr�����Δ�G7�6�k�-���!�����w1�z�.�WF�q���S�����̥k<�x�yճ:�
���g�.�x}v:7nurD�{n��ɠ�]���fn,7G	G[��z�Ivɺ��И���'&ng;��W:¦�\a��!�i��޷
)�.aB�$#�ڵMfŇ��]�F�e7.\/r��y9��ok.-�1��ij�Kf,p�HR��8��rQ�xg�{/^��n.�=�&4�<��]B�W����̲�r�`���@\Y���];����Uٸ���Nzq�"�`���;�[�[kl�;f�@��:eP��q6�X��M���]�v�[4�4Fm�5�v5]<���l�xy�� ��1�����;GV��t����ĳ���.3X�z6/m�����y��kZ��rs�5Ʈ�eJ� eՀͫ3WJm*FoWW��]��B���� ��Qn�ع��+u�\�-v���$�S9�&Nݮ�.���7V��rս�<�^���QD��ݻ���1�ꑛś�ψޡ 3当v�pXCg�9�-�#�	P�ǋ��6�ژ6����h��c��1u���e�뚺b�����U�l��;�{W3OJ1�ny��#����Y�E�/��-R[t󡵲iWm[�����#s͆�A��ܽ�P낫=[�5x#S�tpb��suz��u6��Ę���ʤ�e����o��=���-ۂꞷE۠�mڻ"]V,l����a(��JFgTbˌ*����yjtq�R���\�u�lM��K��S]�HƮ��](��T�h&�X���ߓ�~���K߿�0�ÐI��D��>�8;&�Ѿ�k�S��@���Nׅ�AxxTg���_�kj�8��Ÿy-d�>8�/0�5;�ީ�I�����{2��R��&8��KX����xu�We�ֆ�^���bI��&�G�s�]����";�$k�%�������x/4M5��[dM)��>�	3�#YAgDd����X�`_]�u�}�LM����藆��w;�X�Y��	ݧ�m����{��_e�2F�̰�,P��(�o��ܜ��JG�(6ƶ�IK7i�U�v�;\�`���ZcUY-��j��>���_�:�,�רn���v)��O0g	%���  ��F��e���j�I_D���N�����V��3�Ϋ�h���V)�ݹ�t���S��8'����˸����&i�O%�\�'���p�^{C�׽�+���ѿ�$�&!(1���$#�<�Ա��ϓB7"r�=1�T�/��$��7�x�P�)B���'܃�4���wʋ�U�`)�Dށ��@�W;R蹇�8֮�ɚr,��j�H] ��B	w�bZ��?�$T�=w_���$��yـ��@	�$�vsMt����2��_<K$	�W�5��"���#��H���������<��s<\[V�Qil[�뱘饰���n��A;Ä]�'N���1#�
��)���rY��,���=B(�yZ��^�O��j���ؓB/���:�a�D�fy�T� �޾���N����9_)b&���U
@'d�.�'��Ց����j0�9s"��Ic;�I�V���u>P|Q��W:�=��,�|�"�++&dV�G��ꈇ4���/.��ڋڥ&�'�Pt>��Yj�;�z6��C*��`P��~&�E'�*Kfw���?=�ɜ�������;�w�0�^�ME����]ߩ�[4�10�b�v̔�b��6�<��.7A%�j�U�����<@!č�A���o�Kƽ�=;���}��X�=�� �_�D�E{��.���̼"}������v�T�	k��r+2�h���&Ֆ��?����D��[�T_��̖�Y�Q)��@/�ҽ��������)*��4�9x&U0=}&�wo=����2��Ԑ	 ׺Z-�1"h���r���j9��9؀�@�"dy�_ �F]��6d���H0�=14����@����.9s P��*.�	he`[�I��,��Hj�S�aJ��#�1��^��f�R[��yŰ��`�@k���/���CgUV]�e��o�8�|��5ݸ���t�D��W�<���Qy�x���yט>_��/ۘ��َ�{{$�!
�;G��F���a�}b�ⲋ�CC���;��?�b]�\Bv,ڮ�t4t��B�����wz�����u��@����t2vtH�	�+�rw�CMŹ'��]3l�u�,�ś�%o��^�j�p�"b��$Bx���r"6a��� ��)mmg�*��ɬ�ɻ��͐H���U�"!O#�0芔��$�O��cƯEoEd�vAk�`�-��,�cryh}�a@�T
�3+�m�R!zL2��%�X�� ���y��mO@���}�����DU�59�� ��Ap��$��sN��O��5���A�z��N��BX�ǠK��m�O9~���pC܌z�w��͖��k��4J���M���Aq�w*�t�ͼ�@Y#R$� ��?S�!�
���s.�%�θ)lV�ri�>6S��c��kq�=���V��.�46ْ���c��0�{k�7���]{-ڷ.�G��Y��Q��Y�`��MWc�Tˊ癴]{*�rb�!C��a�Z�I�]�m�)�v,�����#R�ڲ���,%���'��d�� ���t[���a���G��g��Z�W��ϋ���v۫/RFz����Ҷ�ݷd�;��]:-n���[B�����~�[�M�E�4���@�|�i�Ƒ�@��bN��x�S�\�;�vƵV�2]�������$tdV�� ��z�������^"$%g 1���S �'��7^l�x�>���p�"ȫcG�I5w��X�<E�'�>H��۬X[��Am��;y>X�L<�ݑ�پ�����}��!a�{�D�ƻm�c���\�擔�X������!�P#.�#H�c��h������v����L�I;�}�&a�n� .��$(	ܨP���DhW�z{g���:�9�7m�Z�k���,Y�����$��ue���M�x2
�މ�O���)���,��6�x
o�狼#!d]� ���&e����o�C��;$8Ɯ���xq�&6�e��ٌ	��Ki��X'o4sχ�1Gf��3���>;�|��ҝ�]���F�I@"ή��N�}�8�����/O���+`_'���]�=6臇�8��R<��� �^���lL��� �v̂�<ll������p�z����:�͔�cd.�H���(�Th��=]S,H܎P�L;�P�^�H��#��k�	�I�d�]6ԉ�2˺D�D�[�������<�zE99ć7⺪�]v�n�-��!�&ݻ)��۩RW\(�`]�w)�H$���9�� C�5Vl�2�=� �N�� �8�q�x)�䃩WD�E1��C:��h}E<�D]�J[u��8������w�mW�;В�E1�H��PH8=70���썰r=�py�q�.��bUl�6{r}w��E�X/�c���w��$DT��k��y����Z�����+~��j5��Y�fUъÐU"�1a��0��4�ʐHb���\��Awa������s����x@�.�u\����ϫI<���D�I��P1�${�f�[�=�W��}G��+v0�Tب���w�c�^�y���	c��iEot�M�?���N{�8V*q�����`�G 򶇳�4�c�۷	sS�4��,f �P!���{��D�FG���A�$ϼ��"'ݓ �O�q�Ǽ������r	&ڻd'���s�:"@���3"&d��dg�������>�:>K�6w�(Ej%��-���/�!����=�QQ�DH��d"	=��#�V�<x���b4+~0�wL��sl��xt�Ȧ�L��\[ѱ<k����a����ЇvT�$��ŧ_OFH�tݓS����''�&;��Pw'z���O��wǻ�藱�y:-Rw���xi|1˔D)&L����F-�Qi�'�Y�Ł�i�X������C�$8�' 銍�.���ǫ�o}qCyyv(���2ot��?r�{��@�Kx���]���orOS�j5��ysYT��rc�vH/	�ٜ���"�M�Yހ�X�碈$�����P�!6 Or��k��Q3۽d������ͣ�2e���Kl-�,�����A�'{���/{�)�F�!U����:� �I=�Y�;�I�^e�j�	�A�<��5��톂����bJ!�D�tֺ����#�;)�o�A,��?����X��铬8���ޱ����������3�^���M̷��"@#;"�����f��Z%s�5@�+��)p;�(-�uH�=\����0Bti�b�{�e7i�>���������Nu���V����)��9̜�c��[���7%˲q���"�'i�|s=������f�Nl�S�x)'��]��u\��>-ŭ]cF�+��s+3	y����m�#`�l)]�u\B��8(z)\��������vN�����::at�\�T�k#���%�y��v<qf���݅�s���k�5�*,1�֩���x7pC��]�b�[�{o�ڬ/Id��� E&�vGOA�:�a�et���2曊��_ˍ.D@�lz��$	vU�8�d�?��^&(�}��˶��A��ǧ�^Ĺ��!«�V��n�X�'^��H{<
����Ky�ēll�K�1ezG��GLΊz�z�w��9��d�s9j�a �+�$I+/=�GW���>c�]�1��~#=x}Ϯ]B �P7Oq�� ��x�<��9�n?8�{��9^u[�#j���x-J� ]��X`�7�	�����;�G�� ��d@v\�ovG���E{�]�������P�\!�:����;�\˭���uۮyccUj�a3SA��58�A,�O?|������B�|���������}�
��*���� �u?��W�a9��#y�c.�0�1��Ӯ{�#k+v'��{�ל�����'o��`�n�1�Q��:p輋�����&�"bfk ��3�-��
OdLϼ5�Z-�?ud��rH(�`��O�Ν��tz�^GD�3�w����O�Z�>�����tM���7� �DV�c)$ow<	n�� ���i0�h��������0&|��{Z�n�w <�1��޸�5T�2Mݟy��O"�fA,OF�v��Vd�>��É��pKo?��6gu[@ ��C���+���RTB���M+f�bhėR=m�#s���݂.����K�q�ȇ�v� ��"Gp*�$��d	$��/s
�K�aDu�[)���W��pjxpa�.j�݋���'�|��H6�����d������Q}����W]��`H����H��Һ	%�8��_x��
�n��k� c��ܙܺn�V��L¯��7�|�>Y3�voYazB&�1{y���a����<�Զ����qb5{;I�]=�t��ո����(^�՛Ӽ�]��zv �䭝!s'�T3qKd�Vh!����ӟ����7����Q�E����C�x*}��G���a�̾�Kt緗y�vn�����v���������v��흗��E�����sI��Ɇ�+�	WU����ފ�P�����L{B��4p�t�� k�w+�z�v^��F��q�zt��&����˱:[��+��.sI��
)����;��gV��#��+*̹c)��a��ݾT�H�xi݆�|���>��L�v�+k÷�0��\�H|FC⤯��K)b�/v��
�b)�qx��9�s�/�_D�`�e�q�g؀�U�P�b��&;V[��w 
f����OpYw��G����
B���_2ĉ��.݅1zӿj�[��h�jR��AG���O���ّr�p�M�Ҟ5x�B�R�^������2�I��]�7��<3��8��ۛñQ��m��r@��^\yq���ƣ���Ĉ�yL����>l���:^q`2@�xɹ|�]	/2�D#���@X�%���{�a>ıg��$:� �E�ī�"�Hx�?@�n"�1 }�^�zd���$f!�d.x����{Oq!窖	�'+�'�T�u��DEpq\��C�K����xϣ�n?����������d ���hV�$�Ey�9'��b,��商)_���c;'�g��w=�O�͛6l�yj�¥E�R���Ď�T���R7�p���8a&�~��g����㮻>�6lٳy�
9Յ��aTJ��c�@�H��}	 v��b*���������Ա�ٳ�u<�ϧ�f͛6l7����X���f1����Q����)��lnz�u̼���z9�ۯǌ�?߃����}6lٳg9"�8�6V����bc��*�
��s�������G׷���׹�f͚j�grҵ@cmjq�,Z���m`�XYf*1��!��`��7�U��`��+��!c�ܪH��Z�	�X8��R�˄˂�+6�.�Uk�cS����9V�: pLD�`rr��-�*�*"�+�5�)���E�F6�Ir�!XV)�,+.u�m��Ԝ��@��������!����q��L"�-byE�{�(�y됍��59P$�M�bx]�����WḺ�x�L)*���,���J} �xyf�Y {V@]q ��s1ء��H-MA�}��4΀�\e�]�]�������<��h�h��	���W�>���yd�nof�A��L�0Y���(@A��S7�͎l�s�O� � ��4�O�B���Tc%����..���c� ��.�R�$�nePU�M'����G�۾t<�d��� ��]�8Z?y���f��	�����C�8!؊��I~��Yl��H3���OgE4���QK/s� ���6�E���8=~��;^W��2��òb�{Wo{��N�v!����U��/,�S�UYu.�o��f=h���o��=�}.d~�2�!w�]K���o������[IRp�D�H��d�A��Z��!��" <�l�U��B ��ȓV
�x����s����-��G�V2c�RS<N����~�B�'o��nKt�̥�-��n����)�絫�\�xO����N%�.�}�)?a<<�>�1 $j�D�2na����!���r� ������4z�d)��Y�7F��� � ���H9��2Fb<_ι�un�Yw�GV�x'^�H�.�Ct����
_��MMe�=��u?�
d���Y����������Mz���cޑ�a�/˓�P��nI2x.�u'B�S�Ɖn�����膈&0$]�b����K�b�h8e^�S�x��~ ��|0	$M^̜�Iw#�s�ʋ��w��e�v��qv67U�2s�w�'��n�{��O���פ��c)S՘�T���!����t�/,�w�hV"��9h>�ɓD)�$0���y�bi�#5��3A�u��Al�u�xknv󍗻"�n�٭�r�<X�l"z���Ǭ��<������$C:޲�`�֕�A�nI�A�q�8Gd��VNg����ҥ��q�5/��g���w���|6&s�D�`�ۚ�^�u���7�5�����釶�.`�m�R���=U٪w����<�Ah�k�E����o�3�c��mu�U$WQH�3����vc0[fn��؋�ݮ��)!�����,s�bI$d���9���Q��~4�p��Dg��$��ٞ��C����U0'͹�������:u�-�9�|�/2��T� �D��CEq�,���q�K����K������[���lV��;��sܷٝ�a�$����`Be��9{�O��"h��A��E���{�<�3��1 ��TH$G^�e����㫂���q �r�:�N\��D�a�}	 ��B�'f�uO��Bw�H�͙-W��Ko?)�}�J?l��o���5�O�d?�M�Q,�'']�N��J�n���H�6HB�=��"�hˀ��\	E������A�����#=<z��Ɇ8ǖ�,��AI��+@=p�
l��:|�zIp��pJ��n5i6�|֍�k���� �;�7f���ܝ�Q=*�N��k�z�H���>E����$"D�?w�7�mY{���?{����^��j���Ҋ��xxP�L�cA#;�.�U��&+-{�c��u��0ey9���ຈ�	)�r���ez��30�7� �A��M`��f(�$M1%�A��ez�A�=���>l`��1M���x�-�h���4�����2脖h�I�s� �^�b��7��3��/�թ��9E�A�9&��%�'Omײ+۶��k-�6��+V�K|>ϩD@+�3R���d�v<H���)��o���J�!u7L=�[bB��	�YV�bt�!�3}�<��{�Kɔ��ޚ2G��"��ߺ$&�v~���I�Ls�0D\z�������ۻ̷I0�$WY�>�s]#� {���JP^󛻤�[qj_�IN�R�z#����͡-���>�oBjZ���OP&gyڊ~���)��<I#s:�C`�
E�5Ѵ����0���x$�H�f̏$I��W�1��4��@��t���>8/D4ҟze���0�G����".�y��۳2�ۙÓ�]u��#�NT9FAv +���e<��7�eܲ��g��k��x�)ѿO����臈N���V<A,v�"A`Im�^��,A"��e �{w�!$;݇�;�1qB�+2�xA�����դx�I��F)�[��	�(���/wY�N�)�A�$ H�y���[s;��x"c�>�Ngh/B���H�z ��h"67m�~D�&�0�P=ꍚ���	�I�!�%�s�~7�Q��H:@5���܃?�9fN���W��5dt�^H��D*�۬�m�J���~!�bHWr`~M�0���f~��r`�G�d��{� �	A��U-�'P�	3��U
�
"�'�:d�$9��C����g�&zN�t]ͤ�:�����][�0��q�z9��O*Nt���0����� (�-�9�Ļ$�a��	yq��������o�fX�&D�z��&�x�xxsT|]K "n�\�ý�72]`8č�����@��~-O~r�.����ǀ^�42�� z' .���eDN,�S����+D�v�s�'g+U��:H@� 銏OM���`,}�< S�I�ߍ��[��O���6��{7���<�ϧz����a�3��b�]2���K*e���Z�D0@-��y��,��uYJ�&U�P�z6?'�M�>
hL��g��-����B����ln�aGt�+���9%q\�j�cǩ:��-����u������+�`=?�������wf�.��
�]��!/l�d�H5�]�n2����Sk�u���9�Q�WY���;Aq���5V�;FG�Hnv]v�;����y��nwK�\�i��cĜ�`�[m�9:�S#��i1��7:X��0��F���cbzwL�^�;e3���!=��l���;kB0�h6��l�c[caNq�q�X���Fڂ��n��hvL��8k�i�lK�ڑ��E��itlf�᭏�=���	A��f%+l�q��/@D�}��&�5�Q�v��AM\D��r{��WG�p�<<D+��L�Jy5��jM}�$/���i���h���eE��'�<C��sw`�٥�l"�@�mq�)��Q]��X�+��M�wUz͎1T<*���\k[8K$r��2^�ؐX��n����'�hd���PH��:�Ν$ S�퉑����� 8s}s�]	�R`$%ڠ��$�tD�;�a������x&!�V��m<�`�s�������e��dN�X@�	7`���/���.��!?KpTs��Iמ�:�2d��{�f�5P�r�-��v�S���)��4g��'�_!{O�Y��M������y�m9�i��6����po�G�����H$�üS�Y깅������	���(ɱ�������d�\����������F1D
��Iu{�₺�>�����l8OD��a�dăא�S$9Dg��R�k'%כ��.�LI6�w@{��t'�a@�V��~��Dv�$��3� <��^��1N1zl�y�I[�pix������zH�Cl�����DLfod�l�r<��#�R?=O��~�?m��7f�56�lW�s�n��
��`�Ŏ�̮��4"�w�~��.�j3O'�{�G |�|��I��PJy~w�����<��ʣ�2�zp���!z�<�*�$]�Q��n�p��:���z�Y2C�b O.�>_�z�M��N�3��D����<)������}��K �|ʽ�8��ݽZ��A�����r6I!FN��aH�TFA��(��2��y���p�D^䲉��oH�~Ͼ���fTO N$WdBb����1f��)0���^QK�{������=#-K�^�ybIO��K��v��;�*��y�K���{��Nb@q"�Z�D�=yg`����$T�@���8�~�V�V�T�w���~��D�������EDt
sun�9�i3����;�.ō�qHZ9΃A�������Q#��P��nv|�y_�B �g��p�z�`㽦�S�"ܼ`���W�˻� M�ú�gY-d�M�y]]L4�e�Zq��8��tKȠ@���W/J��[Y� ���S,��<��ŧ��x���{�U	`cܺ�I~�K�p�U�tb�N`9��fV_:��'�-��Ϲ	$�ݠ�������ʿS��:w~��Gxn����z��F(�n��c=�^����[n�i�9��o�������8e�ĩ� U������_�=g{T'�Hv�j�d��Alc�"7_H��h�߰ܼ[��;B�M�@��.s��}�Nd�<r�D��7u�U�A9kp*��҅���Ƅ�{���~��GT�w���J�=�4I ��DE2���|3�j�n$�%�{2$%��Βm�b�5d�:i��z�Ω�{Q$�vD�����!�����>S΁�$h��+ 9N�M�=-&�� ~鼙U@��g"۱d0���{� �ɵM�
"
�iO.���z$�E�A�;�Ac���[y������՗D���5�$V��J�LC��c�ڲbZd��d%��h�c�d:z������{�}����������࿧8��A@y��PS�������*�� D9�=GD� �0��d��!�� V$�	@�V @ h %  B $U�  !FP� �%U��! !	 dE���P^q�
�u�!Њ��!�Uz�C�p�J�!( u�`!�"�H�!*(@�	�$@��!" ����H��q8*) '��*%D�! ��!�!(�! y"/ BD!  B%  B%  BT U�8�	@�@� �P� �P��*�!@ BP!@ BUX!@ BP!@ B@$@ BD%  B$ BP	@� �	@� �� �d@!	Ua	� �B @ B!  B   BD$  BD!  � �	@� �	@� �@�V   BX� ��q�d>A�/���"� ��*TA��C����O������c�s����?���� ��#�7���������_�?���~+��@�?�����Ђ*�G�@b�_�?��?'�4�R4���~��C��P_������������z|��?�&�?����p�~ǀ�*��J R�*���(�"�$HH"B
��I�H�&�I�H�heH�"U(� �iR�!�h �%�I �)YR`Re	�%�I I R`�!�hFI!	�e� �e�"��"���P� �"FB(B� �f��f��$�HH`X`�%`�%a�$dH H�$a��V�fQ�$ZQ���f`$ZQ�VQ� E��bQ�RF��daX%H�d�`HVHFaXB��Q�E�%IaX IB�I!X!�Q�E��a$ZQ�T�	FIFHVXFU!Y%$X�d�eT��Q�VdY�bE�X�eE���Z�F!Y�f�U�i� ���`�b�Q��i �RU�hEH� A "����#H����B�JK�B�B�J�J�
  �"���IV:�@�p�������� ���
PP !B""_�~��w��o�������;@��O�}�W?W�P
 ��??�ÿ�?O�����׉�'��������������*��?D?�?�����@���T@O�C�0����};:Q|���BE@t'�����k���9�B��B���������Ӳ���0 U������C����� (��S���>����p?����;�����������`��>P\~�Ĉ���@P����)?z�����p>'�p?�~��4^���}�|�<@|L�	��?zq��?_�:��}_��?)������P�_�q��� �������������~����d�Md���x�f�A@��̟\��|X=@h(��U@i �� օ���@�JU҆��"@$PM�� H�(�JP�$� }
n�Cց@SCl5@  R@U
 �R�$  (T���(�� RE	 @ PhN�                         �      �  �|  �      4����F*'U�
�4D3��"� ������"�s48F�tt�n 5ѧ694�9�H	Z�Q� ��]fˬ�Q�#�c���v�jf����{4����a��u���B�<o ��%@hܰ{J�7��:{���7�h�)=n�޳� �� ���
   >         <���70�ޱл6�Eټƀ�� �h�n��TP�Z^w��z]��Zn�;Վ� ^a�=�:2��o5%�\�U.PuJ�s��J�-:mR�B�^�   �{|�"���J9� ��VFvh�t�!RMj�t���H�� �N�s�4�r�f���'�Ǘ��m�B�H%!E�   >�      >� �*FZEO�WZ��t�K���t:n 	�JY�TP���%v�[]5JvSp #"Ws��ت�gV��!��   u��)ul�ʨU� t��4��-�R�i\��Z���ˡ���.�:�'q�e\�屶���F�t�t$h53��  �   � � �AӨ��nΕ;�l���Ҏj��7W�';����[�#WYҡV�r5p ;����n1�s��
�}�  �!����q�� ��m�F��`�+���U9ػQ�w@W'\�V������:��@�AD�� � �      <׾�]뺋F�������]F��t5��ەu���0��u�Y����f� �͝R���� 
����  �����A(� ��V���:�u�B���uZ�7 �V�j�[lW��pu��΃��OF��RJ4ɀ�!��D�T�@h2d1�ʩL%5@ h5O�)��)   %?R���T2`�тME0� �b{���U�_�wg��c��j��O����3_ $�	' K5��IO��BC��$ I?�B��$ I����������ߩ��څê��4Kn�=��d^��J��˖��V���4ּ�$71C�ꗪ����*�Z�u��f��%n�͚���7Gr�A�I- ���
#3!�oqi���aϐ�L�կ_j���e8ܭ�4�L���!����T�/h���5���q���{��F�>$ϊ�����ʨ���/���GJ�(ˈƭ�
;I�y���Vdj]7�рV�Paz�yq)�U�u����>�R�DR� 7¶���������F���Zf/B�a�2�ڕ��&�n&�(�b*yM
8�iM��f�y���97�$
�;>4���Аɑ`��8�,R1A�v�ٓ-��
(L\����&L�H�9���w��o37�������e�J��!�U��b��d�9��ilq)��]3���y���!�N�ݳ�;9t6Օ6K̫Dmmτ��C�N��k�m7Q�e�ɔ�Qxn������2��ie��
ʷ79Hg���	�w(B�ѽ.��چQ�.�^l"&ޢ3��ܓ�QK7#X�1��u�EWV,MzUK�SB��Ci fMR����y��0q�Zo��otf'�^b��c�(�R�6�o4m�N�3%e�.:�*�uލ�b��RB����,�I[�b(��q���f�!5�K0=�2��+]'�᱔	K7b�P�i����`��b���gW�Qg/ w�]���Q�FQQ5�R�Z9�P�2��ɰ|��ܦ�Zg2ٹ�չ#A��*�L��y�q��2�j���Y#P�'r�I-m-�{����{�*Z�k3(��(��f�F.Ӓ��a�vݛ���u�:�-◸j4����6(*�˭P�ڽ�z	��7�s-�-�!�Y"��3����T������E�D��GskuY��K>�j�Z�V3��5�h+�z�(X���B��0:+w�ɔ��n<��i�^lO웙�Jr�Kv#�b31�F΍�o(�Wj+��K�Y�*;p��	f�(GM^��ɛ��N⑹���zozB��S�Z��$�2��i��&�ؔ��	�f�E��\�E���"�EL���$��Y&T�S>���:9�u[�5��4i76lЎ�K����K��5ʎ�`�b�Sf����P̺�I@�������d�%�w�1bdȤ�Z������@yQ��a\9b@����fVnc�%�F����(��2��v\ezA
��ε���G��dN��j��SsY�7�5��L�v�鵻ȩv#Ш6�1#ck	�T�P|�Y Ҭt��"�`������駘سRʱT�U�֖mĉJŜ��M���Dj�rb$g4����{�{s�qs3&�ތ۳.��E��4�刍:�k^4�ݳV�c([u�M�Ra�Z1i8�L[LC2��X�U�IK~͆�7Y��2�Y�P��	��xD6��PS��k)�����^I"��3���A<��օ�� �j�*�S���k!Ub�^3�r�ME{Y�]�m�nXZ�Q(3��2�� �
"��39uE'	�&eʳB�M�ʰ	�iʕr�ݽ/7�^�~ژt�V�q�tjy ��
��nf&���L��j�_���30Nd��l�2Ѷ��$�Q�L�
He� ʊ^S����J��*$���EWR�배�+�15���Z�H˒����4`Q�ڂ�Fo��*KӴA{`ٷ!XKU,�Nc�2>������}s�b6r<��)eLgkY[j�"����sa�Z���83��S�^Ė�m�"��@��R���*`�d
vh�i�ӟc	�!)eCZܙx�.Y�x�J-�X�el�)V����!ҡܚ�ʹ4&jM%��9"`�lXk,KP%`���RSPqf�MXзM���I[����ot���Y����uml�+6�yLYw��"�\�� [P�I�V���;��5�UW�h�a�T,�pK�����-�l�F���%!+t]i!�\Y��d3N� ��+$m�y�M�6��6��&[�-�j�WB��frM�vH�77/�S�VL�P��'�u��ݸ6���ږ�����oc74hӫh�å�s�"�ֈ�Ѵq]��G/�ᅳ��g�(%��eB�]�[����lW(���ˬ�3)��nOA5"!N]�j��P�A���������Z�^KsX��8ѫ�iӯ(Z2D��e�-��QͧR
۶��O농%�ҳv��|)Tp�*�.໐�.�x�ah���s`ך�W�t7WYHǷ���\��cJ]�N��OMndv�N`��@��f��O׭(�i9�PK*�#SeA��QT8k+M�BY�W2̦� S��2�/�љ��[�EL���h��ӭ��O�{Wy)�3a���ŉe����[%�jw��������_� �+v�ȩV�ˋ64�Bmj��:��$�J�$��!�.���0餟��
ŵ��5+*T3V)U��+�B:�[��+Z���l9�3a��(�[0;6jڨ�Ym UE��������iC.-+�,%M̪ �{!�©1���`�&��u�Q�Qd�d�O2�b���.*7��ѳj�U�n�����U��`���[2�f�^:��tK@$-J)�ܰ�6t�A�w �n�<&�u8�N��JR	��ȥ��;�pZ	��Х�7u���e�I�[t���P^�6`�V*�^MѴ���Z�F��[�4nn=St*����4���xww/E�n�ܵ���l*R�t��[�"؋6�ы7��2h�|--W�7v�[ͧ�*Q!����i�r��.�-l�M�[���=��a��n1z�Tf@tf��}���#[��2���Wzӻe�u) lX�"�is��e��B�kid�n��G�k�W�$m��
����`�Ʉ��)5���ۄ]��EM�$0sJq]z��N9n��3�jiؙ����NbOMk͒�(�������P�	���͗Z��&	GU��(�fF�f�U+�7�4���`�X�a5����;4s)�	OkV֛��i���MniЅH�m2E��T���NPz�	�u� �١[M�6QYl=!R����pI����ಢ�~ZDg ʩRѨ%n�:�*fTD�TنW��WF�L�
sD��R���k{XMק5�r��0Y�dȇ�j7X\�eU[`���j�*��q��C���N�K��xUm�ԋ�[Q�Me���_+����Z��f�킐���Ӻ���×/uLN�ܧ��DE<L��2NJ ��В���L�sj�ͦ�&N,=�1�˄�w�ˍZ9�N�̭.�2�<��w@����t�ȫATR�:�=,^�d�;�<�ZY�efX	D���Ưe4PfS��1[(í�+4Ă�E%M^ZJ��K�i�>t�k�y�,%��:v
4.�+*\H�v|��'�idԚ�:���n�=NJ�Gn[�.�A۬��A��x�Q3��Pō�L�8jn�X�j�8E�L�����l�:LC�Tniu738���;*)DG���sֳ���bMK4Y�	e�tw3oZT�*���[e�nJ�F�B�j��S��Z�.j)�FHR�CR�M�X���槵c턌�֚��
7�m�����&7A��N��X�.�BZq%��kw�OKYKw.�0n��*�b;vLp��Y�'���	3ٺ{e�RqAr�\�,lE������V���BÍދ�;�Vb�M�y��<F��:ʷ%��Rm�0D���A��Up��B����L�`�3>ɚ�L���2Y�l��^�i-StV�(b�M�I�e�y�X��.S8�I�h{biӥ[r�SWM�h��-Q��Ɲ2ڈh���Ō�u�2\�b;�z�&9��7P�6:���/@$U��b��aY�ȼ0ؒ��6Ps�[�їAޓt��-��+�3+o2�ŷEJPk���B����+%8���PR܋�8�l�=⸤9�.q�wj�T�u>ۋP��bZ�:�O���k4F�۰/3ʏs��f^�.PA�fn͍e���ǂ�5'6Xk�{b�c�}� }e�I�]K''�E L�&�M���	�T�'I����M��z�8��
����Խ-VOZ��W��;[�vxQՃX�F�!T��%T`��2�.�U
raظ�5 �(�@Y�59�XJ(�&%{{�#9�U��h)�ZE�|\Z7���������Wo�MS,C�2�P�p-z1X�+)ְ�ĳ.�m��*�� T�ʴ��h��IV*33^�J��E4���F�sN`�8�j2��v1��+�ibb�[�+���U��M��E���rnm�������t��n^��X�pbz�`�Eq�����%d��4+pah8eZ�IX�ݴsq�4��Fŗ2!Ãp��n͇�1؈�Ū%2L�TPX��88*�6D]�V#��*^[-��M�@�B�e�ve�$���8Ŧ�̓F�� Ҫ͙&il)!ƶ�`��z�,(��s3�L\0������t��{F���su̻:�fS/v:fZ2�'��9i��)��]���4�K����63{*H�Vm.�K�i�[���a�♳|����[*�����h��6ʥ�!���@m(�h,��y3~l6#����iS*�j�fc*ж�NPF��ԁ�`�Ad�*��!Y�tvG����V�YJ���E��04J�קi�J�ʆ�fn�B����PlHR�L��2R��Ō��d�SMֲ��|Jv�Xͻ5��u��Jْ�q@�+�qޡ3N4�٥Z/j��-�iÎ��f�@��yr]'��D�j�KbC�0�;�����r�Uorؽ �Y5�/�s₍V��W��7R:%Z������YGD���[�ջ	��n]H����76�D�F]�P���yN��T����&�8��j��vk0I�SurJȄ�T�aCf��̻q��尛��N4���Q���Y�檼�$�H��W�!���E�H�RJ��e�gq�4��U��)�$�b�:�*.�m��V��N���Ka�����A�ȵ.1I��i�+	9�#V�4�3N������&&�FK��]�)�˃p��]��n�h���u��*(�k>��7ñ�ՙ�kX�t��Ӂ�����R���L�@�R:),�kƟ���H�s(���H� aC(�yVd�X��r����M�d
�&n�rll��"m�5�K�jSw�>��z�t* ��N���1F�
٣q�٩�\ԥ���թ ���r�!(*��/ B��.\����@��cʼȴ@�݂A(+���|i��:v�,А�ܩ�����VKp�*���RQ��k2��&�K��gB��{�/&�9��f����©W�q4mA.��oّ����=�6:wZ���i���ZȈ�y����K-����ը���R���s�i7`��F�<��VB1F�tr�%U��+D\���Bq�2�Wv�����N,N*pE���nfk���؁�Ǚm��\:[jT�����(U����ɸn�ܻ�����!T���,�y��4�5fJy.��C-��P� �@PX���Ė�m�ո���6�G�m/1ѧ)�ו�cM�`����u闹J����Z��S(�OoA0��7K�ǨY�DB�ZȥSlf�q������˧�N<1�v,�w6��d��Mj�}s,�7�D�r�AckF0���W�Q�&R�z͵mf��hЩt� �����.ݓ/Y����0ᬘ�`j/m�0Q�&�i��cԅ',iM�̛�JNW5PɻM�D+�n� 9$�31Ѷ1`�r��i��+$�f|a3T��>��𪨋2)1u�f[����[[b�����w�v���-�W)j��ed�R��-鶌�[��M+�-��hDM�t��P��*���3F�[|�Od\�k'1�ҙM@3t]Z�P�����D����3i�.�f����!dԅ.�eқ�-q���m�Ṇ�3'IU۱),�#��`ͥ)m�׻��3�Ta�Ncu6�X�;)���ͫ�@����Ed�R� ��M�V�0M$�ޯ3��֯C|��`�܇1\��^��{�N	`n]�Ԛ;�a�Z^]қV�]�T�Ȁ�ol2#w)Q�`�(�&�m�?��� �B��7I�ͅn������,jcf�D�.?�����J�*t���j�c���H�Q��u��U̹%��?����3P�ӡ ؉��ꪲL�O��7�Ft]�-d:3s)R�y�zş�
��i��%�f�"��r�L�&U��BcLʄk�3DY&0� �Z���.�E���{��ٛIHf�n�M0N����g
I^��,S�u���$�\�6b�Vre��)E�ո$�4�3v�V�R�f
�ڋK
%ʓx���;�)�#d�R���ҵޙP��-���-Q�pZU�r���2D�/&��D̜��,��.6���Hp�Vl'I7w�H���[�J�ow �b����̓5P�f/��Pv��Y��V"�8b����.o6Y��++HU�Q� ��!�.�������z^]n�!欼w��Ϣ��=�tm�B` cV��]fAV٪��H]��w{��W�)V���^����¦.�"�U\җ%������$&D�Z�S� ;��Ӱ��C.�ҭ���i�.*j����dB��b�bl�pt��;��RwT%0�Ӎk̨�[�i_��jF�sYqM `�R���� 4Ν-�wgn��SQI�T�)�f�S��2\C��L�Hw`��#���y2ϖ`���,�M:8��h�!��ր5sj�5gr��V���6�!l8ӻ��\z�;����k̄�,��iВ�r���y�3����D�'P �"� X ���I,���,d	$$$X@@�) � �I �H��B,���B�BAHEI�$ RH(S$��)B��L���R�,��H�RI$$�� ��)%$RI`H��
B �!�
Id	$XH	HIB����B,�B, �2�
 I-�G]v]u�u�qwwEa!)��E���P$�B BJB@��HS�B(%2 B�aHR%2�$�$��! ��S#����븺��軮� �0���HB,!�@�$� R@?� ��x{���~Й����,,�Q��F]�~�@���7���gtU�8/֖�k��k#+bƤu�F�͡vMe+Wbػw�eC}rns�n��Z�Ҫ:�Q��ٲ�h���\���C7aӰ�@f��f�\�zc���Ǩ��øO'3l��.��G2e�J��r�����;d?(����8u�Q�l0�Y�E�Z^^�\�h�WU%ޜ�8�V���b2˺EK����u�T��T���<�m�����ҷ�q�z�t�vA�+�T��r���Qe�v^w.5t�ݮ��ڻۻ�WUU�7��;2��`�;�gn�yrL�&YwK[��+Y�Z�9��(�a곪j���%C��*ゖ����';H���'`]:�ظj�7��;[��5�R�]���j�����o����zT����E&�Λ��šjq��Lz�B�s	ERc�tF�ň3�9R��w͏7F� +�LN�]�gnk�m5w�,Y�fP�sw����RxN���;ZA����{]��w/��ck�R���kǼ�J�pk�Ӿ�[����wi�
t5xd�Z���a�+N��aB��*�l�V�(92�î��VC��ԕ���#Av��}�=]��5�6��=+�M=dJc=)un֐�9��ЬjZ��qw�׈��i^��ooS1d�$���L����������]��V����VNe��6ΉL饓u���Rlz������v���˳��w9�y4��K�hw	�m�Ht}���B�R�x�jʾ�T�U��f�S�Dޜ��t��@���wS�в���b���X}��v嬶߬���k�wo�W7��9��w�ܔVi�N���o6�EBR�cЛҌn����F�{�m^��۳�>�7rb�M������eŜ�;�wzorm�F���tS��4-B�sN����3�u�[Y[2�Y*�dfj�BF�o��,d�<�Ṗ0R�کKq���`s���qN��<�,�g�O�1���{\��0��˶츔Y��r�mj��2)�f�fP�`n�k^�����˥��meE�T㚫���v9J�g;޾�諂�ދ��A�gC�v9�x����*�$�6�Kp]�v;�m�;s��8S�:�A�vF���Ⱦ��g g�]-hZ5�vZ�sg!Vz�guMaoV����	��c�F�����݆��j��T�[O��t,j�Op;�g���{Wye%3�@4��ĭ#u��G����`� h�o����m+�t(��g%�8��r��_oKhU�jy��.Q��/H;���"��˱U�p��G�f: ��ۦ&X̾�b������0[����W��ni�I#�r;]]kU���[�}Ԣ7Ԓ��o�d��oqHq	��(uҔeV�635��U�엣zm黨 9�R���ႍK�	v��0����iY�3����e��mVP��[���ԥ�f�5�ҋW��[���,�TveT��b�Vɻ��×�͗�kU���o/�ٮ��B�w�Y7]/���;�LǢ�Lb�
 m�ѵm�MRj�p�1mLɄ��2�� ��c=��i���*
];B��仺ٱ���5ywwف��2[Dr͝�� �3��|E��[f�m�٥�&�u��V��̖��9��Ml�5�ݥ��*4þ!�J����V�Г�R����xJ	���Gy�[p:�ټ�C@�2���Su���[ưd��)�|#L|�o�X��i�w��N��ڱ(gCh�쎕��刎�+�f
q���HFmϴ� 6.��m;��;oA�z���.ux��pKܷ��ۻSJƩ��\}��)੫؊Z��ؙ�T�w45�-�t�wbym�s�FX�;�f�/.������7��Õ�-`�2Z���+�}�)��۫pP���+�S<n�
Ղ�:t�*��v<@�'w���G���7x.���Xy�C�Q3]G��o5���&Iͩ�h�Zi{.�7FA75�5�ϒ;��O �Lsq�<�
[����eD���^�+���4�y�q3r|2N`�d앢�mLWlW(cZCU%u�`�sSi��Z.V�`ؔq��:a�C��ј�
7�[B���u�����{����i��;��x�8�LL�
��E�{Y��*��Ñ h&�t���[Z3��N���k.��X�����58�4��pm�����̮Ab	�ݴ�5el��:�n��boJ:�qhZ��1�PN�T쮊�e`7�.E�Y�g
��kI�|����\�Uz�����B����7gbm1��[�/^���χ9�2)aҲwM��K�v�L��4+;d�y�<?wTTi
Zo�7+���2f1Ӈd�m+�����)�ќp��Vl*�n���r�
�)��D�n�^E�%<w0��n�vN�Bq`5�4�ߍ�=mq��u����8��ޚ��Y�^Ά��B����1������u���ij� %��p�f1Lh�U��IK0kb�^�t-VJ}�kbJ�ԩ�ݼ���![����	ŷN�X�5���i�ƬА0��]���kU���;^t��yĎ�aPe����ڬ�]a��6��U|�"�P�	9�VxoG��mht����c�����a=8d|E<}W�ݛ�p���NmSW���������[���620�Sh9�;��w��R���Oy2��hh#2��F�0�U�M^�T-�ntç�v3*�k��]ib�2V>�o,�]s[W��=mP��o+7W���t����AaJ��$�R�)	��T���1�ro,��0��L��]@Vi�Dk˵|^�p���������G��4N�)�[��:� :�k����2V���s�)�9x7-�̲�K\�N_�.[(�W�k�`Z�rpr�o^���d��+p9w��ڬV���w��WRWSz���`�lpV��«B�۵�J�	�!�����p��+�}����b��w6�j���^�pc�v�+z��I틠�j�B��ͬ7����pm����}e� �:N7Y]qu���<fWm�ј����)����vh϶����R��M.!_u��iyir���5��c��1�4�lmE�����w��K$��g*���k2nr��*7��mܲ�t�� �7c����HR��D�ق�+��}goc��D8X:�%E�i�C�0�[@��5w�6�5y��SхѮ=���nv��-�MZ�v�.e���he���˻4�8������N������C�2�I��j���϶ef\��q�ۃ�\�D��1
�p�7c��f���/��nK��J;z����y�}%���4>��ڎk�����Q��z��̫��@��Á���om�`pRn;�M�WZwݹ.���:����m���f�컑^Pn�����Lb5F�/q���˭�C�H!�5��Z.�T3;gm��T&�W(s�}�6�fQ�{�u�+ʘ��wdX�0kY��4��K[�e.����ԗ�Eʷ�xK���Ň+G�D�L���ݲFm�֊�vt��Յ-g`͹в�+�O����m�v�_؂���Uіx�ҮH�5]�n,]�޲�U�vI��ۼ�o�^�O/���Z�Ի�r�g+����v���k��B�Y:�D�M�v	�Kh(�LJjj��������ծqv\g��Ylu��÷0VF�b2���aa�&�6��R�����q��=}f������6�k !���G�}�ʕq=��	ح�:"R�W��f�ݚ�(v37�fXM���'Е��nՊ֋���x�m�֓&opg4��o�1\�E��//e�М�@[�A�Ub�cj��w�]�ۘ�D��r]��Zл�w�W@�]���'U�`,���R��6��k�L�}���7JC�;k�/o7WA�ð�2���7G+�Y�i\ܥr�7*��v,t:���bn�-6��Ǝ<�\�vw/�X�oǜ����m
�|d�Y����Ml���Io"�+��3;^rśZ��tw�>u{'=�٨�ٔ�w���t����;�f�J�V����fq�&�Y���SUl[�ѱ�L��
n�#e`�����',��fe�|�_Z��pjW(�ṇ��R�}��`;V��2ļ�8�ո�RF�+q1����l�;�NV�PЁ����%��z��;8���Z�9��Hx*܉m�ٛ�u��w_9��: ����2nV%I���4������L�&<IhN���S.�ݷ�<$���z�:��{��9�ѥB��e�5��5�_F]5r�H�,;Sz�R���2H��ԤY-ռEgM�&�N����3�d���6��ږ�bj"[
vF�0��
�qfR��b㻖������R
�L��(e������LX+���I�xIp`����qݡ���Ҁ�#��X��l�"BI+���eȋ��[��L��5�r��Xe�aΌ�V]��XmP-�(h���VC9unh�#�Ʊ���D��i�k&��P ��=+��-_n�fK}4p����w"*+h�`��pj����q'����^�`XTsL���us�i���â&�,�n�Fj�x��8]]�����;����hU��o�y�ls6�r�N�>�+�2��Wb���Rl'�vV��E�`)���rSF������2�Mz���9kۏq�E`Zo:T��iܲ4I�7���c$k"��u�N%	�F�.��d�2��X�;&R��/������6V��&_]���'�������IMe�U�|��ζ���@$�{��]*�Av;Oj�pA�h]���Qb�a���U^�� T��U���f����|�i�p���33�u����#��t(>ɴ�]����n�N�"�lc3m���d/wnb�Ԕ�"����|�-d;ˍ2��bt;�J�ɽT!�f��a��H�W���9�b`ϩ)��[�։�p�캱&SGY�
9Y�wi��S��mη"g^�����x���V
�]���\虵e}��쫜'pe�	�T�G(I�U'��:po4�c���k��zs�4��C;�{��xR{�s�Y\3vSu|F����������t��7��)_::��q�吖.���cVO�k����p[-�o$ea��;msU���uIL0O�Nj���� ��|u|�:$�%
W^Ռ��)�!+-+��W
��f��v�+����i�+k��r�vgc&�[j���9O�w>͙Ii�ZT�p
�wowr�}uK_T͢m3�hͪ�^��-D����f*�ݝ9�a��K�<W��M�ln��b�^nX�껺c�]���'k��ώB��wW��M�M=���Hf�g$�Q��n�;i�����T�!+h��i�1�}�b4�5�<lqâ��u������!F�hí��W�%�a��W�i)E�==���%f�z����ybMS��.&����hEAW����G=��/e\�R�,����nk8����P&t��m�
7������s�\wV�y���j�L�D#]����I�_*�`�.�9�D8en�0�ENS�
�����`�j���%���y!3�B�`�/r]������R�X��&s�++���9ĝ�x��9j!jޘi�t����//.�f��
8ewQ�x"D�����=��[6^��U�i�2���8�--0�]��`�	��$s�A[�{�E����́跼��cW�U�R�{U(ڥJە4�n�j��VHm��e�Ee��̀�S�YL8�����	CA1��ڊ��7��U��n��w^e�i���d�{*�1RX���5��^�K_I&G�������d�.���^t�E��V2��*Ɍ]�d=�(:�X�����Ul��]�)\���"x��٢'��[x��/V�N��uu�
��˫��l�N�d�X0P1�XU��y��zbD���ԡ��w(D�R%�����h�]/t��s�b�X����/E-WJ5�[�{�bw���W<X��V+9|����M��f�J�	�B�vhU4�j@�4����cYWk��V�B�zo$ֆ�]e����� sd_XXz��z�̺u�]����ɻdQdfo���2�YWk��Xb���fmNU��^�0HNx��ђ���g���E�!���4�����-�%ٳ��|�{`�w-�٥��!�h���,Jb�Z��Y4��ͧ���������3�.d�z�V�N�!�����@�=e�3$b�]��c����x��/�_JB� ��W��sr�V�!k��uu�֮�C#;�rlF��#���7L4��ń�cFқ���*��(�b��VǃN�����c}s�բ�E��-'�i�׭ň\ �s����zs7����++���qos�� b͋dV@��֮�2�����q��Y��*��,X�:��-6�]�j7j�]R75��IDħB�V�����:Mv�ۻ���ƛ�]���{�ͺ�2��X�QK4m��&2Ju&�wY�����o���<����y��k+�[�3����^�H�܉��i��N�۽�xr������	\#w�f�	W5�N�u��'-�{d��L�

�_gT��f	���Y�*j}�0�9qG�2�j=�S��}ί.�)R��ǯz��	���&��y8^��(�
ĕn[s��������4n�Ҙ�ޅ��ܡ��ވ�F�����۝��q��|]$5q��qJ�����v��t2v���t�]�lv>]�
�׌:kJ�4oCdTف���UΆ`DM�P��t{k���G��4�s9�p.�j�@��#��J�QG�]�ٙY��Ҍ����~�~�4'jW�o�F�8Ryu0�����ڶ�N,w$�T9��uRwS����HO~쨡��̺�7M��nXt�nkkn���"0Ĺ�v�Y<�e�KkE��$s;q�s���p���e*�v��Cu��CV2�o�_Wׂ��	!I�$�|ֆ������U-�ٸ^�5�ֱ�W,�6(S<z]�7a���G���6����tp�q��l�s<x]]���jY��a���{<cN�����ǵk�3���[*���2'���z5ЗN흒䃃KbpC���Y��\�-cc�*�W��6��Ÿ�a��Җ��&�;rQ���<l�:���=nK�n�т;]���yV�Τu��e<�&�MĻɽyF�|�+v66C;���nѡ��vĨ��7�gl�:�:����\;j�����ɢ0ZS�M�{h�-�F��y"{ks�v4%�;�u�fqr 	n3�r��n9�Hn�/���1a{<7P{E���᜼���f�,��<��*�WJ�u�q�)g(y��s�t\�Y8㔛����qn(�OT�i������Gq��9z%v����!p.2tv8xs�Y�q�d�V�C��t�.�n���]�J���}��̼����Kt������5����=k����>I�E����\�4�b����^0�vB6�����{qi�%����2���)U��k�G8���q�+Zma��Z{>�����r����pvζ4���U���&�2�:�:�̋�!�J�Krn|f����$��;N<vS���w��u�>�k��'	��uy�<�ۭ�vyN��P��!֡��Ss����a�G�c��c��ܸc���<Y2s�\V0I��e^�m��������s�N�V;A�ƹg��] %۞�n3�tn�u� �����.��ٖ�Y�u�5��q�[m��9͟{;�:��k��`�-ю����nJ�0{nwZnr�]�\��@����9�b5��)j�@Z����[X�Xκ�^ �{lz�{q��&���5nEk�wgrW\e����Ŭs��NYֻvL>�x��v��s��!lۜ6�cfd���d�4'b���wU�ZH�P�Lg��f_eN�ܦ|���ּx���y�s����8}�p�tkN�^$�qu��.O67<lViu�q�<g����6�`�ԛ>On��ۑ�n9�;wh��v�U��N���{{punrm�8=f�Gn�x�<�v�`ʧ2v�0kʽ�_;pb1��]�G����;6�v�����.�(�71\Y�d�<�q���Ԝ�,L,�r�u�m���v}���i��������t�k���G`]�[�n˹0=m�q�]�����O+�7�ؔ$�Z�^�{`���-I���qE���sZ%wo`K[�NS1u�8�����v�sph��;v[Ӑ�ǌ�"�tM�ݬ{f��,��@u�d���>6����;�y��J�[a��`�#76�^y��}���A��5Pz��{y���v�g�� 7U���K/���ly�[YN��A�n����Qiڍg)wj�©��u�94L�Y{��û(ng��m��us����N�>�ƶ��ܫۋ�9ԡ{	0oOn�s:�y�<�.Ӕ!�%�5�̭��lv.wo+�d[�[3����t�+v�Wp&+�7,1^���s���+ν��nH��yZV�d��;�l�xz-�L���%����W4�/��M�.wnp������7��	��-�=�1�F��K�� ��i6�ۗ
���6��pR-ַ=������ hK��n	6�{c3�w�{[���6��mw�v���rv�,�-%w<WKO)p���W;t�=�����٭X�2�w[���;�Dt�kq;N�܋�ݎ8�Ӎێ���u�[�k�e�e.mFG����������nz4�3Ϭ	۬yzssj�O���Epk�e��bҠf-r�l���8�K�=v�e�ܮ��ţp&u�O:V�����qpej91���ƠNK�`ܱS�S۲�[I�y��M�9�3tۍ�xe�N���W^���7��v)��Ճ��g�n�,��S�Y4�8�]��v���ַ���v�灖�`��'^�u�j�]5����y᜽����\n��뗞�
s�ϥ���N�sͪnڴ:��;����k9K.�7/a�u�(�k��^�����ڎU��'�ݞ��pn�T�����msNGG8�p�ݬ^U�)�Di�]��!;]{4n�
8�ַ
p<��b;������.&��{n���[���;"5b]��I��[�m�ݐ�k���[Y��K��^�S�k�.���c����4'�᭏�-��Ǟ=G������}mn�yz���wW��!^l��<�y�:�6;�:N}r:��=�"�rr�۝�4��Y�M��l�@�	����t�<��Z^[����i3��nmr�/�[l�Hx���!��]�'\eO6+������w�u�9w\�����Cf��o-���1�9
[r�\s�oW`��g�o`
㧷�l������<�^�����k[�������^w��6M����ϻ`�#�ݹm��*�N�ms��nNz{h���sٵ�����ǈ^�xe3�H�ބ���%��X����FEA�m����w6��@9���텮�6��N���s��kd�z��:7[��Z�j�=�	uuʜ�by��@'Y�-a�f峮]���we�ɬXH�v��]��z���UػF�Ʋtng�yX��Gus��Y�h8�������)��=n=ԃ�� �N:�p󍝸�\�F�����0��5ڷǇk&6�6��ݵg�'�-t�B.)r�[2܆K�u{��n7`�ԑ]G���.�w&vI��y�^��aݼ��Vݶ◱�VN����l���]J�խ�q��\uv�	��86\3\yՇ��1h9И���f|vY�+�6"sÞ9��x�.M*2q��Z�� �PKu���v���r�Y�m�����8;8���vv�쨼���;'�������q��8��k�X��eƷn�Ec�����:�uל	�n{;`�N-;<v��7g��^u�n|��8Ҟ'�-m֔�^6��i7��wZ�����w,3�9���G��8{w3�N7\��-u��/l[��kwmOgfw2]E+�$��5gͦQ���|/=jwO�e��⫡�;u�`�]�F:w!s�����='dV7:�d��� �cvZu�Ӝ� �Er�F:b�8N�α�WO�/m��d�X�u!�	A�wWQ��h��}�h6n�DPv�獔̰�-���r�Ōn;n��f�%���pא�쐭�k�IܕN}�'ivݸx��wg����1��,*�=��8����N�@l�&1���v�����s�YC��f�K�]Ä��v���3��m�� ��lAn:���v��fv�n=Z:T�pa.}�ݸ;j�n!�4�������W=�㚸/g�F��=N���3��|��v�p�W�����bH����9��]�D��ݴw8zZ�8�Igة��-�����]g�{P��e����csӺz�����Kk�F�nʅe�IJ��TMDQ�X���^b���^3�nܯy�<qY��W'�ְf;D�k��Þy�:�Gō�]�8m���C�d;��MnW��Օ��������F�m��EP�7'B���2X^�������m�q�ggI���s�w&�֬�[���]l�yU��9�{v�璀��%�ss�p�GTs��{<�X���0�3��qrq�9:{'.����ۮm�疉�E�9��NK/&m�X�i%ɝ	m�k^���u�˭�;mۘ��.^:�a),�G�乔�\rZ��B�ێx�rZ^B���rv�n�q=9�\���\�nȹ�yC���k�I��m�ۃz�q�nu݃1��K�컳ue�����z��f�=��A�j�֯������D�a3s�	ۛ����3�7��Y���̗[�4�F��mn��n;l6;tp�� x{���ٱ=Wm���Nƻ]��@�q�j��%�s�X��Rk.�Ӓ���3�;v����Ggl�'��"m���c;6�筚��b]۸�m���wk�!��z�[�7�g��lu����î�=r���O�*w)ѻp�4)v7�����Z�ƶ��s�ou�\�"ζ�C*�늣�v-�v΅������n�;��������i��úy�5���!�B�W����.��wN���ˎ]۶����1Զ��Y����O#�sn�BG2F�K���e6�\f��Q�G�۲��6qٶ��n֝�wn;\��/<���E�|�"���c����zDu���h�b�<⹹^�{q�n[k&��]�92v������y��Fդn{t��M�����X'],�nNQ�pY뛬n��ʡ�m5�ޜ����d���k��5�c��*s�F�ܪ ���&�0�p����rۓ���D��h݌nyhU�s��]�S�Tr�Kc��uQ���ti0�18R�8���5P@-k������e���ۃ
��5]��v���78����яp�FC�nh��͹�&�2^��ls��9�]�6�fm��U���c�'n8�y|�P�����]�m�3�:Y[c,w
�՗t]Vh�V��ḺG3�u�LG��\Җ�͗=v���j�[����^p(���nM��ܺz�\���n{R3a;�`K�p\mpAkp�dy\ud�m��8�|a�k��
�:fN
Yz�w#��ob񞶝66�^�.�8�����8�U����r���<���6`�%�g@�j:Zv�8l�;t��,pv��ڮEz�����(��e�9�dx/"���M6�u�t��0�z���>�{)N�&2v�w\���ms�.�p0k��t*n���R%@-��sQ��m[%]�<�z���C���28Ϸ���w���$n�'���L��۷=x�����ж�y�D�k�$�0s�m���=륂`�g�\,}wqǓ��r]��pq�%�]�w��ࢊJ��j�^fu��e�;f��>���sn}���y��{v�lٜY�	��8�^�wYo��qu���y�qGyݥ_8�xG�y�n�;���+�l��;J�eE�خ"H;�:���<΍:�츬��󳤯m�ue�vy��=��wy�u�����meg������;��QF���.*;���R��g�{_0��{����v׽Y^�v{{{���qw�a�-�;=m�yY�gm���O���-Fm��ZeEZvYm��γ!�{]��j�oe�;���?�}}l��I�N�>|����aW���l�㭋�`s��@���n������l8.�F�����n�Y{vaB�΅�;��<�ݝ��ݷ����}V�nM�\�<�Όh*7k��/��X��A7M�˱��|{�v,���BH�qn*M��k�^������n���v����3��nn�����+�OF�����n"�un�ͧ���X��v9�yl�۲n.���nۋ80��7;��ӻ%pY\�`�gg�]�8�=]�����u���_o]�:ێ�X��;bv�k�ӹd:�f�;u�bd���-�1٨��4�C$���k8���q�\V���6:7;���^U;q0YS�����2m�^�ɇ8r=��n;a�p �uw]l�Zw;��n'�3�cɪ�nrx��%ط+rse��ʽ�ݭ��M�j��mc�$o��h���2�g'R�j��p�����c3�㺡��	<� qu��B:|���v��H�s�|�vt]7-�z{�*ˌ`�$���;<�5b�Gd�J��5�3��f�m�ޱ���jF^�7m�^^���s����y��l��fuĹ�=� �m�)�]q�toF��(�lv�X��@�9�ѻ�F�.af����=�F�iu���2��wM�&�{\yݴO(�7�v�M��ںy�*ݮ7�}�N%����Ζ���yW�y��K�nU�ݰcgu/>��ng�[��e��\��u�c��v��{t˄�n\��u��f��=iw':z��K����C��;A��n��p^��Z�׃0m֞�j���:�۞�=P\;��x�s]ώ��md^��������F�>��ҙS��()(�WB4�-7B;hG�$���m��3f���-���N�<��J����8Ҹ��^���ݧ���[u�ØޛyG�;[ە��/�|�|i�����lb�63w/\8��du�X]ڸ�x[�M:^�W��{��m۝�]�gc�L��&;dw�8v;rs�� �;;���M���8�_gv®�������;;�p��ݻ�{M��M�Ly�z{e�n����˸��9��&Ga�=�����ŀ;n�×8�X��z�ֽ�^����m�Sle��6����;/."�6�&�
A�bm����m=�M�x�k�{裙�ޏ��M��%����֛Y��ZD�ʹ�x�Ki��ߧ�=��b���U��&���lq�P�|�g�|s�ـ�p�{wCI��I>9�,��HRh�}��K��A�����A��,���%�T���@
�+��3;W��0>���ТH�ƨ�*Ȓ���A
��ڶ�M"F�MN�}}z�	�vS�w�z��}UUt(����LB($�EX4���A��������@'�5T(O�����S�+���S�9���%x���{M�U�l�5��;��<"��3ܑ�h�!ĩ�龒�$D�� R��(I ���x�ܱ݂g!r�7oԗ@��h
2�Q"����
@��"%]��u�,�8::�:X:���.�m�7��fBK�m���Դ��J��5X�t��!�J��x�w܈�ЙD��>�;_e����[�	��\^�1x�H']��I�{&��L&z�}J�
���!`ѵLD���j��X�Y�mOlT*ud��I�mP ��,ue���DH�0dEZ�t.���O��F�|y�*��	�X��'���t�z�*�	$�&����ƊJdIJ`D��ҫlX>=�kυЇщ�审@�@|�݂A#�]
5U�57��z��&�ؙ�2�V������.90�k�'=<r�n��7�Kϖ���~_�bA �7�i^� ��s��$��Gjf��ڛ��(��MW�'qs�$�uҪ�:T���n���i�o�%T�7Ox�O��yW�A>��B�n��n�W��^�m[��AjnG.YM�ذA�օx�Y��5�%OJ��ԇ�[�2��2��g^c{�b����t�Le6��i�ˤJ4c�8&B0C�Z�9<л�yR���:d;�v5�UX�gf�]6+m��kr�}��B�	����&HL�&Gk��r��7"�p3�6ŒI׷B���M�+&��"�@$_[v,>ڝ�Pb((2"�<�R�@H��((���rF�{�>'��SB��\���WȆB0f�\di�є�mgb�cg�-��y�d�ܨ��޵95�u&*T���:�$�� �q�V��	׶�DvSB�Y��E��꾈����H��	�,5	 R�"�5z��nS��]�ѽ�-�ʻ>'��uТ	즫��헎�K�|��o1�l�-+"T� R��C$��M
!���Gume��s��Q$vSTO�w�A	"D��by��8��h�ž$�W�$����@P�'����^�s_�V6^.�5�Sڲ`����B]__�� ���d��ޱ��	��m�]L7����,T�o��\�M�l�F:%+�Djv:�%�b��4�+qРO�:�2`$��1"dv�A�yջ��s��|���Ɂ�:]B��v*���W[�/)KqW"�Kۺ�Jg��ݲ���m��s�ɫΜ��ѳ�펶��j;D�KT�=ު�e��Q�w��B�H#3�PF��b��)
�UR/m!�$���D���3jf|��A
�yb�]�)c�R3�m$�|5�׫��]n�v"o�t��%��@�;tXh����bs^�Z�6�ﳹ���͹k}�N�@P���C��Sk��"���*�N�
#{r�UCt:�Y>WR�I�׵`�ݴ��C^Ԟ�ݴZ��
Vތ"��ύՑx�S��*{�R�V��%��v�S)P�3ӝ:�{��C�9	��_��<r�<N�B�(�+&����]��,,���/p[K�
����	�-[�,ҫ���[N�-pX�@0�����3��j���vlPGF�)A��]�#�b{b2�*��F�ד�������Y9��<��gn���5�;c�%Dyz�zN�Bs��r��6;S�Q�l��q�����:�^!��[��#"��q��8§F�Z@������C����.����l����q�3��(��[k���]dy8���x���Õ��-Zݹ��=F�T<<m�aU�v�m/%���V�ۮ��q������g���;$�{�>���DL�O|���馞����}ݵ^����2���`��T��Ρa���aL)AA�au�H(։�j��ZŠ�O-ͫ��HQ
fm;˨s;�i=��Jg�I�(!GRܰ,��=�(�|z2��DMKS��H<�:��Ov�
������1(/D��iv':�_\�����Y �|���I��\B��V�l]�B�*ؚ��R&bAKcm�>'��^")ەz7v���v ��@P7�hE�7���z~k��x��5Wj��|��:wd�v�X��5�wuprl��????K����U���X�|s����H�ۡ^=��A~g�fV$�6 ��P-��r�1""D� _cB�k�-����Ky��R��9��^���P�7/���ݛn���yvd��H�����
��#�C���m��,��&�8�_ {ܕ*��<C��j�^��rV0���"���D]���P$��� l���x#�����  {��@��8�ϒ�PB�J��3}s�˴(�I9��(�Gu�wa�]ԩq����H�04"f�B}2,.k  P�}�碌u�b��T� w���F��w�_\�s�����1?7����\=+Ί�q��r�dm�B@Ɯ-R�K@"�!E&���*�Ӗ�8���ݻ����e�O��$w[wg������L�4+��r���4"&J�ɘ2��s��hh��
�8�/�>�(��@|��X�܌P7���8�ԡ����1
��"F�r`�H<�A�׾��;�gw�Ep�ˮ����{�ě�ɲT(�j��Ά��·t��4V+�u����x��Cn�F��3���.�F��-��:�U���n�>�U�J����n��֍�O^�����үA>����#�����m�$��"��W���13�L�T�	A{�krω�ZUF׹3N؞k(Q$�[x�Xmw�ޖ�eׯf��Ǐ��"F��S\�q��뜁��ض�s��[V�zc�0:��=+u;����!d��'�#~��TA9ێ�>߻(Q�U�GK�P�d��G���v�뮬���G�^�ޖ��̣��s�Nj�u�J���ud��B�F��%�l�|�mV�'��t(0fJ�0eX]�[d�s���bM0��`��ܬg��|��>'���@�LA�&
��d̃u�{(NĴ������c� ��w<���M��h{�[��<�YW�9�ld�`��f�j��	iހh
���3;�d��K��qf�!rv��v�1w
&s'br���i��=�ZAB����"*��t(�O����Ǡ�X�a��c�:>�B�$�ۮZ����3�������%,����v�G�q����:g��84�2��[r�?�_�L�Q�S%8J��9��^O��P�sN������(�� ���U����W��o�a���R����
h���A��U
�$�O�AZ!D���[۽V7а�iLD�H)2
[h`$���x�L&�z2b,�9��/��2Fwu���o痞�M�=bUan+��29]�U�����5� �uvРI#��8� �^$_vרd։��D)�f���ب
�({��Ϡ��p����R�H-cT$���vo*�\oS��W�u{������'�b�1��\�ĤV;Y�}㹒\�7�v���V��û-
���<6Q�s�V�ܷ����ލ��Q�4��n�A���kBu�c���.�Ӷ�7N[]��j(:�T�v�;m�����W=jύ$n�!�!�wF� ���z�wmnΨ*'�!���,`�����p\k�q��C���p�!����v��U�U�㣭�=�_���w�.v丛P)�ɻap���(s��p����(����6��x� y��m�.9���u9��W��33!l�쾮���rnuч*�ɻqd�E�&tcq���=j�Z��Ͽ��ދ�m�
L����֑@�kZ�'{-���\#.�	ݠ[�U-"�H<�U��LM��1J��~��bƙy��dٿm�s����w���A:��Q$�c˲A�ծ0�~������*��e݊6	��B��eY>1qe�궬E�ާ�xAu�Q�cʿ&��
"L$�*�aW�4/��H��U�H �;]�	�������d��|���鵮���"�����w�i�m��>9�6k�Y2��9�I�[^�o��߉ ��Vk�eQS@��)�����c���.x9�:G�6�)�#�t{n�c,�1���J*�V�[${�<���v9����Q�.�$�;�Y�D7+sGJ�Ё}mW� ����{�@�aJ
���i�6��i�mܓK�.l��2��u+��˺��;�@�X��'L�����,B�=N\�R�n�K&�t6�l�4�v�
c����WV�-�>'ċ��w�A>��f�>1+�s���_aP�.�}߫d�O��R���3[K=�6h�@>}�.��<��X�ܻ�ޛ4}��"T$R�&MX5{i�����pg�'�U;�� 5OcjZ�t�}^�.���{18�|�(F[\"iS�� �Y�N�D�e���ؿ}6kĒ]g*2����jfF�0Ȅ�[��4�dD:2p��r�ٻ']�NJ��f�Ҟ�{28��[;�{6��=0׉��(��	[s4�%��v	��z����]�O�>�$&�3~�I�jr�9�qՂA>��f�$��|��MBT&#$v&��G^�z���R*e�U�MH�ڣ�|#�S�Y�Gi{B!Ģ�Jj`�97g��(��V5�2��~Y�s���YƷ���d�����v������������t�o���H�.�1ƍ�Wo�[��Hl*K�XG��+JĸV��b/0�x	
�uoLM�+��o)փ��u�ΰ�;]\��<�l��N5]��Ϯ��U�z^�;�:�[),���īV5
N�.���p-k��"��{n�]��ʝ�č���A=�"�t��ŝ��j�j�R�v;�nȜ�TEn�;=�Ǡ��%��v�6D�Tc2�kn�!)���2�c�bB��k7��ZT��B�56 S�����Q�M���j���q�X��K$aP#a��cI�l����I�.K�Ԯ��}���-�\wO�i�Nw㚍���+T�D�lk��
�a����+��;�n�eR�q�\��Cs#9v��@�-��N�SMlթن7)J��lV�H땯vo^��u�*7	�O]3���>W�p�BU̩�2v��n���Ys0q�>2	P˃kf��e
�ӥ�[@�R��P�81N+�X������f��(0z�uf����w�s�����ԫ��{o7�h�I[�kN^N�n�z�=�5��5$}��t���fR�{��t��T�Av���V��3��a��VZ�#L�H:*K���S��a8�3��I�-ע�m�/2�y�ѥ����t8�sJ��Cjm^m5�P�r���K��sE�;��#J�ժ#[ً��.cۮ���!��ة�����7�ӈ2d���[n�+�u�����y�η��4�Em��GA�n�+��+�u���ggtq��w���{yw�u�[Mͻ./;:�.�ڝ�{۹���.J�:��^g3�Tu��vQ{ۼ�c���+��o^���:����眗�_N��ŖvPY֕�{���h;���������{Y���Zٷf{5y�}�q{�սj���O����[w�y�w�����e�Gw����^�/�w�\Hu��YyѶ����)(�2�Y���Rp��u�eYd�m0B��|5�H�s^i���Y�I'2�Q9����Q�RbJQ���Z��f&�x��ѢI$v_P�A����;f�>9݌�{4E�!�$J��RDɻ5�j�A���v.�����/:�V;xqT٢|H�	=�����3Ϻ��?���v|��!��4�Fs����VNC�vMف�і��J�����kd�g!K���@�Kw���ݍՂ��<�����VZ�D���H���\��PQ2����nm�^���!3���O$�}|�@�ng;�M����VB�Γ��Q����f��6���*� �zM��e��Ԣ־��#A׫�	��w`�}��Җ��#�̺��U#E休LYcu��Av�ݑ�Ӆs�X'4l�y[2�f���ǆ����۾�кUϩ�j��M�`7y�)3h��G9�ͽZ��z��]x�' "rmzbp9Sf^5D�|���Q�% P�۬�$wl��U��S<z'�X��@=�n��=�u>n+�7��]�z��$t�KD���1��T�x]�F���!$�A*h�Eh���[�wzL�*�&N���B�#/�߬O�ya�r����xO�)/P�U�BP{�P����ۥ�[���I���k]�v����'3����F���~��ZL�L�2�1~�W;�Rߵ�cm)Iv~��A;X�-���[h,�~���L
i!U@s��༅��B�`SV{���T�k~ﱏ@S��I@�L;�{x�R
ACQw�o��%0����zDzT�3&k�>u�����_����I�) ��w��H(J@�}�0RD���^g~� c{�+Z�;| �(�0ƹ��t����%�{��������@�i&3�{&D
e2RAu��22R�U�އ�[�p�H,9��>�4�C
aC
II���I2!I��S���ęJ@�o��ǝ׋�e��ش�e�47|v4-�%��ףh���4EnSĖ�pB�եH��eۡFU)�$�|�F;�e����ۄ����7Ni\��MQ��nov�s�n�q���K���9����s�x�[��������vw�Ⲷ�;��@���vTٛ.�&Χ��v'�Z�X�q��;f��u�r�m�0��h�g��muEy����㮐ع��k��������GA�mG�;�P�:N����"�q����Z;���'/BY�.6�����m�S�KlrvN������x�5�t��@�f��6�yvh��k0<Lbg�����Q�*��$�����Z�8|�B���{�0Vh�T��Z�����S(��9��b�7�l
e�����4���P�9��)��o�k�-����-����{߷�%��5��{>����˻�i�����l�%	L�������$4�{�1H9 xF�?�N����<#>N��|V#n����_%�����5�!�M$?��L���s�� )Ĕ�Z�1�5Z9���Y���laL(aI(��7��dB�)��C)���bL� T�ܯX�L���)E� "��Ϩ�t.�E�Nk��[�$*�}ﻂ�D) ����{��`)��IB2�ﹽ�e�y�1�{�nO�
����2	)���o5,���CV�al3S�o��e�$�
IHSs��3L��V��sZ��L�]�����S�k�HJ`SL
iƷ�beQ�!TT=�ox��0)�����]��u[YGnڲ���K�pŎ�2=���sL�O8��-���vm]�S��y��{��R�I(B���y���{�5�&��Je2S�{������%!BJaG}�߆>|>�
���X��]�z�{�I3�JL�FS�w�ęJ@9��L���R��m%�4?���X�����)J���~�����$�����d�]���c�=���O1�;����\��=��`����貢�� Lfr�IƵ� e%�#�@�����߳�
d���L�;�kx��4�HQ�ky�5U������iq5��F��w��,�����m��ֽ�b�"��
a�w[��i ����ן��{��zR�����ﱈ� �D*��5�CI~�U�Lĉ��bJ��C{ﮝ"s�f;E}�s�r�����^��c��Xp�{��a��0�� w��x)&��gU�5_{�{�Ad���C)���1&R�*^<��7j��mU�ՓI�;���L
�$(*��=��RA��v���^��c�0���o�� �P)��緼CI�d�(C��7��Ȓ�������.Ϟy��@	����ӹ- wkY��v��<�Ǵ)�2�[<aNh%~��������롢�ЦaO5�������)�y����J��
J@���7��2%0=}��Ֆo���7�@�Q��UC����i �����[������]�V`i4	1�c�) �#%2�o�^{�4���0hd�*$��w��a��)�F���}�ङB�)�}���}��Tg�_e�x@���Dn��l�"����u��0)����w�ः��SL
s�uU�s�X���T��7q�[��1��"�\j�W\];����ͽe@B�5�M��xiӛ�L�n�֫���޽H)��I�{z�4���P�=�cx)��>w�7@S(�I)7����u���9w��dӸq&D) ��}���4�L�
�*�q�������O����g�?u��1��j�׆5�m�"�VB([!5�Zk�5��ٮiRd)��ʌ��~�0f2RƸk�#���S
3�u��L4)�)%'��o$L�S%�Y�1�144�}���]FfsI�����	�nϬ��c웖��O���;PY�s���'�׹2���x���t�|��=2��)���{f�i-��KB�h��ofQ2��ж�B�5��9�������X�΍b�l8����׹�m�l�-�hZ%�ｼ�beas�٫�ˡ~��h�ΐ�mu�w:B���$�+�����tƀχ׽����G��ZKK�Z\���䴘L�i-�Il��^�1�i]Ы(���yL?����,O�xW׎���O��$�/���$ErTg�4���Q�����_i
fYh[,e�oy�c��-д��0���a�뚫���6�����B�\���`������i-�[�o��4�$��s����������y�aD��^�>�{�W_8���3)-
IH����&P��KB���o��s!I���i)
a�{�ƚ�>��(��v����^�2Ijb��CY;�kiˠB�̈́��D���L����#�,��{�l[�K��m^:�fy�ư�7�g/��=hZJGW��1&���.w����r�[lRcim����y�0t���)%���=��K>dzJ�{ӈ�]�Dy��I�'ѫ.Ť�e-%��Il���߱�iD�*�л*ǻ�m�ah[\ϳ�����6�wپ�^�,	���a�;�[�G3������.�]T2R{�_�U!#-�EO�.����~��ZL!I)
fA����=�C(RJB��%�l,�=��h3�̐$�\}��U�^�"�'�-&sAi)�ZKle�ﻌCI����1��Y[l���i���I��8�{�3����m%���E�|}�c�8x�G��Q2��ж�Z��1�I)
M!h[,N���6�ٱ����Z�k��������7�G���}�(��kQ���չ��6�A���jR�^�0!i,�Ie�[c��4�f�[l��������]��M�;�i0�$�e���s�����tKB�Q-�����Cn�Z�;΅�"+��_(�ƶҍ<��������w�p>C��Z�e�o��c��-д,KB�s��1�4�`���B�Yt=���i3޴mo���|Ͼ�xINFZKm����1&���Ӝ�W�U�����)2��c��1�m�Ke��в薏���y�e�W�V~�M��JB�cY�s!I���i`��l���{�m�l�-%!HZZ=���hdL�l=�ﵛ��g����`6w�^��x�YN�95�]p��+�.��%�]t�� �
E؈��������l�3��#�5z��[��E���ӽ��������r�����vo$s㑎��xŹ7!O9�w;g��K�^zs��|���|��w^j�϶�b�����˞1���k���`�9����Q ��^��K�q�f{`�rq۸L�rӺ������a^9���ۉ�w.�{����O;t����=�,s'�qZ�!["��7+�u�m��� �0� f\�ض3&il�ݜ�Z�J:v�R��9��zOh�ya�,�N��y.��gk�?_������ﾲ��~mu�;�Pt������.��{��1�c6�Ф�����»��d��L�ZKe���gI�����I�:6���1!��Zb�4�>_����\k�>#\����}��]}y���hB����L��i� A�P��V-��~�?x�8�������hX����������JB�lmIH����9����e�������z���ۿ��>!��#�B���dAW��hYDg���;����Ke��Z����X-&��$�$Ϗ��$�?�vz�>7��dغ�s�a�)5�--B�s��1�4ͲжX�Bб-��`�2&P��l���և�h�ΐ���n��c�ώ5ϫ����t���ϻ�i�ͤ��i---%��ϻ���	���Ф��mη�bC�g�����1�WI�)%!Y�gZ�1�6�ah[e���AjrTg�4���Q�����_i
IHS22з��1�C4���|g<�s���IHS����v��lmachZK���`���ZJm���}'1�U�g��=$,���D�q-|����x�9��+5�N��یEX&����\u�uϓ�{p�����ДJ>3(�${H��>�=�ٷi-��KBˢZ>��扔.�%�i)
u���P���%c=��QQ��hS>�w���le�l����ih��k��2���~�o������˼�i��з�ޱ�Ӥ-%�UV+�Fy�ǫ�!���J���V�&��JҘ�zi)W%�w��D!"{���\8ȡՈ�\��v��eN��F'4��̪h��e����,�Uv�X�KB�R��¿{�I0�KIhRJe����c�.�hU�KB�����F߄�|�HY����9(Q2M}��7��C))��घB������)޹�`�f��.%�hZZ�.��:Ϯ��MiuW|@�=>B�Yt<�5��g4��e��)ֹ�Z�c[j5�j]S�"B����m��j%�����lǱ�{�߱�$�>m%�wD�wϳ��D�eж�Z��o��4�$�)4Z���{���s\���Ƿ���fYhZ����pRL!L=��-��i��B�m�-���`4�Ie�ZK.��s��q�q��I�+�m:ҍ��o��Y���V�I0�$�dm%�Ou�c��D�*�D�.�C������l-q�k��;����~�	����NT�pGrc�7Ύz�x*@�\�WL9Zٚ��߿���W+�F��-'��{���B�R�Z�[�1�Hi-BĴ-�������A�Y�� ^BKj0��n��O��:��RL!I)��IhS�w��2�KIis|�N��U�����)4�Ka���ٱ�Ke����u��u��&����
ܢe�%�m�B۝����HRhBд�!h[,O{��6��RͲд1��xU��_w�l�>��!���4��O�μGUn��DƆ�R�Z�0t���)%�Al7��Ӷm%�2�ZX����米���G�uհ�n�x$v��fk��ٻZX��.iV]#PW:�7[\\�C�e\[Ӧ���K�;/pK�ó��u��$�~KIl����{������-
�%�vT?~�;���o�Q�f��ZRF�k�>[ic[M���`����i{/��{~�t0�Y�Zˌ�-��`�f��--IHS�}��hm��B�X��������GS�W�}�q�� AI��C)�KIig���ej�*ߥ5�I>MD��w�m�v�Ф��ˢZ<���I0�^<���x���|��ah[g{�a�)4��i`��l=���IHS62д--��Hd(��O�����_���`���ԉ��i��<������4s�fpqvL�7���u�?�����#��Q�.��-��B�{��!�)&����t���;�;f�[l���$��]�7��a2%��wg9{�7]�w��	>g�w������-
��h[s��4��R!��{�Ij�+"�L�F���i����'"B�l�-��돌����o\���3�cY�-%!HZZÜ�{�!���0�hZJG��X)&fh-%6��I���B֟6w�s��0�D��"{��uߪ�cw��y�M%��{�cl��%���ZtKG��X)&���$�)��>:����w�{9�<�'�-K-e�{��q�6��Z�hZ%��cX)�P�7�9+�JDD� a��$	<�U���s�����Ci,.��Yt��=�!��햒��ZKK+��rRL&D���l�I��9��W�&�k���Y���_"���i����xB�B�l`ؘ&��OE��y��.�B�{nK��ǕdU��v��czV�-ٲ�s���_���+�л*ϻ�m�ah[g��/JYE��Y�-�����O_�oJ�(ee�ж\e�n����2� UF3c��[@�"H|$f�����machZK�C��8)&L�ZJli-�[����4�KIi��u��kw[���֛�/.DA�]��O�(�})��գnk��dƷJ���H�*>%U½��bC�;)��I��8�;�3��Z����Z>���Y(�B�h[q��m��Ϯ�0�`	 I�NK����i��p8�s}���4�2жX�Bд��k4��5�(�Qs��28&'h!C4�����|�0t���t�|�|�������m����CI)��IibZKG��8)&)i-��Ke��k��!�5.�hRJB�gNeWu�^}�c(q��ж��t*������/��C)�-k�I��l�e�l�Z��1�HhKBб-aｬ��u�;�����q%!L;B�Yt<�3��d���)%6�ﱈi4%���|�K��|Ư��)4�0糽�L���~�����5�un�ޤ�8�KBˢZ<���Y(�B�Z���߱�e
IHRh�-�&=��Cl��]�Y�ϐ�0�Bд�~�5���cJ?�;�r�l��։����ۍ(����P���Ai.]�ǹ��N�m%��Μ���㲒a,�ZYX�=��a2%��[i-�6���1!��ZtKB�}���JB�Ƭ����4��ډ'�K��VlDQe�5��fC)ٛ�=ÉX�ޙ}��E�x���.]��
�؉L$��g�8�жx�r�,p��ބ1�>B���TIYJ^i7��Qwz5j5h��Z�U(\o���Y�t��8h{Ww]����m,��W.�<��gZ�Λ{w;kMV�J�A.��ώF va��8�2�w��&#�n�r��]�f�K����ve�_;��d�oZ�)�#5�����·��.�ȳX^�U���P�Q��9r]�$#�b�dΛyר˺�eAU���I�)���s�����]�+���H���^li�s�N�e��i>�t�źE� ��2��u���V�X���{mR�i�����8���(��A�y���=r�P�%9�oi��җ*��a�����*�������,���"]�<&K��q\�t����DZ��Y!]1T�X�Tחl�ԟJ���l�媎*�ɵ��%�F���n�9�����0fh�Cd��v�@-iQ-��|��j���km�	׏o$�}"B�����C=x��-�vT}Ӵ��d�R�uD��a�� J��k� ^K*�zI���K.�[�V,G-��V�XZi�n����ܭ)v�^�y��2i�{����/i��_Txx�ʶ��¾Ιh��+����T7�Qa�EEl�.�[I;X�_d�������b���z��$�����n�M�Q�!���T���2���f*�ԭsؤ��K_�ǔ�nPrt݋yv�qM�BWa«��&Նؗ�OcFZ_�n��������^v��RE'k�K,�f��eo{���=�,����{{����w�٘�۳#"L�ȑ�زˠ���Qm�uy=�KӼ��Ym�����V�	);����.��v`q��y�{ݜ�(��99[F���I�m݄gaBYd{nL�{>vM�xIK8�f�����vV�D��m��\''fqY�ՕaHQ9��i�n�	 ;"�:�$��JC���qm�٤ڷ#�'L�;'��.�0�hNzj�Y�v��6�eklr��@���I��޴yͥ�Y�9���Q$�8͕������"i9sK�ӤH���E	G�[��=�nkgn�sk
I���4�%fCkmcl��ߏѽ�sZ�������7�^��[a�HT���H#s�m���&�v��홳����U��rb-��U�]�l���X�Y�R�f�y�Q;v`�P�u��nM�g������vq�t���ܶ,5�[�=ts���e�b�0c�Wx�w=��û+�m��i^����F���n��7����R�z׷\�����MĽ�����`�����9c\\whQ�`��:Fܝ��=st��u��:�sۮ!�wd���[��E��l�9�i��{k�a�ƶ�s�f����q[\��6D)��u��2��"r�6����1�sІ��3^���|tn 3��X3�����qq�9�ãs��nq�������5מ}�]�f��;u���������ג�*72u�m��j�,�C�Ј�[��v�}v�y�&��@W��-�u���N8��s��t��z�
ksjZ.�I��<�I.�r����m��6Pn���M��m��Wgy�S�Nλy��&wZ浺��2V�/)����۸,���^�ۛ�����5V�˓i�9�9��!����f�.z�n9�.-�=���������=�������*�wc���Cجpn�6m9Qִ�=����Ϟ��l[�U�H��'�؃��6-��uyʘ"ѭ��F�:��n9�a`�w0��n+����:��n�oZ�8;oS٨�uY�==H�=��S�q6�8�����P۷c�|糸���=D�{;��WMu�M]��-��vѵ������j��[tU��G;K=Rq�Nq�ˬ�m�m�v�\iC#��Uv1���c,��$�hrʎó�Sۘ;�f#p{N֝�o��۳(��i1�ccq\�=Y�==ԛ�^`���&x�tq�jq��.�;-�v� �\�;vm����=qɓ.CX�\��kv4��Rś^�{g.�v��㱶yt������v�G�6B}8iS��!g�kvW��#�7v�͙������u�i$��y�,�%�vo����o��;ƣ�k,�Јg3��l�gu����g�+�D�׶���j�O=i]����Xʮ����܈gFdY$���v�.!�c��PB=G�����4��dN��#n;)vα<��u��qb��'��σ��Y��;Ke�^��gN�s;��[=7Wv-�Z���{a-`��ڢ�ɥ��UL�e�Ly��m��υǜl��;b;xZ���Z�xI�9J�p�۵���I�5�x�ex�u��b�˻q*}}�~���������i��B�Ǳ����h[-����;�f��,KBд�-��|����$�W�o��@�=ߴ�$�w���I6����2�[c�={�־[i|5+��DlN;����'ɸ���;��c���Ih;����|�|���>���]�L�vQ-lah[x�=��HRhBд���l����m�l�-�2д.��[�����t�?o��HxL�l/]˻�v�/�]]gH[h[����i����Yt��y�;���$��KIi�uC��W�61�#�CI��2G��q�������h�Zr��{���\|(Ҍ���m���M|�K�B�������fw�����g̴-%!O���L����,ж1����a�mapmIat>�5��s.�n���y[���%!I)�-�=�bM	i-9�`m�1��h��L�L>絼i�v��m��,�%��}��G��=�����WB��=�2|$�&^n��HRj!hZX��l�7����f�hZJB���}�k!��Ø�W���G�Ɯ{��@�������.^ΨGE\�Ů���g�.<m�sh&����}��OM-_�%_T:���<�q��-%!I,�a���Ɛ�Jv�Iiii-.��k%$�f%��s+�7^����T�f����!�5.�hRJB�������q�����5���Ȣ,�r��m��m!h���
L��-��-�������}��:�D��{�����P�m���Y�ۛ
Z�gPz�*;k5f�G/ҩ{r�&�I�Xl&oz_YvϽ�?��|�>C����`��!hZZ��h[�{��a�ж6����{�I3�IM�ZKn�����i�{�bV�Q��Q]>��~���խ�[g~�6ͻIl��ZtKG��X)&��-IHS���}���w�w�ǡ�)6��ib��ӹ�y���le�l�Z��h���
C12����/&)[D(f�Q���(��~֒���w}�wՊ���{� �=>{ΰ�3i-�2�Z\�Z<���I0��Z���籈e��f��}X�vM�I)
�C{�;���cB�/Z�h��ie%ES>Q����J4�o^�Ɩ0�[-e�з�1�C4���py�g���0�D�-�;�wCL6���д�];�`�����)% �o�^Fx�#�F�>3�5��5�Ƶ�6��@Ddm���T�n�r'�����ZM��Χ��޹���ϯ�����67~�w���l1���6;Il�������~�
�D�eд��7�s��4�&��-9�p�g'�a�)����4��і���)KG�wX-�ea|�������2���0�`Hs�UN���t��3�;����xa���cOFm%��Iiq-%��ﻬ��	�-%��i-�ۍs��4��薅]H�}e�����կ���v����>Q�Z���l�(�jaf|��ƶ�Q}�ഘB�R̲зﱃC4��ihZ���@5���u\Ϲ�,SYA�]�`�R����7׶���2�u�
Ot�6Nj��=�~d_�V��������S%h <�w����Ϸ��j��u����;��Cl?Fж6���{~�I��ZJm���e��?}&�I-/�=�V;[~�U�d�O��I���z��e�z�Ǹ�!̏Y�#҅����8-&��KB�Z�=��CI�B��-e��y�chm�}��kxs~�u�;>d��@�W�����J`Vw�U��wuJ�)���|r������7��.�9�9磌O�׹i8�KIiu��̖�RJfF�[-���>���JB�KB����� 2�|$�'W��w�}�"LD#2%x��|���t�5Ż]{H-$U�
�v�>���#������d��~�F���i�gt�_�ice��-��B�g|��4��R���l=�s��a��-�Lk��ù=u���w�y%ˡ���I��ZJle�����<���j	����{+u}>g���Td�&�B[s[�6��i-�6�����3��̼���{~��D�r�h[l-o�߱!���&����y�cHi�e�i)
B��7��m�ld}�$QO���6ʕ( `��_eCL46�����i�IHRK���y�i�f�Z���ZKO��{���ؽ��}����kŤ�hKIl����m�{ϡ�55D�*薅�C��=�����(��~v�"���k�,k0��}��q��=_r�=��Cl�-IHS�{_��BĴ-KB�^���;Cl66���д�����i:)�ܣ���*�NĻb��OƉ�U3S�}�Y�˘h��cVڼj*��P��c^R��3��G����Nѧ�ֳ�ā$3��J���2���5����j5�j+��H�]
b�O��{�y�3��[,m%�atKG��x/4L�yη�v�U�-�0�ah[s�׳�i
IHRiB�i��}���7h[-���ih��o��2�����}е}�{V~o(4�y;����[<���+�oq�=���-�R����W����"`�h���iW���iG�{���ސ���$��-�9��wm%�i---%�׾��ZL&A-%�]�o���w5�u%3@۟{��4���-
�D��
��Մ/��HfS�P�IJ��~/0�4��}����(ee�YO�5L��k&6��� #�wU�d �KB�R�����a��-��д�]���ZL�����$��c��ϱ츬��e����CI�-%����K�Џ�%1�#�F'�o�ϙdzO�6�л�Z<���Y�e��Z�ah[��s����5����ކ��؅�i`��l�1����f�Z���,KG���RL�l,��o�V}�V����0�`2@�����>=BS;+}Ci)
I��-��sv�KB�R������RL&R�Z��cn7�c����s�0WN��:�fQ-��y�~�\k�>g.�-�O�-L$�i����{�I���X�B�A>��`�@�O�E�R6�a�-a��]Ɛ���l,B�]���7��g��i-�[����4F$zHݕ��q��Ԭ�3��2�\þx�-:f��E�Fg,Z	Ɉ���s`_t�g�[V:� �����+\�3;r���K�4�{?�}�_/���� 
K/`z��A�ۇ����X�-��`��vu��c	���֣�%������^�&�q�����0n\q�v��Hk�Tm�w\n3'k�.,mY�h�8zٕ��-��K��g�8MkV�A���^:;�:8x���ғ�l	lno\���g�� j�q^/O1��u��������6,���s�pt�n�ܚֵfv��W*�u<saW�Ի@����m��x�M�ղp������{ה�v���_>2���%��}��l۴��IhX]��߷��D�eж�Z�c|�s!I)
Nk�ʞ�h>Cl���m�l�-�2д���}��D���y������)��:C���n��c�t����$�_gA��j`R�Μ��k_Շ��)%%Ĵ��;}��RO��������m���bCWD�)%!W�9�Qc:XX�-���n����|$�&E߳�����J�S>Q����iF�״Rf!�-�h[,e�n;�c��Q�����H.IN�����Խ�K��h[д�]�cx)'�RJr�Im��o��!�Ж��|���|�DJQ�#�Fx�>��L���W�W?Ht�,�6�Ф�������+4KB�Z�;�g0��������5�cHi����O�︯]�i$�) �̹�4�֚Q������;Q)kS�i��B�{z�C�-%!I.�$�}��a`���&��d������#�G�����9��|�KIl����8�9�C(RJB�D�.��7�m�F�gy��%�3]l�e*��
<nR6	��9�@�;���5X�X�#��e���+D׷���Y�R��'X��kk�C_V�3 �B�l�-���`�4��bZ���l/��������0�1��|�;��=�>I��5�s$�1Ai)����n5�����S�=�j����R�ɤ�&�[s��6��R���rf�;�¹�%�`�&(�4�1`�WGO�q�,ܣ�j�j:�֗^~�-���tQ1�N�M�lLqj+��<��ܵ����^킉����;�Z��G�$ ������_��B�h[cB�~�q�e
M���)�'�s��6͌�-%!H}Gw�j��g���^h?s�C_V��X���1H�2J�C:C�mw�{���t���[k��4�Im�������|�J����}�����'�[.��)ǹ�bCAtKB�(���T;�o��v?�iG>��=,-r�m�g�4���V��c�)<U�z�c5�_He�h[-����=��-�hZж�{}�����l,mIwG���
I��^�)u����e���[�k��4��i-/����o�o戴�$���g�ƙ��Ke�i-.�i����Y�L!e��Mk>���/7�i;ah[f}��0������3Q;����f�h[,e�i)=^��)��-��g�z��y=5��ԉɪI~��D���	�<>�kj�2Eny��Ԯ�����?BU���~��z6������!i,�IwAl;��Ӹͤ��ZKB�Rz��0RO�1-%�5�׾����M3cnw����%�VQ-��9��Cn��F�{�/�d
�R��&�X�Ʒ�J1ϱ����e�l�u]qyJ��M�C��c��Bб-B�-af���;Cl6��������0RL��Sc-%�(��_��Y�1&Ĵ����5�5�o�J�&�|��{��q�m�Ke���.薏��0VJ&P�(���0�-���}�k��ν]��K[#i�ұ8��A���kg��R�k�'a������7b�.�g�^<��^� �s;�d���)��b5<�p�� {�����B��!hZZ���y�cHi���-�2д,KG����SXҏ�=�ٕ��9%Q�ʹ��m8���}��3�sx�̵~���4�렴�t��7�;����Ii`������2RL&bZKe���m��=�CH;���o���V���AIdG���� 2�|$�&~���L$e �B`��JM!i��;��|�3#-e�г���a�$��gMX��;*ބ@d%�l/}�=���mIHRJOW��#��&$D��U����߾ǳλ�]��!�7n�����ۃO]��\-�O%��+�N���rZ�gWT��7-y�]g��� A���� 9����QرN�rk���:��Ȉ��u3J g3LQ0YWX3)�zG��I/�Z����fP��k���n�?Q$��ctH4IV&�$x�u��dܲq�krZ�ǡ�Y$�c�b�Y�yޡ[k��\כ� �K�7���9��	[�̱eqѴG�s���e������$aY?h�\�&j�?zl��ݣi�\��(���K�ϻ��a��fg�m�wW�/DW�չ��X��|^�T�ib�K�d��('�����SS��D����N˕9w'O燇������/���kf���8J�bɈ5�߮` o��~ͭ�����C�VY��Nz$��=��	'�樂H>�VW����?3���1�ҰD��*��c�v��m�C�4�z[.��]W
4��������]5�\���gM@@u�\�@�������;7[��>>̶UY�&)��&o�]پ�(�c{='Вjxz�J/�Z���I$�{�I'��W{��铤��C����(��v�����0l���� BGq��J {۪M��]���|o^���w�����W{��@�9�6�.ϥ����N�2"@oۙ�����w{� z��3����w��>9�r����&"IF���5�f>�A��MQXf�sY�R�z��	���f���j�������֭�v��܎wiFշ?.=@�D��#��L��
".�(N��J�*F��ٻiJ����n��!2^�٧f��< ����� ���F�E`}+>�N0<�1��`8u�;��1g�*�CG^k<i�u�{sV8��֮���4M	4*�N�oI���tx�4��I�t����l�,�n{-i���͸��;Xt�����Y4G�n0��/By}�v��;��b�nSss�Ŷ�*I+��q�{����<^uۄ��r��3���Ս�ٮ���{wH���ٳ��R��ܜ��qэ�s�R2.��p�C���׮��S�����6H܊�֏�A���>� 9��{ zOd�m��k///6y��yэ�$Oձ�H�x�d*�������o�G�=���{W9��̒@����>��v�W�	����{,���5$�M���w3��7�����5C�I���|';˽3`~�Mzl���I��>���~����Kbv����������b�a&������O]��_��}��G ɰS��4��nI	*O+�d�'0��t]����$�1w��2}��@�OG	?_I�J$�I��>�`"O�V�.��y�ҷ�`��L���J$�ڄA0���A��6�ܦ��:��K��G:?�\}v��Y%������l>���T	$�վL:'��VFqw�ٯc�  Dr����+bd%)��[ﮝ���Rh�.����pvL�Y��j"f�w�o�.7Y�es6Ti����s`�bͩ6�D���GG6��b�`��5�k�n􌙼4� ������` /�{�h>9�~����Ms�]�=�/��x�k�ҫ-����?�9�TH��OĒ{;��uX	�ee��� �����`|��$�M���.2�Ź��"��wV�3�s� h��Ud�I$����=�= >>W�iyބ@�55�3|{Z��X��ՠ9���D�}�9ʇX��q[}�O)����+7y$ �똁� �9�fm��y�)5G�[�F�	��YW�#w���^eh�c��vx<7Z�vݗU�T�����J2���L׾2znk��o\��� �۳� )72���)�//mY�Do[���Z��ވZ��dϏw������Nr�=�3Jww��dɐ A�y�7L{�癀DG�D:�l §;&wxi[F�YO�σ[�` �=��� �|�&��T�u5=|���Y��3Uc��!VU(3���\c�]�.EA���1p؝A޳#R��3�D�L��(��.gq��� ���劇L�wZ�N����M�)ZD&f��{��g�v�B;z�]��ѕS]����z�|����b��T���Y��b�3�ԣL)ٷzb���K-�jv�mer��4�������VA³0�Fe��E�����^eu^mP<wi^�n�j�\Js�Ԉ�面�wk�ks:�M�m�f���n;�huk�t�mN�ERY�k�r������i��{k-v<��h�wxJ�����f�jD���`���z�T����̭�X������nN��\��;L�x����Yj��.[z.���uk0���R�mf�!��d`�{tz���|5��lL_Vnk�1}���"�TF��ŭ��̈�zd@.��=���C#s�D�*��t�y��ve�N�x�x4���cY����F=�G��)� wK���ξᔍ��ηm�B�ӚT�����a[(��h,[�%�{�ҡrn�E�|JWn.ǫh�P�,�hq��vЦ��
R�ve��S]�J7�P\o	[�#��Z�w8��ўW��ope��O�ɝ���1�-�Huӑ�6��`h'�P�P��X�6�����b�i���ptE����3�T����݋�Y����O��������6z����֪-�wy�,�f�n���յ0�<i�ٹn�7�F;ۚ��
���S-�v���|3�/�V���3J�eZaUT"�A�5����趵��09f[h{sl3;[-! ;��,��jmh$���$v�vjz�{d'�pf�8!�'=��q;�l����H�
Q��\t������<���IJ�㥙A���"6�2N4(�Lǭ��!�d�l�8盞��l���n�;�����Z�n��W�{y�f�!zݨ��x�&�`輰p^���VLjG��"q�^��	�'���)�� �t���Ӽ׵��v�v��+��	Δr8tIٓ۲ٵ�hP%�a8�I����t��ݣ�μ��Q��q'N�Nqͻ[f�-�ެW�G5���tD-�vݩ�{o#�ȭ�mck�B
E�N�s��Ď@���hr�:��Cn���W�kRp,��[9)�6Ÿ�nOn��W�������$��A�� ����@	$�/y��R����3T�U���37�t���Ke-�)���Y�5�7�+�$�<�qI$��{dQ$��z@^������=|�1��>�q�$�w�iȧ[M�*ʳ5�����|��+��۲�/���9[�s�">�q	�������e�Ue�d5�b�����-�6��>��K��Η6��X�p�c�81�u�;l�=��ҍ9Uڸ��5t���s�����K�6��N���.�˘@{��w���ߍ+\�k
�L��}VI;W�M��.e��}�u��7	?~>��Y X���f�]��^p-O�,T�k�T�������lH=�m�A�9�3��/v�,�{� ������ �v����=)TD�Vܿ�d���/vS�wx��?��9�Bh�O�w	D�5o�_�⮀��g���Of]�kg$��M�W����X�D�}��*Ӯ�F>���7���&��vҌ��o��+@)��'+@�界��G�xy�'�]��3GB��R
$V`'
�/J���I<��f��|*���� ��s��� #޳`ހ9�z� �ڼ��k)�y br8�����6���\���-����n��Q�S��~��^A6��*ߑ39��l;&�� &�o���^����]�����BMOz͚��q�aF��D*�Y�w��x��!qfz{3:�6|���a� ��=s��)��?]g������J��5�#=f�( ��\��o^��()^��7�����I$�{.�Y����>�j�YdL���vt�yW��� ����VI&�5����'�=%��W��{Ӊ5G�\�V�cҖ6H�m��05�z� 7�s~��z�އ�4�G�$��m�TH��n7D�D��������=�7w������!u�t�ժV�Ɛ���5��=���ah�0�d�ͩ[�L˭�u�N�ZaY0��3o����r��9_{� x�� �Pq��"e	#���">���7��Ť�:����Rn��@�}������y6��:���b�.�ם����-��vM�],g'Y����l�/O`�X�7+,n��-�k��x#\Cu[���;c�v6�Ivy�;��\u���$��Ƭ�:����^�j�0����[�՗�ܝcE�g7�\�\Z��;l�r���#ٷ6f�6x�Z�Y�v���]�x��z�p#�x^	敎9��N��Xr�oϯ���-j*6�����Ud�h�)�� �'۳�J$k�c��j�s������7�G��\�ۜ�@�[M�*ʳ	�緽�������W��R^{����@|�Y�wX���g����K��E�@q����{�Px�d�B�՘���X �s���	$*�ܷ�;52�	�$���� �>�sٛA��X�aH�n��k��+ϥ�+`��;-G77��OG1�I4L׾�� ��wG�7�A�}��jz�w��eR4\�{��w�� ���M%I�s�Ä���L:$���B@'�v�z��w���y�)#n=9
�q�������t5��Ȇ���n���^M�\��������8�l�����\X6 �9�f��_zOrF�����_�����>|����;����{�etv�eaMb=���(����j_yp�[Q.G���1r���Z9֯e�(���,��uەHN�8�Ǝ�Yfa%�bM�aUY�7���6�sk���~I%�������� %�{�����G�{&��
�5���6�_)�>'�z�5|G>Ô�|�%B d�H Z}6k�u����/_������ ~nG���m�MI`�]�0;��>;7�P�����k0l@|�ߝ����&�]i��S*�� ��=������e ��:�5���{sT��؇����t�߶��=�I�h���ڬ �7_�:�qh�E�my{�����bȻ��T�V�\�:�S��n�j��kg��F$�\(5(�q8X<�}�=�r�TQ�Q�{�f? ���MP �g���\��=M7�����HI�ڬ'���*0n![,�&��\X;�;��v�]�l��	�I'��۵� ��L�IZAyʼw�I�{}�����Qm�����g>����9t� �9�,��zCc�w��*��a��`���M���V�
�w	;��|�e����fو���p4���K���-�с�oSB����q=�fS��m����ﾩ����I$�?rk�1 >9��s��Rti�*��'Tm>���w�c�y�7�M�=k@wy�c�{�緺���v��)�7jk�9����,��f �m��ݻ�T2�Х��l3f�&���H�s�7� �I���HK3�g'��Z�g:�	���e�0U��n�vEBT��������<ؓ���v~���[8�J��;�#!��PH�~��X ػ�s���i�ZE��D����������J�P��q�m�(ˑ���3�l��a;d�_�Vw�& پ�ڞ%�ۀo�����*w��I�D�j�ϲ�k��� s��l�m+��bN���v� ��Ll�I>پ� �/^�WT��+�3C;7���%-��Q {�� ?�5�7�O�?O��:�'�m���4T(�TwAB� �9�Z���|�k�u�M����v���۾�}8�N�t4���;r������ئ����k��;#� <�|I�F-�l����}b����r�6�~�� �:Om�
��*j[�eF�3��â@ݜ�f���;ɥE-����a��zc�t�/�\I�2u�ݓ��&7goHE��lKvfwvg�P������~�~jK*�\��n����w���� ?I�H����:���f%7��^��I=龒��^#.�f���e��k	��j=�^;��icd3���w{�� �w�IQ���[��:�k��{�֔�\�5-��ra�[�B~$��{ma?|I%�����ދ��{ ����{ z�ҡ��&�j#�;E�]�k����晻{�߃Z�rv��Q&�4^�c;�unc��ʶz��M�I$��U��W�"�0]೅�������I��̩���P�����������{ CܚJ�@#9���1��y�6]�'�LP�v�n��G����{���f��k"���k�QSٕ�xO*[v��"k��*cA"v�{w�[顴�ٝ����x�vUP��#{\9+�I�珁�&�3ێ�Gm�m���R��r��vС�{P<f�؜��;�Ǎ<����W�_��vyP��Y�F��ț����n-�m�l/eݠ'P��q՞��.�K�!ݮ')���b���Ÿ6��sь�%1���Sz���<2�T�v.N-�w68ϡ��qp�Ѹ��]�n` �wO��n��ժ���tj-[��s�u�;�nL/>'I�fs)�7[sq!Nv�O!�a-G�~���mX�uw���w����p=ɪ�g�� {�����~O�$�I����ڪ�w�`7��]�0;�ˋ�Ʒ���剭�[��3>�I�I� 	�z�oo��{կ�;�?5<#.�#+���=��� }�\K ���7��k��c}@��ң =����j�����Ԃ^�V�;i����x��Y$��S��$�/��  ����ξ��b��<C��2ɥC��MZ�g�ŗ^�n,��9��Zc��-fKs`/I�A$����n�$�H�>u%f#x<�7���Lo���2��v ݷ�}�0u0�[\�
�,��;���,�Gep�x�3�= ��\���^����1�^{��i��9�_Q���\π7���L��%0����i�i5w��*!�s.�m��}�y[x���ȡ �\���NDL��]�N�襵���5i��z� �ظ�.���3
1�f�=� <.�#}����y��� ��o�f muF��[佚�t���s�ء���q8�Y��ǎ� t��d�I�v-��$�ǜ�{Ӆ��d� syۘ���o٘�]��aH�����ό���~�f��v�!jєI�_���$�$��m� z�*�������ww1���;er�%ˇ;�f`�y�٪I�ξ�.�7�ja�&�5��m�'�I�Ua�6�s9y�t�ݐ�o��ȫi�Z��'&����;��v�o+�nA�l�w� \��\��ծ6}QlZ�����|���� �&�,��I�D���o|ߵ�@.NXە�ep�?3\8�$j���N���׫ ���� ��WՄ�����i�xǽ'�	�&�w�\Uk>&����m�٪ Z�5{�M:�v�7���?�S���q!Rß�q�:�f�[�ې2o`�`�#����Wr��2U�	��]+��*�;� I��g��UJ����5J��hҦ�͊���զ���י�՛��><@��X��Nl��{��tq\���l�9�{z6ݚUg֪*��b1����A��,7��Gͫ���<�$G���Gk�'�*�r�K�s��Ni�*��hN��i+��m��:{X�y����n��9��L��]��9�����{�9l��ԗ��}�f� ��#oA>���'x#{y�w��w��ͦۢM��;�J�����j�&}U�,��k��:d�/ݔ����*����$�I�7�ڪ$�j�k�0 ��H=����֡:p���Vѻ+�4��p�m�yˋ  �����{S}��q�l��b �3�1�<I~���a3�����{޴�������	 ���� =�佡P����X�l��tD�Y�}��S_�����k�,g7�:+���SV5���쪿m�b�T�EU���}{�w\�B���|ߵV�{��X2X�P)^`~��������Zs^���P����|g6O 3[�� >�����:��Ok;���:�Ϝ|\��v�Nu�G��ݞ�u�/5q�*�_�_��E���UY��{f�>띺m���6���H߅z�@��$�^�l����e�;r\�ӻ�>�A�G!�vb�q�4�b�L2I&����'
x��p�RZq�3r��%m�Cw|��X 9��,� ��g=��d� |f�˘H���f|��᥍����+�3�3���쳸s�/r�� �;��� H�ٺBC�����	$�>��4f�7u�e�R`���M��6"	��J:�l�e�k�{��k�ݚ��fq������3HoӲo!צ��s�%K�e���%,U�x]ة%�awo���^P����F�Y>B�ih��b\Wcy����=v����
�E��L�8���D�9X�.N㜾헤�;���mJ���"u���6�Я
�wR��,�/tnv]CSB�"S��07�cj�/a9Ih�./f��5Zwwhclc��ږ8��zzoٮeD��MT���s](_e����8��ˍa �lv	`��s��UT�����i�<NUPN��Z�V�Zї��d&ѻo-��U�q�m\��4�v�1Ov���ЋO�ZXJ7�D	��^ң�̖��-y�H9�u).�u�퀛˨�zؑ��(L�7(��v�.g4%a����78/z����OW$5�䫮��x�u/�C;˝�֣0�����:��w���&T��l��W�Mml�Y�
kx��� ���.w��[��f;�Fwf��L\x�O��t��
YP��5�vraQ/9@�ROvg:��EL�s{��Z	³��wi���\�*�5e�Ɏ�G��
��iXٜss��H�T�7hZ�����P�jl�y3\�J�������[Y(t�����mu_E}�l���KK�rR�Xf��f�/�s�i��!�v�۳�=�z�xX^�<�BnX�mrB��3������w���;WyS%���9ob1
6Anp ����6L��"��� ��8];Y��Y۳D��Ѭ�g2d��Y]����p�3NiWQ1	�«t1uHsGB�r�[+���yp�dԴ��*��Lx�|I&��f�;�"8pv�6�j��թ�n�[Y��Pm��IK{�� .��<������#�;n�t'���	����"HAe�1�Ch٧96���fY�����́. ��{Z8�:OM���I%�㐝yM�kq/{�r��D���k%�N$[[����)�8�;;fvZN��s-,��1���kD%����8��;mAmd�Є)qv9Om ��̠�=�+l�i.pK��3����Hr^Zv�V���Rm���^qv!�;m��%XE6�"���E�չ��V�<�Om'�d�NN���ȒR�r=,�Mmd��ǘ���!�戽��(�R��'��J F݋��Tt��	M�n�Ĥ�"\8e��:�pa�h�MU����J5���Uc��U\+v���+�8�g"�{-+�v/N{=&.3���ֶu�.؋��]��w8�0�h.-�:_��]WL�r3c��	�0�֢8��3ΌC����yy�c����gp�m�ջn���v���:��.���|W��ܯL��{;v6���1�I��mك������{�N�{nL]�f�E)��J<;n6��^��s��g��!���d#�+Pǭ�O�z�l�p��,gm�m�!�Npӗ����i6= �cn�	^<�&�����a�`�\�7c��g�]�2U�Z� h]B�mؓ<��5J
\��cI�y]q���5	�k��������8{���An��wZ����uSn*c�����+)={o��Gc�7���9�;"u�ό� �gj�vw9n��*�^����_n6��ݞ���͵��$E��t�xz}���us�ۤ��:|N�D����\�y{m���t� ��OL]�ȓK8�lu�mӻ7�n�9㷷9ݞ�ɫDq�';������z�ތ8�SΝ˜�h��ɫ�7SکK��D�v���R)%X��.�Gc�m4��u�S����m��x�q�Wn�,��d]-��G6�LZ������\���6K��h�ܦv�����f0cq��Ӄ����W�a�ǜ�i}�磬�g�A��d�.e�<G�z�y۵�tǏ�[���h鵶�-*Bc��Ja�y�5ܮ�t�z��Iŏi�c�������Wb��y.�qj5�2\�r�N��u���uk�:��ulc"��z]��2vBrQ���v�hN]m�v�h�-����m/nנ���֎x�BOm��ܞ����Y|b��ɶݷr��tW����n,�൹�zr�nr�!��m��n�=��� �N[Gg�랽���&����&��N9we�(�le*�g�KUhl�J))�*�an���e���k�J�p\���v8v6�fz^�Ì;�[ձ�݈CxY*Ͱl���'������ӷ`딗q
V�9x��ˮ�ö�:�D���ww��j�ͷgѝ�9x�l�f��ݫ���xLuە��C���5s��ힵ�d��8�u�����sz�왎�r�plV7Y����T��uة��������ju�ְלM�G��ճ�t��[:�f75�h5��-�Bsە���{��<&[���LN��s��fM��4D���#nW»O
q��G����p�T�U�[�<vN����Z��:M���yx��e_u��R�9��Y�M@q���s����������L����9��ŀ���f ��m�mVw�}~9)�~�#����g��gu����rRJ ��5�9�T2��1�侹� ��fg� <�vj��^m�{��f�q��4E�9)��.\�� y�٪6�P�&��d��r�D����'��;�T���n��ƭv�A���H����$�>��� ��D��'�}������puj��m�'��S E*�حt����J�=����h��s�=b���\�33��ٯ�ā�\�� ]��2���Fo���)���=�֌nN��e@�;q'���c�$u��c�jjYn�����UT
�߾&s�� L�_a$�OܷɆI���sK-�����0 >6�vk�o�{p�d�9S��X���\�A�Xc���˞]sӶ�"sMBJ�aY�����|5o^��)\d�.�Vi�(纬h�lsb��`�)�P�"�Y�(UX�H��ꪯ���ܿ}�t��oG���3�g�z7���.s�ټI�t��A�xh���X����bA�w�Op�6��W%��9�>�wf�����`Zh�lrX��T�;i����U�"u��Ո�p��h�I��j`D�_�5�ϮTF��H��j�ؚ�vش7s�����3���:������&�@")�� �}�́�{)g�5�i��{�B��x� ��P�b,���:���ËVq�
�ӎ�������8Ij7���M��ڭt��3�Ua5D��72I���N�q���n�����߮�|�$]�(�p*�19�ϰ����l֟}�\��7�� �ܺxw���@ߔ�1�j��t��{qCr�(܎��w���`{��g����3�/j��W^`K1�^i-p����ۤ�e�*�dio����;����j6f�={q�P%��$Ƚ�T䋜�ɧs�{����� =�v�|�s?fb{�G4�+����f���έ���r�����;��2h���Ϳ�$����>z�]�>���Ā���ۘ�Rl%�jK��w�[d�'�|CaZ���$�? �{��<@|�K}�s0�G������{�z���
�q��!G�[�:��F�{8��V'�M���ȤRB���7��WDԣ��ѹ�v��潭<@ �ݓD�n��=1�&j��'w
c�c�7j��1s8G�����窿N띸���׳o<�vF�����4m����7�}�$]�(�nU�H��$�D�|ͅ�$��z�fZ o�}�o{�� l���_S��&ꥭ�5���{��_l��'4m� �4I��mQ'�G��\�{쥓Y1&-���[��tu������R)^0��k�U�s�od��{Y�u��zZ�����7g���[{&1��
,Ԝ�����I?������%rQ:����T7������XR`/%��4ea�'��՜X�E��gk^Gb�JD�A�`�"S6M�^gtǅ�շM���\�iq��=r��A'�~���R��]_$o��b� ���*�	�$�'޾��?9��G����^15�k��m�H�٪���j
��I-ǻ�(��k�ڴ��^=�kO����͓H}�f��A�rk���ؽZ�gu� ��k��Tn�k�a�3�z�ɼY �K���|�]w�� 9͑�|G}ټ��|�$]�F�nU��5�e|���{��y�ᤨ ˽�����fS��o��x���{F���=�������tl��q� s��6F��E�V�D�f�Q$�޸�Y�]�ͲW�̚���iW;Ρ�S�	�ͽ1�V�M���ۋ�v�;����puYH���L{S�[/n�xm���a�%���Z�������oמV�Q�F� '���ɻX�m >��Fq����t�!�<��-��p�:'R�8�e�S=��nq`x=mջ]r�����s؆�։84t��P�Æ�t�뫻`�	�ob�:M�lf!��9��cO���q�����A=�!���u�O���e;#��mr�k�Tv=pØ�kp�]�!mŞ�wG<���ݎ^��wu^��j�6��Ҏ�s��Ϩ�˶�J.�u���n��Di��NA��AUZ"���#����u�4�s�#��zoCx���=�̄�ֽW�?g�1U�q_a��q:���}c���ԗ+�e��x�$�1��e���6eo��x�w�<f Y5����n3�ҡ�gsU�b��0�����o���0>���k����	$��ո�	'�ⴀY6k�G~��k�aוg���{��v��؂k7s >�n�f �2Jg�g��D�Sq:�D�k�ˡ���V�f�s  [�ۮ�љۿp���]絍��7ɯĀH{�o_R+=�T��8X4U��d�Y$�� ���C�q���sĸf�ڞ��닥i�������|�Tݎ������ >vk�%�b$���*$&(����:�n��x� ���x�{h�;-`H���-z��D�Nd��b��jUq��������d�sJW�<�F�z
s�n�r���!�����6g'����j��r�6m��#������3�\���@�}=���>!~��ֆ �w��[5�P֋ؠ�J�N��{��f�&ޖ�������l��H�̧D�$��d
��w-jX���%���.�;��[���r{�,  {�ۺ���zY3�v�{����7sfb�3�J5��Mg��^=}� =��Ĳ�jk��i���E���,Ax�D���I'��]���g���%N���!2�
'��.:c������;�؁�}v��Y��x��������F�ac����_���M�Q�������g��"�g��M; XO�e�/ᕗy��XGxh�!�&��pNG7�ǩ�I�MC��I#��S�$��Y���u�;h�]ЍDP���30�G�������Wpw��aYߌ�u�=�� ��KP�Q�aq�e�o���S��1���H<dy^-��f;3č�@F�Wu�~����yެ�@|8�viQ��h���OW��e�؜���y��zv'u�w��*�@�b+	$�Z���Āj��Θ�����	
�鯴o=��KV����{�)�9�{K0SS\ƛ�(i]��� ~���n��F� ���b�}=�=]��TЄ�1�X���pvһ����
��[�R�����UH���%���x����k�x]��^�i�j7�o��,na�4���Rs�m�Os3�ߺ��)\ ���.��0�<��u���W�᯴6 ;{}� }ױf ""2��DN�������~%#+�pan��:�`�\�� $������������������r�>)�7W��U��n���%�7f�$��pN� �k�8�G�_� <h�g-
DN�6��S)�ܤ���A�d1�3v�P�U�����i�X5rs����[d�#�[��v9:�0n��+���I�C������_3%��rK�#��k�O6�ᥢs�~�� �{5�&����$�^=�R;�-ɯC�WݿQk�M�VU�#��d��n��6�Ll�n�Y�
2�d�>N|U(<��uXAڜ),4y�'�dl�W�� ^=� ��j7��R���;��D��pL�9���+ZqR�LkƺW��Mg_�� 7u�vI$�Ը6I$ѯvhHbA��w�7�����y�;�UY�w�<X $~�zZ�z�[�J�����MO%��ѯvhT���3��r����7�f�^��˥���^<�` �{�����d�5{��g�F]h��8���>)�
�[H����9wL���_���$�jnhT� {ϱ?��-��dLR���X[�o�R�V�ߙ]D^Gt:��wN�K̃sz��_R��Z"R'�1n���bj�V���=I�����~Q�Ƭ�0Z2�ɎJJ.P�����!�ŏ\q���u�.-�sn:��bƻk��z�ͮ��.��<��9��1��^Lv�g��Hs���]ln����v����k�nX�oN��"��VD�y�9Ԧ�y���2Y�.Vz�X���r��tX���k�pmî��Ŷg�8�XӬ]��1v��۞v���%�/�m���x�n�{��Zd�8v��h�lWk��I�㷓k��Pў�q��3�jq�����\[��~w��)fx�I/O�;�s`k��zZ ���|s���䷳�H��7�-y �H^��]�viX9]D)
dς����w������]�Q��&�#�4b$�~=��� V����z�n���I��E��թ����0^�ׯ� ������[糜S�$��3�Z���^=-�w^���tw�K���]�k�� �w|���Q'�jհ�4H��� ~�^t����o^!=[��F�3�Z�o�3u���)��n��=�T�X��W�|���4���I$�WM�I'5u
�")��*��mY�������A��{>3�lk2l]���=�ܻwX��s�&�8�$z�ÝCT��-�y����� [����9y�d�;�yȨ�?v�*�^]�|�1 k|��	^v��N)%Do�*�O��C/7ޕ~~�q�H�N���-ifWm���8Qr�c��iR#��۹�gN�<��;[̙�nL�h���e:�!l�CP��a�z��  c�_�  �=마��~ō�l�|��?���H��Z�`^�g���3=�@�3W�6@5D��ϕj��[���I�$�T���g/:n��9~��5+��i�����w[��w��=��I&j��Q������NK�͞�����7��G#�¶4��տ*�&�����5��v
Q/��9� s^Ř ﹥��%�[�}�����S�`y��9:��紪��Z��:�.�;��E+�I}�z&{��V�JS�sSh��r�N�d�I$�����6�k�6w�ӴC����VA�MW�y�uD�M0�� ���tGU���&ӘRFM�Z�v$��:o�M~5��II��:����}��ʸ�"QHH2&ea�=�bŀ���U�� 5���'�`R�����α"ne]N"Y�cPI�"3"&�N�ܙF��	̋lZ���lV5X��{j�ħ�64@�I��;GFWV	�(.�h��+�j<�7��Q|�ba�S�=�K�
޽��.������!�Q��k�2v���T޺��g��=�97�E,�'k�z�<�s�\A����q�f����i���&�C��!�� ue'k4PU���%>[kNk�hf��t�b����N�K]�H6�ڗwȸ���]�FG{�c�^��;�>
@�M�� 壡ǝ{w����j��	��4���M����65�I֌�%��:@K�צ����U��ٮ��q��	�݃Wmh�/!s�q�-r3i�V�:,tw�s5�͝�z������ĎW����⢊ZcҞu:﷎ۼ#*Fz��b��`�iЛs'g`��!Llq]h:��uqn����Q'-�wuy�F�Z
���8I�q���Ys��s:��UĴ��w�h=�s�ӏd��� d�EPf�ݢ�eΤ`�xog]'p�k8�W��Ƅ�ȾM�XSS����z�1��6�ѯ�!�h�'��<�$Y�e�F�̰�TO]-+��7�ğ.������.�X�֬�(E��12�]:�� H��6a�%��M�u�,0D�֓��95r��k7w��i��)�.s�����e�
ua���{ւyنS���Ƀ\&��nӫb�ܛ�d0w��Kl���-8e[pU� \m×V�';��N��X�b�ƍ{)ǬA��A$��(�@\ڳ,�m��Ց�<�A8A8�n*�!AK�����(���ݫ;#�]�ihH����Ge��2�[ZtY����,��ʜ����#�XJJ,���v�ۻ$�t	%�4[�(9�9vt3Q	�6�@畓�kf�G�-�PB�k̹)�Rr��GNu�̠����lu�чc���m��6썬&h۱(�#���m�&�m(\����̃��G9�іGA�mm�DL�g[kNYn��f�Qv��t�{ZI�H�ԁ���A"tH�	{X���� �,�H�a�YZ'6�΅���j$�n�3�
N�!VvE	@���pQ��!�ts��:,�⣬��N�N�kG��4����R	�v�JI"�HL��|��^�5�� s���1 ���iih=u٨�v�;G�b�Ofw�^��X�A}�ig�	 ~�4��0h��c��|�<>;��$��z�1 s��Q�XԮZ�i��Z��7\ڱplj�ȦDvc�d�A�
�>��s{=�jYm�$Gg��ݲug	��۬����A�#1�'^�;Mr�g�	~��uU�#/5ט����a$��?.�&>>��6��>�&[�]�<�x��w{�Lϛu[�)���ǒ�$�g]N�^o!�,��� ��s_ �����b>��;��e�}�z��Yx�T��,�3Xu�ذ�$�D��b :$�k�s��]�X��" ]����o]�n���;��,��	p|��w�qk^������L2@5��^�xy!s�^��U�:9dc;�#�{�}��v��%�FD�W\��v��690̵|�p[�*8e�[Sugh�nT�SƩ\�%�D:��������z�����4�n�º��A����D�&j������I�W�Q'�IOw�g��o�i���}���������'Q+��z��K�va��,��{sc�q��uBKQ��|C��",-a�Y4��=��TI�O��x6On���e��~��|c����Vn����UY�]��O<�7�5XrdϠ �?y0�?g%��j��m;�ߦ{vrv���k��R�JSX�k۸�I;�����X�CTa=Dg�s3�7�{b�mp�u�ZܖQ�5�6s�Z�Oik>@|;��߻��>߻'o����M�#Y칈�<�Z��H8K�#��� >۽*��.x���{{��>{��� >=�8iC����k�=O��x3m��7ikki�ہZ�WA�1��q��5�-��E�
���{����[���}"
$��&Sۧ��ywdvKt��͎C%[��9����h69��m�F��ɵ��e䛷n6�w9nZ���t���:z]� �;�m&�&*��<x������Q�m��6��g%�<h^6Nypm���{>�͸#��h�j[���d5u�x�n��9�4T��/.G�6w3�n6���X�[(2��''9�rn���z.ծPE�p�Y�6����Wm��t"�/A�����u���N��ݵ�
�z~A��]<��<�:dI��i(���-ȶ���  ��f,�>;�a�,�)k�{vt���ߤ���e��@ ��`o�@۽*���}��'N����5��@����Uf}�=<��8j	&��8/aƦ���e���2I'���� r�P=�F�v:"R��~s(��w���+�zz{Y&�qg�d��� ���ˎ]�1��K� �}���7��8WYkr�f��]�`�D����������W�W����Q'��� w�p�����ܹ�=_�uS�.�����P��m�����,C�Y��Ʌ�\dl>[m��F�lQG`���õ:�B��G��c��o������ ^����[~�>��~��pl�I�������t��Wc�F|��s� ���ښ���������:8e������u��	�0O�	=\�j�M�w�P�R3,Z�솶���ѫU���t����  ?~���oG��˘֝ﹴ�lo�P�u�>�|�H&�aJ��3״m� �{��|�L^]�H�5�{ �����sܺ�>�z�8������]L�ۜ����oa@D}~���D�}ɆI��S�P>�sҤ:������SH�g[�L�����m?c�@$� 3���NȈO���� �I��tH{7x���ߟ�܏�r;]H���E�C]�v�v	�9����O<�bU�ز\��g���_���ځ��4����n}��7����E��6sz3ܽ���>���I��n7D�q?nj��i��9��`|�Ͻ�n��f�.іI&�?750�I��tH�ݙK�ʟb�|U���W�/2;+���yܸ�9�]��S���p޽w�H�\�uшı��	l�5��v��'��\�RQ�;;�c�X��I�ov�֎!��D��v���{XN�������)����| o���H��Ǧ�vwY`���	��^��&���}��TOI�>���������^�����m��n���G�+�'Uk_k�0$��w�UY�0��6�c�'�-Տ w��` ��8j��=iݵ�;����ܦnSN�ǵ�\�k@W�/7^-U�գmUY �/��p��m2�"Ҝ�=��`��o` ���xn���AMۋ���$�v�c��f\�J�WyX1&y�ª�������>\�0|﹥�� o�p҃>๦
uj�Ǒ�i:��Uм�"�cy�Hi'�g��� Y�Ɨ,���;۪�ϟ�|�1cy�߬���-),�(���Vl���մ+&�`�J�ב_sK v��6����|�qͶiFAܣ5�WOud��$]sXz���UCO���2u�K�H���7�u)`���p�nx[�]���;B��Ʌ��2��fc@�ybw ��w_���{Z�7Ib�v���'�$�$��������ݯ�.�>���|ޓ���=��� m�߬Åk����þ�V�kr�\K�:y��3�[��Wd9���\, Os�MW�����~{Vp=uߞ���qi��'|� >�s~�<A�h�����s]6I��g���&���X�G`o�m�cd��|�2�m�5�Հ�	��oH�G��\�g��;L�o\:����)��" nf�)J�J���5*������E�Vq�6�����v���w똀Z��sJ'/ŎYq��{x��l��4�� �N��A���O T}�O7V�O�<7�6�YzUY?_����e��в���wq` ���ٮ��JJ�zjU4p鹞%I'�7�&����Q#u�g�׊K��	;�Ͳ����O�c.�L#4S�Y�����M�'��4�GoK�norӭK;�(wX+[�	"��d"�#o�I{������	�BY�웰�l���aWt�i.�u��ܼ@t]�դ _+��A��nυ`3tN����=v[�24�]�=y�n��V,u�x��4��:���yV�l`��;��
��㇈�bn�O8��K�!s�/"�᭼ݐ}v�V��ޛ��w [F �r��j��<6{p�:[�w$v�ݲ�ތE���?�U��4ڎjX�m
�c)�m����Kq�ny�8�[\Wf#�\:��w������iQ�U�?�vΚ��7����6|��o���H�;���*e��� Fon<@.�uiE��X�Uc��Ϙ7�ش�vV��,�I'�ژ�1�<��:~8<�\��,�LWzz���V�o�YR�Wk��w.��� �z��� <�:�>w'aϐ{}��H���mvM��J�J����7Q��{����{�o��\X �_=b nt�
�>{]�p��8!<�vD
��s_E/�:���u�� ��ɯ��Y��s�[�7�Ě��L2I>}�I��zrj��w·f��==�5h�pLz�ێа!�R���m���H�nS�/��$m���}~w�,�JZ]6����7�n��X $=9�̔���3GNӹ�\ā�y�W'cj�S�)	�R	b.zvhLY�Y^���\5~)���,�=!X��\�aũ�ʚ/����Si�v���t�w�ZEz�
9[V85�e��y����}9#�ϗ�=�����ww�� ��riA��5�z��{��Q����qUVa��y�� NNM( <��x��p��}ň��D{{+M�D�zr����d���h�׬A3=t�PM�o� �o�< �׸UQ ��c}�L�&�ğ�r�n��J�1�HJ���|ɻ� ��tܽ��Җ�{|�$����~$u�+ ��o�03慛���$b�7.�]r��G�qT��c0o��C���;78�z������HH���R��o:�D� ��T$ ���X�y,��o1��o�� l�r�@�uw�,��Z\y�{�2I~�T�m.�S�! �$�p�$�&�l�6H$����"���^�̶Ϝ�8ݪי�g�h��~�q DG�+�v���[�����b̢�;��qwO�˾}W���);�MԤZ���sil�� *W��I�8�oP{�������g3U����S���_j��~�� =9t�ρ���]g�{����)I�!.��qy�����@�3�@��Y �z�uD�&zg�#f)qgy�π=794��e�l�5U����K�>d�H�3�P�(��h��'�5��k������7���1:?>K��t_�N��f�e �8�Ud��]���$Tt'j�!�M�>�����e�uHJ�����5����K� ΋���C6	0ѿe�@TI>��x��.�(���)U�9�ko z򹽁�70O%�.*`�" �n���DL��@S{]����W_�Փr��V�i,)	q�{}����n��7��}�����|�|�ys�����0���l��"�cǯIӝ����*���_[� �5�0 M���Mh�e����{�w��*����.�e���4$vQ�*=X����������ʗ�3���ʸf�����4�(<���M�	�f�Fk��+&L@����賳�}�~��q9��=����@[�UV�y��>��;�8i(E͝���}'��TO�g��'�����oZ彜���'�N�9-"c<;8:N��MS7��-�cMQ��CC`*䬲[��=S�檷�_5�|�7���Ń`O�ٚJ�|(�;��U��=�S@/mv��%N�䪻�̛����t��s\�]����?  ���f F�g(0+��)9��{^��@Z��0�WE$U[0�zw��y�7�I�P6�9ބC������No�1 ��߬�uw����\x��s�]�^��� ��s0r�z�z�z�RȒ2�pBO�}=l�_�����"�c�����_@��Ng����ϐ��V_BL�=m�����$����0�Z��z�5ӷ��B��f�` �������Œ�ajK�P�D�I�U`��^�9)�p�֌U����A�;�5h曂#R��Z(.]��N�:ޖ`l7�.��wZ��ok���ʧA�F��;���
���n1�!K�Ai������kA�[*i�w�+��`<��Aۭl��Y2��Z�ã��"��v����޷��Ե�1Y�+0L��fĀ3���2�zc��[��\/7{���9`��ܠ�c��һ��09&P�!Z�%MqZ�C���I��t/#�쭚ƢU;>B��[�dy[����$��a#!ԝFwde��wV�k$ʴ�pb�Z�����ڑ>��]K��*Fλ�:���<s	T�Y��^�8�Sj,�L��fT�XrT�Bd2���7���7.��dc�ǨR��Yw��82$aݙ�cŰ�6XfDcƵ(W�sP]�>��yfT���foꅳ5�������sZ�g n�2��sOp�ڀN��W���*;%�ұ�Z�=
��eX�18�-�&�]Ʉ���c$W6U�s�����ރ:(61\�������7l�<1��	�ll�h��L׽�s���h�_f!��*�SZ�v�B��
.w�����lcV�]k8۳�����)*w콀�ٜ���2)D=��&')�6��6��.����G����SVd�7c�}r"ufu&L�����F�L�e���L�R��JR��FT����i�Ώe�t�.���q
��>�-y���6*��}�ّw^��ʵ[y:u[�R�o3Yb1�	$��đ�і�FaDSk.'(�#2����8��+��ʀ8H���r����wg'fI�V�Y�$Qe��Y��X۳�"����8yYW�ZI�G�s�ͦ�����ν�D��d��:-� ��ۮ8��A:(�/:󻎀��^ݠ%�tu�
tq�rrY���E�Y��ĝ�ۻ��e�A�ӑm���2.r���
r�;���Dw��Gm�.$�88�..K��I�eF�'9(����۳��,��)�=�t�҃3�D�m��{k���r#����{v2ݝ�N'9�Rq��tU��u�bⓜ�f�;��{ wv=����![yD����s�K���g��eq�;{��v��7���R��Cl7���:�gģUsa˩aw�;m٬�x���Q��neݞ=];n�W��<��v�غ��&�����y�z��	L�F�s����G@w
ݺ��i��8�p�v�v�%c>6ζ.yg�v�٠ˢ�5�im[q�nz�E\�t9d�����;v6R�ۭ˷sǴ�����-�޳���[X�v��5�{��x���]�%�m�*,��ק��W�ĉ��ݵ�������X�]b�G�3o!��Ez����4��閉!�U��g�������:��myE;u�f��A��ݧyxU�[�v���ے��ݳ�����=�̈́4�ѹa�-�J1��Nծݭ3��&�.�͍�4t�s��c"lc,g�jmE��5u��e�m{t��ێ3x^:�&L��d
8��݃y�8�m�)����g�Go�]����n�v�k��9���W�7bE.s�uؽ�Xüm�V�p�`j��ݮx�:ݻ�Y�7�����A��ki�T��Ur����9�0��S�����.���ϝ�Zo��0%Yj ��QA�y]��ǟl�O��[m`�Z�%�\�.�۫���]�.��:�;�;�g7*Xݫ��p�wP�wm�,\�XwY� �] s��8���@l�
( ����5���ٔ�c��.�����v�����%R>ygPp�Wc>*�6wVƸ���nL���n�\���mt�k����=l�A.�q�h��N��I��NۭWV�<7I�N2�fZ�nx^BV��n��Nc�.�
��Z����r�˘�ݞ�s��%�R����ƺ�����q�ݚr��p��CJv<�Z)�<m��k��W!�k�-�^�+o%u����$���� �]��T���Қn'Y!��
=�h��S�=\�O��o�q!\y��iӋ��g5�gr�l�Ĳf���z7k�zو�bw��M����K���经���qqnQ�T�,��7;v;A��맜�����kq�/N��gscAF9ꍤ�[qn�P9��4�N�<8�nd��pj��E��&����\� �z5hyۭ�e�s��M��ַ8͞3�U�;�������� �l�M�ys�����pm�½]�r��qy����Ęϡ�!�`�.��<x�`
g�4�Kga,u�V�Cۚ���ڧ;8˼DWctJ�^S{u�ܪIK����u��u=�e�����E�n�ԕ���2^vg� �{n��$���k X����U;��nf �������X��V��Vט~��v0b��J�����+l>�N�A� >;�NfA�=9����>��Vw�}����n���W��M�@�g4` �Jԝ��~�^Nve����w�6޾=�N`�k�YYJ�!3q~�<�[��ۛ�#��l�G au#�ŝ���A���ִ�k�o��.^v�J��}x�\v�Ѳ�q�{۝Ő�s~��Gl5�;4捞�m�I/$�;����ߦ`(���s�Og|�MCl�)�%�¸�8�MZ�b}@f�K[,�AZ��:�%��{��O���v�_|d9٤� �{��d A��֟���V*��U�+�!�^�V����hmE\�:��K�L�H=�c��r�g��96�NX*��;!�تu=����UIV9��y@��^q����9������I��Y�g��ǋdk�Ygo��h5���	 ���`�{:��$����r9�+w7N({<�7W510QX��[^b	���#m���3�.���/-�3���	���� �&��zۢ��du�ЕW2��a��gW;�����ߐj�{@ ���k���'���Y�+���y��M䕊։E�0��71`|����<�r��w�{Z�G���.s.����f` #sӓ^�14�Z�}�1WY�2�!G�{�k>��k�2�|/ݷ�B"�Q6�el�HU[��:���--u2�z��s�� 9�L�@I2��e�Q���K���n� {=3 ��2�v:0�Z��Ӱmݮn�{HZ}Xf�n��$=�Mg� K�� �7�k~N�mz/g����W Cq��ՏD�g�@C��T@U��djҼ3&�V�͓oe�˸Ч�	\yք�	�D4&ѼYJ��6���rl�ې�EJ����B��Ovo}�q٘����3=���O�����g�]}A{��)$jW�Vט=�2�w�Ŕ��LX6 r{�i>��sS�<���}pi&���m�=�"�]pN�TsW�7u���>wn6zi��a�W�~T�|I�z�l ĉ���A$������wa�ʍ7p'����}}刺^�>uyfK�6�d��p�j#OB;Qʎ�n8r�%���v�~w�����(�k5<zs91,���9koH�����%������_��  	�6��DY�9�(��>��t�#�uoQ~�Հ =�[������6����u�U��{���ղ)HQ��ּH����d~�L�I>��f$u�T ~�.�1 ��=q�\������FP���s]��n���u�ww� ������f�O> �{�A��o��wy��o}G� ]�4�u��]���y�l�]�]�6��'ju�r�|��#�����.�EJ��@��2��7p�7��m�2��Tw:U��F��}�}��)>�¦ݵ�f�t����m�34m�	o�`a %3 TI���l�I���N�Ivw�ivf�I�6��v3�=��)��ޑ��g��8�nܸ�*� ���V]{k�x��*GTgo�������}��e��m�6�@�l�F��]h`7���}��nJ�k��L����0+�{�w��΢oվ��� ���0�I���l��^֫X��{9��{�����RU.<A��w :{��� s�h�=�[��[���{��,o��&���dR�X�*��{6���q
U��)�5��b�F�s�$�E�k$.r�&r�����`3��s�M���k��>� ��_+\���$��n�	�h�	<q�B�#ֈy�"�:�Q'���k����q�9P��&��74��v�ZY��;P�U�;w:Y�'m惄��k5Y|�5|���=��ctd�5V�@0PD'{e��ԥ�������z��-*<oB�v|t����W���;/�؇���m���Y����F1�m�۝�.L��㝷�.�Ӱ%�tr�v�]���<��n�-�t�%7�Svkd�<=��/^��w�5�^���_-5�k�lvX�Q�ѳ����v����-K��x6.�M۷a���:�J]�[ۧ]�9���1ˣ��M���zܰ`:سNv�틶�٫sDE�R���M'Y��69�s��T�T[}�!L	Fa�#�������"����uו�eF��z7y�N���'ݸ�ᐔ(
$�&.�5�H�%��k��o#k��{m  𛪲�+	ɯ-��,�b=�����%l���}���'��H�#n��\c�8��kk�Ap��|I��G�/'��S("��V;k��~�Y��<�� ���>��|�^�E�6�ŭ�7W�/,���^<w6�� �u�jO@��P3A"�+��$���BA's�.�X�C�؅��f�=;���k��S���M��v1���^|]���淧S�[S�ͯ��VT+�a���o�(8}�| zy�cU��8�}8�z�
k��۠����J��+�s�����>�{UY��fV�!�r�T	�'�Df��{ �ӝj�NZ�SZ�wb�*>
��M\!�o �#��»���mD��gj�� �Gd� ��zؠO��j5�����"��0e�eX-��B��窘޽�ލ���a�i(�k��sb=�����"����a[�����t ��n���WWԧrYb���~s2�Ϭ����b�$=�h���X��T�t'C��� �<�� ���T ƽ}����- &��%�U4���S���Ӹ����M�+v���#@�,v�����"��7%V?=����$孊 
�����f�=4���;v��>ctTg�̑$`+����$'?D�t��A=�N����j�	Y��5�`�uOLnפ��P2	EB%BD���Ť��_�G\)��$�p��<�+�Kk�(��ɛ��r�G����f�b���-��:�72��Z���������uk�Y��+�f�����쥬SB�g;�n�9��\�z�#���wd��sy� ��NB���
LPJ+_f���)���%��v��j�$��A��F��~�e^�7����GRCI��wI����3&�Vn�QɠV�)WU��Q��g4�f��Y��y�|���4ԥd�,�u۷`�P�6tn��1I	t#�ݐHpv9A���Ԥ�B�BI��B�mu�F��Do�W��[��R}�݋$�օlK��$)1
��VXT7ǵU���M=ϝˌT����O� ��T	���^�AZ��e����nq�'�тA�>��0�7ת���!�i�3�|q�g�$諅N��$dc�"�j���JQ����{v�23�:P�N�� +x�4��Q�o-W�b�֨�ǤS�Neme���Э�!������8�󒯯�=X��7"�:�+#�ڵ����|���~S��Tr�,5�8�˵Q�̜V0e`9x:��@Uw(�w�c��9$��j�>'�61АA>��˰MUh�r\\���8����ժ���U�d�÷�-m��u��v� ��͍�k�[������F�zB3]�P$�1ԂO�:���e�+X�`7�?H�3jN���(��2��7x�s��u�����o��� ��g@�QS�]�<t$��-�/�0Ȑ���
Mx��u$�ά�,�(��QB���^���v�TO�r3�H>'ݝYw�Xգ�}$`+��Զ���H+b���-�e� �sy�{>�o�cI�4w4��9�i��N�����.��$�����Em���2���D�m;�H$�j�Wݦ��#'V�g"�v��ݓ[�S��Ǯa�ת�C�ISP��D_��X�1T���U�!R��v��� /+J����=}�F����>\6��RK�vy���0��vy���y��=v���y��b�6�ݸ��g����iN5�ۉ�0�\��<O&_]q���h��׳�s�Šz��k����:�==p�ݻ�nohz�Ӵo������%5c�t�l�&���ih�9��g�6��e���v���֯%�OSs�n�;d���t[=����v{k4Z�t9�#�>ٸ���5�Q↴����۶^��Zn���~q�!�����J�,����T�j4�;�N���^:(��d�w``_;�� \�Q�Fd&&+ū�C���{�^�( 7ݭ�� ��}B��9�k�w|[ٽo�׮g�,�XX�Ism�زH!�j���V����A#s�ݒ	79
�Yi0����F�PrN�Xw7��n�$��H=��Q'�cYz9�r�������co��j�5���&=:e!R��#;��$*����W�g��* �{b�	�s�vUw����V��5S�J�@1ƌa8��;N�U۳ֺ�3��6������_�����!(�(��-̫$���ē�������j���݂	�T	o��!4�������Qkǳ6��q���pf�+{�B���縏'�����w��R}�\tu���k��ѯ�q#�Ζ���h[�")���2�V�Sl��}d�AݮTO�퇔$£�j���lU'�$�((��w�Q��b�Q�ueM[�:m�K4��	<�믛���ޣ�����ҷ����9��6�nq�Kư�$뽸�X}�kF�&jڢ@螜*D�LH0�Rhۓ�qu����#�z���_T	:�4({<�|h��`CM�^��C���Z^G��)��턓�u�����:h�vv��ίs�N ��[X�y�yۤ�>9�9^�O��.�v�ƕ.��zޠ5�ۂ75Z*&IS1*	�h�.ό���fһ�S��}\���}oVWg�7T (��E&\/�����8�d/J�B�����5ب�|y=ʰI�M�����S"nS\���p��Yzu�����۷Y����%�bdo*���5=y��,ޔ���/�{���������9וf�]��UgL4�:���ePɗ��T�&{��pW8������q�Q	��{/[ѭ�kw�eb6�T����L�Bd��4
T�ƥ�w-˭!�^�J��s�[&BN��3��!�EP	Q������d�vm�\<��E�oFl�6<����mSl[kY6�I��i�wf���e��j)䜘{" ]�v�l���3gSvE��j��au,xUa]} ��v�WE����/�,-u�AI]��o�%������++�hr����1n>�ڸ���l+�R^*r�Lx����N�:����Ӿk���!]�CÛA�*�i��d�ٻ�j�I�{�w��0u���-�
�m��Nb�μ�Ǳ��ރ*�����%JXR��ՈY�}؁;�w۽��Fvp���ئ��6lg!��G��륥����3�U�BV-��周���:�`n.y�Ԑ�X�*Eݦ6��oK��1-%!���rZh7�Ib�{v��m�y:�����c����˷�˹��\5�⥉թ�����eܔ3�=�yv�y��i`�7q�;�8�P�Ǆ��_o�%Cˎ�F�����	��Z�;��zt3��;o�'�����޾׈vh�S��z;� ��Box�m� �W#
��-�b�m�^ꂤ����ڤ��uV�f5�E��ӓ���浹��
K�;R^��K��X��x��O���DE�Q�Ta��z�$Eaqmi��u��rG��'ZDqt^Y�u�@��%G�t%֬Β�r(���3��A��A�FX\��P\Ei ⼼�;���
=����gVZR��L�8:=�W�u�۳�$��(����,�˵9��;� ����3��:�(�ζǚE�E=����*��++%��%����qE�YC�[o4�,�:��{�+�b;�;�b:3����q�dVQVU�ppu펲�㻎����YIŕE��w[k��tV�>T�X�d�>m+st$w* ���d؎˓�
$�*&>�o�3�! �$���$�4�݂|H<���@���Z#���`rrР.hV(2!��&e]��œ�ݥ^=�WCtؼ��� s��@	w��`�H<��r�ɒ.��H!�(�"J[\��;k��VB�F���-Kv�\:�N��i����0Q1 �EI�\�
e�:�I:�� E��8����N���$�e�;�Hcj��d%$`+�{-�@��!��v��Z�Ē	�� �|y�*��헽���5�mw����n�ES��.�c�T	��MX[��H��	���H:���|2�J$��4Kt9��C٩Mf�N���� ]�m�{������w���$h�!�\�]�ad`/s5�IqmX�&����t��V7���\r�Î����{%m��.���ժ��|�lFEc���2eAQ1@�n*$�b�R�R%i��o�[��*{� �LT9��h����?�X`�vsݹ:U烈ֺ�[�Gg��6{.�i�m l���Ua����픊����xY�>#�үA<�(Q����1����A�{Ԩ����
`�"A���;�S$���+��aK��u��A��^�{�����<�Q�&{���V��]Y�$����춨H̽T	�ë��7}�$���* �yޡٳ2�L�&Bf+;B��)���0Ik�	�2���l�m��=עQ�vN�x�k9լ޺�ƥ�;b�泷I4���틹::�uQ��z
'��b�A��A'�vݞ�)��bT#"N�98I�;')w]�X��R�C�3�]m*�� &�4s�\�U��s.��X���s֤��Qۼ���G &�@���2���/���O2oW�7A�]g�WK跓ci9l���t�r�ݺ�۰�\.������Ì�L��L���<��Z�p�1v���5͎�[P�����U�`uۃ\��s����]�ӫT��}����\�s����|���{E�K�u�g�n^�uϭ����-�q�v�EەN6�on��P���t�p�a3o�r��Cc�杻V������7,�/=�:�:�����������:ą����Q�l���+��J�:=���(J��5������NX�� >�K���'���i�����T	*��RS"`L�涷��D��t��ĺkIn�P�F�{�� ���ۮ,�js���r\�!A��RkǯZ�A'*�߬3�v��C��jd^�* ���vHcj�"$�TB�skjD8�;k�׻w�͂L�5D�C�ޱdw-Oܣ������7�|��Z��ɴA��A�5�o4½��tk���;�"�@E�[�<}��	�)���-�߰��Նޑ��ƌ��]���QQ�׬q/��w5BԒ��~��K*e��N�';��&��j���
��Z��>�=�U�cLj�$�u����ȟL���A!1�v�|�a���z���/�ɸ�Xi�Z���J���!:3:Ka�NX[������ſ�5��4�X���x/q5[�ip$ݻڲ@:{j}�nL�Vd�yY���Ҭ�@̥0&ʫ.�m��>/�j(O���<��<*������fw>��ut��AX��]�_�h=���z�����&��п}�z�n�(��"v���]ՀK��"@5f��m���i�	���r;����@�۫� �|��$7j�ue�'��kMm�jE��%bv���[�^���ێ�n�.��TÕ�*��h�2��w�'���pQ� ����9�4h�H'���V�"z�भݓ�@Ǫ�u��*P0�$"hFݬ$�gT%knψ�٣^$��ڠA$Õx�i��V�970D�(J�=6p��^�٧W�͆ �������/�&.ѻ�R������;�]����RkL�L�)�4W_kgk�u!�n���%d�z��|(}7��	��MQ>�V#aI32��12���u�$�;���ZE�N�$Ct�P�����ãW��w����=���".��as؀�^Z����A�S�ƴ�$yw* �]N�ǵƞ�
/#;���j(�q�Ωm��>1�;\!�h��F5.��['�8�j���?&(VX�;w��q �怮]N��vv���۲_�6y4���.�o��. #���}��7�܌�ν�j�p�.u�'�ʝ�$�"���u3����L��
�m��b�{qsb� �ԯϼk�J��OU�Ἡݛ��2�E����"�<>]P�~��� (Wn.�$�'\��̒��,ڥ�0ܨo�/��1�1wc���w��s�ܕ���v�W��7SS��r'�nr3z:=�l
�q �:>�Ww��e]��:۰K�(�=�U#za:5t��V݀H�i
5gU�4%��f�r�m��U�������m�RZ��fs�g�UNq�k����[Z�~}�yu�i���Nł#�j��]�,�l���n�A>��ߋXv�aRTMX�n����O[}u��I��S���-6�J��^v�7�y�H
�T�r?��^��@�s��$f���pD�t(��VвGOm
����dJH��/�GbtX��z��ї���,/W�ON5Tƕ���>��۰lN\�HL��
i�m
$�ӭ
��#sE� ��n�Hs�B�5뛕,�M�=@x8��m!�l4�oV�I�ƫ�{#k�bG9�3W����0�0X�ʝ]�}z~��0KP���U��3e*.�E�3r�"�w>1s�wo�:��vA.{p����m��c'mycq��v�Q�\�-��s�7+.�'>���u����6m�-�e�Ǩq��Ls���WnլJ'g�v��Ϋnwm׃�b��m��k]=nn�]Q��m�m��x�;Rt��['�W�z�4v�-͛�h�[��1��>7h\��̤�+��7�-������������ލ��N�: �G��,C�]��3�>*�p�i^E;jFz��pv9A�9���)%��Gu�{^��?��(A>$�u�1Rx!��Tݾ���yR�+^Q?�I0]���$�#"ƽΪJ�+�$�<��'�5G�9:��t�:��'�Lĉ�*D)*&
�Nb�@�!��ReO#U����Ă��(H=��'�*k���2�D�z�����v�n�M��I>$cN�D����
կ��1R�- H���D����D���*Q��n�W� ��Dbs���^�����	e* �]�'�<�0m��n�t��$B�$��ƪܹ�E�r��}>�����9�;k�e��3cv�s5�d$&RE=�r�A>/���>$��Ԟt�b�/ĂAn�Q>��B�	�����[��e�u h�h���Ff:����3�1��;,9oSb��C�x(�y���$\�Vk�@G��a�or{9έj[4��J�O�iТN�yV	�{u����y��7��*��PZ�z~�9V�9<� ���3�X�A'5ڠA'��o1��=��E,AU&_gj!��39R���AŴ�ĂA#�o.�=۔6^��>�/��M;���|�,������0 ��ϒ�^�٥N��=�B�${yV	�=۔(�|�Y3�����=q�����s��̨����W�8�7<Mչ'�bƄ����Nu�-A-�ɞ����A'^�]�I۔(�
q�><f ��|���q0�P4l�{U���d{w\CY�� 
��Ͻ�R� �K�9�My+��n����.���Ϲ� �HP����Y��:��^T��=X<�W��Vap�֪9�w_u���a!Lu��.��5��cv�F��j��CL:��	�+'C�V8�K��������wzZo�.U�@ak#�}������9�+L�%��b���
z��3�sv�"��0IS{�~%�y�MՑytNVn��/���b���=����݀K�̫�۸�xO��ƫ��=�7��N�^:��q��� �	�|@/`8���3,H�����7[x��������}��$p��xW�`�w��,h3s�eLr�˲I�(Q63! �RHL݃5z����<A{���bI-�P�H���(|4��S�V��֗|44����2��=V�x�OV�Db9��$�ٺ��f�[(P�������]_]�3%��
�v�e;:3�������@�5R ���³��Z|V��j�(]�__�+���ԋ�sY�'�C�w;䂲sU��!}$�k�s_+��w�ia&��'H:�}M�p�&=g	 ��l��ۈ �Su��C]�pQ�A���(���@A;β��r������u����ߚ�R�m� �ywd[�&��8��ͫn���gT������/+��AD�U�У���@�	�u�~9)�r[@�O}�N� I �j��p���Ț���l!�OU%t�׌򰯳�@^��(���*����7t�M�Gv��s2%�Bf��ު$9�]��&�>T�}F�����q�*�y�݃b��@��B�S%5�YCYI<�ˁ=j��Ov�]���3}#E���ʀ	�樐�E�ɉ��D�a��o���!^!�j�j����T��)�Tl +���y��Q���8ɭ2��� �-bmȉ}{U��k���B3S��5��YC��{X��[r�u��5�Bm��g���CٜqH6���K����K�E��5{��H�)���%��³O/��Z��TiK�S΋��Zޥ/1�@k�U}�.�oJu}[�4��b���/�\$ �����J�}Eg qv��k�}�Oz��g
=i؛3ج����#��2�dJ�\2��QK�{&#�4κ\�Մr�B�VL�;�������m-�c-BT3v/n��X�9��˭ڗ omQH�2oQ=��
^��u2�
��&_'ǵ�tMa���i]�졣%�ա���J��غ�3/	���\��f�7-q���Fqඦ!��ӆX��I�oMl�~nҩcj�L�ɏ"������nܷ6�HE�B���\��E��"f*�X#0(ͩs#X��ͫ��+)-��BV�Bc��!���C��{'n6��R�]�ϖ&V�A��˷RW6���9 K��8��8=Ύ\�eg%|��u���&o���2v�i�����mр�s*���E�.�j��j[��.Kc��hj�����3�m�t�4/mv�V�����Y��(ޭ7�k�ؙ�p��'0��E�8���j�� c'H4oqO�ɨb)m�un�K���gk�~���j%��K��ITt��y�x��m\O-]�=�ͅ�e��Xp](��0j^�iËy�̣�>W�J�;$�}��|��C�5Ѭ�\c�;j䏡�;_�̬���gE�e�E�Tu�fuVYQGivVtgQ�w?sڋ���Yu9��A�}���JK�
��.;��m�wYM�����(��;��.���̬���vy��ո�m��� �:)���pu�wِu5����Q�q��U�w��rq|�S�:�*�����%����������:��wλ˽�:��{v��Ԕwwy՝�+;��	�q@GIQq$wV۶���ȣ�$��+��
..$���+THYXq݇Vt!�w|��'t��N�&�m6�r�7UM�"6�D��۱�4��v�Ȋ� a��B)�w"�f��=�ٖ�wll��IU�N��H��ƶ:��FL��wnE����[K����Z�6�k�i�n压����k�7�:�c5�*��1�b���mn�y殕�غ��������[n�\��o�r���WFnϴ�up���[�&"Rֵ�{�j���˦���s�U�Q��t�����G�a�v�g�wW*q�6�k�x�7�D���]ݰc�yJ���:��sQՍ�c��;5�8�a*D�Y�D��@j'ە糮x����bdܪ���W�k��<������m�N�k:��׬p���b��U
h,�G=<4=dX0�4Z�:�˹��������[/�huŜ^-�T�R[����V��۶�5��ݵΨ���$9�p��b�r��C�X�v��۲�m��Ƶ���:.u1��;ٓs�5؁��{pd`	�ܙݜ�mb^X��]j�D%ۭ��m��M�K���t�bX���n�7�zu��j��n�0V<�
ܵ.��7�{yۨ�n���;�s�2�Tק<�{�R%�砇��m����Ǝ�Î�m�:�]��n��LN��]WY�-e1g�vD���!����n<qŰ�y�M���ˀ�m�rA���`�.��
1$�����/_mVA��<�9N9��i�[�G-���S�[���|�����b�nå	��{F�4�Yn����r̽���᳆�Oi8.I���(d�F�X��*pu�R�z&�{t���·�n=nV�mۺ��ʝ/h��Y�iv{5ěKn���4�Y��=>����'0��<���=��$]���y[����n��<%��ޗ�U�ѻu9x��5���8W҆�w<i�� j�N9��Q�����QcyG��s���۹�O���dǰu�k�f�c�h���:��cb#o\�uGY�β�n�lԼ�[�]=Cih����9�qڅ;M�]/��ڭ4������k����z/
q�oF���n3 �u�Gk� m��)��.��h�=]���n.��G��O�ӳ�۟U�mm�3�S�4���٣�r:��8��>����.�vv��[/n\��l��Yu������fh'�3��ѻu�DGK��Q1n�x�K)I�On�N4�g<u�F��G������k[X9�$��9�G��~}���]1�SBQ�֨�I�u�d�9�P�b�W:����I. ��_:˿���drB�
�3���GI������T��$v�eX'Ď}�b/�2[rǠsq}@Oq�_a`]�Q6>O]0�s_����w���à�M=���$��D�v8K��(�JR
,Em�t��Yd4 �um��_^Р@��0Vǽpd���w6:Q�@�
aD��n]
� �{^*�w�'=��b
ϗʅzl��G�6��:��v�XR�F���C�TmM���l;g�e��s�y#�8��G	~�Ӟ������x�w]�$�|��#��
/�8�l,��|� V����ʳ��A9���Ť�F#�7��N*5:�]�r]����WB����~��8����aMљ|�b�ES�̮Vv���w��@�0B{F����I
�O�j�<H��(�;*�1d�8S�h����kjg|29!b�T�u�U��g3qQ$�v�����s4>�}B��<T	�s�6��&fP��*}y�2�彪��ZQ�eV�O�� =�^ ���&�^l����UA��J���]W�2$$�J���7ب�>���5�IT��vH�]B�>�>��W�$���y�y2gj�~��U/̴��B�Ӟ�
��.,Ӓ:�8�l���W���pR�]�����3�S
$ ���ˡ@�@;�A'{o(Oc�S�l�W�h���
���)W�P��!\ğ���cO�	�a���Smc��/Ă��A�yvH;�����~-X��;uP��Ц��w̤	�q�1@��Ľ~�Go)�)�zv��\�����`�����i�_'����.������*�6���ͱ�5X���zO�6���?.�Ǜ.�x�m�U�	;�ya���&f!H�A\��W�[~��g�\�r�B��R�	�n��(��lW�k�Fۉ��n���&���N�{�e*Q�b��|y�K���'B�v�*C�G~���h�8�if���=���Gkey�v6rnz%˶ʛOQ��$�_f��
Z�WN��^��>��Ֆ,����
/:`����x�/���H�Yv	�[p(��2J��T;k(�}7{�����	�˿#_e
�%RG3˸��i, ����Y@,��\^��Z�o����m2X'NO	����4�q�˲N����Me�c2�$��p����-n�&����$�}�/�A ��	�'��e!��i�M	Y�L��7����yuk�s��mŚE�oeD�ыs8����G^���YO��<��F|�7��GuU{[WYMj�]n_o��6��{�) �Y�o�+h
 H�*ӝ���|�P	cm� {z*T =��XV��	c	�,�l�uv���Ek҅�<��:K 5F�&#:��0���ߏ���D�k�3����$��^�O�n��5��t�}yUw~$��B��p-I%)�QQw�5s�k���bdB��
��,�{z�  ��R�N�{cG�o�:�#��(�*B	P�D���r��@$�=p�{bj��=�I �f�[�!IJb���b{�}+�(�	��	�w�a�Q�QШ*���:Ս�llЦ�}��j&���i{�_f)�ڹNb��]�!D�H:��H ���7B�n���xd��s�+�:�ΰ��	��Uc�E3F�ln�jx'e�l��P�W�C��_*�&.�IS:m�qd��ѫ�w*�uSKSCo�q[�2b��<��guÖ��k��x�	��+�'��5Q�kU��s��t�k�eWq o��エ�s���O���Wkt��u-1�ݮ;u]���n��
5z{=�n��Em�Ź���5����I.�y���9�Ӵ[��]�N�%y���m���=jCS�w#��.�z:�8�U&�\w�����ϳ��W4�nnƝ�}�{Bi�//\t��X�s�ssظ��F�+��7g��zNd9l���}q�Z�;��F�JN��Y��i���ޡ� �w[˰��u����
�{�b���[�	�y�M����AF�ק�����9}!�=���^�Z.�[��uB]<'k�	jfdH�-дz+P=��`2�`;0kc'�<�H'��U�-��f&$)�$Uڲ�����]M��АA#��.�'_]	���
P�(!J����)0d+��v��Z{-�X91+���>��o���񰼲��������L�<��T)b����Gq����Z۝���wK�v�d�߹����B�}�Г�Aͷ��O���Q��)��3[}���7��k=��X���6�4H�,��m���R�>S�V�9�2�� 9d1x��)a���&�+��Wl���#�oy�v^U��a��+(�.�(�����5���8��xo=���(��t v�*�m�ֈ����>�*o�"AJT����a>=�HQ$�!�~��rs0 =��t^�%HE� i�2&0BF�Q�.�Y�F!����d�F��
$t<}�K�bGC�Dm#~�sGy+H���U}ٕm���yBf*δ�������H��_
'��{�]�����7އ
���h��{�n������n��k����F�$Os��B�43����)(�WŽW�|[�B�Č�y	̃Ne?Z��߉�ۡGTe$�RL��Pf��;B�����r�__`�A-�ר��*A7���ߋWk�RNg{�O�\�X"F䲖�M?r��Eb� �����|�\Oq��������5'n�P]��n']Yg��6,M��x�_s�͵�/1�=ݞ�sP	{��J�&W!���9�����
�|s��M晛D(�BXM��ɉ��'+�� �L�@T��4A������gv�h~t��x���.N_�j����_5�o���k-��fW%��5{^�N�^פ7�݈xβz_nK��s��"�$-���5-�����TzY!x"	�7-�тr*)3�}�`I2�Awj�H'Ƕ-АA��u`���
(�P����.��Q��[�$���ԭ�h2�|�םō�g��[�{��L�� [�K�>���LY[�&��F���g�'�{V�Y,�����<�$R��gX�1qx&U�I%�^פH��w`�1X�"L�2���]����5�v�3��Q����g���"��v�*���.ЮfOY�;�fj]y}�B�UH6�*���;�v�E6�Q�asQ)®D��3�ጻ/XyS��V^����؊C�"()�����++�_����P����Ggs,�n�
���w�=wغ�
�V�� � >��V�5�yDDH��H�(ɘ^��{^ͻJ���n۴@ݜr�46�v6P��c�C=ޡx(d^����+{��nV߬�I��P=�k���5��F�����@�$������/�s�N��N��Ce��2��I#_U
$�w�H��1
������L!*L�W�z�]���R	$���s��$��]b�O��W�5+Ad(�K4�Ӝޖ�����t�~��$����B�$s�s��8�v�H�n���� �fRP�*U�x]�nɛ8�q.Q�}{@������U
�A�/M��w�]7#qy���:C�:y�9"�r��p�U�L���3��]-�sOi&v�����H���9��f�z�c�ruZ�]n�o*�t\:�я���`*��q�y�U�>��k�Z|d.�9�/<�țWm�չmm>-��ۙ�\Շ����q��=�ƃM�ui�@����{mY�kg�SȻ�z��KGR89)d�vi�x�̝�t�� ���\8{kN)�3�3�[�vk�vz�n{ggZ���=ɱF�'+��*��ba�ܺ0���WTr\�r��[sxV��=�u��ng붊 ��
��l����u�Y�m�p�Q�n�=���%���_lT���W�N�y�����	�M�7o�b�Nk:�V�.�$�����!�*���R`ҋ���UDfe"���o�	#w��x�s��	�6�V��N�+*��I[�������{�zZ���|��m�9��kɈ�s������UG:-פ���� PE�*���H�UA���A'/�>$GF[�G�)�x�f^��5;��i&�Y}j �a*�鳭���)�A�����:�(Q ��_H�w���~����ƪ��Qw����;;��8���d�a����� ��	ˆ�u�l����l߻�	���rk�k����@"�I'���]����+r�*�РI �w�(���jP�!D���`oywXLh⑳r��9Fͷ��lwv�	k�)gU3���	6�Љv�]�U��ej[�d�]/�i��m�����Z��wX��Hm��48�N��I�N�p侐�[QN.����A�"�9�tإ�ʐ�>�sgęy�R늚��$��2A��'��N�RQ�" D)F#*�(]P�4�'M^R$���ڲA�ԅ��U�C�B��&�PT�vA2�!	(D�T+���R����8%q�q��^�	�ܭ�$���5}���s�̬���ߦ7n��k�\>|s��\�:����v�N��Qj	jh��X�}���PTF��U#����A��-ݐO���B�5��ajm�:3�A;�}B��zf�&eL)E]���R���'f����� �=t���*M�s��^�[F�oINqsVZ(K(��e��۴�|H/@�����B95f�٨�2�}h���lB��2�32��V���+.%�kVԫT�&�;��9}�p�z1��;
�KY7Zƃ˂�%�5���؝�cw�*p�'ltQ,�ee��ẉ�n鲶��kc���dyx%��.�¶��Q>F])�YoJ�s��^�Y�U�S�4Q�ջ�c�ͻK���r���a�7��5Ɗ�gr�0����sn���1��9 n�h�0A2���#�k��m�'j��٘�B��R<�A˧w���<W'o6�	���{����E��<�gJ�
"�Cy����Fڸ�%$&5��t�?��x������U�7CJ���b���{����#c����S�8`�|����qҪ�JVXq!Vl˙7\d�,�v.kWF�`�P񓞚0t����ɜ�e��\6'�6�(��/.�d�t$:�1�F��ׂީ]ۧn�6�<��YTtt��"4L�՝�����h�����:���'�m����@w�G�m��.�R��� ��6e;�V���O\�c�2��4h�)2�j�Y�����e�Ĺd�*��2��Y�hs�Aa�����۰O��[�ҡ߅�mX�ެpVa�MK���6V���
4;�
�Cd�y���P���4[u�%jp-��cf	�A>7�Wn뻎�;��b�{I��"�<.�N7d�r�4����i4Xܶ�n�lZ�z��7��\ʳ]ڑ��sNc�Ǻ���2�6������-)"�����4H�0Ι�u�w&�(2��kɺ��W���0�I�
X���.Ns����#���:������A�~Nө:�:�o�gD��GT�A�J��*N��wzG{nf����^�VRtt]q̸��*λ(�⋸���袲�+��u��w�(�ˣn�<�.+�u���%dQY�ag��u�YY�s�ɵeY�xu'A�\G\]��8]y�׶�����:�+.󳠳;;����#�(�O;����^^egW�IPpO���e�GW�<�~J8�q廲���Fu�C�P`H��T��5�20���Ȓ���]�H���x�p�4*;7�س��H�׶s�@��B���]�i��~���B�HP�GLLu���Œ�P�|I�zR��͵�.wF�v�ڧ|�Qd��6A9�77�=�ƙM���v��n�3�Q��\��z��?O��TD/J&d��Z�����(�H'���W���Pꛛ�������沩J"D�$�&��u#1؉zJ�ڇ78��� �H��B� ��T�r�d��>��>ᆁ�"��^O�
$̍�H'���Ί\��َ�[�|N��
$�P���R�T�a)(Q�y�v���jb�(��"uu�|q�/Q��Tw�ֹV�=ꔭ{d��-�uۆݾ�����G���F/�7u���&�;-uJc�Lql��2ҩ�_����Tj�n�Kx{*�vȩ	��8A����Iд}� �O7��M�j���?��׼�
��U���v���{(dj��3��BH�(%���8�CD���yN��r��Nw'[48������B��]���]�"Guۦ 8�}�k�5���=��X�'>8���/f�b��`�R�[a����>$�o&��]��A���t�DX��}��Z�(D���&�!�^�$�wn�i���*Te�ڱ����H'��Ղ|���BP�E].hv�}^���ѽ�펪An]��$�;�T��eR���بϼ�Õ�,�3.����C�dl|�,�@�yâ���h�r(�w������wpgl>*DeљR�T��&{F�0����t�����Y��e�T��)��=x�9�%g*�8w8����A�������'oNh�uw4ew���UⰉ�S����g�W��ۣCY���n�my�t��͒m`�;�4r�֯W[����	�#��e�su���o������z=�p�Y�#)i�p��g�r��˭\���<X�mɧ���U���َx�݅�2�"9�������n���6�3��c�Y:�$[��N֗�åS��]�NM�;��v�Yk]s��a{[z˦�p9'l׫"�nNݯԼ��]�i�JmZ�	Iw��/B�Q6�]��;�F��3<����P첀a���=g�� }�y�ě�V��l�PXUy�o���lr�����o���� ��l���T���wڧ�f�Se\�[QR�
��t�������K�2�euwF�H$۽�`oU
 ��U)B&A2��B�*�;�H�^z�wi�z��0'��!B��͏����t h����H�($�������u΅Ndf��8�<C��o-^�9��@n�T� ��.1������^�S�r+k�N瞗qp��=�b�Ӛ��W,,eꬵ��*�g����X�I
PC��]� �۴�D��p
�a�u!��ܻ����x��;�1"*mX��wܦ��������ȥ	�m�%�*#��bsѓ�h�c�� k5Mf��9��k���J��"+�+j�H���{�L�t��	�YH
���i(��ʃ�;;�4/���Z�ޣ`Y,a\���z�KM?��L���s��9�<g�;���ݪ	��4{�
���VK�k���v	'ǭ�HfM�Qwe;�o�j!��F6Tx��W�ZꚔf&A� �&�/���	�S�]�*�+[U/N$�}B�>$�E����v
��\�<�Q�5L�#	�2����z�յ�s�(���&ψm�R�9�xm��t���
H0$#)B{ʞר�o"��$����E�y��iЯI��'׃h�R
I
PB�zv���Kj�'��S S��� ��kt�J&�X� Y+:P�pxS�@��U�Q{Rh=6 �_��9^���Y����z������ՙ��^>��!�����9|��i��iǹIc�V:]ٸo�W]ҏ�������:���%^̯�s�tZm{��1f��4�,��+�_u����J�ꆨ Q^V }7@|9�!b^�"F���\fԑ4/2`D(B$J��_m��ԅ f/3�c2Ӱϣ����U ����%J�gY8��u0m�HHzIU�Z�U��p*�m�rd/�gt�U�*B�v��&o����D�I���^�N��~�I�ԅ1�Y>��k�>7�[w�Cù�	&��E	�\�`������ܸ��I$3��œ�|�* u=�����A��-�yF���D(!@��]�#�iz�	NK��T⩇Q`N_Vݒ�ԅC���D�HR.�3QzW��*�~wY�,�y�!Dط�Suw�c��GF�.���ޥc���e-��Ь=k|�=ra�ړ7�艀�En�8wt���̣��g�i{�;�������]�U��|����c�^.o2�S۲�ڡ@I�u;qQGI���77m��K�\oO�ƹMtv�I��[�+u�J�c(>�u��euQE.�3�׫��,��=�i@�$�&)�b�Z��� +��R5k+��9D���{�u�'ǇS��ƥ*8�1u�vH#_%K����_]a` )�5��
��pl�>#1*BFDՅ����@9�[RI��])�|�9υ����
��+Uʜ��E%����'�\��N��ݬ��h7ݔ�  ���T9{Z�N���8���9�B� n�QQd$����$�"�6� C.�%\׼�*��T�J�Q�n���s˰p�����%1wt�|�Yt��W��PJ����s*�V����)Z���B�r��V�i��Ɣ�-[�^^�����#D6���{b��Ӹ�Ձ�ar��{a1�su�i�|v�5��hܼ�y���s��<���7+���z���y�u�pn{l�7+ v�d�ӥf+7ctrα��������7���
j�:�׌�	7OU�?ߝ������8/>K]��ڣ���|�w.��E��e<;c�ru�ep�����]p:z���]s͆��Ɏ�Yk�X��ͮ��ns�`^x�PLU))��7SB�L�{=�%��"��ӻ��M���%I��|��΁�uÁw^�H6:�I$;�"@�$ʻ��l���Y&�fS�9����A#6v�$us˲|D�Ozo�gm��_,m{����!%�e�Eю��OSy~�1anld;'�7T��^s ��t$GW<��/:7T�Ib*�d��V���YW&�^96���8�X�
��/�W{���(_s�����3s=F۽3Z�5���9$��*�{m)LP=�����CĉcwS=x�Q!�n]�I<��P1���
v�X��I��=����I]%�/nKqVwcDX��c�p2���X��y�P��b�|�oQ�NV�X��|O��У�f����7�7�>�{�҄�(B���+����ޖ��4uDt`�3�q$��suX;�T+n4s�n��?8��P��[���l�z%�s�xO,J�Ԏ��3n��>��3˝�}f���V��X����z7D�H��B�'3����{W�7w�'.T�o`�	`L�*��OnՂ1��D�����ݭm��>�0+��R�D�W�J1�8k���9yյ����̓�ӱdH��W�$���3jwml�dM{GSݻ'ݏu)(�B��ȋ�vРO��9��RߜP��4?3^��%��(Gl<�%eu7�1Ti�&
��1��\:|���N8Kit穝��Of��u��tnlv�����$RIcRUW��\�X�=�(�H'�^@�c�V/�U��0���x�>��L��E�Ȼ�����kyX]]�ז���{vר;a�>ϟ�k�w���iY}��Ee����A��'�T�A���24.�yf��V����<�ͪ�źƨX�W >�6P�uy���]F�_S�ٖ7�D���a����g`5���Y�|�G�x��օ A<��II����	�2���n۰{Μ�v�w)
 �A#�� �z�s�B�;y��y������jM5@��2G>t�5I���b��Z��f�d��B����	��;��(�.w�x�1�x�$:�TD`��X�dܻ��07��p���n��_[��u��?_Ͽ��KlU���ܾT)���C�����'������ �o��	>����bL�RDJ�U�|MNDt�T�Y�m
� ��7�^�}ݎ��$1L]�L��tFu��/4��d���V(��$��۱dA��;��A����I����N�;�M�K��"�;-��ʹ�ξ{ӲO�%�zP$��RA �x��O>j�,]��7�W���Y�7��Ŵ}�ý����N������z�Ն�uf��S�Z4��="��Pc����=�`��'�fR�n�]{���b�7u bșU�j��Z���vvi��	��3�+���^�]�'���C��v�kk��~r��|�q ��d\���!Y;7'`��TY��UO^�ȗT������;m�LfL��s� �O<w~�>'�]z�s�[C7��랯@$��ۻ��j��	(E�n�{�!D������9�{�>�vmسϭz�z�z*u�=][U
n�,TLI����A{cj���>=�k�	 �ڥ�c��/�	��wd5�׫ټ0K�2�"��Ȱ��\J
/�8��֯n�%��I�,JY�QJ~D�[�qRr� �iKkv�޻��M�����M��u�| �TIP{��@�f��	!I�@�$�� �$����$�B��@�$��	!I�`IO�H@��B����$����$��IN�$ I*��$�H@�`$�	'�H@�`$�	'�H@��$�	'�$ I5H@���
�2�������������>������ =       ] � ���Q"��	R��J�!H��QB�@RJ���@     *�      @�  h�xDT�th�lU���$�r�ک��:�6�p�]i t�J�r�J> ;�  5C��
�XCn�o

�;�4z ��z��U��@t����
�|�����t��)l���B�  ���Xu�t���lڜڴ�m.f�� }޽mZ>��՘m�pvv`���Q%U> x  �^ӳV�����ph
@�s���!�%<9����@h��[��.ؐ:4$%x�@ =�h��E�al��[iw``@��5�� N����'���V�\�[��]e@(lb|     S�R���� �    ��L$�I@�� Ɉ��# O�*��(@�     ��4R�@       %<��M3T@ 4     Id�4��a�i�S�ښz��<Ԟ�i�zOu��&=�W��5����5�,�>h��>����-�UC�T���iJ��7@��s�Ň�ڟ�\z�A1�*�*J�*@E� Y (H��(`z�y����?�����m���D�B��l]�"$���O�>9]Xhh�u�珅�~�3��nk��tܙ�x�&*d�����=M�HS�d��ʹB6���r��<F�w��eh����]زK�7H�:����������u��'4X�(f����
���x\&q���9$�iP�R���#j�U���LV�o9��L�׉ׄd�Q�V���v�98�:�^q\���W:�z��g�}=�绻yy��N8╣ĭCޗ4Ѭޮ6(,��SѦ��#����q��,�Gy�ϖtrG�e�i����Q55�[�˰��X���k�H'���IK� Z]����{f��Nc���n�I_���Q���
�/ZC���[c�YI�;��睚�3�;^-9vn��vq����C�yMuk��+��s����e�����H�1�=#`���>ΚM�B1�Hk (�뼍�rC�ˉ��Ӈ;�C�-&	A$��h�^�D��;Q<Fk|P/�;;&�}�{/L�k둵��-)�7��ߋwU�x�`8���#(uV7t�>�؝��L���Zx\����Z3���w�Ok����M�����E&�Ч�����[��q����K�v[�g8:tͧ�����G:��/ ��Y���.�_���n��$">��gc�V����*��Bn.���4E���,6����b�v<)"V�u+��Ql�)g%�yt��ݗ)2odW�1��ש,�uF3��O`j>��$������Tk��W�*�u��淋��1�ۼ�[4�nlx���Yρ�t�]۬F�{�t����sj��N+��3N������tn3�[���{2�QÎ��9	��$�����vK��}�Yp5�7��\�(^hM_ݝ�`�ocw2����w���X?�Xu2̸�kX0j)�v#�O
3�7����`�:Q��nKcO�0�{_-�������81hLb��5��	�� \�d3A��,��%v�cÃ��`���vh��. �C�M��;Vq1��`c6ɐ=o����C�{P��5��Ēv��qS���u�u\K"X�[U��aW�v��p��`�f�j]JC)��&v��-q���z��P�Ӛ��`����8���qB�eh�y�z�Xk�<hHwkt���UI�p`��zϩ��^^չ$���趌j�otQ�F��sv6%�	VL�z�5TB��n��\�_�4�ۇ�ӹGK�fNΏ(��BYc�VN��ć����n����o7���B]�=��ٚ��܉��-tUߘ��\A�h�<��So�q��=���!����'����P@糛��"E95���&��@W�^.�2F�a��|s��O��nY�1T�����s -F<���t�jъb[�+yWx6^-�iD�f���g����sp-dNg^���Tue6��Gwsn ��~��{1�'�Q��'^�j�kl~����K���no%f��H�pW�mΚ�k{��0��x��9[ݥʳz���.'�s#<��h�k�FԞXf��/4��oί��F��,�=`��\�eɧ��δ,z,r]Q�A'POzp[���8仚T��̽֙u�����f�э�L���wr����5�g%F�D������P���37�.��`�ť���)��{"w���S�#�Z��͑G��C���kj���G+ޡqR�֘�4�)Ʀ[�(`�tٝy�C���Yw;
K�a]��p����^��M{�:���+���uѫMT�r���Qm��m��M�EuB�f��nj����pgk������ȳ�m��bYg)f��D�ۺ��=�"{[DA�U�xv3۲Ǹ4�+gZ燗��R���욺��Y�v�7�g������jɻ�(�!�����8�z��;�a�ۿ�Z�X��]ѝ����"9��RK;)��#�7��b��!�]�X�-m��s�.�A�ka���U��ظ!G�3r����QځZ��(]��[:p,� �8o)�û.Br�M�b%e��n���0�=g\q������u�F���G{�Tr��`/������#mkx�K9X7��.+BP:&VH-�Z�#��#Gٿ���p�7�.�7F��R ���e�+;��S�����wQ��#c�u�r��	KN�pfřY�q?�����ԙ
6oQ �� 1'���D0~���x274I��Up��m%��gK�o:E��!xT��)��`ǡh�|[vj!��7��T�z��y@Fv%���{�5��;�'�3����:�JW7T� �;v�݂ƙ�n�ܑ��̘H�) .p�B{pd'L��Dwi����Ɬ��J�n����rIe�,P�Q��4�t�K�(������P��3�854��yEgf�W:կO~�9U����ol]���R{;�F�9Be�S�q�1#�.���J�����U��M�A"���1�݉��"��JyC2�n�h�t�9�7��vw*�Lvf��=�FL*F���nA:jZ�v����� 0q�p�hCfN�zFF]���ov&!��Ǔ����~�������t]�{��Y�HYIrD�Z�	��à��q�Z7�؝����"�[(��:�F�<�td��B�^\��͋on0;T_��\�oa�v���g]����{.gm����&r�&ѸV���h�|1U�V{��=��fz}eN��
<I�I��=]�;'���ޢ�� ) H,����j(EZ��Ȩ�����"5V��H�$�T@��� ��2 �@j*"��%DQ
��  �DQ**���� ��2*H��$���
�" "
�� �(�J�/�����?0��z���]���
6����{ͬ"��:8m�.��>�<=�����Ľ[��3꾱���:��r�XNXt��}F?:3��Ì���3�V�흠�Ue����s59�8'�����XwrBh�����7��v9G)\Szh_�C��"Pq
���hR,�A����iج�MP�������Ob�q�o�wKz}O�7�i<w��+ܞ���Լ�譟t����ݹ���Ԗ5k\I,�˺!��)&���j�=}�{��\f�W�1n���s�B`��W��bP�oNV�rD�L)+�B���1�4���*3�����y�S�^KF��'�wtգ�n�)��UY�QaS@ܮmإi�_N����0p�?I�(z=�(�=~�jM�r�ޠ���ô�^�3`r���'Z�� �U��Qs�M�{}�j�S�8����I$s�a�V�Q��*@��Qd�����^X��s\�ݲ�Y6��X�;�v�N��?��=�pb�����@��Dr��&��}�b��e:�s��Zt����s�8�ݭ̔���ɘ+u.�;����e]	�?/o9��{�X�ߛ�#�]V��oA�0N�8�3�B����=��G��ͷ`��k�����{._��dYQi]�h�z��]]ݰ���Sv��:E�Rs��]�'C{�qC8�9P�x���CT\��a��/C�X�#%';u]k�&�֛�>���J��Eݶ�Wܗ�'c���pĶ�s7��0f�1����S���(�e�BVwC7��v>{�z�Rs�4���r�{�՗��>M~�[Z�^A�&���M.�e�w�c���cv��ޞ������&v?	ߥ�pH^������n<G�5��e�6��*����M�}PV��͠�sC��o�E����������,�z���c	<P�hvi�o X{�m-e`�dwU�A��+%���] �G�qx��wN����v7�i1
U(��qꞲ;|�7B�����N�]��3դS���ݠ�/�n{*]��"-����	c7,�E��J�����m	��I�Eq�aSmeAĲߟRt�|{۷܌��InS��A7F�wbg�7M��E�[�_a¥�l�`����\�b��z �E��Nlo����nA�6r�yB:C�vm��#:�f4Fn�er�ю��)��m�;X�V���K�S(:�7"W-�8[�T7(I����1_'Uw7lj1�4�u#dŧ�XnP���	��N��wV��`�j��>�-�>�YK4^`�;Q�iN1�v��Mv!o.g۳��,`�7t!�����f���P�w��U�V*�V�P�_nn�#K"��e��_<�^)��4{����\rl�r�^��C�^�}VN4r�9��_��ЉK��^Q�M��鬏B����f����.µR��4�X΃40�4�C��S/��Z �㎒5�u�'��,8=Rˏ'��=�S�l8�4{+���ܩ=���`��w$���q��Ɔ%�8c�qʤ���9)�.���3�GP!���c��+Z(�Ę��y�)2ا}������͆b$f��#�̡����W�.���^=����p�\0⏸����X/0\��mʣ�V��zO,V�b�.f��wv��F��ۻ#=�{�^����9�����M�/rb���!��x����ȸ:n�(7d����Oԅ}�P����U�+B.�o3�L��U�5�G���Ʃ���i�ys5u�\3e4���}���h2����.�[�F(���u��}x]�tM;z��3���!�����^�!��&ór<�7&y�-��^��/j� _�i_���{�+m��墽Т1,>/�uW�p���.�e���zf�읧�gl�ۻq���MNN�h�*I�j%<���~�Y�ϭ�rzRG�P�ܕ1(暱�hj�1�1z����k8��ow��7��9D�3��Wr=�t3ft�N_!-c%�	����a�S��Wۭ����_�;6��9�&Q��сu�>�L5swAP'"d���Ƴ�%\1a�|
nhlbu��o���J��E^�EE�AB4H�|�u��5�0g�������}YX���q�ݘ+cJ@���a3Bܨ�h2|O;<�v�l���^-��ͩ����x/��,��ťi�w޾�g�T%nh��z�`�S󵂵H?r��{���؁(w��d�s��������L�s����+�4ЏQղ�q3���oN��`����Ë,ˣxi��w0ǁ�P-Ľ�twj��0WOz�}䓓��ŏ;���@�#����O����se���:���u�Ϊ�gx�ǦF��N�q�-ʪ��b�߀�����<������&�<�{����`Q�����nd�����3P%�@�j�\�F���j�es���DWs��@䠅u��YǪ�vk#
V�Ȧ7ʤ����-�[繍��]AEAWb��t���͕���v��;��pv`i�-�b"�ig;Q��a��2�%�E�5X�yⲲTb������:�	
/;צ�%��r� �r����Y9���j=��gg&+����N�ZVD��S�U�e���kE屍ý���w-�L�]�/� b���]�ߺR_z�v���w�bn���u��>4�K��|��cW`I�1�tw:��>��;�f�ԗc�+Yw��.�bJZ��6>J@B��Z0�}��we�z
穃�Nr�d;���h��7��ܾs9��qN��&��ϐ�Fs�.����ծW�烈����a�����ɻ�U�%��
��JN��h��p�tgr%�Լ�~&��F���\�ݶ��Y_���hV5��8�DZN6������f�������	 ��C�R]	��x������~x��b�Ix݊맒6�u�{c7i��h&�-������יG���O3O7r��3Ǝ��8��\on�]]�Igm[M����S��iLle���[Y{c��3�Iω^���[�g���ni�^{t��-�-�9�-�x{k�Nɶ�w3�6�Ǻ��F<fF�[�ήڮz��`�m����"&x:$���.�ɳܼ��*�g$�<�a���9x|���ؙ�%�-����h�������8׎.۞���7;n���g�ٸ�i��t��V�<Σu���+Nևy�7..c�k��ζ�`Ʈӭ�̂pz�@���#�R��A��̱s���<\��s�&�1e�..-����8'��86ۗGZ����L�ʱ�⍤`��"�Z2[d� :�s����$�'=r��tt��w\m����ڻI����*trO=���%�uJ(�H��N�I��9�f�ѱ`�Y����J㢸Nq�<�N�Ϛx�k�[v֗-���tF]��$�]�H��3T�][�M5k���3�56x�&:�Ղ�ZMW���A�Z'Z^݆��G.Ce*�)�Du��GN��n�ოö�(���)�9w��y�.��pѻ;l�V�]�N�h�ʕ�kŴX������.�sz�Wn��Վ�Jk\�S��7���Kp��.1[4k�b݌\n�qk<{]��z�ݚܪ�k���u
g���s�l��������s�9ۮ|[�[�+8Nѥ�pXg�l�s!�\�lv��ݸp�r����l��ٺ���E����n�1z,�g�ԥu˶uk�un��0�o�ہ69�쥺�4�l<p[�2���:<v{'Z�e�I�4����^{v�G\��-�u��B�tMZ4�v�m�9����u�r�vkÊ�����&��,>���nx��}��y;�ѳΤ��J�a:�%�6ssd���	�=.�t�H�,�M�6�D7�"pC̷1�{q�/��d���S�۝�	���ڱ��D�JY�c��;fi��X7��;%�˽�;vɐ\q��/ktA�Cv�<��Æ�ī��GVN;a]����ފ��J����"�&Lx�P�Jmޜ��=�{�x�]��^�i���x��9�oz�T��m�F��g����Wj�.���ۚ�aɰ��5q���n��k����%������{f�t��z���M�n9}����>k�����R���l[f���Ӄt��cj�]D6�vE��%5M��v�Eϭ�Ym4M��Թ�&�%�����mz�v�N�jsv�k�4(m����nu�Q����l�Rx�٧k�r�=8�v�;<�r�6ݔ��ݬQ1�I�S4���v����,�8.x�n�m��d��ݑ£ky��U���G.5�ěZ.��6�:1�e���\�������V��t�G��T`y�ݻ���)<9:���.����N3�S�Q��o� x���Lv{e�k�n�p��<n
����9�-�l�R�v�cZ�+�\&�D�N�^��K�g�Ȇx:�U��MI�<��F�rnu�#GA���-�霝]t��c��9��z=ts�'u����G5���[��o����m���i��ssE	V9�띱<�b���&x�uʘ���.��:B�fM�Wv�1�<;^#��oS��ƕm��zr�F�\]��9�75�Z�[�ݓ'AiK������qp��b],#�ٌǗ]c;����zlv8G�
�qtjnT����O	s��l=oT�8&������`���Vƞ����63��sV�&T�[qq� ��1+��jޢمv���s�GOV��;�x霮�(��yk<�rOk<M�]Udj�`������ѝ��v��$������bH�k�����x8���mӖ;([ۇ��Gn�FK�l;Tb���ݝ��7gٻ�p���1Ús�z���b!�ͶW��m��P������]t��[ai�.��=r˳�,���p��s�j��m�ݮ����j����ߞ-�����9Rz^j��y^W�s*!=CP�t�/$H��1��^�f#ԯ:Y�$�D�g�{\c
�=��2�7U�L�"��"�Ir�Cه�,��s"��{� y�0��9�Q#ė:��b!G�T^��x��7\��fʢ��.�P���&t4�ș!үK���"�SH(�Y�mh�̏m.+�xS
��_|����ֳ�e�X��JQ��;�v�]�����=x97!k=�z6՛��Wo���o2k�q�W7s��=f��/�|A�=��s)�:���K��@�=��ҋ�xq������;�p)���O[nK���I��\۠r�p\\��yᠹ�֝�p���I�w�k�7n��pt�<A�l�N{3��lZ%�Kk��m��X�u��n�V����X!��yih�\��*�{X��0v�1n��v�eQ��r9�|�s�]��5��[�:�̙�2<7Nֵ��ε���a��!�@��n'����0��e�Ʈ�9+c��v]kg$݃��׽�]����'6��R�١�g.����2ڿ�c����%�fk�L8z�l�mԝ����m�{93�66Ԟd�;{���)�lm�L�"c��-F���e�l;g���9�cm����S��ԷN7m�2lB��f��vib�d�Ռ��vF-;�������������r��]؏q����������
u{q�J��5-�A�&I�A�Ŕ��9X�*��u��������XI����j�J�˿�!��7��9�x�d�FTl��_B%�\�^깙BR��o��96���h�����$��0"�%���K�<���g��"���3%i��ő�Q���Z��n
���W�j��OMܝ�*�(��mu��]w��#|�?w0���.�UI�+ٺ
uy~l��>�ќ��$���H2&Obf���Um� ��'�a���t\W��r��St�J�A[=��vg�$��O�鯝�{��k�(���EmqJ)]�����9��*�m��}�A�}N���?H����T���}+l�_�9�>��tC}��(a�Dв;j2bd��񴢝�,�n���RI��K��6�n��N$�wϼ�/�h)�e�ze�ME�����)�􌍇��`�&G��F�1��D��L���|�%FŃ��ۊ�m��{=<��v2�׾`���+w[t_X�a��/C��> ���,"����/��?dJ�XS_�`�_��װ����D<�M#���Qo|rg/����$�+q�^���$�b��}�~~�}XOo��(%E���>�N�/�dNV���}���;�^���|�[Qm�ڔM�k�u��}���P���hY����u��&A��L��St��&��ˌ��L�����oG=d�����A��2g_����mvz$�XPfشIq?��[�uA���2�4�UY��R�w��9|T@^!d�l���{�S7�th�tV�%��`oM��K|�vI�qde- �2���:X�/�nݜ��gVm���u7����5i�9���^\��õѝ۬� tX:;c.�ں��{�z|[�����Fm5<ܹ�j�+`W��@�fu8]yk5�?�F��u[l2A�O������&aq��`�v6?w6GfR�Y���S�c�Y##Q�g�H �A��4�Y!���k��a������*���Ku�e/�!��O�e��s��
5GD���!�,��+t�f/Gj�k͂s[$�5}.���=��h)����h��r�IrK׹>��U���ᛰ�T�#��o�����$�&��#�B=��a���6�j	��o5�W���~�J�+�&n�*�d�l�o<���r ��1k��Ӹ.I��Ȅ�{䔯�Z����Z�جbbv��+]o��as�?X6��5���c��2dl��F���d��bE��\�#�S�L��
u}���	�69�u�U{����(�W/������q��n%U��<��:58=h��&��00N?�0���^��}�%m+�־ȕ!gb���'5��CQd������\�Y@V�>#e��y�E[�͵{�y�v���=�cat��*f�k;�`��r	��a��מ��j��D�Xd�f�^\�H=���-�M:ʋ�WU�c���A���YA ��;�X��+�b.c�G��y�UV��a�ٽu}Y����c־�Bt8ׅ1b4,��#��>H^x$lծ��G����1���}���6�)���hn����>��:͆W��k>�2dl����5���[���`�r&A9���W��}��#��;���ۖ	�����+�j��&�e�w�N��i�o�*Gbd~��0wn�xd��1���D�����׶Ly�b�Ѷ=)u�q3Y�����?gН��ly�B��^Jk�9�N3mt\��EPv���ӯ�r�V�k&4�rg�8�su�%\=�{
`Q�8���[y�mX�94�{tӸ�������)�L���[�����'��L�i�I�§�x6I�L+=
�K��ت��$�L�N�@���I���:��H5$�N��� �#ݾ���ܱ	4�dN_w,���b�-b#U^5��zXuT�ifhM�"wo�ң�E�@�q�bR����B�ؼ��C����r�I5l0�C�I�=�V�Genio���_�hY�<��T�-՛ذ�׃m���!7����kW��t�k�}�������O�>|�M����d��꿌���� ��:4�rֳ3��W���$���P�x��${�g�3Onn��տ�XZ��� ��;�U�����W�sd�ژ �`�םX�����g�N��i?j�f�dMF��� ��rA{��I�|�����A�����������,���9�ʑ�i㜮0Ž���wq�.{������K�S��]�;���`��gf�f�1�W'�F��r��꫸>dZn9�Jg�����Z8s�+\c7���η�V���Mf����R�r]b��#GU��̳��#�p݌a�=K�M\➾�OL�|{�sz�X9�]��_lͻ:�7ܖ��=�U.�o{z��V㗷S�IӜ')��
��w����ŉ���]�QC���G׶u=��s��H���
�B����O��v9�#�/E1���:���tكy~��L����6����'�Aҙ�s�Ԯ�\�j{FC:�Z�qK1Q��+ə�Ld�&�R��ߣ�
3ļ���.�掑]�djtm�cC�D��B�����"g��A9I%QA���EC<J���mq����<�u�^NG-*"X2ɘUD^Qh���HQS[�.s��;�}�����]������:X%�W�J{��:~3r�m��_��y/��CSx=���o�|>�`o;a���<�E��&���m@9c@9o{��0��2}�D��;Tqi���t5���hW�mz(�L���!�$wX���I:̨��jd���VA�2Ore�C�I���U���w[f���b�T<+���-ޣ�� Ś�����1��Y1��g�j��N���dQl�i��$���z�������(���BU�I(���Z�[�M�
�-xH7��}�r���t�OZa{w��Y��&�S�eb�	�L���`�|my���Ui���VI���XV��sezdI:���c�� ș`�@��2������ �Z�{�űz��`�����1���W�	k/�]����*�γ��3�����jk*�>�+!�/����ۣaŭzw�d�G#�o�I���\��S�b�sz牟��w<�ƕ-�軋��t�M;���ݻ\�l89��qC� �~��_���J�־������u	=��wF�t,sa��mky������d���l���א4�hi��(��uVsI=ɂ�l�(pUT+��v��\mw���{9��F�}���.�|!�}���t{��#z#��\��(�*���#+`��Z�s���]ן�h��x4$ldl����ӥ�V���p#פyY�N����ݖi��w��t*D,��u~_f��	����o�r��!)bT9���a�ٟ�k�Aq�A'9�����Y��$���'5�-����2��`UU��o�j�|3ޏa5�޵߼-m>�.��`�$�[Kd�Z�+�B�ds���u��y��}LqI���fF��`�=hwYo፜�2���l��P��у'��$���Y^4de�,�˪������n˩u�}��O�����<&��qKV˰�הE���Y ȭ�7ۀ��SwCN�>/�$���<U���;�;���o9����)XC�EH�W��t׳˪[|���� �� �rh0y}ܴ��zhI�8�]�mzy�n� �6H1�cg2� k1���{ �����F�d��<��M:V%w���Ey�EZ`����ٿ{��Gߵ3����U�3��*�����o����	��	���*��֐~�#����\��@f��4��.�X����8(��3���� iօըx�50j�r~͸��Vq����r�����H�lOr6Mٕ��8$����$�r��UwW��硼�Zda�Ojg���B�����VǞxAN��R����nwL�D,�L���`����q�Ṳ�վ�]�spa�W*^T6��������7H'�c�Ԓ>���*� �l��� j�wqy{��q���#�Ku�۞׮x��uu�2;��9wY�m��#���c��k:����I]q�
��-�3��Z�r�d���Oj��_a�Fv�4�������I�/���ګz���hy�c${[$]�])� �v6	�~�Г�qKv��sQ�$^�Ւ
�ޯqSI���n	��=t֨4�d�hW:�V�YjU�~!,c�r���^T�~~�6��6�\�'ɷ�b���N�T9�#�{����W��vw1_�n��p�a��|��>�i�r;����}��w�!�r/��N�h}�\�ʼ���Y���M�2	��-����96��j��ۤ�[����٨&����۫.{t$�ZI&swvZ��Ma)�q	���k�e���D���V�"u�BKJ���y�<������}�e<�l�{2��E:V=KA���,�BfD1�|^%�c����\��D=8���aߣ�Jנ|�}�����g�[5&��Y�ڷ�����<3������x�|4��{P�n��:?8sE�N�gR���T��&H3R�^�q�267���Bװ^��BE�$�*	�����*[{3��>�A��A���,���B���i����5�j�A&��sPg���v�yႝ+��2!��d�w[�u���UB��n�����$��3����u���+Z���y7��YjΜtJ��?�������T���Ӭ�_���_���0Ol�A����#��_��寭,-R[[��(���j��;�����N�ͧ��m��>7sf��<Є{��aw������1�z�d�0�ٳ��ʋNՆ�S��� ��2';їӾ܍�;�~���:X%zP�a�H������_(�%�����[����V:?���H�����~tu��W���W.b�w��;��Kv�`����x*�K�]�������e���z�l�ʥ]�������0���N�*�u�Ӛ��]
�ڧ�nS3�{��M˥Q����G_m�΋z,�k��5�_tw��D\ݒ�P�.�Z�	ߛ��EE�~��4^V�w�}����u-m����}5Nٗ�&ů���Ŝq��]ʑx��l�ڱ�w��_5�>>k��!�N�ֆ	7��X�b��vK�lk�{px���������v.d>�������f�V�?1�Րa����;Ǆ>�׍��EUU*��$#V�]F�F瑎�Y���f��D^C$*j̸�u&aG��P�3��&���p�<N�R�=A��{J3�j37Wg����i��܊������V��v\l/Y��5�\5����9��g(�c+ڹSghӹ��Uȕ����HT�$L7�6��O�o��#_�i��]���Z�<S�t�N&�k�\]��	Ƀ�x�[yǱn�;7\nͼ�uqQ�97<豌�p;��͒+t��P�F独U�U$ݸ�w׋��n�u�dsq���f�e����gk0�מ��w:!N��=�&vBP{0�������=<`���3�m�t�fNu��z�\�3�K��cn3Ħ�&��r]xxخ\&��[�u����W�cFץ��M�a]�xӶ׃f.��q��x�;��<����:4�w=C]-����e�m�e�ݬ�z˞:.S�wu�E��U��r4��E��U�^�tqΎ:��6Ln�Ci���c��#e�<�p���ld�۱ˍx����� 9�)��\/\�3p�6[5�;]����[ٶc�^�۴{o#��<z����|c��z���{={ �[��.�{���x,�׳A����c��c���H#�[�픊 
|+k��\|��r'XeՎ*����mL�e<�u�X�M__�����Z����Hr-!N�r����V	��UA���m��fD��"��5ez�"�^8�"kw��H>�d�}��ZQ�:��({��{���1�=�}O��4]w��t�uk�m��+�Mk��y�z\����b�VQ�*��A[e�
�.o�}���hmk��@��F�⪋� Ț���f�f����XH���
����:����.�1�uK�?����u��$�o͒}�l��1��V��_b[�̨�	4?���騷X�������i�y	��kF��Oʸ-�LKC�[���dl�D�)k�v�'J�D�C��Ҏ��v�"�-��|�YMy恦���l�jt+��3�i{N�T.[duċ�l�-Os��թ=�ť��<[u��}^_qϲ����m-T�����;T�=�ڳ������q��kT�|>��k��_�y���j�>�;o䩒;Pw@y���r�ǁ���*��m��M7�Iu�)�}�7U�7U�W
�VZ����]<��>���Mo��;���F�>��];�-3%]u���3Pg�U�1ڿ�K�b5CԾ�~_{k�V�I�F�׻�[w���|��O�:0{ڻ�}�?�;=p�ܣ�,3���Uݷo��z��=�Þ�{�_��ճ�	�[Q�-��L���V�����p^��I�M���B�2�G-rJ�e�o=хב����m=�^��o2,kz�SڴY���,�Zi�hA�L�n�]�<����B��O�z]�]�A�y{u%T:�R����/��j�qt�^��X��~@���X�C	�����.�bY��s�<�u��{mƸא}�a#(��o9����}���QBX��ln&���֎��fP�ĉ���,�x����w��!&��=��^�D�-��Y<Ze^e�.y;`�2�U�S`����\�6��B�\C�;�'�m���&��m���=�>ڔ
�	��y�ki�c�d`޺�C�b5���y�ESЀ�L��p)��d_M^{4�t�VMU�W��@l`�Y�5%U�]�^�����H��w��Ƃ�Emn&)P�ݮȊ��s�R���䇻�N!%��`�S~��^q�0�|i]��JώE��L�R�틡��������q����_�x�tfK@fs�ݯ�������~��;�����0Rˆ��r��$�5�BD$�[W��3���a�T�7Z
�p`�]V�tIU{m�v������o����)�[��wt_��_|����.bOi�9�y���ӐA�k���S�<��fPf����;�>��������!�}����v���rݢ�Cu�p:*��}ء�]���|>����c��HVZ�WW��qrLi�����%��9��$�� �vD�j��k(�@/z���w��K� ����j_�\&�ƩS�-$3�!h$�wk��M�5W�MZ�|�[t�_t��S�_��g��8	h�!|R����-���c�l��m�wݸg��D�P����	�Ȗ��T����w�%Տ�}ɮ������~I�=����[�
)؞"�����]r�־ +t����x��������)�&3H���4 oT8�Z���n��oRK�v�ku�--��O��|�&��bDEީDHgv�u&��m�P�	 ct�g��z���l�s�H�y��[���� �� ��H��(�z�s���w�MT���P����"H'V���M0uH���P؂B��έj�P7z�=��])x$`�*Z)��KA$G��V�Ư�K@��m�[\'E�n��P������7Ց,E$:�-�T6�s�w޻ͻ��o[ޛՃ���y(�:ѨV�G�2�_P�������MTQ�	0�A���,��q󈞸n=qr6۬��ֽY�v�����^%�᳓���KL;v-�+��n��gxpqm�+�:u��Yy�zFvK]�p�늎*[�}���_����|��"�i!�I�XKE%c���L7�:� �W�h���W��� �P����]R�%c}��/PN_�r^�{`L��(-y�-��룭^�Ё��.������K� ��[�9��9�i �]Y��R7(LEz�'{ѻZ��5�PZ"�tZ)�g�`HE!��KDHCy�~�b�.�����֖�-��T���������[읗��~�,D\RA!�Y���Z�_*j�h$��t6"����KZ�0m�A�\�3�*�g�h�Y�<�������'���s][�9؀'�<uFH��i�C|�A;��v�V�)m�����M��1�WPCz�k��7딡h$��Rv��/V�����_8��E�Qȉ ��D�R�(w��u�N�U�m�7���� :�+����3<Ʒ֔�o�D��(@�(��+���v�N�L�ebɮ¦��}�wkU�@��;���#b"oT	-JHkT�$��R�l�M��D����E9����	��D�)�r���Ku�]�����y��7եZ� �t��!�Qh$�B	�����ޯ�2h�pW�HӦش	�l�#�ړD�E�N�'<ﲛ�N=(�u�Xv�rL��6-ږ��P/�lU�c�A�^����ݕ{\�ߺ+�����,_k;���*�Y�x䜸?V��i��ra������ �o��;�ڹ�� \/��z�}�޳٠�J���[��Skvv�D�jCO���L\�T}&�y��\�7{�^��Q��c�A�M���h��[7{c+%���ݛE�˱|���Z]}"lW�9*�eKd�]�1�S���e�]Rj^`0p�٬�]{m�0ނmoC��P��هEcn�,n���}�o�i~Yv��U�O�	�YWb1+�T��M�8։==�e�}l�3SD1Qxo>�'6EV�u�]U.���s{G���<�{B.�/"�Xպy�8s-�'���>�W���)\)��:HJ"�SV����}먔3���k[�q���kh�<�{�a��&�<2����Ĵ�T�!kT����5�+��H���A'/͓W��7Alw�ԐC�R6���	b*ot�;��g)z �ߝn^�{`L��b$ �0N��o�"Wt���:�[@�)ڶ�w�����E��.��C��7��;�{��Pv�I�TY�H�5݄�S���;�2� _t;�f�j���Ah�������9Օm�@X�H$�����s�񰮩5��������w;�S��&b;�Z+���)[�z��_ �}u,��H�7E��)'7H�`;�!|ߪƵY�Uu�C��9�6	�&m�iy�-_��|�}P�`��tM�_�A�) �y�qZ�][�^�k4�u�\A(��~�_|��n���C��g����^�@���$R@7�-u�D�q�߻�(�T�ryH�nuR������9��r�,A&ya,E${�]Z^�Z�	޸j֫�w��"�tY�B"g2���3/��A֩lA;�{&����1�}�"a��h��w�R�C��;�nn�1]�,W3�E��ș�~R���U�7�D����7� �v�o6�/�ۘ;��:����k���?��| �����ƙ9��ΰ眻Gq뛱]�����5��W��Y�:�l��&�Ō��{\��Ŷ�-��%x̕A�]����-ƻQ�ϊ�B�X�k�p��]lݤo����}�_�<A�t��f��E&{���[X��GzG9�:�H$���ٿ}j�V����к"��;+& ��b�h�|�8������������D3��I�bb��D�?}��_|����6�%O�3��������.��Uh8*��1��Ř���7����2�$ˌ��K�5�����y��BbF��;ϳ��������=W��H�tp�k��h�*w?��  ���BE�"_���I��)LF��{
�}��i�j���pm ��R���ڬ~�2MxQBnmf�̘����t.q�<��
�[%?_���>�R���dn����W��[��@��4'֜��_G��&�����s�q���}<�׮���iZe�}��Q�� �;��ھ��n�N���wU��b�K�6�a��*�#U��16��[�߯{;��8{�
I]���LQR�"��~���o*��WW;v,Y�k�+�xU)����� �r��D����[������)���WvW������ ��%f�Ҏ{A~ԽMe�#}�y���z�q'g���,����g���������]Ty�/��-���f���s�Z�%�Čt��`k����G��ex��c��3��W)�u"s���O��bOx�|G�/}f$m??fm0�W3�4��97Dߟ=-ot��:�DH���j=��K��οk�x��݉t���mݽ��x���?}�F{38w'��%��w�"�GU����)��K�R}�p�4dY�z��۶㙢��{1On�c�n����C<l�ח�����Gdu�-�Ż���v�dܽ���6ۥi���T8�ҹK�=���z~K����'8>��BW��>�������Wa�v��[0��4�j�V��4��<������.��[���z�7�ѤL�.�toE\QWTtB�:Ԕ����o۾'�k݋�r1���:�g=e�u֊���W�w;���~�"�aTS���t+^&�1�X�7���������j��������j���a�O�ӱ����V�-�{��}�Z�n1����S���R�o��3{��<ɖ$]�[��o��ߏH�������F'bb����n��z�w�^�:|�����k��_���ٞ~���<���3UR�}�}��r�Ҿ�_�'�j�*��_:�齱5_��K�� ��'�g�1��3�y�W3�,U �?��[��V/��}��
������m�oF�XZ��r*����T�Q����>JO5|=�ep���:��`-��Y���lCuyy�e�{W���]~����W�H��u�U�����N�]h��`*��0��U�i���aN�|u;Y����~���~���~1��j���}�"�^��^���N�e�*����Q�,�@�[�w�y�rQ}ۭ���2���:*�ɦ�������Cj�=�}���Oz�H;��c����/����}l�'����F�k2 ͓��^��sV�x-���N��u��e��:���;�Kyڳ:�K8�{R�^킸�M�d�%�s������h�s�0YwS����vr�\gdDX��Yt��n��Փ.������;�LwT�����&d0bS �2�n*�:�%f�R�`A�oU��Pfn[�"K.(z���j�X�\�v�0�#��D�[�x���u���~�6h����/���f�ޖ�_��;F�Í����u��k.5K�f�� �_<��Zy������+2����8�����k��|�:�f^d�x�Ns=XoF�BA	�fS�D�ʜ���I"w����?���H��jYQ3}(%ʨ���BA5�Ծ���H}������xxFj{6s�|�l+��F�9U�Un�܉-ӥ�����f�.A�Ġ�L|90By�J�h�D�)���)����%�+Wpq�y8��D���i��y��ר�K׭�_{۵��S��DԏY���(�[��rz5v�7�g̫{�.����a<$^�x���.eI�V��^'��k���Rჭh3�8cU�h"��,A���η�I#�\�-�C/j�d�NӃ;�N7�0���'Im��\�(�h���^ruGV۝�F.�stU=�v��q�<���9Omq�KhOv!dGzƨ���!��7e���㑗���n��j���V�k���5vۊ�X7n{��<�H�;y��X�
3��7n�9�:��f�;��~[i۳1��%n{I�s�'^a��捳հ�
�q1;q�ܦ ��rIᷬv��Ѽ�봒�wc�� �u�c�o����v�Vy�]Ŷn�ϤspZ�r�=�έ�sÃ�2���]�������rv.�������'��7vɶ���lV�8�W��1Jz��s�II&c�Kt��<�4�ż�c����î��$˶<�;�h٢vB7��w{���g\4�1qZ��[r��d�f�s�N����iî�<����=���"�8ۮ��7=H�3�߇���G�ں��[ݱ��ڸɕ,���t�"��M����A`��}}����}?�s��T���V����+u�2L��U� պ
�G�E�i⽫՞�?y}��O��Wv�RT�k</uX�Н�Wq/������˹I����]�꾠�,j�#�5Qc�UKn�N�o4{��7�K���S�<W��P2����+v�]<��R�K$�'E4�J������~�1ܒ��[T{���\��
����y��W�b�δ$S;�I�w��>}��~�w/��S&�����Tk���ۨ����>�>Ay�����5��o2��MA.{4Zr���}ܻ5�<<��UQԒ����f��8�ׇ�ٻ�(>��r�Ϡ�P������/��_{�+`Z*���η�|�s����W`��I�M���[�cv-?sD׶xe
B��� �RKJ�S͓ķ^�]z�E�e�G֘�<��*�G~��/�~�7>��/Ҫ9r<�^
�Y\����eW}�{�
u�?} ��'�L�^�W��9���^�ny��}�c�|���\��m.J.�������x�-�������x���}����}met*����<g��u����u��{�MDn��}Wȷ]���:	��b�t_��W]�z�u�ߺ�dw���Y������ss�a�}�@_�����;Eז
��=�Q�P��%g��
��9K���0��P�Oz�Y�	�����OZ��� WK�QuT��/������;�}�u{k�[�l�6�z�٩1n�{ˠ�wT���̹$�!`vN[.�ɝGm����rck�p�YԷ���[���pJ����Z��{�y��9�{Ղ	��{���܌s'�G����r��<���F��9����S�����>�((��Vl����45��4�+�[Sv��Q�{��▬H����
�Z��(��e�߽�aw=s8k�����e����V��oۗS6U�y�<3z��ݲ�,Mŉ��y�|g�o�~������96���{�W.ӽ|�u��Ӯ>�󶗱{ܫw-׉�5׃�s��+i�f(i����ɷilܶ���L�rTl����%����F�[x>��GS�?�mͥ�F��e�|j�����* {�?L)��On��2q�;�}�Zb�]b�^7��bj��������׿3�վ�Ի��w��O�lE�se��[�]�Y;{���mVGꎈV�ZnZ;lﱿWo9|��zg11f�=�u�=-���>?�8b�p���i��?,�e}܅�@����k�ʭݞ�A�|��~a�xdUg���n��,�ym�۷Ǥ���~�0:SFEț-~���w��������R�]@���L�U:-���-Ӟ�@LU�|��I�V擔j�h��rK�����׸`�R�������)��IՎd�卋�ջ;��1w��j��¢�v�K:$[.>��e����>�Y�tL��R�����;���*lݐ(�+ARP�� �pU��,���v8h�i^2mó��\<t�����l���V��q���˶���\�d�w r�mv��<�[s2��z�ְN��ޟ��)��r�bg:�z�3��7S\p��<�FRB~��<IlAW��t��9��rb��{�c���P�[-,~V�u<�?�vixr��d�����.]l��3V�{.&��}}��5�Qv�8/�>@�#�q^/s��g���>���2�Y��'�Ek�u.�4��Tqn_�˿}<��LK�~q���[�Ҵtw�.�z�����x��[|�>��n�Ö}'7z�ū�έbtYE�>^w��]��TE2�;Y(+`�+v�{=�a{��~��}�,�<���j�/��rw�K>�2R0:R}��`+^���W��������͑`3��#iVqހ�{�i��.I����g���QO���,����4��};.�Z��d��a�|L��2W0}G�i��b����뗚O
��=ȸ;�I����K�v��9_�/{���w�N�q�tu�WeH���9�[X�*��@����d�G2�����ID�p�pc;R��݇���釸��"r3�{N�Bg��-�39��T�	�fe�/���5ՙ��1ᇦ���:�{q9�Z�y�#��?o��? �����\�A
O�����;��������|���o.��3])!���c5:o���P?-�����=+z���DL9��BTU���9��6njx]P*���@�fyAW̵�B<��`�Ts�
����(�W�W++�����.����q�é1B�z�U�W�2� ����r�3��TAEU�=U0�ʢ����k�E�Q��nVd�5.����b^_=g��O�?
��y�t���ꥭ|����Ʒ�w����UH��+߹��@G=G-=�?v=뗚E>�&'l��+j��`��V��}�TgR��"�,�{�S��M���. �}H��j=�{[*�����O{��y��;T���|�칵�
fL\2�l����w��_� s;�-���gٯ��h�@K�_$��<�}�Q���e@�ݥ��(��3U��15^�:����<���;}B߷&-\�J��}�֔uNӋ�^���_wq���3�m�P*P��]��k�-�;R����ܤ�c�=���^�m՛��T��~ �m�/|�XM-�It��"�ϓu����%¼a�>uL�b�^ޭ`uN�U�#m���������Hh6���s��`ɸ�u�z�\�TH;Zߢ)�l��߽�0�?��Bb�]���An��j�g�x�w��~�.�#�)���A����c��r_zҎ����'2q�fa����n�4j��}�yf|�y��R XH��Z18"�d-���}E�o&mu�9A��q�����z��4�3�O�|����b�n��3E� ܼ�{^��S���rj����j�������f!��)�v;P�3����E�uǨ��>���{��;v����^m�AU
��G��5k�_s=Gz�\�]�+��ƪ������򄛹T3Wِ��lL��W�E/d�:���
���5�^
f�����f&���w�=ډ��w���~���ߐ���j��_�;ܲ#y�����ˋT��%)�)����^��{�r��P�T��u:�-B����g�}�}ro5Ҕ,\��f���}�vؘ*,�;��þ&�T~Y�p��ḏ�|�uuЯ�}��p�^���2�����I�i��WثTw*�twczq��������o�MU~����-��8�|�?��@�+R)�L���@�X�d���G�}�ś�k�5����=A_���\��{r}�_w/�=�+G��3Z���=��S���<*��t�2���z�Ezof����[���s�mmZ�}��b��{��o4�xǙ��[���K�ϫ��O���.��૳<��]IТ+d�<�F�����+��{c��:p����K�>�y�.�^v��u��r��]���Z���k�p��%��͙��'J:!Z�M�Q����w�З��E��\�EG=ҕNy���)GӬ������z5�X*%�ʾ�_f����u�hy�q�A~��!(π����<o=b4r%�>�'�_{k5ݑM}U��;��H�p�2��\�}__O�Qwr�.�!"�X����P�>tUM����lt�w��S��J�.������;�W�-��:��3#I�����ևW��N՚☀�W0m�����k�Ra���h�]ׇ�S�)���b�dv:���6�UYn�������Y���g�d���-Ӛ��̹h^���G��Q5U�־�,�1�{'�7ѱ�����Y�t^׽ݯV잉r鹸y��_��˻�����=w�o�#yc�M/�mpuq�\��Tku^��L�Q�R�E��	�����|r��ϫȾ\'�!�==Kr̕+���j�Ļ�v+ĳ���n�gZ��NP�}9,�X���'�Vs���>���z(YUWa�>�dn�j�p�tM��U0wDp��G��@�:��}1\��g*/�d��P�0eDeE;T�p����<�����Z}����f�ϯ�v��·�&C�}�BF�ϾkY�i~���e�|W�������m�hm%����^�gb�),�m9k���,\;޷���H5���S˟s�H����orFMc��V�ȳ���X��Ǥ�5}��/���w(�|�����+Mv��:>P�w�Q�ܭ{@.{<�z��{�R	d'��r�g��`I�9w����B�1�Ϟަ�#.G�ܻsk���$�j5�p��VMo:Z�2�5_ά�3��
�ac��o�k����l����^黻�rE.�7�.^�n��{ �Rxt��(<�xq��sJɴf�sel�
���]Mz*Cۚ�%~p�XֽB���N��;@�G�孲��]��������2�r%[�\z5d����Ӛ�͒j��L?��T��)D��#�"�}]��_�Wm"u�0#�K]B�Y.M�XYD�"��nyU�}u�iE�E^QD�<�]k8�b�Y�5���"��ES�J>I��r��*��a,J��j|�*<���'׮�垁�D�����zs�d�^B�맹�y�*};|�Pΰ�͛$�ܻ��������.;T�ɹ��[��j�M�Ńv�nKbTzۈ�5R�[�|��ң���s��R��y�m�z�X���=�s�u�$m�\'gP��֘�����Վy��]]�.��c��H"�98y�\�V�LG^­���A耜��l���c�e��Ro�d󗸐�63�sOR�,n^vZ��߿�v��	��!ɌZ�	���'Y[����-O�|u�7���oN6��|n��ل�U����>��U,��i�wl�d�6����;"6�nf3=�<:zr�n:y�lB\�)u��r���.QG���gh�d�8^��v�5�=+�zV�\ROc[��
yg��v#��d&gy�(z�t��d��-5m�O:�ul��=^�q�v��V8��v�H��tۑ�j�|�\�,����εn8{u�qqX3������Y�kE�z��;d��15iu�)��3�ҽ�
���5���PH��%�6�\Ϯ�<J�'d+j�k�����;�O��73S]�4[�ϻ�^�z˫�_y�]���1�\�#�"5�Ծ�½���{�y}�����ޞY��R�.s~Pz�n�J���!_]���#�m��0h:4�L@�*��9ctv�;��;{�QkwB�vgq˲晋�̞��
5�k:ϑ�u��ur�nb����߾��߈ݵ^�tj��,��'��X�ظە�)�s��e�K�f�9l�`_j��[���M.�W�EK۩m���2�=��k�3;.O<�����j�k;ν���ߧ�|*^֎��{2�F�w�F9:�\FG�����y��y~�B~K�^���5���ʈ���Y�X��d!O"��|�q���ҕ�4Q����bǚG���7����T����c��X��߯�n��|���ނy|�A�Kz��j��h�;[��}_OV��U��nLµ}�|/�Z�<G���]��k&��ޟ��>�M)�;bR���W�|˰�*�篇��F���+7m'f36:�|�w�F��j��-�׾5��{ͮ��^ �t�p�ߍ�r-��k�'�����D�GY�܏���פ��l�1g+oS�f�q�~>��J�bd����[A��2M��_��q�>�_��r�-u���ћ�<�Oo0�k���ʭ�j����{C�]��7F�a��g�w���rP[���"��vл(��t��ڸȶ�nj�u�.�����h���]�qu�����[qi�v�:�l/{�,�?>Y����ь���'u�J��氍�R�*���"F���7u]�M-��@��Whd_3��;�A20�?H�%y�"�U���;���2&H$͔%��aK�<�]�q�鎇R�OǱ29̓{>s��b���V��(�uV{�����#�2	�!<N�u"�o��ϝ*X#C���=}����6P�V4���L'�u=�ү۶��y+��y�2&AkR�z�X(T��l�\�%�wE>�W�$M^Y
��A�ݽ�ED� ��$������u�E��xA|�M�I�_=�#�ؤ�T�l��K=>[M�_����L�ޯH�A���y�a��W��٘��]��Y s�#50C\�u�~�|�R�>�$ߓ!�l�k_��_�����o���,���R�}�c�;����
�j4/��a1�U&A?��.)CL�ž��UV`7g�?n&g/���r`���~����*��vA	�H��;Ua�g}Dw�#�f�øe[lܙ/���k/�A�z�>c\D!��'��L�AO��阃bd�/UZ�ٜD�� � Þ�Ε,�q�ͱ����$��2$��YS=8�N�4K��Sn��@i:W�Cp���9��I�L�`��A6�93��o~����KEjdvXӌ*�XU\/{��9n+����_2}���l�Y�s�ux�"�U�������S$��ODn���"<�^v����n�̋�z �A�Tp�R��0i��v��������V�)ӥb5�N~Ֆ:�0h�������/��zR��_o���F?(��h�>�8|9\���g-���mА ��:��t��X7O�[����4V�z�U�>��GF���ż�M����&�^�I[3�f;t�<���ϰ��t�d��k��EY��Q�i�%R���n������`���y�w����Ǿ%�3翶뽀��x��^�궴�=i�ND����
���꡾l����ʶ�{>�����!��:�fMg�"���'m}����x��v�{���^0M�?�L��$�F���&���(�ژ�����V�tM:�:*�K~d.&I�&rEs`wA�"`����h[������*Q��풺�87�����x��ʹ+s����Տ}��H�|č��x�����
��^��#ڙ���{~�z�$�y��������G�^�I}���sJ���H`{�F3Y��2&7��i���g�7�{Mֻ�S�buZ
���ڵ�J�n��O���͟k'��b�k`���*{�U:X#Zd߯76,�D�:0� �?��%�D!�W�j&H5��P�[��C<�}���տ�[�r�?���I���,Ҏa�����Wb�J^�٣hȭ?� W$��i���ͼ����A{��de���bے>��ڦ�8Kラ�`�Ii˃�ۖ�e	0�i�݇/-o��B��S�=���KnUO���g)��]�+b���pd7<�xC.����v�㺹\z���wJ�1�<��&N�]�=i>�f���b���}�ۃ��C0�GIVB�39�����M�T	�c�YH.�X��<;�,��ܡӸ��y۰,�C{q�Q雇��1g(2��d]Z*�0�d�7sk�-���H"	�Dx���G�$�Iӫ�//l/=���Ux�$��'(�'(��2((�B� �(�"���&�UxH�^T^��yU	�J�����WW\��=�U����䞠��(�J�*!������&AUE]1 ����0�ؾ�2A��+�
��Q!|��Ț�$�և��c��o�ݪS~��S�Bm�"{����琝V�JE��+�7Gn��G�\��	�5�I���ܴ�Mr�
���y�KI#���\���}�	[<yҧ����2E�/��`oG�J��\��EvI�l"dH��C=�Rծ�&u�jȊ��U�>��k���V�b��'�÷��UU��f��t^]1��{���Ϭk�f����F����5d�Z;e��������� �`⣭}��������k��-i ��;ɐ�-��De�$���1��J� ����_{��4���0]`g��MD�$�=��w\���"43���Y!��$w?��H�[�~�Or����v�V�Q���&�x�����[�_o�[��(�d#s��m���x��س7�z�Vb���'Z
ȼ���n\&[��q�\�غN��ϣ=��kclԧM�=b�t�]D��Ӷ���VB�o��t�W�ɭv	���9����ȅ<k#���hi�����H�$��	�=�(>���Y�`�����;	7�	^�n�!����>iBA�d���}�*�Kh�_S`�~5�x^i�	"E��_n{K�]|����J��ʂZ�-m
�n�!�����0�5����&W�`�#d�e��'��X+�ü�0R�-��=~�[�Y����[B	ff������h?<���]��U`�lf��=�?_ ��aoy�r6�աf[T_f�9U*�F~��6}��	��*>T:+��H��H��pU�UD�,��h��p��~{}Ep��A&�`�H��L����A����h\��-O,�O��s,��-ǳA�X*-"����޲ڞ�^�OWlW7Є�w7�wƳg��|0v?���Q�"�P��j_L�Ⱦ@o.vK0gw�=�����Si�^���b�276�g����T��4-���kL���u>�Z��ϛ�3�B1�Z	&F�%�j�O���㻕���rd�wWԩ��&�=L�hc@8���������>�q�xu���մw��[���KӇM"u[��{*el.S�,�jǆ]�M��=�;&ԧy$-FO�����.��i�z	�����5m��V�,U
��er��ޏȺ��Bk9��>]f�Z���:���1 ǡ���ћ��D��'b�8�7%���K��f)�� ߛ$�E@H��#d��gY�����B��2���Oxv�k��
N�?!����^[7b�A�35�S�ū�ǳ�yu��M�e�{}��&t�󋻷U����>���9Jac�zu��P=x��n��g\n�>�����.�5h��m�]�����㌋]/t�u�t��j|���<\ƍ/I�Tl�g��ƈ_F�W��$ꃞ���S7���S_^�%��:eŤ�/���B�c�_H���(�d�x*���>� ��GW����B߼yuY��'o��'c`�-���@r@��c49�\��\B�I}�K���w�7��R�Z�,nA�Yk�Y������}��i�r.o�+רq�O�R�֓�,~�~y���oWϏ��\4�����<�D劳ZO��؆��셯y�S�����F&k�+n��o��N�a�A�4�^�h�fD�"�L�!�{�@�ke�R������:�dS���A���M��m��@��jES�C�n�������Q+�������$K����"�)��:mDn�b��A�_/a����S2�5��uA�0O���Fuy_�N⥥^%��5�Ү�F
k���Uc�<��Oy}�B��#��\GQ$�_15�wU�ژ�����Q�+p0O�|��8`ζ��_w+PT*��)�#Z�K�t�ʚ��������Y��L�1�� ��g���69/�����z�hajm���81��[#�����?)�*�>��"��k>�����F�K��N��wNܳ󵠃1�'�l�~(�gqd�9�n�&v�����d)	������{mX�s�C���
���u�3�0I��.���9�s���'������ۄ.�Rm�]���v{��B��ؾ`���׵�}�m�<f�n�z���~��#Ͼd���$��|��w{ń|9�44Jl�\�ۼ�h�H�l�2/#���^�K�ޡ��ɂsK�������'Uf��'9xc�vq�m�g!tЪD�{}����X�+�a{H���ﻢ�ӱ^2U��,�ys��u��������
d�t&���h�p24c���6�TWdbw���u�g)����R�0��]�]]J�._w{ҽ=��׃/���w���d���.�hǉ�	��!-o{�c��q5^y�^l!k���u�My����qC���Y��-���ef=�������mj�|���{vq�۳�%nr(��OI��=r�ͳ��:.W �H
�ԪXU�U[{*`�>c���LJ�W}�0��&N��.�B��n��wV�滅�8xwnu $lp4��j��$���\�t~��"����<��2�ȣ�xɖ�XN���$Z��xfv9�"�]�}P�K�)<����K�I/����za^Uf�Q��ET���>���tt"�lA%�0(й2(a�Q��QW8E���)12 ��0��ESE̳%7SL3<��Y-H�o�_���9�g^�E�m�\�K�y�h��خ��G�PۛI���,/���ǥ��/]�t���-�{v�8�ι�O6-s՞�
C{��r]�y�śv0�Mm�j�tQ�9wOt����v���b��&�х��zݻ\�n�������z�0�ɷ;�l{v�N+���C�qm��'��=\7�;U��R�mڋ��[��e,�@nz�1�:{<��"N��[Ń��Od�ݍ0f�樰�v�|7���9�s��.`	n؋�[vX���HsV�kc�ya�m�j�$�:��s=��U�=�y�S^��P�zG��6�굻i8%v-V��!�&���nL7���5��i6�[����Y������퉭=/M��U[bv�]n��S͙:z�d��x�8�ݫ-��=lse�$���'�Wj���;[m�8�ye�3=�6��7Z,9ǜ��mC�XƯ�fr��O��V`��v+B��
6+l���J�22��E��V�+N����G�\�bY������=;(\�� ș~�r�!^X
��nj��M���	�a��{����JC�i'��&���"r��#�Q��O�LQ�^�Gb�����3$	VkA�U�PW��;���jm�ɘ�v���&s!�mѽv�ի���N�z�I�l�5�z+E�4�έ�V��hu��8ԗ��y����������pK�꺵]�X�-u��!�E�d��$�2��V��إ���A��	)�b��E�`sX����:�+}~���&�L��H��¾���-A�B��H�ì+\.�Q�I3_�Ȫ��Yy���r�([$���:�M�U�}�"�k�\A�5=�%�+B��XR�:�c��7�?dlwy����ahuuL���������s<�!u�~�r��Z9�U��QY�:�9��23S.p/+7�Έ��`������Z�X-(O����`�/�|��z�����'�C��~���Yu�&'A�X[����o�*!�+W��+%;�U�3�H�fb�w�V#�~+p+���
$ș �������͠U.�'N�F����#�in�n�����A����2��n��$�b�y�]]�a2�k��x��^���[����E!�kNy���^w@��&mY��mf�$��|sG�8#Խ\�V��v��EkVЬq���=�[n���Y���:�g��F�9%��T/����t��|�$��$�U�Ì�"J���"s_w���ȶ���&�㐢06���LA�z��'�2WN
Y�?Mm�����7ɒj�`���o[�BM�o)*n�%��{�޲�Yli�&d沮�h�f�Q7P|Z�2.��̻eH��Q�狐��Cη^�I][�}=������j��J�\��jw[�Qg�����������]S�ڡYw��Ϋ�?���sWK9�Frg�ݴ�UX��h�yD��l�w��ixG��a�a�O3��}=o��w�"�d�^�������oS�գ�xxb�r�>[N�>���Kf_XQ70K9���t�}�!�n�T��L=v���5Y2�?_���֯Gkr&��隣d�z�/4�����"�fI[=�2"��;Ա7W�?1R��wb�<mфß}$�dgz:U}��Uf���"���4&���d��5�T9-�9_._U�d��J�����gwRU��Cߡ�ޞ��b�M���y����kK>R��TU˜�}$-�&Gkd�5	���'�N�:e�q?���g����Ȅ��콻�S+�T����$+guw�wg�[�i�y���P5���M/{�/� �у&����.�OZ����Mg����z���Z���P�a$����r�pi7�m�i��&�U�q�K+���J���XW\.����.y�PkY>�"T��'�(I>�Ǒ$�א�ږhH�$�9���ά��uw�>$�5�A��9�\ZA26%pYF���B���?u� �3g5y>�y2;��,��.̱L��/r�h�8:ٻ��Ϲ}*өH:����la�9��K`�8W��c�q����J��<�	E󁯭���U� ����D̛S������IVR������9�� ��������$�Մg6Hv7s��I;9��k.�2=�~W�$�0�>�'�o+I����
p.�HTZD� �`�d���=ɝ ���-xݚoc����Q�'s�ĵ�^�}�b�B�a�v'gZmn9r5<�Ņm��0�]�v�N�r�Iv.J������k$C�mA�>ݝ�1��,��kdY�vq�q.��n��<��ٻhd��y�G*Y�6������I��)~���3�L���dlda��sШD�]���U�#<�#"d��ETNgR��ĕX��	����_��$ȃj.y�'U`�t�a�;��0�.�}��.�3�dMl�S2���׍�9�����J�:P�!z��ڈz�7�|}��/� �� �H��>��׋�z�ul�Z���nѢsW�hz�H��_��3'(v�j�]"ߘ'��ȀBzK���� �Q8,�}���I�l��w$�����~�$i�A �Pd���mi�7�B�'pCkx��<p�o��� ��`�}��}^[����.�&�Q��hF�KX��V����B<��O�|�F�+�����B����L����O�D0G���VAG��S]gr���m�FE��a��[�,9��}ı��NJ���˗{�o�3�:ݙ$�]��u}k���v�c�u�ܕ{Ù|��y�ڹ�^Z��d���Y��Qe��eʥ��ަ�3j�a��z�<����U�Ǹr��Vyv��v�ǭ�U{��р\H���]y��&�|�����2������.�I��̕�&�w�a��	�=֭�J�Uǫy<ޑS�$�ĳA�YS�����3{aՑ@������o��Mn�Vj��Y��u���Xۂ�\f�\�/��B>����}m�f��(��Ւ]�݂��Ee�j�MX$b$�Xl�����G�"�� �SU	x��>�_� �A�k��餕Yx�E$�*yje�Y%J��HF~����4B%+D�'4R4�(���PḌ��O	L�]5W*<J��aF�V��E��FB�yIbIREI��k��P�R��$X�jQj�$W�+���F��D5����)����E�
�jW�xi��Ta��I��Qy��*�J�	 DEG�=�����}l���=
�$+�W���M��' ��EU]�A�G��y��n'���]
j��_v�'��U��oZ%7%���������B�U_�y$���GkMB`��V��_o���Me���6IDZ��,�q�Os�_�ڽ�?yx�h[T��X	>��q��Вw#bs�Rt�L�������g���� ���Ol�lr���u�I���)u�;��Hx�&		A�B�l�+ɔ-2~�a��6���f�&�Aj�)
�S�ͅ��5P���W��;�s�i���4�u{�Gsd��q$ꃘ�(`�T�m�pi���ɜ�٤˞�au��Ƨ6v�W�r�~$�ǫ�ʤ���^e ���_>��ƙ��&O��Q�K0m�5{6�^"~�7�$������^Wo�C����cC(����ۮ�XJɭii���#��Q25l
�Т�uα-�mV����vs�gug.]5�`u�̪��ݒ<ycv��9�vz���p�<v�ގ�=���n.��r��۴S�N�N4���E�٢8�S`�+[$��bo��ܚ�"ck���j��-3W����}��dL�w=��`~PY䓪�Z�$�6H��į^߯�� ���=��Qn��;n��`���5unt�JT��`��M=`�����r��y��o�`�o޷թ�mr'TU��cUX�M׷��i����$����=��2 ����Q��xs۸H��9�vrR�d����t7��E�&�X+:���D����I�%�ՉJ. ��>	�7@�;�@?l�N��./�d���3�A���6�Oo�^���kŃ��\X 	ۢ��1-�4=�/��趢��K絪���?����U����5�{�;�y��&��|��G]+�-}�n�������#5�����qX�xP�M�EF�"���w�NB.�ڽޘ˝�b¡.���������A�a�������v|s$�$4��m<ȹ6�'y0�䅨��6�r��+�D���X���3ҰLY*�Q���]��b5�������:����s��L�˱�6�XO�^�A�pYT�����w�ˤ4��Z#d��-Voe�G�lF�,�־���f�Ώ������pP\�V�MJ�}�0A#q��9sh���13Rn����i�Y�t������ui�ʫ�����2�dL�>�������Ǚo�&׼{�>z/rw��S���$�rY"��Orw�N�8��j`�r6P����Z��Y*{��3鍑����s�W2	܃$Mop�:�e�L�*��q}QY$\!��5ɒN�s�t�L�<K�݌�L����4a�L���`�r��1{to���4Vt~�د$��p^�����m���������J�#[޿}�Ɍ8+��6P�*-P/g�<�٭�6�jm���S��f�n�%��D��ힰ��vk퓲���I�^�m��Q��¹�p�`��ݓs����[=%f���'F+]�<�2���M�"]��es��!����E�a�CK[�R�4.�df��]b�`�^�__6~��$�{;d�Z�>�*�ِ��g�PцH����KI���i���_{9����Л{�z�����RZ� c���Z0�����];^\�������yi$��~�T�^S���Bæ�ߩ*�?��3�]�N�@�(B>1ץ��ی2G���xui*]EڎM���7��VV�I�>`��w����ko�ƽC���zK5����vU$*c$�i�Y�b�l�M���8wN�wzR;l���T���;h*u}��4�g��2&���3��Ħ���B����A��XOĎ��I��)�ܽ�|��b����"�`�IS��Y�|���E��V#SӉ��qh�e}	��lq�&I�L��Ⱥ�5�1O=}m��l�d�^����5�x��6	Nn�l;䷎���0&�&^{�m���:P@�k��	P�jjҢ��)�dW'�y�6��E��U܇72�5t�z�1���q7h2Or�za�W�Љ}���@��U_>@^��ʓ��)��-��I��L��1�2;Y�i�u�s^7����zO����f��}�}mͻ6���"��&�V�-�w��O~����^�������Q���:���cI�:�["v�s��S��k�~�Ț�����M�g����QVo��-��n��D_&=�0g�7�5��J����������� ��5�^�B��g����5>�a��m����e���.$��'Q�w�+������y�?��C�/��$��*I$�rJEQ�����T@~��
v
��ޏ�d�`��kU㢋�~^����d�!�n]�l�*�E�XDUAP�	 P�T�YO3�S����V ��ik��=r�D� ��Q���>��������{���c+�z\�=�k��p5��f5��������ך���u�7��T@x���o����~`�4�Ԁ
��!�@P�_@	��������=(=����A� �0Q��[�������0>�!�J=��
�����X~�� =�m�!d\{�2�Zs�&�� �`~��h�_��֫�P��_������a#��.|�?�3V�w�,
�7�ȷݫ�s�HO}� ����
 UB� v2�H.�4X�yV�5k}?Lc�<��s����� >N��
��}�8�=�?p��Jgʞ��y�^վ�/`���_�O��P��?y�����?Ə��"����i���a���>�?�}��{9/G�C՟:��(
+��+��������`40�������o|��?��c��|�T@}O��u��{FA��y� u��z�!�iG2�G�Hy"��e��
����Xu��Ƃ�K�`o�9`�G�F��!�.O��!��i$#�͉렟��)�PE�H`�=��d0�-����J�$?T�&d3�>���RoF0_�-�.*��������=T@e��/���?P�����;9�x�=���������� ��'��G�����"}���}��-�=��K��B�T@~�����y�4Y>�*��}��$������?XΛ��C�7�����8��6<���xL&�9�R}�;�A�����y@q�!��;�c? 6A�����_�ucN�f<����*��ܾ����u���U﹔�٤������~�z�>(׻5���\��_k�� P�b��=`'�~/��OS�Ow� (�a�֑r���hr8�24�Lj�;?+[@�!"�Շ������=���.�p� 
-��