BZh91AY&SY�Sc�A߀`q���"� ����bI~�     �G� 61�RThـֲ�V�hH�4��EK6��i��#mH��R3l�e� hTkJ+T҂�Z
��dB��5J�V����i�l4���M�X�(��R�j�խ�Qd�
����cIH
�T*I��(�ZQ[�V�� ��)[4�fQ]�>��A}�4�݄�I"P'�t���T0�6B�)Z�XƒM�5(IF[e[Tm�`U[[fʶ�)��[jѶ4��m�U�L�[aF���j�j��3%7�  3��f�)��%Um�J�\ګ�f��4�-����v��1�F�+v�:���TP���@�v:ZiF�[4�[e�c6̦�   �{���tzh�Ü�=�{��\�ܡJ
�۞u��Ӯ՝)�d�rE4��Ǫ�Y��m��݀�W�{<ҔUS��׷�{�J@����m��lK\�'f�3kX�6�kh�%H�|   ]�v�V�jK,��zU=)Tu�&�{`4깯n4um��U�ZSv��s�T�s�>�/���������}��V����D@+鯾�}ﻡR���-���i$l�m���  ��Ҁ}R�m�|��CJ}m��Oﾺi��vw�<�S�Mow}{���yS�i-5��/���}���Y	�R��ow),������N��>��^�W�[<��|zcm��_=O5hI�Z�5�)��4��  �>{��K���篶�7��|������z��ޞ[�g�4�_M}��^_<4>��
}�O���n����}{o��8�|���z�ޛ|���nh��_{��JW��n�J+LT�k6�l��R��  ���e>�T�����{R�����wv�֔�4���z�J}SM.|���/�����s�RS��O*�Δ)�p�u�m�Һz�uz�]�l�����=���[jk���[m5TSMI+mM�|   n]��.��Cmz���gU�;�z�駪S���*=��s��q��j{M�+�F�A���yέj�z�Xv� y�� yˏ@ �{l�-f�֪�kl�-j�   ;< 6���=�^�A��vu:l`���U���:�۵gS�F�i0 ӯy��h gvqTh+�qz�JJbJ��IY��  e�GA�-v���v�5
�\�g��n��(���=^ނ����� ��;���b�ʻנ���@�ՑA�a�V�  3�(jb�N7N W_]]�Ѣ�7]�  �,t+��=�4 �{��Ӡxs��=h{W���oT�     ��2�*@L��0 �L�#LE=��R��� jA�i��"�����H h     5S� SUJ@     �� ����?j���̦#�F# ����&����jG�A�@4~���>O�?���>���,�&��NX�xїq�����9���||W�=����*+����U�*���**�������������T��
*+�qU�p�`�	S�`DW���_��G�ߩ��$�`��)��Ι^���I]���� n�^��+��1��:H�It��.C��d�� t�7L��Q�dN�p�9� p��`zH� �p����2�$n��:B�2=%wL�H[��.�:Ip�l`N���+p����0� �@�"��p����2�$nN���+p���0I[� � n����+� �2�$n����t�.��a�%� t��2=$n^�#�0<%.���G��p��7L��V�:@��8@!�P�2'H�zH郄!�V�8@&� ��*t�.��HD�"#�@R�T�*��a:B�\0��%7L�S���
	�StȈt��dA:@�n� N���H Ct�"la�
��HU�(��TB�P�"	�eA:J(\0
!A7L��IE� Ĩ�Ht�t��`:@�n� N�"��HDM� 	�P�� ��aA������ !�d@:B \2���tʣ�Q�^���z@�\0�%�2���F�G�� ��@�"p��t�Gt��dzH��7/I]�+�F��;�Sc#�V��+�dzJ�2�$� t��e���\08��!Θ��� t�7L��P�d���:B!��2��[������ t��2�!n���S���)�t�u����=|�>oPo��u[�t�Wŵ_˖��B03�E�0��n���v�&޸iK0*�&�dŴ�ɺ0l��Ѕ�!�c��g]���(��o�0:��H��n	�㳖�c7����+B+5�Hh�"�V�5W����ŭ��x@�8�U�8I�՗��Z]��s��#C��V^��Җ%�`��q�3A@��Eb7{X-�UZ=���ƀF�I�!;b��)L����F\p���I�e�К�X��#��f��5�������,�afH)�s,=�53%�	�MND�V�o]_�E�u���m�� ���[�!��q;V"��XkA�ZVV��!� T�hR��w��3>��ֆ j�,�1�6�l�a��
M���X�#~6n��y��z7o�[x�R��6<��� �T���W�ۍɬM�ō�҉�m^9�r��.����W���6��f|X/W�$i�ˆ�� ��@N��YB8��T��C�N��*��o+6n[�p�[Z�ҊG5$��Ͷ���	�i�e���JrC�h�(64�m�˥B�j�ZךԗQ�f��@�m��f����ٌ�.��)����b\��k�E�㳸��r46�Ӫ5�bVq,!������vӚ$�J����ڭ�b��Q�̶k�[��	2[�cz1��m`x�-��tm۹Cr�o�B�䩦�ӁJV���l�َe�J̈�*��V\��I�.Z#�)�w�0����d�L��(P����jc����C3�k��ĸ��I��|y�����4 �#�g@؄�oP��Kˑh�vȻM7�=�KM
ܤ��5c�a#���m�By�4-+��uY,�����e-�gr�Pm��ӹ#����'Ҵ���Y)��A|�r�X��u�~�oFM7�Ţ����P0�A��1gQm�1�;��ǘ�ڸ���v ��-*�l
�[t7�aYI֗n�/6m&�9�T8-`�0<��<c�n�˱R������	TP��m5�U0]����B%�Za��$6]�����f�ҫvz�r�9&r�Ȧ��n���`���i�a#.��51����2�Cg-��/sv,J�$R �q��va̕����b	c����Z"�5ҋoLF؆؆�9]�+
↺���}�:g{��:�ۢ�ěx���m�vQ@���j��<��1����%yj%&c�o����Xw9�/�3�%��U	Yu��jk:w5[Ȟ�ee��>/��J�G��+M��M�9Oi�Ͷ5�kl��� ��hSe�~5!�Bd����k�,?�lT�F^�qG�l��r֙(�#*�=�2Ҽ�5�ռ�R;x0l��6��m�[z�^�	im)$����&��c�C--�N�ڡ�f�=E;V4s�7[Ƒc�ڼ���tuc��1R�͒'E�� C���ѯvaPŮ��%d�xRN�e�����7���2����ɦ+pY�&�7[E�Z�I���n��:m���u�k�K.��+ɻ�Eĉ5ݹ�mo_\���N����5%i��f-�o��ii���Pwb�YfQS`1x�h*�0�;�)�zu���r���O��'żr�:ʡ�	])�k�\-|>ə���nl�n*��ш�SqeM?��Z��.��3rܖaֳW�Y7r��+����2QŶ�Y��E�$���.�q�{[n����lm# ��/,��!��B��7����P}����[b餵�jhh�Y2�=9z%��piDY�ma؉�\3�ݑ��T+��i�Ϡ�dfi�\�hYz/S�	jۥ�A��7Pdln�M��6T�}���Eze���\�/V���q$qmi��R�t*׭AXZU[�-܅XBRT�E�{��:���[����	���	�M&�9 �)ea�z�b���K���CJ�S?q޺Xl%�b���R���*�^�]<?,������dƨ�s����$<��Q\,øk1E!���íx�n�7��)KXA҅b�����B�*��>�Z3Dg�����m��,U��L"�k�����.on�����u}vF�M���ؽE�zj��K+$�P��҃>���E{F����x$�ROF^S;Q�u�	^S����@Ф��R`v�6m3OZ������S!�*A5<�ӂ:�f(�lh�����#��Y�/�����6K�M�����=nT̰�XHR{lҠ�Xi^T�N�W����h�&�@ -�GVI�{����'��8���`�i�PCX{�R��6kpX[�<�!�ұy��a�̛ktf����bԷ;��B�S*���/�Lͳ��# ʸdGs�y{�v#SSM�5`�Vɢ e&P*���]��v�9�2���Z��z�V�s$
av^���r�r)j���MX��Y��O�����m�D2X�|K���Ҕ�RDY�e�t�2Qs���[7n4<|+]�Z�c5ʹ�2l�i,��sui�Jkn�\Q���b�Ǌ\�f�A�5���0��k,��VD�r��8�fI���N1Z��-MGVG�NR��rd�	4�=���-�*Pf� 2:p,Uz��óM���a�����1�]l�cUp�p�ikK�kk)L����DMal_�Zڎen����\ ��ld�ۄK�L7a+{[G14��a3b�����V�}��i����5��kst�//4�h�g����X_^����z.�!�5cI�\�1F��1����K$�v��9�R�E��7hR&V�d�k��E�Քsj5v��cOS�=��B���ӘѽGr��͸d$]���;��V��`Xv�"��ou��*�m-�nm�ݵ�۫q�]�6f �R.c�u�4T"h|�b���\B=��F,�
r�J�v���̩Pm�L��%�Q����hLT�N�Ѣ�t���Rx3wahbt��ЯM��F�!Qf����W��<�Y�zq�̮���}��J�X����d2ooK<����܆�*"��p�=�c7n^�br��u��Ֆ�$�1f$��_\�`���_fe�Z�{\P��3z�����4�g���`0w����Vܴ)=�B�mi�(ͫݡ�e���Id��xa�[�.�d�i����{��ÙFYlErG����.[�;"��+�/��: <S�3�Em�v� ����UeV<��X��d�P3��� Kcum���	�L,G_�J+��l�S�4��c8>�0�j53�L*�mܶsL�� V���v��Q�5�Ul"j��9r���*'���Hڳ��m6�)�Y�h�Kv���ݺXt��9ڽ4�Ӧ�If�]�j܄f� �f�J�5��ˣi�r7m��jKCܬ)\���"�VE%�!VֺQ��֎��J9wpJ�1���,F8�2���t�GMRZ)��!V�M��gQ�CcFQ+4-�ךm
�D� K�z\��QRfɈ��l�k6TX��&û �����M%��op0�]X�����J̸�ÕG��Z��9�K�c��-<��u�ɲ�Oa�:��	�q�ej9J=˵���.�È�_n	)|�i\�f�z{Y�F���5��|.B���;���(�ʟc7VZ�i�N^e]L�H��H@K��F^���ś0�R_�P�4e�w�t�mZE�j��r��ő2�]<�5y��q�3N���c��JGT ͥ�*��{������+H�t2�a#���a!6���ܭWq50Kn(q��f�x�KUv1i�џ'J�G":R�/J�F���C ���X��[qۅ�Nn�[0Zj[����ж�jU�*�\�U��a<�5#��اx�[�.[�x����`�ol�Uj���uuy2��1Қ�-:��U�Y
ߖ){(�`��M�»b"tA�����Q7EP��bb��G�^E��xV��h����� Z\	*Z�㸮P��,�E8��/E��7qU*�F�5�FFqk�,��ȷ���]GY�I����dt/Jf��TyxL�5MN�^����Y_�K������p���dj2me^ǧn��ۘ]�.nd�Rߋ�	�`���Xܢݛ��b�G4h6ʶ�դ���!��{��*-�gC�Vm�=���l[�g�&�2������T�?��͛��h��4 #%��LW�Ľ�.�N�啡$�6����l�Cr)6�f����=���;�t���y��/Wېm*
ؘ�^̰0\l�cW�n��R���.���Y\�+�n�9�՛ݨ+(�����O^eBH���)2�m�y���'�k(�b,ܗf�������z��[t�2K�k6$���Y�N��R���V�K�N�͉��CB��X��Qȳ0<Q�5�50<j�6��MtVn��'P;�V�\��������ŋ�n��� j-ikpTͤ�O���@�������@�e���g$�i�lhQ�s%f�HM
 1T���Q�ǵ����S'o[�V�;�v<��lZ@�SF�V��v%��0P-J$,����u�*�u��+y���#BKE94ޛnż	J�u�h	�eպ(�*:��e���ͦń�Q��l̳R��1,х�_�i��դ3�J� ��O+�T/p켨���{r�-%M����˶���Q-U��2���M��zݔ^��,f��ݤE���K�S7Al@^k�.��5mm]��k=�J�E�,u��a,�[�<}���ٳOIky��-lu/oU+�NaG�B�$�Pb��ð�Z�H�4�A���q^��<���r�ǥU�FE]��mm��Q�y :%��,e+X^����F�9�E��Kp���2��Ȧ��:j�F�xAA*Y6�MŅ��r�T�.����TC�+f���M��/J�)m��vY�.iv3s5�"��*v��,0��J]��]]ة���Z2i�oL7g.;T��/0jx�݀�6���(Y��c/p���������d���ާ/R����֫Gn*�(�p\�Rףel����H��3P�҆ݸ����So^kݭ����6a7sBq���^�P��h��0�<l�C^��K���YBm�$�35eX�`��ޭlw�Pǭ�n�o��-�i;�?=e�yF���r�f��0"����V���`����cTw���:ď^X7�}�&�6�v� m��{��T6�۵�]gR���v�Q��M/�����P�.Y����*�/q�;;Kqf�[�jBΰ��ݸ�:Sе��ed�a!qĤ[�pi�'�@��!�Kw����X�45��h��I*)W���OL�홆�b�ܭ��Q�nVRX��*L[��S�fMf�5��a$L��J��Pe�v�LWn,u/cջbZ��U�U&��1�eni�n��	+4����l/Ǖ��W�)^�n�Hò�Vm��p�)=�V�Z��kL���;cu;��%OF�6����У�թn������9dV�S�,|�f�Uw��C1+M-��qCo6�u�H��b��Jǋ�V#F&�U���I-��hPz�n�ݷ�"��Lh3x#�kjU��.��yH<xU�,�86ص[���f8��q`�B+Y���r�4[.ޛ	T�fV9lcp��n�؄6jG�5����6hf^i�Ŏ64�����cxXa�.`�(�j;!�h��i�IGh�Rn��֯h;�"Q�{�w{������ⷻ���QZC�R��,ޙy��M�{����K{I�'m�h��RW������T��hmc׬�k��DX�E)4�V�U�ni�Nn6�+�i�δ���\o]�hQjnY�2Jk.�q�b���F�ϣ�3b�7o\�nV}�[bP˘�y���2�8n:yI�݂�(��aK�t�ə���Q���ZԤܹIi�un�4�b�l���`r�;јo\�X0Ƃ�Y5��*͂�31%J���Mi�y.8A�u,�n���l��BlY�
�BG�nYNݬ����K�Vsi��@?^�t�����p�S#Q�Ņ�&n��zг�v�����-�딪�"aͥ��L
Z1�0�&a!"1�E^�
��Qā���F���Z���"㥛&@w**����s	v�����Z�Z�
J��! ����nX��z�ޢX�K��m>z�|�@��`�`'�2������ڪ�nQ�Gu�Hl3�����a�o/f[wq��՗4�Y�e^��&�\!Qn�[��U{V�C:�搑sh{���CE�.�,�쫒��F���-�0Zˋ�P�Y��n2��b����h]	wF���L�c4�����udoa�f^�h^�WM,dM��<�7�2�h��[�C�ǳztmS8�v<�6ܭ���Ԑ�����:x��G/-������1"��.8t)Y��X��e�N���z�Z6��YJ`G,v�
'��as �s7��L�'ں1��PG>��(��M�SoY�۲r$�����R�k�,����.���6TD�̴���ۼ�$m1�ȡ�]E�^�Ph�A�����U'��MA\8S5)]Ay�*����jdv�2���U�y��4��w+�L`S,p;�D����>Vkv��n���/�"y���*7�JB�6l&�;�	�(Mݝ�Q��{s)�8uJ�a��1��jx���^]�y]V��b�� �˒�f�������B������P�L_+�f����;�r����]w�{]l��:Їu�@jPu3�� /JzK휏D�:�s
w+��F��M���g�M�~��㔟-�Ϗ��e�`�^�D���*�f�wev���Z��z#�RD$z����q����dvrJc�r�G�����'��W�}���v��� ���^��(��#�皯���ߝs���ޓ[t�5������l���\�E���m���5��sU����k���r[���(���U������0dy�<��u��I@�f�$0�cJ1<�2�����YW�{i3�ě�z��k젥�s݋X��Y�E't�L�K���j���i�;�p��ص�{)�)�Y��Xgsf�}�����Xݺa��ذ|d
^�qd��j>�:�4��&*iv�lk8�=�F�e���4�{jl�:D��P�UɁ�"\*Ժ�:n�QA	-B�͎����sn��j=H��xY�[�+t5U��r�E�Z�l��(��)�mK��ic-y[�n�=-Lm�L��o��c�cnZ���e��I'c��*hfX�/���ਕ횔��V�5h�|y�Y�ݴ��g2����ܽ�l���y[z�qM;S��}\R]�oˢ\E�w�$TeΒmN�MlQj*}�K�NUH5r�uo0͐�㬫ɰ�^�o\7�m:^N�!^�V�H8��"vحɓ�u��Ca�I��˝!۱1Q3�>��gw�5	�t��u�ˤ��g�Sr^d}G��cӸ�*'��̬��EB���SǄ?������;,j�X0�Iq��Ԓ繆)���8pІ�v��tSE=m��M�P]ҩ	���<n�Ү�d--B�t�]])�;1�y2hJ�<�X��mШ�;d�ٛ�* _
ٮ!O�+ڤ3v�MB�2�����0$�f�K�Ы�w��@ğ-����
u�Cm
�wI4R�z�clv]�7f���p#R1���hp����s��v��yWQ���]Z�ݬl���&�;Z���zث������]����#Ɉ�Į�'{����FI��R��\J|���`��yi��ح\��d�o4��L��v)mQf9��G�͊�ϲoc��ZjIF�����]�R��.A3jw�}i#��WX۽��?��6���B�?KTM�K=��0&�F;S�,���"�#��ˍ�
1P��vN�t\����p�
�U�n�W�_�Z��]��$��2v���|�+���MN���n��}\i�7J��է6���1�Skk�չy@┱.Á>�s���SH,�K����:�]��/�;4�Ex�DA��3��P��t-_:�MQ=��[�VAӲ7W}���A�jnm�lM#��ئ#&]���[���`<}���C��4�r	�ή"�趯�\���4[�*cj0�ϵ�έ<�yz�U��fu��oKH��a�q�Y��|MZ�)�9�!��D��.z����fa���kl�`cf;��E_�zx�F嚆p��Sy�]cim�̫a�Ǚn1C;,6�\��D�u���+���ck�Im�/���׃�U֑X D�X35L�hc\����k�5f��I�w�{Z�&g'�n��6SJ롰�=�o��+E��0�&�Jv��Kf�����!�RIUv/r�Mp��2g/{F�ؚ�w�*.���u�ҧn �9��!�ʀ��Y/k�u��5Xz���̳&��ĕ��K{�Y��
�/�uq���K�ֵ̏��W�B�Ez�1����r{M�m��b�?e��o���9��P���5��W�x[���܄��ѿ��X�2Ό,S�'"R�V;QJ��x�����u��/l��w)�*8�\�N�{\iJ�xR�Ps�'r�k[�$����n���i�r��Y�Rwr2w��/x�&өs箧3uһui#L�mtaPT[����+Y�_KG�d��d� =ҹ���=wV7��]+�1*w��}�&d`��m����˭���oL�]�%� ����ˤ�3�Nx�7m����*'����̩��v��
˜#�pmѫmj׳
�N�U3��ƻ�Oj|I:�8}6L�#/r�mS�	�OJʴ9��l坜�y��TXWDn���&ZC���cC��hP���(�z��^���LV��Mug!����sM=09w�yW�*Yn��&�&��I��w�ƦO�!E�l
�KS���o��a��[Ǒ�,}�!�X����i ��,8,���bU�v�a�S<&�L�&v���9ci��	A��������u�r��Y�:��G4u�9s��҄�`b��j`�f���W؞���B���i�ť�6B�SC�]gc�g%�th����Z�j���QCQ�'���W�f>"j��,,ݝ|eȯ3��6�,���K�f�{J>��[y}
��Hz�iɚ��;���|;M�^b�ۗk�����_AA,A[q/:����gw�T)�سnˡhS�&����e�Ʒ` g���m<�]l&�K���q��Оζ^x����!�+j�}~�D��Գ�&�<�g-���ev�Aܫw���h]GG�t��3�Udi��b�|�P���rfm�:�����X����z�� ��X������ol�<�h����b�᲎<s�]�f�߶V���utܪRtǂ.ڒ�N�X�DI%�VuA�:ѡY"����i�n�᜴�hɳ	�".���gV�;�<{�t��X��ّۛ�C�e�:��G0�f���{:T?L�����6z:Vζw�U���O��8�oC�	~+W
�n_GQ�؇	�֞�m$� ��^f��.L��B���\��*���a���s:e`���5WY�+eÊfL6��\�C�ʝ{D�@�P�U��&Η
�K.GL��V5 Ul�tg�Ʒ������0�E������E۵ֹgQ�kR�o�v4�l.��ǧ>�(v����{�ڏ���6͹�<�5�kEJ%�~����aL�yQ�v�b�q닶�Йwu(L��T�&c�Ψ�N�����y����Dc*jͫ�h&�9�h����N���;�e�ܲ���[����ȥ�v����ZJ���>���GQ|�:j�3 ��X��09�L8���|�x�;_]Y���P��7}�#�uպ�L{;Q��|^��QjZ�݉]�v	G����!��+WXC@�i��A`�zv�˘ ��gY8�:n�r���o�q
�'R���t�:���.k�.�"%�j�f��&�,���@5dF�d��3��)��E	+1�o<�4e����tW)��ޮGt��ͳ�h����;!�\�M�-�&���p��]��^������-NxI5lɷq㱌sCv+������{՚��&�d#h���;��EiM�C���r^�^��c�0a9R�
�WI�Y�y�,6��|1�OEo� [�\��f�p���G��i������U���j�Z%BC��.���81����fe-�/�J$��p��W�I�/WĝZ��sf�+[��sR�O��c�7�Ae���K$U�F-�vL�4s���iD��*�� ����̰��B�t�m�.D�޹A���k�.��A��R�;�c���L�g@5�9�¶8��&j���<_f	�^�(u6:݉������e�̣�̲m�\,�r����"g�gA���x�m���i�6��������������aރ}��+v��^P�8�8��B]�!�8G8�zs�pHOb�
�rq��}.�eY��;|wsZ8���o�_�%F�P���їp��=C�H��H<`P:��gi鱜̏5U�zɊ���g��s�]�YU��6f2�«:��/�(5���֎	��x$���z�k����R	�\��K�{��wR�x���!���U�3�ے��!��`uh�D��=��dsyײ��*Y.P��ES��t�g!%*�9SoWn5H|%�*�dU�Z��=�^�S(`Gvg*���L��8��&���������;���Pn���ue�[7��R�U�x����O7���P�ߧW3�G�f�w�NJ֐���	��p�J���4��iQ9��J��^
o2;����gi�]u�b}d��p:NZ̷)��*�Y�q��:�������Vg� ���Ǘ[����{λ��'2�e0�I3������l�2��!����(���8�ǚ��7�4	O��0V./�m���tu}�
嘮`�X���v��d��fp��`�6���_nS�e*��܌R�����T�
:�E��]���Q���&�:V�|��#���y(�5�����[{�r�m�1�J�J��>��qXk@:Ηx�1����z����&��ɼ�L�f�j֚V�L�w�n����K�Q_>@jg�rr��M��Y���s\�䛑+�ݬA����Ż�����ǀ%��9�"wF�(��f!��t^XZ{/�}�u sS�����Sӝ����ٸ��n������]�T�4��F����NX)�S�o8Ҭ���n�w�i��iM�Ӓ��F�4�\(�lF�PcH�Kzv�ԊS�ϩs�zu�C.��&c9}�'_w�ΰ,[姇AE�����t�I�p���*�M�&&�����35���4�^,@�P�y�f�N�k&&4(�5Y���K��5Y'�}oL'����[K�/��59�)�a2�0���J�}i���e6�b�٧Cx�(���l�{t� �&l\��߇[AŽF���b��^�.��7ܝ�l=C^Z�v���9J��a��[ќ鍩�@ ��,�w�,F�}@���`�ͬ��+e�����16剶�w>���±h�V��F�ӭ�����$Z��$.I' +@��v��튇����(���4+h��/]����7��	'1�T�=��Բ���y��0;d{{we�䲌S��j�̄�kwYa������ՔkQ̺=>�{g�p�s�H{6M��]g�g`ϧ[Nt�0�`|������X�Ygo�zܚ�t*�%��'��f��c<�>{�$�wQB,�G)M�kC�HNV&�ژ1�'8o��ԸV8��i�A��)�#��ʺ�8/�{az鿃N�Uݓb���:�ݖY���	�`	
����v�-Vup�o�&��u�d)�U��K�ORJ[Ш2��}�8v��h�7�2V�є���"c��'^ݜT~�ގ����Yg5t�A*���x^����5%���m>d	]N�v��Wn�B��0[W�]�Q���R�5{an�ա��9�uu����X�*�N��N3\s0S�� ��V@9;�z�#�����c�\��ֵ�
��e�n���53��������0��-i)c�FW*\�1i��65N��J�� B;��U�M�s4w��Il��[�m��T��3���̅���]����y|
5�sSC]�6hv��
*9u��Ue����5������[r��n�7o�p{;�m
�O������$S�W��H�"䕗�OW^\�w�鰺���6���<�e�Y+��t�-�BsO<%��Ioi��@�s������%evl8e�أ}H�Ur�:lN8W�^�V-��vY�E<\o�O.T��[9H�B�h��ͤT�e��{IS�p}G�N�6���:���l�e%I�s���o�-��Z��Yg]�[��s�CC��b��9�P�q!j{m�`�):}p�؟A8��9��WIr�a�,G4��e:�����f������FD)C�F���r�:ne܉�tV42�2��Vd5��o8��I*��g6�;�ȁ:�T���78�n �F���{lۼec�	��n;�L*������ɪҫPY��7-V�z9�zܝwe���tqXْ�r�^u�WԢ�SR[:m�C����Y�Z;�́摑���7�8�Kی��;Zci���-�����VS�wήWm�>�<a�۠���IU�q�̰�d�J�M�]j̔�N%��or�h6�*Gi(�MR�������mj->w��Kn^����!rY;W[�S{U��>(���r��}���Ӿӣ���_ $�٦L�2έ�<�Sj�Y��r,�ZQV(�L8//���-s�%:���6�&}�R9��Uml��x����Ajs�,UI��A��%a�F�hk,B�ݩ]rl. ��a�B#�Yv�Kw:o�N-��-wV�*�МY���{���6����ˎ������R�2u���9�Zc�&1���}cjYk��e����}H%'�(�n�s��+�6�P�C�H �R74;�Y��a�P39ޥ�������ؖv;�%���u��{K]�ѕ&����+��v�̸@�� ơ1=Ǵ.
���`��U֡�ar�	�r�oY�Z��%���]]��Ѽ�X&%��0������v�k�����M��wo��H!��j5��&uG��d�5ř[kqቓ<���M�dQ��]򫋅왰�=o�z�ND�8T����][��ҿ�����ⷵ��ZIg*=ݾ�gGh+��axTo$.������C�_G���z�QМ�<kt+�%��#Yݎ|9�8WflU���x�p]�j�P�Y[�B��f��}�񱃌koc�i�˳[� A%z�v�@]3�8Є��څ �9n�Ƈ��B����+�<�)NUv�q{����!��xmp.���b�q�H�\ͭ�Q�<ҿ"n���0���X�%���t�yk�S�����`�=��r'p}ܣC��
�V!݃:�R��7KD�;V�]�L�MV�lj͋ͩ'Ow\%�5�6S�fKw��n�I"����cL*I!��w�I(-Ïv�f��`�K��_�tm�J�a
�=�6A�A�]u̠c6t n�U�Հ�Wr�'�����'���(��y��@Y���P!�(R����q~�-۠��V(S)	K�޲٥Nl�"ܦ(�	3�,���������v�JQD��#d���	@��vU%a4ԟ�R���D�;��m (*1�*�0DP������
;#�l�+�y��*��m
��ü{#`H��|f���=�x�{�?H/��  ���?ϟ~
���(�����0/��~�����|;�>�K&���&�GxAV;]��6̸�eJB��B��z�N�E���h�/{
N9���W�Է�����ӓ�����)KL������p����n����P`�d,�y`�M��T��	+�.p�c:V�̍[8smG��[vU �ֈl�I��KE8q��y+��Hf�2�t�|���!��(u�|5���[��(!�K��6%!o�P�h�Doeh�sv}��'E7�p������_c0H����ȺM�SV���s�8u_n57��ھ���w�T:�2Z��ؾ��6�T��pH6\�=9���,]���>�3;J�(��7���Z/��\�ҷ9�s�Ռ��ڤn��N�ۨ����ngNߔ��6�,�VK>�w2G\�̒+� �����gn\��o`jΌ'L�N�u
���"��ݶ�e�)GHauۙ:�݂z���G����b�q��/M��,�ݱ�C�z�i�s�ӹok�ba�f��M@��G&b�Q�I��mެ"�,�8k*i���W ƿ�!Ml���^m�m�(Jfd�u>�J�VgՂJ�3���&�Y
`8*Ac0]n!���r�s#ë�Ej�*L�ZuGa�:�4�\�;��Q|�n�f��`9�������;!쑕zI�g$�6/t�V]8�s���\\m�=QU޳�ݭ�AT*����wLw\�����}>���}�O��=��o����o�����}��o��{}�����=�>�O�����}�=��o=��oo������}>�:�_��O�����Ҟ���sU�r������Է!���OQ�"׽�^��
M-	�]�/"TG�NK�w������+��io����E�XM�]�2R�%�噵�5���si�������%�k�!״����������n�灉Ux��f�9պ{Lb%f�;��!��o�r�Dj�u����#����ѓ��T���|.t�6ƻS��PK��ovyB���8�����pY�Oq(rR�Uһ��p�����gRX�%�>�d�3Q���d�7XÎ���$ڱuVc��!brwu�:4e�j�pA���e�pΰ"�eUNy�Љ�(�v�rE36k9�kS�49�m�Qb�5��Y��q�����C���'��&'ڋnP�X�j�h�YJ� �fmmH�ŝ��es�	j�gf,��ǌUǐ�wPR&on���ƻ|�ᶰ7�ņ��h�fd@7e]��5����Q�]�%r������q��Q���n16��|�e�e!��ֈ�DwTB[oNۡ���r]�YV&������JZs��QT5[����W���>;����f��
��G�ٚ�{0�6Mn�(da��w�sod�j�w��T#�
�x�5��=�o$ـ����fq�+�u���=�h����
��W%hO�50³vk]��G#�f����/l��o�N�R�<�I�;�%H<�G�Kk�9Zw'��3l�&E�޾߇�=������}�ߓ�>�o�����~=���}��^�o���A���}��o��������}��g�����}>�l{}��o��tWD$��K'� �C�b}»�j�s�[�`l�b!$+{7gN^�Ӓ�6��wn�pUR��S'V��H�1�{ݣ^N�yJ�S�v����Lu)ɓ5s�}��Wܴ
Z�R�>ǿ]�ӬB��8w�Q��ѡ�D�����wt)֪�\MbwfVw��G�բ�UM7��=)/�<��:���4&8m��pN��.5q��Wh�*�)���6�.i����<.�'�PCՔإ�s��ɫ����X#N�U�逞����[�w|5�����>6�!yy�=("�^����W	�8�wD')\��ű*��N�����R�F4�m[[�hw��c��h��
ε�%�wd�tH=4�N��U)`��Y�1wU5�&z�k_ZQ�Gq��|{����o	�滳ڶD���9:�b �4Z�[4�Q�9/��٥�b@��F�]���X�8ֵĊ+�;4��зr�m��m��`��۽�b����bC���+G5/j���݈��3� �c߫d\�Җ3a�Cn�ٯ{�r�;�Z���.XѬ�Ej��=C�'�-R�I.c�RK���w���k���g-mv�V�ˍ��<�:w9O���T�����P����Ie_,�V��h<��,�eq�Zs ���Ç8p�Çp�Ç0p�Ç8P�C��p�Ç8p�Á8p�Ç8p�Ç�Ph7X�f*{�Ƀ.����>��c1��D�ϱ��I���ep ��v�0B���N��Aj�����hmA��$M�!\�X�=j���M�W3�n�r�ǐ��}}�"7�7�庴z����M��G˵5;~�7M]����o�*�z\��{z8c��B��X;&T���;�ū{�ݻ0�ɵ�[o{K:��Hdڸ0���"����c��IM�n�Gd��Zu���\�F�S�m�ux��ܮB뎛:�Y5}�o��k�l�.��8;�3��^]�s��I�jZ�v:�k7J��6ȸ�x���z�^gb�k}v��j*xP��ܶ���A���`�V3+3OT��a�@���0uV�ԕC��ڴUm,K.A�c�6
u���R8�՚"��F:�ҜfX8����;8�m@�m}�N?C�giQ�t>�����ZEu�Uލ���.�(�W�_D.���}xw*ִ�K�u}�Rn�,p�{��Ј�i�R��DWnk���q ;�.� �_'��Y5.^�d�j�a�����`�d��7z C�3JRi��ssjp�#��	w�NH��ݲ�PP��l�تk\�4�t�R���\0�2٥���ͼ��Bu728�Kg�-:%���fA�-�˹D�c���T���k
m�ʅ�m��ol"<ڥT`����`!� �0h�Ç8p�Ç8p�Â8p�Å
(P��p�Ç8p�Ç �*T�[R�J�*V��r�}gsi}��v�3@+�F[ںiA]��g.�@T��:o>R�S���v�g����.��#�і̽�ݒC{F��R<N]�0-$h�)Wj�܄^�'2��˽�8v����T�x���S۔581�+�0[�R:��5����˦k��5�����bق�H,5�GUu �	R��Kv.�S{��]�o*n�
9+m�ط`7�k6�YX*r�eH�6����l���ޫ;�%h册�x�K�b��xm��M�3#�p	��q�+'uR��u��$P���3|Nm񧼳�2.�)5}�A�d&�X��<sw�w���=��V^ibdvqt��+�;�zfZ����=jf>��ʘ��Ԥ��(�l٩Vv���4��E�� ���1c�� �ԜР����p�.D�Q:��+t��a�x��FL�l쫠5�W,c��� *JRf�`\"��ז����n!��`�q��7wLBfվ�����1��#W(�L�%��O�$x��78u�B�L�W�!+�;�e�"d��(����]$c����{eJȱ����qu^���:aI�D[[�̭9P%n�;�oEp�H��Lvr�	C� ��1A}�5����&�^����K�����u�-#��Sx��{�4[л��=�v���<��ݱJS\�Q�]����:g�iB�����0V�M�
֑�5��V֭`�xÚyn<��g.�M}X�=����(5hU1��wM�7'820 7�����C%7�K�is��>p��V�u�u�v�X�5�*��,]��Z�2����SB���ʎk���h۫{���\2V�ء$�<m�������8f�o���Y�fB�ֈ�@tܪ�n#��'�b����;����yk�d���4,����GF ���ʾ��B�T�$v!�*K�>,��TXB�b7���Λċ�כ���w�tNM";�K9KV�[)��H�o@�H��(*�غ�n�XGc�5�&���؃K�p������[u*�:%v��E���&4˰��L*�#yvS�DԞ1��f�U�:8��ڱv�˚c�qV��.{(��m�Ͷ����u6�*��]v��$��GQ��+c'h̆���U�v��H�"��A�k��^�"��̆���&$�-� r��M9��Iն)��5ӹ�x�yi7)�N򔌅Ћ`��� �[�.���<ѽ�,�G*��N�"T��M4��p�[Yhk���18����|���m�<�!n��eX9{����l�RK;���M������2��l�.�)�$��r�������:7Z��T��;u��n)]�sJ���6	�O���2v͵�Cs��eU]'�A��n�HެI��lq�t(�%r���#-Q�sW�*�7��|�E�8^���&�4�w�bv
�k�c+�l�9�ഁd�X�Cզ����q��uX8Vh�A�u�m���	��g��^�2g�޷n(�JՏ�0n�t�����Nh��sY6e�;�uҕ����ˀ��J�ڵ3�Jm�����K ْtBI�K�Yw��5����)dgv��}��/�h�XtGH{�E��u8^)�nf����͇PcV]<������[+��/��#��*Vc��LT�������; H�9��_v�3�ۮ���Jy�J���r��z�=��eW
t��/[v��t��u��έH7c�;�8AZ�%�;c��Xu��:/�4ovW��C2j��ub��s�=zp�@��K���n#���
>Z��S�h=�ͱ1�\�ط���]���3A�t�KM�Ƣy��ޫ��7����pQ����Q���8�ǉ�ʣԂ�(���y��h�mHh�Y�wU�!R�xd��Ǫ�%�����5��U����C��5�R���ڸ0��ˀ-�$�w��=Fg�L�W5�GC5�t�PWɆ�]�(�t�F���S-.xu�Nt���B���]�.����/b�Y���n6�*騱]ћ�X��U�K���|W
�	e-�L3�.Cc�f�	����GH����|;�qǐ`
͗����`�[+ѥ�d�KK2�g!W�{���)��݈5�JEY����AN���OV���鲞u����;��wXPF��xlګ�HBp�+*oe�\�rjR�U�$�mi��
�	wV!��9��fܚ�WL��C�V�տtQ�Ԏ�}|-�$���a���Xw����>V���om'd[
��u]H&]=�v�:�ǈ�*���F�B%�;9�&�vn�є�M�.�.��qu�uW��7�Z�:����.��4�4B��g�#
q��٬ͳ.�kX�u�%���ƭQSy�-NY����D8$;�+�dw�nڬ�T`tǶ��z��l�͛�t�A�N��ۭ)�R$/��&��y���³�)��\���ʥ���F�%ތ�S�j����֔95Ei��L���.K�ژ}Y�޼��}[nj�yg	\��tٺԠW6�������x.�0��zRU�#�a:r> :Jڳ��K��gu�d�����;I�H�ݛ�%RCcHsc�/1Pꊅ*sK���'H��:F��AYT��!UF�*���;>���W5�Ȟ���e��s@�u 8V[�D����a�r�GQ�'T��1��;����y���7)図��;�U�GrN_d#vR/-�ʙ�h;6�,Am�%'��u��H�G�Y�1��.��t��\70�]20�P���Hv��ԥ�6�J�:^�"�p\���\�8��Gd��Ka���֪�U2�.�U��]\�}�/�-b��oP}گ3Qv)-W˵�ݮ"�2�m�?}ӆ�A��84V&�� �z���h��y��5ֺ�����d=�چf�SB��GjU��5&^��{�,�(�1"�����0�AL|V�`v�0��f�]#�i����x屘�h�xB�&5u6�C��q��\�t�t�2o��`U>ޫ�bQ\ ]>��9��V՛ߗ<��&�[ۋ&��)\7z	�r����%�#0��=) ��n+fŹ�.>�-abˮ����ú�.����F���N�1��In�[�ǯyӣWY$�����Թ�Z^]��s���=�#})U��Ѳ�PZ��t&pк�����;7w&𔛙�%�p��t�k��ʘ�3n�G��B{a6H�6��%[ZyR��R٭]!֎��q�fGCz����1BaAc�Li�+;q��]�������١���a�h��[�������C#"K���C;��g	�p��,����^}#�rSlM��K�����
u�s��h�5sF��(u,ȃ����p{�q�����	�U�AB%h!�Ha�r�#�uQE�v�Ctr��M�h�w�a�.Sy�=w/hF-�q)*ٗA�x������}fM��V���(�ql�Y�#E�S���' D��0�����2^6�J�pnʉ�Zp(d&�&�����%c*�m��h��T3���΅����Û6��;.ڹ,��f�h�p�!b�m�wd�^�������ӛV�dK���μ�ݑL�F��l�{�Br<U%����N�C������u�\S���,m雍T�Wz�MaWe�FCӰ�b����2�i��ޠ��/pc0�+jC+t�ݕ��f:�o���b�ӫ� �8h��]"��FG�ōU���B�;V]����J����9Y��F'��T�/��@��s�# i���P[Q9Zlp�#oZ�����/�(��A�mh�k�����M]�E@9��ђ��Y);�]�1t���>�Ÿ��]}(��?��|��z�`�^�	>����`��T{'��@[��f�'(eg�����ڣ}�Uw����,|�f}�-��B��e���w�S�'{4��u"kB/nʘy���݉xݳ�:5�� 2�rwpӉ�Vﲈ�A�QM��c�#��vFk���}V)�dX#G1��'��uq9y�nP���ђ��g
ۍ���fr�s8D�c��:+������{j�e<0���Z��կ����V�䆵]���U:����Wmt'�I���>�wf��t�����;���S����s9�;����\s��ޢ71��P�'�ę:�������x)�Qfwi�i����j�]�m�Z���	�+���m�cBU�����x{������������>�{�����}�R����L�^AM�#
g��K�E���dPQ��������_�m��ik{�w�J�-�K[B�ls�X�OYǉ�9�X�VE�
�bp�zqb[��^FG't��[��� &h�B������L�%j�]�V�DEl="�S��pU��0q�Ag	�i]�IĨ˨;{����t���űu���%�G��-���5�E��f͎c'4�"���K,U�-�dj�|VlV7���g�Vw�"��N���vaU��2H(�ҮW,���	�/�tL+M��)v���g��N�s۝��U��k��X�_bz\5@^vWQB��B�?)��R�2�SLU�d�"�Wi���%���������n�[�hs�p-������D��[L�4�(v���;0���N�xn����2�B�z����s �ͦ(n��Mm��v��ss��"S�öZ�1Q��O�\������_t&���kj�=��d�W�aoh21�.��!|��h,촱,7���o>t3�=�d��3�6��@*�l�^o�ĩ��=���%��֭�R���x�:���Iq�!�s8O%�1z |��ېI۷j ���ZǮY�1�L�������d���T�L��c�ޛS*U�x2�n6��ĠB M��2nq樗��b��4�*��p$;��~�k ��%ٰ�QH�t(�%��4QM3��  �����W�͹�Kx�[�ĻxQg�^m�*�5T�1QU��؊��UIeԆ��(+C��64�kj��<~o������i�Ӊ�-�A5N�إ�ֵb��F�l�T�2h�A��QS��>>>>>>�"u[V��J(���F����(�6��͢6pV��ڶ��7�C�QQhìC��ƳMEu1SY؇VqQD���m��xxxxx�E4Q4ETy9('�65��c[d��"��+�5�nL��4�F,AN٢5�N��խ����p�mb�H��u�ƴQA$��Nն��h�h�h����6؇�6�Z�&�k&�N�*�kA�"LmV�m�j*�cU�j�PkQ�Չ�Nئ����ؚ�5Y���X��X�kh�ű;h�651��AqA�:�*�;c�(�m��9�c��h��[U�Ph�Nբg\�$ALns�ܸU-D�`���ns��3�f+��X˷US��u�w���\�����˝\���}H߇�5�����a:3|�EL٪��<��t�
��"`r��)���K��D {����UO�t�(��������R��tV�+P�tTC����ے{�t`���k�ڵ��(�񮌭����?/�{����P�x<�u�'0�n�m�E��vS9\Lz�n�����?F�yv}���:뻴Gwy�tjmK:Gq�g��/pSw��U���;>�G��n�~�n��	���h�5����8��v�w���y���!�������~}�|sݴ *�����6n!�P<�y����9�����ۖ;��u畘+�}���=�R��6y��=�����A�I� ��shA�h�����S��k(e����}M�\���/,���}&U	<�+�ON�5��Ev>�uvjɳ�n��bi�P��n���s����*Df��zM�;���%��g�\3���5�S��oM�;�����b�ȧ;�O(���Ӿ7^�7����VH��i�غX�q[I��$��n�����(��<��	V�G�sP6s�8i?�,Mb�ڕ�ߌ��@���������i�E^��u�w�Kz��7���c6�r�xΔ�1�9�jc��XY5���L��)��1��I�t�M�̇s=S�֍?���!V��Z�5�����O�~��I߶l����ٸc��~���C���EW5|�|)
�{�%]_����+�k��iёkO�3����v}�S76��f�uzO�1P䦰�z�-�9���J�U:���n��j��<}}�~4��}c�?A=�v�iroa�݉Vw��=��>��$�o�Y��*����|�q�G��N�~�{D	����Z���Z�w���uU��Z�xl��U=�*�F��y���z������"��uF[�����:��=��z�R���-y!��NGy�ʝ�:K�b�G,zSg��ڷ�������89���_�s�9㽒O�3�yd[�r��8��,�<�gXn�xb��߶a��뛙��9SV4�	���rn�	�������Rp[~��k�]�f�\[�˩�z��~��,_wV:�N�� -"�,.y{�� ڭ��cyѺ)F�!�d�:������s�:�eѐ���*Q�eī%]�K��ָ������=T�y�W�&r��L;�&�N;�\�U,^��>�pl���q9#�4û�gվ�O��nzo�==�x%���M����Iw6��3����Rn�z��h��/V��X�|��OOo��~v��ְ�\�zk\9yy����gԽ�^նG�8���'��a��=���SU�D^Õy^�נ�^�᲍�}y�GqV}q�4k1�oۺ����
�i+���tw]������^����ھ���x:�۳+�Q�i������܂.�������5�ܰOT�-	�wҥ�P�|�_}v-;�Z�J��}}y��\����ﲓ���5�j	���]*a���[?L��B�����������͊�����>����|��{�;�z�{}����2�Vz�6���T������&]�8��TS�:�Z�Gۢ����Xјn�e����g�z��0Y����6���9��L��\�}?9u*���S�]e�h}b������n�ǊG"����w�����X�P�v;�����_5�1���ۯy���uq&>�g���ժ\x��!^ֱ��:���9[���S�q����3�)���Ƴ�^�Ef�`�����εds4[�c���9�$ksns��΀��	z�4������'�-��M�d��O��t����Sg�{�&bs�}+P���JJ���3�Sȭ�ӏx�����X�*5r�����+.���s~/p�h�=���n�� �9��ɐ,�Ǫ�L�>�d�A�sKK͝�k�#�������缺��&�{x׻�M:�Z�vo��M	�����{�$��.�����\Ⱦ��3I��tO�GfD�CE�Н'*m���3b�;w^�{�ۙg���>�2�4��M�iOu�[O�/�n-�U����=������}R�H�yy���WH-��3���g����e�W�<%�[�ѫ�Lh�T�y8������7�z�Ѩ��/ɜ	�
��:A�c��<�>:J�~��~���Ƿ����Pײͩ�k���6��I�����5�X�z���=�fU<pԑyw��vם��O���U�6i9�|ã7ݻ{���=�a����5�#ܰ6��qC�31D�S�ޑ��Sh�0���Y&�{�I>�v�%��hX��xT� �R��לz$6�ht�A��ݜw��Fvַp�?ROl���v-e(fۍ6t@��9��k+M;3;5�A��$��n���ʹ륯����G���ӊ�b��e���ڶ�ܽ�ԙ�=sjӥ�B����c1t9^Y�z��^9ּo#�j%/u������W���y��W��T�9�6�����A��Oj�us|i��c+ٞ�awN��V�����t���ƞZ��b���`��܉��=�+ڗr��׉y��Z���Dg�]��u��~�@v��/�.rƖ���g���5�ͣ9w���}1��&.��sD����mY�h��{�������ﯷ/�H�j���@݃t7H;G$� s1�Eh��3��
�xj>U�K���� 2�+�M[8�O���(�H}����f���Ecg�k��^�km���z9w�V�>��So�{��J�[������$e�M��П���=�I��j?{�{�M�?K� �\}�+�;nq�0,Xqv�NF=pgH�v0�R�jl�2����c����X�^�ˎ9zq��XUx�ۻr\Z����7`F#J����U�rè8�Z�N9���\~W����+��|n|�+!�K#���9-J�:�L�yv3tüȳ�L�!�T�P���"����s4g�{����~s��y;Gw	7��-�<����m�Y�O������9�7��=�T��������I��	=/ϻڥGg�&{`E0�L�Z�s'B��W�����g�)w��a1 �9�o�u���ݗ�t1�̲g0�i"��y�ݬ�xDi���3��|��kH�/K��{��S/N��9��YV�����߲��2��:�M�6��sa��!yo���]%��Td�_�e
B���r�ӑ�9�}����#���r�<����w�9���p��X��g�M��s�ؑ��G��U�Ta�,�c^���n�m�bw���?O��9��J�*�+���ع�����FV/3������9ch��7A��Ce����G[e�xٳ3�q�գ�>�X�Kޔ���99fz��W��z����{��ԭ��'�	�Nɽ������Z�q�tG�(�7Z�c����o,��(�@;ƚ��ڭ�vSZ�0��0���݌�s�`�č�R�)�{;�Ǌ0f<rn�7�3I�딹S�[���͚b}7���j���Ffr�2�Kk6��#z���Wcm��"�w��e�[ɥW��z�����s�k�8}1���3ز����6D�9�Xm� �vU@n���3{�r>9�.����t�g_�'mR�{}���˗�w�}��נ}�a��/FP>r�3g����aJ{���}MЮ����U��]S��9{Q�r5Roa����Y���b��R����T����|�v�'���^Ne��9��<&$�>��{K>���ص�	����X����O+G���y�?`�����L�>�$Vn�GʹT�s��Sj��K((��2s<��<[�]sɜ���v��O	Fۮj�4�|N㴑R76D���3��4����n4�ma�}��.0p!7���>�<v+��Y�+�'{]Ui�U�Cw{/�$�}�r`e����	��Q���F��c���.��x��|��P�ѧ�΂���y����iE��}�F��tWm���t�ý�F��F8 �g�{ɼJ��&�^d��l|+a߼U-G���$��o��V��}��N�L�8�V;�gvj�XR�e�5���+zd�Jk�X��#.a-�o^�躯����̼��RM�������e.�z��:�{���u@�ˍ��W��`�J�.�j�＜�켒��z�m+σ�r��P���o�=���+��L�����n��/��FN�v	���DD~F�W�ݴ7_�����r��&���j������Y){�����[��궳Ь�+9��x��7�$��y-Ɂ�d�LEqw ~�%#^��{n��@�f����WT��X�)�+˒Nuڻ>��vr�4&��99G�f�;�,vCO��y�=��;��Ƚ�~]�깖MN�\f��n���v��;G2��ɦq�g�w����6yq��?T�%�[�j��߳�[���{'{����)���8��b��w��QR�<�֚��-��政�WJR~�߭�������D&���b�{�q��N��{�j�<@�����][��_JzR�Υ�AW��Ȼ���p�q딫r������ۄE�dJw)Ȭ�}���ɖ�s����=�h0v�Lu�&\�M���qwcR8�l�f��U���ƾ��֥�u���{K�>�`�����ɮ��1e�
#9_ngpfd��h��~/TOc�@$ܿh���f��}�(|�g���'��/����B�l������v﬊iC�l�7��mG��WD���O�������7jO{��7�랙�fѪ�'�N���4��������h\��j�==�=�C���'����g�	^C
��w�p�����1�GS;q��q�<Ĵ�2�����>r��nh�e�*�:=������Y���5���N�^�T�꩙�,`���@�-�|WwsclN����*;�x�d���㮡���B��ҕ��X.-S�ƶ��&����U��xL�7}��'���q� �1�Phl2��*�{}S){nz\���Ջ����$w'�1^sUy��_���g�|Α9(W��O�׻7��ZHg�GuG/�V���W�������j�~�;q^�kĳ����w��b��gv�y]���=�	fSsI|r��n�Ŧuu��O� 9[�$�9}99���t	B��h|�6����"C� ��W��3;�m�l��j0)�<i*z`Э�.�cE��M�zuFC��7�ԭ��c��������n��KHf��z��[>�~�#^�<�8`��j�j��6i*�[�=��B���$B��u���7���<�*5<�H��vb>Ǖs5�=���m�^o�z��7����K^��Ӿ���I� �p���O�4ѕ{����_�y���������K�W]7`�G�1Y��}�y��e�!в����o{/�}=(y��|�5=���҅�w��ݩ}��L�tn�Iڔ3���י���>�ϩ�HF�������4i{�"��Ookw�\��-fveX�H_���%Ճ�Oh�]�UE����d�]�hi�y��ng�����l��TI\v3�Ѭ��DX�5���V�Ӹj��6*�9�佗�lN�	*x�/nO���/*�z�}���HD�O�K{�=��������h�'u���|f#���'���߀\ݨP������{Ȟ�+�R�7:��a�u3��
Q��A�Zz�2:&�ٟ*B�݌�wb�xl�Fs:�ٍ�Aq縆zݾ�VšJ{}A�b-Ϟ���p5.�l��sY��4;{+�B�ڮ���Ul���0e*�wH���:��4�o��裧�s����=�QQ�1ڀ�x��1�J�*�S�!�I��5Jj<�0e��W5�uit
BvS�5�QY�4�=��:�B�c��@��Ø0���R�J�umoK�>ܒ]����}�nhB�W�IG^Qq�lAn�n����[��'S��@��e��c�ӑ�N�]��h���NN���L���ֻ�X���1���7S/�b��0��|-5���I���p�4!�gU���s�����NE7�7D�����;��Hq�-v�m�رD8'��i��F��|zvg1֯�@�S��T"�b`��7�H{4Fh^<��k�Q5zj�F�LKt�vTO-�r��5/�wU+n�� �&L��ۼo�p���Y���,�%��tȬc����,������޺�/���dE:8;���f��JBJS\��EY��t�ۮrv���D�;8�� ��pUݵ�ô�4�8��1�2,<�2�b����QX��eX˼�-��K�t�]�4�-���m2��H]ٛ��`i4�1I2蛆���Y�BT�ڝr3�X�*\H�6�-x�%ܻ��Y�v�q�Y[a�:����FG��1T���+NtS�I�����y���cr�
=�X���gTbqRa4{�V|/۠Vgtm�@m�>����<��͑��*���0i�y��.u�ٴA�b�XC�%EoC�s+��!ќ"s�h�\�v*GaSe��Ф��/�hA�G����O�v�U�oH�U%g��������f�ո�([��+{7S�z�\�Ю�>���ΐC䷣,H2h�,Gs�_G���έ]_����=Jb*�K�%+M���z�&�f��l$�xy�9Ҷ�#R������N�5�����n]�=��U�!�U�`���m$����)S=׊�.y�@9���d2DC�t7�DTM%�U��NUƭ�7*{� �܍%�˗���̤��Δ&�J�+79I3F���Hl3��Vf��g�Rv҆�yR��6�:��-���`�q:��%����uB2Cb���q��Ea��f�A^ۧ�sd���&��ݧ��hX��9{�K�����ӈ!�\���Ob�Ku3PvЮ����Wqt�qδ�'m枬��z��p2���r��3����:��4��ɽ9N�91�;�K��6��|�e���x�bF��wB�4�}:��V�!�8:©�&Uyܺ.}�,x�ֈ�|�X��1��7f�[]7#������Z ���܁1Y����0k���^D��eJQ�(�%3E�t-���%aN�|��Ne=�f��ݳ̋�u�,�˗�2��_YRU����b��! �T�G�*�-rW˕AUlns���sh�<*����v�9�D���f֌Ox��?M��&�������ޘ���tkS�IE<��消�.s�Es�&�&�nnnr��Q�3ǯ��|w�M�s��9�p6y�Z*�k[\������*ŷ#��(���#ɢ9�5�pṹ͊9�`�������+9���sA����À^DPyh�9��QQs��̘��9��n&LN���kh��<�y��sF�kQm���δ��ES��<<r�^s�j��\��r�pr�������lQ4[;T����Q�i�0sn[�&LbK��mQ�\v��dͳQ��EV��yX�MEU"�s�-�ˆ�p��Ӫ��h涪��[p-r�V#s[snl�M3���W#N�X���"d�#�-�l�3s��×#<ع���V�jۜ�E\.m[��r���M�9�gj��y�D\�\��M1���p�"k\�"`��;�,bkI����i��kC7-m�g�9�\�
{ݶ��`���sZq݈9j��4�sj�����J�s�w��ͬp�DA���`���v�\ڒ(�1D�.G�l��HD~I7�"@�w~��q$y�> �8����n�Re��5R���턶S�C6a��Z%h'fz� �W�p��#��/�Sљ�MT�����.dh�>�Y�{�VV��o�||�*V�D�1�W�1I�W����;y��+3�,�ѳ��a���ؤ��v������m"F0i�Si���:}1fzeYw��[)6��敒Q���'���)1���0��4������Ɲ��T��^F_�1�DKQ��:�MQ:�k���7s�&�:�X_�,��ii�1j.���[_WG�C��_d�:��^6n����A�gM��s����	g/IDV�Jfq��z�>c˕"�ѓLÎ/��pGDVgfOD[V�Dn���6��b�:%�ol��e|n��cL�v^�N��#*#�N�c��c&yK�n.��C�{�H3�o]�I�>�I�6�E6P*o,CX*rZ��ʨ4z1J�L�f�SSҖ��d�6;��[��Ћ��U�GѠ�I����Qi��"��V0֠	��r(pPd�9I��o$��'�W�g�` }�~���m~�����0}��Qϐ�PR�m<n ��w��xjv[����eE��ދ��w��ysЗ!����ɧo�]�nr�h�eK�Uj����Q9�ѿ
�f:��A{(�r;���l���kz�M���+4u���v1w��J��t�V�|S4�z�;.^�*��&&��q�Y�-�A��m�6Xy�H,9�JY�k\�v�i�5m>9WQ�̕l]l�X��p��␱&D����x�{Uo{4�r��ʓvx=�����t2T��eB`k���#XsPu�[+�~���T���P��25��m�]w�~�k_�w7�ok���L~�QC�#�P��P:*ז�Y�>}3Y�"���Y]٫$[4�]����-��])��[<О�l�≊�v�>����c0��pjv��5J5��T8d���.��R�4���}��2|��l�N9���p�=�`(�j	i������)!{�vUevoq����p�&D����%~�66=�oP��7�;<^=��@��@��qcg�
�FT_*��y��Dm3�/���@���"��A�x���N_�o7�~��3���aY�x^��J�VW �CY�,i+N��y0{N�dDʝa"&�)��m4xϷ"m�t���,�ܬՏ-T��g
���j��+�T�K!��?�|�jj���Й>�m8♅2ܽ�E>:��QGy�V��r@�z��x1�L�^�qB��w};7���#�T��Mh��8�V)��Hz՗P-
���Y��7:W=��-z"�해*5�5%�;�ظtT7�� ��đW�aոs:�[���a��VV�;�~o�Q��};ݖ��3��������E �*顶#�:ʳ�(-nZܻk@�1Z̩�Sڛ&)�.�."�ڒ:���_F� y��NQ����.ͱB��_P|q{�"�Y[�)�h�~N�5C^�����r[G:e�K"�탻B�Ҭא�R������U����G=J���.ǃ����Y�hE�(O�[��Vh�?}�w�~AF�īȮ2�Kd�+�O�c�g+7[��聖�,�`AT1�]�m�5ߜg��Ǒ.C.��h�3N�^b���9�/�y9�vn����?h��W�PڟK��q��`&�Ƽ}��_��Пg\����9s���Vs�o���]x:ԩ0�r�MED(�L�?O6�JV�ˋK͖� ��@B�ﶱis���[��Dԡ�=�G���4e��\���^s<�qC[>� _�����jBV���̸k�,���1SZ��{jf
su��ƅ`%R����j;�e���Za��-g�k/��ދ���Y;9x�S��C
D�}�[��@C���h�����璓-G5�]����l%�^7��U�a�K���*�{���0mx�����L0���dƺ�s1z��rn��U�Nާ�'Z:Է?G'�k��UO����P��w��K�@��3�y��d8����&��a6Rw��B�Կ���,о�;�3%(�b��f�%4<i�������$�poY��i�J���3�\�]\�F.�z�!��^���ŧ9X�k9F��Ά�M爐�KٸwD�3��x��u�a�z���f�;Lm�l�Wջ\�?oz��u�聚άq�Y������Y/P�j����s���g�I��=N�F;���~��݇{-�j�-C��m��^�D�^�$`*)�#Ο���T��qG�߽r�yG�N�$Y�Qܩ	���`c�)�ڦ��/a1���0f�B^��p���w	��Uj8���Wf���7�N܀�`<Z����u��u�]��0�DҞ�&W�WB��UZ��\秱��"�)�3Z����ٵ��F�F%f��ޖh4:��c�Ls�ǹ����9�,ƪ��s�E�Fq�3�C�����?u�^P��Ե�o�4b&���9.�^
A��M�[�7��P�����m�3��N0@i�M��e�?���]W�:��2�9����N[�dc2os9��\^��Z�׹G��B��r�h�ן�S��y��*��A�ү���Ƙ�b�k}�'�޽��5ۻ������m�	�Շ(=v�.-R���E'�\���JV�5�*�|=��OK/)�C_/)�;����c>㙌kCy3k���,g݊���LH��%W'N���?�nk�>��{��-�,��<<�2������V��ي�+Pyk�Wqʏ0�ʱ��#GL-��7ɛ��M%c(;K�ò�.g �CK�d' �[���:�]���ه��p�+�.��d��w#�k�);���Ҵt���<}\��V����s�_	UA	Ӥ횲�Eц�C_�s�θP���L�	��4�Sm��V[5)3�X�aE�&7C��3����:�vS*n�~�|`σQߐ'x���]�)���ʄS������|���{�m����]�.g^׵Ԧ��>f�&�
�A��0nc ��L���E�]���J$[4�f��w8���I�Z�eQ��=��"��0e���'%��Ũ��ݛBr�n��ߦ)wF��&�i�������W
�򥑗��u�1�Ӊ@��{�U�׋�a���3H�(m�wm�W۝�a��M3�Қ��#���f�{��t������9���L6�R�
�����P�:��	�!7,VY)$��쿡�T$��5�/'�љyw-�a�
�'/!qi�O�7j9���-���0�;���M?n�H�"�;�ʦ��uq6�k��>���J�����tt����Ǆ
�fנ���z��jط�q>Ƅ�T2�N��	��������֌��Pۅ��lef�@�v:�!�AdK&�	mSm�-�k�j������$S�LW����	�ʗu�:��ך�m�g�@ݩ���D�E�-���iKL{�R�%c��1��8�UU�bw2���I�R��ӴŬ�1-�SEp�����2��L��ۛ�3�ey+�u��|�C�Y�h[}x8�o��.YY7�-ޅ�Ȯ��
���#º/���9R���/_t��q�0�N��tI����@��{�T�l�{6�E�B<��Yr&�!-�]��Dį 2�����dn�6:���}�6�R�T_�j�m��5�,�����&���̉{lV�F#����L�Q|K{I`�lTs4vuC;H�J�[���M��n����2>/�1):��r�!�y-��]C	<�/��1��x\��%ȇ�vM>��i��*����<iW!qu[d_u<-��j�tߡ@�A.��;�y����X�/�~������v�g�ɿ]E�TT��N�e'(��=��Πmp�E�O���t�����N�N5$��`��@��8��y=	����9�n��K��qe�(��L6����P����3\�<�+�.�wb��y�Oe����I�df"���C�ˬz/>&�P���q��j��h�V���_�<we�w��/F��
>H��W����$:�8�àor�K�nH�/4�\d��O֖��~�]~�CgI��͕��	�-\_�7�SQ�`z��|~�d'�o~?I���r�}"�����@_��Ѫ�`�X��&PTJ*��y]��\A��Õip��C[pхP������^�2��4+������C3\ul�d��2�H��n��D*�̻�K9�\�;�䙋�
4�'˻���w�C��:���@��]�es0���}]ɓ��}s�A|�.--�ST>����H�;=�b�?����Гɻu/��=y�m~.�[�� ��k��Y�������]�9�kP뉇��Y-�(����V��nn-o��w�Em���e$�8s��׊�h#!ľP��y�7 uC��h�2����ɬF�vO[ޡj#��������S	��4��s��B������Fm���,�����+e�b��]��j��ͦ��6�1�Yտ���w��>�ƷW��Scz��˞��'�[�/c�s��#"Ԛ���VDb�q�Î����ȯC���oi�.��r�ċp5ژbٱ���
Sb��H��y���6�4���aX���G3(m�q��|mw���K���K�˨d�;�k�EN$Q�5wٹ��,�y�.�]3+�`O�<�Sp"�d@�}y�hņ�G�5�<}��\���z+��xٯ�7�t�s�,��O!�÷U��LSߔT�	�y�9����hCs,D�Oh�M��6�� ����B�0�Z �o�yOъ$V2a���E��6�*�a�y���QIǞr�}�.��*�5�A���T55��,��� ��s��Y��̛��Y�'��O��Ԑj�e/�e/ga�#�uR�oڐd����J�U������]�� )�+K*�����4-�`Ỉ���0��ђR�E1������D	�]����R��#�T�w`9�[&as��y�aR��PY�	�s��T�<�7m�y�u���1{�l�*_�1s`@1��-��u�S1���S)�eu��uP�J@�ȋ��ٵ}u�VԮr�P�لY���xW�ܐ+��"O�|�`~ A����1�ԫ����'�5�s�;sO8^*5���}z5Rf4!�����4u5�rlϕD|��h�xsҫ�0�Z��rxR�ց�j�DA���,�ĉ�P��TP^��_�f�!�5��|D�^�'%�긺b$���]���fD`�}�X����;���zY #6Ξ�a��n^(�4ͳ��I�Ç6&C�;�o�F���	]�g���զ�팻V�1�>* !��!"g5V;������Z����VNг�̏lhߩd���*leO�\sS�M7�R�kl�q�*Ԅ�VY�RzPb�1g���&8]�����OQ�f_/b���Rd��k�>t6J�Cz��>-=Ҩl���Q�����\�n|]oے:�Ϯ�ԉ�W\3'�.�*�	#&|p�Jyq��/I�1�WE��"�S�1��9�re����Ƽ1Dh�n=�����1��9�l��@�)![c6��#�Z���T�y����t�;N�	�mC��y��;�+���b.�3pU�0���7[��*;$�\/so'_F�KV�:��6���~�;�^�f� �1)�{T�e�
�d\�	�cT�E����D	��FQ���nߞ\��j^����:럃g�b�,cz�=���������t�R��|y4�����]Q�q�9~Y&b������[�S��z��@��<�EŹ�E>(�����y?6�
�Z�1�vi�6�W�uhB��>���x�O�Ra���D�Tn����#|J�O� �ꫮ�Ȫ���C�޶����zX(JC��}K���,cj2��m��F����}���T4��B���ߨ�J�vںi���k��?���F|�;�B��A)�e���GN]����}v<T������h��˵m�@�-�@Z�3T�%�޷�y�v�H�͆�t_g�@̘})N�U�0���iy�X��vh-��mΙ���=�Ͼɐ�f'āP���\�C6��%�o�4ٔ.�M��z���\�C��Xk:$����F�+��߹܎=CE}%|�ʁD�mAem�g�ۻ���pr�Ey����ckCO��KT�£�fSy����i����C����V��5@�5��WV��tqԩ�PEgt͞S�_^��.�^���M�f!�6��ڦ�'v�1'm�i-H5�mv
�d�.��/���|Ѣ��P�Z/8�P���c1�ծD�x-r�FG*�+���={J��.�B_p�8n�,5����%lC��a�[�{a�0�P �t���.����g������U��2<p�I{�e��|:�$y�ƌӕ<l�.(.�Fݔ�f÷,.�v&i¦_�-ڝ��7�EpW�x��Pxv�J�3�~���=��4�mx��R���Ք��&i�)��R-�����z�^n46bQ}�\�]��Ѩ
}�Κ�~b1�,�-�m������9"�2�f�|+`�)�����j��Q����M��o��p���>Fm:́
�OZ�cm9����r=t9���j3u~�B���B�t����������0/A��&�|�Qi��T/}\e��M���t��y�̋>߮dT7X��
�,>�8mc����Kz�\���=Ӧ�rZ�D�eu^[5��V&��}��5��As�Y#��e�jހ�0���:ױ.Cs[g��Esö��8X����Yڃ^��{�<:�t��YmmF�7�F˰ēdYp���q��f&-�+C�^A���-ll�Ygo_a�^:�SWd�4�jB���ڽ�����t�P�$vd�ฃ����#�X�e\.��L����ާ�۱)l��X�3��>�Y�o9�d�ec"�֤��q)|NBke�I���?��	��+q��c���bȎoMö	��!PU����#+�1PWI�&٫+�����Gv��#.��Ӣ�ݧ0j�Hp5xgV��ʛ��]�g%M
r�b��A@���lİ�3F1#��f��K�ɣs-v�����}x7HŰ�mU	�h)�kj�%J�ʬy�-�Ve�iL޽�j��%��N0�oo�e�*u�jU�-%Y���i�.� A�|�c����je9�ɺ��n1j�v�D�QCnH�T���A���F�u9c�7j�Y�%oj�j�Sx��Ő�Q�J*��m.F�h�������^�Y8j���XQ�+�!=��+/�֋s3�*'�u�#�yP꾑�xB{F�4*�fT�08���mr
EB��|^rc$;.��B�r�[@���Ԇ9����C)l��R����@W�Nf��{�������yԚ��[CQ�5}.YF�} -�5��klKu2���w�z�󐰊�%CJ�8t�X3�5�:o&�p8.�H�;Dp�i6V�Əf���i�[Y�,�����؊��n��!����3SU�6�+�Vs\��H_'�hOX�Fi�1��C�d^�9���:�D@p޶�㬿�i�TI+1w5+V�&:���F�2�K<+p*�]  ���R���������3@]9��-�j�v�B�kh���6��7/����|��ID"�J�[8p��U�7ƅX����}Ͻ��Q��Z��=�@�I�ȋ��6�C�ky��LE'������)Z�K�z�Μ�.��
��Y���&t�i�����-���*�Z�Y<����A4�8�N��,��5��iꋝi�k9��;(�Z�0�;Ύ��r�;qѰ���'[�α#X6{��e�5�&_l�*�C�;�mᆜ�<��,�d��3H'�3����ݳb����W_�dnTξ���-���s���V��]�0S�6�sR�/������b\�5��Bد*�4	����d.�yak"͸��v�wd&�;[������G��DkvѬ���2�Bz�C���٪��M�^|�j��huN̦���R�I��z��@�n�n^w��Q�kwE�-Q[}��u�Mi���;X���.T#���$�F޸n!�I�q(�:fq��:��V)�i9[f��yg�se_�j�a���ݙ�T�/5��<u�@ҹ�Y�ZX�M� �*{ʥW,��F]�C��kF$7I9�L3I���f3$���]w�C�>�O2���T��Ҫ����U�Xi���}m�?��c#xX�T�B���lu�4ܧ����q�5��8+iB�a���)�L�b21�nU�Y�aNv�[Se�K][��w%�+�Q�b�*�oE n�V���5eS�XZ�i͕��6MO3�rкۙ.К,����N\��F���`���G*c���'D�����-'Y�5�#T]	��RG( Ml(�Z��a��.��]o�.\��S���W�yȦ��.ڢ6ڈ3Zӧ4F�֚J9��O�����5�^ZӢ�Ɗ"i툍�ݬ�$�#�͢*��QDEh�m�CD�D����8������<��(���8Z�O6����A���J��FgZMh���<�DUF�ZME�j��mZ���7.���M$�"�f�"��b*�" �N �l���%�b+lj�*{�PT�M1U�������Th�#S������EW1�6�D�m�����TQQE���-j�������(�������U5�$�AO6� ��76i��D��֜�1LE�TE��h�5lNت-kmT�ULLJTP�Tm�F �4j�*��(�#d�4k{�TU%UDT��PTE1�]�
c��6�D�T�]ت���y�D��&��A����~����u��8e�������Ƌ+k����Js���Aan����bv������Ԥ*wCp<dvc��"D���C�=���7 ;T�	y�I�O`�I��[<О�l�옞c�`�����C�%կ��w����~�����N��_.,�g�qW���P��}(o�ԮE�-�����v��d���mꭷ�KE��j�D,4L��E�/i֛�P����V9��ͱş)�h�-D��jy���'v=���B��F'K}_�`�ay�Xz��ެ���_TݯQX���bf��}���,�W-w(k�bP7�����ǖ��nl,��j����M"n�y0���%�:sPw]���]o�0�x��!�C�*6�,�͞J�;���/Ɔ�hU%�;���?k���]�`~-�&+�����֮�K�qmWp��z�1�⌠�\t>h�8��E4�����I�Ы�}�ˑ�ٹ��M�����*�{Z�X�ԥ�DL���X΄C�]�t��l���5�)��ه�7�ݸw()~f]����j4�l�8ZΔr�J�ۯq����\z�R~W�<��8���z���n��B�Y�.��jKƏ�E����fa�,?�P���X�M:V��e� ���Q�Fl�5�Yu�־\���YJ�N'x���Fm��;�s��J& ޜ�5�.�o��L�;5��vƳ�}[����������ql��[�IݰFN��%;�׆��n��0�ou�q!)x��z�]���R�A5}4�ug3�Ku�{�Y��FW��~ 5wbEʌɵ���F|��B���Y�B�gT[��+HAp�j�uJ���"�٥��֮hW��q��9��(3)�4i�9N�x�<��O�B�v6U�ss];:����-�Q��t"����N;l�[z'���~�)����:y�ˏ�-֣��e�uM�cg]�;��^�:���j`s"�1�{uE�a��(�\��2Y,f9ÌP�ϭCF,�Ʀyj�N������E{�Bͽ>����O��v����b�J_����G�B��_b]پ��z���ڧWbõ��T��HT�z.��(�מ��}{rϫ����?Y$�3��妕]{x�c��1�u��F�$�g��UM�\cyN�����ʐ���7�r����Owa��r���gf�î!k-�6\X���s>��-NlD~�	ߖ������6g���{ҾS����YZz�ാ�C�23u_5����n�0�A,���!��h�T��\�����lD{k$9��
����5vW�\J1
���~
n)!���߀���������*m�#ΟG�tS-x-)�_"oI�o�!�.f��G7Ϻ�o�b�2	^�G!t�rb�������~������pI���l���2�C:����]Ï�R� y�巖����;7n���C4�����SpЋ�y�SǸ�0�H�˘e��o�IM.��ƍ΁s������7��sQ���Y��1�Ĕlb�-���T�cȬ���lм�,a� پ�$Iv�V6Rx�n�2w��;���(�Y�9���|�����.9���1������	�{�,��@f��N�yg#ƥ�D5��P�9[�	7XX!Pa�w�>���_Q��*��P ��8��SS%�or����嬼�YY��S��_tԉ��e&��V�R!�'����O��[��4����ǒY�l��p9�'�`Bw�J��9��m�eM�q�2�'`X}�S����/��	��������Nĉ�����}�@�Ty��$�a`���ܕ[m�[�6�^	{�X݆������.�n5��Cj�LvK��zP��^�	��y���J*�)��"�����9����p�q!N��v.���G��b�f��!{�:����Eı�S� �<���7#��,T՝�q=.�_u���F75x�>��cp�I�!�G�0#~;���;���+Y��b�:�kq'n�kX�j����|{�����������z�s=>�S�h/��qL��=�2��4��Le�ֺX����i�ː����R��������z1�~� �f���W[�nv��-�}V2>AJ,�ú�8�n�}U��ٮfqH��@�wֹ�t��ݨ�\}�'�@�.�=�6�gm<�N��w����0J�����A�`�2�Ե%����S}ҍ[^���b�-6���3�CKd�71���~2,b����
���n��5N��>��z���N��B��<~�Ǡ��p�*�8ۿ5�bv6�{#�c�F�Tk\p��3Jf���c!��Bz0�v�J�P��s#��&gK�����f���S�D�Z��P�/�v���͐�hi��ZaQ՚��2�I4��{(m��m
��|��{P���Z��AS|��6L,Q�Ҳ�&4�N&-�y3�^[6)�ŋ�uP�3��_|A���s��6-�.�|�U�s�,���8ޘnX]+�b6�;���*��u��ɕ6]A ���]'o��CQ���c�2xJ2r�%������iLϊ�Q�UI����|������\��ք�!0����ޅZ�΃&V�Ű��M�l�U{�<5�nQV(lE"�F����G3��<,mX r�2�%;5���B`��x:���s���l	k���1	�����Ԏ���9��%��e�^2;0z�BS!�tn)��dHW�'�C��Z�='�p��.�)�t�K���C*�*��7�=4�qR�*A@>n�+�R^ߝY(��I^>w3��BoC�\�$h���D^Μ�����V*��w�!шoR�K3+����Euyjw�/�<�c/�TΚﲳ9H�9������:Kk����6R�����wz�!�����3y���=[�t�W���%��U�P*�1�����y?���,���^���o;�%���l	�Էgss� ��E;�&����hu�WBA���&q��K��K�Ť[�&��T�����T�e�+��E2vGR�j�r��O�b�tkey#�ȁ��#M���-���M�}�7<�v�MVT*��B�I}ݠ�[As�|r�4�����q��=�I#o�k�B��S;'����WfX(�%ᠺ/����8ȢT���r5���="f���>3�+�͙L�Ef�>W^d�=�aJNOm)�y���q�cx(2jF�z"�R)�{ �ubfx��K�-����]�>�r �$���
y#j�>,b���#T��U��{��L���2�f��?�GOc��Z�FK�j�\���{�.�5�\�m8���LM:��I��pw�1�p^�vD�7��ź/�/��8��Ԯ=������;���Pmg+�bt�Jhְf�1�r�FҍY�w3�}�~�X�Bi�^�{���)���ˣ-��3ڄ���v[����j�l�GmҶ�v���#������ܹ���T�[g!;�0�L�vh��Gáb���hT%�ݎ�:\%P�:�{:�5�fn���k��[�j-���ؕ�:����v�VY폦l\�I�z-=QPBM�)���P�C�TS 0`<<z{L�i����ޛ��B^�ŵ�d��uUC����&,7%�oKI@;��g�u���}��緎��V����Ϻ
���le�O�[P����vs�y���W>޸q`��X�O�ʹ<_>��e*nr�vl;2|�v<�/E0��؝(qͼ�S����~4gٍǱ^f�>7����[��WuQ�{H�Ҧ��o�mC	��;j��oi��l�H8�[�h�)�,�,�4?E=R TZ�VOL\vUb�^s2�tjQ��F+���F�啲���%�#$$����2ݮ�J➢��]����!
��6��^~�)��Ly�
�l�f�!Ҧ�#|\�S��1��u*�u��i��ǰ���{}wjPK=�jg��^�<�g��e0�MJb�������m ��p���n���Dqc�f�[�j�s��O�ɾl�����&����֠l���L�7Ju�d�X�0�r
w�:�NNu^�.<YV|5b�N|�c�_���#�#b�}ӜhQ*T��[�	��U\�L+z�u��8��#�W8Č�	�<�=J�BQ5�
�A�� ���k�=^����(��sZ���!�(P�Ʃ�n��΀��W��z�9%�l̮���u_Zє��������5�xvVGׅ&���f{w�\���o	g�k |��F��v�y��Gl_o`.h��[�{*�U2�7����W�QJu�5�ܹ(C��e�����;(w��||z���^���C�`I��!V�=ڎq�c�������)Q�i���̶6���_�������*_����_yh��u�Ř'�~w��Ւ}��VWV�[8��-/�q�m�3[ؗc^�JD�=�Il��$��9�V�TVƮwm~a"����֯2#Y��xY�q���L�cP���,��i�+D�u]%��*$�'	��;.�ؼԤD�ِ����W	Z�t�W6��b���4V��Z��SӦjq�Iՙ����o�̭�] cZ�M����F��0⿭�Ň�vB��0�T ڤt=��7%�%Iv�8��ΊH'͘c��m�3�pV��#b���,
��VOz�1q��l�~�}�B��a��R5���cެi5�*!��,��0@;�b#\���~�ǒݨjme	[ڵ�sp�5/@r�Xפ�'��:�Ϯ�ԉ��e&�^�k�J�?�PZ�Kδ�Ξ���Qy5�i�Ok��q����;����UL�����e[
*-���V���M@��,��Г����!��X�����J���D�L,����i^4�Y'_��}ƛ��.�z����@�M3�U�ݲ��(�>}�2#����UL���s�yoE?��ԶJ'�4��.Y��2ui`3�ד>ږ�\�������{u%��lep
�})� �[���j����z��b�D�G�'B����f���*<���)$��**� A�Y�����!KL�����M����Z��[��l�ay�Ɣ��RSڈ�*�L�#���[�~�u��>�m�Q��{����XFAM�Ir�!񍬁Q,z1T��%�Fc�jv�(M\?I����r�-�#��t�N������q��{Ȥ����]�}B'�Fߎ�����{ݜ�[�:�k��Z��^��+q��}�9�l:r݈\�m `3O��<�����=���U�L�1ə��7�{�r���ˮ7��y>�g�3�i��Z��[%�}���`�����3D�ϼ>x#�mpBUB���P����01��UV��������f'��nYܳ�ge]2�V��^������+@4��� k��O�����T:�s:Ú�Fzz��:���E�U�v�Wwh~�6h�b�;	9#/k$)�~0���_�v1��ﻨ;i=������'��pk��7o�d�Z�zH�םACl���+.cN
�LY(M�Q�n�G���60�̘Y�����{*v��$6�2�1�.Y�˰M<��h���ILQv����XG��FO�����6�	]KB�eS�i���Mg�����A��
�=v���.k�t�p�<i�����t)8�hӸn
z�&��o�_�!`׏s��&z�jX�y���gfutw�7CW��Ǥ���Q���Jb��|���|���#c_h�h�B��%�
_<�������������ǟ!�[����;���:��ת��'�*S6��3��}P�q�ҙ�b��R5K�hv74sd1ttu�Wn1IB�!Ƨ���ǻ�U��B��ȖM�䶩���ֵꋇ�t���Y�m�LS�8�V��q�h�&9��[�RF;�ii�q����4r�]��ge��O�9i+�T��fR�ʍd�:�V���-�/Z��̍�^���1L�mPK����Z��U05$�P:�z;��O~�<����c��~���e ��}4�@��k�s4nuC;jGs	�stW]d�r֛3�usC��Z��/ݪA����jD6 ����u��xE�z]-<x(}��XW]�oV�B��C1;zY�t[gu�.���ݞ�8cq�$v�����������w4*�5T��n�b�q]5�R���f�8~N2��j�a�/G.SJ{,���ZN�\�$tKX�;���M����!��������%�n/��dU*���ͩ�ly�A3\�B�Zs�T䬼1g��<��e[�����{��t2��S�P:x��/ө��F�6srC[�0V�����ڝ�j�2�K[�y��G��Z���u����''V���JVԶ����n�b�}5�orMs{��{ʱ�=\Q����W������V[�ջj9�&}����J��:�JX�7d��	�s��bJ�n�[�8淃�C+�����&�V%
PV�>������������55�����v��͓�ϼ�����X�r=�}��e��r�����4b�<w�O��m�.(t�i�\�oԋS^a��*�����A�W���̯Ѧ�O���������𼭂ru5j[�L�[��c�ZJ��e�8�v�=x%f��n&�w���V!5�^�?�3f~���pLg���/��>J��r��\�mQ]�U$bf�&^�Wjޖ|@F:jEק�W=	zǖ��2��.����>�6�FD�P�6��=�'4vTe'�<l�#u�L<2ڇ�T�l������֕�A�zz�_���,��]ې��2�MT��n�n}����;=�WF��]>�����p%U���,��������DB���h��U�[���٭���讛NpnH��Uaqv6{n���O	���Ϳ��g����O:n���[�g���jz�1o��3�A����x��&�X�zY�Coܲ�_]ĳS�*ݳ�m�Q�;[��k��n�)9�eVd3H��\�����1�8T�eY�{F�f,C�=��z����O3*{����'�d=�����kU�[���`z���uA�hT��A�L� �<{�����@������x�\$�r�k�#����-&�Ⴧ�Pw8����9���&���YN�n�3'"�jd[NY�*��U�9���#,��ns�kv"�&.w4��^m:Z�s��$�7��+-hsjM+��K�ƷP%�r6s��ּ�����ǹIElǘ�X5��7Sn�>g�f0�9�{����gT�����Q�:��#{ow:��}�Di�ѹP�N��<xٗߌuQ��l�."a#��uz�$xQ�B�ꮡ�8�X�ܱ+&Y�rbf5@���L����7Y��Z'p�D��;gX���y���[|��^�����b�Xƞ�&��D��_</�'it�k��m�b�:����[�nb�-|���Lk��H���O`ˢ���wv��ت�뽀qk%+��-C���Y��w�M�H�
�{C�)�� �Sd���b�ҭ��7�SY} `�*A����4l祒���=,�ZKBqc�7�v����ް���`z�:��r0���:�dkcy�4𺻜h���{�]a��Z:%��"�xXt��:��A�0�CԳl�޽;v��"m��F..�i��+@Vv/�������A �b�h�)����f�t4��{�P�םϮ=�os-��NTt�[z���.��s��s3]�x&�J��;�m�E�2�]lZ�Vf=ID��t����wC�' �k|�;r�����RU
w� ��t��I̗��w/O{Z��˚��©��������[�²7Q�N�6�:��t�ZwYT�PL���i:���8N�ۺ�&�ݛƥ#��Y1�1�7NY���:*���&�F����S�J�	�cX�I�X�z/5��|k�Xa)ú��Xm'��E�p@B��-hd��5�sG�\��z���f��լ-jt�\�)��J�oI�z�c}��Ĕ�i��DG��M�y���������y��
����%���V^}���FC��E���pWJ��yKS���c��l1-��{%d�j�uё�Θv2�Bb��VӮ��(�]M�6{�R<�V��:���l��wm�ս�L�e\���+�y��%HZE�{a��Yd�c`��/Q̈�\����-���;�%q���sN`{���xF��&�O��O��l;�v�I/_L}ټ��b�s�]���b�Z�:�nt<����"P�j��|Lߐ[ڢuq���aR��{��4Cn����1�Z��y�C���[�W&� �BLkm�j�.�c�0<+�3{qT��	��ٴ ��O���Y�nY�զ�����_�	O����ͺ��0�lY���_�j�&�򄅕��l�An��!����q�h���mM�m���*(���J"�d�&6l�f���>>>4xAUDQPQ$SW�5DA%]�*�����#sfbN�|||||/^n�G,TD�F�0L�MUS��b ���n�����oF8t����UI��ִ�QALML����f�H�j����E54�������(��`��R&�H��E�f�Z���F�X �(���*"#F�ff���#s�&"*(������8S��QA�QTL�V�$UD�1A������6�"(��5Eh�4�8���kEچ(�)�"��֢�b��*�5EDL�A$U3��k�F�W6"�j�cSUSh���""*b�(�:��\��*���B�P��~=d�f����o��kɷ�E;�3T���gWB ��< ��s1����K��5(5إ���ċ���ڼ4ے������}|ҁ2��Ш�_=�=�u��߂�Կ��z�0�v��׆�cɊt�	��~�m�T�p�^�A1t��*���9Qx[��\��T&l=�&�`&���y��y]�hӋ Ҟa@��nZ�n�X'��bg6oqV1��Dw���Zc-�	��E����k2�s/���6,�*\b�s��$�t�Ot֘�^J7�e�����SN�`���$o��32y�ɘ���ʹXhd�g���tkv�H�3J��J�cs��z��tj���q�h/E�7�� �`<h���/y�L��<�o�j��;p%ST��dƺ�sW��q~&5�����j��6%��@f��!�\��.���j�����x\����U�K
�A���\��J��,����;P]&�7,G��4��ߝ#��/x3�|ʥ����;��9�Sߵ�\fd;^���`��oƭfm�����z��p���|R������C�Z��7����g�b�Jw�9Xpu��ŇSW����s|�O~�)��W ���֌�CR�T��k�z({�\~9;���:�Q��>�U!Ơ�(���%w��`,� ��C���ݣw.�&��oN�z���묾O75w����\
��ѝ}�k'�b�i�ٵ"�j�S=*q�.�%k'��A{Ӡ�pV��C=
��]��܈ᠿ����/M��!�.Ǻ���
`to�3��{���7�_??�|��ߐ(~P �	�D�-""���x��{���+��8�֏�eP>Np	�&*�0Ug��_�J͓�tQ
���X%pɥQ�kN]]�o1���C������~��L��ַ��W�/LC�8��	��\�Ks��_����Ùq�!��j:$��L���<��]6ڲ���sj���.�����z/9;��7.�B`&���5����Vi�s�t�QU)���l�򄢱9֠˲z���뼹��D�YȫP�A+4z#��G	M�P@�/!��.,9�E=�s>�4�5Wز!�V���,�^���7X�=����c�T\��$�}~Zjs:���,{uT��A�!�[��Ք�Ke���OaD���^�����}��|WZ�Iq���z0P&8�R����3Cr`�R�TZ��R�e�6��f����'zƂ{�U��Ǫ��g��5{�8�5tB�:~Vc��5���vr����*�y�j�j���ñ.����0݈d��߳�W�W�ϕT
��LO*�%�V�_y]��R�1;��;z>ۅ`�Ŏ��1��}���7�͗N��g�e@���>Z��V��A�44���g��*7-ᖅ-���{��] �b���x2���4 �7b����s�t���%��
��voiT�u
�b�Oo*��.P�*���U��u9�Sj�,[g/k_U��d��`�{�ܫ]���P�K �_濑?&I�B%@�� ������� ��n�a�Ct[�grߜ�c�d��\DWZ��j�}�ASk�����nn �}ZlpT�ql�f%��������ҫƂ�`�&��z�d�.Z�|��X�mEeC���v~�8Zy�8Į�wnc��/4�9Ԅܥ���<�[�V'J��&4�N&-�y`��c�_�e������pUc��^�:�i�1{��Bt1��v����<����W*K}A15@1G��ut:���׽�ʚ�S�V�MG��_Mc��>��ב��;U�cޢ6�����0+�b����N�����Ҡ�k��]������s�4��`a{���j%k��A�O�Ĳl�;T�`��k���0���D��.;���g=l�5�z�@4RF�>z��-�%n'�֧���V�DI*��wE��V��z�"ڐJo��Iȭk}�c5�����}%K����7(E�%3!�B�>L��Q�7��ב�NNx�c&�kI7&^���]x�N���}"2:��;'/�S�1���չ����iC;,)W5��T_�EP1��*�Ab��P3�oA��x�����~p�;�w���sr �R��[�ظ���Z�껔}b���ϛ��}�-�;k��W���r.lŵ�ZV��͐��WU$Ų�v.�ᤣ��a�\)ǙHh�\���6,m�&�3%����i�
���<��G����o^��P�E�� "i!Z�R�J�{���E+-�ePhkgno��˷g)�&�s�������tke��6�䓇�k"������s���Id��f�R�qԀ�ζ�R'��@���&^�r�4��
2Yn3�A��.��F��U�����`i���В2������
�VA{/T�V���4,�)��y�=[>{��/F[O8���.��l�e�7���a,%�|P;�������6�?N��B�"�g(�詞�|�e��
��"�n5������	l
�N�C)-R��G�'��C*{US�w3�u�!���(��{9���Qq�lE>|b[����ly�V��=����{��D2˾�[Y�X�����W�̛�v}�礮q�Rp7\���/����1:W�2�ǰ��3������%.�Y�⌱v}��������P����}�F3O���y�7�����x�e,��.i����f����Gy~�]���u"��3����1����򠌉lkv{��{���|����!O:K�^Y1w��T���l�����b�S�V�"�ޞ�y������s�CX8���#�C���x<�h��i�n�����;�P�z���{j���)�����}**���{90w_Q5�4/;zw|�=��{�l|�-O��$�Tl�i�RX̲��zUK���ҽ�-�1[��˾���.�����3����[�P3L�fD�2�>>|���!��Be`V%�`����� 3 7�QM�l��������zY�/�S��^���+�_���^_yfF��]<o��;������ߓ�蕍L���'�s�)�s$VY�.��i� �h���?��fa��(r����vGB�]�Vo(���u,Ǣ��g����2S�%>H%�6/�Y�ClrʿN�ʴ��R���w�Z������4��RR�1܀�`��+5Q��ja:��Ly�
�l�Y�rf�b�N�۩�f��ϱ�K7t����mZ�<Ai�L�ЗA���<��/��`L�b�<�cͱ��7!�s�xe�ݗ;�ۂ[�D<�xZP�L^u	����^Ǟy����<�r�s�̠�&�BΣ�K����m�/O�F�ӟ�Z�a!�Ћ�OP�]H�������;;��h��z)��.?�m�h��N�\^�1έGs��T���ڭ�2�<�#�$�T��l�Ä�]Om�n�B��ҩ7�f��Nz�ڎk�3����^�]�q�����Ĉ ��XǾ-/y�/�������ƼcٕlY]���(�Ʒ�ƹ�^�S�-���e�Ejl{��{h��z�e1e"l����}�\ѥkV�B������0\��]�IX�{p[bW��ۺ��H�׳7G�V,(˱�9Ң�����]��M���@��[R;P\z`�f���B�mCñ��xb��&sB��y�9��>�gO^�~ �2+@�2��(1*4���D�ШP+@�B�{������~���������pL��&O�XB�*���ܢ{����/��� ���k�b ^��w5�=+�m�{\+�o?�~a؞��Px��V+�A�*�𵚖(Y��~�Ɔ~�����Yo[���v��(i�`ߪwxT��G�S�:F{�mO,W�ͽ��-������6�>,�)_��:�k�	����<�:a��i�6��aW�1-��o��z��v�4�lCyU6��	�(Z��ht+��a��g��P�m3)YE����\��>���}�w��S�d�ָ<��^^/iNV�=�O��'����%h��z7���T�rI�.Y[}x�F�.J���]���<-l�Q�%�tBe�L���Y��]a�c~������7����~�1����-8+ţ�|}������CϾ~�.�YU)���"L� �l�m?Lej.tM,kK'��ʛ�Ƣ���!�-��T�kG�:n�d݅�=��H�S�Kxrj�͜:�re��:
"��Y��ԡc���>e@1]@��������:�m��l��׹4z:`����B������8��a�>�'y0�pr6 �ݳF#(ۛo.��}��ê!ԖgG����4��*�P�G�=�ռ�ǾZ�k��z����V���]1p�����
bYէ��K��)��}!YYI#�4���G{���) �rc%II�>�������� �R`��
$D� $�JDP���uUn}E,n5�R���%"�F�����Wm(�jG*8t�[2�a���pj^9��|�\�t[���,#���niSV���8�6�S��%R�rG7-�Rނӈ\�mx�fސ����0ږy�F�{0*�m��joG�}\`:sf��i��O'���-B�
�W�5Z�Ų]�k[�g�_�7��c�> ѿ6(����h<�
���@��a8�Tn��e�����lE%���4�6NZ��f9����r��pv�N��^c���2/�jz펧���,`Xݎk,ۭ�b������u]=mc]�&�4��^�;
[G:�'>_��r!�y�v�Ǧ�}�E�ză�����f�dz�h���h�y��u�%GLi�S���6��gL<����2r�s+1�ƛ�>֌̪���۴X*t6ׂ2�1���"��÷*�+�Z���U��K
g{#�A-w8��pSׄ�{n���a��ª�|a�Ą��'��\�e��v^�#/ql\��Ι���F�`�;IE$fWyw8�L�!����e_ �دW7������[T�	ޮ�͓O�����#o��mR�qc盕�M�\�tf�V1�\޿�\��!h}�d��q��$�]�o��^�X�]����\EYR���d���/F�;����َf���;�W�lY<��^��+y4�:S�bd��놀� '�RdP�@")H�}��������ox<�FQJ3��6�;i��������3�Hߐ���x8�;���~��o.Xgb��U�˔����s�ȦĢ�銸�~�l=:��b��(f�Ƞ��ΟX=���i5�cr*����}���3�訴���B��V0֢nr_���] ��EK�=�Ęd����T���9z�5m�:�cܪ�E�u�| �R�������y�,[C�U�0��/�4F8&uqj73�.��.�۵�jqȗ����4����P�MB��^�܌`�ؑ�;�̬�^놤=�&��cTU'`��网t�.z���fs���B��0��J~=��Ϙ#w��BM34��s�D�c�eN��$��6ua�٩�b�V!F'ʌ�����/�5�:}�B��CmN�^-���/��?��`+Gb��eݱ,g)�C�ҟ�O`��JLQ׍���J�W]��-�.�V��&E��C�x�E���P+V�i"hĉ�m6�u-{����i�����Փ�({4������/N��2Xm�.)͉r�lT'��$��(3^��M}�&Oa���;~�~��Ț]u�	���qA�H�ʺ+9� �S��/����Υ�a�+����k7��Ӊi��S-C�E"�L)�?*YفP3��P9ȫ��>$^�;�� ���:-� l�mc�'��cz�q�c����`45a�������&PY�F!$E�xx{����a���0��c��b��A_=�n�����Ԟ,	�xb���VUBlsΞ���J�C&�ی���r�+���wBmڌ^�%��Dű/x���ȧi�<Ył�Y��"р3HIe�9��ɉV���g�y�f{ی�D�5��QN���\�'��E����2���z���*m�ϳ\m�A�ыK�և+�����P�h����!��M�S�VJk���)��JV��MS�U�������0Z˥�\�im
�f�Kn+����˩��R5��JW��;[�X�VN�Z=�HiV܄����0Ysߖ�'��]�3�M늯b^ۖ��C�{M4[#Sܢs�Y7��Su���C��重�k�ߥRm�ʼ���*�@W{Cy\佚I��ob�n(���;��4w���&:v��b��f��'�=�钝b�b\�d*7c��ōj�UqO.���2?Zr�&����ܪ/��X_���S'&MJm/��J�R+���������.��w�2���w=���I������ǚ=��wg���� }�|��Y�>��9H┫�?�sMV�H�w3���[��[������p�0.�g�bp�^�3����oS8�{�g���W3F�A&��-m�Hz�7
�eJ�u��nIY�z�=[�La��f��[j7���ԚD��K��'m7�s��1�^��?���W��)2 Ģ�@� �P!A���s���׿__gǜ���>	)L�y��	�l��_]�<�1�F�P��~j�������ٲq�tc�̜%����U�qٽ<��Gs�����<*-_��4?�q�缏�v�#��[����-����]�!QL��=E�^$걸��ȫQ��@�SkW��4��n,��d��9�e5,��h���A�o�K
�Y��ncCzՖ�1z�L��3c
�����ts'}a��.��I5T�ޮ��<	��Ѥ��@��L򨏖�,+=�駒�[����m����=F����[��}ڸ:A��v�J�9µ�D{F(@J�.(Md���}q9��v��bY���'4�mS��gp�����d�tW�tkW�7Ï�#Y�1JT�����.~T/ �ρ�������1O\"���O���8���H��U���wL1����g4�+yIT�mUN7S�u=��n�B�њm��T���Bh�R*]
ǿjƑU�*!�����=6v���.��;oZ����zC�j��5���8��:!�dsg[�>*͋���0��i� �[ml�B�](ڸ{�u!cB�EqI����8]s�1��5��_!G'*�@��ǉm�U��Dc��'Bf]��7��[.�Z�p��K��>�I @�쮡cy\yb
Pz�F���\����Vlӱ[�'�T�a�%�0k�[�L����@�n�gG\�Z�J�ɕ�]��k���]�����\�Ĥ]`__lޛDdݬ�]�S	��J�RWH�o��W"(����q�L��ﻺ�]�hU�+�$��8�i͔L�%<�xv���"���{f�|���0i؏qn�tE�e�2m�WE4�n�n��?��ׁ��Zf�@͡{��[#�u�ل�X��6�;H��f��|;E��ύ�40!������|7e�5��A�d�ӆy�I���y��i}ɋ�|��f�v��f�3�^��۠�� ՘�����f�y� 86�zoP<Ҽ.�1 �3\��$�X��Xf���l���5��V�5V,Tfҕ9����-����&�,"N�15�9��;�J��­i#Rq3+^\�J��W��j՜�KVK��C���i���;�^�@M�V�Cw�<�:/��3��&U?�[]�\h�+�Ӓ=���յ���ms�(�(l�o��Q�,�ܝ��`d��x��Lۈ���z+�I��Ǖ��1̩��+Eӧ4o6^u����%D�S�Lk��b�ۛ�ݒ(�=+h�kp�ˡ>�VZO7�<U�7���&����W�.���u�s��Ɏ��t]1�j���L����	뼠́T����-�=v��H��-u�[z�a���N=u�Jz��^xZ1�:5��7QM�E�v401챹��3�2nt2��n�|�t :��2��G͒(SG4��p�ۈ'�T8{Fe��7��A�����DQ���!ꗂ���A��
��[�iu��t�/����!�p`�\B����)|p1�C|nZ��#2���и���Y�#@����؟]�[Z��q������|��S�������3���K�-����.��)���V�7MN뽩�\�HS�xVC]�L�K�ka�F㎯maz��Wm,�`(����Vw9��]dzV�C�#�DE��^bŲr댪��݁D��&��9�t�b.��Nfl�3]X荝S�<x ������w����o^�1g:��8����ʒ��}��q�L�C*%rȷ�E�";�O;km��N��;k�ƝǤ>�z���Z7-��U�ClD�$4�ؐ���@�=��C���-t�V��FV��.���h�|:Y�j�κ���ˊV�ӕ��T�({�q��qn���Ҿ��]�Nh��+�I�j�r�v��ΰ��L�}���<�]��,�.���Ȩ��V�I:I�x�f��j�'Nu�r�(Z�[�fu��[rV!<���*l�y2�u��!�L�8��Õ2����67�C	o��AX�C6�g����M�b��f�G�]�w97�0D���4��T�4�[j���*�(���%�3JED�F���=|}�>>�ƨ"i��(���-�EELRMRD�nmMQ1PO�[������j�f�)����*"� ���h�[��ͨ���b8xz<<<O�g��QL�CSTi�MUS�����E38�������.c���""���TgcQ<� �!��( ��V�"�U͉�SLA�PSEIL3U1-D�E5���Ƙ����塢���i�mM�V�IUM�TSU@S�
M��F��QCZtj6��i�c!��KAEThڬFهc%0�T��UŧIL@ME1Z�1�$QQTUk�,QTUh(M��i�(4h���

f4hִj�����9�*"��ED���ĺ)�4�,L�R��÷�����2i��[kSUs@��Xz���#I��xU���]��c�D{ؕM��ޕ9b��s0L��ļ���J�vHo���~zsp9s���7?!A�d
�(�"U�	 ��A��������wׯ�EO�=nK�]��5��Z.\�.���<����UL��]6۴������Nl��ved_B<7�y�j�['�\G(F>>����
�z7��WɌt�kȤ�eoE�6!ֵj�V�G$����X�/~�&����/���ǋ�����0�2ݠ�ɜ�{��P�םp��'��nOaDR}k=�^*V�5�*�y��
�?�@���P�:�/�Z����gz��VA�����:��T�zQϧ��z����wv�����Y���[���NYӤ����,�oE��z�s�-M�R�j l()��dPZF!r�m�Z�\>/@��2���Ows��A�':٪<��i�Nl�^<���Y^�}1�j��D��V����pE4�����c;�(�#�"���	c��&4?|��,����ks����}F}�ςb����wMQ��P��Ύ~�uǁ:���u�2��p��!A���69�ڨu�zm�5*Y�MZ˷C[�d<f���4a���|�D�߇H��V"9<�����d_߳���)o�ڗ.~K�Er����w�o�̔�r�B��]4�ܺ�/���`��|Ị+�/}�S�lx���Y,��{�Z�HN���r{թ��9�a��5�bG�te���t�_�GWv�CM��iuv�;+,�3�����7w������s�]�~Af	�"�
"ZYP+��0o{�3�xq�]Ȯ��	L��7���ip�7Yx���$6�CD�O��Z`I������3���u2m����+�ľ5�[	�e��PջƝ��*A��"MvJp����	_K�b.e�y�n{~�߃�୍����T��*��l	��+��|e��$�3s��O����aH��u��L�T�?L�v�\隋�_/5��]�.��(�H �_�\^O��}2jYɵY�e��+�%�ck\T:��r�n|���ynV���9"�1�&2��
K#�����if�j�@?ń�F8�i��1o�����7��n ��<ғ}-l��L�L�Y�	I�%K�ײ �˰]�(�qj!�����f�)�!Q��8�d��)�9�R+Ͷ���K�}��]���h׫o�׬NxP�^6j����miM/�,݊a����b�EE�DQ}ܾJ�x�GPMr-��ڹ۸1tS#R�h��׀�ٴ'����.C&�xbۙ�.ۜ�Z�M��Z�<lŁ�A#��ݬL?u����z��Iw�� ��c��:n���͘p�����&\�BiO��'<�̈{<�k��~z����@z�of��SjW,ꄘ\��&/.C��f������-�A�E	�W�υ��g��A鎠��+�M�19A�ې�on_
-���\�ݧ}Bu($9s���ً7��|K|�29��#�J��)�W;���X��}{ٰ3k��y����������,JP	- ��H�*�),(R�y������������_{�}��w���a���A���e�	���%����Q�ES08U��T���� �(�Ee.k�'#�Zbu��|g�urVN���}��g�����+w��SQ�<��1R�-u:�nx�.�Oܨ�W�T�~�^���C�$V߳.������w�z1���sjB�z[J}��ks{W���m���k�lw�B��F'J�`mCD��cg�C�Q�Ы�"��^��Pʤp����zJ��!X�+^����O(+�v�l>�]W���?4��	�j �5����}�ӗ<:����3o��g�,'L���Z5E�[��/��,i�ۼޮ�;#���ý-��9�;���~b��~�B���<jj^:��	W�/Λ��؇��e�j�{ZR��@%6��8�é�u�ZG���4=��4����܋��6(�]�J/������Y���.�CL!۞�E'��+(V�5�)��C��˳�i��^p3�֙e�ixۜ�ɘ�[���9�l��4hb�ؠu4r������y��+nXP݌e46q��V���s�o��η�-9�t0�G7�qG&%�,*�n̲{{aĿA�L����;{6�;��Kl���ݸ`��Hz+ 6�Y�k���;v��gnKE<�}6��Ս3G��Q}oS\����_�ik��֒�T'ݿ�� �|h�|{�w~={>O�@?��J�H4� P�Ѓ^��7�������V��Z�.K8�[�h�q�Tl�sX~�6n���J���LG�jJ����ą�<����8���pY?@�0���'��4f6j�ϯ�%:��Ly�S�	���;�|V�s�Y<7ߣ�nlj��'܇��,�����A�I�x���<������<���ε��M�J�!G4;����o<	������g��Oxd͒:�Nl�,;Y�r��˅��ʹ�����:׈*�2U��h��@Q<J��
6�� �b�}g�d)|��}�Ջ�azP�F��SL�l�uj;��PXN!R��>D�cC+�%��T��<��^��Ϊ��{��*)�GIo_�y`��L�Oǁw����k|�..�E�fg��D��:~���xk�8��/Z/����r�'Vny���8�x�6=��}y �In|z FѪ���Z��7�i�'b���]����7�>Y�� �/Wរg63ְ灅��0n{m��c-b�#��Т}ު�_�\)up�^���>a��ϐ��VO��@GP�Ɗ /��Op��]�����k���[UMP\mvnt�tv��+��*%N�ô�ӣ̩ld�2t�$�4l��yQ��Z9Bx71ퟵ� �'�eN�B���qs��2�����!)��P��^�t�N�:n m�(�P��: ����	0���(Ĩ�ЩB�$�������������������n'ȗx�D�@�#QL�3l��t�몈��l���
��Qg"�4��N���[V{g�z!;b���ƿ2�|�8�xr'hr�wML0��v2�9?�����-?Kn�w^zp�;c���p��T�@{�������BSEZ���6ǉYb��$UYQ#���˨;�gI�x�5y[��
�vų���@Kv'Ź�Sp�R����2�[Z��*�şz	�	�e����vm��hŉQ&eJB[�3ƥx-1��E�����M�y%^s����DoctB�����.1��}N�[yzK��؍Tc�ܨb�,Y�7:���0�!���]�|�c!^�0K�Km�4�@����3m���j����*]��xBn���UP7�뚧e�6e��A��p�uJ�|Q������	J��%@0�!�ux�DB}m���M).;{{�8�_����!4�>�޹oa9"	S�הA`YP;��2_��:P�:oޓ��|)=g~�pN��
�(�	�_�e�w���T��]AO��#�b�*���E�cq���e[q��NL7hu�d����C�w��c�i��Ov�c$�K����xIjk�SM4^�j�T�N�p��)��"���U^�ȝ �g'*���"����66��Ȍ�k�	F�l�b4+�3����j���ͮh���������@D�P�H�׸��b��3�<
�Hq��%�5K�kH�ޫk���<嶩O��`'9�y��q_udt�)d
l�m�9�<3��cK��C��*Y�1W�쮠�wF'��M�n�c&�V��b�^vH����u�d�|��&�MC;������C�lPZY��
����lt��>,��1�&�]�n��A�� �j|�@#�4W��_���DA���I��~>PP�G�|k.b��Z�=�>�˫�v��P���f%{;7�r�v��	�D�ASiú�r�Nɍ�r�����a��tM�i�3�ol� ����Y�����a�n�h�� ��>��>�[��9��ʙ0P���r���vK�lnv�[�&J�*a�[y3�u]���Jk�|e��P���sM�)��F�	csE��5�v�a�ӰC|E���ӟC����
��1����?r�Zם2kƍ��'Z��{����sR�����ֻ�U���n�H����m����i�l�A�6���5F��0{_�x��[n�E+�}�����[�4�@�z6�#�~����KQ������K��i-DUU��->zh<��o�����)�@׈8oV�f�ׄ`O�������R�[����Ϙ�&D;�C�hf} �������͍Hp}�af����_ב�"m���k[�[Z����K���=e�YH5;�;�g�D�0��0�"D R(%(,"|y߿��~�}��Hn���L�8��*���ӓ��^�YX�Z�71�^;ʦx��R��uj�m�����͈�>Q���4Ψo;N�TZØ��(�/��P<��m��E����?m^F�}"uy������76S�&���.���U-Dܢ�<�=܌�1ͯ�|�ZV*�rY���Ȋt-	�)&a_�m��M����͑s1V(��d��T&���\_:��֤�'+�Q�۸�f�]��̻_���g·Մߩ�$m+�|"<�٩�b�V!F'�ͬ�Aw���2p�\��i�v�XZ�)�ʯ�?+��8��Z¿@8#������<;LZ�.;ERa\=a��Ce�==ݑ)׫i�Ԯq�4-��H�뵧>��P>/�C� gȑ�y�x�5*�'[��l��5��8�5X<�i�p3&�J3_���-��Tbt�^	��n���̈ˋlbˁ��"�f��p�ϖͷ��^��V��5��
�M�l+
\<�r���a��Q,҃���'����yX��vf8���)��~'U��,�2�yu3�M��ݘ���)_�bφ��IႴ����듦.U8�_��Wx���b����v�mK�$�JF Ѵ��]��Ψ#���):���'nVu�l�q�7��X���w�%nv���AgEI��^=�8����x��V-���1��9�v��s3BlW�*G|��_�UW�*�	�I�"��R��h��W�=�|�{�ϣ������O�Q��~ޖ�P����55@�Й>�v^�Ԋ��g���b>�&����߻J�Xáj42���l�Sn�#��<4��T�/L��8�f���!=o[��f�S
�ٵb��h�qi���a,0^�Rq�a�C�yOC4��]�m���Y1��˃�^y�۷�p\��`nkCC����r�L���F�ݘ�����2籉���ic;*�qv5mC	��mZ� �7&���^�Ιy6�^;�8�.�q"ܳG�N1j���k~�I�<T�c�^=,̡����%3�}sV�e�:��M �p�B����	t{ �,�f�f�4��:��*�ΝB7�a�_��Ÿ�!�ﺷ�om���*g��p�"��.=�h9�^ǔ��1A댦b|C#���˲w_E�u���E�%��9)X�)v�}3U�������W�S��K'�>߂�ݝ���s��� ��R�ăv�XX����ؾ�Y�p�5��S	%�|��*g_��Z��H2Ӈ�ٖ��fm�*��Q�x��R��_�˧�Q����
�U}�������|���WW���J�>����Yu���M�˻�ѣqY��55z�C�9��竜��<�{k;9�s�5���Шn&n�
�0�@چv���Txa�wN�;�3&�D����M�e3�̙��m�WV�}ݗ��)��S�������s�߮k��D��;��"dI�"hRI�
�Z�)i.����!�,3yko��az1`'R�݃��7�ĝV7Rwӳ~�S��fe���c<���A���Z�����U��i�^�???0��[��@��2�@��Ol���_xʐ)g��;EnP[޼�F�cCq��[!Ѹ�p�����h�-�Sʈ�`�{+��$6�����dD7e>_����H��^�0�\�ь�Z�ޱZ�^c��x��S�F��A�^��9zL����8߉��K�c���^�$`��V0���:y��NbY��04�iP)�̬�7.�'�v5��dn�SCU�8&,�A��BD��۸|����öxl��VD���GUVw	�u���ni�4�����Sk_����@Z��ht+Ƭi��!�i�@�U��o:�o���Y&�~R�#�S�~�lO�I2��2}+f�u��ol�������7S��v��M��6�?�R]�<���zki���t��kd:$��5R�f��g40*�s��7E�co��6O��p�T^L�yO����p�0.z���`[
ϗ��+.��ݔ�5*���G�DZ��0;�;;,Q�����I��̃A]!�X5���FD'q�՛X#�͜#��ոGi�Ȱ�u�h���2A]&�J�$�Ցۊ*O�z����åU��3��Cy1��V��ڹl˃ȋ�C?����>|�JD�"4�R}����(�-[yN�_�1)���R���M6HW'����EC�,�J���:h	������������;�6�K!��(=r�\W�Ү/�1B��=�\�F�5�P����j�}�/���It�v��'z�~���v���eئ�dķ�	*�=�D��u#��S��s���pkT^ܘ��7�5�׿s�:O��\��� m��^]SmRZ���J�n�&��9�l:rڴT�G_<�M^̮[dtNԆ@f͉�}�!��&^s�46oU��=O�t���U;2�i�ci�kk3���l1�5!��y���a�G��5�����&Msϔ��v�P�,u���ܩﰴ�����,e����l�_?nG��׬�q����wT�΄qrF�,m!�+��BB�/Q��'I'+q�͘�꾩Mo+uP��9�a��Fӽq�(�/NdL��i$gm��ӷ��ט�g-��n�����~���h;_r�v��q�~�N���׹��Z�n��T��~�3��}c�<+������[X=)�خ���̈́[y��v�Ѕ��� �x=Y�7�~<n���7/Iz��HZ�Σ�18h���}2uur`l^4R$o� �P������A�����`M��K�s��{w��;m^o7��%w�S�^�R�N?��b�;v����H@�]-^>�WY�n]sm�na�n�&Mc�(��(a���q��/�L�gPz��1ۄ2�ț�8B������|�v�'zVu��& 7(�`�Zt*:�[������݉A�̮Mo.
�	+�n漽���
$���Ǘ�o �)-�3������1T\y��RP���X6�x4�AW�U��b\,b�SrK�ʅ��.�x�h��w66A��ޔ�r����Ց�tp���r������N�7{��Np]���f���<'�V'�C�3��k�\5���(�]s�ur�{�t�ۧ1vB4BXƊ"D6����n�s���?�n�̑ ��V�,��|��YI�ذٗ&��MܢՓ��@*��v[��]�ӽ�-�ʱ���PЭY�cD��%��z�YX�M=uД$�N�6f\���&�Uݶ�Y;)�����đJ���pP�z�=vjm⏉D�WW
���@`쥉���e��j#Ҋ5�2�ݘŬC�<���Wc
u�k���͖-b��S�ut!��5��-tz;	t5�DZm��[��v�t>S���5�1;O&D#z��mY�bv�V�����%d�0���V�%c�iv�;qq�����I�[.�l�C8�s�.U��[�G�֩w\(�1���~n����h��9�j�	�|��V[a{ݻ�0�A'�o���䓚@w��^R��h:�9�peY�pz�2P[R�EKT�I"��oZ۶��-���ThXX�z�IwdЛֈ�yj�y�L�\;��M,�U6	��v�f�U$�ϻ��ɵ�E�OgZ��m��|�N�a���g;�ZS�+ δ]oD����Wk\��7ёu��+.�c�j��cn���Յ�Sa~壹J���W��W5�s�����ɘn��`�,R�W��H���ظ�����q�x%���x�Y�M8KۻpG�ߚ�rɲ�Vf��F�Sv��jV�Q���+Xg^�-8�R�3(��m T����$�UǬ1v`1 �f^s�Jr���c;b��F�|��������Xlk:t�e�V�-M�u�YOA"��4iKM"�&D�1�M�*���/�����-�WS��i�k�F˖��2V쭙�r�4���������w�,�/1k�]�iP�N��qU^�u�κ`�rum��s.�䫝f�0��-��g]F7zѺA�S�Y��3-,���mIxh��`I����y3T�V�ۿ᧥�XG�'�=�!��k��47�K��U��bwc���:�ϑ�qYRS����7�KEm��������:���s��8/�&�J�Z��*/S���
���.FmE5�-$���o$�К"�����]%4�70�ZJ
t8���s�����y��y�)-gh�nG&(��yR�u�1m�������䖌RD�b���!��t4�EAM�.K�(墝b
��v1�������T/�Q\�1[�����M4�QED�6*b�����sh(�j�&���Z��Q4I14m���ss�UD��r9p���Slj�
(&�h�I�Y��ĥ&�h��"[Z��r����s�98�6s1N�%4%Dm�h�����
9����
(��"�'d�R[<�጖Ψ)����QE3H�4U:t44�UL�t�h40Nh*�ր> � P#�2ˀ��ܨm���U��϶��.G�1�#�Hu�AѠ�

8�s�*�*i���U_���e	�"@��R��R���©�6�|�x�/�)�E���MG���{��¼o0�O�2y�N��E#�+�CJ����~�r�'�3��H��;m�T��SY�/��b��|���gX�^���aL����x��l�k��Z�Z��7bٖ�	e{x�YL+��Vn���}I��<P�+~��:vz؊�ʵ;����]Y>b��-z���u�)���)�%Vk�zlه��쭅��&LI练o���������/h&�����N���d���/eE��U�+ki79/���5�Q�mOwR���X�Db�FcO�2snY��Ψgi��)VZ����_���H��dw8�j6�_u�n�!��Z���L'�L��- ό���#����P�����I�]�e�l�l���:����3߽��bt	#�HG�P�J�L�?��=�E7a�.�x���1�S�j��wW5+�y�H�e�c�hE;�tc���������͚�dЗj�
1c��z��u&��U��d�sE<���I��g�׭l��&k����?�pv���Iи�����|����L���
�[jl~q�sff�.hP���L���͝�&�8����ڹ��o��}���c�fa�(E+�Ͷ����~c�L�M+������ȳ�:�D��jS�,os��x�΄n�:|�3D}DY�z��,%�+��˩V?� �? ?�(B H�ZZJQ�����߿������"&>Ǥ�����p$hcU���C�އ�,�|]x� g�?K�&��~��z�{'�u�G�[р�e-�M����������z�<�h�փ����3���ىȝ�z�#��(]lX`��|$:b�C619���i���.�	�l�a6����}�5�j�it��E���X�U(�'J���U�ߞ�vv��W�~��3%3Cu��Ѱ]�S����oiWkE�,���f�n��1.�͊:�p�\Ly���:�B��r'�%sV̈����D���B.��Cd:��y�{\9��yI?��Y1�J��7��w�DA�����O��n�&��wWn���t�	c���e@Z�O�\���SV,����˨4cc���k��v�(��ܡ���{��t�5��ӵ����Ǝb�ִ-�Oַh^�U�����2nCVR�;��Gy���������	�|LR�b�2v�鯦�)>�*|��0ض�_j�p˹�?5I&�dg��|����R�w��Q|��A�����f�<��钝^�e�F^�U�Q2,oc����)@��/�]t�;\�^���=�o����=	-XY&�#�#��ݖ�u�ٶv_(k��]AU�nNpLq��f2;XD��C�w��[���O\K�I��&���R	�%]����RU�$P�nsC�o�I��ٻ�������Ϯ7]Ɯs��~ f�&X����� �f]��)�aCm>|�^��7c�G\��ƹ$��^>�R�?��V5OO����ˌf~Iv~|߅�WDy]~�UJm/�1R�~�mJ8�Q������a7��^=�1��)swQy>aU���oj츣z��Sӯf��U�hˊ-W0(�nC�X!����mw���Ү��,e�0��FWU�w��ڹl�ϔ�G
�N;z5='�q|c�,N j3Oă�]��w�ī����l�bn��G�L��k߄�.su���u�N��ۉ�z�ĳ=Ѫ�֞�X�q�3��:�U��^.� ��^�j��,@}k�d�:�s�/\Q0Z�r�yk��j3p�m��=��y��C��tm�Љ�>F|�z�����:��g�o�����rH��M��{N����v��r���/J�9
%��8��r�rb�m�z�ָ�Q��M�N�k��ܷ�v��oD]���/͞N��܆�� ���21L�wF�z�p�8�>���[;�E��K��0Fz���Bj72/*1�nmSc_��r��B�@�X�y]C	�eL4����>$f�coF�'y�w�6<
���+�;��N㻭��B�͕@Y.�G@����k�!(�AS��HN	�ؤ��,�C�˗Yó8P��Nk��Ř�#�l{��ޑ���]���}e��{�� ��Q�ݫ��d�&!�~������^}���_����8-w�
�;�=��ۿ�'��M����WB��[@�(�`�W�e]�k����8,�?Q0@7ɉ�5�^P
i>- we+���8�%�I��a-��f ؑ7���n|�M�C�e��dS�˲�j�c���I�-�Y�L{�hh�A�GD����z;j�^c�ɵ�փ��d\�F����IQ}0*�[BTZ�]7�D0�ج�0̂����_73�u3F�=��s]0�
�MݞJ���us�b�!�3#Y�[G�hs�rV������b��&�ѷ�>F��qc�<��z��\`sJ�>(�O�k��R���	��K��xM���J����+K��kp���ak��@Lƿ5	0��dK)�5��&(F�U�A.�R;_S��'!3�� ��v.�;B+�0���c�A���	�hT�d�sʋ[Je���
(݊.$?S�����nѬ���������	�DƂ�t�??3OB^y�CCk_�w���;��~2`���4TUiɞB���"�PS�i�UXտ��~��x�cK��25�9g����͝ez8*�sq��D�Q����� ��LX�~���nu��P/7���	BK��>�>�M���;�� �^������Q�)������Y�lж��ulW��\#rK{��mZOj�tq]K]ztM��`�w*�1�w�G�_?>���瞻��`��"(_3{�q7�;�&�C��6��:�v3�s`��~���.5�GWѲu�?����ᧃ��;�7�]�D�T�^C|�~��\����za�q48P٪-Nb�8@5����L���1)�U��e�=��׆[�ig�6a��y���d�;l8��;P!��x���c9M���ٽ�M������[�Q9as��c ݦ2'���W�l����w{�Y��!�0�-�{[�.��=٣���N���ｵ�>I-�	���Q���*��uи�aؔO���'�׬�ϕ�&�J�ُ�o7o�����+����3�m���Pʩ8X7�T���*��q5iRc���k��y�66��C����ɶ�YT���V�ߵNC�M�e�.��!��ʈ�wk�.W]V8�ꥺ�+2�	c�����=o~�N��<��E6P<ҙy镚��>O�؞E)iV���7m�=,w�R�]���A��k}Ri���Z�='<}�����5�s��͉�b7�We�Μ�|^�,�$B֑��d�o��7:���y*-{B�����T	D����Y^o
��K�p���z�r��R;����vٛi�4��������މpj{3�Ƿw�:W3�:�T���\��Lq<��e.�2��m��$�jQ�ծ���\Z�����v��W��;w{�<���^��u>N��uW�T݂�~y �o0`�`����q��75Pc�B����{��!�?r���.>3��s�s����ܢ�m0� �6��c���۹
&����L
�,��q�6b���f�H�y�E6+Jz��`��7|����gh]n�a��.���օ6�����*�jIvh���\�C��P��v�y��X�����O_d��|��){t�@0�����kg�	��5BcY�^;s���Y��&�׸�Ό�V���^��)O'ͮ6&���l$hcP��T���1�ܱ�p��R��/4ZLF��Z���w�hT:�����D]>�u�����Z)8N�~zW=���-$��6R�+���TK6�W�Ej�Y�@_�ް.���W>��5�Y�өev�|h�4���2W��0���}޹�ꢹg��M?W킒y�OL!5g�����1�S�~���u(E�9OԠ��G���Afׯ$ь����3�Fm�WG�QB^���>��+f��U�Y۸�՜�X����ܼ���#��i���PC(z(A�# �V��w�ޖ�0v\m}V��/!+u�u�zE�[X���i�T��ph]8�?���kJ�)\[\ȩ�xd��vv�y�o�)4�e�W��P�l9�W�a�CQ�_-���q�ז������c �J���w/0>/�e���DJ*9m�������C��]pUھ����#e�������`�X�8�����́?
�op�÷�c޺�е�l�(V��VF��dmO�Mj�̰��?2��,�v��D,mL�_�j�	<�ƷP��M�}Йs�ؤ�kv��Sx�4�Ly���~�O̍ԏg��?����~�8�NY�Ʒ6F�W5�锟q)�&�����Kgf�[k�O��A@�����q�=�¡��e�2A`3G�T�v��I���,�1�Sgy���e��
�l����mϥ��.9j�o�h�� ~��[��DƸ��X([��Z뾾�NC��^��b���L��u�X���C��E*9@:n8���tSM�VM�隼Zj�jP��u{_���a�.R�`et��9�P�ύE˳�f�iW ��p��+w�o��-HLF9j����=���6.�T���ިO^��0�,8b/�v�/6�e�{a*�����S��@�g�̝s��jsu�}�]d��y��F)踲�����Yʰd��Otdt�����r ����}�E����G�q�|���)�z�	ֲ�ԖK��pQQwR�hs]:YR�̣ �n`Z�%λ(v��Z[����2Oki��.��[{�d�u�g�1NSI;�*���		�;�D�5=:��W�ֻ���"�a�0�nƝ�غ��Q����N�YB�#˚��Y���k��=�8t�ɓ�a��O3�����h4~���(��׾�ɳ>U��%�xș|x�*�1����I�k/uL��tN���zc�yl�K�1V�ٽlk\4�S������-uGx��W�y�Ү�vN#3%�F���`Ǡ��"��*m�H�y+�2V��fsq��G[j;��a�M;9�ES�x�5�s+��Ň����f�x�>*eC��9^�X��L0��]EA1����}#���x����ϙ��=����oB\�����SkX�"SExZ��h��X����`�t��m�ܵ0w@�I(�2}P�JL���e�K��o;�Ċb�Цڷ��~�t0Ԇ�2ё&`ŕ����0k����)���+2�߱mD<�T��UI�Pd�-�f=�4�a�pe�6"��Fb㲩k�ۈ��8�Y��چ^���//�~�a*/~��W�e�Ʀ����[�T��Ҳ��Ԇ�:�L�龧��S�W��mY�L�{^�M�u��۞�z��7�9o1�le: ��@M�Pz�(��4���Kά<p���Ve��&*o&�Z�g��7���w��wh����L���^�޿^}  �VϮo�s'v���sj�+{D�M���k�
n�����;,�%��᜺Fw��\��)����t�s���V��_�+��R�u+��d��˯���(D�o{������y	w�3_.��a�]���7�%h2����Ȗ=�c���^DH��{ �m.q��c;V�t͎���3$��>�$�cD�Wڇ�\BK�-���E��J����uxP���,R������fn���>���`Ev�A��>}���QC���fᡢ�(��9��V�_B�|@t&{�U�j�z�|�Kd���dDh�C�l"�.��\Ķ�����t/sb{�!e:;J�k��:��&}��B�HأQ^�M�;��v�4��A`%*����d����~�]&����c�:���W�����˾������oş)@���|�����y��c�;��;L��N���fM��B!��36Iѝa�;�S�Yx�\D��*�\9Ry��¦vbaT�v�!���C�2�=��u��C�yI��c'�9�#�F�v��R�l�j��}�畺���;1.DA�w�)@Q�튽�3^��)a1q��_�V.&�u{��]�Ў�VgeL�����p��f�3Q-kڲ��'�����Q�T}G�& S2��5N�^1��+Ej#�o��%_�`�ՠ��1�}��n�����q�MQԔ?ym���IBU�缄q� {��g��`2�(ݜ���kE�m�uٗ%p����G6d�/�MtGEuNާ�gI��V0;��,���ݵͮ��'�n��[ٔ��[�OY$��킖�[��U�Uwo;f��.G!�$둬�2bD�m�V�nW�X�!�[���C���4��7�qX��v��e��wjC`k@vGW��V<���Ӭ|��u�!���*�UC����I�K�M�尡���̼Co�h	�~�T��K�'k'��������q��ik�)��o�Ed����3k�u�)��\�"���o??9�.����P�O�A�O�q�ѻ�r��9)-N`.1`�����{�g
=:{�n#����h�u8�ƈ�����R�75��k��(����ೢ�nUV/}���sz�_u�L-�������\�i.���wpl�6��l�|u��͑s1%���r[�,���qS.�Ti�\�'⌖[�}?1~���#�h5�?FDϾ_{=3ԅ�i�v욳�r�)�aF.���R(�)�/-�hOV�|�D�sw�pf��I4�pF�M��V���[eo��r�.{�Ǣ�L8�9�1i�XK�cU�B�u���%�Ʃ�ڪł���k��p� �!"c*�H����~T���i�ڬw=�ݡ����C�����Y��:���oedJ�n������U���9�t���I�ZWu��4�V��Պ�	@�oI�(taS�mW��Gܻ"l�#	�*��E[���������;�Ƅ�iW)�v�1��
w�ql�ŉ�>��V��<}u�[���ud(�ɭY�0��j��,�WL���C�����Ԉ}4gd�s���*L{/o���g��V�"���9p�]'��0��k�D�J�	�9N�E8�ݽ^��I�>��������Y�7Y����,n6.8c9n�߸���jiv���P��b�R'R�9�*«D%R�Co�y�y�޽�Ԟ�u��s+d���V�o4%��A����m�.�M�ဋ��vNhu�Y]��"J
m^m+�=��ə���h�'\�r�ɔ�ON�H-齁�df��kry^4Z��F[����Y��\�n��ðc1��Ҷ$��BEjg6#JuBG=>�}ܚ���1�RG��u�[�P���srs䙬��0αϑ�h�m+�e�+5˸D�6��b����.�K��K�+��j��BJ�%���!����p�A��
>uƧ�9ԠQ��el�urݮ+� 2�K�����it�j��>
y����'1;�/�-Ι�Sj�Twxk�C�X�KV��=0�_>}�U�pZ-u1��aS����W��2.˛WbV��Ԡc۲��d{�Z4�^0�^n`"ُ�ق�4r�9�[�(��a\F�l�ܔ�Z3E롗۷M��b��9�KPXУ���KPb����҅��q�P!����l��)��.���5�è�s�����"�X�FD��@i��8���dÉP@�������Q�����zU̱G�1[��oh�LW|���	T�7V��M����v�qc�`�r��{.l{��[��r�8,��Ņ������w7�4�ںY�Ҍ&�t��Oj��X�0l����Q�
[�ǀ��u�S/l+O�b��I�f&�V��Wt�OSkkNt��o"�1��Ī�t����m`IPy��K�y��y��
�Ow�w�g�[Vr�+C�µ]�mt�9f䮲�� ����U�c�u��
��R�Ȋ�������wJ�/VVYK�y��d�7[��D�^�S%J3�B��F�S���ے1��J��e���ƞڢ��ʛ��QaP@������.sʾmQp���L����d�0ޓl�ߕ��,���<�V����<롎�3�'�!ˌ"��J�|C�r�L�7z�v���:оJ^�Z��_!��Bt�2����ȃ��x-��y�q��&��p̤�Υ:1��o7M����]�q��^.7�!��R�s���R�֩9c��[v�t�Q8�|����7}��dR�*�"��<�7��]j�k�A�����t�lDjպi�9[35"�V���:U��K�M���R��j�
nذX$G��5��;pو�1�X(bt�!�1hW���6SIkLUIQ1L��6ƈ�h�5"Ơ���bs��?/���b�j�gmTU�*��J�˜֐խ�h���k�m͜Z+�C4AD������<��E!3pQm��&���Q:��M6Ƃ**-�E�N�5>X�qEMcY�EM�UUEN��U;mV*��DBV٩�+Z��
���4d�tj��F��ԔUU���6��Z�1cc���:�V5��km�MEQUk0��A5BN��캊�։ �(��g؉
�j"*�m:hgY�d��jb������d�DZōc:1��V2b �5@���刈���6�Ah4V�E5TUkM[��9����k9�����PMUT�b�T��j���1�L�4ES��/V.N����:��(�H������clֱQ���  ��h��x٪�_���˨;9���ͺp�射�W�Wi�]΢�>�)�J�Zr�ְ��L�g8�;������K�VlU��U��_K�z3.om�?��E����И:����3-�N(��z�J8^=v�a���[����GQd	r�jis���ip�rp�lύ �vW�Q-����,� ��D1m���{��&��U��V���#���ZP���M�Ҥ��tWcB]kƵ�2{N뉀���[:0�%�%��r�bfV�8��ہ�#3���k��J�PȖ�����O�h�+�8|�K���j�{ߴn��r��
w�P-
���1L,0���eVzl�`Y"w��	l:��sz]�x�V��\3.��>C>��^��J�gJ#�y8����71���ܧî)?X[�/n�
vb9�/3��;7T�[j���w�L��G�@�?���/�(M�f�T������gP�ɶ1��vBɅ�w��gA��g�$7V-V^�̡�����!�M�aR���2���ݑ���&fw4���aw:�x��3ɠ孭����vd\��Ӵ{�	����L�r�~�c�w�禝��K������}�5�a1OaEJ�9�ӏX��u�m�pf�jV�ߧp�J��C2�l�pNN��v]�@�]&M�B��俐��&\睲�c�D�#��|�VW��r�����{���g�r����
�_��f�=����"��;�n�6���VQ��fEx��T����>�I��7z�Ҫ-ۚ2�����q	�3획�a��U�l���x�i�Ϧ�/X�B��+�ɗ,ڮ`Q�˗�s
;S>�lv{����/�ږ|�/{�[0��1��0���G�;8ػ�R�moT'�Q�
���c�B����OQSS�%�
D��7��`̃o%�:��S^t���N��I���{]���H�SW��xgC��h}UGo</�_"}`�a|>0(��:o�\���~��q:��c��2�����C禧�������_:�{�3iy�;s2"}�0؊I偸)���e�ѕy�w�����:�t@����F�
'z���.���ZԽrl��L��1�{�ȣ˫{_�0�T\)���>�m
�dg�m��)���rvPq��CJ3l��æ]
3�9;����č_io��~"��Ê�����V�B��1��R��ԉ�Sn��2�>칃jq�&m}Ӿ3��G�th����8ܨ��V��q�O ]շW��kj��MjBmAt�X��/3�7���_������EW�=�#���(� �޸��0c��߯�K�?Ex�T�f��t�7Rש'x��n�=�;b�7X\�də��e��:�1�ķ��v���`߲m�{J)"�3Ƈ9>}����݌�b��4�ި4Ֆܦu��kr��^s���u���15}�����;���Z%u><����v��Ls�������Lz�V���̱7r�ԚK�_�UI�Pd�,ҧ��4��ՠ������,�|�6��M��禋1�2�?.�m��XQy0*�vo�.�~D[䇉�ҽ��w�ߥ��d!����gd<�Թ���h�a�����E^7gA�0��K�ק���V�I&/}z������Ǳ�ߝ\gȸ��q|1����9�����n1���޹ZW�C�wݽr�i~�:����DG>�	0������{l�H�	U��� ��UyC�ض$�r��z�*���J�|��Ñ�Y�4@Wڇ̮"�x$���e�6��%�����-�GPlfn�Vfv^I�n�#������^��Y��\��ʀ޺*���T_����i���c��wr֙��j��,m�ҧ���-}j��RMV�-��k�71�"� �d<��.C��̮��WC�]�=��%��c�}�R9��F'ɏg�d�}�%�ϻ.R�6�"oMU�2۲َr�YY��;^\$tazP��H��)[�.ކ��Ջ���Z���
��Y�;5���/���"X\�g�]��@\� �����"t\ϭ<�.�/�҆�8,&�NýM�_oE�:��yv���.�pi��Yݨq���Gf��C��z��3 ��9�ܲ��=u��S3O*j}���/%�Wch��˕M�����*���2=�</}b��Z]��
���#<�����} �3��<D� en꘷�����z�o�l��{ͳ
�bt��I�8*y1p���յ��1��^Ln	�����y�Ό�#<;�|wz����F���z"3B��{]_�|(�z�Lv����c�*��oBj=�B�m�$���Uǻq�Vfov��W+0.R���d�mz�W4�~Ք�'¹���b��U��N��L58�:_���l.�:�ͣrofU۠i�{��Κ�|�A�+xd��&[8��k��!�qj"E=����;��q��C����+�Ͱ���g-��M��ٍ�Ǝ[h�m��U��ͷfND���]R3w���~Fg�/���+�S����/Ѭ%�I��&��OI���BϹƌ����"G3���x�d�al��������0E���쟤\[4��v�7�����n���\S�79�Zг��5�F��X�Gp�t!���O�3�|/��e|�:�}3��a���y�����^e���Pu�g�����I�l���+���A�]���X8��a�ٟ�r���ղ�9(�}g���ݾͷ�WF/�F�x�+��~��:���ԿOV��^�O?'��,�|w~;2�f���V�W��GH���3LϷr[/%ûo*&H4з�J��.����� S�r��֝iV&�I킲�SF��Қuz�4�_/xC1Y�Y���a�)��`��[|����9F�^c�ZN�]�ͳ��?0ʹ㐕��W�fj6^v��s�cTˡ/6��u�-={���	T�m���	��σ���x���lL�����k�?�I���$�NWJe�:��Trq�{'V�����ƿ&��'h�U�N{�S���(͞���U�N`V��A��	Mi��0��Hu�kv}����4��,�N�/R���n��B�����p�B<��r�o����W� ^?z�Bp�;v<W���r�w��ʙ�Ķ�Bm�oC�`4>�O��ٰ��r�W�bj���3�$��D���U6��8;m�{�����׽�N�����]y�p�ǥ�U��b�k�-�
���V��M�2��b��1l����R��-��p��>�CP����*m���l�Sn�#��&.2R޺�x6�y]��v	k����4G�7 �$]Dml�Q��3*m�N���P���h�(��X'���l��nrڊh��va��c�v{Ũל���vɧy��C;���g��۹�-r�7��A�=��ݶ��U��� yxk��q�o[�c+t��c���np�M,l��+�����I,g�������=�o�!ު����XX�/Mդ�vGiWVL���'d�K���\W ��Tm���:�r�(�os���M�͊�dnm�5�5�F���?_{�۝�P�^&�\]�چ�;��m���iƩ>�L�س])�����t�gb�mLp:kJ':��6��FG�g=��q�>�V�,̡��+e���}-�>@�����\�
:��6��q{i^V%����e��']��)��x�\��H���v6����s��U�`�׏�>�|õ�s�}ޙ}�4ۡ�<�=���=2�H&�7�*Q����І���8V�)c��F���;2/�9;�*�5)x�ژȽ{4Es��x�O�hˊ�j��F.^s<�F(kg�y�Wn �T^��ʞ�]����gN�Y�5Ʋ��O�a1�*=�����ҭS��oO'�Q���L6��B
�7y�2�k ���a���ă�И���	��y�LƧ6*)�����z�:�d�3ے-�����'���3�yUSkP��^� V���|}��sm���+3��xd�$��}j�6���z���Q����u�&v�j6!�����0&�;#i�k�p��� ���hv��o�YY����!�����!���~�^�z ��%]&�7,�v�4C���g�ݶ�����=��W������yfb��8u�۫C��▯�\��őƒ���D���gji�NMڲU+�46��ɡ�O���܌k�Y����5�o P�8۽�X���u�RN3��g7��:�����P�g�x���5xNN���JOu�Ѱs%�tk���]�k�q0�m�(�gO�[�F�}�2�����3�W�,�n���@ɨ��x��#wj��`���T �_��	��sȏ�w�ᩗ/&��牤�ѡW]��Z��+������s��U���G�ސ���	����{�"�crk�ݳ��sB�ۡ\��EPdcD?4�ᴬً�,��\���ޟ�9���= �E�SXGjv��M��C��O�bYob�o_t��]P̤�]��,���%�o���4&"1ݕ3���wV-Ȑ]u�/����2�n%Tȹ��m�*m��� P�ꡛ��1�Q�![���b-|���_��,���c�x`�ԯ����y�98�C��ۮ[���~���4�*�m�BPZ�l�w�ҏvh<Q��+����W�ݷ3,2g������]�\Y�r�c=l��l���dZ�=���%r�ʮ���9Sg�81�����7U�,����ޘ��Bccmi�j��㼘ov�1�Cq�[y]ȧj����j<X��j�v�l,f]�D2fpz�y�p���s��j�S9'\�9S�����+�j�ъ"�8"�l�LW)L���0�j3+2��W<�������Z������&�Y�n�u��*.�dkUN�l`���&�%ڻ.��gL��y����ʔǤ�Ớ.2F�չgA�h�x��eF<z���
5�M�ӹ@�W)|���2}�}�9�0jI?n(ln����
*�[.�4+*h�c�����~]�N��z[>%�6�{N�F�c	h�F�o8\�e=��Z��J�������l-�bz��H��m���3���e3b����|�왕u�T
��;{��w9��P�=u*qT�m�_;غ�q#��[>m"߫��Hx�k/�<W*{7v_�ɻ0Ц���b�H��"΃�̯�h�����#�F��`��ɒ�zjlHlz��N�C���i�>�!?y,SՌT˕;��k �����j���o�˺��h�lSHI��d�r��>�g���R
�4�̋T��ګXH�v��}�9K���/v@g"dF-oO��g�X$��Y+k�e�^Q���NB��{ǳi�y]���������$R��0oJK��;���G���A\��.�q�zgV)y,��|���z�P��7��A�'���?pr�'X��Vs��e�{�8w!�)������K!�@��nț�]6=Y
�F�Z����4,^+�4}<l�Kth{���̟U5�Mu�U���]<�^�#�Uw�X��2�c,������Q֮�RI���[���̶d9Ms-��5մ�~s-�3l��m�4�K���Ā[{�j�����=�g��L�"�@�&;��B�`�ݩ��e��}�Ǵ�޾tQ���	��]�6NHe�>�\��r��l�%�O��ژ�>�~odYW�LV
�r,{m
��C��;G��=<U��7���u�x�y�H�3�]{z�����+2���G[[;#�wϸ�*�ͪ��Ι�oM��a�b`k��+%GG�Xֲy]Z�y��v�<׊Z2�k�A1�Q��}���{!�sO�;�]5���]%��b[�*Y�g���V���3��o�{���ጆ;���d� ���@J=B�aw	�������;ͯ��k.j����o+��n�aя�恀�e���Q$��B��40�{��b��v嶸�mTůE��dRׄx���O{�>}c�
\�ۺ�{A��>�p�٠�S��6*�e��u����l�I�G�g:)��W6��P��Id�Pr*���z����o�}I��{���E�NV���y�[���-b
��Y^��!�IyN	�j��������l��숚Wu���/>�E� �oNV�f�r�G^b̖�6�M�Փu��ً�#҅�Q"�?D���[Y�'����%�殳o���fX���<6Y
��b�G���Oَ��J]�-��s)V0���s<��n�Σ�p7���e����!��e
��&@�
Xo�▁�r'�����۪���w��[7Ul�Uq>�cB�g&Ʉ�2��e�ٞz��캛��M#N����i��|Vʳ{@A����G���i��������f�g���e�7y"eS������U��n:�J���"l��^�h��P�a��Gz��*}j��f��+U��+{�l�}�dK��қ�"�ڈl�`�G�P���uN��j���J'�����N����(@�w��S���84u}�����)U��m�W^֊�&X}���P/"���c�mGpV�,�涸��@��[f�\��&�;
�åV�Kz��z�s�ق>�0S�$�p��ق��EE�IFis4�;�h	<�fd2�s��캖�p�̶$���qǛ( *v��F��}��"��P&�\�]����otb�<�7�We)EI����\%�ȗ>&�����>�)�vM�w����]�>��Ky{kuJWP���k���ۣ�LV��b�]��Sw/n:�@ҹY|���g!�+sr=�.�"�"E�%����e�j��.ma��Vt̴yC9<:�"þص��?�o)fͺ�@u��ύF6�ʇ�Μu�:n��sR�G��&��t�Z.1ܚ�]p�A������J�t��b�"�O#5��Yo��hX��ū:�sr��F�ӑN�ط����V)��bm9(�q�[�{�r��~Q���k�"�W}�@���Wd���gFĵ9�Y�i�[L����1܏X9���������)�Y�`�T��l�����ҥG���ʒ�]7��5v��3P*;�L���2컱;�8�CC䉮���}��7{s�v����q��5���CO�9��� 4������n
�q�gC/���<T���k��Y���f;��-�ԣ����E	Z�l�C\([����� �k:��q���CSʕ��3NoSL^'��I�ER�v(��r�kiԼ[��<l�H@�pi\�	=��)Sn�BkbH��B��pU��.��0�0�u���SѸ�6+P-�T�����PGƦ��9�|%ol�J\�J�(L5)����{y�c#��Q��7d�w^YN�1\q!\r����P�9���r��<C�I^w`2��c�tSsyS���ww�VYn��o{��bZu�r1��a�Y�������7�u�n�PQ��.��w+S%��7(*W*�c/��ۣZ�w�VM����*�ڠo��i�/�R�/��vDYg��E� ',��v��EVf�J.��H�Z����-�ݤ�2�cYt��s�xeK���i����v�ظp��rtw��/��u�ˮ��B�<���F��!%�E�5�իuGU���
��ͥ'v��L�JΜJ�%�<�����Ϸ]�Y�:�2w|���2`�M-np/����	�r�$�YDl/������1���%��5r�u,V��Se�i>��"V�^6��*_[&�w;
�5>�v���:�t�Xe��ڔ�(+Zn#&�1�����yWs]�\���+)k��ޙ8����Q䳨J�7.2�L�+Z�I�L�evw!��{�t��g)�Z������ȹ��씫��[ÛY�'-�U"Z<|������r�ֱK�#�ĔEaڴ��x	���[g2m<�ubD��j�Jeq�^�\��|�w����;��ʠ��)��S���mQQ���35�(*��E�U[b'���}�>>4�Z�b
)bcY���j�דȪ�����媦*4jx�����MEAUq�EQkQ�`�(�(э�MPQZ1�������h�QElV����5�*&j �X���J�(֢5�
	� �������*&ō���b��=��(ƭLQ�����I�"*+lh��M����ة(��UKF �ش�c6í[QV��US�IAkmY�mgV�N��h�Il�5�EI�X�V3� ��,juT�����I��(�TUU5�٪4�v�m�SAQ�V (�Q�ӭ� �EU4Rm��E;
���hձ�A�c-.&�(��b�h�Mh1ɝ�(j����:���c���Yc&�M�`Y�lt�x3���^ }v�`So��D�3:ĭ�m��
)�A񭜸#U~�5���ܴ���ta�}^a�����tF\�w{�w�j��I�|�d�ȮӒ7�A>�١��Ĥ@��$�3��$\T�n�j/݂b��#�q�b������A���� o�i��B0f�=�իO�|؝��Ue'��+^Q��ȏ`l- �"J�!�����I���2-����x�<p��8b�<ҧ�h͋zw��n�_sH�~�K�{NN�T�^w6U�N��ZN�\0{��N��"l�z�32_4�����]mk�K⢶�`���Nf��u#e���G��=r��4��j���C(a��M7��G*0s�%��3U5��n�F|�p�H{�t����ڇ��k�*���V�6R�n���&㲀G�w8+w�P[��U�p0�n�ǭk�]���CJ^˳;��9P�H׊��MϹU��W��N�]��S1���f�ccC/5��9eE��4xv����;�3������}RH4�� 2$����=nt���3�3k<���fT|���&a��В��q�;xwt�ډ'�n����N�*J�@l�\�CGBCIR	(�wӖ�	�Хd�x�;��{���{��Cj�dB+���~m���Ϊ�Z-qU7��^;-����p�/�v��Z���-��]B��z�<�G�� ns����.%�Ҙ/$�c'��ͣ4�ex�ܯF�;��Y��X.!k\rǺ�d���Yp��s8'�f'v��0�'r�ΟQ�h���w[���1,�U�^��_��Kc��/:���֔*�]�/Ξ��{}M�!�·8qٶ��e�o�ca�����{���ɏnK�n珖Q�s"��^&x�SX�f��F�}�IL�˯����2#���=��y�ՐO_P�Ͳft�dnQ~�a�E2�h֚m�Kzv*HJ3Ұ�j���Wf��c7(����2�k�ח��ӍK���m�˝�c�p�����qȫ�f�/ݧjn�sD�j�ܓ�˩� q���R6�d�x���f�����4�ͤ����0f���2�}[��ʔa�� b�І���w�]na��[Qw�E;�ܕ��u9�Dx���me_F���Xػ�i�E���v���V1��J)b�㥣���\���8��:ᴞu��T�������UϘ
�\��B���/r|!@�HIuo	U��NИi,	!�æ�H�$m{�d���<9S��(x�j5>9�դf���;�f��l���y��%�#kP/�!�Qx��*w���g�]����e�W�,=������x��WS��"�YW�$�iY9A�C%��2*�FFI�y0k�=�}�ɧO�.<�P�er�[��
�+ ��a��4�9�椤aL㹛�f[N��Z������p?�_������g�����Ǐ1V���u�T�)��7����f$ڐ����5ȂH�Ṝ0�Xz�#S�#�tpݭӤ�5e�]�1KM���~+t�GR�;��3�Kf�7��y*�Kڻ�+r�mF�7���t(�:\��rR9.[D����9�5\	}����w_cCJ�U���N���=�L�JJ��~�-
l��k��P7j���UN����+3b�\��3�������Ҙ�[�[��{M�͔7G�$׍	�V�wX�ʻJU�<�II�n4�1L�K� �^M66j�&̷򭆃�Z�~�tO��Vo_���X}�b���טr��+�Q�83{��=&X]Bp}��q��q9<5S�S��QV��VR�8�w���M��+yd������K�x�
dy�Qђ�:xׇu��N��D���+�T����)����/^f���>�R��*p����\�.!�^'],�W&��˷� ^��Wj�GHn�G�4ÍvXRٷ�*��	<sN�~�����wv%g
���:��4x@�FCr�T:L���˱U��+��ǈ��;�FVJB'/h�l������D^w5��+t��u�t�ԩ�AǄq��=Ol�ÓJ��􍽖�&�p�<�+U�*������a4�r�7{׷<7n�CO����!�G��Kک=M5:�jY,"��n��M������s�����O��v�� ��>;b{��~��Qr�_����j��\�f~�nJ޴��bݠ��:�e��j����DI�V&�)Bu�g7sos��oH}����8�M�U�ꯕ\P{sx�Z9������3��5�����7k0N����R��ER�Ijb�I����n�'U��_ِ������Ϲ��J���ӽ@��TE�̔��n��iqM��� ���]��n۩6��[4�)� �.껛����P^p�t޼&��UU5!�nw���{ph����G�����*�Iݾ+g���y༆��6�z�D�h�9�4�+�<֮�ţ��s��F=��Q4����[�!��I�X^�KP�j�u��V��nh�b�5>g���i�=��Z��y@�����kYLn��lu���^J��X�Q���d�����F��?{�nz|�c&z��������w�-#؄�����G�����S�D]\�ʍS��t�\��ZV��]�B��s��8����n,1,���7��g{3{�u�D̪�2�2Fƕ@���z�Ux��M�����4�CY�/����h��g�e|&�K�܈jE�1��y�{�,ԍQ��������=�z��k�r��I|�v�eI������X���l�T5Y�q���?ۯ�]����HZŊ$���{�����l�Y"&����܄������u��T���}خ�o�Ǆ*�</�V�HU�jǼq[3� �f�\�#��U�Y�;b{�����?:���!F��Ѳe��*�؜
1ݽ3t�	���M͋��/z���Pk�fE$��l�Z�6�m�|(o�<.l'��^�aϠO�j���;�E��(��"0tS3	���ti����7�c��z�ɮWa��;��Q�����;����*���3���ˤ�-��c�Ǉl�����	Ŵ̪�����D�dol6,��K�[h?k_)�;�q�ǝ+*8��n@�V���䫞aWU�Vf�zl�jh��Z�;Y��i���W���K�Ҭf�X�=����n�t裙/Dv�\H�u,��_�c�٫P5��j~���˯�]r����9w�ܭrXT��-)_:.Ou�Y�u����5��������&~���oүR��Ij/��%l�<���m�[�:�hzhr��nR���'צw0��P+��˨�%�v�|��˴qǄx�騩"{_7��6'fLE�_����vR����&�_M��6`�����x�����ڲ_#�qĐK$
������[LY�:�F�*� ز��F�\OL@拁=��*�x7m���5o��@ܵL-ܡb�d�=Ң���R[]
��y���
N��t���X�qΜ���rc����VVBʖdL���,�՘n\�+�Lܫ��2�"�##JhZ"XUj�ȹX��_=�kh޹��d|J�zr������c�Z��ybL�OlSq�p���J�L�Xn�m�y�;�^�c��w|Zb�Ȃv�v���GbH�����(jK�6v�
�9F#'D�f��Ϫ���kq�]��D|�ݠ}f��s�<ʟ�i�{1o`�YB[M⛼�5��{yK���$�c�e����G*u>��K?���a��^��R�CT�"�T��;W����2�	O���(�Ky��E��]���*Ӑ�:��ڱ�M�����[@���%sۛ�r㌟=!!�s�w��3���zms���g�\Vm�~u]�g�u�5��g^=�E�3^����݁���I^Uo��h6�k�)���zU���ԞX��wK2�;Ks����on�f�M���"Aݩkp�;\���+����{,����mÒU#�Y ������Vz,A�1���{���[r���T�5��O����ݗI^r��a�Pz�5Ѥ��� ��ռ���m
�<�"[�/_V�j�u&�����kU�ʋ/��15��n�����{A�=[�<�Rw56�mx	�v���h9��'jm�hĀ��C>2[MP�]S�w;��5���"R���Vѷ���I��a$[�����������Wl��UV��u�x>����7eWa1��**���OHK[[*!e8M���Y1��7uY�����]�=����\9��\υ�8�����u9u�r�`]N��+��0�6�b��Q������Ňr_t�U;�e��<Rm�)��m�G{L8�m�6&
���$�
j�C�.ȇ�-���[�����s�r�w3ș�C�1��d���{�g�J%�+�T�f��.�]ӿM�`��p�u�|U ��[�sdi��<��M�����j��m!i`�31�56���eWy�#l�7�\��fJV��+6v7ݞ1\��
�:���]��/5���R�=�S�2��.�b_#� ���U4�V�h���<y�:V3G;�ů�M'f���vq��<H�i�Ř^f}��O_m��b�:#���ҭ�\j�H�1�L:�&��L�2'�S��)��\�G��N���F��k��e)��*9�AL�������p���磅�2?<��t���T��R#���v�Ym�'���5_��t��o��7�mo�����f�����EHHǮ;.c��4�阩��|��k�� o$z��\��=E8��î����$_k����ͼW^+s��HUo��.6v�ɺ��⬟+��/SLc�{��9jn��9���f�zu��j�5ɤj=-�Un�?��*��P2o#S��鶘�C��n��5�}�U�B] ^ #����*� ���q�"�6�|2͹Ǎ�V�\\%�8�gdt̲�jz�tZ��=:V*��4�s�ҵk\wS�f9*q^�C5�	Y���WGnn#O�)O��orU�o�/I��ˮ��ŷ�b�]hCb#6���he��Ř�k�B��͈���=��'��{J]��J^��J�����4y�p-���j{k�%��2ξ���,+eAԻm�]�3LW�7{e�v���WL���YۜBY�!���՝x�	lo;��}�ܿ�)^�>[��:v�`6�]���T%:�x�M�f��˓ul��=��vv�o���E!ٽe��W�U�K��ͭ�{��~��J�r���ms�+')��_D���[KV�˫
�At����m��3z�pmPqH�V��s��T~s���u���tO��/ti�ᣨ3�hf�kL�	zV��Yb���E7=s�:E]�-���r�dJT� ���݃�� g�]�J�7W�wr�N^camR0OE4��gr�����1qi�4ө�l3猀��7'�J�o�����t,�ry[���"��}���!�[^%em�0���w���e���ʒ���[dUB����y�p2�M-5�ί;�S�'lY rX�}�k��fh�t��f�Ϳuk��Ȋ���C�.IzXd>�Җ�ҩ3�7 G(������{'S����%_{��D��1ԙn�q����lrW����j����Ґ�S��p�ᄝ�3���s���x����m�ܑ�9�Ft[�[���y�Ű�v�;)�8GYrt��᛼��o	Us*�(����7j���H�+�r�T�(���I�u��mc���-�s.�>�s���F��u���nK�a�jͮ`]�Q�0����2����{��Zm�w�wGSS5�2�R�S|Cjj7X�⽧�Y��M��[8�[�
�zu�Z�
�P�ʽ�,ڀ�{z��K�.i炎m'��H��	,�w�v]�z��b�o�I��,����H}pI0=�k��]G�����T�j�,���؊�ZZ��Yiݴ�W��>;�6ԣ��]���Ö�ggn�y(ZW|Za�}Vsf�D���j�+;e淂i.�drεỹCTl^,��P�/g+Eչ�A��,Z���5�'p�xB�j�
T�9$������$�I�ܧßێ�a��Z�c���Sv���u>G���b�'KrN�Rn�l�@i���&��e@�\�ŷ� ��n86�B���aV�s!m�n���|V��/q>:�B�^qѵ��{zR��t�v��m��#��r�J�O���u��b*�r멝�m�lۆ�);Y;I��Ŝ��g��▇�'չ34��z����cn՝x��C5N��j��f2��v蝂��0�؆��Hʺ��#3#���IKF�8���x�#Fm�j`۾�VM�(Jܡ��,�	��D�]g��lM7���{���h�c�˜i�+_�N��KD����Sq�B�6*K��ے<�f�=����C(���j��|��d3u�>��-f��.�Z�1����p��$�3Ƣ������=DK҉�D���=؜'/)bゐ�Øph1eR��!R�qWKH��{xm���0�¢;0E��J�8qx��]�ȵ���<V��)]W�������_Ϣh�yn�a�	���;�j8Wn�]�oui��������x�+��nV������y�;�:Xg�k�8�-Y���1. ��*�7O�N��[���Qe��@;����S!&Һ#7#�jG���Ǯ�B;���L�Rw�A<�Z]ي:n�[˭Ǣ�$�x�OU[�^M��1eZ�b�y*�&�o}���>���]��t0:��1^S]8{c�́\�j�f��.�qVH�T�gk`�+,����ԉ�.+\�$^^���2�K�6d��$���� D��qb���+�n�
ɋ�IO��\2D�W���1���cu�h�ctH#�oA�������!nP�#;}P'� �r\Lz8�_\��9L��z�X�"��:j%; YӾ�.�9��-�!�R�|��;1�ځP5�i��������ȧ�U�k�f����V�M�1j��=`���Wv�l��c�w�h1b��(���m�*�oS�J:[J��j�����z�;����y�.�+nm�u�5���1+�[Ky���w�k~.��WQ_S��2�e��
Ak��F����+X�G-(��r��Wl�l���b"A?�2�Z
��Z���E[l)"�*h
��'���O���PZ*��(kF�Ui�V�(ִM���v�4v��9������
���k�l4y�P14scAZ4њ����ր��NګA�QG-.���m���-(Ѥ(+TUS�bujgdщ5C�c�����Ƃ#�`��;�\TUAm�t�M����N٭�Emd��QjΨ��F�mQ��H��:�'V���EA��؈��@PZ��l5Al���ڰi)�)�Ō���N�hѫm�U���1�Z-��ڶq&��51i�`�l�E�A�qh��ƵA3ZB6(4m�E�TPbѝ�v3��6�lִh�t�:�Y�b���m��P�Q��!CBkE8�&��cF*XѪڈ����II4S�� ��%��o�l��+�ʞ���;h�NJMv���t��2�Z6�պ]��>G	��U�}��c�\噒���8����d��U,���LI��MND�m����j�GO�y�W�{d$��|<���G����"�9�b��b��ӟ�gg���{	�A.S��Ɵ�䕝G��6�y�m�^���A���Su�ʫ6�j��@�3��IAEv��f[t%�}��۫d�}����;��`ߑ/9���s����T�������!h�Ӿf��W�o�y�4]T6�ʼ�Oa�\�����/��O��;��s<�wM�ma���H��80�ݾ���@Xg٘db��;���"�Q���ǘ�ݕ�?}��s�?�|􆳱
G�/WOϑX2
��WNY�)�pʚ�����ͯٵ�u��#JX�)�lR���H����2��W]����9tf��F��QO2�	7��*u=^lR�#�mc�?rv�ڋ�<+-�J�]"&��dP����m�>j�^��ޯU�s�Er��ͼ)%J�ue��4�,G���,|n6&�%s�ٹ[;#yY/k����������ј�!ulv�V���$i}��u�o��,���k�<�Nε��|�^��<n�zZ�ԝ�{;��)`�Uq����$}A���7����P;���L��ԲE>�U��Ҫ�xx(uN8��|Ν�������I=����g��<̃��.��J������Qjz�7u9 �^�sU^�+�+�.�3�2�H�oi��)	��J���pfL�M7$S�٦m벶wHg;��4f��[\�"|wjX�����-�zM�����i៮�z��I*�$��p�X�GVd�[���/��r��3n;V����>���
��R;�q�])��ב� ��
2�݈����X/q~3�\g�m(�v��w����j��[�׳ٍ��;R�f5��b���Pfu�׆�w"����4?����cgUuG��ܭ�5����߻[$w�a�;h�+�Gron���Ov�%xA�ޑ�I����7^��#	YV���m�m�}��q��sF�Rb�R[����f���nL�>���*Jv�x���2�
οy�Oe�~AlƦ�l�@���K6���,tF D�&���ɷ(I�r2�_*���,A���y{1�T���D���,�b����G��X�Wm��aA�9|���RĦ��0hَ�ʬ�eW)�I$�3�?�z?%��uI[��\џ1��G-!���8|ҡ~��\{�9���㑱�:��Ry[[?ʤ��Q���H� �C��'l,n+��=�������-�g)�M��1���ͼ����kRCKdŝ���N��7q�^SC.Me�������u\��0�'	y�Ò
Γ3~�B�-c��)��:�v7r��٠q����!�@b�C٩�t��ׅ��k���Ӑ;���E]���p���a�U�X�-�h��9���^���ن��+�;�nHi�9��~�V�$�Y� WU�8�ot����(%f+��ӻ���/n���/��n�Y|R&Ϋں��m}��6�ڕDZ[�]<�ܬ����&8��.�4�G���U{L��Vr�����
��_�s��/x$���@�{��G�i��]�y-&�V�Vɭu�D�f����7"Cpp
�u<&:%�ib���,h��dL]Lu�r{W�i�fL�g��@�<7���+6u=bb�C����Z�Y���v����QT�9,�*�mB5Im�I�QȞ�2���"�[+#���7J���ɘ�HB�?	m��~��r}��vLڸ����9=Coa���,��oA��HK�.��{ �3�`�2Α��WX�؜Os�uڞ�ͬ��=��CdUY��0o�㺲�Q"u
n�7�y��ZX�a�y��V��Zv���W\��ܞW�VW��㾣�uj�<�mW���6��G���O�%�3l���b׊`3�s��5��쏮;�x���j�o������1I�_�y����H���G��5_c�n��|�7����X�I�}jA��د;�>���7̰r�X´Z����}>y����$@�L��%���.CNobc,��x��wH����5^���y^�k�ܚ��o/Hm��r5-�H��.Ӵ4�v[>Pe-\�4���J��YD��V曺�u��uf^�����W9��b�y��5wY�~�Y�}.���ٻ�t�a�?�oV-�dv@�G���i/5�q��
���a�j���D��5�]�-����Н.a'��'�A����p;B��m%��Ps��fi�b��ے:�l"�n�ì�jup�]j�3���K�v�xv7�Ȧ�P��E�BV�85��ٷE���PA���ݾgr���������;=��uB�� pr�x���˙��vS��0s����9gi��d��[�ajXi�8��Z�+��y�����{��.�"~��x�W��|MN��/���o�Q��Wh��X�75n-�Sp��k_Mg]gt�w)��ئn
�ժ<79�-��6Ɱ/*qo,�y�C��y8�.�IgW�"C�pafڃ-�;l���S�-9QK���2*H�.�݈Ò�pO�Ge`%gP#������*tc�dm�9�5�'e/Df�
=�f_m��t��*]�H�BZ�Sf�3=F勼��f�����NoM�t����sC����uP�ܖ�ނ@)�3�9������:���Sr�V��`b���?�|?g��Sg2Si��ʱ�O]�%�j�����3ܾ�C_
Θ�fQ4g���/y�L��f�>�1;�p8�w��Hv�Ƭ�1C�:F�n����1�c��9&�pf)ěaN�Ա���Y)��n��WWt�_y��ަ�/m[���cN_m�~�hz���N��(j+�&]ڴ��*vu��j�oM���G�R�ΡI)��ּvu��j�7j�l�wT�;���=���n��F�gK�vL�u]"9�^[CrHVgU���؁2g0푺9֚$`��HcL�a�K�C_;I��-���/d^��z�j>�o���RH��w�IDd�e��۔�����f8���s��M�m��5*�ò"ns�4{B~�e������K+Vl�;L6�g'�r3=�e��Nc_���<��P�š�rW^�@�Y+jxLs!*b�?3�Z�9;�H�)�7r^qқ��e��b���י���o��o#c픓��}��I5@����;�����QV�*�h5���
h�u5?'�Q5~�K�L������weq�h{�Y^��e�W�'c�B�1TH�t��t��DY�70�Ǥ7$�hY�V*���u(��mRᚙ�V�SUc�OӜ&����C)o��o���\lI~ܔ��CLN�<lTlv���"���-�Y�.6|Vi42#8��6ue
�<��N̮�V��:Z͂:Z�)�(p��뛛�u�_Sf�{H�Z,e�4�=�ڟD��yt�Ok"��wLo��68��KL��9�����X.�䭇�t�:����Jf��bN��un�Q������-����B�>��m*�v�3p���I����ͻq�k9�~��_$%���5���~���1׵zn��#i��UE	)�l�-��Z��8�Ӎ-����03hv+�Gb5��/j|fܢ"���M\ᓄ��٪8p�qՔ,�l�3� �n��0�a�o46(J_.��MӶ����{Ǯv��
��4qa��O$�I릑��h~?_�·���X��q��M���ݸ#֯E��1B�Z2;��V٘�`Z�؁��'��g�m[ͻ����ato44�Ikǈ�S��@`˻j��\��&����������gwG��@��7���!L��K?�'�@����c0��a/\ʜ�͙�<,�Fh�9�ٳ�?;Ycx�T��L�D�m�O�ɧ
�z�q�m����G<�''�M�UC;�KlJ����:Ϸ�����l��u���u�l����(�z��W�J��e��h�P�#H�b�um�Oj��3����MRD�[Pkei��4S�����o%�Z4�m�ڕ��a.gk_i�ڈ%��ʎ���2���Ik�s��&�T0Oq��s��3i��=��~]keuY���ͺ��]!��3j��Y�{��u���iݦ��Py�Jح�:wa,�)x�$w|���N[�H�͗i�ՙz`�_oEK�w`-��5?�K6H'b�q\Z=ڏSt^���+c����C�<7-�p�N��mc��k�&+�����`�}��Y���H�u�1!ś��gKte�Y�m9N��ݮ��oo�yWO��Y�g��(Wכ;h\���Uw-Tq�y��O��%�f	��C�r����nfj�j�����5��	�F��.W�w�wmxb�$gG�`��c2�I�tc�[/��F;�i1�c���b�H�Ȥ&;�$f�ؚ�`�f���LY�V�mYZd����`U��RT!���u �1:��N���͕*{n�3��g�f�Ǜ`2M�n�b�7�s{��ϨҘ������Gy������] �N�*�_h�SqFn�kʳܭ]z �ߟ���V�S$U��d�At�6�V+OtQ���>�vn�K���Q,��^7�-�nL�7�ȧ:�v�6�+�EJW&'l ڛP�2ڋ;���ώ����]Μ��?���y�t�s��xw��@kQ��$���ʬ~�~�a�s8�4�ם�M:������,@�I�ڎ2�7C@���L�8����unD3��s��kz#�^�r�!�k���F�u#���x�e6�Gm�l��v3���͏�F�������%�Ga��,Ӽ#{��j�y~�\�V���߻�}�h����RMO��S}CT,���\�qm/ٍ�9�Z���������>��M������V��xb�g��%����d���0L�����H���!�߾���+�7k�j>����U^��ҫ���z�$������F\�jKM�qM�UW;�yb�����H�Y�F�r%r�h����[}M��}��ͯy�^'rA':������f|�y�.��˪�}�~�{�f^��\��W�nP�ts���.x����j_�^��>�u�t�U��D�٘!4V���s�)ǻK:).�����)��[��yW����Ff,l�SB��~#:]�2�'@���*&��TtV�}�f�*�D,-[�(��J{��|��7�},s.���t�^Jz�f��A���g��[�CnMqN��V�P��:���>#�n�r�2v��-�P5lv�}��v����,��bJ���T�tfd�C�jz�r�wo~7��=���i�(h����0#��!��h,�yӇ"r(;J�"�p���5���݃���ݗt�#a-�H�9�C�6����n��;Om�q�|�G�4�D���6:r ʹ'!��0���wp�a��U�����yku붉 JCe;�C�-h�e�s�3ܞ��[��Di�����]�ݗ�����(�%��v�.�>3kYE���f�h��aZ^&1�T�Eｕw}����Ha���j�=p%'�Ωy�˨�ծ�U�ٖ����L��UƜ�DǱ%�/P+�ac5[|K��iw��:��yD��Iʡ�ݑ��)weQ�r&Krqkx�	���M��ƥn���<�!7câ>���Y�JY��,�&��ٷN�cW�q�eÓ]��c	�8D�5�c���LB����W.�X��_�t&�t@5�����d׊��ם�h�B��V�X�;�&kO$��
3B�s3�t��n)�Z0˔r�u�n,eG,S6��L\x�Pn<�$�\�y{kb�!`&D`l�h��j��Аe��_)��G����:x����h���ؔ�㙃�ރ�Ky���R>���/��cc�P���3��V��3݂�&�7.��C(ϲ��'R�1e-�툡��.�yf��[A�.���M��7���۽�}��CM.�`��wK)m]K��{�j���;3��z��{u��7Y�n�pa���B�jϖ�V��Z�����pV̴Q�x١I}�ˮ��Y�q���]:ssR�W�:����� �ݨ�Io:\��Uw�M@�!K��R��(����lJxx+/�&j4�w�ݝr�[u�L�>�I1��i�;z�r:,[7��aƵˤ$�
PV���g�ިf\�P:s�]��)� S\�R\�������M�X19�D�t��)Z\;�ǲ�;m��������ԫm4y٭}�خ��:)`[�r�Q?IxR�I� �CW�θ��Z8D�����B|�M�z��Nf��6e�%���hkT.�e��k�dc��QA͇���ܧ��"mt��la�Us��y�B����W}�M� jKU�.,�ī�v����:��J;���6q���f�J��X� �<9[�!	d�ٙ��ś��z*u�R<쬲v ��L��Է�k$��W=K�Z�f�3����n'��`��c��%S��B��G��}2�M�� a��F+��Vf�9g;"p»9�[�]u�P{�YBHֵel�&
�apα��?��ޅ��^�Ў�P��l�Z�q����Qja��Ď��A6�8;G8Of�64E�z��l:N�;{v㝌�}�(/o�<C����|��D������9���oo45�=��Z\n���;#���P�#ۑ,��ח�k�1ɣ͓����:�a�uu�0-���ja"B��z.vݷ�̌+�k(�S�%3y|`4Y���9���	f�Yu:̣�fv��낥�ř��H�κ#E�[p�]���z)����c,�:�m��fVe���wk��8�O�B�;x�ꊡ�λɂ>��J�	]�*Z���sG'wi*4��ü+V�4�
�i�� Q�V�Wn!�eA��c����4���c�	�`�m�;9"���E3�!�:]N�+2<1mW7���C[�CE���>���7��y4��R�,�n|k�\���"��6GQՍ�	� �o]�;������ �nW �r���5}e�<ki�6��5�K�}O���-�P���_ם\Mw~~z|����9�m4�X����t��!��l%:�5U��֪���k g����||*�������1VmQ��Emk`�@ɣcS�6uSh'�����Ȗ�B#�4�m4hӭlm��j�h(5�*Ɗ�>DQy���
j�14��,cm�(V�"�gMhՍ����<<<<<=y��6�V�l��jmQlX3�5���6v�cl��cT��4lQ�F�v����gkjkY��"��KÊ(��b���A���Z�kTiqM3�SE���[d"��m6�h�Dm:�h4h�&j
�"��J*)��A[j�f�mE���1�*Ѧ��%�F�#:0M%4TŲh**��ض ��Fm����Ƃ��Ӷ�kVڡi*�kX��h�[��&�UQlkZ��N�M��5�ҽ�" ҏ��z�+�9���#�t���W1;�I���ҤK^f�V�Z FQE\�+�
W:��i��\������)!����㽿�s���>q~Tg
��V�g�_M5�,
hO��9�S,����˫���N��=Ý+ԗu��T�U=���m�ss�D�U��ͽx�HF�-���u7$��'��edyWVP��.�q܍ݭ�SY�I�Z�\�s%M��ng +�q,�G��rn�����+ko^vHqs؀���ӓ�8����J����t�9��U���?l
5N;�l�%ew�m���~��1y�sM�J}������T��!GYۭz<q��@�fǟ=��ڊ�Դ���M�WvL\�A�8��'�е����6�=�1�ᷚA�ņP����s�[%��M�J�������@��h�cA�3��#88�f���Ս���u��@iO/��X���w,n���<lG*$�,/ �64̙�L�lײ��8�X�,231K��g�j�s�P�{�C	��I�j�<wk���6o�`�8I��v�TaL�q=��������ygG����w�����}���[]�y�h�/���t<r�����CR��2umh�o���٭�YwV^+����m��<��)3��՚Ղ��c>U���v��;H7�ĉ�m�jm3獀�a짊ꨭ�/f����2W��o�-y����5kE)�M��*2}�ٹKц��R�g��&S��e���3���	j;-d��x�$rkU�V(�DO�[c�Un\�w�i�C<���ܾMmQ�v���ۛ̀�V� �ݥU=fr�tX��d{7{wu��e�!�I�&~<����P�K+�\�d���`�:u-ͺ;�}�̪C[�lr���Šn�=~�aB�|b��~|��5SG�k�I��!�%J	nW�����YÉq�d��i���w�ݍ�(�$Wr�:7�Zj�Ϲ綉���6������\=�;��c��5���j�(�YUxv���9��&t�@QD�˻�1^ώ�?��y�a���OA{�bÏ�FCJ�u���I���j��z�{��7 {<i�{���!<M���p���,�Ϲ����#��,ȋ
}~݈=��2Sˀ�Y�C/��s@\3W ��ێ��Y�f�m�I�nM�I+5�;���*�oaF����EAw,_�o�y�!�:G���U��tI�vu��]��ߙ���c�u�p
��H�Af�ΡM�ocશf��kd���w�8df&^k�1;�>w.�ŉ"�HE����Yi�t��@�s6��m7������Z�6�nT��u�a���8�:�7Z�Ué���΍�ȸ ��c��(�	��2 +3b�qo7^w�Ͷ������mhW�僌���Y��ȼ�*��v�|$�ku^w�g����|�M�T9����&�m����ʶk�?}�k�����~�/3���љQ�T�s1\��E�l�P�N�e���m�p//~"=P������u��������%3�����
����T�9o0�q�YE4ms�Y�W �(���{���u5�ח(תo �?���0�d�e?{fs�K�Ħ}�k��Xz�S�ʮ_S7�C&�Q�X[_�����f�����w[�j5�p���O\�''-��F<I^���al�+ ���l��C�������ig.%u��:��c��k�����H������N_]��\�@|y]�En��s��L���"nt��]q��;8��˲���u�s�̳�e�Ėk9�����1WcJie��K��pq��B�ּݥ�X��u��0�A��V�%Y>Wy�=�5!�W�'���=����L,�� ]�jﷷ*mԬ����Ƌ��`%�),�E����!���κظ���-<�n�͑:މ7�s�9)�:|�A�.IYǙ��xr��_����)F�7�ɍ&/�U��!�LBޡ�; n)�]��eB+�[$�-�k6�S��њ{���i�}�=��Ԣ6�gz�ܕɼ~���|�;{I���Mt@����?jz��|��$g��f�k�����LBڼ�Uݭ6���5������;�	F.�g���]]y�|��>�E��]H���Q������]10o;M��l5��Ne���l��vL�.Mh���#��*>�hd�)���m��s�xX�?\I�P7%�D1�g�D6�ъ̈���/q@"�3<�bw��/F-���"!����k�l|k�K8�\-{sO����X���O}�?i�w2���9���JTNJ&�`�A���|R��[O,g�c���F�;�\�k��d9���;\�
[�2.�t�bZ_t�.����|��\�����ї�����p�xy�ڧf��Ѥ>K��;r�]��n5������ԪDYS蛩�VБw��8(��f��ٝ�B�2��0���<u�u�.4�}uވU��^��4�D�$�Y��"��%k5����i�К���Id����S".��n��\�}9�)�؞�]���+o����{I;@䝣�����(�xx�'�K5�x��eV��nn���2���'�j��;BYe�����[\�"N�T˅�i�����"&��1��dY6�@�K���%~O'v�X��{P��}���F+�j��D(Yג�d vb�J�n�\;�q�K�U<�k�mC�v�r�"��̗M��TO�gH�]0����S�z2d!��(����n��u5��M���6H�fv��f���Hi�zi��y�Y��6���N��JӮ�OkG�:$m ���[�s�o��`���Pf���i�;=g��5��<:����e��ھc�3}_j��JZ0�ʇ(:ɷҴ�]y;�srh�{W�����y�GFOd��:�7�h����C���	#�q�s*F/���]m��*�'�ռ�������4�H��|C�]v��lܼlA�9ǲ��L�\���=ܲ�<���m�fv@&ۻ�q�����a�'����^����#k��3ںK��<��i�Ӗf��sa� �_�w~n��q77�\g�Ӥ8�I�:��*=B�^d{H'�&�����"�n&5I��py��*8b��:�i��ϡY�/�X2���㾨�h%b�:���c�@�=h��b0��ljmR� k0�?��"<gp�U��(�gǊ���T���{x^��ِ�O t5�s���=�/p�p��2UV��әYo��	^���'V���jn�UX�ߡ��U9��Ҩ�]f�m����2�'\t
ݕ�4��ITfH/^^,{W�7S�'z5Z;���7�7Z�) ֣*��ɮQ,2�#v������b7�v!�����M/\��[��jǿ�#n�������Wx
���,\��� wB���B���7�5��P�mm��&�V{�n���%����e�G�:*5{��K�#n��I]a��9�y�K�[�;iԥ��'��򒑪cBL�DE闟}z&Y|JfE����[�	�o�e�װV�wŧQ��t������ ���$�#�'ҶM���[��G����������G�B���ʾ�j�����K���ջ{�N*��l��2�ռb�ʹ��V�k�T�z^v�i�֩w%l��دO��48d�*���������-B�~�K$;�l%�d�'�V�*{�
<!-�q�o(�>8�ɞ�}���Ik��@��·���B����X�-|�"�#:"�l�w�&��3�{�(�`P�i���0Į�H*=�)�i嵹�	["�S�ۦ����Dt�{v�t���ԁ��m�P��7���ɸAv�6v�U��z@�w9O�3Z���,h4����"����^�3�Tי��[q�r^�M7��/�#xX�T�|��e�M,T�P鏨$���L����@�qԽ��+�^����V� ��ΰ����;�[!��I[��cN�7Nlڛ��]M��(�g�ڊ�XL�Fbu�.,8Eá�zc�P��%�ok�l�y:�t�p�|c�x6u�C%��F����Y���A�}�n�s;�=��s#���$E�o�����am;@�N�e��?M�y��3o�m<C����P{t]��7�Y��͔v����mBK��:��@�Wn���m���kҝ���i����,U����i�8�;%�k4����7�iZ7r����P�T�W/��BN,3���7s��,�;?x'
|^�}+��O<�=��y��U,��T�[r8LiZ&�xQ�39,Ѥ7j���YT��U�W���Ƥ5[�ս��]��p�#;2�M��f����qDr�['�Ē����楀�s�^�u���j���_��~����s�<�W �,�=o�%^�B�P\u�=���Y�ɳ���[f^ύK�1
����b���#��TWu�\�����Y���숢H�3���U�ᯠ:�!�Ϝ��mx�s;��HDQ���N�ϵ	��)�oV�99;L6�kti��z�n'z�n�ǳ�q��Ln���0ckd(ra>ݵ[��d�(@J�ԥv�o1vь���;v�Ū��֟h8��.R��ګG�i�%v�8]mq�ǝ��{8�����"{�j���c�lN�i���g�[G{6�y��3�ð��m�G3w���O4��$��.^ۅ��u�>��g�g'��t��ٚ�̻�ш�f���m��Y�~ϳ!��"bW�tż����0��=y�3]-T϶9�&`k�v�n,I���.����\����l����d�$X��������cv8�\?,��}�;ذ$%� 2o<G(x�V{FfKϷIQ'�`J�t�3�E0g3Mi�ɇl�z:3c�J��|dA�e�WbQ�2��l�O:��[L�q��,�f�'cdi�R;e*�5��#y����,�T'�l�i����M��ydoʖO��ox��J�/ԓ�tퟩ�f}���ׇ�d*�ʼ�wWlKx�;?GU�Y �4�YA+ʢ�⭖�-���h��k����:��׽lQ��P"��
�7��В���c&�Ӭ�� �|�m�qM��y7���� �ɺ�W)1L))��Sg���;�Dm���nuv���1�`�ۏN�����9G��"��6�+�u��58ps�5F�6�k�Ν�����}-m�Dp��Xf�\�qӔ��k����zLխ�,����~�ƹAlH�8�CrH�y;����[5�hˉ�s��g5�ˋ�j�Ӄe:[0F��P��6�&�4�=b�4=]�Q�/�:�2���K'�����y^xY�˪�`m�Yܢ1T�m�P��9�RĲ�������w~�!g4��N;	G��a�>́��7��Eم �l�ʸ��t��/OU���̠J̽=�VmEum|�������K��y�I���B�4J�Ou��OB�\�fgd��g�������-�i/ת;���d�}u�
����x��]�i����,�q6g�1#f�d��p�'����(+���wn-E��fLfLЇ�ȶ��]��2���C��H.V:.ܻ·@l��6dD�*��.� t�֑PE���lΘ���橼ɰ��$�#��43MiOf��"����}ߧ���{R���x{��+��A@Q�~_���R����	����9�f"A"��!!AIBD��!$H|`T$*�H�0��9�x��b" !$ I �(.ia �	� �M��pN
���� 9�<�@a0 �o3�� !%@H@i(�@ (� &� �fPbQ ���   "A ��d�Da��idPh%@	���D(�  "$`�P ���� !�� &��UX
$@Ii`@I@i` h$@H@ �� &�@@ ��@ ��P �� !  a- IV�%�@! AITC�y��� Ǘ��E �A(D�?��o���������
�����>������g�� O���ִ}�	~�������`EE�?����� �����
*+�?���@�i�K����r� ����� ��y��� 7�~��>�?�?�O������?u�ߣ�PXThA%HUT�V� "@ �U`�  � "V` a $Ud! %Ud$U`eUe� %�U�$ 	 �U�! IYY�$�.Y  � $`Ue$ 	UYH@ aUa� "P �@ � aUh$ � "P "  �@�T�W�!�����I�h(
-�@�+J��>�����??�(=�/�:�?���o��*+���~����?/�	�����P?�������?�TW�~�$�O?T��QQ_���?F���Ew�?x���QQ_ ������C��80�7�='�xz����:PQQ[�C��?���(���	@y�<������;������I���?�|EE|�C������z��:���~�����?�����{� }'��I���AEE}'�P�|�2��|A�����?i�� PDW��`�>�����/��O���d?z�b��L��(���� � ���fO� ď7�w�J�+�UU)J�"�m�����D�)T�H*��cm[2������"�"k%l҅(J�TM�R@	PD"�@�RD#݇�$
$��).�P�L��j�(@�UUR@*)QIUH��!(*��DT��T�+}�!R(H�!B��R���E�J�U)*�����TQ��UQTT
ٖ�)�
�E��!	%$��@]�*�Qx   -U�g�wR�P(]��Ι:�ZC-�[\ҭ���mu�
U�b�)�J���k54զT��C@mm��(�v����(�D��QI�   v$v�	
(P�
{bD�)T$;^N
(P�B�u:(^�y^ٕaAlf�,Y��m�/l:���`]�S�eb�hh;�fـ%��Z�$��T�:h�m�  �U�A�������$�i���;s��h�N�v��[TmSm��T�cj0ƚ���j�VI�4����4��R��
�%(��   a�ZkZ=:�T� L�K$�i�wmf�m��Ҩ����l�.� �n�WU`ʨ�a��TmL-����#R���B +����6�B(��  �������2����5Y@�0TU�����ka2B��XP*�iX�X�$�h��UR(P�����t��  �$(�iR���j��JP-� m��ATB��R @"��!V�U(	��j����:*��URt�T��J@m�[�  s� -ƅ(ZV �L Aa�j�Z+U%BV%�THŀ  �� �X  {��h S&�0IE��  ޼  ���@F  4j�  40  # U @�  �i`���` (�  ��T@�D��H�G�  �  ;
 P�  
m�  ��8  	�a@ 3  b` �� kjj  �*$J��(R"$��   ׃@ ��  5� m��@ � iXP jX  
��@0� �f�6�@ �S�)JR �Oh�JJT� h �O�j�P4 E?�$1 �ڍ*���� �)PLU)� �bl�o��M�lL��d�MT%�L$+*�-����G/v�mC������_��G��o}�o����6ްll���1��~��1��C`���lm������b�?������f'�;v�H1{�a,Z𧕷�lh�┡t�8�9 �N�%E�����P�u�$�j�ti�`���i n<��V�'�z�&5u���3�'�c��'�Z�W�+BV��s���pe���s&��!�$��<��`$���Q6�hn`n)lm�p'yD�vd�f���<Tv��,$�Wf�Z�6�Tܼh�V�v���0��' Á�k�=�FŤfX�w�b��m�m�'H����f�Hʸ��P����F����� ��`
��AVC`T��ښ�<��ޚn�q���ۤ/{4a@����m��i����k��p���F��\+\2�W[�Q9�NK�V�1�لEM��Z�zᘭ3W�`u���M+7N�**��0�+�/V�[LmS�F�c����XzuB��Q�YKR�-u1����(ҪplKi�Y6��%�x��`���-���`ŧTO(�v�JnDq��	���T@�Bi�X�w5���<w�`R�'��Si$�k"Z����"7��`�YqU�b�jP`q`ł&1��no��3]�AGv��@�ծ�P;[Aj4��xg�cR��*2�`:�u�Ʋ9,ɵ�"�J������A� ԂRZ��s\��������N&omHn^ʉ}iV���� X1�Z������`��J�U�cd�6��̡��"��/EڶM�m@��e[�J��#�7���,��q�rR���k V4[��#1VY����׶q�Ь)6�f�K\�5�f��P^I]���(8��s@3-)Xb������ ����!�4mWV� �X�������7؋إ��>X�Xi�V�V�܈��M*�h�Բ��Vj
�Ry��4��:o)�!,'�7jP���N�˫z�!�0劙�)Y��1]�]�N��Cv�э��%h��]�Vn�2��;�vm�@�������	j^%R]�l(�[JH�Mե�xdX;��xY0ŗ0�H8��`��� ��mQ�d����J�������$z�
�p�J:6=�R�Ɇ���(�E�y�NR�:��V�so0�c�Lrԙ>�{�XV��84E���Ԣvm �	*�a�8�pR�չ
��e�X��ܰ,��(�+A߱��2���ZN�ض��(�s�1�Ҍ:Ʈ�a�լ��)��-rT�;����a��Z�z�C��1X��s�1=�
u���O*�c�ޫ�q����+Kz��s �೨�+wb�z��R�I+�w�SRW��ܺ,�X�D�4�S0L�^�i����	Y�V�V�@�xkP�!�hC+r��툫~�!֢���0j��H�$�r��r�Q��#:�+pkW�z���%��m��nI��w1� V�u�l)���@jQyf��e#+FH^ـ�<��d��VI�QyM�,�B䵗��m+.\�E+��a�7\C�A��{�Ŋ�tI�k�,|�Z6\)H�y@��ؼn���H���^:�v[��f�d��!�V�m&�5�)j�BW+G��n䫐�:E�R�]]f
.���l��Fݧ.`ң��ke��X�s"�-K6V!4Xe=V+�D����Z�lQp��(�w��҅T��!F�m��(d�Ӄ.��e�u�S8c�p���wqT���T6���m"&�F���k�r�)�vb�%�i]�A6�襁�4vV<�,��e�U?�6
imw��d����F���)B�ܛ�J��H��cY��4ו�ZU�k�b�1eێ�A&2�fA�Nƌlb�,���	jS�`���n�l���om˦����F*ݢy�������i�ɢ�[���:�*L�ZWq�e��x
J���S�R��� �Cj��y�l&����2"R��p&[����E0j-O"B�,ŘY�:�ɛQ�(յ���?��Q�3r؁eE��׌[�*˻��G4b��m�m7 ͳ���%����`?���)kin]��]iq����b��� �LV�t��y�d��Z�ca�#�R��՚����ȟ.��~�]j8kcjӑ�&,�Mx,vm���
��J���'l��KB	a@��gs3"Y����-��l��T�V~�14�0m]Y1M�8m� �/6�E�����S�����c�ط%n�eW���5��CR�(��^�PaRAҼ3$�6���a�E����Q�s�Xenh*�!�i��G2hA6�J6㌂v�d�T۫��.�lT4M�Иu�1��^L�ea��� R�^�SWEkx��!D5GT)LP��4�!���4]V×��/ 4m�j�7��c6���������/N�4F!�3l�P��]Ϣ��ՀQ���
k�&m-�p�b�{{��j�	����ٯ��hf"� �nе^�����&YkZ���5���;Z�*r��MLAT�J���b!ܻlA��YMTË6˦e�v�X�d�A�5l�0dFc�D�ʲ�Ӭ#���D��pӵGK^Y�4�P=WF��,f���H)h)k-��/-�N�f	�"����T��֊D?��,���:C�1�{.��jXL���T�l�)#��Uko*^:�,�]k7�ȝԢZ��[�TMc���&��)v\kXKquZ4���c
�i�{�7���8	�b;{b�۹	!�X��?򦉹�Yq��Ĝ�s��ehٹ�d��jٖ��+�VVژ�5�h���`�2�x����w+\���U�eK�c�H�U�Q��O2��-w��X
���� [h�4��[4��mR���� Q�ę!̕�7z3lr�<��pV�ײ�K�"f����c
�k6�lfnF����mZ�8I۸Uhjm+O�H�˶����۹*l�l���%i����.WB���Y�a���Շq��,fkX[�� 7+�{�ZR�hY�M�h�T*�JRm5�[�%�ٙ�i�dL�a91�x&�@�ac#	�J� /�c�S���1�ۧh�:�`T��Ӕ�+�f�����Ot�I}L������"^��flL��.�#yՁ����/Ĭ�ͺP+�Z3q�*az�齻eX�݂�A3B�Bk2���YRK�k�p����X|T���*��h����cA��i�X��6 ��u4�%��iT؂�.j`2*��YSpJ6����^�k&�A�ÁA��l�wpd�"��n)��k�,�ېg:Ѵ�oX��,�Q�3p!j�v��(@�Ŭ
�m���E){6�=)X�����CQ�A�ş��Yg,��t��mC���15aDk֊��Z�b%V렳<�<
U��i�Ȯ�I1D`Y6�Қ��n�y�;�N�R�]�zfVS)b�YvJc��V�T艒 �����5�e�
E��GJ�Vى\�S3�D*Ќ��%`2�]��p�m��T�EB��Ť����m#�f5�Rd#n��Į�M�,� F��<��[h��u-7��,qãS��aJ��^]�,*[�����Rm�o�a�".h<k4(T�B��JG���%��q%j^'p5al5�Z%g*�R]Ae��Tp�նD"|p;SX(=�Cc�g,"6.��d� �o�R��);�I�����K��&�ˢc*�7,�hb�e�DϮ�#w�i=��*:�s�٫�N�!b�)�J�l�*��(%%R�^V�[
B�`fS��CՒ�9�,�u&H�J�71m�A�@�C��f�oq��`ڵ� �7qlܨ@��h�շ�X�=Û����x�H{V�����^�pU�p�7X4Ÿ��і��FB.��jԼ4��OY�6�	� 6n�j4����7]L��]�l<t[�/PbHE� �zhS��!��N�1��,R/����3�D��72�wj��kj��iVT�Q�ȝ<iX�� ,����T�o5j�E�ERc�~T�I� ٩*b3X��T,<ddl�dX�U�	Em9tq�����g�%�V㵋ujT��<`�h�zT{�W�y{�r[��Ư���$5��j@�Z2ٔ��S�7^܈�{laY��N����Y��4݅�Q�����'c
+ ���:�}�$7p���Ԣ���t�H!�3Mm�/^��+
�)�Ԥ���퐚vr乇kP��k�U�!DT�Qvl^���)ú$��6]�0�Bӕ�mCn}�,�6�2�v6��	���w�v��5��r��)2��m�+6��9.�ڔ����b�`	�Ӡ E=Vl[�XN�ں`���'w��^�l%i㡗���#n L��W���YC)J�8��������eT��j�నn��*�KQ�{��ڲۧ0�u#��V;�ec�WY��d��ҏ^�4ȅdw����f˚%�h�����>64�m@6g�
�Oq^[��Ɯv�-�5'(�/R@��
�=��mK5�#b�U��l�X�2I;H]�U��x쫨�GkLe,�e� x�V'J��I���f
�Ƈ��sn�@U���d����i3a۠��XrXEj�Ch'i�/�)��J�,K�S1QwL
Mk���-6l�oQ��"�73b
Wc�7��նaxx̩�Y���.�2�:�Qa�e�V��i�i�tO�;�[o!&�"�n��Z��@\��M�5CSQ��x�5�[�B5��f��ڻ�5D��T#2���MsoT�����@<��[�v���Ø�t��+_ma�1WM�^};fA��(�Y��"�t�����;��df�wNS��i���Ȳ^�n��y�X�Ŷr�������.ux��j�B�S���kl�
sn�bʏ4�Hh�iM�)�Ǝ��
zT��5���H�-���뤭M�6�G*F��ֈdUݧv�(.�ܳ*bF�V*��tä��$�t��l&)q�2]�V�˅1&�)���!��jI���yq��ݔZ@7uum�bA��)f�7�9sQڻ�f���WK-R̰�.��Y�܎](*��d[����՜lm[��ڔt,�3.Is��z�_j�H�Z�E��x��7��n7Q�� U3>kZ�]D�F����`�ɹ��!p\c��f�4n�K��lj��O��o�{�P��X����������l��RҶ2h�n��H�6ˠ��[�b^4a����M���,��b�JFK�[TW`J�n�OT��eK�v���\Q��c����Z�2 �4,�G]k�,l����m�Nee@�m��E9��&���[��al���Cr��P�ĥ�,IE��vȩd<�en j�<a�
��Hķ����ht�G����z�+�N���23�.�AZ��`����9��Abī-Ø��a���aso6񈮦壩A.���ɷ2��1m3�&��X�o^�b"6/4�4�k��]�u*�Y�7y��eʏ5��R�%��
x�lņ���2�Bf'`ӽ�HŻ�F�-ׂ�D�q�ײ���7�v��L�ل��UFejV�BGS�ʎ:�]f\Ү8�i����n�14nlX�Fَ��[��J�nt<��[��kA8oT�E5,��j�HJ�^n�O6���Z)��c�N��T�_ي:`Pg(Q�oI�I'Lw1V`-��4��@�gX�v�!b����2�*R���U�ٷSsh�d���-L��58Nз��k�f��+r�2b�����̧�i	Z\jd�֢�4Ǵi�!�F�`
4ᬋS�SJ<Y�ʚ��%m�6!�v��kl$�۱G���h���h@%N���$������P�V���CZ��iZ(�m�6�LN��X�<k���b�Y�E��'E3R��N�lL��q��:�0^tӦΨ���,�!9e�ATܨ����zQM�i�,�[��)����֨��VokZ�����3N���V��T0�3pN�A���۴
���h(f��� �gG̅�F+b�� ��$Uts��vTԐ�q���@��$5Y��� �R��4��qd��f޼�@P��"���w�3�]��=�:�
�1h@+w��+�m,�wiڣh�����sX��X2�g� ��˺'c����q��S_8.���^a�:�>ݪv互�f�w��(L�Wg*��2�FJ)i!�VF���+R{�(mқ�4�O�6|m[���;kJj��8��T �,=7� i����(�e��w��t=U�n��d)�I�k�F�5�k-^��.�K��;�f0aʍ�zm�6)�r��Ȇi���'F�2�H��!R�w ��2�6��j���®���4����c��G�X�nEB�2�Z�h˳��UӔѰ�L�aQ�m⎤է��{3Ei����L�X�!�_e]��A�J��eAv6�#�7/m*�0��F���A"w5�n"�bǻ����r5ge�5�R�u��̳%�~��kn�TÎ!�T؁�)I#�nk��!�,�4ѧJ����j�d�r�L@8h,�.�����oM���ư�Ej�;#E
�6��-5���m�TՂ�A*ܫ�t�E�@����8�X$[`�P൪A�8f�A�{��zrM%2;��ҬM�s��Y��t�ɕ��`���>[��o+\0��kj���uj�i�������2`d��%�Ο�֜�b��0����ČfxTm�	3d�X4`����$$s2=O.�IGu�J�t��&+�I�bYj�]�$��(�I�G�dal�ύ�qE{zJ�:�`,0�vMүk�-��J"Sm\Yt]�aJ�e�QW�xf���);�_t���](�E�㣻�t[:��.ge�As���lU�N�֙�B<�+�8��{��G:w]G6�:qO�H/3[��[ͼߊ�HN�=���6���Fh�s �Z�G��ĭDL���*}�)]���ȓB�[��i����iT|�  ��+�`ǧ�S���so2�:u9�7��+@�s}�H��{����}�+< ܒ�hD�{6<\���ޮ�*�X�W�SivΔ7t�h�1R�,����
�n���z�D��㉭�)��u�����5�u4��ъY����u�y�r�0��"�j�\����ςѶ�{�7�!G;�|w�/3i_D]�u�X�#|�1�'ޣ�M��J�\�/u��zޠ{U��wR�C�}���hT�
$v�yl�+mm�`��m�/�}IxH]�օ�۬�ՄK%5��4����)HT�ј�?���Y��,^n+۽*��8����>c�Η�'G�-:��w-q\kZ����4��7y�t㨾L,��ůgQ������Gqe�S�)�o4z�>C\7���R����1w�{8�i�����V����&qӦ�`o�pV1��̦�з�0���*��Zcg��5E�3�7/����WlQWQ��
n��v�k(�];��w�:�7F�M�S�O�u8�yH�{8V�����`�q`�|����﹃V��L�@�{��WY5���Y>â�
J�n�d��S��6�;)�U��{bY��I����jr�-���=�W�\�vk����ܬU.`�y�ƭߙ�쏩��0ŏf��\a�lη$����9��gJ�leVKXzrj�]A:���n3��
��y��Z�{�dj��w+�ֽ���i�u0b}�s92�'�d�miT�X7K4i&��}vh�Q���"�S#�qC�\}A���[��WhIh�������d%�ݘ�'�wa�d�����Z�Zw�F�1wL��R����s���*��{v��|���)�½����`�CD�vc^���c'0���;,��Vd�G�o�=�܎h�E���V��+���� �Y��ݗ٩�I��-�Ks=����:.u���g!�
�:���s@eqX��C��]��TI�Hg�N"@�sza����C!|���^D���+�4� F�y�3��V��Vm��L�q���{��3rK�͹E��է�7 ����U�L�碘�b��C�&42�d�[�`�P�e��?gf�J�ç�v.��C��Lt�uua�}Q�6��bG������ٷܗػ��37l�����B8�!4g@�9���zuv�!����2pJ"S��Y��ں��/d�b���=��q]�W)ju�����b�o�&'j��C�l�:&�n֣�n�mtIf&b�Ϲ��|齂k���|)�/,"�yq�Օ�T�*�3ֈ��X�Gn�1�Z��n�䯇$\��ŝ��F�D��c��Dz���l����]H��0�՟s~{}��jA��Q5���mr�X��D���:�m��PsG-i���-�q �5��G�M�O��IkݚD:7z��!Y�]9`es��^e!s	§k��)h��E�Vե��M�"�H'֚0%�b�H�҂����F�����ɩ�I+�����.f�{����$��*Ayɑ�6�ݮ[$:�ȼ9�Xt.ˮ.�I�)\{������1�އɆQw��<��@�Rƃ �b�%տ���<��hwGϖ@�vLY�V+i�n�a����y#��M�=F[To�� m#�ua��@�Y������2--����ѽ9++�F��cC3��$�n�zz�x9���Jb��2��!�s^��������똛�x�)�gY2�i����~f%ə�6�:���M�j���/6v�Fɲh9k���J2Xܘs�Y�9)Y�4�vz3��uK؍�F�]Ynq�[�\�#�n��ү2=[>��;�X��j���Q������u7�dZ���h��I)���^2������`�QB�5gaMh��
��c��V*y-?��Lb;2���nQ��:����r�7Û�q��^�.���%9ܭ\
� �T��w�q�8Ff;V'!�T����r��3^���L�Y�Ko;' k �*���̎�tj����QJ�Y�;�ۦ��޷R��V�����(oM��A�+8֧C |[�G%Y5ӯ�8�>�+��zh�N)0�NfȬ҅��]p�]di0����_F�e�U���A��׵��4�3_f�n���)���>��;b�����+
�r�i��F���P帩Ա�+5;\N,���>�4��H٬����;�%6�ɘ���y����Դ�<{�t��2^2n��p��l,ܛ��h����KNΨX{1�6��
��g.y�h��W��oRb�uy]��wYq���6R:�:�@��P��x�(־�RJ�k:q�a5D��Dm�hs���N��2�P��u�Q�K{�r���\o��γQ�u��w������l�X�ɮ��]�ysS�A�}��:m��q^^,�].K�w_%p�Y�Ȼʱ2��(���ǣ@�M8����B�vO.�י��H/��d���ͅ���B�p�=��F";�n�[Miv��g��u����1�)����6���6U���fK��Eean���ܖ��ĝm&��K�V�٤�kI:�j���:�T��WA�&��� �c�ַ%���Etꄻ#��ʂ���W���V��aG[�|���(��vx������Ϧ�S���!�\��Y���}ًAㅐ�0�T:��Ȑ�]]F�������8�a��Sqn�O��%���Pc���KO���o����"	��z��s)��7��|� /e\ܙ�"�Ecp��N�mXH�E�`�МGgs�j	֫� ����}9	i�-<O��a&��v3NR�ʙ#�}�M�/V&�R\���{;�'��m��z6�\����m�7#v�&��}�������Y[i�1{gj�益�ӧ�a�yw+�۸Ȯ�B����a�ҡF.�e��ˈ�����,��E�	�Y���{�(l���r���*�vD��>���D��9x�Рh9�{��D����r���W�3�$��|��T�ID�>�)�غ����aƩt����Mg/�Mݩ)}�%�8����4��u�n��-8,��,iE�zܢ"�� ���]��٭����ع�T��[�l�W\tcw}ϛ��}�'����~Ky��T&i|q[��
�jn���#�3�a���rq�Ӱ�{�N1�%�Q��]0uYk�tۈ��z��I���B�f�o�0�ڰq��7�|V&�dK�H�f�]��7o����vьZ�E�p�1ÇnP�ݫ��)����|xV�55��p�5�ŕ�����A=�y�e����4�gnGWfѹ.Y=}�t�x�w*��]�S5h��.!Z[G0gn�t�gq����mu[�-�k�w,i�����m�f��W�#���7�P��$�`k��:|0���r��:���߽O�˷�:���/@).M�7o����b_�7V���灲(D��
��Z�;J�,���rWu�&��F=N�����=X��QN�Mvm��m��#�Ȟ���7y+AU�e�k���I��U��rqG���\�m��֛��Nһ�')�w&:s/ �:3�c�"h�2Qf�Otw����U�e����uL}�d��t���є�Y�i�m��ǛJ�������u�b�Y՝]�Z���i���;&�kP:���vA���s8q���[Ѳ�;��/Tg��,O�r���	���'r�̃��w����V���"!Ӗ����#��VZs�uZ]]-�z�ҼA�{�ȴ�U������2z.������TW\I�Y���|��)bU���!����r�-6�{�7��٧�a愂�ǏL��jחn��o���1Ôc���w���֙����
�;�%��7�'nmuŚ�fQC�����d�Y*<o��b��b�aG7��v��i�����жx��� �WV~�^�hwR`�vUG�.����S9F��W]����$�B�U��T=�ފ;��)k�P�f��1�"���MKk0�s�9:o8`���<G��xT��r n���`PgVne�k��XY��� �E�[l	ۜ�;`��e�.��Hق�6��W��D{��<���m
{\�2�8:��@�ܒ��uxepUete���=���^7ofvy˰�t��:��
�WzY�ˆ�R1��)�׉���NS�n��֔|��ֶ.RJ��;\�h�2��(��{쳹�igu)p����L�}�*��Eug.�^�Rf>�EuIٽz�ۺ�Q���{>���G�[�(�b]��$ˏC�A�����Ҵ����)�ͅLeu�st��6b��{P�4�3Fx�+�v�[܄���!�F��"椞�tŎ���C�;���V	�H]w;|zo���ţ�(��
���n�f�ޣ�&�1�5�EB�b2]�K�����ɸŬ���At�w3Օ�R�1�3c��z��\ksC��ڽ<�5�(+d`M.O�E�̭Š�[�*�E⧃%�h����^I�hޤS�VP}�I�P"6�/��[굪��sS�:쭹��ާ�ze��M�s��
��@8���;��]9v������f���8�á�pW75�P������M�egs�_�kt�p^���W]�Z����JtO_p9\�!N�,�o��w�����"e��(:J�f�=]��ʜ7�6�kVh���*|�����N�,N�}l��GzJ ��;C�v�g����T�Y5��۬��D��ۗ�����lf��t�B�:���ŭ!��R�*[af��ՌP����
�B������j�:�)V��y5W\X�(%9�S��R�of�5й�tZ�us�ϭ�O�Gd�gD���D�k}`mpx���FN����#%��:{)Eq�Z�x�u�h�����D���rYHk��4lx�K#~��9v>���ո�NaF0u�/뱄d��Î5u����%�VH���Rt�dhHY{��)�[�)QE&d��hٽpt�]6��N�"�k����7�P�0��A��fT_f��_��R�!�gb����K'�����#q������=h��^F��-���{�Om�-�mI�}�����D�P�{*�Śy��g(0�3s{K�"�54%^}YƳ�m�p�3�bR�www۽���x�}�n�``�"����v��:��[�O���o�y�o:U�����VV�&f�9�!r*Q���9���.�Ґh��Юf%�����^P|I�k�у�	̷*P>��s,�WVh�������͝x�#k�r��J���O��Z�Z�Z[٘3vgY�R<�Eoܷ��7Q2�e��Ժ�=P��\F2�pcUb�i��E�j�\4gGCzF��!�Y�V�5����{BF��`�m
��ba���am��2ú'��3-V����k�!���H/��wy�0���奼����3�5�o�L� �WVݰCFm����sQ����Ŏh03Á�����7�v�U�ƗVc��|��n}%5�U�3���B�x�*�w��[���2��ة�=w�̢��g9��v����T*�м��)𛛋�,��yF��xIt�V�G�=�u��Ti�r}O��v�H����Y���yeP269�Fc��/oe��e��on�]` �o�(�H���/��]K6�i��1W�I�
ƻ�� L�}����-w-���v�`μ�4;��4xT��]�y����k
���1&*�� ��Z�]^殫���݀`�zW%��6t���Bmm��2�<�-L��OMb\4�3Kه�-̇c,�v
u�3�W*�f$x����B��SY����uO[�ƄS�d2yŹ�%c�yV��7/{P��r\����`�]*k�U�G�t{11hޙ�Q�cw���E�N���:��; w|j��[�(u-�򊉦��eh[ڱ��5��rإ�v_v�S����>�/��p˃�9��j�����4�������Oj�\�t=k�@��Ѵ��ghDoR�w�뮋J�}C��ۜ��������r�$\�CWA7gl��\O��0j�4e�=��/�0�C��T��p��\���%s��	�%] >{F�ȝ��W�C+7�D�*�A��f]�\Yt�la�4oQe8e�p\���;Jժ/�EfQ���<z�Pk���M�a�7%5m���]q��A���lP�0�G{�UY��f���rx_{�~��~M�/es��u�gPl��Nc:�����IڅnbvE���(Y��g#z�	�ڎ��{�%-��άt�}��*�}x�!�	Cwz8�u1��J��[�oV��NoVD#j�%�������{�����_,؄;Wے[w:d
��à��o9�T���[�<�oƂ��x'��V�U&���v�Ӣ���Vv�ZXwxpk\yT8�V�CQU�m�Qh����En��N�Z�7�Rv+K���G��C����u�����xP���ވ��Cѥ0�:�EV*�Hs��Y�c�f&��3��jJ������Q}�A�6n��4���W&:��;��J�)s��;Ν�;�T��Y��Ԗ�cL�D[�x�ݏ7�,oIE�Ggh_Gd�38��
]t0����萧�Su�n��ź�)p��Mk�ɤS'p��=Ik>���4��=*h�u����5C��m�mm6k]������`�؅5 ���2� o*�Y��حY�۶۝]���8;���ˬ�����ɳa�Y'n-�s��J���n�s�}3���B���3N��;�	�ۂ���-ON��n^�1ڹט`��)���%�u:�z�9��c�,���J,]�B��F<�;w��PpS��\i�_S��hu��y��[}N�w�
�V����m���lm�k��������ן-5��;H�ZgGV���S7��u�T�J�ݨG:�����9�`:����>�{������Bl�6y+��.�<��3�z��*f��R�2]v�t.t�B�� *�]�݉�Y�ōG{]�N7yY�ݭl��=glU�WOf�S��l������26�f۵�.k1���)N�XUwR�T�2'oJv��7%p��X��YX�p&%��+zW|�,EΎ+����3jt4zn�{y$՝M��l:��L��=���ݱ�nFA�q�������2��U�M^��_�������7Mݿ��B{EwWi���Z�3k�"���A�x�6z�WI�r�c �Q�C���;,�΍g�A���f���Q�&�4���[�`����K��Zu�K�lJū\��N�gu���fR�6������)0����]{$nZ���Kr5�+>�%
��mK��F�X�Y�W#R�yݢ8��X����b���B��&���q��*��mht���zMc{�,��Z�s].pĊ��R]��"�������� �U�^*����i��+�[�l�n]E�J�b*y���C�V�/��h�N{��fj�qrcs8�Tn-6��"o����K�L#���-�|���b�kw�G�n�}��v��>�ջ�]շ���s7�$��W�w�� ��������g�**
���&Ae�7%��ƴ�Jɜ���P�wÊ��h���WMQX΃��+�@I5 ��)�� �6����m������x �o%�����H��XhIWw�F%[]��Τ�xoNn���9᷸�'��\�;L�;^���#R�§B�2��S<;�8�ԨⒸ�&; /a஥�%hì���g0�LT��;�Gl,��O i餶������-�\]�h��Q�#t���gW*x��hE��i|4d7��Q7�އ��������1�9y��uB�k.�lR�r��O*�Z�5ܛ���nvm�}(!i�u�4�������f	���[_#��	���pؠ���7%E�mI�ݡv�`�*˵�׶� ��en�0oz�&�mZ���+!l�Lc�<W�+ް�́v`�h�x�<���wCC�Z����m�u��mYީ%�r�"N�]�nwr�(��D|����1������k��9��nu��#Y���W\4��k�h8m*�:�Ҝ����X�䮌�,^le�Ɨ�Kw�1ٝDh�A�{�1�x
��^PI�M�y�F���aT�E�8�\�k�8Q3N�;k]��`�Ow�����ծE��mu+W.�YNTtE�eӓ���R)-@�F��:�^���{�N �����x3>+:��3ko��v������Y��-3��s��]�&�;NU>�rm�Cf�*�P���7Ʀ�& m�yP2.�K����\L���̿�	�h�H���-uϻuɃ�v/)v[ǯ'�;���D��{z�s�6Ex�8���b]��|�9)3��uP�R��oSwX�_<�D�\�̶�y;��9v�Uc��;�q�zw]�.�4u�9�h�j�(d��	]+��'ba��hZx��ƃ��t,��.��u*�f]ţ�5]�O_;iΛP�N
�4>7�:�
�L<n�qfޔ�>����v�S�tbS�9�A��{G�Ҭ�X����rL�hڂ�*C�@����cr�$�{�WB��	�rW
�w"�3xN���N�+3��]��[�Jf�Uq��]�}Cx��CJ�jW��6�ڑ�h�o�C����uq�����X��ibY�v�(�Ջnh�2��9�8��� ���Ť�k��\X숖 �$�/{���>h}7�*\Oquj�da��B^�Bb�"�1�����T-�;/!���q6)ڕ��+�6��`-�e��hr!�au\����2�.ꛗ���{y�^ˮp��C�
��R�b� =}��Y�'��.+6�I�*���Q'[`:3'u6f� ʀ�r����X�;�C�1ȩW�\�rl��,dzN���]e�w��M͋:�vK�J�ɼ�[OiA����
R�:�C��mm$�q��)��h��g�V򩄦�(�].Ѝ�M���̫�{�6�p���(�W�<��h��ϴ+�,�c.�:�m֙��b���J�#�pr��v(FoM��К*�䗛uԁ���My�dZܽ�
���Q�[:u��3s�D�B�ǽ��pR�̚��uv�s�t�.�n)�a_S���@��*/m�/c�8mN�p6B[��v7v-s ]4�!BZ�8����:�Cloeݮ̓�#�ׁ�q*��s6,���.A�A}���2'�]�i�|��x4�,	�'t͜�Ԯ���yZ��K_]���Bj���HY��uѮ���[(̭��C��3cR�
F�+��w:�Vҗ7VZ���˃4�\뺻_W�.H60�g�%n�����脧�n�'V�\�r���v��)��s(b)�(^z��)�zf��z�������3e���+��j����
��K��c���:��&�p�*(婭BK��o�aah�z�X����4E+�f�9�<�^���I���,+�m��8���#R��q� ]��w��(¹
좣�7zt���o-�mc��ᒬ[�&M��_2�"�H��K]�\�4��m����x�t�ϖ�+�V-Ɋ�j���_w]n>�UevW`[Hf*5ӛβ^��Z��wJ/5�}6�"%띊�E��wQ�C��!fgf����r��k>�\;4����Z<!A���:�r[�����϶�h��ں��a!����vշ�f�]/�}���.�<�S��/��.�pЬn�N�[�i�ʹW@���Qa��>�%M��n򹗨��^�q��$=]p0:�v�s;�=z���v��oY�{"��>3�fh}�����������ǫ�0V+�W@���4]Kݱ��+���sz�q��r-��G(�9�}�b�o��C�^U��x2�0Won��Y��]���/�F�YJL蜬��Iwf���R���gD6Z*'Ig.�BZ��!%[ �h��xJ6P���q]M�wu�dp��jP5��%��R���;��d�_I��ؑ>���œ8U�P�Wx���^��;[w�ۭ�T�ӷ��i���ܭ|��(���W��N��GȾ���4U�g!�Q_!�shO5=1�=��5ne>�f����U�R�Mp�w>k�dn:w�r������e& �ƪ�"m�O��#[-�l��&�DHu�dm3�

��>j�U��UY��<��!Ԙ�e��o�Yp�A���޼�i�a� b�E^,仵���Rζ�<�Gx!�gl�S���ի,�ݵ��uXR�w�!���}m���K����դ��)fQ�WRa�R=��h������}��$�k�����m�;�R���}��93z�$ooc���m�w��,�"����F�*���칽5H�i]��Z��M�&�xT(L!�z#�f��fۮ�B�Ar�%���eѹ:ke���sZ����#�3���eiWS�)����.[�/p��j��}q�#�I��-c���S��R�ǀ��b�\^�츸�ԝ^����hS4�wC6r������4�'b��l����
I��U���5���(2�w]�j�;���]�]@ $�K�{dr�$%��H�+tm?�hݫ���N �z�]��(��LPͽE���fdQ��ڣ'RK���Z[AM��w�,$��-����h��t5�����L�Yor�9m#���*Q����ܳ�veY�����Me�}\�2^8���ɚ'��$�Oi�qR�˶j�.��;�K�za�^��ͷ[w���c����5���*˝wV]N�%����b����Jg����[ޚ��)+y�z���]J)묦Tbf�3:��� 3�5H+������܊�Y��Y���o�&Mj�V��%']fw=�Ճ��D[L�)V�+M�s{�[;�[ݻ�]@�;�`���5�L�\�����h��ʃ��S"ʒe����e:�b�j�۾�Z4�wK9^_0�.gdp�����{l�X�W,g�b��e3�;��5��-���d����-Ou�d]������lF��7�_K�DԶa�R|�S�����s�]ƻ�"�f��dg!]n��b���Rc:����6�okf㷉R�+����\���L��;����;���&�mi/�U&.���η�u��d��A0��^��W�z�hZh��&m[EϏ��wD���9i��//@��Y��c���굦(Ë�9�yd�q�3Emw^�=�Ws�͌ю�[���[�!"�6ë�ʸ�Ǝ1,���E��P�ͬ�[/��#��br��̎>���d��=�ܵ��f�jJ�Y���7I=����zM>]@o�%l��d*�\D�TWtdB�a��U���Y�����kX��uC|�5�.]{ӵ�<n�uy�9p������U�{�L	z��E�!V,�{���M�X��ڝ��R���ȼ���׶m��n��`�h��8��i�\#+'Wl���NB�1r�8���ˣ����s�Õ�v޹r�"����3�uX��s����5�*���Wa�f�t��h`�vr#-�n����_4�W�U:��ݎ���2��bt��<���b�Z��'�o�TK��W�>��k� Z�T��1E+����!΃���y\����,*o�s�.bZ�{����ݫ\�_PC.@�W�x�W@:a\�V\l����X���Q�\��N*u�0�R6ۘ7Y�=A�w�aՂ��șK7��0u��	�J�N`wJ�k*�S��ې��P޾�j�<�[�o:��pL����L�]�S��@�`�X�ms���]c��pV�WYtEtr�jT����)�p�1��Q��`*�FUa<Ħ>x;z�3���:�pf�;(�n)���]�����vI����'�A�WK����AXH�٨���%�i��j��*��͗&�ZF��r��ޛ�j]5A�Xo�p�y�v&�����6���Ү&[�w���*H��V�^ mw>����6�µ�#�L>TX�k���[KT`+��o�JK��i��劐=�i�@)t �Y2�7N辦�O�+o�;�W*�3T��ve>�1+Y+h�:FaC�[ٻG��p|z�FS�諥v.�]:�y�]�AʖqGM�B�L���t�uۅ�]J���MM�߻��z���n�W,r�z���&T�J}��GpU��jCܳ%�خ�p��77�*Z��*��XlԌS��1m�A����^nfi����֫=g���%C�^��u��͉۩����h.o��q��C9� _>����wb�Ql�M�$2����ދU��a�G�b*:�'���^������[S����|�|k�y[Au�
��4s�`�2�C����I{B��;5  �ʳ�T][ �Jt���Z�S�ܳR{Fh�x�zP"S�y����'V�Pz�IH�n�u㮨	�	*�/9�K
���w�CW*�>©�����R�u�o�q�ͪ��H;:J��6�v���GT�(�,���L�s�/�Bʳwk�%�2cud�)�q����ھ�Bh�1܅�E@���y�i��(��/-*\\DR�g]�^�խg{l_'�PiB�luk'gE�h��X�P
���h�:8*4zAӶ�sgn{6'��
8(m���e�[�2���Z�C0M�҄oV��
̕�s�N�fe:c�+����gw�:�|�6%�ɘ��.�iuM�w���ؑ"K6���ˠ�I O�z�i��18���w�z,�-f`U�ՃKPB�R��=�ͫ����Ff_\r�z��Z=������jm�_O�z�1D�x�9�Z������m���A+ڃ���J��G��-K�_|��A*�]�f���N0�w��}M�̓�r�T���N��t�"�2M���f^雄���ڼ�8�I�ő�t��1[q�����o+X����颬
8%�v��"�2�ٖ���r7W�/Y�z��B��5z�R��S���5�D*�&�� լ�*h�_n_R�w;:wK�;����{�'�8��	�F�����4-�ut��U��������F�.�[p��ٺov�fgɕ|�N]��j] Y�sB�L��-捙D�~;$������!��kSJgt;T������":lқ�xQj�Ո��������S����+����V �
��|T�C2>����{��Q��ͺ2T��� ��LE�8�)�һ�H���SmË��o(��F�[��g��q<�G->�˦ẑ��f��Ε]�mN�h�eoR��];��Dh��ǈ���M�WH]�Z%Y�S,:]Mem�[���	�U���6��+�����u�8LRӘu�\k���fv��f��5&�oD�:���k�k+�ȉA�@���6~�W�w.gEsv�^�R(s� ���TI,�Z�fT��_t꓊`	�6�Bd�{(P��H6�,:�p���p�z�M����IAԂ�\�`u��V�u��$kD#ee������Rް�l�Ф���ۡ�j��k�F��M�WZ* �ǚt7�0��|e�z�6�Sl�3�+C�4F��c��˥�:ɖ��,��H��l�Ў���t�ʠ��[v-#��z��7�[t�9�-hN��Wmq^˜��h*��	r^���]b��$�ܼ=���m�X�ԣl��VG_κ���[V��Er硃�XB�QV�q�ٵ}����[ܱ/�r�	r�%�����Э�԰����z�L�S��V��c�FC�b����Ѻ3)3��G�-&oZ����ƪ�_:�f��^+�k�L6�¥b����
��SQ.ݾ{v��r3Q�g��Us�[l�v]ٓr���r�]n_?��G��G���[:A���]�2�b�&��A�a��5�m��w��pc��ul�(Q՝t���i]<t�4�w�AFUK��8+V������<՚���)������.���1��yU�J��U14�����6��cl�49=�Wɤ�1uE���3#������J��ș����L'����L�y�k������&M*�o��e�'���t�{4P��*(_,�&�����T�X�R��(����{��vʹ�ev�D��)�c.�Z��f�r��q7է�1��7����a�nn�C]!X�l��iG�T�����n�}�ʥgA|���h:N��P�]�rWN�\��l�)f����v]
���u���f�4��k[�ֺ�:�Iyhۅ�L��v��o!>�j������pirQ��M���s��v"�{��^G�b2N޺�k����N�v���L����C\�0�g�0N��R��q|;'Y]����,��	�E\u0�rf��܏;���p�׀���X�5K���Qr��۰h+߸rẟL�m�b}3E6{�t�(u\�n����I���^����ے�A�v�[Jn����&aLH�z�+�1��e�f�n��D��o���Kt�39_e2�=v�P���2k�S��]�ێ��P����L1����{y����/d�������9����s3.�q�I ��+sF��u��`���>!eB�Z=��*0�;�AE�]+���2� �D���,�R��	��! ��"��!3����E��I��Z%r΅(ШuS΅�L�QATF�t�^X��y�q�;V�s��ҺU)f\�"UС̢��#������az�^�;er(�
�� �*�TU�2s����AЬ����,UEhE�"�08�,":a��XW%"C�4����Pj��=��EE����!Cws��=�1�\NidL�y
�㻁�ܬ�r8��\�W��YMr�Z�uT�I!��u���$9fE��r���UI�$a�\$��
(������wJ�X�$�����<���R�ԉ�rJ��s�1s��99�2#��s�:s�r*͜�և+�3ʈ�9�(ֱ�Ze��̮��R�Q%0��Ȋ�0��ńVe��y	�G=H�W't.��P�Q�P�G�)�R���l���<�6�f@���l��en�c��VP����w�=�%�}��l��l��<y�04����rU��UCq��K�mAHV_��.�0訷�,��R�ҝ{[\��j�커�i�|�'��B�+��5=S�Y�̲.� I�3Y_p���F���"��3>�U��*k��{���w���y�q^�f�qS3�
�&Z�Oh(F����8��:��
T�X<�L⏕-t$�{��\\f�����X�pV��"��5���{M:6�zQ����l�7���Lwd[	1ϩ�\(E��e��@L}��jr�Dt5'MCܫ7�t��@Oi�1�/��+Q�R�skJ�څthqs��l�F9}{H
�<)9!S�B��l�~s~w����nU�+Os��:/C޾�VT�mh���g�k��o���>\���^�y���|f^��~�y�/1C��]�PS(pp�E}Qrx�(Y�أ��+��F3���H�F/;|q��iGH��W����S:�w�q���8^��<0敖��a(�s5Y�;�2�fZ��z����Yp��{�W�V���Vs��gրZ_�泮���;(�7ؼ�y5�:����"�R�U=.��U/���bo�m�u����6�dN�;��ڥ�9]��|����m򆙱t��_]�(�ԥݽG����*ϧuk[<5���z7��\�ڥɩÙ�aKXyq;OE�G<��vj
�Y� X�*|��v�66�^UH�|�}<Z69��i�n_�F����\��
%Q��󍋣�vC!���+6��D8&0q5���w>]DD�u���M_׮'��|X%�j�j�b�?,ʴ�/i�{��[������]WQ�)�ÐLpwknT,��"�[����@�� 1���L9mE��k�­h[2��B�������2.
�x@H�r5��Wn�&p^T��¬���.���i��wv��tD"T����8ED(1��;�0��ȀB��_eb�[��.���V���{ʣ��מq�9J 5�ހ?����]�⏅:��G:�[g�H����г���,�:��U�����aT%L���s��j��;(�MK%i"8f��B�:�_�����He�twKWWZ/֬j.�xY1?v��Y,\!LW�ڡ&+�m��d�"�|��h1�y�#s���Tn�ʒ�����<;�A�ܸ@
�ޖD�),����#�2j���{Ui������y�^|dK��X�ʿmy�_���Uep�{zcV�E���Q�ax6^ ���.�6I]IL�.X�M���NRU�5�|��G�Q[B����T��Fe�����XΥ=qvU:x0f�(,0�k�&9<�M�ќ�fӒM�T���3j1���R�ukbX���f��<��H1�VE'u����VN:����Ϲp���ѫ�Ы��E:�e��<%W�~��V�,����9<���/=�SK�k�z��Y���ي�����Y=!�TxF���u�W�f���;�DE�<`"�GG�D�����*U�59�3F��cΛ7�d��z��_����d���m��^���E���@���a�uܥx���*������R���1ImOq=QA\q�l���K��Ƨ�i�̏�]K��)��/�FkI;�9|���T�+�0�vUG..�,a�c�\a������j)��7u�7�0�2Fs���)Wq��[����Wۏ�@s��36�S.�Rp)־��)ˣ� ��/�x�t��F+�s��H�5����\6̙����oJ���f���VnE��/N
�v�E�U+�n`���G����W�(R� Myh��ފe�j��\a\�*�u�7�1�8S�C
ȇt@�T��C*bc�}uĘCg{��2�xgQ\��9f3eD$�s*�p'3q.b:���5ji��r$���AKR�F�Fۼ��jiޤ��v/E��d���Q���"���o��J�~��/{4�x��/)�Ze��&k�c�E�r�nk��}<P��G�Wk�L��Ej�{�_
�:�w[R�ܒ93c��Pn%`g����.T�Բ8��9(��<�&)������#"��.w��9t%M���.��.�jʬ���[+��o��O/pB�e�ՇjIo0��"��
�}��ށ�O��\Cj�|*f�����ڮTs��sG�� ,@���*	cr�3c���څy���1���f�̶&�he�9J:{q���=P����뒞�0��kD�:̤i������=�7u��_c��Oe�Ĭ�Q++.G9�E�7'�����6r8�c1��')���\�I|��⚭P9ڽ�<-�F��ΦdB�b3�0u��l�׷�**���mAv��!�p&�fh��e�v�W� d���ɍ���s�������3�s�n�.*�28UK	��l�=�Ωg`[u��*�/��:�_J��eQ�,U�kKF8[�tÔˌ�n�7����C�K��O�Ij�_A�u�+$r*�[w	����p5�����9yrb�]W=O)vD��[�?�9���Ed��V�Hp�xV�;ǧܩ����^��'��Z򔵩Ժ�3�U�]@h��j;YjP���f2Q8���`��<��P���ue�FN��Ѿ˵�/�`�k{3٦C�����O�ƹ_Àҟ00�o�{6�/7�%Ȟ;��� 9��b��������畜��v�)�w��n*Gp��5ݥwS�Խs����~aq�(D��ldt�V!0v@޿��
*P��bv�yU:��@np�0�ӣ��u'iϹ¤�F��M9B.J⾃��򵲄����9�V(��/�ܖOq�#�1]��OU}!��C{\T湀5�e�DҔLv���u1��T���ug>����<�&\�1�t<7���\oM �5����M�
������	�j�^�ݷ���D,����D����]OK��񙆘��0�o&+E�}V�7Y��99��v��mm�8X��O�_ZtD
�m����������gr���z�U�;��s��n��2�O5Y�pԀ�g�m���IU�^'r��X8k���Tqxc������D�Ξ�ι�Z�gF�w6�
1OTT�on���p����4ͮ��y�vd7�k}��y�zoج1N���V<���W�S�r8Cd��Κq	�0���Ʀ㮮�ލ�;���{������(XVj1��e��'$Z{H@jpf���D_Z�c�b�
:
��:+ΥE�P�X�4OY���f��ȕ����4��&W���E4&�t��Ox	����L�n�6q�֫ۊ9/��Nw��]���'�M��M��Ij��n�Zq��.Y���w���O$	�^�n�<H'/e��7���-&_<���6�A�	zo�/Y_X��9�;P�|f���k��x6a}Oض���cǯ��̔�>�dF🦸O%�;9j������k�[���E�)�I��Ƴ,���8��+�������م�؎���
���o�_Mw	F�Y'yL��wn��6�IRȝ.%�x+!KK	��F���ģ7�"��'��<�@M�b���]F��Jo��ܛ84B��	r��-�2�6ܾ6���!��Up#� �ȫ�ͼ�ֆ�@�uR&	��9��������B�|�ϰv��a����0��j��H����N�e(Zo����7�z�:;��n������u�
�wo��Θ��W5w�����j��ab�01��"��3p��шH�z����b]�w��{۲��TGOLWX��U����f'HY����5�u^�B�-F%Å3G��\�����+���7Zz�K�ü�w4z�h������.q$��;�o,f �Uv�-p��Du��^J{<��A���8H�F�����&`��Gk%"Of&�N��A�̅]+z�K��<e�]2�j��X��mr?W�vz�7�%���:��\��6����1ӗ���ԽF�V�3ӵ�8�S�#��WV�Ђ�����N�Ƿ�O�/(�R�^�UѾ
�9�a���z�b����L����CmP�ʄ����n~|nWV@y�a7�V�Lh�ٺ����(G�V�x��f�'�	 ��Ki_m�x+��&;e�h�:��R$����¹ �s��㛜_k �\�gnu��ٮ���^y`)�\ U[��<.���FyP�{����"����λ�U��j����ƺ�3�0���ߴ��9;��i߯������Ҝ&s�m���<��C~����ݗj�V��|V,�Kԟ,�4�R�ڇu0^9BL[u}Δ���<޶M��	=�;���֟�����H��b�$�u5�tX9�{c:�)���f�f+㪾�����6��+����j�_ϳD��H���̶]�h���n�qs8Y9�{�ۮ"z�������M����2����G��������o�\�+���Y���C�v��siǙ��A�=,`�z%����ɢpVY_KƗs׻ܰu��,Lq�d)��&#]D���*�n0�+r"t}�U��y}��R�WA:x�чT4l(j��K/G�]�9|wXu��C�k½]��^��߇<}�fcB�ay*]!#��E�΋N'��*o�38�������f[��9K�CNK��^J�4�q�Fmea����s�ܢ5Θ�7݉���%�\\��p�t{�G ���Г��FQ��@�8s��=`���WCC���(�L:�lu�>�KV?���< ��ꞥbsևy*#h�k�Txs��Ty{M �a��糣дv����^�$o�z��Y�)�.cDh�{�Y�~�D�3�hƩV�*��o{5��/�.s4%�Nc�*V�^�\���0��[��S7�GKwpj��p���z+�J���5���Y�b{�$wإ���Hm����sL��59b�r�X��D�_svw���x佧%R��e[�?9刼�¼�m1��X�.��"��\�\�{-�H�@��r�`�x#��Q<2�Po����'�a�+�5mw���no�FW���H����i�L�z=��k��p}a{���Cm�2��U��%��H�u�A��[�c����h���䧆)�9��]C`ޞ%2��O���s�n8�cD8eD�!�n*x�o/j���؛vlM��5��gJ�5\1�ɴtn���K�i��V�v���V�Չ�B�[�C)VV(0�wր9g���,�5v�aQ{Z
#��}x���\��
b�[�c�T���	��yY�Ğ��2�R�����]�s��T��uu[�]��IY����c�4�u�y��W#/��z��Ԫ�UQ;:%�^����s���i���$P�=��m�]>���l	�v�������@kX�*���M��V���f�V�NӚ�B�N��8�������	��ϬJ�Xz6�����GùD��K<��m��X�w�������a]��K��欓t[}R�v�cB��A�!l)z�3�k����0�e�E�Fa��5�8b�D����z�c�Y��0�6t|����(E9�lVuPE\!0r@޸�v�z�vgn6���>�!IG.���qϨ�g���I�F9g���!��%0W4U�q���lw�5=�I�.	�+AS]����MC��x\7��Nk���FM��������0e��9������G���GC���p(>���X�SC�����C��/y� �n��e�J�2auS�R��k�f�̕��
{����c�%��}�t��3C�ͻ�hz�����BN�"���W�1�-����"�.���"�-@�݂2vAM��q�~�Cs���ɀ-W�{�z�|uu2��띳��8��s�]R8�8=��a���A��E�N���� u��I�!\`��fܮ5z��\}���Ӂ�o�ji���T�J&5Qܤþ\�j�� �c��[֭񸀺=�����^������j@h��o�6B�\N�<*�|��o�����'�bTeԾ��q��X4��},;O3>�j`�TL�o*����8o� �RWFޡ`����gr69��;Qs��b,ߧ{��1��mƊ�tk�Za:��5��3��13�������ΐUa�ʄ*�iB09qP��6
NH��m1���ѳ��f��piJƕ���"��7`v�\Ϸ�U楖���X���+�ڕ���H�E����v�^����S�!җ�ע��I�W����s�Y�)�.'�t���"�Ij�Ew7ӟ����*��q�[�a���Zj9�.�z6�"xh9>o�S=+�>6L��$��i����aU���f'��} �����e#�Cɍ���U@G�$	�Q; C1m��x���*���[�S˺�'/���A�YU!�X���g�� ^ck���k�Ժz�ymZ~�0%8�w�����\��UH���CI�y�����n�Pi��Ӂ ,D}��V��w�B�	x�G�B7�_Q�=
%��S泩_3�n3��s�q|l�듩�؞�jR1ݣ-$;�J��V���&W'�I1gr	)�������Y���wV��F�;C�%"�:+�kp,7BNU�o4���J��艬S�>��T/��&��W�;��g��i� 5[�ѻ�k��r4�WZ��ئ�ӊٺk��p�@MYx4�\mҨ�V|��Ty�V�%�>̬�X�˫|�r�Jܑ����a��7�b�˭֝��w�	ݦc�|��q��;�;rX�Ԡ/x����ts��/����
��q� ��b���	�+m�U��̰#Tz�Sc�	���M%ژk}k��[�0Q�$��Rz��7��Y5��R���2�ywt���[��@�)�\n���\���L�u*��9a蒐J��oj�]-��;.��6�5�;��XE_=���e��c�w(q�m���k�sܑ�x�%�-9w��1�O,6�b���|�e��u�(���еI��ղ��;Ps۰����	�M���K�)�׃��������&��%-Dp����:�z�ҭ&[ɩ���"�䱊�f��-�iB�7�Ii^�[�mc=CO��p��rVėX��S�^�5�+TF��n�39T6q�]˹^Ҹ7Fa�49�Eب�L��|��x���V�b;�^Ro\[�#���W��U|�u�u;QPu�3��超qmd��t���&<��/-h�#��HerZ��,}��w�e��?$��0o�nqy%:�ݽ޷}wTa�`�<:l���$k ��ùI]������Ng|��)&����ǫE]p���[�hf�{�Y����lXiu.G%��b��o��`���'��]��7�de���$����ڱ�V7�쬛�K\����F~��Z��8�\) (��K�1Y�i��N�.��,
�e7��A =]�>�Ś��x���f	�\���GQ�f�\ʆ�zMa�zv��	�oL{��	�S�J���8k��o
Š��-�>�\L::k��9V*���X��*�4qk�Z̹S&tqr�u>����$i#��%c���H�x�p�W�gS�
cu�v��Qq���E���#Z��:F�u�%�n�����#u��[��}�
3M�a�m�};���[�SQ�8����[���� R�ep����(��MV�G8N��]�5����a}ո@���e�}$�B�2+/H���ig���m2�t-�j�,��%��f�ɛ�q⌜�ޞ]>_:˨�J6���i ����QgLx��GX�y�G���b��^�5L��n,s�ճI�:w��՟j��P�F�F�]\bɄoN}.��V>5�.�^m�iLI�swg�L��O;��*�f]m��ml��v��ᗺ��7��]J=���m���|��|�����T���޺�d�5���=wW>F��;<,Ew����D^�`�-'uF�hP��P�I2WQ3�H�����3�)�uhfs7$�xZ���&棞:ք�d-B�GH�(�Cd�R0�s�w�.r�@iQ����2�j�k����+5%V�QiTC��8DK�)��pّ�+2Cr	�+��]�<�1�e�,�U�**����[�Nf�z��.#����S���괊�G:S���*�=��W7nl�PY��Efs�C��&C��y܉ՒQ����IӢ�rD�r�Sw]ʩ�y�"��B�4�2��3���A���5���K�k��H���!�<�t2�Ow
�c�PQ�%��	���C��T-Q
'<�V�/7%�\��:���u̪.r��xTI��W���Kr4uݮ�g+�PS/$���L��P.��<�Ȃ��HV��E�B��W*N��J�sAgW<"rB���8USs<�ʪ�Vg)���JM�=KR�Zc�*.�˄E�vfPNv[L.�HU��fQJ�z�Hi;��Dd�D�5��rQ:u����n��ke��6�����0�
[q\ɜD�R�r5qv�R�f�w�3N���yy��S҇�O-���-Nu�)(�zF�hfN��%�V�.�C�����|�;�aT]�7��7�����}O���yw�S���!�>��C���7�C�?!������c�O��һ�i�I��?&��F>�DAXzeD��C�`E:��uk�ҥ��O�!�NTߋ�i7�'{v�����˼;N�������0��{�rH~w*o�W��}N}�����;��'���97���}C��8}�9�� }�� ��7i뙛sԽ���*;�H�#�b=s" ��#�v�w���S!'?{���&�Bt�+���׀<��'u�ǌs�ŷ���;��R~;H�weۓ}B�o&���@���3�T������Ʊ�_��a~E{}���",}$G�#H�9�� ��#��GtS
����ɿ!8?�x��ϸ��z|8���ݷ�yv�;������������r�M}���ׄ��On��2"���A��Ї�w�띗'����x����=���oL�<�{y\�|o�x}���?���ݷ�>���=n����]��߱��n|��a���<`Dߟ��z<}�>�C�z/���s�N~���x}""D1�"Dn��8����gM�٫o����DP"G�D1� �_h'�ݼ����>����i�Oܟڃ��]H|��ɾ�?����|����ף��ˉ��L.���m�$?�ʛ�����p)�����(��74�羛+w(o���>��D�?ݤ$���!������?������0�o����i�L/����~���?�����	9���S}Bq8�o�<x I�!'����\y|}��"�D���ExC�ڗ���=�i�����I�����ρw�i7�/??{��*�]�}��C�A���N9C�&���?��]�7��^�~��®�P{O	��&��~���!��C����!A|G�A��e�s����~Ij��#�M!!���׃yW}MF��߽�&O�n?��M��O{��6��ݧ~^�����v�tro�O�o�ϭ��`�����=���S�;�<~������P#:>�9�v������������={��������C˿8��o��ӽ;���;���aT?�I�~���|C�a|��~���%w�i���zOri��ݻ׎7�<!�5ԞOܛ���G�-OE^��j�dӃ(GnP�r�El��ٕu�H˙Ԇ�%Z�\�lѻ�st.�L�ag��`�����ƅ�8��ނ���>]o��}S�o3�r�����bC� �ϱ���]-�]�����+S���֯�״�Qx�+p`�6{��!��r�������`�����"DF��G�1���_GϜ~v���'��!�0���>��~ON?8�@���������7������w�>;���~����������or|C�u/����۽|�?ޣ�y@e[����G�""D|EQ�#G���Ǵ��[͎M�����}�6�w�=w�����K�]�&�~����o�ֽ��Ͻ/F�x�5{�j=�x�:�쫲�����Ły��|�D�� �?|H��D<e���9��y�o(�v��ώ���ܚBO>�9���<�����>���?x=~��n@��������>�t�DEc"�:���u���$q^[��`�!����/f�k1�b4��v�>Ǆ����
ro��ro���������r}O�xw�����7;�!�c>�ݤ����ʏ�#�½9n_l���5?Nr�]c)��} ��|G��S�B!������q�4���k��޼����w���}���P�8��| I;��I��y��90�����9��Ό>c�B$}h
kб�0�j�>�<V��� �DE�G��b��@���>7�zC�}C���[���?Sw������y��׏�ޓxBt��~�yIM�<��'����<YM�"��D��|D}�0�{x�0���_�_�����ן������S!{���|�?x���?<�������aw�.�o&��p~����$�����᝽�!�������;z�㷇}|&��y�}"����t׌?nU�I�m��ǯ�>�����O��ǏPrn@���v����>�X�������z�;�S1F��ṏ���|�}��}�x��|�����}����{<F���y��#�DD,��M������'yƚ��_}���?߼����zq���x��~w�9>;׋�S�����>��90���P��ʻ�i�C׾������>'�c�o�H{C����ě���~v���}#���X��|G�����G�����R�7�NNz ��� ��{��@G�DI�����Ï�'���7�?!�9��z�zO)��P��^��'��Sϫ�����8��~��_����ߜz@��o�/_>�=3��ߐ����|%�?���>���<3ql{׶�K���x��x��Z��dc���U\Hos,�<������}/\{f�a��9p�W5H�V#/r:Źy��m����w5��ʞ8�V�	�WԆ=��K%���`���]u��%o�=�ݘ\O��gvjٟ��� ��+�ՙΪ��������>}�9I��>���xEӴ��!�m�ܮ=�Aɾ�[{OAׇӂC��'�����S���v?�)�|���:Wo�r��?x�y�uX����E<���} X�0DH�%1�F= ~Iǽ�<;ÿ���4����L*�i�߾�������xC�i7���]�3�8��7�$����׎�
o�O�zC�x}8$>���~���hk�'#��IO�0p��f(}���;_c||;�z=��<+��|���ޓ�7���<>P�O�s�����������'��׀�C�aT<��{�)�{C�>%��!ʇ�Ё�$?�O���Xg�~������t���O��}B �������8������כۃ�[�~v�@?�z=��xw�i$>>���Ҧ���\��~Nq��y���������]�'���(����9?����zN/Y��3s5-yg%W�B>#�")<!���[w�����^,(M�<z�	���ɾ�>���ǅ N��s����c�}���{C�i�����_��.����}��y�m�ܮ�}���� ���#���S>���gv��`� �������ǤܟS�
z�{M>}�8��yI7��ż&�����ˎ@����~���˼?Ss�G��
����F��&׿�߼������nr���u��N�wy��[t}� ��{w�8<�����x��U����?~��i<��	�ѹ���xv�N��|���O�®O?��0�P��s!�>����������0��!޼�q�^�VpMV��s=2�;Ѣ#DF�G�|q��Hro��px~!��+�!���<�~I����^�ޓ}BC��ǿ'�p)��}�����|@�xC�4������s��I'�1��U7�A GԻ�0uQSg/lzb��yr^����zNq�������ӂC�����z����aw�S���@���xM�����{߿x1�H.�z��oHRM�w����&����t�+�~�"(}}r?,zDxoM�yuy(�ϟ�~������oۣ�x��]&��o�_,~q���ɹ����?�	����I������|��)��S}�'���Woi8���}C�a~�gޜ���C�A��������%��� ���Μ�{Z�a����U�Q?R���O�e�)�-Q�`�f�5���	aо�.��8ۗ�x�'9�u�\37.�T2�d�$�Q��[F�\Tu\��\�9����]v���'zZU!+��/���rK��`�ɩ�g���˿�����(raW'�;�or��~��n�����o��o��O����o�I����?xޕ���￼r�v���pI��~M����cÏG{����|x���b�E`��δk�ϯ�=��{>~�aWe޽�7�w���OTe�>'�9���S��;�oQ�>��ra|�8����{�m��>8�w��|�RC�[����O��#�"߽s���#�".+Oyr���ɯq[H�^�"$}C���~�ɧN>>�����]��y=w��ܮ��*�7�����o��	�'y=v?:O	�������yC�z��ʛ�?��=;�)���A{�>����%����A���b����~C�{;rf���'���>�}BI~�z�P��ϰ~O;H�C��)�![|O'^�������o������M������'�S8)�E�G+�_	��>�`�m�;����ǅv�I�O߻(xL/����=;�ӎ@�~�����t��������)�]������r������s�|��Ǿ� }Io�O5��M�	>$��}�eo��tw,�9K��χ }{��H��D|��=u�G�G��ޚ"�Y�����<�w�۽�v�~q�O�x}">�~J؈�0DX�"$}����`������b,D����! ,6G����"*+����UpT��3
�����,��	��yd5[q�2���ہ�ǸȊN�_zw!�a�f���#Z-�+u��>��P���+�Q`�j���P�S5[SQV�:��g!����?����N��O���3�G�����UR�s>�Euݞt;^&�Wp�-R!1�������%��-�N�CU<0k��}":n%��(Ώ:���*�n\t�VZ�hޝ�J���Z�&��y�C�p�������C���1����w�Z�4��	�>��!;�t,��RM;�.��|�<&����_̉]�^��q�*3;��p��H4�c�|��V�}*��cV*叕�-m8�d�7�:�s�����Nr�e�R��ߙ�\:���(h�}�x�l� 8Ȫ@A�̗QHGۗm�˷��QN6gLp��	���V��7)���ɍ��W+9���L��*�M^�����T�g�����O"�UHw;�����r\q���T��V*�C�)4�i!ذ!�q=F�쁪�@�I��<�����֊5_/���7�gQ�Yԧ/s�K&��WJ�m��>H����޳N����&�zJ�u��Ё�.�[���{`�&���8K�&��4��4\	F�Ct���C1�b3�tТ��9��9p���m�V����K�G[�L�AwXg�ހ"����(#�jeP`�����+�+WM���T���o�����8XRb~����>GW[g�p�򡤿���y;��x�n���o�J��d�S��;�RX/���1e1�e�<�Lo)f�;�~l�j��$��䨣��l۫�z�cX��%��5�Rn�mT�xb.�-�����b���+��	1�//��h8Ժ���ծx��W��]$e��ĕ.Y��A׌��?zY�YA�"���zr���m��RkKg(�/
2��n����;jK��!���[iԵ:f��/�����E7�Z4�r"�;��&
�NGx�ZX���yh_8���Ӱ��jjEZIbZ��R���ܢ����rW��Evk�׬�Vy`)�\ [��<wĄD���i❾�=V�=F���ʐ���?���/).ӓ厺̿k�Y����8���Γȶ��+���+W� ����]�VyV�3�Q����@X�M��xOT�p�X�[�]�RЫ�Out���g��*��굿)����	�S����e!��g��F͉K��*�\��yA<���9�qY���!�:����/e3�W���n�|���(�YX�ܑt���9��׍�ԾB�e��o@_TU���J����z:�wJ7���>?W�=�*C��D��&��M��T�����MV��d!�骤��,G߻.�At�c ����iײ�<bɶ7WH[�'�8ݖ6�Uw��RMA1�'� �)Wxy����m�cf��ruE饝ؔe^�?�nጃ�Lv�΀�?Syp���������A�6R�aː1؏?K����O��B���.��Crr7�'�U#[�� �ؘ(%3�lT=�=K[�Ï��;�x嬤G	ؑ��Y)Pf�6�䈁͉�'0��c�p��T�Ĳ��i�^�(ǹ�FnS�}$D�mf�EEW�X6�������9��7��oܗ�r>w�]e6ﻟf�w've�ʞ�c��p4 Y�'��:�k�c���J�}[�=�F/�1�i̍��Ī(-�y�pC>r��_�!S��3{����B<㝳�J#=T�W��|J���,C�jV��-'Hv:�nc �	��K��6F�*7&ss[���`�s�����1�]{+�~O���xf_۪p���awy��7����Ѽ�gl�Β��j,}I��j"e��S�s�nvN!��c��{��N�3ZÈa���sT�n�0��'L"Pܳ69��څ�/N�"�����=0N����\�FǾӴ�?y��1��K"�8>��UB��G
�+b&P��WY��^k뷛�O�v�����]�Zn#K�o�鈘��p�3��*!�0m������A�)]�:�ȚT�y��(HN]h�ɡ�X�7�F���@v��#�ub<�{��)wjfnvZI�)�CI�HIB\D�1sXP�a�� b��<�٪��**|b�,m�Ԫ2d��9�9w>z�ܼ�	��^����#����CX��[G*s7��?v���c5=�D�܆�KVJ03ִM[-(���}l�O.4���H��eY[炷��3�{]/LAvfAڮ���VI�8��U��e����l�Z�:�>�z*=���n���Ńx�[����n�ͻӍ��U�MM/��5N�l�҃�
�j����z/O��v�����un7�G*��g��
��"zHA)3�lN�� �T;Z:�Jؾ�/�	dV���U�@�^�s��_ޏ��6pw�6c��_�X�)��4}�Wy��"��+�I[u�LO
�x��>�y�鳑~c��(GD5V�Y�R@P9�q͵yS���͵��j��o8�t(���_E��[$uBT�
��;H�8�l��Į�k�;G:��5c�ݼ�u�d�:�?)�uP�y�ÅL1v��V�_�P�5��Ra�^m��Z}��?w�ӱ��v�zn�7����F���"�/�p�[�y|��%*꯯�נ����[M5���LU�4�o����+Ƽ*|OiȐ���T���fa�0y{o:��3��lw3s$l�q{��\7�l��
�x@�z�!�;̊׆����c�[#�У�CǼ��Df��ioL��[.�B1�yD®���ϵ���&O��$���xLk�κw1�(�=� �|� ��oy,u����#5���5�t�ӻ���(��8v۸y�$�lŲ.}E����m��Gu���ئ��ǰ��W��^����1(�o*���5��璥(?\�cw�Z�y*�n�=�M�[�����]�HE��;�;�;BE��æ>����L�}��f�1���euYs��2�+<���K����g���GUwcj4��� }��F*K����.pP��,��� +��yb��B/��O�C�˾�;~��=��ّt�S�ߪs2
^W�F�[�n�A�<*� +�c��C�"���Vbn/���^;��P�V/ջs�e�bV�Y�#�}�|�Ե]Qn���f�y���ڟ%�*P�<K�8�v­0�����	���6J:�/�K��L���!o�O=�[�J�OA�C -.$�1���9���ξ�5�P�q��϶D�du8bz�蟦�u���a��{��6�c#L&j']Xy ��rY�+��
�.��P8�)8rSʳ�-0?FTK&���� (�@�q(	������tBʩ�;������G��r���T�0��:+K���^����َ��U��6	�M3̭�K�����m5>p;�mblU*�Nԥ�3<xb$c�v��~*=�Xt.�[DQ�WYa�o���w	�Mu�v7��.�PS��-��*O�/����ܳQ��mA�H�թ�G���J[=�&GZ�n�Mѡ����7
�]7���!t������|�f�<��뤥���],t�����_�v�uQ�k0�񼑲�3t.������o���W��-ÿ%�*_��F���v��.�)Zɮ34m�q�@���.�o��YC��@X�(����U�+�
M��~й%q�f5��{!��U��+ऩ�7(p���A�
B}�k�{gUmƊ��>t���} �wN@!�I�����/��rr%e��Qn`/�q�w/�7n��Ӻ���S�+I	�c����9�ei���c+����==�@s,(�m'��۳����K��D�9&8mD�B�ʌ
�'~`"c�Pwʬ�!��&�|�styj��#�%�C�{�����Ū��ȁ�?c߽��W�^�� ]��3of����|�j8�p̙[���5ו B�v�����v��,��/M��m��u�Q��{�g�r��^Ǡ�5W2�e/����d٠8?�V�^ �ߘ<p;��ʫ+b�#�+:"-����n�J��q̿����C�5Ӟ�XlD]�t�|�D^v;�n7�)�A1�sXz�g\Ʋ�=��܍�l<� XZi�W�J��P;Cf��χ(�T;�,C�x�r��E^!7�J���K]1�g�~��v���{�*L�D�A3���웑
��9a�h� �j��#_���ۭ�؉,i�����5v95敺�t-�����iRm��q�L���7Z���ԕ�i�ǲ��뉨྇"Ɇ6F��Ne�OWb3&T6��[�qi���`6oqh��2��͞�-�����OS�x�5
��!�k�ɮ�zq�L�M{�p� vi���luM�Ҭ��'��ů�"��]���}�RZIHۭ�t�A�&��&N}7*�Op֖��˄��Y��ƈ�����԰���!<�C{��_7v���L���ۙ�e4q��6{@=��s���L��&�\�#a�<��+���{��f-3F����̮xK�:ԧy�_����^T��ٯD_J��Q�V푒Σc���Ryj��R��ykj�i���9���ܾ9���Ns��i��B������q��,�z�$�������|]tB�Jo
� ������"��2�R
o��e�[���ڴ$�0�y���>�m�T6��PE��:�]Q���2����޾����|E#3@�9�j{�*�䫺��T�^e�L04��:�7�X�����ڡw�6:\�)�(���Y#m>}E�9��j"�Xb�0W5��R�-.��ۋ��Mdc�w{����9�3�oQ[2���{1�ZC/��y��<�*8��.�ꚟ7w.��k���v(�%r5egDg4p��Ŵ鏸�VhP٦����A��z��TC���E���^S�A�e���05ׁLF�mS&��c/E��v.m<f�n�Eҕ��(��f`Z��jҹJ�i�(s�a��wuSe]dB�)��S��6.�;a��V�*U��0],kf��UA���uj�A��]�ceh�9A(�}�u�.���k(�5�E�)�Dݣ%$ő�9��5�ZB�ut��nѭN�0ufk�u��Tyѥ)U�zO9�yw3z�mr9�Y�om�+Jn�&�#Mۥ:!X�ILq�̼�vl)�rf�y�t�̭Z��-��I�{]2]�m�Vi�\�++{�D����˜ݎQ3Z�JR�q��"Iy��(1p@�+��tr��R�;��`Y�]�@��ud�T��c���	��X���A��V5>��,�lY+��5 ,ElZ�hN�Y���b�f���Z.��ط��%�LP�v���(R�en�X���^��f�M����7��i�]�:v�c�]���w�3��tn�=��� ������,vԵd�q����R�8m���}Lѣ��&�q� J hu�=dhR)&�*�B��Ӟ�NY��#|���*��c��F��>M;Ere�GXr��r��w�/�y9�z��ׇ<��K $�:�0�:%�J�}���e�J1�����z2qӣ��K�7%o�"M�ڜ���ہ�t�s�uw.Մ�݁�PI��&^k��%���R�(
Q�2J�9��+p�b*̤"�2k:�ZD�Pt�Gq�V�fN�[7\.Q���uIwePPTDz�\�'��In�&W�\If)r��ML̕I2�QR�.��tH�<-���1�Ȍu�T;��s)B�OG:�Z�edD��\#���$R��D���鲨�DC��]�U:`���(s ���<����9:�Hx�)��N�ZW��IHT�YD����$��W�&�����iUBqSd��ꑫ*�RHs��BN���"ʌ70�ʣ�0��YW
�wK�"��2=B��%u�<�U"wp"�r5+�s\�p�I"�h�ER����0����z�KAdl�M[�9Uf�:�n�K��r<�u��e!F�	�w'<T�f$�N;�wq�!9�^��<�rv^$[׏Q��^��C�����\%s��Cd멕�(�9����E1�&�Z]�Z�}ʎv%�h[�g���������/.��~�ZO�ה��#�ƾT*^U״�t� ����kt���xy{����� �q�=�y������&�
_xz���L(1��>�9�*�����]�I�a�V���7-��T�Uʋ�GU��8�ݸy������]�����&��"��~'@F*\�6�󧧜o��W��wN�yM����@�����;H����Z�bsփ�7Dt�@��yC�+�r��z��%�|t'��H�.y�v��i3o[���:S7�h�܌*�ǖA�A�����Y6��O\9��-��mD��u���4���1��m�w#��=Nb�L�u3��n��s��ǖ���q��yH�~�v���;�8:r��ς.�j%_Yz�W�J���DT���;R���agU�$ŀ�:�>k�h8���v��?eO,E��^Z�18�����_rY�t,8��-��dC�Rw�n`��LI� !��ls7�n�";E�<[�J��s��Gp�70�%�l73,�b,i]�6w��p�T��Yڏ�������� FV��ɵXN�r�^Lޛ&��|l6�6�r�eaw��)Q��]��b�U�w�Q]��w7F�;������/,���u�w]3����֧�`,�dri!�r���� �ʸ�w���l5�gv��YX#����9b;�ﾯ�����]~m�y��s�7�᥏^<�I�鈛�w;��x� igm}P�ЅM��-o˽5N��~���`��`��[�r����f}|�yK��l�5\1&��r����R��w�s6]OR�"���'LẂ�j$��"a_D��x:��u�o�|�(y�������31��^������_]o3Ɵ�B�1������2��}��f�L�F��0���U|��	�f�|s�n�u,oB���\7��vFȞ��J	M���:�m��h ��c֬*��r�%5?\k����1��Е_F6���� ��V�L��^����u���_�Ԩ	S#�Yh���ơ/uÄ��O�v��r�T9�lgNQE"*Zb3�2'�-�W+�G V�ԇ�Ph�|�H�S�D�$�6cV*L柰nrnkZ�����uW��uZ�F�٤K`�j���'��8T��XJ��i�j<+m,v8��wwW>����8�[���pU><MnU
=�"�[��|M/���3�{M\�+��U`{�?-Mdn.��]I%Z��`�G��ji\�#z'iY��xf)���%�Q:��`�uà����ǶP�E��gF�<j��S�g��]*NFee�b�f�\oT=�Ih[Ǚ9�Ӗ㥭�ٴ�-�[��p2�`'���U�Ra=aN��᷄��6G�}|f�u6%�Cjp���J�E�{(��V�AfY�pJ㤁�rx*T�Z.���b�w~�r���ګ��|�qb퉎0�ŷ�l�n�����:�o�_ZtD
0�e��N�հ1E]\��ߴ�r�#�Eh�5���u�5V�����n����0����s��^��y����ޜs:����o�q_�p�o_x��o�b����p��Î��s���YuU6�V.�m;
�H�6\�_D��(���aUs��Tb����yd5[q���|���u�:N�۾���վ�p�� �=5�ͪ�u��,+.�N�i �QM�Mޝ��\��u*���k�,o��>C�@n��/��W]���7��au���6�l�M��"���yt>�N�(E#����W�]pѐ�E}:e�\,�S:=���({���&���i<W??���Qe@�l)1���x�߸����p����{�t�}��w�s��X��w}sw���x _�o�SvWJ���f7ά<����С��
�Zj��%>��_{XŬ^wGv��GN�no]Y�-]U�謪T��U�FX�0����b6k�)�z뚬��c���X�ޔr�(o�50y��/'0�q#�u3F�������r�|����4W\��P�X�Ҳ�����]�*�@I͗5qō���+ꪪ���s�t�`P8�Ф	�S�*�`Q�rl�B7��Cj���|lr!�ӯDiN�J����RM��E�v;��#�c����H�$\4�g���]DB�:6�%��������@t��'�?��gA��-�wi�k��,��1G�,9�w�:7b܊��R�e5ͼ�4�-�B-S��Cr����6*9@!����願k�+���P��-�1w�vY=�w>f�a��)��2�/+Aۯz`��dW�Qϒᢛ�%en���V;ŀ�N(|�rw`<���,)1?ki\1�gY�7�����X�ѢL
͡��<�e�R�K�0���E�=�u�z}}7�O,~:�^�nb�n~|^�Tz���+'*��<���<22Ox����#Z1��U����6MiCI�=�Ud�Oa�s.����%/w����
�q�]�0��ӫ�� z��@�ϼ�$+��+�k�;o���8�p"���[�yJ( �+'�t�����E	X��p�}2����,7���u��Ȍ+w}��)��}n��k���v/���$7º_�rʞ�v��2�uɆ�ݼ'TT�m��={�Z�Ƅ��HF�q���_�αEq�!��Bj�\�re������jpq��Ǭ@. p6��k��En���}}_=��'���BM^�?�/$��O�S��}�+ݳzX�lX�M���gon�f�i�؇�����i�&穊��3�lӞ�&�g����x�����iz�{�e�/+�OE"��d���G�+��\ۚ®2g\�ꐌQ�_e��v�e3�TY����������c��H�-w}��N�*
�-y@r7�(�Ã�%}�o#���[}H{�كQ��y�QRr�̌Ű��|`�L^7�Y��p��MU '�k4��������AW�w���(��8A�C���
ˈT���'!�?���5�P+��>x�k3��C1f�HY��{�����<�'P��c�5�)��b��(�)@F6I��ӓ��Qr�d������qz�����}��B�]�!�9lN�6uPBYu�b���[�k�����.&Qs$��1p!�{�I����gBd3#��r0�����a��<�ԭOb������R��IO�xX�|��p�/Rv�gΩ[��T����Ӊ=�4��h
��r��1W4�V�*��i�f�L����N��7Y�/z�Cn[��`x���ژ!���15u�'�k����o<����	]-Z˔��h��Vg\��][��ۦ�K)r��f�x���=*W	~�#��1.�+ӳ�vg�NLB��������t�q������T����̺�7����m���O�œ'�u�򗮲냌�WF��@<�:�>�����2�u�-���"/���}M�4qdzfq���j�FKݾ-�ţ"mHyN]�0��Г�*	Cr�3c��=5�c���wb/���ހ�;���+�e����!���T(�e~�Y����]��Ԣ�GX�}c�����X�L<=�J�UJ��J��y<���rx�@���'t�<�5�˩|�g}YȓV-���\�LV���ٳ������UC�[X��5u���}��'ְTڳ��v�>}15�GLWȁv]#½��\"����*�w��]�,w�1�E�Ӓ���t=[� q���q`�^��u��xԫ���F��t�w�����Nb�ْ_������M�σcDfr��Ʃ�3��뒾y::�D���)3�f�	кW|�W^㷕khfLS���ymT&O>���5���cS�cE�����["�W ��z�ik����;�#hT�ʝRH���Y̓ث��g�]ˣ!�Q@�K)�97��=��V�����D��*@�^�:�2wI��o\�eF\!=�;��h'2
�_v���I���o]��ٙY��ފn�6�����KPt�BT'�G�}������ J�}G��ڄ"��2���Oj%9l�0���P�sNМm�Gw*J��&ef��BI6���"�Я�� W�(4b�l��
xh�I�F29¤μ	7uB�e���K+'�7%w�7NJ`�j��PO3�s�P�eS�_yM�0
)c9�z��c�=5�5�pN�|yz������Q�ˉ���qȩG;�Le���]Ÿq3#��`8���m��ݮ���Y�u�z�y�@����J��L���a���r�,��Gi����+�G��m���]t~���[9::�) +2ȸNH�1�{�c5&�|�$3�������9�/a�3�V_o *�w��y����!Q$����4�4�k�����:xk�����+�N�)8��}��d3x�g�Nm��a��������6R�p]uv��W�οWg�V�U|�
j���+��rE�/]^"�|���� ��5�^�g6�}�d8j{�[�W�֋j�pp�,+.�.���sYD������b�=i��X�%)X��M�<q�Yϳ����M��g�M�Ӓ�Bͫ��J�ZNZ��V��MT�hM�v<z�+ˬ�u���8@�l�xJ��� ��m�����oa��md��0`Q��
Q�"��F��co��ݿs�*H��v["�)��u���b-��o�}�}�Ր�no=���<pV)"�:��2���ٳ�e�bm��e#�}�|��6+��Ć��U�w��(j��{�|L�S�e���O�tz0{l/�ԸY̗�7k��=�=�9yxw(�Bޝߝ��6g�J���ҟL0����`ߞ�<�x�7Y�Vf�}��(�$8'C�Up���(��bYs��nS)��ƈ��b�i���V�]���g���8���b����f�7��Y3!����t�pE���V�"��=��#і�!�{�O��P�u��*N��7���1�I�y���Ȋ�l�~c\��֠�](M�f�X���?C�j�6�}�>H��Ȫ�1Py�B��3V�v�C�#�K����m��Sѻpz���	��qoe9@t�E7L�,3_�����{^E�O/d8-RÄ�;��|�D=h�U��L�C��9@�RDi;=&=�B��ov�KU��wv� !�G����9���8XRb~����͢��Ҳ��V�Ψ�ӼT�9�ֺs�䛣sx7��]bĵ_u�h�2��ӻ��Ỵ��t��{�w�������k7;��,�=gs���3�$��j]�v{�)�]���u�Yhl=��<Z�1`��]��b�D��@1]4U�Q�菢#�)7�<;ֈ��� 2.7�t�[$-��a�ok=�U��l��e\�]U�h�i�Y\�L�[t,�<N��[�$�',��h֌i����?���X�`��n.�=jg���Z�Q��:@�
b��sӭ���(u�u^�و�������[�Hؼ�y"o��N�w���U�`�D�)<�AQ����ٱ2R]�"�]e�{�?>���H�;��yV�ު�Ua�g�qK��_Y|@�ޘ��PY\<%w	5z�9j�L<én(�N/�x�k��p,R.T�ˈ�ۇ����LF3K��ۍ<��S;��A5}qGb��ɲ�:z`��u�K �$���A:3eY8����?^B�l���:\��#�nb�Yv9�:}*�m�?1[�>^P��
����sjx+����p��P��p�w�XUڻjgO���qM���Q=�m�~��5�U
��N��5�@��j�H�4-k���6ժev�W���������.!�cT�pTxL#JB�#Y�E�{�j�׎徒����"��c#݌t�Ք/��s�7xBŒ!�C�nax�o!F��KGM��ƭ�L3/��R�n��p��j�K�g:��ԙ�v��}�:�zY�ާI�ړ�?ϗ����r�C^�OP��gm@�����JGj� YϖA�E��}��}U[�M�����w,'��!W���{P�'Q��D�;�Ց���CvJ*��U[T��С���O���֘�tS��Ơ_t�����܁�86)ҩ)�xM�Ğw1���[c�@ųs�����%K��7v�e�nb�N�f���&�S�10%�3:k���֧/��<�w,�s.H�p�9��H�=f;�!���;.���2*"f��i!���W��ܑ���ޒ����&���u��\�bb�TH�X�f�x��s{����o"�snż�`���xΕ!��ց��>�^��ϒ���:�o0�
��\����ԃ���TsGn���<#������X�.�Sj�}�r�1�����u�������A���J?'�����6^��1��eBf�̶1��dXjf�p�c��,l�fU��B���$?D�a"<*���d�l��C�3�q�5��r��Q-���.}nb�AߦjS��]������r�NI1����t��i����/��)Uz��Ҽ*US���t#--��\Z[}�Eawx�:��k_U�CI^�I�]:*R�e���.ƹ�w<�e
Љ8���A��=�]�N��j`ڋR����W��V�N�.�oq\�H���8�[��������p͖o,����������w�[������G�O!�H�����n}��k�+y+Ň.�r�\���x2�[S*�o)l�SX���%�f�g�����0-�I5�Y1R2�cU]L(����Y�%�n=C����Y�]�o�
E�o3�r��tF&��ڑ�` ����콵t��+{\@��q,cI��P���=���s�'wV�x>��ك���ڊ���:��
���C�m�Y�o0hn��s��k8]GyL]�u^���w4P��(�H�5���^N�Be>���s0Ql�!ˈ�,0�*�^��C��폥7�ݛ'U!�O������yˀ����:�Y3 �%.��"�-a���>���I8��]v�=�l���;siA�ݗ��Mo	;��s���u�٣0&���r�ŝ��x�or.owXϲ����K���M3�	QpI��]ww���1�����|s��q|�����i+H��^�5,\8����L�T_/��!T���j���bҮ1K2�lZ�R�G�9k�R�o#�B���^e<ʾkuwdkI����ۚ�Sv��Ɯ�)�-�N�&�Sﳝ݌话Y�|��<�	G�9_Q	�rۈһ����ʃ�VŉaN�c%X�!:��\\-�f����ǧk�Xy�[��v��k��yA��P��Ic��@֊Q4��Z�S��a���(��/_�U�<F�����"�������+��$N�#o���;վ���\��j��f��5z
�K�ymb�2�{�����a���c:ݗ��Z��/�x��f��3�-V�yZ��L�E�@"V��s�V,I�:ƴ���#w�n���Rc��ɩ��uaJ�%�=�Vf�Y�^�ї�f>�>b�2���t�*�^�U}%Qw{Ջ�䛚Z:�n ��X�ӓ0Y����݉/h�lc{f�\���Mom�sk����̌�3mܫ�lK�XL5[.�����9I�[���\��x��w;�Y֧Fp)�ˮ�r��8�Δ�Kt-��]"k�[��ZΉ�۰7�ˀE{3e1m�9��O1t%�}�������i^^AȄJۮ}&:��_���l���w~�"%X���(eu��n��?X��S-f�]�G� {
��R���H��:����S3���H�ln'Вf��iK(�ո&>��q$8-��-����0)����F�L�.�ᡜ�披9ll��"˹��[OF#�$���k�Em����&��5x��@v:�u<�Y���˺xU�3��2�u�Z;��A4,Y�{��8E{�XU���0#$�4��E��8�$GV�w<�RON�T�:q����$e�{��TR�^:㧗�z	Z�jHz#����2��wK�&W+R�QG13tOH�5���2#s=D�,��ҺQe�IR�-N���)�G1�\��7:�VjDJ�����T��UUj�-�IG",ʕ%��%�-,��G��b�*2͖rԲ��D�J�u���(�]iz�',�t�̴3J2��!C'@�e�)�L�H��%���H�LȊ1-Z�FwX�V�DZD�"�wQ��4$�<w1		M�Rº�,��.YUYQ����I$�D�����]�DRU%udiUk*�D�,���u�5IVfeU%e�"Dh�WP�J�D���r��HW��y���|��sך�ee����Kќu��ݜ�a��xj�1�I��wIuW�G��Ǌ�7�j�5}��9UU}_U,ҟ�s~V��#�I����*+�m3O���t�
�ʥ\"���-*�uW�U*1qWk�q���U:��{a6���/���C[���[e���o�j
ƕw��k<7^��푘�=���9]Z6�Os?h��Ÿ��k�kunUx��'�g�W�� �:��v�FT7.R�rkv��[u;�����g"SW���/K♍u(1J�o�GNQ��k��ǯ��|��� V5y�|��Vyp�()>�k��6t|����]K5=���8��˼d|�Sݸ�!0r@޺wB�*P��(4a}�GUrс?�w����`�\A�v��d}�劂{K���b�rxg�#F�T�9���)|��IC�(�OS<e�Gf�|д��qs�Ok���#K��]<�A�ao��&(���a��N; �mۧϒ��1k���t��}4"��+cw�;�� 3F��9�|��7qV�8g5�����T�ע-�*7���0�oܘ���(�@G���b;Ȋ�T|v�Q�u�����U�����5�at�#�������sY�5��l��"�(i��r�^'{�Hfn��Y�k�(ȡQN�r�� @�+�,u���a|v� �P]>6�k�>Q�6#qR��QwJ:��ZJ��|im,�]�ce�R}Y��c�B�W�����J����W6�\�Sqz��z#��">���x�N{�~�+�-�9�.����ܫ��@F�'f͵ 6n����ZN���WG5�Hq�:J܃(F����Y�grP�3Q�(;�<��ᩂ�_c\ݡi����9f.Qp�n�`yG�8@f�J�
`�aVpH��R��� �S]�&__6�w�T�pu�{��6���m=��,�o�1�*r�J0N;�^lkKZ���Jc��/+@��7$Z{H@jpf�쿤R��Um��eR=g�t��z���DS~S;�o;�*!RE����3ڈ��s�ei����ˣ]�rӗ�el��U�8�_��#��z��]x7=��sT'�c���r$)1x������~�.>�(hW�p%��I]�w3�K�Ł	��� H�xp;uH	���,%c��&nRw��Cr�H��oo!�:{f������u���5zji�U���^'��Nw�����W�*�;i���,|rV���X���w�kU��6i��N_�U�}>�0W
�Թ�G��5�	x�9�}�r�̗��*�2�k��[t��+��6ժ�����+Ss�=W�g]�Z����[��v���n�����v��y�B��t��;
�4>�^����NU�����u�����}��rTy��Ƹ�Z��OxN�6�K�[+M�xs����}���}�%]=�����V�h��78���`n�ã�LW�>H��}ٓ%�P��v�y��3�d����=вㄊ�N��7ԉ�� `��L���n��w)��:�T��.q��ш���_R�G3���Ҩ�uP���o�[� 4���4\�h��ަ�J�����e�"�0x1��;�2		�ӑ�5��7�\8���q�fC%<��Ǽ�M�v��VXn`,��7)G�Ȏf����_�_�W�(�^�S�ͮ��~Xu��BC����_n����z�E	u�^'���֌t���n�s����|���'��9��3UoU�b�銆�	1���Ѕ��k2"N��}��쎂�U85ArrP�SP����S�z���j���0�K_�UJ�8� ن�(Hj����	�3�}�E-�λO���ޏv�noΪZ�������W�qx�6�i�oL�J@�2Vj�K�חP�s�v���@0W�6P;.��\�v�*����.�:d��Gu��EDD�1T
����,@��z�MKL����3U\�u9��Ƴ�f��λ[��F[��pW:���[��Éۗ��d{%�v+e
bD�u�T�Vr�t���$NB#�.H�R<��K���"��0ɻ������YMld���>��U�}�}W�.���w9*�2D���`���8���u�b#�(���˅���DS<KJA���pw"X���� �wo��3A[��P�7�*��Ã�_y]<�Bx�&�������.��<�֚������Ũol����"����DL������;���رJ]����dL�W�*}ݗu0+v���̬�1�bC�v+P�O�ͳ˶��U�eio'G���|�C71�wP���Wg �f��M�H�G$:3`��,1S���h�/.�(��W֜�m�!�Qr�]�P1M-�ݿx��[�^ݑv��P oZ�J���*_�:�om&n�qW:8��ɗ���8�R�3�",z;daW�-L�@��Z1�U�q�)���٩��Y_'�5���hi��aR�e�9�b#r��%�y�{OE��/J�k�(i��&�`�6g[�]|��oMp�bDX�Iճ��I@=�� �Zb�_ٺ�͇�`Z����J�#,ʺ�\3�s�93��+)��(PYO�6	��gu�v��7F�hn�A�sن�\·j8p¹��{��f��vsXB�����yX��r�Fd����:���t��������7�� ��֑'v�9��M髶J��Y��Ru.Y�0;�G
�Tl���>�>�O�w0��t�O�G�b�^R��Xu��
�x� �9˱B� 	<`ŉ9w�kޒ"�͝m���7 Met���0V�3�	���-�J�Yt}�b��Uw��e�*�j��n¾R4e��Lxe�^fR5���zU�x��(�]S��w�(8ֹ�Ei�_�>/�<e�E�}�_'s�w�p��A�Q9He�M�,M���s�Pms�*��c��*zC;�F��z�� 5^�ƴ��b�He�½�W�vxKJ����kyUoe��h^e����X�ҩ��j_�s�[y|;�(�X)�#j&a3��e�*��ns�8�I�U<�`,ϼ��}���n��t�Z���\7��vFȞ�Ζ^�uì�W�1����5����Y#�Kj�2�5\e��rQ�NXЧ���{UW��Kx�VKQذ!�'@��:����UE}�<��3�$���r�z~c��9�、ٖ�4���V!��J��s�QX���7�)� ���5�H����΅v)n�[�7��C�z76҄������{%����:���5�ʐ�A��j��l�J^Q��ާ�WL�1uo��+���[�ڕ���ӁT�o<!I7�$�����S�ޝ���,�[��I�3��U��r�N��m�u֮��|z
�6P�����>�+sy��eL����9��#EE�!TC;NJD@�(S�h�g��a�N	�ȼn�oWgc��l^o��nu��:��h}
)!Q� �;q11���U��F&���`q�j����sLe�2������U��
���;�#b̳"�\v`0�E��t�e��%�qq�&&)�m�L!�|j��L_��]�n@�PP�7!��^rP������D菉ݡ~}�Z"��5ۢ����l��X����z��h�Re}�ٳpڠ1U;�:�<�ԓ���Ve���I��(��P�!�+�QyLN4��wJ�I��ҷ[���+��b��<��Ki褥`C���������	s*"N���P���sj�Tb���͙l݅y�R�,��g:ێ�8^\Х�1p��nLpÓdYzPN�w{Wq��ԕ��H��5������/yu�3�Y����f��\�-��Ӗ�igq=K;v\�`M�o5�k��c�k�֤,���r�|c5�v&���z�o�rRZk���M��=;�]G�<碝'];;{Rh���ط�~�nz�/��^W\���C;4��:�o������e������,{K7i����8���Ƿ`h�]�J��x2�Q�YيHG[�a"&r[U�,)ø�w��>�菱4mpk [����l:�J�]{n9T�{����7k.�3�*�hL^��%5��y�2O�pډQZ�E�Ml��:q�^AW/��Ը�T���ڙ��j�Ӛ���_B�L�:~�ΡX�L�����KJ��M��̗!+�P��	�j�'�g��J���Gf�S!F��@�}ҭ�@r�u���7s�������f��&��S+���6SS\z�u]���M��S:-�����MI�L���ϐy�����-�Q�Ū��&�N���]Y��fLWL��w�ٗS��Қs��y���Cr�@T�u�ݭ���թ�T���u�O��V�\�.#�V�Иن����WUQ�NV˶��l��kg�K��!Xw�c�Y��ڋaO��2�/3,�&/�ڞ���ͧ[9p��B�����W��c�~/��.�����R�y?������.ʣ2��Ρ�ec�Ӗm3�f3��ѭ"��b�-���lffW;��tK�E*kA}.��T��3z;�(4{��6�Y���qukȍ���t�;�� *L��G�#�����g)��lt�5��P^d)��W<�q`�뢷+���7ۡ2�^�j�+#;_ٝ��A��q=���5%p��������e|�9<f�{`L9��k��+�r{��v�~�+���lή��;�.�7�����)���zq�]N򑢜m��Z���"�:���X�.q�͊ykv8��ոۂ8�|y��-e�o^{���Cih�<��}gb�Tu�d�²ӭ6��Լ��Ϣ�ߣ�����w�r��M�}��gV�r!w�K�6�x:��\�Ώf���n����6��O��Q���=%�7:����ӊ���pbY+�e��W0�5[ǡnsok���u���B��}�R�k==�맫%���3܏;����pSJ���q�Jw�)n�3EVn��<;�X�sc�f�ֹ��GJ��R����Gj%�S n�WL�j�
��v9$;����W��8	�������G2z��F@��\y�I%� %_MZ"Z2�������n���f�,��\7Ew}������U��
[N��ꖡV�MN�
�P�'��Jo@�^������=�M�9YQ�s���*�%��7>���:}��_0q2_QK��wԲ�"�j�Wp�)�b��K�G<�V��Ķ���0���#���x���g��w�>��ނ����]�S²W��HO%�©��^L���wd@w<�*�ԝ�5�w�1�=��32
-��E(�Oyf�9)B����QkL�,sK��r�뜅Pڇ�Խ��̛4��3��&�Α=�n@�YPi�E�:�{�A���?����M���F9kP�o�Ya�9]���:�/���Yk*;��c�X�w�4���3}㾏��.�qI�oφ�=���^4�A}���߭�V(ǦhFk��gn�v�{J�;;�[v���碘Y��--�q��q^÷�R��y&ߓv�@|]'���Ҟ��w��[���~�����hq�Y�w�%�W������+=� զ��`�s7fM����
3�rHn�i1�G?m�T��X�v�}��[���
�=��t��7��.���Z�L�yZ�`��N�ӧf�XK-�N�����re�{�o�7��b��V�O����������(����԰=���AMF��e{��������V�o'L��1d�X��'<_w���<����T�:��Z�N�>q��c���..�_(��n>6��׫�&UO۝C����䫖�W	󨁯��9{e����;s��3��n�ڷm�Е]
7�%̄�mQ�r<�A�os�p��O|�E:TÞ��K\v�qr��
G�JD$�����������{���q��Cz�\A���o��q���R�\]�c�E�X**�V�r��08���7�/�u�������[�?R�xקU�wkخٞ����B]s��,VF�Wy�|_&6�5n=�v�eH3X�W��,;ֈ�f�`>���ڈ�O�s��}ɋy��5�R��A��}w��e��X��2�;Zc���4���}x�,*>�}���ᾣ�+L����}o�	]�T��3JW*1��=�<�ԧsI�	˗�����|[��;��F�j�ǳzt1R�Q��6%&��0�\�A#��
�Z���m$ ��_U�p������WQv�J,��"wBv�0�,W˥�
���&�k9�LwgH�^m��C��<�)���sK�+a/{�e�g@Y�;��}uH��VF#���1u@�O)9�s��e'�nL��c(���4E��
7�>	M��V��ѽ�³�3rŵ��#�C�u0���t�鋂���Iܦ=��lp],TCnnn$�Yk^ʗ7�1��'	���ˡ�oK�걭�KxR��]B�w_2�oup�M^�������qي�7%n�	�V��&U!���-�x8��luw�-��9]}\��A�'(.�:��"�{N����eK_K�}��fPğS��9��Ը蛻��rr-Cu��y�Mw.�����h�k���q0��[��[dn[K�
���{trJ��r*4��XD�5��bx��̎�YǪ<�L��Hẓ�f�+[��e,��}EI�w%0Q�wlR��<ei��y��="�L�t�Ӿ�[���ˉ���2�ŘB�кRP�ω�Z����z�V�v��*��`��1�6(�|;��$r�4݇ݫR�y"(�W/�"cǡBr�7����l�06���rNS��j��yM��̋�V�����UM��gE}zڬ�H��,� uΧ<�L��'���M^6��S��Au�u;��m�v���qT�8�����_eXz�\=�͡����tvd�ܤ��S���ixw�^r|	����2���-u&�_=����J�p
 [�l��L���X���1��N�1�1.c����AS�tcM��*^̕�p�:��Z�oE���uA`m�ו�[��1�6��ޤ���D%�o!ݦ�n�j)}����(��V����	�ns���6)ۘsPTh�M^h"�|��v��e�����K���1� ���.����9wT�o�v�q�e%�����z�3����܍L��Z#�nT���I�|��L3������6,�n+�T�W�O�@��P�9��z�ln�u{s"�-�mKAa���r�8{�b��s9.����.�ǁ�m�/^Z���ޙ�x1�h
3��#tF����v�r5s�e�#�����)ͦ�/{,aX���8�}YJ�Γ��js���eS�@߹�ܧ��ù5Z��bv� ��>�]ܒl�RU�<�V=��}�NZzA��wFt��4�s���zB� وw4�T��׋s3u'}J�v�Wm�P��ǺC��lQ묝(��t��E��Oc��i4Kxu��I�Ս��O!����`S�:�u)��Sr�b��ǫt>���,c�(��(�'��%�j���[��]]�V�|K����q퍮�ʵ9�	%�@_{�p���]l�j������&Gi��9%�s�Vi��):NS���id�U�Z���Wػ�t��+��׎Д"���"	s��k0�J�.J�HQ�r�م](�a�e�-,)B,*���D�D$�V��U�e�I"��%Z$�gJ�$�D�$�$J�ȫ(���.H���Ia�]vz��hi�Ed��bmM�)j�Y"ZT��*�s��bJDThR[6Z���.t����YI,#E@�ht!.�)RTX��$J��V���P�%�ȕ4�2�
2,�)N��ԥB�J�Vf����e�!��X%�����QV�Q"$ �2���Y)�,�T�BY-8f�T��ˑ�����UI��C3��*��p�K5	,�C-,�R���TL��(�%�a\+H�\�+�\KD*$S2��A9�����RtVr�e�d�fDWN&�
�%Z̈�BB�K����h����#BJB��=[��II]�ʝ�^W]v�o]v$���Y�%�]f��䳤Jj��ڻPhF*
T#|	�����d%l��r��������a|�?z��=���o����~��m_K>�s]P�.���JĴ\]�b���5ݵ�MGEf�!�oN>�{u5�7�)��vQ�|���&��)����h�Rx���_V��<�pk3\��*������Z��;$�Z�bK='qɾ��p����.�ɨ��U�Y�oCW�=����]Qպ��Z����ae����]gD[�U��Yk����kqr��)p�b��/��������1�7�B`����Z�ȉ�5�{Ƈ:yf$�K�M�����M\���jgm�so�>SZ�5`]�8dc�Q;�g�|����Q�n�	>jaSq��Bz�����B���)���am(S027�J�"�ji�o���7��w;�[�4�Bp�m��|�:�l���{�):�͛&*c_,k�-�q923U��֎�}�P��_���X���"rj���6��^{_Rż�q�r����0�x���C-��2��Y9-�+��Y���Rݓ;`��ʖ�ƕf��ࣞ��]Ǟ1�n�6 =��{,����Ҝ�԰[��+Oj|j+hY��;E���ci"��l�㘖h/�W�U}�gJa_!3T�xC{F��阀���]��SZ�穠�f�ޣ�7pX�*�T�q��7h2��]�Ϣ�Jܼ��e��1�+�rF��i��vk��\l��n�"��ύ-���]�#=�ziWMj��C���W��N��Ԙ����)�
��&�e�}�Wgט�X����
y;�m��<��./8������J�<�Ư��z]ã���wGF�䣓�s<�>L�ﾌ�u���A�Q��ە2�t66~jm��2�vK��NbK�%{� ��׃R�ד���Q�Ԣ���f�����z��9zNg��k~񴶇Z�G>���~5=K>3޽溻5��=�x�y�m����S��]����o��_A~�Y�zӶ�m��Fj�uT�"�S�7���'ګ3~n��ϰlcwA�u�{�?uI����`���.�خ���/�f�P�;>�}s�J�;���*���ƃ<ݚ��	ϲ��5�U��*���I�B�J�"���9�Ԗԣ�����γy�7�[ɕ����ӭ|ܖ�f�f�0dVB,�nr`�E�VA��u�_�}U_}��>�#��v���[�hI�
�-��[���D%V�ս��r����'�;��;��I��3�ۉ���<����?y;��W�罛8���E��#��T���k����K���DOA��¢���Z:a[�|So#u��c�UM��ٮf
Q���=}�gn-�^�s�	L��1�.|zy���2gI�־Ѯ9(��|���*�
׻NQ�nYV!-���ڌ�G��a���-���ܪ�
r���8,y���R�W.�1�b���vv��@[�MN��M��s�o�Þ�q�f����e)g��Wh��A������H����N������|g`������R�q2-�8V�ۛ�މ��x�����E�;Zw9�YϮ��U�NZ����l�Q�=���y^�v�<����k�E�*�{_j�S��s~ϫ܏T6Vԑ��W��Ӟy��Y6-RAū�z������[��ǻ�D+:�ѠsK^ZݽY�ƨnR�8�s:WtE҇6�\2��¥��k]g���-\�h9g�ӖF_�������40Ah��
��o%�i�ǜ�Ws��f�Nj�_=�����W�<�������^�v�C�X��yX�]�ub�ߘ����y�VxAꃔ�Ų��nt�UϺq!؞VJ��e|��_eWg;c�s���vd[Fi.��Up�����ا��_���n���`T�bU�]�E�;�{�;���}Hs�R�����N{�WW�5�zo�/3m�M�V��b,^����Ty���_��uq�)��]��1�S�>�~^�s��ʮ͊�=����sKc�rZs��fw��u���_ܺ��>t5��֛J\�����ٽ�NR�~�
���)��=V�=���]D�2���U(�BO�F�VWVnu��	�}лo�sM�	\J~��B\-5bf�qy0����T���k/��}�W�M+�ƵP-�#�w�,u�"�;���F�X�ˋ�ڎΦ���K9ڡ��#b��v&������>�j�����Ί�!�9�EfS��C�@e!��^1nǀ�j��?�f2�b~��\�pNE�xՇ�#�-e�>��r�_P��G�y���X�t��b�A��}��t���`}���N��mڇ�7y����h+{*�F�%MKb�`�K����#����Sԡ�_b��b_+��8'ͥ�R��0�p�S�7������\�(�6oh�l�%nMF'��^�cj�w�}�Q�9�FM���ԵNftu� ���
������՗2��eQ\��r��|����W ��Oy��={B�c�	g�d��i���4��K���\�O����f��3m��3�I���9JWr�7���w��.ӱ�LVE�л{�V����v<�R�c��m�|�46a�˦�3~��W`}²�Q�]�Y.{�����JM��/Q�ި��L'kC�����[�7L�;j���#}y7���З���(�Χ���]�1i��v�F�>���^�x��x��yH�,�z�W4��G{�Oa��D/o��;C�F���ICۦ�\�{T�/3���ojx��7�B`�oj��V�s�w�+���w<X�ʖ����N��tX%E�cF�~6����=�V�����Ǿ��}��&9�ˏK���O�-�ݷ(���I���sR����#�S�/:�CT}Y��zf3����N{�N�Sˮd�hf���7��m�f=�{���܆8��p���ꯪ�ұ�.����Ĳ�svCz�u�
*�ç�ΡX箴P�ӈ<�~w���v[�ɽ���8毞��6���wl-��)����@c+gA��5V�E���,Mp�\��Z:U����W�;��[�:ʼ��W'Zv_^^R�e��\�O��.w|�*�㴟uCy�/Q�YO�s�;�x�O,�����8���`������ .̿��M�,�rd�|�����Oe-5=#F�B���Evф��+s.y�ª�g -�me�h�U��B{ʥ�g���������
���ȶ�Wa�R�hYvꋓeJǩ\�u?��St2�&)�x��
@����`��j2�%S�YQ���zk�gc��8��N�䬻�Ӊ�z!)n� �����v��|e{�y~^�ZTIAw8��ux��^�X�;���Z9��{s.~{me��e<�s�P�r"�N(e�|�Ee�H0���U����q�T�L�[��uWL�Tup\��#Z��4qS�N��+��M7Yq=��{}�����9B�X��;(fTg-%Գ�UЛ�X�(������c�1�ǝ7n�t�IN�Os\�Y��}D|�P���'�uGE��uW`�Y��Uy9P1=:�k�Ef�.��%�F�4�_[��Se��K1�*���v�8���K�{k���½��o8�S�����{�&����V�K~m�����׮YX�xD����3��(�^���O��Q|�[x�9W��6��wCr%Bi�j�9����fSҵ\NW1�W|1�m>����k��� �aa5WMl�{�}֧W=�C$��~��[:����or!�5��}J�yV�Y]
:��ie'���l�q����K��Wдt�z� &��c��/:6�	J��3�y�j��fO$(w8����\�@K�}���8ɐ1�St�ﴧ��0�/u{���a�3�+�Y�a)����]��y#f�6n���7�FT�|c��}��w���]��4��]y9��<�v)�*fZ iVp=���u.sJ�����tBC㡬�%p�>��ި5^˄���.oԭ�x�wq7x��O[�QM�}�V���5Σ��ytK��P״y�ڢsml��#��Z�gJL��ȥ��,p�;�j���!��Z�GvF�����}�r��of�eߵ�ۄ����i¶�Ak!_���"� ���Or&���x��3����3���q<͎+*9Pʄ�;C낮| En�+�䝾�|����y����\�W��sڎ�a�!L6��<����Unմ��J�)MFX0:��Ϣ�^=�ՠ�Չ�Wl���3�gY��mg'�{v�EؽU<�X�_�Ye��n��Db��9ٙ�ڇ����\�8���VV;�u����;f����@nT�G�\�So��qt&��G^��V�q�3�Te�a�����}}5��X̢�������ɘ���Cʜ`O]�B�^���ζ����R��u�P��/�ے��*]�>y���D�rï�����8�7$�Q�2���}{C�����s����bS�� ���jT�Z�<���N�<獿yI�u��ͽ�U��dl�.t�f6��AQ�=,dƇu�4dU�à!����𞜭;Z:�ˉ枭������Y��ʄ�L��x�0r��4r�S:���� �ڗm<�r{�:��I��.�����X��Ow��xڃ7�n��$�|y�e�?�����8S��[�Ē��Y=����)�vN��㕞t������+���&�ۀt~��o<�J���>ʷ�̧�!(��ȗ0�
���g�3�t꯵�]{ك\;�I�z�_��&�%q�*�BS�ͼ� ���+�:=��!7'��~�G�%zD��
��T�O)f7w�IlVD�Q�2��ƫ�e}����������/�u��z�;C���d@S�U:���V��Bf�`.������?Jܚ�O����i��ݓ�������JF+Yۍ\Kc�jĬ���O�,s]�xT�N�s���Q?j�īRBg!U�C�S.m1�pWh����*�g-��:cbr�d��ukc�,O;��۸�q5�'y�S��2��
��ώ'�w�f��z4�os�����}���1X�[�i_h�p�^����[�����#%����K�fn���1��X�>�yu�"��9ӵ�ނ�BJ��b����qR�Yfhz���2`���nZܒ{�QT�v'��h�$t�̮���y��\��7����iQ8���Q��e=]��*����}0�St�22�N��d������}�ͮ{�/�T�Aj��]E��c�w�7�޴�D'��S�:u�O	\N7�\�RC�F�����.�.qT[�]G��(���G��Zs�Pk�r���<�%N��\߉������'��_Y�n9tU�`Jx�&���ܞ�]�v�Ѻ����M,��7� ��\6�T�֪"�&-u���9�մ�ݝp{��5|�k����MvMƨ]_d��F��ǩ��{ѯ�u��ǧv���z���w	󡯲և�ی���4-�
PqT�MIӲ:n4��n�[�o8�E���Z:a[٨i�q�;���1�w�����xHO���#8�0�WK��N�zAs�Z:RĪ�/����G5��"��:��7��z���eq���U����%5�!k��/�t�R��C��ܿ�n���=S�95Lf!��y
�-؟�J<,�ڃ	�W+s.y�跐m^Z}r�@�;�)�lF�Fe��nE����	�Y���cveL�m#%���*�3��>�k4k��t=u�m
�T/�֗�q��l����}��F�^����s$�:&��أc�Y��j��;z�m>�%�7z����nԉC���[�Y9��k�ZFsQV7��l��ԁ��btL�9o.�;|�ۧ<�魫ʘ�Z��-��}�6��G��b�w�b����=�.�U�)GC�E��3�>ՙ�)�}ڨ�LV�#ʳ��Z6.�┢u��ޮ.X��If�4-��fƠ����ϒK�J��b�lL]+��-Z,Ǣ�����u�Ѣ�!#�{x锸���������v ����CN�XU^]�U�ćH�8-����z�����o3�Qoe�@h�=wcA���D��`o)��e<�T�|��6�7���wUL4�z;(��_�fH��W���O.ZQF��o(��v��3o������[K��]M�}��V���9f�sy���tk����B�Y�5����wCW��P�tT^��/�1#�f�U�-��x���l����A��֣NmeM]�off�?�)ie�j8����κ�QKAM���������í�DE�h��_qf��ޮdbZQUOix�,4�� |�rj��E���h̫CXosiѮξ4_zP�rDܗ9��+�{�և�O���q����A�^?�hn>ސ��%MN-�4��{;rc!������Z�HޖU�35�b���e�J���je%b%,�'u@°����R#xt]v���Nnnf��'�r<��Na�����T�VT����]������u� �HG������:��A�x6N�������M�#���R�%����D�r��n���v������o7���՝j(%�����j���G�fQ7��NMڢh�<P���}wJ����RUx���\�J�
&�IX�<Ǽ6�Y��9�ښ�d\�ΠP ���;�2����`)%jT��.�q�;�٬8�P\<�M3��ٛ�����ˋ���T�a�V�b�i'��ŋ�ZF��V�:keGB�o[��=��5��K��u%8G�ٵ�\��i�CN$/~��uw��-�u�}}X
.q裖����RQ��ɴtoWhR�<x)A��j�waζ8-R�Li`�h�*
/j Goe�������rW��*���N+�eu�	���w,�d@���B)�<��.�k��:XL�E{[�T�2��4�^9���WQ8u�$2�`Wf�\���V�2���(��x#xMWfT���+t����O#Ѫ�ٰ����D����`����/E!������WW���{Q�+��Vfs�w�XTp���J�սPn�aꜲoe��j�����2�n���C�؏4�Xʘz�1�h�"�Z�ui�;J�X�7{y|R��r7;���]�B�I �(P!-a֤Ta��P6�P��e�fR�P��J4�j�kb�-*$z�p�B��ʸY&�a�	���L����H�de�.FE�5
�PwwK�DQ�R�515D�VhX�*�(!FQRl�U%�s�'B.���HQ�S
NRfSZ�4�r�:b$�<�ܩfD�\�ڨT�R���,������,Z�)HfHI*t�J�2�#�!�D�fPh�YZ� e�4��%�йTHr�!t�K]G3hi�(���Y����H��3(��=\�f�3L�"$�$�)5.�MPD�VeUVZ�.�\*���;HT�f�ATY&VVT�J�s@��Ӊ���ן>޼���c�꼡]��f+��m�����Mv�Ƒ�=Y$R�m+�%eoJ��J!����G�Y�7����wl[t�m��W�}mb�QO77������J�L��tsu���vQ������I��Ԭ3�Q�����]=�^W*I1Tڇ�T8R��������|��i�;�B)g,y��zg1ڝG*���m�;���\o��l�@�^r|� �7�Q��Ux����;��]%���a�D�]g&���1M���k�l��[Aq>}>+��0_S3z�q-i&��}&����z1���v��"�i�eu�ʂ��UF��ͨ����8���Κ�*�?�{�U�,��]P���=��C/>*ƞy��!�����`gAU�)[��ak�ꬸ\ا����n־������m�>/_j��9��W��'೟T�n���{�Rhά��>W�l̚&���n��ԯ��<��uD��Wer�-�n��]���R�]80��/�V,yJ�=]��7z����+��%���.��eN^�vmu����[��QM[���p�(U��՚9���Pz���r����"����B�!��h�R��+uݟ�<�.�BU׬k����ʒ�`���Oiv>�v㜏 �EQ��⻱]Z)���}�f�V�8�>��n<���׫��?�Y�/h��i�?+z�M*��g3x'�
N�q���9O����S��J��2�_Z熹�.(&+��\�uk>��3�RȺӎ�c����4ܲ�K4�S�t������]W��^ai�yY��7qڏS���E慐��P.��K7��:�fKz�+_9�0?��e�K2�����=N�<L�Q�݉�R��/&�	.'�+5�R󟌱�H�~]���rq�~�������Н���J̑����9�� y���Q������}��y��:�r;���9$�S�ײ����f��x@ug�nT�Qy��/�ڴ��>�,x�oZ��~����O|��u��g�3�X2��|�ൕq�_��P����rͯmsY���8�M�s��C;緳M�ʈh��Ū�ql���>r�w<����2%�;v_]�N�f�ۏX9Mugb�_�x���u��<�ض,[W�v�[��]�N�yQ�m�{՞��Eq�@^����]ٝʵfm�4]3��"T>c�uu%Ϯ�'z�8pw����N�sݭ�vޠ����M���$�4^|��]D̨+�l4��Cd5�o����f�k��ۯ]]_�2r�f�;�Td��b�e����4{�䴩0�m߶�����bF.ꓨʧ�g;"�:��:��9�O�ϕ��wۙ]�ym�m6j��F��{��|f���׎�}�~>��ƅBm��qUyO�y�+72�8�]_n+�댃���PgZ���\-��>hѼ��]0�s<��O��|��b�Af�='c]J�I��I����m�AᓈΜ�v�s��:ﻜ$�n>�k9�77�t�_%�27�3�6z�&)wU�_'�W݁�Ֆ�t��I�q�_��&)�W�*���O�oAU�������gܝ���v;ZӾ�nuu�����-�4�|*ymn+Ǽ�Y�ڈ1�b���/
��	����;�̴;x�mۙ��r��OFo7��Y�+�Bܦ����8+Q��.��,?x��@�}�²��U�g:���$�^ �5���ұ7������Q�0u��V䷜�.�y#F�H�������j�=R� �7���Źh��%�8�е���"0�;�3�]ˍ7K&�I�n�3�s�}�|������N������-d+wbb�*�4���u<7����;���������]6�Oٌ�7�PӇ֦\*�c��+��.���'�cO���A�l7]�y��������+�pԕP�Aڈo)�V.��uv
q-�&��Ggkg�9��=I&P*�x�����Bs���n����/T�LLdӡ$����ޠ^7���M}��j�R��Քf���w�K�%�X�D�T�c�7�5t.f����3(����J���ogqF*�ӕ��C�\K��2���z��
w�w5\�*�ڻ��V6���R��㯭�$F�]��s�y\�+H*����z�����s���u��x.���Z҄g"�=�x���9��aWvㇽr��r�5����ñ���k�ꋃ���x��ۜ��a���T�������,��|㚾zm�oQ������V��R��^f��X���zZ��u���:��vJ����ã�bS�eoQL)����҉��Ë�&Naq%�+#�yf���Iq��y�ɹ��ܓ��C{@�y6�<׏"��y�6=G*��N�5�:v���Z;��U�$�Ȩ��%o$]��ܒ������罋e�/�}_T�V���b�ܖ>�����ו,q�#1��m���ٜ�\�uZ��/�
��2��}Y�]�y��2f�zJ��D�娹�yn䑹�n�#Pܲ�C[F�6����ˎ)��|���	���k��k#���1�o�
�S�b��B����'�\%n\�-�� 
�Vs�|�Ս�����7\u|���I�We|ime�:˺|m`�ܿkJ��Q,�v�Ӷ�$�<j(.�-�i��J[�	+��1���V�+�R�<�.V2��oܨ:�!T6��;�K
�Nm�[���f��+�#@q��/r��;�[���נ�m����jO F
3�j5<�����}�~��y6jf�
�.:|�~��oԻ�m��>�;��~C_������^��;5%��^w*����m�h��Q��.V7/7L e�m�Ź�l�^�W��x��ZV�6ᆰ�������mn=�ƽ3��Ol[�YX�\{���x��]k*hwm�T�j���H	�=hn�e��Gi��|���]A��F��@uK{�k;9Pۜ����t)���F_X���^�Իr�yE����r���_5}4��X̨*���<��;������|a�5�Z��ع�V�|u�Z��D<O�!^�t�~}���t�(7�t���u��,��;I�
E����q����W�T�5��kq����ac�&`;�t��|7�Py�άr�\��N߇��m���;���J+;C�)WwbH�̺Xg
�B�����A�K�_5�Gt+z�A��Mz��y[�jt(j�cW|�H�u�C�)�r�I�ٗ#���ˬ�����m�Q���*����7�z����,�)�1Q���	eA��"�e�Z�Y�Fm���˧e��S��MAz�:����bb���L�d���
���\���*ľW�f_����eL�>L�Q�М�D�I���I�Z��+J@v�,pk����ɬOv���"�'N�P�t���_�k���L{�y�N�i���zju9�<V]n�6����ɯ��;K���>[�	���Y��;�>�pɋW=���^v&2mIw��zp�|�V$to:�I������<�qc=Ћ8��=�]�����Y�!�@�-f:n�K��)����V���_[3���zv�j���wّw!����	��>�4���:�ޙ�1c��7���b��^��\fbT��y�5�R� +�:�
ܣ\��E��ՠ���Y�k����E���x�`�����:��/�,�-ewQ~�aA��x��䭷�]f5��Ԕ�5i�Pb���S�����_Bw�𬆀̨��K�L������Ig	��=^��8���z��g}��yK���>����7�h�7h[Ҹ��<�w�w9�Z���b����n�F*�O;��l_7|�>��ip��T"�hY�'�������S�&�߇{Y�39U�ی)��s]���M^�w�{�<��Ȗ��f�k�W"��t�k:�?uE�J�m&>�| 8�k�<�쪶��-�7��Zⓕu{�#�T�=�"T�&%ʛ�[WS���ʑ���R5�o2��o��ic��o�|曾65uݕn���q�[yc7�0��X6R�FQ��Ԝ���w�Hf2@��:�w4�P���I���Q"v�k��-b�}���2�"�W=�� ��(�Sws�a�(/�������}����&w��Î�˱���D-I��}���$AKY�.5�9ҷvĺ��^��՞��}�_$ҽNys+�r��m	u<�VЋ�;�s���r�����f}v;�Z�Cĥ�]��q�1�4����Fm?�-/{�r�}u��:��G<��bV���/zS�����ִ�r��5�`��>oμm�<8�����ɬOv���#b�Y�OtO;CHN7�t5z
��n����
��4o=*�o�I����&����=,f�y��L��S
���첻k�K��uаev�/�Y�љ�s���W+�mIOT��b��6�V@��ʅ̻��gp*q�(�N ��-՛�l���M��և�a�9]S��`����	q���xq�E�U���(���'��L\Bx�Kd���ˆ��^+o9�,�ސ��j����8��qv�|�WR����Y��]V�ְU�m�EV6���7X)��VY���O/�]GW��]+�ދ8��:���T���l@�����2�EsFS��`���p&������k���j�o������Y:����sB�,�=B�3���s�`w��6�������9p���*ƞy��+̻�V�[�+;)����n;������}��{��f���]�-ueL�C(*e�ݶ���7��9�ki;<��5|�k��Ԧ�o�x���B�����eg�G����>����Fw���j�eO�Sk-��mf��o�R�� �����"�}s�]RccQ�C毡h�V������h�X���tT*��J��[�j��7l؛WReZ�6�ٟ\�������}�A�k�$#3}x��9f��8�֡t�4��P��F�W�����C���޶z�= ��w7��U���s����n�[���W`�s���=�n�����6�\���1�W)6�U8�p]¨|~�� ��읜 �ʱ��*�i1��v+����?_'��*P���=�@��$�+���ОRQ���Ɯ�+�o���"]��,Ŏ�.;���Ip����Ҙi^12�����
{�\�tM������W�bn�w�5M���9k{R�1���G'w,A��ԇ��[� F�����Ԥ%��'v'kI�������J0��u�^���ͭ�WFs���c1��V��Bb��ݨ��귦c-����*-
��ӻs;��k�b�r�<�i�pJ����2��w�^z����쪓}닃�B����⚤�6F��7o;�w�l�]��-R��*��-=1�س��&����[�^��Y�=,�Rt3q��(��샊��M8�żWOW����ꭊ��F��͊yko��i����Q�3+�OL��m
�Ռ���\T�X���ak��\ئ�>܆�����Xͨq���<�cJ��!<2�q=Z�O���VuUD,k-��㷢���R�0��5<��T1)|�n�y��zN����ڔަ7�Y�l�����=9l��y�T�#:ƅ���ю����c/�����{�*n�>{��x�me�����m�<�n���a+�	H�����@.��@��qq 'VY�lfA:�Z"���p�Y� �!Jy+�-ǖ�=��EYZ��:�i���;pn�R�-Բ����? ����)�l�ݽ�܊$��gd���v�z��@��W��UgP���똮	� \�"�E�uf�dm�m�ow�d�Ɯ���5���e��)3���ͰV0Q�ags�����%b�|�S}�9����cr�;d�����v�,��������s��S2�ٴ�/;�ɬ�RP٤���7�(,���wQv��m.�ا�S�E��NaH$
p'��I�y71b=k��ʳ��y-�7��;N%�E��cVMb���8�^x�C���X4�:3�Cir�m�������h����\�F�{�dw����"�N�SQ���F��80�D��l��)\w.��]H-���w�����Z��WoR�sj�$� !����్��3Xʕ?�ś/+(TvrΘ�����	z�rk�gf�=gZ���i�7S5�t�n��.�����q�����Ce�|cv$A��Π�p\n�h���fZ|���:Wmĺ�6o��������@k�uՕN�x���R�&�]��R��Kc </)M����-�F����i��%s�v�"�N�8]�ZOו'bxs�a��#jkg�J�c��X��wF�VmM׸�WVe쳜���R���ju�㽈iT�5N32��uj)�r����Y�록�}2�*����D�<��z/̹��f;�Bxfs��J��B_|z�v��֞���nk����Q#Ts����2d4��i/�^sJ�5�#98�n�=���E�L^�+qE8=��gl�TY�����Q�vV��f�4tm={�j=���V-=2�bD�[}y�6�s��:��sx9"�|��`|XYdwP���ժ�K;��@�ëR�M���4�-��i������2���ޏ�'�.l��"��a�AHR�̇�+��K�2�\�8i[����K@;R���,����w�1���n�r����	��L�B�4�ˎWV�0�=�����t�������.6�+�+��BՎ��䚭���V�[Łg6�5��q�=c�N�b���X��+���y�ج���;];�GM�ۮ8��@�8�/��͛�m-����Ρ���m-��ǰ(R��4�P=i��9�#���_o]}ЊzLͭ�DW.��By��)��g0!��>+2gv����yv���`�ĶY��e��-���H���O���S�V�q�g�]��&JP �fj�5�-�cv�ܭ4.�]3�AvN�U���P�T�����³�#F�t��Lm!������iS}��ý��W|1]�2��y��D��_mi��뼚䖶Z�Q�J���<w��z��:�Ic�B����v�BCY��.Ų�ƲTrv�sI�{|:��^k�/o�R!�-�6r����<�k����jʺ�>�x��Ns���:�!Sg(P��B#��D��&Q&�d�+��vEh�Dʌ�!*Ek�ҭT��IQ�E2��K�DE��:-*db�eR"Hg0�ӉJ�T��#3��\0�̴)$��LebÐ�ISX�UT�4���E
()5+Q#i�"J0+!"���2V�@U��*N��HҥJ,+��Y����ʢ#8�

.hG
.\1g2
�K�e�d�\#P�e&���$��r.�k(�-QCZAV�J�b��f�dU �H���Ԕ0�I(�$��!f"EEX�4*�����(���*��]9e���2�r����^�ʊ��3�Y�Z�	!č�{���׺�v�a��J��R��O+����H]�暾�Y�5\OR�}&EvnfTyMK$����*&���!U�jt�J:f��;�����M+��ٿw������#d�:M�+�B[F��<��cPqչƎjwl��C5���P�)��Sw��!��n�R�GS���p��R)nޠϥz�S��Q���G�m��Oo���)[��b�Gj��NRM.��q���좶b�2�&�1=ێ71��$��p�b�6�p��r��m��q.&>N����P_eA���OE�s_w-��.�o�ݎ�:���s�a/���jȃR�-a�뢷*s��Vޡ&vw�+�e.Q#tV`.3�����K�z2a��B�~	e����f.�GD����`�#�@�jbr�n�����t���К?5�4�����(ň��/5�8�N���l�}�A�QYɊ�\�6��}}"����apx�9�����b���tQ�~���+|���v�����{��H�@\����饙�&vPlI{V�WE]��U���SQ�.�h�n�@*+UÞL�D���vQ;������
_hThf�ks�4�e��Sޡ̪�,�u=��#"4pn���@d�憇d�o��V���hz�Ej�����*G|"�d�Z�S��Tx�OJ*w�-��������)�]T7�S5�2X���>��p�Ǐf�����sor)u��ou�A邸IP~�}Qgy�&)�Ŵ;MH��ǘ����Ѻ�j���.�v���`���z����k:�h=����u�T�f�t�=����\d�I�PO5k��p����ul.�Dє�����n<����7�OLf��o���l���I�q�;��qm�O+���Sy�e���ξR��窺f\�&����ӵ��{�{Ņ���V�P��g�/�'�v�}�lqz!o�\ek�]w�4��Q��U#(�����#כ������������hG�9�SV�'wh°�NM�g9�λ�y��N-�p������y
݀bS*\������4��+V����a.-oS�ʆRLU|ڇȽ
����GGnw�y]���n}u�V�7����B1�ٌ��\�}V����Ʊ��\1�;`��s�%���*��
w�Jњ��2����Ԡ�Q<�3x]ڵ��WR��V�a�åa��ǲ3Ձnȷ��-K�Ey��5$F��]UI�#1���N�S����ۃ��R�7�nr�`�I�K�ikTS�k7W{V�0kg��ݵ+����V.�s�[�sZ��\�X�@c����x�9�b�^^?>����\v���Qr)^UjƆ�A�nT7\k��FXT�
���7�>{�R�^�'.�'&�G}��L�گ#U�'�c��ͽ��������IX.�3�- ���gR�<q�{�>=��#��w��B��],u{��W[k0|d���O���wЩ��9+o�"κ�cT��־m4���}c���ӱ�vH�YZuwqu�D�ڨ������S��|�8�{���ᷪ�*3g5���|�m
a�9#UH�ݢ�5�Gr��4����ʮ����)mL��{��	�w��TGs��[�o�`�ޝu�����k�ǖN� Vd�B�^-|k�Hw4�Ty��n9�jv����n�q%s�W��&	O/�V��2a��u�s<�9at�Ӻ�Cݵ�t�Hz!�_n7�f�YԻ���Dխ֮�lq��;w��Q�Z�S
�T�H/��o/�����3��y�	.;��3�uw>�P<�,�N�w�k*�#M�+զ�7yysr�a�5.;PS�Nm��o�Q����G_��*�biJ<,�ڃ&sQ����eco*��*���/�ʄ��C}N����k![�Lp,�JDoL20u�VkKuE�%k��'l�E���em��mD'-8y��Cz&0�&~Qe�����Dh7��אim^gU�3����\�>d(�7C&��ӭsm��[��ۥ�LC@u��nTsv���F�b��<\�z���M��b�	g>�	���M�b���tZ���8~���0ٮ$�zf�-��y}8�f�ZϹ���ʔ�~����87i�U�f���uk���au�_G�����?(z�zk��sV��m&hq]꾺]Q��g�S�'P���^SH^�p�k��\ا����n��T�Κ%�A���Y�l}�b-�5�M�]��1.}�uN�Y� �X���b�;c;���R��RsC���Y���V�*�h���kӻ��3�b��l�����E��Rڙ8] �4Pm�L��ĺ(��,8quu%@�f��
�����"P�}��z�s�c;�=Ρ��nUꕍ^�6��e�ro�Z�j������Bq�{���PrK�5=�����Ou͚�a��~�Ϣ��NS��]��ڈS\�PX�Eŵ�~�=zg���,X�Rc�>�=��^�I2�����X���3QҺ�G)���\��+�):$���G{>�`�ޓ�;�4�T7l��B[�4���9uռ�b���s?�]�v��)����p�)�NĎ8*�9b&�w�i*�ԵÜ�Q�_���Nb���/�z9�$�\9�v!�{W���S���[7ٱ�6�2�+�������&��O�>w�GwE�{�^��o�wzx)�zԩ<]���1�5xim^t�<3��s���0����|3�R�٧{A�[P���;��	�������\���Jg:��Ll�8�kO�S}X�ZhL��s��\9�͋&gr���I'� ֯�ˤ+y�,k���3�wX��|���ZC
�9�}�W�[}��>��(%ye���ݍ��u�K� VY�1�ƺ�z��f���V���]��,j�&�G2y̬���֮U_vN��S�w��D5'��+��^g�+��߰�����J._���):��$���w�Sr�NqpƆ��3ش[*���q��[��λˆs��7vw�+Y��{��N�TM�&��i��+��.�Vnj��p��:u[۞�9S�X�.u��Oz��v���+�d��s3Y���'������Oa{7����29�y��V�8sI몾a\����cP��bzD~���iP���y���0/Pk��0罕e��[W9��u�8�j�:�@�������Mv�6�������ei��c��\�n�zW	��:���5�r�N�����;�0�۝�Z�z9�L�_�ͬ��:^�C�8�o�_�5���^�ϫnEw��:��K��9#�G���8x'���%1�1ϫ�wzxɜ=��ix�h��Z)?wCAZLU�0�WIsQ8�<<���x��P�Iߨ�4����HG3	B�R�nb}���㖟X�p	�f`:����DE��T��C��7�a+u�8�:)U�^Tqd�Ң�^q�[��K�gR�Ovs�ضv��;sK�����&��v2iП��z�.�1κ�k���2�☱1ם�@��C����H�K^�SP�n�l[�1�h�=�_�1ĭ˻J��[<:)���W�뻻q���cil�\�q�����&8T��=�zld������lD	^��ҥg�KJ/l���Y��+�p:�3��ar�����4e4��ى7��<����k�'��p\����:jJ�mA��]���� �����u;
�H��@uP^��uw�V�&}�;��䩡_}�6��hq싢{t�K���t���8;�Z+��ʾ�hw��
��>�(7t��cR<�>sgg_�������*=��B��Z.Iӷ,g�Ė.���^O���/*�=��ށ=U�nZQ����+j6�5��M���[��{#��W�zv;$�����G����6e����eS��	��2�b��������^����ZvOq���o}�Q��F[;��Q�em\������y�vY���q���뙱;��W����Q�x>��>F�o�u���+�qάYbS_!��Pf77݉���:�_\U�F�z.;@.�P�r�E��kO��zp��}���®���O5�w/�ߜi��]wA�뺚	�ۓw��W~@��� ��t�i~�mm��@�3ü�����^����/E������g�Gb��?(��Q'Ý�U�(�>&�e�{w��#�{޽�_��Cñ��g�2�z�8�/������
�%�w�j<&)�D����G#O=�o��>�Rd���޻�j���Q>�>�|���_��xZ��ˀ�����[��}�=ӎ�G����ojY�a���A���qW��֑�zB)���N���n��ޯ� �N�Z�@_�}'}��c�~�7��w������ߎA���G��<}�n�\9�*H���Y�ڪhԞ-�#u�����}��ﲰ��JgF+N���ߩ���W�=�O�9>���=�;�g:�o�ߠ��v����8\�jMr�3�&��I�:jc�c)�yVѸ�>��p��'�C�׍���Mj�~>�)�C���ov�/p�dP����#�u���
���kK��j�8\'b�+��.��O�On�ޞ��>�TY��^�"�<Ĕp�;4ͅ�q���k�o��e�l�u1�m���182�QS��} �y�ժ�6CrJ�2�g����l�+Ì�'+}r�^��2��iN��d�X+�v��f*��D[՗���]@�Fw�ٮ����w%Wֺcv����5]���a��␊wt�j� �.>.��|�+��"Oz���դ~�̿W�e�=P4�{��=���yQ�X�'�=ZǞ?X�[uk��5��R�^V��P�L�د��~�e�y�����l�CǧDO��"�:W����R��r6���<'"1ϳ����x��3��z�}�=j�j��0��]M�ء�v=]����$]�s</�5��'|{��@s^��F*��\�����?v�T�UG�y�3�T����[e��)�K�zf���鋈ɝg��p��f5������ZQ"e��f�uk<v��Ԏz;+Û��4z�xr��������Wz���)�p����Пe�z+��T��裪�Dx�_d{-����b���d9U�;�tXM߁�/�l�9�p��3]��yi�nՉ�q�y\{�6s���|^��_�}
r�. ��]��3���=Ȗ�%\lO�} q�&���|��O�Z��_�c �u�:��5�w����K�"6�&����_yQf>�]* ?d2�ml�/{]�W>�e{%9�(ͼ�V8[JQ��Ǵ����_1�x�WV�h�gkU����AMZ�7��1e��-J�D5.�lkk��c��GhD��Y10���C\���l̅��i
x�7�Jݦ��;��]Qu�J+��2X6�<a��=u-��mf�������/���[=z�9A�Qɚ��h�x�V��KyZ�����L?@-���^��LM>�i�Z;�K��#����Y��w�.)�0�/��ַ�bZA�P9�V ������x��-���d��dE>��������=5�;t_��5~�観����G'V�A�<�����Qo�Q$�,�y$%���O����B��6%_:��K����}��H�y٨�^��~O���5�q��&��//�>����om���X'��zk+#<�fO	�l�i���Ǯ!<̏y�˘Q�u<o�۸�;�g~��K/K�rz6��`����^�Qz��E�<;�;���:+M��|��*,�ǆ�V�:���~[x*���_�7%�.W����"��o��F�'�nKgnv���{��Zu�3��l
�Uo�C�K�f}3/'��t�����r���=�u�}��_���Ló�[P�3��o\���j�f:c�:�tЅy���J����O�]����Ӥ4_���\.#2J;s,a�(z��<'}.j8�y_���=�^+�l^���ӛw�����}/��ǲ�x��;�Y�8��@.exh;)���_��QQ��*�+ÂzV�Ks����⎔�zp%�R�YWٙC��s�z�itl�-l	��
��f5���*jf\Yx_�AJ۔�\.�w�����n�d��_N��s��)-K�u;O��V�U�)@�<��ޢ�LL5>�'`�1Dލ�k�c�0|��FӮ��i?G�Z
�����(�	g��.F�������|�U����+������E뵋@�̨��8LΨ%����!�����e�{�(gh�[w��(����h5�7�}S-EDh�k�MM�Yo�%�����CR��)�Bx2���zu����Ֆ�V�o��,�D��KT��8�%uok���7�JՂ��LԷ�'ҴGQ}ĵKd�d��Y�����1�#r���ՎS�7�gXUm�Jm_
wy�K�3t�;b��hp�B�#[Ϧ2l,KL�F>��u�)^�Q���@�Cz��~���]��]�n����w't��Z��*�bW���G-,k�WN��n�1�+�(^W^��A��V]�M$%Uر7�ܣg �ɍ��A۶`�GA�Nu0l!ב�|w��k��+��e1�ō[r\���S�Ϻ�����T���q��:d���86!��.۠�|�\��YuXc+wKU����%bh6�]��t�U�_N�jmV�7�_Vn����\z�f�;{]@]��QH��Y�����.�0�X�kwi^�u75�_7}ڀ����!{m*�r�A�k��W
�oQ��8TB��Uf�/�T�n�|~���Ր�v�m@�9��b�2��%]q��2��N��
��`��$KI��N�\�N��M8�����/x��KR��i��(���g��j��]	��v�����t�5α�2�����$�`�f ��Ѯ�y�;�,^ )=��u����hVK�3��/1�짙 --���{��¸nP3e�p֊z������W�IV���u��V� ��������Ľ��Lw��TZ�K᫝�ѳ�����*
�bq�'���903o'j��(�u�t��r�:fPxz�ã��n6� Χ���r���{�W���LT5�,ū�h�@�Q�Yp�^7Cu��U�E�����5V�:�+M�.g��]g��+ivX�������1�iS��Dj�۩V���� ެv��x�t�f���0NY��Wa���B����QWfnӤ�Ѯ�S�EN�J�w�}�7��EJ�o2�D˖"p ���&����3��������$6�#s�����8>��y�N�C�_@�1���O1��n_K����qۜ�o+�\3�:,К���jy�oZ\oG���*�mGX��눌��A8�6MGq��W�L�Ŝ$��;y�I�ê>�6��)X�Õ�4��尧���;�e���n)���p̄������XC�Zm�����6ͪͽ����H�(�xP�@���}�p�� ���8s�9
�Ȃ$Ȋ2I%@�%����d��R��XAM�t�UJ���r��p�j\���%�U�e���U��r�NP\.�D�E�N$�r�(�$R�(NUQG.dY�9\�$�V�Up�'9h�#�TXES��\�<M���PE�ʙI�%�ݸW�339�$�(�A8kL���kMX�Hqe�I��	��$%Z-Y��r�*I5.��V�EG�B�&A��ՑDr���EX�d$Qj@f��" ��"YV%&�;�K(��$�Q$��\mRI�*�:q�d��\:�E9T�s�EH�YFEE	#�8Xl��4"�T J��.]_y��P������}�҇�_Fz�.@'����9O�4�RQ��ڪ=��� ۼs1���*%i}�qw�,�:&�姝%�V��3ε��u��CѾ���ޗ���g�q{j�z����š�F���ڡn(~�@O�S�ɼ�<��۩����쀧��Ϸ��q�z}��_�=j�='*&�hy��'���0��F���;�]
���&����T����Θ��D��D�wG9{���m/�ͷ��C���|O�*���K[ڃ����,��z���q�S�˾Z��չ7>�>�WS���E��H�z�n|󞹐5jhW�_W�����[��z����+7ڪ+��k���\{���]6-�*M�L���D�c������*�Q�����͞g=�s��wN}�i�o£��y]���Ӭ�Iw .���5���RI��X�z�Ñ�P�{��Wk���D:�zdTk����cS�Q��x���|�y��I����^�ryL��;�刏i4ϢO3�7P��fއq���j;�p3�Ǻ�'��>����	�6���߫���y�«S���vQ? U��/���B��V�q��7ޞj/m�)+�����>F���1�l�k"���*�/�:��s�V+�է|X�oK�V���l�������^�T^����2���Y����oWK�o5
.ȁ����i�c������=�|6��N2�a�W�u�=�y����t�Pfv���;���xvt��=.l����o��6o�~ͭ�$��Z8ra���T;ͪӡ���wj*o�lU��N����^������h�����ݝt�N�d�;q2�x�챗���`���Of�����Z�)���x�)c�W��߶q����7x�*�ݤA���+���]�&�'D��˷���3��3�b�7�����l5>������д}����-��G�ܳ�}o^w+ԡ�i��~��1s��a:�*+n�y��<�>gF}���������9��\I�Mu�{ݹڬb�:�'a�W���5'�T�Sb���9�2�mT?Yu��fO~N��~4������ʌM{�l���(�CU�����9��'��\MCܢv0������@V
��k��zVbQ�~��Õ6w�|;To��_��!NQe�!��x��4(�H{�Cr���������$5�;ޏ%�Y��j9�R*�C�3���^�s.O�sq0Xs~�a��㇖�޳]>AV��G�>��g��Zs>]^���Q^������%�zF�y�*�S��r�9�}��g-1����2�9��)VH��~���y��I���EvٖÎ�%Z;��~t���;M���,[�P�ul�m0����{"�d�ff_:����5X鑔+N	��E�ͽ|�S}K��V��\���maa������o0������l�`��E�&~�=��i�F^�����?L����/�7�Z��bb{�����sXw�Gz�7��nKgML>���14�mg�u	cBud��W�����)�����C|�'l�j�};8�� ����>GML>ܭ�
�=]&��>���Á��)T���g%߽�i�,�p�o��������>�Dk�(�,vl��sra�f׸�M��>�':�(�J:^�3�˅�������Qϼ�����=��>@�o�e���e���o�.&Pˏj��&���3�o�ݪ�pv|L�1j���Nk|Q2����W~Tp�#�wMռ䢷,�/z��Ez����f�
�o�o��:Xq�灿mc<�;��<�\W�n��&�P�Y���ށ�Z��1�����^�|/c&��q�;�z�v�{0r>�#�����^w����K��~���8v���R���1Y;�~.���{�G	��F3$�����@�������E��wz��l{+î]��>��R"6D����Sq5	��ÿ��\%Q�$;��y��a9P->�[���o�9�����uj���*�]5+��!ee0���;J/��|�������t��e�ۑjpշ�P�Zpm�H��+V�h!:W\��tWW vc�s��t�{+c�|)݇w;�
5���r��es�tO?&��u��T���W����_��L��e��n�[��3��%W�g@�M�`!#�k�TzbgN��.}���·c/��>�6yq����q쀽M��H�\s���7�_�B���ρ�}���>N/8�HԳq!��ש]
��̛�c���!/�+�W��1��ߎ��t�_��;����I��=Օ܈O�����L'_E��D��#e���>���g�y<T���Wz�\��n��_�NE�x^�̂*/������10�WH����� 5�����z[<:tq"��v�>�}ղ�ώ�0V|���=��+�׍�r&Z=s >7�b_NQ��wr;�d���.b{���>���r݅�H��)q�/�� �����Y��QD�Dς��͆;6HHl1�R��%\��ƴ5̟a\U#�)И���l�{΀�.n�=��&��;�L�."���VW{�˯��y����̜�#8^'���\'ۻ~�>��8�{n���'-���x�A>y���֣��^$g���6�~���Zo\�j���%~��ȏ:׈���}I)�]�'@Ć~,��5�f�-��+�����M}n���x<I͹טAƴ��̹`Xm�͝�G)�wέ=�Au�6�v,[]-br��j�ڑ\o�՗�P�����tnZ�(�,9��Ұ�F:6��rKN�= e�屃���aW��6�LrCܹp��^�q��{�؈J�>Gn"v���W��q�Zo�� o�:����H(3�{,�m�v{V�N�>�]Lu�8_����`��q%��f�&Fz�β17J��k|���ZS�0���7���^��y��<�R�Q�X�ӱEWخ���Nv�܊�{u�H�P��v}�Q��U׫�W���~>]ˍ�p���9�(��'����#��)%����Q��2e)���O�>����z}��W���V�79�SJG�ڥLU�_bY�V������T���y�M�ٷ�R=q���VJ�3�>�9Zo�o��削u�o׻ηs��=��Ag��&t���]��+���[(�¼^�Ϭ���}��lb�?�e�[}~���cҊݐ1:wyNx�<������F*
�,9�}��
MG�8�[~�͎�%�ޞ41Ҧ����/#�����쑐嚏_��)w 6k�SB���:�33I��Ԑ�m�����n����G�x�޽ ;��e�Vꜩ9,.70X�E����� �U����V�֫�{�,�w��z�\�$�>�D�tmeĪ��b���N|U�ˤ�M*�ĎfvN�v���;���|�"K��>�Y��7��ԃxwk[��uub�F�9���E݊�^�+�y���[I�ʸ����������Ok;&��T������T�{�@��j������O�Y��>���tI�|J<����T�m$��uG�$�D�0����i��;���p�������/�t<�>u9�m{�r��X��¥VN��}}(�i�>G�&���.φ�Z�A��]�{�>����h��9���}�E�s���^'
��+�/���^���0�g�z;���}���UR���Ȓ��9��3��T�GuT�'!�#�#�˱B���Z<�<o�e��f���uC��j��_�`��¿6��C�ǳ�&e��ԧ���|-�+����d��2�x�=e@[��
�Y�M~DOt7h���ާf��7�5>�׫��o�8�v��\$o�<W��<{�Y$n��67�/ٓ���v�X�s�k�X:�ɭ+	�1��	������^�q�v<W7OG���GO���[c��ý����8O���*p��`O�=����T_�#jPw<������:�=_a��R�F�X���3���^�}�}q��e�Y�2�EN�Sb���7Sson��9�><z�d�u��1V~�V��p�q��v��ҬW�b�t(Vj
����(88o^����mE�W�f���|ĵH�6�I3��2/�WNx�[e^�U'��!�p�A�|0-n���yz��m";bz�Yb�.��pԹm�5�Q�!W��6Pӳ��&�V~���-��X�Pc��w�C���o�P�Sr��+��;��1uU�2e��T�z)8(�!$�=�ґ����wdk�4S���+>�Tvnk�t���M=W�g=y��/��>���ﺠ��%qW�ZG>�zB)��~�r.=�Ix��GS����>޴�F._{C��P��L���u?�{����+����(�{�4���Y7�Tpn �xz�������p�;�&�Ց4�t�;�e���l,�U+��|}��3��D�]羵�����g]���k�Q9Z<ja��W��jv��k�q�FX�\�	��oH��9w���o���g�F�P���@8�Q\y�S�#����J3��kK���>HH�+|k<U��𧙾�c�fئ/Ψ�~�<����ϋ�DTy�(������7&����c�uF�S��3��d��G�k�o2�uS��;���UEk�8k�IG	aa����Ng[��:��zU��+��kG_�;[7�i~=&�3��Q�����e���׻:���:T}���:أjI�gyJ�B͐]�gh��M
�J���Iո�v�BUvұD�e}cM��`����z�f�WB7=l;M@�"��ޭ0��{�hv>��]�ۼ�H�*$AOS\��k�vkz��H�Аǜ��Q�G[�$Q�V�O��[�Ab��%%�
��Ň"kE1\�Zxc߬s���t3�Z��	l�V�0��!V}��Y�3���;#��y6�{��;T��sZ�v_F:��^��ڰez3�vV���'t��>S,Zɭ,\d��� c�k�c�U{Č/�ۀ{�.�_-��8]#�������Z�Q��%"C�j�}���&u�N�Bm�=٦7�-��4�n�럖���������x��rǪ�1X(r��=5%���j�w����yz����VX���aWyq�o]Ǚȕ�q��w��w�2��/Ã�T�B���c�%W�x��Gs�M�d�S���1E.��*끼���|}�~W�^�ίH�|w���J�x\)�,�������qX�S��r��xG�} b�R2
����c��>�C�|*�[f;Ч�q��6>�^{
M��*��put]��q���x~4x[�J��z����%[�>����(uD��xwbo�^#4~�[���~�������۸�nY�V �*�baz��D��O��r	h��#Lx�&o��k��K�BR�5Ζ:T�>��i��=��� ���x�>�h��2�W�1?S��=��=��-�`m�BFl䜠I��osiou�_ �<f�1t�˱wR�p����o$�w"����~x�T>����w���*�z�/5/[鳸�}/J�2��%����C9��l�z��e����E�Ƕ����!�,~He��5M�{���3�>t��� ��,��~�����l1�~��'�u5��յ�ױ9�|F���Rj4��Q����Tm�?Y��9�T:˸��I���Ľ�EM��D��^�ͩ~e{�h��Fmh�fp��eB�~7�y��[��1��t���+�ķ[�ŕo��F����$~g:'k����Y��S��q���=p߽�Nߜ�|f��9\�"��şweX���<�=���-;0�c+�X�͚�z���[~/(ĥ7�k�����ҫ=[�JH{���G���J9�
�,�nK��U}�����^5fQ��Q�o0H۾��z���t#n1��K�~;�����#�-Z)@��g�	�}��[�%p�ܿ(�eW5���V�Fx��ƽ~�o�����\o��ǜ7�l�+>�U"�i�t�<��[Y�y܆r�1 ׾�@M�\+ɕ��ϟ]?ߪ�(}�����d�7
�\j���������gd�Łx�� ��OH�|EO/I��A�p��G��և�3�=
{M��G'N��(����ɐ3���(-�B����ccl��º��U��Ι
�7�['�˩z6Q}Ջx�#�*�-�#m�D���v
�SQ�����t��Y�v2�K�9t��Ꙙ+�s ��r[eb���}��۾�B;��W;�St�:���U�Piwm�H⼿[>�q���(��%ѯ�H�*�F�l�o
�ȇ�B���B� �_'{���ĳ�{���S���'޿d1�٨�7 t��Q���K��yu6��������Ͱ�m�ׯ��~�RG>���/#}`h�S���L�;L�ٯ�M:`k�0z�����s�]�>�L�{���_{�\U�k=g>^�@�	���&)�9Rr&X|q����݇��`���6��K�`wrD��s�
gt�B�zm�
���y]����>�]�����7C=bj��3��$�h��3gn&��TC��V����ϡt���\u�����?X�"=��U�	������)̿(�g+	���>�q}�\�CW��]��t�gA�]lzӫ'��{z�c�����w{����^ЯG�]	�^ɡ�(�+�	Xn$�:va{�����ͯq���2�Oo��q�^W�+)z��y���L�)/�B��n`��<��<��9s-���v�Ḍ�T?{����O��
���7[�[�g���ζ ����NC��(��=��m��N���c<g��7чy�A����5�-��Q��x.'Q�6��(���:�z�g
U�Ê�ĩ>��V`u!��g�4��
�Y.�S���92f	�;�Zܥ.����涴�-n�����tE��x5�s{�-_`(]�Of�!�$
��Yu�,+��z�����T��Ӂ��p��\��k�A7M�X����l���lU&��vr��$Ƴ�:�ot^p���z��\{���6�d�pD�J$��/�(j��͠bPn����#Q�RT.�L���<� W���8k}���#�Y�T�I`��O_j���h�<=��95I���X�I]�NM���L�-HjgL����Ȱ� i���K:�ُ����(��
���B1���gX��.�ۮ=|����*|W ����:�����Xưܐ��y��f\<%���M��v���(����&R� �)��H��k����n5p��F������|�m����7�w��W8��.�7w|�KɆ�Sֱw�X&J0d�w�v�٢>��4)�f�p�oC-��g����	��6Ov�k2	YEBZ�����z�G1�n������.>�o3v���t��1��U&c	���ܗ*^�jά��_-�볻bU��ؕ���,�m<s!`���ݾ�4;{x}u��4����'z��ԗnwN�
	�;ᲅH0�eԄ��QVjNڽ���%���v�s����:�r�4 E���m�b�ˤ��"��g��,,�g|��f�R�E��֕ y�f��g뤼l��6�Y5h��+�K�j� Z�sϱ����R�Q5Lҁn��ON;�f��?^���ެG�	�s��CR�5"cj<ڻ��� �U��6��=��A����{����A���7���s{g�C����#����[)�r�v�p�l!��en՜{ǹ]�wx��1�ָ6����Ԋv[�l�]�k�B��^��[��n�ӎ�-�s�m�{��݆��p�Ԝs�pPG�{�]��T��{�]�p	��E^K�Ϣ�t�T�����@]I}�_c�<�\n_dzS���u(Ρ�"���t3����f���AS3%|��XuGXx�`�(��9۔�y�39%��A�ǖAM{�o�S��cT�����˃s/oY��%+��Cmۧh}"Ģ�7���N��o�kv�5aͬzƎg^�a:N�IKg]�u !e-2��J�o0�=r�k8�����f�)�	���uec�K�w7&_d{���p'��@�������$� �4�4(q>k�:I2����-1����SÐ���U/�V&�m�	��h�9���64u�iktx�k_׼ 9�=�F|8�w�q}���Y�w9��
���RE�V����Vgd��D$�֑F-dR���;�r���РкW�s�G�PP����s��۝/[N���t�(���,�@�%�DNM9N���UA��D�*�K]܂��U*U:	Z��TYDEr��\*.AQ9%s����S")��\�PTTR�W<��Ȋ��9��
(�mts0�Ӥ����Y'#�A�e7!8U���r�ӪӖBr�*�:L�Rs�%r���ʹvI!q&�%J�ܓ��vDY��	ЙqE�h�^�9Y�T]�K�uu܊�F�g/8��G,Ȉ��UbE˦y�B��";"�����$�l�J������ �YQWN'���:!y��EN�NJ#��DA\<$�(�G�U*�D �J���?�{��{j�4���,��>��^�T��G+m��}��uڼb���^������	N��p�-KJ�wN�<�Ot��C����_U-f��gq�������z�~&�����!��i���v����Ty���]��sUk�x�����}qT�������k���}=걹z��i��;'���_��cɼ�Q�:�^j�=R1z�=���a�R7>����7=���οN+�9��3��Y�bYA{�^mt���Dw���u��G�A<H�=*��G��6-eT/v��f��{�VW�+�wx�w�N�V{��{=��ut����!���w�Á��"Lo
q5��cs-�՞r��-9۵����,��~���|g��E}�_��!NQe�@!��x�+�����5&n��ъ(���z�@�H��.%qW�ZG>��"���D误��G�3�/V� #g�(���>���)�L��P�����Ӌ�����w�c��'8�}�<^ړ��m:�w��oS'Đ�͉��ꋤLӞ�џJӨ3�o���ʯL*����c2��5X2m����u�>���[�d�5�(��-����>&7覫h���û�7�Pz1�꼸W�em�T�ׁ��}S-���̳��E�{��;+c��W|���:�V,���,�v��������YQ��u�]�Uټ�&�u�Q��6� ��MX��Җ�mf�g;
ƗJ�T����h��N�EZF��Y
vra] �7k��
����}��.��2���En�igqʴo��=�ܝZ9|�y�ě��d_y�R�#��M�>���==$�a�Rd��=�����q>�*�t`n���uG���@y3uCË�DW���\L��pf�~���=�|�廘5y��:��D�1�������~-�ׇ�̮����w�2=��0�Q�����}Үw��W��G�S>�}(e���z�v�t1���p*3��=�mJ�)<}��w|inv��}���|�k6|��%�0��_}�ZU��V��#}7�t�:�5<�7�g�J�`q5�Ϟ�Io�V��3脱\U�����w�/�}Le}�ZX����\����X�x�{����ίW=�^g��^�ք���1f	H��ت�㊥������|�2���X�k�8�~������w��~�^g�s�]��s�z%�;X�7�MC6z�گuJ�[�r����F��E��?��dD�w�=�_N������^�(��!��Tt�����Y7�j����9L�ժ�7+Ž��~��M��=�F�_�U��62�䊏MG?�u�k@�M�aj���7��@U��<��J�t���i,ڽۭ|Vr/qI�n0�U�W���g7`��-���jJ�E0��Ҕ�Y0�g���Ԝ޺�G��э�`��ؾC����=�`ܻ�ۏ�ޭq�����;�e�x��9�z�Qr�7�Ǚ�MY�R���1pw��ȸ0�|�/w�/>G*O�v۸�|:\���"ba��' �ⰆW�������ڏ)�.�֨�����\�n]z���ѫi�;�5�{2��L�,Z=s�H����:KGt.�W>$F�~��tW�o|��]l!�S��qR�Q�V ��p@���|�2�ۙ��a\��ځ9w|͞B��a�=��x�=7	�W��_��=�̀9��,��ߨ�ng�l.��mdx1ٙig!��64?}�Dz��������;s^�Þ����U��Q&��o/Uy��wv��(��/�gC�D��+ͭþ3�l��f�KN����U.b��⧍����:u��vNzލ���J��ݝ��g�e7�/��$��;>�'t��ðu��f�i�0��#�4�ٿp��5[圞�+������G��� ��-����y��,(͚Ӭ���S
N_z����73�-��׵z䌈^�h��~YhP�}��Z�;��$�>YUN�50�O�j6qݝG�7t�y%yhd���a�t��ꋅ�v�J�šOm�[���T�RhA�:qmm,����ܬ�/\GWl��|�;��?nr��d��ۘ �|֖7��Y7��Q%��Gm��mܼ(-/��C������g�w�*�Ӈ�gH���[��/W���Nx��z�W���^J
#0JKzw��<�7}/�g�Cfp�HW�P��L���	��wq��^�q���.7��c��QT��f[$��靭~�O��A�_�^o�Ǯ2e9�}R�Ozh?D�[���_��/�z0��}f����sݪƯC�'a�����늦�S��o%ͽ�������
|Ό��7�|g*I���J�U:�2�>����U���\�c\%��9\EW��-�N����x3ylL;~�ǥn����P��v�C^�l�;����ǂ7�P�!��'�72��D�X]x��ę>��ڹ�[�~Vu{��_}촍�^��G�ԁy��4_�ԍ�z�n<�d�ᠬ�l
>�Ǿ�r܏u,8O#���{��n��ޮ���\
�{��dnV
�T�I�z}��yl�(z%���"b���Ȁ_��ϹU>8׍G{�|C7��>�Y@.���<���k��8x�}�(�a��7Lu���E��"��;�،��	ظ�n�nc�Fx��Zvw��V��ߩQ�΀���t{����\9V�s�ꆽ�+9x�[�VzLh���f.Ι1f�Zř �����]��I���"�\�¬���t�=�͎��)�%��˼N�Y�r���5�Ν0C��Su�>L�v��.ĵ�1R���w>[ܨdO]E���O����<���R��՞Yc��xS�jr��M}�>%i#��M�5��_FO�I�t��Ǿܶ`è�}k3�|���D�ݐ�=�#\��Տd�A�y+ė�n'j�+tü��R���7�;'T\�Oi8��h3WX �{���ȏ:�jN}�Dw�uB�y��$��Z9�;P��x��e3R��}��v2�fd�F�#�Fu�f�y�v=s�I��ƣ{�B�	���9��>>�leR����H
�[ٞqܣ�)�OO������\���|}^�_��l�=��\$|�TW9%^��{Td�>��Z���=�C�J��|=��Z]���b�З7�zhm�5��7�����LLꫯm�W=k�R��4�>��򒊳Ĥn}8]Sb�X�u�Um�"y݇��ht���x���v�]aV5�}<l{��W��e{��:�q��m�Y(ԟ"���`LT� U�EDoo� �Kƽ�}A<��Ew���(�������[�T�Q�N���C��'@���GF��#���n{λ������낋�uG�~��o�|�o��_��!NQe�ɛ�VV��&�`�=P;�q^;�ʵT<�mҡx�[B�3SC�&o_<Z���[�Ewi�[Ο��,o
NX�\e>Ua�V!��T8{J�J�#�K�y|�tvp�L�K�3�qT�}s�sf���9Ιn�w�
�ȝ��+�&�ŵ�
X�9�,S:�X�)�҈�����·�u���a��WM
��L����!��F�x��5^�˃��S>�c��~�d����1��q� ]�Nv{�ew(^�; [>�(:�T* ��9����|����[��OS�_N�(�1~�F��[�V��Q�}{�)�_�U;,��Ϥ���z�&�.�3�9�}+N�X�oև��r�jU��7^��5�0��53�T��<��9�I�s�-����ו�b~��h�>�/ޫ
EKzLc�[�^�|U�o�_�6����>t<�>�8����?
@�L����^V���6:�J9�����G}R}R*���8'B|)z��q���>j�0xx���J9s,v��݆��LӽE�����NxbT�!����j=y��7��3Q{p�m����B�T5ywɳ�Q�[q����L�Y攍2_�x=7�챗�G����=�7��1{����Q9RY�n�ԏfO���V�'5s�Fv����{}�Co蝦2�kJ��|+N�3�ѝ,�����[l���9��W�[�t���}�uw��W~����vK��LeFMib�&w��\��k��ۿn�١Y��y#�D��T��XJ��-�m�-^�1���Z;���!;s����g@݊}
��S����������e�<��3y]n���-[M9����5	+�y�cܝ��<�X4�.���<pv*Qve��K�t�/��mu��9;�:��uF�]n./$����U&H���+��:7�=�hvG��F/0JF��𞺨~8�X��t�K&�u^ӕ>�qq���왏u��f7>\���s�3����uv�����H,ؙF���Ǒ�FC���Z����p��|����^W�������Z߽��8[�LZ���E�������sם/yCw�|9��Ȥ���FJe�}x%�w�q���2<wOF�}�vM�L��k�޾�Z{�{��>���9O�F-y,y�ϟQ	��߭�g}���Q;�[���{֥,��>\}�#M_��<����3�� Cy��W��^6�W�������7G7�5ZY��^��(6x��g�iW�.��S7>Z=q10�WH����,���z�+-V]q��B^����A\{��C>�*���i������d_[�@��2�뉐~������3�9��N�FG��J��l�b5�p��Z�y���O�	�H ���E�Idꣀ�����'/+�˧uC�/��î3h�[����}G��-;��h���#�:��x_)�S���77jG��U�[A|�W����xu��f۷�e� �J��ی'X*��=ؒ]b��Eܡ�Gm����-PӁ�@�B������i��5����Wu��6p�Ag)��&�g1h�z��$b��,{�]�����7�v[���9��h>OMς��kCþ3�,i�\X�'����T�`�X���	�[���w�6��3��+�M���,�9'������d�\FN��q�5{lw�ꗼ�]�K�`5Yy�y;Ӫ}n�+�}��Q�ʱW���t��=��KGn'j\e{��l֔��0fi��r��`>�FN�F��zH�d�K�=U�B��֋X't�Ix|���rR;W����Iss�[>�̕Gڤ�U"2��%�����	�
�����PQ�%�M(�#,y[��w��o(�j}GTg]¼��M���7<��r�_����~>틨�j!?k�>�{v���t����ءA� ��`��So�p�&S��/���X��=9��/Ţ���q���d~Nć��d��U���ώ� ���7�[ߑ���6sjt{�ԇ���梊�*&��gs���C���>������adC�th���D�)&�W��1�}���^�[�c��Fz�����3��JG�����_�=GxT;74N�n�ߣ�]zW������ԥu_����P6�e������Tw�:������U��=�"�\fY��ఁ��:��M�fL�Ee�Z���(��.��Ӛ}����=����)�Kծ��q�iu�)r�ƥ��Y!�9R�ȴ��I��r��P��Sї`q,�2�ޣ'�#����������^��{�H������߯Fz|j�.X�0`-Imx{��B�Q�9�FlЯ��SÄ�f\q�~-�TR�u�>��VG�z w��!����Y�x4�fOw�B�sr}2��q0|=jH�{p/�t�zm��p�<��|>�Mq����u�-�����ѫ,
�O�F��0���&鎼��땦E}�wǐ,g'b�H��,���?G�w��g���f��O�S�=a�j<�ĭ9��#���CW�V�w>&�\�3��ʝ��D�c���}s��~�ͫ%��;##�A�^sC��W��ܖ2��^���0����k%���8��;c�wKK}L�5Kj����_�G�T�'#ʈ����P�=����9s-�+wo�WT����i
�j>�uT+ͪ�z_�M�u�Db�`&m<�dN���T���+C�>�+��PU��.���ŗ�Yt�`��v֝f.�V�P�r���d�;�7Q�|��Y�t4���{��G�gV����[`x����Y�]�L�5������ަ���9m���X����è�R=�~� ��$s��m���u�	y�`[� ��x�W,�n5N�G/�ʵG��a��Y��<��kx�`(�֛���h�(!��u�\%a�2�w�(lܱ�E�kB6L�jG;$E^iރ������'v^���+��YY9N���4�qs=����E�U�y�EF%"Y�ze��=���L���V� ����9fyOU���+��I��>gs�O���q���|af��5|�����5<��#���^�{��z���*�Ӟͻ�,>�#ᇽ�ў�-���Ü� �)��;!ĺ4O�Ѫ��Ѧw�v����E@�S�D�h�Ϯ
4�|�<ǧ�>��^��0?W����(��Kڙ�VZ��c�]�U>�|��20�R�Z>�}pQx�EtC�ZG=��w�pt��ؤ��r��d�Z�@�G*d������õ20��9�i�ޗ��J����Y�u����=�뒥���Z�t�9�~����:�$E��/l]"f����>��P,eۅ(����3˼'�����S�1�}��3�>����˃V�%�Z=q7P��LM5[E�	�!zI����}�/��;;�d𿟦�Q~�[=�:�<r�����D�C�ץNG������r=���7iI���>���G|���^�,���,�9v<3��Q�y�(���+�o�����DWn�7�ڌ�z7�٧(�]�d:�r��C:�����V�%�_R�uJ7v�Yev�Q�U+�{����m��x���r,Ůp�n��WS��*�u��͂�AX�n�����vU[j��/�k�4Go�V�p%(N}�[�E7fek�
��YS"�L��N�S�����L��NW���r�&�X �`K���ುr���[�(�ڼ���Ik)��G�^����ޗ����\��Q��Z�O(���P	�3�\w4�ڝyc�<-�71pܽ��7nvI��b���kWj�x���or��CP������[Ө7s�^
�ȕݞ�gc@��Ï�;m�b�;����Ռ)�Z!=r�ѹu:�g�O&-�hm����襻��޾g$B:��j�\�-�!�(du/^�� ��)<}-���N�7|(�֔��;	т�`/'1�x��[v=���$�p��Wt����6+h��<-�}X�<j�"�͎Q�Э�T�n'2>���oJǯ���Et�cXj5����6�q��t4mlp����Ü�Z�u]��+D�-�t��t0�����hCu�#m�θ��f�Ep�Յ�&�p�N��"4���(��؟@���l���4��^*h��5!�l�����w�gj��#s�e��3���%�a�"���.0{�^c��$ھV�Ӥ��z�����u���(�5U��!�(�;R���%����P�&4gD@f��r��+��5��vv�o
���}8V��suѥk4v	+����j_?����/�n��Q^N�y�4B#Q��_.�+xsƘ����&oe�5�x}l�-��=���������N��\Dm��U�\/7����3q�9:�RY��,�n���֗p}�N�E^�<�|G��pV��{%�@]��6ب�l��ҽޭπ�F@��j2twcRթ�sgp�H�=�\0p*GzE��ê��� S�Qę}a��v���3F���	��_q�X޼�8�)��T����7C�Z�N���|�U�盉�]B�Cw���U�;�u�
��T��d:ئ��Ԭ����I��#�U��rU�}��*��;Ր>�LG6�;J]@rʎ�A|���Q��Q��b�y�m�Ngi��f]
���=f r�Y���Y��{M���;)�P�Hq���������u�no�EE�&��cT�Cv؃1!�JJ�A�EP��M����n5K��}�VMe�Ն�Fb�0}�K�R[b����(y�G'b�;�t�.�,s���;��>�dr�)��O*�@`#��=Q�i��a�i7w�����J�����8�m.�qq�JT�������2�- �Z)s�$��ā�+��A�:6�^�
��X;�TS��%A�Z���.�W�OX�X�1N���x+6g5�@� �{�c�w2�6�x1ڃ3���pk��aBt�/@Ƴ��^��9`�H�W�r�GgH�V��9�.w�A�Y����f��I$�)P��%$L�RiE���Q@Qr5aZ�N�Qp�r*�A��Qd�nAQ9�DD^��J�N�I'f)�����۪*r!v�R땞NuH����w=Ȫ�D�2'\�*�Z�;V�9�s�$Z��F%C�9:�T�C����O2��������u
�e�+B!1�����",�R������L��I�S�ّ"�����*(�;��a:�Q���M$�* ���i���p�+��哊z�q�qˑ�̣�]\�͕ATy�=�������n��ܩ$�u]l��U=ZAK��y냦S�Q�z�wRI�y''.�h�{s���&(�*u9�Z�Z.Zjh)Y�+��Ķ\��
��Ȫ!6(���$)�r']RB�ԮD�FAeqɻ��u�8W2]J���5ng=���r',�8t���Q!ŔQj�f�e/�������γ[����۰���ېt�o�5��^������םV���X�޾�!�oi3V��s�����!Ө���s2�r�����K�f�G7&}�O����3Q{p�n����~�>#LZ=�qw���n'�.��n¾Q��=���2��t�{�zp:�����,{�o:X�����8�ח�N��x@Gs{���l�ɽ�g���N}߲2����~\2R��r�<=*ׅi�Fz{:X��{��a5�k����u-]�з׾(��*9*���g�\,�Hv|����:X�s�-���O��^B:Ϋ��l^g�}y�C}��$\{]y�y\:��;�(�`���0�e���m=�9��ڲ��fzǺe���n⽑J�m�����s�u�{�du�����!(, �l�����^U��f�xv��<�T�蚆�K��^/>}wį*�F�^o�2����հ=���D�f������\=�z:@��<)�,	�n��Ojģ4��+!z�7���������3�y��n�l��=�3�4ˀg���}R-��c���!'��S�j���cDG�M�B��g���:L�F�F������9^��A��!��J�D�V.W�㓳�n��sp��;%*�Y<ܒ�:�;�ܖ;E�j�.9���og4��rB�뷚�E.�cD!�P{�7v����q�A;p�ΚX���9�s������y���.P��ۀ����)hZ���W�[�nj�A��rZM)�j)v��B��ث��������ِ`T[b�\-0a{n�123Ӆ�U���bz���ZeVz�����G�1�z�(g�U��m0V{נ<���n�m�-���<���h�=�~��N<3��^U�oJg�	���������<��TG�Őb�m�ld�ڭ����g� 3Ɖ����:�͢E��Mf���8��P���q��l�{΀�#�쎞OD����3��NeExnQ&��J܃,.7r¸����3k�j6X�3K��\'���{�|i���h�m�ğq��d�Ǿ�qS�ym�z,ݕ�%��>��v�k����\d�7k���Rc#�}�ݎ'��`{��#�#ӊ�9�G�G�*�\?m�1~@Oi���ۉڇ�^��D�p�c=]ˌ^S�[�g�k�5\g[׽$w��M��\:���B���Z/�wMė�ɭ�9Z�'�8B�Է���oAG�u�q����j�F�a�l��5�2�aև_ye�c#�E!(v�@�{B͟{�bj��w��L��鸢��Wp�2g}7��7��7���}�����Q�uT�F��4�g
����{\��0Uɩ�ܩy�E'��.e�uZ�o�b9Z�^����v�h�DZ�}kEMn"ߓ�EdëUs��V����5+����ڑ�}޺"]oN�τޫY�\�1g&�q���O7nb.�Gw��\Vj���)�����Y�ڨb����+6@�Pg��T����p�3j����N�h?#���z�"+��{�=�M���`��H���7)Te��,��d	F����S�/I��A���G�I��δ�5�}�����=��L�ϣ�.>�����Ǳ��v8�F����I)%,�w�F?�eY3�Y���H_�Nw���3�h!��:b��o�Dm��p�f�� �h��M@d99�q[;+�ܘ��aωH�2\P��4/�^��{�H���4U��ȿ���w9�
�M��fv�]Y�<6�{�5�Z��]^Ä�wP�~*<��d_�W���x�� �2�ew�[�N��P�@�F�3�$�����W�j��s�w �Q/C~q���~�g���}? '����v���������X��I��a��t�^z�u���#^φ�#,nY�rط5���{9+Hz�70��zPP�}�I���/��q7P��m�w���z�^���WG���Evv	�o!ӏ�}y|;ޚ'×�;���	���h�*<���������/.��U[K���▻�~ͬ�}p��vDhfwH�:���4��o��{1Y������
��ڕ�]n��#H�J�6�7 l�_mXK���V����{zA�W����1�-��m�X�ө�����f�7����T�.N�t����-�N�3heup��e
h;ζ��ڎ���G{��=��f���R�_�CUS�'�Ԏ_?mؑp�N
�!'N/�텗M�(�c&L-7;�Z�ڌ-G���O�}1��ZoO�zs��;�3h��j����C�=�]~�=��V;�`�Fd�v�P�nvX��ۅy>W7�����Z�@���5�E��o���;ت�R�;��&{yEEW��,;���_�Ǌ��L\k���Oz�n#�|Z񳛦��n��Vq����c�=��=�w��Q�8JD�`��0&�X�ɝ~���'(�BO��1��W[��މJ�{#�W�������S�V�6�ޱ�
�be�>�e�q��j�yV���U���=�@��{���������	h��>�]��)��;!�u3��=o��o�x���tDV�2n0���낋�uG��l�j�W�[գE{���sX߼*g�#Ti��ǻ����Y�7�D�	��W��An�;�����E�Uνix�y�����| �A���nf�r;YQ�=���3�-@ 7�LZ�\��XZqt�������Pg��^/�vh)%bH��NS1s�n�������I6�o�];K<�:G3�;��� =ݚQ������Y���#�n�V�LT6o-v����r��G�0�F����n�]�۵���D�tīFwd��pΨR�f
�aW�rI�\)'ϗv5�??|&k%��Q��۬n����\LL/TE�&i�x�+D��r�V�ʻ���n�L�ge�x��zg>�N ��̃���(���ۛ�}q��a���Mb��x^z��=(wg�5���[�_���� �z��3�7�L�.+:���>���g1|�/F�mn��9�=^�U�W���Z�_�D?U2���AZ(���=��*9�1�~���p1�D/�8��l{�7&=ћ^�q|L�׷������E�{���s�n5�}y���j�S{~��죅���ς�q;,eǧ��*��ic�3gK��Y�\3D#,�n=H�.�}��W��N�x�5uF���gM��{M�O���c.2kJ��
�z�o�ޕ�8�;���5���ki;��������+��ܸ֚�dAG��f�K��Led֖���6�.��Ozp��{���U�.5�2�΍^�ZϹQF*�JF�K�zc��g`�jk�w�=S����A�[��,��[�<��"�B�o�{�y�߽������h��ꗏ{}������-���H�VY>[u��S��6���n�F���t��9[�����:��������Q�;sO+;�}��ᵒ�kٮ�B��6]-��F+�X��6_[��u��)�PRnw$3 ���{�U�cɭn��J<'��P���G5���
e�}wķ�qN{��9�}��c��g2'<n��&�8�9���T5:���*�����n��Ojģm�\{ /����Ә{�����^��jg�Z�w^R>��O��k���r�/�Pz@�>���_d��w!��״����O����O�
��<������0�����qE��FF�I���J�X{їfyf�p��X�~:���=���]�W>�e�{i9��5�{2���7�\LL/El��+����_�\��������Rӛ3˧�W��$|2=J��{����`?uA)׍�.�����XG�\�~���o�vTa��+� y��ؘ��մn#O�{����?
�~���>t�X [��R�+_�;�A��yG �x�v�I,,�3a���!T_�d�z}G�j��|�Lms��'�^������vπ�}����G�֒Ǌ�%���y���N��Dl�&M|�X��W���:j'7�[���=�p��U>���*x����ǳ���~���G�Ó����Z=d�5�.����'ēfz�ݷ5�*�P��L�*��P:��1r����7Y~qР2��k3���]O���g^�P��I����y��Z��vq����TX�_f�2;�z��&�Ɩof�c@����<get�`g^a��<��n�CaW9q(��~v3��{|�����h),��eX���Θ� '�ܖ���C��^�t���iq���r/�ef�i��]�u�SO�C�J�\y����B���Eh��wI�f�z�"��޵oS���.��Tn�ڏ^:�7��5�R#63��m�e'<9y;C��>�ǉ����.A�֨h��vIgIB�N�b���d��o�&o�wq�z��=��_f�>#�U�GsR[�|Vnez>��|2!���϶D�Q3���`L_z��L�>�_��M1XZ�����]w���ƻI�������ǳ�8۵Q��Yeg� J5�z�S��o�'սS��g$��V�y�Wo�w��C���=��������q�ȅ4�p\���+���k��	��eMwf_?v��#���=��u��>y��B���2;�)ȍ����~���9�p��Cs3;WP97�Z�yC0�Vъ;���Ĵ}��
P��f�C�Sg�(����j�_���fp���׵�^��܀X}������ё��{A-�F�����w��~(�k�Z���v��ʟ�t_�����\�^�j>�wB]؊�Dn��S�81})Z�4��D�,���fr�Z�,9<)��fPx��|�5[ӻ{f>�]�z�w��<�.����J�q
��!U��䷪6������*j��&�%ޛ��Ot,�ܦ�<�x�R���=��e�__��*I,-&��S�ӹ �ӟ)����p�'{���z��kh��	�����5&��O�`[>%�3����I��ZdW��|z=hlP�ӌ�}{����	���x����:S�� z��$����D�#�u\en�";��i�~��l&���G�*O���3}^����I��F������V)� ��V����w��p�'�-��ҳ�	q�ѵ�cכK��ޞoi�6�_�}�U-I��:�=�/�Eh���>����u����	^��%�g�t�Ǭ������mV��g���lq�݁l�SWA��MO1��fiq�����w�枻?�N���3��b�쭸W�VoK}7�S�q�~&c�'�*�B��\�w�J�����|��F��\U���<md��K6lER��kK���L_��'-vv	J�qW����P~��V���?�l�5��yՔQ��Ĥn%��L=����S
��]���ʃծ�*�N���ۯ�<�����tg����ǲ���ի�Ͻ��`�v��ǔ�eLDWd�G,CG���czIOvk3�J��u��XE!���$�rLU��u�Mn<��;H��l��!K(�K�]���f�Kﳻ]s�s��!�AM�'��\WA�%�u8y�H������w6ӮN�U�w`}i�����e���3O���d�zsjaz�>�q�Ϗ?^���Selw�Ë���w�/=Xn�N��/��P¹�>}MB�?S�"o�+��D>�(��Ty|������]��0Ll���S`8o���t�=�������Cr���zhQn�7����&�7�Ts�RFL���Nz�z]L�.K&e�+Ok��{oף#�>��r`0�-U
����[/��)��,��Fz&}ۓv��㾊��H� �w�G=�]���"��S���G�&&�QN{�BY�nϧF���5���y��4ﾎ3�|���D��c�*~����
��̃V�%�Z=M�>�y];�	�zӊ��~�K��Q����=\e�Nh�����)Ϣ\�������	�t�s[�}���%�&�7�#+tüu�j#O������'b�.�ܳ�@�'.�xnN��-��"{�"�V��V��f�Y�L�v��l/�ڇf׸�}��3Q{p�[���ΪY��ڏ(�Q�f������6�}�۪��죆���r���ZnvX�~��鿴��y��_U~�}�&+��dc�lIz5�k�Lռ@K�(5���1f7�7��r���نc�,u���C��-�bu�+$D�S��F
.jg6��X��׵F�P��
�y�h����݈�����H7��
��>�sX��P�6��w#�V���N����,���%/1���E��>���Z;�]��7���&����6���2�~\2|��\�oJ��<=�?�����s'������6/<O�O����m�g���Wq���qO���wM�x|�*��j|����'7�|]v�ok+c�F��e�� o��X�S��ב�y\:�^�C��Z�e������>�<���d��-wS�^���ݥ҇z��bݨ��+1��SӜS9��W�Z��4�4JZ��u{�U�V�Qذ!��B�=5%�桁1޸w�A\-w�"W�ǰw��s})���%݂]���0�fW�1�꾿��Qg� �t��������7��v��J7�y��Q��9@�N��ᥫ2^����;�#�i��[������ 4z@�u�h��c�둚ϧ)�s�K;�/<E�/��U���1�ޅI��H�__��:��׉`@l��ʕ��1��]K�l�Ƒ�,��s�����b�)K��È~�gӇgF�wpDש����D{��^�����U������*����Դ�Ĵwq�Q�G��,�|��{�}����<����m����m���m�o��m�kcl����1��S`����6����lm�o�1�m����m��cl����cm�cl�[`���1�m����1��3`���66������6��cl����1����m��b��L��:S3
	�� � ���{ϻ ���Ø��� ��� $�

U %	IE ��*�
 (R� PP�*�R�QE�oCT�	UD���	B��T%D�T��QB�T)BJP��*���(�m-�BV���UP����EI�
Gf��QUTBUR*Q(�Q��J�H����ER�%*$��T�� 6��	��V�d�U�@�!��T(ѩAY�jh�`U@PRi@IV���  wC�RTMbU�`
��8wg@
 ����h��E ���t 5c@�@Z�5$RiB����B�  )QW&)(��UE(�,hRJ�ִi�-+���)l�1�Z�j�TT�A ���  p�]�Pi��&�� ����5��&Rj�[&��5Y1h([f�TѫP�V�I���TJ�   ���mj� �b#ki`�4h�������f�A�AM�` kM� ��3 P��m��*EER)  �j���VP���@i��0QZ��U�5�`�Z�CMl��cF�dcH��f�hF��T����� �Ցl4-X
�d� �-QAFV�h��ԭh[[Xf�(1b��	��j��X�P��H�P �� ��b�(T kk�[EF0�TM�h �5h
*��*�$֫F�*mQ��AB��
�R�� w3T
إ��P�Z��1�FV�h� Ѷ�U�j���f�)j��� ڬ����h0՛P�EQE��� u	!ђ Z*HTE�m�dM��kJj���,լ� �w�  P S�2�JR�@`��d�����)�@d�=@�L�  s �	������`���`E?�$z��L��a4�L!���A��@�L@CFSL�y#ȞSFcT�R	4�UJ  4    ���n�
�+����~��;�Xܡ���kԦ�"R��=h����� PESq���F���oU&�ЅERbį�>�����~���P0�P@ER	@\��L��D�b�""*����ۥ�jQ����ͷU/!��Ju�-!���P�Dr�a6L� ���G���f������5��0�b�R��Ga���6J�i���.�j�	�Y��$1�t��{&�ˎ����ї��m���Ҷ�b�]�� m��{{��p#JֆQe'[c�t�X�enV�f�Y���yYL�����X�LPb�'@B�呙P:��j�����Y�0@^��/p��4�5��ͧ�R��5�����$��W#x36�h̚-] ����Gh�3j-Ԅ�P��&�B��.�L�ee�(�V$� �o�A���\�"�q3��E��VR,e�V����tF�b�4�^��v��Y�Q��R'�V�`�l�M��.B&:4#*	[�O6��wkC-S�
7C2��i�Ō��@v���Vێ�Z���b�m����Z��k>c�9U՗J�4����>,���]�<xP奴�£؎�}�^=����Ml�8̬�c��V�-Cu��w ���i/�=�v\�~�9N^\�%ʫo �v��i���1�ԧ/E�ۣr���Y�v����>7[�l�r�hv��$ڢ�K=Z���սXL�"�s�ϋ�ur��0�t�ȵab6��P���KZ2�� �r�P�z�Ma��	zUelZ[͊n����^â�0٦�^�Q��ne�)h��K&�Ѵ�^V���C�}�U��Zc���B�*���Xd���2��)`<DK�x��`�Y��6��В)�Bv��,�tQ�IX+yZ�G�Z-ڦNŹ�f��5mЉ%�G7/oeA��"��w��EмGJ� ��0T ���ۗ��m�W2K_a�D:�!�&��W�&�ۡ�6 �[I@��WQ�Ӷ�m]^	��6��	��ƳQ 3Y�A;f�N��}W)Ԕm�U�~8��^e�D�V�=M�3c���[�R�IlW��ѥkX4��E1G,�[R�H�m^"��!#CF�"D��P��f-e;셙wzUf�t)Pǡ'�b�:��n�vY4��.�=��ح�<e�ֵ�N��H�6�5�2e����M�ܭH8qx
�A�MZ�gt!�lP���u��.�^k$�.۽쿳s▅K�kX�t@(��7����L�� �ٌ�^�p�`%X�Tǰ�-aƓvt�f@������v7���!��rek�}\�ŧ4|ţ�1�j�.]����0�
��4�J��������_�]-�&���̔#f�G>��l��S݉X����e�Dɚ-�%����"�`]�yńm��@S��%iu�Eon%�3rZ�ʸ�M@�]hn&�e�j*#v�죴���m��J���RQeۻ��.��K��K-+�l�v�̑`�)��Rf�vp�k*�ݩCr�V?�\үn�*	�J��n�ͤ���*7�ֳ�ոy�������-�ߘZZ�Q\��&@C��%��4bs*�ʲ*Acr�v���� p=ҖD���(���ȵ���
��k��s��YcJI��`�V�)Y���t+GU=�E���W��S�,٬z)6�弴Q�j���I�m�è����D�����/=w{�2�e�c�j���n(nfg�0:uKa�׸V�8
s�[��fj��s.��k,7��MD�@���Y��J�wjӸ�VX]�ն���0���ia�d��k�^��-E���z����CX2�Ͳ�ܔdj�J+t��jS*�Kub0�C�@]��1�dz�0��{M`��D��
��;�R�cPF�9h{p���-�JnZh�Rj���h����f��ٌfS��y�*����V���7�S�r(�d�1�͎�B���%k��p!��C��M�%{%�%����έ*�2�4��TPŇ@� :�aṂRQE*\
�|�!�����Pa��Yw
7�#s]j{`�A�޺O6��o�K���/
(��[��{�R	����N���T�R4�;9�8�v�pH�GN �����LU�c	2Ε�BбN�Vy���F��l65�^V�s�D�����t.�`�[{�򛉕L56������[/еmU/��H
�v��C8 ��b�mf���T��rU��p��#��Au%ޛl�[K#U�`�A��z����+	c�ȣT�ky/�[����G�Q� Fi���r��Rm�wc�R��a�ަάH�gl���c����	hH���G���TGX&���F�o(RP*6��Z_ő�B��'�j
�R"�����q����kI�"I�oq�a�a�$nQ4Uuw����>ޭ۱+]\��ni���٢є��@���h���sܴhe-|��GK�؅+ͭ��K�R�/���P��Z�,L���׻� 'v80�F6)+*����RH����Ӗ��`�
�c�`Х�l��ȱ!�´��Cby]A�dv��9����v�Sĕե�7g!V�n<ud�n){Y����8P®��nȖ�J:HvDk��EU�tFK�A͗eV���m����J���T�u������f֣�͠qc����m�Y�b��>ʂ�n/��pBի%�e8��u
me��=!��-�tȳp�[��mA�����{sA׸]K̅Ʊ�.�yN����6����ys5�s�i��?c�K�w�E�t�ZL�]Dby��`jլa�ֻ�DӂQ�h$\1M]mR,�JEbk�X�T�ӵSR�N���ur��A*4�&��%ɗ�pn����#�UG����ּ��H-5v�/�a��T�V�E�*�.��K :�͜�tc�yX��rL��a�����g}}ϫj5���ᗂ��"�l�`�)�Ek�pfQ`���=ێIO��W�VN�]����`*���;VYBW�/.��le��1�N��Zy�&���-_(��¾4��Z�-[����7IL��A$�j!��vPf�j�A9�L5Uֱy����ҜH��׋��:Q�H2���f����!V��ZǨ+5�N�u�f>�f�n���60�e�5a�����f,�Iv�-�a�v�i;e���7	��:���F�ٙ�m��L�Q��@4ԦO_��U�����c cjiB�p�Ef��ܱ�t��n�.�M�s%��3����Ren��.�y*-�s�0��x��IՕe�y5g+��<�����ڂ�c�u�.V��ӳ��%������I><Jf�7���G��o@3jbǵ��]N�^mm%JA<��{-*j�-�����sr�h^ɥT!e��N��}�4��ݻn��9E�:	*�J;[��nPI�e^|��k�T&�� L"VP�a�v�w�41�4n��p���3�zR�D"�h��3���5�X����Mݦ+I��/e�����-���MbR;�f��y,�yJ��K
���/�GF�#pę��X^᦯`��={ ��em`��sb{���c ��p��Y{Mf$j��Xէ,�]�G�=da��0V�$��V�ҵ�Cl:����5�u5�Ў�K�����ܕ����ê�੃r���k�ܩ�r+�$#�� �T�j�jN��j�lM4v��nt���"U��"Fm@��� zE�Ci�5j��X�>�N��+,�k7B�t��ڴ�/eJ#Uf�U��1���,fU�NڎD�54�ʛ>�pF�ܣ���j�������X���6��)��代�>�5Z�N�vIʰ���]u�,f<�x���غTn�f������(�R��ر�tH�S34�Ŏ�і�D]�$Omqo���V�V+����J���wp����Zl��dă��ѡP���iǎ�$zl������4tJ�Al�#�1�;�cSjJy���nk2�Gu�D�(;�R9 n���(���Ӭ�
x�`�����2%)��Mc�Q�&�A���X�3n�;�A܋u�]��Z�6v�����f�˙KW�l2�UH
�&��߲��n:��HB���2]���-�W�&�1�8h����gD���4M�f�c�	�*��#*֡���Zޫd��8����b��]
QőL�U���2���n�u���*m�uV֔���o7N�͉�ri���f�X�1s�N^����h35�Õ5�m;r��r�B�]�{2��5�f��ͺк���f�ko)�a-yN�5K�Se\6��7p-�(XU�����&^�!͘7&�XU�35�4&^��7&Q���̕#V����k둨�T.����+ �m�S�9HTY�Ee#0b%�B�V�-��\� Y� ᱊�R�&�� ��4�ܭ�	�>�
���U�,�պ�i�W�s[�԰v�0�ӷig�|l�ܦmJ�5����v�N�l�]`*�h�]�������9����bc�X6*8-6��˩���� �	�;i�NWe�,����@|��][k�^�;m8��kp�Г�!�v�h~���rN i,!Wn��1d�X�B
0LO4io��n+�xK-Ʀd�E�#%��s6�� �v���V��p�)�L�5��- *dhy����X}��*6�w���4�%j�/�W����2��{th�Է#��k3q�����'i䠅�H��^X�p��.�
�N���\�"8T���om�K�dڰ�/��Y�˫"��`�@����ɮ7�����L���u�U���n$��Xm�V7Q��X�I0�=Mn��iv�=�O�1�v_ZU@f��)J�E�]��m��D�m^m6�Tf�):�>��+�o#�:�z�n�LShX�K3/)��2�Ʋz���o5
�r3�0X���:�,��IZ�����	�R�����7Z5�Ce�J�+Պo+6�������Uwj�'5��	-��T"���A�wvk4]�uv"��.<���Vp�n`��!�ڛR���bS�-R� n�,T�Ճ�l��f����V��SR�r�X�P��Jݞ�40Z��GS�i������	|d�-��t�ʙ�ռ�N쳅7G W�=���n�C�S��{K1Hq�t���0jZ�]�������I��5����b�"�_[p��eM7l�K��H6��r�I�CVEyI���hU�۫�l�d�1����$XVF�
�w�ތ&�{�.�B�r��9��D�R��<��0��ڲ�sD���h�VrL���ڲ�=�`݌:kU3q�F|�H-�xl���f�Y�8<�/6�d[��t��u��e k)i]	B�/Q����]����X�REw��orve���c�]j�VX������2�Q	6G4��c�%��Rg5�zE!��Z�8�P��nbuxj 2n�H���h �}�u���W��Z��w~�u���ퟟ���'�D��^�G�M�9��W��������l����M�_v[��%Cj�Aq��w[�\^�F��ZN4ۭMl��ݜ#B�{�5[�Wzn���=9�P�3)=�I.ǺW�k�����O�Ͱt=��WhC@�{FY��~jzX*�<�S��%&�r]��0�c�:�.�R���Ar�C6�,<u�)�����h�'���ʠ��5z�1��X˹yd�p�j�l��G4Lo���$�˝qh����m|]De��Y�6�/ �J���>v,�\�����t�
̆[��ˮ�'ds��Y���屁FJ��� �8�K{�x�N,ם�5:G���wo����a���Rj�LX�i�4io�v.S���]`��44S.�>�xX��}
nfBY�|B��PUǵ�7r�f�	�8���3 ��v��傃�k��\
p̃����k�7p���e1�ݍ2�M�l#�!mڮ�'Q]U�MFHkf�ↅ����{i�!�%�\S�o�,����u��6���!���Nem�;��+MऔIޚ$���0��H�d��y�]"r�rf`���e�W��q��Jf6�t����A�e4�̭y����֯q���}LƜ(҉���$[��M׽�Fd�Ѯ�>��k�z�dd�89��聎o>�*ص����NH�^�uׅ�lx��Z�2cH�U�wzk�ԕdWy^v�q�<�ݣ��d\d�Z�����������'l��L��7�^�m7YD2�X�ИӜ :fQ}_u�`�� R�_b��w�A���X�Q�Q�`v����M�/9��ݼ���g��:���w��-V������;c{�+�s;�;�UfPJ��܁��x�<�o����ka��k�T�v����Ja�殄neē��ѫ�����r>[1��B�Y�3\i]�Ų������0)*MK_f�B�̺��c�ǋ �ۧ��680qv4؂`�TB&��v�̃��5�O���(K[h��e��j�K�#��nLf�d�j��/y%N�Z���])=��gs�*��_;�m�wه�4�L�J.�i��T��ª�����ژ�H��a�����յl�����i=��f��*��G�՗��G=��<�����>�鵯6�=U�S�qs:d�T�G�#+��/^ҫY�*
-��f�s����n�*r&����S�����qvn��K�{(�p�(Xkt�Z,��7/���v���&�7EndDH[t��ݩvڦY�7rRoKw9�33r]Ѷ����m�h��C��v�]]���DVŒ4 -�B�[u���9��ˎs��J��[*��zX�l���nY�¾�5���#�^9ֲ4�'o$����N�h��pE��������j�*��9f��[P�8^��=K����D��-Yn՘z�o����:�h9�5,����k�x�k�u�+���7�l�90
n�aŊ�]����n�+q|p�wX�'VS�E	��-g[a��l�9��[����U��b����fm�5�q��=մ*������O�o���/r����cv�4�Z�i�p�]�޶�ʷ2��<.���յ�=&��jQ,2R�X�۸5��jh�)i[}C�B�n
�B�aS�`pħvo�M�i��F�=w�%d��@h�8;=h�!зp�ӥXP=�*y�;��Zp�YӪ^�^ǹО����^���]2��[,≗'mgF�0�����{ljӆ�в��V��vˡ�V9�t݄j�7���6��nP@m��ҭ���T���*�P�亻�:�鴉ɩR`��[�ЯFr��ېM�16���� #+����)�����W�9=�ɖ��&�k��;$�9`x�R�퀤�ch�n�ip�_\ʗ���^>7˜�B���ȂRCiN7��D�f�=�w�(5j��&_9�X����7���=�ܙV�a��*V�f��-�'s��1�2�"��δ�0.7��1w<Ј�Wݘ���+kC"�e���U4NY,��y�ta�ec5�� ����N@Q�ṁ(\�Ru.�WV�j#{QxuI;LrȽ�u�iھ�:0��� �T��f�\�bU�u��(�gd����Jw;_g�uw}3y<�}-��mޙ�e���&�M�é.�f�{��f���u�%�n(���HE�䷴Y]�8uGuc�vJ�L���ʧ�myct��b�l���0��+�r����]4wF$ѨQ�'��+N3UCҦv�h�����gK\������C���j]�F��z�u��^�5ȓ�h���V2��9V^���2>kc*�
�z�z���}���y}X��!1�mLk֥}��Z���ݩ�81���9�(gtpY��{387��Gm`�7�z�bRl�e�P�s3q[��c�o*X���TQ�ga�ʫ���A;&wې�K�)CV,��E�� �o͂�+/iАI�W��e���V��J\v��0.�I� ���wg7\��b�B5�S�T1䖐��5J��N�7n�wmkmBt[��r��q��\+jZ�D�a=p��ږ�}����Sh��:�����%=���kDx�WIj��qV��Qmɽ�P�u��@"2���KW����b8~z����7m=�4��s����ao���kG>eF
4�M�5z������m���c�a���cwB$����+�#���E��Ѐ���>Ϋ��n�7���#����8niB���m���Sv� A`gT�����Z��7�%�h"죁����f%b*�.#Hݣ�����3�7�Ž���z]�}(���E��ۦ�p�^��p5*MŻύ8e�<�0���8��.��z�g,ɋ+ji��v��G�"��6�W��UX���p�\i���+�.�R�����A�KOZEݾ��Ǯ� @���Wt����@��0�񥴹���)�Umt��`���h�Y[�#è�-\�6q���V+(�9��LKr9�7�6�<�M9��X���]M�� ���V��m�m]��ʧ�k�%��'��kGy��<��Y#cl�ȹyF�yp�X�]0�������DR�zu��Wc�I]i̼���E$@9�d�Հ-1��}�R�t�M��E�wK7dí�$�:�����l��oh0�1�*�c�i���"Q�Q����(sz�ׄ=>��V�cB�-�8&��jVl"午rV���N�ƫ3��z�V�v�k�.�:U73�(�����gO���Ĳ�1Fȭ�t��K:E0	�Y�!ی�3c��\��~ �b�PV�;��_d�:X�dL�+�%ۑ���@�*�9vX4�SՔ��%��v?�:3��ַ�1�!�u�n�ښ	[9��{p6��lԈ��r���І�`Ǡ���i4��Q��{׵������Xpۄ�.5���{Z���Wb��W:��(�n�Vm3�p��U9L|ﵼԦ�A0��uȎ��������E��S#���ۺ]7��*|+��ӰdaÏ{�Ƥ�jZ�n�f{��Sp�+P.���\�M�-��o1���p{Q��%��")ƙ;y	��+���/�
,v��W�!%�1e�˝hh��b�ԣBbv�A��Y2Ac/�TČ����򳜦s�v��
��37l�1�;��{k��]k�
s�֐��<V��i��:��I���Vʱ�+2Q�A���s�j�ń���� ��5��� �S�=���@��V��Y 2�:�ve��]CL.��M�s�cea<����Z��M���9�Ω����;����+	P�@�Y|�oK5,�΁<����{�b4�f��w���r���w2�|û�����|w5`�����\���G\�D�iY3I�佂��k22뚻��0n^�8� K=8�Y��ƺP�f
��f�Z�5�y;���zq��g5����l
K�M��'��L;k9MNAu���c�5C;���P'\�<ƣg޹��;7j^�r��\Ց�7fL�Dk4�;��g�l�q�B�%�Gg�u�	H%��uv��c��Z����u<�'u�;:�"����S��ԛ�J��	"'�i/KWӻ�� �NS�m�ј�6i�ݠ]k&�1ܝ����k��]֛�����H�(v�Pԫ����v��}��KwQw�*!ū},�����Q���7�����{�$x�u�RX6�g�_��ykד�F�N��&G�m��%�S8�+jQ���;YueN�M�d;f�]_�ӎ7W܂�����x��/
؄��4e����)`�d�����+�*���	�������F2�;�]*�����tաm�KEԹS�`x�5qsf�K��dB݁��ڏ�*]_
�mrr�%ʏ_1�v��1�I��)����j���jQ���Z�^[=;�ppѨ�Ȳ^��J:��R��#�0$�ߍ�ǈY�ӱ�/���(%Z�X傋%��Cb�tY��md�퀫 �\��.!Yw,�e�db4��t|�{o�sP1.l��X�V��\$��|kqC;/Af;�(�Ť��*�{&��n%�u{��f��ڀ�����TnjD��k;����t����,�����U'��^=�o{��rb
�x�����[T����^�����{G����-:O1�3�
`57���������WC�����C2ʜBM�*D_AyN��ɦFLO�j�q�����}�g�(`T�A����\���)��.�7�"5��D��N�(g,@}ת��e�I��@u���ìR>kh��}��o.q��n(-����M:�v랹FH��p3%���ݏ�"��b�fh�n�|��奛s��R�X9���,�454��6#B�����u�l%u4S{��*�:p���5�c-s���h�S��K՛w�%�O$�"(��E��O*�oIy�A����r�+xJQa�����}O)�[���x��󚧘.t�9��%`���q�$�,�C�^Wx�wMmL��
��&�i֌�����,��#L\Ó9���D�^�:�Y�ѭy\+��[�Sd�|x�����,�
��vx��Lt���a���[���\�������LzjL���o+!60�^���r>�Λ���PvPe�x�)�{n�lV�E!F=�x�fS<���O�M�I��Ŷ�^���vb��+@x�Q�P[E�6�˝V�x�oh��0��%��S��CS��i�R�Of+
{�[�F:٩
Xo�����;���q��i��:G�T ���4Kߥ�ȧ�9��[�d�t���Z���?,}�wbhw�3F�|U^�A� �釾,��*��J"�t*�T�r��F�O�װ�c5�9看{ESMI�<j"�gk�8%�e��p=72�3�[�!~`_�if��ۥ{����Q�f<��p��`�,��v����b�F���oL7Z�n�X��q'(ȃ���#�'_o+�k6����25���;�����茠�Ȝ� �ֻ�����o OJ
��(q''a}��L���[1Vm�r��i&���hU��Wp����������/:��kª�lw>Bq��vɦ�7b�!&�2��{��U�[�Ye�\��.�C���ʉ�����-9������[2V\��0ݨ���i΁LT�ө�U�|����n�uև�b����vw"���
��ר(�g��;��d_,
�9+(.;�c=%����ϱ�!o0�#W)m�-��) �����@��������&.�H����-�nu�Nrl!,�Z.Ĥ�|���ˮ�YC����F�����<J��n�*%��
��P"�2
3qmr뮅��*6u�QN��r��ri�	�qe*��'�(�%_O�Q>��F���������TY�X�����K�k��Lb�PY)�Ԋd�o:�a633�oQ��k43��Z�F�6`��/���*����t�;�:eM.�ۓ#�&-G;>��q�+�7��$�i�y>(<b�(��=�<�kbT����)m۽����1b�Cņ-uy�'J&)�j����v��:��;�%v�-AY*�<���v�"����viF�Ȇ��U�J
 ��1Z��n�-�X=AQfu��^
����m:��7��̙s�oÖaS]nҰ����iN�S�)���\	��>xf��5�\m�YOQ�"Q���9.Zѳd;îݙ͛R�e���4�;�{�TwE+U�Aַ���Wf_X�D�K�[�Y���b�O��8uk�:.���/�t��7N��W6�����̩H]���l	�2f�GWd�*�Z���`���
��{-�rp�B���Ӧ]��n��T�f#EbK��jm6,�ed�\�9�l��N��A�/q=96�yb��(mf��+̅	�}�t�)�6���2}w�:u���ޠ��1�q��m��0e���6��/\�ݘ- ��Ζ�7�[��%+��8�4�x�j�[6أ6�`���u)�P����w;B��ke�rY!��5��Y7oA���y5��V�1�^.�x�ThQ�Q З�jN"�i�p��.f�Bd�G��O�|�B,�:�5��h�ر���5|�*��O�Փ� ^��+�h�ɕw���Ħ�s�����]`f}yv�Cv�f�v��7���۱��A�:%� �3��a��M�Vf��%������1+yMȞ���:�O�QN��ssbC784����f�V0i�<���[��i�"��֖	�{�Ī&�3lؕ�i[[NZ�����٩CoR��2���<_�WY	�������N�"���e��{Qv7����̔�!2��}f"� Ѵj#��k_
{ENf&k������솈tz�[Ve�Ыm�7�m��MkQ��S�{V��?E�-�L���������-���2렦�{,��˷B�}qGOF�NX�Ƥ�Z��M�J����q:��z1��7���\b���ʦ�w�#�����gS�PX��;���vŜ�{־s^�[��[��8�fm>���/��Rnvo�.�հ�1��R�ZY9���"��ͭ#�ͨWd�0:�W*�s]�Pp�Q��;]9OK��X���54�
��m�ܙ`9F�lE�(P��p�l�qI�>y ��L���P1;v|l�i�%a���Ӡ�(,�|���A=[i�K0!��1�:���3W��Wo��}-g*�`u�P�7���
g2s������R�uZ݌�� J��\�l�jM�g*��J�+�<;��Mu,��sc��̮�����:b��Baڕ6����L�j�}zݵ8���7=@#��܊Y�4��*�=���Y������۱m����"[�\��}�`Ɨ`Z$&inX�oWf.u�3tR�����qDU��9��sl���H�oJ̈́�l�'�{��F;��xݧ(�5�����E`/5��YK�.��ȫR��h\rٵ@�jQ	�"��Kko4��S)
j���l�^�͝���E ݂ӫ��{1��"���ò��8���FE�]�
8%������+7��P�d��+2��(-�nXs������t8@n�p��:Uf�*�Qҗ�H+[�,2��Զ�;ل7Ue�Y!E�G�u�T�W��@����;���J��$F�P�}۴�u����-�;ra�a�N6�r�v���cd@�lX=S��.����F�]�#]��WV
V����cE��>�F'ٱȿ��
�%���ܡ�\E�E�1�����"���՟.���'z��g�,ٹR�B�xIP�C6��U^���5[�IV�����`�cTV>����	�r&�Ի�1ݬ]}������i��ڽ��*�ȑ��{��3Q�Q�ږ�vv��vÂ�rb���*�\)t��v�/nք�Nv`���z3�k]f�T������ E�C����/hH������+z>cr:䴼z%W�N�&L�j�wx\p5�n��m��Ur�gef�$YK���;�2z��#5�:�=2Pp�O.w�[]�ΞW����J��i��z�%�%���1�N!q��������������ݶ����W�WB�r���N��h�e�m�y�	+�9�̧��ȡ�`$���b�D����ē��M��I�t:e,�4k,���m4��7wY�3[̱��>�w����71	��xb�G7R[J������&�_!�M�����h�s��	����I+��"zIY��T많�t��4w�S���͵0l;6�;���}P�g[�x[��Zme.�؜�����2�$�	�SoOu]�n���U�z\�̥�-aX�r�Z�vb8IW��rX8�Z���%��pG2=��":v�[�ԃV��`ж��j�ݶ��Ҧ���s�X9!tAm@�6��p�|�>5�Y@�h�1v�ZwYZ�)������U̜G[�aŧ��06�y�/�z�aU�!G�c�5��)�;��s��7����;J�on�z�������\D���-�r��,vا���K�F�ݓ]ΣET[�c:�ܷ@�h�]LQ�|�\G�f��ą�Э{�E�^��1��ج��(14�[�ܼ���h�_/��wC|м��l�a��L�w\�@T�����j�j!J�\�/��zt�R��|q�y���X��pm�O �_ e�n�1��� E�j����**/%$�1]�ב��ŷ����Wp��z-�F�mT��]i]�=Y�y�(��Ցތ�4#qAb�PǱ�7.ًm�=�:����;dfӴX��]�j��h
�hֹ��[q��>� �H���/��M�e��)F�*��{͋�r�Ol�σ.�+h��t����CP�#J�3`3�7vɵVmټ2$�U,X,�(뙺��\W�"�-��F���MGحF��\�޵��n���i�	́�+z�n�Zѣ��2dR����( ��v�\��­���bŒ�bC)��ڴ�d�6u�
=׺�j7�w&��r�͓�ߵu�ӬiI�MCyV���ef*��Gp�,�gnVC����2zڂ|.�J�a�_Q���mw,Gm�r�[(&�>��ϻN�{\'bv��FBT�5�/��>�R�*��w���WML�if��4�B���q2��z��Iw����`v��RdY��ꛨ5,����pJ�9d�v*=�a�Yݠ�|�p�sI�"ۜ�+j�ֻ��A�ѩ��������f��n�ī++CWwǞ;v"�45�`�.v��{�����ol�;����ϕ=r�C�߯^��Khq��^��)kd�v��Eo��]>�o�DnD,��b�v���7v�G�;9aJT��a��ᓬ��/�Ӽ�%PӲ��� Zy�篮�1Hr�J�Ǫ�r.�M.gL��:��V�)b�`�JU�U9w�)C6^U�A�B0R,t�+[���m�y �T�r�!۳���\��]�22C,Й��f�N�M]:�t�횕x�����M��4^�h?3�����=$D*
���� �(�+7��p:v�L��+n���$���i��M���d1!Vf�2����*���W0N�˨�p���mJ�k�;q�����X{I�����N8��"Φ+Dـ'DZ��W.��BeՊ�ܧv�4��7�:�x;���`���� -y9%2���E��I�J���jQ�`5��Lެ�.t���ұ#��b��μ��k���-X�	᪦R�g�.�h0�f­̴>ɲ@�]/�j���α�(���d�����i����>�E9�A��c��u�Vu�^�ꚭ�u�^md��H�N��[[E]X˼Iخ��c@����vaO� �R���U����.��I��1�3����a60m�l7L
��%��ƅoduy��%��nfB�K�+�K��%�nZub��kr�Q%l��lt���e�b�����D��/������$��[�[#�U]0l�� �<�Xr�Q����][xIgE!�f���eѭ�@�+7Oh�i&�c-�㺇*d��;�+�9v���Mg//o��}�:	�[�v!X�W��m)u��bgb6u�#'��$��I�,лD�'�B� /i���ֹ�CB�#�|�nu�h�J�J��D݉��a���`ő����qE:7crtٵ��z0r�'Pׇi��e���#{�CQ!C�W.�	�X��Pb]YX�t��]��NE���
m��(�$MI�XSpwm��[��-]�s�"���7LR�V�LUɭ��y)Y��5�;�: \![Z��[ċ�%B��M>��ӳ�Y*�=|�md����%47-JU��15q����ٕy�Q�n2f��a{F ��٦���[/�v.�W2�����EWS@��b��ڭAs4�+���o�R{c�k�TΠ2 ��A)��,ÿF�X%K1<]j���� �������:�:&Q$M*�s�����V�d7H����m��Z�:�'��}����HY������ tR�ٴwΓ��&fQp�utӔ{2r;���M��j��,����P5��E�F��H���.\ϱ�Ѻ�Y��ቀ���*��Ə<�&CJ��9�
�1#׬��eZ�#oyeJ�x_1�� �1cB,"���[a�O�ټxڢK��gp��] �봛��
Yn�������9�d�����ꪨI �,�`rL�yː�*08w�H����2�~G�b�����s_\����c�e�-\�t
\��@E�u��q�zx�%"{T
���c-K�YO1���Y{W���n*�[{,LwQ���;�<����Lg��l��PVL�\�lƠ��j���U\��#z�3��g=�ݳ>����/Y�C���*ly�cJ�^$z�CK��S�R�'uJ�ޓ�}\�W����ި���;}��	D����/���-�LEiޖ�L��>Gs#,nVu��&&���<��Z����zV���ٕ$=5�&��6;���J�+En������2;��\o ���e�FA|��p�Yus,�԰>\�tR��V�gf�w�]-�n�$���\4T栗h_@� *qÎ�`�V\��+:��v���#E�X��5���C�g��Krn
�"�]躺f�D-#f���.5��S-^�Q̤��C��5P7[|��.0���8E7�Z���CGp�-h�w�u<ʴ��O|�9�v���ǜ�|eY�ҰNm�jh���P�/�D�:/�o2�n�:9��zkEX�y�Z���ox)AqqY������L9�2s�Z�۩�9���Q�l{Ȧ]�;���#"�U��b,TF(cr�-Sm��J$eJV�0fefY[j��-.dZ�E ��AB�1QK���T�*b�/GF����YmF[J����mEq(ff%e��KkZ�`�mk��9eh4VJ%1�1(��J�*��T�s
���U�����bE`����uh��er�I����b����m�H�jcD�T�1�[h1���2�b�YEUb"�رDZ�#m�EK+*�m�X\BԖj�YUPr�˔m�YKh������[-��QPY-3�EUX#i(̵�ڻ��/�_��_�3|R���ONQ�ᓛ��U�����`������'u�약����u��c��,msJm}e6��[�{?���?>��k�eJ?w�w�v�з?�l�|�����o{�h߼�����f�ٝ���I�R����C�f����^Y���KT�	���K��K:�hz
��?б��U�s.�]wts'��xV��д��ø�1��JtyW��rz���:&l&�2i���^g��"d�~�<�l�I�Ѿ�f�s\����2i�АG�<t��k��yThf���>��.	�ؑ�}1\�P����1�j���z���~����:ޖ�H��zvW���d�zeH��^5����)p���t;�\޼龇����o��"����G�v��(���0�CG2 �n!��J�2^�.��-�R5���ġ��E}��noe����:�*�a��S�;�|�V7�2��O�s�CF��0jDbO6o��Ě�7+��gvq8�bL򫬆_�~��Ԍ��������W�k1uNe;��X��S�۝�����M~Jm�ߵ�9�2`�s{�6�#�+A
���D1��mZ����K�fn�vz��ڣ&5�ue�+C\�vy�x�9;��m�Q{6�Y�55�o9S�J�'l/T��zN�r��zP�ƶ�]k�����I�H*G����r�c���=��'
�w�26�?�$3S��������\ĸQgw!l�nt�dnx���_���*F���~�Q�ۣ���'����hP�
1]a�:LMg{�M��YS�c�t��\�����ɯ�p�b�h���฾_7-CN�ՙ�Yޱ��3�n�VͰ/%tY���wWx��Q٘��MIN}�E��C%���.b�>g(��}�tՇ��k,&�	Νӛ8pϱ�]��5u%
��63�C7�ޤ�����H���7�*b׽$�%�rA��Ƴ+�S��F�F؏����uy��y�u��Z�u.��P���p�|b�H�k��e�\���<繣68k��*=<2�s\*�~������q�����ݙ@���Ndc=��R�DȽy��ر�O�[�"�=���YU�OD�=f�)YR��I�=�tg�<���A�ܮ����tc����V��7&E�J�/Mq��3�;��w�-}��<53�`����XF{8�=�U�Z=��o�6�p��H��k�_�kM_[Ac
�}7�߲��k���`�W����x���X�P����k^e_�>žӧ+������7W���F�=�(�D��3s3�̜e��ij�[]b���q�$���$o_n
ndɤP��m������V{z��ӑ����,��w��5%˞�u5o�ڌfx��6��ٕh[�x�uǏ��	7�#�b�%��:6�w`�({}yu��{��'�,t��x+[B��6)��gm3[\4��F�c.]�Y�4�u��k��f�<lhjvg��cݾ~��.1{�u	I])����s���ٻ��Q�]�6Gr���x+�ҫ�U��Nw��]�I�ܥ��Q��ᝬ�ݺ����`�2�b���L�t�i�1\�]M��6����%�ځ�-Q<�1u3�WAΨ9n�9��*���qTW�p�Tޑ�����Bg����<������Ƹ�xtm��E]T�+>��.�iv��5WIʳ�Cxj�f¨�m�6�Z�����]�3I�Zjggw�z���h�TƄ���wzh\��T��/��쬹���t�$P�څ�ÎG���BM0���QR��|��/��9�>z�ŗW��c�^^~�䛂k��[�v-�p!N��9*w��Gvyz���f���et�i�[�=3���i�����d+�5YuU���)ʞ�>�C��G�=��[�r��S��9�z���1�d���}3��oH��χ����<�7�y+�9�����'x�o�N}^�>W���寺|)ӳ�d�y��'���u���/�t�sYjAG��>{�B����[���^�O4:Y���γ:���֧��'@p�Q�{z�b0�ew�3���ӏ���P�M�I�C�y�Ͻ�VE8��{�v���6kwp_��~�Ʌ��w�w�3�mJ��_4u��3][�*r����c9B��wk4R��M�%�Dmqy!�yv�u�B&��zv �\�ݣY�:�����ղ0Mv��i�PX}8c���ӂx��*�n]T�{seΑ��vKHU�=��f�}1_Ӊ]1Wg�{y��M��F�����%�����]_r��ܖ�%���;��}k:"�W��T���o�,Eq���_oet�5��O}��zwn�{��o�ز�I���Ӳ���{	��2C�\C��{���k�gf}|�N_[�c͙�����3i��-M���o�~{|x��w��ZmV�/7ʰ���3Xzz���{#;��Bՙ]s�u��;��2}�?��_<f�LXL���H7�Κ�~�՝�ÆV׎�_ۋS�g�-�o��0J��=���N�S�ѲMz�]J��ܵ	�U��[Q��އ�j��
��N̙)��|�f�c�O^ƯZpU���O-i�.�c��H�љ����_S����k��L��ɸK!��Wo����3Nl��2!���\����I�w2���>�]�i�n��Ee|�}�!�B���v ��z\c�JV/hE���ך���>�D�|`r/
y�
��b��t�B�gB7b���T�/l\�-����n�u��d���Wn&��3/�Zϼ�p\&1��;�F�aG�%%����n^�ކ�ղy;<=�]q���.��j9��W�Ӻ'g�3�;�j��Q��]�.5Ҕ���gt�"gs-�O�+��f���e�,F1��{lf����8{��ُ����Ƽt��۟S�{�U<H¯|�n��A��lH�>���k�m2��J���ʹ�����C׵t�v�K�i�=[�qhJD0�[l��*(fgˮo�Q��ep�~����F�C�zQ��1ꐎc^I݆���sz:͆R�~�e.�}Z�7��o�P�K}���{LҼ3ګ�;[��?o�_4�C�vpo�}�țn	�
��Us�ɋh5y��po�=��d^�>�/L3��<��K�ãB���aͦ_�>þ�:Zf���W������)���9}�/�u��}��֭�бQ}�N(n�����xx��]D?3���<o�ٶ�f�G�;�V�{9�S��o+xq�x������;�b�-���m$��n�{�4�y�(d��>\���������a�����^���EF|{���}b�c���Y�a���ez��s���h��h(%��"�t���y�ɲ�ez��6��$᭫��&�d���2��˅���Bh`����ٍ�<k-��k���'���]wf�c��dsƟ|�Ѓv�ooM$bp�yE�����k�C�W����<RI�%���5���Q�;]*��B�V�<ݐ���������d�;ԪN=%�}8����w�tky׌0�^M�ˎ\�M˖#���2�"�쏵��'VΙ��Ƹn������ɡ�n����K�����]���@ߘ�^�IH=m��o"K�gz��.�-�������n��5	PK�| �7��-ulQpﻊ���������I<��s%W������˫Onu[�C%�R~�7/����z�3�j#f���F�U����w^7���v�_�~�W���v[��|�7�]b��B���g��7�X�̧��g��1�r����Ǹ֍�9yF|�T�m�6y]_��}[���NT�,JAv�*�>�f�Xu�b���}on[tn�p4��py0�	�fv5+l>���ٟf���ӡ���(�'&Y������&���gm�$mBJ�jD.�����߀C��>��]yf ��p���9;k���vL�|`�ɍ'N���1
�|�~4��"(1�\C���Hx虮+��%���3�/f���ٵB�ܭ�׫w�G���S�)И��bp���f�n��ϼ{���c=o��{>D<�p���G�h�*���e��~;kW��;󩝕*���Bkg�/N'� ^�e,�{���Y�ɷWN��U�w1�JNOG�)s�Üssʭ�Zy�L�<1��ܩp��1c=Щ��x�^�둻���+Љe�M�����/~U&��+5�||;hvZǽ7��3���;~yجu�}����A���l�h��D>�_��7J4?����mW���:��,��P���k���3��L���i�u��ݦP��{��\��$T�>Q^V�������mf��ZE`�.�VA��I���m�{D��N�uΰ��w+5�%>
����5���ά7Z~Ӧ79Y$j�2;�vp�F�kd@ri�v`�H[��_UY��U��ݡ\1�'�>ۼ&o�>D�t���I�⺣��ٖ�V(�ԛ����ו���T��#<�yI�Ø��e޵�4k}ͦ�����Hc��l�4]T�ݨ�+�ИyJ,���u�Dq��H�νW�7��WM�I�W��3\���]�yLR�rp"梅,�ܟq `]ȴ�ld����BMNغR�Y�(l;x)�lK*ʬ諥w`r� ^S�."ȭ���Q<��8gX��E\ѥа�ZqdP�M����W+_m-�r/Of�giV6A�;Y-Y�����0^���d<�V�HSS����ը��fŶ�Q��x�*��iLg+a�#� �i��!�/;P�B��ᐍm�����Rg1\z뭜���CY}�%�����?*{SI�hM��.=��C��:�l��=;i+����s�Y���~���hP��G����!T�N�6��bҬ`ݢ��Z��r�Y
�_a���� �J�h��Y"ʩ�j��'"��$��:U�J��:�ve1feM�Y�t�Q^Jr#xnf)0����H�%���+((R>;Rj�l?������;� �(��zU�9�v�e�'�֊)ў_u-qF@d�;�ʈB�N��n���l��F��d�FVT�� <:�@�H[�=���&��b�]r�d�6Z���j�V�YN��l%oR]g�k�K�7cB+`@qVZ�!
g�Ac6A�gUՙEp=�r�.�%��Yӳf%Fk��B�2�!͍U�F9M^;�OA�����tub]9t��(WKW�Mp�EVYU�Z�u�.��ӻ2�O�2f���ۭ3���\ѧ�S\�v��-�Nh:��t��r�ح;̦��]�;�]a�v�#	d��,��>ec �튽�l��6��ȍ�i���d�^�cq-s�M��&�y��v!���3vx"��/�~��H����u����o��,�C���p�N�{3��?(�$�I?~!"�R�Z�U���O�aX�X�+i���QAp���kEU
����c�kF�Z��6�k"e+��5�\�+2"3+K�U" ���mr��ګZ�h[TQ�.Dem�QU�m�bD-(e�QUQ�Fe,UjQC-@�bV�e���pD�J�\sKK2�8�c�2X�j9�L���b6�mAA(�c[mY��ն��UX�J�R�Ѫ�#R�j2�J�T��)m(--��K,Z��ѵ�m)IT�KV�5�)TEpZZP���ES-���q��T�n9�LK2э*V��%
�V�U`�J���K[mr�jܸ�qir�`�*�mh�\���)��m1���R&c�����-�(ѣR�.\TDX�7m�m`�r�Ō�̹q�e0f%s2Ui�~�����W����q��d�s^b�ח����1�s���v�<pJฆ&0�^��׸�K����m�e0��&7æ2hn!3�q���؟��[%�홷����*>�{��l#u�j�����yz��O{zd^����zK��)�\����U�����_�3�����9�YKEz������N���y����ق߻��h��C�/j�P�پw���\�'�l;LQ����N�}%.�]�_��ÞC;s����e��m8��8.W�o���F����	���:8��Mkڅ��k��[��1�¤��IYf���.��N$�tBu��;lP�dӑa-�x���]e��������5�7C�/8r-�ih����p߽ǓkSnG�N�VL��J��t�b�Z�̡+����%�2�l�J��Mm���ʋ�!J�n_o���Blp��nmSQ��95�<�!�/��h糖�r;��anV:�>�z�=Ϲ���\÷�U�묌p�Vر�L������׾z���J�il��dMj���}KJ������u�ܩ�Q�o�=���B��+������ң��r��>��^UOϵ���[������F\��^��g��3֊�ڎe>�W������`�<�vx�=�&��py1K�\�۝��<;����:Rۥz]��߳zϷ�!�g@^
��5y]���~�2c���8�2'�9q/gn3�W�y�Z��ڗv�����y���<7��ީu���h������E�I�'_����\�y~W�֡J��w|v�������+��z=	S.�
1/7A���|�3_	��/���jP��eL�����kW�u��{����r�L����v|�v��3-�:m�)a��n�A��\�62��sNI�.}V�O����'�;�hP���}Q�'�v�{��'���ʦ���XΡ�}'�|��n����gٻ��xN�kšA^�s�O
b�f�]�F{�Ӎ9���E�X�x�朦�Gx�j��W3~�95�p{��d�fwk�W��mU���\rk�)��g��6*q����g�^34�[���;�OM���tR���Lt9�9r���+��&���ʌ��UV�9�x�bw�:ʝ�~ކ�Jy��uYCI8�+k켘k�c3@�tzQ~�Z|������j;x[�X����w�؝dE�{lS�.��U<��b�y�}f����煹�i���z�DoS��X^K� �)vn�#�����e���N�)>��1t�;ӣ���ܶ�֒�%�۬k�ќ�؎^+/7����-�Tkkc�Ir��ɵ2`��&W�Z����Zeօ2��c�O`��)fN��޹���"o���6o�����4�K�gۑg#�����:���5����U�t+^��6���Y�t� ��y ��ڳ��W&��&�I�����O���P[��
�i��4ϔ�G��ғO/LqD�ؘ�aW�W��+:�g8fo�sL�r�z§7��^��^�w�/��$؅d�s�N$�La���C��Y���l;5b�ԓ}f@�%x��ud��	�!��m }�����=�����\�\�����l��r��d�N�6��,j��%�=��Hq���7��q�LXbz�o��3�2|�߮��N����L��������~G�Rp`v�2i���M��VϨm����՝�q�-n�,��zԓ��E��Ci�׷��]�ݽ{��o\ε�M;`i�i�_a�6ΐ��읲m&�{>��M�O�6�+0���M���޲C�<LC��d
��w
���^Ľ]��P�Y������܇Z�P�/Zkg0���z��|GJr˥���ܝ�@����γ0���L�E��T�|�V��5�6�gBsel鹬�����l���NK�?c�!ϩ8͡8�L�����w����`|�'A�0q''HOMXs�$�u�$��y����t�������>`m'�Hp�$;p<����3L"���{��N�$ҲN�y��&�d�	�->5a;d�5�����_����8?��?b�~?N2�{��a��d�2M��E^�z�Ԇ��,��t���:�|��Y6�I��M�r��7�3K�{��s�y���l�Zs��C�<v�v���L2o��$��]Y;d�|XN�0�I��I�Qd���[z�޷�/{��y��Z䞲N�{d�'�����q�i��!�L�;x�7>�<g��F��`����I�{�)�{`c'Ȱ����>9�{�\��Rszz��K�����+��ǟ|�����i!ú`m'oL�����z����3l�O5���Xu��6�>�k�g_w����k�lY=T"�zɴXs(�0�u$���7�|�i����i�g�6�|�$4�|��>�>w�z��w��U��/Ĝg_�HS�}�hV�� ��d�C���v�ՠ|��N������<I4�w�I�'��I�=O�a9���}�ﯽ�[柹
��<溓�<d<5Bm
ɇ{�E�q�ɶ��H��Rwht�K�Bi��߸N� �d:g��m3��~s�o5޵�5�4�1�2x�8sy�@�Yd���}�d�u��M�����O2�Ԛd��`;�����}���<��t���N���4��Xh,�p<f�O�i����M��PZO]�n�&���7��1����S�|�ꮫD*Am�"���`���?+��v�-hF���*�.+����^��:��yNᏎ���1��g4Z{6>��$�<�g�� P�<8�^Xc&�!��I�LE�u��@P�v9d�a�Y=a6�2���N$�=���9�����7�}k�bϨO�9Agl���d2�d�!Y�P� Ұ�&�`kVCl��h���*f�=
���Y2�g]unW�.1ۜ�=3�]��?$�ṕ�M��4�+;:�i��'a�04�,�N���mI��m��C5�
����5�u�}�߽]��w�{���Ç~}�XM2w�):~I:��v�׶`s�Cl'���Ć�t�Ld�=}�E&�=��IPs����_��g~������~� q&0���d��7��C��<g�M'a������3�d�П2VM*��;I�M��lּ�6_��s}�w��!S�V�b��i��v����6sY�����{�x�E��<��2O뾲M�k����O�y����d���<~����G�O�6�}a���T8���N��Xd�9�'�����(N00���!�T'�c'<:��ow�<�s��c&�{�z�I�ԟ2q��OXm����ЇL�6�v����N�!=��$�D|��Y �$|4���k����7���~k��Re@+''5��=I���M�O���&�7l��	�m�2`m2j�o<g�O~溒m����������|�W]}��'=,'i0+'�ü�=I�N��aֲM�$��'4��yCI0�8�손��!���e�w�O���I	�W��k�xsk
p�}��}��+�.`�G����û��_#@�m��IH���dr\u}Pu�x���˔����t,tD���ޗwq,wh�S��o.�m�h��'����|f�襁�w�Ԉ������{�i�|��O�L�q'��T��a6����'�d�����N�0;�Xi��'���/I��^f�ځ�$�4��Nr��C�s	=B���h{��"�Y���q�̠ii:�Y�>�Z�_#���~��徠��~Y�򥱭߷� i���@�NRa3�q	��k$��|7�@Xw�(�M��V)=I2ߐ=d�(@�L��C?N���yO;����x����@8��03,�$�6��d�:���!��d1��0��hVN��Y7E��a=֞���y�5�i޳�p��2m��I�C�;Nˬ���O�C�CL��Y'�6�@�$�s��6�쾯�#�~��$SC�	�w����u��{��ˬ�^�����pwd�I͖-��,RWL�VM0=d��!�C���I�:�I�C�I�2e�4��� ��ŝܬ�)�f9�?c�������9>�@�a����}E�I�	�`z��d��S;��$:�i$��LBq� )ïy[�:�������*,�[$�	�7��i�-�A�� T.褜d�)1�$�Н3�N��C�IY�쐼��q��������{�������k{u�O�1^w�$�8ΐ��Ͱ9l�F����d�s|�HT6����'�V�M�FP�!�N�Rl9�^s�u�:���{�y��d<a9�;C�O�P<I�&���4�2�1�a�M�!�d�x��k VJ�X�`f�;g�M�Z�Y������Lp7��ki�˼ ��PN���AC.%���c����cx07hJ��ۂR�؍�{�:�V�ӝ��@�b��fRǗ�|�T�02�êYs���]e����<9C��I����*M���z�������}�O�}�����I�Y=�$�'�XO8�j�ޘ�8ä�!�7��I��s	�{�xo7�Z������	�Ol$=B�0�O�@���4�I�(m�ć�=@�'-4�v������0�I��C�}�~�u�k<�_��rI�+k��I�h��=C�Cl�d��,�ԝ�ɴRO|�$�'-��I�04�j�i!�ߞ�=�]]��oZ�V�f9��p��+y)�)�exW9�hcY�<gG�R�0���:d�'s)�m���Bu����>|d�&���~;_LϽ�sz��nԞ='hM08�rÌ��:��z�oWI����|�=N�C��'�4��>I�N�|�&��ٽ���t�h>����~�����ߐ��ô���P��;x���L�	�MOl��M}�	�
��T�0�Y<E�I>I�K�o���k���������'�k2I�Y�&�M���$����<g�X0��4�$2|��?{�@P��ȫ$����w4>��~Ϲ���d�"��'��@��Nw̄�C��t�a6�uI=`a�d�g��}��{fК@��Y'�vɌ7����~���o��'�*�b�@��Om$�/�2}l��$�N��o�M0;���Cl:���l�Y�������I��:�㯼�<��k���ā��rd�LE��hVOf���6ãv)>k	X0��'s�M0=I���I����??��o�����Q�뷘z���_���GN����='���FR����<�dݷIR���N��w�5���~�H����iBG�6Ja�*��ÜR�rT�
�ָ�(���}��k�~�c
���'7C>E��ԚI��î��6�X]��$��M����']Ye��'̇���X���-*ɋ��ǘ� ��Q���@S<��Y&����&�`kT&�-����+�,'<Ջ��}��2k�߳�������j2JϏ>�C9N�z��N������I����j�0��rН�����hvn����q��o}�����=ߜֻ���\O�XN��M��@󯰆Нj��� ��2O8�H�$�$�g�d��r�`m���d8ô�>ѳ]�r��y��u���+��km'��	��d�8�:a�RBy�>E�����I�w9Bx���|?Z����vz��n��y߷fo�o��B��	�t클��!�{�Cǣ�(M�3T�3��Bx�`u/�d��J�0�xN2mN�i&�9i�_tz��=�~r�	�N�4�v�\���L�=��a�9�x�9߹!���!�<�!�2t�@>I�|�6�I��fz�~̓��zzS���b_��|��NZw��2}g�O�vd�!�ߚ�I�1�z�$�u��C��ua�$���I/zc��{�y���7����I�Ny�:��I�$�;Bq���l��i��y�=x�>3�Ck>d�����i�z��C�����7�;�u��}ߜ�k�5�2m�CĜI�a���_{�Y�����oG�L���I��uͬ▫��M���e�4��!Δ���w�4���;�����os5���avز�%�.�[f�u땆>��,�D��X�ꃷ3#�͔'>�^��v�j�mtI�꾯��o޷<T?��}�j�x�D������*�9u�Sgr�2���,�c����F��N�l󢈣��f�������~�������ƥ${�l%o!~�}�+�ӵz���<���[/k���z��cJO�����^�q���8rOu'���ӾA))*�BJɮ���a��${Խ4�s��6�V/�6���T̘�꼐ٗx����Ã�Ga{���gd����u^Q�/*8������у�!'��?Qb�?�N�I�?���3�^���ؙ0S�ܾS��ϯ8��S�ڸp�����Zy�J|�͡I�_�GA�L�;F���/�O�~t�)�g,��C�i��m63hi;s�-H�;��T�/y���	u���5.�{��m1[G�ˤ=u3��a%W��=��E8�u,�+n�J�@͇�.W�j+#Z�m�ƩrB�`��V0E�V�4HB�$��Fܧ���E0s^��7�f!mv���֦Fxj�&�pc::�njOlpmZ������ͫ�7k�ݻ3bU�@5����qMⓨ<��_>��o#v�$h�Y��biՑ)Iם[�*$m���/;���a*���&n�(��8�r�{zzh!�|����������OH+4m������j�����8��C
B��ٺ��)rg�Y6�qw��z�i�軽��D�1Z 
�a�MYn�3%Ji��2�7܄�����&����h	� ��WsVm�޼g��vwc�Ku.�=rZjR�V�؊'�;F���+�vJ�c��JY��Xw�k!��׈Ia��-J#egd�E��/�n�Q.�5"�������[�-P6GT�.�9[����YA�i]EuFU�3s+l�[Sk0�R�+�����m�P�bƩ 7f�[�梵�׳%d��2i���?s%��T��K���\B�U�*��&�ʹ}D�������}c��h�}�+L
�&�:�*�oUJvl$t�5�|e�aU�Idg�в����{a�vȅg׊<$P�$��cvMZ�.�� 
1u/%o1v%FEv���7�\�4�W�))�r���KiR�=��QVn���c��݉H
%�*˂�&��s��ˡa������p� -���#j�n6�m}�����:�}�D�8t^�Jdm��C��	�q��>X��v�ɢ��nn�X�"q�A
1�vE+����m�b�]DQ�+X�յ�����	�#��ܔ
*�u�`��#����
B�J�^��M��On䣲Z=`Q��`\����Cy���glHRI���J�7�еCVvC�4i!"�Q�9P`A�<�ȵ�ι�x�b�����ݤ�K\�;z����yRWd8��ˤ�n�#����%qn�)�k�n���*�����'K��C!N�A�O`ڽ�;BN��+5֒�L��':0���f���/4>��'���|k�&<�gXJ��sl.�q�c7p[y������M����w�?����]A� ��c�K-FQ��Q�Tm�╭���	2�)U�Qb��J�2���ش����)s0ȃ-*�L�2f\Lfe3!J�*�ks&eImm��f8#m�J�TTƢ�e��YZR����`�����UT�\C3pm��F��DU���&��Ŷ��լ�����.e)��,��1kUb�[Yb5�Z�F�ɑ�`��l��"�h4-UnZ�j�m-��fR���DPLj&[�*bT˘Tp�\���\�V ��3nY��Z�\����-�f[LqV�ʵ��%���"�F#ZX�-���Q�-�[F���[�0mU�E�jԭ��\pTZ�YJֆZ���fW3-��j��b,b���*8�rLE\p�Y��r̹\�LL2�-E�V"�l�0̢Z��ە�r��Uq��e��z��Y��[�-fQJ���-oN����!����fD�o\n\!M�,<'���;�I�}U�ٱ�����4k��x�D7��O�O�;�{���~B�R�y�ի��
���~ĩ��T��Ϧ�{�v���{�����:fYr)K�����<�r�����MJ�7�{��ϷB���V51_/J����\��S_L��}s{ڷ�s����$W"7E�p��{�g��f����įDf������b�a|�Ћ��:����!����=^*n�~��٦� }G{�o�6����Ӣ��~��
e�<���_[��e.�zEy����������W����,ϕ�=��%��x�����U��
�S*	i��J�5�]s>��|����}'���R{��竆�,�=y[xǚ,�� ����c����U�xm�j�D�tn4U`�C^vRE����vwpm�6t�펒݄FlK&V�C�a���8�6Q[��-�odC7Y������??x�%y�f�}��k֍0��ε�(н��`C�Q��䃁�{_����LJ��z���9O��8��M��ܨ1A���|b��Q��Z�C5)X��ꂖ&��n{T~>�ªp�|�KQ�>�������~�]Vg�Tw�fE۫�3��˞ꃗ.C;�6�g�B\�֮~�\��l�������m!�0��׸6L�"p/(��X`�����ˌVt5�zsDH�Am=���c��Sfi�k���yʕhG2˒������ф�M�My���ϔru.9�r^�pU�4������M�����7�\�������Rk(�y�6���������`2�Ď��}����@�Lo&V�!Y4[::no	�4ң��T��!N��9]؋�]×Fb�L�t�Rd�����\OiB�����7�Sʈ�4ڗ���YQXQ��F������~k�=�oKS�Z%�c�^�N��Ƣ?DWnl=C��=�:�z��_�j{3�}�Ut�GD��n��s�{�ܓ��Fk�W^�<n���p��m�+�u��7�m����m����1��Wz��(^��[P?^���jI�̞������3A1N���KL�A<�jW�gOSj`�&�d@�*t��|���j�wJ�c�;S�lw���kڻ��	h�3����я��=���Õ�Ȍñ�Z5�̪��$Ϟ�V�u��ɣޗj\�W]����{�u�:����mؙ�W��ut��{bfԸ����d��}y㒼��21�Y����v�$����O�%�H��3��ެ����Q�������%��)U��WUk�ot�T�B�9��#Vo����,��ݥ���Ӄ�l�&���fg-3�v'S��R�_~�����{ͼ�֍S���:��M};'�a/hvx�̥rT�6���'��7��_�:�7&_��yּ:�B����n	y=�^�:�����>ٴ�ϟ{+[��{�w��g>2Mc�,D��͡n����<�v�=���v�Ȥ�����xY�����ޕ4y�g\����J���>;ރܓ��1��-Æ��� v	oXԀ.�ezui",�&�����۹!�J��G����G{3Z�s������l{ޡ��ό�>�]eyK��cN�֧a3������c/�亅_���Y(JtX�m}Z	Ó&o���syڛ������Y�fG���'wI��R���t�:l�61t�bd����ӳ<�$hE�r�)4^�o(��R�0[�A�bT��_>ݽ����lw�(����S�@�h�kN�U)����غ�K��޽Z����؛���_}T����2�X�r�����5�6v������^�ᱽ���og�)͗K`ۈ�a���j�ܩ����<��R�};e0e2�i��*�J�G�sݿ+�֪:D?eLS�{[��)�+�T.`�f�����@������7�O{}=�ߟt�@L���S7��K�ߚ�=�����k�����'Bg�hy%�sf��ǔ\��3W9Vè��Վ=.g=�R���A�6��C�_:��zƕ�$����nA���Ck�]b�=�.�rr��fiMʧ���S��7����7�k���[av�ky9����^�L}◶��\yDʎ:_N�g���ٺ��;���M���/� �����L�ʶ�� �%Ї�^�}]�s�g�N�$
�Qluʊ]���Lɕ��4��]��dJ�k��;+b�Ѓ�=�Hq��
�6�*o�oc�?���^�q��1��붫o�oת�r������ڧNI��=�<���?g��>?��V�ۅf.�^|����琼�,e�ߴw���Q�g��A����v���7�:���%L��ށG0�ǹ��Ã	��e]뜨_P�'��/hYν1��&���6��C_&*�Vu����n�_�잨�1��l�8��F8|������v:��;���zM՝�yo�����(���1ٝ�k��J�{϶�d����-t��t?h�ž��٥a@����c�Q�����WWI�~�2{<�Qd����-E�{��u����XХ��I~ކ�z!t����`raeb�xf�>堟Y4���vW��5#�����^�α\ˡ�R��R0ŏэ*��\�=.�EQEǺ#+��7s�`j�43[j.Xڎ���]ٙ�'{�:��uE��"��?���U}l�S&\$�����w��#n�
��$�c�.1YЕ\��	��Uޅ�^�<�ӟ*�F՗%oq�5���틯x�ُ�M<~�O�Tn�#u�Yu���7���ѹ=�=��kv6kڛ�ٙ/m�6n��rb'�kW�ʞ��?q��o��i{�R���,��.CO��q,��u���Ы�yi��U�1�7����!p\���gF��Oؠ��c�<R��`�����ʍ���߭�w�#>1�i��O

Y���JW}h3��*g3f�1٨��el}��LW�l�|�	�v8s���U8�e��6��q�c�A�V��-�̚�I��5<|о�·���f��?|�,�Ǣ�;ͥj���!L�����"��K�9c�FNW'�(\�J�n�㭇�vf�3ծ �nh3k_١-wWY6�k!���a���Zpm�J�g�C�3g���/��-'(��ե�����T:c��}��g~s�\�[ý_�3�[�����=\�k��j���_5y]�֦b�rB������ݾ45��h,�R�0����M��N�|f�9���mP���s�=Μ����t���j�!<�b���pO*�4�����EƜ��^N����-��P�r߼g\���u�����)�w�Z��'7x�<J�|�������xҫgw��3�EK~�	�����=���Kv;z�d��Wwe�K;�O/�I�����}�*��Vŕ�[>����4��R�Kٯ��3"Q�$�|��P�)[a���ϳʏ���>Ì�*Nt��X����>8���^��u6|K�}f�J�ԛ�2�J�z#�tU������g1��-ku�,�u���6��U�#��Z���nH5�o�2=;���U}X[��<f����i���O����q!�P|����&\�[��2��A�Ԫ�G^������*k4�tƛ����x��WL7�wT.U륎����khUp�x�z�;��(��;=�H�OpM����
j<5������2e��{d�1�l�;a�hY�^���t����%e˯�E�������
+�7.�W���A�MU��v��5�Jj�{��w�EW��``7|��S�_G��=���챜��Uq[~}=O��.��~)8��&VM]��NЬ�4�g��_{����_Ac:��|��r�~�&_q��>�[�m��y4t�w�,�̮�?9�l�;X�~��Yy=��U������ �Hm++EDt��`,�?��qN��' ha�~�۪5#y�v�wVըc��4s9���+��&�>�\ޕ�������vI���E���l�\W��9���W��|�����Oo��:��Ǡ����<���/G&E��.n���[ڟkA�����^��aWC�2s�Yӂ8��^�#4��&>���ʍ^S}���Ŧ�V�j�s���Y�RF�fǷ\s���>\`q�Z��*C��s�����/~�L��'�C[�m�� ���b���]������^ۑR��TE�t�7�t��@���ＹNW���όߋ(-ݰ�`�B��w�</��%6�}��'�`�3�n��:6>�c9��1�bJnA��	.C�.J(x=�+�,++:׌�^���QS���j���4v|[�-G�΁����S�@#�~�e��z�C[�EF�^�
�G|ɮ���Uu���Хm^w9j�^ki�eRz�!�ӫu�ҼW 3W}ԦK�J�H`���i�]�c�F�ħ���Py/@]u4�9]���a�%�^`_
��b�X{�`q�Y*	�j�c�f=��,��WEc`*By�ѽ_k֎���
��-P ��=���V^HX]�Z��0�arى�[@5R;���ҵK��N��f
O�y��P��.|9���}��\�KZ5��+'\����F��.b޾2�r;S"�N�hv}�J�h���]K-�_=�R��E;�D�+�Σ6����$��'�ǻ+z{��fGO8!=��U��k}Ht����n�R�f��E�e�zMhB5�q��n��n�u$������q�H1�}�#�~X����2�:Ѕ�l�z�,v�q�W@�L�j����VB�r�M'yٔ��(�a�ɶ��L��d�\��`_u�ka�uI�ݡ����3��%]7�.`����Y�M�YlǗ�Ֆ�ɑ<��J"b�0��E;d}a��Zd����6�WbBλQl27���2���e�ST6�ot!�)��rʴ�ve%v�B�������->�XG�%T,��{+w!������m�Dih�B�48��_ׇC��:JóČ�[�J��Wk>���H4�V���6���ZR�!'��`&�V�X���U�Ltͩwat��z��iИ�v��MhTv���i��fZ�2��p�>�|���6*�˱yiT�[/I!BD%e`e�#[�pF��+2A ���hչk0�-R�v��d�*˷iv����6��O���B�*<y{]�V�2��2��3yp$���b���[lX8�=Q�i��b�*ԯ,�
�����ԝ�h<I岭��-c뼺^[Q�a�V���:�S��a�f����A��{8��j�R��c��y�[ڞ���H��}u�f���Ϋ��0�}#�j�Gp��s���ɳNh����r�g7F�>̑��:l�����X�[��*,�L䅗da�`.rޜK�r;X�ZL��"L�u���x^�kl�3+[KC�c-�*TT���3��B�Ī��*+��e�X6���q+���˕p��a��Rڪ,A��%[QR�%����3�F9lĹJ8�h�Y��(Z�����V72��Ib��UƢ�b�TƊVZܴe�q̮&ekeJ�3nU��9�Dip��ʨ�-i\k�U�p�2�R�2�d-�1b�\��kZf\��l�lR��Z��\0nd�S,��r�`�bEVQ\�T\e��iQ�" ��k�e�`�1̶Ũ"�*�Ppˌ[����QѴ��Ƞ(c�1�X5+\�S.&"�i��n8.[B����\V�s[q�������JɎ65��BٙE���F��	mAF�\��kQ2�6��)Gj\�.\Y�W30��`���cb-�EFZڵDR�kC���o�zݾ�z�]�8���nҢ6����M|��]Ko�}&nk�t�e�<����l���>���g���%�����W��boC��gY~�T�v�zwvIx� U*Z�=�ws��k�R2�Z�a���9%'~~���`��^C��t.�̚'���Js8�Y��j~�:;҉+��ޯjp��::.d�ބ��U����l��yQ�\���دy���U��PȫQ>�;��%!&���3���O����A>�$�ϥ�����?y�	���W��i��S㑻�)�޽���^V��'������<���~�b���[�����u���8���� s=jJ�]*�s�gog܅k��^!&ȧ�K{,���q������<�o�BE<�!צ�Et��.(�z���rAW3D꽽E��V��U��hfʪ"̸.̷/�2��9g����&N��vj\.SZb,ҫ�cF�=�/�m�ړ!0��w]��a�w`��Y`�C�u������j��Ζ��s8��Y���7�����������Gݥ�n3��؟�����N�����{U;���t5d%��5�H�mb�%C)]���xI�]���$9'��=~�v�%�&�y��1ќ�[<v{`qߟ���pj�v��ء�ɩ!���a>뮭��{X���}ab�Ya�����������Y"��~�&>-;B�Oc�®ƴ+�صV�h{�'P,o���h�#(Iد�ɖ���L��U��l�ݗű���NxfJ��	%��N��}�Ó�f�u�}Q1�������-V��w�������	dpn��/TP�����c����-���T��^��W7��v�Nv�c6�䞅��}�*���Tu[�+���@jo�0W_�f��_��=���O�rJ��rr����}U�Uo8�<'���̶sޥ��Td��}�4��x�q�R����s�Of��]�y&(�b��k��&���w���ӏ��� z� �t<��o����-r�؛��o���״��3G�N2�D�yͺџ��ޫڬ>��c�[�͟Wm
/N�6IO^}��J]l�>���T�Q�ӫ�����:�]qՇf�/����_Mf�c����/�.]gg{�7�My�ڀ�_^�,t(��m�Y���K���o�޿g����
�=ڴ�,VwɂPxPZ6&���U�X�g��p�����^���u	`Y�R����N�L)�G���F��X�Z��*���ٝ����w\���-��3)�6�H�p�p��Kow���[���֏�|�^^��s��ٳI�Qt0mCG/WD@�붛��;�%E�n�W3X�k���O`�������J~��� =�|Է�_��0�w8��N2h<(m�Z��V������Wp�א���^��J�4���Q��<���#%fd��[�t����K���*>�.���-/^��<�R�����ܥ]&Qn���k[�j7!y�S��v_�{�Z�������΅�c�wx��}|���xD-�����<���ʛ��E0���1��>~��W������)&�1�ʑ�t��q5�f��G�3٭鴯ܷ��7?>)ƪ,V㮫ʞ=�]���$ƞ9�oJ�= �x�a٠�H��۷Ќugg%ps�l~���w^��5g�ζ�WXc�מn�.�p׳c�Ԝ������|��<���<��p�5������C*e�Ү�h�4�G^{��'Z4�C%���A�:�-���E���P�`U��+�@��e�;�M��w�qZ<�)������}�=�m�7<}�<l.Ϳ�K;t��:zגl��t~���?W��@ԯm-{V�kmS��SM�_
]�����n���[K�,-+8���u���7!��}Xy�z��`��X�m�n減^�s�����ݞ���T#'����z�j�'��J��p^z�9cuh�#Ź��J�T$��8$9���{s��ڝ���f��u���E���L�viQ�w�#�bg'�-����I{�y�Vq��%�yz�.xէ���c���ُjGr���$�z/��t=��4�߹��M��q�ޏ��}�>A�^��ZŞ�ꇹ���C���&��ig8aȯyoX�9�T3��lde�r���ف����fm`"j���"�C����
/�ը̌�
�2m�v�hSҎ�ø�d�ҒI�M�l����gT�A���A�E�Jqn�w.K)���]%G��?}UUU�w�~�m����jѨ�f~��3�D|Z~�f����/ѝ�X��'�s�����{�︮)2,��	��J�{�緳��2t�G�3%����u��{�my}h��Ή7̥�꺺���*��^Z��L��Xl��_���<�a�g�#�c[��/>��F�\�ney�;�}�x�Kv�VE��B&�-m�l�4����� q�C���w�ҽ�Ө<~�~�qt�/u�u��b���=6N��k���~��5[�|��d�xMx'm�v��e�%22�C�J���X����@��Ukhe[�w��o����/Q$^�Șޛ���D=h3C���xF�~�f%�!�>�[�X��+�>^��G�SG�e�y�����5=~��~c�a����D�X��Gw��9w��D��D���?����T��c����]����i�m,*�Z*��"/����
�i��xV��軑G$��t:���X:�s(7*�8g!gG�g����5��͡7y��ߙ�'����,��.(4:VE'm��"`Ad5�aճs�o��j�Վ�\u^8��x� ��c����uN�y9�ܩ�����9��9�?YB��-eC}q���x�1-"���Zz�z��M�Y����$�Y�h��B�<ur�(
#(*F����ϹD��J��)�>����l���&�z��~y2��'S7�\U�x�G�
N�TǆR�j��̢{����:adxoP�P�t���y�����ap$����V͢:���-���N�4}c���ylB������]j�Q�<�^�G@[8LR�=���+�8�/�pU���%�C�5R�o�|�4��k��^C���m�p�6m�½I���z��t��f�����㑈��<��]Y�^��@�彽�gτX1"P��`$��ɔ�{0*��)B(�|���PkJ��c�0��/Ey��vbf��z�� ��W��-���q��4�S�"�P�*,n�Ѓ�Ԗ�^+��y�I���{�^V�7=�ۢ3� �8WlWR���B�������a���w���������O�~,��Bu~*�1V4��ߪ�+T�+��ȯ��A�*�O�����m�g��b�Z4�x=и"�ҩu�<�Vı0��5��tZ�\��׈��w���),Ĩ>5\�E�,?V�x�f��w�Xۮ����j40��[ ���E��ʱRS4r�-gӍ����g�U·���F�ç�aܺ=L��&3ڨ>S%vЃ�����*��{�����e҅��
��|�ؕ��u���=��_ǟ��R��r�gT��ՉP덆B�v�(�<���N�TJ{����M��M�8�x����m���<��0�L$t�}lW٭e�ȼ �q�:BoVg�ux��#��nX�2�F���+&[@a7�"�ŵi����6n�Rƕ�R�Ã��7�jY줕��[�7�Z/�N�
�G������n��G���W=�O���W��1���ض�o��zT�Y�B,����c��V	L�@��L���B��*�?UzO_���+t��C�XY��}x�O���Y3�p��o����c�(Y�����*�P���>�?1j�x4h,SЬ����ՏTX�N]�?����ά&|yx:3���,R%�V��������)���=������AB]�*ZE�J�m���/�6<Y�>��#�/.X�#���MAy+u)U�੼t�B��+&�#g�u<�W�*��w�/5��z�������A�*�i��S����3LRkJ�󺻥;�w�����3S:<�*r�4���ʄ6T4�B��
�%�J�m�J^��K�z�qFT�(н��B��m�ag�C�P��%a�(��a?<JT��f��e�>B�YUJ�nU�ѵ�]��#Y�'�X�YN$������7��{���7M� �f7����H���v�ϧ�vr)�Q�n�S�j`��9���h����nq앵f:Zlɥv*=l����QN~�����eG��V(�;3���*����,�JG�/�6�Hxe	������<ײo}�2�¶���F�ʥ�<;�xhߍcKh}�wj��l�=�U���t�=զ,��/�P����
�,����
xpu�K���]���|�=u�������l7�8�:�lJ뱥�ev���/=�K��xϒ�f�b�[�F���+�K���l�,r��k��g�o���JrA��?1��1`ډh�s˃��ċ4���:Ϭ���wּ�S�}�zm�g$�PE�tJb�mq�TΊ������Gּ~�q,R���M�ߓ"Y�ʁ���y}�B	c*���k5q�n�(v��0��sQ�3�����P"��g>���4ʰ�8~ӺQ!Ԋ������gs�~�ʠ��G��.�y}��Oct�s�=|�If�ajZ>��jm�8�o�[x����- ��1	��:O%IT���m.[ٗ��舫S�����n�M�#�T1b�n�����[�B��_h��m�olS�O�����m��h�-�<C{vKA��~|�:�r�u�޵}s�NH�b�o���KlK�7��dm�ƥ�O��\/��2&�l�B� "&.�:촕���G���t)����C�s�	�'ûtBP�S�yul�#5��x��r��w���
��c��嗫��a&��YW���iۨ���Ѷ���}8�9V8Gwe+P�<��qV�$U�#�_WgG���q��l4��r�N��Z��u�j���cO:/�����t��  -Yw���8fn��z�4$���6����n�إB�"�����u��֒_���
�7Ch
)����7���ɼ�u�
ۀ+r�U�f�Z�N*�n�~\O=L�V�Wϋ���}j�C���k6L[*�J6N��r��˫Z�lڒ<��P78ϧ��=�,�f�@��S��v�NvvN��vED�Wv^*���O^�oE�V�(���:9�hJ���[���HKe#'��
��E.�F��Fyi�!َ��נs�5��&p�}�q�Z�Y }�*��L��-���Վ�\pȃ��%���{B�[5��)ؙ�pŰ�iK��`�J���[
�R\�i�Ҟ�#w��S��nIU5=M�oe���͞�p'�%ږ�F�S����I+s�h��iq<��f9yj�b \����;�`����b�ϓ��m�ڷ���N�W)4���GG���x�q��KU!����pJy����+��|Af�J�ܗ��ӹQ�it0�Foa
�`�Wv�ϖ*-	h����n]�uoCHU�#�NLO��K	!`�ޒg��g���KYYt%�l۝����f�_�i���@�3G@xA�:7kt��WHi��K`r�/m:��%}���C!ɗ�hm�i��$���bqsg#��*A�(�iF���YU}�-��[KzM��nG�JԪ�Vema����I�L\�|BoaO>1�h�FѨ{V̝����.��Ìuv5Fnml<NwThYw[�qΔ��S�3�v�d$�a萷/z.��2�h5-Z,̅V
���"��R�h*�"�d��%¥��7�V��r��9U�����AKiR�2��bT)��3710�s&a�mS3Uq�*�n"aUs���4Bʡ��ۘ�G&�U�Z�jf\W-q30m����B��p-*Z�Z6c�[X*���*Ym�q�d�-+(.)���i���2�e��\nZ51Z�[UTq���a��Ja���ɉ�.dq��9�ѣ�W,�L�s1���2.%��ˌˎeQ�n3,�̴2�+�[h�.f+��ne���92���lnf8R�LfZP��J8�ap�R�X�JR�f\ks2Ֆ��j�K��WJ#J墔̕s��8fZ��0�W*Z�rb"��Ul��e�J��5m��őAF��1�ecm�rւ(�-,��je�B�9����)��)\A��4WS9��\.R���L��[r�ke��F�ƙmeT�2	F�۔�̶�(�թ*�q0r��W#S&b>4I�@J��yR��;A�3�W[��E�[�N=Ƕv��8�%A���[�kWw�\A���j*����/��+^Y;K�U�/�Xe�2�����P�`��Q��['��/Oo�����]WE
D�:oC�X�g>�ʼ�+jm��d$��d��i��(��4WyrR��l0�THx�]W�
�(��O%��;��& e�d�n먫���������^.�Q�+��Fܙ2�ͮ�﫺�M	�Q2.(���Q�eN�WG�D_z����r�e�Ҷ;��eZ���Z�����OO�@uKT\PȰÆ}�Y�	��W��T�x	qY�SP�N��Ҭ���#Y��<p�W��(��,yo���z�KN%��Ŧ�`�E	5���X;hK���tW�(nd��n�xz����?YT�е���|/��w�%cP�ܴ�uH;gy��j�G�L��1qd=$]k�W(�
��.y`u5x�6T9�Ո橖kԃ<��+~^��T*�n���Q�
x�D����M��f�W:�g4������zf�����6qe�q�I�R(d-��:�=���ԥ�~3�X�t�E�,�Kx-&N�p4��'���ꪮ�<ؔ6$�h6o�7�ڵ^�3�L�H/('A�g�B�X�����)A�x��:g+�zP��Et���y�����a�ND��EZ;��]n��D��G��ג�mg��U2k�J��ߗ����C�J��b�]־��?p�1`�|�>^[>	$��B�T����uea�eK��M�y=��%;Equ$����yh���ƿ�`�D>U����uͫ>���l�\� l
�d�A�ZY��Q�0y3MB��y]��9����]��*|�Ei�7�A�i�eX�*ƃ^C��]N��~�D;�^b߻:\�����R�O��,�\gq�iJ<�a�Zl%g��,3zf�/�,���*��TX��Tؑf%�>5\�Ea��v��܌GU��jKƷ���2�4/��0�b��_:�V*ܶlء�T�X0Z�'��S^�s�,��GGi�Z����M�9�9���.M\����A�M�fC��V�PW������X��:���gvY$n�����Y�^���t�c(`׼���.}�{3�
(n"���U}��Y��{�+�tl*!_z�8�#��:��IQq�ʃ��f1#盵<��N�k�H>B�C��~���Z�<7�����.��N���g��e3�*b�ج[��Pb�;o�EChU�|�05垾WY%��>R��z�*���Ea���
ڬU\�оҺ�Ge:�{��|/پ�����(K͸}��-��3�SU�늱%��(!�nX����������A�j���� D��n׃���Aܿ�#(���f��2"��C(x������s���(`��C���ϻ�����}��Wp�y7
Q��Շ�&P�+I奥��Ccx:�Y�!��Gs�`��W���^��	�E����C+�zpWS8"��K�f�����sΫR<\��@�!W�B���j�+څ�DY䆌��OU�;��ʽ�%���8u��g������@t�%���N����O:�j:������gEr�J��be�y��V�e�{#�S��B�]A���#��kdr�5͵�����~����mks��Q�6��_y��P�i��l�j��IѤ,GOmEW��nטŌh�%��K�W�<�0#J���>�"��f��t�(��T�!w;/C��h�E��(պ�a�ޡL+~�E0��'
V$���#p�����gw&�ƚHИj:f��a!f��[�b�ǄA���?:�/��i�!K��t�U�r ����>�~7ʘ"��.C},u����e�]������#���G���J��,=�Q�,�$�Ŭ��r�)�=^3�P���C�rVo��7�M����t+V+���nz�$<�4�c�3�h��Yp��-c��=�^:#�o:��v<f�N��"r�l�����Tb\t܂�\�F��侕+�:��l�(j���	�)���p��T���}��|4��,��L��M/G���Q���x��v���	+.�t�_a|��S�vʹcJ�x2��=��ce�,�J��H쩩����˽���bGeFƱn$��)傎�=ɼI��X��;S3O7����J;K<ܟ�����'��H^�}���������[\b\T\\��>��៽���3����J�9�-6�#�P83~���#? ���.b�v}ͮoR�hc���M���+,TI�Y뗑�ڷr�WK �����$��-4���t����5�!����g��N���Ԃ�L��{nƉwr���{x7�N�^)� LJ��<k�!@��e3O�jWH `���ڶ#�|W��`�b�T�����t�f��e����f��h�-�����T�k�B"�:i]1P�kTHa�Ap�X�x�(�N�v��e����*�"�H�8Ҋ�c�b0�Z؄�Ul���ޖ۷�����g�6�F������ux��h�����[�W+�3
�s���}c������E0!��T�FÕ����ڪtxf�z]H��́%�`�jŨ������cX�g�r��{Y̶���N�*�j��I�u^�;����1����AԤf+��M�ʥ<��.;7Q��+{��ȷ�m1Ҵ���I��W�U}U�)�1�o@I��"�=�LP��>#����|���+"ǻaI�.Y�1V�]�[$1�1�T�Er�b^4x��LBMb�|W�Ϻ��3:x����JfU���hᕲ�?��!�F.����xp��>�в���85~�d�5'���v�so�{
��:��,kN��34;�d嬞�=����2u��W�뢻�PK0iM3ƒ>�{��yo��/�:T�Y�z��B;���l__[/��Pΰ���`���}��f�x����wK���P������ֵz�f��dP�mu�GP�2�:wr�6�}��B�,`_ �-[<,F���i��m����56��0�����m2�����0���R�g>U/��_P6x�hxR��g+sk���o[i�6W���!u�F*�����E�r�_��O��6����C��NUkj�%n��+Y9%U��K��>�3	�_lU�*C�IXΫ�]���B�b��*ӜE���/rL��n�x�G�y��3����]�5�2�:�N{��gN��}UU�Vgn�&�=z���U�aPL�t�&���%f֡zr�f/" {r/.t���!BѥQԄM|�3}ƙ�(�֌<)i�3-���A�{[n��4�/�s.��*,r/}���K�vT5:�Gv��}���oY���l�f
�=}C�χ]��	_:*�_M�L{��-�^{�"^���^V*�#1����^9H`��X�=A�j+1�
�߷�bg<&)���K��R�P��
�����ؼ<+9sK��C�y�1��xqA_uǰJ�P�XV�w�a��_��E����oF{2j/\��N�M�>թ@7�������ǻi�a印�49S�n�(�_�73����".�҆����O�����jҘ����n>�벳�~c��ia!�]Qn��7�\z,�]�j��+Q�4��f��7yO7�S�`o��V�2S%d,/t�`���\��T\@]��1�3vgf�m�}�B��ٮ����3 �2�#��$Grsv��JeZ�0�l�="��F�}�� =~q��=����v֛�
V��0�;�aU��m�����&�h&Iz��H�t���-7�';�'�����-C�c�o:���*8_A�{�V�{�y���f���u�e��A\A�M�C��AvV���s>2��+c*��l�o0���<ZP�(��5Ɔ�pu
#o��A)Ghd�?_���1�js�E��q����aP�Z`�i���eX���<������緇������ť�ϼ�*�,l �P�f����m����L��(�	�+"�"���iF��S����L+����$��[�{S�>�<�=�QQ�4��>N&�? _���PbMG���O�˲�(xN���RF��=b�0V*u�,��S���4|�	�Yo�L���Z��B�7��\�3Ș_�j�i=�N�;�>[����P�����C����R����{�.�v�Q׭V͢5�Ԓ)����atc#.��̶4s�������&��x��]�zw-���X��գj�k�,(l���i��>����ﾪ���u�nK��?mV���S:�Zt�j,N��0yYU:���<%>�+|%�=5/s�z��AHō8X#ع�`�Eܸý�za��hJ�y�EV��_�0x,-�$���DH���+��r����r�ֱd�a�]��n�W'�H�bA����U������Qӣv)u'^_I޿vΔП,���M�V�qi��4�bej�%�9�JfT��)t�����q���ں�����4�U+��}�@�w�:�_x��U���c�4��<�����q[L�D&�XB��g-��Y[��#�$a�1�ʺ��NW�8ʉ	v��y�p��t���ȡ4]��}l�^�߰�s�{Y'���JT#X-�yR��d:r�$�^K�d�ɾ�xm�=S/�Lx�kU������\Q�_:h	�%�{���~��E[)[�"��Wv�k�'ʺ���N�nDwYpq��6�ZIV�Ĕ/ާU�k�Fk�(�}�r��X\�r�V&��JWv�[i����x�n���"�"�fs>w��3; S����G���o�;y�L�(��lv)����V�Hx�]@_�Wƌ<MV�q�y�R4X����WQBH��i�W�]P�+�}(mnW��^��x�{'OS�y]�����(��dQ.��8�oֈ��^,>�-]u���s������d�P���ê�8m�|p�iYaʆ�XY�9:qP�{��l-���5�%���"���<��_XȬ8z+��W�=���כ���{�N��K����U�f��rTBO|-y�KH����uK����d���W���f�t�0~F3N�Z=�t>>���H���ᕚ���{'���+��[��c�B׎�R�FPHޗ���>��Rd{m�2��%�
޾9�Pٰ��/;n�5�P	�4���'A�����W�Α[`�]�em��ȳe�=L��-�B��+G��#G��R�Q��{ښ�[��8�Coܕ*_p�B�R�vUc96���[zX3�m����N�rЩ�T�����%��!�4�]���'Łv�V�٬ �]��S26��}"֒����pս9˛�Kcc4���ms�vNՌ��x���|Og'��Ɗ�u�A��Z&���m�H�	�jF�R�����(J��Ggr\;��^�\��d�X�aY�&�J.�K��+��������U�ǚ�65�8���5o&�ug!"�,���k[¦g�Y��7�8n!C�)\�1*8@o�vc)�Ưiq�V�6;V���Fq�Z�v��A<�ߞf�r�ȭ&�n�޴{+���J�g�nb�
U��,I�M�֓�m�%P��oz��`���ږbع�S�u���/h\���=;� �M�U�=��43^Y��ܵv�*�/��AZV��Ըu�<�����Wc{-�8[7�RY����*<�aX��d��R�]�[o�91�pŖ�yvR�����ܶK{W��l̳ʚ5���ɧ��q�t>�e���aւ|�sgP͹6!�E�t��
��}
܍�؉�e2
��u�T �H�aT;�O�oS�PZqV**��?H��Y�1|H(��U��p���j�w�o{��v�k���i�vCf��3.͑wb�@��x_�.6V�:�����8_�� �̧B�ǁ[�5�����Vb��J���n���/an�F���C�O:���b�w�7t�[y�b���3��0��Բ���-�8n��]�Q���.��viY�n�ۮ��<�.�"d��诛<C�!��{�,v�`L�RT���ڴ�:��[U��͋+']�nd�3�c#��Ú�D�5V�g�W;]3K��B�m�FE�X�乱���hR׋�5���݈���e*{|��X�%]�M�X���Jc}΀��)�ݼ;�X�Aq��5�%�}�j̾�C"4�[P
4U�pǣ+�g {!�dE[���i�wu"N.X
���Af��<��Z���*�D[�h��K4����Xg��� 1P4y$$&��vn��ûD��0ؾ�L�
y����nK[� �upV{5^�>T��٣R��ٝ�f�q��ZBS�b�1㤺L}v�wQ�ԣxv�X �(^鮛T�t�|�q�*�o�5՛�7<ls=s���p�;��Jҋk�N���9N�ys�����^\q�26��KJ��չE�ams�*J�p*�V�UR�,��aV�9F�ZbS
[Je1�-�*9Dc�D̵U+r����\+TE�"��e\*�%��1DLa��[am���lK[`�Lr�-�1�ʹqȨ��r-k*X�(Z�[s(�c1.YYUP�\bZffP�E����)����ƶ#��eXҕ.YEC*�ʶ��9�-�[k�de
���P�bUK�j�q�b�R�Ee��*"%K\�9q�U�m���kPbU�Z�H�YiX�XQXQk�[�4Xm���L�p*K����V[P��c�Q0J����9B�K�6�amQ�kZ���VB�F�J�Ԩ�m�Ҫڪ��'�g�����u~���?Gֿ}�����@�t�L���<�â�+��U5Ieay5��9m��j����|³_I��0����@��a_b�x:���k���2��嶃�ٖt���L���_���}(+�2\>��-���X4<�P�������}�)c0_U�,7b% P�u.+O��IA/�,k5������0���=ޣZސt,����[@�b�<+��J�wP�������5s�	���<p�C��cP�L��L���)�f/^�%L�KY3�&`��5�\��HF���|�]l\	`G�F��y��yU���u��z�V�h���(D��p�����픈f$�1ɸ4�OFA����J?�V)���0�OW��>_5ҬV��j�X�|�c�"f�Ʒ�Z~CF��3
��<��Cëj�p#�.���x�:6�Ӽ5>�V!v�d�2��3�@��>d�C|��U��,zy�G�1��������OLT��N�Flޫ>������F�uO�Q�����p��f�CbK���l�z4PhY*�8N1JJw�����C��-7z�&�F���8�D��S��U���f����M�,+�-�m����z�谂����`�N��>E�X{���~���{+K6=�����)�׏�+��w[��h�9F��G36������H��W��Co��(nt�E�p���*��fI��g���{����=Zxz�:TF���P���Xx�]��}
�xB��>v��s�y��� =���\	�L�fuC�����S�϶yk}O��}^���i*9�����+�%��B���W�LK�:���9���WK�
����7<_#�Ze��c��/�Z
�h2)��q>(g�޽9]L�9z�	�*��穵�yi���o��Ъf��㼬ojءtسb�n,w��jۿ5���+�=ɑ�2���&K	!���u�j��l��s��7&��5��_�@#Ǡ^K�]k��=���BJ���P�zD+uC�ۥJ�ur�zmN���|1��؃^݇t7��2�*Ե�w������#��J���~�S���Ay�8�m�sK�y��J�b�'b�-�c{�Dǌ;�\.��a�q:�{��f�9A*5n&`���Hd�ӧ��V\)`�Q�+�od#s�{y���{ծI.c��i/Q�PT68+"��x��RP߭B�eQ`�H�vI��.79�E�b�H�T|#4�@|4`��*p��^ZdLC��U��'q��G�:lOP�*�T$����=U��*��Ѡ�yC���B�5����/�M����2���..&cR�����^�,z��0ЛP��u��
ͻ�V;�PvЫ��~�PﶸŁߌj2+#��aW:�cEq�	o��:y����r}T*��XӅ�/�K��=0���z%�ݽ"c�rfR��7�A�5�I�Ͼ�P�r�����"ψ��*�Q:{���8_{�фn�űX��+lY�R�`ډh���ǉ���ؾ7�����>+இkj�KW�1 �]Ax	v(pV��L�K|=�"et{ޏ����Z �VX�p\��CYTϝh��P��(��A��~~�����W*���J-D9��v�ӷH0��«1)�;�G����KVh�/��m����N^�{ى�n�4��������:Zs�΀�Pw��1/�����b�(Y�}VGU� �!���<c�ur���$Cg��Hm�Bf�g5f��}Z�6�X�v��y<�#����i%�-J� N�BZ�(W��÷=l�CRM��5K�qν��h3�ڊ�J��.��2긢*�(��CBf��ڮ�z�Ӟ�g�ر/Ↄ_N�WD�S��Tʡ�9QT��廐r�u�%l�ޤ�p���Q���<�$Wi�EX�,���C�E�\ˇ0�{9s��P6�:6x�K��Q�D�B��֊�ֈ��S۾�nGɻƫJ�g!x]�/��lbȦ0�޹��}5pH�g��^i���C�F���`d��EJ���8GC�2+�8R<3����H�~�%�a�=�����k(i�o����[���&�x�)=usN�z;����E؍n�e���%��<�l�2Tw1J�{�TW��]�u ���֟4��(�CP"	�x7}^��D�ۛ��xU��?�Vo�l/�{]�%]�����`�]ǜ�綹�Io� ���6��l/མ=��k9��c��"#S��]��:��;�M���љ%���PFP�]���|�t��F�U2�(>(4oMn����w��9ܴ��\�9����P�Ɔ���ᮙ��0%�4�ho>R�1{�o���I��ʄ����6VE�nX�L�:zŽ�^j�*��3�v�uGWsS��t,��p5�^$��C/崾2����[���n�Eb�u&Jo�Rc�w$�v��PN�Q�O�.4�-a���Zx���7J�]-<T~��V���[/<޴_h��M۫(=���C�^,�¥q�+⨱���۬Vȶ����_Q<���ʸ���S!u�aP~�ZY\�^�}�fй5���9$��
�hwN��J�P�FЂ� k�q-u7O�v�ev����tU��%h(.["�h3X�*�K!��>N���Lҹ`P�ڤe��6g���r\AL=�G��6^�J�k�.񴂛3F9�M;����h޼'�+O��^\��ˁ)�v�8��#��kbs*R��Ը�ۖ��YO�+d��}խ�27�?W�W�o��sM?�]CiY�\h[�E̻�7j�\[<1.м[���6�z�4g�=�ʫ"�Ғ�εT	�pw*����Ϧ�C/$kT,���_'Rz�xt<#3�e6@c�MPg�	��.�U�'�d�^���������Ժ>P��
����MI�]�{�˧����ǎ�&%��e3��C��x�������|>x��<Y���u�`�!
��-,���˰݁�:�#��r�Ly zkS�-Տ}CSo]�5�j�"��+�27%q�Pܒ����SU	F���)�eB��J1δ���TF��l_�	r���:}5VI˾*��������<��A�|�i�T�8�(��[�z祬�K��Z��},`�����=�UY�P|���%��7�����wQ�&wc��Zۯ5�괶�#ӲP�ӻ����*�5���X��2z�-�Ӹ
�/������ڽ��#�y�"۝*&����d�b�::�3��q���V�\eoe1���n;V�s%IML�d�KJ�5_0����qn\O�wqu��	�@�Ü��i���v�뫰l�������T=]B�S�d7���U�cZ�W7ԥ<�K8�!��~�mٹ�><�.@�%z�*����DV�wiB�f"%m�9��>(JMJ��ζF&p��P��AX:u�j�zu7�dtvv{}:������)1�d�j�����8JR N@���S���6��싏q��P�L����*଀��V�m�����)�X}S��Wou���!pA��V�j���!�P���b�^/�ة\y���9q�t魿p��r���!P��B�T�V}"��h��P�/��h�9�w}����:D)���(_}+�Xu-\B�.O\�2�D½b�=��/��6'+c2��shW�T��"����'�a��nJ�-����u[U-���3����M��ŦxU
�౦�0Eb�U�=_Wo�/M�(�7�a.�Cִ�V���)6�Y;K���R�f/��H�&r�kZ��%綥ߍ�lVpQ睽��tg:�j���nKK�&9gqr@S�W̽��^�z�u�SYd�0�T!$o�����eh�0z����F�t����q�����/Uś�L�M-��i�����[�ǯ�V.4��"�R�j�TºυW�>�;4����y_�6l�D�)}ł����m���*�~�����G2�vnN���|ʉ8�3x�"��֚�҄ޡZ�f�j�<YX��{�}�]�u�O�"BNiV�o��}��
B]ex��'���Q͓.�\�-*&I����@��8�����+��jZ�3��z=�����^!ix��S�QPUB�Ze�Z�A 3�(pޡ�٨��z�8{#�o���u��*�ߘP�kG�fQ�s(kV�L���mz�ի��ꀲ�#;�:*�����ؐ[�1U]3g�k�x�M�m���ްw��1�}W$�nt�Y�L�t��u�gAwk�S�)o���#��S��io4ֻJ<�ͮ(����5�� �pO
�vS�3��~�Z�L��-�?1m1�GNRon)�ҹ��B��2)!,��K�P��Tt0�����Ю�dW���u,�V��\\LӔ2�]�,mWx�(E����ဋ.m�#�7Ӈ7uT��Uޭ$��m2*��A�8��XدZ���eeܻ�9�2l�n_������S�cm+?	����Ԍ��H̻��^���5�_:�GG�MU�g��#��ݴ�	~Z��t�i�1k��Ŝ��!Z�=�p�w2�o�����Ǫ�ҥ�P�6���x��_�y�w�p:`�M.86S>�:�3�ݸ��%�\�ҵ9r���8�!Ѐ�?j�V5:Ը���l����/�ŵW�NT�7ͺ��ۅv����%�I��.+�[C�m�ᮇ�>�dWU��ܭ�`߫d�$,�`ͯb�S(�������u���mu3�ҳ=�u�2�=���<כ���j�VS�߸��Ev��,��1Y������j���݋��|�:zN�p��,��k[����!:ߎ`\�yܶ�]��㐤�,u;A���eJ(����.����*��TP�B%�'����*��ig>�\s
���w�/��v�6\L��,.ꡚ����d n����X|�^��N�9�YJ���g�}s��f�.6<4a�T*�QL�u�Y'�)�LU���~��wnܙ����ʦ�]�
��Ȅ3؍-k
���'L��"&��j�U^׻��g1Dt�0Au��VsWN�&]Ãʋ�b��R0��p��gk��L�K0�j	�(���b��)di�<8en'�e��a-#��7�S[�F�]�|��ء���VVQ��Hy�V<3�"��w���=��*S����$�X_5C�L��IZg��f���P���4K�����R�R��O���u�wZWo�PŁߍbke��=~#�Lu�z��N]18X��m�������(�x���:w�K��C2S2ï�bz����j��E��xz�S����l�)�,�F��˛�n�(�Seuh$m�]�$�k6�_e��&� 2��>ډqt2��r��-��$�Vc�]T��P���KL������F�����;�O��[؍eI�B��<�ž�촭�
lQ1��kRZ#��@�#;k�Ե����ѧ�%�����ȁ����6r��f;��/bNm�]��+�����m����J���7Gʐ��';4+7�V�����I(@Vr5x�{����٭�椺�ۦ����6�|)I�(�l=Sp��w�)e��ػp��Rλ����{�1�]�@Di���W��}w7�G��.�WXd�7]��}�eo@��M"��m���cj���kW�mj�,���2�d�
�;d��t��.%�z^��!;�% �|{�X�ޢ�T�մ�jx��g2��4%,^>>�v뛶�*�F$�S�B������Br�|�OX����g	���/�Qh��)x���.�~^��xx�vo=���G{���.��J���oH�D�`��ڮ�ބ�s���rU��# �T��6�p�Q�4������	
@UޡKxXN�2�Tպ���vb'9}Z�+��Ǭ@*��Qs"��ڼU�P���t0�t���
�P6&X9N+'� �I*���n��˘fXrY�4�ub���*�� �oc�?!��Z�Sv$5}�S��YJvt� �S����
��R�������z�O0��ʒ�&��fYv��Õ"Kr4�HU�h�v�C-��� E�v���圶�fe�B����*���b�K�C+_٘*WYV/��m���f�e+�o(-�#0�R�<�d�:��G�1:@��[���.%��m����U+{�W6����,;��ۧ�1�a�d��75V�ɓ�pHz�^:�F�N�S�4Y����۵��4.���Ѣ���qԑ#���m�0��DĆ��	�p&�"#+g����-��[[2�����}VqwWi�C��\�٦��W.[�΢�W"p���)�©᫦R��YwMW��spm��n�]�gkjL�rq ��i�:�m�j���zӍ̮�Jш-2jZ�y��_t���̾]b
������YE��bG'���\�d6�3�Q����� ���1�PZ["ʲ�U�[V7(e�"�UQ��(�V �b��U�T�*![R�kPPY��Qm��Z�*TR�m�QR�����%AIKb�Q�+X*�Ū����%E"%J�)U�R�"4e-�mѵ�jV[-*TP�J��TUFT�F�T��%F+*X�Q�m
��U�
4B�l�R[aX���ETJ�b��(�"�Z�b��)m�V�-Q�@�Uڂ��-T�+���V����1Z��V�ҪԶ��,�)F�Z�lF�Z��DBҕ+j�ԩEKK*UF�m��J�E�
���YV�Z��EJ��cVԅ-�Ѩ�ER�)F֡@h�-$�V�t�G���K"^��ÊI�.���PB�k4s�)-X��s=�k�a�9X����[2wm��U��8�4&�P<��b< M^D�t]�^v��N����0ӕl,�p/��X��ϘLz���t��q�7)�܋��}f+�=�ƥ�:P#C����/�HV��W���tl��Y :J��I��bKv^o���ţ���O����>Tt֙�j���f�+<_�ff���*�yl^u_Yv��l�C�3����t
�4��ċP���}C�z��2ۻ��l�I��yp��V�lz�EG�R��Y�Y�upP�2e�a��u3p
v͟k�N��Q�J"�]�C��w�=fj={��v�����cH�	�ŵ�;�S#pz��/�C��Y�T��㐣OY�Sy�MW���^a�)�ia:ڠ:&�φ�RP$S���x����?c��2,P�ZZ�J
fS
ଇ!g(z��__�T��ݷw�J��gg�l�'�)���������T��i�T>奺J�5��c�`���Ξ�b������٭�O�_��o]�A�fVS�N��p��}\���GG&��WA1h-�$.�)Rɚ�@NJ�l�Xƕ���o7w��ʳo���x��J��c���L�-s���kڡ�s����z�ڣOU�}�S3%x����C6#��+�v=H���ϻ��礳�|r�ڽ�-(�G��ŏ�L�>2+?,���^o''7{Ն�u��H_^֗�^7`�,q�X!Zp���[���1�������B�TCz������gN�j�8}�Vo䴳H+��G_ަʝ�v�<����^�~h{.�ed��>yS\@��yg�{��������~�T�~Z�c�[����|g��b��mp�퍮k��\�<G����0y]J�_����3R��\�zb�?��+�Z����	n����SH�R�/3$H{�}`�|ʉf��w
j⇾̭7�c���;q��T�ׯ�k���*>�� (h��5���ZL��/�f��]sgu��(�G�A�80V�-wW1Jl�����J]�fa� o=��wB�zi*R�Vӭ�%��Qškr�hW{�o;:��F�TڙHL�ȴ��#o�œW�yޭ�odC52�s�:Ԗ�d�V�o^Vr�p���Dk�ሺ����-��ϔ�N{<�����$��o��⡗.l
��ai��WBii���y���z,�f��.!�ڃE8�%t��,�:�x���[�fV[�q�0��<n֖|
9ș_v��$��4諎�����dŹ��2oL���ޯ)dW"�v��p���]}��2(��40�o�
����~���i/&"���Y�g��c��.(5.���0->���~��rySU�Qf����~	�{Zm/EcS>7�ŉ�0w�8BK���+*�[^���+��(],7�:�,���C��C����h������pu�x�ݗwv�������k_��͕�ۋ�ь蔭0v{u�U�s�x�z���3�1-�,�uſ/�c��y�]dT��ϋ���}�ɨ���ݓ�Jq���t�F�
��ra	�j�4��ͭ�Jj�T�*ˣ�׮`�����\�s];���8Z�ֱ������H牜k���{ʸ�fw���9^�kz�ߘ����,Z*��I���l�%����V��i�b`�ⶄM�w]w�|����E���T���u�\v,��P��2:mql][�L����Gs�ќ�����,2��|�i&�\՞�����B�f��Uon�-Onx�yȦG� �CK2�B�E�?�'ZZ�L�7��dm(s;u��Unܑ�ߟ��^>j	(gU3�n��`N����$��ʋ���u��x�����y�a�t��>4U\i�����!|�@7[�9�0%�o'���YZו�j�v���5��P�@�ƦY&멕뼮�ùJ�p��y��I�aЃ����U����W�dz �F�L��04<a��[�9���ON��#�t�)z�H�X�b�_.���K(u>Tb����Ω^�y��ؙ	a�C\�E��^m`���^<3b}E+�z�XW�8�������c�1�萾2����IE��pn��>�Q Ħ[�&Q�\�M)VTڜ�-*�#����]cU7N��]��Γ����j�uns�:���4��.����[̽�&W��V+ҚT{�>��q��8J!�lx^r�r6��+O����]:�t�A���6"�/�X���Y%i���3P��hb���!W`���zn�x������Zjfިb�~"�z��y8z�!��~�\{^��N�2��7.�QGz��N�TK�C.S2�a�7������+��ǡO��=��ț9�V��K��=���_�����'Y��U��o��]�1tV�!�]3���f|�Iz���"�=��&b�H�b��+e�L#(��i���N�ę�qݳ�agu}���{��}�ˮŧ�>�V���փ��mQ43���h'������[I�}aP�U��~L�mq��"%G
tΥ�yq뾽9AB���6ؽ��K�w�>��^O��V�+��Cc���/���^
�),��S$h�u���,W�'�}u�wYxKuyL�v�=T͞���q>��
�a�����|�Vm<�m�/�j�!��)2���U���!��3.<Q9JRf2�oSk�Υ�Vs�ֻe^e���]��NSX>�T�k�0"�)�>%>��C��J�S,��2�{gSm��tUg/�p6��xALX��XO�T�+��t���iA�_w\�u�� R�ս���&�A�z���4�0��P�f��bY�D�j�^u���)Z��6�*?Q4��1B�p�m�EId�#@�c��\_fV𗚚�EǙ�=&���a�*���,c�]�!P�B��J{�w��13��r�ZK:���VlAH	�U��hz��9�T/��0)K"a����������~�&��_��NO�O�(x�m3�R�W��]S_�"`�W�ߌ��C��S��R{�i�"z݅=烴�WO�I[/ޥZk�S��eс�����42��%��o/�.g��Е�ٞ:p0�hfՒt� [o��t�$j�7K��ԛ1�"�{;�X9VΜ4f��©}�\T��(m_�qg>�4j��n@�w4]��w����A'�������%���+^v'�f��k(���gx�p��έ~;ā���S�����ݵ���7-�ZާY�s�n"믍#Ϧwg��D&�6\܉oL��{���N�I�>���{k��+la�v�}�#�z���:G �eV9O�3�\帴]P9�����
w���)�:8i�lf�܆�����S�>
B�ƻ�>`�sJ&E�w�*VE�i��	�)�}P����a�\��ֹ����fR��[�5����P��ƾ�Ɍ�Z�WN�����V락&����%ޜ���ʰ�%����#�3���(XT��>�j�S��.p��{�*�{6�(}�R*}p�b���Ze�qD&���x/q	J���ːG����U�(�}�C�VSJ꩛����v=9���/�v�U���Y���"_��L�6�����9gٝ[�9�h�*���>�B�g��L��G��_��F�����u滙��o7�j֊�=���GVEnP���"���x�(0!��;9c2�u��uA
�Y�3�[1�L�u�Xq1�*/�+]u�Ac1���hv��b��Pp�	-���]z�%�V(���#X�x��܋wG.9��0��-���_J��E�RZ�JMA8p��w�^��o�����u��c��.}N�{u87��'/r9��p�(SP���E�=�
��0�~����G�V�7�g��Kڙ5˧Ƀ<�7�B�4%}�ҮQ�~]z��͖�����gC�N�<n:�w�����4˿T1+�b�:Wc���^L�<�鮳��cW���x�Mc<`!
/V�����$�l�lzT8q�5ޭ<ps�-��
Cu�o������e@�����@� 8~k��u�=�N��.���:b�����2��S��><zj�+�B�p4�i$�tu��:ۦ�yV[{#�$�:�Tw7���y^"Bn�z*�����N���dY��ʈ�ͬ�#�7-3�#����W΅fݳ.U�7��>�X1%�=ʲ�����q�3�v�4,,:GyR�.��	�l*��@讪
��:���
U�n�J�ڙ*��q�i)H�w��^ڧ��W����,�c�C8h<���ne�z���"��7�����A��`︬w��7�4A}A�<)�R�����zcv��F�=�-H��:�/կ���Ｘ�G6<4r$U|�/���cS,���nJ\��[{����+��F�C������"�)_:EP0x����2��\i_��"�~�a���H
XtOޞ��P�\�M9{ga�}�I��(n�rԨ	ơ�Ԋ>�
�u��tJz�T��J���	�{��=��8p� ����b�9m+ �(}g�fQ�􇮩+wyF`����k^�y�3�
Sצ�hE�_:�`>��P�˺�hz��P�A?k��Ku)���P��C�)XG�9,�����Xl.��#����/��1�+�P�w
Th�G�\��z�^ިa�#�!�t��Ye�L��F������t6��x��agԸ��+���P��:�+���ve:{�6�X��t�dO��0���f��<z��i�.3{2�؎����fh9@�B��͋�%´���w�4b�R��k�CX�Vl��� >-��Վ�$b��������}b�����4���56'x���қ���� s���iNzv&9nӛ2��gfy�mo�佨>X<�y&���Ap4�3*��t��t��n9����z�Zg�9�Ƴ�����3���p���@��D5�uy%9_�g�H���*�:����ύӦwƼ)�έ7A_����s����{��'�H.�rG�7ҡ�^0����`��iD%8m]K�M����^���
��գggp�C˅?�Z����P�z����}6&ٲR�F�Z�x��xO�1��%���@��L�[�}������'�I0�uq�4P��P�jV)�Q��1P����9C���7t���Zg���o��	�Zw>�\$��(D�V��T��!H�~5.>���U��<��K���f���=�61ae�mit%FP�����:EYUO]ie��^��sͥTgڣ>�_�7�C��C(]��Ҽ�y��*��0à<kA����̾G��!�X�szο�ɱp�i.�dnj�8�8�&���tMlj�k�e���I�:��{c)#�e�Q�gQ�\Vo�Ֆl��y����r�v���ts8����%b���V)�5����O6e\Ô+�c�!M��"���АY�v�I�,��H�j��h���3��ʤ*��D��i�]n8�z����k�x��/@|�B"�5۽��D"�]e��i-ޡ��`�}:hCff���c�닱V�m���y�
��8��l M��L��-�jH4X��>y�t�vM����I�صz7'������O�����ά�WN�GxlA��Y��W$z�����e�X^u-Fl�x�&�h�2u�H"u���Űb���ۛ5�n����&�cf*L�O�y�Y3^���D�}3�~�FK��q�=���ja�F�n��8�ux�as�] �[s���w�VۼZ_
*�+�g&�s�������}�&f�TYZz7W{�ZE�q��"��wA.%�	�l��z��F��{C��n����XDN��Cqi����;��B�,_s���v�Q}t;\�~̧��+�aGn���.�n>./7q{��Jݺ�tT̙��(�V�/�U�+l*��\����h��h̀wj'(���y�f�GJ�KI$n]J)� %�S��.�4�a��[�p���i3i��>�-l�ҽ�WF��6U�x��W��D�(5B	��ۣ�x�,M�t�0j���%+���8�u���C-ҹK�e
yX��,�I�M�����&���2R4�镒��MN5#��D�E�d�G�J�|c-���y���ļ�l�"�s��ꢲv���;��\WY�u�u�n��D
�U��ѻ�L.���Տm:7�B{�3Xp��iU^(D�6��)��bY��s��m[�Ci٣��mՊh�fܳ�Vے����\��h&G~-,�Q:����n�pх��u�,���4�T���!�z����hl�7z���b��R��[d'��h#5�����2'��7��X�R�)�V:��B�.����S#�M!��q[�VIqٻ����܍���˨ͽ}ڮ���-�]�^<M�&k-�=���ocቌ��;�)�6
d���zӭe�]�ޛ�x�,�k+�E���++��kPDX���em�T�E���D���F��Zҍ���%aZ�b��ԵV
���*�*��J6ث"�����l�V�ص�@P*5�V�kPm(��X���(��֡P[l)i
��B����(+m-"��Z�e�Z�U
�
��UjҌe�J��D��V��eJ ���Z�ajQdF"�Eh�E��"��*�Ph0�
���V�%h�Z��(�EX�ZP�U!Q`�Z��*�l��*UX��`�+m�R�V�ص[lA��b-�~�^k�>~<��������\�Ƌ�;�]-sB��A�2r<0�*ð�m8�u^���jB$MM�&zp��&��Yw�ʅo�
[j��B�Q`�)�~��;�C��[�B{_F�b/��+"�Ϳ�:��D�{Z^
���7��(bp�|�<}3"��:i��PID��g���vy��:Mu�>�,`�F�d��r
�|3�tb����׺Wҝh#ǫ�Ɍ��\�@A�����g����O�k'\���+q��Z`�M'�Yg|����B�w�KIᢲ�&��~m�����b[���ى2�fA��o�=�jݭ�j��~��n��V=��L}ɽ*?�3���U���j��dP�֚��7��\y�=#_{7��></���Y[��0�����*���8��r٣~N�#l�5�l�o��zy����:�n�^{l�L������-R��U���͎��v���:��d�����"����p�ai�U��u��S�B���W���y��=��+X�>ov׭�/����rU�77�*2̂���^=�EN�� �h*z�T�Ǐ!���P�K3��39B�K3���3�f���V��ѓ4��%͌���ZH��0�T]a��xٶ�E����A��Q$�T<�[<or��=LV�g�
���f|
9ȗC��v
d�]Ɲ���̾v����=�g<�8$F���Y��Z�+����g�,.��F��G
���>g�\`D�+�=U0���gy�VEnP����X������y���5�<T�v��u�,ٜ���	����^2���,M���V���>�}R�p�p�f}/�j�Ua���=�
�"_�C�����f�M��c��~�Z	��O�4�dH;��!�*�/i`��+���#�������r�j���{L������،Wj�J�[\_y�C�4{S�$Y'��efn�r��AB��!�y��+NWSI�a����ߙ�n��]uܮ/L~�������43�n��@�8C*�����.9���*_8�!��s/�ʺv>��\u��G��TYIz�@��]?v��l�^o4�'��9�YV�D�Hŋ���8��7�X�ģ#8Q;�=��BM���p]�m���5��\��t��$�l�E�2_]{L�}����l;],Cl&)ZI���]K��){���;�ٰ��yG<]gj�-�\"��8�:�]
�����	֖��"˯?z�>�jW��;y̦���\n��Jk�g]�MQC�7�%��@�.�^˺��wVޘ�Y�,�m�dq���Z|hVQ.�\f�ae�2)�y��쓴^R�y�y���=�<|�D��J*�V&Y8��ࡣ��T:�e���>;セ/|�<oŒemB�
��^�~��U�U�t͸@g��iP�H��!Zy~{6"�|`��V�B('�F�u�ҳ�1h)��Oѿ�Ӱ����]�;����B�b�	,ĩ�j�Z(�XD,�q�u����4m�>�����Q�b��r��y:OW%�^����VU�﮻��Vd���|{\Nfŗ-���ަ`���;s���X$�3�ByG)T³'� �\8�Y�ʯ�fK�4�^�����I`x(^�Z#r�Xz�e@���O2�[E�z�= ���զ�A�M�|�e�љ�P��WЅ][;&k5�/�hI�\�3wz����{�
���è��}���o\1xV�)������D�O�:�t�7�uL}���N�.�WY�p���\���z�W�Pș��lk��_����ׯ�Ί��O��2�wYZ%_�Sה���]�ӯva�&��x�;o���K����I�����Z`Ϫ��ʢ8��Y���)ͷ�-����Ve��A��g_w�I���I֙���ܻ���t����r���u�4vg�>BJ��){Ӆ��x:�H7�]e���i����eZ<L��C����+��1a�\2����ʾ�9Az��C���w'��" ���B�o�R��C�(lᇀ{KS:f��rr<�{\���׭��Qޫ���}ʐ�|�DY�ђP��NU��גBo,�Wn���Vb��l�.	�����3�P�,sK	�4Qh����3�ՙf���޹n���h�^>�,��57�Q�+]f�d��/N2�����Eþ��|%�g��9k���^Ru7��o$��%)��x&��$MC�N��3nM[8��Zf��Jƹ���tg؍*�l15+�E<�!g*�[�ɓ�=�z�z�aG��զ`�I��#<�
�¬>�%rF�~*��U���_��|�e��T�kC���ؘu\@��Hx>����T�ug���4}w�~7��#�*b#�졔���n�����U�P�s�&G��fS�p	,z������9Km^�uL`�L��=�hM��^��5Ӭ5gDܠ�]�������]%a�z��b`�9�WK=��GMa���j	|`{�x'���]yN��	[F�~V{��:l���Y��H�]
��5��U�ӄӚ^r�T�*�J��Xm��J�I���~w��^,��4.SK�<r�<R|���m3ê�,��c��쮾͆7�~"If/���S.��zb�_29`��Xޫh��g�7���j �Γ�ݗ�y��-�ᶳsR��{Q�g�́ YN���Z˱�9*G�5�[�ӛ�̾;(�.TT����[{���K�&M]Z[Ge
���Lò�6�Pۊ�f�W�drn�n�Xv9���>Ut�U���j�,�P�^5��	��P��5n3S=�l���6-��8·%�a}D
#E�,��chu2zpΦ%�.�뻞�Q�=���딮��d=���_;�B��E�Y�|��A!���M�*��3&��5��8�C�&��SK���p�b��g Z`S�J�����%��(�]H�,�p�b%�׊������WD���43��\���adR%V7ƌ�o��Ǉ�I��=C���t��My�Ǜ��Y�EM@��X��Z���)e�&k��Kg�!���ʰD۬;w�DAz��^�U\�EP�؈�-/�VE`',{>��rL{�ǽ��sH�Y�`����XlIP�XYßN�p��L��>�/ci�����Z���>c�l������԰�Y��
�"X�k6�����,ӛ玄K/n��2v�,��rGθ]h2�X��L(�Z�Av����C�֣�,��hKɘ�s���������W4�%)VP�د
����zV�JK�h�w���Rl�����8�px���f\m�`�Iå�����fe}��/i`��i>��3�t_�+��5G�qȡ~PĽ�Y�Zz?\M��y~�:\����b8�U��(+�`�/5�-:3�$�
�p�Pٶ��@�s���p=�>0g[8�$��
���`���T7+�R�+�/<��<k#�����
���*=�8�C3�ʸ�v!`�>R��iqg��{|{=���zOG2�fp���ά�v=ަE�͇ո��ʸQ���>N�hz�O�뮛w�ފC�x!��t����ʔ��GɃV'X�\�T;�	J�^����g�7��+ZY\��l/�!�ƅ,.��:��2''>9+NLuޝ1�ˤ�6��^�����	�vx;���>*��p^�ǲH�ewH��p�d��I��n�j�>K����p���4�
j��vh���Yz-景����L�"�c	�F�#5����,�}��8��JFuL�˲uy/�	m����N0^��ja�r^*3�Q�ƠO��n����?��He��(u����+9��4�Y�+��V9`[{6�Ǥ�ێ�#�ܦ�"ڙ
E~A���ʆ���~�a�Zm+9{\U�dL�̬no=R�n{(J*���xĩ�ju"��XD,�q�u�����$��'���95C\f��p/!���b��i[O��������:t�]-}1�Q�{zPᒫ�3�eЭ�B����2�P��Ϝ�3�^��n���wG�z�O
�_3@����|]h/T0�T1I~#�%�K���:4��b<램+�Vm�(��$��)����֡��r�Z�t�����7>ZG�L��T4�p�m[)q��
9���xos7�1�B�����!Q�w�r[�WJ��O��S��W�<�z9�l�J(��a�V�}��?oc v⡉X}��P\�R�D�=�%g3z����7�B;)����Ũ�Mt�!�����)}�ʠ���N�g7s`��m$Ѹ4���}��9b[v���Y�SW:�%��՘�QEQ_na
�R߽Wi�Ǵ��a�)\iA������w�����~�����R�J��:���tm�a����iK�3S�F�N�ϻs���B��_��V��T9�ʇ�;��]:� F��=���q`�DU9|h`��\�D;tt�T�Y��kz��먉m:w�=@���=��~��%)�4��7�֙��tW�L�"ϋ�U�J@���{�$����7�g�WF�G@�����CJ�Q�����d1W=;��9�2�����z:_u�,�D��HS`�`��Q�D�pD$!�Sk����[� ��gG�T�cD	���bb8uq��TB�2�dWer޼��:vG��wUR)w����)���-ۃ(Aüt���"�m�؛X�d����\t3Șd��8)m��B����wd�,n�Ț �M{��=z<t߼%�����{ W�x=6������^�*��}�_.��-}[� ���'ᇱv��3�͚D��]�bܺ��#}�h��mH�H����EM��S�x@gv �Ե�K���h�LN}O)u\۴*�@e�Z;�m���x�q��wl�c�sr9W^!C�M`�,��3�.4<��%UY����Vx��1y�y�o�^e{�9x�<sBfc�G_�2�D�_x�Ɍ�������em
�x�'R}-8�P7�o�Ք��L�M'�C7�O:F����Ά[z\�U�_]���^l���B���(
��yP�9�L��g��Xwɚ���k�삱y���ƅz�2��Y�!9}���Q;�ٷ|r�dP�֟Vo�ȫ=�=<����8�f���ŘUc�0F>�����Y��z>���|����a_-_*��^ĸ-�­z�G�Q�U.TF�����}�n>�����{+Z��5+�T���Gj*�Q�������ݍ7���jUqDP�H�:q��C��&��_S�45�h��5�)��5��tb��}(r
6\�ZvA�蠴���P@�=e%��oE֓��[W��-�WL*���
�#�ס��L&��,�������_>���O+{k�opl�����٬��u:�
.�_R�V��ᙎܟn�w3�V`\}l�&Z�i2VN�|�R�eV5׻����9D��E��]A��]���@ތ���g@����2���e��bu5ܮ�+���6aպK��SGS�[��x1��`Jty}.	�Dą����겤�4պ�R�o�-S�+K�ʒ�����>�"�4x,�oX�f�;v"�!��Α������ׁ��e�h��wvw�<����;[Č���D�L���dz���^Br
��N�>+�\�Z-�i���E�I�W�Ρ����rD��\6�G�-4�A�*�'����T��R�ZT���;b�D�]a�ڼ�g�oBM�Yn� ��t�����f�.�K�q�����Q��49�\�i�w~��y5n>!�+����rU�e�r�Z��e�����Ý�L{�:�w:�gd��#ot`���R��J���[��K�k&�Ӛ�j�V�FXڨDgI�����%�m��r��k
Ѫ���T���S���.�rRe�dR��p����e�/Ye882��B�[-Ca%��|�����4C9B���X��m�a�&Q�������]�������i&���h4l�
�e�{I��F�۠%|��Э�řp+��l�I�k*+��/*B�D�+I��+�����²�����of񐏺R�,�R=E�X��8Y�6���⽳[F�҇X얱�6�JT,��������FJ�f�8HE0���F.\2�r=�dW5wlv�ҧذ��]�L���Ob�������8zm����qi�7r����{{SL��t���z�l���v�j�9�魨h;�����W0x.=�F�Ɲ�-�1��
b���4�-eJ}Ytx�J[{���;�#��<ga�gGXP��<�6q��ay��!���ŦvԖZmkb�T�o�wK2�ǜ�E���>λ̊�/�="M�:���m���8��t���+8�N�+D��WJ��ز���Q���[T�F�����ڊ)�Z�V��V#��J��Z�)jl���֤����[KR#��Uh��h�b�E�������ʈ ������-��*�+KlJȢ��Q������)V(�m�HVV��X,U���ڂ�Q�YQJ�lb��d�ְ�`T��U���6��F����ªj�F*��V�R�������EQ��P�-�DEP��EV��СVʵ�F���+�QE��iaBЭk
ʨ���m�F�+Kh�U�V�h�m-�Ҩ�iQT`��QE�Z ~	�K�A$�L�3�q�V���{;��tJ���2��#}�:�n�&nB��80V�FȂ��r�N/���ޱ2��.ٱQ�Ò�`�/���^�Ȳ�п�9��۞�e5�j&pЎ�+�3C\�EG�Dv/Ԕ�u�Un�~��x�W8��>}�g�y1�a|�*8�lE��3�6w�xn A�<-&qܘ�[�Ç�:mA�P��(b�����ů�a_҆,xT#��'Er��ݭGX�^.U3f��W����	6���Ϛ��g��qX~�K��HNg�{5�<��C��)KP�*>���62T//n�B˷Z_���\��D��W���f��|A���Ơ��O�^j�1ZlgTI�*ҡ�O�����J�ݯ,�P�:�z늰���QЁh0p%�m��Ը���?{%����ǜ�^�)��&(GOW|���/���t!`�8�2M�ŻG���;�N�4}�5�#U���}K�G�m��3��b�}B����q�ul;��Lr:kȐ�c��7�骱ާ;���皕���Ɠ3!�'Z���d�Y0E��K�_Bۗ�!R�_��6��q�>\&h�T|�#'�����:b���dD8A+$$�4=$�,�S*��8x��U/vl���y#Sl�	��[�%�?^z�oh�1 �-��*�K�|�5�U�n�dD=$w劣��x�\��#�hq�K�Uƾj�^��9�L�Ys{���� `�P4$bpZ�5�Dߕ'k�捞<,�e���v^�v��O�~2�$Ю��]1V,4o�[���*)��N�k��/p�'�������d�U!��Z�;�3J��!����u��@�����s5��QÒ/=�zf�,pC��R4Y�sf��]b߇]z��W-��@��[m�v�h�eڨ��C%|�*��iY�P���c-tܽ����3�K���a�]
�e��I�6�f5B��*�>���^}���ۥ���!�	�1|�ؑ�XQ�tOT0��Pł_�;[�%U��f���}��fM�%�a�,#�ͻ�Cg�[N�/I��{���S;�����댲��uAN��{��Ea�8W}�Q;��	�9������8�0���s�S%M��Z�S���8�<�i�3	���sg�]+6�|�l�{���5�V�G����L�G{d�߻;�yn��mjX�95�"�S<f���Ժ�PAt�0Y��eW��oޛ"������wC����Z������|��Q3���j�Dc�~p�W�6�x�2y�4t����i�U�l����i#�/
L�2x�.��e(��զ%��8�;�XC�Ug���L����K#-��oC�t\^7�`�A��#9(Wm�Iu3qB�x�c�꼛�x��ʠ��9ޞk�7>ZQf�Z�W�����HW>��Ҥl�tΌ�����KN6�yN��=r���~?o*������g)��Z��(S9��F�^�y^�	�1��/i��yT�k�bT�5+�S0�B��S;�ݽ�����*,���B�B��/=D�
�D��(P��O���wmY]G��&H��v�D��f^\��j�|���%��.�g}����bCl�]����9O�И�����khZ�Ncj#6�w�*��xGJ�s�GV�*iU���ˇ�v��ט��b�������w=��a�T6"�.�^ ͜��3�ug>,4KԈDX�p�����c��׵�	�eU�I'<��9�R���e
�1�.��e������/3Q<|~��~�ǯh�_���KmlC�]SW��H73=36��])�,=w�/VN�fĕ�\����a�D�ť�XoSW��n�h����u+o����v�#�r�������^u�Xg�������װ�3������׾�^<mF/������&u`>:{3�r��X��^�k9�R�]_R��LmJKG��\��zb�8:�]��TD1nym���W��{Yw�U�X��������<�	I����R����@���3w7�2Cu�K�xKzFW�N�T*8D����/���RAO���w�N~g�_�zg�\5�P�Q՝,«�a`�0��i	o�fX��יC��$~��y�3� v4t>f���Ԕr�g+vM�*]��7嫉{�Z���4/��n&�*�Ck%�B�h|��V��޹q��F�;3��X��d�� \�-Òeu��},�`Cb���Bz�<j�����,��|�h/
+U���|:��{��s�
y\�hj^�P�P�"���z���s�~���Xv�aC/�(��H�8x���1�Lv�������n<�y��fgN���4S�JAU��THx�.v�>�o�F�"X�ͨ_�)��7�b~@�,�+h�tG�h�T=�,�臭k��d��o���^4&Q2��Q�%�40��EzOb"�ե�VEa����);n�N~�\�DK���Lj]}�-QqC�,,�>�� wG��X�cw����)�i����^��@w�8lu����Xlv�ؽ�L����C��
�/#����`���V�65i��>6�$il�D�/��2������ܻ~�5��͗V��[�����gD�i��KD���6��ռ�ޮ/�L؝���k�z�r�yW�ِ�ûj�d-ZC���P�,sV�[�mۮ�j�j	��O�k=�|�q��ϊ̭� ��
Q���v7z�R�2۬��J��r���ʹ����7�?�s��Œ\�D���9-9ωk[�ݝOu�7��<���]���C�C����i�2��Ʃ`@#��歅�s�$���=SP]�}�w��5bǆ��X�3�C�Z��F5K(R���}��V�y7{��\����n��o=V��j�Pl�^�C�V�n��9W~v!�AJ�M�r��=�����p*�u퉂�rVt=�i��Ա���#ឱ{G�g��o��m�A�1V`YZbH��C`�n����=��sݗ�e�߭jZ�^yj��B�J=����MieE���h�,�6pu��(���yu��П4W/7g)ׂ�25N���c�Z�5�EQi�~�dKڣCֱ�HHZqMY�v,K�غ4p)j�Z�N�QvkbX|�졚v]{<v�9iH�^����16m�L�j�aDh<s���6nX(Byh�e#�{:��շ{�{���s�l�.��(���1l	�KC�P��:�F"pL�Y�X[�s���W����Ew�r�f�;�r"���CM\�tP�rw�໵�8�zZGLKkWV�n�wq@�̾�.'�N��i1$n1�z�y3q�LYmz�����ڶyx�.m��*n[J���l�^�.�|��x��6>p�Ҳ͍u�yt+��BǖI��c�X{1d�˻uz䘛[վ^/.������f��T1׍���t�{��m謠��O{��)�"Lۇ}�N�6'��^����۸pR�E�=@\��eV]�k�==%��Jui�%3,:�6'�Nޮk��|��V�}D�l�8I��[�o��%��O�҄��Ȗr�&	|a��Ca��X�j�[:pPC���딛˾>�|�^�,q!^v�U������AP�v��� g[��>��ԅuݏ*;AX6%���7�"Ǝ�l>'�~
ƹ����B��~�2�k�����W
�'��N�桫��T||+����v*�yߤ�؟�T�}�]Cl,��������Z���g0ʆ�V������k�F�,�|�lz��_-32*��
�;����T<�W�/�uW�Y(���_fW*0���Nq_Ƿ��'9���� Θ�Yg'��[�z�]�No=�Js�1A�2�8fb�Y/�C.Z�u��l���h"tt����\w+����k�˛'OS��D��7���:E2�I��g	�����3�U
b�o���l����ߟjN]UmClJ�Ǒ�"���8�t�(̕�L�/ݲ��y�X�:�Q���_�5N���L&I�(TN�滿d�o����MRQ�D/��U�px�P�-�p{�p��:%��w8���g2t�{6B��2��%ͪ�kJs�賞P�/�ЫTY���x秇:W{��t_���%;U�σ���q��!o�p�Զ��+���=�ck��o�u�4��n���Z�mC ��[�|nJ�,?z�jux����z���s&��fT��U�����jB��r��q� �ZnJ�bzX�`3�H�[[x��o�O1X`�U�	q�bA\l�H�:io�Bc���\�,r�Y��{ ��\w&������{��-��i���;E�yq����N�
,S��J�2��G0�}1;��{c�(�V5���9$�U���͡�A��{TKp܊��1h�.��VK��X��׭7�� j����Qb}Uś�L�Ji>Yf���=���[����ѿ����
O�w��Y��xK@ A.�P5x����㒩��L�L�vd������X��X������Z�?e
xN1�1�yu�ʳ�'�|�lp��u�u�����4cV[P���������W{ٙ5���;����Z�W�:�K"mW�VhV��d�^T��(�6�h�R�˛�7�AYA��z��������WEW�����JwT���M^F��/5|���䴢JDaヂ�D�Q׊N���]�s�+=7z��.#A�6�EF�Z)��q���Uq�t�*��ś��,߂���%⁬�Ǐ�/N����P����hv�a�*�J�X�B������*�=}N��+3ㆌ(�[L�@IQ+�j��ET~�E��Kʬ�'�UJ�켏��&r�*�ﻥ��~x2bí�>���D�a}�Jr��K{��ن���8J��ǃ��5�{J���\�ݷ��/&lDcz��Y݄�3�� L��������;^�s�Ej�eC}�A��5�����^��Ua��0�PXi|���^ ���� utx�ϛR�^�N�$N^5��"��lX��7�=B����"���5Cˮ����zg1����2l>^�
|(O8s��b��(p�ǆ��2oN^>��J�g�eq�|=��y����S��F��k�n���-�$֮�Pu���K5�ޛ�<.����})6f����||��4R��F��u\2�n��Ɗ����_���k�[/a�����ڦ��A^}�c�^w�5��T
L�^�s�gz�$5fʥ���ZX��&Ǐk��w����O�ʴ���Ǽ��M`�Pn���O�Z������o-�D�i���ƕ�~�����?gz�1�
��=Ys|w�
X���
o�v,GgJ�q:뼖r�y+V�W!���h���ե*Kϖ������e%�ս*pR��c�ՙ­fPnr+�w����P%u:G���]SY���d1�A��l�+kF��#����o�q��9� hv/���F�{W,��j*�l�E�,(I��1���T���n)��]�� �d��SF[�*��������ԬMak9]8g�-f R|;+{� 1rZB�;Y��K��a{j^�f_ӝ^���%mDr;��&T�2T��mr����tuؽd��z�R��WB�fH�21�6e*������s
���K��R-�WSt�]cFF��߳����#��i�՛A!� �6��?H,�9J�)�;^����ص�*��}(U��tr�j��ki������4o�Ҏ��fͱjf l�]a�*�V���r���@�Qob����$�r��եi���%������geK2:�d�Y���8�w(J���b�B���2U����&�[X�ݩ`�����rN�u{'�G��6ɕ�^�I�+��������WjC��n!��U:��Tk,���L;�]O1�C�5���O�sR�����}y-Gᇈ0�⺒CY���n��n�'�#*���إ�Ci���p�ۻ\,�V�����k�d��s\.��jvWr�'˒k���s����5ܨ�rč��ؖ|5�[:�u�l�y�C)�#í�TC8�:�����q�z�/��� +�"[Y���H�"��W
I�J�vU�+K�x��s�(�8�R��|"�Q�+k;�v<l�G��Yܧi���F��g'Ʋ���^o=*�,�!d"�V�nP����W�.x.ΣN��],���5Cv�[/����S��RG��
�;]�;�i
��[�lT83��J�E���׊��迥��Vl��N�c8b�ǍزNk �/5�fs$�YEu�����Y�v���_m��5%5�H�-����ܵ�Ii��'I�s3�z��[���w2�����P�n2�W\�0lFg�$�Kq������%���;�*>!*������dX)l���]�yk�z��:>�X�F�iJ
ղ�J+U�h�A*Z����m���UF"���Zq1"8�.32�Q"�[,Te��Tˌ�q�,�mm3
,��m�m��iJ\�̶()1��m���ZQ�QAk�,�-E)�4ņe�Ve�R��b�(,���
��[1�E��˙G0�-�̆(�¥H���%f"!�2W9f&e�eaU�Z��f`��
�-jE�XUd�*b"��*UKJ	im��`�bֵ�1��KV������R�"�dh�1�ƫmnZ��̈��jDV)r��Z�(֮Y\UY+�࢙ed��kO�<�{h魊�rd]�GR�P��}��S�f<��V-�'�1�^�o���=iCd�I�#�]�u��)ץ�Ӹ��,���痨����I�|9�=ͣb��	�г����{˳^n�Ȭ0�I�v�沺�n�N���Ѡ�F���������z-�F���1=�v�-��*�K���Aqz絝��h�����GCn�e�64:R�g��˦�Җok�7��u�LO{�|~S�N�tw���zT|����-�'����G;=���^�`��H��BzLf_�ץ>��ޫ�>�t�ް���k{%����%�c�w#�cچ<���sےJ��o��*8��cOk�;�k!��M�����#�ѿC�����r8i񍰦��Na~ˤ3�=�5����潭qE���iV��x��=Ik�#"����c,%2��]n���m`�9�S�i6�U�n����C�W\:v�b���9�+erk�Vr�L(����֡�]�r(;݂�\]Jq��^�}s�g���S\]f�V�{{��O����~��W=Ǿӧ�(T౬w�7�>G����:4*���[�k��z��ҋ{�ѕ���΍��v�&�^!��.�6y��c@Ë�Lnv��{�+"�;Rj���.���lx�^;R�]\\��c��1��{����d9��t�p�is'��~�%Cٽ��R>�~��q�@�z���/��`-�ţ�Gk���;ϜO��Ł���W�ゼ�������lxOO1�l��y���
o�Xᮕ]kˏî���y��x_73�z邹);MN��N'�%�vyڈy�����N:U��+ʜ1ـ�j�����W�un^(| �.�ά���h��|'!�kT�Ϋ�a�<pFru�	wZh8\�J���:�Y],�;:=�˾*�$�̩%��w���;\�JP��]fB�������JB�ۙ���<}��An\������_5cе�o_;�>��)~b�ٮ�[�_t�o�4'd����׃ո�{v&�	�ćկ՝=y�;������5p�hgh�,����s�J�2`�6�Ԝ�ܖ��Gd"�W<^d�|�=c�R*��
�B�elW��F�7q��M�{o�ܝ)��u�v�#�w�=�Vڛ�����v��>A��1�=�&�o9St���וi��E��s�����ބǾ��5Չ����m��(��_1�UWR�8�Y�ٿ��o���Xo{È{\��F�bOI��[{m�k ���v.۲С}W��3а����a�^	�Mo
��
P�;�\��+so��>h�9��ĐC��e�\���zt�!��#2�n��^c���+NH��@�j����<+l\IӋ�����BZ�fop�uCn+G�%9ױG�7�	^
AN�y��i�MV��VXq���yM�sL��o���A�>&����g���t������1b'�;�~�=�]b��^8�+9�'�#��]�|x@���N&<87=Ӌ��l6����~ws��j��TcDk�*q��Y8���	��b���F�����m<��=���E��t����/6��Wˬ�K+3>�����ke�(l�'���Y��6'�&K��w��U������Cd�=��f��β�G2z^cn��j�Va�Xw�̊{Ӷ-��K+���i�c6�khR����,yN�T�{%f���RA]���K�r�.���)�/;N�Jd�z���h7�X�ƤZ��7������9�|�ww�+��S3,un�\$�ok���ёuj���	U/h=���˚7�NA�z��a+/&V��e>���(�R�r�{[V��3޾�^����Öl����i����v�2+�U����x�H�2��_7��x�Hw����蠦/.���&�h�̠��h�f��vc�x򹓓���-��Ix� ��� ���A�N����]�9iDɳ/��)��b4�b�[V:�4�@h��^2ݨ�Ώ��l{���CN����-�A17����ĥ�w����5*qU�:��p�l|b�^ݪ���ϲ����dղ��U��d�Zw���t�S/�V�R�����i�9�Ԍ����Q_4ѓ���u��{M�I�ޜuӪ�/)~D������[������~�,dfv�.2O��@][JM�v���:�!3g)+���*�X�U�����Z�WU���`X�:qq�(��L�$�L�smL�1�W���2�ę�&=YT1�Z4l��g5vw��M_d���+�7S�?a��dc+�d�~��r1�>�p ��c��rU�����o����^�:T�y�rv�r��t��n���o�o8��{�ۮ��s�2rd�^%W63[�{^��ﺍ�⽺�Gy���Siü�ԃ��YWG�t������{�X��z��.S��[��=�0נ����"�ϸx r�����!ki,�N{�����5�c�g��ݾWPbU~C�,��ы���r8��ɡX�hUk4��i���s/���w�<�����~'�c�u�b��8�8QyG��~{�v�����S�d�/&p��F۫�)Tyz�V5W'y�3w�������Q������l"�g�Q�ea��!�����Oz,kegI+���TI��{%�b�Y�M@�["sfn���{���ޟ1!��PW�450J�plU^N�q�܄���й�b��ׁ>����>��z%��7�2�$<�b<3�k*���z�y��zv���ҷ{���Bc2�Z���ԍ���Qs��x��淹��S��b]�K}q�<�ף�������^����~-ɝ�#*߹����-�O�J���4'da]��f�g�Z{~�4t�+r�YU��m�}��㣢ܙa�N�oxU�~�3��f�}�-�TJ���X�y�a���1���;��=P�kr;.��:v�ھ����W�=�>{�d��◼�W#5thUΕ��� ����tF/b,7%6g���T���VzҗnV��WY#k��c�NYL	�����Q+sfJͰӹփ4�R�0�G�r�Ο;U��=���_s
bW�a$;
,�s=�hcwd���8��r^2�RvǨ�>9�^�cXp�Ҧ�}��yU��2^n��ճz���t�w�ם>��nh㾿�R	��;Td�/�
ý�]jꮢ>>���������`2�yn���L03�U
��~3ڜ��W�O
�L&�;<Ι��;���z���֋Ȩz<�w���F�|c�c�(G&*��az+8�pl}�*.�9����h�-�qh�a}�~2�Vѫ��>�)[�UJF��/}��w���{+�4b�Z"f8s�l�}�G���]�F��w��U���3$å';�tɔv/���q�*1�r����ut/V�җǼ5{4�Tez��,Q�,��-W5�idA�*��޻��&�H��ZE�v�,�8���Q��b��-Mı�r�¤�ו0W5�Ƅylڳ\3o���j��]�b�e�َ��2�j��C��k��)�=������s�x�����"BE�e�=�{���O{nLʞL��yIL�]/��y\.�q8U��w�*�嚉��`��:Wd����bau�Vd�gn�<}�$ޒ�����ϯ���me�Uq���)�3zW�{��>�o��:1�N'Dx���5�q��빃�s���k�]�=��x'�w�խnxѻ��[�y��>�7!�҅�U����ۣs'��U�����'�";x���)vh<�ѡx�;]3�l�u��l�A(q�T��о�/(/��H�^��v���z�V=�9�OYlV�is>LV��>�������ő��`�T췇U�'"8�B4-w2�����u�2L�^Ӝk���5�\Peq�#���Ԣ�u(�-;u�;E�&��]/�ϒ��^�݉�r�k=��7����NS����@���6�&���*��Z4#�
.]�U`�_�$~�*h���*�|�
���"�n��7\s���-n�ݗl��]m��ڻx>��Gw��KJ7C�u��6��-�m�U��P�Ӽv�wj��T��l��V���T�5%N��*K�;��ec%J"�Viw����O��zv��l���mFޛ�o�Vr���Ǡ��k��q��֫:z󏞷�}�OT���O�%^�<�M��ڸ*C��k%��;z��ɻ�J�Mqk��>�|񛭣��h���V�_5�tG���i� ���[�M�#��g��E�|���.�D�����W������S�Z�����HcO��p�"��ܒqU2i#��>��*e���"��t<hV�5@^O�*̦�p�� �A�f�Z8C�	9�J�4jd��A����"�� b3��1����ҿ|�� ���Z�9N�Z�7�3���0�Z�$ZYݙlr��a�$�Ra������*��j���ΝL~ ES�6U?pތBIfq2��Ni�A�?��6�<�H��;�S�#�W�G�H��U/��_y�8��F~�`��f@Y�d[�� J�b��U�/Ҕ	K�vB��s���sƔ�7����?���HƱ���[(xN�P@ER�TwE��H��1�ș*�,!e9�<�`������@ES6�h[�sM�w�f��h�od��O�!)������/3�?���i�2DU+���&&�C֚[�?���5��X��t�Su,���>�2��ȷ����mZ��<]w�'��xq�=nÐ "��� !�������gT�ڷ�t����C�!�QT�{Oc����N��.ٍ.F���s� L���c�"�`��q0>��26H#�\t�QH!jHj`@���`��׉��2�,�>�;��@��~�3Z��V�/0�{�
*����aۈ����@T�}gXL	[ �	�|4~F��`|�F����0N}{�:I�����q^���YD'�xw-٘=�J �������#Ԓ�%yz}�t�@ "�%�[���>�i�c�#���Ԛ�7h34�N��S4���"�@MgR�{ǗnX�m�H}?��Ww���uҺu�TT��o*�7�H���d�n"x�mS��9�æ��r�Ad	Qz��$ �*����wG���5�o��T��RlH3�ttHl֬Y�܄+����9ԲhA@A�$/fY������"�(HL/t�