BZh91AY&SY9��p��߀`q���&� ����b@��    }�-���h�(h�mMk@i�MV��k6��Udm�5"��5��B��@)Ehbѡ���U-�5Tҭ�kV�؉��(��sa�Zb����6�j�[VL��2S��m����V��Vɦ�j�
m���jŐ�U��5[ZȚ�Z�R�ka�U����VM�)��}�/[T1BԖ�2L4�ę���&F*@�m�l̈́6Q���k-jͫhY[Q*l0Sfd֛lJ����kZҥm�im�)%�i[,�ٳ�{�SZ�mSk�  6�>�V���@�mtWwV��@+��f��@�E�ݥS�6j�u�jݪ�sV�eʹе�Ҷ�a�����ZsQ�5 =��,jJP��f���T�٦�   {����
T�{^:zSt�R���z6&ն�\�x�zb�Fw���S��+{���[joy�*@�&��s��f�ɳw����˪�5۵���̡{3F㽫m+l�f�ml�%�Z[)Qo� >��K[lD}����j���������a��v[����yYMU<�w%zʕ:˽���f$
����ŵm�*�<��m�j6n�5��P����I�{�O���
K�VmkEm�Tm�V�  s��T����k���+т����}}1-�J��>s�]v��z�8����J��\��>���ۻ����=�V��v_z��vʯ�]4o�}�W�ݪ#m;�\��:�W��礡mJ�Dց-$V�  ;�����v���Wά���4T���}�}��_J�뷽�^��M6��������&�ޖ�i��>�����m�g�'^�ԯeXmm�<^�9=4��˼�S�Sx�͖�Y�����ִ0_  n��zݵ]]�gw��J��[M�^^���w9V���]�{=p�+�^�k����:�����s�z�]�w@7��Wh��쌣l�oz��`���u�ۼ�m2+���4�d��j�ckR6M��n   MϷ�Uk��Q�=kWf���^����[9���zk�4����{�U�`֝�X{ZB�2�<�{�m{�:�=�;�Ӫ<���]{��l�W�/.ƒUk!�iT!D���  �>�֦��h��)磧����p^�[��ު�� 3�9�TU��o�k�N��t���U7����w�)ת���z4��B�6cEPl�kL�  ן��׽����.�A�Nn�P��TUܯyѧ���w���
;ʷ@��y�Q��{�-�W��22cV�Z�m�Tď� ���vb��{�sv�@{o{�[��L'�����Qpw��{N��h�x8�X����:�:;����G]ޕ�� ��      �*R�0#  CLL S�R�T�� d  ��{%*J�      T�U* �    �@�HO(2�2h��R�ުcE<�FP��M3H����|����MM?���%���>�����[���������>~�AW���� *�
���P_�
 *��������?�O� �
��Q�. A*�����w��߻���<��dՀ>O�~Y_�W���L/�e� &W�W�S���=e}e}e~_X_Y_X_X����=e}dY_YC�=e}`X9�����������=aX_��1�+� z�����/�/�����������#�+��	���z��Ǭ��+�_X_X�������>���W��W���C2�������������Yz� zʈzʀzʢzz�z� z���`�C� C�XUXTYAXYXQXT�e��@�� ���@��@����P������O�XAXYX��TC��C�_P=`P=d=`=dD=aQ=` ~�_YPI��QS�S��D��S�S��0 �� >��<ʊ�� ̂���'�(0z�
zzªz�
zªz����*�D=e &ES�}dOXC���=aY>�_X���<dX���=e<`=`OYG��`O�@�aO�P�dO�d��`O���}dOX��2'�3�*zȾ�'�!�z���}0������Oo~���J��_9S��QI�*�����^��!���*�&H̤i�˝�8[Y���MUލ�-��[ѵ��ʹ�L�2n-��IL�u,�'�,f�Y����Jסk�5�E�̍�/mܨj ��2Qƫ&�਩^ɕ�$c�WD<6��nw;v�۹m�]�Z��A��+r��`��V�FeU'[Ka�'�F�m���YzČ1��\˳{���[b�̱�ֲ��;�;��e���j���*`c����!C��|��]��*6����u�������:w��ʊـ�ɴ�L��I�DlTrC��)]ń��1�O���yyoi镏k8����,ݗ�6EV����kX�R7#R�f��^���!�%�h@0���-�U�׋(�X�+�t,4�ͬ���:/[J�`�Ǌݴ#�V�[y���.2��2Lʥ�Y���;��J"�ǋt"7*��*A�q%��0�iAZ8�a��f�V�#MIf\Ĳ�q+4l��w���wgY�t��5��̼4�l��(P�ù���爽����� 8�nv�MY6327m�7I�"�/tm1�p�+ra�l��Y�d�BM]cr�R�$d�l	�Vv���X30LT�	��*�,چ���iu�]���<9�����{@����C0�v�Н�&��kv0��"�4��F��~5�Co	�̻���f�-�e�H�Ԫ�nR�n�����x�Ɖ�N�9J�ic����E��"�n�����[{�Ll�sxk*��w�1�
�Z�' ���[u��FS��r�Sq�Լ������Si�M���܇�:�טҷ(ݬA̍b��ȑ
Vfv���T*V�r��GL�>�V�1�6k�y�o6�8��,�.V����E%L�E��1��FûқU�MRr�b��
OE:ڼ[�r�b��ݧl�%F��$�����{��1B���ʩ��PX��j�5Ra��|~7z���(iujӴ�u����xA�jۦn��)�(����{$���	qW��y,ţrG�Uf2Y���d���`��E��	d�:�©��^���]���Z�r�Վɸ�
J�����/,YY�>w����%�9b�޼!f8q�,�qU��͕B����p̳��1)�Xn��	e=W�
֐���t��F�i���F������v =�+7P��6튷g�L䘲/���d:�s��$w[EVpd��^����X�ͭ*�i�oر���[7�ƦM�����z�A�C��;�P�R����jh��hB�n��GV��&-wz��B��M��-��
��]��ʞ���9� �gm�-�ٹ�q'(��kpP{�ۻ�N���gPC�$�dn�Ʒk2b'X�3L�x�Cz�Y Xoct�EF�[wڭ˻�9
�]����,�uJ1�a�I�����n��[�W�ͻ�P�*��]"`�"Ll�6�i�k�+F�9�����[�ӌK��@��VeP�0d�0��r���".� %j��JJ:��9��g��ʭ���mZ���+Mrh�64%����R[�P�0m�oR�ڵD`�p�*P�6�M�M	P�62� �*�;D��+u��*�ˁ�0���h޵e�(Ѻ��	��"��IѼx3��x鯋��2A�vp۔M�������Өc���4e�Z��V6��W$M�ڦ��нh�lP���@�[5�	�EnYVAue@iF()�[��z�Ix�/V�Jz&T�����w�Vf1I�&}������ھy���W�;��n �,��9�	e�!W�N�#c���{����V@�Ư.���o�6�K4���HQ��[}Lh��m��IW�nM�ŴQ�ہ�����Ҫ�NމR�4B!�Vl���2�b3jVf�R�#6]�������h�ݚ�YV�حu�=����I1!�gv�!,��YxXR�;KM�N����LBeb;�J��72�A��b.;��U.��XM�������˖E�4{�:
ĀԂ�Շ^'���q���:�ib��x�I��g
{J�)��jb����ə�M��H+�h��u�XT�z�jO�����-Y,�t^;u���,B���уfV��W���h�n��v�E7(,�k]��Y���s1�U���O3�Ӝ�>�I�8lf�����x>����׈Py���4ʛ�UÄ�9Q�����"�6�j�n�Tƚn���+�;a�ږ7n��4���{�F�:�h_2�,=�V���a.{j�`�MbۅA*�4-�M\VM�A�d��F	��4�oh`h�0=���2^�����Ʋ��	[�jR��6@V����-\��qR�x[WU�^��J3��s��^3w91�¢ܭr]�;�j���Nm���P�Zȗf�[�� ��r���n@
ˤ6�c����Yl^scz�j�3�p��S��M�����oA�7���A��q+M�N,�7�m�8N����zor�a�rΙR��e� ��sm��ޙ*�S���>z\.��%�;�����t(�-zܑ�$(�oAI\Z�n�{RkAdr�n��bwm�-�[���-��y�0�[��YA�l�l
�upT�"��uc<եx�7C�[c1[�9s��sGI�I+����=a���W>�[�/�@r��ƃ��r�A�M"�`l�Nm��f!I֝t�*��΋�6@�n�7�a,�ȓ0]eɊ}�Ͷ�I�úؗvF�0L�K&��?�V`ڏռ�y0n�nLz��;`,1���6�\4$�/bSoCqn\!�-J ����g
�/nd��:�Zn�n�I��:1�V�Zh�䑆%f^=^�ԩ�A��+whՑh�LSf�0����z��z�ۙ�$��X��vV�U�����m`a�u�֐m�0X�ǥ��*m+5�^bS6H���FV��

��%n�V��yaT�Ůŵ�^���.^���[ ��Ԣ�[%�NR���L��Uݲm��0�i��r�:X"�0�*R6��S%e���EZQ�aO%��Ki�j&��ض��fх�5�g%�Dl��߆�t^V4^f�f�7f
��sNAN�Qu�\C#ћYhӂ��~�&��en\��q�uHҒ�;��!n\��#d�1<s%���5!ɕg�e]�����>6�M��h.�H=8��@�ڈ��¶��,�f����Ǣ�R@kư�]��Z�SR��.^�q#��J�oeP{�Iy,�eǰc2�]D.Ց�V�`T㙋��������pV�Cm^��{�-+i6΄5#�&�[@2�j^U��z����w�����i܊��1G-#�l+J����nL��#R:]i@�L�4AW���*��t�-Y-3^+ҩ�!D�D�Qb�=��^�l�bX�<r�Z�
V�;F0�wb]`Í1�/�1�����{�a��n��c3j�ɦ����*�J�R�q�v���ڋR0I���[i��oa�V�2x�T�)S�֨���)Z�9ޚ��+�Si&�ExÉG[�1�����F�-�֥�ϱ&-
f9�$/6�t�i���銛����2�|�m0%��yAn(sfB���n���I��-�d�]k�^�kAX�br���U���6l����$xo僘I!�����M�u�c�<��QBތőU�.��������mՇ�B�-Y$Ǜ���qi�+V!l���hQ2��zh�&T�R��r���ҔP����T	��;G1�5���ͩ�e^ö��yA�_e�6�L0�6I��&���F�"eϗ�P��&4��bE?��� ��jYb���ndtݓ�R��9�	�n��OK.3�Y��Y��R�3I�+mˠy�l�-���|{��w�Mˉ#S��20~td��L����%�jq�9���l�M.X
��]ś@o�m ��%fR�����X�qI vޣ��쒠9�Aa���ͷpfT�$�f�)=�����E��m�Y�2�i����!D��U�6��j�v� ��+�M�ȐT8�+�9W�d��/!r{���f��D	4��C-��th�R/R��f��&����),���	ZƒR^�r�R)��f
�L�׹��P޻�n@NBa�+.`D�Q�b7n,%�����,=
�������w����ە������o52��^+a��҆�%�=�����u'%iœ(㠩{i����L�f��F��7�w��m�HW,�&)���j,K��e��9
�9��R0�ش-r������-ǿE�[r��&�j�4�Q�Y�K�0��Ż�0)*�E�2�/j�"��	M!<N�
OKq������@q�j�me�l��d��lͫ�Ia�2��Y�R�U��^�p���Zd�In�k�f��;Lna:��1��Z���ל����ʖ��i-�".�e������&����vv���Ӑ�ODZl�9h�qm�"�v֨n�FRyTF��2�ԭÅh7y#*:N`�md��L�Y`�S%]X�[��J�G׳0Mؼ{q�p��ax���x�
��Az��:́���ɨB⻅�L������SNTu�Q˳���f���`4��b��Yy-��Ďmj���un�w���IL��m0��Gv����Fn�ȳFDďml��/+UDr�T��wN6$y���Y���C�	��n��Dve��Z�ϊb��L�w�=ag'��u'OBսQ;����&w���&=w�/���0�4���Z7#L䬵���Cswj=Ԝͦ֋��� #��8��pZ`���땦�A�m�����qQ��\�=klރ��Лu����lD�;c0�3��J,U)ީV%vB3v��(�ƀ��i�AY"�z��1f�N�5�#�,�A�<V7�u����-[�:j���W�n1Zf�#75Ef��
�p��k�U��25�DW�q弔XIǷ�\��G\�����Tm���`����Ih�Z/ �U�P{r:��mL��h��E4´1R�E��tm�n�[���Qy���,��n�Mǻ,�ۃuҭ�]"4��&=��h��������@o�އ�v��D���Ӧ�j�sJu1a��13��m�xv;���Z��p��j�w}�(����GѴ!�q���otՁ�/oZV��U��[ۃ��=.��v��!V�E8���[�h�+�V��9�g��ݻ;ܖ+l,K]�k*fg��6�+�����<�y�ⷺJ��5k�][9��ɻt��9|���������tom9Q������CE���B����՚�
��B̍��)�x�4�sD�{�@ܱQ}Dɴ�:���(��L�X�󻭣Z��Ƀ�7&�Xh��l�=�SD��%�:ګ�x�ms|������ԫ6�������k0���Oic3j��B��L�,�w(f^�72\���Z�!�+V���X�Q���mې�����`2ty�{MV�
��]�����Vc���t� ܽ_&���`�P�u���x��"��w�R6>�wX�Cw6����>�p@d"�!�PFb�͙�R�u��
���5)��U=��9w��!l��µͭ��E����f�f���2tᛪ�l(�zӱ|��{�<���YVUm=����t���W�Jݪ
�)�+v�	C�Zn��{4
�5:��d�� .���Ӵf�4ʙ*]�!w�K���Ӹ�����VU:�I�w����]&(���W�Evd#9�ü��1FL�f�
Sp幕���d�Y��kf��4��L��hM��N��K5���Z�a�Y�b��EaݏE6ͤ�G�m���L�aLsۤ*Ӯ�b&�h[�t8��_i�t��9��� �˄�J��YJ�j�hB�9���R��������ZE�h���;���c�am��Cn���1[��Σ m�{��9r�=�k�*ݭ��^�cx�_="�!�6�
���n�U�7SՔ�=ɚ�����Xycj�bи����A��*�e�PY$������n`�L\&�/���sy=K����J���|3@h3�#�Ln���"�N�"�(��P/���j��V5��:�����U|��朄X.�[��*�*�FLע�b�Y*���7r�m(3��+P��Й���*Z�i;��Dje�dܣd�JPV��q1njtƬ�9[Hb-V�Ԁ%�|�i7��ZF��PE�Y�:��kN�E�f
͝�D����f[�{�*�p�^k��-Cf��;�]k�̚Ri�H��U��w6,M��e9x��v8��Y����3+q��X��H�Q���4q^ā��¬�Y��U����[ڬ"��k4�f�&ԲM���H�p�ԩH�?���ƽ��5CC�[Sf^٩���GI��S`�by�$��T:/3(`s.��	a��Y��F��FP�`"�(k�a:�4�m z�O%�m���Z~Wݪ�t�f�jX[��&̵MnV�f�)��GJY�4�d]\��^������F�a�v�K�k]fǰ���e�S6nP�d��r?�D������Z�k- 6��\W{l�H�,�3
[2��ab�jPݔ�`\����t&iy���6R)(s!�h;�^cv6)�h0uQړS+$��m^���VuG�����x0b-�/��� ���x���
�X�ؾ٫r�m��(,��$f3F)]'X��tk�f�>��v��9ɩ�����f�����	�x�H�L�\!1����ދ$`���PjWQwN�gj�c��M�AoHE�$��_
 �WuwQ�.j�4��f�ɟS�gi=Ԋ�nj�O-�9�wNR�Ź ���-�>�L��رӳ�	�ZҤ{�D���XvoZ9T�pO9J;�ox֢��Z�%nV���1]��p�ks��o	�᩷�c��N_gj�Ap][��F*�V+3#yX*��pJ Ucw�t�{��cmo]�2��5�����|������X(>^���� eo��
�|��N���8��ۋ��rO�̚��S�ty�ML˟vʻ3�˜�851���V�L��4�ͬx��<ٝ+�*dCCU,�f�ղ���������sneA�ր�m_E�z��T�p۵�Y�: �/4w2[c¸�L6���(�囥��
�$�[L�{I�W��;j�}�X3SB&9ǂ���V���r�M����F�h�0�tJ�ʠ����n�i1�+�����6�=1��2��`g�tj/��fK[xe��s.Љ���-�1��2tY��-fJ�)m`/U_S\A#T=��$���
�\)fS����/tj&�S*��/Cy���۽.3Se�o�[�m��/�L�k.��F/��-@80ynj:��p"��Y�{�������m�c�H��8Y��(q�w�a;����5��K,����n��f�Yޤ@��I*���� ���Y�5x���y���o������-+'��vts��C��eй�hj��U5�3�7�sENҊ�&��5�ǩ�Tɖ�T.\�u���)��8ܱ]�v�2oj�S����_�,���<��� k\�G�+�U�h��橚�yS[5'�d8��%=Lq�(���j,��]0�݆]�EG}�4eZUҔ����ΛS��P�7�Y���"V!9��x8㮖�:Y�pa��,Id���:�[��]>����V�� �s��[�2N��݆��FdԠ�ar��,N�O��O����e���f�����Cu	�\}W����h�Fl�=��`J7øĔb�����&�r�2��8G��Z��wg�#�wU�}�s ��d���k�<;�tN�-b��9q\�Ɗ���IbҀD{[�N�[Dc�V�Vf���+6�Yr��x=w�؄��vi�o���Q�jZæ��ȋf!�{h�/�|O[��b(��lWU�z���{��ط�6c=������)8�˧�5HMT2�u�]ܓ2w�:_L�܋q�d�٭eΛ3v��w�dY/`���Λ�������AN��$s��k!��Z�:mS���+c��a���_on�5024�ш҄�8,y����*��2Vj��;��cVX\���:"b&���q.N��x>���jĻ������*{Y'���G�n�V�dO�m�Ս�u*o_u��;#�"cզ�']� ��])���}6!�oMoJv�G�+7K�(܊�,}f����+�ڼE��I���u�����F����!��]V �\*�W��!Y|�0���M�:̮�����V^_��;�2_kv��];���ՆQ����]����I^ay'+k^Ar�����Wa��Ӑ�G��E;��i뫢��ѣ��*���4��{Ma,�P��&;�k�B᫻��p�̕�$�����\2��z�+��K"1�7�|�ݸ�*8ؒ�u�Ef�SC�DL���m�'b��Mo Z�-O����i��}���V�V�h�q�K���6T*��ݕsW[�Ƞ�v�1����j:,���
�-�q�BaD���x�$u��ۧ�p:�[vwz��G'}�Aۛ|�5���%�:#Lw��*x�k���3x�4�:X��S����|X��LV��$s�*����F\�7���w;&*]ni�����u$re��;���u����RQ�f�������L�~Ǧ���W�򃥙8vs�)1�*hi���Z��q
2�ۤ�ԩf�Fa �l`��ݙ��7Qv�lu�i�u��e��uI�ظ6Q.��X�5�c.\6�\��O]h�)���b*/��/k������h�lk ̻�3��.���$Ol<9[�V��\���[�+ɚU8h��]fI�JYM=:U�7Y�)u%,�2�\|V���x��x�6a}���\OY���Zv�T��lسy��N`����Γ4\�fG����OS�pB�wU�Ydkݖ�	c%s3^�
��#�v��Ek/�W�#��p��]n�c���]��'R4]C��,����f���2�.Lq<���hU�����j1T��M%�W��
[0�����	J�41?�Q�Ҏ����#	��1:�h��Tʦ ,�7�ss��j�Z����S���oP%�r1=�����Z�ܱb,�or�l,��=��)�"����N�[L\
�;�	s�D�ve�a\���e���R�z�V~p�Ox]�V�@m%��D�D�N�vgZ�n���~y������*1���a����ݺL�	u3q��aܣ}k��\Q�YHu���8w+u����Lb��ŀ���0lcn���T��ɞX��AovWN+�*��!c�B�$��Z���;�I�Y�A���^��	a������k1�x� �d[ڛF�;J�3S!е�\�x*�n�h,1؆MȻeq%7���m�"�7+t�TN�%��t`��d��wS���/,�&C�3�*F��D}x,ݍ[O}X�L����I�[�/d��@�� ��M�j�����LP�pM�뫜��Z��+/�+z`����6:��g]����b�6e�)��!;aw\x�V>[�'*����F���dx�ۛ��|;�0V����f�zã\w����:k��֯�����fr���zy^%]�v���7M�KTΑ�����]���%G� n��9��|�9�\w
3/9����ݢ�k
��	4�t���Z�7����LO�3�V��Y+�=�#8):�����8x�V�����:�-PބM��w�"̼Hv��?#n�m庶�j�B6���H���d񄧲�X[2��De�4+&s�g	j��2Z��|�Ҽ�Ʊ�gP��k����O`��I���vf�Z%;p����V���l}e\�K[|�9&bn�EK)*B���镈Jʷ�b콾��,�TB��1�N�T-E��2ni	^&᫴��᝝� E42尺�»z�N{.>���Cܴl[rj!�����y'X���:�O@���E�&�wt�C]�0��9�5f����Fz��v��T⥁az@y-ŕ�ݓ+u�ʫ�ZV�}�ӛZjf���̹�&#\��vާ��&��*��xcY��_{8JL��ڵ�T�߬y����s���&
c5�)��� ��;Ñ��q8#�I��v��u8_]�Ǽ��:�MleŦ�(�1wH�����N�XQ����>�0����#���'2vw���7E��X����1q�����R-���\Ċ�0>�X���LFm�Ъk\j�v�f�E�����k�K��r�qo3K�u��w�c��ꔥe�gc/5�>��j�'Dr�{kD��*��침

�G((n��ַ^��)��x�Z�b�ۭLr3����:=x��hD��ٚ@V�	�.	��X�I��n� �.Wc�4T��o49��N��r�	CvKu�N�1_n�qn���%K��.�.��c~�'<~�]&�\"���*�w��K��&��."7C�I��wb0R��}��ǅ(�����;ݤ�
+��[K.�6mv�;N�Ñ��Q�y+s�'z��5��X�Yp�ۜn9k,V��Er���p��i��a�쵒�`CJ6eP��$���oq�˼�)!yݰg|�>P�^<���.���[�KT�k�m�'.Ո-�`u��K�z�hŦ���ޅ�*�!#0�&�{/�M}"��l�E�7{�T�����_-��YcMiM=!,F��]���7�i����m.�ʹ��� �NVq�
����J��>ɔ����ާ��+p��fb����Qd�<L��	2�'8fD23I5�؎R.S�dJ���|��`S����V�^Qpor�U(�"��U�V�w(�o��k��K��[xU(��p	��e���٭��ڦ�ou<��-��׮D�gY-A0,�%I��1A��.<���wҾ}�p��}.)��Y{9���X�W�Ю�愋[_e���jvR8�.E�k;��6����$E����sl��੍�*�d�I��ib�,�5�:@��qrճn�Y3�!�d�gr���I�Ť��W��<��-yS��hx��]�O�%�\�Q�7�$��)V6��Ǹ��>I�x����Z��1S�I��3�4��M}�M�VN�l;�q�i67�^'}�fQkfp��AP��7|�j.K��Y�d���ӳ��]�� 
{j���%pV.��Ό}G�M�����R�&[���P��7�l�{�qqª\�V����CW��쬶����L7b�V�7{5|5dS.��}p��-����kV�j�t^����S�n �] ݶ���*�Ol��ݷ\^es�8���xT�Z�aS)J�=E�8��(۵NB�ksʩ����\eaV�|��Ő.�Q�޼�N�/�:���O+�.��"�����Ir�r�< �4��Wv`W��^��լ����Mv�͕�o#�u&k�AVm�6�N��T�p|{�>��P��vNc��9"\��1v�:ވ�#r��o�v�{�˝S3b�isr
�J-�Hi�����сœyqT6�]R�S�Wq)�M���.%b߻M��$�9	/��^�m(�N"�9��5J�Q�ZN���lf�]{ۊwt�U|0��&΃�GUs���;:F"��.H��(����L�m]`Iv�[�1n饳�h������<�3Jw�s/ �K9��J�s)��EZo��ˮ}y�Dq����ڵ"ɗ�{��V��tWw�$�͘��a�����wl�1b�����P6Qɨs�/p�Ǳ�Z��^$x�Tv�=�aZ�-��Ż%�q�TN�ՙ�I���aOHi�&��i��ob9#�VW�k���o�%ˡ3@���,-��t�w\�����	��[�_X�RJ\�:��R�L
D���]"���1wZ���G#[w-fC/uU���J	X܄t�M�_�-[�X�L�$�]kY>��Y�\����;y����\�0�~���Gd��_ea(P5@m�K���d�.���7Z��W�!+A�J����Vsqb/`���Iږn��o|1V��z�s�t�rQۙ�`d����X޻w�X�@���bʂNP�1*Nr���,���`�I,x�a-
3kAt�*Ұ¶�0ꏑ[r7f��%t[��{ҳt�R�L�y��:�:������n����dC���,n�����8�,)��ۇX�_^�Ή�;���M��ѢS7�wX����Y�WKO�uө)foө�C�����u��Q�;��s����d����yge��kw�eFOXba��Ps��3��ٹ�.q)#CL}��pۨ�7V�Z1<#��C,GP��8��f!#���1�o��B��b�r�G(j��9GIf�'�����@�"�NY���nv�,����KdR�2ST�@}q��ٱ�K�)������&!��^Lx�B���A����S�"�]X��I>ɖ9�Dg17�]�.գ���շ0�@�8՗]Lg|a�3l�u�hQ���;���FV�9�kn+��l+	�0�r�bp��T�8�cP�ǯa���V��rj�R��5b$�&��sv�P�b��\q��AA7M�F�9��{�He�e���8L�l$�u�ᣞ�n^�[M��� ��8�P��I�m��Q�+})���'(%{����0��yy:�
��=�t��}�ʹ;yS�we*Q2��r�CZ7&�$ɕ�GE��.�7������}4P�GO=�wM��ql]��U2u�[��]��p�}��ǐ3���t|kO��g�%�=B퉟H���0�B;�J��|%&D�wŇ��Z�br=7z��ם��M]���%��lm��u��̮M	��QP���ñ�N�m;��5{��CƛU�"��Ot��(�0м�O;���t����&|n����N�I�=Yn�z·�nl�,はֺ�e�]�����"a��
ۉ�&�Σ"+��w>"p�`HϚ\oy}�{V#[2�+f�S�� �A�CM��8\�T�߈^�z]�p5����;[a�x��Y�GQh�9k3��Ľ�ƺ��-�4<;�uzΌ�ͨ9MK��H(M���=MPy;�V�F�v���v8V�z������q�R�J{4�wS+.}���o��O��zܕTnغ4�I��M�9�a����4�Fxt2���=3q��kB^�
�1�����,zH}���f���!�%��	$MA]귙�k�SPj�yV������V�T��*��(��I�1{e����D�l�ջl�{��N�(Bl��O�abt��P-H^*n˫X��ͣʷ{ju�k�,���(8��W>��Y�]w%v��<�^����KxH<ۺ��˹:t�3�4&�Θ^	��y��`Σ�`6��Iqz�U�)طM:0Ty����Uľ�7t�޹��}Lfc�:�P�T�Wh��Y��.�_'0-ᵘΣ�g@����+t-b�'B�ٛ��*�9�.b.N�f��rf]=�u���R*�-8Y��k�n|0n��33#�-�Z6^W��;8����)��u�u&�&��ky�sj��MJ����m0��_D�gL�k�ٝ�9�'�����
�R�n^�W%���嚣�	�Γ֩�)��{q��]�������q
F���{�4�Z�w+3�&�ʗ��[�H�]�0C{˞��ڞ;���v���E(��$n�a�} �Q���k+D��u3������U5�c6D�&yX�uF�{�7�d����&�"�295���.
+"�U�����aDP��5�Xm$���9�qt. ��UG��ҡN:���B�d�dF@�!+2:�aL�n���ج�M.��(Y͢jYh��$��4۲��"�Ek�;RK.3�x"�X:�q]����M(}j��5���_[�~M��ww�����/����_�� ���Q�N�����DTQ��7�?���|�����~M�5�?9�ә3�f!�A���ǅ�f�������I|R�r�W�V&�k/AO����r�XP�#{]9�}ZN�Ά �5����#�+{�u�w�i]�o�0�u�2�ޮ ���a6��B\�������4�iH�{cU��MwX�`G�n�ݻ�R5�K8{_Z�,�^�<�Qz�sX��#� �bIglH(û:-x�;��o�������E��kɫ%�.�V����o��:8�ҁ��dj����]��r�����t��Fv4��[�0�[�����R��X��)v�7jlѼ�F�[��dٓ+�vC���WHR��a$������koFH@���sBZN-�L{�w��#�[��F�������'L�M)�˦����2������a-��ݷ�����.�Vu��,6L��p��؍�H�<��)Iu�n/��J}u�ae�x��ټ����'D�;]-����:�j��f9�{uH2�f��;�1��Fe��Ul��a!�Q�mu%�С�Rr��n�ya��S�y�(ѩ��+�Vg��2e�벳^�eVB6 �ElJe�A�R�
��N��]�_'J��Y��4 #���\��K�d��jm-4����ح���ĩn�XFu��+GB��.,����M��+����`��U��:�W6;$V�r��i&��-%�nd?kҮ�ࢤ3Ri&*#۽�g`�a�i4�.����O8{1�T1i-f�T�m�d�m���sG�1+��i<���ջsr�e!d���ۭp��ֱv6�^/�� ���,����-�2�:l��E�LIBnk2��SY+0�*'F�F
ݒw�U,��
��u2��1Ġ�l���R·��ǖi��J��jո�+{���3p��Q��'����x��*�Y��l��4Ƹ��ݴ���p��h���w��F�ﳦ���V'w|�nS�fb���fG�Y�S2��4A�H��D�L9G���&� {���ب��G7cQ��h����U$pƝ��Mkbr�84���v��B2��b���[�!v:��z
�R�"p�F�UXP�R��y/�.�6��/j,�Z�FФ�]�a�U���m-�P�#hWhU�G�u�V����.֬�́�Y�rK�z��un@>�A듶Kۃ��CR°�b`��vZ������ǅ�wM���9E,�����E\Bya#�tph�CYA�QwZ�+_v�Ww�;.�o����h�.�@P���N"M��/A�X�)lo&����X���	K1�ۺ׸�Ů��r��P��f�T;ί����2�O�z�ao':8�#�k�r�]W�NZ;`�R��Ρ1��ũ:ʁ�W|�N��;�EL��t�lϊ�����Tۀ��lwZ���1��q��f'pU���#\\��������y�E��`s�#��7����e�j5������%L��4i`��3��<>����+j�b��{7%��*�����:+�=�&�]a�&����nL�B��/����ڴ x��
p�@*�Y@f��j[�EWBc��.A�f
Ml�!�:�0(�غ��B�;��*Y��6�Yj�u�P�X�� `����k�l�[���r'aRKoa���uu�|74�C��6�ͽ��|��q�����[�f��K��H����D��8��Ă'!<��y���7ΐ�h�0�459�ED�^.(Jtf����c�}>ם'+�j�ˎ��'��d�dv��(����{3\ ea����j�F��6�7k�0��1rf��N�����#�M�-n�
���Q������;@b��{Ɔ e:sGZhh���*�5���e��d��չ�Ea];�Q����Թ�y���ز�nb������e����n�s�T��I�|��;�unФ�먻�Q�N&m�k�w"]z���t�wB�Ka��;I�� �kOk4#Ǒ�-�.6��j���eDܒ�������-��; n��Ӹ8Q��anA}�-Ҵ�V�ӯ�f9��劆�jt����7�m�	8�D厣o��]|2e�)��z�֫��J���.
�_.��7r8E���!�k�p�Us^ؗ�ǔK�K���4��c��!wP�\ ��r�T��:|��`����a���mF��}NH'zü��pAwb�rT�0�(:�	c}Y/*Y�.GT�5C5-�:b$N��.�g!.�m���3F�0�����6�+[�V�oulTE=�ZFl+٣��n���s=oN��I8�b��DwtXյO]B�^�S�:Y٦������C��������u�,�8�D���>@:�Ṫ9���5:խ`�+5+xw�m�t^0�Xr>q7۲�;�̦9}M�v��M��*J-�����sz���`,��<�{��P�7��_2��V�}�-v�Y�'X�]
�l��cf��%�fi��SV��o2*��]l�FR=��+81<� �l'Ǔڀۡ�)i0��z�����߃)��ܟaǥܣo7��^��r�7u����~%'���Nk�:�4%=�)�1:����^|��0�P������R�[u�ȭX��{ZM�97EX{nF���U�@7�c'V_,�P7��n]��=��Wm�2��ޒ��qu��D��@�#@�C3s��:i�w��b�\=5ۻ�s;�q hϦ��Z�N�U��e��I�
U(���^#�F�b�a��Ό��)�._Tҷ�ٵ5��$<]K��<�r�*i�oX�6F�4;��=5u6�H����mu͖Y���ݨS5#��2�/U$[��P��Cn�T��rҬ���0nt"ˤ�n�£�q��
O10�y�լ �q�BX�c�o3��Dtx˧W��-(�㔆�(*��\�N@I�1g7o2���!i���b��V�/��.�/��.� ��9�j�"��џ���<�$ڬ�X�f>����&C3(5�i<H�Z��ݩ�V�E@�x��y���"���O�v��oU�H䄶��*��9�����ަ�;Ϥ��]D=�gUNlӲ�Ճ�ݡ{��u³h[��u��f�;ۤ5bȶ�3w����0�j��H�k�-��G�N&vǪ�.��`˱�)	��Qt�u-�{��u��Xr��Хy�,Gطu�{��	�#��9x+0S�,t��?ma\x�b]}>���XF���� v����s[=5�˳o h���buo*r��DN��='��I�&j�ʻz����'N��:�k�H��tE�ˮ*�.u9d@W��`3�c�A��V�)���T��5»2H��,�O�� Α[�s�fTW�Q��|�U�1N�^f�#��Lܳ+2�:V��A�c�82m:2\��,N��^<tYE>�rv���x�<�Ŧ�MAb���8��(C}�K�S�]�j��c�]�,6Z� :�u�`es �ߣ�N��;��&��M��$���v���7X�Xr�fG�9�\�P���ٱ�+4"A9�l�6W.	>�v�q�M�w��,MsWn[����>a���r�\�}�7���r�Mxf�E�CոW�unbk���١�i8Oj��.�j�7H��C�-hm������^�W���~qA,�s�ﶦ<�Op�[2��Iݩ.�v��ɳ$1Y�����v�J+Z��X���j�V3�XzH�f�ʮq���y�e�[S�Z-��1�,#V�қ�>��A5O;!!����:�P׭�uF�9�	g<�;˩�A�5�����5�U�}�d�D�T8�ۊu��Z��$j�s9�f����+b�WV�\ZF�BZ�Kk�����u�WA*�����ʾ)�P�+���5�7�5�3�O������q�쉴q�1�u���_WM/+0�I��y�h`����Y.~�HA��a �PP��W�R�� �M�3�I�b�	Cm�o�]�9��J� {�\��lF�G�ES;r���ԭ��|�6��_+���4����l����m�|튅�`�����hj֊s��¹�qph��0�E�+�q�aV��S:i,�6/�(��kw�ɹi'�P8Z=�_VF�p�lל,E�-n"��Q��ڀ�s�&+�|�ܨhdN�ͳ���2��9e�ր^�=�N��ta�̸��q詍�t��&�E�ws�:�Z���4$����z+��L��
ҙ���^SG*9X^��"-8�AipG�W]�|c'%ḛ�M�x�;�eu����\��t|sJ/qS�D/�+����z�d֓����7\���%4>�uv}!l>VgBbu��dQ��c��j�Y0��i<�h�֠�vdy����n#}6
D	�s�F���1��M�Xm֘�^��;�0cK �XE,�,Kv�ޓ�#��t�[�Pf��ogj����IU���[t�U}�Fg)atlPu�%&8�[ݧ?p��0��W�I�G�J�1�7.��y ��c��Yf��8�̝�'��O ÷w��A��'Oǁ����v�������6�f��a;��侣Ogo��v�â�6��tJr�5.B�Ƨ��P���{��n�bQm��ٸ�n;R��A`æ,�cw�(����`�Z����nr2�Pάg�X�ُ��6tF�Z�]P7�NQ	C6]�]��h�7�k|��|�싩]�tilzY�:�q9���3��#P�nC5�5������E��X�_:�[9/�n�+�mѠ�㤮����3uG	�r�F�'��g�,m�@X�[�������X���L݀�#��w{�.����Z�Ӕ╧Bw恢�3{2X�B% M�eM���Gv�E5-^�EpE1��f>k(�09�9��kA�u�ρ�X��z22��qQ�I�ϳ��%�Z��K�X��(��;����.ȩ>�f�E)N��En�s��~�ו�z���w9�Eu�C��C������/��f}S�Aw�"�d�		m��� -�\�"��b�5Z��ld.6�ʋ��Qܤ������dT����Z0��x�]LM����R�j#��+��F��r��Y�(�Z��r`�a��G�Rݫ�J����br�w�K�(�����Ë�b��Pf:���A\)b������߮�E��\8�U�@t3>F�(��i��K{	�~T���V�U�3BuF��k��x���l�r �l�	�	w7^M��iv��Ӝ�J�K���uf}mC����tc0��md��#�����Л 鴩C�-��~r��U��v�d�����O'gI�k��+��|�"�7J��P�I�J�;��.���Y�2ZWnP�\d�\S�:Ƙ�ѻ�IX�.�
m��k�=�&��+U�5ր���Sr��^�֖�*��v���B���F]t�hM,!�"��� �UT�+	��ݦA"��U�,�"�k�Iu�l9���8Й��m�1쥷���N_��:cZ�7m}�Hĭ60\0(z�	Զb�bވ�:n"���a#v�Ԙ�י��j�o�WA�`����
Z���Ӕ���OI���_^���QM=��F���w#W�'-�1�$ަ՞�1t�Z'J��d�X�]3�������)ԭx���_rTժ4���w%�2��pd�0��n��G�������;X[[$�g:cP�o���ln�(\}ۍ̮�\Cg;�[��k	��]��yI�u���m+��4E��(�)�K�drU�/���RH�n+���;X{�����v�}:�۸���Y[/]�ɀi�é��#{I�����I�i�u��S�.Co��Yw4�7 �5],�2�Yv0�i�<��v�w:��Dmq�v�ol�!�&��]6��U�
a\��H���nV-*|g�e�ыW'h�+��N��"�a�Id���Z�-8�w窻�6�d6����Z�u�#��J=�`ޭ�4枡)���W;���Ա�؛�'&
�@�+U�nK˵'L����:���J����Ak���Ih5��ԕ�7��ch���=݌��!�x6�<����OsU|D�W���29�R&S\�wX
�{KZ�WF��9�ӈC]�5����łr�L]�SJ��p緐e�z�Wf�`��k�X�P��VgS��+l.�X�R��̚��:�9}"�0+,]"��:��C�m'��DY�^����̪�
+v�q$�>������(^%���v��Y����1�� �1�p���U!��6�k�y6�
�\W�!u�b�Cq��6֚wT��ͺE�|kWTR�����N��v�Źmȕ��ޗ��3���j�
�dz;Q�T:�k{�M<!�����h,D[�/��[]uhx^��9��InN�X��R鎲p����gd8t��-GZ�e�f#�#r��g�tr�Lv�V�َ�!p<��wґ���@��ݢ�ɐ�K�S_A�g���, a9[YE��j�NI�)��ż��T�˧�i	�g\ǃ����*�Mn�+��S��4-WTђ��s�gMĕ�y�Ʃa�CZ�<w��p�e��tM.� -41P��2��e�z�+H��ꉩ��s�r\xl�RGt�2=wΰ��M8/�j�	h����=�Y}���*�o
\��-�s���	��;�O�Z�e�w=J�C�#�Хoj⽪�rav�HY|I�{��{B���3& *vm6�������E�-Ŝ
��f��JQ����υ%l��B�a��ibw�T{��5�]c�-����>�;U`�ac�ǣ��N�<-�?�w8u]�6��*�T8�^�8�Ud������Z��g��o.*Vt_E�YH+��G�d1"�B�L����z1u�z�����]V�I c�^�H���L+��5����}��!sM�k���;Y�bѷ[�4����%ʜG4s�ֲ�eC]Z[�3��q��/'�}����37������`3~G�O�������?��_���W����~�?O�~ٜ���c�;�!Sf�B�z�ȱ�<��w�G�9��eS&����[a�ʱ���c0�����Zr��{�r�p�67M��ujJ�xv�|:,&P˻��[�2]N5S�e���e�j@kzՋM�.*�1��x$��r���^Pr�Eh��QYjy2�gXr�n6�Z�{S�9!�i��	�n��Z�����M(6�2���ݫ�w���Q6b��nنh_=ɓ.V2,�#5άxe�����ܛ,�b�,\�z���as�NW*%�+���\�8�J��\���Ŝ��5�I,����\�c�A)v�T!3�R5ct�h�=|�ڕ)�*%���Az) q���#�cnp��\Y�GQ}`�)��B��~��^a�+s�q�yN�+�jYh�%?i�r�0��h����0L/+EMW��Q����NS�78i�F���.�F�Րi���<�
c�F@5M֯tQ�/��N���Vƨ֬h�v��R��uбn�i*GR���j����o�)�I���EE��9*�3a ���V�'��ue�������{qL�p�}$<�m
�z��qn�P�HT�d�mNJ>Kx�\+B�Yg8m�m,�ƫF�%��[<�7F����`���S.�T���n:���X^�1Ew�#i�St��Y�Ԙ�6OM���A���� 	����Єo�����|��=:N��O}�<����y��6�RŤ���5�t�y�aД�a�m��<��{f�J6h+ATRi���i��'KGA����=���zRWO]%	֩4E���]!��/OH���Z6Ǜ'���2y�:ҝ�풞���^���c�zZ:t�WCBhd(�R&��E!ON����U)[w��������t��Б-@P:�F��):�Ka4%&���[AlP�F��E������
6���4�4�G��I�֊R��6��Ѕ�5�Q���mA�
tuA��n0�`�h�S@���-/���(�:z�|���I�F��Eh�^�CK���
+K��n�'GK��i
B���ɦ�I�"m��+AA����������|�r_9bHoTxevbN�n��m3_���<��d�L<�Q$�ȵS���Ԏc�"P�X�k Ϟ�9S +���Û�_w�83����%���^3} N�=<���[;�u�V�'�oTx]�/#N�}���j=�^���i=0ts����G�u�^�G�����Uf�/�]7~�^��ە�/�zWV�v=�\�P7�s�l�a����yez�)VĭxwJ�HL�e���/z��q�ʰ����*˒\�w~��/W�EY��r�*�3�����N�{s}�'oWE���>����׹&�����A����f�<�U��3C�x��y�R^j��� �q�=Fg���A%�'3z(t�%��p�H$��v��;!����ڒH�2{�Jny��4���t������q�?h��}G�����0+��ӑ�&9Z�^��f�Mt�/��=�Bc ^gu��c$�/�D5�f�;w��ڠ�1�%�/�g¾�^~��C3f��N���p�<�4p7��������n[����u��b��;8�
c���x⎓�N<�w[�����<����"ws��s!ӊYϐ�7�"Ҍ�/:��e9��̇��y�..]���T����]�a�o�
8��w�TR�!r�>���x9�'�֬\�]w�n|��4�^�t�r�*-_;o��t���/A�y����8�zF�Z9]�M�3��i�WL��t���{@+�vW�69�t�3������[����sP�/�����c���X6E��+���F� �cٝ�:q�@nސ7��ޯ�O��2�ټ�x|Y�F*��j޾U�<[�T���!k3z��<F�MFf��|�}{g�0�5/G����������"{Wb������W��������%ϗz�y޿���V��?b�������*���w�������a7��y�cknz�w��zP��S�c�fH<�¬w����k�x��S��`�7.ߗc�pL*IE
}��z�(��H���&_����m���9k����?M��_��s ��pc�L�qk$�����2^��{.γ�5u�y{�L<x[���8'h�T[�/�_d����bI�ֹ}�/�����	mn�7�X�Ơ箓ܪ>�Z�
�=�2��07���E���h]�iw:�Ou�ZP�%v4�|��o�и��5���$˂m
ܔG%%�ǗF2�&�v�˴��e�uA�9C��U4ݳI�n<h�ل���sf?;�S�A"�ʰ�͞Y��Y�ޱ��#ե���-s��==)zϞ���y�ں��ܗ��}�s��ր�ϩH����6Z�wq|�<�����sҠ�+ o�� ��G���m.Y_G�|�U��߳.eHe�y8Ϗ$��߽�y��	�{��c��\/��wG����>����/���)�d#r�2E�3�%�{�f��9�>��S�Eq	�������[=34����/Mo�N�����5>���6��XP�ջl�9���<�ԫV��Uפ���ѹ��9{R{|���rǚ���it����r���������f����R����mgi�e�{-��q<+��/(�ўi����U��bt�9T�#��p��.��
�0)3�Q���9����:��/#ޗ[�q�%�����}d�y�I}��â	�T�Fk�o�3�1�G �,!�w/G>�e��O��g$᡺J�A�����vsK^�ـ��O�Wv�N��.��2��ʒkvޗX�ِ�+u�1��ޗ��?�bt�����uK]z���α[���k�ײ|^�e����Q99Zrg�-�6X���j���'���"Nם|{��)�}T�x2������t��롚N׎I���}�;�w���E�T��;�6?{�w���H�W�c����	�N�Y��wh����I��g�K��;=C�K]��/����O7�tA$����=��K��&���9[���'c�;��eP<'���K=�F���a8$���ڼ�md��9:����{�y��Ab�y�Y�U����.����v�i~r����9��^��������ެ)��5C��U�����Wf��	�K\$M���n��QeƿP9{tNv�����sԭ��W����������P���>�7:�s>�w�}��1j�t��� ��Y]����x{�;@H�wS�BF���S�5�	���!��[�^�n1���V�ͬ��[HU��f>��7�5��*�ux�H�+s���w���K�E_b���^�p0r%���kn��ǹ�%s]x�)���NL<n�@���n���.�C�y�������a��];4�������5��q	�=7>5�YӽߐR�t<4g�Cr�/�c���+<�����~�4VOa�k��ޔ����y�ft�^ºa7ɇ�����Q�|6M�Z���C����e	+���j�M���������-t}����]q}����|�#�ݞ��f���^�/�E��5�qX��N�_x�1&��CK��m|s�j�m{<��f���t�b�w���ħ��uau^�������>���{7(������%�k������N�������Z[ݻ�����o��M�A�V�?eN��l�W�p3��#AU������`̚�si��a�۰O'����������^T �9�UU��ת�!��FR��r��<�Y�g�?]��~���N��Y���7�A[���NS{_g�G
wRx�&�e�Z>ۺ�2�����kd��s�
Yp|�A�u��"nT ���$�	塱�|��Bׅ�X���/��s�������,J��ם��"�'@"�m��S��\9^�pT�3�����XW��Ndv�*m��x��R2{�q��#�e�ĺoU��6�bp��߄�Oux�{K�|�}��_��Ӯ�s����ש'/z{�Qp��o}&�Z��t<���6�����Cr���<I�7�vD�,O�_�l4d��g��	�8�I�9~1���ޮY}����{}���=p�Ƽ�	ֆ���qs�6gۧN߰�Y&��������>x�͘E�f<��!��~s��^m��g�:̋�����vn�d��n�՞[���Ҏv���φ}['л�ړhI�g@q�Ǜ/����H9�]�I��ކq�������7a�O1;@��ʂc��!hr�5~ͶF�RP���{Zb��R�,Z��x�i��F��ޯC�G*U୕�j`[Fg{��S�xݟ��Θ�� �8�r��K�wβ]	�cK~�ؽ���+���2�����j�~�I����x�??�ڤߗ�i�Ym�ϑ}���z���
U<�a5�_��`ݮ�<7e�������s����e3s���ϯ�em^�8�:��K���z�|,��YI�-���,�ln���j�pa2��ț�`,�]Z��=;͘r);�6\��{q�5Z����j�^��x�
�J�yK����?af��h�s�yyԣ7�kצ��֪=��;D����>&'!�[h�;��Հ�i���]�'l����zG�p�L�:^ۯ;��@ɱ�Ӝ"�$��d�6�H^�D�x���	ˮ��ۮ�)��w8WݕJ'��J�G�G�$jg�h�>����G)��=	h���6sp�D��deP��e��i�Cf�3=C������,�x<������.9��^�x����6�y���iȺz���|"�7�~sr���9d��h��$���=��<��l������=V7+�_�th<�+�Vc�X�xzZ���>A�k|�y�}Yފ�����^���/~͂}�k��w�����O$��)ܖ�S@����l��}S����=���l�����B�Fε��8��b4]���7���Ba���_����F[Z*�����{ˋ�r�]<�E_���q�M��Ϧl��r}����k��q��R-1�e-኶e*;Hf��G�녍�&����Z׍i�p��ѩpq{[���s��A���KS;�s��qEHvބ�7����э��LU]{�Ww��~yP�O�E�|%Ψr�˥���tz�{^z/c=%��;ƴ����Ԟή��[})���U%uj�N[���L�y��rn1�67v�o���1X��bW^�7�����?�f��Fp���M2Շ���AU%C?O|=N��v~
���V{�|���������?x�o���/�Xϫ�OT9��?�Y�&u�Cy �P��u�uR�Q5�u��<��'�0����ȷ�O�g�j��cϨw�S15g����D���ҧ�~�'�޼�=��[�Z����n�q�D�t%ef�>�]�w3GO{<g�����L}���+���S�C�;���<���'�������"���wY�v}r��J]���uO�� �\��򉧬����5�fo�r�'�\*�TT4=��Η����Ѕ_Ҳz�u7.���4�S��<N�L��K7j�+�jR�i ���w(b&�HdU���l�N_O���Z�ٚ7C\���Ӭ1�++-E�m�2	�#�
�ca*P㵷a��o�9g:��F�� d1)�ևY���-V���/ VD�Ρ=��]��|x�&���<�Z	7 w��ubj#ڨ�x�D�8�z73��	�k>�=B��@���	�wi�D�OΕ�hz�O�E{�˳��tKO�G�;�}��b4�����Wq1tq�X��D�,�K��oCH�R�=r����^��^Q=�Wq�k����W���|���1Q�8;������*.�=���)W�[a�el��=^�;$Ã{d׶��I�캽����f�Mиxh�0� }ɜ��װ�zjL���<�3����N����Am��1��N����P�c��|P���NEN�����3׽C݃ջ�p$^i#�o�|b���l2����յ�P���u�y�Wj�RF��U�A�]�{��Jߪ�/p���v�+X���6�o�����ѡ�����U7��W�b����f���T�Z�g)?D��s���'����1�s����tݘ`Jt?���U���#`��x],g.
±Dz��t7oscf�Q����{!��GA�m*�.$P����v��87Wu�!�rc6��J��RY)�
k���"�T���S�Ke��*�^p>��6�wརX��-}^�&��%��Q�x�v:ۯy�}�9b�^�<�Sے72 \���\��t�r�QO��T?b?-ڏ�e��{ܼ�`2o��~�f�~�z�<�q���9�G��:�: ؍�=��{2������H�9�>��g�.��NW�7/�t���k���v%D�����}����н�X�s�I~s���^k'��m�t�ݬ��vh�G�?j�=ro,��!߾��I�r�_�>���y���B%�Є�s<�)A7�y91ͭZ*�j��I��Z��zn���߼���y.�`�gGLɫ$~�sfWU��T��:`�p��W�I�����uxb��ON�q�|4;�S�.�ŏÄ�89��O�_��xl��e�&�+�#��x������M*f\�B?�TP�T*���'�������~���~_��������s9�oV �7�Z�:>�tF̸�,�קtF5ʦ��Sq�n�� �{��|/"x-�4���l93�"�{lG���l&�u�2�:Kv(;2�m����r��*79e ��8Z|�̝i��r�ak�;�:"��2��:w(K˱S����j����Y&ɜ�7���aCEح��(�;pv��{�^f�lr��.f:�9����hT�GWj�H�[L�s���K������O�!�#�D�T*,4:j�&��{�&#r;�w�g�]�/.6
r��
;- ��#Ϳ>��m�1NJ�ԯ`՜Պ&flء=���Sє�V:�3ҞL��w$�{l]��n�[c(�K�5��Ɯ�g�Y[��:˥��p��E���Л��Z73�q���5Z���vk�.�v�@�괈f�˰�
$�-�[�H��mJ�I���Q�]�c2��'ɲ*�ݭ�2s��O���ׯP�3t��f�o��Ԩ��u�s@h�s�Wy�b�H�Ј?[:)��X�bu�s+oGr٧�t+���b��Z(iL$jJr}N�95�YO3E������]�/��nV�J�$@�G���$�:����E�(�y��P�B�^|�duݝP���L�a�`7:��\Ȕ��{����U���֧��B�P��T�bn����+d���x����W^���WT�@(��ݩ5/f��+@ܚ��X�g�!��vH����ޡ�lIW�孜�y���4ݶ��tlн,��yU�|+��i�xrEP��`�9�wd��+u�?��H&͚�J֖���_~�x��G��g���4�
��z"��s�D�E���(�N�1Qͽ��C�,u���G)t�\�#��[�� zS�aht]�K��h����PE���ԍ�w����J��8e�,7�u��<�j}d���9�<����j����n�o�N�s���Ou8����n�[�\..�N�ml�n�itܬ���+��Q5��e�%`�5���W ��c�<HiP��z��|6�/�Bm�JK�o.���N����ޓ`��դ����%������`�i��OtQȆ�S���ڌ�E˗���+�^����W��VH7LKAS�m�1�n�����Lf����M3M�\<�}�����N�9xn�h�cV#��*�>m���F#�����E��.ݾ!-;�nԽ���q
"��0 ��丳oiL��
:kY���W�wPE��<`��(�R)�%_:�lq537ɩ���Y�Wʫ;Bց\Y�
��7/��X5��<�R"n��
�*��
����/l���5��
qkdd�h��Y� (�(ͺ�OhWY�4�5(��|23�4�kV}vi�98�Z�4e��Q��H��7�j�$E1:������]զ�=�k����@n�&�j�FlL���g^����6B�V�o�1�j�����W5oK�˞>�%N�}P�(�<�*h� ]��x'b�6�}+Ep���
��h��Ҙ�
O;�:�m��p��)���JV�l���I�E-��Ut7mt���ꍶ-j��y�m��F��u��QF���|�]:4�#�4uE<A�A���l�]�y��Cӳ��Q���D;F�/ ��kC���D�i)�OĻ��:#���E[h�����Lh�k�NJ����M�lqZ���ڍ�ŰTmG��%<�Ͱ�)4������k=�7m�G��:�i�v������y��4�'��T�]4yb�-�PSO�i��w���-;�	��Svu�4�]P��ڟ�ǐ|N��tu��1�c�;�u������a��/BQUۍt�U8��#���.�:�.���t�V��y�<��u����O��5ב�-�wq�ݸ�z��OEww%o��+�-���|@ty�Ϙ�|�!�����\AQO.��q����4�ݴ=���8��@V��G^A��8�--yɮ�����<��w��Ƽ��^��8|�`�z�m&��Q[�p���r�&t՛��C�)��[NaÇ�헄Š�#�j��j|�(� ��q���A�κ%��������ƇPW�g�b�{�7�\��E�ΣK�%>,0W�����v"���I��~�#}�O�pNN��������� Z��g�;�ӷXc ��D��N�˧��1p���nn�Rt����q-�Yq\{�ٱ�O�Ws037���%ɆKj��޽���
YsI�_6�{Z"�Dk�U���Z΁��P�N�{�����ר[Ͱ�$?�����K�֧EWu��v�հPfU���wm��]�;�z�8�!ʟ�FM0Yb�� ��M�P,**ʋ,^z����5����'x�ndl�L[�-�l���]�.�w��q�F)�$2������z�N���p�4y�O-�z���x�zފ/] b�����T]�T�>��ʨ�=R��d=CD���E��n�+���NG/[���0�0�=�E��Īk���x�T/k�+kQr���K6bl��>����'X#�HG.�4��Ef�R)��o��K�%#��z�<���Rg���Y�8�oK�&�نq��v�bl����3�<�D5FV�"2�L�u�&����֊T��XM���K���ܔ�׺�k&-__Q4����+%ڠ�R��ٙS�:V�n��rG�w���{(��z&������3�t�ʼ��cZ�,�����un톪�4nZz�Z�1Kظ��9�
aTS��F�+1q5���<C�Źz��F|��}|���|	�G�n_Jm'$����w�̶�~��%弛���|��B؏��L��{�kb��gD�S�t˗OO1�_��i[���������T"��@#�{��{l�fƺk���x
.\�B�.T�m��:z�͟\�1\�0�c8��v�����G��vE�$�gNR�2��I���ЎR:����v�"�U��C��z�0KD��n`%�wHܟDr�yoU�0�
�3$�4�D���Տ�KMme���6�w&9����[v�W)Ƨ60�e��ݗaE:D�i0u5������x���Bp��e?Z%�C~���"	����_�l�<��$����4�+�r�oԘ��y�b}4��g�V?e���rμG~:���g9^L�D�
���Gd�s�U�>*}@��(����9�0ƺ�ߑƃ#��٧���bZ���h���8*T��Qf�#�tE0�N�:�E��W<��a�˿��"�Wj��&ȍl��\`��G�!Q��;*@���.|��˞�E�d�Zr�T�iض1x����y8p%q5��*g�1�~:��V�*+�;��+�SwMoR���@��	j ʖ��\X����z��rgf�Lc���v��gW%��� ��"9����j�Ѷ��'��A�oe��[$��;uѺ��֑R+���E/��$��&���YПi����TA�2c[��}4�[9�L��<��v��zT�8�mrs�<BW1Q*��u�x��ᗒrHvjvΡ&
@�3Q�mֱj�F�g�� ��Q���^����,1�W5gnGK	�	t�2��Meν�}��?���2�2� ��2�w)^@4�aa��z���|��׻�
�qDȼ��{e�}���Ɏ��}�H&��Ai�<@c�l:3#4���sj�{��8��f��1����݇�W��p]~]8�}��P�����ά��L����Zz+�a��ⓟ<+�k�)򃰼��pї�f�s�]��˴��&ӄ�ga�nu�9�b��­���
iBb5��L�.n�������K��W�G�*��j�J845��8jm���D�]Uy��{pt�Q!���_������E2��[��J�k¤�j8S�@m
4N�l���kEf�X$%���ȃޟ�Q�?�_�-7�r�-�Gy�ϵy����+pU�_I��y<8�4�S������	�(���?�3�d��3�!Ƃ�󷝗q+<"F�I5AyFO�y�x��D��fdy��+�}O�JҶU���{$�c� m*&�K?$�|]�
r��w���*��C)��+	��(����'eZ��6/&���:h��^��+�l����zKZ2*�������OZT�r�J�߯��.���s���g�����W�T�:�K>���c�+ҧ��El�m�NB� ���SN�W�P(V�ن�wF�~{s �9>�hjnO!�.���F��L>K�m}�m�R��nI/%�μ�B��;M�C5N�%�m��lO�[2&C��~�"�f�&�Uc�yF��)	 ���Q���>����qW� ,�����T"jRi���]���&���U䲅c�T|���[1Iq�)��U2��xy�<�a�� ���A�Nܬ��n��j͚�#�N����sk�]f��x�G��\=R�-J�ܳCQ�q.���ki�Z�C]��03mtwFOf�m��m9f�1�`E���#Fe�)��������#4���nU8)���,���/a�X<.b�쮜��׽��b��7���4KߌD�L/����o`J����=���ma�!fBݚ�0_��]���P�t���v��1d"pJn����v��q�./Ɣ�����ת9�(V�Мt?����Z���e�lv�^��( _���1�0�u�N������Y巔�5⟸����H�oY
���y/�9��sF�t��u4k\��й��u0�����p�̪ͬ�}��C�^����.^�Vv�wL������p��Ws�L��y.���Fӡ��1Q��f���xB���勛s��or�R|��Z���� �Y46G�z�Ps��P�ن�Ç��P��t<Ɖ���P����޺�����_�pJKZq��'{c��Pr����H}�����U��G�?g�Dv�s�	މ����e^���t�/-���@�7!Ս<E��/�ȧ�m_<��]�6���ӦL7�9����~Aq� M��G_�T%۟�9�
�1U-7y�L\I:�>��6M}�c�L��; � j+�M�;����p2|�j�X����O9Y�^b�
A�^��6:�v��y�Ək��O;�'���,�V;׋�g�8��v��I�R]3qӓ�{b�3�L�_��P��k�^� -��X�p�TG�ۨԕ�M	E"��!�� e���Y�2�R:S#؆%�Ű�.JGZ%�uկO�C^^UH�>@��P�a޸��Z��uw��K�U��W�w�eLV�����%��#�$k#��ע_�S�x��>X�}��_rH�<��L�좮�fТ雔p��fId��m����z�$�󛷗*E�d�k�\�h�I����E[�m�#E\���:�t ɩdK��[2���N
�[K��㰯(���/8!��[��������D����.�wTu;c&׍<�қ�E�$�U޷�nb��+hrD�j�;��^�ܩ@_�+��+�b�QW�4��[˒-�R�3#���6���Ε2��O��<&�4�*��ԍ@�p��<�����"=7�=Xy�3�	��{nv�}��0?�o{�:�_�ۻO�@����uxGD�{����uϋ���چ�r��.�W(��f�̔��z��@]��Zg6�ۛɕ��c��o���
�Qqf%R��TZ~9�����0r�v�}p,NKw4N*�}w�f�>(��]I!�2��o%�m��Cf�%��TZ�����C���{�_�u��C�Om�g�@��#���BO0�\!��F^����n�s��^f�#r��}���<���<��ع�YM�[I,05��۹�@}�,^C�R��)�[�ʃ���1s ���7��f��4�ԺT��\e&��-,����S�k�3�GCK��8��[����K�2�Y�\	��u�q|�H��L6��t��g�u�J�_���_�ut�"��y�|�H��o�{1@��YZy����hu��q8�	�k�>�5U�^&03�w�=�T��fM^v�a�?��$C3���!�9���3��.�P8�wގau+��P.�jh�\�Y¤�8AE�W(���S���,=wʿ@�>��@�>R{0W�����{��zn��΋hW�_~w����dd�+�"�]4���
���݌���9ך0/Z�sd�m`��-�CF=^H���B:"#�N�77JΣ����\��h*�*�Q<b�خ�qC�����G�d�����������.�c��ժh6�f^*�6؏�I��g��� �`��q>TW�9O~o���s�;�M"}ܞ�[G��ٮC�CL�=Uj3��d�9������a�3��4ˢ�R����5��������Ejj�t�u=ռ9�U8�^W$^mT�^�a�$�jvq6آ�0ˢ�q��l3�4?��]a
($wnw]Y�o����U�nb�O��T��tC�W�m-�YZ�H��p�n�O������f\k�us="3�~�h�irb��6��.�l�@ �������՘j�#I�C�Ld��KU�R[W.*܍�`�=�A�\@�5�Ֆ�<�7�������3ӳg���bie����~�^ζ�2fP��'+e��X58�*_��e� ���n�4�\l*m�m�_r�1T�iBT��%ք�L��Q��g,mɛɊ��� � �������80@ø�k�ε�l�H��ޤ�|aF��5�t^�N�-�<��cvZgWu�c��)�k�;��x��,��ǔ�;(��2a�S�7�Q4Y�-CS���sH�ߌ#�+��d����!Y��V񻟋��f��/8��>ІN%�xI�7�k�WY���Azͬki��kSu>b��py�_^*��e����2Q��؋�E��6�����k�l�P&��9�f�ۛ}L�+�u��&�rڜs��|Eu���X��,���]53�ߪ=����0*eki����q����F�K���7quْ�]iE[�C�jp���
��`��G���#[����JF_��|�*d���d��G�8�?V��e�L�=���7e|�� �@6�y_���������?>�q�z!��~�1&�ʜ,�|W���8z!�_�SA���P��ޕ���g�'��u�'���lb9Nd�=|���!�V�����^s9.-�*��-�:i��O��-����{�r|�* ���Eo>��}�!��Ia���g���~��jhnQA�.��Ü*t>r��:����fʱ�S�b1k��K�Sء��0��z�PCmr&�Uc�{�wP�;{;�=�Q�2��@;�v���4�^O�ж���AmbbF�Q�o3����'�'s��.��>U9�ú�u��?�[��6`�P�xp�=�6�M��`��D����*���T����s�C(؊�l����&��SM������Ԗe�θw9�6J�-���Qŋ�j�0��R�j�O��$Y�;e6�|��',:�����#Yݻi�`�uӾ�-��4>w\dV�\�(����x�gl��[BT�t۔��RL��K����Վ��A#''��Iݸ��;A��\C��sQ�hj�D�U��9L�{sSʜ��-�͘�ܽM��q��)�����!\t�8���gТK1	�2�_��X�y�l ��|ثƾ�B��dG^�k���O��r��!��b�C���4XƑ{1������TK_+���'��%���P��9}(�=�]���-��U2�h~g-� ���w�"��Ң�TEk�	�{M�Q�td�rٍ6(N�R[%78(�X?r�N����z9�W�3�A<���P⫓�r_+/"�E�Y�'7���c��l���B}�i������h/����ͩ����Ģ���e�\ֳV��:e�ט^&%��L�B��y��Lh-�;�*?OӼ�|�:&�:c�=���d��ҟo�n^��j4S��O��ު��h�G���cI�0������ћ���EQY�����]'�|��S����/�w���@�^?e��߳��O	��z���2��������fH̭A�Hd�s��Z=閲,��T.1��s��z�E��#�1Dk�T �g�VF�d�R#�%�ƈ5>��dg��9�3��=��Op>c�hq,0��� �5h:b�^��{˭���k��ge�m���`�6� �O��� �M�WT�QA�O���Fm
�3�F U=a_�FSR��[��Q1qȯp�Xs�}��-�V�fnGZ�o7�
�� [��f�=�D�V,�#R�;5�{_ʯ��i�OJ�k=W������ɳ:`� O��\CG?"�l{���;��a��4縋�����4�5	U\ė�
Cb:Y�7u4�t��X��|0ӵ���L���
�^���K��@�ùݳB�fy��2����ŗ�&ޘ�tزHhX�]�A5����Ϝ�Q�)���v������N>�����9�6:=;n��d�ķ1���6�+'S-�%�Q`�ᘚ�w[T٩Z`�a��t釾C]̻�,������C���yN�ɏ�3i��-r
���X�O���(��?\���������mS�.�Y����IO�E�㚨[{�ے��=
�W��a�� ����T;_�)��~��?-�s��Y�
;��*L���1���S'i\D^���J�|�4�\�Ŵ:9]	l�\!��.��z0���l�0E��6<�'�ݺD(jw�N��EW���<�=��������$�VF���=Q>�B)��f.�T�P��so�uh�?YLh�s����St���,�����zL�M�dH�!��c�������������_�����}���������r:�KlC����q��?QnDP��Ne��K�qӦƵa��d��]�a�Gs����@�:�L���+pq��}ɍpA�
��|�mlo�.3P;ti�"rj��zCP3~s��p��A��J=��tyZ�6����^�^�m�����	Nj���aZ�
���Ö�C@��-���ڃ�%uP9��N��a-�)\0�x	h���|�uX��nfX�ء	y�3���w&����V��ۚfV�j�ʊqZ�GVt�Y�v�%$&�y����BR���q�������{G���`�f0�.6xtX�S'v�8�&U�Z&������Ϋ����Y2�E���	N�;;rv�m�Ԋ
�����P��^�s,um��[)dz������4��Mp�`�+	V��D�H��GV,�{��D�t���0%����Phg+�v��$�WX�^�/��X����,��@�{c����qA1Y��OQ=ݵ��E�(��N��Cة���u�L��{�Fk[d.�o;.�j��B��3��6�kKyo:
XOT�׶:���_Y��"ZF�J�mA/�N�0��qV�h��"�,]�f�"�ũ�U׵,774Ю�У�v(Z�C-(zcz��^=E��j����-�,�g]��ti�1(��s��VR}�Rg&�sn���ֹk ���i��ju]�����߰�9X)�ۀ����PGU�Dk�R�LF�$����6���9�`*t�t��[��S$Ȧ��QwO;�X��9�Q8��컙8�
�yku�Th�$�Y�8����M�k�:����[1��[��hM��f�t:Fo�'�/�G��nƻ�]oZblK��$�_v�db�5�J�P�]�>Õ��}a�b�-j/Z����(��cw����.e�ە�;�µ��)w^��{�O��A�;E��U�6Z�k��[�Tw32�yGD��Z��&�W	�����N�7�K���ӷ�v:Սo�xڏ^�ǹ0�3P1M����[b�
��X�nbs��j�z�>݉�^��6tS����I�N�K�-Cդ�]4�iu;�V!�%-|$��5uXD����D~���]u��n�eJv-u�=}xd�>F�(%v`�EJ���˥��,pU���٘�����
j
Su:6Ϊ��W��ƾ�-l���fAʑ!�2/̇�
Y�Q�1��K�'��Չz�4f����m���룏{�م\8��Izoa85��ƹق�1JWT4�r��yS��ӓ��w4\�4/�q�(ǡ>���i�P<Ea�V=�)�qޘeݵ�ڍ�'-A�	{7��ww�~f���+W��	��7C&)��cSP\)�:�L�����c���C�4ĭ�h5��������qK+��U�zc���bӒ�����i��M i�dw��,I�����8/�ˊ�H[�c0�-�jJQ��ٜ%��@ɳ�r�i#rn���l��]tD�t�4z1|Fa�}/�A��'�&k}P�����ЗNK�.�2'�t�r�{����{��	�s)��Ֆ�$��� �1�Ae�RBv��u��?_S���@��Tzwc�I���DS�כ��]��#�<�@y��Mh4u�ձ����u]�::qV���<��N��GJt= t��dհѡ�@[֚ѣZ,mkB�y'p`Ҕh�F����u�"�hղ��X��O$��t�F�y&�7�@v�B�l:)�I]!ݩ���k�4�%��/A�Mi���;:J��1 �))�4�f�B�����7p�@�ДŦ��ѻ���i� :�N�Z"b�$�;��I�C��rkAQD�j��d+Il�â#ۼ�GZ�h(�آ���:�3���߃�w��/����eu}��WC1K��mH�ru� Ȕ=��#$�\j�hL�|�ɼ���8�z�ߺs�t��\�Dvl[ ��;�/�C����u�#GvZ������-<�g��U&x����Y����43��_�uuَ�|����0�=&��0��XR(_��Zyk2�>�Km��K�2�����j��h����D�Ȋ��U��ek�`d�D0���܂�D��[s���������Sh�s�e�ɧ�gq,ja����Xʄ.a�E��+�����K}I�������P�&*�KW��l�:��&�}0� s.�L�,'��&|� ��жc�@�:`��A굃�8�Y�;�:�����\�Ƞ�s���/R����n� �P�a�L�r� ǗE��brȞv��S�FW5T�j;�Y�d�3e�MS�W���L	�tÜ�%Иm{��V'�J����j��܉��Yؐ�r��q�/T����2�B��\�K��^�t �(z]�e���
~Sl%�n�c�r̫[KU����`"��].B�����a�}Ly��㨜l�#cK�C4���0��IȽf�Z�ˮ|U<dN�Ħ�^>�٤�Ŷ+>�dzmP�?p��}��,�6�k��&�{���<j�jm�^Xu���o�N�&`|q�w&EĬ3��xoU���C�a9a�u��aSC�._[��z���w��i����V�`t�3��n��ֺ3y=���쫊�Kz멦r���Z�1Ҭ��W5�}y�v�%�Sq��Q��{��r�9�}�x6�}8�{���MVg���UE��8KH�N�����ƞW�-�����O�����O~�7��S�0���,����l��危&o&9�T�Mr��Uc�}]��T�@�N�u�O%�݉�<��L-+�b�<���(�p��ue���rE��s����pF�xT�����ܑ�P��`	���Ǝ|�f��x`�mW0H�e��a#53��!�&9d����ͩ���&��Bb9�Tɔ��=�}���*���ٿt��A/�����4%�M<삷���dD����
3�!�(b���`9���s9ȁ%����j:e��$ّI��r��*;����>F���t�Sk"��-D�LG� u�B�j���)�u2rwec�_g<��4�>�ˣ�QjZ�(���p�L�	c��GO���:���9�l�(0��dm.��5[�ϲ�Sp&s���@��,��[p��%R���*[^���͌p3���Q�/�Gjދr\@py��>��fE�è�:�:9��uCSG(��;�(�30 �a�N#ǡ�e�Ӿ����|���UtS[p���e��C�c�8��|0ax�Y���VII*�c�c�����m���R����Pmu�h�2�;8�zi��캶�ntd�`��%(��E#:�5M9v�lL��/k����/AY�,���U�W�t���n�\��u��%�[�X;a02j,�O�.q����[^�2�ba7W��-w2ʉ�͈y��P^��U%��RE.D^s�x�Ǽ%�c>B����n_�^)������7K�F�W��eW���:���}=7%8%m
8�6b�[4N�ٿ�	�_��o�ή�����(��;���nN8����V���+�j�Z�w0�l��I�0L��w���F5�@�{���V":s��m��dgj�F��wAU2S#G�v'�{�w6S�����~��U�m����{�F}��^�20S�3��c��p���.�0�YN.�t���NA��6�/s��Or"�2���@d�9x;�+\�.1��ͻ ���<�E�RS��(�5�Tsn�\�n��SVe��Jdg�q�)06��Q,Y��Giv���PG����Y�J�Nm��֓�1�9c�^~�]�X��>�Vx��.I0u���ꏈ`Gt3k�2=�����횘��^�,��||حV:�	��$�5c�(~i����'zƂ�3ҿC���._w���?
����&�عm�<�sUb����2�� ް��DՒ�z��.'�g�
f����N!�g����5�]��q�߉����+Jm�;���9�N�ݠ��rU��n��Щv��c]���v8vVXy�-\s�+�Ĝ���x{������%��9^8�pR-��UU���W7f�,�K+� 3�H�|r�4ʻ��ѽͻ؁�����k�삠�)�<a�a��ϵ�)k�n�m��3|��}�E`u���潑�}&e�S���"q@sA�����i�{F���|\���&w����3E�r��ҥ�K�aM�o����d}�ѿRd�??_���/�;Ď{۴c��H��x��nɧzЬ�mN�B���Z����x�["僔KL	3�|�/|�S��o�U�4�E[d�t-d�}h��C�[�'� j�;`˪J#�ͯ$⠘���(���|�S���3�'����-b�5nH�|RӫS^�����9�"M��!�c�w�2Mq"��1�Kv�Rƃ�F��n�Y�Kd8�t.jF�t��W��!*�\�df�ȱ+�qtY�FpR���ǉ�n��QX��p
�4�H�j��a�Y��Y�הV�Z�_�)�ENc����T���ڝC��%���H�^`��2M
����[������\[���0����Վ4� �0d��Y�k����.ݑ�p7s/�Wj�5
��᪄V�ѧ�V�u3Ѯ�c�y��� ��������ъ���:��c�KY�M�O^I���2.�n��폞=A��!\�x'>���Ņ-̠�6]H:�V��F��d�%�A9��Kf�d`g�{�M�� �7��E*s�z��� *St�2�^��e������{�G���97p�B΋U�b�^7����r��:]�7:���"�� 땋ht*�އ��/��1��K��K��"���f���B�1cn�;��8D/+�P�	�E� �=���F�$r��09�`�#L}�y�ܢ����쾷X��"��{�R'�{tж���Y�M	���s���3�7>ǲH��0S$C!
(�N���*���!�#�k�gL{g�%Ja��Y˥�>��L�=�b��*K%��M�[Y���s!���\s8/�[ ��+��wz`���	b)l���%J���*9N����n�&��^����i4;�9��6����s��7|�Dy�3�:s�osT2Ͱӻ���l\��c\�t�--��x�^���.υاbϏZf��Z���]o���_qT�r%��~��_����ɖ΀;��Y�B��s�(�i���y��"$J�a��][�#�oMeX�T�pq��ʹk��%�O�����3��ItQ*Z�<
xf�$���Z6�J��n�_p�f1�aouS�6#w�2_�
��9��i����Mb_*T���w��|�`�&����xw�N�sm�/W{h8���v4�u��C��x�F�i�1�vM�T�lL���j�~�ٍ�ފ��c���!M��ڎD_�MNkץ�[]8�/T�����N�f�gm�,���q0-og2QP�bw"��cF�.]�C:���I�7�nb�Nj����2�!dQ}���liF8O�-|.�PD�lHomI���~Yva�*lS�0Q>���#��\>��}X��t��ŧ*h�I����j.��6�-�{�sV�ʆy ;j��oi��l��Aċ}�v�ث�:/�Mq7�ާ��t�k�Y(��~ħˎ*o�Y�Clr��60��mopАsf0X��a�޵���9r,/4�\�0�.5��V��X{ J}��卹3q�K-��#[*B�� ������5N�(�B\�E�S���/�&MJb�T�G��m%+\P���H2�'I��^�Ҭ�q[��x�l���p[�ϭ��4	Æ���6��_�2Y1<���v����1Z��s�� �H�ؖ��|0�D�?'7[>�ƅQ*�����=uZ*���<�)��'�S�h]��>��Ur �bm�^`t0�>���EA���vx{�Z����<%�K�>.:�6k�?CJn%�;��崦��X���ƴp�R���Z*g@��=��`q	��P	�-��Z�f���Vk��o���T��vi�cF�]F8�4��T��3VN�t�t�5v3��nzf֐�M�չyo�:�s��c+)�Mv�����}�W�_� ��� ������4'⅊��C?Gs��(�e�@�}�@�!��x�.�d<��M�"�_&5q���rQ�v3����E���H����a@�-O^�\�
��O^��s�'U/��(�f��Co=R�+3TQ^�8���cAEf�	����m��g9��y*�'Ǧ*[���[Y���1��s��Y^�'`pL�|�~���W�֫5��7rw���3�q8���ޝ2��\��EU�kT�vxV����fw��g�i;o�b�E�|n�ݪhj�z���� �\�O�s
�=5%�o}6KlڒD��ϊg,���?bdq��T�v�j�mm�'4�����gg	й�# ���-+���!�|���ئ%��g�6�8�g�
[ew�q�317���.8E�h�}�9@G��D��jp{'�]�U5��sl��|M�E���7!�*��O��s���U.�CFay����p��\�TSg[��z���9�)�9�$�%�Q4+2%2��u���	�=k��;Vy��,{"S�
�C6Қ,�;��6o��z����ȩ��zQ*���vYZ����*�W^�h�S���nY/vV�BVQǕ���C��f�����J�Ÿ�uxQ?{k��1��ڰ��R�8/3�jt�%(m��klC�n�X+KA�
&��1��۫|��[Y����������o ��  �k']댋�!f�Vk�Έ�|�h�Ŏ�(5f�)-]*9N��B�T/ mX�%��^�5"g��Ap�>��pg�KM	ɭ]8}/��g�w��|j���p�O7�g2it�l����@����.ۦё�ٻ��G�g���^h/��(f��櫓�:�Y<Mј���_�PK�8�J:��7-��-#�v�����1��݆0�>�8
t���(U�+�[Ͳ�2A��?V��Y�;Ѩ�~��|D�-���������`.sd��sY)X��/O@�B#�,3��M~��i���?=!��MzI�grч���D'3[y*�j�8�"H����ʴ�-υ���r������3����r#ř��9�&1H�U�2w�+G�:������8j��� _C_e3���71u:��y��ݑ���,�i�{��+�3T�T�T3�t�1&r��󆀤��
Q�n�O�����6�;x�@��R�kΞ�����M;Ex�!��)f��J̱��(�i�mN�4��5�i5{W~t*-$�2?e7�䯄b�cs��uXߗ��*���N���n�ti?�F=��@ۏ/!�_���JX��'�>$�H�*k=�IM��Ȅ����Zy���ٕ���p���VS2�����m���zq���d<�}�7�}q��<��8Q�;�>;�U��L�(5�n��
m��:f�c�2x䣀�,�ċ�b�!�c�w��*�⑋�Z�4�rvrnp�/���EȦ�q�m��a�V�,;��L�o�W�,�\�pUyla.mv�V,�vҞ��Tj�	��'�C	�s�H��v��ke��QŢM��yEiZa��ؔ55�B�3�yݳ(�]3�]L	���3x�mO��8�4��yy�->�������T��lBe��2�m���Y�7��T�k�銓~�v���S3���#�t��Ml!�s:�/�p�*>5�B)�ru�_w�R��r7@�t!�8��4F84%�sԹ�\(vF�C
1�ѹ�d�.k_"�n�0Dz�����wmi�G��r�[p���`�����}u�3rp�����Լ�0 �	�4-��&�T ���Zc���$ܶ=�F8����}`��ڹ��U�S�3��=";}F|�cOq�3�ze��R��t�0l�.���*��{�I�f��~�hB���b(�3���	�0#�}���̧�Ƈ1i�p	Yaa����AJS���5ڣDL.��̛V�p5;q���TLW*�y�
x��5�O5���G�y1F�4�^�qNp5@a)����Jswa�E/{p����/��*�k]�vR!k/z����l>�鯯Z�|H�0�V���:���{P�x&������ȳDbc?s�s����z��C��1��$O��,��k_G�5[p��܉��5�Q��*���T�c�;�3�C��.+������K}I����0=wɃ������a曘�m(���O�vԁ�i=�0��P��GC����0���v3�-��g.�35��^Py�񬽃��葙 m��9:fגDi*���#6��mQ$l�Ι�a�=Nݤ�:��=䋯I��B^��5]�&�\TAz���|���P�*[Y&�FYu�)��zE�p�n��
�p�\ѹ�ن(i&��U���,P��iL�
��S�N����k�q��̾�蛦���+T�	׳�e���-�Q�x&Q��}�����/�����ca��nJV:^]P�)b�Go2n|�����p�f���r@���Z�?��Z֝�.�W��}y\��&"�M��c��(��T�q�B����6�,���c�B�[`��b���垩�u��ri��0w�|�h�j�QvwI�g��~)O�U�����7{1b���G���<��?O���?O�������L����m����w��T���������p�˹+���|��X��[�nV��;.�<A�7�-���:�������Ei͛f��J!�Ts�f75N��kan	�{f�7(nLNc[�ldh�	��p��¸n�I>t7Ʈ���Cq�o{��`TS�s�}P�;�ۮ�+s�ۀ�����j�H�엝��vڛy�ɕ7�v��ew�l�1���҂���rdϬ��;���0���3gkCE.���n�W��纼���2X� �dخ�7�T�؃{�ZGvK[�n���M=ZV�J6�Z6K��A#���Θ�v@�nbdS�U"�w׏��SփĮL,D�t�(%�TW-wA�X�N��4��������m�c������_aL��î+�ѵs�U�n�-;���P���7vT�޸�Sc��41�p��h<٩b�h��Gq�u��.�YJoA,oS�t;���C���l</`�J1�ӆ�3��U��*�kOi��ƌ����Mc�	[�|�4ض�^t纎�,iѩAcz�8��|�t�߸���lf͌�F�˘�n���fb��M��j��r�nm��ڵ�%6�����-�V��=j��_L+�)�-���Y�u���7��*�mXA�ݣF֋�Jie��
�sB�u�]��ޓ�l�ҁ����w��:띐C�a�S��;�#�|�t�,Z2T�9N�P.[�!,ק�[ݮB=&�p�DyRy���c�Y�Z*ݦ���;meh�&{\�����T=�8�r��v����.�V.M��1�/�Il���17Yy�S�|ֻ���\S%L�ze(:gbx�!$�n����t�u��\*v��f�/Ӽ�X��jO�a=ã����wb����Z���0�ھÔ�f�ǁ����5�Ôrr7)���k7IbF��9��U��Boƈ@�N4݆.�Z���b��lW���e�O��ie&��\on��܋f�A�V���W�.��\[�b[��70 �����Z����s����.]9L��f]��IݕXVޜ6�.
����٭�0���
�eP;m���j-��=���:�\�����sNeiؓ:�;Ydѫ�=Ɔ�G{�thT��έ�néܺ� ֘�"����$�b�ɁS�Z�/��ܓ:V��4� �$�ċ���R�4]�l.^8s�i|6��Lڶ���]�3.�6��n����>�*v��<&��4����9è	k��N�;�r����h��{5�QH�DR�S;�����4ŚtD[}6ީ�Hq W�56&�
����m�ǯ�Z�a�s�n���b�A+���粕 ���qWx��&��4����+"u�X�q6�e�N����5�oE��N��sR��YC���K�4�(�����C�Ӧ!�Ϊ�4nƘ��h"��Pv�Z2SC��F� ��렣��AM%/c%PPQU@[��h�cF��QUt��ڊZ�N��OA��M!F�L�[�@UD�E����&�lSj6�E=V�6u%%�qARu�EPE5��PG�I���[VX��+N��S���v��R��";�,cIZ��I��I���K�=:�RjL�A�ASbL��٢�i�Ov.K-���@b�GwqTRl`��U$T�D͌��ĄAA�IM�Z�f5��vJ�4đ���C$���~1�N�{�\�TL���}�[e�컣6���HV��KW�N���gc:q�A���B�[[�8a{2؝�<���������U�(��"PJ
R�R#�{�q����u�������K�s�0��x����^�R���)<��_E�#�*�ӿ_��t��b"%3y�	Ls��[�u ��yǑ�ɨX;��iO0����nْ��1(�M�kԚ�'
�9�, �g�2X�:!�"sb���l]��K��Oڛ_���ǬeDb0{��j�}\��m!�l0!���C,�>iw6�g��'���#��������w[��6d3��R����C(��W�⮄������ȃށl	&8��	YŚ�}2js�Q5�Y�+*ε��r�SM�'�sP0f���3��c�iZ�z�x�^��~�	�$N�U��2Τ��u��	�F�hX_�B8)����.$6��ى���`c2U)��H%_�+Cf���YP����n���3������>k�o�Jݙ��fd��%۞���8�$E�q���T��N�����6(�l㓇q��dx[���1�b�����a�+�̓ن����/u�	�(F��q�-��]�ua��뺱 ��t���G=C�`C���^��֕4��¾����}��U�*}Vr�beiY���b��0q�Ğ,�Cp�R�9X��]��,��� *%-������G��	�I����+�z��~��Y��ˮZ���<����r����͝%hز|zhL�v�������X�(�پ�͡��tA����+����������f���'��)�\�ߜ�Ih�V�-��&޽�ERܧ����
(��[d�����<�[��R�Hs�����e�U�i���0�0}�AeZ��d�骭\��i��nV� �ۇZ��u-��Q�����p����(d��d*��,(oL�[�U2�:��9fV0��� M�hg���;nrq�i��w�=���(z`<��Cn��g�/~��S	�y*�զ�a��1��Z0��/B�[Kw�԰w�g��ϭ��~O�&h��<��H�c*JR�!�#���uG���h+������)���@J�a�C�t�2"!>�OCk�{"X�ڮ�g�Lsjqk�\#:P�T��u��u#��j�nj/������-���wC5��9�X���g)���m�tF&�_��P���Rv�^J m����-4���͆.�����Mgq;<#F��[���F;>������\��5�_��O#���6�ǈ��&�Z�H�v40nb%w2���\�$x�aM�1��0�3�#M�6e��l��I�ۄ׺��z���׀\�t)2����H[���M�A�IO��d�(����B	Au���V/�����@e�ǵQ��-��k8��j>Wo�8��P�[�k����{%^�S�n/﭅���{7�m5�:U�y��6�:8��b#;2P��[/��FPэ-5ؓ��7���^�\b��}����|�>�<�w�(��!B�B�������o 7�*��Yb��w��LE�$dPks������Ϛȳٚ��05����s�\1�=r�6�V��w�C�Zk��`� ���N/tO�KT�¢���l�k�DX �l̉�h��a��:�q��b�v���T��N���F[L���ၝ.F�^�^D�D���2���F��X\�$O�� ��0�f� 7�B!��]RQ��$�.Ӯ��j�r�'��������5UxU8
j<or&��oMzӲ|��K6��j�6,��Y���4_��R6�q�gK���uz;��|�P}(�dF=��c��M.}d1
�[� G&[4%��t$2�̹7e�6WUm���s
�p�ӰV�@�P�.�$����Qy��ۉ�7���4��=f�S[�%�"�&,���)7l]�Ѷ������&E�(#%�������P��֬7<M�6#��<��Qi���c:�M�֟re��e�<c	SO�A�O���֙�3pnC�Qtۚ0��.X[�!lS�r{
"����^����1ށq��t��o�k$�`��M�[�p'�ٓ;.�ܺ�����]��Y݄{5��Lݘ��~�&*����R� �!�$uk�@]�F:��gC�u�r�����P��V�<]�r
Q��GFҨ�[�Mme;7�l7A,O����>��{��ߟ��?�(ҪP�P(��R�AH�@�_�ǿ���ȊE��"�D6�0DV�K�n��_�vq����v�vSud�i&��!>��W]���n����#�	R����	�NL��|�R)�v2�,ܦ����Qe�/��$�ft�wє_rԄs��ѻUM+�"I�	�à��Ǒc�q�3��3���%Ra���Ӑ�������t<���IIxu��\X>��#�@5�A�:6��C�q��S�_x�^T<��3�����2]�y�%��!��3fW=�:8,�-��D1�Q�Z
��o�I>Dx@�=Sֳ4���c�xa`�6�>��s��I^Cʃz�(������;@���*��2�DS�V���\*��UvA1{2<���5��w@��Bj񈶄��yw�A�O{�i��CTV3&xo�w���� q��+���U�m��YQ�,�jg�#�ItV��<w?n�UYT���{Vz���(y��rE���:�
����#3�!+GU������?o��VЗ���Kn��^�ܿL8�o� ~�� mk#2~���T�3��Jgh�C�hX�a��t�9��6�àu����X7�2��3k}H�%�� �5/nʕJ���c�?�z/>9��/� �Q���.�X�:l;��U7\z�%҅�W5�';fw�M��V��YܰIo4��6�m��ڃ[yG���n��c�0�;+6�'�LX'8�ib�䝘N��mJ2�_k������
()"Ai�F�Fo{����ڐ�vL1�X{�5u���D2��ڃi�_A�9
����}	�PS�ݩ��~oTǱ�s��F@�,�0h���l��@��<�ؤ�cнJsVb�p��!kΐ�2 [�My��&&�CA�dՅ\�"vb���Ĕ���B�k&Q~���q�����ߕfP�G)��s�l����6M7)�ֻ6.`F�h$2��i`3E�*Upæui�s�Q��g,m�3y0���F�
؃�љ��C�L]�Cy�	�a�g�a���|i0�MJb�T�G��i5����۟��HӜ����g������t��u	x-�&n/@c�<�jz~�'\W�ڮa1z�`�ri��Ɍ.!�?+j��>"~�3Ei��QM!���秪7��	K�P`T{��С��`v���u��+��ţ.)��=�����Ш|^_��!��\A,/�z�=�z��s����K�ۙV�T����)m�O�B��)�C���x�7�����w��E����*`�Xq�XUM�N�騑�P��n�	���cހ�\ϯF�$���h#�����j�#Y��z�[ű���}��\5Ո,4{��px��g�����
isU��8���H��r�����I}��R�I�:��()���{���q�9M
Lܷ��bQ�ʵ'4%z�eq�N�*��� h����>���JQ
iPia�y�������Ψ��B�9�軡�Ŝ��؅��E璚C�����u�m�k<�J�)��c�K�0���e�%cͦw%��P���l2"D����yE:�CX���%�\����Pg�i����In���[E�z��5��(��=�ǃ�h��?a����h�/�A�P����ұ��*���߿{���+���fCj"V{Uc�tj]�C�Wf�h���y
�������ͻ�%�e~n"�>ͧ�+����=��<����?^W�%��i�X�CL��.kL����>�xp{����8��Ӗ׏
�wS'l�/�ٱ�b�Tyc�7I�z�UKJkW.�=F��v�5Pzvz��-�kr'�WM�q�-��l70X`��ʧ[ ��\�=�0�m�������t]���˚�,놕�P�⽰�'A"���a��m�J�\���UJm擡�Ls�ʓO	�p�Wtn.|�?y-@����GMN�Ռ|X�/!�����;��]�,��;x���@j{U�'y�:�J�ђ̔,:+Н���:�;,��˄pN��h�8��9��&**W�A�CakM����o�r�{_+{���=�'����k0f�|�9�&�r���f>W�I<�+�"A�<��.S����24�$�����U��E�c�ZWOc'�Z��yGӫ%^܄����!مJD��j�����o�ܕ���k����ĩ��=̡�dg�������ZJZ@�F�F���)V�~������������x4U'oY�#�x�\��A.��������'�� }�y��R���9�&���|=zWh��g�B�N̎�� gZS}I�
yd�F�{e�-4����`5SI�1L��Ӫ�̪Ϸ��O�^�B��ؑ{�1��ϕψ� ��j��c(j���a-G^^�����|آ�́@|�ʄG�yW�U�M� :���{޿�����v�%X��z�F��/��.	��5�'ß���`U�S�c�9���u�F���p���zZ2�SM��׸�:K��T"ƶ�u~L�/hO�x�_��{�FO`VGN�f���ۢ�aqײF/�2y�����E�肎�&�x� ֗�"^��Z��*�Y$��(\�XKU����!�~akT �1K��4���-�I�%�0�	�%H��&�d�=u�lųMA==���/�S�x��>~�5��p�ǹF���q"�I��o,@kB;��LOk�>�O���H���]�A�n�c�R�A�'܄��_�]0Cl��x�L��ao;O@��S�E���t��������:+��ӛ�N�,�mVwf�Y��A�3�9}�уQ�`Y��;V�؉IR�E^����3�8�C�~��8��ӮX��(��ᖢ[u��T�ql��;��9؀���'ό:v�QC+/QB�*�v�uwo���~>�>�4?9T
DhE�ZP7����;�u&z�Ui��*��X7s�"o�T5�;�*Y;*�F���Y�f�����vY;Iᴞ���n��iZ��z����Opv�̕>w�f�y%����`7�B���P������;�v��*��d��K��Mr������,�f�=���u>�1�����Fn�a�z�R�n"��7T9�5^�T��ȨN�_q)�|�m�������/��F���ݚ�y0n�.ì�H��A�	���Ō_D�o(���.s��O����iMKn3t�LJ�(N0vd��QOZH���S+�}��]A9N�����?5^�MD7�2Ynx9�gizG�Ĳ�gm�<�a9�	#���9�������`ƕƚL�6��V�f0���(�\���E�����0Թܚ���U�:�y, ~�*�1���C���Ն���4�c����H�
F;����6w �j�ů.T1�Z��Uk�&03������f�$ڎ��Y�AՎ��܇���/ݲLL:�Z��cK�nGpcN��2Xe3E�{�lK�����D�ǂ�4	oz�Y񜵒�.q�on`�UG	m���޼NV1<v�ts)�k��r����U�f<�ϟ��ˌ7����[%d˙��MD+�AxQ�w��{[Ji�m�-�d���6�R�2�m�lq�� �`��"�M%ݔ��?N��~Ђ�-H+;g9�+j��ʉe���gM���_�_|*)�A��������o�߯�}~9E?���dߝ�=^�1��Y�]�&@�ʡ	�;�toCr���4����+{�AM|Q��x�����n��6/"��v8��(,��!� ���L��!T
��L�;+���j=p�����ӟ�Z�!J���a�R��g�A����=%6�)�J�M-W�o��T!��bJ~ޖ�3���}M���[^��1P�'�|�Bӷ�gY}hR3�Y�r+��oӼiX��1E��KhV�-\;��r�{_��6�&c��=��ru�e	�rc���֘�5Z��!<p�^�t����[M{l�,�ڟT�k�ː�X=;{:�X��3����Ys3W�M��z�^X�	���R�6�u&�<�ȭ�4����ߑ��|mw��s�4��9i�f�Ȇ�	e˗��e� ���d3H�R�߁���`�l���G�WU�0��P>�R������_t��G�ђ�b��3�m�:-��1[��=b��}���LS�T�:��u�V�_��de-Y1��H�i�,���Hq�&Ƹ(nò�}f7|�n�4�vOAo��u���è��y&���(�����1�<9@��������;/�;��B;�v�����K�
���/]� ������tM�[�ۖ�j�h88�n�Nҳ3/eÚ�h�#V�=T0S�5��(��4x(��9N	�v�nZ��Օ�%���wC��e_� �xea�zS3�,��T���|��(jg֡�C(���w�}8�F�q�$~�zk��a�j�Ub�����lB��Q����ו��k�%=i����6�3��������nA}�;���J�ͼ�ȦՏj���4�oP�qX�*K�P�N'�2�L��
gǠx��z�8��]Z�C"�,�]��0�A���
騑��њ��P�z+�?�7����]n��!~�;(]D�����b�0%3�%��g�Qh��E1���0ck�_1���z����a3w�[V)�!<�nsI��x��0	�.���va��-
2�KD�r�:��8i"GU6�x�\ю��}?zՕy�uo<��z�`��p��A�ޖWʽ��
�x߃C�I�����8'�5�U������z��j�B��9̶��;]��K;�bAO�t��9�N��|�=%�2�%%�\�����	�:5m��M�ca"D�r9�%�+�զ
���&��Ia���eUc-��6|�ҶI�ý�2�e[��[Ǹ^����(��l�{g[�!+6.���Dz<�g�����z�^�_���=�^o7��]�˚�Q�X����T�ptΫ(Dk�Hl�*�UY7�+U��z��##��H�����u�aMp�;�/Xz^�h�n�r��M�iO^��^��j��v:F:�z��N�*U����Rs�um!y9R,b7ՠ�/{v}pލ��%n8u(CyOS[��	Bj��y��]�U�ݩ�c��oB�7:;���N�"V�B�X���I��ᗊ�Ncp�PV2����	ض�}��
��}�i�ڙw\�Lo쥴o7nP���n^���z8�[f܇WT˙ڲ��:���6wcUg8�5�� -��y+q2�3K��G'�I6D��K�J��_�nR	���IX�̴�� �&	K�8�r��QZ�m���R�����-X����q�N�#��l!pEt~��Π�.C����;`��� �����xu\�������H͙X�2�3�p�f=��N��:S]2M�lg46��b��ڹ ܶ[�2���i�@���X�����H���T8�'d�Q��q�hXݸȔ���j���)}�,�F#���|��@Ba�Y#Qˮ[i�gpm��33�9|�X7�A'+/6sK���̷�bT�m�,wy����˽R��9�&u�PG�dgD�{�kj��S5N�W#=�=���R��5�v�r���@�[Dܢ�m�)cR��<��Ja�������V%n2�P0��-4�2�E��.@�	E^5S���u[B֩�}ջVF��Y��+Eq�ۚ��[z@��Ϸ]��mM��]�8NT����J��c���Ek`�ut��z9�6���9D<0]\[���O���EQ����JYJ-\���rs{\�]w�t��C��Y��X�ѷf�\eLK�7EB�(��n���=����Z��y����˫��z�H���̂vt#aL����vn�s��y+]����m2v�l��7YDV�kW:���t���@�<L�hbw1W0��z�B�K��M�ȫ��z�ݻWn껣r�Ym����	�$NsZ*�6��E�� ��0M����oiz�)��_����0ۙL4^c�,_�Z�k*��հyɺ����g��B��n�@qa%��6��U���eLr_�.�cS��/i]�\y���@��E�M]�DT�2��D�:��f
�Y�ONe>��8��P���#Z�=YX��g��ݧB9|H�i���rۊ�O~k4�oPpؕ������_uV�����F�G-�}�� )�v+����ȶ=�v��^�IѤ�Vt���U�G�c��w�*j�3�d,H\����r/�+��I���Uf\R�m���'O6-�6�@��.-5rM�u��m���C�ք�ۜ�h%�Գm���U��\#���Rw�u��-o���;hVs�p�PI�M��Gr�>�%��Ä�S���eJ9�m�!-�D�8-�FPJ�c㷗y��ȫ����quvZN�h�b��A��MQNՊ(i�Altl�ִ�j6J(�A�m&c[�F���l�b4FɈ�V�ڞ�h��9+�ښ�l�"
i�m���cC[[Z�+��SV���2D;cl�Vڄ�� Ѣ"��&"�A��"�������]wm�S0h�.ɪb*��pDT5��Q��j��FڝԽ�F&���"��6��vsѪ*j��ڍA0b���b�h����{j���u���u�)*�э�F�4h��5�V�0MӪ
��X���b����Z�TK0b?!�������:��R>�Z���G�[ݑcr�?�s�]�����
y5wJRWe]d�,�e��D	��ٔj��y�;�.�0�}o�>_8���/;���'�(
�-��0o32����dɭ?/�a��B��=������7�x,'ze2Y⪙s���p��eV>�1�UgAhz�y�L��6(^5���eť�]����c��X9�����jb]�V;ҍ��6K{���Wj� ������<������K����b��Y��,���b�5�v���ح�����F�\4��(���c�|v���W�T �K���S��m��wE����=��z_v0"%7bK�c.�a)���Q��p'N(�����"��p�p@�|Ρꯙ�W���he;��(��&�L���Qkc��HzN�S�$�5c�<7֚`���`1�d��o�hB�͝�#
n`���f����<%���s6�[n��v�p7>W>"a��p9�J7/��I6M>h�̸zt�)��6!�xYॎ�RY���n�	������g�������|����vg��d�11��1>�^�P�b0�����`@O����g9P��T\�-�K��L����5�/>�s�="ƙ�'��|��E��9ɏ参=<(�����q�Ǻ�v���i��f��V�����w{�W�����N�S���4й�O��>����nⲆ��ḑ�AFh�����҉�r,��ޤ��i����әi�'�u��]=줅��r�V�l����ر�97��},�w��9�}������ ����x�|�It��3n��X�'�w1�[hw� �|��T����~��L�7���ߔ%4;˸��?&��g���f��O��^eT��T��ʐn���U4�#t�랝�!��1&\-�l�ev�{�4�p)�6�MG�W���l.��|e����s�Y�^���E�˕�t^gh*Uc�p��xL�]�q�o�C�Y���U��
7Q���/.�>MY�V�`������i&��������ה�&M�����c	qA�k�K����$mDwk�2h��GD�yÔ5q�&��޹SEM���cN&kP�/�E١��Ǫ܅Rŷ�I�-���^F���vg���fa�� o�2+zS���+^ʋNN{U�YX�Z�79.u�t����x`xL��3=3�׍�|zr�_�PY��;o<��TX�h�jJ��C��W"��g�-���ɬ[�c��wYhM���!@��W�$K^��MB.���7#tkm$v��,�)���g{+Tl;�6�<S�� ������/%��H�y�R)��ɗ�P��H������mi������Bu�=�H��r�C+q���G������<$��{���<�^x_����ji ���b��g���[�G:�8��Ι�@�ss�eL��P�Q�l}��h��| �۹�.̱[ӑ�*n"2�pj+mf�䃷#`!�z"�դD(�r�AyVN]�_^y������Υ���(��>�/?"�~}��_y��=�����CW���O����/<��n/��rÍ��|ãj1���Z�[��U���H�\�N�[>���v�8�����ø����E�ufQ����r!'�u�MS�;f�m=!��N'���]!�Uk��r����<`m� �V�D���������V�s^3oG����'f3�;���z�<�r����z�Nq�,���rO9��s�J�5J�� �8������HC��܏>�E���9��<�a��T-�Nl<�c�l8䧠��ẫ>P�27�@>�k���y�Y�Lt+1�p�oVdԭ��\���+�c�O׼QBʣX��4�[�*۾x��u��aw]:g��;���g+׎�ʭ~��q�ܰ �� 6�숑��Y��ZW<��>� ��]/��ύ�y:U4f�Wщ-��(!���E��[B��V�F�ϲ6��h��^�z��8���޲]L�Lu���~�WD�}k^4Sg:e���>hv�킫u��jˆ��C�mS�>��a�~����a����I:_r�����c���H]�h��6i��N�ְVd�&�Z�w��j����n�
a�	|
'�v�\��eĀy��%M�.���YOz� �R�)�A�ai�I��Ś�����	�������sKY�����������P�����0o0���ї��"U��а|ATP�++g�7�YHeH&jx�Go�yoW����Wu���<�N�P�w �;p��4�'�0�|xb���Cv�ܡq��H�E�-;iG�pD����z(k5�Ͻ�PЯ9M��w��7u@>02�l<�χ0�1F���z�lbjS��l:�Z�v��b��mMX���C'�,,Q�����$�p]�vCx�Y�1��!�7VokM,PFU\v�q{ܩ�!�їmRa~H�dp�a8���ƾ@kQCg��:#�·t��79�������O����J\m�b�r�>�ܰ��~#>֬�;�1����Zҏ#<���M���L\��t&`��yc�;���q8�nc"��=L��ƠKǨ����z{� �Ԓv�����s����A��=T���	����U�1N��6�3X�Lk[�3���T� �N��5"N�s=�w���e����	�P4u6)C<z2/��GCU���j0G�ݺ���/�1�?�t2Uh��kW�E�D�Գ�[P���
������pO�y
�J{>����<��1��1<�]v����s_��a��l�}b��6}��?ni}��k�8a�H�AGy�^{�{���������严W �""�3t�*�!Q��2�S��nM��Չ�,rT�Mu�%�l�����N��V�6Cw�Ah����;otE_ʯ��"
J�*Ij��I<<���<vZ��T䦘[���<��%�4542QA��Q�&��x-�1����S��,�8���#8I����0�Pq��s�d�0S����S�l�0θ��Eth�p�+�+8v���>>�گ��[٦.�V�M�Ly�"Gnl@�����p�2W,��7��Ҳ����$��\�*aD��^aQ2�W��EP�dQ�tgݳ^-]
m��2}��2ڵ8=����\��t�����1�qF=��w�"�s�x�f�j���~����j]&*�
�3<��?=z��+�yk��ϴ&W	쨠�ٯFݥ�����ns�ȹ�d��~a�Mj�*���$C��p���l��Tƌ�d�E�\n�Ţ���-b`;Ї�`}b�����Q���BQ�/q�����u�}�)�^F�e�ҧ��'y�i�z�,:*�8#KF�wO��(�
�T��ۉ��7b;b���zB�Qp�vm8���\���D#�Vu�-;�	�hh�:Ixc�6̱�$)��'&�M^@[.$�^9�����S-��h��ԦY0�0��m;\��PW��zu{g�<��[�_�bY�i��h��]G�����.�eK�N�6Ҝcʌnʺ4%�ݙ�+&��k��2�i���0��"�{eL�GR�J�V�Ֆ��k�
bu9���[���u�n�b�9�n.��}�ual'��;|w����ߏ���O̡�%i��*��
��$�|����|������Wߟ�X9�`|>�0co΄fČ�Jy���tP�5��ۉx�
�H]3�����q��-��~�A�����z��z�n|/@c�y�Π�^�O��3P*��C���k�]vi���ׇ��@���p��_��?2ԡ�5\��o�����,�[W2�(�e��w�8��+Ì������˨`�fl�a���b��	�8�hW�c��v]��MMpY0�PY��gpKW-�n�C�ٺ����E"�_�J2ׯ$��05i�:�wE<��e�L�L�TTK�������w��D$�f��G�+2ǥ�<�j��"L�7�����6�350]Jp�-^�#1/����h6�+Q>���� T�Y���d�c�̶d�e!M����`��U|���omSO�K }�W�6H��L�#
��{:d�zޥ��:('k������C��ֽ�j�l����E�'�9�P:������e,�uKjɲ���6����ޛ'�οk��I��)�^*s��e��6���v�rMH9�3˥��́�i��ѵ�P?<�w2���=�b;j��"�f3M�@�ݎ�So���W���Yذ ��{�je'�v{%��f��^��<Ѳ=��uԏ�o^�T�ev���V�Ծ�u�/�F<����w7�-�8���Þ\ ��������������y������΀�� �������W%Ǔ,�V>�RXK�\X1*�I���)j���;�ލ������I�7<r��v^���NU�<?1�P��i���n���˓�a�J[�ϕ���UB_voPt�Ϡ�Lf=�gσ�KP���O��x�I��z�2��CQ7(���=����a�VaU{��[ξ�kM�Iv�;u�}����̩i�>��6�:ܺ�o�y����%N-�����Z=���3�7:��=`h,.|D��}������U�t�P����h�c�5����n+�<�,)����=�:�Ń���v<�`;}zJ�%���<���ܨ\Wuan}�G ��;(X�,�-��A��=X=瀯*D,$N2��5K��P���/��펰�z��[��5��@�����۽��E����qNlA�-�	Λ���LN���.�Ύ�a� ��!B��W�:bse�i�����e���?g��ބ�}O�+Fj_!5�n�-��X~)��K�p,�l�C<GF�����[k��ĸ�;���N���c�`tת������򋯟�4����T������a�s\�բ�Mݳ��yO8��\&�8�Z��vF�#���Բ�	�Bc!5�!�U��m 9.�;����LɆ�[�3r�X-���m����C��7mwek�x5�(�ucE̴�i�ށ���{�UB��|3x3 ���� ~ÛМ�B�����f�X_f�:���⪈Z	�Q��{�t���w�0�C��v�ln���''8B��2��
Y�C@��I�.�%�l���"=p�H�n]G[����A�KwT�k���m�t�i}!��Ga�)�s��x�W��p4�kW�=��-cb�t�m\����𺉫-v�v.�K� :5>�;��xP�(,)c�9Mk��׶ʧ0�g�x�߽�oQ��ُ���^A�8�#�KP�H8��Af�ث���/���S���+f�zY�Cv��r�W"��_F����
6�z*��V�E�~���f��T���BP�'�e��[r�ɗBz�﫟")���ݛ�;#��\zL�{pZ\sì�am��;΃W.��/,/�ۻ��ڷ7!`�)�EN����.(VZT(p���4�]�l�Cf��6Jm��0����m�#�����0�hڭa~D�dp�a#53�W-E;la0��ޮ;v߬}w��j�4��)���l�+�C�+e˫9��s�nkMPpސ��㮷@R�7�J>P��	�b�t�M���VP�|k�
�]>��-5����-w�a��ͫ�>PK��A�=r��#2�-Z�
uY�!w�����;%�e��C4��K�S�kиAbs'zA]Ӑ�\��Vӹ���+�*�s 8LyjCF���6�wG鹈@���Ы�x|�`���7���TyJ�����<���:�
=�6�礷��T1 �vjO��4)�b{���Kj8�Pɰc7v��[��ax�	!c����୚���-���ps�;��ޝ���̪ɚU�NEU�x�\�άK�Vt�(5D��1&��#��'�
�gO��&����ZMKu��<�7Z�.��y5뵁�<$��%f���y�6lɱ0���D�r5�a�,�kF�=�!�{��{:n!{S�������hj��
��i�<�T���f@����y���o=2V��fy������_�ڻ0���̈.��s��N�d�hh��6Ke�$4l9��^�,Y��=��Ooyq��q���W��9B�m|�w繟�`,�=�m:�n�\�ٯb�2��謮��Q��Z�I��i<���<���cǋXeV5��,�߂٦]v��gK�x�ЊN�>�u����e�b�r\�'t�7f��L҆��Y ��%���x�S�t���������l���%���M��s
	E�@�g�-k��9�F>?r����;=��;^�1<��G�, ��W-}��n��T�Md��I�zU:�+�q2���dᝌ�J;6{�zj��-d 0�{�^P�����*�<�)}]�0�7�-��S��2a���n�/u��qM���\����)u厮��W�#B�7��������o�x��E!V�r�t7�b�C{H�Ug*6(\��&����q��iݻ��e��t�]UՄ����1A�L��Ү/��R~e�����R��\�!�Dt��`�(���Bg����*a�w9��@���oI��xg��:�1O�V��gՈ�`�Mǉ&��Fq�Az[��j�l��!7xE���/���=3njde��/�*�Me�1�I�ucߝ?"�>��&��en^L��iDRN�^�l`�l1�ϼe�Ɣ&ϙ�B�uF#��8��Ҧa�=��@���wYf#��yڕ�l,���l�]4q-�X�C��\e��7�}fQ�݁�wz�d8��|��;����#�s�����Θ�wK�x[k���av)�	��HQ�u/��z�ŧ��X�)�6���Ck��u�5��1���,i��*z!,h���5�d�??hJ��/�Kݦ����O�l}M�~��l;o۲��e;ig�}�N�"��r�=A�t��N�i8�DQ]1�$��LYq�4T�c �#����2�a�ۼi�+�I��@j��1>�w������}^�O������^M�������h��]�5��Pf�sT��;��ژi(����>c���u�O��'f��w�}�Bn�ذ�G�k�k!�͑
9����K�u�c,��Jh9s�+��1
���.I8���x�]����%�p��7�x��!��(���nՈ�o_n��,v�˺�noGS�e�Λ�3�t+j����1�#Xy��3k<*G�]�*[�h�N�چ+�̜s_v�w�R7.Fb�9|K�㏜�.���*g��v�5�7�I�B�_q�WCU���X�wI���Գo'֜�����:���B�٧�;[i�SiLol����Mko��MS��]�M�Ko��3��V� 5��٫�2)@k%.U��h�)L��CJ��Y،+]���C�C�tN��j�Ы<w��.��?e�����w;�iٲ�>�)R�Fڡ��u鵔j�I�14��k0�䴡oV���&����G�1�Yc�Z�]+�&M\N��^��,A���ˣv�x�7�Y%�]o@���|V�x�E`f��ӽ+lj�E����2fr�Ab�x�R.�d��۾2���2�StJ;�%{	cS�η.�P��:��9{F�+c�U6��襲ol\��K�*��Ao���=��Q�m�k٠�;r�˶ѣ���-3]'&�L����0]��9��&h��yj:ʽ�F��͜��GueZK��v�|��+��"s�6J��*���@ԲK���)��F�5Ư+Nñ�fUǅにX�5*��7[ptM���N��8b�!�|eENûtxI�^���y�.6_ �5Pe�`�;��k����'u�-�h99b��0���w�c\N�p�܈�(7Gsa�3���X̋e\A��(>D|e���j����e:�P�@��!�j����Ͷ���3�s�;�Y6L@dL�ou��qm��8�� v����[�LMJ����ZmM�kf���|c�����_K�/�\�
슟o8���E��z��u���j���u��,��T��RC�����z��p��M<mܭ��iӛY����imf�y�)�]�i��F[�q����9�J�3�c���Sv���VVk}ԫ�RG?��̍����n-e�WSʺ�t��3x^ճ�p<ĝ��$�A>���iTz�wOP���˓.�a�֔��ѧ	�R���%ω\���c�IO�m9��Z��ͱ}H��k�� Y����h��w�Ҵ���#h,g[�Y̮�X���[����˻CK�
�Ur�����N�Kf��[����M�y�F7���P����q;�����	-m�7ƖJ��ϙ�ƕ�d
3Jɚb�E���;#<�r����n=I7��]e�wd��vg@J��9�W]�w�P�w�O�RE� � �g����hJ{je���F��F!�i�b�-DSE�f�*��#1�-�ENثc]�=h����袨��
+�vh�]���i���vgF�0Ln��q�ELEM��	�*-��DMcj ��;h�65b�LMk4Q[��h"&6��']h����J"��cl�TE;�y�.��Q��m1S�F�XثVLř�EѠ���WF�Z��&	�b���ݺ�]��ӭ%1TƋ&�!�#���cZ#����ES]X$��b����Q�;�tqkQ�G@tQ��`����m�ݓZΌEE1Sv֍u���]!�GAT�DD�3kh{��4��ѧN"j��1QX���vr�y� �nG�E�i^a���-�i���9A��1�Ƿ��TÛID�c��n1+�.L��_W�s�穼aD���N���5�Kd\|^�&��m^���׫y�.���g[��G�#��A;R�ZŒCF��w�2M"Eٷ*E�@��q���t���K����r+�D�Ƀkkw$�+a��^�w��+���V��_s�+6=l�9��$n�vC��b���bDD>/<�4md&��޴�'I�.�O׊E6P%V���W�����w�Z�s|}pl�G�f��A�����<�4���a|�w���l|��{U�+kP�r�^�|;�o}(¦���,j���z<����`��v�Wq�,-���ń�_RR	u}p�����_6���8^I��r�TO�T^��i������s��lz�⩑f'�������Ϻ)pіv)���v���}T�M1���zU��A~��T�*��ʝ��<������PaMX����IL�B.ߧ֘ķ<I��/���?�yP�r���*� �!9w��kU�3zŽ!hb4�e5��Q�+�d�/��5����a�k� ;c>�����K:7��GYV&��U�Yԋ�/���y�-<NV��^�O'Hy�4kL�S���߾xoˆ�cP߳_��9�烾޷y5
#Yz��N��Y�ײG+6K�oX�k���*5� �l��q(�7Y#{6�Q��q�����A�!�ްtM��V�}��#OQ��"����>��֜�'��C����F��%�3���� r���.DÃ
����`���Bc��!�9��-9X�.khw1��^�<�(��qA͉r�a����!k+ܻ��f�s�
6Ab��a�����}���vf�/��	�l˫�A�/N�Ze�Z���=���y',�hچx��i}���_��?ٙ)���_����/��a��ۻ�םoVM�Jl��#v����J��i��/k�N�~��FZ�i�u׽��^�������{G��~��8�\��	��b&�Ea��(��6Mz#�T���7��s<�	�:��m1�-��l$wGc�� ���)>�	d��3j�"�;���!l��vєE���ػǿm�s|n/����Ī�����RϯX�l�Ai�X�U�����n����2��Y3�ҕ�s(�sl���@4���Y�hE�(K��`������g��>���"qP�uC��F:xډ�7����jP�VV��>��i{� a2��.C.�m��7T.4Ǣ(7��Ec����������Y�}��ޥN�F}hANd��e/�k�T�1-{�ŝ��9C���W��V	ˇ��}��K��*�r��;��W�#3^Cp��w(�I��j���G�8���r� �����+�ট �Pv���G��w���<�\x�4B���"'���b�y��v�R��x��x ��xd��t5���l>��s��*�/���z،���B"1�2�.Cs{��<���1A�M��ЯY��06j�c���؆E�*�2O��Jdp>ƌ��aigO�Ɇ=��^.�:`�-09�� ���m׵[IT�̞�{��;:���6��XH�nY���$b��Zhr:Ha,���P�����<�vi9�Քr��ƧS���gt�T�HޞEY�-Z�ph��#�3Q&���=����i�����d0Ɲ#1�T
٣��z����F��7���U6�]�ck�M��;��'���]����L&�_\K&;;��Xs�(8���������nE;0g�:-�B�-����w�:�_zٞT"?--P��|Cfgti�UP��ʎ3	�A�!�AA���=0��S�8z]�p�dDʜ."r
w�GH�Нj&���sY���F��������S�|w!�����!tH(�l9¥�5�q&���]w~�3ww��z�!5�9�^�ڑ��e�):a���	i�jlS���]R����/�~����Y�յ�	�ũ��oZ�A����r��Gwu�����ϛ��2.��^��'�C�+��}V7f�ۭ���y����֒M]��2��$�c/g"��j���Q)��k\��P^�=�0�#a�z���"G6}?���Z����g����3�|j�:�%�i�T�26��sX�D&Ր9�J�=�Z�+%>����u1%�V���\\�d���$ذ7EC�L�FM���]*��r�Nid����IDD���4�z3����v�J�v0F]��;�6K��@�D�2���Y�K�k~����U5�{
,ұz��L��p*��.)��� U�9�ɷ}h�]����\��rfZ�s�B�6�d�X�Z�P��:�\i����Z�T!��H�o��ܽ�;8��iq�e��-+�IDr;uy��e�����q<��j4��2��*"��_�@ڔ,~n�g��؂=��_ߞ(��7�pT������ڥC42%�3��Nޞ�b�qS��>��^*t�b{.{^ʞx�����F+�OK�(봵�x�߃��͙�����nĦ������O�*��8sH
U��7���p������b3���?��1��z���3�	h�<�;;ucu>#�L����U�lڑ��B��i(��=���\��ns�:<����@����9g�U��?��Jh�m5�z_Ӕq�X���J�v�d`�zt'_��/��C�D�ק<��8׭��מ�������!��٫5co:���7 (Θj���s����;��(=�?��\�;S���6s+��@�6e��|�5�\�ި�Y�Z��mζ�8	�2���$�|8������tk�+��L���:�'_������N��%.��g���}��憙#��a��<�U�uu<|��đ�(
�:z"�MG���̸=+��j��z9D���h �:Q�]P�<��=u���P�'�M�Bӧ�e�V�L@]��z�)�%�c�!7�V\?�l�/c��O���sv�Z���4HJHe^�,��B��;��ܷW���|0L���'�%��]�1�i���}���A�|�O�y�/�c{K
x�W�B�l�0R[q6k{b"{]��į����At�Q@F;��j[pvz	Y�S�E���[e�t1k	�m �U7X+kZ�yt�2�����.*�EX���n+�/ߏ{Y�!?nV��M�c�g>�A�>s�o)��-yGm8��Y�.�W(�8/	
�TX�����+ЬɺQ���'�W�O���l���0e�y�U(qq̥k�*-99���
X�ن����2׸ܻ�����Stۯ~��)���g��ϖ����s��GrTZ�̄TbzO�|����O�zO�?Hc�
|�U-�Zs��+�i֪��bȻgKvn�C���qI�!LE�[��j��wҤ��e׈ʏ�ψ��Ыmh\9\Ov�3w[���m�ang��]��vVEk��[w��Z�F�Y���0g1��q�WX���m��ﾪ�s�4޷���©�xw�/=�g\gE�_CxG��C*�ץ��:bķuBⲡS$8�M�e��TսQ���}�p�a6W��t�+H�������U�w��_�BI^J�a3��(�ub��V��y��wQk�&%��e��=&y&��#	�S�b��W�,���mQ��z�u��Z�T�j�����g�4LW5Cav�`�X;��8��U���&_c0�b6ч��L[O:�_q��3�Ɣd[p�C�UZ�L`w-CL0`��Qc�A��g,WC��ƾm^��$��WN��;��J�O*�}@I�M	}��lW9���}X�A�`u�u{!M�22R0M�vPb=
�>��K C٪>�~��L��N9�̑��)n�͜!�[��U�0��g:I��
I瘐O����,�yw���roV���?5��|�.}"٤���B3n�ͪ4yן=�1qȸ�-"j����x���n5��MQ��5c�	̤醢�'�%k�.9�n�����HCPoZqϋ* �9!���u�y,��l����y�ehw籍ݔ�J�R��rŸu<�CAvMӹ��< 2m�	��K3�Iw\������ \V�:]ݚm�֜��P#�f�9��+�v�y[݄��O3�Z_q��d|z��5�t���gb�͉�wwx������8N�͒*��?�r�*2�nb�a0q�P�,�/��Э��8D���s.p�#sS()�U��F�P^��=������nԿx��bk>�)6f�Myc�9^��Ք����u��-�d��׻�̧�k��8bǣӠ=��gi<W8f�t��\w}���7���C�wDmwY��%X�M�uUCj޹8g�p�����A�>��۷0��`5�T.#��[dm�+f29�����n���ث�[2:*��h�7��b8L�s�k�Y�rފ��k��{����5:og� MJb���Ȳ2[S�q���i@��*	�=B'���T�8O
gV�b�yq3��L�4۠�+��\��1�[}5�֫C(J�L_C;Rq ؖä�-`=Cظ�T�ǧ���v��mT����fsb����b��K��b�r��;�aPXp�K�Αӎ�����#��o�n/e�_����~ ���Kߩ�(���e"3����S�2�T��P���L�L�LC�\ټ�k��2����C��`�k��_�F��4ɍzyW5x3z�	zW�-�����c�VN�6�B���e�}9}��~�t�ϱ���P���8V��*t��z­�a�f)]�\��6Fl���C�k��>�*��ΰ�n�3J�+	#{�������z���hi���PČ�n>�ٓ�hމ�ʝn�b�d�/2gb���U�,��^��n��8�j��V���AzY���`��`���@����.8h� 	���'��!ñʈY�q��G�R�MNji�o��Z�_����r}3�-P��>�����*�`��'/�/�*�����s6��$X������:z��N�ۭ���HB.��J3�FP��!w�*j/�,|e;��m-~�,a��T9h�lSd��]RCC����DYF=N�cVѭ��/��@������FZ������:��Z��^Y ��r&޲�~|W�W����'�d&��ܼ�$؏A蒺(� �'nY��z�(Kn��m���$���tm<om��4�֣�{ٖ.��r�Vq-�kY��ey��ֶ�zC6	e׼������,�����@Xw�EWQA�3N���!սx������vд�Zs��w�l�4��:C��A�x�B�3M�{/)����Jhd���;M���jޠ�uY���KF�z��QQTF�8/E����`H-#�LPz;(��4����/́?6$�]�Ѫ��z��Q�;G��`#Ҷ�5�.v̻��û�>�cb��z`�}�S�Į�L!N��i~�>�[xܔ�cM�s�[�Q�GZУ|{j;u������t��t�Q����WgC[�0�"pح�;1U�F悳���2)��=�_uh�x/z4�zӣ��3���tP��vm�t5l�q�����<��hNۇOϬ��d�U,Vo��P���L��
�P�����O
���?*v��yr#%���.��n����ir2�a�;��b��b���,�����opgǯdup{)���%�3k�+�k���S�&7fpjjr����j�d8�E�K�8]h7X'�q׉���S�dʔu�r��C`���&}��B�Hد��5�[3�3���g�!�lW��CWm��)�Q�����_���4:�����3�螡��͗.�u;���-+���lv����_g�N5�y�''����e#��sm"E��Y.U�9�mKV��u����%fkp�l�^�O�e���^eT�n�h�%(6�j��D�bs�L���lTHU�!�^T�3�I�>�i���Ŀ��Ƈ��F�O>�̰~�7���g
�-�d�kבɦ�մ��k���ʒ�*��b�/�0^!\c�~�~�}��r����~��>T��7is�fU)�0&��'8�tP��'�M���_���{���n���j
�i�y���v���Ɲe����6C�p�0\�|��`�ZT��R�DF�LHj8̡���j�Z4B���{hw]{�H��̴�ƴ����_��^ǜ׌������|ĝ{�t ɩdK�L�m���F,�%�3Q`�٠�P�7ڠa���P��ٓr�	�;p���蓏{�I�>y6�s�!��7���>��.m̕tݕ����MSSC.wEY��f���������CKP���1*��g��'9][e���^y��U�L�F�Y���qC��?�����8����#��O�>^m@"u(�<��S�q�o&  ��P�0���t�,��2�$�w�hy��#=�_P-���ܪ/�Zg�Z`���.:Â�5�d�9)vwEJ�r�O�b�[($v��09��ZF���=Q>�QO�z��3\�^��������.n�s:eЖU��]���	�=���pl�A��ptk��H���4?yL�:~G0j� �}ӷ��暰%��Al���~P�}�Pl�Q��*�<� 5�C63��6�g�1�ΝB1�4U��A��g^g�~j�V=��l^���WPƫ]!�Uk��/Q@�c�U�Tf�Ⱥ�`�D rIV�!�9���23���gr�XcN�`�����s��}~_������g�����{^aWX����ح�L���OYA`��M�ڣ�x+�W�l!��s�,�dީH�n�O��ws��T��: ��w���]gh �D�]�ӂS�m���S��'��	p"1���<�Jװpۻ�����J�]�T��TvnA�w�ؔ�V�P��`0jo��/���ժ�ͣغ�P�Y8
����p��c{F��n���J���SA-��Q����2N�y>Y�:{��M<Xd|�kz�і(qz�V�(ƣ;gnb��J5��C�1�:��q嫵:�.�Bn��1:��o����]cIvf㍝��'����]�P'��t:�+ ��.���wV��7u��m2.dZ�VGm�(�\C���]mm[��#o�su��=a���;��}��Px�N�/]�1�x.d땤�v k��ޭ�D�O�0���\SR����B��f�N��0�A�t�m"Rut,W����5�)ʯOn���:;���PY�it�=B;2����vX��k}��uU.����7��[�rS��h�<��<��MgJ	c0��N��+��4l`��&��ZK,^ʝ�N
v�<��ؔ��r��`�S5ȨЩ�]����km�iھ����/�ك-u<s"]"ǝ��u����ʄ�+���ՁX��H����w+����\Bkϰf�F���E�H�B7����8i�f�A�p�r���L��ד/aw�Rٮ�P\3���PT�d�V6=���k)E�jw�����PT�Q#P�%�mK�qvX6ze���Y��ݤpk�&���Mm;�5�M��'�������|�L�m�ff�����N����wv��sF�����2b\��u�����"|5�u��M��gA�EU:1Z8d\d��:�>��BؽU+y��46K�S;z�C��=���Wp6OTka��\9�8��qr[k)oO��0���Jc�rs�r��J:�u�c��@_��e,�935�o\uת�),d���4�!�1�`��M�N�ؚ��C��1��P��L����;F�E�[�;����h�+��Y=�("z��ѪS�e��A#x���R�l�S�C�C<�z�V��ͮs�J�N��0JrfG�P�Z�`���!]-Pw�Һ�̴�P*�Cd!x�S���^vs8wzDg(E+iZŤ�#z�]�sdA�i����Ke�s������(���}BeQ���A�_/��t"K-ڥ�V� �$n�ਣ��q�]N�,�v)�[rK�"��s����R*U�spuM<��2��|靘���ऻ�d�(��;��b�����j��SL>���Gp�xcy,�br��mF�̭�I=��KlY�L��Fξ4�/5A�"�C
�bn�\�huַr�M�tﶹ*����XP�p��1Ѓ��c����:�iTo[�9]�<X;�YV�\ �N���`�ӗ�j9�}��C�]˶�#��{sm"���g�L2���>�.��A�m�01�]���S?|}�SM3STZ�l8�c[:;���qC��Lƃv7d�MS�ZT��;��5.�)��mѩj���A��")"b혒 ��Ę���c�ƶ�n�F((�u�Pj��u���bb`��i&�h�B�9)��"���������T��SUME5ljJ#F��l��-�4QQ%5Om0th��ZLSEIQk��S�QQST�SMUP�CF�%Wcli�b:�Κ��"��l�b�����{h��Y�����""�cX�kl��TMACDQU%I8�*#�j(�")�cUEU�TQEQT�Q%EUq���U�EQ�MAEQ���H�&���I��mSEM���D1D�DDo7EI1N����U,GZo3����&*h�l1�&v_�󗖩��fM����]���EOw1��X:���mMLV�=ox��C*�
ZX�u�y�a�Py-�S%7u�߾����++7��_���K�4Q��n��(��jzC��觱�5q���Y���h�td��{ c�~8<ݗ�ܢ[�LMP,�	�� ��k�(����n��3��<,:�<_cq�q�?p2;��[S=�H0�(�-����a��M��dq���/�j�蠮�[ �O�3n���cY'�S����I\�K��h�;���my7�3I�m���B�E���sO�*(4�ug}V]0N{q�o�CEΩ��%����xj���H�+33j	�G��~9 +�~��J����4��i�p�ބ�=��)>�Ŵ/m� g'��aJ��Z��&�%T���Y�4U������E��A�G����l���E�pX��l�h��6�r��z�b�5�pu�W��f�3(m�'/a�mᅰ�*_�]� ����@b��ς��W��&;���U���jZ@uk��s��E�,*��{uKc��C�Db���ת_�n��J5�*p�mt��;3�a)�#b� ��G�<��M�E�(XZr C^=9�ccn��4�f0�}�w�@ k����u!��ጹ4�����v�[�JwtИ*��[ώ�-T����۬��{��Z`
����T|�K�:�gA��c+��.����Y�}���{4od����{���8f��}�<�2ݝ9ϐ�Z�Y/9���b��ߞ�uOgw���c-��y/"�i�_i�.��\��2Y湅�,��8��5�3��.j��Nr�77 �>��E�"8��R7۾�ަ��R��U���_c�C/�O��$u:�4bs:�]�¸�яYo���o5P��-���ƕ�&�����KYY�O�}��*.g�xV��(�qf7��Mq��:�" ��}@\���N��՞�"�Ю$Z[%5�s<R�,��;��j���K�">���;�?���>���^9C?*���X�WT~��Z����X)yj�KZc��]�A���g<�T�,z`�^�����g���*6��/�z�� ���q�237^�t��a��M	EˢAF[a�єV��]7rk&��{u�Pk�a0��A���Y�;>̘V�r��k��@oՉ�����91�MU�ݧ�"(r*��q�ꌴ�&j$m�)�S�U��(,��c&�����U'�&��n��?ϟ�ڍi����4��iw(��b����4�R���Ƣm����i�����i��2�e��~�Wk9&	62o��;�<%5����jB�e�̭�,�z�7H3���Q�!L�>9��aۜ0hf'�m�s��9�c�(L�n������T�7�h�/-L���jE*�6Q�&=z5�g�d�?۸ƽ޾:�_6�|��wX�Z��	-���b��%�*	f(�04x���>wS��7î��n��ѐ��B���!2�U2Np{T�j˛a�J/"�uqA,,o�#���݋�;���eZ���J<ϑ��4��7a�u�#�,{"S�UJm�J���:N���c ��{���L�'|S'n�d�]��!3�A1��Zf���8�.+�iW'.�[�G6�%��C�zX���/��� 6I,�8<u�jX�wӁ�;E�nڗ��xg��:�x��8�%+ �����T�9�JF����4���������ں�>�$vbS �����L�j����:�B5,��lg�
H�.]��3ohLh'��G��U��:n�O{��_nN���6���Fּ+k=_P�%�)eyڤ��j$d���dDh���an3z�`R�Y�k�ep�	��\��d�U�O��->�g�`>h��$�1�QίPl�ꢃZ�WΨ|E[]��ˬ��̩��Ӱ+�g=zq��Q�P�z�
;��Okǅ6t�q�d@EO �������-��y�RcC�L�.����f�m��]�����T�����S���̤�,}��B�Kjor:��f^��V��/7��]SU���9�}��(;oqӣ]"��׏� oi�R�2�cq�����>���r�<�����
�^n��v�6��E'cy���c�CB�M�\aQC%Ⱦ��>#ss���do474�A����_;scE޳ʛ,S3��fp�8 �x�Oj�x��i��d�o��d��Ϸ��h㽁����4,��Qe���`Ψ�΄�0o{^��R��O����|�m".z��{��&�)�fE5@�3S1�sc�s����b�C��6�Wמմ�J�i����df���Q�qS��{���7'!��;tӚ_^�ۍ�T�獳c�!̩�h�]�#)���U�u����W��eJ�>�)���ܱ�{��5z!S�f��/�BoP�'��Ruς�M��FE6r�Ǣ��rGs��*X����jadmi�Erh!���OE���.�C#�Ga�aO�s���J���TZ~85P�����ᆸԨ�Å�+-��ʢ��>�z�|Y�3�����M�-��4�O
nwe��"q���E�4��3Ri[����Asז-��%]i<�e&�TO�U���~0m����g�ᔲ]��0���7�\��=˞����9I-�U�v�K�8���l�(�w��?:8$e���mP���aSM�(+�(7����[R]�V:?Z�ID���h�,;��5;'-���=��
h�9g�Dʠ����/o�o�/\�K���r�6��qZ@u*5Ѽo��,)��Ƿk�����vmfJK���3s9��"/\�{Z>�@�b��u�n��K�����r2)���z9r�S�G������&0M�8�C�0v)�1.k&��-��k�n���O\佊z/&xл�L7s:rc��Mߛ��u�a�`�9�ú���/*\U�^���0�0��`S�({�>Q�a�:[xs�-{���5���Uc�cAe9w��tsV?S'�aAI�	���b���G��ڨs \���_)�R���q�{7�y��R��E|IX�-�ʹD��	����E�_�.T _}Y	��3��!UwS1�D�tW+�%�uk�@k�s�0�a��|hy�/�_�(���T�����H����b����~3�exUz'h������VLY#�#����ʤ���S����c�v���&Ü2���~�Z�nk5l�l�	�v�k��q>�tÜ�N�d� ��*qEatQ.#e͞�:^��&,#�&&��8Y;s��Y\����2ľɊ��:�a�؄��A�0�JW-;�a�g��xq��n�ک�mtHu �-���y�x&g���2ف��>�!B���a�l7�n�a/Pbmօ�S��Ф0�w槸����]^�e]��ג�5���vP,m�b���y|�=y�Y�Q��
�<����I�}���%�j�|��%dW;����[$�6�8R"�
 �	����HҴ�e��;�Օ�B�EJ����"��70Wnc"i VO���tT�oc7I�@v���m�aƠZ�߀��8cld�8WW���\���Bl��ȇV���d���V��̲��l�]s�f�������Gl�0�؏.�r׆�sbq�w4C2�I{fRu�'�e��G����6�yLE�����m�#���?eJ�[�;��ӑp`4떎t;uE�2�0���s� ���h���N�����rc�q�j��^���Ǧ�G)iR��hL��b��%�
h�N*2″j�����G<b44CZ�@�Q���68_
�V�{*W�hſ�wҳ�#�	�����j�vr�%�5�2��6"릅�b���+ѻ�ڇ8d���gG��3���昇��c¢�=�QoJE�=�2v�	x���U�1��n��m�)�fF	\�W�~�A^���.�
����-7�r~��]���,�CL����>V���-�g�hߗM�[�c����:[]��$ztdw��uiu�����{k��Y�gm�-/LnkWd�5����|�^&3%0��pJ�ؐ\���{y9�{��ȓ����߸��SQ�Eez��d1����Dp�p���P"�:+�ma;q7h���UӃ}�Pt�f&�x���خoV��%[��Z�.ˁ;8�������N�,��7��nv����B*����3NWc�{��U��"�;g�3{�
S���Y(��k���l���|�m��H�;�<�`��'zҾ�m���[N�?��I���H�����)߱�Ň�vB�^�cA(A�������=���&�2�2�I�X�U$4VL�-q ���bǩ28̩(�����i�6xO����Oe���8�q�n��t�)�_]
ǰ;���ܤ��,1+6b凜C�v��{�XWޱ�'~;A:Ȝ�����3����U�ܶ�Yթ�씮骖\�1F�Ze���Ǥ�A�����w��S֟�M�,c����+zd���UL��j�*�l4��z6�[�/,M��[:;v�]���VNf'�#��C��]���ނ.��W��/�_�޸v���:4:]�Y[��uU�8��9x;����욼C��p���^C��iҢ��w�:��x4�I�W�&��{N�����:v��_�IG4k�;-y�S{;	�^⫓�}s�Y���&M";�uO=���X�-����]�`h��\g�"!o���L������ت��Q�>T��qu�yՉ��j%Zߘ�{[��y:�
��P�~ s�se ��MÉW�|ww�[��I�$�� Q��VmX�c������!�\����J���T�V��c���ڄ��d]��؛���cQ؆BT��9[��/)�JZzB�W��.[�y���a�ȧK��,u�<�Ls��n�4�w@�?>������0u������b�hdz���eZ֩�U��)�>އ;��V}R�',+�ݖ��q}D&Eζ��n�}۶��y�|fvI��G{H@�uM>M>go*��-ƈ�DZ���7����w�������r	����4D�Fe�;M8rc����쓺�����=��m�7�]�F�,Ų��=,�(�����O�zW�P:,�ILM��,�nn�e���&"�j�_����c�p��g����k��~F�KlQ�����z�_N�*�.�h����ͣfU�	��2R��V�|���u���6k0��n��"oT[ޯVMms���@�񅲕�w+-�i6�`��I����f�ΊǾ\CƊ�r֖�5yҖ��;eM�Y��ǖӐ��u��P��g=�.E՛%vW���T��ŷr�T]��Ru�P&�G�P�82�P�w1��oSW�jE*����<���E(»�,�����$�/h��P�I��X�,�������Iw?�֏�1j=�>�F���ڽ\�͇$���8��֩yy�-�
-��з��:LCA��L��;����<��(��/ړ׌#���yLjzF[U
�:ٛ�Zk���x�^ wr���["�=Wsj]w7';k�y�z�$�S,�����֧��:�l��<��2��7�����g�²lZ����cߘ��35{��g�GM��r|�Ψ<���]���?q��~�8��fVt��q��ѡͯ}Z�;s��&8N�#���Эl�z�۞���u-�R�>E<�ĞÓ�Ґ�ΟD"jZyǶ4Էr+H�U�����B�tN�GV�a��\���?�n��;�1��z#�p�p�㥹]����Z�~����q���4����<l6�o�@ȯ<h�yFf�8w�ˤ�^����Z���\��o,@�ŝp1��z�㳗ƿ{��#�>2�f���4m���M��{֟"�#MʝwCi�c�znw�����3�	�p��o�u�a��)G6��e��C��v��o+��ܾ�����f� ݭ.��L���M����j��w����dq�z��Z����\�(��bo��ʓZ���Ճ��o���;��|tJR����K0I5	���הA�2�JnI��P�Lк�jmZ_�N#�\5I3*�U���K���y��0�mE]�a��`��xf�fұ�(���fv] �1؀�N�ƛOm�<������*�5Y��꧍��mg �|�y����]y=�z�P�=^Kñ_�~�{�v�N��+����8��۵�)��a��
�7ُ���l������ėq�C��lt�g���ZL͝|�n��\8��OS^�3�a:R+6nV�5oV�X���u_��_���c��S�	׈_M��c��l����נ���f�ΛIn�:�r�������~6�.Yv���*ӯR~��������wy%��Y�}��u��Y�����'���۞�U3}�����^J='�*��ɭ�bܵ���×�Ek]���y�í�,�zD>�Fu����v��O�^����=��O�����=�������	�����B�Q {#�	����e]�u��w �	�O�62\�gΌ�B�YN��&�f�L���}{�N��-p�.�Y&�-��u����r�H<B�췘�p��{ w����ɕ˕ob��q)�:���a�w~�z^}r��!73[����C��W�yR�&Cq�뼽c�ǫp�$y���9^0/��r�F�I'g_e�f��-��5Q�=�K�v-Rd޳��hm�a��%!4kE� ��ڲ[Op��=��͸Sۜ	ΧG+onQ+TH�:im#��հf�X�;W�1�����K�}��	ři�%�|��r�o�@��+IlWnH��6���Ҷ_M� H��{Y�ٽyR�K�ɛ��{�۳s�8td��B�>,S�<w��(R��\X�	6�n�QP卭;�R����X�,���;��Xt1}�0wuE7�R���٘e�}9�,�@�����ׂ�<�d��5�\���N������o�
(5�.�ò�њ0V����:l�K�S� {@%9����e�P�`�Z�'F���z�@u�wQ4�((�e2��W)�=�hhh)��������Jd�ٯ���4>˖�j��N��9��}���ct��q<�x�k�릜7N�'�pc<V�z�oN�0#څ�q�fo
�Gj$��_J���7V�:�kC}m�J-_�bk��`�ͬ��u0����'Ok�	p��vJ�@.U|��\�pk���g�{c��L��Y=ƭolth�x	�)d�x��.����Shӽ��I��u̸w��[l
��_q�j�6��v���v_��Y�����3�:�ҫ��{8�SJ��bT�����Z�-�>�
a��Kf��g-��jR�ha��L/�����4�u��\��Ӯ��"�Q��W|����4�|�F���X���g�ԹQ����&�8�;��T��v�a벒J�	���]�*Fŭ����jm���ۼA9���}1p��ao��]qh�P]צT�N��ۂ�Wx����@�$��ubh���7,�)��(��[�d����0�N�+ϓ���$�����]����v��`T��t&�kk��|Q1(�����C��v�a��VZDt W-��i�Q�=x&K,��u�:����1��}4�]������;�g�vj�th�iV��YX�)�Z���h	4�C�q�h8+ 1�|.�T��>��2��L�" ������2�tW$�+��{mZ���];4��
�iZ�9�w�lR�#��p-��B�]�P�ݴQ߀˫�.�:$v
�0Z�Jf�N���YNT���y�IW�q9����d�Z��-	[��49�;��3����)��:�,�OA��{$����Sz�u�'�����ܐ:&R��\-��B�G#�c��,B7V��V��]�{t/^Y̬�Y]B_��
]	��f��q`Z5��M��-e�.�����t%5�tv���f��|�P|��A��QPM��R]�4Utf*��Š��4W�44�T�QIO������.�"������,&�(b����A��$QAD�E��Z���#Ͷu�(��:(���h�������0ձ�mD���kZ�bJ(�q���i�0�X��v� �JJ�h��Em�&)֨ѡ�δy8""�,��t�t>cT@t����B��(��*��q%D�4�ABQAIV؂��ij�R�`�ӎ5��1���"t�+�@RT1%�AM�AAAMDQOFf	�(�-#AA�2��O����]4�OX�����`�X$�sqi"K��TI�+lR]���h���k]�y���&�L�DSO��C ?��ԡ����D��jʆe�٦j1 ��U��l�m�' ���>ض�A���X٨�Cܮmm"B՝���R73olEthx�s���%�G{6�v�`���,%K��6��ގY<%�&�r��h��n�z���H霐;�9���b�F�qiG���s����PV,0m�{$�Ӓ5�-X'i��cɘ2�A�H~ti��YV����7�nؿ�uy���\o$/���u�abt�	Z��a�GCa̭n�	z�k��&ޮ�ٶ�E5k�b/N`��g����A����PFTy�R{�������[U�*��E��a�%� �R#��7@]�fNTf�HB꭭���3�{�w__�(eNHy!G���{Sk��{fTOk�s�tﱠ����_*WW���JQ�L�V��FqH}]��=�T�5L� "����dN�dQ��u�n�Ec��w �����Y,�ܬ�bB�����;�Ғ���5fƙ�˹��	���d�~1�P*V���,t��-֏v�6F��F��t�)�1��u��L�K�EQC�%v �k�.���mz��İ]tu{x�N�X��f�Qv����׶%��,��i�u�m�^'��[��9<��Yz��{1����=�0�!�#5�;]�u)W�&���>w�j�w8כ�x��7H���a�y�=j]a��\UƫJ�B�����oAx��P�x]߾������.��-�5�{�[��i�נ<�HĲ����4�契����9ƪ�5��~wW)ޟ=�b-O�gX���uq	kIc�G����kh�eϹ^�h^�}�4��p������sU�)�0nc��1Q&��^�0�PK�]1FS@�B�x�m,�{X�Z��O���Cz%)���-⫸��gXύ��6���'Ɉ�����,��(�k���`V}�z�����ֲ�5�n�͚��6�Y��fj��9����}�r�b�9G�ٛ��l�~���9�$���'��x�K4<D�����&/D1I���|[��5�#�U�_dӍ�u�s}�ܳ��2k���n�޸�Ŗ�Ո���qj۳
��R�][��U�r���a*��yƦk�Wr*w�Vu e�{����ھgl��EkU�X�xPA.��u�@�;Y��X`F��q���k2m-�N&������wB��:��T����J���-���s�Ñ@�s�ܫ,��ۢŇ2vP�K{��1X���c�S�<���� fed�����+ځ����=�{RSzʦde�D<d�R"�iF����ۻ�zW3Y�U^Ott� �RCy�M��T��y�Ʋ�j�F���lg_m�S��J�B{`TL�e��N�K'(��^�j�qB���i�5[o�TD&�M��m���[����ƥ��&��Y]Y�����$^?	�~y93I���@�mЫM5Ϡ��ᔳ�a���Y�:��ŷ(M�;Ў��&����6^N����t�>�/�y�Ԭ:*��3�o7ү��O\_i.�E�^jYUה#�>���r�G��8̋y�v�HWQ�.�+sD�=k5ǝ������~n�H����rYg>��+�̊�8oF@��1��A�g����g�R����V�6X�f����Q�:zw��[�p>i�1�LA&��oMWr(���+��':ǰ.Mn�!�=;��OS�^�:�퓀>��eEV�Yz1�
���m���x���c`��|pۣ�>mWE7���/�Z�1`nt�s���IX:o X\����N'K�oV{���7}(]���H]L�6-�ǝ+�ӠL0����iE/�|�)��a�8d����j9�q��H�,Ƭͪ�0�1�^m�d�[��6�ZH����>�=�L3[��6(�]\����ו`�����M�"vS��a���n�f$�4��0�c�I���^���}
�$�N�v��_������Q~�Au�k>��m*�/StP�t�Z9D	�7o4��6�ƹ{��O\�i�/.�)�|B᳚Y�*h�	�8�CL#A��C^����^g)MWv�佣X<���M�+ ���i�$�vT��@�sbZ�����^Hu�����GK@�a[!f���@�~��,��s՜ё���\�������3{Z�e&%��YF�}_1o��[l��T9�08�ʛΣS
�{�.w�ҫ��n�v����6�L��"�m�ػ�S�Ԉ6xDd�s#z	���*�s4�h���k��]��7�b_h����<5~����9H�*Φ//�2�}��s3����|�=R�x���Oo������"�Y��K�� ��T�u����ԛ�o#Y{ܦt��fܬcV��)N9G`��Z`F=���۴f�}>�C(X�J%0wDr-�sv��/9Ϩ"l��W�D 9GfVϕ��ห��ӛF�m�g������9�:Hu[��,�Yv��J��Rh9�w6�-�����neMK�no��>G㲠H�n0}��o��w�<l�O��j��<����T(�Ӵ`��wn�|���i� F��l��y�k��u	�/Q�R�����[?^n��vփ�I+,`{��3`>m恮�D����
s��&7D�i�ۈTz�/��X�^>��>š�+��qʹ3�I[��et6��7[/��60�_�M��m��2�im2l*����EKښ�M���6Z��-����y�Β�� ��!+R�C6۶p��8�$�ed�e�W���9
E����}$v�ޝ�Bi6�?��u�qh���T�i�vC\���T��7}����4���5���_�cE4��_o.;{CΦ��
�:��
w�g�z��e�J����o�{*�B�G�����YT�;^�q��M�i���0�lG}�swk��z�5E�vH{E��N�|��5{tK����թRu1�Uy�\�����M���ag����/�W6L�/�O:�ޞ1�=��G��^Ў�Y�:���g��'�Ʃ�D����m�Ċ�{�/�ۆ���;2���.j�����N-��ܬ�m��;	�x30U�qY}t�t�::��5�mvw��wЖ�*R�n*��JY*����j�7:�,fؽ渡:�-S�hg��ڗP�U�U-�J�NMM�ҭ��5���k�0��W�ls��Y\N,���tY�a��6���k�1���ڽ8�R�t\�w\�{3�u�[+�A��)�S�z#f�t���|�s��@Ӵ��qe�G��6�2�5����B���N٦�oE\F��l���4��foMa-T��Z16l�8�-.Hyy�����1���=s��0��J�2cb����6�@6����j�������1�Ӷm�;T�ǀ�,�~��]+w�ޞ�����ї�z!�o4=|�u�>�ǺU;��=�c�s�Lm�Ew+z#�Z��x8z��2�_j�6���땋>r�	oY7�˔�\����+I�7$	6��r`�pu�e�l}[��`��4�����>���w�� �rcp��R��'�k��6�3;�keH��G�v�B���^��p�l�L��"���|��W��ahO��5��7}�f�^����'ኂ��Wb5䇛f�+��)��o3�;���������U���!��.��H��R8�_S�0�J�/:�<�m=40b���v4�+�����J���+�lЍ2�;�d��6(��5���#��WdAU"��ޞ���Dd�#��m���Jp/�.�!�N���x����'�_�C�뉎Ҳ��,��\Yd���Ό����E�͞�3�n�
X�{����u��j<�gt?B��Kh���]�9��_y�v�u��4n#m�u{N�Wz�Yl8�Hz~B's�)d߱�vS�L��ӣ��lh����6j����yv��&k�ǫ����U�1)9g���ɨ�Ap:��t[�@�ldΠ�U.��u�;�(ʝ�<]�x��Z�Y�:S'���[[�1�ޒ�,�H��+:<Gm��ޝ|�}BK��q��f抇;׷s�e��!�Nv��aA�=µ[O9"VL�5�ײ��\�cwv�l�w2I&�xz��6������}?���^�񝕖)�8�/slŇq
�j�m��>����E�#r��y�s+q�=�ZX:��YY�{�[�^��2r�c�eU�`ܥ�Wq6�!-b������]o.�ڙ�`��HB��Q�˼5ÑY@Z�Rov��3v�^�W���N=�>ч�~���+�;Q�d�~�'��coC���1a��-��L�e�{L8���0p����Lıh~j��WB���49�p3ln�y6܇�Ǵz'�t��־�&�W��͔���ݧ7�)����I/�o�=�z	��?K��m�]�0��ّ�Ɯ��?@��nb�H�������;ɺ���Ð�*�.�Q"N��/�}����P�����Bw"�H�3<�y���L�~P|l�N^y�b�H0�}F�]-��k]oj�lݕK��[.m��Nzj���ǒ��x�\��
M�4�r�w�'
�fۤr��s�)2��r�n�zk��KSA����/.LӜoxYZ�I�����>Gc��p�ބ�˹���왹t�dU��R�c��n)&K ����G��C����Y��t諚���6������Sن?�Q��tk�\�xM�s�jf�����5h:�#˓��M�s��0�ݍA���0�� �z [+j�d����:�x˅�ʷ)�ȷx$a�8��YL] ��}���=�	I�ו噒��m�/7Z�Wi���M����Y��*�O6��d_벚�#,a*�U��_*��M�+�����ݧ�����q���T��h]>���4����iq�^{%fZp'_MngN�Ol�"/K�$��C�Q��϶�C�͟[���1;�caZ��
��[^Wܻ�?����g�`\�����ܮ�/�ٽF����j2��m�M\t�Y�F0Nb��c����m��l3����	U�PX\9�m�g̸���=���\�gZ�r��#7��֟1���[=f���5P�ɚ��w�7]-t"�F��{�d��M�=:w�MLd���	��L v�1�l˸k6��P���gV�_F!�:�p�K�G��:�n���� �7��NcO��A)�RW[|��"��]D�õr=w��R�ޥ��]r�՛';�f�Д	JE�C���H���u��	��[H�3�ѱ�[4����G�x[�-3]��M�';s�����kg�q���#^��B���R��鳭7ѕ�XXr9�6E�xC���U�.�"�����_��� ��kg��|����℃�I��n�m�{�bSf�뻇����
-Q�������t��$��%�Ϩ����s��x��F+�o��pI�Wn�2�G����ZAyQ�VNu�2�� OC��p�O2�@��A�9����M����Α�;�]�=�iVy%j��CY��Sb����7<6�U�m����xC+2hʲ��Hޔ��4�[Mo/�:����r!s*ʸ��wq�K6l�T0EF�8(u�j]<�yZT�|�������������-����i��Y�j~$V��v�� |��������}>�O����/7��u�L��ᆼ�֡����R�+/)�fN$r�4gq�O�%�1JG�օ�ݹ	0��I��/���1�VoS�l^h^(��7vt�m�<rkq�.+�ON6����,�&�1�r]� �r]�E�_q��Eu�qÅ7x��
���{����3��[8�vN�~����jj�Y��J-3*��gSj^lt�v�=AV@�g%i�;.���a�Z����Ox�&�gY�K��A��1h�Պ��W��Zz�B�n���X�i.�ݻZ�̸�j�q�5�9�fcpuc��9Mȱ&T3~��ɱ�����r�\q�S��4��w�t����è�Ue��ɽ|��Nk�bf*�K�b�,�8�"�m�v��n��.�I8�y���ݱ�k��L���;fSV�E��S��9Y����A�oV�\WH,���]v�Y�z��l@��M����.��y�K>�v<�G�*#��Z�H5�)3ǜS��)���0T��vܺH��7G��_
�'�]�<馎q����/-��
8�JB�{��t���d�!7�;2���Xu�8^|�6�ڵ�׵yzH�/<�od'S�V�tr�e��]�ץ����Eƫcb�0Y�Li�ԨvG8�wϕ���@�	[*R(�'-�#`<۱�w�����F>�:���yL`x�"#�NQA)�f$�:��ei�.S5ͬδ�㽻���]�npd�sl*Y'J��׮r���I�-Gç�����`d^���`�)l�s�Z�ﲅtU�͵3G6�=2�G-cn��y>�.�/-������[��L�4v3���a��w�X|A]�4f�VWm|��sm���'v�K���h�e#Nq|Nu��oV�/W���]!f�1ëqI�,���8y����ԗv�g,���=�� ��z�5�G�fn�5ayQ�q�Uc��q��ۖ�6i�F�6R�C0R\�9�n2���]�%�VrB��B'*�Rv�y�A �6��5[ժ�w}+��E��N��Ō��N�X��tPN�Kȯ��̜uvnjYK-�8�N��n�m����>n$����ۖjZ���N�m��vH�X�AΞ���S�w�o/��V����`Y�W�
ޭ�z��L��)�Us��X�*��(#�S�E�K ��Gm��O��K�D]A�~�U\��b�2:t��C�f�}�Z���1�(e�0�2,\Vޙg�����٪�tw5�L�4f�2Lo��<�p$�١w�8E�4�2=N�b�ڱy��XA�4d�;�Y��8Ʊ�Q��f�vf��M�ݑѨ������-�܂+���J��)w[u����~���Z�F�Q�A���*U��n�����b7\�Θ�'6��J��I|7N�:db���@�YCEwL��6�g��gu��\uŹ�+%h�E�؟>љmW;3�nA�F���V W���%�3���B�:[M�a�"�����;L���D�EB�T�AP'P٧M0�L���A��ֵ���4ih��(*$�T��CA�5��(����:4TB�PR���&�`ב�15u�)�QPDã]'KB�D5vJi4S�C�OZ*��4�$ON��(ۻIGV�v�<HQAMD'lR�u�3��;n��Mi���*�;b������+Z����d����Jh�t�y�-iאi�4����]%4�F|�
bh�!��R3�P�AETu���
�STh�RU	E)�y˯)�-۠�$���:�#�	E� 4�yhnƩ�MR�HPMHyh
J�t�)I2u���v��C���i՝!��(���:Z�����*)j�
���P����܎�������n��tot�w"��"���c�� [��)f���ty僘V@K�-��[�1*�Q�4C.T�ɝ{ǅ�7�on	���^s�� $��s>n��{2!ֿ�W�#O��e7�66�<����ԅ����q�������2�V��&�������������x�H�KuX]�A�V�(^G�6��j���e����t��,$�����޻⮎1޴� ; -��Ћf��lw{+oV����Ulրǌ�:�ܨ�~Y�	����"�!h��4��{��Ha�}��� (�n�lE��e�j��kY�w�rw)��O��Y���h���ȶ�9@���:\`M���Ȫ��m�Xv���@N��wu���%����w��T�ƙN�8G�9����]�C����*|�S����p3��a����h	p:B��T���Zӱ{�����LK�����gի�w�"n��Z����#i=@�L���_c��\#���s/��RPۻ�.�ʙo,KOc}�����/jι�)�"�岥�2��<��/P�*s�
P�vwaS��x�♵���ί����f�d���yY43�tmkleH0�hZKV��r�����o+:����v��i��ܤ�~��/�Cҫ��W5��ns�����y�-Z�fڧ�ѽ��L&�:������M�!��Un��� �[��,��,nY-[rZ�K�~�"ʬ�Y�@W�n��[�6:�b�8��>wK�E��=)����g��;���@q:j�\�v��9��l�S\�v[��ݚ7w��!nf��D'����%I�ⴲ�\�lPgY�s�� �[4v�<�{��Zg�����S����V�a�и�Er~�=H9�k@��u/S�3R�M^�����"'-C�"���8=�LH鼒]Ǐ��Z�-�o<�1K�q��d4
j�fM~pF(7��1��5^�Em�E�DDc?X�i4��$6�k����_ex�F5w����C%����P��VJm��m�͞9�=���h�+*m8�ygdMѾ�r�ǰ�l�����.Ӂ�D^��f0a���òv�x�g��-u)37C�l<�۝K��3eЇD(�ҹ������x��_ On�a���<5�N��+hΜ;v�C��㤢F>���i�'Z�iG�4箱*vk�X�"�6�Nmm�*rd�y��,"#8��[���QM�C�B|�oM:�3��\�)������v��2�c>�c�OP�-�=-8z���56\k�08Уb�j��Ŷ����p9I�U6�z��B��B�e6�ow>Ѷ��q�E��}��0.�n�nI��P��#u�f�9�d�{Y�IM�>x�jʘ�멓s�E��_�Ճb�tƉڹ��@��d'�Xٲ\R�=n9H���~��V�@���FŶKUpy������NP՝T������]����+��E��Bܶݳ��$�z���Է�VD�-fJWuVmԁx˅ݍ���N%�b�jC+I��/�0�"o�����G,qK��W�wQ�j}�B-��t]0O{uf�f8�n��A;7��s��1���3A+d+9��G\r���>�>]�E4�G⩀�������.�3y*�*��N���'Ȟ�w��v�D�A]夌�ڧF� �یLB��v�AD�VhL�|�]]3'M�)��eŜ�@7-�wYfh�j�J�ǥb�wî��C3��[����1J4��9�2��ܐA���ݺjވ2�,�`QS1v�Y4�PS.�V�o/�L��9Ǔ�v�����{CQ�	}��~�<��O3S��Ağ�O*ě���ty��V�I"���{Y�X��za�<O-��~�@꜓ݐ�V�O{�$�\��1"�7I;�/�����|��He�j�z�u�.&/[0�^tq���?�q�TW5���rw�A�W��ǟrDcˀ���r�qK���&Ty��*~�ӓ�}�o��cQ��3'�6ڷ9`��D�޾Le�n�l��>�HX�d���;`l�'H04��*�^n�h�,F�'x���}>u�����"3�t�����g�_cmP[��i����U����M`�+0�O��zD�D٪�㚪mC�j���F[q�/�]�yq��F�&�kR��d(��ܰS�w���F�Y2�{=�������-��Z$�rR��[f���<LI�i���y4ףKL����cV>}�F�Kq����]i^�C<n���O�*���!ntE��K�x�:��{��*��U��A6�>���-=m�&�ػպ��Y�u/�2R��}n��+���`�9H1,���[��(��/�����q��݀d�ݴ�=�b�$�ő������f���Q�[zz.5N�YC����ǎ����B�g��"9�j��f����m���ʮ_5�B�+Zp�;^ޔ��Y�����莖���f�'��Z����\��z���"l3�����w@ĺ���a�vҁ�r�5E��hU>�����k��m٧�QPM;A�u��+����P��jQ9�v���^�Hbx�/=��]�G�M���t����d
v�G
��Cbu0���o^�g����R78��+��>��J�$w�d2�#2�o.k�1�g��}�t�F�So�}��'ռ���U׊2�Z�ľ�蜳g��6��"��f������{��J��v�
i�gI�h�dk]\w/��������u��(ϣ���)};#��]wmnP����,Eq�z"�h�n�S�6/P��1�i���W�43���Pze�b��^ E��W�L&��@�)�+5�Y��V#��n�OF��=u*k�ai�*brU�5n`�8�s�Y��ʀ�pTn8��!��L2��ؖw|h|��J�ƺ!I���=�p�]��$�-�rlEwM��|��d�qFd�p�>������};K��s���8��G"�Dk��^��U�[m��L2ȣ�}�F�r�D���*Ա�R:9P8np�U�o��9���f����>���hǯ2b@��ґ:B�[4i�C*$u�h��ч;��-�Q�TNM�ݣa?Wq

���1���s�l݂�x�g�G,���#��W�t&��R�jW@^�U,�;ܶl��.;�k�zIɜ���=o=dgd�ܶx�ǅ݁���!��jY�w!^d�44���F���W\����F0��N��Y^K2��ɠ�<8�t��~A�XU%x��	Wn����t;�ܤ���P%+�w��`7kWMn̘ny
���q�s6��x��-{�|�xBQ�r�-
�+!W^P��;�G��q������Oݏ���%t��WO����o����t.=��ݷ�#�z�/-��g���I9YuW���T�l���#y�����%�H�#x$i�J829/Ws_\=i+�ç�{�:}� X;w��G���;��(V�3�,��r��EY|(nk^ˈJ��n��-�@j��=s�oz��d�,D1���yU�io{fwD
%��os�.ɺj[O������J��&nԷI~��v��u����g�@���T}��L�`���oH���}��wȬ�ҫ*�E�w{8�.�4�lh=�_��-�;��00m�t�Kb^W� ͓���t-әZ�޽��m�W>����l�L:Q`Ô�Ǝ-"�vSU����	�������m���T��Nv��Md���O���4e�2/��a2'%04f�w�^V����8��P���>�:�^/|��l@�m�V���:�]����[y�S���[1�A�>��5������#����9x32��)biɸA�A�Ms��<���=O�H������^k;��{aF�����P�&�g����i�wc4M���r<�T��2#���FK"�<��W5��_at^�㣞A���77��ztb�x-�%��ȷGKT�^�0�x<0˨���m+����e�h*k�Y{sA�P�j��1nZ���/�q7�WP�U�/��dR|{����9;#}5���]c��r�]���f�U�˞��e`�Jx�5�Fx�n����SӠ��pg'/��),2t�/e�o�U�ԗX[+m]�WuBͺ�p
����"h���Ŵj�L�AV��o�79��G/�\lb��+��E�\(��8��^+6n.��ms������f�'c�C��-><��0�(9�I\��v���0.6Q�ȼ����U�=S��0���p]!�)��h��H��\c&��*{����w�3��ue��K�7f�:��6�F yCce�*d���hcNov�ek�u��)�5�G�͇8��y�ڶ�V!밝V*�o`��]�|u�g"����,c$�ڿ`b�#�t�`�y���)@A�74³��y�6���Di����;�-(�r�����pI�HDH�7�q�U����:��#�C�������d�~���p�'X�T���
��ϕ��h�I-��O&�^q��Jl�Vp׫y�Ο1�b�d�R���������+��1��SB�0M�,�G���*n�[Z�M���M�w+*W=<�yL[��4�#�f��L>N��V:T�O�a�T�wҦ7Rry� i�v�;���*������b�Q]�8���k�B*g4�<�Oj�6�:�K��m��B`�:�j�ʣ�0T�����ؼ��vXH����P�k����^��)������h�� ����A2���R:`3�5wL"�&ͺ�|�nut�ƾ�(G=&b}���	!�9
�T�����Y�(�W=^d�n����������+��D��Uv���g����]m����U�4
���ǾR|�z뉁q�w�e����	p1:Wrّn���M������G�T]��5�(��}��^�Kt�,��{u�A��ܠ��Bgc�m��dNj��� Q�h6.v��n��1����������t���M�U\�u�P50�<�4y�,�Z��î�~�)�Ǚ>V�ۯ�i��:�<3vof�E, ��M��%̷W���r��q�9�=���ًwK�TT�����(8Z���t���O���>�2�L~sWW���Q��6���6NcR����ʳc�2�=�I�ҮKUpp��Ux]a��6q;��۟qr����C�}�Vg!7yt!�{
���R�K���`�8�v��m���1[��q<��Ǌ��1ޤ�ꝥ�Z��;^K�Y���Sl��]8�R���sHC���t|����;s�cv��^3��ډĈ��}��YX�S���m���jO��y9~k����Ŵz�Ͱ-3����F#l�*�Ɲ��س��U�[�J��4g/��.�v����u0��Pj,�ŕv�z�Z7�K�DjKP�γ����5�r�=m t�1�����B������F�b�����w}Rl��G��8��(aT��i��bg����'�Z�Ҧ6D�fCw9��z�h��LH��ґ#HW>*١d�3g^A���5�F�7{v�� 6W݂.�E+�:�f���0ܹ�#�n2��K�{z��7V��g�k6���z��d��e�ne�*.�R7��Z)qvv� �u��rIeP�j��T��4�Z�����W������z�>�O��������������ߒF�De(��^h+Y��+8�3�9}�c�I�\k�����X�r�3o�nM���5�:�03a�s㓾����ȵc��P�4KwR���*����l�E��π�
�pHxoYT`�kv��7y5�ٍ^����$o��Tw|��Ao��jħ�o����Pw�����Lgr�S�]X���a�G'V=y�%�\�t[�â����+�{\�����-J��Z�c;�KŢ�X! 4�����7�@o5�E�]r��.��j����^����w�Q��«S`�t�]��vL�i�faw�ӯ`������9^#�jB�`����#��;U��fڙF�7�{EӉ�����]�{>��:�ޭyRV<4���3��u 8b�ofs)��ɾ}̰z]�#yK�:���4w�eq�畧]�"F]%���lIM�6s!_)v�<B��ɼ��q
�z��y�O��" ����<�1QT��{�wq�:8���Ѽ�CZpJ���Gwm�w&ofCC���tu�
�M��[� ��{`���p��y@�?.Y�G������X^�B,9}s�*�f	st�3(��Лfڏ�s}�2Q��Ѿ��r�&1b��Ą��.�H��ٕ%]M�^hᔌ�Q�Gv�����bh-�p�^��T죷p�NtT�� �2u�G/(ӌ���<��!m�&��Y �Gf�\����6m��9ʹu����e�oA;i�qE��s�w.Ӭw��
��\VU�Bj�#WS�ÌN#㝱�]��#u{O�_M6�P�5t�`b�����=�`�����B�$J�7uGM�0�{zS��B��.�E�Sxg,�ݻ��`��W%����y��c*���L�s�������K/*
�T��]�zy�ە692���a�պ����库�����|aXb�l���EY"�=c/��C�OM�wΛV&!��b����I��c�`^!i��_QN�ȳ�>�=�-_5��:Q���i����;+sSS�B�4�#7-�:9§+U��R���A�Ѥ�kNqC29+[Y�)�.�8�S��/��'$1�'Mw[��6�"jlA�8-r�Dz�Z�Ekv�D� �;a�9
�NU��`_з	YЍe�ƴ tfm��7��]�Q�\��Rǚ�l �:[.a�\,q|������v���J�O5�حL�y'Mh3	s��\9AF��E�'A�[�E*�鲺5H]uYx:D��y��8���6ws��|(�G�}i��*��hΚ��rs����`�]8b1a[��
�aq�1e�#�1�2���w�� ȱ�׷J�I�M�1B7�TK��҆7��1��,��. ��V��w0P���-��\�5يZt����6+�|�����f2t97���=�m�]ҡK�Pl�3�l�flC�������;u������9�/PX(;��y�����J&Z(�N�4`J/��F&�J��vB.���J��5u��,ILM5�lW���T���F�1����ԴD�4� ]�A7�B�yE�F������B����B�d���th)�i��"�N�B��<��@gO�a�
iO!5BR�:�/-�d�j����e7`�hN��Kl��t𞎪�Y��/�OLGC��1R�P�4S�BU-�:N���֗N��w�N�HPv�Ay�CHQH�ͺZ6�1)ւ�5��j�%�:_%5K�i#�4��B�Uu������"-=!N���&�CѠ�(J�
���x�:O���yY�\� e��S�yl�����ͩ����+*���קn�Pː������s���-ƱS��Wm�T�mm.�*���O{�����s锫d��x�[-�1q���
m���]]V]?vg-,�&ċ��K�I��9i,��n�X�E[vd5١6p� �Uo�����70	z,-�|�o�Թx���G��^�YUוJ2�p�`a~�b��\��쫔�bO�����vj��[��o*�ܼE��4K����Y��޵��1;<V�\0W��V��'3)*�v�n�}��ͷ�խp��4�z�;
-	l����;����8'��M��yW�c=�ӻZ$�|������s��{��c~�r�g�n.�XT�B�� ��B������_����uW@Z�y�'�z|����)�[�q�I=����O��� U���zA:޿vC@��k��xz��GQ·1~��Q��lW�q�Jxkd@=�~�he����H�b4P�΃2Ъ+]�Ӌ�캾�}4�2��{�1��Q�w�2e�Hm�+o+ƺ�**G���P�ѷze0 �1�hu+q-�����,��wi��y}���P�xvgt���ʛ���DŲ��2��n���=u��	��׸s��V�3�*����
�ܮ�������K��_�R���Vr��wxa���	�+���ײ�M=��Y����i.���]A�Qٿ� ��o�_���&����nv�~��3���}V+_��\��j�h�G�5��s��)��O1�WM�;���f�L�|�����~^�vo�{��6��,w���j��r��zn�aၤJT3z5�Ӹ�f����l�n:�RJ��V׬�{+�fU�n�۸�n�0��[HyxL���*@�bAm��C&�q��׮:cƽΎW��Ю�L�����y8����$��n3Sd�+dY6����F�:R9I����ͽC��][#�^�J����q���_�VLp]6�e�7��w�+�w�M����U�~�f�[[/�q)ѯW��e��XY,����-�k�G3W�f�f��c&i�j9���y�:�"WXu݊�s������̍����M��T���=95��ǶY�N_-��i�6d.(A�wv����З�m7
�'�w"��Pjns�1���{D�#79�s�t=�.u�r�����WZnkNM=��=�r�������)K��Y@�&�״@J����m�:��ڻ�DY��m�.�hy��?tª�)D��2	�XQ��Su��m	S;0:�Fߍ����0���� �|���b���ki����Y���U(�5��c*��_Fd�a���U�}���=��#{hܔf^�LeSX���y��d6��Hq���f�"��ճ��z`�4���\��S���]��:-��+�D��,����E��*E�d7��o�+�c��hG����|�r:4 �L������ 5wH�hQS\�C�K4�z'c2t:�sd��x�D��f�Mj@v퐣��ڇ�.�u����u51x)Y��17�dƬO��N��vK%qkh��`5�l��{%F�\��o��R�T��&�jW*7՗���Z�)<s�qn���v�I��g'o�8��z��g��mU�\���!'��?A�����?oem����ϫ����0�VB��2�N�V����6�\���;-4���k)��ز��
s�?_���9/Wc���ݡ@��Pd>M�os&)W'w�(lv�w�r���2�9ʎ�:Hm��C9k7��V�����\ti��aJ^	��Z���y��%&�s˼�~��ɲnԂ���g��?%�3���P�E�^�D��s����%�XҜZ㔫$+����Sl��h~ٰGS�����ɬ�ٰ�v� Rv��9q�^{��d�uzs-���fX^��
��Y�t�jG�9*��59�QS�-��s���(zv"�W��om4ƴ��8���T;�l�>>R��Z�K3��#-��Iﻻ3�9ôq�B�cX��b�O�g�W�z;'M߹+�Q�9�W�O]\��0�u�z�(�襤[@�f��@m�	G@�P�s'�׬�� �i;[G��<�b0���>�<�|�3=��;+溓7�����Z�szOL��z�:���u|�$˚3�!��6s�4�u�N�k��pʵ�H7��w�d2���v��<�r��`�,eX�y��:%�E:��)�nL��ф^d�i=â��Uq<�3b8�/��5�EA�r�ُ�tJ�"�P���M2�����i�y���Ь���y|vr��g&��kz��[[�����r_��<�
�E�h�{�e���X���S��8�CT���߮��{����D_��B\.{K�Y
���L�A��)ݖ�fh�6�y)M�f&��v+�]c[>	�|Y��5z���QV8Ʋz���*ޖ: ?G^��|㥾`�Ա��c�4R�s�I~��۲j&Ƥ���Emm��WL��w 1�n����;�i!��ձ���#��N0f׬nz�7I�9'*ʬ��eO���e6�K5�w����}7��Nq�}@��2���&��[e����W��.��Bݧ�v'3*�=u���\st�K%�|6�V�-�)$���J���ջ����e��G�ϱ/�7���#��7P�����g��q�]T��i9�N����DF4�J=�.�Dx6NKvt��K��㣯�W�	��z�1ۊ�Y{6m�r�Y�OX�Q�Bs�ی���l�������|%ok��%x��8;Q��9W�b��9'V3����Ë�r;�3?O	Ԏy�`����}!k�������a��q{u�ɯ�����n��[��%��Us�9��#�Υ\�ZB�wE�`� �Af�ڒ�j�չ��9Sك��DN7E\[ԡǏ�x����v�$�i�-�A���]�\6u�*�{9e��
*P�ޭ�&v��q�k�'�gdM�;�a���Y��S��%lY�S�`kn��] 5�e4�i�3FX�m,���>�kʭ;�h��ٹEĿ����fD1B�.�@�E��r��7��h�w�[:��OE�F`��᥅"����f���%�a��%
u^���7��{v��c:�T������^~�
՟)=ֹ�{[D�A�q'3�����M���TV��F�CYc��|�j��v)OL8���U��he�BZ{��q	�_d�su�V,w���i�����a=�k�հ�R*��ӧ�el�Җ��z�d��ꅛt�R�aP�Kݵ��iƫj����[g��8�Zh?Cx���Ҏ_����V`��<�$��X{f�65�ʳ�g�5f(O�!�A���6�5��e3�'�*���neԋ�bw�*�\G�"����cV0YV�5�� ¾J��A(��3���X,HY�-�ֲ��M�}耘�^e*V��Ɔ����'mPh��4�ʬǄ��E�Ys��;�s�.bvw�&W�ռ������w6L%�E�����xDR���34�`g�n��؋-Ww�����&���?�'�w��CJ+��t�[\E8��X����k��&�.R�W����̸e�j]i22<��j�}��{�,��iGۘ������9fy�Ku*fv��N�[?���n�M��C19k�Ά;�w����vRyV�<{uaG�	m�_؊I���KotoV�nI֎�4 �T���a��b�nZ*<�Bײbo{��[a��o`mK��I{:\2M�H���� >�i��#@�%�y����	~�ݟ�b͑zIomz%2C�αۂ-�_�Q�׫mJdwq��Q��r�����i��o7��=bAV���5��E�h����쥖�4ԙ��5�>Mf�kt�ĕ��7J^���de��0��P���7\�Qw�W��U[e0�cO8�G!ˊ����L�<��h��ӊC��s���+dv@�\��Q�d��Ȋ	oJ��ܶ���5���^�I����0��x�'��ݘ��\D<B���B�Y��փ��_NOQȬ����Y|C�h��� Gr|5d/DO�;W��wU���ČČ$�h�+�Q�e;-�m�\v��R=��ݶj-�j�Ë�.��Q\�ZBy�h�����U��D~��{.nn��v�ݩ��q�(2R�/�P̹�1��r
U�d��욬�͊��Ή�x.�UT,��[q�&[f��p�b���6{�!�ޕ��}�������������P*�/N3dj�Kf�j,�w3V����p]pw�7;H�U�Kz�+�YI���S˲�WG�	�4X��'&\Ufl��<ӑm�3�'�Q�1[F�������^�#[�:�n��]�(���9I����WW�ɀܥ~3�e'����$}�U�vѹ~�YT��Ԉ�Lj%U.�ٞ�4� v3�Ѯ� ߷�G���-vMqN����g����p��fp��v�ĐtKp�	����F�Bgcѳ�}�Z���]�3<A�`�N�����S:套�s��L`n[�א���S�	ce[�����M���ӝ��4B� �9п���w+����ρ˭[Va�ڵ�|r���g��4�Z�����3aZ��f�����l#j���Q��Z��y���j�������c�kH�U���4?�.w���uѝ�<�M;m�>��88�f"�`����Ec ��z�8ȣ�쉑�z9�꣘NL+�ϧ�{�~-��K��l�����9��.k�yga���h�%�Tۻ��Y���rq��,&���n8��t�# U)�2�۹ͦ1��]9��������{t#7n��ޖ�Ãt���B��wm��<^e�v��pȖe�4�#l<dx5*��S��po�%"��Q1�1<dY����_3%�wVX�銫v[����;�!*~6�U8���6����w�nw3�:4:�{�<tr��v�W>�q��v��
�a���,<;҆|�ԦK�;�l7�b��O]�[>�Ue�3�~+/t�튚ފ��x|�q:ɺv�� �G�C�V��$�"��<o&�ƩeNl!�e�N��u��ش��	S(�8\=�'Í�7�jL��8�|��4r�#�|�Dyk4A���>��)�_���aݐ�!�}y-uG7%l�Y�Č�І��}&��e�ܝE,�-��x�*`[Q�Y�AmP|	���]G�ZB�Y���k&�^5+w����h�O�qt��J�y7��r�m���S���ay��q��Q ������#M���|m}��p���6`7=�%�{���ꍯ���k���ǭ���������V�:ށq���V]Q\�3r�c2M�}��#d�'w��B�B['k����mE�o;�N��W�lt���{�S%n�`*̺��qm��7g�|6�c��3��i��hu��my���Yer���D�&����z.�4i����+'����,(�q�i�OAs6z�n��MV*��;�ջ�d�����xV�3I
#�}�B��G��M��^��2�_Pˡ,��+��F�g9q1��U�_S�����7����U�]�r=y��:����퉩�Ptd��}-Q�����\b*�����������U��#��@]��������q�L�#������#��?'o�Pp2�0,2,0,0��� L�!̫02��(C(C �C(���8e a eUa�U� ���~~( C |a����� v�@:� ��@��e a t�PPDDD  � �Q � @�D�@�D@�T � �� �� ª� C  C  C C*���2��Ȁ0��� � ª�*�� ��"�*���ʰ�0,0,0�� �aX`XVVV� !�a�a�a�a�a�a�a������}}A������4
 *L"
L����_������_����?��y���0��������p�A�������|�>}�_� *�`g��?�A��� �
������@�؟��i�`��C�@ ����~���7�H�/�O��o�����x�?�?�E�ߵ� ����$,� � �  D�H @�J � � $ !  B� � � ��0���+  J��H\�*�H �*�0�
��c��b��?���������H�P4+B ��?`o��?��?@�������>����@^����'���'�x��x��c���<?���@_���J^���"�
�� U��?k���*�"���{�!PW����L���ྸ0`�ho��O�x��_��@[�C��g�B ��C�(�������i�Cϧ��?��$������ ������W�����I����L~�,I��?����������}~τW�>b�����L����?����/��~�� ������x
 ���?�?���_�2��b��L��/�3�gų � ���fO� ā�����QU"�RE@���)E)$�JHQ!P�*��J@%*()DQ"��)PUH��UQB���I"�AP��@���T� ��BT�T�*�ER�IB!)U*D%EDT���T�*UTR(RI%R��IJ�u	JJR���UUU
��%**��BQUJ�*�D*�R"RRR�H�$�*��RH$�	RJ�D���TU(��  c�mF�akX�P�Pk1e �4�L�Jl�6�!4jj�P�e�XV�Y�����j5�ZU�J�S*��m�Sj
AH!R�THT�IW  �
(P�
7(�4:(P�B�paС��
 P�UaC�B�
�UrʹР�T�մ�	M2����Z����i5Mj �kiY+iJ����(R�%��DN  6��H*��ɍR�+M`Z��mJD�
����4�*�*m�Cl���1�m����im�)F��j��[bm-Lha�-�5�)UUEQ%\  1�[f���6��-��*���*3(�j���5Y*��� mj���@6ְR����(R�� �T%TI � �"�  ut�ֆ�`�i����()�Y�@!�L���m@�4�����ٍ4j�iY�
H ��RR!(�	
P8  �B� ��T�@�f U�IX�j�A�5XP� ��k1U�ژj�aJ��EP*D�"��  	� h+V5  fҢ�j ���h�4�0R�2��jр4 6��)�	��hM�DD����R�\   �  �6�@ ְP m6��,V� @�P �ʘР�6�� �5`  �� h&����P����  1�  .E�	�@6j�  ZX ��  1��44 )�  m�X
 
m  �(�B!R��P�  �@tV Cd`  )�h &� �6R�  
 �X F`  Y   E=�b��A�� Oh�JJ�L����a4��M0O��D�  Sɔ�@d  	4�i6UH� ����8�Ȏp��2�ɘQ]IБƞ�3�n��m<�ӎf��ɿ�!$I=�����IM�$$���r@����$�	'���$��������O⡫.]�?��泉������@�[�죯2�&�
���i�r#z�6�5{3Sێ��um�.�J`��ཨ��kH !�e��%�w���Hn�7�ՉH�-�3u���e���ڱ#kq�� ��ō�Lb�f����,yE�-�͊��LgZ�e�:63f�`�@��z5�L_���|���cC�٘5iꗑL���F�յ�m���^cWP�����&�3+u��hK�2��P��m��HkUf�z�ʄy��N�dt�[n[�ZP�"�Y��C6Z�#��0�r��OU̰f���Rs;��3M=��z��A�0�df�Y��g[t���h�z�
��Z΀nŽ���Q�k�teaA��F^��+��^ͻ`Z
�dѮ�f1QE�Y��U�P�bH!z��K�j`I�IJ3S�,��Yx����z*X��S	w25AUz�͕Oh�9��n'�hТ����d.�`�5H�B�f�r�"I��.��r���`�u�ie�P@q��Zn7���]��^0�S�ޔ�G#�T�(��ځ쁣����im��t�ֹ����BX2]ЖJ��+)^�H0���3GY�f��µD��oVҭq��*h�;�5�v=shT��4�*�ǁ�Z�eR1L����A�V��k$��	z��MA!�0����s`�U��T�9�K6A�a�Tɀa�7h6�K]ͬ�f��ǴlH���Tx�ژ W��n����2��(!�T5SYj���qPt1�ͭ+N]@"ո�IV��bΦw�޻4��Mf��a�m���f�b� 4����sD����],�a��sl����&�َdT�!<jYy�������t47���[Z�
�'N޼k7hc�2�;l��wW�j�,4����!+��@֙���i,J]電R�JR�
8h�(]�Z5���Z��˺�c�K��򍹘����p%��f̩�O�u��t���ʚ�(6�`�%bu�[�)��f�&�A�j���Yuu�1���4�6���Xܬ�BTD^j�PijA�\ۘ���v�>�iy���r�y������e����p�0K$�캁^��	E������*�`ku�U��$�b�c9O[Q��ͫ��T�:���l���6��2!�1�z��L��^)H�����e;kO��2����;߭�Z�3-�ୡ���%z͇����d�{{����N�����Vof��!p���XӑL����*yY!��e�4nT���F�۠UiE�;>�
�9��ˊ��Y�J�V�ݸ1s\�MelRi���JY��6�U*�.��v�(k%��	b�����,G)���r9V�^�5�U1�TUv;�YN�f�4�Ʀ�8,����nPh��u�v(�!��{��ۈT�$����--��%��l�ٴXb�R�l�A25y�����X%��B��J�kF#��jZr�{Oc�������X��\ZƸf�J=@���K,�Eہ����D������1Gm�c���*E�`���f\/��ݨOnd��:�U��E�"�X�L��s��GI��a��]+�	���^�?��f��3o�	d�f���C.�L�ʷ�-_1YX�A�E����j½�v^�3YBS�q�t3 ��j�1�<�Pe�i,�B���nZ� �3H��L�m�[��t�Q"�8��$�vR�m�Y�5)hZ�J��i�ͤ1�
Gréws�>Y����l��nJr���E2%
˖�lCM�u�]9����*�JS��q�*�e�eV�Z���6�hm3���N�&��@��ܻ
�Tm�����2�jfQ7�,`aM+�U���q �#[�Px*�.JR]f���ڼ�V�h=P]��4���aB�i�Z�^�oc�.��E�ښf�Մ372��b��nY�VjU&꧚U �e����$��������ɦv�޶	Z[�`Ke���uq�3E&��
1]e�7m��J����F�n\�j��"�v3^
uP�,f��M:��0��������,t��&��ܿ�$v-�x�PS��n���Wq�@^1n�j��um`%Xٖ�I ��Kb���a�����S�S���4*�`+ղoۢ q�����ČjݘDI�-"0YQ</&X�2���̲҈J�V��乲�6�h�v��&�̳W��-��:�*�a�ۦR��!��V#�t��I��hXp�-��r����y� iM�0^ӡa�);�v���5�B�^]�l�܋UИB@�譧�Fy��^� "�.�Y���)"��S�-�3&�Bƃ��#�f`�$VeH����^�u���%7�èږ1��ضڨ���;�1֤K�C2�Xi�,�0[��%thٕ�)���v�ذ[f��"��Y@���p
�[��ͳ�;��HJ�/Įի�����x�*(@�J��
��A2��u�CZ&�ǔ��K2�j4.lz%b�	����
��#+-*�3TG]b�t���L��]�(�טח�u���S(k��qa`eLiY�p�m^)U��*���I]���,�n)�6\�23kK��à�-C6�|�ne�Z�1��Z�l����mbF�̼.�+Wc�n�@Ї,R��1�h�B
4�7gtn,����bG`xcGt*)������$��T�JN&� W�fc9�
�E�WY+*ӥX��k��
KgJ��e� h� ����r���koqހNc`V-R�n�c��4�i�`b�fj��	�zEV���{��cn�t�b8pkkv����՛Q*e���մ2�÷!����"5`�TD�fD�`;k�B�
9q�F�����2W�5��2I��T9v2�j��7MnQ��%҄��ݜ��-��Z.��KM�D�Ў��,��(i����L���Wn���l��t�\݅=*:'"&��5&�1l���dۚ]6�YF�I�q�d���re[����b[�A;��5b�ZV[�KpT��k��N�Nn6��y��5�XہJf�ꢮ­�唃���P
5��+Š���)E(TH�N�V2��8���Q�3.���u��)�oT�5�y�7v���!vB��`�7Pb�vT5tvȆP��V9�c����RJ�L07r*��.�����g�ͤ�r�ݐI�e��w#[�;pMP��1K*|uꛔ�X��-oe���i�i�ǴA�z�	1mͬ�#�E[��N��+n�D�k*RSz	5Gr���64��.�m;t��nC ��m���Rܘu�+2f\�TR����[��CZ�:�������E��S�t�S�w�2 0݆/$׷v��MR�;E��.\�R�t� s@�`&A�2�n�y(�(P;j�g
��X�hۙ{�3)}�Ԧ˕����[��yBۣ��`k\-K[[���B]�&\���4�=� �/B͗G�2���ܟ0��N�zwYԲˡ�"�i$��S8���%	Z��	��3Z���ayL��^�)�PG�^�w�GBr<���Q�E^�H�ƻ��!X�ݫ��& �;2��\���%�n�af��Opb��W�H.cT�m՗/J�si$�qQN�ؿ����{)Iq^j��40�bkP�)�#i&9�51��F�`�B��
�՘f�m��
J��2��el�H�YiX휅=�4z��à�*7�k�'^���r*�Z
@<���e��ܡg,T��Gu�\�aǈ��r�>%�7�V;�S\5���j�s�j�c�B�$��nh8�]���l-�"����g(E���B1�r�ylѷ l�ҏ(k��M�����-�5%�6f
mݝ9��
;x�;V� NYW�
 �.&l��{���� ����(�b��P`��0���޼߈��g�J�"�]m��S�#wojV��Ƚ�!�Q��L��c�WK^���-��\�+f��iHt��AY�l�yx�խ6�w��l}�2��y��Y�q�T3c�D
v��b��w�o��.�U��d��,(�% UnKS>w�e�qԤ0l�R�Y�X�FE�T�P;(Q{͙���,\r��$p�}�̰��J{!i�o!� �:SSڰ���S��&0��v]���ݣ2�ұ%��B�V1�R�[8P��	�~�׉$(]jB�[�zn�$�B�KT
��k
ae��sKN��n�AA[f���I,�n��͵q�tEGwI�̴l
�N����Z��Ǥ�vbAk�&
ѹ�RjdX��*�lj,�#���Xnd�OT�5�;Ԫ� �s[e�otZIQX-�9*�Tr�%�hZ�@6��o4
+m��xλ�x�Y�¨حL&:b�ս/e�Uq*�* �(�p�&w�i�ܠ�ޗe)$p#n��f��5v~���hb9Z�i
�.�ٸ�<Ʈ�P��.�<�Yy(��U.��l41�E*�N�e���4�d�[�Yr��&AH^��u���g\�4/И$P-�\Uj��J� ݢH��c���+�J�ǚ�/b&����S��DR�Oj�F��c�]�B�lA �[gh`�Wڏ2m#�Oflv�v)BCW��U�ղ���"�@v0�WEbu��������c�0�\LeF�{t�j�z>ܠ�e؆)�A��j�+3뉘�PR�Mt�d�隋Ɉ���"��-���9h&u����6�;�x��sK/�H⬉�[�%����V��dQ��`�QM����U����`�h��/I&i�
�^�.h��ܡeI�ҕ��3���J"��L�&�0q�.��r��GR�l�rZ���֜īb�He�5꩑@[j�k>ۊ%�VF�{��"LĎ��.�h4䢑�$�T7I��6G:!���M�4ĺp�׊�N�)ͤhy,f��a��i�.��Ȩ����pnCf��؎�u4�Z�Zh3�c��6��+K�����\Ū�AD��.����NQǥ��溕���ߵ;Q�p^�x��b�"�sw,S,V.Au�2���e�����&|]�[�#H*��(tvć��m]G��KhCm���:ٛ�ne�SÓ:0�*GD��rT5{���� AAdk`�D�"�ƎQ�C3�������wu���ꊥ�Jj�"Sى�W#���:AP�b�[��رX1V�	��@�����R��lK�D�m���ìl��8�J^)&�DBU��mÊ���[j�d��:���4�=^na
��z�b
M�B̧�Z����3�f�X�,_Ρ�n�r��^���h�%n3�)%�2����z��n�Gnd1�'b��f�b!f�-;,u�cR^�r��f\�YQ���qY�m-d%�=����=�H��Vkr�E� ���haY�M�]Nӹ�С���
�)V1Գ�)�R�pց�cܤ,*A]^�ۡ�(�7teB2#A�&��A��K%�̰���-�s� �t�\�u�nE�R�OǠJ��߰�^�6�]�4@I(1���d0��
(�n
��2~���;�uc]1���.$寨l��Umi�2П"�S���[�>ǹ�޺���ѵl� ���ԧ�G2��
KsE
�ڙW��ʂ��6%�P��Āt���-�d� �Gv5��ʕ�L����L_T�1�|�Y�+(�F�'6��#XwU'B���{m�F�;o+F�ef��VՇhm'��R����X�-���=v��XiU�P��Ү�M�f`�5�¼���#��d�O2���-K��D����8�"��J\7�T̈́����{z���
si��ݕ���b�]������ґ�8F�H6�,k9��&�e�+)k�v5�y��c2�mΥ�V��,�t�ךD�^V����ەx� f�{��s&��9
��i�h\1U����d�`j45�J��ԁ?���ur�eD1�&	Z�VF�J&�]dV�[M�IY����˄%�M
Z��T�
�,�����D6O�̧W�l���n�dd�U+�m������Iں%ړ&��ws�U� ��u��U�P1.\l�x�Ȏ��A`Y�QkP�L�b�*׹y�	o	[Z���YBѧ���QC��kLc�5歋~���5���yIC5,�kf0�7U���A��2����s�8k� ���b��5���R��mZe�pM�ߦ���
�$�h��R�T�̶"�S۹�^�H��w�����hH�l0�V)9�9/Lی����"���d�kX"�]r�dr�"�阵Ɏh��iASwp�eU9�-܈4�B���_Ņ�2��I��xp��^Q��slb��TYY z��/h�u{K^ ��g[%m����Z���K.� �FZ�ç>z�&q��#��$�8��4�QE��d�m���P��{Ck�61 ��MnX�^��?i����q2��gC�d�Me�[u&"\Vܶ��~7��h'mսTAj��,=˭%�@fQ��.�(E���IY��1w*5y��ٍJ�=�i�����Ez�L���4u�XĖ>Źm!x����B�V+cSr��X�xh�����b4�-U��e!�YT���YBVe����i̫���W
�H�)Z҉r���ë�րb�CwhS���J���
r�w\��;8{x[�#�Ur��)ޥ v-J6� �47V<�V�K�A)n�7�;b|�ɭ *����//��WWZv]�b�Y�%�D�ݥ�b�c��n�Z4J��t��u+	:�m�"�hCn�Vj)TX@��ĺΜ:{a�4G)���~"���le3��RJ����7����^�Yׄ��SP�6¢����?��G��*��H�|L��n��y���WJ������|⹖���ѭ/�GYY@[�����N�\��U�6_|��w�k6��IL�vy�W�xe��i��,}u������f
�*�������%#��ޭ��hT|g�:���33(����+�[-ʃVq�y�����O��$X_�.��E�6�3��b��k�)���r��ݺ�;`=+�s�G�H����)\�vκE�*�i��-w^�w:dD3���;����!��R��熘@��u�Ji�݄��9b
�tV�nm�P�����qܱ9���1�7Ұ���5O�[��7BMj¡�۾}E�QVr:i�Xh��K��Y�^�h�߶�g�w���s��P��n�"����@G���A,	\;
(��������.��D�5�]:
�\�1iR�&�۱w�i�����Z��h���Sx�mz{3'U��ހf>k����%]@D�r���Q��22�ۦP�p�Y^Э�����E��vV�i��*y���s;&"�U���9%Z����Wdn�|^Q[ƺ���s���$�����Ygp�w�L�!�.�t��� vc�e�ӒU�!qi��F�n�Az�VЮ�qum��(k�s�eD�.�i+A]���gs/j1O�VLb�o*Tܷ3xu�ʺQ��� ���;��}x3�M>�Ngm�����:Ie�K(ݸ6�ڑ��U�1�K#	�ڎVc�D�7�޾&��:E�Ŕ���zK����,`c�N⩩ټˬ]:0迥�;����4�`u
��[;���s�U�͎���1o�˘W-����}a��,y�K{�.S��mj\}GK;�O�״�+�<	��1-�TgN�Qe����.,.�4xcǘ�jh
�B6��ɚQ�z����'��jW����}7%�a����@� �������ך�ć$�Nu�0�t�Q��PI�ws�Nf
�o�X7���J�ɢ��z�s���%sh�jI��9,�)- y�7��&Va��;����ټ��㽍m#h�aA�э�7�V�����s�i^������*����L9z��3AB�}z9$	��NZ�C�C%_w,G&�Y�Iݜ�tn�sl�]���;Z�5���+v�.,v�U��u�( �m�Y�`�!�����7�P̨��F�j�u�U���b�����U���*i��tB��
I�:Z$�D�ZVO{�95zshxy�g88�{�����i����c���_<�=�ܩ�N�(��!�o��o]�p��;RB�؉��n�9Zթ��]�2�`{��HhmA�d�%^��+��ux>�S��S;A|��1T����Hk.��ku�C��]�	������-r<Cy��Z��h�hosʥQ��d25�2��ذ�pg�c��U7�c���^B,XqΫ}��On*Ȏ�z�\�եܚ���fN�mf�g�Ы��Ӷ�;��I9�����S�b,��r;ɴK�Z]�,����X_h��V䨺�f�Vts+t:f�_n�V��ʁ���u��K��XŋhW� yM���v�׸ϖ����=Qlގ��^_�щp؝x;����-������"H�l�;�q��6D��Q�1L�rl�j,�.�,p��%Lg1�V�WU�{�j�d����8Ŧ���D�o���{���C�[I�xwgW:�M�LfT�k���6�pd��}���@��u�sG#�70<U-8���P�s#㖚)��Rvz:u�����bo�2��e�{�}ɍ����,�U�FŎ�Vj4"���2�`(�k��mֶ�!����U�[�mr�hıx��^kʰJ�@��Νz����t�M�0lv��A�툅m�>q>�K,nnU�WD�VBٳ[h�)�/����Z�B3teoj?^��'5�L�<�j�_s�1Ld�(�7�RGn:ɬ�A�4K=Z�)|�L�}!n�00,��+:��	�*O�N��\��y�Ž\Lcq���ƩS�|0i
&�M��V���j���C�R��`]�y�;�����%�K��03�\����t���J�"��7;�n�6d[֢�$��V��V-)֭.V��b�=�/\�w�l�j1��&�;-	�Ko�� ��%š��;����E汭�`�{jtś{\ŭsK��cc�.�T�e�?^�Pl&z���-��:��@M�-
�2��5l�����k�:f͘�Ir
�L�$;��9�4�콛!K�E6�r=�u)K/mJ�fVTy���{�V6k���]6�/�.ՎEX�}͛���Ʃ.IKw�tif�]{Ec��H.��K��oo�e�2h��l�V��Kŗ�l��5��u��t� u�r�lL>(���r�oky�;,1�M���*:u�)F�.v��5��a�V������yb��q��BE�YM݉�� AIָ
���ھu��G�Q^r���n�tS���,���k�v>�f���kR	A�k2�.�i��V�\z'�)�᝗L;<���W��Ԕ/ �;d<k��� �Z�>Y��)2�KC7�hێ�^"��Э�:{�f�n.����e�e���;;�Eؾ+2�܆��t.���]-^�f���?!i�g�o���{;D�Dt��fȭk��΃��gf����:�֔��q��|�7F@ %Li�/��+>���\�j�Eg OAw8^�`�}{2f��!f��Һ��T��3z�-�f�Eh2�Zz�n>�y����9ֻK�]�b4d��a��"�չs�Ѯ&ؽr�bK�E���)ơXy ��7���]#�ꋸd�w��q=�^$>P��z�V��hm�p�h$x�Ƶ�ޥ3�n�1 ;"t�2��:׶[I!"���D���6��v�Z�u�&�RK(֧��j�VSܸ/����ұi���8��h��Z{r�x�ZLWZ�GI��s�u�m'�Ƞ/DʛǑ<���Xڻ�l����z�W�r��[���#l*b{&�L���`�.�dT��_*�Z-:��l�e50Y���[u�v�Wm������G}2V��hZ��&�����$S]#Uyb�M���b�m�1���{��z�n�V�&3o�z9�#�a��\���5�3w��fm6m"�,�����y ;D��9ꂹ�j�+��{��v����i讦�*M�a޻�����]�v���pT�:���},��5Xc��^Ω�\^�x�#:�Vp�9�b��&+{�+[�R�����V�6�>�|�����׽X.u�����9�r�A-��Wy�_˶r���\�A��>&Ѭ�w��|joA�P�(���ʍ��N�b�e�)��z���Sr����e�����;����riR*L�Y��W�j�Q�sub�$��o�Vm�&�(�q\5w�>H���0�Xk	;�{P'��u�Lʝ��<�q�Sp��t�n��-��Իa�;ws_;<"�b�0��0��I^d�Ht��׷�B�3�C���`�{��L��7�Z`���V6M$5ܡ����o#o��w@Bҝ���U�Jٝ[.���WcT��Q��(|���!�R�L��9��y��ܷQJB�R���S���q�t�|N���7j���s�\it�RΦ(?z�~� '�Ǡ���y�e3�+-����>]I�mV7c��%* l+���������|G|��w��+�)�i�zkH�8�=��1v�U��U��)!������I%yxǋ�[Ё�]ν�y��0`��L��(5�Kn��wn�^Ε���o�HoO�\]ps�ұ�U����{S���5W���}�n,��pJ���s��������lͣ�;�����aJ�|)RĀ�2�SBHỤ�jNY�sx�R�c��vsFPv��}�w���:P{YB�uYͽޛ��A2��/��U��HHȭn���ȁ׫T��9��;��T�r���Q��;�$vY�n��=�ӵ��IDNRe��n�t�پGD���ݕ{�
WO����M���z�kci�<뺎L�*�j���&f��.jJE�)v��8�o!T*f�2�-��淵.����8F��P��4�r��8e��6�H;3���Ԥ�t�(p�s3���{��X Y�YO�] u������nuF�Ʀ��<Ɔ��s���o��I��me�4sg&�1�I.s�8�6����K�e0���U�a�${ś�0����$s���U��3���w�߃`��JC5'0Ga����nҠa��Í��`�Rr���MܥC.����R��#���.��jWF�d;����^��v��R�;U��p�"� �vk��`!�����|1�c$b4ot۳�{��.H�u��x(�ƍ\��-�)�C �ʭ=e���5�wf��]+��l9���;.�h�N�BZ|�6��X��*�W<�Sr��F�f�Q]�{}�H/��D�t;D�7����vK"D��YG�*zݡʞ81���[��:���.H�b�c6���qY�_T]�9��jl��m��q�����M��xL�n�X��5�gWBCf�Uq�g:�^t�烫y��}����Mή�Q�٢��9�vq"�N��H #���wi���툂jv����cr��if���T1����:p�@WP}�F�m<��ݻwY� �a��c�( ��.�$�+�`� �N�V%'v�9k:�.�4u]�up�Ė�م#1�ԫ^4���-�b� ���J�R)C���[��l@��?s�0�y��cO�G���y۬H�p�!��-Tۮz����ʀ8z|):bdi��qR#+�}��J� o!�4��f�,�|:��P\�H���h �5ڀ|Ʋ�r���+'lcׯl�G.�^�Z��B���&�Gzy�R��څ�o4@>�_Q�&�t��e���ooJ�3^��,p�h���ڠ��b�TӶ3�#��
}6Ō��h���q�S ȕ0X�䮮as2���@G���fVwQ��i�}8V3k#��ϱ>ò��9�
�6�)�n���VXz��%NR�:��p�M����N��[�\�����FC�u�����{OpZ[CuJM+��,�we�HԜ�k���؝N"�\�C5�Մ��p>Y�������:�t+W��G[�9���i������Ɂr��������c�Y,�	(PHp�ɼuH�T×s[���~�o��b�#���Z��>�Gp��G���_L�;\=�>u-u�Ef��Վ����ck�-�̷Oxp���f�.5��y������s����vD.�l����"������r�x!�q8�� ��B�t�vnX�t�lŷ���s�f�;��x�w��l�Gn��l����ObrJH,�z�ݦ��ڊ��t���Tb>�4�r����;/�-W2�St�#d5�U��4��P$��#G�ơu}eĲ���{]֐�n�2�*�3�W �4B[��00�l� �'������<6V�5��yK$���I�*H�	� |o�N��f�>�l!�\b��4׻6�-P����:����r�|�G�E�0�o4g]Agw�uHN��	��&�H��Y{=u�uZ'N=��n�A�����a3T����Df��$L�q7\r�PN���f0�,Z��(i�h�U|�9�yʶl��ۛ�5ڟp�� ��F��f�G =�f��|c���7Luv˝�[����9�Ҷ��&�9���}5�l����[u.��QԸ]��n(WRܶ�F�����P�Y��>�|t^��C��|��#~���lً��v�ܚ��1E/�b�m3�eШ�<��d��4�5^�Ykv��p����]vg�+"�lDmچ��C�1�bn\���X:� �e&멇��+�a��\y�M,�y�;8�������ՙ5%9O��U�4�QK�3�!�)��cm�(�瀻�o6i|@��QK��Ŏ;�j����ΰ�N�1 ��6� �������[�Ƿ�oz�l2a�eA�(�}Q#%�4P��ɝ�B*�Mr�=�S
Y׫7���+�J�\�:��
o�E;�آ;��w!=��٩P�B����-`��m라��q����)���k19O����q�'����ф^�=Ch�Х���u�79S��xێ��i��b�^(�39)�[y�Hvc�lg]�ʊ�����1-]^���X���Rwh�K��=���M/k����ѻ��b}���/'-�Ǚ���뮺���l�,Qޝ�K�AVӈևWzG'�����i>W\�\�Ս���|�4�<�on���r��DΣ!X5cԨ]�<;R��Tk݌�����q�ڂg+���SU���wBb�>����;K�6�v�]�b|�񁛹��:�)Ǐ�$��|����޼���d^������)wr���0FW^��J��ڡv5J�����p7�K�:�vVY��oHt�C=×��o���f���65J�MU�]3)Hc� ��Ƞ2S�Z��Ób��ٮ �/�̤���*�`u�y��wa{���\4:����gGu�]�E�d����>kN�+raﻣ��Ԩ1�&�Y�k+�ܗ�:����5|mNr�d��H͠N�!�*�tw}Z�%;�Hf�v,�id�6�@)���Z-�e
`�<�'I����]��y�2�w3%t�,�%�X���Q�o@��>�9��_[��{��GA�=�[�ru^,w�_9��c���){��\���֧`���n힤�{��ý��]�.����((W;y�Y���n^7:��x��&n��h�X简��r��� �<����3�������3�_r�kjWM]2Ds���8M��hs���;[�Ε���3�ӎ��qI��6�u-��l�Z��u��K_~���w_����|~���ۯ�BI	�B}�G���W��������ڛ�T�j���僡�J�.����X<% j�M��7�mj[;�����E����r�i�>���O�P�ë;�D�K9���vm[�jiִ	���/S o�7�w}.����d6)+���,[yG�� eӷc8��J}����ns�P��z2�eHJ{��`r�"��v�LB�z{���Ī��w��tT�x��w%������]dd�q��݁m�i*��4~�T8ȑ��7���m,^<�׃����m�/]s�^�+�������oK�P��\��B[lp%*A8/�bX=k~�j0I��lf.�֖�S@f�4*:ͣM��k��[t��)��O���ҥ��f]��n�ѣ[����\:�.�P}Ή��Ij�:�'�nu��V*��@[iVV��Z�"�&�ú���*�
#�f���^<�Zmɛv8�w���a� )hǓE7��
ںi�.,��ԕ������ζv`��u��{j��r�q�p���B�m�v���O�m�2��5ѭvm��#����w͆��x�7_d��b�֩����ȃt؆��c�9f�˴��4�t0��tih��beļ,JB�H�IeN��ՁAV�[[`5���<q,o(d5:�v��e�K�e2i'LuU��oܜ��l��ݰ���3�V��ѳ�PIo=\6隁��s�wXk� �7v����v� ���6�ᬭD\��g�9���,��چ�'�]���E���}K%F� �o.�>��!�LVA��}3��:^����*�8ؙ�wmM��2r͙}��uJu���ex3#Ύ��W�h���z� \t�3З�WSݽ�re���c:�4m�%�/fh�|�cԯM�6���+>*U�o\��f��]SWd���I!]�r�t�A/6�ֵ5�	��>9b9��y�̖B���Ad̮}3b�-[#��͍�Ę_>�qM��sF�V7R��U����h��k��X�H��|g֡b���gdw^|SLV�{L�tl�3�Z6<ue�m��-�O�GLݏP��;��ѭ�v8\�nAZA�,_E���6����D��BK�WE�X��G���)wT�J��w�����ԉ�$pV��n��TMͻ)�U�DjA��"�$B�T���PJhqh�̶.�QL��mຘ��Ǻ� i�5��0��͕:����P�njb����H�7�V�-[�����ErQQ1W62�fV���I1����B�%|�_�R�S���weP�6U��;��Qvm���9�\ӳ����ݛ���A�roc���h�ͩS �1��ًn�:�IP�Ј�G*E͂�[�T4�,|�\NCc���ҝ��6��d���!$�	��l�ŃK2����n�R�����"��^$�����e���nх�k^s:V�r���� 9�ۖ��R�&�f �m�����U��U9��3[�l�Y�u�(<뫷,z*��@N�*�}{�u��sy��8�t �c@���X|�A#�H�+��e����ȫ��/	P�CK���[�`�]�0#D]$.ڔ���b��(Q�-O��$\Hm�s&0B��/�]W·V-��wG�N�_W�	2���j��i��mbU�vFS�j��M;�{)���M�%<|1�4KS�b��4sH��2���ԫxb<tp�[����fG��S�`��YS&z��J H��#�9{/VpU�t+�S�t�7\v��-�y��E�a�!�'|�͋�m��2WmmC\7��j�񳝘�Y��JƜ%�_1�̽Ko�Q(��X�Yה��Y��8e����:��>�)uN&��O%iۃ�]�P�V�Q��j��ӫ��VV�n�wx�;Ru�r� VV(;Eu�����rb�y�Jh#R��u+5�"5�t-*�����u��h�ik�;�eˤ+����kz��f�y��V+�_X�Ⓕ�D�	%�s(\dK_FbY�T�]�{ji]���i���؉����1�	cO�����rM��we�l]�WhZ��<�7�i�jzS#m�{�&��{��Yr0-.���Y+6�Ö�G(��]w��ϵ�cfv����}�↞s�
�52�ѩ1��MU��i:�лrۺ:'���x��f��D����� ;��$��dN����[�%�Y�gj�[i��ű����q+�j�Okŕ�N���5�ņe�U�1>�wi��[��+�x2-y�E���\lR�9�ݻ��f��ў������
�>�z�n]��I�n��!��lM;�8�mxܷA��ܣw�3C� ��[8��C.�u�#���Go��'gn�f�-,\㮓l^e�Ts�y�o�f�I��%{p
N��|�{7��	(*��8e�˘ R�b�'v�Wm��1ǯ솉G�YT�V,k��HS��`�Q���6eT9��+ޱ D�����;m�ncN� u�Fee١��b��B70�9���J�՚[ؗL�
��$
"6�	{����+����z�f�#��F1I��x��M�@���$#X:v9�e�����t�����R�4�͸;b�--�v�Es����c�գ�\E(��
�u e%:�g/��!م����oe�Y1����1v"�����"�5undH�G�7�f��a�P-6��b�w7V��+��S-�ie�P!�e\\M*X��ǩn(����Z���t>q�K�q]Ɵn�4�x&rJ����>�ʻ1�ӫ��<��3�,��@�+*�k��ս���Λ�N��U�&�7������\�^H�>$]�"�v "�aѦ�+�Uw��ݭ2�u(���@��J@ ��j�Y��{|6���@KK�����/-������[m��b*p& p�]5cڲDW��������v��a	��7l'u��"lcm�l��uw[�6��30�F�y�(���`�3��-�=]}��=i��rW
ܭ��[�D]tX�2�-[ܒW����ܣ6۝yH;�Ozu�u�gr�S|�H���5��Z�Syurٴ/�eC5�Yy�F
�U���aaK����vQu����vd�Gk��O�V㾋mw,!�{	�PZs�=��ȾO�@N��ft��M*��:^r�w��⫐���8FV3���95�%�ʴ�86��ȸ].�sڝq�gvBo�&W)B�'����Л,=4�o:�S����y�G�wL�gܤ��h�u_H��c$��th�Z%e[�o�f!.�W��o����/�ѕ7�#��B�Xz���Jܧ�NY��S��Ts7�(N���1ُ�����qm�Ĥ��p-��*����ٯ6>�e�gF�ֆΏ2c�HhB�����0����Vl�WaY\��(�Z�+}����0vְiiȞ>�y �i�B3�-,��ux5ޱ��Pë��-r<V�{vV=g���lD��>n����F����K�>J
�^85��n����m�n��<d\�OZ��M�4C�Ɇ�la����偒��:3�bͩ�]5{���Z�����WD�+�Pۘn�5x�["ߙ�O�u|.�V�z�Dn�r�S0�qs�jو��Ss�T"g�@�G/�!�M��$��[�v���DƜy�[(i�zu$���+cz�A���mwu�3k��J\��5�/���|ͮEX����mį)\y���du�=7�V�lʏ����P04��;+��jJ�N\d�9hB�ʥ�N��Ʊ�ɜ2 ���_]t�ϵ�LnIK�8w��tp;^��ޮOe��kkZ
x��F�Tvp"�f�I������7���ш]��{S*,t�m�3ݯ\r�t��w4��#r ���k=�\���o��-��_4l6���������Ɇ��X$[�p^�}� �eu���
U�8"	�K	|*� �{�a��Б�A	zhq-����E�)��F���Fc�8��w�<�C��J/v�^X�]WR��tn��H�Dᝮ�i�y�:�)�J�f�����(��mL20�&��c��R��먪ֵwλ(d�&Z�R��p��P�8"�,. PS�w#ϸrmS��d�{E�3��0�m�x�`�}e�5�5<��p����9`7Ykh�hJP&Z�!��w5��D�W^V��3�1�J.S�}�Ɲ��(�줸i�·���Li��i(Ǳei/�'uT�g.�Z��u����<�5)��(.ZѮ�{�����k�x��ڡú�髶R�]u�O �ޜ���1[
`�%R��2共V�a-q�WrU�� P��m«ww[E�2�N;ݢ���4Ҡ�y�\�'��d��U�,7��.�)Cw�кݜ<��#���E}�rje�ٴF���V�r�y�	W�qc[}�h��y�ͽL@Ŵ��\{q��Q�$��T�6R�p�P]���=�N��u��5��'�14��f��C.�weܔcIZZ�J�Q��'8ث�&��yRQ}���It����^d6�G�JC�Y�t�DWF����S�ZضP��FLeR���h%Q�~}Q��ť�n}i�v�'C���V]�`�f��>�y����ᜟA��Po�C+y��t�<��f���R�(n��f����]��j�u�[���RL�6n0��~�;�u�m�0^��p�\M\e��5`c��5�Ԉ�z�Bw�m�׳��	�&+c��C;N��!�X@ˁ��V���Y������+�)���8#:�-Ca��wڦ�����T�v��H�]���\*�bO������ғY���}O4.\
��z�+f��i�m���g+q�7]����o#�,bt��K�qJA&��<���,8�dJ��S�¸0�ƜG^ 3[)��g-V������
y	\{�[�|x�FJ{N�-i�3�qOo_�R�:�n)g폷��P������nsm�eWj9��s��"<�%�[Ҕ�^�qw[`Bʵ�@֬�Zo%Y�R���-�r�<e�k����	X�*Nu�*���Df��+؀��h\�?o 虨۽KKڽCwS��8*k%B��v���'i��W5ED%;kr�ip�@Y�yHf�Jq�P���Z��X�v�n��η���t�6�wd'���%E'-��ۉ���#{�1���*�&����T2�r��K�2iɼ�>�0�F�odpv7�z�m�ӛC�Z�-\��ׂV���ݽ�W]�I-1a�6�v���;(��v�0X�
u�5CWu���w�0��tR+�w
�z�Sv�eu�R�-�=���˶��IZ�u�[u�)�����#�4����ƍqpB�p��zp�ɝ�}j�?�˸�&_R����'F6���avjt�-��NZ0��Jq�`��v&�p'l,lR��'�]����&���:��4�<��sJ�ю������C7��T8x
N��-�7}ǫ7�$����D!
�dšP�չ,�
���������F������`��u7W�ѩY��UG��Ju��8�-�:�;�uյ]��L�7�I��X�E�}���&c@S�=��y�L�N\�r�ݨ�YJ-��MTR{c�f�>�e[�	����O%[�j�4�����'{���ӭm�yx6�w4���
Q�{Yo�&��	��t7���>o��^�[2�A�7�>g1[�!5wُ,�|��R���\���3]���M�+��N�ֺ�(No.��nB[܃z�j,ZՕ�8�,B�gn]sp��u��P$ @h��n�'�Z��.̻���	���:��:!�|�����W�,}d��VL�̮���`�+�#�.�oG�����K����"C+�<�&�@sxZ���4�F����N��n�k��� v�_k�ڔ\��D*4-1�����Bn�v�%�`�WP;�bL��@�I3.F����m�8+Uh)=ۂ�֨-���ڱ�������R�L
m:my�++)���яT{Y�lٴ��m�-��ۏ;C�9cy�qo��Zv���J�>��=�o������'��i*뽼�Q�͊�sk�<�Nd �	
kI��XU*H5�:���8Z9T�N��1�p�> 켼t^�6u����\.��I�UՕ�\���H���۬]�fj���5(Z�xS�޵��C��41�=�g0�v�R[JWG��w�;%�U�;��Q�\��R�-���s+j%��tU3K��|_%�V&3u�t��.��@Ɏ����� �d�������S��Z�QyYY��Ɵ��ѹ*���7W"D\�v%n>n8���x�����7��u�R�ٵu8��^,=����7�-»����h��q�v��t����hǶ���tv-,^�QsV��+~CZ뇂/`��.�ԅ��Z�����ܫZ�e�F��U��k-v'ۺ�0fGaȣ:�n!��,�/E�n}�Mc���Zjdx��xEtbVn��3i�7��䢣�|w�N[�:epu�Q��(p�;la�2M�5ho
�:��Ԁ�[۽x�
�T�����h+kw.�ѶH��X�6ry$t�@�f*_!!�}����y�
�F^���ފ�d���Ն��Q�ʱen��(�Ҁ��d8,J�;eE��Ʌ[��z�' �lR�)�jf��
�q�z�e�5Վ��,.�I��^��6ɫj���_�Hh���*���P
��Wc��`r��Y�>/H��Q�w���m�5�n�5�Gcpri�V��&�{�<���v�N|�ۡu�APTl���m��W3� &z80�T�q`���䠾�ę{[.s"E%���ͻO�-K!e�6���%�Qn����H7nf@4�R��rW��kλ�L1��m�vZ�n�>A��N���ͨ�>l5t��0�t�;)P���n�YebX��eZ	�I{Ў k��E�,��
K�t����_�������ﶪ�N�{^�=nS�^�Q����$��]:���K�V��[���>`�rB�I�Ml 06]�J��*���غ�o�F7��j�&�k=X�Br�8��Y���[�gv_MI*�S�ۇZ��%����T5�Wsy�)GwlJ<�K�n�Yr������|�8`���P挮��>܊�9R�b��c�'_o^�����PW�GQa�9�{o'�Gi�ź���U�^]�R�"#:�S6]>̧������[J�{ڪT�.�v�mc�f���K8�*?3����q$�L�Y���+�b����iu�1��&O���ܻ����#�`2{���Y���Us\9k^�ј��TR���w���87k]N����|\#0a1q�&V
�v��?Z�R�a�V;��ouVwP�;7�|�U[V N+�3蘤,v]ҧ0��m��pCN�h���(��Mj0�L������D��N'��^*�c��;SS���;cu��� -�T�V�7�Y�@}m��-nYY��[�\~]�)����ƺP aeB�mv=K(�Yz����
ܭ�B����})�(qI݂u�]�NvG�<�_1{Z��m��P������L:�;n����p�o��5ؚ���7s#�Ijնt���t:�X�P}K0�D��Lw��i�9Vq�mG]}��� �um�:��v�ń8�w�l��E��jChԂ�P<��&�e��ձb���>H`��1 �d�c���+
�ʖ�YYR������%aKT*(4�([J���Q��P�J�%@�C��R�Y+Y"�H,*(V,ZZ�B�T����UC*務Q���Z �lY+�J���4j���QIP+����\Ld��
��R�B�R�q*c+
�T�1��&$�%�.X����J�IQAE ���ԨAdb�
Ŭ*J$���d
��D�,&3Lb��B��[eJ�J�T�Yj�1	�+�*���X�YQJ֤XW�2�%H#r��`�� ��ZʂńDPR�+L�E�i����f[�QaXTe��d�"�@���=�߷��)��Q˜��u^gWp=�ʇ���B��s���u�G8�x,a[g{���i����⺪�uo-]�EX���%�]Q v��?-�lخy���^�7���� ���i@�V��:]N�>��{"���p��DPTk�h?p˖��S�uX{��ܫ "��o�}� �0�ۢ/_>;CC��`w�o�0UW�x�ˢ�+p���G�!��e�3*u���׊�����7�v���Kj����籚�Ƌ�"��:
�:��RC�~��1F\���O�ʘpU)u�fj	Ű�~j� �'A}��y��4x	�9��p��fi�q��ԣ%����֋�u"����4�Ȏ~����`�f��:��Ou�Tn�k��Ş�1��T����y�����
�m�*fqys�����w)�.�G	�>5}^`@i/�����]�ΤGMĸYĆ�e_I�j�],�sS������E�i�GaZ��6�'�qӞ��4����#����J6�r�Bc!8���
����p�d����0��n�#r3�;- �� W���Y�E�s���|��|��
؝��{T��ۙ��ӱqc{OQ�`�5&�J�����Q��I��˝�7��������sN��"�=�Wk��X���_a;�-.�[q�eΒ�m����:��_>����]�5�Υ8�]{�|J�"�-�p�o:��v0�f��q-��-t^>�Rb7S��n�I-������bP<1�d$_�ٱW
Σ����`���>�:�"v9'���#����r4&֝���mg��34xv�3;I��rF�Kp��w)M-O�v�z|O��o�wϬ�]�]��� �O+v�O�H�beɭ�q9�ȥy����g,����p��b6�BBȩ��މ���B�r�W꠱RZ��v�=���'���L�g������eR\4S�G��.9fX=�6D�I���VT�̻L����'>r�ׄ��w��������yPYU�n|��Ny��[g�[8�]zt��n�����Ds�v]H������|ȋ��:2K�/�mх*�폛x0+Φ.���-��+>P'��&�Ĺ�"�R�UXL��Qq��z�g�f�dM�����R�F�lS�;e�Evb	�S����ڇØ�ݹ
fo�9r�¨1:�n��W���j�
�5�����烁@�c��/M�h��7[֦d�ڦb�z6��թ{�jϧ<)ѐ�������'�G�>�%�kCe�r���>˂�M|��ޤ{of4rs���ǆ�m+�6#S�oC���ν�%���rv�T��
�ob����*lb�.���t����aIK�)*7��%]����yLj��^�k�t���(��Gh����&7�^������<���#f��<g���V�V�^���uڼ2���G�h�۬!n�����>�OŚ��WN����ty�����*��3E��}د�%�=�6"yW��i㑏�0H����z��v�"c&	��v�M�Fq��љ�ga�=U9��W�h��k�F�m����F�dj3b�}�� Ɋ���_խQ<�Ff�s�^�!t��f���F�r��Br��嚧;/�-~n� ������b=�wh3���N�K�I�N!T��#��|�E%d�4m">S���_K�3p͹�a���{�ܬ��/�N	���Ü��y"Q���S���H�R!��#���H��nb�ɮq���U��@�"�L�0{�:1=�莠u��G�:�*h*dFL):3;m�Ұ�}�x�[[�h8�m�[�n�b:`̷S�w�,L�,�� 5��СS��=�]]�7�B;do4��}�&_���D9�I⓴�c�߀�N�)�A�o2�"�C�k���_������
�w��s|��	��3���N@{,��m�S�*M���W��}�ǙY���H��{�2��TP���]�9�j����{-�Xg ��McC�nĮ�(�|76�H�5ۉݎ��Qd�}����!��ש�\��F{��pV��M�=�Z�ϕE�l�]�	ӹ�_�������?{����CÑ�%�9u�~~;@ƅ0��sӐVM��*aJj�_�l�^m`���Z��^��������=mnx��O})����U�wښ���뙂εG��9�vВ��.�Ȭ��4_��B�ʧ+@�s{��w�����f*�b��v�Y�S����U��Yb�A ��u}�Z�#&���S�*`�u,��ȭz3/gIR�Z���U����U`��#a�$d5��3~;���*a�ϰ;���{g�n�{���U���Pf��BgZ/.x�ۘ����|#VWOd'�d��D�9���
�4ʝ��d�&�2�P{ٟ,��nF�x�����o��3��M-O 6�/�������\6bSG���ig�t�[ǝvII����/@�u;S�)�=�N��z�ib���2�ͩ*���b��6+�s�}L�	�
p������ECW[��c�z���8�V��EѮ���Dp��u)Clӓ{��)����o���v�{,�B�f�ʉ�.�m����8,J���Գ���/�4ఋ����a��Q.un����L���@�q���u(�������N�"�����+�s�c��m�@�9D�a�J����M�ǻ�@��Oч�T�$VEv�`M��f�l�w�I��w�W<HF�ԫ,lp�f�ҘX�[��`@H���BwY���{��hf3^��C �tJ��˭�|��0�9)��˰���\�J�.&�Xǜ%[S�bm�����!��� E�J�� ���jԽ沥K"�:%`rw�)L,���N{�����f�9�DTX+>�s��S�R}��^zp��c{�K�}������_}�ū�����a�w���TW�1�-��y��;�U.��O��(%���X��mLƸ����aE=��>#$I�5C=t���+~��)�$�����=��)"��FV}	��ň�!�Л��{�ƌ"&N(�߆җ"�Atξ[x^N=��驇�����s$�w^���]�C��1s��᩾p�r^D���"��4�9
S��S��93�Y_ +Φ>�j��Dw�p���x2}����8^�E����=NM}Z�ze!�m��h�U��A5]:R�Oh���YD�<ӫ�'[�ڎH^!۞���I2:bp�֖*B��w"�l������PK�(3f�ƣͻ��q�.�V����E-����l���)f�ƉE�˹%*uK�����=���(lW9�ŋ�ׯ����`U�!�@�L+74���]RTì�z4f���E�K��$4zsl5~.�^��G��ȯ_�|�UЇ�,՗�%S̤� �j��B �ˆz�z�jk�'�����3ҺU�Ƽ5��q�o���e�1D?�K͛��|1��#{��G��Ph�w��KX��:K�s�^�` �q���;QT��&a���x�ϞDI��α(�22�ό�ޅ����ml��`Lhqu��+��s6�]��� ��av��b��捻��|��<;~u:*-={c�rR�k/Y�ѫ�B�Q g�~�(%eٱ �Z6 �/2dkr��+vH�Lڑ9/iСӁ�K���[�;.z��[�WȖ#�BB��̮���� OM|�l��褶.�fQ\&��L%���}�B�< S�j!G�#).)ѣ����U��W�	�|_e�o�mYU��[�zp�Κ��n�X���Rۙ9��C��@itUv��><H�ܫ�@�SR�S>1;��,���X�Ա�ǈٗ���\��u�h[�w/�Vե���]:�-P^���%Y�]L�0�ꊘ`e�↳5���v3�B�a��,�t�*�)J��5�o��v�c���H)��"������	0?�����-G�.[,�:����GЉ���֮�gM٫x�=��آTw%��*Lv�=��n6Ҷ2�����^���b�(GI��]�"���''5'��S���\l��S�.\쉨=J^AW�9ȉu*��sB���p;�,o�dWȥ��H��z��D|���7��!f�>�H��.̓��ɇH��<����9����f,���{��{�K��j��v�?��rzo�Ee+�;���]�խ����:���F���l��tܫd���,tă��@+ڇ�Y�8��Z�D=ے��^]�^ɣ97�I��Ӵ��_o�8/��y��g�e/+�D��0y�W�"�8F���_'ƕ*��I<�������֘$tNOpO���X#".�ԃk;��5�>s��#Ŝ��ڙpj:zp*��Y�EJ1)��D&����ג�D������!���D+��&o��VR�|���<L�I�ȦU�R�S����O�ct箤��lu�2f���Y�^��O`q5G[�wVG1������~3_,}���y��n7���Ԁ�ѳciG�W��#Q�ADI��-U���y�ǚ_n>��H�W�.�tz��9u"��Ժ�u+ћ��/D<��`Z���_���`�Q�h�����{O�&V�)b��гU��3ogv�]��wz%�DE���WVt�]=X1�����$�)	������N�ƟԼ�C��..��~G !���p�˹�T6^.���6���ebf�+f�n�N����V
�s�9Yy���e�g�=@��|֦[<9l):�6��m�V@�	�������Y���7nՄ�3�U�5Q9�u#�����'Qӳ�S�aNtjOnN��n�^S���"Cy�.1[ i�ti��[��]���oHN+/�E��}��uW��z_��_��s��5r�	��u]-�n�s��͐z3Z��D}�X~|���J:�~�刼�¼���,:ށ�M��xX�=�x�pt}��<o��Qp~�� B|0P�#����s��������N�ej��
�z;��V���(����Eg�о]��̈́~���2��Z2=�;�NV�0���VK����߮, f.�-��)�q��\.���rj�pg��f�e��孯�oZw6��$%�cv5�y�d�ǡLc�ћё���di�2y\9���aW���{��d)�v���ei �6������N��jRߒg�^3.��>X2�.�6�u���׷»q�M ~"��=��v�;��湉�-uYٓ����x3��}�-t��A��:��b�Ƨ�1��MMoW9�goX�~�V"���ZU��_/�}[��֩��2M�O�˷�	N�pפ�Y~!��a�*٬�{���+%^b��aM��Z���ϖ�b7"5<Do���꺥���8�b���T�T�os�}a�۬���ùbQ��u��o���1��ς�iV*=C�4��%����̈́ �NL��2�m����h�
�u�� ��
p�|m�5�۳jG:+s�l��H��'���N�=0����Jb���xK�[z��Bn��bzن��6�l�+/u��R�]\�
�s���@�N��!J�a�s��nӘq��R~	V�3TK!�wA����t�\�=C����c�U��@�B}d*�u$=1��Ǐ:�eJ]�[K:�؞C\TT%yh�/F ��ψ�/>i�a�R���
A7���$�ޮ��KW��K�'v� �t ����ep��S�x��^��.�S����=e�&)��3	vGkH��*�c�9ə6�f�y�@W�˪+��5���^��w�]	�����-f������w>�,�<�����:�8B$X���[L=]�յ��T�6;@�Ƃ
�0=v��Q?mh�M�+�2���ʶD�f+I^r���}��:4�;"S����Դ����e��>d�u���q�8�����3��#�`94�9�|bT����7R�&'e����+�S1��`�șd8��>ϐ��xW���׷�7���Z�yz��֎(VH�(�(U2iK�Ow~��%�|��c}�e�DL�AS��A�bK�=�v�~Űw�e�8�1N�xՎQ8��W�c~/,pϞ��6lh�Rkwi^$N^Ե������9ѵn^�&'f�\m+���L��	e���ϡ���u�KN/`31�W}�{��n�螰��Y���T6+���!���B8�}����y��%u}巢{���c��o,��I����'�K��Hh�_��K����l�Y�:��}�9�qx���^㿗��Sӌ�ٓ��A�A�T� �g�u�ɏV/9YƑ�kuuX���AC(��{�-	�a!���͡dF�8���q]S0�	e*�N�<�퇻������廨ͣ*b��Լx���%Scga�`��>/�s��X`����Yn��fN���vZ1xC��e�Q�� C��,.F���N�jp���fh��fvc���cT����T��5�J���٨(��h$Ьo�
�<�&#]��s���;]��td�����)A۠bv�+{�.m
룍;�f�>I+U����6L��ɸ|��z'��]�fsyW�/��V&�4���bsYh�n�˼P:��n�ش�v��ҎsAZk'<@����:�Z0�.E�6!�
�3oyoWv���nó��uԈ2�Էkb��HZ��f�*�"��1xw��.֫��~bgQ|_ O��H��
�3���bm�v�Y�ᚬ��hR��ُ�X��نI]ą!y��^*��_�p⣽�k�#�9ʵnKaQ-�@��[{̲�+ŝ!_t7FY�Z�ec	mDFK�,���x9����&��^Y2�W��:X� �vPs-��7t��Rt���&͇(%��F��(���c��^�M+I��I�H��OQ]ӎ���,�z���Y��3n��=�7do����j�NU�q��`����;�ū�TԚ���<��Yo*Y+0�6��k!�V�&��B���x�I�N�ûv'�䭁AR5)�����3�}����A����u��{���|˪EZ����%^˚�449f������m�c��	wa�RE����u�[BC��!�iw=V2�'$���E�e�\{ewJT��>Ѝ�����=<�lM�%�m���Odz 2�,�7�]hU�Z��[���\d33{�'V8��i E��g]JZ��Nqg1p�R��!=V(^V����;��r'B_u�&.�ۆf�km&�����<�DٝRC-Mw�Ԝ�06��@����=w�a��+K6삲��K`��iQ����WG���M���L�M��X,i�`���(�Z�Z�C5)����F��e����BQ7����#�ôq������)��L�$uj��7�|������"��vx^`O���)}���̺�ݘ�X���tR*���n�3u��Wc���oj�`���˛��1����gY�Ҏ�X\4sb�<�6�Ӭ��dG����W(czV^>Z�yX@�ҾVu�X,��C5��:�	��:�#o;V$ ���ٺ���)*C���\*v9���]ì,�5:�$Ɗ �s^Y�̢�ƅ
�]rݻ��!Ε���gwM�}�:-c.ɼ��$yR��������j�֬��r��Du��:��%%Sc0v���:,1y*M]�qs�(��ki���P-��������1r�\�V����c��x�ի�"9$<d(GE���ݫѿ�t�=�+f���)w#�.�n��WV�o4�;D��/�	���R���0��L=�-�]�\{I�K��{KIUլ��5�~�X�i����#��ɤ���&뭠8��o�!
��[I�e&�� hh��V{r�!����7���4��m���x,q�RM9�Y
\h��˩Z&��'6��چ�Dd��t��
>9�d:��K�l��1�^������J�%�������(A���I�b�&0XZ,V�
$Y��V��P�b`�U
��b�6����E-"��aD
��"ȌB������iIjR��c1��E!��+RKm���U1���$�*)+d@�"� �U�((�ʂ�Y"��Z�P��V�Q mX�əa1���IRVA-Q@DF�`ȊԅTĘ���(�+$�YF�@F�(�J�IUJ�(�)Q1��ưX-e@Z��VTQB�U�*Ь+YX,�(�FKl��%@X��)�jV�*�1�T����(�bV���V�b��f26�T���̳F�ʕ��E��Ŋ�Q���z��zL�����n�K.兇�i%]h�a�v�{Q�!ٍ6�L"���R�+���Ki�c���HK��-b]��"�5��Ͷg`����
���G�b��]}���H*�["$��bMCX'~S�|��Ă����C����~�LT>aS�o��<H?�>C�{�V|��i*y�oGRm�q�ϵ�����C�wuD߼����#f#&"�*fc�G�"�hVz�|��\`x�2Vy���uӴ��'����b���e`)8�LtyC�|`Vy��~Ou��$�(c8��~O���g�Ru��ҭ�5�?g��1���mmQ��1�f>��}�Y��Ldٝ�Sğ����=�si?!YY*���b����1欟&��nj� q+�%FزT�B��r�0��Xa��5���1����bNg�ꝡ�~>/�1~�51���b��Ğ�·����AVOɉ:�`}��n���6�=�2O��%eg��D���!��;f+*K�Lf�]$���>�>2i�Qa܍U�c����o{G3�&~���1�?)�'����1�!����d�C�+��2yi�����0��H.��Z��:��f�̓N�����<f0����i�f!��?!���tKF���e��,�w��3g�N���x�_���=��g�*��P�J�M2b~�8�Cԗ-CG߲I�+�M��拻�C�.��OW��7;̓IP��T�w���mX
K��}�<�q��+���;�nn�wJ��3+�
��ʅLa�m1��:�C�nk��Rq<����bAx�{CH,��&!��M$��Lt���Ȥ��au����
��T�y��:����k���۷�Nw�/��@�]�t��4,����RViX=�����c�5CHu��$����a�Agz�l;�
��t=M$�
����P�?:Cq���s~�O�`��-:5�H����7Ěx��:sh�+>I~����&���&�~I�J���%k=d�>|C=qY*T�B�2u1�5�@�I_Sg�~��>g�gi99?\�uoI�Q�ڜ[��\�.������<~f=?{�4�P���u�������l�����g{�H*��*y�w���Hw7����+'���������a8���%�S+_p�#�}_s����g���m���ݭ#F��i��^���� Jݡ7tZcn�喈sU��5HO��E}��ϝ����Sv�X��u��m�6;MJ}�G��N{��!��/���)i7w��)]"��Aʺ;����&��mZȟQ!�ͽd>�����}\����?!�SZ�~x� ����d�T4�Vn��H)=��u<a������C���O�מ�3�>f!����Ad���4�'�c����Ag��1�5M���wY�5k3���{��Ͽ{�z��J��Ձ�����'�l��o�N0�n�O���O��Ì�$�}̇�q��=g�7�W������X��s�hҔ���O�S>�^�ϐĂ�rȦ$�ZE�'Ɍ�4�Y��Vk�d�����17��K�{�Ci�u��}�����J�ֳl��w�|&"�����m�����yoI���g�Rm
�ɟ�����i%{}�5�i ��PSI8��I�PĂ$��1R�����g�11���ϙ�3����eH,>a~��u�F�}>�o��J��3��yۊr}�O��ϒV9�J�C�+�~a���6��P������$��'��Ry������Vx��)����C��|��:��

q8������?9��O������jھz��y]��>����bt����AC���S��N!���ُ�*>x�7�t�I�<��6��+*o��x���yi�+
�OSN�b�8��y�$��?|&>��xzX˸�}�`���7,�>�|�`t�I��'��{>��!�q{N�SĂ�!�5��s�1�{q�T�!S���k'��q߽�P�%d�ɦq�$�/ư�S�>}��:;��y�{u�ˤ�(��R�q8�_�bL@��H�u������������)8�v���a���g�3�O<�4�^�h��9I�L���1E'Ύ��M����Wiq=8����{(�8�ڊ�)�ٍ!���&& V|�!���5v�����ݚ�&!�^g����$��߹'�u%~O����N!P�k�B���O��Y<���w8�'�?G�M�}�(��Dv�fŞ�^���>d�P�:~�4��*Au��%O|¸͚��C���f��Ă�!�7=��~C
x��4������x �f��s�6�ԩ?!v}�k'�:�fxg���z��uOuuo�=��͔�-�k�[�=�R�)�b�r�h�Y3ǫ���C���l�Ԁ^0Be�J̿��2�Lۭ�9�����8�Or��4�kz$�vtd#Χ)`�Δ����>��,Q�c�bOkZWW�f��A&���N��wj�$���aXW��K��F!�J�įC7�iVJ��y�CYd���<2�$�����eӶC�q7���<H,���ĝ��2|ʬ���Ɉ��b
�10G^(����eO�d19��v��%a��i�g�1�Ou� �?$��~hm �N]�14��T�����|�m�&$�>dێ[I�+�?�����Ps�k��0��z��m��Mz"���<�~��2^R|�M���`"��3i�Oy�4�����0����i�ϐ�y��$Cӝ�P�4��b�{a�b����hJ�
���L�t¤ʫ��3/?!���|�M!P�qլ'�wL���}`c���dՠ~z�~��q��C��?sZ6�:�Tv�M�S~a\~;@������O�i�!���!��H?yu�|���t��߾����$��z�C��t���^��@�T�M�&�Y1'���4�J������c
¾��s�wA�IP>}����J�+%|�!�l����yI�}�8}���p�>����v�����s�T8ÿ}�����7��%t����1�VO����4�y@�g���� q+<��<a�4�&=C���<H*�!�3���!��g��ì�����~�%禅y��j*�,f�^+�@��eg�y��N!S�M���X
M�_w�IS������Md���'�՘�2^Rq�c���LC��i �C���>N!�����m!3�1�uc��5��b���X�?t���AT��0�
�C�1'P��8����wxx�Ԩ|�����&�q
��5��R~��2�]_�<�t�䕕�箓~P1�d�S��4�:�T�s�u�Y�����۟k����w��'�c��������i��Y�|�$u9i�i'���tUI�T?'�3��tCN0�,ם�|�hJ�ٟ�4��ɉ:�-1����te��
¿���oy�$���^'�;�5��D9���1��� �[���ʓ�wI>B�ì1]�~�4��P�g2|�0*g�s�I��bA��5*N>$��1=?f �'�Xk��!�Axɲ��!���Ļ4"a����5j���(5�j��t�g׼�f��#I��+�<��_uU�kڸ9�y���g��\��~��e��MH���q��%�� [�1p��ú4YR�mۮg ��� �3��E+�w(;���ɲ�s=�h��[mu;3�<�x��ݳ�;�of���>#�+�8�ՊH*�SS��I��R�'Y3�I�d�b,�k<~��I:�O�w���OU���ʿ2u1��;N���&r�a��������'z�Wߝ~���~�%w6���� �C���m�� �M�E�:�C�7��Ag��y7O�b�]y��T������0�f���`i�P��{�<N2bN!_Mw'y�X�]az=����5���SG�X�"��2\�I�߲m�++����z�Y��<7��u������I��1���՚k��?&y��YSI��3�?'�c�*��*����0�>��?@���ǝ�q����~�X�g����iYӟ���6��dğ���c
«���$�
����&'�bJ�'(u4�%E�e�N�Y>O2�X
N!S��Ԟe!P��u1񘹊��M0�MZ���0��=����I�s�߾�+'��w"����é�bm� nw���%eg^$��w�Chm �9|�\��1'����2g(~a�ˤ�E��S�o��L|� L)��!���כY8?~��qX
O���H���?~�Aԕ��5M&��g���v��6�U����hI^�~�\@_�?!�����m6�Y�6w�&!���J�	������.���S�{X���J]�v�b���HJ�yA}N��mt��xzE�2I�lzZ����T8[��5{����j����|��@�6��R5�ڷ\>��P���+�f֧�Dw�p����V�@�<v󮕖@�%����N}v�p��pȠ�4��]KU���ϑ���힇��r�eU��yv0�8q\н�Lf��	�j�E��n��s�K��Q�w�|������u�lF��&;3��客]-�r��|�r��� z�_5��=�xщ��U�X���*�5k���o1R���髅x�~�1�z$
cypU8����:ܾ�"	"��:Cg�q�2I]+!&�l�o���fVRI�]�oM�|i��y�uـ�
Cy��B�Hv�M�qA؍�a<dt1{]}�e{���Ν�@ /���k��BS.S���I����kUDC���	���%�@-�&��͡dF�|�� ���dc/��F��.r칂⫦j.���e�Zۺ�ӿ��M�`�H�����Zy��ʅKQ��}\���j�n�D���S�<&y�Z˙�R@�ݢ�=��E�}58[Y�34xr�}�+<Z_N��ůz�qvmݿ&R�,j"�)d]�q �Z6 �/\anA���P�ջa�S��s3\��!�mH���d�.w���B��#f! ����]oF�	�!<����imvqKf���q��*���y{ �y�3����:�<4U�<<���Ui�ɣi��h�ĆGpؑ/E�$��Lӓ� �oԶ�ND'�@\c���T"5�챤I�x�d�縌�0�	�!���V۞�"��@+&��
�2���q�"^}', ]Y�����H������u8��|�xcM׶}n�s��u�dM�/
��1*��SB � w���H�?;�M�^N��ջSR�g�̦�3޵��^����Y�<<-��
�-�+�m���j�%�����ӣ�qN�*���f�Zfnp7��-�}H�5�Oz��;o6�1�v.�+X�'2#)�!��麗J	?n�DZ�/(4�Z���z8eԉ�.f����0��:8��4��ƿc��+��UG5˗T��sh�8H��i�û(8*�k�*B^���8^R]�*�s�����i�y~��#�t����p���_P� SZ��U{ʸi��F��zbA�܀��؍�tO	�)Z�v����N�OWZ�������G�(���P��	�l�zl�0V��fĥ��"[��}���od�������j�Tes�B0s���nC�(w��!=Y�C=`�*�c�݅�4wR��)���d��Eٙ�
T�eV�[}�em%��Y��4�J�F>��m��Ӊz�M�F��ðl֡��j&Wv�k�!��
Q�����h9f����c�bX���obU>ԭ#"�C�ţ"�4p��lr���4Vz�}�$���h,.خ��ӝ5sY&wLi�a�<ޥ���Jytv[��󹝚�c܅:6�"D�W )�"��B@�8w��#~q�����p,��SG 1�H��;$&�q��+�͌�y�#� wb���Lch!)�ڞ-˻�j���t�N!wGE��\D����I\$6��N��O`�yjh$�	kUg����[]��3}��6�b��+�Ǣ���jJ��yj۫r���ŐDtI�W6�\{]o�Wj�Op[kH�j:�Hpt��B�e1����٧,�h���<X�W�IQ2��{�T\���FF�2�n�u&.#Y#�bY��2��:�	�	�j�������YK�m����1��R��lb�����B�p��'b��uJuYN�
&-���c�M��j����Z�V_݁�h�T�wz8�);"�2h�xƄ��We��Et��Q��MX������
����O��j�ŭ������gM��W\�}kk��q�N��!A겅`u�s���h^��mPmnx&��'����w�`GR&�,����A�MF��>�r����4�fCؕ�49�7�JN���
po$w�5�n�ѽͬJ3���M�ग़�""�;�ӫ��#����������0&`�%t�M#�ýT��V��:��ٗ�3�}z�����.���;A�e,��}�E�4���2����!�!2�_�:`��S�W�NNЇ7���Ո��;ۘ��z����])_pX�bR��9Jq�p�ߒ8�vq"�ˤ��kQ�D����t�����6�>�^���,q��ܺ���DA��؞<x���{���P�G��g请֓�Ws���Q��%��W���k�m�.�wt*F���[6ۭ�cxab�5d#��G\=z+���F�u�ckz��]������,��_)LWJ�����2_ﾪ�������w*�����L������6e�� �#���O�Y�]tH�=����t�<���P5\V���プ�Qb�?�͜�́X���U��Q��,|���
�u&��G�:a����$�Cؔ�D�Ó�5Ҙ��x��G�ÕX���R�sý�K�<��o}��>���:�PE��jWb#Y�塪v��62#G�5��-��5�%�[��aKf��l� �r��Uf�l�ѡT9�]nV|�g�n��3�	�����mi�ϩ�5�F孪���s��H90��e�"�t� "#L�-�@��˗Z+#��s�V�]�Zf��^|9�!�P��;M�$a��oMz1^��q�.y���ʚ�䎍�V��j2a�)���������)����C�w�Ƽ6���]Kdl��
ynw4�����!�ߐ���B�)�Ѭ��lm��� ߓ�v�9���X��I끢�2�q�8�f�8�o�yZ�\m>��JZy��Au�>QU��~dו�h@U�c2��O؁v�1�!��[���ttŎqw �r���f7�f�'57y!]\t	��ZmK�(Ҳ�FKy/6�s�m�`���yec�ua*w��U��nr�sQ��#����n�S�ޱ����}�+1D��I�	�����(�F���͊h�K�W���K�u�'f&nǢ�16��,zU�/�<ݞ���j�V�{�#��&N�J=�J��tq��u��%�܊�׫�p�F�[�[��}��X0� W�鏀y�vo&�6��6�i�<��u~����oȯ��t���}-W9�ʤx}]�`��g"���N�iVn`��u9`dk�`��w½�G���x���%��$4{/��Gdc��Z8V��氨H?�(��]�)�#c�C�ξ��)��g�v:��P
L�5z��}SQ��S��T�j�qǲ}�vD)��y+`��N鄁b���q��PHjя��Y[��v���L�)��hg>��h2�UT�U���hl��J�7L��S�m��k4��j�k~��c�BpL�7n��) n����1�t����r�3��=��z���a<��Uc<9	��o!��� (���؋�Ѱy�.�����t��ӵ�q��sR�,��ٴ��
����~R��5��U�^�<�^x�M3���&��nW��A�N9���y�q>�w�4���QT�q�u�u؂Bm>��i��5�"��9]���n���5'Re0T͠���`���T��oDOI�R=�9�!�^����R��hpW�uw�w�������`�
����^N��w��_W�������5�RY����_��+jz2�9Z���h�h��{T����O1��<������a+��ؑ+E����Lۜ��Cim̜��0�>ʻ�)ޞ�ZJ�y��\�N�R��U�eр\t*!�R�/��9�U}�+m#���X��Q.7��N�K7�Uږ'To��`|{aV
��ez/�Ҿqxb,p�F����y�|+�r��[EK^�5߄��޽�@�{��d�1�C���D�:q��ߨ�B�
����ͪ;]w~�w/���h4I���m�˗�5��o�������uY�pȗiȱ� ~^���V+ˮ�ѬU��|�=�g��aL�$��v�f�r�00��$cYEϦ$rƲlՓ�x�< zyz�vw��꓋Ǫ�i5��b�q=�^0#f�����6]aO*:z �	��Xm��U̧=���ۧ�1~���ig�E��ρ/>�E㑛E��brO��g�Y5�6wV��_sh��C��Ɇ�ҨO��U���J����z:ֺc�U�h}���G(��Q�F�緗�n�ST2���G&Sea`�̙�|r���Ӻ�ʵb�v[��y��uI��c��۩��b*q��Q�G�N]O�=�P	}��Y$��Z�5ٓi9E�gu[Y$mVÏ��$����{�z��$�[XTb��ϞjS[����/-���@.���n��@s\�&�W�s]`I�]�sߣ�����f�Nul�[)X��gm�2Yy�5.�N��>:޳p�-Ś���f^��ܥX�dw�L�EH���`�(Q������Eu��^��<�F���; �h��w_<yA�w�>���	���cgi�RS�BzO,�*æ�����ܫ6Uӣ����ۗV���A�m�{v���oo��h��{X�SB�"���L��вDk)_W_!�QYf�r�VB�j���L
6D��쫔T��²�k^�,ȯ/e-*꣏�#���CoP�X\1�%'�H�
���[��� xe���&P�%�����`r��E��8�vm���"��̡G�n��S�T�v��z�Qի4uJꂦG��»�9X:��u�4&طϫuV����BAΖ�9�t��{v�����|=��+zR66�݅.b� D��������֍�gx�<[��������@n�-{��_ZY���6S(;�+���m�QL��}�S!ʺ�`堊\��/x)�jzcKEb</.��ERB��b�}%ҹ8���YQ���h�*g�#M,t��XU3�7�j⦔-�с��p���y|�K`=�r^���.̳|9��'������;&H�f5������l��F�Vĥ�iKNn���Fk�q�`l�J�oK���Dԩ�\WHZ�*Dde2�U�ܻ���U��@Խ�i^�e�*^ܐ��Kz�PyX*�A|���s�l"�N��^c\z���7��� ��,��٥���g�4��0�e��67��m�X"��jn�
�+CB�(T�т�,��7��Fk`@�:��d��b����,0g>�Q�LIN��)�O�x2�z��yrEV��Z��,R���8��6;C�G2_���gBk6���;dTREYA%}J��Q�6ᭌ��}�u�(ج9�h��+en�܁���ռ9����԰.���r�ik��C�e����B���tȠ�e8��D>]���0ʒ�Tz�����r�\�w��|��{(:!Ȟw �.MeN����'j.�Ypf	]������om���d}xoe8����bG�˴++m4��m�K7��f�b[�Jѯ�*J�;��Y�9ma�M=�I�I�əV�+G/�F��k��`��c��J#�h|2�H�ֳ��B��@=/fm{s9���r���3�92�>#x^��ME�.��Ҁ_"J������f����U�Z4�J�1�1I�1��7�*,��8�(+j��M�]}�]U�U���(�X�V1bWC)���-,EdY+*Tm�2��r�Yr��--�QER(��Ă�,�Y��QE�B�VbV@Y�AT���8ԶV�fPkAdr�QE-��$��6хT�["�XH��1�*(Ub�R�X���X�TưS-�ш�Dm%�*�Um��1�T�6�Jʂ[X��#"5
����X(�4p`�3*�A�R�D��kXc��J,�[@cU�h6����e��ZɎJZhF(6��"ʒ��
�J��+*��e`T+c�Y+b�@X("(��*���Z�)[+*,�ڵ*�
�����w1�V�l���7u��]�+�v��]�;�z��'i�B=K1"��Z���݀򱻪�#���g%JN\D��}�F�|�;}��G羚j7"�}��L2U)�C&.��4�R��C�u�N���R����_i�	��L,�'!�:#��|�i* d���J�KX�_mn���:~�q��B���}4���ɞ��<�sf�PQ2� :e�u�Z�=�s�%v��h�]�E�p����Ht7DWxϭ[��R�y�#��#�+�v;���6*�b�w�ނY�2����i1
N��֘���(�1,GL-�g�_�8c��%���z�ݝ�8��H��J���C�^_��lԭ�\2gz!����T<�y$g����� ���k�����3���B�I^+�b=ǥ(��U��O���{_եp��r��ٕ5:w����]2�jUǐq ��jꑨ���x=�i��vϭ��u�.4)�Cd�t�}Ȥyt��峊v�)�G?b��=��;�[����G[V6�M�v����(��iA�f�;h�aƈS�n	f[��wa�6�6Co2�+lh��
p'Z��9�"_�1���q�g�S���o���}������ٖn�SATY���z����K[�gb	�U8��rҔ�5����n���v���O���גs=�ϸ�ft�Ct�n��.w�P���jf�{mfH�ޗò������DD|*�#����f�ez;�e����	�C>�Qi�>�N�@���Z���On�*ȝu%�f��qś� ˝�;u���[s��ٗ�g���p+:W�:���H�n�^���lb�㮹.pk���:i��v]#�^�\*��^�w�L��/.N.�12����V
��*�����V���ٓ��)[XB1HHLU�U�,k<�+����v��Gh�s����������;�27��3�߆��s��Fn �4xw)T��Vy�@��S�S�s�kOT�ifACb(&���OF>��t礕��%`���S4dt�:�h����������}�y\t��c�
�����R��6"za���LXv�������� L0t���'���V� =q�a���A�\=Ƨb#G�]Rz؎���>ّ��/D9׷1�zm��rOn����:'�_+� X:6�s��ܬ|��b9=2C.z���{�25�\]P�N���LU_ϗ[*�ӓ�J�Σ�i��@DF�J]D@�JK�ymEo.�����9��^~VLٟk��� ���YΨKי�����4�b��X�2�́��a&�E�n�lt�걇��s��`��a��ER�(�_d2��Lʸ�n͢syP:M:�5Պ�Oq��H��i��\j���V.�LU��xs�����,'��n�!�0l�+����R����W�Ou��Y��r$a������#��N���ֈ�:aN�3slJ�k�7G�`VC� 7�"���E_�Ŵ3�*�תʾ��[��T��4.�Dv��]��y���Y�
���wk��.�>� �j�wg�׆1ǚ����;r�뮲�9��`�%�������F!��\۸}7�,�s�-��˥�Vq*be`��ȉ����7B��S��C%L��ǰ�Z��3U;�ǹF�����O"n=�i�~Zl�V�++D�V냇�xAaYw�
�ε3�Y�QFmsb�&��[���P�z�P��9�~���ñ�����u���,0��Fb��c@,�s��0��=39y�.~p��!��;���1e��꽸ΪDt�K��R���85�E�GJ�{~qj�$��J�qȽhw�|��C�F|�}�8����j*c��ӻyd��W*FUtˌ+!��T�9�!0���s,����u;b���Y�d~z3�uԺ�1�tO�n$��p&���2��,�;�o������o���%��<�F)Grk_p��md�5Xo��|�{�8��- 1h�7�����q��ק]vb���k�K��k�:+T=�7KZ��/�VLձ��P���ctz���}U_U}쳨 �5�dD���~�ꙅqJf�C�0N�ܺ*�NC#$�,w	�����rB�<�
.�}A��*ߩs/���M��Mp�\;�Y}��O��)d����g�1�ha?8Fip�fu;yH�/�?$* 蔲�؋�ѱ A��E�	���fczl��Ie��;n]:H&�H�����Vn�Ssp��b5�j����`M��o �m�;Gg�=�r;�8!ݨ_�m��/>wp��o�m׽0Nz2�yj2�ᢷ���^7G^��5{�o���O����f�!1�6D����4���Pp�L�O.eWF�v��&�M>htL�
���¦�=�kl���_�]i\2Q�[�leF|�|�=9�jYj���շ������.'��Z/u�-Վ��類�"ゖUXq�ܹ��!݊�wcr�G:v���M�ok��ؑ4��z���8��B����v3���c`w(Kj�1s2�����45�L�6�=�/���{Iv�8��ϯ��6�+�����߽+������H*s�.��>�V��iM����u�5�ż��ޜ4��l���X�..�q���%({gPp�Ow���f���-���:Y�;0�d�:��e,�[k�jk���+�����o�۞�
���_UW�^X}��=e����|�C�GZ���M!3_o*ѦWl�e���R�ذ�b6h���ք�i���w��3��;�y+�Z���r4�{"8�`d����|f�ÑX�f:a�	�����1��ԥ��)j�CG�\N�Y9�Z���S�\�^�!��hQ9:B\�uo�:�gt��޺o7�Wn3�P�+t����TU��}�#����Lt���뒷��>w������^��E"�pm��F7�<~ﮍhB��So�T�i
ѻ���k��M	9���d����)���Z".�}e��^�@�ʲr������}�RV@e
gŘ=�tz���Κ���_�d=�N�N>�r{y��JwP䌠�_H���2�tC׮t��X�F��좃�G !q����ʝ�5:[�}}�x%�v%{����8E4������^��@f�4 �TT������B���Lo'7#�Ҙ��6`�7S�^�A���j׮ڵ��'}�T焀�kE��_�d
�P�g :: �)��'�Ht��;���,�&H�u#9v�� ��T����1�t.�����R�<�c�
���wb�Е�QO�ѡ�w���L���f��<?_@i#w**+C(�Z��9uԎ��;�<+��Фׄ�]�vM�'�U�Ὧy�������ovuu���HP_������7;s���b���{��vVd�ğ��H�9����x�O�����z_���*Gy�l#�ڷ���]!P{������r���
��}��z���'�(�[�?OE-��tm���u�oq��3N	�=%�Ӓ�L)��0=����� ��4�`���Q�cJ��7ŵ��բ�L��Lb+�\�5��?d����d���#�S��9;�{&��d����W]�A�S���^F�_V}�U�j"���{�u|�׽��^}�୏��I��{��n��kO��5a�-�~-1Z��v2#i\�ɸՐ�.
����V�]��ٚl�rn4=3�U�X��e�>픫��Y�ZU����q{�h(0��U[e���u@�g�&\�p�y]<�Y�-FF��C"�d�new����@\:�F�T=�¾���Ik�p4�Ɏ����C�[��Y���b�ǃ�v�~�b��Ɉ�'���Kc�U���p�fBc~�Mg���B9C�rg��:�lLvB���u�.f��I�O��U�z7������x���wn���/��q�gXh0@�C7N6�!�=Ѧ2Ⱥ�p�}G��gw;���Te��Xs�.���%�C��8���j����c��Ž�p���{���&�N�;��Mg��c,m?�v�W�}�}Q-���|Zݙ�U=3�p�/ad*��E�L�=�N[����0�+맏T�^��ޤ�%���6�'p�@g�>�:�˅�\=Ƨ݈����)�B5�VX�Z�\��ȸ3]]�M���^ul��cmPS� $,@�R�b� �tlu+�;���\CӟT㹎����2�����Xq�TZ.	gu$d�P��+�Y㒕*�E���8=fQ=(��x���\�`1�Z��zv�sT�SW���L�׻f�)���{MĀ�3��x��T+P��7����M���<.�r6Z}x��N�c�o t���EF�3res���eܭ�{��c���-�)⾡G��Ȅ��?�yW��Y�{��uK�����$,��1�wCo*�é�'g��Xc����^V�Z��&����w|�%?C�[�&/�1�Z���<^8=�s�l�K׶͘<(���i�\<*�쨬1O����b����z�=�K��Y~oBԺ{���p��o&��#����(A�����E�e����7W��P�V��g�8Sa&쓕ds��ژ��z�/��A���~�����`;����(�����jz�!7�d���j�y�+;��g�c��9�������GiL̨��KH����>���cU���i�] Yٷ������G�65pT�!��-̶�R��듶B[�T�9y�����>���I;��h����hO�y����v�z��sW��Ex�5���/����ܤj1?y;��������M�C��]���6�q�[���j���@�\��YŮ����{}���})�T��>��F�0(���B1AOΡ��O>�1;6�� �t�)Jl'��'��z��;�`8�7�)�)dF�!p�0��y 0td'I��c�3Ywb1��mO����U��.!r;- ��X��ip	��#gG
ߺ۩x�ϞI���h`
�&g+X��u��̴��X#D��u�}��څ1��:&t�����3�_�o����K��R��z�D�r�W�r{�_pI�ߩ�q�ר47��I��rF���=�Q��@p���Vukz��\�Feڜz��|�[pf���$jfԉ��S=7��UR�1p�e��"�b��9�[�:����fN�� P��B�so���7	�����*~���ur1v�D|�N-�i�h�+d�8�� �ԇh��Cc�lD�Zs_wɛ�2Š�[s%�5ݹ���č�_(��T���5ܶ��^*u�mMj潆,�n]l��TH�]��(�\�xSx�bn�z_U�ɖ���,�t�}{Z�m�ɻ[[E�4��j̥�Xn���|���Y�#;�+�5�������>�$4��(Z�w��9P.��i���<��kl��j�`�;r!_ܖ1�(23��w���O^�s��G���}���y�*���{��hvݺ���b88X!n%-��WLƷWW�x�\k@�q;S�	�׺/�頻h��hlϑ�9?���B�����}5C��*{�4�NR�Y�32�җ9
�J��D��n.vr���y2R]�"�]d3����y�m�5���*z_��UXug�qO�'�[��U�L�tl�����l׎s��}8���.�w:�󻕲�6���;�}��i����F��q;�;`8b5��{~�ʧ�QVB��W���%y�c;w�HU�Vr#���`��<9�N�J���A�_
��~Fw��y�x6���P��$2�]ܭ�p�Ǔ?��Ѻ�m/(%�\U����k�����Z�'�c5��.�5�rk�uC����u��n��^�C��ЭB��S��Mf�7�2F����W� �oKF�.x�f��;���>�\#>n��B��+B��S�}��
���>�d�������j���MA|lPxhҗʦ[��β���q��7§<���[]�v���<2�MVo��YP���:��9�.������c��Zx�kmc�jr�A	��l��]w��t��}5x*g��}x��_�pT#���Rm�W��aQf�}�w'd$�n�#���G�}��dκ-1��up�(>�D|����%;�9���qy2g#^\9�+�v�4�N� ��e�,�_2�?�W�<��������H��;$&�!�~�a׮tcl����2����Qo��TE�zѡ�}QR�����m� ��3����dWZc��3s��`������k;��oȁ+�h�B�� TE��;8�D)ԝ����+T2"���������j��Uo���y'Q�;c����T��/[|�3�L����u��"^_k~�E�*~�q��ġ/�P�2�>b�O�ӛ22*��V\#�m��v7 ����lj8�IY��0�S��VM��B��j�}Ù7�_U�*�=ׂ
�:�YSWծ��9<���M��뇛��30;�ۄ�%��v�N@3��CWp�OX�xx�q�*����y����2s�Ul�F}B<#��c��X�J8�~Ԯ��z�+���|���A].j�����)j7�v���0��I���[�r����ve��zx��^>�y^<|�M!����u��ל8<Wm�@�Ő�Q��W��4��j䶂�P��Nh�,���$K�L���ba����h�6��sv�2��d��,��Bk�m��g�wMRz�b��!w����X�Ƶ�r� ܉�ї [�H.k
�엿����� U�/����J��B��!��X��ku4�L���W`�X�����B�P�*Tv��bo2��$�8�ufR�L�@�^�١)Y8�pf�W՘d��l��/���2��0nSB,ր�Ex0�J������:;G0娩Mmκ���+C{2<��W78�z�SQc����V�}��z'Crƫ��uڊV��ú�k2�}�Q�4vҺ̭{BV�2���Ӣ��.L4�HH�	�����IOqr��V��o�Ts+q�0[0���x9�s#�zC��[Thf-*�6"�gtK���嚬cz"�B�l�J擘Gv=�"���kr[І.<��b�n�Ȫ����2Vd�R�o��ptz� /�T��>A�WK�j27)�Z�o����^7�1��T�}O����;��:h�O�^	SE]gL�����{Uf�b9A�w9jkR9�3���v��r2�?��$�մ���x��C郷)9�:�sh�'XNX�-Z�gD)
]j��:V��!U�v��T�w����<��P�@�|+M]���.��%�N-�vCe����ڮ�L�E9O켼ʝ������s�l-HgP��*#����zx��]XUř8����j�$d�ؠ�xrL\ef��YٲQ�N_9���-6x����$�t�Zv��o[³E��H�d�����l<�����
�7�;^z���{\|j;<��c��Ǯ�p�;g|�N�[�5�i�)p��1���\�s��&ˑ��l�vTW��p�ǫ�J�iN����0ړB���>�S�#���:Û�*������w= .��]�\9�@�em���
B��o�f*˒��-�˝�5K��F�xT�_�I���Ts!%#�Wn�O`�v��Vr�r��ھA�P�S��K+(���=�fd��E� �FIJ�|�tlf�.����XQ�j]�����'Ka�moy9�� ���t�V��:æi�!u!�"Q�#����yv���mܝ��60d6G`���$���h
ˠq0#�2p�3+���I�Ivv-��'��u6]�aD/�;�{����5������b�8?e=�;@���
�5jq�;�PT��l��3��R�s)]1K�`���Nrh�ɗl�tsc�;�	P�]�y����O
��,��qj;�@=���CwB~�k)��{j`]�zNm��M������\Y�I�(��ӗuǫ�����U�ye�=[X%�U���d�DU��(���"��.-�	(,PX�2���
�TQc["�
���T�`��6�Fҫ-�KZ�i�J	�R-k�V�*DTPTDR�dR�6ƅ�e��#1V"�Y�Q�e�5�T��B�A+PR�Q�
���Z�Db�e�-�DE`�Q��mQU�Z"Ȍ�m*��()#VF�	U���F0B�Z��b1���lD��b���(ŶR�T���D-JQU-��B�U�AH��*��ŕ*+im
�",QEhʨ���`�mQU,E1F�J*�QZ�QUF*J���dTTUQ�Y|�_�~޳~5	�C���u+V-v&�c�����G:�\o 4�l����wj�M�x��N���\���{�U_UU}�%ڪ�m飣$~���U�ȳ���4�v_��l�\"��vxKJ�� jJ
�6���k�Ƹ���9<�s7i����'�d�G��I��FLp��6���܄�璛�Nk4'w���ݐ6]������t�:S�!^��9�͙;�TE�)T��Ƴ�b�n�7�����뎙�!-��ÊMg��!1AJ��;魱1�u��|$�����v�<W��(΀��xS�
>U ���k�N��{A��J`��� ��\ۗ�Ԧ��%ef_��Z<m�)�0�..�q�3���zj�z��wx���O�����9���y��
��Tl�a_�e�
w� �p |���O���^��=|���@]9��x�$�U��.�!V�!�md�U����G��T�}WT�Y��h���n�֭ZHF��2���
r���������y����9����UL����=2�;`'�rގz�!�jՌ��{���1��q3xƆ�f;���i��7����ľ.I`LR͞��r͙F����q�;N��pT�A�"�)q�7��X�ٌ��Cԇ&ȣW��fv�8��P.Ү�񴎀^,QnL4�:���i�d^pZ����̙]Z8;xu��l���H�]�\��s3�;L�f�{�PU��2��[G�R�@\�¥~�">��,�9w�m��b�w�+��1�9�8=���r�����b�f�[A��N��ٗܪ����`̩�$�l�1����'6�V1�?m)�Udҗ�'��dAu�L���	wWͳ7�6� �ݧ�Z�uw4:��V�AgCWg�V���V}J��﮸NwWyy��''-��{v�����K�U��cj�1s��p���g�֋uJ�pT>��'f�b����\vބXu�\=h�T�����6�	�O�LN}_Og��>��U�`_�[���F���$�n3����������u?Q�h"�<js2���z�r��ׂ=�͌bʺ�b��eR:e�cd�j���F�u��J�ҝ�
#�C�������W��w7y�[Y����s�,Y����<4�� ���]*�.5�/�w�\�lއ'E�I��N�z7�ټf�a֏}�W���_�Ϫ�KX��4����}u��w/ƽ�?y�s��)\P-��98�09gx�R����b�VJ�\�8�͔��kF�wǳ��ݞ�AS��&O�������K�6
۬�N��t��䫮����V���c4U�:g���!s�mAcd=�l�bΣa��K/U���D�$���!a�M^R/�=�q<�J������]C0���[4we8_l1�r�ow��}G�kG��h��&;�H��x��@s3�	��x6���'�|ĥ�]�{��X2J*P�[ܴ{��`A���[pf���$l&m��zn]���팅,F�
w��JӺ��z	f#�p�\���z7�څ�崮,û�ĵ�d$�f*ٱ74bf��}��1̬9�~�K&Ɗ8o����,��wh����֙�s�b���=�;y���e��/�ˀ9�@ieW���G§���?*�W����ԜZ��Ͷ��l���VwXچ�|�Ȯ���%����7H֌)Wmպ��/�q*vDѤ�a=,�kٞg��dٜ�{\'��ʟ��#N�����?h8:~ǿ{h�B� 1ê�߳\u=�1�aP��ypff��R���֨U�:at��#�D�Nc=;����Nޘ���~ߊ�W����]�ړ�yW8�i�1 �yb/{G���9kG8��/��fQHh��pȭ�h�f�j�{��*����U�珀?Z��2�����P���zaWb��:U6J�JW��o�ֽ�}���H ��^p�S	�v��P�g�Wr9���8z�	�C��4�����B�WV��gIC��'RK�������S��^Γ���l�������=�����_UUU|���o��y��~x���xഁ�;�e��W�wUS�<�P��_f�'�DN�9�OB#j+�l�N����zYҿ���g�T�].PK���Ä&��j�G�� �'��e���ޭ�L^HH|�V��ȁ]Q��������t� ��� ��&Y◸��.~�m�cz�䣒����.%n.�R��k60J�cd�i ����T����B<~ŏ)�iG���y���!p�/���󏙇�)�)}!�i�y3�i�Ü�[a�MwVX�(�Z�:�t;���Ӏ���� �dnR!���@B�0$��N���$/)��4��UZ�޷}��US/��P o�EG�:��Ty{MA\6̐z��Ȭ��1e<��ȴw�~�{��4�1﷐��W��s|��h�Fܲ�rv��2�:�gt��\��[�{ݏ��C���ڎ�P��uT� 珤���3�=Ǣ��E�iS�t�ہ}�8�S�����	Ry�jy����[5r�mɗp�����6deS!�;]��ݹ\��#�V���OP�.��v=立GP\�����̻0���=!����>���Zm��9��2M����w "��C-�yX�S� �/{m\=3�b���Ϲ��a����TіV*ˤ��y)�4���|2��p���(�Ҙ,���pt�_g��ﾈ�f8�g����Ja�A�;7dۓ"a�zne�̔%�pGM����il�Xն��v>�s���}k*JOz	t�Y]�%��t������i�̄��bᯢ�@���a��Yjx��j�}T�h[����ZǊV�)o]S�W�z}�O8�Ã��N���mWp�����W�q]����xh���(V�^���i�2m	��,bT��y��8�d��xXv;�ؕ<���@1[P]�7]z
��G5��+���"]�!2��r�h�H�<&o���'~f��L�T�FB��9�-m�#2A!}B2c����(�Y���� W阘5X�~�W0QiX�����Żrq^��-�ў1�4hIo�u϶(��9i�=wۃ>�b�\h	,,]�	��Mg���G'NL�+'��a�ޘ�}�S���5$dI�z� ��V���.�:�v��
"i��r�v�؞�rxq�.s&4���!�u��Q���3���Q�l~�3˅q��b#]ӁT%����E�6h�m��o�)V�k��<9�Unu�O74��R�`��1Ǝx,��9�a�K��<f�dW;���hK�|�ث�h9v(�F��`�!q5����!j*��/�29kW>6˴:K�9�q=�N��.�H� �����W�M\����興͹��.1��!��vX�u�M�0��t�J@� |�`��
��8Kz+�g����{KY6nO?k�\��O��[ΦKڹ�6қ���7�������E�s�'M�YɧF�d�&x�����ݤ���K���fQ׻rCf8G�L�t�.|�Dΐ�ME[w�3�9��.��)��m^PlL�0�̛��`��u竟\�Z
[IZ�&%��{b�sٴ%v;��pv2�鲪f6�<3��̴*l�?�5�i��cl���wEp�1�_�������\0��WN��3�ہ�.[)ҳZ��{�J�SIE�UC2�ƌ�zbe`������
Hq
�������W��4�W�r)9K�y�`��5}�f5�e\޷�8F|X[�R5����pu��C�fMZ!�~鶍�����A�s0��LɚN��}lP��b���D�X����zϺX�.D��Nޗg=���s��8~�*k��5��.��v[���~��|��U����42�
Oz^�{Է
Zm���u�6}c'vqˉ6�<K}�n���Tk	A1qްl�p�M��un\8�-��5�{�����:>��ݕ!x�,hf��"Y(�꾹��!�6e�}J;ڇUp/�8G�jՉ�_�������Z��W&P��N����^�ϯk��J��O@�����?t
T�Z�(>P�^����OF�u���X�AQ<4�S7��-�B�j�L��:
ù��o�GBN8���:�v���Dnr��v$���.o�Kl=��nsxT�8�s����h�a���oj�cQrs�*��Q����2�%����'%q\:ӄ�U���i3'tƸڄ�!xq�뺝wR��h�.����/QQ�"�{�3AOw��5��j�T�ęR�sz!M����_bwz�2�nJ,�1�8�W�Q��J;�Sl�p듇�%��;=���sYZ��ۧ���vv\�glCufiv��J{���Ny>�U*��5�\��]ћ%�b�hp	�y�*!93Ao_��^9U����}�-H������Ϋ�ƒŪ4N�ޛ��3�d;��^��}��/�\��7(]&�-��#G�ʹ�D�ܻ�]���ݷ��b�|�U��:�d�h>#�nC�j��v�=X����7�]�r�߂�TU���.�ss�.���:�x���N����4e�����|0��>�����u���sz��|�+���ne6`���C��̜�٣Kd^�\�N���v���ר	�}"���A6�bWI���������=�H��c;_d��z6���+�&9e�.w��ގ���Ϣި8�o��́�J�3�湪]�F Z�[p;�5�=���j�v���-���w:ܢ�`:�\���	�ޣU����8�ڬ�Ë��Y�ju��Xe����W��{T�ީ|Z�ִ��k�7�M����(�^N��w�����3|��g:7���>M3��Vv���`�> (�Q�b$VL��ؼ��UӨ�����e��>�;����y�ݜxM�uvnji]�dpꌮ<_>������+���Z�IKY��SI�8cjt�,�n0���6�s����'�)�BwN�#;�"�t�]�B�NBrJ�b���bm��v9wLP"�Ŭf�̃^�VH�m>r���ҿ��6��B0+���Z�����A�����W_���]�)�x���h��uy���-�U�{u�tɵ$#v��M�����m�k����k6pP<�9˹\���EB"M�S��a?]����荭=�[�ܷu��ИA|���Y��S9�J;��_c*F;RN��e�d�ζ�u�u��N�9�s�Z�!#���""�=Ȗwb6�XP��;.��GW,W�sۇi��yἘ�NL�Gf�n9�sֳ�����iq�cl��YE\�S�0�C9�M|�d|ӓ7����˗֫$�v!j��ݚ�����p�Z��\��.�\&�����!�p̋�us��{\�R�[������'O������fm�|���Y��M�b}{�*�iI������x5�5����y����.3�W�m��n�ҳъ1��O��'=P�:������;cV\ei��[k�zj��7V�֜��M�Aڶ����<���x��#��z����,g>����8j��t��Y�����r)�cNA*�7{��y�\[���g�\�nM���c��8�o�n�!5��c��8�:�i8p�j6�Eғ�6����x�
��Tq�u$xP}Z�LM��Qv+�=cL�\h�u�cU�<-�wIk����b9�n�V
��|��s��f$��軑M�j�8cs�l��8lͼ��i��WQK*�\�;�ﾈ�5��@�a�/D.�����;ot���.�ͫ��{<mw̰���zl�ٝ��ѡ���1�W5x
Y�<��������}�IP)��D�<�_mp���5c�Q�RNn0�ivR�L��'�;϶�����e^��ŭ�R6�.3��<o>���aQ�b�TJFn15�����(�:��x�����u�C2ydk��yig�ư�鄪&DdIg$Z��1w�	׋Iz��/�w�w<��M�Z�Q�|��ݶ+|q��TRB=`N��	�/U�R�O�r$�����H���y�Iϛ�X�v�0g.BW�{u(y�m�X�'y1��2)v��}�VtANz���ǲ���F
�	R-ݠ,�ҳq	q�\�@'n Z�͓QoF�u��ʹ������/E��Q[�,�]�rf����!Ws�����q���X�["�'Q	��y=����*u�`yV��!�S��]��{C�:& �|�\����e
/zO���7�l][����bn��%,�/�Bк䄽�Z����}��]g�X���������i)4iP˕Ӫpx�L���620��k�������{�q�nj���
W��46�T�����S���tY����ܻMP&�z��y��yPI�6�M%ތ>4U��R�gb0���
�73��(_*�1��W���Wgs�mj
��_�Xһ��wT�j��"��$m��#��V	`�p�����r�0�]�MKHm�dKW�JR2z�D;"�)��c���v��B��5y֒��.���w�t���N�#��:a��ֳ���v^�hI��#�32gu�"���y:Z�7�؝�*Z�i�� �f�'qkc��÷��7��^��+���(k����yml�r;ć��DΎc�U�t������J�w9V/2����w��8KtC���u�ͺer����D��ev��d�<�+UU����	�+e�x�E����)n�$�=yC�S�$�Z�T V�����mQWE�ΒN'��B���K�LxƩ5��N��;m�LhUygw�T��%����P�[EڮS[�:!ن� ��01�� $�]e�B����(D/9�N'���#Z�Z�&��lP錼'��a�h�l����+{U��@��vZ��U�w�-��c�;�YW�{�!�I9]*�.�T1�S)�ps�Uc�u�=��ݰ�#��3z�[��4W`�gg0ڃ��gn�C����:�I�&Wi�Q�ź�|�̾{ʹVgpλ3S�B�$�  �
�k;q���#GۼN�W0���
 �veB���V�79V����.�D��%`��׃(r��kk!wv�vE���9���%�2֥�Ϋ�	'S2�k��
�Y;~N]X�=y���1�)�����[yYw_�K���i�ʺsB�JU1��0��o�T#H A���c�����5Bŭ��I��k�['[
��re���*���<��fڡ31텋7n2��f�W�h�p*Sa�����e��ʠ��
��DUA��uɼհ�{dv^�70E'J�mc԰P˛���Ze�h)�Dj�;7)�iU�n㜥v��an��^ì��.����y�^��w`|���H�o�^m�b�f�uW<pɐ�����f��7�WG�vTc:V�VJqN&M��vNzk�������]_������۵X������4��cOQ�v������U{�͘0P ��k��k#ƬW��D�&��*6����y�����p�&]���7�wS��|8;�r	C��|�+��ʍ,˺�{�n��\\��ǹ���c�O067jުl���9x�u�=��-�6.� ��8u���κU|��f�<3B�G3�-��tJH�W,\�΄���	�	]Ղ���V�����2f���u�������V�"%B��*��`�*>ڊ"� ��V
�E�������#2Ѭ��"*5%F*-��YX�h�UKlb�[
����X"*"��)iEQ[b�bV�F�DTDb�bX�*����"��lF1AX"�-�b��)m��Z�Ŗ�LB��p�* ���U����$E��ڢ��X���k*)m���"���JR� ����E�*(�(�H�EF�E��
+Q��(������-��T���Q�k*�R*�,�#��E��*#j�dEU��Ub
(��mDb(���J�����EDPETdX�U���EA�-��l3(<.�>�ݍ�i�u+�=�Į�?�$����I��(��q��h�0�%��5+}9��%Л�N�����9I0ɹ�G�O~d����#z�.���m�җmQX���4[��6��'Նc���d?���4F>���di׽b�xe��m�}$�Z�L,"�mۻ"�\�K�Ǫ��[�1���(�)��-ws�5зv������z�,<U�eΛ&�Ë����<�&�M��Kr
F���-U,�YV-���$f�Z�{`���%Xm^v1�Y��{��dkL��UW"��.Ett�s�!f�E$��vD�N}��=��E�Y%<T[;���ϓ��kiX��g�>$.Ǐ���;m�\���9��s
:�����v������
��p6{��C��^�}p�xjZ�U��L��z�/���M��H��E>��5����=�w�'pF0�&
�ڋ�1��z5�s��0Y�(��E���	�Tɟw�GK�b���=�����0���*�U{��.���Wi��q4{"��t�ӈ��$&�����(R�{'����2�R�m
�RoJ�$�T�e��[X��ѥF��d2�,��Z= �ZԮ�˪�=<��dQ���(�.�R�VK�bӸ.���sF�q�T)�}��o(U������Y�\��?I�CL>NΔ-�ⷥ�{MNh
�5u��F�v�[�c����	ՙR�ܔ�L���!s&ʽ��c��P ��I�F@y�ȫNL�Q^sG��U��r����nkX��*��7O�G�^i�����Pݺ{q��{��~�h���n�L�2mb�}K�YH��mH��*�*��Au*�P9׺ߧB���{/�1�,z�| ث�>}�1�=ڮ3_\s��(�o>6�Q��NB���U�}eLEg7鮗痹���Tc�+�˼��_VEj
ó�Υw��N������h���N텊�jˌ�8�tw(�\g}��3��㣪wv�r��J�vӋL��	J[ʒ�������qv��k�v��4��1,��ՙ���F�/�GssoS�՝���g��d�ad�Q\�^T�zWAt*U�J5�++s���P�ǫ�f�m�n�{��A��:��Krh����~�w�ű��)�ِu�+���Id;��d'mfIoT�ґ�;����%B��
�9b��)E�t0E�H�ݙ�¦��
Sw���c7�9(Ɛ�$�Fq��}�X�M�͔�z���K��ֶ�Mv���+���Yؓ/�M�}Ng���� ��Z�C�wE^�gl���y��J�m��U��d�:kk�9���gq%،_8�n+��3e�;<�c璓o{�q�2����C�����yS���q��L5_N�W�:����؋܅�j-/�L������{�u>�"B��m[�.��oJ��&n�?N�b�j�k���l��F)I�.��{�����rV��W�j�!�G�Auf�<��ޞ흞WY{Y:k��3�s��9E2�6��x���w;j�3��׀j8��c
�mU��O#��>��W:S�e�}�
�y5sM92J�������Yy��߸�;��w�k[E/a��u-,�R�����sq��M-].H�fGN���J]�Ρ.-L����ie�ʩ~ǝ��w�}�zo�ﮈgCgK��w���ow�����mu����Y5䔎�Vd���i�$z��M]r�_@�9�����I�j|�gN�L,�����#q���%b�jR�Z���}G���l/�6a�0Y<V3�D�.�)Ws���k�0늡VAY�D+�����/J���j�s�ۗ��r��Kpym�yq�w�[q��,���cF[�H���4�t��	���U�:���t���;:�c+M�@Z׻�<�i�۸���E�j��iͽ�ӟ7�s�.l���ȥ�1��j��4ޛ��9�F��p���Ks�B�{�����5oI��af[���"���[���So���k'_�84��KTkL��f�a�m)}7�Ty��>�[XೢJj��t�����H�e��7�YM,��u�=)�ţ|�eM�ݽN'��_������)2�_#nCTAv;`�7G�4e�ֺ�;o�K"a*��7�:���&�8K+k(N>�'p����5p��Q���:.�9W0UL%D��wgZ��78�w)�.$���OR�u��'�Vk�W�&�R�tf���D��ZZ��k����@��cU��|�[]S��:�^}�æ�wg�N{�=x6-���
A�d6��H��tMފ�N�qT�F$,�f7i�O ��o%��*!V���3�"�ӕ�>�4Ӻ�E�S���{p�B�Z�YS��P�MwE΂�P���ο�D}��z��7�1��̊)�D���Bw�i��X�藎VCp�&�L�E��7<�îR�F�������s3��""�m^�݄-)��f�D��pI[W�p,�8�޼�1o�յ&l#��*�cU?YR�<��֫y����7'�{w��;]���%(E�SP�dCNN�z�Z9��5��[ �Fm9���5���ݱ��If�e�)Ao��x�p��w5���f����=nf��"����*�ũ�g!>��ҧa�����y7o�s�q�_L���5f�o��s��}��3ko\k��vӜO��k���˕�u#��4o�Vݩ�~�k�l�x��Z�]ƨ�h������ۅr�C�)�?bL��%x��s�D�[C���'���6���N4j5���T�x����u�J3��9i^kk3�x��4����ʈ��\�����rjۼ��e�(F��yf穃|���-u7����7-�w2H���c�r�(!X�������vX�o�:U��hSr(ր�őWn�G�>N�	������NИ*�V=��|��+�d��=�r!�L���cN�.�19�&f�G�}N	8�����߾���6;�Tb/��4�Kt��:�c����7pg�����z8�>/v3Zne�D��>}(�6�����9+{�
�"z8�̌�B�%��̋V1!;��^ӝݛ���.�Q�-������K���9����b ��tr�g�J+\K��ꤳ�(��H�g�L����V' ��6��g79�T�����n��u�W]�fg����D��iS^J}�_'�tW�?�Ǹ�b���/g�j� fQلՙE.�ϥ=�+6����F�[���:�*v��u4�����y�����]x�TY���$�L�c�CD#���Aۂ�u'5�6���,�r�f�rw 3��o���<�Q�B)�%s��P�{ �g���0��t1�r�D��A���#��knI��X)�R�y�n3__>�z��m�R����T7�Ok'��*n�Lc�hl�8:O'�	o�E�����:51Յv1�7��I���}z!Hd�W<��jB	W4Z���/!]�t���建�Co'ҳO>���U���BЌ��[��'�K�w��!s;�Wh��f�م�U��ۗ?}uy�8s�ʓ�Ҳ�;p5e��y����}B�ޭN>��|N�;�v�<×ޛw�Ԛc},�}��>ڠ���7�,��v���S�]��QF���j�@a�}m��I����V�������죋������d߽��b�~��n����aOU��Y��{.I�'�)A�.���t<s��%W|���y�V�y��k"45��ڞ2�ߛ�gbJ��0�&����:OǺ˞O�^�R�[6v����ƛ�y��7����6*���An+U9�(�)�U9���Z�I�c�	��K<����3��!Eu�������k&�����BFwu��q�D�xF��q��b 3�'�c��\&�Oxv���L,�+�%_Y���dJ;��۹�î8�%��Ԗ]s����
�<��%��cLU�1E�.��NU-|��gm��q�P���0o�^��h�^�}�ls�/������]����t�uܳX�A���J(��i�Ȓ؝��|���X��3jV�%`�x��4��-{�F�Z�ۏ0i��ۚ~Ӈ�%��MESj������oӽ�wq����A4�>M���D�ld@/ad1yh0f���U�*�iظ��&���H����=ވ!m�W;pS�C���^�D,���Q��)�^ZV�*{�_�������7V>�����nerj�u��[�׃:�\	�9�bYsp�2��m�~+�i󱚻�]���ů)������ݽ��Ν�	N�yk$���in@kg]�{]�����![��ٍ���þ̥\�Rt�?���Ȧ�Q�q�W/z	��l�m����猉Z���:�=W�\U8F5^r�Ҝ������M/��k?e� �X�ޔ�Vŭ�Fh+q՛q�M�Q�>�]�.nn>z�v�,D�;ό�Q}��Q,�e�\�S��9=t�}���5\�#Mn���L��f�����s�l+h��8��i��F�2������,]i����������)��!�`�ߙ'0'yX^ݎ�<�[�T@+74|�dJ��"������D<��&��+]�Ӏuk6%�G���Y*5���+�6#�I����+�����-�==`v�-k��+����t���;)><�`�U֕�ad�^p�f�}�-�`e��I^��7�W��R�P@��qJ)';R����T�/#�)�;�ﬦ9Z��z�1�]q�xF�Y��U����U������ˑ�ƚ歎5���Ob���x\�fN��6�yid1�,�a*�a.��qw��c8s�]�s��$������5̤�^t�	����h�s�[$uv���¦�u6Q��LFmE�|�"Q��!;m#��y/������N8�J��1�u�0�����;q[���m^jd�J�)˴��ɨWώv�v��bi5Q��r��h�/�>�e�9cU?Y��]�+�lZ�p���֔`�x�n�5�Nб59;�������X:����������=�j2�(ݧbh��}��K����V\v��1Ѳ�W�%%��/yd��/�f%!޸�����gZ���um���9��j'���v��l[y^¼�n9ID�<�u
�K|���y���uMŃ���*V�
�:�k��I���4{m։���R��K��Z��%{������љ9�8�&�\W�d�F��o��K���wT�S1Wi�.*`���1tɜ�3�U��Ș�7ﾈ�X⹶(�^��.1s����Tk�Q�t�s�����󃘫n�vs��W%�/R�j��m��C���ݪ]K��-������j���|_T�C�1�ި�f�Esj���q�#�6�v��pU�W��[r�r0�V���7P��.��\#��2u|�g�Ğ��3��(�\`)�
��f���h¾Hq�`�9�-��&��/��r�v$�G3��q������QHv��\]��e4�_O3���Ȃ���7�D���P��������t���\���QHLgh���MZ|i&d�k��N۹��B��Jlh�ml��`��(��E�B�+VC&�4eN�o�s�;�K�q�Z�G>��i�"a���}f����o�F�����ֻ��@I�\3�>ƺ&�8��N|���sH!�+�|k����.��]���b��b�5��E�d땐����TM|U�г��CS��ua��C�M���aZ�gZt ��,")Ǳ)�Cw��� s;�MZi]��B�(,W1���ʻ��;T�=��^VK�d�=��*��3�,X|;t!�t�unV&���u��{�+�ϻ-\]z�f�r�� �3q���c�
ᐲb��G5Ot
��)������͝$���A�Y�Ng"��7o��Rw�T�ZF#]�B��	F�gk"��dDY��B��� �Y\�����֪�w\�r�f������c]ֽ��l̨�I__]�8��v"ņ�6���v�2O`�VV`4p��@lx�Z(Wj���o�˨J@��W��o� #ۨ
ef��˨�u�_N.Xv�0PȐξAKԅ{q�# �"�Y��ⶲ�pॺ_f��Z4q.̵�����Y��U w��W՘v�b�Ct+n銧��3�O��jvt�/o��F��!m�8�ݗ��\����D��預��i�SAW:�O/A��c+~�c�H&�%>���̮#� �z�k��gZ}tʤ7P���f���Y�]���G�չ���|���8	9�*98��/+f"�[X�١�3kV%�73"i�'���u$�ˋ�+��)@h][0�-=���S���8��Ջ˹���u^�v���1*�ڜ��*�X���y�t�ɬ=�ň��[�#�(�XsS�6����ʾ�*�4�Oqq�x��$H�vТ�z�RM�g��܉����V���{.��m�U�X���&u����Kŕ+�Wj��-.���h�T���q"��8h|:�/�Euh�Q}�Y�6+�Tޡ�*��H85>�o����5�-����v�����$�=��R�շƜR�Q�Ŵ{�r��Q�jCuo9�{��*[�m��fX�J�HpI���J��B���mD�f�,���޷�6��#.ϵnQ|et<��ǩ]�FR�kjS����u�@vӜ�uY�m˨1��̩��TgR��[�a�V�=������6�4e���p��t���2�&W%�A�wC�W�Ev���ZV��lp�����QQ2�>�۽l4,��)��]�:m v��wK��c�4J�"��R��t8J���+l��:K����r������H�R%��PbJ��.yi]�jV=6&�%��u=h��Z�f�B��ph����`���S��r��8�7ە�C���2����2=60��RI�Yu}KhG��?hT�ƆkvN�u�m�
H��-;�7�Z�{JC�X�e�࣪�Z���d�xiWɩJ��y�� \�w/�v�*�&��ܬ�v$,m�|;8�]*����$�{����Ƿ�G��mꬶ%?��_V�o��p��m�k���z�\�Z��0uٽo��g�7V�<�E��]۴F_a/�˥v��;#B����B��G�M0�ڻk�̹vz�.[��+b}imD��QQDDF1��UDb+"�����DR#R���U
�FT�"�R������TUKK���%j
ZV
��X#l,DU)�X��Er�AH�"��V&%�"�������TQQ�QE�**�TU�4W-&0�Qf%F�EU-DH��#�TT�UV(�Ġ�"��������ʗ-)X��DDDX1QQf�q���­j�X��UE+EE"��U��P+L��T1Q�PUFV���"��+X�0X��R
�(����� �V�ڪ�c
����U�"Ŗ¢("%�����X�L�&*�Lj
*��MZD~�˾���*�t��Eu�K��ҹ��m��,�FLV;�����N쫆:��:���Y�S���UT7�F�Mv~����O�U��;g�b3�%�-0~���-93+��-u��VK�X�����"���kHh�p�>2���_$���mC9d;�s-99��jY���nu_ I|�M��o�y{h���dA���]�R�!�QGӿ�"rzn��қSI��Q�9N=������_\O>�q�6�!/�����ɐ�k�g���z3�&�o������Q��+�.�_V�Y�F�{��QS�d[~���qKjKhq���N)��v�F��k��f;N�<��'��\�E�ƽm�YY�6�vG>��s��d��u����Xkqm�O[�I1�8��{�77S�W������9rO@Y<+�v��ɷZx�P�����JE���F�k��uŷJ��7��wTV�+���ͩ�ܔ�b��l\Q��*��;e�e쵏�һ�{B._|�ܕ�WouL֍uI�&M��|�K��Ha���d�)�}~*t��W�d܅���ƣ�s���8��];�v���;��%�'s���.��N+�l��\��8�̄_p�P�?��T�Z;��Q̝�(��Zj;��s�M��ӟ!�r�:���������/iV2�����uÇQ��b�����n��c����"U4��pU��qb�|U)�����I��K�`��H1�JFn1�����#9Իg:�發��Q��G�CrJϣ\m�C[��o|!+#"S9U��83c)3v��xs�t���yT��M�Δa8.��D$O@��ĵ;�v`|1t�X��ݹ)���&��f�}/A��j�0e8x����c�/���Q;�k��_Ԏַ�eb%d�|��qCw�o`8IU᜹�;j��f���\R�s<�E����c�Q�]"����X�5�Tn���W*u!b����/+����^O/�]�W���_^�ڃp8`��s��s����\���k�i\I����܀�λ�����ӛ��tl�V:� r����h8IE}����Q�.:�gSy9�\��gn�c�k]+5k�
��;���bR�ݳ"TC�bN�Һ�[ק��̜�F4��t�#��	u��v��R�ձ	A�X0�d�Z���o�ww.�## e�#��pY���U!-����H�hp�xm@�g�]��JK�A��Lν�}���b��:�I�����L����.���R�0��]f����!s������5�k�q�S�[��)��/�=�;�[E�uݘv[�J�V�FV���uF%εB��ާݰ���=�զH�n�;�v�:�3S�d�*綛�6�up��@�9��%��|���+m��d������M���iP5.)@�j�K!u������c�[�ɄiP�iԮ�Vu��VVD��D���(���K�}�5�P���h��ܘ�;JI�M���u����ύBW0�};n)֬�\�TY���t���g�����t�}����3'�F��yic�ȘK���m,�z������J0S��9;�]�\�Ԩ��reK߻y^<��I 7��{m��*��.�UE�K��F�{�%:l�,�?K�'��ݞ~�Lkзū��ِ?:��+�o�VsX��89mT�[�B͞
mܵ����V��s�+�m��ۯ]�2���UӶ 'T'�#|R�@b�����1�3���ũ��\��!��O3_X�1�����d�b*u4���gcyu����T���@�fmLCf�Fs�|�7#Lq���|�&�93a��k��͓_[�Q�]^���DN��#qű�+6��f{��v:�۸��3�;�,M4��@G�Z7�n���@�eE����K<F�����DR�(m��������#��q-��kuE��+/�S}��koS�Q�	�l�u�N�������F������u*ɣ&8�ڛ�5��z�mmƨ�g(�;i�|�#-n��{sz��x�cO���z72s��ݿ��CYą��u.ޘ���|J���~�q�o���W.�y�;�i�ȳe}�Ή����؞Tf������z��x���kKGv�Gs}�>��z����=$�lQ����9�ʦ�A��ou�Uv��J����܍M4�"�uZ�X�����s[m����ri�u��oyN�V��>��*��w2��-nC�G����V�����u5[t�TI�z�gy[.z��c��ý�e�R�@JK��>�����J�!��o����:�gB��nsr	h�	��]������ø��כ!�c��rĺޤf=Y]���e��Ex{jug���|W��c�%��VX;�c�6d����;ቾ�c;�.���>�E�]$�L�%��q��f��
��$��[����{[*��*�v�5Q%�Ȕ^.�aa4�'¶.����ۧ�iv(T�Q�աp�0�&鄶"�TJ��J;��	�/���o�.4��%b��Vh�r��n��n!M�M�N��.�F�94�j.�t�7Mo_3:�������ͼ�x�� ���W֜��s`Z����&{ %t�iZ9%���j�v^Tr�'6��e:��Zs�=��V�:D^\^⻊���le�1��Xʨ��S�]�R���k)���̈́����:���2�_f�J�u_ٯ�􎏻9E�og��[Ե�T�u|��Z�rx�v|ϑ��[O����v����]�7������K8"�.�jx&��0b�W{;�.�qcg ��m-}��N)�}4}^T��"�z�0� ���E{���S�ە'� +%�B�����%�s��/ݸ7�
8�u=[B�M��V�m{�,��ٌ�D�=�2�4b��R�S8e����4�*�&��.��γ�ʴSֲ�%��c������eZ{Z������.�`���'7DU.�ܲ���4��t���۟7Ȼ#�l��rwe\�����΍Rǽ�o�ϓ)�~����n� ����}��S���y�d�nw�B{�f_6fm��FO&:{������8�l�m��V�C[ɇڡ�P��VqVZ��S�^��X�/�0H
2��gch���.���6vaWNF��Z�e�Yu_<�2_d|�U}=��#7���]&�>b!<R惓�;#sd�1�񶭵�S���j�wPU*�3�.Gzd����Q�G�����o��@�&q�Jsڌk��v�\6�_�	m�J��s͝�ڪup��{i�5l�Wo9gs'q��Ϙޓ��+ǓQj������R�k���и�Y�M�E��s8���6�Һ��LXyἒ`��R���g;�ٱ�;�e�'��i֧ݟ�૝�)��jE4��+7����B��)	�l���=�b����i	�D����9���J6o��x;/�V�l�m�������N^巗�V��-���r�U:�|���^�x���_]I]�CE-ݧPE�he]$�hsw��p��)�q�fg�iw%X���Ƶ�v�Y�RF*��N�Oz�6F�/�Lh�~뗿�ho2�1�k�E��+%������e��\����F����&��9av�.�3u\Fk�]#@�y��jD�Iǋ0�u*.N�Yj��ߚ[���{�}���j{�w��|��I�ND�y99����g\7�����v�[����T��˝5�Iiq\��?�k�5��^r������.����w�2u��J3��eN�p�}O+�Y:�j�X���E��-궘��/3RZ�i�l�9e��2��7�Gc��:�hp�5S���00Y�}�wwP�F��V��e�K��Ĳ{�'��.����,�u�<����qSBt�j��9���[�e4v-��y�*Nt(&9�E(����A�hu�e����G[�l�j$��K�1�u���l��	GG�W��ԛ�}A�MDk阍�zㆸ�n-��խ���
���<{R�-6��q�s�!���{Gk����V3�V�/n]r�%x0��[Rj�c��Sf�k�a#9��Rt}.T�2,�u;D��]j�6�B]�����F2������o�Z����ݜ�+w����ibjQ};��+�c]p�̽��35mnH�cO�kC��dJ/1sWR�u��'�V��'�f�mkN�-�K5L>���U�ȥ�rQ��i<i}N k̚��o2N�$�B���aFV43aq�]�n��K�ܾ;�'N�~����$�(�8���y�>���x&�93vi4Ṷ�1���vz��J��ݧ�8�����{"���7�;�Pӓ������&�%�Q	mv7����#^��=�_�f2Ģ�@�om�}+'-���'�M��Q��Ŋ(n��)��4�3u�ߵ�z��	��)��g�ƽUG6��+������jwQpy�E���d쓛�ח�\f��w�	�Nr���1$��i����p�=��lùP�Z<}qË����R�]���/��g��Vf����4���*�o<-Bi\��Lhr&r��9�+d�iVzk�LY����ؼ������9��{՜ 6i��%ut�,̾��S����L�&u��4t��ĺ��՛�����79Շ�t#j�����Iڀ�Wy��}���s.)�7�}�wo�9�_ϥ�&�ڡ�؞_Q�������<^-G.�Bot_�i*�;�^��o�Ze��S��~��5nP�os�/58f�}�н��t��=�ܜ.���]��n&�.�J�v��s`�˼�Ҡw&��QDl:ԧG��2����D6�����9g�k7c�Ў��H��(uQ=��I�Z��t����ᦖ|���ӸL����ƽ��ͧ�OWcPY��QА#�K9�J/1t���f���mN��(����������p��h4g醺�BUf�W<�Gt�Qw�v(m�̵�\��N�W'�/zNC{
��ť&z;0�٘�Mڠt1{��M3�^���^�{��$��Me��LK�O�w�ߨw-��"�=�r�]h�~�
�<�>�V�V�}�BҪs~����jȃҼ�s+}���k�E����Thm���wxX,�.�h�S}�]�2c2���!`��K�a�b{,�sp�Δ�T)�Ӧ��Ś�*0|K
�����ɝY��Y��(U7,b�K��j�F�W<��0>x�.&.Ώp�El���\��f[��Y�I��'jY����Q��u�V5�T�8�1~����{-ʊ��s�w7U��Z�A�L�W.��|Ӏbqr�;�K��eu�q��l۹yavΗٺ�5��ϤU�i����Zv���v�u&sgnZS�	��Y8�����o�q�>}�bڥ�b��y�F����R���ړ����⌂���4y(;oTv�������j�ԇ�ɥ��޳�i)��	q�����ކ̞�����Z8ۋ�h[l��e����6�[��:ͽ���P]�9��&�ᮗݩ�4��l��0��˨t"�u(�T���� �rG��m�X9Z����i�v��e|��o`�},��U��0��_��u�$���'��:*��MWVv��������E�^,+"'�m��UD��q�RFo[��J�Մ�)���-�G:�.K=��6�;o ��Wr]Ωy/�v�}X
��?^�n4����j�e�h��]��P�*�e����P��yL�k4B��5s:��Z��=��5���̵>ۨ\�9��ˬ.|�[�M%��P;�GB���מ��N.٫b���Θ4F�4��c:�W�!�w������=��R����W1Sq�sލ�\T��m�R��U��5��Ϯ��%�sH�ב9k+X��H�vT��h@u�0�z�Y��+�֩���.ń7,_�����p��`��f�ݡ@�+Y�þ��Q��L�^���͋ mF��7y\�N���o��GG2B��]���1��g>�Z���#�U��
����f'����`&c�IN%˴��u�R��V�Q�-.��S��^*j��bV�i�t�P��
WD��PC{h�.�/���Z�nA٫3��o;pr���Ѩ"ͺ���#%����Gj��KG�@��n�� <ǜ/��}�A�]1�amȓR�V��N�����b�ٜ�yޤ�B٘�ˎ����'�K�.ep�b��W�5 � �m�3P�k��WAC$�P5�bn_/�e�k���$�����u�T�o�*���Mb���/w��S�MM8*�W*��
V)�o9�Uօ.���ռ��a���awT�6����{3�������g���r�T�Ώ{]���*�P��p��=���
���*�]�(m9=�: 	�]�T�1+g�Ɣ���vA��͵�	��0Z�c +L�6����:��W�KN�.Y��\�u�MN�Y��"�C8��e*z��dǚe�wֵ��{Μ�(_W�/w|Ձ3X��ױ�ό���������`
C ���nle%��,�.�}P���Y�C�W]-}7k/L�]X�W�E����I�,ͽ���mҺ�s�X�ռ��ˍ��cd����n!��4f�o^�(�����)ᤕR�J����2�tN7�yT����N��s9���t6�Y���^�K[��WF��c�]�Z��;[mw�7c���M��4;yڤ�S��]݀GO�!1tC�v�
N��o����H�B)��&�2S��¹r�J�]���,N]�� �JZ!:1��D��*�;�h�$�Q�#�E��B�@�r���w<�v�yJS]�/,+[��w��#��XL�i��2Xά�O��Z�0D����h]��Cuv�`���6��*<ӕn��5S0�Ѥ�b��\�&��Å�r��\!��p��j���l�%��9����� ���s�j8��x{Es�Sx66A57������G;6쳭�g�`e�i5b^��s�3��U־��Ɲ�����qW,l�����.I7�[�תU�����{��IvY�!�S��ueN�4l���%Y��R��@NXs+qq��w�blU�q���f�WD�O���2��c|��gb5��I���b�誯�t:`�����0�zv}t�5�CI�X�5==v�L�gt����To�����*Zᜲ�6&�!���d�]��1b�TR#ZȤU"ȣb��(*"�UUQb�UJ�*�UX"D`��B�kQYZ��b�M���B��ł%LpV"��*�UAs.DRc*�)U�
��FEU�Tb�l.P�ETE,��Y$Q,b2�bE�l�aPDX�X�E����1cX���EX���V0X,D1PUX�DUH��Dc��ATAE�U������`�d�(�V��D�b�*+l�r�Ab2,,�*�+iQTY1�be��*,��,��"H��j�4��b�Er�U�DH�"ȱE"����d�X�T����H"
V�����0H(���"��V��\J���Q��E���B)�J ���E�TF#�M|ET� J���V⻘�k��*xE���w���d9�-��J�<�����V�� ٍ�W�X��$:��(.��*:C+��DgAMo.�Z��v/Д�I*�ܓ�K5�ջBۦ�oJ�t���	�~��a�:����ϢK����4��czNCq���y5j��9�z�T���=��'��Xy�"w����E>[�,��o�8X�'`�M���x���b�y;��)�ǥL��O{�Gj�S���s��N�����K0�	�w(��B�2�n5�bZrf_a�k�3t�>��"�t s׊��u��ib�'�O\7��N��yhs[Cg��]�W�p��ox����2Fa�]:*�Y�d8�U�<�U./�ӵ�Yk"NN_��Y�^_p������k�ϳ)Wn��[����S�����j3�\u}6�3`��?A\����(�S��V��u��5�r��No0��~�?.6Gc7[�=��)@��/���8Y+lv����d���V|��ϗ7/������|u�_�W5�8���%1۽��\eP&)E��c/VL�wx]jn����J���ٵq����z�mA/i���b�����V]]�:�㰳�6�W�-Ќ}͓�5M�����o��-J���Ŷ��6S�E<9Ps���أ�0���U{��꫓2�3�C�~�͢nK��U��3{H]d8�)����dP(��+T�i��,���	6�m����C}$�I�$\R�\�IJ+�LT�����ǟ)^0[]-��=��\i���
��"�'�5g�ĉ�7��l��t��E<�kJL�i�Գ�[�;�2RȘ*��?&��ىv��1\YQI�TqS����]&�a�)����\gD<���{q	��5���^�\+[5C\D�u" �f%���|�'�*le+����Oz+���xcrԈ��^\0B��M����2>��a�!;m"z(��Q|��ݕ�a�2�d��<��W�&�`�z�B��܊]�q��-�9�`	ׁ>�S�ܚ;|�5)9��7a����DRrf�[p-u��&���x�x��UojZi"C���+x����P�}SSBq�'e_t�ͽT�'��b��V����"�ĸ��u����]mZI\W&:���(u�9���*�.���EY���aU��U�p�]7JT�;H2�%�(��bZ��&���N �ӣ�{p۝e=�V�玀g3{�\�2���9;��{���E|y;��wA6�sj�ħ�pwz2�ĥwz��p"�mq�]4����W���QD�y�U�����v"�l�řǰq�����ol�����vƬ��+�6��uF��ͧ2#���%Q8�af�a�������fq�I�ʎ�ڡ���ñ���ƷE�Le��\̖�5ƿz��#�nW�����ߡ��q�'��7S�A8pgW[���I0�qρ/;Su��ޫ��Ooϸ�A5�P̬Bc.�s����(q��#W��� r��hks��9�]�d�4�d��{W��g"n��W��)�on+�W%7�+�m��e�-��G�!��c�g����1@r�t���}P��;���OK-a�t����!��ݭ+���s�qagSU�.�3Q�frOL���6�������n������pTu�А����}�ep�'��7	�IZo;��4S]�ة��7ir����\�0z���yk���hGq��rZ*	�3V固���4���i���S�B4��b�Z���[O��YVT�wg���&�6dי�q��si�3���|�FQㅴ��wU�A��10v�W�W=��q8�.a*{��Q�ޤž���ƙ5Ы�ȗ�'>oU�<�A2�O�9����&q:]�R�nBY�����6�%�c{	��rf�=���a;���V�e��Mv��Ȯ�X��4�#���'U�NI�Z&���Oxe,*���n2�-l��vž��7�Tn1Py;*�%L����z�v��{V��κ��	jd���%�^b��__.�z�K��� ��-M&\=�q��-/�R���T7���G�xlg�پ���p��ka��K�Q��� ��get�՜,�j����7�X�~{�B��L�S�|��&�1F;��:��� �����=��g�㓻1&��N�U�l_4QZ�T/la}�]��
�;�)�z��Y�i�Β�ޑ�.���3ml��d����X[5հtۏ�7T9�Q�Y�U�����.!�8�2&�M����Wf���Z8��uSgb���Ռ�R�R���zj]��|��J�5.����n9($bV{�����Y�Z���ًfV�2Q�Vn�D⾂�urHȞk%�����"��������Y�*��bgѓna��sɫ6����S<��S�8[�fv��l��h��u|M��+e�`^*����g�nsm�Պ��ܛ�
��"��Q"���ѥ�����PN�����*aR׵]�������M,p��c}p�1Vi+�*���AЪ��]ѳ}�a/��#���qz�I�f�&N|����u��߫�>~��xPx�θ��+��Y��5U)�Ğy�N�A�(��X������8��d��V,}j,BUfE.{�D�gI|�G!ѷ�/T���UY:j���B�yq��욷D�vV��">��W��;����rr�k��s���6{m�[U��In�a��4����[/������S���o�J)�_9�;��m�xnj9�W	�fVS�0M|���4Y���6��(h9B�
��x��]8���G�v�[k�K�r���vIe��:��j�����Ӳ��C)���<m�R�*�D�b�r���+���M�6��lhA����#����yЙ@���;�eF8h�\ ��f������]M�R��mn
]��N�.���\�)�jE}��*��ԗӚ�n-�̸�Kp�Xg�0*Ǝ��x��]V�>�y���ި�m��.�q��
o'. 3s-�ݦ5Ek�}�P!���^��}�_��uF>�QQJr�l�?_&������׏M�=�$t}���VV�[�qTj�]�|����{e��*�N���'�\���7�&�s�o�Ǯ�3H���.�ڴ�	����K'r��s}��g��h��o��J�χK�B�zno;wI���4oB��m�Vu¢���^��(�x������]���έ�f�N_C�
����d��;;c�	x��$��V�D2�!�vGJ�Oc0c|�F����
?���38�������ҿ�Ou�D��l�����K�KY��ޒ�M��s	TJTMT�s"Qy�.4���M�6�\5w:Ѱ�jw��h�s�]*�Y��S"�1���Ϻ������"��Z��̫�'"S+H��u��<�Vǂ��us�Xܼ�Hb�K�Ty	��6.+��y ݮ�m�U�x,ɮ��N���#��Y��"�{`wmr���:�GTZ�,*=��.�,���!�!7��}���;�-9����i�$��¼y5j����]�Ȋ]�/-��d���K�����ޅԯ�E<��
v'bӓ3ׂ����W
�,];�^�eIp��]�Kۂ��_fD&�LA&�Rw%����DK��֥Z��'�ڼͼHV��Q�*�R���o)�,��i�vD큼P��-���K�ɻ�ƥq��x��'S�q�m�Jڛ�0n���4�����w5j�M_C�:y�+�T�7]�ں���_��7��qZ��I���]p؅�-��v9��5T��S��ɰ
�W�a�7�z,������	��)U�y���'�w�_��U���/g��#:�8���zSk}��S���pԆ���}%<�b�g����\��Hˇ��((sL��qF���9��ۗ�WTnj*�;hh��S��v���L�Ȧ@μ=�y��k�Iܽ��zk��Nq��|n��+��+%����ޙs�%��	:���'+����}7�L,m?�MoVG;��yM���%n�핑����w4˦��F�݋�㏅�.3[Q3ˣ���/"����E��0��d{#����`{:v<f��g�6��ˬ�}�b���d�}G2=8�g��)X� ̗�
J����������!���G��G{bԛi|ׅ�Z�>�&s�_�҆P�%R�:e*��\�@^�9ތ��ҼZ�=ku�jJ���{"��Ć��)Lw�p��z %~��� t6���5������M�5��V�*W(��B��%O�Ǜ�>�o�W�����M�O:�J��Ph'$�*�7����m�>8Q�C�z�
�Oç`:��B��C~�/ԯ�{m��b�[�츚�/F�ϔi>�����a��蠼;+.<v��f�����>*iΔ�hu��}�S�Vt���p�cK�|�o�=�$M�yM�Ȁ<�ee�;]��Y�p��Z8�ӟ'�~�#'��1+��������ݍ�����̜~����C�&��h!�9;�*��n�=��2`���G�Nנ��lW��p��4�8�w��T����u\{
�8 ��6���� I�W6Ҹ�9�^S�)�����ˌ�6w8��<�A��;�s�:nr�3L�]:J���؎�*l-�q��������C�ztr�q���Y��󂒓�ݸ�̬�JEQ'ѳ�q�Y����#�wq��{8}AϪ����s}pĹt��di�f��a��("�n�J�F�s7��c�|��NEdB}��>Bxl���\F���]�2�������y�қ��S���s'��H^�����Y#c�n*���D�9��~����S�c�C%vEߥ^��s�U�D��{����u�/U{�y�1wp'�i���ut�GC���W6�A_������j�a�a���9�/�3!=����\)��N���a������K�����VC������eZSG�uJN���ҝC�zvfBc#�����÷������/�o���+W���9�Y�C(1�L���VXS5ig�Y;��]��q�0�X;�}\��/x�yD�[c~���߻��p���JA�2О&�'�����:3���f�ڰ�K�h�26���fī�elQ~��O�������<����t=:3���u�]S{��^+�x����e�>�c`*>�9�yZ�u\�z��U��T�g>�#��~��-��tU��)���~��/o���)K�w�	�	w)�1�ǒࣝ��nմ37p���w `�^�Jjr�V�G���81�������8T�/�p��Wի�<�= �ۄ�� 锾tf^��:��o&���c�XǕ����U:���'�G����	�FZ-����:��v�)��~C��n�4w��k�^j��]pv5�%^\�G�o�}�d	�^dtU6UC"����U�}c>��	SQ��!��=�#����zuF��Ͼ��y�>u3�Y3-������UzWg²\�޸W����Ч�a�Fw�l,��\��A���i�웋�^�c>+ހ>7��+���o	��|W�i�.��g]D��Oo�{ڽR�ڛ���Up���!�ݏl/]�Q�48y��>�V�џ���o�]�7�s+��g�[���9~�6�g�O��t֎��zE�u���{cҟ��\��TX�~]�C3��dxw���V�8�#��ip��Ϣ��0{������g��q���$�m�x��^�LV�Hk�Y/�0�W�J×�S�鸵�[�({G���ѵ������S<��`����i�����k����7jI���������z%]�œ�(���J�����Tk�ef�����_y�V��3�O�~�� ���:s}�	��S� ]ʪ��<����/�{Rv�uh�I�Yu�>ۿ׎��W���hr=]p9b�ǻ;e��Tv5\���g���%w����Ӯ�%��Wim��k�`��2�olQ�/��SBCS]f�v#�!��uM�Q�
�O�.�ҡ(�/�Vv�ډj�>;3���5�3[�����<HN��u.�2�*�Lȸ��E
7u|s�&�zm5�~�N60(���qt9|�2�n��i+�5Ap��lޭ��b��*Z�R[LZ�nZ�([�_.�Os��S:�)-}m<��4�]�R����`:�n�;�0e��T��拚��fu[��|�o�&��ַ��ɉ��V��dMW���:���]�t�IjZ���Su�Q3���726�x C��c��q�����Bg]dp���bV���T��zqѺٹ��F�'bܜ�3���>ƺ��V0@��󮙝�d�LL�wW|��a��*i��YJ�T�>���=�Y3P��Ҵ���d/uVg7�4F�.�#]���8e�.N����FI��T�Zή���.n�;�-x�e*�͝��J��3�ů-Iد#�F�wR\߁��/�N�Bo@ O%]] ^FM��#���N��4�R�u���7o��N\ZGks�k�;5�^���p/]5o6��6�,�ड़.�H�ieG��`��Wt�niƭ^Yk)Iy�v�:�m^��\N�+��%%h�vRʹ�S6�u��g[�Eq d�=N��y]�V��k��%�j�R�hn(3�=Y��a]���:��"�Z'�"�����3W�t�M�OTzzh�(F�N���L�����[<_4�b����{u�U��s�tMj�ZUn��5f����oqD{��L���rХF�o��v�e�"���;o�hs��r�1�L����
�˗бX�=l�����G�����Q�Q�Z��2Q�
�_TV6&/�`?�~�[on�>��>�n88�;Yآh'���.]>�*�7�{����^��,ENK����I�\#�/���y
Ⱦk	�r��r�Q�t%h7�C�L&K������Gp�eV(���+/����2��w����J��i@��r�졉��On�a�Y&�g"&RJ�]�A4��)P ��lF� �eEB�d֯,X�[0����ٜ��*��yV���0fL|��p�T�;�m��P�*���i��@��v�F8�3P
�Bxy�f�=���	���M�+d�h�V�/-)��P�8�ƹ�NfX)
w�y��ewt$�iF�E�y�;YL��pM6ޡ�&L�T�]��ك�nKy}Rw#��yC���IbJp=�!��88�Z[Qa����,��M�*�`V��'�^���J}*��h����j�WH�Z�Wlt�]au4���Y�Q�3��eKte]�=l)f����IS7�����.Y��S��հ]e��K�fC�;���tZR8�Z'@���o�1TD�~��`����Y"�(ϒ�R"�X�Qb���Edk`�d�P��ȱ`�0�"���D*Q*X
��1Qb
1I�TQH�aU��T�HfQEF�r����Db�*"��Le�
(����
Q�d][ ��1`���J�"�����EVcm����P�RE�E�*������TPVЪ�V,Z��X��X���
�4Q�����,H(�A@b�X"H�����P%IUdKaQk%eB�b�m����E�E ���(��Ab�bCV�`V"�%���ŭ`��
�" ��� )Z�Ab�b���2�+QH�Y�J������E�ز�VF:Lf�im%a�H���JAUA*�i�!YkE$R,=�?kY��>�����z������z�����ΚM�]f���;���+@\�4��J����X���氂���ĸ�������`���Ω*������C�t�y���C���25���h1�L���.�2%
�^~s�Y^��U�>�L�(ϐ]uS�߱O�Uy�Ͻ������+��;L8�v�z���Ջ�}�#���.���ys �@f�J܅�$�B��S�����x�(ҭ��V�r��X{qy<�L�����z��!�L���õb. /ZѠ4=��B{I�K���1��y3��=(�.��>Hې���L���X�^�Y
&Z�5S+��f�� ��*_�����c;�ծIm��=��#k��!g��f^F�pL�  ���>y�1�[晻�.s4e���0��w��<�p@{A��M��~Y����ʙ-�r���x*Uw�E�/n�Xd5�׮�
S�,�	^�|*o�}~����by9�x]A������y�U ��ϟnǅl����J�t��|V\��X����ȳN|S��NAw>�ȏy�ѩ�;Q�2|:O���K@��'������-[߮�8=8�����iԵ����
L� :���~���������B�[f�l_c�$�m�ϷcU�Y��aL��ԶL���oe��x�Nȗ�X�X�U��*���7�'VtxX��k���f[��1���t<���̱h�JO�8��v��)�ƥ;oMu
��t�U���u-4w��Dݮኬ���K���=؞���nٵU�=w?�=��my�M�4�����{�ط�1h�}�^s3��g��o���8w��OB�M��-�ò���eu9��o�ic�@O���HU�x���J\Ϊ�BU�<�~G���}�B��q�5�2 ?r�óY�V&յ�t�K7��v|��-������Q�\�W�h��{a:�zF�޷�����\?j�{�p!;WM�{-�dQ����t���4|�6=F�BȻS5�Xs��\�[}����/xW����~@�G������֢m�w�yQ�*˅~��|!dtU!t
�"���(x��޻��u��߷��~�7��w4?F#<{,e�|�}z1*3ވ�j}9򭗐�K��3'¡ɶ���x>f�!܅�)T�0fF���o˱z�-�FF�(>������=7��{=:��0�e�0�n��W6�"2��_a���ԋ����g��	����*n;"�!����zF��糧~uN���-:Ϫ����������u���>��$n�!O�n����7�y�8�4z���ǽS���������o^��Fl{g�͋���TV�^�un;kj��R̉��<�ɯU�b�Vuu5F81V�nU�і;�b�/�)��p���ݣ5�1�zQ��h����Ӯ��Sܚ�s�FE��J�]K����|�$-�Ѳ��d|��oRV�m��L�S�mZ��n������QQ�q�@���c�G�p�)�-��)����y���}2�k���*����
P�����w�x���;+.<s�����^�w�B��'xNC~���O*]��+�Q���Iuu�q~Z��~2 G��.~K����m��=]AG�׍g�����8s}e��Ǝ�Lh�t��G��s4[��Iu��3�����VJ��چcz�F�2���W��^Ǹ�m^����/n�b!z�0�ǖ@#�˸�}/lh�>����h��s���^��"�e��%��٣
�{��;�<���}2�{c����hqܲ+������#���6=�9m$q�~��jw>���썯M���Oz�4ә9�'���c�{������Ŧjw;�FG�v-��eR���[4�g����;qW��mWxg���y���n��u�>�Oû��2݈�<y����d�6P��٤�E���~�-΁�ԣ�.�N�ts�ǁ9,D���� ������}��J�w���c��+��F(9J���E�d<��L;۠�sʱ_�*��6�Z�r��6uQu���P]�^oh��'�v;�ʒ�z<eEB�>7��1��0X�.���5��j�=� ��#��<C��t���r��ao.\�+�P��JJ�wx�;��3Mrˁ����lZ����K0�i��(����^�C�*��#���;��~�t�w\�����V����y�:��2���\p���{J����#Κ}W4�o�#��m�<�z�^�g�Uu��H�l��*k�NkՕ�5�E�qH�g�e̓I��m9��	K�5�����x\g��1�t?�j�n�y͔�W��O��r**��e���X;����5�w�X����S���t=��W�%�.}�9ׄ�具�^�-�q��2��**�2�_[7��uv�N}��������7>7�c�vj��{��nCߓ���ofGM���1Hڦ�ʩ�E�zj+�f��K��[�����p�����5�G��3��_���ߨ�~�!��:OR_�d����g׌�I��s�t���RE��,z�D%L��<��ϋ���|���������_�~�'�c`#���Ż��7��b��/%���}�]�W����4�ؙ���?]�Tg:�3����<��S������o_�#�������?E�p��/6�`٭�u�Eg[�����z�t/\���{�N~��TF�U��3�1�Z���qx,-癲�Y��f�Y*̈�w�;�S�;v��5f��y��H��E�48�{
��Ÿ�Ȱ<W[-��q8�f.��C�b�޴{�(dW��!����E�mt��Q�n��k釟K���E�{�g"��֦���p�9A��;"���F߈s��W�>�S=�ӎf�Q�~�(Ϗ�r^�;X��W�mZ���}��Jܒ�NɈg��r�w/���z.6���F����s<����~�eS����j�ق;�������y{���RE�~����9�|�Ϊ�J�μ�LW���9zEwoqgͺ�k�4��]�'���߃G�nG��k�N�T9S4lS� ����#�����G����' �mQT�a���Kד���a���C��^C�������v�W��z��ǧJ�Y�ޙ8=�z�}��ٙ�[��m)lc캟g����U�6Tz.�_���������\�xwW��*���E;�d��P�lh^������/y��z� D�ycF��v��>����g��^�lzvw�CߤKu`o"�X�ִhk7\s�1��6?vG_oms\ux��ϱ�c��ԇ������r�Q"|��T�c��k�&���F�U���xb�6;��p�3���/+���m�c�Ι��o��;�J��S�F}P�;�iQ_��e1OŸh���WZ\z֩�x�Oڐ��+/�}J�뜲�xF�Gjy��1�Y]�%�w�:3��<��y��R5�145�5C�6�����n�x����vɺ�uΠy �mn�e�.�"�������δ_t��Ur������D����X�'�����O����ߦ������;��z��T�Q�`c� �&b�
W���{0J�H����O��b��z5X�q��T�w��
����n;����O�/��ϸ��g�5���q�=�'�W���z��:�=�b(y��Y���I�~�]"�i�>�V��z��K��$.׽Q�c.fe��d��v�87���O��e#�9)c��"6��<���}FE\gc�����۩Oٙ�s���)�UD����7�nd��y��NP#r*�:������U������l��z9-�=�W��s3�Y������a���ke-�ò"���r�7|�fz�}��C6uEk�Ǫ�Mu�}�z��������w����"�ǰ�	��W�4��ve_���h�+�"|�eV�{j�=�Pb�ܧ[�^Oj~�H�;���8�~o ��P󝚗���j+��C�hc"�l��v�k���>��~���R�(��{�
��N�?;����A_���x�������}�?v�k��Ǆ�T�� �"���(x�	���p�.���ǌiRs��뫌I npn�oh��0Gq��aZ�7�K� �����pM����K;�L�oH��:��
�˴0:��0@�D�����E@h5���-�l����ė�]k�i;�k�U���ܣ�]��SA11:��֞B����n����-Y&fh(\j�鸷����H;П���<�.s�F^A؇R�2}�Wm�@th^���m�^JO�%�/E�~�G�}I�==ǽ�=7�g�ӛ�sc�ҁ�d���&/wMN֭���>�p����!�=]p��Rȷ^����&7��WM�{T�{�~��f[����1O��v��Z	F�����
���+��#o�!����W������f"�\!α�ȏjJ���d�ǳ��0�4Hy!/}��[��ӣԸr��K~�+kֳ��m�U+PG�Q��W��پ3=�;�/=hE!�Yp�Dm��j��1�~B��B/49nz���ƽ^�9���+ڇ�4�hץL��"o�?M��_��Q׶U[�5����U��9X"p���vd�����>2g��/]�3��s>[�d�w�Z,M��7>�rzE��ﷺ��2�M3�p$���\Z-��^`Vu�a����O0x1��$3��Ȭfƃ���{��UgLmw>1Z��K����#k��8?C"4ә��g�=��� 6��iȬ����!�����SU����>�����q:-W�х@!����S�Y�L����BR�&�HcL�SX"C���W�^u�dʼ$�%�S�`Z��V���y��t9�b=Kh�ਡ'`��EѾ�uL��ֺ�+�HT�fV��v\]V�+��p�W��n �b?E[zv>B��]10Zݴ�1G\/�K�������}`bC�Ns�W��mzo�1;�5���ߒ{��֠�g���I��1mƮs:�'�\/A��#�#�	�v�oj�9ȍ����s<�!�nIf��'{��;~`fpy9^���ޓ���WO{�qI�#��ݚHdE2o����=�\Ƕ;3!3-�V#w����מY,����g��>w�ez}q�f�O�B�[SF�(9j�*�����^1C��g�T�ޫ��ˣ��⏫�{� �=�q���p؏L%�����w�ꭰ�bd#�2}^�@Q.}X������CJ{O,ng�G���,{z�yo�#ڽm�^V<��x����Ӑ�l0�YExL^��蜟l����G�:��z�_Q����ȍ�>c��*پ�C~��yJ���T�DGt����s��%���Y����xV�P�=U	\FY�pc'>
���/aR��w|���>�y3W�]������c+���_�������Y"**댴W��������-ϗN�)F��C��~��j���莵y�u�c�Ιy�݁7�����~��f��T��0����lQ�c�r�W��6��S&�NU�>�ў��>}\)���f�4�?^��h=�B��Z�ݨ�}������<y̚:	+�F����
��s�����������ŢR�>3�j���ƥݽ��֡�<�=�.KޜS�U~��{`;ٙY���c��}^���'nlԀ���*�޽��H���+�ڡ|X�J�FBy7_�X/��|��>̏o�m��^�}��d�IS��ybܼ���<��g}���k���sª�~�{�ص���7·��dy)�&���7{J��z�Oex!����o�?1ë��?mwdmt��9���ng�K=���;�As�E�Cl�T=[w�i*��O̫���`���C�v}]p�6�C��Z;�L��4���Q]q���ϧ7
_+�n���H�<2v=����)���[5��UP�(���{�69���c{A~����\Ο�1���x�����إy��?G�M�Ϸh!�Nt�S��ͱus
bj
�0���}�+����� ]�i���#�����#���צ{�E��3K�vv��7�m;�]�.F�����������~߳f����lx?F�k�d+őѹtI���5㞴4�m?:��.�L��]����Pͥ-��U>>~�>�U�:w�]�Vz���4P����^���.E�o�r�yIc�����js���<�v�Υs��ck�y�����-�ەu�->|�f�}~-o��w����Ïm�o
�Npn�3'0�3(Tݍ�m�Z�ݶ'k�Ζ���HwA�u˥^o-�Z��z�L�����wL&����\��ɽ����Q�����X���:�g���X����м뵛���M�=���_{rf��Ec=7��>m|&p���;���lH���2�R��K��k��8�����'1w�ooiK/���7*�=�ԇ��ɓ7�yS8���D��dUL�1
�0�s�5�]��*W+�2��� OD�?��ȼ�mo�y�)�>����Bi�:��r�I�P��״,�e����6��lK��	U>�n?,��c�7�{s+�(�M��7�Q������n�_�=�xvV_��j�>��T�G:��ʭ�j�Ɨ^��>~ɵX��E��=������cS�7X���Y�\5�m��Fפоu�*�G�"�ө������s!w{cr�<QΝ�{��T����z�~�C��NO�c��.��<����dV@�:�ѓ��j��KTI�Lϣ7�����y��]*��ݻ9:�kd��T���o�ë���(���'�y��k/���0�5����B�y�6������9S���N|���K�����E�4���i���x��Wb�R�1)���\�����������GQ˔s���v�j�_PP�V4[�YA�$·GJ���v'L�g<�y��]��+��CU�f�H�lpt����V�;��ݝ�W1�\�8kp�̼9iw>��T�}O���g �&�G��Ɣ1��Ku���7ڹj+{˺m�u;�ԥ�"w��,S��W�oI�i����?h��mIV��[��S4J��;��:�2#�� j�⑧[�ky�m��੮�V�̽=�Eaʁw^P*����*���i+	譙xUgq5���Fa�J��q�7)Kɹf��V+����LCD6�<BX��	�C:DD�F�Zt����UbM���-�����U���`�;�Y��&Z���	ή�3t�m�m]�Q���袆M����Z�ą�n��k��x��S�wa���X���h��t,UV�n,���� ��8//��`D�c������}���R�W�����8���q�E��oms�o�B�R�cG+.qr9a"���Z�ޣG�;x��{ۗ����\���bܩ�,��9V�X��Kb\�{vk�ˌVs��3{�9�!@`j���"�������6��5s$ǙԳ���e����vc�bv�&���Z�5�X컱�p+!Ճۯ�8[|�<��<M���l�\ե���ҘG����4 ���fS�k�v�Ӣ2��#�"<��D)��=��k{��A�j�����P�r�u%0���+7���Y�&����T ���k
�ISx�W����k�
��Z��2��磞EZ��b�<�f�pw��:U�������F
���w�l��4�e&��鳫:���ݽ�����-Q���LԵvT�V��1|gL`�畈5]�Ԙ�'t����Ǌ��q��U��]a΁���nV�g
\2���К��B�5q>�:�,�\Vծ�X'��*�/1w7X=�XG̡%ؗ��h��S��Wr��g8^���Ci��M��_gLF�̮��{��ۀ���B�����Q�'U^'s=O1�5wn�#"B��.��n��3�8I}�]�GCw��b���J�����:,�0��]�M�ۻj�p�/�� v�غ��-ƴ7Q�寖�(h��M.��4f���k�L�j�*���R��rQ���%�,X����n&�J�W�U���{*=��Ѝ.H�n�cVM[�4VL�	�����I܀F��U��Y͍B�8麷�WuwN��'C&#��i���-��k��9�݋���s"	I΋PI]�m։��S-��*�|r ;4ЭsdӖ���v5>J�s�Nk�Qstk{�� �����ٷٟ@}T|�>"«ATQAV,X���
Ŋ
E�����[4Ll��&���P�dP� �Ea4�"��X�"��Vk5�P�U
��(�"�@Z��ETT1̠���²LH�"�(���ŋ-�R�`V)"�dU4�D��AEPEI�L�DjQ�
��H��V��
AVCI&8jʂ�i
�ʩc1�`�PEC�Q�Z�ZY"ŀ��DX���1��� ��(E"ȂAdEdY�*"YVVCV�,%B�i
*,��\�0�Yt�@�dX,QJ�X�2J��X��YU������\�P V1X�E�,��C.�0Ab�R

C�"�4�@���H�#"+"$D@L��E�B"(��g�׺�N��|�<���f�o���
��-��o:����'9uY�hcjܐtR��9�1�O�r����ާ]3�q������;m����=}��i,��'�2!���������a#����MTo�lp��&�[fW_z*q�ж����$���K�����A��r�m^O'����߁!��)fa5C1���54���f)�>��3F��ȧ[ �]����>t~�|�����}#�l��s���8�~��g�݁z=��C��q����6*���aV]����kn�y9�^�p��8���}�2|�t�x�4��_��yj\ꮗ�uԻ��2}�p�۴�}~���΃��w��i\�r/�����J;�ɞ����P�'�n�L�t�}�^���W�WE:u�Ѹ�ej�O�fFF�cݿ3��z�E�bC_� ���Et�{T�w���=u�t�$��g9P�S��]���yߤ9\5~=��^}�_��3ީ�{��3�~'}�ڷy=+�d�m���슊��2���>3�iB��~�%W�g�7�6M�͞~�#�[�9}Y$�_Uz��g�	����~�A��Yp�F߀�j�Ʊ��_!n{��/نϩ���-,���q�����o�x�UJ�־C�^�vp�%��0�p�([�3c=����a�W��������\e�Bm֌S���QҰvn�l�P��2e�9�8�Z�F:������9\R�ՆFC����:���}3�w9{�;�[F��}�HNT-�}.Ǣ���j�'^F����R��L������]C&}q�r�Mǟ�Ԍ��!�����o��QT<����3*��
����y7��.�xdC�){w>��E��9���S���W���|�u;̠��Cмݲ2��3��C{���^�P�+�EǼ�v=�;[��!�N|K{rȇ�s�{����-�Q�;���]}Y�O�V}[N&�<���W �ϼ�p�������`(Y�ݿ��{���|���T�������zkB�Sެ�Nd���{��2==�R������G�Υ���ǣV���{�f��P��-��V�	������`g�ߣ�ֶ�~�ޜg������|������?n{����nHH�= ��?Ֆ�6���ߙV��V�ѭ���K��/g���{��F�w�������{�zǽI]SJ����sk�u��Ƙ��.������(�vy���A����w�?��N���U-Q��J��zP��igh��<cY���Lg|�m׬�����мڹ��~�^�����Dlw�����zn#%x����Đ�L��ڰ��*d:6��S)�y��z�]$�4�n��������!�Q��9��
u$�mnkE�o�֞S*E��\�1FM��g-���3��0��Z�ɩ|�4�ގ��p��k�j�rDVV�T����q&v<������ }&_��2}N�e�@{N|�k/*^iX����#"��(z���R2�^�e�Ik;#�&�9A��e�+�`��xn�7�y�kp�F*�sy1o۽',���z�U��L���݁7팅�!�r��z��l״p��q@V�66����U7ɮ�d�Աʟz�匏*r}>�t���d	����"R^��@�����e� x������!v�lz<<�:�Ǹd'�9���`y�ώ�w�2��F	�� ='k+���{-���k�se����1�P���z�%L���n;	~ѣa��3Hcwq���O��j�B���N�F�*�@�����+7���mw�_S�H�>)��yz�:����F�Nt�����ZhlU��-���DI�2#���C�vEu�h�1��|3���H���s)_�=&�#� ��;ľ���G�~�?m\׺�
�?^6`��?c��5KA�)�~~˞��9����z���f]�=m{��f�7B}�@^vd�n)��g��ql�p#���n�e��^׀�U�m��T$��h�fH2o*�c����)rk������5���6�-e;���F+bo\-�ܫ�O�����R�F�� ��i�,��5��v����:@��[�]_IVT��q��A��$��%)�r6=��F^�E���vjQw>����ݳ<�RǢ�x�����R���T��i|%�\0�um{��_���<|��d����]�{j�P��x(��#�����&{�nG�z���,�-7���#f_��3��L��
��jf����T�zw�r߆����xc#��#c�^��=�W%̋ǘ����+�y>#�f�&K�s&�Pͥ-�}�S�?b�lD��+�T�=��p\��&�*�gj*���h�3H�������a�.�A����C@l 2#B�|͉^̀�18�X�2	�4�վ���ږФA�<-�=��C|.�-��[ϮՈ��kD�,����͓�<w5o����G5�H��ZA��Ho��&o��<��~�VCؑ>t@�ldv�K`@F�{}�Z�u����.���Ū���m�~^�����e�����*����т��Ϯ��ye��%�T&�X��G�lH��pԮ��~���U�,g��z�������{��Ɨ{�xO�p��vV_���Ļ�\*o�u�a
s؞NG7^P�����˅DeX|vL�b�)�s�!�����m�i�z�3Ӵ��	R*�;�>�ɋJ�˰�,z�f���%E#j�)S�b�I�?���Ĝ�AΚ������E`4��<����#�H�ōR<�w�������w�l���יSc6�h�/�@�h�a\�2���o"�L�˴'}ܬ~����Q���t�^p�8]C+o�=�@�:������(b;W`,�����77ް:}�7+#<�yמ�Ϗ��ĉ�򙥣(2;>��^����z�EC�t=�Z��O�qܑ^2+�㙛>Ǟ��<���bMǽ��s���M��P#r3=���{^A�����5�[�nޣ�Uz7�]���֛����y�=��ho��\��N/t�NB�8б�������Z=i#�Ǣ�)��o�=�^YY��=��j�'>����w��ڲ*��En�dn��k|�����O�Пp�U�S���<}P;��*p}W<���7�k����r<;b}*i܌Z�����6<^���XB�0 ^��r.��}�|��K��/h��~i\��Z��d�\[�H�m{X��>���m�w�#�=���z*��AUS�غ(x�Ba��/g�<M�.R�o#�����+��ߍ��ӱ���{=+kَj�+w!Ի��O�*���i�~u��T��G���x������@B���{b_���3^@�w�g�����ߕu��"[�F;v1	����k�j�Ji��U���ֱ�00Z��[�g��wK�%��=ٸ�1�����֑�q%�:h��Ǘ��c��c�VU��&f-fp�����匘�}S�<�FI�s0)�˅i�h��`S�Y��K%��x�w������g.�1�T��o��7�o��+d��s)�!S�w����3p_=K"˿ca�=EǢrO�=�ڜ�nZF�����q�����U�H�~u�P�US�א݈��p݄m�g���Ͻg��W7^ˠ��վ'���+^zE>�N���	��ݻ�@�EB��*����Z �Hs��~�>�1~���w���R�>U����U�2�G�@�w��Ee�9��"ڮ��ν$���,�c��kh�����t���xNG����w>5��f}��"n<�6�dUyϫ.������xF	����kNZM���Cן.Z�N����B��c!{�3堳�>���.�C:*��Y>0�gۙ9�з�(�Ej-xOx~�=q����p���~��zv!z�0��yd.=�̏lCu���(�9�\���8�����[>�]^��[>?mu�g>5[.g���tz��G�:���!:�2�W�#9�/�����@�t��S��Z��M��u=����{��zI���/�H��욓���{���{a͚�v[8k�WXY�|����o��Zx|'֖~1g�ꒌ�w�FT�	��f����Eۋ�0��wN�~�a�E�Fw��f�HU�3��.����c��HOgõv����ص��gpI��5�t���K��B�a����ȱwd��c+��P�Z���t������S&�D�c]s�6W;���Ro��Y��3~ �������8��٤�E��~���]�
�#Q�kV�IrN�>��+>�o�#�����yߐ=����{�x_߿`|:��K��GùWn�p8,���'���9�.쇛E��? �nK����I����&]�R��D֖���+re�(�>�9��ue�3Qo��I�ټ�aG�<�=��H>ø�z9*�|!�7�+��&�i��ef_��1q�d���\�Ѵ��s4%,k�C~��P���/�iS��8��*C��z��z�p�9^������Z� �����3~�}�c�A�O��o���ɿG��wΐu�o�x,�{�&��[
%�Ƣ�z��V���{��H����T�ݻL�#8�Ɏ�|E��C�����y�>�r�{2�����-H��>��du-5��#}���>�:9�G�yڱ��*j���qNǛ���S��*�̯{�c�����]N�����ܷ-�e���L��Lc��q��=c�F'�q�_�`��s>C~�ّ�:)4^Ѽ�qTn!d�m��401�nH�ڤw,�RO�#Q�_�.�^�ֺAǕТ�2��gAy̫���	�L�X����0�HbºKj�;9�Kz��WfN���Wk�fMAl-�->\6 �<�̠zU�V7�s��B�uq������>�u�{�W��Ee9Y���k�*�&ܑU�C�Z{�Ԟ`�@����zus���3&�|	8�
�h�븯5cG��D��~ǿ��������ްj����m}2#֤������7{�Ou1��
x֜2<�rE�㷓y���8FA����]p�6�C���wO�C���т`���ͯD�����y�P���I�������^➝��}+$v�/�T<>����t/��T��M�7Е��L�5��~g��2#�]�Ez��縤��ytڜݠ�\P^V�m��o�ςE�b��:MƬ�y�]�����6(���A�<GA�?{��-����>��OG���·/��BrF�J&|e�T�)
} �]���쇑�IקY�~Kד���|6��$呱j�t�[zGm�<��T^1~�=��v��`�[�3H]�>Ȼs6
��-�������O��ɛɩ�_���{��3���U�2��=�m�!l8�b����.�b�l 3B�|�\
���r�[��I�_��j�9��{��yM"�z�z�~�l{���p�D��8=��7��}�l8?v'��g2G�\�&6�xG䔃�
��O���[O+����=�%I�:�h�-m��n��\�j�@���W�t�]�wp)�c�U�R�ږ�;�M��z���鬜�˶ۙ�'מYegnʰ�=V#��i�Wj����{���1.렮% �zE�,�
�Kr���P�Cۿ6�)�$:L;��5�ڐ�9�fT�ײc��p�$O�8U���>��c�=|�j�g�)�W6�h�s��\?�ײ/"�q�O������y��5�q���\���Bk�]C�]>#"�z}b�6��!�w�a���[��߆G�c��ЯW�.c��0k��=�}!͍���x� ��7�(�6_�G�T]�O1�P�<����B��	�ܛ�
����{�o�mC�Uϕ��2��� �lP�"+.���6�&��κEs� ��sW��q�J���k�N}沞ǘ��c��O�۩�2��l���F�p�|{��	�yȹ|��3�V=��R*�Lͥ��O�U3AyX��e���M��������Ͻ��^��/����c��7�����nfO˱�ߟ���Ǳ�WY��mM�����Sj��z� =���`O��C��+n|���2�At�`tB��;~n��Wo��`^�Bv� �'k<�{'���ފ�=��М������֞J����w��-��{b�z@|�G[y�#�}�.:��O��w.%��RI�*���o^�,DMk�>���{.���*_�v\�,v'�FK�A����Ȝ{)D{,Y�ufC�)͝��u��iƼ�oX~��_-y����K`�.#+��muH��a�#�Q���tF�����+.���*�CM������@���r���,�dG���=6P�@1�Eۙ�����#j���/�ԵoMz��@��ＲW��M�������^c��~#!^,��~��:*��t]���(x�=E��ZK��=�Q� ��!��^���i�v=�������®��u�;�d��ޭ��u�����r垇>���>�X�l3��g��=��~����w3�Q�{鮰����~�HX�x�a���!>�}:�e��׬�ͅ�R3i��f� ���Y�;�$6� �߻�]9p��',߷����U��}l��-�dT.���@u�7�9\5~Ԯ-;9��mFՁJStM�~������������bk�n�	�������t|:v�p�!�ߥ#~U�2���VuG_�w��s���^��^�\�w�A��Yp�׀�j�Ż(����ˮ�;��ܞ�q�RO���??U�d*~ɳ[�]3�͑9�NE�x��Yp�E�9�=���p��7��yЅ��P��>�k=&S��J�PAyT�>�>̟N��bn<��}���4ǿf=Q�-'V��OL����xM]ZU���'�&��p[��<���W�f\����8.G%�&��i�TU3wݗ�J3��������{VgA�M
���I��We3���\rp����(��+H���kA�8����R#+�^g���ռ�z.����b\�wd�͜{lM!F�a��ޛfZ7�E�v*r�~�{Sj:�(��g"َs����׿9ټ�� ��e_ab�k�{9Q���J�z��;�F0�RK��X���N�0��fRW	���8�hx)��9;�M�����-+��-�W
���O�Pŗ��cu�DnJc�MV�/��v��Fң�2݊�X�B�q�y;f@�S%�+S�}E��a����It�WVN�g.G2�5i�ʋǮ��܉�o���'��Zkl��)�0�m�k67��{�� P(�j�o N���-���w�i��$�J0�!T�A�BB��8��&����{vTޮ��K�@�&ʂU�N���b���4��r�jԏ*�&�EK���-��E��zڵ��|(Q9˘j��HJ��Tn_P�k����2��:s���5��2��j�v#��Y��;��\��7z�vu����, ���Ւ�����c=���T�w���[Y��M^��u���n�qq����b��r��y��`Yl#�TuՋB�7����5`�b�`�˯;��X7�yJ(
#R�t�ɜ��MZx����w����
��F���8�D9����H��uuՙ`m�q_ڷ�}��F�W4
�`���Uޓa�+�5�������L���)�Ӌe�v`W�c[��<ؕ��;����tFh#-�=�����\o��v�Y8����=�����m&a�o&�ZgD��s��D��5q��{�Սl�aBj���5P[�TxlRa���s��h��34�W�b�)F�t3��]'T:m���d舼�c0gFF�����{�}�i�h�՚=J�m�lc��RA>\�ZR
C{���\�)C�lP�[{J�SO���ɜgU�7�o�C%�����*]�����eԛ��M���c����<R¢����ɜ; wϰt�,Ko0k=.�]��E��bK��+C\�6:|�woV�e���:�|Y�u�x��C��෮���;�H֟4��^j_s�C(1�s5��<��bib�ewc����nml��mQ�x�53�r2ޕ�W���/�1$�S��&��h<u��@��k(��(s��Cuf�H�޾k#���6�����F)QӜ���*�wS��t[���4�����;4辜;3,��@ncU+1,m+�ܬ�YDw�nQ`/�_0ެ�ʓ�!�(p.��*��z9�g^���qf�
��oj�o:��L�
I��l�+qw�)ݳ�����yHxu�ڳ�LLd��6�]��u�:�&J�Ǖj��M�ØEtk:��,y-�����哂��~m�v�Em�K���\��H��)��xf��Ӈ�tt	&e�k�a�!d}c��B�-���:�fsM�md�aQX�S0�*Q�As����q�ҩH�*��j�Q���UXE��

�1��
"
�1m+2UJ�U[T�"bն�E��"�(E��t�
"�,ZJ���ED`TLJ5����"�"�R���"Ŋ��*�2�l1d��(�2
�Y`��1`,D1* �H�\W� ��X)�
��T�$*��b�B�**VJ2c �E"�T�
b�
Ab�"�� 9d�EdP��,�R)+`\lPRED��bR�k�`�bхVJ�Ę�d�ʨ�XT�$XĶ�)+H��d�=���_��B9b��vdEok�&mAѐ�6�L����.�o3)�.R�FuA����)([���fV7՜�q\p�����u�����o��@��Fou�ȍ�dd
1��>�����c��7ǽ�̊]ʵ*�Vfx�U�����`Zqҟ)�>���U|2+���z�^�]��g�i��j�l{~~�a ���G�N��̨#�竇��n�ܓ5��s8����f��u��;s�W�dmzo�s��VF�s'�j�j]k"r��Mn��������
U�lp��k�	x<�۝�ھs��	~����~��g�T�9�:V\���x	�:�Ol��~�Rv<�##vi!��r.�����13�?I}8�t�7��v-�؃n��~�F�yߐ=�d�Ͻ�.�p\6}h-MJ�Vb����Y�~�-=}����'+�U����Y#ix<g2��O�#�z��cƓ	w�=*s�x��A��K,lΏy�D���1���'�W�U3J�Q�>����m���L7�sH�~{�/[c>���yHv�՛�b�7��V;C��nw�W��$L�/�jd������@dm9��ؕx���
�W]�y�쨒c�i�R�1���ǐ�<6�A����9�e�� ����xlz���c���q:�Y�IB�%����qv�G؞!���N�of]�L&o�	5|��j��b�*��1�^O�5�*W���޼�m͸�<�3��ȑ�>�ei���eG��a�}٤��JŊ��g.!#5*s;+�9"(吶E�t��F��ݼAY�ju��r_�����May��=�do�g�}�'����ި�^���ǏJ9�b�Of�os�|{�G��ݿ!n}����y^xO����^̯Do�`M�;��#b��Fr���;eH����>��=�5�}c"8?v!���ٜ��y�>.�|_¶fU�!�e���\y�\�����P� z��ݐ+'�w�K9��������<����~w3�:�~�=��z��\i>���m���x��J Xr��޾��^���ER�iϳ��v=t��<����ܽ�GTy�tC����`�
?�>C�vEu�f�p�Dmt��_�T�w�O�O�2k�u�H����=��a�<r4����~� �MA���so�9��"�՜��q�Ӿ>��c�5S<��8�n5^?P����' �qJہ��afH����>�'�sPk���od��)�z����l��g|���s�k��7��{�_K�-�.|�iO8c*UV�Տi�`9��,��U9Ы,z]�̇�mWz���)��/2;a?g���{�q�!�}��<wp�������b�r��у�tr�Yo~��Y�.� ٔZb��o?d���OL�;�+޽��7��k�Ǘ5qLMb���Xw�L����&<xu�R�Ӿ;���M��_S|(��:����yħ�I�}��en̉����{�I�8�a�4l0��f��*A�3����ӯO|n��>��c�y�8ρ�U1Pb�5��e�O��5G�+��>�>!F�O�.��]������.���#���@����a9��OW����h��z�@w�)�G7�\S%g�칰B��� ���g���s�1�r�x��I����ȁ�6H=��s=y��Ý��d�hL�n_�%��cp������4"{��L�y���縐��~���R��d��g��NG����w���P�=�O��*�rW����O�S;���͏����ꚇ��?{��G�g�g�td,�{:fZ�Nϖ���ʾ={t�:��3�z=@O�w����bm��z$?᪩�ϡ�M����cw5]s�}�����%���oy���mRۙ�G��@\c�@hoDV[��o�K���
����:�9��=�0<Z���]����[Q�?z�g�0�����C�ȡ�Ee�Y���k�hFh����tȠ w��H���^R+�ᗋ׀zs�;##�w4k>������R&��f����������ng��ih���Ba#\x��o<��8�ٝwd@�e���'��2�_VsK�GZ*彥�<���w]��ې(�sk+�.K���"�v>�$��e�z@�&�wi��Q��Z�r)KZ��t�Q�(nr�Y�Wm�6��b�=����/{$���>�"�:�35	g�ӿ5w^T<�ԕ����s��l�P�t��?M��b��x�){�?E��#Y��o]����Zm��]�<�Qa;�����L����)�3�����62�ɟt��#����s��셣���s=�t���z�Ƕ��W�v����_w��k=�k�;�����p����9�ڟh� �Tu%�R�����k��4�N9���U��o[�ƚ���$d?k�;�p!�F�!��d�s8������c;�!��o��ή��Nz(��[��`Ϙ�����x�:�=�Y�T���>�s8�3Q��ʌɏ_i��9�E�����d?K�!��gNǌ�@�~��O1K��]/ �:�uL���ݒ�[Y���fߪ��YV��^T3�{�q��m�+ҋ�}=7�����Vg�d5ng���/
[#��K�\ f_�/�sp�#����(cJ����~��`���+n'&X��Voo����xϾӝ�9��۠��-�._}������Hr�j4�����B��W�:�qYD$�x���d��!�ִ+/��g�aJD.6�X�\E�r�eg�JФ����T��ng�slyIn��U2��Rj2��ºv�'���ژU<��έr$���v$�<�e���P�#Wbgp`� �ƶ��e�EX\nQ\b]~Z<s��rG���^�;A�sꊅ��@U�>;��.�8��1;��xU�����N��{޺�����>oުدV̬�{v�;���ˆr#o�G��yf/B��Uyj<B\Y��z������ ��Oמ<�|h1�>?xfT���?M��W��+b�������(ͭ>�x�}���=�k�B�>�������o��T��L����}=�&�b�9MV�^��9,��>3�Tg݂�Z�p�z�A�@�ۇ��e�|�vC|�o�ʕ��y՞��mv#�}�6�G�a���+�WS��V˼۲3����Nf�Q�txAĊŗyY~�1Gw4�����C�T�}�3������l��Z4�X����Sޮԩ�z1���#�|B��L��y둑�������jȬg�f�����ݹ�����3�nW݈��/�Ǣ��&J��������'/<�?=�'��J��\b�Hg��c{�'Go��3�UvP>�8�=�Y��j�:߻2�zM;ǟ����w���%;�Sӿ{�/�$z����j��-VV��T����R�nS;n�NJ�k9�#�Z�3s�0u�(�W�-�C���:bt���b$f�ce�[g;�� ~S����L҂��=K���歛�|�a�Ȏ_ga���9���[��M�u���Zl{Մ���MY&G(�j��p{���OU	�n�A��Y�C��L<g2�O�"��{�ǂa��I�N�y������J'�fw�o�*����W+�K���j��H϶�"^M!��d{ez�U}�S�/�'*$�ͽ�z���C�E{=��6�H�lI%u�.e����s�;~fġ~&~�;�y���5��{_�t@Z�����y�����t=9 4TT7b˛��ѻC�`��_L�:N�ڏX��/n}�o�9���aK�R��g���n��t��1!�sꊅ�ݐ����<򶮢�iOi��~�0#�����^4z$9��IJ�+�����>��_L���V������C_�=���wj�D���2xY��پ��=�N��'�9?+�w3��̯F�y�}zo�N	�؇��>��2���Y>���bU篨_��2+hlC���/�0_ީ�������#���ޒ���:=�݅�3o	�x�>W�7�Qxt�x=*�~)�/p.�>�f����t{/}��,��7:�ЏUQ�tFG�ّ��^�џ��>cLW_���l��t�	'J*�	�3,c�e��{bh�X.�����h'y4�K���;��pV��X�Z�q	�ֹ�_�I�f���)Sw5�b�F4����2���C�joA���X��iՍrμ���k���2нcrR*����G��M'd�{��yb���2Ԋ�B8�n�_G���s� ���㷓y���8FMZ��]�b}9�s6�@�ؽ~v��_����mu��	~�d�fNA�⚜�zo�!l�p9hWU�O�����.�0��w�{}q����L�0�{g���w�+�vdߓ�&j;z�	��fmV�+i�H�����hxvU)�k"×z�!�UW�ƏJc"�̎ߋ�x��S�D�z�<�D/w�fa�O;:+���kӆu#a��4�9REۙ���T�zu���R�������ڂ4xzbn�J�ȕ՞x=�5�����F�kb:�i�S'��~5��V�{���������m���
����g���!����H�:��<�G�aU�q�;:�J˿X+n=Ð���b6���n��A��cݰ�	V��f�����M"�w�g����U�~�-����׵+��d�Z��n�X.��@h{v�	���K�RC�yҐ�}�=7�T�����|�wue�ڪ�w���G*�[��Y�`�څ���y��ȯ~�fB�eE0b{$��G����u���)���y&qf��r��+�e�p��fz�BKf<���&	����ز��z���ab�[i;J�%c�7'7�bL?9�q�Q��7�X<���R���Տ�+��$�Np�u
�}-���I]�?Xp�Wɝ���?0�ݸC����o�#"�9��+_[�öC��
�����9	����HVOxś��c�������U2��ܠ/x0T4;"+-��P�r�
��u�܄��5����@��=���Y7�}leFG��|�i�ϲ%�/�:����>�ˆ�o�1�����"����G��]}�[�yԴ�����{#�w��U��y6�	�G��-�G'%Cu�k��ks�=���o_��>�"����W���UH����7��M�y��O�Mx�m������Uo�euǴf�p�7��g�k>q��G,y�7�Pc>����)V��H�R����Z��z&��|{��#�C�eS�`ps�[p��ll���"��lF�ۺ�s��߬~wu�ڕx�̌��!!�'�"���D�Df�ܪo��V�J����w�8̌��w����>�k���~���~ב��	����5Ngr����z~�����-�(�۬��ѪW]+�Gْ��y���^#������dvǽ�<+�γ8m`�ñ~�A=��W�]��h\ѿ1�|�9B.v����K��źyGk4���{o\�5#O�oj+v����v��y=�P�>&�d�u���Y���%uЮg��m���޺귘���]7���vC����l��\�o��_
��8W<D����k���ܯ�g��@Ȏ�)��]C�~!�ײ��h.�I�V��B����j��[���'y�+d]n���>����zgݕpf���+���C��9ߥ���5�G{�3ӕт.�|5��H_qKz��{�w>��:�:e�ϯ�s-ґ���l��c"5+��~Ą�o\���aQ����'�
�x=^�3�^ɏUz�ȑ2ӡ��+����nć+��O���f�?y߄,�ű��t�x�mm�/�m�>=\@Ccީ��������۰�ؠ�9QP�x�M[��ӯ�}��>~>�oc�<�1@/���������Wꌁ�o�C�&Q�{v� �Ƞ�쬸f+ԍ��fԻ4`ng�mg��mZ��ޯv!
��'xNG����|�}Ԣ�lϽ7u"v#��jDo-\�S��oR�ږ�~����o�A�F����k=&rɿO/]��L�������ኝvw{�z!<���C�mH`{}�[��z����y����������]��C���|rƤ9K%���=��ޜ���]7"�Ҹŋ��=�EoT���Q�U��
��~���W�kڵ�Q�u�M9����S�gW&�9�L��{�1R�3'mv���.�3��N.1Z����Y�Js�����Gݲ���٣̔�^�����G(a��|5�1N�:feɏ���� ����I^9�	�kl7�ӳ���5:�5�?W~��w?{u�>��������W�O�9ѷ}+>���S>�~ɇ:Vz�$��ޜU��o���_^���2<�d[;`�+f��}A��ػs�.9�`<�q�y۱H���GO�Ur��{��^ܓ�߼�߈<�̜w��'��dn�$(���".GVxQ/7b���UF��j�s�U����OBX�B/���^���_��+�S�{a468K�OA�f���򖄅^�R���3Qg�6����!��q�S��	��q;5=9�wY�e�<�>�7�=;�ǁbd#�2}U.gb��Hͤ��דHd7�[���@���΁#ǧU����=!�=>�i��N������-�"d��e͇M�Ϙ����ϟ���oj.��O����g����R��qީិp����9ȁ��QP��Z�o�6ܪ������E#�H�ACA��� ץ���X���^{�y[�[<��	����vC�}���.� �����F%\WZ&I�jTH�R���y�y���h��!$I?�BH��!$I?�BH�Y	 BI��IO�!$I?�BH�b@����$�	'�HIO���$��BH�rBH�Y	 BI�BH�I	 BI��$�	'���$��BH�i	 BI��IOHIO�1AY&SY	�i2 �s߀RY��=�ݐ?���`w��
EP)*
 JD�i	@
RRH*@���T�JEP�E)7wRp] �Ј�)(-�Ł��G%H�� 7J$�(���.�l)TEbU�����sY�����Wwt��;��k�)v�
�.�PD��;[[j,rP��� ���V�6ff��Z�lʡ*�l1U	C���*J��J�d$(C�0("�i���E�5 Sp�J(H�JR���:    4�$�*0      S�0��*40  ��& �0	����L&i��S�A*�       �`&F F&&	�bi��ID���D�5'�����F1M�'����}��W���� �Ɇ)	 	�?�%!5!$�@�I	 &H1! 0��?��?�?����?��`M� ��O��� '� ��0�CH@��>.=���j?���?/g2 '4����}�NZϵ>�aŖR����ϳƪG��k��
�(ܗb�7�NU-aǎ�j��-X{Y��ڎ�bv��B�)4�"�7%�VȜ��J�Ug`��Q�X.�Ё;ӹR�����B/aRx��D���`r�67n�CYqm���#M���3Va�*��B� �F��ʎ�n�ךR;Kc"��͆�5�zu]ں4��-��E��bD&�J���X��b��4�d����v�W�2�ڛN���R�r�(f̫`���,�SL��Z��d�*4���T
���S]����82�&ɴ��D�1�/�i;�JZ����2�KQ�5���۸�*�2����jb�Ɩ�N�2�f0u�f���Pmmm-�e�Q!Y��$�mbR�S4 �˫����ҧ�n��&�U^��k���ą`AU��ap��L�I撷u-�Z�x-L��kp�=Ѹ��[5nY�弧Y1!`k(7T���H�2t��6�e �'`1�]�m�%&]��,����8�%c@���,-�#EٽQB�Y��ɥ��L�u�ik�����SU9SVC*�6|��$Z�700��������ԖTǶ����%StR�3��.�F�Fl7��'l��F2+��l1��*�G햶Ma�9�I,��c%�Q`�Z��@(f021x]�Ĩ�.YZv��8�E�s*�W�V�xn��Xy�$8���r2�A&f��7��Ĩ�AŻy�^�'q�#!sr���*@틽���[p�pU��.�4�s)�͈!>����m�R��+\��L�x�bnb�z}� ��z.j�tNT##Tn��-6��ڼ�3��5Y�neK{D,�.k9��p�[�k٤'�I&Z�1y	%�n����VǈȦ�eD���V/p��مC4�Ra�p�(�`Wr�!�C]� ��Ōz`q\����t�\x��@��S.�3/5�#���U�J���>	^Ӈl	M�u{2�<�B�r��֗��YL��j׳e2�)q�WP^��`� ݇j-e�^�ѵQ���ɤ����E��ep���6	.��7�m�M�f��*�f���:w�D�8��ZM(PGo.����kjm3Ŗ]��HA����`��om�X���Zj]�"�[7�b�hǵ)Y�U<�଑!�4L�7u�O�L"7e�ˤ#������������YG~6��*�酥�ӸQ����l8�lf����,M����q�4a"#�IdU�В���p��4��8RT�c�0��c+t��l���=kp]�,	B���TY e�7��K�DPj�@������m�.�x䇁�R��N�J�&����C��B�H�ܫXp �'+��5��ъ��Z��	�z���j�#$+U��k������Ϗ/чI��)�{�R:����a�_�C3��7���u�w�6� �=s�]����m�]׽Fv�M�x�FZђY��*�&D��M�s:�@��^ut�M)���xЍSV� 杲��_��V;W_m j��ow:9�P����Ŭ��-�+S�ٛ� r�rk����HM�r��C)�r�tq`�ܡM�HY���a �}0�RD�%�[��4VT���
���:��.��&v��k�;
�z$�ޠ��醥gL眍���]8��%�4%�T�E��{�_v�ga��Ɲ ��t41e��qe�s���uh�`8 �X{mb��yMEh�۶6�m�Si��n�����:�rtF�+s�>ސk���⺖�������=ؙ:I��(,[s�|�t�b��h��{��;qvA��gj>�o)vRV:`�:���H���J�:7+ƌ�����X�Ԫx襹Pofk�/�jJ�<c7*(�t��a0�l���Y�j�[oa��l�(f���3'n$�:3s!��w�I�;r�*\S��I�ν�S�vG��D[n拰��ud[y9� A-�^r��z#�0�u�*�c��uyu9u+(t{5�9�&0����
�7vW�N��o+&����6]E2l���b���	��e�`/�RO#�����璔��W�j��a��j�o;p�u�շf^�B�����OoF�q7�i���N�q���4�N�^ڷBV�y@r5��Ϩ�e�u��A����!�O�ȑ��+���;��:CO��(�}��$��j������|�w}�:C�vu�1NU�圗%��A@m�\�E

�T��L�@U��V!��ɜ�݅AC�Β�����/^���>��KX	���f>]'Wt�\��;y%�A�rn��2ìw�-͵�%Ի����(��]����tS׫7������"�� ��WN��:������/o��gL���N���g�
�8�B���Uo	RF�g�V�0�i���f멮΅xҝ�i���Eg��k&�T_jX��&�{u�ڥ5q���uի���a쉋��z�ӣ4E5>�d�{l�|��$��rM�������hp���v�*��߻v�����]����g|O,x컛��r��K]�2q���� n�:�N��eA_B�%1R��k4>7%mq��,��飜�T�7���g�TX�J �n�/z��:BV��Y�p��N�0G��SmȦ|��jr�ܘ��ws�x(�%s})��^!�ͮ&�U��cO�o)���t��ԋ�u�j�N��-�OJ��97��CunƦ>p�-�VTXqr|���*�D��oT�pH6�����νB�����0g[1 �c����:��v��������˓�[�o���� $ '�pL�q��	��@>�r|�p����gG��Q�]x���7n��F�F4�<s׶��x\��(] mG��2�r�N�LQ}���.
�Kɫ��quk���g]F�"�K��~s���嘆��������mƶ^ތ��}p�]��[AŹR�\6C�.�t+��b�=`�`���!����Wۑu�*�p�SUpr�Yk���Bh�3E�D팡�kSVP}����`,��qdV��oi3����m�+��~���q|3����K�g���*��%��s@�A�k���w`b�a�]"��K���Ô�H.j�J�:���N���Uؗ���ˮh͚�b�X�V���X�G: �Tr�V�^�I4|Gn޵(�mr	����`��eѰ��)�ѹ�].�w�m���{D]����v��
�1���nBu3��gEXy�e��fb�j�˫�3���ݴ��e�z���'na�z,�n�\�h[�j	pn^��+�z��ǹk����2�s��-�:.͙���)��um<�lЩ��}M<�l���r�c�U0��.:��=�����Av�eC����&����*�w��R�b)����٫�7��0EiżC׏j͠Fީ�m�ǯ����)u`��Cתܦ�N=o
�`�{v+�H�#l!#NҤ���ԢWp�	��:a�w9wT��m.�7��\WR��Ps�z���u�'Yy@�b9�"�^:O�"㽙a�W��uN��YJ޽w����DL�-�%U�r�i0�z�î]�$��|���V�:cf�ܫjJ�|�&��̥����j����� �*��G�-է�Y�l1���r�]�Ҷ����"�;4��J}ç��Wem�<�٬����n>]��/r�H�[��l2�YpD�"��Y�*���p���H}�3��o�4�������gR���Dw�]K#d�vwR�<+P"�Ed���r��硁�K���Z��\�VdK4�X��9wR�O�Fwn\�Iu|�^󱧰���(�hpJ����0�ŷ��W^Z�K�w0x�zw~ʵ�a�N�n��m���sNq�؈��̾,rf�x0l��:�6Р�]�H����:F^�אo8d+���Qܐ%�I�Mټ�M\'�nn�U�L
�R�����M�->*�i�*�D0٠:�*�b��\�RG]1Q7���+��e��Y�9���[L_.���>�#e����wy�b�>���C���3�� � ��mf�\�ҫ���yV�Z�/�^s�{��z�4��,����(�˔qr]f.@.�Ю������M�����p�戲d�b��|w�t�B���{�G���@i�Gkb6��h�MV����/��mʻ!�W(�ִ�5������j�����p��L�I���t�r9�}�N�	� @ �� y3��Kk�XS��}�_���30�Y��0����hK�I���d����u˶�z�J�Ŋp �;n:޲@�qXZ��,��׼k-P=g"���+U�Aj�:G�)���e���Ug~/k77�i���`��C�W���ALw!�k/�]I�������U��n������w�iF
�V�S4�qF5.��f�4�WU�I�r�$Ӆ���l�(��Z���ޛK��jk,�i��T�u��X�+��)�����[��2��UL��������=����3��L��������+�e]����_��Ll����8odNf�������]&V`��'�%�x�(U���B�D{ʤY~����zIlZY���+��p�O3�?4�z�������8��j:M��㑣ӻ���w�z��gq�
�����דP��q
ne�+^;���vs�����^�8R����ē�!�j���F
��k�o�[��;��=�"�b=�C;������=�4�JG/��~$��e���c󬺘2��b\�a۫���}��ŭ���}���
��r?��U���v�uijQ�}M��"��^��ʱ��e��C�̲���WVN��T�������]�l�<^D_�P^^6��]i�~H�Z��ҭi[�>��E��^���:�f�����z��ez�w�ֆ�N�5���j����8o8�� �{���}�-�Lt+9�S,�{ۏUkݨ�έע��(W��>�6c�z��t���%z��:�H�����E�D������ے�u%F���vU��:���pl����h���<cŔH��p+����ܦc�Um6G�U�;��ױD�@AX�,;UW�.*d��@vѹ����F ]`�,��Ouz����G��fQ�܃�Y��ct\u�V�[��8��vz>��QF:��ُ���`�n��{������4|�ӛ>:1[��	`홊ލc�罋�z%"HP0�uvxe/v��w�,H\�]]�e=��`l����+�mΔ�Z�5����X���������צt��Q{9����<7F��]�o{~�h��&�<Ys:��Z�l��t�Ɠ�kNGk��dZj�]��O����{7ڦ^��Ӣ��m����~�V�{o��K���k�Oxld��yޛ��ɵ�����^'Z�b��Yjx�����㷉����3wX0Y���{�Cc��ul�Xٹ�=yO:u՞Ί�C�bDY���<=�`�O:���9?�p�]NO�ٜ��3�*��ڎ�=�fc�n����_L�{�*s����rOwI{�o��6����4)
U��6���ף�ːś��7u#����B���z�p������WʏZ�ߖMse'!�1��;��u5�k�7ox�ҹ�#�]p�5��x�6:D^���\�j��l��$�e�U-�]t�������/Mgk�&��ˮ�eǤ�8���\�`��:���7z�u'I��ݼ�uyS��S	�b`M"�p�k���'��|���j?���8˰2��lf��2R��6�U��2�y���%��P�:X-X��#�&)Ö��ӷ�`"�jʂ���Ne&~1��bf]R��r�2Yő��� ��GB�)2S�pf`E$�b��36�J���@�@Q\�µ|!�mQL�L��ikI������Zۘ]j�:L��ѩj�V���nSUm��:���Em�3-j�Z"ں�ĭMeU֨"i֒�YL�����AX�f9K�h;��倫C�������P\�e�$ΥW9E�V'�B��3����uO��LY}���T��/��}S&�B{C�;��G<P�Q�j	o�h�e80���B��v�����t�WWCR�Z҄�N�Ys���v�i���[�v �r��5G�:��e]�rS���[ �;�==^�@�1��Z��)�:P��'��b��Ǔ��sB�l�`;TT�/6oԨI�nx�o�U��S2_��)�	崞�r��d=�u�z�	8�N��.�D�3T�Ξ�"��������<��2�xvӃ�r~�|e�X�2����!j�㢘N��~�1��jN�v��A�D��_kǫ��vѿl����"���h���>��^`�Myw��ex��鼞z�e�ˡ~��w0mn��}�:��'I����$��x��	�]О�,<0&Ї)$7�ﻮ8$"�Iިxd��:@<��I!��ǝ�� hH�9`NXm o�!��;a�Ϟ<y�x<�F���US���&�{�'q9��̥�[�=�ߜBP�Y �Đ�gv��<s��,�i$���d���:d��sְ��R�C�I�B���m�LB0'�Hs�$8d��I޹�{7$8d�T��m�g,��$6�5d`���[��i!��m :�Y$�I6��!���͒H0�ᄞY	� i�!���$8��Y�d��<0��RI��Hp�BCM����{�̐�RC�	� t�&�I�r�O	8`2C;�^w	d��xd��RB�Y!u@�@�y�:ץ����{{��&9��\��m#}i޹L����N�g�hC"[�o���7t���B���Um֗kvg�
�T7V��fN>���f��s>��/^�-�m���i+�~t4�@��F%C��(j@�$���|&��ys����,U�V`#^_�����;J�@ly}� ��i��U�A�0�r��`
X�Q���a��2�w��-�R��5����l���˯K��tԥՊ�ϋ(���*ڒ�X�G�>%�{���u��Df��Wl�%]�n�T�����N���˘���U��8C>�=�����z]��1:�Q��S�%��`Ӟf��]��ek������6G�Bmy�I��]�:����Q{u�ڶ�ZǄ���g�e��p-��9�]�l��-g����"xQ95�x@���P��c��s�Sr��-�c�ҹ��\od-��|��T=�n_�R�<��ۆ���T���j�W��#(]�Ɋ�Yt^o֓��*�a+��!�V�u\�U(&���x'#�*���ec��?g�I�;���(>�t)�k�{Y�WI���/w^�+c�MY˟t��7�!`�a�)e=��z��Pu��Yґ�6�
Y�F-ڒ�]�hn뾛[*��l2Sհ�(�����
�g��,#�U�}N;��`��v�ҨE�׸��Ȥ��}��y��]�y�=����� � �s9Bܖ-�wY3h��T���j�K�0�"���)us+�T����2&q٩gV���[)�����q�,��)+,ӹx,U�i�D�6�*W�B�]&s1J����*h��DVVT��U���=�B��?İ7.V�8嵫\���b��B�k-mV�����R�l(�m�DP�TcaZj��JʅB��R�m�"��V�T˙uB�`�č��Dm��T++0LDF��xmߞ)�����*�T�z������:�~n.����l��˺Z�I�6%��yU����Aj�}
�z���
i�y��C�у��̤u�H�'��c�*���ǻ�I���&�ئ�ru�>����=�ۍ�'V��� Ctw�t\T�ק�X����A��s=;��`1�!e	�=�ҹ��sx�VF���8�e#����7��4��~�5y��_b������|n{+�-���t{7��0>+���3Y�r������x�Kߥ��˴b�
���S.+�C��/��x��r�=�7�{e>Z��k�֮�j��)uIn1�º+*%V�ß�z{7ўٯ=۽��~���rv�g[RN9?_UW��/�b�E�\x�ⅼS�O�!�������T��s8��&1F�e�=ZWo= }~�y������h�[�\9���R�~�ķ���.K<�k��FiO3�%�"�N^��[�L����I+��0`-�8���ɸ��w�(���B���;�xwz&� �ʉae�)��/��㹔Y׽g��}���f��x�T�5��-\dʃ5	Iϳ�ޣ������>�󉁗�6�h��.���ժ�gwѥ��^�a�ߐ��)�F
��>|7�V�7A����ȭ��f󮏥��M�����z���/~gjƳ�����:�� ߖ���Rt�f9�BPx�o�EMPF_iN��mi�[�;i]����Fv_GM��D�rL9�#.^�1~Ʈ⾌���&���%�dC8_�n�~�wm���.i�[TG�}����Ӫ���OB�#�ݯ�h��u*�e�p�+�CV�ڼQ܅��i�,Uj�	In��|� ���c=��_����W�����v��`�粤�Z�i��.��ͺ4�)gzԞX{frc�eT�謏����k��,�^�.�����y�P�MvC��  ?K�b��~1ۧ�Z;%��o𰑊i�:�� ���r����H!���3]I���ew��Ry�4���%:T)y�&��~9]��
��W���yK����q�?_Üt�\{8���`Ք������:ǵ<�' ��{����4�im/��P��K����}�`�/ZcF����'�w��S��u�V^hÕ�˚���Zj}����9��an���D@�X5v�����WlQ[/G�b���J�ʢ'Qgox�$Ԗ��
τ\��Ī�״c�#TۖWq�J�-uj���4w��o[�S��i4�+yZ{5�vs�����8г�4�6��:=����gUjON}��gz���l!Qe��n����X�s�1,��1� ND����'7X23hVd�,F�)�7J�wM�T��]�X�T��G�����D`I�-R���&JMI�p�R��u^�zdY%b#l[-*�mDTe�EPPF,R�(�EbfX(*ڵai@��mR6�LE��TFTTe�E���J�KJ+eB��e��H�S��+�b����������U��-���}���
���2��d��o;x.���뱷FXZD��V�S|YkYɴ��dA,a�I�����/z�=3o��ޗ�w��	��z��w�3#�jX�pjx.C��Cp��%l�Q��
�R�[��{:��vFʡf��ao�G	�(�i��.�;�fnq�C�����,�30v���i7H��=��4��JZ�^�Z��5I�==TDaf��:���&'�0g��
�zߎ2���ֱ��q�z���lW��<�ml�v�91u3�e/z�_dO{�F�"g^ؕ�����|4�o�N�s/>�9^D~��Y��/P��\xt��ǽĮ���ů�f�uX�xގJ�{%��y�r|.z;�;���\��|^\Y�g�y������pfz��i�W�p�C)���w����\3{(Z�a�_}���Q����F`쑮Z_1�q"�ٹ��)mπf`;�}q�����3�$�o�7ޠG��-o17^���\e]�='bwk���^tۚJ�p���0�jPz.�yj=�nW��;��ҝ,�ѣyd�a���(����Э/n��.�xGu��Y�4㰜�^���0fl����1Jnjݽ{O�c��%�k�������Ҙ�e׉��}O=�Ri��jP�m�ڍ���u��A�71H���`�\\;F���qq�tj���Ub{�0`)�̨�W�:�7s���<�iQ�£��陘�؇,�����yM�o<��I+�c�)aO"&M����X�s�4Z�%k-�˅��Am�Z�3؂��DQ����.DB׷����@�8�m6l��Y��,H��vZ4��ډ�yW����ʂ�>;��P��˝�O��n�������jF-D4ȋ�w��Z�p(��i�����F�x6�q�s�fُL�9Qul(�&i��v�Վ�N����0�yO�]uxH,�|a�<'WNM�C6�K8#O�4�C�!�<͡�sލ���ӄ1�;M�V��]��0���1T�����}���Y�L���h��yN[��7�wd�U���,�#���)8Zȇ���N܌��\{M3��T狷�J��D��u<�E���q���������Z�v� �'Kz�$M��Ka�.)�uf3�P۶`��1��#�[���ΑC�Tz�❦�Z�o\�6�0�*o�r�3����t�
¦��^}kr��[���(�Nr�U[;Uπ,�G�����E�����vnXr ������9awH��bF-��DYfxʖ��x�l=Oe��,'r�8-��D�|qR�]Nj�4�tɂ8�e<�
"w**�C�5�"����s|�)���T��N'=�s�����Ir��E�<!�t�t�;v�飜n����v������>��K�5|۹�bL��d���ug�ls`ݮA���k*�@=�
=�o�k?'֭�wy�N��"���fp��WY�1��(w}��C�)�Γ{�1�qS6�'^�A�꒹�8ge������I��I=rnK����fn)��:� �j���c<���>q��
��
�Du\�������j�Q�;lo=�v֗��ߣ��������s�ZS�8����V�6����i�rZMð)�C5e���]V�s�e���!�-����u:o{��)`���zp����V�N���J��f#l�V(咤PUU����m%m(��ѴQQH���Q�K,f%T"��Q�J�QJ��1��V"�H$�ɀbk^ѡIS��*�*��3nu7�t8ab �%8��g#��AH:�:j��������u�9��h[��E�#��@E�W<���c��i��>��E'k�o>�َр�nN#p��g�S�x�oo<C�"�"�*
��\�b_U A������kjg\"��Āc�<C�Cj��m�w|�~�闥U�-�M�fan	���77UFW�fn�,���\=8���C�����,����=C�+w,�[q��$<8�q �ײ2n����%�E��:B��Z���"��!��S�AES�j-$m���%��k���.(��I2a�Q]��I�ql��	Hj!���#g@~���Ep�WW=r���o����V�1]Ʒ)ʮĵm�f��$�ͯ ����,<��V���9��3�9yH/,��|�~x�
��'I1��9��3z���w��7=j6R�f��Dal��q]@��tY�9k1�4�g=�1��r���fY�<�޶m�4�Nu|3�i��N톑��$A�(���!�@��Y�D�/����x����L?M%cb�[�M��5��d�ũO���� ����2}����,Hg,�>:-E3�F�T��zs|�v�Nݧ,��FҬ%�V>(�Dq� ����곐c����$�},C�6!�.l�e�8NS���bt��l�ӷ^)�t��-�P���6�	-��in�y�Y���;2�b:w�!�9��iͣ{{jJ�����b�;i]���E�
K�,���q5��Dk�$Qg,�x�˨�{φ6c�j�`KL;A���$	"��0��'^��_%���G��"�^,�9���e�
��ɨ�����r�$;�ߋ^Si����|��T�*�m�m��4ZӋ�a���heE3��m"�O�DC�tՖ;�	���^�g����}�T�/���l�,崎Y�)������Ь����x�tW��5iΩ^Xm�\l�
�)�ϝ�jc:�a�1��﫣��E�FP�t��yS���ak���$<8�i�l�e.,�$q��й��a�˦r���՝%M���Mqf5b�����7e��#{��ȴ��=�_�Tjˉ��S��~�bt���"��m��4�*��Oo,��'�IӦ�������<ka˴�l��j��<'BAd�{u�8|&�l��Ζ6�m"�k�"�h,7^��tg�|�o������8f��4�Hq�6��6����4�-�.�r���՗���[Ow֯�W�4D(�朐���K�r��/4�U�> [��G�0[�7K�a��0���$I��"�)˒Z���"*�Qh"OF�3S�9j +�j��\���XA�̋A��](g��3�LA�Q6��>8޹͋�9I��v��\(�6B!�war��>�<��8`^�֦���:�����3��2bw��[W��]ζ�2�N�n*�ݽ�����^��a��DZ<�YFC��)�f�,��Y4p�"�J�aQ`yØ-P�)'�進vY���-ś%�>)a��d(q$6�޻���8Fӄ�v�ʜ��i�"���SL��=��`-Ų�	"_8��ål��K� �I����ۧ�l��6��(ʿuxߜ:k �ꏃ�I��
�}Zv'�����8U8�8�%8g�Xy���	�I���u�'p�����;Jq	��v�&���Lo;Ç��k18�Y��Q׌uy�tp�Rp���Ӯyw�ی�ӔX�5���7���qxִt��@��!a���YEԉ$����	��UƬ��W��K}�F���tѐT8�_�۱�\�{t���`mt�֑u���V��l���Gtɵ0R��xG#�;���	o�o�����c��i_X��ϓ�LU�ц�oL��qDj�G�(C+A�;Us��s����/��$˾@k]-�^�,9�S1�zv�:���^��On�5+�,å�����*d+��1N�h-m�.�j�s�U��Ea�r��2�'݈��)]�̀�k���.��,k��_b�Vd.����
��g�[P��/��y�/(�|6vٛJ
��][�CO"K;!��d����'�VRF��G@�l�9֛�zj;�+E%�%���Qm(�8�,U�D*˖�1���X��[YLh�j�1�&9�b�\�"�"���������s�:{SSn�;��3���,TJf��ϣ*�q��͆��M֦�2E�.-�4r�4������}޻�,e/���?C9��ڻ2�B*/_t��w^�T�--]�P�ǜf��\��(c��	������u�;2��i���^���i�i-չ�n�Y{.��3���c�=�^��oVs��T����d��N���;oL����Sy��.^�^������ܯ$��*�}�KX1���O_UѴ%�����ao��΍p���=�w�'j~o^��y��)�>�Zx��Y�����-iȈ��w$�U��N���^�u����S@�-��Ӣ{�/��g�����lf�(�꣩!.v�c��?��:��լyL#��ѹ�|M����d�c��H�o���]M5ˤ^~��\��-
�p��(�bO�ۚ�u .���U�c�ǃ�ȿ�V�_��&��vF'��u�[h���k���;��35v<}B�g�I��s�����h�f�r�,��%w�o��;3�fS��T�J�������,v�a�F�U7�BӴ�e�MV�e%��|�g)��ʽ�He\*��s��4 NأO��z�������<�w/X�sz��P@ua�zZ�0��C�f߽�/0l;�ہ]֤ks��S�f�K���S���Zit��kWG��I۩:P26��ъ���Z0`%-r����N���
ٳ��eU�}�f,����w���2{g��)uQa>��u�4��V���ۗ�f�i�>n��A\>���J5R��;�O	���`�	�T���@�,�Ӯ��n~�pg�����X��5)��{ш0��G�K8eא{�H���M�]��3��)S��g^j�=!֩�3b�:�I�vj�+D�ս�CT[��J�*��y�}2k/y��'�ܡ]B���
��0�0�����.��8|����F���7+=�́��G�.�^)����t�X50�j�;z�F��{׃ȟg����K�Y��ѓ������U��Õ�^�F����$TD_��?�9�&�TҾ�)��x��HO]bS�ʻ��䈍=�I��k��72�Ċ�+j̋9�p��#�/!��}jMzr��\��@F����x��:)�3�O#Ԩ_QW¤�k�=�Dh��a�^й\�-�K;&?�WIٓ�w^�Qp��ޚ�޶����{a�F)\��ԔW����,���#n��՗�3y��7����J�5f���SQ,�]rZ��Y���Rc��Sᖱ]���(".�nr�ʸ�� G�.'��<��V�90��eѲŴ�X�����k2"�2��S�N���5,�Yf�IjJu��n�f}V�*� v�љy1�������fZ%Qf��WT+�2�%�-�ʑ0Y�e�8��	��Օ��ID�8R$�)
�r�[iU�B����-����(�V��
�4�110V�eD�" �lLZW�ҸX���UG[h��6դVю9L��V�q�J�_�Mq����}��\�JuC)d�}("��V��ߙ���q]��ޔ�/�!j��|P�~}��>�=��HH���P��ߖz��ƎvT�p�A�qڑ^��k�ŉ�;6��v��%���jgΪpH�z����3v5G��g➺�J�ˤ�X)����xi��g�e����Z��x}��:�ȁ�����or���J`�⢮���gz+������ې��.�P���A]�Z��Z�,o�gNK�W�����g��o䶴7
Uf#�tn5�ʯ���V�������t%\q�h'Vl���{����`���A�H�V�vV#Z"4uS=�3
��;�Wi�|�mV�C}�l�+��wyN�f�0��w�=�;/t�Ӭ�=U把�w�CޛC}�<r��yNZ�S.�y{sp����ڏ�S������v��p�[���0OM,�f�/M��[��4^�ce�&�C9���'l\�.Gی��(k<=��6�Gڒ�|f{�͙\��o���s`�Y�'+�����oF�1Z��d�i���=9��mp����`b������٨�A��/<G�C���3�gH��k��;�69}�m+^R��B���E�Y�f%m��F�ٗ����[���:�ѥb
�C��^v����c���hK��V�4m"8���,(���{�	2q̫k�k<���<�Vmo{h��b�iҒ���s�gt����2�k�����v�޵}�Uy��m;���T�2��I��s�Ck�g��-��h��!7aVW�l���зW/�� �����t�8�ua��v���X*�V��>X����3�E���ЧǼ|8��XZ�{[�kB&�ӋM�a��Ȇw�^5�6M_�m�L�Jj�/< �9Z�s�2iVz��I���O6�۹F�Yk9	7ԩ�v��A���
��m�u��m��f�L�S��7:�/�j�(�����{�^���z�β���O'�-����*[z�K�4�	����k5����e�^@4v����oa)c�6�!�˕:�ڛ�����Їu��ܺ�c��>���{ɜ�3��T_7KYc�6��f���٤�r�r�ˍ��^����{z��>޳�Y�2����)x��S�pr��!6��y�<=���I�M�F_�_B�S(
�v�ܔF3l��9TrJ��1��C�r��ȖR������<Q�GwPdSq��]�i���תn[ �t�l����O>n���7:Ի���άo	��9	r�e&��:�v7�	E�:��P���2�;t�T88����j�XA�o�a��\xy�U�x�<+�>�q^a�i�{t��F�-W�:Mbut��T�sl� .�,�N��@�0�Ecy>n��(P�Z���H�N2�M��@`d;�E�%\�c�V�\,U��(��0�ݐ��2�ܩd���t]k�WA��TBSS�(եR���)m�*�̵�Ъ\kGm�Z�,���ҕƬqKr��qh�L\�kP�FŬiiJ��j���*�Eʕ2̕�h�m��8$���SE!���5M��K3����?>�b]�h�8efL��t����:��a�~�o�3�|*��1�9;��ܐ����Ү�3A9B��d��7*q;�٢��}����P�N�vY/^�@�}X��Z��y�������Ef����%/|��7ᷡ�&��ր���% PE U���¯��,�j�{D'�2�=��F]��{:=Zx����25� ��o�����x�z���ys)'@�����������%�kj�=�V]�b����z�S.�/� vkY�YB��>�!o�7��E�(��׼y���pB��t6S��~��X�z�X́�Q�$Z�0n�&���������~���'?S��t a��h��t����6{��7�����D>��:Z�N:�y~�&�mT�q����)�-O]�-�L���j�b5��!��k|��ӺU���ivvc�[hw��ҁ��_�k	��m
���w�y�˵%��&�w�~�.��V�������S�����N��y��ԉ���	elo���O1@3����Y�{���dV٤Ue�i������b�
��3��	+u3V#�0���iVGP��NΌ�Ό$�ӆ�ד8돻m�^8��U�Kٶ���y^��~��̯iYˊ����ɠ��@L~<��>G��w���&�\�SCX��������7����ry�|�N��/#��]S�1J�:��Ի��q��w%r��F|emu<����k]�y�G�f]RY��W@�vѶ��ni�Z��S�b��ڄ���z��1�z��
��^њ�v�U�s��V�jܜ][��A�� X}dfj�WQa7��ʙt�]�g�����ᶹ-Wճf��L�`�4�Dg:�g���2�͌�5������x�����]=���F�<���j����<����-��0I��j�\��#v:�T��5� �>�i��;����f�~s=�1�y��AQ�1���5[W'!�Mw��O�nR��Q���7DV��26�G)�-y�*�9w����]�V� 	�#������sg��B�6=��h�ܮu6�^S�a"fyC5n�/K��+ko�������+�X`�..�5��#[��q󵶑t�͖�pW����f�J��Fn玔ú��~�MZ��'���OS� Dξy��ȥ������߰Zusש��C��3=���}�w*��vf�lx$k:��v��-�CP_h�4%pӐK��B� hV���V0s6R38MP����18��q����5�@�,/h@[ɌPTbxk�`��7d+ �j��j�)�����sv��J< �`�Z�*�c/;%�Ү�b�H!�;Q�SH�f�Ѣ�˲n�a�RА�3�	P��� �}y3`L,b�x�0�7Q:#%��9c�R��h�]dDʌdͫ U(�TGƘ��%-T*�ŕ�q
��e�R����ZŅ�B�(
�e���P���q����UUTV%�X,A�����V�U�W>:�T�=�"tٝ9oE�U~��WȨ��N�ތ�úU�>���J�3/�	1,ӌ«/���2;���ݵ�u]�XW1[I�[��g��}j�M��j��3�s����] ���fכ����'�7E��ͫnL���cQ���{v��xvn�g�LƁ�\\�.��y�d�bK�e�z!I��t�|ӽ`�+�Q�4���:�ڷ������=���}��^r�ԁ��ʛ����;������v�H�~�o3
�OzY�LR��U�����e�?_�^���#c�מ�	󹻙\I�\@n��:���t#8���f�mО�f���iU�z�Twc��.�2���{�Ӎx�x�
���1��=|VQ�}�ӥ�{��l�i��{�X3|.,�iP��|3��v`B�1�+���jvw�����GeL��.ضN��O�ؕ��#���ӔR�tk�CG��<���]�R(�a�q��MT-�/��w]�в}1���@N�H8v�:vw-�������n��wk�%��P�'�w�.�ϲ��2�fR髐��x��$4n�|N�%Fq	�I����sܗ[�R,�gUˮ�\�'L�.���K��o]�T�ӷ�tx�ln���	�����#�;'�i���w�����h,���fK�OůM`�LضJ����a�)�~�LP:�����ߢ�U~�K�`�����2p���I��(7]�ʗ ^f�ɥ_��m{jG����}W�,�ea��A�Pf�	[k����<��Ԫ��PLѽz`\��bK\�:��;7$8^�TE��]p��×-�;n��$�|�ĥ6W�fj/^~���,�|5�~e�#m�~���9�R�ӛ�����}�>M�;�4�Iysk��-����r�y~�oH�"��߆.}:�o2K��vҎ�q-)[��/}�x�Z^��"�c�L��0�1�Lꬆl�`��z�ϫ�j�7ZY)꾌:�j�����ˉ�^��1��z�%Ji��T%O���Q&�Gj�
��o�[C���I�#�<h�ɒ��y5������w��r��Eb�ckB�g��x�v5�ك����Qk�:~Ȳ_�TΙ�z��*����U�zێ·a�7��b�0b}2�ly]T-�t��l�6&���ub8\��>�<�dx�zp��`��/��z�*x׺y�����S����L�m�!\�f:2���Wn����n�0�O�鵷:|�ݼEά|N%�*�*rS]��<�40=�Gi�� cs�0�c��T�Q�{	�)��2ը~��t���gv��F�/Zw��Ɋ�S��Cb��7;����;�b<�]���R]��mr{�����B�W���ds@{6�j���%����/L��#��ed�b-.[����blVWL�%��z�.�29ᵑ,۩�ӥty�U��T���w�j�I_vK���u��tnu��R��*.U�Rj�P��eL�	$� ��!��4pR��ը����iZ�LJX��H�0�J\q1-��UAĠ�[V,��YU��%�VX-��YR噔p��r��M*�	a+tTŬn��{F���x����<4J�Lk��p�I�2���0k#��p���]}|���
%Z���yҹBb��oZ����e��������y��4�\�ץo=oҎ�`�zG�>P�x�&b��J�{3��j.$��3��. #�R�0{{7B����M�i�������yb-�^xz6yX��&�V�eG�,�������9�՝	� ��;˺`������S!}��NR�NB�*�y�;�U�|�C|����-W�:�:�>a�+�{���折��!�W����\��1�<�K�d�9��*�;(��d� dcp��4<�+jI-�[#�̩������+x^���~��:�cH����Tz�[��&��A�m�n��rp(Z�]2�v���f�笿>l�e��*�Lf� [�w��1��n���h�;�=	?D�(�⬣��P���I�i�B�����/�`fn�bݽj�Op��ps�'VWy[��G�r' u�pok�����f>�;�nJDm�z�D�4���73=�ks	�wNG~���˺��'N�uD|�ٻmq� ��o1�S�!�bj�m��	{�`�Z�Kz$����uݏ��9����S-{3,�9.j������o�Oʆ]vS�0_�s8*6F����R��ٕ�+-̼<^[�cf�٥���lj��V�լ�+�m�{;^��e>9L�F�YO�1.��%'9��6&��<�����`�F�w��vGLa�n�׌�k{]��]+B��%{�����]�^U���D/��Q�Sss��+r0���sۗs�B뗴ff0m�����eJ�;ޏՇ��n.��	=˗i_9�'#Z�8�Y\����a���Y�׼��^������`�;�w\;V)���*�X��l�n־e��}S����Z�t��^����g:��#+�*�ׅ��y��['b�2M��s��9m�����T͞�.��G��票�Imd�N�u�*aNa--4�j�z#�l�7�Q�����s�%+&�;������m�Sf�x��<�"V?s��]8�Q8�xU�L'f�2.J<y�k�ם������t�{���-u%Q,H@�2���:G��Y,=&+lb�٣=���̲�ư-\bW��_�b+���l�8�����>��T�R�UU~�[ @cO�� ?�w @y������c.�/7Ӣ����z?=�ׄ:B ���xk��6�B�n��<!�����њ߫!6�K�ā 	����o��_w|z���a�=�9�{���{��p���Ӷ����[�Z��g��vcB �
l�3\� @x���ߦ����I�@�$�$��@��,,�}G������C�����	�C��O��ο���O����O���� :��~w�d�>�*O;&~GD���38�d����$7�~��$��u���� 3~�q�C����������q��!'��� ��C]��h�����!��{��qҬ�{%0��^Y.g����=�����G�� ='�B��>p����q�I���P����:�����y!��W�I���9�?y)����ǟ�q�t��,� 	��Y��$��퇫��?�������pj�ޞ�=�'�(r������8�>��p�ɰ?�������Y��q�}_��g'�� =s� ǯ���g��OMî��X)�XS���|)=P� &�� ?I��'N�Fe+d��5�����G&<�'�p� ��F$��Ƀ��3�z�`B Dd�I��$���6M~����Z�	���7<C q�>�f0��of���� ;�_����Ot=� G_���bA�ϳ����B��Ǵ��p��Ol0!������}(����������a��� ~���^�C���� >��=����/�K$�~��A�H �O�a�������;��?�>_��z��=�0���<C�Ñ�d)������z�o�'����o������ܿ������w�=��_\�l� 	�|y���}��9�C�>�B���z��x�B{zS���Ѱ�%�$���� � ?�$���{��}������$ '����d�5��}?M'{�����9������=B(O������	��9��rE8P��Q7~