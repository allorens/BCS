BZh91AY&SY�5�yߔpy����߰����  a>               $     � (      �   3��QF��{^\| �@ }�U*�� K�7*�w�5��;�c��{=��t�zg������l����ϧ W^��� {���Gv��r �Ԩ��o��:�ݏ�<��s�ѫ��������� ��z �е7{Ĩ��>�O�(�a���{==�����ǟc���y��Wa����|�](p C<���܅}=w���[ݫףT��������2�o�N�rIz�jx ΊO�8v�R������g+������ý���o=}:z�ٯ������`��x0�5�x�;��W����������f�o��ۻ�z����z�n�� ��a��ѹ���^�����n���&�}�on�`�<�^�!���ޞ <!{����k��sԶ������ͼ��>cĽ|���jKZ��  zQ�Ɂp�� �:�=ϯ'w�.Z�s�>Ǔ7�;��w���z�|��	�wU��9����<�{=�������������w�{�z��                         �A��*�4��&&�� 	�`h�L �R��42 h&C@h�"{J�hb� �dC 4	S�)�T�F��0   �����h��➌SL��h�ښ��i�iS@��T�a��FF��o�}�_qXAK������ӣ���ؠ*o���D^DE��"����2*(/�xT3Z���O����������l=����}�D p?ݴP\^ ���/��}^�"��$�>��x	t�UUU�P�C���7���Wݯ�����@֎#f��t�� �;�d���#Ј�<u ��$��DD�z�N�8'DJO���b"y(��""M�K6"t��f�N�I:'DDN	��$O
\�&�M�����^��:�UhWk�vh�	p�����슫cr��U]z�z@��y�Ula�����r9�S�J�W{��x�T+����t��eW�+kcr��\2��.ƖU*_���p^Vˁ�_'l@�]������.�%j�+n�
LL1"�W��l�v!`^pt���0z9ŝ1���z���ޅv�m}�ܜe�d���
�n=�b!���^�,X�s�@�+���-���T	�{���=�m�{�nq�j����ؑx/�m�o��C�zq�o�R./o���!�M�[C��'"�x�m��ea�WT�s� ^酱��5�zpm���*�PP��"" �Ո������lDؐ"P���'J�$���6"$�b"&�K$DG�"pA�v$����Q%"p؈��xDKH(�'Mȉb:�	,Dy������$G[����%�'�B"'4�""'DDu�6%�%�D���bDDH�tIDO �lD�s��� DGI�:<�"xD��%�6"$�c�K�$�b"s�"lH;�А����""pu�,J$DD����P�B'DJb$����A$D؈�"x�	�N�bx�$DD��#��"tDD��B"#��� �w��� ��{b"pJK"'�Dؕ�8$��d�7$�:B���DIb����RQ$��:""pA9�DD��%�d�"D�I��K)(؜�J; ��'&<z�����>��l7�6l��p�$�C#G8Mi��b�����cB��Uݎ�ڲU�;ld��Úuj�E^NB�lnU�UdR5r�F��͎�U�-��^ˣj�8*�����bϺȪ�t��/I^�]�[�M�y]�c*��0/��+�Z�ӧ��Ҿu�^
�d�e�7�}vpJ�{��t�9�B�#��,�+^<���R�93����E��DC�`i=cK�E��l��Â�l$�I3�6"ON	��D�E1�W����}ƅ��W��v8�j�|؉�vN���@��x%xM��$G�:��2/�N�z�g|At-��"\��D�8��*��	����ȶ��Q�ĭ�O'��q9:}�|t�Ǵ�B�A���D���U�خ�iy�;
�;�`x+᳭mם{O�v�"�OCd��|4-����c��D-�N,���S�^�t��Ye�8^���DOX�%;<t��#�"P�$D�&ĲDJ���'K/Ǆ؉�PK�9���BQ$���,D���DDNxDD�ӣ؄D�J D�����"%��&͈��b"a�a�t��v������Z��͊��Ӧ�b$w+��m^
�]0*в�"��ܫ�VN:��O+�[
��>&v*�Uh^xz�q�W���J�*ȧW��ܬ�E^X��Y����{UN*��D��<͎�,J$DJ؈�d�&9B%�8$@�����H�<Z	"$xDM��""pDI�D�+�%���"%'�$Ux���LB�zаG����_���LD���l�M31VU�-+^I���vq9�:[�NH�C��N�N�(�o�:CᡱI�RM�%�>,�Ŝb�b%�I8"sH���DD�DDN�Ԉ���z�D��DDD�	B'G]ȉ�g=�����r9<6��ú������u�#F��֜�����=	�	x��pAlwǇlx���;ߵOc�ݱ����h�۫_<����"�����$��vq�!�/�&�A��VnK+���p#`�zKJ�'M�=ġ;�P�#�����z��t��S���By=�Lk���O�N�t����-�[�	H�淾t��x)��NOB��b9c�t�4;w�N�b�x(��쒯Gφ�]��{k���$�!lz5�H;{vo��4u��K��+�:_;��)ru6rz'*,�x�J*N���&��i9"""U�bob"'�,��I:"tM�'DuP��N��bQ�g�����D؉""t��D�%,؉R"'HK�B%��'(|@�Hb""[T�ڼӧT��y,R�Cd�q����F<�7��3B�c������ˉi�+b���aa�h��!Onv0�N�����G��|��'���TxW{!U��J�h]�mW��W�ʓd���Y��U{�v���/W�����2¯%�v�����>�m��&�����J��[��x[�7��:�k[�+{��{���Gclv:zzp���lR��jxLG���y��o�����)���k]7�q��N���n��**�	��#[���:q*#��e����h�7�L44Z�,6|�Ǆ�8����}��а�e �!+���0��wǰ^��șayp�z[	c��9qZ��ޥz1�n��=dn�.��֞��!�1������������:l���p�Y'����խ��<05P�)�H-&����BUshp��,�lؽ:T��M������5�&5Z`��T����G�誖�m ��ؑ�|pW��+ǎ��аp�x>�-_
�4��#���C4��i���v_o�D0;9\��cc�ZL��#�]���y�x�W}�,��1p2\�$m'�',O"\��i�IpQ�v=���Q�����#�����_ɴ���3�P��DK�Yo�7
����,g-�O��O�?����IlvA4�qc���.�*a
�i%"S��ݰ��������idR�LB��~^(ɓ�3RI]�Pm-q0���#�h	؁2$��/v׊��U��%b�D!vr�;��&ēHv��H�>�7fЉ�6�4��Jv��#���s�td�b+t[H-?&z�ivA@��/���:T:w��ئ�%�wcXy��n��Lnji8�����3�ߏ���!�y��76�5,��l�u��"��A�o�y;U�c�a2$u�ZG��Y�+��R��ѳ�!�N60���U���fOe�ݠ���ㅔFZ�z��s��L�j]��1�2�8��2�A�tZ��v�8\�,C3%0�c���0�y�f�Vx������L�8���8\�-@�M춦���)p�pw/k�B#�`E����8|tߛW�?)���s�f|���g���c�5��fd���3��^�i}�9�9�`6,�a��	��Us�=�Lz��>ћi��,�홗hy�������>-u���e�"%�	R��;�+�y;������}�9�=q�SV�X�I%�ٙ��A�8���sU�Vg��I%���9�>`�۲��ƴ� $��$[z���Yqe�::�>3���!�McSNf��3�C�R<y�L��(��G*�`QYӍ����b9qt��2���ߖ���L!�:I�̳ʈ$n�lçS8cd�[�8\L�@�*�G	7#�_Er��捥�=h�VN�:T6VjE��Rq�q�����B!�Na�*0�cӐS��f�nt�f���.nR��?^�2kX�L��o�Òp����|��M��Pi�����n�$uHa*ԓ-�<p�
"�,c���dx�ƶ�$߉XZKzm筳��Ma��>�+�	$�ٳ��;e2�V��vm'�' ��.c��x���kN4�$	Y����T�i�
��1���u�1�l�AX�!2O�>�V����Q���8kȡ����dd��ݼ&D��J$\)�,M=�MSZu�h�ٰ(�.׌��w���R]ΡD�ʻ`HH��`���0�^�]���mbV��#�
���g[�M�~��)��R(^@OJH���Y��؝"���i$4��ދ���#iݍDK!xQ��a�|���)�M��I��$��"R����0��)�çK:r[�$�*y��8���wg5h�/��3O��|}��+�G��eb�V_zt<�9���d�zIG
-]��t��i��|t��r�,�BHq�杤aG���7}�xq�,�|x��P|z7}z;|w
8G�9F|�kEp-�����CP�� �	�6�9�I$�4p�r۞(���!.�cyhsl�R������o�c\t�l�d����K�����SD���X"�f��v���	<t��H��F{Rkuz4���H�z�����8/nL<YE�5���ف�ZM5���>>q�{]e��<\Y$�uF�䄵x�+k���"�5f(��دVb�#��l��5a���6�rI�)�&e�k?���df��l���ҵa670�1��o{�A��U�1Bt��F���1:0�tS7-Iٷ�1�<�E�,yK��Q0���^f P�XgJ*�ڢ��	��j;�H�>�E�	{aí�|�����$��h��Cy��Cb��r͟,�ic�[lri���<�� �$���:Lm���A��D"}$Gl'J��
�JQJN�ㅖp^�%�:Q��D$��ɥl��O��²�̷ַo/�����n����6|Ov���y��=z���e���)�f8�P����%Եe��v�+;��ޘd��j4Aa$��^��/#qaeQ���"p����lj�#�.A^((��x��xI��0�l�p%����dm�f堤s]KE-0�f�VG-DY�_6�H$���(��g��26�o &;TmN�A�,=H|���g�{�mW��a-3��nݻ���񝬙���$�%�I�� ���ٹ:I5��+�1GnI�[X�E[=lr�[�ŷ"�x`�U�TU؎�
�fBO�(������M)�,.��kC�!ُ�����t
�b����ń�����[�g��<a�{֑֠�Cz����@a�x7�s��Ǯ ���[�e0�-�ư�g��$����a�쫢��L<�"u�"$��	Y�zYD����[�����>VI�}燈�y>	�k>��,��!.p+P��0��>I��Ŭh��P49i�nʶ��kE��xyt�
l
R4�q�4��\m�<�m�q��J��N޻`�z|I�!�ud��qCm�.)x�鲉%Yեv;[ɗw���c)��%}��:I%�	�@�D7WqXT����+7���^�TE��}�O;-�Y$�}��w�4˵�ׯdNݏQx� ���׉+H��Re���Zmy��;�L�8��f"�Y~�=l�Ğ2�7��6`�T�g1���Å�蒉bs���l+>'������93�/~�Пt��R�ZS�&�3ǟo�(초�O��+Hzsz�:QG���a%E!�.�!YiYb$VXa�o,u��sFf�̻dZ�!�a����8;����=zt��z�L��0�����A��g��9kV���f��x�,nl���ⷺw�r�Rz�V@e����睌�{�.!^&��3�ٝ!D��4�*�^��x\K�I6Q����%�d��~L�6]���"򬫊��٘�IvٲY-�:n� I#R�۝��O��:F�Hs�x��V!�qi�4[��{v�����q�0�T#��̫���t^�8q3ۯ���x�����bZ��2dQOؽ���DkVg�n�a5�x�1�^aN�e�U��"Η�װ��`-	n�^,��͏q�\�hf��Y�ΜX	�t�RA�f�6�h���p����N����ֱ։�[�Hŕ|�瞞�r�-�,*��DÑ�
n��$4���j�&�_Zak&�P�I��O���e\k����m-@���7��vNB�­�_�h揉 �Ҷ<�|�����j��v����m?`���;���W�^��Â{t���d�%�$&;%�a�$:I�b�@�]i�����}��~�����_�֋}��g��Nď��}���:>����~�a��0��85��H1�y�%�����8�Dq�S:��7|p�"PV�z��q�uc��8�ث<�FN'&�suHu����;uW(v��g��bt�![B;��y5�T�;�'��i�.,+�n��n�q�z���b�z5�s��ݷ]�L뎺׶��7 -�km�VI���E�m]m�NL��c��wAÍ���a�����B�sgے�qӡ�Ms�^\M�B�u#����3�h�4��%�kd>Ʊ#puv��Q`87��:�Bg��psWY�QZ�8�,s�{q��MZکGs����p�+U���s�m��nv�cb�f�a�gS�;�ģ�r���=�ݼe�7h��O$�ll����n��;kj�t���b���ݓ���Ƹ��q�6V1g%���wF�C��P�5J�$v��yr�r��1F���[�8���ݹˆ�ú�܇����^��I"����w"q������C@#-T ? ���t E����
�9�M� ��͒T3J���+="��&��B��YF�<��>�����]*��PA{t7#�B��%���  ��B��р���s�|��t�T:��������D�:sY�SX^�y��P�ٛ.01��5Ο\j���CNג6ׅIg=e����&��m&����gמ�8˳�����ߓ�_}m�uN.ڬ!$�'!���|<{�������x��S���*���=>��3|r�?�F������O�>�����������!�X`�1������?1���N���"""%"""'�D؈����"&�D�< �B""P�"""'DDN���8""'DD興��b""pDDN����: ���tDD�������""'DDN���:p�ÇDā���""xDM����8"xxxxl�����E�@)ThN!)��P����DDD�DDD���� DDDD�DDDJ$DDN���DDDK DDDDD�$DDD�""""%�"""""����"H����b$���"&�H �DDDDJ$DDDDKDDDD�:t�ӇDD�(D��DDDDKDDDKuj#^�@((C�d�-b'�'p�N�x�g�'��(D�<"tN��$DDDJDDDD�DDD����6"""xDI�H,DI�H:""pKDDDDKDM���bQ"$""@����b$����"$����G	ӧM����8""'DD舉��$����"@����!܏R�P�J�	@;�!�83P�"�����#@��dR+@4P�R�I�9J�@�)�b4 R�H�
�j�i������R��)������o�*
(,%�����O����}�������GO�6~I�'�?i�ʪ��E���]>Sb��:Uw�^QG�"'Q:""Q�"""xD��- DDD�K.ѥ]�`Wʨ®�E�S��'�"+N�,
�B�DDD�"'�9��Vފ�Uxp�׏:L�1Xd��6���/%�i��E�}ప5�m��6'�D�%�wu]��eWbʯ��yᣫz���N�հ;x4�^Z��n�8g��͎�Z���J��ʲ��2\/V�ЁB>2r=��R�[/�h4�@m����U/�/Elc�����U�R��Npd֑^�u�M��eg��y[kj�S���v0tK1�����wZ\��rVk
�ǿu��/�0k���\��K%��f�H��k�]j���i��x)��t����s�uhڼ���$��f7I���;���qsҽ�I񇶜`�=x��u���D���Mrې����A�1�2�L=T�	2�3rcf����"-�їX���cq]b�%�����݂%��k���f��m�-SY�������mQ�u�ģ�C�����nɢ1�v܁�B��n��������B��ZQI���[��i[��H8x7I�Whŉ�.�e�6ۍ���/Y�c2lZ�[�9��"�6�#�חT��0��*��@���������v��~4�jU�\�����[�eƸ�$*�x��{8�� e*zo"�\�]6^�ކ�Xw=�&ի�^�N��٫a0+�M�q���b�du�ڗ���&�M��V��.%1ݝ5���mȆ{lg�#lcv��mwI�r�x��բ\��-<�#5�y.���w�r�e�o�y�@���\�N]
aJjk+��^<l�\�j�{�ӧse�zr��O:[���]���4�uڶ{v�1�J��k54�v�m��B�7�����c���>��틷m<N�B���y��S�)�[�Z�����vRm*v01闣/I�6c��{y�<nL~G��nx�!���Ese���f��cOGd0���7ct=:dH�\7�rc�{g��y��;�޻�3�9�b��叾G�Ŧs�*��k�p���d�=�$�sWAG�v���R������_��u�>Ç��us j�Hy��8���t[��:ݛ֋�s��1�`�]�5�39��=��k�٩��D�䛞�Sg/oKh܊�n.�E� �%�)1`�G��1�������g��BP~~""%�Y��I�"��3��3ǄDD��8'I:t�h�0�,�0�,��	ӦΘkF�Z4x��3�%x�a.��آ��A���}�������Ŝ�J��OeG�M��D�pՂ��8��JJ�ۑ�;��#<�n�Ì�Hƅcf�9�������q���S���t���-�B:
�Ab�&$��7+o7j��=<���<:Ȱ�ؚ��ONmI��Q4�<��
G�.y�.�7.���sϗ�g�A!!Yܲ�;m*I����a-W$ű�U�I
M�&B��	�{���U{�M�͢�f�B���7�l)�,�x��Af�8˦Yg��ʾ.�(���S�+=C�٤$�i㡾� �K ���wR�4վe�Z��LV�N��a�`�V JM�-#)u��B<lY|5 a��< �5dA�Ju(JC��I���[n.�\2��V�9�<5Y�e�,c��������A�0mז�������r&9՟Y�1��g
<e��i�lQh|I���q�d@�>��Z<y�b�����J4iפ����A��4[I�ч��	����`���SF�<��a�\(4�,�`龎��\D������ڤ�D��I�����N��O�E�x@�tD�����bAHk�Įج�f�F9ɾ4p�w:H�<�0��`��M�vΒ�^�(��l%�x[ZGy�|�h�@h�kZփК""'��a�nk�L
݌KH��q���.H�����M��c*�P���T�t�x1���p�h�bR�5�0¯j͒ɢ��$R���*&�Y8^X:j�nn�i�ˆ�䳆TQ�Aq�vz	V��G�E�d"bGd�QfV����q:㲂V�F�!�M�?!f�El���Q(ӑ��A�oDkZ�g<_��<6�]�����p��,�*�f"��!G�`�<{v�kA�*�0!��5X �R��٦�PBHR��
��پ�c1�#v2��D�I$�a�M�%�SE!G���Nɱa0 �F�%R!ܼߌr��:l٣����h��÷���@@�zR��u���D �0���9��DI��Q��N}�Q�-��Ob�C�H�6o�Α���7��,�P�m���V�ΏmQ���sBͺ���Fv����M�!�HY�t��yfŎM�;�D�Қ�������Q�<�N�Ud�9Kt�RY����F �Y{��~��� �ɓ�}�f]��)2ȰE�d�6�j8������h�%;��8���^ �5�(!R�@�@:LH6.6����⥹�0+M�\�J*�$Oo|[6GLF( (�4o���&�<�&���J%���92+�E�@��FDQ�.*3�\��j���Vf�P!d9h�{+���C��:�a����R6�X��=�'w���
�v���đ�l���D��x""<�1����9�}���:3ЅAb,z���_�J�Dlm��OaH��V}����0 Ά*�B1H��g����S�ޱ"����;12��RQI���8'�e���Pц�$9r���{�IF�f&�r	�u�8x��#9�LڕGExQ#�3F����
(�E�x[�đ�K�D�J""<����{Ę�p��~Yk6��a��Bd�����0�Q
�x�t�9JT1zW�fz� /�$>c��Uy_2�C���XE�s&j�N���a1ǎ�K&)��`�:IGj2wvf`�B�Ng�`�0*T�.���� �9E#Lh�h�!��A�^��xaEH�Ocb���;͜�ꈲ��DDD����Ν�ΰ�Z0sd�/X��ս��"�)Hx(�M�N&�l���wwl�b]�H�+��0�̩�8r��V_���p�1��Ns�֍$vh�#��v�;�qF�P�g�ol�0�(=s�J_�u��h� ,{[�c �\0���i�ll��H�6s�O~/��'��W����dqX����x���R���Vl6�t�bZy9�7p�99���x��d�e��e%<��sR׶�I�������{��)>�����L^i��I�˾E`�y�L��h7o:E ��J�2�Ȁ�6x�܍��d=�^��b��H��<e���	�x:���ʙ�~�	WP1����;�i7�X��X�m[�*�S"���	3ӊ4��C«�W������R��miA{V6� O�ԧ�*��j�I����H@��L1���*������C�gȚ�+�2�\�h�a�%հ���.��aB�?�I<,�5��/ՀWL/Z��+��dID�vVZaEH�Oc�;X@�Ğ��r�`� �V5�c�2�Pb�Fs��N�
��-\B�U��S�@��3Zq�~�T����\�8rʖj��X���t>Q@�	��H-kY6��������_wJ�U��N�\fG!����]�y�:[E�`��U|z����i���Pq�"�#BŉK����Uw��>���8QG�>'�<8���D�����
v�)'#�$o
�ܜ��%���nF���'D:IÄ�##.F2F2Kc(��)��#5�H�Q�`�2F8���c$b�F!�c$c$Òj��$0��7'n{Y8.�r46�=27#@�b�4t4tr�P�y��,�fK�4!90r44>������1C#�2�2K#Ⱒ܆!���M����܏	0�A�&�H�Hʒ�D��9%�C���:��2K@J4@��$44b
q!�!Ȅ4>�C��I�4rSt4y�u��zF!�G���H�I���}TH�v7#G�'}��|�Cr7#r>C��-�#�ԃFF�C:H�tA�!�Y!�Gb)p���9*I-�F���r4prc�9:�/�R��C��_�Û{���'>ٞx�eJk3ȁ���D(��Ϲf 	 ���Q#I�z������mNz�NDt�3�$R|�PTȡև/P�
k�$�޳#-N�Ø:��M����*�R<o���Hv�՛��%���|w�tW�p��F3ቄ��eQ�I��sZ<a�x�0�,��0�(� 4c(c81���c<x�Ӈ1�i�����3���w�4��{�t�4T�9�^gGq3��I!����zvW�����a�bM
k���F��q'�C�8��E��C���\a(8�S�OH6�#�CM%G0d�d�R�fEp�h��^#�����ˎM�b��d̦�~`c sçIuΔ�:$�5/��h���%
���)ZK0��,X[1��󁫞i���(�y���7��s��L��x��cĆ�୚�p���4�^M�h� �5�O' m��N��j�	>un�f�w'��(: �0� aJ5T�`�a�ڎ�o��w�dMH�o��ε��s�,:pu(d!٧� n��Aݐ �n��Q��ʚ���Ixxj3��{��O����H@D!�����!��t=6��ZsC���n!�e}D��d��)�8��pOLD'�;�ӆG�\�&�D�a"�bQN���a!FʨB�5��8��� ��u�a�N	ש��7�`Gf��>����V�p��p�3�����Al���/f�fWD���8Cr-A�b���釓1����l�Jj�|y+a�-��*�a�q��:�k�s���`6C�ɉ�)�d0�ġ|��í��z�}��p�#L�?=�W �$�:�`8A�Ʀ.5��l�|/�QF*9w�{��v�`,��ع���
�`��~5,.�n��!���,�k�)'�\j���2v&�r	w�I���q9ׯ#��Xr�)��Υ�l��<��z�u@GN�64��ܰW��8�8��$ƹv%Ɩ�S��ϏD�8Q4E@����/�|�[L܏�Zf|K��X�c�����L,�My�hL(����6��Cw�7�[�������;G��M���ts���!�'���;�7ދ3O1�I�5�h&��"L���tnrB�d��i��N~[ֳZ8_ߘ.�W��{���#�'��l��
"|�ԯ���"�P����!�����y'�Bw�̈́���w�����9�,�YW m�d'D��v�8:�9��I�{�'3�d�A����|R샫�a�����᢫!p]aα��Eф�����t���p�Dp@bj$6m)�7���~�d(:8Ɂצ'�d�1>�}�4:��X�|QE�\�ƞ�Op���!Ned�@�D�=��W$<$��2Ozm����ݞs��-�M�Bq�ܞ�sGXLL:��U����J�ɒm�D�e٬]O||�ְѣ�}#�@��V��$���/F�ve�����܏���G����rx����28����I��1�	�>eP�L�TLm��e&��8�Wk�e�[_Qb^ /��3T,�2���ch)/}��%���w�-fzl:��;��a�#��Y�o��d�x��ј�eb�˂�Ǭ��ދD�$���9�h�%�Ͼ�,���.m<-���c��{Ѿ:�{��O�"������Bh�{���NI����-#�+G�������\h�<;a�^��7;H�{�\��L�=G�����bD:aÈ@q{�q��W޵�	���Q�T`��3�T�TEh~�ML��%9kk�w��3Q��Q��Ҝ�vAŸ<�a� o��|Y8�b��:".��8�ffVp��"4�۬]B<s��;#�A��-#�8m�N7�'Lro�:dx�����%>F�]K�����b��b;6bq��G���|���_�ޟ��gN�>�.m<-���f�����/��w�����A2Z�'���|`Z����8N	�|e{�d�F�v�lşz����=|��֭NZ{%�"NNw���{�~���s���9O%d�`8��oHx˨��Jq��02��00����p��#���9eN��k��~py�;�H�Ą0�Z�,�N�W��̛�4�.7g\n�v4�/}�`a<�11����s=��L�돗��kV�NX5�3��M�ĉ}1ρ�F�^�آYD�� w����@�
z��J#�@1�V�c-��Du�aV�Ye�\�x[/����+�.{lx4���H+.�H�D�a@��N��~N�_���:����{�Č��҃�+�ӎ%��LW���cM����z�ٱL�R�	D����+�4Ӈ��;�s*��D@�(D[�����o�j�Ē��[L��0�rEDE� �v��]�۽;܌�x{=k>������^Oz��_n�=m��}:t����6k�^8��4����]>۝u֓ۼ�Ӄ�>@�:.�c��|x�(��\Ӂ�0��{/�ǗFivF�_N�5���q�����7n%{���( p�И�E"������̸��G�<�#f9�W�o�5����I�w!L��B�N�_9�x)�O8R<S����kX`T\h(�wT���;�������qm�&��sp��\0��U�@�Q�Ox�-�	Ib:�ԅ�QM�־>,�ϳ�i�l��Ӹ:B�3,��NF��h����l��㲱�˘6�&�V`
�^Ƽ֪�8.�W	|닾D�c�N�wᖵ����N�VI%ۢ��A���vlwj���(�i�4;#��g��3����y���U��k�"�H)���IC�t�8��	�Z�6a��Y�b(��{��y��C��~�fj�h@M���:<E��Ʌ4��|��#�Ƀ��*1 Әt������8e'�.8����C�^H�<�E�>F�2�w���
����DIt7ʆ2�YD
f�]����>,�ϳ0�Nx[���f�����ߠd>���"�e#W&f*@���p�� �up�d]m��	��[��wpOHzF2�8>���<����vO�M���L/<�GXG'��t{�W�"H��x�#���)�3@Q)���P�P�q�/L�L�8h��x؝N��s�8��`��::g�E�5G|A���?t�̾0�X�����瓇�L����U��Q�C��ZOq��~ٲMj0�=�-�tI�/�'d��JL��|�.9&g\�t��Jl���/S�O���߽x|t�Ѷ���g���wN��
r��(��wf��D3+�d=pUٙ5Y�,!×5,�l�z��Zd�z��ܞA��`���φk1�L�2�gy�t�G�o�)n��ǎ6kO1C��-p�^��zI��~�����᎙藸�qŚ8_�&�`} ә��2q|��X��D���g��m��Ѿ�!����i�K�3Q�
�2`���VY�#���P�sT��BgI��D�Q����a0s!2������`a^���f��G	��nO�rx��� >~w�΋�я�y�19Ml��n�I�F|I��GF��c���hnF�nN�~${%!���t<,x�h�客܇dt7#����t�'Np� �1�2�C##6N���H͑��$��`��,c(�H�H�d��<2F2F"��1�u�o��������#CC���#�`��i�O�Q�< ������"%�&H���&���C�N��:98�C#�H�Hq�����1�2仓Lt7#��nF䑺�a��=(��1*JEp��9$���X��c$b-(��4	5�h�$��D9;D�zMCC��#A�I�K�C$~$�C1�1�3�xG���H�,���?p�}'�I��}D�L�d�h���NL�!�dh: � 4qGPqF*X���4!�R]!���#^P��]d��S�C$�;[��J~��UNZ��/�ܼ�Ƽvu��I�C�sCi�R�0 r)X�P�#Yy���f�3^����n��l�&�cF�-!.�K	jgn�T�E�s^;Z��Մ�1$wq�����a`o3���cl��3�-���|�K����<�e�r0Z�,��r�)���E��ޙd��塑5�.�J�IHf#�q�6Z��ʳwp��v�� A,/z1�
����ߓ�6�,!,jҿtv�Ńm�mn���cP��Aw�T�ŧ�	HG��Z�Q,�Ǉz�=m��$�r�3%�K�����Y�KzIp�Y�=X�^���ucGR$ 9 ��2�Xm}��!����;�w�6�ﾔw�[S y�0�T��"Bj���Q�`l�z�]o�ī���_;���8�q���r�iݖP��B�@���v��bd�c2����=��-���SL�Y�Ĩc@��7�'f�L��uw�7���GՉ�e�dH��J�1nō��,\�N�Vձ�+�Ŭƪf�f���ja�9�$�8�3����C�ɻeQ�7�n7=�V���T9���@�m>��a3��8�xM�	QUUW}�8x��|3�O�1�gN�8xc4�K0F�c��1�c���4�4c��0؉�`��Q�<x�׳(�KK,�30oV2_�雂'�;ÿ�[a�i�&�3��X�j�m��0'L] �N6&u�g<���9�vzX���:�Buc�v9�-�fŖTe�Q^B���kR��'#��dv*D���W3���Ҧ����oe��9�aȓ-϶�*t�ü��'RL��P.��5�=���G�9k�G���W9\��m��נH�ó�ug�c^��o��N<Ck��W��;��Ut��e�K�٧+E%�K|�,y��mE�1�ov�r_��&A�n�<,�J_i��㓲9�b2ofRA�0���GD�Ɵ�����v�@tG��d<;��7�P�G�k���>;0�@q�0���pC0|G���,9<�<�",�"0�H��CQ����IZ��[�H8������980��f������8�Z�gD�Ɇ��X��0�&���e�ˎ�y!�y9�޳��ټ!�1�E:q����A{�>�<1�.��{G.��O��q����=�� 3˼�j.G8��^/,����33���l��f���̳8�tD�&��B"(!�e{ۆ�:�wavǾq:g�YѬ5=���G���1�v`�[.I6T(�T�$@�T�2���;ӐR	��:l𳉭�Gd=�V����X2l�{�l;��O������&.��t|p��^����H���}�{���h�	evV̮x�mR��2���E��#�A��C�G����pHټ-o͝O+��gF�������R# �$<!Ժ��x!�Ϻ�~f\p|������2C�]%?5�'��z6Yff`�x[W��f���������"�gұC����M��W��	|gLh��{�pV�{>�Y���|��᳾����ru3
D�EF���<"
����.��y����u���6F>g������]�����,׬�p���HP��{\8�l��
ɒ;�JB��EI
8b�
�r��(d��B��H�*��XigX4Όm��	�4i����;d��<<����o_i�vO���x���<����ff��l]_�雂'��þ��y���AD�>ɓ1߹�sW�'��=A3�^��M��pH#�Ǔ��$�\m�Lk�K),�L�(z�m�~_}���@U����Î��4Xܜ��me�ߛOzq����'`�!6a��Mfg;�VY��������c,Ύ�V��0��`�z$Sβ�g{��A�@L��.3����u���q�z�莏�m!�l�&R *5�Ovu����D��v��4�(�
(l���.����������=��T�%͗-�"Z�m���N�1�7BH�u��:����GPU5�tvl��l읙��k,U�V&��qj��.c\NA7��"�~��KX���ܘ��J�ZKv����EH�W�C�
n��,�\=ט� ���Y�r�۩h"��>Dz��Hz�3i�9|p�x�����>x��=�����f&����&@����"Vt@�8Is@Ȝ��Qu�x~������ԁ4h� �R,��Ӫ��e�0Z�iQ�4:ݻe&Ɲ�*�4k����� �5�2<�_�.��ͪjV���q����]���$> �Tk����9~���ſ��ȃ�j�����(s3��e���_L�Y����F����%���}���J4k���r	��-���F�J���}�綥UѬ�A�m�^��x�Ϣ��;6�e|Ŏ�:I���6ٯ~U4q�F�����d�ÈB�%0$��*F���]7�[�N���P��~d�������
��{,L�NIN�vm��gl�>�ث�O�8y��y�7��;�pt���3�kE6P!%��<,�u�G%;�<�gç�L�V����2�?�P��F�~�V��%���\h��i3�;Ï��ǘ�3:ϋ����˒�r�I Y�����7s�ԇ�����K�khP����a�h��痓�OO����t볷������16���ò�x�۟Y�����s|=�����&�;�����β��6١��D�EDH�g
珼ώ�8w���3F�?Gt��I̓2�=jd�	i�K3˜��p��wL��a��aɅ
-�>x
?��L�7Uj��o-�&�D�fʤ��J��a��#{6��.�f}g�<Ît`a�w��<&?/�7���>_9fw�2x���q�h1���fG÷��Öz��3����;��o����3�7=�g�ߦIȒ�^�>��B*�Q��΢�ŔQ�f�Y�c��}3s$��u������,�[�u4u�F(�v�E���t��`ݥG����+;\������ŃmPٵ���wWH��,DlS6f�[u�Ň��Q�I_������R�����#���7�mu)�!�9���r4���mz����������ݻ�&���}�f�]����C� �@�\�F�J��;լ�F|:>x���(�\��ٌ��^jI:��J���WGF�[��c�@���Q�I��4`8A�tm�:�0�'�0.J='Lܠ��9+~�N���ݞf�Bh��|DČ� �\'�����������AU�
�LtHT?m*;@���{7��gլ��e���,��������u��A]�oЗ��՚�T�rK5�N{���Ͻ$�u�i׽���"U����T���H|�! Eo�$�����WS��;�Ń��,v�����G,��3|�������Ϗ��c��^T�ѣ��м�w��-n�5J[�"E�5��7����hje_�h��0uo������PS	b3B@�|G���Y�V�׬�w���8p�:lI��A�o	9H܎]�܍�y�3ãU'nN9������̏�H�������t��:p��	���1�d��N1�12F3�1�2�!��X�82�f��D1�3���1d���b#����I�w$m>�Cr4=���h�!����1 �|�vC�D��	H�.F�$�r>��P?4q��2F!���t2I�!���h����t:�����C��4�L0��$�����R)�#B�I�(��H�e�A�T.F�NF�CE�!�CC�F���0G�nF�G�4y��P�!C�$�����8vO�H�v000?I�}��L�3$̓,j��P|���|��L>��p�N�>����5�1q�R1d�B��,r4X�����'����<͢rF�!�T4)8.+K�EG��P7�l�7Â�j��%!����>o=~~"qܞ�c�5�B�ή[F�}��3璿Y�5�9��8?R()�H
(��{
��qQd����$� a�/#k���`�tWy}��G��	g�>8Q���DO�Θa�Ǐ0�8""lDD��<t���M3FpcC�x���f��<x�Ӛ�l�2�K:po͏�}��wS$�I��B�h��:��{3{�M��>{��1[��TYΑ;����IK�G¤��ʃ�E!P����F����Nc��R�>�mѱ��FI����-������4����p�;GZ��⋐yc���ɶ-pJД*��z:��M��Su,�fG}^����>��	F�OE+EJ���tߐ`_�}��˕%��)WJ��������"ˏna�:t�ߛ��?�p��I̓9�LAJ �9�!��q���Xl�	�첒�x�{ن#������嫕i#��I��Yo�Ao��Q�5�Ii3����f$����q{l��ü���ZB~��HH�X "Xd���V;���a�?���ct��B��p������$,�9�����p8OO�t��Qo
yv|H�~����4D�6Q��,�1L��O����y����'���&�����ݸ�;����6ڌ�!�VcP'pZ���
yY�j4썷X̩�a.����N�'Rr��f֦ٲ��k3+�k��"�T)�a��k%�#n�'�FDZj�<�}���DY����}ً�밈�cd$
W��.���&! ��&��L����F�!p����$�8�R�>=e�����C�+��{�udKB���'��BA���=`J�U���D�ÿ8<��Xtk9��P�=';w_j�	��6h�9�9�4Ɵug���@TaF�		0�`��4�j��¡�Fm�E%Je)Q�������C��Yff#����x_GY�oxo��fbh�Dǁ��:ZqC٘�<\"��;��f�yQ0�4���;p߆e��c�Ϝ�^�q��E�p}���x���^*�D�48�U��=��G����j#-�V1%x��)���#��Q�D��wԭI���(�#=G8�J�G��(���\�w�&�����ӣm��c~<7��z�I̓7���M]#��D(F��S1ぱ`�VI
��>�'U��Z_��Ԥ�/>�)rUU>,k��G�#���(��iBG���Y&��f��mn��h��¦�w6��/�8|
<h�G ��V��>�D�;�f#�>;K$��CK0�_#E���D�}-�Gz�$p�%TE����#��%��%
����"Cy�O�Ӄ�,�30o0�L�4�x;�'���kE���rCDt�q����!�z�e��`�,�mn�I+�$}�%w��V���l�%�%&<o����=���Ņ�/P�����6Y忿�Q�7��!���\ξ=ꤷ#����)�u9d��8æu.F�����0���[t����S����\x��P$_O��f͡$�8z*uETB}�����\�t�mLL>�K,��L�L�4�x^�I�d�>m�E$�%��+&r��.ڴHD��;��`}�q����q�l�JY����v���7�����քN&t\�X��c{%S����'����|����5���}�c���IM�2��JD��2�o=��=��q�w��u�q*�������t�N=�p�*&	�I=�u W̮Y�	���Pb��DO��e����R��N�h�h�}���+�a(��膉ԑ���Q��G�^���g6SSf���IiB�0~���-�@�3�·{�r1�?�^X���M��fbY�����{�G�/��Ag����� ��atP��Y��e����k�ziv����T�iA�@!����F\�-�Z$i�NI�a�T:��=������x��i�+F��g�?G�5Ī�*���$�iT-�d;��A^7̖@��Aa`U����c���}��ɶ[i/��M	��U(C,��u>�t�ʝ4�(^Pن��B8J�F��agQ�>�/E�T��GŘ|Ϳ����H�ؼ��0Ĳ��pQl��5�܄�aޟx�Eǀ�"qI���,��&�~����d���4th$*���(q|Kz:#��N��0�v����%g��=��bU�#��hB6��D�� �n&�I���]�b�L
�;U��`�F�n�����>�nRB��ǌxD�G����D���ilƖ��`�p���"�F�ME��
��JU�����āoD[���:a�����tq��~��~c��tm��jd��3�J�r�:�!�f���,3�ebVY�Q���,󁾍8�����'/�Ѽ��6�XFI���<�#��F�~����1TȔ���}^{N�x\���%��8����ď�**��pԕ@��E�Y�Z.*����Q��\8m\���cG�2������IHF>�\���ݥB�;��YFQ�Q_a��<Y^;�(�<+"�׍->_�;���^е�=�U�QQG��b'Q8"Z@��H�"""JP�"m�O%���7u�]�$*�Ү��P�u=	�:yU|u[�8��B")"Jor��UVEzt�Ã�D��P�`]�H�	bq�sF��n��췅mh^7�N�ä�""'�����w�fHfb�BȬ�f��Q�gl�>�{�����k�ؼ엷ǐ:��c�Z�w"���bD�u��k�໅����[(��wՙ���+~i�}M�����&�_g%�Y��n��RF�Wc&f]�fa��H��r�7���J����g�m��Y$�]�di&6�I�%#p�7�Koĕ��	�g-e�u���d^�AH�w�j�$g+�F5��JP ��=c2��d�����ːHH�:$�^yD�02�RIS)��
���f�E�ʢS�n@���-�-���E�x�`G�"������G`�i[� ^K�b���l����4���-S�ƥE�r$R�Z�-��<������k>r�'V�D����e���G$5�E��嶙k <�i,�f��l�'X�"�1+ˀ�J;.Xa����<�g�s��'��i��v�ՠ�n�[�����g[m�`�<���4[r��s��s���hv;P�X����G��v'q2ݝe�J&����/�ם~k��m�x�.}y]�l�Δ�����B�O��Q��X���fx���0������fx���0������0D����x{'(�,�,��E�3���A� �м8�x�$r6��8�ջfj۹�Im^DX�c��z�꽙-��&r2��Q�=.L��7<c�n;�bsk�>"q�x��n�S�c�^��3��)ۥ����zy���aE�-�u�Z����V%0]<͒�6��S'nԺ��J,�f��6��٦�L���Hє�L̛a�(�V�zm��7�v+�<�iF�R7X��9��D⅟{��'����o'�E�!�ɝ�O.Q��&�\Ul��+2I�����L����-�[����w�\��m�	z���F�e�BD�o�=�u|ꉴMsx�CA ����Ă�hB2���ƝM)kDi[e"Qn;�Zc�Q�W�Q���z�i������z�q!^rR$H���>��IC���*��"x��۷�Ƨ^ٞ��aE�BO	>\��t���>b���4JP0҇0<�g\=!���J�*�G�C)�0l��xK31�0[�ΏN�d��N���Ƶ�^e9��D�ێ��=#Q¢َIy|3Ƞ�#�ҡTp�;gاb||.��%_��$v9��R8��Y�ヮ�k���pfWJ�h���46��pQU���4LB�]�̌���M|��$�"�^H���r�D�Pr�@��B0����UЀ�%-^��L��n����p�^x�����6?t����*d��1���F!���4�5t"��U2J�M�F�;B(�s0vZ/�5��H�<�5ƞ����iB H��#�\	�mqmWB���B��<?_�'�
f�s�,5&'�K�0��(�w�w�t��}f����35TQ�$�aFl4zXg��h����SPA�d�x�%3��%��"@�(�O��X�e�%���a��fgG�w2Ow��z�g�iT�D3�:�!�v=����t(���R"�~ �y�����1Ro�I/�u5. \h�$ ������%m��F=]�M%-(�����>��$!G�0Xdf�}&[��d����z�^�B�9	��1�9."��T�YS@��!_�:D�zV�"��iIN��,����^�c��s���4=|<����̣��%���a��fgG�w2N���'nܿzf�Ҵ�	Z�:���v|�{;F��l�Y�J'z��6s�붏�s7�H�%�3�y�.�$��a2��1�J�Dz)�R�����ߦC���v�Ƙ"�����, |O��w,�dP�1�_'���L�6±��0ÎH�Q���1dk����0Q�z�^����Y4_{�L%�8�ԧM��:ң iH��,��$=�]�l�QhE]�{U������͉Bw�a��+�J#G���&!���X�`���\�A��R����h%g��RGHMq�;�c���l�<�H���I����fh�hn=��h��G�Q2Y	�Z��2�K3�<���vy�z�3{�{x����y�.B �h�à�㏇'ǃ"I���|�,"�����z���0�4�FtU�#��$�|�	�Z;B��j�$�h�"l7�_N���'H���r��*�.C��s>s�+��D�5Sp�8�6{`�%&|Eن�IB�8�hɊ$u_I(E�Y$��L�=�p;�����,����0̱F��*d��3��	�W��H�B����&xlҮ(��#�ԑ?s�~�C�"};�ӄ1��c;KX�!Y�tH��,���4h�5p��������o-�K���t�Yj3퍳��)r;ՇLu2����#���_�{L �i0\����0e�&�8,)bW%�|r����8w��J�L��J8�%<I�`�ei$ٳ�N)�(��,�\3�}=᷇�ʙ'2L�	,�����%Hσ��HB���G�i����Z��y�k�{�����#��|a���h�C�+V����NA��`��G�R�y�%L���t�6��+��L��ɯk����QQ�_������N!�"�����(�qd̔"�Q���Ѕ�!|r�i&a�2gׂaEن&.���ftl[H+�.�ˁH�re�@�]��{���5�P�Y$��a$�Eӷ��2dk9]�zi���N�~�z�����Ik�n�]p�t�[��\t��r�����߇�D8�Ϗ}�ݴ��r<��4�#��b��}����EK	�cc.xt�ް�}�Y���}i����р��,	�Q�0t�eL���\h>�1�$X�K�4L"P�{��Ԩ�6OH(D�d����7�#-dd�]��A�H$]P8��v��M�2b}L�çF"ѱ��"D�WP�1)��.��A֣�B�\xyG�}e����G��(��>��������(�OT�W�9������L�S3:=;��{�;'cF� ��N��E� Q�qST4���TQ�z>e��R[�/�B=��C�0��r+�J�`�I7K�`E��OBix�j.$�(ۙ(�	e��?%Sb�4Q#D�.(���"��9��H�h��nf�����IV%�Eu+7�fU�a�|��i1�Т�}QE�|uDѤ���1��><s�}���#Wuw�D�Q��I*�4� �t��^		f��W���V�M�i����m�
���(�[,�e�"'�b":DDKHh�"'�D�%��ѻڪ�k�J���P�u=�:X���z�$�":DK"$��*��Wg��:p��&eөXd�"$Мg	�ͺ��2v[¶����I��'�U��K��p�f*���,�by2��Þ�o"�����V�Ž�㮟Oo۳�_'��y�rx$#qK%��M[�;���d���0�9=�
K!����C�y��G�S�kuW$2!���,�D6�ѡ1��D��n�-VY#Wr9D������Ic!�J�	���$����N�,@��Ǎ��"Yg�$�'�<a�a"""'DD��$�<x��x�0�L0�D��e�`�ag�6{3yEQ�a�b�ߏxm��2�I̓?�I��D$Y㤘���LN3F�J�I��V�,�������F#���4��~#�zq�Q�ǋ��L�2|���U!e)(����l�����bC�}�͝���h�x�`�ivH��o=h��%�4�.H�� �&d��1�S���v�#���$��<�C�Q����<Ty�	$\/�_x�3\2��S3:=;��{�;QB�*{;�� �Ԛ�PD&HjEԺ�.N� �h��prt`%$h�x4|25K��X ��T0!�~�!~'���l��L�bP�g���Ǎ�v�� �À����$w��]�=T��j������I��0χFH�0~�sr���%>�Xz0g!H�	�� ֑ߪ�Vҳ��A�IL=}�#�c�RM.#�(����#ĢO��e��:���|1�P�b�f"�����̓����O;li8��BG G�k�+J���sy2/�=ni�������#JܮԺ��"\�l�y�q�"�S�^�a�Y������Z��vRF���O��S�N�n��+�������30��Ld��a����� a��Ǧ����a�����US3|ztwOϚd9>9�f��R�`s��V��4ϕI>tz:b����oя�4鸄��t�D�Q�V�BF�$w�)P'�c�� �!yS_T����Q<I��*M%��v7?uIOO6/*�a,��pxJ=�d�l�L�ޝ`p�{I�o�,��>p��3x{��s$΄��p����B"+������QH��>#NȮmL�-J:����Q�$���%�P�ІLb�
T�����qE��J�~��I(B*W
�X�\I�gm
�Ј�iW�	��;�A!���S10�6���BVin�d��t�X���?h�]����?0`����ʁ�I��G �j&4�-0�&<D�"���+G�i��*z�ifw��t����|1��}g�6��3$�e=s"�,�A�H�M𦪋��W�3O-�"����R{��=�
��A�CK)�M�.�9��	v�5*��3���w�D�Z��-U����In+Uwk�G�G������m�B�Z��̫
����֑�S�&u`rl��o�j�p�,����W1��Ƥ�;�@ˎG���we$)�#��ZQ���7���&����3�{���Ѷ?�i�L�9�G":�Hhr�tCF�����)���}f#� �@�p]A��=��2|�E���˒[���?'>I<�x:���Ta�@]���P�F�+�>����y��	>��ך[�~ �Q�
�\2J�*�.!�/ y	�R�a|秅'7z��*�#HH7�,�ML"�_�p�_���H�k��<_h8!�`����9϶�EQ��e��bfc�d��{O��=�V5~�m�kd�_���l�{fѨ����m�iHM�R�Rò�b��;�ӽyz�\�����S�W�vn�6�����D8�w�o��������"��S!ْ;��GQ�e�!�ՒA����M�/LO�{f�ӕl���V��9�T�v}ѓ��	�H��.�2M�%
,E��Da�
Ԫ�yZ����!#�}�l|�u�3\��`��<��v!(�'U��(�oD$p���`@|/���'����&ѷ��X��Q��$�]h.�C(��ta���BW߄�7�%P�8.ff����ə'�ގ@��h�"�����mC����j`�;2�9��{*���8�P��ǿ�����|5��:Jυ�u�ʒK��U���c��Q�}�2�է��,��5�՞K!L�hh���	�K����쳗i,�-��tR����'����þ����R�XQ��c��/)��.\rbW�>+�G�ȵz1�G7����]m����F�p������>�:�y��ll�~���s2�*�,�
!*�Zt�K����T"��#)7�ߟ
��gN��N��z.���4u����h��v<	�~ͣGǎ=�4�a&��<F����������:\�I�j��k�����ਡfC�P����c�ç�/Vf�Ye(p�V���\'�S귰|1X�[�����ct���W]'症Fp���;��1�m��o�as2NfQ�8�S�b%+%JJ��"q���Fs��P�{�qѾ�xt�̥�&�����S�|����?�ޚ�/S��bH5u�@��:/G�I�o{J�7>��Vd"�ѓ�~���@��ω�d{2H��Y��1�|�$���o!M���w�No��f�^1�qú�7�E�q��վIn~ f��k���*��Y����e��s�{[���,�ôa���Jг�^+B��Ȼد�R�6�
�G�QCe�W�M����"":DDKH8��"tDD�#˾�>����da`W��Z+J�S��ӥdU<+|D�6���e�o{u�UU�=:t���"L˧J�����=�Ǆ\8뗬�36fWIVůqӤ���DD�M���̼�Ff*��
Ȯ�>�ٙO��+���3X�����{�����Ɡ�0�z(�-#��d�6���>>���m������;.����&�@i�FVG
Wb���*ya�l�,�Fj�p�C���a�+6X2$z��4����!���<�ĩv�VW���^�4NХ�es'dy�cK�t]�1�b**u��Ǽl�l����
w'S�Ǟ��o��1�	�X�f�e��À�0,0�h@P�o�㱘!�\�.b�F�B�8]+��B)��8�y-+�%CQ��<j�V]9m���+x�t��v=ի�u�Z�\L/�|��eۣ�;��~E5T���.���e��af�|�D����`Ȭ������v��wǒ�$�ys\yCV��CHp�vm����"
�n9��]-�֞�����sj�Xk����$��&x�T�	���^�Fnp��[2Vl��{�>z�Z8=��g<�Y��	�:�"b��vrݼ/M�S�"��a�7f#q�{��7�x��$��DD��e�|QӧL00�4��N��0�1���1�g�O�Yft��ffg(��(�:�y��ll�~���s2��,ĮWM덛@N:}��F�,Iђݽ��ye\#�IťɥRח�%�Mʦ!K\<K�z67�6���˞vUC��w=l'@K �N��5�֚v�G��A��d�rH�V
�ƷV�h�n��A7&ɸ+؎�a2X��е��*l�2�u��:{na	:8)@�G;�=ms��C��.�n�v5�7+b;�n�Dx=�����Ե�?E������x��v=��DNm�,�*g.�i;I�K�_���..��W��ݰ���(�&�����_
�R"G ��L.:�&8�T���4���V3GR(]�B趏��JY���L/f�zln�R�lH�^�R��t>.����'�A��S�^*��߇�n��~�q{���>t�'�d��\����m�c�Fn�i��G�80Ԡ�*�F��cL�}:�Cs�l�����ŔQ��x+F�����3$�e!9�W2��BNraA\��8u���h9����,���\;�8}�<W���Vw�UC�VL�O�T�`#S�G!���퓂vL%���"���߅g������gt9?ud)�K��c8�bjz{�����(��w��#�"�܉���ܐ��\-��E�T澞���O�>�pi��O<a�}�^�Y��`�>:rfI�e�!<,@�P,���JQ�Iw���]o{ú>�x��zO3ZG;][��xKөg>GǦ,��1�Ю5{x�B��c*%��uK�s7VQ)�N&CH�lY�FV� l�>��f�BF��Qm)�L,��*-����tʊ}�Ġ�}���PH!y�T�a��\/E���� q�95S����|�2
:{e���,������,����|t�Bw��u���=�o �#�"�~\�W!�%%�J���nڒ&�E�RcgY!��p$�D�Q�þ
���,EK����b,����k�\�:�3�M�H3�m��?�F�~#t�WG�*�NA�IXr=���d������Ǖ�j�Q$��?~l,L�(:>�h�O����,�{�g�p����c��<���$ݱy�����8�Ẹ́E�����Ť����%%����g;`�[=;
�"�'�k�I|�VX�s�`+#rK(�y53m͔��t�� ���u�9��!�H��x1���fk�����@4nXI;��A!-�f�x��0v�����|=_i��.'�;P��致���Q������&3�O�.p�U�,��|b8����t�3���4�R�A�E
g�Y�XY��i�ͭ���V!�����ۣ�r.��W��|8,0'Dt��-ē� �E�a���h�o]�i5��K�y��B�	�}����B�)J6/7zv�(�%�8Y���V>:rfI�{������̔5�ֶl� �.���� h�O޻e$JB��c�M��*^��[.�=�O��z&�Q���8Y��RqV#��Q吶�R�k?�ہ�gX���/7�_;��Y�=e��Y4�С���㤼��Tp�0�N �K��IF�3�/�Q�Ƃ�O���t�{JA���'�|{��oS�%}�K�~,���+4���i?=(������X�����#ݟ�D��OVU�����~�G�!��E�U���S1z۰=G�;�!���!�:�Z=D6U&��\�Pҍ0�J���!88p�+D���*������dL��^qA��>u���e^�UV�©���i	B�8!u�3Ҳ�~ԈCDkկ��U�ݣt������E�.���3�|t�̓��e�~@P$�DG�瀞UN}W�}�R��C��=I���W��jBIA���a~I+����^�#���;8��uڧ�TǾ�����bwE14-TIދ�*̊ذ¢�Q?OJG��6ay�Ը�P�R�I��&�9�FEV���x�gc�+��e�F±�I���P���z�P"���F�Q�g� X2_����|�.����2��ӓ2O{'w3��	L��mD�a�m�����w`�k!�m�ݬ^,c9w��IS���a%����5-�ۯ{'^�8��lm��3d1G�*���|���� ���䔬�Ņ��x�����Dx�p;����H3��,�"��7/���r��{5�P:H��z�6���()���V�3��9�"����H�
p��Q(�t����9��_
l���}��Q3FI 2����w�(�\��ÄD�ؙ�+[LN�h���z&Bå�������$)�L�!	-��B�Ňf4�%#���Ӏ��r&73�G���Ec�F�3�=x{��s$�8�0�B,5:鈒f{�,�ٰ��Bʆ�&��6���_v���!�$�@'G���i��<��TR?
����|���]]f��0L-�|S����p̉ײ,�´Z[A�l�r}u�w��+�ͮ����Ϗ�X�h��E�G!XE�LPs���,��I^�q�v(,��a�����N
�YVەhT�4��_VS��"�E<x��R&͈����DD�DDD���"'舖�l]ؗ
��,�.���Z�r:t�*�k�DM����HD�˥UZYU���ӧH�=7�N��;6H���N3wz����f��t��ŭ�Ӥ؈���DٗT���̬��f*����_hn�Y�{n��A�́��z-%�[�z�#�1.�3�[��ha��@��	���;���D���b��6�B��S��Oe��K��eI�0�^[���l^nj�7����@���""'�K,�
:t�af""""P�Yf:t�a�����%�Y����:wQ�32�=Efu.ѣ�3���ͤ��M� ���);��k���\6쳞��yA����<|v���qBKbt��~��?��(O�Nj��r�`4�(�O�V��ZW�r�_�ˎ<��W��u37��,�E��OO}aؙ	�ظ�4:�숨���Q:>�?z~?��]J&�U��~��>=EcԻF�30p�gG�72O{'\�1�Iыg'DD�"����1\��(�ouE�����>,��~S����pF�R��8bD`����K���]c�3,�����N�j(�7��Ό����0 ���`�C��&T՘���Th�z����Đ?V��fR���!7X���&~�³��:g�$�c��#�e���V���Th�[N�uzJ����QE=K�h����=���N�'�^F����U�o=R����/�˗\�ێ�-�<��`.x��zۈ���z8�lv-g��I��Y/��"#�׭��|�����=���!صc���؟�r�e��ñ�q�.n��<-1AqG�K�d��Gn�A)k�WEUF�£G��T�(���G �n[KW��g%)s�lp��G��
&ji�>�	2Az�V毶�ϴdx�%��F��R�����1�bD����\'ѫ��Gs�w��;�-Y��=�+>-[&���잣����QE�.ѣ�3�tzss$���Th=�^`d/�S�8a��]��~��)��I#cH��B]��ա�0�
�F�P'�'�顇Nǡc�͎���s����W���ϙ
П'��U�Ё�@��3�F��*�)D�*"�Q'	
��+�)r�5����QA��G���)8s��x}6>ݷ3|ȿ��Dk�>�9�D�P�N�Ǹ{��x��S$�\e�B���	F�f�}ZA���!m_
�ʴ�A�ؘDs���7�$}X�c4A�E��O�}�?A�j��Ј�W6d8f`-9=���"������W~W�F�D��������{�UM%ϸ��Rn���~�eӤ����F�b>h���$Я��&�a�j��|I�_���o[�"<M��z�(^�ߏp�<Ǐau2Nd���!B��$�y���膏�%�K�x��e
��n�^g<L�e%���5�B�u�_W���kl������w1�`�׸룇6�KM-#)�L�)i�%����q٫͏t޳����'E���\��~<ß����3���*���A�V�u.�&}��w�#Y��kq<&�݌�>lJ*��v��`���c�#H+��>B&ɉ���4Tl��T��PE8�WX�wn���G+��w[���O�ԓ�g�q��;̐��1��Y�ic0�A/�""<NwFPVK�}��R%h&����Mq�������h7`�HE*fK�}47���jxs�v�Fe��8/�B{��f'�g�q�#�#H����%��pӜ똟C��%>ܪ,"�3���b�c4�����9���F\��}\�Q�U������q2ex����_ST�w��;�}_Q�i���C$���5��-"���f�͙�8�+�Q`5'�9��S'��w��TJ*��v���y����d��5s4Nݗ�B7.<��t���]�£��g�H�~w�w�6�2�'u�V�gz����E|����A�/í?;�A:mO$���(�g���#���l)�yJP$D�&HE�.W�/�v��9^usY��^��X�Ľ���=��WS��
��R� ��՛��DnqzaF˽�}�z7%t�ا�E�.ѣ���1���]L���"Q�1A
�� т��lh��ǁ�w�DU/Vz��|�"�ͅXx�y��f����E�d��0��l)W���Q�Pi�L&F�a"�(�Ҋ6����&�m>G� �%��#Oj��%���ZPϣ�0�v���镚� ���!Ȼ)՞�+�(�K��h�����*��<W���FU|�.ѡR��2z=6�
�ȍ�0ٗz0A=Y���R�����=şO�_L3a����d�MC� �D$�Ck��׎�S�_G�IJTi���3�.�7�M�K�37�����#6M_0@��*�b���d����x��~�d�[�{ơ�pme}��EP�0��k�&  ��u��	%�YG��ŉ�
�Wb�U�V��KllW´���;j�<x��KHč"""J"""P��DN���%�*7~t��P��͋�hZ(V�Ԙt�����U�"&���l���7��U��U���:lD�M�ޝ+��$DD�#�a�i��p��ffa�>�:M���O"&̻�n��fd�3i�
�^�|X�>������ȃ5�f���z��K�]�����)ی�s-]��p!g���A_IcM��"[��i���`�q�v��ǿ/gmE�a�]���m�q:��{,�03��c�scs����>P0pቲg;�M�Mm@��w�1��7/�F�ǐ�Ȇ(~����U)�^�a��#�FB���H-�]��OԆyS+X�8_�(a�af�7��;9^[ˈ*�"��m���>�h��JQN�S-�cv�4e����(F�3]'l<�ۣ�͗N��<���Ks�����IÙ�`�6]��:D�髄��6+�{eK	�z;�6�;0$$�d�n�ZM��<傂S�aM�M��,�ǔ�h��.D�bnl��cv���[)�cI���cMGMuI{�ݥ.}���i�O�H�w3%���)eM�/��+�ںҮ�t�n�H�קA'/�q�O���� <�[����8 ��N{Z1��#u�螳��=�#���X]��ۇ��I��]��N;mZպ����qV���'=n�@����{�vhhܺ��=��=��;l��2�#~�/.L�lf�TcT�����~?�x��Ŕa��"%	e�`a�N�a� ����BYe�a��:a�a�����BYe�a��:t���YEQF<K�h��w��=�Tɕ����Q54���X�ȫ`�9�����ty]�\b�#���]�g���֛���v�;t�C�tr�������W�ն��t�c�����5C��!�q�Lp��<�n��l��d���z�\vݻL�^����N��v<��5N퐱�t7l�{ui��x�cYtSlzް ��"�ɗj����c�]���,m�Ȏ�"�����1I�ks3��DA��?m�rƋv�B��m��m�X�ˁ~Ө�����w=��Hd6�i��U�[��/N���<@��|'Gٰ^�[
ziC����}"���&x�N�Rͭ�z�0 �v�~��[�;��O���M��	0Pೈ]��!_�.���IU;�&����燜L�~��Fv#b�eU#4���Px�9�x'ux�^k����a���P���@��t�\.0%�^��O}��⊢�x�hЩi�=��ɕ�QU ��!B�c�3�:J2ϡ:(q�.�����U9y��v2�d_6���NYk����@WG�3,������gD���F/�H�y/Z��87��C�q��7$>����>B9�o7�8�a����ǽy�^��=ى����mc/JȞY�ӧ��L��Ä���C�����,F�q��Mt��1>ϱ�F;K�hT��2zDrN5�b��S�	�&B��9""&����W'�,dV] :]�R�*��壙%��m�ٮ���w�Y����+�/%fj6¤����H1�m:�w���-]��I/y��ӏ�鸨�4{w�Q��^_~��3"xpB�.��͞�vT�Q����G���_lugvgk>,��Q�F�KL3'�G$�������y��EB�Bľ�9>����T,e0���GV)n� �����B Ah)*މp�����Q.%�6O�w�o�Z������Y4<4= ��x��״�<�m�A�����\�zd��zpa�$�E�C���K�'�
�������F��&k���ۺ�t��Ϗ�<U�.ѡR��2zDrNo���A�U�<\Wr8 ME���ɉ�x�[����!nl
��P?W��>�i�����|#��OZ�7�oV�ͭky�{�h�����/��������-�;��ę-[y�����9���ɝ���H�|V�L��Y��W3��#qꚽ1����t�bҖ�j�����5�e]�ʷu���T��J����P�&-�x�>�ev�s��ʖH���}&al(����hPmV��x�%���J7^����D6e����>��x�6�R��}��=�����ҫ[98eK���z��͋��{��O�ޢ����H¢�
&4�����l������
<U��F�KL3'�G$��|��#ӗ<�!
��E�GA��K#�<$��AH_t�q�]��0JQ��ͷb�����C=J�y~
�w0�$�H0wh�}�O��u1��������r�I��]�O�,�\sӾ�<:v�Gw�2|�R���:���L2�6LTE��%B裠}�H�(}�#Tt��bYG��v�i�����cs�W%���E!���B'��L�Я�#�D��vB�6��(X|w��$Yӡݿ,_?�X�C�����~�s�ݣ�-!��2��)��$F&i��NT=G*WW�J�6N9�&�J�{2�>�"�N�Qf�$J.�jUL�8�S��ʭ4+'�A�������FLr-^G�.�a\>~�>(�T|�.�©i�d���.vs�,���pB�(T{Gc�kC8D:����YV���8��P$�-�&ڦ�5M3D�vd*��2�'L]�E��zT��㽊9ņ鱅�&0�Ý���lnPv�`.z��'���Jk���p��J�C0�%�\Q�p�O%L=MVg=r�9��ۤJFA�lXg8�����B�(��$
�n�(�ⱔ�O
����t5���>z��ɰ��.���e}�_<o�η��\x��9:��v�}�-ۅ��|=V��|=�����䏞]����B���nw	J�l���v^���A�����5���޾����v�,�X"}�X�v���Y��Ɩ��O}{�c��3�|>>#��C��1I�֣�xz�՗)��Q����褤��'����9=SÎϮ#��q{�J¡�KU�;%@���⠸����/��v-y��*�O�I�ErP�ˇqw`��,
�ď�G#��� -��%	�~���@���������٧�I�9'3�0�Ǌ�R�<*�����k��?{�����7ӲB��B��@���d���I�c5QG��R�/W���O/��W~�X�I�꺡��$�-�Q3�I
DtY
��Yћ�������/y�E��e˰XƁ FJ\&6Ca�68¢�==陸��Yk,��/���u>�ɗ���}�j!�h6J�;Ky�D�P�^:>���� �WJ�ȴ,�iM��V���/|QF���c�Dt����$�""xJD�<��(K�ma�,
ڶ,�#]([(���":t�*�
�8���DDM�{^
�U^�:lD��˭�`]�͒""t�m��b�Zt��v=��ffs�i6""'- ˻�n���ff���偅�xh}���No��&�d�;���K[t��A^�4��P�<j��%B$r�Z�Ks[Eڻw7<_c�0��І�i��f��_�'��1�x]S���$��>L��+e����\�SV�Ă!�����3�HA��Х��za���((DDDD��,�:t��0�DDDD��,��t���0�DDDK,��0�'N�;�32�(��c)v���cX%wE\�!B�F��"n�J�a���S6	Q�P#�9
<�ýP����ߓ�	ACΫ�qҌA�ƃ][M���V�$����UeK�)�4c10��A�z�h$���ah�����$�������c����S4�SG��"�H{G�K�	,�+%��c�D�%��d�G�p�
�
(�_2�i�T�~2:%wE_�e�B�>�_%�r���#�HęnW��OA��
T����e�"0���T����������(�/�6�8Ò)El�
ðG�M�СG
u�Y{�����)>�����t�L���װ|Ll@R�'�Mc��Z~|�3Y�eNj;y����pP��3����"���3�9�O���"��#�پX do�j`��I�i53�{8�b=��"��ēA�gb�[��]%t)I��g*,j��ͮ�;Ayh��`�tv�Ė��)�lf�һztDDx��d�d�r�qy�����B�&D�2����!Y�&j��)��>�5�Sl]*2�vr9�9��Q��dK���3.�՜��°g<.c��}Q���H�4C�`�1��]�5���q��ٰv�H���ǂ��p�"O�#��#�fx�#���ޜ�~rim쏆<���;��3������X��6,:��!aH�Ip�pb���*�C�i]�G��Y�$>�+z���]�QG��R�<*�=�5�YtU��b��V�!B���9�*��4,�{p+��.�$_Ǎ�
*����Wp��C���+��v�g���7�
u� ���[I�.�?v�w����af��!F�e..�SSm��h̺$��cBs�
�}�ur��o;;,t����쐓�� A9���Ag�I�n�z����+��N���<V2�i�TE�#��R�y��(/1�DG��F�����g�VX���˽.(��
�!^C�i��i]�T(f�x��|ѓEԪ��X��Y�������>����uuG�R����9��I��7�*>د�Gŝ&=F��]�/��c!��D�F��`v&�`O��&���Ty����q�(��c)v�D\3��.��=%D��!A��f��Uǿz�g�%*��uK�ʺ���\��x˰ݖ��&I�^ޥ�o����^c���$��-ʃ��>�*W�tC�U���Ih�+��K�z�$�v�������Ju,S���>�.����&��G���")%U�@�d\ ���^-�8z:M�=Ԯ�	E+K��(�g�#��7W�/��.ID�v��h�k��bV~��7�Q�[������9��{	i%�Y�wJt���z��/:�n{�*��ɦy%�Fn6I��+�6�~L=?����g�`�}�p%H�|��<��CZ|��Dh����Rd���u{,�/��%^�Lg��]��>��J�p9���G��J��Q܏��.��Zc.��b'����<�h�J�z����`���6�3!L����mO�R�.����J�h&]��w����uu���N ������h���H� �,
KQY�x��NßJR�^��#5�~��p��<V2�i�lQp�Gy�|���� �.�`�g]F%w��<0Z���$�h�#?n���G��x��������huEi����4��[t���=��`_[��)
D�A�,��ë-�d��ӽ��n��^}:���!�!o����凉�Yz-,�I�y��ll��{G��T�"Qܳ製Ý~,����i�lQ~3đ�l�r��e����A�dSIC�T�`�Y����/�S���~��JkC�jG�����W�O�QA���n����z�,�$��,����;O��v��|cs+�b�S4�N����G��i�B>�m�r0�-�W�h��(6� ��h�1
�Xyle|4:I�������~���O=�%���+z7��Æ����Ob��x�;͛��u��<A(�!�}�R�Ns�5�2I�8��q�Z�'����$��&*����ƚ���L���~��!�Ǿ�]��*,(*"�Q:�J��H!��P��HZI&�q|B�����l��v�	��F��a��?�]eb��]y���]������A��iCI_uTUU����?������������E�a"*'�����^��	�7ɦ��p$ � �{��LL�!0̳�2���0L�,�=�c0J�0�L��2L+�L�0�!0L2�L�L3�0L��$���J���112�̓ĬL�3���30L���30�L���+�L�$���10C�Q����&&I���fV	���bb`���ebbfb`���%bf`��&�d�&e`��	�d�!���BI�I���&	Y�&&���`�a��ba&&&��a���&���bb`���fb`��&	��d!�G	�b`�e�&�f	Za�	��fb`�&b`���&ff%a�`�f&&&	�bV�	�bb`�i�V��&Bbb`����f`�	��a�����i��fb`���%d�&f	�a��&�fbd��&fa�b@ �&Y�`�f&	��%e�f	�fa�&	�`��d�&	�a��&Y�V&	�b`�f&	�e��b���

J	((����)(���
JJ

(h(�������
Z
	)((������F



Z


	V
JJ
)i(�������
()h�����������FJ
Z()h���$d����
Z

�����Z
($a�������(��������


	h(�������F(i()((((i%X((())((()d`�����
(�����h($`���������F(h((h����F


B���
	(h(����Xb"*��Y(�&��Y�f`0�q()���������"��*b�(Xh�*�(��F)h���(h�F))���)(��
h�����I(h����Jdb��J(�)��F(��������Z�44SAM4PH�MRQ@P��%RPQC#�3,T��%�RJ�E$M4RBԕTLA#R��LMPRH�M4R�E%23M���䣃E%AMD��SDC+D��R0QMQCEPT�MQMM4��STQR2SAQ$��T�AA#PRPPU--�AIAAIIA��:
)���P���
�0!*�°2�(0�#ƺ4D�,�B8*@¤����(�����$"@ʰ� �
ʰ�0�C �2��oP��H`ax�paHade`Yub2�0�3+�C �0�0�:�4!!,0��`�Ù��B8�C��Ä��B@����2CC4�@0CD$�$)$D�Aː�B�LA�AA0DA@AB�AAA$AA#�DAB�AA!I
AC$A0K��I�A�AA
PLCA0DA0CI�AA0I�CP�0D��DA,B�LAA�0"!H �	�`��`�`�H�(" �"`�H�F
`�(%��"�� �"	 �� ��!���
 �� �X&	`� ��HR  � �`�	!�RH!�X �B	`� ��HY�e� �X$�!�  ��	`�`� �	 �R �X%�!�"	�aH� �	�%� �	�!I �  �"	 �" ��	 � � �	� �
�& � �&� �&	`�	`�& �	`��	�f&	�bd��dH��f	�f	�f`��	�bd��fI����&`���&&�fd�"bd�&	�`�&��&d��f�d�&I�I��	�ffa�D��	���bfd���a�f`��dI�I��ba��&��d�&�&a���X&	��fd���Bed�&i�i�V�I�ff���bfbfd�f	X�a��f&!	�f`��b����`���"i��f�fbVf	$&a
fbfBiY�bBi��.1Gi���H`�iY��&�	�`�V�&I�	��bb`���i��f&�&%f`�`�����&e`�&�f&HB&I��f&	X�&	�`�d�&IY'X�2L��4̬,�34���3 �0̓3���0J�,��4��4�K��0�L3,��0LJ�LL�L��+�$�4��33+�112M0�3��0�2�M0�L2�0M10LM0L����0LL��4�$�10L��L(z����z0�~o>��}qL���}`�̂��2"�Ģ!@n���%�?�?���w����������Z�?���7��>���ϼ����׏�k�6����a����lpZ�߿��S���a�?N5�E�|����8;��)���
l>�'������DP_���_�y���~��@���!��=C�$��� �3����a>���\���������.A���>�/��!��0��=>���؈����~��Ԃ�}���L?����������"}�����9��d����_�I���������Ǟz����'�O���:��}�]���IO�����u��\�� g٣B#�@8�Qӡq@U&P�D=E\dQAD���DN:6g�``�u���3X��~��pt;�����i���O�0��1  ���!C�1�P�(*�����������'"��S������w����=��'�t�0f��7�_ڄ�'���W/��0�(.'��ai~��C����/g�?�����A���o����8Cݙ؏����r���?�'�D���G�����>��?g��oG�>��(��h�0$��W�Z?��?o�g�xtx�?_K��U�l��(�����VW�o?��������mO����v����|;K��0��?\ACn�>ꈢ�:*��8	�&��UT `�~�O�t��v�|���?ޘ࿇(��skˮ0��A��?���j�{���TP\P�?w�E__���ToǄ7�������lO��7�� �����?�?��|�?���O�?���It)���Y~q�A��O�/��>�����
~s��������D�8E���� K��W�J��a�������������a���ȿA8�o�?g���iC*Q���� A<����?L��C��G�������C��bh�\�?E����u翔99AE��o�~����1������?Q��@|~��{����������
3�Nj��)����N�>Ϣ}�� ���YOۯ�Gڽ����~G������
�18\����F/'��y�1>���6���Y���4��@����W���H�
a���