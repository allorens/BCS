BZh91AY&SY8���ܩ߀`q����� ����b)       ,                                    ��
� ����   P   (   T �          �       �h  ]� �Q�@     �  
  @  �   P�@  �  74   
�� }�B�mq�)يse9��g6骦W :��Nv���n�鱵�;R�Q���J���lޚ֝��-��1|�   �   �>����zδ�U��j�M�c"�Y|�x�������wׯmm��qwӟ6�t�XR����Pun ��v�E��u�O6�)����SҼ�E P �  ���    P  ݀�}(;y��5=�����ú�=:&���@w���g�t��1������=���<ҟ|�e��˥*�޴�� � �   GzS���w<�R��� ���-c��v�4�aGZf�����B��x ^�U)u���4�5+�j�A��^    =|   b�   
 
 >�ON��{����z�-os������Xz4�+��
t7YT)���xPZk� ����h  �_   ����y�������M�� �`t;Pq�� ��8��֥ ���'T�    {�   Y@   �@(|
�z�J�gZ�j��S����{� �P)�M��6
wr֠/x =���W�@���z�  |  ^��9j��S�x 
�\���]g@H����� �QKXt���4� -`Q��@P��� (@

  

�
Mx�4�`t邝v�S� q@�wS�кԮ@�aA�����{oP*�<Z��    /� �/�(y��P� ���N� �+��9� q��(��j�u����:i���        S�JT�i�F40�#F)�)*� 4ɠ @  5<j��*T @    ��U*!M�       %<��A*       �4)MM�E=1#54�M4ѡ�'�}���Ϯ��?ju�#���pA�<�����Ԡ���?X�*+�>J�����G��W�}�`����?w�?�|��v~G��?���T�QVኪ�8QE~�M���rJ���_����9 _ɕ��eQ&EG�eP~�E�dP&�Q�d@vʀdv���Q�*��(�E�
��PGl��*"m�6��a�.�Wl�2��l+�U����"�v»e9`�.�l��(��;a]��Q� �»d]�.�Wl�m�{`]���l/��Gl��"����E� ����"m�6dM�&�l���(�v�2&�Sl��T�*m�6dl)��g��"m�6�;aM�&���"m�6��`��"m�6e�����v�;d2�e���l+�Q�"���d6���l��(�v�;e]���6��`]���l�A��v�;`��Sl�a��l��A� �v�;a�p�2�Sl�� �6ʛeM��2�eL0�l�� �v�;`�'��Q� ��;eM���A�*m�6�;a�6e��XSl#��*m�6țdza6�e�*m�v��eM��l���m�v��`���A���;eM�8av��e���l��� �� m�0�;d���Sl��Q�*m���
m�6șaM�&�Sl	��
m�`���l��T�v�;eM��0�a�&�Sl)�D�"m�<dM��	�T�"m�6��dM�&�l#�A�dI�6�;d���l��@6���e��G,��Q�"�v��yal(��.�Wl��
�v��6Ȼ`]��l��� d0dI���l�A� ��������YGl���"�v»a�<��Gl��� dC�E�"dL2aSl(�XT^Q^]���eDv�����@���4G���\�:z�UPm�Ji-Q�v��(�I�D�0�%�d�Y`��@���jjN����g���7���Em� �����q�wk�n.D�t��s��YF4���y7��M�+&�Dm��n^�|���WLY�cqO�S�us��P廧r 8���vW+UO�0��R���٩�n�o5��e&7��R�N	s�k��ž7YrS֢a$�?�O��nn%��)�f��䂣�&�����B%^�n�BRygJ�3��!��ـ��n���)Q��ނs��B�-e��y�9�Bcv@y9`is؇jU�C�]g�MLo\�;�[Q�0�X��5.�M��ٰ,ް��:j���8.�'85��4�X��\�[;"�h��k���p��u\X+?h�q��c�!��U��d��S��,���轝u�͑%��ۙ�U@m��Ծ�G��-�vr܉͖�坢,{��"r����T���d�f�:V,8Zf����\�#c� �4j�S�P�e��� ����l���ک���TE�1J˳�x�������}Í�%����v�kB�}���r�3r�BM��/�"Պdl�(0�W�LM�ǵmZN�Œ>���t��M�w~\�M�cwU�9{�Z��ߔ87��6�S�����Z\�a�j�-\or��p��sG�0��Pyڸv���u�I�d�Y���s�I���r�8g%���eݝ�����Uz���Cw�w`h�8;�ZĲ�'tՎ-���&k��,=�\|�̧3F���qK��c��0LczѺ��2܎�w������۴��%�jl���C��a�\����%צ��C��j�P�	�s���bh�0�[�;���E��j$[޸���#ѽ�X��a�	9�K�o�
\V�ۯp�ڧbo�9�w��S���cwR=#���7[�r�W�Aو̨n�Ѯ�X�o-���|��B�P����m�Vn��I����.��/F��'���\�svp��|9�}o=7�Ns�M�N��#�#ю�����I��-�L�ww��<H�+KM�4��s��zo)��k�\z��Q�}��;��%3���x�i#��i�ÖR�0	J�X�j���p����$�{�Q�=���F^��]�����_l�P��M�ý7)��6��C��7�xн�n<�h.V\]�����u,�]O��F�c��G0�Fኲy7K9�Cb߹f��2�����C���`Q�&V!�u�;�����uɼ��Y�zD&(��Y�"	�9;,;��F�@��Ig;^�h�\5����M����EED�s'.�Q�,�_pyT�u��;;�ѥ�f�о�,�ETb� �Ụ�K4ͽ�X�����m�
�r9�-Ëm×c��R{)9F�j���I\��˗* ��F����p���x�:s�6�78���d����=s���gC�.�� gW�ٜ�Z�h���]W:�O���m�/0;�t���؎�m��8F�pj�ӣA豕�r=J�[�9�j�8�:�d��ﭙ(Z��v;�;H�c2�>�+N��$���[ׯ_\!9�C��¸m#�暱	ٽ�t���{�����=�tǞ��v��ӂ�k.-=[��ʖPO0��<vI�s��X7�e�ɝ�͕��GT=Xzu�v�8��nf�[�պӮuϖ'�q�X�$����@���p�L�	gW��A��͈�v�� nG�{�[8�.�G�t	��;&]X���t�2E�Z�]�z��H滲4��*F-�6NS�[C �{�/����;Q:C�r����r��-ۈ��RB���&��3C�3���`�ŦrEmg$��u:����P�F\���2�2�wVv�aw�.w6���<�2+��M�D�W=��
jR��-�"�N��Lt=Ӧ%�����H�*x`�p+��C3�Pr�0��8���sƥʹ�o��N���Ӹ�F%���c����{LĪrNݝ_���@#s�Z���9]ِ���;��F�O	.����\��[a;��QJ>
�t]d.�x^�*��������P��wp]s�QGm㙬װq��y.�w��K :���؜4��@N�	w9�w��s]��g����1�98�=�(��ok�]���m�rq�~�ͤ9�&�e���N��n(2�;�����=⩛��>w�<Fo�����.���@-��j;K���wE:���y]�'#͢��ެFv֮洁Y�����Ky��}�,զ�wz�4K��{�\s�����F�w*h,=92�y7H�-נp�g U�Rb�0[���%�pE�u@�軍��1�3���7�위-�]��Kw
�A�C��^MD[���7Wi���{FX�\s^ɷ"�pѫ�#f;3z��gd-������6Vow�~i[&�\-��j\#w��͎��p��'ˠ���(\|K��gJ�X�B�|gJ���c�T��&�&� �kچ��Z�-dnr��;(ӏ�J��+�ݳ�ˊ�KYz�.�0�1�Eѝ9�t�r�,Rv 6�»��f�v@k�݌�+�1Q�|�e1�h��R���8�TخޕQ�S�2�\ﴖ��S;[�:�H���5���g�"y�{{t���m������w�������q,�3GY�T���ͭ�m|��[�n.�N"�c棜�M�s���x	�iSc
� ��^��Qɼ�`��e[�ou�ա	��^�]��{�r�]�\nv��ؘ�$!;��e�6ׅo.8�h���Y@�7-BN������.��Mʢ֥�	g�]�E���Ϧ#��;��'����e˶�` ��=�2�8���sj��ݰ�i��X��He��mE�v;�Ӄe7Tuv08����%�]��u�9����V؎�q�V�t�:qQ����yj�r`�f�B�����h�,��V��5ovuܬ�ê�(�q�з	g2,�f��LC��m����sr�R�i[��7�Yծ='rcFI�.UJ�3wT�D.[3��3�nB����n��{�ݜW,�]�>���+��ۻE݋��Ӈn��'�M���6�R޸cǏ�38��A�X�L9��������R��6<=þ�wj�[z.�6���њ�9�n��*�Vm7-ZY�1C;h�:���vw$&C1��W,/P�uQ:�Ir�'d��ʵ�75�49=��Mt�j�v�T��P�z��q�瓅bN��7Dj泺�ݯ/b�%Ĳ��[f���-�������� ��Hy�w#�8U.)0�o�vi>E3�zM�������NOS�T�v���jǓ���V��b�.��~]��\b\��:�{v����82^	��ǄS �����Wr�]��?Mܓ�?/o/��X��gx�A�S�1�5�X�9��1v������v\��:C15#΁�����u�ƶ`M���b%�dvb2�$������ݡ��3WM.w��P���,��kνV��j�z�s�o>mgg.�#�˫�@��@���.���[�m����4�	7:�$�Jd�Έ%s�f5z��)�Ζ�e�泧X9�s��k\z��]@�Gv�����;D7�Eth:�4ʥ���Ǔ�e1b��)#y�x����z��s�������w^��F0l��TҪ̛f���:u;�.��kA%�pwg-�@�?����8�����ZwNcL�Z����8�����dPV�����Àq|�st�0�˳A��J��D�ë��]�)�c���-��NȖ��0�C��N=�A_A6�����t띻kiķ��3���XԞ�H�v���3$\%��qZ������Tu�{Rp�.�΃�ߏ.�G��qNgL�oZ��1\��(�S���;��稌ة�8�{ع�o� @��;��@$�7���=ڻv��;�6:-K�<X�ʌ�D�.��J�޹Z�8�8�����P�_>5[x\y9�]���})�sgh�OVTSa�cg3�I�:���%'� �;��%���;wT!�EHg��r!5�ٳ�Ը1qh��/��5���۬b��xՖ������y�93R��M�����Z�]�e�Oe����%6�we����KY�Ok�R��{#���R�[�4n�-3�;��Bh�����	��ڸ`wV�t�!�����/H����ݬ!��/�$#O�P��/��x�1����l{D4�c�[n|���W�[ D$m|f�y��y�[�6)��a�=�Hܖ�]1 ���5���z��=��"���؞�x��7�Fkn�l�cwx�f]�
U�M��N�`��:K>���<t�q��״XI��Y�3t`��p�p�� sex���FcOw:�ǻ����Qۍ3�nV���BQ<��r�h ) h��������f�x{�/v\�d05�"��꧜0�F������(�%�z���Lm�����s�$��ę�m���N�yi��S�T5]��(�f���des'��:���'9ͽ��nV�Zv���Ev��[:.h)*�ePR/<�t¹-=�2�l����3���������K9�S��Q��V���w�e�6�`������ŝ�iݸ�7z.�7�Ԙ��-9���w�-�j�F�0K�z�b��nHX�n�^�����+���,��IE�W0��׈D�r�fֺ�G59�Rˢݥ�Ǡ��7�&+��;���f���1�X��ɂj���ɼQ��
�Ó�W/oyQ�> #š�t�+dL]�y��n�݋�C�Q �s{�ۚ���v���e%>Gp�bڦ��a;�A����hmQ�����('f�GT�I��u\�7���=��m2lp��}��_c��5s�7d�UD{�����=׵���nn�%R7J�=�)���s#��Ϣ����6�9��Mk4;��q}0Rd�wݑq�:󕌇雸7W=u���m�s����i�@������ᜪ��楢��E�g`��ӗí���zٶ|oi
 aN.DِriswF�ҵ�7��[_X�ds�3a��.�H�P�&	ȳ��su���WM^�{�C��\�Ӌ�]��JR�s#<��&���%c97�A� ��]�F�f!�v�*�N�in�4������sXq��<կX�[ޮ������\{4S7��M>A��V
"Ŝ�#������)<��n�%́�]��w�C�/�	�ͤ�o���y)V���䄪��U����å����;�A�x�#�wn8r8�#\np$�!�7-&�t;��÷/U��v"�M�N�`6�td�3��0Y�tf�/`��H��nu����p}c�G>շYI�fs"�B�h�2��G<ųS�5R��۫�8�ص7��y��F�)��5(�c���3b�����(��K�i��c��5+(q+P�n*ɥ�����:���t`[İĝ���C�*�C[��4���3⥄ݚ���Վf���8\&n�/`��4?�n���v�N�*ӛM4���u
7f�!7y��K�5�о��8��ջ��+���r��ƴX�n����c�m��ijk�hNq84�S�B�����ɜ�\�|�H�w^庖�X��K�ͧ�N�9�O��KFN��/f��5����9���jY�V�h��@��R�*Z����S�ml�l}�l�5{)wr�&U�����M$K�4�{(n�tۅ��z̭nXͼq.���K4��=񳶍�T ;�sqsj<�P�%i�v����,�\��W�|���'�Ң�r�ۆ�7��q��K�ZKg����;:�l0e�Z
%�ɤΡ^>�La;�-�G`نm����ȐÅ}��0�x��1E��>5��$u�1�R��iy���zU�i*n�@�Ok�y�2хf���wN�xv7�cVTW+��\�t�Kx����S���̡��Lѹ_n���8�S[-i�kz�;�7.ۏGt�7^�1�;.d���@��)�K�8�qT�N���/,r���i��r��;x�YΕ���f�{GTx���i$N* zl��v����S\ty'�s˲��8���/5�PX���X�7�����T���)�Y��dA��P,U�p�8>Zm��F�qG��WE75�.�f�Ϊ����D}�!��;�8��3�\�uҨC�v2�}A������('�YLG�u��]��։���=�B@�Z<t��2ڃT��e9"�ˌV,�����M�qL�7	�l�Ğ��[�s�_ȣ����W����tPB���\Q=��~�ǡ�6Rr�,�3*Բ������
LZS5�>�®�Ǜ��U[D=�rq�U���k|H�ݜq��v�M����$�"_{��܇2Y����{�zq>>�i^��� Ƀ�������{��-ʣ
�J-K�jT)4���#3�B���X*�Z�E��e�v�D��Ƕz�W�:��X�O�x�4Nƫ�zק��w��^V�&���2��m�L���x�^�� ������e/T�����E��}����@�
U�Nc-�V�7ȃ쵉Ȝ����O`�߽��ʖ)[\��G�{"G�������_����	�_y�Z|L�||\0x�����ˀk޳��# �Y<~��x�gN�7wS��9s����]Q��؁��Hu9��v�>���G��t��M9�j�^�N��^�3���7�dU�	:�����#g'����ߎG�6��:���O�"%"�	�@*��UJJTZUV��\@�@� �Q� ZE
J� �@(!JZ�$Ċ�$�(@�8���U)D�(()D
@)q*)J ҂8��B�G
�ThT � i@iE�(� )� �P(\@&$��
!H*Ы�(LJ���F��ihi( (J�� �AJ�b�Q(L@�b
A�ZQB�F�T�R�D�*8��
�U(�)iPV���B���"�_�}��8�k�u�Y���Q�?��13�,.zY5�+�D0	q���^h�S�y>q�R�\˂� ���~6#PWخ��`��77#ܭ��n��F�	"�M�_u���FⴒL9@r.����r�o��*���r�Y����%rx·�&i��b�ĞVĊ�g��O�E$�?HT��4�+c�#~���w/�ț�Q�P$�����cJ��>IÃll(�l Y[:~7�>�}����0���ҏ�ᔅ�@�}]�����5�ɝt��_�oo�|%M���7�����ε���˂��8��U����}�QD���E��{�'�}��? ��=���/��1��;��?��[����O�z�v8���Soe���`B#���8ޤf�E�sܛ눤���0�y�K���<�ٛ�ϖr�g��}4���|6�æ4���R��s�/MMb���%���Y�
����1�{|<{z�W�s����'����1�y��m|��{�&]P�#7��L�y)�xK8.�j��m&��,�Z��wp�=��D|vs�c�P޳�ӛ�J7��{��z�iC�`���=ا�y[9�
�͈`�+�٨MXv�Kx7����~�v��a
U��$��b�z�c{��g��������.����g�����������{ncө���ͣ&����e~;j/f�����.��y��<"�Gj��<�<L�Տ��T��r��]��0�+��W%ܻi]�2�y�j���yz{�A�ʶ�f����+O�*R�n����~����G��7�z����iWx�P�x�s��"/�t��$��o/�ۣr-������:���]�N�Öb����W��>˨�u�ᄋ�ش���"[#s�3ׯ([ b����]�u�l9��k�l/>��i���}%V�άA�Bc�g"���;��g��x/g��BkW,r�l-w#��T�W�W��^≾�qj�tcŃ")bݿ]����},�{�^B��u�3z����=������G�����k��5����;Akw;5�e�z!H̃fj^����4˭x�oN���MZ:,|�)���Oۚ����F^�8T쾏��-�x�g��S&�e��-*�/�	�>�?z�.n:;�oo��ӿ|8Ş]G�+��\�{*l����{'i۝Ï_�wk����-��#���jh��%ȹi�w�����eP�3����}�0��wU	͏�$���b�k�������+����by���C��a�&���noB��慔���q˟U׉8w�;˯Ӹ�SpS�i�F�
_J���GKwя-�-Q��p����v훽�����.A/{(��#�yw�M�aq��]ʕ�|~��@��Q�0q��l�Y�������k��.q����s�U���U23�}��}���u�G[�S}�������Oq�L�!�=�:�B�����{��'����z�y����$�17v3_��״������&�����F_?p�
�P{����3�-���G8�w��*0"�ԗ���s&n�M����}�b����k�W���G���w��&j3�����9�h��o��u��[�{��=�T��ǅ�:�r����O{s=�.�w%���TZ07d���sva��s�Gob͐�X��<���i�sE3Nx{�FUWG	.T�=�'bp�{�5��-]���`�.h�5� C������{�ww<�F���6z��C�`�\]�F��`|�m�,��0f]��ǡ;�}�Fyk�*�v��߃9_5�u6�Ռjͭ��z�`k�9N����H�?a���=26ߗ6���ޗ
��0�Ktnxv����L�t?v��"w
&�{���\�~hz��=f��vEm@P0�Y��A��l珰Es��a������4�rx�ҧ�����=*�b���*���ރ���i���;�� �I�)'�wuz/5�ow�Y���/`��[��B�z����--�O9�|�M�)��vŊ���h�������&�S~!f׳'9����n3F�i�\�#��&�5K��1��Շ�H%k��ޕy��a�8�E�):�g���L8�r�Y�o#ܰм#̝��j�d)͢�9v�i�9̜�nҏb9�s$h�7p�.��e�{o%���oȬj��nE~�پ�3�l9�#f��{<��� �{:��s����bu�{'Ǧ��#�N[�;=�������hS�z���L.�s=���,k�?/P��<Gv�Y�3�r��3_q��;@��gL#�}q�ڵ�7���R�ݗ��q��[�q�!A�)�K��`�>���*aЧ��]}w�:��aQ��QnS���C�V�� �;�շ5���� ���!���[_N�\+�W�zgfR���T�A�Ki ��ˣ�U�Ǽ����|�������=��m�7���㾣pZ����<�?`�.�xl.�wC�r����\۽:�~����7ۗ]��#Ɉˍ������E}IZ�r��+4�����8�$���@�����M98s.-�Ɇ���#@�폷�q�wz���nO��3�n.r�5�-�fU+j�L���E���`�"�]|��רx��[�9j��j����?{f<�*��=;_{y�˚3���8=�h�4�O�ۋ�Y�C㜨���ğ���:B(F���uz�>�s�\{p������6p��;���ы�=Q<�3vL̳�����'f�c���4��g��cU�b�,����U�'�Y��b�T?�R�>M�9�#;5a�q��e���/�x�;V\��@�Y&�;k�H�6\�ߵ��4�˽!g���f��re�����&����W������î��E�gf;r�Gn=w�ދC�F�A���t�����L:S�8wT8xps9��j��^�O���ξ���&3���NP�G��gI M,�M����7�m�2[A|ɛ,�ߔ�R����Y~��K�o����{�Z���u�o�'���ck����w�+����} ;������-���b�*Obڤ/	҃z��W/���޼�l����VA�@��xb�����Y:����g���Ԇ�H8��OŢ��э�ە\��o��~��|*����|�����l�]�ɾ]�L���f!��[N��/R��"�wn{iVҪ�b{<�y��w�G���2Z�/�8�9=��t{��G�����zG�^%��(7ڸ�;�N|pK�p��Cb@�z�=~�^TN�c4�{����u��r���]F���b���$�y�����=X�sFU8t8&�a[.ga��z����sSr���%�I��.�͞��nX�o׽���(-)=�J%,���aH-��n����X���=e��������#�-�&���z\��`�v�ӆTgA���c�:j��E�_��\�I{�F{��{*Y�y�0��=aY,pӷX���/[ΞgW���B�v�vz�*�9{�!� -W��|tM�u���>>�B�r���e�t�d���ߎ�U:��$p�⎮ng��{7)8��H��^�|������C�_��m 1\J�Bؽ��O�'W���$�,ɉ�\fL�3V.��nSW+1+��F;��q�A�}ޛ�ݗ�+^��Qv��wY��ȩs��X��Kgj^��|ŷ�X���8!p����I�{u�'�.�Y�o���X(�5nx<5����N�������OoA�5���Y�_;�1�Z3o�r����k���;�����n��=Ӈ����1w��{LJq��w{��x&?k�Nѝ���W��n@�/L�(S6�f���s�jxި�Dj��l�ϗE����^��/����y�4upoS�����#�N��C���2�@5�ٻԓQ'5��a��p��8%����ѭv�ؗ��h��9�G�H��/��Ww�����v�=�Ϣl<�9�$��^X�ׯ�϶�$����s�/0�a�p �`1���{���\��r�}Q�^��'����'�;N�ֽ�݋��b����\�5���<}1��z�����8��|�׻��={9�k�sq!�ܧ}�b[�~�3�;Z���W9�<�6{�u�m��8+Cx8|�>P{�SR�HdRd5��y�^x	��+_�YSq�Nnu����wHZ��P��r�,����ǣ.�{ޱ���(.��;�=>����:W|�Yh��e��{�'�c#���j��4�{��ǧ|ώ����yS�%U�づ]�/.�X�V�)ɧ����_}|-[���8�J�{�g�����;���_N
��#��x�n�9�v�C�+���}qs{ޣ��䞞�5z�L�9Y{|^\�=�^z�:����ewY�>����7�� {G�ztv��	���{�^��}�f�ՙ�}����$U0�b:�rZi�{�P���}�kJ�jǓʣ�^O.=H��E5�j9��oԶG�������<X{��W;�%�f��p۳1K�_�^��[�wn�1o=�D̻���;�]5/D�ư�<��t��}ޣ�ʋ=�.r�����F/ayt�<dl1�r��S�����sw<��0��ּ�^'�+��@���9�9�ޚh� �t�(;��%ٓ.�T»W��MN©�i�ό/%q||v�x���~C��Bc/�������8�݅����_e+�0�^��>/�.������H�v<�J} ��oV��n�o>�E��:��n׾�P�Z۠���c����jy�1��X��T]�c{���x$M�]��xe�wq��1d���л����'�������K=��*XLד8����n���^�M��)eI�/U�
��OƟw��{®�Qa����-[s��V�� MNY�$:a��aU7k^���C�kTl��ua����K���ec~>:�lq�T�z�v_%ϼ�sUy�FzAݓ����O�=g7t#pqmr���K�w<������y6]��L ʵ s��{N"�o&����ݝ�{
�u��c��ۣ{�{�!����k�G���M�	 �坼4&^,�x��no��R�F��^���^��_��]8��ڧN�?<6T���g;�Dz��|�������b�4b��1�	�k	Nb�V�e�{�b����{y�%���b�<p'��=Zu)�1y:���3W��ӔՉ��<�V7�2#1ڰլV2�����
z���}�Ǐ��;3�u!aX����;G�m8w����m����g]&z_�%�8�bx��¼���H�!��Y������c[�G�Z���ɯ�q�j�����������tʼ�^5�Ͻ����>~��������Y[oۄ�g���CW�||�ܺ6.����_�O:�w����'x۸;|i^#�i�(�庫��}�
�Ž{�QѲQ�����}u������w����E�c�Ѽ��m����8���h;d\��
��)v�`]�M�����l��9��7Q^��5�;���r֟������J�����L��+���ת�۰q�e9�ݙh7Ӈ�t��Dv㍧p�!sw��=�Ps|/]6B'g�J�W��m�q}��0n�0�$s��Xp,��oN*S�/?v[Q[��T�p�>��r���Y��X�zmN������9��������"����������O�|oקN���>�OC::�=���G�omg/
�{���� ��\�=*�C�\o��	`�>���[��OH��\�v;���Ѭ�yh���ַ_gQr��[��5���[�_ll�c{+�=M�VZݎ,�Y��_]��J��Zȓ�zY(��&OYO�x�Vo�m��_�T��ՙᾄ����Ν�g�0b�ܑ�=�pc���}ӥ� ���9�v�sG
�{i�s���M���~��b���=�B�{��իފ���7��ޯ�&�FJS�=7sV�A�&���)�e@���7��.O"b����<�î<]&�׷<�y��-GK����ʨq��/%��T�*�z~�n^�3���~��vz���^�E$j�{I�k�Id�}�Y��M'�<��}���`����v�ɾ�áw�8Ǯnش��Y�P��	���4������L���:�`B�B�o������ؼm�VM��E��e�ɾC��/|�^}0��F)t_dD�H��;��se��`�����h��F�d�©<g4���d��ۚ�����~SB����ݲ�LdY���S��ӏ�����(|�-C/��>���W��f��_
���0���!�[��6]�&x{�==��t��xn٢�S�9d�#���@o�L�e�^I������f	��G���>��3V�{C஌
��T��bbaK��noQ�U&{7=H�Y��W&��}|�Ӛw��в���7׊�<�ޔ>g=<��8&uϻ�<y{��^ydvQ���o��~x���t5��zv��j�DFWK{x�v-�7+f�g�ݝV/��2ߒQl�'O�_g��y=S~� G*i�q��y��qo��poc��]�gg����?C+[�a� ��#�S�����r��8`�p�����/{���>���O_p�w��}�ikB�����&R"�T3F9��e�U�j�^+q�w3^E���;�g%ٲ�=� ���J�%�	���H��}�>�R5"徽�)�&�H��Q=��FUjίW����:<�ޕ�Y�����]*oe�CfJM=��	4�^Q�>����~�����>81)��Lג�?{b�q���i����7�v�p�Z`�)�w���1{��p*�r��V��/����͝�<+|��1�=�[����ˎ�׶zmWt��3�=�k37P���Z�ɀ_����{ܣ��>��]��gVI���K�}]���k��g�(����ˉYS��N�j��&w{'d��'� ���ݧ��y,���;�b<�;6켟��Y}���g-Xs���a�yp]�^om~~�g����e]1���=���ax��#�=L�Y�Q�f;�~9���x�J\��2���ɝ�x:��Z����ϰvu���؍C�bh�S�ƜI}ҏ{R��z�=1e�N7�m���W�||���c�k����'��q�<y��怢���?g����������~��~��~�������������ӧN�:t���t�ӧN_��x�����1c<����n�/<�~%�� ����ϔ��U�?�����;�-aq�YNё�'2X��-���6���x��HS�l�y�^:0-�m��N:+:⺑|�u;v�gE{w@��%��ۆ�ɎV�u���8C�qq���0=�,�1��\�@RE���ۧrn�n"�X�'9����u�ۓ"�v��\���g�6}��k�sX<�mɲj����.vœéV�W�O9�+�6��v��SLV�(ۂN��Z�Z%^S�Psnxܜ�,v{��:��z�u��mr�>�a�Vf���Jt�N�pv�"ۋפ4X2[�eǸ��<O��b�y�%�lC
Q������ �����&��ޫ����`�%�z�ұ��m�����$��/F;/;&culOr�o>�,��E'/<��\���pmv	�k���u>a3N�oU�]�g�h|>֧����q���s�3Վ;s�`�][�n�:���S�ǡ�=��lڝ�eqZI'nx���G:̠��JD��T(�V9kQ�F9<��<�\��$麸������$���\]��#C�,;��^x�N)�;��}F��]��nŌ8���C6���;�g8�j��8�g��[<u��e��n���l=�+xLDWQ"������uƸ����ܨ�G"<W!W���ݦ��n���H&�\���g�v���Gg����e��U3�{nӪ!ty���0��[k������)s�+��;���\�F��v�&['r ;IOpv�����n/X�H��BLv�;�pk�'�cs]����d{r�������NtiKIf�Ky靀;m���`̪�����0Rn7	n�F4� ���H'e<8+�����-n�z�x�^9u�j��5��,ݓ[-�/h�����penm��u����ܚp�gn+�V9��@��.�mpl���tvY14q��z�.xY�t܎�ͣ�¡oZ�=\h��bш��p�pjõ�\Ěa9���ĚC�ssiŶ�G��̬�u�H�y\�������4:�Λ.-�b+��cv���su�����qn���\T���7>���������9:�幣Q����d�6wnX̐�ѵ�iĀoc�Q��]ۦ��4[xw��;nzCZ�&7��!ۆ�b�c�n�^�ޥD����eFX�I�qٮv�<�+��!�#{ps�>ێ��y�����{1<�<٣ju����w'&�����=�U�ė^�w p�'`��M�<{rp'E��n6*D�y�u����'&@{���/r���M���hy��r�o�a�ۡ-���`��GednQ�۲�\@/$�he�۲�m���T6�g<�'��85r���c�:��`jx��i;\�nȈ�N����d]í�g����z���<���2���olm[�W�;OBì���(�k��ܑ�ݝ���o@r3�/>Q�{Gk�aٸ��&q�V/#���)�v_,�v��΃8����N����r�6z�z�7p�Gf�͐���箭�#��y�ەn^�3�k��^)�ַg�:�1m�`���e�$��H��^���;���v�]���*yh���%���٣��$��l��m�c^{���#��[<�����9�a66p��k�ݎ
Rr�<��i�p �:��λ����t8�Ju��i�0�g�7n�a��	̝�X�!���+�r���k��Bݒ����{e��s��6�!�n��'9*p�x.7N'�`7+�᰼l�;�!^#��P��m]ix�;w!����fr��!������}���wi���quwav˵�'�|1뎺]�\���F}�u՞�Yc��\��u8����x'n1�]��9��b�]���p=C��c�۷;u�tg�[SY�}���gɻ��=��8�m�*���1���&�S7��@F�����p�[z��۲ɂ�g3��l�=����6��8�n����;��B=ɭ��;G[m�mmׅ�n�����k�tc�v$�tu"�[�Lz�eO<���=��颡'y�ꐙ0�K���Ǭ��2�lµOZ��WH�������"��9���r6U*�ry�Z	�v�l��#��v������x*K���87��Z�uk�F^dn:6V"�m�c��X6�s�댷@�g�
������R�6"�X�ֳ�Pێ�pq�y��Fy��F�ݵ���OlhLm��l�8��㶫�bp���r�!���s���.1�s��E^j^�<��񵒌8oc��͕v!=��[,��9�x�F�6�";�h�p�ua-���<˱Yh���uۮ*1�ujQ��]2ۯ�����ښ7����䣮v�Պ&�up���)���=�v�pU��hx�[��Bu�\��`��8�\5�ͻunT�Ͱ�m�(⓵h�Bt���$�u�'�+c�<�x�{]��h�w�{g��R5It��s�N�;]���5��.x���븫�n�j��R2�f�tu����6��me7v��;tk��2n�^�)�fN���"[l�wv:�O����YF3�nι�y���u�Z:z��N8��ivn��Mѷ�ii]�Ԏ��][lo{��Ƿ<v��;���q �%q7X��4\h�vG��G]�9�B���lX�f8���d�F�@r㎥H�q]FǮܯI�e6�&Pέ�ݮ��{5�6���;�͎9�A..�0rXUI�w��{x��55��L�]�((��X�E�����^y{l;�3��"�Nʏ��p�g]c��c�'+�4��q���tn="�u��n���М���yqv���7d=n\i������\n���F'7��`�m�m�L�k;u����c�v��$֣�n��+n���>��<'��Om M�ۭ���h��uś�7b�N��s�Gf�����h�V+��I��n|7ɼ-�4�3�y{�]Ֆ�41��[��ks��5�@��mz���={0 �{!��[;��+.*r�==v���y����x���c�ڰ��ɳo��l���sa�1����޽�.��o4F��C�$Y���u����v��㋮�FWa����u�������/���c���fָ{\U��g�P[c���!u��0D�7Ou�.�����-�C`��N����+��hq���s�"�нo��зn�k�۞�K�n8�2��٬q��SX�팕]����8�1u�"�r�u˸t���8�n�-�	{7b �ۭ�����ܜ�e�ט�;<�<�7lu�tG�m��Fp�ܼ�N��NsS@��3��Q9/H��7�^��L��W�u��pk�5s��aM�r1��$+�\����u;k;�T�)z1r%̉;������g�Gfo&����-	�Oq��|;��U�ʹmF�z�{j��wl��ܣ��#W";�mqs��u�����Z��͗�!�n���_\��>9�=t=�y�w�U�z��5���Y�7]��O��چ�9L�w=1������OG�<(b<s�r�OFs��n�ٻ��[p��/E�۟ۏ6���ލv�i�n6<���b���:k@&�fP�v���I'l!
�ά�r�k���
=ql�Y�$��졧���8�"-uv�cmь�kq��s�\��l7m����#��ͱ̽�x�;��$'mn;n{�����X#Y��J�ϻVg�q�\/7�XE�ɺp��/n��mu6�[Qi��*�G%<�u�R�ˎ�pr����l��ݍ�ƭ�6�[v��޶6�WM�t��s3���Ad�nR��57n�<��N�����M�2�GNtv�I�_-��^r�>�.�=��uG�cr�K�l;��fۻ=�uI�2Y����gv�V�X�jw)�7"\�}=���Ү�p�DS�F�9qv����\��eqҵm����[����8Eè�\�� >wc��Om��#��m.��k�pw&qgN����X����u6�R�»F.:..[��ux��]�{m*>�޼9����q�6.�I��9�i{k��[��k-��{:E�e��c�g��!ݲ��s�b'��=�l(��&Od��i��W�^�6�X����"�{�5�{��nk{q�kŐ{^ѻ�z�t�nw��צ^����� u� �C������WO	6�|#��:�w�ݮ.FZ��1��1���Dk���7���n%��%@fz��v�䋝ӺՍ�ڌ�5�f=]��y�:۵nl�����m�-'�g׋$�DvRq����'9�ϙ�,N�^��s\n�q�Їl�cNW��;�u�l�xMے�b��.�q�=u5�����\�;%�K�1Ÿ^��[�)��8kFV�[�,�>�Wm��Dg��هs֨��dl淞��n9�!�݁��؉�t�ġ���CPSGeކE�6��V5����ݫ���|�==Fc����3�骵t6�ͣy�6�J�w��-���ϛ�H΍{r��C�����<+�ft#!m½�s�m�
��`��ۮɝ��]F6덷m.������X��s��u�������zݕ��b䃮|��ӥ�]k�Y]��[1<Ź���-���ط	t:[R�i��v���q\Oe������������5�	A2��2���p�E\�qVZֹ[��UT���K�稈�0�P,��ЮQP�jyy>���0$��q�|���9�A^m�D����4��00Lb	<�f�H�aĀKNt�R�~��y�Y���f�]���O�C!0�@��x�7$�	�B�M��؇Z6���ص(�d��[h��6�E�Y�j{�!��E%�^�h��Z��qA��$/8K:݀^�m���Fl��k6bZ62�H�xQ����re^Q.��j�UQh�Zb�l�Ur��&p�nBE�H�V#h����j�T��T���!=:�X�����6؜��ݞ'V���!i^H�͙&{�PԠ�N3�Z���0�EQ3�r��J���D���TK+�U1/(����y������V���bR�U��.L�Fъ�II$R�ui'��䇦�n�W&�]HCTQ-t���b�-H��(�e6ݎ��/W�������m,��@�uC(�<���m����(�5���oƚ�Gm�I
���lB��fwU����8F�ت��aٽ����q�Ժ�N(��,��7�&/�c7�a��N�62�mO���D�����s��������]��h�.�[#5Fg�nwmg��r���.�m����	��Sۮ�v�u�=	*=xR��p���tt��g�]��gv;ju��'`1`K=y����i��Cg�_M�����n<g�vvͺ/h�<�Y�y+t�\;�z�[�w�y����nu���/l�[n�:-nGEh�y�}�y�hL�}}��i6wom��.���W�n���|+/8��[����d����q	�p'���I���gbg�������.y^��fqV���Üo3{OS�dM��3�7$c�+==����#$۱�g�"A�]��]�q�[\�#y���k��W�m���(�L�t�ۣ��vwuq��ݱÝc]�=��M�tx��[S���c<q�\�7�-�U��6��S�ۍ���써آ�Lv�h1��u��᭲���d�o7=�f6]����ά�9�p.ۍ��îdP����t�wc�A�=�%V�/�f��-�2z����g�N4tP�Fv�m�����nξ^����6��(�;Q�k"�O@�p��q��|<�T�ph�rv��n]�-�I.냦�E�y��E�+�.�cv�X�(J�9��ASĠ�p)g���A5uB*��ܱ�H�8Lb���ٷrJ]=4�beݝ��˜٫̷u��ݛ�x�%��� R(�贑��7���o#�X�G"n�;6�z\zcr$��76�n�z,r����u��h��b����z�pv�=1�f�s���]ouD��on�wl۾~�1���nn��F�3g�g��!��a��P�5b�ػr�z���5��rLu�؅qWI��f���ԟ�wǏ{h�\n�r�>#�q.ml��D8�M#��6ɚFt5&�m;mL��a�f5"�ְ��W3ͭmX�f�l��6�ؑ�n��dۙ\g���� ���cm�f�0��]���IL��[9#Z[b�U��h�1&�؜���2�K6��.m�u��ʙW����N�EH6���1����[g66��ge5nX����e��h���gs���IYN�#]�R��ăp�O�+n�2?9��GcL������.�;��>�k	��I�|�5�G�!n�� ϏϹ|]w&^L�7���x�@!R ���yx �V�d A�U�����g�ys���I�UZ�	��{0O��C1�'r�'t\�Q׉tQ;4�ޠ��v�/�mv�<����3*��f�NO�n�"���<$2AFF�9���%�����m�������f�	�z�$��^��A���|�1/gb%Y��RB���Z�z���ܳ�#zJ��Z7�$�ك7HUe�2W����p�Z�#-�뗜�2�ۛ��cXm��_]�S/(ןM!�7 ��8��T��&Sj�_f�+�p�}�e�1ߔ�:�"�������{�*dj۾��)�/�K����;�%�#��[�g��tR�`��^7���gM������|&2���o����M��`	;�� �l���h�Őգ٩�`�`�gE����d�e�	"u���H9p�ks%���w��S�s+)���N��77��
����μ�;i6��aW�$���yI7��	N��]A�����&[:�7�; F;�8d���H���um���(2�j�O����<�>۰"��H�m� �I�%�L�w[usi�K��@<��ͷe	����խZ+`�k��ih��
0�ü�̦�MogL��p�f݈+e�T�L�@�A>m���?�"�S���'Eٚ��v Mb�#K4T^��>#i��nǠ)�2�w߻����]��q �o���tYD��2@ G�
�`�K&���Bf-W��34=�5+Oy�mD�l�-���l��	��� v��eyg�z�A�4�����/�`=��~`��6��%��VZv�$�g[]|��ؤ�@�����&S�G*���8Bba��I
��A ,ײϮ2��2k��"܍xM�7nNq8�B�)��h�M�;���VM	�n)�-KKA�{q�mܘ^(�>c�f=~P�^�N�b'r�"��9�?��ث�l��0n�)������-�����]�Em����ߖ�:��d�w�r%�@*�^	�Y�f<VN��͕ �a��7�cKO�=��+$aw�Ce��5��ۉ���ǉ� �+���||H{/�8k�`Bn5�ӻ^������Ϧ"���L����=A5nA���H6�%5�1�zZ�?����'ĕU���Nς�^/���K��M��Xi�63��dR��}��-��cĒ��`�K��s?o�s��]y^��$��g?YzAd"ł}y��{q����)�ߴ?o�{�'��������ֻ��y���Y��6��B�_I
��Q3�z�6��$�:����5�;
�x���^ǠkS�	5��������e`vˏ�~߳f1Ye�-�����ۍ��sv@����k�Ң(�!\�X�B�xk\5�(�|k�I+�n��4n9ٙe���7Oo�z9����?�7<}q���+ClK�$�ڸAE���$���g�#��澼x�P.q�ܘ�P���t@�zd�Ed���)���8���vt�x�S�j���z� �e��ǉ�'u�����T��U���Jb>����V�m���ǆ���'_<O� ��s���Sd�;9�����<�ڛM39�+-q�a
��z�	� ����M��e>*���o�m�)�A܌x$��M[���H'���ؖ/����[��]n����h�ޙHkCSxzC0n��U�<����Oq�� �<
R.s�7ib�� μ�Eɾ{we�K��s�x�HaD��`�	�9�Aʇ���y1�X��t=p���W�f?����g�g/Q���ҙ�-�/7n��>a+�1r
8(��G�ԧfS[��|������n�@�X�3��1��;m���N��uc��c��	�\OC�6�bO�c����nzFפ�	cck.�Q��t��ۙ��y����f�{��ɷZ#8v�&'s�E�:@;m^���eス9�N�W�i֘����JD"����+C����!Y]�J^.N_�}ċ��p�m��/��ݺɩ�}0H$;��Rm�E�*B�)=tгgݝ�[�^g+\�{a�|x$���*7kS̴b=_*(��덢-�·���]w �n�� ��fa1T��l��x�`�wg����E���VH(�~M����mk5U8��9!�r��Cǉ$�n�Vj�V����/ ����>�u�0�t�KxZ*�	{�`~\8~���Kȴ	Z���A'Z�y��k0\lȶ�S�m5�`kHH@e����#�Ƌ���fh��u�l�/n7Lڛ��Q��hO��;YS��(��}�g	��n�ek	�}�q&���q�Rj��f��)�b3�ײ»��_N�-���CS�� H+ɩy�`��a~,S���Q���u��3��t���aFX�����r���������ŵpք�1�d�SU&�Ϗo>;��܈'ą;p �"���?]?j־�<9#�q��m1>ר	[x�A"��>�<Lm��"���Ma�+{�������HTv��wZN�:u7Z2.��ß5_���< ��H5^B��i�����+�_�w��9i�p++t�"����Y����MՔ�r 6��	'�3 A �s_�͚!*x$��� 	���J%���e���s�7]u��Gr
�I[ !�]�}vZ�,��l۰ �m��H$�<��v���b1=�� ���_w��%:@��_ߖk� ��j5N�ur�� ��9p 	 澼|
+#m䈝�P��u �AX����>��y��_|p�m'�1ۻ��~����dF]�]�;.�J2���9��y�8e&s��n=;���7�îU�v�t4����b�R���� �����{� N��Ot�l�*aL������[��z�������[�/�ǂn�Lwa�S(Gͻ�������=��e"�-��ǰO�*�`F�Q22A�FQ0"^2��&�-��
ͷַ�{e�s1�<H?O����v�&�
Ư8��Ld��y���-Ѯ�h5c�H�lAD��ܜ�h2AGJ��O�]�<�I[�V��/mWH\���I�ޜ2����ۮ�k���Zr�^<n�HU���Y9��}�{�$���� �A�v`6�1OEX�3a!�1I+v�����.��\ߦ�T, ��^���?{�A�����֫�����5o�>Y���'���;�I� S3��!{�o��wd�uԏ��9�>el@$��n</�\�fS�CF��.@���P����l>kwob�a_.l���0�C��r�+=A.����Z��ӳ���x�p���/s�?�����n��MB�(���}��q&��e1x5�].���(�x�
���u&m�]��'g�\�Ǎ��)%���)J������2�fm����]�l�T�TR��d`����w����t\�h4�/�O��؃��@�6���5��7C�c���߉�0.�$�x���*���9���xyަxw�>��2y��I!]\@�$Hl܁'�EC��珼�|$�	�h�B_�& U�|p�d�68^����Dy���p �Ԏ�$3�.���mk���dj���$��A'ą6�g�A>;�������{�70^ِc�Â�^"L�5yl9~'?'�C���_M��׀I+i������ /o�����ڐ�{�]�u���o�{ۯ9m���������ԥ���Y���'"�6`�8����,��ލ}:3����7����"�s����XF��K*���YS�:�5���b�4E]�ݰ[P�1nw]�l*Bk�g���C�����N˸���6$�c^�Ŧ�����ي)���=�LyO\�u�����%��b���ܼ�j�;%��ύ����Ѵ )%'
(4����c��.|��sxk�g��^�z՘��ݍWQ��l28�y2C��8q=��ܩi:v�l1�W�d�ʿz�Y�/�guqɪNY�t�b�t>x�Ymւ�\Bw�M�x�-B�(���gރ�J�l���$3b�wy�OZ�w��&���`@`�=�"�E��Q׉x�|j6�C�����I5���gn^Z��5�r]�<���Qh��GK���{�m5�N�8l�V[���A[�I'�u��n�8���wĒA<M(K��1��r���~�/@-Z�I-��q�F�5�eO�w���8�l���Ǌ�Yû��A �u�����5e
9�rbu��V��I'v#4�@À�SL�f�<��8ãtr�q�G+YT�&�Q��,e�5�v.��Xܤ���{~�#m&���o����I�5����%l"b�{"�@'�p�6�u6���*8}��¸��l�6�d��ՆB0$=�W;{hM8-H�g�P�}SO~��ۺ;�ȯWv�߆��9��0���u1��κۚ�RST��|j���n��Eyi��k�{5D�����#6�tn��d阰�٥���W~� ��<��k���ٕq#o�{��ݻ\*%��Y�[�7:�z��|���x��c�A7������1Z̚_'f�3���g�+�؎$�	�h�W�ޟd�����;o���-6�O�]lz%^>����s!�m��K3��HcN6ݍ46=��q�������+�0	]�)s��x�[�V��]N��mM��r��$�q"�y�@��l�u4쳂I*6��bgP�N哆D�u#}l�m7�Y�fbdč�`|�T	�q�V�郞5J&A��)kH�$~+�#E�U�S�O��ڜ��cm�cO�.߇��n9||||}}|v흺t�ӧN��:t���q�Fu��1�soc��mPq �^`�b�2��EåUs�l�ۄ�q{�D�� �����{=�;`ћ��h��nnٚ&h�z5�S��N(;�JY�ޞ��>���y��F+�m��������<�͙o����U/�L�|7(5u^�������{����v'�`O}|}���F�b� .��D9�3�8�{��=��ݧ���~!���I�{�h���(��1@������N�}��|��jRCńqo=k����
b�2�!�ק��W9���꽞^�{nK<��w�y!��bGwxgOb�ǝ�Ss�L3}k> E�F�h���;y����-��c�&/a�n���P��L�#w����qr}��'&E�z��r~�n{�,׈��i��D?F<�ш��L�{���1�-�q�z]FS��jOBֹy��v��a�:��`��<�jwm��{Vy�{sh:.���]`�偃k�%¦�G��F=��מ�,�wz���Yz�9m]�?	�K}��i/e˿�Dխ�7���ڼ_��8�������>] uS�}�d��K�b#�n���ȧ=�䇽�5�D߼�O/6��,g�j��Rs���[���|�G��~�ow^��=��_.������g�����o���"bǹX�y?z_b��/{g�/F[DK��z*ns���
���5NXWvw�{�xwE眩Ŵmg�燇{��;�Ěd�I��Lۚ'w���G�i�y��6إ �6��U#l������%MQ������m��������PI��a�Y��eT��
H�(%��I]L(��#RH�FnIJ�D奚.Iy�A�4��z��(���Y�ꛙ"Y)A��Y�E�hy���TXI���Y�k�yE�@���:Q4��UCB�BIgq�J�N^�V�0�b�^\�+�T�/m)�劚	%��yִaPUTTT�F͢�e�%��YA��G2$�U	<��&g7#G4��R0�t��*/s����ʜ���n����]"�����J���tF�E��v��t�]$#�5
�)r=�Y�*�4�<�ll�C�5¥q
��L�H���ܠԢS\����
������T)2��SȖ�so�)�7������|h�ۼ�]�\���g'a<��ԋ�����K93��x��pm�B"���� �Km��x�n�;ˑ�|#ű�|�����{��yW2�۠s
E�8xY؉�MsK�gN��Ny{M��*J���5EV=��i�����%)Lc�̥̉)]0q�}�p֓�NE��{~��E�X_5��z�f9�������O�%(�~��鞣�8	x�8��u�;�q)JV1�<O{�����fH[���iT���>c�!��	I
��5�wmbw���}��_^�|�T����N�w0G� =G(�L�o`O��"��D/s׾�'Q�t�q<���ϼ� �\A�\A�q�u��� .y����q�����o�$^u:Pn�V�F�%m�w-�5��s��u���	�el[�a�o�V+l�,���R�q�e=$�\A�pA�8׹�/L�!�ĆĎ��9��'� �-3;�<6t��>�А��q�2���8��yGD�#�W^V���e�7��XN��0��IG�]n���8�^�6����9w/R��!Ĝy�w����8��������9��1 >Dt��A��]�����	�"H�۝u��V9)u�X_8�t�p�������70��Bb0����<ϯ}�Z��������SIk�V��μ�|�!h���	q9�G�&~�}�j+AM,F�����؀g����c���xY������
�y���C�b��s�NlJR�	�����{p���U�����?�k�Ƭ��=�f�<�f�y�y�^R���M6nV�'��
m����!�1��F<�\�FC*��-SL�q��({�}�O���؈���1��"�u;�N�����	�v�{���y���`������I ��靱.Gv'���<��*＃�)@�=�� e`b ƽ�@�k	qs�����j,j��c�Eh%�ht<��հ[)s�78�1�J�*��n�YId���t�#��xk�<+����<a7�*�]��}�J蜲�Hb0��y�I��uP�ደV ��'r.�O�B�	;������|�~�k��x�q�l�I���D�^��&��N���<���3'��:�q!�1)B`��g�NlBbĦ8��r'2���r4��nھWp��Ȍ>�H��i�:y�����!)�J8��2���	q&!���g}/�ǽ�!9lG���Mg�3/0bN��x�����'0��8���fN��h�
(�[�� (c�5�mZ�R�1�1�#�{�7!	���Hb8�~dNa=lOdx���G>��|����F�q�%�3���G�޳�x�q��_P`�����|�[�vai�i�>����n�G�1�5
�6ys�̥	�{�a9lJP��=�yBn���)X���ϼ�#�C�d	���y���S�Q�b��8s3	�)�|vQ�ާ�v��5v�{���(�xOs�����0�����W3XȾ�qq�;d�ّ�!����/p���_YWz�N��\�q�dl����,���Z�U�q��u�u�Kjl㣶�8�ln��r�U�!�W�v���w���sq��ry�ㄵT#�.8�n]{{� ��ٗf�[;n6e1Ƴ�KE��f�F��\����˔Nu�P[�]X�M�.�r�a��u�:���6S&Ǝ�N�MOGb�"b,�x�4&�@t=�;�s��d�����^g��+�::쨕F�K"�� }��{HRZT"��<%Ƽ�P���ᤣ�$ �.#:�ܽ�)I�q&7�}�qRbC��ε\���q�Իg���^`�� ��@��F}�Y�:�s�ӹ��A:YTt�kiǅ}����q)�ﾵ��bY�Y͢!1��a��7�7q�!��8ÏW����D
�����>�k�1̔Y�K6�95�x]Z����u�{<��ʁ���E��I�����$�R�������1��G����CZ��r��|<���R���)�`���:��bs�=��֞�ER��wߓ��W�Dx�w#ʱڶ-�> �<�`�ǻ�/D�JR������=I�q8߾�0�Ϙ��w�|g�a�D�=e��#���C���&���{+`�rR��������y�ӯT�	w��q�9���L���߽{ȝB��'q�����q�F��}�xYk��՟xE�#��pbw��C�M�2s�6۠�W���_j6��9�@��.����D��x�mk���R�K�1'�}��x��#�0Dx/.�#�G����y\yH�p�N��w�JQ�{�C��9l^���o?g	F���E��;>IiP�4��k�~���Ё'n��7�����n�<�0�.��
z c@���^=
��`@��|yv��L{P�=�kɛ!��=�gz�/MY�-�^⮳��$C濾>�P`���8�㟎��&!Ę����w>�'����Ν��N
#z>Z������%�GMak<.7�w�t\K�/S��o�s��C�,�D#��2���o\/��l�=��p��<ϼ�%(:	q!ǽ�xYx^ï
��~�UYe@�e�clz�|�� ƽ��[<)G��,�38�u)JR{���.�O[�)�J�~�NK�ێ%(Ϟ{����:���:�J�&$���#�J;E����wH�!�$��J�<a7�0�R��g^y��^����o=��~.dԜ7puϜ����LC�LK�q�u���. 0�$0�#�}�"s#չ-��#d�$��9���?��Wkƞ<Wa
N�W�8��gF�bk�V�Y��ܕ��V9)}ְ�����y��u�
)1�10%��n`+-��a��#;�܉�u!�{�rW��u��,q߼���R��\A�q�����b�F|"ϝ򾌃����,F���糳�_</�����]�㣚}`a����G�w�O$�E�����q��{�����	��Q�_����6ó9f��*����#<#j�.��샇u#���y 18 1\G{�^�^��.%)I�޼������Z�tp����нW=�ݾҁ��{D��yo�Zi�����/#��ߟ?��~����z9e�D3[=�Nz������<f���>�$W����q8߻�e)JR�u��6�-��h�"�t�5���a��{��A�w�Rjs+NbIy#]�焐I ��nD�I%�|��G��+-�*($��蘓���X�+��]݄��ҊI%6sdO��a���/�P��Iy7vH�(�A�_�|������Dd�{����|�\�cu��b��	�\{���FN�l�J(��TAA��[]]�W|�2zć6���vdI�%7s��O��1�4�&�h�RH&�������s�v,�2)3��]��5̲I{у&����m/��	G��|�ѹ�&R^	0�[t)Iz|�}�3�������z��oz�������JJ�.$̰fA'�n�d�^	 ��5>݌��	�ȗ����i$u�T���,s�c�� �[ړ��S-V�߯�ͤ��35�LI���I �o��$JK��Ǐ��`����N'�pɢ"�y�j���s�R��������rzz���*��]���(���^s%�ayc��p+�.E9y�1"M�5i����bO�}"E&��/��^����K�_֢p�� } �����t�]��	o*]ϲ���̼���B>�7�8��x�LN��=&���4��:��}��]��{M�c��\�p���$@!Z>�}�IeTT��?o�L�LO���I��!I=��H\ڻ��魠��$H�IS����¤��H�����˧�)?sG�/$}�9?{XF�R�l؈�(�f�v^��K�-�h�PH
��m�:6T�����䐫����1d�I��]���y��Iy#W�H�O�D^��Mu��_�I&�ǃ)N����r���������g�I�3k��ּǢ��os�Iwv�)k�Z'�y��fL����}�A������v�4�ݜ�p�Q��M BA$��2}k9'�($���I���H%٭ B$����H����=�v���B�x��j�2v_��L�0���Q��x'��тR̪��Ӧ���8��ӡ�b�U���Q!4�³��ܛ�*�����rK*�fg���|��쪱�-N�R&�v���4��<�oHs��up��w���q�.3��5�z��Y�Y.c��vq�ݰ����h�6|�=�F�g�q��g8U{f�7]����7���c�;���nݢ�t�uq袒�w�A]On��:�\ TYe�m�ik�b���s��q��>v@v7�v��\�=W 6����,�Xx7;v��[\ןg!=ur�uG`�6g��h�V����&q�H7�wߠ�Z���{�L�?bF��Hﵢ	$���dL��	.ޗ��ug�~�뷽� �! 	��	�ȣ��L�Y�;&��$���$�M;}�dK�d�lL�JI-�h��I��"|%��u���Y�]��>�0����]w(�!����4BQ�f�]q �	/$|�\Aڼn�˹��  y&	os90As�șKC�}��N��]�ٖ��dLlZ��[�o2=��=	y$��>��PIs�����/{��C�T$��BE�����;�AӼ����)$�ds� T_!a6��R=2�I���t��Ƀ$c�L�#�MM�0�h��ؘxO#
L��f�\kf�/Q�5�j2�vݔ��yvf2;aw�v�o>?VX�yoؓg�8Y�?"��L������&R>/����V�����I5��Aqv8?<i�R�Rv�v���D�����u�)��׎�`���V4�v�������}�W~ǐ?�/����˵9&m�<}Ӆ~����]�Y����f��g��I`������Kd5�J���$6;�I2���FD��f	��P�b������g5�z�'��	�h��%��(��Na>��p
I�	�mQ�!����X��+���:Q��d�I'}M�bš:g.�+OZ��ӣ	�3$�I�v&�2�'bL��H����9")�b���'XC�B���K�6DYi�fI�&u3��-�zY��I�h�}{�/B8�⹭��$�k$L�J܎�2$��h�����f�?�{�����+y��\;G�9K��;�6����W�焤��2*��
�y�_@����rY�q �	$�#^'��bI;��>Hݼ69OD�f�~�(��c^���o��u�A� ���>śĞ�nq���Ϲ؆�'��<��^2H�f>^܎�2�	 �w4E$��M8�2��&:��I]�x�h���տ�����H ����	$�#����m�R�mh&.������+$�$�E}g�o�G��s�j_��U;�/!t�ۻ��K��L}�	8v��)��7�1ɛ��7�j#��Q()Y���Y5᎞�ﶚ$�I%i}�4�Џ���l�`Rb��;&�$�[ M�Q�q4ea���<�O�̋�[��	��d���M�m��'��m�9ok�ג��SJCޣn\�q ����\DO�G��#�W�2I&R�֏B)�� A&�mD���bx��.�(򜝻0���ǡM�q����n:�km�) Q�Ѱ\^�݂��F┛���vi��H���e���;$L���nH��]_}�=I1$����̚�������D
c�vE��H�{�;t��~Su�U�E�d4`�n]�&QA#孆ļ��e{Y�����*�
Q��'9ĺw��(�`��7ϒ���q��d��X�ž h$��=��_�%��+Z�_��WJ[-VZ]iOg>4�-��e�D�Y:�����y��D��I���C����N�N�Ab��Y�ZK�����Cޞ黮�{O���z<]�R��ٳ"�Y�9R�]OE��:��ʦ��:��.������q��~$JPJ��I%����?Ӈ��g	�5��'{�)/��ǉ	 ��b�pY>��Mr�	$���2�(7�WD�O����m����0H&��x�vvb���z��3筽=�����池lP�l��n�P<�˵�ж�ە��3��x̊H���gI=H��!�d$|ɳ��y����[8�Ɓ�䒷��>�����3$�:�����g� ���U�A�,��l$�K��r&|�30힉2|��d^�kk5cr{��,Ȟ��
Ub j�No;�Β3[���@ d���vm=�l}	��@$���"@E[3f�D�	N���i���f��������t�I����h
@7�K���&BH$�[���.R"�넹>Y�I�zD�Q�Xs�t�Rkw�?��I w��!J���YN��Đ��^��V�{v$�I$M{�99��맷���N�_^�:t�۷nݻv����ӧO��s�\���]kA�3�_�e�|z,�Yw�j������]O�'�����(�t�N��_t��g��<=��hNL���~�8�n�~A��-���r俜�Q�����d�<�M8��w���vU�.�B������k�h��ǬG�׫���{���{k�\����#��r���]\y)��˧}���r��}�e]:�{�֜�w��54_jj�:D�eV&���k�ߡ�o�{��|~މ�(=�A�=�w�[�{���p�ł[��!9fz��4t���R�l�b��o�_g���[��!��9����
Δ��SF�O�\���w��_�K}�s�rM�!��}�R��ּ�H���~���g5A�6L.̹�?�;�����y�|<����O�f��g��e�x��t3{�.���ؽ��6�_"w =��mVw\�(̽�z��y�)�uc���*�N2��6EyU��/N!U��W��ݺy��n�(���[ѣ��g�g�n�Տ�V�8=���7��뾩n��=�1�=5hW�ѻ�&YF���q�y]��^�i{W�2ukf�q�;��p�=�0�	~�>�MgY�<�\���S;����us��76�������~��'�4�ெ�G=2g`��".�Lcu�B4~�(8aT+1��vq�U"�[7���-`�9����fڽ�L��u�i��?���vF��-Fb�~���?9�GY�=���vw���a���\�o�F�N�9�A����<=���p%=��[������㊞���яf+֌��}��|���w�tg��#���#8K���o�YI"PĎy,��m��E�CE�TCy(x_ ��;*��C�?�����Ơ�0��ɖ�Om�J�*Y!Vz���XOP{�{*(�>O��yP�y0�=�l;�$(�y!�Cq�{�x��p�vG�g��l+!v��yqr�����<�0�\>�u=L�n0��{w�ϮwhtKT��B�y�t\`�S(�c8�ݬ>{��np3�z^�WWt ���t���fH�	].�����>���d�DDh{ѫ�D�]�¬��|���$ݭB9�Ԁ��P����I�EJH$S̆
��G���/�OD*�n��uz�*Nүa�P����Y^�2��EE��9�u yķ�|�܂���":�D%������q���.઀<���e�y}��ܔ�L��w��$8�D��cA=�G���{Q˞ɓW�)��ɞG����\���@�Bm�h�{i}��oA�r!�
lC�%Oz�{{w�'���2����2K�.Lɑ�[B
fx+n�܉A3Tg�:���1,LI"����A�dϞ�B�T/(��I�O�\�#�'^eP�<��5/�*����dQ���ˠ�^�ύ��]i�<��{��Y\���"<d��fL��'�U_A'xd<ʯ��w�z��~ݶ7",R��c��G:8���`�nw����fأ\F�R��Zz6����;Z��x�mї�n{n���n�ci��l����l'[�냤�&S�#���)P�m�=J>$in,�1Z�=v;F-�8�R����������V�Q��o��s=y�[pb��ͫ������l�;yy���Y自Y:.��uHC43�����6N��K�r����u<�iJ1^��v����N;qR��L�1Öl����xu��]�-b���[��N����^*x}�p��e�Ŵl5ݺ��Vc.5��BL5Ԏ��@�e�v��m�W>����ۻf��X+]7F=�tod�2��.�n=�E�{.���Ý뭦��v����s<������z�5r5+�C���nst�n�<��Lq���d\e*붍��5�I�0cam�"�J������������]hk���v��魵Î��#t]�<���&ƞ�I�j���D���mМ���gn8�D9��A�M�T<lO[��m�����d;rv��q�)�F؎��l&c�,�a�m���;89,$�۞���]@�[���L�_n�θ�K�؎hu4FV( D����N#rk�Ǉ'm��g���W�|*<��qq8vl���v���$����V{=�����`��l\]��yU��	�m˳�m��a��[ݏZ�;�L�d3<W�v�N�x��75�U]+��u�k�6�-c@@Xy2�
4�G	��2�M��1��g��d���u�lf��n�yU�v�7<�p�W��^yl�h������mI�xݪ��10�l�l���4q�tD۶x�Jh5�f�n�<=>��r�pg�c�m^��u��qGg���ƹ��X^zd���v���V���plpu�ܤa<�)�Kv�ۜ%��m�ֆ�Ԏn
�M��۶�Y觶�M5��/��w�wr���1% Ҫ�\1��=pg8�I��[(eG����mły�Ϭ����x��pM��N㋃����X�<��Ev�����K����i��Y�ӻr��"��.��z����3[{��Vf.:�?�=�ю�sp��5��`{v����Z��9��*�0����OM��L2�Nx|tb��ܜln��D����m�<z�#������켢�6�Bx3ѫ�^�����u�sĢj�L��%��V��������3��W�Q0���I,�ǌ�U�I.�h$�~��-A�ZX.��u73�R	'��ߥ Y;��A�Ra%U%�Z=	y#��PzV�?�RH%�aӏe#�R	osG�&�y�:��mg<M'���;=���H�@8S7��߹�H	z�$��y��0c��|���	e�ֈ&���͉2A%��v�G�ʦ�ӹ��N���� u�r�:���`�+���H�W��k $�As�φ&6�uuU���'d�j�2Jj3X&wvw!�;�Is�D$!�������77B�Ռ��#�L�#�
^J�Ʉ�\��'Ҁ��7�uk6,LNYG����G��p��:瑝n�����-F�m��7η��Jv�N��T*�W8��a\��Jc�W��<�I$���	��7�;dL�}������[z$wX��2�	/%���l�:�$��'d�Tw� �$�G��n��XG��1�8��mm���;A�������{"U�}���%>�n�w W&�&-+�}�,��
u��>�6�>� 4�� %
�J(�)�y��͗�m��Y���K3#��@�L����Ix���z'M �Ɔ�ֲ��	h�R��3$����@2�D�s�v'h�v�\q�%f`	��G�+�%��"e*vu�&H�(&uUA5����і.ꆅ�A#�-|%�$�>Et^șI$��"I�x����fWƔ�I�v�)���@h)U�Ӽ�=oQ`�?0f�7�	�};Z�����o�|��޼L���%���/R<�o)��;ŏ�O�X�7H��q\,j�5VY�q��%΃��+k%���ETo��T-�(�<��:n��I&�w:ORH��k�D�O���b Xy�@�t�5�I$�����jkѧWKerZ]?S�R�K�9�ghcl�N�c��	 ��̑$�������ϒ^H��^�L���C��Z܄����(,OIn�����I��x�$��32��������?37A�6��$��1��\�qV�̸��@��Nnfn�*��{K!l@W��r��	��7&CU�Q�kYd��A�< ���JU
H��iT)�T���
j�����>k��8���/Z�bI����=I1�kC�^��$���~����u1�F1����$�깉�W�C�$�>I�������i��t�f�U|���6��Q`AL�UPO{�3,�2I#V�:>vqkY��0k0�UUP!{��^I��>Iy$�ֈG�h�L�Ƭ����!��BJ����Q�Ŏ+n��akć��y�9�A�E�=�����V"��w��ȱ�)$���Ą�&�/-�h����W��&f�fo^��q"_̙$*/�L��k��i�*O��I�w+2H�;��窆E�˪��潋2�I$=�I��H����y0d��Y��So=t��9����\��X++���X�3�Z�&�R;�h��3}�WL�gL=+R%��V�I���J<����*��8y���8weU~I�� pխ�]�%\�S�`ʢu���>I$�n�BI#�� ���)a���y/�1�\�c��EXHG��f8���o����C�����/�>�I�����w��nC��7��<�2�A�O9����뿅�F���P��R��%
 iR` �Y�JV�I���
JQ)I�ˏ����_��ٌs�X��t������%���*I'�{Ξ�=ߧO#��w�I����)/"�Wz��������%�m�y��{KQ^ր�a�/C��u���;=����-���svn�mrՀL��c�f(�(u����sɔ%�^��I$��dL�@�/TN��!-}w�Qs�{�@=�HN����M3��-�!*踐e�e��!�^'B1�z1"W�+�h��H����D��a48e�k��9���>�KLQR|��O�YH$�k�Ip���i뢡�l�D���4B(�I��{ƀ�h�4���p�2,��@+~��9�m���I#�-�C�7W@�H���O���g^�E���{䀶����) �,OIn�ķ��$q� �AG����	/*�h���̐O}�$J)$>�J������܌���kӵs��C�.iUE\�Fg%��z�/��z�Q+.:<���ě'�uޙ̟a>��
�}\/==˸�-g�y1՝Z�jiŗ�B'3O���_���ZP)iF�B��	�R��)d�Q�i@�)(i���P��~�W�׵�lI����M��+=��V��^��7FS]�bhMO�]�v3[�Ź���W)kp�w�p;/XS�G0sѲ�w3��!ڎj��S�64�ysm�^$��<���f�8Ǝ_-�7n��t����\���hwO9��&�[��k�-`�_'S�Cdx�����cy7��g]��q<vrR��wI��1���]G<��9D���k��w=h�c��盍�k ��wϵ�����WsI{˜��D]��|d�C���|�Q��WC�L�����H&�%/P��4;�b�Y�U%�~��%䀦c�m���g�d5�I��%%�>�I��	U�u\����y9݆�VdO����(X��R}��I��	k��HI$	 d��8��1��Lr��/�ۡ$�M��&QI,}�2E��y���B�T�\�$�csK�+zfZ�m� A4C��$ϒI�����5�Qh��� ��M��$My�y�/U^
�c��|�M�֤�H��~�ϡE�cX���2�37�����L�$��=�&R�7��������,}�2����Z�jG��d�ì˕ˑ�:1I$xM����*m��ݔѪ��HV���}���-n�P0����2��@-|ǉH���� $����y��Ӗ�Ģ����(���}����Wsw%��s"�����>�O| ���0�����W���B��.w���W�085Oyn���ݦ�n��������軹M[[y�j��|�u�*��R��"PbDtCۉ���1��H��e�) �J(�`T�@Z@J& Y$ `�=���z1��;��qф�@& %�s�Kޤ���\4�߰_�|��z�9vf.PA�UPM��2�$��@�J	kC��K��cǒ�����jjH���O{�9��t�*��yi�U�0��K�T��L�8@%n�"}�d�AgkD$JM��ᱏ	��E]�	!��r��Uf�wNY���P�u����y��{މO�j�*�ˢj�����W��ޖ,I�fs�H�=*��z﮽���Q��5ێXYhbG_E����&�(,uٱ���D�&Q���o�=��pV+gn�Σf]$�^�}�"H�?vP�	g�:�_woo���X�Iy.�g1���fH�f�ݙ��$�e���� Ԏ��[PĐ	�W��	��L�#����Hܹ�/y�I(�8�hgL�X������$�U��Iy#�����n4'~=�.Y��K9��s
�A7��1��N�bL{Eŗ�;ڻ�x�U��t�<c�V�t6�÷��7��nl�wԽ����Od` �B`� ��&AY���B�
&
P�T	ǻ׼���p�\W���I&�nD�R�o��vf.PA�]�m]r�e�����!^��	�h����)$�{"g�$�a���� ��CXvWi�I�G����:V"�q%�DX3�K���R���/&g/����� A�
g�!$�M9�'ҊH��$}7�];����4E��	�&�a�3�h,����^�a��>]�YGl"u�c\�8�A�`'Wޓ��q�$�K�w:PI$�������]t�ͼ�d�u��)$�ﴵ��q���Ub��]}<(��D�9>]��i��j(y&��),�3��}�jI$}��n��F8�k�>jG���wЫ4�,K6�VIf̀0�
��䮈�K��j��5"��I$��dL��E�[�{ΌB8�LL����]�b�޿��	�1T^D�)_��!���ғ�&�]|�����繎��N��*���@�dQ�ǻ98��V������
�e�Xtc��b��s�GW���1�;p{��d�ݖ��@}�
Q����R	�	�Xf(�A%���c<��GGX��`�zy˳1r���WQ��^Q�_f���k�0��t�����2I��`���@%���|�nzߞfp=S�W�wlp~;�[ύ�W#�n������d:��0<�{pƫ���U�!P����H`�"�2��%ٕ'�P�b]/�G{�� �P��u%�d�����).�L���������:��oja����;#ƺՈ��*e���2�K�O���)��	 �v4B$�u����#�-�lA��a�s*�X�.��	�kX$ĉI7=�<�$����3}��'����%�͖��@.n��vH1��Qb�Y�vt�w�;�@	`��g�=�i��	d)�c) ���1�To�@g����w�L��C���mWn��?Z��>��h��U�\$@$�W����jN&7��ZI^�Դ��G���D"J6�H�J ��})ss�է�����<]�<�L��z�:��\oh������X_���n�j-?F�K�@�x���8�Rc��mG���&���dǁ0a�c��/�@�)@I($��L��*4�$"�<{����]x;; g���/GY�*�\�Y:εm�Gev��v�;qq�����L=r�&z��lk�A�t�c8�<q��[`^���Qb����W�8�ɺ�ԝ��E[X�kdv���]l�<f��U��{�/;�>�0�t�o;qyاt`#1�b�bk�2�W�Nr�7a�;q;Z�{�Jct�m��=�W��R�����`3z��9%.q�:s��\�޹�Dw`�"�Em�	�����]ի��3: �J��:^I�f���H����I򧽮��ȁ:�7�Cm�Ғ)Ӽ�O)���C B�SCz�Z]q�Fܭ�*.��Ӫ��D���� $�I�:D�S��e;���(��L���qY�z���:ϗϰ�me(|�'���މ2JK9@��*�D$ד�My$���B(�M��$JC��r�E�ڌ�~��|��g�f��.��JR� �K�&��) �]�,�������e0	 ����CW�FV�Ř���隨�m�j���K%nD�E�]�����fa�֢<�$�n�� J)%��������˔��d��c��*�%�,%a����mǔ�m�{:q��k�.�Y����\q��G�'edT�����̒KϷ�%�O�I$���2��ƪk���c�;L��PI�]>�H
K�9vftA�UPM��X���y��t���Ta��������O�+��9����tM���?�~m�	�2j��ڧ�M���H&m��Gr�f�Y�3DC��)����9缜c�>$P�Q�FIJ�d�	� �Pߝ���BA$^i�2A%�7}-),I���7�{8�!�>b�wx�R�Qwzr���I%г�����1����Tc�F�-��(&�ɿ�	 :[�n��;Ͻ�����i6�O�7������Ami�I��<���1-�ܖ��I%��y���c;bs���䉕;s��ڬV;J����g��$�H��h� �%k�YtZK�;�$�q��18�����a�,��Y1m��4 o!L�੷>5���z��&��;�֪qQ���V���=��]������H�t�ܓ���tI"�H.�h����u����Օs�@ �7���'$C�?؃A�M�T�&�h���;�`�[StƙI��דu#qI�z�ˎI;�w�_��h
S�'FγX�Z�˳3��ꪂk]s���^H��9��J����=~�O������~�_���ӧN�:t�ӧ�N�ӷn�\��Lv�8��Z'vI�r�<��	HzMلD�s�;�Jc�ǈ�&� q�ˋ��|w<y�w*y���V���m���]�,=�g�o����N��[�r]�н[̞�٥eNU1���*�(ͽ�]����k��w�۞�/�e�'.��\@����u�t�*��̪���s`�f�ZXە���q!����� �:��3�Y�T.��Fg0�*M�u[�!�v11��Ob,z�ǝ<�o�睳�?q:|`��e۩a�[�Er��yw@V�>ų���tںw�j����8��[ 	���{�wW��j?e�U�vԐ=��u4U����8���K᧞��wCMN�R��A�vrt6��;P2r%��L�]�*,g�$��ЏN�٪s��B��)-��=�PHB�W�������@Qs�Û��y�=�<��oN��%��Wl)�Pt��������o��S�w�ɲz�e���=�r
`����?HG8�!�C�1ڱg(�N�������v{U�n����ߟx3��>��r�c���Gk�嚬���g��W��s.����ա�0�y�9���x����\M��u�uS9�p[�!��R���S�Ƿ;]�,�Uk�e�q=�q�r֩W{q���ܻ���bg�6��5W2o�Γ�=�}q�w��{��;��qQi����k�ׂ�iÏJ�<���b��ʉr���Q�����#�XJ����o'�;��c����<WX<���5�>s���{��"7��}'��QW?�����k��D��������^��yE
��Op�tʃ�=3��_%��GE���e{V�BsbI��d��DS=�*{K�R�Je!|2�ٮZ0�Uyb�D�$א�@�N���9!D�[����E��S�Њ��}X�QH������$*� �\� �
,��ș0���r(��{�}F�E���:������P�������>�1��4u**�<��
����[U�HC<�+� ���(����'i�{�reCED��UQ�Dw#\L=�2�y�bT���Tu
/g�U6�]\������I
�.�1�2򼆸�'9�Yx���D��h!PfDB��U{k�)���*�/���K�Or=r�T�O�J���[eH�Z*�E���ȋ��(�E:��w����DU}�2,��҂d�UO�8L<�lgE�J�
)����C��8~4ʇ(��)J%%*�� R��H�"���	HP*8x�U"�}�`ɝ}�����f ��$Ri߷��C
Uj`lܛ�w�~�%�)]m'/��I\��� �+�3!$-�����n4���eCu��� <�����C%f����ws�1$��)9�όؙ���t�kOKHH��ƈEy$m�"V�<j��A̐�$x�7l�v��#0$���kpSK���L�B\g�������-O�c�j�X�/�6L�U�H���!/$�H��N��g�wN�RĒOf6Ho�Ge�阳������N�� A_���i���"��H$��!$Z<�Ͳ&RE �{O�Cf�OW5���J��;�P�'����$��'�x)��Km����#X��%����I&���J�W2�,�΂;���uA�7���e�H$b���"Y�:D�I �ͯ�||}�|h��⧹=n�x��xrsCx5�0ޝv㥼=��r>xgU�y��l%�H�n������S��7	�`�{��䳣�;��+� �
*(R	J�*��J(�/8�~R7��ѭ�7��Җ��7�>�w��I�g�.����։�Ē��Iy$��$L�
Iy���\��]pӻ-<	.�>M��t�E�禞9�T�3��8;%��ݕi�v;V��s��L�`�Jέ�o�i��H$��+�O��-!!�<_--eo�*�h�~H��?nH�+}�c���2�3��M��X�I��f�'l�7��غ��Iy��D�M�f>�-)#�c�x�/�w>��sD���s�h��"R�����GLH2��I�_D��($i��G=\��}@�Kv�	�RI�����%��%�X��i+�������j]o?I1&�&$�I�SwKHH�f����?h~�Q[f^��$��̈3����&gA�U+u]2 ��̎t3��i	��-��-�	F�H�	$�kv�H�f	���������ښa���#,�ĺ/1K�#7^�0��tF�<׳|���)Mƣ��f��'[���O��uj7m �s��P���ҏ��Q�C��ws���D"��x�S��$���q�$ �� ��E(��(;�;�x���_1�c�čf�y�q�f쏺��à.9�1�Gm�uy+���n�4wF���2Qۈm������ΐ���]���,�A�k2�n���e��H��/p5<�u��7L��76n.�0mpp��\��K�]���ۍ����y���:���&�Jqm��O�иS�G��)���A�kV�ł^�y�v鎓X��@.��=����&�/{�{�����v�f�Uv,�;4��q��Z����~u�qU ����$�9%%䚗lHt���K˻�!,�ܦ� �7MȐ%�ɂH漖�f���L�`�J�-|�=��������_z�o$e�^ƈRKy7��2�|�	$���'̀a,͛��=
Z�L��J=�c���2�3Ǟ�>���I$���rI;} ���2�.�I&�>I���@
��ً�����4��tb�W���J��	�"C�"%ye�D$N����,�s��q�
I����ԓ/e}����$�gYͤKv\I��X���Y�@LK�SPHRYz�+�`��o4?t�/���9�Wە�"�+� llJ
X(/��ўͲtu���ݜ�D��Q@R�(|�վp��\�p�WL�I$��֏BI ���%z|�,��3e��c`~i�c��D��q�� ���A�'r��wx���95�+�/�?���S�t�B1�c�Le[dcR�H�U/�i��1t�GxS���*GN���0��3���m��9� ���{>�s�s���'ʿ	�����Aa�x���6
H�O��A��fS3*��ǚIa6�KM��)J#�]u�y�?q��c�|�)!?�t��I���h���r�1��W����C��ʈ V2V}��ؐ��s�5y�y(Έ�ey$S�NJ.WuQP��Z�I ��4B+�/&��+hm���s)b(�[>���nϾRO�R����#@���H�s9����$�nDכ�۲�)��M�����c� 5rs��y���IK(+{�$�}��=I"R]Y� :����h�a���x�@$M{�&QI ����z�.�r�2�~_��[�q�џ'�9n5��iٷ�cN�n�K����H���W�����f�)�rg2bI#v\HRH�swKO����m&g60]�J��Q�E �	�nD��`��˝3��Bb��:��t�@���nh��jX!J�]􉔒H66��1�Nl�n��͏k>��v{2_6�]�]T��P�o3]����H[�lHt_ɼ����؞׭��WoW��<O7�`#S���k��zB&�v��h4�L�	{;T�Rzh���f��g��rԯ$��*3�]ڨN��j�%��b��-G�x�xb�o�����*���KZ�I1}}�U��k�f.]1y@-��&�8U=��Hk�'�6�\єI ����I��ӐE�2Zu{r<�̒��>��1[K�`ɊL��!/76�K��G��<!^�I�fu�!$!�L���y��!�g����KzYy�
���!.C�K��0�p]]ɱ�����˦��uֹh�r5Y!X���k�����i)e�����gI�)"��o���m<�$�#���BI�8=��f1�Kχ��NbI}{�V��Ϫ�u��h[�|}%=b%�`�V��F�ۚ���7��OKzR%u��sO�������\`�(�9��wgw@���	�Y
�X�D��h��7��ܭ��I��h��=<*�)$�ZBK�$�����$��w��]��w{rs�����}��IL�Ȑ��o1G�%{��	$����=^�Rkf�"DS�bd!�i����L�&ڻ�ލ�͇r�5����ڽ�ݛ����5���y��B_u+��d��%���r�^�=��'h���{��o_���دa��L�ު��T�V|�����d�Io�����V�n�`\5L� H	]�I/&��oD�޶�sB� �(��$o�;�ڵ�G�o��y��eۮ͎�V
많&di������v�X��KK�K��kN�%�g4H�M��"BB�Z��TOnWO�i�i�H$�U|�΢�_��3�gwj�
<��@�-t�3�9�-�&����y��L����I.�h��@ �z�L����w����)�%�vX��b��h[��'�ܬ�$��Ξ��)��x��v��H$�]��!I��D�R�����\�������t��k�l�O��$k9�А	$�{�D��I76��:���uqX9Э�-�Mvљ1�����+*fғ��󧨛̊ŝ=U����.�d�]�� $��n�>�IM��->@#�����2*j,~/Ω��������Z��������xd�\�<�����yC���h��Fv3O�B���{��� Dl۸����'P�d,��8�Y�6�^uհ�9r�vWv�eH��>Z[s�8���p���.��2���;C���@�p�:v����7�[�<y�4�\�z݌OX�Ǟj��O6z)�/b�n���]�kZ��y�X}zh�;=N㓌6ݼ��d��l��X�ɉ�3-�i�P��X�<ۍ��3U�;c����[v,�y���v�[n�`���'3���Y6�_=�7�138+��ky"׊gd�kj���v7]h,�k���$%eu��ߢȶ���3>G@�e%���E��s�ccp���J{=��n��m��ɥ�LRfv�M�:gΗ�MSfk`a�q�盄G��#�S�����2A����$���)AZ���s�fD@��(J�����Ǧ䗓�ΰI$Rw2 ĺ����1%�w\g�R($��:ZT��h���W����ٵ!�^o�S�T�,ҹ�N�͏%$@76��"4���ӛ�K�N)�$�ʼ�2��9�N': 1�+V��Nfgz�S���M�9��I�8i��U>�f�R$�g���$&BIsw(���:��Q���Di�d��C0�j�G]T��o&��U��T�Ü���֤u�X������l�,*���l\I�y�����C�I+k��1�jە�%&���@�J)$�ײ��4��w�U �*W���}9�$xx��11�K��:��Q��m��mPd^>�,�+6'���w�2�)`*Yz��W<��[�pR�-���V���n�$�������_nl|ex+�3$#:ZR���c�~Q�D�/6�� ���~���ԋ��N[���Iiu�{3�h1dĵZ�Q	��v�X,���Iԓ�oKk<L9'o�3�ɵ�_�P�(J��wދ�=��2�`�eBK�(�5 Q���JƌPk�Y$��9���o�Z]Vo�����',G��؁�M%U�){��	$��udO�;��z��'f^�Ơ����%��$�`�On4D���L�Z�T�ǽ��SR�,�R�%8z��܆��+����td〉�Z�����	A��f����J�������D�6����D��&��)gV.����k��nS�KHI ��N{�+3�6݌,(�&��{;�q��8��u��.S�Jj1�$�
��#�$@D&��%O��K�%)�(Mo=��_���H�\f���9��瘨����%�����A��G<덣���R���Ϻ'4��i��î)�:nA�@��=�.Z�����n����m�dP�#-�#[v�aӼW�Y�U�d��?�~x�|^I���"�I7�t�R�[�Z�݃��������s#��	Z�I����L��)���Q4��iLm��'�g:1��N�J�u���Ξ��K�^f6m�=s��I�=m��S���"���m��R�.��>�ܯ<�R,pp�ؘ,n|��������C ��k���)�+Y�m_~m�<~����-��R^���H�1I��Xz�L@m��RP.�v�Ά���I�Ʉ�l��"Vݛ�ݘ;�34��^�L��̈́[��9���Hg��$�dI2�]��Gl�*o30E`�]����w�w�$�����N��n��II��q �)&�n���32�wTN�����Iy"��e䗛u�T���=��;�H;�A�]��m�alٌ�U�i$�#�O�'�$m��D�!-�o�#����j[���k��v��2�z|���!�ͫ�Z�$��W����ojb����e3��;���*���F�RaѼqI��/	�<��v �S0����?����	R��9�V�N���L��I��I$����^S2�ͼل�>@�Iy$�o��&|��3�u�^��Y�$�F��n6{VG�i�fI����w�7b�4�-[c[8Vumo�TЖ��ސ7��=E3�`�=�a�D��g�%�"Wo
��f|�<��dA3���͍�!%��A����Uq�[ww%�(�w�n/sZ��i=t��"#=�Q�)%����TAw��&�g$�쌦�"�f�5˼��K�wL���	���s0&�k�e"Of�zI$;1X�'�I�D�I�n��j%qj�%'��f4E����!iF���������;�����j=�"m�e�$��g$����S|�cB���u�~d�9�T��ς�N��P{it[@��H�x��ؐf2�A�ږ���%Ͱ�^�e䷱�$�w@�Y�����v���������.�:t�˧N�:yt珳����g6�F��&��I��IM!��;}穄}�;�O�/9�xh��]���=����]gpi{6x�����ozcDp��}_M�Q�ǒ#��!�q%3���Ԍ:��<]=<=�����YX-Ƀ�Y���t�������ְ��ug�Y��a��k8v�,^Ξ/پ{7���n�|��Dޙ;8����8	�l���$~��L�{��2�x������\� �����n����:S��.�G�3�LC~��H����W�rG�/^�x�z5( _e �<uh�Tɚ�]���[c�_I��=�鍟Q��+[�jÞ���l�'�p#��W��*��̄���ro���.����,�c�2��H :%���h��bd��#�.�]���t>����{��M��;W�Z�����Jg!��V�(}7F/]כ�zy׉{��(�O7z��iv??o��>���}��f�掻*ۆQ�g���J����A�e�}g����z���{���5�;~�#��7�	����+�Py��S�}�����<�݀]ҍ
�Ng47ԩ�OzO�������=ץ�|yo�[���jݾ��A�cF(0a�>i�q�~�k��YO�a'ѽ�v�����b'���;"����Q��n�9)P�����s�y�w,�Z9��xw=����]{7��:g\�+p��V�p�6n
, E�>�ُ�� B�F����w�=ϭ���k��y�^=]r_`�g�{ޏ ����IÊ�ݒ8�)8i�g�x�A���W���<���D�'
~ܷ����� |�n)�������7|'����<7n�T6c@����0 ԱE�3�����
)�T�^�ZQDT	���V��Y�h�x�x3.!{�oއ��uP>Q��*𼙎��	��k�EN�}6�an��u����}l^A�E�N���I2EQ�J	hH�{yI'���+�	�:9�)��Ha^Y*9F�!W������j��aV�d����n��1�Y<�@��'D@��e�痗�xS㇌�<z�Ćz�2�a�Z�`J���dj����Odez�Z�Y�z�yU*(�HQU�d��=�]�+�r�� /3I"�(pH�̈��rR�$ ��]��/L��I����UQ3ȓ�(����'i�I	�Y�k�	>3ƢIP�I�xQd�K�/
�(x׻C�OU2Q\�bain��2O/(�J�V�b$HnQy	�N}+�
�����"*
)2�K3�$5[��u����a�{�K���m�V���g)�mgnܽ���wh�^�pޔ�ۗ���tL�]J��݁�彏;#:}�z���Æ�xۮqÊ��ĦB�ی�T�R�b!�[�Ӻ�,P����v������\_���|{<{��ݘ��&8�vw����u�gw[nn2��h�-��ŗ��f8��/S��G���<�a��dخ.6�Ѻ��ˎ�s�P]���ޘz-�/ݳ�T�D���,�/���$u�<h���s�b8�&�]r��Su�>1��牮��6\F�֞�$�M͂�v���u<}Ʈ�8���՚֎N��^��I��W;`�Gg�-�a)�n.0�3z����o�\�.�ݱq6�\�Mn�v��;pe��!�Q�.6z�>�8�ڤFm<n̳��Z�:����7R�j8���;�Y�(5ٚ������J����ƛ����ٞ��u����̎�i̫���pː~�7�z�ӑu��[pEuۄ7J����1��6�1ϒH6-�Յ<��)��3�FmнP�r��N������X��\c�{s$�������Q�&ػ;�����@��RvЦ7f��]ru;�T�=�\��,�ַ8��O¯�y�NK]q�<�Mb��s��㳴\�x$��^�垸�7��%�9ryFޞٓ.�j�%#C[ٝ%����v�rͷ1f۰�QP�pa^�Yg��ݖ��(��=m�q���k�ݑ�v�rr��O@���3gi6.�/.��N8�:��<�s�7�F�ڎ�K�^��+���v�`�:�nݻ Ѯ�ѬBns�nx�9�a���<86۳�M���1)�N��f��tB6����O��K��=�\]� m�vPz��@6NC{0���oc��y�K)�.�K�kj�Ĉp�g��cu�Ӗ6(�Dnl5��ļ�:�
h�ɍ���{�7&�`�\�U�u�1�dNv9z�w�����_F���s���cnnE�%�a�w�|xʘ����F!q�>^Ѓ�Lu�������9yw��9���ם^��M��9y�;],��l@r�7u������\���vg �m{{ �k�Ʒ��=)�2�הMɵ�k�����q.]a���.�sjk�bN6�ud�=�}�^�q̽��zVm����:��=�6|�Oav콲1���V�n�Ofw���˩�9��y7v#�@��V�����u����Û.��2A%��4xB^Iy%���>@-l2Ɠ6��g[ԩ�K�$���д�H��ޜ@V�.�ݻ�z��j����,n�\Pd�A$���y���O�2 �JG	5���nkE���ʺ��%�C<�;w(��M�fiˉ2��2-.l����D��Sg(��RKɷ�D�^��NG;޾�҅�#R���{}��Z~���w
�-��H�]j=	I ݝ"d$�M���<^�,��Uq�a$����Oo �-&�	�]�w��pQ�����r�L2Q�YTM�t���Iy6wH�@2��z$ϒj��ϱ�N�!52tX58R#/2%�X�B�({,U�ʣ�!��a��P�|��;�H3�A�A<�Z�	$���}(2%�}�x1�QG��h甴�s�HϮ#��D���w	3<k��G����yR�ϧI�_����d�����e\>E'1�Bi�15x�&ړ�z�Ⱥ=���o[9�{�ʰ��6f��={��"�� =�|����ې O���ْ@%��g�[�f1��r����v������M������i4۲�+c��o����@�W��ŷ{�Kzb��rɝ����ɗl��tFo�^-���-=y@$�n�ti�4�g��uI���ك�E1s R���Aٰ#��7SU�y���)��@'�<�n�ٟ�)�_l��EK�͕�:��ؒ!��?^B����N��=�Nzݍ��Lb�;m�sA<�`cR��Z�<�d-��y�f�	�%m�����������Am{j�{/'.xO�������`�vIv(<��}9@5����9�p�G�!u�D�s�{�@<��"���^>�=�	�]*]����Mϵ"I*��> G��ט"��b'&���K�Vb�'�e�ܨd$oQ���X�N;盝�G�wk�Ў�~<�Ұ�}�C�4��
q��̙��p�5K:�("-;�=�����$�B��ْA ��_=�K��V�.����}�~��ǧ�Nu����O�$+ɳ���s��r�����"Dî83"�;3O�]� �G6[�)���]�Y�z$@+���[�_8���C��_,��*(�d�Hn�μ)
b�a�z<���M�8��:BVWE+q�S��k���!�)���m���$�ۛ>��;��/L�9�s�~�x��>'��nt�E�=�����P5���fSo�����:8nkDG�(�"<�A>��	F����Z}D�c�`�vIv(<�񮋀 m��<H�u؍�8���||��'��=��N�%@�g)3�M�71�m[��r;sՙ��� ���A �^��H$���z��=�Q\�������ĵ�x-����C��WU��n-�!P,�USZ9��>�x3U�������OQ�x�����|������ +�Zr��e�ۛ���M��j_c�o$	���w�N���.�3Mє�3@&i��4	&b�v�w���u�[�p��ڈ��v��h����Uy[+��^N�w(�m>ٟ�QDH�w:d�b�� ��g�X9wO��	n�lUn��;�S1 Sw\� 3C�z\"E��P�#��n��|Vv�I�s@�$��{UVh�3�*��b����'���M�9����m6���h��m�ё�� �w�-�A$�ooKxϫ�rwt�Ȣ������]���z��	0�O �G��^w�ؕ�-���l
��Y�C��rz<�i'%�1%��N�2���~3����#u�{�Ő
!��H�΁�V�d� �Am����z<��jY�4C9Sme�*�#�-����;q��w���^K���������'����=Ԣ]o�:ڞxɢr�k=&�n3\)Pvp��q��3���<�ڄ���a�Y�n׮[���m�n�ρ�(;V�=��[�\;�8�Ҟ�����=l�I�2���s���lfp�~���n�p�]�3<e�v�9�=��q.�:|���v۴�:˞ý��݁%�u�i&K�K���/.�ǋ>{j囂v6�Q��;��;eۡ��<�[��p��댧6��]�7jw�=���Z�����βMlzt�=e3�k�gy��Iq���~T���`;B�÷�2�m��ݘΒo����Λ���4N�@��^M[|/�2�0�̈vd욼����o0���[n�A'˳rkԈ'��w=x�9��i�~��`���g)9sT��L��A}͈ �9W��*��š����L_}�e6����e��뻎��9@��ֽ��dV�owQ���~k���O�$>�Dx�.�q�$F��
�"�rA���}L{�� �:W����y�MM�§˚4��_�Ot�Q$=�8�[�<cF���i���t�B�\R�DP$"�ӹ���<�N�e���(��U�l�#MT �ͽ��V�Gc��?N��>!�#˻����;0�Z^�eT�����]L��sng[�j����3�@�(��<�>�O��)�礪��or���r�i�v���F�3j[7F1*�k��+����~��w�����������1��y-6�Z�.m[�
�T����CA��|��xxO�z���|>�b<H���H�ŻM2�7��,��XzL�+���˥'}Ŗ�iOsfSM�(i;I�G.f����+{�A;�6.��vt�)˘m��Bɫ��k��ͬ�N����Kx�C�\xA ���=QU�/��.|B>5�� �5h�.왜�;<�5�O��M��V+a�Q���3O$�@����3�X���,�o]��AO���HeE
�P�d��z]�[���6y�s��#]��Z#)�s��#R��zA�9	 ��x���1��oH�tt���A�4�*�#�VI�
Q.�;:w�P�ꉜ$�2��w�흸�>$�y� 	3�d��jrb:z�ϳ�j+��2�xm����k�4��������!+2��%��.A�g"_���_|�����-wn��%�A���;�ތDI9O:��f�+����c�
�u+'}f �z�5O��� xK�}�]��$��}��$g��Xn%����5Qf�֔�,$��o�\@����HD1��x��Pjr��`���X���H�.j�d@/ٱt�-�6��� ���� ��|W�&����wl"84��T��1�$n��9���w�6�^������l�j��ŭJH�:�������B[FR�[᧏p��~�آ|O�{���|�ުzn��f���I!�3fI�9��wtBgE�&�-�=U��}`F���	$7VlϋyyQ�� ��;�aY30GB�+h��D�F$�w.�&:cf[� I{�A'��I��s����$5m��m�{����OٺP+J:N�����o5��� 羉$��ǀ	�!v� /��N���Z�*GA���2�Y}Ϋ'����KxU�l�F\F*ҫ��9S��dY�R�<"�ø�l$+��Lo/&�گ� |L������D��Y�	ػ&�,�\A$�c��aetTeU>�zA|���[��(sW��Zǵ�[�+�rZ[dtl��4�Az;i��"��չc�����Z��Q4Wa ����t�Z�Θ�A9s��m˙$�Q���/+���L<��wR���{72�M��{�K/\�yd$�`SZ���K� �b~�ۮ��{	�$��
���J��u���,�=��x'7d��A�I���&��^��$�Y!�7���X5䣷\@*w�@ #�d��T�`�ýTt�Os�n��qx��>=�1���_l-�]��������=Mw������Α(0�5�o<e4�y�� ��lI��t�(�G4=�7�#��b*s�A �-���?��"|�I�Bw:rz�f��T��ggU��{ /����xڹ ����]��s�[�ZE�������x'�Ŀ�m��O�E��:�g�����R]a�9� ���m��m׏a��pw�|���l��6��/J�G�ὒ�ڱ+��ʮ��.�=\�݈:�v��*�9��Ou����;O�H�.�k��������{][рI��8T��/%���������^��n�J�<�5z��k�gu�-�6m�9�-�[.	�ݶ���j�l֘�zN��'Ynm�v�Gb;<,�Z���ӷ\�s�=��+��O��=�~�Z}�uc��N�{s�to%�/78e����V��9���Ȋ�\����9`�yn �
�މj���f�����p �B��vt��)˙����� ����׎ �I��@�Wf�� �m��e���g����X��:�t��5��Ǿ2�m�{���6�F!�����8W��ay�n=>+3z4�mYl����(<�񾋾�ۆ��A ��<x�	!ufL�������+{�}����O���fj�`��=P���A>/}�"��x'������|S��>'�?ww��Y�<�̊'�ƪ��ak�������\�Q�g7g�j�V�$`)##+yzo�����'���c���u��M���ry@�22�kF�������彽2e�ާm����Ғ��Smc8����GM�1_�ݺc��@Z3c�s���ͽ���WDJ'�k+��o:�?�t�7�-j7[���?$�c|�
�z.�\��1���&W� =��6�H$�}#�}�o�A�!�E�t��v��n	oLuuݝ�:E9sUx�s>$c�c��S��{��A�� ���#�os��8�t����<ɮ�x��3�o����܁$���<�@އ��>[�6��"���>�4���'wD'tPy�{"�e:��F5�I非C�#*�O�H;;� ���� M�΂x�$�!/\Y��<sB�F��$��Re^�J�x:�I�J;(��-�w.�3�Ld��$o���p'�W�Wt�5J��wsD�\�zB$��_<{6���[ZZv����}�{��td$.s"	��� ؛�j�㢓vh�-`�2Aػ��)��@��^g�6�ƀ���xv�ӧ��ǧ�o��:t�˧N�:yt�ӇN���V�1�^eAFR᜻=�"��,��������z���g-�x���!1��-Δ� 9!�o�sw�q�I.)���ꗏ�u��w���y���1�#wX�әA��1��0<)��ON��mw�v��a�ĞQ{o�|��3�� �g������B�P����<��7�+�5y�	*&���F�
�ƈ�uw����xA��x[��m��8�,���zE���䠁��~����ϧ�.��]��s��^�P��Gf���xn�[��j��Ox����4�o��]~3����h$���*�r9
eBGsȒ����	����*�������>�����x� |}8M��ўj�/=y��&OyDW�����!�|<��<�L8�>b�u?!-Nq��)��M��w��oMА��l�s��Q(J�����-�g���Ǣ��Ϯ�,���y���]ؽt竕ڱI��݋^�DܾÊ/7;���{&KI�}#�����g�ܢ��:`/(�.��/�����m����|�z�������O�>�}_��t:���n��zc�Z��p�:�I�@ז��}�=��ۇ\1�����6�X���_!����W�u\���n{x��gs��|Xٔn�Q�g���p��g*h?�X���=m�5)~��S��,n���o��S����号��}���l�3�I��/�Y�?�ǖ�Ż� �+�@m�Uʆ_ޯH�;"@���N!����w��ZX7R��=Bh r´�~�\o �]���E�S][y��1)�!�'��ğ"�l�*d$垕�UQ����T�59�VI��W�RZ�
瀓���.=b��H_"_?,2(���>�9Ug�\g����z��RDg�YQ�TG��x�UNJ.E�j�N�����-\����K<��%T�EWM)!<+�#�̋ʲ��<�u0���
Zޣ�՜�+�E�h�.�Ta�UW��DQ�j�J����)ʈ��B}EuY�9�Rg!�*�
痡Fz<�i����$*^T=y�UEޣ�"�("���")̗C/2�"����C)�(�����J�H��3J"�*�"�� "(1TUҕҨ�����7(�2��J��U5�ߗ��y^x�9����Q�J#�^���$�� �fIVFX�	�d����zx^V�N�nG�B�(��j�E�RAW�GA���{b@����gM��A>;?s�%��	ȣH73;�t�r�@�^?\���F�A�I�͏A'�]s�=�o�+^+x����ݘ�7�̬�{[{U�����2kf\@$�:$�����i>d���O�n��j��T��Z�BF5/�����0����q'k�$��n�;���:�ف��M�i�U
�[קz��G��w��)���� KV�L�5�W�����%�OQ�1�O�m؏=�/�4��vd�	�����n���=8'"I7Y���5�������G<���D�<�Y��,+�?� +Bei[���$G}�gO���M`�ʔ�m��T�@�Ij������v"0�:N_{�j>�|*���.�a��	�vfO���������+I������ǩ����1O�"�iڳ�+�>#��h�0�w�3�qŞ�o_U��ku���n�tW�"Bq������Ϣ~���|>$7o@�rQ���"������$��_Fl�ޡUX���+w�<@�A!��g|E�Ҏ��i���m���Q_�'�����5�[�X}����+pi��{m��n��0Ic	j'�߹:�#%��������<o�_�I$�~��c{Й�� ��A���^21�p�wdBg)�v=f�Q-��v[�����c�����S�lͥ��K���vӴ<�������|�2p^g�Q;2H�$S��.aUq�[�ǖs��$�}����OǼ^|����;&V���	_�V|��έ�ǣ�'q��A �m�<H'[���LL7����O�fq�q�\��-��[�s-<-^l��\S�������L��oy�}��<G��=q��fD�'�JU�&^g5^E�rr~�C�eߧ���D��N�ǌ���&��}|�!L���AQ�2�R�yql׆oz=Ǻt�i��`�k/�8u��gߍkԞ��F���n7m՗��盕�z���n(���>����R�wp�YR#r7f'v�����'H����_4pQu����i��7EW=�W�����i��5��^�q�-e��;[��j4�4C��'v�q�Z�����Ϛ-�S�/.��y��i�t���c��z��J;������t�V۳��<���p��8�kGV�B�/u��ö�7m�v�F3n9�����2�쪎J����]󾕅D���}ƹ�}��	>�vǄ u��s�o�U�t� ���D�/�.��N�<�������L/����F�m���A�ܿD�I���$�q�-4�ل��k��wH��Y�7��9>�M�s��/*O���fgOu�}��r< O��l ���x�:.̜�Q=/1�j�	���>$�n�	$svt�Ċw��λ�c��Z�L奿-�F@E	�9{�-�@��ؓUY�:n��Q�Wy 5�:d�٧�F�d�P>-N���3�m��ݶ���^1��}vQWU#*b�b�+A�^�}\�v�[�a��ee�Ӟ���4�w:g��Y�e4'ɳ�}��� ��(Ss1w`�$���Uے$y��y��&��7FS��Z��y���=��y�E��{�g<fR��*��*4�}��mK)^�G���tB1l�7�Վ�����f���� ���߄A+/ ���ddoYY�)��,Ǫ؟@�Ձ�$铺gO Q��q��y�$�W3����tg	3Ϟ9���nΙ�ŸK;�Qg,����p��`�4���x�E�kă5��F�o"	�2	�Oݼ�s���`پ,>�f]ϣӡG"Z|�2p^�T:�dy r;�7j�{a�^�#v:�2�}"I_��ƽ��dw���Ş�O�E&rWU(��Ջ^!s��Z���u&�.M��m�t���(�E	��m׀k�[�DO�>$s�D����#�ѯ�<IzMf���Xb��N��%�� �_m�.Xμkf�C�$H���H���@ �|��"$X��	*A��b�ˠ��3'ʻr'���������e�7a�7����5��3�����[�Vnn��V���7k�F[19w�P�h�e������K2�&&.�������|E6��!(�A�>��+�&�`gI;2wN��G9��:go�y�Ex����{˷\`���*���Y��if�$t�L���pwI �Y��踎��o�^EU���%���4ٙ2O��n�q�wlx@��&�q�����۟�<Z�L�@�=��6�����<��������A�߽��,=�k:Do��|Wv���r8u7��EH�HD�wD���^�!"��ƒ���^׽���SL�\`$O����$���L�$η7f_��{���LM�XK1N�'vhu�n<��Tt�ܾ{��H-ٰ#�ol3�73N]���$*��փ�GmI����W]��A sv���oo�~����N��O���I���A���� #�E�۫��[�ݣ^i��k����	i�	��}��V}�ܞ7�ֿc	~����e�+>�$��!2k藂M�ϑ�Ǫ�`k���y ���A*�a�`�N��L��sH�G�̯�i;h�<�j��uz9�9�v�q�e8�l�r���#e�s��R�� v#����yYm��9����o����[f��>G�����/�"��D��U{jk�Hf�cݛ��$�e��6�H��Sw��^�������-���h�Cl&͡,׀I �m݁!��0�����/�l�H]w#���|�h�Eqd�;�٦AM�S��]�gU�x�[�� $���ِo�x�wB�h}�﹙S�/�#�:x�lf.��	9sU�dxn��xtYctuH&�.=�wd� ����ޏ7�5ݳ$�c����H�w��E][0���[��uX0=s�����ܔԅI�o��f�?��y�A�_��=�n=x�m�靽��45+��{�ߋ�o�� ���<���F7v�.8���u[�Y��{[v4sZy,K�Zd���G���8��x6����n��׶z�v�c#�l=b��y��C�.sv�۶�u���1�r{�-��=c)����U������h���w �ckn�89������\�=8׭�ٰ��v��!q˸��)�+�ݓ=��.�ы{;/m��}������a�cs��w�T켲�:�CP�3F������'�$���i��|�t,�߮���6�j���2Yn�u�ى�G7l$m��>�g6���Ӡ�ƺ*����4�f��m�R��v��	-�� ��ZQM7C�,Q"�i��|���i��'Ė��	9}}��+�D&����c���U�^A K�DA�e�'E��;��f�x�!U��=#w�*��$���"+{`>�D�k2�8&.��|
�Ue��@�+_,:w�Y�xs���Ǽf��&�Cu��8�UI ��@���{`H=-S��ܿ��3�䢉)�7&9/dk��^xz�1�1�V��֭@�$k��Y�[�$������p� �ݚ�H�� ����{Ζ�ѓ�U �W���7� ���ؙ)"�l�n��&��۔�G�?�F��?���%w�ɠo#t֖�guyuAܴn)�|mg��J�y`j/�)�Z�v��@����"�C��1�g�U�}�I�!�>��w��c�)-#�uS�kFt��mְ��$��v9�F�r ��U���,)�^��q'{�I �g8�w@�E�)4��)Â�*:'��r��HEm�Că��% O�%�"H[�Ӗ:jͥ*�����uD�:P��`]i;}�e?�$���t�Y^�v�T@9s��ٮ,�B�ޞ��x4��O��rD��wi�A��`'0�%�S<y(�au��^3H�V[KE\�ڥ��=Ϧ�
尪@��Sn��,�p;���'(���g�gxsØ=�egbE�#�=*!H��s6��2H�*b%�q�İ�y͖ �J���An���FE�_>��+�ӀA���	-�V��KO�kFSi�����oog�j���c�f�J �x'1�qS6�V]�t�S�.i'�l!���F�Rn*_Ӯ�w�)27Pi8�0&���N
�e�}�$��ހ����D����a3:I3���<�5�Щ��\��$����	��bI���s��'�/��7D$��A'
���� ��;�D�ޑpNv�z<H�� H ���1��c�˹������mJ�%n���¤GEO�3�8l�� ֍�X]F RF�VkK�_BXV�}�/:e�i��$�I�wkz �I�:""�t�Y�Nϧ½��Hw?�&��V���O��Nn�tuw�95t�c�q�� �,Ͻ�+��v�#G]o���H9Cm��L΂L\ٞ� �ۛ��A_�=�AϞ�/װ�>/ݱ� ^�N�3;g� �Ļg�Z�Or~�GQ%<�Ă}�H��؏W���py��M4æ[r�Z��U��N%���A��g�촪wN�cu���S������=�LasXAQw�`̦��.���[ݻ�M�Z�x�3:I3����=Ǡ���x3�y����'׻S3�A ��D	ݱ癶X���
bQ�dPd�b���#�z-�wF�h�:E�¹��/u�eԙ$���Sg��\ݓ�>$�K^s����m[��8��>e̙���;��]��°,�s�1�fJ���{z%�T�x���I ���H'��� V�}�%\���k�I����k��尪@�TSW<A�x$��j�E��RP�)�,;�;_Dx'���:��7�"�L΂L\�z�ػ&߽B�nO� �>�x�{���� �G��;�`��.��2I3�@�	�fd�ü��}SI�G��sv$�ؾ��P���nCUݽuEq����T{��ޏ�_\=>�>>>>=>>�xt�ӧN�]:t�˧N�<}�߶N����O緄��1�"__C�����y�@C�`�C��-����Uņ�ʰ�V�q���GS�i��K۹s"�^��3���Um>�#�|e	e����������l��{��S�N�s;��������w��ׯQ���8�2)�e�O`Fg`"k�
}��r�h��S��B���3G�-���e�gz��{y<'i�{k����3]\��F�M�몭c�W��v-��mz�0�ww�\���ڻE�N@��Ո5�׻�%����t�j�ܼ�aȞԳpΧr����5ӑ�ٯ��7x��|u�7!B�7f��wbO�\nK�u�<��Q~��Ӣ^@v���<r��S.�N����|����� ��޾�Y鎻qzcɚn��\��l���Sہ]��G�(�n�U�L�4h�f�S~���\ܽ~����Zس�}�75�h���s�ސ��=f�L�;u�3�ݼ�ډ���c}ۥ��� �o���D����0z{�c��?yo��ۚV�<z!t�ē7�k��� �^^��T�
�{7w9�w1��w1�ӝ�l��lrxd�&�*��]K 'x�٫����3�f�{f�|�k>����}��|�ӈxnB�;"�q��{�@=�X�d�%����5�o�!�V���G}}�w��j�1������{��/I��k���{�1H�����zQg�B����j�j���"O��!�ף���s9]�i �"�~~尴�@x]Slݡ��6d�`���s�^��v$�J��M\���J'��Жa�Ԋھ�I�n�ߟ�����Q�W�E�b	V��@QQ�n^EVa{�:2H�/#�O+RǑsؘ��R�RY!ET.���ܬ2��ʏ
"*�U	5t<�W)�hD��L=M�""�]+�I^^2Ђ#�0O3J��*m/PS�Y�G��'(h������y�G�O=:
E�<���/d�m���]�ʈ�/Kq��aAS= ���C3��H�(
���Ͷ�
����UUL�T�t�"��]3"!=@0L��4]�Ą�/Ҽ��4*�3>��/#�RrO"� ���SȷR�]s���
�g"��A��-��f�E�E�sv��!H��h�^F��9���Q��Z�̈��"�M̒�W+�;��W�!�#��<�+���R�N�k޾���̀�rZ�픏\n��pom��v��m�>9۴�l���
Q���K�R1@T�Ĩ���QBs�ݎ��z����-]v2\������Ce�]�zヷ]t�j�)*�0�7��iĝu�kA�$� ��<�/m{���#cj�.Mf�f7<�s��-も�"���;���q�{@�]�mm�u�m�YB�uǋqnTJ���?��>��q����a<��Xt��=ZL�=�ضݝLmg1�K�+�CV����P���&�.9ދ�u=�஻U�Ζ��t"���D�ֽ�\.ܝ�u���EۤI��(�:�n7k����-�+b����<�,�g��i��%Wctov6��|S�q��b������E;��m���W���c���/�D{=�rq$ή��f۠��tPsȼ`f�v4=7W�b.Ly�D�V���w"�����[qnM�Rr��%p�\�m�#�	��ޕ@�yr\�x�COl�Zwg��3��.T7]=�s�ݯ�vm���܊��<V�C���q�[��\��c��q�PSL�k��gIr%3�t�ˡ�;v�g��OOWc�b�g!e�N�v���\���g�[�0񃈳V���v�dgmK��n]��M!��ݧ��Q;hWY'����Sc٥d]���c�<{v'�v�A�)�;�gq��*�8�.�s���x;�7��=�>�]���6��Le��@�㮭ּ�o�ے��]z�v�go����a�����|>�ڶ.Gu�a�㲹�c�떔�G>1͗��nyk���ݔ�q\�S�ems��у�_V��u'<t�)��]\�>�i؝�u��	�b��A%�7����r+�B�e��ct(�Ǣ��66��Ҟ������Έ��n��v;v�1����>���ۙ�v�.\�b^k ��n�k��0\NB�9���X��]v&��l5�9;���sv�^���C�U@��D�67��m��_k��Luʼ)������V�j8�Q�L���d�5y$���2�J���͜�	x:����v��t:����=��d8SRm��zD�<�cs�kC�p���!����{R��NwQL̥�X�>~� �:�1s\�^�yd]��L=qȅ+���Ʃ綳9\1�b���ݷ��jzԵx(�a9ob�E��M�끚������j*�C����$����c|� ��Ug?�č~ޙ��z݃˗>h�軈<�{H�$��%5y�L��U�ى��KyD�o�|��}�Am�	�}ޙ+����)�'gN�3��.���M?vߦ���"DJ�cv症��	�!f� �H����"���a�nt����/})ɡ���g�3�y���|G?n̐�-�̘��J��Hk����L3:2s2�w&I ���(�l����� @$Ϸ��$���D7���WwT�Ҩv�ňp������`�$�6��=�>J�e��q�o�hɴx�J�"�_-/��	-�tw�{��e���E�D�������rɕO��t������Ii�������Ih���y���ꅲ��6�O/.v�2몼�A��^\�z��O%q�Gu������}8M�Ř��K1l���r�I�H�ذ)�_g�m[1���Xc��0��M�_羋���$)�zk�<��x�� ��3�����M�4��L�R���>�>!_s�(�d���iƿT�CK�=�i����es���BXR���|�>�70�g�l����s�o�#��D�؁�-΁�h)*��.4�z�Ǜ'���Y��9*��-����[o��
�U�F�����ueL��I-W� ���{+)�|�̻����O{�hL���a���x�`b|��^y}�H,T�TP���H�t9��o-�ٙ���r�� �	-�� O��΁~*��F�wNLܼ�ĂHl�A�/}���,&�{�?�c�2v����c{`檨��H�%��؂I��t	��
�|��桩��q��w��v�w�ZI
& �>�� �A��q �z��tI�WŌ
=��x=v^��D>»}׬��m0�xj2�9��������%������LL�.��iә�E��4i_�P��+�>_�}� G���ϤI66����A0g	L�t����ո��X�ȝڗ	���/B�-}ާ���p���ǩ�=ռ�B:RRJ\�8{��o���t�q&xl�De�'� �~ޙ��k�i��0���%�����e�`���6�.]ڱ�õ�O��rUH�؁����D9���x$��.���U�A��V<x�K��w��(�c%��C��q����w+�#)���3'`S'5^]{�$����<dq�N�y��H��[.	wLgT��[��o.����9q!e}�(Ik���+��^^$��Ή ���spb��m�@%6�7w�e7q'}�{KK<9��ZI dw �ǚ����+�x���l��< H��>�H'������y{��d0P���-���U����Gp�B ��&$���{�;%yR=��z�7qi;��^>� �ku0X[C4S�
#,%A��oP���|@w�s� �ޜu����&�(���#�s�+$��z��ʇ�;6D����e�W&�S����$&�����5�s�Kc��<�J���¹
�M3QƊ��;����vtΓ;p-��/���GLz<doJ�M"��f�iE��h���s gGt�1,k�E�Eݚ$n�EyCX��ŐW\�\��$�f�rdx���l��bv��zۻ�S���3;&��N`U܌���旎�F2�q�s;|$���N�lzz��	�f,�˽P=�.d�+}1���F{��q|�H'�ݐ�5³��56<B�'_*u��qÛ��@_a|�xk+-6����jr��)�Z�ꛃ�<�>=� ����W�
8�-�[,�� 8'I`����ˢ$;�̏OW(�/)8���ޝ�G �q�|�^S���x޲�?{ʜ���Ρ��7��nڳef53��`�1��ùZ��J�kB��[�}^OUF��D��ۓG:�Y���컅ʻ���m�Y6��:y=�tֳ7n��pn��ڐ6�:7]��s�G��Gu�������s�.;4�Ÿ8��c�js�q͎`��^�n5�ܒr]2����n�-��Fx�s��\1�Q��K��l��[Q���\[���.�>�ţV�i��v��v�n�ۆ�x����T]��p^v��V��;H��uEjtR&�24�B.�K�KX���vd�@ ~׀I+� o�)f��Hs��ڧ9S�/R ���C� �֧�E�R�l�tSx��w~�ڛ𚡍Vb���g��==� �J��	�xa�����y�%z�d��%�.��4��Ͼ�$^�  �8|G��3�1��þ##�c�Q 3V@��
�\���`S'2{:��bּ����'�����n�q �A�}��MU���Ϣ�����r�,�s�Uih0ְ��e6��΁.w#q��c��ح��U�#��A>�|�w'v��"�?5�C>IN�r�֨�u�o&�W;�#i��콱�e�\�����(S��w��W v���~�~��m��x�$���D��mM��غ���yq$,����d��|�&b�G<�H�}���7Pװ�N���W4�YV����Ӆ=���E^yԲ�4^���~Xj:��|"���4�:�tՀ���v�Ƨ���� ����>{��	U�%����F}R	 �����ۣ�_��^�Gɧ�s���R����+�I�� �c�Ă_�K�*���7J7�/�U]��k�L�" �n�y��vi���lw���Z�-�AU��'�&�#fH'��%���ұ�&�.�q��&��N`���x�O>k�`��O4��`@>Y���{�R~舨5TZpL<�;���E�$�DMĢ���&.*p<��I�\���m8��P%ut>[[��$���a�����>�.�}�$os��x�s��wv��Lz[�����ŸY3�N�]��z���ąOƌ�F�x��|��wG�{v�,[�t�M84�O�^�
��A3:%Uk���$	/y�����8C��2�#�ɲ������������}�ۏ�ooksvA���!�ϽN���}�������U���?y�}�p>[A�/�xV6p��璾��I$��{+/����~"�����+5�YL���g�+D$�؈���	 �[w`@%wd���ݲ@>{���lzfN��X7��wf�V�$��o fy�.�k9̉Ż��gĀH-�� �V�@��Y�Det���*����]��6�d,�N�.��&��<�7Av;vJ�B��j�h,���'W���HV��̜�.�ɒs���z	>$-� �����������7���dl��+p'I�gd�]�=k:)����\6�xB�ێ���6�J�xy���	/��ivF�T�3S�S����q��H_#)�gYK-��t�i'yzv�����|H�j܈!wd'�}Cr�T�:	3�UsDtH��ğ/T�kz��������^�@��������N���׶��.�vX��fK�ke
�ƕ6�`�h��H��^�������A,�߳����ݻ�۲&=�q���S�f�|a���m�po�"Z�����v�����d8c�xGZ��9E3&aw��?}�r�:r�:;�t��@�n�H5����yB����ͮ�#{č���H:ܭ��DwF��T+޺���)-��8�k��q��I��-�nF .�
3;-�H�RW(�G:�ھN��6;7v�~�A>:ۏ�����<U���K�S5�gM�߻���v�
A�`�!uuƑ(˦�_Ih��K�=��W� ��E�t����$��<eWT�'Z��V��: V�vE�gd�]��^8�/y"v�:$F��\�P�VI#��@'9��A>����G{�L�:N��F�ּ`�&_8kݰ�>}� �I#m�&H%��;Q/1�Z\B�~%=T�:��'g(�IS<�;2A�k툉�8��Z�*�`Lo\-��T_L�In�H�O��{zce�SEw3��&�..�a��j�.m�}q��Щ	c��/�=d�����t�Rb���y���ǝ���pM\ǖ`�(6�l������8�^���5��f�Nk�n.�q��jL��]�&��c� _"��G��<�4���������WZ2\ez��˳��kq�1mq�r�8w^C�\k��$�u��mwh���	�.���xn!3�n�BXMA>�[�td�R�|�`|d����}]J$n7Qn����'��۟b�k���������;�Ro/>�Z�m*�vǛl�����P��@�nu��a�c������$t	Ie{��>����{�Gy"]�b<lk�θ<��`Ƕ́��S�L���4�`�g%ݚdݱប{I��/h��n��fS�$���$�Kol@>)���IZ:�_����
�:pY�fNj��ܙ�$a�b	&=�]"���V>�O��2dK��G������qU)`0��?p�c�Fe6ë@犸����#��v@ŗ'3u�y��|ٟ)���Y�ft��ĉ���@�^/�=� �\�j~��n�5O72O�y��I�7d-}rm�r�;���P���mpM�]�ϛvɛg�nd��UT���v�VV:���m��2Wv<�H�K^tA$y� {�y����O���M�ӻ�s�p��$`�0Θ{\G����a�a�#
�ٲ̠p�W��kPߗ~��~tGZ�Ȯ�<t�mQ��F"����/;^���o9��R C�9�Ne��ש������Ik�x�����A��+]�\�>I��s��x�Wl-֜�����̒-�V�k!�얎��rwA��D@$���0��gN8L��eu�N��~.Pq}�`{4�k��J	�� �g_zM�\���Z|I���A^���'v.�ި��	��|�F׳c��P������s�D���J�$�{���-�s�V��.�^E.-�F��{o:়]��ή��U
�z���tn�@���\�g���;Ͻ3�v�C��@��gY1� �O5�y�h^�TY� S�%/U�����'��WW�׽��-��H�}�N���v�끑�<���"�P��t�x�i�����I�&�q��;xr��o��_YӧN�:t���{<��g������(�ȫha����hisN9�_��<2.�ӻK ��i��<P��̥*f�()��7����I���a�!;a�����x�+}��aC��R���|���l�g��8��{9�+����V{����V�:P=�fe(9��.Ɨ7��w��ܵ,4�����A}+�"KI�ws\}����T��^�A��]f/TϚ�r)���s�xlK� �{��C��ۥ�8������=���x2�Z}�B!Ӓ�[������/GS3}k"=���pc�*������ 8&���0�M��x��C�tH��ܻ�����a��{������0_��}�� ������������<�z�/i�Ϥ9p�R�w�}�hxzZv�M�C�~��P���i
;�s�Gn͋�F߄�|�Df�=���N]���!�8�[���������^�r������T����Ћ��4_8X�n��^�0�m�v��ǭU�A�+ޞk�2�'/�[=�St�X��{��X>Fu�9�2������m�����u�(�k�R,��l<�<y��a|���pn[�st�;W_N4|�6g8� t
{eo{��B����������g�W�}[9�"�1{�՛�n{4�I�
�pv��L{����l�����_{g�'�.^3�6][����g�k��%F��~�|���L����4���r�pN$�>T�=�>���8@�zN�8��"�'ĜX�)�E?�dxQX�$�DɎ%v\��1���q
=�y���RW�AJ�S�A�["�<K0'�,���
����)�>l/z�U!	h%j����_��E^^y{�Qw��o�9:<��<:%�QB}l+=*35���{c|xʂ�z|��(��9AL#,�W*�Q��C�>T�*	�����G�vN\��t�#��\�]J5����J���	�V���I����Iii����$�^yRdb�FWVh�AZRŕ��t,�D(��8H��Aε�TT�ax���IU9g�I��E�4g��Uj��0�#�**�*I�y�F"�!W���'��d����W*
�=��4L(�*��מG���ʡ�q��q ��s�L�FI��� 1<�o��?Ѿ�S}��f@I��q��ށ ���;��z�q�S˔M���r��jc�����)襠��� j�B<�{�&���F���M`&� A ���A~�C�ysY�Ó�t�m�ɥUO��["���I)6������.2�0㱷`�$$�&&V�q|�Ρ�T
A;����c��o'�A$����sx�ŕ�Q�y���=ѳ>'f�EܖgIݜH�n��� �w�A���y H�͌����ͳyY�	{��nz��E;$w$��P���C�lA�h��Ͳ���т��E��̐F��]OV��3�~@#a��=��}ߩ��4�H-�O���D@"}�� 	���z��l�304!�H�mC*+����DoG����h@螉�b_��+�F�+6x{����vG߿uѨ��h����2�_����[�>&G����an���������o���t��*��m�C�v̒Im��kvG��v���<1>�Ь)e��U4��UF3	�h|�z��ǽ�{�CJ)M�7k�ݯJ�:+h�=��ݳ$�/o� ��5� @'�cM��\�� �KWt0 var�`�:w����O�T�����Ȏ�a"��< W��� ���p̈́y��F�ȋ����w%��wg�h�D@���x�c/.������6s�@DE����#�Ǭ^	T�v!'rKU{�g�]N�q�EA�����n�	����W�[qӟ���s��8�_p���#a�7}׀H7��٘�oL᭦b!S�z.\A>��� ��(.��^�z�o�n}����-�\��ogO?y�m��]�eYg�w4�`���`���1�I�]������p}�%���ݼ׳�����"�mw��^[v9H�*mU(�6�.'�^W������b:k�D�G�x���p�uJ!��u�ɉo���}���sd+G]=^ >�Uڱcnt�'�'Tu<���U��v��k!Ѭ\���^��O'l��k�K�2t�Yu��n8<�6����&�]Plmػ�N���;�;4����:�y��)����k�[+�:9�:y�c]H=l���Z��X���n���fm:9C'Y^v���]v�H<�mt�Re�V�o�������a/ߝ��V^�-��My/v�t��UT�	�4��5��	����"����ᙝ��]��$e�7��o��%� @$;r:gƼ�aΑŷr�6�b��ʊ�q{���@XP���M��I�|ϲ��&��ι�"+�'8�v�N��{}(�홙 `l�p;���;���=�4(�)d��R'g��Y,����z;va�6�d9��u{��n+�M� ���v!'pCU���Ϗ�;��f)֗Q�,�����@&�"J�<��{b+#U�����$���EŲ����.]E����W<��n�7]q$�k;��Q`�a�����V��~�����'Ě΍�$_�$t��W)_v�ʁ�Zj�_6��Λ�r��R
*&�M+{b ��Vlwu�{LO(���*��&{:ż�������y��ǨM�����|Q��<T�����?�V��'� M�H"p�4vy��<O�')�f|H����>xK�
m#:R�����c���Z]�{�5����ދ%{�f���ꢴ�E��CD��p�o�'M�KM��e��J����'�|w�]w�x1ˆ��'!�b�>$y�����#���A{��`����t�C���<�\ɠ���w%3��� W�s<<�����<J>��"b��I�>4�� �G7dWdS����L��?1�qQ�\𛁞;N��g�Wv�Pd݉�<>[�g-�U�	��.��u��H�]���Ǡ��ݐ |yd����A�e��w g�		dc�����d�\�BgvwD�����	3&�6⧞j0�E���$;��SM�q�璽�1�p��܎
�&�I���e'�H��2e<%�4���ׂ �wa.g��ܻeI1ϑL�wZ�K�+΋��:l��T���,RkS�Wh}ڳ�V�k��}��{UN��aBԪ0��g.�bbj�/�ż���q��� ���W��p���u�L�w�Tٔ��ff��oS�>'�k @	�|�z=p5�c&&�ɪ���d�h/��DR�,(kK�pє�x}��gO|t�r�z�#�������8�+z/�@5������s��sq�|�"��Kk�@�:�󍫞�������s+�:�lB�����O��iݜw�k�*��	�$���� �7\�aq�w��X2�q� �v@�b�CJ)������ց���?Y��б�퇒D�5޸�I ���wԏ�+ơ���sR�ٚ����.g�gvr�������I�~�D=8ގ��i�Ю�6�$�ˌ3�J�tc�����Nœ��gŹ�o�3��z�n�������@&��bI�$��^^;�Y�챗�h��=%fCd��AdiBMj�,Lm�IX��;���[�g��t3����)�ۛn�/�U����-t'�k�I��E	�l�9,�#����v$��1pɝ�H��"I�5�纣�\v�G^d� �e��ə$����;_)붳n��^����Kє�[��O���޷I�l�+1v�sPI]@�5���DH�aC:O����	>Ͻ	 �GDW�7d����И3���x�3���[Ok=�|@ܣ�Eb��x�W�A~w�I�}ȿPD���<��nAL��tVŜ9d�i�ز|���#�D2�j�6M���7"��bA>$~�wճ!.wg.�W���cD�N��s��'ĂA"ߺu� lFu4dv6h9Q�D@�p'b��wM2Y�`A"=ϗg���d���A�Ș��AQ� Cy��G��^�f*�=�!
n�1�U��i��ұM����l�gݪ#M�Px��c?><���t�~�jq�#4.��֋�yLp�C�/���*�qB�����K��~K���6,�r`M�<[S�kb��5�ȓ�63���Y��Ƌ f��4m6wB�k��]w�u��ts���S���N�Ƈy�ϱ���N��rg�/���0n�a��x���v6{=v��
�����c��z�^�8�U[N����<rcv
`�S��GXpn5���]����fx6�y����nq�#A딌�c�i��ro/m& ��-m۳�����Ю��� �h��--�q�:��&wʯ2dO>�z	'[����ѐ�\�z(>W� �A]�:L�d��d��<�+m�S�T��SQ	��{�@:ݏ���N�Ms�,�X��	_+�>F�P(����/Yi�4�=�	 ������j�=>D�����F{t�LS�,��UO3ґ������>H�OD�� N��K\���A�\�[O��&W��kQΘ`Q���a����I5ϻݼ �зg3��N@�O��#����萼��a��ƖsĒBj4�Rk,�*,��ƤA9���_O	N8�JMv˔R:ܮRP�|��_�P%�^ �v����	$�Ή=���|�2�'����� ����39f.3��]{�$��_���Vo��zz��b���<1�¬UL�k��{}zQ��e�n1^������g��]��|tw�]���[7d�ZE�g	��渾���nG����oHHT���ن��Y��A�v�.�3�b��#�����<���57M[О���p������F��L��+���.�p���{��@͙=�#�8���G�1��M�Amt�x�)_7hU�ᤆ��H��
Qv,Y3�g��=3�H��YCwV�Jm��H���O��Ft� �O��M;P��;u����'+N �D
�LBP���9�����ke��q�"0�����0(�C+��ߢcb@$��	'���/޸��q�w��5�T$�lȂ\<�"��D͹��sn���ŝ�Od��Y��� �F�dz=���Nd�3�j�7G��&d����1pɝ�hU��$/!��>I�7��h8�0��"�v:�!<�U�4[��wz���'����g5{}���à%�۾�Z�:�Z!���Z��1������ԸR	�m��~�Mk�G���@���.�3�b��2[˽<1�h�"�<����@��q����Vcׁ���)�"�-�b4f�L����vk91q��4ɭ�wk^X����0��+�d�|y����~��H먳"0�T\��$��	'����q�۠����+�:�Un`N;@V�:��>� �d�Hn�yʑ$[g<	��|� Ÿ#VH��W�52I n؎z�%��]ݜ�t�&�]�\@�=�7Qy�U�U=E�D�@�̀ 7�$P��#�[;��n�-��ikj�(W`�K�'���t�g��>�	��/._���bC�Rg����$JnȀA;�p �Nq���`�;��U쁕�Eݝ�7tVtG�c�z<NoFϼ}^~��]$5'�k��,�x���f�lK�Ek�c�6���>�1�wPeYX����6��̫�fͱ�H�%�{a���uGK�E��-�X�Sg�OTC�t�`��I蹁�&E�����س;Хp��]�Y82�u��M�w9D��� �[�z}>G{�e�**&6�u�>��6`�7b�R��)iЗr�]�N:�PN��;ufB�q�[QT*_qs̄et�8q�y� +�\@#{�b|{�r�-s�C����6�t7op ���6�;�,�膐+_��A%Od�i��O1@�{�|�bH�;2s�]沲U�d�A��%��Yݜ�t�`�G<A���	 ck�k|醸"���A9�3��#j�(WaK�'/��d�*��ao����	��H'[��K�`㡅�(����]ɞ:�&3��m^̂I�v#}�z�=�2��D{Y�}[ֹ�]�u�F;zv���||||||||}|}gN�:t�ӧ�N�:t�ӧ.�f.}�,� �d���˿�gy��i����b%W�ڌD�}��Ѹ����F����D�oq�1o<,��4#0*����`�v�5�ze���l��X}�L�������vY�����Xj��w^ʉ�{��A����nw�om^��[�g�O7��v�|=�Gb+eͲZ�_!�O�wE��岉��(g���[,����t9~���G�K/����L��{7*��ݐt�(g�n *��HM-�w��<m۞��#����_x@�vj��p���x����p�8�U���S��rl�z�X��bj+!��9�z��^�v���{�j�.G5��i��;�q�r�0{�x����}t�����Rʎ[�=��c�Nd���X��{wG>�qI����։X	��,);9=�8pn�Y�{�9����{�׋��"�hCk,���9왽}�Y�i]zyy��%z��[�r�ٯ:�5���0(Q���o	���jPiX�k���ü��tf�C��j`!u%�^���a���&�s؋:�ݻZA�`o����x�?�Pu&b��=#�Y�<@��#�OE7��qYlw_M�<=|�_x�L�w�{�j�ze��{�{ƹ��D~�y�3�6	��^܇G��k�iͦ��\9�s^�^���$%�Ӌ��ӏ#�}���w�����4��>�8�#gd[\W�u�n\K�>���`�7Ɔ�wk��=Sچ�a�/n7Y[����T�1�~Jd�E���\	��86^k�8%��(.V�K�݋<v����v�1'��l���5�7�IS��qZ������Q������=��^�Y��p��CC�
!�*�1����H��`��X�G���Uާ���Ո�YTQykn��R*�m�r)�"���Ik�zf��ȕ�i�8̙�OeXe��zrez�W�KR�
Tˡ��![,��k4�{)���-�J��"�`��ع�k9E��H��3h�[dgb%XtlQ�v�rT:$���r�O����ɄZ�1�*ƙE�%i�b*�&ѷΒ��!�it�:v1���vy�3��xk��{r�L<:&W��ɜ�4:��ڕs�/U����c8]�yXFX�'�!�i$�ճI&W�U6��!v��GU�0̓��n����鳗�㚵�:�(�B�z	�^v�nL%��2%�x�G�:z{(ܜ���۵��gs��;P�1m���7���/��ǯK%���qtq�Gի�feW�Aо�������ѡ�뗧&���p��.�c�b0����u�"=�\�u�����8U�;\��Q��){�����ovv�kl�(<d�xG�U�NIj�C�w{��e�܂��n�Y69����=�>�z���ȍh=�*nr\Znq����-��i��	�lݭ��-�۩H��77e�vn+�s��3����Ux��i��3<�.�qw+�m�m;7Y����Ϡ�d+�nݓ�����m�^�x�N����rz������2nқ�5�.��ݳ�[�J��A��"�k;T�oK�n-�xcʗ9�\���o+�Z�kz�9����,��P�CջOAc���]Yz77���"�퇬u׮ӣ�ݶ9�{=�����1�C�#&խ�z
ݪ��h�F�uH�m.�oeOs�ֻuێ�{�I�s�{y"��9ry�9����̻s�O
�Y��hp��w&�[s�t�u��cZ���GV��sS��yqN�eM�$���ݣ�c��+�e�����q��j��^v�M�pYݬ;��c��7�k6me�=@;s�]l܊7պ*w�;sѷn��Z�`ܞ��g��}HSΔ���/;m�sUӔv`؅�n���@�n���:�̽��]wF{i�Y���cڇ/ki��9��v�ێr��A8x4�M��D��&��5�a�2��ɱsvN��zR'e �n2�c��mQ��g��V��6�3�C��g�v�m{q6q����kSn������tn�u�b��8�8V��zȻ�kt�@�[�	Y)����u�ތy����:���{v�u���mh�s�X�u�vDNֹ�w	au��;c�OQ�	�n:dڂ�M.f�6��t��"�C���/Roxa���۫���z�<�˷�6?s]�g����n��q��ۤ|l�<O\�O.�[�et�V���\�ιy���a�t�l�l�A}�c�;^y�4W��ŷ<�<�t��p���ݞq���5�VG�֡�7��TZ�\�m���< 6��^��1p��݀�p쵞9bY��8���P��v�d�-�F�u�Ѷ���\�ۃ8�l�@�6���H��c�9E$��RH�k��*�T(�=��_VA+�=�9�h�m�ﻞ�M&��##�� |Cw3{KdʬSz�= �k�:O�ptfN�����O��.	��]w/�}L��̂<ݐ<�W��-�K>�>����ܱfgD4�#_j�I$�v��%��U�4sN��=��KI��}�*�̷|aУ�����x1�ϵbwUG��n�sۇ��L�e�wh�k�����T��ǂv,�t�/�7v� �k�Ǐ)�6ov6ҳ={�Ǚ�$�u��'y�+�A�����[5����U�X0�u��<ղ��y��ޤ��|�dvU�R�J0i���}�}��R�YAw؜����m>��+-�?xثҵ<�Ƶ���稛��ms�LFJl��Whi?��i��oƼ���sF���Ļxd��Tك6o�Y�,�����zhՂ�{��q[l�ɻ�W@��=�+=����{y�᠓dX}MF۾�p ��n�y��Ann�Aۛ�G}�̿-�Q2Q�i?l�V[i��^<I�g���a{�{��:ّ �F�\67"ٙ��ftCD���SZ�fݢ�O���#��./`O�g�������1�.|����-�s���D2�=��"�'bO@w�Zذ<��@�$Ot@ �my>'w�fM(�6p��ue�n)���c�#��B���4{a�&+Ǻ��gd�����0-�X��w��U�B��\�6c��[��Ѳ���tAh����^H�K9;c���&w .������w&��+�	"�Z��� �tl{�I{���f�[s�bd���û�L�� ��x�A��ؒA'�^�t�`��w-ܕC��ZnTd�Ľ7�(��w�/�n-�x{V���¨�[!�����O=��̪�z�ʹ�#��
%߸��]<c�n��{'l�N�L�D���Ų27A�h'��a��H��ِ��b�ڤ_���".�x��l�;Y��8�3�O�����ڤ��O�|H<ݱ,�8l#��O{u��Oo^pj�K�3)����Z�����lpp���K0�0�h����{Χ��B2�>�<2�p粴��o��ʱ�c�	�:A�g�-�A-�$O��c�;�]9i���=/q��Q��I�>�|�H:ݑ �s{�Ю��v	�"}0M��`�;��W{3�<۰�j G�9�9��>$g=��Sv9�Yޓ�!
 ���?]��\���������y�0$A<ב���� W����F6��L:���)m�ul�pg-ϵ���q����1+�c]�p��$�n���v��SN�mX�y������a�&t�d��Y8vp]��
;o @�I�}x43�Ө�VH�{2I'[5��Cz2X"��Ş��a�+L�nF�v�	�xӷԩÆ$����F)۱1a���_-}�Y)\v�5|�s�g�m����H'���u�s=XW3�$�9���X��S�`�)��n��Z}���tG�DOFx�$�~�����
�
�j�f:��zˬ�wޙ����K9t�U~��v=�/�C�KP�ʤ;��ǎ�|m�"$�Gtd�0�UX)�,�gqޤ�v5��|�\�gl0@$�F��Os�FH��~��k�Le��\���T%����w�-��w*k;��}�M���1�	�C::+}�-�'�^�KWF}��P�!��FU��`1kd���)ɰz�����gV�1�Y6�J����B�F�~|� u՞
 ��� ?Gq"@�D�x%<$�.9�N�v�h�����2=�;�v)�8��)��n��6�;%�l݉�%w[+�vvc\	�:� ձvpj��]s{{\���lJ��yS>��x�8l��;�������҈�n��Y��u`�G@q cz�o��	��zl��l�n(�)��7��\va�ۇRC�ўݖd1�8��Ǥ�6^޺Y��d荱 ��-ˋ.vn���ܝ�Ԇ�����<�"����F��!I��:�]+(�i=��r/������w:{s�^l[��{�|B�� �c:)2gb�3:!���;Q�"o�;�0�^K��$����C�/gGt� �S�p[^�i�]0����S�(�COľ�E�6��9�&I�޾��SWD����/.��-��Nĳ�NZ��v���ұ�VmQ���V��|I"��&I$��4�/zl?���� A C�]�& ��Y��ςۭ��O6�7~���z� B�D{�7��kv�vgm-��������&��W��$��g��Ǎ8U���OE�u�qk����UTN�u;�KEBYh{Ϸ�x$�k�q�"�&�� ��|��9,+W���m�p�u��}<�+(�i2����2 �M�j��v�{z���L�6��Ƽ�x_Z�"*hAC&�gf�qf�m}ߘ�������4��P~�Y,��g�V��'��,%��%��C>>�@��Î$&�vd�u� @'��"]o-�����V;'&NfgD4
���$�q��{$"�ä=���Ҟo�Y&��b@m��<{����K����C��v����2v;s��̬���7�'#&�}��F�ʴ�hF���|H����9tŤ�b �u�z��y�j�����kȀIݑ�n�Is���k�S��e�"�䘮��'dpg^*���tnB��b���*��0AB�Z���u[�Tݠ��WY3�I<۰ �A!��"NU��H�.��?{Zx������J�h�K-#=}c�6�6T��}��	4�� ���<O�˳�գ\�-��$u:���aD�I��>��u�1"~7�8m6���D���;����(�;�D|q
`�{{z�UQw�#�2�ͳWo�����3�^��y����5��s$/k���3!F�c�7�Ēu�"�$kv@�[��$�άE�8%���b�g��U�C;��bj�����I�q���o��7��On����e�� �uŝ��٘�Ovz#�s��ߕ�[q�y�b�i��e� A ����3r*���n��v	mqoệ(B�L�8����$h�/������i�9��Wi����_�*td���r��K"�m�I�$�>t�4����a䉇����	�΁ ��x��03x�Y��R�ۙ�"��_^����砓�m����^M�@P�/�E����\���Ĭ��[��DM�^�����\�����P�Z#oO~$�z�:$�M�� �D����$Վ �ѝ2HNwJL읜��>�h��q��;5�:a�Ē�y�bA �~�o&�ݞ���z�scB����.�o������n�&��-��L��1�Ϗ�[��ۿ���%OmK��3nƻuw��*�aüH��@�Ń8%���8�=>��o�"�ڼ�O��`��3ϹH$�v�v�k�R~Ҙy0,�$����v���v�ܭ�f�;����CژM7n3D5��!�4w��}�(��ey0��	��݉$�[�b	�Uo9��1�w�Y��I�}�sH2��N���c[�E�c�A~s�g}�wq~$�羙W�Oݰ ����*y˿`�Y����`Jgq~���������NC1�\f��)�7�N[�O��[�^籘�38gtə�d��}��Y�r�﫲��x���H$��v �F�d�8 �0��̙����``���L&��{������!���+x&;���1��\��gĂn��A+{ A��=~��s�
v%磃haq�[Ŕ��a��>e��՛z8Οo����$�}���g�-$��x� �;��7�^���x�����ko�G�+O>��1�͹6��:1�y���h\�v�ͻ{ ����HqܧA2�{.�Lu�����s۸����.y�t���!�7Y�a:9��G��z�98��)j�ʑ'i��ݻn�' 8&����;;���^=�cNώ�5�cGu�⚭�p��H�M�����Qp-���ˑX`�l��BR)&,����d�*,�41�B&ך5{�%c׶������j����ʋ�Cz�;@V��|�����'h��W��g\��I*�A$�-�-酡�۴t̐L��o�]�r7a�|x�M����śkn��B�����#Ă���=wd�CD
�܊v��fP*�g�n�H;�'�x��٠�Wf7��~�M����	v�w{'�ۜ�b��^�%y/~�A>�k�A�~�:�R�J��T����4�Q���p�Y-i'��i������ڛ,�u����Bʸ�g:;�����V��<{�>v`]�[J�a
��9��͏%�3�T��R�& EM�P�z�ܲ�ju7z���]c��$��ό6P���K]Ǐ�����@'u�fg%�@�f�ۙ<}���WM͌Ze���d#� f�y����Y����#���@��~]y�ԗ��sO�&3Z�7�{r��h6k�4{_����d�Dci�w�B��=��� �f��"�z5޵����_̮� ��kI��L�	����k�ɟ+{� �9� @$���'�a7"��g.���)���\�we6ۄ���>�gv$J��Z��L>0�/���������pJgq2]tϯ�{<�/��u��NUϰ#꜈	&y�A��#"O��:�!�VԱ��D�vB����eS�z��W�ۀ����P� *�Tν�T�)HI%�����i�bA!��y �`6P��v���KV��@>&���H�i �Q�,��˄����т	��
<�"s�A$�:�2gĒ<Wv��A�&�"���/b#Ee�fg%�o����`$/#��R�����ۧ�۷O������]�:t�Ӟ�g�����{=��?��M�qk2��ٲ�k��ਫ}��>y���^�{�ǰX��Y}���vM��3w�����=sOn.�]�V��Y�Y�i�;N�O�^߯[�s�����緷W�oP�����8�RM�$^��Ez�����yM^�)�n=�{���ݽo�!�49U�ҒAo�}����ySf����)*	���c�΍.��SK=��;<��"�ó��T ��ە�s���Z��r�?o��V-f����B��U�����'��<G�ù3��o��1�1��z���5ó�N[�z6P�z�.��X�f���k@��{7�lP��d=;x�����l}�[	޹�/c�O�վg8���1!�5�.P�:�Ɔ��{��G����p7D��皗@}�k�E�Ө�`ɝ:���`Ҟv��@7���z5�����t�[��[5{�����d~QP=�.yn��F!9`�Ӆ��6=�l}s��@�1�P(�}@���to��<��㾱�4n=�&�L�nm��
|�ˣ��C��|ϻ��� �������U����?c���w���V�c�fM�S�y��/�o�k����=N��o��K4	c��I��͊���N�	����5�%�����ϬZ��u��|M�T~c����W�Ǿ�������7���y�0G�6�S��6��n'�!��j|��y{��֓�}��s7թae*�'����m��{����g��y�����7w���_v
��؞5�Cޫ~�&FS��͸�+Z>��,0>ш�ـ�EH����_� P�lB�AyLQ�c�l�d�E�6Qs�f����+$$�m+V{�.�c
/h�˧9{
��Kd�\�.ښ�YS#�],RF��9�q�z�eP������d��{;��$Ѷх��Q6�ȍ
-6w�L��u���d�]����7k�F�t]I-(V�;�Q��Kl]�Ƚ����#P��T'I���;+C,�R�TJ�oQ��ee<�L;dNĴ	Jw/V�Ńc��s��ّ�m�Ҋ��,�*.�ն0���h�Wk
%mag���59[GV��Q�*�6s����xn�̦��U��(�yj�s�]�E�$StI%h�D��U�V�U�$�T�f��"W�v�߿�ڿ�������6��{�Yk�=r�J�/S���Z�n��Y���ˀv�O���`mڻZU����=׭� ��Z)�r�L���A$��x+s���j1�mM?C�����nf@$�k�q �n�_>������}�o�� ���ӑ[�y];��k^� �VJ1���{��
��S;��w��d�
�؂	�n���@�'�����NH�IW����l
vggL�L�2Uu<��c%4u��h��@�;b	$k�:/+��ӪF���=k\�0��=���� g}s�g���HA�U;�(ޣz.v��y����q���8)�-�L�YdԻ����!}��>'č}��RB�����eJ�ϱ ��cO�

����=���d��3��g���=s�\An�������֯�N���r˪>e��VΩ�yƼ��N�zt�� � �m>�5�S%Gj�6$��O�5l$�C���A��hnc���Wa�-��v�s�~��aֶ�F^w/J�8��M�N�;=vn��KcT�����}*���g�^s+'��m��	�����q�2�R��)���9���E���{j�Q�jPY_}{/�A>��;��nkr�"D
�`A$�?t�$�����\��=t���7��N���)��6[� ��퉴���t�v�$�l�#�}��$�=u+�k�\'N�(n�9hI��1��⁫�x�$[�D�H+�Z��f��zV0��$	m��@�`��f`��N�j�x��$G�nΘ;�;���	y]��ߩ[���(�nj�q���5��`�7��T�:�u��[n3V��4Êƹ��w�������a:�j�ki�\G�*��Է<W!���p�Ƴh$�d2l<(�lw���Gnv�3�>��}�4�'
n�N��;!���n���rMeM�Ũv�nψ��1�іZ�8�l�3������X�[����P����kw�8�7	rٷJl��;;���N�v���Ǟ��^7�:z,ę�K&tu��t�k��1ڋ�g�yƛ7���c{��2ZF2qcM���9#lv�p��1��TB�R�J�P�@UTt鎰7Ňwu��-������$a����E���_6�O���؀^L�{��9':�@$���I"2D&�Rr�Ӧe3�$y� ��MX��(�z��I$|+z6g�<���ws�=V�xŻ�(��#f;Ԛ�p�rBgq�����H��Έ�FsM�?D�������Otd�o��#�|��l
N΋�I3�ɦ�x�3����9�q>$7�����4A���CE�ND��s��=��� �[�i��� �k�1F���&�>]�3> ��� �u��X�F�9�K}bӤ�����HC5�&6;Y�kR��8�k�YS����G�Q�۪1��r���N�n�}���$��͈�����ݝVc�>ʙ�l������������5�����V�i{o9o�꘻�����Mv��:���������,��,S�^u�L�N�LU�-��1U͒���E35�I�4"��k�����d�Pb*�\�r� y���t$O��c|dx���I����,2�]�V�&}1�U�I9d��2�)���	W��qX��%���x�t��D܈%w\�5瑗Ŝ8Eܐ��U.��Z��,��cN�r��]�fޠ�d0'�א O��8�zK�V͓g�1��EDD}�Z�N΋�I3�
]Od��ѱ^6�<�Q}����#9��Wv8�I�~��X'D��As�v�6m��ۜ�FIo2�����%�g�/�E�4T*V�oo����ъ߼8����I>�~���x�wȝû`�T��e\ ����L����r�C�.�A%��M���}�y�^����'�/u]--G��A����RAF_|�{�-4���=�7��Iz\�_<��� �qH%�*7n#�-6ږ��My<���F���86ź�#��*��l��Kp���|=�^te�猔���}��i�eq��}ͼ�ǆ���;s�u�y�Fv{�H���$��t]���Sw\󋈈1�!��|HQ�-��$���6��l��[�<[�\A*;&�F�Ƶ}��Zm���eg�5�s�1Vˇk�ȋ������"�&1��Q&��!+f �H.�)3�.��pRz�N�P�u��˰�Q�D�o�>zG
GU�3?qǭx<W�z�v4�$��?d��^ȉ���;m<���]AD�z>�.7&I���i,��N���m�wX%�6/ϙv׭���.�S�o6L�"pQ	�g��35n��n6N����>��l����r�C�:�I[gG���ű�(w��A�W�'�dO�7s���%���ӧI�.�@�t�wm:�b:�Ƽ]�f8�	[r ����+�F�֑lBz�>NU��b�6_w;׌���W���ׁ���������6�Ov.�c}��=@�W$�R���n03Z$�G{�g&|b:�H�L�fh�w��< 
��'�e��X��D�Ge��Ē
kȀ@+o�@8�ӎϫߋ�w��\i�Թ�d��F����g�2�� �tF�/G#!H��GD!�L-�DlP>}��y&߯xg��=�g~�Է�YS�>�m�"��ē����&g�4�� �xq#�LC�tY �l�J����ѕ�GS^^����,�8N���M �J�ǂ	�6�8pv�D��m}�_@�K��jL\0)�-29�Xa���E�jV����HY�$�����v-�<�6`�b�d��Ӥ�y�gK�$k�v$�������-	Syx�st�� /p�]��qK�$�0��jj��w������ӚǇ�����yo����={�7b����y��)V�x:i�Ox�4�A��F1�� �� ��ug@� ��6�m�Q���Xu�;�m��y�
s�ٮ�s������g�hy�n��v�<�vc�=���Rj�y�Ϡw����OGrÃ�d�g<��8��(�&^ӻZ��۶�9��Σ���縔��q��uՅ$ݺ�T�]ˮ�s�3�������RݟV\�m��v�q���Į:��yxh݈�W�
�w���,5ۤ��6�㷶kn���v���Uu��p*9%���S�^�y'���fh��� @>*�$�wzvd�|;2�֚w]\�3s� �|��<^us3�໒���]��WQ!=��}���0I%]�� 3�vd���9uF���&�l���-3�'����a�w]Κi��s'l�t�G�_�G=��7���l� _���w�zc�+u��x-����z������Ă|wnv$�A��̞����D�ɞ� �F8�k�6;�
wE�@��~�� �m���p��M4�O⼽�"$	��ِw�w�0���Ӭ�2��"��2�����n4)Q�Z��"YHD�F:L11\�Ӝ�ܺNw�-�o$�Wѱ$O7tA�nֈ�\f%�H��Ș�� W��%�3'I��2ۭ;}�崌Խ;��B�����G��LS��c���3~��5z#=sDl�]��'�_o�@�~tm@h��P��X�I�3� �oeC�yy띙�$�n�i�������mKD�;(��6��=�kM?��w��i��p~�	�5W�]�A'��+6z����~1���s��a�KM�W�x9VҤy�*	1Q{��>�y�"��Vfҳ��[$5>��!y�[��`B���w��Þ�L�?n���f�鲟��H.���D�v@�f��,s�TL����em4��Ӓ�a��@���l6|�ٲ�[Inݸ��3Ʈ�N!�,�%������X�r�9n���	6��#�W�n{�96�;45�L��G�߶ �ڔk$�ܺNw�U�:�	�ۆς��f4�6ב�2	n� w��l������#��d�N��5P,��W��$
���_�ʿc�~{��]�����V���(�X���3��n�6�n6����v-:5��2�)2:2rH��f��TD�IS��m���2��������>��V&���轚M��K��]u�^A4MǠ��= ;�6r�"i�H\���"etz'�80��Ӣ��L�4�ۉ��s�6'�DL��	G>��J��	���闟���7}�yù=�k���`��6VP��c��u��Xjv ʢ��� �b�!
���s�N�P���ޚ�~��n���mލ�.'6�u��ϙb. ��E���^FcJgE�L�9i�~�� �y�k��Uv�	 �.���}X�y�||�����N._Nj� d��7���u��� ���'żP9]�\x���=��C_l$�q�$��XnvI1d�3@�,�յ�D�5E���/b�A�llI�${�=j��Z�P{���i.9CQzv��n�?b��8v��Ӎ��ݤ�l��K(�&ꎢ�I�v�����-��	QUl�Ed*��*��V=xP���,{���}�l��0m kX����6ݗ��G�����	ly�O��9A |H��DZ�����T
�RJ!;;p��mZ�teN���lS��d�*#���cL[ǝ�m��B�fx)�߁$����=��y��� �=o\�)Ss�"��J�<�+8�'N� پ�� /%[�-m�ק�y��	w3�G�+{��.�{�7��Ja����:�S;2E;��}��R��A>$_F?U��9fA�
tg��\n�q�i�3��2AF�w���Ӎ�24�ˁ ��w���nr�T�����woH�x�lvI�2t]����	_[�x���33xL�]L�	+� G�k/�}?��/�#�PQEq� � �����?�¢��T   �x��OG�(a	QfY�e�QfY�e�QfY	QfY�aE�fY�eE�fXb`E�QfPY�Ve�QfY�V`E�a�Y�`E�QfPY�Ve�AfTY�aQ�Y��Y��Y����Hi��Y��Y��Y����	I����Y����Y���Y��I������Y��fV`fRefRaf`fVe!���I������Y��Hz�ȊFBefRefRa	����I��Y��I��I��I��Y��aI��I��I��Y��Y��Xde&afRefefR`f���I������Y��A&�I������I��HeefRef`fVe&Ve&����&afefRea�	��Qa�P�� C 	
�2"�u �� �UXdU�P@d 9���� !� ��
�0�� C"p %��ʀC
�0 ȀC (0 Ȁq�� �P@e@!�@�Pa !��p0 �. �X` !� �UX`@!� �D a 8��  C(.\��8�S,2��(,0
�(,0�Èp�*,��2���
,�+2�̠� ���=����h !B�"L� �D/��=�����yT�����?�����Xp���h���2c��?�?W_�{��PQE~�������T^|HEE�����|@�������s��h~�
(����"�A�X�:�����́����?U���QDAbTA�PB�B�� 
` &UY@BYaHP	 �VD  $P$@$T! %H@� �$@!	@		�Q�$���pE��O���O�*��Р�@�P �%���?o�����P{��� �����q(�������������pg�?�������ݤ����}B
(���C�O�׏�<�Q_���+�?bi�����N^~A�	QE�~�ܘ���C���y����I���&N'����� r
(��>�����D?�9QE~���}��ó��|����u����	?�����c���Q]G�G�������W���&���:
L/�?zp} �'��~G��v|������"
(�)�T����&?`d��8���}p���@ ���9`�|s�U W�^�9��!����PVI��Oq���6kV` ����������                  }                   � �      ��  �4  @� (�    �� (     
 
PӾ                                     @         R�W�fz:�rj�f�ڊ � �
�1��U� j*ɥQ�� v����`�y��    �����!3j�)� ��)Ɉ
d5T��P�.YW,(z1� ΅
��YE�^1���H0j�����i@P� � �H� z	         @ 12��OA�y��СNl���)�x =(S6̑HW3@\��W,
R�YW-J:� ]B�*f��K��PPB��  �^g����h�� TS��4U�Ӑ���zֵ� �ڢ��z����3G�T�4:� 	  x   <         pٞ�m4g3]e�i���3��Mjm� ,���4ܺ�����vngN�Y� �;e���4�rs@(  <   ;��:ͭ�:�ԍ� ���al9�DE-����3mN��\ 4v����U.wtl��ͮde�;�m%Xh  �  ��      ���.\��5�7)q��;tQ\nv�6p .(��]V�q۪Mf�g@Dc��ґ� mUnq݂�r��
@�  ��7.��s;m� �Q���jk5���K(�ݴ,�sk�-5�� X����S4���Cb��H�M4�A�� �         nU�\�\�X��ʮ�F���`ڶ��t% *�aswR�ն�k����scs5�*� �S�q7V�s�@�JR�� = s��T�Y+�� ��ɕ2��fh����7 �:4�ʨ��]nf�Q,Ύ��O&�����4?�i�)T�1 ���=��  =��FjRP# #T��i2�* �M$ML�*S@ �$
�)����7A[`yD�Zd$N���$���0$�	&��BC��IO�H@��B�$�x9��w�����ZɪO�3Sx��T������i�V��@�@mm���v�`��u�#94i:���Ǐ-��2�;�9��7}�敊�������|w�C���N��zw.��A�ښX��I�s�ḕ#�jYO.u��7ON�5�9�E��h����!�n^�W`���;�Py�R�H���{��[�b��T5���K �+��J����WKyuئ=D3�h	���Zj[�)���ε������q�p�wW�ɵ��e��w$�f��m�NŻ�9.+Fոw;{�p*�f^Xaj��f�ˈ��L3@}q�͸�M"Gս�՟�;Wb�7'z�N{�vg�S�����^�n�b���Pk�5rA��n��ӝ�oJ��E��ifv-I�*��$Nb2��u�7w�Y4jG@yr�wV��ݱ�zV� �;w�}v�]����s�l�2���f����i�#Ss^7NU�jx����|��V"=���&��ët�����n,	5�t�a��	85Mۯ��y�%�an��[;�ww�}�~O���šW�:���j���K�G+��x�Űݚ^L]�A'J�HT�Q�	�F�]ެeg���窪M|�B$p0�k��۝��v����p�Ҙ���
�e��e�@�w�i՝ߞ�OV��^5�T�֢C$6� ��k������nC-�$.��o��1�c�{��.A�9bWww7����띥�+d��]�gQ߁�&ɋ�ï ��6*�*����#�	C{-���ب�i�����bHL=�bGSx	�Ճ��ƌ��@��V�	jc.�v�u��{��B9@z�0^����8p97ɽy���R�zq�R�-p-Y�XfHuiܪXV���w�$:�ck#lt{'o�3H/#=�,j�-��٪���A8#\h�y�^�[��D���\�0�T���v���� u�e4ю\��[On�W����"N���zgc��J`��l�g]p�2�ӝ�stf��%�� cv�98�y��)��M����>U*�Oq��]4n�0H�q��^�]j"��b1F�>�M�7;�aa
����X�ee{p�sΘ�O9���C�l�ӳ\�kӽ�k�F`���{����!�(�8�i=�R�.�LR�7�Mc�;�:4����c1�v S�6�5���1��5u!^�U�1����-3��e�b�h��rb+9ז���(���S�tJO�.���·�7t��p�݁�;���_wu���軲-�6�P��{�-~��us�1p^�$^ڝa��"��lQ�D<�ny#����(_(@�_T�<���t'��#f�<C����f�3.<��$żs�6�Jն�ҕۮ�S�n��5v��'�;�<���'j��xs����qnu��܏����&r]�ڸZ�����.�Z�Q������[��J����,n��r���9{9֍��&mC���d�냞��r��T�L4�;ENdD4b��=�q��.v�	�zi�NM�\�إ/uIύȋ����9W��eaW�!5q�S]|����|��̑J��D�N@�b����ם/oT�Ǜ�4�����|e�X��b�ݴe�,F�Ω�:-���a�*�&��0+��<X�0<����aMt�]��d�5�3�C�6\ֱ��\+_W�"�0&�b�Q}�v���z�LҚ!�ݓtץD�֋������J��b���hL5���P�idќ�F\\u�tv���׳��(�֋�т_ʋa�]��M��w��ŅwYT���H>�7f%�9^A���;��1��Iwq=�)�`5J��fot��y���F����f�/-bĒ��_m��[�T���ҝw8k���#���vG���:�ȧ���䶃����=�w!-�G�\�����gCp�Q����Oy����tq�O����Ɇvt��7']�8k����;�odҠb�>�����]nZ��ri��\7��ϩ����c��(�ؒI�ݜ6B��o~YѸ�Ɩ���k�ح	@���6�*��7�,Zvi������O[�q�Upp�Ov�$P�Qfn�ݠ�G���J��n��-�Փ 2��Zꉋ:�O]sz�y�11;�&r��7�n,���X��0��[��N?���INYޥ�?@�vďMi�dZE\ڍ�C�;�8q��]ŀ��4�7^��{1�\�Dag��q�	p�w*ۓ{��RUͤgaJ��iCn��^E�P���7"��.4���/0r�<o�9���;���UXUGan��K�b��5Z`Vj�1��z��ĽK�]z�{��� ���_�N��fp��gP��qw2|�Y�ܚ��j7���s��憞�m]��R��$rS�֜�@�0hˎ�ޑ���"����2���Wk����!e-]M��k M�m�r=~)��]�A�{���(����FS�d���/.�% ��T�9��h&�!�"d�fZӊpW�ܣ�s0i;�U!��՜wۨ~[�Zi#Ϊ�+mmȸ,t��40�f�M�u�X�4�h�}���V������t��]��K'M�w��%��Nv�%�������������8��n���GX󵄷��\�eV�l������wDJ��q�f��ٳn�G<n �~u����^,85oF��W���F��p�k���.E�O.�y�(p^Ma�ќ�c�c;��ۀ�B�ݣ��r���en�r���xA3$\m��J��Ƅ°���iJdѺU���NҔon���U5�1n4�ɗ6U��[�:���f��ȃݻ�\'8��d�����õ�uY���p����Z�y<�^��?F�4�1s���H	GK�-�n-y�M����93_�B�V�9������LO��F�Ov�����>ݷ�E����4z�0���y�������C�m[�!��1L��Mc�Ni�Y�v��(t�U���#9��ug��P�ōũX[9�+��:�[�{�X�G��Y��z��osڦun-��x:^��H��*R�X��t>���c��G���,.GtG@���=����Ό�T�^����ҍ�l;�{{Xbt�<5�2�c�:�����v�1]7��'LX�u��%�f@�/�&UE�,c[˖5GA���D��斮A(�C��*(�(���(�E��4�yݜ ���X�1d��2�z�7o��"�{�����{�����iξו�+��*`�*�$�dG-4m���9"k�6dT-i ���p<�6v�r��^��j�?�xM�)x���� �h��B\��v�9q�I���u���nM"���&��ޏ����h ��rU܀�/JS$fl;K:ևZdw���l�k��%�����#2�dnv��=Qs����B��^Qh��Ž�ڊ�Z��V�A{���k�ygn:\9s����紓@��x!�%�aa=95��1��)m��&�3v��[w|�ÏsbR���,k�9c{%�.��y���	[�x���٣�$/T���c�;7�4�,,���5ל���/��,� <m�I�X���h��M��E C�hn����[��0��hݸ�]�}�ܧa����mkT�G(�v�f�Q���{g�ꅎ%Cv�gn�`�t\�g�����E��NX�M�Fg����Y�ZGu�)���dn��Zmb:.�$�*��Xx9���!���%e��QA�Gf΋7�y�F���ݜ�º���\8��Ғ#��H8ov,2�"�����<�mż�`	q��c�N٤Y�������`4��f�t��r��:`�Y��`o�c�u/��4n�{n��Cӝ��t1�����i/9�ڟ+x�2aL�-�IC��h��ۺ�jMf���Ԏ���.0�n��ݑ Bw{��/d,퀴�o�6��:2&8A_��=��ۧ��1��9l�`kZ�LjM�m�t�0�� n������+�� U!�Z��І����SA�w{d*�e���B8���Q;Û�P-Ju��+V��oQ��"�<��]�������%19���92.?�nR�w�}��2��"r~v��fE{�6P�B]�_rgD̴��$@�iks�1��&�]��w&���>qm��3�d=�giz	і����%Ϛ�ׁ��jx(.��4��X�l�~х�%7l�J��wc��`�osg1���*2��q�o]�rn>FcỬ`Xx'����iܟ��@d� %��2�һ�6�Y�:n�9?�^�^qü��ū�[�Gg�kW��B�э�0WRW.��)�3�,�u�b�zrm�-��y�f��/!|C����grJ�D�&��!����vQ=�f��t�Mu��_>M�!�Q�3fL�tx�������0��3] ��h�Mm�������x���,�ӳ�uv���Bz����7PS��S&���Q��M��(������Q�;�"���ǲ���N�TW.;gg>4�z��nI�#Лa�����A�-dĎ۶^��VT3�g8J���Dp��Y�.[أ��X���%�:�7��q�S����s�9ݓ���ƻ�ΐ!�j�V��6����whC�e}�=:�`Dnx��Kq�
G��7.sǿ�r$'!,@(.$�Y����˻�٬��"�β�6�����vr�;�y�ٗ�V�U����o���2����2����}2)[���q�p\y'e?�}ǉG[��[Xި#Yh�R�c�T�=�Q	����'d�.d���ɜ����h;���+4e��$��'�=� S��9��v����*4��(��2���s��Vv�wR��w\�u�){��L^�ɨ�3p����9��*��e��C[����oQ^�,�3w��ڏZ���v0;pv+H�V����M�T�#p����i��1��\�d��Xo`O�=�cn��ί�U���7��Z�[��(���f$uG��x�
2��Q��ʻ�+.��`x��4gU�c8�5l.e�ݚ m����2�/RòsWIhr�o�7M����)���n[oe�r��ӝ��0Y��1P0�FI�2e�?�[��y�h�x7;�b��0��R�{V-0�b�Dˢ���X�Wf�����h_ƌ䍘�	�=�^����l���ЪoL=��wZ��r��*��tD>���|�d���v�T��S�^���`@�:���L{H���c�+8�9F��ۜ����i���'4�z�А��	ܱ�1HwI]�#��BgW��hy�c,f������:�&H\U�z���4h*�F��:�ڳ��׸����객�E�.c��p�qh�A�Q�(�ی��x���D=1U7m�]Vk�'3��志`�ª�wn��*��4�i�ɖӌ#�"��wR�w;K3�q��#X�=&9���a]My�����0�FC�T���!�Z�������1,�O1H<�+��ׯdVq�F=d�V��aȴq�I1Jս��G���m��6��KIqn�3����'q{��.��;8)2蜳��{��rs��&��.'���ݏp�M���'��o�wW���᪨��}����8s��٣�׻f7^�ZxK	�]��g>��[҇���Bor$��p���y�;���rHa{4�nu
-s������m�'8�^�.oN�D�j.-;��_E�x2���`6��n�NZŒ<"S�=�gN�Y仩� �Pe��ot��, ۂSQ���ˁ���=�d$��Ͱ;�15ߦt�3�M��;����9ѭ������}O�W�q���?jg�'�M���r]��s�����[�zmm�,���5�guC:n��5����9��g/:��F:]Ngd� ]m�^��Kxn�%�5Y�Ux��0VA�]�7GۋB�s�	��/]՚:a�F�;��%��:�[��j��F%�Nƕ�N�9���)d��D!ㄭ��f����T��e� ����epǇA��D��lś�?U����o�`;J�������e��i����7�Y(K��]��攲$@����Ot���պ��Զ%rދ�-�ѫ��a��.q֬�k d۷s�՛×	ݸ��'i��.�Ѽ�������r捁���ن����w]���(�ћ&.�;�sz\}��@�0bɵ]{z��7kº���aӝ\VK^ӫ�c�9��s8�ܸ2f9��aMi[��̵�[��,�/�S���h-��`� �@���\�Zņf�('* ����[����a%�+'曝��Ї��{y�4���3w�O�n�?Vf�ĸ�V��m� Ð�F���fo⪕�������.�"�}sL<�K\d/�կ��j�B�l�cyHO.��nu`�9��ho�*�-��w��w��? �\���<FU��g!~"^hi#G"��j��6Z�ѵ�/wnA5�2u��m�te�P Y��wi���	��5�̉�Á˛����l1z(�Z��a/��Ρ��m���qcW���ĉ�:��Y�q�
�<�be,Č���ew��Ͻ��H`H�$�XB(E��P��BH�HH,�
�$**I �HVBIR�I$P�V* �IBT �
A`@@���H��� � , ,�"�`I$�� ,�B(���P�,�
�T`H
B+	
�)%d�*B@ 
�d�@��+$��I%a!"�"�$�!���!!X �d��H
YH,$�T�aEY �Y$ �B@XB
HAH �d	"���I�YB�J����a!"���	`AH�B�@�$�@�B
B�a� � P�`XH(��� )I�I @$$?Đ��$��߹�i޷�;������D���Q�S�S;=��]�����4#���:nAi���1�6r�OYXiѾ�x�3Pͻ'�I���<Y��򻿎޶.Y���Gn�'���M����0�_�k7=�@�2I�WOk��X|�m�z�|D���{�����_��'�{nQkbS�n7���af�>��a�Ґ����ok�su6���pU���>�K,�@Nŭ��R�v��˼��~�N{�=Og`����0�������%��q��H���vp�;��=�:�0��.-:�;�o��}�uyII���t��?�\����*ni���=��{�Gӟ��v��8|��[�P�ōN-5���u}�L���{xo������(�<�3&���w�K^�A����06��6�#u�3v�����`5�G�>�
a����E�,��T�(16+�7QE-н}x�>���j�g&�_.C7f\��vǩ0��Z��L��,;����MI���z�#�|?�:'���k��W�y6�x"v�����=�e�o�rU=�c"z;'�Ɯȸ��44�c���G���t���@ƽO5����w�#s[Gz�]�tO�w
�3ߕ�c��ʯ7�N�dkݤ"���˧g�����c�׶���u${+Í㉬�ti�]���U�+�3�&��{s�җ�N�Gnm^��H���i���z9�Uو������[�pԸ�w�'��#�w���$_���Y��w���l����&��<v�s�/��_���,���$����~�7up����un�>�8�����蟡��9���~�nD�04{�h4y��vC���j��6a��Q��}���n_'�-w�y�2�x�IH������z�16��dV����w���v���~�'h�s����(9`m�j�W��.�'����Z�M��̾�ܙ�ˤ�9T9�O^{:�9Sp��B�� {|=ŋ\��w�u����F^�����5
�_wf������\��ʔ�n�"������,�r�L;�yw@�'�a�]+}�z�Ԛ����o����}�����6�h���R�,���zԻR���u#Ѿ!��A��?	��5f��^!�0��w��f˸frX�~����y��[�l�݌�2�ٛ�픰��{��X9{t���f��Lב�y���	�>Y�U�cDL/�a�[���I��n�\��2i��1�xt�zq�Un�}�����^�sԗ��������7�#U�3!c�[��a���eX�U��2"6�r�h����7�;K	���U��-+nD޾�����#����
�A��[٩n�P�e� �;�����1x2S��жv�`�po�޶#�1@=�φ��zf�𰊂��{.Uf�r���K��˸$�&���O��������t�S��"zi���݌�����)�{l0�{ޣ*H�Fɾ��������;=���3���MC��W@?��of�v�0�k緸���I�Θ�����7'��]�wb������YÂك���$(�*{�k��ɜb�^�tk@�@3����j���^�.�`N9�=�w��?1�	�wG�]�I�ǀo�!��n;��;����gm�ۖ{�-���)s�P����)���[�!��x>����r�}���W��=Ķ_�/nm��"r-���sd��Æ��{5���<���<ҽ��gp,)��>�9v�X��
�]E���{�q�(I>^�N�i�sD>��������Y��vMh��g07d�� ���n�/�%���}`I�{=��c+���_�4]��wu7����O����ء��˽^p ��{V��y\YYw���o�j�d����̚��}�gW��>�����PDM�E���λ�T�^�N{�_�z���j�g}��{�R�j'4=���tE�I�w���:�,,����>��׷���^�=��}�7ˍW��0$zm��J��ɇ=r1ge���te���o����I}�2y������F�CS�I�1����|���ON9�F���ח���^-���֛��Ëe}����o���oq����r�=��/qM����K�4/Tf�4�{[d�>������qj>վ�9;�	E�����f�d7<�þ��]6b%��lcc���K�u��F�6���B�ݩ�qm('��&�H���RM��n��Z{�y��S5�ݩz7+G�^�]�1�Ǟq}���0��v��,L�ŷ�c*WΣ�c���޵������mK��{:?%��{$]wX
��������ga%����� �z��lW�J��N{ϩ��s_��!Td)=s�پ�sFx�}�e��̚V{��.D֧��5�{��C��8%��l�×�����|��գ=�6���͛�g�kv�s�jzt���5f�η�������|��y:�x���q�A���{bY������Îm�{�pZ�tz��3Op��v�8@�r??HĹ��JP�o$q�M����;K��D5��8F���x���@�<��V�p������n���s�d����Κ�����ͷ�jn��Ç�~�b��cܦȳ�����������e���x�=#���^zs39��I�"�}|�X����s�=���4�1H��^��j�ȼ���Ra�[V����x5v��2x��#��NIj�dJhE1}��=�=6Y�>����@���p�L��LO�3ϖ��1{ؽ]n&�:��'�LH��óÉO��x���7�LK&�}�Ow��qxY �ѱ����KΤl]�OM����w��Xݓ����Z��z���`�-��ỗU����d�Ů��=�tȆoOj�(v���0<Q�y����gB�i�H#3�K�!�Na���y���<�Ӏv��]����LOe�M��x�:��4���K��W�����=(��'��.�;���	���=��x?$q䜜8��r���o�:�bH��NG��_�ܙ�gd9����{���8��1/F3�n��۞�ӴL�W�_���{�8��]������Ÿ,G4��}����Ľ\x�o�t���#X�c�pʛ]����������싼��P��5���n���|Lf9���!�D�p�7ղ|:�fo ���{Q�'�#}�����Mjjz��'f�:y�:=+ɨ��� ����g�m��+�ǽ�r0�u�,�9���r:=l�.vn�޾2U�����We���g�x3�&��<�Է��p��S^=�=2[���2bߏ��W��7��}��g��#��a�IS�íMu�_�uz��s����������^t����/mqJ��??c����Ӫ�F�&^�e	�#3onLzPŪc�u�`B�ɫ���0�l��"椮��q��?��yg�̵x������w�����&���<p�x`X�S���Z{�[��A�0��3����.������=�����[+�^���o�\���<�AI�U���&����W���C��\�m��ݴ�w7\��6׽�h?��^��c$��\=�m�ջ�|���v�4���)��V8K�gnZ�W�����3�ny`�wWb�g�nyl�ܾͧn�����;hu�����|7J���8〜�{��;�����w��)�-�jƊ��)��w�\<�2���q��j�3}�f\�/���xp��ż�/s��e;�J���"0�7���O_Ox"��9���:�t=�|v�{�vL����o��S]����u�IH�h�}����D�����>ҖC/��f{�h��@�n�(E�o�VxkڇQ|{֦/��Ҍ�۝���<l\ꫥ�ԝ �:=��k=b}�s?�x.�BQ;z��E��t3מ�x_31ޏ���ϔ����$q����Y���ǂɔij��>���u�6��sE�;|�3��%��Ï%ۨgr����o.���vrB��U��~k��ۜt����_;��w�jՔp�:e��7�.��������������w׷#މ92f��2�,s�s�q�9��y ����{:{b�NM��wM<,�sog�q�p�Cso����jl���s���������ե3�\y��<�}�7��o����9̓'�K�:����P٨q@�m��v���O@�cF�>�����uy>3���F�^I� g�N~>�AOwI�Bw=��F���C�do���o)���j��'TF�.�[�{Y'^vm�;V�o_7W�=2��޿�x���8޻��y�gK��������� {�\�n�Qk-f�Y;<��*L�׆C鞜�����<5w�W%-��mf�nީ��[5}�����5�b�5OC�ϊ�y@]"lq=���ͳ�s���Y��=�Ō���z���֪}<�xv��/� ����tw�2�_Z6o��K��֟c�Id<0��j�6��}��l�$�̂&���RVE�Π&���Ý�;�eJu����aXg��ms�E�W+W�~����m��19�!��޾�=�pf��>��u�4����P���܍���CqL���;z.#�{jG%LaEmj���z�ݾw�̯�/�v�7�W���K�e����A%�.wNV�i[!ѿ�g��`g�/˹�=�S�n��9��VkcK��zl�=G�{O���vW_u��{}��&��lɖ=�eJ7����חy���T�y�N�X��g�e�7g��xO����HL��v�xx��Z��x�o��)���+\��I3����㯫�p?N��y'` �w�����/x�N`�<F�O}��U=W��V��./u�}K��g��ۀGu�ko|�+G1�*vo��8��]8�B���[f�D�7(n�ZV��$�x��G��{����vr�<=��s�K�܏y��y�-9Y�'��֠f�>���S(�{*]��ʽ��;׍�%F�B�֍=�u��x��615AY"��0�۫4���pѝ�{����~^�ɳܦ0��\�0��1�s�3�������[�c}�J����)�{��-��]��w<*���2��u���8<=?zMyc���������o5�\��N<V#�V0ߠ�׹b97�����ŧ��e����{=������{;�S�!�c7^�s��=:�;��s��{p�u���! ����/Ow���c�!�N.�_��]���m��;����Y��,�#��X�����Y�F�bن'���%Z.���%8ti���d��/y��O���C(�u!�5���r7Xz���,#��B��wc�ř�ʭ�v�=�8)3^��=��*�"�O�	��䟞l����_5����޺��%���fٺ�>�7G �y�x�f�Ť� :��V��{eQ�ɟ]�Z��xx����}ӽ Ɨt���������u�T��x1��df�����sT;�Y&�0 =/�o�bO��ɻ
s7=� t+��0�����׽�e�=��+����1�������.�Ƕ����9�=�d(���V����Q�f��S~��ا^7�o���Zr��d�-�w{;������7���6+<�Ո�ە����]�\k��lA=�m여��8�?-�L������n#��]�zX����('�]yС�^���{ؽ|O�?n[��r���vpW|=�I!W�HW��������ۂJ���V�������������Ň�Kn�>�wc�Lkd7h����GH����p'eZ�`u^�A���k��;+�����e�����[�����`?{�5�z;�{p��uH�V�𺷍ef��=ܸ���E���d�ӺD���vM}n�vK��E�^����r�Җ֕x���k�6P���c<[K����"�
����2A���nX4#��,@���'���Ʒ�m����i�ǒ�\���9��t��V�-ܡ�зظ(�<;j�:M��V��՛ow���N�=�==x�9=$�q�9�ΖN��٣=�M�C��
��޾Zvh���S�E�/E��sWX``kk/��o���b�xOE۶W��
�к!z��/�'����M��ȼGMC��>׫޳���g3��;T���;�{p�Ϋ���y��5:v͈�ݶ��֎�3��)綠0�p�+�/�>�+�p3�_�s�/�v��9�y?ۑHoyf��7&�S�_~��؄w���&-�X}"�8�3<}��xبԨK��'��K�~O{�c��f��G�zb<g�P{9g��!B�rNΫ�1�n������_��w���E��=�FDcE����᎜l{��U���f{.�[$g�D۩�L�5�׿�oJ���o�����{���f�w�y��xsc�G�g~(s�pG��bd�������_��/6��Cp�����MG=����{ܺ��-��P�m`mi� r��Ӻ�:��E���x�w�x>����<�����c�2���7�Wq�܇���\���睠�yg~?�49��o�;yC5h����d�
#���_����)��{�E�>SMuj��������{��{}�@���^wr��L��D� /x���+_�%F8�o]e��N�|�֭째7�X���5�O����ij;�[�)��7��-���E�śv�.�5�ͺv*�����]���D�zxM�e����T����fm�)d�<��΢�f��U���S�Qk����d�����||=�����^����z��3�R�ɾ�c�軹�O�t���U�=��^�m6c�*Ss���5a��:��<}}���~NK䯮����q�n�z/mތrwn��
�"��z�nY�}��|�.�>���^B������ �wU����	;z3Ӕ@����������$�	&I.s7����9�'mm�q�;���qn�ъ0<Ʋz�`�w'�)r7W>��m��gl��p�O,s���:ѵC\�fǐ6�mכZɮEIa�t��-��۫h͛��kn�����h�^y{a���7I�l\���k�r���p��6:�G;X[���:�ٸ�Ԃ4�|mSn��o<�ǉ���ս����ٶ�x�-�g[�;�z6S�iBup��5�՘���&[t����i��/x:�ngv�u�u��[Ÿ6�k�p�y�n��u��ю0�nk݃^m}s��;n=�\\ݗ�73�q�h��m�v�n�[N��>5\�7��X]�4ݺ�F���ҧDw������:��t��{r]����]0�[��ϳ��8-��vGn��z��w��\�+����n�q':�b�#�s�����l�y�Kی�N�Ҽ�x�W5�$m3�Z�5K�w�=��xMu=������c����A��\���k�<J�um[M��T�M=m��<���Otb�y�����Ƕ;-������1kg�K�Of��s�{P��V�����W]�Wֻo\M�����h�<�VM�v����㫫c�rq�gq۲��.�As<q�[�m�D�'��2���ܺ�ۨ^ ��&�B-�gQ��-rs�ڌ���n�����۷��`�E�k���.C6��=3q�;��̝��v)�c�^Mv;O	t�-ȭ�t�S�n��^�w.ݠ��b���Vpn�Z���b��aln�`+�=��<{B
=�6k�
%����v�9�����
��v����S��+�fn���6�v�e{��v��-ӣnvxn���B�^�I�;��4�p<svU��::�ܜּ�w;�Ӫ�2���v�-<󠰅ۇ�=G��ǌu(;��v�2g�6��ݗf#��r��\u��M���kDr�Xuvs�n�87��V,�vK:ļ^�#�ʺ������-S��w<��1�8�=��f2��]��`���ק��N=v[�g�5���f�9w��u�������sY�.���܆��}��0!���'2�5=�r�����;,��z�m��sn�X�.f4=��G�t���f�c/#���+����&�	۞�r��q�,�sm ��'r��Γ�:7��8�y���z���s=�#� W�<�k���u9���[nO-]�:ಘ�� �<�
ݮ�t=��st�MtS�m�J�2m��؎:U�6���ٲ�����|7�ux�Ug{h��nS7g���ǻ\�1�8}/<2�	q[,�G:�v��[�w<��qۣ�����=�c�o)�N��3�q�����9�4�ǚ9\8�دO.�y���',tL�j�]�sz��]�7;]m����T��윽��v�SY��:�9�ݳ�H^�`�'P+����4�<iT�u;N�x��pX�S��#8���m)��}L���Ob������s��pi���6�U�bC]p���n@˵ځ�	���a���g��ΰ��G[�\�8�t{lV�k��7U��m.ѻ9�EmF�t3ʏ#���vUk�`6��x{c�;�\�RKHU���Յ��ƶtF|��\���7n�˄�<�s�(tnY����Ƹ�uW�3�I�{�	n�n�g�'.Nݻ�[9���Fd�!�#�Y϶�wf�v���tnl�uǷO G��[tc�S%�ñ������m��јr���n�W����M����7]db��d�47:�t�7=s�p������W#�(����^��0"�^:���|mٹ��f�Mp��8K��Ӹ�nk�wF�d,��g��8ۖ��p�g-[ŷrV�2t�d�vtj��1ϰC��'��ۊsn9d7nv���[�9�8&�\q�.0��x��EW�0�s�6�ӭ]�:��wf�weq��V�ny�ݛ��ݺU��*f�gp.��ϭ�n��7m����6h�����F�]��9�)v��.�ԇ���ͬ�W\�tu���:8��6Ɨ���@�,���{nF����q=��ք�V��;]���^�r�W'��3]��c]̑�{[�������Uh�m�enV�Q���V�a��n:��Qc��x��ݖ�睂�`��mUú�wN������5�7u�kv��ҺvH��rb�+�{/W��1�8^s��r셱��G'���q�l��5ͭ8�K�n��p`;L�V%<���E�1u��ۮ9�^���ضz������f�v��y9�xvN����lX]��^���ӻ�^\u&�.�f{\Ns��pt�f�;q��u��e=�-�Ny�����é5ɷ<�pv���k\�GZ�/Ǝ �eϡ���="y��a���i�Q�y)���xx,vT  �"�{$s'i�s����;P�<n5�F�!뇞y�Z^m����f�K����s���q�
8{v[�s��b�5��3�k�d�+l+�1�l��ќ�;�<k���S�g����\Q̌��.P;Ű&+��=tۍ�N��;m��n�Ck�ջ:8^#���s�4rk�u��t\\�{=�+�c�,*�C�v1���8;e힌���h��퍮1:��[g��)rk���^x�� ��wv3�K�3�:{=�{nt��e��ݹƱ;l<g\����9�K���}�vw]t뗃Σ�C*&���N죳��v�x8u�����;���Ɇ��[���;7vN�m��H���؆�kcM!����8���TƼmۇU@�ܽ��:�6݂d����<.7
u�}<��t�S��\s&]�n�hS�v^S�����Q���mӢ{$+��ɷnULi�N1ˮ�[(W���7��C�;D$s�Ӯ�22K�E�@�%l�o/gf����5�;u����3������7d��d�O+q���^�T�x��mۍt��ͷ �g�tܻfɋN���|
N� ��9�v�1	�k�,����5.�\��ۺ��ݭ�i��j7����cZ��f��L�V|v�
[f˝�hT7����rqm�&�vݫ�60<auvM��a4Zi�N�����:���l�\��u�8���\\�6b�sīف�d����p;Z.�0�+�՜ɰ�Km��z�qvЋ��ف�R�v��C�y�7r���X=���%ą���V��+�7ʦ8�6�۞���6:F��;�,�8�˲f�[��S��+)��6{�C�CqV#��ݹ��OT�;7��]u���7�Z��m`��v8�dv����nĬ{;)˽X�\�؁�0�s�v����R�Lgv�
�	�-���q�\��5��tn7�H4g�b��ܽ[n����t'n_%m�X���9�t�Z���\ufGt�Q�Z7 ������Ѳn��c�Z�U��hM�:�.��= �����W9y'�����u���;rz.{C���X��'V"w;v��Ө7�5^�u�Q��Π�p<�x��}��-n7gC����gr�rs�]3�Y��f�D���;�6
��Gf�rc���6ڣ�a��A�G-�i�nз&�t�ܷx�nm��y[��\�$A+vt<w9�={:.�G�ٷ�x�ݹlYz�u՘ձ��x����Þ6ƶ*v�`喦�+�8��@��t��'h��=�uڨ:�	�8�s�n�d^��7O(�9=<�1ͷK��tv�����Kq{n;�v뜾�)v;s�onk��jݞ���I6۞|`"^��Zㅹ筵v��u��'c��<�=gm��Wn�J�ӏ768A
�[��սv`�\�����a�ɳ�5��vuax^������+��p7$�m7��(m�,vS�부�nx+>��,��s��oZ�k�Y��v�kC��Uˡb�:����o[N��y��q�u�T5h�\�1���r�Nۜ�6u���s���[�.&�qcȆx�:�#��j���qU�O\E�WQ[klk�k�a���\�Ń�`⣧s�^m�d�"�x��
���R_\u��l{][�v��<g��v<;�m;��c��zJ��a`�nS1��˛����&��	�Mq��F�<�\�����c�W�,ў�ak�����q���嵋u�;l��l��M�c\q����j�ҽ���.�G�u�0q[�\[8�l�&��3�u��b�1�I�xM���N�6뭺����v�Ƒ��-��^��Mn�\67n'=!��f���3٫��
���j���a=�p;;��j������h'%�ۧ�r��Ȝ�9"���]���-�Qq�d�ٯdk�y���F��%���ݹ�8n�c<�vیs�3F9:ԕ���aK��\�#gv�8��v�u�u��G"��Z����l.�����8ׅ���g5U\��%�玷f)q���u���'�I�T��θؓ���NA[�η���q�Y�,�k���4�Qku����'=s�<v*z���s�յ�uƍ�v��=s��$�����]�X�Yi�(O#�zܗ��Glu��X�^��؛�꧷���nܰ�)�Ő���,��s�'.�N`��Ԋ��G��W��Yw���6+=���T�]�[p����8�>��۳�6�s>g-�w���y��Kg�E�惈�Q�ه�c�C�W�g����N�6nePT�C	�G]�۰��lj�m��u^�Z�r�!]�����.g�9�ۀ���;��x=�]w#m1�xҷC�g�����]9�7�z<�+�W]�`ިV1 �P���:���7co^����c������Y:ݩ���3bL�b�Ţ��=y�N�j�6�v{f�<s��f�
W�ݍ���=�-���$X��v����̇=�U����y�8�1��z���v3�����7p�:�Fp��&7;{]��3�j��(��T�j��UuNJ�=M�mV����V�Pi�.� 1T��s%V9q�TLj��Tc��h�ҮUŴ�bT���Kl�P�!��b�̲*9Yd���Df\@\X�Q̸"�PU��f\�j�k.*�����cA�[��VХh啔L¢�ib�e�Pb9q�˔*�[QJ��ZfRڹ�pk�"9J��0��n*b�E�2�X���Ujc���T��Y�Q+D�`+Fi����A�Ut�"�b&	m�T�A��mm*��Z�����2�˂��q��EX��J�Le���`�
&\�T��2�*�[LJ21�������+*8���b��Z�i�R�S)m*�e��Z�G)�r�PQE�)�nQ-m�E��Lr�+��R��L˃Z��.a�s,DAQX�iRR�V�ыD̷3#�Tql�W"�-�-J��m�qq-��4QTA�˫4�u�4Tm�*[LLV	+E�W\�j��bQfb⍵���e��0r��i�0�"�_n�+��{��t��n������[q���������jͤ�+����듶�r�\Z��S��m�؎�&O���2������ �<�qB�����
ʧGe]A�R݇�a���q�4{c��T��C�s�:�1�Lz�ģ�����|ۄ�"iַ�Śݽ���xw�����{�uѢx��G+���["v�Z�O��#��㰾��Z�k��f��g[��"��|�8c����֝o���yô���,���v=�mۮt�ۇ���=n�<F�6�-�ۋ܏u��Oj�s��^���H��
�Ս���u�Bv\���ecl�n�ۄ|x{q���띳�� ���u��v��)k��6.I:�csp]�W�����W<�W]��*)����c�ܳ�\a�ƺ3�64�/��pѹ��4]O/k����n��yz5�:�(�sq��/p��;d��I�^1ϐ��S���.��Ѩx�yۇy���/qZ:�ڝ�q����q�;�(��8���wm�����m'\����'���nP��ur��/o=N:�c5�`�7%�7ot�w5ѽ�\��bjޣ�Mɻ��:����;'/������9���>.SuvG���F��8vx\��q�m�Cӻy�Gg����g�`I��+�^x6��rl��x�h��^�mf��9�ܤ]�g�jޚ:L���;�C]���ݶ	�\8v��r��zz�ae^���^���ݸ��M�S���K�m�=�ѹ�nW£:�㮸���<e�k���J��E��8��ŭ��Q����Fk���lPػ�*i��0���%���s\o��<�>����i�/�/�8��k85��.�v���v�k�������mCv\s����ձ�7G�q�૳�,�N+{]�v�n|��1�2�\f�ܚsi�$oa��O4mE׎�nwm�ڼr�cu从����#�xb����8�(��n���]3W3�W�S2�;e]�m����r�L'#���M�ar��9C�kU�n\*bej\3-�)\�ǀ��ey�"���s���<��7h�n�FP�܊pg<���s��*'ga�㘎e�h�Qm��q�0�ULL�l�{v�6˷g<q��û�v�m�{ �l�\<y�㌡�J�VZR�j�c��q��a�����{�U����ձvĜ�͚$�V�&��;�q�mvNFuwU|:�kN��I�>�`�(�,�"����A ���D���� ˰��w!NS���h��e&�!3T:����z6X�J�lW1��CN�9ʿ	��T	$�9rH���p�m�����ݤm�1�ý�_T�>7�dO��9��<�Ng���}�L�h��D��" NL�'z?���~�l��ٻ���@�zL?
��pa&&���]�_l���D�~���!DA#�=��C�k	h붹���ݕ�k�/^�v!�~�{�qL$�m���Y }u���}���N�kL���&` ~�@��쭼i�T�I����N�q<��D���9��M�]�/]�U�>����̞�O�<8�9Q�;}$����û�}�)2��:�xq[}sԝM}�K˽���<	�>%f̉$�w�TI�Ვ-�� ��g̔�E�%�Vo?��ڢ	6�hSj�`�����ݗ> ����n���,��&g�k�EL�q}�52f��A�{�(�ޒ�q�ނ_|���r����K)��xڈS��uGĜ��3�Vi�ׁ���� ��2H��uP0n��r5Y��Y��zF}�k�oe���+k6��g��y�JLT�.�k�!''}���M�H�{�7{NA>$�� ��Ϊ5�(�}.A���sr���PL6�m�����t8�A�sQ22���$@��$�6o������vKru�}6�����*oe�E��w}>�A����$f[�镱�\��ё3|	�}}�#7�K��h<��͐�����/8,��L��hF�w������eQ�el��DD��Rvo�k��/�M��I��.�k�P�*D�'����s��O�kڷ���p�t�s��6�����ϝ�W��3��P��2�n���"{�d	=�T	$�u98�T��C9g_ ��<���9!� \��;�1��2�5��T��7+..Aa����)��x�H��o� aw��G����ҜUЩ�(m�L�K���2�H2�������~z �6?���w�	 �}�4	$�����q�y��f��ڞ$
T
�>P�n6�滪�$����D�������Hw��0 ?���X�%McL������9��"��iz�o0�I$��"I�!f���a�����]モ������E^J����������Et�#&,݂Ev,!9'3 rJ�Ikxv�8���t�u>�'�������J$��� ����h�{0C���Fm�P$���⳺F^�M
a�7\���ㇲi�mq��#�eQa��E���l�l�u�S�Il� 6{����,��9ѝ�B�'\�,ޙ+E�l�`�veW��_O17G��-C�`6Y�AoM�j�����1�f�$���Y�Āl���Vtt�30�TT��	���>$g9$�ʳ��h�q��ĂK�� �Vo9'�O��6b�s�&:���W���SH$+Ι�۝=�N��d�A�x�ܜ��6ӈ,���7u�$�@/�zkǓ̌��3(�m�O�VoL�A!��PJ�DM�b���xLͽ�ݽ:�;"�=R �I������~�1���Oe��ta��9?:�b�־��}'q�����Mt�����M$I��7�~#
X�f4�Q�q�Ҫ�b��a9�5t�Mɮ���0A����4��uN���rJt��ue�z"�.�5�x��기,�8w>���՜!�^��u���m��r��r� ��у�]�us�lp������w%�kY�����.�s�݇v5�3�I��<;�L��:纶qv�t^�v5�;T���O5ȼ$�Ԑ�q.k���%vΝVۥ6��F������B�֝�N
ï�?�����mL��m�$��vD�^�t�3��]�9�y�"������_l�5�	�m�X��Ę���  y��F���E����B��$�s��E<���>^nm�$��:��C-�6H�1�S ���H$�Q�֌�E��R4�Wf̂{��D�hJh��!�wϜU�';]r���vD�H$=�ڢI�s��Ux��n���\��o/M-��~�0 05�{�[���Eښ�	ں�'ć{�T|��KK��=���o/v`)��m ��:v�l��K��8y�u�ٵ�B�,i�qջ"�;����O6ӈ,��w��l����'���}�U�;���Ĺ";:d���j�#(i&�g`�}~�qo�����Xw�=�v�8�jb�/�YSE�޹b�s���r�\��m(��ݹ�n�;�kb̈́��Sn&�B���T������A��rA�86ugUs�a�5�V��F���)�d��.��� �g1 ���Q�uTNi>/3zh�A��r��(6[��l�P��ꌿ@��Ѡ��[SD���bA$�ޙr�/�Йܶ��ɿOI�Kp��V$�x�	Ƀ�y��|Ug;���]3V�*������$�f��5d[�s�C��0r3&�@��V���bS�U��nn���\=�-۫r�ܝ�V�c��Gߋl0���.��@ �����>$,��B,b��l��5B�>1�\d�ke�e�Λ�����ͦyRA�WH�LFl�$��D��s���ag�Y���;�{Ai�[8� ��f�H+�dI$}��/�λ 䋳��GZ���xc��,���v�"�}U���fnl~ه;z7��n`PɌ�A����4w;m���Wە9�<�弞 ��� ��$ݙ5�����UQ=�L��osP�x��?O�
�$I"7���w����l�	�b}�mJ!�%��
A]�2|DvgMi;��Jn���t�D�I!v��1��Tr1'S_ӏ������\n�+/N�s�O�^$�/^3�e0����ϟ/��2s��5��������f���rI/dI'Ĉ���6EZf*���s�Awk����S��!�ā]W�^"�lu,���\��
��H$���)��઎�D������Zb���L�LgwM I>3bR.�ک��c	%u��'Ĉ��[��
p�I�I�V�>�Y���� e�M���vl�$���)ښ�&�T�7#2.x὜�Gۄ���NНɱ��y�;<=�x��1G��	~q��f�I5 �g�M���U9��b�!ޚ[ơ�	�dp����N%�N��`	_����s��_y}�d_M�"�:�b;��m��\/NPߛ965�G��>6�ֺ@r{xm�kS����Ë�%6�i܄#��-(e��Y����D��� ���)v�6�ffI �Ee��'�èR�M� ��Ͼz tdӑ�K:n����#w6������]��˝�.j."��
S�M*�O�6�M�����I� 0%�z ϳ�ֽf^��v��<��Dnf�x�A��rO�a����h�y3��=b�N���� �V��$Dn�>$�΍��f1dD�A#zw��7��M���Pm;$����4�n�..���
Dw0%ot��Y�[��;u�r�%�s����on@��-{�}���z���{y��9ޑ?Lж�%�"r~���U����}��h.������)$Z7�1�
+�Y�Y�0�,�����	:��r9����*b73�L�\��in�ϗ"B>s�B��7W8ͻK��s�^6yّ������=U�ݓ�l�6ۮ,�7u�z�K�ٶ�y:��{qA���@���xJ���j�s��봻�*��lf�v�ú�����c�m�û\��W����yۺ-�rw����V�'>�F��;8/p�9ͺE��L�1��c٣`�Ƕ��t�������t�bz����@b3\�A]�2%��3۲o�'ޟ��^�$�P��a̂���If�U;��#I�>�$.ޙ	w�p��\��vm�ZQ�� ߅��A+�\�A�q>��;,�ۀ�I^u��a��n�,��{�M��2�{�W��ΙK�,��q%�K�	ٳ �H���ۤ���SAQ��� Ց5���ne�&��˙�wt����QNsRز
�ɐI";�j���ɠ���`7�?�Hbh$^?Ų�8=HЈ�󜓎����n���8vz�翟��pUM�n����r	!Vs��;�j��Vw:w(��u�>+7�A"�J�.e8�Z�=�U��S+Hђ*�lU��k2�B�1l=v�َ�^y��޻��]�>�N�v��=5�NC�d��rY������;������ն�lH��������/�v�VɵBr�3n�T��#d�P�!�f
jJ}�H��٠I��X�Eu�(�Y�I&;�j��v0r!&�L:o�ͧQܲc8LV[�|H��ڢA�9�����#X�7āUuD��-��m �M=��N� >n����}���׳^ �{�@��� ߭�{�|����g�s4cF��.:�e�����52zΨ!���ca�n^�������8�]Lg콯Q!���$���0#m�Ȋ�״-��;�r��	�uW���ҋm��$��>]�s �C��ꀪ:gA%�ޚ$����*�]�I5U���#��F�2�J-Uz&嬨>'�!�	�s�mi�\�dELdX��F-'|�ޙN�=��sܴ\;x�8\���.�!�I�r��^.{)d���<�=f���}�<���C_��ڽ���
���&T�7�WE�Ԅ�����b$#�W���Sx��.��l�|2���4g�/O��w�{w�1��y����{-��P����nZNS�9%���#l��3� ���Aࡶ��զ����2^��$,�N��a���xwN�s�.��؆ܒ� i��� ���� 2f���3�WH��W�~��+�w�b��%����%�gxW�x�k�ݗIs|ߺe�v��~�*{���Cï��B��i�s;��ȑ��O+G>���'�_<��Y���lO������<sX��Z����Q�pF������|�{C�_��!��3\�4�Y��gf�!���/K 7R;�����3��~�y7���'�^'�4rΨt�z�n�9�>�A��hoM�ۛ�g�����wdg�e�{ޒ怜��>[�^?��^��t�J�e8g��	:����F~SR�4�k�=�0e�}���\5K�yk�K�����o�G���Q�3���2�^z�b�Es�ù�8�f�N�դ��v�����r���֫�����O�ս�9���=7���;�:=�-��������ŀ���q��{��ӊ>��}���b�����eW-��Uny���Y�R�?kl�����i,pc;��{�(����gf��xx！W��h���g��춟��
vty��c�'�m�G�7�g������Ǟ��5p��H�z,go���  0~m̸��
�Q]8�e*fS)nf"���,D�dƈ�iKh�kD���2Te�p���rə�an0PZ⊘�,QL�EEm�rхe�mjj�na���U(R��BѬ��2��r��9j�-�-��5�LkFҔF���
��TS)Ym�c�E�QE��1�ԋY�S�5UD�sY%CZU�6�h(,�+l��ʃ�m*�UFDV��JՅ�UDU�
�V
\(dV,\�8��-kWM-�]8��+��b%���j�qɖZ�h���[A*V�j�4�1�7-c�-`cdոZ"*�`�:��˘9K"�Eĥ`\mj5-Lr2�,XQRT�TƊ:��T��0*V���fd��w��gxݰx�pa���흋*��ˤ����]d)�����%Q+�jZ��E�T�V�FM7V�[Me�-���W��<��{;�O�N�"�+�,��Z[+[KkB$�� � ����H$<y�D�z9�Mj(��I2�g���_\L�u��C<D�ʚ��<~�H[��.��\�6'�zh�pU �p�Ú�yω��z����~���pN��D_WUx�H;��%n���L��nr�;���}{�ۀ�a�8v��'�	ڍQU�y��cv��[9�쥇����S廒f�;+��H;�>[��^3Vp�T��`>N���7��p����/&w]��&�p¥&�6/�	$��D�ol�LQx��!/(�MmFyCj2!�TH;nI�$[�@W�΢�B�4��H�r �-���U�0�L�Qj��5}Q59'�s���ē�@Y��D>��crv,C�򂪼߆nP�Շ݆�=�q���p�����i�=��l�;���>^Y�_�Y�tS;���q�N��q[f�bMzA�@�&��b���t{QGq60��"ւ��Ex�;4dn���%wRvvP6O�.�I$��ڠ1o&I�yJ(����;�����e�c��ή�蘭�oo=���=D��犑��A�-a,,/��A�<H��<�H+�:��|LvN��g�
Y�|����0e�-�d��M9��m� ~��%�d[�vIvoUx�ӳ@�s�,���j~�;^zxf��p����,U�Ϊ$�͞�Q����t2\���G(�>O�]����ڢ}�P��Cl��
� �e��X�=F'��P ���@�A�c}wQ5�u�ti9�TtN�kp�a�
-J����>$�W97s�8{���'ʫ.��H���H��\���KD�N?R����խ���Y�|��~����#U���<�z�~��:7��z�p�G
�ۘ���F��7����v��R�lg:W�@B�f2�s�vI����{S�,�v��zv�����q�q�����w��5�;,u�sof�����wZ���ZSu�qƅ��cv���t�\�y��q9xے��3z{��=Yt��������T�������!��n�Z�=��ծ9�%��2�9����x�8^t��}�;����rC�'V�l����<<���nM�c�z��b�[vќ	c't؋�l�h��N�ۨ�nls�10)�V��.8f���ck�+�0�&�?w��'�kp��G��}sD���CĂEt�$��E�ՙ��v���	�";�j���A��R�M[_C���;�l�]*f��ݒH��گ	 �W9�p��v��oe��o�v�0�h��-=���Q�V9$�7�(�F'���� ��=B���r	�2w"�p�q	����S�u���n>�~$E�t� �J����z��<@zm���^�4�cx�I��	^��uZ]P��a��O��r���Z�	w��wzv�p���)�ZW��:�D,�d�76^ɣl������C����Il�"<:�9�?4[@��tUoU	��z���O�>]��G;+�ㆲ�� ::�cj(�$���Z�_��	᫓���]tN��r�@�<t9���3ߒ��l���V��r��e
�ˈ,Zֲ������J���&&�q�{#	�)� ���U�L�q�s��i���v��pD1:�b�\�]{�@�6�Q���D��un� �f�9� �O���@��+e�pb!��ϯz���-)�+��n�r�� �J�ͪ ��N��˙�����ٙ	w�6X�J8ZGH��;�� 0;��9WB�-��`�빹	�WwUx�H��ڠv'�S���9����i�2U�K���gYq*���[�,�Y}s��I������*��s�ؒ��
 �L�N�@��&\�b�s.H>%gn�}���j�e�Q.�M_UA��}`ggf⚶;�-��H&{��`s���J,W�`�����N$����O��N�B��ыR��E��&��f������9��	�JU��f�Xe[a1�9��g���H�s���<vgé�;�Bv�]�����qdA��V;��{j� �"���8"��W��d�����'`��!RT+}��l��2PP(��}�;��	Rƻ�{��V����Y?v�����4	�{9�<�
����/�t��ִ�<���I��~�g82VVJ�]�{<J�w��?s^�{����D���}�y0�
°�,O;�l�NVJ��c+�w�>���w���G��0�2CM��l��rrr�'d����+��k!6�v����gi��n.c�����fw��0+RZ�}�vy�B�B�`Wz�� H�@�ߵ|�!x��O����<gᒤ*~���Ăß��u��k��0�y�oa�
��R;�y�zw��>�g=�ݟFq����{����A`q���{��Ry���<gx*n��̓��6w�sQ�i�����L����ed�����x�P���D������}������|�۞}0�
�RX�w���$�����2��;�����_33�n�6��xi�+������G���~��+珫�R
����<�H[HV�+C_���@S�
���}�~�8}_؍�B3b(�G��V��7"����_F���}����t�ʕ�o~���������G����p��ӭg�>�&mM�nڹ�ʜ�b�����������D9�9ݜH,9��o1�f:���u�8�]y�w���IP�,B��w�8�{U���;�D��@W}�B����`X�]���- �B��;�~�,����z>�OT|���M�x�I�h���`숚�67d�q���g��v��5��
����>m2���H�쯷dYed����{��<IXg~�ۇ�80�>�ߟ|��i3�{�Ğ�+%Y++����'�P=�����Lֆ��tl��V����q�AHy��ٙ����z'�3�EpC�$<@ �9�<���J VQ3��ۇ�d��%A�]��zp����g�tIX|W���f��sKw0�0�;���x¤�B���߷82�Q*.n�����������D�
5�`�_�����)B�>�~�8�^O��/�C�ϒ׀�,�Gכ"��xxl^Tי�;����L�������*IP�%aL��~�a��aRT����8�;�7�~�L�Y,ew����"F߇3.b�*jSU	&�3�;�p�Ƥ~�y���矻�闄8�`V�����<@�P+*g?w�É�d�T5����!ĕ�ǽ��}M�ͨY��� �p�W�b'.c�[HĒ!wv�c�s3X5W�P*���U��uy׻V�K��@�ko��t��L.��:F>���s�X�I�p`�ti{se��Tn��ҙ��-����m[��w �Գ���	�n�;휯��m��\F�Q���4^�$k�ݸ�����n<`�ݑ��bѺ�g**�2Y5�����7�ێ���Mm×m\78�q�^����ۗ;��p���{{m�/���p4�i����e��=;o%�'au�Ի ˮ�|9��l:5ܷK]q��n#�����=��c��a��H۶!�����ahi���������,�h�.c��q��a]���a�
�RQ
�=����8�P(�����ÈG�}����=�P~���8{:�|$���=��nH/��w��:��.kk<���$��8�@�����9��^������>{�=�βT*J�XS9���q ��
�����6q'����ѵ5{��O|f~�y3>��^��
kZ-u�����?s�{��x��H[@�{�l󒐩�
�����6��{�~���(�Xg?w��Ă�FJ����6x�V�WY�kX�4�>�P>�ד T�M�8�!���IA
��>�ݜg+*�P.��y��%`Q��|��Y��np�w��oH)�{翹�q���x���52�Lqu� ]���<OD
�*As�;��A�����߻���I�	+
k�~��q�#
*��l�'
�YY++��ܞ%@���~���?o�s?������׫l�y�<���j�͠�� �՞�xx��Ch�.�����T��r?�I���y��0,jB������<H<��l`V��;�� Tϳ�����M��?2���y�É�d�T5��"�G��W��H�L8h����υ�f�� H�#�m�`��\S��#yq�C�Q9��ç�����Pf,�Z>�	_�����0�r�������(!6V3 aR"6bbj�N�̹�|�d�g+*A@��o���A`q����{��i ��3����f�n6�D�1�N(L��$�#��gI��e+)+���T*Jýz�?y�����}�
AI��~�gq
�FVK\�{���%@���Ym�����dd#��� }��m��k* ^��_���$�m��BФ+Fu�}��)��R�S�D}��>}y�d��tnc�D��H�$	 ?�rE�,�#�A�\6����Ƙx¼󿷰�0�,B��
�;�zE�Y��w_T�����K} ����}��+�`Q���w�ZA�x$�#����̀|=B��d�D��{����8��)��n�\o7l���Yi�EN��;�s\poc�M��߿���~������������~��$pd�޽�{���*$�.}���8Ì+�W���w���m�k�vx�Y8��ew����P<��D�H�ę@��fd�0�ؿ�����g�"����S���� � }[�H�< �V�+�w�� �y>�~�8�2VX�P�w|٣�����o�6~Cؒ��=^�_K�Y������a���w{T�!RT+���g�J�x ������lH��菃!�9n횰�2���_x��s=�T��?jwO����C}���y,�r���K9R1|Tv�GA�|�W��ۏk��@��
`Q�������l�-��߾��`�N�Sm�ш�ˈ�$P#��۲,��������| G�}�|�}+���{<d�
���>�{�8Ñ�H)*k��8��G~�{����~d�ed�+���ܞ%@�>}y�5u�-5m���%a����
A@��yݞp�.~7ˣ9Ϯ���!��+�|��H)�e;��ng*AB�5��݋#��>�0��;S�)�9����(WfU�kq��uaq��[�ې�����z��}�����5�k��H/����:0�* �����83��e@�P.��;��D���=jo�`~k�����H6���?w߷<�q�۝�ѫu�:�.��ݞ'�e��������~���@�����}�@@�"#��(���0�

�������N!Y(>Gގ�ڇ�*�Gy|}[}�7��>��J�g<����2�FkW�@�+�Ͽl8<H)
Z��>��!HZR�jz�>ov;�7�=�	�O��߾�<gJ�*��;��8��������N�\�א�0��~����qv��s�H� @Dyx���gղ,[%�*J�M{��xq�X�⌿���ޗ�����n�!�D��V>������5��vw��A�����Wlf搠����0~�%��/z������+�w,ZF(U�m�>�]��y�AH>Xo����q������b#M%!�Q^H���G�>��&X�]�����d�o��_���~&!�+�{���
°���}�Ĝ+%Y,ew��{�Ĩ�=�����}��߽�v^=w;k�&�<n͎�����;��i/۴n-M5s��0׿����F�E�[tt��Vw��l8�A�
Z����󒐩��[�}�<���>����矯?Y�>矻�q�++%@��y��|g�~.��kX�4��i��
��wr��� "<��������K����s�}��q���*�}�� q+ư+]���p<��m!}����ʣ����ߡ�>>���9Clt9�'�<����q��J�+�w���d�Q%B��9��y�M�����߻�;V0�(&~����N!Y++%]���ry�s�;���ֲ��WYs6bAau�;���ֿ���c�gy�?~��g�`pjB�o|��Ă�^�׾�p�*T
ʚ�}����U���V�==_.���x�Ȁ���'?/>_GE֝\���!Ă��op��RQ
�]��l�g6{��}�_ƿM T�����A`q�޿w{����;�{�x�d�s��|C2�pY���̏��!^<���B��Nr��	�|h���Z.ޞ��n���ⱺm����Tm�u)��Is{�<���A}��l�{��H��I��h`ޜt,D��~ۉ�r�w�����5v~�v-��rG���'���������==�6Z���9�T��S=�®�y��&r�]&w{!:N�\|@�i�q���l�����p���M���z��Ab,�L�ߒ��H�I�.>�/pjb�t{_�^>�.������V=������w)Qx>�/'��[�ב�[�(ٺi�6�Lض\So=wK�����m&Y�O�w��ٸj�1����R74�C��W�ί3x}�6��	�Ox��-��]���*��x�{�S<��l� ��<n��Ӧ���,�)�=d��t���&����k�����c�s���O)mB�� -�8�H\�;8���ڎw�p�s�����,lN�o��	[o~^��<�H¼����6��F{y��}�wp�{�[|Q��1M��@�U��SH���i晛wz"�z��{*4��m�ᕬ��$�Kؽ�y�U��x�{�9忏]%v&:l���F.�]|$�>��OV�uv��R
�~����Q�{�^����n��bY��k�	�ޡ�st�ԍ����xʸ�W��foM�h�uIŔt��ȥ�[[��N�ɺ��ٽD�4rH�T��oϏA���2����,o��������PZ�g���A]1����1��w��%�eb���8}��]�����?x��<��$��Z4�KF�,�Jֈ*6±�DkE��ֵi[[J�հ��m-���N �B�4�"�+Zbb�FҴ�Z%XV�#l�TD�6�nTkE�R��m������j\�2�*V՗2�\�(e1�YufV �me4�0m�QbU�lYmE�W)TT��*�F��U�K�fUW-Q�f8�lV��X�rܵ(��
�-��mDM5\��Z��,�3%J�ТRآ�����ɆQ�ڥ��R�kb�&��q�w;��I�;* �i[J1��1E*6�0B��![,�V-)\�ƒ����Q-*�B��Y�0��*)X�����KQ�q���141�J�%`����m����ņ^v7m����9�Î1�v�Pq�q����jmkh��Q�WLu�clWT��-Z5�m���Ҫ�k�¬Z[DeJ�kY���6Ֆ��-��%j�Z��Dij¡m���.`���ew���G��=.��E��q@q�ٸ�;��ǆ����\��v���l��c�scA���ķ7�p���Euy�%�Xٱ�]�:-�쓇��Ӝ�uO/��nc&]qЪެs��l�㧚�p�F��qF
�yvÉ�3���^i�=�1����v4밭˼�m���Cŵ�����`=��cq���ۇ�	������V��]{n�\n���Apn��&ݳ�JK�l�����s�p�]�2���Ѩ����s�F������]����I�y�o=�=����0������ᶍ	�l�Z�B���������g۞Ɋɵ�bxڋ�Z6\�j9G�E�[�|.���С����j�t�۝`��sێd��j�G\V��#$ȧ)�U��/$�2Þ�;����k�����w���h2
t��:����h8
*Nݮj<���hNjܽ�x���P���(�Q��@�����c�+�۶vyN=9;;��[3זd{Q��1\�i	aN n'��糮9��́���2]��g3�95�ն�,p�$l>�� ��3�9p�9y�Tm��[����v���78�SΫ��Yx��b��S�9�v��Qmۄ��'�+oq9ڍf�]��r�W���\o&�8��0�F��1��kf�{w�m�u�k�Ltq���M�5N.��qc�N#v6�0x��s�;�.;�3����*W
p;����\�N�ky��S�6W��k�R����n���\n��q�݅����[���ݶ�%��q���ƴ�A�=]�x\[qbg<˅��d��/'6��8��]����b���9�i�v�I��v���^9�m��b�����ۛ�%�n\��G��q��.�g���^'#�V�nm����Վ.\�;�+��#y�=�v��[<u���n�[�:漈[e�l���N8�K���j�s�H��^5�t1�Nm���qm����F2�H�n#��[p{v��`u��۝׋��x�8j�)��{�����Z�n 8�Fj��uOln�:�8����;yؓOFǻRl�B�7�;'��|�$:�u�X��n;UFp��=\sO���ٲ�v��1���롎�NC�ݚ�\ݕ��pj[O�����B����Ŷ�\��[g��l�����p��w��X-��8ݻA���E��mg�K�Z��=n��6�;�s=j�<�n{�&�8kd:^��-�:��s���v��ں�Z3�����m��ճ�A������E�k.��fk5s�@���{�}���@�����޽�{<*%B��5�}���+~o���<{�����'�~�vq'���������*���y�iu�.9m���%a�������R����������6y�BҐ�����<���J VQ3���Ì�2VQ���y�~�~ú�5����ĕ���狭kZэ�-�a�¼󿷰�0�* ������� �y_w{n�������O��V�X��߷�ZA������Ï��>��˝�Ѭ��4S<����<�}�����3���~g*A~��7��J�IP�J�߻�8À°� g{�l�#�<������y�zɡ�����s{��*�y����j��c�\��������px�Dx/$ ���V�Nf����X�<��o�~�@R
Aay��n3ᒤ(!��y��������������?u;��1�] �9�,n�v�G#��8��iѝ-�x,�?6����hբU�����»���a�
��R���g �2VT
%@���y��	X3��}C�s�1��Q��3�	�K�>߾�6|(-�J#&��ᨯ)�$�{�ݜNA������x�����JǏU�����]�{�ퟗ�
gEW���uZ� �byA�Ǚ��9�[9o:�j�vko�nk�0�!��5�7�g���!?��������%B��YVg���|�q�H(���g�8!Y(���~���s��O��;��O�1������֛�[tl� ���w݇��Ƥ-�g�w�<�H[HV�
��w�&gu����_;���
�@�be9���8�FJ��P�g{�l�IX�G*�[m�C%W�>|���{����&TNx=�����Ϸ�Y�,e@�P,3�{� q+�`�3��|
ո��yш\������K����~>����a�l�J>��;���
��YA����wg��A ����5��x<H�>_�w^a��aRX���sgr!Y,Y(��}�w�_y��i���\��R��qp�u�wi��w]hx����R3w%�I���y:�uƓ_�����2I1ҟ�w{�����p�ѩ-=��l�!l�+X"��_��D'	"���I���π��ɯ|��Ì�d��d�PC?}�6qD��?/:���Z]k.f�r0��滰�a�(�I����/+���OB���{�g��d��%@�����8��Z��]���xe �=�����vV_�_x}su>l �[��FD&��3Z�� m<s�{���@����2Wz���&!D�
��d���o��|�ʟ��t�Y�0�����Ͱ�X��lnx?_y#�ӼG���1��s�o/ݤ��������ou)�u�V��k� #�y��a�+
¤��}�vq'*Ad�����I�x�}�+��a���  �|3����y�9��<��Ձ�R
���l󒐩��������
� VX����Ìd���i��$�����<��^.fen-���sA�F�߾�Ov�M������g䂁ɯ?{�ÈJ���
�Z�u�) ����p��y��ך�9����k��c��kZ�r��Q��t���m�n:_I@<�j�r������~��kI��v��I�}��8�@��d�����!D� ��;���8�X8_ψ=�:�Ox2=�#rn�Y��ed�+�w�I�� s��wNk.��5Mf]�����o���x��ԇ߽�)����3^y��ԅH-`V��}��
����w�ngJ�2T<�O��p�٠�28�|+�G,6N���zº�ϴA��(�IP�3��ݜg
A@ߚ���_�;��������Ο p�+R�{��m �R�w��p�������g3.��ֲ��	"���l�"����c��<k�Q���Wz���m�
$�.{�{�8Ì*AIbk��vq&��w��w2�Ur
u�w_�E�@7�X�3��5�糟�/
��x��PD ��`L3Ud����:���L}�w <=��d�2�Q����w'�i��SϽZ\Ӫem���%a�������i$ ���EZ>�'o�u�8|hs���@Ă��~���<H,��P���ݜC�+f}��s7ߴc���j�2lN�jܬ3��\�Ƌ�qL�f/7���4�X����������c���}�;�a�$�
�=��9R
7���@�Vw�t����s���3�?w�k���w�R)K����f����ȏ�4�6C%�DY<���8�++%f�����Y���i�����IP�J��w�q�V�ISz�{��8T��u��M�ze'~�9'���z�T�p�qCZ̾��V������R�7���$JB�`U�u�=���;����1;*T
�	���w3����T*�{ݜC�JÇ�=���4hֲ����0��g;��7�}�����u
��V�?{���%��J�M���È�Rƺ�w���s�����O����!ia�o����}�;�_4���<���'<��vq8 VPd����t��dΜ�ϫG��G�zfw�C�8°�*���l�'
�FVK]k;����@Ϸ��/������6�v��K��ݧWa ����}�cN\���>�x�F�ՋQ���ڈn�G�<m���t'Y�7*���j�?�K��{���������;[m�f7>i�t��\n�T�ۮwǅ�P��p.�-��On/6�A�O���Œ�/UL�NͳR�ݑ�7	�U��%��J>{n��q��2=���tzU �%��ή�y2��m��gF�@���֊��<F�U�R��v�$��7g���5�lq�u�8z�F�������-��S]΄�;�g����i�^��4�-��j[s�r]�Nq���-�T�N���i#%<n�=�k?7~��p�w����>�ﻰ�<`Q�
Z�����
B�R �kZ�|��7��m�Ϸ��τ���p�AgJ�Co~�@�G��\#VPi�Ä�����0�<���x4��T���{|�����k�Cl5�{ݟ�%e@�P)�}�|8�Xkƻ�w���A��.d�Gl�o�}3�������D}	�5M3�ND���;��ȁYY+(�]�?wg��HQ%B�+������OK�}���aXV%z���ĜB�VVK]�;���'�7w��Ӛ�э8�B�G�>��@�����B5�Ӭ��������9HT�с[�k����+*g~�w3����������~d�Qo�vq ��x��F��2漇��϶��AH,����Gޞ��9N����!�YG9�k��n��A��-,3��É������w���.����;s����{#�\lmƣ+���k�^��pݻ\#� ����
%�$�����g82T��y�ہ�x��D��w��p������sN��x���{�~�Ă��ed�+��nO"i������uq��<@�J��?w�<H�����W�|D��yk�Y����in����;$w�ރ#T
{�D�S��wc��w�:�T���l�틚^!יs��3��$o������H[)
�l�����1<�( VX����w�g�������rw�+�����Y�<������m(d��dx�{�4��RT+�~�g�JʁR�}���������D�
��y�w�j�m!ia����8�[#�p�L��W�� Y\�"����߻�������s��<4�IP�+3����q �� o_}ݞ$����n��h}���������>��eJ���a�0�j 
#�u�`��G�H/��hx%D9+�����*����2|(wd�xE!x VX�����8�2T���o_}ݜA`�#�V��[c��ZPS.n������lG��vƤ68�H���j�m��4��ޓk�;�}�th֝f\�aĂ�k���:�ID+������$
����� ! ��!G��"������nH?�e�s���ǌ
�}�;�_.�����s�O��������Yc%f��>����Od��;�l�ɈT� ������0�+
��o_}ݜI�+%Y?y���3]���ُ�s[ܟ���zzasN�-�� pJ��?w�jB������)
�S���g/�v�J�3c��g���5���������!uo(�k����:�J8a������W�p���������^2Э��$p��������y�O�R�V����<H,�%B�K��H���|��A�&�i@aW�#������g v����K�x2=> $�
��~�7
�{��xq '�_�> Q���|����k����B��wϷ<��{gmu�ֵt�3�NL��;���d���޿?�W������֠.=Dy7���!ĂÌ*J���������-���z�� �>����zQ���c[Y�h�K�� g�[ڍY��Nv��)�#h�Jm��Y�08�P�p� ��|#{2C��jB�@����<�!RFu�뻁R
v�vs��o���m3�����r2VQ��P��{ݜC�J��߽o�WF�i�e�y0�º��wa�ID*O/=�?w�>��>����ќd�*�P.��xq�V�`Q����|z�)C��~���:Ǿmώ>�+K������sYnyi���}�vq9*Ae+�w_l����O"#��7�][��:�j�����>�X¤�o~�ݜI�
�c*As]�w�xzo����sN�-�� q+ם�k������5��H�� �eȫ)
�Z0+L���*AO
�>��|(����8�R0����8˸�)F��ѥ��W�FC�����@�f�)����'.����ɣ���f�*"��*"��Kr����=�����ިT?�s��8�V�3���˚����|��x»���l<a�(!R����}�T�;���x�@k�DD�
5�Z��w̤��;���Q� �����A�_eL+��L@�68�<vl�����Xh�p�������\�ɻc���ļ����5�l��B;�Q��ϤY������~�ہR
Aa~���
>|�n>�ts�#�E=ߤY��d�+%��k��ܞ& Y����5��ѭ\�|1�+�~�q�� J��}�s}Sd_ ���	<���~�|�R
Ag�3����q����o<��uy������$�7�[�ѣZu�s^C�8+�|�v1 ��V�ﻸx�P8�>�ߟ�߾�_�������8��+ư+\���p<�A�!Xg~����~��9Z-A�P�1>H�믾�B۸������ށ�x2VVJ�����LB���3߻���F��*J&�߻��?|�������[�~�N����]�
��M�z~4]hu��U���?s�{���Z������vx�o�o�_w�f�_�?8��?w]�
� T�������gJ�*�wg�JÃ�.����������&"3-\Ș0#�D�ɡ��K����냝�H���o{�K=�s����<inB�?M"K��#S�3T^~�� gu0�'Y��Z$�J���^Յ6���烒�������棦�1�]���1Mt��yJj�g�k��Fj8m�
썷K���������w>��c�omحc98���W�n3u�[�X��SG8��N�뚛y���'F�\����t�1o ;��9J�ܝqeyb�ˮ��$�j�F�.j��laLǛh˝��rsr�u$F��i3��J=\�]n���L���'u��.�tF�6z;�>!Ap���<���Fw�H0Ă��+������%��	���@B>h:�;�Tg�i>�O�e �B�a����Ï���_��\u�7E)�@�q&{����AgJ�9��w{���}�_l�2bIP�%as����q�T������vq ����}�GǾ��}9�-����'�ջ]f�4kW.]��ؕ�}�߶�
5!m}�l󔅴�k�qw������r�� �� D @��t�[82T���|��8�"J7�o�� 6�DC�>�96��;C�ޅ]tյ����G����|6��E�}�JʁD��Ͼ���+X(���> �h���*[��	�5�\Ï_�/�_(�.e˪��m<I�y�vq8 VVJ�J滯�xɈs����?k�-��IĂ���>��!�aXQ�@���<Iȅd����+��><�g�ggh�Ș�~�M@��7j�8�g���<s��=ll޳��n^��������:�۪���J��{�vx��H(��wg��-�+X�o��*P Eg�G5���}�	>����>��Yc%B�k��8�Xs�7�y�Y�ܺ�)|��x»�u�a��Q
��b���7�4���W;=��[]����s����1�/9c��o��~��܋N%X����Ѵf��B�)Mh�jk��������t�Q�@�߿eQ�?���H������v����[w�	+G �6�AA��8	��"C��(�����4�s@�Ao���Fll��i<l�����JC��n�Oz�3g>$�8ψ>oz�,ٺ��4A��l��Kō��Og�\^� ��2j�ç��n�ﭲ�f��^[{�@ƌL�34�� a��H��v.^ӱ���.����ruݕ.=�R�mAv�g[_�{��\�p�&�>���UA ����>%u�U X���o��� a�����x�(�E"����{��;#:��ed� �D<|gĒ��P'�4M�~+�v3��r�<��R)�+�&�\��J��M�f��W��6�mn���d�Sk�~�[s�<�z ��e�~�c���s�G,����ݼ^՛��C����M^�ۥ�r�����wpa�<5 &��,^��!'S���K3ǧ��s�I�r�� �Sӻ�Xca��zn����Ǧ�#"m��-�a���uqH�>����ye�����7F��Јy/<�wW������˖�y��5�U|2�N�|�� �[�Bv��<�y;��s7C�+_\E�{���vlp�*��1�\�����h;��0i�����E�m�V謝��`������<t����c�<�+��l��"܀��;ݰv�u�ϱ�3��ݧ�ǯ��@�^�i��Nk�ϸ-Wzo��y�gwnv��{����Y����ZJǇ����{�w^��Kz�9�ʙ]�w_��������=���fxO����QP�l9�zPE�H�q������l�/��V�3��[���N����Y�/�F��ׅ�糦�ș�S���	a'a�V5{�����&L��VT��Wta:�£=ǋ��e�z��e�����J8�����ӡh�{wx�83��}�����S	�'O��x�}�/8KX��'�'7Y4o�Ǥ?q��#y��yE�0,�Vm�0y�9M������ �wU �_+��y/3���`~�hw���O.����>��8b>�7E���Խ�������ӻ�ɪ���"�vh:|^�ى��PE��B�+�.\�&+�)klJfa��q���JR:���X�b���.����M@����.(:�9VhʰfXQ�ض��22�R�,,n�Ĉ��`¶�.�`SY�����q*1�
*�Jʕ���k����VZfYm����eeU��f$KV�F	��2�JXղ�[k�-j"�ZXѪ�QU��%EW��DXV�F�e�sb�2[s-hb�Z��Z�9�TU
�@���-��J�D��(֒�#keF��+R��N8�+l��Ym���U)]Y`���Zб�QjҨ��Ve�"�PUĕm*��qb�J2jbH���(��*�Ԣ(�T��Ub���1m�J5*QKe��[`�ƍ�*#*�Ī�Ҋ�J�mmD(���DKV���+AU[�G#\r僅V�er6�X�����[ll���L������Z��D��b��AH.�l�UA�����$�xnu�{�a�(����,TrCi�)1���v�Ñ�b��?,�@J�Ϊ$=�Hs>��1�J̋�C����O	��?O�@ �߻g��A���u��>��FI%_oUI�=�9�'�T�՞���2F/��a%wq��㛀��hޯ7::�)۳���"�x,�~v�.`�ڈ�zLi�	f�P�	<��k�**�ͱ��d A>U۵D��Ib��	(����Em���m��� ��ίtoT�/�ᘽ�[j�L8�F���4\AI�Tf�:�O����$���uQ+VN�_["��TI1����p*�6)�+#�F߼}����1��G���u@�F��	�r.&K�9�|�O ��m�}W���U���z��ճ���P�n̽���DVxNP�>����^�
��=�9%ӽ��b~��< ���uuD��G �2�P�P���a�t�������� S�##+�Q>������a�l��*V��2G��}���Yo�x�67]l��'H�Ig��6�=��8�:�M�����t3�q]t(��6�$C��+N����W#�#^u�b7��0CmDD9�eGHD���H�W-���h�I��uD���d |gT�U�z�"�����	ƁE�����&��^�"H<,���crstOFu�	0�6Q��a�È%2j�����:���`�d����@��|��$|6/���+&�+9J� Ϸ�&L�$~��i$ajv.B$��y�DX��K��Xo���$����$���F:w�j�:�C��͉z��Z��F�Ir/�x���~�tr�����k��ˀ��O��1v�F��3j^؝�Hۅ�K���ϟ}���`�,����g�\�\k��,d;a�G	�'j�:�:O&�k�Ց��[�����+\�kFnŮ^��tʾÔ��F�h;,��{�c���b�A�<�#d�:팛%'h`P�Vg;BQ�	�g��k�N���Vێ����nf��-�`�'��l=�*�m/����ܣ���NN�7FD��mك5��v�c;;Nv	Z�z-/"�	�ي��4�t��l%��jÉ����������8�բB3�u�
�&�H$���
����h�n����0~	��p8�Ϙ8�/
	����� s��.�ǲ5�� �I��ĀA�TH1��:��*�>{�����#�<�)$��
Ϟ��om
 �Նx��YMv�
6�A;�T	�9DхH$�ч>�ʚ�F8$��$�|Wnt�$����ؗ~H�ݯ����e��\/��a�U�u��D��sF�W.W�-��&�$�+�ڢI�޺�Q��u��n��_�j��	�8b܉������v�V��z�RԼ���V-;����͠�a�rzؒJ�͡D	�T<p�̍5�.�2|� ���4V<B�f!����& (��P�`r(i�E﹍���p䈋>��b�h�g��!נ<�K���=��xl��1x�w����y�{>)����X'��|<���1�>$,߾�$�z�'{L�uVlD���.��4�!�GA�}3 �3�:�I'�=�)�mN�$U��P �{� �w��x��)ɁX��(xސ����v�Q$C��ج���lE����zL�P1a,Rd'�wz��H0�6|������X2�u
 ���u^$a�t�z�k�ܶ�l,6�

�Z�8���83��5��t�t��.n��F������l�\A�d��ݵDN�u�x�H&w)3}5h��'[�6H9�"�$lō�Pm
��ӱ��?z�U5:I tmuP$��tǧ\A���̑}}U�'�X��!e��]�8A�M_O��K��jO��G��f]���*�&���_� ���?.���6��>��r��϶{�&h�UyA-CV^WFgA&p����:�j����Q��x�� �����s�w�"�u{��ך}�p���1!O����.w'!�o�#3f�$���'�'ʻ��r�s3&���s~�@7z�8[�ZE9���� [��*]�x��i��=�g�6��H*��%V���1��`<�6�%0�>�[��v����\`��M��qp�jW����[���a�	tL�Q�}�W�D��n�@%Wv�x�Y��wO9��UD���60&M'
!�T�����gH�|��M�Z����x�	���B��E�9Ν{���y@��@l��D��R��*�:�@���\xL�ٝ��e��A �+������H��0�
L��}>A��ǍOP2i�f	 ��m
�+����n͙�܋u�ϧ�ws{�Y}s���~~p��+��$�I�b� W�~ѣ����0��A1�������2����'N�5�ΎS� =�<�f�����8A�MB�
���� ���hi�#i��ās�A$�of�T�t�:�� �ġ��}���Z��ci ���F<g��s��	m���Du�!��:�R� ƈw/���e�(u��j��>'�v��HS��D�`jq���oڰf o�}2ÈFE����9��ʠH:'D�/�%�y�����t�'���W��qy��zaӝ��n��v�`pM&b!�B�$iO;��shkS��Q0.�ТB�ު�Tn�F�jj(�b�M��;=�S�*}�B�TgmQ ���co�o�``��>���X��e"���  6���w�onҝ̙�;�^$��٠H1Gu��X�wku��!��8�]lTfΠ�g�:�:&��@�q��J��&���Jw	�������Zv�6����l���{�{+}6�Q�J ��,��:t��v�ݨ;���tk��S���S'�\���l�۟n�14.��S����۞m�������:c5�x���\j��;x�(oem�]���+�[�d#���8m�S�\=i�
C��3��@�\Vy��pkU�������,s�Z�!�<![��9g9#�պ9q��V���q<�jV7j^�����R�b���N⣥��L���p�yT���qQ������1��R$
?���?o� �3 ����{*�rY���u|�ܿcMD)��6L���QM��MB�TZ���q���z����~� V� ��}�p`�]�ͧ�.o�T��p�:73���Eq)�뗾� ?�^�  ��ӽ6�MT߈!��P�K}dX���0�L��MW����-���2�]�����w�(@0�0����#E����/_��zL�?vr3��$�g	Z9�\�.��꒝�c��B�MENP�a�d�Iw��X��{7gp�,Bb �OHl�7unջc��Vw������۞M��76����${HBa�����TI�4�$���]jQ=��Ê��D��A�ђ�:��X��)Q%�~�� �T�����
���.:<@)����^� K��˻�>l��?B&���q�[w��Xv-{p�ڽ�<���k~� C\�{��[���q������}>	k����?@	/6K(� ]Q�$��ڣ�Ayu9���2Z�� ���@�@[��D��F�	�
 �@u]�	GW��/���G�y�U�A!�������66F vf2Q��Q��a�Q���� �ϺhŅ]gF+��_�$���B�	} ����)~3�u��?F���A:���r�j.8�g�}�����wgv��t���y뾌��a����A(��b��^mz�$��=ToP�de��� ��T� A]{�^'k3�!�ZP�UgT�P"�f�bWV��LQ�IW���y��^$�K*ϻ�N4;�o��j����:?4�%QJ��]^�C��� �Y���K���(���ㄼwg�B�!�G���/r����o�����!f�"�+�M�.1�p'iz���{���x{�*���'��nwUI�y��Q"0��RPm&�C���"f��)�`��ͪ$�|�Q%OGX�u�x\���w�on���H�4a�0��9�گJ��'�x�����
��j�)��X1dWd�{�U���>���'�灲�/�I<�N�MŇ�+���uZ�=ll���g=}���������&��Ρ@���t�'��J�|d�U�s��35�kޙ�@'�=]TtRW�h�L3����?�o������?�W,>$�U�@�U��I$Y!��6osN��Gm�v�#��!��j!Es�r0AUq���9�P�ukF	�n�Iͷͨ���!S�.>����	K�V�%(웚'���r+��O�.���+S�vT�:�q2Td�*s �_�����o�y<�*秸>VS�^~�@o,�|��oj�k���Ί��m�� xx����ᝲRPL�QO`V/�� �o���>�%�}��޻ �ڝ��A���$��y�D�Z����zn*g�J
?�(	�N	D�x���=�[lp��;�ܩt�:�tu�����&��;* �����ĂA����DA#��;잰�u\l@3wTO�19(��,�ɖb!�U�W��(�&9�P�	f��UCv�:tO���׆|A�B�ryt��u�f\H��@��8J��?�o�$�ݯQ�>�Xb&�J�R��$bz:P ���B���� �/�A���[6HCb��u����'�#eJ��^'�z�r���i�'����wQ��ۋ�ꪩ*$	.}�5޾�q�Y���X��&[� ��Ϊ�{g�h�˲�q��	o�}�[ϟ�{�c��'a|<��ۛ��1�7��f�-{���uO�nf�NYX-�j��'B�/���s����T�w��6���ض���(���,�yA��ǶS'��G?+�{\��O؏����� z����܈Mbp�˹q`��O�Z��˝ `��2�^Sg3�=���6x<	�=sW��s�o,>�����06�f�0U�ߔ��i��@��+� *�<�����gg���� ܈�3�q�8)�.T���a,�}�,y�s�������n���4ؚzG���:�9�HG���w��{�D�_��=ь��x���;G���]�s��|��M��ܢsۭ�ͨ	��л{<�(hɞxʎwBZ�Z�Yps��"n�ҜA"2�F��c1vl����!ҹ�"�1�VZ�X�P�r3���3�ԧma��;��'����y�^�������{G=�vmS^\���=�жHoj���4ܵ���'C��^��{ɺ�{F����}��;
���V�`���Ck�������С���wn\�{�$v �b��u����w���N#�;_6����9Ӟ�fvt/�4XNky0|Pٮg�ߞ��l��.��������x=>�
��jI\P�������,���Z��!V����<�5���3=}�W�����8�о�jqh�׽��'c���Q��<�a5y@r�/��j�&6������6��ѧ�^���Q�j��u[�u��q����wwd, �z����[�w��Tu���;y�t�씠0�7����S&�x�d�A��EQ�PUR(�%�0����G-L��\l�ejA�H� �0E
6c�1B�e��B�.k2
i*CX�EV&Z�m�e��VED��-�W��eJ�����N(��MIZ�cj�AK���F,Xa�LC0�ڹlbVܸ�,PX��X�Eh�A�U���je�YV�Z�ʠ�Qee��U1��ik�a�t�R���e���m�PQb	*UEV��+��k*V�Q�ҴR�[eKK�m�`���[ekV.e[*Vm�*Ҩ6��� ����(�R�%j��h(�b�]3���j"�"���%Ed��V��kd�Km���Ƞ�QDG[YP�(*%JԊQ�h�E�[�ZZ�[lJ����Ŋ�R��m�UlB�QRҪ�D�U(���-�b�q�ڕ*1��YPZ����L�֋*
�`�h���*���j4�iX��V�K[eEQeHĭX�«i@��oq���w��;U�+�Ш^9�KrJݘ��\P��йݼm��/[��=�[�U�9+�֡�ZBp�lL�V���:m����/GMڞk����8�ե���n����6�l��9�	ӞC�2f	����U�w6�ڱ��"F�Ǘg��۲ݓ��<s���<I�s�˼`�Uy��r�t�`L�n�.��N�F�s�n�9;{
�G1��H�v���c������1Q�\���6���9���oh�u�N���+;�v1�^6l�۳�,�'�X�DF����$=u��$Vsޚ��Еz%�V���J�{Im�\��n^����N�n������n�̹3�<�x��rqu2nqV
�lm55og^z0j�<I���]��l�]�����;#�Cc�Nn�"��Tq�(���ڃ�G��q5)�l��JI�ƹӱ�x�):���^����i_G&��9�7+�6NU�I�\�Fr\�x�����Z���85�Y�=cѹ�vm��z�ܼ�N�ƪܛ�;���ӎ�+�ܗ,����SjZ3ln-��d��	ls��{��қ��Rwm��'���i'�ֶM�b樹G�Ξ'�+�ݺGg���۴W��=�j�����m�g��{T݃[������������=��\�r���s�,m�r����r�9��m/a8���Y�{n�=cs�c�C�t�n;�����/�[v�H�#u��Z�t:��"	�g\s���eS���v�k����VӮ	��&:����p�ƹJ����b59;��<��}�ɮe�v����c���R�
�4;N,�����7c���'ـ�Rt�@���f5F"��z(�6w>(��W�*�����d݋'^��S�}�PM���J]�;#v����3�J��8�3���7&�[FӶ����4��S��[Ӻyy��� �Nl3r��t�;\=�7X�l����v����}<nˣc.��rkdʛ)�8�4lO^R�6�u&��)ĭ]UE�w{����6v��o�����>h^�;8���'B�Oڮ�{I�vd���Zgܓ��˅���gj���
�'5�q7v�������$5�g��m��q�ݺ{
Y{9ST������\uu�+(��<�Ν͛�	�����m�z�#�pv��Z��m���<U�T���+�|��t�(sk��k.1�tP�;x��3�Ŵ�b�'��p��X��õ�eY�m���qϔ۱�V���v������H@a�Z�?Q�!f�W��Ol�ׯk��[u7�Uta	����f��D���X�=W�T ��SYtf��,����$�ٛB�ힺ�@9�9y%�e|�%p�Yp�~�C�L�]]���ޞ���Qb_U���_ �@[��^�{�4�Jp�e"!��Q ��^N\�Ԭ����P%�v��h	��mРD>�f`HT��+<�}q/�����uy�~jETG^�D;��-]5H��w���Κ �}q�u^��a�t���O��w{%�|P ��+xF��|R9l��s ]As�ူ�n:��������߻��A@0���]WP�O�Fm�@$�D�CEN�;<�܆��U�A<#���e����ULQ$��A^}M0@�
w��.|b�GMg� �Ț�sv�`g�����;���(+؝��O�p��q���f�X�Z�-ܺS��tNhsq�S��� ��o����"�߱� ���M�x��+����3��o��ݘI��"1sQH<SFwf_��]��L:���8'f�o-���{� �ݍ��E�u6�+D?C!�8]+��(�r��1W%� s�m2" ����@ �}ݙ;;y;�ݼ�`��r����5P^��@����M=�\0O{y��ۙM������'߬�!#v׳� ��~�N�L�L�$}��T�xKxQ��y��9�d��gch�Y{�u�/��������
�E}D�'�R��L Au�M�;����171\�[�\r=�[x��L�I�u��'{���h�@"

����|t�Z62���0��u�$��nw]ߒ@$"a�N��nd����#/��US%M�cڸh��g	8��1����6���ZO��o|5b����=��ħ�т��7�Y�&]Ӊ�S�����c��W]<����)TI��9w8�ީ�bc��*��{�|�^���� u��DA=�ݙ� �U��(�)�;��qy�����9�&�^w����Nosq�B��f����1�O ���sI.GN+D?7�3R��Fgv�, >7�m�6o7���π׎� ���fg� 7��I��W�O0�j��A �Sk
X�]n�=��r����V��u���c��Zz��������QP#����\?�	�o<�@ �o��E-p)�c���m Oovf ��r���E}A2��9���+����pg٧&�I(�޻$�B'��Ixn�����ߟ���b���)��	��'�;1`�)��l ������Zݍ���H��� B���?2���ED�TM��}_M�49��^�s����@ ���m *����L�c����Q>��ݱ�����	>s��0l=���F�\��t�A�ֽ<Yu�o��f�w6X���a�Ub�we�}�����n���Y0���Q��"��� ������{rm�x�;33)�sl�UwS���޼��/�>o����Y��8�:;Z��N�y�c��,/]n��7OH-/1�^�z7���~���GK*w�gv�`| )��` Wu����ؼ���d��٘���-NM�6�`�߹�Na?�:~o��z������H��{�� |UwS`$RC8��/\L�d�=��ҩ���W�����9�"*��p�@ݺ��w/q���|)~��U�M����@�%�$§��@6�:�y�����s�o�	 W��0 ���K8�!%Q�SQ0����&��F��j��b���¯6�`�DN�sň�FIs�[���9�$>ʚ�H$���U�$"��� �:��"��'G9�N�3��R��z����IwN��&ym�v�����7���E#]]���V�n�4m�1����V����L0La�w�%Nc��8g��{s�=�(�[n-s�n0e&���ӻ<�qL��M��v�nAdD�옘�s����nڎR���n�����Z,����N�w[.�H��E�<�lT�������\A���C��PV�#���ЮĮ�p\t�q�䶶kes[�n,��p�ri�3�<�72��uI9��C��bۮ�c�&��F�ѭ����l�g���n�¹���]�^��(�cw�|#߁-���r�d����  �s{�0"���۩�*���dDu�6����)M�jT:h���q��]n��hk;=x��U��p� ';���^0�2-�.}p�,����l!0�������x� @����t���}Q�w�l @)�ko�>�[c�ED���I-�K�پ���?I��	�ڸ� ������R�^����k]l�XD�?{���_XP��$ XP���>���@���L����������}>�[��}=��Ȍ�����ϦQ�^>�c�f^2�C�G ��Oo=ss��9���"�r�|��~m�7m&�7������`��M{k�L'����� R�n�B�Dl�d���ӽ���$����"Ј"�����4goݶ����Ii}��u��R��Mau&3k<��*�l��6�A�P+d���lX{zy����}VxB8=�ow�ͭ^����_/���u�������x� R�[�h�����}��H�r�'u(t�3�w` ��[I�~gUD��7z��;���s��0 ����50����5.�����[.���� ���Ł�	 �_��H""���Z0s<��eDe�	-&ލ����4�RK�y��0 +��q�흌�Y�n�و���� ��� A��m��/�������H�<a�1~M2��ԣkv���;��PI��[��u�s�ѹ�T~}�߉�ch0�aC���O��@�=퐀p���IwI�����w���d�Iy�飦���q�XƓE���=	���6w��}�I�rV{u�� �_���}(�J�v���Kt���`	,G0"0�-$^)�;}ۢ�$��^�$A���z#9�����p;�^���-��u��:o?w����o��1�>��{�}�g%�[;D��{��Yi�[���ݗr0�a�����Fng�H�"{�k�$��:�XM��bF8.����'u�Gv��銜pI͹��U��0 ����Bꮷ�wQH��4Nȍ��L0p�	��a$'�y�î3�޿k���!��m �7q�BA$#{z����������MƙL�g�6z�v�B���j����9Ng���c���SR)����B�R�J�$�|)���EW�[������A]�T����.�5 Ut�!�t9*��R���;3��.~��_?f']w�| 
�������� O�2�1S1����^�vCz#��2�H��_E����<K  �e���U�M�W�� �WO�� >��vf|�ZC��$���,�˺�)��;�^�%��r|N��dF )��+kT�����:Z����r�+���#Z��ߕ5~]����+NN�ge괏���PHk�����TX�2)��O�/���&���9��tmP�����$CSPD�ԩu�?y���
^���76�����T��h��lh '�ݙ�����!Z�C뾇r��nx X�(�@6�`�=yV�j(@g�����v��uF�݀y�\���j���u�<�}dC	�w<� (����Y���q���T���:�$ףs���f���@L�)lS����+�����ͩ�4�wfb )}Ͳ����'���2���Q9�����,$$*}�wg�K� ʽ;��5����^� '���� ���pױ���"���f��l+��%s��d{�
~�y��(���> ���x`��Ą��>뻴��#x!p�I�BaT�s�2p$�o�hTggV;]=U�y;�D�
_s���*�zړn-׵�7�+5�|e��Oז2q�o1������{�����J(��<j�􃳔��W�u�s}R��J�F<�o�NLy�Va׹O� �"����%�ˁ�U�����W�0nѹV�l���:�����m�y�7	�p�uѣh�t���[�n�Y�^�����]�#��ʝ�Z�lޜCk�9��VLgn���`����{u�fy�g��[-��J�Kbǫ���ɤM�� lȍ��v��6ۚ�Z������gq�n �I�W�����v��g��ێ��w`l׶ɼ���j	N�A������ݺښ�s�ۛ�۩8�2O&���y*!�&�vky�p�%����<8�M5��{�d �o���� |�����꼭ʟ�;;����� ����j檨!T!�}>i�G��̅^�owgy��	 
_m� ���dC�A�^����vnp
�ssR�R���I-�O���H^�iȀA鰏^L��u=��
_kl� Ut�jB�a��Q_T� 	��}����9�:��Mw] >��2h$�M�d�H�_w]���������'#�&Br�f���16�!��}M0@ ���3]�;��7�Q[m�@ ���7�@��s{�8��O��
z Y)���	 /���� �v�\���f��盲u�q���u����F���y7��3%!�$�gy�0�v�`s���$�IUs��ȅ�5F��h$[ݫ`}�2�*�h�R陾��� 2�/O>��(�VK<a��Lc$��bkf���oj�My�5u9����[�w��r�}��P@��s��S�%z����T�ҭQbH�����w*�~�M�9&	Nw�������n^�Ͼ������>&�B���� O{���dw�u���e{� -���H8���1 �-�%AQ*�@�e�O�y��M?n5	�Q���0 ���ɿ$�s��r*β�ĝ�Il�:&��C�¢��R@�w;٘ _Nە8�K8ɽ��a%];4I����Q6�_O7#�o��7��T����E*��HwAv��1�n�nztc>.�z�3�N�T��ܽ�L!P��RG�c�i�=[����_W1�!��U�_÷����ջ��f��C���������c��r'+�ў}�z���e��$����π@"��6��'2ӽ����>Nm���f��pHeCNS3}}Z- |�z܇� ��_��ҳ{֯�����Y�f{��+=�+���������&��}�k:_�����`����rL1^�w�e���W��J>6+I{gÞK6p�<�^hqy�,�Ѱ⠋�}���`���4�s����˫.��U�l���&0B�u�����h��sYoyg�����RoN=���xIOL5Q���o��c�����|<����)nr�T�ʈDv�q�����~�/��u��6 ����|��1qNd"H��]�PW�ov���0��ܭŏ6�w�؜�\�B��t�L/A��ך�����T�k҇��+�fCK,���g���e9�4�!�ӗ^�P�n.�������0�~��x�S~�����%\V���m���J^���#�A����'d8��ػ ���K��?��w�]������l��~^�sg�Wr"q��DuH컇B�1�u:ѽ��+l(��v�q:���%���L�÷���7�ΞfP�{}u�S�������g=�6>�~��pyv�R��l��-YIf1G	n�!8=��r�wTŤ�k�]��l�������^�����B�κ�<�Yʍ+��zvhս���>����,ўx;��R�Ý�i̘3��ox1v$�{�<�:���}zA�P�,n��[S�'ǻ���<��(���$��f$'l7�=Fo����A'�HEZ��op=�� ߽�L�7�(4L�G���ޝ��'���Z���G[��w�M��~��Y��Ǆ��j�ýV��)�ڛms<��H�b0^5e��DE"5(�m-[J�Kmy�\���-�NaZ�Z�h�-k��\�ư[B��QQQX* ���PV�D�M6:h"Db*:���U����m��F�Ƹʊ
�UE��*J��iZ ����iT[J��m���QQ�[�l�M4DH�bԪ6DU���F։j�b1TE*
%V�QKk-�n2�Q���"�Z�ت(� �V�ck*�Q��[Zэj(�KB�Zf\�XU�U�E��B�,F��*%�E�%lQ(�l�B�-��k�b��*5ZEPF�Q�5�+)YYF����UD)J-�`��R�m��b����P�V�(�)U���X���[F���Z5UKaDڥh�ZV����%b��Pf5�*�X���U����+F�)h��[kKQ�Ū�1�UEb����kiUV�j��E�Z�[k-��������J�U�\qDPb�R�Zv�_s�����|���3�!���檔T)*�v�z�7�Y.�V��c��  >�:�0��r��n�6���&`����]ߒW����q�xCP��$�'n��d6�:R��o9����=nH��HHJ/�������ZEa����BE�k᥮�b��6�` C�.[�M|���w�(��B� ��FVw�� +\� �_^ۆiJ���� 3}=^��0�ζ��W�L �
�RC^u\D}���sO���߯{�ƀ�U��������@b�D�����m_��NR;�"2�a���6����"I]v���2$�<��^����pDs�dC ���Dd>�U�5��f����M�e��Ó�$�뎚���u\?�@.�ofk��Fj���7�#ߠ��\���X���U{��iD���z�~z4JT:po�wW��L9�c!	��Rk7dk���ʇ��l|�/26�4�Ѫ�M@�l1���O�;�Ů�����Vw[z{�T�t�a$��r ?���ww�Q���j�@�:���o��<�K�v��gl�8��7�4� �	�C���_]c�7��~~�����9_rD��d?�D]{j�D﷛ς-�ݞ��ǞN7�� ��u6��0�D�&JW�u�]�I+	�1f�����#��|����@ '}����o�Bo������LT�%wfw�Ra�pa��ֺ�I1��W�H$L�9k;fcw���@'_|�$ qz���$���M��E�}���g�P5+���d  %>��f$ �y�zߋ�zb/��H����Ng�|1�F4�-���f}�
�=nC�P�5�y��ۚ���uq�����3�s�mI'w���M�����b�^���xإbA�7xov7���K��e#��ũ^Z~�ϻ7�i�+2���yV���!�?>�W&4Z������{��Ypt�6}!�6Fr�ۻ�˝�+Ӻ��_@p�,���7`��tv�3u�h�x\S�wf�rG�=v��[:��E{������W�,��類E�q=���3q�[٢1�-�Fj)�����Wll��Ogc�^�a�ȝ>L�;�{n��Ø�Y�8���;.)�1���[!�{u�[������a�wn8���خ�v�p�۳�+Xm2ƈqn{a��ڛ7m������n����ls�z�F�6S��ϻ9pl0S�PY?%���H���6|�zƂ�EY7}��V?"��m�ﻳ"1��q5T�D*��D�O7!���m��,��]6 ��}�٘�W9��<𬩌N�*���/�ɇ
&�EDJa�N�{3 ��s�Ԃ 6��E�Y��==w��$绳1�s�o�fE��W�UL��'/��T���S{���y�  }^ü`"뺙���ƫ�'��r����i�"6�a$��6a�y��>�m6,ͳ_�sb=�؃�Ǚ�� V��J� .���wI�*1��=�׈� �i����`��2��Z����[�\�+�;�l=��������J�s������i�WMy�IQ=�F�\��������f�g� W��ѱnb�DȊ�R3$��yI �����4��2���!��Z�'P�v�?[-�}��o��{�נ��麽3��{���Pnտ;Vx�&�̝���/��u�>� �U��9` ���M���Q��o��c����H�"�[%���o�M0����6���ا�y�"V��  /���gz4`L``,$�����.�n��&h�$��w8^H���p�N�{3��P9G�~0����b�߈������A���`��'���`�W���%�S���:}�X "o�M��'���|��s8w*#�}��ڶ=����;n� ��X��!����9���m~E ^,o�Z6�`������z���[���@Nv�f|�nT\�Y/�Y����O�t(�3��)�������(-m y�w���m�@ 
�:�4s��"1��ʪ��96��<��($QS@�A��M�>��� �7�6"�>/���:��mӿprg�}}�0�̹wy����|7�g�
����˟���O0M����qgo���E��e�[}�������o7�� �S �;fDW-���*U"�I�%��A7xV���^DjA���`�	��7� \g\b��Ὰ �'0͟8��*�c�(	��c�� �m�F��B�Is�=}�p�N��f|\g7Be��>P}��*2�Ł�CH��N3��p���kb&�[<\�.fa����[�-SY]w�{���c�Z��O�k�`��y�@*��9i'$�8鵎��&�@k��I{Q���M��/���Ǭ���v{��o�s2��X� ��ovf �
�����й�=��;����҅��[��M*t�7��f,�+Ou� V�j���E��x�@uv�dF >+�sj�in��$�)MD�}�����St���׋�	����`�������۫­�y�=�S���ໃ�3�����z�*�=7����^���[ɽ����o��jp�R��b�*/U�t�����C�wc�*�b�� �?�����~4�p��RKh�~�Ң Aw��f�S�D?�s��� 	ӵ�  ���wq�{.�}�N�z��UD�����/n�;�v�u����id݋��76�tn@�������cO�K&Jr���`Z^H�ջ4�]�U�Au7Y1Y~�;����| Dr�5�a�p|Yn!%T���&��fr�d��	B����o0"tݹ�a}�m ��G��6���`�=٨
GP���O@�3a�ݻ��I/�n���3�j����ݹ�"cw[�	Jg��5��Hna���:���ۛ�f�^�ۿ ��om�����p�@ >����%�7ʮ���@�o?i�{c ��`������	$�{�,-�:��=qur���u���=��V�fD=���ɫ��۲��Wok��5:��B��=�����vŞ.�2=�G�QKZX��\U�4hZ�t�TA7���ˬ�Fjُ�}����������^Ռ5��W��v��ŷg��rX���GR�<���960�Њ����I�xN*]R�n�ݭZ�v�VM��N�8��S�oY�Н��;Wt4�sغ}\�[0<��v��$'R�`�{k�n��l0)�Hݽm�:n�l������5�Zm��c�wϟ7l<�%��":ؓ��k8�M��m�mN��O><�+vwd;m��ݘׅ����4Y���;�&��n�uq���B^�rv� ;��52s������=q�9�"a�����\?�@Nwvf F��pG=���/Ϫ��Y�f�DJ�E &-��vbX m�Uӕ�������q�����@ �a�^�YB�w��������0�H�0��� w����j��-��S�u�Q���m �9�ٙ�#މ#�U3Jf`�;�;��3�6Πnn��A$"���l�*1���=�	8zo�O��C<���M�t��ۿZA"`�dԡXym\ ݠ[{�F��1��Ua"Lrܚh�S�l��_���ri���m��l�n�r-����]�wN7] �"$��@c��k. ��
��{\��>�sϰD
zw�XY�9n���a�d�"���go]�I��ߜ�DL)��,�s�ن�}�j��;���\�\+Tò���y�Zo�]��:�m������Ob��ۡ�<k'}�=�OD�G��i������_ģާ/�r ����� 	�|ڢ �2�=�}����G�� X�2L6�o{3 �O� ���%��vb ��ݙ� ��}mPgyz,h��I!/j�����~���g�%��};�, /���Q9�fnY�ݼ&sϾ��|�Zi<����홧�ڠ�����֊�<�}��� ��;�� ���ԑ&�n��������PX�0c	�����-srz���&��\[�p��]����˅�z��7��w}�ul�9{�]iy$�]�M �*g�R'f�������ׯ�[��n�h=��JË7���ˮD1���U�U33���`�	N�y��������&�{�=�#m��꽼��Z�ڪ��j"aH�����@ ]�zƀ�,�C�r��#�k�r�5�d��ב�~�1R��^QB��'8�w٫{z��˫`B߰z��"��Y�p{[�7����ً���+��I䒎]�^h����<ڐ��.�����(�&D���ͮ퍑�"�cl��<{o�"��cHD�"���Dm�w�=U�5$ҽ�43�,h��I!.����}��\S�8����7��	��r�@"�'�RA�Nwsq�6ݺ���5T�PG����n;x.���6�F�sv�p93Qt�kmcu���4Zx�7�>��&2I$���r Nwvf ���2G����H� �ڽ"'�<L#>xa�����s���J�ǎ:�yv��D��t�i%��dߒ��R:7v�1�z��h床�T)T�R������@�}��>�"#۪����evN��{:��@�{�vM�xl�o� 1B���)v�=�%�3|`�I����%$�sz�I�)L�+�3�	�F�?.�n�
U������ӂ���w]���\Gޣ٦l�b짠�=�L^Tng�5>��Y�I��1�al�)X�n�qY��V��{�I�k��I{����J@���"x�[�U�y�8�z�� �r�� 
3�������eSCe3Ѥ#y��g~n��ِ�,뎜`��qA�9��q@nH����mL��C-br}��!/���D߉}��1�'w��� ==�,;+��R�qP�9��M$�vo]�KI�0���x��|m�$�|�q�n��s|��fg��z�36ɗ�(��b�iR#�-2�lӯ+���@|�n��2����yzr@ '7�3 @�y��z�EA*�PU4��ʷ��{�x�<&��������D��ܨ&�IL�uf^�s��y$6�=��+ն�W�2�c���,�mQ�GP��=w._QU�v<����M����D率�~]t���a�FG1fd�s�n�;C�,=�6c#y��-���~I������G��d���M���n>}+ݝ�}��s�������_����\�..���9�y�w"pnn�Y:XH�ʜ"w.Nʈ�N�^��o�9���w4J����y��f�A��G��l֖��]1Oz�,��.�=Tg�|,������J0�A[���rv
I��ك7�ÉҸ`ʟo�f���1���d�<��O����9Ok�s�w����S�ؼ@ݨZ��%*E(�;;�3%Fm��b�0�<;��;N����ZQ�-�{�>�Zbز����i.�����n{���s˷6�$g�����<]đ�j��H�w9�yuf�6!���c�*[��l�ts�nM\�.8f,��hQ{����Y��G�����q�s6�L�p'��sb��yI�[��G�y��$'v3�Q�ye�`�����E"�E�p�~�6v՝z��{��{�ǭ{^G�r��Sa�El�?<ޞy=oU�7Zz�Í��sIg�J\������=��������5�����0�s��ò�^~���Y�v����ܢi�P�~|�᧵��s�����Iԗ�9!�������̓�Ղ������'<O��2�K�3��"�;<��dM��_xO@^���dղo_`��G�z�w�[�y�^�D�ev�`��E+/��i�-v��#���.��Xxǳ���*�{Gg���r��ؕk��}}���5M�����ӳ=�p�N��mV�X�oh=�l��Й��������T��Ԣ�lQl�+ij%�ڥVҨU���m���(��j�jԨ��ڈ��im���jKj����3�kj6�4mHZYmb�Q��*�T�����J֠������Vэ�b��F�
�R�lkbA`�[Pm(4�Kj��E�ҹq�ATm**�U(��
Z0Q�m*ň*�Tm�-������ʥeKeEm��
��PP����`���V�UZ��k*Ŗ� �[V"�m-V֡[�V���	X5�R�"��T���Z�Q�jUm�YmcRUj�J�b��(�s2`[V5��m-A#hUAe�b�PUZ��������l�EYm��Jc�-�U��F�F�Ҩ��UP�B�h�F��b���ڋm Ƥh��,m�m��Ԫ�bԱ�0��eB֋J�0H�ZT����Aj)E���X�j�Dm%`�EF����b6�loxߟ8��V*�l��UƗT��g��]���mB�eu�]['q��{%����l�ޠ;]	���UFn!v��ܖ蓷�{��v��n��a�\����I��g�m�d7=:HM����M�d���@>T���]a1�ηi��jr=�S�kqu����g��_5���nM�[9�vN�&�c'���{fύ�����tK��.D�v�9Q]�u04R�QQ՚ˤ��3�+��\�����[������Omr��¹�>��b�lK�R]�q�p�k���|τ�9��K��..G�L6��u��<;��6��a�2y���kN�kÞ:�cV�]�������v���ۮ=L�f�X���k�u�=��W���"���zOX5\�x���W
b�{\9��Z�z8�iݓ���ض�N�Z�<�
K�m��>��=��j4
<b��X!����^��۞�;8���|���'���2p[{`���{{=����h��Fr���uɲ�۳����/\���:��ogf:�v�ڱ��̻mu�A�n�c�+�0[v��	�z��ه�]���X��Q�y�ܝ�����ӡ{-�5��ۢ_cq���iE���Sb��'Q/%��<i;c+���{YGn�6��'����[s�ZĎ�X���.�z�yA��9�!�#�˴(�rc�7n���	���vRx���$%ջs͝���� �����mO��/kO��άm�@a9@K�X�;M-�Y�}[u��˓��Y�j4LU]u��pg�͜=�����Q������qm�[�	9��1��.��q�m��i�7�n�rѺH�歳�vݿ��>|�q�wY�����v��#|�۩�aG�m�<�<,lun�c��:�,�û�a���)�϶�=vzݮ��`snb�Y����vB4���Ghf��멗��Pk��mq��j���u�s�Z��E��/��;t��6�7��4򝲗`d3�!`�����ڴ��J��H��Gnڣ3MU����=����v�1u�]��8��'9�1iy��{jm�죐U�'�+�t<�t�u�����,'%�^��L�����F|�N��;v5���H����;w8|s�X�������wI�e��Ϝ��\f�΢1��7n5��9W�n�Bq��'\g�&�9B*�u�nq�N�#1��J��;�r�$v����p�K[��wnq�m�cs78cRK�%Bʚ�b$����9�p�vfy��0qr�p�k������}R@�D����@龶� 	w��h!�D��w�Q�~��zN�I'
���%��!/���D�������Z�1�{����I^_X� w�ͥ$&���O��v�G�a4�4tw�v�I'	��zDI�o�]��;�/u$ �;T@��GR41ZT��Y��u�w���nz��Ek��'�v�.�>�� _k����ћYt �=)#��&���i��T)T�R.���7 :�y��GJ�_�5�T�l�ս^O��@ ]��B($���&�E�LJ̶#��T��qu�\J[9ܚ�۷	Hq�v8�^,�y�\���o����Bg��y$��^�$�y߾��M�r��iuV~.�� L$�;�z7��he�IBR�w�D�CY��ځ�S�
��AQl�i,��[����(W+/�{CMw*X^���O�Ķ>�v���:��2����k˭��}�{!Ⱦ�^݌|�~��������|��k@|���߻2#hlޚ����A/o���f	�
���q띳� �V�<��{�(c71��Z'H)����+�w^bi�FTMM)����gz|�c�*O�� |Ny��@ >����@|��v���\�$���4�f�
**%L�tљ��� ��[�T׽�]��G(ֻ`$�K�D�QݽwiW�.�0�|�*�#��ac_�%Wb�-;�&�D.�n9�z3�5�Ưd�����������L 0�y'�U$Ln�U�| Ouc�F�>��/cQ�s��i>�����m����U1�Il��ڨDʹ�3����N���uz��Q��� >�{�RA�v�Zl�;5����� ��e�EÃ���A�蹯BI$�-��s��i�Od�� ���u{Ȱ7!����C�{8'����ޏ���;��{��	��3iK;����>{"w=��;)��?�2޿3� '�~��$�{���u3CmBJ�,���ظ�8w�Q,%}�0 �	ެcA}<�:㕳wbtBm����x�9����h���� 
��iʷt�Q߻�1��g�"���nM�&h�Y��sA�߲x�l�ìuF�m����۱�}678�g-���3($��]��c�i�`D1O����1` �9m)�
����٩7�u�:<z���$��v�D�;� ���JU!������r���!N5f>���  %;Ռ@U��rDF�meu��}Xۈ����Q
�T��Im�^� ����G� nk��>��q���� '�q��� �W�ͩy��(��RR &'��KW�>���<πH<�}d0�����s��̨'E��s]{?.^i���ݷ��W/~���9h��Y��!�s�s�_\ޜcFܽOu��H2D�{.^a!�4@-�ۻ��n2o���f�@$u��jAv�`��ĩ�UTH�y�X�HQ��U�����}���K.�$�/�R` U��"w�٘����Ô�����뿑��\m�՝�!�9퇞�pm��@�����(�@��my=??�7풝Z���j���I���&�I��b��j��7o���H� ��}"4q3_`e�$�\����vh���{6n�� �W�� �w����|
��{"�O��!�;�Z�م��J�q=9��<��k�m�3�׌H�����r@�S����-�T�jD!
*���6�tqBs:��R!�9��rD�o7�  �����F�]3�[�ې��%�*���	���}�� H'�9mI��d���E�~��|緳"0N��rWlǶ�EH���c��ﲋw˵d�w�𸚫����ݓ��ڸ��y>��8Gk�l���V�X�ll-�L}�(�Q	dv���+�7m��Y^!�<�i�����X�_������s�#�|��N<m9J��8���i7^N^�E�{>��z;5v`ڴF��]��q�'v7t�=�=	�p���SeT��m��#�!ɒW8�;v���b�L���';R�\�Ҏ�<3�/���q��/n��*�Ŏ&Ν���������NN��
��!�y[��]�q�sf9�����-�X��&��}T�랜4ݹ�+�_����٣���%��
U�%Q�P�Q��y������0�?\:�5���7�-�$	>�vf|0�2�*�*����3:|�aK�#ݘ�D?\�r Q۽w~I$cz.kЊK]�|�doFMz}�������h�3I�Fgv�%� Ol��Q��U��Uv����f` |�ޜd=<^TI10M@E�WO��[3���8� <���� @}=��`�W�Ϯ�d�z/۰�N�����m���L)��D�/B ��{W�O�+��.�K�[�&��uD�V�T��H��t�,�=o�Ӫ�~ݿ>c�o���&�����ػQ�����z��;��\9��������;S��&=��>�XDDO�r��A ����4����
j*[����"Lv��z�vB)@���AJ�Ș�I�L������F�v�E,�v���H�B*nn"�P���2���V�ul��g�W���n���#;_?7��������Y}��  O���D?�E���"I�{�o�����[����4� [a�Y7q��}@�Awӯ� 	�LR�=P�ڞ�'1˲k�����	{�z�銥%'L��n]��x�m�`_���]@	���� BW}���������k?����L���$�����J�P^^L`��@gNk�� "��������f`ef���9������j����Y��g�[�:;ut�xI�7m��;v��\�߿�������[���Qڹd�	L�m
�I���Iل���xx�����"]��r	�a5U0B/%	
�O��q9����.Y��-��;-� ���1�ӝݙ� �1/}���W��f����9Xq �i[S��!���<XD3���ݭgrj����o+E�.�k�U�ԴWuA��}�|߾��Z]��{��읹��=Y�p��wu�N����������is_�AL�m"i%��d��
E��a�X���Ģ�q���D���K�OX��'�y�A�ux߳j*j=ѱ���̆���v�鉨���f�u߭$�I�ܖt�T��!�lŘx����;�٘�"��ͫ:6Gl���ܙK��8)�""	d`C瓶�Q��ۚ�.����Y8�Q�L�la������ds�Q�'�>iȂ"}��>� ����{���2l�Eק��A=������������"��P�����3�7�T��9�c��@$�����Tn��de�<Y�wj�+W�v|ڐ{�L'QS!J`&�߰>G��Ց�^T�O,=.�?��	�wfb >*;����,�P�"��f��9�;��3�[(�����Q���利_{�xs�؟DQ�W��|kӹ��i�ÚS�yq~�c�,��Y^I�V>��g<ܳv��4t{�yaÐ'�q^��fo�OܘlLDr^x�3>Ǘ�P0*iMQ@�2�����[�S��'sE��#�{����w�� ����d���q�+����X����n�o��.z���ⳝa��ٟVZ�C�.̵�p�/_���~q��=f�cynfuش��,��ԤD��t�ZeU�';b��ۻ&��g�&�-X�,"�0HdM �ˬG	�Y���/�f��q��t��"率�HV�F�7d��ٱ��K�A�Q���d@~����/�]��h瞼� �����I�/��;�/�cA"^ J��/�1�T�,���1�+�+�ݑ }Z�ӛ��g��{�뜰8tw��nq���X���5����DN��ϰ���3ir�̎�����@$�ߧ[� ������_��w�����{��}`��.�~�`qg���[ֽ�Ǹ�!�����q"�9��9�4�ϔ4L��\��Gq�|���$�{7[e�pu��m���:�ɨ쵊{k�m��Վ'{cm���>f� {r
�v�tv�46�c��"�p�um�-sx���['�3#�'<���+um��=b�e�6Pn���Wl���I���]��:�v�Nݬ��Z��*^�s�r���\��b�۩��T[SWt������tk��痥�v�z�8����n1�K�V�9�
Q���[A!�v�'#�p�v�֍wn�_�u�un���5���w�x���� �|�q��n�E�ο��9����)Cqٷ��J�����oi �U�6"""v�ꉨ��陾��ޞ{=>HWA5�\[��w��D?�s��π@�vE������/��`��L��E'm�O��D������\ןK���U���E�O��"9�٘�6!�Siy�0��=[=�=3�Fչ����>i��N�vf ���b��d��E���^Q�U�		���CU12��0�/{3>�� ��zڲ�zI��"h%s�r�"T^o]�D����3J�X�b��<1��4O���.��3�tҹ�\�F��v�m����wL��߽�w�T��UET�#��zȆ�ww�`| 
��:i���븝�؉Z�[� ��������J��EQ@��u�v�{�L�/{���B���R�<$�8��R�]��g��-O���=P���.�X�(F�ݞ�C�ٺ����vf��q�ۚ��9�s{�π@�o� H:1f���OY�d��'�D��
N�7=X Go��`�A[}Q�U~�xy �s�٘�@|���9�����"�Lɠr�uá]kޙF ���q� �uʾ�l�/���Ũ���/�Iy����IN��.^aQE���JI�GP��]�����2=�,��fg�|EG�΢�}<ڑFIي�O�gd��T�rNK���zm���A�۵�ja�v�D>����u�)o�g��S!_I�o� *=�5(�s�ҫ�<��w����ݹwi �	��𕝃��@e��ג�9朁�.7�wUy�{���D Q��L.�y�$DEY}>��o|���eKOe�6a���� o��  ��GL����@)�	sڰ�V�Z���{�,;�G�o�����7{�ꌧ���p���^���M��9��)ϸ��΁�$]��q�_??{s)��loZ��z^�C�<�T�R<fuy;v5DG�V1؞�������ޯ	��8�� ��x0\ܫ��wwn!=���D��<��i|*�X��݅���+ج�{m^�	�z��ٖ��w�{�¢��(J��	WJE_t�nV��P��{���f��M޾>Ь��]�����G�����,@{�;��bi�SnnR}t5����1���{����Ϯ��n�g��HF鹰�wU`�b�����܀��n��W����i�K�s}9���wT7�ox{�||�/zз��(�)�Ӗ��]�M�}�]9=�y.=W��Ћ�����\����n�u�3�q��mh>��o�C2�Qї�����W�C,ɸ���tl�+����S��s:��J �z\��DB�7gF����S�"��l�o#�y��1<��&�o�w�7=�[��%P���p��g�!�`Qz��]�����5�Y��3N�C�/l�2Io������a��ץ�z���2E���[���*�;u@rᗗS�@N�4q�=���#�X���z�v)�ud˺�2����xs�M�ע���=��F��dC��.�Gn���!<Q������H���ot�w/h_�N9;���->�&�+�+\�"ۃu�ކ�9�Q�\[��sס��������ف:�!�w���_��>x�E�o¾�KF�[k*��R�*�TV+nҦ1�J��*�d�+mյ�F���KiFTm!TX�q��b6ԵJVTk(�,T�(�)*4�%E���"֠�Kj�ڥ�h��Bѵ��1b�[l�bV�b�TZ��Ԥ�$��,kEkm�ՋR�VTT����LL`cA���Q�J
�,j-EX��H�
"��[-*�[KE�Jԥh�6����Yj,U��m(�(�Q*J��ڴU�jZXʕP�--�V*
Ɩ�5�5�++EVҌ�R)e+kKm��V�aKj�յih�e��m�W*�KQ��E�
4�Z�ZX��AElFV�-���X ���T��[ikR����ک
#d��� Q��iY@"率�����p��-�LS7�]X!�%l�:�|E^�V���D?�S���q�f�����G��<4�d�%Q���+g�0O�������{�<Vy�C�"��D4��fb���Z&M��y"0���Z/
Ƃ\�<��pTZ����G�O*�,�y�\XX������ͭ*��$�"a�6���N�� ��z엯!oS�@,3�U(���r:����Ppb~�`�(�뻴H��#�Q�d϶7� .�v� Nv�f ��������=Ď��Iη���UR���|=n����7�{n�9���|Sˬ��Dfy����޻�$���Q�bM�
���̨����V��z� �Zt| 
}�ٖ�I�vV���`��oJ��\���/{���KT�gI<?X�����{=�+�t~ �M�]Z��<'��l-���o�3,��z<G z��Ҡ]�C]54W�UL�F>|�h+�e�B�r���o���=�_����1 �+��j�վkUPn���3$%S��q9֍�l:�#���P��s��5z���GÀ��-��K$�-��"cw��Z%$��:�)*xg�w:�Pe�!��t@�J{��1 巊j*
��T��[D��� ̬ǯ6C�ܽ�; ����f  +���2=\�X��j/��D�B/Ќ����3��
�r� \�����#�*�����!��w�"0��n����D�
UET�!����s^���w�;׏�+����;�Z�A�/7�p������w��V	<-��ه�#*�$IL����Pv�fv�0�/o"3�
�N7$ ����GnVF�*����ó�=��x��2Sf&ly���t0N����11&�6l_N��S�	��!��f�}:�iz7�w2�jX�d��������D<Xc/k�Da/]�(:��M�.�+8cՎ�r���g�<��[�����[�W�ݸ��P\����=v�D��MOl�=Z�lV�Ykv�L�Ux����ʤ���k��zf��G	�"�F%�Qۮ�p�!���`vo\Rnv�Jh���یX�J���[2�v�Ywc�N���rC��*���p8��b(�˷��7��.�p\��рȦK7m�^܈ӱ�ێ�ngn�y���7/f��7�n������54W�UL�w�ggc�{�,��@+��r��Y��U-�����s0 �|��Ȝ��
E��ɰ�g�1��N�����nw���G$�>��.���uW��ߡ����1����a��6���
�/I��	�7��3�6C��]�=��>� '�|Ȇ.���湙��I�J�p__:�쪲;m�vj�{=mH|]�s�$���ft�F"�j9D7����٘����2����" ���J��U�ip�y+�=�|�ȹU�H̫�iQs{�1{3�p�u�,��N�6׎�@��%��= n�g#��`�Ɂk;.nv���z}��9�a'������ڬ��$Eپi: A9���u� ��TG�o�����~�L���am���/#����L��}`���n���Ф���/�'��w�����VGz|PE��EcD����v�cc+��f&�fZ��ӖeS�}��<l-����_jsg��w�d��� s�倐����߱]0o�{�[{�'�q��
H V2 x��;�:> '����]J�b�"�DSͱ�Afu�DD
sw�0	���6S@��J+�ktٽ7�7�9�x���: ��vf ]����w��q+����U=���X�`��#� ;魯�� ;�{���Nd���dNTRD��޻&�A=��E��k�p/g��@$?�cƞ)��7r�N�>�s�9�MU�9���j~pg��&�߽���&�*��T��|�t|ӣ�{w�|� Oy�*�C*�X˼�����7�(b�{��'=r��"a'���ݘ{�VLA�wW;����r;�  S��̈πEoO�R@����y�bM�������� �̖�y�{��tI�_�VhBA$V��}:����k���y�7���/������"{9�_hoq����h�#_��9/8��Kù"��ڳ0v2���giN���7W$�N{y���EoO�i�%�3$�B�N���QN�u�q�h�~n1�H<ה���	�GT��n	�S�;Y�_��7�~T�J&
�&1$��=����W��>�վ������n����$+�>dC���r[f���v#����|�T`9�z$��'W16%g]m�6�Lf�Nu��g4�>�}�#vy�q;��� �l�  ���0͎޻�,p���I��΋����4� b�X��	V/�dD�}t� q������ W������m) 	�κu�"c��ov�m�o�CpZ��6&j"�j&��gz|�R �O� �Y���H��w}���| wN6�� ��o�b��U�LUC������j�Q>+@A���Ґ��W1��Iz77��A'Xo�V`�KMi�̙m�ݼ����NAf�Χ��'2��ۏ6�v�۝ǧ�~�.����ɝ:{���d���j7���b��q�Pə��J!E+��et�ƀ	�w<X=��Ō[~�Ĝ��C	 �ݫ� �ﻀ������^���~m�
ebă|�f�[�>�z͓j� ��Pu�;6�۬�rV9�;���4LTL"bI�/g,���N��W����}�!���������aw�ͩ�5̧EHQ
%L6��������0Kˬ�d�Y�虿BA$Bg�X�O{{3,�����Q׸]M�3�@�BPce�$HJ�}3"?�>��� e��D=O�LM��x������ ���x����P�R����
l=�V{Q�>��Ef�/?Ĝ'ί�T�Q��wi�}�u����������f"r��1��-�sw��wI%ߗi��~�Լ�����UѠ
ww�0 [Ӎ��fMd�D�?k�a�փ�s���{�lc����Vn���wZ���GpZ!��Wy���	=���3Bo	���/���b�^�r⅏xb�
����,(��&����v�s�ڕ��� wE�9�m��8���@F�]�t-�x�F��g�,Z��7�u��z�9-N፞܏*��Gm���A����9x�ܽ�{Wl����8�ͪ0t뫞��D�`�i��Űm���������˞��Ӹ���{j�7M�6��E����:��Ž=����tu�8��u�Ka0n��n�ƹ�X.�v�/&v��@�݄a��mš�]����'�*ۖն(��䞩x��E&F�~�U�" 	�w<X����0=y����{ބ�7��
}������{3D�UD�&$��%��iH�2���ࢧ��=9 �c;���^I���"J���K���.>^�����#-�H�X�ӛq��9nH��Z��'%���`���vA$ދ��$2��1IA&1�� j�������};�Ā��� 
��� ���1��5�iC@w�w3F��R������l�Ud�D� =�Y�5�kG� 	�߮f`�9nH E_O6����G)ϧ�Ϯ������m�f�vnzƶcc�;�.Ź)��&�������ܽ~�}���u���~W#s�ى` �Ӗԑ}=cA�O�����3���� �SH��-) �P���	E�e
�w�n³�R승��뫳�������bə�i+ݣ���[�j�02w��s����Em;�ɔ�]91�C�K8+�a��]�>n�jÙ5$^��r�$�O�.Q$�Nz:�B+�<3�[��$�\+j
uD�&$��%��j@~�i�@��o�B��d6����@ 
�nH����ޅH��8!!_w�ߘ�u�Ek��e�0�d�܀W��4���g�vɭqA��8ڐ[���K
 ,i�2�_i�I%_{��~�$��y�z��"�gͥ$;��w��AnN���I��6�(��c�	xݱ�T��c�z�.W�짶7]���6�5�����F|�$�i0���꬟� �+"$�P���	? ]��W
G�6�$�ѓ�"pA�?,_�%!�/��HM\�����_MM���k��D����	ʽ��pЏܻ��}��R)20<�0�~VDI}~�AĀ�o��ٯf�syow����<y��'��A����������z�'6֢����~b[��7�c����}�kB:z�u�g��ս���Vg�@/�H���I 	N�{2#���LTT"bIo�_N�|t��`|�q� ���Ȍ ���W.�_���2`$���GR4�҃E��M#�b�}�ٜ@$���b:�w޳��V '�ݙ�$Wt������m/�	��~i��b�NpN˫��ݫZ.����cvr���^���R_??��I$D�����ܐN�Z�w�` ����4rQgT���T@���������JJ����tѝ��r	/����������ݙ���8ڒ"+nT����پJ��FɟR��EL���3��0>��N[R	 �8�Vj��;����`����$_�.�O���	20<�#�T\5�׌^�N{9�� >���4 ����������u�&	C�����!���Fn8��E�}gn�вe"��(�CG`��u[;��_}���uP_�XG_Gué	��vL�����o{3 ���B�
��DĒ�ľ�n@g��&��ݯuzoٱ�{s"3�+�8ڒ.���T]�����ߛU>9ۤ@��t�N���P�0vk�@���v6���.[�v�>�w���U�{J��'3�`n�[�w=�b8�ی��5�z ����>�tA��$�4�FOĪgڡ78o��ҹ��YF���� oV1�E��o� Ab�ʷN��uݷ۸�� ωt���&�u�9~R ��\��J��.;7�/�$�	���$�S+��y���I�UEASC�fnvK�fu��D� o\�jH���}�-�N�y����#�߉?���"?d"�20<����t �{������d�������n� ���dF��v��ۿK���޷.=�'����a{�7�8�w̻��#�(@��ʪ�ܛ9����w�xЕ輄����.�!wy�����ox�y��l��[�|����.(��껷���Wl7�x���@=>��"%3.�������E��u��~��"G�j3t��<Eu��]�Fm��,^������{�k�5�{�$
9�R%�޾�Z�Lڡ͝���6z56N���}��������}�wR�Ní�{��NqbcHf�Yod #�l����x&�q���;�@�b�S<��4�3��駟�T�\�]�%������� 5�{Y���Q>+|{y�y�[�˳E���swֿ�YH���Y���pgV��a%�1�,���cW|�����&�o�#�x�f���1�$�� 	w"Zp��:mW}=��\P�e�V�7���+���zK,�|%����2g�:��l�Q��n���g�x���t䟭��<��ӻ@�iu��f���Y�����O~�I��A�&zT����+�R����^�ɗV��^�/%<B^~"I���sP�n�NoH�Z�*"�k�+wf��^12�*����9��9p;
9���r��]�e�5�Ź�O�w�}*��/x���>�͛S\'�I'�>�㻊��}�'!͞��8�S=�w�'.�L!�y���.w|��43����j��Q���&O;���sǴx��-qxx�Ƅ��o��m7{Im4sr�5w���y����miE��V���*U�cl��J��XZ�khV��ƹkF�j"�ձ��J�h(�m([
���FVږ�F� Z�-�֒�V �ƕm��J�Z5-(ֵ��*,A
Ƌ(���DH��,QekQA��ch����U�X���R�j��U�������Qm��q��5�0`�	R��)r5���K�UR�F��Tuf6˅����ҋ�5nb�(ᘨ�(�E�9�㔸�0iX�QT6�d�=����w<���v4�iV�PF��h�KZ�QUJ�D2���\)j�6�P��R��qF12�2�+.b�[kr��2�s�e1��B֨��r�T�
�,��`(eu�]1r�#FV�*��H��AUS-m���\kR�iTD�F�1�R� ��
�eX�V�Ŷ�[B�[3*+B��K-R��Ng�w��[<s�Ҿ�kqrT`��r��M�r��$���a���`�z���v<�]'��0>�c�C]�ݞ�,�:.��K<���݋�z[�}��1ˑz���Ѻ⣌�ay���0�nݭ��ն��ɪj��<5�u�.5�؂�p���+lRFa�]�G�ʷcͳq��nÅ�� ��uӚt�ܧ��.-ͳ�����u�����z֑g=�3��3�ћ�m�]p�kW`��=t��p*�2���&z��v�7�{!����k��I�{t��W<sԫ�E�'"���uv8n4q�nv��cgq��u=g/Q�=��6�!�,�a"�i٭�i�-dx�m�׶4���6���7��*�J ��)u���E�y��ˁBy0 �7mӐn^v��a�!��V�M��/\���`g��Z���c��/�f��k�c�uq��%���1�z<�㝷t�y[Û���Ԙn�m	�۸�q(��é.������n�0=�P�]ۣg�qzM����v!8��ݞ�v�g��Wa:;n�>���x[����8��\J]��N��<�k�.뫸W������9���������v�B񻃳V�^���69M��S���5G����U�]l[�ը8T�cr&yv�C�Y��ݶ׭�F��E��(�vg���uh���z�vz�G=8ۭ���O�@W<#�P:\^��k��aLh�v��v�ج��a����;;q�yD����VW�+�)�Ǡ��n����|�;�uu�Wg�x�۷��1y&y�V9l9�@d�6h�d���#h�����;h�]&-!:�prg�خ�I�S\s�]k^\�nF�}��Kkg3۱s�:=b�.ݥ�K�{J�97F��"q=8��WU�Oݧ�N;6�Hv����S�'�ڂsx�^��Q�=k�(�n7j�y��4����j�M�c���'��ł9��wN����p�6zʼbI��sF�Bۄ9c�J���R㞹Q�����q��ͬs�eW�Ӟ����u��K�� �y���Lyu�a�Y�편ڽp���]q�a�s���]���Hj�7cuv�]��GO8uLV8Ź�k��
��M�cc!sn��۷��k')�v<n��ܝu{��Afp� �K,j������Ӳ\������;s�;$�r#յ�Q^y�c�=�3�Ѯ^ѥi덄�3ї��Ϯ��fs����\8A�I�W�oe�A�M��W�§˛�@��n��A;���W�cU7�����䤀����;͇.T���R+� ?O����%��ߏ�qa�ܳ�ԇ� ���\��'}���%<��Yc�=�{�?�|�"�i �%b��SA%�7z�։'܇]��5�� Eټ�!�'}���}���H6S.9���Y}���� ��	$�-�����>�wvf| ����Y��S��ٻ�ì�d�O�#��,��i5��{8�p�~]���g���@MM������� ����z�ܽ�}x�I���BtZ����t�681�v���z��`@n^��}�`���$�-��I�sz��$��c�V��u�;V�ν����3� �of`>WZ�MTL�T"bI��/�j�/%�]�*[�.��m���}}*8�;�o>︮���������=�}�s��wr��� |���U�'L�ؚ�ή������{zx���Q�k�˥uަJIz/;��"P�躡�ܾFV���9�,Q�-&�+H�����	�r�$I����̩߀_��7��N6�=��rH�UJ��'��kGv^��z���H��1�������{�ȉ��8I����$��ߗ7� �L��}˧"I�]�N��U.�~u]w~I�v��&�AL���슈��}{Y���7Wn"�����9��3X#t�"ϐ]�m�ֺ��8	�V�Q��	x������;��� A>��jAAw=�XC[Y5���5U�|�|�nCO9t���)����9������y߻��Ӹ�=Ӗ4�"��n�>���g_e�7�����.=�"6�RaO�[�H|���N�
�o���Nx�up#t:,��?4���VFv�\�{�}o������zc�g��S:Q��ì��b�7�׈����7��N���؎ �l�r@vw[T�\�RT�MIX�BL+�p[����$z�H` �;�- �����N���wd�q�o�=� ��[�3���E��T����I�	��<K�4���^!,�{J��&evM4PIF�uݥ�H �;����g:LӢ���#�S3e�b����m��lM#���v]9���|�������-�H�z|ڐ@پ�` ��ݙ��m�;1����Ivg6����S-7�+���#�i��߶4W���}���I�I��l@BW�sx�SzUA�p�k2C�r�&f	�");��7<� ۼ�` �:�7N���Dp	gkQ �����/H���j��`&�%��G=��<��t�4� '���  D�N8��<���T����oB��$����������S�,u&)����oR1LaW�3����P��΀��]62s�ܱG���l�D!�ߥ�'��9nI��7�V� �����"'7���Iv)1׍Eq��#A�%\��Eӱ\���w'fr	�n�HGd�s[9O�˵?9��"*H��@l~�E��%H?�+G��G�IFwuQ&�Q�*�0oGF�͜*��DAٺ�$o�gӒ��S4S�񝑕P�D̍ݐ����vo����gwUg���N2!��ngoo��{]+�o��d�� � e Xe���{8�}ӖDC	��?Q9=s���fDg�"{�RyˢBI�h��N���w�����w�V�|��`|)�c�gsͪ�rܶ���\\R	����߉9>c|CI�����0���"p��~�����3�z�~�,������Ԑ .���S۝��O�n�m����@�:aY��)���u��.{��=�_�P���w���^�������O�ϱ�Q���qf�^���s�1�.2m*�г�d��s�2s��k=z�99����M���㝺4�=��&!I����z�{h۶:�[���	s'kF�Z�X\��!���:{y6n�᱘Xfr]�$p퀬���;07ny�ɻ����������q�|7nk�v��G7���˸M��y�,lU���X�xx8��lb�+�ӋO[<n6۷nf4��p�l�=�����'��8X�Gn�Ul�tg>ä]β�t��6O�{���-2�XHB�f�w,""'vrڐ���9�y�ѽ9�:�v�Y�ۙ� ���7'��=�8�e��0�L�F����4Yhط�����c��;�� ��w�������	�˖&�l�^����G����t$��=#��w�'@(΋�^Ḫ首+$�	i�-����׼7�����I��d?�Hw=�b��َ�r�_�c	b�^�Z@�8�|s�D�10M!E'mQ���Wn�ϰ��Fo{{,sq�ekD	gkt@��o	�N)���w�LH���8�7��X�jg[��ڣ����܁t=��g�۱����X��Ϧ�I������K��jA f�t V�uQ!�]��ȋ�ʋ���"JS+����E�Ka2���Ҿ��w�'	[n��ՒH��v�)��f���K���E�t_T�17Q�%�z����B�o�/����u��ۃo������I��&I�1u�=��{���fTW�I'�ݙ� ��!�w���ݑ^�R���@�0�O�#8H�� v+�/�c�(��Ơ>gsiQ�|�;��a*�TL�4��Wَ�g4�J���S� �=�А V�vf@���k�y=<;�z��Kʱu���Y ����SQ�=�����J�sلؐ漽���;s�d�ܿ��^�u݄��J;��/�
ӂg�W �BF�ɱ�6�v�	�*��ݶzqs9�j�t��-�ղ8O%�y�
��y7�k=�@L%��UH�#��%y�bS����L.�2 8��}�}�W�i4S�@��D��l ��َ�'.:���ЀAY���`��� U����ϭtU\��oe���aa!	0���f��[�������0�zA�ڭ�&U�wD&�wJ%���g�+n�y�����ۯ��y?_/��%j�6z�@K9�.y�U�<��P'{�(����I�ou�6�Q�n�%�O2�BN�(�1��z�]�L�{�>Iy/f�`  �ܷvo]���Ο��t�;��Iw�w`$;W�0��$�WL����� Avg4�lZ�9�׻3{�&���| �{��D0��z��*�_�S�ڰ��'� ���	��b6xKnq�L�j �VT�ѭs��r����l~�ݕ�����r7=ێ0�ʸ���ޘ'9��uQ�W�h���۲m$���D4��D�ʘ&�����(�:>	/}�U��v�]�s٭��N�[� �7�T@��i����uE߬����r��f���TL�/��� �;_΀>��V��7\z���$'�)�� ]�����[�u051QJ1tu�\�{�\'�u�.'gi�5�	
�s\� 
��ي�t�}��y��5�Tgu�h�WAiI�>߳�/�s�����2�.�����+�/�=�Ms\��!���(°�&��\�b�V��� �}�����I��jf`�¼v4� �osł�~*{j��r˨�0�;q�.�:ܐ �}ݙWĿ+ے|�R�ٺ?��l�,�/nz�d��rP�ssX^7#�v�.�s@s��5�������f)ULM�7��m �N�'�]���	6}��fwn�]穴�+"&���~HMGw��g�>T�)cSe9�V����� �A�w]�Iy(���Z0�Lh[}r� ts�D�ʘ&����A���0Wn�� D;]���Uït��� ���7�� +}ݙ��E�S3TT�(�[D��c��r�%��v�@A{��� @}[�ّ�'�)̓�:�{��$��\y v�S`+Ŧ: ��*)@��u�b�I����If�L縌�؍�~���>����H�D�:l+�.
�C����$�V����,�9Q`�w,�s�K��zQ�J�f�>�	� ֳ����rA���Rxn��=å�f�	AJG�����6V< �9�[[ke����x|O\�+*m9������,����n.b�Gq�9���J��=�����K���-��ϬZāx+�s�vj^��@.L��ŝ�������5�O�-���n�n�s�4��yݽ��u8-�Qy�n9�m�G/�<Y�v�b�5!�ܼ��k�p�1�9�y�VN�8�v=��uPN����b�7kp5��v/;7&����Ռb����K���E??6����AIeq�^�Ȁ+���`$�)�v�c�!�"H���y\��t��޻���*�"e�M9t��Iuon;��7��� |��o�=ΜA&��8*����`�8IaC��fonb�H�umA�1�̙K�lA>�߀W�{2#�{�6�z(�	~���l'�|���ת�K ;�n5 �S������rU�9 }~����#��l���+fa/�M���m4��UNeTF}Y�٘� ���M� "�z�_B��Wo�e7���~|[�������Ɲ�U�U��8)�4�;��e�m�qr�p��������=���oq� 뚰^٨�qG]�ۘ�z����'��h���R%"�- ����9	%��o��fu����TA�P����t
k�ld̒��w�����5q~�>��W�ʽ�;�"of��4%�����R�N��^�غˢ�5� 	�vကE��7�@�I��Q�S��$���1D�������;ަ� ��:�L>��r�=vy��x�=���q�w�M��"�"J�RT陝ۅ�*׷��׮g�>�uo��>�z�� +�{2��O�ujK��$����'��F�K ����n+^
D���ޫ�
;�G[���
���0�>.�i��
��������Ԟ;�Q�����Ä��&f��i�u���1k��gtlǊ.�l�k#��6L�߿���35EMB��'`�ھ@$�w�W
������2=��_nӈ��E߽M�x�q2QB��l���ŀ~jz��g��� �@]�ۆ�]��v��G��md�gE�ט�d��E��ePBB]�9� ;��N�$�.j��g8G�� ���MWS��8��v���q��w��{U�ݓ���@��]ç����:��6����rnE�D�Kݸ�2�ތ��bwPUvj�v�{ۻ��<�9��C�<_��C�}��2�ҧ�W���������6ʳ��v���Bl�y@��-ͥ[���d��Cd�匝<X�y��{w�:�ZO�ȁz=��bɼ�k9�B,b��wȇ��>�>7���T}m��ݴ��2���az�{��n*��F{����ޫ�ܩx��ܼj��`��Ell������Y�F�C��Z�D2��H�3Қ�OC���K��)���
w�4��O՚�E��ޙ�P!�λ�b��\�0�{��fɞuu�n�M�$Խ��7ý�]������wv�6a>�Dz�M����+v�oN�T�4��TKW�{m��ح�Pt�Ǽxs[������3��ֿnFV�f�kF{^�g6caM���� �V��i��k�����(#�s���"�׌1;Z�Y܊��A �{j7N;���̽A��כU��9�x�ֳ��;	}wEMw��m����o����z�w'��<
g$˶=���ș���mn�/)]x�[�҅:��^R��� ���k��Ӌ�Ʌܔ���D��`�Ba�q�v\�1x�s�o3�p��]��J+:�%`��zH�
�~wO����x��{y��/~��G=�U��z�����'�q���*�#��J/ɖf����Fm���6�kQ9��ʫ�Kޯ���-��񇴪�#1�X����
�-�l��!\sDU��b��35�W"��F(#m�b�ٖ[faV+Z�0�2Ҍ3pJV����[�b����q�[[*�h�QVV�1b���8�	[[e�q����U����UEfd�ض�UJ�kQ�na�r����,a��\�ĵVa�1�RQQEEQ4�f��q@jTG*��dr���+�UAQU(�J6���XTb�S,�#�����&aFe��u�CUJ*��X��PA���Qe�Ɣ�\LLQƘ�J(���[,DPr��N��s���S����۞�V�dG�UEF��n[#1,\�r�PDĬ\d�R��bTQGMĢ:�R�E�QK[�e-�U�UZ���"2����V�ĭ*�[2��r�#��j�¬UET��+iDT���c��1�� ��F ���E-�������"媉�UX1o��8�����M� V��f|�L@��T�ĕ%9��ʹoۇu�R��wm6�H'��4AwK&z��O=��eU��
p8����U�J��$�V̕Q�X&//���ު$⻥�����o��o��Ѓ����cŭ��>#O�^��\�]c�i�HKv�c�����ߧ��r��@����I{��+��O�tȓ��׏�����wuD����B���8I��$�/�}�f���#�~��$���"�]�� �'2�7]N��}��7츤Ra�����Fx��e� ��̵U�j��3Ē�;����.A=�p��I��(!�w��^�a��8��9�� ���D�A 7�ՐE<[�)��Ყ��D���zogL,�d�#1]�����	t�:j��]tm�F�k��ٰ,�P�;��J�b��߄s�3���@:�g3��E��w�� H!��5ˆ�lc0/Ʈ�6�z��A]��Io7��M�Ȍ��|+r|���9��S1�nx9M��kr�����nǞ�vV�.��* �0ck��'�1��N��0����w�H9>�8��z����0�{��~D�Ki�^�*�.�x�с��S2�joĒO�lϤ���@�c�f��gl���}D�~,��E�%�V��翀 7���/*3(E��f���@$�Vl� ��aU{���=���TP�@����S��6$�l��k�A7]�(�������\�C���$�W9$uF�&�C�\(2b���	�wH�(�r��v�2d�9S>�[��A!�oPɆ�u�ģD\ 9��g��E�:��'��]T��׋��{%�cݕ���\$B���c��5�ǯ@^��>�ƃ��L������^��]��r�k���`;/dRb�N����a��8P�ƭ��ق����--���.���nl��P�b쉪ָnŷ���Ш�m�<퍒6V���:�p��<K�tg��m�H��y�`wc<u��;�-���r��a$;�O�b�jM���:��i�S���� �L�8Ϛ'��`��ۚ�F΍n�Yc�xѸ���۳��6�n��F������ů�h���1 ��_�ws����I������u=;5:�e�;��7{��� ��͠	6����7dt�F�F�$���W��{z�Ăi���O����L��m�&�`<�)�MK�ޚ�����ݵ*t�p�H-�l�$���������I��A��yq#N䈨�s@�=��D�|ﻫ�Wt��t�Dr��|EΎ�"�g*���lP��i��B&�پ�$Wl�%��LD潽꺖"{����]���>'�wK�e혼��6:�J�S"�l@:�wD�2Ԝ�p�r��Nݘ������.�M~�߁��1qB͜��Iy��(�J�z{b�,�eUE]��
%�oU/p#81���$����3�"�,�{XY�+;�\}����@���<���~���1��oϲ��
�Z\�4���w�޾z����Ϣ��O}���wO����A�B������+���Q���)������*�>$�,H$�qxt֥ZA���I+z\��ݺn@0�K-OX����e���]MB��$�}7�Ob��r��H���~=���,���+�� �{�*�WAy"s�ox�uY�D�I[����y�TN�r.Ȫ"&+I�	@P�*琎'�LN�Gj�qV���}��v�;V	��fioz�8C���P������	 ��rH$���
ehM%b���;9�T	���s�@�<�JL(��qd��]xQ"q���6n�)���,ّ ��}�TS6guEʓ����4��)V`���N������<��$���*��4���i���	1����Eo}"��<W�����uM��ׂAa�C�蛉Ԝ*{C�J���f���5�^�}��=$J��Ô)=*�`(��	*�\�I����`y C�͠ě{����b4x�$œ��<Hv����u�4A�ooT��S��7P7].I�e�q`6Z`2$���� }�`�$:��<T�E�� �}s*� ���ު���g˫�#~���&��- �6�ƻ[k#6�]f�n����.�@����Ğt�:����u���I��-�|An�LwoM�*������nO[� ������?.��i�B��������e�K�A���z�����1JF�c�jO#R�
!�\(2�����{�� ͉��Ή�Bv���H��ʢI[��D^�&P����˓����o�8ɔ�'s:�$�۽TH$�9d$����>�gN���j�{oU�����g|��_V��9|ӵ�>�+p�{���䄽��~o���y�l�U�⣹�>�ewLZ�&;:�=pJʄ����6��*�O��˓*iM���f�9Q>|��'��UI �9r1�i0�/��UF?>�\���q������=�J��\�N��p���I�1��$�nK��4���L �}��{�+ݏzk�|7�Ȓ/��D�v
�1 �_T� x���O�����pY	2��n�<li�4�]����;Ϻ�	yː}��7W/{�{N�t���zvن`�,�Pu^�w�^'�g9s�	v����˃�!W9�|Nl�P�N�\����H4P����p��s�u�O���2$	󞾠s|%�=��ڍ� �E!SHJ�����" ���#�+`�U�u����A�\�Is��@��iսG�A�=R4�K�s�'��'�_s�Դ�ekI:�"�-��
�5*�gx	��	yF����e-��sw��މo��EF��S;ݳE����@;���u�]���d�䰞���\�]���6�֬�c<�Ik���n���n��\a�ֱ���nrۓ��T�nV-�X޺�����N�<�Z��������]��m6��kG6m-v�e�k��4J�����l�M������n�#�^3]��J-�x��qf<�I����g���x��I�F���N3;�;ջg��h�	�{�x�S�a�9s�ݺ�5�Åb >�%oAD7�Q��neP���� �����7�;��7�*372��>�^��3&O�i�6�`�`�wUƏV��9��);٢H�rĒ	s��^#G^����bη�|	�n䊘�APF��W
��Zp�"�-�P���{E�w����o��O�ĝ��!�&`�t�t��+�;p H=}.I!�v�{�zP�۶0�٘��,r5$�I�4.��2�~�`˳kq&B��1dH$�+���ު���A�m�6%����3	�N��ݒ�W)͵�f��7*lg]@���ۤ��ߠ~~�!6JF��5�nH%�^ТGt�M c&j=[#�0\^9��7}T	.	]0Q��)6���� ����o��[�����G��&�k�s�x{���P�!bW���0@��|��f���GEÔb�����~Sj���J;S��p�����Ϊ$F�oUxD^���>��g���=3}amaX�)�$�*��A'�������0�Q�^�ۿY>��ʯ�[�D��p���I��A��s�4��m$F�w�u��y{��>'��Q>=�]]^�y�&œ�W����!�L�Pu��0�r�3ON�B�켩�E�oUx�H=�\�ѵk�;���s�0`��2��T ��2]����s{3S���X��8����o�Mr�\
U�]D�����}��@�2o�����<��$��ު��J���`s>�: �Xfs��B���mOewUw9rA)؋ZL�pˊ��=�w8���o_��'� �׸�0U�8��b��Þ�u�w�h̋�S�8I��w���&ؽ=2�����94L��bH	��z��=Y��t�.�r�n��y[�^$;��О�M�+	5�䂮�ܑ����������gd� �9�$����C�s�H���)�����EF�(*b�@M���r$�9�Tfs3�'t�5��@�w�^���~{=��
::O�ʝ�P�Op�p�!;��ӹF� S즒��q��p�<iյ�@��t���eD2A�z��U�r�	�oM�b��^v�ܾ��$�|�����>,��A��Gps�t�M�qKշqs��'ē��2$\�����l��s��7ޠg��g-�\������2�΀�����$�o\��淪��T�DM�m�?��wǏM��@�����@.v�h�GuoU�zbR���݋��_QWL���-ۋ������]�<r���c4jX%{5��c�Ӣ'���j�	
�e��ӵ��.k�aC-D8���}5�;kzhĹ�;��Ý"r�"̉ �Ho��]��T��vى��8&y20�%�A�m�F���;Tj�N:ۜ�T�n:T�Z;h�������~�I8,��1���rA*s���N�oUx��h.��]���'�)��O����54!
��Y����hM����W�����^=ս4Bv���b�#*�x��Zj7�j!
�ڜ�>9��"�&v��n�"��+�IN�P�w�zh��>"pA��@	�����}���b��'���ʢ	�9��U�=/z�؆)�\�����O`?n Bi��M����B� �t������Q$���$�9�����ށ$ I?���$�Ē$��H@�Y!!I�d��	'�$ I?���!!I�d��	'���$��H@��	!I��IN�$ I,���$�I	O�H@��$�	'��$ I?�	!I�@�$��$$ I9$$ I?�b��L��h�D���� � ���fO� �H_,  @P*� �P        �@

 PP             � 9UF%l4UJ��*T��P��USA���D�QB��Z�TR�F����J�(�*�;7l�eQ�*TT��                                     �  �      ����1�a�9i鵚n`4�c� n��0 D�ﻡM����pu�`��݀�� 	���ngt���=5��IE��|   ��|�t�M��L� �:������B�5\�Z�68��N vk���Zf����<�'L�{F�2�l�|   �       � |ꏪ�s�(9'`}���X�S��x  ѐ��nj<f��Vmˊ���S��� ϠG���)K�4$��v*�ٵ��   :
^` is�t�4��J^�� ��,�����4�'��)�Ҕ�/{�� ҄�w�� A�)V0wy�4���Iy�:
|A�C+,QɥP�*�HZkm
��   �        z�V`�}��@>L�^Y@qHT�ʹ�P��]8 >��>���b�{�M^f��{<��M� ��{�z�O�|�e @�5��  =��0:} Ǹ 5C��zǡ��a��s��7�u��� .��ɮ�)��Z@7,�N{��-�Q�           ���WJ���=h��@ � wQC�g�`}���*����
{� �
�m=�t�uO^�KF� ��  ���(���K� �ӛ\������[��GZr��S. e �{��k�ҫ�ɪS���5@��hh��d�  �        �Ñ�uT���F�ZA���� ���t�C�5�i��Z"����{� �z�3{V�s`{ȅEd��  9����x�t�� <�8����\Z@��y�T��w���Ǽ�\�yt�:��x��M_ � �M'� �)�4�)*Pd ѡ�������L�  ��UR�@ ��~�	�*Pb I��&�)����������_x����F����ͷ���x��$�	��XB�R�HH�	!I�B��@�$����x{����;��.?��2��d�F��`K	W{USIy)~�[���~+���u��7sS7@嗞ݵ��ִ�c�x���Q��kZ� )yj�iI���Gt�������$e�F���Nƻqtwf���FB:A��:λ8�ǵ��d�`u���x�[�-N�!��U\��c5��&��6^��b�F{ya`�@wc=�yp�z�V\����'��l�= �=�A-=����Q+0���B��_-HW��+��=�r�Y�m��p�VC�E�����8ƒ�=x ʛ�f�m��bh|#)�3����`�]�����2�ʉgWJu�Bf�H;p�H����};zYޛ��I���A���7��C����J�
˸Gb��m�Wt
x/.Y�K䪬�JB�y��˭����.�?�T�j#k�8*v�m=�İ횶� z����Gt�{n��$�N81&����k��OwW'gt��d,�PC�Z`J`8N������/���i�y�1r�!F�B@�P��{%��c�k�X��+�}�VE��xp���{���rf�x���B�&�s�gXqM:�$>c/2�CU}׾Z[�ؖ>睏���m�5nW�<x��}7{bk��w��`E��R�*s�	�u�:;�{�jM�7�0��0���n��$ �F��6"q{3�����=
����"��lM�eow��}�x����b����:�\Y�n$q�|x(���bWx����fH�xv�;:��p�0W�rh�h�WkK����l�X�����k�S0��T<):�:G��Y��������A��,Ӽ_f��b)��:%�7��C���0��KO Ϳ^�Y��xr�{�)�jո&�.���1O���fwg�V���;rّ2M�D�<��f��Z#��0���U9�x_X�k
�3�(���}:��.�\�U�^���y���#	��
h��1@������.�H��&>�.�rmsusڑ%h�ز�tC{���P��0/�ټ��ۜ���r!���H����-s���&�����{f��<}ۭ7���Oh	ЏW�3�)������+�J�[������Y��5��Y6��2�o7q4� �C�b�n��8Ɋ�[��-�W�ǹ�M��!����w����]{���a���s������mogy����|w8s4
��#�ν��1h�ˍD�,�LZ�jN��M9.��}�/9o9v�3�>5��7'ܲn�V ����5�U���p�Pf��۠h!�o�����"-���|�͑�z�!oB1���e;��85cё#.���PXX����
^9�,�ޛܖ\ь�:����*�3n-�������ˋz*]�N�K������c�פl}�\K`��-�"wS��[n���0X8:�r6���9�#��v(J�w�6�C:�
���,�6���xs�F������We�=*�����tV��6�_<�=�!�+t:�r�fEܓ 7�P5td��=�����.�oj���3A=9nYTBv��\�P���)�\�Y�"䥜��-ssdŝN�e�V�
�n�igqiڮ�W|ؕ�x�V3�uq�F~��Z�p��
�sC���� Fɯy����т@��Y@q�)[&������ ێm�a�.pX�"����wo�e¬d؎�n�"x�r�8`H&�0�saN�vb�g R�꩘����2=x�C7L �N]�h*X��Q�g2��|7t�۽�>�l�*6��%5<*\��A�Ҕ�eZ,\�udx�<��:�<����$wE���NT���H�/r��i8�]�7����C�u�p���0���\O��t���v�0;&��vS�Ϸ;P���U�k�Z��f�LR�0�t�;��뙽��M�Ç����p�o:y��8[�=�����^];�lͧ��O��8\X��c�F���`b�;�=L�q�B��m"8�5ۨv�9���ð{�[���v��)���N&hģ7��:�EU|*��z�si�����s{&[WS��zt-q'ٱ>ȸ�{I4aP���gm��nѻb��CE�1l���.���ty8�5�L֯%�Mȍ&�4��ݖ�f�閞�5�P[�5�T%C�oÐw{��]�x��kO��N^/	X���ݫ���*_
X��˰�Y�u�q$����&��i�'�����;�wH�m�w�,ɵf]���"��� .h�x�jΥ�v똍��B#Cq��Z7:]�hg�*�/ot3�^+����T;���g׾���T�{'!|���Z[`���k�m=��@�dIjᲩ�d������/>������՝n]�+/���+ !�T�CS��Y|f��`�[��%�.G��r��$�^
�U7��2���U�;�%fۮvL��xv�bA���d ��8��%:�sR5�"tŰ��ƌlq$N�����GN�c��QݜY2�& U�
w:���w=�Բ����6,�A�3Х����{,���f�HS���K'Y6=ٻ���e�zv�N:Ps��X�V�f���"�o �!Tf�zF:u���Ջ;���UL]p�ov�T�����t%Q�G�k�jPή���^��l�Bj�L��s`���/7þv��q�s٭a�:�79�e�CѶ�i�{:���ׇ"�^vp����Ta|f�ni�=!.����٫�c[,���ҥFhC:!�J��gm���G>AV�Tm��<��[�M��_�&"B�Ys�p��r�D�׎���ӓ�Ƀ�g)3��3�⹞�]���&���=�;�Z©nP�^�`ZEѓnI��ˬȱ�+�C��|�p��q|	�X؅�cD�*rӽpm�Ӹj0��w�7�BTl���wZ@UYd�5l�q��.,/B�WR�cs��Zq�Z�ӵΧt}g�^�^�_,���pBժ�ә���y_^䖗X�ɽ݇ ���{	۽�߯v��<��Th���Vެ���sK���|����n�_+��V���	�BݸT �����9v���꽳F�)ʣtb{8��{2f�7�R]' :On�T��`3tl�.䑘���&Y���C��׮okѣ��LO:kf
�=��s��+���RvX 1�4i1�9<�ΓB@�an�)G���m�2V� �Ӧס��rُ+[b�ej�#X�z����2V��x�����=�В�T}��
otuڦ����N�¢;�:2;rf��'�x��(�~p�&�Ѻ�I�6U�����;�d�3q�Ѧ�C���ϰ@8#K7RU���ڒ�jgZ��\H�����Ǔ���]O,�91�Ռq;m��(ܛ�j	��]Y�/ �mB��"���SsNN�q17�e"�������ZnHq��	
D$�O��G gF�݃��n��8���Iu�a\P�ݒ b���V��M��,� �z���Î�+.YWC�2��n�L�s\���T��l�!̛����NQ�K3w	S8�w��C�`�Ag"�Ϸ�w��l�|nɀ�5�՝�#��~��N������J.t��!�$�%_|�<�goh	l�ɦ�9+pX��ËhZ�DC�Ӭ��+�s�=�Z]p�:4,���M^�fsz��Xj�J��f\'����<�Ҋw ��x��Q��N�r�O_�)ǰ��Q��	�Y�;t,��c�twB�&�XJ�N����i<D�u�OoÝ!��d�2Dk]��cS-VX��i�3�YO&�>�8������{��g%q:͹�r[6G5)��6����sG���掼2���!$�y�y��ε��E���Ș�i1�ܧ�(�P�v��]�Z���-\�؃��ub��۝j��M�����`�仰�{9^ã���7�ˤ0B�0	X!�*�z�G�j���gdA$&�s�-2���k�P3fv]YX��&��բ��:��C�N�w��a.�Q�*h����B���,�`Z&�d���܊L�FLSg"	�U�i�P�H�4�Z1Y����Lz��xJ���ץs6�i6l�2L�ܱK�5`�Һ�;Ce��5���c�6��;`ĸn�4ahN�>��3��3<�y���狼��gA<=��!v7��{/�gd�e��ޏ���& �`�2��m���þG�M��E;J�8~��#</�,�%����!�9��UT-�p K���٫;f����]�S.��*�Xr�b'��m��f�ğ-p=zk�	��^1�W���i�wwL��7�k��9d�� [!�n��"�:�uA�^�6��	h��%��y6:�lF�x�#��oàᢾ������q8���ѫE}��ub�\��{����lh���;;.�u�+7�E�}6.��lv ��h�=Q:yuHD�t����ם6aw;:�e�2�
��=y���Λ�Tr\Ӈr�'C/j�&n@/d#����Cq�[��uw]|�V98S^���n���V�(�ѽV��K�:��f��UT����M�ܞr5Cݫp&Y�����5r����c'�����mR䜛�8J�%��V��=��6��2L�Y���Du��A�J�� ���O�lЅ�:L/;Yy�0(��j�za=@BȊ�f�Fcq�d�����h�T=׮�1���|�p�ڥ�[k��	4!K$�������;����w�b�pLl��{�ع�+������pݕ���X���L�o�fi���P4<(��o�m�<�a�o���Gz�3`ou�C�c3L��Wr��u1U���X7uNո�`�*{��0N$�;D���ڴ��R�S�xx��ϛC6�9�aq8�̙wfvh:�}�4�S1n@��rk�n��m
]-���qx�Nl��F�N�Sn��%���r��{7�q�R�5MV�O��� :�Z�`�!��Ca��ΫI���w˶u��k}@�;�ۼ���i398Y8��Ȧp��Ğ+ۍ���9	8u�.yw8
��XX	��o5HW��;�R ������&��t���I0.�]��n#���u�/9s���ۯ
W8"��^�!��c77��8�;97�u8��h�����:�ԑVh(���ƙ����iR�-er�{d*�-��t�a��f�^�ܶœ'Y�O;z��������Hmq��ηN�#�Y�����]���S8\�f��c��p<y�v�i�r�B�l�����b��6�3J+7!q���u�~�\]8n )}��Xd2��v[��a8k��}5����B4����p���}J@�u@�u�*d������/gm-�3u�Y&��A,�y���+�p�9O]U.��Zr����"���@�v��s�n,i��<P Hof��s`!�8��X��{G4�ZB��k;��^"_�Õqw_n�����܂Xx��e녓�d僡�`�tP7MaFa�9�3r=#r�4t/�:H���P���0n>�᝗|6%�k+�o>C_o�dn�ܗ۲�؊�M��#\um�A7�듣��yT�ND�5E���Q�WC�������5a]K�L���2)z�p��� �n�6h��ꁣ4�;r��E���)�00噲F�g9$���w� ۛ�2�O4�W�	C�4lC�J˸r�0\-칬��m߄]�A�o7D��ww�Vy,�N���,�F\�9ׁ'�қy��Jɮ��eq�����Ge��Q���f���8%���J+�N���p����zc�Y�d�͚x;��MOK�G{LY^K9?�Q�m����6/�

��0d�1&b���(�j"��v-�f�Tn�a�.����L9[�9m��-�w��בױ�xW
�ǵs���[��IЬ媦�]�F�K��תz�,�[����HO	���A��8�r����3����(aﺼ"����*��z0�,6����	���7<�0P-C
��f�1����pBY��_�ʺr�a�.md'l���ޙ,I�V�[{�����D��p��ۼ�t`M�5"�,�=�<5�w\��Հ��g)��"9�y5:F��3Q8 �w���HM����ʎM���{S�ΰ�(cf$�G'l����E��s���з���7��'ø֮+4M�I��[D�HQbj�3����QVFZu4OJ[��u���ƾ�ӹ˯`��xe���٧��MX�ږhw-F���ܧ�E��w!M���.�U�ډ��(�|�v>����&��E�lҍ"�x7��Ȧv��9Թf���	��څ֮�I�N�hJ����{�r+�����Ǧ:ro^�_a!8��:�·P�ŗ�X�����|��Y݌`�B%9'���r�|;�`/�t`�n�r�	�xp[7;y��Χ��"�}����f�˥�z��!��6��p�9�J��n�6�Ѻuk*��Nc6�Ǉ��>�����@�@3�w�tl��� ��-��F����N[{`�v�ׄ�S7z3�� :q+&��f��O겡�JZ����a��P��	9���  x	 ��
��HT�AHA`�H,�B
d!T ,��Y	 E$ YAd����X��+	,�d!"�B� �"��B��
��I�PY ���� �$PHT�$a�� $�, ��J�V@R
�*�d )!��, Y�I�$�IT�@) �! P)	*IP�E�@@	� T� 
 (@P�,�E�	P!J���H@ � ��HE�"���B�B,��T!%I$+��XRRH��	 P!HE�H�HAB �`ABHB���$RI"����! ��� IN���?~�q���x������vK�<.fr~]F�cC����k�'<�opg����,op���V̷O�@h&6�xvy&��gn��{���o��/��$�ӆ#ݥ�=R��:����os8���N����d��v��z��[�ꭠ7d8�r����1\s���D^�'�xl7ޛvϸ���r[��O{�8w�o/(O!tk�<�z�}|#o����;���������}�S�*>S �Y���$��ߑ���"�sx�m�<x�^�t~^�+״H#�F�f���]��2q�=�xu	ܣϘ��04��/NL�s�Cz�u��:�l���~�,G��k�2o���{=�˼��Nݰ�?n��sF��' E�8�Hנ��>j���jP{�c�[Hm�����zN�+&{7����lnE�@7�gq����-��\�.��Kb������<�j������y{��݄��lah��ɏf^�j� *FMQ�JS�3���;]~��+�˜6N�
���Q�)c{������׾0;t��ۓ�r��;;��E�X�|Xѡ���9�{�8��=n;��{$i5��4vm<Z<��fk�x�������Ut��������v]��`�F�I�n�;N��8c���;�^����d>�<�5{�:�˧U�eQ�d�O�@��o7]�n�%S�T� �,���������7}�p^��6�17e���$��2<��a�y��X�[��� '^���4̅��� =>�߹��﬍��t��u����0�{/�+�*�BO�N'��p�zX\��X�p�+u�������BÒ� �'Y���MX���|��}�q��	[�2��ٵP��C�u7��w�g)�
z#םio��r���۹�k�_�h�F��"xw�fy��x��>�X��~�qo�'|���}��g8����6ٶoiВ�'Yr�[��,weB���3�؇��M;��A<���ub1�|��fVX��o��s��S5@�tvkֱ�I>i
���Z���s������:�q;���v!�܈����+F�����Pm!YUex��7���;ӥ*@3�#[�������,�69z>�0<��Ϙ��# ]��З�b�����tmiR2��˪�(��>��^��m����Ϭ�1��yL#y���.����9�|�{6<(�X15�bm��H�k�6�,mŨ�)�z|�2�P�n{:�t�Ƚ��K�59q��h�ͣX�kGZ�(����_��Fg����p��;��&��{]/�m�^i77{p>��Z�@��=Fz�@�G��M ��~�R\��5v� �)��@)�Xc�~���$>�w_ze$���n�������=��m䧎$� �j���.��7��Ű���c���(�S=��m�f�����g��U�6f<�vr�J[��G��<|��,��dj�n�����ny�6l d��R
�<^zIcbZ���R{p�ś��=��:K)��B=�R��B�ɖ���S��O��I���s�o�:J;�o��un�Έ�`&�:��&ݦ���Gs���ѵ��X�w��b`Z�K�/����4<�"J�1��~%��y���7W���ɜ���+��ݮ�;�T��t���[�
H}�ܙN���c��|����xc1kO�w��<�c���jSظ�8u�g+Oe^'�E�^��U=r���u
ںL�U7Q:q�+�F�a�u����F���p�/���oY�=�f�cyC��B�5��3�|X����0&�9�x3鹴��*��Yw��l�-�.+�f� m^�n�7��N�pJ*�mZ��l�޴׉c��֜��vP�B�>�K��ظ�!�Dxa��`z]:$��I�]ܚ��_������f��o
�=<��y纯�t�i�6=�|��`*�+�z|2u���UR�g���kWYUr,}=XWx4�'e憽ї��{����-�7;<}��(:����b>|���5���i$���zC0��ИG�Jˋ~/Vx����TwA�nMO�Qk��c:����sݛ]�~+�.�dܺ<���L��|���C��-X��g6y-����L�,�|j#���p��۲l~�/{���z`�G�{�p%W{l���|�z`�wؗc�}�-�2�{�e�����/kۧ�V<���\9@�vB�lћ��mw��R���OS红������b_�ش��v����Ȅ\�^{&��܀��t��̺��x�ît/�6?.����.���b�E��w]踑�i|�[��UH}ͬ>wi�ϓ��x_q?s�����_���/{ų���m{���w�ܽmh�z�6=m-�q|uM�C���\_A��P�P�z��1��:%��I�Fr��|	S��8��S��C���T��9���v����H��������k���Nkp�z��мFu�3{+�_\������'g2}�Ϻh���\_F���ꠙj�D�_[���{&�9zb�r!��9�����q�Y�=��t�Ը����C-���@�יZΠ��X��mXw���v{B��4�kR��L������ɢ��C��(�i����n���Ȧ\���Ae�l�H�={7�q \ĞL��C�Ap�	 �j�E� �o�T�9�xD����=<Y�ϼ����H�H������9�\���.�:
�ҧ:O3:��[�O�ݙ^�ݒ��kr�c��h����y���%�<�c�X~w{Dr\��E�Y^{��S��x��.�u?ow��f�Nk�;�&��vY�����g���$U9#9T;�F?{p�{ �:Ӝ.�����y#�����U��`�cf�[4	qZe�+a������q���S�LL-�V��1ص�{�~Ow�F��ї�>�v^��snD;�a��kn�k��W�8�|��{�>�[��9ֽ�p&N�wg�>8�W_W�3u�|R^�K<�7_�ce������l?��'���{'��W�~��0�'�%ϱ�������#~��=�j�������������|�N� �N^p�}oܹxa����Y��H.�o���kc�,���r�;�0�}�9��[խ�;������z����vR3׽�V���1iI�[)%���k����giѕ��bC���t뻞�M�*Q��xΆ\�c�����\�7#PP�xN��4[��v�.+$6�O��F�i�|�p�|&zo��'޵�Y�QCB���!ű#xW��f�IŎ���ŴF���$��(ҁy�\Xtl���X}3&�'�=^�xS�cש�Z۰����97.�]�8	��ξ�۽oCTj��]p�^�ѫ�e|�>�-��p�N��_�_��D��Tk'1敹�[d���Y�zag5�!X�9�׾�*c�˹pfm�6�����+ �Sn��=�������!�i�Xɡ���q(h���@ídB{�轝���Q�^����w���6�V5�m᭸��u,fLp(���9���٬ǳ�����9O_�Ξ��_\���<�+��6��H����0y�7A���Ԫ�f#�¬�h���hI�;Z:��D�]���_Uނ%����:�\���/+��9�+�6������i���\d�_�ٞ�GA��n�S�+-kw����D�=iVe-'��\(����GC3f�Gc� ���+,�w9�0�o������8�������sO��6�9�b}~W��q�k4M8����B���b��'z��~��ĩ�����<o��y��;|���p����ݖ�)�� �w]�����~�$o}ፁ/�`�l��C�5��K���U����̿f��t�J��foj2Q`c�"{7��~�2��=���l^��k`�Aq5�]]�z�U����T(��4n��Ӧ�Y�6GE��� ��گn&Љ��'� �LO�h�+�&�/�$�ǯ�B���f�^��|��мyٲR���#���/A,�z�x���7Zݯ�p�`�r^�=�
>�9���O���l�_�|<��$�^��Ȅ}nw�j��ɞ�x�/��^`��h}�����=�T�� xW*ϙ�^x=�y�mo�THS�[q���rl�eԘ�ǆ�����i#|v���d|��R�j�;=ξ����ܾ�
�6={@���~�Lbp���8���% ��;��wI�5�pKr1�C�����օ�u�p��6�By���]�yrV���ѭz�"��;^z!z��E�}����]��Ԟ�����ڡMn\1�p�ܠ�f�jꍍI�!��r<��f��W�~Yֻ3�܋��͍���$��#��w�D�o���	��G��M��n�bI�X��(<��z|\�gG��+�{�e�C^����A��`���{̷���#��ȓ!��p+U��İ3QZ�ĳ��LG�
{/M�ȏ˯C��}��p�G��5�>a\~{OJ�:!��Q�.ݙ�X�xzn��wm�� ���MDۛ$�x����k<{�oxM�������ƛ��N2�Ӝq�~AY��Ԏ��ё���8<$G+{Y`>��j�.��X�\��<��#0,�'\�OF=��y�$4���Y%���9W�$���5�����a�J馩NcǮ�N�,������ �Fsn`�߻g��8���b�:d�K}��|�e��{Ɨ׷�6�A������5�[o�G��x]�pmLy1��;��\�p�{:��5�XA�`�p�����Q��7$�"�w��^�S���;�]�?���ޤs�2��X�.>� �.�ag�>硳z���"w�6���m�+���l�<<�1��G�l����ޅ^�YY�]tg/=WJ������rz��@�=��۵�'"}7�l����w�wx����¦f�7*��c$g �Qho]w�I"v�p��^�����7�g����9�x�c}�Ҿ�����E���l�[Z���z���ϰ_�����'ýN�;Sf"�
v�����k��z{���~B�������ǣ����O@qw�v�]l]�3s�˚ѕ�!�s`�$���ot$�<Ǉ��Y��t�/���{��˪CU�����f�xQ8�zv��/�A�i�xz��*u��c�/�m�����W�lj�n�;S�Dl-^=r�b�/{sp�G��{�R�z�-�Yc���D	���5ޝ��No?M]�E0��;��/A�8�|!8�t�%�խ��3���ܙ��y������AS��"�?T l�(�F�qq�T+Eӵ�%���wus�����m\���߶�ꐭv�dZ1W������;���q��S��ܷ����g���<��ԥg��4dT�T��G���ݽ���5�+t֎�{�^������r"��zo�o<*g7���oZ�^�f���*���>&�5o1.��
X�}_.�L�"���W��=e���Jr�(,�w�-���$�sdh0�õKjA��«�Q���E��ZC[ٸ�J��13d�����#����k^���}�|�����:����-�o;�c4^�P稝�P֖.4n[�8��&��_p�dO��W��N+D��W����T�z�_�vu��W���y�;��N�w�Xv��duՔ����u��k<����/��P��j�������`�{��rW��g�mKk��z�	�.!�ا��Κ�9ץ>u��mw�������O:Q;�옻-���~�ms3,<S[�t��F��()��^��u�"U{xzm j�徛%�v����S����������p��\���ۍ�9��n��s�gB|̭�i�'�kO1@ۙ�Z��ٶ�M265���<X� ��˧�>'e��o�We��/�ŵ�;o�1Vff�,#}yXH� �H��{a�UcQ�^��x��L��{�`{�랴x��#f�|T��������5�6�%��Bƺ��lY��8�������@���:�psf�v�]��k[þݣ}�����C9�*�o��a�� ����Ӧ�y��2�|��� �籷��(qΊ�klgi��<�J������l�9�T|�3Bv��nУ���* �M���Lqz��tjH�^��y�j��3�ܼ����{�K��	⻔4��wB4�~�8+��+��ܣ9�}љϻ�����9&��i�5A�W�0���2.���
�ɓ�a����=�A<��w��y�����E�i*^~��G�qs��1�j<�=��3�<=!�֒�Z��4����<��dY��y��6���[�OA�`�Ozl�/D� �wo����qG��O�|}��/b��4�Y���Yk6Eh3�LA�7GaR�h(M�w �h#����J$F&')O���]��oy�|���a�I�!/<�#:�s�����ab	�)�{���7�[xq�:�F	�վ�k�:�q�E�L��p��U���#/��@*�,|7�䭶w~���,[',A��$����j��4v�t���m�7��̋q?h�kkĬ+�oOM�V�W��<(�����\���m n�����a�M �į>8�~�e��p;��)*��v����p��j��!�&�k��l3npE�#9S����o>���8��4��l]#���;����� {�z����}s��Ռ��� ��WO��_�x�P� )�&����M�u�zrO:�p=w��"�{;D�nk�&43�{�A���!m	���pD��ӷ����V3^�]&{�]�Z�<|��0$�	&I39��7�k�7�/^\N�kl�DJѱ��1ٶ�q�gug�;nqG#Ѕ�.7��<m���F����F1�7:�.۶�ۣK�c���#.ʎ��4�Ţ�hR�;q��ٛ��f�d�Yk]��ů5v9,������ltc:���9�ke�籮�����'����a҆x��q�<��h��է���5��-E�)�l�7<����n�l�z�r���]��]������;k�1ж�o:;��6)���}H�m�,q����ͷ�ݽOGa{�=� d����/Xgr������ZO��[�'W"���k����9�=�7e\\�:���q�a[�m�k�J�w8�x�y�C�e��v�)�b��k��ଜ�޷���ʶ� G�q���_Wc��:5�n��ޞ�q۱��k=v+��ݭl��U`�M��ے�tmn1s���u�.g:�����9�z�jW�8�]����5s�6��ua��Wc�˗�c6�l;����M71vz�k��'�!�l�ғύR;:]�xW\�eƷmrt�0�u[n���^y����N��P�1�XK{c&��ft�vws��;ke���_f55��&]�+]����Ӽ/6,���o/vs��w��u/G���6�띱�;vlm���epi8�7�8xՑ8��=����C��=��ܽ��2�m�=���ܓ��d�@Gs\6���xMў�mm�v�9Gm]�cr��)1���;�מ.^=�y��:��Wc�7 =DK�trk���g�5oV�p���q�q�.���x�z�v��;)��:�n:-l��n�����;y�mZoW��d$�q�*�cns�,��y��Og��!SF:��vS�t��>V��;�(O[�D�mg"\�cQ;��`;L�p����na�6ͧfLpemJ{�\8��`���*P�
6m����h&y�5���#j7��H�D������Nl��c�j�Y�/Z/F�Ъ�!ݍ�ݷn�N�����n��'U���>C��u��۵����ٱ�Y��n��N\r�vuk����a�M����q��u7Te6�X�r���v��6:���W	v�.<loo7Wm�+�)8��8:�ͨa�+��݃]y�z]�n3�(A�Ls��S�'lv�h��b���s�۱g���g��$��n{���9ݭ�v4��qi�wlu�9��G9�q�z�;6"���r�Rܺ�y����8�;aW)1�,	�Vla6θP �ێD)�����[6�-�� ݽ�,�rW1���#�m��vl�g<K�\Oe�P�Ź�M��ɋ�ݗ�̐v����g#nҩ������wmoO����{']ţ��l��ݮ����vܱ�{{k=��8燧۳�[;��懋�D��k\�[�'v���+O3�x�kQ��t���]C�յ��v0�f7l��wc�y���;<�:��n�{HStOe�H�O����6��;!���·؃�6�M���]����&�ڼ�uw1��9
@��b��9A��z�/�����y�tiɷ
��Vx��κ�9�#�&'-Cix��:[c#`�f�;l�Ol䘂t��n��l<Nn� f�ˊ��n�����n�j�сF�Zk�ΰ�� ���#u�]�OV�<�^2���m���n4qՔ�}vM�8|OR�I�)}�l����s��5c���oc��g��[q�'�Mœ�1K����a6�B3��X���W,p޷�S۷���m]�toXnz�Ё.61=����nV[۷��7G���mi#�n����ܰա��x�7m�:X�Ƽ��=���`R�nǎ�n��k�<P�h���[�gs�:Ճ�y�og�m훁mdn�c���X�ޤy�b��Ni�c�0&�[����{c��^�^#�G�h�z}V�)�n�+��7p���<�oi� '�)7����\㶣��:]���.��v�qqa�t�3+�v�����8E��[Ÿ�*�1]��kc�w[q��V'nwlg)�Z�W'I{Tq[���y�h��i�lO]#Ɲ��p{`���ok8�m�O�F�On��n���m�����l��9.弋�&�8��u�'���I�����gN稹�#���v<6E�p-�lV�N����ds6ݭ�N
�e�M�������פ�[
�f��ۭ==�ͽtv:T����yx�ܐ��/���&�0�u�ē�Pm���S��x�^�����VLv��<�vp�\�u�^������v�pvm�V�wl��8�m�r"F9v#�t����n7�v�q�[cscnK�a����]��nX��Ƈ�N�۴���DV���uk��s���<vpe}�E���v������s:�9�1��FC�ps��g\��u��.ܘ�c>�n7F��C�<㧢:
�ۆk�`%8�Nݓݥ��pi��e�д9[�U��X�7���B7���$]�%w78<`Z���N�����۩��:�7)^3�v;<���ܒ��q�rٙ{�����=w\�����OG��l�=�g�J��]v솱�Y^�=c�7NCq=�Mi��]^���R0ǂ���q�\)+�.���m��\QmSr��C����c<�c��9�6Z�vG;���s
8�s�:�W��qIɛ���v��Tb��nza��֮6��ur6�8���F�w:Kx3�]�U�و5Ҟ�ug��;�䮸�ٍ�e�����F��ssn�K��p\��<y�r�ݬ�k��]��e��m�^�[��5�:�F�;;���q	E���u�ɇ���	�`�{)��:gr�*b;k��7���:uv���v���^�QN�ێ��tx�GQ���5�=���<��8I펽�nyv�v���̉�LCX9���u�h쓨�OY#�u�nɈ�(�!����(�[��1�ڇ;v������vY�m�n�#v�/�e��암��m�D���&[��^�I��MJ{���L�y�N�퇥����:�x���<d�ih�a�`�7�;4���M�(��� �6N�c/j�%j�g����v���f܄��Ӷ�3�t)��!�у�=PfC�mvf�;%����ʩ�q�23S��a��7]sny��+OM�nC���=�Wy���N�(iySY��'I�c�Mn�Ѥqu�q�[m�ֺ��G�pj�0��Y+�>W�C�k��cr�K'�RȽu��=�כ���{];/c]��v]�y9л�x6���d{7�{j�Z'r=�%EYʽ���m���cmh���]��p��1���n5K���9c{�ѹ=XbDy�Ϗ$��4�j읱](nŐ�:Χ[t��������ꈵؖm�{O<v�&Y� 9�!p�gsC��\����{v���g���U.����F�k+�t'U'`�����o@7`��b�
��6��Y|�R�\v��Ws��6-�����eݝ������$`}�ZN����g���t��%�q�)�:�1�:;����5�9z� \��`<��c�>96w�7����SÓ�@�؀f�ݽ��8�F:�,�]�y���7m��5�rv��_6n��[z�ݷ�ݶ�r���F�ކ�kdO`�ㅝ�%�5^9����냳z{;G�t���&��ai�3���N�xwc��n �<ރ��jE�;q�:n��aG���uU���b�Y\�@��.ϵh�c�6M���ҾY*{��oUr�9�:�KU8��[O�5���Qt�b�O�u\r��;�G�����l�6�K��ZA����n˘����\�<�݂��&8횂��1�y��v�|v. �`9 8��YwD2�1�^:I�Q�Yq;Yt��U��@+-n�5E����ݜ��0����9i�YӟH�8�����]��l=�s�ݧ�Y瓱��mv�gn̦��ʖЉ7#�1{Z��]�ǻ]1���x��{okn..y1�������g;���C�&�d�w؍���vLw'1g�z�����b]ͮ{xq��9��zf��Aۓm�/aIޣ�g�=�]ݻ<]G�"�$�q��l������k��c9�ކA��\�#\#��Yݞ�=4t���Tr<t���`���n����n�z�i�w�z�sW v��ڈ�w�ֲ���m��&3�s�x[Kv�9oOR���`��;�r�+�g�G��Q���Ȧ��]���۞�TZ�]+�톍q�5��ׂ�G�uε�˛`�z�dA��uQ`vm/ݧ�pM\�&ݞ�oa�1��f�Z�w8N���zfU���Q�����Ǎ<i5�����n�-q� r�#{vB�֋�������Iָ�]�\��uU���Y����A*�r���&����;v�u=c�����mlcD�#g���۳ȼb��#�=F���컂�s�˺`գ�{T�I�N����5��5PP<��l:㇃��Yѣz���5f۞�o��fv�4�����B����y�)�.Mt��a���s�X94�1sݺ
�u:7'n�	�2�����ې��9\�U�Hd�v7Y2�a��޳�ɷݦ�[��.��\D����&2���ppVz��h�TX���I�#Lw�ӎ�f�f��T��Cۘ�ix:�[��l6�;���!5Ƅn7�&6��=H[�M�[ֻ^��	�v�f�t����!�9N����j�V�<�9���Sv��u�-ۘ�}�WR���^L�N���ۣ�-j�Z�W(�Mμ���l�;@��ة�68�q�ú��q��}�j�ND1�{f����6+C�s׫�)�V�:��+LViz��(l�箝T���.�:7W=W1��ק7j�j�;=+;e�7>���V��qu㮍0�6c\�E5ӛ���u�qu�\񮽛����ɸ+��x�aԖ�bo�Y{{{��������R��7qƕ+UQe����"Z�R%,�V�-Ycm+�KQPհ�LKh*�11U̸R�XũK.4r�FR�%T�R�pc��Kb��Q�5��i�*��F"�T-��+Ab[F���T�ƩF���F�+(�-ZPRT���c[-������ ۤ3�K��ET-)RUk��0�,Zֵ��RT+
��"[Xe�Z4����lB��!D�(�,і�EV�(��՘�KTk)m�WMF`�E���
�VVZY*Ƣ�iLje����"�-��3�T�T����*UJ�9qU1��ˊ��[TD����Tm"�֖ʪ��3.8�i+�jVV����F6���ѩV�DUA
ԣU��*�KkR�il��rI'8oF9�nb���]C�t��V�QP����U��scQΗ���6P.�]�q�L�n�]tk�*y; 6� ���}u��1�R�9.���g��g�֚�ά�cn���k/N�mPj����6y����� q�3�\ �us�:��=�z�lc;�W'at����=؇���n����7:�g=�t���k�:������c�#���y�qWV����vT:�on�8v������gl��n]�����{	����ױT
vw���u�힗���Kۃ软�����>����G=Xn���g�cɇ��tp����z��t�u��ra�٬f�k�n�$f�<w8���(]�p\�]^�ў��N�]�OTru�Ԋg%sWlr�@�P��[DA����y�����dVCq����l/Q��e�Y���wOlq��61/[��;gx��͌�.ڇ�	��ec.q��n��]��81��(@d�5��y۳�H��;[�y���E�;�ћ��4��}3�sb5xZ��y��l�<�l�t�.;Q�7��8�l++�l�|�b|�q�K��b��ݲ%W)[c�V�*k�3�N��]�{K�s�9qӸ�'=v;����ɷM�v�I�m��9W����&�cr̅�n�R��s�N�lm8��w!��lW���q�X�e0=�S�`�B5���!���<&��-#�/h7]�;m�m٪��N�Ss;[�m��n���ۏY�^��c����z����}g�����O\[��X��t�x���.�ý=��4�-�8�N]���&�sq؋�u�#�+)��գs��:kjmnw6����s�t�<�"8u�"ka�v{��Ѩ�(SC9�y���}+�le��Hz�1v���5�c�v7%�5��i�v9��d6�v��=�V�)�dy����9Nz��j��okh���5�3���v�+���l�U�-�(Wg*�7U��uS�����v���@���Z�(�0�C0l[�\v�m�9��Ñ2�1����;
�U\����������[�Җ֘�PX��)K1��p�pr��aNw/'ݰ���O9ANǲ�x��V�1l��[�.QG���� m��m���lp�9��+�{l=��	��q��+��e��{
��0�
��'<=��vp*>.ݗ��~�����?�'�[�V ��M ��$�p�a�9Ӟ�(,}��Qy+Q � �U�b�b� ����agN�ܝ�%z�v���(w��2�
�q�37gr�J'��[^�A�����K���L6��ꗻ��r��� �݁��P���OڛXB,�ߧu�l��z��@����`<gL:����W�;mtm���Z�=��W��7В+u�+}��W����j���ˉ티>tgTd��ީ5c93�v���	"��]��*���0��>la����w9�0�q\�xs �/q3J����0s���]t�� W�vܓ��/cu�r ׅeū�ћP��܄��Q��&��i,�S����\�/��b𯏒�q���^�}w{ �U����5��l�mژ�V��YM���+�N.�|ם�ʳ�r� H8͘t�@{�M�wQי����y�Z� �1���ؾ���@_z�����=�o}1��\ ,��Hu{�N+��-�C� �P���{{�zbH��1D�oLP |U�۶�~���\iuE[��YR�6�W6؜��rZ���T)/$���ܯMewI}����6e�{92� *�ݖ�y�m��ՙV��*+;P�R}�dȈ�$D�2Z�#��x��E�݋t�K���g]Wmj������5�=nfd����'2f� +��X  ��A)'mu�ٜ�[;0e"R���I��(��0�~��8�d�}U�*o��K����� U~���>�tݍ�'��a�O����C�Ğ�Ƶ�PO»'�{����uՀ�&�������yn�=���2[~��.kv6��ٻm>�w��)��Sn�{4~]���4.�D��nC��<�u��-�#&0cv�5F�A'�INn�����>��j�H)�%D���L㭊ܧ�n�5i {;/�>9�&$�O܆ �>�/�� f�l�@S�i���I���$]�}{��Y��zf��uD�NG�*�s3��͊�(-��2��+c1��v��ߝ�f�Z���d����NGc����v�۸���%�������n�w�wv�%������Ιt�vf�������9�6n�3|g�m+��C��Q/虘".l+rf����M�,q��w����lݠ> ��_ �(�:I��滽}�B�8Z��2&Z6���>��L�6D9���a�3״I$�^Gz�%-��$̼]P��p�'�]�l��J�f�ݭ�~��u:��| >�zҫl#��.����F��t#3(E��&��X��:['*k5�9��Z����^��1�XN��<��V-M�{L��f_�j`�!��{�����Q�f�j$i���Y�I{�V�A���a˻�6�f�@���x�5�Vw����_|�M�݀��.� �ٽv��%�'�����}���_��X\C�R���x0u��]����=lNqŞz���n�>�e�!��^��V �� l�f�cc�o]�躺�޹���;6���N8��4)R�9,�����m��>�DE��-���V lFg�] >���o ۇ���οGU�=OoC\�Q/虘".[���@ o��x����ʩ|m�X6$fuK�@#=�ً�]�+�(�1D�B��8ڿt�_�D_�� }�3_ ���;s0��t��㽎����ɗ@}Q�\�ħ���o�k��`؁�{��؛��L�z��uZ��.�z�w3 ~�ekP\�odA�c�E�y��L��]wV��[�ۦ��ݝ���8�1G�.SԨ,�o{����^�8Nb��}jL��S��E"v�0������s�u�4��9��wY�:u�ֹ`�$�s۞;��h*��^�-�������Y�tt�\`�;x��=x�uq8�糑�Y9x�M�����j�r�bv{pqix9���9�!ٝ����H���Nې-ʙ2��/3��84���˕���"����Zn3u�:���ni���2�Gn{d�W��6g�0n:�j�@m�6v���ݝl(��R�l^,PD����6�'(Q1��r�B��G/��zg���u���ߺi�8��lw?su�2� ��nfQx�P}$�RC�.���Z�Aw�����_�z�u w�� �o�7��A��t�.�
|�y��)R�9,�W�ݙ�����������s�J�{�-���=٘1 �o�6�^�9R�_�2I���37�S��n2�/��|��Ͷݛ�R�����x��H���ń���J�e��`��v���t�$�[+-V�O�~�����f| 6��v6�s�[}m�:���Vw���_�vv��GY���i�6n�����F����ݴ��+�5V����g��|����e�V㳍���x�@��֪���T��4�;n�s���޽�o��tݞ1Z��"���#I��p��'+6�"]�{r�n��]�'"�^@q�X��;����o8��ȍ���f&���U9����Qq�1t,��^ĭ���Vﯖ >6��v�m���$OFwG�jsj}3�b�u�S�Ϧ%K��voz�� ���4���s���^�����M�=Ιt���hN[R�9(�W�ݖ���`]����'��� ٵ.� /��D���Ƹ�N��k��HmZ`0��Ďa��V��|@ ��m��=�s�h[���uޛ���ˠ 2�ݙ��Z/�s= �:t�[���kf�p�����Y���u�e�\��v�M�����B�CL��8z�ҫ ٳ4�A%䮳z��5���>�:މܙ	LV��8I�l����"���V��Üͪ��Xom�4�ꍧW�� �������� �a� S��`��ۉ� r�ݝ� ���i���S���e	��{2EY	�1�b/�s�ǔ`K��j@����0unM�S����VD�=ض_s�J�W5�5]"OF��z�[�H���ń_�$�)q*\䊰{{�=�y�i�Xs�t�,�LR ����@ �o�4��̞t�ݶ�wP����͡9mKp��+���X�v�jj	�:��}0#XIc覥"R:�ۘ�m�6��j����/c6d�F-D�7�k֤�q�ݚ��;�9ۍ��g�s��ￛ����o6�w���~  ����։I �/��-��v���ح�[����٘�ĮP�P�,n����A^�ʫlLd ^v�` �gM����{��SκOn�`��n&!2e�U�z��3 {��l��ꃑ[�sp7����%� �7��j�z3�$C��ʗvm�p��t�m��=��^Ej 3�r�� ���"8�[�Q�9V��*��Ũ��8W7:���8�V��D��(r�����ˍPd"����ds ʽ]���������b���9"�|�:���"<R��X��u�6-���� A�Κn��rg����Gv�_����(m���Y�0�^q��H����9����v�=nA�6���7|�>p����6�}���fګ�#�po�˫��=����`�޽�##R�F��31�S�p�������!�s�f��+�Bs�Oğ����!�lgT: 4�$V�dx�zk����q�5B�CL��dz�� 4Θn�7[<�T)+�*�� >�tڱ�-��@T<뙙��b&Z�F�_f�_u@w;7����6�s��̌�� _���8�c�� ���6�Fe�!�ʗvl_L7_ {�x-ty㙐��t=y�$��Z�a�d$����W��]~�	1����L˸��E)�cj�:��Þ��P�Tt�hAm��]��D����.��m�dڙ��w������&�|�	NPy�y�H̺���5�(�&�wE�ͩ�t���v.��:)��ɨ���y���wU�TnCQ�uǠ/ov���ċ��it[�K�v��V�{����t�v�y�n8-N;���<��#>ϋ6�lpt�/^\G���6�ݽ��v����{p����5m�̈́���l)�'�tm��NqZ�V�k��]���!뗷�Fg�n5��n煋����&=d:���ы�#�ٗ��ߧ��Ź��K�m�ߺ��<g�� ^�of`:eH��E'U�6��M��0Θu��VF��pe�쭴H�˾������N����tg� ���y��$t�ۤ�vg��$rq-�`8>pc����[�I��<���Ѐ �"__3:�g5 ў�m�@�wf,!��9B��L1�dz��FU�u��u���Qy1_ �-����>��л���ηz�1n�Y&D�Sq���
C6os�&B$z�ϛ�iX=|}TgL:@|2�ݖ��o��գ�^&gT���t�Y�CPZl���t]�����۞D��1��釛�m�'<����߀R7Ɇ�K�6/f(Aw���  >7��v���[.s0�ݨm�@��y�>O�x�(f�CNj�"�~y��:�^����W��v�'C����Q���\�4��I t~��z��Lu7�A�V��oV���
h�rdw�{�7f"뮶��nJ�	<�v4^�{�כ�m���7c=z󫼣��|������r����e������|76j� *k�W����a� /��3 p�'����|�BЏڂCO&{l[�5ݎGom��� ��e�� f���� ؾ�u�4ڞ����;�����<F�Q?q-�e��ۚ�/����.��< ;�;36 �{fՌH�/��\��Tgl}�T�r8�H���ӺB�E�6ݴ�e���zE%�a�[p�����q	p�0�/��ۢI&��k@@l_T:	��n�ۭ�e����ϰb�f�tɉmF�K�6/�+���g>Ι��z�}����vt�� nz�_ ��޷pg�⻻R�o�$�Ȣe�K����s��@ �Ǥn�)%W��S*'x��ޫ'�5w63��.�5�>j�Ⱥ��e���U�.�u21ݳ��@��
��[�#](u�1{!���]`���U�rg�&9����U�u`n{fPu��^��E�����Iq��z��m����o��r��g���SmxZ��91^�{��Aܷ��4\��Ln���C�=¼/����v>�v��i�<BO��I�Y'fʳQUU�I�:���N�J�>�g���˷�Ta�!ST�j�3G�V(�/
��np��j۾�d�����j���&P�C�J@��b���{���,�M�a��⋄N�g�;�KC3�f�ck* � k����8�r���ڟ0�<x8�޾�G�oi�&!��}��om�e�=��=3����W��{� �m�^$�wz7�z7i���K�uj����ɰZ��Lѹy{ڽݔ�A�O2��oy��ݣ��(�TN��v�֩�}�1w������=�;��nv^Iӂ^@o}8�?iEr^ɇu9�/w����sL�L ��Sٽ��=4ÃM���u�����Y���r��U�f�����O-�z�}=:+������^Ƀ7f.���Qo9��r��{h�B��^��'���|#L�<���FR��,HNXV�e��Z��527`�w*�8++x*3e��gۖ�)!���%#'�����[��z`{-tUb=z��B�܄5L$�VeG2�,-�'���v�h�j��c�c{s�B�;�Y��pt��s�R���0Ohuf�;��Hfi1�3�IA��$�j-�D��P���������V�E�K[h�ml(�T� �jҷ��k1�ӅKU��U4��Z�(Q���iej5+Z�PVҵ�e`֨%h#�,�Zʴ�j�naQ�U�`�J#J(ūcJ�5
�Xk�"�D�T���K-PkT��յE)JZ"��m�hQ.a1��&3�&��V��
%�mE[f����H�R�"%�,TeK�ps)�bņ	��pUKu��kX����#lZ��ֶ�J�B�+�J[Ik[jVT����kJ�%m�Z4���b�[Eqզ
!K,j5�)�qL��-���uqT�U*�[j꘹R�T���R�,E&UTR�L1Db��j�.���)U�[mKh���ƈ�"�J�)��e���*�EQ�i[����,Z�����Ɗ�T���(,D�V�
TSI��Ң�B�V1Z�	RյJ6Yt����-+KB�Z��mӂ�"�ke���"���*�ZV�j�-�`��1�-��
UckmZ���"�m-*���Dff�f�aKm�#ij� 6�m?��@�b��]�� ��j� ێ��Rx1��N�(�e����ل���J� 8ͻ�m� ��ht ��{<�H�W*�og�{��O��d�����(��$4��U 		mfuX��z���]���wrK����w��\�������ϰP�78C{�����*֗xj�3�d�j���y��ru5����!@�3V�\r��7�~8(�]����% ���v��WtD�^Y8�:tN�e��u���(y[2L�&!9�A	��f���9W��}S#��DV�) � �s�:@|���[x
�)�\�z�5�'.ΘRX�@X�x5�=�@]�m�X6 ��r��i�"�*3A�u��R z�ݘ���(x�Q2�A�tN-��QC��8��8 odI�����P6��w�1a��ѩ!�Ne�;���y ��ȩWR�'���[�1j��͊�ݛ�L�S���&n��z�p9n�P�Jpi�w���Ψ׆Iy]3aH�x�[�R��]�ս�Ճmٹ�7�)��lgD��إ�!$��'����$�/l��Y�qz����~W�v����۬b��[N��n<�>mp�\u�V�V��7ձ�����|Y<�	�k������� >�q��m߲'7�yp%W3�H
��e����D�Ķ�����Z����'-�4��#�� �~�fb�E��E�
�w�kZͯ^ׂ�u�$��b��
�U�b���jl��������� �*��1,�E��E�d\�Q	`�`A���&��A�"����u�� 
�ٱv�ng�q{�A3Q�Z���
s�)�Ċ#5l�}?<L�'	�v��fm��݂���vFW�_�31��#�bՌ@-��
�b-�	�.:ڸu���qYy]�Nss��B�TN�K��t�h���4��։��շ[7Q��I
/W�<\�n;1<�P��@��nF���,Mc�6�m��� ��Kr�v�wE�뉵��ͥ;�b�A��`�@H��sf.{L{v����<q�Gp:��(������ǂ�㎺�fێk5o<�=>.���UG9��2l{*�m���G]��`s���rq��Gk����q���m��Z���m���1n�v��`��덞�l��]�W(�ۮf�+]7f ��V��<�ɐy��m ��h_�[�.������>n��X�(Q.�Ewv�,�ڛ�m��6�3mU�(\DӾ��� ��t]�wQLD��LASezc
�۵�T'p�=]z�>�������2�i�S=׼�P[��G;e�aǈ�Ki�h(���6�8�  \��vOFM������g{f�b@-����z`�LBs!V7}����ί_���$�2���<�w�����{��ĕ�l����2.�s2�� �K�6�8t�^������(4��u���2%�{	>�{�0�R�z���u���N�x��!��Yy�(�v�5t\v[a�R�:�6$�Br����S�j!D��@�s��� �[x�4�D�nuU��T�0����'��i���g��9O�sc�R�(�e���n�i%�����A�s٧Q"T�f��md������(ȐY�d����޸kez���5�q�s���ʔ��Ww@�6\¨������~$�g�_b=��f,��,��׳��xdF�Z�Nj!��0}�T�ع0 ��ט ����D�幛�^�7�Q���v�@|�o�3��8�
'�'�v6����1���q�ǐ�S-��g{s0�{��;���<Ím��ʦۥQ�z`�LBs#��jo�Bs	?�o��`�������i!��$�L����b�IY��ԫ^Fqvd�[��eCC�'�\!��K�aF�����˙�h��0�\��9�_���6���)�K�{R����,�c��F��Q�y9S�O$�Iv�mш��E��IC�q^7:�π�:�]��5_���]� {���� ��{�Ռoy�>�U^e��7�r���� �(Q.���ۘ� A���W�*4u�Q���7rֵW�<��z������^kAW:���}��M��q��%@oYwݽ�� cbӸ{D�0�C��|@�7�y� Fǽ�j�ϴq�1�
f��ܩ}�f{��]���"� #��x�=�n�{:��<����z��Q�	����cq�(�"Pݍ��b�>��2�G�����n�n�+�����(-y��	!��M�|���v����!/�Jr��������#�魵�!�BaziYWn��ι�L��Q1��0L�&!����F�f��5fuz)$N��FB]���5�ި�͓!	&��0� ԰����X�3�
|I#��8n�ޚ72j6�m/$��ٱm�nGH���MF�z�͊�"�-�g`����ʿC�C.�	j��Sg� �G��7I�,�����<۞��>#�����G$���%H@82�gvS�ηwWٝ^�l
/=h3&t(>=}���W��
��fc�lV\<k�\V��WRфnI�흳�GDQ�5���$)`���n	0����@��P{� DotS���8ؘ�pӅ3sh��¾���o=ט?k�2^GT^e����o��n�&t(^�vf��z�4aﳧ����*�%
*[V��ˇ�9�U��M�n�<����{:%����ߧ��ظn6�	���>ȍH �{��ʎ����"{"Ս�nL�) �$��&G�ĈWi�����_�f��#3�l �3�@�W����A��%�����Wu��̺�uҒ;�!v���)@ n�{o�_ٓ�[��ُp��g�H u�w^`N}�g�!�e�uA-[}��3��8h�J��)@؂��������hj=睳u3ι�ff��
F�NLL'�(�e��ݹ� �L͊�g���6���z@�D`P����� lft]��J��~_L��I�6o�2���龾�}BՔW��}�:�:�==y����}Zs<ߟ��Ayu���Ӥ�W�hh1���ۻ�&
G�8p|w�!�wgb�yRΞ��\�˵��	�i���}����n��;p獁��:Wg�����y��O�.��W�|{����]v�hx�uXD���]�bK^|tkm۝��:\�k��	>ڍt�hT�8Z�9�y7Np^��ێ�F��=�j���y�ٹ�A��΅�w\p�Ϭ���L㋫>9歳]J6mX��_A�5%lq=�9��Y��C�:��.��<:7Ey��x�SI�� �u_>��CP9�O�V�aP �{��m�����/};t��K���2g���Ww�1`8\a�d�dD��-�6 �gflF����dE��7W��@|���iX�Cf��iyϳ	࿀�.]dA28��$L![��������jlH�#eQ=[��E͆ �n��� x��xz��'P:R[��f�������;�d�0wI��wf��I����7"86�)�vF����m F�vb��3�f}(�0�\]���{7i#��e*I����0����@&pݓbՌnL�PD���6��+�!*�w	�����a�;u{��EfGZ�͸�ܻWd͹�e��k��%ĉ�
%��{���zfmͶ �&x(9l-S����w��o> ��ؿ�>s�tICP9��
v��d��]�!u�т*�ȹY9��B��=�κ�-��x�_gK���e�9�;�Ơ��]�d��Z�&��c�����>�_�  �c3�]� ܙ� w������Y��J񆍒1��迂
�ڛ7"8� #6�����e�=��lF�gE��7&x(�U���b�0�n6{.O ��]T{2�MP8�˛lrg����^�vS\������ȦlR�̄9���r����)@؂�}טt�=F������M�ȎۤW�ݖ�g���ѵĸV����mH�a)Lr�bM���v�絜q�񎹷&��.Gk�l����?�?�W$K��vm͟ �G�@  �����w<��w��.�Նg��A�O�� �oG$O�Q.����f, ���b��g[sb@|ݑ>e$ ���1`���l8�������=Q�f&e��͕�㯠 A���ϰ A�9؋R�Mdo]Ɛ�ɦT�{4�q�=�8r{����� o{��s�:}Q�\ �۪��@�������U������G� #�2�=��U,~���|��^Ώ~@�#�(=~��1`9\x�F2"Pݍ������k#���{��F�� ��fb�c��vU��*T]�8@uD�����tA28&	"a
��Vn[m�2�R���t.y�,Ȝe|����v� ��gE;���>]�ޓ؁k�j	q� �ڭ�H��^%꺽vz�n�v�#Z�0F9���Ϝ�L�����r��d���m� �C^_:��<�'��<'<��L�#U�۷�M�>n3�2���a��EZ�Y���G]DDق9�ty�'+w���؍�gE�}Q��<����g��O���'�(�e����x�=�jm�^{Ϟt�]�۾�g�@/�^{s0b����S�Tr�fe��M�V�a��z�a  ���İl=���_�~囝��X�GէwJ���k�vt8i�@��4n纀��q�b�<�L��LT0<�#��->ݭ��A�����^]�N6ӿ��v�4"��x ���
����ߋ�|�$c"%�i�`�G�r��^�gUt���J�/j�� �ř��V�G%>HGz�D�y��{�A0bj[�9��F�77f+�m��`GC��6��1��+��H%ʒ\K��,㦳s0> 8��)���8���5)�:m{�1`�7m������@�I-�46|��=�� ��3�[����[��?BI ݷ��@ 7&xnc��Ù�zvn{��k���>s(� �qm��6ؐ{"<W� N[F�ۭȽ����I#�3�R)$6�8+�>��Cz�8�8iĻ����>Ͻ]��z��km龭� fL�P	�{����}�̀)�/�x�*.o�In�D%��g��7���9�����o]�]n���>�aՑVѓ�R����^�ۙ��G�"��}�2c���N��j4v�,�o��7�ry�C�VZ�̅=o�R��1q��vx
8n��?,)r�Q��,��bފ�|r�Mʘ�5�w}Y��t�+MC"d��Z��*P�B#䮥��Y��M{Yd47z�eAvA"�A�x0����zy��n^�E�rX"Ga��2���Z>�	�&_m��;%zvC�|B�tV�B(fT������qDX��7�F��ؓ&4'�8�Wq�;�짵��	���S����J�E\��-���oNd������3<H��N���53�7=��}lY;p�Dc>��:��>z_NF��z�5&��щe��/�\Wz7��W���j����S<n\�p�Ȼ' %����oR�ߜ���q�����3��A�oط�}�N-�g�ͣ�[���m] vQ�{��+�:��
���<o� 4 n�G��$�[�M���S��K �d�G=}7,K�l=�j���}�4 �v@wdÛ�f��׵���僸XS�Kj��ܩ��4n��X��^��'M�s�J�T�Ǽ����F㎐�����8{O/���65�I��)��F�ܶ �@%��k���.� g��ݦ���?GJ2����8�f7��A��觯����,����!�&y����$�OW�^�y�.E����3�]��o��N��Ƹ{�$�:+�>��d�,��^)�yr�#�����돠��<�F�ݽ}�8s	'�ik*-Qkv�`�JV�֢�V�+KaTEEŪ(�VK���V��WR�V�VQ�)Zƭ�+E�Z+mQBڥh��JX�mFؖ��(��ZT�[E�r!\F)�G�����e�X��jZ����EKlKUƘU�Qkm��R�iTE-�[h���*�m�X��X0Am�Z��fih��5mb�	X-X����\�[Z4�h-��鱌G*5��DZ%�����ҵ�X�F�hҔR��DiU+j��DeJ��Q̸��m�lb6�бFZ��Ekm*X�P�,F#U�УV�b*��Tb[eK)J�EKh��Z�,��-lm��F��ֵ�2�U�2�TuJ5V�6 �UJ�5�[c,-Z��eVT���V��X��eƘZQjA[h�ӎZ,�+mD-�kj�-A��X*�����b(�k.7.���F�(����DX��E����Z�*R�[mJD����[���TfZ�Rխ�5j�L�������#�R�ڈ�eQT���e�#�l�ƅVTQb"�DlE�*5�",J�)�?7�@�z�ыM��a���g���8���ց��Cj��c;uZQ�D����׋`#��e�lq��5���nM��8����nCCB�i�j܏l��K�3Vӕݡ�Z�kg������V���N|6�vlo����5�;�ޞ��M�ے"������E�6�6�\�׮Jk�{4zx��=s�s3��ɖ��m��NJ�۱a^�kNo��k��rk.�tpfݹ���-&ݰ՝]��[gF�u����\bv�Hm9gN녥�p������S�zT����wN��`��4�I�a���k�ܲ7��޹Ͳ�9滲j�qʼ�՞��ֻ�.�0��;kf/5�b�.:�:�NGnQ�w{�*�)tgQsv��Q<r�"�voSS�:��v+Ѕr�0���3��wM�9�k���t��x�랅l��8�qq���`{��7v�6�ܘ��{��l�u�ld���`�8��N}rۘ�q��|�O3�ٽ���Wm�+��Kx�ڸ�b����E��I9��v���]ym�J�M��j^l���)�,�r��>�޻q�rIEs��0,�gm�|q/%��7cFu��h�ڃt�]gt2<�$	�n���#@k��Y*s��8�lc 7W[��Vk��-�G��^��ֆ���k{AW3ڮm��������b�N�Ɂ9�Ǚ��weG�u%x�8�vq�e��p���b�
�6�9�,v��ۋ�:k��>�%2'ix�kN���������L�ޭ��:������4���q�^��G7�(J�DFܩ��;Y�v���ý�Vޥ�zv�Z�ͮ�̾!Y�c����nS��L����j^{n����l㝕xZ؈�m�BE�<��&u�|�q�:v .�H�N�X�9�۝�9�o/kHwF_2k��=%�(�r�N�kx�x+�3{O�u^C�lCՔ��=ק��;uu����!"85 �D���+==��H�=�\j�MM���V̖�	 ���m�Uu�\�ю]dz=��ECfw�	]):�S�_�u��I���z�V���"n�#�<v�0�M����=��;٩��p�=���[�\����p2���[sg�l��8&N�D�ms:-��==��F]s\M���ƈ����F�А�X8H��ĘKpBr�c�4V��]��۴�{<ld�eιq�NvW\I�j�I�8�k\Tջb|�μ	����V��� ���I�u�\�u�\؈L;s����|>�،��6��)����:���ăݚ���"��n�[= F���RZ5,8����O�8O�ͩ�Wl؀H���P�{;������[��v2sv26!�In�Y��*:= ��m��}el�LwS]�޸����2= ��ى`M}>n172�f �svnu����m�[�>iy"U��]ߒ%�3�nMa���H,��+���C~nH�	ĺ-)����KVfЊ=n�KsJwvl�ϧ`�lE�n巈l{����9�����������.c��:��#D{e3��];m<��`��-�ul~�~o��t0��l�..;����Ł� /�=���]�tt�ٛ�op�����wVd�~o��!���
�`p�=.�Р��}�Gj�Jt�۞]��w,����]F_^����B�4*�%�^�q!ݳ��'3x;v����R�ry>�EE���d��{��L-�K�n���π@���E�Ā(�e۽u=|��%ʂfa��ٳYً O{����e<��\mA� .��3|6=���#,q�ff"�uAk��+ӏ�j�K�������ڱ` q�ث@ �2z
���U6t�+�l��U{s>�QO��M�*d�%��i���� {"<T� ��=1W�}�#��v�� ?͋��}�=C���y�;��=��i�10�̄ ����{T��.nt�;m�nܜ����������������%��ۛ}���lU�����1�J���]�f`ϐG�bՃ��]*"%�R8��+g$n�U��,Ռ�YՆ��em�'_9�����:@|F�2�:�+���o,��<��L0"%��W�&�nGII �}�񯻢+���"`���z��'���I�DZ��P���һ�F�%/XQ+�kC��r�*�a���PՆM�L���L��𫊋���>ϳ���_~@����b���C�F�(�IPLD������:ƞ�܍�h8�ۛ>�d��z�ݕ��Z��U;����l������Q ���;% lA^ͪ~�WR7�UW��`ؽ��:�����ޯ6t���0fi��~+ۘ�$	Ls��!�v�<��[��lų�&�~�����m�1/W� 㳭)�̏H� ���1����?ͅ���vۼ�O���٢7	��"]�W�ݙ��a�{
�A���M�.&~$f�ĀMwߤ�����L�Q6*����Ix��ڑ��\�+I�_@ �oݷ�` %w-;[���Q7��'�� z������=��(n�/�<y�GDh!�c�� �����@ le��yb�)�E�GD��'p@P�^�:�XU�^�T�,�c�GoO���/ޔ�]>18��Ώ�9�/f�4.��H|=�{��~�R��rC^�C�d�LD���گ��� �Og�S}��6��+ 艸�@ y}�y�ǳ�Սx�ޛ�D���. s�9#F{�g�lI^Գ`�s�ua')
j��v�����fp�7�L��D9P��A{����o A�����W�ݑW������e�P	����倢��<%	ĸ�Hs7h4��Sg�ꅪ�E�lx�Cπ@-���π ��tZ��.חïk�x���x�K-C$��ү)�λX  �ٶ��n���1�h�kә� u��f�c��vu�t�bX��J�����J���p����$��mQ߀���ػ@|،��.�R`��y�;� {��^,�� �T��0�'K��I$���tB�]F�iل���� �>=�ݠ6#:"�)\z>��X����h���a�ù������������Z��v��<#5T}��[��͞�Ǉg�Z�.v]2K�㼭R��lFd	��6r�m�}�z����}�<^y�u��ѷ.���9�[��q�m<�����6���q8���6�n�
;��}c���;��r�[lgK��nk���O>8{���n���v�8�<g��]��sn#�[��⇍��Gn�0�5��ؖ��;[+�m�&�m�r�y��v@�nm�&:K2g���������<;�=u��']l[䓏'[q�I]j��7E�������ղ�&�X'	�����r��8J&;�w1LCq09���g������ �Kb3�֧h��'��A�����Fǳ�ՐzȈϡLL�DH�՚��� ����آ�z	���}�ǳ����Ctv�+vܕo��]{VG<%	ĵ,s5a��\�`c=┍�!B��<�wO�b�߀:=�݆��E �p��pL4�쿑^�v,};�}ʺ�����ؐB��L��K�egu�A�'��=�e��##w�v	<����%�P8��)��H��m�׳:�]���>q�����v[ybg`��C��a�B�jE�'N�
c
�k1v�e�.ix^���%��=t����7�|_���s��H ��ٍ�{z͈��F��Wc>?G�Paor0�D�&$B�6��3�Aɽ��Wd�E�~q��ެ��b�(Ł�דk
�t��Ŭ��т����B'S�x����^z[��nS�.�Z��z+��P�����9���=��([K~~�ݶ[o���شRC���|�7SuZ�Ԑo)n��q$��DhoPv"I�_�B~md�^���&>�7�� ���� >�z�����C"P�)q2�3w�Z���l��r#r�Ж�tf+�Ugm^ �G���UUz�m���:|�wYc	d�gŸ2�Vnu߭$�KV^�QC4�v9��m�	!�#��H�vuQ$�ǗνH��]j�}rGZ�Յ"~s��+n������ў���at��=o�c�ۈ�;������^rd��k}?�� ߯ݷ�`| �gE�K��4+C��M�qH���ϰsވ59P���DҠ�U�B(�u�ә���wr�Ój@ ^�s3����j� eϧ,���������$��bM8�74�H#��=U���@ޞε6|����S[I5�@�a+�ڗ�VULd:�S��k��q�ж|�w7�W����}Fې6I�\!3�#z��5r����r�lJp���j�Y�jI��x{�xB͐��$����`>7l�׌���ݟI$�Gt6��Ȫ<2��;؝$��۵G�D���6�}�z�{s�7"�r�,�6��-N�D�8R�e�f� �s�l@�?ygb0��:fs���O� �g��I���W&{�ox�4tq�����+��\R붯c��Sp�GS�A��+9c�sLc��2�$�Z�pu����$�՗�f��P��{ђw���~���gf`�G���S�I3�0pH�l�{J��A厢\�ӎ������ l{:-�Ij�����Q�ڕ�יix��f�*2"Pݍ�z�l��ޕR ����T�W�Cڛ��p ���E7h5��E �� d�P'2�B��=v��s�u�w�@+�*��/�QI$JWY�{;�s5�ȡw�[��uX�&���<c��.��Od-m{5S�}Z��$��yZ�;�/H��&(۷Q̳p�P�V�G���޾4������o�I��"!�l�y|~������M7b�t��������d� $��WY�w�Ca�7ɸˢ��<`�m����A�������l�ѫ�/�K�ãd7�Y���9R�e�f�8��Sg�?zU) >e��3 �Tʙ�Y2������9�Ң�PfC�m��@�4���V�IF�u9\�؝���r4'��lH <w�Ea���ϰb�͝�#"�;�T��#�"y��pMM���*�@�߻o���ED�}h��������;ԡ�@|e��-���j��I�X@e����'���?���7�*�� e�nf  =ol.ل�{[�~yҢ��^d��̹��:������_���O=���|w_fhV҆�e��3 �tP�C1��_F`�7(�Zx��Xt/oy��q����핏vr5E�3<}����gK&��m��ǹ�_f�'�w�j��+��Ż��d�ַ��쐁:s�S�(�F��[u�֪�.Z�vC��-rR��s�Tk�AF�\eH73�`�b���l��$���T��و���n��<q�m���xjϗ'at���;�$g��Eۍ�wv�q�̯Ez����yq���;\<ְrݷ"��[�y�u���Gx�f�@�֭�dw	��G�n��vH{k���m��� �V9i6�<]����P<뜝/*�F`ḙYۗu-���Nۋ��Nx�5�:��юk����/�LL�L�~F��U#b��^` >�YoU-W��wR��^v�`E��J �`2�
1N��إ�Ea�gvW���m��3>σ���� �>��t�<�Ѳ�~~�q��D9M��tY^�췀 {��J��=��&j��.ww*3�m��z�`�o޾��{^O��'�ķse=�[1�nJ�!�o� ʻ�İ @|���݀��:�D�լq��U��u�Dj�s�8%�`�w�X��5�J�����6%U����30��;׳v6Ŧu(��N��_��v�����]�k��9ү/m�Dy�q�8�7rV
S9i;3d�<+�H������˃R�B�����g�	 �����@޼�QH#<�/^>�����ڻ�f� ��Λ��#�𤙉��#���W�>Z�㟳ҟ�o�S�#˓���/��9�Y7Co@�3�Jlc�WW;(9kc= 	�ˆK�y*�u+���T�A����E�Q�1� �Y_~����YY+*_�{�ng++<C��>�?�lY�Jʇ��?�wQ��_����#{/��|>#��� �ABe�cf��Jʗ����m�d�e�əf0����<,�&8�Ɏc&'u��}�=�����̟��q�#����g����t;d�W��pC�y�6,�q�3��_��S0O��^|ϼ����l����ۙ�=�~eg��Cc1/<�:3����J������I83�,��y���}����ogo�%���)S1�13��}�m�u�/��~�Z�J�9��Y4�q�/�9�N;d�d�&6��Gn}�g��^@���&eM���?'�37�<�6ΧF�fc1����سHr3�`�f!�0������a�>��,�ĺ���y�\vng�F�u����P�盷sי���l.�-�1.����s�Zu-�tb�z�I��1.��v3���c&e�������Ͳc�c&2�T���?}�<ed��*�W�i�-g�G��y[��'�k�g�������b�'�L�_�/�un[n�ꗐY�J�����Y臌�b�C|Ѻw��vq�%�|��q�����y�{�4��3c��L2���N{1y�y5�}�s��5}VUp������O�"ϼ�b#�&��B�
*L�N�}~�����Lfd��{�����c%ed��d;ۯ_��;�O �J7lД}b��=��}Tc7�m����"���'�:�L��rQ�����fݩ�Q�LN�Q��;��3��_��������lO`s�hJ|�^���2�	��t��:���3}��n_z]	>`�+�:��V�q��~ �#�V���ޛ��%{����\���_�2��.��K�d,FFq��"��-ژ{�bA��Tʮx�N�ٛ����}k\�gs���?=V�Ң��鍿U��2aMn.�<aT���o�ب���#�p`�J��i�ؔ��s���d�e���[sm�h��*{J8���t@���*Df��Z[��/-���U�����yU㾗�T��Nv�4r���c@%��^\�jݢw5Tc�����X4�Q.Ц��Z~W8��43佔i�*�|t�&Z{Y��"�ѣ��a�R�8�t=�	��D�o�p��I�6��9��˻������l�b2L�ʌ�m�e��y�^|ar�֯u�|^�'��Rv�"r�i���D��N���7-=��]O�!�����`<{��{�Ұ����3mn�%Hv��N��N�نͥ�ޞ�0f���ݭ�o���tn���@�6akh�e��۫���F�=�ۜ��wo:��V\�����O��nQOыM3������?ry�L�g��
�y5�DY2Ay�{^�|�Y3;M{��w�-Ո^�v���{���5����
_d�Je��&Yrw���XM���%�����\��U���ק6������0p�(
EkX�4�(�b��$�V
��hb&)X�Z[J5AX��}�E�X%�F�Ԃ�-ed̹����!P�j
�-�"�"�kb֭�EZ��DA2�Q�(��J�q�m�F��V�fS��
 Ƶ�e��Y+mCJ�`*Ȫ8�,Dc"�DL�\AF���#P�XT��֦R�5�V(�R�6֭��MP��
�ZթV"���J���FbTU�Z����5�d+-�`��
,Q���X�˙eV	m2�b*E,*[dAPU�Uq%�c0b����ZG���C�-��Ƃ�K�E��R�[�(T����(�F��E��)r�Um-�-Z4��ب�����W.���+m
�uh�E2fdW����\@R�Qq��E[J�,b�mKj�d�ʫR���-���V��YZ��)JR��h�j��(QUb���m�C���mUHQQEJ�j��ڥ����j�Z���
L������^�a�u���VV��ob�!�3�`�f2T���o�<O�2k����t�.kMb��Y�ϙ�>������q�����ܳ0�1����c�6Ɍ���Ld��;���x��+%ed��)���ۆ����=�Z�U^vM2�$�c�}��͋4�c13Y��s��ܦ�Y���1:������x�fD1���b_۝"�}G�@��������.*���>�Lf0���9�f�pq�� �1�2�w�o�O<�++%pLL��>�6�}�E\`ϰ�7�_ըIJ�P�D u�KU휜���I�U�4O^�r�']q����϶津m���&��r��lS��Lfe��d�����}|x�q&3#f&L��>�6Χcf3���|�?:���gV����6��9��6,�f3��f!���}�~0�O�2��G��iԹ�уì�:�1.��w����f2y���h��5��u�����f�+�Ld�1;�=�}d�x�&2�VT���ۆ���1�ȓ�<���]�/~��ŚOc1<�^_�ܶ�i�.೉���s�w�<���b�f%��l�g�0f3bc1�|��ޟ�Y�=��f�t�3++&O;�������d�Y���&&~�Ϸ�N�ba�z�5�B��LB�}�>GÕ}2	t�|��[ݜ�c�d��,��2ɉ�����'����La���=��܆���f>d|χ,�d� ]P��Sʉ��$?�L��MZ�v�D.������t�ޖ��
�ܐ!\ы7�>y^�%��P���h�]0�`\eܒ���9�˽��y$���i�!�3��>��߷�N���]?p|֛��sZk�gRtq����ng;�c&L�y|�{m���8|{���������Ȉﳲ���G�2b`�&2���>�6Ν�c+�&3~�}��4��L�_��߷�����f��s�C��{f��Lvh�听UĪ��u�m���WXW������g�-�Ϳ���>�17��~ߌ����f3����;�u����`����Y��,���pV�=�Vf��z<П�>�>��1��Ɍ�~��ۆ���&&_����5�+h旝d�+���x�����n7�U�zȌ��l���2�#͘���{�ۆ�����Ȇ3�_�}͋6���0f3�9�����|���5�7�"x�a���?i֝L�]<:ʓ�3��a��:əf2VV�>�ǅ�d�VJ��ɉ������q��K���|}�#�ϼϑ���h>���ӶLed��!y�6,�pa����yz�us�j��q:0���y��e�_���3_����:�YP��f%�߽��q�d��2&3e���i8�0�2ϙ��{�M�x��i���(�]���'���1�R��ng*f|��즋��8j�q<�0}��ا#�Lf5�3���E�}�g��]V�W['��w��g����~��ng��3��f%�Ϲ�f��1���b|��߾�>|υ}��F���j]�\ܞw.����H�z�2:�����M�Z�{�F��v����7�qm��/-�lזS~c{*�3ۓ����$���>�$��b����\)���Z�1��"$f9�]��v������'	wMx�[jŸg7��}'�t=ֱnݎr�q�5�v}fnj�l��j�����s��sɋbu�>��2�'=i�Z��ey*�<]-��n�=��A�Z��{>���f5q�����m�^���;�q<�-�ڹNC�gk���+#����L�8�;f��@l�WS�z����ۮ�]��nםs���6�#ug���y�s��Y�k��,��]���|��t[(ڴ��m���3��Ϸ����1�,��{��8Ɍ���1�{������,�̎�m+���x��|�A������Lepc1�/�~�śNF�L7���~�fit���u���17��o�y��C�}��[����i�K���g��:�YX`��a���y�f�q�bL�32e=���o�O<�./3�3�TϾo�Npq�Y>p�>�L��|}k��*��/:ɤ�q���sb��1���2ɉ��=�}|�<f9�|�`�3�Do�~�nk��)�_}�'��YY��3�~��6,�%ed��r3�|�����V�~��u�T�����gȏYg̅� �T�����zO�d�e�Ɂ�c~~�śd����������'���<q��������wz��{��.�d����^��lY������y�]\��Z�w�N��o�}��C�c1f!��b_���,������󞅋�a��q�6c����i9f$�q��S��}������d�f2c�����ۆާY0���xzs���jfK��l��Bu�;�Wb�x����v�z� �]�[���/���o��MY�sM�=e`���سl��e��,���Ͽo��<f8$�c%eL{��xI��g��3��u�4�g�_y�6,���Jʆ�����o�x�a��ӕ�F�-˚�Mp�:���1/��}���d̳,�w矓z�뛞��j����ov*2N�ה=n���=�P�.��!_Q�o��8׍�(�|��k�&�֛r�~��s�|�����Y�J�	���1>���o��O#����&3�����u�d��D��s����}��y�:�޷�śOc13Y������f�I�<�Y��5���Y�������￵Q��>g��ϙ�s�%v,�.*私f�tq���c%Oy���'�Y��1�S�}�P�8�S�s����R��<�&�Xn���(�{��<�y�AH~���w��FJ T��y���q��%e��}案fmO�w����{=g�8�f!���o��ߌ<O�2���WZ�\�:0xu�'c���?wA���d̳3,����b�2U��?r���_~��'Ɍ����y��2x�2bc��ʟ�����t;d�Wc1�/�d�"�>��9]E��6���#�X�͵��ٸa�f��Oa6��۴73�6��r�5�s�����p�֭�����'�s���x�fD1���b~�ϴtgY�0f3++��w�f�q�2=2Nf��-3?eG��o�}�޿4;�6|d��1��Ɍ���?jz�d��kǷ/��.�X��d�u���sb������y�Jϧ�?DMg�s�&Í����r��Ԟ3I��Jʙ��~�:ΧF�f!��dO���سHq��C���R�_O@����f�O�0��	�7_4j���[Lٶq'A�b~����Y�L2�d̳y}�{Y�LpLd��g�d*�{�~3]g~���&�#�D���u�L�-tl����:�4�4ivn�/KF�W��/7�־�2��nv ��Y���dTH��n��~  ��~����q�d�fS?���p�;;d�Wc1�?g��سI��L�wܹ�r�8
�5�g��Ȉ��fϾ�'�*�I`f3��d��y����8Ρ��cLf0Ͼ׼�pq��YY0�{������尒�$g����ϼ�#?w�ng*>�����BR��;�&���w?sb�d��Lfd���}�l���f~ڼ��c��O�������������!����w�f!���Cc1f'����"x�a�=�����~~|��w�?�t�On��P�p�8�\FtE��<�\�l�������׳��+���'��b]s��:<gY2e�əf0��{��,�&91���{�~��{�ϼ�J��R�Jz�NF��������p�;;d�W&3y�=�Ř��f&y������ֵh�:�S��M�h a�>d|�ꏊ;�UP��f?O�Ի�����uf3bc1�}�^��I��bLq�əO{��o�N�G�X����=��v��o?�Qus�'��&&����䦍fj��y��N�0��y͊ptɌ̲c0�&'{����'O��<ϙ|ȼ����%�n�c�6�S�������~׼س��f!��f!������~0�'��������p�"O��Yg̅ݟH�ʻ��Lߟ��L�f2VV�s{Y�Lq1�13��߹�'���&&2c�w>�	>������z>Q�2l:����~�ĳS�i{���n.��,�
��"���yQ��{��?����~������5J�HHy�&�Y++����6,������ϲ����֝e5���1:0�߿����x!�1�!��D|�]���'�@܎����ؗ���>�2������4���1���fS����񓬬���������m�d��ߟ7�����~��6|��[�X���L�6㍥�\�9�����a��ִ�9֯�����q�١��M'�0���lS��Led���=����	<f2VT��3=�Ϲ����g&���;�f��}�vVi3�`3�c1=�}�x�3e��/�9�G�xu������͇����y�י���!�͓�Ks}��r/,�&8&2c�c&&O;������d�VJ�2��}�m�d��Rc1�f���|�?E}�g?�B>�>>�������ո:�w�N�����������f3��϶tg�0f3`��a��zs�����eu����Of2VVL�y�~��<,�K��Ɏ!��s��dY����k<�q�0}�"�>�ʐH]|�4��E�q����Ԙ��&&��߷�ȓ�c�Lf&1��g�����:��1��YY��>��i����y�~s/&�'�������~������1�M��-�j�3.�)�gY+*_߻���xβd2�d�,�_}�ǖm�9��_�������l��<>���<O#���8Ɍ��g���p�:vɌ�Lf0�~�{i8��~�����?���o�"�}�j��:p���[�ΝI�ǞT��>���J�J@qy���u�b�� 0�����H�}������ܮ�K�2l	��9�a��u��<�w]�[o�h��:Z\u��07U=Eݶ�Oc8���.z�ۑ�=��Rˋn�Gvӟ\�34e�s��텗�֍茦�#a�n�z�n���<x���t����&����l����aT���N`�u�	�7n���1��C�n9 ���p�9xcOC�:ݭ�۝��걋�;��۵���ۢ-ι����3Gd�-^}q��u��i��~��?ɓZ��֟����S]����?�<f3"�C�Ŀ���Ό�:�Fc1�	��?g���$�f$�횿y|ߙ�1�dٔ�ϻ��d��1��f2c*_���ᷩ�LL/�~��L�JU�:ɦV��A>��#�{��k�ߡA��/�{ڛ�<����x�pI��Jʘg���!�u:���f0�~�{iFc1�������]�Mg�}�z�3e��/�9�G�xu�'\f%�=�ã�u�,�J������yf�1�1�Ld���߻�}�]����'���&&2c0�g�|��m�;d�Wc1����سI��3'�y�0p]\kE^A}dY�duV}8}+����;�*�}'�A��1��K�}��8βVV&3}~�{i'#�Ę3*{�}��������u@�i���>�<���0�؝d��~y�|�h�k5����8�����ا��1�2Ɍ��;��~�_x������T�c�}�I�g̅{>}DX0�c%efD��{͋4�YY+*�{�Ӈ޳�|3qp�K������,�8:�n�>�s����7���nd�-ƺ�Zѹ:6�Ŀ_�� �@&T����[�{�7����݇��u�&Y��e������Y�Lq1�Ld������x��+%Mu�?�]��Y6ʗ��ۆ���&2�	1��C���lY�������>��˭:�kO!�bv0�߿��~3ȇ��c������.�0}���l��K��ɒ�C���2-��Z�'	�k�	���N��w�E~DWb5w�J1�5^���97�f׈�'_{��<� N3����?��u����Lf0��~��i'�0f2fS�����d��1��Y������7͝־K�~�p��:ɉ����Ѧh�*懝d�u���͊r;d�a�Led�������x�q&3�L�������|����=Oц3++1>���b�2VVJʇ#1<�}�:���~���NkS(�P	�gȏX,���n�	�#_�Wfz��e�ɆY�7y��xY�Lr&2c+%L?w�~猞'�����Y�L���>}3��ݏ����3}�>G�G�ǈ�wef��f'���0r:pu�j�8��1?s�~ߌ�����Ŀ��ۆ��4{���߽�f�dLf0����p��N3`8�d�2���~ߌ�O,�K�c&8D��{�ۆމ�LO�����������������Ɨ�Wj�ZJU��q�V.��]��;ڸ對Ҥ[�s?������=u�~�'�������Y�J�e��Y1;߾���u��&3c10�y�܆��J��~�9���1�/��ef�+*�b3�������<f0�s����@��A1�T�ƾ��h��Ԗ;c��^g�T��F���/�
[!A��+%ed���}��<d�<q�Y+0���>}b׼ϑ~#�����;8+��/go��s��G��2!Z�p!��C����f'Xbo��{�:��YP�3�s��:�3�c1��YXw�w��v>�Q&\��0C���6���j�vf%Z��f���F�q3!�e:�z�&皌Iv^�c�|rb�9��G�&���}�mV�>�c�fg��ݱ_�#���bLf2T������'���r�d�T�����oS�������L�JUp����	U!���1��ޣ�vLfd��{�����c�I����K�=��m�N�1��YX~�kݕ�A;Ϸ��߷����1��1��{���x'���x����`����:�1.��vxβVVL�f0�~׻/$���f�o~��|,��!�y�����<Od���&32�����6Ν�c+%epC�}�vVi80�bs�>޵��:oϼ�:�;YmO�:�tƎCf��Jء2�1�uº�E��~~�=�i��� ����'���<C�c0C�c1���{��q��11��?g���f�+*N}o���[�i��ܧ>��w�'YY/�c&8������6�:ɉ�׏._%55�upy�N�\a���vT��a�>�>_8�H�������=���{��I����K�=��m�N�1��YY��>߻+4�YP��f!|����i�u�hʣ���}��ߟ�d�@n��+r��u'G�~����L�1������v^Y�Led�	���������k����}�����q�d�fS>�ng++�&3C�}�vVi80�bi_=�jj��3>|ȳ�ȝ��>k���*u`|���ϙ�3�B��a�gP���a���y�{�4���̏2ϙ��C/����j�m��m������w���{7�.d�?��y~7��{�B���,���ZC��o�M���f��32���T�s1kN&�#D@;��7��z]~�����d����13����6�:ɉ����4n:�sCβi:8×���NGl��2Ɍ��?w����=�̞�����ep��a��ϙ�o�����0�c%ea����,�c1��b�N����"x�a�9����w����ɚV�\�G-֗O�u�z�����g��wB]����v��W�����N�;b����'Ìĺ���u�:əf2fY�=�{��6Ɍ����LL��߾猘F}�E��6�uơA^��A�!O}��l�%e{c1�<�}�ŚN1��>������5�j�:�b{�;��>��O����]�O��>�.F���� �_}��pX�R������l!���ӎ��z3@Wq��'���M{�˗ʎ��N� �v$����b�Y����~��Τ�IXQ�a�{��������o~�a�
��*J����زr2�Q����������;����P�BO�������Uc�����#�@Hx$�eT�4��4`V�*_�������T�o�	>�H�S\ʼ����y�������g�k.��Fk0�<�Xv0��}�èu%��e`�߾��8��=�9TQ��6��G� ����>�5�F�)i��~�`t� �HV�r~��<	v�2�[�ϲ��m�h��{Gd�)m@��`+܎o2�z��Z��pj�n+7{%�,�t`^�K{�[��͕����si���޹�=��p��A�f��N	V@�&�U��t�أ���wH���[�{�3� ��^߶�:���c��~��Iv�ֽ�%����{/
\�2A�~�yv�:����s}��jyݔvT#��:"���}��#!28�]��<����H䖯-ZLɑp���xP9��}�Aރv���y�{�Qa�ظ�9�M�zwT�aǸ�M�f��i�܆�u�2Tf��l#�$����8��_��<�{������%���!v����ݑN�9�i�񓮥,����)�_�ݲ����{M�:��;��_���yZ����z7�h��v��Y�k��c���Ǒ���wqE�#���lI�E��vg���3Kщ�$��Z;o[����3��Łwo�{X~����ǌ�W�v��u�O\�F�\;�}�\@������ ��=��sp��JZ�N�S~�u`g(�_k�ۜ`�-��v\GC]�y��k��߃��ܓ*uzv��g}[H���{���j>�P��>;����!�;��ǯז��6�n��)<S>S��� ��ھP/m�{,��b�	,x�\�}0�Y��v%��<�:���aV	����s/�0��[�X�Mo�;����W7g�����)��9�qx��ƭ~�#�t��{���ԴW��}�
���x�M=7a��������y�w�{��k�Ji��q����LV*�Te�E-�kDH���j�ĴR�PAeE���+EA`�iDE�B*��������+֪V�VT���,
+kV(�A*ĩ-���X���(�b�R*���Q[,�ũZ�1�����,���2���0����ʖ���qʋH�.�,,AQ��i,E-J6��*QA�DkETUk)��YF[jTJ�FQ9�
B�`�b*�ũ[Bł1�V�E���p��t�&2Ѹ�4ʠ�k�-
�VU��EEDF ������"�m�ڊJ���R��b�e�ZVŌ[j�mj"�m�,XȉmX*���mE�(�1Q��ֈ�"�DA��4�b0\aYm���2�J�*0UJ�U�,rˍKF�"�T--JZTR�0�2���Yb�EX�������UUTb�[%A�+1���,X"�<��i�u�c)q�u��A���wg�\Tv4�f��q�v�8���C���ooA7��n|r����5����h{r]l��[�M'�ӽ�m�u��̛n�s�:��Y��]�fŹ�hk��u�<�e�p^'�5�7�֬�6Ru�n����Sq�q�1�nͮN��=��H��lp��T�$xݩغ3��d%c`[���[�V���A�퇗�ݔ(s��Vu퉴p<�Df�u�p���\��km��U�������6�+n���M�k��}��ͣ�����97oNzݭ�닎2�'CX��6(��g���G��;9�7��s��A˹,bm���"Wmv�M���bH,�3�#ƞɋ�uUѰ�x�f��r�+���<�;�ۣ�'#ע;Ѥ��{:ݭ��#;��#s�q��6ҙ;s��:��n���	^���5v�X������y�&7Q��<�pj)����[c�X��[��n�vuv��m��蒣j	�Ӯ��X3�l�z�s�"������	������n��қKI��ݵ� ���@nwT�u�gǃBR��:S���<�]M�Ŧ3��n�y�uF�p������Ǆ�;K�^�3��n���l��'n��t7�ϋ�����kgȞ��N�q�#F^�'g��[�6D�:�ၮ{74a���`�
:�������m�}�f
�1d�۵ScOn�ֳ�g¸�}�OY�衭e��vn7(=�C�3�ͻl����/:N�ny���<(P�&s���ݹ�iz���n�]���q�9K�e���P���n�St���"�^�ɽ���'y����9�4���"��[��чc8:�Mv>���'���u����Q�Q�Q�Ż՗v5�WD�.ju�'L�ۍ5�tl��Q;��F��k�ݩ�<�5ֺ��h��soQ�^����q{=�`��ϐ�5���<�5f�B�ćU���rd�n'sn�/��6�}��:����W����)�dzmj����{�����^�_^|��8�g	�2us��vW���q7h=����E��T�������b�P��t\���B��\cp]n]�y�Lf|�c$u�����Cyȱ�v8���`��)��xy�L�7�;�:͌˛�{m�b=h���1;�WA�s���֗��Z��q�k:�Wv�I�]v_Z�6�]��Sj�.nZz�ù��۝���cI��[e���ǋ����;�9�I�!�TVv�ƴ�.��WK������-ˡ-G4?�'�M��ا�YY*AO��l�N�A%H,7����r0�<��gs�އP3����'���2�Q�?w��l�N�}��m�e���gk^r�
��A!��n*��ž1�x ���
A{�
�>�N�,@�7�����J�P�������>ߜ�Ň�+��;�nM\Y����
��}�`q'D*Aa�����ͲQ��@�����q׽���?H)i������;H6R�3�{�i��5��._*:�֍\��I�Ͻ��o���}�ft
�>��#�}�DvgH�N�0�,�9＆�r0�(�IS߾��O|��~��y�y8��+%eO3odzȲ Q�Z6��mC,�	>�a��߶�)i
Z~���y)
����+:�V�
0|!�m��� D"���{�m �8�����#�Ճg<��:)UA" �D4�\Ӷ���6�ݙ��qWhr)��ۙ���W[������Jh�h����q��¦�}���u �VV�{��3�Ĩ��{�
A`k�_+���wĆ�����6{H6��B���w�y��.eЙQ�����w�6)�d���o��z�����},�~~�F��m$'����?<��p��r����SA
V	�]���ӑu �֊؜��,o��v�����'�����l�I�)T��y���
��RQ=���lY82�X2�7�y��{�'���l���
{��+�l�8�м:�����v$)i��{��)
�[/۽�g>u8�� �@��!eg��l��R
~��lXr0�,����OИ"$x�G��7����Ͽoz��Ĝ�VKX?��휌�%R
������5�`ԅ����`kw�yw��8R�~o��oK3��._*:�֍\��O�}�6)�
�Y`�S����u3�_<����8°���܆�q�IA
���}�6,�ed���eO;��l�����cϷ滜�j}��p�kL�t�1K�x��o/���U�^nYf�.ԯY�t_>����˕.�u��`�翶x����-�{��)���R��}�:�@�ک�3z�����s�O��Q��<������G���6�"�7Ey��
�����:u �S�o|?_/ߺT׳�����ќd�� �S��{��H)i�}����
Al�ꊨϧ����";*|$�>��ߊ2�L�懀bpI���͊q����2T��}�gRu
$��{���us����Qs7�W���'U��;=� ����Ϫ);������S�%3��36�8I9�hf��V%�7�7X���mH�z*����u�� 6]o�|?�T�
������b�R'�<���'D��z����X�B���>6�@�eeLmT�J��d�dxjC��\�yHV�
���C�~��Ԃ���%�}�m�����������=�o����D�
����6T�Þ~ם�7&�	�գ�,8§��~�I�+%��y��8�2~>���~��<@�J�g�w|�XjAH)�|��`t� �B�!|�nx0*}��?sy[�������_�ў�>xZ�e�=]f�E��;��t��H:���7�⟟���'�ݟ-�����|$����eH)�*w�>���'P�J+�����
�}�߯_|���
���������VJ��FR;3z@@��-4�J1BO��|�� Q�<C��
����@{!$��0*S��?}�:�S��B�ϧ�O��Ȁ�G� �}�z;�ˮ�[�!��~}����C�5���~C���V�����%e@�P>ֻ�x���~���Ұ:5 �)i������ �R����᷃�����2�L�懀b������������À}^>�>G�I��϶u'P�*Aaa|��`��$y3������(����V�`���U�8&�mllH�&�a��\NgOp���N��Gx�����|�8w���۫N\���k�;��Bcc��pm~���O���YS}��'D���^_��5�+t/�:5����ᴂ�P=��2B��Fow^�{+�N�0�D_}��'A����ᴂ���wӲ����G)ۿ���g�"���B�Q�b�7!p�U��n�*�2��ݏI�e�:3�����~�˓Z�5��~��S����H,�2�}�Ϸ�pe@�P/��h#�(��5G[��x��A!uy{�����矷��
�?xv��3M��u:��>߻*r VQ�����o��c���Y�H�G��|��y���*K*J�~�~쬜Y(����w矓��������:�w����71˖��\6�X?��퇠� �)h��{����R
>k\}���]d�a���� �@>D-��𔂇"J�C���ݘ�Xs7����ˡ�"�#���� *�����Y��ę�����~�p�'P*T�G�A�@���#���o� �;����=�7��Rȅ�߽�6�R����K�t#�֗�bpI����19�>�>G�Dv��"�G���;z��3s�s��"���aK�~�!�T(W�{�A$�w~ϨV�ʼIL2��43e��k�F��{ܙ�Yy�7�+�5��ۤm)����".�$��㽽���jE������%U�{��N����}�۲�m��q"��k�}S�^%�v�����nM���]Z���z�`�u9+���nv�h�7.8�틴��.�6�U�Z�;)�v��0�=�4�&^����i;iKt(�5�֢�w��qK�/��yn�Ks�L�6��s��۰�����m`��z�u�&{pN���ۻnnPz�.sZڲN��;qd0NC�n������׮�Yw%�D:����i��^.6� ��:��������� �8~�<�"���P	���7Q$��؄�A9��TA���*��Q��|��c�0��C(��u���:�C�׼nm�}�=$x�O�c�R	$�Α^9ٸ��hp�U	U���I�5(*���)��͚�.�P<N��ԮI�e�R�O3sm[�8�ѧIY�.���$w�����PL���	���A ��v
���S֭�����tΒ	C��%�[�������틣Nz6.�V߁<�4� �j���|2��v1��ל�g!iIa#-��M���tp�\t�@�͎{��6��Α:���PL��J��fA ��Κ�|r�AQe���S��Uh���2'w��Q|%r)z`� ��C���Z��p:�:�ۓn�ʃ�s	#��@�X!�1K|�}���ĝ�
�8u�X2���V��(��Sr���5�f�'���7T��	��ﯨP$�D���p�q1�'#-��ez!�A@�OUH#.�'��F����eMge��f��H9w�$.�Ι���P�݋�j\7ae�GO�	P$�쪣�I9w� �H���*�xu�3�<H/kj��
8pSe��b$3+bI ���3�jl昨���O9��Q˽�$�ˎ"�_�}'���������^��hy�����s�n3�v��N_I^|�k]ZF�8pD�=���JI�#��9�ݿ���6�"Iq_!Q^��&���s�Tu���n3J	� ��b	S��ԀH9G[ܝ�E]=iK���Q �@=w�%���s��U�A=<��޾�*� ���|�����痿���g���Gtv��Ut�g[x�[2�4�F@�9��7�"��P�|����A͵��W����j��
�5��!����]��q�:7*��2Z�'Y�s�� Y]�,W���mbϼ��v)��ќ�f��X�������|�H���"�9��$��|�I��㇢�(e�N(h$�;��x���$	qv��g�M;�͵Z1��at�ӣ<I��� ���/O�gg_�ʠ��ɉfY�9t�!?�D�qq�e����9O`՝[��QͶ��=���~��tpSe��b;�wV��m^)�H9�}4�_Q����q �M�RqZf��Đ)r;Q���i���9S��l-}��I�w�|I �m� ����Ū��V�;����s-�&ى������M�}�s�q��v���3o�Q���H�8���'k'����;�x�{��F) �{���e�G'���I��]`�L���?r���y������_rL<ow�j��al�X�tHf���Ò|��q��$:Z{��~�_��u��I����;w���y�������S]˿��۪��R��� �mI$�޽�Q˾�񧱇���o+�"f��;�}z�K�R�[�`�t���m݈��ompؒ�+L|�j&=��C�'?A K��� ���z�$��}f��mdvގ�q�<��͌�T���7t���ك.OH�
��ϳ���ݚs*�O�$�y���� �~\����=Q��[�ڀ˄Ѓ�x��mQ$��ȟx��;�k��R	��u���}NO������i̶WTn/��o�6��v��<H���D�M�U|oI�=��$��U
#/��) �"HהlܒNZ�@_�F��c��$��@�|�N�0Β��X�&��=L��\g�j�����3f�z��.�sa�J�_޷��pv�FԺ�1Q�.V]쒌l]��W��wY�x��ù�H.p��o�_<JG\��q�c�<���Z�\O=�,N8m�'��k�t �F�����B�c���!�^��-�cgC�M��V�9�/i䴆�P��;��s�qy�X�'i�������ǡ�>���]S�����y�Ϋcms�*�u]��M����0m*Z�6�ݎ�۝4Gf*����$䇰lN8q�9��� �r�ۯV��y�X�֮JX�ʻ�2����*�쬧ƛ��$*,/~��"a8�ǝNW��{�@�_)f�i�v�qF�{*��&��i3�+Q��*0�e�����Wm���;wR0�]�H'ċ�|����g9��޽���jI�%�D"~տZ�s���x`�U������^9w�$���|����[j.f#Tc{�.4N��ɛ�"|I�s�$�H�w�H'3s�VnwT�U�WlI'�F�Bb	R#^ڒH���sZӻ�W������O�r�RI>3s�+Fwvq��%I�f!a�!s�t�-���J6�װtttu��=�e۝�|����
]W4����f���l|��뵈��{�o��Ǻ���i6��g�yĠ�@!���㮧�����f�Y��K�"t-�;���K�w�֢��^�%A;5��#̎�����s4DE�!u�ײk�sн�Z�&��fÁ��ϰb���w� �v}T3j��E���&��N&��l��f���5��6�	��ͪ �Sj�NF�ɽ�q|N��S�I'3s�Q�&!4�,G�G�#�\CU5�qf�w�j�A9��5�A7yӼ��\i�JM�Fi_6]dlJ����4�f��>#n�D�6�\�ɶN��R	 ��ٵ@�A����o6�e,�G��~;�'��	�n��-C���p��պ��˂�>�x
N�.߿�?���T�nձ��jԐA���	� ��D�[�.���v��M���m�}��ဉ̸D+�C���]���*�z���|M��W�w}	_h�8z�g���!q5�+�B"P���&���gU&�Yur_�w}���]��Ȟ�M=���{���`K���ܐ4.�� ^4�����PdLۻ�w���r�９���W����;��*�Բ��}��l�ەR]�1�S�K�t�X��)w����MÖ�Q�lK�(Mz���v,��c=�h�y���q{�Kd��m�-�;�!�[�*�ཤ�m�����!n̫Tf����ڝ�B~83<�o;.w�R�-����� ���ӞՍ�R�p��WG�.߸��ԦY�/>v��6��#/���G�*���5�ݻ}�袧�0�����{E���[�>�ך�Y�6|-�s��kX����p v��^�L���=l��9p��N꽨3;����Niy�p�t��{���"9q����+�\�W{�ټ�ږ�n�u�����+`�LE���N�&��4��p�z�&���&�^�i�C���i&�q�TF�.P}�D�-=���	����y��;����7/���-l�p|P������Iw���fX6m:O;u�邫.*��� z���Lr/Mo�S��l��\�bl�w�fX��;
��TZ��G�$o1����l~HOg�;���.�C�4��#��$c�vN��1��d�=���/���i��� ϻ�\J��i������V���p�i��S#�}�������nP�87�L�<�ȵy�	��^)�Uι��NP�1�m�̓O4�٠$Z,�
ќ֕��{R?bv�'�x37wWiKlĨ��FN8���UQb"�#(�إ"�X�A%J�t�b����A�Z�e(���][]YP�b�1�������GHQX ��UKB��m+X�E��Z�-UAUEAE�(�F*��Q�e5�X�0DG��E`ŀ�0��EVi,D���TDb3+�`���MAQ�U�QE�����L�Eiӂ(��b"�ADb"��*̴b��5k`��H�":IDX)��$PQ��e"*""�
��*��������1KfaTE��� �Қ�
�.��Qc,FEF.�G	���D�X���*����mUF*�"+"�P��
����G��T�b��EX�?k<��(�vo�����I����F&��d�K���غg��o"�o���I;w����}�p�[jL<����{���e�(I��y�H#rvd�\��:ᗶΛ�������n�`H'5�)=..���Ł~#�(�wW�Ż��Xո�6㫬óHUvN�=�;mۉ�����O������s���#<���ۼ� �}���u%ۖ2�����������o$k0�D& �"9֩m�����0�-��@��z�A �g>� ���f��HYݵ����/k�m �(�0�7� ���$�H�pF�di7i_nA ��@�׶;�$�ͩa� �(Q��'�Օΐ�A��� �;rfI �ט��Fgg����.f����bMo]GL�WԮZ/'���MQ���h዁�1�)��ټ��
����1N+&/:���[;t��������� �H�z��jo�W�A� �!CJ�����Mng�)��Ō�Ih65��ؐI;��I���Tʶ���ԡ�˨H@%�C�l��i�B�;�3�L�r���7U�.�3����g$�#	��y�qӓ�� �嘤�gv�����G
��)͹��؄�ӹ��5�6���Aܬ�Lnœ5x �I��H$�s;��@����T^��{dhp�D(	J��T�H$�v�z�� Ȱ⨵D-���Gs�BI���ڣ�֎��P!�B*cd���G6���U�|	$]��@�7|�M#��;��,�*�R�RN\�JÄ#�7'�_]UA�w�#k��N�ò	�ա>$�ݪj�T���!�ݟ��mlE�����:_���u�`����k����G����|��Op,�B�ׂ��X��-���_�%~�dLIEH��RC���E��q��� 9���k�D�r��'�.�]�Wofq��9�s�`�6h \�ɓv6(C�z�����rK&�/�z9ʚ\j�vc��.�b�5��!iB�M�5��^C&�`m̍�&˧\t�mt���[wi�`�O�ny�5��ə���M��]��.�Uv��[g�<ln�S�;u֊�Uî�3̓ma3X{�9��������4x�������|�� �QP���[�RO�5��TI���98	�ήY�5C{�,�ݵ�.^I(B0�,G�D��'�>=�v٭ۉ���G(Ť�@'w�j�E��s� p�����fV�@�ġĒ;���wX	�w�����]i;����ݵ^>�3�S�Ǫ$��%s-�=��eW���ji ө��	�w�I"��,�K�>|Y;�r�kě���De��ȶA�PҁAٰ ������`5�^�]��{7B���w�H'¹�))�C`���̡���Hn"N�� Xw3dv��'+3��;Ok�N^��r=#��������9�����8yuB��O��b���C'�ʲ��K��7� �d�������AL�sC-�! Ս�W��bL�9���)ߥb�x��l�og�g�w����������!�BWC��s���>6���sN\�d��=K��2;��1�H$r��> �?�H$�IԹ��ۢ��EFL��'\��\��|	6�%㻞�����rO�j�R	���L0�j%$�ݧ;���˘r�N����x����Gs�R>$���N���[���ˮ\�v4�p�D(	Jz�U�O��n�gni#r"���E=�;RĒ��^�s7�������_�~�ʜ������\-<�ƽ��7�z�\��<�������|��/�B]��b�} ��اĂA#3{j�Ȉ�F�of,��e�'Ċ���}0R��A,�� D�}uB�1W���&��:3��H�w�A$���@��2����{5�f���[L�2aˊ���&��hQ9�s�z�5ag����F���q��=�b���cX1T�
55~7|��/;=���E��^Y]f(�5s)+�cɷ�$>�اĒg�m
!�D���	&y�O���\�ف=��]�'�����|Ewn�x�}j�e�Ȝ��	��X���E(c5a�#�^��6>�%�ս5Ag^�9Uc�I}�B���9͌��������o�kl�ܞ&�{e�nˋ&T���Y��B����y� �Z�����b��[.��n|I �v�
$�F+�~؛�k��)Y�M?��wm[��C�D̊$��TY���]PG�.9K���^�O���ݡ^8n�� ��S84���5����\2��
	e' �d�ۺ���	Q�κ�n�����G�7ݻT��w�|J��M� �P�Xj���(�P/���j�����Fl�\+���_��]��o��x��t��X\��B�qI������6��_`sx���n�Z��ۅqw3u���ǰOs�u<������שO�QPR�[1�i��"�׎AUÙS��"���M�	y�TI�w�@$��r	ک�]P����YcV���S��Ȁ$�$�mn0���ub���q��n���&�G~|�F��j�1��TI:n�D|h���,=�	������?o�)�5�j�p���d����,��T��u�I�8���$��_9$�녷���Hبs�RG:V64*��@�D���0x;s3@�	g��]�	���R���f1L���%6�=��P��;�֮��gg&	 �Y|�Nf��4&uĳ<����0̬B� �h+B�o�� ���P�;�F��sZ*K�U[����$�3;��P��u�n�Am�>��G�FC��E��\����{� ���t�Kc	��k�\�{g��O�i�^J00���T-��֭�hXam~�������n�����#c��vNٰ򅶬]�ap&z6����ls)ˮ�I�iCz�Ku؈�_G\�:����<(O3�-��Ϯ٬-u���)S���u��z�/huu�r�84����X-��/sN���*)wb\N��u�^Om/-�7�Ϋ�A�A+v�x�$!�,�y�eG�����۱�s��z�N���Z+���ϝ����3�4p����(�cκ���G��xx�ve�����ł=y����vD|h��A${3�hTme��;nz��|�x�uIߵa	��1��TAB��WE">�1�^�Iŗ�I$��@�v�ܘ�T�e���Ip�A)��vI �v��kq����{mu�	�w�A$����T�D�S$�=M�Uҽ���ҩMA۷$�I��T#�6ox�r�}Q`�Y8��� �f!2JE�$�^�Ƞp����y�;�Į��^8v-� ����x��'ce�3�J�/�������Z���/8.����΀��6��.ҹ����ng��a���iC0b�ڮ��$�ks:�p��l�ڱ���]:ĒogUK����
~�����KO�w���&����.��(�frz�^+��޲֓��|Ӌ���x��00��m������;��mM�8��pIy���I�{ɜ�z|F���^'���ωi:��d���^Ʒ�o��`B��Y*��f��$�ɂ	����h�+fr��$n�UN+�rO���	�A*}�ݜ�wQy,r��n>=�[T|I#س:)6�XvtQ���������W]�j���e��A�6`PE�_��t��:4�z��r�B� �	���'�����H�Oۚ���n*�����@kRH���V�7'�S�*�&x�Ƥ�n�76q8R/pf!0BE�$��]�8�� ��gB����N�2Zdfe�m�3:)|�u��	��#*�����*g!���b/ft�'���$���>$���"f
����%�R(�a�X�8rx��$W+�$�|n�2;�a�q^t�U��I��.+�1xp���[Q��jM�������B*ٔ��T�뭼3��ݘ8��~j2W� ����w�S��4TOT���2>�)����Wz�㜳�MǺ�#�9%����������z,���O���	9��y��u9Rtp<o��s�'
CpQ��dN���nL�ժ�"#�3���m� �\i	9��B�������엕%����1������чv�lt��[������`���zノ�r&�tߟߧ��r�1�u߼��=�o���I9��C�Ƅ𕳻xNE����3�|�f!0BE�$����t(������Gnx6���>$��q�|O�9��B�"�q�l��"͌�w�|�W�	��#+*�� ���uQ��Q�X�MfX����'= �\i�H��ڣ1q(�ц�b<���h�*�9�a'���$I��ڢA#-�+��Wن1�+o���'1M���t�;�`.]�ޅ�4��uY�;<����g��L�}��}&�l(͑ߤ�{1[�WnZJ���O��g��M���
dP���>���7y"��xg��f��$Mfv�	�w�K[��q�9�ݾG ~A��9trs��na��;�:B�c��&�<�x�K͋����Ϝ1�V��[qfA>'ǳ�f��8���������q�gĂA��ٞ�C�l5��	��m��pȌ�y�Wx���H��ڢI���<o,Jz���z$+��8�7��$\I�j�Dr���H;���j)��`I��ڠ|N[�R	1��1,t���"�/�=]�wW�z� 	vMPI���)�$��q��:jsj�އ�n�v���J(���X�8�����Rw�x��_���ةTM�M��#<Rm��'<}�Ζ�ʃ��ޢ����|�����r
F8qR�י��,:��p��k!�t�)n��ו{�7�k��	�x���9�؎�hBjSr��q3��k�4�x��g���f�Տ䇶t���YW�6T�xyȞ['>è�_r�<ǉ`��g:�*�4���8����n��%�/��!8��]�S���%͏�C˞# F��f��|;�����w�x�=��YtٓO�&_ y�Ɗ�䧻8$����le#D���kQ�8�o���B�u��קE�g�O`�>�����z4��<�V�"D�W7�n����<I����'�.��dD�2e  }�4t0`��"��-�n��� 9Ht��g�Z�l�]�*��k�!2�v����-(�چ���M$?!ϱ/<���{O8i^眾���A�+�?U�<~&\���;�5�@�澼m��W2y'㭻�F���BHFSä���%����rӉv�aQ�u����苝Q��x?M�%f�7N_�g��QNx��o��W��� �p��d�-1iκ�Fo[ �]��l$�F�{7�퇶 �����W+�W��x�sK�K||���]T��W �S����-����E���d��'�6� �o�[ 3�4��^�e�[�#�cJ�)�vaطGKm�;��F�q{��_2?���&c�)�%y�2�g�˖p_��V-�Kοns!�=�8)�TwA���;�9�=��s-��"�" ��UEU�����e�������WAX�X�(���)�2"�Dbł�QF0UV#��"�EV(�Ҥ��$k(�`���1�V*�U��U
�c"e)QU���b*�d���E�"c֢�X*
���ł�"�Uq���EQ2�"�U��TQ�1X�1������Q�kTUKjZTAb�`�"��eEEeaTDc����Q�JEQ�c���,��E��ت��,b�����(1EH*Ȍb�icH�1�(*��2*+"�* �UU�*`��cX��*6�UQ����Qb�,�(�"1�*�(1\���E��e�k��=�.��M�\���筊�{&�=$�!����b-���5�zVxҜ���۱gqq�˶n��Q� �����^��/v�C�n�hy���pS�jk��n^��V紺3�ܕ�̋]l�Ӟ �{Yʞ�?⾾����y|`��!����nx����>���n ;q�4�g�1/\.�����Y�x�ۋ�pv=;��D�"G-��(�y�6M\��hnp7l�L���8��OZ�8b��e�#���rێt��):�����]�1����{r{-�Qv^2�;\��g������Q��(I��0g�A��۞�	�Qـݶݶ�����Zg�.v�n�oZŽ�1q�d�cWlXm�wn�1����<�n��s��Ѷ;�#��wb0��q۔�d���#��}}V�s9�v�rS2��v�q�8�\G1��ol ���D�7	���[�v={c�{nΰT箺��vx]�Z��듴�7>S�#Q�Z��g����s���/[��I۷7�(�F�ؕ�=C�n+�l[v����R<3���Gm�v�=��Ss�l]�ȕŞ������c�3=Y��l탣X��];ۦd9�1[eN;;�l�1��u�l�v���Y��$5���$�����z|���g��u�����+��׷_<#�[��s�uq�/�W��N�uQ�GH�bǫ���p�>��;n�<�ܨ��:�Hs�6{p<�i6]�x�s.�<=�ۙɝ���7m۴rn=���LY��JݣXŌ3Y����\*�[v�{(��0ʽ�+�܁Ī`ǭ��ؙ5��r'��v��»��1�u�>�fѡ�>
�퍼9�,���;:�rG[�:w���v�̾D3�vn�nי���,��nxs���3�k�ǭ�.�WV%onk�y]`]�մ�HT��=�;]����{s����uh�sַmU6��8�Y�h[�NI�]u��s�n���Q�N����t��u���a��z{]���;tj�354�C	58����}�����0V7w�7q�����v��n����	���I�v�&�k��-]k��喭7(f��#�������z���/�m�vN����ˬ���iO=�y�	�պ�m�@�x�u�^{4�bQ�bksυ����Δ�n�u�my#g�q<�S�kr�dw7n3xݳľL�蓵�z0v�svݳ;��K��N�*n�D���u�9��ocI���)0q���j8喫s�����vᵽ��Z��������e����	���nu
$���$?Z��Ě��U����H�w�Iw(7
CpQ��{jI�P�wePQ�����T����H�w�Iг-Y3��y&��(��T5��P �L���p��3�A�W�I�$ڊ�VQɫ�W�4H7k<Wͷ}�Y�K��	�)��'�:����r��d�嚄�:�b�H��ٺ�#�2��>>�sJJ�8,Da�P�M����EonЩFlE��tFj^r�I�Y�I'3�hT�$�Ж��������ߙ���(=u�y�g5d���i���j�J�x+u����z/��>|<C�ۉ����Mr�S�	#3{j����|ڭ&����S��ut�H��7��Q�s�Mof1���'g��];������)����fsl8�۴(��=�%k���[넷�㓶p껠�9a�����4A�j(k��12&����AD�� �KQ? ���帧������J����9�Of7L���z�I$I�"	Rs�R	$����>'���dՑ[��VR�c�S�I���]��4�d�jHr�Ӊ7ǲ�	�V��o�(�$Iw{f�$]��}8^oFJ��Nnowqg<͝��h�)sB���y�"�����3V뭪�UT	�w�I�������ܐ����kܝ� c��$�6�{\z���I�s&�Ƶ��Yc &��`�S������ ���oqH$�wn׽G��n�򓕱�ig^���8�	����fre$X��n	
��=,�n{:��ʉ�9ϖj�x����^$�|��7^vO��_�!GQͣ=}# �e��.�}:	;j�C��Ee�q���xm�+!�	)4����F�'�xL��s��P^�b4ٺ����BTl�䲥 g���B����ߋ�;��x�Ǫ+}���_M��mz�v�� �ݠ�("H���Jz/KsQ�O���	����(|6��H&��*;4�V	��몢+v�M��A؁U��m�$����w��-��X�����@�v��ZM����W�S��c��N�C�!��a;[c��p�c�Kј;v��\��띫n�����{�>��ɸ��' �F'u�A ���Ms�S�V��݂'�uGX39u8��e<ǧ�&%�n�
�M�Y���M���V����[��D�n���E-�r>:;��8���9Fv�ZE�i�P���|O��َI'��t�D�ܿn�Gq$�m�� G��N�6�n �T�޾&��`�Uj4wq �U2 ��� �|s7�f�Kץ���sJ�YF�ʗx7�{շ2k�s]1�戈�&\���@��M���Ԝ�b���e���2~����C섚��87��.�~�w3�R�wb��_��yj|I8�1ρ>#3�hV@WW��=�gR"7R,3	�*
�xLۡl/NS�{l���a�<�@�<!�������L���	����7��ĀO���ڣ=p�+X�1)V,$���� �p�1	g�:㮽^�L��*Z��ω �k��I����B���	q�f, ˫&ÀB�*�����+{v�	 �ɑ��M\�޹C�َH'3{j��*e�ц�q�f(��*`2��A��$H��ڠI"��*ںU[��G�N��AU�I7񾾐�Q,���^1ݝT|H;j�C��1��gn�='T�1$��۵@�E۾S�K�ax$u�7�s�j�K�s�������2͙����⼤,�I����K��a���jI��;-��6)'�Í:1v�t������ʚ�6y-��N���۞��X}��ZyQ�\�շC�x���ϱ�n\�
�'k.����q�n�n��ظ��Q��뗨-�Ή̮���طPl2'7n��nz�$�Y��ã�/eݻ���:M���*�9��{sh0X�{N��B���p�\�ԽlvT�7=ؑ��:^;v�����,�3�'o>���)���"ݟc�起\��#�v�t���_v��;�t�$ϳ��A$9�MDKg�={�~�vׅA�w�M�o8)F�*�F�$m��]�sه��5
U����4�����s^�������ݑ^7j�H$�q��e�s]��Ċ� �p�$1a"d㍺��A�W�$�8���㹝��6�#8��3���Ĉ�Sv���n�Ȕ�[�8�ޡD�O���O��-�u���%2bI4�c&!��q����)�>$=���q9��b��7'���z��I���Ɔ������s¸fUՖSKMf	�]�u��/m��҇���i�B�j3c.����X^�a���(���y 2E�r�Jf�lE�@��mz����$�[�jp�){��� I�������}uF.=\��q�V�o;�]���l��3�#yI�7��X3��.�گu�VB��L���6�3v�R��D��	�ӿQ���T�<M/��$�c!�@��ɞ��1]�����(���T\-�~�w�A ���3;gF���H9j�I$�]|�ċ� �p�$1 �d����r��go,s�MHg��l��I>9���ƍ�&�O�!�) �w�RpB"0�W�c<H5��U'�{Kw�|����>$�s;��z֫g�{c�}փbN��a��íh�s9�.�M�ƣ�U��h!������!LD"&Zd�q[P�n�n9}�ݵ@�^8�v�R��ҢI�]�A>���)�\AP���mwo���)J��[*!g��8������ڠA�4�mt��Yڷǎe�0\8(�T�Y�����|H�kfz����d�k�[�ˠ�N��w+r���w����~^|�r����#�#�O���^�&1�;�0�0�\4��� ��ݳB+��2чy�`Uo�`�x�p��r�T��	����v����; �Cn�r�Os�m�l��Q3㏦���W�m��ƅ�m�I
�J�7}�B��;n�H<�o��U�Loн�I����m�����;u��^6��ܚ�*6��m���ng�����ێ��1���x�k{v�� �� �z���;�e&�m>�ݫU몀�q"e�AI=�]P�>�SϤ�~�p�H �v�
��f	�ّY�L�/nq=&�s�$��H9��u���^K��͞�W���Ok��	�7j�	���+;m�IM#)O����$ܞ�� ��ު z��O��{��a>�uh"#�#�J���zѳ��4��1�(���F��>sn�P�2vّ�we;�;���ʏXT�1�5�,\�����_�8�&S�r�Ӊ7I?Y�)9븍���%�}�m5�¤���7�u�+��y��[v���]v�V�,��ȭZq��8���¾��DL�ڟDLCn�2��>�̵m�֯�2H&��)��Fj�پ뿚̌�RU��B̉�)�WF?&|z'Y�X6��=��S^'Ď�|��U��I3�T
&;ok:��T��$��N ���b��I5V����B%�<6r1f%�X�v��*��#.tBi5\$a��3��#Fj��dN��~#*�L�	9��ePsn�g�O��s�I�6�8C���D��˞j�O7ݷ��;��[��Hv�P�F�G�o;��OfgWUA��$�V%�s��
j㦙�[������S��,h�b`�/:���&Ʒnv��y��,-��k!>���}�� ؝�����xۉn��ѧ���Y2�m� ��2g;,p�x�=��u0dT��u�����:WW�I�e�"��^q����丱��u��$�%�v�����5�	�]���c��n�<dQS�OA�[rk.z�\��g�O����Y-��mN�.�vk��c��pl9Yyu��.=�N��9�<$s��V+��	��:;O�';C�tz�T�k����<z���88��!P�t����rb�yw��b܆I�9<��$�M�v���û�Dl��)6����M�ئ� r������:�Q#���
V�kTm�	7<��$�y��@�3���l�vN^8RTV2���L1Y{D�N�n�E���UF*'s�/T�ӏL�A&�m]ת@�Q"e�AI��p�U��Rqzc-�N�3�|H'7{j�H&v3�)>��e6�nyӟz�Iˉ.�;]�TI3��\og)���u$���2$Vn�xP$��|�����{sj�u�����#�B���f'��˝��NcMkn�p<:�wJ4I$A!)���S26���U|	��gmQ$��|���I3�v�eG)���۸��� L��C�V��7)Cs��f=ވE��\Q*.f}�*��U|�dc�/4��1����,�ݴ>��'t�vy�� �����I�@��(���3mD��F�;xxA����xN��$����!��QR}v�i#	�`DL��:���꾐�$)��,Z�A�	���ڠA"u�)��,��e
aM��Ο<�&G^�E�5�SS^ ��x��T��CyU��빐F�@�ܭ���)f�ëNz��~ 6g�>6
��_^]�@���mUA>�w�A��)Z��O�U��!\�����뉷;E�7 n�M���Rfלd�d���n���v-?w٢I��F	9{$�+�gĚ�܁X��R�Ԩ�����x�ƏN����h�+�M��k�V�6$u �\UQ$�+�$�@�{�|I����M�Wy\^�:%@-��U��r�����O� H��]H�4��;jkf��X�@�*g[ݻ����{g�b�{7�<<�n#Cj�ڮПggP$�GB�j���7q�$�;����<^���lfO5Ԡ����y����P��c3�A�\^��\��Q�	�xr�`-�2�?y�v�y.ҥs��o+��7����bG�]ͯ�i���pcsF7��U�a*��؋�8ϧk��HX}�x3k�.vo�F����o}�w���'����K8�x�}���Nۻ�����b.�־�P�C���'ݍj��:��pD�茗;�Uf������2`Q����"�wIa��{/*��g����o�r�2��ټ���:��k��緒������z�[Ҿ����{o��瓅>��V������"�����q�׻�����y��nl�)��j�����w�wx�� �5�=U�f��[�k�u�"L���{��^�C��t��Y<�28r�N��K���2�"�ծS'�+�hY���^K���=~�N׈=	|��븴-�⻩����M��G	˸�8��9�d��/�Xqj��o�2nH�����QWQ��aM����_7�Ѓgkj����@�����#٨8���Z�M�����ި<����^{6��a�=���J��O�v�J��C���ȶ�>��c��������[����r^֟r�Ҙ�E�=v������:/(3ݓ/d���8aC��42q��)g�������3yν�ߜE UĔdV*����Tb�e���U�"��
�TDQVU��-��F""�F(�E�DE`��(+��X�TU�"�E��U\��2T�DX�Q���A�1��(�V�m�YDF)1�TQUTb��,V(�U`��)��j,EA����,SI(�"+�,J���������s%b���eh�Z�e�b�2��9h�1���J�bő����UX�F((,F�TA�AQrʊ��Z��X*��"3V�#����T"���j�QV�F�+*
DTUX�WEP���i���A*�EX���PUƢ1TE���������Dc�**��T@�
��PDTb��N���W�s�ݧ9qM�E'� �nT���=x+�&ژ�v	�S�A �U��s;�pq�Ra��`�a�xsL�Ո�Ė[��3��$[۵�Vȷư�H�GS�RO��]�I>9��^�j�f��5��:�*x�qm�	{ �q�IM����oM{Y��O��R!МB�oݺ���O|V�P�Tj��$���@��Q���m�7�1j�����mx�د�o��_)  �Q"&$Ux��uQ-�A4f�,1ĵ]��H�׬H$��@���ONP��Z�"!71 �2m�&��{�����v�	�u�P�h'���� �Nf����� ��N���:&��ѤLJ�&Af�ω�$��{j� ��|��<����a���Ё}dK{�m\n��۷`�R*��
����+w-�]צj�ө�ޓ���:�=cN�s�dgG�d�H�p����"
&A�Tr��Q��.�D�6^�����@�������K�wS#�&\D8�rl���9�.��DgJ�)�/hh�@A����?_?���DD���7�Ax�v��$��%�ޱqۯu���@'ă���Ffꉈ�"~�AI��u(i=~�D�*9rI$�w�j�9n�I ��z�iA�3�]G��mE��L@��Q"&%]���Ux���%�I�uX��_t1~"�wj�m{#8T���"s#!��z�:Af�'#� ���'mީ� �R��t5��z1�rݳ��y�]Q�^��J�@��V69N�4��?o`n���&,��5yB�#��)'Ċ[|�s�6�r�Qw��}��HIT��k��ף�5�"C\�
{��!.
!���orG�\�^�!�ڛ���9�n�k����m����g�vY�<� ��L����n۫<\�|ͷ'1�dC>v�MvՓ�m��ڸ��V�;v�Hvv�筻�ܗ�8�[�;Bn��O4��i��G]p^�]���rxzج���es�W���b��
j��;4u���ylp���˥��4q�z���k1��8w&C[�W]/��x�&�n|z��������v�淳�^�;ny�%�ݶ塱���p�u�G#���ϟݾ(hy��m���eH�r��4z��+��ȡ�k�$:�c��gޛ)������4�Ė-���U�<H.�h��˷�ve�o��n��H'Զ��$���p�:�N��}Ff�a�TG�d�;,�M�rO��͞�}�1�yW�	9j�H$G����z!4Zp ��������vt:�$���e�	�w�I���ØxLwln�@ϛ��3EKW6�M�H�D��'nE&	����r{׵J���'��b��I��'�3��U������]��I���Pvg�f�d��ƻ�ϢR�UV��cC]�C��-����*bQ�DJ�0]��i���$	��T
F2�[�OeX�T���E&�lJy�$(S.A��OV|��e�y�;������Cy�G����B�޴�� =�T���rǴt��ܩ�ď��>��?�/ŀ�����X�2��r\c��	�� Z��'ٝ�U�|z��5�����p&xEpPD81\��ω� ��mQ�$�]�	1�ۆ�T�$�����FggW���L6�"���fN��S��$�	,��	$V�uP$��s����y-�|l�*���J�1*�;��Gĝ�y>w/3z�]2���s�6���r3�n����ʌUj:��Taǘ[&g�\x=���:��$t�e��u�I��='�s����#��E]��&	�"�"��>������;=��б*f܀I �fuQ�<�T2bQ�ʵm�4�g69GJu�zi�I����ҮX[��:���V��)��P�Y��&N8��P'm_O���Ω#u�Ly����[XZ٫*��W ���Ǿ`�U��{����+��{�tN���5DQ��m�^[nf"�Dҥq�I��<���ާ�	
z��3O���͡@���'Ӣ.ʀ�"!���N���YY������o��6r�A�[�6�pA�b��s4�Fx�bj�G�;S��� 27�2I�W�K����=`�� z���e< c/�+�ȵꖻ!�d�7�?æ�
;G��:y۳p����޳u[{Uc=�l��Yٱ��_f�a4Zp$a�ߌ�fТO�ڼ�A Ѯ�>*�m���Zf�|n:�v��M��]�	��ȑ����Rm�S����p�+�*l�	n�H��U��
�1���o�����t@eC0(�
�bܳ�N�r�����=���uuv�k�3�|�iY}�I�:����b �D�:㫲��oJ�D��[ 2	'ԫq���om�ܳJ`,���\kEt뎩�QyY���n���J6�n�>��~��~��}�M��^��7�&j�A�����y��D��ˬ��q7�%*��Nc%@��eBݮ/�)���n݌37�'5�qOP�Y�۪�\�A'3�h
�Iz����]�?A�*
�� �K��4��00�]�]:�����;2�~|����N�Y��[ 3��ؐH$���@_�\������T=�|;WW��pD���%U���Z��]�\R��^꾡���� �6�bA �������d�{.~��-&֙K�!71"1G��X$���(���Ss�VgđսH��ݴ�=�!��bQ�ۉI���o:'������ ���9�D�A��&�d�M&�zQ�ܓ
fP@��UG���Ȓ�.���A̞�$�ݴ(H��O,��j��-ٸ2'����k�N�Qw��`<z�,�
L��7O������|\��&	�bD֦\�3&Dd�ݍ�g6�K_�N���:v�M<�i1�wn^�R��6�lج���u�c��!�j�G��{v;%���vv��}����݉�ɝ���vKm'=��g��\���l��F;H�w%9.v+�g�.��6h�����vCF�ۭ�t�����fzzwb%cn�v�-g��+������i�V�J�8�gnp����O�h�G�kkx������զCj�]���0����yu��b���؝�k�� 5Y����`��Q1Z�u��MI2�
s���H�|k{v�DA#o�|��0�Ř�����rMd�I ��ݡDL��7PJr�:I�&�BQ{
9Gi�#�w�ݻ�@v� H$З[ڔZ��{�Ĳ�A>���[%��
���@�v� H$�fʋꨛ���M�vȢF�d��&� ���"�Ret!�s�b�	5�T|I9]�'�U���E���b�'j2��������W�El	�2�"|t���6��	z�A#+#�|O�V�O�S�Y�;~����ˎ���g��ۡ��:B��#ڳr���v+�V4�:��'���󿝡�Q�o�teM|V��I�U�`EMT�ԃݯ���@�}���A"tN�SB�!G+�$�X��Á�1�鳃;Msxޕ� �3�ҝZ=����ko����s��qѬ����Dd��H��s2�D�]h��T�U�����FV��V�	&��-�ݙW=��OULD�@)�p���2�m5w�4�@�u��A6��2�I;]d�|j��I�Ln��-D
p*�v;��z�W�1�f� I��҈$���H$���v72�4<@'��9���#�#���A����>����u[8�v�GAN�G���ؓ��Ϊa�=��������O9���Y;��b����zsm�u+kZ�LlOD��;��������������b)�FWdO� ��Ϊ8 ��围�)����À �c�8�� �0`X.�{�7���-�| �~\��z�@�9��h�ؼ�#'��v�`�QT1W[��� ��3�)���S{��q�{k��o�����E�0���;�)mϹ�49̖#��|��>/C�׹W����}��+/��}��W
�d�2	��f���{�F^]LD�@*F�[�ﵧ.(�y��f1$�y}�@H���w|tڲ����O%�#�7�a��
18E��M�<�w��9��(Y���ےA&��k�'o��/.�`Eԡ�ǹ�ı3 ;t�O/p4�`/q�n�)���!�l��_h��@�fhE�p�*!�V���_mQ�v�0�&	��1RE�/�:�A7y�v�sz"H�D���n6�u��i�tH$�_l���a�	�{C�t�&����'�)!8��t���G�����$ڨ���z8ęUe�\p$�k�v�H��� �'p�6�1q*P����J�Y�R����wͳ�{B�o#��V�X�;bc���7��U�a6�ܩ�'&h^��&6��%�l������Un�)q�c�ݷl�ʹ���Vt��W-����Ó������������0���H6�7?,�9�w5>쮿���Tg|�/�)7O7�������0��0���nn���+���e����x�z^���|�~�|���,B�h�4�O�}B�;x�Q�'w?.�x����+�|��9qL�D2\�����I�\��5��GWm^m�A;{D���>$�d51�Ւ�g�툗�T�"$�Nf�]6��z)7�'�L[ˉZh�Q���I={D�������e�%��Aǈ#S�Q��6�]K��]@��s!O��W�I$��Sj�wxR�~$D\a�D�Pnш�p  �S�RI��B�V�䆍��Q�2�4� �+�>$��]�O�%�v荾'e;���G��Ɏ�W	����,���t�V:x\�զii�L��u�M���s5E���=8u���fw�\v�ai�{������,�;E�.�cGS���<�e}�{Xe{����;���w6>�K=��i�?#��9�v��b�G
�8��^�����=�:��1j��A��������c�7=r����랅Q�A�aR�_�;}X��eGC-ɣ���;��)�F�;��&�~��n�ނ��Ӓ��Ql�0��5�Q-��>��'��e����:��N3|ǐ�3/����_�k�j�/n�y�<*~-F7�L6>�c����=u��-uE��o�Qvo���g>}����º�y��I�k�8��L�+C���PcAUkf�)͜Gd�K�r]F��v�yd��I��Q�$���w�e���ҷn�x'wS绹(][��ވ��|竓)�J��<����/a��!�����gb��}k�p��j�pn��*:1�����t��|��0m�F��É��z����n��O�sޫ�2}@��buǗ��=�ϻ���כ���;�w"��յӽj`]�
���9x��V�7
+�g~�N����Ȼ%�]Jz����{��@���լ
�Ѿg�`?n罸7����Xj֥��ռ�TI3PLUW��juQF7l����_�7��v#��p�I�~rx,v����U�������B��[���;�&\���w'v7D�3_t�cٚB)p����������[�[z2'h�^mP>*
,Qb�j��UV*�m,X�����,`�)Fi���a+hZ�m�(��(��U��
�5R���QcR���X%aF*�QX"�����EҊ��`���M0�Uf�#��
.4�őE�Q�QF8R�#*�X�"1TXkWAkb����Q��8"�\j(�lm+ ��TE�lib�Ъ��1�Z$Z�Z�DYZ1T+X�
�XJ�mEm��H�����CDf�V�"���b�Y)UD�R�b��
	Z���Lbe�T���e�[��i[Md���Ɋ�*��VT6"bJ�ب�E��SHU5K(i��1VF"�4�Yr�b+�-EDUYj�LfeU��X�TKh�**k~�������WI�ȧb��#�n;y}pq+tuN�Lc��q�f�Ľ���.�ͺ�l[�ʓF�:,O�k����n8��OY��S���a�Y5�sV�v�۷q��+�v�u麽�z�x��m��ݹ�ezzIp�◍ع�4����ǌ��B�:���8<�î'�F���9�eg-�G"um��6�{n^��qs����g��
,9�m�'��JV-)�k�ae�N`�>޶��ss�Mmț{�[̮l���v;W���!��t�v2U��Fn�;<6ŷW//1��(�ەp�[b��xs�����������8���%�]��rj0g��/N�v��ez%n�6v�6mi.�p[p'&�\7.ڛ= #���V�ڕf�.��շ�s䍩s�OOgzL���z"{e��\������؅��亻m8�Jv�n5=VS�&:�\(�<�/N�Eh�n�@s�6}�Á㬥�y��x�	�+��u�y�ۅ�ɣt秐'Y�������P�2�Ύ������&�Ѷ�g7k��ع����1wLu��Zz�ג�8ɽm����M�cuQX
-{n�s�gal���Wn����ݓce��1����t��F:<���Ugfw 't�z��ƞ���ptY��:׋��ӳ��a��8�Ms���"p�W�����][��<n���'NmGa���uk�G�����X�6�]�����r�[���܏F{tuҽ�n%�sk2�@�k��aB:�
�nK]6`�zsc�3lOj�Wn���gE��%�rY�̻p8 ��hѫV�.�%r(nMn��{�7@m���k�:Fw�^�N�9���y8Wm���ٹwd��h�ƖH�j)�wO��ri�q�C��)�K��1�k�ݗc�������c�����mX�s磇��·�=������G��Y�;I����8X�JvOG�#LM�WOc#����L^v��R��z8.�Mtv��g�f
�����[�Ybc��IK&3��M�v�&P-7i�u�nP�:��.���N�6����o=�����O93�:�V��n�c�ۣǱs���X��v�9��0�m؀�����k>L`z�&��kcrv��!�Vn�:��v��xܚ�R�������M��:�p�8�n��vg�V#n#��F&ӷ�8NiGy�&���q����6��>z�ݜ��Zn�Y].ܹ�=��ݽ�u{9r�b�^X�a���#���������{"];'~�~��I3J�	�$���=j3*�6#b��w��χC|x�ﰑ��	iՍ����m_^Nw!HT�>$�:���H5��T�>��Q���2v��E
�!�9.�{պ(�A��r���;D �?��W�1��!L5�DIv�����D��}�m<�Z��o3�� N�Fz%�s`�]JG�9��tZ	��d��4O��<�,�պ�|�u=��'m��$����
��k��\���Ib�a4�Ch���]w��9�t�E��E��N�ͮ:0f���n��?_??C|D�����mH$�z�r��I���5����}�I�>�w*�q�B�`��d�79�!<Bܩ݆9D�G6�f͖�r���o	���M{������\HW ��Z��˥]�����c��l�b#;oM�@�+z"�AFɽ�;���^�uz��F �Մ�:z3b��gͥq^��%�0D�[�KS�=�@$�vЪξ�{f'��ͪ��m�x��zg��	�-�(��ݒ@�-�`��{7�� �v�b��M��\8����n}�֭���@��T�"%Ux�*���+�$�"�3{��ι�u<�$�M��O��{�SZA8���wgi�Cvmņ׷m�����ϙ2�Z7$��Ƞ�Q�̷�"R-���V��P>9K�C>'�]oD��;J)�6��P$�=��?�@$�,Ո�����������r��|I#i�)'ě�����OxO�*�rݙw!	���टx�2����DXUEi�*�'L�4���$�X\)Fjޓ�Y�CE�y�|�\:r�����(ϫO&���)v�E0��Wt�q>&��)u�N9á'C��p*���0ꔨ�P(�*�gĒj��@ ���w���ХRl��f��P�2��r�1��>�@;��B���]j�B�\��v�bA$���ҦՑM��i�2��#v�����h������-A�<m�v���e��k=5��-^b�?�?~'��c�����>#����r�:�.ű˳W�8p����M?_t�M�}P�2�(�?	�:�z�Dq�Zz�71:�1�N�tH$���(b�u��u�A�ʲT�D��4v��|I��B�$��e:U���S��f���A��郒�������ЖVX�]�^$���H'�ۛB�o�,R�d�R�U�T�_-q%���7�$�˔�z����p3E���M�d+�i�rn��o��o��l�pb�`���j���7��81�ҳ�t�Ăr'��
�T@�1��^�NZ�Xr�Es��Kc��$W8�s�6Ex��ا�z;t�
�tjd�
+�"�l���V���,]�e�F���[ܽ�5�&j�xhP�2��r�Rn�*�6��fuQ� ��ؤUx�d\��腝O�s�6�Y��j�p��b�3�:��8"��sn� �vl� ������]e����&56�� #"�� �Sb�$��g����B��֝�z$^_l�'�o�O��]��Cd@�0�s�g�`��qY�	��M:�b��w?M2(n�$���
���D6MD�R{ܲE�b�リ��<����N�r�*��:��AR}7�h1WyѾ�2���[=�|�jΙ���ꧼ��}Q����ݻ���&(u{;45��e �'��q���y\�%[��*P�a����Wѓ�.�\�.�{�7q���ƻ[.�'^g)�	�<ڇd�k�wG��Y�-p�q��.��p�R����!Es���tӻCЖm�U�g��8��ə{f��ۍ�o����po=Y�t�'okF�����t�3�ɸ\�[v����h�e8�z�X�ˈS{c�	�e#�.�ۣ�;٤������V�;�������ݎx�wm���uǳ�z�գv�+�Bh듫96���[�������"���{�{-fHd	�{{��(&�Os��~����]���(L�hd9EO���ۚɊ�����w����Io�Ht����L�S���;]�EfZ�y�R-ª.�FʾRH��z*������k�b�A�{�I�'m�Je��A��b�i� �Y�'ŵ�>��EK�RH$��k��%�黯M��ڲT�Dum��d@q	"����پ��E�ˊܻ�$�6_b�H'�/{j�5C$�y]{��ϭ�k���}��N��t�gCGX���A��.�^��(���;��
 �e���nR��[�|I �����F�q���Ԃp�m=�u��u �A�ca{����B��y+��GFB����X�λ��f�YĬ���D�}2w`8��8EDO��3����K}������]�$��p�n �SYlP`�^��flʚ�2>�w��r���Y�iB|M����@\�A!��E3<]J�I>;��^���֒�w<I;OuI �r���G³G�/� �ú�x/�����o}���b*pQ����A�;��T ��إآ:��r�a�[jA>:�"ղIM�`���T	;k�C�R�ݺ�8ܠ	�wJ|A��k�	;o�O��}h�<�O}h�������l3d�^-�Ǜ��V�k�z�_j�vWv�ܜ�d9�M�m���~���w\��ӝRA5��B�'č�ؤ�C�q��9�lv���T��Mv�ר��B��"ԃ���m��U��u.�`�A"�{j� �m��>'Ƭ���s��w��z'��I�e��Tg���Dx�{4f /���?_^�]��8Rk`�B�&�<6ɲ^�';�1ڌͩ[P�~"<k�y5W��=�f78 6a�w�F
���e�&�wdP;K�Se᪛P�2�ȑ�>�ú��1<����ɠA�y�O��}�DK���x�P��?J�c����ڐ@��E�
�|�e+�>:��o@�9�uW��<�$��-� �\�+%�l�� ۄ�:3٘�fݍsp��#��T#]7==��i�Օ�Yz��x��1�x�˪�KrC��>� ���T��v�c�'i�*u^� �@�(���Eq��N�敝���zl�t���ES�R	)�����WI;�~�(��%,Dn��|�i�T��	�%NY��*���'ď\o�o�vwߦ�����d�ʻ{��Q'�%�;B��� ��ڤ�Mgv�b�ᡎb���-;=(B��vv�C͌T���k���۫�s�r޶t*�N��U�Tbu��ި��!ɏ��)�e�C��6�"l��;ƪM�d�C"FFf|�m<�ݨ�١�t1��{�I�[�I�>7��T.f��w�Q^��[�!LĎf��2G�VxG�w��۞z͹+�2gs\����r	�꾿�o����J
	�Y��U����W�O��omP8OcY[�8*�nqH �����
����4ҏ0Aީ�^��^���{(�j�C �z^�H"��hW����aGR�5��(� (���^o��ڴ��fř�(����RO��y�A��m�9�d�2eH�+�;��}�=^dE�� ���٢A#i�,ꄦ�7"̬��s����M���"~�%�*�UwN��Ȓ橻�h]g]��E7Ԥ�I��ڠI�}�g���	��њ$��N��9T��z�Z�:�p0Z��k`Ƀߊ�i��{:M���!ߕ��w�$���.y��'�:�o&�Y�]�Jx�#	|3p�(�E���㎸{_��m��~����7p��s�6���ju�=��ݛnĜJ+��MM�
�i�������w��v� ����1��|'kq��g��b�u��������qo	�=���7*V�<v�z�ݞ{u=������КQã�E����!twZ:���tr9������v�뛍��ۍ�;�#�W�s㮦�ة��n�T��#�ob�;e�%B�v��mv�l��v�,�����w�g��c�_omO�_v�'i�)1q�T|�u��,8ujO��v��87�󆠠��A�;l�0zf�豴�U�}���^$�������c�65{=뎎TH*���h ρ[�uD�v�b�+.���<
}k�/g�v��v�b�3��DJcP�%������������j��P ����A"��)l���L+ӄ�1=֭�^sR�"2�q�Wz�]��.�"�Ɏٟ��ݪ����@���}�Jtc���6)$��2��yc\o;q��vҜˎ���Jó���	��v������v4�-���l��>7J�Y�$�<� ��:NԻ/ܚ��+�]��%խ�&Z)�v�i�],�!y䚥4o~ц�^�n7�G��[��=����figE+����DR�Q��wOpi�\�{؄ټ��j��� �M���I�S�R	7W���B繸�ޣX;sĨs܎"KQ�}5�3�M�1�߉���͕�9��O]�������U��70�.<A�}w7�^d�$P$]i ����M��S�I9�ۉ��O6�lT���R��l��LjB�����H ��mQ��vjޙ�G;�I�W�A>��wmT��bY�JL�6�bq�]N�Z�Sm������n����rN�;F^��q�9%���A�=���Mݝ�m�Fgv��uvn��@Ή� �z��NL���B�

�'g�h��r-n�fe�d$�m=�$�^���XΌ����[��J�X'İ��p���֤H;��TA φk��;�&�*�ڇ�Q%V�$b&���ٖ�vlTl��Rp5ݰ^��4pN��?Q��s}g�{\��=N���+�jc}e�s��i��-?2���o_���`=���쫴�����Z]�e~�x���h.��ekV�M�����&��{P)j���o"͝�2��C�J����V���_����7T����	��#Ox��|q-^�G���q�%�͝����ᛜ㐰i݁�����!�k�p��x�F����{���1{��}}�B��|��2��˳M��m1��]��}��.W%����wD��1E�o��;c��[Y�p���m�-��K=K�<���w�`���}oh��<�i�3h�{��X�#���C��n�q>.��tX�±�I�y]�wplv*�=�{��]�(��r����u���c���Uc���y7y�\���;����wPu��«�胀�gyhN�}�	$�V��:���}��!R��՜�	����Oc�;>Ӑ�/i����#�B��L��[�ns¬1�XF�����3j�cDר�F�I���Q��vB(��:�k�������p������J��O��e�԰���3�g¥[�4�q�a9�}�ֳQ֯:�^�	m��z_Q�6�W��W�\}����1`��]�{��;<}T�
ܣ��F��ū����t7��Fi걿��[�=ρ����}�q�l�+��ʴ�F�֖�cP��W�0OeG�9%��v���-~�<��ӹ�;���w���.*��j��*�2��.R��l�TEuK-�0Q�Ŷ�U+A"�K��X�T`����R����Q�$X�DQ33m���UbZ����X��E�Qb1DEm��2��LaETQU�Z�EA�)R�Z���X�V�33)mFik*KJ�j��(���(�X�Z9lQQE(��ւ�m�k+��1LE��E���PJ�N:n�UTUih�[[X�UA�s0Dkh[���(�(V�()Qj+�T��jժT�F��¦����ZʩK*�U�m��*R�cam,[TF�#iV�Qm�T���F���m��X��ʪ髪TңiDD��%Je��Ym���IR�E��[GYr"6ֱ˂�E1���\R�Z���y�8T�T��N_v�k�x�f&nQ����7:%�1�q��$9/.�ٻH �z����K�\?] 
��/���zZ�q?5e�72��iޘ���J��槲�~��T�݃y��j�$�z��NQ�M�N�D2a.��җ]玝Ӌ�❮tm�=[\kW\t`�-�΍��S��DL�jB�8Y������{���;��FO�U�nŕ(ٞ�j�{��ڰE�rK��%��6;&(��k�]���'���ww"h$�Z�%�d% �lV���W��7������$��*.���]X��<{��6U�{ݱѕ�'p $��mX���T:�5O��&_��d��1�w���q� 9�uՀߏza�@"�w�½���9���o�s�E�x��^Vq�xU����90��Ɇl�f�v{}s�
� ��w�;Sëݛ�p��vI�A> ~�z�mX����*\���*��z;���굎awk����m�d{�� |U�qvJ�<�UK{�}߻��_<u�x��;��%�g����[���������\�\=�~����-�'f���le�}V�x�LP�s�]��^�ha�vK��R+�j܆d$��jn"C��T���$�;$#�e��{٫��}P��7�V1uXKH����K����:B:�J�<5��W��y��z�Ƴ�on�6i�@}���t�;�VK^��~�e
I������J�j��@bۜ�� gv���z��;���w<@(���I�U|�"T�!p��zyX�?v��*'�����`�@Df�:�=s�)����Y�3/���|���Kc��ʱQ2��9��n��/�ե��1�Uǋ���4Z'��)Ԛ���7�����㧵9A����m��뒲�Nm>��F�n퓠j-��I�v�@��2�[f�wmƫ�<G��g{���Qİ���$�%��vW,<�rw.�ֶȕ�:w��ܐ�dm�vn3Ȉe|윺����\�tvdH�����Obڹ�����Yn�<���CWV'm>��<��>���}Fw��:���S$p����v�#�n���;��ݷ:�\���면�i�]�x�;�f9��j��l�q�|��ssmq3�WjƵz$�l�[�ӕ�)���a�W1� >�������_���>s2v�ίG����]�qNԏ^�a	�q?5cl뼫��Xt�����+&J���f���ib2;�/�{������xؤ���%�(��N�Xt����� =�jl@�*3�Z�K�{�6L]z������@$dol]���J���*	��c�"TVh��L�4���`�_��ػ��O���}h]���㣽�j��P��7��(RD��A��E7h<z=�S����mMFʷ\�Iy$目�P�эH�9mo[-j��L��7� V�Đ �a��f�c�$[8S��U�'���^��76�Z���O��&����
�.76-X|����lĶ:}$���}��Z�>=�ݠ�ݱX'��r�9�22\Y1q�CD�[�#H�p!:��B�����ݾ�V�N,���ӌ�U��g=�u�ȓ#:;���_i̍b�*�r�$�˥���I}1%u�S��7����#2:����l[w�c�P��w�;��Wj��^Ǭ$xj�LBi���Ֆ�̹� �N��t�^����N��f��#cwb�`iޘu�*�n���wH_n�f��7��p����\\%cV l^��C� ����w�sj*%���˸��)\��LD������Ɋ� Yy�vS��z}���� Y�@|./�-XZ~w?����o�ߜ9��[��m=��v�Mŷ/�:����a`]������ rB
\��?rs?I2�$K�oJ�����za��_tU���s�����:�lH��8���"�Hw��3d�i�D�h"B�����Y+�[k6������ a�0� .���bu�%r�ʪ�y�K�(��a�a��sÃna� =}� >	�Z�b��{��\wP���/���ĩ����`�����}m�6A�מ�u9���9�-��L�gw�g���k¬dxK���g�  .���%:1�`��q�)PI����3�ȓo����6�n����ة�N��o[;��z2�$E풉��B�GV�݂ 4�m���ݗ�w� +�ڇ@ �z�X�F��;{�wq�w��ύP*u��ٶ�x��n�Te���a��u����k�=�	�2���>w�F9�nZ<��L7�|y�X��티mT뺫U��/��XR�=��>��m�����jl
�����_�=�t� �H���v�틱���엖���\;}��i�D�h"B��~ͻ��~;v*�	���U����V1�j�<��6Js�˙��ɍɈk"5�G���O� V ��b� ��:]j�j�Ε[�ׅC�y�a�K8��Y5׋=��z9��\��5��U�r�W�6�������uZ��x�:u�2/7v0�rIm]URP�8�4AD��VZAf_�`4Θ��{�s���`vߪ� ~7v-X�>�Ψm�
�"�U?��G ��Z��Ia��?jdzv�8{Oiu� 둷Y����������~���]�ۂa�Y���ڰ��6 ��Q�g.FS�USm���ؿ����J���
b&Ivl_L7H9j�~���zoz�����v�7 63�m��n\nq��{���1�?DDa8.�_tU���zb� �+�����^���u�I/+{��^KU�2L��ɶ"T����u���ӷ�j0�@�� >@,��H w}�mWk�Ҵg(�I�6�z�h���&2�`��crb� =}꧲/r��EO���� �3���޻�\Vg�	���|���CT��u��
/���qd��':���˹�/d���'���S�
�Z���J��\Eײ�4^�45���nH&%H���snٲ[���hN��Ҵ.��l����g��.[�E���)Y1�����M���k��ۑ�9ydyv�����=�C�^;`��#av�m�9 L>̻������&����������/r������]Q����<�"�Kٴ;wj����mǛ��\�>�F��h�8�^82GP��<g�h�t�-ۮ�*76&U��	.��/��+A�u��GQ�r��n��K.O�����I�;3�Zp8�e�� ��ي �����
#���U�
�.�2s�v0��P� *=�J&FӈA?B�G���X$�q���e�V�[b3��@"�z���d�_O�.0�je��1����� �uS�>E�m��뼚��3j ��u��
����o�%�-�u�$y�����Dl㰐��LR@؀[~����ol�9�j&ѓ��ː��C���\�b%KAK/���v� �۳Uy���zNU&wGtä ;�ڿ�b��o�.�G�^"����v�,Z���@wmX�;u�u��P:zQ��˼��m���e�s������|چ�p�\����ܘ�=}꿕�� olݠ�8�n��P�m�w���J9���q?5cl�Ub=i�o��)�c8Z�U��1)JN�0��j7���yh��y�\�JJ��f�Q��#�kq�FY����9�A�����c��z&�/�FLp�Y{�v� |�ٻY�j�3�m1;��C�$%��b%��1TO]I&���� >	���n�އ�}�v6��ݱN�<R�2
b	Q%ٱ}1�;�l�u��U���S���`ٱ�P��E.��! ������V!+o�%�-�u���_��10L�(7��q�9f,��]� twlp��h�&Oz�a�'���Cpn��u�����/	��Q�5n��3�m�}du���~~�m1���&�^g]��lA�nm���P���;j���O^z��b=�`��9�R�p�\��1�0� ��iC��}���Y`�cwb� �Kc:��=�u]ד��7#r��Q���ˏ������A�w6|��t�| /-ͮDEx��]u!37Y%�z�q�yurC�}׼��A�x�O�
ѕ
��;��A�J�b)>�f�p��W�O�g�v� ���v3��:a�
=��	����<�y�~���I��o(0���t�m�H�޽Yq���^���͊w���L�B��TIv���ۻ�U�w�'��1}�@*�z�� >�Ψt����+6-�T�U��VS�f��D& �mL����?�$�Ɏg�v�|�gu��.W����˙�Fe����Ϛ_Sv�Epq~��l <g�) >�>�޻���ѥg)��Ǵ�+�!(�q���O���Z/��h-�ݐ�5����l��T:�]�]�Q�/Gvl��7��]ᏼMn!� ����crb����U�a�	:��yw���_�1�@ّ��m� �޻�׆�L|��~j�� 켋��j���O� ��b���:�n�� G�{b~Q]&�ܪO](�]�5XrDUw��6�&�)kQsnl�c�[�B�8^V�R���VE���{�������N~���{��M-x[�s^���e�å�T^Ah����dG������I%�;k�G7˄�[�d��ʇH w~꿕��틱M��e{������������,N�T��Ѯ�m����J�U��l�b���N!������:�����Hؽ�� ��S����Gv��z�w�~�*�<�ϖ��8������笠�����漖���\rWn���.��p�����_z�@�wl]���n{oN������M���8W��Y���'�O����i��z�����Nye냦��}}�M��{b���s�*�s.f���ú�V���;4)JǛ���Iw����B܋2���˵a�.�g(D����VX�۪�RH�W��~�g�8��I�tn�9m-��|�7��|��u-�	!I��B���	!I��	!I`IO��$ I?�	!I�xB���IO�$ I?�H@����$�`$�	'�B���$��IO�H@��B��@�$����$�p$�	'�@�$��$ I?�b��L��;zL�̓� � ���fO� �O�ˀ    �                   =            x  �9	P
=���@ H�T  �Zj�U@iCBTV�(ʍA@�h����C@�J��   �                               @        �@�{С;�49�.��;t��ܵ�[�j�Vm]M�W0�A[��W-\�U)0 j&Mr�˪� 	*BC�   ;�y����m@�7z uU,�yb��#NmUNF媪�W �U��t�R�h���*���U<�$�       P   =L���.!����R�73UT� �U�={�S��d���ڼ�UQۀ �bk��W0��@+o   ZmTS�rj�Om� ��Nm{ Ӌt���b����UJ� j��8��{��yz/
��\� 恶H <  �      H ��!��@wX70��y= v�� �JP�)fvh ��@�b��@ �q�� �v����=�t��AJ iH��©��  	 �4��]��h 
S�� �: ���YJR��R{ ��P)L�4:�y� <��5G6S��@;���c��� 8�  ��@(PW� �       � ���`��2 9� �� ��m���9�8� Gp 8t9W@9p)R�J��  pא=�-tU� ��  2!�;3� ;�  �� 7`9 5F@IRT���   �         G��@ݨk�t�  ݜ �` �r ���.�� 3� ��ju����	�b�   �W���l��w u
=�<�
������l��Ap 3Tڮ�70ӡ��j���7B�����44�* �S�0�)P   �&��P �Ob�Q���  ���b�* �S�D��R����wq�6�h8�U�ks<ؘ�3�Z�Q̫� ��3>�����033`a�f����f��033�p30���S}7�y�6�yʪmY���mYc*b��7P�wiJ&�<d���w^Q��Ƿ��x�Pq�̤�#�X��99k��7�cyie�]�T��W��9��׋�mh�Sxmv��o�gh�ML�EX�Xi�u���2+�T�9��U��j���`�xt滲p	���zq���³���݂�ilUแHJ�#����/Y)�ԫ[t��eܻ̹xd�MI!Wp(��ً�<'u��yM����4���{s�� 6N�Б�Tm�v*j!
H�:��%�7��x��e�CO_�Ap�`!h�t�h��3M}�/�E%Vk]|NH��p%*z�O%�0�ˡ�n@�׈����4v<]�0Nǈ66e�7vcf\��Y�ϻxY���&B�s�t��n�99!��[C���E�+���
fj<{u A�Q�s+pdi��t����
]tD�5&�.ޤbm���Nٺ�RE����&��4� c�����P���R��C�������٧�]]�Xy�,����!�a�NZ����46A�7�P��({�e���X�y�Kӣ��#��1>�u��p���G	�8�����
�q�s�<�[�n�]�w�����Xr��=p9�����ʶ�]	���rv��{99�ʤ��-=l�qt��ո�-�丁��j�O ���u�AW������v���=Ӌ�9�T$�rӷl��i[3J���.��
��;�φ���/*��h�;2� �{�+ػui�f܎φ������w5��K��Nf��0y)�L����a���r�&\�s���XN&-X1�!�+�+�!�up�U�.��w"XI3u�u�y�Q�pR�`!Pk�ӱ:
QI%�s���&-ŬZ�%8uk|���Ѝi;tY
�8<A]\�}(��E:G����8�*���elȸ`Q\��z�sd�А��AC5�[�V-�h��/X�qN�өP��ޗ'�4�n�W[�Ҿ���k�wH���G3]��婉��\*�8v��sW���n3�E�ܒ#�����p�3[-��yC�B��r�gN%�9e,#��6��ƭ�+�,�����:o)ʜc)�c}�H��gxrQMgCh欝y`i�]�5��UR๯�48��5��X4�O���@u�/*4C�(�NO+�^�&oU�_;�������%&
���0Aܚ������X���E�w(>U�.�T]�G$�l���A���*N!+3t9c�K�2Q�U��N�ľw"��[vͧ���mSy��Ů5#wf(��4od�x=�>ܜ�&���Q���gkSA�^���÷�>gaA<�I��8N����U&����0�[}�,R%3V�Δ�.�2��o� �	�k��L��Et���:��݆��M�_σ���O˄eڕ���s��fv�GgU�?�z��!�3�4&�O� �	��F�WL��nK�L�
��x��7SA/���x�ݗ:w8Np$�+�G��`��1��!������ ʱ�yؘ���d+nM3|�4,+���=����5Lɺ/bLl}��՜�KC8�vb F沆u�Z�Θ)��2�MI�=S�ѥ�{fv-�-�@ �u{��JX��-�ۀ��94���Ч���Ѹ;�ȂL�������?m]�dǱv��΃��ꓼ(�B{-sxj� �wU#�qћ��o���cHm�3%�4�#n���)�ֺ�е�L���f=��\{B�^w8V1a�;Bn�\t�jWyTI�ur�wC�"�A���;hg�ݝxj��M�ňVC�aN2�|OoBÅ�ׁ�
	Z3w������ �8����,���4Q,'���b�R��\�/K����0��t*G}�c���Vznq]��xh�L�J��{�,xW^Z�q�F���N�5g 
�8�sYnb��;�U�j��5�9b9�U������b�����V��Ι���0����v�-�vHa�@XO��	�2��ToM`vۥi�nj6TL���L#r�\��`��iȝD�5-$�Hw�^$oM��C�F�pj�4��@B>�vn�FWnꛢ�3�CoG(׳N�h���7��R'6컴�0��'>��-9���m+���ɣ�on�^�}�c|�[���.�9���v�)údQ�JFr�~r���"�O[����$�{k�E#����y�7�����Dn�7A ���&�3rMF,}��=��!=w�\C4�������Y4�������ݹ�jU�Xܛ� "j͝�	\�=���/_d3�bdeTt5 �o�;Ϝ"�5�dѸWoD�SV�u��o�7n��5���]�v:�ɧ7;��n��;��A��JB��w]�gp�]W[us{0����nmh��:�v�}���g!����ui���á�*���ez0��}��l��uLޝ��<��Y�:�V��N8Hِ�ɫ;f�lCnͫF��Ĕ ��5�@����{ǽ:��7n���x��%��:�=u!-/@�Rː$�!ֺNM����N�V���$�[��0y)VNɰ��7&q���#�L��L�ŀF�B�	U�u�J�LG�����^�ɼ��˲s����'�p^BYt��w�x��÷$�g��`R�*�j�9L�gsY�p�<��H��ok��}��V�#��{u�(�y$q懵�a�w%Sr�7{;nLtoeSa�/L�O���i1�xJ۫��%j�nUz��h�KNdPN:�UuonA��T���v��sc5�ѝ��X���z���K��Yح�/rV��U��6�rcKk�{�X���n�g�ǳzD%�f�8%&%�pN�r�ܭλ��7Gں��ư���������tk�����Q��b� �#*L��7F���4m)���Ҝ�ѕ^&���f�$�aq���L�(g�C3y%�'&���v�g/�ˡR)0<ݚ�i`9�)T�q�k5@6A�z8.]
���`�]�s7�Xʮ��u��诎��<*�p�''���eX��Cy�eH}r�n��2܃���j=�у�,Q���|��>#z�{��3A=8z���X��s]/�ҞvhmA��!Y�.}�9�Y �l;^�߻�)��g�\z^g�/�v��4��y2���W>�R8�%n�H7]�Č�H ���TV�A��w7Ϥ����������Zn�
�CK��Vsӈbݧ�XA�$3	����n���9w;��6gn=Bh��h�E�%޵k[`:��wh�򭉁{{���:'���Xu��§K�y���L��=}���M��sT��+��.{ǒ��q��w}�]�c���ucӸ��1�M��N.]nս#�¥�<z%�a�r�' ow�S�]<��/d�zVr�S���p�����c��)Y�׃#�A��͙x��l��kNH��B�q[�5�Or飷#H`�t^������/,S�қq��r���N���K/TU��#��=N�gCY�qq�7P���R���Mn��w&�)4To�Ӯ��8�3K%�%Ůk8w#�Rz@+vOZ�j#�뛙V�5A��C7��$Dా7$��0V���D��v]�:p�J;� ��M��ը�{�'��bgn�!�Ӷ6��f�ț�I���s�@;W$띷-�b��o#�V�O���ݻ��e��nw@�P�Ǉ����Yƕ��{�/}$8A��ݙ��R�)��2jF����� ��5f���Τ.��$h��sQ�V��F��F��o�N�m���(SS��f>YS���Y���]`�]�I��+�X]�~��_3��b�RJ�5�ѯ�a���$*�j�qmӽ���"a�giᷜ���k���aa�]��[�ޡ-��<c^	gn<�,�Νqj�^�����%�� ���7��h���g<R�;��w]�rM��U��1NǤ�9�svk84NR��V�q�ٷ���׭���.x��w#�]���oY=���5N�"�6Lh�ӳ�˸���snA�mR�sxJ�Y�<�-�V�^�� ��'F`Ma��}�$EÉ�qqڥ9Ǝ����8��v?�gL��ݚ���I��.W�Q:���-�*K{�:l]b�YY��n���<:�I���A�ض,�Y3��)��w5n=�ܸk�RV��,��ug��5=��w'#}g
�fl[b���C�Wvq���syc��%��}0��1դ��v�g�n���8�<�{ |q���ڲ��@,s��.��ڭ8LE�6k�ǒkTV�rLX#{�e³�v.��&�urgZ�Fq����x-��а�n-��� uս��:�sW�]��H��b�n �Ӈ$�c��M���yCy�+з��zD͘a��2k���'�Q��{��m�w=���S��d�F�{�,5^*��k��8��ݱ�Z��ײ>���se��W
,T<ii��p�
{��V����x6�v��=g,B�ۚ�׵�ސV7E�(�#Rr��
A0. �!i��{���²s��+���B�6��g:�*6�:��Q�"�Cs��<�ݙ�5�ժ|q�釖�k�w��pp��sb�+��pN
sQ!ؔB�E�tȮV�m*�+A�I�sq�^$ڹ��q�O��;�<���Wpl	�#�t�7sh�u��sug&�繼T��l�P�y2����q�C���͜�ٺ-�r�C���iX�N��aU뗓��ӊ�t3�J���NvK�sA&k���w�v�(�#�-��=��,;��n��&&��R!�zȶV�w(���ܛ��I�c��LŷDŽ�G�s`v>��&!�6�v��d��
ݒ	{ERl�p�����V�V�$@��sn�fd��y�[�;���[z���89Y���"�S��s�O�h��8���m����p%��6w]�
{]G����u�хK�h���3�ǚ_d���ܖN'�C��VkP���&��NA��(\�i�g-�q���,������o�f�78�ǰ�����9�t�IŊ4��m��H���ݛ�_4�{�w�j��]i��b�������^�q���)X1�!��9���1^p�5��r�Ob|�ǯ4oK,��V*Y�i�p��-��x��#��oN� ��g��;�g)�ٝ�t���N��5C�u�x����nWfr�1摈�=����B띝�,�r�+h@�x��p�����Gb��q�]z�*�M-�e;&����5����8����Y䣼6󫼮w�xӣ����`���A���>����P��ؘ��	GkU�ދ��C'{5t���bybL�б����vp�^nL;�V��nof�×^2w��[�mX�#ٗ��KBR�D�Ċ'�����j��r�4N�VN�۬�k��f��Sw�,}���p�og^rV�mG�V�'�v|�~�3�;5C�e��	k(�2Ѽ�CL� ` �s'	pC5ź�gW�iz%g}M�7c�e3*D"�XX!�ѻ�.`'������6��N�t����������!4�x��nʁu��t��ǹwx�C��8 M�L%�(�޻���vZ���NM��u�9����ugd��u���8��@����j�Z �w�vM��9r�Õ��w�w N��� y8���e�.i;��P��W�J�2�l�Ws�Y{[+{�x���	-�kO��޲%'m}{��i�36N��F�}9,}�uKY�{q�s���uf����4�:+��ѐǽ�\�iުhJ�9۵r��ܗtr;Hy�$��v>|��ioI�.����=�b�Mi�%0�iU��J���֣ՠF�.Y1w0s8�3�(�����W�ٷ;;�XD�w5��14��B���O=�����n�-�m���`����<���SE��
S�Ҫ��ݷFD*�����R3i�:�l�� :�Z�����)�yZft�r$]���\��܊���h�~{�HVu	�!�a�����-�"��ל*$8z�3�i�ݳ�f�Xg���q isxȹާ�לr��i�jP��eZ����Ђ8m�/8)�qP� �	;�����n=[:~	��Y�[��ٽ���(�d�3����Φ�k#L/&���v���ak�I^�����G�h8f�}o���Wd݋x�sp�Rk�v�ۜ�2q0r#v�M=9C�]Rb�DL����{�f��}��pnKPc���K�W^�V!�Y��[��tm�_hI��)��37I��l�{�C���:`��n1�F��-Tћw�ܙ��@�_v�L�;56E�۫���ٲn#VV��O�&c�͕o�=p1m"��qeo{Q�.vi�\�f=Pq�6��|{�*���R�fq#�N<2�0N݁�7C��po(���	gkl��
���]8��n2���iW0��=h�z�Y�^᫤WJP|�|�.�jz>�z�+N��9�@)��!�R��ocӗe���o)��:By����X	Z��{�-H���T���[sV�qB�ُ���C�{ˮ`��3������ds0s�3S3�L�\0���C�\�" D0�P�1p�\�f
`.�L����� \�������@����0�000\ ��L\�30��fG3 �031p@0�0P��2&�31L0\#��\33p�C300P�0��"f��\���b�`����C0\���a��#���D�P��fa��G0��G31p�0�� ��dp���0&a�`as �0�\3S ���1C0�@\�L\ �s3 0���S�P�0S�3�p0�f$<�D�D���u�:_i���O�?��צˆ�l�4L�#�:,!f�sH�N_O���=�W�-�QF��e�p�ay�O7������8�U�;"ڼf��V�D�7�5b&�M���%�a���e#5U,7��ux�?-hX@��-��%�8s�""m;���~γ�$]��2gS����(����y��_��ڴq�)�f���v��Nl��Gss�
�ihnörgZ�%P���Y-�)y�%���Hɬ�ڳR"��)�pv�{�@.�2}t|=24j��y�*ּ�ܽ,x��!�tҨȓ{8�=��CS��rܷw�c�Ao;{�X�0�5vB����K,��b��3�#5i�Ar󂩛�6m���y�"D�3o���vu���n{�$��)l�~��1�此OT��.�Ż����j�l�%9{�䑶Kc��ͯ��,��}F}�R�)ޒ�����3�G���MI�ۀ�h�u���㵚2`K��'$ٜ���/:��n�rJ��n[��+���;���/#8��a_K�ݼ�T������Rٞ�Ϸ�՚k�綪ݢ��s3�6��-jo+Rr�2��^B2;�35��A|�x�ib�����)����եޚ�Ϸ%#5����8jǋ�r��C��c9�䎅}���vS�K��t=�a>n�^v��s�h�zL���仼v:�X!R�O劽d�z��9'��EqY0avv��o]���4�͞/�tTE3_�p;�l7=�B���Ua㭑���5U������a-��c��^�H�s�h��Hn�5>rG�+і]�ةOF��6͚SZjǋv�k�2Z�x�w�A;�w���jӐ����x�W{ʱ8�˽[��;��ޞ�:���������Г�{yz;=�}J���T�ǈ/Y5&i�s]LM�j����"��T��CB�mf���i:�����I_-^�[��{3��j3o6�;�"*!�F�rZ�N_��GjN��deNz�Si�5El�y�:{5�XK���2�]�@�8�����/���.�Teg	~YU`�؟{���{y%|�r�2'|�Ed\z��<�VW�$���M{�:W��4}ؔ���o��fGJ�ʲRėq���{�L@G���s�f��:�%;��|{է�yٞ;��Y5Q�ٹ��ps@<~���#{<lC'?���L�^z�E�6b�O�=�=:1��ўh̐]������l^��F:�K����ھҖ �@����:��o��e�e��S�c79{����lm[ʊ�Bxl�;; ���z{4�����yX>pv�D���1�±�����9l�M���}}�H���!�'Y����rn{�St	aA����i����7;:���ը �P^:a��F%+�fb���;
��4�e�1�ݍ��*��sm���уL{��޾�Hg���ڱ����s�C3h�W�q^�*����� + [��&�:�v(ԋ�Gg?��k��&����(0å��Q�xd��^�~�X�l���w��묫��d�^���/]��u�ͺ=��ݾ��钞,�u�.{���g9��V�Xs`�w�7��)�8�'��L��fD\�oTa��(m�,V]����oծ��9��ID���i/Q�'��8nwMY{�׷�X���Ϡ�|�Vskd~�jSh�?r(�'�0y��Yٴ�޷�OY�x.����l�G��=���-�9��{��@���g��B&^�+��������K�F��颏-��˯o��M?n���|f����s�r�gz<�LJ��
�@���4d��GBʼ6��m�YLa�ri%�����h㭺-�F7w�5^�3��Y����]e<Z.a�&�a0�e��9P��E(�$+���Oݮ�tU<�_L�7�/n��p ��t���Ȭbb�^�FbbA8����+�y��Fv�9�5��RJ7���_u�z�/-�.�Q������k�<���%�E�Qޝ�a�`Q�p߉fx�M�^R\��m8��;{}�}�k�e�ʖx&�����҄�Ќ3��:?��h��]��"���o�/���!32?��;������Yn������x�OЎV��X=����[����ႇ{����~�ϯ>������X��W�U���<z������H��sa!.0tx�@h'�l��|����+�oP7x�tOI����U�(��ϱ����3k���cp��ވ�{}�U)��Ʌ���U����9i��{wbѷn�y�[ڈ�N'ppǛ�;_���P^��&^�w�#h�&�v8GZ�c�4kU�֪\�1u�����[�g��s����|	d^�`gc޺5̄d���/=���v���'��ќ���	���~ s2z�ݜ����[���I�-;�7;=���gN���У�|����^��PD��^ٮ?Lb����k�W�h
{��(	�� �eۥW���&���X�p��77Z�ֈ.�{�M����>^�o��֝;�����L\����9�Ϭs��tuׂ��v�&u\S��^����{�aМ�-,�'N��S����]�Ty���<�O{�İ�QY9k`���1F{v2d��^3��z�({�RX�s��	�8󹣸׫J�Pb���1JӇ�X���2�Rl��7��3���R�f��E3
��b�Ά�=$�r��{b޼�2�dI����DVHƩLաt��r�Kz'�~x�E���uD��f��� �fdP�ضd������lDFV�L�sP�l�&���4μsS���-��e�'&���p6��gV^s:~�/���i=̽�1���9>Œɝ�y�'o_��7O�X��NiԟQ�vBs���E(�Hw��l�oN����zuL���5���|j�qePq�hk�g-��fj%�\�$h���/hޮn�U��LӼ�`c�};\?G�LL���ҧ�W�������{FѓP��6om��L����{ �3U՘ui�[i��x�wy����˰�F�9�L�H�3D~�B�]$�zm��X{qu�tXΛ8������E�;T*GR���Ϸ@S~BMw�J����<Z��6�"�޿HuD����(r�v;��N��D%0 ���e�u��޲��Ρpvt���=�:��Mʢ��`˾�,���#��>N�*9��oq�~�OVW]�D��R��	�fwؽ�R���3��e�T{�ٱe��Gg��Af�k�iWژ{��J��+�5ֱ�O�ۉ�xJچ�͈h�!ꫣzȯ+�����E]�1����o҇�b�s..k�*�2BI���W��t]��H�M����p����{�o!۶(J�=d_�����W�C&V�|n��^&�Vj�V$�}��g���^(��;۷I��^mJw�]�Ӹ�w�ˤ���٫���Oc�[��Ci��o�׸h����6oLAی�z6\ �	�e;&>[��=ޛ��|�7*Œ�g`2"�!��ې����{�<��vU�x���6V��cS�|L�f���8~�����?)˂y�o{�ӝ����޲PՓu�S{��%�>���o��\�l��b�$��ԝ��Mf�~��n�{h�6-��nz��6��d��#�9i�g\�a��}ot G�bi���;��$_t�3_�\�N�G�y�Xr���}�{����;��po��=���'� �yP�;/�/��7�K�ŗ��V؊�v2�p�`�+�'f+��#����U�?���@�zf�H�����l�d9���pnn��'O�#��8/���k����;=���;�p�mL�S8��f���x1ʽ��9��LC�K[���sn�]S��N��!��v�+7���ubއ� ��+��g�r�^�(q�E܈�'}��Y+�6�T�h`����<��|��Q���J]�`{�_���W9gzu5��m80�����W��J�;۾H��mY��P\���1��unoe�Gr�{���8��7���n�����U�+w"q�ni�#Z��!&���~�H��#�g/C}�'8���<�K}qm
�=�|v��X�r�^��q�\>`�}�no������ۋ�W*/e�
�r�Q��i���7sX�W�<��J;��F��gE;�d��re�����y՗kY)�2��w�Q�q���*��VBPde��*+Zctk�c=�ξbt���:�<^SqS��{q���������.�Xk�3�7���W�������!�id��O+;�9��_	�,�����0���>�~��;Po���I�#�]R�)��V�M���<t�L����ː�^����ݏ	�6':��ˉ'�Sq+T�y��q���z���da�g'_�;���X��Ȍ�b�Cnu)ɡ9Y$�v!�y:���Ll�#*���1$�'9�r�-�Z�Q񆘖�ѧ�P����(Dᑖ��̆&�M%}}G3���wgL��8}�g�r��ɥk[׺I=�4D�xk���g	/g�����ٛ�DXv���T�M��7�S�g���V�%��i�lG��nu���ތ�����g�]LM���<�sx�Td�}p���� W&�3Wc�����673�w�c�px/tl�=w�}o�_�Kwu�OG�Q0�!.!Oyr�g`��.�ZVG����o-�D5��]WK�T��UN�o����؂�F���ff��2��a2���]���X��Yz�էܥ��[�^�(���خ�[��]z	wW��KO��|2�����x�7��o��3��׾.U�TVH��x�ۀ��׷�9���Ϗ�p]E"CE�5�ی�������C�;}⽽qH=�tm���<���ٹ��;�_f�R�[��Tg�4;��!�ӻ�{54���R��u縃����0}��_o�N>G�d��"cG�.p�m�}���3g����:hԦ�['.k�]��v*^�S��wwWru+��l<Ĥe]��"�+�[�n�N�6Z�W��R�x%nU���2g�-'�ܺxo�^;���w�(A8���v��c��fs��޼�"�e�?M��ם����1j�q���4=7ohݞOCS����]�܀��Xu\N_im��3_ϼ���<N�������m8~���e	Be��4�D�މ����d'����<���e֌V����x�T2�qn�]������$f�V�C���^s�*����U��.$��i[��o�.��"K���v7��:�Gψ�c8q<-��,�6�{�N����
���)]��"��u���u�����z��b��c��`��t:{���>�ٌb$�y[����ݾ���'-��|:�	����{�ˬٯ�r)�T�EJ��>�㏮ӈ�X�,*?\륈S�5��3�'l(�TȌƯi�F�X�!�;���e:S��kiӻV�F��7$mo���n�r�Ό�ܰ�-�2�ƭ����"��D��Y���孵˛��g1�4���ه�����ܹ�ѕ����+�=�7u�VB�'�e�4\)�\
�+ȍ����4�;�2�r"DFd�]ٗ욣[��(Aj҉�wx�4�fR[~ޡm���诗{��<�Y{,���xr�v7HRo�{�qz��>�D�z~��gq郉��U��G*��sY4��1t�,Ppø�y�uUJ�W홡�y
����g)D�r��>)`��t,�Z��GϽ۞W��������iZ-0�]�7<�H�s�4�Ec-����k�{(>��=<ߜ»=�n���e�^��^�=Wd���	K5:0VD���""uT�ױor�7�)�EFF[�>�$�4	vfI�a@�b��a��_��5i�q�y��@p%�b7%s�P�ge}�j	`M܎!��=�-����L��{�Y�/c�l+�p�,�LY�@�C�OA�1jFm��������� ���Rm�]�H�rz-�� �Q!��mߵz�'䤍T�Nf3\U%!M��]�q�4F;8t���{E�c�,z�аʗI�N����y����f���1έ̌^�Z��5���\�:n坞\�voX�����6i'��e�Iw%<%�7-Gy�Cz9h����/�˛;��}�-�:��o����8�����>Vdf��}�W�z&��ԫͻn��.�T3t�xD�L����s��{�@��٨�M�-�c�� ��9ƃ�w8��]�d����Iú�����od�A��wE�}p��5|O�_�����p��,�zO
:�"*��罾�{�5�e��h�Av��4&�vrp��2)��qQ_�p('1��]���YZ3f1���q;�z�4+^,������mM~>�9\�d�^��W���[(>��U��Q�?|�f��o�X�f{�J���we�l�+���.ǭB��(Zy�L��_Ty7�jW�؞�C�\�O�K��MK�h�FL�	�S���^�B0m��/�G�q��p���-��Ϸ��	�w�<߁6���=��wŷ|�M���u9�4��Ϻ�Q�tj�pkzkY�V,*�?[^��7���{��pV�D�ow�'-��;}�Q��1����H6�aJj]m�䫒�{al��� i1� 6�$G�gw)숞a���4
�la�po�쳹`F��׆_�Fi�+�\S^R�'�������T��	��w�e1�9t�t�����vGe}�]Xf��Ʈ��<�ӓ�%9B=!�fī�M���6�W����u�䱻n�-K�&�G���W�H�M^�#��˯v������1�ai���'b5L�z����ݲӪ�wuM�T:=!�����b(�E���E� ���*�*b��U��Df���V��%&v��V����v����W��Wn�g=�9���]#�s���g���rsэ����\�k(��:]vu�;nա��w������=�d˯g�WĴv8�nv��c�/<��]�ۢ���W`ټnƇhAxz�]�m��x�FێT�T۴�d��[�ݴ;V�4��lh&6Cc�m�[V�'��Nb���ԕ���ivݣ3�qv�q�o./��y�f��]�C�%*!�K��л�;e���۶��&��c��ѵ�N魫���Iׄj�HFw#�/-���f��̎�q��6���g��;۔{*�7�oY63�L��X�t!����=1ۙ+a��^�[V[Սf�G[C�%e�û�v-؊wm�[��n�z��ۘ]lt'Bh���Xb�v-���P�����m�ژ��s���s��͜��z[m[�����wlv�;��뀜�6�<n���<'V�;8���y��s�"�O��C��縶���нr�9�ܴ���ڥ)�ܵڍ�n�q�+]�s.k뇺��=���Z��nYm)�$�����6���qGy��]��J��mԍU�uA�L�m�#ɛ�<�ZJ�#�<����Z��&��_2�:xw+��7a�gtR�]�=�Jm�!����ɞ��۞-��n{'s�N�1͋��bhmEr�]Q��Z�,�)-̝dx���d�.5�x�F����䃀�n����Nw\�<�Ά�a7a#��d��qv��^˩=��\�t�琸�:��t������[��Ő4�����=�whi��K�n�]3S�Il�.Uެv��z�X��rq�k=��<mY,�����;��f��;�n��^u�K;1&4�;�'U�Kg��.@Y���W���y�	�\�6�<�����:u��8�nќ��]��Ѽzv���n�9���Mc�Nݵ���I�M�2�V6e#��;'U;Z���#v��Vީ㜴vrnxJ�B�a����4�<	<ѻta�ծ��Oa��>ג���N��g�d5ӗtMv9�[���W����SCun�U9�͹Nѓ]�cmklWn��$����<=(����W���CA���
���i���f���x{q�FV�N�jщ9w�[����'[t��l���7n�Fx��z����{jKR�{[�n��n�r��!�t�Cݺ�6n�V���[;r��G��U����=�q{���λ[�ub�8��N�.x����蹧�fw]�Y8�vu�v�[w��H���9��jwU�oe�sӐ�q�le�w����w��w�nM�M��:zv�i�ټk�D��s=�ܶѝb2죒�&��GR�g�6�[�]�쫻(z^=���\W<�n�ݽ�r��q(����*vxݸ�9�WI���;u6.nݷZz�d+���G��:�=��^���P<�}.+]pmtq��壙덝S��P��E���Gagl��.��8�x4v�1��l9ke�=N�ݣ�A�7i��Z�Ƕ�͞���m�ф��u�;�8gW v��z��.'ƶݻpm��u��$�}��j���W=����lm���{!�p��ǷnwK�4+�p�m�E��κݻ:���s�
�{=0U���t�����8��c�΍�rHs��ۤz!yN7l�n�0uK�J�u<[�h�������\��=V7/��X^lm��yrlm���q\�n|��m�R�!��mbc�c��1;��Y ݵ�3ͧ�m��ʋ��ɞ���cݰ�)Ό�왆����ƅ-v�n���6
�ӌC��AJ������mz2��ݣ��ZƱ����Y��{vy�����p8<��j�kx���s���j�������oodq�vSl����d.�cs����F:Ƕm���s͝�=BN��Zp`��aM��zH�wZ�d�Dct�r`b��:7m�;`z��ɻ�ǡ��[N�gl�X�ن�{O;�㓨�YT'7N��v-�ŭq�Z��A�Ẁ�z�n{Y�wm����8��9����F�=�M�j��n�w5ȵ+�N�7��q�����n���N1gSK��CV�R2z����k��q�[�%���]r���{F����{��+���u�Ҽ�ۄ��n�YQombʫi8ç�'zD��v�63�����u�\�n��������E�٤xA�b�m�؃����B�I�W�>V�AR���ـ�,Ev��4��ֶ{�����ai���Ŵ�������nz٘�cm�b�9��5�W��8�ㅗ�λE\WI������έ�7J�$1�9���]5w/\b�[��܎�5�9N��V�3pq.�h�n�[�n#��֞���n{vXpWm)���έ��@�Z�jޜ�)�&�t\lm8]��*�\S;6�zcZ�3�g��ø��k�C��%��D�,'=�]Ӭ\�i,v�8ӧ��X�^�����vk���9��(�'.:��3v�3�\p�o'.:`�n�^^v���\(�5Mk5�ie`6�xWv�k��`�kiy2;�bv:����ӎ3���2wݗFl���v'��N���y�ks�<����^�o k�Oh{E�k���1�Qݱ���\rvu�7n�ƶ�vCq��::vi�6�s��c��C�睤�	�]�.�KHm��x�vک:v�]u�e�F�q��{t�i�n0q�c�q�]h��mՍ���k<�ڗq��hd�vN������ё��j��C7���gN3�W���.�s7�u��.��:�h��pgsnø��s���%�-�F6�˺����:lu����tpt�:q�u<�[�z�uĀ�6����6Mcp�^"8�0c���rt��3�Vn:�%���Z�^����g{q�a�2A��>n�\y����tv�G
(�a9���ʎ�{v{�[[�n�;pG�|�7R��W�/A���[]��8M��m۶�`�kj7��<��]m�7V.�s�mu��c��Π���xGq��;l8�Ӫ���ۛr&�p��7&o+�ux9�́wm���`Ú��	�ų��v뛭�ў='n�E�O��]ն�iW�+n��c�zvnP�Y��|[x�[�x�2���>s�Ch.:�h�۔	�U�e�y#<u���WWA�ѸvQ��t�۷�c���W;�9w�ܘԽT����ngsl���ɠ!뗋�Ov7箷������E[�������9�fz..��/j������[��_:�Z6�[�;[Q��4-��g�ݴ�\w8��r�}b��+�������yi��xxÎ�nm�\>��N��A��^��[Ay�{t�,����0��d��[�Znq˘n�q��h�z�����Wu��r�u�iB�n��	��۳<� ���Т7V|���;���j��vۚ�rgl#�{;��ؗF�r��ݸ8뀀l�pKý'��5۱@��A���uP/C�Lk�r�v\��띕������[�-�xoE����Au���1�luچ��۞mB���g؝�݃OV����G��&��]��vrV+�Hs��lv�<<F7z2���R��v��βƧ�\;h����:�#�����ݳ����d��m���nJ��(	@�۫��\::;���{/f�X�ܑ�G={im��,u�X��x�=�g�ǈ���/Y-��1��^lr<�u݀ua����=�3�M�S6��ܗV�p��vN!��B�m�^�^n�Q��㮣�`p��x�u�gض�=��qlƙ�'&���m���#�4��8<�n��	��qۻ��v.�|���O �����9��L����ˍ��ɕ99�ݬ�{'��m�m�
��]�tv��/����C�^�ɓ��kt�n�l�N9���q���ܲ�\��5F��֢��-�.�&;F���g�^�W3۷v�s����<��vM�����:��gs�c����I4m����Q���\FsǴu����=��Ƴ�=�b��u�h,�!k�W�� N�v�/oX����!sq�#�Hp�q2�k��e��:�G-wK�]��>��m�wQQ�u��>��Ǝ��vMn��s��l\v�"d��Q{V+�J��Rn���`����1;��ә�c/Om���f��P��5��3�Dݷl�ź�;]�bC�\��\�
�V�S��.
wnꔫ�m�l%��v׮%{*`7]aݺ�8�Zu�X�K[������<��]����s�Y�>�e`0��R����sgt�a�mع�N�'FTW�e�Re�MlMX�:��\�t�✜+�s�<!n�]���������I�w8��y�������ٓ��6�xGV5t �Ms��r!��o:<��.,�>G��E)�k�+�]�m��q�\���{�mn�I�z�v�xK���NĻ�!#=�n�ZEۙ���rr���Rƽ�9��9��GlN�D�^:;g�9ōu�燤Ѯ	�Y/�Wn��M��eʆ{7 h�ԃ&�	T�{����zp�"�>�u����gvq�i�ۈ^z$���م!	�<]�i�5�:������8u��/���X_O9�HL���3A5��4���
����i�)�6]ۃôg<kQ�cku�ˈ�n+��L<�ێ��n7Qv:�"#�pΡ�3<��Gn�q��\���躆��[�X6��ي�';�=s=i�E؞gm�����3�y�58�a�8�#O�s�ɜ �0�<^ݽU{�v���Uv��۠ޭYx�=n��a�-��{q�	֨ScZp���[shm�oU�m��=���zݝ�\Fz�\�s$s*ƻ][4�4]4�V:�lC�e�����X�����u���R�v�Kq6��u^Ѳ��M����k3�qT� �㨜`��.���qܘ�1;r��n^͓�\�]���[��M����z��c%���s`��$���i{,o�v�u�c��aH�c�IQB(���!q�Tq�V�H�X�A��"�b���D����P�*#��T� ��P�1&ID0Gqq�."��D�*9�)Qb,����BD�I���X�����BH�$E���#�T$�#�"�HAEŌ�2(�0��8�b�����8,�GUULQ��B*������R���`�
Ɍ��1����G		B �L�n8���8"�H��U��Y&c�(��ノ
	���RI"�eJ��(���"��,�Y#
�����B1�$�XU�ČQUG�\��*���X*��ジ������
�L\�ŋ�"�F8���!!2H
2E�r0V0U���(ɄDDF1qP�$�$UY$dI$UX��V)!�I�����8"��� ���$E�U"A3�U$W�#�D��r."�����b��1pX�+��*�$qUWG#�"�$�Bb�
�������xffx���*��8�U����5���k�a�m�=�
G�3��G��u�XM��L��ۋ�wE��Q�\���n6˭�f��A�����ؘY8_]b-&[�
����9�.;uzxK:��iTK���=Bn<���X��։���t;��u:���c���v�Fݔ+;�^����G�vss�ێ|R�s<���`��pao0{n��oOf��a�5�M��g���wWgZ!�"�WL�&7�)ѓ��x
%���1�=�{��x��⧒�u���/c�k8{n���cB�;���-�9X��;C�񋶺��Q�a���,r�����k�Wus�3�A���z��{%�d<d<O<[�uӷ	<���E)�Ӊp���.�y���%�����m�f*���5�\F)�k�v8�ۙ��5�z���h,l��Z+q�;^��u�p<}03sە3ӯM!�HwC�E۵�}z�웒����9X���vϝ�V���\��{Vݢ0[v�*�q6�;��gm�;��v��k&��9:{�yL�������7d:s�֮>�r'Khd���ڻ\����o
���wg�w�H�hɷg�Y���\{[v�]���K��s��]t�)��<WQi;�R���:�h�^eʛN]�G�"�5�}�����;[\�2ջ\qh�`�ܛ��¦���r��n�;�d�a�{��6�'�r�N�i�������Q���W;��gl��:x��r�ڶ�H]�`�::øxxtiFn惚0�T����:��c��u��`;g����1l�R9�(%�gbl���'<�u�q�.�ۄg�[�ys��a�Nh�eֶ��&�W(�f���6�R�4�kC���7�FT_�5���Y������HE�̝>�ݧ+�4\�V絧�Kv�8��}sqxkqײ��<�^�����/��K��=�n�ح��痬n��`	lnL��qȫu��{���`^<m˃˟(�;"�r�8�����(U�(��YQ��6ڶZXBY)b�D��%jĊ��$��ZR��IAe���Rd��p�h��I�PX�J��ՖYVe��,!���dk%��KX�U��ù�q�Dðn7���}���*����!,D�-E�"H�U�� �D��b,d�;�����#ۜ�g�
6R6^{�~��SQ5�L����m�nR�9n�
+�0U8��S��J�}���d����Â]g�e�T
F���e��[|���	�(�v��In�!�j@���i��d��;U*��2*������}:P"�5*hD�n�mv߉'"�e	���₤�)��$;����8T'��~Q1S:�!%�z�A�t��oq��t����Rי��"�J��T����FjIS���A �����m�#(��.��nt�6�Z�H���`�Ν[�Nl���
��[������t��OM�:]�`�Z��gmzf
�;9���9�7}ƹ"T�� 9��4I>9{<�O����f(L�9���%E\&٨ 0y�����Wۣ�|p��j���ee-�ך:0�sTŝf�����c�+m&̻�Q')�jiT��-g1�39�z��[9qׂ��P���䏄���'��N(�_��yl�d�����7��XVtzlU[�=ɽA�sƮ�GM&�
f��2��A �wsyY�1�;�d]� E�>��+�XSa��S��e�oS��S�*�H)\�	>/q��|��d�zo�A�)��J9�K�	��QB&(Q���v8o�Q��< �6���I��vO�/�P6�Q蹾/�>w޽V8xd.�<�w��9�c��=��>��n61\n.�[�� r�v���Ԧ��$9:nM�I9ݝw�o�P7|.�M�e�e�:� ���{�.>��5��Y )��+�k�@4�nmdAS�6�݁��pA� �ky�d�_l�@:�uk6�nMt�#8H�A)� *ݾ��	B�{�	|Ŧ���TwRv��p���l��d�O9\*�̺�W���ϱ���0���ӥ5��hbRMx��5M����1!.��R̀I;��ł@.�h*��h��4(W�j�����xw�^̂A�Y��>#��"Im��Ev���%~w�|-)���a��l��oЉ%�N�,ƄrB\0M-���|v�iH�s�27�ٮ֡��\P#A�<�'f�\�۲x7s��Ю�x���Z݆�� sy�s٧�p;ٺ{8_�#��0���O�$m��c���F��+]�'Į��_%���M9mJj\�����y��"�h��L�U���﶑ �����[y�q��V�k��Ā���a�)��]��J�'�J;qE�{s�N�c��<v�i�6��-����a�!���k��y�tV:�
	{ZW���u�T�\���5'�A�+&��v�4��}���ޟk�s�j��Yݨ��e�I����|���k�VWd�T��.��17V��AW��$R|�&�
�M]���B;�����1QdR�9�<A9y-@ ��u_ʳz7<�W��3=|��.P�%L ��u���X�Νp/c�u������\s^q�������߆��L51-���t�%}8�$�=�vg''f�ܨ���9\vS$���
u����hn&GU��__֔���m��(U�ՂH>�I"�]�A�V�P�՝B�pSUURdњ�5�H@>9o��|{�6en)Yx�A ���||��;�/�[kFD��!)�����-�ܛU#IVO( �O��s�$��v����پۛ�{!���g����a���s �Fwz�|�.U�5�z�S8Hy��Fmq^�}v��Y!��i_a�	�!T�(�w�v`����f��w6��u�(�m�;�p]#\��m��Nf�4n�s1�;�do����b�(��7�Lj��a0�bj>�g����a���l�l:ٻnka8�7�;���;�+�x;"2��9ڡ�g��<ȏk%��Uݜ�X� +��Tc۱�r�A^�`Fv�T������ݴ��&�ۡ+u9�Pv�w.�]�s�����:�չr�F��瞬�ŗf��p��A�����z^����.8��m�����B;.�s)��ݭ����q���n;lpV3r-��C����׫=E��DU�1��֧����[0�2�L?�w3k�����i$���G-@��gJ���gO�w����p��Æ�%���1��/'4{�׎�h>��<O���w]��+�W����E��I4�N��*��Ї)���.����/�|I�]��j0���9���t�m�mڅ�욅)��K"\����驮3�H��~$���A ���I>;n{
���ו_,�&V#�P$����D��+�k�
�'�W蕄��0��]v	un�v�yz$A��t1�FP�w^�ǘ���k[�^�qf�����q�ki:x(u���$O���P@��1#:��Q(�{A|H���"���cDum
�On�*!k�qP�:0�r�S��A.�L���Zޜ��M�^F;���	��n]����}�tvn��+��C's�dS�3X�ۂ0XZ�"����N���[A�\�H���N��`/[� _�����߶��H[�:Tta�J/ei������[��B@�}:�"[� �y��kT�� �c�1҅�������C�@�J��W�{��r��Vj'V��~$�HH'��*J��޹+�Hʩ��	�,J����m�Rȗ?!2�gMP�%��닧p�tB�rWR$�{-v�]�w�*ݸםe�a}cb��h�d-��{�;wZ8��uϮ7f�$�k���4�J�%������#��UA"�0��D����n���3a�k���"�Ԯ� ����A�&+H�3BI"b���,��T��J���ud�Iw�ϭs��C"��W��V��J�4�r�Si�����	%�۷�/�v�s���/#���[h⋘��BZ�a{M��|r}�.�DQ�:_I��V�jݙ���2Ӛy1��Tj���yU��v�V6�>��6�h,dP��Y�޺���!x�k�]�<.6��L�4dMT {iRH���+��u�����[ܬ��붯eUM���7�0�# c*mx�S&�������Y�F�'~����Iv���f\6X$�k�����c�Suy���Q�̘��̦�f&T�M��6� ��q�n�V(�t��`���`��
����󪪓5j|`�qo�/A'���Y]��Om2�}S:�k`�y��SGI%
,7	��K�7������wvi$���� �]v��z�t�/3�f�Vd���9�P�Wu�dGS�@�|Ui�m�W��.�g $��zŒ]v�$R�*Lɪ.%ݢ\���}��b�"-{_e��$:��$ⷧ�{8�F��Ș��_S���:LT������y����ݴl�f�m�]�J7�vn{{`Z/w6��������A��.�Kw&U�kn�r&����J̋��m�r51-��-�!$�S��!�&���32�%fw_+ �]=�⒅Y��ss�*^j^��)AܡY��t�XY1�Ǵ�t`׀��
�Fx�������0bj���3^|f�_��H��A%k�+��\˽�T�;�H=[��Ip�nT���2����(~���^=��ʷ.�`��]v�$����'3�zv�;�	S�XI(P9`����V�|�g��Vͻ-�R�"l�맀��㤒�Y���賄�D�\JP�$e���@�d/�H�I\�O�����S�yΌ��N�*@�R|:$T�$�pA.��2�P�,�ݸ�z;����>��@��T��'o��@>'�m�ٜ*sr5V���	�nA����#yl&n+���N����L�d�aL#ę4������ʄ�d��<~���;�;w?/��> �]�\t\�9+��/qtn;(��������8!ɩꍴ;'v�{3�?��||C��z�h�Gr��G�E�v���R�h�Zؼvsݸ�4�g���f��nێ�ŗ۵��1��!|���Y�;���ü��ܗ3�qm�bz�����t��]�c���͗ul����sC�#c�FO�F�tI�j�W�s;�tk��=^=$s;p�|��x��G����[���v�����ے�?����-$�<������\�H.��I$����[4h#�+fq��ΤI>=y<������&��yX;��vA=]a���WN��<]��D�v�]�L�6jaq��)�͹�J�"�r�n&\��L���UIz�z��:���o���*k��:�u@ ���eSEĒ��Jj�Ev���7��)W�b_��/k����%��뿒Q���x+ͣ�hp��g��I����jFR2��-A ����dkZkx�ZW�$m�wd�mHϲ�'����LD	72j$�0s۱&�n1�����ڵ6'���g�v�=�y�*f&f�	5��(z���$�|Z�4o����8}�$X�ər���B�t�F�@a��z�m���m���5!�w@�7�����c��kڇH&�p_j�X��}�|!�����bn��z���^�Ab�w+J���v�j��i5�k÷��aϧT).MP�5&k�~��]�O���H�L�lh�518z�*(H����!��D��j��35!��*�M^r����'c��k�괠���� ���Ѿވ��D;���go����3!�����ي�%���)o��+��R���x
�i�R���	|�}=P{��J�}���R�@��.g��m��,ĝ��\����q`�Y�rdx�X�Ի�H�ĥR3���J5^��P���q�ZG�k{UݒN���B�8�a̓2��S.��=PC�� �g�}˘�	�#"�� �2�y�V*�-�D<�=w%q�[3 8s"NXV��Q �}:W�9[�1���]p�U��~��xu�x��1MwS��]�Ǟ�=�g�[����%��dk���;90�;軽C˾xx��e�QZ���K���wn@��e��R�����l���B��g�a�R��5u�چ����vϯ�Z�S<w>�{/��\�|�=thw�չ��i�\�Ş�Zp	���W 1� ׏'c��N��F��6�P�]�lW|��^�w-ɫ=}O7z^7֝��=K�B��y-6�hѫC��b������J�xl��[�G���n{w�Y�;j���7��0��r�
s�0Z�{4_7��헏�N�^|�SZq��'x�wQ�Ǎb��o���U��'�PZBr(!g�'{����&|�J��5[Y�Ķ�ݽJ� �'<v��xn\�G��{��b0Xr�*}��ٴzX>����-<�$�p�A:����T�Lb���I���9��]���7�Fs��ޘ=|�hr�I1�^���q*se�MS�ؑ�j�S����a��l�:�f�MB��C���KFhs���Ԋ��F�1�}�?H>Q�u���{�a@�u8-^��})��8ԛ|l}O�g�:{���^/f��M��r�y:-�N�䄥#1�#	"�^�jd����ID�HMLHpi]Ӱ��⵴P��M��wCw�{��������1v\�:F���i�MV�öe�~��7�[��C%���>'���︭2ll�8민q Tm�X�z�����5��>����p������>W�x눸�*��"�Y�DQ��s�qpA��� ��Fd�"D�QcA�b"�**�A�f*��$$�1ATTD$&$E!(�จ�+��9���㈢� ��Gp\Q� ��(�����r
8�"�� F(�f1���GB
*���b�*#��$�$�QqqDpTE3DY2"������	UQTQQ�1Y�qH���(���&"�� ��(�dqE�bGU9G"AQEq�WDUEQQE�qPPTQQ�Y&Fb���fG�$���*c��d�LPU����������(��� �$���DP�WE� �2AY*&8 �DbDE�GqG�qF.db$Ȩ(��ALp��RI$T�WEŊ�TS#UGEQ\qEDPQB+�8��(+�"
��I0���!$$�EW1AUd���`�(I\\��E�
��!�TU�T�UDEd$��U\U0���GB_q]�J���:�ԑ-�HdLW����J�6\ҙ��T	,��@	�/�J� .����̉8����u�
�lje�7?eB�٥P��������A��Q����P�]��+Cȯl?\gGuCgɦR'1'ɯ&�=7����'�֎��n}3�^�@逞������*)�'xD.�@M��O��w+:�SYǬ��"3nP�nZM�kH2&���b���'5ﳱ�fea��$��q��V<H8�P��.�V�J�8�s$�l�L��N\�@�(Y}�v��H]C7}V2���d�|z��.�����M�!Ùr�;�߭�/�;v�2NnN�O�����=�i����?��8�������Yԙ�R���O�#�I1�H�c�!�<P�-��]\�+�w��8�Y�&{�߷J�i�B%�P귒S-ʒ?��y�]�FOm f^�����*r��Iw��� �94iў/����5����=Pa�.�N=g� �]<���h� ڼ��wD����9���j_�&r�ɪ�$�z��Am".C��'�,Σ����+�nեS�d�2|9dv�{Z$�m�]m�"j�����d�a��$���6:���Y�L�"��0j&*1��Y���@�O�1'9en��.k��Dp;zڲ|I��Ay-�"�bf�*LLՉ�����^��|O�5�vA �gwiO����5{}�â�(��3]��1����gn�x���.@k��F�ع�aY"��]�	�{H�ko�}��Y����P�Vhem�ꫣvX����fc@����C��ʎ5�v��ǃ>Ǿ�,>W����/d=������	�n�52�dĨ �:��^���r<��g��A��-B�#aVE�L�(�֖�ف5��q]�)ӓvWg�3ƋvZ1��[C����N{����9��9�łX�v�%����nR����[�&�a�y�8m��N0�r�%u��;����sv6ϯ(imGkW))�uc���yl7F�U�����[40v.Ʋ��{=��4Nj�<o��]�2v��X�c�]cR��d�Ӗ�˺p�n�8��㣢���n�Y��I����"�� s7r�FS�HZ�(��uݒ!��� �z�i��l�������2�^ޚ�B���s�%��vA ���yx�s�@ ��b�sg˟�ДS�Z�fO�,��n�x�>*�yG��;2���6�-�	9[��+��=P%|��
a�)	�2��W]�����t�$�s�"E��m9�)M��~��o��P�I3�L˻�7=B��Y]�q`��34��H�S��A ����&�>��#��D�ʍ�����.2�+�'��A��Wn\=��f�n�h�E��LD�!�����ٗp�HM�w˱ӠA�]�ЂI>�����1H���� I ���!%̓3U3MH5�5v^����ET�S�)t�S�4�����u컊�[�����X�!r�G��غk}�����f�s&���������fʔ��W��>������ mWĂI_mq-s��������̫�IB�l�k��c�Dʅ��I/Vo\E��-� ���Q7T�IVt�K�޻����pL��,
n��.u�
N�حY���<B�!�޻'����x��q�f�������K}	�CjQ�b��_��	u=�"�Dx�+t*�kzp�|H����.�i]0eG�vD���KD���!"�F�Y�nNθ��w^l�͌u�.K9�^Na�������LS2�
fo���v��Q��� ��"A��z�l��q=�O���fh��U0UAG��{�y]�D�o�.{�F�|��O���Ň���������>K����T�^�=}���2�iH*�����;�)IÓ���F��e����{���7M�^�'�ֶ����65�3���/g.���0�SH�kc�.�m������{���~ �O��>�_m/Abj'd���*�2j�Ҏ�ެ���'�*�]��Wm 	$���Mm�U#В˽봩�ȸS*�N�[�|n�x�m���`���dS�@�N۞P^�ݍØ�SIz�����$MEq[�s�8�6KƎ�n=��f��Bۨ:�!�6d�~{�P�R�#:��W�{��(P|6����*z�d�
k����r�h'Y�2B%�'2�ӗ=BD	/��m��i�ω�')�";ny@#����]�nz*��i_��L��ȓlQ�-�$��J �vi�옼�WuWf�x��\�%����C��"In(O��.�E.l���f A$J�H|H'/k��$v�^s��Ŕ$].�%:3To���g�C6�՗|,2�M�ɵ+����uw^O�����_���+��1.-�9'0�|=��_��	�,I��>����L��~ߥ( ��X�yU�ڷncSr��x�	9}- �.���R�����Y)br����%L��{l��:Eud�h��:{�lu�Vj{u������e�ih��O��$��N�I+�޻L�d�T�W�ޮ�	�'ǯ'W��|MiE5(!�2���v�(s�J���脡$C��W�'�|��Ăq���'`<���r�c�YK$"[bs.�I�^J_n���b��6ug*�A ��� n�밗���&a��m��]�O�l����e�7ф��-A�G[ޱ`��:��z��+�zu��_��%��i?��w���O��Τ
᪨�r�p�E�]i@	��߁�Υ��ng/�U�gA_��9~�r6 y�x���O�v�d��Z��UW�P�j����f�R��E��GI�_�x�N/ju���˝[}Jp�|=���\zG�2d���UU�����#�8ysƶ�E�<StնP�p n�Ht�&E��vx9	4���y��]-��E9��l���j��������hsɉ��1�6��덋�6�������nN�,r�ݴ��ۇ�y
3��pؑm����e���ZF,���s�����6l�ܠ���ӹk<���u��{���h�P��m����\V@ld��+-Ӵ��5�M��vїI��v!�n�r�ۇl�˻N�M�5����Q������e3���j����uŨJ.s�y�	o^�nV�z��%N�i"~��!;�Eg8�Y��Tۓo������v$�9ԉ4��`G��n�F�]_)��2�FV��jQӎ�>#h�,yc���̼�G^7w�FϹ�%�]�$"[bd������-F�z�"�4��˻ �zwh"|v��HQj�Fda!�޻��R�EA�������T0�}��6�]�8�jo ¿X� 	��b_�r�3 j9�?��?]�yϣ�'�����8�����Ɯ������a�`&Z��J}��D�����˽[�,�A=��$�������KOn�]�J==�+岠~HP�m�2�Ks�"A�q�8�LMÍ�	Z��.LV^�Vr8�>���̦����L��4:�z�Բ������N-��G���x��,�(^���F+j�Ś��<< �:��޳�A��� ���ROSd�I�^=2�{m*�Y��KSN����I9{ԁf�s<���շ�w�;;�*�����K�a��53.r![�.'6Ǫ㲯�$]�H$ݽ��&�7��w���w���^��P���%��B�EU�34�x�F����z���	��D���m A�7����jf�A+o��tˁ���?��")��2��E�r�*��N�(Z6�p9��q������z4����!FU|I%��@�@$^c�r4�Ow#F���}�y5HN[��ى���C��*��b���)X�T߾��I.� �>$^gu�$��v�1W1W.&�րH�AL�4j�k�&�x��HI8����vL�GE�̢̝�+Ę����%��p��	v���a�ڼ�F��ie�F�,�b�(q
�È�X���.�͙cex���������|O� ��"@������ň�њ�$L���Cc�>� .�D|l���$��6�QcGw��liu~!�(�uxȡ�Q���u�Z>#�� l������]\Q �e�w�/�hf�zo?}�9���ﭤ֨��#t�)����n6�k6w\�\���A)�BK���*�M��ڗK!6�8����O!����j�O��u�H��fzhLCVM� �}��E����Pfdp&�T.�N���M{kj^�T8�}9��>���I�m"A;���x!�ڣ��({�x$�0?��(�Y��\Z��Wm"5T�CPOU�y����5���Z�W�ʄ�!4ۗ��dn�ot�9#��>ݻ$�z�iA>;q܅���69U��p�7�t�1T�8��f�b7���C|gs'Tj2�R��t�kS�7�=s�8)raKb���	~xx{�> ���aW���������_�҄�g��t��璱n���N���D���ӗ֧N/*�f^ʎ�����1$7.[�!hh|��m�ǳ�:^��΀mnEA�5�����~�z�\Yf��5�~�A^�$v��#�y;5G�Ƴ�N.������!�v&��Bh��+31�	'�'KJ�d9�����@%���$N�>BA �����i��fN^y/�����̎�
�M$�-��Q'Ă�fЙ����2��	ȭ�^�����Y3.`!��Y��T���؊��� �x��^ ��݀�H�o�����K��{�4�A��mBM�L�خRA>9z��q\t����#�u� �N\kR	7|������L�Z��_.�W�=��;�⿐�wa)��R蜊m��ʆ�u�"�.��e/&q��}�MSn~�1F�����R�{������=�6�]	@��(��*��qƴ�Z��[O���y{f�f	U(���8.i�
Yf�&��9�I�SK7!V����7���*2Y�i�Ud�4r�y}�^_;����nj��)�|ߡ)�*�����J�s�#�w��G��y��������`:�{�������^Y��t��.��#绶7���\����#D��6
�b�z�	R�;�Ϩ��wc�ܥJ���?�[�Ú���Vi�s4���&P�h�v�eHyNw����w/HN�<w�g�m����]�e����9k�����8=x�֡�*�H�4���c�f-񼺜�~і�sdhR�T��؝��[ǒ�hY9qT����;6��6\U;i	�s�[��}�:���|X���۪��t=��竼�G��}X����'��S����S���b��~�<��ִJ�Sj)ԘwpM<�)�H:�Kt�8���C4f�c�cٔ{J�;�콧��{6�,���s��jH���R��` ���x�Z���G�g+Ù� ��A�O���zLH�KՃ(���m؛Qj^čr&n1��M[�fl���YT�h]�9��0��)<í���Cw���=�W��,�ʐe�no�sy�.�eU���6j]a�$І��'	����2I$#����̒QGqW$�"Fb����",XEPT,�*8$I!L���	�"�� ����.+���&$�D�r0DGE�����*��⪃⪨�"Iq$&."�rH�TqH�8���$�Y""#$��U�H�GEX�UUU���U�"�0��9I��F0��#&"&*�H�E��b�)!!�0$dV(�UpT�(ɒ1QD\VFb�DP�TQTES�U\Q���8�#2"���EE$ ����"EY��X��DpL\E$Ɋ��*�8�, LUT�"�!�q\�E�UȂ$�Dd��*���(**��ɒH�a!E\��qqUQd � �(�,!QB+QQTLSY28�`��D��.
��"����
��$�DQ�d&&"�����qH�\S#��	2�+�EA�����,�I /c���5o.��.����uC달���4(��1Q���k��S'2��F"k'X�)�pw�ɵ�
�f�m�jFvl��=͙����q;n�����f7n�*�6�����h�6���m�U�j�.v.u��c�6�[����BlmA�2�m���mk��r���&���ɔ9��zq�۱��f�]�ki��t���|�5ώ\�:87ptg��N�;%��>�Nó�h2vm���xy�p=�&A��}=u���ca�r��n�T���k�l�Z-γ���=\�v��O9-�ɇ�vy�[�.� �ײ�zǷ%�]f5�v:�5�u�]�p�Y���Jq��nqu��n��n�rW�p���������j�@&�j�\�ް�hy���K/n5�n^ҰJu۠�f�\�P��N�o<��(8w�e�u6�Xx�>;I���Qbf�:���7V�n4�"��_n4��h��,`�m��l�v��k���=��2cJ��Gd���V�Xܲv�GD�ư�:9{vyۚ7dv��dx�9;m�غG�瓯Q�nc����%�K�lH*h�SL)��6�n�b3r�W:\��l��Y�E�q�|�S�S��R]nձ�
�cn��M���Mυ�����Q��1�qr�On��v����<��֘W��Vé�9��:��nui���ׇ(��v�u����U�#n�^6g˴�";v���k'��]��m�F;%�Sy�wF���}����pz�7=ssd@� 3Yۭ�98mb�dp#���pdS�8�Y�e�׫+c�מ��^�6q�'Tm�ܙ��]�Num�MvA�����csuj���q��n���5�&��'&�^�Y+�+q�0۶ŃtA���m�4vm�'`�q��˭���0�u�����7��K�g�&{!n��7zWnp.���壷f�mɷ8v�omˎ��k���Qۡ���:Q��n�[l��v���S�v�w���]�s)����j����n-Hە�p�Ck���w7c�]Z�����z��망�
U�&�,�q�)��\�W\6nss�ǌ���ֹ����v��r�ێ��n-��&�i�b8���&s��n��,v.�Q�\�{;tݭ���ص�����;u���)k�����p��8�����8x�j-^ݣ�B���ͧmힵk��;c�G��P��ɭ8�*΃ۛ� K���{qCz̸ݻ;�J��2����s�W�XI�����������D
�ȅ�(e�5$�E�>��2�i��LV��&�W��$q�I7�b�&	��̹����wOۣ�+��P�$]�l H�c�J�����{/��(pl�	�	�SUvfa��$ocv,�\]���9ͺ�	�%����/׹�ȤRH�M��'*}|xw��qy	;җ�w3]߈g���L�'����J!Wd�|'��3.`!��]ٞ� ����v)	��I�7��$��<�QӗN�*�$��`Ѫ�<��ۢQ7Y󝄛�\�.�RF����v�&;Avc �&"�UMzd�p-��D���u�Y$��P2و�>��6�uΡ ��Qp߶�2�jH`C��:�b�qs��-EcI�.�<���ݫ��=������yl������0%c u9~��dj����a�m��QF�������gO��;s�$~[(T7#5�[����3Ú�B܍/�a��L˚��X�H<]�Hw��'n���b�Go�;O�u�H�,cBh�Bh��]�fzS���gco�k��G^�'ăw���΅�n�~:7�f��+�e9$	�I���M%	B��:�'�&o��j�]�A�Hﺐ:��Q[5Z~}3�����x������ ��պ���;k�����6zi0s��ߟ߽��+&��~}ٹ{~�	8]�>$]� �V-��v{j3�����$�n��1�Aa�5U5�P�wk��q�t#�W$�1ڰ#a=�}v�����'V�^8}w�f��<WP��!���?
�Ͻ��a��t���Qk;kՏ�q�.�fN�,�
.�6SZ��HY�K�컕Hv[(�#0d���g�e=w�<(\=8�&�`������Mo�$����$B����P�х�L8&[��N�w��S=p�v-9��'���Aw�A}{�����ARTf^5jx)�&I1&&Re�I9�vŎ=��.gzTs�	�W��x�x�	���vkNd�W���<�BO�|K-ӫ���6j�-^��&���:�]�j&!?�>I��+ٳ��$R�&�tq�� I�Τ	�@�|��Dl�<(M-e^0}s	,��I�Ez&eȟ�[DU����~*/ww���H`�n��@�y��i%~�����e���
4��ۢ&M@̗\I'�b�%��mw��U;�$�.��JW��v����fFC>b�v�jv/��<��!(]��BIBQ��ݐ|��f�]��� 븬�:&�9k�en��94>�t���K˲_9��B'Ik�n��b��P؝�\�d��cEO����uj����Q�{� _ĝ���-xȡ��L�H����>$6�Gd�X��W�6�N;� �}���쑆��\����啐�B����22�5�b�ݭ������c���\��e{�����߼¨Bh��g����ۻ$8��^5�.f��\#��X�"	#u�vM�d� �$p&�r�s�IntϞ��Puk\iM�i��5d_l�Aӥ�*�߮���'�虗"p"[DU���ˋI7�!
��Ưt�f�2c��v �c=��i%_d�_*RC�m��e2��*���y�U�:���~�I�q}��
﹛LLl��7���q�I�>pEY3�wĒr��<�e(�*;���J��|	7}Ԍ��";�ٳ`�׹=��&�L�[�FsY2��$z �]F����_iY9���x]bRF*���FIٗ��9��w�Ge��0~���<�W�|5)�����Kr+(�f�驻mk�t�F
c�k�a�]�9ɣ��9�������ݵ�;��t�Z����{9^ɼ�y�)7^r������6��Zϭ*�m������!����B��êv�vz�f�:���I�u�mG�n
#�>!����:�\���;Lv�����7o]޺v���o6����^6��&�[�ۏ�ѻ�c�����%۳m�؛����z���պ����Jgs!~�	L8��2e��
{��׼H,����$����p�MN,ށ�=j��#!=�	��&��B���]���D��a���2�`��{!x�n�R ��wooT�ٶ/{;A9�jbfL���A�Ҕ	m�R$�)�S��Į尥��`�}��e�.�R$V��S2�I�K`��Xﰝ��P�N�K�Tv�W�%�m	�6�;D�Qc)8�j��{�* �Q�9�ۆ�S+哚�"|s�48�u���;�=�^$��t�(W��Q9o#Ւ����L@ؓJe+r�71�dKz�ESc�X�������% �����)�r��ħ��<٨I%���I}�Ղ�AeY��1�(�	-��$�p4L�B�f�Q���~9Xb�k6��]�[X���rm�/��(G�=�3ל���^/.�7ߚ_����Ú��]�ٟ5	�m�Uq��B���� w�ߗ�(#��=ٱW;߽��qvd{i��=u�C�m&'dw`åH�I��Ղ'D]��TV�oT��-�s�_/����-�<�%"Dڄ�
��S�{� 5~�H7��Aww;�I(��M��Ͳ<�1���\�t�eȍzf�`���V ��^&��3��$�ւ$��ۻ� �lWl�x#|�vo߿O��M%м��'v�m�g�B��2 ݈���k�k��'m�����~��ꮲ�8��@�osVH'b�e�n���,<̭o6��%鋘2*�(��&��W9]&�:d�]t�'Ē;�w`�C��Că����Ox���V�w�	�2 P����f�u��:��D��җ���5K��y9�!�6nd�7���w�����Q��)��5�?��U�V�Zۛ9.�S�24F�V�_v�5�E{G������8O����H$��i'���8�p����W�ȗ�s��ti��-z��ş�At��$�Ouz�x&v��gU�Y�k%JS"mBm�B�j�'�����232cN�/�̖u���$�=�	$ݹ�������n�Gu"z��|��sv�"�5�R�q�n�`��L�㩔���ԃR$�Y����L^���/�{Vm�$���H@'���ULN�K;��b6���J�c�B��S �o�2�K3�[���̫'�;��ԴO�Wm"B���!B�u�a4���bD��r)��i�5מ�{��?_�^$��B�Ns��I���	�s�	�P&hȁB�f�Q��䌺����*��H$2���o���{Շ�����Ȉ(ֱ����{�4��f<ryj�EK$���ƕWK�j��d�h00�b�{}Y�%����Q��Ef�����v��W�w��˄Ĝ9N�.z���ۻvf���B�����K ��t�I ������n��ڎY^�W��	��M����p'n:���[Q��P�c���Du�8���n�1�{��3��UQ�T� �nZI�{�칊��1�O*�喯iw��?lz=29!?�nEW/�.--u��#g�c��$�E�WA�|���<���y�o�OДj��0�9�j�Y�)@'[�ę�z2�Ꞥ	�%۝�__������\�a�$R���1yB�Gz�t����'Ăﱋ�1tꇮz�P�R�J�p�e��ݾ�O�oiat:��`�j�x��珝��.�ix����]:�&�X�3&���a�}��O��E�u����7����/$V�����o0��z=�l��p7�D�zi6�M���w����7�m����O]a�Utv����3��f����R�l�������j����Ŷ�t�\�b=��k���W�p;c�/6ݱ�q,�u�e���n0����[u�W��%��9���ϖ絜<u���1m�7<��rm����a�ݺ3�m�wN�K���k��R�؃s�nZ�m�u���ilW=j�cۺϖ�l�68���.`v2��piүA����ڗ�O��n���`7l�Gk���,^y��L�`a�X�z7�g�������v�A�����>$�o;� �}��d���r��vt�d�k�j���6&aL��	���t�ES)��������ĂC��vI ���6�qT�;��ڌT��[�L�L^���7e�{b�e��$�j�Ts�*�!�|�ذIw�@��T�EH���H�8�r�W�z�p�1� ���UݐI%�:w�\��2���E"�uߌ,f#"$TT
��&�3����q��)p�9C�|�I}yw~$���^'����t)}�w�=������;��]�nZM����\G�p海l��۶�j�e��dx٭������n,�Ш���3�}~�H!�:^$�n��2�BQ����=뻰I'�:�VgDD���!8�;�D��%D+޽���-bu'&nD��W0ov7��MB��M�B�d�y��t����g]>���{���l쑇<l������x����3�E�V����gR'ăw|��CLV�r�ϧisw��{Z��țP�aK�Ө$���o&�.��yu߉ �{3�T%
��+��A�ND��n\�O��ˑQԞ�pL O�f�J$�6��s{k�d��Ħb��]�BL�QS 66���j7y�If�m�ra���fL�n�#>��R� ���^�|H�|��u��sS�oמ�[�>�$�51?|q��e���1�ۓ��mdv��[��ۮ �Fg�������TL�5�"�G�q����}��ح��a"�˅�(�|]��!�5"��4*&j�-w]��Pp��7rw�I�{�Nos��V�=59Y��VNHέ�1-&�É�D��%��v��I=��x"q7!h���ڕ�Ҙd��u�~3a5��?Q���N�H�m�4ȫ��s���4�0eX�-���M�~����@d��V�Ёѩ&�Y�<~�(���h،�%vH��J�˴�<�ө�C���EF��e�Є��瘆l9f�;{%�Ԏ��m�?f�F��OT(�-��}�ɮK4�6w��o3�<���w/��\uRw<��S-��@��g�({��Mk�ӻ�NEy|5��c倍�|(8,�<C[&�<�տ��{ɸǽ7=�&�5oy�X��k��9�fh��`�!��oh�y$��k�a`>���Ct��y�.1�W��@a�xqQY7]|���z0��klJ#��P%I_�����<q��,/Wq��w�R{�]�����LI�6��xV��b�nY�y"��� ������[}���yٮ>K�xĤ!ܺ���V{޺+�N��hx̸��o��w����r�{��4�	���ß}��c�Nф����iz�b�n�L�{����n�`�����;k��DG&�:w��\ڣSn��ẒaVMe��T�����)��'}�]�<!E�w�u�w�f���o�6�O��֖���z/�&����� LqJ[�-�/l�65�®�d�ڱ2��&�aU�#(k7n��{�*�z�u�5
w��{|�Ko��݆m�l�Gm~�6��xd��0��,��6�y8zJ-��A��4j=K�G�)�z��k�a��6�F1��86��l&����p_A58$�=pj㺼��}����8L�ȓK���e�*6�)�����V�zjqZ��ZNz�'���I$+�6DU�L�����**
����TE�+1Z���UBa+W�
F*�V���PFG1\E1I&+��"#2&
�e�l�DpEG9�U\qEEr2@ ��#\�*����(,b��AH��r�#8��F$H�*�q�WH��%�K!*���,p�F#d0Qd"�
�ArHɋ#�DDEW�m��B
���"�."F*$�"�2b5� ��LG$f@c����#� ���1q�qH�19�C$�#FI�LG�EI"�8��%�V�A �TG1��T`�1��Q�Eq�A����`(����U�d`����sL�Qqŋ�a1r�R����D���"+�+���c�
�E�Er ��$�d�DH�q�rH8�"8�A,�"�p��  �<���=n~^$f���_I�#	��j�{�bc�Q�)GvO�A��n�Iw�UWX�E��͑~/.Z�OA��j���UML]�}{b�$�����S\�&��
ެ+�ݼ���﶐&Ȧ˫�#����$���r��]h�=�[ɂç�1�Gu��ۙK!�Dv8�U{5GL�Ӗ�dK]w&���;{n�!�m"Jw-�F�v���W��K��ݻ�"�PZ&��L����%���M[s[<�Ƿ�� �}��7�W��5q6���q��C	��2e�@�]�du��	��"�d�lU�7�@$k���$�﶐'س�ɪ��B`��&��kr�FN�A��v=gē���t���h�S\�}z�Bdu�/E&'-��q~���̳6U��8ur³R*,Iݤ�6)^L2�*�o*A97��n�獇>������1��?�=�_�{g�$&`mBr¾_�Ӥ�������5�վ'�f݂I.�i|I�}C/��I^�"!�D��xт�E�3 ]z���`ݞX<����8)�ݱ����nMTꊩ�㗷�`����$O���7��C��E��gH���v,�z�%��́�2%�,ΧP����1ߢc�	'b�e I>7}Ԉ �7�����gVWz+u�0��bdwp���A�ޤ �T��ҳ�r�c��'��&�(I]�:���'"�I�&[u__l75upeg�<w2P$�w�AM���X�(H�R՝�&MH4EQR'p��脒�������������W+ĂAw�HA�|՚���E�UrnM���a��b�2�S�Qp�>���ȭGf�6��	�w^s�κim�Ff��ؔ����	Sk_��n�C�|<<<���3Q&b���dL�R�.y(�#�,
��xѝc#�!<:��Y�,��_7:�T�^��p��$:뫩���"���=�-�G&t�u@�$x�M۬���[F�Mη��V=]�v�ں;�l�=�ڐZ��\�%����h��X��{;Yn�W\!v.�����.Q��c���[�q��O���n��ܯS�����0�K.��qn�'9��`�wh;[\c�ۏ"�&�;�p�vf͓�^��}��~��1d��Y5u'�.��G�>�[�����{vm�m҂��3�lVܢA �����/A�H1���U��qj��s.�̆��, �]�A��Ւܵ��_�{a;���R���rϙ�.Ϊ^�K}�X$"�����-*�R�*2�]D/�g���!(/u�0��S%]�"�Ȫs�B2�w{vO�+�D�Is�$��;g"�H9\�Jk��ܕ)�$��Hۥλ���.^ܘs��A���%Oj����n� gl�e�*r��X��q��^�#�Rh�(�{�<1�X�%==�;�c˓u�c/&�u��}����r�Ci1?r�x�J�n\Z�J!�+�8%u���Fj�W�H��}�iG��B%12���]��%�\��M��f����?D*�lZ�y�������V���$�}tDw���18��C���y���5<os��髝��X#+�WuB�Fd�? <<��u�~��v	�>/>��pNd�K���FkeU��8
�1ꙩ���z��Fgm I �ȃJ������łA=���A>/;h!�#2f&���� syVS��ĸ<����D�A��"���jb�7�6�j҂�PzI�35`�:�|IY�H�ә�{L@ي'�+�${�@�U����mBw,M_���������,۱��5�j��ثn���\���4���\�E������w�5a*�ݿo���$<{^D����іi[�۴�Iw�%�WfB&!�����e���2���Z�5� ��� '�܄(Yy��^Q:�sΪ�U��^�!3/�����+;]%
/�����'�'�y�,ַ�O���ܽ/��e���N���|LZ�g�du�Ǜ=LǸ�����l��RD��sU˜ܺ(�e}��k[�$�^=�H����Z8X6̗3^��{��=�V��J9�$��Ax�N�v�sy���dvP��T�I�>d7��N*[��qzF�2�Kk�'_���)5H�U�"}�ݗ�Bu�����;1�T��T8D���NHn��c�����[��	�ݮzݵ��'������%Kjf^�k��(J!W�]%� �>�f2���F>��)+�`��D�ΉTD��A�1UA�'�Ƌ<�����[��J}� �7m�4bGr��g2��k;^�B]]��4&�bw`��R'�^�m�$�*��ֽ�����W~�P�,��ե��$���.XW˝*�3"vj����|y��	�����9(�=|.�kD'LN�n�?�x{�Hxn��}��	�t	Um��m*��.�W����|�o�J�ѫR���؆��">�{�^>�H��(�+ƪ�n�5�vI#3�`(�2zv�F�2�ւ�@����!([��I��C-;�*�����H�)^F�<r�m����.'�ۆ�]�:�� �P�I��jy�	阁5U�^��Đ�s�d;i�c��[�e�����׼�\^��Kl��p���Jo#Z��1�"���	�|������I=�B詳w-�Q�9*��2�G
F�)޾�$����A]�i�]�9[�>��wi%o��ug�L�ځ6�����[��w nRwdH.�h"|n��p�ˁ���ꎷ	V=븄�=�@)&f%�.XGl��_e����ի3�~}weV�M�[vA�v� �n�����n���6H���u��wNw��.]�A�v��ʗ4Z��!�)����>�nS",V���������kц[�Y���=���ݷ~���e���ş�/͸����x��M��({tm����c� y�p�����<������8F��{"��g<=F�s����͹�p�]��<L��}�v��g��%����Ts�g�{d�p\v��hx��c[2���Җ�r���m�\����ġ��Q��tmv��ώ3���Gaw�:ݧs�2�M��1��������q��Ź�%�pg7`է�w	v�ton�����u;y�m<��~�����Z݋ڡ��ݻ'�}�� ���"���Q�'d�'+-��'o��>��ɉ���L
���*@�b�����m�]�,��N�m/I�}^@��7-�͙�ܲaf�<D��Q.Iwh}�����9��%	�iT��9Y��Ւ	��_m"|I����
��2�M��u�������=��6�W����w���2�S�{�r�-�S��{��a� M��D�u�>$��v��wq���WH�6�����5`�[��9y�& Xb��&b��z5��|�_��أ����q�差Hc/�vu-ƥKw���IR��,"�-��mā{���c�[d��L���X.�i��H�N�UG�W�Q��ivݐn���rx7�j��́�Xo93��o�~��ǽ��|5g����w(\�DN�c�;�޻�{Ծ��p�I-�9E)bQpȃ=VK� �Wx�O�c^D����$wJÀC����b�L�	g�Cq_,�P�,����&�����3��R�y�>7���ĉY�Dy7.`�rK�C�d���<��䗚�J)��yoR$7�]�$�l_l�<����U�������_o�EM@�%6D�F{�.�$��e�.�L�c�2�(?	۽vI##�eӲ��f�b#z��S{��Ǟ[2�n�K��!!$��y���a�cg��NnR�!�w���8�������zc�Z��όW*@��w��	�(��ܪܔ���(J#��n�g[2IR��,(8t��6�1Ҫ����y݂I�5
/:A�ݩ��#c��W,�ɴ��N��d��;ex�	5�����N�h�Tz�U��$!��2y	͝7�~[熔o�?l��w���)z�q3ϸ�O6/Y�ثƟd�$\^���������������犼���??���f�j
����O�:ŉ����$63vQ>$�v���Dn ��z�}�`��U5"����Es�>gc�n�;�;�$7���_l�H7�ԁ�������������-`�u8�}��Pmqۑ�9%�;c��ev�O�r&{�f�����߶�A����Y�ͽ�A �Π�mL� ���/�jnf"fgɴ���s�P��ޗ=)�����~쿔i{�P���s��2u�r���u�>�{䯲�-�����\ǒY��I|�+��q]F�M�X�}�}�� ���@Ύ]+ƥ9��}�S����BJT�M%�IwO����������p�A7l��@�ޙ4��yy�-�*��Z�@�qPc�j��{�eڸ're�?55�oiõn�'�1Wo>�� 	���v��~*BGș���g<��%����>�7���H؝R��gR �	��wk�/z77���	�m���cL�R����f���n;����Fs�ǖ��qL�9�������H�515�"+�B'�;I ^���g�u���Lv�@�o1�8h��"&	M8!�P�{�M'��#P냶y�@�k�p�z}�6��gw����/!36s���d���D��Nջ� 0�lҸ �J����.�,��� �Ղǻ�� ���@�S-����\�#�=SVw�G��N��� oy݄@$G���v I�.3۝}��s�� ';��p���"ځ��9��2}��W |ɦ}�>�����j�]��%pO���  �;&��#渚�^���?t�!+;��gި���/���X�<!I��O>~׾� �9�ɂ	D �����D�{P��P)��=����v;8���c �(9C6��6m�ѩy�֑Or��p�N�+�˯��-�nG�fsT/[ɛಊ�?u�Ӌ���?1_���6-s���}���פj�7ă���y�Hz��*���gi�ޮ��7��
a�<�T=��F=ؐ�R�4� ��N�.����5[��tZ:j�:�I�}�\��k���͈4gu/�Z�2D��W�{L��ݺ�Ӷ��>�,)��*:E �Bɽ��7j���2�n����٬��ˤ&q��q���iPgY�拍-jyz�vۋ�\ܺ���=��gQ4P+�;"��'NQ���(���i�"�?y�Gw�0˚�y搞w�&�ҶM��F���v��Ƕ��=Aq�-^�"����hG��pP˞�V����Y���%:|�N�6n�>��r����Jvxe�Z0�N��v]���7ة�䵻�˴p2�{�}��LB�؃[(���.��Lټ��x����s~��,�]��hO��O�x>���/�{�5
^�C�hM!}R�z�}���M�x���IBv��*�ۚ�x��Щ��t�z��܊)����xd��;���={;|f�l!�:f��_X����ܛĭ�P���{���/(���h��p�V]V�����R�H"[�Vď��Vr���(�����OĿo�����S�xEk�3��9?{�o���y�=�����$G
b#$��"#�EBb���D�������I�DV�Eʄ�Q1H�2���(����$�Q��B#�$b�EZ�TUl�HH�#H���Lq�fF@���GDQ�WD�J�WT*�U�pUX�d�G +�
Ԉ� ����-�,�8�� ���!1AČbD$���#�I�X"86G"�(���*(Ԉ8��Ɋ &(�FDEL����1#���$#�A�pU\DR!\qE�E�,����JF
�AE\l��d�S$� )2��-�$UEQI#�⨂�E1�"�FY0\U28�9+a���d�d�1�WU�TIY��Z�UU���Ő��TQ�G
��֍A�a�5�U�kZ��cƏ[5��u���l�5\�����O��3ѓ��7[�v4Z�]�i��nn6
����y�v�rF�9z6�Xѱإ�|���F�mm����b���˞�-�o>n9�ϱ��,�<Nc\Ş�:9ݒ+������*õ��'1nv�K�&kb�'^����j�{D�ٲe�lf���]��kc���
�mQ�z�vN����n��x�[]���8�Mj�Z��O?���dy���tsj�۲B�v��4�a��ng�㗲�Zۧ>U4�R������Վ�r����mŹ��'�q��B���m�h:[n}��
��4fe�-ľ�7c�6����9���k ���[�mY�Q�����>���&;'���+yR()1�-v�/��Ҽ��z��>�W@q͵�Hp[��s��7Y�l��9��c���m�^��@�4�����秓cn���n�M���͐���]����S�z�\�x����ga�穱�q�v4Rkvې^��M�q��z��o^%3ƺ[��ۑ�]�g�r��N6�>�0���ψ�c���vq��>7k�{ip-�g=����L���%�Z]�5�QU��B ƷZ���)���:�\A֛v�j�x�)�q|��7�s�~/��D����F2�V<�5ͩݮ����l��]�aۅ��ʍ��?5���aRШ���	ɵeH;6���_!�D��d8��׮��nk��蠭y���]U��N@�J�u�6�@f��3ıUh�����xM6n�,h�ח+műm ��ۓ����0	��Lp]r\A�I׳v�SOR�'I�v�����ܙ�懞��q��`��vݗ���ד>;j����x]h�pm�k>+��M��-ۓ��8������C���<��i���x�e ���d��4M<���c�{)��/)�f�V��X��{K��ϴ��Cqb���|>o����mM�i 6��cp�6m�=Y{��y�j��\#�d��X�KtCP��30�Nm��Z�Qѫ�tY8��8N˳{jT�(����m�&F:���P�+�$�A$iSE*�4���0unK�.���7�9{;g[����6��rG�<�s�ky�օ|#�W%z��qn\�{Tg�<�����}!ЗWL`��i>���Yw`���0$V{m���O/l
�n�%��<�{OO20'm.�8ὤ��-۳���v�0���KiQ��<�]�7mŞ�Y��s�63�#]�ԧ�ߗ��$p�Cz��ϵ�X {zn,>� �ɞɚ���G�<����m[����gM�>�j���r���휆7�Rpom�X��gM� 'd��Io���gk�&6{�M��HvGEcP��ۻ���M�@�_0ܯ{7���y�a`@q�髀H2Nɨa{�J�C�5-�L݄�MΞ8^�c�]o<���>e\�X|@3�3_ �}Ϋ�w��2z<&]Y����ũ�o�$�^�v�2ۙ�[e���>����p�#:r��~6M�%��� �7&��#�7���
R�G�v��=��̿�4K�"�]]x���p�c���V�V}���w\�m�_~�w�bw���\���nM�|��ܚ� �괔��<�68��L��SU�v	ɹ5$դ!\H�$��%�����gG?k۫�y�Ws�fz��&f�O*���M-tr,_��E���⧺'�ꔩʩÍn83�nP��3S�#��T���"">�rG�?���6g�L�$|{���� 3�����'�
no�s^��Ģ�1��iĎnɓve%P�k� +-F;���DmW��|@l��L@/o��W�gF�cPK7i�ze�9�zzװ�K�*j F~�0�8I���ב��$ x���K��r���-�9��t�`�7fdg�i��� ��뙠 ���w`��ݳI{�<�����<���s𡉌 �6�t���<����K�d<������������73��˞��u5 �s�� <wlՂ^]�[>o:����65H_NC��݁�/a�҇�q.l�2o�o� =9������'�a�$G��V� �==�7q�M^_ze���+��B����I�Kg9�XD wl�X|��Et߫gY�=ʏ!dV�y�W7�=�*v�Z4���0������]:��^}rG�r����Kݞno�mA�+8>������ �w"t{� -�ٟ��k�@���w ��zHr��p�G5'l�Љ��i*u뿬 '{f���o�=ꎼmh��v���j`�c�wp9��  87&�����ʺ���t� �7�j� �t�����6�[yI�Q�7�ݣ�{��k�V�M�vv�Qs�[��ӺG�7[\aɹ�~�B���-�9��[� 훱$�;&j y9ْg����>2svn�Ι���%�3��ʛ�:GS_1/j�� Q۔��� }���w D��J�ޙQ=/�����}E� ��P�N%͗��Mń ɔ����~�����7�o���7f� ��eTB�0H.PډR4�Xf_8ݎ��S�
u� i[�E� �4 }��{�2��{��r|S�̇q�^�&��b����Te\<�fa���Т`��q��M���f�T	��;7a�`�U��"��4g=sI�=��f}�<W�o���x7�����5��57�'l�K��]���V=Eң�U> d�Tw���Y��������G��Uz�8��]�olyg=eB5��W=p�L�13���JX���tz�n, �47&� }w�V�ޘ9y�Z�;^���ɲl��0�W�#��B���s#iK�H��� L<�'�8��{g�a @l�d� w��%a�EB�l'ܻm��{�O}0Kng�m�7��j������>|�sn��{� �$̙J����;�}&��%͗M�OW���5���� |ݞʴ�^;�kwr����e�q &��^f�H�RډR4�Xuf�� 4�ٸ�'!�=t��]�yj��D��w���B&D'!�	>?}ʈG�� ��f�x�&Jg�|p��� [�w��?�.�[/�z`\���ky=���-��)#��]����M)���ᠤ�"M���y{n���T��ﾈ�|� I\���5l���pnU6��zx�ۮuKs��ۤ���8�ja�q�V���L���6ٸ�wk�l�V�g�t"�\�����rλ݄.Kc���n�)Tk>D�i�u�[I��h�v�Nyq�x�+�㣏v"W�ͷ[`��@iy��m����vi�q�u���Wmson4�i{�W lV�t;���@]vݞ�nS�v�L�zڍ��wn�&�i���ݹ�n�E��Ԭ�i��]�Gl��l�i�>��>��Z��Z,��¡�T֯�l�x!�+�ʅr�T+���oxx�C��
�J�p��~׈x���W~�������@��)��+��=D#�l�������!"s���{�	j�Mּ6�����}�u�8�2�Z�P�m��������<ȩ��
�ȁ3�
�
�~����!"8�B�D���\C�qʅr�P�v����OwO&X�;��@�O���	����]in��p��+����8<B�D"e�+����x�������.��|_wϹ;Ҡl8�c���{�\�	��~�Xx�/���M�d%���L��E�I�bl���W+�
���og�2!��
�~��o�qÃP��T˖�w�(�U�KGΦ�X�A�}$zL��y���xq8%L�I�~/2ɬ�.��*q+�y�u�8+���
XeF���U�D	co�LG�쁣̀����V����B&D"dB9�N����s�T+�r�S"{o���	�$�e��/�V�M�5�N��E&���
s�ymѳ���K�l�"c�����n����k9���V{[�%lӮ���j���{��"g,
�K�}����2<r�T��2��Z��&i<�W>�����29��;���C�P�P�a�~�\C�0p�V���K��԰���^aP�pB��}��&i��n��|�~S�џLf[eS����Ԝ�8�ǒ���W�w��П+��ܰNRP�]4\u�Ogo��1{jY�)4���m��D�3?��W����9�*dB!A*�����*p�5
�Z�L����B���H��G��\a8>���Or�������8�%L�C�y=Մ��N�k^L�q+���wu#�jeB�eN�����mHeB�p�U��[��>�_?a�"pB�R�T+�>�}�u&D"dB!�J���ݚC�6�p��߽SZ֫]in��L�F�~oa��}ޓ�O�w�οD6���S)`W�kϷ^q2�ʙR�Tʔ���L�x�2�#�󿻽��'�|y��|�p��DȄ�a�o�n�ǎ
���f�섺֭�u��8���T�W~l�x�ЮPr�\��
����xx�B]O�9����<B��
�M�����5
�Z�L�����f�4�L��T��+Ͽw{É�*eM�xy�߰�U�2H��?"\�&`H���b�<�λ!��㞹y��t�<��:獏����d�[��\���L�G���ۮw&W(�ʅ������^͡l2�Z�P��w�0���$	# }\�ol�m$�[���C�?9P�QʅB�N��ݚC��óo�Y��Z�,ӭ��L�G��H���� A�'��AA8�ON޾����+\��(�2������i3HD�����󿻽��9a�	a��?t�g��n���z�¡[u��r麺e$��
�"[~�f��ChW(9P�Pr�_����q�!S"�P��=��z�oN?�><��1�ם����u��鋖Gآ~��#�C�6���32���Ƣ�9kd���2�U�d�sn��0+}��gN�{� �}���T?85
���=����g��S#\����y���{É�J�R�����V��tCZ��g������o��qJ��i��2G��3�C���i3HDȄ|*����xx�N!P�P�W��~�C�?yy�糵���i&D"J���6ihW
~�����kZհ֖��!�5
��9��1�2�S.X��u߷^9��߼���}iJ��Q$zH�]U�#�G�S+�jer�y��w�8��K�ʅ�����ۨq��P�>7?s����?Q�-����o���ùx�.�ONu�L��>����ɍ����/������pԾn���i:�Oڻ�f��6�r�P�W*���og8�B�P�PJ�p��w��<p�P��s�w�~C��l<��vi3HD���L��}�����S*Ro�Z�Id�MWWÉ�8%p�����8�2�Z�P������y�l��"}o{�^�6��2�Z�P������B&D"dB9�?}����"�T*�g�s���w�ԟ_l�M�\)˷꼖�kR��u��j��~�Ï����w]�u�L���(�2�ݿo�v^�����?w�I�B&G?S*�߽���a���a�����8�p�V���K���ut�I5�'��^��H�[j���i���B�qʅy�{���T*dB8w��ۨx��j@�=>�����9Yξ�Tn-��2�k�~�����+�$�=om���f��,����R���=ɮ�,��7H'�߄���lv?}�o��}�y��T�S�}�k�0�&G�ʙZ�{�﷼8�L����{uiIlՒ:׆�8��o�|�����L�Dȝ��vj�y%���:�C��zP>@�'7�<�!�
�B�\��{���s��
�r�P�S�^��Hy��+�����^�]�磯m�l�Ц���ه�ݼ�ti޻NgV��8���e돞������Y�ՓN�u��8��B���Ã�*e�S,
���~ޞq2�ʙR�S*{o}٤�'�T���������o�ɟ9�5�?s{Èr�*�*�������<p�V��f�섺֭�u��8���T��٤���9P�k�:�?{����>{ϻ���
%B�q*÷߾ސ�À�+��L���ݚL�2>�2����?H�י�w����|�2����^i,�ɪ��q2�0J�������+����S���f��fд�T+G
�{���p�����y�B'��B�B�\�~׽�zC�qʅr�P�Q*{��vihW۷Ҝ��WV��u��2@��� :*
�������F[�n�����s���TʄL����f�4�%L�V�W+^����!�y��t���2!<�k\���<p�V�^�_�)���U���Hq8!SZ�}�I�B�\�TȄ{�ﷳ�q
�i�}����q��*÷~�zC�5
�F�S)a�����g��24���W�ߵ�����L������w���^���w�F�t�l�Rg��̩T02Ne�y�$�fD�M���:�Oj!����n�=�Ɖ�U�<ܣ����N��^��w�OW��4�u�O�����|;��p����?�>�8��|��x���L�L���Oo�3u>�j�r��]�+�7i��n� ==i�v��.���3�uq��#����Cƈ����	^SgW㎝��^�8�k-���Iד!u>7v�[��a4]h�i����D�Qh�㛲g��gv��K��]���Ƿ� ǚ�m�s�{��.��a�nۦ�v�}���Q��ˇ>��h�v����P���}�w�����5���=B8j�Ϸ�<L��jeB&D�߽ٯ!�B�eB�*�~������$�$EZ}�s�w�s����������
�r�P��;���4���B�_~�ӑ���Z�N�u���^��oaǈTȄL��&�5x�ﾆ�'�o���9���*eJ�2�>ֻ4�bT��jer�_�~������ C�MAs=�q���;��D=�
���_�Y5�S,ѭ��NT�_<ٴ�!�r�S"����xx�C�P�Q*�~����~xw[��߾���C��p��*e,/��vm3�����9S+G+������pJ�R�<{S�F�e�u|8�S�\/�w����8���M� A��"*SA4��P���{��<ÈD��BH� �A�|� a�Z�����=� RdB!�*_��l�&Ю�zS��ն��u��j�}��ǈT˖L�`W	���{C�Ȳ�瓾~�޾���>ʙ�2%/����4�	S+�jeB=����!��*�ʅ��N~��J#�>@�~��X<y��J[�ݮ��n8x�Tq�F���o=�=[@�)s�b6��K�}��r���eX��4���*]^�f���\�T+�r�^�����9�*J�B�B�R��}�hqÌ�$�_V�Q���w�@�=sz~�������L�r�~������2��}��STe�U�k^L�s�]���h,�A�]�^�ꬃ�����תf��޾�ޝ�n������Oc��q���ޞ�7w<f����|D]��r��^Фˀ^H�9*`\l)����g��%���N[�ݚ�fз!�
���y�B'**
�Ŀ�������W+�
��?y������EN�G������2L���TEF��!�B������������������&V�S*T��<��}��w�Ɠ4�	S*29F�����C��T%�T-�a}߷�8�p�V����H�]�u]y��s�ڛ�(�gk�:�������| Q����{=s�T.%B�D#���{��C�jB�R��^��I���_��pWS�8�A�}$zL�I���1���?�p��Yu]_&T�����=�������P��T�o}ٯ�.�w?g)w�_��L�z�*����a�"q
�K�T+��߾�����
��T.%Ou{��!�m{�������5}GA��f��mr7O.{2u�pn9����ݱ��'Nܢ�f���ߜ��n�e��N��ø5
������T�`T�`W	�{���s���Tʕ*eK��|4����W/�q�����7~�ݦm�Z���oxq���T-Ʌ�}��ǃ�B�.�zsW)�ji�c�0�N�Mj��O6�r���'չCb����ʙ�2���C���(\J�B�B�_u�����p�B�D����I��S#Aʙ_�pS�����Q�z��!�$zH��g&�)e�Udּ4���W���zs��2�Z�P��T�{�I�BxC*���$��!�]�u];�K\䗡�Ab\z$��*e�I��ƌ��˫Ѕ*��;ͫ�=�gymۥ��*V��a�����q�$l�����/���Ixr#;R��K���$d{����X�hs� �4�6<^�d��
㷸�W � 4��W���?�iC<p����.�N-܇}0�L<i���ݣʽn����s�g�aa��j�'s/U+�5+ܲ*J�,�1��
R@z�n;w���t�wo���|��Z<55�{z�n��e��X�nݜӰ�ISf��}�d�v��ـg��n�_E�%M(�b�E
���1밌�NZ�5�`�zV����v(m�>=�o3/�Խf�Wڽ�Okׇ6�b���=�ZXN��HRӮ��Z�}��<��d��V������[z�⏜]�W���#�з�ᶽ��|ڜ���k�'�K��wj��x@w�>͘�4@93��o�:t���ǽ�~���J:^�]��=k�l[ �n��!r��������v��~��:�7;�5z�Bv�O�؁�g��mx�l�n�����
]c]����?V��q�N�w��ᚫ�a��W�ȁ�T���4��c;�����R���u�]��{���{�VD4+3w�J��i��7�Vy�������EG`���;(���/��"�_,S��ܢ����\���B�O�=�؎��^��tӉ�N:��<FVX͔��H��"�:I�
�dETTk�1qm�!
�k��TXF
%��H�ڒA��W$�c�E�VH"6FZT*W*�qEQQUK�#I�$+�I�Z�%�El��"��Q$��\j�U$"�r*#�*$H���E�Zb"���f�\�	
�Y�Q\�B*)X���Yl�+ek$c
�UbȠ�-���)UrȮ.*"��6a+TA\W�JF1�#V��*�YD���B���Gq,�k\e�2�-l*U��H�$A�Q��H8�&2"I1E,��8���.-m��F&9H̆X	(�L���(�����BU�f*(�0�DR�U�?�}���?!�B�R�P�T����oHq�9P�\r�P�T�W�ݚC���}��ژ����Pf��|0$	5��@=ե��t=:~����& �=3 I�R��O1�&T"dK�S*^�^���'�S+��W+^w�w�8��|��ߝO�z��2�i0�[���<*�ν��E���˪��8���Tl�x�ЮW*��B�������!P�Z�>��u�C�J�p���w�!�Ȅp�P����_}٤�!#�9S+q�󿻽��"dG|���������&�����G-�O*�c��]q�q�q�Cq�[��.�k�;�]Y]~��j���.����ʝĮ��=ޜ�����T)a�?[��5�C6��ʅh�P��w�|�!� IH�'~9�f��y}< a��6���!�8�B�pr�P�%N����&i���o�5��jY	4��!8�)v�H8@�=3 I?Z��R�~�����r��oHx�Õ2��T���}��f�ĩ���;���!��"G�zH�x��mg@��{����¡[�_w�Eֵ4�1טi'��^��I�!�*dB&D#�����9�*dB!R�\'�v'���y���!�dB8~�L�a�W���g��S#\���W����'�T�{���Y�bb�`���a����Q�`|�A�y�o���g�652�K��y��&i	�2�Z
����a�"pB�R�P�\O��~ސ㝷^w�_^M{��?�^�Cx��Nt�s�:���I��xL~&[a� ��'��#g���y�/�����=����������đ�\�0�Ӛ���94�>����H@�$�sYP�E��+�vr�L���Jb�zC��]w�oaǈT�X2�'����>�=&�N����2=� D��7�s���4�%L�Q���5翻���8P�P�&��~ސ�dA�ʈ#�~��jH�	>�RE�x��!��l����g���TԺI�&j� 4�7�~��E�Zԙu�]Èi2'��{4�ChW(�B�\�W����q�!P�P��>6����|0�O�{rO���T>���*g�j���&y�2!#A������N%L�C��گu�U���eNWu�}ޜ��2�"׾���O�Ig�|��|ٯr�*dB4p�V�w�|�!�
�
�r��]���s�T+��T5w�[�ǿo��/��l�&Ю��[��d$ӭ��p��+���{�*e�*dB8}�w�׀�+\��.	S*y=��Y����S��Ͻ�zi3HDȄL�G�y����zXeBP�T-&��~�C�
�m��:�]i֥�5<�Hq2&���4����{�ٯ+��P�o�W+�
�w{8���������*p�5
�Z�L���ݚL�������3�zG����}�xq8�2����q���,ձu��q9�\7��q�er�L�Dȝ��v*�y&�.�mPK�(�DX>@��s���8�N
�B�\����ۨq�9P�QʅB�Ou{��&i�#�>���������}%�J�c՚Eo��R�~�S|CT����r���IحN�F�柲i�5[�I�sy�dĺ|�]1�R�V �SہK��s�������^�֮zt�������ط�v|�^ʱ�L�9�1���uǳ;�ق�oOo��͝�o3��R�3[K睎���;�lr�a�g�.8��A�n-A���{]���<x�]���K�҅�*����re�A��V��[h�y_<,[] s��=����T�y����ۀn.��a�t�o@μpqf�Vێ�n{v9����\vw0����b���f��8rng_>�w�.�uu�%�t���
��9���3�`TȄp��w�׎q2�r�T��2��Z�L�x%L�=w��N:վ���s�]~�w�8��DȄ�}�~�C�
�iν��A��ՙu�^a�4�B�u|�f�4�s�*�qc>������Co��w����T�T(%B�_��yP��L�D�a���P�� A�ՙ1~ݫj]�Q�������*eK��m�#��)�����ʜ�y���s��2�q��a�?[�vk�fд�T+G
�tn����]%����a�>�T��B�S���ۨq��
��T.%Ou{��!��B�v���SSR�I�[����}���a�'�����6��`T�`Ww\����&T"dJ�2��{��&i<J�\����������߻�;{���O��ʄL�Gk\��=�¡[}�:�Zue�5<�Hq8!Sz��f��ChW+�
�r�_����ps�T=��Ϝ�>��D8�ĨWw^su85
�����_�٤�!#�9S+G+������S*^~&��m�ܦ�|�� 8�ܹj$�@ѻ6�)������,T��Ip����}�~�g���ֺm3���}�;��&W(�ʅ�ʟ[��5�3h[�V�T+s�w�<ÈD��B����_��W>����wP�r�\��B�R�u~�f��hW���xK�kWU��]y�8�ơ]w��Ø�
�l
�����Y�Q>^)S8�jf2l�"�Q0���ݹ�����>�-��7K�V���݆��=�/�X��ͧ	�럫�����59�lՄ��2~��M�/ÜL�r�T"dK�Z��&i<�W+S+��;�w�8��K�_�o�g��vs�j�$?�$	3��-՚֦]iטq'����l�x!�*dB9G*�����s�T(�	#�@���MZ�����eW���!��T�a��g��27����{����2�9w�g$�,Ҏ��X�=$a|���꛳u�g�W�4~���9֦T"dO����xC6�L�F�B����!�
�
�O����$>����4��Ͻ�#�A"v��l�	�+��7�Mf����M:�DȄ{�����T�X2�\>����8�]x���U�����<L��J�R�k\��I�O���L�V���w�8�L�Nd2�hL?}����
����~|��9�&�֤���X���j�=���s-�}l�8Ρ�ϭ�<��u���}u�WUԚ��~�Hz�B��}�f��6�r�P�Qʅ}�����!P�P�T�W����*p��+�埼��t_�;����"Oo�m3HD��9S+\�߾�{É�*eJ{����]h���.���!5�y��=x�\�OI���9Q]<ȏ�5G��@��%2!��w�<B'�T��B�D�����8�*��B�|.���{��Fup$%9���"��~6"h�Tԛ�%��j����x�L�`T˖p��w�׃�L�r�T��2�靏�һON^��ԏ�6�or2!"Kث�HzjE�L[����b�n~�����uw�;HjM�U9Yp�y}�y��:m3I�J�\�L�Pk������8P�!�I��߷P��¡[�����Y�je֝y��pB����ͦ�}�?|o��!�r�\�T+��~�����S"����C��p��*e���}ٴ��6o�����O�i��9S+G+�߿oxq8�2���m��h�J:ө��ʜJ������9�+��P��'��vo�fз�';?~���;*����B'�T��B�~���9�*�� I�#g� X!$��Q�k�!�������g�n�lR��eź���s��\ u7k�f�U��ۗ�߿w߽y#\��k��:�+�ϻ��1�2�L�`W������&V�TʔJ�R����Dz��D��>�f�+�����{��O�~�{Èp�ʄ�2�i��}�u<*���~�mt]3T�O�i'1
�w�l�xm
�r�\������_�}�C��;��z��T�TȄp��w��L�GP��'��vm3�p��2��Iؾ1�q�#*#���\���=N�Tʞ���ɩ��V�ֶm3�#��|�􇉑���ʓ���7�3hZC*�
��������u���k��_��������B�\��׽�zC�pr�\�T**_׾��bm
�}����t�j�VK�4�"��� ք�zlJT}O�G�� I�÷�~ޞq2�ʙP��-�_{��'�T��ƦW(ם��Ba�?F�_m>�/M�SN�}&���̲�c&"$��]��Y]tX� 썕5<V�ܺ�c!��8AF���)	���m	��ZL;����L�G�������u�L�ѯ0�Nb/��6m<ChW+�
������8��}ѓ�ϔ;�$G������]0�g��W
5
�~��f�4�L���L��+���a�<L�����Z�}�u�8���rs;��t��%|��]�:����ѣsZg�{�������=ծ�٥i���eN�\;�=�zs�+��P�a�'��vo�fз!�
�
�i�����8��T����ֿK�ٮ߽�-��oHx�1ʅr�T*J���vm�o^zk,�t5f�y�#��W�;����&R���w��sF�p��oO�q2�ʙR�L�K�]��i�B&G<jer��{���C*�*	�e>�������Dxᱵ�&�ɢ�MR�>a��K=�A�9�r9�r8s�h��	����Ͻ���v���w������5
�l/o���g��S#qʙZ�y���8���)��xcb�i̤��(�� _C�������m<��J��3�~jeB�a�'/~ٿ!�B�P�*������8�B�R�
�O��~ސ�{�}c?k���:�:��"R����͡�m
�Lwg%���&�%�Q_G�R�%>��!��`TȄp��߷���+����sI����#�=$H�Yv�<J�P���5����8�C*�� I���Q�	 I���sB�S%�o.���#2���~��o����򾆓��P����l/�a�!������O|��J1Rk��G�t ����rV�=�vȽA�fthJ�=����v3�|���8�3�8�p��En���t�,�F#���Fu{a��8�uK�vzRs�.��{v:�	��]p�Nk�bһ�� �b����9�0=���e;K1��q�˛����x�z��>u�7�R�Q�5�l�ysڃ������㷶�ܭ�ڻn.5݃��#��Į��n5�6�:�"��8�	=�3��ݞ�h;�OZ��w/glb��9���~~�x�G���{��b/��6�!�+�ʅL�G�~�{89�**
�
�O��~� a�i�ܱ�b`N�b�xnL�D�������xq8%L��]�0cjA!�*-GҢ�l�즾ߗ���H2G�����GG��"z�yV���ma�
�¡[�~��0�8�B��W*~�{���
�r�I���?>0w�,��M����@��ߓ�Df��)�k�!85
��}��!S"2�\>�����8�Z�L�Dț�~/���t��5���4�J�\��ʄ{��!��*�*����oHx������E�9�����(�P9������^Y�4��T+�ʅ}����8�L�D(�
�s����i8pjB�D��}ٴ�5����w�8�9S+\�^�^F$�Ivt��&f�H�Uf�8�Į�y����ʄL�P�zH��h+<�����׬{G��?y���a�"s�T�
��_w��&D#�r�P�T��}ٴ<����>�������IN��I�%�ubrtcmǌ%�g��sg0��N��Bu��6����'�Y<*���A����������$���aǈT�X2��\;}�����&T"dJ%L�?^��i�O���~�"~�z:)|G�����^@Ɂ� D�*�;����8T+��߮�:�Z��]�!���K��͛O6�L� _n��z{��7;������^�#��V�65�ſl�yM�N����[����{�=��N�9Zb`�Y��Yy�[�t���g�^@��� J*������4�8�+��L���{�ͦi���������w￱g}�{���%L�s�}�f�պ�4jxq2�+����w�8�2�F�T"dI��ݛ��-!�
�*�??���������D�
�J!P������
���'��vm3HG3���De���i�8�p�5K�y "���O8��u��L$z��w�ޞq2���(�2�/�{��4�%L�Q���ןw�� �=���MN�&��ra�s�ސ�dB<�߼]6�7Rj�i�!��!R���ͧ�B�qʅr�T+�����s�T?z����_�O������P���w�<p�P�j2$��ݛL��
�T����������%L�*�_��W�B�A�s2�,��[M��[�u�+�9�{^�e��]��������P�������}�[t�ֺm3���z���Hx��S*2$���ͦi	�2�Z8T+y���q�B�R�q�m�_���s��
�r�P��/����f��{��W���j��i���!�5
���{���';9߿2����p������d~*eB&D�����f�����\�^w��xqXe@��� L�Y�-G���;�H���|%
���_:�Z��]�!���K��͛O6�r�P�Qʅ}���g8�B�T*dB8~�N���v��w���ϑ���k������ ��ǒ�Ux���nQ�����^w:�kޡ����V���2��ѣl�������9Τ|�{�y�5��}�����jB�D�^��i��S#G*eh�y������Tʗ9w��jM[�`�F��*a|%��#��W���o�>���,2��w�����*�
��}�����T��B�R��~����\�9���8��|�B�q*^^��hx&Ю;|��KlҷM5��j���oa��2!"�}���p����<��8��#̎"H��"j���i<J�\�S*��}���XeB\�T-�_����y�
�>��_��nT��^��#P��6ē�K/d��ׯ<&���u�XI:Ӟ�t����~�v�ef�&��?'D*]��f��6�L�G(�B�����s�T.%B�D#�����m&D#�y������F���[�6m3�25ʙZ9_߻����Tʔ��'�5���L�Mk�i�NbW��ۜ���52�������;����^sf��fжP������xx�NT*dB9A/����&D#��*w^������O9u��C�m
�O����]j��i���!�`�+�>��x�L�L�`W	��{C�����.%L���W������o�7�?L�z%L�Q����������9�P�P������p�w��MD�N[��.��qTͪ�~��Kw+ ��q`�����K�c}�vj�L���S��d%B2Eom!�(V)=w�rg/��$�)�l�����Ǝ�;���1k�N�v�\��6�1w��ֲ�[~���L�u� }���u�c2� C�Y��`����;5^}�c�L@�˫W ��u ��c�fUu׳�
�&!�O1�>�h��ٚ�y�C�-s���fg���-�;��K��f���2H���KD=In�X@��w`	-;�?Ur��Lh�Mz�{�D gv���uW�)nT�˘����!�e׮�š��n���n����N�)W��q��i�[��6)��jZ�m�S��,I%��P��y35���]Q�ܳ��\Ƿ�݀	i��!��l*��62G$�t�=Oʢ�啞��Mv;��H2{�Aw���o��ܮ�w$�Us��>�Z�p��Ԧ�ù�*�C���;�fʞ�zE�|T_� ��u�� | q��� ���U��ʶ�\�Ϋ��~��Fl��<b����C�o��`��=W)�$�ux���.M�r�ZL�������~��}]���/�rn$iɇ��wtH�OE\X�N��������nK����LVS�9!��9�p��m�˃�
�
�1����vs�O�Wcvi��qK}P�@����!��k�g����`N&]�\��A;y�����a�ˬ���%�����m���x�v�(E�v�u]���O�����^����G��\5$9c�󻐃2wy输���Y�q�����ӵ���x��o�e���xz	T9뾧	����L����巩#g���7o��X1����8� �&���=*P�^�Km���'�Q������ˉ�U,SVe��M�����p!I��+���4��-��� �VV������i����՜��=�1S�+O�~p<��㮮�6�X:�}�ǡ� {�����740�$T��lU�^R�a�8�2Lc�3WN���!��M���zph��;v�l��:����:V-1Ḵ�s��|��Z�{;�s��Ȃk�R~ܖ�Y����,Į=����Z0��gƼ3��keѮ��u�t���>�M4�yt>�һv���d���hI�&p9WUd�Ҕ'5�=����y�ڕ�ڀ�M��e���2�0n�K�4�����qK~�͹9�k�ϟ��|��9l^�!��!���S���Ljۂ#�(4.Ɂ��Nr��Fd��a*�.JCP�otUVh�Ҫe��מ>����`����
L\I2��(�aJd�8*V���Ԍ\.I"�G
�	��WU$$Lb�ɎLF5+�q�%��DQX̰�$��E�#�c\ȑ%��TQ$## ��9�PG�eTWԖłL�hR@UG
��T�#���b�(�\+K0$��S+ldQdJ�bBB�$���(��-I$bG�@�@��[Q�2
��$�D$��-�U�+���@�!E0�GF�DQp��2,e�Yh�q�)AI�ĎG20H�F�DUn@GbRL�.�(D���ȫ�$��*�"��ɀ�LR
�B�Ȋdc��̊0�)dV(�X��\,����,�S������|���e�����O\T֕:�8@ҝ�'Xܮ�u��z���`�t��F�<�%D�CK7V39��Ri-�����\��S\�[�R.͆ק/��j��5q��vy,x�x�	��k�`�c�y���c#7g;q�֕b^e�r�c��w�|D�&h��n8Y�H���Dn��^�i�D6Mv�;|�p�K밝����oG\�حɧs��ƃ���S�ԛm`5��]6n�vu�lW�a���bi�s�멱��by:w��ng�rvѼ�n� һ!WYyy�=�� ��>��0F�z{x�{N��v磷F�KH�a:a-뀛�����b+���uݶ,�kd��P'(j�s�im���<�^@����x=��ݜ��'n�5�yƧ���	�N�g۲yh�c���K�nͫ��;�]��P�("�uˇIb:S�8}x��ݻ�/gu��5�q�	g��[m�����cxs�"=�v���uV�΄/W��gq���n�I�P�y�ݵ�^�k�[������|�s�
�9�*���G�������q���x�7���Ͳ�8Y֫����h��8�u���z]c��kSM�O^�[�S�<6�v�`\��-�.�lD���k��/t�����4��nA��a�N��t�ۭ�خ��e�gs�x1���s��Sl'6͍��80����7<��y�JՆ�
W��x\�v�;Z��T����S��{H6{q�J����[
���S/�	��[l�#�",�嵳�y�y�:��ѷ.Bk������/A;]\��Q<%��^}�ו[�F�8���vv.�tv5��#�h��[�A�{n(�C��v�9M�O��ݨ�5q2x�1e:�Xα':��s�1�\;��ʶ��m�tv�n|��n���kq�ٺ�#0�÷��=��v����ӌ7�vpL�ۀ�|O�����'K��3���hx9�Q��<m��1��tt�d��;'����K�KBڗŚ<�x+����a�e�x���'m�g[p�8�5����r� �G�0t�Њk֍WK�b�<kM���u��ti�u�x1�/����kX�휙
�c�^��.$�l���vV5dK��3���s�@�������C^vȹ�ƎMЂ{n�w�*�k�Px�={`�0p0�D�Y'�ݹ��`����B*�&����Q�nGrn�8�^c"j2�q.�)����Fe�|�V��/�@���}�j�)�2��-�T��]��"-30�����ID��jaڰ��:W �}�{8�o^��� �q�| ���^��N4�or���@�½*F�2K�CE�;\��ל�," j��������G���b .���~�6-���9�nn�_>���b7��e�� ���|� "�z�_��{{]��7��o4��p�'��0��V&�4ڑ�2������%����B�=�7&&�A-�(�:�z�"D�{�]��Q^������/�wxd9p�����F�����p�1ڱ�u��.�U�ʤt,\i�o?z{�	6ӑ�p�z�i�� ��ˋ���Ε��X[����5ꈬ��& z�9w%��H��d�Æ��2�ͲI��_/x�g�h�s:X�{�ۻR�����0�{�(?��QU�ՙb�db�7��^�m�!U��X#�߳4��8I��y�@���VJ��0SKzi�H+�֜�(��mL;W�ӗ)$��]+�-Otqx�}9'�lK~���� ������ey�4��ܒ9-)�ץgOg�O�)��]��뻀> 7�k5��+����c9.�1{9po��J��q-8s ���>�wa��q�I���\K�26+����Ē���݀	oN:����z�u�Y�p$9��v��N&��;�rpDq��7b.�t�Ós:��\&�Sm�e�$K�Q�G��;]� @�M%2��U]������{���D@{�]����i�M��j\;���ү�c�ښ�){nj�� �;u�W����$�Ӭ6;�feg�ޜ�_�e��0r�J��v_���w`�ct ��ՓU�ڮ�s��b�חI6�-��$`f���;Fy>$ߝ2 ņ���'�Ot�e�}��K���;_`걡j��f�S� �{]_�| ocu -��9�Q-Bm�%�w�e7�՛~W]����)��"]�ԯ��Q����IW�%}%Ӕ��.fG%w��[� ���5Es:WF]f�s �3]%`@w���D�7�ٗ�5^{��as�66/L����[h x}�C�=�D�U襧 zK�d��߲V�C�i���t��qa� ���U ]��,j�~s�������9����u��م����@�n�'��r�3X{ֲ&��חwk�#���U ]���X.q�܊��U�9���~���$�NF�ù��M� ~���	���R�]�t��׉{�>{�|
離����ˑ9l%@�.z�ת���u�w���IUct	��%`|f��'��N�qn�^lP��<[�s�n+�FE�iPi�l�uBԅ��ɹu�V���aܪ�	��*���"�L�r���Z�<T����K���s�c���Z��!ڰ����� |w�Ҥ��g$��ȱ�� �s��| �N]Ȉ ��v�%���O@]E��n[�M�J�r�v�c��æ�t����q)�V�kT�#n��ܟ{�ƛM�eK����| ��ۋ� ok�Μ�x���ڟ|��@#�_OX��e�l�Àp77`���X@j�;�ߩB��_�z�� |e��� ��݂O_M{s׹�ý���^�p&��7v�n�� gk���	�]���rl}s�%� ]�r�D����wa���ӄ���Z��.r��#]���s9m���.  ��wp ӎ�*��5�M��W�7WYzM̦�	P�7b\��,�95&�ꌝ��Üdm���q  {7]�����5�:/ۏ�_qp��{P��q6krvn�E�K��C�6�b^�ޑ�gJ�I������I����o�E������,�/}"ʧ39�������k�,vv�'�ۜH�>�O�=bn�S�͍f��p����'m���Mًԗ2ۊlķI�k�cj{u붽�võ��u�3�^��Y�r�n���һV�&���zL�l&kWW���v�{[��1=�َ�I���2����XxjR�L��a�e윽�z��T��睍���iy{�����[5v���g�;��g�uA�:�ݺ��ح�(��x����z"��]��9���K<Hۗ10����c����B�?/����,�ov��� ٞɚ��g�r1��9w�H�>=����+��6Ɯʗ3W��횆%�ϥB�Ś�_WM�p v봒�6Nɨb ;�^~-Ů���gwyM��Ĵ���Þ��IXpnM0���$&y�-ӽ�G��Nv��A�vM}#w2n�N\ ��	}7�8��{"�.*���&]l�X GL�L�@w�֭r�9��~����(��j��b��%.�j\;���� ~���\�L��ȝ$�̀6z�n�>:Lɨ�" �溺]G�/�{�0����	ăp53.�b���N�r�:���vG=sk v[����c���~}W�6�JjIx���݄ ɨ`wϬ�����}V�7��������5�]Ym��2�1-���3==~��D=���o����!$��'b�RoY�z�^�d����8&�o��z�Q�Ll��8Rqs�1�K{�C��(D��Q*�ݞ�Hٝɚ� ���� 2L����d����a&^����ݹ�T�����Ԅ�z�v�� ����F磽[n�4 ���Ԉ��OU�}��)���Ď��s��#f�Kk��[p�F�� >�N� �y�ʞ+:ݞǂ"d۩%�ٱBK�#wa/f�� 0�ٿ���YJ/lI�NV@$A����� N�����.WC���#z�~�J	RԄȜJ�W>lK��9�b����F�n�)�v�d��:��{�p��n[�p���5 D ~����==�6��O���.�ɳ�s_]�r�B����6�JjIv���M���;:=�i��-� "�Ϭ�H��l��%���I�ҽv�.]Y6�[�!ڰ���ܐ i��q` LC�Vh��u�q^��Cv�r��L.�7=P!�b7�CQhl�F�t��Q�w�lJP6
�0rT�ɳCe��$ b�ٽz�2v���W@~���� z{�m+�kW336��ӆ2n�=�vi�礹�� ���� >����� ����v_�ۿS\ ���q!��i��-�ķ6�}ӑ` q��s})�5ө^�� ���쿀�On����c����mS�^l��R�.�N�pm�Ͷ��i�ܯ��뛴�8cn����s�����	hCp��M����t%pv�݇�@=�*��u����y��}^�D|�wf���Ci�m�m:�:j��Di'<��+�¼s.#��*�a�s@�	�S��Z��Μ�R˙����)�%����c� ���Zd
f���Kޛ�6s�n��s�sٷ$��Ȗ�Նa�j���ƪ���� 3of�p�6U� ������<ۼ�tc��f_:7my�O��=�`$�=�ع�1�Z�o��K#o�8��V���Z��Ɵ#ެ?rz�Y�Wy��%�DϷf�4Ȳ�(n\L1�W��5 @�;n�d��{�+�=]5`t�������훓+��{�~m��f�Y��nݣ���m968�Ɲ����d5i�˳�C%��߿��h�*��?�x��Q$���N�Eܾ�'��Y�2�W�sѓ��w ���� ��ɸ%��H��K:�R��b���/���{&�Ā{��� .�� %z���z�{w�齀��i��m�i��:n�,��v�>��{����2�r >�7@��.��{>����2��]�6z�5��w�3� ���� � ��͹J�2w�l���nU�Ը �� �ϦܒKc"[D;In����ٸ�R7Qq��5��]-��]��f\�gv����5Q==�z&�aZ�E��UY�h�laQ-f�owU�;X�0�P���uL-��%���`�b���4�J��9Qn�o��^��p�����&����3�6ܫ��m�v�^ �tە�-��ۇ�m�a��A;rxRR���9c�ka��J��{\d������v|2O��0Q�F�:^��n��&��<u�Y��s�t���n�s����^�st�cO�]�7l�@sõx�1=���%�nܡ�����燘����9u��ۅݻ�lo����׬
k����f�Ȏz��Z�j8�Z�mpJdM�kk ���9�
��w:�!/V�������K�r�ˉ�2}��t �;jR��gv�����y�jړ��n� A�nܫ��L�LlM�LK���u��,K�[��V:bɦ� l�RM���Ε� ���2z�_8���{ٸ%��H�����$����  3��:*.Cţ�2�m$��f����� ���Lq ��m�;�t���~ff�����:����{;]�����7o{Y�d�TO8�6n�7��w�d��	�7P�6�V���~���=�7� ��w� ����
�:��*u���%>��v���q\+=]leu��k�.sɺx`�ٱ�]	�T�8	CD�{u���nSR�!���=�m#��{f���> �u5A3=E���̓�eܥ`GNn��{Ejܡˉhs7p9�� #r�๺5.a]GT����<��Æ�ⷞ\����J\{eYӽ��L�f+}(|o�+^��Q/SN�����lW�hH�p<)~�W]�� Dd��݁��m%_�s�s��޺f�q��1���5hT��n��t�X�.���P��5�f�N{��} ��5`D����2j�D�s#u�}:�&�g����G{4�� �[IP�]�r�2(j��{�7`G_e&8�p�p�sp麀HW�]k���8�e�\�n�  7�� ��{�Q9�&}���Ӱ@�W�A0��,�M�����紜��^�&zՠz�4�٧.��;_~���4�)�%��ӷ� ���	^����u2����� ;��@^��&[�d��v� 1ge��;�����\z�}b@��� Aj��ℑ��ǊOLվ��s 7�j����n�st �y�@�9��k��T-�U�r%����&�0�`�M��(�9h�Rwa+�P�
c��9ykR����an���I����n�l	�}�Ky;��+M~�v�C*����s��L�ЏP���-�J�ǩ^��Cvv�s�l��/�
�N�F��~�ܢ���b�.�\N	����n��\��([x�\�S:x�ŶS2�=���p'�Ì�p��2x�g�Q��K��z����[�{Mp�3�+�������>�ݚ{Ɨ�H7�T���X��(k�0^�cD�,YUV��%C{Z�I���f<�4{=�4��s�q~�=|�]`[[�ge3�&<|��ԙ���7/������p��3���V��[�pϤ�oMz�si�����ʊE%Il�*�E��2��~��𗷃\=���-V`�����b�LyvPD�Mkoa0d��P���/*.1�����B�=��b>�.�GF6��k�OY�T� 8̇W�B4��>�'�;�ӏݸ�[3�����E���~ܞ��_l=��f7��|��R���U�O�J��k�|��wT���qc34�d�������G;�D]��,�&��7]ۇ�젮��i���y���bb�o���<e)���ߍ���M�S�AO��*���@��zm� ���Z�6ض0;���-�{^t�#��9��I.�ۆM-�j��(�{�J���b�wl���n�0�@�m��P��gi_6.��˛o��y\Y����}}P��� �[�Y�2�Ft�稅{lIeH�$���\q&,G�)$ ��"����j,�V[J91�#2E#���2䂤���1a�L��HA�2b�a��	B��F3�RY��HB�m̵Y�9I����$��m��d�\%��-q�2,Q)b�[H0��e+I2Kjr�dA��T����VfD�ۖ�T���U��HH�B)��$�(��$1�E�$�	
�Aƶ�"�� ��2$rF#$qT�dc �q�Ƞ�fA����2,�	FGH�rI��"ɒ�����a%���"ce �W20$b�H�BU�dH"���"�����B$�W�BA�bErH��0F��#B+E���XBB,Q��1$E��	���#��#E��=���$�s�ky#3 ���]�Fv�6�p9pD�nɚ��]=tIw�K:��  #Kܶ�����}tBsw�.�H�n� �ܶ��CLP������� ;w_̪�k�� ���/�$���"�Ov����&����0�/��g^�n������xg�ƣ��"�s�k�]�]�mه���r'p�p������ Wӽ�ii���uR����@����[W��W�R�mL�i��\A���`�^�j�Ez�ّΙ�#���� �����$z{�n� ,Ο8���� ����6���e����"iXb�ۋ���M훋��umtIK��z�D|b�u�����l݁�V�p!�r�9��}����Z��ni`D/fӿ��Nnͤ�ü�k�����0n{��Қ˲�X�I�D鈹�}����;Բ���`~ڰ��Tܬ�4��n�	!��P�y-����X9������e�\��U�G��M�d6��(c��&k�n�=�jzf� #V�* �wm� �ݛ��>2}�jU[��=*�*�n\�RCc{��Y_:�޼�1��n�.�t����ο�~���lc�J#~�����;vn, �=�%DlX���=|���{�x��PO��v�_�G_������6�[���]�	8M�[{�?z��xyI� I3}�f�>6}�h��R�[���U9���}"�S2�d�KN��Y �s��I+�6[��~����5`@-=�j ����[�N\2&��b��/iFlmk^��o�� ����P�Z��kw:����������/-�V?���0s4��r�D Y�/���RJHK:]��� A��s@� �y����#0�7�j��S�љ���Q��q��/&�u#t�8��ͬ�L6�\�*�=�����W��JԱ��T2P�O��j+50�j\��@d��.�xN"�hu����&
6�y�b�7l�&�����=vyy�'gחV�]8tc̝m�؍�=�8���+�]N�ez��K�Md껟Bě�����U�pTVSlu�:^�*�v�R���Y8�y�h���c��i�XCs�Cnr���扷9Bo1�c���PC�"v��ԗ!�����Hq%�'Ksл�Fa�'ؼ���c����X$��6����U���Ƀ�nHx�ź�4���I��&k�iX%ǵ�  w�݅�~z�n�h�D�m��Ϲ�@�����"ZP���	W]w@mNA�wx]������}a >�P��]�J�f譾��|�`��tԤ�bq-�m�q˧)P��wI �O�W��z�$�z}�k���]�o�nO ڙ��%�Kz����{ڽ��0��)P G�p	���=�QI.&�����%����"mXj���$���wdV�c��~��ΩT yo��V7���|m�<��Vf�{�ͶƓjR�-1<�d�wFwX57����E����Ң�˭�m�~����m�hrg|9�s@��y^m� ����$��@�N9���L�ǧq�J�W�wA�u��@�p�ZQ$���5��,0����,�߄�!q�S��K:pn��go��g;ط[�h1�G,X���Mi>�ˠ��c��>�`Sbٳ�����L��r���x�⻥e딺 �<{�n�Yݮ���M��췙>ȭ�U�z�+��$60S�H�w���w@ ��]ń��=���}]�+�	��n�Igv�J������$��[p۲ΗNT��B����p�}qt��vn�� �'����{��1ע��J}�q蚒�nBa��v���M��x�s_ǳz��Ԋ�軈��`@�ݛ� �Oc�	�󬓞{O���g�˙%���9���]�;5��`��Iz�wF�fj9����}�ƴ-Cr�H�\U�N��{f�> ��T��iE�>�FosM{�^��@ӝ�i\A�]��nSC��s��$��z����NymU�$��J�x�sP	(޿'�'ܽ���{#�l��)Ĵ�I��f���W��� &����Ⱥo�s.;/Ywk��#�Y{��S�����gn.9M����r��k�fG�u��Ǧ~[���/�z�72kc%�3{��ޛ�" ��ٴ��Oc��73�[s���n���=vՑU72 ���, ���I%E��yT1��߹y��]^�I_��M&I	Ķ�e�5NRJ�<v]�ێ��!bۈ[����c��@^��ܕQ��U-��o��Y	T��*66��i�=�sm�]�E��'\��ld�ո<n_]����&x1L53/=��c���H�/��9�A*�'_eZ�:��i\@d�9�����	���q$M+����R;){\��n���7��" �z��Jo�n	$7�r��wS������?[m49.�=�j  =�9\�����D���w� l�9�@^��܇��*־�q-(d��@Mw6�.��{Вy�@��j ����,�>3{]��'��z=����U<�^p_��r�1���Ad;
���G0����i`�θ;s��nΣB�e�28z"\�ԡ��J5R&Ey�n�����܀��t���\-��׌8�r� {g,I+�7���lt,���g߿ݸ��U��1�5�	bY�WF��x�J윰�m��M�I_������S����?A�t� 7�9\�����"��'�JKg����@" 3�r���Ҫf�c�˵a���X�m��ߣ����7�Nz � ���Y ݮ����)d��^�sP.~��	���q$M����ۋ��[ݮ�����R]E�5���� }��q#���w�ya�0'.[MK��s���9������h�t��H ݺ�+���5�Ϯw�X�@��lW��,���ZPɛ��z��X} ��4{�sT�Oe^S=p�>�������O��S��+ine����ͿSN=�B��Sgݽ�W�>�NoB��W�lM5�d�Qr�9�y��+[�'E-v�n]��18%@uzԓ�NL����9�u�@��|��;u�É�YU��=�l*��ؖ븛��n��y69��8�����z�ֳ���PrNp۱���2.�0�k�δ$n�)�Dq�\��q�q�.y�׉8���x�{F*Ћ��[l佧��ݵvS�{t���R��]ڻ n��Ȇ���5mb{s�s�)r����s�ʵ�k!&ո�;���띷.����i�ɷl������.W�u�ٶ�Z0L;���>l���j]-�L���n�|��t\@���� ���R�.sz+�r�<e9���븑 D��Ҹ�Y�*ۆݗl�s_R��vlQ#67����	fn��H���r����r�S՘��5��J����.��k�w`���n�">����Ys��  n��� {��vR-�fZ�2�H�Ic�o쉯���[0���������A}��;N���Y�� �y��ń]Ȅ��i��W��n� �ݸ�,#�J��6uGu�{y�)��V^�7P	"��w��,�:{ջ2�"�"i�.�Srڗۣon��p��ϕ��rz�#�*.�?~�c�st���;�5����[�n� ��Wo��������v���n���#"�e��S��n�:��Kb"�b�>@���ov���zv��F��aNP��ܻѿn��O5��қ��{���wǕ��7m6laNUՕ�Y��� ��U @^�;��zJ�����/7����������T%��/��M� {�ҰJ�j'{;S����/���@�����ҿ�ґV)l	j	�j�z�ڇ(/lw ����  ��W� |gv��.�j��B�Ux�� �ԋh�o�.��Ik�{ ���wd�����w�� �1݂ 3�]��>�J_8��i'�h�\�dɨ�:r�;#�p%ܑ����miFjF�ț�<��8ۖԡ����@ ��q��wk���ԭf$j��=�OL��u��Ҹɼ���Ē�HU@=٨�+�
�e����ǂ��z	�c�p ,��V	v^���ő/3��#ّ�q2��)��7w��qa ��w C20��]_t��ٺ�����O ���.�?+>��Ѭ���1��N��N�zܞm��CS��.1��J�Թ�i/ {=���f������y8�Knt_�Λ�F���*�~\�� ���wa�$�w]\@g���VT�ԗ�� �o;J�ґv)l	���j�;��ŀ���vvN�/%��w�ks��_U��>3w]�Y�n��^�֣{�)�M�U����i�^��ݬiUp�35�ۚ$p�a���G53-�2�ʉ���z�"� [��� �>7�MT[���˷++>7;�$����jWhn[R�%\�n�	ǳ}yyy��z��E�$ۮ�  7��I,'�kb��^�<Ȁ;�l��-6���%��s��#�]�n����^{�D�?[��堑v���sivdz*&[�%?���"]�a^˪�
�� [��� ���I*/}��r�*�m�;�j�)ެ�(�4�ZԪv���Ak��N��2�!)��O�XV5&��]�SԊ���<Zy+f��Nz.��؃|zvX���ۆ�鴫� 3����غ���̶�� |M���$����� ��;Iy���陹�Isb�t�f�)I��Dٶ{IˑӶ�sn���Z#��F]�P�Gݰ��6��&^.m[�p /{[J����U��tnnz��6�z.�w��+ ;�� �i�s�ˇ�����J����<{��g�WW<� ��� /���S1���ݞ���y jYar	���]�9�� g��XG��5�M^����E�Ĭ����G���i_�ζY��KI�K���jjZ)���+d }�� ��U��f���q��ksѰ_Fc�S�U�w7Ay�"�e��S�6��	��v	-��qd�j�n��4�U|ڨ�H����J�3������{.i$�y`s5����F�����5�P�N��G���t߽�~�s�ĝ��M޵�}�{��I���ogw��;f�c}��:<H����!�z٤�nU�"���:�ǵ�3G��x�5�cǅG��.�{�zN?x���c��� vE���`�&E{pޡ��.c�[���z6U�Gz�`�`��}R;J�qt��j~-+�!�ʭ�x�ٸ��r�� ͹�%�@�EҤ��;+*�!�]I���F�n�F��4�n�v��5���=N�o�F�^R���4wmfmޓ�%�-C�}beu�f.S�q(�u~��h���������ƞ�Ira('*T��,ǯ��8����,7T��t���rKD=38.9����qFC:�ز/�9�D�;�3���"�;5?*��1�W3%c�u�Ș3N]��Uc�W'w���u�y��w���B;u炙��x�eM�$�f�B��]30���hV�mȅ2�Ȩ*�ʽ�D�L�D�,������ǀ]���ώ���Cqdi|���:n^a���t�'�68�sO�O�5��	r�|�냦�z�b>�k�o�����+�Nn���!��y'�\���F��;w'�Y����M�.'�m3}�_��ˇ����ۨq(S7�>[8&̶��ݼu�Yt�ՌԽ�g�cto*4/MԽ���=�yk1��8���_i�e@7(���^��1nq�]!<����\�ɞ�'Q��f%�����=]M~޽�٩%�Ud�H*�#"�ɒb���Œ,�8B1"���ҋd�B+ �WD�UH�r$�`�*AI1"L�(��)2&rGE�"�	3VL��2d�F1$�$UH1PWI2[��fB1dI��Db9 ���$"����$d$`�H8�H�0�1$ (�#1�����9���$%�[!XđH�B6ҡ�$��GDRqI��1!$9	&ATH�V��Ȓ(�bE�F3d!!"`�����$qdd�W#�@��,Y"�*HGc��- �Dc1QE��"I!1�(ŐqE�$��B
�c9H"�0b�HFQ"�pc&* ���bL"T�Kj�EaY�"HA�Œ)!2Q�H�c	H�W1D�iG�FE1d���L������bA�TQs&A�dq�*KL�#�H�d����G$�q��$�	d��2B#dD\\�Ab��"bK(%�Q�I��BE�"��� �.*2$��V�߼�n�,�E� ��mkz9E�e�v��觶�l�;0$=���l�B��k��U�����<d3��.�c����7����ͻk��in^��yLm�oZ�9U#Cn'n8�fn�=��,=v�ˡ��:w+�WV���F�ɮR��v붙�1�����.�c ���'\-�k�.wk�ա��]�v�/��s�r@�c��N:��B ���N���N�{u�X��=#�99���/dm�g�����<pv�Q�-��;X�{sv �\r[S���0py���/'<n0qڹ�s�.��\U�3�n=)v�nb7=gb��cn-΃������N�3=�C��ytc���a潣1	ێM����n�{=YNǶ�����@AȌ�׶u�#��gmy{Xe�ɜ��.�7���\ۏb^&km�q�v�氷j��۬r��c3�c+�-�vLl�"����z�
R��ܼ�^ͱ�Z��{�`�<��屻2�Jntk\cq��x�ݺ��K��\�I�!������9!z�x,og���Nǳ�v�gl�s��F7e۬��+�Y7'f���q�K�:��̹���O������`�G���;`z��:�ب�omt���$�ۈv]s����'��!m��Uր��6v�Y;;Iɱ�n5�<F�m;3���+i�۹���U��g&Ӽ��u˹ʹvKv����2���v�Y^��j��ۃsb�7V����ݻ�+<�x�g�ݵ����9�n^�y�3R���j�k��N��N�x�cmط�cn��Xw]DN�GC�i��p�K]��k��=���㋂��l�q��(!'o[ӫ{u��s�h�-���ktm�m�1�h�ѭ���M��uƵ�kv	t��2ޝ����۬��m�^�i�$�dۣ�nً[��7�sc�F���zo3�kӽ��K]�vDW��mVڧ��cE�{nV\���%��A����t����[]��1��X�ݸ��1�`e3�F�����q ¼��k^F�����W>�u�Y����;��)�#�;���Wm���OY{og@٭(hLd��1۫���F��!��Iş3�zc7j(S����=t�a�Nk8�������	�9��1��Χ�z=�U>�TY�#��;=��+դu�Ղ���*f�5%qft���K�x�	��n���+��+����n=[�s�1��3��ÉƠK�c��0i�!���nt�0���g����`��9۸���Z�-�ڶ�\S�;��e�ʉq-�m��:n���1�X|	ok��6z�{�*L��n��s��}0����˵a�V���WQ�So'��V'�=��� nnU���3{]� ���X����
�_{�[izz�˒e�L�r�mXv޻� �k��� n����QU��@ �w$� �7��W�[h��6K`�%�<��t�T鑝^u�0;�qa� A��w`@%�sz��-�^XԵ1 Dw���{,��c%��%�>�$D�kt?m������v[���{7]�$�����~1��Ͽ�>�[vySI��8�筱s�j0�.ㄬn9��+wc�&��������\ӂS�6��Ezk�R v뤕��SI[+�7}�ܿfO�f��WA��w}+�,�H�ۆݖ�� ��t�΃8��=�(�OY��=�t*��R,��b�&c���.��˞79��W/�Kt��k[c���<�o��VN����|9)�5�l�,��ğ�8s�]� 	{��|�=�r���3
̸a{0�\̸r��&]��3��� ��� �{��^z{/&}^�� 3;]��^�7P�b��2ϥ��Dҿ�8�'��w{8�u�� � �e5@_��n�r�s��R�����6&:չ���[ ]�<��  =�ež�?7W�Ǣ���MX {�I��w�:ʚ�̙�G�f�Q��ӻ���prر=��oȹ����'S;&��FL���ϛ���&g5�7�� ���U��1ӌx�8�{jz}�M�  g���#}�cp�?�i���+��g�,���Fz�Y����H�SU�Ǻ�!�"}��)��WMz/#���3�[pۡ-��P��M�eZ�	�xn��v�%��]q=���y�Nl��%Ýa�a�O�ۂ���LL��:����h��ng��*����4�ZUV��a��\A$絺�=�*��]�ˇ2ԥ2�-9��_U,����f[iP ^Ϻ�� ��ٻ��td7�`@U�u�V9	k�m9R���4�]�����!�����^��?��~\ D��?'� wk�OO*��]zc����Ci�n͵���c�9ݵ�k����ۯ&�gT�]wA�pnZ&���\�b[�l�a�u��>a�i A����J��^+�?�n���=�p��z���&�Ua5���6�{ӕ䀵��� @�u͂G�ok� +���WH��h�O6���3"܍�9b��n�&�ꛀIon��ď��������> �˶" �;�݄w����f%Ķ�B[-�Oj)��nԥov�J�,�U'�f#!����{P����n*y{{�拳znK�qKÏj���!1�1W83q���Y�y�k��L�	&�`9`��"�-T�R2�Oʆ���R=�2��q)L�W�V�"� ^�7PuPr,L����+���w �Y�n�ǺR����:���Ù�vs�����ȝX���}���G��,�ڞ&��ێo{�چ)k��r�@{��l�ov��ď��=��DlV��y{_���뻈b>��i\dLo����Cs �Ҝ�������pc�=^���@��v�{�IPzp���������=�Z��%�[��*�:��K �[J���rA�4��@ٺ��� �7Qލȧ#sX�6��	���آ�D5{%� *�[��#�>���T|{���N�$�7���W�nT���[p۲Ý6�Yǲ��7���L�e�� �{�G���� A|{���e��lnG�^+W'��礻��Si�ۺ�[��?~~_8+:{1���)�6��i��y�4ܗ�5���=���nx�Ǩ�o޸ڛ=c8�S�~!LH�+�ݰ�p��s�!ss��qz��ƋU�v`�}��sg/���"g&q���^����fm�nû�%��Վ�ݵC���N��q�nH�g{���u����d�nu�y��@�w>7��v����]��5��..G�%�n��ͦ���6Qh޿�7��"v��7�V8�9�:�ƚ�֢h��-�$ ��k9G=vN0�
�Ž��]�=sN����jS]�)s���5��}v<��}~�t�JS/���X�������T�"=-]�]�,�{���	%���"}hb��m6����3��Ų67���Q���XD�WǺ�����a��#i��j}ާ�g��Zr�saW �J�aS��/gѝ�fc�-���J���w�3j���Jn\�h�v��yͥL�k�=f�J}ͥ@�z}�)_�A���j66�݃@T �/#�-�l��6���emM� �;]������q�}�xH�MT ��r��,��V}��T;�Uj��H��bO�{_2|(��\ݯn9�ݹ^����n�"�B�h䵪������t���[p۳�y�u @i츶 ��]$k���<�ޖ�{z���" ;Omʸ��K��K�-ĥ2�\�[��%{O�ۧ�}PG$���u�������E�8ƕ��ǭ��ŋ�s�XA�F��!�s���<�f�7���tZ��|>���bf��w�OĜ%�?-J���w ]��q��ꄷm�|>��17ᶂ*o��7�l �k��6N���.{\V<ֶ ���b 3�]�q�1��r���0���7���E���3�Mw�Ion��H�3�ޛ��݊�:����\��YA*�k�݀}��@M�P����f���� �7�7���v�� |d���s絰���)w��w"��wv{z%�����[���Td�zD���Р'�7bz%�d�s�l��d@��7b@>�P��w�n�%���7�ۿ����5p��=�ʙ�8�.v_�˧4��������4���`;�7q @O��|�V򠪛�fK�sr_J�>cp帔�]��g���H�4�B���"{��@s��Αp��9ag�����LiG'3)b�S�(s��v�{ۓ��/��|��!^\ݵNm��L�>ӝE���� ��ݛJ� ��9��m����)i�.o��/s_{�TL=�Y�i8���&��� 0�9U ��9�2�P�*�L�훰>Ș�V9hpK�C��s��> =�TT�_���V��יul��$A��9I$��yt�4S�N�
&���2�[����o[X8^�����F.9ӣS�
�2]~>�����V	�@���$���)%_�̠��s�>~���O��� � ����#��7,�r��ӛH�������/��׳� "�k����%A�jf�;��4�����nT̉Ĺp۱i-Ϡ 8ʊ�.�0ě���M�\@�c�D�|u
�eY:���LL�KNu=O�t�@'k��D���FC�ʙ�C��Е��f���Hpyá��OoNZ�����/�76������j��\O�{wR�����'�&X�������<e�J�N�Z��q.G*.l7K�� '0�o����<xM��AP�MhY �zu	Px�ɤ��:b�7^�c����x�����|r�kpe�O=���Y^uױ���&Ԏ2&�z.=��-	sa��9���a�R���wq�[�l��U�$��r�� �6�B=Փm�� �	����w%b�O�����V�*�H�2v��wc��]��o����+�-D�BM�7a6u}  ���X FW�I�9�����It�ڨ������c�ܩ��r�e�t�r�K�"�c�>
�Y@@{ݎ��> ��9�ϫj��a�J`��:��"�*��7[�beڸڷv$@x�9��nȜ�eg�DONQ@ n�;����s��*>��'�w�w}��soj�T�j����b�0C�F7�}�Ugr=�b��1��[�f[L�c:�nG��~����	��N�����pc��j&�0A�}5	 rq�V�q���炸6f��Ս����ɮ�g+�8��v9��:�{gF�7i�KX��Uސ�=n�[�	���ݎ'4<J{>����[����\z-��b�ܮ������v�M.�j���A.��z�t�i�=�e��7e{\�דnm=�rC�'�>��k��"eܛ��;^��8��z�vS����k��#���ۮ�5�]�C���`ݴpWV^�L��y�Ck�M�������~�8o��q+g������ �q݉ ��ڨ ��Z�Ҷ0��*�$@+��W lLm��8%�!��<��J�5.E����l l�d�V���IGf��7�=�^є��8ЈMU�5�7b@.��@S�Wu�{Q������}�7`�w���.;0�%�NT��sw6u�����^3�QT p���H� ���� ��pd^F#���=ݠn�ٽ�*���R�� �f��+|�!9�8��$�Ԉ �y�����O~iv:��IЭtL�����W@��sn���n�xym$�${q�S*f	��cb�:�_e�׈ ���r.�ɛ��B��s�����P8n&bq*�g]�\���`;W�H��q/\��Qg#dFUONֺ�f�G	;Z.�\��Vs&Е��پm=#��<j�s�Oh	���)����	��Dy� s�/j�j��{9Υm*�8%�!�.��ss�>'��.J��o9�Dgg:��/��K�̶����\s�޽�{6t�M
X�7sR����d�zoo��_Q>2�&���&��F�y	g�� ����c4�V�'�Z�@�3�R�$��푺aF�Nq_^>���3K�͖��e#-���rc��� ds۲u�fQ+�ڹ�}��sɯg���}�N�"��Ъ���vjG�����e r)��;�2F�t�A��B��]Q��5^�5Gu)D�ݣ����f�uP�A/���C��rλr�m�2a4���T$TP5�-�R�p�l�}�2�E�ir�YV#,��PÓ�ْ.-N��2{���-`̓�'_�1������}���t�ŞQ|�:��<��;�J���nI�L^߼�=��Vxd�kCvn�wK���y�7�Y�2{S�J�S:5��R��4׼�
}6�=�wy�s�7籞�ܽ�}�v�{��hN�U�퍢R˪�ocS!�70��ٳ	LN�����\��l
��4��7ݕ�o�eB1^Xgn/{|�8����z����F	 ؈=ǻvd�|�z�{9�\���*诃3�W��Y)W�I�����Z�x�}ou�r]��W�܂w���8`���Z��BGrW(���g�V��{b�;����oQd>��y_a��f���5���x�{�YN���^l�q��=�`���}Vғ�:�DVj*E3��h�m��V F�r�!-�:"h[)��]	]9�gu�^t=z�{���5�ڷ~�z�kR�ڪ�~�s!�>����ÐdB@��{��m�зj���+�xԿjLj��j6ݻ�OK�<�Lq�F�ʦϒ������Q���	��=�\e��1Ou1��4�b�-��f�ub//"��8�[��2µ!DZl���h�ۃNsȧ�f��-�9�<��y����9��:�s�g���%�7�i������fS��=��뇋C���=���R��շ�Ws��$דR�q9�x)T��Teέl�qD3'a�h�q�E�ɹ5]��{%�5��~�x<�5e���z{/�|pAF��j
��<��wQ��ތ�6��{���瞛�rI�8�[R
���!$\#��Q��U"�$�Y#	B1�Ȃ��DFI���U`��AR ���VH��"@Ql��XF*2̨#d�EQ�qQ�$`A��H���1�*��#�p!�H��b��H�U"�Aq"AcmJ���%�kE��AE�QZ�TTE��d�"9$�q\b��2̘�\*��)�DAc�Q$d�bE�0�AW"��1d	��*����XI�q!	�)��� GE ɑ�&8���9d�H�E\"���Y ���"1�(� .
�$�eR@��1d�R"62IR8�HF �G�X��$�dHBDq�#�$�rL�3! �dPc!&��LR2+pI$b8$�őfdA�I"�,I"��Ă��f
đŉ"��2F1X�a�"�AD\cQc�ATEI3�I	2
@r
� ɑ��U�D,�d&0��Q"�H1d�1�Y �#�Y�!0��ŒEFH��c�$���D�/�P�������f���v���2����FD"F���>$�ݲ��&�u#�n�h��J�3��T{h�n`bChD'w]�Q	B��m#59c'�3ąU�xv9쁎��+-.��*ɮ�3"~q)Ԥ	�b���dΌ��m��㳚z���燄x�[�����~��hDĊ�Re���{(�1�P^*OLn��>��H	�(�|6����*\�mݩ�N�]��Í�-!�IAӝ��>�s��=O:�.r��%h�9Tj��W�MQCaҔI>/3� I'*9q�:z��I;�W�������D×
�&�s���y*��Q}��$�Ƽ�6�QbLmn;�Έ��{�R^+7ľ~ʼ����)�}��܊�.�����������~�S8W��4;���ʌ���������ֻW|�E�5!G�P僅.a*��D�s{W�I8*;��tO�璉� �Υ�'��j@�A����OZ�+4�󭵎:��{:;l/G,tݷ�<����5,8��Sy��sHЈS��Wt�I��A�j^.rf:u���َ�YÛT��m��(���1"�ԣ� f�3%^��m#��� ��@(�:{)�7p���5��0�G.%����*@I��H�ҳ#��Nh��ɑ�U7H�@/si	7ݨ$��uF���z���U(\���H1-R� �_n� }��HtۭqRr��]H��EP��ߎ�bD�3{ix�	
4=��1�E�jĞǴ��}���k��u���|i���x܋(�g����F����_"i!*�����̧��Ў]�3�����~�W����_��~���|�q�^�c�u%5��\�����xƧ4�̻�:;u���!{��c��6=�벦pDpV�7��m��ܦ���7���l�H����\f8Ch�̚[M\�9=��N��)�G9w���9�ò���գU��n`:�<��ޒ�k�q�m�;m7mb�q�=>� 9�`�6�h�c��F�cV���\�q>���ɶ�-��&7T�W\۝�u�r�����s��my7���,�9���*��qh���.NZ�)I9�i	��	FZ��n����u
_^�TW��q�&Hp�:�A�%71H�N\�R'ē盩x�H9ݴ�mM�ݼ�1b�:��;Ix54j&bEI�^0�H�C紁 �p�t�d��1x>$gv�I'm����DÙ�������:��(R��K��D��y�"�������H���	��F���z���j��w3�G���ՆB��H�M���"�u�Of뿣��Ӗ��9�]Y5&�)!iKJ�v�KXw`�;n���,��O���Ru�o�??v�ͻH�$���me/Fk�@�"�9D#39F͹ԹUi��m/�Z%UT$ML�����nR�<n�ףq�w5ʧ�	��2��cp)��v��i~��7�W�Ps̈��=rG�G��B�Vn��)��dД���v- ==}0�>���s���~D�H-�� ��������W=�L���tk�&H�	�Kt�>'���y��$ou�5�*"
�@	��H���#|�f��LD��Rs��q���h�A�ԉ�ޠ� �o�r��Uu�Ɖ�ڥKč�a��D�L�ķw��:��Yَ�z�q��Q�BWt� �o�� ��j@�b�W��k|�>I�g�iJ�E:֯��Vn����s�bٵ���漜o/�ǃ��~~o��uz��u*@�{/�A$�}�f���Ӝ*�33�H�K��@­d��U�R(I2��V ��fP���@o���H��@^oeF�Y�G�t�~��.���)�1jax�gR �7�ŒA��r	��J����ڲ�ٹ��:W��ܕ���6v
J�r;����.t��!�ӓm��Uc{C�Bsr�=�eJ�\A:�i|M��w�Vҍ��3*j@�� ��[oU]���"|^]ב9���[�W�p_Y��C�'��n�"f�ԑ"�J�}�,�B紼Wf&҂mV��>9�I#7[�d¬�q�y�B�����a*[�����|Z�Չ��6۳�]k���hG�����֧���}����a2ɉn�B�:u
,�ݻI%
�������\v�ˆrw)I���"�M�m97�ڥ���U>���f��G�Q���'���7u��I ���6�ܥ^��}��!"�rP�7�N��{�n�!gm/AD�o<<�)�I/�w`	omA-F�LE&�;Yն&\fޭ��t����ZD.NŐH!gm"A ۾�9���\f�;�
�ەZd����tdΣ[c�qNz젂�I���F�.�TQ�7�v��62 �ϋ���=���GU�l�}F˛��>[�d\rU��qq^ts�T��	�*y�� �\�9�|��vl�L^�m`%��݃�ix�H6����q�f!_���ۮ�"����yݞ�k-�I�-�p=Z۶��c��H��b�@�=��trR��A"p����,B紉"����Du�'��m׵Y���
[�M�˻��N�����	#J��t��<�$�nm"I6������^�˸���#עl�Q��^�5E c��D��:�"r^���y�&�ŷ݁�ssi9}ԼO�,d��U�&�w��{|�^�B��G�yב��AA7�z���sױ�z�3Q�o�SYn���-�CiÐp�\����$Ǐ�[1���TD�q�ď��@F_m/I���dr�9���SL�����3��,�����F����M����vٱ�d�ԑ4��Ux���\��T�VlS��ܖ��i[x�ݘNۉD�����,�#5��e��(nd��@CՏg�����E7Z��	�r	��ȡ:�GcmI�^6��c��ض�a�*�{v�ՓFy<c����sq�E}n-�k�A��틋�7�>|;w=������1�q-b�b��-$�̞��Y����^�Z6� t[W�����m�xN����t�����һt��m�����q���N�v�+n�bS��5J[g�;m�k���g��rzuŭ��U@K�������1SP"K�k�|H7mא'׹�vF�pL�P=V�O���@`�&j�2'�F��|�U=�ݳ�ݥ	x���� ���/Ɖ7��]��ҙb��)��|�	%3ݷp���҉�/"p��eH.�ix�	���o���Ff(Uz����WC�)�Ӵ�&ﶗ�$����ĂK]��*�e �h$���	��hК"f��Dݝ���]�'3#Y���(���@��'Ď�}v	5�H�Y�r���	͛]0{�������caqk�;c��W����cg�v�9`�����Z�������H-��>$�m m��FR��"����P���m�%���$��9dvas�H3�m)�����"0�.sj��4� �ʫ����8��٩��҉@�_׿s���R�r��~4��A����7wQCC�J�z���.��ŀIk�� ��bVD�I��X-LЈ�I�B��Yܞ��$��Y�b��4�i'�����[|#f��5F�5W`̮��\-�ݪYԻă����'ă��/I�}Z�-�]��Ъ�`���^]��^	�LP��Ъ(�t�$����u��'ѽyb���K��6�R;W��~"��&���H4�SK'鞧�s���{M�A �6N��-�����������!4D�+���ۿY� �OiN����Ɋ��V�i[���˿H-=�Y'QU5*b��50�޺^$��$,x�(����	�'V�/F���31�-Vg�]�{tk�TJd"	�Ev���H��Z�m>
Ҳk`�E���J�ˆ�et�-�6���y��v�p���HJ�T}BR
�_��2g�.T `����}�4�1_��'���ݤI>;}ԍ�:�"�W���P�k�6�A5�'Da ��T�H$�;�Ax�}w���<Brz�6G�ԉ�rҙM��ڙ�qP�,��_R��e���t� 	�w����w����6�m^	�f���7)A�s	�e���8^Α���W�bح�{<�C�N�0���~w��n��B����]/>.���A7z�����v��<��J�7��@$��D�[��P�2f��;y֬�K����q�	�V|O�^�����,��a�h�f��q�.(�-�j\���g[��9m�A5��<��l�R���v�ξ_]��_�=�5�*%�)��ν�c��2H�AS�K�$	�w�ذO�]�g�]��;5u�$�p��;KrM�$x���dc����\�|�߂�գ�#�S���u~�*;.wVK�	8�K1�t�wS��Ys�5�(f���1?�!�!v_w֒�{�$��#������y�ՀH!�m#9�s����_�g�_cQ�-`�Rk�.�������7m�k/7=p��:eO�k���}���l����}�]H�;s��	w�H��-Uҹ]E���D�t�[��J�&2��7�:�D�F9��l^�FC��������C��@�z��y��71Ұ2�d�P�15&Mz���v��2�iEF�)�	��uG���~��}�� ���r�MK��rT-Λ�YW�gvĦ����	#o������'�zz���.W�u�w�Q�u<��ؐ��'���/��B;�
L��D��Ix�AՙCb�<�~���`fg����3?�`fa����3̀fa����f�f��`fa����f����031�@30�����fa���큙�f|f� ��3<030�������^�* ��
�+���
�AQwAQsAQ�PVI��g��2 v` ���������  }�PP �   �J�   �4 @           
 �
h�  �R��TR�
�R�m�4"�ET�Ե��]m1	Qm�F�ARk
��W``[ٮڨ���AB
����J��U�                                    	J       ��Ϫj�Z����w�N�.T=����)L�zԡr{�ݵ�^A�ս��4)��� 7�I2˼�f���*	)%]�   {B���_L��N��� /y�*嗞qԷ�����x��rS��ɭL� R�LۯsT�y��y�o"���{�-+���IRQ�(�e�   |         o�iA�w}q%y��=���ʕ=3�)֩{�� ����z���^7�#L�#T��cR�s� �$������-��b�z����c�   9�o��Ҭ��1��)�� ��J�6��T�n���Q��ڲ��퍶��� xt�eɮZ��י��y w׹���	�u��;��V�   �       :�ON �@�� }��  F� �]��t=y�yp  ه�� δ4��>   :�h/`���� �@b� wcW!��.n  $9]`r��px�%�7��Y]�Q� �        J%B�T{2%*�b��d�W-T�G{�O��PO\ 2UIUe�r�����J�n���҅/���(��}w��%T��g�U)Ur�%^�kR���>�   zR�����ܫ�Ԕ*�w� x���,`��:)B��9�zX���  ;d�q � p�����x � @        �#݀�B��{@v� @]����]�u�&�C  ��$���[�eْT��m�>�@+�Ю�q�a�p 7K���w>�O�{&ԯ3^��g6U*��x �Ӽ�v�&�����C�Ne��T��O&���M=M h��b��@  S��=5R�4��ت�jRP# #T��i2�R ` M$�)H�������̯��{�0)�l�' ����?�3y��@�$��<޿�H@�nB		�$ I?�H@��	!H��BC��������k_�뎞?˾�Zy�������u��;�nS��8Qc[���V��t�͜�)��F�)�pi��d���;%s7%�؀w�A0ƾJ��qCr��PN�Nw&�ݝ�х6�x�s�� ?&,��[���|�vc�V�w7FYq6H��<j�:T�A@�e���L��,�xg.,1E�rϷ�4	1wd-ⶾ��,,�ƻ��j=ɴ�oB6F���W02U{�{;���Q���2� ��w{q��׻x�����<R�G�Ĉ��FQ{�/��$�$K�3���M�X����w���/�jk��g������$�$�k[���I���9�T��[�Gj�E�5nn���0 ����q!�َ�� =�!� ]_�:���X��nږ�l�Yw�CX��G���H�Z��E)no�v�z�h<w�aFW���x׻-�X��Q�75m�E`��ϰs�<Q���ORZ��EVk��{78'uliÞ�{I�Ց�B��gOQV�7�����}�=U1b'��4�7r�������s�H�vY3����4식h�Nr!����My��΢G�fǚB�xtv�>F�X�K[ݪn�� ݼ/'��θ�uֵ7P'�-�Ϧ��/NӎL7(�wBj��}5���26�Pޫ����`�|��6&x��'�3V�X�x�YnM\�s�0��7�v擧�ѱ%z�)����,7�hL���L݆9�ûD"����gG����+;�'H��Ê��І�0��VM3���0�{6��XBݢ��wovo>�WV�z �7 )��Ҹ�pꬣ6���D�'��j�3�Qc*�!����E=߹�P��*��Ɂ��i�B	:`˸��֨�w'8�a)0�*gv����S,r̀0�7���!v�.��B[4��5
��4Yߖ���2 �p�^aưo�H�w�ݖ�xo0�bt|�l���r����7��Su�V�[F�����L����h94��l�C�}���<��7�q�8W9��1H)�nI�1�j/�y½�9�kYZ��E٬U�u�o����y�rX�.�㫵U0��]Zt^<�:����M=3�G��SwH�x;K[��OǶ|�I�q��Z�A�j�m2�XDp�$0.�EEf�8[T�&�>s*�|����Ѯ��;�O�w�1�c1�ԯL/�.o���ܜ�\�U����8��J�h�x��vn9OKrC�k������ݴV�"�,�.;_-ȴa�䳀�|5��a<���,.2!91�bcch�.,�pp��9��O�r�Kфf�z����7�ũ+�3նp��x>�ѹ�A�#0�:���1���G�1�홮�����_j��G�6�����;��L��ݛ�2:Sv��kY��,O'�&�v�����N۷���mq@ޜ'K�n���m;�i݂��X�<.��m��V�1���&�8��=fh�8��ޗ�Z2
���OL3�fhι7J{�uW0����R��`�;� ^c�.�F�k�Ǐ_u���j�m�x
���rV�9����]� u]�ln��l��,�=ޥӜ�b����r����Hٝn��.U�����1tcF�:-�����sE9(���B�0��:�!oq���}خ��cѨ1n�5QC�ꛨH.�IU��� ��ǷLFr}��N8�b��w	�>�h�y�3Q�]�-�J]���5.�쳻�A3�fCJ��7��J?^��{2y��������EN ��5�v5�u�ǃn�(ٻϜ��K�wІ������!g�y�٭���f5eQ�^u]�fKՒ�Y���L�o�ȋF�ől�s���y1�w��U9pX��tNv;��@��REg{M���t���PBl:'Bw�%���s�Ah�%��������%Ԏ�qE��зd��Ǭ�s��(��:{�v�tr+��wp�9I:�g������o;Ŷ�|�=(�00�PHt[ �|�Jw6H��h�n9����{��^�Ȕ=��21�f���[�5xk�_�s�Ԍl�	����Qu���vN���)�n`��)vr�@�k2]�3wp,*.n椺٧�1](�ۏ�HdX�,u`wS�i��? ���f�m�0�I8�U޹"�yҏS4��s6L:������1Ou�I�t���wV��؊�9+���3����f$�����Dp�y��@�G���暈�LpD^/�����%�|�2q�#��˸"Z��qW`��u^���	�א��@���l1�ێ�+�o�c���;���2�D��h����6X�ti��J�I��!�n�\ ����+z�n��+?��c�^k��Alt9p��D�M��+i�#"�u]��v�n���y�cq7�ӂ���L�s{�X����g���h�:Zr�WoY_]������"�9Ӆp�m+x�<9��:��wy�n��Ol�jд���WQ�a���%���Чf�Io!��{UP��Yʣk֖���(��Tc6���x��!zڋɇ9D���pY��7�lˌl����^��@d�c��:��4$w��.^�8`�'X�*p�NM�ɝ�ֻ(<���oU�pXAǣhy��7g�J��P���Md�>e��t�B닖��׭�7�Y{���7��@�X��F����*�u�8�
�-�jK�ۑ��6�����W�;wu�6#�㘻���ƨ'w���Sߙ��t[���L��K�K���t�����3I���9a��I{�wS�3v�Gu���H�N�J���=�0�5E͌�9ކ���J"5M1n����Q�»bM�����4�x��g%3kqS���R��g�p���^]�)Q�U/��b���|�a���K9�:�3oo���fs���z�{���w�\2���a�hWq��g	�˵�2!L+�z������� �"��D�L�F�%��3Qu"�Љ2X3����;4w����}���#�ќ�������f�9B����ց�@p��5���+q��Bn.�Wu�o)); (��gjiQ��բT��,�㝛J�ߖ�{�@�~W��6;M��%��&b=F]�SS���E�8�w��t��؃*�,QRR^ѯ�%3юk�p�2��{H���;��x{v�3R�!Z����b�3�q�r)ň�{����3�$�8xc�='�ͣ=�P���ѭ��e���@�,ݻ��YH�������0�������Qc�����AJ��O�$c�8DR��Z��3�Ӏ�˸㜒��>�4�$�sg΄MW@�l\�i�<��9Tx	;@�6;>XV��k�Qi����o3��C�z�� tq�2�����L�.k���Okt�&�[z;r5�"��`yۗ�ݗ׃R{sr�jC��њ��߮���z����|�.o�����a�5�øIǩd*�������զs��Z�_i'����wd�����Q���m��L"]x��o6'+.M�S�.��(��笎-q�9�w`l7�k[�ǁ΀�,�x3���õ���-A���_3�߸F��l	A�����x����*v@�7�˴�爹�Z/=����%;������&�ٷ5NL����+��ᇐ�¸K�hrD�
ڏ����ڞԟs,���pѳvQG}V���JȆ���;��+�D܌'���+�h|����ڹa�������R٩��}[$#���c�p�Mܸ��Xy�]�;% �}��<��h�gonv�K).|�Ö�m��C+'��FBp:wN�Q��[�"}�`��愗��V�r��L��wi.�L��D{��$])��%fؘ��;F�=�Qk��`��+tR5ܣ�0v��7�I/s��3�|9�a�)T���M;Oѭ�Z�4$�m(�κ�r 'Er��.4��1�ۘ!'�⡫f����8��jZ	̳S�\���`����t�O���S�ΚH�Ҧ���k�f=�z�͙nUþ�.F��2�y�Ӳv��mݝ�+�ơ�t�(tI�<�w;9�m2\�z#���@D298�[m	u�p�+������5�K$�\�����'N,g��f��z9�*8w� N��yj���U�}ȗ[S��;e�n9�r6�%��4�ق�t�	��7oJf�X2j����� 	�>οk�x%7������q\�uh���OTz�F�ͪ.r��q�z�N]�����:0�]Aӄ�u����dk��3� ��9.��q�+66�f��L��M��|{n=�]�t1��bg�p5���ya��\��G�ꅔ����I��;#_s����{�I�7Itc��	;�N z�6�	ˢ�u{�tn�gs����{4��K^��R�e�E�f�{�ͬ�7`FMb,z��x���� wq�z��!ՑX1�����VG�:�=�v������@��&���[s[� <��n�wr�>X����iww4T��5�S�E���1�{�Q)�#^�˜��S���v1(t�;;E|��Z�)@���β���\��$�RV���]�w�LZ�b�%7�Ϗ��B;n��ზ�֏C�q�d�vP���9���f��aҟ(E�o]���۽��[��h$v�ц������Pi� ��S;{�]���\Wp��y�}�^�U�B� A0&q������=�xnrt�@����.�zqoZ1�/h�6��5 �b���O^왩(�mޭ�^��19�W>��[rީ�Հ���h�0�g�&�i5�����F�h>W�&<����3��W" ���Kv������M�8���r����K7I�٬9�-�G�r��?9�j���7f�!�-�[�l�ϖ8��cz-��Ş�n�)�5�5:�8�=}�ݨ���;��c�u��<���=Ia�;!�};8�S�9-�����?Hx��<���ç����a}N/Uw����j1���"�>-��5nk*o+�܀�9�[�	���),y`��L���\WL}���&�焬��f鯬�,=\%�u�#8�f�����E�\��;���wnCȳ�����M��޼�T1󒇻PQ�GGn��3�-͟pdU�S������sM�yC��(�^�iv
��)�H�n븺��h����vNx'4�b�=r�J�"KSK��v��4΢qyn���},��j᲍P�����ߓ4�;gJ��h�q�s��^���sAW�����5�Շ�;�˸����p�'7����p����E>Y��2F�'D}�5i��^o^\�P\'�8�圗x�˛��@K�\��gM�2,�1s��&�@,!�<7�عkw
ǎ'&��a�]c8S�4��f����\�Ip>����6n1������ۡSʍ��'��HdY���p;4v�!�|q��o1�k����K���VmK���B����]�<�/���2'i������֙BsN;�fG�$;yǆn��*6k]���&��$4��n��uH��/=!x���<������!=�"+��XnU�,5`��v=,o ��#��`�=	���>�!M���"��xлL$�ڨi�`9sakD[��ъ�����^0�vp�gbQ�N!&ay�����ڸ�H�W^�.�Z������F�q�ۣ�\��]ͮc�H��iw@����v�4nM�u�@��i�9֡�.݄�� صbD���L����JC��䔞C�<#��u��c�u�1��7:�û�,zN�(����&�1e�Ҳ�����˜���A�|�i���j�f�K�6>�x�9���W,��@�z<tcWvD�Ue:oNB�qF�t��]ůr��]<�\0��lQ�'l���y5k'e�C�fhhj�5�\	W���,�����b!g��B'�}��	���t���;	XN��Y6�H�Y�pP�j�5�Q�{q��X��O�ت8G�h���FO\t�u7���{P=�uΪ��:�݂*�;���2 �䌉'S��|�w��E�;�EV�<b��ԧ��]���3�>L�m���V0�|oomPN]�G:��.��|1���W�ܢ�xhDe��Oq���.-u��6�I��w����wk�[B���p��hq�CG#�`��6o�Ҹ��93���Yǃ`oo4��(`�x�u������wE�n����VA�B�Ą��=�|z�ޮ���Y��������kB�p�2T�	�d��V9�HpExݓ���	�1�m�.f��5lVVhr@u])��Wf�y��{MU���p	a[���]�;Xv�78��Xgi��[U-r f���BߑʯQYp]��*O,�w�q��pS;�agi�7�;e'qM�W&�Upf �{�Υ�,��i�q�֔s[G���z��!��;��f��S��OgB�i�;���DY�0L�{��Z��%'v�z֌X�!!��x¹tQ*8I�om�t��+����i�y���$�=d��� X E��)$��!+!"�%d	X+$���X
IY	Q�"��d�, �V*XH �� $RB ���� TJ�IB$�(@�H	 (� �!!XI XBHVHBE�($�B�HIY�AHHB� +$�BJ�	����+J�I+ (HE�� ,�B
 ( �  ���P�"��I$RI"��$�H
 �d��!
�
� %` V(�RH �@ � Aa �J� a��Y J�H,$�!���(��J���d�� �!'��HB"�@�$���$�����+����u���p<R	U�Q��Z�A-%�¸�˲��L]Įu�w=��wu��f���,���<�l��!��;�}����W}�7�����&�E�=�#i���gq�E�\�׻��e�VQZ�ǅ3#�4dx��[K��@��o�\���PX��C�vΧ�כceNʵ�fψs��͈��k�׮p���_R��y�,g& ;���.vJ)N7-;��"]MfJ���Q�M׾~Y��+���4�RP����H9�v�=lO0�z��K����R��M�L5h��ԍ��J�$��/Y�����uh9�W���z�s�ܚ0néB���6��p^Rx���24������ �{B;ʓ4�����n���A�^Iu��z������y����wϳl�W)엑���U��;�7���v��*��^���=)��X�i�9����kB(a�&��Fx���\/l�~�� K�{�k�nb��^���Mc�ۓK	󡹾�GBr�l^Ɂ�6{9���}���-�f۠��W:�|��y`v}m���J�`������'.��]�������q{˽����øb���p�3���Ջ	�ś��rN�a����/�θ[~��d��෻:�����bN�9s���opz�Qb]=|����#�)˪]ڄ�	����gVoj@G���ǺNc/*���ױI=�|���TQ���=~���k׸�і-Ѧ�8%.[ᓢ,�Ad�ө����N��$fc�s�h����>A�=�����,�T�1of��A�?�O-D�4E��̄R�D�4gU=�7T���8`�z֜�;X�o�q1r1<{�瘫͓�_@<���9�����5���}�S(�G�:D�V]�A�G���1Y�W�6��ay���<]�n�9q�w 86<׾�[�u��I�X��6gby6D#y�L��p#�E�ۧW��̈́���a��g���S�A��3uR���ӕi��t��1s!��e��:����۳�� kܪ����E�w�x�nE��n"W���!�읂��nnTt�^�d���>8&.���%��Ug��X�Ɍ�=b�=� �o�w�X�ӻr�������[���j0�O]8Q\�?3���H�՜v����x��簻u���{={o���61.�0b�Ezҫ{��k��|]�ww١���o��ɚr���Ă�̺Vx�ݨ+c^�3f�V�O=�/\��eO��}|&��݇����zcDT|U�/��s՜�u�R�7W����Y���ls�K�w<�viVi�漾S���T����ީ�/OT;�D�z;����	��|�Q>���T�译#yYu#��r������p�*d�꼬�Ͻ�˛�Ni�X��\H9��i�^*��/��t��09����]�c�Q����O')L�O�����#�4�[܆pؼ�?"�Ѝ�Т'u�7:q`g�ı�:�B�'�uN"��7[�-�f��j��3j�۠�h-^�9�yOzu���7ܖh�L�3��L�o_����0{�8�|�E?&PXwI�b9���b�?0_�y8u��N��1մ!N��s���Q���om^�hX�&�Y����3Ooݞ�.<�-�AF�K�c�i��)��i�k�/�~����̵���h��{���y�K��,�a�7��L�����z7���P���\��R�r������Ȼ�Sa+��\��><a��k~���Kj|p���y���~�A��<���b���<x\Vy��	t~����d�W;i�����=�H�����Y�b�LߏR^{�F�������g�^�㞆�ze�f��0n4ߧ��5���i*h��]zǛN;�dͶ3V�w����7� ���"�����(��Y؃<^�ћ�Oy{8����y���F��V��St�9������K�b3�U�C�]�,e�m1J;q��&�黋��w��v���^-�Er
Q�aiz{�^N�Y{~4��@b^�C���׊�Ĝ��;�����{6��M���Kv�9xnp#�{��y��������˽^r�ٲ7���y�yJ��e�%w�=��t�.�bRkv�wU�O�yT@hz��)؉Y=c{�ڏ��n�B�|��$��ab��;Q�4=G�y7��(ق*s�>��	�YWW�=�8���&�onD���p�+�g����0��OK�ʥ+�W���5e���<���۷�M�{;6�]�6��cs�߼KጰX�d�	�s�P���3ޢ��^����Q]'���6Jp\}���Dy�A�C4�k,�5�GAKk��{�o}#��u��D�&N��b1��(V�+b�o���-�&>ڍM�ܛC/��ק�8��Ҝ�n��
��Դ�DB`c����ܾ����78\�	��^�|ڞ����(މ�H��4�V�n�*XxGb��X�|�>5ʮ�Rs/�z�b⡷�&�^H�Jv`iAP�nS�;+���ށ�]sr����x��2�˭���f�綫:f�����g+�ܱ�+��xi��e�+�����{Qe��Y-˃��q�&=�پ�=[,YR��wM���je̘��1��y��&'�x� ��ǲ^��y���O��=�˲Еۣ����n��P>�p)S��w<7%I���pwc:�$����������Z�E���2"��V�g1���wx�{$f,�b*�3f�y�6���緂C�����g��/���Kc���wڷF����ܣ�x<��>
�s�jn*EB��{r��Ӈy��c���#�H�$�90N�:t�ik��y��ɬ�g�k������v6��[���x�ýӝ$�=������}�Hۯ����Z-/e�Ҭ3���6h�&h4]z����b�ı�kG�*	�u�O1�M��^�*��ܐ����^���j�/d�8/����מ��
 y�Vu���w����N{�^��Q���d����=Ot��t4j����w��; {ޛ��Y����]�S8ý�5�W�{�#�{H�:��W�ˬ`-�=iyF��V���;1?�r�z���5H���]�=��<ĺѹs�rnt��!R��7��M]�3}���}Gۍc��.�`^#�./,Ӗ��2g.?�'��	��Oo�m�����G�؅sz�	��q�n6�|M���yaw��\Z�ۂ�~6�(����u�د8�b��,7��'�	�Ј-c�^j�o�	d̾=�/�sm�%��R5Ojw�=���)Y�#�K�<�6�Ss�YN��d���+3��]�۾��E}U�'�{���-��WD�W�"��^+�T�Yo�μ���i#�t{͎�Ӧ=� [e3o�O�����uTv����M�C��)�U&5e��l�z,3N����,�2���}J�K���v5Þ�� ��A��گ�[��wB�`��:΍3-iw��j��4��}Vn3�;�4��&���8���2S�hOql�7xV ���G{��OT_�7�������}���Z"ջ�3ڻsa�Tۃk[pr��*��$�5�oidz��C=6��.������y�^�xi��̋L���UK��S7{k���b��K��3>>�{u�t�vqq�An����_{�Ń0U�X���v�<B4�owFF�[��n!����~�\5t����e��F�5�+��n��w�X�Ӛ`�5��)�9�9�wx�1l���u��o��8�{�6�,�<��:�'��}�!��imD�2#�_p���N{zq�g��Q����[��K�gLh��[[�^W�rtǺ֓�����z>�g���B��x>_>�!�{��ܷ��35������Y�3�"؉��)O����v��#���-,̃�<T�e��������G�����V��|�q�r��78{�,t"�Kv�r|;$�µ(RѾIq���������n�>�ܹ�f�O܌5�{<��nV�]�p��^������m"��ʩ��zK��kxf���1���.��){Vj[�ws��r���YвxB�? ;/�7|�"�sP�3N�^�x=0O�������T�e��wҔ.�!y9F �ݺ�0�7��\opk���d(g����hb�m��@���De��`>��!ٯ6��j��i(ԙ�t1^�4Ǐw�O{^�\�u���m�n���8�e�3W��b�������1s��&�[��2U�vSpr��#�m�v��!��I�)��P�Wl�j)��ir�<f����}z��nud���=����:{^G�a��A���v#�R��r�愝��<�x:o�sz�y�-cxZX��</s�=|7��)o���<��{���#[of��/)��=è�*ϣ��k�pk9'G%�=ȎWj�<�5]~A�����t�F:w ��7O�1?QO޾����{r�4V�k�O�-.����Å��r�������a0�9��Ci%&<��zH���4�����aE�p[�y}_6����	��hx/��k��Qɱx�}�9�3��/g�P�U,��9��Q�w�)0�{f��[��ۓ�s1���H�6���W���,�_]���(Z�H�;x����}�5D���#<ͩD��|eS9���p�I;��}nn�.m��!�&���vA���Ta�������/:�f�!�*cH�vC��jt�ض�j=*O���B���(���Vv�}�
�=#	��n��a����m��gQ�ݪ���]*_��q]';
A��'�����;�T���T��;N;ࠌT	Ӊi�0��Hց��uD��{I��v^�y�u��(2Z}��E��!Vs�9���炇�r{l}��u�!�h�����_a�_���&�V#��+�x���~�e���+�<2�����/�>�sϨ��3�8���5��7̿�v��t�>��A�k�n1��o'����O��x�G������'3�����S��=�>q?6���vD�4,�
M�&/*��~Y��a�V����:�tz�F�v�ibd��	1(ѳ(�v��d�~Όg�8�0AԱ�,Bx/4�l���X�BK���r����q<@c;�ݛ\>%�d�T�Y�r���zufC�/�?&w{���d]�SAA^�̀ɓ�e�{��A�aR��cR[�E�}i���ƣ�{�`7oK��%N��}��t�_���5��OԽϐ�����M����n�|慭
�;k���gs��p:�/b��9��b��e��y�����/	����g��z���lѽ�bh��l��ּ�{<�Q���<�^��1��-��83φ�]��Q�w9�%%��,�ip��&�Rn>l6����oPW�x����L�1�&�,�úc��=o=-b�s�vX�o�>����L+��B��
�W����_���o���vnz���έ�a�V��۵�>�:��t�J�)L�n�X�3n�'x�i�����m����S;F��/�	��{Hר��;'��;6��Z���
�y��&�#8��)����s�o��k��
O���Ϲh9qi���у<WMY���t�6�
� ��{(��x�܋���QI���v�Vo�e4�
0t����jXx�5�it!T\<L��1�&�PX˭*���q{����#�n�Ɓ� �<0g��V��P�f�,���}J+����8r��:V����ZI�����*և?k��n�q%�{Yͻ ֽf�bÁ�.�z�Fi]t�C=��D��Ò��)��޾[��ݹ|����/�U�����hq��yϛ�k ��w��������z����0��8��x�j��Cż��}����+�8W쪣�����{��ћ�y�۷5��f�a�pS�g���9�M����&w�ד��߆%���L��;�#^X���\4<z3��'t����<\�NR��w�\����7�J�g.L}�7�tgx��)�v�Rݖn����ҵ���@���%1 ף����	,ŷ$}��M+���}�8�� �?]� ���:
�S��n&�}�jm���h1�{�y�츯=L��j�"�1����7	/yxr���h��V��EN�Ծ��߸��{o{!K�Z�5�Kۢ��h���q��|��~�.�]�G�O���D��[!=�{�rI�.��7�|���)��|,�`�p@`w�s������e��#<�a�ѷ��;���#{y���c��EW��W98����9����MqxF1������P޾h�'���{s����o'��5d�!�����O��'�xM�qxd{�yD�]��dG��VE\�wv>"�0�{E�[�~^�.�̃i>��ȼ��x�uݳ�����r&���
��V��`�O^��X�4�e���M�����41g�e�h��B=i�d�7������y���ۅ��}�^�4�*a�y.`_(�5l{������B�>wj:�צb�7j޻��[��sp�ug!�倽J'�'Yh�z���dgLԇuz�N�r��-�������}k��G9nv���O	��2c��##�8���(oΉhz�꘻��CPMO�[��S�Ϣа���>QglO�j������s��=��=�@��h�z�E�MΏ�T�K�v���cN2����[��{O�Ot�/Ec�w��bz_�4{����)e:!�N?}F{Lv��^~3]{��f��f.˾g�p[����-��Ơ�^�T���5��O���$�$�5��3C��r�Q�β�F�^;:��d�z-�k���z-Ҵ�%Ùn-w#�s*�9��"˱uݑS����.��d679.�u�崾8���g��u�d��	��۝��m�8���1��rm =m=�m�훋8�t���mƓF�����x��v��q��=�3��]6�گՕ�mnT7B]��w.�����p�糷�{'9��s�<@y%R�%�M�۶Lp�g>@PG���Fs����#'��a75��#�u�7^0���v����Ϯg�����lrIq�-����۞�h�Obx�zw���[m<�[;OO�۶v_]Ǒ�x���is�����Jn;x��˺hTPj�c���p>��YȺ񞨊��<b�>�9���v�g��vA�k���f�^z9�d�m�p]��S��&���r�ϐ����qq��;2����<*n�{�\:��N���+��o�&�wA���H�ֶ�d�݀m�1غ&7 �81n3Ŏ'��5�]���c��n�'d�}�v4&�:4��r�ܚ�nhP�mc�]'q̆�M���n���gzά�8�V-�:�p�÷$v8�n�Q���c�c9z�V�]5�cs8;D�8-�ůbێ�J�cdѭ���v�	��W%���>��]����;m۵s7��m�F��Ύ��t�׶M�i܍u�۸3�:�o!o/�<�:�a�u���G�q�:��;sݑ�3�c�]n��Ür2K�As:NX�㷁�d�=t���ʦۮ��:�aɈ���l�P�F9�ݍ��Okl,��U�.�ۘ��&��<��}�f�7��=���K��=(�����[H&nu'�/=��ے�:)�9���w��f:u�G�5�YON�D�nK�l�n��W7yS���N�9��N��2��
�s�\��]�LO�!d��v\�۝�s׎�7Y<4mN���:07cn.s�٠,<oFn�d��#&��ԓ��,[��ł���O.��͓d�nx�"�{L;ƫ��Ӵ���a�K60ە�hɫ�
��l�s ��x��^�:�^.J�'^�+I���,m)�t7�9|q�����Î�u�<ێ8����ή`� u�[��eZp�z*{`<8s!3k��Ňݝ��J�m�ݮcsq��y�Eѭ�÷��,7on7xd�woG7%�xۮ�����ыv���:��]v�ם���=�#�����<ݸOn�vƳ�8��kM�Yy��*/�=��]q䱕�����nH�v[�.<���pn;n;v��[Mcq�.��1a���&�2�����w=��<�6{p�ӂ�n3ͭ�^�W]��vۙy�ڑ��ۙ���X�m�y�@[���>H-�v�'m��nMӮ���{=��&�'�8�gf$8�IΞb����'�]����{feq�gL=�g0��'A�݉���=��sM`�Gc�7P��=����u�sW;Պ�Mأl=�X9�!7u�ۉ�孷]c$���g�^�y�9�ܯc��uμ*Ʃ��/Y6�k�piz��;���ۋk�X�N�e�΂z�o/ka8=t��I�}�C�&v��ݝ�CZ�1�x
��N̳윆7n�9�3Kn�Y�Ls<�6x���:ɇ�]�o<�%ێ2m=]���y�]�;s�s=�lz�z݇�K\'o:�G	Wv��%�C��tpj�%��2���I��_Fd��lu���]\l��m��ɪ������=���^�`�ֵ�=Z�a�{kh7��60�S��V���lm�ݭ��D
�S���>y���=�Y���9�F�]a1�u�m���\�a��e5�-���m���Ÿ���un��bw��V8�jty]��7ln���;<l4Y8���{�nxV��d�7�p�͌`�9:_/V��Y�b�5�^]�9ưࡳ���5vֵ���Mwd#[a[���wT��8Xy
�u��<�J�j��ɷ�����u�u�.|�.�*v.�Ӎm�ΚT�k[�'n��	-
ۍ���r�dl��ؖ9�,v
�ݡ����������{=8�m�g���k��qkt��6�	��㧲�㶐Њ\c��փ[nk��[jO������m����H��vu�/n����}�h�ܨ8�]z�9������Hs֝�9uѧ۶�vt��]�[��xz���^�{n�z��\����6ی�u�鍵�nZvӺ���WF��G\��O����b�t%��y��r���m�Ir�#jv�8��W����e�n7pG�6kn��y��6z�.۶ɂ]�" �;6dG!��p��vMI�^�n7C�,��p3�펹sh��ꨃgseЀ0��1Z&�/��u��ݮ�zƨQ�z�f�q�z�ۇ 5���Q\rW�Ȧ�KUn�m۞�.�<���O=s7�����)����Н��rX�ǎ�\�F�wx{�(`�5��9;�*�c������;�Ѯ�	ݠ�,�/3�j@�g�鮶[��AZ���q��Ԫ�l%ޝ�F��NS���S������1Z@�p��t�/������,����M�g/r<k���[�v�c��d{+�����ϧd���{<�2�cy7<vV1��e�ݔ�����.K:�\u�n{�=�U4��T�GLp[N��݋;�1��Yyϋ���-n:�N.��%OKO��ލh�Y�כvz�I�ݴ�9w\vAǺ]��ە�׮v��)�!�k8ͥ�8!��; q�Vfz������!����H)n�9�mf�zݴ^�b��{1ӄȂm�k8�p�l�d1�Z�v�����ݗu����k��gv�T��u>y�����k��mɒS��GY�U��t���0r���W�n�M��mڙ�q�go;��/�[pȣ]i�=t.�[Wg��[��*�t��	���m��xV9�Cv��e�W�� l����u�f$s۲hN���nyFIuq���N���غ�i���v#x�v����i�ݣ&h�Wn�V��r!V뮌�8G�ֺ��y����n0g�9��H����4����Wr�:��Y)���ې{V�qt�q۞���7�f���1�9���AQq����հknmqX�lH�Ib�����ѮKn��0���Mq�rwjy�ܾ����z�r�,��v�n�N{ݬ`���c{]���]��2q��;qn��ܥ�hyH!:�%��۞=Sֹp <��9� �j�p[����Y���`��l\��u�6A�L�s!��:���6�E�٥_�k�c=$�`�ܼܙJvֳM�s۫gvǴ+�&^�@Wc�=j����3ݗ���9�+���bz}��������i#f���;)lh�\h�sk<��,]x��m[������mk���t�tn���d��̖��Ү6�mWm��u��gs<�S�u�d�Λ[�o[��M��`;��o�V� �,(<W6 �5�n}����k���U��Ytm�vz0vO�[���h6����v'q��qn��܅tt8��uc#6C����qzvXt����Z��Du���N�8X���a��&��rqi�(^u��[ks���]f�g�,]pqm�<3Yn�B%�%�շY�@�(�d��u��<�r�<6׃�U7�M�Y�ȼ�]s��/D�\��6gu���3�=^1kPk>��	���m�t.^nl9�:�''d���V9��#���|�ۣ�����F�r�1&Δ�mc�&�z�>���q�l�sV{(S���Qܽ�[�}�6j��s�W<C����Y�y�n��C3�vla�չ��INq��܉ۋ���D��)�d|=�M�vq��g��\s�*��)5.��{]� 6�=�ee1!�[c���S��&5n��e���K�POV{su��Bj]Ъ ��&]������8�n
%<��N;,-�:��;d��69����nx8k���M<쩍����ݓs���I�k���.N�J!���ݞ������d���=�ndS����.�3�{\KN$��i1<�]��u���N�j���rQ��;q°k�Lk��l�;��oF��ʛ�q�$�^��{6����!���f��5�rk���N2t-���m��m��j6���=��s�۝���Zι��@n�m7�:��⫈�˴X�-�b���L��I��˸L��(���8�ͺ�Ƣ�qk�=��xKXe��ݣ^Оe��v���X�h�N�wnٶ���T�\�.�{v���kq�:CW.$���sۘG���8�$�ugf�tZ��k�
ں޸w=;p ����ñur����2�/+\nH�X���GSq�-�����vN�����t���Ŏ-g
>����g�c��qг]t��մ��t�yb�c�l�u�oE��Dl:�y����;���o5��y�3�!5=�5�Ĝ�1�1���9��{N��I9���B	p�����{=��TpvѮ��8v��3�S�[��:�ݍ�݇]�:�t�I^7�����Vj�F�m�/]��m�]s���� �k��:N]�{P�^5��n����g�6��hvݶ�{i����q�:݅m����.�6Z���.���XW�8�xmt>�A�4��`�xCKs�u��]��a��o Z�6�R6|��z���[n���^���	����|����u�.��v'�l�z9�:������%���ࢷb�A�6n�]gn��J4mw�m�wf�b�'y��Г6�ю֊m�n/t��l�槷Xn�whl.���nz�[�Vx�:����7f���-m�ZI�܌X����5nӵ����ꂇ^�t��]�井K����=d��<F�=Es��x�1�Ҧ�Fι���=]�{�v�Գ�6��w���;E�Qj�m�V�V�m
�V�6��,�R�����Cjǌ�6�G���vv;*4�֊Q�q�"ڵ���cb�3
V�-�2�)R��W��=�vx��Y�̩J�����b"�ij��Pl���˙,���DR�k�pL��[[Y5��t��R�+B��E���*��Z����(���x�v7:���;&�w�e�J��\J�����XҦ��Zi��D-�Z�Z�U���*-�c�V,�Vcn\PFP�*K��V��Z�c4�ո5�E(��(��F��R���fQSF��DkXԢJe�+DTQ�f���3"�4՘ʨ��T��J�2�1�\V�5������E�T����kʨ�D�.��4�ʔB֥j��ֱs3���uj�԰�F(�
�n�#��[J��jYj�h�a[�I��j����sJܩ��8撶�M����^ۨ��vv�)���;\���뾽�}8�=5�82u���V^B��mxN.ɱ�,<��n��{	�ۍ�-�띹���ŋ۷9��iM��/��\�unh�E�p}}Q��Bp�}u�9CvK�W�Sî�oӝ�y�*�88���%��:���uq��;yݫ{'+Ϣ���물��9���u��q��h�	��gm� �p��n�����;>���4����9l�ю���o\�Ǭ��Y����UK���6�:�ێ�n�x�;r�
���<��P�2'gBn$7;<�1ѬS��v�q�8�G�yN��Ε�n�ד��'���g�I:��x�W98�rŷ9ݭ�䵞[�;=�ϸ'��cH�ӷb�۝;;��q;���o���n�������td�F��af�8{F2Z�s�b��P�n�;�J�k�O�>��/�n6\h�kk��+��d��ka�(ӶS^g39�ttkͭ�+Y9� ��i4�7��ܘ볻O=�@���8�Mv����$�њ�j3հ�X��s��j����q��箜Ħ�9� �j5�t�Ld�Y�5��a�Î]�E��6��=�iz��7Gs��0h�b���g��`�o�m�=���x�ۧ���:�Vm��q�㳗�L�k٭��j����<%��]O�x�ڵ�h���� �#[v3�l�=v�v�;=��Odն�[��[���۸��<O�e�l�^7\���θ��n͝�(onȺ�{�M��m�1w5ío(4��a=qב�'��֔]���ݎ9�0m��<�:���c7`����ZF��#�+Ƒ]mm��v�q�H���C��ZHa��e�e�.��m���7pp���q ���WN��A)�(<n��<]���$L\맛pv{[q������te�2���N���ہ7j�rq�N���3O]U`�.�����Y͛ԒI������`���r(�GnM�x��9�a�c�nW��9;a1r�2c�����WlK����#܆���˄�r�^Wc�ۏ�����a�+Ǐnpp����q��8S���ù�;��&yA����98�<m��Q�m-*�h�cqJeS)�82�\��siC`¡�r쁻;og;�*<.�ɸ ��i����e�0�1�EN��߭�D��X 3]���~_����!gw!��� mvSL,�dLDR��*u$�>�A���{Dt�kؽo�� �F��8��dw���A����T�Y�o���b$-�N�;��S/�G�<ձ ����iX W)mg��߱{;w3�_GWe\C�;�逊�܊�8ja��ު7��*ؔ��H�vU�>i�c��۽���_��By	$�3�
G���	���L�=�~�@wo<XeFnJ�� ����;��@on�g�QQ��Y�^E��|���ۍ���Ë��ND�7�z�P�ܛ)��s�s�c��������g��u�y��6�#c}�Ցۼ�){�6�uV=��(j�d��-مUI%+<_s�ϰ��ߣ�#�J1v:��M1�3b�D�:�&C7��w��
?I����u���A�џ�4{r���`B僚'(Yˣβ0b~*�OWY�	 ��tɠ�{w����q�]E�*��f�R�o��Ip_�Pۙ����P���=��Wh��γ]�ϖ���O$N˗^H����v�9�jL5�RZ������'U���63�`�Dn��y� �����oh��:I^I�˖M ����8.2�.u�v-/$I���dJ��tk��$Ǯ�#;��a��۪B�K����Y��YI T@h In�uׇ��e�f➫mՍ��U�{^�N�%�VV��Oň&�ٞR$��oS�� ��V�	�A�Q��yKg���a$v�]�KGlF3�,�pX5^H��a��W
����g������	n�7� kr�d ��;�iR6�^� �u�UD�QD�RcF�y��@��ճ�?<ȳ����g�W���&5�M�_������c�~�2%��O�.H5���7�u].�
�L���3���O*���\�k�A#;w�=h��K^ۡIG��D������Ll:��'��w7ص�$��� �r���w�����:�خ������R	Ĵ#�A\_ď)^s A��e�g�t��1�6�,���D`��M2�t����*9��Ͽ����Jڴ�qxA��[�LsLy7[W�8�MY��i\2�}���|s:F���~}�c�@ ��ƭ�,;������&^���0�+6��A$�=�$�Ky��Oň&p&{j�R	L��d����}Tp  =]����˦��n�o��W�-%ö#��L�pX4Iwӂi$�lo�݂ <�p�wY�۞A �vSL�2;�t��vmETMMI%&4s�|zj;m��S;�y� E{��l@G{.� {w�w+��TQ~�M�C%�sbX}�y=�g��<5Gi���}���xM�H�ȟ'���*(��x+�@`,��h77�!��̒y)��B��e"�1�5������v ���㓿{T��W{Ԃ;�U��@i��Q�ݻٟaV�??�֎���i�t��Z��Ƚ].�n�v6ƫ9�	1u�2I�߿���;�H��)��2�Z�|��[JȈ���oo/+_GJ;�Y)��d ~���2I��D'N�Z�Akg?~�!8J�~���nK�̚%%�r�I%ݻ�~�PKg�|z�wޗd��`�PrϪ������6Tn��> ;ݼ�` QӖf.�ٳyJ�o.���w�����v������bP�j������d�<c�S݌��D��ɡ(�����l$��Z�o=SX��[�d��*��^	{�^�*���jd�����3�m=j�Uz��ڕ��Zvk������̄$����Z��:�8�4Ԧ���
x���<�p��i�sC��Ɔ�����|p����gf�?����'l���tiCl���#K^pI%5������WRݰݕ�9�����)�cd��u[����ٹ�0o��?A?^Sg��7��3"��K�������sє�8�o�n��͛�k�x9x��Q�wk5U�x$�t�-�����gF�7kY]q�m�fkF�8N��[,�ㄸ�XC�n0�������:������n�gн�c���֭Y)n�q��+��=����:�p��۰筍����c�cѶ����|��"LA~MCo$᧓��^J�w���%䗖��T�ndV��2VW�v�:�D��ޫ��c,�l��a��*�:�*i8�S�饞|��ܜt�l�V�X {������� AWf�����Wu]j�с3*jb������Հ��|� �WK-O�Ww��A��v-�K]k�F�X/ͦR~,A3EGk`�{z�/�<XD#i�[@ 0�7J��W��7����5��ͬ�#�fP�j�3s�i%����f�ޢ/�������@F�u6@���[��ݚl�&-Q�/%����Y��(��5�n\8�xox-���<���SmD6�P��o*j�ZI ���j؀�u~�]ma�Ӄ�1��D�I-w����r���1�4�u'L��s�^qĺ�uIɆ�m*���&ܹu>��p�X�q-/�=�O��h�L]�*GZǸ�-�Ი��8�蛿����� l�l��ü�&�������y�f���Q,�Ø�)�4��T�>�󺈆
��9��'������t��a�n�H���TDp\(e��R�zěfjZ�I^�������;��|f��kSOٵ�Ϧ3����A�>�*��S�EGkmX >A���b���M�*k\�� �w���A��Wk��l�ӎ8����-� ��\um/*�mw#��g&��Ա�`��ծf*ߟ}��#��fP�d���:^I��T�I$��{z��C2^�M���h�{�$��[L��oe�RZu"�ұ�}�9&C����enbT�w��� ���h�V�F�W��1����"& �&�n�����W��Y��V- "�ΰ�x_�i�Ou�Ȓ�k+���̴n采�����2qg/%��)^#���R�T���Me�"��N�E��>s�7�R]������u:_��IY�L�	�ު6!��"YPR�Ȧ4V�ʪ�ط��6��� Ts��a���{3 � l׶W��ޅY���$�K�u�:�I�GYN C��C..�{1` �J�:{�t�!��Q��O]DD4g�{1a@|l׶Ze�eO�*.fZ�/���A����`���P��4��cJ���f�;an��M���;��[7�N;�=)�[۽TI���y�D���+2�.�M�Y۽w�H-�#Y���j��s���%1ҥ�����E�����Ivv��$�Q{�D�˸�ȍ)L[����%ؤ`��B��������`| iY����}z۳7��'oo]�h���ý�5��#� ��Լ��C}�ݱ�e�Ǩ�/�[���٬�o�dw�׋�^����&�rͼ���ļ�_��+w2,"�.����\=n�;
�6֬��Y�OE��#�����b�'�̮:�/X\��'��������n�3SIL��M���d�)C��@�v�,�M�ߤO�?o �?WΒ�}��x`f�T�a��`>r�뮽���cbۋ���G���c�xb�.����~�2��
&�e�>}���J|� ��
+Y���>w��I'uF�F�dZ"d��b	�	��mX�7�%�\E��9�XD�ܖ�Ddw�������y�F��e��`#��3ꉕUQ3SDCafst�lo�ڰ@ n�dN�nS��o��4'��Ey$-v]:I{v$`0�1�d��}m�Н�ٹ�N�l�s� �t����쎴��.���@)n��M[�Eŀn��ҊO����8�ۼ�aV��{7P	�_�� �=�� ۽������:����۟��H�*_���ww��M`Pa���$�5�e���u��r�D�b�TL���Y�[�@I�q�l��v���a���g	���F�nǥڥϳ��ٺ�9�v튡:�g1j�ktk\���w7Q�DZ�lf:�ٶ.�u�;cs�&��9��)�q�ݍŧ��F��n��7;<�ś������v�v}�y���t�uU��s�d����l>�f�u��FCZk7n���g���Z�v��ۄ�=�sAm��nr&�&q��ۗ�,��1��GZ�d��:��]�d@�p[n�U�z�[���iƃ�,1�5uƆ\��Cp��bD4}	�'Vs� �ܷ`ۼ� ��ک}�֟�S�&�x��Lk^�&eMLMD�d���wk�1g���� x��M �;�{3{sж�s��ל��WE�!�Kd& �0sfpJA%�;y��H ��O�f�]��9���PI���z�H.�"0DÈm�h���.lwY�u�����(�Y��w`�GMnNO�=��unN� ����myD�3TMRc9�����'�N�A���#3�a�t�'sw��h��]n$�sN�
xLS^1�(Pa�%�/K�ZH��`�Z�[��gh���n Cnj�ƲIP_�&��హڡ(�o�y�� 8�ɷ�'��^����zT_��F�oc�}SU(�����0%��W��f����U�"|��u*�&��v��!�_QGo������/G��Ch��7_��{�85�/W�5��wF�����X����Li��"}Q�|��oV��C���\��γ����]������b*����Z +�m�S���=�22�ը ���n#MnK`e��1TET"���m�ܚ��~��'	���'�A���I��ﮧ/f�
y�[�ґ�ڷ���I�U*���!�Q�~����o����Q�,3���Dq]�������7s��f���~�`B�����/,��B�,yM.۠]�β��7<�G b!�+;���,8m6����ڻ�I+q� ���;��eǶ
���wj���Z($��}qT���I*��U�Bۿ;���r��8�9]ٍ�  Kf�%�� ��c�8�r����[�'���-��D1Bt��rw�S�,�e�� ����>֢n6j�3�Ԗ�{�4�_ٹǙ�l��-�T�~z�4�����q�kpz"��J���9�vOY���2����-����WH�82��e��G�'p
���6�{���������զ�{G�]ۏ��[ gjk�D��x�n$(G͓��x��>����ǜ����.�"�b�a�y�9'Y���FWP��]��Lxgy���KUM���~ٗ��Su�;��k�n2����F��doA���d�=���#�p[JC�Q�9�\�s�W�u͇y�#�?��9�)b�x*�ܷ�>Q��9�M��~U\�<�+���
$9,�p�{��g�^l�P��ĳ�����
���]�� &�{�Fn�:��'�vnoQݜ�L���/�Y�pt�*J��\�',�꾨)�`�4�����{�n_J�U&�����Jm`R�+7����ӤW�o�St��`�Ӌ��&�&g�-����Y�a8F�]�i;�g��vM�^���	�㫞i1���v�z���^.����=�}p�λ�¹Rn��,^�r�O\��dq�g<���]s���8�{P���zM3.k�< {��
nj�����轫�2��u����x�������=c[u�k�c����
,/+���}5�L��m�^�,�)��nZ�a���1spa�X�v��BY�K|��<;�V]CiN
cIk�.%�x��#ĥ�.��|��Q�vx�� t�^����Sͤ�����4I�O2�C�$�P($�!I�F���U��-*")mն�Tm[+T�T�ATF�kJ�ږYYU�muq�VW[�X��VҊƃ*�E�PUn�5�-�����J�[V6�Q���e]Z�ZT[em%�*��P�",J6Vi��TD�S6�JG)F�j ʶ��B�am�EDE��kX�$QF1kEjQ�U�DTJ��Z�F*�b�Ьb�ʕJ���+Y�j4�eQQ�*�Q-��m��V����� �`��aDQ����X֪�4T�3�IR��j�R����iUDD2��iJcUr��h����F9� �%�Z�m�T��Z	DUX�-�b��EL�8Q�E`��R�-�j6[��b88��#��X�����(V�Q�jҕiD�ZQ��J�X���+m�����%a[ab�U�´��m(�:j���J�m�(�U)K���MY**�ʕ��h֋m�� ����kkF��6��QF%m�,+
�AjZ�a\��b��
#�>��| ��l����`�{&y8)�f"�(�޳�5��ʸh��@ �޵L�{���wn󍇾~��#���؈	�}-�:�e��"�JbB��� �o7��"A�(<�Nw2[@�w�������Gu�[m=�;���6���Y0�ƍ����gnS�X�3���d�x����W&q�u��ߟ�N��T�U�g���� [��l������8��vR#�w��@�ܺ�Iؑ��,8m6��K���"�wۯ���N�{�V5L�{}����K�w��z*�njک�ؓ��2�<"b��(�vж���� �;w�,�	��������O�� ��˶�@$wn�ݥ�c,��� �0Ȅ�P	jw���Ƚ�]f��[̶�A��w�3�A%����3l8��ԩ�-N�[r���f�l�|���Ҵ騔n��s�J���Ά�b�[��l�Sr&����p`(�ذ�k|$��H��ԒGR�13�T�D�L߉罙�A�v:y������_��וV� �ki� ��f${�bgo�$�������H�ݛ7n.�!�0˞.KE�t�#�uub��rv�/����(��!���L �7ݼ� "#kr��;v���q���O�߀�����X��I>Q153UDCa�ݱz��ޙ��|���q�v�7�H�zkdv�mP��'���'Bo�ע&��MQU35c6��b��V��� gO*�7Q~��=�H�����h�u=��HGs���4�u$l������H+m��"+�m�A�g{��� ��c}��[�Sj�fI�P��Dq/�T��w��dl��� =}����MnKd��o���eq�}1��n=3g�G�y<�\������8�t�ߥɛ���X��H+�o�Q�r��޲�����B5JQ{�N�c�3���@Fe1/8�l����;�&�oZy,�=OV�w<c��L�vͷ�ۋa:s�b��/e�{M��T��/nw(GC�Wn<�<]����&�g�v���\��=��U�c�ign-=c7h��v�+�Nl�jՊy���Z�v�7Z�>�k�.�Ÿn5����=�c�Jv�f�e�8�C��������P7Nco��j����ȝ����ñ�nz�,f��B�vϳrb�&�B�Z�ںW��n��1.
j���o]�%%��ӥ�NpO�>d��v��Y������d0|�]��e��
bj�jQJbv�p�v�����_���a�[�؉^7�u4^J��)g`k��ܚ��\7�d����&�#7�Bi �#w.�`��2�=Q,���U�۞F��W�H�e��	v�L6���qĦ��y�d�\�(i�|�A��[D��v�ۼ��c-����"5 ��u�J3X�b ?&�n�闓�  �n�q~�,^y���=^�6�	i�d�Iݻ�D�-6�vxVJlΈ�B'R�]{�u;	í�\�3B���. ����{�"!C�-9\��z�#���> ��{3x�ٙ�g*�ȇ~_��d	���:h.�옙�pQpʊ�.u�tm'y�q��K1G	���%�u��v,9N*�ٽ����m�|�j>��>��\�@�4v&���� �Rm�"�\[�{��ݜ��ի����:��g	�Y��' Gv�c���z硓�X��ʡUR�S�EF�mY$ݼ�` Owx��|V���h=�u�;�yشtv#�Fp�h����Tc�tL΋/Ӡ ����a� w�{3  ��}:w�DI�Z]\	+YwN�Hf�8Km�n!�Tޫ�$ߒ:����/I��d^c,;|�Dgn�ń �|�g���؞���ӫ��E����i�f펝�w5�e���..4j��l�1��xzb ?&�o$ᗓҒI-�ޫ�@mnSvfgU콿l�/]D4�,�޻����D(~e�H��Y��$�{n����㷯l�w��1$�K�-{nI'���Ʊ�ڊ�Z�"�ʂ����pʉ�-u�v- �H�멢W��=[�\D����йr4�lU�R�W.������&�]kʗ��6�R�o��y�l9a�u���5��v��5.l"�&q�P��H�+�K�e�W,�	/.�޻�IIk�rin*��-6����j�=�P��N@�fzq��Ww�x���N!��{o��=.#OH�I�����#j �	iI�GO��/$N�˚�x�eE�d�$���wd�K�չM�$�w���)Dz�wѭ�LGϯ��[��p��P�t>oVۛk��;�K��\�K�̓ɷا�������j�,Է8���� F��[@��u�?a��>N/�d]{y��H �nSL%oE��e��ii�ʡ)���ھ�Qo�+Ν��` ]���{��3�j�y;07�s:����"p�(�"#����[�� �s�7��9��{���2�t�8ȬiA%���K�o]�Ȯ"2wg� ���|�{.�{w������gv~����to�y�7�H�7pw�9Ɓ������/�#��2�9aś'�ufg���f�v���j��kcY�l^<�UUOS�=��c�9�7q� w�6I�.$p%�%�Vhh�����s�y����y���-�q ��t�"�}�������	��$�騼�a�t���==\=WH�;\�m�!kQ���b����3��d�E�M�L�	�$�K���4�	.�޻���6Yn�[��@�	V~M�I?d6ƞW�7�3SUS4�h���İQ�ۍ�Okq����K��r��H��ݽ�~�R\$�WS6So�������a�h�[n��l;�j���x��ֽg��+�w��]��{0 7��3�	U��V��Hb�@�Z8������� lU�a�v�fb l���VV��zIMN�:$�ȮD���%���f` �K웅9S��F�L2F2gڳ2�4�]��wh�uN�I}$�7���iR��Q���b`����ro�Z�p�=���fF�թ]����y4�[`�'q�iG�޿pmC1��"j]��#t������$R��=��#����gD��;;\;�ƪ>�����:W/n�7���.���ЇZ���M�i۟.��u�!W���v{�8d��C��'H��<����sV�-8r��N[{HE���5��r��k�t����ڲ@�����^��KY#���v#�{gh���x�ok�v�qM�76��Bp����r"my�d��jԅ��X��֖����hy	���Uݬ�%z¬�6��5�'��yw͠a�. & ����%$��������&�Tz=A�>�ę[tɤ��n�]�:;�#�M�L�V{�Tσr��|N̨�*=N�� >v�vf|���M�?����*����A��0Mcưl���*>��ŀ�4���0 ���c_��c�	$�n�Ua$�'n$�3�Y��TUU;h�_����~����|�7�-�:}�}���0�Qޤc�ς���i@��%'�!��*KS��S ��mP���X�1<�1�nf ���M�?�8�\�c�wft*�2�dE;n��#�O�ӵݺ��.�����������A]ޣ�PB��*+�:��X_c� 3���"��&��p�_��	"��׌�>[QS*�&!�W�J�3&��q�����E�[�MK�w�������ە�|g(q�������`u-ؼ�:���&Y�2������1�� ��o� K?O���~�ٛ��Mol�S��i�p���00�F{������n�"1�WK�8�4L���D��=q$�J�2�	��0l���*�Oz��qE�����xɠeoM�v}�Z@ ���E��ɱ��'���[�T���� '�[n����� ^K�{����C6LO���/V�g���d� {Oe� nwu�����o��P�L%	��u¥��X���n-@뱭5uƋOa���?~<3%T*��9 ҳ]0��mP|[���āMs�w[h�z�(��i� �����6�~T�d���%���f` 5~�MKҺ��� >ݟc��#}�٘DD�ũ�%u��Goe���U
&��&*�b+�m� ��x�>�m���aڒ�Cl��K��\��R�<4L��G��͖҇��S�/꯳��5
_+˕���To~��oGNPUٌ��� dM�|%f�]E$�K���i-�d��ن�&�{��k_�U���o�t�������1| �狀&���[<��IvD�E{�(�q��0S��7R���Y'М$�i��\>b�����sz�Gn�<� ��Kf{�zⵟO���~��:vU�x�����G8cF�s��#�V��N]���.��p�W�}��ߎ�狭�UW}��^�@���y����K%���w�1�PI'7�k�!2�MB0�	���+sΗ���U���vM;�4˿}A� f�vdF$�{�i�|�}^U��sy�N�7{������A*�I���m��3�" ۞�RπAVEe4fN����	 K�{��h����`���hD���TLC��n����V�a{$@ �_kq� ��=��>6~��_Fs�w߁і���m�0N6v�F�z;������0aF�v���s�U}q-�J1��-��'�.;T�v��$'��[o?w���������!���.��`'޻9��]mw���?�f7�|�[�L��V1��e��hMF>��1�Xp�~�AN]���C���9x��we:�@\�1\��j��?�>?�b)�n�%}哹wv�'�7hE/$�;Ռ�����l�%=��o�$�_j�I��,@��S^[SU�	%W&&.��.�S�m�]Q��+�/�o� ��c�Fʜ��:S�U�<�^S(&�l��s�Ej�	 λ9擄�&�]o��勦�%�$�ۭ����c*��S$�UA-���u�w�r���i����D4����|Mϗ{шf��B��Up�Pᴠ�`�1�9�	x�f�sϰ�#�Y�nZ6b'�UOF�D3Ռ�h}�ٟ`�MyV���s��y\ד&����|��.��Q������g����[e���hU�v�ꚛ:���=����\��B�j&���W.��^�q�6Y�.����`�}���_���±�2J@��}(�ol3������V���O�L�3Q�z��R�#wۻs��I�o��B��k��[��m}JX�~`x�o�Ǫۋ�w�ݺ�n��stO%C��Y�j�]��;q�̅v�@+�z�P��m�my�:�0�ph]�����V?*�PЁ���XM������1�?R��Fg�ש[��}�� ����5ж�n��W��1���=����^Tn�����J��w��k��v�˚�.v!��\t���įu��7v<9k��ގ����E�䌽n9�XyT��T��Rd�Lόi����a$ԙ-W��#~�p�����5nV�=;���:�hf��p�eɝ��2�<g��>i�D��nn���sȓ����e`ʵ=j��n��K���;`�u������M�%o�������Ν�۷+�ũ�4�̇J�H��ʝS5�	^5�$�Z�{��;N�4�U񍾝�MoQ�w��{_B�Jk���}q[�y��9 OkQx������R�[���|�;�1�{�l�"�H���Z���כ�z�(�L�*��f�F]�Rt-��U*�ֵ�s`�#� ���=���&���gv��W�#JG�b!�z㳌�j5HXu�ǡ�*���tY(�/Rҫ�E����#EDU�A��TQ�Ī"��
�V��#m4�X�TDkA-lRTX�֢Ŷ�X�R�mډR�kX�6��Q�)���R�����Z�WV�(�a�F
,TTr�D�QQX�
�b�V�*.��T-��E"1�6�TQ�j墩*V+�m�R�*���բ�2�B�TX���-�b ��*E12�dUXڵ�b�J[K�()�`����[n-�X����s-R(�T�m��K��E��#DQ�*�*[V+�TUƨ�6�"���UQUEQ�mb��E���R҉YUTb �F�m�b�-++
��,A�,QVE��+���2�,���`�Z�EZҲ��b��Dm���FڤDQbʍ���1%,h�
Ȱ����j&6Ej[liR�U��t�1Q]SI�4�F(�b,
��+-���X�1R���F[AJ�A�EB��X������&��͑�M�Y�d�{7:N��-�f��^.�ugZ���F�Sy�*�O��h�r��li�sX���.73��)��]����6:��\��ռu����'.�	z��vn�l�=���TAE^y���	���s�՜�[���-w;�����j�7l�@ c�m�k+�h�ˇJW�����޸��@6zJ؏!�n��y�q���g�Ƈ .ˊ'T%�(����\6�=vÏ[j�ވW���]���E��)rsk��l��9��.7�'6�C=�CQa�ݻI��`+6���Ld�q���8�n��'l���rWQ;c���xWpne{%V�]n8����=ͼX�0ыTcU���tٮ��+tamNۑ��Y���=v�pi�9�*�G�^Aof���[O ��;'@�9�.���I���\7n9]t<[����c�&�d����<�v� u���Ű�#ռe���U��cX�t�d,��:���;�N�7`sp��=�Nx��L^:��{��r�;Z-^��9�1r�m�>�s�6*Ⳡ9{���ꎣ���Z�8�^8�75�3�g�;mxv�Ƴ�;]��:S�����8�nƱ6���	���n���U�ۛps��L�ۣ���݆F¢O=w=�J�1��v�[�֝����v77������-Ϩmm�v�����AN�:*V9mX�.�g��]�N��lٻ9tvܾ�]�h��y��y�6}`,�sV�����kIs�����܇ZU�z"�v��v��k'��q�ӻ��C�h⛝m��U:a*.6�d#��yu�d��ʐ�6;A����c]����:��֩��<��k��zy�6k`-���b6��k)���Ex����1;jz�\<�g�ڽq��[^�l��rl����'c���h��n5����%��:�Wh�5H퀹�p4�m���'��n���y�����X,��L�9^M�t��WWD�e�2U�\T�1�7f�������_���ۇ�<��B��{#�݃OZv�o����gxpu��ru��#WU�a��~�뺱-���>ޮ���k�;-�q��#��g��ӷ�v�6;]��m��Y�O�՞6�:�2{q(G�K�jٝne祻@���-	wKZ
�GY�v$���,�:�n{j�;n�������v,��kZ��H����̸����MkV�96���a|�ۣ��Gtv��;�\�\���l���ɜZ���|���\g�5�s�J�:�E/$N���D��gw]�.'�o�\��혾��sk�S�,�ZRԵc/���2K�s�)W���N{e�|g�����X@��ۖ��/k*�v����#��"���6���" ��� \��9S9yۜ7> ���D��̴�򤠚0h&S���8�t	롺����ϭ� ������u�\(�EC�f�y�K���Sq���S$�UA-��ݎ1�m�kR��5O��ת+�:��~�_��W1���٘@�:ovZe];�4�W�̽
 �o�{^M��{W\�ui�k�Wb�z9��T�C٨�õ�q�I%>��55PIU���m�$�w7 ��e��͹ƍ�R=﷝s� �����#�1D�E*�*��6{��@��i=�zf�Eם-������5O����D���p�%C�0Lb���n�E��f��I=��0��k�����=�<3�p������"d��=� =q31S�"W�C���H��e��{T�/�<����(��IU5SI�}���@ ��_��;յ����ܩC.����ݙ�$���z����(A�0�!��N�y1��*�ӳ���Y��V-���D��0 Y��r�I�����x��s0���E*��T��e� �޶�A]"a�.#��	d�mQ$�Y[� �=떂���:�}�Ϻ���&�;�s\r�ɸN��`�8ݸ��q:���9x�y��C����ȳ��Tg)�����=j��D��9h=uJ;����9�;6�Z)$��k�R;��Fl�&�&Lrٜ�H$�M6���N��g� �{V�,����?��VM;����K����,7	���K��I�6����&f`�ɨ�쿠Uœ��p)�˿C�m,[�7|��9��:s&����3mPj�/��;H����L�3u����D�<��{����f~@ ��4Ȉ?z}�-��R.)�i���^[=�wO��%T���A^��������>���i.����RGVM�^�$B%L)���_�^i�KsrkԦL[��$v�L�:�����Z@ �ݸ�8��&�{��}��}|�mJ�΃���%�������Fqp�8���i���{����8��������zձGi�[�A}�ݹ�6k�#&r3#�8j���:�I�Y��&�C��
!�Q4�����JεM��1$V��u�V�6}�,�3{���"�WY*�9�I=j�Fl��a�<��[j�� n�kŁ�	���򉥒�Yy>` z}�/��ݗ�ilr�cXE��6X5IJ�S�,���ۘ���@{�s0 >6v�=\-;�j&ť��$" E�X1�6l��.=8���|cER�5�aQQ�2{�����q�o�����\���h�3�ܜI�hm�������l��َʊ	!k��!8��i�T��ٙ�������;�� ;�z堈���<�"l��1���S�\=���Y,컌�md'�.v��a�]�s�m�16K�F�y���p�ܡ�����iN�	���  >�ײ�}u*�9ʊ��c�������S�X"�M*%9h5\�:Igw\�i9x9��1ے�f�I��{�1 �6u�DFZ����}����K&��ML�I2EUA-�����O���焀��`���5��޽�	$��ً4ײ�$o�ʢ"h�Q1A5A>[T�	��L<�ok/[{A �:��0 l��o���9���VS��� �����-V��7	�R�h,�mS H7Oz�.��^�ELv-Y�Ϸ33� =<�n!��=��[q����*�m>�i��0���;�<K�[�ғ���~Т��lzs�s6[��܆=�;��8f��?o.�鿈$��^bS1�eJ!���{uݱ�mŹ�^ݴl]j�z�s�<nΰm�696[�붰�	<V�K��vr���%v��C��;:�'�R�qΛyǏ<m��>ݳ&�v�^�*�kG���nN���A�V��4�_ml��`〷Gn&!��]���cAonn.{cb�n9��,u�γ v�G�.bv�*��Acm�L&ٻi#��`7F��R����s��<I��ݓV���.cՇr������Npfo����!8��i�_��w~�I:����x$�gO��#��d��z�j�D�f�, @ѵ�&�`�,(a��u4���Lz��V�׊k)��y�� t��m �K��4/x��7>��)�Ŋ)TҢQPS��L�t�����A"b�\��ec�nr�����I����d	��:h���U2T�$T�%�Ϻ��nrо!T�rD¹�t�'f]0�3��"mc���s묊@"�ߥ�3�*jJ**�L�)�l��m� �����P��NU��|�[@��Κ gwvb�3w��&�k��&8��lN�a-�mȣ�k��)�qˣ����:��,� �$��5	�Z�ɦ�%�M��JVsj��Dto�n� wwfb��	�n:^Ūj�ߙ ���?�;�-��%L�UE&3o���7;�9�*��}F錾:��u���o�)����{w�X˭%
s��$)3��e��b�2��S��/uHj"�F�{����m���:%�;�.�I#}�TM���g�r� ��[��u(/(%�4�UU�l]m�X v�<X "�˓��ҭH�k�)�I gw]�P.p�fi��s[q;��p�;1��qo��	��٘� 7i��U��'%u�2h�ŲI	�E6�wݘ�7����S����i��t�(.�I;�X�R� ���ÿ�7���K�n���<$ X�\n�݉^�g�p�cWM�M����?��չf��{�Q��V����0�i��]��������`�.֞~I+�����cMKf,���[� �e?BƳ�+b�'n�X| ��ّ�	��?��W:�+��������Z�56����e݋D�����D˛9{�w�~�f��')5��".��v��x�1��������9�zg5�~�vmV)�d�0��4]5[e���Z��3��=����S'<�����&�H-�X�RP0_L(%�2����a޺.<�b�A����`/�@-�~C�;�uuP�:=��Ԁ9��ZP.t���-��uۉ�I"p�dԭ<��<�!N�$��컴�K�u?�ý�M���آ#H�*fbq����ͮܵ�)>M�
��gb��C����˪iS3ܻ��!RL���O�<�ۙ� 7���,@G{�L	/��K�ɿ)�F<�{� �~`��Cʙ����U���f���_NK��Le�Ǹ ��6� 2;޺`������ٞ���itj�	�a�ن��&v������� �>��*����c��ڀ� ��~��,;�t�S��Pড��b���;�+|�$�ڧ >�}�O�;���;5rˁ{ٵz�;�ub�_o�vոb!��T^\�g���h�TF��*U��\�Qs(W�t�����(}��~�[�'C��{������q��T����`R�J�UU;b��[` ~��x�U�j����@9��������� �wvf�s)��a�۩SS�E
`S��㭷\6'��w��-u�֎`�U]q���j~�7ω�[I��,���KU���I!��4)J��w]ߒ�.kN����t]\P�RK�32���Q�BN@NN�K���^�y�W��l�ߕ�������I-���IV%���2�u�/#za�L�LUB��Sm
�[i����sϰ��Yď�O��S` #w�v�Iy$�w]������%��o���z���vYw� +��� ��{�1���Q���K}��ɘ#P	��U�E���P�e�1��e݁i|�~j�Dz��|,��w�{�v�(.�RD��9 ����Ġw|�Y��_A>�ֺ$P�o�e�3��;^>���y߷zxl���.��<S.��������I$���Wҙ�����Y�^wWn�����x�ڧv�m��ݗ�]�Q��;	�wx&�z��\�rf1{z4�x[]��>-T�/��.�US퇌i����ǯ<���b�.�1�W�6W����lt��r�ζ/gn-�$ݳ΍����-�pg�f��u��;u�S>]�L�����njq�+��N8z\���A�L'nn���j"MGV���]���$ �/=�������3�/l���C�8y���߻��&�!��~NN�
H$��n�������\�^Ft�o�*�� f�mݨv�C
M�eD����lF�FD&�wu�R^H����d�H���i2��"���9N�[�� �`�D�I2��E[9�vg�	 �7��� ��#k^۳}S�$�����h��Kv�ש �	�q`�bd��3�o��[���5�� �<��F���I�H��|m�:���w�z�M��Ѿ�Y��&�-�l�j�H�mT�I-�z�2��/�(S�K���0A��M� �;�v�w^�݉察��w��ۭ���9��.�qO#���9�e�)n-+����������$���������I��p��μ� �k�Kxߪ�����N���"7_����W}*�KĒ|�y��d�"�p�n~���&��#�yۚ/�g���s�fq�;wP��U֎�m*���AVg\_]�O�r�ܷ��y�6g8(�� ��f{"	��I|�t�����G~~�` ���;` Wϻkz�hQT����k<�mL�QJ*	r�i�����{�� 9���uWN����H��w�xI�������wp�.�q��S�������%�^]
q�Fw�����}�ٹ�๟�C�z4����ڊ�]�յ��a��6Tn�Ղ =���`�.`��e�+��K`��:` �wfa�L{�~p}�~��垟^���KkD�h7%݂���EN��x8�yy۫g:���~�t�n՚�Fr@���$�[���wvf|��]M�滔��6@������'v FApa�i�ؘ�'��v-,�|�Fk�^M禉I!�Y�N�^I.�PKo��F֚L����K�f�}�&�B��v�:�X ��x� *���"Mm�3�7"�D���E���Nz�NfH��%=ubhMʔ�`�'?��|g������p��6��`�.q��/�fT	�I�}�&�����a0����1_D�xw��x�����-j����o=�sOh�04C����KB��<�8.9Ӻ~��h�3Դ:k��׸���z4�˞P��	໖�*�-6l-Z;�d�4Rz�������ub���}^"��#Gc��l����ݑ_564Ч�G���F}�1��XE�'����|���gT}\����N�͛w�'�nm��C�=��A�E���[�t���pp�Ci�W�v	����E���[M���v����:>��@�4�t�v��Űz���k=�;�_l��\|��IU:�pH�0i�!ˬ5���3�����yx�������g3J��TQ�rJ��� d~]��_)�݀�m�$/N躃U�7����_1C�J��������by��{o�׭O9�۞���9��[Kk*rTEJ�tUkPb��יT��;}�x��>aH^Pn�Y�W=$�B�(�e�7~Pּ��Z
q�)�}�y���P0Y�����oF��wpy8}�ߜN�Ż��N2}i�;gc�<��Qv.�$����>�ղC����#	�;��B�r%����~��_�x�sɕ����t�t>9�eq�/��P5�!�f����Ưv�xz� ��e"�7x�4j�xo_a\�c�����uְp��E2��,��P�DjJ���A����S�`��ZѪQ"*�\ɕ±1�j�[���
"�1�&�r�m�dDV,V(�[�U�J%(�Q-�b#D`�����ڈ��Ub��"84�Y�j��j�Uej�p��2�Z������QTjU�W5�#�Yq(��LsV�L��Tb�L��%A��Ո���e�Q�\�Re)R�����*VEV�PJ�b�����J�5EQImuk�Q�A���
��Z�"�˙QQH��,�b�cQ�`��PT(���X�c3%ST��l�
�Ŋ(���
ŋ��f�����(�dEHAJ��Z��J�ŎX����iF6�AbZ���DE�$�J�X��ZZ�QEb��5�X�eeE�֬�b��JȱTR�*�R�JU��"�IQ1U� V�4���Ōf
�UJ� ��+F�UH� �Ԩ��j�q)e�5(���"�*������(���>����\��%䗾[�N��(.ϻ��ü"M4�eEE����Oc�k�f��"�m�`� �ovf  k�Fa���H�*�:��l9��=�F�'WVDȗ9'r��c]y.7=t�@���XA��~�ɍ�}C������̹�~��J&b�4޺^�]����=�I��fhn�S�$K�����!G7:��|Tz���������N�Ka���姫ϕ$m������ۋt� H���	g��L�l[}h�k�������ox�鸇��,[�֮4���>|Hx�FApa�i��r���f, i���L� b����]x ���� ���i��`*�a6�SAi����\L��Ti�L����o� �~�� ,;<���r�����$8�5�g%�}�i~�^̬���A��ۃ��O42��UBS�Q�)�b�6�j���ʾ����$�s]�~����D�M&�h�%�2��������fYUye�o��w��3 ��4Ȉ����KIMLS����O{A�O�AGD"p�x�9�uZ7On���zt�jw���Q�鳞_���>w����*�O���ŀ F��[H�t�KN2ҪkfH{����<{���l>3S'&Bd�1SED6Tu�d�n���z�e�%l���o�SP
3���p���>�ꬎ��q��1DBl��M���5�U4J	�ɪI! ���]���={�@|��i��ד5��q �a�i�ب����/��J{�Μ��HDE�� �-���DC;�ݞgs���.�}��^[����a��d6��93���K�.��y��zm�v_{ʈ�7yN!�g���� �v�`�2U-�{��j����[��wػ܇b�A��O����5u�7��P���Y1w�z�:�)�2c�-��0Lҧ��� �}B�ND¼q�S��ݟ7�z\m�ϓ��o�m���/]�Sm.���Rm��~���wu���ܻ���p��'n� DK';�%9=H�yٰ�lxv�\����'lf�R�uۥy7�D���
��瓉Cc\U<�������Z���N�*|<�/m�������`#���4�t��$x��z@wnn��F��v
:ꀸ���{Ok	�ꋝgu�S�B�q�:��J��ˮ���2W����q���D\X~���zձ�.���0 K}ݹ���1�����2	'0OZ��r��	D(	�b�S�OUlk6]�L
=��+` G��;a��y� ��&�k��ù}�)�Q	%	�[i�4�;�� ��x� �8�ySݷW�G��v� �ݹ��u�&biDS)�ª	�������9q��l$"���Ȁ����b ����Q4TbI9YSI>؈7�Cp[b]y=�����U��WO���{�F_�� #7�^, ��4�ۨ�~��Q$�ѝ&]�c��H��;n��8�Ѷ�e��q���M5;��0�l2o'��ڪ�$ H7w���@��M��c^]���3k���&���W��tlD�!�iQE*�K��z��j�}�޳1yYp\ҋ���w\�`�U:�����6}�o�� ga�<p���o���މJ�"֒D�ڪL��{�� O
���ȁ ���ky���U�4�$ŝ�Ѳ� �ZmhT�j@-�v�y������ g���Nq3�O���DF�ݽ��3�{s��#5p 0�i�Ѫ\jv��������N���_^cq� �y5h 4̹YUٛ�;�&6�^_ueݬ�YaD`��a���C�ul�ѹ�iY��_�|��z@]}��� ��U�4����6s_'3���������.5��|�\㴜�h�v��wwAm��Kڴ���Vpfo�ߟ��՘Y)g����I${ҿ��p���ɓՄ���w��[����f >��\?��!��%6�SAIͪ�J@%쌕]���.}Y��� �vz�!���t�$�gf��_M�W_z҉�*C�ˆ�p�h#���b :���<�����>�rC����7tf��x���)�&�L�^~=Y�Ƶ�W����w8��6tz��b`����M��(ٱ���hY;�GW}�<<<#��a9�?vz� @}�~�����U2���Q.9��nW�j9vz"PFw��| ^�2k�%�����$tLf ��Ix%�<��#' �QED6tS�����y�s�ϥ��A<��M��%���0 F�{ٟ`�!�"+-t�lDB{��Y����ӱ܍���ѵ(�a�n���N٭آJ�ǵ14�*��T����ݱ�Xg�Y&�I�컰��sN듚��� �{M&DA��?���r"�QS3R6ĺOo���AoE<�#]��kث|� {{��0(�Z�r��u��r��,\'��o�ub�'��|N����ʻI"t�����Ǖ5���f{�"/�t� ����ޯ��0�(�����9�@C�	$�ͻiXA���f  A��TM�c.jK��;��[��qY�6g,Ӓ8�Y�k��L��c����Ynt>����:)ԉ0�CD�֓�p>7�2�c���xxd�����e:I �6�T$*e��@����f ����������ӹ���|退;w���!�x�R��
���|�Ģ�M'
���t0�r2ɝѱi���WaW�q\�FΛ=M��%��dE#�m�!ζ��K���y� {s��'�	�'X��K��c�ji$���ʣc9��
�f�F�}��!���J=Q�� n��|I$�Sd'���v2Ć9�=��o�r1E���6�3]U��H�#w<ո�����Pr���~�{{٘A�=��i���;�LҨEU]�_����p�+��_�0/���a$�J��$�G�k�%do�X(�zi'�3��v���a�Yp���OS�h�=��t�*��z���^�s~��&�T� ����i���m�'��^�=�@����|<�{��T7=����٢g6:3�x��
g
~��~�O��0�҂�2Ta����z��\�Σ�!��:Wu.en[s.��aw�9��m��'d:;m˵:��kmۍ9��;��DG�`��8L���z�����v ;v��M:ێ1��[��iL��;&�;�rqˎ8�Ӗ0^���l�c�w78xۇ1Մ��ǀ-�Q��p�m�L�,y-�dм���;`E.�%��&��ݵs̛C�v�q맻��a.Wj�lu�H�9�=��rݔ�������H�[8.�t:�q����v��I��W_����c�D��P?��=��7��[ |����u�y�qQ��4�s$�������594��*�l]O]�
�[}�*=uS�ٯR� ��8���?;_ ��Uk�߽<G��n�Bo�n)�&������o���ݰ�}m�Dc��t���{o0"�og�� >�v�d����7�wRВƙ^��]������]�$U��I$����$�ٽ��]�$��8�Њ���C3J�T�_�����<X��<�����~��!y�����f,8�x�,�*��6 �N0�@�-�.��a�����Ԛ�Z��v���=����~o�,������	�^HmnL�i-��&i��{��u��2��3�+ԉ#��>;�
�"QT�qϯ^�]�����Ov]���p��tD��0��ݘm��suSE%;�f�wc��u�[r<���Q���4~�~�t=(�3����4��S��߼ � \a��� >Q����#�����]�v�������q&���hE���U�S�� ��y� [�7��:�i ��}�o� ��o{3�=в�D(~-�pZS^J�m;ڍ��vg��D-��i� 7��� ����diSl��7q���wq�"��� t��lS�'��wiy$�����,��oFf�'�U��m �3���X@�<nzk԰<�Wж��GA�A��$\R-z9^R;3�p�Ϯ��6�xw!�^E4�Gg���~���┓UL�]�u������ �s��-T��_S�˕��w� ��˱i2Ć�e�p�
*	�Obp%>��������Y2k�$��7����[y�NHș����u𨚮���I�	�P�瓀�j�z&�]�쌎Ԫ"N�39������ۍ)vca�&��F��kI�0x�Ϥ�I�q��o����sF��lEA��3K[�Đ �3���_}���೷�;��?zi�R-��M�]/g[��g�i8(��ɼ��$�T����GvVV�!OsS5.�V H�h
#:Ѕ
�3JL��vmd�on�;}KN�����&�&��Ē	��ʢ��r|I���$3��厮y_)�ڝ�[Ǻm�^�������yn�]@Cp�f��Cfm�HWY?Qq��}���0r�q�:X'#s$W����%+(����=ɜ ��cb��P�p۬����D�t�\H'���+(P;2�gi���!0w��칩բ�pla�i��Q�� ��$�`Em⢽��t߉'ڧ�'��{����mb��Є`B-�z�v�m�ps��&��2A���I��Έ<�{svǝ�ϯ跎�{ܧkM{�k�v�=�7O{ޮ)P�˖�8���G��尿��mA����[�<�d^Y��������'�6~���f��>y\�۪�i��P�N�	7~���Z�p����9P'Ċ��Of�J�����������,u�Cp H@�'�ܶ��Q�
��t/��N�*u���r#{6��紞ɐ�$ͼ� �;7���@U�gf�bo����	���ῠ��4�IKPZ���}?>�]��q>��Ŵ`�~�� �� !����v�x\kO\Y%h���(l�!�#gv�� ��eQ ���6�>�d�w������@N��M��pl��a:�t��qΣ��nm��H.v�h�@;��5�E���Ք��(�������;�B��`=];5�N��;��֞��$�����I=�~������?��ǭ����]��,�e&�Z#�d�������5�m�H�h�����0C�pԨ�ql����f���>{"�wqy�H��W0
�'V���W�?�vb[�0���u�������m��R+�1��s���68�;���b�z|-�w]�=O}D�@�u��7�DF[j&=^�-��%��F{K�n�?��k�UnH/G�In$[F.}�5���XO��^�s(ju���ޗ����cYx�C�x=3*E��ǵ.�V=�"�X��nu��P�:�5Z�ث-�CǴ�r�('KV�o�����M�ݪ�zF��Lcem�ϰi� �n��bT�"Xǔ��J-�a�y�v§��z��9^��o�[#��4S(̣7ZV17e~sZm��ӻ�udD̎t�s��<Fc�8�!��Zf��J�
s�8��b�v�N?o� ����*�<��&�d�/GI����������A�/y)"��i�{Ixy����U)X�3�\L��Am��~ȸ�C)vMA ���߾������x�B!0��8A��~��<��f���=P��g��Sz%�G��v���`;���Ű��{ԑzz�=�6oX���7����=�T�ɣ���z��}����Y4Su���.�F�/=�?c��{�J���Ygtk $C��RAi�����2�$������M+��Ni{4CE�xV�j4{�|��瞝��7\�[�h.ލT�c��zf�/��wM��V�ʕ}�묲�n�v�lz��Ѣ�ʩ��ٯ!�,!���k��*��}�=��~M�UEU*��h�^S=iL��P��Z��A`�,��a�ZTe���8���B�b�9�UkD�*�R���W�j�Um���b��4�R,A�TD�ƥTP���jR*� Qm�*���em*Qĕ�R.%�!X�.%U�Y-�Ab�R"�F-��£F�,0�l4�ձb������X�U�:j�Q\B��TU��Dq���jfQ���P�V,*�(���[AkV�4�"�*���������iFj�Tu�hV*$Ģ�rب�
 �(\-q�Kdk
��e�(�mU(�E""����X�QkKb�*��DV*ưK
0Kek`�R��գ-�`��ulW-b�-WY�ZV��[P�±b�*�ȫ+*�cJ:Kb��Kh��-)D�Zj����EH(i�A"�ZU����T���e5J))b��+�X[�#V� �V���WMt�f ���5�h��W-ueb�"�T�LZU%�E-h���~�~�g�0�uڥ�v��v��m��og�v����.뾋����p���5ƺ� �v�tS��!U�j��,nn0K7%���r��Ӷ����ճ�u6s�5ܐ��d�9�خ{e�ns��L�o:�T�wn��d*�We�n5�Jݷb��.ϟ{c���G;��6���s�މ]�̶��O<kF�6ꃰ�{wG.���ѷ\����.�l.랮Z����s�B��;U0�[N��'���Iûlb�^���e���n����^\���#����N�Op�wm�pj�V�v����8y�k��֪@w-�n�&�V�Ƭ�(Y�U9���b�a��q͇��Ɲo8�/bN�r]slԝ�ڨ��c��4�E�h[,ܷ`���g��s�V]�R'7�\[��1cv�Z�.��,��n�f:Þ3{�1���8�����غ]�,2ˮn1i���q�oe�ukC�����������ͪ9����q��vػ. ���4zWp��띟(R$$h�bx�yK��9�^Ă�m<��u����9̫9�q���N�X���y�]]gt�������e���Z*��]۬6/`:�N�)���h�ܐkjy.n5�]�뷨.ݤ��v�c��ph������y�@�����ծT��^���%=��L�P^���V��1z��e���<�q��[�sɯ�hι��[�*F��7�c�7��Wu^4�/gn'����ۊƠw���6�N�ƭ�Y����vλj�"�<�l���cn�W�Bm��S�����[��O�ۇ�듦�
�\fLT��o]g��6gw3�J��lN��q�xn�GN�/�E�ؑ��������9�)����q=�y�z���˶f6睶�7��H�]�teۊ�uX{��N���k>a7��ڷ���pb�m�%k�F��	�m�9M<���wv�l�� h���V��q�e�:�U���s׭��nS�L���E���p�+7�Xr�Y�@!77�)�\rZ��WY���u^�%.	������ӷ[={c�O�>�3���k���$���y��G��h��;�[;g�<s]��渐ݷq�b�f����h�U����	=9���A���n�X��q�]ŮX�ob-��<���Z��ne�M��{K�A�v�&�v=�a+��qg�N{�:9����맻��a�y��j��-�j�mʯh6|�cs�x�ۋ@�����ȩ�-mE,��]|������tCj��#*z�|s���A�U�Kc!�TE��6��	�{*���t!B��M%��8z�b��^fAG��"�Θ0a��ɠH&�UĒ��7�j���6��Le��b%��N���pQ�'NU�>#��k5OE�
ood������%X��1 �l�!��vf�V�Q�:����D���� �e�Jv���qmGo��:�-CC`���i��`�}��ry�/J`�w9TA�U���	��ʠy	���ھ�2�H�$C~np"�.�5�+��]�#m��q[��q�v;5��ۗ�+����?�G<��6q��٠	8v�Y �Gv^U�E��]ˉ����k���]WH�� ���b)j���o ��پU��N~�ɼ��溮�)͡=g<\�(Hl.�S��٥Oz�臏G�F�f�����/#j�mf�Mԭ��M�]T�=�������H��$�	}��(iln���Μ�ɬ�WB(~��p�S�'�y`��� �G�O����wտ����=�yB����,4�p�W����S\�˕pH:ĭA�y4>=��ʊ�ߏQ�� ��/ �3�>��Va)9;�T	� ��e
�.f	��j�v H��>$᝷�@�I��ʨQ��sG.6�z^���z�V�f�X��YqtY��æ ��svQ��2Q��ߟ;�6�1�]?7���Y��y"����.���Mծ���ו@�:2Z�P�$���$T�}!r5p�*,��g���_u�Q �{7�EWT�£ݳ�3+z���Y��n��uN�f�eQ�jrԸ���=vfbGm��P�C5#&^�]Z�ڧxe͑R.���N���we�Κ�R��i�O(�Qi����4 �;Q����L��$>μ��;7�F�Єb�i�M)2w$�(SlΪ���>ݚ��H��TI"�U�fP����*q3c�l�虥 ��Ս����l`t�\��bmY�x�x ���@����񧵻�J�5�d�E��j�5�`�3�9�Oc�]���Τ�<�Ѳ*i����A*!���l��Q$���eQ$�YW��"o;Ud;�[AM�Я���E`�!�4!6U���g�мge�G8Korda ��ݕ^ �ʸ�D(~���vn�	����-�AQ���Ӳ(;W!��{�ɉA����H��q ���Y����z+�i�޽�M���'�+hQ�z�������C�C�0��N�9r��HsG%΁�N1��w�����y�G��ל��������j�_��tAY�u�wh���
�?{����̻�#�لb�i�M)Od� ����n*�lf.������T �]W	 �[וF��Ù�h�;��Q��H��!�ǩk\uڮ"^؍����tLK���a�Q~����%��N�:��Q��*�3�A��ɣ�3=bD����M�
��j�A ��������A.��#o����p�O��.����޼��#�}Ow�W�5�vw��CD2C����EW��Og��v�M�H7uHn��@��iڸ�F�^Mx�ђYL��!�1>=]={��=��M���3�A7�yTA;��X����)T�H�3�mi�l4���{ngj������K!�Sn�į'0H����2�ĂA�ok�>�8�=�p�k�>�uH�˱�ڡi�G��8gz�y�}8�}<�vP�(A��6i���r�(����<�����m�wS�20��{�������@�m���Q��8�.���v<=]�A�n��y7d���nR��*�����{t��m�W_\o�}l��3�W=�Y��!֧�u�n#�d���[�<jՃBoJ���Ͳ���W����'�xy�M�l�t�����lۄ3]&3��^Cg����F0h�4��=�u�qk������v��.���0�;V�98:�9��klu�M���p�9����%˚���T���f����?�3[�) ����l�d}��(�;7����F�)��ߚw�$ݬ� ���6!�,4�p��1��4M�Ҋ+c�9�A �/6���A�������{��+-$ DC�n#�&sĒ���|O�E��x��f��.���W"Ay�TFA�!�5P�i�����V�bL>ښ$�ٽ�^$�YW�Q��S��[u@�gIe3R�� Ğ��� �p�\��|�ɋYz(.<'��U�A ��e
�YWF�}jM�=�2p"��n�%K�l��'�K8褐��l��jj�4��]����pXi�g���I7{*�$�ʸMl���j搞�ʯH7��@Q����6BM7	� �ܘ�^:�_�s��w��q��F����� ���[�C��I�u��k���+���C<|O��sg�Q/iG��g[�(<�1�������*�$�YWIs�j
��ۻ��Du���8��n��1��5�@:r�|� t��#���g�7��B�6r�$
�tZH@�� �n'�v�{[��F�ӗ�����'ǻ/&tQ��ܘ=� $���F�܍�-�6�P�1��$�\�NI�� �wd��d�I �;�����������?���ma�c��F}+���D��vu��]լ�1�������|�B�Vx��{TA'M�$�v^P��m(� �MРI�����.x¶�7�ꝡE�c�S�o��hN.�� �e�� �����G������U�Se�M)N��$��m�׉�3p�]뙖�ޜ�۵��-������:��n����7[��,��m�1�m���ˡV!�G7`�Z��������V�-��9�Ϳ������q�Q� ��yTH���Xna�[�*���O��2d��H(�\��A��ɢA �wd-Κơ^�X�H�΢A�m"�!���ڪ�;w����e�К+"���{A>��ʢA �weNn�YKV���	<��=�m��]��{%㉬\����bl�����CL�JqZwGAaڂ�P���Oy ���0���yw�o���������I��ʠD��-&�
J!�b|z�mQ*b�oT��5���oo*�>$�weP>7�w��OF�n�q6�U�m��Sm��ꝡ^#7�*��7U�]�]�H'/�*� �ݓ^�B�I6QN�ғ'rI[��Ct�Au�sD���U>����<�s� ����3Ѷ畼{�U��^z������I�#�3���[*'�ċ�
�l��j)�N����s!U_��΅AB���$8��AL�����Ļ�����+E��L4�p�q?�c��-����������q��ݕ^>7�nN�\Է�͕@�]ɵ�v�H�8�p�Ϯ��Ů3�ٱg�Bc6�0��ӈ�D@����K����{+�A$��M�=�{%4��:�ʢ=��^��r:��څ4�{2Oըk���[��&Ϗ�w��x��ےAَ������"ll��q�h1۔A>#6nd��������]O	���� %����j�qhH�r�s���쉳�g�gVe
��t����;9w{/�,Ę��^@܊�M4�m����D�d�H'ǳk$jlӋCY��$lM]P$����7����{���t�u;�>�+��v�ƨ�ݍ/�Otޖ��<si9�B���X���|C�Non�_vzj˷7(:oY침��U�Q�[�يG�x���2s�d��9nҫ�"v�у�Yv뙚��r��5�o��W���n�6���u�&=;��ęٷ'`ם�u���o*�M�E;c@n��Ʈ�z�1�;;�PH�<d{M#vvm����x��O��Lt��n:�7S���;�%�5��N�z���8^��&lb�����2[arƜs���Nx��g���ap�=�F����]�<I�+솸�g-���nWu���-:[-��u�I6�v���4a�-���T(�GVT��VUx�щ��~1S[@P ���$��ȓ~����3��XxVu�u\ms�s���S�쬪"�sq\�s��'��7�`�	��˃Tݹr	�k$P$��GEZȅ5ٛ\��\��VUx�gFĢK�0�C@���zw#{�0��*��I���D�O�o_^m�n�ܦw||O���r	�}IÆ���M�j�S�D�H9�}T]�܃;z^�!x��9 ��n#���������q�X찉�QGW��^'�������;f�\�<�NG��Tvӳ�p_n��Zi�T6�4����I;�Y4A����ѭ6�<vn܂MwNMx#��0�አczn��v�=�qGc��Kl�v����q�g/�@T�$�*��gS�c�v?��x�1u`��,3��*�{�^�����~ 2�~I$}�9TH$��_P�A2+�b�-�%`a����њ�H=�U�|I�����H9��@�����1�'�{9T	#w��Q�]��0ل�pj�F뺑����c>Y.�W�'7��Q ��2�N����)�ڠD昘$���Q'��M�{"d��xs��)�Ԓ^Y�|"k��g_W�O���>%����<R
D-(Ec	�.�v�7)7:[c�ۈ:�E.����.��~~�p��Sm��FT�Q�$\V1���Ұ��A�`N^�e�
$�u�z����M4��چ��4��5ڊ�'�t� �7v��ď�c�J�E_:��ĚɱQ�V��q�b��7�<`}�v /����=U�Zw�%1�]���d>�Zkۭg�;R��[4�;��I�E\��߯N�7�,xgF�Q.=|n���ݽ����gv(at��;jrb��Bs{�M�U��g�25?v/!��<�s�ד#]�&2��+�n7�o���	;���[����}T�Ӑ��ig���Y;_$���i��9Ӄ��ӡ=�:s؁�}������F/[ݵg��0�
��%��؞G��|=ҭ��7�ڟ�����������A���< �C˻������+�y;y5�Ⱥ�D�/�����8E9]��]��C�!|����n\~(���<3�]�
����+!�.��]��΃}W�}q�.�G7���Z��Qy��t��_ q�%�W/��[�ӝ�=�S͉7+�4����z�~=����Y~o��r���4�;��<���eo��ZF�^�d�mJ\���Ʌ<EW���[7���*cGݞ��=�ܩ}ǥG����-}e�l�n'�-]���L�O���?��?6��z6x�7)پ����4�~,�����5���d�(0e���x^W�aݳ�\�J��i��M!A���K�3e��3޷���X��6�m�L��ԗh;A^ɫ�r�� =��I���nB��,�J����>oc��yr7[;a޵c���y�ص�ޭɹec�ݣv�^�!��͆oQ�佫�:�-�ȟ���Y��z˵x�~�������@��s5�+���snz�-�kZ��1S�0�ˍh�e�ٙ)Z�,��*��S"�1u�USV�$TF(�[Eb��e�X����"1QkEX��c�f2��P\��#YMZ
��UJ(�Vڶ��X��%j�U�� ��q�J���uJckb���%,V.Z��Ub*E����h*VTQ"1UX��eɎ&
�p�V
)��V.5q*TYX�+m�QFF�1jV4�UEDA�.�,Z�J ԕ�T����1UQEYDKaUT�3T�&������QDEX��M��!�YQ�A���
���������2�%J�eEQV1ATQ`�YPb("�)�U�X�keeTKeUErء��dF**�i���K�̶Ш*�6��E�AU,TMAb���!X.5R1ť�X���2�5�2��q���UXT��eJ:KEV8�R�ڲ�U�lPU*X�1*��%j���+QQ��b�h����} ������>��8*=������_�DCD7:w*�]T���6�x�r�:��	��b|OvVR���x	�����<�a�ӃT�~\	���ok񿮅�xg��l|n6ܒO��VU��FӸ;<e�PPC�E՟/7o���<��q�9��=[>�c���n����Z�	6�Qǩ�ТH##nd�OvVU�h�)�=;���@z2,챿V��B@��o>�`
���Kr]wfz���q��I����
��V!�^)�ꣻi'�%CmCKιؒ �md��taf�R�$�vL�$�m9$���@�GYZ,4a�አc��j��s���Ǔ$@��ʢ	���_�;���5���{q�xtJx��>�Un�'cb��C��,z�0����{��Æ��uP�����GI���꼅�9zF�:>���}�A��rI�#h��ۉ�*��Oݽ�]�gC<⺄x�^9�O�v���I��ʫ���\r���0A.  �2[d��;-�B���ú���+K&9+뿿?��6�nУ�S�$��$�w{���z���'��5�۹Օ@���Ř���s�� �)�`��7N�M7�A$�ueQ ovP�L��;���7Y/@'�u\�p�p[)��P��گO�gvP�F\�ܖ-� o���~�Y��D��vP��تE&�$�6�4g�M��b�el�#	=�[5�@'�w�&�$��TqMt�0Vڎ�'#7�W�,��q�a���m8����v���y�Q�s`�O�wvUE��B;c��ۘ����F�NUC���c蚻���O�&��|wz,�M3�3�<r/����u���]ԃ4��u�	s��7�V;�0;���5a�/z�E��[=�`��Gg�:����c��m���Z�̖Og����`د[c��[�Ќ)���[m��Sc[��;��w㶋˹Ô�����
R� Ƣ�5�9v;m��Ҳ�݀��9냝�x�+��x'Q����PrF�=��b�3��t'C\�qђqw:�q�j�a�v�űPs�o���C�\h�^���=f�v��l�d�:�p]p���c�tv��[�=�:􀊚k��Q�"�q�^�Uooe
��\$��,� ���ͰK�ձDU�ȅ�Dle�񚊴�6b1���` [��o U�\��ˑ0'���A&{`�Yb�~�7��(�FT� ��ήX8���qop�M��H�H�c�3ɤ�e6٪���ھ�{�_\��;��(��u�|A�vNT��1	N��c�;�UW�Q�tU�M
���$����{j�mm��]�����{f�'��[�H${�+*�$���~�/|6' ^ε�o![\[j�A�f�f��{g�c�.��&�6�/�������a�bs��A��Ioee�2 eM����Ut(om��ܢQ�D�p|ۉ�UD�]zc��L��{#�fԊ��.�:�n�ӆ�Eu����M�)��t�m�M�M��|w���I��r��c�g.��WT$�������=ZCƿ���#�	���>�+(P53�w2����"���CP�j!1^ܧ�A&�k&�!�wf��,�|���>�$�ed�&qh� ��5�܃��zm��`��L�l�ԆH"�k*���숤oda���L�ۉ �9��l���l��{#	9��*\&Ň	��$A#3+*�$���S�s�C��V�$Y:v@{1�#te�ۦ�����X��E��� ��=��	�&7
<�}Fg^M	#�{*�o!�2��+)��˺bA&�&�m��a�[@n��1;�4 y��e�a�	'�/*� �oez�&�M8��E͙Tw6=Ѡ�H���9�:'��*���[=�$��Ȏ�?����X׻�����N�ļ�e�]�:����ʟ0�nV�Ww��&p�T�fR��*�X>i�mc���������yTI �o�40E�����Bb���x>�e�lN�@#��&�����l���oغ��@���W�p��,�D?7'��hP'��辆/$S��� �_~�s{�?v �O����6.E�y��=V1��':��7�F�ظ�S1�;SW��ϟ���Ն�9ގ��'3{$P�U������0�]`���ݝ${w��z�]�MJB���:�C �2n�J*�����oeQ>'ֲ�$�!8���d�1�62�E�I�L7POzpQ$9W!�IȮ=(�s����Sk�$n�H�E���� ��Q�D�pCi��UW͙�evv�'��wT(�@'V�ĀI����&!'�t��u�
[��<�>wf�|=^5Z��XySW.�WH��i����d�Z��&��bۘ��q6�����~���	5s�B�E�0a@��Bbh5�>�o�U����d�D���A#]Ă|H�yT)=!�E���F��/"Z!�a��`��C΄R�;d՗�t�"��{V��������Yb��o�U����� �ݒ����l�����k���Ԭ�x(���2�iC��M�j�#�v�e@�3T'�#z&r��8���ݗ�D����{ �>���Iܺ��i�	C�Pѐd�ȐH;�y4	� �N���k_8xÕq>$켚$G^(�i"�i�ኣ]K�<S��ѾA>8o�C��wo*����z`_A`�$�]�	4�l#"�f}����$��ݔ+�����=cK&�m��H��ʢI�{��Xr��� [���)7C��`y2N#?{��Q}�e����j�'f\�6�uz���*����OH{<��q��u8�-���4���P�a$qH��k�9��=�랷nxnݜ��f�
u���l��<v�v��{7���]�o'3�j���gi�$#&2�#�����ܻ��σݙ��7�g�Ol���IvG��y^2�%����ٸѝd�u���0d��u��vS�^[��lpy�Y[��\�q�¡;��n�u�u�ul�cI��u�ݝԛ�K���/j��� �q���f�������5�[�&ӊ���ەamyi炨���G!0�1	��魙� �{��D�A����뙞��+��Q�	$켪&P�2�,��i����g���B�Z/+|��/v�{w��z0����S	�s�P+��sJe�i6٪�;T	'���e
$�Ww��vov����A"��*�I'�{*�n��e�҇��>N��ܥ5�#$��@��F��U��q5=�R���$�˽� �G^��i&�0وb���9w!�![�����|y�٢|O���H�g.�9Z���+,��$J�IKL
 8#�b��V�'���Ϯ��î8{9=��:U	�ۓ5|������6��y�B���(Q �Z˸s.�Z�2���H=��8��0��!�æ�g���� �a���ə@}��B+FW�8
��yj���)�w4l;��i����pQ�}��2"AÀ����i��u臦�4uVE�}��6O� ���*��"�]Ē[��ƪ�\���L�xeYa�	�nG��Nȯx�۸ON��0��ElUoNx�ww��	��$��r9��e�i�l�G\�F���sL��q�S^' �o ?~��՛�V.��@��ޮ_�i�҇���2y�	�o&��j���O)��w�e�M|M���$=���DEf�3x���?�n�H��lIڅ��nӝ�����lt�h���<7a��
&!�j����l�1��c/���.�2 �켪��2��b��v�S��@��n��
4�m3|�j�Aج���`c=ތ d6M��~����&:V�7����b�a��CG�l�d���$:�Ɨ0/~�����'Y?գ�5�އ��Y��r7+���ĆG����og���������(̞�Z?o2JE��<� |���A��$G}��FH�2�,�ۄ�7'����8.�n��|Qw��H��ʢI��1���s*=x�ؐKܑ��~��Nf�G\�P$��ݕBtn�6���D�͉���;{��S7�W�󕙤y!�	�8m�s�%�}s���e�۔r�ػ/�W�{S��ߟއPZ�f"<Y�$x�m��'ĀO�{��>8�Lګ�an��켪�1׊.H�b!�LP[�3��ڌg=X����ث�> �׷�D�OovH��3ոY8�v
6�����ڪ ��۽�D�w�wEL�������MO�Dw}�������,0��>��{�6��R����x�ݤ�����)
�k���~�u:�Q>@���>}}]4�y�𨎪/���{)�Q/+"j4?f�ᚩ�v7���El��s޵�W����7���wxd�-佽�A��g:�/�떜��gǟ�}�����J�C_���ΰ�°�0���GN�f���6Ã
�����u%��e`����9�O������f�0J�߾�͜`u�
ԅ����`t� ��_�~��m��^���O��/�`�.|�c�s�
�R�;���W;U���tlk��ѵ��ز�������uiZw�����^~��:�+(�YA���{��:$�%aF�������*K�^c�4y��N	��~��N��VVJ�G���#�E�v\�T�Q�C2�Q�3Ӳ#�y!�3bz�b�ygi��S�5���$��Z��C�>����R*_�~��m�d�PIP�3k������_�0�a�G�y�j��U���2��:ì*k��wa�:�����}���g
A@����f�����y�N0?`Q�?}��l������߷�)}߂_�ᙚ�SE4�	�����Y��w��~��0d���;���Τ�IXX°���ra��IP�(�}��6u�~�f��||k6y��c'̬��?~�϶N�P,�����c�F�ff�`u�{�6�
B����y���+�ߺ��p8�0*Y�~�� �u�+��p�82T,IP�{�����V	'��$����ɸ�9p]P!�e�
���$�@�1-(�{�Ŧn,���c�J�z=��VM�j�O�No[DD�
2	ܓ�I��i�Վ#d=�B�������"Q͕W&�w�\X�8�nYu�N�7�q�y�������w��)��%Z�|d=��,[g�U��J?w��<=6%e�$oZ�߼����u�Ə�#�Cǖ���ΞU�������:]�5�9�̏y������5v9qD.�;�=G����v��t�*��g���JT�W���l}�e�4��V ��j�g5��0��<^�G���=��dhxMZ��ɭx�i��p��]���L)\���{�{6_����B� ��4{�7�{��Q����L�cY�&�������_�G�����wnb�8��
�N�`\=���S��r�FN|�v����S�LÒ�����>�5@��̟;�ߺ1Fֵ����1g���������T.Xw��~2�����}&w3��^&�o�Jוl��D�p^�efщ9��a{xt�Iy����IS��gxcV�0{�GJj9������Q���ҵ�j�I��;����ݭ��j%a���×/G�x�m�hM�]C �������]�:.-�������������ߛ�8[��cL�$��'��`�ӯ��Ǔ�OL0:����Ə����U_��>&S����|<�x�i��8;ݶm�*=�m|�Փ��3���W���1�\���,��ö��ˇ<羽0?������+��GE�6/������`K2tE����j��Z��X����W��kb�LaikS�\�-�EP[�TU`�1Ac
�Z1�E�a��Ģ��DU����X����D,u�d�\�Ī*�TV
bQ��6�e*�*�����YU����G%�"����V�q�Z���-��+TF*6¨�����#)F#F*�TA��F3Z�f�2�����m��Z��(�!mE��ȶъ����W-P[eD[m�m
"Qhե�T�QE����A[L�`ċb�eEdU��
���ETcQQ2մh[aU��"
*"�*��f�%�
����q*��VĎ[K[R�pc����7�m����q���d�&�PTdUUJ�!�X���ER�Wv�m޵�6��1L�[���j£KJ�wJ��W+&Z*�Sn*���WHb"e(��Yhv���}���F���V�O����u\��؛8z��8�l�c��\ݹm�]���s�6u^��7�Su�{Gk�xyݍ�g��v�n\v�=:�A�ǳ��c�����h��kL��
�����\tw�]th��^�77+��2u����[�d�2�E�7��2w'y������;m��N�y�y!��cn�$_F���⻳kWor5k�����=�)�K��y���GC�<��t]���(���=5��Ytg��9��"{�=$"n�-��L7��1�K��;NR��m�I;�񎶠#��;=��ľ�o������N����ڮ��2�u;f��N�M�=;S���y�5�^fv�q��F|����-�����ċ��)�]��tr�'K'����nlj�������{��ݻ�{c���v�D��C�]����K<P�u�k��pހۺ��vyŋt6���::��q-�,�/nt=q]��m���7e�>�ۣ�սE��u�ٞ+�����˫�+�7jZ9[��.��û]x�Nۃocմ�F�r�nb�_V_� Y���+�l� #�M>ۗ!i�[�76:�Ӳ�n�m��X�mچ�g��͵�Y��F�s����"���3�͛�''Hn�����92��[�����'n�!7N�4�E�;��65����[R���u�]'h��Dc��x��]���瞃��Bm�7;˨v<�9S�^���>�dْ�����ϲ���˭��M���[^���u�㛜82h��u=���$�2����ۄ��m�ݷ^2���Ԣ��ۡ�/��Z�1��6ƞ��x���8�m�s�{b���'6�̅6�{-�	��	�F3� �����6�륋M�۪{s��y�'�*c8\�3v:����<���+��;X�=W\ݱ���s����\S�xH�`Y���˝k��v�'ewfhv#��]��Ohގe'�v��Q�wW���Z�<�Ѻ�j��Mt�u�'�{�yowѹU�.6k��N��Km9{6ݸnq!øs��;G�sہ��aL[���G������J�����o�k����;Џs8�l#��ո�<݊�4�
��.�k.�aZ��Jݶ·lgG��k��V��{F���p�2��ۧm�7��[�cZ�t;�,iܚ:7A����[зf�/`6���)ے9z���B�0
��NRuO3��`NqͶ�3�u�76�)�s��}<]q�ɻ/Wb-�ٕ����w�ݭt����AO|����u%B�VV�����A@�P,��?yì�`{�s��r�u �}��l{H)��3'�M �^��=6l���
�E���WH�/� ��'ݗǳ>�%+�9�js\�vu'P�+
°�����Cl8¤�T~���8�ѕ��VO���G�¾W��%��(�4}�t!(M����<+�`�����ą��������g;HV�
�M~뿯��&��^�o�=O*X VT�}���r2T���6E��5FC)'D1	���`�"g� b�J*�e�p�"2Q���;�ᴂ�P8w�yì�>��I��� w^�k��:�/��7�`T������3Z�f��N$��{ݝN� ���~�`q��r��߹�o��Aa��w�y��T�!RQ=���l�'YY++%��}�=dY }����,�H٨��i��\��nz"��p6���9�۳����=I���1�V�p���8���""�Q�`���q�B������y���*AW��D.�� Y�o%����L~盆�
����~�gu�a}Q�)Yl�E�u�$x>��H�����Ot9Ѡ���qd����D�eN�T�߶��sW:t�8�B��ba1.ٓ�����L���U�c��o{��9��O������g�8�FT
��{��8u�ְ+R������l!�����Z��{jOd��y�	��O�#�����ae�D8T �,�?sݝN�VQ���T�߾�gD�H)����=��W��������x¤=���8�ѕ���VT���d�u ��
!6aD3�G�QG�WN�����y���G�#Ò 9��G�=`T�����y�:�@�P+*~�;s�Ϡ9�F�ܩ��_�W}�Y����dY�X�Ϣ2I8bpX�$ϻ�6u �X����;��6�S���V:������d��7k�Q�������~�́Ă�X~�MO�;��Ob��F�S��A��Og�0�F��.��Xȼ�Ľ��m��l��s���8UMW��!h&Cp�4� ">#�]�"��@�������}��:$�AaF���s���r0�0�ߙ��~�
O�w��ݝd���YY,eO���6N���H�6I�DDC(��GÕ�H�
C�<���������s[��9�HV�+FJ}�y�:�S�a�����@��@���|���4	�ڑgÏ�>
�8R �ه��$�Q�Ds���tC�*���<��8�%eG� �Ⱦ����~[�;/*#e@Z�[����`^�%�������˝������lT��K ��:	��z;V
����f�jp���$��?�XH)
Z}���l��l�+A��wp���"%�/�&�0ˈ�p�DYet�"�4���i�|��Շ7> 2<	�y��6�
��w��F<��;�͑Gޛo�8ym՜��3�I�#�����G�� ���8�	��fE`r5����Ï��-�=���#���؊t�}A<Q�;���x*6�@�t*Ae���6�FJ��  @�6E��O���=����)�*9ݺ��ú���,���ט��6���s�Bkr�sQP�A6�U�F�)'Cxq���$ן��èu%��e`��;�m��D �D�nl�>�>t*W��F��Hv�����8�R�/�w���B���!`&Cp�4� �����r:��ed�O;������H���l�IԂ°�-�����*K��#�6E�zϑ��>Gި�&�u�?;�Du}�#��,�5�\��i6H��bGk��͇ � �)h����9�B�`V�*gߛ���sZ��{�O�K"eK���r2T(��A���G�>Q�E [MC�M�^a��O��}�}��;t=����?$���������6�FT
%@��y��`u� ��}��s��oy�9����ƽ��M�F&@�P��~&E�?r>S�f]��H{�}���O���a��!�R���+�Yq�/I��{���R���nH)�{���Z+�u�3V��Rk��=���e+,dDo��dX#�@���:Iߖ��� �&���y0�0�*%O?{�͝d���YY+*}��y�tN�{��������~~}~��3���/F��8�i��ti��
��і˩TY��[H������D�t�V�`�Ϲ��� �)hy��6s��k�`T�߾�`q: T]�W<8ؗ�{��pd�X��H�fȲ<	��]!���!���T�~���u%���}�y�7�9��?}��8�2VT���|���0:Ԃ����~�́���+�ܾ�=�����]��'A����!`&Cp�4�
�I�>��:�Y��YA���{����F�w�����[�m��������c
��RX����6u����2���ȏ���G�� �B[��""!�|�|\��z;pO7ݒs�+�#�KH[@�|�ݜ�!Z0+X)�~��E�!>D,ܩ�峷��1��M��w\�8ì+
s>ߵ�֮�k2�F���§�o���u%B�VV�����'��������w���bT
o�}�`u�
5!B��=���읤HV�?sp���S�~�}�|�ZK���|�Lޏ�Fj={�Ql��9��3w���]��}6{m���L�ٶ���<�ǧ�����?���������ǭ`�E�����.WW�˩,���l���q�1�鹎:�d����^6�л<��R���3q�B�E���v�4._��#à���yaf:��w�b�[k�n\v-�v�pS���G��E�=K۱ہ��\��ɽE�G=�e��9;�;$mf�U��c�!vxѫ�^��y��gl�L&�1��8�Z�<�Z����h̽Iͨ��.E�shW��^��t�#�>;f�F'e��\Yz��������%q���j��<O�&���vu:�R+%O<��6�J°��~��aRy�>����_�ĚL���βu� �VR7��dD�jQP��	fB#��=� p��I�s�S�G�p���g;HV�
�S�~�́��J�%����H(pIPw��\�y��6�zWnH��g��\c	(�f�c����5߾���N�Y(1ۗ>}�>D �D z8)����y_w�0?`XԂ�{��l��m!J��>h�B�礕��ۈ[�@�}]�"�חg��>�}�|�J��9ݝ�:���aXR����a�%�('�y�͝d����~�����G�>�"3&�G�d��Ж��֔��ѳ����w�Ï�
>��G�;����Ei��Ϗ�DT�t��AN�V�;��l��P�IP>�sdQ�|��ڑ�70�`��k�niz��e��.û:!{<��+iRꔨ�WgȠ�MBp[�$�||�:C��J2�|�����d��B �ۛB��'�|����(��x$�s�߶N���`��;�m���w�?.��5CJ�E��?��E�`���G�In�u
�*�"_jO�@�E�O�#�R��{j��җ�,zg���s�?����M~�[�rζc�4�ˌR���f~���{�E�w�?$�%H,}�w��B�}���6q��ed���׿W��Y�{�}��'S���~��f�����s4�F�y���r<HR��>���l�JB��Z����|��=v�w���@����ᴂ�T*}��6u ���WB��I61���g���n@��ν߿o����Ad�V��83����@����l��H)
Z{��y�;{~Xc�=�pƠp�4��>�6|$�>�= ����� AG���GS�����J�y��l蓨n���}yM���'c
���!��*K�~���8�ѕ���VT��~�d�E��m�a��u�~��P�~��QA�tz��t�p����M6P�Ŧ�J�t��エ���~��E֔��i��������aǉ
ZB��}���$�
сR����p�`�'n�j;�S�\ ��,����l�%B��Q߼��ΰ�°^���nC��u�'�D|��tB�sZ�<��ks��|��g+*�P/���8u�ְ(ԅ->��� Q���:�Լ���Deτ��"sؾ	C(�5CJ�@�>��x�2VVJ�}��l�N�by�O���_��$�؇N\��I�n��/1��u�e�4�Է�V�IM)�ý�V�שM�%��<%vny��Q14���t�ժ�1����.s��?0���{��$N��Q���w�#��,���)6�-A�f�`pß��߿~�ɼN�
ZB��oyݜ�!Z��/�����H,�?o��g{ߒ��k?k�]?I��Ͽ}�ΰ�°����_����F��:9��¦����;�K��^>Gçm��}蝞��1�7~� �J�y�}��:5�Z�����́Ӵ�e!Z����C�;��ߟz_r���������c\t<sz��������r��v�rlBig6��__�9�y����O�w�{ݝN�VPd���>�߼�C�+
0�,��;�q�T�����y��]�<$�?~�l�'YY(��`ʌ��G�d ���kL&�١g����jHp��I�?}�z�ןl������!ă;���aח��J�Qu�,�h>� +��&�ff���6À§����:!Ԃ�YXy�{��8�YP(�\�����y�}N~�5��Ӊ������{��������;�q�`T�����4�3V
���(�#랑Dg�W��uSV ���T�>�͝�:�IR>���8�RpB����w͝d�uϧ�v����횋�����q�3�J��	��6��I��zf���3ٛ�wMUs�f��u�Xd��ߝ�g"΍9'!�0�����i�ߏ�W�#�E����m�Z)�!�� �w���?ąHR�?���l�C������G|�D!�� -;*P@��K��wp�AC�%@@���{"��'�k���L��r�䑿�t!�X���/`aS����ηlp]E�,;Wf�7B0�m��܅���m��xQ��
����a�C������vpg(ʁR�S߼�:�X	�m�g�}��%�u��vC��JB�!}���I�|!�H+(Ciǡ� ��{�vu:���8�����M�������X���+�����0�,B��{���gY:2�VVN�����F{H����,�>v���	�DfkN�0:���ą��-��{"�!���"<	�lW/�`��+,K���p�8�P�*C���|,�#��c��ۈ�h�xI�|}7���E�
/�{�|�z�*A`�>�g�d��J�O?{�8u �;����~�́������������!X<�nH)�o߯����4�sV��bM{����t@�����T�Ͼ�gRuy�&�{���i�aXYy�<�6Ã
��RT��{�βted�����>���;��|�����~����^���]1��L
�6��`Twwi��A�zc��2$���V���<�FL�hw'��z|X/�P��0^��(��,�~N28^���\tN��t�΅�s٭(��y� d��s�;Q��mѥ�v4�떥H��]f��	��^�>ۓy�ҚA��T2�m\K��oa����`+�N�͔����ێ.(;n�d��u��}Y���K��e+;U�q�k�����'6�\���ݱ$�nu7���GO:��{���$����g6�[J���$��dmgs����P��oH�e�
��~��ݣ�˚�����ﹰ�x����{�6s��l`V�*_���8R
�e�������k'�O�yD}��#��g+�)�j �^G�"+�@G�>������v�Yn/Ɍ��6x3��P=��|��Z��H)��}���A�+��yw� �O��>�># T�4�I�=�:�++%e��>�߼��=dG��@�#�x��O9��n��o�m��¤�T���w͝d�S��y";��dDz�}5�d��lг�,��y���G	9չ$x<(-���͜�HV�+FO|��6
AgD���w���_`��8�(u%B�k��ΰ�
����}0�ֳ.iu�\��r0�����:��VJ2�|���g5����w���M m*7�<��X�`Q�i������i���|�᷃�����[�s�����˹�7l�<��E�WM�o\k�[�����ѱe�������`�g;���^~��:�@��2T��~�gbN�D� �����6Ñ�I����ׁԝNo�?l�'YR%S��̀� ���i�L�1
��������(�$<7��٘w�1_r�]�7t��Q������;V�~}/���homٓz�TУ#�e��Z��52�!���n�S@F���_��� C����R�
���a��������@��w��g*AC3W�����e���N������>��X��H��QG!�aS]���:!ԔB�Q���ۑ@����>Dx }�7;SA����䂐R�}��l��m!Z!w��H(��'s)n:�5L�l }=�"�����8 '�}�|����w'D�B�+
°���{�m�%�(�}�|��M��?f;�H,�eG�}�=~"�v���	�DD6hY�:���ą-!K@����g;H��f�Kk��H�$}wu 
#@ *e�w��g*%B���{"υ�|3#�ϫK�5Uv+��2�J򖬏]��E��͸Gn�[�� �竳�]�d8Dv�n!C���g�������݁ĝB�Q���}��3��� ��>�odQ���f��_f�����`t� Ґ�B����6�wZ~��PҠ�}s�(�� #�}�}zb���`����"�n�p$�IR~���6Ì*J�ID��;�βted�������|�y�s��)��#�E�OF	�Sf!C4��~������-���͜H&���|"��}����?]C��u���e�rhݵ�eΝx:�{@~���;cZ�vA�p���/i?4O�afg9bQ|[ߒ9�G�#�R�<�q�Y��<�h�����r�������}��T�����%b�O��&��&u>��Mw�G�+����9��ךL�;b^t=&V�/f�sp��Ϩ~kݰ��8�mg��C=��/�{���[ �0)�g���	i>��i��B������{|��vs�1`-�0����\|���c6��ζ��@����s��*�a�C��{P��U�2zT�fE���2� R�V�+bn��<=����V�<D�����[�mR���\5�s��#^,���G=�4��3�����?Wȕ��)���2N�����2��Z��}k�y���MΞ���l:��;��{v.�<���|,ǃ� өzA�y�Z*����`�Du1��|�K�����
n��k-kp���:F����z���n_l�B���򎂸]g�Վf��=v�xEן�����e��뮢�gF��^��{qv���*3��7�7,/{'�x����/�	�ݤ�e�����x�n�|r��������O��%���ˢV�U����at&�@J�* �[�*�I����-Օg�����P�w�k�?I�.��;�)��Wx�	�<ךV��9q��a�zu�-��Z� �Α�W�&��J�ab;�l6ۥ�6	��ޜp9�rB�u)���ߖ�̝�s׷&�spb�Yl0��Q����}7�́���۷�F�l-*�^��;�ܧ{�5�ẙ�ME��a�U��Q�E�(���*�GƋ������Ń[Y�b�6"
�J�E]R\�T�R��\AQF�Ʌ��St�WY�m4�2��B�����MEŵ`���f#��V9H�zU��V%e7iĺs�YX��X�#���1cmt�mm��
��QQ�`�����`��*�Z��E���E�Q��Ȫ��-T�
���r�,QՕ4R��Kh�WIW
�eS3f�(�Wy,GM�XċUQQ�*Ķ��#�\���Q�\p��QQ�ҫL˂�cv�X�**�F��Ur�L�j�e�D[���b*;��ADImUU-��A+]�1�1.bd���U�UR�bkEQ����i�Պ�Yf2��,�c1�b�DB�M���PVh�
AE4ֵM�Q������nO�>��/������D�
}���gR������@M�
 �^|,�"����jgs�t��ԘVJ���~�g�J�%@����:��X5!Rw�l�;�c����dPq)�G�4@����6�S�����\na�3Xf��i8��}�vu: VVJ�S��͝u�wI�����7�I���>|4
��T�'�}�6u��eH,��=��G��Y nvv�2H�$�FKeCj �>�B����h�;<��ͶO=ԝ�М��fe�3}}�>�<u�օ��i��A`��y��x�����~�����)
���=���G�!�:�����s�I/�	>��P�%B�{���gXv0�-����k2�Z5�i�>�}�a���
����5�ۯ�k�瓬����q��*J�}�|��cX5!m>���� �HW:a����|\�翷��"M�5PJT �,�{����v VVJ�2T�Ͼ�`q��#����ϧ08w�}^�S�xI��H(��|��N��VVJʞ���l z]xr���5�9�eH,���;�[������{�� �;-�s��9�B��*_�����:�YR���6͍�5`�bL[���P�E�na��0���C�8L��Х��=N粴# �gh�������xvɿ���`�/�M��˝w̹��}�<	 WeԎ0�aX_?y{�����Zr�:9��¦����u��VJ����wgq�p�����$��@��H��,�AH)��}����A�![���w�>����=���|04SP0�1qIX��k�����c��lc�ܽ��{;���I������s��5���$���ݝN��2T�����l�I�($�+
��^�x3�@�"=����>Yt&\�G\�F���L��?y�βu���������~� Q Xە򅩰[�Cf���O�(��4#���inR/2~T t�l粐������u: T����;�i�*$�~缻u�,D{c����"φ|�>��m����ra��O��}�u�����{��6�YP*T�|�>��|ϝp�gޟ0?F�+R-?}��l��RD?g|�ᧃ���>�sZ-�Z�T �,�?��E��d�s'�'�}��2T�sݝ�:�V0�)�wۯ|+���H���}�G2�v���VO̬�eO�w��:~�~�����4����w���!m!m���ȫC�����1�J>����@N�T��O��{�i�*%A>�odY�|1��s�<������[���;��~�k��m��xϝb���/>��w4M�.W�������Ϲ��Bd������mm��rl�s�E8j�\�qvU:m���i��0q�v�v]ێva
�t\Mq[t���V6�%��붕�	��������)�طjwO=��:�
��N�s[����۵Q弒�q�
�c��m�)\sݞv�g��{.�`SY.���ڒݑ:�n�x����n-9w�W�|�\��x���=aC�9�� ���N�]�j�����s�;v*�O�[�^����]ۜ�����|Ն!�uں9�BpaD>�����"��vC�(!Ro|��3l�e@����y�8u�ְ7�ۿ[�=�~�>���x��5�w݁��A���边�dx+��$�B�D8��$���ݝH,��Y����[�y߹��&%־�`q ���a����a��Ib%O��l�Ad��ɝ����ru7��r=�� �+��`�$�6�>�kn��Î���-���͜�HT�%�oo~�߅�A"F5�p���+*y�󻆙���RT(���{"υ����
�A�6��0\P�*}��������3�^�I�B�Pea��|��m��*A@�߽�:�,��E���}� }�o,�M��J���dx5�ߙP�JiCW`q<k���gS�ed���<���ԝC�;�o�3G~�J��°�y���i�T�!RX�~��l�'YY(|���|����dz�@;�S�����ÿ�c������3�dh"��(�]>xݮQ)�c.My뭤K��~��񭝆S�|�w���oa󴅖�P<��|���B��Z0*_���8R
}��}u���=g��;�ۆ��d�Q%B���w͝a�°������Z�ֱ�̺9��
���wa����>���w��/)��"�µA��S[F�eZ������}qo�²?j`=�0>��sK�|`�A���N�;φX��1�n��6|ͤ
%@����8u ���{�߶�i�B�����{��[�n��dσ4|!yf�TB�D8��u�������J�S��͝I�,IXPaX8�~�~�7��}���}0�0�(�IS�>�:��T�ȁ�#��@@�v�P�!��u�Ѭu�6����v���>����JB��Z0*S���Ԃ�@�����O����ٗ*��_N+�{H����϶q���aK�~ϫ�ֵ�f�Xk��F=�}�a؇RQ
�c+����l�o�o���|?�M�|	P/�￸u �:5!e��{���i��E^��I� ��������#\ݘӞk�Z�6ޒA��ɦ���ca.�����(q5ھq؄�i6�� 띑D}+(�YFJ�y��l�N�RVaXP���y��¤�{�����}&�y�{�βu� �Xʞy��l�N�{]�v�\[�̦i�X�`����@�K��cO>U]2�*F�A����M�S�|j�t�^��{3"���z�*�EP�DD&*�b��k�����A&�qr��9����~���1��Έ��������E������}��&�[����e��T�s�r3{$�&�(d��Z�-9�<	#7�*�$��$ېJ�Q�����Tane��v��8F�]H�I��rH'��YS��(��k�)���0�1�T�$�}��@��sKO��w*���m1$��9�@�6�S+*�m�~]�����n�![u���_n]vvx6��%q#�Tt�a��@�5�"	m��`�;�����2��A'�s*�X����H}WL�x�L�$�e1O%kp��Sh�謝�}���hiy{�I#���$�NeW���`����;_��m��/��@n���dψ�ٙ ��;�D�|o��f�b�tF�í�$���>$�Nd�$u�W�0���P�����ʘ�1ۃ�F͆Y�$��	ޝʯI�*����27�t��ܽ�1���Xww�+&�
�>@��kX��h�WaJ�}w����EҖ�;���Dbq�L����J��w�(��� �o�O� �,(pDN;�$v�Э�vF�Ђ�|]9rH=ӹ4��\�w�_������ׅ!x����ԓ�8QI���]����d��V�������?"ٶ�Q��S������ �N�WP�5��^�F"ke��$��Od�$�\p��!��8����;�ej�|4zU�0�/gr��|wz��{E�VR�"����.m��i�f��hQ'3��
>$�����O4ޒ	��ʠI ��t��c"ɀTC�!�&M�ٞ��}�+�o�H)��H'ٝ]TI Z���TVɂ:���
��=k�e&l �:��++��W��ɗ���2�َ��H=�]"��Y1'x:#�*�3E�ʹ�-��-��wL��٦��9���:�0�cr �훣�����V8��{�Ks�<�����c!��t�$j����xn/dz��F�ی�\1��v���p�D�d�zsK�F���lsy���.ƺ��ع�96�ݚ�<��\^���<���=m�sk������A������v�:�[�E���5�X�cY�.��a�Jղ��������a����l�.8x�j�Cx*E�&L�dt�c r�8��[s�hI:�l�#�۶t`�\su�K��n/6Ʒ�V{u�Z�v|&��$����������GSݪ�I=�]T���Ɂ��in�<tH7=U�A&�z�
>�ep�h1��UGLVHd���l�}�S@�I>�I�*'���=y��C����1������A�u�@����2H9Y�n�Ϋ�{f�gA$��o]
��ʁ59K�m���m��[B`J�\�a�Jy\�Is}TAU��7�2uoeA�1��4OD�|b�r�DE��0
�O�ɓ&�bA �ܚ�i�r�$_����� >�QZIF?������m�������;c%�,�^��1�q�[���<�i�&ձUf�����1�\(�O�1]�B�Ʋ�|O���M�OS���qܛ7��=U���ډ$x�X�DAB0�q<�j�^�텝4����WX��ƨrǨj՝1hq��n�17i�Y�����ު:M�2�b�W��@ݾ����~�a�ƕ����٢8e��P���X���\��@8kj$�t�Mx��݊���]�
�e`�h1������$�ܚ ���N����YQ$wNd�$�\h��!��8����}R7{�X,��$39&�w&����_Nc��ȝb� b�Ȑoj�DF���n�s���$fw]P�{������"|I��ɢ|Gouש��&���L֚�&J6-�M��vB3�A#ۆ�\sM��M!��'��5��ߟ;��_�'����'nw&�$�{{�kǽ��.���m*�>'���I�4�L@I&'v���[�yW7<���~'���TH$��]P ��U9F֝��#:��"
��ˈ���UA��B� ��^$S�Z8�Ú�~��:�{e#-�z?:���~!NŅz��U��(Oa(d�8�Nk���mo_����͘���VNG��Mx�A��zcA�`��T������7е�� ��d׉'���]Q$��]Dܝ��w.O]_M|g�pBnC�p;�s �	8v�C����B+���s�U�A ��]P>&�]D��xF��m8���s�ԡ;���u���n�zL�7b�e�q�ź����=A)�����Cm�J�lEw�WU��s�$s.��5C�R/62�vdO�fu���(	(��ɐD�L�5]�
{31FxX����$H��TH$�]1>;-�wu��2������Gbрa��(LU�T(�A�R$��F{Ǫ�C��Y��H7�N|E��D!�	��{2�wt���$��ڢ	'�v���ٓCw-;K��k&�`��G:����sxc�ڽ/�8=����ɭ�f�ڴ��z��~*�ީ�&�=clS���w�&�7��r��1�!�6�Pu��$_n1��=������	�]]u@O���;ٓ'�NHt�z����~_Ÿ����Ӯ�v�J�e͌�m�}�6��7k°Z��������ꜷg��[T#6��#�1�J�C����nU	;�N@&�ilCP�M��b(�������̗�t(�A �]9���$��[��޾����v�D��4�$���d�ܙI'�q�$�bȒh��'�]NH��s�A wfH�:��F��p�1AOt�j=����Ok\A ��.|A�ܙ�A��D�)��ƒ�|���bD��a2�"F>��I=��^��ݙ��)m�9�}Y�3�A's��S ZeH�;��f�Y��͡��v{��ɚ�0k���ο=���%�~�e��9G�u[��]�o�O�Y���ߕ��m�M}�����w\�3��<�N�|JԖ�9�9�o˕`�8R2�à���r����i��a��q�����>����Hˍ��.�K�ķ�g����&u�xI�_,LcE���ȯ��OMtp�,�Tsۀ�t��T/M��)�{�����Nۮ�;b��A�w\�C�\J44'<�.7MTH�nf�U�*�,��{|~�z�T�3���TŃ{� �	��ڱQ�~9R��2����s�Y�Ͻ�9�2F'y�q��N�q�F�X��t�z�97L�qf��fA� ��z�et�1nzc���8���������2;��n��[�P���o^�ʣ�zy�l�w|�YT^���;	���4uvF�4r�z�i����Y�r��=g���䮁VMH����i�R�����1��Jq���ǎ�7����� )��5 {8*��qM��F��>ZJ��a���<k�ܧ"�z�s`��߆y�n�o���w�~:r��@'�5�ܱ�)��ܦ���ч�Ǉ��Ө.~j��ny���پԲ�a���9t���9����x���d����m�s�Ҿw;+���9��a�������+{���j��m���=�!�Vͯ���[���n�;����p�M�̽g�P�9[�Hj�*Ƚ�df�f�T`j�I@���j��J��V�(Z�1��X)Z���EQek*9pf9k��*%h�������,�����EDF�A���QF&Yr�LfSɘ6��c���2�W
8˕h�UkehUe���l��lƩr∹h�lıdKi������n�ATb�q��P��3˘QƂ)��:AF�n�悊e3)��J"V�l�ůs�;��B��Ѽ=���ݱ���V:B�;rn�r�q��8�����������̠U��L�q��	�������"Q���7i��ڭ����b�����Gy3�̦cl���3+*:�Z���`.P��kH�ңV���P�ݸ��\�J�[E���ۙ+�(#b�B�X6�\f�L�T�.��W-feŋ���nZ�p�aDV,UV�z����f�a-��9��\w]�U�]�[����:�sgtu����vzՎ�-p�^��s��꽨n�+��HDy��g��m���>��{6�)�N�]ls���K�͚�ˮK&۝�8�g�.�����/�"ݱ�ۖ�i7[p�5���[�PY�:�'��Wg3^�l�v�9PS˓��۠2�u��v�=v���z�{mֱFN�Ơ�:�r��BΟl�*�n�gn:�e֛s[B�g�oB�gjn;{a�f�[��ln�N��l���эv�eznn�H�]�W\v�(��8�
���c�R%��͋��;v��s�pj�RݣA���(v�JŎm��=���ہ��\���R��W&��n}�M67�V�ۇv�B�r\���}t�v^��1�%6瀳�m�۸;�]��y;<r��.ݍ�1����Ν��>w����sf1�RM������Ҽ�`ƶ��m�Xax�3v˞I��z����[�����d�z<՞�F�f�x�]�B��B�Sqdx�lULi�y�ܦ�[�;��:㙣!;m�Yq�WV����(
�o3F�p��!�pA�u�<;��r����\��l;sq�g]<��;<���3W�]������D-�n��nX�nm�������,��>�	��z���5���9�{g[��r�)�nv��c�luI�'�V�&�}��p3��{!�ϋv`��*�f�N��rrW=��j�%�0q�D���lu�;V�Qθ�e�����d�f�V!V��(\�0/M䓨عxX�7�f��1�T�U�ӳ�.u���͹]q��
��.��lڎαǫe[���o;C���{kWcZ�=A�}�k�8N#�m�&���vz��5�.r����\�'�v�O���q���خ-����<g�<���&M݃8�6n=6��[AuWm�u�]�&���YkٗX��a8jc��%�5�Z���6�{�r�ic>N����9��g�"���#<ݦ��ڠ,ݪ��u��'�Os�ɭ�gviP+�^0�s6���pa��lU�\�ꗣ��:�{F����x�(�v&���(��:�tiݩv:��W��瞯�s8��s���}}Wѩ5�7;���Mӫ�5`�S�g��Sʜ��mm9J�끜Ul�#c��ͬq���0�N5�䒒s��y8���ܘ�n�ݣ�6���:�g�;:�V�n�v*D�ĥ�:N�μ!����B�B5�;K� �n��b!CmO����A>7یO��v�P�.T��"Me�[=�	 ��ɟ��Ҁۃ�L����+�|Cp���Rjnom�1�	 �o7&O�;n��6Th-�0ޓw4� �!8h&؊���$�s;��Dc.��v��A���Ăk�$O�;��@Q0ʦ`�	%œ ��C��{���` �_�� OѮ�� 3�����S[�.�����Bb���Q�7.�zneʁ�O����ْ	����/����r�Ff쮄T/�q �F{4NnZ����Lv�F�Gbx��l�k ��q��8D(P&.";^̉#;6�Q$�o����eov�2[Z�U�� ���u��g��4�P�S@��D��W�k���@�T3��W֑:=��{�v�1{?[��_{�G��Ȏ��'�+ou�v��Dp2[��rRcv�5H���#�I��T	$�$�ګTtN��������4��0S.$���
 �λr	,h�U���E�ٯO��޺�|H7�nA5�K�'�G�^�v�d����J��> ��vĂ}ݙ5;��[��%~��ʚ=��3@I&�,���,H={�N�4:�͝�K�S]�D�F�ے�d�n�Y���[4��Bb	8,�!Z��p�1v(��{�vGU|�q����@���	���UDF��N�dό{oq6�b��;2�Q&���$�X��C-L���{2$�b����{�$��˷>�3��{� ��~mkV�����1��0B�ڪ�og�|O���A�%��N=��>�aR3j��LӋ��;7ˮެ���#P���:4�*7���]z�G����h��<�aMt�5N�L&XP�r�]�A'����2gė���P\O��λ���o�6�d�	�ܐ;3����J͔��ė.|O�d�NU)m����we�k]��R�+ô�W��*�����3�I7��B��B��?߷� l&�����C���Y���*�ũ��l�#7"�ջH�Ͽ���g	�V��Nt�� ��9 �|O��n�c���4p)7w�H��s�@��v�Pl�cy�_�Ͱ�ǜ�l���E@������u@�徵�xۍ��tI��!B��a2�##[�A��^�O�#f���t�	{� �H;��B��k�F75`é"��U`ܐ��&tˀ	�� �A;��B�O�����]�1��XE�,��jc!�&#79eBsN�믌2�͙M8�4����V#��Q��c�␍'o�i�����֤������rq\�p���v��Q��u>��*�9�Y�D�G_\�$|k�n�A��c���\��⦱iE�p[����^&O ��ɲ��4�k�9e���P���}�n�����ï�Ngu���s��o3�4[=j��d	�:�Q0ʦ`�E�� ��J69ýJ��wut�	&�z�$��$K�:��%Ҕ���V#�Z�a�D&&�V�H�/ $9��W�f�Lpuo���͹	 �]1 �X��B�Z0�qѭ�V�Ran�`�y=t(eӐAٓ�/�칺�D���T*����!CmM:�H��M��h���{/eI#bz�P$۔�7�&A�G�\u��w5жh�.ɥ��B�����k}��������sL�=3����:59����W��姅\��&�v��ǹHVq���	�j���ε�g�8r��:�]e�nn�����;v�c�����K�<�/W`9��&νtdv����8�zr=����qӝ5l!��t7VvlO\���Ɲ��9��������9�7A�k�a����:���U/e'���p��ۉMu�v*Gr�zPK�Y��n1�`�qgv���K��x;.�6�U�+���-v�k^��N��VMl�1�-�n�IMo�Оp�0i푶� cp���$�V�&�@���ȗ�1��>5n���FvT�$���ɟ.S��TJ�/�*���e9��49�M�a��W�N̒�Ξxm�L��e9'��fL�|F���^h5��n�dn�T"�l���'vfH"�q�A���@���>�sR,NvS�I=ٓ �b;d�
a�Bbh}�N9����H٩�I��rd�A��rn�-��	v�|s�J0aC-L����	 �f�U��}a�Ud���NA y�2O�����d�Dv�B��y�dD4�@�6IEq�1�"�^��`���6�jݬ3�{�������(m��6޹�'sq� 	���0Q����&0~�́��7B8����E���$㻏�`t���Ȧ�l��[w���m�".'�>���j��k�o�5��n�Q�r��w��?RW�2��HS��.���	��ɒ;��>N4Y{˷]��#Ph��fptN̂|I�H���K��V���A�_d� ���u�'p�QM�dL��}7tRo�܌d�2�܂	�A��ꍄ�]H�
�HU�"F�ዃ�e�	��b�������fj� �$wM̂@$�v�^"�]D���g�����I�����$s6���h��ݸ�v觝�veU��9�&f�����疀i�"�fI�$�ۚ�k��J��pNՊ���I��ͺD�z!jd�	"�`����پ~��	��ro�ko|H$���� �o���C.K�DMdLUg���H��D&@q'u�PA>#:�d��fzM-���Kf��ɤc�3
���[�<�����LaM����{+�������Y,h1��
j���V�{�ͬ��^�ޫڳ�#�3ׁ�R��S&nNe���$��۪o���2�֔�.a�tN��۶�n9]�{@�0���$�˦$ݛ�	�Kz�Z�VVېB����TP��)&�,�!�L�$������.��X�ݝ�(��t�Ovn���:r����QD�w#��q��x�<%�9s��Ӄ�<�b�m���6���όr0�8�LHS�?
�u2|O��n�<�n:��ʴ�����T�@���{.IF��&�Q�ff�$�u�yX3�-T�[�=�	̺rI;ٻB���f���v�M���=��B�`��T�x�}��@�	,+��a>ܼ����$�ݪ�0��1ă��$6��kf;f��T�$uWH�I��ڢI�v�&&8L`��N�.�g�S�"^79YZ%�Njק5˼L/=�?�{/�A�]�������fΧ���v�!��P�霪4�8=��L�w��e����aA�	��6P[=�D�=t)�Rݙ5qB�L�g���I>�f��=��;yA��b\\�*�C�C�����B}�(�s�P�2b�=$�mi䖌�|�����# ���>ɟ	���$Gl�����F�O8�\��Of����8�e���g1��|�; Si5"y�Y�=��U�A'�v� ���	�OD�U�Y/I;�$�6�M��1�UB�흺	�ݙ��d��֫m�$��;j�>'Ƕv����!C��<�y�Ϋf��Oo)$��t�$�Fl��xI��ldw[�ڍ�b"���!Sv�-��K�-�'[��4��_�"���?vP$��Q��rl�+�g]�;�ȅE�Zp���ÞΜ�}���"M�2"�Ʋf1ɾ���d��;˺U����*�h���(�5Q�]��7��w5Vǵ�p��q���ns4ن��#m�>mnnWuhX�d�݃�ś���h;�q\�98�Ǯ �nާ�gc'Eۿў���e�������󶭰.6�w�]i.�o@�n�.Zї�t��Os�5�n;n��\���M��+$��K��'���e���{s�����q���&���х�.�ڍgp�jՓ��s��ƻ�m�	�i���qz�q��Z�j�'<�A3w�w �����{��$�{�T| �>4aT]��7ә��<�����P�&�I�&|C�2兴�)-��a��v���I_u� A7�O�#�Lڕ[�	��PpC�l0�!1Tc/��GĂ7j�I�!���dM�k�w�Y>:����'�r�`&�Bi����Q�s���㄃�U�(H;�NI=ٻ;rl�	���SI��z�WD�����/�n_�`����d���{�� �wu6 
7�����RH�TY�joѮ�j8�Q��5�uۮҩ��&S�v-۬#j�,��`�ˀ�7ջ##"-H��( =�m2 @-���OT�ΗQrTD�M$d��� �nc��oDT�&*UKϻ3 :���.iӾ��<R���F���Iۉg�<:��u���u�����jN�rQQ	-+��6�g�{�a�j��ѡ::���b {2��ݎ""/�I���7��2.�]��,�h�� �h��3'Ivwu]�I��m��l��S��of;` ����F���)���J�d��~�}�v���� �wp���{��o�e�nӍF�$�Is�5�vQ(�ND4ڈ��-��� s�җ.��>'36�P
7���7���`�n�vwS����:!�GU��=����8�3�^#���=�Nyٝf������s�0�	�q1�eζ�|���� f�%�5;��c�N��wm  ����Ł.�732U)�+7t'�	�N��K������Y�U�L��ݙ� >��l���r���ԏ�A8"5�q%l�=�` [��E��ϵGV�c&hB�\G�g�k��.��Q}�� ���8�c�g�#�z�on�2�K.���[W�KM��y؃#����M#��3���us�C�0e� �.u��e���GT���� �z��6�];��yJM�m}�ؓō�x1�,'ua��[��}	��n�xma��ݷ������V�h��/b��yԽ0��?[���I�ݬo�>�3�V��ȻhW�����{|KTE:�]ӡ2�զ��K�P�>�ܭn���{^o��[�����W	'G��A���������z ;�/j�3-�O&<Esp�	n{M�x�׏���>g{<�GK�m��l=�cE2m��>�����bͨ�@{(�!�ý��Ô���yӷh�ү��`�o�+"���ܜ�/0�[w
<�om&Ȟ�*�u6f>�Y���>=��U�Nq=�C�o�`��o;����^��٭t~ޔ/���z��f����~��7�����)�����ri�5}�|�=�4�UyW��Ό���9޻w�;�z�,%���8�����מ[�����w�<�[��s�yJ#=�p�|��d]I)�@�!;֠��)��ww�CΜ=<���r_u��y��g���ʂ��ٗ��S�wt-�@W�<�����ۚ�Yr;������>7����]���ج�r�Nc��7�_+�����6*Oh��Y����5ZT21q]��@p��Y��G�����ET<+�liR�9y�I���y&0�I) |	$�
E�\F �3���J��(������DUV���Z*X�iRm%Yf��uK��#�6)P��;��t��6�}����E*�iF�	��ĶՌT\��QEW�3%�E���e��h�-)R�-��f5�b(�mm�QL�V�����4mZ�.L����Lj�-EQ�e��n��gu��4<�:
�m�;g�iz�5a�n��aM�+n�m̬�R�ۃ)Yk-�m�҂5*f�jT[�k0Rڛ�5t�Le�uE�7Yq�j4��H�lB�ILQ�U�E��Eԭ�f"�h��0X��ՊYZ���W-Z�q�Q��FQ�t�ڱp�*aQhʳ(��#l�fv��7-u�@wq�xܜ���\�+j5��5���շ���� @ �ܦ��=�=�DU
(�!�L�2"zN�v��T�L��s:� [�N"!e��َf���n �ݻ�H-�Pq�a����	��̐3�ӛ>��߫��b���Y'ğ�
��2 X�.���l�_Q�1�����9F��Z�Q��\v�2��MmN.Hٞ�A�����>v���W�߷�����	_nU��F>�l)�sӽ�7������{�M0比�Z����yUH�����M��U�~�����6���>��=0�\t���L�T�biD�N_���q�e�+6���fT�T�wDj +{)�D@�c��d7�$���8�
:���	���6)L�� �6�l@ #㶀� wovF#�~��@����F��<=M�2���}i鑝����i�7���Ql����(���=�SPm�Pɻ���;�c���y�{� ��rip�0�ɢR~b	�t̜I%���F2��0q�i �k)� -}�l"oovff���n}����쫯;q��K'O�{;9�\7�1��R�6{)��/8φ�6�/�����-5k�K����[!kܶ����$���Rۥ���!��� F��o�v��	�����jfX��ٙ�` �����mYt�:��n F=�l�Gv�fa t�ޙ�j��W��2g\Ӝ�F�UMK�.��l>�����R��}rk6cӲI÷�RM��{����廧P�	�S�H�����S��7�^��@���L>@$����@ >���{�"1�Q��v��?J
�jh��U-���ݎ3�6�*弿,Z���Y��o���nb��ONۡK^�cw-ܓ�)���ƫ/�q��Q��ț7x�}^l�?�x�l����=���:��L�������2��^g^ڠFMz���n���hÙ�>���	��L���n�k�yuR��txޝ/:�۵v6�8�i�$�N�_Fcb�]v��"�''<�'�/:��m��8�C�2�٫�������뚻{E��)�8�N���͸8��;{n�q����^#��m�	�מ4<u�0䶬;�@\A��,v��W��]�ێ�/�C�%�ݤG��}���a�]�<Z�;n-�k���;WqĆxرqv3n&fGR���n^{uce�����
���M��M��� �����sܦÊ� ��+k(�z�f�%���F��:b�m�Xn!0j�F�����W�b�;v��0 �v�b�{��d	9�槠�����> �Ct%���l�����" �{�[ Aq�k�#bnz�ޠ =���� sܦ�v\tīn2JnTPB6��s7]oj�<�=Oq� sܫ�;�y�>p�m�@!���4���&�f*�&Js�W_�?���٨�6w��zBO��Y'� �׹M2<�v��k�Z��W������>zbI�-��@4���6Qv�^X�y�%b��aA����?~=�sP����?>��� ����l�@��c��E�U�c%��3>_e6F/8�>(�*Hb	��]UB�J���Y�4��,�N����lKH�S��s��1�e�w�<������'��I�p�yY��}9q���<�����f�����݄@�^�8��
v;�i�(���l.�5G�:c��pp�5IΪ� 	�忓���:��~�� A"vvܒH���$�wn�F�-�L��4u�fF���}�\�RA��l��{��� ���M�ʛw]%7I��rz)pPpa�\6����ʓ@�;{[�������j�}{�hkr�H ���q�{q�c�^S�+]O|��vc���E�u��[�S���6틱���l�i�Q9y�}�c���6]]��߁O]� Oݖ� ��ۙ���f�(k���dr�;�$�Y�ѐ�P\WOuh��S�$�u-��,�e3� _Fgc��H������}�Z]���A_~,]����#B���D<ٜ�J	vwuX����F��e\*�7��tuG�Q0�+�����:�����BԳocp�y�u�=���P��C�qXɮyhC��мq����f+.�v�C�7� v{���]�=�L`p��	�4�,�멜]�� )��0��w7���'c�@����Iٯ$��۩����%fl��b�����"yN�B��ڇ�{Q���v� o��3 GM�M���'���7��<�b(p�*k�M���ݮw.R�ɚ�x��O�oE�wk�����˾��(������]� 7��� �]7�-���UY>�w��;��� ��뢢���P�An
��0%��D�S��U^���v;#в�׬����	����\XR0N���0�gDT��*UM�i�f, K�t�>
�w��5����� ��٘A)tN�I�cj�!0S��j���Tg�w8���E��� 1�<� ���o>$���0�"�
�����Ϲ����v���;�|-4`m��钫��͛%��P)���v_j6y8]P^A�Vr� �v�֏��6À��`�x%K:��( ��˨�͙�w֎:y�S��������C@%�v:a�EKu��̂)��~q�1Ѻ�.�[���۴ǝ�Ë�3��獄�2!p������I�\�m�b��^�|�@a���%6˵�6*#���}� ��ܖ�%��H�b%�m�PZ]�P�O`���˜��|���M�>���g\]�W��N\�V�P��4���*��J�?�� �ge�� A=s��o�O^lG�7�/�@�;4�1�Z��!��8*�:޹[�{�67����N~�` >񝎟�|�7�{����^X��I2��$��W��LAb"Eǵ�d@�;���vy�viʾ��ǀW7ޗ��L�t� on�8��=��^_�-u�]��yn�>�nu,��A�I�����L��w\�lś��� ��R\�i�OB8_0jp��9�X`��5�#��I��	��!!ۓ����WY��[�q�\ �u�q7�9�X���)7&6y�玓h���F^I�̠3ry-�O'n����ͧ�m���y��p��\��e{���۫n[�u��O-����e0q7�u�f��y6c�N���8�'[k�B㮸zӧ�s�����b��wm����{�;��p�v{z�]�Z:�U���_Bw�ۓ^�y�yD�kr��rrj8�LQp!��l=s�fF�����ꉚ�B���Q����L@/��7-�  ���ȅ��۵��wn�ߴGNy�L� ������@MD���(�ƾ/��b�"E]��f{	�j�@��;D0���y�T�OhS�N��1VhJR,@d���3�+'�I���i @�UH��Fӏ{�;%��� <gc� ����
�+�&�f����dG�w���c���}�Ұ ���π���iYn\�y�<�K�wT�$gR�E�0�p�Ak��~Iy-O�&�^�;�2��	Y��M@{�{1aBAt=���o���e3"���[t�U����n�O[*<�Ӈ�9��C�Ih���[��L"���ꪔJ	_v�^ ��%�C�� �oŶ�!�wn�- �vDc*���}8�y.��~��N�M�D��2��*�*���@:�EyX׍���'����%6n[�܀{��4������s�偹�&��y��9�o����m���� :kr_ɐ �uט��oc��Y��^�^A5QU@IJ�_s���[�[ �i�Bh�o�~yZ Gn�<X@ unSI�,�PXE*���j��6+<�&K%�D4�7�� uvS`|Xgc�=���Syf��ǹ ��ݺ67�e��i1*#�򦗉$�?N|qTCǥ��h��ĕ�~��� �unSL� ���L�GϏ��οo�e]�_�`��xb띻KP�1�`��ƀ���L��Yu����1s��R�_�ێ1 �6��πA���M ��m��UG4�>Ǹ��ݹ�@���6I���>�(��g���� ��)�W.���԰ �mnSFFu�&�F���{=wi.�ʆ�e7�D�}94�@���ץ �H������l��B�����Q���:ܱIN��wԜ�U�U��W�}�9���3:��/��	U���Ǟ�:���ֶ`�
�&gm�p�r� @%�v:�F� ���5PRcG>y���p�&^��h"!��ձ  \o��$�[۽}\ܭܺhh�˳`$���u�K�O0�a�ۧKM�UJA$���~s!:*�=A�I8gV����07�y��z�
��j��ۍnvr*w����n:�cW+e��m�J��USʝ�v�m%g����i�5??���|��ع��m�?u� �̷`��w�07ѵ����s�=���i2 >�s0>+�
STT�*���罘��X��:��̽��.1��[ KN�:i �;�{(��R�_<�Yuǲ��=����+E�!T(�S�q��J����� ^��ɍ�|��e�'�Hj̺tI#ݻ�F֎،eC`�����K���:���l��ݚ���߀H=��������ɰ�	k�ln
�Y	ո�P����i]KT�nla�Jm@�wr�f�z^�<g-��\��e��ڨ�YӪ<g�9Ҡ���cn�v���=2y�L~�O�XІ��k�&��b�$����f%��H#kq�n�U8����;n�wv�H^���/f�ţ�C���G����c���6����0=��^�uz�I���P��m�`C�·	�D�ߋ�m���i�@ۼ�`mnS�#}ώ��yv�j�WN�@�7w�0��zK��D�%SF�y�lAh�͙1����a�X����� �H6�)�DEz�b;5�y��I��.�p�K�of` �����g�L�)̻�8����Ey$���&��Z/�	���S�*;[�����'A �uc��>�չM���]uGT�3�����Iݽ�b�X;c)�0SpX5^J/9�`��-�)*y�~��a%����-[ny���r����~�$ I?�H@�� �$��@�$���$�p$�	'�@�$���$ I?�	!I��B��P$�	'��$�	'�@�$���$���$�H@��	!I��$�	'���$��H@��	!I��IN�$ I?�b��L����΂n^� � ���{ϻ ������ �                     0 ` R� 
P
 R�((��JPD$�)A@ ) (gx���*���"���QUR�*�P�*�T�QT�*��(H�, ��)J*�*�����N'@g�@]�T�Tq�u�Lç.�	��/9*�)��y�tk��� ӆ����J��y���o{8)���z0��rU��b���F��\U]@ �}��RR��AJEw�M���7����s�ná���{:tn�.�t�uޤ=�k^�W{���(| ��OZ�M�
=@�r�D`P�����gl��R�(x�|)D��� �C�T�� 붐V���jC:��z׬)Z ztz=;��s�\�R�9T)A|t����-j�c���@i�@��r��ڎ���T����@h���)J���B�TR�H���}j���Ǭ���������փv]�9���$�O@��)@/��(�>�Q�wbG}䋏T�bf}�� ��z��|���}��U�}Av)�;�;����^���� �
)@c�E �UT�T�(V z�E@ƅ�P=����}��*�ޢ<<:U��f��9���Vy+CA� *�_� g���	��3�wn���Zyu���מRa�m�U٧����iG�     S� )I$��   ���JT�i� 20  14�OF����R14bi��@d1@@��UJO)��       5O�!�U4�L&���LLC���i"j�4FC)�4OT�&��z56���~��o���I?�Ɤ���v��>��$�?H�$���K 5��H$ k��?�$�� no�g������� �A1c $	�<�?�� ���!�`�@P0 !�`I v���N���H����~������@�<�!>v`Qή�>�3G�-&O���PO����YK����>���۟]w�u����fvbd�����(�*��F�ٯhZ�y.���� aN��o�&�F�"2��k��vi�Ƈ��wu�IO�M�u=�4	��$�.��K���Vrky��]����$�lk:��H	t�wO��9hǓhC��KHo�~�6����77E{*�yU�F��5N;���;�ۀVr�);O`��u1f<Bٵ��}t�m�]����)rT��H��'� �^hA��,�[�w��2���p�W9S��:՘�n�FI*O�w���Ӵ��Ph�0-��}x���nOS@�PZA�;���P9����%��;6b;��t�������;�3��0gr	�`̙��S;��gr�n��2�R�c�sXu���p[���7m�
���87O7���&)u��rPE��t�����8�7/gq/�'��	\ٙtv��n�X�aF�F=Ӛ�m
!��øWM1u�ڼqY�\�.:��Jt���2Y�~gV�^X��5�IEEԗ�7Cw �1����9�s����BG���0�\�f�渁�j�c��6���A[&�!F��dn�S�6R��n���(	��v+�N,�EŝB���w^��ǃ�yٌ@�=��]��x!oAm�9�6;�!I:\ko�b��nP ��=6�����&��Xo(��$<a�e�Xq�"���b�5��.MTͦ$֤tc�)m��L���ʷ��t@��<w:n쫶��P�������S;Q2�@c�t�C��p��)v�ԁ,q�vغY�M|U1J���,ټth�tMqы�9��lz��7n��n�d��ܨ���`�O��m�y$��~~�=��5]��-B��������8I�r1\�3��3;�8��Qq����xe�{pk���G^q��S�)�Gv<�n�M�'��"aAa�L|���[/mH��d=W5�t6����KWk��Žw7��@:bWv��w�=�uћ;��w8�ď�����׬�A�g� .%g;�ck(d+�'�;/0f�wWj���t�|���{m���X�1"�3-�׮|5� ���M��GBf��uRZ0e���\��O���
����UC{)YݠU.���|w��Mo�ib�V;�$��L勑�f��.Ŏ�]e�j�:B�Ǚs:��p�A��"�Bb�6q���(uu����f���¢�U�f�u�=� ɝ����@�P#9>jin��ҁ�Y�����V1���0�S[�.op��T��eg��f�T��ԮA븰ޫ�8+��A��qWܔ�[�̉�s�T�qӝ#�U6�P��ձ���f�5��]�GɮӶ*�-� ��a*i���\[Lٗ����}�����i�׃	gPe8�5(-剜/"���58�^��2Gy���r�W�%�P=9�/2���۝�oF5�sfd\�Rӧm+w���M\��^Xì�Űi�1���:L��/6X�7NZ��\+�dyb��|yi׫6TD�m(��@6���{w���b��[3�G���xmn2npY��٭#�w2n��ԓrh�^�q�m���;;P���ֳ�-aYt=�|��^J8el���+~�0�ۆ�m2I�Ƀ0�<�֬�6�����P0`��U�:�W��ܪi�A˝�������\�c��<�ۺF�f)F�	U:G�4�g�^ј:.�$,�N%�d�f�r��.U�{c���^�Ȝeμ���gZ�y]�N	��U\a���4��ӸbU�6WI}v7�`��F��n�  MQ�zhر��q�����S�$��on�#7w�o9�:I�ʻ�o��33R���#�ѣ�̳���/nf���.>��vl v�3T�<��fp*v���6���~��@�wm���[ۺB�O�ܧ�Bgs��5=�"���cue���x-��e�^�׼��(���܇^-��{h:�-)JwnD��j����1�G뢬g�)�Vi %�`mS2�{�e2�:���p�14���lI�G�wl"m;�{]�Ǔ��r]ܗ*75� 7�k�r`hF3��:!�h;�;�ssrN�Y�6V�;�G
�c���ƨ5�]aX���!F�U�(0b�{�i�#�e�ŗ�5�v��O9�xD��A�`y�	*�G@>�X3��j5	H�5�b���&v>V��]�-���=�X�d����ǝ7������`;Ɇ8vu����v��y23l����N��.��� �#n�ͺ�k.��T�
"��P�F��)ή�t��ڜP�ieI~����Y�^8mLF�8�c�LkqӰ|�.x��w":���:�����gU��f�f<�Y�0�7l���cC��O�����5.�dá��䳇�e�T�*��w��?�/͗`�;�K����0�]��N=�s��_>�0ϐ����֎݂�ܙEiU�&M�X�Sy�R�:�.�ߓ�3��՜	����wze7�l��B�f���0�+ndū{���=���e�q.3+���{I��w��Q<7���p8��W&�q;�!fiD�i�c;���c��pl�4M�)5X��n����+[;�C���g��'B;�r�`���۴l
��yAO���N�@:���E��;;;��8λڤ�As-��O�;8�j����ƽ�a��� cu�[HӤ�Xr^��u�ٺ�Ļ�x5��ۼ*էK��Ow�y�3�P�Xׂ�/�d�FQ4�\��m�o���B-@���\tˊ�7r�jѬ\�8�v��{e�O�����%��n���L@�޺�'u`)A���-HJ4����0��N�v��+�c@���.y�EoWU��n�ӹB�qQ�v*��S�e�n���G�^]'.K��~��&��j�5��x*ANܜ�a��͝�N-�";5�
d��`�WJ�wG#�N����z	Ǜ���ü[�敆/M�2�+����9�Be�:���`��>�G#9��죦�������L���$�םz�}+�3��޴b�����$�`��x�(��D2�O,o���/�;	X�#S��]7��뺇v����5���(0L`7�I�2�Rz�_W�h��E�o0�T�X�թ*�Qt���>���N���sbG��7��S��ɻ�(pL<,��z9���Ǭr�qو;��U��ޥ���*�9�.�`9FmñǷ����e��G0�;���7��ٴP"U�h'b��D�MM�zA��F���8��F�R�la�fX�f�%W�̩��w��78����s����{]��������4��j����;�l�(xF	�pC�sxze���0+�����7��P5� ��cP��Qx�z�a��'tDh��b�ҍ�wtwf�A��v�B�L2����k��!
�%�rh��1S�8��aT�{{uM��g,���"��w;R�ɷ[c �`��A��4���u���c�u�hq�#t̷�CV��Q������V�M�ХAo݆�f� ��{ x݁bM���P8�����N�[��n�>�.}�P�����;[ĩ��Wf�GS�>�871cܳ:����q��9��q�|��N�һ��UЬ���8�Q��{��o�/�Q'hV(�Wl���;wjr>�C�=��Zi�x�u$�YD�rsNm�qv��6���h�O-�#��obX��3~T��ыwjք讓ٷ����=��M�v�)칥`)J����*&�0����5�AH��l��f�ݣuf�4�7s�����d�C.���jj���r[��;O�y%Ť�v�o՝v�Ưe�p=�WK�� 8���E�K��}�g
{A=\X{���U��CK#��Z#�qj�©:!�k�"���� �.��k`'0l�Ƈ!۪�5�KL�0N�gsN�.|q�C`#��*��2�Fy���k�{L�On��3xE��ɻ�Z�[0�\^ҁ�2�4�*l:��P�Tה�S7R��<z�l'9�u��;L��Þ��j�ɑMoG}EE�t��r�C�,�;� @;��'+���<�L�lZ/t����<�v����W\����I��[��|r:xr��0�8(f��<�;a�\�˳!��:;c�$��n��<�ю�θ�T���9�ϊ��U�rM;���ٔ�k7�poR���b�#8WKC[ߎ��׷)܈��s�<�����y��<޹����g�:��:�Fd�P��~����a�����wGOׇ��̈́{�� �XH�$`H,�(�(Ad�E�� @�P����H
HY	%HBV@��	 �@
Ȱ�E!TVHB��B�
 ,
��X@��X@*I,��R@$�H��PP	�$�d�I*B`I
�(Ha$�d��!R@YABB,,�E ��I! ,� ��`�$!P!$�,�I$������~χ��o�>ߴ���؉�$H�&��nBI! }�|� O��8%S�S��nH����3�������C���Wd���%17�%.�TR��
L��B���e=�Ǩ'�l`bh�q���bz�݆R��>������Qb׹bR�A��]�k�tS}GW��\�y+c�{�8��X�b��w�E�}�D��3B�#._nz��ףݽ|�q8��Rr��������;�����!쌁/n�����˜�@���3��!D�P&rbw��A��{uy��_��3e��)<~%��Z44f�Wܘ��z��8׼�f�\��|�~~Z�g�������d��yq��Y��<�g{�8��w:�_r�Ɨ���`=پ��=����|�^|^��G4�%�u�j3����a��0��ӯ]��j��_`k|����[�eY5a�����Gw|`�%��3m�&�@�w7'��9��p����8|_�ݺ^�{��E�y�&�˷B:x̜�J.iS�Q�;ޝ%�q�A��y��@��.��Fe�`��BV�9s=�|�c�v˷��E�DB}���c�~ثp�#�-�6J���"��#wڔl�#�έ�r`Ι�L,N��Oe��O2�1�2��3_�W��'�9�ta)�����Q6�V7���x��t>ܽ��̷�q��n�ܞ︕�ų�d��<����Y�����v�U$ܻ�|_vV|wx)�Kz-h��']��ťp"�S��X�5���ަiԗ��`i�#�l����hYXۚ}稛;�w�F�7yxM��}쇆 ��r�w�p<�A&��M����sn�
}˼f�azZ|��iq����q��1�\��O�{�C�����{��'N{���ކ��X�����9!�)�p��}��sG�g8&�A���y��^/k���ó���1{c��Ro[�=�dsټ�Tw�"�ddm@n[o9��>�R��=�9�V.>MA���3�x-��/qVc�Y>�:��G�o�O�z{K�=Gю��_OE��K(q������f��$EfT�Q��Қ��Y��7s�ݍ3����v-Ұ��W�1����^�����pܾ�w��4�����u���૦��Gvu�#H�p��50���&�B��}T�L��EC�B��xZԚ;㢼�P��O��̞�Ro�_�힧Oq4��	c�^������Ĩ��S�=����t�cd$מ�6�Y�!d�=�����KqW�+�f�2u��<�x��aF�ӹj-L&�Ap������#�� ή��;pvu�r��� C��F�Gd�S�U��R���FNKŗ�&݌�y�ﮗ���{
�{{���'�o}�ˋO�&'��᫼9��/pxȊ���rݕ���F��梓g���F{�T���ݻ�*:���:4�a>���DSsa�G��5u�.��;�e:�`\]Ӷ���(Ōw�z�v��_0�ZQ;���ty��ct���]�[��d8���;�����y�^~��/��<� 
:�W-�{���Xvf�=�
w��{p�������t�.� j��X��\B�}����]�ռ�n�;M�^V��K��vYp�r�`�Q{�#dB7i#kN8/��]�팫f4�
�����魳�ޞ����׬�C���u���[��1��,j�g�&g`]J{u��z�%��{g����{��K�]����=�̫ �Ԍ��'��އH/Z���EJ�,	(~;�
^EbX�d��{'����Jcս����u��(���)�3�=��c�HY{T�Y����D��Fm�r���z��hl��Psjq~^�L`�;,g����r����p��Z��NNZ��R���{u�>G�O{��\�������&o	��L�Gb�G�����36y'���߅�JP�MWb�P1xS��{�<X0��H��OD�=���[��2�jem'��ϊ=|�K�v�u�y����z���������_�__;�Z�'��.��8ߊ�r�%_{^)�=���sz\YԐ��B��ۋ�X���#]c��r}��W/N�5x�O��'`�I�e~��Q�I��R�%<G�x��UZ\�����1�[�:r��u���T��t���a���+�B]ᾗ֐w���/&��q�(����S��Cټp�,"���u��e��6禒�
t�^�P�`�����>�ۡ���Pa�����K�y�D���!�}=*FzN����<��6�g�r��i���oW�Z�Jq�z��=�?5d�sf�+���k�ql��=�w��rJ�F=ŻF�F�{��2��U��B}U��(�[��DX�� ͿWM�^��٦��{pۡ������]�Ō�I4�휝�:��l����q!�<���[�}u�F:7�u�GD��F��,=�ܽG�z��9��.�^M�'��ZC��2��oH#��rv��«�ݡy���{�P�#}����ݝzow�������,A�˱P�($qb�ϒ�w����E�GgQ�C��ѩ,Jab�df�}�랏�wb��+�~��u�W$7ǚ�F^ �O ~����
�Ĕ��)y�x��ԁ5�e�@�p�Y�ṙ5\���
-
n�鼍�9٧8�}����ܺ��@i���SV3�}٥h�|�h<� �S雭�Rp�uc�(�7-��,�)# #Q�M��	 ��s�<�2�������Tl�`@�ɓ�6(��R�"q���9��^�7�*p����_�M'sOsu@ڹ��b˽�b5mӨKa��F6֭յ�՛ݍ����G#MŚ�Y���(4�ƑJg/[k7a���m�=.@�Y˟�K��m�h���oM�B�o�Qzxeͭ{/��I��e��������g>��q����<	���rdl����r��ym\��[2���J�;�țں�/3]0ѲE��*1m�����jt�H����9���ID�f���4�r�辫��w.>�=��:�\l`ޅ�S�Ռ@��Y[��F���F�������5M��t�ͧזyG؁ːo]��3*���
��yH,}����,O��d!l̅'`ݛ0^٧K�fw_���icɂh����}�R%c.����gr}6e�|R
���f�=B�GzgI�vJI[����� ��X�=�!�� ��5��ť��p�47r����d12*�u�b�T���G�95�����{���Pk7|>�1醟h<��(��rԴ�������u��BNd�6�5w:�9�~�"�䛃�a�qۦ�O��C�t{�w���p�\�(��	.��������`g =
�u���(�>=�8��޲�	��X6�TY�o� "+_kq�^��-�V'B��[1�yd�*�wr�P^����^c�K���E�IQ\��S�'����Q������˽_��x���{}�uq��I۩�٧��,�Q��.AǴ^����3����ɏK=i�}x��b��W�3��g���-� =���΢n�V8{ ��s�6]}�Ӈ��-q:�ˀ=���Nk���o�'��w��h��H�}��Z!v�8t�#��:�f���yt���L�M昸��*���ɜ�� ���,��3�J�����^:���YMC@�k�o�������Cw��zQ�?ei�{�M�NP*7w�=��w"��i��^:��W��|�龻�9��Й�����/hZ��ת�JG��<��\�q~�<w�v:�e�q���9�v�!g�".v����λ���{4��|�ԯ{˨^w`Y��y��g�����:>H6��/71Ճ/�WàocȬEd{E:A	s,d��888�zw��5WȲ�(nn�n'���c|tr/�o"�K�cې?y��mY�;{���R�a�nQ
􊵷X3R�bhR']�L�x��˘��]c~�>w���!�z�!��X|�g��n{:ν���ٰ�|ڎ��c<b�.����'���\u��7@Bx���ٺ��IǶn{WzhZskfa�����y���5;�ӘG�e^��U��4�A�ɘ1�|��=��^��þ���df�f[L9N�I'qǒ�����r*ӱ%Η�8�Y��v�͉K9j���W(?q��ؑ*]������|�Ӏ|���g!L��e�(}�\t�J�g�p�:p�N5�/k"�Sw/L{�d�}��m�c�/�%SN��A��ԕ����e�u${�u�%���~'ݴbR���G��Ȁ�a�۪l,��uyO"_�熟>5w����e����k�d�%��$9Y
��b�u�;��[��:^xJ9=�_bX�/W�7�����z����>��S��T��Ӹ��[� �{��a�Gp����wO,�~K���c����(i���뿝���}o�O� �$B/��!.�X`���>|=0�`e�v�}ʰ�3v3Hک6�tq�uW6.��p�4��!���q�l���39"�\t���ݪj�h!�J�:z�Q!����ISk*��ͥ�`�\>M<��t�ꨂ��vMyp�1+aͫN��Α�#�����Is�T���{I��^����j�ۄ�R/I�b��������Y��1�\����J[�l�d�X���s��]�6	�xJy�p���g"��V��]C�V��Tm��s)�����ٱOm�C���[Q�ʈ1��Y�[N!h;��Kb��2��4)sԚ�n.�s�o<�
W�>�g�y���t�m�qX�1iv��]��v��F��D���`f�j�nqHjB��ۆCǎ���6��g�zt�dq��м�]��'&х��d���<=�{�8k�����-��gGZ�8�Z�B�gR�x�u�f7W%��0k�E< �o n�v��֡/Y��@��T���ˠ,��f2[�Xns�c�dwm;�`VJ5�j��PLt! ��#]�nu�=���WG+v�t,cu2ј� l��!]I�.͔�d���+l.%ɭ)�bĶ3U��KM�-��Pa0jZ���ئ��ba�A�X�i���m΅vM� lmt��jPL�:���,cP�0 ����D[�b=M�8�[&�6綍`���;M�zK.�]q�������;R��5IPQ�l��5Ѝ��^��+m�����ͱ�)+�UAx�Zjͬ�.��Xd;S���v�<R��t7;�'u�OB�f��`�a����=�wS����V:�4t�e��6�Hlk���5[!m��L=t�r��.��#�j���;v��+`���\G�4�-��0�%YGA�M��˒\ŋh��D#�u*�F���;�^�g��/��q�4�Dn`�ݝ�w�n.�:JE[�d�-]���kC�����2ݎ�wJݽ�Q鰇>�1��z�j����+z]�g��=;pn)��\3����T��5[p=T�۱syn8��!a�c�
����!�iMKv*>�y�k����wv��3��ۙ9��2�iH����9]W�lG�ַ#tv�]�ݒ�//-��ϳ�d�.���{��㌖7��Ŋ������l�l�a����fKڸ�:�,, f���lP�4�f^N�3�wGnծ��8zg�q��6xw����mv�m`0�[6��nH[%E^Iq��v�.���v�����m��7`6Nm�c�v񹵌�\��Dt��`�	j�R��ls�K&��y������>�H��F�T�j�0��mьGn��m��y8���&b��l��,1�fĳ.��}�����+ ��Wh�	�C�4��\�t�fc�A��[Ecn�Ȯ�8�9��u�'v3!R-j�6q��4׊#�CjNo�P�:���C��8;Y`�m��p�{psv�8i͚iQ���&Ύ5�l��8�Z��:]�n���qf:
z�ub���-�X�YZ]2ػW�Ԅs�@=�"�����ִ7u�Le�Zɚ���vx�8MއFɪ�E�R�`���:gMFj��5��3P�^��2%���F7��v3�]��.c(UN6���4�h�*��-��P����Kq�öp���Ή���&�ԗ�BQ��.X�+!d��^��0��!a��`���f�+5��64W�B�!p@Ь�ZW+��vWj�i ��"�v�cv��x^�=�H����%uka�m,�m�`P�Yf�# ���]�k��ͭ-G�7�� 5�L8:�+ě�\��:�9EQv��ۮ9.��ޝE�m�%@�WK��P�Q�:�L���ӭ���(g�-i��*[-W�u6*Bf�]i��9z�\m9�����iJR	e"�v̔Z�Wr4l���h�`�F���f�6������Ρv��,�&0=��v�L5�nK���ƞ��bN��v�tT�Kt(��"f�m JҊ���$ܸ;�6:y1`#�#ź�Q��=�;��'F�N!�[��-V�Tk:��|#I7/ldzm��d]�X&݄]��V��)��Z������uv�9eݳY��M��P�-�m�+,�`E3*U��4ZӲV;@��7��Xp����']�<Zx���t���hx�;er]lɝ�F7�v؎�&���̪����k��lqɴx�y�W$���#-�k,�fS���aq�<��l�=��玶.�7`�����3��6,g�G6�X�����aAж1v7�"�Gm�z2�['�D�0��6�q4�ƱVk!��؍`������۴�tX6+�g�Lݖd�RaC�M ��zɬc���fl�c	m�2��kb�f�Ǫ=���ζ��ON�O>��\c-.�6l�A�Z�1�D�w\r�w �1�3��Z�v��0@�;bcV9ի�q�q���[��TY��e8����k�lr�u���\���,�6064e�e�n�Ĕyj���ru�n�C�ny糟n2�\�!�6І�%���P%l
f̅�kIT�X$%.f��e�ιgZ(����cm�X��˛�\-�K�����#7ew6۴=0���`��;��c�芋,���mk�@�tu�B�:�
AiԆ�c�[B���%ѵnA��Z����&�weF.�Å�vBu�6��cQ#`�F�031%�.��I���պ�u)�mU��HTV:.&�F:�8�[��监�st4UMLRR�V�yp���+[���L��6��PXd��Q�XL��[s�#Y���(!4�k�۵ͷV���N�3\�[�NE"��j��j��f�����=�mE��jr�ۡ�b;�ە٘�k�M]������8�Gn5�'b�(U�n�[�E�k�+��Bج�kp::鎃<X�:�){k�U�b��h�f�W*����ґڊcJ��d0͠�J��i��mY�S�p���څ[g1�9��xI�6�s�$�ې��fm��嶆�u��1	�]�If4�&6�X�q�,��\%	j�)fKq�ڇ��N���{v�g�9�ɚd�J�J��UUU~����^ppz��(��J�01ue�r�-�F6��\LƱ�2��m�T��WXe���X�����FեB�kS2Pm
�)�������J�Q��#�Eƪ-ۀ�""*�LkVX1AUE4�B�*��1)2���Eذ;j�"�rأdZ�*��cZ���v�I�T-�Ub�1X�U�YRQUV+c���R
�Q��TXe���lDAb���s02�,b�,-�+�Ŷ�E����F ��AX�UQEI�b�Q[J(#��b�`���D��wN��ɾ��,����`P�u�toE�pA��;z�e���{W<U�t8��J��I�b��`��'oj�b:La2ݞ֒�ħj�5���7����){�Oa�1��u�ٻq�Әx}X�n5[��4�B.I�s�a�c1-�
C�H\՘����(4^������/Gb"�f�2v����8|F��]��9Nh;�x^��lօ;��n�56��Gk��Ig���#S4޵��5��֓vq�à���tٮ�Rh�����F�N��a�4����|׾p�ۅ|��GbN���C�)�/=[Jb]!�RcWj���LXm)/J�����Y=<���;�[[�q7Wrb�Vc�eZP��A%6�m�&sq�zu:Nc�9l�7#O28H��m�;���q�W�o9�y��j�6�;\�)b^��h��	�?3�o�_V�z	��6�Et�����!���[oh�D1�5���1n�t��6�6��a�`�F^p-��yr0�U%�,��ny��6lH��W`�l�٢�.@��K�pWm��CqWM#Ul]qpW`��gi�P�-A�w/��KZ]N���q1�EF��t}I���s4�^�g��`�ƛ[��^���L�Lm).������րX\�r��7*�3�r���)�vxq˅�ܠ�vx_n��;�#��n�]�9xNWm�vy=�A�/�8x�����˳�ʣ��"gl&�xN�8x8]۱�z%	$����?/��P�R�E�c�W n�U�2�J_t́�H�ٲR(4�}4�R��NC��nH ��@�s����k�M��3EA�ڪ.`"OO0�1äSɞ����@�F�-��R��BB��9�y����ѓ����5v��ԭV"	}��;P��;8��_={^��7��ʰ@scM ���g�J��i����f̱��\��.����i�Ȏ�U_>~y��#��=����??���W1#�$I�����V��7�?/g�q,D�z��1�P�b���`?�x�񽣚�K�_��~�,�7��O9����@�#��L���$��y��	NZ��A���TD�s�
,�u�Y���%��3%!��.���U�o|��1��y���;�Y�=�>%�͹I��U��c�ł��e���ǃ�)#�����#so�tʷB(�aa����h�$(-Ƹ�n�U���|��mX�!��$��$�����K��;"�W�;zD��h(��$ܝ�@	���Ι ��O��B$�����0bV�ª=ՎA W�H2*��ƕ6.��6�)fݠ��CV[�\r��P(�m�L��Vll�סmyl�*'�w�"H��FY�RPH8h>���r�⳺D�H̅`I;���m���o�g���+�]m���dmuT�fJ��#L�x�}���a֩�%�=�భ�&�qAU5~}��}/�=��]� �;�I����p�u-���|Bz��ݢ��oTs���=�7�Ēz�"Nw ˊu�Y�Ӓr��U��Mώl H"z�;����V Az�o0Ȭ�c,5�C�m�R��`JӰ<�}������^*�iU��B�7��ɽ��r��'f\;��K+G�.�TEω4�M���	���[�<Pé�v�n@�r�D�	+�LS�:�2cgO���S�@��t]⒵���Xh�v��EU~O�Ҡ�m`N8GO??ow1o�&&0�B D�[\��/[�����&}�+��Ԕ��[���9�ίP�Ut�9�U�MB=93-���n�q f���`ox������J�p���̡fq�G{&`�W�� ���h����M�� ��b�G�_�����$�=0*�}��O��nc���k.5E��[�S:2�j�k�o�MTd���tqBP� B!�0�~M�����ؽ���2ۉ��!�4U�9��ug�gA�x��u��"4h��q�ͫݮ����;K�O��bT��։q�i�*J�X� �����B�a�G��k%�g44PK���`�0vp�.��c�jd`XZ��5n�����ʹ}�/ϗM�]�^DB��Ł�� �[��!ܴ�I��E0��E[w��ʰ��yr��؀$�qb�Z@����L�Y:��r�z�
���D�H#z$�����z����� =*��[�U�M�'����Z�.�1b�h>Io8����cY{MI6;`Ӂ��Q�Q�g�c�F��9��\����y��b!A��Onq�I�ص�]�5Ȕ'�m�5�#42��md��f��h׫&]��\z���&,!��ѮH8ht��6ll�F�M�����n(�En��{Bx������_(����c%Q��4��ޒI7P ��l˱����;$�z:�BkXϵF�D��d��y| ���\�^7H�����}��aW�A�\�lzL�|m{5:{���,�>��wM7��:�I����ƈB�"s�����f"��Ք�y��P�0w�mR>�ah�h����U����z��I��Ɵ r�M��������pY�����3)�G��}"E҃dH ����3�d�zn��hef�h�����L2I�ޟI"r��G/N��}A�Y:�e��D�j��yx�);�l�{,Tk�Ė�X��P-�$�k9y�wK}�xu��&�2�tQ���xI���N� �C��O�K	����Yx�"���f��_;űg\��vy�x�@�"��8��E�)4�a��\ZAJKftnr�3]���7|�l�{���GGكq�-���ɐj␈��I�Q
�?V��ʘ��<�G�+��Ru3�tE�E6"�t�zH"͐��F.2����h�� �v8�x65�	�Q��3��d�g
$�sx���)�R(R��u���	�+워��v�%��H��s��r���f����ĵ��H�ywA���X� ��/ә�u�٘"T-{ѧ���=�ϝ������Y�E�npRh$m��u���0�qS��ă�D��+�v�S�֤����%x@�4�������TJ�	-�(񲏻y�I�qy�	��ob����I�|���W"],��\�&��I���'ႛC�m���sA�CAGJ$��A���9y��jL>����NQʙV�ӧkٚЌ�G�k�X��h �����<��ӻT�R�i�^����\�mNl��z�j��h�eu�W�MDfw���i�AI!aIp�D��N��p\�KCY���z�O�p�K(d����n�kĻCe���b<]�Np��
�u�T��Xږ�31�؃��	��k���y�=q��ۧ=/=1��҆�4vt4P��.U����T��lOC`���0\Z4�K��6����{�<\��󧫂�?F��L�_9��r���ag�)\rA4�D(�>�w�r�>��A���2y<MeXq�x�\҈JnB����}"}7;�|!�� ��k����>5u������p�,2�;��Sm�n�ԓ�����J����� �6Er�k�=�� �^1$��#x?�������ү냪�5�-�e�Y�lV�����a��6�F����B͞��	�u��6��NN��Z��n��{��b>󣏽>��?�]ّR}?yz��Q��]�qTuނ�!N�9G��5)s^���"N�(�VOMR�ήh)NB�%d��H�/��]\��=����s��J���.��o5ET��:�Xe���R�P$��ط��vh@����@�T�E�
��}ڇ��7l\���������9��`̝̈́���B'�e��H� ��՛Q��l
�7k����>|�-�\ͬbM�(�o6
��34��s��Iåx��N�A���a�u�f������(�{y�U�B�ʬ]۔&����m�ܬ,@�R�?�Y�߼|Ndw�Bp�#�_�;L<YJmf��N�����_`��Ž��X�t���ݝ����E���GRY\ݝ�,���+��r{���	�wC�Z�U�G;|�O��
No��$bn>�����=<�����{)�~�:ʹ��4��Ax�tU�ص����z	y�x��VL8=��|�-zm����M�"���cv��Kv��n�6�I�3��:B�������VXo������8	�؃D���s���T��D���bA��S�+������G8n�����8�����Xxw�޾7��v��gm�~��-���{Z��_nnz4#�+^�oK�g,]�l���aq�m��T���\ݨ�ｎ/k�i�-\f���N+�{�zu�k
�u<����%׉i�� |��1d'��!����'��6�0��|��IO�ޝ��+�t�ǣ�߽�i���>y�Һop���tak��[k�B�D�%;�}'=�1���f��g�x�G]>?5�>zpd�
du�R,AO�Q�ڈ,D<e`�F9j,��T��UZ�",��q�"���5S��cYm"�؊�"��B�b(��c��Z�X����̕PX��QU30�Qb��,҈��kĪ�����[���J�Ls��"1M4V�)�Ym�lq�U��D�֬��h*�����-Be*!�feQ�F�w��̪V���a�����T\�E��Jʁ��X*��6�Lt��KK��U"t��$��a�r4�;Q`��b,TQ٤��ʆ88�F"��q4���5�TO����(�~���H)E����j����������G�}��~�� (��y4�!CU��'�O�_Lث�FM�TzD�A���&�D��ѫ��!/�k���4��ٛ�RԚ�RM6�w�b>M}����S�$�y�3�P��U�F�>'��S���-�g =�c�kx�68e�2Q��=��I��s��N�A���O̒��x��c�o'(���=����S��{�Xgol�Vi��h�3 68�"L��PZ"#O�v�0��GK7{Q5sfn!����\n�C�U9�8Sm�l��M8y�R�М"o��(��IS�H�H?� �����[�4�A�l�,(٧9�4��|*�����Fw%q�z��6�q�s� ��n�7�D(a�/�$o_H�I'�/U1���ۙ"|*�Q���$�ށ`��.�1WW+	$��Gt"JM�5���Y8*,r��&��VL��ʰ����s70;ε�IVw��jA��L�c]Zr�'\��>��H$��+�M;_\�!wa��न)�@'#r�"���ꦎr</z��o]]h�隚)�<�F�i�y3^��t@{��y���H媻'3��9t��r��_�K�ێ�?�����������ƺ�F��h��d�G���P7�5���轍tp�n�ol,c
lI��cc�:Όvڗ��\OWW�̥$����u�빺�;[D�Zl�ʦd�7=,�z�Anj�$1tf63�"�[+%u����Z�0R*̴Ur����M�Ut��w0��V F���w⫯�&��)*�}3sn���w�����Í�]�rA'�.�$�s*}f�}������b,8I47��'�� ���a+Y�w��M�  �sdN
��Ű�D��xC�瞰]_�!nF�}&��6a�����2N�P�e82��{�(H��LQ����7��$�wH�1�	�ݮ�>dXG���DCE�Kb^.����QS__����Fi�7PF��b�7���J߁쵑��f!G��<3�y9�f���{[�Ɛ�?L��ze����o��T�qc����$��oğ��8��L�"E]�(�P�UE� �u��A ���7)�@�;����V��E�	&��FL�˻�H>�� ��ݨڼ|��+͢A��ϯEE�E�d�ޫ�>��U�{��zq��G��X��d����l>��_jd��f��U��9��/C�t(�5������Yn��֚���$�2��Z9/�6w0.zQZ����Zn߼���]y2'�=:�SS�J��h)NB� �Ι$�;�D����EF+���t�97w�Цʻ�����ٌ�7c��TV��[�}_㽜�'���Q���.�Y04�9�H��D�HrU�zOl�=�z����:�t��'I(��@�:q���	[nQ3���
� ��n�X,ls��S%)G�%;,��,�݋I��!0؆�۾�	��r���f�D��B�S�{��jj}>�����A2�����X�=v����}��b=-4j��k�!ӰJ�褡��uBbJ�������Y��; ��(�N�0�H)NB� ��5�q���(�H$f����?�J�#��@�qW&n���o��֍��/��Op�,�=ʹ1yY�kj��sP%v�dn��cN���M(�Pý�9A?93.���ך
T- �-2{��N�eOZ���i�,C���h�p�����mn~��vlQ�����"�zCݛ3�K�$�'�Q�Qp�5Gz�D�ד�Y�[g
�$�u��{{��.���=�xlD�իe��۶��6G�_������<g�h�9�3+��wwM6��Vz-���0)���*�q�Rk>ˎ�;e�����XY�r>z�nr�g9 �<Q�}t��+nҭ�S�4���6�(ݡY�⛮p�&6ݑ8,��M�fe�,{@��'v�3ns��|��J�cKqX�b�Y����Iv��M8�Ɗ�^������H����Ʊ4-+.�̶��ȍ#�Y��gh�4�kDt�L�J��"Fl:���#��k�Gn�Ş3�5���Ԁu��K<��Ank�+�#�x��qh2ˆUl�f���5K��\�	���3�_��a�Gu�	��~Fw���'��d�07�Kh��V}*v��uQf�}���Ā�,���Y���u����I��;׎Al�C̹�gK�Z��6dt�^9�����L�9�{T�r<@�X�V�E���EWd���)Ba��p�Ir78�'�-z���w70�։�ߝ�o��ogV�����.uX�s�4Kr�®_��|��K����Cł �6S{���z#�/���BL5!w`~k3���΃�Y��k�^�c�R�7�6ǧ�Y���yf/JP���xf�������� 弎��ttEE�-(�:l�zq2@+�;*�b���$�qd�OD�xX���M����FD�K L����h)$˧}6r�=��h��'��[�3:���rfnKA>����;$�ι7�j:a�Hi2�1������!je��������n�z�D �-�{�b�O�9�}ue�k�lbA������}$�m67b�s�"�Aܶ�7��A&�eU��۹�f��T�!&�/y�N�� ��B7H�-mx���C���\��E��(:�#M E�E]�)m�oᙧ�H"��#>��B�*.	iDOG�y&���2D�6�9�5�*ƮwϽHۍ>EQ�Qi83Gz�D�l�@�fbjFw-�M�������0e
����cc��t�^�<]���jm���Ij��.�F6{0B>�AC(�Rq��I֫�V]մ�y߲��s�/����� �+
řے���ySB[h�HIS�2:x�H,fy�gven Nw0P����ꪭ�[���6���w�W;1b,�v�/??�g_\�i��CW���1=��-��s37bEX��wi*6cF�O=9FwV��|���d��(��%�#�� �8��~�U�s{�M�#��3����4LyB�p��pPP�*'0���,�(�7��}��0�d^]�$�6Q$���l�T�W:�������=�;V��	��g�}���y{W��w !��|zKM~p~wn��'�Jۺ��ow�,Ѱ>*1Nrs�NM	�wdq҉�'{���	m�aZ���;��9�FX!}���#�;Z�+�xH�¼L��8��Ê�_bb������5�"�6F��{�j��g+Փ�ɟ��.K����gh�v�=�dm^�zQ^�ݥ�^�e���h���-d�v0�.��P4��K���=�=�H�q5�{ǽ�����}���
p6�a[��3�r�K���v�X���s.�x�(��[��4n�������綻������Uf���X�s����=�<�zh�j�<�r�0ĳ���+���������V���4�^�w2Q>��be�pâ{E�(��P��p��{�U���A��=�v>�uw���M�wFj���ʞ%:�:��=�{�2��C��3��>Y��]�� �s�����;f��7r���%}������7�^p���o�4���@SX�\x(��>�ǚ�6����TV	P{��W���ό�
�{�;i�
HNxz<�g�y��6Z�s���9�{��j_,�CY�8󋇺�IQ�
^*�>������V�Ҹ������K)�]Ñ=�~@�0��~��O�^xN��Qr���	��x}b��h�����H(�_�PƤ��EH�ˈ)������)Y�b���ա&5�`�eul5��ƶ،���bS�SB��TY+�X�,:'J�N����&9�S�z�����+U"���[l��%�T
�œL1R�Em15�`[AN5�hTZ�VDU@QB���Y�-E�!�Ƞ�Ӛ������+UU`���e�bu$Є�� �'JI�%,�Yԑ�XH	&�q�:����Ѷ�!UR�a��1�%VLnXVeU�%O>y��a4c�+��՚ۚ�㌜��-����U��*y�7N�a�kq�����
�
�4l[ׯ)1�#qק��8�,�D����n{M�
��n{q�nr脰��<���q)����q��9����!�$d���W2<</\\���ֱ�Û&�(/P����g2f	����W<��M-��E1A��g�6�
�Y�ɝ���B"�.�j#D�6�Uf:�Et�TT�������9Ԩ�sNlq�A۫��츉Q4ٕiP`���dp�Ӎ3ӪU1�[A�=[v1Н+�	*�i��\3�n���bW�X���q���
a!%�Z��Yk�m�[��U�q��0*i�B�-���'��I�sq�%0�3.���l��4�a��)����;��q��Ʋʍ�kp��p�y����;3���^��2��p���:qv^�q�����Y�\�A��g�H�X]��쁷�����' b2�Iu��>|����6�@�E���.ŚcB�*�bѻ�a��Y��b&�Q&ed˨i�;\1H��/q+�/���Ӯ�F��]qZznf�\V�h��F��Vٚ��V��Nâ�V�'ݻ6�X�}pMB�%�Y-��䪅bL(�SM)Yy��IaLC%�������m[Kݶ�C�^s�VUE�k���s-�����B���@b
k�����u���^;7�=i��6��Je�"ʆ�RcN1e��Vpu��K<��+j����8�S�-}?L��z湍�c��m�۟ {]k+55���������� ���D��ц;�j"H@���ŝһѺ�tn�rw1mRrK��p`���hD���^��V��8h<D���u��m�2rf �aͯy�`����4��$��*J�T&$����E�#26|�ɟB��G�`��o��v�HIS�ĝ<Q�jr�����R3ݓ$�(�aדՊo����� �w+0�j5�-���x�V�9'�UU��ݶ�&, ��$��[}�g{s�A�qj ��'c��Ȇh��:Ի�J�K�p^�����mޟ#jj-�g�z�ׯ��߻����������� #1st�iwϱ����$����'đw[��|��ےw3���Aޣ���n���lښ]Q���,I��w��c=3R'U�ġ6[uF�<��nE!���c�Xʰ��֨��[V�˦��L�V<F�i]Aũ҈�p[m��odii�0�⮐~#:�wS񪊄�uY �f�˥Pb&��a�Odu�W!��K�<���%�v-Lb�*w���ԥ� ��� �zq�H��x���Y���˘�Iْx]j��w��g����-"�W�#�DmfY6*q��s�=�V��A�'{�����P��Tk����hp���Za�y��&sYf�IVbݲ���&]����/8I˿u2�B&q��w̟��|����i7�.�ɥ5�W5g͙ܥ5��������}M��B���#d�5*u�W$�TS��smף��ERď^�J�zL����wsd������a��MwR�1	���D�&OE�̧�v��	���P�*��	(�v�#�*�\�"��۶ ��u,�Ոa��y��f��=�?y�N�>�t�x�&k�^0�y,���^�5�#���
���r�C�4>�������M���$�ȟ�X~ݤv�b;%�	,��J������{�����?y��}�����2ʘ��\����>{�*��~��A'j�'۰����d�z�~"v�$��С0�t���Ω1��;Q�}V��d��̭��E]�D{iI_iͺs��}���h��rwoh���n�K�����}q�� �j���J5�1܃�i�J$�vE��I��쭺s�[7��>���I=������R ���bkټ5�9�{�)7��YQY'4��a�U�����:tv�'ޱ��SU61p�#��e�M��l��	�ّ�u���
(z�����v7$u�㣎�X�=����Ç���83���k�x�lռ�u�Zyb��Y�:������j�M�6Z��\�[��'��*��$U��D�Z:8��!	�m�m��4}�(I��;�0H��A��cj��P���f�!td�m��H;4��W�&�q�p��[�\�� woyC��$\�,�	���3*�>���5�yd�Y��V}���"�D�ۃ		]l�J�	ؠH �sd��\����7{� �@��R"
aą}��'y����A�D��7�35�co;����b.(A�d�7v�8�b�ʗ7B2Tm��ϡ���NQ�v$����dA;�����,y$T�wY�6;
P��Tk��L���v�Y�0r=8W��;^�3x�{�Npb>�"�8?-�H�p��_N��UZ/sg-��3#�{��;����7�O��Ǭ;
�C0\l��%��
;V���㨛8�4Aݦ��7����_B��m� j`ظZ1+��~g���� D�3WM����W8`�h�^�4�#v�3�I���$��d� ��[�6/I�B!f�HR�(X�f�Z�����a�?3���L8��A>3���$��65E��T'�X'��&E)��p���&j��g�n�� 7�l ��7�-���C�jdN�$���l�H���HI��K6##5��)���DE_v�6k4q��z��Oc�,^������TP��D�� )��?_͒O��܊�i6�j���[[���B� ����wu2v/�&uF�>$x������Z߀���v7%�޾���ߊ+��j]��u7SĽ�x9ͷm���nʻP��=[���{�C!]�;�02U�����Um:�C����RVt���"JV�=h@��i�Dk�+h�"��I8I@΋� ��oѶ��VIz IV�f,�;Wuv��F�{�/	�p�Հ���^��3�7�/� JX��@ܔ�֊0)Vi����K��#ƾƵ?,��}TwW� y|I˄kx�8M�a@�*�]��C������m���e�?��%���c��A[kL��p<e�#W��$�2�$JM�ۚ��*a�]�SV��� ;#E�+�x��Ѓ=�dn-��%햨�o�ׂ��]ĒK�l��O�Yѻ1}�_EQ1	�[��_����0S�un� r?��_sd�E'-$�%�=��T\�,���`�'[�dO�վ�����Y�2���[͂ET E<����3�ߏ��L�Ճ�;f�b�\
��9�6u��`�q�I��}���n�g��V��*ͬ66*��� <*t�2r0;rdƝ�1�}k6��]^�%�X�I���YCM������N��+ϓ����.�\��-
�hR,��Δʕ0മ�����U�4[!�uq[��%7\���.l�ɮ��)'���E����J�']U��U��LP���v��Z����^�m���ďf�7��$vU�wx��V�U��l�Ƀ}Q��0ۚ�$+��T]r�/�?Fl^�둏����b���j!/s�D���D�J���ҳI�c`�s`.슠`�P]�a�cM��Ip������͌�-$�%:,t�aE�u�Q��D�l�g�H;Xq8�Z���`1����y{�.�W[v���B�M�Ow��'x�kET{ʊ���NF����+�V�
�Qʢ���D�'p��u���YC*�E�yY��&q���ܜ�OS�1j�a��8�� ���U|�$���{yO(r��7k�Ԏ���j7*�Nr�e��1t�O\ H'���e���i���&��R�GV�����7��;xaK�H��	�ت
a�}����>#�����9#h=%�n>>ߣ�??/�����k�85!ϲ��,,�h��r�}�~��v��_���D�Ӌ�nk�{v/ē�;��#�$�'��!tv�{!lq$:����y\�S�'ӔcfLQ'��~���
ڮ�)�v_l�H��m�q�s�]��Y*$���炵=�O���;�ݖ�a;�K��Ж߬�ڣKd!"C����##tR�$V=���Ha���n�d�6Ivݹp�!�r�Z�Ԩ�3cn+6�Y�ڝ~����Ah$)���ۭ��"iV�F��[/LdƦcgVӄظ#-��s��9g�����D��RLm��p.�8{���z� 7=���������]�zrݯ:F8���_{C[�����4�Vƿ,��Y�3��Bc}��Ǿ��Jpi�cΉ�j��냸��f�� ��߭���,�cր����:��&���0w��3���tv]'�������JT<?��{u41����r�����O�x�|��$j��P���I���ƣ�n���!�2'wm��f�a�G����Ǝ<{����T7��='|��0��;��$gg�d?_|�kՏT7��|֌\���DI"o�	�[��c�S�������~{Пi��"���b�*�lD_�
�T+ ��i�����E��kZ֬m���8��(f\AU	R��AD�X\���f0X��Ab��R騢�ȥ�י4ņ�L,�R#�Hi��X(��e���@F-�-���1�1�f"�WH��ulU�2�$���CY`�*Ⱥh�DB�aF����a��R��Db��"���-B��WT���� ��_/�W�;�K��9����6ꁩ�3O��XF�|I;���}!ٺj=��N��p�fri�}��̀Hۧ��@n�1�{D���K���C]\�5�v�@d4 �,���o���(�_��m{Ԯ��I�ǽ�M [�l�"���p���ɮSt�7@`�G_6	#v'si���]�(����� [�hB%�]���y��]Q�p�`�٫�쨹�D�i�Ol H$��٪Yv�C�n��U�c�uop�:V�K|�������t蛘霆fA��\����'ݸ���5�t�otܫ�s񧷾�>V�N6 ��'sT�+cy�Bt���N"p#t,��Z;���+����vG8i�	�`����wu?9OV�d����QL8��6"��%]�δ ���A;h+�yW���hF5-C���H$��~��{]��{����vF�Sy�UۣVH�6������!mՂ���v9������Ε�-�E]b&m�	�_�s��Y�
x:V)���FΦK�ٳa��눎Ġ`���ͼY9`��z��ME�魥k6^8����
�����]v�غ3h�P��`4��-�We��v�;�np�1�%�b��cC����cq�y.�l�x����W����i)k���읷=����A��3�+�q+k,Ptn�sa�8��
ؤ��ڸ6Wq�;��ء3�+v�YY�r6jGt(n����߃�L'U��d�s������<H"v�ĸi�	k�+':)�c�^��Fq���ےQL8�؃�^-��>��u1�ԵQ�tz�%�cj��{��t��}8(d݄�pf{�UO(���>�w,\�'�8V�FzӘ��0%	��}�c']�K�4��S{@�^��Vf;C�L'�4=gM��f�ڑ#�ڐ����^n\���Q�n�rԲ���;�)��X$�s��� /���������u��l�\�眇�k��{���ݫ�9d�e0�;�����W�®��٭S��ݹޝ�0M5MC�����ӊ;��e/s��˻S�t`=q5�ȨH(�gX9![bdή�e�h"�i�ӆ�n��hj!'&����z�l=�Urb�M�S�H	���F�@��uZ��.�Nm�F���`p�	�����aӸ.6)F�Y�Ft�	}�#n�ZԮ&���8��އ���LD#Y��Ш>9;�|pg�xx��}X����Z;-��CR��:���և�y{{n�Uv�0T��`��q>Y�g����|3�x_r��92�vrL��b���0�k!X��s	���Ѷ�v;qs)��e�8���%T+��N�Va(h����S�r�9Ս�^��K�ξ�њ68�p���h=�YUͣ�=����Y/�8i��ȍ31~º��u_wr@}�n�����b�_1�/��.C���j�R��E5a��Fy�M�]���,Y{����R�
�ۈil׃�ˋ�"�M_b��*�l^�}��5�u���\%�Y�XJP�l8m6�;}�YL8����@v�j�g�q3H6��S))Y������Cך�^���0�pf����@r��9]�]�wP�m�`��6&�.��B��f�շ�9���f�8i��f���B���oG{w��&�ܧ߶�s[�~�O�.��,��q����o���ڽ��������Җ��Gɪ��2Kt&Bٺ� |=�  �DA��������'^�p��-�36nca7r�hB���n|̶�/�wV��g6T�Z�4 �l�Ԇ��Y[�+f��י1z�؇h�e�[�ipv��ЄXh�p�c��6㋮ ��I�T�V��v�F�9��؞��Sv������Ϊk���M7���'ڇ�u{"�	���v�6�Y0YL8���:k�о���P�-V�NČ���J3o�8��(�k�ֽu{�A���$҇�r�"�K㺀ˤ��Ab���]�#��R6i�Z{da���b@vr��]´�;�};��3�M�ח�Z/"AP!��"Rm��Q7�4�}sH=�oF�������f*��8i���f�j�i�	�NJ��mBj^d��\�j(��=	`�+���p��L�SY�/*`�spl��<��{���vo�߹o�Mܺ�͹���S#z�����jȝ���^N5)-[��n &|m���׻;[Ӯ_GH\�Va��L�=G""���A� ;y/\�:3"dr���XƮ�%�uC�����Z���p��̶"���^��uc�+#�xeZ��	��9}H7 ݢ ��]�U@G;�f'��CK�g���8�چ�Lڴ ��� ߎK8+,��ܥ�r�7�)�����A�f���޸�h]�{��ʺ~O�/�I	$.�����1]ߛ?n���q��̊��|�� ��>���xc'z׈�����e%��g[B&�����WJ�#�����jf�*���=	�"�ʀ���U�X��kb�nV�מ_~D�R���� ��l�A7�����x�˄	�&��gl\q�[
�Ǫ�ajNnYQ� ��Y�`�$0�H�-��8�0.�|SM�q �����!���Z�r��r4Ѓ�6ՙ�Tۺw�f����$����=�3��:����n`s<�@�B�"2�)ĔQ31�p�'� '���Xt�UB,Ȉ�
X��/����@��qW��lt������+����A��؍��%"�SS��w�ߗ׭�3z^��W-��P�qv΁�.C,��m��O�Dpl$�㓬1&��>��9�?wE���B���g{O�*ۺ��U�/h�0�fFߎ_6A6 օ����ot\q�[W�f�4�j��Ѿ��V��_���5`��M6a�]3�;ׅ�z�2I;�$��d�o.3'p3ː��m�jl�@@��n�E,Q4v�0H$��Dfy'���M�c��0��o��kL��5�����0�bC �����*�NMjk|�u��S=�˕k��=�}޹�v��	zz�������'5�^�t�昙�J�e���W�	�O\��|"���u�����h��:H�(ӹ�f٤:����;H�5{�	E��LY�4��ʁMКѕ���D��YL��_Nseɾ�ώ��B�>ޖk���,��ϻ^�rY��
N��^^}�jȷޙ��*O!nW}3}��6�^BB����ա����n��h�=Ӷ��B�Q� �ӵ���g��zg9`���T|��\{PC�]�ս��vI�3}��@��Wg\�u�|�U�3����*������ݘ}[�X�ү�|�ָ�u�y�:	>���]��5�a�P����0�r� ����,��qi=��g��W}�(���!ݽ�I��9m���cP�q�'|�o�~|��ft����<9���w��o�ϴ:�%eߙP޳
�VЋZ�R�Qqg�X�Ld���J��Ɨ.&8�ٌ4�PU2i�m*c
�����+4�.\T�Y
̹�əI�V���̵b���QV(��q�*i0dĨi���8�
ܰ���*c�	R(i�V�Vi*�i�jQ�	N
u�RI��bR�Ȝ�.�b2Q�f-��6�bT�ə`)�r�� T����N�X�
_sO�?a���ʹ��Ue�0bb�����l�X���'����fxM�y��j�t�m�&� ����7`�w�J�/pf[����U��������*R1C^������lI��U��]v�]	P���=�C�T� !Tcmlu�8��Y0�;gZ�q�-���}f��g9�:�����f�����{a�Q�W�5�]��-Q�2d0�&���:�X�Ĥ�6�o⻎/n=��쯞��)Q���i���+E^*���v�+��pk8rS�1�ͦdn���f��)P���&�3���9^+׶�-jEa��vb Y���wO�Y.y뷣���l&.z]��;��"v �1�^w+d�q��ks8�xc\���p�NNDSu��hm݊�e0p�9�98�ݣ���YM�/����-멋\˙�^R�٭� �n.���q�:����r��_6�=�ۥ�	��G\vkz. ��:Ks����o�oZ�.�&�1��p`�#.��6�#H;�0qc�I�E���]�J���n}�J8�\ݪ��.����i�k���5UV���۵N!�5�/.��$n�3z��l[����0Kv=��6�GB�����t��H�m�.�z���.v��Pf��8��vD��Bfk��{[��r���Q��#���x�Na�i�"���y�;j��l�-�2����������OMQO���y3&N��b�8��&1IQa�%{B�]��-��.9WJ��Kqc�������,�\z2���΀�;P;�nF���<=�ZƮ�u%��e���z���>��)��A%�rs��]�Uo%Z,�lS��ǟi��>#����m��B�;W�r�BL`���P����$��c,`��>5O�B��;l�X��l����o���%_�H3�߻y"�Wn��F��pa' ��jhJ��f�L�eW+���6�5]�U��0|wu0k==J���A�����t�-���X���x-�,��_v��c����3)C-�I�y���䗗!�a�"���p;6�lb��{��
�8�a���6D��گ�(�tgR�e�
����z��	*�I�y� [��	���V<L�C��M�''�'�Ͷqc�5��A�g��}�|/7M,�$�ٺl6Tf����Z;���5UMi��6�	)�mk4�N�{dA� ���V$;!���U�K�ժ��O}�T�+�F�6 �JFk��x���f���fn�5P$^��^\���֚��U��L<?Eǎ^Q��cc���� �h@���٘�o��1q�3(��ҔwLyN�����C��)U�����&E󎑍��7qj�����y#�{�2|G�@@13��,(UGgcDf�3�2Ip$���s�:4MU�=�[����(M�7 �B��[��>u�{�C���"J��]��{�)��h�D@Q0шE4�1�(d����͢XݮU����|>�P��U�	"� �39��Xl�'{�$meXo���Sm�:��l�ݻ���W�NS@uEI����/wP�X&u�m�j��W��u��t/X�vy�~7j�\�Q/��_T�zr�u:"A�ș�a���fv����O ���ٰ�!�WAa�����"b�{{7��L�W9fѮ��8��[��{�x���B�ΣL��Mx��~���y6!M� ܺ`����q����H����؁=l!긒Z����&��S{g��MD6+#�g��	���Q�/V��A.��t.8�m�
��[&�����t\ĐI��vk�o�o��Mr��sΆ۪u���$i��9Y�Y�.6�8�w1�I��5�gY�ۧx�)��\��A�����|��י���Y�n��N�#g��G;"���d�F]�:�a�t.���(!�bkM���N��G0�+�һT�O@�6nj�P��г����b�W���F��"")
� ��=�5\/j۳��9����@=s��̽u�m��	�PjF�4G#Y�''o��%��q�d�o�.����fm�4Յ�sΞ�i�sv��Ѻ�lU�\�)!��nJ�e	�&J����d�Ke�n!zCQ��z75e�
�;:� �k�N�
ch*.�-���H�<��P�!�=�X9]���*� �Z`�t I�;t�K��h4ʅ#��3�Bݫ -�g������g|؏����t��E��5c�W��q`�"r�sм����q�y�^מbI��P5P�$��w�/7��� �s�a�|Iks��:cB��c�c˸y�^���z��\�=7N�}[��eX!��m�#���E�"�͢�0�H׸Ϗ*�(��j�Gdֹ5v�5��Wdf�P(�m�Umj���ԧvIg�r�"�ȱ����=���NO�Ϲz�>�vm����Sx�C�FMi� `�]�t)ZX ��a��o"�7
�0�:D� N�H&�X��rk"���!l�Z�SmӬ��3��z+�r��V�] �O�5��(B��� KZ�� �,�I��+�ݺ�\��ƵS>�{��	���(�H������b稚(WsgʗÇ��eN�쳹K�e�ڃ:�#f՗}H�4Z1A�
h�Lz��Mzƨ@⭭Qbܩ�������x��<U[�#�#���\�MTX�j�y��ew����|��Lȿ�%3�1
.ޗ|Uh0v�0I;r�H���4�Y�̎�w-�n*4�&M�1�rH�ߟw?i�-*Kb�Ě�Y�\�3L���mq԰�2�J
M�ۛ�҆ۇT�~���'�VF�z���v��+�-D&]�0������y{��!v���eN���2��(�K��A]����$�Mgm0H5��#J$0��(T5��%21أ�-�H'cJۺ.�Fg �E�6����'˱
����{o�&<|E;@����]���QU+/tڥw���,|!V�	��Y)���tq~�w/��tEX�9͒x�ۭ�Ƭ]��	_���*\��-���(0�L��o�\g3	�զE(�3PEU��V�-�p�V1�Jn`涮���N�Z�
T/�@�#]�{�������+�n�Ak��� <�� �W�2{D�N��w9���KI��}RW�+�߬f�|�l\��9��&Y>)�,:�b�
�{�v�����ߌ� 6�ry�a��sΎ�uW �[]����|����C�=���[��~T�ؤ���)Z�i[������/����Ӽ"�5%��鸙���=�6Ȇ���1͓m���P���.4C�M-f��R%�G5pT*�b��K�:����<|09wn>sʆW��r��(�77�iΘ.xt���\qu��--�m�����F\��!���F�+ `�h7
!6�>}�L�7�w`/�0�E�6q8�(l�$��S��)�E��հ��ˑ�ŒA��'����&��M^�
�+�&�p�}M�I��Jܮb,M�B$��^cs['ա�T�L�A�4r���]
d�V� ��l�Gt8ؓj.��0�6}��KI��z7�����ͩ�,H��~=v���`t�$�2������,�ĐZ���ǂܐ%�bʈ��r�O�?1|(S����� ��F.��M3���u��"��[
��o$a���zi[Tf�e�렬�JS�`��2�04)n�����#&6.�4�< :���ϱ�I?t"I>��	n�fpdm���5�ټ`v� ��j\Ϛ�7�$��5qh��8������x	3\����{֣��_C�8�n����V�G���kC��
O4��j� 9%ƣ6��T���h%(0(��D��v���R�	tµ__G�x�8V[���^'ĂF���sU���6�`&���C� �
wr�X}[���B��N�����ł�P�΁d��R`���q��w#�Q�J���(�
�����Z[�.�[Tn�Nd\ŋ�s�t_\qq���v���~���NЁ��<t%�<���`�{���%�My�v�2B�`{L�h���7��������ɲ,0�{���>YC�������&3�)>�<1ISs*GcF��PZgl�����;_������-B�2���um�Si�;c�\�v[<���/糺�����^A�O��=ڴ�|^������߬�OyZ�={H�,�c��x�~�͛�p��p7N�[q�w(6B�;V�W^��Y�T�������{!-l~0U���p+ě<i������3k2ED�C)%�� Х4��Z��E{;ݛ.�Qp��F���t@޲��K����b�nԞEaKHg޳7�e�V���C���H���s��+&�E��=��ް<��n}��ɹ��u��;B*�'7a��̍wo��}��YO��> �ʊ,�-���R�T1�゘�([sm�!�E�14��"�]�&j�`�9Q�lY q���!����׉h-�TmAff8VE�Aclh�8@��f�E�0�ʉejf����b̴*1���ܵD��HFi4�LAH��Kl����ȥjTr�S�i�0���!oi���d��̑@�R�1Fi1	�T֬K�e�P�8\Hۃ
֪c[��S�I�KK�Hs�t�ɉP�ō������� ���G�Ϡ">��9�q��
h�W�կ̼C3��*�	�m�Δ�:@K�Ω|pӅ_S�;ɭ������sS4�G8Z��Ԣ�a�R���x!b��궪��~w��Z�&[�3P�$�^cw[9*��%�n�g� �G*a��p$��ɞ5yj�0@�N�h=�6��+��-g%�����/�	�i�g&�^������'cO��]7w3q��9l����^*��s+"mv���3_��	��2fvq��R��kBC��ҕD�ѝdL]]D�����*u_���щMhd�4Qۑ1�谹��Ad�4BV���c~b���qX��M�]��pԢlԥnt�6��{÷N�]+�F�6���9�Pvh�S��;����*P�-�2}���ש�0>��`z�Z �;��+������~����>Ƣ��� }=R8�h�|A��N�<��}k;A�4���Є{����^��[����`�7�M�D�7u�5�ꢍ�/<�!o-Q�n���oJ�2�e���̣#6&{b��,�m�*�'�ldd��:�B>l���Yes3U��%�.���`մm/e{q���tQq�B%{kI�騛P�B
�֬;M�w]<�Nv��f �e�V�Ͱ��E��`n����:�\�۱��J6K���-��=7<���+������l�R�i�N�;pdf�jx۲�69�����q�P�p�`�\�I����ZdQ�� ��ɂX���e1�-�DƔO�F>-8m�R�a�b0�%t\r	��>7����!�7q�f�#}8J!8n�b�>����CyP{S�G�9�[���]�ۥ�Ȼu O+Ă�#٨2w5�|�\k�B�#U�P��N�Fֿ;�Uɿ^ �Ɣ	#&�35�.:�F�oH����Ӎp�����f%���he4�۱�8h-�Ɣ	�=I�A7��4��D��ϯƯT���щ5�bz"d���m+����N�&x�੘�w�Ӝn�w���㸖z��4�~�GO��;[$�����O~Z(�H���	�A�w�O��)'���o�vsl�F���յ�w�����m
N6 ,�[�F#���຦���d��NʼU����*��H΄a�ڝ8���VV�[�{G +�k��0`AE�`��O;`h\P�����'kS$��z�\��n��,�A�E��!ںn�«����k\ΰG�[F�H2���"������)���[g�Q��$�[��a�1�!̙��j�DS����6
�P��3�wuZ�;mVoR;�n��5)���|	���#��5c~a�ۈH.�FU����� �H貉$�u��<���Q�@-~lu�l�t�7����di���7��-�N�I ��U�Mn�B�p��a�{M'3#��F�.��|��|0��7���:B���YSgs[����V�R�M]^�2[��%���s�LBk���A��q˹�Հ�m����|��&I��4fi�}Q�A��6.q�Fݕ�ٽ�S�E`�m	#�7ڙ�wr^����ߝ5�W��.���\3ş�����!�9:�S��e����>���n!)�{I�g�a�8��ݼM�A5Tߍ�V����|gY�i�e��J+��&xtf��P�۶��T�N�o��,�g�0On�^6�ZFH��F�(��+��:���2}�Zh;#O㗞{<(ƪ��`�(T�^���T+imi�u�{SEB�h(n}���y�H�ӈ3�i�I���ѻW�1x�}m�m�$tj�fy͸ �h�x8��H5Z��;EթǕkWm9�f�ѴM̙W���j�w8t��j�V2����hY�;�	wU���ث�{�2�����<K-�:�l�/�,\X�ۮZ�1p�Lΰ���o�Is���LkDu�Gf����gA�7R��t=���ݎ#gVi�0m3�ԓS�����5�kf-�XHX+���o��i��S8��+����sGQj�8���-K]���_'矑����7��oǣ�*z`����s~7��=�5T4���(�v2�y�[=��w��c�DT)���bYE��bE����ľ�R��W=��#N���"�
��c�N.�?��,��PN~*KgN��uj�P ��JV����r0���m_@F�Б�Xe��󂛆�-�k2�B�6vE�U��>|�%э�m�F�>"�XVl8��;���:Q5�:C���G5�Q����f��d�X� ���}�<�d��'���~��:���cV���yH�_���������{�rw�ؗ3�>=n:�8M�s^���>$��Ȭ{4ʰ	}�z�Na�n�����p�2��(A0H$M�d��Ut� �i��!^�$��ku���rp�� I���&�X͌/��t���(�'��J -<X5`���[���<>�ϑ�$�#�4�� ��g6�v㾍!'1��v�4�EM�i��A�s�׼t�!>KhD�m�M��ֲ�`-��!�ۈjOU7��l�۲�J�hv]OBu.�O<P*2&�d�rVȥkaN�fj�A�0�, �4Ȏ'� x�v�~��7l��n�2R�F��ɒ+A��$�o���q�\fŃ�l�֬.e�p��@��ωOsi��~=6�$��a���r�ؚ���LC�vW��OV��\�X��`B����Yi4�M��@�P��^�~���'N��=n�w0�':�u��,(A&�lq��ngi��o��x�DA����u��X�V�m$��U��&�2�Un�����;Q��6Sq	�uO:��8�`�h���=���;�b�Ө[�8����f��u���F"d�ױ����2:��cR���k�������6�e7�
�(�_s,m�݃7��p�@�sXy�FN��"$A�C=�vU�\�[t+�^E���_i��z.�0O!{5�.���W=�2FƔ	l�DE"Q}�i{=z��#)�O�(�I���8/w�*�)Y;��,$�M��ҁ$t�dK�����-c�$�ti�n�sb�`i���;V�/��X��	_rdn�y\�+�}х�^�l��$73S�$i�ܝzū*�9�;���B�Q��l	R�Fv�a:�d��	s��97B݊�{��M���
�	���^{/+�3}Zӛ����/֩4�c[c6&lEYݜ���j�y��\�.Z%wK�/M�îX��=�ue����q��wp����Ў��v?lׯ6�M�����yA��#�·��>���~�;y�{&�ArƸ��,2+�0s;f�E�֒�{���7nV��x9x��(:�c�w��[��>�ܝt�<*�CT ���L�1	�F�*�XV�e�+.h���;�-��ў*t��ɉ���q�ۅ��=�,��N8}�u��^0%�5�mlT��1�tm�,$�;����b�����z�*�o�n���=IadnMh��{�`&:v�*�Y�C%�6t'� �˚o4��������J~�G^_��7��0ƏEeMvrh�����z)��l�°GH�����d�@��t�'1���!;ⴏt����C� [��jsS�d���y�r��BÑ�)���KKZѬ;B�Y+|�k\,�VڹA�`�1-.%��fR�F�3X7IX��3*�[ؘ�	��&�,d�1ׄ�aE�)b.821��]Y��b�%Յjb�bkE�i��B�ZVm����e�J�)��X�0���B���s*��+�9q���[d��Um-��e�������H�L�q��[j����V����3xu�5��ة�D̤\C*�X�V�s����X�ː����p!�us)��E��1��c\5�1l]�y��X��k��[���^~c�[�xT�-��ڶ�s��Ld�),��ZG�mj�#"]b�av����:�Ҹ͚��.����ƋbK1��K41�؆�ܗ[�f�BS�..���d.c���=Õx�\���1!k۱4;B�d�5�:��i�֎16T�wo6p�7�����k<�c���E�y輙�\3&չ�v�5;�\vy�k�%��ś!(1�16���3P-cms��sꞡ�l8��Q��!��ՖZ��(�f�X�Yu������� K4����R��M٥#uBYB�����6��#�Z=E�1�۟ �.�$�y;8�(A�*f��1Hj�ti男�.�<��ǩ�L�.���\a��>�cG\=v��vc ���nsK�jF��ɝnuK�`@�q*OOϟ>|Ls�7i�RM�#�ol.��W���նZRRV��[-uY��f+�8��uC����� Nbv�Š�\�{uG�3�'^�Hے7\g��۷-����ݻY�Ci�UlV
V⒂���vF�kH2��&�ڮ��!=�n*۴�6�n�8.�Y8����]���AƸZ]l����O^�c=X'�#��j����\�u%����Ijr6!���;E=̯m��F!����=�ٱ��#�<�a���qɹ��Ó�;]�3Gb��kyJ؝d �V ��ڋt�0��qӮ$k3\��b��x9Y�Ъ=um��s��џ!�*��W��?M�U6j�~���0 ��d�wuP��Lu�Ό(��L�l6�I]͆��݋���&�2A;��$
��M��g2Pb!PY��#k[$������&wW�5Y5讋	"�r:8�L\1�'��~��tqSZ���.J��a��ָ4�IU�6�i��Um|{��.*�Ml	��� ���]�y��CDq�$F�
�	pg]��/�)R�	E_��s�M����=��A��1 z���ר$9�$��c�r�l�ṱ4�$lԛ��P��a��2U����W2r���ҚM�R��2U�]5uV�x�f���3,��g��%\|�LA�}�~4�	PVd�ݖ�+�_�d�m��z7��A�`/N͚P������z����يd�*��a��'-?v����_]�@���l��$�M�@�GU6����2��Mj���qq�\:E�`D�jx۲�;W�5y;r�8Jn��CM4���*�"� D��l���Ǒ�+wi���Ǖ`�\6ʻS3X�H#�7۷�Y�����B+l�FP���������榗�%��(�Id�o��6nq=�<�p�A�`3��D,���0H�*q�{M���%�ˎ5�s��[_���m��%D=v�+�"H����W,Z�f�D�e �Y�������LOV��B�m��4 3�2E���L���P	鄃���%����B�l%��ӆ�n���R�����zi�G��km�;�~/���li�+�N����3m9b�R^G�-4I���Xxj�]h�Km�hl�A��"��uK�R�H�� �jgq�l��s��W&�$�u�d�7��s�x�/�O�/���|��u;�tlM�v��x�������;uU�J����Y��ψ���~fa�Q��VI����;v�}'l���J�y5S��J[ ɱ狻m�O���9-#��{�:
�LB��9�kS�uz�ӎ6iM�f��E5`�	7��&�h���d���?�B����*���؂�	y�6�C� :K�L�v�N���ʆ�mI��Gn)W�7i�}րF�\;>;�n�R�i8N\��H!��gffA�F��i�NҰH������,�����n�����ج:{�9�I��T����4��$ˍ�Xw�������EA�R�s�O[3ԋ���v��"sgrhU�c�:������ �賗<6ѝ�>
�,�P��q�jm��{Up���)s�ή�.��n{^�s��(�Ty�Y�,.��:uŖ�-�"�I<sDv�7��3��+�b]k�m�V�~��(�V~0N�I ��l�29i�ێ��v�v�=,�RɈSE�&��Om�Mv�Al�E��20S�{V	�F��.��x��f��,
����ɫ@�p��N�7�KP%�2$ǉD�!x��A��{U0HQ$!��ی�m��u�����fˠUPV����uv�b�L�E��!BA2�`�2�i�m�q�֪gټ���8O:b�$�^rd�;u�������3�Rh4�I]͈��\�Q[�fA�8Sl]���$Nk�p4��[�B���^��{1����[��Vf��xz��Iϱ�wy0|b"�D�Hzl�)D�)
�aZ�"������I$�A�{͚$Tu��$�� la�H=x�'{�څ�j!�J�j���o|�P%礿!�	n9=�锶�^����tٚEoL��N&��pX6��֍j�lt��`��Sm͋�eCl���oӼ��G�hXͽ9 �K�x��z� �e9��>7}��]�5@�Fg??w//W|��c2�i�ҏE��|I�{�gbŗ����dl��3���(A�<xge�X]ϵ ߽����g+l�/�|�Y[���{�lD��i���U=���tJ�S�[�B�lf�D���mW�nE|��&`��d�I7#�xtҸ��J��^ nڿ�^��c���JEPlo���l��37%��i�J
M&[���v���F�۶�$�@D�O�u���t1]��]�0��9���7|D�l"ϡ���z������ ���>&j��s���<��p�Nh�D�S$�۞́YqZ'z��a�q��ҏGu��`]Q ����������z.��xW���oh>'-w�g^�{�.7�������
a��Kw�=��'��1MA�Rn|��n��Nb������̓㽨V0nt��6�DA���,COДxe�V8̊������C�~�e��D�M?2I���w#\����x��LWw�i3C���m��L���H$�u���wu�/khe�\T0oGbh�h��L�"{����u����č�l��)��e:b���5��^y��$��:��:���!�K��J=�$��@�]g\��LT�I3z�٧p[o��c�~�)H4k���L>믇f��=��;���jeF��>M�Uv=�W�_/���*���6wbe��+-�%L�C;���i�v%P���*}���;�Ŝ��&��wE��rǃ2���ً	�I�M4m�mHVfku��y�Q��0������< �vŭ�Y��Z���ZԶH�m7r��Wֳ֛\���� �'ka*���U�����[�~�����k`�w`9��gd��^boXu�&I�;��^̼UJ�$���a�w��z��Mҍ�����4���;v��$U@D%��D�F�0wa�ښ0�-�=4���^�d��l�	=�$�v���n��0�S�T�i��9�D>�K�ܝ��m��� E�4*����>}w�C�B��Hf���.u�ZF�T�aZ������tv�~���Gl"=��ܤbT��`�7a5��T�A�u�p�/Q�-vṾ����.�Cg����v${֋���'g��I���"	���fo�' ��.,XI$�ދ$��L���#�̭�W>��s��5�CI��÷t�,��|�� ��L2Fn�dc;�0�Ԏ�ц�mI٥����2�2�`��Ēj�y��o���ֲ�JX�h5N.n�^G�y���ੵ�m6�!j�S�3O�� ���r��˄	Os���P$#O�]����~�����
�Wǫ���1MA�U^.��I��� �ק��}|/���ڂ��+�s<�q�d��Ww=��~��V螗��
5��L��9�mhw��8���g�x����vI��X�=��e��2�g�w���3�� ��}4�S<=;nwuv?�ۊ?%�ܺ���������$���y��?O4�yQ;O�ZcRaWk����A�*Z�Ө����TI=��I�h�;��
��A�4�o�\h�ۨ:��MLeaD�$��R�#8����{�â�-9᫗qx)����}c���b����1$�o	<{�'�8���u��V$l��N�A@���3KTv���Fm���j���ry���]f�p����0���Ay:x��E�x��=�<�;���)Sw�(��B�$� ��r��N���:�f�>>�s�~���)����%E�o��Tw+����zO?IK^M���r�����Q
w���a�R^^þ���S�~]eѶ�p����]@�_��Fz��y�ۆ]�;�	 �0D
 Ia �R�dq�PndU��U���(�E4����2��YU*[�,���,PR*y������Z�iP������&7-q+�S��N.��D5�/;�-9.�
�v�mx�1�0���f�T���9JԱ%d��Z�q#�nXZ��TU%E��M(H�Bɮ�D��΁(�
��Lš���%d.*\KTC:n��ډ���pI�1�K6;7��ΰS7�a�^蜚R��mcl� �|��۴��"%m1ۄ�m�c���dEtјe�"��Fi���1L��[��sW�*�Ϟ���܄���A$�v{�qYc n���WJ`��L�3cz�h����w0��7 4���n�'�M@�a��`����z�g7� ��Q���0�)(�1���:9���!t��m�T��)��ד�!d��JZ���r��+$g=J�i2�Q�����W$�����^� ̲��k�J���h$��AE���@�A�q�eQN�d����q!H[�grg*�h9�� �[�ow܏z�(��Ѭ�Ff����./՝C����	es��&ee����o�P���g=����Mώ}�KNG\��x�sd�� I����F�c2�Ì(L'�&�;������cnz�B�E~����'Vʭ\݌X!�j��z��7��N_F�fE�9�A�����ǝLH�EI����wQ%��1s㹒���2�Ш��$�����޸o=SP����q]8�Zut��<�X<@Ch{�?���ʝ7�{�B��@�q!PY�ω=Z��n�Q�]0�E�I5�����,*��y#��^5}�S�`WF�Yٕse���8�j���^��荞�w������$�@S@$��*BĉTV�ڲQ��;E�nD�����[��Uw`�u��N�:'R���;n�jm�2�����9��{T� 6�l�X*V8!��V�9�@����m��kU0:n:��e�Kd�CC�HFڻz����;cE�F�X�jg5U~���$��la�=T�7���Sˤ���&�pˊ!ru�Z^@p����HkVs�j����X�#3�>:�+.�i	��Á�*]��n�ʹ̑�!oh���$����l杚h(L�4*(��5�m�G$l�Gӽi�jf��X;��F�6�p�IW�̒t�&� O�kd��Lv4�O@ȦУ%z �h�aB5�)���� �@E�`��N��=� �+��[$mj��@�B��"`H)k`��L�f�҆��D��uD��=���.,mR����D�кk����Âz6.�ӕ�2��lg^8S�ˣPX�`�j��I��ϧ�Y7���b�#��'M��Sw�fՂ'y�8�N�G�3ҭ�]�M���7N�����M�` 6RD���qn5㠉{l?m��h(L�TT IuT�ICwUd�@�sW!��o{��y��]gk��l��4�n
d��,ңW*����������!h>���<���B��WK6��ꊫ�C�i?�|�}���>��z����X����XjB�{܀0<	��������xi@������e�@m:d�9� �5T�}ᴛB����z�������V!A�	��_���n�e���p�J�B�A���C�7ۺ��P8b���kz�7�C�O� �<��d�*A@�T�9�i�߇���kF]��X{�xg�[}$9i���� ������H)���rB�]�D�AB��=ʐX|���3eֱַ$�
���m����^�!����_/f�7��H)!�Ӝ���
Aj�2H(���gi��Fd\�K`����!�zm�q�Zm��㹭	����TR�x
����m
$�+
���u�؅I��^�_�6x2|��k*AH(J��M���{ֵq�����5�06�!m!׺����u��r�T����P*s��&�
��YS�}�l_ _ K_�.o>_�ˡ|��zR7������
���bd�����9/�Ė
����=7���Jp�|�AHxZw׸��a��4�S}q���:�]t���ί��H�q�����i�J+�9�m ����z������ͥ�[��@����G�5��hG�h�1OɊto�E�F�����߇�G�"���?�:3�/Z2����>�y��i �:��H.��{+|���x�S�����Y+�s!����J������V��[}Ͽt>�92M�Mc�E�k	����c��U_��/��%\/�D'��]�n!�J��YXu�2@�T
%`_s��5���Fy�|�i-9�p���
�<�2H)��>����5�tl��w*z}�/|�L�0�I�*J°�9ϙ$�B�T�s*Ad�*z��>�,�� ��[�KFI�`�=��H[H,^eH)4�S��[�9��r��6�++%e��>d6�R
a�9���V~�G��inu�
>��#��\��Ͻ'�}��|>�P�͠Q*J���ޫMH)
Zy�p�q��7�� ��[�i ��;��~��]�����i���T*J��H|;z��d� ��뚆�lB�������M2�Q��Q�|���>��}�S�mU�:����Di�F��7����D�E[������zx�=Ԃ��V��$3PXp���Ւ5�K��nEְR���面���Fa0FK���lc���:;k�4��+R�H���%�vq��S�fO(�7vWqt�=�����nmd�U���%�;,Ձ�����u�&1Q�j�hne��]��j�}{��Ϛf�x��X{�$7i
[��C��R�T���bf����ORVQ=�����IP�*az�1 ���9y��u�u������X�;Y)�k�p��'l=��CH%@�X�f$��)i�=�7�AH.k�oWF�����	*�9|��M�Ii�F�ؾJAH)�}��M��a����޼��]��I>!RQ
�D�w�ɡ����9�a6&�pֵֹpu�KF���g4�}
�^"<,D|��t��`T�,��h�����d4�\����xO�C��y�5V{�ʽ��Ku�;I�7��6��YX{߸m�@��|���zqԬ��k� ��{�ot��Xy�#��?g�C���P�2�D˄�]8�\�hAdTu�V��떾z��]z��3���*J�;��6�R��6�hT�痽���2xʐR
y�M�����Ϙ9����X{�v������T�q�x>��NU�A�Ϯv"v�/FQ3\k8+�س9�2��˓%��0��_�_H�����*KןM��͌��'�~���%H(l뾵}�#�����P��7^�G�H JAH,:�2H(J���+Ky��:k�!Ii�y�i ��2_ ]��NW,*�oR\>G�si�Nw�RVc%H)�^ᴛB������B�J�=�dߧ:��{��T��S�o	����\�5pu�K���9��i!m��\u�_=�7�����4�beJ��s!�6$�T���n$��O�Nx���]i��k��Q�D�<�c�M���A=� D>�=����$�Y++w��
� �>{q �'ξs�|;��u��u� �ݯFe������!��Ooz�����&�Vߟ5�؅ID+�
A@޾x�}�vx����χ/���h��ma�<�i!�H,�Xϒ����P��y�������~ݝ�mZ��4�o)+������6�Y�9�/p��˷�N��˼{���޼ߠ|N VR2VT��2H(n$�X���1��V��>�u\պ�P�ANo�����5�i��� ����c6�D�J���kk�!e�� B�Ϥ�U��[����O}��I��S��=���kZ�'c%�Ă�2T(����m޾g9}���m��°��5��B��VJ%��M2�VT
�>s�M���|߿>'�Qn�����Zͧ���mSi�\��G���?t�Ͻ�r�������M�Vf��m�1�������c�f$7�u{�V��v��*o�`d�+&��W�{��,;�}h��$
��o�kjAH[Oy�I �L���@T���� �#k`D�-(t ��f3���+%Nw����q�a�l���>�o�u���%��K��bAH(���i������e�њ�cXs�>h��vo��R
B��y�c�h��P*_�|�H	��A�x���~@z>��Y�N�����[�y������w�4�=��$�$nLy�v�x2燨��#�@�|#m#�����|q#Aׄ��H}Hm���Q��]��Ft�����]
iX�汁��+R
o��� �����t�S�Zt��|��y�\�Y�>ӻ)��CŹ;����d��M��^F�a��#��E�I ���=�n$�V�aOy�n$�
���s}������1 �i� �]y��m�|�����c����|�g�KM��/zzߤ�~~~|�]f?#��Ns�I�����O9�j!�J�IP��뾻���wV~�^�z�[���NЩι��6�Rs�h� T�+�z�׿&��ι�
AH)�s ��AH,9�sP�t�S��R���e���t�y��s�;Ϛܛg���RT�]a��i ���9�m ��
�R󙌗_<�W:�ɶT
�7��`y����e�h�o��Ü��#�B����~f:`V���~|�_<���9�6�@�����Cht$����Ă��k�~=
��b����%�'v`HGqM<dl���uFT`����ʉw�	'����k�x{�<F�=Ө���,i�j8�o'�I�����l�N�י�Һ���@(�����ʻ��a��T��^�ՎZ����=��K����V�;�˜��2,n;v���������uG�0�JlZ7���>����]�\n����T�z�x��TvW�9�oY�����5�UO_��L8U�7��]U�$.��)�H�ƌ��{ؒ��"�t�i������L�',�˟xz�t�Q��<������T��:9�$���e�vv�[��V�#�N{�{4$�Y�9� gs�;���ذ�|�k�#�|�k}ؕQ�u46��9�6���]>1{6�_w��{�����}��5�����j��� 1�1����Oe��x�L_0�9�|��������;���{s.�0�<��^�z�B��~���Ѿ��ˊ����v�PE�����S��kI�ca5������+35��R�`�c�DdEj)pɩ)�m�'\Jq6V��޺�JJ��d鋯XujIH�� ��	b�n��Z�J0ui!�݀]�@I���`�%�94�r��զ-��V2�CM`"�F�r���h��V� �kP�ur2'p����"���(Ԫ��+��EQm�UZ�AQT5V
EYn��"4�(����1r�b**��*,�ulTQ��Ta����"�%J*����""*�"(bEEdA�-**:����("ċ"��[�b����pp�a�����&����ً�/gq7+��RkK��ٺ�����nXJn�$M�X��u����
MdH�3p�K�-ע�f�S��ѐ�V�lc8�ۭS�f���t������Ɗ�6sYŭ���b50mJ==�� ��)[�k/I�uJN!Z79KMt���1v�"���`�]t���aR�Lt�*�ErU'����Paam�,4�ae̔��e�-��З3e�b
v�k�'�q�3��`� T�IǙ$79�r���A+5H]�Z�.ƺ���\�YB	���m�p]�5�`;��oZ�c�A�Gf�ph���`�و`�M)cG\.K��KM-��BQ�1qۮ�9���n�#��6�|�w&�����e�]�́�]��,��-{uJ´m4HM�UZk(��H��<g�޺6ɞ��+:�Y�@�ʧo"�d�GCA\�����ۧgjB���[�d���\{�&��+�6Ҽ.����k��\�m��I�bs���d�O/<���']=�'�fBz�]�g�V�/M��4b��ݹ�+�]�\TU����0������4S]HOn֮��mPpĽ��[u�kAudW�����mF�C!�ј�C�[J̡U~��_�o����bI�ضg���k<�k������(WU�8������nlYm���\y
�lc�5�>3�)=dy'g���wԘ���N���T�t�
nhK�0=.��Z�e�PK��Xײ����'-�f�c����Ά�mE���������W�鴟b7�x�
Aa�|桴�T��y�Ă�������y�w�ANw��t��Z!�|�P� �\9�w�[�����;/}f$���3�g��D�\�m ��
���|�:I� �T��c&�Y(ʁ�����i�s	�&�4�W�j��v�:k�jHui-����C�����G����ed��y�5��%B�*ay��aXP߾W�޲��v���}_ /v���� Ͻ���O��kΐ*T
����cMH)i�s ��x���/l
�7���t� T����3<f]tӦK�f3L��2T��s�6�hs�o��E �������N��*����M2�Pe@�T��!�"O���x�X���ӧ�
 V�8*8�E�71���y��
3m:���	8a?��|2�#�"�l�30*AH)��4�Y�O}u枤�9ε�蒡RV߹������3�\�P�N���w�i�l��{�����>>3w����U�E�PFD�M��p�˚z~X;�S|%��Z�+�Ua�Y[��B}��ރ�y6���G�#�`R��X�R
AO�� �A{�ꍹ���߅�H�|r�)� -���Ă��*%Nu�I��V���x���Y�>$�!RT+%K���M2�
�9�007�O7{�[�����Xo��A�G�3{�AH,�f$��SӮy�6�++%a�s�����>f��^�P�+�3haX{���an��
{�p>m������:@s�o��f�:J���k
AH)�<�4�R9�jN A�m
�Q����1�m�!5 ��#m��x���f�����������p��f$��S~��m ��+��p� ���o�t&%�4��A��S���n�&��sG�i���f�	#�����t����
�R�9��I�
�YD���$�T�;�_����f0�¤��o�oN.�[��t�N���6�c+%ea�~�P�IP �>����>=X%���>[9[���--�r�.=���+Gܽ˺��>����dsq���յ[�v��O��$�߸��j�9�t�A�8}����dY���#�X;�D=��AH)�o �AH,>s�9�t��*Ad�y��F��޷N�R
s�``o�r��5n�^���[��Ǥ���X9��W���g�����I�Js���h�����>sP� ��$�V�f0�
�:���Ӯ��%�/�6�!`5��$�sYAj�)-����ܚB!��{�ը	��VVJ���y�Ci���f � �ϻ���N��B *� dx'�A�_��(�E��%��I�X9��+(�P�}y�~��~��a�M��a��{�m'B%���d���YP9��W���m7�a:M�*�^�ѻx/�|��:��4_ _!���c�h��P*[��=��<׀m<@����O<�5�
	+���4°��ǘoN.�[��
o�`:u�}o��1���uδu�A@�X�����HR��y�s3�ggi�%��lU���ۧ�c�Y�dT��lD����a�"�$H����#�x���C{��C���p����5�ti�%��i���T*J����m��ќy�^�_�����ޡ���Y>%�eH)=��M����|/���ԡO�s��렺Ō��ʫ����_ĭ����7�t��C7}�"I��F�T�I�ٶŜr.W���X\#��A���G6����)�qh%A�ݷ�z��[!'/=+/�@��v�>��o{|4�{�s����]v��dR� N�F�s��ٸfÂH���z�e���ɶ�͓2����B���A�}��3�v�fF�ng�Ɗ}v7�bȾ�{�B���rs�9dp�ϥ^�AWbch\p��wV-[�v[j�X�R��ˠ%�]5�RI%p[��s�ª:X�K��6d��Va� �R�WZk\��p�7����	ɯ	`�q�yB. ���e+��.� ���r~����*�����)UU��c�-Jttɷb�<��ْB8�j+U�<���52�&���h)$�C�^��\kz����Kk�)���WK�fp��S���I�f����b_v�\�3�nۻUOt���$�xU��=+Q ��l{;�S�A*M�����(�����sI�5�6/(S�$���h�V\0ຣ�y2O��5u�Ыw�$��2	o@����n5��Ob���l���lt�	��{Vye�A�������Dͅdwu�U_1:3��*
m��D���æ;� ,n��'U�ffKۢẑ1r75�&p�j��p�ݎx�n}l}�y2��ۗ9\�o��ZЊnE���&,
J���^�/���w$IބKڃT�B!���!���pfG�#���j�wޓ3�]�s0���%a�I��Az�n��4�	�ϰ�V �4��R���1k�U�>�kpj��dF���r2�Ni�ᚴ�`��nձ���Ăwcixa�oZ9�\���R�N����ZjL�0�
���wV� �A9��wKK���x��5�m��_Y26e�{���Z"9����[�wI��1�*(�Ʌ��j�b�WUr�t&�*ha':�Lj�*eD(�}�����|2� ���$���L���p�^EE&Јr9��O�u�V���	���L�������]*��Sfm���fr���u:C5	�f!CI&��6��6	��rj����#��wcf�v+q귀�Yx�=+�����6	��0�7JX�4���P��5���2�=ݹZ�h;�#�&��5��o�W��Ͷ �93>))��:��� =F����������3S�<we�VmlS�i��]��g�n�k��I��;_4!S*!G��vI}�;iۊ'��ɾ�H;ЋˌsXH�9�|;��s�%� ����o�M6�{��ܒls�9:�� �_1 ��@����������k��A��cz�I��e��+ӗ�3�	ބC�/��S�7U��
�u^I�$U�� �\��̷�	'��}%Xs�%��v������_~+1� ����x
�/�����'�[Z�5�`���]_�ݧ&�`
JW��˔�õ^/ȼ'��'�U�C�%��8�*��m`ke	d��Wm�
�>�ՙx�g�5�Gx��7`�pW][�C/ldyxl���::��/Y(��5�&i���5���2��cB��+��J)���;�QQp�퇧F9�zF�JL�&�.*#s7�ma��rʂ��m"K��]DѮ72㜰��}g��U?���!s*!@��.|$���͟�Z�rv��2��}QT�lt>}��S��V�Gv�,繋�#eY����.��02�j����oʰMi��Dzfbf�$|{aI �r�Ê�0�R;�����(^>>{͂;7����IJ�Ӈ-�S�i�54�bȻ,����F\ I%�0�=��_�V\�&�2c�n�Ҝ)��Fz^=ۉ6�D��M����L%!(�	̈́	9��A�]&t�@�	u�f�4!S*!G�޹ �Q��ͻSJ��za�&й����!���.A�2�ݗNb�U4����yP��[A����>r�	���UD6�%C�c$��}2HȪ�ܮ���2��CI�wt��J�[-BlwB]٬>�y���2A>�� ��	A�R�!^/�<�8�bT7��A"���2B�ݸ)44�^�'�wB3+m�'/��q����]�;-�I�瘄d��P�p�M�lrC�i�3�i��b����.w��L�@s�����J��	�Tf`#{0��1έ��t��I��s��(T���*d�K��;��E��˕�Ս����p�I$���`�w�>&��N��`za��o	�^A�o�b:��⻏�9���)s���0�:���g���9�w��<�;m�^�/oe����E�f����FGG=�R�r����\�������^{8{�e�����I���j��h���3�ޫ�pԵ���Fx}�w��P��x:�=�N]�x�֊��a��_5���h�zk/�?����|Ƀȓ�y�� vEܵ�JW)��u���va�Kr_j��&�1�1#��e�����ٽF���3�<>gP�vuk�»�-�Ma���.
�fM4s ˼�9�R���Y�9T��/g�!�v�98�b}����b�X���j��4�X7��d�������}�z�2��9�<ݔW��b�s�M�[���<��Y{t�v��^S��2���.�����(Gp��=�|���{��uP�"gkhe9<#��C���Eb�UL��Y--J+��)MZ���CV�U��DD���Օ��PJ�Q"�F(��q�#��DX��ER*�Q�1TQ5J�"(*���V#mAUT�e�*e�Bd�e��@����d�5�0Yns"�B�eb���-TV1��Թim�kj�e¶ʬV:�Qb���b���h�Um,D�)��(9lV�U[j�(W2�Q�]j���*!l���X�$KIAm��*6���KmJ�iUX�h5�b�ڈ(х�5�E5mV�V�**
*V����ۧ1b1Ye�j��ei�;�����،y�@�5T��!)��:k��scIl�L�|H=�����'n�K�$n�[�PU2%}�&����^�ٛ��U��îU�ovb�h�!b��6�CG�O�/�89�|B�S}U�Z�1+�so�U� �wy�u��of�N�ͼ� ����a�4�}(J�T�Óy�R	'6�s`���\K�k�����mPn=G��>>�{���m�u����Oں�L�	y>��!L�WR�I�|�ﻧvMH�Z�'�ۛ���e�n���9b��c�޵���O�9{u�����>��zeCL�R>{��_O�n� ӴM�p�I�{�	�ޙ=�a�7=�-�J05�i8f������+q�f��X���m��]�;�mw� �ɯ� w�����񒕁�[[�v늚��t��2��u�����L���$��n�r����KCN�ۼ3���f J4�Ez�KP#26���L^�˼n����3*�،��R�`�I3!IK=��n�	Ͷ��W�.��!�,���WO��r�¤l��y�=*��U]-y���)����!�F�A��-��2�cUB��9
`�����y�Zf�����_Q��a+����.=�B`�2�c"ZX�p�K��hu�6*-خ0��j'��Fz��F{y��]\ћP����%���u��ʡeyK��1����26+�V�(���;T&�̳E�J��&L�9��Ĩ�r�k]
8��	���i����f����N��I;мE͡���뱉�J�[-Bo	*�|�s�m��G���#�|�y��n`�J�1*�y U�$����UL�?__l�Ot���!���\��8ȂN.�$��@�H=���.A�]�r������R�D&܆�a ��ז�ܹ3�D�h�%�F��/�U��/Y�$�q�m���[�iu�YV�W+����m��<_~�G�U���{ޙ�/w� #��@�mR�����O68S����<�JSbUD8��:2v�VR�]�n���a�5m�3�U��]��O�ޏ#�͂C95�a4::Ƹ�!Pi$ޞ�g��V��=7�$�I��V3�C
p�^_ ��ٽ9@(��$or���P͜��D��D��ZC�i��U�t��̻��� � ��A���'rv�e{_~���szIm��8bG �mɞ(�O)j��?>���j��u S<�)$�&��e{�}[�]Z O��N�C)S&!! ��$�^��.Q;�>�<���@V���շ-�`9g&�$�Jh��d������7�O��1����\�uUe�[4�l��ֽ<��_�3��?w�ӔN��jj8�Aw��f���A��c�,�\����dm0G����IR^�{�?sL3��z���0�oU�E�y�u��Y�A�&I;ۓ I�	�oqM�/p~�/���Qe/sh�8�h����\���߻應G;�׿�0A��rI�#�܌b�!��gH�م-�Cm�0�S�Q.�yQWvϤ�B#/��-O+�]�L����c�E�V��]��C����ܞ�>�JOƼ��aw�L�(��9u�3��JJ�A��qo'+�!�����e��9stԻ��&��]�/\�����!nO�軖)�!
�I&��z��t�����o93�6U�dn���'��S)��o8��,��6����I2�6�}��.ahݫ|	]�$�wy���t�r���4:�̍AÈ-5&z�-ƪ�y�2�넒I5������+�fl�=�s:�Sq�uFf$��F�9�.ԙ���� �ꐊM�����Uu��I ��^ ���;��ENT����%��viBL����6�3ow�{��3��2� ٭�	�ޙv^������ڨZIj<��G�ns=���d���-�.�z�"E܊����,��G��1Ftf����Ӑ@�(�Z���Ѕ D��ͦ�cH	�X���1��R9�����Ye
��q3�6p�!�QxGj��N��8ͷ[�KCX�Hk��f⻞�z{����n-g�X�H��T&�n9��\�Utyfz�c�f�ԧ�����Q��%a����:6�M�N��i$��݄I'*�d�/w�r�ށ�1p��Um������0��z��R.g������`�/7�IΠb媪裹��8q���Sd����L�:���B���@NɊOm^7UV���_fY :9��H|�L>�� =+֯my������r�w�*��!͘�F�Pn���i�]��$oB�
��ۂ4���P��M�	8M�6pAJB�ѹ����~yᶌo筡M� ��⳵Sh����N1VI7'�={���qn��X�D8�aVvf")�ӵF�F�OE�t�fX�����e�Ŝ|Nv��$��D�yP8�WP���#٣1[p���^����*�Z�'2��}6��H�ܟH=�3.93Ai��)����];�f` ��}���Z�s��-�Bm���g��%n�`��U� ���%�^�%Q�
V���Q5Ή麊D���2�/:�M��aKC	yd��I��$��l�K��*C��@�%Ṣ�5C�,�+_�����Ұ$���8�/���G_$
��I���z�f�����oN>���n�fa��r��t^o��yOv\��uޫp�I�jk�d��I9��zqZp�T:z�ԇ۞�+���l������(�r�꒮�v�� 2r;ޜ�X Eʴ��a�gs�zQ���h���xÀ�N��v����rUe�j[}��rQ�t�1�0N�s�j���T�`I����2�SUWk6f,�mxwJ:�|䶄}�&`G|)�L7�wK�M;�&y���1,��2���)\߳���x�*�I&��Dť<���I9��$�;�»Y�M
��3Y;�Wnbz���1⧓�ɝ��g��.���Y@�C(ڼ��S�ϻ8��(aU��A$U���A�٬ �K�`n�� %Z5M��3f�b����\��-�e�gs�-�L5�������\gi���� �f�p��Zh'y�ςE���j���	�^wJ۞���*�dH#z=[�r7M;f�C)Pb!!%�t�IV��Ί.w9ú֠������QI����vE�� UgL����7�:��	]�"�$
��I�9��&z����tb���	���ֿ��G�?�$��*}��EUPY��� H���� H����� $	�V�0Fu?�)��fa�L��@���� �Mߢo�^��|Ja��uКλ3{���$@�7B���!~��g��,�Fk�_��6%�X���� �$�$_��������u�����8�0;����DΉ�a�hC'�A���@�?�u�x'}Lᇒ���/rw�
���a�����	@�|��~�~��O��@�'rOȐ$	��'`@�?��XY0���?�u��? ������?��������?�~�s��~r����� x�!���2~���D�܆a��C$!��$:��%:�����? �M���Z�[�L�H���y�!��F2w~��������̏�$��� $	<>ݖ{o�\6��n�0?�w�B@�$A��#�XΉf6B��\�����Sr}�'��8d �$��Ht"���΃��y��������7�������?��}�7�}Ƥ�����������ߏ�u�:}?"2�	@��%����?�C�:?(�$��8o�aѠ��O�:��	�B�����~?������}d܇���O��?�}��I'�:��?���g�~`� }��FF>~����i��<<���������e�5�@ ������� �?ğ��;?Ő��-!��M|?��>�$�����P!��2N�� $� t�b �A'�Ƀ�RD?�xO�/d ! X2l��;�>����5���!�V�� {�6�$�gZC�����Ƚ��� �$�������{}�� H�����8�D>����O�S��B�>��S�C���?�i>�0~�>�>�������~���l?��g���!��}�Hx�g�J H�?I���}_����ZY$����!�� $	��v~��0��Y?���O������>�L>���w������C�M"!��C�>�&���~���������g�?�������C�|=����ϳ`� u��$��'P�����-C�?aD�C��>���0��}
w��~��Ԓ��Cp���}̂H���D��̟̘����?�>���?/��$	�'�~�}�a�4@�?Ɠ��ǩI<���ِ?L͝� �d��%�?>B�Y���]��BAά�