BZh91AY&SY��v��߀py����߰����aS�z�@  �� �� �@   �C@T  U�sb$�GFQ�Vӭ�Uj�Z���uMj��b�F�6��J�TG:`WM	
t  C�l��
4� �@   @ (       �  �ו]����t����ǆzN^�u�sW9�v�zP�}z�����f-��*�N��У�}vޛn�����k�}ݻTweOg�{z�ݷw�nݫ���P9m�V��������\v� p /b��%mc` �v�����;�F�a�;�Fۼ�s�h��z�WO��n�l;�n7`��vJ���z/�ϗ��/���<���B��R�{}� ӛr�g^� v�sQv;w+"���Gs���U�Żrksv�9��j��۝�ȪPG` z
�|{���k̻=}�}�ݍ�O�W^��V�ۻ��`������wf�]� ���%s����Kރk�@vg&����9���'��vm�uʗwsN� g��y�; �  �����w:���;Ѯ�����Wxk��(�n��s��]:W��W�pd� o(�{��qGs���u��gkw4�uܓa�T�k=��e�w;�� ��!�  ���{l����n�o�/^���V��UݷjMwn�;�ioJ� ހ�;�{c�P�vݛn�k��U����jQ���띱�@                 
��*%
 @             ��z�JH���� 2d4�  )����S�hd�� 1 L �i�)�$���0 &     ���R��Q�h��H@@�d�2H����5O
zSɀQ����=G�@���*J�1�0L��@di��o����U?_촸��I��&%ԡlKp�A�8�I�?@�z�d?5P�8����l0|�l�~s0���?��P�H%������_�c�!��+����o꟒ة+aޛz���Q��������U��z�m��i��O�����$$����Ȳ�@E�?�7�?�����<c�����,���y�L��t~�bߗ
�-�S~�~r�m(o7�e��d-Y+!T)B�V,�E�����m�t�)?e%�B�=o؝�t�Dګh��iܹ�=J�*Ҝ�ʪ��R�P���ߴB��S[�Ŋ=~1�-�M���n��1J��oU+�b�I��(�D	�-�)�z��g�&�B�IjQ�jTG+Q�P��.D1Lp!Y~jU!Z.�Rh�&��-�hZc�r'�x��-J%�X6�#�t�<�#�!d�-J��V���P��"�f8��S��B1�\{��l8�))���8��b��,PC�
�q�V�b���B��?1
�p!��?w�p!R��Zy��K�V��<k�
v\Z�B�q���q��N)5���8�+�>V��<-J��B�\\S�R���x���B��P�8���q�Ƹ�ešQ�*�R8�x���B�j�ǟ+�(�㘫dqI��m�P6�S+:#���rp��1G�z��n�"��*��b�_D����Ūn���&�������S����i�$(h�<��:"=�1�
�p |��8�4�#��+�:��	��OE1n<�U��)oC,1��qQ���w��4t��#[z�m�R�m�cb!�����V��V���h<����{�����mh�����m���q��*s۶.Ә��}����;ER9H���FU��1Ép(-��\ec�5�<��_8��v�p�Ÿ�"1Y�(�s�<�R����	q��Vk����qk(q�7L�u����g;�m�r�Ҳ��� �^�2�D��ڿ��ulW�]rk�_zl����7j�h�g���=5�{��ߣwئt�~W�Wø���+~x�p�V���><Z'��L.�y������|#y����lVZy(ZRy*�O9X'BL�Qi��QID�bbb��c]�|��ҞB���\jf(]�P�y_�4Н
�Oh]�g�i�]�Z��ض�T�W'��iυ!;jĲ��c��d��n�M�_�oX���B���{9�kS1�-z&�|6�Yy(Y#y*�o5^��.��lk�޿Qdf�gC=����٩���r8��o�p�;ü>V�k�j)��1p��cL�rz'"=�LG�	�	��CMw�Bb�
�P�#±
��w���*�{�#؄�>}��i�.]�E�B����l�B��,񭋔��SG�iI�MJ��J���d	��LX���X.X���ht�#�'MS�b��+�)�P!m	�Q�1r|'�Ք�Χ(Ciڴ���B�����
$LB�G+P���YBb�B�j�^�+�µQ�1Jd��k��b��LB�劳S���'iZ�P&!f	�O��r�!<V���!�v�D��Q�bx�U*􊐚�G+P�N!�Tu;�WM&#�u�z8���ū8Oҹ�ڔSO���	�!4!;M_�!Z�dLGrx�M<����HZ.ڈZ�bt�łն�y��jiϜ7m5"X���	���X�|���7�DiYq�iL�t�B�Q-j�]m�Ś&,!w,B�mR����=��.��Z1b�c��5�ĴB\��:D�X��LE�P6���b2�ZV�z���&.WL]OU	j|�C���Iʑ�fCڏUӥTC�o�ƞ��-5��b�T�� ~�dC�10�6��=�)X�`�T-JBܕ+lQ���G�j��J}T6!p�v��܅�P'�Z��R�IӤ[2�Q/Wj�3�(W�C�#m|�ʇ�?��Vb�ȸ�v�xC�6�f�=uI�#ֵ�D\=X��b,��m�+S&�wQn��[2!�V��=��}V�X�4��2�#b@�jG搑o�\��b�C�R���s�,U�q��^C�m
�����b����a��6,D��4c��X���gC�b�$�r��!b)Bh��!��*p���I�_� w�BC�"��F�!��Z�ZlB56-@��j%�FL16�ʂ!f�4s�B�Ä!�1��!T��47�%��\��a����C�я��+E\1
��B���|��~#&�����*�!f�Z�{��I0�b���bIG���q؄���,���~�B��:R�Kb-��a�e&��M
�7��r�s����?GU}�&�/����D�u���wX��p��w�Y(E�]]�Y�Cb-�ѹ�.\�dt1t�;Z��b�rl\���z�̇�����%�OP�>j�r-�z�R�~�[�]$;���c�ʩ��'�V<}+��I�%�2a��K���F�X�+n�D0ld?P.B�x��M1b�
�Q���\�cp�s�C�4c�O�	Q��[X���T���	��L�I�Ƿ�:�oq�F�6v�P˘fL1C���d;��S*a�P̨fl8�oC8��O+o�7��&�R�pʸf�0�p\8��!Ŧ�M���چv�5��y<�̇��aP����<���P��*���G�����ki̻Tت�S�d�O�f���}��Z��f5~{�h����O®u�[�MԳ�0�f��[sŰ�lZ�f��L�i��l�Y;�*��8���s��U)ڇݱE���]C2��Q�ۆk�C�|�{f���e�;3��\�� �M[3<�M��2!���~1��[pC�p��/q���<þgs#p��!�569p�a�.��.���<���]�1T�o��>PM�����Ч�k�
����\��=��R�b���&�!�!X8�+�q�*Q2��9��b�CoB<!j������Ǐl8�))��aN ��E<B9�!^�5J��B7�ZhCV�3�ULQ,Bϔ#|��!��%8�mA.9b'x�)�qhTc�
������ǣ�N)5���8�+�>V���%J��B�\\S�R���x���%�Zy��㕢qǏ�B���F8�H���Rk�8q�T��ϔӔk��[�O��mځ�"�B��`��������h�L=XܫES�S�ň��-�#V���+n��ʡ�aҜb9�b�J~Ա6�6��6#ǂ#ֵ������HTk��.��)���q��ξ�<�����ؑ�5�{V7h���gb-���Ƚ���b�tD�ͽX6�j��9E<V؈x��w8B�Z8�j��h�(B�v>D�D�],G��h�G6����m���q��;���8Z�y_��W�d<j�ᇎCơ�{�1�cq����Qn(�l��ofc��q����k�^�sݎ{��M�X񋻌�qF85�0d�!.o��S�}�ޯ���ޭJ�Q-ڵ��e��S�HB�y|���V8�B�f�^��s��ָƭ�iO�R��:�e5lƱ�����B݄�z�5^��3�*��9���T�����XS���O������n�������԰��X��h�O�¹YZ��z�9����)ӽ�,�a�zE��4��p5$,M+�Sٳ�ͲE��_B����";��Ի����ߙ�[zWV�v�5�	f��S��׏Zv.�I�Y[t�\����<�4���ݾֵ�����5=k>�scS���;���ޭ�j�,k,k��R�ȧ�UkL�<ľm����;�߹����n\�t�~�[>����o6�L���
<�I�P[�c>��Jõ�ʽz��[ն�Cߙ�j������RzFl��%����}&��X���m��L�v��z"5�k陨�o'}�}>J):���'�_1 �y5I�o��
���[�U�7�T&��I�,��V����~d@��&�;���yqcY���o&�.Z�$.�ރ�(׷|��j�^w�M���u���J�N ���vN=���i��Ò�"��(�%,{���ޚ��e���|�����_^ݬΥ΢�F�f�7�+������l��Yc�Q-{KȽ�׹}����H����sv=���&#ʞ��W-n)������e�$�˳����#;��yu�m�IñS�Buϯ�^���aWV��2q�.�^.���XN��|�W�9"U>�����$�y9s3�~��S*����s����mj�$��}���NU3Vg=d�͒^N�MYՙ��D����{Uʌ�]��9�{����z�E�yd\�I��浞F������aYv��s֒�=���Qs�}j&=z�/(�r������o89]���qfu%���4�>y�g5��SM�:t�����^<m��ݷ�Һc�o8m���ʋ�z�>t��7�0�}�Ϣ\GL<W�P�.�ԛHc�p۩���Pʓ�y��&�Y�͍��Iq��!kϓ_/$���S�#"lJ�<����P�a-p��ײN6����z<xۖ�<uW+W(�ѯa<��ny� ��RMERI%RZ�u�j�{{5"q�~��n\9�GZq~��gu|�k�'�Ar�}+d9ԭbkiSs�@��N�%�>���3�*2�;�-�8�ev�H(��Ѿ�����]�!^�<hc*��+�RHs��;�"V{m@ַ��^(�)���u�gS�Vm�J�+��=�Y�5���=�1���9>��`^���g3d��cؗ��9C��1w��zn��;x����n8�p���j5��[�Ipz�B����X���5�.s���h�������X�j�A�9����+4�ʯJ���qJյՙ�>Y��Y��ט�|�+�*�Q�Z��u;����L=�8����up"<����Vo^yי՜FsX�#p�)uE�͔�c�j;��.!�a��fG�)�Lz��cT-�+W\+�RbE�ƊI�]���nn}��fC�D��Ð~�3�[�eeY�I���5%�kfi�$�X��;����R�9���x��(�R�eJ�^u+>&YVgX��
���n�]j�+h��Ԩ�E��g�egk�۝AWx�V�ް�-�c�s�H̕�Z�mk�ε�\�u2����ƽ+�oi�&��z�Z��W��e}�nĞk�]�u=��ʐ~kz3�_�/>Q%IU��p��H��n��{e\1�y	�~fᛧq�uG��Q|i�����N�eI!|��cr�s��rU�v:�\���pC���W�DkK$��ֱn~�ǫ8��/va��4׺���,�W�;�1��^{�u�%fV
�S������mK�u�{7S�/����?{"!���c��&Tc�>��5ucMg���"q�Vw^ë�y�Y4��%nd�^���S3ؒ��.#�;ݣ���t�\�3̕�Y+%���<w��}c�̋�$�<��݃�,�;���a�˯�*���e8�k��5�������4(�Ql~J��Z�����j������;C���)�~Y�:�ʱ,�,�1��?\k��MC{}+O�z�9e�38F��������x���9r-X������4��L��Vq=���Hl�WRF�,��_|ϋ�ȳ˫2,�5YND�:����e{�_[����ML�$v][u���l�S�Y������&jʲ��gz�G����#qg{ ��ff��#{)�Q�9P�D5��Wf!�d9�R��Y%2J�ܫ������䯻!��gX�Y���GՉ%�]X�qĬP�77rQ��G?j�NGSQ���Υ9֭���-B��.�m�o�;��J�}�H�}짳q��s�j��~]X�G�E�qeIcIeS�ի9ƹ(.S��s��~}+Q��zy�V"v9�.���t�t���Q.:��h�"�,h��ך��q���kȵcl��Q�;øJ�(�a9I��;����uFGp���;�f5Fኣ�1�du����MGQ�j5���ԭ��[��5��e6٬jBq���+E;���j3�H�b;�oE�=�a�S��5��LS:][Q�d{��֊�~��S'��7�sG�w4�9÷s	q��N���7G1����K^��Z��8����������j��$�"��:G��/t�拑5�����wơ\�p��P��n��g��6<����1gV5��L�U�ʸZ��N��%d��Ƹ��jJ�|�S�ug`�o<�$������+S�k��jC�Y�]�ֽ^�y�x5na9M3q�qһ�[�	��q�wa�	�{�\��7�������y�dD|��x�yc��+�si���q!��(�'fJ�v�C�O|��;K�������FJ�e��gɾ�ƻĖ�J=���O�����֡�ɮ�17�ZԦd�Bk����Hͯ"�#�yX�C�*�i>G?b^�"��A��:�"Ȏy7����W!�'z���A�l��I�&ǯ<�{D�4^Tg۽���^��[����E�a���i�-.��1Fڸg�Y���.}��t�!V6�Ȝf��F���È��r�F�Ϛ�/h�Y�-}�]����h�2��Q�VY�gȨ��,�z2m&$�kMrP�� _���0�S�׸>!��Yތߞj3�,�G���;Mkb+FJ�w�'%N}a������L>�<k!x����;c�A�[�ċWi�i��:h��W�]��[cן,K7�ȱ��i5��I�����=^j�pid��ϛ����jx������|�'U���!�v�	u���JDC-aJ�=������c��~ƛFt̓���͛�L+���DMnL��O�,�������������VHg$�?g���_�uH~�	���w�Q�g�qo�&r��S���\�*��y݊:VDƩױ=;�����v��yC���'~����k�a%���2�kp�y^���ut����TUޝ�\��U��yN.�j��8k��#�z�����aaV)Z�k����I���鼾e~�W�'��ռů�;(�S��{��/���N׵-��w_]�'=��NG8��Ӝ�.ף[��R��ڍ�'f��V�Zl8�q�m6�g'�}��Rox��99��!n��QM�q.hS��(����gg}��Ժ�}�M,�/8��{��4�[��=��vo�L����{9-�n����DU�ME_b��ͩ�:O���s��vp�g_��y�^8��과������ټZve�������]���w���}&��|����ͫ�n.Ε�7�}���g�/{��I�qwЇ���s�2o�̺��Dc��d(�}zN��QOUtl�{���j��f/6���'�rg���_��WoR���=M�dI�a4o��^�*$wNr���wwKw����x׷ם��w�{�ŲBTm�r����G�}{5�z�M�$��q+{;͟�_xo�Q����Ys���.�������������s���1f~�C���M�bBI��m�n����`�s�.,�+�]�ܗM���`���fk��quTj�$M]-�Ycv��Tڪ6�l�Z���Kߑ��b�`���U�Y;"S�֑Ēm8��2�WGjL�%�cYQ#*=�D�KqL����gVd[]�m*��Gd�l�ŉJҹH��FĐ�H�ɶcC@h�_��9��EQP#�*ƭJJ�Ƥu8B)"j�<D2$��de�h�q���cbzÇ���8>"奥G�?�seQ8�Xܑ�-m'�%W(���`4dQ��Q�MV�(�k2�Q�(�j�?-EMU5�h(����=K�ں.E(d�n�s[���V"+*ʀI�TFn�G5ŕ �Vd�AQ3^qYF7��^{^���Q�Xbr�u�{F�%S2P�)Ss&�G ]�j�+I�XFMa$&u	f%-%X�&6�U��Q����qq�LkDnW�BYZ`*�x��<,U֠G\2���b�dY�Y�j��D�B̒J ��2(�=XD&����Z�\^�N"Oүo���.: ޲�*�eXQ��vex��B����"Ŵn�X!f��L`7f���$x0H�	,�܀{��9���@մf��5���IcY#ͩ�h�l�b$���*�liD	4A	4*ХxVҨh2"��/�aQ�����39����~9�8J��!�@�I|(�e�E���w0(f��gk<yV�%�#�W"&`�a��_3e����c4��$'(��>�=�jr�END�ʪQ��� �d�%�Pܙ�J��D��op�q㙟7�9���+��$�@�O�����b �hq�]�{��h��DSP�SqyD�������Ȗz�뙾�:�wUs�$8B�Ī��̗(�ح®�雤7�[�݆���J�T5ˋ�`8����9Tbf!��%�L�
�8��Ê*�#8��<�V��������'�4���
�c��~?�����8�~�>���|?�������C��"/�Q�0�$$�߫?���?O�������v  p�  @      � X X H `� I@�� 8@  @
 , D  p� 4  @$i  h@ �  �	*�N    � p� 4  B~ֳB�Ov�5�YJ�V���ej��3
�Ւem��m%F��-M��ڛSifՏPr6Vȃ-ljw�m5��s6�.           �  0 0	  Ѐ 0	  � �
 � � B4@  ,�
 , D    Ѐ�  � �  Ѐ���   h�  �   ��k�7�y	�y(i��	�&�U���V�D�0��M���l�ֶj52��3���j5�k�'��~IK^�� i� �  �` P`@        � 0   ��  �  hT�` P`@  �    �� 8@u��`  @` �@ ����SVm�q5jnY����R�oП��W}���@��P X  h@ � X �  h0  �    0 0	 ( �   �  �@    � �
 ( �`U�d� h@ �  Ѐ �
  �����n,rܩɽ�3��G�w0����ٵ(�A����2��QQ�n"����G ��ڶi
�)����F��u���Jo��������@H��G������+��)X�����A���6��m���hҟ�D)�Dq��HDFQ�#��"<��GͲ�!�B"2�ZF�DmD|�#��<��<�#��<�:�"#�:�>R"2��""<���M2��">DG��*U|�#h�6Ӎ)�F��Du�S�B"2����m%WQ�m�ڕQ�QM2�FT��Ub�8D���F�H�(�6�2��:뎢=�̡Dy�#��"<��GͲ�!�!C��x��Q�]��s�K��/�b0�ٖH=�"�P�
���KE�D6�J!WnK�%�c,��1��2LenKa^"(�q�%i�d#��dQA�M$AB�UڊK$
AX䥤JDDY1��ƫ*Bd�F���~�18ܑ��U�FX0�����R8�$�@��X��J��(�5+�*VTZ`�H�-1�D�#���#J8��[#%.X�fW%�J���N�C*��e"���'k�K�qҼHHdq:���R��Q� �R@������rh�B�����6EY[")�e,t��¢���(8Z�Y�*�� ƔUdx�JZ�-�5cn1��D2Hԕ��XJ�PpP�c��"�q2G-x±I" ��)FX	%ZM*,���
$�VT���HM!JI��6P�(�!��D�<��	:�5jE%H����LcQ�KJI����EhՑ��b���@�&J�x�Y,�E�R���&5]�CĄ㔧m�Q�N�W �R1�pp��Ѳ���F�J�@V8R D�b�Ƣ	UBK�pU��R�:<�7��k)+X�J�
�rO�]�3FHQ
cC"�Q�!c!2���bb+�R�:&B�2K��hPiJQ�hX�A���Ae��e�v�
I2"dj�0�1�J*�����H��RD�[7X�G�u�2b�(�9%!X��p����J�I�Ѕ������%H�BTLEX��"Q��u8R���aKEJ*�0R*Er��f����U;��&DU%r��pM�(�r�,�:R���
ZA��JZ
�W��@��dvdqO�8J(k�P�����Eplv�Q+q!�<B�o"!E
Zơ)YJ�Bє��H���	)Qi."��䒴2��k)f*<�p�%��VŨ0�=nH54F��$C�ho*���6"��B4��Lc�M�A���Q��D���i�4TE��V!�e��R��b�e̹F��'J�R�"��yE��UB��S[�+���e�v�A�ʐ�)�)Ih�X���K
���Z&5*�E!.,ES�,.&A���R�WP�$������cPԭ�Ye$"d�$Yq�,�$��c��K��1�ӑ�2�hrb.'
ǎ��Yqc+$C��r�F�i�2d��d���c�K1�#��y��e�V1�A��c� �#�*��������cɔb��DA�N�D�KEA�����%V&,e��cPɕB�&z8A��ܰiU�"Q��Q&1c�X��	ć�$"!R�G�M+��f��r�b�[���B��q�#�lopD�,YD[PɈ�Y)b�@�,�,P�q����6�QQbY*�$c��!�(�0��e��aD�+Q�Ld%
��,�V1��"+�D"�Q��T�+m,B�H\�X�ҎcV�����B ��LP�R��+��(\Lx2����&"��(?����Pǌ�1���P�4B���#�M��ŉziX۶4�
Ld2��Wj5
2��* �]�eH!�$ǈ��CBKB;B�EYD��q��Lh�u[PHQ�-�¢�#C#l�_M"�Ğ�������������R����B�ݒF��!h�"�B��孨�7$���ȇ!EU�!aidn�;TU֛��\n�(���)&6�hHHV�2��%b���Wlc�nإx�%"r�����r�Y%%�bL��W-U�1�6ӭ4�ʊ���-V����ɢJYR�-���Rѡ�F�+�k�+q�dI:��r¦���W�S64�Z��4��?���q����Z�:�q(�J��U��(�T!1X�ȉ`��M$��B�-k�P�*mF5jJI�vʬEm��P�V��(�j)F9�D�t�FEI(�!Z܂l�!�ZJ��Qd��IY��bJ�F�H+iF�))ia"�G�e"�;Q���t�iT�XU�F�#H�uĪ��r(�.'R�F�iXۑX����"V'Z�DVڶ&䒢�f,U��R���!ĩ�!�-#�n+�i�11K%��*&�8���R;J�VcM��t�D���R��@��%
��Q4:�V�UKI7jQ#-u&�Lv�ӉHV�m��v:�j6dN���$I�Q��,s*(�r�mpV�݅Q5�7Zz�4���$�C$Rԋ�!ZL�j��Q�D��'S$r�[RT-*��,�UF8��F��#Q�l���q�U���m&���R"Jݿ- �l؅"BP��)#m��2d�܊����2�2���T�fYk���tr:�jb�'T!Y$����Im�� �j�a-�]�k���i��+P�P��.X:��8�i[#�8�rʒT���r>�"�x֩Dڈ�i	���v�������%1�%Z�2�n'SMQ���akTn
Eh�l��SY�ȫ�ڣM;�"��dIX�j;j���cdN�, ��/�����߸  ����^���� h0 UUG|�����@� � *���{� �� z$�o{��1�KZ�����Z��Dy|��O<�\iޯ��x��(ձ����p��1DڪH��VƄ�t�6**+�8�UT��T%F[�� X��)D�+m�P+jT4�*��X��F�D��Ĉ8���E1J��;����JTT��x�R�E��P�
1��M*&X��AB��L%+ �k1ђ�D�W!(�!H�eT"e��40D����m��K�.9� �\��*1ܤyY%C���)���\e^F!!�YQ��F8��AT�h�JQN��af%�D��#c$n�E+!,(�!�؄Q�V4�D�Q�hŐP�:�	0��D�`�R"H+�X>����z�+ FQ��tj�ЫT��p��I"��Y ��(�P���-N�"���R+T�F��*�h�+#�$�UUQX+Sj�E��I8�R`��V��r$Li�u
�	��̶b-��c��R9����ʡDK�\���kCc�R�Gq49U
+[�Id�:�%cVD��[I-������t��ϯY��{���i�oiBq���:�}�k���ij)YKɼx�v��%�����}õx�i��y+׹wy{W{7���.Ů���j[�_����:i�I���ӈ���9?���ѳ���0RT�T�����g�a����� �q��$�޼�:���Bj9w:i�����@Q�P䎜�41���aI�y�)p8a�88H���r�HL���Q �oG�p˿�$9���J�=P�����8a�,�Oͼ��"#��8�2��uƛ��]��c|`�+qh��u��ӲI$��=088n<1�1��LIʻ]%x�����ɖLs���7%�Ԗ}�$�wK�X�[0�x�f�	� N�WaeX5ey�Y�ڽ&�jce���>^6���D����M�u3����H颫3�K���lܟ!�C����@�9�����;��c<uO�i֖�-DG�:x���t�,ɍdj���DTa��-�Pj̢T٩$�""���rB:�:A	=~��ʌ�&%�O�Zc��.�i��tk�$!)�ʸ�GFhÓ#��0Auf������g��ᧆ�XLuN�����S��?����$2���0��<h�p��C�"���rA#�޵���s8PA�4���B��ے���ό�����ˎ�~n�Z��U�aF�S���N6���DyGF^yN�Ӿ�r�r�)M3�	����k/1;7d���I#� 3�M���ep���Q���]Q�>̩�lߨ�Nn�D��t�`�J�����g�ף�4�Pb&0૓f@yM˚w7G��bz}�w�*��a%J�և���)���Oƚ�޼h��KRf܄֨�X�p��c��i����i�-ƞiD[����O8xN�!�e�����Eu&l��
p��.M|�T�7���˺.Q.ueQX^.u9h㉲7ҫ�[��$QօĒI;���_G�Gr{�/,�P'G=�Ւ�TSS�-W*�a8�uj�m骖W'�)�[�,�
�ȕ��O�R�!5J������G�E)R� �!�l�k~�}��2b��5t��0�Gڗ���x�%�j����xG�lx�HD,h�ۃr�A8l�^�s �{i,�ʔ6�D�H���jVL,>M�
։­���Ow9P����ܐ��p,�:NBcI"D�RJ:<t�6�u��!3�5�֭��t>:����Ô�C��!	$p06ƞ���0\I�M���Y?�MaM��CU�����#��u����5�.B�с�I�.g#!��Jm֟4���8��#����������IlD���>�$�FǕ�Xh��Y!pv0��6G�QJ8��,%�36��t�E��_��x�����wΏqT�L���W7&�CGyLY�ð��N�J)P&��.����1���89��GJ!� X� vM��/�L8E���`v�Oh�ͭh�"<�#���yN��Z8��V����1׀�F�ĒI�F��x�A�Ӫ�<~�C�|$!�$f���:�S	 ���4	J��+�� Gh9��8X����ee4S���׼l�oUy~�x#�/C����\:��3C�8[��L��Y�1qEH�M�)��44��z�������(��N�af��M�P[�*M�ǘ��2����8�ַ�yu��uƙ��v�[T��|����y!��o��=$�C����� ��8�m�ղ��]+�`{��nI��cu�j�#Wš����T���1�c4�i�74��K�9L��@������$x�>����R[9*�l��9]��EH�Y[�X�Q�������t�uT�'��S�䑓��H6PT�����O1!��ਝ�l7Z��E�lçODG��u<�q�j�3�)[ѠK.�(�jZ�\�.���tC���2�q>4�a"�v�ku%NN�i��k2|�+�
��m�Oai���cƜF��Zm�}��8}�����D}ax���,5}�c4���{�v��[i����X�J�b��VvD�4c���D���g���ᴜn�gnMG$���yY����q��˝��ܗ�J�]�.4�,����m�����2t:p�G-�!XSRHI-�����N^4dr1�$�k�H@�>�NU$d^��F\;8g��ĐR����y("��L�1��w�2��g ��=�����O	b3�W�w�:����Z8㔮\�vֹ#`���h��HIp ��MҚm�y��8��#��<y�8B������OK��H$�Hl;ZL*`%"�>�0�RB�Y��$���_l��u��ǣNGCz��\�j(�T3D�x������)�N�Ą!�n�,�ߊU2�R����%�_���[6�'��ȳ����Q��_f��$�������wRK3��:e:!��p^�ӏ�� ���s��$�m�t���x5�ˢI��Nz�ߪ��<�Z���2��O���L�mL���m�mKU�5�ڵZ�l�ճKf�m3k�U��f����j�eof���qO���f���-J^j���x[�/+OŸ�O��L��q���S�Z�[+S����>U�岊��f�h�֬�Z�h��j���V��+���5�Z�V�6�m�mK&+�_�g*���_�e�4���mV�U�Wj�-�qV���qV��[?�g���Z��;S*�W�~R�U����U�ͪ��f�e���U��-�U�ͪך���O����#�>�f�3������x�j�u\^"���s��%��I�I�Osx�.���x��u���yl���v��1QQ��u�mV��x���[6����y���ٵ<��Z��V����ql�O��U�<姊yʖ�K�xO��KxF�a� BƏ�9Tk��g������̪�Ϸk��!����������q���ꋧ9?R�{hyi���B�~G]va�Ɇx���;Ǧ'���i�l��O�~}�%��Oq�u��R:�3h�!{�v��z�ЧZ��R����V?Vb�f�E�3S��L��ytmr�?M���~�����巅�K}��^Ω�|��r9^�m�m5�״ܶ����L��~$�O����J��������}�����?���.�www}��kZԿg8c�]�}��}�A��}��w��fd��������� ���_}��3?}�{��]��}�3$�]��wzֵ~�a��<��i�m��DyGQ��F^i�1��	�EEEhH*wŧl���wR86B0N-�p?</>�����p�l�Y��:��� ��~��h�j9rzo=�]7��YFHd�d��*��.aq-���,`�lW,]A���Y��X�#c�J���a.[b2������t��@4�CCLA8pr��^zH�넢'���,3ϋ<0i�ш/����`� ` �^�҉�,$!
� �&��p����[��]� � �:?
�*x��4>��A�@�Ѷ	�(�CQZ�G�4��┨Y�,�����y�^u�C�F^i���O��v]oQQZj�BU�dɚ^�CM��#p�c �ZR�tk�0\�6@����$���f�=Ĕ&'��B3x���Hm�!G���4@��cX��ÊNV�1�>��{J�9��3�2�������&K�@QD�����'
���=��\��i������U`M P�5�\�n���k�oe	�/Ñ�O�D�����ҍw�)��Q0.NO������ָ��mD|���h�UX��ѲG�ad�mH��im����<��������� иv���d�O���͙�չ��K�E�����[\s�h��9ȥvQ�]���WK[�9�y�c��{�\:h��db�Fھ\�Y׈u)¥5�w�br�w+v�i�p���ɜ��$�:X�dR�T�����w{4����X�.�_D���3�Z��؛���]M�.��#2��GG9��N��eo8�9o�7��:�'Ŕ�CٺZf���y
���O�Aq0�M4rE��B��DDy�T�� �!�4@ʁ#��&	)� ���SL4� ѡ��X����=d���gd�&��77�GD����M�����4~R%�r-�5��`p�W��׵�4A�-b>!�Q��C� ���F^�d��������$��L�r���r1���>���:���gs�l�ɖ�HIC*�� h��GuD�4i�r0Q��i�X�96���Z:Z'sݳ�GQ�;h&�MBz�tv���}	������Қ�C�u柚u��?8��#��<y����s��Vq����\7X�c|8�;WhՍh���f�P��c,|QJc��5t�u�6�� �h����C� ���\s��:o�ۇ�6�)�oi�;�UV`d�5�y�S �7s���||�o���H��A ��C�������h�Cl@o⋃n�K�By�� QP� Mz��D����p˼(�p�&�w��ކpB1�&��Zb��OP�0�Q�0J��`8��2@/2B4k�`Q#��:����~槳�~��)Oi����#3�.�$W^�M�A"����8����G�6��i����ߜDG��x��[β�.��y�j�}f�Bl���QQPHԄ�������:!�Q�4��1��o����tt�Y2Gvέ�ڍL�8��q��9���'��9���t�xcXq��E�J���� ĸC×e�0	�)������ƴQ)*�)�j(H�N��I�~4��o��"ǃ@\
 k�:�sp$��(����*�G�0QX��)��L�D0��/���Kr��&!��!d* {�C� HXCM�!�)�q��d��]m
8��&3M�@�!X$v%����5m�D,�ݬ�Q95V���p8�i�4��O���8��"#����?��2¬�xE�GD�4�*��7���f����KaD:(���44��ۣ4q3��n����ݐ說J�(7V&�L ]x�,b��g妎r�|n�83\�4�.�9�L�Zy��{onr�ن!�E.���*�5Uh� |:L!#NT���  �)�@�.V��|�k�
��O�j�i�`d�Xm�d�Y�cM45vx�H+u R@� J�a!��#DB����h��[sY��"&�u9g,����ȍ�J���B�.��ʰ�G���XtA���҆Q���m��
`�C�40�40�im-o���DG��x��p��9��ql���:CS@��<�_.CN�᣼V񜏛�&ʷ3���k���K�{���Ğ��/I|;�TTT{���r���˟��y�7HH����޳�"z-|��%t�O��\޿�t�-3��wa�Hxe����j�8(.����=Hphg>�U�̛��٦��\W�ջI�)�E�~�5'���8R�ٻ�7���������P�tc�2����l v�|�C��m�@�2!�T7]�cC�l(n$�DS�O���1#M-#� �IT��0�%�IL�6t�	c�x�Ic���,ǰ|��0b�q$C��:A/�O��®���%����.��{S�(�9W$�P�87E4l�ٿ�h�SF�	Dz	\�	�r�P�%p���P����EA4@� ��84SM�!u�Z_!�Fjh�V�HO���cVV�M3ٺ<m猠{�pGqp4Ѧ/4�����Ò8
�n�0SL^2}�U1Jp��yƞi�??8��"#�����Qw������.�:#No7�[=�u����***	 ��{	��Շ겴RB���� �l$)�Ħ1�\6�M�<���|�ٗe�ܡ˔<3V�ٳ�t:^	�OG!���f��u��d:d�~�Ѧ�����ˠ������#�����#4ǟ�4��s���+S"NT�?���,^'��l�Y��r����5yђ����� C�%��=����> =)Ԭ��!	U�B�a�A���kE��aa�.t�i�@�@��s����u����%�MX^�l�O�6Yoϟ��DG��x��un����D�W*K2ғX4�s��1QV0��y����0ִ<�h<}�ͷ�L&�~����7BBÔ����l�iCoR��2�Ci����S<����(,l�$n`l+Ēo^ܕ˺�3g
�Ԇ:wr0��w\k�c(k9_�
ɔ�D�Ce���)�1�
C�:0&���7C�l���m�{ύ�``���:$�(�x�7YUuxRR%5�ډMUZ�Q �^N8m�9l��9p��~$F
$�DL��nb���5n�m�h�X-�kXc�o}�U`�q�x�<[����<�O4��o�"#Ȉ�<y�:�E��3�� �˘�ɔ��ޑb�9�Wo��c�0����i����Hpx9z>r�d@�릩��6�c��{���������"����4o&=�������䁒0�h2X�aX�k_I�	&���@6�i�e5cC�ܰM�9��a~��O�I8692a��[o���P�Jqd�mӆǆ���M��K P��c6:0���������"Q��6@:���?4�$07�ۋ"�A�-�:�n��RYC�?��"�V<���6�_?2�M��Sj���bٵ[Y�fך�V�6�6���Yf�Kf�m/Uhի�3jZf��j�eŲ��ⱵiV�U��UU���j��YKU)j�-KS*�c�ږ�8��il��Z�-���VqjuQQ^[(���R�eee�EE-QV��mQjf+��[4�U��[V�q�U�ԵE[��KU�Km���Z�[^j�V�*Ե-�-][8�[w5l��qV��ڼ���Z�l��g�o�?+�"5�_�f*�g*���Z�Z[6�q�[6��U�[.��U�V��̶�q�Z��i���`�R><dɆ�%�!$�D'��I��'�����oI���V-��uV�yo�|�_*7����F|�6�TU��e�U-�U��T[YWͪ�5V�U�ѕ�ˋg�|�)j^�W����x���yPc���F���'㣓�s�g6��ѯ=:�F�MQ�un�voW{v�>>�������\�k���s�a�>/'3nj|���:�WE�<�;a�f!�Ӛ;��{��ɮO)|��ޱ�O�϶7����*�!s�ڛ�6%6�7oO�i��Tt�=�&髗��p��.t������ʹ�ͩ��t�]Lߞt�5��s/-��9���qF,S;~۷>X]:���r.��I�����3����-�'�NcIX�O&�SNߏ��zp�]�d:�����̍�빨�Ξ�6nf5b�-���+��)�b���{�Ӻ�z���fqѹ��g��^�}��Roq���ۗ��S.K���x�'�e�N������w����w1����1��#�ƚ���'ej܍Q[mJ(�CA鶷��H�4VY�2F��M1�k����&ґU\���L��t��[Q��k�a����4���O�� � �����L���wwuww�X�>�멟�{�������$ 0]U}~����ﾰ	 �U__�\�y�<�O4�ϖ���":�<#���N��D;"T4njpM�I�홦��2�liQ	;$N�EK!-U�22�*AY"�b�Ak(����Ұp�����J$I`;1	��TA�Liڲ!�d+�PT�����)pL��
"4"�P�L�
��kCͬ����#���)l�)Mb&i�X���HHc�x�+�W4�,N�(n�EdzA��d��:E(�򐌢r���Up,+��W�7KJ�!".m6����b)*�J1TQ&(Ȧ���oXB	�d�ۄ��L��mA��n��Y�h�e#cf,A�\�岃��jD`�I�i=)EP�Zܣ,�����q�-��ּ��+�l�IXݲ��JD7jmT���4�e����$��w$�GGl�	W�R�RI*ڤ�n�l����P�ȥ�K"���6���WtL��������/e����:Ԋ�9+�ئ�i+M�r
"���j5~Ļ�1��/�n��o���zs�7ioB=Ss��TB4"x���NuD�s�������������t��NJ�ZS2�лur�6��b�Z�R�+U)��mܛ!��0I;�Q��˔>̦욚n���O-��'2ǯ�m,��i_77��2���W�9�QjM�����x����qD!ƃ���\�p6�~�k9��W8u�;�QXQ�#�ʚ)������:C�A�(`�l��M��(�������v���^�<. gL���C��
(��m���|I<A202@(���ac�a������~l�$����$�?B5�	;�aL��v`2@��ɛ�4���x���,�g�%Xc׿b�/��&���8!�U��G�_�9F`ș`�c�w�xي��D�!O�OB����	���Z-K%�ixp���y�S��M�J2Qki���>~[�DyG�<��<z���-el�e�=�2�@�@��P�]��_�F:��Y,���8�X�7ͱ�`ʍ(NM���EJ���
�4[�Z��J2�&���;�\�>`}��w�����M=
B��v4�H��Yb��vOP��e§�$�y�g4�A
6q �G~2�.a�ǘ�g���rDE��4�2'j�j��BW�,�M@8A�8\��8p2X":Ԍ�6@��0���h�<��.�h��)�~�
e�M=w���G%�|4|6:�}�I)����5�h)�,�e����[���"#�����S*���*e��2K�����蘪2��Hi��c�@�P6�݉��d,��n6h�g�
�,�CYl�t�C�)�e��	�.|4�`B#�e93����m��cdi���Q���.�щ�+*�G�C�Ȳ���ミO�I���Ӈ�Υ�ʹtax�7@l*��j��s�9��26k�J�Zp�B"K�ܻphB�v�~���S��5�:4�,� �p���$�l�c�@��8��QDG���=;pqms}�Jt���Q��;�40�|#Pp@�!0ȍ�a�4į�%�M��		�T~�R���"��6C�u��a���e�w
n*5���]ƍ�Q�s���<�̙m�om�e�S5�#4D3L�!x�O�:��o�-�Du<�qg���.�#%9���1�`$�?-�l��0�O��J d �08(t�װB�#LFdF������d"Q�[�ݜ��h�-�MoM��y��"�8!萄��9��BHe��2A,ǘ5��cP����v�/�C�f4�I��6��� ��l�Y�OxG�7CE�)����)�C�d$V��Q$W��W��Y
�"!�
��VӤI��A�Zt0`ql�B:(t0�<�Be��rH0���!],84� A��c�3��1�� )��`B0�i��mm">~~qh�"#���t��!/�|�6��n��9��>�N��9ZH��YWS���j:���r�*�"����}�j&�i�� �SNp�C�?=:.�7��D�w�-�ͺv-<���o?�8w��Â��68{N�/�NrI�ݾ�@�x�C��=t�biʔ�i�\�����t�m�Y_f����U��%D�ne:�&^SV�U���6+���Tz3���~�>�ׅ������7l�=�A�`g��f+G�^��k4B"�@�`e�ˏ��U��0@<=hp��a��FF���`B�D$;�#Aa��`aYFRh�,C���#}\+G&��M6RX��'a&�N�g��ju)�s���n�;}#���!Dvv�#
�CY5ѷ	 h�B�HgrG�%J�艦�p�ZE��Zp�>~��>g�8ub!c
6SP,��CT��!t��s��
!h�R���Ǯ��=���8�����aQ��Ô[ t"@�l���Ě��.�InLa�4E���ͼ��|���yG�<�\Y�W�4������휳<��.1�c	
7��<a٢~ pFq<� >�?���Ĝ
qe�YƔ>�W,۬��kQ�֝#�TT�K1�~2��p������D���gV�TY���X���C�Pi�F"�%��H��m[
|p�/M��_1R�>~�������!���3�ێq��z[��n�:A7����ayc��o��ur�,������̹����S�_6>���G(Ƌ�� �B�e�ҡ�&O�!��M�PB�db`��A���8��<\�d� AOc2�HA�)0۪u���k[����yG�����Ǟ��l��BoTM4�N0 ���"-�m��lCeZ����+T��X�Q��tg����WFm,x_���+� ������44x���n>#��x29 �G���F~�?<)����Zp�X(a����IRۗh�ht���\)3�荒��gC�D�(vF周>�v�� q�Y!!I�?>���W�S棴�	��*�rH����.�B��6q���B97�*����fH&G{��Ά�` L?b��
^��ꉋ�v�83�D�Vw�h���s��L���7�p�&agG#�� Y �`�Gfl~j�ђϽ$!!0�{{�.��)u�m�[�Z<����Ǆt�R~[ǖ���!��Z�XHf�w{��c�0IR���?���%:!خ��P��H4�I=�'��9�5�pA��j|MD2�M�+>�/K�C!w��u��������2��'a,��4Ah ��)�^�2�t�s�å�pF �2j�RQg�UI�d�
u�ǣƀ�T����P�}�<O�\1�����H�[U	TX%$�M�~�U0:Q�T�:0-�j�G
y��v�t�5��rgH��!��K�C�Y�V��u�]�#D�&�z6��pnҡ���cX�Ҵ�F�R6�oͣ�����yG�<�V�>��ֳ7_�W�8pۭ8��b��۽헣㛐��kɮ(�{7�L#��1��]�P��Ie�J�J&�i�� �p��򧿾��d='_�c5��i���=�7G�Z�{�ۧ!��n�d�\S����&0�����g9�`�v&�+V�<�f�ԯ�ܽ�B2�dڎ*
X�:�1s\�΋����.�(�j�3<��ɇ��x᤺�Z��"��O�E�Uh�#flcY(���T?0�̌��怲��k��p|���o��>�qg�|#�g|�۶v����;�8�v�kn��<A� ���j�9/���)!}�uL���Z7
7PW��ē��� ���TB�'�0���>���3��&0��t�[�� g0W�bd��8��l͔?��
0rK͔#Ih|��4�H��n���� ����Ϲy«��ɴN%tYeYwtJ�>	��|A�4|A�A�2'X��ӆ[3�cwB �C�L�H�ʊ!�3�Uhlӊy�m��[����yG�<�V�+m�X3L/ZkU��"1����BFd[M4�M4F�«,:��������m�1��N�>Z�uL���v�I'���Cp��r[�:�C�a������u�{Y���7��x�
�մ?h�I���7��aSc��p��@^��C��n��L��zm���!Æ�w����%]��3���6���>!�v@�ԡ�����C������41]:���U��»H��ӎ��c)k�5E����p�G�pşbǀC�vGdA��}&�e�C��4>�F��3�鿍� �rP�6fQ�!�!�.�2�y�b&�nGP0@�!ci�fu2���PaA-cy�>!��88g#/���m_�ڳUl�ٵ[Y�^�ٵ[�ڭR��5L�j��k�imZ�\[6�L���3j�e~V\u�'i��W���[�'��|8ͪ��R�ʭN)�-�q���>U��ejZ�����c�f�ʢ���ѕ�6���-����*-�TZ5�m�~[4���Ζϕn3j�Z�QK�J�Z��6�m�Rյ��Z��6����U�W�-N���qn3�uV�+��y��Uj��g�gkf�j�-m�QV����gKfյ[�?����*�j���_��[9��U��m�wUl��SWU�*�gj��-�;N��%��4�R{Rx��*�jʭKV��j�V�Z��+V-�V�8���o5k�[6��?��3V���ԥ�k�imZ�\[6�L���U���>����V�x���R�U�T�)o	◊O��ڗIRK?���^�Ü\O�����D�7�����ZD���:�y#�N�΋�o��s!�N]My붣*v&"T.P�y8��P�ĺ��F��w39�3b�[�껵}�|]�*����+7|�ǖ:Q��8�+��U{;iĻ�����$�u0G��Ήۼ���˪ދ�������yH��Nr%:�n��'�W/�ט���.�����=���٤�<h��B�7���I���ߟ~P�몯�������� P`@W�U�.������ ( � +������}�}@ }u_R�%˓\�r�ʗ.V�V�֏"#�����ꭳY�u��c�hHl���˦SHˏ�dv(���<4x����P �h�1He%w�3N�b?��
2d=��L�3��)�4X@����oF��wV�Hn���L\?��Q�EJ�����k�o�1�N!��x�yv��2�db2����#�O"th���`��$���&��v7;�[��ȵ��!��[���7����e�!����
�v�s�=w�i�}v<!�ࠢy#6E^�c$"Zw`N,�>�L��|1<F�0���4����Ϥ˟^�(���R`p������iJeju���mh�ߜZ��Du<�Z�~�3�j�K��5��\ʓ{�TTV����))JM��4G�.U����x�D���b�!�����p�aD^*;1,n)H��h�D��xi�Kf��Z�fs�d�6d�a����<d>�����f�>�P��h�'4�>�Iw3Dr@������4m2Ro��Љ
s���Q �#����F���g�@B;�Y��p��$�9Ì��K�g3^�a��%cd��lpB��c�͡k�͚!��	HO�����m��u��tp8��:�UO4R��R���U�b�֘�1ǘ�~�>)��<�M�o?8��-kyG�<�V�;K�9�w[/*���s������0�G�jy-��O9�.�쳾��%n�nNv�j:�	z�q�9����cV��Ϸ���~����~�Ӯ��Ky���W��KX��K�B����)��;C��OgIʹ/�.�*<A��	
�8��wz��w�oqF%<���ߋ���t���j����[Z��z"D�	Wu,�y�����g���#Y���|8&�ڡ�@��k�K��!�Γ����FƸ��Y�OA���ǘ��!o^l~7a���*��e�T�E�h�U��h`�>���à��q��ٝ�D.�8�rW0���H<p9�l����r�$���K�Á����2?@��E�h�¿"S�°���L&eRB$?8�Yv8��U%�,CI�,-Yӆg��̆�������$���O�vK���h���qa���(񦑧��[�Z�h��ǞS���'�n���@$��\�**+B@?s�
��%@��Z>��B48�WR�:=d�q�h�[������~��!�j��X"�"����G-]��C��Ą!gOV�{���C�Jt��i�B��T��M!ԧ{�a�H� �~��l�뜪H~�B��D��p���xtX�gr�`tl�f�ڄBH�Cp�:r^0�0e��5���q�p�3.��`�}����޵&�Bp����I)<lż)�l��o�:��-�庵��t��x�����?bIBC�J\�lR���Էw�TTV��9�V-�QEP9ٿ��G^��Ӄ�نwą�d6G�x����M7Ph4C@4�
�8yI�ǋ�|�NW��O����i��6��9�p�#}��o�_3�m�]'f^�wZ�;�N.W܏�f��ɝ���^����2nx������60�}~tp�4Bv;�r1��T��9*FtB��8�y��O�Op�8x�9_�v[%7q�g���Ύ]S���
!�k�W&7�``p�Fj�B�2Q�E�,�Ə:����<y�:���1�c:d�>�QQZ+��4}�?=.Z9!��p���ن��h�!/Ñ�@��Y<x��R`���!���.���e�D��`��{�1�}L��"�x�7�q�rLw$>ly���'O�����rW߿*E�2�r�����&!���8$6l�������(2C�lm�cp7�#������[!�9cf�A��@�e2�L���ӫu�庵��:|x<xGJU��v�R�ꅥ�z�v�f�n�w~��w�FE$���e��+����**+BC^��}�n��s�N���P��֨�Q��J�G�A3մ�M��z�[�T�5O��)��GM�;>Oq��G�KD�Zv*�|�b�Zޅ�������lUS�яȾ�tT��=���|���/U�{��ض�y¬�G�RSS״�8��<�2�C$"�t���d�H�`��ݾ d��0C����!�*9	N��;s͍�4͹�#|�7Ij,y#�����=p!��pb���|gJ�@B9Đ��H/��5?D�l��zt4C���c��h���nT`�RT*�O B�1�'������eZiaGm�6�A&A[y�嫆���4�m�V>c��Ҳ�\gd�M2��ki�u�~ukZ-h�<y�:�>�cU��e�oY��G>p���Ã�Ɓ�d�Y�c�|����$>���d#z�M�?l���'���J�L
!�t8!a��3߀��ҙ�❊�ǊS++Yi�{��b*��U�M�UT�UV��T�>�Ƙ�H~ C���:#g[e�<e#���'�/+#���s#��?wW����;��K!�r]68J4ph��?���x\24C��{�M�P��u�y2u�L�il���??:��|x��Ӥ8q�au"_͢���$!�$���S���Ѻ�Y������(S8d1r.!����T�&��`lv:
!�<�'��l�!��ߙy���l���\�B?�٥F��M����`��`
!Ĩ�8{�D�vn�%h4MI��Տ�G�>8pɁ��4l�p��20r:"N¡.��q��(2k���TP�0�^��d�BU�	C��<����a��ɕ;�4Ř����>4m�:�ͭ�����խh���N���YR�#>UY��}s��{ǐ{1,u��Ԗ���؊��А�]B��i��l�20������*w�x��˕J������HW��$q��3��Ȏ/F:|eJ��4�����<l,���Ӵ��<� ��Ӗ�)��JS]+
ێ�W�|��q�{�/K�.��]`�Ҹ>�~������
!��^��F� Q���a���4't��Kv!�,l��w���0R�Q l��m��|�)��|��f��Y��U��m^�6ժ�o3k�y���U�J����m�6�U����E����gڬ۹���K���y�x��'�U���Z�j]V�n�l�W̛�ej|�R�g����:�q峏*�J�Z2��Z2�E-Ql�KT[8�fћF|�<�ʳ�یښ�g�[�ڭlڼ�*�JZ��MZ��--�V��Z��1V��R)ų�W*����q�m]W��l�*Z��Z�mlڭV�|�VTU�g+f�U�U�����[][+W�Q�R-�F\��m\�>�BY�O�f�3��ӧ�%��x����I�R��x���x��2O�6`�<xp���a<_�/��x�><?������W�~e�U��|��j�W��T[+^j��Wڬ�Ul��*V�e,����T�I�o�Rx�$�q'@�& �/����5~fږ���{��}���񇕷�}���}��Cv��;��R�@:U�m�NT��T�U���F(�ݷܠ:�:˩
����MꝌqw
�1�u�.�4��^򽋝����5����8)�Gן=��K���9ݲ������<W~�e��%�;��:E]��$�S�\�i���S��8]���F�tf�t�B�u{������}��|��3K�X�r"ek׵��[�ɚ�Z�T��iQ�U���4����Y�NF�龽D��ߴw��i������ֿW���(.H�[O�8�Y;
wK}�<�1G �'��I=�㔷{��KU�4�RV�jZ���%ۉY,�b��,ߓ���b�U���NƄ����mi��Q�#f�s6CG]r*4�p��Wm�r�"�"������;�(z��c�*�o3������.������ﾐ� ��믧������@�(J����������  �	*��ް���o6�o<�n�խh�~?::#��1��s(�mX�e�5[r+�sW$��[�'�*EN#�;�chܮƓ�(9U�ZZ�aYwf
��CTPN�V	�i�[j��[	%�p�;�$Ȉ2\���i���+r2��K-�����!2�2cq&*VE^I3Er[�1��P�
Z���$K`�L��3#h�G(�*e�9I��nQ���'�c"VQ!����ʌ��N��T�EA6�m���$�DPde!-ē."��
6\����<5�����(�E/9HAL8�H��J� �
T�,h�R2���B��{Dޖ
�q�,�x㮹%c�Rj������i�Iu�$T&�ɈWL��B��L�C�H:�,`�V�o-��h�؊C�%Sh��]�mr� E%P���!�HM�f9W�Q�#�ƛS���1��BƵ��V2Y-�-c���X�$���'%�]�q���rW�����$3�t���G�����O�˻�����ӝ��<��$�ʽ�{��_xwv�KΌ�p�}i�)�V���Q���N�V����r��*J5N���lb���1;xqN>mB�j�)ε9�k�
�)�D�=�=,{+DJ��v����ud�mB�|8�l�BsG�b���o4l2CΛ��<H�AD=����,�l���ِ�/�"�>�NG���+�sc����ܥ��ӣ�Y4�K!�&�����)W�շ���o<}7�6R�sNB��1�U��7��=���:N����|w�/i���'R��ᙗF���2!��e�&�ĩ��:�O6���uo��~ukZ-kuӮ���Z�4ֵ�Wi�Q�����**+BBʺNWN+Ea�u���)�x��1�O��Ɣ�o~j��L�vz�l����Jw�Ot��p!���,�ሸPB?����"| ��ۑ���L�^s�Q{�1�S���]��v�R����v�B+�f�z�^(�/��r���wٕ!~J���T������f.4�6�(��?6�kmk|���ZϏ88Cbb2�,���[���QQZ��I$�:jIS�M�7ʨ���A�����u��y2@����f$����/^�x��W)��V��C�>��_�b�a��L�+���������'iW��d��Ök��
π��Ar��`r��2_�}���ٱ�@����i�o:�$��d�is�^3�χ���#��Q�.·�^oI�+뇓v�Ɲze�>2e�<�Ϳ6����~ukZ?��N�N����|�Ē*�XE\Q�P����!��D�H�P��Gm�
g{���o� ��B%��Ş㲰Pd��<S��B�����O��HN���8�>�2C�:`pP���.�4C�I��}���Nc����r��UJF����C�E�Kh���M*�ɪ莁���fl�4dl������=���A��4�{���<Y�B��<(�E��cჷO=*;�֯��Sm��ͭo���Z�k[��N����y�MUn�/=����v��t|�ֺ$�.-}�*���Sm��n�%.G/&f�בQQZ6f������s?g������_�^A;x��x�ì\��x�eC\��YE�Lf���s姾_k�"����KE�[ϥ:��7��Z��_�n{*e��������G��*��V��)���8i�Mn�����<$���8��!0�n�Hm ���g.�U�
��͎}�0�>��z$�:���|��!O`ٳ�����G�o�ԹiQ$uā+�y>vl=��+cZ�!��th�O�d�t�g��s�Hz���7��`���-�F��[�À�8��=4��'�ߎr�Ä8����&;��4<u�]��eT�@'��0�7���
d�J���ѫ,v?%�K�Z@��$:`��G�ο:������T�~���`�f���J������А��rBL�HC�'GFyۢ���>�u��#Ύ��I���ƹ�x�)�4��m��gL����<j
#�a��/�8�d��B���	�ۦG/;豳d:�����FJ8f�~��Ђ4�a#��҅;%?l�^���8$���GL�0S��C���#�A	#����jQ%N���P���8d%!b'��Vn�*��%���m�n�:������T���:uq�7m�w3	q[��EEEhHp�F0Ѫ�ɲ�t�ܐ��(��0^(,����V8:�xU[e������uOۥV+�k�8Qe(��s�|���¤�YݚF�j�%#rr���BI����s�Ac���͝l�&Ð�-a�PY?�����`\�ذ��t��C�Y�dD���p����`��'秜;�l��#-�}�7X*��ڥkLu��>R�|�ͺ󖮿:���uӮ�ʗ�I�dFU�b���ID>08=��F��ād�C�)��j���z�D�*3zBFJ�����8�a�Ƀ!�6Q~6E�hp}�h�0�{���2B>�G&�GcN�#���GF�6lv�)�tG��t�8zD�`ʇ��}��=X��lx><6;�N�x=u���ӆ``�GN���d`oÇ����c�,q:�N<��[[��?:���uӮ��/f�������Z�ӕ�AJB�J�s��x+c��.9���iXY.wo!���!~��9M�'̶�Ц���`�t�;N���ӛ�h����oi�a��Q��e۾���z��N�*<{�M�6�J�z1KZ��o�Sچݷ���"oI�6|A�:�9<��'���T~m{�ֺw�{��}�>��"��n�d�e����-��N��6B2q�6!���6����!�}E�{]��9���:;4m�Jʟ�d�p�eC$��!�c����،g�U^��G�/G�4�6���dʆ�o��y�q<ƈ����I�)�('ap?��ä�!���8�<�8q�.Q�����n��a�A�T�[u��6���uխh�����Yq��n����U���"����׈��d@K�x���А��I���_W
�� %(�)U�2��h�]c���7�-8�a�:��8��+�h<{�c��|uO�o��o��u�Jx��h�x����Xh(�ɦ�f\�������;���ۉwj|_n�lT����j����-3���fo�!a�l��h�t	!d0�6I�s��ٲ�����Xz'Y�X�������g����,���x�,���"#����E"#n"#��Ȉ�����l��!B�F��TmF�"8�#��<�yG��yG��G��\i�yeȨ���E#M"#�"8�<�>D|����Gq�")�F�Du�#h�"6�#�"�G��U�6��F���#-#Hʐ�:��iH�"��GDy�|��4�Dy��Z��ֵֶ������8�6eB�!jS,���4��U��{j����j9�C�����g���v��v�>v�gr�S�΋���[**)WT�'���o��j���Y�~Q�M�{G��R�.!��<�K��ʶ�dN�c��Yr�	��jٹl��8�m��{���c��-5���y�|ձ��~+���s6��_5Lt�ys���D�v�nd�h8�6�#{fy��U��7w�Fuu�I*Y�Uvk�q�7�JLd�����{8�@�(J����������  �	*���;����� ,�$��������߾� �
 *����{�&�C�4���yn��V��֎��g��W��TTV��뾆��a���/���q��4^^���oMd�Y%��g��q��_8�h�!��&HC�g����֤4UQ�ǚph�t ����m�J�����=9�Y9�G�eK�?b�Cę���Oŕ�/%pl��SrB2O(p�2h�x�������ّ~6��o�������X/d�6w���%UJ���(�Ŷ0�����9>|��qƟ?6����kE�u�:˘�3EW+O���)%8��9�����	���{D�;t�$�.�8�{�v�I$��|y����t�0`bW�'��8C�WT����%��#���~<G����M៩�����?%���C�6�v�,p���4h�!���`�ۗ���L,�$-vfI$�:t��hr:4!���
ۡ;2J��a�x�}=+/���$�Ã��`�C.�8p,�؄�k��f�8�L���;�-x�ͫI�u�:���?6�?:��Z�kG]uN�����y3����Mzn���J��';���]���vv�G[J��PWq��Ҋ��А���>8n���>����~2u�U�\j�ŵT�Zz�7�ZN�R{���l=9gџO��S��;È��G�9<p�==�B�-
��j�Xf]�kXA[.xˋ���{�!B�;S��ޮ)���F\e,nv������'N��}=�s�����=vP=�cc���`Y�:2���>)O٬#m���[)O�Sf��h�vC�Dx�Dr䦝l�UT��К!F�A���$�ヰ�)���z5�ݳ�����0���;�(,��:ū��Ob�Ɋ.���+�eI!$���v6z������A��(w�w.$��|�B	�Q֟#o":��Z�kG]tGFp��Ú�MPeYۏ�ͱQQZբ�~���!쐠�=*D��G�g!����H����Ҵ9�"HH���*�R+����w2�Nģ�'}&����qz�;63�� I6�9�XY��>0?;��3��C�X���ѷ%l���w��t���_��Z~0@���2tw�h�dӉ	 +�a��U}��a��A��_�>*J����&03��w���T�v(�Ju���6��:�]Z֋Z:�tMԪ7l2��L�E�F�`S��=����О�Ye�e]�q��<x8�m��Q�F�T�!�kSalu���y	��J0[a�F�/�Զ(D4$���W�:�F�۲��>!ܦ}�1�3��4;C!�9�%nz=8h1���A����}�\�,��![�CGN���h��\��`Yۯ�UYz�$<8r6d�A�a�䧡���4��q�n�6ҟ�|���m�_�ukZ-h뮩�\��^�cU�h;f����ԡ������'p �X�2�M �H2`�M��=A*-F?-��Hp|[�q8,H��l�v��)e�n㕔��ّ�lru}��nil�a!C���G
3�G�����s7.�^�ުj��p+�<�X˒�[u��q�Ћ��MMx[��6QF��6m8�,ٔ�p��u��M�����4�q�,�b�1�mO�[�-�ߟ���-h�"�u�:˘�����ε�S��IH��T��y��\P�,�ڒA�N�&^�v1���􊊊Л>�6w������������i�֫:��~0ߓ�8�/s�:�S�>89�N>�pB^߻�$/V)��M�B��T���k4����^��կR�SXjt��Y�Os�Qi���^�F����%���FrR�P�6�&R�҉i\z��8U��~3�7q��~�K���3���t�.��C�;��	ӣ�4y�F��B@�>�ohra뗹m���G��óƞ;���s�<�Ҡ�꿿d����F�m�qS�K󝲱��A�$�q}r}��@�tC�l���;.B�66����$$!=���i�u�[��kE�u�:3���������>��%�*�%�[�y�0>��||r�l�O�*�,1��BM����i�p%��w?g��Μ_Z�I&)-�l�K�)=^�J�j����c�kǓ��l���п\�}�ip`"�x;6C&:BI$�٢�:>\D�du*ya3�޲Rn��JX-6���i��c�l��[�媪ꪱߜ<�`��{��o F���M=!&�9N(�6{�`�(��ύ<p�պ���Z��S�����Z���5����d�S3Gy�TTV�޾�oԣt��v���ss�g�q/f���T����O�������M���WD6s�	�)�#ݞ���f�ܔ�ae�G��	u�G�C��v�Y.u$��J�@�Iа�J��v���G�O��ܧS���nx41���!�'���a������p<V\�J��Q�����]���K��J�����c����&�oٜ�У$:QÅ�,��ߝ~un�h���:�Yq��~c_�9ūa�7^�Ђ��4TСB\&j��EEEhL*�Y�&�ϵ'�9�r;!�!�CY4uF����	#~�`�>�z�ѸH�fj7n��� l �J�.h��g����9݅�g�;�4�`���2`z��1�9Дw�\�������:����Ǟc�����[,�CM�u�3תP��H���#��	��Y'C����ƃ�A����VƲ���e���m�7���o�<DDiGYB"��Dq�DGN���L�C(B�#�#M4��H�#�G�uG�F�Dy#��<�����Q��m��#�!�|��H�8�#��#H�6�W�mH�U�#h���:���>F��G��G�|��y���em�!C�!H�"2�#�"<�l��N�<�֋y���"#h��ִZַ��|��B�!E�~H~>�����9��DM�ݿ����=7c�k�^��؝���q�UV%[�z�_O�^U"�_9�q�ݒ�y�����ӝ;>~G�����FZH�DE8���v{g7#�=����Ϲ�}|�*���>.!Z�,'����i����5quUʲV�ކ�=��˯PFlf�"e9\+߸o�����}E�۟z�����TK�"b~mS�n�*kL�5jgZ4{�#�Gz�C:�N��'x��bݍm�H�^���E����q�M�w�~���å�댫�6ḎJdnCw�ey���>�w���s�^�v�}��O���������]��BF.B��k5dԐ�R*r�*�m4J��2:�D����㉉$�ݹ������)E+N�G骪i�,NV�u]���8���)׮�w�s�]a��@ �U_��wwwwo�@ �UU�ϻ���~�  �$ ����}����w� @
����yO2��<ӏ<�V��Z���|x���O����&��+-�&�	j<CD��$�-CM�*(�(P���I(��4R)kc��+�C���-+��+ ��
$*��tU�Ɋu\�B�Z�q;\b�"�BFT��X�L��c�ҵ��e$,-)��oA�1��&�X�Q�1$�"-��A!.��H��e2�1�N�����m�*)1���,
Qc�����"#���F�1��
��(��(�Cpy�AI�x���2���"�]�K
�##�2d�F�rZ�Yk�ad�m"+B$�It�e���!D1Ԑ��A7*".1��2�K!m��Bj�4�jHCƈ7����+�����QV9HU���'dN�k�qF��K�L�V1ˍ�e+���uA�bu)��"�$WQ�ERmUciҊ5m�-�Ve�)ERH�Z�b��j,��"�X�؜h�H��M'2(��$)$I�� ���1�4���di���Y+�Z6B9G-�tq�:���8̐d�\��q3"�zu�TgV�S�Lȵ�)XAi��U�V�|��/V�T�T��jU�
�MJ�T-��b��_{��"�P�VK��U-�Ӈ�d��<�K�]�;�lW��\*\��OLkYDBݦ䌖�֫j���%a�i�=�d[��v��:�v	|<8�s>��k�Ч���l���{�I��� �+�Ѣ�;l4c�C'��$l;�ph�
|{Rᦙ�Y�Re���<�f��YQc,����.JvN_����rh�v������%~Ͼ�x<^C?7�I1bHB����ݥ80�k渗8R<I�<��6`hx�/UU�a�7�|�Y[�?4�ߟ�Z�Uխ|x�ӄ8&��Q-O��m��f7P֯Fk���H>�"���'F��L�4`�tI\xŘ�P�B��+�E"�������#9X����a!,,�ǸK������!�|S i��!�4I�r�:jOd�IJ��f����ܽ�2H}f�v*l������)]|6�ُt�3��Oo����fxtO�^�뷁��!F�:p=:l8p���'��:���ṥ��m|��ӏ��?4�����qkE�y�:ɳ��'�D�E��Ċ߽�TTV����DV	)��}I��Ex��$�|�jI�D3�D�%l(��݆̍����x`z8e|H$3J^��|%�p|^�K_���ą�$0QUESF��CmG��o�My!っ��!;=��g��>�L8ovMnI�(t�xa?l��$��L�64
U
V|�Ú�����Q�(���iE����Z�kG^uN��X��)TQ�N�jl���T8�4���ИW�9�}i'J��+ԝ[l(�I0����ό�V��w�x�Qo?�h����5usl��5jo�0�&�V�m��FD%P����I��`^�lr��Xl����k��9��M��a�F/g7��,�%ZJ*�~�=9��#���泶+~)��*��G�~['�pXJ�*OdزBCeXl�%�1��:����o�2�4�<�?:���֋Z:�u��:L�������#���%��F�j����CM�f��؞q���J���H�j�Ibr�􄚗�clm�Ζٲ���k7vE�M�k��Q+S��'��]��r�r��M�p�)���ϕ�R�55px��K^���KU*=�8x�H:���9��+��t�3��/Χ�ld��;r�X�7(Bp36��=}�^=�B��i�� ���W���(i4?vMSAc�!���2���l0cs�+�a���Z�CC�����1p%FA~<�����5^��e����{(vs&L���}�x��lu��,ɗ�k�YU��h�rE�N�K1;q�!ӏ�������xџ4�c��2י���J��o9�Ut�*u���<�?:���V�Z:��u��s�dn�X4�֫��K��r�CJ���(���%�M��۱�Wa����>dK��7�t 3��*�{��שͼ�����G#�;D���0�|hv:%�4��N�L)�z�s�>��O��X�c��HvHd�,��r�������$�px���L2bvz��şu�M�
3�BO�cC�͎J(6d6�Տ�u�9/�ʺ�^?ci�8ˎ��H��խ庴Z�מS�����k*iE�G��\EEEhN�{�.U.d��5�X�ҩ�C����t4�S�?tX��:SHf��zh�gGJ�B���d,�g��^��KG ��֟C累M���o �[���gϘgq'�
]��,2q�fy�#&��`p�:�:J�h�r� x8w���8�>�Q�3�@�3�!)�^vs��t=.����2d,ʛeo4�H���~[�[�����!�63M#q��.@��f�QQZ�V�M�����k�/q,H'�:cN��q�Gdk���k5��8ʯ��?���?�24&��"S�v��C2]3�������&G��:P厭��`ٍfU;�?�*�_��·G����h�����F��8�d�s>�d�`S���͍rL��9�%HBN��3;���`"��:i���yn�-��Z�מS̸�+U��e�6ٻ�5m��!�I��kÜG{��vޥ�S��#wdd��A�h�����f�g��TTV��a���׆��_���]��r�����6x����w�Į�=:]�A�;���i�Z�r�sk�9��CI�fɅ� �m�C�<�m��>:\�÷�G\!ʨ��*�*i�U6�q:#`s�7=~��nd��g����K�v�r��n��6���O�?�t�i�*#�3�ÓH[��A���$�8l3��0>w݇�4��mt�&�Ag�<B�K����
49�S�6�t��ӣÃ�c��Qa�Jx��Y�bx�6���x��O��R��O���S�&��8�`�8d
b4�M�4��Q��;��ǂa~}$����Sl��-��矝Z�Z�E���Ǆxg�c\�T��Ћ0hS��**+B4��et�?�
���r���O�=�c�OBu_d��(�LF��	�aӠtw�B����l�T`vx�$	2�mz�$�)�F��z��Ap�gO�V�$8���z�'N�6J	&\(�vsm�:ss��7zZp�ӧJ(#i�6��|�p�s��L�S@�t��]�49,�ɣ�!�M����s��v~3�'�vp�hv�,�����y��:��h�l�E"#h���:����#��"":�#�m�HBB�|����TiD|��9*�����<�F��yDDy�u�(�DF�2��#�!R#H�>De|��#��6��m#��DSh��"'����H��")�G��U�|��Y�YF��#j�X�!��4De�#�"<�l��n����[̬��h��#��""��qo�2��,�!������[�n}�������X_G��ۨ����S�=~=�����P~�N����2&jn�z�-Sy����z��[SnZ�9�̍w˓��ve�
�|��u�̺y���|�s�'N���=�-V�y��a�7fym)���~Y�}��6����Vn~*����1U+��w��F㌙���G~������7�]��[Q7�����o��F�{�j�zЧ{ճ�͚�S�*��þ`  UUW�>����� � UU.����� � UU.���� � [����>W�y��yn�o-n����N��쟽�EEEh������C��`�ίv�^��B���7�lm���]�Ui���_���Y#���:��0���c��S*7.~$��/qmə��Mb������-���r'zHBzgr�W�٦��u|J/�a����ѓ�'ܓ<��x�{:ie���G+�gSl�W�<��<��-��Z�מS��\�;��h�TXE�`$~xА"
8R)0+��q�g듒���[��+er=��O����m��5}�k�ލ���wzq�g:���oW�a�C���؉
O��%Uf�A��������#QZ�����>�����|Ph~<�`x��hf
b��]��C�>5϶N0�9��t�
�C�����c�c��FBBHG�����z?9)�{AFHd��E�0t���_����-h��)�x�kI�/��;���ZA;'g
����ڹ����U*�m�ܕ�H�T��d$�y���7�rA��j�{�sGx���I��j�}�d6tL>�<[�9�RmU��i�{I�8�|��o�2����)j;Ww��[�W+9S]�t��*g�"�K�ֹ�]]��jR����g��'�ۓX)֪����$��k�x��8\��0Ͼ��v$���t�v7$��	P�ĖWs�ҷН�ؒ�,me���82�,r`vi����}�����U[��gC���:.�j�i(�T�qD���'e�x���V�,v0:1ˋ|v�RO�u�#<W�[kZ��張��[㧏��-��Nϐ�*y��ݔ�3R�Sk���**+FS��^���A�D6�p�C�ۇ'�����a$ ����~�ÏjQ��2�$7��8�K��$���>x��nP�''��m���_ΔE���S�UuO�i�I�f������F��g>����i�)�UR��<tu�΍�������8��8�S*y���N����խ��Z��Ǆx|�*�K؆�F4�	���**+G
�]h�[+�ep>�YG	$�:�B@~��QX�a��^�h��aX,c����Ӑ��L����p��Q!7�x·q<!4��<0ہ��ɢꤪ(6	�v�O�0C�W����]�ٟ3��GRcCgh�����Ie�U^/�]2���I�C�!�٬9�܌p�i���N�����-�Z�מS��\�ٺz���f���1�i/5>�"���`B�Y�*��o6�v��>m���>c��I�+�q�#B���~B���wu(e��Ϣpc���u˲����#�*�d���6�Srz_]ň@��p�<��ǩ�wnmv�ѨSK��e�d'���^�]�1
AΚ|��Tu��f��f����۽���	�ϴI�e6���#̾a��*Fb��6���~[�Z8�����U��ߔ��ՂQ*�����jeIE�������cݖ�/ �K��U4�#`4ђ�u�%��U]��ʷq���clm��QY�ֺrs��R٩�5m�,��C�T'3J�,Řjp�^n��*t(V�������RO���}�����U��~(��Q��ֻ]�L+��R�g��Z֟�w���bV$�y��+��Ò���O>;�s�yb�P�f�*��;0�ڣo5d�89�$��S��?�C�/،��h(eϽxی�ś�ď�,���lk�^)�T�V��c�J���>$d2cd�:`0`��m�z�[t}�h~t.x���1w���i�el�^����hp��Hɝ0��������r�>iG2�]�[f*��-�k�bˉG�G�����W�L��������6���n�-�Z�Z�ŭy�<�xn󥤩w���˯f"���|W�+՗���r!"jf��j���g=-������3&]�6h}�UV�BI0���_��g������
l�� ����*K
G7*?@�`����]6�	�R��0EJ�IS��/�G��Âѡk�^X'6>r�n3��F{]����ஸ*T48��6�����W���zh,�+j�Hۨ��?-�Z�מS��sx�Ub�ݐٱҢ	4�s��clm��s|�OZM��RY�8|ƙ�)^bֳ�3���=o8�UU4p���ۤ�mu�zbw;-a����9N�cd���cωw��Ĥ���M��뗘̧��"g�fGe�wM�$�������73��<��&�B������\C<���2*V�º_����׃�~�_����Y�1�qN3�F��y帋[�Z8���<���t��]%
���Ɯ��kclm��~�q�F���}�z�&�;���1e�\}��$PHg�0y��g�GD���l�C��FISfJˠ��;�'�8�߉�.=�(á���8�Q��pxȉ���vi�Ѵ'5�<��	C�烦�~���BP|VM{~�w�~#߂�8W�j[�&6�5�[o��:���C甈���q�")DDuDDq�>G�2�B��B�<�"6�2���qy�yu�x�#��"#Σ��DFQDD{j�GYB8�F�DDڼ�D>G�mF�eR)i>����8����#��<�#���ѵ4�i�iT�ڥV!C�"2�"�O�F���e�]|�Z�n��֥�DDuDDq�>G�m��ҖYe�YՔ�3+ϕ���}�97�է[��n�����os��A"�ٿTҽ�>��6����Y�g�:rH����o4͸uy���|�!�G���q/w�oY�)��j��j�4���F᯿s{z�J#빨���z��|�J��M�M�ٍ]����[Qv3��-�f���ʋ*o�Uo�MM\�y*z�*WA��a�T��j�0��Lɻؙu~�27��+ٹY-fv�ogN�#=B�N*�ƘG_��ڪ|Н(M��ec��e�Sme�FEv#�KZ�&kbI;b���oy�E����t�p��r�&�s�+ܫ���;�ϙH��Em��;'Ї�G�%�|M�*ݱ%Z�T���;"x��vՒ&�n��H�UB	�F�U�TK���R6'aT���Qy�[CIE�q�[v�,�T�R�W��)�J���jj%�]�~��m}��~~ B 
��>�wwww�  �UT}����� � *��������|  � UUQ��˓\�J�+��yn"��֎-h��)�*;���lI��+E�Z�w�QdL��H�R�HB6ŕ!;�PHC�(�1��(�E��X�G"YV%l���)DQE1F!�!��!I�&����H�"��%&,j<�q(',I�Q1�Ą�YB7��j-qm1$�D����F$Q��6R�T���![,�<+%dQ�*ʠ�RF7bE)����1��<�YV:�*XZI�\���X��:U���G��r����J��KJ�-(�
��� EE�V�$�Ċ)F���FZ�cC�XX"*he,Ɯ!F��B�< �R`��Yl��*R)JJ��H����\%��ڲ������)�m��Im"I�k$�Ud�9OMuBR5H����7
\�T�n"Yb���JD�%�j�d�������cr��ܔv��J�+�WVF�DV��ԕe�ӐR$�eq�\�ˎ7�:�,c��"�[%n[����6����e�����y�<��'�x�Ν�|�Wtb�T�ј��K[K%.f���l�S���b�X��N(�\�w���߈t+-��ҩчz�9�8]������WsWXŽ58���i��Ώ�^a�Ս��֙�8�9�nr�u�(Ȉ�W�SO�}��N�2In��i�����#ǃ�����xO=0�vR[��CG��~�}�e-��i��Z[`���;���M�&'1]�C
(ʊ�%��=��S�����x~x�rLK���L�_��X�f��o[���39�tz��Ezh��-��k�R/5��c��Ոm�:�H�ͼ���o-h�V���t����k�f���|�wr��d��m�O��hHKgC�ٖ��O�8o�])Kű�:�i�¹�B��+T�)'�7*�����<I%�ck�2Ki�!�µ$~�*����L*@	"����t_�+|�M?��/7U�'U\���T8|� ��C�&+����Ӄ�fUQ�`oa���e��N9a�{�O4�ߚ~i~Z�Z��֋qh��)�Zsػ��ri�g�O�			(krI>����A"�,6j�P٧�c�	�{[,�x����ڲ>z�v>6�����n{G����:��C���������f��O���M��j����&*3�Gr.45�o>�������˾IW	>���5��a�Ѣ�4=+�Sa��9ѧ#C��9�Y��Ju��ӭ�<�-kykE��u��<t���^m귄i������y�g�q�}7�����|�sթ}��h~3��L{�g�"ݚ��1�I
����vB�<3:w}l���6�������G>Ζt(����~X�c���pѣ�,Mj,Ó"j}aSj�Q����A���L���$�Ѱѿ�����Ij�""#3L�2
,�L��iJx�M1֞i��Z�Z��֋qh��(�������� ���a�ƒz�c�wo5>�w"X�h����T�j-�I"E[���P����{�zJt�~E������=�g������UN�r�T��5��*K{2'���*Uq�8�*�\������;�׳V�N=��Wr�/dP�P�96M�M��o��m;��-���i��-���PO���(�C<������l��@��M��tHy�ht7�����0<��c��N/�s�<����eMs����t}� �Ua\�O�tM��6:>l���F��2�W��3�Y���y�����e0g8������Z(ц~<�˓0�x I�6��q�G�����֋qh���<t���U걖���B��ʞ�h�4$$%��X��Ӄ�4�퇰}�U3c#�Df�G$ BI$��h4:�Ƶ�^J�ٷ�/�d~5���$��<+5*�X�۪<X@��!a�����ϳ�aюof��c.�s{���Eۥ3�g����0�>idX@��p��͊f,��iИ4FC��&����8�3�����VV�j�~���~�����٧�~mk~q�kykE��u��'�l�ǒ	�bDX4�	0��!!%�I�QT�֤�!�6�p6ޏC��y<��㸌� �!Y�N>��Sc���r�G�<��T$���<��}�x����}�⻼F��~-��vF�D�ݒ�����$r��>3���>1���}%|i�UA��M:0y�hh~��$>a��\��X$��*͵[%׺lQ�}��K��'�!	2`z86Q6�4�����ַ��[�G^yO!uqyɌLMDg�����Xp��Y6ƍ5�7���<�����j~�D�eū.Ėu���;b��B����ٽyy�u��u��3��"4<:�!��a׼4�r��6}f� X�pz����$K��t|l<t���뗏|!$,�����%E�����z&��B�0a�.tS,h,-���'}��Hm~i���������Z:��x�K�{�l�hX�r�_yvKk����]>��v{��QV&񦆔q޵0���%�����9�P����}��۫�5��NP��Utv��Pj�-�tҁl���z�R��#.%B�H��m-R#���ն�R��
U�5ښ�\����E�F��ٲ�]��f�wm������p&;����F�oq_r�YJ2�+8gf}��#�P�03D��F�a�E�<�.�d�f�l9��x��*�?��d=6:��a��ǂ��ތ8N|�!n�1&�ͽ&��͜>%�8�Lx��w��?+[ޫoլ|�kZ[8M�>s���3���CE��I`��P�*�:F<SJm֝i�ֈ��-��h��)�Zp�R��R!X��*�V��BBBXw�I9m�$���;6d�ô�s"ʒ:�+[��v�[��I�����va���c�C����3�!L!'á����2LT�����Z��'>�����}�}���pu���L1���6BϠ�r=�1��}�:h�a�������ZY��j2����6}��;�.�������L1����iǑ�|���|�H�̼�DGȈ�#��DGȎ�<��:�#�F!B�"�F���TmDm�#���Σ��<�#ȧ��yy�u�(��#h����uHG�Di":�"#M���F��V��FYDR#������3U�DOUF�G��|�h�H�"��eR6�U�B���n�Iʨ�4�2�κ��QkE���Z�Z��#��"<��G���P��Ye�Yn)�+R�Y����3���=���ϹL�y|�/�9��M�ut�rڜ�SY�yu5���w̡�F�Vђu'�����Ujsm��Q�/-̩7�21��xFF���v'��p+jf����쵹TZ�0:k��P�Cq�w,W�J�݊{I��-�٘k�k�^��w��Wk�,�b�Y\;����n���:��i7�QuN-NG�	�����<�M�\��z*���؇fT}CyɕKi�xp ���� �#%�O�ܜgS��J�����Ev\[���eB����M���  �UT|������@  ����}�����   UUG������  ����.\���^i��yn-Z֋mh��)�K4x�VG�����<��7�l���[��i��5�1�Y����
6~�::2`W��@�t�bhr6q�������˪:|Q��-��R�ۡ���3@b��)�3P����"W~U�V&|����d����D>�l�7�|Q'G�	�-��0B�*���Ȝ�#A�������A����
(�M|ӭ����ukZ-���<��h����-���(D2��I$�#)��Қ8;��z65�w����_��˫��q�ah'�������34��nM8q����!���~ӓp_�&��L�{!$a㛢�&77��%����vC鬎��?�%p:*X���5�xnôU<�}�8g0��'(��C�<S��qh�-h�����u�|�h�ol�����y�Q�U�xK{�*;���sH�K�M�8�j�V(�����7�~ԒI����!/Ŝ'���ҽS�p���׫˥<�t�E��ҭZ_a�g��y��Otd7��o������{۱/?I:������TK����q��㻻:�?!�R�(��dMfLA�w�Z��f������;�O���8�~�����O�|܋�����C�7��5��֯e\-�Ig9�3�ˏ�=s���M���;��@�����A�c����	]��g-��R��e��Բ؏+s
aC&<·|/~x��B}9���KcH��,�]��d:29g��)��`z�.�x`�f�j�i�B�t�n4������Z�kGμ�t����~@/Ѝ�.�z8����)$�6!�+eY��!�Uf�>�zQT|QOK�x=�R�� �}�H�DWvF�V��N�L�����!�h���y��î{SD����m��ǎ�3���M�.dq��M��˳E���;t�s����w{�l�#���]V{{���Fx�l���f[[Dw�JR��b�����\���l-�E!!��p;�U;���)��q��G�q�E��|��)�Zo�+*�ך�h�B�RI${���Ĉ%�)�J����q!	>:gБ��|n:���p�L����c�=�G�|˜�b��,�1	(�y܅�	�����R�*J�D�rI443���o��G�'L�sϨ �'�W��!�)FAY�!5q����Bq��6?-d�>`t�|9)�S$eO�i֝m�����֋Z4���<t��ڞ�jb�4�[�$v�$��n׽2���2�8!����$>>�K"Kۿi#�&���-�U�rz��p��m4�� uѓ��N�0�lj3ch ��o�nHk�����9��x���h�U+3��N��j�m�
�&ޙk2��O���d&����(��$I�dKEw�2�m��&�C��:im��~GQ�z��uƞp����*<���}Ȼ�9��T����}��9�u��F$�q�:�;Y��R�H(��׺��$�Gi�v��=���n�l*�#��\�S��j���S��� �n��g�a�S;��xH5i6sp��A�վ����i�8t�2�v%�{!�ڡҐ��G+9c,�WV�^Y��vb>����	s,햅Sx}ɮ�otsO?{�o��&�w��i7�M$�MY�G���~̔���d��΅�>v�~2pi��I�&�{ϣUV�<���0�^���D�����§J�$��'ƝƂ�l�	����7�e�˃c���'��~0p�b���[�z�p@͛�jOD��x��"��G��b��(��i1�6��iu������E��[o:�\!2�ߍ�4�9v��9�;�$��M��d�r:6h�3	?FI i������lt���w�w!�4�>Af
��b�|hzk��m���	Ҵo#�K��(~ ૘��g@�4]�';S-���;>-��	t���rcTg&��'��L�8�!	6��͒jUB�e4W�~4T'�|8|=-��������_��!����fD�c�b>CM����i�ߑ����E��[o:�\i�U�j�+��?,I�*∈�aTA��$�Hퟎ�v�*����\�=�i�K.|}��4�f�-�̐e�\�;�\�_����r�Y�E˪^5B�g0�:w���S�esc��ҥ5���A�6V��\�����f���ʂʐ��V�㵢qڒk(�{!��4�g�����vRJ�3�+�5��*BB�:^T!%�Q����*���JyƟ�[h���=U�>,��6YMҌnĴ���d�H{����%�*�+�d�b��2I	��Ϟ�}�X���%�eݚ�ƴ�C�W,���n|̇p�͗�b|T����
����k�$8��Ó&Gc���0��O������ٚ������q+�=��COG�ت��kf��h��W���L%��m�h�g[9�o�ÿ��r�R���UV�4cl���oѿ`�+�Z��|+����ݓ��D@E��f����-�*������ �������7m5���DD����E�h��-�ZZDŢ&�h���DD�DKH���"h��&����"h�dM--c�ni4ZMI!,�MM-)i4-�I�D�i���4R�i���M�&�[KI���4��hI-;�4��KM��Y-��I-!,�h��PD�Z�kD�I-"M$�md�i�HI,�m	$$id�D���M���$$�H�I6��$�$�$�%��I!$��i�&�I,�I4�KH�M$�I4�I$�&�Nq�$I��Y-�M�$��I�HK$-��i�$�$�%���BI		$��m4�	$i$$�H�BI	$$��BI�$�H�I!$��i!$�I!!$�i!$�D��I��!$��i%���Z[Ki"�4�i&֖I��i%��L�6q��ZZZD�kKH�D��i�i-�id�Ih��mh��$��� ���H��MM��I&�I�"ēi���I���I��ZY&�ZkH��-5I-$Z(��l�%���ZIi���4�M,�%�4��4�iiE���4Z-"$��i�ih�Y�m,�D���KKDI--6��ih���$����&�q6sKB��KD�MLMH��i��i$�LMIE���i�LM4�4MI�h��bi����4��M���Ѡ�4h��5�̍lF�#[d9���CF�#Y��#Lu�p����fC��gM��#FF��fF�h�4kkl�3B���t�I-����3F��Lѣh�#M���CF�F��#8m��dh�5�۴m�[l�3F��X#i��q���`�6�ш�24b426��m���٣F�Ѵh�h�k6�m�m3F��F�h�25�F�F�h���Xѭ�4؍F��4��dkm�[dmfF��`�l#L#Y�ki��f#Y�ml���5�5�4̍�L��5�#Y��1b͐�гd,4!�&�m���&446�b̄�B�m����f�Y��ݹ$��4؄��LІBm����B�B6@�ͦ���5��m����i���&ɶ�hi�ɬi�ɬɭ��&���bk4�[i����kk	�&��-��d����5�Ma5�4m5��2l�����&���kf�6�̚2kg2n6I��M	��M�k&�Bl�M4�M4�5��Bi6I�4�I��M	��i�&�i4�ɤКMi��;�m�i�I��Ml�M&���M&�M4M4�4&�	�M	�КM	��l��i����&��M4�l�[&�Bi4&�M7�i�ȚM	�4�M4�4�D�4�4�[M4�4�I�4M�MM4M4��M4M4�l��i4&�Bi4&�L�"hM&�h�I��&��s96D�MM4M	�КM	�M	��&�Zi5����dѤ֚$B-FMD�"�"i����kE�!4dD�D�"��dMd["h��Z&�E�--�D�CZ&��!4&�#&�E�4,�i����\FH�YBȲD��,��E��mD���HkD��ȴ(�։���d&��&�"h�E�4Z2D�"�hM	�ё�B"Bі�D"h�E�֋DE�h��	���nhZ"$Z��h�&��hDd�дj��@�#Z6�F�F�F�B�m4&�	�4m4&�	�4m4&���4uӻ�(��8Ѧ�Ѧ��B�4i�i��4,��MM	�4kCMh�!h�дkBѵ�Z��ѭ	�Z4F�4B�h�DkE�u6�#Z4D�2-�ZCDkB��h&�BдD-1i�b�DZD��-55���DE�� ��5�&-KD[����>�s�1t��iM4�c����~�(��2�6ٳ),z�}۟�������k�g5���m~��/���O��Q��u����q��?� ��������!��h��Zy���V�O���'�G�+��=o�5�w���'�`����d�x����#/����g� ?���W��O�@�������ُ�l�f����o�Xf?�n$�����[����3�~�?����D��W�������?���o�He�?&����\`}�g�����j��lzK�fı�����D[g�/"a`��?�9�?��h����N��F��Z�];��S���P����`e1�d������]y�����@P@k��,P� R��hU@�q@JX�
?���rٶ�m����wO�24���� λ�S����+	����z���߆�o��������f͛���m�-F�5	33$6�P����P������~�-xM�_�o/� ?Q����C���'�!?��W ���g�}�}��1~`m���o��w}o���0* R��B��o����������?O��'d��^��Z���G�G�_��F@�����
`�H?�|���?�����Q����M��g��@ ?Z�D#:���G�����]��~��c�ߖٶ������������������R��~�!������|��c������l���)9Z��B��nB?���"��!H��ۣ��e�Ж0:q(������4���إ�DT>O1G�cq��-4݊\����A?�<T (��@�~�����,����H���*#?�M����u����G��O�~�~���~������-.��=���]O�?�~���?��|3���EO�Q�D��h��o�'Çq \��v����!�c�:��ɷ��暚�5jj�VՕ���V�JիQZ�jը��+�(�YEb��)�V��jթ�
Ԣ�(�ڵ(���L�++V�j�)����Օ�����5Sj(+�
�b�+�


��b�AJ�b�X�V(+�V+��b�X���V+��b�X�V+��b��X�V+��b�X��+V�V�jVQF����)Z�e+QYEmJe(V�
P����VՔVVՔS(�QL��S��+(����VԦR���)B������MEmY[R�(V�[R��[j�VVVVSR����Z����YYB�������������YYYB�ee)�
�XVVVV����YMYZ��b����+VV��j�j�յj�
յ(P��j+VըP��B�B�B�2�Z�2��2�
ڲ�emZ�mYB���YJj(���++++V����YYYZ���ej���Օ�+V���X�Ejڲ��++QZ��[V��VV�Օ�V���j+jյjڵmZ�mZ�Z�յe�����mZ���Z���J��jVQYEeb�55j�l�����V++j�b�V+�j��+�V+j�V+��b�E5eb�X���b�X�V+
�+V��5�X�Q�Պ+j
ڶV�ڶ(�QL�V��5��MJ5jef�����f���څ��mY����+emZ�����+e2���e
���e1[V��+V�YZ�5j(��jՔVV���[SV+V��5jmYYZ�SQX����J)��S++
�+j5jj��
�e

b��+)�mMF��V�
�m[PV+�X�V+�X�V+j+�
�+��+��b��X�V+��m[(ՊV+�V��b�[V���b�X��jQF��e5jjmYX��ڵ)�������ղ�mZ��[QL�����ڲ��+(�SP��VS(���)����Z�Օ��SV��MZ�E
(VQB��emZ�ee5j+SS(�El��յ+�Q[R����������++j������+++QYYYZ������YYMYYYB���5el�����+VՔP��Յ6�S(���)��)�je2�l�Eee�e2�l�L�SV����L�VVV��+5j+j�SVڵm�Sjڂ�X��V()��PQ��)LV�V+�55b�X�V+j�
�b�X�V+���X�V+�V+��b�Y[V+��b�X�V+j�R�(յ2��(Օ��P�e)��Ee�S)[)B�)L����ڲ����)�S(�R�ئ)���VQYEe�S)[)B�)Z�VVՔ�EeeemJ�J�J�5b��������eemYYY[VVVVSVVVVVVVR���e����++++6VԬ�YZ���ejSR���
SR�����)��ը�ի+W�~����ߏ�����C� ���_��G�N?�?`y�������yi"�"2������8�!�C��ő[d����W���m��?�������;�;�)�yL��-���2�* i?�~�?0?�
j�������E-��,?;�?���g��=z��O�HFF���2�������S��/��?���D������́������S�|mDԟ�%w�?�K��kSm'�?{��#�O���������P��b���N��rE8P���v�