BZh91AY&SYcs�� �ߔryc����߰����  `a>� 
t����{�D�  *��`��|{��n}R	I;�� ���Rf� �  �5��� H �!F� -���4��� 
 ���� ̀ i'��A D �� K��� 6��q�� 3��@     � �  
  ���g����&���0 �F� ���%)&HC  ��h   j~�U* 2hhh  @� �� �) 4bh4�����#@ *(�i12'�I�d��)� 6��<�h�"4�$�  0&A�  ���wӻW)Hm��ra�D��7�S$�"I	9�D�̉��_������BC�?'���4�����_��~k�G��2�~f���ȱ����XK-R&�&��HTeFΛLa�[ncq��D���I�)&�6/5��m��mH��8�l�"N5�>=��������+����u�{����&��k��g?��|b9<��G�:��L����c�Ӳ��0HRN�N$N',�rw�W���zp|L��z߰�7Cpa�K�=��3���KK���K��pQ�Q��lv;3d��C�����9�a���f��6>��8ṟ�犖c�0���ft��83ө�h%%Tpe!1��1�Q����q�Llfxɖ1��%\��vs�U:�(b�ur��x3#�ce�r�e3�W��n��w�U1��(�Nl�`GM�vS.�gJg(�pf%Χ%X�E;)(*:��
��c�&�яM�e�c3�1!���%Χ'6�w��UGV��2�TV��e��\C#3۪�s,#1��2q.v���������cĮG��j�u;;7Į��s�T��r�[�������.T���pCN���L���g��|U�ʬ+#�L���{�W��3�׵�f����I|��|OW�o �|��;�i�5Z�zv��Y��S��3mQ����e8\lcE��+Y�W#eF��X��Ξ�ԓ�.ԗjK�%ꐘ��IR��C�fseV
q;֪��+: ��Gi��lS#���,'l%���ai@�+L�W3��됹u-��R�ͳ�!sڹ�K��,���_cE�d�2^T:N\�d�#0jٽ�`I�4j�F		U̓7�U19C�b] y�<�?3����e��i�p��r�Z+*�*�*�L�]�+<���t�NS�g3��˦��dB��_%�s*)�J�[�eFT�s����^�o���x���;�'[�.�s�Uԯ5Q.$�\K2��&t���1�՜h�w�)�F>29�i�Fb\�R�7c-J�݄y�T�c�#����\�:p�V%\璨��!}���3���t�tf���](aКK]K�%�yT��^%sȐy�<R����3L��2���o��7����6�||.	�(�t���;�;�����=Pz��q��+n�T���6Aӄ�dH3�<4=p�W�VU ��Ҁeb}�L��u��e�N7�Ux�ǩ���Xfa�T����?!�~�Uj��i�g�_��u�yW|�nB��k��t���(>�����	�/�۾�m>�n� i���a��E����f��km��y�!����ު�M�ۉ�G�ݻ�l�p�|1t����*�	%��$��-p�$|�pt������֖�����7�rK�2wx�O1�k{Х	�jv��K+&�mέ��k����c=�]�ʍ馌7D� �"b���I���2icJoD٦�8#h���`*�^dy���$f]�N������4��a:f�B-A�a7Om��1<ţo.��z�>��/m�+}o/�y�Pk���#���ZW�=(����t�Hn���O�h�ɹ��u�G-t-��<ū&6v�~l��1��� �(���g{�����K��6}��ׁi̭k��j�����'���ϟ2�{�_��� ��2뱛\o�y�0�> ={~� a�P������^��,�OO�%��سS�@�&	=q��7	��po�������
\Ui�O��͝�X{���6a��O1	aT��K��4w��w�mÖ�$�c��9|���r"BOӠ�*�H�����t��a$�ק��B<����Or}��t�3ʆ7(���X�l�.�yM7'jΪzT
Ο��=�tt�0�p�R�60ֈ���+v������W��F�%(�����GE�{���>��,��u��{�^�dl��I�mz����I�c���c�y
	�3�a���ޞ�z��z���:���i[��q �)�c.����'���ޡv�zT8L(��u�) C鷹�}��&��V�ʡ9SǦRQ��RAm��o�)����ffl�H��])���4��1���w#��zų��sT)�2�b��X��=��c�F<����lí?�:�s����6s�����kܭ�i���I�N���NgZm?u?nN�<)���^�����l��s���v�i�H{� �,���qCz�-4L���/�5�lԭ�C�͇v���J�8t\�SGj�a�]y$cݐ�i�&�QҚ���s8s5�y�hY���B�x����;���S���?��q-}߶k�k�b��g+�U׫.���y�8Ƃ�����o��9�1'��|�-:�7�щ19��ҹ4v��6Ah�}���<!o�l��dS���k��i褃Dj��%���m��H�a���F�1*����B��J�[���F����؊�ܐ�G�@�j��X`�!�C��a#���p��r�lR�Q8hQ�H-iF��e�#�ˬJ`��M��1�F�U(�#Pҵ��!bȔ@���-@ƨ�NId#��|"��ML@w�W��C�[r&��!��A�T����Ƞ042i�R�B�<Qp��I���K-���Jqm��M+c�� ��i�U�"U��^�K{k��d@���F��ᑯ�m���d4���[� ���%��<i�c�
�3
T$�Rez L@~{��H�,�A�q�p%��'�Ć&ۚ4���ӛ�k���V����	!H��������q$ ���\Ϩ��ԗO���{g��漟��}k�ӆ,��g,�!���{��~����kJ�^�бUmkUV֕�@���M�j�U���:�UU�U^��Z�TUU�*��b��ĳU{�r���k<��۽���TU^��Z�TUU�*���I�k���kf�SRl��5EQH!5J�����8���튾_+�j�V�U�U�;�Ɩ�I�i��-1��4�h4�hi�	1(i�#��\��Wj��*���j�W^*�V�U�}�<h$	��x�Q�$��%j��F��$�H�W����W�*���;�*�Ux��U�{�L�M�"�C�KR�h!�`3mSH�b��� '����s��^��ZUVحS�U_+�U�{��{�Zim������%5�Q�<ت��ڮ�W�.ꘪ�kJ��]��4x���՜��KQjb�d��M,h�����#[&��qu:~�d��	*R��KV����|~>���7�;�����a�`�U��w���������[�'a0c7�Brn1����a;9;9ّ�*\c23#�F3'��:Y��t��1%Ѣ,�����׬��^o�N�����`����!��=b�<�V��5唶�q!���/ʍ���[KP6ڵ�Ѐ�feѕPQ��R�+](����C��F�D��,�B��#TfD+[��4�d�*���gj�ƣ�*�ձ���)\4/,d��-��ӗD,K��f�p�;-�ֻYb�4�q�3.n(ۢKbQ)bl�f'A����\m�^K�)76[A��U`xUٽMX�ӲK$lp
>�[ItK���L��r7 �r��l�#�8U���׉�F�] �Y	�(hQ��*��)ܥF�l���B�(�$nƘ��C^k�ƅ��Z4mˋ �ٚ�-ma�cGA��U��ĺ�B`�]x�!"�;"�U�Z�8"��SM�+R>.��-��sKWwwwz֮�����I%���ޤ������@��{����	Io{��{��{���Ԡ��	4M���vL�T���9y�����/ͥ��&#���6�����,�<3nk�欪)-�|Zo�<�N�h�D�4G��mRn�n!�a��oG�����^DC.�!M�ܧ���<iRB'G�R���`�m%8=��:[mđ�G�Z2N�nΚ�хh(�V�TG���H�b����8�ꖆ����.��4z�E�pa�vF�D�Ș�U�K�9�Q�������.�l������D�#Mh��6"�b�åL�6�A.a�Ç)�PY;[\m��JթD�7�ZEY[��Nh(��$�,���V��e�S�o�I�&�{-L�%T���fj��<�l�:��.����QbUA�uH�*Nˍb�Q2fQ�7	.��A"�*�f3����9Zp�j��w����`�0���MI+@x^Nn����	!�6�o��RN7QL�M��pф�
3|dzc�ѡ�y�;��>b��!-��f8�5���d��TET@6����t�-���.�g�"�8a%(�m8��I�-4ɴ3/p��q
%Z��LK�mJ���Rqܭ�iU$�g	,(�'����!�Wś;�"�2������T�����دk4�p���F�! �X��!�BO���'��m8F$ nRrY�؛\7T���l��ѵ�H�Ʃ��V�S���=yx�_�&� ��0���N�
T.�h)r!,�&-R,�,FpVw��s��LZ��$�A2�3m��$�a��yh�4N=ᣤ������7��>��!���A����Ql�pᄖ<��Ƀ�3�3�x�~<IG�(��(�0v<�Ѣ,��n�p�|#�H��g��?#��ٲ,��!crA����7�_����ps0����N7M��A+ϗ陣s�W{�f�.����)	�_q5���(��6��������{�!����4W�W�����z@)�ۜ�[l� ��k��X []��[]�� �P��`��`���p�NF��Wd�!-� �m%hijNM���Iith�м5R�<��մƑ����u}cdJX��5 5ѦQ�� ���jb��JH8��D5:��"��k�\�D�qH%0�ڕ���= �B�j�B[�����hڥ�KLA�P)LF&���r6HC0!>.:錬m���fdb�����c5EQq-u@�ddi�F�"5�H������R/&0.�P��Z�Le+�L[��b���F�d�fg	�T�~�- Ɩժ����Np��1�J83��,,��-�m��l��kj
L!�mA�R���BQ�i��r*� i4�d V.�4zf�±��a,SK��DC"��c!�%�U �f�:Q�ߙ�="f��h���#��T"IP�cK�A�)�!4��m�D��0����
P������GF��-2����KyאЈ͍�H��1��c� ��A<oQ�"�i-5�����sn"C��vY��h>�l��7�f�M��B���#��4M,LK�ڒ-��>8A�m(,��J6�Q��,(��3�8m���p"4<��{��a�h�&r0X��&��U[x��;z�yYrf+<"ND��vdƃ��F�B�7�
��]in���-ȴ4q�z�J
h�KM�J�%^�f?8�I=��<�i�4���L��A�������0O�(�Ɔe(GG�DX�6���`�0�kK�ºD�T#҃<�ْ̆D�p�K����:��)����d�A��Ξ)�m��:}����]m�`š��ͭ�\LAu4AJZ5b8��K��4ܪ�!qBM5�а�6�b�FR(C[F�}D"Ap����Ha
	�֠K��0�aD���^""!q%k��i�5V��K]!u0k����]Pd'و�����-�����d�J�� m4J�SJ({�>D.��.vt��gHc4>2���|#
2^�`ꇃ�Q�3<!�F&����vEa89�����4l��g�^8x�p��H��0�a�`�#F���P�L?C�9�Q������\<��$R�R1�u�ڐ��ႛ�Iŝmy���{U�3�S����|����ה�x�<Eγ2����0�nagb��n">��O�d�0c0�{����/1t�w���LJvm�[�L�	1HD�!�?�V��iQD��TDk��]�]]�Z�;���&���X?\Y^R�4�.��#��s���.[l�m���[l�m����W ��j��W A(�,K]~� ��
�����誶�	�~�t���A��h���AAY&��M�YqdMK%Lj�	��c��DHl@	�@⟘�C<s3}^�b�s�f���M4��D��!��r�n�D�U��l�t�:ZP}#i��dAQ&Cf�(1��t�Iг��XM�3���-P[
MqFuP5��!f��[R�^TyH�y��"C��P�M)V�� ��M�!ڽ	J�*66�-qN�XR��(=Y!�t��=�	^THY�H4�#��Ʌ�\$��$�YF��:P-��8qŨF���FH=("�	J�$'j���!2��(���i\-�:P�C�t�PU��������;�sI�31p�q��7U�S&$�I���qZ����E����5��S�=i�C[6�"c�!yuq�Z:�C�{,"�!kk$&X�n`�d�<��D+��e��N����3A+I��F�DC�1l]{����Nݨ	��RV�qZ(/M�*uQ�7n�AMŽg�0m<N�b�S!Lk��0g	:Q�|R
k�N�΢Q��v5�Ճ<>��D�J��{n<i/!��m�	���%WY�w����h�l�8I&���6�����([16���1��	��h6�@e1ܣk:�A<���@�+�Xz|�T��J�9� �OI��2p����w����v@Z��b`��c���g�yXkPw�.�RCx&�#��D�Z�k ��8T)W� .�ǜ�Q0�W+�Vߌ�A�q-�. l8�����:l�K&�L�,q
*�Ě;þV�����PF����h�/Hޕ��P=����Q.b$u
	;�qG�[p��ഃ� :iY^R�Ae�� x6h�3C8A�X�>���G�<O���ÄI�]�K0�aD<4M!P�(�(� x3!���,�6F��p�'�#�H��2�����pѲ`�,ra3#��yM���H����d?f?�w;�Ŭǫ;����E��{��Aջ��FM�~�7�f����@~�����p[l�[m�E�ܤm�H�۔�m�H�۔����0.�8D7������p|�4�&[M�}VWx��&�^�.���]RR�xf�$=�Å+V�lc��ވD�e�N�6I�H,,��"Pƕ.d����G O����IB�����x��h3H�XuSUa��z=�F����.���8�<kō���dqpᆍ�A��6��qҪb-����DV�q�Z)m

��3u�t`x/K$�ZX�zDK.1�[��ha=eu:Keh˰��Ah�
ES�zb6�
݊�÷�R\�Ea7�mVYђl�H4]�;�[�I	Q�:0�e�!6�sjNA�Y۠�h��;a66�.f���Ë�ì�GIF��p(�B��0�GJ �Y���4
Uv�n��G���1��t��<�b{Z0ֹs-�1�f(���7)�#F.$�B� 7���	��2��f4x����4����N�e0���-�<PuX�ͬ\ءrL-�Ѣ�[[��u�%Ci��${�	P���'��b
< C�`�N!=��i%�²��b�IťȂc�ܩ�F���1�^����(h�
�&���49�d��ln	�<[Z!Yih�=(�I��Ies�i�LX3�c�hٴz��:��ÇN�Q��bydz*Js�֔]:�If��J	P:��7�[S��Ԍ�g�!��cg�QÈ�]�h��b��nZ-��m�w1��0�X�a�T�������5�t�D�mh�ȵ�����Ұ��N#%��Z��/���%tvJRX�h���/�XG:Q�:sٙ��cwS)�3�H�M���H�GN�����Ҵ�i��\��(�/f��y����b-�(���'��"��Q�Ign�t����L��8<����	��	�!����vx�x�0x�œF�(e"�#@�f����h�F7�	Xx�|a���<<A����{#`�0�tA���0�C��YD��� U�?�O�����t�>���R�J��E�&�⸄햘W%n�(Wm�31�I�︹ӡ�Z��q��.�&Z���kJ��(��D�P`�k*=9�p�ܱ��]�m9�ߍb�q:$���Zi�L�w�,Y�ƈ�60�L&*��'�ܾ��i��m��ym��m��m��m��(b��0e��0\�Ƌq���!�����835k�I�Z�4�R�J���#4�K+X��M�1s�p;�v�A� �E#��H�^I�D7�!��ܳ�+m�d�@����3�	)&�3���\�T�YGL}Gy��aTQ�4v�Sib(�$�m��f5��x�Z�J�#��4P����;0ۓB:.��IY�yI|PJ!5%�/s�'�ǳ��4qm5�b�ו�|�7l�f��-�\5Ʈ��1�D�FaH�v�l-�'�3�d�!�ƄJ�4�9�qR5&��d�Ø�A�\8���8���k�*��y.΢7Zs�h��E�6�:h���E����h��i�~���sUTD�-�sJh�W4AC���\mZ&qZc٣�BR{4�$�Xl�FB���!$�a%�B�Gb�2�v��plD���M�z&źV��g.tER�rS�������e�Co�zu!�����D��jMoc6�b�"S�8Q�[�(�(k	�m���Z:�g�fѣ:t�����z\�'�V���0�quJ%RA���=.(�P��P����!�
� �4AȒ�Aj��㤛��~�lF�"[ �H8�!1҃kG�1C�������m:4��'��G�(�Ác�˱(�h�үY�7�8�6å����:�6A.��[K�_L8-��f�I�lT����Fl�%���>a�f�46}$����s�E926���c�6�1<o�I���؂H�r	)Z�E
�'#�
�x�5�D�Ѥ��o�p�c�^(�4��a�-P2��$鏄6�sCp�n"%x�SDxn��8I��Z�ƈ#SU�S+B8zGj�G�5H�_��kNMi�F��h��_Y����J2ԑ��Cm����4i]�F�.l��
6t��@�lv��8�#����a�0Ä�ht`A�f&�N	(�5���
0�ǈ���F���=#���{<I��xx����?��ㄛ���'S�������>��� ���o�y��z���8������6��g���Ո�|(x�_Yw-��m��)��m��m��m��m�"�P0�3�pL�������(F͏�Cr��H�$��o��h´q��q�ᥴZ�taV�5H��p�M�˶�9RL�-i�o�7�J�A�-(Xn���yT�F��T�����]��T�Y��t��)u55�h�qZ���
$�q,P�q��F�[v\p&<c�L�Emb���{ZO�65���p�o[�%��Mm���ޖ#��ůGBXފ:�ۥ�`Q͘��]LՏkT�&k�u����G'H�f�#�5F�$�p,Ō툢|έ�Hc��LGQ���=��N���DiVY�a�,�7�
�:�jո�2����ږ���d�PXQdrH�S#Q7���4h�j��Ν�����|�1�� 	��2�ke�&R�u����a�b�l�d�
<u��K۵�+fT�d���"Vq��h��fP���J����4iזԦR�G����P0;����<IH�q/���e�1��4Ey��ZN0�f����U
�t�Z��Ҹ��%)#5U	n֎�%��J!F�#E"�g�>��
��E��Q�F����ލu=׏Q��Q�1�C��h�d��Y�0kh�R�����ҥ�DL�}!� R��V��fq�M8�Z!pkʍ(�Z�$�F&I'B����n]:��k\�Vti]�����uH������aQ2���6u-�( ��� �����84wE	���ݭa҃�F�0�d��:�PB:����t��G`�1�zqB�1�#��1O8�qi_#�i�R�qEB���!�Gt�I���1�3C��p>��aF#/æ�Ɂ1�p�N2]M���(���4n^���l�c�Ğ:F��x~����0{6z^���A'�$����{�{�l��� �0����V/��Ix���Ai.T��3�CJI 4�
H�d"��	S��׸����H�*(���0w���6|��b�x�	�2����û��13�X3�}jU�yL{��y�LP��)绛�S���gP�M�Y�-��\O���t�XQ�c���oK�i�8����sv���,�MG�d%r(���/Mb�G2lӫ�4?N"I�/ϋ�~���m��m�ۖ�e��e��m��QD ����r� Ùqx�ֹ�u�1j	0�6�
XחM1�#���H�6Z��[l�MKm8��>$�5�;�{�{~��0Ә�C%F�	EǷw�������!����\F��9��*7OÍ%��I���q��a�;$��V,[^]C�gL6
[��u0P�,)>��)Y�t;������������"I"
��xF'��\���Z,�ӧ��ve7�b��;]S��r���d97�L��.��{VJk���&D��-�m�m"�(�AaFj}UD`5��R��66�ъ�u+P��׼��4!f֔huZ�Vqb 5|F-��8x���i�7���os;�w�ͷr��w��c�rf�v�X��J$Y+�ߕ���.=P5�f�H�c:�ړ(�<��p�H�|�������o�J�'����V7l�4���T�MF�������h��5���pǐm6�D'H:�lꕳh�E/	Q��(�h9����PZy��Ҭ6BX�u��%�|�~�t"5�r�z�y6��-��#J����x�e:�F�,�h"�F6�-�ͽ��.#Q Tw��!�:�m�فK��Dmx�Z����aGtwF)�m�x�G�wۓ������ ٰ�Ӭ!��'�52��'r
��_���1 C5�F>>� �9������ ��'-�(�wu�֠��/l�><�U�'m��*����g:xjy���-�<D�a�kd�;KF�4Q�����4x������C}d��'`6���1�*xNl�8�is^g��L��g��۔@AH�*8IH��5�R��2.zk��m��gF3�1�xG�4a<0�0�L���a�	������(x8F��#cٲ<p�����G�`������0|6G����t3ĐadP��(�~�O#T�ߘ7��U�� W���g=W�v��ݧ0{w�b���k������J�f�gaY�[�G[�J��fm��E��m��m��m��m�ܶ�� �3�� n��5f�J!kT�/�;M�p�ԥ��m*6�Lp�5�p��8m#u�8��#����AD4��frJ��CU��%�AOonfe�c�aK���Q����^R�K\��v���HI0v��x!@�~|�E{�z�[�ê�y-�B4Z����0�lD�)�#Qy'$m��i���C���pY9��[D"�Zm7{��-#��|>
�;J��ILiuq.#KJ���M�t��s��rz	t��FJ:����X��.p�,�h��Z�c���X��"��-������WQܭ2�f��)�6Xp.�-R��7��`�MF����)VF�9=�������"�IAm�Kt�߆���>2���0�a}��H�u/%Ը��d6���x�P����j��9�Q���[5�J'�����0sX��-m����Und�1`�2c�E��U(F�����k����$���z��861�cƏ�D�iF#�<��>x��Sݣ���$j��È���1	���N��LE"n2�2s��>���(�i��J��z�Q҈m�c��Q�q�l��iix�qWolz�i�pڃ���*��سp\
��٣�Xt*w<rK��[�MIͭRzW�]T��i���p�Ds�k���M��&
�YťP�;���D�ΐA���a�M���cf��it�4E#�:B�;+jx�6SM̑xxȨ&&Sp��\?#��H����*��\FѤk�:\�W��6tp�i�X�l�?$�2�'����	����0� ���M�DE��#(�� z� �4x�����<>��0x?#����>#��B�$ܑ��G��/H���^�@�����S$�(1���z��0�U��s��˽��|�ǳooI�΂5�V�!9�2h*�}=�;��z{�Й�3txt{U��zR��3	k& �*��!qbE�xI�0�-7I(���]*���oV�/P�׹5�x=��������
8�y�Mqʁ�R����NɊX���*��HWjE���UV*�6'��?3����m��m��m��m��m��e��m�!F�~� x����
H�	MhM���zq��ݐt)n���MJ����]��ji�B�k�F*��.���%�F�Q���;0ż3uͶ�`�a�� fx����*2�Q�AE&�U������#&�[����GI��k���Nբ�$'>'IY��KT���(kM�g�ť~��s�(�z�U8��C���=L�-�m��#��:cy�Q��W�4�R��t�i&��tgH:A�ad���Kx�4f�P@RΨ[[�udg��j�����g�3����G���4k���{o�GPױ.!��'G� �aj���]��<^*7k~g�Y3L��D�L��ytZ�:.��\[L���i��W�Ό�yI�ĐY��ߗrE���"Up#3#�٘��8�j�V;�$�l*#y�dYrdOV�^)3���=i4��K�wE�e��6=��u��D��qE9�Nv��E&Y&�,�Y��Bs��Ki�<4��U��N4.얫 ��l�p[U'��3j"�O�7�QG��I2�ɂY�� �xo!xk�D�ȏ.�D,R����˂��4#�Z7�k�E�&���^�񸥩^Z��A�Ag���h�޸����-4��D���(X�Z����W"��Z�8���63��ꥨ��m�4t���n�<�I��-ۘ3�	�e�Q��[U�����ԏ�n8�:�j�j���3��#xy���Z�iq@t�Je�b���$��刔\��έ��wh׮�و��f$��Z\캨���P�.��9�ymJ��+X�e*�)gr�yDQU5D
�W�I�uq�$�[Pt�GFt��A�F|��\��ndga�1�t�C(��J:QGFYe�a��6a�:açL0�:l�fat��˸��Π�I�˕��O].>������N���:��M>�ed�޳����ԍ&��L��p{{��dުn���2�w{�Y��ɼ���2���c�L��-���m��m��m��m��m��m��o�� .�����2�hڟ)R��p�1�J" �:��_�ߌ6�H]1M#���Y�Ɣ�#�L4IaFm�r}�ln�#j�|���W�Ȉ�!�ȂB�+�{Z��V��t��U�F�\XW�p��d�J�����v�����%��[t�Q��,I�4)ר�ko$�ID;Ge=�SdD����V��ﴹp���a�ACr�����uC�sM�8I'��S��֑I���0Y��޸�gW���8p@���Śm���O}�"QkI�Y'B��f��#H��w�15p����i����)�8l�MZ6t�,�d�D����E�(���k1���E�to:��[�]�G%�r�e���#�j��ݛ���cd����.�i�hrB���;���$�IAD�Q�Q'*��8�]őyJZ�c��&���̎�D��K!$�/n.g>vc�&"��qJ����{�p^�������l���[A,0�5�ukp/wȪzd�Ň
:IADS����!_Q�8���#��b!�8�%��TDt�l��ӂ�*����<�%s�X�y�6�q�m��:��#G��$�Q���:s��lo@G����*���w���fS�v͘�F�G�����6�W�u:�\�gO$�� �4�8��J�¦V1�F�z�3*_Ə����6������\6qM����=�AZ���]�9Mc~����u�Z�g�ܖ�v�
�����m���1$2�~�|󽯥�N+t�U��e�lAɲI`����� J��(N��n�)��Jsi"�6��AjKBԵ
ol�gl&$��7ق�K!JE,IK
P��))�&"R���)aJ��J��)aLRb���*JX���%,JY
X)�LK)��H�����0Y
Y%,E3I��RR�R�)d��R�)RR�K0��$�bR��
R)B�%,��
Y%3I�R�)�*)d����)D�)1$�JX��J����)bR�LRbIJ�(�����%,���JY%
R��`��)E*���݃\�-쪦,��KKKal�Jb,����)�aKH�,��iTT��E"�&��3(YIb�#B�)1(��KJ��&s�eKJ��RU-�T�RX��Z+83C*YER�T�K1R0���,QE�m�KV�Z��2��RYbb�bQ,Q���F���,P��YEQe*��J����*QeK�X�*UYJ�R�KT�E�=�jҩ���V*�X��%���(���e(�H�E�E�K*Y\(bT��T�V*J��,T�P�R�K�,R�b�b��eK,[+�1*YE�-R���E�ʲ��Z-K�RʑeK*�YP��U,�(��*)eK�IbSm����RXRT��RP��)*JK"�Ȥ�RT���Ib�R�R�R��R�J��%)��JJT��R���J\��aR�T��)aK
X�X��)d��Ko�(ˢ�(詛��e0�7�7kP�k	@�(A�Rо�	�*�*IUQ�I��b1��1����q��p�������c�����?��{Z��ݬp<�ǆ����U|g�6��C��M84���W7�a��{����O�ou2��˫Mu�z��I���˛&�|�Ť������9l�Ǘ�e;x����0�$?�9�ރ��{�xZ��������"OЧ"wQK	?8�K*�YS��O�O*}W��G�u�<����Xđ�̞����N����RdÓ��g��첼N.��^�G���D�B���O�,g<?��R��;>e���74Mq��ިhN���6ZL�B�e���8#���D"(��M  .�
������Ƀ�z������̚ƕ��Օe���{��O���j��9"$VZ�/ա2Cb�!L�#C�̑;,�b,��,��Y1D��LTC"F��n�j����M���d�ɤ�<_�V�Rl�<��^�Jh�2Xr,�@�D��U�HKJ�%�TI#��R$LR�.^G��z�zS���J��'��o�'�������jq�l��,|,�KS^Q&�O��:�C'�t74��,{����8����,%����y��+s0�L>���;Ѻ|I���{�ԍ���9���:7>vy��`�4�=���sV���OR(�et;c��:�g�G�o���7����ܞh�Ht�
���,%%��O/���%+�sc�ɸ������G��܌1dU{{�؈�!U��	��O�E�w�����G���2;�5G���Ԛ�8j�ä���2�y:p�"MSX�y�[�ڜ�+n&Y��NXJ4r��H`�����=�blI�#x�Y8�Jh��Lb0��1$�1���8#X�R��)��)%�lKH���e�����#��$0FQ����m�|Yx�{(/��4����i�m�T����=z��C�i��o��n�#���d�N����2�������	}/�`���O�8'�=G��1`h��Ƒ_S��i�?��I��� ��h�6vvS��U/�J�z~$�S�	�CX���i������:O����|��H�D�m��9�C|Yd��E��v��M5��K5[V�цP�_/4��:�ߧ�Ň����'O#�,�QI�š9��7�M�٫��87�T�F��9��OV��	���v��Ƒ����a֎��1&CS�Lc�v'eE��i���n���cω=-e�^ݱ�ũ4�0�~%�j'�>g����ÄvG�B�"M	Rg�4�@�yQ�˓"<"��zo�Q�℉:ϋ��6��9�g���w��͇����<b�^���4�J��z��i������H�
nv�