BZh91AY&SY��Q���_�Rq���b� ����bI��| B*���D�Q����RP�(TAR"���TI*TA*
)D��$HAB��T(�J��*�TQPP��4�	ET�J�P�DBEIU*�( �%�A*U"*(�"�%$����*�@�HEBT*J��y���OQ�Q%����Dc5)%�AX�JH�
TB	((�"�I��RR��(QPATD��*	!$��   �|�����ҋY�Y�����m[kmM"�V�ֶU5JM����P���Mi�VaU��յ���*�k"¢�RJ*��RE*�p   �j���3�
��T @�  l7@4 J` h5]� ��0 -�Z��@Fj� ��R��JH�
0   -nh  v  Җ�M 4��C�3p  �w  �� � �M݀ �q��:� .W�y��Ҁ	�U*�H!*��%   =��ٴ��@ 	�w �����z0��(8���@rU�� d��  n{�@�W}��
G�%(TJ��Q
�)�  �q��E,�����ҹƥA�	�� 4��\�� ,� �y�W�P��k� (6U�R(�;��Ȃ"I I*�*�U	p  3�t(� (v�M #  
L��uUSl�6���Z 1�$
 �;�  �IR
�(HB�"�   ����L  �� P��  ,��
�e  5��� �
 �� b�@�PUT(U )PDK�  8�+ 45iK�5X � ����@4L4 6���j j����H��JUH	J�K�  �  ��)� ɀC4F�  6,45�1�  6)� Kj����JJ�P�HT�K�  �  �X 1j ��F� ( F� f� 4Q�0(�,5��4c@4��P� O�2�@ �*R�L��a0M4�d��0��{FR���ddha�M �4( #Q��	�h"= �Fѵ=B)� ��(����M2h�44�=I�ު�Ji�2=@  44���ID��(  @   �G�����*��k��癜�<��֚\kt��6�f��V���Ζ�=�UQ\�QTW��A�-�PT���*���TW��]=�l��������UDpQE`~ԒI&=M�EQ_���O�?��`�d8"�
�=5��J~w��K�H�(�Ɋъ��[1[1[0[gm�{;od����d�{&d7����=������;��6�q��ogm�{8�ɷ���og��vq��gm�{8�����=�vL{ v����{&ǳ��@=�og�m�Y6�v�����v���� �{&���od��{ �7�m�����,�d��=���0{&ǳ��@=�og�g8�ɷ�m��q��od���{&dÝ����{&���������p9��=�c�6=��c{;k>�� ��ogla�����{8�d�c�0�=�c��`; =���%��%��%���
4`+f f
+V )f*�f`�pl��`�od���1�{;d6���{&�d ǲ����{ ,��ɰc�0`������0`�U@�@��@��@��,�E,�,�P,�E,�,�D,�E,�T,�9��M�ɰ��`�v0b*b��b�` b�gbɍ���� vv0�TK1U0l�E�F��@�U[0Q�EK0d��� ���{& =�`d�m�c{8�ɷ��7��og�{;ogm��{&�ɷ�m���ǳ��vݝ�����ogm��od۳�Y6�v����ǲaɷ���@=�od��6�pY�v=�����ɏg���C{&��og���{>�Ð�ɷ���C{&��7��fY�bG�:�䖎W��cx�:�γlN���Lsf]��	�ӏCLf��(V|Ѫ]�O�%���#���եw��?me���oPXZ�_�I���#�|ZT� ���h:��&�e�wW��X�lP�c����%Uf:Fɚ��2�ʖ�(i�w��V�]�8�=
ӯ�^m[�mS{��m ]�����G7nM���ū,���nYz15Vڼ�i[�Md}-��[�&aئ����m��ʧC�j"�Q�0l\5r�%l�X3C�X��Kݨł�j{L��w[t�)*▕��"tT�fX�H�ۖ��Jbp�.b-ʫ��ZBv�(=Sa�Q�`��)}^�բb�����B��U���� M���h��e� � d�K4X�;������̶VɎ���o�ř�9���j����]-T�M��j�c�bQ6�Ôpe['f]�'W�(M�M�T��O ��wM���\�U&^�tv���w�"#7LEi�֪��-=ӱk��j{[���6��N�M���3i�8p�9x��&:�xh`*�uy���F�a����K#�a���+5۪X�.LΉ
�2��h��a�	���ZsP��P�b�Z�^Pgi�T� Õ��~H.����ǗV�"1i�b���_h4��ZD�C2�6�ݬ$�t�f5��9�`f�vw5pU�/n�B�Q
YX7n�DR�ܟ��J�K���
��-|Eڑ�ؽ�wV��d���[J\��pB�n@W���r�un��L�W&���X6܎��{���t���I[%Xw3P��m3vL;HnL��Lъi��1�wR��إYff�t��r��u�t)#qMN%#�a9J�g,G�h5e�wvۖ�X`�;ǩ�L�^�)-����a1c+)�e��U�HN��-j�������+�N�wi�[��iˈJ�v��� mj)
Y�t��$j����//hۦvl�f$i��:�Y�:�y�&�%�+��W���,�)�|6�<S �����x�9�, �P�a�f;���rFpFv���E��R��sA@;�ʇl��)Z�h86�HQ�����!�6mZ�܅Bj*b�l��[N���S	�<��p<,:M�H}E`�-u�Gܵ����7n�p� V6n#Ժxl]$�7Z�,.|�A��o�(Y�!���M�E��p�&X��NF��<���Q����v�P�όx�[�%�AL��1�g.Pְƶ��i���B�j���n�x^�&5�\Gc%��E֘j4��jv���(�T�KV��	ĉ@��{N�pR�e-���{�I�.���� S��i8�AZv��"D� .oĳO3Y� z��%h:��0�7h����f�\4p;�0X!+XYe�yv@N�����}�'y!ҭaZ�9��y��6�	�Q=(I	�V�W1V�u�n�A&�䵁�6#��x(�F[n*T�&��4%Г.�N6����ݢ����mA��-�Z��m��@�h�%��M���˧k)S��%IOn������*H��n�G�d�V�0p���ut�ܧV���Ӳ��.�,�-�v�F��B�4 {L�J�]���n��z�1Ky�>pA��G�zjvfmA�-]���
�NԘ0j�op�e,׫*�)�+��U��[�[��h4q�cں�̨sXq��P�ZU=;�*&�8ҧ4��ReZDa�Y��e��&����M�n�Ȯ�i&�a��(G�2#y�,b9��v�f�^۽JL'C�����R�P�&�Ҧ �kv��E�$�lw�-�-��i����=�j1f�wo����i;ʇ7 �j�2�c Hr*�@�GYZ���n�Y-� Uš�zD �M�z��Z��!PP�]�W�������ĩ�E勸Jן<+s	�E� ��6. �$�[@��ef��H�,��wa*V�AY5�zq��;�������M�x̲#���S�r�-9{0��	�庒�V��Z��5�L+\�K#����9���:ɻ�6 �&[�R���6�ꖾ�p���J5�kn�L5�4��t��� �s*�G�P�jZ�3o֭85�F<��@����72�e��ҤqR!���Xr3�!�4���	`^krIF���Q]�5�'�����[��դ�Dּ���V-�@)��{�)&���ͳ�5�Z�ۡrm�&6��4�*��)�~JH-�$Gk".�w[F�ƙ��]��T�� �(ZĐ��E/��'�R��ː�G!���o�E[4 ��0�v�Ol�YYB�˸7e�Ս���C*Ŧ����CSu��-��Xi�Jɡv��yM��"m(�0ڴ.XCS�Q��F�W���Le �ْ^����m7[��b�S	��<-)j�p�J6\�r�d6���i�zX�Kon��zN2��ҵ�I���8�^����T s ),��K�Y��]dJ2\u�j�6V�kh���ASj*��TwmS�ݻ�/q�0m�Ow���_�z�pՄ�3W��B�&%�
OC�D��M�eI�)M���	 x����QG��ǴU���Y&4�2�Y��ѵ6�Rǰh��Dixt�m:PbD�]���2�V+us_Ąn�W�"���[ES:X�J� M4%^���" �i�Y{u��7j-��kA{.�n-�6�K��[�nYD� ��jaMKT�`K���v��(�HrS�v�52�#�ۑS�0-ː��M٬�B�J�f�P2-�>!��@�q�Vb�`�2�Ղv�]��H7P��2Q�b�])p�@Pm���;��V�]^�/&�Ӏf⦒nB)�7osB���BՕtou�j9N�WzTTV��2a݂���Y�7@KY4�4�Z֧����G�Q��b�@&��n�K�i�\�RK[���\MiM���&J�Y��K��1Lmӹ�3�kM͚��Պ]b;X��ʇS%7���b���7YsUGx�lBI��hV�<Sa�um���IaB9ݧy�����
/N��F|,	&��ܭtd�M��*�̸c�1e-�N�ff&"�N��T��D$��*�OD�ɬ�r:ؖu���YoDE'��4ʷ��bWy�U줭C�i�AVզu��$H�����K�B2�ܖ�B��չ@
��1z�.���լ���.�p��ז�7b�/V)�G&�F�"��&ֻ�E�@�۬�КJ���XYz	ŉ)�`&䷸��f��Z�!#u�*9��L��Z�4��yV�B�1eb֬V���P$Q͛Q���ΑW^�����c\B�����ue]�&���f7 1�����6�B�e�	�$��2$���Igx,'Sɒ,���D]@r��,V�guP�"^c@��=GVլS����:��0IQ�c#d#�����= j�=�{[ئ[�X�NлI�B0,�WZI���f�Z�R�^V)xB6�����5�u�m����wqD�6vL��L�V����l�w,�2Q�.�H=F�Z��/,!jG�բ�Ѵ-��ݥ=�1�zp,J�+8v�&5�,����
�5n�w��ޔۤ�3[��B4`3��A�[�Sh�Z�h;t2�C/-�ķq�yz�r��yR��Ń(y)���8S�-�������J� A�d$,��Zܹ��"����͂��(�n��v��� g3ۚ����AV�L{{��O �"��� �D�z~Z��hǱ��m��3�V�Dv�U��Iޙ�C�L�4���EJĩ�u�ۈ
�u��xVv�0=��(�A겆PK5Kݭ�b���;b�%WH5H�&���2d����W 5�Эݴ�¤knY1�.�VR�e��B����ւ����V��K�M�t���+ܬ��̲�-:�c� ֊��dm�oN�5(sUK/�/IV��Od�h,��8�;�]%u��*�O$��ڵ�w lm�K�5�҅�rU�{`66�����	����d�8;�*����Q<�mY��_$6k�h7�]�8�G� �F��h4�H!`X5(K6
ӳ��+.��Z؇*�m8�Ŕ�^�*�ˣj�i���`������+V*3,�w{�<�t�D��RMb駈k�;j:�M�������S.Rr�Ņ3P��K�B]e�-��ϥ��`ؘ�X�
Zܵ�"(\�-ȥG�Y��h�X��p��vG�6�gSZL���7LS�7A�ƞʸ�b��6!���Z��Fr�˰%:�C��4h޶��w��f4�ZРb1y�ƅ����%y�D��Z*�ЫU�ۡ�"y��	R�&��[Q����1bmI86�7�.�#9W�� 9I�À�vwYI�	�RO�p�8�fkR�V�Bi�$�(��y)�v�ϴ�Z����՗-�Ҕ1t�[u
Lb�B�5�;�ٴd ,`�#X�)eW�V���n�EX�ϣ;iA`1a���jm,��� �7+4j�Զ��x靧��mZ���=��	7!Y f���
�C]6��ZN�A���j�WX�U#S.؅a.d�M�&�=3֑��$��%�9r��ӣ(${�[k���mnL��փ�["��7d6�Ƶ�΀hi����R�5ô�T��{�RPK��⭡V%cT�;Q�y�j��ĺ���6��8#6��mTJ������+R�ŕ��e]���w�Y�b#�5n ��A��&�Yt��+*#��X@J��Y-��_ݹ&$Ԥg$�.��x#(eef��1<��f1*n��w���p;�Q�G[Wi�������$���c��A#Q�7��nШ����c��'��u>����h�+-4^[T{nt�S��S:PR�Uc�qʰ���2��rjm�Q�S�r�)2�&��r@��g���ۼ�.л�6<�H|s\����Qɸ݂=B�T���X5e���*�֌�J-F���!��B�2��`�Zz��V11A��m�Y0�����2�{y)�����jVS;�&�-v�k F�:��5z-�7�	,��d*)(��ਚu�'����1U�b�)ww2� �*j �L(�X QZ��6�z7s]Ja�K6�E�����q],� �6�V\B��[�9��`(p*x���n��f�S>���F�ד`K]������wB)�;[X�"`����B�L�i[�	L�henZ/F���+m\	rR�{��v�	pTy�*�b�,�Ɯ�����Sn-�mJ��&��.�8>��^��[Iѽ�� N��� �pJ�YMLK4��� r�ۻ0�ۄ^��c�^MQ��Y�Հ���.��)�nQ�k��f��a�M���,�s�խ�f��n��`tv�N�뤲�+E
�K��m�(:�͓���n�*�6�6�+u��{���QqJ4�͔[;):��:�����n R�3Y��Ҥ,P36n�t��U��K�q�{��ݫҳ(�"b|����%^�x��1JnAT�쳶*S��j +*�^ca�ZD]���yx[ߍ�Y��I�0\Pۦv��s5�� ���ڋY�&���8��N��7Qv�Ƚv�]a0�X�b����:�@���*�ѫ��0�Z��E�eYĝöҐ�0Zk���t�^Se�;���Y����E�]��j��ᤩ!p�G̩���3�w���I
HҘ�#�,���v������˽�(�#��-X�łPw�e$�;��rw�J�ؔ�;�oc���5��=��Y�U��bu�S�1K��F�Yz1X)b���wy��N�#P �ZD�7�a]�a���n$-��[&D�����lD����ʸ�A�>���lYX5mb@}&k��.���S[fe�d-g�njڸR�J�Ԋ�3#7�wV��ʎ�&�y J���ֶ�1K!m��_�l�ɀZaI�f<��������P��Y!���7�K-�ʼB|�cz�7�l;2Ckk��YnaqU��=�p%�n�-śNűxa͸�%�˕n�3S�fMX��-m�p*�ֶE���y�yk� N�1���Z�@�O(E��mKW.X�)�IZ�3��9��ʂ�5V���7

P�5gv3e�b� �r�U���SV��tB�&IAVqh�W[�"��t1d��ZX��U-*AO]�hEv�f/�%�9�6�	�ǀB��7h��`�b��`�"Re��r�K��0����A�9WzVh틴JJ�Cul�ֱ%"���u�KlMڸ��bĉx�&����q�
{��5f��f��C����V����l�-R5v.efm�[�;� ��ͅe2�(�v/1�1�֫q�2�%Z�:t�X$V��n��. ��d}��(M��ƞ,O�Ӭ�d�,�I�u�]�ӭ�s�.����V<�q}h��On���Us!�Zr�N�)e+��=wn6���E�LAR^:��-�'.f����	�FrD��̂��B�o3[a�u������E�ea�*�R�M����^Z���L�3]���c �G��"Um��Im]Y�~(Y�u�Q�tUaj�Ym.:�	0X����s�����k�L��@�u��DOX6�ޛA.��IY�}�i���������f=[�H"���fq��'d�qҪR���˹�d���w�TŨ�!W����e��[%P�z��y��ótʧ��3m��$�̢j�Tl�(*zjT�t���;�)�b��;B�UnL�t����;��:�]�͸�ݺA�KQT�v�"�hw�.�b1R�'�e�	�oq�h�4��
-⡱ZJA��:!��12���pη2�L�U4�Ɲ�V���8r(��:��� Tv��%���u�b\�Cu&U�ٮ�S��wuwN�ȕE�;��Z�ǅ���(><� O2T ����ko�`�K�w�a*7SFY
�j�K[O>�2,�)n�{�n�W3>~��i��=j�`����J���r�"<z�~Ic����Χu�WDgk���M�\`�h�9տ;�r�ځ���g�m,���]L��s���+��3�8�U�]R3�N�)ە����|�>�=���iN[D@E�����'N�b��7�x��z���'Lj�ԋ���#��@Z�yz�S.;�כ��/z�vB1H�� �!1�9�˫y�ʶɱ[ô�V�\.��wH�:��3�sBދw��KV-��Vu>JKuq�ZpJ���[b��8}�����V�-�L�����k�,�2�);%�}N�x�.Kz�IY^����򒬤ܮڦ�*i�G��+�t�f.��
5������֬œi��&��rS�OP��'E�.�ڳ���X�v㈀T�'״�n���f�]Z� �Ν-j�����cG�^����}�򭑚�.̉`�NQ{j�ܼ2#�B�^]N2u53�ɠ-k�u�]Ckfr
�k$U{�����h�]u����`��j�e�M+W�b>��3��
�*�k��Gv�u΍9��w���C���7�Y��S4��bvy�a�	l��ev��A���	�yI�R�u>�.���EM��p���8M\�`���0I�>xr�u�Vk�&S��3#ӕ��k����:zl����է�sOq0�EZ�.��[�����x�2s,���}4XZ�c��J_: �+��lt���ۚjh����}�,��4⼉�Y��'Jt�ik�6L����Y��y]Bb��X>�de�]J�\�P�nZ�܊wv�B�#3O-��x��2��L"﷣�t>ԫ�m���b��>u=�5G���B���|��xb�5��u7:�?�oU�(�v*�r��Pg n,���
�ŦwJ�cp}�SGQ���u�(���Ck����jV��Rr�p�;wrl�^�4E�A7���X�VRݰ5驩�֞���Y<_�L@����zk�i�u��ҭ^2��U��o��L�njLL��WZ�r[���Qt��[�3���4-���S��xR�̨|`𥍻��
[K�Tb�,gbU��[�+�d�\�g5�)T����g�裱�Y����(����sj&�-���ƌ�LIS0%�{5@�%�>�pY�z!�ֳ��$��B��N��ק�c��@�p���}z����t��0|4�MYn��p���]���4WN�FͶ/4�1tX;�'�.^t�/�]t�Xt5��1�g�X��>
� e��ͬ��f*���$�9���r�kPŗ��Mn��MҬJ>+X̬�Z�>ط�z��+a����K;�Z�����a�~Ҵlٞ�����)Xދ_}�&�J�q.��=�U}q�4���)Ŭ#����t�e+�o_s�/�PNn�;�3G�K�p�}��h�\��v��sK�yB�{��cAUu���%!�v��zK"v�#6NW�c��%1�Ŗ3i�:�a�FY��n������j��vQU�b�T�!M��g��פq�n���H��4s��C3;�P�
T��N�6پ���net�T���kI]'V��C�u���h�C!u��2
uH��C�׌G��ѫׁ43fYi�O��t��;��
�Uץ���Ɛ{¶G��Zlj��Y�*Z�I�9��!��+�K ��*�R���:�K�}�WZ2�c5w9$/�44�ˢ5�*U��-�f�>Y.��].�nA��H�6�"	�hAɇH��3�_�T���seg^^�b��!W�-�!��I��x��rs�]�i�����6[8z1�����M�ԋlS�W���w��@�vǆ�5��ٷ�p�cr���]�Y��W�KN3Ebn�s�z8�ꊺw+��Xf�����_f��\���>��t�o=tu͊�5�s��j��V�X���]�7�8��A�BfW,Ćr|��.lISIh������@�[�WXʳK/����}i֞����:�{�t��֥So��Z��8�Gf
��S�Js�J7�E/�z"�p�2텰b�Z:�!B��C���������X�J�2���V��|�oG;��	��2�ǁDh���s4zQ�(�
�8`�EWi��d㥨�q��F����ulV3��t�a���.���rĎ�8��2؃*늌̢�Yj��J�L��hk�³����}M���3��� �Qϸ=���m���ؠ�;�����J��/3�R����I1es�nD�$�N�v�hV���eړ����|��*A�G�btU��Z��sȾ��IX�o,z\���ܭ9��B�+F1��$�����/�m��rWs}�>&�|�=<�1�Z5�sWo)���Z�W��5�*�X��Ò�f��˖>�caY���K�W�u���6��/7L�c�muJ�b;1'���e�.W�<.����"�Z�S�UM�p7�qǓl�^�N���ꏥZ�(,�#�vM]���+�n��k�����[aE����v��K��k�5H֎nɱi�6�VYG��V>��<�f��r��#�7��!E.���,�a{��T{�_+�5�5�b�Vڕ64�.9�X��8{�piJ�/%���绔U7%>��u��c\�ڰ�|*rھ����cӶ�/�s:lj�A�m�R�nb}���khJY��% �r7��ԙV�=��4ڀQF1z_(uͮ
������/�^�������W�eJK=��F���{����h�y�M�k�5\n�d+�+����J�oq�*\�P�\�h��F�䵭y�9�{b��J��k�%���Y�g�f���@e@25���Zݤ�����s�ѥ�C[P�Z�5.Mv�������֡c�YQ�2{�c��0嫙Sp��wR��k�F�J���͡q��_wTI�k�Z5v̇/[��D:_i�����B��2�cB!ub:�<&�*�Fo�9A��"��v�:oJ�|�邱�hg[�mg��X�30�]���z_P\�R�%@m�#��bY:�-tq0D�L�uf������rHC&
���� R�iI��웒�`���>��y�v͇L�o�b��ƴ�"7*�+��K2#�v_K(�l�U�X%ݥ���4_�v�4����
M��/�����w(w��J�mDRV��A,7u�4'�U�`�w�\iJ��qa���7e�#K�ٱ� ���;�Ve��.��k�j�w"m�Yۦ�oE]��D��z��.�q^я�L5��mʵ%v՗��ևtRe,۴6����<q�z�ǀ2b�J���}ap��;}���1C����WV(f�������Zֻ��{#7GA���7"�AJ��*̏2�o#��"���3i���4�[i�Jwt�M�8%��w��Q��X�m ���n#Q	k�h��T;L}��u����D����d�\��'����H�: ��כ���[Au��O;/H�5*fN�,��ø@��F�!�Bٜ�X��.�)��j�e!:D���^i�����4�^��J3d����s�Qk/����y٨!��	\�k����uu�M7 ��Ͳ$׏-���H��T<�x���+�to�}��_=l��.C�!�Ji��t^T]�&�=YL��ϰL2�a����<�8���v��Q�Ѡ�:);׭Z:�Y˻k|�޲.�M2s^E�yù�;�ԪYn��iQӽ����mLS�:��%���	ui-�3�����A���&ܝ����a�w�
�=��te��iGtEܴIdu�8Җ荾c6`�k%4�����D��Cfo~�872;*ao�5w!�v���u�]̮������3�G�[{��� ���ˡD��c��o>ot�׻繥�U��T]�s��Ǯ��f�����h�.�r	bYڷWT�z���N��Ɨ�geL�u[m���̴!��fiQT<�{���&o�g��w)�x�����X�V/2��#ڙ����P��e��_E%:����o�j���a-|�C�{��0��y6Y��rcv�!���L�ks�]ܭu����V��d�f�����4X�ܑ��rԮYy�㬔�����k�$�hZ�cF�@��]��ZkJ]չ��u��F XĆT�v�ec�jog_����╗u��*�tSA�m^�w��+AE� �w�a �U7]f��R��eW[A�Ȝ��5m]ra( +��הO����Ds:�tj��]�À�ݮ�|s���o{jkSs:�^��:�:.2]�:�wӱ����|N��ӧ�o�/��)\���N��wWhc�PTs�i7%M�+b䢪k%���\t�0i��u�%������Ey/��ŉ��`��)��ژ�!��&�>��Ru��1��r�j�+�M��m�/�٩�h�{����*v�ّn�H<hwRz��u��Ӭy� ��ۗ�++"7M5hN)�!�<��Q���[V�*I��Й��wh��P��-VFCU6���{��8�+�oY&th� #zm���>̩��:���9��LD�r+�3��vi
|��S�w���٬��N٠b��X��n�s/���NV�+�}�$^2�l�g3;��۸`y��ք;	��t�&�;rPē���ީs��⡞�ţ�f�$�i��1)�M��"˼���t��ż�TT:�@rJt&�fV�k4��sat #�z��U��:�3��ї�d�\v�V_j�8l;�r��i6���@n��骺����*�]z��lu|�u`m�b|�=#�f3���W�.�AJqU u)�s7;q1l��lwF�Tk�%X�V";i���ŷ2�C��-���"��VT6u��/l����y0��<99Z\�h:�G���VQ�-�yi���,�wK"���>��=�C��i��Q��1�*�v/��6�!l��;�+��"��J5�h`�vvb�p�q��o��]lwZoi�xML��lp�����z�z��ݙ{/T�`U����;�(]f�k�/1�c�����/ԩ�6��u�3�⳺*"�ye�a�@��S��E���7����r��4��Mvo|t���p 襗g�^h������V�·RN�
�����;P��⨞�P��'4WL��	|e�㮞��|1Ỳғt��d����h�&�����_qCw_'tm<{�27F&�.�Ũ@"U�]ZR�4Fm��'�F�eeI,����VQ�[�g)Uqeo"�A�����G#U�br��"]�l�ĸ�&ok�:�i����m��Μ��s*Ǜkk�U��_NUax�u��rXFPMS��a������#;Mj�qU�ۇ���M�q[Y������n�������N�V9�RJ��5�U�yu�\��^����zt�}�:SY�	
�� Rn��qڼ"��������ǈ�2���`6��'���C�ض8��gi!=��$+��Ƴ��3
�|�t���fP��Mռ�}d_<ؘf��{���z��h1����\�l��#U�]�G�{0�=e�x���~�*��Ek�n6��&�},�<��:��z�mu@)=��-X��k�)MȚ
�#�����g�Z�ou��ye;,=�5}��h|PV��"���x7\�5<�s@��f��5\�>X3{%m�L�6�յ��R:[�s������R���;�l��-7DcI��/mPWV�s)|�����MҪI��r�*b�v�Җ
��e�5�ΎM�n��I��}J����:��UK��n�(�ǃ��/��ϫlrۚ(m.T-����ghLS3��lK1�+���gd��T�^ 3�׎oUռm�R�1.J��)Ѕ�\�J�t� ����JO�֬�*�d��s[��T�����Ȃ�q]��G�ε��Ļ撛�EBM�ޱq15�/3W��h�/��N��);��Sz��2�^t3]���Qr����dy��#��-������>h�����r�'�M��`��<�ʾ�M��/j�rҪ��3���ho�C�:t����s�)��Ǽ%��v��W��.�5�9�FG}'kaх��!��R�vd���Z��Fǌ��l��h�˻�T�Cnf�jcIpKԍ���__�C9�;	4�T
�D��Kם�|O'S_v�+L�z�{����-�(�M�;j��)�Uq���ZqJ�>Xse���M����tH1�F�yy�_Gˮ�)�/ܴV�21V���b_ :��˥�BBwb�Nº+o3�[��;�ȅ��	��[�,̝�T9j�[���[��'_j/��F�LdV>�αZ:�W:�ԶdGd.dl)]n�A�mVL����i�WJ�%�暽����3�v�S���������s�m�_t
PwVdb�7����Sz���u����R�Ep�`���7[��4m�]�v�i<�d��3�̽�=�N��J����}����k�ǔ�왰7fu֛�� �]��l��Ytz�+h����zUa�[f���F�W>Z����S��z3M�I �Kr��.����-VS�͒b��ڜ�ᣈ����n
Hs�άe�|5v�\����7�q��]�9�����l���ki΄q-�h���o`�Ou�ӝv��v=�ip\���]��zOW�Մy�$z�gQ���u�5��wQr����-:�Ňk�9]�dJ��Ӻ����/�z�t-�X��2��%
��A"Q���:�B˽�Y�ZYn�
[5߉t;(�e٢Ś�>"R�r@
 �L�D( 	蘠"��H����WXS��&�	�6���Q���Sl�w�]2��n»ԙ�6�*aGJ���%2@f�h��|>'�*(������Vi4�-�
���l�L�	#���u�l	Rm��� ��(�z� ���|E�
�<+m��$0���P��!"«��h�^���\ǽ{���=���c1��߇G�͊���m���ֺsm�/���9���}<����N֥�r�����.c8�W�
u��dY����f´�ov]i�7j�o�!i�[��x�d
T�O�&���m���jL#}/"��!�A��it��<u�I&Y��uh
��N��uN��cDtT��Ńr��A���r�ԑ��eu��9�1Wn`�9P(�����h���%��
6Y��Q�8�X��f�f�\i����;�؁I2��1��[�]b�t&=�fZ��,]��A�m��y Ԯ��6��q.\�EZx�{��t���A'�k�*sP�]֛�R�8�Y9Z�hk�ۺN�A��!�]��{ʲ�7r�NBj��ʸ�q��y�T��vl_�}���b�����Ʋ�P�N��n��om5(bԬ�Ց��n�R�)Z1�ytU�qY�c�
Î���}I�m�Y}�V�h�5!T�_@x�O��w�#���Ѽ��[q�V#�:�1�5��qW���S�6�u���������qƐ�d<�*
��)�:��Z��ZҸ|�7W׃`�[�#�H�q�)���LlG�`ᷜ��(�R�+�4����졋�"��Z�-&gP{���l�<Uժީ�3�i�x ��I�ë7�|4sagF0�=\�5����U5Hm�����O"��JK�t5l��2aʕlJ5m�����G%�w�cדr�.���4WR�m�ν�|*me��N�kt8޵�g9f��6p��80"""""0"&DDDDK"""hDJ&�r�R����;����U�,+�[�l
��ҕ����\���Eֶ�Q `�ޖ�U� hRa��èt��;�\Y�;�`��IT�W�z]k��Ӵ��]���S�0>����84ucMp��W>�ME�[a�T�:�!�V1���1Zo�Ȗ��� �j����]z��G;W|��-U@VN��]{L[�;��<�,���7s_R�+a; �q����_s����ڛW�pT1,�W�S����~�.|����>�pR� |��B���I������5|�,l��ʴv���!�����"�e�9WB Yi`��ʓy�Kb�G��t�("r�u7c�t���r���f�]Z�rm��S��%[[(B���YVĥG�H�R���#�w��3vڭm0~����gS@\q�gu�����W(����i��u�R�(0�m��F��]�R�����/����UV��ዢ#"�L׬-|j�Q%�@�r��n��$�c7ki����U���>[�ذF�C�i��kn�A�e+��yD��C�)y��Lv�4�^L:�;ʮ��,5q+��Y׺Ì�����XH��˯#�9*5��ֱ/(Z�x��Ux��8,�����z1wqU��t�M,�j,ۭѲ��5F\��:����2��f���td]%$t�5��x�_a�=�v��}��uK6��Pa�n�}�\n��f�ۻ_����FN�K,�;Ј�8"H�F��B""&�DJ6""P���kW�������.#D�ȓ��T�ٙe��쇅+�d��do,��(�rU�)���
�u�*|�Fm��/qh����me{]m Y��$,V�_v��̈�T08z�&����+h���Q�V���XDx��U
���>��"��]u�����)\�i��N�H��;U���u2�G�m�_��+Lqǯy�#�.�)�v���4��ʇ6���O����b<%e�ɛж�"I�\S[��MC�rwHG&����wZ�����Q�JCj���o���p6�iⶕ|b��璵[�x�j�U(&fTd|;�#��_B`��_r���î�u>�m�sv�n����N���UG�삻-`:�z�u��[�[��થ6r�{�1+�Vq�
����C�rH���Bӣ�Du�0q(B���C�u�lD��a�	.��tv�����;���z��`*��^Ֆ�}�IEݦ��3��nns�
�Ee;�\F��Lά����{K�+r��\��n��vH��Q$����¶�G�W%&�9vU�.}LMTGD����M��Bn,��Ҕ��c;���MK��	ut�.{��o�?�)u�2^����x���}07�T�EY�j����v�����땳nG��\�WT1vmL�&o��Kmк���+@61ܸsi�3d��`-`���t�
��5�g;���FKe�8p�b%���4"&�2Q�B"&DDDM����_w��}Սn:�����'dL彥�"�`�%Y8�[G%�������P*md'���Rj�&��k�6l;p��n�ub���e�\T�)��������v/��q�3�.�U���H�Sd��t�^��]XF����$��t΅��fQ[е}ٽk^@`Nj���4�d�=D!�4r�� �^M�]>�Se_(�k��VK��û]���8�]���ռ�*�X�z�D��27�4MyF,^�fe�[q!�D"����6/>�==�:V+��*%���W�Gq�*�9�K�]�����`��xw�����d��y%�i��r�7N��\{f:g��X;�C&oh�vG����H5�ј�QV��e�Q����������0be;&����zŖ�X�[LV�흕;rZ��(��\ �1p���u&gM��΀�colҵ0t���{��B�MUV�]M�3(��V�ވ��	R����'kw(І�;%[��XR���cT) ��vD�R��mXzț/t6�P��m샮���ݱ����.�Wl7��֑���r�6	��J�Y1��:c�AGܩ�N��4���w�E]�4qj�Z�}q��]1r�iU�DZ�5*B^ˎ��E�Zz��M�����=��"ک����,��k��]��Z[���io���$��$f��L���;:����pe<�zĥkl�wX}V�n����iAv�/	N^늦����4Ve�i𖻪vͫ8��+�4��bٳ�͈�bH�����DJ(��DDDD�$DDDDKDDDDDL�'W�ᨯ���E����s���#���2��v�aiK�e�K���Ԕv��}t��7�7�*[�̪г��U��5
w�
=)���H���T�5ӄ���<+O.3(,oF_h�s.�X![)���^�O]k��WP/��R�ި�fY��o��9�ʐP�fۃ�����]4����IQT��]^>�]:(�YU6azEvoK���ήr�r��ʘ�ve�Vywm-Q��gd;��;��ǁ�Ga�I�\�5P��$���()X���h�����ym�Va՛}YP�U
Q��Zkq_�(�,�T�=�s�>ʒh�l�}�ђ��5h>"�j��eWQ��]Il����Τ��+C����:�J5����*�Ļc��.$+�	����&ʻ�ً���:�(�����<��	La��cE�f^���i#��a�R�Y4���z�76�T�u��MBS�M7�xj�m���7�+T�����p�ָu�����5pA˥wLҚV�v��2h��_w44G��9˷
�U�L˳� �Ǎav��1V���ڦL<.>����l�+ ��ܕ�Mnۖ1X����G��opө����׫����a��PY]���A�>���H�3-��u�u�Spr@���
��2�n�KK��e�G(��B�;16�7o8py6�H�����A7.��oq7!�}Q"��V�q���Hݍ��U�	�X7hj�ˏ��+�w���}�Z*��l��:�3�W�:2-�tJs�9Q��ݴ�7�cP��Y����4�����ɿ�&{������㏮�D�Y�.�
-�+ݾ2ӔB+�w-�eX9���jVTvX?h���:�:���&�oEtOt�3�bt�Y%�{��N}79a����WU���u��C��J��Ѿ�P���9f)��,����S'�����L���E_R�՛w|�����1��9 �@Hf,k2$_h�nc0�v��'*u��X�7\���oz�Q��v�N/-�4r�X��\I�c)��y4S!H�A}�-$����k�UswNU��V���i�} ��y#Z�&��2	i��u��{��*K�oO�Y{R�iݬ׍�+jq��k'i����`�i��2��o:Vr5�Zչk��u\��oہ���
�m���c��X�@�#����@`��`�)�����+r�J��,$����S���s�'�θj�b�x�2��s;2o8.[b�.\2��Y��T�� \��r� NŖh�Z��cC36����o���ݔy����3Py�*$���9w�fռ�˽�ZS�	E�(�T�x4dUd6�	��"]vU؎����3PϚ��:��$7���y$a$.��W�w�Y�:5���h�9к�+����a����@7E�7|�J���|�3V|�6+O74�Oz�yB���� ��N�+�Q�1��\�eԌ��t�Q«�AD������{R�Z�[b_[7M�����.������j�L�"薛�ޑZ$P��lW����\Պ�	���涺�,�Eј�Y����4�
EؠZ٭B�=�IW�X(�[{5�}��=��r�oDi���f|����a\�p48
�j��A�n�"�n4s�W!�f1�P��ҫ_v�en>�Lp4v��u����k�h<Y��u�$�WB�C����b�g�t�m�3��_ҋ�t�[<��kr1bl�]����>�m"�r�"�g>d�麒f�Qg_YaQd���΃-�}^]�˫0�����=c~t�Ь�u�2�	�ϲ���˥�o�L���׺C� 刮���u �2{�WCP_R�Õt6����'[r՞���bb��\ܝ2���rʉ���bE��mj/���Ὂ����=�9V�ݰ�U2_J	��-cxh�[X�`�Fہ7>�O4����>�b��v�����Uv�!A;���vFv���;����Il��(G�$�qeD�
9���'Q��ct᧧>�V5G�d��#��d�mދ�t�a=n��hh��v28C��;��n����
�Gk��FҐj�皶=��`q�sk.(j�Is(��E�v�l[H��7!�K�r���v�Wɺ0
��x�i�7���wXJT�l�\��+�ѴE ��K2d�t��Ә�;ʇ5#Yc�3(�����t����k)yVyr���:�ۼ�Kم;o����R�U��Co)�5���=q1-���eA��zS�N����y����B/��g�{-�B$/` ��V~Ÿ�_*άW�1�֤{�"��PE������O.�ZE��Ft������-bw��-�ۚ��y1��V�;Wr�e'���g=�(��E�L}����أ�� ̺3�b�7�5%�iK��4����_V��ۊ��P4�M�*m�M!�����a����ҪeOn�05͌����fh�-N�E��*_�PS�!�ڷ�'3(qF��s]u�_k�u�q��f����Bܽ�K�X�̃n�#jJ���!�1����[g�/,��\t�;��xfI[C�M�M�u�S�c�,>WA��M��W[���+3z#�lNFhM�3)����7֯dՀv��A7Q��K�Z�s��R���'�V�y�r,r�u�7��fSf��亯�zɻ�bb@s���u2/��T�z���Ӕ�a�Va��L�6���X�h��-��΃��{,8e������g+��6�m�8q7OD@�J'vh$��B��$��//^�:,	��m���:6I��ޙ��z7�̞���ņV�qXMu��c���wI��Cϝ�;��=ac�u���BU��zp1o:�Gp[j�nVn��:�1���b�U�s�<�v�n�IRt���J�v2(��2��gǈU�*��]�WV'���`��g��.)t�oZȄ9��������ۻް�uJ�)�j�d�L��rZ�h:���r���8��y�*�&�oJ-eE�'_^s�eq����\��j��j�`Q���7
���1����)��	�5TF
10�ۗu72Ո9e*K=[�-��j_����6�W�{\n#��.TM$0N,��%�g}ݝ�c�&��o��I\z>�o'�+/#J�rw���νA�X�R���>
)��efvi�Y%�Rq�˷�붫69�.Wj�xZ���u�kvԡ�]�
��0���ï�R�U^�����I+h�@�/���}y��ͣ�upS��1�V(�Q�ϊ�2�����ka�(#�#s@�^H��!�jS�L,�/r�~�:1W�����F�-"���y>
gS�ʇg]e>��(	�[�x��-[y�'��dә󠬖j. ��O�,�u�ƨ	6��˜�"�6��e�ml���ء��)X���V掾��^����:�#8oǛ�Գ6^��H��ٽu�����N���[Ğúgₒ�LŃ_ί�����=���C�B�m�������v{٤[�X�p�O6�Ij�s�����gtƨ.s �Q����w�ph���),:HNF񦂕��8)Y�/:�(�"X�m��w��J	��=y�E�s:�ܽ�9�A�6H��]]dgB8�Xȫ�Ev��K����U��3��cZ0A\S�ʟ$�gͬ���a����b
Zm+"\��Z�
]"�;�eG��[ٷ3 �<����7� ��wwpA��2�e�X�Rm�G$0��ۻV�r"���6��%9�����f6\�ǬJXl	5b��]�v�n��(c���s�i%�
;�WV3��$F�ʜZ���j��eX��@H�
D���Rt���K����c�����YH��F�R�e�N*A��|�I�J�V�uI3Ot:����h
��F��kP�$Ƭl-�,Q{pWp���[Ys��Uٱ,�b[�eުTa���%���b��f��0z�e�x���V�qI�t�)�a����Z����9�޸�����ĉ�9'ΉOY��{ys:�����}�_����*��1���������!�~;<ے�S����������U�l���4���C��_�O��|����S�ְ�D9W0�C��A��	Ku��>����|�]����u�Ь̘�%J�b�`�5c9�\+3��j�G�^�]|�
(���뷫�S�7|{�9۶�}@�ݭoE�s����qFY�*��٥�˵5�u��.�2�:@;�{{�����y���	ޏd�H9�_U������EԞ���}]��g��d���OI;� �j�K��'c��F�ɉ�F��p�B�*dRݹx(뎐���oz�cN����fQC�5!Ȼ�+t�̚֋�����h�(Z��<t���Xλb��^��5k8_X񎮼.]��V8�\p�]7��^S)�ѣ�"z3���V,�0�	�{(����K��wM�\6��0�O��ڛ�n@M�S��Gc�[eq���|(�j��6���%.�ky����̡��{�;{]�R�$w.�jUczP�Wjc%�	Uz��=�ν�.Kd���1g�ܮk����Ӗ'	���芾6딩�ZMuK��Q��:ۋ2���PW|��]��|�V�ͩ4��u.����r�=|p n��\���I�G)d�]�,��`�[�T��K M�i�=�ѧ�������+�9n�lv�=0D��8F2EE��Ŝb�۳�]*s�͒!�ն�r�k���#�P�|I)kb��J�ZL2hQ�Q���
Eh��m�T��(�.�ݰ%������W7wu<-q܎�o�@�"�^YG���9�G<�З'w'	����G	�\�n��Gz<��s�T�o���w��25��(�GYx��B���{���a��z_0�G0p^Z��c�U���	!��7�';�oy��S�v��{}�w��}ʴT�0�$�ؾ������R�r9鉑�yT��z��<�֘UT�[�V�M@��6i�{{}�w��}ߑ�)��Z��4ߔwW�*$ܑ��͏�x�T�����gB��p#�2+���~o����!��]ҽ���:W"�Y���YJ\p�sr�k��w�˖��$뻺#�^y�̙}hOw���g�۹�]�2<"����uD+�<
2U��9����.U:��J|��&�{����q
8��:,B>�u'W�S�G'K~�-�K4��y�s�UL���
T��^���ny)iX��u#�<��D�8�#�S�[�z���p�z��4!/����|��%H�Qq����w�7]���I�*(�1|�G|c�)���W����p��K���L�߾���e�
�U�;^	���vj�����չ�c�lejw����X.�.=h$w:e�&䤮���-��q�9�'@,��L�WpUf���bô�-�ή�Ga�wK�p����,�\Y���5v0?O����W<�y�x1������/�&:����_��m1��qz�2�37�񈑦=�.@�D�(�?WJ���������뗌s��i,���5�'� ���,���C��nu{"�����rO{���PÌ�H��W��ǅ�a����C�mZ!m7�Ԉ����.z6.�MZ]/U�r3gb>!�~����l�l���e�pA�;L���j��ַ�T��e�9�r��<}�~���_�B���+~�{^�D��A�eC�|8��QRgL�vU{��Q�1Ʒ_�W1���b9�`ޏw7�S!���5�a.e����������<緤U^���+�����P�I�<l\]�1Di���g��0��]�[��~�7�^}�/�|�ϐـ�ny���$������!�
�OQ���G$�6�����9{��j4M���͂��r]ʸ��ʹ A���'�2��Rm:�D�k�'t4'YzP��ܤ]�L�v3�hKU����Մna���n�1tթ|�-���K�>�鳠�鋩4hd��9������g�*eT^黮
lx�����^�x�嫸V�JGj�ɖ=\.φy��B��O]vp�1";�Y�b�wm{�p����ZX�6�X��ٞ�֓}^v�~8#��9Z�x��Fwmw��}�/>�϶a��7�ޯ=�+���;G����ML�����$�����o�9�i����s��U�U������Y�w�l=�����\u�^���q�O���zj�P����Ps�.��3�_�E�*į%@�ՏϫB�߮z�T_��������{㝞��O}{���ރ\��cL��� �r��eh�d�M{Y�'n:��^tؼ��t^;&Gj�����]F�ڿz�c�5�c�2M誖��q�"6I6�'��ɳۣ�s�X�*{#�0t�!�h%�zC�T1fT'Wf��O	�Ǻ��8�� ��II�'7K˖m
Ỉi��J�ac��:g���Q�8�m�����co��yʱ�4f;�J�]O���-u>������=S�H�:�dT:���YK�]�^u����S�qtJu�u�eC��g}]b0�Y�ޓ�X�H��OC�ǖ$Y��kn�=�[:]�מ�l��rvv��ڡ�[�,㘐	݁'z��}��Z�s�'�|�b�ۗR^ԧ2�K�NU7g�3�Wg"d���O�+5y����bw˻9�%�M�On���r��N�Oݿd������:#FW���}����YM�Y�����5S*ѩ�өc��e��Z4��H��7=|vD���|��v:�S�}(����AaԻCrĶfu�z_7ʯ<0�k�����2��ݽ[�uv};�+��G'�Z_�rn�n.<x��w�����=�M,�q}��P�;�{�յS�u���P�.�!l���1��E>t5X1���Tz"co2.�"x����67҉��/����z���T������ﮅ�����d��vU&�e��ѦS��{V���;�i�C)���s%�Y���|/u�����R��pc��Mն$�r��}5݋W�i�3A�*
[�<ͫJ=0wAvۧ��죱R��vX����AT|���9���k�k���k6���96��r���&��0�5;�oV��I�{�y�{��ҾZG�{Y�幒�n�I��a�n���avGkt�VzMx2veָ|���\hy˲sv�|E!O��[�����z�0a�V�6�#�춒g×�*������ض��ZF�{��G�s����9�u>߳�2��YT�߳wh�4�-�x�v\sM����T��Rj�{ڝ̧�J���W��,��E�"�����MC�wꑮ`E�>�������|>z�h�B��������^�Z��g����fx����4VgĹ�7�=�G:hq�{��k��� `v<�y�4�ztb�+6+ϽeH��ny�d�N�u���~���:�+>]Y�f��� "���X9=�������:`�Ў�v�7���]1�ڹ>ݝ�&����h�~,����(��]�m�#�oN{{L�����;'M�Rg<��^�vV�8�_ub5�WEy�P�5�4�(�j�.��C(���Ʊ�Z�T8�F�b�o	��)��!l���Orũj���c{	L���= A�j�s�����y�Yb�No5�������� -�g_=�	v����o��B��PJ�N���up�*��W�����0����jJ�\�w��us,��<񫖗�|gL��9Ed�1���x��ӣNP��RG�A����S��4�^��ʌZ����o<�n: ��vI�(���<�pCS����ۯ�R�<����jȓ�"�	26)̍�{�	�璺�3���O�J���|{F�ջ�������U��޶���;6!&�c�%�� �-�.��!�a�U�&��<�s���q3G�ў��p�g�0F>ݜӵW�n�ƍ��GrF�l��o�tO?�g_G�����oh��l� v[슶�\H��Ǵ[{�{o�n�'o�o�5+}1�n���~ާZ��L�/��$���5S���8d'���h�|��{F����<�p�ojs���A&l�l�ڦ^a�����m��z���i����C�r��%�Ks[�� ��(+�;�#(��{�P'�xLS|�ʿ �:/k�:�b�JӾ�{�|7��ڍ�}��Z��8a#�ѽ|U��En]%E�֧�T���1#�кu��s���c;�عu;/�N����kφ�r�ͣ��������Q�?]G�}�^���'�������C�و��=������K�;�(ԛ�����9q�����c>���]xG�هLᡳ�K��ݧhXwTW��3��r�'��dJ�~�}u�,WT�O�A[MM������5�L�ܓ�R��E��������q��@�Pn�4s8�{(c\^צ�t�)'�-$���{�.5�I��{����o�\��2���Cv�ׂ���s&��k�Qa-�PյR��@�W�.��7{���p���vȞ�Cq1��o�p�S�d�~�	}�S�����x����]��߽�/>j���s|���ihK�wo8=򨗆�ƻ��}̸��$��32<z�b��O<}/;ӷ}'�f�ר�~�)�o@Q�}ɡ���q+z7/���F�)�:�E��+u��`��q!���c+����.ʈ�l��{����Fz�y�~s�N�}%g)���Gt;V��-����=�k(�e��C�}��E. f�q</�c�ͨL�w���vS��2o�ܾ�'V;�k��`j?z���t+~:G��z���a��4���/J{���O8�q�7ǜ񇄚��^��h&���}���@�c����LՋ�s�.�ޏ�E�h�_g�l7A5'\Q�q7T�l�ә��
�ہ�z�F�sl{�m/gRϼ���EᛳǇA�|�&l��ut�������2���5����[�T*�?nu6�y�?��8�y}~�~�E����wm������o��WG�����0=��a�О~�߼��|c}fyX�)�6��u���<ٮn ���xp͏0�`w���ix�}��K7���K��ZZ}�9���o����v�'�M��ꃪv
~�.9f��pe	.q��,�E��Ξ/�d8n���Ttk��R�]_o
W�,���������t6��w���>i����=��y�L�ur��:V��V*��[$��{��V�V�r�fq��C}�ېW|��l*ʖ4 :�8:�^�+I궒�F�XKc�L�,�x���g��m��C�˻�}OoU��c~���
��oc8��!Y	�R�ۮv����^(zw�u��C��r����ו�CJp���;`}wS��9�z7�j�R>�/_��ʖ.���O�oV�uv};�9����og��F����qz�O�f����
�M	��_H=BN��oQl�m�>��%cs:�{�D;��:�u�VD��t�����i{��y�>;�=0��N�r��(�N�m3��U6��WW�����7�v[�G�Qrq�l�p3]�v2�q7kÏkwMg�i�E ���
:�fޯ�W1?>~-W��B�ί3�I�g��1��\���^6D��\�m������tГO�Ȍ��b m��I4��'�ɗև�ݫ����"`]�:ɜ���='Օ�Y����f�c�x��o�ǈ�!��۴�{j�;1���\���w�����˔�P�(�{Z��[c��[|v�y�)WV��v��N�o7I����<��ώ׫�(p�2�=&vv����݉cW[>܂��樆��q���������SǕ@�*�X�=����ê|�8��&묞B��v�������s"�4�e�܋k��R�e\C��\e���8�>�� �L���opW^�]X�|��]q,nU����Ԍ�6*:؈s.�E���3U��l��n��3
�7��#���'�@=� ��5k>�O�K��xx�oq�9@:���>�a/}�GŚ�q'�ݧ�{�����1]?��|���d��A��?yP~]��5;�F�`��i��=�@���"�x��������1nI���>�c��7�Eɕ�g8���Y�uc��8mG�uӣ�2�fw�(v{�(yy]^���5����%H�
|8uF�+��7*��8�*;K���n=�(���C8#�>t�>��r��x�Y��*y-�SLM����j�H�4�G�_�Y��~e��/�S�����w�ɗ��5e��g�{��];�յ;����hk鶫�/(~��e�s�����>���v�m��i9|A51��kHͨ�����w��A�:��9�VQ�z�g�z�/z}� �u�����zM=u����[�:�u��Ӎ���b����w�}���=vg	���+�M�9y���m�ֺ�s�W���E�p,��C�b���{M��$v�M����{�4]1�Z���!����X�qeA޽�Ђ��L�^j�l;�h�$��p�G��b��&q����4ڧ��ؽu����Ѥ����0l3Q:e��6d`ۧ���@/�6���&Ub����J�����������.��Co�r��<��uQl�&�l��d6�ϩڜ�c���z�� �_���>�*ks�Z��c�\�zdȳͲ;���8a/^�Rg#gY�{M���&;��U^ͳ{��OYؚ�:Owx�>Ɇ��ƙ���n��VN=�s���fM�d��7�k�2~��vmI�?xɵ^P��NK;9�Zn&�:o�@f���`��6����U��>��ݾ���ލ5�@�1��c7nP8d��I��[�|�5�p�a��V��P���֦L�c_?~�Q-�ў���϶���W�R��S�vk��vrsM����G�;G�xIz��y9q'|Ĉ�\��iA��?�^�`~�>���>-�;�<==�ٌ������.���e���Ou����-1t��m�Zjd�&�f�У(t�qHQ�����8��2��vS�*:#.(*��v`ɢ'��c4�+��Fˀ�KQ
f�	ގ����pg{'i��o�R��	QS]�����A���:��k���N�t�{�fs�(B�̨��\�Hs��[�=�x^�� 2rU�{�q�!�BJ���۶g+Y؜I��.�|jS��>��@�Y�v#�H��[S�t��`W�xqSR�t�h�g��-�W��\�vK3���:q�$6��̾,�n���j6��n�߯ɠY����j[�wEm���!+y�1�:�ʌŗ��=#�g
��������1�ƅc۶��K�����J"��:�����	���3�yy�R���fn:V�(.bԧ��F��]w�$�MB��;3�6_=롻1
�0R�����#To���3��\:���ū������[M�[�N��v�=ð(�}���8�Vg}*֌Փ5r���Yӽ�+<�ʴ�6��>�+fU�K{L��'��38�Y�_�f��C�#�!�`����v���g6��$���[��$�[f^w0�ͣ����m`�5+�b�{%
[�5��$t�=���eb:�չ�y[ٌZ��Oi`��$�gǸߕ�����7�!�r���ZV�q�YǬm��kv�	ȭGcIN�Pm��On��L;���֣ê�guP��z��^���w{򥔨|y[)�wt[|�+�铪W#�}�r���d8L���	J��[���^��[�Ë��q�uG�{KF��6�s�=-h��v�jgww_c��uu�<��3Y��Z�X�����y|i�ԕ�@!�hϞ"�w��R#i���*���պ�I���>��-DUҗ@����D�r�v�����U�bR���w���Jqɖi7��o�Q̲e�*�FX΄�Z��0�I�P��]m�c���̠>=-�GR�EC����S�[�������0l��Ibpyu�2�\����Yo
�g���n�Q}�Rh���Wp<�ZhЁ���GXط��a��0�wqx,Zr�if��
��OzS�B�-�0�-2����7�[@ޑ9�6ȐCu�cmК务¯�������zp`n��k�L)��'�)�Hh�����q�j����f��)V^�	���c�<�h[{eK�G�Ɏ�+��9��w���/��˿<��G�5�~ �wSb^Q�mNSz�tՁH:�gV�� c
�ywq��B�v�\���z���ʺs��"�um��YM���&\Y�t�˹\�Q���NJ;��ͫeD��R�0vtyf�W\Z�k�Ջ�&�wژ�pYPmp�\i7���'sz�V�S�Z�Z��m��h��ÉA���8�]�Sꆺ�m�=�������3<�\����|d�B�y��x�76������HR�ݑ]�(ϻ^g{���+�έo�������q~|޽�T�=br�ڧ�s�;$*��#�㢒��"�ǟ%Wر�qЎO�<\|�p��T�����o��|�u���O��/6���x�QTB��N�5�NK��`x�	�C,!a��x��u�]ۺz:�=��|��w��}�1_i>��a1	|t���v�'�O/x�ry$\s�.\' y�}�K�,��g�>�I��<qq��)�=��v=�.�7oo�����r��Q�f��q;����<��Ǻ}S/:W�K�3��p�U貔�v"DE9�]�'H}����<T��]���񷓞N}��wy^Tn�Ϲ�כ��w�ς����j.Q$�;�V�⤃���*5� �K��B봼��|��~/��|��$��*���{����g�H���(5!38��	��{�n�DNt?I��>|�c���+M9�9�h�E'w<�~%�N�
y�{�U:SID4���"';�^���>V�{�¨�u<�O	u��8ܩP�ZF�D���'w�ϑ�4��o[��}��;����u��CM��SC;��ƣ��[˂�ʛ�*��죻��h��vՉ"]�2�p�v�j�4,�|�.W%�U}+��y;�\�9��eF�A��n�0v�p	��HM;�O��f`�6ޖ��ĳ��iw:��M>CY�MlZ���Ί�߻�`���z ����~l��>�ͧ�ʃ�v��[�[}Y��#�a�^�_�4pd>�����ۓ6�5%@3m�2�*�7ޯ@L�ݸ�Κf��	��9���c�@����M�h���a�yq��R�%s�^��g�ɳv�r�R��Ξع67�3H�5jә�?x�]��b`�H3©6;��_,.@��հ��\�B�M���������,�� `��%�&�)�d�Jj�����l��w�J��yç{;�kY���KK����O�Sw������%8	>9�N�@�@qJ�[\u�5x>Eë��aLգ
[&�jm^�ء)��z/��)S	��;.�O�J��JN1I��7H��K?����/��+C��oM�
3(��3��}o�Ȃ�^����ܞi/��c�����Z~XH-��Y�/y��d�̉���O��1,P���[>`�Za����յ�M���\�`�/�0d����|��`�l��y��؍(�v�ec߮�C):��e���˾l�|��R�d���Rv�U},�-��i�T�'+w�2��3mԉ)k��x����R��7�>�8�L#gh4yu�0�&�\�>��D������<L�?=�i/nD��	���M�����<;�{c�@C`t���L;'��"yј��I:���
6ws6n�s�x{�2�����]#%+!@�Q�y�C���w#�ۦ朶�����y=��t���S�����H�m�Q@sQ}����!ۤ{����73����c�H�/�����q�����>1�R�ν�y[y�����ߙ�H���+���-E�;���X�|�i�]�wu9��u�	L�	���s~�ԍd�ú�?D�B( Qv�	�b��0]��M�4�3�s[	�ݸL5��B���T�>A�4������N��q�����4y�o�l�V�Q��<����f���<?�m��dX�8�P�b��=��M���
FՏ�7R[�u��KcwScC󺎵�� �#;(�p� �M^*�(ų�E2op�Ο�]�`t�}���{`o�].
/i�z����Qhu!9^���a��]���ȣ:��o�YQp����P+�\���7�F�d�U=wcoh/�*#��켶tM@�	�E��`e�`����
V��
j
��x�mt���~�~��G`���ۘOK���NWYi��/�M��fJ˾���V\����VD�i�a���Y��qW9�6����3o�w�Z�<8{6��
}:���+�%9�wsNj$�N�hv��y ���"s���10@�t��5��lШG7���5��.ӹ.�'�KsOЙ'�1)դhZS)8�[��#s˫�gN_2���m���ޑ����؆W��q0���L0��2��b�6���>�S�Z�5k��n��C1*
��6^����}�B1���'�pG>v@�U�>-#��k�Ɗ�:i�ﳕmj6��fۓ��sN"�6�vk�����kd-}�!���.�.^��Yc��������c?�w���(�.y`�"���z�U��!<;��Tx��q]�U��Hl��t����^��k�Br+_l*���$��3Ī�-t� �T�/vZ���Ƹ`Ћ���^�jJ�s	�
�S�O�?7P�ʹ	��VJ�~�W=���G0�z���k�~��1�%Yٲ-�J�0r#�Ϡ�0 >'46��m�,9��T��t]�1�;#K/�ó[4ɫZ�fm[S/Z�z��
 3� ?�!끀�0���~Ɇd��f�g�ń�l5�p����ym�Z�e���30��D�qL��\	w��02*�F��y���j־��M�qCi�Ά���}�16��}�����Z*ή
l��>6��� �����J�Ш�R�G�6e�ڵ���+��J�F����G��uJ��hp�Q��bŖ:C�K�Z}'Y�F�s��+v��<C{��\�^@zH����&,� �^�!���$=�r2�>:"�s�8��f`0&@B,�bKB5�[�4d<�R�t�/Z����C�P��׊�"g͢�i�WL\8�Y��_`�\���%Vi�
�*��D]��UF5Ɇ�<^���,�`�u���0��Ej�ͫ!L�ܮμ]�� ��r��L&�q����3���jc��q�4!1�F�'��k��x�mz�|ĝ���1x�cռ0Ol� ?0e6ԜI�&C�|Cu���������>�G7Qm\����w����MAJT.�l�=k�<'�p1�[@N�|�L��hU]�w��|{��f2�SE�C���;Ϙ�%�u��L��0�?B���̘����	�@�L=�j��E=��EKcܓ�K�plC-�NR��y�I�L,jQu�n�eX���
:�;;��`���׀ޣ'Y�u���� ��kg���1��B�����P8���f ���P�����ĸv��Kzu�DE,�s��xA�p�kkP��hLJu��m:v�.�%Q���Τ����E�cv�6�����5Sԡ�ll��(˗�p�]x8���Ij=���s��94E����	ϧ-��+3T��7��q�A���Y�E��"su)���p�
�*Uc�]-�7�5�&���1��78w<�"�IBfc�74���v�F����������Ҋ_��w������"�����p~����'�h��PښmV:����OZ��-z���bb+�kpUͷ�1���:ˍi�f����0`(p���p�]6���q�nt�'�TίX��m��G#�\��c�Ӂ�ǣ}�3<�Xu�1��g�3���	�Y�5����Jm�*���^������C6�Y$���I�(��� ��b�:�;�x9a��v�V
:����C��D�c�ҝ~���k�{�ҼMx1�n�0v����"��W��v-��{v(�{��y��$��gu9�xH�ii�Й�ۓ�Qx�pwP֚�sL�B�KE]Ԍp�f,͈�Ӊ�n:�xi�,Bii&��(6*���Crf�RR͖a=́�yrL'��o;Ws��Xk-����Yٺ��z|zo^*��w��ŴxXt�	�\zxB�`�	دɲ��f�O�9�}�vyy��͞�р%?x*3�(�Ƕ�x/���xA@��f0ʈ��:�܉�	���/�ow��љE��	���Y'���+T�5����c�� U=�e?�vc��Yj�&��لQ�
|F<�r؆2��/*=h9tĮc[� �rw㵴��ݽ�$�����V��"���[l��4��G�f/��C��R��.��ݺ�e�P�d2���8��d�&P�t�%k���%!��D��P���S�ʜ�_`��&zs+GkV���}�� 7�7���T�8�bzvj�c�d��!	��|ޱ}4�㘔��H�U�&��G\�W� �Oٺ�"MH���Q���//H�f���̨L�{%��H�$�4��:z�) �"�),9�T�`f��m���꾭���/�b�>G����#�C�����ܞ`(���a��&�z����`ͻ�����dlr"�
�^�M#���z<��"����s���-z����U�y4�#z���L>�Z�Mwttޢޖ�*�kzGs��q������¼���`�w;�'リ�s��悒���y���Y|B��NV5��Rr،y>W>U0 u��_څ���P��>�3��djmg7�&w�u����i�K��L:��5�=�x�����[m���B�z5ͭ2�:黈��y��PPΨE�i�؞�ڀ�׻U�i'���0�_�՘�j/�ܶ�Q�[,����L0�5֎�p�GCS�,�=3� �W��XT�s�R5��wPns�g�4f�� L�3�����-��֙k�.�Hz��x9�@��4\sLI��uc�q��s��Fe�f��peM,�邤*�[���T��t֊K;����b��V�])en����]b��������K<�G��η���e)��`zO+�w6M�y���!�e�i���wR,�]�ҕk}}��3z�S�m�D�S;��\l��'K��A��<�裻��x<޾^���{����z�WE�?�ɑ� �{ �^B[#<�mv��m�j$˴��Z3���5�%eyS�`�FՏ�5W%��`�/��|Fe�����g�5��\�,MA�3��3f�Vo�cBz���X02@��g�����+1_I�{a�,�ȫj����0�	�8�M�(γю�ƯeEÛp�Ӈ�;����U��T)B�M�U��iӬg�\��2ǲb���J�RaMAu�6�r�\+��q/$�wmU���{g@@�=�P2dm�L,v��.�'�SsP~��=���i<_�4,}��9o���������[�g���.x��m]8ސC�X�H8���ۃm�Cp�I�୯,(ZY��3�3���%���(�Ě�`A�/N�o$n@A�v!?p�s��%�ナ9��^���f�^�B������6Ⱥ�^4�E��vk���3��p���-y�7s���f�����,;e�(5Ƹ�,��y�&�b�,'�J疠r�'�_����lB��V�8Y��s�8�ih���:�-�
ZЅ�Ƚ���uf��� ĝqd�,Zq��vU�W\�B{����4Y����"<g��#���kr�\�4 ��Cќ�c�kêQH�L��ox���{-�dS����#m�(��[\��2\��Î���z��_2�k��]��%[��s�M�t�U�q��
�ssF�+��/4�]Y��0�y��� y�=�9]<(#�`�z��`�Ť@��]09��Ȥ^8�<��{J	{kU s�{��y���Va��*d-�;�	�2�# G��!�Z`?s��f���E�5�Psi��]��<;j�NZk��.J�;n����mj=Ӗ��pȗx�����8x���fI��n�wf�sm�{����eE�,aX����7c�30�����-���;�@���^})�T샞��[j�d��^F�����wH$9Nm r2�t;z�s�MĴ���f|��c�Y�$gvVl�	��J{�/��c1�����*�!H��O�6�5�����Bv!~WQm{�����*���?}t�R���iһs�}u
�:�y�+ܤ-|.��]
6Up����Rxi�ţVL�'~s��>�|���� �4��i��՟L2Q���~"Se�d&O%��`6��o-��`ѝ���
�YG(]���4��]=��x�ҜI�&C�}�!��օIyܻ��n�NK7�k���"uՕ%�jR�}���5�з�x���2A� �'�;N��֦����,?+����ƌͷ�5p���Qvi���Ue<������ZX�o�}^��p��.�]N�J���TT�I�{;� R���d}:�ڬ�<=/��^�W)�e�����M�N��|bwE
�5b�pn��]W�n��e���>�xy������y��xx,�ǈΫIS�>���):�1,���tS"�����v��+N���!�9n�~�ؿ"qx�&�l�jN<9�N4�U�J{"���"�7E2�e۸4����u���d��eCU���9�AkH�f�Q�9�L��
:R�����Y�O�b����)�~`3	�������v�6 �t)@{��<`0rڼ�%�5鉷T:��-^:v�߉Td�Q��e�'�]0�\��h�ѻѝ.���@r�m ����� ä0�������WL��J����S�³�rv��"og�C6��K�ָ?]�6W+y�@�r��K�Z#O��"7��_�m�$�X���R��s�1Fv������&}:��3<Ǫ�z�H0�{���t6�dd�n�C��� b��wR0�]mC����	~����Y&+��-�P��g��.s���mC]���ɹG/��v���LN����f�8M O�k;O����o���p�۰��1�����W*�Mu�����a�\K<p�ii# ���$���gui��L�}�*�r�6H쩺wq���N�-%��I=�R~X��<1�f'�y_&l�W��{�Ƽ��W���RU�̛=^��#���ր���'\}6pMZ�4WwEh@��*	E>$Z�y�{;$|U�-^J��WG3�1��'z��n�����7���� �`<=ॕ��(�h�0��o�)�z�eZX*�x0�_��)j�q��㛓6ڒ�l�}c�����]�rܓ!��b�'{�+�{�!�e��W:���5aU�E�.==R�%&�hȕt��N�.������W�g	��0�& Z3I�w�]/{�(c���e7C.����C"��ߞ��s��_f�Q��③�b�f�!8��=�$f�_�*Mv":��=���On�S�ї� �!�-����3BPՑ<����!�<��	�v��.�L��5��\�Z�0u���m��e�,��=��)
��vm�	��vK�R;$É�I>y�T�(*[�R&�M�\-�������N`Yz�Zv����f�G���M�1��۹<�_�)�v!7K�ǱѝΦ��M�vcO3Z�{��	u������	=�XE�2�F�Ñ�$C�-z���6W6k�[#q(ս��ܮE:|���61��Λ�h1.�c!��0~�vd�p��i���lT�+�G!��O�6�R@�k��2m��Ϡ�f�طvm���o�h����`Ư]�߿���#￿����e�g��eԜw���!����L0��oi:�/E�x]� m�CG�Cx/cx	��U:RQx
E�X���p+�c�������P���w�]��"wV�|�5�d�Oe7�kF�Ѩڧ�]6��.�[(+��*��^A��u��B#��3�ͦ�h��c��D�t�H2�z�B�u���Ҷ��I�&��0e4�1�3v��{xct�=�]�an�u�9�U��Ts[;K�߮p�CP���OlT� &�K�V��XZ���vN�8]ep"[5�^�4M��Ѿ����|�1g����]˛�C&�z�q�fU��-lu��w7R�mBV��P����wgB��h�Q��9[K�5�%Jk��d��h��fKz�loj�#�L=��]ec���k}��}��N��+���4�̺����FQ\�9����G:m��^�������o
�cyR.S��d�7o]u����cխ����˹�eL�o�p�v�[�����W������[�tN��c��̇�j ���:����&E(�\i[T(��lv�
\x ����J�t���4�˦�)*躣3���*P�G>����7�g9���jP9Z棥���kj�bƴ�/�XWӻǯ缯L�ۥ�x�u$������V%��7G�]a	�s���Yd�f�(�:�eD�g.e�v����j�r�����X�fH��5���h]��F�17�R��ܔ%_&6����Q-����[N���5k��W8�8yuT`M6	z,&�	ҊU���
�J/�$�%�x� v�1����-��|jJ5o��n�K����`qU����Q��{˓�B�p�������	Ʉ��+�����}ɽZ�uy�+�G2%;l�0M#,4�R�=7�S�ܬu"��S5�ܸ��vpQ��;�E�P�u]]#C���q�U���\����]j׽u���x�=�gq��T�ZB�6T>�y��2��\Wv��_�8wu-����0LL#Ԧ�5�����y<�qV�/�Y���>�'F��o�[U�m-9��
H��\��c��e�!5��w�|�ǁ��&b��r<ˈ��'¦8*�%f�\q�S.�S&x���Xv��1q�s�X#��d�l�2�,�M��->�dN0����p\Y��<N�$��t9�+fр�r�&P�u�݇m-r�W��Vqڌ	\��x��X�e&$��B@j�n�\V��p���a�p�˧�P����̮�E�j'����ь4,Y#��e�Gq��p��ǡ�(1׏���R[Q�Ŕ$�o_"�E���Y���Ů��D��qt��l�65]����9�Qzh8�KwQ�*�$'��IT=|��w[0Q�s������E{�O����TڮƜd�g&�{"��C�%m� uđ|0�W$y�a�u���E�v0��k]�㱮����w���s�WW]>���zF��hG�Ra"��=�a8RU�]����|$��{����{���o�B�i><�9WY�Ae��s�n�Ąx���"�(��t4r��)Ց�������o��I&\I$��9�Ww#̫+�e(�O��><K�3��E^I9�Bi�����}�w��J�ԗ��X�~?{��l���fj_6�N�d��M8] ����ꉑR��oo�����&WEo�#��"8�F�QJ�<���}F�=�+���S�u�R�9d'�^���o����o�RT

�^r�K�$�r}t�AAt�<��y��P��g����T�W���8A+��/!�K��RO]�G=H��nxaRj/<<�9E"�(�R����E
�J�9⤊5i�T�����5 �2�<�aܟ8�P�(9�a9�S"'<�P�M.�,�T]�r�(�EQL��q*�#���$��!�))�,ȭe�0�����y�}@��L+R��OVEvE{��)�t:v�s[wS��7t-�E�E ��\�q]~���J��k���ݜagMf]Z5:��ځge�ӡ�H.LT`�ۤ����om�0v:���� �G�~}���{�����v��9����{�{��R�|*�cU��v�8���{M�'S,;�c��ǥ�´����G�tH۞��nq��i�Kf�����p�δF74��g=�d�@v��e'���0�p, �q��zS�6����صڻ")@os[+{��<{�v���g�X�6�k%c��s�;��]��m���aZ��c�s��YV�w�&���x[ἁ�	i�Ag�X�=�8�}�9�>��
��L�c�E�TJ[ѳҙ�z�u;RSl�PE��M����x86E;�."��aql��Q~�,m`{����}���ƑY�I�����Pb�[>�ٶT2���s��D��E9p;��F[k�����k�
��	\�U�{L �Z�A=�%��k9~��̨�sG��U�!�_����������q�&$�H�;>��!s�:��b���#B����M�H4�= ����yD�7�cW2ʋ��|g�s��2��!�v�;%؉����	�{bS��shX+X����[p�]�:q�c�A��� �4�t��bmC��Θl�+\��,�I�K�L���o2�f���s�]����|�yB��̕ DG�P����'7E � J��g_<�J���&c�N)�c5�y�x��Y?O���r��H�P��i,o�l�������!�#u���m+���x �o{���y�����-��%wY����`쭺E'�
&��A�/A�-��@AƿC���`χ�[�ѢdY��2����ٓ�0K�Ͳ.���#i@��;�?<�m8�-�h�l2��=t����5�]B��v�
�rW<��I����4��0��ٷ��i��EY�UH�;!cO�۝ƶ�Ƽ�]6bN��%QaV�y�ں�^���r��X=��ae�͑h�u.3���0r�� M����dROj�/ҹ��A/m���r��tMki���z�Q��t��I�Ã���~k��Pc�R̶��E�1Ԥam��A�Q�B-a��7�tm�t3a�w��si�^�^�9�����x���fIъf�N�ō�c!�x��f�;2�����1�+����m�c�k~¼x"U�YF��`��'�aF�eC����ޟ#��ny�����7u�ay�] ��
��r0�:�ҹ;({M$~$��@�9}��GP���<�L�ݢ�Tf����4�BA��/@rDϚ�%�g�� �%��}�AC��_�G-L�/�Y���uwv�:!C��ϸ��թQ�q�B��
�뢥
�}D'ҧ5�퇲��G�
K��r�����iUc��NI�j�Ku���3�+�e�h������Ƈ3O5�I*Z�{��;�2��Ws��݈gz��ѯ-��v]�|=�}��o0��y��� �� ���F���~��}�*��p�W4^��NT���c�t��B�z�\�6lU���g\:�6����lS<p��c`�-p�9�c%�v������</.���y�~��x����A����+�d��W��f����m%���866����w�	Ջٵ5�w�Z��G7��&Sԥ*u�S�~VЬ������胝p�K�mR��|��Սeb�Ot�N�1�d�`n�dR�ß���]D'�}f�6CZ��Q�r[
�|N�	Lܢ-�ǡ/��}��$�I��y.�/b7J�ctS*�;u�����s�Ht�6(��|q̠��8}h��͍"8G7C��}�b�iC����^�ŧ洣|\�v�|M55/�Ĭ��<p�N)w,���x�}�����֘� ku	�.�:�-~�;B����
��,��h���M�[�䬺	=,�� �8x���#Xt�G�í~�6��U̖�W�r�vXsw*��\�|��K炸%�^¸�n�k��?O�H`�9���ݛ]3ஶ�`��?M��i�X�
�c�yW�5�W�LDռx�FZ,��ד�,8�Ƌ���,�̻<���r��;0A3is9D��s��;-�����o�W�L2�ĵSXv�kD�Q�o���MmL�}�7��a�в����B��1�7�3me�QZ�cU�N+m�K|i���u&�&$ox����W�]&ʍNՏ�Xf۬)T��x�}�g�N�3<�\��s���~�`>���m.�k����S�u.��۲�{%�c�^�"�&+���-���
Y�a�H�F�:��˩=��W;��l ��q1=6_e�]"M3�������D8�vX�����_^n'�09��DT>P1,��K�[=l��T^=��ٖe���$� и'Ek%�����3vz�0c�л$��<�����A֖�����f��H�|w")�t�H=�i��Z^��wN�Jf��!��6�5r��o{��i�h��[G�:/".==���}��BB��\�S*����Jr(w��!)��A�Fi=�Q��>�L�`C<�sF��E>�>����C��X���'a(Da��n�B�b�j�� �P&%�t�K%&KR�G[�P�t��5V����i�琮���k���.A��f�o9`pv4�'�Iz�)�|s�Z�ʇ�T���o^;���ػ6a�mRͯP��y�t3[HT�mLpe#�]��;��.��'*��]��t�����ڴVKa�̢8}���'+��hZB��o?z��:����(��0�a���%��Ǣ�~�@Ռ�t�N�Pi�D�k�U3*Kv�� �v1ftü�uKVn��U��ˠ�j�"nhҧ:·lމ��T�����;����m����v&���߈]��	�!�߷i0-^F,�>G�d4[A�;	�D�L��KV9��R7�fnҡYy��i�t3 �$(�.h�3L$���[,kH�s�ge�g�gw<�6y���FR����vvWx�X���/IGs�	��t��v��vW�y�\�l93*)�I�+�B���=�L�v�U
��7�Θ5�}й���d�ͅs� �K6W�-ݛga�oj�����v媫)a퐮<�X|O>�n~Ǡ'����ȥΥ0�c���V�5\����wY3����4��Gf�_�J��7�	�<D&,�����{L��;I86#4$@9Y��gf��5�F^�F^n51���{� �x��сAi0���H�J��79���ҙ�m�Q���9�kc�og{r�����`���:"��<����%�q���	:�m�7s̛�i��ld�+CK�p��^f�JNԔ� �9v�}kO\�o�E;�.!�2�m��1.g�gWd0���U\���mcbr�ϛE�A�QW3��g�fͲ�Ο=;�ӎ��=a����nW�[�m
����SI�e	���=;�c��c����,�nd�������O%�e�n��rw0p]hF?�;�j���{��2�T㜲�*�W50��v�.Kv��u�j֞��q�Z.M���8���������������9 �Ó B��oR*�R�(F�ϡ��P��ߧ"��i��at����Q�g��|k��Ѻ�5�@��{�^.��p�..����*by�F��M^���oЃ,~�ؤ��hR+F�WX�B��nԻ����v�R����Qp�B��D&�Y��0���K�	��I���2Ovp�]d=�>\��)&7���m��hZ�`�j�]�N0��Шt�zA|gd���F����l���Q�.߶�Z�;�y�z�ekv �b�7L5'�Ba�&�������n���P�4}_�5qM1k~�9t�HᎲ�Ke�P�;*Jz�6Ⱥ�^4�-#=�U��w�~vlb3�!��8�����:hhB��><�%��R>�o`�&r<��I���Ƃ;P�Bxwfm2�n5�n�&QxF�S��N1�0~nwܟ�W:�WB̓u�߁*�
����Oa]kZC���׾q#�«�9j9��^��X0i������p�1��#�k�еaD�qź��p��w5�TD�]�B�uv��*5�����A߳�0~��69�@}O�61��{'�pd!����D��֠_�I[o�g 5bhnP<,�ȥ;��x�b,';��V�.+�gT��ISź5M���?����ve7�k�}��������h� ���f	���D��æ�]�]��S' �5.M�4ǚ�.聫��c7�{x�5�5� FZ�����a�rʘg��Ss�R0��� =�&���]hg�f��f��q�nc��E���Lw�8�	�����;�X@o�*�i��)]驚��.�n��E�/�A2͞,��fA�Ƴ�#���xC N7U���m,�gOXO.��V?0���Ywt�̋/;��Or2� �eC�mኛ�6�t��/�۱]ѓSs���fq!���1�t����{m׶�tC�� �Uz[�3�4��D3�Bw��Q'�ቋ�T���1p�@�3�t�)����{��j��-o��B׽0�y��~[�r�;��S�[~�#ނ�Ꝫ�T�C�ئxM�>�0Za�s�(�K�jo���_7y(�9V�^h�*{�����Ods*�hR{
�P��5�cռ4�{gh@Ųa�&C��f�U5/�4��y�=y���]�%�9BSbS�JKԥ*b6o����z��y-��TLxb"5�%��M���5!0Ǖ�	�5��):�ĲN���L��I�y�+�5�Bu�*.\�{�ܻ��gP�f��SЗ!�{{�J����dQt��]&�U�ӷ]bN^����o�![F=��&z���e���z�5��'�M�m�\x6�k�ݹ�������ʉ\���G�L�8vP�(���nG��F�d<����S�2,�rWQ�Zr�Q=0$��75����$,�p5#v�t�35�m��a��_��>��`<� b(�"e])�6�Z뮣/���8�+kPъ��]5_��a�F�҇@⮗�f-?4�6�����R�;�[�lY����w�p���sP������$������h^�f����4�W\]-�ͧ���E�m]�@����r���a�G��k���ԙC79ͮz{�W+y�+gkXP+�sߊ�^��+�cu���f��y�k��#�߭;��T���,�n6�L��q�,3l�T�ߓ�S�>�z�3�G�Y����A��;f˘׺	&��o*2��;zC�P�O"y�=�hb���z���b�=%�H@[^	EzB�šv�n��t�B�'l��tt� A�8��6^��f�D�b@ݬ`�#�	@����f�=e��3�k���G��a;/
t,���G���M����F���}�^�s��v�z ��PV��K�������ݔ��/^]+�dÇ�ٴ���6��5���CW�P���\ટO<��ٻ�v�)�5v����g�27z���)A�SlnC��y��V�S�-�â��X<@朥�ld\iܘ���/YSk��8��M���֥A�j�6�G
����լN׫0S�]�cyB���wU˗����:9�2&H��3mD6��!8�t��ωګ� �+�R6>�x�TݻqmN�o��]���֦l��nѝ8�7n���y����{��=�La��;������~���~~�����+ӟ	�,9X����D���Z��4�I�a����[ռ��sW�ks������W\j��
�K>�^m��z����?B	��@��I�$��ߕ*Mv";}�����J.��S�t�f�\ϏM	��Y���2|��_�`hz�c�z%:N��:[X��j��&a޺^+g3Xҵ��?U.��dV+g����^@Xt�sfژ��@엇	�d��;��N�I�~���M����[¡U=��(�,9��ŗ���솋a!�9�hD��86�ڞj.^�,�ː�z�/v�On�����e蘴����^���9�z�l�
5��p�{1�)�@�^�U��L�n���z���vQyu�$k*~�Q����%ݣ����LjG&n��i����E�8ۡ��Ȟu�5"�׌�ƻ��I�`ԥ[��\�T�exl[�6�9ՕRD���Ti�w��e��@��^D;s�z���C�кLJa��{��x��������^��ɨ}���
����p*���3���ŧ���^�u��w��i��vRpO��
YE~�ߔ�mޓ�j�ߞ�2qF�|���3�e+	��0 FU����#��m#[�z�����N�2����3{C�[�����ۊ�&��	N����]6���;�q��=QL
I��i�J,�F瑊�b�����'�DGi0@I �"��#�8�fi\�֚�L��ò+Z��MZXFq>���Ds;`NZ�ac�ڑ����ϝ����̱���M��g_��;�8��4������~�V^���l�wA����D�N�m|�h�_ٮ#*��T�ƽ~HϠfZ�h��$�W��d�v�}kO\�o����B�^m��Ae�_��ҋ�N��������#$|�2,UA�Q�g�ٶT�F3����cogc�Պpbٹ�������Ի�G0�
��@�כkNB|e�O^YYg�D�t�U�Ki[�ȹ���=s���ʫ"�zU� �yU����4������F<.x~�c�1Iյ���,]޶v'��p�����t+U�\�WT\9oU�3�rޯ(2�t�Nӹ.�;!71�d�>�Vښ]�ki�v��sǤT
���,GN0�ȶ�^��cz}@�4�t���!�6��hE�Q��W���;��0��k�@2�0�aS�D�6#�˳e<0��g�[q�a�2�Z	�ڇ{M�3�����#qk���8�}�RQ�^z�"����o�#N���w�~}�����U���<����&���~�׸�}VYL_U�o���ΏOb.߈[�)}��¨�E�����4>�͛�@�0��ڠ����L�N��ڟ5��+�mD��4zci���d��N�βi�'#'��n���(���O�ll�R��r�f5�B�f�3V.Hn��Ռ�;��j�uF��o�t�ʊ�f��.��BL��@�4�T�B>�4o�ř���4M��V��\X�h��o2����x�:��mfd!��kj5�S"�{β4�@��o5�N����^����t��f���ϙ*���ù«��T�7�wL(:��0'!�E:������/�b�qʵ-���OP��0bF�wT�Os:V����
mЏ*\�9��MW+��H�:�=9��t#������㦝��J�e���ww8��/Tf�/�W91�u2ա�&����H.®j:﫺�v��*k`�}R�h�ܦ�FR�u�z�����z��V_�s.��v�ƩX��Ԫ���f��u:�ct��Q��1o̧��K���Il�9w(;c^�2�y�o+�GSw�gp���&:ˋ�QC�+\�F0�8��k��e˂gJ�HS�ԑ�si���S��SGo(vRN��ȁ5�	O)����y�H\v]��Wlݍ�k�_3�]U3kǆ��p,�6Wd�.�
���(�KqqV��H��l)W���[�T���)i��$>ᵺ�S�[K�X�9uy���71:��\�L��R��a�Qb6ЪPhc�|���Mc�\
O<�K�)׷TO�_u�S_P�2V�GtWs*�n(N��Zw_6�pk*�.юU��8��u	�˙�AI�w��vF�q�\�cZ��O.]����ϥ���Aݝh�j^=����BƙR�ƣ��ε}�yҖH��9�z�8� yU�.�5���i��F�����Ǜ'1b��w8�qE�G���a �G*V�%�q��NM��0�w4�0����o���'��V��5�m��I��U�\��V �\H����z���i�|�G~�8�m����s0JU����]����ś����7�Q����|�����:��f+v��;�/C��}�ls�&R�Z��Q(.�L.�qE[}�:�RW��,�Po�٥ِ�+ǵ�,e�.��Э���.r	,�
4e�� ��Txf�	��1Tƹ|�h��x2�3�8�%Qq��-D��.ۣ1E��k�����.J�9�.�}mVYb�|3|��Uc���XG̀�I���eF�X�dכ�j7�r�r�o��.GJ��� 
��<V_l�{3s04����.9֖��>Z/wR��C�1��5�F"�4�۹��eZz����;>�W��1���ۺ�p l�|�l��Q�Xg]fk�,�L˫��$�1���Rۮ�q�ze�P��kw�����U�:gR�;js�0�g�d���u�UG���B�W�-���c�nr���3
ÅY	h��TH�@�����o����9t4�4)�E��%AC��ʃ�w�"���Ժo�#�'�������|ߛ���w܊e�?x9�ȋ3��C�]3���p�4H�
����K��������wo����>����¢��ގJ,��Iy�2�(�%E(�9O<��.�{[�����rs"I6p���Z�ej	��Ib~S��>���J�QQPd�a	}n��"*��R�qu+��9D��AI'XF`�ՙ����0)qs�\�gS�V%l����v�P$�E�;s#�$���Y(�G^�xBr��̢�c�\:��\r���"�0�!e���t������dI��+�i�$����J�u��D�5����R�W�:p�2%j��!�87	#K�R>�H<Y�bаZXs�iF����I9�J&�Z�t~xasDm�_�����w!�ۙ�8\'24��~��9�{�ņ�;��oZ��s�֤응���(Iv/�L3�\Z~��ﾣs1BAV1 DQM/5���'�\ߞ���ȇ�ܞ���yO�Q�F��aTrW<��I�}~J��ͨa;W6u�*C^T�c�ɕ�ݑh��)K����)`�D@M��OEs�����q�i*�
�y���5� ����v-����i$Տ�`��٢��B��@����sH�a1��#�k�еaD�q�]nC1خy�����Y�Ƌ�����G0�z��sPw���#��k�T�涥�j`�P��R:��9p�{ݣ��pY��[�A&�}&�k�j[��@��{�L�w�\=�V��<2���u�E�gcwO(�+jY�9��,�w$�%㝏�2��g���~�V=>�V������^�P�讷��3}�ʃ!ʄv��tz1��j��a̋/� ��A� ��˴��-��-��E�H�KwnP�%����Ѱ&Ae��BO��/��cs ���/���T3�
�-��ts�UF�7�>eQz���z}�����K�����TN;<���s����)�G��:onon�unI�ؽ�t(�oM��skb��!	�]�L�C��lQ�2U'�*���U�h����fč�Y��Oߋ\���j��<f$�cw�@���:���5I�>�ʉ����z0���t�ڞ�Rl�/,9C+�ıg�,ê�����ңz���%��ݒ^���O���0 Q���:������$Gzm�/L����ި؃ �F �b����{��71�m��jo�����L��hR{Tr��=��w�cռ4��; ^��q%�eZne�`l��].������
򽁤�y�?)��1)ե%�j
R4��1��Z����u�����ԇ�V]oM�k,}����^{a�H�I�1,��n�dR>����.3iU���Z��T�����v��V�B�l��&�41�;D��cz���Ȣ酣R�Ŗ7E2��mi��~���=u���%;$޸T�;�ׇM3c?M��7p�4(��'�*�yҌ�F��c��]����j��l&U�K�5'��d0�ty��֘��Bo�EՎ�,1�U�9n��]�N�w QޣB�w:�WC��di���܀��a�G�8u��S�O=FN�MJ�*�wd�j�Qkn��V��ҹ����W�ܳm{��: ����{�s��Ӯ�4�O��;[�t�ۏ�pͱ���Ze��:�	�F>���5x׹���1a����u�V�"�S�op���P��{�υ�j�PݐͲ;%�1�Iz�"�&+��ۑ�a/�W�Z0~Z��)�U�v�k���Wp�7�p�tԷr��{�^���B�0�n��A��,뉗b���~~�7��u�N��)�`T� ����i�':��R�}���u�.�8�O�8Y�����𮱹F=)n�Y�eAȱ�a��冟.��{D��Q��� X�A� f��0 D3N'�ӋVDK�.lo��;l�Ļ��円���J�/�����c#v����A!�՜��p�Új�hR[�\�CB�i�i/����0���,�D���-0��={�/�{���3oK�E;�T��d)m�5U2wz6zS4!y<�PJ�!Hɇ7�i�m�k�<�,�t�Nj]�s���"ݵ�K�R�'��T���%LۆdE��	���^�C�ٵP���t	w��Ŵ�hm�J�W�MTv�{B}u
=78�.����	M���d�њOj��
���^=oV�^w��s�����X�,뺡����a"A�V�y��N*�>B	�/����V*MsΜe�Ab�j�̭��r�������WιV:��25�W�;A�'��~�N�㘔���@�ƁAU6?-�o�3&��s�O�p�� f��	K6��S��v
Gd�q\�a_�9{�R�u��[������(���%Z�a�|LYv���y���%#��M�0Cw����A�^Z��y׻�a���/�꼣�e"�׵��İ������`��k���ϯ���.��\=S�-�ev��C��/�(!r�7���C��k;r�����A��~�3����|�L��9gԑ����sc��U�p|y��/�%n�*L��uh9�e�QV9 �J�����g�+��=�����g�_����m��Cs�3�D0@FDTu�����3]pֆ>�<7[ҭ�e`v����E�H�R��w:lw�%ݵ����b�%��2�y�H7S���"Д>�����:�W:�jE1�d�0}ғ���ɷ��>�je�89�[��iƭ�[�7��wf�P���9a �ö����|�Cׇi�j�Ja��\O2�Č��ލ-}�)䨒ٗ0�����(�1瑱����R!V@��x<p���/�F9l�����%�ٮ�"�9�9-��7u֎�r�^+�W5�-��؇9��v�`PY���`��̔�
��ܥPz��j���E��˼�<x���5�,����1��|tE��x;��-���{
;�L�=u�
������k�#��uݿ3컎��8���Sl�W�v�}kO\�o�c�P��~��l-�)m�T�#��Ao�-�=���-ئ�P�qB� Ũr�P(�3�͛eK6�+dw��k�C��І��V<����s)�u�_��>��B}k�'��%�x��S���艨�I�Dܭg�4��*.m�5���v��&'��ڧY5FB�tX~�k�3L�޾��깝�W]�㼍���:�N��"�:#�)5ÝY��c��gme��,Xk)ՇK/e(�q�XF,WΑϹ/��/��::�Tڗ�n*�N[���)��ڵ�e�5�]���,�+n�)ug��iJ�踞�{ӏ
��5v�2ܢ��1�2 b��*���������B�x���B�{��~
�0�]Qm���\c<H�ހ��5צv��v���-F�j��]�Mx�K �����:�W*�qw8�}�Шt࿅?�y1�_�� 2fѯ�z�ģz���r큧��wJ�˶���5H��Q5�lA�.͔����W��Vd�DY]�wk;�y��ą��`�И9����jGeI�Ͳ.��i���Z�P����z�e��i�X��ڼX������v��8%ݸ7s�A~�B���B�7P��	Ibm���o��a���v��~B�T(����th��(�� &��'��њ�GA�:������nQnMR�Q�q��[U6R�ٺ�ɘ���P���9���,➀N`uH�m�lbf�֐�@�g�5Sij��K�X�=�r��%�ʢ�I��C�ÿO��f69��s�pYJ��6�����LՈ,�Ú����9��a�l�c�����1e�3Ԡ�
Bp���r*��*�Y��f>�	�'��}��Y�:��f��ܢ1%ځ2�u�2�~�V=+�X>'�?*�:~���b�*��%k��7Z�����N���qu���j�+,K�=�t���-�֝~��D�4_���V�U�ΙJwN�e�_���1�Q��"f�}Y'N3��6�K.�<��駘�(5y݈��l���(��=����>�R��7����*b�F(�"���7��,�8��X���E@���C�>0��qu����f�Ȳ�@wH$9Nm��ݼf�猥����l��xl@�f��D�\M	̤�T^�{lcfz�|�^*�=It˄/B=xw�C��z�ך�e�����u�,�,"ä�b�h���Ʈ��K[;���SA)�Ǩ6x��!X�6eAeФT�p�7��:��>�~P'����5��\D�3��⚦�=�7�Q;xL���^��cN�r����L�ѡI�ʎP�=9�C
����v@�2c�km��=�=Y�GU�����:'ڵ����<�����oJ��	����|�bvr޵��ח����6�o�Z��s���C�;;z{�Ru�c�:�ˊT�P������5N���O�e�ᶢ1�}h:�b�\�%�n���%P�>�.�XF�YO=rZL�T����V1����n̻q~��f �����!7T�M�;
'eC�s�L���n5e_i��5.���Z�T5�K�{�ѨJ������(��B�Դti��7�����o�pf�yA^R�)�n�~��0�����8�{Y^���Rx�v��X�R��e-y�ne������T��cNpo��{p=�w���6�b�C�Ҿ�vή�gU�]2��}n
�4�բ]�H+�{H��.V.�H�L������JB�%��N�����}��M�r`�v�Q��0���`=�@ڠ��&�͵�&����XK}��B����Y����K s�����;����͘�q���A��!	��eM6퀪�[%
q��ҹ��W�ip��uW+y�C�&-'�����o����?�~U��߰_�����6��I��<u>Y3�ס�g��C1�6�
%�G�gb�Z!��TgA@r�:�^������>�_��c�^�	F`Ѡ�e�˚0�ΙhR���ƠlC��tK� C���Se�^��$�c>ݬ`�
��kH��E����չFt:�@"I4�>/��o���Ց,�9hjd�{d������,�|lt!���i�ץ�id/3��(Y���*�!Hɇ"�m=y���k�=�憠�����
�iz-�Ye4r5�k���Ҫ�Jz�ɛj�U2~�SA�[��	����Λ�ƚxX:E;��ab&+�,p��Yeq��$!����1q����pn5��q�.�qH2k�i:��A�y>�l�K���qge�^1��<A�l|,;�S!Py�A#sP~��&%�{�Fi�Z�0�˭X��N�2uEh��%׻z���\iY[���˔#ڢ�:��}�� �nn#�nX8<�|+N��)��>>ǋ�0RQ56��������T���g]�X�#�]�WF<�L���z��v�dfm>Lv����W�31�U��_ 4�.��}U�|a��g!��@� ����0���0��Aw�Ny&h�R��2K[�W��?<�{w��bx.�z&#��=�y���)�{34��렮�q+cM�F��`KR�����oP�W���CW����mLpe1�N���* %.��D�k��㲷z+	�ޣY[Ϟs����T����,Q1e����[xBG��D&ەlv�${Yޙ�r�:�B�؆ܖ�{Zf='%7K����e ��E�r1,0��A�Uü�S��39��������\O�᰽m)���U�ga�H�R�G����=;��b]�`}�8/��2��s�C;�
���;tC�3�U�b�ј���j#�Rr׈ɷ�Q�{4�ɦ�$��^�|��\r@la��T[�2N�����C�y�mt^�����i�kPJa�����{̛,f���n�Pw�����Z@/��:�;t�a�>��xB�C�az�u�'�=����}Qx�v�e�q�&͚`HpoG�b�)�o��w�� h�gh������7�0�Ո�SX�7eҳ�(Sn���!�0Ж�/%�A2�Zx�w���9����T<���^:�-��6��	��d�;;C�>�(ŉ� !���@02�A��[��'V�v�N�˲ӺsW��qT	��h�N(�yu�{M�T�͆�<�	��}���Qw��Ӹ�bt;,)���f�stS�K, ��A�o9�u�N7�O/R�9�X�:�@v��(s�e�Aǀ�{���f��4�ýX�Xe-�L[���W8�n��}2�3E�%ڼT� ܌;h�ִ��y��QK�T�S&n2{;���m�ڕ���s��V�yUH]�SP�qe�b�Tȣ8Α��؞g`�����1:�[���;���d�0i)ݷ^X`����U��A>4�q�V1�nTdg5��Y�l[����S�fTZ��ۆk��Iq���תu�>:텆��p/�ST�5wL�����m�֎a]X�hRS%����ƯuEë|g�"z Pe���a'eX.deCR��쨌��*��
��
��5 �$��%:HȤeRN.����$vE�*���H1�٬sXv�Z�˧��ݘ�mEC��!���^v[�a�vҤ��LU�H�� �l�����E�~�G��u�3c����Շ�^�Ѯ�`; K*��4�����b�H��7��z������M��C-��^wL��5�pq��Cw=z^S�I�'A�L*�J疠r�'�G!�_�&�����f��;S[�l�3xwf�wǷ����s�M��y��f�I�0T�`�EP�ZZ[���u3t��Y"=z���)��W��U�{���Ns-ڧ�\V��v�����R�>�35>⚺���3���"��n�a�]�f-e�}D���������z�C�[���xc�F2?����к#�;�?/������vÜ�(l���$ c[�:e�p��f�*a�a�e*�Xi{�֮{p�5ݜ1��>�0�8:�sma��&��u:#7�p��B�؝�	7B�I���Q�'ǬK�_��B��28"<��65�E4t�ơQ�hL��N�.�fޠ�a�GR�StN>��f��5-�^=�׋�g2dK�1{7ĺ�z�U�ٝ��^����nwiĻry݆m �QaDėj�2�u�30��Ǆ�[Ftwj���Wk��Z�=D��!@�����³i�V�:M3�z�]�	L�-B��.���і�-���[^!���B���e�@�B,�|�I�UE��X݌îC�_K�n+�����#.��we)�ח �My�\m:j�:�!�tS<x`��a�q"��{�Teyۯ2L�Q7����aN����n�E�����~�2�]w��	Ty����	��T9זt5��rֱ����g
Y�pش7]�l��0�����`i.(&z�
OaQ�~=9��0�C`���3�i7t�ʝ�s��)�A[��U遼'ݕ�Gb�j~BSbS��JK��B�b�׼!�x4ؗgcC����~$RA��ͮ�8���&�)��pX0��u�ov1^^��~y��7���4J[7��pq}L^ֵ��}SXIKm;�1�Uhw�i�����5�,B����p\p�X:F�9��(�8��F�>W\�d.�RL�� s#��V��b�k6�����Wͤ���	��:�Ҏ+Q�o&�X/�K��4v�wh���K�6���r�׊zJ`���՞��
7�4ҥ�+�]���Ϣ�u-B_gSn
�B�����ϴօ�u̡t��-�ݰ�Uy(X��S� �\9�HWR)ƭ�]����6��bTٕ��`�(�Y�z�ރ7[�.�,35�Z/��m75�3&,h�͗��g$��D�e���o) �(5]V+Rs��/�j��<�C7n���>�FVP�)w�O,�Şw�\�[��;�5�`���[ۙ���Й7�ڴ&b�"1�R�[��� ��Y�Vi̎���Q\�+.�00��q��)��c��&'n��r:�;+�դ��uu�P`\m�M�:Ѧ�D�\S~̫�љթ�����\�1��ޱ���t�颯 �i�[�ʉ",�!/vM��-V����h�eeH|7��vl�L�|�n;rR:�IA3���k�	����kNS�.���|m0	j���ғ ���E��]J۰�?|N��`j���z(�dPogn^�6�w��ӂ���fh>\/�y#R���9	��,�֮�V�̩Qr��_1 �͂/��X��V�i�2�>�<�*u���,AU�b��\m����ʸ�:��6��9�7�~C�]j��%-��^)�{w���hb=�th����W�"_b�@c��VZ�5P+G`��8�<��2ַ֗t�q$fԩ�w��t�	h�(t�4 ����j3��gq�5��Hm^M���U.nP�=�v��B�ʗّjv�@v��z!뾺!f��Νהy�o{�y[�c�_f��^�K��z���n-/����t[t���O�z�];�+���a6gv���q��
��]=pSY�������Bpٯe���s��\D���y�	�ʾ��Z��W[;Dns��"ޮ�[����"c�J�Z��hϡ۬�c�Xm�g_��&K�>�OpD��#jge��R�k�NU��8�^��<:�����¢�M	��Pe�og�]1o��Ր�Ž�	&��~���`�3�!�,��U�'�i	V��(�tw`@�y����$+Y���y�����@�!ĳ'[iҊ�R�]�J�ߟ;�AZ�2��Տ��v�SY6�Fif����`���d�6gt-���N���@u�h\Cz�j��ל�w�̉J��7c9
Ի��+�º���9�n�[����]��
�y��SY��[�:��wx�Y��trd���b���q���P�֎�ʟF�U�5�*	��h�F�V��:FM���T\�Z�b���B90*�{��W���A��VZ�s�f��q�9gs;ͩ�����TPM�����������~��⧺<���r{��؟rE�Gߑ�?{�JNUh�;C2��iQӚs*��v$�<s��*'jl�坘���!	����������$�K:hXhʠ��(��24��0�J��Y�TXdҬ6�J��w��|�w��\N\HN]_nQw:���� H�d]�T�s����A�����������#�^��I*9�e�8r����#����!;�©�!ɦ�������=��NN{��]D(����rj�$S*�+7CD��G=�狮��8DU.�G*�Z�M\���$9��r�8�B�⦅�.f�ue���ѹ��.x��r�����"�Ef:r�q+�.�Q��wn�Yiȸ^y�4��vAj�Y���u^�Z4��%S�aȋPЫ�h�Ba'*��Ξ�'�^s�R�ē��H�W�k�d����/�p)̲@�EZs�ͽ��y8�ȍ$7A�puC�(~Å�b)P�^{����5f�n�i��n�������81�z�V��F�)�M�;���Yl�������fցg�'P��a���h`T,�@����}��a�6� Urm��< ���o0���+{)�Kƿ�>;�al�y!�y�hOa�H�I�1�d�`n�e��-�eѺ��ӫ[����_�n��4�T���+��>�;D��a�(�a�P�Stu!v��g-�7�c����lS�N�F9foװ=43cH��O�ꀘ�͠{�K^��%�+�?�AN���W~]h"ˉ�����^�%ߚ��w���G�M�"8F�e,/��fݸ��5�H�|{F��֥�h]�Ta����+��a�^0��D+����KEt���T���L?u�wXs���?R����%���8� OJ�T�/a\sH7rʹ=�l����E����Sgob\�!�R�-ǃX��2�9�����~��WC�L�u�q��Ǭ�g ɽT��g6D�龆��]�����Ԝ3W��!�h�]�1��d�@n�f�����1�I}ݸ��-7�V�;N�E�|{s��hz�m�_vS�]��0ʪ%�r�4>
,�mFk����;�nf�Ԗ���f�+>�,�di^H@"GN����b*�dK< �����l��
v�Qd�g����#p7WI?͊�V]]��lPz��JlĆ����`s*a];S��'�ܮ�e���?�}���=�Ӡ����������Ї'�<�f�$����/u⼢�	�H�:�Kzftr3��I�h�J�⯳S��_u���W������;89M�<�0����uWJ�*�c�#2�Y��}%��
�R2a���'��6�Ӯ�Ut�0"��O_疍w�X�韟�o�s9}��U>���٥*f��(2�jm�b��}͛OX�o��P�X�>��}�tC��G�}瘸�����	\�W���Jl�(2j�f��TgP����/��?~Қ��_����(d�R�)�γX�����ul�(F*���'LK$�*�f"(AsXл�c��˞�jQo��L����H02TIvl���&��iH����^X蹜�s3)g�Z^���O:]Yp)Rkk�u�5ȸu��٩�(fΘ��hG+��c�ec�H���؛�[��r99	�)?9�NP��Ԡb�Ú��.���<�l  �0�e���=ZǤ�yx�����&l�,�jOgT�t�/�b���N�P%�yH�Fi�����p�eg5g5W3��G7�\�UP�^�z��UC�϶s���Ӆ���h������%��BlwQM{�q����˪ȿ��C���������<ò~47��˫�׌�ƾ�I��&�oZ���~Ø������ץ�_���R����io�{����&��p�L��5v2(:��:�fc�,�3z����"�'�k��v�J��rNx��u�w��d�}ٵ��0�rD*�T�G̫w��v���9�j�mIx�K�/�w�߿�?����w뾟῀�g8�p����rm���m��}��������������̳
-ݘφ���~���OC���hZO	�Hi��f����哨������E���GP�n�������/����<f�?!o����j��K�����|�����23L(� ���~�3�e���&�}��ip#+���j����v��b��7��->ƫ�ywPny;��P&h�Ÿ�;ǘ��ge{U"_�-\��&(�,��7򦩜E0b!��4���u��N{����i�+úIv*)�n]��Z��E�͙
d���n����#����2�1�=Ų/3Q��ݬlN�qE�nbU�t��Co�`s0�/1��Yг*�yJ���*�{)������m҄�f�ζav{�u~�u9Q��x��Z��rL�u�X�Z�^1���T\9����A@��d��S���nwuo۱,�U70ox)�P���۾��b��F�*����ڂ˜jQp��3���Pe����<�45��;m�]��p�`��^~��=��%:�$hZ��JN+���e棱�C��E�V��W�c��Kn��V.6��/�H��6mlרVd�1Хj�u�=/���8�X��2[=9+0��+�=�x��}�دn�+]o^��ˬ]���V����>�若�A��L���Ⱥ�5Ss��f��~ܑ�"���[6���p
 ���C.�\\�)�\(�[�	c>Z�4b���ס��+ѡ�r�m�ن��F�,�	���"��D�7�3e��\u݊�?6X�έ'�%���`��\:�@L9����3�����b�H�mT`�B��iTDd�[�^�l@k�
���z霻�A��v!�_��?W��
6�aUe�+�[����[)��9\���l�T��0��٣rC����M��7��u`�гz������+�t�R%�/a�-�k�u}���˺��HK5�
�uc�%��/��Lr��i�ϔ�5Y=��H�İо�J\R���\�/d�I�_�h=a���r�G�|1?Y�!V��:Z��|�����>�0���%��:���q�Ӽf���@��3���LOdG
2��b���v����H���aa�;�ږmN�wK7H;�XQ1%ؘf8�8��_t������n
<.��(�olE8\֮���yw�����]��ٹ�Gu3�dYx�� ��{֨F*�.��Ѓ�{�s�L�H:"۫�ohlg�`L� ���T^=���5{�ƥ�_oS�$��h���$�١�zf��.v��ڟNF�I@�f^�Rk|3�g[
q��^����mx���c7�����b��[�;���Au`․c6���v���(���)��k���:���p,�\�C��y��fr4[��݉�=�j�s{�m1h���}���~���8Ó� 8v9@�q�vl�m� ��q��j"�������6�����C��W!LϘ>��m�WL\:��a�q".���v$��b���C��QsL�)^����Yt)X*�8zޛa71LkbY�t��e�kRj���s�m����8�v�����ږ��%6_���Z2%? ���zs_iᶨ�6];�Y7o ڻ���L��S��ʘ		�ex��v)�����ħW䤰MJR4�}�e)�x�����O�F_��a��@j����5��f���O�n����,n:�q�;l,-c[��n�j�b����=�eJ{��$(fɈ����(���Tz�V�.����6���lK���aa&ܵ��7<L�;65��	��n�ԳyU:�U^{�|m�2��)��](➗�Y�O�~JT�~j	Ļ�l�?��M�b.�%(-YQ2�^un6��mjby�y�j ��c��Ab���V��z sIzp��[i�5�U�ݹD̊ʓ�N�Xɩ��0m��ښmV:��>3�Ju��.:�=�^��\sI��m�0�fYX΂�h_��o��:�g�9���>5~5	��I6������X3=�ci�J�n��g"�LL�"��D	��S-⯰l�鄩a-���_��s]�Ҭ�ݧT�ʝ�T��K�eH�����۬��B���`N4z�����������̘�L)��Wd\Ce��&˃�?��߯�������C����O��]4�C����M��*�OO�L�u�J��P$^�q[)�1�2�/��J��C6 ���0n�����y���6����
��l�����v� ��u���}}�8�y����ϰx�b��!��D��9aC�p����f�L����3�2�w��*�tŠچeci���0� ���C�ڳ�J#��L����b�5�7��AP�z�U'k�@]E����ӻ�����zKee)t�p��I�sͼ4��;��
�2i�鞇u�#R�d0֑N�cП7f� ԕ3m�2�*���	�r���'W�]<�4f�k2������:�K��Ô����J�`��v+��Bk�(2j�f��.��sti�`�f"�X+Qx��oV��m��8(>���� ���#s7:	�3X|��<�,�մV;�*Qk�Y�i��J�[�S�`�ΞE=�ă�vl�0�)�i�1NY�l�2�(�T�oM\R�-x��cžk�ħK�K.*Mmb:癱�s�D�ύBR�n�zxLji}"����FoQ����{F��=h ��L��0�,!|�&����Z��ѕ��\WW�;�S,��'e8^�i9���"{�U�[ǖa��q�Z�]�.�*d�,^u�B��7e��A�fFY�2��-º�H$@�U��.;9C
.2����x�D�V�6}�.�$,�'��$�^S���R�1Qa�K�}|�>���s���W�,[˻��;)׾�F�brSQ{:�A�M��8ŧ�P��/�������3�^uiN6"�t�tXt���9ó����������E��������޽�覉U��?�����g�N�.HgA��Us�=̟���EҘ���j>�wl��h�v��b&'=*�מho�ߕll�j�@���@���G�Z#O���������lP�Q���ʺv��w�)��+Ϛ�MG�8U�>���GP��DP�mz���3�P����7�p����ѢV�ܛӲ��PXh?-����0$87�b���nZ�{�9�C�;,ji�a4�;e�I��Y��_�H�J�;�79�2#A3Eڏ��b���:��<��Lxc��v�Z��5�mwRCG����u}S���=�2�3E�%ڽe8�d�v�����.y�ia����v�q���w�
�� a�������mcH΄��.�*�Jw��/�t/(���t�7��YZ*h6���\�]�(C�wcڊ�o;�OtkT�,S��S�%�
av���{����{+F9�����w�:1���]&��K*�3l����up`�W���:No6V�(�JgQ���`�n�8~yS��_��&�CM�(� ��oy���j��9M��C}�g�6m���Ο�]��!'�C�=0�3r�bUk¬:��M����E=�f������.��ʁF���u�5eEÚ��P-�'�Y|G`�`�����sV��~쁮ᝮ�4�259����X�hR�T�SP��X�:�"=
�ϧZ$P^a�\:��;ʏ�ȳ��g�=�ݡ�jBc��B�vC�s7:d]y�Jt��J�␎�a��Йu�y�w�Ƽc�k�xz�sy
-�s��Ð�v��=��s�Gu*L���X�t�O^(���'�kX7׏e�o%u�2�t����|r<#��v!?d�#�}}YWa�i�)��E���v;��&�$�8�c�6;H���2i�u��~g����8Q���!����?P�4(ޞ��{1�C[������-��5e�V6�����a;�h)�qq����Q /�#�P��(��*�;�S�\뮱��y~yu\nGn�U�|�/����­t�)������}j���\0b[���ύ]X�ek'v�d�cwXemk*F��2)r�Z�t-~J	{e/�~m�O5[�w��.�/�Lu�*��fRSi�ʱ
��a{}�����$���]܊��xJ��:ȳ�*<{���r`=ꠚ�3�o���}:$��y�
ʻ��3fb�nM�ӻ+��ֵ���e���I���w��ٗ�ת��ĭ�%�d��zv�s�/�]��_�߿~r�������||?��L�0�3��vr`S\`������������qf3X^f�`�L��z꽵,�hv�a�GR�o�?Mk�&�x�76��e�穏M���ݻ���
�.�P����c*Y�u�%۸�,	x.�L�x@�'��m�/XNΩi�P�Rm�`5�vO:�� �g�#
�g����Z����� ��1�
�5�Z>��a�#`�^���Bt:�i�v:�`���Z���M��~4s��jExlYo�s��W���~������,��Bq��
�W�5曍�M����s���8h���i���N�myY�J^Ӫ��Mq0���FBױ�eAeХeQ�Cy��c1���2�%J��0L���M�^��Q�>��5�w�+��nj�Jl�!4�Z4)=����Nk��1k��OV�v�������ۇ=��_(	����ا������ħV��18�yI��-0�37��ų3��hG�	��z/��^��;Ǥ?��d��8!?{��#�פwL����p|�M�N*��.(�����TR����y��׵��H0͎���r�v4�K�sF���Џ�ʉ�3ȺB�i�(��ˀ�s4W1aɼN"Z��'e�h�.��")a��K]`А8�r��ߴ��Ȫ,Y���i51�Y��D�e�$[|9�T�,��l�[I��˛���^�G��@�`��c�y���֩Ǝc��>�_��������e9@\� � �0
��Q�[��ч��V>��5(���.��n���=�7>�|j3kH���m�g��],r�;�Z>���sZ�B���0���^�ŧ���T~n	Ļ�l�a��k�ȇ�	س]�-l����za0,p�<Uu��ꊺ�K sH/N���Uj"��j�D��i�p��L:C�g�@��T6��U�QkeaJ�a@���~*	�^�+�luGWcL�^�'7U�5>�j+�`�|�0gt�,Iz�Κca۱�pͱo\)�����=�3*jw��M����{5׻#���<��Q��H�����y��|/{P��uP�]ר�ܜ��R
�����{�h���n�N� ��r��z@:"����}������𸘕6^D�0����~*����g���|h1�������D'��i�[�F�T?PȖxBK(ͩF���E^�&�)em�Խc����=�����������d÷���m?4S�:��s`rWSr�$�2��	M-#�ƴ�22j:*���@nL�jJY����SlnC�V�;ӭ�YS�uw^\t����׬"sgY�:�\��r�3�w�R�wf\��5�@��H�u�o�۩X����ƍ]/�xV@�8���q�X��<�=���	�~Z	�6��(2�k��"��hk����#�t��Q6k�$�hѼ�+���GN����M��M.�f��/V[��a�Mm��iuqS�*媊&uo)�����:)8�`G�=�)_md[��q�%�o�a6��y9 �ӃAa�)^�m��Ҟl5�D�I�����E,�jlL�4�L�ؕf��^����1��P�sl��Pɉ�O�Tˢ���-M�k�G�ȌK~�*nCz��8[�5���ȯ�l��mX`Et�����%�J�Ҙ�{��du�f�6�J�H��s32R�e��F"k�t,u��*����c������V�����U�� ��D�|����QpKfmZ��+"hL�u��#ҭ<F�
�hQP���n�H;�F�#s�r�_�X��=�BZ"[�۽+:��k���mSC�ի�:1�Y�t������TΞ�ю��R� �q�`5�|#ʒuC#����A�T�o��W���B� ur�Ώ����٬v
������U�mT�4R)�Y\�r��K�4�N�WiFIV��4���+�Qu4�ڸ^35GE��_��y��F<1���W�!y�֐��i���M�v��ʱa��m'܂]����ۣ{�֣�3z�vao���b�:�9�'2��A��b����,;u�Դs��ؤl�� u����b���.Y�Pk���?8+��C���G�:1���sT΋FP�	/_iSy ����8��4�	3/��O.�1�O��{��
��Y91usك��w(������7��ʓ��`œ.{\���XJ�H��=aT]�{��o�r˶�:�9bb�̾��Ǟk{
Ր��!��ɾe+����ox�ҵ�"�Q\�1���ȝT��w��"��]`�G�{�%��]�VWH��[�Ƨ�b��{�`�g:�i��LذFh�;�b~T�{��}{��f��12Y�*.Ǻjd��Ga��Nb{Y�r/F��:ɬ΃�R`Q�c�:������� <U'�J���Z�1S�7�]���D@�6���V��-��{$��m��fE��D�	�(Sq8����@�K�f(.4v)GCdK.����Wd�#���4�
����H�N��#}P�%�	��������.�۸�K���|8ZyB�h�x<�Dɶ��^淋,��K���(��II����%�M7��OR�kE@i�{�G�ٹ��4p]���R��B�Bt�Q�Wٝ0Q�ٖ�Uƶ�H۲�)�i���
��*�#��Z��9ld�U.,F�we�%R�,֞ѯ�5���U��KE������`�t�/X�;�-��y} �WY�4��'tX�\��vwgI�;����u�T^u�s�͙�/v!�l��uV�hQ
'}V�(U9aV��r'*�R���Q9${|�����o�]�U�NW�ww��M"T�{�����k<�Qr���o������4T�C3�"|����dgN����-/#nC��&��/o������~�M|�rQ=�aGf��t	%�Ǟ�Qs{�'9�R�Qެ�9C��������+���rS��Ҫ �x�U��d];U,B�̫D�r|�䟜O2�{�5��"uoS���)RT��^l�.W�c��w{��M2)���y�I�p+B�+�$��G�n�xs�ZX䇕���{55�"�t"y<I%z�E&�˧�<(��U��#¨*�r#X�Q9�Q�p��<�	�)K�r��G�."--"H&] �0����.�U.R(YT�r�If�}C�$�(|E��i)�v�,��+��9Ĥmg��}7��g�����\�+��g ��50�fJF�W}��߯�����_����� ���L��L�8�vr`��������������{�-��j��ȷx����q{q�0�%�N�zxs�)�ɔ3�bN��˞��2����8E�з�xOB��N2�D���zdG.���s�v�8r�uws}M�kMl�)¼�mOe�V�Rkw�{l�Ξ���H02TIvl���>մ���/Ik�d�f��!�r/� �%:O�bS��%��'��X���ȸ?��t������x���U�ۆU���}R&�K&l^�!�|�]��vI>�	����'+�R�TXsQ1e�ϭF\칡9Vf{�R�(?��eCn���uL4�[���^��)���E�vM^������wW,k^�,$�r�����G8vvZ��n�S�\�E�H�R�'V^'&bi���6��1���V:��kߊ$MX���\���D~=�]%Nuf�SMc^[���R�"Ö�|s[ws[�6Q�a��2m�T{ U2͚��ͺE�G�/�{Ţ4��㮗W�<�3�j����5E���B��ʀe:�^�OO�oƫ�|_�?��C�O��q���<D&,�/Z"�hb�K�c�ݒ�+���Ɩڃ�6t<Tp,���g{<=B�%�y�!���dX#�Tu��E���d�e��\��&�ӛEgeG6���St���87�b�orK�����h6�6�� �f�,�^�ܹ�ۖ6\Q���j����}������W������dw_�;g=˶�2~;I87J��D�EsP/�ܵ�}'��&�-/������NNfaR�����11��ޱ�Y��A�4 ���&Y�H��I�_�f��`]=��*h4���1D`�%�P�� `q\��)���m�8;����i�	�.�T� �B��,���\�t��eN������l�w��Ey�ol�હ�u������!q��OÝE��#W���IP~h����ų�l��Ս����K��qy�y��zap	�X8���c7�7.t<�Y#��s,��ϭx��C-�o�������j�?��ut��e�=�ځ��7b�ꈷǎ���Kq�^Jmj���^~�c�1I��4)Z�L)�u�4s�EK���{�ՙb^z�*Оk]wUM�?�����ir]���M�A�$�ħV��j�*�qw������>�6�N�.�Κ���q�cL9!�C��f�7vl�Ou*L��`&*��"��,�v������!9As];�0��=��Ƙr�L9�C,� T7d�OO�5c��~�0��n~���ee`� n�d�P7].�Y�v�gV�X;	��N��^���7ƣc<�ۖ;�e��&M�7_��ӊ5q*\�sBR(�Yɀ��1����f�o>;��z�;��v��"/P��[�ze#�PY�8��׮� �y�{F�X6��%M���_υg(��9��_���}������_~v���2�xOm�I��؀�o��^|!�n�yO�����=t�uu{�z��근;۔�WӼ��jy�������_�$��h��P���~]��äH{��c�}U�\�أ��{aD�qd�,)lk^WZ�|^��֯�!C ���\�Y�W�W�)2�h{W���`�k8����Pf��"� �V��/ҹ��J	{e/�7���֯s�w�/�5LTSţL�� ����h����[R̶��Ø�R	�~��%٣7�Ks#�^�?���B�M���a�]g����|�K��>�Y����R�2No����rKėj6�'#����ky�m�6�vL�I�˜S:�F�Ӽ �@��^a�>0ب�G���E2l��#z�Uk^��D��}�i�pr\ˑ�c�����463��B,��̔��΁��*YYMAUu��hl�p��-�i��<5}�U�B�&��q���1s0�tS;z=��?��HY9[��i��p�П\([4����T�ӷ��!k��2���R���ދ�3*.���!�s�@v-`V�b�~'��y�uo͝b��`b����|�*+�r���o��K�Q�%��W�w����	����}���du����\���ي��%�����U��lBm�sS�����vrٯ���-EeK9���C	��ai�W���a��f�;Pԭt���������v�3��l�sk��M��L���)=�G(\B�g� ��ٴ���Ve�ek.�Y�x��-�`趟s�O��!�vW�i�S�܄?��c���թ�.��r"�Cj�����ǯk�<�o��!ݭ�:A�	������^�T�'V����rԨ�5����ܝ`n����
T�1y.� ��k�D��"!0\��7?
Lƻx��,,���Sy�p�_vNC���,��E��U�F���r���wv-~(fƺ�7�!��������������09�BΡH�q&�캳�kJ�%ߚ��K�k��
ثw~���&�"t�ێ�νi��SL�<]0X>:v��RaϖGs�U#��� s3���A�Ҳj�աd�u*�B`���@p�^��S@6����vkv�V�V0�ҹ�%�]��l�h�f��#T�eֲ���[3�3��@x ���ͮ��<??����α�?��Υآ�'�"���NVl�u�Dsi�b^�<1�����x!�y����d�m����.Z��+EL&G��>�d�Rɠ�W�:U��-��1؍���tO ����͡�=<�H҃�~��>A�S�A���.�*�#A�6���7iұ(�Y��܄��7��q��6�ӻ��=D���C5ۜ9BN]�#��Yf���;����������|�������&s���/���Ӄ��/�z�3w\^9�c�>�$@;\b�}C�M�5�!���x�����\?`���E͵��۱���<�����I�č���;���H�F�q4�m���Dzb,��If={�(}�o�ϼ��n�Wz��,��v�����g;�kH��L�^�X])0���m?t�9\r�n�!�y�<����ӄt����|�U>�}ȊmIK6/a�W���	�{H|iv̛��W���3q�u&c:1��7:E;�[E�E��q�����	_�b�#��]����4OY� ��YucoVd)L�:h��3�(�^=[ռ�|wA8���" F��C�m�u7��S��{�ל���`��1,��Fi��(NK���\l�&�yV~5K�~�9;�
h�a���!,��ޠ�S������H�TR�����"��tx�moJ��p�e]��K72},�S��]���&H�I;���%��jŗ؞�N�4�)uڱ�x��y��p!�^r �И��;��E�S>�M��Z~X�A.�M[�<B�z����}-��`�u�H`���9���q?��lg��v�����g'du4
�����I����'.�X\�E+`��:��ʙȣ�������`rv�*�	T).7{\�6�rtz�xrA� u���[I���o�QC],Z��������]o7��7��Q҉X�'!�y��%�XE�3�
5����^��M7X�U�v�E��DcŞ�,�-�sۑ-���z�O���v�61��x!�:X?s�;'�]T+�X5"��T2���zӪ�{��޺=�u��[ܩ�:7��{�o7�S����a njz�
U�=�����u����������~Qn�����5���zG�oƫ�A~����!ۤl0C��՟�o��ٻdI���]~#�ݮ�Ͻ�C�x�$���s4������S��Ǫχ��F���O�#�ߣ���p���e�d�����Ƿd6��Ώr�� ��`puǅE޾���L8��"΢u��.�V�o��߸8���	:��8�npwO�� �4W�t��0�WT�* ��@�����ܫ3�_�'M�qvW��l�%ӯ*n�R�J��nM�*�}]~ݬl�H�!C�E���DVq1��^A��*���|ئ[�-�<�zw�\e���@��z`i:�)E�ћ'�8ߛ�q��ּ0�H72(�3�u�5{*.׮2	žb�pt�ߣ�{-n[� ��J�+�x���7+_6�<�����^;d�0fS�>�V&S���\j�f���:�D��Rgz��C��6C�6\��t��*�,DP�7\�u!�t/!�^��UJ����ˍvW�ԷP|���3���9M����
�|>�������R�}�z'�s��bq�|�u�P����e�K�tF#B������A���?g���  5�&��,m~�-`w�G�C�q����~'�q��$��%:�.4-X�I8�7��)���9�YJ�v�X�)E�ex��	�Pp�C+ۗn#s�Gu*L�1�����d�K��-¶ؾ�;!������,Y{w�xa#r�1���'uy��7�%�a�g�c}�M��7��i5u�#[Z��/fͷ'X��s�"�6��s�s?>l��p�7sԼ��V��������j��1���ޮaTrW<����R�nH�C		�ݚ7!����F��:n��R���]5�ؕ�x7��k�Br+�oʮ��$닲U�9��+�a%��Z�=�x��B�p�^:��~�<�Ż��]{�[�^����:�G>Ǉi�j�J�e�W=�����G0�z��`����3�42�¦ȼ�"иX�3h/�P�ږe��XsFG$�5�`�ft��4Y��s�3�����V��֠^��̙� p0<4Bax���ʖe*v]��g�A
;_�X�1�NJUܢ�;�ݼk&��h��T��PN$���lY�⋞��qhw+�S�G0>6��)�4�;�wJ���?��g�m�t��d�Վ�d�;�~Ҽ�&Ȳ���xw�Ѵ�@��cԋH��o��s���5L�7_�W�몿������ox3xJ=�;7֖�)�o�y,�^���H:"����^u��0&tF�T�'��s����␚�x�Sr���Zf
�/�+��C�*#��iD[.x��:�p>B,��������[�7K2��0��n�WN�4�|���4�28���� �x���y^iN���gF��)��Ѐ�|Wo�����)��5�]��r)�;���km&��a�U��J�Tu��N�t:��E��U���wiQ��'��rk�g�DscO�L&�C�G;a�d�ӵ-�O�Jl�d&UhФ�+B[|���/�y��.0�C�xcռ55���
-�8��S�HWUx��ا�����p6uFGQu��79�E��H���X&�)P��x�5�ׅ�;����t��L�cFy�|�=o1���.�VG^ik�^���}^c�:��U�R����0Q	�_Z��1	��筲�nLa�-m���=�Ժ����'OC�dRt��]y9���4���]�S6SLNN�E�tiGd��:tBf�C�bmz`k�T(�;JQ�=/�b��$��%ߚ��I��BT�yw�`[!Ne��vrYX�O��}���^�7#ظ��Z�}}�������$�}��4��]��1.�˗�O(+V�5����]J�z�I�u�{����Sݴ�G�͸��^qb��������U˱ήs)�w8$��4Q�ɹc@y���M<>��x7����i�!%��A���=�>����Ʀ%?;0ef�:rEh,_ʌ=,��U~WC��c�0�'t�\�j�K��ÿ��4��h��Ю_#G������~���Z������f\������s.�]�����^��]�6�����P5�ʏ�=�@�ܿ������z��?m
 |���Y��'����
��dϧ^���P=r�_�f�;���p�0 ���ξd��\��x�f�ë��rћ�ϸ�^�FC1��K���=%� ��+�tF[6�;;��^A�f�(�6Ô���ֹ��XO.7=�j�5��h1��X��{���	�e�<_j������>0:J=�h�֛�2{_�:"�Z|8t&�{nO^�ǳ�����w3E_I`J�hFL8~y&p�3Ks�:�uo6���=�MC���No�R=<�7&m�j>ML�xe]a��e�;A�m�v�O���Xk/Ô�͛�cռ*�S��a�y��OB�`�N�x�����5���N�M�6Hd��Fi=�3�=w�7�ྲྀ���/�D������6*�˾Bfu}����
�����Ike�����w֒���Dumn�\*'w��rI��=vWתt��k�A핳Y�۸�	��w�i3��i��e.�'V�K%�[��m��vJ�/�]g#��[�N�;]\=����|�����};������`��Yy0�7i)��>�I�� ���:U�b��I�[�o�@�����xŊA7��OZ֯q�jzvjS�4:���4�'�1)ͮ�L��I��:皟"������h�eT�t�kΧ��G8Y^o
��A�fژ!��K����0�{��O�b��:���摶$��י5�IM�.�O��2-��r!6И��"�W5��yLG�}o����'$�	d��2|��Ь{��5�L$����|�F����<2ׯmt�u��潕����f�䊬nb;�]��^�4�$kr���>;���v��ga��n�˽zdO:�UK۳��E�cU�Z|B������2���`�̨��l��wf��`�C���L��P�jS@[:���3�n��__mq�h�&��3������U� �X|�
�X�n�`��Q��©�i�Q��Π��P�d�!��=mC�]����x�)q�9�`Hpsx�s�NZ�/oP�-If(��w
^�	��N��L�s�jF2V;�7<��hEx���@,Ÿ ��#rviPU&dKPý&��E�=��4�bc>���W�E�ITU�c3��YY�&�T�zX#�J�E��܏��-�F��XAJ�I�����&����Ho\:�����Is�욗q�6�#z=������n�X���;:�Y]f�
8j�v�H�bc�Nȡ�Y�� Zk_Wb"�|��=KE�0n�jT�.�ët&��`bp���9�M��T�*c[K�>�b��n��[*!�a<,Yư^��ᾷ��D�����Ɉky�5�0T�R�3+{��V�Cv���u���ʁ��sGh���>-��!�DՈ;^��ݷ��ŶiŴ�@�Co�6�_0x.��
� F&�r��[[���|�1Q�p3+3#����O*/�;+Ǽ��>^a°�B���4����y˶�a�q�7'ҝ�_:�3(���U��3�I�9[Gy�f\|�[SN^V�u��[FZ[�����v,|���Jv�jW)3��F�,��������}\�0�IQr.�FŔf�IW�1--}ɮ�0Yt�a��I]�7������rhQ��]���[J���]��Y(<2�78g/�}����i��im�֞Ʃm��0�.Yc�O�B)�^IO.n5� r��A��B��^N���%㏻:��\�d|r�X-o
�P,}�mj��Ե3�0���3u�d���HvYi�9�!�r)��롑��^�9O���|�6�$�:\�h���n�]��d:��� ��5�C���v7н�	�^G�Y蓫t��X9����ł�[v��@b�wl]1VҥL� w۰�N��x{�ti��z�w�O>y�דu���W���(w>�k��OB�=�����	[�W+�CP��)r���pt<����m���t����/^�4{�&�Uh����}��Mg|�-)	78lv�[P��ؑe�ԄSS�=��\���Ǳ�#��>��oE�D��Ikf�X�� }jqT��������Q}��κ�����d!�����6QdKw3��jw���;�I9r�J$&�v�T,�*������x�M2�yk�������Z�����H>�'��c��XF"��A�룂����hf)m��q܌r=�ۊQk����ۦl�Y�����%�U�0��5�����&�d�G6�m��9���.�!$W��6ls&,4����Q��Y�}����t���mؚ��<�|���y�;u���g�ʻt�LЮ���0�z�Ʌ#�K�S����b����c���e�P#�
}��;�9o^
U5�gN=\]�[�v��Ѱ.SS[Qk�5�k�
�sXyL]�{���j �<R�(�e�K��s^����a.�ͻ�ʘ�P����|U��!����w*�G{o���v=�,��Ҹ�=��-��٪]����l��:<s�^�ֱ��U��њ�`��xn��Nt��]0�g<�|YW�/����)�y��D�^�S��|���W�����*y���|���:�N]T�����*W0�Qk�D�����o�������F��OH�fj�ӯ&.EC���2I�G^�fb�]9,��KI,�������~�ER��f�rHJYS��Ҕ�]�Ve\�K#C�%��;��;������O��D��vdUD��q�����XEu��r�^�x|=��]����w��|�p�}�����^�g%�����R@�r,��j�����K3��/A�L�<��9��V�{�YR9�l�]��C�zUQ!Z���!r��t5$���Nl�H�]�Uz�8ŕfT�G����(�K�;�EjH�$U*��j]:�k5Y��aZ����y.'���/����OZ}b\�-��u����WR����W	����^�z�W��u�* ��\��i�nnB��&�;�Iu
(���̹\tB�U�n*!ϓr�@����fq��?T�Q�V��B��M���͢���VV&2`�ݾ���=��wKT#A�����s^5L�Ž�]ܗ�~������8�&�_�`�ˑ����(䥦�¨q�-�z��l�w�Co���4��N�uN6۞���4��O��z�q�7���)�ey6�1&�Y���.�R��P��P�?R�J�����ߤs�vyO���o�������h^Fpzf`�-@����y˲���z�`d���Wc?7��V��}�Y��TK��#�ȫmNB|n�A=,�,�kY����5��.��fj3�o����-�HE�pW�+հ��L�c!s�� ��1I��4)Z�L)�.��q-�ݯ�z�]-��Nf�V�q�H�o@0e��L$� nK��MͯЙ'��%:���k��ͬYf��<oO.,�*e�/GN0�r-��1��c;$X� �O�GPu���t�?ѝ:3]��S�'
�%��m�E�4��/A�-��@� �cH�'� �{��L�	r�71�ȹ��ջ�b��2�S��}���"�x؋@�f��ߙ������`�݈n��!춗��T�.����hЭ���
�J疯Y����%%�#�'�����F�	�����#[^9��s
��;5C�� �	��P�35�gk1>w;�4+�f�f�T�y��B#c�Ӳ��k�T��ƹ�9:���T���^;�ԼS���J�ݦ�\�@�������r�}ѳ�tŁI�W���ك�>R
һ*T�.�ʼ�v#+���<������{ƨ��,B��K_���ЕίƮ��$닿���]<�l+�a>/v����ے�ܹ��Jl޲2��X>�g��=�#�k�е~Q+\qn��%���Ts~�%����Q4YEv�O�S!oa�'(f��0�ږe��E�5J���4��]�4E�g˘���(��L��s��@��^�9��w�\=���m�_���'W�,��,�VS���ffz3�����bS�%,�^��i��ƽ�-����0�� `LЌ/0�vMn2�UX�5�D����D���+l��i�@�i⻤���O#.�C�.x��<�fq�听�O+&A�$N^Vl�|�T8P�Jy��zmǶ��D<5�_�W!
��H m:j�L\:ض9�O>h�|��	n�VΤE��p}��5zs&��1��&�+S�As�t�t)'9a9�0Ѧ��u��nnt~s�a�|O,�DƜ	�C��iϧ+�,$�%6_���(kװN���C��{�c��t2�UC�\������
�^Vߍ1d׽[�~�\_�^)��R ��+7i��$�\�g;�m���ٹsN��[5����ݖ����խ�ˏ���X���w�wt��e�T>��wsh��5�jY<�=گ�/g.���j��ig,Y���ps�e��/{/�f�.���qQ4{��9��q��������{���Y\r�h�U��S~ȝu~*Kԥ*q�x����i��Cj	���'���je���Sۇ��0!ە�̤��IϗE2�R��W8k���� f����(ӏ�[�٪�0�u.Cd�i
Gd�y�E��5(���M��##��r��]cY�Ţ#p!�Lc���7Ak/P�f����٬(6u
Vv�88|���'z��IAc^��.�ܯ��SKt���%���-%Ô�<a��cL�!�:����;Vл�F�F��6T%���1���V:� ��=8}���ǁ�:|tz:��ښm]2%��7~qity�l�l���w5�sg�]�&^��Z��*�X���Рk�ʗ���O�~��m�ȇ
�T(熼�j�]Ϝi���
�Ƨ��3�ׯq��z囚C;u��3h�$B.Ŧܽ�����v�q��I�9�T ��^[/�v��_�1�KH�+�Uo)�Wm(8JۤF�K�x>��݌��Yk�'`���q D��=���F���'k;Ot���N�_E��bF˿��d�)�N�����k���LDE�2��=�;�MLr�%K��[n���ڰ������ֈ3�9Ef�����K�'c���0�;�LŔ�Q�JΨ�G�3��nǼn��߫[����Y��[o�&��7�t�Ԭ\���g3*���g�>�����y������<�PqL�>~�g��E�i�Y'�uFk�=>�f����%��tT���f�����ɧ�,��vPxX7G�	���W����㶔��~�{л���k��[�w�W8�4�&��q9A�6m={���w�-�:N�����oC �n:1捾�,�v���:k���	��JPdԆD��Q�`yϯ#q�1�[�:
ȱ���pnش
����ss���^)Q���?A	��?$����B��=�{gO"���}B0�Z�����L���Lk�hgd�zЙ'b���H�TL&���+kz�Utt���-����#��C�?�3[90�`C�e;r��rzO��RO��#�d:�槈���|�.j����8�8Mi�>���ŷ�p"=Ȅ�Bc�l��^�b�i��^��yV6�ų��f���s!��F�٦'�t��>0�s;�����t�v0l/'T,~���8������9_N��x��^�[��zO���-�[��<���s��K���f׵�g0j�sX_ V}�Հ��rk�/Ǽ4j���,��x�����b9��i��p\�J\�J���2t�ԛ�n��bUKM ��W��5�z��X�kM5�i���n�[<������E�����Jn��4,�ZYu!��r��h]:Sx�^U�۴w�4�Wk�%%~����R���vUd�����ġ��U"�iI�k��)8�]=�QY�S��Y��E��c0iXn�ٴ�[�C��O>�v�|&t!�ܗ�Q͵�hZO	�pcYk�=>��އ�x����F�r��Y�]�U4�D����P3�ni�۾辸d�@�P�;)=��'�������g�Z.�?��y��pW��TzŎY��G��y�o�0$}�A���B��.�'Q�-�F&uMm��z�ȧ�_��3kN?;��-=s�:�l�w���l��	=lŶ'9�>��ȇvx�sQ8J����
�t�PJB>�eض�'�y�����E����i���I4����m�tůjf���+���)7�Pj�F@^�?q��a*���)4:����7�ahO��q備�[�NE[it��A=H�V
5��`ۉ1P��n'��,�w�w3�@������q0�]��2m�����e�c�開F�+
����2���5�h�~�U[��+[W�qZ.}��|�~`\k���5*}��)��>Bd^�ħA6򈼝��+C0�V�mO3����6��6u<\,�M�xV퐫�%׉1wEj����Wߒ�ٯ�p�����C4�;���P/k�ռL���D�j�����qd8���0�vnr���P�,��p��[�F��\Vf���b�!�����Ѽ���=�H�[��F(�%��l�	�mр7�56�C)�ۗne~9㞨����X�(Ϳq�rE����Ħ���&������ݼ0��"1�C��B`��=N�O\'�R��1�x��4��JO~F)�u��7xb->Gf���6�8zhA��q��t���N�����Z�ΡJ��aTrW<�7):NX�����̶���|K�g�h���NV.��B��������6��H'�d닰J�­t�)U:�}��76���o�]r���ݛ�h�u.3�匆X@pa7l��Z;MV�V��zW:NK�L��g��=z�*����t��̓ۿs��7�6*9�6'��+r��jR�z�~ٛ-�Ѻ9[u�N�r��{6�ʥ��ǠYz�{�ǃ5p0C�#-�&�wkX�^u;���3v��0C�Iv�e���� �c�)��?D��{��8���˗v
���vFw0�J0��\��oWs�v���y��]�g��W�>���J��jvP�+�B =�ֹ�ٌ�Q�;v�Щ�v?l�oLt��#�'�u9���~�/�����ғ����m���{��hw9�v)c;t|���M�I�e��Ǯ��R���;�:w����W;���Yђ�閣�{���;wb�1���q�{}s��}����"�̅��/�x�g�٧�AX �ǚ-�>uE��X݌l�$<6��%�rDϛn6�3\��/�M��^�����.����LF0�~N&.�ߪ�OV�K[jP��Uj�\���h�ڙ挌��M�.1�W�ce��?�g���1b] F�*,8���J�"��ga˕5W��H�r*i̊�p��&ؑcV8����������-��WzK`�5���'|O%JR�٫4�����d$Fw�j�-���t^n�v{������	.^�ɟq%S�t��u� CY�S�3�K݌�'wr$Hƕ�D��n�{k�I�z��os�ęMy�_��v�H�9Yۏҙ���?�❁j9wa�JХ9���ޢ��`$M���zk��S���v�1Lx���ty����T����Y;�(��l�g����T��s�t�<\M�u-@��oS���fuW�enFrkm�h�G�Xn[8�t��G}C4�]��\����zg;��O'W�i]�tcM[�4y�=����y�	�1M�Y��������q���/h��W˱\ܻ�Vz��*$��M;z.3�R�w07s�����ǚ~(�dp�ns1W��=�#�4���Nr�9]��_oqD�pT��oH�������� 8�g7_���4�]�f�)Y��d��N����N��'�G�Cl{[��s]1]����u3\���w|��K�l��ܑ��g��==���ɽ(��_]G�; �������.��Ɓ)p�x�5��W�tl���f�)�V	H-<�}V������Y�^-Ʃy{��:��+��$G��m����}�=����be�qޯ9���0V�C��קX�8��'T�	����N�[N#���u�DA����gg���4��4�қ�Q��Մa���B���nوN�g/w�/eEPYD��\{���7�]붴�Q0���Ӛ��ǭ�d�2��6!n�kF�V��IT����\���9�Rb�*�.�{K�	��25�>
~G�p�;H�t�	V����f������i�=Vk��9�Z}�c&B�V���{�����ydуq��zP�:"��pP��7�s��h7�E�C���w�:ξwLT2��ZeR�p@�x�m�NH۝��n*2�p�z�C\x4wVT5�.���M��.�7���g˜(vu.\
�8E�?��U��{���e�R�K���
q��q�J�����R79�wJ��}�}���ܵ蔮�$�	=Hs�%�h#df=�Ab�p���i�1�9;a휃}��l���F�{2��ֶۢOd���-���r7���v퓰!V�\�ȹ�j�����Y�3}�"GZJi.�u(�,�F[\3|�0�)}n���K*�qƪ����%9]�p��b���d��3�BQ����Bv����"��&�c��F�@�]A��'�La;C��x�ѫT4<�o�_s���l�b46B��d�<[a;򩥠�j{���u�f:&�M�4s��G6O]�$��t�.������i��FM�㹁��V9H$�zX��g@��𔍊�O����6����O_>������>$QD@�Z
�U�ng�X1 !F?�c����v�^��d�!�[k���L���|�'��`2�4�\�_�T�0kׄ�2g����~{V�p�[�5�4�
��Ž��^���ښέ�!����5���z	����l|]��3���}AK��ﳉuv6�	R�X�^����&�w�����|�Ҫ�T����� Ȃ��ed�T� �a��f��05;�)Г�w�)�aDWr���%e_djU��{�L^E�L�UB�/w:��k����:���*�#b5�
�f�I{�9y�cZ�:��K�\,V�$�<Lz�8.�\�HF��;ާ⨇�O�S�p�*2y�w#-	���x��5O��V��fJ��u䐹�?eTW�h�e�6տ̐���]8u8=��9$�t�(����t�9���软9���>H�x&�ў[wJ�S򟷏��넰.���ҟb,�ˤ�=�/`p޷讉���з�)��ٍ=j;;�DѤ�.����}���F_H��Z[b:���N�Xo�%��F�Tf��s���r�ܡNd�m!M�O����۽����Lh���zr{U�J��X{VO����߷_�<ʒ੗�P��T�*�&(\-۽Ij���,x��΅ПG]�c�ص�[��k�Կ�zy�Ԃ�Lz��]���	܂7A�g
�!͍�LL_q���}4��ɷ��g�����q�6kH�D�x�XsWuv�6�C�e�FE�'}(_=3�E�%w@�6���u�L�3���]9�-N�L\{}x�u�;#s�t�<9:<��A�z�Rf)��j�����{�q�S���y7f�f({1p��gI*|�G���^f��0X��(]���SQ�vEŜ�ިs\L �!��OH���|nV �s�s����b˜��OkZ���&d�9�yO[�	�,�.��g
�d̦�7�k�d��$���5|;'T�n��_}���u�b����o��I���aM�8���\���bS*.��J�S�r���		�b� sZ�(�H%8pt���#���/����ű��>���j�_�H:ߞ�
A"�jų�z�+u����K]�䝚��S�z�pu�������iY\���ȩ�;�V�a�f^����Y9%kP�5�vY���j)���L�F9v�$%vv7��^�yK���W�:U��,=�U��B�"��[�� ӗۯS
!/H�n���V�)�f��V2i�|��c2�T8omo7�t�!i�����
��۔ih�犮E28;7Hs^^N}}�U�w)9����7Yԓvd�Vu��}�����Ð+�Z��5�̝��|��M��5	��;o��r�K��3.0�\F?����ՙ���1ν���ۮl�p�g���}ݖ��Z��MT��r
���4�Qn�]��7;jI8�Cgy�ۺs-,�&�WNQv5������u��}B�ok�nܙ�I��=bK�wp����ۊ5\Y�\0��|��z���u�\��tJZ����9ȃx���A��X���+�0W5}Cp���Z�o�sSxabt�>���ô,˝���V��,�ݤ�E:��ÅW#F^��IޞbG���!���CE�n�xkK[��-�Z)��Dj՝֯�uk����[�9u`Žtj����]b�@1���)Ld��He���;�xԈ3�l��Fe��SRk�0/i�]��2<un]r�n�I��KJ�%Jm�wYT�WMmuՆʺ�YV^d�Ŋ��G;���51&�Ek��e��w;��6-�PhBA=Wٮ�x.f6�bt4!�׸�݆��1�-V*��Z���.�%�,!��I���\Uo�U}*�Kͺ6+*N��������$�ڱ���29a��:�{X��	���mx"T��(��j��+�>�gJ+��.�i�!H�@Fr�^@hPSVi��t�����l3�M��op��v^��P��QU�Ȱ�����F-qp�Bwu̗���w��[5�:�;����Nc��0w��7k�C��^-�D�����?
�+�H�EEW<����y<�Ȩ�y�p܇�N	!��^��j������~���}�QD~�����)��jF^�Q�w|�J+�<��RU���Z�A�M-�Q�Rݾo�����#R},4(���J.IV��P�5Cs�J�sȢ���)������v�������eY:mL
���t]>�竺ou��̧1���w^�<�[�٢G�<�>Tn��g3#�������QI!��u�<��������TU��\�T0��x�<�z/0U��U�fIB���	�����R�+��g)C�r���I$b��B蕒T躁�=ww��DUQQ"��\�+Γ�Qʫ:&B�LBsw{����Gs�Rw\�!�S	%�8��W]ۄ\*���0�̏��E]�8��*����|�qyS�Sq{���8�1V$Q{���Eʢ�fJu�k��U�N�-{�'S%��O>�q/8븙�=t���9�V�oO"�P+.��]=詌 ��s19�/fT��[/�_&�V�͛\�׎u3�}�^1(�����˃a[K�c�������� =[qm��n=V����Cdu7o�s!���S*^��B����������w@���N/��t��4l1�G������aY��F�V�n���� �r&�H9#�v��nyژ `�hr��;�c�l��ѝ=a��q�%�љmw�H�H�%��ח����_����A������	��Up�x�r�l�Wn��0��\zyQ�ܛ�8MV��t����j)㡞�P��w&�c����[xPV�.EO����u��>e��yJE�:�jS���p�X�FE\��)��{k<�ʪi�����6E��@�p���՟\Ϫ&�����nC��g=�]��=M{//��ܥ�;0Ϙ��:;�y%	Kd��78�x�g��H�����&˕i��]�s��>f1�m����Gt���%^['�+����t�B�/�������l�v�8R
��۾�sS.�V:��U!�\�^>�������7�hqc'�U�S�;h�{�W�\s0
�zr���w&���R�7��;���h-�\�2qκ�,K���g����gNPD�A�Ք�:5�v�Y�����Q�5��-ĈO�I:�G�Y}��D:�]�<6�!�L�A�|��!�aO�C��Dj��&�'�kb}�GVwr	�+e����X�\D�\?�]�5����W@`���C'����Ҫ���1T����.��p�^����PV�k���d3�����PՕLԂ��7mW���鸻U�?�QD�W�8d^J}��9�GTft6w�5�����֐�m�X@�NVȎ�3]�vw�?t�Ά��?�εtW;ٛ�� D�0�g v`�M��OS�=îF�oh�!3����+ފ�|��肢�P���%^� vYy�$I �j���u��c�r����2E)�xM�K�"�o���ڙ�锑� g�צ��.I��ܨX�ydI%�VR�6)����dy�x�۽�'{��W��
����}���*[�r�4�Dl��n<{��+�K�K��y�^Xn"�݄@
Uݽ0��5*:�_���E��j�i��.�M�����b��b�Z�HIYۖ�:}�+��WB��S�wdg6\�q��j����2�J��5�Mj�wx�)ogJy�V�9��!�E"�޺)��ړ���	� �&� #my+��F�=���Z\[��h�h�b�.�z,⨸��B�P\�3Ǳ��.i̊>l��&rNVK�y��u�T%�:(Fh���C��m@�&R����2՞���VD��)�~�����*�:����]��b�mH�tJ�C���y���UOs�Ԭ%�.!{����c�A��P�mR79�wJI[�u���	���H����1�ܺɳ>l��m2��-�#�D<��%�ۙOӛ�~��$�9<'Vl�4���c֩��k�v��n�0�ӑ��5Q�ު�3B%�(��[��Dt��鞳�D�����r�| ;�k�3p��kY�L�^�%sp�,+4�z7 �4J�\��rSKt�zJ�R2F�
���̧����.�v��
�@�8�Y��>�4��]Vc_ˬ��3Ϊ_�H3?7.TEU�'
8k��`�� ;:R�7�qZq���U���.s]��`$]qE�p���J�eu^�ƺ����A�x��D�,��Q��Zo�����mPX&v�����lv�93xtl�ӑ�A��`�+�i�K~���t?0fQŮ/���j}
��z||� �?b5퐶{��z�쩺}ƽg���@�bu��4��H�#�2�i9�p�u�IX��T�RجFbȺ�W�]f�8H�D�â�K�y�|���`�y�fX5c�UQ�&f�4�Q�k��w$Dxi�[j�E��^�c)��]c�5Ze�Xd�d��
�xL��{2��Ȏ���H�`�>�]6�#�!��J����6�vUy�����R��7�Q�S�,� �*�GY�5<D-vl�hϲۛ���f��$a�z��?mu����<-Z:#!Q+�y�Xh�_C���x��y�sʏU�駚j�("���6�7���c����g#6:�	��j�l�TQY�M���ߧ� H�I�(].��DS`WF^**��.�w�m�$��T�L���j���a���#fU:yR~���Gr�Oܳn�qd޻��{y�S�Ε-]��S`_d������>��8#�8�z�x�$���v�t8�-6m�����A�s_�U�t�n��M-��T�u|��'���yFI�R۾\J�/�buԏ.���q��n�G)uC�����%Q���k��rU.��Y.�"�'w���[ml�<�3T�b���Y�C�Ô����J�](�Iw/�����KF�E��@fÓ�U����pò�	q�6��9�UܹU����[����ݷ��&-�*&��a�7۾`WO�_�G�M*
4*��[.��۾������zx�oR�����}/�~+�z����|l~�2_rI���W��9�*	�r�FO��{M�7�����f#Nݫ�U��b�q�W>q�H���o=܀�2A �q��`������0�:Xǎ����A���Գ��u~��]c�t{2�7{�F�%��k�7���Xx���j�{:��>R�<p؀F��l�ѽ��ԃ�Qp�l�/c�F��u�3c���\&@R����(:<BP�rb��s+T��,��S��T͆J1�<��^Y���Z���M�+��n�͠���Q�יX�)a2�?s��|X�m���]o���jޡ-���L��m��'uqu���^���2(d���L�0��Y]:���7���΁�4��5�,�I��*�{jw+�L���66YЪ�~��X�Eg,~�PO5A;�"�H3|E]���<��FU)7'j�%͊�@�yd��lvi3ٖ�ФB0��ݛ����Z'qt���'�y"���Q�o`���~��!��
��M˜f���l����N4���9�IU��XIl;�?W;9ɹ똗��j��Ñ���%�܎��Q�Q�_v9-�*ۥ^�ȥ�^	���5øNO4g������,�ղ�I�������pZ1�n�d��������� �j-Ҍǻ[a�t0Y~�U�5���t6:6轓�r���6��'t��4�������{1J{�;����\�l�wd<zo�$��Z���&ԩ�Y��g��r��Wow�%��w��q\�Лss��Xy��w)�/�P��MU��0�B����)Vh��U��t^�I�*�ӷ���Fݏ%��HF:�ba�'K�����{ad��i��=@�R�g+(*���WZ᠕��z1�Er���i_2�EŻ/8�]�!���鯵MS�8V���A��1���LԽ�:�X���3�0P��Ώ��s������?Um_#��f��=��y�L���;ѹ��$�����Y����h�~vp4r��xVkg��7���q"J��UUr�h���/�n2/X�
S��;W�wWC�J��yG���d9���
��	��ݓ{hz���%hH�E�^ҟtS�%��B�C�#QWi�{*C���[a���;�(,�<����i*(�Nm+�W��(�;��rü�Z�KcM[m,�����L�6Ҩ��(+�%V�=ǱW�^H��3�g~9[�͏��+3�X>�f "Ȏ#N��{[>m@��I\��{{�o2�Y��6k{/�t���H�g�� �T"����;`��I��.3'"d��/y��w�5�;�L���N��"���e6���y�L�ګ��L����٤��� ;�6e�5�h!��������n��cJ��ι�Ԃi�V��9�ѽ@�ms���[E�v�b����onk��'ܽ��ԟ�Zv9��k::]�h�9��h���^%��Ν\�	z�.�c�Tw���wLRz$Z)�JP���b��`���]W��+�4�M�T�v�z�E�+�;��֒�2�׼_ Y��Y*{����-P����,��;p=L%;�#;$
�du��i)���.ǂ�e��P��P6�6/�0��u7��hP���Vaٝ5�D����n��(��^����h��בٝ�|)�_0�.���
=z�@+���m Ou=V�P�g�k�*�n�깂$�JCv�7��t?b;n�����ԍ&�V�ⱙ�{��]d�WJW�l򎓴g�1�t6�i���꺮y$���J1�*y�Z�U�����e���#t?'$�g�Lc!��������^���#�<����.:�-���P��8��l��h�-̍�r#^^��,g�����#R+���)w�"nv�,�:��|
�$�+%A��1�1��=Y�ع�T������u�N�Ej*��wZ�S�U-;-pH���������-�!�}6�h;�@�H��.��Z�mΎ����1t���;�x�{g*�G�9��� �]c~�u�o<�e�2'+�J_^��|�X���K}:Miה�#3�/�
EM�rb��Ʋ�q��WrV��!�>����hGI�}(�;�-R�[��+X==!Gq6{��h;��Z��y4b�n!ZSY�c��[etӽ�m��m�;�~}�u���&��S�w��y�e�6!�s����]�-y�|ֳ��I"��I|�#r�H��-��P�{�؟-�&��.�R�7ѻ�nI+Ҥ��6��j�3��Q���$E?<�뻾Y�`H�羹��Z��ax뒨.���ґ���;<�v2��O0Tn՝�2��f��#�u���n�	=��h�T���;a��`���猨u.�u� �}�>�z�%��9�]�x�*��t)971E�߼�dO4��&[*r�R<��4�q���l������4����q��L�U'�z2��/0�{�Z���6GSt��l,��b�/�Yo.(��Rj�M�F���u�	�r�Fo>��6h�c7���s�úMG��S{���iY�r]�z�
TWf��u7���o�w����X�l��C��OD���p$:t�Y}}/ ͡�58c��n��5���[����������uڡ'=搚�J�iY���7�Kk�ک�I�^�I]C���ս���/y��T[���6���y>�es��C�ܓ�{hӉ��V��gtig�W��o�tf[F�p�D�{�F�~�O�$7e�3J��)�M�	Zg@"�f@{J}�WY`n��C����Z9GZ3Zf�������o�O�k��"Wv~�ߕ�����*�K�5���z��zvyV!���+]m7���4�}�΅?�#�8W+�i�t���2������!��3ܒ6���s�u��[:���)��:}�zÍ���9���غCr
A�F��JUAC����,���q���}xz��B���	���m���IX{Ғ�WR�R\�/:0�G]�b�g��~��Ca����__K�0K�h(l����䑔Sds�	�4>��-�x[�+�ǧ�l�0��7��ղ�I�O��#5�a�pG@�<)��y�X�t������J�
�1'�tQ���e���I�mms�qI��\�}�7��hݲ6��)�,��]������Z����3�a�(�r��Z
��>���`���D�1'OH�:��]Y�{�P8"[�J�U�H��6�������A=��3N�aWb����è���I@�W�2#u6�u}-Ⱦ����hbnNMgW2��˝-+C��=�X*L�WG+��d2+f*��u(�����Um�Õ�ɫf�W{�����˴�1��nr]k������= �pv�[�֮�7Iw&���%�2ҋFY�|X?�B���G��z������$���Y�9�K�Z��YaɷL��@LN�؜��R�'`,�	&��\8���WX�I����m6xP�n�&�Н���,�E��Ǽ)���B�F�>2wXw{y�Fs�;y*� ��#�J�'�.��3�6�����.����ouY�Z�}{�]J]�ٙƁ���=�HU��e�>$g>�Գ)��)Y܍G��I�yA�G��i���Ȏ]v ���-�Ȼ�w�r�����/W�}�8��vY[6` �yBL��]u�.4�t��gݕ8m�F���C�VE��#j�����Y~Y^7�Z<_?>��Ɩ06�S�}�}�)S��v� `�zcA���V����Ό��ա�R�
ֱΦ��D��k���G.}�D�A���-��9o�2ۊ�&��S]@���nՍ=�M��ml���\�|����^h��L��P�d$�DU��b*�|:��&3>ʑK���Yd|(�,�J�z�`7):������O��]��[��5;.&�.�=W�\Y���j���=�76>{���:[��]y�R��+fV�4N��v���ܣ��w�[�k�۬�:ҽy]K�lNb����D۝͞n�݉[YsX}Km�{(�R��%�Gw��Y|`����Y϶.!5��r�L楹�YW���{(E��=]���,àD���VVkU;2WR�}F�vp8���]�����ċ�_h�����խU�K����)��c��]��Ҿ}eLFU�W��,}�Mn`PR��+��Þp���ק� �C�áW��IeE+".�U]j��:[R*ޔK��q��,R�%DA�0:{�tK��Ӓ؂�,{ΨX�K<���!�o1�����Q���-��LXqV�m��1K�����j�,%DJ�u������M�.�ޜ��MJB�,���ˡ�����E�c�Ӵ���ku��Z�ɶ]�X3�+�`�&�%����u�˘��f�*}X{YG%�ѽ��K\f�V�umr*�f�o+�S��0"���۝�����D��V�EG��Z�%p�8X5
��,L
���\9���;�d'��[�X���p�S���"4����+�#���1�+��cO>�zv��Q�v_\�/&���}FھVw�����ZEgը�iD�hz=���wO����>�~�������}{=����������t��7�S֚�Ԍ���Ǔ���ȥy�s�\���s��}�}�������� ����	��4���{�T��]-�t�u�*���Vm]����o����o�3��r+�}������%=y9p��9���(��z8�J���ѹ��w���}��E\��I���9E�A�}N�HU�q���Ά��[�G�
�tu(΅�����}�w��(�y�k�9;�V�#�;����wq]�R���uwqtʲ�<j��G5�b{���r*��S��9^��q޼�V�/��0ݻ����<��ws�	��ȹ�z��A�{�=��qʜ5]Y��+"�#���G��zU��Hώ�wwrs��J���s��d��QN�y�Z�o^�pꆽ�"9�!ZTw�;J4=nz;����χI֖�W(�׼]��
��u-���$)�'tr#Γ��ܨq_��M��PQ���r�87Ty/�D��
�7kN�j��<��VѸ����^�R�O+.y��2��k0�j<+)�e`���j)щzx���?����`�gQnF,v��
�C��w*���+sv��MkU�ڌ��7v��0��� �3V��F�?�ހ�����ߋ�k�h�-B�j�]a����P�2::�亊&������to���L�s�-l�֫���dT���6�y>�{pҠ�l����S�����a�.<o�	����Y��\/�I�g&r^~�~�m��am��z�t ��優�d�,ƫqN�gr��[!Pg�g;�`F��ītl{�˘�F��T�׈Q}7ӽ�Q�
�����%_�XM�P�g��rR���,�v�=EVdL��枑s�y�
�W|}���W~B�ȵz���p�P�b8#�b�Uu�~ܖ�7G'�b*LʕAd\�E	�@��4��6l��[��AvL�s��/��kw�t��{���&�\d�$,b\W�\����K���<X�w�^��t>c,%�T��]=�Ϻƌۂ�����65+�E�c�y��<�+��S�V�n��eیw`wm�M�\�;��{�v��d���J��¹އ��N�^���j��3=)S��I���;x��R�i�$ڼ���6���̧+D��5��6�M���U1s�\#V��l��
&�2��VsZ�k���w7O��4\Y���`�;m{^="Q�>�J�ۆ���ԏ=Aܶy�igf�3l���7����J�9�7O�4�.<��@�mB����9y6u=g9��Ͷ�ƃl�<����}����y
zޑ���zsl���피�-����h��p,)r����{%H�n�j��r���EE'0��7[|7{DSHԄF�ʞ�ا�loZJm'�~Q�a�~� �15���"qp�:-����0&�3�lΪ�I�@�ʠ;���b
Ιe�&�T�ĥ���D̰#��F.��#>~���iW������L�.��$Ym�P������;A������#��~����q��^�V;��w��伃�[D�v�`�ͣ���gG3�A�r��?k�����YH�h�����pβ�v�qޥd��:��Q�t��"��Ң]��Ƈ%Yw\qr�C�/A���4�����{2�L�{�������ֵ�xYJue���g,8�Q�"���ِ'v��9&@Ә
��]�q�ΆJΜ���N��D�t�՘�YgG	Ì�X�c���t��eCt�3���3g�4'���d���!�<H)\ĝ�=9�n�p�a������^�Y����I�P�M)Z\:��X�BJ�L�R�b:]���2#g���|�)[���=��P�S�͞�ȩ�\�U��><޽�h��Z�+9��5�֓���R0���Ú��h�.|*�*4��]^j��h^i�Q�5�<��_D�����	�PEȄ��l�D�#l�V���ǥ�6��rH�c	PH�$�]-��2E��]�e�R�u�5�f>�������|�Nɍ�H�g��Ht-�(����ʆ���-7���u3�zrr	k�}kT����u�TJ㬗{mS��C^f��ˍDd�|�ל��v_��.�]�2hJ�]�	1��sc(��vgv�M5z�5���V*������QEX���{V�N5�	����RK{`Gz#���.�Τp���N"NG���Pe�iw%oE��7�����+ظ7n����J�����jv��Xz� 1�Cҭ�ol>��f�����dU�R �q��k�!�oP����9�N"�MF�5vH���&����J@fQ@*ݓ{��r�9�k�t�K��u�j��7{jjxfe�\�ၡ�x�fO;@��W�]=Cz[�٣����b.�M�]#c��r��C�e���R4��zɝ���F��a�a��i4�s�3M�r]�n�h���гN��^&H�P��F�3Q�f�h�o�n&���}�h�E�
�AIa�QȬG��2�7{��D����-���9�#wgWK\�)"���L�B`��&�n��Hw��gs�rz��cUS�%�;���T��e��� ����A({�5�鵭�3�{2e�c���7���=�^b�4��SU�ۚ�쳄*�+q��~�Z����:�V�W���5�tx�-J:����M9�U�xQԯAy�����^/!QV�_���Dxc��7���;e�N�>���w0�9�z�"��)�=�n���yp}ܝ!�D5`���O�.Ǹc��ޙ�3�� ��!Ϋ|q���j����7�H�Ǉ-�X|7oz�[Y�u����Zw��ngv��
�iL��P�i���(R��onwO�S>���G4F�!#�t� ��h�PR�W�j����EȖg�������e�RV>�����$BQ��@|dwJJ��T�ME��}���_;o�*��1q	�3���-�|5�
�ElpX:�@�/ n�$�ÈL�F[פt�Ԛ�oꉹ<1���}���L)�25n�A�h�8YHʛ˾�|��ܾu9y�GRD�j-�Ŏ���
�����pӫ�Y�6m���#b������O-���P%W�4����X.��{4�h��,1L��v���)t�L�t���:�w%�1ΪT��O�/a>��z�{{<���Π�uLknN�Q�9[<��9}*v��sr}!�eIب�2����7^�v�\��o'!6 �>ٜ��p������Y�rX�:��ۇ�i0��Y���9����7��V�k1�Oӥ-ǅh:RZ��p�+�eu�Χy]��7Q�ʙ��n�(L�2�w�̇\ ��떯Z7��t��:,���%r�����ή����&4{��QO��^E8Զ*7� c�Qt,�JP�ώ"�6���ڱ�{9��%d��v]�4f���{���zB@����(�ا��g��!\ܒ98��At��NjH2*����n�H<�1Ű�F�#���<�G���Z}7�-c�2�v#��{����Ξ��1�'�*�*�l\�(MrI��6݌6��e2aٺ��Β�A�wn�OS���N��oME�H�Y@��\{!;(L��v��=X�MζlĽ�A�m@�
�A��O���jP&RV�A�9�µ�hө��n�`��ϵ[��[@2�R!#q�Gb�3j��ɓZe�'�Wf��n:��x�\RT�6:���x[$(?��?S��ތ������Y�e�ǂe$|���ǻ�z̶c��p�Ϝe>Z��{��Y���M��F���/�EMir��Z���Y�ܻn����4�&̮��q,O�[�щ���Gm�#�lO��R�w.Ǜ����̶�m��[0����,����Ү%��1,!��n�\�\��Z�РpqF�Vl��vY�i��y4�ol�K	PZ[Y��<\��s����m�}��e�]f�m3�mT'Rj󷫊�m�YZ�^�D��Dy�w���	}��anߓ�����-��%2�{3��I�FU�p�U���;����F=i	2�`��7����Fz{'pҠ`����Q�0��M�o0�I���;�N~&�l��Ẁm���0๻͐��đlF�t�e������'���%�Q ����ߺG4�YN^�Fʜ��m"�1��50��#%6;�A�2<z8Op�Ic�����CӀh�����`�d�V���=Ar�u���*��=�d<�$�7�j��?��b�W,%���~�o�g>��G
V����̸�B��%R����q��c�f�n�p�����K?�	S�OW�l��ͅ�á��4�w���g���7Fۻ�&�,ȓ\N����p���,Af�6����fZ��91��:s�U��L��&9W��4�4΁�
�8�j��`i�\��݂j:�y`�=�|�84굡��	�q�z�w�GvX3)��ra����Q��G��M�N��*�f��}�u_
�z3��R=C�	�+�	��Ŝ!�h��m+}*]
�LC*��u��!��+��=slZ�������*I�w�������v �Ѩ���%A"��5O��)�̲��dX���=y�[tL��*�'���#o���Q���*J$lj|!�����Άl�b��v?zyx�� B�H�6 �2�v��%R�\u��Ηb����"�W&/9-�Q�>a��t#����X�k�R�G@2�� ��\D5�͂�������2w�O�0}���v#ϫz�
��_)�}���ʬ��չ]�o��]�(*ݓ{�N#q����?�#��yٺ��.Z�L�)9�%V��,�P'�$L�;�#��o�y�)�zl�O%ڻO;b��8�����:���9G�$oFǻM�����2�pZ��1�N{NFy�Ũ��^ײB9�0m�4L� �r}�/+i�U0���0�˷�#��hҷ� �?��<*5�x����h��=�2���P���k�C�~Z�dO�S,H�i&_c�oj�1#ڴݽt�G�Zи�	ĺ���v�5�O����A��m�H���v�,�ʒ��-`[K�ԏ�ds;�Շ9VXD�����y��'�u3�l*�q�SÊ1+b&�S�ĺt1��c'K��.�]�w�Р+�f �1�R�ih �������1Y��vj�H��e�C�1=����W��7����t���ՒP�6����K�Ogf�M'��w���*{J[~PSJ�����V\ә��:�폗Գ�v2�oVm��6��(J�I��PTy#4zM=r�ȩ�+2�QVɗ|��w���^10�a�5fx��D7B��Y��5e4�;�ꜣtok�_6�k��S���<7�Ʉ����6��������Ѽi����߲��'��r������:+jx(�e�]���A���i�c��K��HO��|��V�{gAl,)x!!�,�պ=�X^U��`�)�d7�UحO�lE�Ӌ�k��ߟ���kٹ�E�WK����?W���FS�Kz�S6Iq*r{�F���'@�^����U��.j����G�@:Gx�]�۸輸p��|�`��賬����m����;�Y�
4�w+�4�J���b�W�]=�����}'���z��ΐgg2�5�H&�����w]�G��dں�EM����t�;&��קE_K�"}w0gQ�_9�"����7vvgWD,~n�]�u��S}�J<���2��N�W�w���^p%�#b5�$��Z���ν�,q��[���[v��l���鋹Th��L�K0/��3�H��Gb<�AxO��۝��ӳ�P��oF���GPg�vY�휄�_[�x�'��6�8����O<I	=��� v
:��y�t+�E��M6s=�y�a�6�7Or�okmk��"��>��
�9�VR��G��ߊ��߶�\��V%q���Vn�w�"�v�T��r5$&� IW�8�3i9�hv��vEL��Ý���P�̈�%��Q
�%!\ΞL�ƌ4�͆&����\bB�䋚~�C���熍Z���P)��5�O�DNN��%󰋞�7�&�������[8)����*�[� W��A��Wfc�s��vJa֓�옘�5�9s[ ���̻T�A��jh�DhWm+�M����ߧ���k����C%n��"!�G��m��K���M;:���d�g>�c9��`��']�7�a�6��� Xa�>���F�)PKs���w�S��W�39ڰ:��U�d�Хu�u(�l�i�h�O
�X��	;NI��f\�ZN�\���N�R�=ܾX�W���J�r���6�u��/C���+� ��&7'vs�[٣c�������e�;1}e������:Ď��O.���,S��2����#�_�fJ�[tI�YN��j��T�]`KG�
��>\������k������X5ϕo�Jߞ��B��u�@�sv�Dq����ZWn�1P�����L�7@��:�s��ˍ�;P��C��\�U�hӱh��}���'%���g�^.Y�#uڢ��W|�j�-_D���j˸$����*R�Zd#�W�:��>c�՝٩�&%X2\}�I��8�6X�&��� ���,hrk�����wf�O�W q��P���R����K~��X�r�9���,��
[FfQ�9ǆ��炎����k��W%|�P|w�-��'*�ʯ���Iq}Ko^��6��̍�}�.[,�=�J�s�Q��}�=jv�ZF^~�|��k���\P�ͺf
1J�zR��j��Z�=��,#��guC
ӛl�ZF�gk�4���I�=(�9�{��5��ס�T�q�:�VZ��`��ˉO�V�t�]�z�򗣻��owf�����-����7cD �T��l�}��x.}���B��7f��G�D�'9$���0��A���J���Ë_hW7���oԻ�'�����ޒ�(HykOm5NK��� ؼ6k�&��-�N�v-hӯv�Q,S�S�h��˳��c�\c�IfulΊ��4}db��a#�u�ݎ�Q���ۭ��+�Z�z����J��K�*S�k� �Xo\��)�s���&5J�9w)�JKl���w����;��P�J��*jYh��p�t�m��r9c��!w�K�͗���Z��ʃ����|BκۣD{�������HIW���� ���bW�-8v�G�G��&��h��x��p�aO'ێ�k�mИ����]�R��(���n�k�E�r���W+���f)_H���̨����d�Cu��kӑ�4���� uY�A.�Z���k�d�3ϑx�[t�������qq�����>f������%t	��(��p�a�A&n�V%�E#R��}v�=�\�Ҹq��լ����2Sq	U�GV�9���̪�WF�/��������{i�o:$r�����x5w|�����Ӂ���vI����6m���l�둾k�
:+T@|H�@]����%3����E*���+"-).�>���:��v����}�w�7߷��C���^��:QUr"�*���Y�{��̧z�T�X�ǟzUp�.��w��}�w�~�S^{�E
�R$����:]d��Y}Y�
(�72�A/{��˽��������k�*�I��\�$��w}�=��ݤ^��9㲻��������E��������E��#�c�_Bz�T��N���z.���GtH�k·ͅ_'��{�'�xwIi����w3ժrI
�G8�wI�W�C��H/����9�TDD!6�&�(���\�V�x�(�d^��>��{�!S�m�w�g�I��9��9,w=�p�n:yV�8y�*�n���k��TQH�!��"	���L:}׽x��G��^^����TT��t������5��i8듆>�Ǹ���<�y�l#T�g����I%����=H�R��'��r,�twk�:��x�{���;z��9x��`{R��G��@$=�Q�������j�)c��\G�m�[f�̂����cJ�};�;��m�ɣ��/.�����s��"K�vNn��t�O��O�}�����T
K}o�5.���`�d�T5y�[2_�=0\�����oOཋ-�$,/�RVܸ�m�Ǘq6d6c횎Ĝe���UD����91�cn;l��T�4�_��l�vJw�[cZ�D]��������Ѫ���OPn�kcGZJi.���3cn.mi�xlO�R����m��\_cS�9���՞<�<�yn�gV	��#K��ʜ�6���F�
���0f����}�Ԣ��n�jMN��|�X��v���푛!�=�}�t����I�ۺͪ�U����&�7� �=@�ʢA�c����oá��2��d�.oy�OXc�zܣ+���:<r̀z8H�x�����u1��/*^ȸ����5��׌`(��<wHثF�Ne���H�W�*{�|&G� ?Z�M����e�2覐���4kUm; _R�j��|/�C/y~9dvomph+��PÃ{v�1ۜ:R����g���F���m��gۗS+��R\��b�ܮ�\2��\��RiK7�Ck>��O6,�Ã��c��Iφ/����}���`=�4&j�3}z1W��n��iki2�s_Sc��²6�[��g���MU~����ȭ�ni�]G[�]���;Շ7A6��:���Op�
��`83&.�O-}ӊ�&﷥�ݔ�d��ۤўU@��D�][ {,ha(m
�-$W>jz��ӭ"O��A� m��ԑ�K�0MW�)w��Cz��zĶ'���z�z�R�
pg�C���n�<�@ݔ��+��7J��Q;~�/S�y(��lڿB��,e)xД:�F�a}�q���V�k �1����n:24�ֱ]�^4����A�>~�GY��ؕn99��Q���������uJ���{��:�L%���5��d?-�+�"�D��+q����+M�eoF�r�
�g��:X8�`�f��pp+��Kµz��!Ƽ3y8�p]A49*ĠE�bȌҳ[Ka�Ƚ��(�}��s�ܨA����اU�}r�U��Kc^�}�
��V����WΧ=\3]�ڤ�4o(hq}.������%X)�p�F�m�"�'��V��b[�97u�")��.�%��Z*�˱���,@�)EW��F��Cj{���H=�h��V���Ʀ�i'a�Fg���W��M�̅Pv�{n����<���+ǣ$oF��7w��ڞ/n=R�%n�!|H���Y���|��	p�6���mtj]��h������S�-uH��V띨���f£@d�#c�tf[bf�|��N��Et�G-�L#h���϶
�k������Y��RU隺�]��ȧ悋&-oUm0M�7MY���VI�U!+����R:)�a�w �%L�L�{V��Tц볨��I0d�T�<���p��U����yJni��u)��J�ծ�3nXex�=XL�c)���%��uܒ�hʠ�ܝ����5sZ=O#��7;0z�]/�p냓l����غ|܂�Ѝz���ۋ�F��k��f�����[g�N��\���[�ǽ�*�����ѷu�#���O1{�j߻�v�����Ŝ/�J�l���m�i3˛z�Q�����-�es::�3܏4|��:*k&K�'��o:�w�����n��:�*.��Y��ɹ!�L�FT�@���>�� Δz�7�(&���ӣ:���}Q��~��{��zst�u�P�<{��_e4Qݞ}ZĿ�wLNs��WƑV�H��>-����L��<5�s�~�=�yOy[к�ٝ�,/6�'��uZD��[������"���^�~���V��#������l�h;T	F$+��wd\e�꽴���@7�-���;a��q��^ӊ�s2�tu��r]EQJ�l����ƻ�w�ûݐ��&e ��s�� q����nu*r�������%!`�J����(?v��CY]�ru��Al��$n��E��.�y5�d�B��-jgĎ���l���U�x��wh]o
��6��S�kkp���}[����Z6<r�o?q#A ���;�ا��A�K#Kk�D��cMۛY��u|i	ayJ�^�y�M�;O"�yJ,yo.Q��	h_�wl ��q��TK�)]{���W�K*!�V�Vڴ���L#u�Aʚ��e)��jD�U�|��R���)��K*���m�6��R�/DU	�Ï�n��F-�4�-�I�i
��ጞ��)<N/�|��x���.g��-=�ј�s�+��zED�U�^���ǭI\��� ��>��
<�;K6N���Ys5�p���̵����q�����q��D,%%��!��&V�b8��3e]��G�$\ө � �nx_��S絰��a���1љ��vI�����U⌥3�j�S��g�]9 B(a�h��-#P���1=ټٜeD@h�<��I����w�J����N�iq �A؍���Ѭd�Mz��E���./;)���.6��N�(�	Z��q2���=ɞ�++�
F����)i��l�4M._�E���Sr��[�u���姶Nv�~�1L/�m#y�m����3#�'��VaY7Ҭ�t�����r�ד�q���l0\ˋ�j��X5�������:�0���w4I͞��΂$�5#6Xg��f�#zg���S3pg�驺��z'e3����7��,y��)���κ�DU�^G��7gđK4�n�����.���L�Ys�q�aK����%m
[L_.]�gWQhQ}�d�N���\��a�j��)���hvR*���H�Ǉr��x���M�(�iU�W;���/dg�*O�I�3��2��n�t?���p����'v���=9z4�y�r#�V-�G��U�H;<c�{g�J�*h���
<�H�s7�T�!��F��F�$w9d����8��^�%����.q_��dL3�P}!��HثF�����Np��姬�}M�K{����1*��~�{;B�ߧE���	���˴�����}Ot���E�_B�ʁ���N�
�:��t���T�S��<�R�(�f�����;ר��33r�d�&Ԛ�GZAꊉs8Y�����k=�NM����U�^>*�]<�+�Q�&Mx�*�ם�4�se�j"	��bi��v�]��ƅ>����nǨ>��K�*|`�l������ƬP/����5��T��D�r��� m��w��%mҟ�X�����r��ɰY�Q��X滬�`�}Q,�yz^W��I`��KZ�t㖻�N���!�vs��\�,���}��;�F�k�l���v�R<��"(�\��1���h$�_e]�=FB�C��)s�s�����s��q�,b����{���]CNr����X韁T(�a�V����������tp�t�A��6+L����%Oq��X��)~6��[1���f��8Kl�����L�n�B�a�����6�]��{�w+�!}�F���;δ(`����6����{��e�m�-��j�Od��eW�q�V��)Ѭ4��K�`�e{N�&��l���m����	w��C	�+U�J����f��J�����u7I�֭h���T��6i��ӧ<\&ѝN7a���:���;_�'��?	��ƶ�}�/�}��p��(@��Q��Ώz��T6BS�޿>��'OA��ph�H��AG.;n3O�"=�(Ϋs�ԁ}Y��M�7�9T���̝�*��9�'�*o_�}[^(���tTk��|ψ��\=$����DtC�5CHʣg���%�٘�|ǧ��(SgN�觍�z�6?;V*�խW�'xZX���qʏ07�V��2p	�m�c��0�.ק�=��	�^��LG�E��By
h�}��߱��{<�U V:7X�u<�z��Y� ���Ä:���{�ea|*��6�X�����ӛ��ͼ��5S�6�&�K�]w�--o��[������5�s��&��JVx��/)M�9���B��I�����L�@���^�Ī2 v���$mJV*�37��k*���N���V�V��}�lH�XD����v�
OB7��ݢ-�������n��5@�^P�k��|��)XɄ�u��Ž=᥯~����з�Q|O�y<}7��%P~���N�Y��[S�&�SS=K1Ok��������;��h�*��M����[a� �@z���y�S�^�9׎M[���'���ޣ��H�E�#����5Ul-�Byk{��B�Ws�������ӓ�9.�Yf'���6�},����V��evu_��Jg�	C��oN��腞f���(���O��kpm���g�������g�nK�c����k�
�ɳ���Ʉ_�3���]��j����vސ���)Ɣx6Z�R�Xq�Ͳ��R�A�ȫ�a͊ծn����@]od�AEWPN��%'��SA�`��/7�pk���S�H��;Ҏ�{y���,��S௴#'�������{�+�i��bH���v��������k+��Nj���Bx���$,����w���ܧ�-�^��c�xGl}�:��Ѳ=�+��A������{��5�.�v��X��Ϝ���ѻ��O}�	G�����X���~_�t�H��ǿ�w�v*?�WEd����2�yĚZ9�++��w1`����1�P���D}]On�L�ü�S���8dF��T�G)=�|;��&���f9�oQ;9�X��e]Y"�=�/A]�w�w3�VME�j!_o����%���T����?��ڣ;��M����*��0xF�Ut���n+��q��u5gAv1q��#*����s��U��= ��Q/�|�.�Ǯ��]���j�@X�iG[��T�%T�B,2�4��lK�O3ԝ�V���!�C`ܖG/��t���ˍ6ɞ<��6W�z�����������P׷��z��1v%��X��5%AX����*��Y&'��C)���Y�W�K��c�f[��j���n�����RFN�P�H��V�k�,��Jn����òi5f�/�F��%�^�GtNX�4p�mս��<�O?lAێ����xd��ir���w��3wD�DT�m񇜆�(ʔ��0�-�L�"!h�������v{9�4N�H?�ǻ�h��gR�v>�2��!���s��I�"��a-Om""���T�b9]�o����TzP����1�F�8(��)d�i��o6�U�f���o�h�]^/�h{�ƿ�^�m��������*�;6;�����6�Xz�J�7mv����P�J�d��;FG��e������U0NvcY��emr�Vuw���T���|0Kuy��h?/�[�Z�v�S��(
k�iB�����Z�h��9�C�q#`5է��:$S���Ɏ��oW�>�r����m�>^����H>�ϨV�ݥS5uY�|4�Ȇ/A��\�Oa�ـ�|#��ܙ�ndCP΅�4��r��{�Ӥ���~�?TK�����UA}q�V� d����!C ���������@R1T 0AB 1T��q���62�!�m����b� ���}���dL��F 3��d3�0 A�@�h2 A�  ���b e3� ����s� r�v�  p.C 	��`� �`2���	�˓`ˑ3� ;����s��.G;�dr�r�˝� s�˗!�e�8�	�;c ���`.L��`ˑː0cY��c 9Ô�0 �8��93��g�� �`� d � ����r� !�`� � � �`������3�����(�Z��
�V��C�0��|)@��~}A@#@@"jq�C��1��u�w�r"��'�O�<���~~_�ֈ����c�8��1狌�y�N��=;��zl��`�U��{P@���"����EQX��!�\9��A]���������i��C�"*��OwW�ݻ���
�:归N!L�g�����j�����ho�;�iBvӉD^�Q�� ��}H� �   �� 
  . � � M���ɀm�A0 E��H*� D`�0 !� � l�n�Z � +  �l�& �` L� ����� &�l�� #� )�p & ��2;  ��aL �6�lc1QP���(J�$�*���R�  �H��c�8���_�
@��r<�]Zh*��x|��\�QEj%���-�5׆�t2��	�)�3���цO�a���9:��+��;� ����{��oz�2�M��@UE`��+ԇ1�Qf!��b�(��!��p��jiQX�o/jU9���� e`�� ��гζ:cX�l�`�(�@�DU�����N�>��������A�d8�����/i�v�S�@n�������u����5����}����(���=pC��Ӓ��+���1�3ʇ�D1A�s�
4���m�tT<���-Rb�1Ĩف�p��3�*"��\�30��qԀ�:�a��������o`p��^�̼@QA^�����`�b�(�
��������
[���
!�� ���PVI��aJ�!�"@` ���������x        @      @   (  @ 
   (�     �fѳ)-�Z&k6�f�ڭ��S6�Tʲ�lU4��6�^��5���۶��ٲ�Eh4��W%��X����VVړR���U��m��ki�:�+&IZ��e5KVV��5c2���6(�Me��e���j͵-l��MI���c-��[(I[j���ͪ6��f�M�ٳVe����t��M���R�   ������J]�X:A�:�#A�N[Z5J�mt��ښ�6�i�Ɣֻv]B��iл��U�R��
���4����[ci�B���ckJ�+b�>  �8}
#�f�(P�|8t��m��6��Q�_{��c�
2(V��}�x�B�@��|�N�R�20=����(�Vwn�+N�I��ui[eP�s�����-v�hi�i�N�i��j�6�ܵ�RV�   Z�=�b�f��.�j_m
]z7i��TՃU5��֮`�Uv�M&����ӫ�^]\U-�Z[gs\4[
�[r���U����/:�J�G.٭��	Vf�h�6m��|   �������t�Y��q�amV�r�ų@mݣ��:)T)K�隡M��]ͮ
(�V��5�-�j�-��f�Z5�]�[cb���[)m��3ZYm��  �j"�ymX�}�
v�r�UP.G���Z���kb������@����ёU�:0u�U˽��PR�Z�f�)cV��+f��u���  <�bZ��V��\Z
۵c�7��]�eUT�=��	n�]/sE�+oNz��MA@���uj��[�l��2�ӻf6�	�%Ti�   1�u��{�pP4j㺪�*�Z�R��ٹ��QY��몠�[\�S5��zW�(PH�sǇTU*�w���u��%wy�Vf6Ȓ�m���k`�|   L��)P�a;��PR�T{ގyI��t�*�)��(��yNzѨ�U��s�@�w��z�U%!�z�(zR�Uw�oz�!����Si�M��lT��T�  �}J�/{�o{l�T����RB�y�6�ԩR�^����{���UI�h��ުR@�;����K���zT�l��z�6���"�{3J�,��i�)�խ+�  ۾T4���QG�y�)R�LrzjT���u�1(��N�R�	;�wWc6�{�/y@�%N����J��4�J����*��h�)�)IT� ��F�O�Ĕ�b0 �b)�A�J��#@M�R��@h�0I��L*�  ���������&�F�����{��1]y
��0؂*m��󳂵�v�Y����}�W���?^���}����1��clm����m�cm��m�cm���`����6����?��������V�&��Тt^�����)���=�{{6����f�;�G��W[�u�.&��b�Jv�9r�=.������8Lo�=��l{iCs�q�a�:�0tp��6�R�;ږ�.�`{�&����pY55�U�.Y��Z@ޝ	�.�d�
���c��p��HU�*�V�"n�y-��f��F��U�pm��̣Nsm�NLC�M�.�ˢ�;m+���J0���c]�S�c��}���1X{i��q8��W
<�[�\����r�5L�̽��q�dR�/��p<�wˋ\ҽ�,��=�;�8i;��ai���Bl�����0��ՍN��ػ����w��vo�`�R�7����R��1@X1��*�������pbO[��Z��Y�[;�Q���ۡg��9E�t]>��ǽ ��QG�ނ�]B���s.H)��7p8p�:%M�:C,�roՃ��0�؞5`��>S�}�s��9��.+�%WZ��'>Ԥ��\I�ҭ�yE�����E���\���z)����ɑ�Y��wv]Nk
&�f̌|����I���F�Ty�R4-l��	3C��CP!oRQ�^"�/ ����k%D�Y�.���h'�m�l�	�8n�i㧒Q$V+gܭ�>no`<���J7��78������b	u�p�9sx�� 8��-���׈�݆���ǋ�={���d��z��S5�騅��9d�tj�{5v��"d��uN���}	xr���U���f;;�i;1C`�LL\�YiY::��@F/�!J0�	���j�x�;(�I9�彐U��Kl�8Hct��/�s��'�/n���xQ��:S:.��ڮj�M��,
LM< �b�л�w6p���zͮ
�x4'����-��mƝ·��v)Z2E�\�ћ��#�AS�$�7v卜6^&��Ļ�.+��#���bOZ�#ѫc��sJm���F�fN��'_�OF�����BS;�<u����o���6h��q�h��C�t�齘��RK�8Jvf)��i��`ܱv�+�R�i�J���&݀�x*(�&��5=�c��6Ey�F%υ�4�I���s.,\�<�_^$Ûp�Y8��t�.hZEK���?\���y#��&�0��Ÿ6U)���D"���|CJd�C�ۍ�݆|����b4k��g3	����_��!��'����D<�#\���r�iɗ)��6nJ��i��$��sx���K��dZ�@����k�hŧ�=���nA�{�n1�*.�k� ��Y^���zzٳM�_fsؐ�L�y�㑜�-�\�]Z�ogj̷]�۴w;;ܝݱ���@ZwL���������Rݛv���8ah�2�;��][�O�ȸrp4[��.�����
�,�r�z����B�⹔;!B�� ]N��c7��:���;�Y�kdR�:v}z;�^�uQ�3�|x^�;n�1+h�U�u�s�����vf�f��v��ӳd�P4�(lB;��՝ي�K�>Cp�u�RY�z�s��5��1Q����6w��{�m��s%l�;U/���ovc���"&w�9�ŞJ�dl�@:�,�,�s��"C���p�$�5E�[�]�o(��h}��O+m�CX�aCJyS9�V��J<Z��B��G��嗞0��tpyٰwe(�sxs�k{�	�H{�Q'Y�h�p��OA'\����؈���;�F�������1bgjݟ,1v+��s�q:5g|��&�"�{�Kj��ӂ1���iژ�;9���'t�f��s:��S���`����׼r�2�xy��ڞ
�DHzt�xb�\|�!����m+�w6�J7V�u����vQw��^����j�+s�̌P�mxS=�;f�w����'��Ԃ���T &��̂��~YϪ�p��o��mn؃';�;��&���f��i�Z]z
v�'�{�Uɲ��^d$�7&���\��K\+f��˽���G�,��{y����2#�A<�[�w����՛n�#f�7M1��Ǚy�����H%�F�b�jwL�Jܴ|�E�0��y�5i͸A4I�����;P�d���TC{���s��P!JW�;�
f����;M=�闬Z��xp��en�-a@n��;d1#�mZsx
��4������L�XJ�(Y�S����������5j���Y�yrq��G>¯[�D�9X��0�'q�������zoG�ם���@5)/p���G9�f�fhYo2���.]3K�E+Fk�k6;�Ժ��ע�u2֥p2o
��Fo3[�tP{9Sz>��>�0�dSyuC���Pq-Sx���V�с-���\�I�;�-�E�����0�E��p}���z�c��t��	e�1�Z��tt.�C�V����SZ{'u�o2}z�����s�+FZ!�W��m#�Ӈ�w�'l՜�4�M˔�u���bw�d��:����`(k�z�a�.�k˕̽J�L8��;̮���ol�)6�D������^�	%��}{�H��:5��0�U�{�]̍W!�-^��{�ܗ�,�x���ǵM�ξl�u��q���eMe���A�����լ��㢱d{�=����3@R[�{vwn�P�ԈDq���gAK�+cёf��L, �����)v%����[v�����-p���S����?w�t��#�>���X����b�����-�ña{݉f��ݹd�ƺ�}�%��A����#�ҏh�7'Z�Q��iפ.	���a��1Y0�{��ӣ�M	���� �Ǹ�֨]�$�i.#�)�'�9������%�0��?t��K�VH�#@Sh�mg��&j��p�t3�; ͯ����t=2��`�g]��k�^����dX��zG��w�>��
� �@��.;�JgMm�Y���	��D��]&w:��Y;��,c4h����RT۴��5��{z@�1WC�:;I]�w������]� z��D���*�vݗ�㣤���,�gs.!��0ہn���x�-��T
�	�e�Y�{�~��:-6��}ۺ�<���!��(�ۣ��6rޘ+�ۏ*:IW ��<s{r'ns�l��,��-�l�
�1��C�u��a�H[$��.�P�-j��;�P��GK�4������0�|���B�"l^ĸci�a�l�cl"^ѕu�N��^8�i��r���͚�nr̼:��a4=�NY��M��n�ѝ�<�5I��D�w��/2�֕1D����;y)M[c��<��ٻ�S��F��:�ЯQ��<c���j[[ķ/tqLp艠�cJ�n��an����!yܳ�M�e=󧔵.F���Q��ˌ��yh7����j;6�YrB����ti�'w��m{���v�@��qIk*"QmuG�4�E���d�W�R�ږ�{h�EEg.�;x);6�f��[��%n�泞�\'�*Ǝ��zpS
ewC�V���D���������)�&��ݒ�unU�;T[�{��:��Ź°����i�w�YعU��-�T���,q#��"�QcStFW8{��Bw:��*Ύ	�@3���]�'�{n��-ej�6�(��\y%�fᙧ7M�G�$���j!u�l�|5�a#/K3�tUdN)�ɲ3�SX7R���b9��Bu.X���'V�n�����EaB��'Js��m��**������O{�G����`o|�[v�(�N{ �E1�����M]`�WAQh�/ Ky:S��4��pNҴp�6�1�h׌.pE�����W,F�3H�-q��gV�tV;:nZwr�ey��5W���9E�'W,�&�{[v\�u��2�ٗA�X����>�;��B�2�³�7��`iq��tш�!��`X�[�cw��̝GQ�\B���T��#J�����;B)<�"Ör���I1�j��[��3D|�Utp������7��}yn�~�Fף���gqH�Ʈ�����y=����{}q��Ń+W�wd�Ik��(���J�%����Yݱӵ,=�Hj�'� X��4b}Y���7;`�����=k)}���ܪ�X�u3��,���6�R9�Hp�X&�R� t��A't��؋s"�i�Ar�X��Y��8#���=��dt{)<�K�����$������u��|���NJ�kE��ɑ�2�7&U�q}�lᏏbTň�!��Z�7�E�t��Zp(���C��i��M��"O�E�ĳ�v3y���.���%tV���-�nc��M��L�n\ۇ�i�OBr��r]�M�oK�J{U:�n�I�F��7t�L, ��̶�Q�<Γ��d��n��Z����y�G>�~��d��ե�-ٚsn������Z�I�oj���1C;��[Z�q�.�[��9�x���}z>WQ	���<S�o.�ω)���؀�'�*����]��{�Z0�����4púw �YN/S�����GI���xv��wN�f�-Xɒk��blQ�,�s�Lh�t��d',b�f#�Ń҅���S��-�{TYk���PU� gK�)�뷔\A�F�݂n���׺���.�Xv섕q��;+�mfv��l�Qnh��٣$�X�׷��a+�Ŏ�r�s���k�/�QN{�"��	��
l�6�~c2W��wy�w���v���Ƿ���6Tg`��	��	���.Ī?�{��'my�\|1��!�ovL�
L��/WvV����dVEЌ1 ��fq; 'y�흑M0g5��;�Qh��~�p+/^׸
�^�������{7�"���+7o�%7{Ӌs�f�(�4��Κù���d�5��r���^�۵�����Ll��1��6�H��;/a/�$1�[����o]f��ޢ4M8�|�Yy�6����J�sK�x1�D��\{�p*�V��sý��K^Psq���p8�v�_!F��U��!�E��x�פ����I��t��L��m���nt$՚���{�$�+�-F�UZJ�[��CtD2a�3��u>�u�,Tt�w!���Ho����;�=����jW{��x���z��R�Et�1�fvЮ�DQ�F�C�4cu�1N\O&ڦ �d,#�Sd ��ޅ�n�����F����Z�k#�ݍ^�4	�N�-�V��.gN�"� 5���e��v$�y
2�+'nNJ�۷�y���j�;N�w���6=ɣD7����M�����r�Ԕv5� �Fü��e�7V���c�[�I1���֛vq���aɀߣ���Vc���ZQ15@Un\srq'��	��r=o*��g��5���g̭o5�_i���6���:�9�s������s~�G�s��@Y�	c ���P7:d�1���Vṣ����w�1�@�m�%6�з�a
3��Ӝ��><�uжMA��w-��`�J�o�v�'�)`t��n��^�gu[�t��!�V���_Lj��ò��8R�wwu��4�"6Nr�s[�I�J-�0��5��j�X�8��;��R��PU-P��� �u�0��89h�ꡜ���O�WvY���^�g>�����i%��oe�i�B 9Ĝ]�.���um��3Fٺ'M�6�oC��z}��f²����K�ձ��]��"�����^)(�>WF����v�Y�0�C�5�O*��y0����B�}tiY��d�`ލκB��h`+������պ�� ,{���N�7�k�)MJ1�p���N� Do^����A�H��T�%����[��gx�$Y+����h���)?�=@f�4����p'��	��t�S0������L��do���0_�����g2�`Uj�n7{��U��K=��ۣX�Ÿ������d�<�p��`���6�9{C����o-A������j��g	+��q�^͟���s�ntq;�`����}Y�5�E�砥ˈ@�C�h�k�4Վ�I���ũv�|ow+-�������ӕ�I�b��X�'ۭ���Ѿ=~�=2n9�;��S�=�� ��:O�xs��כ��co�0뎣#T�3�i:�kw��I�<��ܝ`3�WѴ}z�4u]�C��):�=�f!ľ�AN:��LK!����yk �\yҬ��MKK `)s5�r������x uch!�|sN���� ���y������n�I���x��\k� ��RvZ	�nd{7�n�Ao���{��>\��e����3uw+w��Y�y�8�]�Kg���]:�.��o.h��⨍<˯�G��;EǺ��b�h�9۹�p�7��oga�	?*x�v���t�+DL��_57/<Ռ�U#��P�s��Q�o=�\������W�'���Ơ��Z�O�s�w��|�j�4��#a;�u�mA�Gi߲��`�وa`�Y�Y�pۗ�1��8P�h�Ќ]�X�Q�t<�T�r�>�a}���,'f���H��)�QN��܅��d�ڤ����u�	�%�4�F-��.OJU�m��7"P���΀��Y�c�#�BX�W�q-$��,���1�뭈<���K�Z��V��ݵl��\�W�,"��T�L��9�ZG�H�yk�����}/������q��l�t8�0�=t^ �u��/iç�F�"����N��#���˂����4މB	7�9L�p�Ô��-���Z�rGfYm���d��]��`o#�ܩ:�dԆ��y��J�����烰��:(:f\>k^���ђ�{���h��ǌ��ԕ>��.��[*���/M*]f�ق����>�޸�0���[��nq��-��X�<�oHvG�[w�I�C��[�a�Lhɕu ��H���M�1TIGF�P��&��I�]"fn!���!�/e���!j�[�傥Y�r!1�,"�[�o�R�� p:S���uk�.���;u��-.c�z+7�*݃+������@�tlp��pn<����q�$��]�+�P��#r��\���w.YY��I�ks���m�
��Bi�G�y�k�5sQC��s�{Pl�,sr��ݕ�P��ŐI˻8��(�!���Lt(vfWK����W�VB�7=Y��ޯ[vy�{����k�p�:f�hƫ9�da�gX���i����4��)ŮƗբcI��=	n�'��1,���n�9��Nh���ѭf�Xos�����n�����y��;��ҳ�D���(�F�g=�YG�t�3��ғ�r��wE���]�J��+�Õu�����Ϥ�Pc����{��ǵ�m\<��	7o����<+���Mٗ��K7�Xx�ɗ�P:z�G�M[����f2;m�W`雛Ӛ}�=+Ȓۘwg<�\���!�ó��$�MI�I���r������q��|5�^rW�&r�����b��2��J��J�C����J��e�$}m����'7�CƜ��G+O!>Zd�݄������9��˕���T�ݦ��g�wa]˥@�Y�1}�,�N�\�2k����t9x�EB�M��Z���%�gk9bt�K�������o�S��a����V�4�Y�H�����JV�&�S��2S�#r�Qn9MV��eY.�g�ԟ��w�Vϩ�{/�I͙b~�u���q�`�=�;6p��捥�����R�P�qf�i���(�^�X��$����1{8h9aѸ��g��G\P��¼�'F���Wx+�T�@��۞��h;�{^�.'��⋫�!:��kX�멙�=�,��w�RP���`8;n\`��|j��}ȇY�GT�SE��3S���*几�s
�b�I͓b��܍pD����K1A ��b�Ky�t����$v���ѨiՎ+hL�V��e��}F�Twj�����թ�=��^�Ǘ�7��,}��#pV�	��%�]���A�=�[泰1�g>u�e=��a�豚Eg:�JD5ވ|���=~��Z��v�ݪxyrH�y�i2[:O!���)�a����}��#$�3���(.3�y�uL� �.�����x��`�xќ�3�,(��v�2-��=`4p܅�1ml�X@Q���q�]�X.�U1�	_zxdwb���p�3� ��e��܇�W�������^��{�j�E�b�oA�-�ed����2d�!4�,��Tmc��+�7*�����
�7��&DK�K�=t���y������^��Xq��Vl9"���/"�&G�e9ΣXה���Dܒzʙ[��,�e�1�V6��N���3ݚ����f�pv\m�+#^4��c�j�;�#�qӾ_b�H7��X<�2<+��wyd Aē�wLq�b��h�5�@YÊ���X;~�,]	���&Pp��)�u�����`VՊ�n���n��Cv��%�p�<3�/o��!��{�{SˌmݗW+5�;��w����i�f��V_K�0��G�Ur��眤�I%I��$e"�pǂub�C�=�TF3z�xsI�* 5X\:tW�w�-ܒ�ܬ)=��|����a�c��Y�b�*��Z�ato�i����2�t���n!�vX��n�H:^'w@�O)%��8I$�x\��G�u�d�H���K���n������(%���<|l�77k�����B$x_7v�^�0��$���E���sY}���b����� eq]k�3j)F��󭧖�1��ՋX����n�f�(p�X�����<�ng+�t�3�WAgi���K9Ϻ�)keo:\����y���v�z��)LŤ��Ix	:�fW�n��}5�j-��tN�4^9 �2���ڼu}�H�_b�����^,����z�ȷ�"-z=�\1h�ʁ��|�[ep?u�%��Hk��fJC�k)օ���v|�X�>]L5����o��Y���o����ˑ�^H��}*�M���|3���{���I��o%�6M��z��������l�o(�݅-�9��L�z�&5G5W�VbP�1�������;�~
��M��E����Y������Ao��+���̂i�/��x���1m:���-�Е*T��I��Nb�,��}�^î1ϐn�#�F��{�{R�_1���w;Տ[暜���}���;Z�~c�k�Ml��jp`U��(��*�쨔#K��wt	�`�uND�&f�;[x�Rئ��YG�����y{{�0T~�"Y��6�vy���d�k��VLջR���oA����ɨ�^�yxp|��/j�/�����6��=��F�e:j��J*Bn�ނ#ɽp��v?�������QQ=|��fE���P���n�[&-uz�jNY�Z�	a�Rj�;�4K]N�ĸ6ss��e��ڐ;��-P�c�Z3�u%�9ls�:�k��W��]D��L��؞�x�F�<E�X�=���F�i�����`����+o�s�.`���VwU��� �S�H�,����|�R�x�(J��r�;�"��|�;��v�c��TY�O�G��Ӣ92�NM����
��+�GAԭns�m�k/XSn�j����M��eqۻf�c�Qƹ��y�]oh�4��y�(���\�dk�S�lė�&��i��}�!�#�	��8ꙻϊ�}��_:�o�x�7h<'�Վz�rw��U��U�0�����$�DLY�^��s<�J�q@y��bb�u����<��mk��������*^��)�)�Mڣ4k�6�g�X��8�|FWU�]3؞˯X~=!c�`4��ݑ��u�m�՘D�H$�^l��Y��|(ɮV�c���.��{y��_qL�\�r[�S9/C�8���J0mk����=s�數ob�XR���!N�����@῵�tvh�����릧�1F�n��j��&-�1ڍ���;�n-${-�{u��z�p[o�
۬�#B፜ψ����2s���5��+��"�0�l�MQ�I�3�F�^_Wz�N?�8󪥸@�mt�����`�+����P-�EJϟ`����v�=�Fs΋K�u͛'����״�n��k>5�+3��8+�ZjoJfW
�$�lĆ���`�Q[����t��J���[�Q�wO^\~���=0���!�d�is;�Խ��&�c�u��c�8o�"t�/"ig4�Щ��8y�`��;I�՚f�weZu��˵�\ºu#i�nk�]5�E�Wѹ��5��oQ�{�^s�qx��� �o\}L�4�y yF4�T%J����������s*��'��n�{9�i��,��p�)�k���z��p�'�W��t��睴ɶ6�9g�!\ށ� ^�r��@=���e�T�x�=��z�ڠ��]'h�TaT���^�jM!���ɫ{S�]��o��Q�m�-^�ݛ�f�C�mC�� xp3�at�:r�2	G����\{vK���01LI�gN��,ޥJ ��Y�4�RS����^6��R��"+h����lPʑX�s"�v��@�@;i}��^���WgnΒ5i4� ���)n�}��lk�͔w\�{̧��i|� ++O�'���Fj}텢6��Iz�R�9RQ'w-e�#��G!��V�b�ѓZ��|e޻�d�H��Ț��?j3e
�%��>����oF���'�uߔՑS&=����v�!*����nQ����ثC�טQ%>�y�Et]w*���Ba:�q*n��v�)�e�S�P��(΄B�6AU��J��6I��V��[)\"��[]+�x�7�kx^]L!�B��=7NT���ah�;+e���:�C!��xs�2�����>oI�{4<�^K7`=�M�����+����a�,Z�������iS��1�B]r.�i�,�3&���id��H�ч�s�x��?g6{�=�mN�Eæ��X�C�3�,�"&�l((�*�n۪��ﳜn��oc���ge,׵̧���k��$�H��L%�k��hw���ꥷ]�b��=眐a�3�v�pN
q����U7g���/=�un����_n�|D���W�8�!����ʒ�^�06��E^��#�˾=���Om�Mв^ޏ�kl٣�]i��b��Ы���M���	gEt��AL/�HӬ�n�k:.	���1�6���7LLͰ7�hѾ;�$��J�5��|F{��f���%p��B
�{㙫(���5��X���X�E�;�7�;����bk��wG��O%�Y��..,[j�Y�Ιc�j� �A���ss@"y�IxќV��:�ޫH���MI�G`�ۼ�CU'�t�ۼ��W��c�9w����'�_-`ew�^����8��&Y&oN�e�-��OD!w�E0{9nA�oj��rÊ��u*��@uؓ�̓(`N�K��:G����:�+�=鳥Z�쳥�����
�7N�CS��Y[Igm�m7�����S�{D|�!+�U�Q����u�ב]� �d�Bv��԰<t*'0G��1C�S�:v�C�[������oq�fS,Q�9�ّ,�ق�gl��ؖ�<3]l���mJMq�p�>T�;R�lJ��X����v�7�KUZ�PX����qc��Ma�$Q�&��z�����C��wڝ�VmË
�gٺ�"����0� �$g"e�Y�j�k�n�5�8V�-ZDPCkd����o(�1��)/d{F�m��m�ؐ���wV�(�뾬'��I��6Mờ�	�&=���6�u�
�I���G�qn�؅�A�F�HT�w�g�ܮ������\B�<����3f"��q�U&-�6]J�ǈ�C�w%����۔ZZ�15Z�n���ݩY���{\kqJkv�	��YAA%9�&�.�U��6���q�m�E�]̃ٙA�M�g�"ݚ�T\>���������MM��Ow��J��OmOWz�ּ�#�_vnC���o,P��IL��Q�rR�>�����;��M��;���tڧ�Z�"�08�{[���IMm�̳S�ݩ}k/h�g��ݼ�.�Կ��)*�l֧?�W�������i���~�V��lf�pc{՘2���C";x�wp��
쀠��U*��%5΃���vBKgv��{Km�]���N흾YOn��]**<I���Ǎ��.-�+-*�[�x��{�h6��3J���7,@G*�N�_&<F���gU�q�7f�ଷ\�dnڙ���9��}��y�A�	�)4�Y�p������v>vxE�\ԟ{��φIQ�zK<jBi�nKhN�ڼ-�4Qjк>~��A�t�ٲ�>�5�û�1�O�*����p��0�����!��8�tm]�s�ɋ�����k����Y�<��e׎��5�ؑ��
�1�y��φ,N�(`�c�O�?+6T9ͻ�=�v�.ko�㧨��渾�r�=Xm�1�e.w������ͫd��j��"=��F�l�^�09:�����0����M���T�y�&x���*0�|�w>wpe6�ݴ����:>e�
�ׁ�]%مϩV2Iq-��f�7R����b���,��0<�%۞Hsy���/WG�]��
��~6GJ���K��r����
2��gh{ws�ӗ7"n�b��<xlT�N��	�HO�wJR�U5�D�woq��}�{��&��p�lԱ
���y�u{fy���eÑ&*Q,H�h�@�-N��	���Gg��fÀ��p�ɛ�0W_y�	}��BܽQ2��3)�p�9�L��L��w�����9t�ڗ0ǑV��N]�IJ3��%�ݭ-c�ݮ	�HGX. ��޻YS�gG�6�-� +V����e����9;WX[D�UH6���[䇾[���s\����%Wݏq #����:a�}W�u�'x*���74!��;�ŭ��&ϩ��U}8C��M�n�㠫z]����.[G\��/+�i-���r�x�{ڏW�{]]|�c<����{>�Kx+{�#6�Q抗!�Kv:�iǞ��4/B{&��gT�drHCZ���{*��Q�фÕ�QR��6;Wwӎ@ ,һ�T�D�ݚ�ۮ�[����U�b�-�ۜ�/���k�Nܭi���М�}�����|��<�>���E��4%��m��v���������7z��������]c��\�t�bKB�u���1m���㳬��%�/cT?�2�u6mA��
dY��ո��l��#,&��Z���]I��'wK��]EI�u2Z�5u�_U�5��k��G�R;�*u�w!�w�|�Mf?Yn���cK�9r��x����S����uo��il�<�r��/X�L6KY�촞h�	��%^R}R����0�,;w�k�;=���hR��F���P�i��D�Gm^5�ٰ*p�9��־i�2�u��${��9�Z�e��cD\ǃOG��㲕=�Z���\�x)\�}P%��	��I�I�z����������o{��7���ը�1dbv�����Ǆ���	g����lvoC<��n�� Ƚ�2q9�{��yH��1����C��D�U �7J��Е������1�C=�e'a�#��ѓ5Lm��q0
���ad�U���mڏm�}t{!�y+�n�5Ґ�׫�򸍊{o�	���8f��K1p�;����;%��1�Sٝ�o��"�pI���;y�"7]j�W��C�To��a���"�X��
7&૖+:������6���+����ԑ�.j�g���wO�UŹ�/��M��;|���Y���f��>.M�"O�Zߐ��,s�fG�a^s
e*	��MRwf=�������7����,�9k���0�ti4ODķcX���vN 1��nt�j��unak������(���5�U�g����v]I9:
:��WG��XN A��D��M9wY�#��ə�{�j�(;d��b聲��+yq*�=+ �-�B�(0�3h��S7p*�W0�7�m���q��HvwOkJ��"��&PO��]��hEY���}�>��g�����Onּ|�-�ɉ��ʱ�B�KL���؂���gA���,�ݿU��g�P9���
�% yr� ݮ�]�4�:.�ʔ��L�ӳ���Nױw��w��;J�i4��[�T�X��H^�֚�}�opK�A��$us��;v�臐[��3����Bk��r<׵�M�i��P�	dI����l�%�%�w��mf8p�9�t, T�&���Eb�#j{��wf��i[�ݤ�$*�ț��[{JhU���c{/�EQGN�ry�3�e�GvV�S�{��Ӯ�:0�śq�x�{j�0F A)���Y�f�֍�Jeo�D���u�Ǔj�q�z��T*:<	��lwvE[�]t�Qf#���`Jw͜|��u҃� ����A�����T�Q�"J�*�b���*=K'ӯ&��	6��6VU��-�w;W*�f��0F����2w�t��޵��N�!���+8 �ӛ�� pZ;#Ɏ�����-��7��gz��o�r����8��u�4vQ}FeŢr��Q��G��ڕ�\��c����L�����TX-�W7"nf����,ݯg�Ă�b�����F��/Z�i;�[V0�WO�W�a�u�r`>t���z�tݫWw@��<��C�7��oF��'�$ߚ}�L�I�m+a���n�ݫ�$�9e݄A�(��9}�Kz��ݹ�X6�y(g�)���C��/v�]��n��
�����>c��e۝�����˽'�%�ňi�J/��d��\h���جlL^3��<�+����(5���#f�-��x�t�y�b���#����&�� �LS3���7r��I��V6� V��Rh��E��<�L�eK{��A�ݼ͚ �J�H16�)Ÿ��؛{Kszf�Y\V�װJۺ�F��)���u�8���"ԧ�4�[[K�G-](���,z�^�ɇ����Ŧ�;�%�/g�%��Pۆ$���E�{�r��$�#������\�&�3nDDt���:��3AkɆȋ��oOds|���9��h�FP\^�@�wݤ!�rᚗ�OD������=�"I�w<۫��7*�XQ�/\�[v��<�R�������V�w��Lu2,���;b�35.ln�)�w\k�ڙ�ךR��w �c]���Ό�f���N�7��B��{��@�61f�[�eɔ��N<��*��y��zX��Q�Z-��O,j��vx��f�ɗ\�p��wMD�`}2���!�m�s��f�xn]ʶ$ї���G"�ܴ$L�"q�ή�F3��>ڰ�+����,l���o(죋�,��;�6^�q[B�N�@js+z�@\`#C���P��c�YKrZ�(Vb�T���S1��n:zqs��#+�37�7�Ѹ| �5w��c�8�������<2ٙ�ש��%���.����t��ҫ�.7�ϊ�x:��[��M�m�ng��;1��h�b{;�@oب����x�-˚�o���ӳ釥0��-�j�0j�	�3�K���1I��^��2�rou��i��o��m�jK����3]���qBH�i�ȅ7 ���� �!qR�>��h���h��>o����'�c��o�����~\;f���9����F�Kr4�HK��q�q��GG���g��� �oe^Զ)�#�f �H�����N�ྼ�է<_h=���bD:	�H-c�p�kE_/�P���:��f��x�r��{B���3�hx�X� �RV�I��ܠ�j�p[�ʗ!��i��	!Y�E]��\�zq���`�%�yȽ#ˁ��������Q����a�Wݣ:B[��^�H� &U���kT��������E/�.�0]װG/
��	�8�z0���xD���V���aY�=��m7�����t5�g��7C��kY��x$�$ڇ��V�]>eJMO%J���-䜶�f���w+�m����A��x�]�'���n�M�8���=:mo�p�v&���Z�Ļ��Նm�!�n���2��l>\�Mv�Fޱ!���K&�/���(��i�Q�g +����p�������ٖrc���Sw1�4,*�[f�Z\�H��Z�uCw�4��Wy�WC��B�p�t9�/~�燸u2M|�#�U�q�q!������j����n�m@Zr������1{��1��>�caf�+���i��s8uq�rg�������T�6p���lL���̃�"gAu̬����ϕ':2n�wYRO��%c���A��l��@1�Zf(vr;J����Te�y��8ǙG��������
�s%ں�l��7K$b��YcZ�L��sz��J�in�����촙YR�Y�2[����ʹ�h@	h˓L�H�	fyȁj,�����ћR�WF�JDJ�Z_>�~�x泏�j����l�\��lq�`aU�C�Xj�]}S8�Y�k��*��)�������<$�q�[�Mm6��}:x�2m��\�[o�@�����n%h(�,헳�_��H���͈tT�݇����#ǭ�q����V*V�X/z��=�:u��:���~�#&��8�X��@��qų���L !��Zg��#u\�5��^k�e�f�G5��NC"R���r�0ݚn��t ����i�@$�8`��e>Z$� 7>]MK�F[�GFj�z!�c�4%�x����mU�3����y
Y{Ӯ��Z^��oǨP�8�k�T1�kR�w��f�3&%�5f�N������Z.���cs�.	������O��h>ɭ�m�5l3�oǑ�cm�Gz�s:$�֟N �ù{dR��A�(�{�Tڴ\��媻9l�N�.�W9yI�~5�j�$J����u����l�qD!�4�����'m�m*��F&=YH�+�����8��܃c1��˲a,�@MOZ����<�w�k�i�ڻ����8�w��l2�(��1�&W0	(�O	����{�:L5��rCGsd��}�*.)��S��Bٌ���`ӝ�iY\�V�[ueQ(�F8V:̸��af�G��vG�e�W�������o{7~Vw�$�R�˂��ٖ�� ��v����.�yn �XUْ���9��I);7��awKTwЁ@J ��Ihto;���.�=�1[.���G���ޗg��
p�wљ2$5�Lv4�����ا�q��ɹ7ȻQ7&M��d�
�n|ޝO[V�]^���V�����-���h����,�Pp�pp;sku���v�Q��pf�	�y\���s��J�����Q���W'�5{o�y��m�g��Z1S�0����fyC��#�TgZaɂ�	��C'��]t�'����m ��o��g'�ށk�a��#�\h���t6<ǽ�������a�8��^HY��j�[2��;�L�Y��ٌ}cg����w2f'��>�4�ٝ�b��8�]���B�����&)ʅb��z����D��6/A|[�-��ܣ|�v3�l H��ygK��H3*	ES�v�K�ŅW����籨�\/�wq���F��
�B2J�Nn�#�y`��t�������~DZxE�{�3{��m�
���ѵ�wm��5���,��mj��{�ݮ!��\	x�n���%pFa���my.���G�{�G=�}��)�`g	{��,�Պ�%�9֞;�2/m���O�)q��n^S�w*��:����ᵥ�K�74�f���>U{��N�G��][N^ȟ:�u�e{�N����k��d��O� -���:j��\�v����밎A�{��;ܢ$.�PS�E~gNŲ���kY��]��u���ݴ�n�I9��2���i���&��@��{��SI���Ĺ��ܼb)S����@��v֞��<md���nn�G.��+"���:��p�����=0����=)�v��v���z�FV;��8K��%ȺA,�=�O�w����q-;�'LD�r�p(h�۴yۗq�:篷`]���;����FwE6i���r�z̭���h*�C׷�滲�1|�S�N��kV�\N*��7:�r�f�!���5�R-��]h5�]�z��7�fx�G*���C\�ɽ���|���5���x��7�#Sz�Ssg��Z�i�e+
�]��U�!{3�	Ì��E�+^�n{=��%�,��|�x\*w=.����wHو���*��gmI�F�N�6d��v�r�^WN3�5�-���V"�����(�����=��������p�*��Y�NU�o��9���Ϡq��{��0�_���1=�sh��u-�`�ۗ��,�*�g}Fkx��yʬ�|��RF��[u���Hp�D�'1֯U���/`�8�Lc��&��s���D�ZYr��y�u7������p���5o���-���Sx6>b��7�t���U�Pq�ڳ�5Ⱥ�qm��1���qi�Ɓ��Y+~�1�ׯk�����l�4),���wep�%1�F��4gL7%���4K6�U�T[
R��͕X"���م��M->>��w�[�r�}��^o�N 6�!�l�Ng��b��iRw�NwH���m����w���y*c���WM�������1�c�8���A�+��1L�[�{��o2K�a�t`�T�h�_����U���tz�=�,t3��8`��<�|��w0�"/i&�V��{�gt�8�Ưŗ�|7=f<�b�ub��]&��l��*�QҾ7�g^^�3��mA�0 m�+@��ͭ��uuJI:5���9v!
r��=����9����{<�z̕%�įH8�W�.R��TW�Y��GEk-
�:�c�v�w�g��*;ΘV �t����u���Ҧ��_K���á�@�fI�pY�����/�Ȗ�o޳W�5��iѻ�o�������;�#��3�mQ�6�w�ƙ�+ ����Goku�]
����.9nt��v�m"7����y���@��O3�⫅h1��5G{�$��%��4K�6���T���t��%�^��1��&����r�<��<�6�q�ӛ��?��؈֭xK9v���1>�F���+2��1ɭ���z��=���}sp�����%uun՟��2=�V�v5\@��|�Pwu1����;f��q�5$�u���^�cx/. |�}��=���t\�C�-Spxܥ{��7`�ՉU�#�X��`��c�g+Qnd�n�z�.���μ�dA�5-����oR� �q�Lee=w[�Y�鵓wl�٩A0ݪ!���#u���_+��8�E_o> ���2��z�,}���ڎ�toQ��P��3idڕv��l��l�q&(�b5G!�ݷ��u����6����;Y�E0��g�K���3�[ct嘦Ǯ��^0�F�e|}�4�tL-��\Ή�U�q�F�T6e]�Z�Vk�+��\��
���*�5�:�荣x8��fF�5U��y;A`���B�H�^<3�P,�\�G{͏f���D�����K�]���K�):
���W�^�L���9s��aTs�NoH�Ö��]۰+�x�&�ܔF��*����ݴ'뚏U���툄~�͎۫b_��k�l��W=u�(��v�l�oi��شĔ������/`�p���0p�[���o.��¬�L+f�:���[�|���9K�T"`���hH���������7�k�A]Y)�Ԇ�f�5�M�]�I�!Ӓ`j;����~\��IM�G���毉�b�|���J�W"�t�֌�*G?�����J�k(��e+FvL}���+��̀U�>��mk��ep��%	3F �[ݯ+k|h/����3pP����6v�ֲ��\�4����,��i��&�#�4��.�V��n<�|�%;I���6=VG��G�!�+������G���$.YwՅ�J���v6�k����U-��]t{F\̝�N7���<�m}�1mK�t�U�r�v�w}�v�0a;��a9��Y�A��:M1�v�N�TZ��.�&��u�	��)T�Z<Q�>�}Oj v��6n�\yί_�rN�NU�s�9no>U:������j�Z��'�h��8K�������ef�7��V˜�R�g=oaS�:J[3�h��U�Jz��Z[��yd�91J�s�מ�>�y$7��G��T���)���%�aQoee`�����EM:���&�/*.�IQ�+ڪ�#.��gY����l�珻
���[A6t�3y,x�@�ǿf+�����{�f�{ޏz����|u�2����[U�;*&��ԣr�l�c�֗k�6�L�$J���k#�j����SN�f�����0� ^~` # ������0?Dl��b��y�:��el�s�Yw\s�'�A�����:mbH����q�d^���w|��$]^[����C)�۹�Z�]��q���T�_@d}2�)ow�rN�h�)�FMᲷx5݅����v�2؍q�CW�mS.�^�fh\�;���m�L�G6���͜��ŞXu����1��#;Pu�ȳ5�i=�19�λs����f�"FG�<�����u_d�qa�:���u\�~�g`�e����w0W�.x�,�|��T��U�e���S.s��Sk@��QG��v�u�Z�ɰ��^�24{k+��ǧ�hU�9m�޺~�++��*�5v�_:'i]1�����}�{U�h�_dĜ����$�
V�pk�B��/��}�vf�)����Sv&3�����{j��g�̖�����N�s����s���F�Q�䚾/"��vcg}�-$�N  ��-t�a���.�Gb',�;�b�Lu}�gUཝU�y	�v�uf��%�d�z����REnr9���6#v� �/=l^�>����3y&���'k�*���|�i��Հ�*����k�ʡa;�i�%��o���b�{�{X��9��|0�j��q+���xs�:�ú�]�ҧ�< ��n��69��H�]w����Ak���UE�
��wn܌۞�x��$%E:�{��99�Uz)��[�{�^㈻��+]\��D�U��-�-r��6���i��<�%M�N�QRN圼R��*Y��RWr��!:���e�:n�54��J��9E;���EwP�4��]�E�<��\���)�<*5Λ��,���B�U���ЭJ��*����O �XGN�*�I���!��4����si��A�E,� %��+��d99穘x�"!N��x�Yr��z�N��zZ�2�K1H����UE��y+J̈����\��G(�Vs�I%�A!U4��9�p�0��]���zQ+@�Q-�9{�x�RuBȬ$+�^��"\ƈ��|���̧���V���RK@����UM�;m�P������<G���d���]30ͦ�f鼍�Fܭ�y,q�oW�g3�0L�h*?��,���<�|z�}�s�-�p�n����_\��a#棽��X�0�芰4߇�ر,�(O:��qX�~{�ީ���5�<V+wΝ!f��198�Ċ�2����7����˱zf%�j
�6����/�V�2�9��@��D�G���9�e���$������N��+�+a'��S�*�Fi�F,5�(��0�ʳ��F��}~�tʓ�J�c�aa�����\0�]+�#=.q�Ȇ��gӜȝ�;ꂮɛެ�|7�O,v{�$��U�>�=T)��t�<(�����T���I;�M��+�f��y\�Pn%5��,�Gؑ�=^REg�Vt�,��"tW��\]=�	0sc�.DE,�J{a�1
Şl�#}X���v�؃=�Ϋ��Βt��3���5�44(O��\,�Ξ�s�r�e���a���]���uG#!Ҧ;"�GT@8M/��I�`T=Υ���Ƅ5�,�{�X��N�yO��	�6��K����熈ck���&�V�ƣ���T9w��>���{/�%��9���_��_o.�1���XU��z��⮝�ʵ{�%��J�7�3 �,�E��_���Վ��Ǳ�.���!xUr�(^���zv>9�sl�R���i�[Z4�j��m����.�p� �c��f�
m��|=�I��JIoa�G�#�V���zi�0_��i�5'J�d��f����]�LP����Z��v�a�cf7I�5;�N����M_��(gy��&���K1��B�37��]���:ȡ��.&�R�|��\=�#����O+C"�Dų+�;�.�Q[]{PN�ľ1YV��$@f; |��E�����JG�*�
!Q��7[�2'Kj�`ۥѽl���6i�8Xc S*L�J'�@��8�fk�Ѯ��v�yN$b�B\���s�M�v��Ϫ�[�ɓm���<�uƙ%Uj�u3��:#k��t;:�k�7 z���B�{�V-�ai�ח9;�1��̚�.�N��fl�q�:E�.��dR�q�hyS��yӫ�F�f��t��(1�h0ڧ��0���é��p�*p�vΩu��~�"��2�|3�	0TAU�9yրz��
\�3��s1q�hf���w{�9}����P������wu"�5x�ۢ���E�R�X$���
�_Id_˕HH9�\�`8��5��S�n�;��oB7�U��6���Y��/��Q9���iK��`u)$@��������]Ƽ�D;����u��9NVȪ#0�Ϻ�f�ѱ����󵩳+� ��Ge%��s�n��f���(�+�t5���}-띦ȉ�ۮ~k+��:rLUO��XYZ뗒�_*�CQ��Y%��8�{���	2N��{\[�0��Ϳw��Vr�t=$������4�ʳkwmw�� w��(ܦlL�*E�OWֽ�`2����L�v��f+L�x�R�є��Võ˞���@�8����E����)��;c��:C1�v�5p��1#���!+�72	猳*�x�!��Zk]�K�K8H�U.����AF������!�۵ǯͤ�if[�����|٪^�τ���)�Bj����=�~�u;�a�0��jxK��kS�.{�`�R08�%T�G10�JtҸ���ң��vu)t����j�5�[���;X�n��+TH��#!߉�|'�
k��^U�� mS��}Z�qk��g(����'���71��s8�p� ؅4�@Ӑfc����O\�5�)�Z�VwF�BC����Έw_�'fJf#x*����vd���p�lS��ٮ����S�n� ��{�y���.�$��y�n�7��%�
v3�[5���/�Җ�pQ4M����4$R1gD���y�]#Sf��*�Z�5zl`y�y��7ܝ��'�Ƹ��c̡j�K������c!j�7*oV�����d�N�)՝5-p���z��Fr��L7ժ��:��/B�d9�� �jpz�k`�}L��e'���0��y�׉��H�y.����ƌE�����NC3��/��u���z�dh8\4����������+��h�1�,vʌ�V�1�C��dM
�;g�%]�rB�\%^|n5]Aۅ���ɂ.�:X8b��>���WwP����U�}�@��CϤ:`����fy�K��\6��p�o���oi�	|o3��G]i>]����v���J����@-F�<�\�yD��ޣ���Q��h�yR�%�X�.'w��ˀ��a~��P�����.�,��<P��#����_+l�3r>����xU�_���������+���7�,}ι�؎�۽�L1�d����mȳ
����:>�?B=�nKu�0~�< �+�1QS*C��wK�陧�QG�:k�����ޖ_1���p����#:W�DD���ܝ# T"�
�RՑ��7:��zM��Y��1,]��9��W�P;H�@�Pr��kZ�*u���=<����A�O��J���&����uo+a�f�O*ܶ����p��0ƺ;��K���ţ��������޾���fԋ\�m9c��w�̊S�X�Wl���j���^����v��$� ��Q0��pܑm��N��)uǏ�JG����<�~ʇ}:&�IvY����||��5J��c͔�y���M��T̄IG>��Gaj^T����qg��>���J]4%��1�GG����Z��1���DQ9T�%�5Ex�M�3,q�g��UҌ�YH舫3�=�y��*!��Q�JY-���Q�PQ4`Gi[aD�jF3��5PDLiD�!i��un��etFm�^\���mU�����n�,�{[u��b����Jχ�ؿ���r�<�饜V:ߞ�{��@�̥u��?Qꈞ����0E>}w�=��M�쨎Yv4+��F�EQ'ʽ7Lf��	ә(�}X�k͊��t��)�η~�*aዄ�V��9��W�4����A�\�}[����z�B��*UT���v��z�C.���.q�����5|�^�T�ȸ�t�Y��MV�:��.�d ���bbs(M�Ñ.�b��̉\���!�T��i�����g��4>Ψ&Qб빺�a)Q�9k]nV��S4on8� �#�9/�C_m�흪����������	�Z��Ƀ��sn�ˌ����Pt�������n���c �j�8eks�)�h�p��:�c)!j�Bj �E��؟f��u�{��0Ho��֖�!=�+��tTt|�0$�͊���Ȼ#(�\�T��aN�^����9�W�˭���Z�N��=���t�{���P0����Խ��:��o�}Myxc1��=�LJ����h�ɉ�'j&PT+��F:�p�dd�f[���Q�
�%�ZhM&���jK/�xh�6�:���p�=@�`��WI+�m����ӝ�.�e��H��V���zj���5��-��d�쨇0�*G��ߜ�Z�w��G��蟮����H�����S�+�1�W�/J��iT5���w^E������q�fD@j��0yOQ��aLZ��pF
I�C�D��7����h���/��`�\7ՠ_Z����Hx�!|��3>R����u���2*��ɪ�q�pQ���s0���@�f���!�LB�Rg�& ���i���~E��,X	���GѬ�����MTV�2d��k��
�1D�5����LxX�5/��>��MWK�.qR`�l ;��ZZ��-��q�%i8u%G�y�W&u��Z��D�^�w��y[�4�Y[4tP<�d.�nY���^��J��V�{�P7j˴�h#;�M�B.UlI <~����zF��;�ӷ�"�6;w7�R���)���{�w���\F�^\,�N�f��&�ܸm;�7ő�u1Wnw�:	�~���.�v���Tj~�0����W:�b��(;;F�Kێ��q��|7�����י\���McUV����'v�g�0a�qSLp�δ ��P��R���Y�W5�+q2��h�?)Y��Ք=K�~;���O<N�S��?��XRJx��
��FD�[d%��e�jNɑvT�}G�_�]w��W^��_���ω�� �^�b}Z��h���g�,�H�zl�F
�'��V��~a_�����p��M����x~Е�!C���:�6�G%���LW��(�,s��἞���;�@��� �����j�����Զ- ��	r�����)��;c��:C��tBj���}�a�qy7�߰�q&�W ��HtMv��WQ.�,�!Ib��[M��p��\b�
.�y�B�m�j⅃e�Ub�P=�0R�$�U�U���Ĺu'4'Be0�����:���i����2Ȯ��j�]�j�BIԻ݇���"�F�`�%�+ �v�͂�Ղ̽w��#Q�%������Օ���8�l��Q��Q��kV����bq��%�$+�ty���_���e�M�5%�s��(��''՞T�(TH���mQ��7Ჸ��>�3�)�yW|�j�X,�gֲy�tCg"�`7���Ђ�%i�R�hBx�N�_�������[�X��n��8
S1�[[NJF4B�2^Z)�H�`i�3�D��DAi������8���+��zcx�=�Έw�1P�vd�Bs��FE{eْ}:�Q�.�zma<J�}���b��/�F�!����N��	��j�"jq�]a�9���M�?�-�]j�<�*�]P[�����+��ͦ0X�,?5T�������dk]�\�E�^�+|�,.��0�붅:�0�c���YM�����e3�U�Lj�c������_�Z t���;h)�/�}1Q�x4Ǭ�?�	<oM�D^��؍��ܼ͞o�oA�D��?<j�䩮e��F1��������3��9%��U�cFm��l�uE�&#��;At���5E5<�)�ed����Q��`鎎Be����ݱ}*w�;�3G��݆OV�̠�j�ȝX�v��i��t:J��l�'(�fCb���=�H�
[����7�7/�=<���Hz�7�Wܮ(���VY�LJ�R��a\I�R�-�x��.M=ܤc'Wn�=	�ECi��6��V*?QZ-�@�|.��5�b���k� �9B9�L�;�[�@�Ѽ���Yt��Y��*Q�� F�s2g�	'����W���G`mތ|&�r-@d��ۼ�{r�n�ó$������RkG]G�I�W�h{�Fʐ�v]ĳqEi�4�B��c������ �����.�-��.n�6�hk���F �E^�Ԇni^qJܗN�w(B�Y}���B��wfY�,�c��7$GU�de��f��"&:��.��UY�C��QL�]��u�-n���@%��)�,Fx1�kغ�v*vٌ6R8�V
����Pq#�]�O�N]�-Д������?�'�s�ОSg#,;s��Mu��9j�9 �d�� �Rw�њy�˜o�uĶg$��L�V'��zN�&��q��oR���g���,�TJ�v�p7���s*@�b��MltE.>'_�
M�c��=ӏUxk⺥���޴�0��M��)��t_���K�jŇg�zY=P�u��"��z\�>�Lݜ��x�Q}0:�V���sn=�
����x���)~���Z��2ygV��6�L��G��})���t��Ղ�k�,y�}��K�|E����ѹ��T�X`T:sQ��Kx�J��S(��z��0����擇f��%��[H�ȡ՗��u�sۤ5=�~F>s;ѱG�Lg�Qů��ݪJ����b�V��y-v¾�Sd��ޔ�u:�F�i8�es���ӣ4�#c��! ���=�Q����U;�+b厺���<9�(�k!���WFD��{����1b�s���ʑ9�y��}jϾ�3U�U
�|;O��.��̌�I߁r��]�p���7�Uj��zh/Z�OY�1��A%����:*:?�����9��"#0;��GxŔ�K���xkyl�t�b��=���hm��N�H������^�CB�Qu�N�P�&j�^u�{����5ON�ǵ	�s҆����b}�N��`>�I*���H�y=˼��8���L`qJ`3P9�S��Ie��!��[�.	�U�`��e��u)W{��t����}q����n�5X���i���%�eC�B gi�x%���^>��3��@�WvO�����jr8���p�����8n�����d�f8���u�**��"��7�Z{�n<���������j� �*F?W�Q�Ir_>��m����Xm�6�R�c��7 ������]sbK����YY�[��pec�$�ڬ]]���NJ��륄�4',�O�K���Z���8��O3b~0�J�<�kc׭���M6e���JugS��i�����fgf��ó�A�\��-�.�j�;7kC��%�F�E��qͬCE�-���h�*>>Px,Ք_��<^���=v�n��@G�\�ʎ�����dM�r��U��8�2���������ȯjn�S煖.M���ʉTt{֯cT{��jq�n�9cVjb����0��f2����t;��,,�H�{�$���5q����!�����z6�'s���u#�v��*H�s罷[]/+c��D�$q �\+�ݏ�hm�K�܃��a�R���<��/4_��c;.�P��.q/4��*�2}ӳ����7�J
L�0U�)������Ö���tp���<.�.^�=�7���A��d9N57{7�M.<����I�W}ĪZ*��.��ܬT��6Ϋ\Tm�����2�t�^P�0������;ӹ�vĮob�ͻ\/��Ԃ]^5W{xkz�d+��xZ\��Ǫ�6nXH�h�{ �ʲ��b�}��壮E�����t4���=q��5�`�wLC�$ov]�vU�`��-�A4�#�����+�����=���C���)> {�T��������D�ƥ���g�s�[չ��j���e�}!�vaR겵)��^�Y�ϳ�gأ�+�*�m�܄��'
����ɶ�Vv��5��6��]��[����h6����+�rW�)�=��>~x�ՆGX��kB�wn�Qgyt�K@�nqC�g�pqgL��`����������7R
V4MkdM����
�DuLGV�S��D��v��Oyk&�/�r�v]y�̯/�ݱ�J��G\��⭮�G�����޹Zì��A���K��-�qnB�p��DjM��{5�[	+bҕ:�˝�&�u���b��{��okNv�[��^���Z�G�";m��������0#���	�1�g�%��γ� ���k�R*v)yv�M>0��� ��<W7��8�z��]�9�yk���/g=^��o��IaYf����|�N)�M���R��F��ebs9�m^��qU��{�T���Q.���*�aݰq����I7&{MT���f�
�l���Q�5e'�B�6iI^���o�ZC4���s[��{�;A�N�5�WŒ�u��#��Lڇdm�tX���W�|�����o�ћpTk�N�F�����vu�8wo>H�*ߗL����j��dZ��# =�i �6w,tɸ�ov+J����\0̼�v�WOL��ax�p.��JJ����%���"�nL�t'u�XɄ��81nӛZt�j\8�Pӿ�4�%��g�Z���S�"S*��ȩfEȋ9�*�GP�ws°�/!�ďSn��bQ{�\���)0N%TYQ*#=pNV�г5G</ip��E�u%E�N�E蚄L��"SU�y�I�N\�˻�:d��J�FHE!$z���J5�-��AAzģ�9���m'uÖ�E�\��%��Z�J��UN%�D(XPQ�t�%wk�瓲�"�6�Fd�U��:��HA
 W0�"Tȑ
�Q�P��g"����I��D�ŕ�*�6r���=H%I0��1DH�]��B��ԡ:�YkNVI�D�Ȋ+M8���B(".G���LLȽ[<��Ri!RHd�*s�#J�# 8 �0 8@}�4��8����R�X]+P��e��Tp�l7+���f��]����n>g�)db�v]����nt�"	����-t����>�s����lx~!ɅS��c�BO�ro�:�];��9���Ʌ��G���~F�!�<��xT��~������>�|=���w;H�'��������_��{�Dt	B�����[�Z��{C��ۓ�7��M���v��?�~�c˽�U�o�z'���	8hߞr�?��7߰s������>��ǔ���ro^~pxw��������ww�v�x�Yy�2��c}�'+����bC�a��������s�;y���yw�k��7����7�'N��}_x	7�N��/���!����rמp�GN�o��9�{q��\|:b8E���f"	���J���27�K�n�=����=�!�H��b$}�O�(y�=�������
��}���yM�N;����7�99��ϯ߻o����O����������|�rrnw�w����ob��GG�1UPQ��7-P���+V~���v>s���d�������t�=${���\����~w��o�^�{���7��>����yL.���|����ǧ��_���Ǎ�P���;��n�l�w?����O�޷h3_,�Hoc�C���4=�!�.�w9)�����#�,�DH0���?xW;HS��~v�y���y<�����۷'*���c�o�O���6���y��?�/��{�������ҧo4o�9w�{��p)�q��};׿?3�՚'�TVޑ���qC�=�=}�?��ǔ��9G����9=����	�]�ǂ��q��&��y�	��{v�<���9���[�_�;zM�	ӵ�����.7�$~�m���7�9�"���+�F����ѿ[��~�X��H���q��]����;�}��yW�?�����^�z�xw�9܇�=�Ʌ�P���?;�S
���=!�7�o'�>���'?=(RpG���@�k������Is�z+`��{{M�H~��������ݤ�����<z>}�y@����ｏ�yw�iǣ�����o�v��97�sɾ!^�����y���i�0��c�yq�1#��s9�����y˔w�e<'��;�`���t�ϣ���s�ۓ��������o����U?;_#����a��n�|���]��v󿯉�=;xy�ݯ^�����'*x�m�<�A��|5(�ߌ��2+��X�odu.TѻQ�f�}�-�G�ecp{|@�{��<�	Qg�����\'�=��Dvj�����������L0�"vVg�l��{������W���^�����28�N�巊�B��|�&���-�;���^7{�]a����~��ŷ��<&������h��y��x��aM��}��]�����9t��r}M����`�}O�9>'�޸����z�e�������pI���#�|��#l5�}��{�̪���z���#���L��������i�;z<���m?y����I��������'��{��@{�#�9�=�1���������>a��S�c�"$G�����7���7!���<�o�q8�w�ܛ���@s���s�;����������=;㴁�/�.��[������5!��;x��Үf���8�Q�۸;8+��b���oc��87�;�<�Cÿ'��ﯺI��?P��
��㿺�~�.�����o/�nNC���]���}�������C�:���#�(�<�{��/)�W-�6�����w�?�̙L{��_�O�����yM�	���ރ���HO����x������<[s�< y��ڣ}y����aC���`��n��(�c�
��B�
��о?�-���}���1FB�o3���_�ɖl�C�S��ݚ��-�r�b����)�N�`��t�ތe���˿���G�����o�N���cǨě���<'�n{�o�s'�n@��!�#H}@|G�_���Jٔi�ٝ�3/�b��/��e*%���]�ٵ����v���r��raw�?}��˿;�����xM�	7�$�����7�99���}�y@���>����ۓ�*��Wԁ}�:�Nqd>���)� ���]_��B=K�"Ǵ{�DG���<ߝ;ô�׮��;巷s�{��xM���M������щߓ_�w8��	Ʌ��������r���x@Qb8G� ����>�V�-<�U '=�����G���MχnNOߠ9��m�,y��<&{C�[���&���o
�Nӿ�����<��oo;��v�P�o�Q떷o3�x�0{bT���t���O� {���]�����4o�qV�2�^�x��;Tny?z����&ϻ}A�����nw���{�������{C��S���x�!�=y����	2�O�?����������>=o�C�������m���U�T4�<f�w���2g��q���u���3O�u�U�%����]���yyd�>�w1�-�.�w��G��8n�+jfLk�⭴�&��l��wX�9�{�ʮ��}8r`�WM�X�8���J�w\��;�/�!$�/�qU'ҟnwt�p�^�������,���O�;�N�� s���>����w�i?#�zO.<8�ǟ�97���?�-�1;����t{C�yL.���m��.���T��e[_0բ���EQ�.��l������Y�NX`�͸����f��ާfo�8��xğ��nM�����)�~�|N����oHyL={O�='�{v�{��<��ޜy=Ǆ�P���ܾ{�rf=�DEɏ�Ei�Ac�+cp(���U��23�x�������d�1/��d�����۽��E��x������䙟S��;z?�Ѵ!����=��֔3=&O��?}�y�����zv@�}񺊪�
b���}���:^�1J��5�9��c��ك��&��]��Λ��۷�����cώ?;y��������]�7����˿;J�����&��w�k��y��yw���뿎���raw�{OG�ݽ'�>�ɇ���_��T�%��r{S�*~c�G���#��!&_��<���w�B��onܛ��9ۿS�w{��<$��������N���������t�>O�݉?'�\J�X����7�����?��?���6VM��`-w��Lz� �yC�raO�����þ��=�r���{|u���7�;��x~;y@���y�<'��8�{��&�m���kv��0v�?	O����������\�i��kx!�%y��3����$a�)�������7�<��c�=�'|}�O����O��}q��9���®�)��|C��w��xw��n~;��^I��?[w��yn����˩�}���.��gwvM���W!ɿ���:?;r�ۏG�|y@�󷷟_߸���7!>�����7� �ϗnN�`�|�:v�o���C�;�A⏯�.��*o�?|8O��CxɬF�������!����o����bw��������=&xK�v9>!�@��x�»�i������L������z@���G�<y��nM�<������p�$���x�������Ԡ��d�l�e�f��?����_o���o%��&����}q(�.b ���B$D^�Q�F=y��W�!��ɇ�{�����]�O���¸�Bq�������ѽ����<���DE4���.b�B�t@����z����9m3g#������@�w����*��9/'2�]ۻnq��f�v3ZY1'�d��3ug
diwX^���T���77p����N�dJ���uV��B����TW�h�"�m�j���HԢ�s6	��h�f�"�ބ="E�zG����E� �>'&�$G���o���]����m�<�ߝ;���ɿ!~���|�p)����<zM��bO�~M����$z>3>�=�����t\u�m0s-�T����#���0������������w�9���hz��<&|�c֣����ra|��=�_�xC��Ϯ�������.�����'�o_�}����&��>*}� D�62�?Uԛ���������ߏh?�;����xw�j���_�]�ڣ���.]�ҡ��M���{C�n���=��[����<�y<}��)�hs��Ͼǅw���ň����,�[��4Tv�e�*������ٚ݃�x�>�X���޳��x	ӵ��<���~BI��߯������zv��P~}<�p�C�|��ߓ��|C�r��S�ry��M�яAB2,���"8Dp���%`Ǘ��g���������=�!H��!?��Ǵ'y�﷤<���~�����ې=��Ǉ�?>��X���Wտ>�'�ސ�z=��o�o	��ɽc��C��I�u���o�_ |{~~�����o��h������Ǹ�#�$B#����*5>�os������퍽�([gR�\Asa�����V���s�4��-159rrN��Ʋ��a�pt������H
�k!��K�p�m��n�og][�k�#/F�p��&b��Èy�:m�0cϊsXo�*�b�0 &"�ZfFDRN�$��8T����,-s��)��v�P�����;�w%�W���G�qocL������\���gH5$8�+��źbˮv*]��nZ�� @[�42o���9}^C���_NanZ�g���*��[���L}�r�]i'���`o��Q�Ѕ��5��|nk�u$3TZ�p��{��GD���Ğuy��r]���w�Xgn喉�,�C38���iE��Ȼr��S��2��w�q�&Q��)N�nqV̡�ۛ�%<��htK0��-u+��|���q.�`� ���q�^4C-����ñ[���6M.0u�PT��������9��$�9��$dND.V��5%��4C�o��&�W���5���D�؉���2�0�H��f��[>���Z�C�^�r�	k���Rt��K�=0\�I.��Y=�q<:]u;�Q@�H{�g�F'<09}^l�6�kAK��R���M�79D�6�����	�iR�>f�*����M���t9u��R;_R��r��!TA�����&.��Mցp��H��t$z�����㽝g��U����-yⰾ��w��m�u�m�ؖ �X3�eGJ'��Bf�O���z`��[�����ѫ��1���+��'��MQ�d�����l>4�*�T:�Y噔/�_?y{�ۜ+�4X��]��K;nâis�.�G'w�3\��l����6���Y��7rn�1ۥ��ـ:}�X���<8'��1��(;;F���F�#Lw��%��	:����2��@���X��o�1�������;�u՗���[�h���$V����Z��� s����x4�ǜ_C����J)غ���4�P��6Lg2R\�̥pQ�x��}�� ��Y8�q��]��)�Ɩv"���V�7��pܞcPdo�����۹��&ׅ}��<�g�w�ǟN~ 5�^U�k�{�ߕ�>֦���I��_��{���ܾ�y K�T�ϣ��XJx���?r����K[/�Z�� �{�E�T�D�AB/�t�E{�h���uL��iL/��a�{.yv�a���Ҟzj�hcRv\pK,�jy����r�<#6��!Y���w��N�b������s��d'g�T�S\��yX�Ls���L��n��+M{UU��oQ��2�;��#�A�<H< �!zy�뒊�Sys�=p�:C1�w`{c$ 
��6b�a�
3�EeB�kO���x��Ψ���ɮ���[��%�C�L`�Ԝ���v�CV�sN4^Wa�ܜ=pX�p�*U
��F<�=a@��i G2��{�M��_l���r���z0��%�W\1nr��n��o��PY1p CX<>-/k��w��o�Or�ᕈ�b}��c�^�$�"���v��n��6 ʙ%q�R�v�k\�"y1��K4ԅY������4���W;EZ�����u+�����|}��r�%'�֗g��1k�Q�N�������[/q֪ɺgrƚz�:��j�a~C�S�Mͣ��_W3uϭ=� �٘��5�cIbt"�y_j��2�R��G����m��a@@�6"��#�c�e�o�S�ٍz��x�e��N	��M���w��������S�U�߃��cx�<����Rb�N̛�Nb5�у��~��$�Z�yz
=F�z0lV}� f*WT`8��0�(��~A'T��ˢ��u�m�,��dZ��z�� ������[@��=�N�t��^Y��$!�o[64r���[:�6�E�p�~�U�/�̬�,4��
���XQ8��lw���u.���.�߄���K�:�U�Ƭأ48�r��͵lg��xMě�c�N������|��8K�q�!�"w�
�ܕ�%��S�F�S)�����j�g�d�1�����~j�����,G�"���+Qs�@��l�����%�?��8.���4�$����<�\�y��1��l�G8��E�ic���5O�W�w:���
�'�2uPEhsA(��<P�ʬ̝�jU���WE��:��k��]�(Ѐ7(�<Q\࿚]��>�\خ���1���P~G��֖k�W�V�81��孑n#���{L�`Wy����xz��
�����ͩc3���1�"P'�>�B�-A��o4PN����v�%;e����3uk����A�q�å;�xm�9��c�K땜�"T��v�L(-M��ӷ�;V�~����H�����,�h�e��!�u燦�GX�<x"D�_y
�a��Jyk1�L����2
Ț/�u�2���jK1�d�����W҂'��=�R0��巗����/�㛬G�)�:��e5Q ��\9�c��rDu[vF\9�f��A#���'FD�D��%��~���(�K����P���΍P��f2͔�&,joh'�9�Y�����=�Kǥ��_���ך�?��|�NL]>��6���>�u��C���������J�h�9��JqףJ���2�����w{:GG�n��N�y���K#��Y� "�Zbb�r��s(��j�JȆe��(?�<��	�	�z��0�5����0(�})�Wթn�}�	��o��bj�M�`,.M�	�d�@>Zh����a�8
'�ƞ��I�j�S�])H�v9Lh�ۨ넝ޜ��'>��y��p�#�Ҽ����~*#}t�+fk�'gΦ錸������L�}������z�xD��Bv+(
�n��FG�C��3���7.u����t�=���g���|k^T`Ѓ�<�Bl�;�dc�PCYi��G�l^���>9˺��QN�wI��}���w�g��
�-�^���_{�Z�M�wZa��V��w(E�,��Y{_���}�R'_0ꙸ�l��(�ʃ:`d�wꜣ������@U�Y*��Q.q�V�7��c��y:�nZVW�^��\�5���h�U@�W����iῚ��r�>�:xe����ڲ	�)T�C
F)�����go���:�;�uW%���GUGT|�0$�]�;+�ik�jX�e�5��>rEC�֧��1
�����[Cn֒t��9�����6湥����.
f�����Ξ��;P��3�1�7Z:�&&8K *�7^�ڗ��e[+O:<����du�M-5�q��		��~��%�� h�6�o��H�ٹ{�w�'+����eÂ p�#;�R>��Z�C�^��,p��:\W���eX��x�0����]O7�It�}~�(+�h��� w�I��N�S�+�zo��x�uό&��!OQ���Tu�M��<`��`#�@K�1>�u���\=�\AA\�9ܛ�]降�/$�-gR�]"a����Mցp��M,�T��E�J�tu��3�z��IA����j%�qh��ly+Ua�א�۽�Y�k� ��+�2�C�`%��>��qr
F��Lzy��Z�I���*���s}���7�Aʎ�|��"�r�{�l*y�/s���]�рd5�d
�*)j[G1�q�����W�S+���{	�:�{]�
��*7��'�u��f���!�(�E>P��'�������<w���a/	�N�;F�z_��_�5DTZ�ɓm��@uCo�1d��p�˹iduR������q�K��DP�aI�>�Ƕōyu���rw|c#\��l�;��o^I��S��|߲�$z�<F����_��F�t��(1�h0��>�{����z���)�	�c_�����a�v���L'v诼�0Ժj���/ѝh�i^�0'���m�-���1łv(?;9�S�fs��!�?�՗m�P�ۢ�auG��l���9�4]�vm�\�zJ'�`	�mY��P�9���~MWj��1�Y<2�2����[��k�.V��S�S��t�!#qe�WK,��2�E��
���ۈ�p�{:nN��<���m�b͡�~��5�Ѯ�Pz�S�[�0Mbs����U�nS+��.��r0:��X�u�;]�{d�|=���n� �G�� !���ܔU)�s�=σ�1�Aw����.cej���+ �tm�,)4�)��{��F��D�����������k�p2��sa׵�F̏7�o.SE;F�r����MLkO��`�2�����V�e��2��-�U3gz��ĝ
-�5��гz9��|�&�wZ��4���d��KQ �<ow.�	���X�+���N�GE;��rL���mm4��&�u)�jC=Rt�Too�VO� �B��֚˜cܦ��aa>���@�󜺌jPฃ�U]��0�����+X|7����ëE�=ŭ\�#� �� �#X�u)������fE�)���`�DI$-]|{�E�����d�m�t����j![�7}Q�:�Z?Yv�ҷ{-��Ɩ6�|:gv]��2uW;����t7���mm{Z���[N��{S��k��Ըʋ1��z����tf����C�¨��*���NV�曎m��������쏮��n��L"Sq�7iIzt��V��2��$h��2�e��O�tk�[�Z�i]={�nm��<�;KIFQm �[U������]ZE>Xw��������괿D�"Pݮ7M�]��P�c(��f��C���{p��I�[�QC��{;\F,6���3)��X�L���r@)�<2�w�&�ވ;�+B]㧓1aU׷)wv�� $t{E���zCW9FU��=���\�oӻM�,��:��^�V+��9o�۬���ۀ��0��H ���ejծn����f�nV0cN�ϋ���s�V�k���f��F��Z�>}7.j�ں�OQ"�y�|_���Q+�G��l��nP
� 橷Z�n&��8�/���D�2�L��]���m�H����u�7/�V�]����� NM�c������_�8p�rH0���#m���ۮ���u[鷓���kIu{F���=���!˷�NA:R��A���T�̹D�TUP�������M�C^<�{t׎��9���^�26�eY��>�1�9vQ1'�9ڸ�io6���ZƩR���ޔ�c*ւd���/e��7.v���vwpҴ/��m ���*[������@�4�ҁ�#j��T���	��ZɻH�%
�,�ހ+'*+c6�̫��X�,�L��w���6�(��9Vicj
�ss`�f ���jj�;�c'�z�y:fG]X'^k[5�\9��ê#����܏��uEs�m��+z�X2�[�����З���q���y��nX��͑�U�z���.t�˥��EݭqVmu�dkM�=/��,q�;s3C��A���q��
0q���V�]��կ'��8h�Fy���{�O��Y,��g��G�ష�0U��ӭ�ok��r����ZWs�w���k����*r�k��MJ-���2�x����A�gT;[E]����|��%��*��Q󃓪비Q�(�{����G8�
�CȔH�5�BT!2֔\��21J�*�DQ��*G$%��1sL�(�*I!�*��r�Yj�ʒ�AI��kTHwwV�5*"��&Q�AP��R(�@C�^�A��.DL�H��*��VI*	!U��re'#
N��^��EU)Qh��9,3�j���Hd�b�I�
Q��"�WT.�dVt
9		EEu1i.�(��DP]��*�ҬB�2��Ds�G.Y!'hIXr��9J�TUUET�%Bejs%�F��MaEr�H�H�g8r�B��Ud�$\��R�d�l�����Q�k6�f��H%ʊ(ʩ*,:�CR�Yr�%:Z�HDE%�]9�jF�MP�LSe�Q�*��ʒ�4�Q�N&�VH�m	"�C�j�$�.U"��@��y[֡�yܹ���H�¹T�Q`��mz`�m/t0u�\_��n>�b��Q`��EzGn���N�)����	~�DG�;u����٨o�{q݆m�����OQ��=Ċ.aq�u�D��K8Hqt@�ȡ���½��� ���ms1����,p8iR�V.J5��L%*�l��V[��h=��|�718��!��q6��pf��Ά�&������H���!�<>�v��!�0��k���ז��w�똘�W�
�>ԝ$q���C������qL������UF�Ş�bnYZ���b/���,Ezz_S1�Z�%����&�/��f���殍� S��q�[����4fa����R��B��5u�����G���F����TLsy���ۖu�h�m���YOT��q�<�b�]P>�MNu��G�7��Νw�N=6�;�x$��cYf��5�E�羶�z�O1��X[�漳��>Wl�za���7]�w�0V
&�����x��K����yS�hS�0�:߇PKjf����/�S�ġ�]��E�L��i�Vm�c �J���s����np�y0E�O���6�ϖ�쥱Rkc�ٶ��ʳ��']/8�8\�ul-�A��)�8ኃ��q�|�}0����+A���y����&�X��F������h��Z|�t�導�Ugf���>"{B|�lb�O�@�vcҎW][|c0RX���ģ��#��i}�����nX��eV��L�%�و��j�䩮e��c}�N����.����1�k1r~�ɕ�S�ڎ�JuA/�LG1j�:�
��1e���eN��1e�q�(Ի]��g�����>��ra��M��-�+LM/
uKc̭>v&��k��uw�;���Qvh)�5�g���v|U�;���Z��<U�����Q��.�3|#b��;�$;n;x�L<"���>���{iߞ��&�u�G��	1���5+z��$q:M��b��g=�#*�W��7GJ�eIf6��N>�3�W�x'�� �cu���.VfyK�Y�<�C�h�U�\ʼUcx�+j��=�����!�":�m�ni�O2P�,��Vr�y��
�D?8#�.%:��)�#��5�]\;";l�^�E9��ʘ��l!�9��4�Q�W�⃮H����BG��B�Z��E��[k���:�u8f5�21U��j0�(��L:�"�&㊈턫��h�G>v�wU���US���e���[��M��Wc��mL/��al�!���M�6���ػq);�׳��Ro�m�i2������,��~`�[���i8̈́�e��>j��p!���kB��5-���ה���2Ir�__�ൾ�c�i�~6�F���ib����+����w�1�|�Q?q�>��2^C2���!:�)WN�"i�Z�<�REz��f�vN�[��kb�8e8�q�*<�15W&�# 0�`a|Ջτ�K'����~���k��`�j���V<Da5�go:aՖ+]wK�u���V>���ZI�\<�
�$o�/{X���a�3R��u.'��L�{:��ʘxa'���wH����a��j�
�eo17�b����89���\ENQ�7�(�ֲ�t��U��l�a$�{'i�5��m��9�]H�W �5Яq���<7MF��� �����k��;\�h��kl�qM+�t��W^�7�p���qe��>�d�^.���m׵�c9��SV"���Pb.7$T=�n{b�1
�.�1�W}����@�XYٷf*��~-n��еy�Lb5���UB����!����3T��7Z:�&&ԋ�;�����2#�;���I`
��9�a��逍�	���jK:.C\ۮ?�x\�1�h����o�RS-�d���W��%x
����%W��jN\�"�˞짜����y0V���/���j����}���+���=����k��[l8@-T��
�}��P����J5+k��c�nA3u O���M����Xj'�k��=��c4>��M��+�6
5�K|:y��2���ڭg���C�8`���Fi�U�щM�S�S��"����t����b�u^��c����ZH���N�)��N�h�9qׯgL\>�*�hՐs<��,ny��&�1����K>�`#>� %I��z�uk�w�ٗ�[*=T���w�Kذu]8{pFڤS��f02i7Z�Q+�CՏ�A`�U�ºD6H��H��T��;�muy�&1�9T2[s��� p�0	UJL�D�C<ݱwd��L���GC���}��j��Y��S����~MTh�L�ԁ��T4w��6����;g ���]0��\m�����[�����޾5A\Cc����|>�V� ��kٛo
Tf{F���i��&����M�V$�^Á��I�����6<9�F���6�F���>YS�zGC�,�^^{x,+��9��pg�`�S�+�m�������еއ���o��\�3��s1|�i�}��˺B�BwA�g(�?�"f��u��qZڨ�ؘ�F���}�s6x�S;6Is��s�zg�>���hu�S�JW$^r��V�YH�OPu�Y��\vY9u�;`U�El��m^���H�ll��1�6,�X �=|5+<�=��g�sJ
���lT֍���?�ff}����MQ׻���2�+"� M�VE��l���b�&��[Y\/:rLW��xcHf�̩�q���ru��s�]B��n+�!�ge�VK,��2�[�0��͸�p����eS6�9��*�M�}qi}D�F�>�[O���'�ҵ���ea�7)��ƺ�P���H�`bW��"x�i��E9 �(�,D���9W��6��w������p��\��-����&�g��>+�{*��*��ϕN7�n���/�����n�=�A�$8ڞ�hª�#���p8]GK�Z0��{��AѓP����^��Lo=w� ����y��O�%˨��r�؆�&���^n���q CR٥B�{/�ֻ��x�emh0�eb���X�גr�NgD6s��k�&6 �Y96���w��3dm���=T7uwO��?�zW��3cx��]nKf8C�D��4'���5���/53�sH���,�]��QW�~=����>�Έv_�7 ע�����ry����\�JIF��������aĈ��M�yf�׮��'�>�b/h���\T]Al���JS*M%*+�x��H��f�5d"��,�r鞜�A��9�9��_@��^��X-Ru���K�z��F��y����t,�qmVB_D{ވ�,�֘�8'{��9��a�e:��(�����T�ӪS�`9��l��T�lM[á:��m(�'=A��t,6C���MCS���wRl�z�T}x��s�H�bg��$�r���yEw�z����mU1��g���K�T������q�6;�(�����Q<�-��8�,��٪�̣tm�<&m�c	JX����:���&����<� ���gFKYgF.�A����Zn*g�(����j�g�d�1��j��L�	Jt��9��J'�#���q�W���k�
 �c<G�Z!H����s�ce �4�1O2�Fy���F|�]-.��`���b��w�ƊN�1�EAt�2�^��!����8�:{n�6@�q�s���#:A��d�ܦ{+��{���N�v5٠+W������¬l��xm�u��	Q�Kl;�[�w�b@��C�a�Oh��מ��q}��b &���z+(�O/���-�k֤�tgt��WpQ����.��RY����~@���n�*��xd��:d�so�]�"Hhxg~��*�kn���Hv��T���~����:&���1F9d�[e�^��1vk����˾�E�t�tkٝ�e�ː���)_2j�f%.4�0I/��_S��E$�XyI��]M�x����F�1�v���T<%h=��{�yH��Y�R [$`D�B4CeZ��y[W=ǜ�1�s���ݑ�qr��ө]��{%��^�@�]Di�K̅�)��S��3�.�Щ�g��R-��6����͟_y�R'*9�n!&�
��y�пV��6a���-�;Uv��Y����p�Էe��+�y�J����*#����YT��"��+v�OF��2���vBKH��`��}Ր��=G�*d�fX�½�Ju�>b ��\C���S�~-{}�3s�9b���1�y�E.ylbj�M�`)�`ixՋτ�K'��@gV�����������#mz��C�V6$
�XhF��ޜ��&����On�_u�����<b�h��������錸�����ޔ��[�YS\$ⵕq{.�B�Vi�Z�T�;0qı��#V�Za5��_X%������s�%ۮ^��]d��R��c���ڟ5''`�=8�743y��b�s*tߑ�3P*�0++
1᪅tEJz���	�rk�+-��� "�%�7p��e���=&��Z�Wv�{6k��QQۙ��6�Y�J��
?;�1X�x�
��WV� ]�u1�����Z��5h�r5��5%�T=����zҹ��RXubSx��/f��N^Q;Z�$r�{��DxNg>�T�Q�D;��dg��~.�=��٦��W��T��HPD-�u|ԍ�����׺���;�H	F̄!�nH�����o��
���xv}��u�6�֒t��H��ǹ��u���(�3��0����,�-Wp���1�V��&b�Ҧ;&�GX���s�}N��2�%�j�q0�	1�P=μ���6�*�!a9���+���6��hӴG�j6��Qp������l= 2	@Gf`$}ݕI��n�,����λw�8�.7R����yۺ[rt���c�^sB�RQ��u��������8!��'�D̛�h�Z��_ ��|����
Ѫn�����ϥ��:Ls����l��g�gܙ�obN�Ծ���]�#$ա�]"b���M�����A��ux$u����N�s���尨�[YFY�v�+���Tm�d�6�y�0B��UJL���#9vY�J�&�������/��>�	i���H�ޕ�����j`��)�&�t8�ř&7��n���|'�YPW��b��F�r�P�f�V�6�Li���d<t=$�:������Tգ	Y˄��$q�uazڮ��VuZmi�f��.9�"���%��MA�\���Ӗ�Mj��<z?4 ���Z�S*��"ʹ�y�fb��oX�:�Tׅ3������������Q�|k�d�^C�����6����"������B�P���dr���wM�.������B߸�UO) ��'{g��6w���\	�
�<&��@W/β�>̰�̔�t���9�vFF�C�,�^��PWs6p"	t3�e�EL�1��t��zwa3y�)pY�$�;j��L �)s��D7\�]w��*���u�m�P��jY��J���(}�#�I9���e����ya�&�+"�Cd�"��&��_����/
=�	^��e��x�/���L,�uH�t�4l�Y-ek���
���Sx��^���3�.���_U�W��x]^�M"xy�KD�i{�[�@��N�� k�����xw���|̃ӴB3�{�|�V��0��[0X�TTP>����U�3���G�&���zF�q����A�~hu1�`3���}�fو�82Ow��& �E�Yy���Qm�S@EY��K�����KF>������R�Q(�@�>,�Y�Cq/��m���;}�p�2�v� ���&�M4�}Ps<�(�Ŋ���x�G��x��BNO	[{�i����!��x�Dl.3�C�|5A�uh��c��.�� ~y륐���s���H�[�g>'t�:�o)vT=�l�����������;ќ�`-D��c���^�X�\K�Qá�S��%{�N�	D�$�sݎ���F��<�� �^���Gu�n�j�>��Ʊq�RN�,��Nv������Ή��Է!����`�RѲ`<"�zW�:S7�e5��n��\+�.�ح�Z��\���{��Q`�Oć-Q��]�����-���+M��D7�b�j�_Z�� X7Ku)� ��3S�%���ԭ^��|a<�b�X>�N�Nu��^�n`��f�J�廸�a�%ۻ���UL�2�`MNV���Y=P2au�N��Qyq4��ỺݭOkWB��<xB���CE�,_��b/�̢��jyS�B�''_Z�Mk
����7�M�c3v-u�;�e4d��;
efڶ0�J���s�������O|h?5���x����e�݃��W�X"��]�z��zm��&���vz]{=���L��v�}����F�J���R���Vy��
�5��]�p����%�4��j1�YGT_�]xQ��+�3<����ɴ�����J��:jN���jx��*�z� �۹��޲��k;�L��{��yG٧��mh�R��S`D`*��U1��(�9�onVQn�2=�b�6�
�m�{��3�[�\���٬M.��z-����*Q�u��*Pv(�qͺ�����򁺀Ʉ�R��۔���<7Ǔ\�yƅ�)���p't1;�S�wc�W����d��|sx�=}���8_9�i��R;���/��\	9F�+��F�Sbs$�k����lK��;۹�4��]�!��Au��U��*|��TUlu.�5���<�S���� �X�vj���ް�;��"H��JL���U�!�VN��_�f���V��GU�)��T/D��/w���w]�]�s���n��֨��s��-�(�Y:P�vmP���������	�{��z���NowЪ'!�9@'��U"b�e���)��&X���=���x�����ԡn�'�ŗy��	8/�j��*T$b����U�҇�_�{��ՓL��v2�Q��[�T��L2���Ֆ�r�H�yw��D�r���R���z�,<4����@Uћ;Qý׵�ٹ��]��=٧W�z�f���>iݲ�<9w%MƱ���C<q�x'�Vxo1h=�"�x;���s���՗����e^"xA
<���m2���G%+w�W'RZ7��$��,��y�z� �3}\�Y�+<�ٶ���]CQ�}KY�ַ��2�w`lƝh�rB=;��t��)��uGj�e^r�9�9�X�O&��pY��%I�opwv���Z�U���k����-ͫZ�'�ϟ�<����M�#�!����(f����x?\J���έHx�RO������WԐ	K$v;��r|��!IKhZ�v�u˸f�p�`���
c��4<�ò��oB�t-�L���߳a�4m�&f��,Z���r�|cf�Nwa��j��C[���v��n����s����E���&6 �WO������8���d�:f���w	�K�3\���]sY����SN�?�n�W7�V��&�A��V���e&�l"� �u�v}��[yB�Z3x��Z:Һ������j�h7sޥx�M�$�zz��w��Z��,��x��u�^V�k����P�:����7q�������#�)�3Bu-p��=����6弭Ĭb8(�t�_���ͦe-��Tu�����+���/�����qy�Gݛ�� e5�ްuڣ��]}�#]I�=͑������̹wj�'l��*,�.�Y�z�uqw>7A�\w�n���.��_n.�Fa��;����%,�U�Qֈ�����̫�;L�,VJݘ-id���1�|wބ���2��{�s��w`�.��X.�m� �le�wc{�9�!��L<;���p,����N�w�zx��������w��"��Z�)Q(T��
��*ե!H�aV�Re(�fm���,�N�4#"�L�%L�a
i�5L�CaAF"I�F)�*�:��W3,���fؐa[B�P\���KP�"IM
�� V�;hW4��P4H3�r��T�jdb&e-$*j�Q"�Tb��R8�*��H,2T��NӕI�kMfb�9\T����KB�+bd�"�ٖˡ�&��ҍMS9��R*NQ(�j���dZH�\�,0즈i	)��PE$�AM-�Ι!EGI��+�	$e�]4�JH�D�b��fB�$*Y$���DC)H�9ɥY�!�r$����D�AfI)�4Q,��Ԫ�K5�VAp���X��3��iV�*�eI�Y�*ڦ*AA�i$����ȫ�µd(:B%$y���|=>=��zv��t\(+�0���ζ���.�N˜���BNT"P�|O�Ɍ�_	�R�e�:��Ҷ:���������I�5����8��L�<b�|��1��Ӣ�+����m/
t�1��"���)Eɦ�mggZ�$�����:B.��dE:������ F�&g�z�5W�DSu���b���4�j�؅�`z!n�n�=7R�����b $��#kk��ټ����1�(Σ���(�QZ}P�SÐԖcm��ߣQ�|��4��{)��t:���:���'\9 -����0�V�H�SC8�({�9�c��H�T�:ᴐq{G����#�fj�"'�8�^d%#�1�x��ǫ��t^~�Z�*=�sy.���~��R�ٍf0E6�ߝS2+�d�P�H�H#�M	�0�0����L�ܭa�u��|�$�U��8rՖ`d���:N�����J��Avt��"�w�5�����fv�}�Uh�7��_�+!��z���*d��fX�W�����d-8%�7Ph���[	(sn�NEl�Y�GB��y5W' 1�nX\,Lh����uSzT�u2�<�/]W�z�=���Vrq�5(�����3�6�h|���]D�յ9�(�G��1ʝG�.��4C�V�F�U���Ѿ%J;�f�q�
^^�0�+�Ƣڻ\����
]/;�zn�S���4�h�r�╺�oh�t	e��{��U]�pY��'�b_o��t�V�����1���lG_�wzr5:ɿa��m���E��l�c�9����f%�k¸*6����[�˪|��7�3q�n�eL<>.�.�����n��Ҝ�Y�ZwpU�tf�F,5�G~/�A���|p;����d��;(V�Mc�=��O�NdX*z��8�8�dCuc{<��1q��:P�.��4C�/j��H."x�6>�]�yq��n��!��3"Ru��g���٦��W��A���=8�ʚ�X�V9�}
�S���J�KU=��g���[�!\���d*��yuԍa�֍L�׻�ß�	��7��G��>��M��Рj!j���9�ӃD0��Bf:U�αc��p�mM�]�ۂPdס���/ �Nu.�Pׅ�>T!bB�G;�LbN�Qn�N'��O f3r��o����&�W �<z  ��:̨#��eRg���N$Qݎ׋�� ����ړ�\d��sB��RQ��uρ������N�ǷBuz��=sri't�40����Ü#�W	s`�W��k�#�h3gN�8c����m�re<��-�����t/k��w�U�Ϻ�a�u��]��i�����Y��*I�V�*�!ӹd�oH���y�x�5M�����䱾�����MW���5~�3�P܈n����n��ϐ���q�	�}�O(md8κ�z�ou��Q~�1��@u�Tc|�V�.Q0�XD�S�*U��f;(fl��J�n�k�W��_�I)tr+��א����Lg)�Km���.���7a��v����.��<Ｐ��'��3^t�w��u���Ou��	��*-JdɗC,��te�-�@�vw�Q�m�T7�Q'�3��%�Xu=����t-5���-�:K�CN��e�I<�ÎS�M[� �{f��
�|hB�N�
�GF����zyeiQe�~�UeGq���Č���A�>��N�Y�ÞՊ2��pPϽ�`�Qg�g�z���b�gql(�.e����^�UB.l��AJ�!F��=ۗ�@	���us�;�e�{WN�}�j�?�It'�� &�+"�Cd�b1t�j�CW<,�p�ko5���̓�(���N���L,��;�T���b7e�@2��jy��~��'���\��p��2�4�7�~�:1�t�e�.�P�4�y�]�n��Vy8�������\3z�BSY�ͧ��J�ө�C8-퉥ն;��O��]��ra�9��б��Ģ�B栄��:�َTͮ�}�*m���ݔ�I���V�&�0��_}���}n��K��"&����q�:6/d�O�Y2�b�b�:�r��Ǣ�n��n�� TWv��٨��S)�h�����ӈ���
��.|�OU�j�we�����$�v=Gӥ�o��1��&�g��>�
�c�$�(ā�o�a�G=y�8�lGY^Wn�[���b9�q��ȍf���~$O��nFkէ�$�]�Ʊ��� ��>У뉿:w.�>:���m��R�uh���܊I��Uf�c{��~d�$p�)փqeq{�Ǘuz����y���9��q�i푕�Z�t�#�Nk�b�0lA�Ib��?#q�/���\tn�t�c]�����!f>��1M�0�;���'J �p�=Q,�2���'	Z���J��v�����Cp?ǩǗ���{����E��<Jխ	�-����&��7���]P����Y�O1���j��X1O`AnfVQ�����í{�a�0���!p���	��[(Wq��A���0�Sp޺Φi�ԤXs�\,ՏL	��K9�����;u���ʜ��7��Н(�*i"�����0�gn��ʭ���|�,̸�W�{��U#Sޙu{Y񃐒&��1sų��#��pNwؘMh�9dx��C�F�D�o#'�R����������N��X}��zw�)bdo[/�j����'��WG����Tí�hQTWh��4:�d��-�%8��ݨwYM�#Gl�o6�� �d�T�4s����f�2�B�8wS���}�]l�tL���_��m.�L9GUR���y*k�d¹=�������`u����7~�8��1���×(eD	�uJ�8�{�Q� �i#3���u�=Or4�V�1"9\P9鲄��n��6�+»�P[i��^��ޕz�d��c�\��B�8fh;���T,
�E���g������R�7 �2�N��b6�=맩j����*gY�Q��+�V��(����a�{$<���M����B��n,,���7����|��$����qF[=��pY�����J��<Ԗcn�M��#\P�ܟHQ�[�܋���Ɏ� w&��B*�U��*�U��ڸ�2�q�3v�.ȴg2�6q;ӈ��VF_M3(�D_Ay�@H�����B��s�ܜ��Wy�G�~�2,����i
G�Au��vz�ct���i��t��W-��J���ش�6}5P胫v�/��U�	!uJ��R^�a���Bd���eN#r�˛K��n��]��l6V�glrK�K����'Q������bi��
�1��-s1�)7Pv�����*�!P�7��m����O�~�r_<���/b��P�>�[Hp~rՖr�Vz&���2`]y��׌��b�~���$��:5%ӝF*�]0���Y1�}�ҦK�e��{ ����N��g��������˱Ñ~=�/�vv�Wf������p�6�]�)*���[��ӭ��H��b�^���*;㐝�3_g���^��Ns�8f�8 �B��[���Q�<��j����c�[ꁘ��~�K������z��$/�$���E��M�^������V�S�v�d��3��jn#߄'�U��M�j���'��e&%f�\�c"^>��6�oTe���0��'e_�n��{*zj��ߛм�Fź��ees��5%�d��|U{���m1�XM�� !RYֻo/p_C��@<��u��e��������4�ľ}~R]��u�����@Z��ٟn:R����-���l͎nWo�k�@7_j���ɨ��͸{9f��8�ZO����`��O(X9A}����e��w�d���!�B��;巶��Z]��y���wj�ON��xR�i�}O���u�J�#�5�A4 ]G��G�=�fw����R5�R�W�y�ꀔ-T�ky~z�z���p���4ӧ�Z`g+�Վ-�C�9��T�TII�WPU)Q\�;�'Cw�m�d��9f�]�l=�[��IT
>���>n����/l�־�'<��m�b��`�.2w��ֻ!�ζ�딪1��0�KE *�Va˱s\
k�K���J��mÖ��9�[����r�����$��y)���R�[�qV����횖��V��$�a�k���اL�~YN�؜�f�Wiy����yT	�SS˶��:��6��3P���q�"�y��Ε�ڼ�[�t{`����'"o������D&����
���Lc��.��F�k�&9�@��~�n2w�����v����<��gOW	9O�V�7շi<��voX�k�a�Ǹf�����/˭�ٲ���9cT�<n��6�W���|��ȓ�s�Vg�Q�`Z��
�獖1y�u<y詨1�w��06a�/u���	�q#�ui֫%;�:5��Wk�X���DlWw��f95]�zb�b��*j����k����w;�)u+��^�z<��ʱ���*xo�Ө��vԽ�N5�r7��UzټB�<y�S̼[V3,mϷ��-�)*��3��V4��K����M*2�tk�r?�ޣ������/���j�np��lQ7�
�ϛ/Zk{K��q��@�����j�W���*�ި�=S��p�0���6k#&��9Z�өxg{\:y��*�γ����y��>�P��y�cZ[��we>��Q� �q��\Bi���o��k���v�V�_���VT�3�v��w_����h'蕴So:�އ��{f��C�#�>*/\����+xgf�7���;PR�=�p��������5�v>�o�"��	T��3ݍ�X���r�4��\�5
���`Y���9}�[���EE�7PW�393=���\T72+pv��8��َ����
?p��1��zO_/{kά�+�0� B)����{�'ػ)T]:�5��Y�dU����c�0��C�2I�"�Ym��*�(jZ���Ǘ*y��Gx(0�l;��ӆ��+n�� ��;T�����"*e��Į7��Z�Ι�v^C\5Ap��!@�rW��DG�ݩ}F����7�Ԋ_JT4����F��my;!���=�Dn�Թ�RAEƦ¶q�
��=H�xp���<�5��Cz7�{���FF�Z�Z5��ZL�n5¸�tD������j��r�!N��+[w6d۝]#~���潨]V�'SV�3Pہ�eW���c��3z=l؛��-�Ujp5���yk�׊/j���{x�3nE�b9�oZ9E���[;�k�zYϯ�߬���}Q+W��:��wK�i=i�D����95J���Z�˓�E��^���s�Us�{����}��s��@O�t�{&�b�p�~�|��W�P�u�����K�#+��᩿nf[�����*��mꝼ^oFu��[hN�R�y�X��a����j3��i��Ho��~m>�|�V�Q�� 4��lI4ME;W�n�2�Og\؞�ii�5v͐�9(	�!Y�]x"����#�z��i��λkcp�ÃRrv��.��ܷ=gu�X?)�9�~]�`��ή=}�:�AȦv	�[�U�o4�),�vj:���WW�J�at���/��������Ǒ��0��IJ�i�t�+���e����=<�jyeR��t�3��k:pwޯ@2OA�IK�+�2���R�\4ۈz��ʉ\'�1�1<��m�u
=���"OZd���]G�N���Zyk�ٶ���5�n0^vc�lg[b��2�]�f�]zE{V��5p��d�C�F�-��qd�N6u;�sRc,l&�ל�>D)�	T��6�Q��+���>�[µbc�c�mk����0�ȟE
��;C��ݥ���~j���jOQ��7�+cy:|����CI�l��
��_S��=i��fH�&�ʽTw�,Éevjڅ��j���6�_�^�٘ٮ��FR��2[TD�1��kk�/�Vb�iſr�}����<��x�}O�$���D�qp�#���J5��}C1T���8�qS��WJ{�4A�f&��-�~h�ϲ�]�'ly�Y���<����T��y��HI2�֛:��b�m_iu��9�^�p]��h�}s�q�܏�V,F�8���Ib���Ѱ�g���`ڕ	=�t�Lq�&���0��N�yP~��)�V����ZgL�ǤϦ;�����-�����s�ͭ}A|�Z۳i�c(�F-�Du1�d�����N�����쇈93�3��[�����7�Z��Dl6��^�׽m��e��7��-f�-g2�#�J<��
���b�`�]�1l�y�"���&�a�Y\��cݥ�]E�<]]��l��A������=�EԞoqLc
ȏʺݝ!�c�1U���GZ��̮���{��'����eg��yci�'�U�jU �����r*��n7�߻´����b�^�
�vw� ��n�D��N����ṱ3�����X�+su�&�i�Rʕ�9u���5�ڮ.�KE��V�	�n^e[Pfoe���8��
*)�|l��q8V���;@tM]�A�3�7}N���k郇L�O���6N�bc����3����$�z�3v�x�c2n�����4�S����g��������5�~AlQ�����Z��dID��D;�|��Ɩ� ^����wn u��6��E��t���ދ`;MkX�� /�:	ك�Wu��6[��%�v��)U�׼��\��\{x9�s�h�%��۩9�˖7�_:	W���:��=F75����v���� D�^��Zȹsڕ2�k�q��}������%��Uų��j����[��I��^�c�&ǻ6Q�um"ţrsw�`�[KF�ۚjm���+�X�f��O��G�/���ۛխ�o,�ѹ��n��Ͱ��<q����s����jN���1p��Aι��F�����Td�=�`���M�x,�h_��o{��H��b�^K�o_)9^�:$�s����*Z�R���c�f������Jgjk�ǧt�Y�-�$V�K�U�2�L�0�U�Se���ΠuV�bI����gX-��duv(�G�m���c-��&8���ҋ���cBH�۶��}���'���o�K�U|��v��OAߜל8U}�[/����#��Ӓ�T.�Ћ�k%L�(�xi)z�$�u�!��5�gn�K>/i�3��������]�nCA�z��J�=�n�}X����5����s�L�ߡ�l�2moooHo�l�`�:�/%�l�����޴��\&Ԋ�ZX�k��}�5ɿ�ŷn��އV���y��N�SU{�t�ɽ�c��}N����`SWjg�j�9Xr2�F�^�,�~o�b��s��5å���}|R=�D�fC�l���K�wv�6n���C��s�7�2��R=���o��=���}���%��B������>�e��%���^�.ҩ�F��ؓ�.��Р �4P|> �
C3�����aDĐ�H�.Y!�R��tʂ�2������b�AE�,�rQ"ʑY��R4��2"i�$E��i԰Ȱ�fˑ�l����I��hjI�B�P��r�PP���KD"��%�Z�U(�(��,�W)9Q$��*�2�A3.��Gf�.ZQWT�r�
�5�L�Y[�N�
�r�I3!�I-L��	g���ZҐ���+<��39JVDX"(��#2�at�#9i��)�Z�Qt���E�Ee�*�5�-B5Zb�;��Z�i��\��\���t�A�Q�IF"�&g5�p��l��4*�*)*%Wt�!�2A9T�l(��Y'=ܠ�Ni��=Gx�x�cf9�w���{7rh�����xc�3��V�1%q�tĬ�M}�$Z�A\+|o�4|ѳ�y�ؑ��+�3��A��ڭ^8�N��.w-7�Dk����[S�vҖN��&�>�R#z�����oCΉ(k�Ⱨ�O62%����_'�{��,���O5��׭m%=�^�L���M�Y�s��jK�9����/h�
=�r�5ۛ�W�VN�no���@+���'\%p6Z��{���4����]V���#�g�r둞�Y��79��D����Z�F�|�7�e"{�	���;{9����bg���P��#�#��"n+�"���c�n�F�̴�݅��D��sۇ��E�[f��C�ϰ�w
�ݣr��|�v�Aۼ��\v���ֹ�/��ֻ��T9J���������B�����7X	ໞC��b}��p�j�o�TE�5�q�#�%�z'5F�H��*�~�ƂsT��s܀�V.9I4����8�o"߼�ۮ{�;!��ŗSh��aZ�
�~$Q�,���e/y���#�چՖ�v�u�:�>j���)�Y�ʋ�����T3���鄪kXn�h�i��`Ө�#�n|�h�a�Hyr�����S�'�2�{ *��wc�y�[#A앁qr�=��'��ꪯ���3޳����(Q߁}^�jyv��ru��mG.f�|�tW#��7wGR�m�MԘ�pD�<���m\�57�w�8������K�x{��Ö=���A�y��b�6���tZ�t���D�^�v�`�,�&�iy�C�fi���q8f����\F�7Q�t�]��W�M9�k��{��7�99��p4����jɣLfyq���W�����;L�{��R��r�Wt�32���SojK���&�7g��Hc�SJ���Y�7{�be��j���8ތʃ�0:��ʒ���o��6�\tf��bq�u��B��5n1�γ��`U{b\�zuCW\,�Ȕst�nw/m����4笪��7��-�v�?eXSpy�)W5�״#$�/0ӹ���b�$����x�m>�I������Т��:�3{2�
x��;L����B��N wCn��76�d+Y�/�)���7��ǝ-ͅ��|����ϒ��#����˽��ݲ��/�ޯ|���M���m��]\J߄h�#���ܓ��
U	w�Τ�c��+�t���炻��DG����\��kŧ�/��m�>e��{I��Z�C��w�cΎ�&��[	�R�z���U�>��%-(�{k]�|3��)C�P ]�C=�y'k;p��8K�?fL�=��̀���Q_s�;����f�5�~p����]�b�[�3�.�XE{j?p��1��zBc�����SYY��`�\����اL���@�7i��)B�e�^|�c����`�H�Y��o�b�}dLB�'�H�@�_[��E��%h�ob��q%�)�V,�{i�>���`�n5�Y�r�}}�����3����}e�H��̿N7�q��t��I��E��6�kW:能�ۄ(��+����&�e����Q�� fuz^a�z7���[����'�[���	�x�]�X�3n���#v�ٺ�2/�@�F�o��qڝE�'~*^�!�Ldh�k�'�˃3�p"�7�����*^[�<��d������ֺ�T�3�,9X��"��!J��r�D0�aōrM 9]@���_N��D\�����;y�^�nɐq���Q���t;k��i#%,��`���k:��G�@�h5ʤ���_}�،G��o��w7}�����r��3��f����є���:Q���[��$:�;Iy�x����oTe�ʎc2�Uρި�9K$��&Vn�^���|�l7�a�l(��)���x�ѝge�킯^M'��7F�=-��V)�]
ӓ�^��-�ZB��.��i�ľ{~7��{VȦ��޶I��?\z�����ָeӑ��=[���i����;��7ppmbe�\�;� |}F��?�:�1�I-4�<�h5��� �Ҕݞ�z�o���-o���邠�$�iI\b�s<�ݷB�tp�������X��x{��Ψ�leC�f
}��������1����O��&�^,nZV�jY�
�M�e��!q	d
��Ծ�����n��)q+9�x6�1��k��2�;�gVD�F}��B�wC�R�D��˯l����xvJy�&k^��q�{�� +���5yY7sO��b���5�����,^�ּ��PZ:8���F�EoT�z�b�9��p���ӹ'�`���z�5�\��ܐN�	.�&���/��_���1d��rT���m|RsQ6�j��|��O��4�vˍv@6+��]�3m���Y���ϕ/�U��o���{W���Sƚ�֜"t(�!���;~7p�إ��~�y/�2�_�uC-�5�/4᜷�v���j��>ca�+sT"��:�N�u�L}P3�gV������b�/�[��K��Cs^>�3�����DV���Y7;�����.� �f���{���Ile���;�<�.޷7�oV]��C2'=8ح�0y=G�Es2z�[��ø=Qє���mIo$��k+�����zձr*�,�;�<��<���;漹��%�^�y��i�s%$UP�}�5�
\G4�V����,9�<qUI�l�����\Ҙ�7��z��~i>�I��{���/���(��GH��|��>��ܮ�[l��S��Ȏ���
��X51ֻ�tY�E,���&a��T�
ԯ@1��>�s�m&r�P@,�����1��9�v�;�����>��7�m�1>TJy�9<9��îN��$�ޘ��o�Pl�R�$�;����x
�_}�UU������;�����z��i*�C���J��F�� ���*����z�����T�i��K��>�ؽr�HW��(���H=o-[����x�&;tT�f@Y؟gD9i\3�����r�-Y)������]핒f}��g�:Z��x,U��$�ahN�-{pƫ0�^�����ߌV\8u�x��ʼ4\_���Ʒ������3Y�0CZVض��+g��ˍW�!/��	�Z��Dps��I�v}x_����!��:��`��Ϩ�L��k�
r���C��趯���=��+���<�{Ǌ�q��z���}V�9ΌN��f��Q��׷�룻�fyb�w��O���P�VDDhe�u�MqX��k#]{s��ͪ��7�5��9+q���*pZ��^�[Q%`ˎ��;*^��u���ޡo��-A�z�����bA��3EݥU�381�=�N�9V�'Zn�ۥK��gC�7�f��p��u�
�}��z�i��g�wY{%�U� B���u������	FƢ�-�ݘ�U��7��v�����aEQ�4��wc��諭����5=�%7F�>�m��>F�d��\@���Z*�2�=�N{��s���d�z�ߋභ��*�z�\�N�j5�n��VV^�l�Yͻ妶	����W�6�*γ���e���)�<�*ˮ�P�wи��G`*���lS��_�O�'��c��U 6|Ts��Љuz�\����98�]��ɼzZ���4��5P(ug��B���{A=��r���@M��]R��S��Z�c�^��,��F2/�Շ��V1�?
=�������d"�yU{<�x5�.xNfzZ�<WLor^9���~�fQ
{�H`��T\�*�{F0kc�6�G|�����i3TA�l�4�X؄��z3(�1ҕE�'�7�󻕄��ҽq����_N���o�'��o��gp�1JH�xu�6:���5V���_)m�᠇Zw0��1��c ���7����>(�[s���ycr���Z\�W=�<Ē�����x�YN_>�(;��J�WHa�KQ�&J�XFЃ���\�^��oZ�x&μ�y�qEmnɻ��_UUtO��P��R��_=�o����5&&�]�Y|�U�j���,; �b+����e�����ٗ9�j�V�.�W	:��ᚆ�j�Nثp)�U����6�L{C1ץfZ��y����j^�bpˮ�su���<Ɨ�ڕE�Ь��wj�p�.�_9�U�7;�~����r��^J��ǣ.Nm-U��%�g���u�7Q�ʂ�>�h�D��tisz7mV��m�&S�w�62%���oC[�Ts"9��7�'a���x﯉�M���D�7��+��(�	�k���]�m��;^�9�nR��1�kOf�\�^=a��T놴�Hu��M�����[���yt��䴧�����"�>������2�)*V5��z�����ӽ�!�:w!�
y�bW�]P(t�0:`�>W%.����Җ�R�t:�r�U,)�lS.��CW�kS�u��yc%KF��5Ǿ;m�dG/�JT��^��5���C��@f8�6����LM]
!n�3r�YQ��ʋ��k��!��{uے�WΔ�w�n#�tW6dް���Z/��o�M��d����頻j��N�w��j=o�"���|o�LV���ojM�w
����k�v��0J�;͋}��ί[c)�2�S��0"Z <�b���b���o�i�x�1�j-&/;�3�c5�2���	3�����osO?b���3��΀��|r��̾�a\�1�A�(ࣩ���3�~^��؞���o�j�K��So�t�Qi0�.5��S�0a��Ԩ3�gH�\�]C�艈�6`���"'��ޢ�S��S�B���	�mNe5�c��ǗFs�s1��6|/�՞cǏ�b�Nm��)ڧ��Wf�V$�?s�یn��L��=��voX��Փ7�������W��/\�U��v�q�dF���U��3(��޵:Ԕ��i��>��x듨e�v��i�u����n�m��e��=�� ��_�����-�!�<�i�t(*:<�p�3�~�@E��=�q�zmWq{*��8$����k��f0G��]5�O�V��e���i�yĈ�G֖�(]�^"�ͮHBJ�6h/���ܡ-�M.=B�t	<}�+uC�ܱ��g�^�{ު�����5oИ������>�u�2R�� �r�t]y�E������Va��Z�zp{����;,)��uBV6Z�lt=���b��L���ܼB���ϫ=���a{���g�9�yW��:�-Z�^[�(�UKˍ��g�5�Ɏyp�>��I��މ~���BO�]�a&إ�wk9w(�	r��Bm���������-�IP�x��W� ��(֠ɓ�1�k�2뻜s��>��/��ֻ��S��O�/"�����L�4�˟�i�W�kk2Ψ��n���չ��E[ckT����u�᪔Z�-�����@�s�����q��M+e�uNU�Q��:���V�S!�ɜr��5O 0x=��h%k����W����f��,�gsHfg4r�(ޤ9�q��yJ��Է�߳����]���O[6�֊����5|���4Joru��v��+��,�Aw"Bxo,;���n�OX�#�i��s� �['G��s�eX%�̎:scMt"S������d^^�77��e'O�^Q�@��R� N���H��g�t�ۡA�T:��jS8+�%�S���¾��<�M4��Ad�M�ڣΥa�	vѠM��&!@귷o:��aq��u<��|��>�z�$����u,�X%��j6\V�@oH����i�t&bU�q,��u c0�j�i�%���M��SԈa��Z���o/l�'�0����!�I��l�5mD'iP�L��vÇcñ��,�`��-�JڝM!.dk;r��n�d�tˌ���^d�_`� ]'(��Z�̸����t�;���g&�gr��p�T6�.F�þ�K��;��&��,j'&g3�ŷ%�]��yy�c��A�`^�^v�i�vǾ�s�Բf��3��a�=�@�Zn7�,^�(�j���==h� ��^�e8��c}sS�oN#�`�˒`�7�����ia�x3��lb;�o,��¹j����#!�q������� fX5Ri���r=�9��Z����m9&�m�hm�R��k*J��B�@���T����8�6��daU�2Ժ3؛�Q����0{&��j�z��Y���_t���kI�ln�:�9��EƤ�C����xb�R��S���F3q��(��/k��R�*���֧lr�t�p��2l3�#ٲ�u�-��nh+.���׀��m6n��S�㗕6^8j��ɻ�"��(n�jA�p�.�'0��_eA�`��z��7vV�D��;�	����
���C������!�w��N���݆�ɹ`q���n���ɲ�;l���Lٛ�����C�򃔤���s��v$e	Z.L�Y��jpK^�T�]}2��l�)�WW[��Nf��zK�-�O�t/^O2'��վW|�y�/�8�pݺ
����j�(-uǰ���@>]�ˢA��L�r�ʰ������\o�av������(�:�h$!(�H�)ɞ��K`�6�<ΆKԹ�u���O\�؜���P�X��N(�PE�L�W��n����F�LK_��|�*��{��b2�Iֺ�4��4Fb|�yon��{�<;-�N :E�)���P�
�W�k�}s���a_SI���F�\��ؐ]��חRY�X0|��\n�(;Ѕ�����5B���O[��f�,�\� .h�+:J�2n��t5Ӫۧ7!S��j&��v� 1VȊ�JK�'��{[��{�s�֭j��.�Q�jF12R��Is:�ޓ�;bAZNl�P{2�e9�Q\Q�������U7c^\ժ��l�Rd0΋��@�#i�������Z���K�yZ��c��$�N!��d�v45�P�wl�2��|����i�ӮF��]���s��z�z����xZ˥A�U����$���\�2��d�DL�1J�г�^xy�M�g.Y���,�$�Z`�d"��r����r��
���^�h��@ѥ&�
j[�b�3��-J�*�Yӈwt���+2�S,���P��P���&V�N��N��.b��t�J��W5�ٛ.�*�"@�ti("��Y%��b��WI�k��N�h��6���c��\�+��DZgs8S����'M�S����+�&�
�$R1w+�u'�E�a�P��h�B�БD�V�q=Рs��t�(�Z��;��BL,�䜡ή{�!L��T�;����É2.E�F�sI=�� �3�X���+�aYʪ
4}��||��O�\n�-�nt�[Y�w���"A~����m��%�e�N�K1��g]�u	K��ӳ#�\�B�<{v^�$���}��g݉-�o�H٥�����Qi0i��)���"c��kj��*6�^u�'���l�����յ���u��2�-�Q	�TF�7Z�m���EN։�I���1���y���N����^Zq���Or�N�)��}�oxs;��O,���[�=MJϴ�z��Z�C^��Qx���/#��2{.Ϳ��1і��5k#=o���r^|I�i�J5��Z�<0߫��蟡l�~�[:'eU�ǃ5�CC�:���UW�n�e&%��R|��6�î͸犽�gj"���1ǌj�@3�����ŵ���P'+�5�OYm����5���=(���D"�%�Ԟv�簽7d.s�ͽ|��=M<�i���3)$��Y�m�2`��$�z躔�Ҕ��ֻ鉪>Vǡ؞���U�����*�=��74簙�mĎ���]��ҝ�Ӭ���9${�mPN�Eo;u�\}r�a�+X�`����J��h^�3�S��N�]R�XNpۉwq�u`�̃����=Ћmw,Nw�)�b�a��}@�L��Z5�Q�U��ԕ2f���E�C�]����C��(>��)\����j��nT��_i�Zb���ݠ�8�x�\7�*-��Q�"���1PR�^�����:X�7��%��Y$�ǩ�z�gpT&�*30��y&ڰ'�]��s-�q*�B�{�xV,N w*��2��f����3�;�d�y���~Q��AY�e���T{zul$'�\M����0��:�`�n5�Y��ûջp�{yj�:�W��Їs�W�7�}��A�����ڏzrN��ӆjp5�qc���99��ӑ��D�z,�^���ڲ^��'~����{W�m��.����ku�Q�gRb�蛮>�y�u���۳o����c2:W�u���.;S���� u�f+��$�r��oZ��C���v��|3* ���*��G�wU(���_]�ǭF��8���L#͂�kmo[[�vr����w��ǜDR�G�O9��Ѩq,*�]�?xp�g�sЩ��e孭�s����`�/��s�#���=`�P���8l�P��%��D�+e$Ȍb�gdׂ��el�����f+��da���jI�"�*�NC	H1���\i����w����l`�V������|�t)��T�zN�끎:��1Msb�[}j�5�]�gr�G	�!�`j�*o��V�
u%uD넯L�@��,��O��,,��f�#L�CLn�gr��p�ʪ@h�q �#�"v�W�(��������Un�̻�\1ڰ���~o{D�l
= �e��'.C�I�V׬.K/��jio���^���Z�)D���ࢠ)��BHE��4d��g��'�iJfĪq��j��q��63����r�����&0t�Ī��ԫj��uf� ��y����n���Գ��
����f
�A����i�9�J���/z_�W=�����旙|���;f��J{x�%��a�1Sc�^_���k��]�{��>A�}F�L7���/^.ʛ��RL+�F�|=��c!Wxj�"�o��/�z���O?=ʻe�2-�Z~C�.ɞ���~~�p\��W<��	*��knPR%���Om?S��;�Ͷ��g�wP,���]v�0�bVmup����)(593J�f����M��� }��%�}K�ϋc_OS���[޺8r��w�YI���tTr��q����Ǩ�W�n1�S1���cb�r e�z^eN-}�0n�3���u��K���v�����߱8f��3���ٽc����[xT����^��k�Ӕ�ی�U����y~I���G>��t�%�mc���G��yҶfS�0k��$�}�&��~*[���u��;͔��h�ƹ�˛�7�9k�|լt��X�W���l���8:6���n;��eE�M+V���O�>�?T��ӝ�j�6)f�h��ol�!�k��Y5�-�&���k�u.���,�b]����c�yv��ys1!@>p:x�m>�I����P�@l���˭@*c-���Z�,r�:��F�;�ۇ�����y>[~4�
>�|�T�����Z��AmK���tZ)��"5
Sı�^|3��Z=�n��Y�a�wb���W��R��~n�$pIH��=l��c������5��c�r`i���Az;�r#�K�0,�u8VF�s�# ��',8u��SF�k4��*�w>��\���!���-�d�<-���P��S��+w���  r��6�2�#n���'>U�+�OЛ�Չ�2����[����;	���TQ�P��f+�9Hs��(��:����f1�OI���{����+�(؜�q�)��P附F��75˷�n{/{��Nf��8wx��1_X����o�L�wd"��!� ���'�Ș���y�[Tyn�S��þ�&���O��4�4ۍvN�"y���c����ٖ]�)�*����y�PŚ�r�8f�ہ��Uk�|��a�*�4��fG\���b���EON[��L��=^��d��`:AMq%�\ſ8+O{���!x9ȻF�����b+vT�v`>̡�b3K>�;ݦ�3�ձ��f��*᫃Su'���&�SB�>���Ѷ	�$�v���޶��Fds�'g���e��z����D�|�n)�_�|�ޱ&���N�˨�=ۍM�Pu���y�S	�gj^�����
���v�`��:t�$��+�q��%v(p�t���p����1%ZS[��n$��N�c��p����Φ� �mE�֮ĭ�`�ĩ��*d�&�dᢣ2�.򎴳z�{�w�q�7a�i�o���w״rc0k��ie]���ڼ�ͬSܺ�s�%(X��ا��m=N�ќ�ܳ����eF�'�H	~7����^���so.��އ����	�:Ehz]%<�	
W����K��t]D���a���Fu2�����)�Z^m�]-T
7�d��V�j��z�>'����NÊC����ز�t��3��}�_!r����T���QwV�����#��Ըy��Iy�Ա���͇L�!Lt�P40�)fCۍ)ͫ:[Kun�j	+y�G�n���T5Λ|��!}H��7�j&�g+�w���W��������ܚ��T��I�i1P��vF������,�@K�ʃ�֩�����y�>�v�u6�2�e��{�/%^�#{Ҧ�CkLB�#G;P�5n�7���?wzc=utJ�'k��z�d&��Mjyv��A��[AJ�U���o:t�zԧ�k��Y��e�)@�Ҏ+A��_�.n�7�rťgC�2�q2��zeҬ�kv���-1��;P��G���_��dgAʨ\�V^|=ݵ�/2�\�~���b9S�W���#^��^]��a���]���Lj��=0b�i�b�2���w'�^���@��nㇰ��UgƸT�Z�(u|�Y�k$`P�g��ٌ�z��݅��(�\�<�ȗ���{y�vr��f0+è1
\�c��g�G=Aw?��uH�]p1D�&)�l��*�ۆ�U��U�v�d�v�	r��X;���;%>��	^��������6P��kU��m�v×�|�vʪP_Q�*y��k|&I����%V)ejp��y�B�^w��}t�{I����P��(��{�w=������\k���wv]wc� ��e�a��=j-�R��G\w�IP|9��50cL���vgf�Mv���:�~T�i��knCc:�-��T�
{���E��=.x0�S={y5�J^�r��j��;�B�|2=7b��F�!���:/ v��Ԩ��l����o��O��.L��]o��ВkmY����E>��X<�{�׵�����W~��,[�����"�w��8�t�2�����Q��!��j�9�+ �fD'1oJ��~��ED��^�Fs�RҶsSyca66��EU�m��jn̻�<�n1�'�us�����6�!���8�R����P�} �����L�gk��-ryvV�y:��O�k3{�!�َ��r9�v��pN�Htg?�>RN�[�_�(Do��U����\{K��6I�|��E��n1�*#]1`N\����v^����J�z���X՛Tv���}~I��'׭��	�k�Z���잧~b���מ��x��#꬈�Nѷ��^Ӧ���Z�t:��LB�5X*3`�f�͇�kj�|'�aS-L�]�'���j�Ɵ-�o\7Y�f׶���u�E��d<�^�vfu���M��h���ԇ�X �3���5u��?6�n�Σ���Ruz%�קz��i1O��L���`��j_��V=�pMғ.Y�������>Ε4���\�|��}A�q֋�-[q�ao�g)tfejyz{k z��'��RMG�����d����va�xc������mh�:}ҏPK%aX�:���&���wy<���Ʒƃ�H�B�Z�3��ON��O����X���V&U�^�{e�X�7������P%�}N5�����������l�U�r�\��A������^�SR�O`.����';��|�C��>Yƒ�C�z�b�	5�v�9��x˨Z��pPkk]:)iE;�KZ��:���T>��v�V�L.��X����t�BZ(o5�gV'���g�HU���w]t�ۛ����ki变��l���o�G�n��w,�Ջ���M���y��q����C�gȍ�{���sS˴��u',j����ǝ��I�~�|2�>f�|�/]��*P��6`#)-���&�JPcV;v֬םѩK��j�����}F�L��k�&#]1��u�HzP�}�g����og�m��R���6l����v�3M�I�(�������n�J�q�.�ٔ3�l�V���>��Q���$k�G뱊,ŒܒgZ������U۱nT}DJ50Ǵq@�^S��m�3���MЊnk�I���>y�M9�|���*`q���v�D��W�a�[� �q��VG��q�@��4�>��j����g����v{o5:��w���p�����+)��+}R�gF9k��f�p����j������1X�r*�fq�v.l��*z�%po��"��p�,��^���n�Cs��n��F�$9Ǚn��0L8w�	�bVx��B��zv���"vXNs���|���̥X�Q�0�6���
�]�^���60��
�^Ynť��%#���p1�P�5����|��,�ٞp�z˛���l�pQ�z$�T��OuW6�ކ���=u6�����63�Eb������и�zG�>���$CfO0�ĘP\�]��gO64W]�l>���KbX_y`t-�^��;�1<�2��j>G�=ţI(����}��[cG�����h�`����|��{����eH�4食��A�C�*���՛p^�c��=<��⇉�>3�K��M<��S���heLj���<�9�GP�_9�m`��ħsh>.Hh���U��������Fɡd<[!�P�qf	-f�k �ŧ9[t�+�m*���D�(�{���('��83`V_T��t.E��O/5aeśƗb�|���R��f��)�LT��Ė��d�|n09����K�}^i���>;X\�0�N�ލ����,��ASC"-B�wo��}��B�T�
�CK� Y����g^o˘��u0�k����u5(��w�>5�(4
W���&v�Źw��u:�#AEݕ�Ә�ך�[;��#\��wa2�ɳ{�Z��j����F�����u��'[u9
��ī�%Z1Ӿ��ש1���Ω�R4����bO��)vvm�C�+�Eʯ���l��Vy�z"�j�z�
���9�]/�؈9a[ɩ���'B'zc8e���/��9ʯ���KR�ѯj���=W�T��%����[7I��\���T�+���d�pK�8L��i������N�|:�V����>����l��K��NYN��Bgav.�����X>�Ao^WX��|�NCr]Ԝ�r�Bs��ȿ�aL� ��ݥ"����`F���`Xu����{��!�o�J�*�m3���r����J*�K��c)����$ŮԔ���V�a��r�OzWEf���+�.D�:%��aۧ���澗{	����x��N�t,h죤g m�N���s��J��[�����lqU�jib-���6s���iD��ĕ��7k���ٽ����m5�OQ9Ӕ�\��/ ����-��wUv�N��m�u�RR��a���b���Rs�;!������6�;������%��ѭ���r��|��u&���x�oa�Fn���h#���5bkKf�<���rV߻Gz��KS��gc����2�&,u�蜸(������Ӱeśu|���0��N��7�墨b�=چ�N�c:�-��&�u��[���{Ը'[�(r�*��Y9��e;cN2�)�G(��W�����5=��;f�凨�pLB�oT�X�ޮi)�n��Q�t��t\�g��pnV�I̕�����怵�*M0R���:��J&�ӛkkGZT�_E��l��S�7k.���/O���khA��Dw�\��yp5ݛ���<��� ��i�:�D��D��+-ш�P����'�zu^��b��k��"
r໷6�P�w6�'g�A4��x�L]k9�y*�ԉP�Iim�������[ՙ��u����2e��M� Ϯ,��K���5&	�;]����yc+�/S-^3ziBuE�nJ�/N�ُF+A�cj�����l�����[�+(E+j�F���=�?�>�{�p2�++��R�CKB)J�XF��*��ݛ�����(B�A��
L�i��NpH�ts�2���8ED����E9:�K\�<�t:�*�Y�9Q���� U"#JtB���-<�b�U&�#5
��h�\�
�Mֺ��E4���q%����Q\L�+�!Z�B�l�
�-E�jӅ+Xm�j�c��k*�YµT�PRuZ���U�����U��BQ�nwq1�#��GpwAΞ���3:sB�N�Y$ܓ�\�:�1I+K��]�(��YjrK��\�
�NB�����E�vG�" �p� ���((IdPPG*��
�,��\��-\*���N�EU��ժ[Gp/<4@�A
d�YΒ\��MD�D(���.��L��V�IΝ3!2sJ�\*��k�w[�Uq�>�yw
=3��srp�	�Z��4�b�=��l)i���Fz�63B6�\;/M����ƿ9A�n�\�R]�3��c�׾I�l楐��M�y�(qҖT� U֦;��av���۞�=��:����}s�Ƴ��<�ŗ}Y��5�!7�S�yW��=�j&�&�3y��B}F�L&�`��e㯆D�kf2���!KF�����G�a~[���Ӥ����L�b�yy�S�S���:'c��&�S��k�&#����guq:��F��
��
��O:�Z��}�q��5n�W�e:�a���}��W�KU��X�{q:�ѫ6(�׍:���.��=k#]r^�9��	���G^����>����:����:�Dv8�i�S͌����ڇٵG��\7ޢj�`�X�_��i���G�5uz\�D���_&5�lީ�ǅ�p`y=[�a�/��g]S��g�`�)�zuBW�z��)b�v�w�������
-�ol��� �[AƄ�_������v�mdq�2[+��oB�-Sw�Gm�f(1�l�=r�!6�)K����
����ozu��I��%c��[;'=���@�֙��չ'7h¥hG:��f���*wL��w3���\��9��g�P�l������w�>��?�G8
"������ћ�����9��״�}~5�Q�r�/=�����P��+
��I���	~��0�x�k�-�R���Gy��P��j�^ӛʝ�{��;PH4{�9�ʟMy�ꆱ��c:����BQٚ��fT#���]��Ⱥ7��Nv���G^�r�-+�3�����֓}�jy�Ֆ�qp���(j|4[7���]�Zn�sj���Ξ�.qEؙ���G�����N�3ŝ�y�0����W��>@��'�T^�#���s(�r���dLB���H<�;��s�������
a�l-"��e���ԚO���k�@S�H�j>�P�2EQ5���[Z�K����՝��'9؜3m��O*����F���/W�Ձa`�e���҂P�f��R�hH<l�ޭ9<�h7��M�*,��=�װq
��ա�v��g;דv�L����k� b�;`f	oSRk���k +����yE�v�M�j��=Y���.E���5l�r��^�nP�I��ٰ\x�)�w7��"��(��Y�����N�i�^8��Zȍt:��SQ�ORX�̵��y�s���w��M��+_j��cNʗ��֫�@�f���
+ۏ�ٓ������d��v|#g2Jc�(�HL]B=L�ydT����f�c�.~��ޅ��-���uZ}.xꆀ:�Ҫ�r���O2�Z�0LSPO��覚/�9�(γ��d�u<jܪ�����&�bK!v�J����l<�Ci���}~5��zPެ拽V̮aK����-�nԖ��+�:�������5�C΄�ۃMU5uH��G)&��a�m�0tT�`wmj��ZuJy~kZ�|3�U�vl�B��s��U�G�$'��E�T�Ǧy�7�ҕ�&u�7�I(ޘ��ߪ-���(ϑ
c���`�KED\�"-O��x%kV�Ug�REj��@��f��r��Hn[y0vhh�r��(�������<�{s����A�H�e<u�D���y/�_��1��V�����O5��c�1oǶ��I�p�L ���������	�'{���`2t��������}��N�E�\6N�X��Z�ј��wn,I2����k��
�&�)�3�D.��h��l��Ù�3�7��{­b~ʡ��������=t&R���}�j�^/�x۳}]6��L��6�V�=���y>�^���q��F� ��y�&n��K��M�<��P�ݘq���յ���9:5i�5��
$ˮ��W�q"��Sv��p�o/������'k^e?.Y�^�䰒I	�e�*�}�{d��o:�>��S݆��f���C1W��T��.#�8D8A�B�=[�t�+��b7��>�6��Em>��_q���79��ih�8S��j�>q��nq0�eO62^>��|�ϻ��Y:'_���ybG�_��X��Ц\K�Q'c��8�	�����k+���/B�:��> W
��c�Z����v�L��:�+�.����<c���~c"��F�:�;��+&��n���̨�2�������OdɊ�#+�tOAk�q7/1C�Y��U�F�ɯ��B��K��U�1��o�M��x�qN��@���9����i�x�Y��s;:u�a.N���^)r�L��V�I1iEǶU�K�õ�p�u6��a�nE���Y��p_�z9=�;C�'��w��5�����g6��8�`vhu�o{l��
��*��UX$|�G�$CD�i�v���{�:>QE4�7�F�p�=���KE�> �$�F���[�E'��nvVvcq�
�7��r���}���le9E ����۩�-��{��;{�wX	�^d�^�ݷ
ZV�jLe�M�e��B��P���g�Of��J�@����Ӈ�2��4���3�+���xK��s�vT��xp{V<��vP�ٹѪ��N����Q��hʮ&�,�TN���7&��1��<��Ds����`�OV�B�?h�ݷ�;���k��]����3\3M��
�]��L[P2���TN-}�qព�mO�ٺ)���O���qn�o����'պQ��5Y��Ky}9���C̩S�����[YS�:�{�-<;{q�6O{ E���jfb^�R]��.����Gm,O�V�ׅ:S<�?o��$g��z�$D�0cTf���2�!�}��[��C�^+G�.�nE��~�q��=3�{\	��Z¯j�c�K+1�Ҡ�-MR3)v��r�q���S�i8ֳ]���%�p���sRϒ,�ԡ4�f�U��m�fTR�79Ry�����Ɲ�S͌��}~n�oϷ�K=�g��LL���K��M�̣�03gP��b��I���������'F��z�Qw�ڵ{GS�;c�ys[*KҺ�@��}�^3�$��J��5�-��5r����m�����o�<s���O���O$�>��H=l>YoCYqS�I����:|��ʡ>�Pǹe����0��K"��3󓐹}��X����m���Gw�o�������<�I��Ql˕�Hzߣ*��}=_cX֯>��ʈr��X�u}�aUk���8[~̓���j�Y؟g9i_��[�����K]-Wd�f�8��l��x������f�us�.7��HG�&��\�f(�g��Ԙ̈́�ه2�zpV��y=����nm�#��6 �of���j�q�E�f`�@7���N
m�{�[��37��b������h�5v�+Lr��3Cc�[8_u�F�	�o�����Jwz�`:��h6�Ör!`��h|��N�{��U��
gl���`$S׼i7���x,�R��C`q�}��`��ɜ�c�@������r��ƥ�2�[��NK��P+�А+�*��T8}S'�3��rP�cB�������j��հ�c��|t]o�h^F�>-UK⪴5�
iP*�'EVP�6�b,]����hE뫓ϐ�_d����9�v6��L,���t�f�uM{Un�ّ����P��w�`�w@�H՜��dv��S׷L��,Ve0��/��\-0ge�mw�FS�A�X�C{ί)inMW�G>�x����c4�N\1��M�5,�Us�o�uM/��w�~{�ss�W���'~ ������]8��#���b=v���9Es��%u��L�t�Hgw�xu6�Y烐\�|R�Dr�S�WSf�r�/^�Z5� :e-���y�B��^��n�nV�LFt5J2��SNm�Jp�
�%�F��q�G��3�:;�jbs+�s�d���9EF=�\|#�����n�|~���rp�z���;�Ǽ�/�l�4{Z��Z`��ld��J�ޯ7w����;9.�ejhnp�ݶ�-��@�K�Q�=��ؤ��8�%�f��e������˓/��ڵY���(�����*t��<\�|T���ʓ��.u%�l3��4�b��u7N��a��}?)0�%�%�)tV���RM�Ø*m��G)�3���e�Gw�nON
"P�dƸ���Kz�D�>Ua����Ҿ/t:�F�_��`��%�<n��[�p8���FN���O>�i@|�2^$�����ą��θ�}��fbr����7y�׹�5HL�D���YDf��(��)�t%0�Ih٩l�� �r�ĎdG�:��{�x_9�ҧ����HR�yl�z�
fJ ���@+��r �������J�^#]E��csUMbl+��o-9	zf�3�+z��!�1]U�*D�P��1�����KͻLEś�Z.ѳ��� ^�߆L.���K[z2+]}��7�����1�O�����ܷT�t�5
w���R;�V�����O�/p�i�3t(���[�)��&��oI}���T�7�mۗت,��t&�2�A�b�q��ɧ�Y�#.6Y;^��ݨwY_#~����m��㛹��3��С��*D�{��F:�TdꃺpT����E%�:{��z�:!^��u�]ۖ/����p����p[�U������Qx��jN�/��5�.mȦ7�J+�j��;Y)�j�\��^�f�ӌ*��Yk�\(~:?QUԞ���	�����jXm1ܽ~�P*��QİQ�f�w��<3�e7��1f7�! �a�Y�	�V�'�@B��$i��/F�W�\�`���5���9o�yY�-B��	���S��<2�S`4�R3�'*Rf��5)�Ux�җvs
��6e���ĹK�C �Bܸ��!p��2�u�����JJ9�/Q���-H���8A��g��[�^\}�s*� l�b���$��W]AW�K,B�}���h��j��Y�cCq�u��%�X���u�UZ-�*x+%�,���8~U⌶V,��@[�hR�J�.��uu��rh���	���j��w�t��3%�<�����d�$7_j��Y
�P�s�}�ewoYr�&*i����+�Uw��;F2P0uF}�����3NdT ���1��7�-�٤�{e�^���+Π�_1�g
l=<�fU�$Q�S����!�k�+�]��(��$���C�+�^8�!��a:[����'/jPB�F �=�B���~T���tĴ�1���`T�������7T�(s,��AVݩ֨ZO^�sŰN�'
5Dõ{��˷��S� عњtU��ܝ���sx�x�ʕ�6W!i��֩&%G;�)If�t�� ��aT�g�N�6���gYX.0V�]�^m�l��c$����8�>+�=a*��.�M{��Sp{b�zK��C�⺪4`��%��S�h�x��S�w�K`�5|>��*�P�q�9�A\�;cr9�ͦ:��)��Kt�iǧ�:G��SZR��[9ɧ�Q3��qntSxf��� �+ҝ�������=�[��xa�����*�E�.�Z�a���2��y3�X(��K
f�l�Ͼ�6�l�c�nlj�寉�ξW��h/6
{F�\����ӨmUL9~z5",}+2�,�r��@��^�Ұb�Bs/���.>4�I/�K��#l��I�(�5y~޴�Yo��cvV*T{�����A_���1���'v�c�W�O�X����%�.����_(CܞT�ek�΢�-<M��3��oxj�O�-�����T��ؖ��G��roD˷E>zO'L�^};،��#�\�]�K�o�9\*eHۈ�d�5WƢ�� ����$��޻��M���q!%�L��J�k` r��?�����n�+�l���ٖ�N|���۫^Wr���o��wNZ�S Ag�xL=
��z`��`og8�f@�����s�`�n��9�'^Ż%�XUPa��/A4{�N9�ؾ�!:�c8[��BS?<=����(>z�,t8��QE8�&�%���x�q�Ͳ��{r\���c_3җ�gzdu!]Zz똥�p'h��wQoJd�G�������z��y�<�̜6��knwH�i�g���^�V�>Ժ�i��z�t2��!1��9,�^�����l-Q�)G%�N�K���޾'�)��Z�C����Ebc/��%7_r딎�[�Sl�u���Q��ugU�Z�-h<����s�X�Γ�0hW]�p>���S.fvS�y�p�s�����d�L� `��TA����:(S�=7
#��izb3n`�٧.��q]`
�󍺄kq���'��}�.-�)z��*�=�q�X�r� ���{���H�W�&tu=�+XWe)�:�ahQ�)	�xf���b��t�8oa��㎯#��xܞ���}�K��<����]���[]׶Ԇ<���c��lѨN��ؖ�ã �5ؕM�p����z�Fv�W)IP�lu�1sW�z�4��sѭ*��w)����p�Nz���3��ɣl���ТVG�
*���rՐ�o+
Za���iøm��Sڅ�g��n�����)2��A��1��S���;�e-y�*Ոi3�����z��=��
}��y�ɻ;���o3ڦ0m��5�7�j�m����έ���������M��/��>Yz���;V���Dߏ����@j�{{V���?XPu5����)I�0�v^I�j��v?�
ة!XR�EH��/(�˘ȃ��g�O0�7U��D����4sƻvm#� =������,��䎩�c_���{\}��%yd$���s�k*:��%=�|	��/o��K.�(�Ğ�:�|Vp�@�����LWmA}�н�n��Öe'g��l�X�:��FMnE]R>Fl����c�����-�[���8}&���J���8m�M��m�d��g/n6���Ecj<,xNr����kך�����s�Wn�~�IM�؝�赪�����`��ک�Z�ޮ똪B��u��5ˬ>@B��HZ�)��x��y���⫺���M̏��-��L��M�B�$��{s����[�Q�)���S�{��\Bу���5��t(���{�Q*6�}�]�9��)�pvnJg�ee�ԏ7�Q��E��˵��qf�N�4���;6����ěvv�U�Ur^�w�+H+�n�aة��+����2.-�<������b`����3O�ᾃo,=�[<#ų��C�j�[�{��V�YEy�
G�M{e2�nek��ٛ{d���WV)C���]�XWZ�˲Q�]6u�d��Ѵ;��sb��d���8�	�|0b9�
I��%=ؕ�\@�ey,u��S�yIe���C�FkS(���
]�dȋV�+E9���, ue'
EN���V$�W�ܦX�.\��E�YId%g)'u�����I�9Rz�*�-+T�sM+��ӂrT.�n�mU��@�#$ȡ3 �U�trf�慐�Ζ����kLT3g
��M\�GuSwn����HB��L�$ÅW%Yr�YY�/�*�B
.��B�Sj�҈�Q�9��=�YQ"�V�Q�r&���jЬIs
(�
�J�:����B#�ܪ���N����EA0�s'9�QjY��L(s�̜�$�M-Nr�F��y�Y\ԣ�0��I��;=ݔܝ�/T�&�x���(.��bVQIU�hkQ�УDۛ/5�$������a�G�@�63ٴ�3ݵ��Z8�A7:X��<_z�ں>\׷<4�\�B*�wa5�
0����x�k���d��r'xZ�3�{�s��k���I3OǍ-̺E�l6�K�3l��`���Q����DK�y _MI8�c�t�w:��5��0���	���P�Jy�B�{}GU���iS�@}�,㩹��7��<�����Ƽ���D �ž�,����3�-Z3�W�ˡ{%�=�M�%���E䪑�zh䀗���N�X%��"u'���������cֲF��=�ldLW׀��ܐ�1k�(R@6�F:��:�L�SD���e\!�pzH/��9JZ=s�8u���>@���Y�;rC��	�s�e1]Jy%<�[!)��[9�w�2`G�xD)�t[�xZ�]�ˬ�7�s[y�ҧ����ǖ�+(�@�0PP̼��i\�Ǒ���eݬ�L^$k�?�rO�*���8�JӢ�W[����W����UhkT
�	�m1U��G�[ъ6�\�p��L���1�b߽<g@��l�T׵V�푕��ͅKꃙ�Q��6fA��1��HZ��V=?UL�Љ��3	�	�0�Օ��u��.� �ߝ�U�P���&�#5{#j�$�&�7F�����V����T	�B^��v�L�06�ȝ�f^JIc}�c`�X�VTj��o*��h��ض��$ ]�wo���1@"v��Dɝ�!�����g�F���Oz����,ϭ��-�j�ʓ�Ǳ�SO�LL���i�E���e���7A2��C�^?*�u�Zn*e�J᥎;V(̼j���޹;�W�A�Ɠ��_l[2n�,����$���Js/z�B��1+�F��.��m�v�`��,l&rء�� �T�C�*�l��^���p5� :9�E��YU)=A�Oi�b	��N�p���sl��8Yc�((u��L��"�H�zbѓ�o&�IB7Nv�~lΚD��2���X��T�9�YD�i&i�����Τ�[-�����ɪ��js�k]m6����� p���^2��"@	t�먟���.?�F�/}
�jj��ǫ=�����֧��r����p8�\M���{��p�����jWh�W��Yǰ&��6���%p�Jy�
kJC�yL�� 1~� nGċ��\M�B�n�}�Z�}\�5�a[a��͋��Q*�А>Q������/鿌�9�Z7��m�k�71B�m���3D���J�#_q���L��[)��P+�B�@Z1�w>1$�J��FV=T<F@��;A��ب'"�-�h�rܗ�3<89.�~��5��wFE����\�����ζ&K�X�7�|��*Ǆ�Ŗ�^Ll��4.�\���[x� g:5ֶ#����Jn�>��^+,u�ĭ{�xCD�:m�Y��L���~)WK�G�ףcxK�4ٞ�W�'E1�!��P��@(&|]<���:�:k��0֛(4d��OT@ɇ�'�1Q-m���_q�ަ:᫼d'�܋ڲW�t���'1�1N�b~�EAwU[�櫘q;�g�c����T�
���z���;e�L��-̭�MN�u�g�[6%.��V�E�a]̋��΀p/�ݘ}Y_"kQ�j�t[!�UY�sxУ�бAB���'!a-�b�|�����
�ɾ,8K�}J�x��y���r��Oukrץ&gELG8_�Bg��i���&~H�rϝ�:.�tN�l�1:��;��啟o��&XW꟨踩���r�\iv�R3�'*Rf��7߽S��ʏDT�kY�$�]a�#s)� ;�A{�q�LB�M:e�7�
i�b����I|���Z�mn��wtA�lB�f�|f��B�F��Ğ�,tT�F⻶��;n�~?��廌h?�{��#�`q+�$��e�����.�\Tk�3��$�a���we���ۙ���Y'//4&d޽[d�0]�6{�[޴����Shm���yVi�C����^�B�A��ɴգg{���;�vʎ����Z��v}�v@f<Ȇ�zY/���Od�q�i(�J�4sO������ɜ}}��g��_3������6�Z$)�T�JU,�`#l�C��ޱ�.i�����I	�y�w�eޙ��O�n�q�����7A^�)���%u4R�]�hvd�`��ZT)�I&!��M��<n��e��^T��uM+��,��we�����c8V�}0���Fm1�F��R�=t�mY����՘��}2Qrc�:��)��qI����s����dm��_�����M�{G.���E�	���N���`�E��i��3��`v����R��r����8�ꝝ�Z�s�@��4� �	�9��y*�Kt6\H|G�1���NV������!"�s��VM���e��l��]��i�T;���`i�b�;��[ �|F�
6���fҭ��j��Vr��nY!I�B�{WM�Ī��K��ja����뚈���q�ʹ��l�p�S����T�>BuM7)�=+@њ
�{F�_�ĬJh�8������p�܌�[f��;dO~JS?b3��;:O�gG�S�tT�J/�K��b6���+N2T���a�9��*��L7mnSe�1�|gҎ�h��=�/ǩ��Z�I�|�,n/w�ui�o��/�	�t+�9co�E�2�aN���7��p�@Ƕ�3�s�ԡ��.q
�aZ�I-4�m4rm�=��tQ�U�2�*A�W.�α���G%dܿ����s�+�S����ۃ0���Y5���,�L
����d]Yf�e�ɹ��>�;����jcSϚ-,�z�g\Ɗj�apў�w_U#q\�ݹ;�KU.kkivZ��]t�v��\�=2��cq��toҩ���*F߮Y'�zJ�ѕP�����,0���+;y�wcb�Ù��USf}R�Z��-�+�I��ފ�~�"�'��������i�՗yk9���[jb5G=�T� ���<ih��:/�`!��X�0� �Ց��*�݊�g�{i��8~�j�$})��q���5:��S�4�W>=����X����h{h��l�dZ�i��ҙ!��9�߹ÿyv׆�#��1���W>��)F��r �*^���E�|;�R�o>����`�P���u���TQ���Kp��;Vm� ���b�I�Q�#�# R�w��M��!��=��!�J�D����W��/�^U��v[x%�岸�(�)�
�	N���㻪�~E8�O�����:��*7��f�έ?��7��������X�ս�?k�っ���+�b�z����
�<�	v�����
�YJ�ҭkǥ��ԠZ�N���G�C�#��նh-MM��ͺz��47b:��m�Qb�9e��lk&U��H�.)��;�q=��!�-��h��i��j�Y�R社C�hU.�ukvdZ�"Ν�����x~�\�p/���R�趜[I��6N����7�*�CaM
���V*Mֿ~?������	��;����j�$��^Ѐ���2�g��4�=O�76��ګt���j��x�������w�bL[�'΍EM8�o.j�(nN�0��;��e}��R�A���J���S���2�4�N�p�*u~nScx�˩���Y;��0���T9ɝ4�؍o�}���{y��;�r�Ϣ��>��*y�2�-l��u�g�{h_�N#��&Խ��5�'�K|�s����uu&��S<*LrE���g-��� �T�C��WSf�,���^�Yɍ�A���g[*� %4F���T�z�T�0uD��>�N)d�d���ʍ2��w�4��,��塞?{��7nH=^3�E�*Wǭeo��X�������X�Աu0��,�`��	C���ۉ�R��F��*��$�J]7���'�o^�'��k*�-6�#���[M@Y=a��Դ�c��X�qȗv�����Gjf]>s�]���}�M����C�٪���B���i4\7��,9�N�/��;�0���ҾY�0���*j��:J6� T�/�v��S��Ò̫}ٯ^��c�`��	�K��� ��l�=�ʎ�y� t�C�P�\�i�8��x��x�l�r�����y�z�y]��nT��5SE)]|��2W�Jy�J�/�@1>n�L������J黂>S}%�v�P��c8,�R�°��bU-�FhHc(��R�w�QHA �����:(�b���j�|�(���f�Y	�@x�e<�OJᯭ��|��[)� �@+�g�L����U�:*ڋ&�2����L"u>ͼ��%����ރ����P�*���3b�yw��.��f3�gR���� 6Y��<+--m�s��Q�Lu�WxP�6�dH���o;����=�1	(N�iǧ��s'a��p�i�07B���=B�.[	��%�b̳�a���Mj���2�^.��V�E�O]w0�^� d���)�d��}��+m@Wo��l�r��1	��v	�e?A�X0�v;ͦ�[��'$�����^|HSG��I\P�۬n��RB�O�73��#�/� ��v#L��@��a!��6�3�!�s�Й<�f~���Y�ط��rgn�G��O����r�j#��췖%f�M����(!3�;Y���%��� [G��t�~�x�r�
�;��x�p�*޷�=KpSAvU"����8�=%@⾫��7���˧�b@̥vԦ�9��Jl6�������
/�����#�m/t��#�i�7]2�c�N�@���Îq��'��5yH��ꦀ�i6*�M�s%��Xʀg�S?#u΃/=���o�� ����Bݖ��|����2�(r��U�;����9�^�]���7�PUC<u�9�rIe}��I�Ӣkk�E���E֋��~�=@��$�3��T3��P��0X��������bWTЅ4���Ld��~F1��Qq�gʈ��a��V) |�~�,ċ�V��c_+�E�3�N��2�1/�!d2L�Uwe�v��������)�=[��#���_`Op|���9��>��p7���,n�:��Z�;"}m��Q�D�;�z���>S1�#*3>�_Ω�H�c垁�A�qʹ�E�Oz��i[~�n}���
w�Z�y���el��L�O06�!�S<m�aH�M�튶���R�]i&�D����Ôk���A�֭������	�U��lw���ĳt6\C��L��V	_��f]I���Cݥ\��=��*�]�~��+�u�Y����kaŊ78��7����7v.�Pe����:�9��5oN.���^���-�r����K�Y>�Z��Z[b��:WN�s'V1f�q/ M=�T�Rn���Tp{JهrWk�:/���D�.e)�TU�Է�R�*n�^\���FjE��9*N��|�s'���-Ί[8mfJIɲ��u?K_����1�F#��8��n�%Uh�aR�S5��\r��A���״�r��b���_g=�u·&`a:l�f�GA�0o�6
״i�"��bSN�q�USE�b�Q�%�]�������߿.?���g�����e��gC����1��}�]��Nj��]���!)�}�jm®���|�cռ*�0gN�0����ɭ7R��@�`��hOa�6��.�{d�y�mu(��!��SϚ-�,�zι����l8釕�R=��'f����{�wn�Q�
�
�˲��h=�&7�taO:|拝y��E�x��4�lBɎG�y���v��1��4�,��l&���ꕁh+i��Ra>��}g�7q�&�y����p35�S`�_zg ��P䟜�;֮�7$�<S4�[.���k`!�ֺ��o:�h�Z�����hfGe�}?)/�lj~�	޼��V�$�5:���N�|��h��S�vjo���-}��UX�nM��8ghp�uh_�Aޥu�wM�w�N,jd��[����QJ��ym& �{UZ�S�^WWE�C{��Uo'�D�-�H�S�Ի;�3�C�'wGgNE�'�y��mj��W'z�u����V�ܶt�Y�,nr��X/����F�e7L�ƙ��bTd�}$\���t+�����^E�(��&VZ:D�q�(ͤ���Oh�J�hP���Kpvre�4��;"�v�_5v�t����]Oum�Ό���yf�>=1H�tp	8� &)N����d�2��ٸ=$N�mg��V�uZ���:��Ȃ7�RmT�
f\^[8���)�
Д�����;��-��LV�}7X!R�r����ߓ?AS��?)ǚi��6��A�^<��f`sY���I)w��!�Y����j���w�����İ����U1�1��z��:+Ǫ鍷U��
iP$�໧䧍�י�џJ��@=n���fl��,�P2a�Z���E�'\OoK<��}�e��^Z��������q��TK�Y6����b�6c�����ѳq�'�!�b�/w�Wn�e�;�j[Ԟ�J�B�C�r�|�l�g���a���3�Cغ�Z��pWLw˹�׻��3�ļ�� �M�*y�9�1t�Bn�,����S�z�s�(mG�A����L�����6­��q�ѷ�*��Q�ڋ�U�^���m�
�@fS.i����uD��q����q`�&��;Pr��k�&C�q<�WZ`�D�E=�^�5��f�N��0����PQ��*���Ǘ�-�+W��¾����Ɗ}��ʰ�ӫ^��g��`�Q�.�:R]����	bT��#/Qw=̄�iղ
,��̈́��Zdv�:6U&�vK*$���,v��s�00��՝/�@'s�K������v��~|�,�z)�N�:d�G��;������8�;����͆TB�,��㧃�ܮ!�^��p8N��r�a�F���G^7h��ʡ�]q/��sb�y���۫�s��W.�L`bZ�6�\u�Q���]��6�hr}7�K6�e?��ū����G�]݇,����t�>+�.9(w
G�zy���|��s��=��Y�l������͏�����e7t6��V�b��w�0�[�^ӱP[ =x�E�f;��hИ�E��>����^%Й���0;�������YW.!�G\̾�%ȹ�ɑ\iޒx��B-3y�7n��j73���]֥�L$
 �z���u����3u�W1��훼��պ]��8_6!�w=
�J��.X��U�M(����E�ӛ�M]�p��4Dc6M���ǐ�Q�R��?�]�uTφ�"^��ٝK���z�
�>������"E��5WYػ&���j�Jp7�Q��h��
i�f?uJ��F��rJ�3B��yrȧ�k[sP�X[x��r��.�<n=�|%�G(��sqn2�㥩K)b�.�q�`e�Q!2³ks���ΔQ�o
��Rk�J�|����sM[,�řA*�h	���t)�/4�H>��+s:��u�����0ܓ�	&˫��S@|�
{��`!ό�0Q���Ԋ�Q|�9���-��,�S]BD�%۷����Xⴔ���:�r��%7Z�0+���7hTb��������OPp��+�g]J����z"Ee7,k�=��H�.�a����``=`���yn�s�����\�C�,�=��cƖ���3�+�N������E&�l�^������X7i���f��W}�:.���]���C��Š�h�!*�J)w�f�`ֲ��2��7:�ŋ[ڵ��ɳ�nw%�4��5�;W,��2��G�3��� �����v�h�r 4������S)Х֚�|8SlM�3,7̇�L�I�45h��c9k_Fpb�	L}9�ɛ��z����	F����z��nX��<�W�ܥU�Y>!� 5�ý8Cr�n�U���J]��[��O]�pf���lV�~��9�������1�eJ�ͤ��9�����aw	�hB�7R,���Z5����n�3���t��{��.��u��{��ĥ|op9]�b 0E E1�R�FNt�T]QR-�B�IOs�*�(������lI:�x9��L�7EԨ֑Mȸb2��8��!�l$��&�iΝ�t��E$ETa�\��	�K"�H$��<�3�s9�E�ݖ�N��ӊ`f�Tj�(�g-��N��(稚�2�RQ�K*�J�q:K8�O]۸�.��*�T�W"�b	G<���H��y&l�R��rT]�Թ��s �Ē���P8jEwY�WDw�Dz�*�����]����G<�۫7ws�s��7Ul���6Q�5ܺ܇<!=��7q��r<��g���*���r�!)�m�����㣇"��LL���$n�y��Qb�ܜ����(�5�Gs"���z�8H���"�s���)t���rtq�A���$�aS�L�v�M\�R2�uw@�r'rv���"��$�Ȥ�n�	�ի���k\@�y¼�<]��s�2�)����d��%�w��ã�R���S��݃&uH�i&Jl��J7Ҧ�ژ�<�L�	���y��Al�b�)�k��,��fa��i�x'D�ޛ��9�ܒQ?�g�������:����a�)N)�HA`�d���t�aAq�4����|��3��o���3l��2���$�2��~E��T�4�K=�n�K_W�@ќ������υ�	}6����6�Q�Z�P��.J5�~$�X
D��R��b~މeW����~���t�~bG�\�Fy���+~Tt��P8yӨv.K4���3��\L���gDqf��Zit��zʂ+�:��0���k](�\7)��-}$oG�LM9�� s�nE�� ]l����5��|G�-Wp>��{��j:ј�%Q!z�6q��]��)�����"���apC��t��m�����g�(R�yl�z�
J ��
���ժ3캜r/F-�}4�Yؖʼ�6�5	zf�3�*��'E1�!�]3�*�CAos�"5��w>��� /�M��Ɩ�T r��1���koD럴ڍ�c�S	��J>�qV�y#�A�u�cQ���8�z$G��E���yCc�b���4�����:�<��=G����F�R�w��K�s�N����E�s�~�m��SC\��Mu�sT�V��^����\Q�.�4*�� ����i���飑�v��q粲�����ǧ\��҇Q� \|�E�ﲤ�OĪ����W��N=��f����w���zc��U���U'׽����̭�*]7��Ɗb��_�eH��d��|y^�7��>�|�t��[�w�뙺�ZN����7�n���be��_�԰�c�z���srZjbS��-k\o]pE&�V%�tc�M����pY��]'�@c4�ߊ��Q���
��5�ļ�F�qb�gG��:v�e��3�]O�t]K�򜁐]��N)��ԷCGN *��Lu�;�W�*l�J���g\Ɗj�a�\F���\#L9D��/.O$׹T`<�xr�gH?X#�_�7!�O�>�C�f���G}e�z����T���E�}���n��/����W�5��e;IM�-xHe�l�[EQu�H��z�Ƒd�Pfͫ��?�s�t�j
\90n���f�v�V5���m���\F|���uL;�6J�_3��H*A7t���#@�oS������r9Mu4R�]��F!�1����֕���*7��la�^��	���:P�0��k��/L�w�����p��7ő�X��N��`� m����vw>���"��
"�;������v�)�ub�W}�+��Φ��@�A�´n+Lu�-K�_���.Lk�g��d#�r@U-�Æ�f����_��@�J#�?I�p7���,n�:��T�d:��1�Φ˺ۜ.�s��������J��~��w��26�f�L7c���hdR3�n1�W����nsv���w������/Θ�T�Q�,������n����_A�1�������n7A�2t�[S���̵ېkʵ�������L�G�~�Ȁ�4
]�4����d>#�QcpE��W�{���[x�	�ACj�6��<�S�y#5"ʇu�'}
���׵\�(�J��'GT+�>ߪމΤ��ʯ�s?A���N���\Z<����yp����
�u����N� 5��U�f�����\�
:#�����1���|����h�͂�^ѦV�bV��u����n]]c�2*�ay����&��/_����gn&~� l�w9GEԪ�N���F�;�j��>�m���/2��6/�8M=8�[%4�����W��c7exC���b�kL� |��jb��K����M�
�+��!�r���T�:ٍO>hJ�����q~%+�xA�(9�����`�<��?|^����Z�s�C@!�Ȯ������ї��7�{�	��f�n	l��/�!�二�Vob��r�U�&<}}f���3�-7��<k���%�(���h]�RYJ��nΟ맡��_i��M�;6�5����ֈ��;w�����gpw7��-Kmǡ�j~ZSt�p��ۢ�M�}r���ևâ��~�MB��x��ք�:��?�I��e�&5΁	�\�C�F4�&p�{	�bڡX�[�e��*���1����g���������v]�b	��� ���4�Lx��k� t[-���(�������8�M��c��"�s<�� �2���|f��e��w]�ϯ�B������o.p{���������f�iY��;�a���B�Td�o���Ҿs��Y�Σ�iv�Ţ�$�:��I�Fm�J{@�����R��Y��B"ux��_WQg�4:�Y�geYG�d�k��,��lTغ��阔h��S�+fB1��)�zeJ�'�!Du�!�='~�]�y�6WK6�-[�dT�*8��ަ(S./-�zTIO8V���g���S�/�ҔRk0��П�|�����&��zpT�V���l���PtS1���5P,����IK����Gz�2��޽Y��g���#��WO㒇\���Zt\V�����>7����O�1?s1=S#>�'�}ˤ�h��Q��p�O�Ojn"����o��+��"�{���:�jA'^����M��WRʅi���J�7���m���n��'[ΰ���|��ę���5����rf_$�r�k3�ݾy�ˤ�z��:i�lkwh�y�-�$�R�ѝ��яˠ"���*nF��;B�d�WkC�������c����N�:<�j�(��cӯr��kĥ�A��{�k��DP��ܧ���\-��[I�L���̜����ƀ��M����V#I�ʬB1��@�)���]ԅ�s*FZ�N�0��lq�7�]�g��.�?E}��T�D�����7dy�*�F.�M��=�/T��wݿWl����WI�ʈ���B�ᓰ���	��`R�Dr*d��*�l�MX��{"��Su$��n�����U� �h�t�k������:e��f:���>�N+�$ ���!*�OuV���6!o3���A��Y�i��`@�3�*�ƕ�g���7�9�n����n�FQ�}��r�Q�[l"�cOP8O� I^|���2r�����{����e��������D�ݴ���*ǶGeغF~ϩ��:�K($f�T��5i'��̾ؼ��Ȁ�GpY����a]M�W_:�rSϠU�!���x�
�������/�U��XZY4ͼ"-yj��Çn�� T#��M)5}�sE��/�r�%�E���n`���x���͵�t��9�A_�h�` Ǜ.��EZ;�<�^�j|9�5�t#G�H\��A�.�����8W���?��[z5��q���۬�#��1��zJ��W�܍$};���)��q-���Q*�̢3BA�pR�w�r�M	ތۜp�F��ܡ�l�.�� ͚����D��Rt��ô)�	��#ԠRP�(s�py|/B��R�U}�J�8��L��ǧL�/� u`�s�K�ٞ�V��tS1�!Ж���O&�,�+��E���n�?)1��-�\)��.���"���ɇ�'�1Q-m��V�Z*)�&��P4�k̾��[ʵUo�|�T=5�.�)���6�ǧ��s5��%^t	%����H�˄G�I�9�ܲG�`��f�׽����̭�T�qM8���d�׺�a��`�d�B'��N�u�
��L1K*��b��`�W�i81
��e��[i�a��;������O@��j�ȞﻨʛjN���82�6ĳ��p;�����=��+�� !Cr�D��lw�}79����X�P��w�M����/���
F=z*]���`+���i��������fQ���9��qF�U�ٷ�l���g�R�,e@3ŋ����rf����>���>�ғ��v��J�/ �J���{.�+�d����tLSx�,��*EK�;k6�1&6�:�a���3��'=��z��dԟ�4hY�^$�Z��hP9�ݸ�z�O�>�J!`��[��Nܝk���<V���Y��ض��3��h���d��֪y�[��Q2� l��(H�LW�ے�1�#�}��X�7�UL���ӷ[���k�C-l�[LUZ�~�%�Y%'{�N}
+��Gp�7����X]1gL/���"4�����)����U�F1��C�ֺC���5�C�+�*��%}�>D� �#������	��>�I]M�UwQ�hH��Y������۲(�4���� �(!^����n����,n�9�oZ�;}m��
�Yv�~y�>s�ײ�`���/��)�T�iL�@[t�O�.�x��s	�&�ѱʍE��n-�6�� �g'��d��1 m�Kc<��-��x��L�`�ݗ��Ƶ���ؼZ�l�R[<漸�t�WUC�"e �N���[�S0㛠���!΍l��R����o2�v���7re�9��!!�lٴ�E1唞����VT��JS��ri�\Î��=�4Nd�¾�X]��Di����n�������)z+r����U��
�u���m���d���%�m9�\3:���sB�n;`=��v�	Aҥg:T����t��7��v�[�%���F�&F'O;{q%����3��<���߯�\^�.o3.�Jt@d�k�eL��z2^p��5��c��K����Soh+��f�F.�`������?�D��F9�i�O���t��(U�e~���O�R�[;��W��U���N���f�Bȋ������O�#���2��:�X��m�Ε��}��V=�`�MNwW8M*qJ%�5�uo�6]�`�E��pfT@��b�kOj�>;d���4���6�.�i�Jw�ZTP���ʓ��)�SϚ�����.������Qk�)-;��*��mF�ku&�1� 7�j�+ݑp�Ss�e1������ʑѶ�Do��H�}Gl��8�_� >X^�ʚDw�Y�L�q}R�[-���[LWE�2��:�koX��{����ˮ�{��d�r�'��?!��uL'���SI3Ox��~]��n(�x��ip�����L��v߄R��P@����|f��[,k�ߊ��O<��Y�+~���\l�	��[�ܯ�w�'J��냿L���f���!ǐ'`=�F3�'�O�R��Ȱ<��I��J4^�Fm�J{@�J�hP�%�Y� 4�O�1����~����|�ж���ˡ���iw�����D�3���7W��[l�C����͵����1GC�p`�%>��4w\�b'��5ڭu:�q�Ӯ�^k�f�8G����Ԣ���<C��%�,��Ǯ�0�k^��ܯN�b��B�4�)w?�� ,yW���^�-_1(�{e
x�[�
Q��R���Q�d�ΣzG�;j䞱�u*���� �
E�B|��b�^[+�R�I)�	<'w��-�Z���pz����B�:�V����(Q�hߊ�/�E\VR����/�����ze � m�o�1���2%�����qw2j:c��0��>��V�Z����O��5yp��λ�\\0Dm�𞸀N�[ɥ@��	�mx���a�7~%T�j�mhw?i�t�q=��U��~��8��Y�K̽��[���U[��*V�_��}PuD����ǧ5Q-�|�ܧ���$�[�5k�nV�n=�L)N0��͞����#)��)�L����g�x���0�b �2�;G�����*��L�J����� ���Q�1t�n�,��m��i��^�["�ǐS�#~�ߪ�1���:�U\n�T/K���M��L�bF��'� s9�6J��M4��/��b�x]_"O:����\=m/�R� |�_�a���g�5k��E@Y}��2b���`]�TcG��`��rn����e:���Xɍ�WL����Njt�A������^JAS�)�'���oVH7B�T_^RT����A�֜W.�p���@"�8�Sf;�x���]����.�ƟRVڣ�K�h�����_�d}n��q؄{�qnH=^2�������s�.4�
a���L�v�`<&�h���u%��l�6��L������B?P,"Bh�մe���m��ݚ���KB��z��
�trLˤ`�kS�0W��cL� �� |��r�T
4)��]�f��}�+k����s-�)����R���d�����iH}�S%�]�9VE�L�����Fr�#r�v~*H���p1ţ�([8W���%Q"�Df��2��qv��0��Q{[�}(����g��}6��I��5?���D��HU�*h��
_���*6�j���*ֻdP;��W�`�Ȗ~�g~%�ՠS�d�E���3�鱑.{�Bq��}��]���Њ�����	���#��@jb����L��̶4�*�Ϟ��°����sZ��*�m�XՋ�U���˪���qUP��T���%�<�b�ʐk��U�}:�O{>����\���s���ؚL�
��ZcoR}z�^��{�3+F�u���O]yR3b B�������*��Sϧ2���`���f��ܯI�[����[|)�Ӣ�Ǝ�byXe5�#������X�V���#�L��r�G��i�deu�&V�Yn ������l�T�weC;5B���\���ڨT�t6��<�,�r�̕ŧ��� R�`�-B�)���U���T������i-���3W6���w��|��� �wo;��Z�]]ԛ���M�\%h�O�˴`)ј7{��
����\�;�9��W���v�v��B� �AW����\�H��S�i=j�,z�l��h����\�MXE�X/&t�39geDCEVjQ�5
q(�<��Ұ�b�6�4kkk��fb��9	���o��ȥ�T�ׯ"�f�d[1]�3�^��Vv
���K�I��-�C��+�g���3��}&:@��ҼsX�-�/hY.��%�RGd��j��).*ՙ8��"2٫�
�=�x�Q����ujK3�@���wwzn{`yG�d��lh�f�mm��q�����=Ԡ�q�rPS����!�'LU��'9����̕�	�t�ZZ�^�f�m�>)��Y�v�h�ʃOϲ� 1HVE��7�� �]��C���{��w�G��t�@����}������Ͳ�և�1���	�����ڸ�����U��;��^f����
���&Д�T�k���8�R��[z��^�ַ�����Ȉ@��X�;ePڕ�����OR�y�Q��e�ZN�������۶����(�2�͹�I��|qͷ���Z�RG�M�X��ýuD�{x�����-���ۖ���5X�؇7!�>mԼH��N����^��V˹���@ׅSO�??��Wh/D����2��gn<y���Sc��˚o(�>xx�U:�.P��Z�V��D�y����7Wk��E�K�P-�	b�(1ԳeB�������ӷ���X�@m˨���&�D���H�s
�&�t�8��ڕ�Q˙Q�F�)�V&F]�4.�K:���]M�	]�J-4rMe׷7�0�2��l(��u��w���l��Fk`)3�>�*=�A�*�`ҮW��7[�S|V\��Pˣ7����9o��u�
��|��sLGٯg�.�]�V����5
�M�է�͡�u�ĠgZ}ڊG=�[�^Bk:<�Tܳe���һ�W�.b��EK}�%���W�k2��_ϻ�@<�'�Sߛ�|͛�om.�[��J�,�0{~p-�E����~��G�p�NX�O���t�?1�Ahd�T�h5,�T�\f��ᗟX��e,<o:��;yJ�Ά��L0��t溭j���N���q�f�ł�jT����Z1��=�}�uށQ�w�FG<7�11Jjݞ��|��6e�����n�x�("��\�6s2Z�V�ǯ�Y��˾��u��D`�bV�]Ȋ�����ʒ���8��w$���7�K;�㞡���9�*s]=�y��/D�OD�5̽U�r�rq��J�]p��#&����Rm$̼�iQ����3&j�9��B�=�Q�]L�$��-MJ����(�2��qª��/ZQQ�p�)�njF��G�*F��2�n{�EPN�l���rp,��β��PH�C�"牕rۭKH����+���	���Q=E���㐝�6TyEʯD� p�B��D��$�P`EJN��*�wn��N���]�fi�*�fy��\%D�\Gal��T!Ե(=meGJ��"�]�MԝN�4�wnj�.Wԛ��-'8���rW<

�W��@E�UG.t�D#�繚��2�L�FI^F8y˅�F�sզy�UzR2�2:��]�=�3(�PE�wB�/�������=�i�R�i#p��הˣυM��n3�Y+]�@�G:�wp�����}9�iʹ{]2��N�� �M�F���\�`�HS�eM7+�4��l*��'��2�be��[i�a�`�j3�C&J�rc��s����^�N0e�F9�M��9�Xdy�F�g��/�Ī�Х�c4��ς�wXԎ&)So_���U����^#_�(:$�t�x�G~KH?H&$����N0
\.Rx*R~5�٩M����1��A�L ����b-j�V�G�v�m��G$:i���Jp��ԗĠ���T�q:;nc�P �b�
"�vO�ˡ<�s{tnn�E�LF
a�cuuӷ1Jm���$2��d:�b��є�p�-Kr�߸+x��w3����@᭝��57]SB�'i���cQ��m���E3Z���ݱM�F:�ܞχ9�l�^r JH����-��%�Ai+������1�ӔsOmd`�a;��/�B�F��tJ&!���"�'�"b[�8���9�u�C^��[UA#os���d�3��#p
)S�2�<��D��^}���D�z{�?\�zE5;�A�[��o����+��z��̺=�!�֐m��n�uup;EE�{3����l;[�a�`��}�(�����M��%��k-rl�]YϾ���Rm1Hn��NQy��<�kUz��b�w�<�<㮳L�q�G �1a;���d_C3x�~Ǖk�>�Ԝ�� YDb �:��y�-��<Cr�<m������y^�'f�̬:���M*4�V�N�����tL B���lw�*�Kt7�C(���7֘	hܞ���?�\�]cr9�ͦ:(��Ol���VT��J~O���X���1֠
.$��/�+y���� :Yź�^�&s`:��pʺn�UW*���,��\�S����L55��zn�.����S>F9��O���t��Z��2̦�l��E��ɾ��.�ݼфr���K����+�L�	��>F9����^���=ګa��.��n�\����M
yZq�*q�Ji�muoʨ���fW���C�B���!:�߳S��v˄�s�q����B�O*N/ҥ!�jy�E��ϝQ7��~��^�H˭u9���b��4ӳ$F�wG��e�\nȷ�����)��E}h|;!��cI�̢P�����ȍ�;�PGr��� �>����cR!p�4�pE3a5LoϪV[������Տo����Z����� �1��9��W�>j�{ݍ�ʹ�W.���������s\7{'^in��4p�ci��z�/yW�7{w�oUokD��#^:��\�3��|��쨕9���9�;^�Y��S���ʽiȢ��`�on�(4��ݫ3;zZ%6�f��]<�Ῡ[�@�*��	=Q2���wS-��-]n��~i��Gԥi�G���q����(݅�!��]Lv�Ei�S��`�XAw�~�B+D��C��j�O���FvY�/)�v���Txg�tMiSQ1�=@"y��t�C���8�t�h�&�l�ץ��u갪�׵(�{Q�E���-)a�B��D'���qFUNQ���Qb��.���dSJ���s-������(�tp	8� "��*Tй�d�%m�>���]:�x	��+�Ѹ�-��+���11��z�
�Jy´%;���k���Z�����#��^iJ�ҙ0"}�@בP��/�ENJ��E�]��4�T�w��q�hM�J�׵𻀀�Q�},�x�s&���9(u��p;�Zt]k��^{z��	��ȋ]�v6�{�4�X�i�7.���ؓJ�h&q��(V�b,h��a�d�n��:�\��a���V>|�Ƙ\�R]^�ӧ�#+m��T��9�i�S-�zzf7s+2�����暜��X�j��I��^�Ԓ�̫�8ebv3r�Z��-Fh�	Ppf_Ve�X��jj�����5�Y��|� %�r�H�^��U���K����\z�>��Ec��ǀ��TV���t��ډ��
vo�I��::,�r+q��:����$�rjq�ݴ��k���eV!�N�o���]��M�sk�hmLoc�Q ��\o], ����8�s8*b
��K��_dy�*)�b�MΎ���U����P�9�phܞ���L� ��Q��,�a���6(G �\�)�f�4�UP:�=�e��3�&���Sf�%�_!�xu�$���%����.�˷ߦ����踫շW4�1�F
�&�#A�l�AC�ʍ2�a�xm��T`8���~E��T�.�q� fWf|��m���/L��L�ԗ�e��(�-�Hø�(ב����7�;�ɚ���Ib����G�'uͯ��]�y�E����[#����,o5��(ɖ4�P|Xϓ��.��Aƾ�4�����@����� o��g+����u�ڌ��q�)��+֔�ӽ�U9�/*��Ӝ����2�4���?I��pt�~��u��F�h�D�Q�!vӹ6�a��B�E�	z*ԸIuk�tQ& ��0l�*P��M�K��܅F���j5@c;�T|V����㴎�m 7�����}z����!W[N&�������F��s��']�L� � ���xW�W:iM�g���.҅��/r���L��7�R�v�����m�/,揄sG,E��溸 �s�3�}�=�����'8�J?}3����y?T><��*���<��~,,1�)D�d��E�i�t��̾;�l��]!�������J���Ϫ��cK6¡ Kp kXc��a� #\�.�F!uo�]��ʝ4�+E^l��=Un^���z��.�+�Bw^F���U�8�m�O��e��'�ɽ~W3)���A�I��S�t.�ޤ���{WI푙Z/
�B�}x�M
ۤj�9J�y��9�Z5�H�Q9����;��++�n�^��K��g[��s?a<�F�%�9�|qgˣ0����׈010�k-=��u��P6#�F9���� r����,݈�-�֕�ќ�R����ŋT����3���F�dkxV��znP0e4A{�x�~��R1��]t<���I&�"kv�'��`��RI�1S�'*Rlk��R�!���1���ĥpe��x��v���Xe��>�����4�.��
iͳ���c�/�ACJ��]l"�4�m�p������]�jk�񯕲h!�ǩ�DS4�K]]t��Β�u�Yl�[L�Qu���O¦ZG�I���5O��'��#~3U䏭��t��Zu]���t�]��f酉�YО[N�͙h):�m���YYOjZ�z�QZ9���%e�`f>���oXų*�J�W�]�@&�Fs�pP3F������*c�c�BE(�˕�FI:���+:t�j�3��IϠ�(~UAl�Yw��Z4ɥ��ƭ��������F��ѯFr�������%T) 55X����-���uc���W֑h(�wr%���|%5�,#p/%SZT+�M35dT �����n���7A���-T��m�[.˾j ���v���(��(�L6���b�0���&$�������&l��ow{~�ǚ�h�)�G9�[�i��N^�B�Z���:��yc&Z9���r�q�G)jvWnvxV9�2$2�3�+�q�b���+�OEuT:&�	�U��lw�*�A9��9�Hy�I��zm���|~=r��ݜ�	]�LtW�,�����T���J���6C;Sfk1*����5ڧH�É�@t��Z)�E�T����:�pܫ��%UptiLl�薜[�0mWp�:&�
O��;k���/&r�:X(����r~�J��7��Ms#vc!�Q����U|��15&hQ;���M:��2�W�x���!���	��|�sM1z�ߩ���~�+���բh5���=�1sVa�h�C)��^Ҭ᫸��ae�u��͚[*�{�"�*�P"���+��^�:���ڈHI�������Z#�>��W�K��3�����S��e�ƕ�(���%�FuM���5wP�if���Q�Kd���|E���=��i�J�C��{�eռ��c9'3b��
[�eM������K��F��F'Ezceߺ��S��<R\&�)�[�x����ٍq/*�]m����]��OZ�����v�P��g��p:�B�ݐ��s�\�������<<��|,���ma²�#<�>���t���g�0��5��W�`��+	�cl��`��9�ND�S�Ҹ�`�^�렬Bm����1[�.�&8�	<��~��t��Z�,�7V%�g���UgW.����tO
�&]��~[�]Lv�EhP@�Tx�_��-��G� �&����m���NAyJUs��:���.����*a��2Cz�G3��`�p�JɎ*M>��k��s�L@�r��u��O>?)F��2��/�F�֕0�L�KD��c�lj׾x���U'g��O:]���ݡ�k֮Fo�ldGҧ�Iź ���b���t.�h��Qy�q�SBQ������vT����j�����f���%<�t��ﵒ�͹f�>'��J�!�2����|6ݩN�1�M�F�B��m;ո���G)X;���.���4�n�|v:y6�RNG{2��\�sc�[̣�.��ڛ{pr�rt�)4�ٝl�\Z͝Ҷ�f���rz!Ce���=�.D��ߨ~z%�VUE�</�Tਗբ�%|v�G)|m���VZ�h��eT�'7�Ю���ٰPPC�hU41.9��E���Zt\V�����= ��K廟.��nj[4���
iP)�Bg^*����3B���S3��f�֞�ܥے�����GD���$�f�:���O����¡�G6��Kk���Ŋ�c��yz)�T/n��M%��4ܝ�q�[6uw�FS�A�XDbS�SC4�˩��(���>��+>�F\�}#R�2�Cm���M�ঘ���g�.�1�� ��ɗ1}�;xK���߶�~R�^�
��?�g�����j����ġ�2lK�n�O�<)�v:"��g5�
P��SJ`����f���R�2�u1E�֮7����/T��I�C�<���b��8ݘʕ�x0�w>�ŶK��i�t��B@��zX�a�[�a�nܐz��'���^d8?����ڴE�g=���nB%M<S1�I��s�/��BLQ�[l"�cOP8Kp@͞�j�ߒ|;��×�X�ݢ��M�l;đצ���5��۶ۘ�k�~�Ş\��i�DW<��+����O��:f��J�oW"!�d��ZH�K7��a}�{+{�)��g�&��a��ha���ۃ�ӧ��B��[X�M��+ �fD)� ȥ����9Ċ'WM�w�o8Hr�������]#W�O8�FL�h�Ε.ƺ� \��	�}B�d�2XCk<0*t
��g2�°������FJ��O>��`N�b�d&��t�+�6��S%�Y� (�@����n�-�b��oZ5J�Ddf�d�����f��O5�XG��lㄔ㾨�"|b <)��"�l�4<�^���_q�
T��`�%fq���ΫΫ�zp�&l[Fx�\�1�9��HH��Ff��z\�ƀP:��YYc�1flfv��8)2���\�uT�D�)��Ϫ��cKl*9w�&F��Pw�+V���f�έ��0'�mק�lٲ_h�U�{⪡�u���\|�E�ﲤ�Q�. \OK��]�/�* �s��3t(��д.�oR}z��]'�fV��.�SN0_�d^}C��ئ�b���r1X�;��l�2\[�3%�M�� �v�B�h�{���R�ae#D����ݣSn_d/R�k�r����]{`�����Q�k�s:*b9��2>34����u�E?��@�\L�)���WJ�ˡ_��Y��>�゙�;��[(�M�Q�r�FpU�����EG0ۙc-6����j��K�Ov�������w��}�n��d�z\_^�_5:ý�!�;�Oee�g�s-�f�}��|c�"s�&�E{�/,7�}���ق�MJI~#%F!��6��]��KE������1�K���3�Խ��s�X�[W�y�\qy�^`�;���8�g�N.T�:��Sfߒ�!�:�4SP@I�=eSn�UޣH����>�(�/���.��#8A0�Ц��>)N�:��~JJ~U<뭄V���0���8��+I;�?R��5�� ��2�R7]Rë�����So̵�!��C��Eք�Y��H���%n�𹺝1�ܯ=@"|A ɞ�cM"�mhB����c&�@F2�12T+2:�b��T%�?G�u�g���R �����x�Q��r9O�q?.��s�_c⫤���E�Z1�����*�A����gtV��D�u�߇K�����lW���u%{���*��l��
IY�f�#�F�)a�̦P��1�OL1-�6�Ì�]w��f�Vbt	�u�9<��!	�3-���Rr�.��e�~u-���&Z,uDE�>�E1_�i�R���-1=f+ҕ:7Y-t�r�u���a9�5�N��o��������m�m��m�m��m�o��m�h�m���m���6�6��m�m��m�m����1����1����1�����1��Sm�cm��l�X�`���m�m���l��m�cm���`���M�����6�6��6�6���`����(+$�k/L��&{�B �������)��r�lիX}�V�:���]�i��emmݫ�Vյ4��ֺs�Z��j��JmAѥ����U�TV��Tե5hH�ČH,�V����JV��֊�hU,�Z�������53m�7��b��D�&��[Tld��Z�-��M��+Y��V�j�V���٪�� ���:�Ɲk������@�n�.�� ��9�읶n�y�6}k��wIO� //{�������kN� �:P w��� |�p  �\����
��T���=����| ���wmt���@;��P�hMJ��������{�z"�6Y��Km=� .���΍ikV����ع���\y�M��S������m���sֽTc�N�۰u�֭%Z6��� �M�>�����S^��wp��ݯN�Ūg���l��=n�u���7��Ju���{�m�β�Ƅ��A�� ��Ml�KN�u�T֦��M���	�S����ov��2�o^��d���{ç�H�xkY[,J5_ ���D���w���^�J{�yE{f{��{N�uV{�y�u���5��ڷ��Q]�{�ۻW{��T�j��1&����t���}���ͫݽy��{��T�Տxy�pP�� ���u�.��A�EY��3e� �6O� ���u�=�Ұ`	���U���V�wk�wak�46�c���PȲ��� -���6m�Z�[j2@�� ���j�k;��.�P_      &)MT 2m@ 0�M  OhaJU%       �{F&�UM  h     O�J��� �	����JP���C�2h�0�I ��44�&�=#F����>_�ݎ|����߇<�ξq��:.�y.��$$$����S�@����@4 BB����@k����BH��u�����?����g���v����PI!�@@�!ݐ�� z0�A�h�&�+ �I	 �ۿ����h��������$ I 9�u��fo��C�X����&O��'������Q^��L��?�?72��{v�/l�ƽU1��φr�<���S��.8���q)��-��G3�u�Z;�]�oQχa)�]ou;��\���ʱe+#��uy��Z����v�\�v��`��Vշw�cPE�γ�G�Sf�V,[zr�,C
ι:����ز-����w��*<Y`���6]�֓����Ye�I��Mu�
7Y��;bo,hV��]m��)q���;c^'��l��E��uz��m���rK�+ݡE,���ZV���g�r��ϝ��fUҧD�����Z�!��g�]i�۶���a���[J����=ZSB��u�]��u4�Q?i�zSU�+�ܬ\���>�:���-vkm���|r�
�Zpw[�F���o�+���ǻ�6�Պ���v��N��+b��7h�'R��4V[K(�N|wsh���{׽I���,S@"Y�@�Y�s���÷u��7���f��f��:ŀ�8cAٱǫ�Hcx�X���l�3p`�v��]�ρ)����L��޾;�����NbcoQ.Z0��cQ�Y�%�{̍���7H1�G]_Wk�º���>OEzmYĵ��U��>�\t�z�������:��7B�,���R���lX�ά�zKA��<�6�G7u��֛d�]��z��ga�&GV�oX���YARK��I��*b$�
��Y�����G�DMz���7l��M�V�nά�t��1�B�H�(�Yx�r��z�aWJ�I����T�2�-�h����2Uvoe-;x�]��]'K�m0�o����g����\j��}{���`�B��<�fV�ݏԶޛ� �uc�4��o�V�VVS�k�L Rnլ�W����K',a��cz��oko��6�3i�DYb�Oe����k��Ch����]vΟ���n���7�e�е���A�s�zS�#�~j�^I�S��s���񓪊+,U��b���k9�� �m���U�Gu<���6ޅx�u��>6���}t�!����G��{��m��P���k�oV�v�E��)�k�}����ƦP3`�n��*X�y�Vz`��Qc%�U�<�m��4:�|���C1�Ֆ�#zF���,;4��V��Ҟ�����y��0��M,�V���j�n:v��y�=��Rg`H���"�Ż*�e+;�c0�ܻ�r�n�Eh\�h����U��C8���j��w�0�j_?�wB�Wsս�x�-^}�+�n��yE�v���[��n-��es(�W�pכ�w�g?�Fٶ�2�2��дC�*���X��V�i�p������O�2���\.��5>&�ہv�J�����q��ҭ���l�Ҥ�hn���@e��.�h���*bЋ��#����46p���s�����ﯕU��m�I����+������oUmn%�o�O�������S�i3�hݷH���503@tW�Q`*K�g �n����W�vֳ�-?xopP8�RVƵ��v�Z��mZuŖMZe�[d�7`�n��F���P����EyV���vks���^i�غ�9a�M���C��@����]Y�֌�l���eq����q�}Y񳹛�V���	�}�o0��J�	5�m[Ÿvaos �:!wn������(��@wR*��x�,��-���%7�����J�č��&�27��U���6�m�x��U]W"z�e ��p��[��u��DZ�Y�N�l��/��XvaeI4],���j�^���v��O|���l�"���o�r<���|����oR]�A�N-�Z�7����L�O�|���4"���[U� }�u����6���-�;��"�M�;����ن� �h���֤�A�XQD^5�1���U����Pڽi�k��R<�t����X$f�W�m�8ҮZVR�O����k�n�	@;:�WvY�-R}V�*N��{�����n��޽%�J��f�=��vX������>�l�e����K���Օ[����j�Vj&�mqcس���cU��Zi�Z;��Y�'�6���W���/8�y�i�K�f�o3�E�H��
��ݶ��f�0�V��Ӝoz��`�ͭ�;�cӀ0U0(��v[�ڹv�W�Z�yG��K�8Ѽۢ��4����*�0f]�&�n�Wܩ���b�f�-3u�mhZ44���he� I���l��\y��eصX�轳�o5w0��ī��n���u�n���<�zA���=�6����+o��-PY�w{/�4���Kqh�ܞyd�]�z��]5J�k�/v�R.�rN���L��v��2�/(]h�v��J�e{oih
xP*�.k[Uu��`���cӘ3+m�-�"�V�xl��Z5�N�/���ǎ����t�Oy�x]��{���B�#�/�ZUp���=��:�Iy�S�J���x�x��m����4����7�U��iMY�d>����YL:��u�g��-ֱb�V_�y?.��r�U��Nj�"�km`�B��do`X��R���-��6�ν�v�U�envq�薖*/�z��mj�e��wJ�k���NRڲ�b���]���^����+��4���b�`<�R�v�pʴl,�ծƽ������\��X+R5
+�@Z�P�3⓼'
lVVM�E�ՌU���κ�T0Ҿ۠7oJͫ�h�.�o;�Le�{�Y�뵴Y��n��V��!��XܠÃ��4c�I!n����}�G��EվUv��]�eCl��ޝb�=ϟ������o<*���V�ՙt+�}��;5��
��lV�ʱa�:siuZϛ[�O������ �F�������7v(�5�'@kZ���gX�����-�%Q�T�V�V�Fk�gRN�|3s/���1D�L���u�{��cY���4�l v
{�^�kC��v��cr��Q���h�k>�@���h�Q����������R<^r�פu+��H�i�%|�w�f�`�Y�GX7���q-5Έt���ͤw@��b�i����g9��oP�P�l.�9�>+8Q���'��ioBx����Vu�I�,����i��]�,�̇��hmn�o#ά�]������*�m�9��?i;�|S�Ԃh�v*����66�1$ˡG��hԩ����������b��Ӝ���`nr�V�7ŀ�$M���Mn��`��yZ~8���#2��
ȼ�tnq���������������z�_^S�{v��2]`x;(^���玭垠�-��=yB��
���fe&����i�s�����]��x�{|��˭ <}��Z9VI��Z�Y�s�Y�i���c��X�Y�I|j��/���,�5���j����
�(����J�>�VCy���xuC3�t�	�(���(��k��Ny�(ZaRf�ZkwO{����������L&����P� �W˱���t�qyuոZks�n�<��v�sz(*��k�˲�.i��ͭ�t۲\Ce��Wv�`;\	������ItsN]����:��o��� m-��������*G�~�&|���a���!��i���t�{�GN�x��H�`j�8��C.�
��V~t�t���]�:��7ά�`�|ot�Cm�W��2�v^�I�m!�-&u;V��U�������OW'����74����V��	cF��Y���:t���xW6�*7M��\wJt�]�����r�ӑ�sm�
�l���T�3�iɐ�Z��[��S:��c)P��N��}��Q����� ��p*'S��WON�V*��'��V�X�	>����[7Ռ�/s���vQ[�>k]�����7�6�����g��{�E5:~��A�>{=����¥8���X{���h���gy;d�H�{�K�] ���E5�GR��b�yV�����{)�܌ɻ�9\���LX;�8��|�G�h�M�2N�C�8���jyWWg;T�^u��<����n����sL�j��hWT��fF�m}�AM�^�i�Ow
ȵf�2�=3Vc�U`�� 2*e�H܋��6�=�GC���ǭ�.�$f��o���)��V��ƃ�"�+��g]�n����9��
�C+��$6��t�J0�V�W���_LD��,��n]�2��)^mv�}u�|�����bX�K�U(���
s�Ø�eo^iZ��)���F|���=n�L:������}�Q����mϱ]	��F��/��+����:��4��#&*�s����'[�6]Ѣb}r׈fPͩ�T���1uEN�o3�h�̎��2�8e,�f!�Y�T�s��/r��������%J%�ON�-�y�¦�Ur��n�C��8���A�ۄ`m�Jw-���5��9�N��e���fk��Z*�| �x��a�a�mƅ�c����ȏ$�tt�Jw.M��u񴕗���ݜt��5�9��ݼ��N��͹Չ�x�u�==/Y+���l�Z,�ɚrub�#GTֹhw�ژ�Ŝ��3�s����TVﺋ������%�E�w��S0=���=*��vͤ������Y}�/3��+���f๦�T����1�80:ؕ�%�e�X�D��8�N��b��v��9��� %�[�_j���T���;%2�����f�++6� 5�X�r�$�U���� ��-�}�3��bm�ה1��㣰F�H;^ޚ�/��:V�圌 ���Ů�Q��{��,�T�Z��VWwE�12�����;^��mp��>4c��v�)*me}Xɇ\t�;e8�i����5����Ԫޓ[nM�pδ`R�a�����	���T��=���Y��X���Yb\˓mROr��*�&�ܝ7`5	��C�S��,<�Yҳ��=FM?&+v4һ#�SaŘB��ؖ����ق�_uX�Y[����B�9�;�B�b�tKZWYN��WP��i�����2RC����MԦ�9��o*�Շ�d�(��Y}�ݬn+#/�����a;��z˺HTS�X�i�\��&�#��e��_ �8����\�
�M�>�1-+7�dZ��dМaw�۹G��l�M�ް)Ccө��_����{g�5̫�{�G�<����:%��=ZH6���:�npWH���v:f>^�@E>�f�1d�1�P�����{�����65J�X�(!��ժZ��x�k��o�@E���)��CwFq4o�ze�goq�7��aMȂ��Z�ox6�[=u�[������l��˙ri9eD��6��5�iYf%M�0����w��*�Wfj��n�8,��3���m
�]��q��m�{3�f���@�|Nia��r�u�ă
��];u����NTݭ�2i�и�����؀%�Ҹ�J'BoR� �����-�#*�Y�z��GFN�)u��>�/�
�͙˞���틷Fv��n1�����W�âd�9P6�_e/���8��;���):�P�1�/�����>��� tqi�\Z��f���6�%���3x٩�־�thXC�,R�a�4)���72u�+U�Ѱ���b����H�z	�(�9l`�j��.�r_] l�����kT�8�+�Hjƅ)ݥ]n�Q���#fV+���j��a�%��-����(W>�=��I2w��B�� �+(�u��	�ɼ1[@o	K��.����[���|�Ͻ��������z"��Ⱃ0��kG��^�@3��w;�e�o�j�K$�yxzCGiYo� �m�;����J�.����J�#��]�T�b�S��]LsX�wQ�WPr�%����&]=Iu�`�	���E����2O�ٷ�]�+]��t4���\������ilU1P��|��]zrȳ��s�3����齍�Vdb�(،��KS�bB�5 F�"@�@8`�G�+r��R�����y�V|���H�k���Ã�0TB )�l>�Iv��Q�v�)yR�Z�V�J�f�(9�a9��t	Ȳ9�W2*pW#��\8�E���Z�.����Av/cT����;N=�ɐ�Am:n�k;e.�f&�9�!�w�x���l��JU�K�$Y�MS����Eˡ*!���f<���hRx��*��	�.��O7����i�A9	Vɜ�t�K3^�.�s�Vs��`�q��e)]ij͂��cS8��W�^�h��5oY����/�
�f�͇�.��	�3]���QvNgoA�J��/xoQ�����-�jZ��
^>�
�[i;�Z{��I��7V��96\3�,%��wS��z�Y䍺�\H�8^8�}�������[�Be}`��SP��b�x&e���ơȕx���X�r�E[�|_e��H�3.�@r뷹*�7.�0[	1{\�!�h��?�Ŭ��77�4Uݓ	����JoR��=1f��1��)k�[������­Kיq�T��N�K���D��%k�
�>*��W6��*�qg*K������w۠����t����JP���M_^@��a	t#���'�~���1�rjfZ�Ӱp�RďqR���\�
|��R�7�Y�$.jC��<��@��Z�n�{�)c��J�Oaf�0�Y�Z�����8̠�PaPrlT�����"�!���ʮ��������wz���֎֌�-\b�x��j�����]^�{��r��a�[w)�& �H�Y����[o��sg䮚�c�a+n#�!�L:·k9�K�5-��T�Q��i��!���#����wfHʖz͙�K��B��� �S;��!����a�H]�gWkم<�\eT��\g�����7�Zn59'�֠�R�N�l2�d�w|�n�CB͹ɹ&ir�6ֻ/aG������2�.�����F�-�|\Oa-7��$�X�sX��h!5���å[{!ڐ��rT� �]o+�br$mhOe�1&��箼�h�����|�����J���v�Y׵2��ެ�3�i� �9a�m�K"%�v��k:2P�f��L&�lT���PL}PֺkL�ɲ������H<�Y�&6�
�zVk��ř�{��Ku�$��9nRv���2ӹګtm�*]��ǐ�p�2p�V��v�7��(L{���MϑѤ��+ �ȶ�|�Qشp�9,�. �-c��� ��2t�z�!f���/&-b�`9(��� �fƓ��
�� ��Ho(��g1�6f��+w�T
�>��+��)Fpk[}n��5cf���-h!㦺���&�U���Lr8{�^����*JUku��ǎ���4�B�z�J�PҝvGk��OI�����Hf���`oSN���i�]��0�M'6��V6\m��}��Wۍ����A�sn
+:��F��Q�:�D�8V�Nj�v�J��k&t!�)�[�Kd�	l�GmK㛧�X]+};P��奛�52���	WIZ��r�ǐto���R���iѦVei�.uX���̩�88����;R�E��.�V�8�ȎmlC~��յ��Q���k�l�T쮝��	06�m�S�w۷�[�u��n��MY�SxJn1��]mm@��#�e<�ڌ�Hq��+��S*�4��I\N�(Uuʺ:��`t�̽����c2���؅{ �w����;B�1)�������o��Ԩ��>���G3���@�o�y�䐐 �;�HO���U���h���>���?�c��w��k�	���%�V�g�|�Ӻ�+.�qG��Xx�;"��$��]�8�%�����u���nq�_%V9�[�2Վu�|yҚ�T���� �K8P����]K�θ�%\o�|� ��#'e�`󦇳v�r�g�r^ ,!
;Wk���I�Yy�v���,*B�j7�]leW�	�*�d���5��N��a�sĺ��m�!#��۹7�l:��1{J�ɔ
X�2aܹ{Z5�]�C�bը����Q1�X�<�*����;I˾�S���|EAu+FT&�J�.����(�ԏ��P�L�[-]T-��+�g�ʑ��7��T��b�v�'{`�T2�ao���6Y���@+�c��	�}]:u�jŃ��k�����8��]�\oB�V�Z�AQo[-9`e=�D;�e���TM*si%7�Q�w(���)i��袕ǧef�KC9W��9C-�p��W1�.S��aO�]�"S<���*�18��ɠXU)4,�w�fe &�kx�Ri Q���w��.p�qj�1p҃�mw+Q-�
���ߧ
`t81��.<�o�)6�wK�M+olO+�|fv.gt'f$��a�j���[������;��X��ok��CC����vR��[�hb�JT6���{�o+#1:g�q˔��x �K�ؐ�1حi�\�ty��r㥩ތ6s �Ӹ��jU�kإ�s{��3�j sz���>�m��o'P,��m�p6 M�ݧ�j&�R��9�ͻW����ؽ_Fx)�j�)�K�{n�+QêY7�W&��%əޫ+�N4�o],��1�IjSG-��t63gQ�O�r͇o�gv����@ԶI�uk�²�3����$�����V��2��&�-'�ͩJ��=y)�ff�[Ƹ����hޓ�i������Qa��_ܥ#�Q��R�e������G��ې�_V�ʹ!o^aƋ5�9��߬6�kMs�.�2uۢS��r���9 γ;K{�e�P��B]�����\�^T�M���,����ӻA�/0d��t�lvU�w�i1����F��6����MhB%��Ef��Èk�ә�吪��t�9�ADra�'��*�{nk�	�]v�5�k�2�IP
�9'գ�=���P�ktz|�4mZ�[����`���3)*�cC�� V^28,�n_�| �3���)W�=%�9C4���3�!yI�D���ֹ�&�%�B�2�C�JҖӶ��:Ʊ2R5��W�}��O4�܋z�T���A�]P�z�q�������1��:�f��Ra�iŠ,�Cx�8qF�H�4�rƗ2���vun;1�6�m���ZX�k�"�2OK�N�="������TK:OTw�V�aЬU�φ�聫�Tdl+z����S#�[����o,���Ɍ�.�Z9Q��r\O��l��e����ݢ�dm!i�W�ILC�X��@��B�;��y��͈��t&jt�V+Z�;nP�q����nL��.ō�*я� �e�4��m!��!�Y�z�5�������w���2!���b�d�)��ZE���يf��j鬧�Hp�Mݳ9[�b��'I$�ʨcR�Z7��uo+����vZ'�4պ|΢.ʡ{7+tP8Kc�li\+N�=N�c5y�uN�v�t5��n��K���j�i�uD�)S�x_�� )��:��tEL��mԲD�t��u$_��]q�v���F1����!]���#9 �ϴ��R��Z���O�����e�%��u�^Gd��l�XN}�7{�"9υG3n�[.��; Br�*�����$D�Ǖ!f�n-�uo;mm���魬t�O�}˩�ˋ�+�"�����QԆ��3[���V�d���>�Hw1�@D��U��,��>Rv��F�,��u
'�0Pϭ�R@�}�o/�-u���Mvg4��(fM/j1m�BU��$Ψ�6���^��rn����7A@*TϹe-�V	v�����y�o}��(�y��AjM�P�E�m�j.�&v�W�*R҅M�%�F�\����@Ӵ;�"���j
�Ӓj���8p�e��DB��[F�:��\�n��r]�\�R��d��Xl<�t���bͭ�'µқF]-)7����Wf��9{�:]��%�ˡ��nerK�٤�̝��qah]5�V�m��7�f]h�ĩ�V*��%'�&t�V��JY5�ˍ%f����QQ;�p��Y�E�swn�Z�{-v���t7����-"�	�3��-��ċ��t��d^��V�e��:���W�`N��C�y�]B��"�Q�u�F�x������+*�QZ��ie!�8�s�0V�4�a��Kq*&���u�D3�2��]�G,�n����������]+(m(��{*�IP�Jv�`�Z�'v]��+0� �7��`=Z�m^���	��nS�ҝ7K���n<J��������ۄ^��CL���ɝB�J�;�0�<����t(�9/�}�
�ߙ���A&���A[����ͱ���컬�n>b�f1�w6�-�.�Z#è��"�6�5��{�Py(��%j�]4V�YZp #T���wVR�����33��k��3�Ԧ�h�S~,�=�{��2jF>���W��N��L�	 ���] ]�v�aKͺk�b7�ҳ��ܣ��A��y�R[�H��V8
�,ϐz���=��-�re��lR$�K-��O�(;)fJӺ�\h`Q�p�ܾ`V��t��³��s�lb���GW;�l�����ʘ��P��Z�p����}%�>[w(��hV+
3�Y�}�ڭ���-'�̺J��N�ci�G���$�-c�nauf"�uN�+E"���Uj��U ��F�1���;�EZ/94=����Uqt��g7��E��f�Fn�r�a65�*CVm���g���%���!\�R�n3�9�v�T��/p"7˥��o��烕u����q��ik5�!���@�+;*�ӫ1t��,S�npX��Ao$-.��n�ۤ��ǔ+��!�!���3��d���Z�$�=��]Pu��}�c�狖ֽ�J��ݡx��.�v�I��� �T�Ic�9���]o\�sw�Bi")�H�C���I"0���WV�K�{tv�u��Ӷԭ.ԅ
�fRefZW�*�8p�Q�j�}}��a��}:�d^0hM��W�Q�۲ʱצe2x�w�[l�٧���.�2���Xdx,zKh���̡�V;{�nXvt��(��=�L2��H�"�
)2�P��K5jr�A���@ �<�[©���@��MZ����5%_�P��Wr� JS̷�C��Zo{,�EK�5��/>"�`3&p =��^U�e�����K(B��a[�@o[�I��D�����M�����m�E�>^;f���"�i�9��%%s�K5�h�y���4��+!��2��-��b`�®��`9[���F���2��p/�z,[mq9L����r�p���bN�$�]��or���Uzu�l�A�=ի!��M���ru�9O�:5eޥ>u�⬼�)CM�΅��Ѵ�\�.ڵ���W��$�[ȷ�0w��F��V�}��z�~HZݘcY,�<�oz��8Ҽ��3X� e�s��ڑ:Υ)I-�YG�.�Wj9�-����o�n��]Ӗ�����>�v�0ڔy<�&q����Q%�{�1&��HB�*\B�/,�ѐ� ㌾�)1�T��ݎ��L,r�f �&�t�CCR�;���;2��:��k{S�٬k���{��sUk\]�νD���$ A_��B�����:��0�@S��ߝu��;��'�v�0�F9�y�9G�_U쾘[콓��u�%�oL!�GW;]����$&;t�Wb��X���9H<�;ovР6A�dݛ�&*��'d��FE�M��7�Wѽ��s��G��;�<��w���?IeI�{�j?0V�&I�c)��;(/���~1�W�Ea��q��5�S��yU����wX��m^e�r9�1ӻU��L(b����[=���D��L��b�TN�qxĭ��E���d�u���8�i�����8�n�R�t\DN�xwpI��='U靼#�4V�R�銣 �{�n�G������m�/&��Ef��s���*[]ln�M��rl2�n+|V	�e��ǩ�7��o3�5�uF��
��[R�[&�I+�;��3��Ž���ffN5�Z����e�q].J�����YS0����
&-��qZ6ʥE5����%��4���H���M�J��3-Z.4WV-�ɫ�U˂d��.�pU��Z��`�-��QE���03-n\+[J�̘��Z�-����ċ�2�mc�ff8Z�TE��qP�8&"��bbU�LZ�&�)��*�T���(�-r��r�c��+(�!j�U�4��DEbZi�4a�SCp���)�4�-�j+s3T�4���8
TG3-��I���b������2�����܎ڭ��˰�ou�
G��F�j�$LSl�w$���NFa鿷�~���A_�5�UGV�cD�O�6����{�掋���pO)�����y��sʙ�"�L@��zm[���\Pk�,�U��fuӋ��!��{�Vm����ƒ�	h��Qx4QB�&}7ٮ�)Ӎ�Wv�,�¨��r��y�i�쳶�aQ��9�{�F��JD��^Az���0��GX.��� ��&3m�o�`����:,�F|�f��%�Klo N���(K�f�%��H���}��m~��x�Q�N~�&��&3+2~��:w����L5ιnk�J$�~�qE�;��ְ%P�L�X��U��9ʡ��1�n�����S��R�{+'�;n�F�6��Nh�O<�ū{�j'&���z��ECGݕ�>D6����XG��x�zyO	ֻ�{���e/8��[FLf:�v�鞠g5��U��(dKW�#�]#gn�ucL��A�F�9��V�+��Hz��pO^���X�����S4�/Y�R��{sO��g$�A���䮆J���2�3Kҟ��|��)1d+�fC��w���OR L���� �޻窼,a�����c�V�&J
��l]�m�9�ɛC�Y��a�v�{O�I1�<;�U���g\nq��o$��ot�c8n	�ZR^�i���q��=t�����@'�H9�go��@��}8������T)cí�y!�g��a�qt��j�g��f����P�U��ێ��U�jU�L������Zx0�u�Q��yw"��2�}���������Q���t�ܞ3��"����z8�����3�lh�VF����k3�\�]�ٓ-���gB�*���挋�l��ڣF.���kKڬ�2IQ���y*�5٪�C8ҿF�u��8����W��r�e�i��S��]\��#[��-��Z��%���W�3x�6�Q�2�:wEY���a�bt�M���m���q䓏�ȟ jp�{�\�A����U��k�'�@"W�cczx��V�tɱ�۴�C�D� ��"r:7RF�i��5V28W�̼D����T����<�m�^_�J���5��bv� ��R���@�w�Rl��2T]�jUSQ�#����Ռ*-[mĽ�oP��"�2��7�0��ļZmMܝ{6v��Fm�,nd�O���xS�`<T��V�GDվ��74k��O7�UeE����^JH��Sk�+�~Z��*ˋ��?:(>�<�m�ݶi���B<���
�����ʮN�Z.J*�+��b+�]�w(�Ӛ;���)�%$�u�@Y�縛g�:¹�ݬ�\�s����Y��I5�����_Uj��a:�8��ltq��"MC<׉{,s��lj=Z%���,�2a� [�(@Q�S��G.���\C�JpV��v�;'��[8��T�Ưf�:�$��u�H	�Z1��=#�.a�V�աqH'+�˛��!d5�n�)��pA���v��Gk*8Uڿ,w�Ȋ]�p��?`�3�I��S�=:˩�j���P��n�V���0��J�%��F��g'�k8b�뺖r�M����`q3ӑ�ӈ��a�S/�Y%�[�>��H���\�(�D�������/{���?�1���о��2E�.��ђR���U�Ū�t�|�D쫝�.�L�ӗ(T�gN��b2K��#����C�Rs>�21�VY[:�:"�x��p�g/o�m��:.�݅O\�'tzV���.��e�(��*G�7�>����y�2��@z���c���pP�\�QӷpK��ǚ��ݮ&Ro��c]�*��lr���& Z<���{��lq�{R��^�}����Dl������"s�x����I�^��2���+1�u�25��Z�r2���_����jF�;w���<9��1{�߈W��5�]�\��W&����%F!�+��c@�G(0wV��;�d4�c�V&pD��53�H·I���z����/���˼|g5:1�Ѯˁ��w�����7�f��k|�E�'�kPL��Z/!�{��|.n#��k+zLV�%�\ƴ�WE��q�9
kH�J�;�5u�R)��
���y[��~�PD_[�t0��a�ç��w��{rz�i��j��ծE��4ޭe l��,\��R�XucFJ�19��x^�G��"�Kp�\u��跶�G75FhH�%��$�S�a\�|�tד�nެ�F���F'9��8��ך�W��tL�M�4��ɣywx�ce*�vvor�il��4a��L`��~}�qp��5�j/Zț��4,�aP�r�7�\�A.y�ņ���f��ʜ�l�ޛ�랚 u���H3�ѻ��ؚ��<<����%������CU�e�<a:m�p�����Y�ۊ��b�+w�8ή����h�ܜf2�6E��Z��U�3uf�eu��a��N��Akƍi��%�#z�LO��� �w7)vج�b�7z��gæ�	�M�Ds��*�cW�ܜZ��E97!�9B�{�AJv_�,�/i��H��M�w�Q�L=
n�끒�3^J���<���{�N�!R�r��c��Bk+ǆ)����*���k�nf�F�=L��� �|�6�f]�=[���U�ع���!OP��Q����1{)�2ݜ�6��/C\$�J;���"�i��pg�"]���`��J�.z�}Vu�<�E�	�7zD�1�c(w��9�e�7��ns�$w�JE�t|�����B�r�����\�SQ���y�l�$��A�]ɝ��G���l���f1x��V��{����m&�6��5Kp�]s-u��Kt9���4�ʬ�t.^��ԋ���?Loݸ"�@����-�n��]�X�g�bs:��I�]H����j�����-9�:�{hy���_���-Q��.F�z�����ji�]�o�|�@9��<t�����oz0�r�;�O���h��܌9ܗxc�ֲ�tFr����$�6�w ��kˎ;ի�
��b�k�Ď9�<�{#kӓPMH���l~�v���`g[�Ωƭ�/��9�y�\�5��8��a��["�LS]x��f�<TGQu�(U
�U��+��i�M�n��ѻ��ąӇ}��@�q%vl�a�dA�5�N�X�^]D���J�fc׏�V��J�3-�5�:k��2X�s��(WPZ��	���qkl�0��	��+�U�y�ݮ��-r碮=Ge�T��Y�]J�H�*fp�n:)/
v2�T:WY?I�-WWnh�ZW��Uz�4r�8'b�$V˥�~���;hٹ\����a��w,��픚��5}�.k�G������F���)�9T��ħ�&��o��6�����qW�;��`���e�H}+�	��g������h�dITہ��m@A�+��6)���m�����P3��du�J� �-d����}썏��z�d���l�㇞����@r�)\�t:�b\鞕w�f�=��`8�
�2�=���9'm�	D�l���9N9bd��iX�(T紮	�w���qʷX��چKW]-w��E�gD���t�B���.3����[w}E�4����7�YNPKj�G37oj+R�a�r�zu�Q��Y���8X�
�e_�Q��,�p�ɻC��BrV>�%<zwR��sm���˛����A�)�<�a��a
�!K�&��t�H膅E���4'[�v��v���<6����[SƘ�$���4_5B`�;��V���+]��\q�o&oD��\�����;l�9s�Jt,�-�Ɨ{��VE5lǻ�Y{��=t֮�;��!�Ɯu��N���^Wd�ҷ�&"9j�R�R�ıĪW̹lQ�kT�-��`����5j���X�V��1�(�
�X�)]a�P�����q��-Dimb�KSĴ,LEm`�J�VUb���WL֋l�q�Q��4�++��1���i՚\3ڈ��֮%�A�۬�R�0M8�bVƂ�CU�F�Er�Ģ]\uj��P�X�l��DulV��AKiV����Ӭ-[��f9�*jъ�9���cc�q��c�����1�2VԵ�����Yuun�]f35��ƅ+)Ym11-s0�֜3W��1nf���֮:�Y��h��!qֳ.��^�����9^���q�k`��wf�(�����Z@�� ��y�X�cz��d�����[��B]��'�Og;AP~Glw�����˙fz1�6'�m�_^��}t�ڝ꯳N��<�Q���!{9ߺ��CI��q_ ���9��j�=��v��SR�b/g4;���G$D��$�H�ïp)�LU�J궣��7�딿Ĺ���:�݅W�H��g<C<u-cϼҍ���V��˼u�kU;1p�zMC��G�qi��]��=�|�
�ij,��/2_�>��P�k���Ձݹ�J�[���
Q0����<N>���пi�(Y"?N���&���q�J���#4���a���;ŷz������k ���x���|�\r�,u�
i��o�
y�������V�W����=+[X�j�.�:�4*6�a;Ï�}�wW�&h�
�-�r��ZWzI�Ӈr.b�>W�y�p:������=܀t���*�V$�F�g`.�����E:�Z�l�N��b��[^<�>����ä��8�WV�v����0Y�j2�gf����	��Nx�3���A�y�b'�m\�~�\2���\�� ����רV������)ij��a�u�M�fuـޥ�m|ka�5�MPB���=�y�ם`�_�-�egzCr�Cx������
tu'n��-'"��h�����������=s�r$�vr�Oޣ�Ή\�|�s�uM����r|%�Wii�ă�(�ݕ���m�d8��;�))��#�	s��E��D(6�)0�ݗ�󭏥��%��Ю��$�
n�޲�Y� ��,M7cN�=���[+n���M��qk���w��u���,��n��ꍤ@<��9Br$j�f*/�-�l���T�|Y8[[6�@;]bj�U�[���	�l%t�3�՛N���2.�3�4(JǺ�x�f��cr-��{�{�-������X
��O�y��
��I��n��ˁq�������ް����q;�w_=닜��#����o-�5�G+�����KwR^��z��=��}��c5�+F����a��^�{2�<�'.ves��#���m$��*g&0�v;ME�p�D�O%Hn�q<��;u�|���dP�'��v��Hm���pæC�C���0��k����f������t��݁�V
$�s@:`,����w�,�u`o�!�p���j��y��۽f��ǝ@��C�����)�����逡�AI�&�!�6J��9��	<`e��$ӳ/�^x뾺�;$<��HN�k�d�d�Ht��Rx�8OCo,�N�
�v���I�]RT�x�6�8�:�9�N�Y&��!�fb@ِ���jI�!��٘qNX
9�:a0���'�y�w�w�s������{Cp�Ի��}1m�:4n�Tۅ�Px�[��_3)#��{n�A�
9iz�e;v�B����܎��TzBnԗ)���n��rL���}�`��"��I�H'l�ސ�	���C�N�7C�&��9�Xc$�5�:a�Y��ȱ�|]|�&>��yO����}�C�$�qI�Y&j��<`j��@S���t�t�����Bp��:����p��
G�ޏ����T�=��ĝ�i����6�B�dP�!���L�p�I�L�� u�o�y�m����y��&0� t�êt��tÖt�ēfI��&̓�d�%��*�V���NP�6����<���$8|�����CcVC�Nv�=�,��Nv� :d&��	�C{dYtw��\z�k����y�4���4�2VI�P�<<��'l�yC�Hq��$�\P:{a4uI8N�4ä�������k��;��!�6l�d8a�I7`"I�N��HT:d��P�$���;a8{xa̰;Bt����>^��8��M�;d.�(N\�8I�T����$��a�O�0"�"�=}@�m`w���g�혈b�r�0� �d:d���Hkzp°L�v�XNY7M�l<k � �2y�)���<��t�nÔ��NXN�<���C�k�!�����m��@3{'�2y�c$>:<���Z��֩�MK�����	��ye��,���n�� ���k�AG1��^�a�9��^��\=A�D#N#��Y��:񑶤���(��ȕՅ Ks���5�D���� S�͓�I�*�͂�L�L� �&�'	3�$.ԋ'�Hu���5�~s�rv�i8Bv�xj�;$qBr�i�T�9a�:Hr���I�4����2�7������ܕ�$��"���1�r���;a9aϖ��!���qI�$��Ӵ!��a�a��q�[y���y; �Hp���J��<8��;�5ht�t���
e6ON�lqd1��F�I��ז{ї�t����XA�}3�C5���M�2vɮ��C6�)'I��	��H����,&�T���d;d:��/[�ߝ��r(p¤��)����铧ěu`n�gt�H5I�P5I<`e��I�T���7���y�~p�� y9�!6Bp��8aR�퓷�ǔ�x��Hc�ԓL�,'�Րٚ`f���ߎ�w�6�8����4�c��6��,�$���@���'oL'Y&�	4��y�C��v���<�������&00��$���!�Xr�X�ᇈM22v����ၺI�rI��Nu����\����s�!S���C-�d�jC�:`)� r����5���C�O�ِ�	��I�N����w�����7y~0e��(K�J�5�G,�Va�����e�<�y��E^7B0}J��ǩ�+,JZP;j����n�Ow�Fvi	 ��H���S򘈇>��>��I�fY!M��
��"�t�Y&�8N<�b ��'�i�9I�u�^��kכ��~y$;����v�0��0��I�͐�	����P��X���I��!�6�͸�)��뾼��ٓR
@ǔ+��d�xyd�;a:v� �C���6���ɞP8a����k:��9�N�6O9���MY��Ι'ohle�����X�g'(t�t�0����K�zۮ���IP9���n�c	�m�<I;C]R�d��y@�n%as`��C�k��#�/�뭶�>w�PRw倰�2,�= T� p��s���+���6:��3k�IYP��S�C��7��w�Z���v�N��	� �񀰇�u��{�Nݐ7�Ӳt�r�o��N�'�M���|q��\ss^o���$�9N�C���Xt��57�$�Pqa7`e��i�;d��M��');7�������oso9��VC�i&�醹�� �,��v�r�;d��v��"�t��Bv��հ��M�{6��~��:���r��<8�n��]���gv@�0�Θ!��N��v��I:��$�RN�����N8�y��۷m�뗁�L�PMx�4c
����#�G���L�B.���x���R)�l��ה�;k��,M4����gF��;	FI
�M�Q_z=�艘������?:��b��m�t;d4oa8a�sCogHC<��2v��~�!�����^u�o�<ޡ4���Ƞ�!��!�gLL���$�q�� kk!�L5a7a�wH0�)�'}�N7�F�\u�}s�x��fIӺHy���P�!�IX
�'�����L8I�!�ԁ��s����~�����r�ë�g�����t��n���<��U�?v���}��&l[ܓ}�/����{�C���ͬ~��ka�uf��4�OV����(�%f�ֹ���Vˍ�:T�5$�"��S<���} t$���Q����2��l/�J�+֬ˡK����#*ö�q�57V��Hv�B�cc{�A��/^���x~]�8<���CԒԸQ����u���Ζ�3�|e�*�7�����:�c��Kr봬�atu���T�o"� ����gt���EFn��LB�����f�+�26���H�4�c��q�*Np�9�H�v֨z��c��Eȶ)����l��jґ`��7�X��ɼ��Ж�W�q�e�y\"��R%�˭⋌�^d��S�F��=��������j�'���{�잊U��0^�aJs�g�gY����>G6:���x�i��H��a��5g�q��2.I�O#9SgRa>�qf(���;'�'dh�ƶjm��h��_zA��G�x�ȸY��V�������n!����I �c/掿RYͺwO*�;�����B׮`��N߆֞�)����b���NkI�2j�Z+;�_���C|��'g.O��M4���U�.��pzт�ۿ)��\����>����ͱ=W~Z�xg��\�&���[#l}/!�}�+9�Q#d0�+Y�Κ�o}CN�V�0�I1y�n���M�b��E=���{Y~�s���[J��@��.�c�MD\�u&_9�`D�C6ú��\f�UTe���8.��K�ͿHjm��i\R���-�B`�6���,�ŉ�|*��q�ۜ�\Uw�|��:��ӎ�G@���j/�Df�ߵލ�*��5s��K�E�&Κ;,:i�:��xFͺSTa�9R�X��З�6D��l��;��ҩ���ǧe��lQ�-SV�j�$����͝_j��h9|��w:a�+vF���W�mR��n�8+��j�ǢC+o�u,�٣Kwγv6uÎwQ���X�KY�
c�HPW��F��/��ZH1a�Ycw����)�N�O��L��pQ.^���S��[��^�]�TGщVR���p�t�`�sz�6k��]��'�$�Xr��ض��-��̝͕c5�* �'�nv�q=���n�$Ʋ��:�Ywci�t�1Z��$�+r���0uR�7ܖo!�9M�1�}vܻ��ŕQ0�r�s6	i"/+q�BX�mZ:
�ݶ��[�T���NJ���Q�\
r����M�߾dA����v#���7^�w*�0�]# YI�N!fH;gHքMtZF%�+2Das��(�̥���/jr��aQ}�h�κ�s-��͜���fu�v��2R=�c�t%�5�����u^��%L0A��{��Ң������Z�<G{W9͒3A�S��ӥ��h�|G[$d�)�m��V��6�g�jg�m��⟮ ���sD��*Fw*�+)\��&�l�#+���iw����r���`0��rDL���u���HVz�(��w��y�]՚n�;ɻ�/�S\>����<Jֽ.*ς:�
F�<�9!
{2$@{���t��jF���-�I%mY��F̝�X�2���F���k�d����NƭF%`=ĭ�b��{`1E(����G������x��xܳƖWiuWIr-��]S��U���Z�Қ*��T��)sY�V�i�1D�e�劷W5��!��i������t趗Y�1��f��[�\ʉ�J�3��.e���U֬u�2�EQ���L��-3VQƊ�.kSIfR��5�c��ˤ�W2*�b���9J)mX�A�4�Z �l�\���\u����j�t�,��M�N.�fR�R�m�]iW)U�,R��2��
��X��MeD��miMe]X�e]e�%M5r����PbR��+��0-2�L�tܗ)�"��2�.[�\J��]fe2�0Z�ND�MV�sbx������ӎ|��ݡpkj�g9og.��r��:����Top����~�=R�i�������sު���ߪ
�]�]t
z�P6���'ק����+d[EN�j�x�T��ƻ&�c��"�+�M�O��=��9�ugu�Jڮ�4�Y`)�C�2�imC�?=�Vzؾ9^�,c�f�	��0i�ymcx�#���+*�� Q(燻Q�ε���Yl;��hJ�f����q�o-�8%<.�n�w�5v��lC[sT ��m����ҫ�fs$-uS���)��K/�E�u��{4,���1��$�,�̼��;�_B�4iH8]G�9�<'��ND+u�:ZZ���W,G��-�J��ވV�)�?h1�aT�`덃�Y��&z�c�ES�,F�oʘw���A�Ce��R��[\A���v�ґ��i��9�f���z���x4�M��k0�Ѵ�͞�qX�V���59�����H\�˃�T�D՛��B���:����*'X�֛	�W���9 �U�1Wɩ����-	�ZN�ͮW �L�Ze�c{H9�V�q��f� o�#�L�����A����v�;����T'�|�.rlEP��>�A��uOK��PYp�ا�x}����8f�r�Ӕ��Z?-ߡ��S:�܀��(�B�T��	6���^�)6���%�i9�=�Dy"ZM3?�ja���q����]r9uw�_e�=\|��%���ۊ���V�Y�ѯ{����֛��8ч+Fġ��.j�Z�݉1;��w�s�L��=,�$e5��
��6��2a���Q\��םkp��Q�kтH�m�����n6b���H�rt� .�͙���e�ӎsB��AF��P����1Hc䃂i��"�c�h��V��1!H�h���siv�)��
p����V�ױ��ў�-S7�v��(�7������6c���{՞�\�m��(�5��@��1������v!3I�"Q�#����1�������	�1��7架\lrʎ;U�D]GH�z.�nW��^*�l��l����w[y97xYON��n)������-��X-y���o�l>Ts��64qWó"w�6�)����]b�P^M�Y[�ْ=^>�F�F������NpC6Si��DVѢh�L5 ���6I�r�{�J�W�19�E�$$�� 4�e�_>�Y�ٿ&��f�&�;��⸃Uz���8C^n��{o=9���Z��m���4�"�Ꝙo1��*%4�JҬx�uI@���fSs���jZ�#V��r;�ն�q�[ջ�#G���|�G�?vt
��i��q���"��M�8�a�xw���7ψF�亮u�srcT���`�A�ӯ�42vM�!������{�IdUv��o�f	��*�X��C8�UjI��,�I��̻��q�]ܚ�w��@�/�y��
{^�,���r��5"9��q��SI�=�JZ�j�ad�q]tZk1֝�+4q-����ɬ�&�y���g+d.�����iqc�g2�\��)=����Vf=�,E�����5�"�fK�P3^[���bv;e^;�F�r��.�.��"/$X�ہ�y��[�Ԓ� �CH%}���a�����(d�`C�f�á���?}�z��,f�
rr�S���T�d�5]`3�ۚ��'h�M� Q����dt�-��wtsX�y/G:�T��z�F�٬#��oWF�An��F;�	�|�D}o=�
������O1�l��:ՄR�
t��4��=��^Z�1���$�=��9{��[F���3f�79����g�w���ʛ�(�ɶi�Y�C9���g�L��T�ޞ�W�BK�rbk�eL���{c-6�kZ��ܩ�v��u�۫Y�Mi5b*3.n��/c3rM����URXZM�<N���~�-�7%����ì��a]�b�r���)�kyr/�vErI�C6�'v�;g:5�	��cq�C��y.��,�:�}-�$�=���M��aҧ��W&�(��s7������j=!��ܺ�cD��O2��޺*�.�4h�+Z�(�ޑvt��'G�%@*������`�+$U��=���7a��aη��{VE$:��z�PG���`NÎ��IFT2⦜�e���!T���[��Ht�[w]���v���4uͫQ�w��Cp5�� �?�b��!�����lm�e%����vV�s�l�����z"=�I��Q���y�����,�t`ax;m��̖}+=�1�7*��6����b�i^����!�̑�-����N�+��d�#b4K~R�{Y�:2ݝSo���{ϧZY�+�zv\-�5��e���f�E����j�b��5;ŝ�~�B<�о��¶��ζՍ�p�I�/�,9\�&28�j���P�oz�!c�ݤ�-k��dOTƋsE����=��6pi��t�����#j��,�*(~�4�]�2V\wp�}����t��me�)e<NMvq�㶽Pzx��T�VLU����+g%wMg	/QU힏���	䒟��z" ��YY_A�+7�p��&��LTCB^^N��Lہ�W���.P)A����*e��ɱ<�m����CU� �j��>���I)��WI�7Y�ՙ�8E�Ԣ��-$8"X��t8��j�wY���Fз���ER�	�U��o�WdO�N��θoǜ\7�A܃�lN���;Q�74"��n>�]�5rK��+�,t��Oq�A{'�l�AZ�2O.�Y;��w��mt+)`�]�9f��~�� J�B�YJ�xs[�Ń�}[o*Q`r����n�YYs68��J���1�z�T�ݥY�t�%M�*n�FD\����
�=�DI�M�ѳ��`B�C0���&�e`{��P�3�Rs�u���ك	;�)��/�ڄ���Y6�L1���$��P]��~g���m�Ȋ�n��A�\Bߤ>���Vr���Z�a��=�/<2�c�9�O)O��t$U Mײ��7#�c��y5ء�	R��fU�l��6��:�5s�F�u���&G9��!=|D�z�Ʒ�gfw�t צc\l=��"�n����-�{F�r��L�&�I�~����W}=�tZ�<���
��K�s:X����R�����&I۸/-I�,[�LJ��a�N��,aL�L�	rFU�n�]NK�ܡL�T���*J �)g�%@�ж��R����=��)�W@KI���٬ �sr�s4V�� ����\���[����G�|T���I�W�5���҅����nFF_1[4x�<�|©��|]^2��:�[>����E��J���ѹ�9��^��i����"S$�x�Z�K8��c5�RV���t�t{r�Z+����x	�����JFV��-�ܕp+̳�����zog7�2uWiN�Y����k��&LKj��6�TI�M��*V��/� ���co�Lʼ6�#�i�v�.��uH����3ҹ&�uY�����(�!T\�iWe�nw;yV)֝������ אi^y��AG�_�C1s�Qa\�T�ż����[{���*��[�v�wv*�oJ�����<r5%i%^�t�����"�����E=��Ri�HMyT���(^�\ۓ��j��J�])��9�������H����s1g;@�����ҫq�Q��d�<�i�3u���2_QL[���D&�\�no�dl(�P�v��.�T<h�V6�r4�J�[6�C:��3�G��/v�;��B�R��1��$�-C�n\р��^A��Ũܭ���ʾi�u�/8-�C�];��]��oB��Y׷�fb�M�6I���z�g\�Q�U��3��-��\�����q�̬R�2����8�3[��k`f��9�..��pl��C�U�[ż�U;�$$$Si�(��Y���L��)Z��c�,usV�%Z�Zf\�e�Z��4&-�7e���J�S)U4��ʖ���L�:��`�j���6ڵk�.��jܥh��`��u�11�uJ]\�Km�)Q�-F��J�&����dӣT���iuh8�]-�6:�ulեTh����].i� e+��d3)��0J&8��ʔt���P\��U*�s�WY���q��[��]5um��u��`���.�b����(Q�mE�T����(��SHU��J.�˗�(M�&���T��IN2��X��/Y?�԰rS�ɴ������G�K���{ޒS	�"�aZ��U�k��:AqI��:luw�q7��kE^Z�1�u�1�#�e���Sf2�T���l�l��_����(ͮ�-��n�F�D�Z��#/����Ng��,�	m�G#�<�8�:�9�%n�!�7�6Cz�{B�L�CM�\b�;g���6�|3@&��5���EpL$�c6b��<���f�#�y�����Q�g��hն�wF�
�fs,�Ե0��ώzIRm����'��b�Ui�,Q7�К^�ְe����4����y�O0I|��G���JD6���Qũ��H��oOa8�i*���-'y�%�$��G�=	�)��ǮR'6`qUC�Y�[35�e(���6��� P����x��~�no��LU�ս�s������7��ڵf%����tZ��nMF�Ӄ�V)@v^YgV�1r ���L4�d��/Y�Æ<��ޝ�Pi��S���ݷ�Տ4\�1`$^�2(j��S���{��Ѝ"Ń_O9��z�i�k��>wJ���bր�S݅�9ջ��c�q���[��e\��K�ξ�1� p�h�#:U�t�cw�Ӛ铸Q����iuԔ/�Z�W��kj5o0>��f�l��U�{$�[�ޞ.O�}���Al�[����䏞_U���/��Cz�ݛ�+���Gs���3�E�ޚ��R�]�Ƞ�����";��]r"376	�D����H���:-�L�\e��W7�ϯn(k:���j����f��l���[n5�\f%�at�f#/
/4na���/ �p���Sh�M�+�R����w��6x;� ъ�G,�OL���ye{s̚*ǋ�IR�hJ�òm�ӟ[�_T��)^O�:��[�j�bD�ж�5]��WC�t�祺������\S�@b����lWzA�pù�᝵aaq�:�َ&�꯾���p0�gOƝ�f��� �qe"�w���_S�|�.�;�j�5rK��W�P�l�h4%Ɗ��q��d'�zq$�-�WX�p'l��lr�˹=�b/z0i�X_��CGM�X��� ��P��$EFI�e��i���\��wkLe��m�I$�L�=پ��pS�����G�E��ҳ�z7x���0�o8E�g��s9��w4Y� w�]z�V���t�qZ{y�Z���������G'~~35.fC-��BU�֕(�lD�\��Q뼉.���4��9�xkt$s� �ú�1��
Wz����U;B2s���4�����x�9�����\C��q�����o��WN��(j%���@�H��r�<������{kKR�(��!�y#)i�A�ķ=;�GAɚ�_{΍*c���o7*Wx4�3�!� ��0+2HS��b�X�^���}WQy�j5:bFm�U%���9�����ٌ��"֫���-������C[G'����R�\����ޚ�߲.{�{�\��j��#�Y���^[��x�g�{W�X�vѺiyݰm��>�­Ƿ��#�X�E"n��ܬ5����P2��VV#��K�kw�M����̜FR��1��Y&鉆�N~������A��E��*�4��� o��!�f:�NܪU
�MoMh�$�O�3�a������{Qآ�Kâ����-�^��0��Zڡ9M5�����#���q���8����θVY��A
���4j�
���v�m�4ߖC&M�y*����Jֽ�=7�a�����>�+�\�aHܻ���Y�ډUm�\u��)[XCtn\:밹��܏-R�q�F���
��#�
�4U�c�q��=Z�v#�@�M&���֘ق�̺�w��M�0�_D�SЪ7So*Mx*��Q��767�xK)Oh�Η��NKX�V�ݔ`� r9�w��I&���,n:t�X�'\S!z��O@�	NJڳ�XʠM�������Q��T���JO��{Ƶ��ˑ�,�Syw�|�i�ǨR�Y/ ���u]r�<յ�'��+& ���UT�F�^Us|���)�	��d��j�e��T��>�p��׺����zZ�.*�[�������|O��(�R��+��+��7ݔ�w�5��\��|ډzB}M�T��S�u�����޻��������=>�,�!�Z^9M����\�[z�VL�����rǦ��	q���Ŋ���G�d���������돚��&A��hј@��Nw-5�ߦzJ�ǩvR�g�Ztc�7���Nݻ�b�_D���^���BM
L���<��)kT��<�f�c�&�d�+��a��²1��׎/AI1^8�醫4ս��5%�-d0�gj��)���ڥ%���Ѝ��t3����x^�KTf#9�
���z	��Ù��S$M��,..j%��^����ww|����yd}(�skj~�k�����ED(/j�o��4�a�P��G�
+*>�Ƣ��<��jF��Ō�ju�c���l�SN�n����3&s/�����2���
`��;�n`REk��w�a�5aa�M*P؁�y�d���)Q��gp����-�ʍo��r>j�>3���FXԪ���]\�_����=;(:P%B&�"0Y�ͣ3��2��t�ӏ
`med,(TY���(�U�=�Qp
+�]bՇl��pj�S.F*�f6fA�����3��Y�]{#�'rE��r�$������Z7z�jA{�y��o��7mV���I���m�"w�r)c�0R=2�c��+6�֔��+舏z!-��Oc��%I[jT�wkHߘ���X��gw��f����Ÿ+�j��b9��yoK�c>�jq��ޣ#j.:k��R�b��O��{b�m����pK�M�G�S]+�ʺ�r� �vRmld p��/���˹���� ]FӺ�c�\o(۹���12[u�^���<�������*�p�B�����%��)q}6{�}���љx���m`
O�f��7�9ϓ;�{dt��
�����@-4�%aL,��Uf��f�^���SW|?�4iE\��HSS�*�j�\5=�o��:|��Eq"����/-	�a���TU�N�����ٌW+(��C-���G�2�V�P��q�f�.��}s�@��1
���p ������ ��v-h�5��0�:*�{�n~�����,h��c�I�t�VU�[�ȫ�,�zS#gS&�o����X�j�3:0�1�X�z�v��7��	��E�9.��]Nm���
���OL��vr��	ër,+{����������aL|�OO{ǈb�x�&�;E�#�;���	�Y��"k6��}�[��t&����_6[im��G�Z�\�{ۻ��矹�ړ^�`�o`�R��+�g	��6��6r��/*���V
t*�wr�0j~k�:����װjN0R1��جSM�L��U������Md�ڋ�ʳ^~U�~0Fk�. :�a��zݻ^���ދf��ymk��C)P�Xy��
���ݳ��9�\4+���YI��m��q�����R����_�y_h��淐=.��U�qs�4�Z��ҺG����☵ֳ�f-,͍7H1b�	��u�)��S���V��3\�HMk`�Z��j��j�J��7�WF�ᵸ0��:E0�:d��)J��sU�^R0�{#D^�k���^���SE�k�ڐat*�M?�j��$�˻��Oe¬ 4�{��-:���p@����� ���u���뽚�o�ׂ�4�����v�(U
;����0�U)��e��X�I#7M�`��Mۺ@�#��7��V�-d�Ε�2:�#�HN���@�RR[��!�H���bb��M���A�B�v��ދT3�XR?�TY���~�ނ�w�0]�h��-�����A]�0i�7�	t0V$U�QY�d�G�������]�F��+�+�kʛ��-�f��V
R��=���;��6�{fY�SH��A�x�
g���,i�ښQ��l��U��;u�kR�6$e�d<M�<��ї�R�c(ܜUڋ9���g�L��o7�G��M,ѩ��:�YO
I���h�ZN�˭l�&���`�����l����_$��~����Ì���(|-zf�U���q8*vh�%j����>���>��g%L��#�����]Չ^@�pKZ���۬�̗;u�ռG�a5���bT!�p��N�l&��p]�p�&K�X�e�hF�an�M�W�@q���St����F��ɬ�v�k�W�p_x�T 
����WWY�3(֬2�ˬ5��,�EPDm��7*���31�3T.�J\�L\���TB8����VQ���1&%J���h�8������.�ܩKP�ˊ�Y��1++t�J��0D`�T�q�(`���EڴI�L�F[Q�Pm��0�\����)�7�\L�D���\AL���*RVT���$S�"��c�iLE3�\�T��Ufe�2�0̆J+���V2�[e�3,�*�11ɍ���m2,�rb�ecb#�(��iX�R��2���\�J�ڔ���������]�����0H&6b��Z���:����M㛇���"�^���� &�N#eNf]�~�6��+3{T<W��V%\7Zk�r�~d�z��8�W5`-<}�����y{_
�1�Z������}٨�Xk�������i7K�O��LX���7�3bݛ"���z5��T�����.�/�C1��k+8Z��j�u��9�~���f^Gؔ��.4�ڞT�{�*:�/��2+֕S�k�$�k!����f���g+��r@�<.��F%:�N��xOy|�P��}��N 5�� T���0&pmfB
��,0�ĽO��
!P#@���yT;�[�1�}�rn�̼:/������:vh��� g��Sk9�	Qн���0���g�VL���q��v��Q{Z��Z�<�Q gŘ��3�i4�Kڰ�`�e��ݐ0�EL朕���+��+u���G�މOi�Lo���H��K"%�� U+�wn�
�ܘ�N_7?/��5�l�xM?k�Z��`n�´�����K�����ۅ<�*2o]��fGTgGծ����!�uM�@��
i@��[��y���K^�2�2��q�v��Q� N6*,M���g5���zf�ђV�ק}u�~[li(T�>�f7��Ȅ�8�K�ˋ��oٽ�}P���Ǧ�R�!��>;�Xf��1��lѨ��R�\\s����B�l�R��젪��Y5W�݌�U5޲m��F����F,(�\<�������I= >��]P,<8�Ċ�aiE4��guoS�q=�fVʛ��q41J\�!g�����6��C�۠ ̠!vrm��ݗ��&q�s*X�m�S:�b��ބ2�`Y�(�R�	}�{��YL7�8_���Ȱ��$~�Pq��.����f�鬽��P��(�O�"�L+Z��mpwwssĭ\�ѯ�� {aaB����H��LW�����ޞMd�u�g�+-dd.E�ׂ5D4��b�⽑N��o^m�E��U�4�kK�kL$�g\�n�����-3��2�m\�a^5mN5�V���ט.$�eN�p�vǓjI,�j�+|n{�{��zr���K }Q�,Ƃ�5�_9�k�6e*ۜ��W�w}��|(ƞ?��!Q��{�_�8\�ODZة���جZxb��Wf!L��]>q'�9���׺g��I�[�E�޴W	�=GE�7 �9�oTY�eI]nJ�s�y�X�wX�:�X&����)3v�L���Huh	NwW����L�>���6w�Օr>�4���Y��UXa��.�z�l��/Q��Q����a[C��V�5��;���-G
HTԢ�Ǣz�Sb����Z�š����+�k��̈;�>L�^�ю��jv�RY=Jl��;ii�'������i�O`���2.���ǭ�8$+�0�T���{jLwJ���T+/|;�r�p5O*�ŧ��yz��[W5��k�6r>�+��$�w�Onq�X)�(+\�-qm�S�[������-�w��UZ'��`GUF�b����7N�ʸM:�f�^ov-ip��)QFڼlW��ET+��x⵷�tu��2͍f,��LԌ�l_.ʝ�3���Z���'Z�Ѳ��-uɝ�v��"��1c�q5*귥�fmlB7͍�F��h ���G��l\?���<��CM�1��v�'�A��������f���'�G}
�����n�ở�鍉������}�w>����画U8Rq�� ��TtQ�5xHE�Re��{ف�*�.��2,�~����*��a��|�?{HH��g��SF�j�O(x�4�lǉ�D��[ܡ@H�X, ��X��b�R�,���.XYd2��5Ұ5�7^M�h	��>>M�Gy�VOd�`�K�͹r�ӐiM¨VO���f?��i�U]�͘6*�;�K\a���1�7����W��P�n8�e��y�b�c�M*��
�ھU2�}�~�r��!So��Yn�ykwln$��gk�^\�2S�oQ6��}�/P�R�H󽃍c�,�Y�Q�V��Sظ%��G�������~D³�����\SS�u��;�U���z72�?���._�9�q<-�Aف| ��}��;2{/�
\��h�O6���,�^�����z��=���M�N���+�T(���]� �
�b#3w��&zj�֬�O)�V�,BјV*<�1�7/��L����N7Gˇ����������>zt$TYV�;����������dU-d�Ei����pS��{G��2:����u�/ׇ�/9"]�p���<VoL�n���{Z����&�&ڡiqpsRp��~�k}7�ݦ��X*���~_]q<t{~J�)�WE��acˆ���ΣZu�`{�G��:��w�#i��FS�m]�mS��H�:��ːI��.��
�JVgi��N���Q5ya��J������Ҁ�̆;k�K�8�=#l59W�Q�'�vzNy���$R}ʜkK&��B���1��`����u�»����(�}Q�Q=�&�kJT�}ތ(Xy���ٝ�,W���r��	�PX����s^4D�,��8����&�-����^~n%�r9�MC�<�.����3�|J�س�UόLǈ>Cq��bE����sRk�2��Ln�j�����,L���Li�WJ.�5Ǫ�z���@U�*Z�k�GO5�TBi�eA�ҷ��<���`��?:^0z]c��K�CxT��t̺���Rla��k�YhR�&��k
�ċzk�A�W���C���W���}oС�;/���z|����V�I|.��Ŕ��$w3��v���n��)��u줯V��*k{8 W��Dx�i��F�}18x,��P�C��5��O�O�j«:=��{~����ξ\��= d�v5�6����@��q�fT��nO���"��HR��h��^X8y%�)�&��x�r�k�Z�a���[YMX��
4(X�nN(��ȁ�g�7��W�2;�3L1M��+S��a{n�;w�\��^:�Ƨ_�δ#�	Pf�����˿v�j��/�
�c��8�z����Uv�Tn;��]M/1P�(;�>L�kʼ�'i��Pu��G�6�8�&:�PWS��B�h
��}�W�|s��"�}yd�~"�,����݌�PZ���KW�S!v��r.���e\
h��rt�닀g��*�A��8h�U���(���J+y��گ�u��=�n@�T�p3		8UI3
�+	����z(��i���D�q��7[%W��W
\���VoӀFk��u5�SͫWB�`��\�ZWw{IY��
*e���m_n����	�2E�������7�1s�Z��@�lsi-TዏfB��
E��K��luA���������[�~ƛi�x���iќ���dۨ )�d�90%UA��7)שT7sቪ��\��_��X���u��Q/��ӱ����CRq��A��v+��nÐ�+�!W���!AYw�kϲ�>6s�|��6�ӯ;������ȣ�F��.�c��Y��j�*����,ʾPc�i��Ӗ
Ķ��������O�	����}t��uC�1���{X��Yͷ�6B�᯵�j��s3+�i�$�����J�}=T���v��zsGYҪ�%q�D��́2���UUUT�?v�b?M�F��f8B&���W�'�(�M�FU'��߶�9�,܌!S�t	W�K˦��#xZ\ ur�C����j�e�ߍ��9�:_�(��Dj˾��� ���iR�L�(�b��x�S��1�ű2L`�`T4iZ�AUpح��>Scƭw���N�������.��0�秊-4�m�ֽ�S�c���j��+H�"��|4
��Z9�G�dGq����i�vo����\a��� 
;�
��=��{�Yy��P�Ԙ,�LҎ��/G�|�]H.�6z���s���GFs�1ߐ����n	m�x~F��������{/Ev�~��pP�Z��-���faq��)�]���Y2��*.0�X�nr<iX��-@�_O��͎�y��씎���b�HJW5�˝�/#"&���op9�{r��� !β�JK�ֲ��V^��v ۠w�tЪ5��*�:�F��H����sU٬����$���i��%�Yb@���'�:e�ȝ(�!;27��Fw�w7�Q�n�c\T�L���H�C�uK�:�5//4�:�9�zv��t�(���)�'��^T��YԳ~ox��+)ծ�X�ͱ*9����:N)���O;!f ��N�A{�kEu�w����į{䅑�Q[k6�Xhݳ��i_\̵�[��M���\'�/% � �բ��P�+��y�s�edy�����V��G)-=%�|�<)���)�j[��qo6�p3��s�<"�|HwK{/�N�Y�?���yl,tc�c�O���l��g���o�ں� #c�fec��b�copܺ��q�F�/���0�7E%9`���4_1���c��6�\+y�t�b<���7����5}�³��c�����stqf��yl�:v�ȉ2T�ǝ:��y9�{�4����d��C���1���Lj2é�-dޙ����YUҦ�[��&GK`��<,[���]�rw�;i��,s��Uu�;�%��>&�f���s.��RVk�fr[G��tٌ�=.�X=��u��]�`K�/���f�.t�*kM����3�f=�}��)�ܐ̬���\��ڣc�$2���R��҇KȚ
4��ͨ��m�{`f�z��$,QTUI��Kj6���-nZ`�2��b�--�+l1�-EE���Z�E2�[m�F��X�1
±f0Y��m��ƣ��0R�
�ffLm-q1��EF�����q�L�Y�)�.V���r�#��Ub$e�K&8�\�``�S0̮ZʔmW-jใh��5.GQ�b70��$S2�9j[�˔W(�`�mr�m�UKe�L\1�Lq1Z��(����r�LjT�e�feCj"�.X��\��V�̣�d���*��2-�G-2�e0UYZ6��Fۉ��R���=���o�W�\��0��������sدX�+�#m%����w"�Q�H�i��;3>���ZB֮=^��s^��*5ε�j��^{&r��y3~�%
�&�&�F��rrD��������A�p*�����%MC'1	��������[y��d��m�e�
-���>�\����"Ε��.�o2�fe������I��ikj���R�4���6w�7Vz�E���4�j0d�S���֌yי���mQg7�{c螌,d
5��a�켩�D��Nef�Pq��:�s��Ck�
���{�ڙ����Q���q�k�N�G�d�и��������iT�UU��i����Myr�+�E�J�����z&���5��бv�˻�>[ ݲ�4�dWSsGZ�y�\�c��^��k�C�m�t�s/�%��/�=�a���ُ���X��ې��K0�&H����6OWT��꩸��`"�0�B�Qį\f����fW��Ϻ��J�"�H�b�/_��Z�R�F��;�f���3#Nk	��Ά�	�֡I@)O�at��k��c�q���}��}𸢭�u�}¹u=bRZ��{P�tT���
�s�MK �z�h2��Z�;v����3I+�����lV`�V}�D*0�ޮ�z��/�f��B��K�Zz��P���
�X�~�h�B��7&�{�.��9i|Ro��P��??��B���Ѽm%0�+���m���á8���[C���eW���t��{�
�PN��j�8�Z���X:�s�%^��Ta�v��B��҃uqL��v����r��������9{�x�����%�ӝ��`~d�����g��yWi"�C�2c���[Ƥ/Ƙ����$U@�myhT�1X�y��vn�Bd�WmD�B�jȧb������jّ)dfzw{�׈(���S[m�%�{�))+gz�f�os�|�!��iaK�F����1s]	:5�EgOg;�q5�WCk����T:�"һ��OE�=��<3;���,���B�Z�UG�U��#�z�z�#���G��d%�Y
@��^�Su]3�-��q{�p����Zq�b� S/Q��iњ�F��"�s:�S�S�o?���� ����9M�������ԧ-�;3!s�h�:{%m���2ݨ�^��U�W��7�z�T��*_��n�I�֌Ohܭ���F��@�	_��)������������ib���I�Q�'��Τ��������Y'6��kU�K�?���l.4ܧъ*��~�5�K��iw����qʥ�LK��hw�����o/m��S�kJn�ƚ�b���0�_�q1X���w;�ͽT��oE	[1�jm�yl8�&/�q�z���}<�ጠ�f�
�W��>��Ʈ��j{��{{wW�?�Zh^�E�<�!ߨ�����\8�@�Z��kt�Y3_
d�/f�k�EKLU���d������VدW�
�I�CvK~梚�y�c���Rg��3��fWr������0����]qpOcOK�S�ݴIx����]�gĶ� ��`���;�WEAs~t�f�;�4�]3-t1�WY��u�W��s��M,�7��]��+�{����i��b4u�_�����ѡ��N:;����ض.���]� r������+	��k�S�� ���)vν96o�wW���B��xAŘ�o���a�(��U*sS���w�����C�1��í��oa���)P��)+�G��3�e��}��,8Y�[^�'(T��e�§�
b�'r����u�#�j��Ϡ�&�����2m���$g���è^�2���XU�[�6��ʝ�[��>�۾cj�6��!h0�i�:O.Z=�p�����W��l}�AƱK�F��6��D/y{��<;���d>F��Ǣ��¡b
�^0'�P��1:s����C�D�⦡w��e[Y��tWf���Y���x�棩Y<!�����;��X��}uw�h7��T���Z�1��Wވ�x�����+������|��k4�=���q�NN��	Pׅp��Z�O������/}~�UN�u(0��딶�k^<��\�x�d�7|����~J�^\`��2��V� tp/��q��:���7���lP�/�5���b��]x�CDQ|k0-U���=8�=�LE�*l_hT�yO�VR�m���c��O8T
��z��������*�xV�JD�g��s���s�F*e����^y
>��]�z����]g�x�?�S�U�U�`����>��蚍�^��ƼY������?y�Y�� �`���Z�8���ʛuR9��oM��b�а$����+�:��N���Y��t��J��7��L9���Իv�sO8�gB��U�}K!���#�aX��lU;=�~i�)ƞ?��@=��,S{����V/ؼ)e{�p���6���6����$�V�U�.�`�<���Z �
�8>���<��쫚ߤ�R� ���1�)�
�[�k`>
�\*����=�:1o�ު��� 4��K��G���W�^�C*:����s+�F��b��)�s%���4`y^�v���u6�f�\j:�b8�֮�]_���<7j �d�P���/*���3����j��REo�i5�o��d��k��3Z%��#	�.ͫ�������qoG@�Y&մ��N�B*���Ȫ�4�/�)��C��@���˺�zcmz��fR��7�E��4�
/� T�׊�Y�9��Ү�PlSSVSN�֫F�r+������k�3L���<�0��HI}��vAmv3���U�u���<6�v����0ꜜ���}�~^�V�9	B���F �� ��)o����Q{Xj���H�;0J��4l�x�.l�{-k���<4G
���QځP�~0�q�~�X+m���f�]n�]7���=mz������1ef�S^˪����A&����]g:I�e_/�>�p�s�<3o3y^�}���}%���^��nr!��ooQ�������L�|n�U	�Ԁ�V.��#ޟ*��R����wscm�Ɔ��Ea���x��p	ǖ���ٲU�Yb���]���/
�2����oD�0���J«��k�7�Ö�E�)�:�[��#�8ţ>Y���>��ZU�]1�
NP�u�Co�v�z��)m�� �}�z
%���S�yP�/s҆_�����W������}|�/n�S�u]"�լS&�C�V�W�:ȩ9����7_�=أZ�$VA�q�g��j)�4�)�䭷ٹ�5ӱX�28�]z\�Vd�(�=0h^���w{��T4p���z
xwM��N]Z9����\�����yћ��b�E��B�vy6'������ݯS�B�ك櫟
��χ�]TC�{g^�����q�Q�
w!����r�0���
��c�Ы1�{kx&H��N���HT_�K�)��i���h?1��%�/�]��i��HK�س��ǔy�^�]n�㪙�^^֟w��!�	����nލ��2.�-� ���	��&kVC��B +�:���:ݚ��5`�Ѳ��a��ū���ܟ����Y�s���m��kV�4e[Y�E�W�p�f��g��q5]ݪ냚�vY�&�,`����J;S��9�����k�ǝ�+=���	�za��l�������TX��_��vӺ��f2}��s�ƈu2u�\�%Y����]�(�룼��0��������8<(�b
/x����=�F��P!� %��qF�|�W��7��wm�+,PPYz���E7���E���z��ս�$uŚz���U�X����z\��#��[���p�u�o?"�����xpW�]�"��P�!�v����~�ތ�;�0_��E�a��ky�0�o��r6�|�|��������/+nUu~M��o&ʙ\F�f��;�3>�o�,UɡZ�=��xj�V��dM�[#��Z��6av �R(�r��.�h��Ԩ^.���a.�ۧ+��FP�YWw˫C]`�N�wӷ�=0�B�8�S�k��+�V���8�:u���@62_H�t�>��Y3��,X��ެ,��澩۵҈$⁇N�RϷ��\�޾A#Y�l��β���B��yW��1�w�Lԕ)�v-�$ͬ�n��Й��2��R읡X���i<&��*ƌ���U1S�TL�u�0,Vx��g����t��=f�Ŋ<r39��%r��&{�X+D�)�" ���X;�u%��N݉M��H��L��XT���n\��I|�KܚP����;Ԧ�5��cN��A�L	��zN��'���b��}��F�:�zv�<R�1C(���hm�۽r1Z�\Ӿ�賚�׶�(��c����S�b94��5^���ɠ�%<����H���n[O*1[���M��}��=��E]�p���bXbx(�8T��	k[��6�.��V�RD��/�sM�u,Q7ݨ"4`ذ�����B���B���}&����ah�y����J�R�˚��c��"%� Fh�z�;�m��9�����Q��ez���.k�ݬa��hG� �6rɝ*VH�9��	4���s�/o����A�g'P��cr(�1nf����z��)�7�\���-��+�� e7J���)�j9]s󹧤��ظC��뾌�r.���\s�V%3����a��/u��X��B����e�c*�l�(�³2�qZ�̦
�32�+�9��LJ̍k+(��+JQ�U���嘮*��h���˘Q��ef[�e̅X�"e�8ƋW,̘.Kl-�&.6��2(�)33"�,\����Fҵ\-��KAe�9nD����QV
���)�9f(amCP)qr8�)LnTqr�P�����cS#"�js ��\��4A��D��e����TnfEU�T.R�f`�֖�3.V�*Ȱ�s0����lbO�hhB�3^��͌(�u,m��;�+�|��i�j@�������%�;�Ϫ�9���0��p"�j�=1A_�<�x�&b�뼙ǔ���*�f�IW�b1���[��F���*�U�Ɛ}���W�a-;}�fp�έ�w]�����%����޽ d�1�@���_���WO�9��}P���B�a���k'��ה<cX|a���2�����I��._
��~ƴZJ��)ٕ�˞��kG�W��;�;o��V�p����.��ݕ��y���F����i�i��5c�n:u�����SWQ�=�=�(՛�<��l0JŅڨ]xz\��8�Y�0E�u��\CVx]��<j�p��A��}ȅC��<�˱�y,�^r���҄ �Knk�N�LҶ�,S��,΁�u񠫚��Eة��#��m+��s9r퇋��ͅ�*W�@Jsx����R�-�jp��LA��?Uzz�_EK����œè{����z�����#FLP:�\� ݪ��RE%\kM�{5�I�)�V����k@��1k��fҸ����6:!wW��ڝ/g����9���Q�
�R�nE?���8O��%��Ӹn�:	l�hc�a��F#G�\�]���
��w��[��%^yCaH�	��ܛv;��廥��'�E�Es�]��`�4:
| ( �2�?2<y��}�`P�����<�?�@�L?%2��:6�a�D\S�ʗ^��t*C	�^������h!��]�FBsӤ�� c�k!4q�]��x*wdo�W�������ZZY������awT�v4�������dq���i����9֤��Q^&��̨�ڳh��Ňt�]6�sݶ�5;O$��	|��nv�uԔ3�F~cQ�Fw�
L��6��w�t�}کW%KH�?�T h|j���嫄����E�vN�w�J�{!��=0���Ea�SjEQ���\��껶�B[�&v�Y�*��Ⴎ�Ԡ���Kݹ��=�37�za�i�,�}�XP�V�G���@.k�Q ����o��?r�Щ�SœY篅&�S����$Y�5�;+U-�-~#�B���ݒފb�hu[��9,����jT��{��(=��ʴ� 6ڰ�&�Eö�#������rr�ƢL(���q��߭����pp"�	`�پ��_�j�����g:�������(VZ.�=�d�|�L���E��A�NQ��sû����V}���u��2�f�p�w/P�^[ .��֪;���*�6���H���ڔ� �=��m6��|+�OT��"#!i��Sx�
W�䴪&+��������;脤Ry�!6����n�{t�~�dU{VS���o��r|�N��\$&��d����6�[�O*��v��@�_��s��(0�T�{|���aDՓ��O^f3u�z��:4�,�|�)T�
���)�h`�H���|%�x��%�R��J�D(X�a��S����\�w�}+/����&�(�`��f�Fʓ"R�3("���ɞ�u�֨�lQ=(>���?"��j+�糶��v�lb�p�THGl}�+�������]͘+x��׃�\��q-S&�a���B�N��.{:If�u"�o_�ag�͞���9�>|�]+�2���'e��2��q�X�8�1���*5�p8ٓ�vͶ̮Ch�=)J����<Srf;�7
n�? �	����L2e�*�p]��ŏ1�c��{F� ߭U��YFeW T�v�ʿ�+�p����y�I�:�[�T��P�Z�{��1i���C�����/�X� �GQ�I�z�O}-o5�o����Q�W���n�{qlǟ|*������F*���D:R�Z�<�W���&8��������)����!�,c\�0�j��9ݛ�({�+z�h�1G��4���\��E�.���ݽ��k�Q�ڒ%��tF���ƹhX@*��v�?I���9�1P�az����k3��׾��S�W��o��� z����0+�%ǲy5�!��4������[�Bc�����2h}�wl��7yW
�9,ԯ����u�+�^�{��,�`!�xμ�a׌�U��D��6��)X�B��{w�buײb[�0e�))K1�ĉf(M�5��,��g��5%Dt*�<�N�#�/�ۻm�C���Z����z�f
ӌ�w��ލWah׬إYʕdT�\ :�u܈�,��s���Lr�g�z�"��p�+��:�*��E^�c]����=��|��`�1x`��BڵT}�H�1�=R�FN��eH���;�CI�F�&ġ^Ϊ�k�(-1r��r$�߫��70��Պ7!B4PU�����ʊ�ھ�h�l���E���ưW��5 �Xl5��Ϫlș��ʔ}BeS�}�^XsK�UHS<�/������s��g?����7�^�h��b����bۑ�J�_jT@������-k;��tN��X-���%䉈�(Kqt�㴡5
��!P<	X,�D��]�˸��;)�[g���иh
�]=[J��I�э��m����ƺ�4�i�����^y�Θ3��}��T.�SMK�~M5���*n8�C4Q�߹�ʬ�f��4�y�W�Hme<��&�M�k�������}ط��t
2�\�k����E9tgz P+s}�'�m�w: L�C����%Pg��иѲE���"�3�_����*�yz�
=�ۄ�y�0�M2�)��#;:�z�7�H	�^9C��dǏ|���q���
�2�񂏭q,�w�7�BVy�5��Bϥ�d�ŭs����پ'��/S�!3Wޫ5�{�
�n��T�8y�S8��މ׳�!���|(�W�
n�m���7�E>$R*_���qe{�V����[+{;�L�q �Iz��>�y���5s���t�NGn&���5�>+�aS�Rg�Mʊ��%Cz��).�~�b�U�ڭfԽw�ڹΩ���s�Pmٻe�e���'�,�xӑ�MF�jm�[�I��~�� ��3�'n��Lˆ/ו���P����"��h�fU�c� -3��^t����Q�����Un��P��~Սf�z���KE�a?W�����"���)�+�w���8���DYD�g�W³E}��ݯܮ+׺������W#�Y�+u�!�JǄ%�:`>�>�Y�<���cr�z	Ra�0o�F��~(-5иj j#㶛U[�ۺ�M�-..	j�8Ґ�A��A�itj��2)��e�ڵ�	�{Q��h�a6xm^S�p(���3��;˾kk3*N}���[�U��咛=o����Ѓ�^�72�3w"�t�\ݻ5������a?bzp�R�;���X�MmG�Iܶ(��
�|��x=���WgV.�A��cSfyQE7g�w�8�wƮYǉ���{*Änd�Azj �W"�S&�$�-g�s{&Ֆ-酤k^��Q�륵h��L�^�%��нک_,:A�u�4�U$�2���K��V^���z��9�U�
W;�޶ݞFN7~����*k�P<���z��S+ʼ8N�������A����r-���ϬXL5Q��q�MH�i��$�ᣡ��w*��"�0�Y�5E����cԽ;ܵS�Y����}Y�!��T�c�ަ+,��ʘ��{V7�"�H�[N��wKn�t�
�5��S+����(D0�a�z�P�}��b&H9��rg��y�1WJ�8�Y��b��� +L0WYA������Bk7 �0����;פ�a墼Z=�[���� �X5j�"j��;#F�*����M���&��=���ީ� �����^()2,�ʼ�B��]���ލ��U��Ѽ�jj���>{M�i�z �)�/���ݼ>�����Y��vD�RE;!{���j���6�bfBƇ=�<,a��t�p�U���)ZoJ�'�[����\�9�Uи�a(Z<��1�/���-]������}�}G�[���xj�Ǐ��:��2��B��ohw�x���d��_.��	�49���jA�U]_��WyCgj��Ŵ�;s��w��M�/P����5��y��T� eu5]�k��s+C�td\$n�oWb̼�ԇ�c��_=��z�&��d�,P�<2��"+�x,�Ve�F��U6;��.I��b��1�A�K��yU��x�Z���Y]�ln� �kw�QNf��@����Z�	��Y%�I{�Z<ʡ�]�k��9��ul�CG����Fb[��3'`Xn���6�X Q�2Ŭ����64�и�JY:��"�Z!N�j��~�ҩJ�C���:Mv[,b���X�11z��k���7�ԃ�tb�b��JC�F�8Ş��]+:Ħ^�:��32�RVn'݄]��CUH���R���u*�ݘ.�&vuj����&�n�ݾ��q��u%Dݗ�m�(mu��T)�A=&[�E5���7r��We�bY��{.�U�`���cX���z�i����n�@�m�Nd��Ƴ�;��"���� �h�⻒�Ⱦ���Ql�msXp�C�aY*<Q+٨&r�d[��xa��
�Z����n��Q�d-��Փ���=R�jC*�»5M�n�2A-g�a ~V�J�n�@!h�Eq��%z�Y��#X-�K�x�h��떬~��t�ǔNŵE�9�SI�r��sS6�uݨ�o������raz�+�]�Yg��GR0!��D�0j��	��;%�����OZ3Fu3��]�0wH�Лlk׵�j@�,B՘����,���j�( �S�#�1��h��؈Rs�ѳ�s�F�#��c1&����擕�vK�t��*�t!�i����7QjJ����¯��<�|1\��z�	K���>�:#��r�~���P�%m)mˎVŶ��Z��B��3J�DE�U�1�q�h��J�&#J8�Tk`��s,�����Z�m�.4e--*��s
�Z"%ˊ�5���ٙ(��Qe�F�VA.S��d�q�Sk�rڷ2��.6eƹ[J���1�\s3%ȩlm�e
R�.e�,�Q��U�q�r�Q(�\�
���\�,�r��j�E�UB�Z�j6��V�cnZ1X�S-�1��H-2�N�d�}�ջ���q��(��e)�����/���M�2J�/�CG ��Rf�Y�A�|�]C�+Z&G=;7��\U��*�G��+(֪���D֊U9RR��EX����1�T�A��
Y�p�͢����Y�m��J�^��LT�W&�2U�%9	B�ȒaD��P�={}ݬ`��ĄiUr�����jW�'�]��gU�c�g����E�3E��^�%���A]�hǏ�/��p}�H[I�*ܴ�FF����qb��qI��y�{�$����L�h��@+��x*TȳY*q�闳������X��a���IFw���ne��9�r�:-m�_�[��P�!`k�k@�Ŗ@�D~�3sW63\�O<q�Xh���[��8���obיv���kVz]��ju�Y�WƋ�E�t�/�m�x�쮹���::��LL[��p��n�:�D¢��v#&���م�Wl՛~��FL3ڀ�jOK=�$[o/E��
��7S����{1����?o�4E?
�X���˛�];��\�\�]y��Y�/=q�Pqc��u�V�l')Q��H�
^ij���{��T��D�\4����en��<�e�wTP W���K����A�Y��f��{��6��=T���E�/H>���u�56�R��V�d���wf�7GS����L�:��I��䤠���KZJ)�{h@���|.
����Q�੟+`/{;c��=
#�h�Mt1[��f�:w��R�Y�;s]2/^��[+z>滀���zxM6Eɀ�!�;hA�苃���\V���P8U�P]MZF�pJ��X
+}�lˌ�/!X�ȯLX�(T\	�#��n�����;��FE��|�^CL���09����Y4}�9��=\�ä͋Hv���-s�Ś�W�G�����޶���N"(����Z�/�\��
1���=Ŀ_]Wf
��"q�ёf�������8�Ri�v�ǚ�3��7>xv0��h�/��SF���S8W�ABܽ�T��{;��Q��%���RI7g������ʸ�^zF��ё�4�֊�ak}X��i���]��q�3�'��=|�{N
�5� :��!����&J�Ь	��'�+�-@^*(��.�8�f`�kV)������,���t�X�q8jԓۛ�:�zB\�
�ݍO9���P�5u҅�9��F�MM���^��4��P1xI���ר�I�6M���������:��2����eve��q���[to��χفp�D��� ����i�I����*,��[�z�cTC�K>�ap�z�9T֡�ou�2��{�'������	5CN�\�B����1��~�~~~�u�fVp��/t7����C�z��zn�������IZ�c�E2�N�҅r9T35CS".<���е)7�Q��K�O�^�Jtt�����fWc�]�e��=�R�i�;�1������q��h�7���D��r�Ԑc��>�M��^�eE��1B��p�)�������sɋ����N��ݼ��mt��Z -,JژA4�p���c�ņG������#\����;5WP��m���I�㮥�ǃR/�Suv��T�E�R�ޓWEu�IY.#o�-�n����E��v0[.2�Y����z*�[�z:kv������wZ/k�ո�B��cv�(}\I!j(�z��(7��e� ������iF/���{{z62r	WӀ�|���b��9}ɡ�#Û�TƃM^�%��l��h���+E�W���Sݍ�d���o)i/W-3x9�̱�y=� I��.���kH����ݽI����hI&�d��f�ՠ��+^�Ζ�b���j�5��x��� e��O��B�	��$��٤$��(�,����æ	Ro��׳&jT����X�qD���	d�^��Pe���50!�ʕ������'z�v��e��^l-�%l�$��w��M�TiqOn8׮�ҫ35'��a� *9�,0*j٦�]��:��i��4��t��ۉdV3�.թp������\����S���� E�\�SZ�2H��D�kƆ1�z_�/ӗ�$��dZ\ukK�/�^�Z�x_3�&.B5˼xt:�.b�)4�<�e����.�hQgM�k&R�֯+�+v��Y����zM'X�u�v��m�|�q���C�q�}�T<c��P�x�.���t�7�B.�M������
[S�S��6*��Ma��3���q<�}�H�S'��N�-�q"���d��xv����`ʼ��c&=JOj�!�>�8_w3���pw/C�K\���E�F0�a'���M�7mk)\<3P4�ڬ&�mc�knhA?�c��ѯ��#��㞩����3.zݪ���q �q��8;`����M/C�����-�<1`eD��Ƹ����;�nIVL���+�";�C��w�#�cWf-�d�OM��IL^'a�B�%/7V�D؇8�K�ǈ�R�At0e�
3�M���[C�Wa��CD��MW8��F;AiH�еӈĝ�|J���/w�J4�rK�U�uOW!̦X�q�Rvw"���x	k�����tN��<ӌt�D՛��B�����k�fz��a�ei��
�;��rA���b�\U��Ǯ�$�8�Yګ���|{%J�7ğL�D��:[�2��E�v�9�G��-��Mf�:4؎�ћB�I�,o�����;�Nh��e�2�x�X�f_�A��vÁ@�u�2m���`���vvP=�`�}SQ<��㛴�:���O�����|ZNę)���oM��rZ��zc[�5���c�z{Q��cn�\⹼�;�]lX�uA���AO+�v�ɉ��A����w�7Y��3�Nb� C�`�u�� cD@����5EQ)G�w�ٮ�dn:
��U��z�ĠjsK\���g;/-j5ʡڋ
����i� ��s�nB�j��P���X�;��U�$I�̑��q�h���v�6]�|�sN5P�֭��7�:��OP9��c�s�m>|�Lluz4�u���K�6<�Uլ�[C^��NG:�7�b.�.��7P�P����f��zN�dS9�<i.�{��g�F�p���
𠊼�|��&��ow ld�A<�-��\�X�'�q���\6�o`=����t��0h{\��JzV����#��5�ˌ���NO1N�ǝ�gB�<=O�s����W	d��*:$�%���-��9���+`��4I�銆�mt��˹qЫ؅��G!ҰU���t�9��Cx��e��]+���k�k2oC'E�qݛ��hp]�fgN~j&35�{�y��P'W�[nLu�?/ma�*�ޠ���k��-�]��ա�-�� Gј�2�:%%wG���Z�����+�Z�˪�#ZnE�V�}���
��[x9n�,k����:���ȒgbΠD�>(rvu�a�驕��Cn]%a�òAI��X��f�� s�e�n���^�ZT���m���78L���(��W�����6��4��p�+�n=�K],Y�Lp.�Rp{���H����x�^|�juf̬Q^�-ӥ��g�sx�^T��Q�zƲ�C���
�Wn�DL��c��\���.�v��Ag�x���k����#��곹�E܄��:��vb�,��'N,�!-�5��O����l�S�m�Zqh��Xn������/w�c�c��န�oX�s��:eLt���q١����{kuN�k����&�a��l�jj'H���.0R�^���X���ݝ����vt)vM��L�ǥf�{9J��Buҷ����Zy+$�R���Q�"%�lLb�EP�(޼��v�����"�e����kvh�HV+�SVM(!y`#�aM�@�����3]PPn�B����\5��+�3u���ƙt���U���v �4����˦#��I4W\��;�����9������1=�4���w�nb�����n{z16���dL���P��8o��r��KS0e�aU�6y�7;v=k�t�b�
���:�j�*�n$/3R\����H���Jqh�{��z�E����~we���$��������w=
�q�����wMwY�3[Ru���]w&�%bN��a*\�c��6v�*+�V3$]��Y�1�(�>4I)J6ʥ�V媸�ūZťE���̷��jan1���)iV�U���`�4m�ԉ��p1-10�R�faU��R��2��lƥ�e-�Z#Eh��ɉUr���VۉZ�3.ZT˒�
.UR��5�33%���[�T�7%�ˍ�*#�JR�[K�r��mZ[���\r��q�#�`ࣖ�T�mq����0�-1Q��)\ʶ,I��l�G2Q�)e�p��f\i��1�R��JZ�ffWs
drեr��Pip�̴��e��s����jZf��6��3-��W�ҙ�0���H ���,:�BYݷ#U;�$�ocNBF�?@�א5��P�<�Wd=�t8t8o��9���'/���{������^��IUJDE��s��������AU���RLa]e帳�˴&��k��\���p���y8+�)�hu���Õ�U,�k�rm��ɬ���S%G������V�P��7-"w"��:{��i>,�ɨ�='y���_�ɹ�TO��.���G��)�]�S���Q{��7�5��rꠚ����0�fN��.�WGڡ�[�¶g��x�C��gСu�ҥԹWaG���,�1 �g�.E�"
�����iX�)7�nwIe�N>j7��=F)5vy*ڔ\�".P�[�n����Z�\E��l��&�f��t�#ǹ\��n�)Ȫ��F�8��!ֽ<�+�:b���a���֬���L듙��TɊj5�A��&�k�-��Y��&݋]5@��T\PR�]��X�	��s]]b�3]y�i��$�R�Xo�JR���O)�׾�h�ǉ*JK�Pd�Z�ժ�g:ݿyS���#O���лd9�HW��,�aݓ���d�'�Tlud[�� ���cj����N�KN�b}�R�s�X��V;��G�F��$�4<������37�f䃺'#s�A�q���޼�gZ`��AG�g����dY�7�F�����(��{7R3���>R�FMZ��x{�K����n6�iS�½���z1*.po�p�4T��Z�N9�vCL�ޥĜ�*�X�uq�p��׊;y�Y��HK�`�{b}���<�J��4���� �[F�*�jx��N��je:����`�Q^1��B0 �>��yܹ������:�#0ߙ��N�V���|{&]{PV�V�vV*:�ZN���;Ӽ������~E����.��V�9��n��e*���:�`j=Ǭ��U)ȂRQh��f�^B[��F�~�Nޞ۫vE���ChZ��$r�f4\��I�q�1�GM?Q�K�1�\����(�t��!��pVp�֖�wVN�,��P���Z�p6�p� �{�5�R�ۢ�&�o\�5�!3��m��� ,�xY2ǭ���=/QM�V���J�kV������N)=��[^���mU��ɪc��6v��L䈫][esYLٕ���j	�;�B�Ѷ畓kf=�TŜ�J��_f���9�q�Y]��r�a;SIR�R�\Ueۥ�pَ#�E�eǊs�=v�j�79=�Gyu�nF"�e�(LM8�xse�a�^]�z2C[6 �2ɬ���%���n��:�3B&0�7��n�
�0�}��nѶ7�/_\�e��2�AJ�X'�Ovmą~U�����[l���g�T7�A�d+g_5���>���ʛ�����&j�rK�ꫵ8���p�ȡ98x�ǧRE��_(q���o�*��qyt����J��*1�9��ް�������tJ�XU�=�<���D��Y"S�_F뎾6 �����	𩮑f�n�C�:�Qӷ%��U�*{�Fn!w�A�W�o Skb��b��<�q�Q�	�X�5�L����U�vm����(o��/�Rc����U��I��'iN���]��x��d�{{4Q+�e4�hac�4��H��cT��\�I8�l�k�K���ۉI)��!�l"��eCO8����=S��جf�n=��E�Gq��R�9��m7�mP������E�ze�*j=8;a�ճ��w����������ti7���������g$�}8����kxC��ap�i�����~}�XɁP�z<��Ƣ��ty*WWf	���[���&�C��	���5�k+�=��w{<:�Rj��5(����YފF�NI*�Z�_�F��b�`�=JIü,Y�0.2ӻ��dl�m1��\o���q����yd��U�2R��cf����^���D��}���&�^l<��*mJ-��^�ߗ��~|/,C	���M%v:c�XM�4�v��lm�ӝ��q�z�-\
�5�[�Y�-�\��J.��?z��o���Vy���(�iU�p
~��O�|�䚧-�o�2%�S�|aq9�r�9�>7K:KqU�*wڂo0Kx���}`�Y����s)ˎ+R6nN�	�/�����Y�7��j"�i�x�Me\4z\���W)��H2�Q�7��ĥn�R	_LH��>�����A�؝�v�7�Ӏ�`��V�VA��NTD��s�R��4�K��oU�V��`Eַ�]J�W�"1zw����!�,E�r��Y�U!�e���<��Q�
l�&Alw��ҵsr����^AT����r�����my����Ғ��rR���7�$�j�M�؞���&.�I���r���ZOX
�6;��p݃����~�M���n�ݕ��wSt��vԆ�/��%�}ͮ��b�*<���G|w6�M_n
uf6e�S�vڗoy��fE@^\s�3�7:�v� _u��k�&���Qu�wQ�Nm㙇�,q�Rp+���A�g�]Ae���,���S�*��=߾d.�k����2.z�4_��jT+�n�����s�∸v ���Ŗw6) ���N��9�����I�&��O��Y$���^)w�k�G WJLd�����n��yx0B���mP�j�D^�n��	d�m�<O�Oc��Z`�ya�'�p�(��(gB���j-�t}�Ub�<�g�]��aA]k(�eZ�Wx��1�洛y�z���i=�\0`S��c������9�wN��s�'�M���aMѸu�w�{�\�JU�F&밐�����L���T����͹z'_�܃8�����裇:�+O�3�&��;'��&������Jx�x@��X�b�O4��;r��"z�籜#	��{X,���C�&�Bv�W���r���`|3����RE����]��U�j���u��G����g��ӂ��z����L~�r��U�;�wq�m?��]��G�P|���xdg���r��Vr�;��֦�Z��6T��{y[R���P�c\Y�u�7����l��}�u�]��b�v��Y����Ӽ�S���.�BS4Pn	C+�0n��L��ܩ�h&�u-Q
�(?�$�P��`tp��o�in��m�T\���o����X�i����-��͡J�7��H�׺�h��l�q�,�2�蹘�󩛴�v�\%	�e�({s-\;�m.]КѴ%q6b�����|+Q�<�'ꛣ���7wD7Nmݲ�4z�ãJ%�߻��1Φ���M�4�)�vR,�C��E�͖�+�����B�h��I��'���)�HF�;��Y�Ά�����S��}�bK��#�����bU�j���_vwS�؜�J��N�K���O<��l��:�ܰ�l����:k�"�ä*���P�MF�2N�ȓ�(8�d��:�(��ub��J�I}��������2�3ngoC�9]��%q��obOI�X��w�2nv��o-ԑ�$����q��v�pۊ�q�C��'`֨�X�q܈�mK�&:u�N��4����m	{sz�!��*�[Fi'Ji5�ʾ�3���]��t�:��Rn�Y���V�A�&�]�n�9.e���I�8�9���Ŝ��ni�����Ds���P8`z���d�u�7�L�|�h��kp��^aꊑlV��ݲHo�O���e��������!4�գ�5B �*�}6�w��9����E��:Ӑ.A�¹��ɮR�aqQ=>�JG2[��ӭ�S�ivj.��{Kt�oa�2�.[W��:�;��V��+�H��EZ�|yζ�;�m҂W8�����JU�2�w����q�Y�Kee鷚�b#YP!��pC�ii�\l.U�)�+1�Y\ˍƦ-S2Q�+��#-��f-�p�`�r��R���2�\(�.�j�L��r���ū�)j����c��G)������R�e�-�n\�U���MsL)[mĹ�aZJ��tj��[s3"er�˥��*��r��2��-��]\utZ�m�me��Z���4�[b[cq[�bҹWW5f�-��2�
�-p��Z4]f[�T�\�1̹m�126+LnF�����TŲ�"�f8j�ee����*�J%���k��������5u�8֭Mfj��2�cm���dKQ�o�q�kk�T{�7��ww$����|Hg*�-K%Dsu�Z��$UjI"bD#�d3#���&*/+no-�L�2/�p��V�y5i	{�l�}�K0�s��u��v4I�dk��!�z/c��mk:*�%�%d��٭��a�,���P����B5��9�`�o��Nk���Bķ�\ʿ6��I��P5��6�:&���\^혖/^� �0߇W6�w*3�=j��
�B�b[ͼ�-^\V���d;+Iع��}�"IN�3$;q^i��o@�������CV׺�Ug-L�K�xJ��8�^����9�5yiTp�7j�ב�Z�X��oiD`��J|_���u��zx��� �O���\�K�E޵ϐ;�{��̺�pv�Y!�M����s�lb�vqh(��*Z{����rq���t�v2	<�S���tό�zb������<87o�TZ\�CJ�V$��Y�����Sm4�.�o���I0�)��`�+�D��5M�<1�'	�f.�ۭ���e��%��
��켳��8a<E��Y\���y~�٬�CA�c�e�h!�S�ӛ�����u�w��$>�(�2S�\0�����x�35��n�mJ�����6�̀P};`m�c/t�|��(�٢�Ż���2D�T��1���pѽWx�$�N�W��TLY��C��@1���RO�++ � �����Cj�E�������[{Fβq�)z���}b��m\�ʅT�Q��uY�ry�ee6�gm-IAl�1fDo�P�������
%�{Ϯ*vW{M���w�եZe��Y��͓v>�8���k�w,�|��)]���j�+������F�$A��`m��k
�H� ��u����8L����{�込�S:�I:jܭ�KF�|��1�G�|s�+=�c��RU�/T*!��2���V��7י�-�y&t�'y��Lr|�OU��i�
bx7g����r�Ul��"���5�H�bj�#�[���K�~ �I_zE7�۾̀�z6�����aǑ����@�c����+�)w��H��������U&�[3͡<��%�3��8\ۚ:)����]E�y�X�/��0n
53F�a}ZUk¼�8}<}1I���3 t"��h�D�A'	;V
�u�]\s/��r�Xdl2O>��
8Y�5�-�A.���;��n�3�Zާv���c�E}3=��ԙ��J]m�r�1>��]����9@�WtKf�y���]���á\�i�u6n��M$���qή�p~^�ji;�6�XsY�3OrX�0��k&��Ti�|�����J��������`p����U�z�]���q��B/�wN��6�-��u�F����{��O���&
�[H�r���]����-,��<38g0�A��װ�VV�Ӄ���a[{W���=Nƽ�%-��Jq�3�Z�
��6�t��>gN��ߚVa����*/.ޡ��e�Zr��X3��kX���8�$l�Ϩ��*�y���R����|�,^s�#NZ��xU�D��=���	�$ts6�ޫ�Xڱ��d/��]bn*�K�liCXJE`b����ͮ��[��"s%�M4ח�<Uz��'�O�A��Y�<z�.�Ų��1W���x:��kg����{�53Sy���]Qb)6����f�vԈ�:�i!:qF2�x��)�h�C��Edw)�;��=i�Ù��{�D3i����֟M^�i�iU�箫�u��q�5���
x�<���+Y�]w	�;���ze�@����Z�m\e���KK�
�0c{v-A�A-F��ws��md�+:����L�T�U2����At+`nt�3xl
�}�3;M�\�
��*���M�o��L�qm5�����j��rt���IN�F߫Π�9��^�j����BX�lsFO�e��pk2�1}��_���Om*�m�B� �h�pYf�o>���ѝ��C�/���㚌�Î�f�����,G�G���)$�!Ks=ۋ��en��NpLg.�Ic�E�+j�r.��쬉j��E���x�g�|���^p�꼆����m�Aғ#�e����#$镩�k�l�6̽�����9�1�/��v��o[��Eѫ��cy\�=R=�vXy�m�*��`��*�-j�u&4n|��u}��G;��R�[��)�4^�ع#2��l�w`Q�n�Щ�qG4�ux��|�����L[�N�_g��ej�Xp0I�.I$]��-��1QjV�;댬��7�M�Ī/�d������M�E�!�Q���^��wT�	�&C��&>�n��xo �gc��bN	#���F�[w��M�=t�8ά�f/�ј�~��ڃ�{wKjkc�њ��YT)c8�<9FL�J��$猒�;\N�:����W$�n�k����uf�e�P>{�5v!��G>�+���i�HǊ�8�_X9g:��nu���s�rD�*Rz>h��]���f��2�ZN�1T��,�H����Bm��AntU4�4�MdNNxI�`��f�Zj�ވ�2L���dv��Y��7'��H��^os\���[\R��=SM]a"��|���甡�=�)Z��ĉh�9�oT��Hy�٢���j�\o]��
���Bu�f����Q��7[���6`�'q��|�A.j�0�CS��ɫ�3|4�Jjy�|b�ت.�7��F�������3}V��3���j<��5������Mwz�10�����Z�s}"���\���a���M{�sׅj��̹�;$f���^�x=�������Ժ�&�� ���^N4��]at�ؓp�R�P�(��5y��+W�8�F�f*�[5s����z�o�:�����k�7f:Yé(�ંU��Pܺ���趺=��Q.$c^J?I5�y�n5��͢/���
i�.ky�ھ��w�y�eQ��	��P�����aݞ�ph�����y�;qW��כd;+[ʼL���)���T�t��&��fΒ��5G/5��j��Q�b����~gӇ�y��o���������m�qs�������`C��EOu+QAAUTB��O��!H�}�,:�H�j������0�4f3���w��=f��D�s]��t�* ����!! 	! 
@�D?�f�3n�Dذ���d=$Nҁ�P����}V@�B�{����f0 I >�"���o}����{x�������?B��7�c`���xD6�C�D8�9�qJn3�e-a��żIǶ�w����:$�$ ���q����u`H�p�@� 0d�������a����D=
���?��>��ҟ�������y��=A���>���	 !�?��������鴆!��C	!��O�	&�����a6@H=�e61$/��P��3y"{>_0{��O������\G��ŁH ����;�6�.&?��>@�$ ؟s�d�t�HlK0��z�p06��<D�i�W��sG���$ �I���d��n\hO�y�6��q��B�1��U�`��a�'��l����~�
~_�}����ڞ��a I 6��dgf@��!�7>$?�����a����'�7��	�!C�������|��o�>�����|C���z�=$�)����a��>�$������? �OV���6CO�ϴ>��-�׮BH �`}D I ?�?a?xA:c�22X����5���C�D��`��B�����!���@�p=��,I�0}���r��BBI ,6,��C�{�y6_�GzN�0�+RP>�x!;�!�M��}�bKHu8m���ӝ�$�JS�=��}�d��C���?��$��I"��z@>h��?�П��~��!���t?�z��!�!��!���#��Έ`�O�'��|g[��	�t=���Hs���	 �|��oa�}�F�������q`�� I ,�����3���A����vOYI�a�!���vC���!���~T�Ɂ1�(}g�@��� >G��z!�p|�;���������9	�ٯh��>��o�>�o�0��U�7�9��(���=^О�Ň�z8�o}ܛ����O�zCڄI I ?�#$��O�����	����������}Đ$�L�9����A�����6�;�$�06�>���lo!��A}0O�RC���!<��'��ܑN$=��v@