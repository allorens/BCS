BZh91AY&SY.���]_�`q���#� ?���bC^�  ^}�}m���m�0Q
��$���V��B�Vږ��T�[[ZH�����1(i��ڭm��`I!����T�ҫ)J&�Jԟa��eZ�UUU*6�͔�f���kCMkX�ٶ�P�Vɲ5���؋I�ړm[+4ke*��-��aM�1��4�( o�Ƿ����[j�,�UUk�mF���E��l+�MSj�30��1L���3cT�,ѭF�j���Ya�V���Ul�ն�ڦ��Y�B .�m���  Е }2z�ukX�]V�m���Z����f�ݶ�ڳ:����UwV����Ӫ�6��5ɵ�� v���ӷvhҚ�j��Ų�JT^  c�K��G.�J�ܛ� ���(���G
t���h(SM���u�i@���WGC�MS�ǙY����e�P��V�.  ����P #��

 p���� <Ӡ۴s�V� � ��a�
-�㢀�u{�  oy�� =
9�U�5&�KML�U��h2�  ����>�m#�z �x��Ҟ��[���=�Ǡ)@]z�h]�;� 
 .��  t�ѧq�� ����m����ܪGkd�֥P��6�� �  n}����oK�  ���( -I� ��^� ��=�[����ӇY�.�@iA�W�=^�@MC 5 +ή����F�+ke�6`7�  ��K�.u��@uv� wrۀ�p�:�
�X t���n�� �@��� 6�6iJ雋p U�Iقk[f6Pٛai�e�  ;;�ht�Ӳ��Ew9p
�N�X�
¬t� :�N��Ta��(nk������ٷ���.  ���V��-m�-��V�-3o   �x�'�Q�7T1AJr���:�` ��*α��WrΣ]m�u��] �� �H��eeEk&ֳV��   	�� �FҘ( v�u�h2�@t\ �N �˜ 
3AI�ݠU5v� �e�Ĳ���*�Ux  n�uCC��� �`� n�ۀ��WwZn (v�p tm��s�� 3�\�]��GO�U
P T��fU%U �@ )�4b���OPɠѣM0���T�L��EQ�р�1i�L�j��@��P       �A	'�djb�)�hz�����=5�IS�
S"2h��h4��vt;'_:��J�t�=/�4�5����7����ͱ4��\���])|Z�ɚ[\�UEs��*��QN�TTW��AQ^�����<��y���?ߏiC@�C���T��N򪠨���6<1�QQ]=����
P��L!�m	�����;m �0C��@�;`��!�؇l�`�l��v��!�48��C�!�� B`! !�v1	�� B!�q�B�hv1�6!��"&�	�C�	�C��v1C�h@�4&2;0C���Bc�� bb����6!1�8����q��1�B��b�16C�`!6�Ȇ�!��cC��48��!�b���� dv���6!1�� `4 m��� ��m��q�dvC��;؄�lC��C�� !��!�`�m	��B B B!�M���!6Lb`��!6�~C{_�-�}>J�I�W�[�b����SĦ�ť*Q�Ȭ̄L��%��"�(;v0C3e^�	��
wbXʂ����f�R�N:�֎hԶ\q�[&=ѩd6U+�X��F�PD���#�S9ù��\G3Jߨ�։��9��Ś"���G/�JUJ�ӂ�J8��rՉ�u��dCh%p�ӱ��K!�v�{*J�C�W{t�<V �>&^���!O%��	�#bV��M<ٙb2-����N6�X�Ӹd�
V����������3B����Osq�����8�������Y��l����D^�uL�%���Ju,�'$:Ȥp�E.�bc%�����5�w�;ƥ
�����c4���{���[%�5C�q#�����5]�Cm,7@�{��mH^aYM�0ɉ�HeB�����gVV9�������i�=��I�I�q�u���}���q�{��Mmc�.̶��hSjm^�.8"�0���!$�t�	�
�v�d7�p}>pT�֝f�6UG�#X%�J�jv��d"�y����4��[����PaP�V�q$q���F��0DZ���r��ecw[wu��b?[�J��A\&�QV3Cr�/ F��Fnի�j��å��ނ虆;�33󝹆MTI�]�b�	݄]��`�O%*�u�T:[��GoU���Y�trP�v�)�*��*����D=t�G�#|~ٶJ��s��h���b�9[1�Um��0l̟]��fE��w;��B.��$�N �J��WssJ��[�1�F3U��2�*�!�4����n;�MSB���Z�lDZTHY9��=ڃQX$%�A 0q��F�Gwb�!�p�]Ha:LX�~�be�d��mMQUQe㺪�]Cz(3�%Sմ֧i��c��֌O#�:b�T�<͑����F��k���p���;a����S�����V�C����f^QY��q+4�JGLT9�UXI�惢������sŘ����鑷��5�bA�:4h�z-��Y0����ը՜Mo�ڽݳ�5����(6V�sk0dt�[ae��,��-��
;j�M�`�D�PC	��\�cnA��"�ܱY�����ѳ ��pfTUY��5�ADke�q뵕�jg�"7���r�ʁ@DNcج�滽+*-�!�i̭vB�ш�QL�*P��KR8/IW 6f�&bc(ҎùB��72��H15(^�2��X���U�*w�t�JΙDf�K�`���a���p��0�/ʮ��ڇI°s���Ԛޒ�ʧ�D
�wX�����%���f�h^^�j��r�9t��.�,��tf��O���vP2Y�ZZ{��]�jޗb̵	r���65UOe�����b/e��Z#��͂�9V�t��{��/V����;2��y�/+�iǺ$�I�ſ$�)ݳl��ݖT�(mi�Ot�	��UVb����W�i�1,Ւ�(m&�w�/��@Đ�Q��܆�LG���Y.&����U&\�q���r��X71Ʉ��Dd�Pi��U/A�$l�d�J��6��Ar�j�3e5V����Cq��T�ZN�31�.D1YA�
��D�&9{j����0U/6	U�թ�4�0�rj��r���Rmh�u��-
RT�K���sS
4rY���6٧��D�ڇF��LZr�	
�3��[����Q��J
�m��	�CRU��/5�,�v1U�u�.��6��rԗ/K�vR�W�*�Upb:h�C��[H�bfM{5b������,���%��JT��@��MfT�U�6�Ci���k�������Ov��܂i�<�U�-n���e�t�2�P٭�8�����̷x�G� ��77m�<��]�@c�q���Z�m��%�M��_t���X=������o]��ݹX���y�޵?4!u���qBS!_���WB5���5o/��ȹ�Qɑ��U��ttR�;ܰMNM�0:x5"j��q�;��[��6V�w
<;^�Wn٫�1P "��O��o۽L�d��М5g�A�i��ւ�mWĔ�E�j�&��b�㰃�#$Н��j;���]V�v�`�/�e�������`�~r���P�� ����� �0�-9�*�F2�\���卩����t�d���UA*��3�Z&�Ȟś(���r��7�^LN��E��e�^¯3�e�'qY�l���Tp�58)������c6��bl�ZkB���r�.�8����Q:ơ6�fX�����X�d��a���]�a1˅�v���]��
^U���䛱�ҷ$�V1PTCȷq�+ڙ��{�4�P�z)�1�Ɲ���Ս�1�F� �Lvh()�z�]��N<Z�}������A�dxp;�e�odn�I-���5`���D�f���+6Ea��)3�m���'E �*�-�����N$���H�٪*��6�k4���3d:0[�Q�Zw�X�zې�F�5�F,c1
צ�f���EeXNZ/u�xkNBbas`�Zr
�F����W1v2�u�
o�[ ��'cN�B�����t�i��͂St��+ޫ\^6;����w��=�B�kČ8#�/v�⡉S5�kl^�L&(�@�̧y%�VIV4�*�]u�����O���ΚZeB�6۷�d'#�u���)H�Ơ��7i��l�4�Yq	gvi��Jʲ5#d�BԓAܚ��G)�ʹu2�������Io����O(%C���;�ي�CF��p�&�!�;vM�*mꬸm="<�e�U,�ǭ��hWY�i��x!�oDZ���3���̩Z���0b��s\��n��k�Yko���Z�o]�VY�CVu�M�yG����I�ٮ��3�&D��L)W�2]f�é%�C&WD��y��mX��B�ܗ����3���4m�_�ʘp1�l�Y	e��Sriѥ"�²`5� V��Us	t^U��9SC˖�١��X�f^���{V����c�2�S+3.�Y�KƲ��H�8n�f��V�A��5�_r����a����,��l�x�Ǔ�Q�@��pG0�[��#�+��Y�{�F�ʹ3.��˕�nn�f�z���ͼX�JML�J�K>��rS.�3���Ն�f��/^��tc�ю�e�r����T���DSH��V�ʗ
n�jý��U�a�����9��Pܬ�顁�{�"��������l�)M�MmV��/6�kx�3u�ܛ�M�bպ*ܐ�`��WN2�%�,��j��yH�I�7��P%�6�ѹ�zC���Ŋz�v�d�W�`��+7l�U���1���y�Fm�9vk��Suf�
�UN_wvȥ��c-,�w[b�I����|��]���{�đ:Igi%$�Y݂EXsX7X%mV݇uNR'I]������!z�������a�ٸ�����n���iD��h����1�Un�Qn�a-�z�wS5v�[�~��!��-S�ƃ�mO�fnd����tU!�㫣��`�Nƫ�Zڔsi�\f�2:�IY�>UHM;���D5oj(�U�A�a�v��1� ��ɬ��Q��X2��`l��J*��.�*�̬ѐHT�����ؔyR�:a�+R��&��Y���չ��׎��*kB�����x���5%8Q�#��K񫌆��Ef����ŏa6����܁���'n��w�l��ø�!uE�8u�-mY���F�	�%�k�3/,'Lّ㙉Xyը��ƍ,^�O�݈�	Ӻtu.�
���u.),���%�!�E�$ә����B�W��)7�T�lúU�L�J�77vc:��6��]2- ��B�|[�,1��ђۡ�5M���	//۴2�,FME�����&��:ݰ@{]���qq���<���f��u�5͡Rf�#3$�+s ���GU6p�'.��VEGK�&愖��X�-��B���yl��JYN}M�aW����m��)�{�D^^A�F�0ٶ�Zљ�S�.��)y�dj�,R��֦�o\�j�9��O(K�qͽh�ǯ��^Qf���sm�BDZ���MXE�L����Y�w��!�J%V�E��l0�H-[V�V'��en��s�D�d��i[��6՛��b���s6�#eg.���g�36�Fj���ۢp���HZm�/ȑBX9*��7wG1�[�a��f�q�f�ؙq�G7�U{�j�-����e�#��*^���y�<i�z��7&٘Rڽj71�ٺ��فf���#{0M��փ{���k]�u�iӵ��=U�b��I�v:Q����
MZ�}��V�2�K�<-!������^�dg5]��dcmrAW��@��*�V6i�L׬�,K[���y�obR=��t(�'�n����a��Tr�%e�tZY�v�4�)U�UGi���(;?n��m��ݼ���`a@a�	$��r,���u�QEr�܋w7[��0�yo2(��dU9nL�Uۓ�=��
�-�FmI��7z4��P���n�A5����yP�X�^�˕��X��0��r�,�M	���'��]YoSuc��z�4]�x:��MYX��Δ�\�z�*�ܖq�S6��rM�}�.��K(�i����:b,Xծ���N���s*�k���U�t����Bn�%�� y�M��h�;��h��K�0mSh��	:,|�̵E��֫H��Έ�I�w�+h�ot� 9{�-r�&�@�mX��0�9zv�fh&ܔ�|�Rv���+�kE�ZY9G���g`"f7n]�6�%���u&�8��'�ޱ�}حbAӾ���6��<Zv�	[0&�4�\n�7i�,�x��mL�F� �};�٭y�=���w��*c���̽�n�fn�;xh�+�A�^��o�l��>��`��$�܅i���&K�\Ȯ�C��ً���iG˗�j�W�bb����^�ձF�v)�m����)dw��r�g9\���H'�ҰWk�9��\5���S[�;�+��y���/Hz��qcy�:�� ��T�T�4�R���+ʺ#@�g1�X&�v�Y��w5O�����U����i���a����ͭUd|i%��ͳ܈z$.c@SSuXn[l�ee�.䊴�+f���K��O49���w[T�GLP���@r�X�+E��9M3V���V)���B.�.������T�Z�e�kE��6�%/�f�"�Q9�*"r�m��*VK�[�9*��_V��V潋$�30��v'N�u�l�u/��L��F���WB��C�k3$kX8̴�KF���f:��V���l(M���,��3�[y6r�t$sUʀͣ.Ū{q�����h���SR7)6��eTˎV	�� ��:,�;g5%�D��{Dn�5�5��B��m*�M]�KwA����&�0��V�rmZ�`�$Pf�
nC)�Yj�Y���2E��e��Lr����ފ�VL�+NZ�[B��#�(:pY�N5�X�a�ٮN�Hk���S�*�����/��]:WX�ҵ��ݦ�;h�"6nQ�	:ᄢ�ުm��.�f�t��jQ,�JؚUc�#++v!x%��-��Y��u��	��A���Ǝ
�"Zj�E72K2�8v�S�s�(��4s�v�&��gK�.cG&���-R}v���-ލ��w�7-��e;I�Va�J*�Y-���,p�J��ص�i���n]LƨnMa'u�J�Tܗ�U*�1w$��K7&<��&��&������� �]h��7A�Ƙ,���s��á���Z��m��C��˥V~<�@�7�LԨX���:$`�g^�E�}\���j���p	f�t�#R���sJݬ��K-sRR�\�HE�P�&R�ݲ�M_X��\G�ᄠHŌ�9K��E��鬲�#x)'�$k3b�D�=��j�^b���ԪVI?d&��H��$E͖��VἕV�pU�zflbb7�l7j8��oVW��æm���/,�ؤj�Z���mձ���d�c�[h�Q)�#M]��I���R4]�-�J^Ml�UX*���*�5!����Y/~&6��k�DB�*�ʰ��!fQ�k�a*�{�vc,	��{�l� WCb�#0&G�E9F���Ʊ:�j̴��4��MR�S1l�/,�q=D<��_n_e"��Ύ����=����hi�F6�h�Z+ß�f�sjM[�ͼ���T�c{���Ա�C��	�i�l�OV�i��I�VӲ��p�e:�n��^���#Պ*��HQ�n�	z@x��Av��k��wMQ)�4��L�X����r�l�y�Q��yI^*Jef�W{�+FA�.H%���I�2!�t�ǓfL9�^��-ws]j"�̊����EL5/iT˃����IUmY�-�I��6�x*��Skh�Gp��zv����TSbDq���f�R�Y�&'KZ܂��#��8��#�m�:��iԶVM�6c�-x�Q��E�ksveI3i��^KS,��­�s��1։T�U2ea�&��"�(�vl'#�5.\
�:2i��6"�^cyZ�����Q_i5b1�*
�Y��8l�72��ӄ�&�;x[r�Uc�%nDZbl�N��Z��B��4UfЊ%��{���Lc�B��g�S-���y��Qg��$A������=��;�J�ERR��V��7��%�
��M�k`������m)��Y7f޽�V��r'i�����J�N.J�����ę2�q�6B1�շ�8j���%�m����t2���Z�T�O���t�,�A-�fn�blD�6���ҮY6p^)1�o��mH��(�C6X)6�N��e�%��}���mL�pZo��)iY�V,'��v��*i�.���_2����r�����7�m����w�E܏v.X,���lܖpJ�@�ƥD����a���!w��&`5�'�܍�D�&,rJ�U��)!��k���igt�}����/$#b��މ���?�z����o��,��?�uun+�gu��Y����9��IVu֩�
l�E%��@��X��u�a*��%�)���vM��P�B�ە�ͫ��*����w���/��D��]S�&�����k�{�z�x����wl��E�2�h�M[3z��a�@KʗՃ��n]��9�H���V��+������M�$���TRx��ӢJ����!��&C��Z�X	�J�=L۰H�����W�*W;�Eɬ�S`hvWD�:���o�6�My��J�m�E+Q�F:�5��n]n����l2P�#�:��O� �\ݵ����ϰ���mM��;�]}X��Z����:��.]�h�)�'Yɣ��=|7/1�c1QS� 6}���J��F�q�̈́f��%o|�.*�4ݴ���)\�X�8,�9�a���hMTzP[�M�Hs�­�!\�1��U�Ϻ��Vm��"�"�ݷ+eAnu���c��M�y�O�N��*���[�q#�����z��P�ڹ�*C�����;Eb�k���{!w[ړU��blZF ˹geR.<.ۺ�f}ʡ0�cy�(i��XM
u��s:��%ܸz2E1#ۼ�5ٸX���$����ܷ�3�Z҄���p�z��:I��)ܻ�q*R�\�ensE@վ��㥪ږ_hޤv���8���]]d�[ܻ��R�/�����3��:lݘ�nG5�4\�}�>�f���y��$G��բ�U�U�Ug��й�$5��b�`6��C�:�rL{��W��orɹt�$�h����D}�؛!��;�o���_e%�~�䃤����b�-���CfN��f���+��G,�F��w�{�k5�z�]+��*:�P�"��U��!r�Ai[�܇�d޹[��m�E���f�	X��ͱ��{G!�7���Ll�_�t]K��P�0��n)�u�1����ohS�gJ��̹���Ÿ10��.�;��;�rktQ��hv�yj��ރL�P7]Pe<p-T��[��%��A�@2棖#�!2<gp�\�mS9܊֊v���������8'Q�~T�SږHc �v��ˮbn1�w��fU"!<;�����\��XN�#aM���W��R���o��.�=S�9
�w��)m9�s�1}k�bڭ���f>�b�2�M��X).�����͖�/�|mu��bٕ����O�;o��+��O�Rң�oOr]�ji�Y:*��mlM�u�jDj�j�oig(a�*�K�M�v\�v �)�����J�>"'U)�6����C�2��5�}���:3�K���40��G�ŖȥF�P�(=�Ji�B��Z�Z��(�1)�T�&��4"��Ș�4���`��6m�I���՟�d��)�G`z��*�0��h7��݌q����|��Tǘ\Y�Yݝ.�a3:��Ӻ�=�2���BYˇ6�+�&�#���Gn���
�k��A��YEٲ��ݾz�Εs�~U��jF��QtF
��r�lZ0Yר�����N�(��N��x��GEq������S�d���܊1>2��~s&f��YNJc6��ᮍe9���5(��ߒ��C��Xw��|�2GR� ��7[ڙ��ք��i�x�C2�`��XΔFh�Xn�$)��q��o�\��j�F�W�`]�pY��z�t1�+�]Y�k�ҁ݉��R�q��LJn�������q����;��p����P����qu���+YG,i�Q�v���L�2M�������S��f��ՊԚ���[Αv��[��0gd��a�ٽY��JU�����qR"f%ege�ʔ+j�ï��R����n�����ks��]�I��ʪ�Mt��ZK̪�n�p�i+�k��e�Z�^��s1mC�n���.���+RŚ6���aR�`Lp����ј��P�u�rwo'J_f��x%_Ӊ�\��-�+Yfe�FPOOZ��Ju�,�CMʽ-�d�w@�,x7�rU�K�����%W�OzK톱�p�n��w,B�w^�l�x����-ꏦ\w9�G�\�7[]��篺�$)\���\��jS�w]�W-�D�^�L
eE�SE㩀󻚦v!u��V�����+t8�yfQ�6��q7+Q�ַ�Z��ճp��Wݶ]��ب��[p��jmi_w.t���PX�ҳ�D���^}���������!T���OKk--��VSP4b�-ڎ �vgJ��TsbM��g�X�����#J����]�i��3�x̬��e}x�r����.8���ב#ܞbA^�LrGE՜�h����I��3\�,UX�^n�{M�u�h\�P�M�]�pK��k���b,Ж����ܧB��^	��66�,�A%CP�n����Q�l��WM����&v|'�q�S6��x2�)au)(z�E�h�r�e��3uВ���U��w�k��e��uQ+���(�T"���uhݷ;�e�t���7� �Qػ*�v�n�G�����H1ҝ���V��������B�p��%�wSN�{Ʊx&�v[��U�KI{�l��s�q�0G:��ױ$��fí��j��^��b��V�ɽY:�ys&��o����Њ�ˬ>tv���路e�Z�3�,�*�̤�ڀ��n`�\ˏ��{ŰU�kmCl~���5��l�F&�v�F��օ-O�)��i*l�5�ǔ:�vԻ�A�2B��2J�D^�n'ƍ�e��x�-Q�8�[�8��%*�L
�@-�9ޘ��~Ya�6M�ABi�n�FȆR��yʹ+s4@hr������`�^
�l[�ܙ)@^v��ZSK�Ԧ�1�Q�B�>�J���w��w,P.�@Pgx��ם ����)�8��N���]:c��3�A�nj�}��	�v�p�o���{�z�k5f��VKM�(Y��h�43[}DQ�]�Tiw8ԣ���7��W��]Xvk�������20�K 79pH�%��4�k��5�Q�.�Bt��FB��̽XB�7ZZ]�s�k6���<S;/�YH`ë�ގ����oݮ���ٜq�ճ�<ګ�w�ٵIW8�w�lNv��p}�����cj���*��l5_�l��p����xU��T�lK��nLZ)VL��i��u�&s��oj�vw��Z���YY6��5����S�T���9��&J��yY��U���Z5{0�r���I1�����e-�j�ۇ�Q��h#��S��s�F�A�/����F�ty���˳@��"����3^�\��yg�/���M���K�{Ù�DH�$il[��v�Q�œ�ݻ��n�[�Od�mk�Z��v�����MGfP ��\�|I���{��޼���m=��U�lӧ�J�ݞ�evqsiY6���y҅mr��N���:�1V����,�ͣ���Ȧ�
H౾��������O]����]g���z�Α�5U�I"������g�''}��x�Ox6����B<�Bod�.�v��>�ѝ���snز�p	��aug��&T�c�ѥ���'�����d�-�v�x�׏�.�6�#+NǛ��,*Y�v`:+FH�ɼ�q�E�����c�m� �	��ges� s�j�Ц�]&����zX���녮�.f�-.#�E`:��U�x�,��Xfmo��R���WS�c�����A&I�?��)�4&q������FM�[�=4�71CC�U�n�r�V+��h`�Y�B�P��c�ᄖ��s=^cڐ�/x��3�9oRn�h���p�;g��.j8򞳭ϫ>�Xv[����Y��l꬚&Pf=7����e�S�'!�9��GC�˳3��#�ff[��uU�_�g*�}IZ�Ǩ�����[����
W�V'N	u�1��A ��\��ӵy{b5r�q�UpޑhΑ���k{ub� �](����31����.G6%Z�|�j�/�yJ����ܳ�L�ÖJ�q�h�(p�=O�X;�tQ�M�����mT�:+�����<�[���VaEq#I¥����=�lr�p�r�s��':Nn���C��t���
Ka�y��f�Ri-��en�{�K��f�r7���;Xh7��s��S�<S͂���
�;���\�)�;9�9�
�����킵�ʨ�"6V�E1+:�ڮ�X����4�vXZ_9�]k/L�g��(api�j�[UbbǓw) �*��i�0]:��(�s�}��s��ySn ���M��m��a[*��̪��Y�.q�y\��ej�Νnv<�V���f�����]�-1��]M@8�ң��I=�e�F���n�S��r�F�ϯLKkP�\�afd��i�;�A�,��ϙ\L|��f�n\�%�ss.��Cf��\u�H�8��gS�4�ӱ.�$�����u�i��WDjX������3\���s''v����T\by0��Eb,�Kn�U��њu�z�����[�2����M�ӶN�嗏��V�u�Vc짹5�Y�O4�[-�\)�u������>�[�Z0���v�ݢ��VwC0	<�J��͢��O���꽠���JTq_�y�S��Hs��³{d�bR̔���Zʧ���oH��_!y�c�M�4i�4a_Z�l��K�5i����=mJ�2�f���/
!��t:��f��p�Qn��M�]k-G\��Ҝ���w�mf��]��%ݮ���SUA%r'rħ"�њqh���x�'����nr�o!��S!�:�N�U���0�ǵ����r?C�E>�7��~���+��n�N�y�����Z/U��<#D�}p���V�n�&���6�:: �7c�O\͖��w�.��w�z��MԽc\�fC���.��u&��*3�c��E��5�k�7V�+�=����H�yݘZ�l�Җ"�ݙܴK�[j�N��F @�j��Z���.�ܭ}H�Ι�]FT��{�N��{�L��<浔�\y7�r;�g]�ȭd
k��W���%h��n;�1���Β͌yP�/C��z�rh��ש��uC֪��bz��& �\���j���{��7a���͆�in�һ���GI�t�k���2!&_`��á�3����S,��S�(i�.U�����l�'�5�u����:Hz`Ƶ���1g^2;u��H@۵��:�w,�c����^��F�:�v�S�KB�u-֚���F�y��G���rЈLݩ��%T���	[�������ܜ3�zp�Յ5��#.K�݌a�����}c`��l6f���� �r,\Y���Z��m�=Wh5m�5{%�^I��}�xɣ��@�]���T�\3��3�GU.h��򗵙�d�Mi7���`�x>ª:���v>7��]��F�lv6��rK�DT'*͢�N���vH��m��feY�l��Ofչ�2d/�UY���~�FN�Y�R�q�e.R*U�P9Q7���u}b��������_Ƕ�v�4���$�q��R�(o�^�f�m3QS��*�aسo��ՒҬ;�k����E�Y�{�I��j��KB=�`,̋y�;"l䲮�|��I�yj�v1|�e���g��������e���b���hK��fj���B�ۮ��e�^K�ޠ�#5��	;�[#z�mM����·+Lu�׬˭#�h��)�{�w'�ƀ�c6���8yu2薦=Q�B����֘h�֊�1����4mgr@�
���lC���1��� �&�⎦	v�n�uj�ä[�۰~�e�������oCy�>�͘f�y�Vjܣdg������	�ݤ�a��T�w����5kT�F	;A�����>��i���V�k��T/s2�����J��9��,�-���VN������S9�����u�e��te�D[�!��f֜�u��Z����̶r��w4&��[��*�Hh#�J���<W�BE�iS�(;ܜn,��:���,J�2�n���5�_>%�Z�g�^�\X.�c��e�X�6����CTV,��9L�G���5%0
�GZ�.ӣ�3�����c��_3��3/x>��p���J{J��O	u��.��eu�ut'
W��L1.iŋ2���B���H��?g2�%t�mm�ܘ��/�Krkᷯif���Ѫ(2#Fm���}�୥�f�mY�G��m�]�ܴ`#��	���߰d�ŭ�fM��+��x����lS��%HJj��$�ꭕy/<݊q'���-�UUT�X���.^�qSin=R��N��x�v���\���
����\$ջs��ՃF�Ma��q4"��nR�>�1`��+�E���W2ƽ�l�^�.��J\�n#����������8[���w*ힴ��/�=\�Q{Hf�iec��42>�����K�EgKc�䣚Wk	Yk)�1Rt)m��r��[�ȡ�/Eϔ���[v����'b��[���_�A7���Ѷ)���J��U�ģ�z`���� \�h�oD�#&r���m[æ��LX�A屵�>�p7յ�޵�����w�㝩��`@������/M��f�r���ꋓ!J�; K�umi�ql�mu-���Fk�z�F�&�_{r��vQ�ÖNM ��X]�Ԗ9�2Į�&��2Vd���=�18�lR��f>�..����v˜Y�jqr [ñ뉌�����2�V�T�鐗�CL�{��r�f蚩��*ZQx&B��l��%ݹ��:��z�$L0Q�`b�sn�v�=����
���b��x��}W57)�T�s�.;����zJ��>�6�*?�!���?���$���	%������߫��ǖ����OڹC�}�?�~?���?
f@�~L.=��me/�"��&$p�ҥ��Ä�ai�+kiKB��)H�=�
�+����A@ 2�[�_�3�n(�
�����\�t���W���ǒ�c5���-jkz�J�Z�����e�L1.��\ԣ���C\�L�n��R3v�̡}!�M*��]	�8u��^I�,����[��=�x��fdE��{���-V��ܱ�S�;8١9�A���Jq�q����qӓ�g)�;t�+t*h?f��u0J%��V��r �fe�*����ϖ��lvK=�a�{���/;#�9
�u��)8vcl;�:3j���f=����+)䬒��el��՝�m�ĥ�
�h
�h�z����\x^<��X��G��g9�u�h�`8�G��dt�|���ii����Ӯ�=��b��V��I���u�/4��L��ñ���PȘ�-me`����tu�wesE����(HOm��<��2�n�]�y���9g+������c�+NU��Sc�'Z[*�k(�we-�ܴb5�`�2v����yե�mE�w�hZ-:�!���]s���7T�GE���<:j����q}ʊ9}��x[�d=������Ɇ�6�9�z�p쾣V;]��4������\a0�\,�
�W;�����]�-yϦ�o�IT�V�/.J����d60����k����b���=���]3ˮ㎦�%35���Sk`�sd���V��-�3.�-����jLcj�r���;y��*�]nMځ���"ѕ�rN[q�W;�I#3�7��}��v�/�ta���3�J�naĢ1��/� �8h�C�8AÇ(p��8!Çp8p �8p�Â8p�Å�8pc�8p��#d��>�N������^X7a�T{uA�2;^���"1M)d8�EuӢm����*�Rӽ��Q�ջ@�5�/��vM[�x��U��1�7}&�V�[1-�iF�R4�m�AӃ�h�#�U�y��ֱ�*GrӾ��2��Bf��3^kz��&�U�n�R�`�T�ڛ�h��f�$��wM��!2�NA�Di?�aް�u=��I�GI�\�o۬:�V���1�Z]X9GGR�f��ƣ]��[w/PVV)�&��������5�;(0렘0��.�GNBH�7�,O��������iܮ܈l��.^|E죦L��h����֩�&;��5�q譛��"�z�m���Ӕ��t� �.�Ǒ�̓�+͉�%^�c��<��,H6
!�Mx^���ǖ�U]��9(5f��/`=|��xUf�⥗�왽�1�c���W�:~�֊E�t)��;���\:�D�0�
Y�ڣ�,X�Q���[�ju�X�Mh�m��Ϧ�;,Ҷ��N�)��v<��[ںت�Z�\�Zw|�8.�n���1�;���P˕���h�yQm��o����A[�v��v_R�ӡk38J�:W.���S���Ң�Z�R�2Y�����QdzQ�po'w����4����W,م'՗o*Ѿ۱%�Cx+Q�����W�5CZjj"�Y�������<88p�Ç88p�Ä8pC�a�88p�Ç8Ç8p���U�3*S�GӣD���j�\���L�X8kL[QG��Z.�P��;����(Q=�V�(S�jYm[�XM2둚l�h���Z� J���J��c���3(fؚxhAXέ0�n�ưSat�9̫�b!��[��62+ü��x�P�w&��=]@_�R��ٶ�����=7���۳tr!6�Y�)��wc	�I���Dj����[k��P��晀Ø���UR�Z�r�GɈn�En����0�U��흵��X��f�v(Ss���ҳnP3[t���/a���d[nv��tn�ϦTՁ��`U�,G�D�v!0��f��xJ2�P�ٛ]���O�1��on�Z/����\4J�p���m�i�{�԰*ӳW[V�r�6�*총䎆�玨≠���-��v��*���{M�c]-�,���U0��*��.�.Z�&s��t6�a�������=��kr��]���<���gA�ʄ��Ǐ�ޤ39<�c/��2�Mޱx�t��6��z�֋s�6��.�6rF��S,��@�����Z��/[2�z�K)�i�Q�^����vYN�|��O��W:�U[��j�ڡ��4�K��c)#���7ϫ����PS��㊑�m��܁wIT`c���+K����W�*�7�� ����h��T�0V"�ɀ��̈́��!s:�n���H�Wӂ�Z�Mb�ںw�:G5��<�k-cV�YHV�̓v�WrTe�K:e5�.a*�D�Ds���=��������s׵�吡��X�97{9$��Ϋ0 ��:lw�	�8�7��_�Q+���k:�Nܴ\�b�!��S��v;]ڳ���lZ�����J2�b���c@�:2�:�����[�9u�x�7rC3��77E��D"R�Q#0U�CqmA��+7��?\V�Yګw�v	�Ǔ�Ǵ mܝ�K�`���n��5sd0hpl)�m��UG�TUE�4�;^�B��޷-�)�w�[�t�ԞC�b�`Xf��3$6��T���ެXw���U�����g��rbW��"�w��M ���x,��"Na�����Ğb.�l�ʛ�fdր�L=�c�K��ǯ��u)a�{�A��ų�h�j<���/��b�]K�S�:2��ĮI<H}(��Ď�U/ λ�T�s9ӫ���H�����}�VT<���YCo�/�ww)�Z�sB� �C�jH�(ݐH����'C�J��oh]���V�.�;&����O9���IxsA�	�u��}+X��E#Օ����O'g���ӽ��ۣ��s�O�c�(��L#w� �ͦ�P��3}�&7!�r�7L�wf�k:뜨�#���O�J��$�钕ҁ�����M��mz�;����m��=$�#h3��c��yt�p3%eSd��=�������b��o-��olZmJ�!KA����.�n1ԃ#SaUu�Y�'Z�kk$�u�T�͹k�����7zJ�o�P��ˢBTAV�������r鎝��`;%`д؉aF�Û��o['�Ƒ�r�};j�Z�R�ss&����QⲭMI'���5��7N��;����+[ToK\w���y��N+��B.9A3rsw���3w.�)(�o9mn���E�j�[}�|�T4��Tef����i��v�mg*��n�L})V��jr��m�:������ؕ�"9��Bk[y1*uu�i��k��f�ѧ�V��wf։�^Hf�MKw\z��ԍ���|�^u�	��\�u@��s[0V^.�ꪴu��{�Q�ÓPz�h�R"E�Z]K��j#W�w��Fnk�	���� �x��Ι�`�}�v�#��
.���踷5���N\���B��)D�Ӯ��#�� �AZ�C�XN:,FL�� �1Rf�L��"��V�u�\�p�zP�8�76�n��
j��|V��,N�!��ۯ{ky|�v�Ӻذ��O�U��fX�#�(ܒ����W�\�'q�'i�sK>�J�C_%5�3��ۣ..���7�_`6q#�]�R� :��+��3׻b�H���&bFĒ�j6��3�3r͘�����b|�,�Gy6�}L�:�f��.�8V��'�޴��^ZZ������;j�����Xt��������Ի{�����<5���WN�9V��F�v�Y�:Y�X��Ef�1�[B��4sP�Kr���`���.6վ7�ݱ�k�.�٫��4���WR�R���іӂ�O��|u^d�gG`�����2՛i�:�P���ÍB�mV����	CJ� h$�b�����i������ԥZ��I�P��՝$\^`��Ԯ�鵮
��ủ�B������SU���6.��Xm�E���&�Nm��-�B�0����>�j��pU
E�"���r�<c���x(g�����e9�Vkx�����mkt\
�����m:�b.����⣪�/�(��{��;N���a���zZL����}oH����v��X�Nk;�Y����5��Ir��	����GbFL��Q��IWQ���Xi�<���-Y|]���YJ]чV��FvvjJ��Y��(+��VS���=��F�i��̊F���ΕwZ�1K�O$f�H�e�sM6�k�;@�B"M�~���O��g+_2� /n�W)���٘�IX�ػ`� �Zˑ�V]��r�+��F�#���ڋM�t6��,�h��oz���+�յ;�F���-T/�{J:Tb�w��kT�ܡ��ˣ������h��;�#ݭ蓽
�+Wۭ���u����0q��^4�H��f��^2��ӡ�EG�]N^�c8Du7wʆ����X��d�"�j�[_rKd5�ta���7.��Z��d���p稛�ꨆ��fә�1�c5�\��5�[�h���gԮ&:�uS����:���iX�A�+��E��z�������5$�����l�:�F,�y�,vDѺ��U��-:���R�$8�g�5��ވ��#y!�
HX\{�1r8;U빣�����El犣7٪���Pȩ�["���K�ں�L'Md'�h��Q�ڬ%9�9���W��ȫטA6�e��|��M�m��Z��Hؽ՝���Z�wZG�SK7WYr��&K|�,��������~��[�i�a(��|&hoF�7FM��"oVR&]�߶�M}uc#v+�!�'^�"��V��j�i\�|��V�r��f�GwOd�=�#&(31�8�Z�����ڴ �eđ�����ٻ��Lo�	H����I��d���;o���vZ�;vEG2�mՁkR�rF�J~�����Y�����/������r������j�Y3��.sIX�U8	�)�`Z.C �"�Ҫ��_v�1:��v-hV.@�Y��
F1X��{b�)���9^*Ր��	F�
�a�bi��9��A��+�/9Y�(#En�'��t�Rɘ����e�0�Ƹ��t������E��X��Z-�*
�u���v�q���5��f�2��w�Ϊ�K���o6��V�0͵�u��/�yg����r�F��4n�nbo�4�5�pQ<����<*i���t�wQ̺��l��,��(l�r��an�}Kr�=1CR[-����y�����"և�R7������={	��$��*�v�rIb�V#ӾӼ�;�̷;�B4R:�uw�\���{������t�s���3��6�j-����2�과���Swm�fsݿj�}|Ӻ"�J}5�;�n�rn
�E���tn_�JO�m�����qFt�,�pN�$;��� U��'���:�"��J��:}�����"���鸝q��w�(��R�Y!�1�F�v�b�G�[T�����ݭI.�2��t/h���&`�W.v�;��K�\�{p܍I�~�.��������NñsrtD��r��s;��:�ƽ�W51��N̟+���悷:ݒȳ����t�S����g�{&�|s�:�m
7��u��P�V����}G��ie���G��B�9�J+8'Qe��Ni�w��x~�C��F�D��o�e#zέ,MM썛E��W^��F5x�v�Ų�hŎ]�u���[�v;�("Te�좏t�޸7s�43�K5N�z*��Wtm�sha�s�u|j�Q9T�g�����5��0�Rӫ�*��	P۳��6j�"]A��E���Y��d�W��6��5	p"n���L�u:J�f%bo|����PG�q`ʫ�@�wx	��/_��P��h��ذ��:gtќ3�9d�9���ې˖1�V��¹2����y�G)ǕoSu��3�C��1;�-��dWDCͼ����]hł�wa�{��V��㜾��Εf�'f��7GMI(v��S���DU��*� ��wDv�F�K۲��GK��vrJ��R(�	p]��.yǎ9c�B�/x�mT������;�eaRjN��Gs��;ːG�w[��Z�,L�3���x���eqB��jo�B���3y�۫�Щ�/�Q*�[2;�=K�#D�`�j]��Q��ݶ�vWf>)�sNĥ]M�����]���W�Gg�z��צ]Q%t��4⭀N������.�7�D�Ȟ*��q"�w�F�Tɫ0J�u}X&�lt8��}�a�����!b�ѠsNURs�FΙN�!�r���p�>wX�q�G1�����)3t=2V���Iv��O5�xN��p��v1W&�/�m`�^N��lǄ8/2�v�1ȵ�V�����fb�{��,���1Q�˽����Acwi��]s�e�Z�C�p�q^񱋯9�.�o9���_)�T��R�	]���o��dd�b�^U�]��}W�L�E�����8�L�t�G�x��Ƌ�����k��eP	en"�ͥ�spc���`�|���8{&
ӊm	r�Wݮ��n;�q��tR#�r��b��0����ppZ��CĺJ�(w}�7���X�V���0(��1��w r��a";��as�)w3:{7+9�z:�4;z��K�)����X�����M��^0��{�V\U��p��n�-��2�J��y��V�fv1O:�ĩ�ڿ�|5�і9�k����w�&r�#9�ɲG�"F&H�z��s�Y�Ժ���w��rj%�.e��M]�a�tr�����n���ٷ�Gp�(����j�H\�k�jg^]L�Q�-��ʖ,̎W>�����䛺꾎���s�{��o��C+MuoG[݇C��C�=ve����ߋeb�VE	�.���N4�� k^�MW��4��>ɍV��̈́���b�Ik�ɗx����v�{m����
�Rh��*�fl�B�z�l�v�f,�t�p��&�N�-)�w�����u��1��yR����m�6��� �_8%3�����jJ�R�%����6��̳P���5�gJd�\��+��2�Ѕ�[N�`�9�pٺ�4���..��H�:�-�ô��s3w����sA��b�n�H��)31�o�F<�_�?�>PTW�=>�'���{=iؿl6� �u���Ki+�����m��o����o�ޙ��X���)*2���z���r��>�R�`�ŝ���Gn	z��k"�uX�5<�\�U����ÅO��p��u��ת���vK"��}66j��H�t7ug��B�����J����W��wOo^���ջ%kl�2�;��	��_�t^ٗ*��C֓��M�W1������<N���VŴH�{N�1[������tvq��EΨ9.��f0%�Z�o;e�6l�g��-������f�'#ٴT���gh�v���<��s`�r\�Y|k�x����"���']˞B��U�n����3���upN7v7��v�f͢��S�Z^_;��g'�Y˂��u��X�r�n+��m�ߨ="�;��V��"��ou�a	�;�8����iۺ/I��v#��lb����V*��s��U��4Kj�T�#�#S�ߚu)��m��&o�Պ�	qH�����v	كH�J���E�N|��p���Dlv�k�3VSV�]�����B܋�F�k�0��!��O:��(�m;�y�]-�o	x�k&Gq�\�%��q1ύ�B���Tޭ��U��F�*���<�ֽ:�S��������R�+�u�Xy�&k]��%�9�c�H� t�չ����r�õ檐��c
�� r '���C��-����.n��/wQ�xi����o\���A��*�ʢ�!u�(TIHi-�J�����ϟν����3
�(3M�e̪�*�LB`���4�s.��"n�;(��bs��Ⱦ���FF�+=[�r,�����2��~Ϗ���JU�L9E(�EQ�t�9~V�2^I�.j��C�q����������g.UZ���NQD�$Zʄ�F�DPQAT�'�9�ܪ:IW-i�D�u6��)�.ED^��9UȢ�J��Qr�TW�tB����#��TzӔs�PQEZ$V"��.\�!�ub��P��z	�+���C�z������9U:��:��Ϻޕ�E�떫�T��S*4B�"��!'���t�Q�0���h�TԊ���G�"���U�AjDQQ���"�B�P�D]�d!��<��G>dZ��ދ(�#�#�'��B�y��UAG��u�=��������_�����?�a���F����C�w]ϫKݜ��!��|ܾɼ#��<�:'6���+.d��}l��n4�kG���pe��6>�Ov>S�0V/�A����J��g�Ee>��"lM��.��.���dN����ͣ�J{i�߫�~s� ?u��^��fEg<�V\}�2��Ad���U��l<$�������v��'�������)�c��Ց��H�>�;*eoxb�����:WxH)p����+\l{ި<�1K����T�yU�ǔ>�Gd>�<���֑9R�+��|̨j+���8��:oS>({�y�Ǧ?t/��>P3Q�n��+������3��d���j�tn��*H@��z��'}�67<jO8$�eו���.��{r[�}P�K����'��Q�u�Xw�&���y��>l׻Y�mЦ���.��B����K��iw��"��G�D�o�ʵ	f��$���
]���BvsW��{�W�P��^.����u;��R�vR��������3�c�>��t6����,]�M�Y�˼��\��;<vT��*a��f�/�}y���ԆUUsCq����}h�d�;�aށ�ݣ9��̼��R�o�M����ε5y�l�ew7�.�!����Hu��{ݦ�>�-<�����e��Q%Rn1�(�jVe�oDf��1���]�Ǝ��܁Y9����T�_��j���Xh�5i����z�{et�����خ�����`�����#�ޝ��S;��2�?E1��.����� �CW����x��Ƀ�2�6�xC�<\��壵z�����ɯV�I+C�.�����fG�(ު���l�G�����q���8N@��k�Kϻ���O�U���]q឵&���C�M�ڰ�I��c��6>U�
�s>�������@�Az� ]JOn}㱴IC�U��~�1ļ�K��r�D ^���\�{o�>~�� X��5Ps�=�7�ݿ0�̓�X�^_[�쿊�#^��</p2��FYX*��&{"��{��{5}�WX[]A.W`ͯ��d��H���F&��}��Fg}�d��W��uL�\���>����y���q쭾W[�Z~��<�+᷶�-a�s\�u��l�9Z�|IN�u��S)o�
�^f.��V��gܱ�E��HU�����F�t��hh�I�tn�����qh�<�H�m=o`}U��l$�!x��[k�Fr��ɳFo�6ÞE8��ח��WĘz��3Q,A����0�W�P{l,�ݖ�>���C�0i���}�'���@pn%�W}*�UN�g�<'V�Pƨf#�V%�al�M�ݮ����P�m����ܛ�[l�ju�r�z�V]9�M�8Y/�dBMݤ���3j��Z��F�W����1.G���ߖ�%���^�3�K���4i��\�w3�1��fyV���{f>J?Zo�FV�ϙ�i�[ߟ��c�^�AtQvb��+L�{o���<�y��%��.���ԧ�-��^�>�&%%U��XḖ��*�3Z����-ѻ�vr�T����ݥq1�̮�08ڭݲN�s�J ^5CL���Og7����>�@r�)w�J�g{�J�+�����{�D��]��h��*ֽ3��<:xu�|�"��	�>����lC+��+5������ۦ:8=�1��������V�e��3�c�d_E3(��M�=A�x�-F�[u��_:����C�졞�w�L���H��K�-���S8G��co~Ue�SA�Uޚ�Zy��PCS�w��Y���%��LS�e�m¥J�7��׽@[�N3��t:<�}�<�[��������q�e�����i��E�����y�>��D:+�̓������l1y�9u��nw�$���􆠕��{ӽ���[��t{}Ie�c�i�n_��s���[3zk���
�u)+~��*EoR;���U�]NA��	�9c�O��!u�=����྽��It.Hi�Iot�b��=�.�o.�t�'�X����pu+�J�,ʆ,��ZϽ�&�{��} )v������+q<ӟdX�v�Bp����m߹��������jL�+�ژ�-~ga�������}��h�TB��({Q[յZ�]Ndi�KՈ����+B}��������Xۼ��g����C7c{Xy��L՞����=�QM������������=�m�˾�MPEu��6�����g��4�#RSSӼ��x3ӽ�,�d�>,+��X������o7{�訊�l��ް2��9�ە��U����oG,��O������|#�j�dV�Җ�m��l6hC�&
���C��V�/.���0q]D[��(��h1�i��ܹ'��(�"j��86i.r��0uu	Fu�]�&k%=��~��C�`�
�ڸ;�{�T����w���<`�Z3�����o�Q��P���柯�v�ӏ����Ͷ)���X�{�:�6���hC�OA~���*K����ހ�[�~�u.JEF�ps[��a���b
�X�.�7�Zh��j"�Qu�@�:�m�������Ҝ�����X��G�-������ފ�R}�n
7�hZP�=@�M�wg��A�r,�@{�����j߫�\�����}��ۿF��s��r(xF�y%��+r�e��JB��վ҂�eu����Qc�qخ.�m/����/2r����1W���X�o=�k�}�����P��H�-j����j�$�G_W�v{���%-���W���φ��hg��W��K�ˏ�Ԕ�`�]A{���"�:�Ri�0��o�k0�K��q�co"�*'ȑi�.R@��j�㾏k�����g���o,������7)�!׌MN�R���U�^��S�Sy��sY��ZK��t��*��m�~fg�J�d�d�l�u��z\q0wmږNX�z�q'R�R��۵k<�Aaܸͦ�'g�5[7�jzC^p3캊����H��aF�˞��+'��#��b�;\��<�7�.�����.��:�8=��`x��*��;Դ��j���4礼ѝ7cUH�U�^��ꥷ���}^�.���)r�}s�T�Xg�� /R����;��)�|�2�ס���S�j�zp-v�^g�<y����7��/zo��_t�HJ�?[�&g�
���/�Q�ӂry�`�]�y�N9Ք������b�x�8s�c�䆤ձ��r����W2�x�h�;A���x �]��<�w���׫};�?{��~�k�[�T�A>��N�W��� ��M�!~��D�'�
�CUZ��8�^��zuڿ.O�� ��^Xz'����膕A���wI̭��_ީ�ڂ��Ae+G���q����͈�C.f��by�(ceT�ڽa-v�-��"�Kn�=�.�4�����T��x���Xԭ��{X�^�7�s<�4:���>Њ�(�Qq9�B��ͮq[譶�v����S��aVWX��;2egu�sc��!\�o��-�:<C�~��P/K���/fp����)O:���@*[��N9ʑ����O�}sh��)���q�zo���ʠZv���|�!u������y,������.U����dQ��p�;�O�@�Px=+��~�ٴ%Np��:E��q��>�^?y6j>���	V�V<Lͥ�9��PzD���W>Ck����#��MoZՁy��t��&�W�<�u���wIhC���P�ڏ��K۩�Ϧ�\�q�M:��P~�T�n�=�V�|�����W�̺o(W�,��2/���V����&������E'6s���+��n�|���9��h�z��9�W7����������/vԌ��&8�s5m�~B�ܯ*��o�Y[�J�v�w��Hz@��K�R���$yxZ�� ��<c��{ҽ¢U�^15��km2��,�n��9~b�oz�q��Qsλ��Q�ci��F�3N�Z���cҏI@���G=$��=�{�cZ�J��kn�O���[bR4��T2ƷOsb�6sZS��Sa��h����Ppn��,�����{q�t2rv���*�^�/P��Uyu���U��
	+�����^�Qe{n��':�R,?}�j�%l�>���Oco�핅9*{}^��0�٧Etr�q/ݽ� ��>�t`�"������{^~{�=��fg��۳c�]�~�GwJ�1��׵U��{��ޫ�+l�3쾥&�_I^V����S�y֥PKr+����*�U�+�y!��~�.F�Ko'=Uׅ��b.����\>��K����^]ŝ?o_�Ut&w,���mo�*�ĭ8���Y���KG]a%h�U�r~���j�=��������W�B��Ǽ���>z8&��g���O+��<��~�K<����~����O=�ٗ�FP�<<#�����݇�w����zޙ�Z�=~��6�6+n 5����{*(�������xS��M��{ht�Ϙl���emz���a2�|�����wN5B�¡��;�^t������¥)�׽G�g�+��J�Ÿ�	W�k<g'�76��-1g�������ؘ� g�@���e!�b��S�e�Ύ���%�z�d�U-�D��=��������s��d��\���;MoC���o��=!����~�QP����G��7Y�S�3ظ���a�~�ٴ[�z�73~>^���+îߠx{U H���#r.҅��ީ���Z����j���u�һ�4᫋��{[Y[�9�S��O�+w$�W��q�����g�}^�j{$��.�qd����U��������^@d�(#�׷�PI^����,oW�M*Tww�G��;τSE��d��^X�����C׊�݀f�$�N�dس���.p�Sk=^jT���	S�|~y�*�W�f��E�,̈���{�33���C=�Ob	+��R��eV�u���g���l������v�V��[�UϦ�R�� ����z(nM��૥���A>[��0�oN	��y/I��,[�Z�[�j.+��B/v���c�����1-�
�9���G6���,�}�;&��R��%,h�][S���C�y�z^zК�7�3%��Or�c� m����w;��u ��O�����WcH���o+�g���I���'X�YGC�ka�යZ�`]���U��w^�V��|%Ĥ7��	�[������Y^yE���^�����߁����3�Qz#�s땕�{w�{\A%:�4z7��4���B:u,��$�Fދ����G���̰��ntꘟq~�=�_��9X����6����y�G���ʧs�]�ޯW
�Ϙ�T�"�{�B�vR�}�qk���l����y���ˡ�V��B��ꢧ\X�z����puJo~�g�U��.��\j��M�ݠ���)#���K�*v�{Ҧ��xw���D{��k$�W���~�q�o���w��#B��b��)LSӘ��_�����Fy}�I������j�+k���O���-����g���j)�s*U��zX];�F��ݱ��B��ݤ��?o5p�� 7�e���/���v������,}���礑���k(����YZҝz�"�mbq��fQ�B9�����jݽ��#��������*UM�+�aA��sm�s���C&m�sm뛒�|+��T��v�NS���q�V�<�9De]��L.7v�
��<[L��L��	��cǦ�.��.�.+w��׼�X=
����%�m�yX�-���$h��)љ1pw�[��9��f^�L�"N�rc�6R)���Fl�~��(9iu+�J��CR]���ؑfGi6�M����QI�9�1,/;e�8X�b����{��n�j��(�஫	 �Eo���)���Y�ՉEqǒ�U0�Ռ����(��S@�&s�Gr�m�^���Y�#�xT�a�̣V,쬚�6َ��aκ[9�y��IZ�Ipj���[ˤ����p�n��}9��}���՜`�Gj!0���г�[�T����P�[�uʭ�:R$rt$Ю�Lu��5����7W;�����2L*�J|�����qbӬ�x9W%�n��@�m��3��F��u#Ot�^ܙ �8^7w�ַL�v��t`u>a
�gQ��RI:,��^��1�Q����wy����R��j�5�M�,M���+�-�^y��=��hQ~Q�=Kk����ݩ��N<�uU4�Vg./0ɚ�8M����jȫCV�-޷!v�j4n�<J��.]ی:i��*B�W![37�+[�իJzNmgQq�a��B�n%v�ŹH����/,���㗗N�6�k4ڎ��᱂a�ȯD�h2� ��`��I���0S���=)�wp;٭�((�+����u�[�4>7%-8+��q�ր�̌���ܶ=4��������ɰ&��,���ge�o�@��Mۥ86��}�iL3E��nu�i�A/��dpL��CBSW��w�]EB��yYh<m���DT���J�D(�֬��b��"Tn_U"Xǜ�7�6Q{C��O�z2��6�x̽�^�V�]��G<��(��{�u�����D�\w���q{�%H�)uԴ�Y;��vۈ���Ħ���WWc���ow�`ط����w��C����TnCH�0���;���f�x]}\1ğ�U1��B��8:��5��nt���
�Oa�Fb  u�_�:r��}��2�OA�h;�(>P�!��X���_WEBC�6�:����EWԆ�$/��/�io�>�n�痖@\L��ST��{C.�=���<���QP����;5����H<�8�ܘ�᪸d��R�-��saz�:�`X�x���n�q�}>3%��I����x�o7����r�m�q��k�rl��	N4�LZw��xO�Q{��%�F�m"ݩ��X�ۃ�r>�jawaq�+�]I�f�yˈ��R����Z�� \����zt���W��]>�d��o=&�$
�+2�2/L��l��k��*�^����s�7��w����|���9_���ZQ��,��
�1~�E:�E\�����~����'�\����E��	S�2�\�'�(�:t��✊�������|9Qr�*�QDD��*�AAU���*4 �����D���r�^��N��� �DW��ZE'@�B���Dp�Μ��t".T����D���\+Ԣ����wP�$�̢��e�!�.AL��YUQ��
����G.�G[�5ȼ�PPE.S��y�U2�����E� ��m:�OF�wSVPP�
�+��as6S)����ʫ�vQ�Q�"U�©*B�}�̄�wu�S8UUʩ��{�G�QEEU�l��(�<�Qʹ@$��	��</�r��Ҙ�Q8P�#r� ���w�V]n�ųY
�v+i��@�:���5+����
�.�֩�\��\2n��������2�m�+��mϑO�X��~���ܥ�o��	�u# ��k��5�1¥�{���Uz��o˭#��J/��L�\�N/.�����V�No(1�x��^��d>X�N#�A{~��&�穟�
P�Ś����Y2װJ��+���Dki�v1נ(�tGlI��v2�~��%��}�sŜN��NH�#_O�__�����|��q���qB(��WpP���8UՇ.3�5��K����7�Q�>%�G��	���U �=퐃����d��DӬ��VsP�ٖ4��5m��ϩ�q�3�>�r5g	�
\m�3H�{������R��A^�S��z^@�<��C:R::f�l�)�ec�6���}=�迏�$�?z��#��^����V^xo�l��Мz�!o�UT�[�ǾS6�~�v��E��|���>R;Fy�Q�N�p9������B\m�����h��k��E�I߹N3�ąG`�+���ᑥzK��5%�g��� ���>��g��8�ښ��_��s��E�+�:;D���M^y�+!YӇ"S��V��[����]���8��A��|�QQ�Wp`������oK������gseJ�����ȥ�30�m�)��%��i�2���eaT)>&oiyζ	p���{e�׶z�ȸ쵍IX������ٝ�IY���WJ�yr�+�}hz=%��p_�����������0D^��>���ʑP��,�?~��;4�v�&��/��ߠ�N�O���')Q2
ആ8-�GR�*���Ы}�/�͸����Чa����wԦ�,#ق'��c����v��~��^=��+��$�s7�v��+��m�������sj,xx���G��$txЭ���r�����=�&�x�ۡ��u��yy[���c17Q8����9K+�_��F}�uf���}��"O�����T|��:����_�����ܡ8�/^d����*���R^Y�s!�z3�kM�ܥ���)'�������_�q�>�9PyU�3{������J��ݪ�q���'�BS�:���H���\l��xτ��X��l{|�zc.��צg�ak��,%(3��-��r*���(��\�c$DÑ�=��7LuB���eR3ϣ�A���5�^��ꖍ�zX����ZU�p2���r+�rK�)�F�՞Ñ79�3�г�W#L�5����ě�E^��Y�Y}��Y�ٕ�:4c�[����I6��]����KJ�v�s7��G_�b;kW����ky��=�Π;k."�P�Y}x�>c2�ۦ8���|����18/Dy��ͮ:��wKq�~ `���J޿~$�_��J���2���Q��Vu(Qc�\6qL�+>m�ǔ�23��sɨ�:�~������T��2��~ه�px`k� ��!�uD!r�u�p�2|����S��Fh�����W:�v0��O�,��#`�3����A�'`ǃ=�#kdT;^w1�1o���F-��}��ۖ���e�Q��>[WƮg����D�|jJq�ɶR�=�j�E�@9�ǹ�N{�!r�J�����D�U-���W}���&�=�b��~=a�OJ�R�z���B��{�����#�ij�`c©i����>��T�`hg,�,q��#�s*��l�36���y�c��pdC�﫨tu���c���v}��̆�#���"�=	�z�
�<et��[�O5"�?D�ң�#̯��{������t���V��+�]�d�SL���'5�z��U �Q3�H3�\'p�}먆�����������,��pD�Iջ�N��0�TB��Ҫ����V:FAF��,"&�O��3�V˘~�y�G�ѳ�S��ͱK�xi�t�36�͘��?��r.T6�:%	{ؐ9�-^&CE��{=�h�'�1��:(�f��j���&�\��l�'s;�SUܮ�����Xw�P����5l6�IX6P`���0��Tnk׵�՝��v�·��$�C�$[y�^Fx�[�;��܆"���P��:7�� Dx2&h�=�xs�9��b��ږQ�Y�~�Ts����V���-�Qk��6ߨ14�诲vˋ��rK��pS�[ȅ�Rh�[���Y��0�|���]\�[U�Q���:N-�!����7֐oz�T<���g��}�؃_gn�*sY�:)����~3��'#C]l7�wP�9�q��Aüj��p�4��q��ɼ�jݯ�Ko�f��BcV���c>��"�"�>Cc��@B�t��s�7�Dm�>��#�׎>﫠8�iл&b�[���Z����_��,|;�!KK=2b�ՏoDxz9X���]<+Ц���7	�N��,�T�Z� �'#�(��>ܴ��p��fϟ�s���ޥ&��.���08�°��c�OYQ`�Di�A�Yy��z��c���棷�	q
ؕ��nP��m�bw�qg��NT+��R~Q�� �-{��j��~#H�����5������<'a_¶����d<��f}�ړc�Y�c������_���kw{ؗ`��*ম��A�� �^K����M�����˯רνʔvA
5t��QDL��vkn��/Ot�A[�A��U��ͧ��Q���;0h[p\�`<�ǻa:�:x�̔�eG"
ي�/��U���'�A(Rb���&ŗ����\�#�'���9A��G�����^�ښ�{]j2Kw��u=(W�w�k&sG�Y�,�Y�{�_ת�/\�v�� J������hI�.+�1�o���59Tb�DZ�滗����s�:zϰ%_W�ܦz5vTB�8!O0J������˺�*�[�qmx��o8-�36�J}��B�T��?R��;֔����Q�X&�h����h�'މ�Ie�BU�n�x�76�w>��*��ߠ:7�[�bC�>��:0�[3r~�Kf:��P�=~w���ĳ�>���L<.*nr8:�V��ѝn:/{]�U�S��Xb�:D�;]��	����`���ޯf��KL��a}@h��{8J���U^��q�X��3��s��*��f��/9�
���`��\�!p��u�J�D���s¸:�@mm����c�tu�Ek��7}���G�N�P�r�W�X]>�7��<�z��|�L�@�tF MyEL�[z;��ϲ���j,)���E�5	�V�2g�}�g	�
\o��v.4�oec�n&�9��]A؅���	�{�}��9�S�h!��m�4�{|���S*i��m-�o�.��\��.��~;��E�F��>+Mv�D����lu�Ve�	u�2�{u�mp�>�����hP3�;�@��\K�����	:r;.y�Tt��W�V�����X�F:2�m�ފP��(��4�g�)�ec�
�V�#>��tX>���׼�H��#�{�������LE�J������~Ub�H]N�(����Bݽ�������_Nv`�+DZn-E�����X�,��d1������6p=v�E���Ţ�d�GU������<�K�[�xF��Ycy
�U��]@�}~��=�7jj���q��[��w�~��O���榵��e��CФ�)�_J�h������=\G?]T+��'�0�l�Z��;�ds��35Rg�����[��;�����&#k�T(�������Ǌ��6Þ����x��N@P�W0˿���Nv	u}{�R��{���c��yUS�+{3�"dn�v�S�,xMÊ�OG��ۘGK�lL;��m����b��nmE����c{��H_�g�xC�3�\Њ����Y�Ca��k���^'X�[u�]���,w#�\���ϩ�+B�_R�����k���m�u>���g�\E-\Di*���́�Ӛdk�$"�/2�m	�P�l��3����/��f�,W�M�-:�p��s�^�WV��M�7����Ʋ�y[sp.��kl��Z�뼼��ڒ�Ω4��[�C�k~SV�ݑS���=�"��.���*s0��U�����A��>��0��Ѣ-%Sk圥����
I������Y��?]瀿���v��M�k{ϫL�;��\��b_�?R&�`���Y�\|8�W�y����;�?~�
G���6�x�0.��K>���\Xg��e�o�@}�V^}�~�v׫��M*���xP7�՚��`C�MiQ����b�������=<�2��b�<��(rr��o7S�6h�.�f^I�:}E	��z]Dd�l������G��f�X۱�)=����ہU~��+��uo�uh_�f���gL?�� ��&��~�c:b��Tb��nG�ӭ���3ֳ��O��E��l�.V��t�3���b}��렂6�EC��I�)
�/��/9�=���X�d4_�I�x�_��(7��)��\�8h|���#���Ś��.��ϗ���Q���vځw�*|f,b�l�|�(V9�	5\F%|A��
w�I�����5���j:���M���/>W�1B��/y;P1���WN���C��W��V⎫�*���H�G�;��kKvy�h�e݅���i9��R=���`�EX�"Xl�E�8�e�#�3�2�^�f�a�iP�O<��l�n��*uTa�˜9N�Zj�Kk-���31�w͚�a�SV�quo*���f���7��u��D�S+����b���I�^��Wё�č��tm�ڬc�/�p{??ܤr0S����8D{C8�v��sG{�V���%��D���X�QBA�*��D=�R���M�X=W❕��8���>4i�����a�q��Q�|¡�x�+�=!@*�0��]���/vb4��� �݋^W��ޘ�r�L����S3�h��}# �_i�g���<�j|���?��8~'=�]�q��&g$S��ƺ���oH\
����T��7�5�ao����W�'�����m�o���8�k����i���/M�l�B�b�{a����;E�I����2��l�Ҳ��;]���`��OŅ��y�W��W8߮mC����>�~�b���xݭ �C[��7�G���o��H?��Tܗc����%Ǣ�*T<c7�l7�n�X<�8�R:��ٙ�!�_�}��������ymwH[Ho���S�L�@��T�����"��tnxwTD���[���f�S����L35��n��B�O��7�|e���?K`�����<��W2�{�<'j����x2�v��"\˽x�'�e$�zV�J�9�GsR�Oۂ���U��;��<^D$VCUr��U=��9*>��ͮ����ϪH�XpJ�e�� ����Ž�|ȷ��P튳PqJ��N=�����+ �(ͮ���nV���Z?����m�:��k�w�����/Ц���#��6���5�T��߿hZX�̜����f2�m^��N�-�tX�B6��
V�ɬ�\�t�~f�X{�1֧�����˽�t6���I~�8϶�P��႙8hK��WPp�nX�-�$]�N�M��q��	ʄ�T��U\���{*:")D?bJ���� ��}
6,K��[V��U�P���7V1=�%s�Uf*��� �;�쭝��=e�H�o�8A�� �O@T t� C��SQ��u��e���v�5�gyi��j�79�,y�G,��ڥ�1�N@*���:A��F�Ɨ��4u|�M��W�at�����s��<�������U�k��6 ���V�hԼ��h�-y��θkA��:o�E^��Ζ�~�W#J����;>5�`��M.�W�?uV��WVN�B�A�"����;G4��J�/mz����o�Ć9��:0�O;K�ox��x7b3\�/%�Y���<%EB*<&�!��sM���c��Q��p ��c�[��y�MS���ي�ŷ��w�[�'o?g\�W�^X�ʿ?F��rgh�Σ���һ�^罂?'Q�c�Ʊ��M�ܾ���D��r+���X���xo���e�ޗ,|����qfɁ�1�2�NC#�Ɯ��ҸY�����[������,����}"4gd�7�W���oOᦰ�V�S0N4k����̵����|�8l$��u.�9��"�ez(��+)��`g�(u?{��x���^
���%}��H`-�z���`7�s��P�
�ǫ׾�hO���|�ln|�1,j��pS����60�G#���#�`?qg�EOmKV>>�?���R�ꦙ�V�*�,�a�r���nj����~���Y�g	�8Y����\d5�ڶ�H�1�3H�z`���3�#c�i�ϔ�2�>�p��n23��WC�.h:������;߱�����cY6W�d�	�N��0)d�ԩ��S��S��f��V�ɉ�}�ѻ�	v$*�����,���
P@x~���_~�Z�Woݷ)���:��R��f@<ނ|�;���^9�8Ƞ����hz�U���.�z�N�Gόxrc��WՒ�h�[��e�m��B9y��-�B�GI�;ϹP�bVz��"���Ø��B�H�<�Lc�JRf1<���%||i�Q�P��'��fwSg�����[��uQ���Կ�~�#B�#� ��g�����x����h�T�6��y�<zn��Ǧ��t-��qR�|Q�=xdGf|�C�=ϗn_�x�"��M;gΗ�`��e��B�����'���\��#�*�YB�e��)s-)צ������O���2=հQ���o$���eTQ�㛱���q��A��]M̚�*�2��d���y78uu?���mm_#�J��r�	��SU}5����+��뎑����+x�*e�����5c��$�L�̋��M�/bDTQX؍��_����U0��X�VT�[�xZ6���WՎ
ǫ[��ĒC�o@Y�Z��e��&����'Y�2�S�s���
����F�)��;f�(��T���S�Jl���q����Qnu�l��c3'�[�ŭr)��+3b���lqu��������!�sH3�Vt7%c���v��SaC3d�X��.Z"ˡ)u���g�%�l��\���98#��g;0Y��Ì�7���b�Wro�>��m��4���F���H�
��wj!�����=�����q�ʈ���ݛ�����$���v�iY��5r�^P�SV%�����C/��j�]յJ�:�LYj�E)T�Ҋx/���]�;b�H�٫ru�Ea8����� ����梸-�Q�f�r6���\�&Mn�ݹu�X=])�e�삾tPD�<���4�N�r�J��i�Ր�]l�W�G[���-�/��$m-l�z ���&%!uL A}Ö���vݣ ��R�yE9���keJ!�&�5�׹�m��ihحƸB�ѫ���`j�S��\5�ɿ��Q��jb8B�c���Y!�O���5/UJ��A��EQu�Wݭ���J�0�<�:����݋	<V�z�)�i��v�kWo=�[n��V��� \�e.����P|��X�BX���cU:Rm�������1��;s�J0�Q�2�<�n�t�tÓb28;�7^�T&I$s�������%����Th͝%E�����Mi_K�
4W!1�o�s:�]��b�fot֘�jh�y9��{���m��WN�U�C�X;cT��yfĂ�#j���jdQݵ��y�#u���t	�%�,v*�*�C�f�����Eww-[:�e� ������9B�pSn}F�S��9.�L�v�u�o�A8�U��v��
�������^8�������-����g3���|p&�(���w��$	d+�!�9q�S<+.��N³/u��m�<[{|�
�rֺ���=�O���U��m�$�zbH�b]	}�Enh��M��9,V��{r�WnnI�5�ta�#b���^'�;��և�LEX1�*�ֆB�w2��x��ٝ/d��z�}[;��=�ܟ
7;�Ty���le�.�ڨ�鍔��o���,�ٶ�]q^1�=7{�]{�<�:U�Zm�Ai�&�t|������'�G�\��]���,��p�,Hd(&eQQvD�7�3�������*9,f�r ��I.���ɡ®W*� ��������$>gaEDQr��A��CD$8Eg *젹E<ޤ)���"�r���BL)�*.s�I�aQk��%q��$U�'�wf�fgI�����[+��QAa���*�(-������Ҡ��ʸ����(QT
9D3��SrbAjߝܢ쪈/8�M�$�$��	e���SC�E�C�Qw�S��;*����T(*�.5�t���98d	3S��NU\�>�9�^L����I�����ʨ)���$G��9\�
�g�� J���H�Ĕ� 1/`�;�/WR�uu7yaǼ�������b�s�W-/�Ni�(��/�/i�kQ[���[� Z"Z$f�;� �Ж�oc�nY�W����~�'���ߟ�����A�L�r��`��>P��h����Lx�����v�j�����S��q.��r��E�{��X�;t-�0�N�xf�C3�8��:t�,i�>;Yޠ�����z��U�y�lP[mͨ[W�D�X�yҞTe��g*�Ʈ?V)���E�~5�Կ���P�<<����u��CV��}Rᝡۯ�>��~&�ݏ�2 �q��Xe��L�D����7R�}S��+v~�|�>�����UF��O���1�c�E�4�b����l#Xe^вdx)��V����?
�r�ېf]Q�w���3�/4���SZ��
-?�HBj}���;Y�\|;䚠�y�[W����?o�T�����X�Ox���{`s�5q�Xgc>e�o��m��
=�#(ܕ��Ƙȭ�By��-n!�D1�HU��5�Y����b�հ��Z:zX��9M��=V-�P�`�W\�̒k̰���n��뜓���4G��Qte��1�@Χ
8��S4��y����.�Ѝ���[��_[%R�-�'��(��~��0�b�5��	���P��/����ϝRU_���+�Oy�N���D����?{,MbS��!��:me-��C�����h�C�g5V7�r6��U.4�)��}�aJ�N\�3?!�ro�D39��S-��������Nw��u"]bS�}X`�cSac{�Ǉm�0��`�5o7�BNﻶF�D�b�a'I���og�F�FGCyƅ��*��	��_h���'�_IA��:� ��53�Ч�۷��=����琘Lw+��WI�Jn-�dq���k�+����P ���r�Gb��Ǎ����]�*��ͣ��_�Z[Nwة񘱋)�X��с��&"{�|c�kZ�N;cUv�t8#jd(�6:���Y���ZFrt� 1�t(��`W�僱�¦��qu�u�k;ޕ����*�Ð�+��������c ]?��>�����,yl�N�P>��=xg<��?��S��q�J��@�~�cOF	̫�n�ߺ��M�V$��rCʁ>�>�S������b/���P��gQ�PT(����fw`��l���<�d�ԣY�Ǯ�ҕ��G=�n���1a*����)h���\}��%�Dމ�>9�<�P�����	�^�Q�l��6��'���zqW�A l7!�k�c��r�#���+�7����Ti��^��=�$[��8�7�Rg��s�9;e������,3m�E�3��_�Y;e���Mc���3�jmA�1M6t�巟y�PKe�yBE��$8$o�2���uj^e�ƭ;�fY���i�U�Z�|��'(��8�E��O-G�L.R4�l��7Gx)j��Tw+��$���_X���˙�"�F���n`�$�A�8���u�qZpp��dQ�BA��)M��}��]�"g����D����Z/�+��Y[u�\�=8���[���2�ɏ=�E�yV�;�uD�^��jJ϶n�%ǣ�J��H�1c]l7�n�Y�+��j���:�S�σ��F��x�����}�HYti}��U���p"=���{��+�kܺǫsF+9�2���3�3��*p��>�xޝ�r<L��%�}b�{�_�v�J��+:����8��bw����3P�	gVB��ہ��,�T�cA�~|=L�Cљrn9�m�����5���cnP�alP�azܚ�:m��KE��n��$�.��0#���4DMb9��F��CFC�������Ӓ+�;�61N3щʄc�l�\�s��ĕs���3p���A��w����O	��\��
�����ړ��޸:nE��ox�Y�=Ӵ���ٿ��gA� �bz��t����n�5�R�����bry��;Y�8��Gk��@c�RӍ�G,�R��~ʈ�"n�* � �R8$Ɨ�}�oDezv��^�^{��C�Ͱt.��Nĉe�.��o*�ev�y.�U{=X�4��Ub�vuN�e}9p�ـd���ne�mN�\ř�d�<���!��QPc{,^�n]�}%RG� ���R�4.-��p#��r�֨�99w���>?ʯ�U��@���D���to�Ӕѷ(��y�C)ӄ�9�>��}^7�*��]���8 ¯���� 㻡C4�Q|����R�N����I�<�s���B#k����B��alH�XJo�Z'!GX&x�:�eut�n([�������-p$`<ȯ��c86��[J�%�@to��"&���l��]A��]0g8ŷ�ν~c�7'�zj�x�𛜆�uϴ����E��wV��{��cW��ɺ�-�Kք�_>ܞh(�_��)i��aqg�ˍ�M���z���7�U�{;Ϊ��(�\���O�wzcs��9��p��r��5��۟��~c����BSށ,K��/�\�=�|��ڕ8+�cz�j��=������lWF�!ž�E�O��-t��"�&���8Ñ�F�ˢ\w����w�����[T�����w�İ��SP��up�
j�a=�#�r8$5�w���2&s�]�<��0)����F#�@~�w��,u/&Yl�
f�Y��
�j�dE4Hר��DU
cyqT��?~X��ɳ�Bv��8��`=�L�@.�m�)�e9-�ʇ���m�z��s��S���dt�vfǝ¨ۤ���]��;���(��lj���5~�z�O�X+n�X���qmEW3�`��,�Ժu�ӯE��S\͈7�^ӫ���
4E�=���
�0S����������w$H�O#�]vT����V?���ʿ�}>����.�v�lA���߹�@�O�����l1?H(K��[\P�k�Ƿ���p�׋r�#�%��l��%�Nqo��	|�}5|���>��e�}E�E|8�{�u�}X�k���U��P��;�����Caɴ��g��u���&'~c�*q��u�����<���q0�Ų��^2})_�0r��F5KS���#+��H���;n���?/��pŹ}���A�H1�K=�k$���v1×�>t?!�����l�&϶n����s����������3�����3��Pℝ�#�a���V'��+l���\��r�!s�y�0Zx��5���wey�B,3�`H?�L�����~1��/XڃO�X�k�/+q{�{�W0���WꈜpsϺ���Y���PJzH��q��a�m
&X"btd�T��e�u��a[�e��O��s(I���vi�����q�)����X*��;�Dٕ�,��R*��@��l�Jʾ�l�e��ދ����������k#V�`�^�!E�����l��C����d��'����M�QR�sM�F+��Y�I+�&�P�f׫��w<v���qo�g�A{��b��N�V�E�x�Ϥ�:Ȱ��uyn���û�k���k���g
�ǆ���"���㚡��ca�
��sG,�7��.��l?�郏�^�_K"������@��|8_�����`y���9Ƅ��w��ټ���v0-���EC��_�ڞ��5'�X����a�4�����}�D?�:FP&�q�fm��l8������=89M����_�c��������"�{t�hn\P2��W������(?�|�	������ȏ/��ƀ��?|��2k�oMz���_�ʘ�'p9��vд�;L����
�ND����O��`���=�0�C^u���ټ���s0���(!�lq�l��*����0����%{698�6<ό���Sg�X��)
���+���^	VCE�##��25zkMw�g���yk�uJ�������LP������W��Ӂ\1S�1x��5�'J=�Y�b3/7�]�*lEz���8f�Ő\�"�ڙ
9���o����1aT����@��>��X-���"����!ύO��8���O�ՠ� A�t������}Bt~�c�������G�Ƅ�3Whn��:��a��DX	`��G*����~cg����V��=����ٹ�*���+܂p��{)Ÿ&�ٝc;ξ��t��8f�{�8���f���8��W�9����v94�9d�'��8�z�Z-�b3l��V��ں��7�	M�#t��=Ͱ�λ��h�+�S���Q�\����ftg�{}ݞ�� �������1	k�\߳������~�E���E��1� �"I�
A��K� ��<^>��3�h{^�q���#������TOb���hv}C�����t�1g2��{,�=�'�x������ѫv��	��HH��E5�1K�r�0�+��\ϟ�C1]w�؇����%؝d��#��}�#>핧�[���,37�[J��z6sӹh�Q�E;�G����(O����7'�j�6A�eZ/��tb�ۨ�Z�A�ϖ�ۅ�^Ww���2��U|/8��c�֐��Y�:k��E?���#�#������׵U��]Gջ�0����U�w�Q����S�X�W^��7�b����8�������A��>�Q8�W��jY��B�T��R�8J��:p_�ӱvL�_�n'�X�}���W���ǫ��w�8�q�!7�x�H�w���e�Fj/��p�T�q��"2�Y̮�J���w_�p�J�s�2�$o�b��B��[�Y�l��Z/`�sz�;�|�C]IpC�QA7�u��f\�6��l]�4;�w;�)��b�7�°þ��l��� O�^f�5ی)�-�ra�.��~:2��j�K�1��3���b�1��zΥ������-��4�E�%vq�7�z&�s�A��8��=�Q�͎2��������]}_� |>و}4�l[���n'GLG��	q�+�8V�,Z��ܑv1;�7�q����f�
T�C��d�z�o�?�|���A1�al���B�韟��ݗ��
u�<�P��)�}���y�j1u|�j�#rG=����.�[��_��*,�ݲ�����?@���m�������l�ϳ'#�l�Ըn��=��V@���x7)��ڥ�TGZ��UBæbyV��	M�F�N?8Ӑ��!#}���Yzϰ%_W��U]�b�8  �DU�u��{sj��z��H�H�5��v�#�7hDnt�{�)��7�$w�����NB�ݹIB2�q�s��02h��\	�}�TӬG>۟io�X��@tw��7�lHdeB�n���	RM�ov��J1q����Lܗ�0q	QPǊ��l��s�8�S�������7�N�7���8sg{��嬁o�?X�iR���o�a�����=×7������.r�䝿y�:]o{��s�k�#���<s�o�[���s�c�w!d�Ԣ ?�z���Β�,g���_�{�YW&�|{㧂�E� N��t��t�":����gyc�dA�ʍ�̎��ś�{fp��E{L�+�!�Y�3$_jtD�e|��Ja;��ĭ;P�	+���u�/�n潔ݺ�C"Wk}4�s��ppDFPG�_m��m44���"6��;�m��As�ps�!���U��S����9fQ���v�Vz��ed�������y�b_�&�/_�T9c����w�}2�"�)�-m��ϩ�q�&{��mx�~��OS�����M<�%��	�C����f#�F\މnu$o[>S4���.u��{2/}#3���լz�^FC�wձgӒ]���d�	n�6�����0Tɑc��_��o�WS3+^n�'���<���@��O������`����:�k"����5��	�c=�ɼ�0����6�4����>��+�����P���ui�2:.�_�5�w�Y��>��<_�*�`��3<��61��rl'=��s�r;�&8��!lI�i�ɹ�4��oo"�ŗ����J��)U��z�=�a�[���uQ��p����fR�̡���&<�C��H�}�RcO3
�<v�j����;��W׸)M�B��:.{�fo{G{���~c�$ïL��K�$�yۘgl{���*l����{oԓ�(���$|u��~V�vQ�zG���[~'��F��&׮{���U�X-�!I��n�-M�Y�5�a�I�wd�)t�Y�-���S�;eTZJq����Wݳ��i}x��b�Ї;sar���g7L����,w����Iɷ}��J�2��D!u�����jo���1��kc�q�����H�0t����5/�f���wX�8S��''nK��Q:��=��lՈņ�!�5=$R�8��2�D��ѓ�Bn������z�yVFt{=���38�-r��=��*��$b�u�b-�S0�c=fVȢw�H�w��#��p�E�F��=Y����k#B�lk��8���!j��n���O2ub��2��U-��C�I``�
���fvwN@uT=a�W7�k��v3��8Șz�_ނ.�!�E��1���Bn=g$��pR2�M"�r��1ޝ�ꖍ�zX��9M��!�ׇ��^g[��p����0:�@��ݷ0�Tײ���C��M������C:�(ӽuP��F�<�ޝ>ԡ"��ix���>�i��=^�]c�b]�z>�O��`��jP�ԓ��1=瞀��/8u4��#��	R���#!�y�ͷ�Ǘ;�Բ�"h��|����%�����/x_��=i��!���	y����t٬J�/�##��27V��z��7=�1n��k/2�4�o���v.z�P�r���aιK�Y�aՎ�=��F`�ݣ�]o��.�=<]�EM��ʝ�鼺�g,�J��%�.F\��Κog;s.��Hc7U6�'+zƸ�_X����V3
�A�� l�C�8�k(:E;�Jvrn�/nEm��	�sU7�j��v�֌��}AdUu�Jd
����-n��*�Z�*^Mɲ�]��W�ߎ�URUsh;��/Y�ec��e,¬7@n�2���U���;��m��u�/�}i[=��]�y��S^F�V�N.�w������>�6�c����6�^3tfGm«&4؝�Y�)S3i��}�Jfz���=�])�������v�BދUD��[���F62+i�ǋ���fT֭��Yd.�a�լӚ�'C��-�	͡�k'hVP0�5�]�u��e�`H�S��M'�wG��w���P�0�r�,��c0ˎT��� +����zw��q��*�]6z�D=�v��2��Y�ʰ_-��e���84��w��vB__Zֈs��tqe�=��*l������{5���n��gXu�\�g��m����~�J��ܣ�\�eN�Ws�I��u�g��+Q�M��nuY�y����!Iv�c]�0�WY˵�&5j҃gB��I�G��i��R�F�e�+#T��N�c{�he�K��`�m��N�>�X�ov���ne�Vqվ�ڴ�ܙۺ�z�#��Pk�k��$�K!H��Q�ۧI�}��v$�y�$;;d��=�e5�y�zֵ����z�%ّ�E8u
6kL���Ьj2�q�����uW����ݡv�u��0�/��٥���)Ԩ�r�����}�Yi:Tif񻾾n�[2J����t9�a̸��O/�vs�V.j�i�xHP�.��`��G)��
g9pK���rL�+�&x��RJ�H��O���Wu�Kl
��5���f�tr�̓���.M��nơH�H\��N�t�䝔.������x��+�
N����(-\�ѷݦ���S��Y3�-���e*�P�W�";�%���_c 8��7^k��z3�d��WL��N�!��Å�U[���)�:�B���2�T��(���T�-��xnS�O�vR/]�s(���6��Sp�hh)���ܹ�Z��1y��mQϢ����Ti:�n�Ҩ8W��+ՙ��%M�~�ޔm'y��[6�f�)�yN�擭zu�/��sw`9[�kq��L�g?�a.c��d���eK{,�i���#::����ef�jԚc�s���''���CCB]�����!r��x�~�[O6�(���Ψ����s�7�� �d2�N�(%Ip��(T._=J�v�ǝ�	]ό�݈Vҋ`i��/4%��f"v����=����$�$�G��f���4뼎S���J]���S K[r��mI�ݏ�>���q�$����^o$��Gi,���t3�'N�S�iN�����?G��ƿ#�<&�껳w��8��I~8������·�N�[�"����ۣ��Ǐ����!�޲�5S�<;���\**��Y����<���2�EY:p���wwq�y�2(��jQ�޷"*���]]�ċ���8���>�*:Atqr�]ɕ��
��p�w;����6h�'��6�#�d�L�a����F���z$8�@���8D{�;��3/P�rs��~z<���2�I��OP����zRT�Z8y�	�()!99�*��i���΄=%G�ayS������Ú����5z�r�=�'*.*����x��*�<�
�Q植�W/*/DΒ~�UOS�<�VxC�J�S.�Y���e�Iݙ\�!!!'8!U:)��*(�����P�TY�6����t�ฯ�k<�;u(.Wo�����,��h��d��^�"��V�/ˌފ���Ny�Zf�뮹�%s��H�U!pcp��05�x~4$����6��~�k�p.�S�1��\�(V9��ES4ERW�y�.��>rp�c���d8�o�o�ς�XŅR�3 ��@�}]
����4���5��s��?@~*�qzp�?i �;P�E}!˅b����P��/�؇<;����U3�C��Eq�`S����
�p�B�'��J��wJ���!��Ǆ٪�w�qx���vo�@�du����) �D_ZwP��Σ�
R$���t�j�B��؛woҁ�{gۨ�����P/��1a*���꘯����̮��~`��[q/b��x�ˀP���ؓH���C|u�	=8��ޠ�6܆"�k�ax���f1��D�1U��Zȼu�c�'DЈ�B}�*o�z�5G4�ol�6�[����̀ߨ19SqD���H-�^B���.:��ڜ������6FO���]\�Z�T�9.t�v�E݊���;��b����Z�J֐o����Tܕl�K8f�`���k~�~���#�PO�X���� �S���پ�w4�����i1niVr��mc�j���/�!��H�!�j��;��:յh�9�%�7���hxJ��֟�^�
Q]]8A��k������+q��ڱ��s�̖egW��dz��Y��O�m�����9�+���BTD�7��7��Xb��(��b�79Pp�cV-��ޱ���M��xf(9%�9�|�=��D=3�j;3�Nѣ�"3�W�C<���X� Fi��Ӏ��c2}^����1����tD�+^�kߛ��|$1�Xm�R8#c������z����3P�~���ڧ�Nq�3��~71n�&�'19���:b=S*�c�P��$K��rhgM��s�h�8�¨�q��1TK/7VD��cg��"i�7�A�G������%�B���$]�w�j�qW��5m�؋뷩FT����t�vR��l� ��h@��~�\lT�ښEʜ��StT�7=��n�c�ړ��H[��l?H�6���"X���������[x`ּk��v[�~��+m�C)�@�]ON�#�rڥ�TG#p
�ʄ��;��C��V��Zj�6!�&0���LB�U��Jv�d9�>�%^��Uк�!hS�%W���ꉠ�q³��0OA|(<�SVr���˫vv_O�{!Oԁ�Q#�a)���<���n�=ي�ԋ�ֿ��<��T��.1���f�l9������P��X�)��l�=�3�����݅�����γ�[޶����`[yc<���gH����'bvM	
zk���A�M�8Zg���gr�̊Dv�=���S�7����Jt��s��`�<(DF��k��,��У�݂L:���bA�7[����J�/mz������z� ������)nv��'<��j�)~��{q���a���R���Ny��[�s�u�7;�{���v8�a�l�PcZ�$����ư�Ph�,p�����d�^˦Gp�7[\�zg��^,%U��;���m1�:�k���f�o��Y3�FE��S�V��g�r�g��̯��b��U2\hm��K�����cSL�����O�la�2�4�!�6z���� k�lqƎp�U`��B.�%�E�SP���\<���o��r��
D�C��`�x����Z��$����n|���WdPC:R<L��jf�[�}�c>�0���fp��[��#>��t_�ӒW�B����Ń���C�m�S$]�{<R1��#|}9��kW�o����}��3|[��=���.�#g�����	a��.QfU���z?ގ�J-��˒�	�,��I��r��)�y�3A"��>�!��]��M!@Gύ��(���]��tr�F�R�w0<�:ؾ��ؿe�;R�}_��i�.pm�)P�9��i�KO3`�lѾ\%�?^"D�����A�*�3=+gk�a�Z����4M�9�!�y���v�pB�޵PQ�C����7��3%9G�d�ɶ�Dҋu���_6ӁQ��� �WKL�]��Z�~z(��SP��_��gk���*h�㡰����q�ω�
fɄz��NG��.���c<�8�LB+�:�_���JW����6z0y�Xk>�_O��=U����������7]Z�b9���~�y*cKFl�;���<Ӂ���;�]_n}�ܑ��g1�>/՛�M��ϱu��m��+�������D_,*=C7�N��H�L6�DUQ#3!����6�z?!A�'X��C�b��H�8��ŏ*�ⶤz]~�ۈ�Z^���ٽǺ�}�G��w�xu�ņ�!�5=$W�D�=fW��,1 h��Ty��R3��=����c��������Dm�RF-��1ҩ����l5�U�'�!S��}�=��0-�c�����g~~����5�o��"���-?R��A��r�הu���Mֿ$c�>/��#���}�)��vwN@~��Κ��],3��e�lc�P�q~�}�R��c���͞�V��|�ń�t��H�(9X&�q�fm#�[.K�K��:s|l@&��D]���E��vf²缾e
�˭[����X��\϶>��^Ê�٪��a��	P]f���	.<�{���2۳W�n����S�)dH�����G�Q5;YZ�Գj����N��T����Ӕ4�k�kG=����9�Ygf��N^c��W»�aT�nMw�;�}��5��t����ZuJC��G��/��*>��TF]ٍ�1�[����V)A��t-��5?�eƣ�f�M�Чi��=XD�v_����_|6��^�=�C�}�����cB+9Q��ݸ~FC��q�l�|�,��#d����b7����+�=q|���xxP{(qǷAV�0�:�C:����PGG��ճ\k6��=5���f!�aԐ�jAؐ0�L!�îm��+��X���T��XŔ٬	҄7����옦����US�G�ji��X�@BQ�2r7�\���~��
��f��Ѩ��9'�+���>�=��/m���]��r���Ax-=���ly�}Bt{��~�&�uw�(_q��;�Ƒ�-8|)��S����WB��D�?D6z+���%�z�#X��{v5u��q�]n�m�X�U���"�:�Q��c6�)H�lpR�X��0,���`�p��-��$Z��<�j�F��àr����rpQI�|-}^���2���3՞��̩��O{O���eh��(���>I-Zb
�`�ɟT���Q���:���U&56��s�sh*��1����k���/�l'��p5y�-#m��Q�Zk�{G�	�{wz�We,g��Z���VZ������������E}���@�}���cFc��1���AH��&%�@����k���-�	m�b+�}Fuy�Ӌ�Z22:�"/���y��Zg�k���$�>���+�U<�q��^���`�/X��,���ň��Ie�y���y_�C'l�_T�Ơ焨!�0	��x����ŕ�Q�c/B�WU]qX��t���;�jxCǔ)��ߵCzY\t׫]���p��"2:0[�?:@��߻7��I9&�gyߟｷP��ܤ8LcV-��S�X���7�b����vj�N��Uz���j��q�`4$���_p��s�����p�g�j�Y�t�8�i���}^���2�6s#�g�!J5���b<�,`"�Ԕ���HA����U����/��h�}7
�j�w���$�< DA������~��3���v'�1%@|z��[)��l��M��s�h��o� e��*z�F���[��aZ�����\Sc�O��u
��X�ܑ~Z!j�뼪R�O��Hx���-zs��S�
�R��a�D[ ��}6.xN�^�Z/j+������b�4̽���h�w�9'����1�j9��!Ej�:�(��Յ>���nu �csk�މ��o\m�)����z�4�L�uѵ�&��_�m�8:�Jƣ�Gv���jp*�cr<�6��o �9����w_E�d٧��|e��>��ￕU}��#���˂K��&�y���X�7)61�X�W�v;M����G3� �a
P}��P�̡���b-Z���c�{⺦�'�+Q��u�9l�ܤr�5*;�쨎�9 ��P�Ws��2:�Y�}��0^��hI�z(T�o��󬇂S�3�sBU�x��U�avTB�l��@��ЏA���%o���R"���)�kO�͹�z�hDm}�M�(PF� ��v�q��]�'v_נ�t=�&�&~`����E	�X�}[>��T!!�@t|�.9����F�1"����C�B�8ȿ�����n��,���79���i�]�ζ�S�)�Ǖ��]ލ�5j]q/S��Xbڥ$����k�����QL9qN�WL�B�l��q��ut�G�V��\�!x{i�w��E��`���3~7�]��d�}��K�Qv%���<�LxEx��ޯ��]����.b�ns�!Ōj��s�O��,���o=@���:��{����8X����=_xM@~!�{=!�;迺e�E��j8۫�)m����'�cMX�v�D�e�L�\EN�1�:��̽����6�u����L�g&����U�A�F<ɳ��E֓�pW2t@Ώ;b&v'%1\������c�Vz�O-Ζ�'5��M�,S�;Z#��wmlkG����k���ZZhZ�s�����
��F��}��'S�񎬗q��w��zrp���L�1�F\c�Δ���2٬����y�͆ǻz=3]��!��q���ôռ#'�]}9%�O��ȱ���v
�B6�р���'6�,Kn��6���{���D��|��Ͳ�D�}������6}?��`�e	q�W��5&c�1Tm[��Y9J�s�G;ULb.:N��g��f�F�3C���p&����?x>��$̚)��`�jl"(mMBg>��\vv�衙���f��C���s�m����&.�Vt��' X�5�ܣ�c�f���i���<��W�R�p��J�3�6z0y�Xj���Q��z&J����ۙ_��37�#Ӆ�0h�P=C��&4�n�O�;U�G��t�+��~=���H�R2 d�Ʒ89;F5��1���~�����eՇB_��E'c����;~�bz��d:�2�#�I���Vc��G1�pbB�f�h��������и�C��8����<��A���n��ٙޣ~�\:^�f�C���p��#�D�68�["Ib��'��^��� ³���dJ�1���v�ƾyEÚ3���ЭNn.��P�VD�=�MۗWn�!��-dv�h�)T�He���^hۭ�Ҫ1嗝Z��o��]mq�o�zs��t�/Si�Y
��'��;�F�t�1:�\��L�\��W�5�mmm�c�(�DD�C���N�n�bE���S|w��n���~�b����K�[u�b/�LW�}́ưʘ�n�D3n%�n[w�s���X5��F���8�_ϧjyO�ڿ~?bbXOԄ_ɪ�5j=������9�G����?��dhi�p2=��[5;;� ?���
ټ���v1l����MGq��&�=����^�~�W����.�DA��#+�.7,ͣ��qީh��}n*����n=C�tZ��ګM�B�nm�U�x���{��:�$����*>��TFXe�;2d�K����xeg��ޥʆ� �i���cS��̞�@���K���O��DP�p`E��wG�����jlF�z�!���}�n�58M�ƅ�`7�����:0L���F�(5n��Lvo3^՜<9��RX⯮���ם�Pκl��!�R��{���H��o����M&�5��rt��S���x� ��#�:}E��7�6�ϕ�Ŭ�m�c>31e6k���ܻ�By
��}ʎ��~�}ޤD��'�,W��a���Ǽ��o����(R�E�Uz�c!�+{��٤�ae��E��k%��-٘9���cy����X1�������b�-�F)K�S��(�eiA���K��r(�l���*�V�������9�7ڙ�R3O	g�{��g]�����}:���U����/�߀�> �a�=m�N"�����WC�_V��p-9��OP �=���y������4�DkwS�ja�_�J~���c9�ԼBϡu=9�r���NR"�k�C��^�`������_p���\jӎ؟v�q��BW�jE�7ad>��^n�/o��E��1�G�I5�w�����0^���$� ����O|���= �ex���5ވ���U0����Ѫ} �!w��7�t-_
Q+ �C�Q���(l���guzqW�A l7!��/�8�Sxw����q.ﳻ\��B�hTw�Zg�@�
E0q�7�[g��}�#l�7��[��Q��3�A�9Fo��Yo���U�h��.:M�~�3���!�2}�^"�����A�{B7]*g��j�n���j.�Ҵ�~�o���ʛ��B���8`��\�Gó�[kR�%^��]G��0��a,n�:/��S��T;Ƭ[&_e��պlx��rP���aB���+;�����~����xw��"�s"�/��p�f�x�8N�������ս���=�3y&N5���Eo*�/qB�_�.!��i�j[v�3���&C�󠂩t�o��UG�c�(F'�!ܻ�r�5�/�]��fB)$�%���]�Cջz}�h�̇��w��M�����:�����0-����Eh%�B���6v��$願�~�4��*����\��7�Ō����Ac%#k4j�>��kuaPe��ì,ː
���1�*">�ɼC���Қ��l���D�jVs�GЊ��C.���r�Ǝ%,���;�2x�|��VB� ��Pk%�c��S	)���>z�O�WIt���v�C��5�^���TQ�ve��xw8��5���\����Iu)�w	�!�P�c�
�e�}}C%=���QY�*`yׄ*ҝ/D��L�7��ڈ��6��
��x+��6�B����=+�4'����Y�7WoG��K��XI�{;-�t�f^h���0�K�w9���ן+WҕJ�?sqoL$L�h���u;:js�n�t��@L�c��s�p����&(W��F��+(J�<���롈s���xQ�կUǃ nQ�7�;�8�8���̥'gaw�k���v�>r���/�^��'�ٽ��!�f�9�.�z���n��˅��n�۲D��ԁ�'z�<�������Ì��9jr�ۅ�ѕ�j���-�[%�Qp�(`�quv\PfU�����[z�j;��K�����y5[�v �J1���:����Kl��v�LE2�KQ"��F��d�7Xa��y;,ع�]�*rͮ�������KR�*�u:�]�n͑�N�2�ʃ�6��2Z�����2�uv[p��T긔A��4�{2ɘ]����C��a�f
�̅c��`-���Uj��W�'s����8����3�k��6��ot�)��;u�	�&���-�2��b$lIR�-�b^�)]l�B��n��֭����m{���&ꨱҥ�	����c�{��/�������_gTnKTT�uc�#Ί����]��^��f��Dq���j��Es�M�� �gk
[p�ef��
���ͧȉp��u�f�wY�ne���u&l��n�a�8U�=yV�,q��S�O7�g]�1Z������ؼ�n�*�l���5�6n�l�W��o-Ve+g�)��E�Ʈӵ���2�aJm�bn7�ʼnS���{�6��o�`�ŧ�'P��hӊ�BMͽ�2�7��r�k��fNB�T&�us��6�yp����:�S�Ν�6u6e�}6V�+9��0b}���ِ��=�RV\#Sf���ұ���L27�;��ۛyʯ�-�f���m���v�̈́Ǣe�-Ću�Og�����BA��u6��R�f�Q�|�����st%�nޝ��o�=oqr�j��m��R/Dcl#���������27��m�J�Z�Ӥ�n�j-b��:�t�����n�̊&�q�k�P�ծ���ԻȜg)%�>��Ꟛ���i9��H$~$��vVaUE2�?I�£ò��TbE);��v�T;�8������ʔ�p@�����L8%�B�Qt�,@$�(�hF�q�A$���>>>>>�EGN�Q(:YE$TR�.�yҥD9C��Al�$�I��a�9�$'Qiˉb���q�$�9/sǨ�*��y!E8VEi�r��k�)�\BԊJ�u���$�QK:J���/��%��	�p��S���*"C�*t�c��-e��'��զ�3ֹ��Z�I3���:D�y�h�d����z�*�y�.�gԻ�*�e���l�*tX��TAG��J��2�,�� (�C�?���$���9��H�!Њ.hUȊYfH3��0�e#���2�D��pYzlO���wR�XH�
�8s͡��$�jT������¸OGv�+M���'8��F�l�K(�1�9����
���u۸�p���ͩ���G{@���1ěMO����c|yV��Q�����Ѓ&s��DMȢ�"*�rgL�]��s���ba�3g#��
/Z�!l�HC9W��-��f��|p�✏k�wgz�U����s*Y���H��#�&\���W�ءN�+d���\��-i�1eʻ~kIځO0��-W1������A�Cb='������,Z��26��SwdǄ��gܮf�"���I�m��NT+�I迚��-�?���:`|���F�Q���e���x}4��O� t1�^���ړ��H[��l?H�6�iXO@W�r{^�@�)֭�D��D��T�wN�E�b[�p#]ON�#�i�Q�?eDr7 ��=�<P.�=�5��A�6b��\fB;���K>�����Բ��?7��e��rKXN~�h�z��᧔F���:�dDR�ѡ&���na�ݑ������H1L���p�{�;�wOe�O���t!߇���]4M�bT��.oN�ϴ��Z\�F�<�K���Ħ7�@�-���bC�}ԏ��_�[����?g�?;?|�C�~�cj���Xޮc3d���N[ڹ��O�ҭ7��Y>t��R���i��5U�E�3)>���=��g���9��x1|7}�Z���a+���	rp�������T�|s-�:�����Kv�rv�eU�rEm+|�4��񌔾���5�N�B
aF_��O�:����;�TN�����z��a���RA��kѝ7�1C�A�	�Tl�C��W}���^<�-�"�C����=5?K7�9���#�-�!�:��k���fǍ�Tg:����������<Ē��F�������������%Ƿ�1/�j�������C���@�$��xw0p����2���<�	��A�o����N�,t���5x7蔼�~+cj��V!��~���زwC��AF��3����#�.�ފPΤ���r\����v�۪��]��nf���\+m[��ޮ���rK����1-�F�mp��/z�^�g
�ގ���
`']H�A+V��S7NS�4-������7���v�	�����{�-	����ig���=t�m���s�����8�8�g_�f�FƧC��\	�����u�(�3b�5�CP1���BKFɘ|}�����3<��7��Ó'=��>'#�/��-�/�E�G��~uR/��\�:F���g�uؾ/*
�ҕ�f�l�g�����!�����~Y��������լ�=������:�T4�[�����`A}#��:�o���&����32�a�d��.Juaې�1��u��)b��J->lB��Өe�p��Kш�S�d�]g*a�3�@a�#8Oe�j:="�� �}�|>� 7�5�u6�'�"<����!���b:��b:��Lii>K��o�_־����9��2�k�χ8�ƣQy���9��G��u�*a#8B���\(����#cna�4�qʡ���q�]��ٿ'��Ȅ�Up ؠ��sj-�.X$gÌ���zx2����w���z���Ǌ����q��P�wX�4<����N����D8�����qt��`�]�_]��^2�0ڷ�o�A�G��JE��F�^�z��3خ"�z���z�*���ь�`���;�]�@��wr��u�|����B}Med4j�~�����!x�9?Rڅ��]o��
�1���1Yr�ά���#(F��3���z���Ӻn߮��xl�E��ؓ���n/��#^wBt�Yc�EG_$l��}>��IV2DAa��&�q�>�6�X�V�q�plG�μS�a�={q���q$X;,F��Sl���2��@���+�b�*d�������\����Kϖ{=�"*wsiک����c�Υ
/�\6s�3O�t-�N��Z�7���u]0���9�q��e�%E�� ��w?Z	^���%#�b�#��`k��{4���3{�,�ǳ_<��=�2҄ю�aʐ��+��W�����z����l��2�stf�Ѷ�k�Hva}ĚVc������Wa*�m�Ӽ��y�� �@�?��������0'��Pڔ!X�Q�"����v��#!�})�o�����%�Z�wG��S>ܞ��q���ht�'�BJ���A["��:���l�t�.)�#������Tn�I��ځ�yE�}�5`L�4A�O��Ԕ#���sl�YB�����T��oC��3N�-�z�����޳��}������
�&#��gO� �_��d8�lu��x��1�x�+v��H��<�Q�x�"��v�X��Ы-��Q��E�ti ��T��B.��aSrU>�wVt�����p���Sӟ7)����E��WE��U"���S��ڍ1�1B�l=@�wEqJ�!y�u�<������W�n�/o��C�-��5�[N
�`�����1�%�:A��v�Vz�!����Q^^�������x��HͣU�W����!7p�yE׳W-���{# ��$�
EV��5&�����5��qFzqV7�$
{���#�ٱ�]y�笼τ�{��T{9�L��k��H�"fSg���NFv�Ӏ}6K�i�C[��^��*�´��/Z��˻���8�����#�w�g uZ��}���h�v�F�	�[�v5 ح�	����u����{�̭ZeJ7��b��b�a�N��qMK'�5����j����:^5�;��M36�/1��8�6�V_��@�� ����Y�_������7�N�[�h+�(d�&���>�N�>��~���$W��f�w�}KᰵҺ�E��=9��b���-�v��iY�!^�A�%�ƙ�+ʶ#��U)��;����S�5�1�"�ŭ�����b\{~�A�ƨS<)��fպlx�������Ī��Ç�OEx�@��Ŏ���Vs���b�,�Rr�8Rӱ��ʎR��qFz��W�>�g	��$�,EH����p�޿��)Ц��[n�����9=�M�~��.����[���(+���8 �' �Gܨu?��B����/�:2�D����+��]���v�@kn��0�z�J���$F�f�Н4����tm��ybG�#m���G=�Ra+rE������8�F'*�����H8�Aځ?t���W;:d<���+-<��w�hw	�uxzT�<��f}�ړc��>�c��|u ��A�_��W>�Q����y`{�?@���W�
�q��7^�@r�zp5)��ڥ�㜨��p#;F�זK�x�Ӕ<��<7��\�67{�Wbt:��a�pP���JWU��_JMܱ5�s(�˄_8�����RH1�a���H3.��hib�d���n�����s��2���[��Q[	����Fl���K�b�*�{���41j�җ��l�:�\��9�8����(�M�N>-:��~T A�3���hI�.(z�#|o}Ր�S�9�>ϒ��Ʋ���F]߳d_�N��d��~�똎c�U�x)tKF�֟#�m�3׻B#hgSG�ǥg��W<����e��v>SR�9
/�I�]��2�P'A�"����/�m�Z�y�N�6���!��@�)��Ć+�}fh����=�0p1**+�=*2Ѿ���^�z(]O{{r�����(?�V��{���E��wV��v��-�RA��X�Dؘ٘9�١w���
�+�so�a�����S+�\��(�uW����#�-�!����Zk��k���s}���I���Z���-֙��L��D�G�&};���ꭀ��no��s�s�t�8�j���d����4eW�;�����t?	�0��p�!�2r=^P�EPl��S���^I5Ial�{��d����UÖ����L�����!.la�3Aϣl7<��'�Wa��3>�6����̯�+pop�ĸ��4Σ��2�>�p�T�㾞�tX>�����B�����#\��۱v�/]��'�ͳ���j@��0�<]f�4'ϣ��;L�	YG��R�j�ߦ�j lg����J��
 U�\�l�K���x���6��̗�^5EgP�$�Q'o��mQ��mw�3�Xֹ{�:�AwΒ�3�J׾�=��|>�#���  >�{��kΧ�@���ʌC:�"��v��S�����u0=�<X�lPR�ۓ9����
������(R��4%Fz�D-��s宦+��6�^f_�f�F�:>��3�jC���#;�{�Da����1��ة(q�5�VMGh�wљ��4g��'�N{���7R}S��Yu
���ގ4蛏0�ɉ��8��@=Ƅ�g��ףq~��p�Uq~����Ři��27�С^��Frg���kJ�te(Q;?�����]�GW�T'5�hv��9�'ؼϜ�s����{�@�㱸XK���F�5�~�:ę<G}0 ���\(Ϥ�yb=�ߣ��͸��U	Ly�d,eU�xb��nmE��_	�OC��Y�����5z��O!�M�x��O��q＼���u����D8h���q�Xe5�=x�'��;)m��p�8�P�Pd�)�ףp��_O��WV7�q����1U1Y�x Sg<�T*��:�7��6g_킒x>bO��n��Z*�~���Xk����q���s���v{��q��w�et����6oޯg5Ή�Fk[��:���4��溵�>��Gc�f^�Lk�>���I��o�ާ^=�p�ۛ7y��5��r�����鲂��|.��In����7����r�0�RG��ݜ�@��?��������^&���.�~�[�������d���z�%�S��r���l�B�{�;�
Ug�ǵj�l���GaqЍ�&o��mOx�/�\�y"!�FX&�q����������F��f����v����0�R6
���4�OU�x����?l���5��YE��tkug@/���vs�m��b*V���B���GᲉ�y�۱�)�da���9�o�x����:�ʵ�����Ó�@�ڔ!����Ȋ��Nd8O8жl7��mwT�>�D:7�4_�b2��xzF�ђPg����[ �-y�ƌ��`j�.SU�`c��[���C{ɍ�v��(7�r�,/��O̡��\�+�Ŭ[n�7��k��e�N������h�!�bt�k�0��ƱO�,;�Ǡ��ytS�Ë,�u�t굍��Au�o1�OH�iځx��`�{�僱`q���@����v:Z�:�YF\��p~����)�
wP�
V��/��l�n�)�WE���_)9B��l���IA0�	̻x�_�kF�Y����'R��B�k2m���ؤ��	!s�hf�0}fѢ�[��;>W�b���D���M|8ly�Y���(�sT�t�<K�MP�Z��nt�˸��KrV9Ne��V�L�޶��Y���G����W��BK`ء�s�v��/bR�쟾��q_H>ӷ�Q}��tp�n�������N�k�ɕQu�ꏕ���>}Ӌ��K���?(��_�m�C��wTGW��@�e�Tc�oa��\wu]��L�e�<�9H�,�I;�
EP���5>XE�0���C�����k��$Ũ��
�-��X{#�P��b�X��s���`�Aσ�!fW�,�h���$FǞ�q�W�z�w������Q��j���6�/����\_T�Ơ��H�["��~7O���Vo�0�ȼ~�����ŕ�.�ы��>��;�����i�� VTܕ{7}�}�F}^,^h9o�ם�p5�ᑊF,j�@��mл�� ���T<j�3z�`�t��y��x�C,�gj�x�ld�����S�!�w��"��tX,S���V��q׽��R�:�ibv�㱸e�'E�	-�느�6;�!
�W���-��⊕Cn}짳<�}���Ѹu�
nn����t��?hZX�̜�����o�W��>�@�kT+���*�6i��u��%ܯa��9	�5xo�#AW�]Cڒ�
��|���V��n��"ħ���t�[�Ʊ�����EJ������ҭԻsP��	�����Y6��$���m���f!W�s�nj˫.b�����qX�}}w�Ϫ��W�}�}��<{�䃘�h�ٳl��r�h�q��E����OYQ`�g�İ�#��p�������Z�}T��1���v��$]���I��)�z19P�J���I�Ё?pՍ��]�'��E�p��=�5�1J�E�/X���I��{���w�3������1��C�ǽ�>Cuy�8������uq�+�FCϥ��]/ǾnR9f���Ҝ�r��Q�y�����k>������_X/���K�FN�۝.)ۅ���>9(d�lbQ��jsz7�s�~�]��ݦO�P(����p�	�yF���~][�����e��ܯ�W]޹�+1�<�t�LpGbF�Ah���`�
�h�`�4"��k�^q�n�}Jv=��ݟ��w���v!׶���lĆ+�Y�~�jO`�� 1**.�PuQ�Q������k�1�1��}�}]>Ӌ�u�Q{��"�/S��Xa�RA��/���1M���1�+۷��2��e�|`��-s��忯��7q�-�!���XMz�?����ϫ�'�X�RX�����=k^����T���G�V��l�q�7
�΅͵��R;�����{��iq4�m7���f�q��5,�c	6��z�!.K�!���m{�f�������oP�GA]�]�YT�$��M���"����F����]���j�_3�V��3�d1UƂJw=3I\9�V�L.A`���24+�v�!V[�&��*A����6g[�"_q6)�@��sXr�k��,gZ�ǵ.%��Y�{r�݋�TcÕ
�Uw3f5��H�n��e��0�����+.�3lM��᱙ne0]Ö4_x���Nt3z�|�3}Zr��G�kَ$/_@�7���=�MD�^�W��]��i7(r�!�A�EH�8�g^��Q�0�*)�kU��f�Lۀ�{B�K�[�������E�R�0�f�X�:����.���;�M�9ܖ� ���_�)2=���u���-��uꕺ6�M+(w#[}#�ٔ-�Xp��cl�g@A�#m���&�㲹܊����w����;m>��\h��/w�E7t�Ծ�U��ڶ^[yhWJ9��A�a�_V�kT��j�e2I��|e��h�m=&��E��|��kʅM�'WYT9ۘ�#�2.�z	�M�X9+���s"3�W�+�oE��'%LzD=��a�o���%3��Aq��g]��\�
6�T��7l-�Y�q���ɵM^�%�U�}jlؔ�7�(��)���I�O��ظe�n�u���=A��u:�<��r��h�r��y�f�x�M&F�;[C�/�#���x���S�vhh��A&̍�˳lQ�nN���C���km����v!4��k9�D�v�rI�w�9�l��\�
�T�!$�ȸ�ҥ�dW9b���i���m�
<�-q�o;�^�[͆��b�Y��q�so�]�ݮf>��j�!�9�s�R�r�z�kM#ܟ*����Q�x�7UYPs��N���<v(,�sQt��&É��t׼��1�L̈�OJ/�}6�7\���"p 9b�Y)�@��������S:y��&[�T�����U��tʯ�8�c��:�|i�������0�L�S�ͷ�pt�P:��-�q��Jھ�	������B����G+`ׁ��"�U3� NC7�m\����"ѹ�l��|����0?�"�t���X�:Z�N03|Yp���jH-j�U�X��p��+ځ�fV^��&��F���(�۲����Kb�v�Md4��Q!a�ǜc)��*��p����wb�4k;/��P(�e�����8��p�
�f�)�J����v�����Z�+
}���GZ�).wy���Z;�EZ�؛v�ٱ0��H�R6��y��EƟe�vi?N����akkD�ם�l��2+	�nY��+�7s��l̈́"�c�#y<��t�O�o-t����#MvYܫ���ދ��F��5�����X¤sr�n�ÇUgn�� ��:���	(���Ȕ��s1�gJ&'(H+�Rt�L��%NF��-����>>>��vYQF��RY����~\�dM�
���w )�h�L��|~|�p��H��e���f��[(uO?'*L�(.Y���P��/�	��Qq�Q��o'���L��.��V`�\�H�J�$�VQDEˡ���(��"����z��V�	�9=�rϙS���)ss��p���2�b%@TuA*(J&]$�BE���V��\Ӆ9�"�u�.�N�Cs�̇�S0����.Q�߂ܴ���0���I���]�/B�ps�QWp쫷jS�P��ӔD��$���8��E�p��i�Y�B!;��6��*���+��<���\"��g�K�t�MZBI�t�TB,��n��nLL�H�E9SC�wƆ�R%a�σ(o���U�H/Olx�T���v�SZ��ō/s��%���d�Wk���&���-�}��K���:4��b>��W)o�r���~�e[+����C��6�/������mЫ���qٮ��+.^Ռ����*�36�����ӘX�xe�|L�
��7����;�A�}�r���X̋��~[��Ӛ�D0��k8up��=���,�Y6<,*qv��'(D�#����i%/��h�]�7�VzA��K���E�s�m��P���>4x�8�T����y�g^|[�y}����B��tY�Dfۈ���`-�P�L�K��g�L�)��w����|��}?���{����g�����b~����n����r)�Z�b�����<�������V��7��&�E�CƵ���q��@���,q�5�VMGw�lZTћ�l93^��)���kr�\#|�e�(��c�ɉ��`��:B� ��/��ʑP�R��Ǹ?z'R���s�Y��7ҡ{��ӷ_K��r��H��k �#�������%�J��5Q2)e��V
�>Ѫ;c�X�g�@W��~8���)����P&;�����/���{�2��R�O���|��x{��'��Z(Ю#ۼ�K�h�z�nn
�r�ܔ-�s5T�]3s2)Ε.ֱ2��@�;�QTs�K6fC��1-CGY�(=Oh��c,��uj����WV�b2��*�vfP����?���}�
����5���b���a}����[d,��b��nmC�\hG"G��9�^V�ňN&���<�?���{n��Y�b8����:�bۨ�D{~>�����Lzp˪X�7�t'����K�2Ƌ|`v*{��]L;kٽ_H�b����\b�n�CL҄�=Y�!v�{j�^U��ō7
���d��T���YY�W�ݦ�5�Ց�D�*�T�0ǅ�r<*����<�\"�^�Vk���W�~�&,y��_|�׺r���l7и%/�q��i���������P㱀-��r*���S�>���9%aÑ�0M"�rG�' �]�lJ��aꭅꔌqb��Sl�z�[uJF��^�뜒���4�}C�E߽�%w���p��|�J��By�I�;=OA�$�l�V|v1�i����z>�*_�t���W��޿D��W������T��H���w�z�!�LwS�	�!�y�ϫ����N1W�m��yX�9U�6O��
="CV��A�a]��L5��u�f��νE�De*��˴`�Y�9OaF�]��{9�ݸ���'lϲ�}ҽ�ww����Q���8m�o�d�+egޱ�Q�U��Mծ��p~�N�9��(%�X������+O>�Wp���H|��Nic\<0M����/wG!/&V��"{��D��@���p���I�9���t��B��Q����)D�600G�В�wsl��_�Z�Z�-�}nn�"݋/�#�2��Ov���b�l�'J�{d��i����/�O͏�y_�
������'������Z���o�1GJ��;P/WB���
�v/�8A�"�<��>r�
������C��r.|6)PQ��B�����}ON���FS��j��j8	S�����o���6;<�o@�����P�{����V׺���n��}W����	�B���_!b8Т����q�v��i���B���R�L�����Ce�uDu/Z�c��0]`����f�{_a��f/�tɇ�'!�H�,��D�
EP�>Dĳ����k��*a>���K��9��]�]Q�k�������P��b���;5�ai�U18��7�[g�U�S֎%���կ��3�vT1�V��L�^��ߨ1`4�诲vˋ꜒���*`@�����n�X}��׆W�~�[�v�y]�
ۨ�X\��ZX��~�o>M�H,o\�KM��z�T$Syc��s7���F�C��f3O��|mv�/rDl�t��c��*m�-�[�Y;f�o�Z��J�rj�k�Yg������Jf�λ=wyۇ���׼��r����e[�5ɠ�93"�E[j�S���m�wcy�k�0��Ó4��:�EEþ�������[y��`��$�`�H�b��[���tY�)���8w�X�e�P���i�G�<���`�yE���rN���X>�����W�F�:���8J�����bw�^1��p.��lf	�{�cp������lة3w�B3���}{�6b2��O;��;��:8�j)�M�mӁoH�R��ؑALG�e�|o�P�y�3���}��w�]Nz�؉Ziy�4_��7���u��
,�dİ�8n��*��CC�����N�C>�2F�[�-g�m���I�m���
�R���I�;�!U��.q{03~����0?�蘸bP�����^
U�
/�z�g'jN3�US��X~��cP��1]0ssŪ��9�"F	�� )�A��׿WZ���[�@�]OKe#vc�s��4xyϗ;��?C��!��@*�P�p�i��l	�'������*�y��n��T��dE�����O��m���u�x�3ѡvTB��T�G Ήh�kO��6����
2�S��>4]���w�C7�"����L!�y	�ȼW�#�f7D��Z������MA[7a��[�q��M�=L"-����ݍ�7���\��jj�m�e�}�C'K����%�^�����G6 ˗9l<71Ȯ�<�
$�1\CF�E��۽y������|>�Üw�����؃���_�w��,3��w�Q#������Q�	��Iߝ����BS�^VQWS��<wmz�Jیw��[>E?|��U�@tls���Ć+�Y�,��3rzǦ�蓞;&��q�{�q��:4Y�ss������^�X�n����(
����$ͬe���������@�9�0Ś�?`~0��L�k�*~���L?w�Bw��b�@Q�؅J�B
9�m�#/����qc�{��pPu��6e��`�`7�k��S���.a���$�c�C`c�[����.���Ӑ7����xe|L��{�������{n\gҠ��%�Xz�	��1�,i��g�n�M[�'��{�9��'()�4�G�y�X����`��{=NѯK�ǔPB�Τ���2�D�𔚡��ڷR�]������}��n֟Ms$�ɞ��X�����U��B��`:��)u�l�)�e?q�m�t��8�G�x߬�	��~�5�{��`�?O�	q�S����V���.5�Jq�n$$c�i����_�+����n�Z]�j��ɍL���Kc2H��3[�0�
Hbi��>k',���y��g���{�_g&�m�g�%%xb*�=$�Wp[9n*s-�Al㫊��"�z!띅���ѻ|���v�iM����۪��邨\�wqj�����U
��A���l�,w�W N��@�@U�=�~��|z�j;Gk���*h�c�*"��4G{�ޕ�>�=���ٴ|H�
h����0$1�:��LC<��W�P�Y�=[ې^���>�5��#��Y�n�w3�8LF��!�$ ycKF��lʸM���;_g���Y������P5�S��p%���}Jo����bLu�t�Ž�m�9��7e��{�����������l;���po+��m���W�b���(����E�O�k�Ox.빕`��4��1�C���~0b��i��)��s���1�1�`g�����Ώ;�1UhM�P��{��2���(h��b���e�Tҭ���˽�g\>���z��;a�Xk������ϙ����̵��W�R���dϰy����r�x�o/��v���/��m��'
����]F�^1/�D(��!��W�s}YE���m'c�d�(��#�#{>Y5�=3���~����[<jᄥv0-�"��!ÿ����O{��\�y�@İ�z�ﮱ����?~��p�����uc#�Uoi{�e�ȯ���ү�!ڍ�9��G1p�)PIV��V&����Ls.��ͽ�����{1���EL9���И�Ɯ�`��'o2�"�Grֶc�u]�����U%y7��jL�s0��־ǽ�#��?��(W��M-2��:x����1aml(��Rѳ��=9�)�^�ȋx���r��\��o֌�g(���뵶��A``�H�U�T�1c}F8gJ��4%�E��g��n�9t�*��5>�^�So�<}��v���K�S���^�� }�"�ڔ!���0�P�Tb�u�p���:�3%ue�Sy�7�Wc
����ϧ���'�fh�a��W�Pg����["�����"�3)[�D�M{��ӷ-i�<�#�~�觨���m_�4"X!�4(R�}�6���lA畆o>��ި9�b�����O�Ł�)�X�(W�=�D&�/��P��<��������[�٥�6-�6����<��ZF`Iځc��U�[���(�|8�	�@�����+\�׸�{ﷳ��nʎ�u���v1�t�G`���nR9)�D5bz�t��hŠ[��>�V���"�G�D� ��{u��mQM�^���S^�������ef��\��sHu��#�ޜU �Q3� �.�3�{=u�}��3�^"�i�K���W�j��<�>w��lzP�u6[/x���8��hf �P�
욡���n�#e�e(���J����<;M����yG3�xQ,���ԟ�xd��R�x�2�^X)�Ϥ��v�-r:S�����a��ӛE�Fs�j�]:i���u��eB���(P�� 1�Ɩ��������^69UZg1eyMQ'��hy��,"�\�WC�c�Hc�+�]�>��{��t���܆"����XZ'!��k�_�"#��+�#�R�7M�^�z�~��g�./i]ϑ���+M�l�E��a�������-g�>���'Fq���4�E��,Գ��g�ahU�Gٕ,��מI��nC�al��?X��������]����t��ϼ�?�����>8p2�=R+�X�[�ۺ���%�>�B���W�Wʖf�w�ϝ��П�v���nX�=��o���U����E�������]��8Yz�U��莘Oѻ�=-x���^��{�cp�;����%�|$���D�0,z�p��LK�cùD_��Ǻ��^����#��X�p,��s,��;��$K���H�b"7�m��H�}�yyM?��<�δMw��p3������w�{�1֧�����\uVg)K�{��^��o
�@����ܱkے.�;�7�q��ʄ�ϩI�Ȣp�r�槦����f���am5Ts�cZ�O�}�ᘍw�y�7�4<(W!������(����oQk{$=��Pm+�%юogg�_ �!�r�ƅ��V�JNR�-�qEl����0���P�@��o��:�� ����Or �jQ�4^]>��]}WW_}_c�>l�(c5�߄	��@>�E	Bv���R�@Q~K�3'jM�t+������9s����-�]®���5��~- ϶A8O@U������u֣!�	n��u=6b�[�O�P#�磻���o�����u㼨���W���.����;��:Y������~�W]��
䧶� ����������N7~��uX�_)pR��Z&'O����F+�7��36�Jz�D,R����H�Gy#_�=�	����GӜI��<(K7�{$k��Ɓ�%��$;��j癖sO4�`��ߠ:<�`�͉s�1�ta���Msr�c=���ʾ��~��|a��K�g!����8���E{|�"�w�@V��1mR�ʙ�J.ȭ�n�ȿot���j���U�����S&Z�~�?N7�U�|�Do-�!����k=�=�^�s~w�B��ݞ�͹Ō.����_`##4s��������no�嬚����F߼��<=��5\!��Ul���a�v��O�Zğ��2�W� ��m�����?�e�>w��(,oۀ�S�yH׽)���l�x�Tk�f�9�I������gp}%�%nX&�J�=�$�N���m�ۧF�m�{m�ht���BHr��|7즜�b���W��;��l���R��3n�
�VT��޹��k�Ƀ��?�� �:�i����!�*V���������W5n3�x�/�9�P��#����o$�%��g�ػF:2�m��PB�Φ���2���f�X�
�j�dg�Gz�#�亏lϙu/1]g���9�*�s����LE�	]QV��m�B�t�)�e>�߫`lw��`�X���b;��ƺ�}?P'0_h�?H	q�R�-�vע�Ů�+�e#l�W=L��p���Q��o�1�X��a��A��@_3ѲP�(mMC�ՓQ��[Sg��?C1�pk�֔���ƴ��6�N{��|H�SD���	cdu} �ܣG�ޠ:�W/��s�Њ�{}E@�M��'��;�qlT���R���[��}M���H��Y|���93�艔��w�1�ƜFx�SU�p�����?�.��e�߁S���X�]0 ̸��C���¨C�,h��:=��s�О��m���U\�����8ap}�=C#ܱ�T���;Ջ�!��`�1xt�W�R�Vԍ���#���
�UhťQ
 ]�3�-�t��<*��w�1���6E�<b�:��T�41v���r#��������:�io�F��U��⥶��y٤t���8�௜��I�]�"Օ��]�I����t��	@�݁��8��r���_vP��N�w|�Kr�XJ|�NƥVS4�N���n+��FΏL;�L���� 3ޭ��Ƭ�e����I5gZѻGf�CZe;��dj�s��e[z٩ҮWV;9�����R�'h>v)#{d��X�%#V�_�Ӹ�	�k�ro>��fQb�o{�E���e�l��gi��:� ��u�&��s�ȕ���xa�cp;�])� h9x����fg^�yQ�H��YF�J��ͥ��{o�2gDu|i���0͓e;@�S�XRm6��p��v�[ڳ��髡1�p�5��zq@&Pv��gUG���"sxK'��
����u�ս�QWP��9��Ci����yw1��ӝ4�ui�5�@�٧l/�$kH�R�X�׹+۹1��p�6WJXO�g���4�.u(�"E�Tu�OW)W�F
"J�QVۋ!��3p~�������������d�NɁIt{i���a�[���P���ܬ��7�.9WƝ�V���}1\���ք�;�+jsʼ����t��ӗh���^���w=���ҿ&0F�ũ,��G)��f-�pUM|�DX:Cڸm��3��z�=t�Iuf�(u�#�ܻvCq��smb�N]st��C�[�R���u+(t,&��R��k�5�1k��9��*ua`�pp��Q�Cs�+�1h��ŖE>Afc�y"�{/���\]�w<��#���˳4V�*[�t�j�G��L�=�5�E�ɂ�4hEV%�2V��:����ooM�f���k��a��IŜYh���4t�۶����4�F�b�0s�䀌cw�B���H ��w�X������L�NH��Va��x�����6��켢P��-���t^R�R��[F�d��!Ά�7a��5l�3)T��U�ؚ�&4�f=!������wu�A�ۼ�D�}�8��W��ŷ������,����J����L�ia1P��v��5b�r�����E*�C�L*O��Mi}�MH=�3�mm�]=�W�iU;�%�?Q7x8@�e	��hu��J"L/�o^CBʭ�[r��/�h3C��,岂o7��]*�R�ꡰNL�PN��gT�l��җ�5�L�����|A},&wn���O���t��^�PI�W��D�-�2a�׳5��M0B�&w���{N�8�omܷKj��Ll��o�=�W������!3#YVh�E�ޙ�4U�'nB�^Xos�o.�-Y�29��̋�9���kVImr�g�:pط�خBBv�2�1��Y�'G�IK"�[۳���S�OZ��(�fs�;Û����$�t�Ƙ�z�P~�����9�����|ۺ8�hʔ�&�{L�u��i7W���j��Lw�y�d&�E˲x���|}�2�?RL� ��2˗I��<�ț�N�UvR�*&q(��㓊�q������~AyU	ıby1�p��d(m	��E�(�gd�j�6$�;��AT$�2�o3�N*G��(�*�.NDZ��2��97.��.U/s��(�e��݈yM��2hM9jS��*z	z��g �*��U'nv�N�rI;mQ4\� ��%�$�yqՎN����듪�T�s�S=�(H�؜�I&U��8�!� �^v���DL���N<�Nu�!޹��V�xfM�t�\��a�ۑ�z���F�w2�Iu%1+VQ��z$z�I,�'*��N�r2(���@�P��d� d�ď�/�#�V��ǯ׹[���Nݸ�w��8s�˲vR��M�Y�b/n,fP�!��S�9���cOYŹ��ܻ3��U�^UdRUӌ:-�+�� � ��<�{S�u$�8��2��D�`��2z(MKe��F�K��\��vZ�{��K�$��ߺ�<=�B���?�ף�$�cp�1�k��d���_�r�&�~����|�s��y���g��Y�j;���\��bXoԄZj��g'k!ߤdk�6L�R=^َ���c�B�r��a��y�����	el�E��Xgc [g�EC���U~��Xr*k�-�L����P9�;��Ψ���0gL1��_ީh�=,CӃ��/���1@��ez&Cw��Y&{��Obp���%���1X4�%�å�G����1¾���e�g�2��cg&��	~Ψ�������w�3��iv;-�W�V��� k�c���Q�"��Tb��ۆ�>���<��Y����1�>4-����=8��}�`h��a��T��렂6Ȩu���DŻ;�^�=��/ r0�������a�46����<hr$0G�VU�3�z���X�w��#fGXVQ��߬Z��P.��O�N*��pN�+��فL�1ޓ�=�%m)���EC���L�MWjS���#��������k���.<L�+�� i���c���
d���*�x�.>зf|4C��Y�ֱ��%��{��{|�lvW�kocO�+�S�}˘�Z|���//k*jnTw2�Yv���r:��kO�����+�r>=���C�D���ݕ���XŅR�3v�^>��Yn�r�ؾ8Aѽ�{n�����.b0�qu���}R:T;�:6ǹXǅ�������F�}NR"�`.���f��e�G��E���Ӏ�_h�'���"<�ژ����Ǔv}5�ֹP��X�K���5�#;�SwH�o�pAT
&x)Ap,���=u�_XО�^�w�LR4=����s s�>�f/�^7�UF)h��c�dv$���"�D�i�@|O�G�`�Ύ�ə�W��3ӌ��A m�G>�^��t��l���T��y����{��ш/,����j�x�>�zo�-�Qk��6ߨ1a�Ed��9%���ڳ�Ҧ�j.�mZ�Zs���u���v��{���~5�<��~�ov�����u�r�G2+:����'dO��z�$��l��G���\b��l7�wQ�`b�nr���߫�+�Z�FZ��m��K��K����6����P��as�Ȕ	!���_�E};��Vt,�0�9�x��=r�c�Yg�u��޲�]�h[At̮�܀Z�{ʵ���_�;�s��o%ZW\!Sw���ᛧnr5����(m!lH.8��)�7\�G7�U���kN8�{i�/d_�Ǯ��-+�WwX�Ȓ?����䟖��^�A;�\/��5��t�8���c2}^�;�,�x���*B�ӎ�oNS���wg"�<� ���C?�����e��5�80�mہ`��E��R��;ALG����D���N��_�,{��#VĉZ1[&��M��s�h�8�á��3�]���ՙw����)�ž����05�G���'��Hp�nX��m�bw�o�q��NT'Ҥ�oy�6�l�|�򘍘��v�?[As�r�O�0
���'c��^|)W�(��c9:RP�=�TP�9Q�q>�jm���C�_ڤc?_ �l�%��
�GO����6����^6~��Մ�p|�N���%B�k5��z�r��9nz)��F�M��� ���&<yF������_{k��q>������������	�nC�]��J��7���u�B�8 ¯����H3�Z9q]��d��U��=��t��y��HA���M���L�;�S_��;>5�>��R��}H=��&��L��|�9��+H3�~.�}��%b{o�e�y�!���b�GF���kaRf����[T�mg�轉�1/f�wV�ͥn�L�V���~�6����^��Ʊ�����*wf��a��ߓ�Ϯrb5�2$.�Ç����I*����{F+�����[�8<��r12��R�;��M_l�3�����?������ȼ��w�욃>���CҢ���[5�t�N/�:({|�"�Ҡ$����<v����g���jج�RA}������3��B�����`��-{*��ʯ��>n�;v�<VM{�Զ����Qǻ�VS���@�Ie��g����(��#"K�(���ֆw����o�`��1/��Az'��Z��<�T�8��U���W�X]>�ȫ2����e�#���D?H8���V�G�1���p���`t����4y�W5n3>��E�� �Va/�#��;���#����
��W�U�Fz���A�Τ����[>�L�+P�M�qpw'c}U�*!.��1���p�ߟ����6b2+�N�6vxCմ`:�L����e �o�~��n�#�1���<w[1��롵�o,��8�;����%����@�o���Z�c�)q�_�EtŻ�2/�����I�w�|h&l>f�_��\	��T	��=$��V��>8:�W�ɒc�d8���r�9�[�ќr6�	�q�ωAM}�5����'�ނ'�X�+�3جmfA����̻n�_�=:��������ׯ����3+@]W��=�M*J U���խ��5������^d���%e��'ٌ����c�;"hV�e��U�u�]�m�i�f���^�������x��sㆲ�R+o�f�ԭh��J�����B~�{����p|2.x�<��foSg� �T��|-���,i�b7FL(����s�9��u��1{�x�>�uL����a��J_�e�>�V�~��#]޿	o[�.x��6����d��P���7�ۘgoܬO_�V�Up|ؠ��\�G����ܩ�X�(��u ��@VRc>��'�J�%��m��o;�G���X�V�z(ܡ��;���pu7���2s\E���*H��'�2�D���&4a�ɩl����+��}x99.GZ赭O{Tn���`>�F��#ZU1_a�c68�V6��#�H�b}Med4s���{�3�Wz��zf}O���)�E����,C�����A�md;��6L��H��w���xd	�ו<����N�p=U��¶o"��a��l�͌r*���7�S�>�Q�*�
���EFtߝ���
����,�|5�Ë�z��`��NSl�z�[uJ��W9Z�\�e�S-p��W��2���B����������-����+��q�ĸl�S4�,�,J�������{��=O0��P�Iw��w�Ӡ�,B�!�C�+[l|��0��f7pV�=�S�Mc�Px6�x�_��yp�Pbb�%onG�a���=b�������;awHF��u4wbiE�;۽s�Q��L����bgu��?����߽����Z�o�����ӑ*���}4�E}%�E�B��������bC;g�-w�7��F������4-�o���OW��}�`h�1�+b��V���>��g/N\�Ld�~�꣞Ba>�s�+��`	VCE��dtPQ��f��=�|Aȟ�!����q�qUi����>��Z"��\�;���-`[n��c�Ŕ٬	҅c�فL�1�|O�����/��l���cq�
�\^�����*��;P/WB�u�]語���V_�m
�Jb*}�;�}�- ���@;�.���T-�.������vp�#��uѪ�z�pO�y�ș�~!��N,#��_)	� ���E	̫ۨ����tw�_7a{+O�e�i���{��=ܧ�6���1�����\E��U �Q3�H3��p$��Ͻu�o[;<* $$fE�櫯k��9�����摎Rc��2a-���dk�4L��U<��4�^ӮxԘ2_��>���ڨk)B}�/�i�	a�Es�'����ϫX'?�=�I�S�|�(}u�T'��v�e
���8���u/��a��q�"��*�oi'��X�,��n��뫼��{����$��Z�%�|�;}"S�����˾3U��<�o���e�pJ�����E�&��K7�t7#U$��N���j�`Z��8�7�Rf���v��{e�j-zXf��/����\{}J1V4�v��_^w�%�g���`~!�I�}�U�4}�^��E�n�Ҵ��P�-���B����S�H�s���d�m�㦽C]���?`���NG~{��c�b\nVw�ۣ����gi�WLd[�m��R�X�][��Vf2�A�aNE2)	!��_!�b��Ș��/ժ;x�g%(O����]�Ӏ�Ĵ�]����n'�kp!�(���e�ϟy0������o+��4q��81����z����)�h�ơpmہ��#.g�V� ���Oq�z��y�z3�b�'	��}�<"�z$*��Mi�TU+�_q��~��c�16�rb�+���#K ����A�\w��8W�ܱk>[nH����b�g�r�P�]s�䨅��P3n��`qL�d���l_��v:��^.������G'jM	l�Ed�s"7����Y��Ӵ�l6l/H�7�8A����@��H/O^�\k��_��y/{�zD�� E����C�+�ck���/���lp6KA������a'�k��ܣ�x:LM����)$4���U�OB������w<����.���|<��W^��l���3j^-O�V6�Y�E:ye��Ԯ���������=7�bN>��ͯ�T�'?x3�y@�r��>nR9g-�E<���9 �u
�0���(���VY�����9���a]�q�βJ����9�>�U��_��q��'��y�(�~���
��#r�ʝ��;͎�weɫ<�;�g�v�F�����ҁ�n/������Qc�I������U��.Ꮙh~�u�SN��n}��}�,5���ѿ�)llLb�������e-�1��b��<���ZQ��)�g�?�Ӳٞ9����ꈤ;Ԡ,�8�����:	�^>��Nx�A���$ͬ�`q�L�ڡLX|a������2e�eT�9P���z�lB��x�ϻ�-��w�ۡ��ۤ#oz�	�X7���3c��˾�d�@ȱ��k������A���+���k�ϩ���sW�!N7:b^5V�}_���\.��8J�?!��6�To�ӛ{�w���n*��6����w�İ��f��'M[�ɞ��X�Y^�FL�W�U��<��X��z�4�G��2�;��Δ����[>S4�}"�7�Ə��^{��C �7������9>��j�rM�/r{�%ن�_Щ������Sc�8)�C��u=�X8z׆zl:�jyt�T^��-L��ZJIoQ��-�����̣X�sQ��bz�vd��r��8�A�R%O;����I�_W�6�g��{{�1I�o�~^5�5�Ls&���N��8C��Q��L�Au�l�L�)�E���Ws�7��\c
�ڭ�Qk�����v��9CO�
�n��m}���G���_ƽt5N�)�Gӥ��ر�}㬿��#o�3A#a�49��	�˨��Ϡ9�%"�����G�����x�,�˪'=��w*ؼR��c����:�9�>$u)�bz}�6GT�oH�7{c˽����q�Wb�R�T=��f��v�����}!�TG�g	��ف�^Iz�Mz<'ܼ��(>���Ra���tv��v��X���t*Q�OCN���l�~������~��#W��XQ������A�}��Mu�z���\<��N�N�9���N���:�����<�e��Z�� b�4�q��&9I�������5� �M�� �7�~E�6Uza�tgx�n���Z?s?<�wnJP4�{�x�}�o`pw.�x�.��X�+�Q�ct��/�B�,��v�hh��+6_�˫�+�*����y�Ս���̭���q6m=�/�uC,�k��F���n�^e��M+��k�����d�Fū!���_(q�[S�X,�op�Z�I�hj��c���:�%LY�Y�E<�t��o;��}I�?^��g�C`�a6�_'��~���=Z�N�FM�;��y�4_�����w��5�X~� ��N���z)va3����ig_|�A�����
����$�_I�~k�Ma�SK�+�d�˔db��'�"������\�~��mY�����R[��p��ӥ6�7�s�f4G���FN�^�J�vw�]�M= �2��uބ<��]NC��tBJ#=о�-���i��N���w:�����a�YA���VFOf��zT�����%�;��77�\m��|����P�������:�#׾�{�C�ͅ�ڮw���u�������^��^�A��ȼ�3cX��~��C\��UsSt��]뿻�;�ܦ^�^����Y��\]u{�q���u�9!�#��@�����~�n�y�o���>�4�WH� �u�@�%{W���:j������[���)]����5s��K�f�㈗�ېk�v�Mytݤo;{S��𾑄���[�vY��7 ��y�6�r_hȄ�v�nrj�8@�c��0���@�/d�ݤ����xvJg��á�"�^0����Vgt]F�/qĒ��C�j+�Q�]Q�oj�z����5:�U4���s���u)K���䕹ٴx�m��)�c�]�;9ES�-W�ډ>r�4��8�����=q�&�V�uj$m 3��/��0�[�p�[#\�v��&NV^H'm��+3����vJ{U�D�+j�慚Ӌ�����F)[�yS�O��I�w�\ʗ���/�9��B��˧Y�+���5f��L��ܷ�qX��l��Tz��b��Աj���ٺU��#&�9���̃hۑEX���ٱ�ZF�}Z�o��]����y�����\.y��%��rY�����qop:�������7s���Yz(j1�#vs�ʐ��N��G:�n�%��(���`)�N��5lW+�
���U��t�-+�uѫ����9��fx^�n�b�莩<�t�6�9��eyǢ�H���SV(����魏z;p�[X̏��ϒ�/��Ѭ�*i(TDÂ��ar�wj�Ź� p�t�>MՕ���E��0Q�{�2}ե۱�u�z�4$0\�}�l��Z��:.�{1�=�C-3�9z���Z2�rK'D�y�������W�(�
3*��2��~�c�.P�<�*���NUұ	I��@��U���s\{��F�U�r���]_:�gR��ٷ����qKN���X���2�-��:xM������� K���[iԠ� �C)^"2��!��}OS�"�nG�j�u�Y��"7E�����H��9�gSB�f#,���w�bv��mQy�e���%�Y{6T�}�pV(K6+l���p�����ӎ��n٦\ـwi�-�v���5�{����^�ϦL���Y7;�My5��0�����l$S��}s���e��$�z���ȉh0fJ�E��gf��7k��BЦ6��H��Y�����W�t�s�uk�Ј+^��de��n���b!�Y:Q.�5������^ꭥwe��D$,v
��;�7������q(jvCCF���!ԷU�u�I�&���5V�s��̥�ɼ�2�}&M&�چ��w�/d��(� 7���	��լ�eK�R�@��2�%�I0��Xo8u�Ǟv�] }T���(p��0��F.w�ΰҁ@X��j���w[{_�0H'�;��۳�pE�8�!��ƭ̾�:�7gdiN��q;J��6�fV�f�#[1�P�)��x_^��{gaU��GCk���arY�����˒�%��U�`�,�E��c�t-.M��n���4o�:ur���U_U|hf��st���ݜ�R>��^I�k��q�N�U���?�ʢ�_��$��S���Ha��$9ٴ)�#҂�I4+�������ߔ�,���YO
��v:�j�C0(	ZBW(3��2�N�I�(�^N�j�a�D"���(�L�hXWщ*:�&h$�����DF!��t������̊�A·�'�ʢ"+�*+,�����'��'/���E˔�3�r��s��Q>��r�Y�;�>���Q�t�鞈T}�9��q�GJ�"	�N^��y��yXTtٝ8\�Չ*4��ʑP)���)T�+@�I��2��%e=w�ls���*
��ʸT�tz��
(���*�\�L�kE9y��,�"�#�r�Ŝ����.��ےr��Z�|�*��E�P�S"��Qt�C
�9I�W�y#�J"�
����B(����, �QDD�99�ET��\���/V�w~$R�6�&^�e]R�޿i8��A@�.�k���[f�S�t��2�Sǽ
Jn�ȳ�c�$�%pGtLRG'u��7š�/G���oz�=�yO��|�����R;�Р����R<����%��a��"i������uh����r���׊�H���R�u�_8:]=���w1Գ��a��!��Af,J�R�(�H�}�ի
�����r��ǴP��]�5q��<�w�3؄��H6��ϢB�Ɗy7Yk۪8W���!����~5��U���^��lJ�����8�Q�⪱�����1:o�h��������k׫�NNP�����_�_M�Gq\���$;������n���PXy8%Iή�[�T��_�\Q�������\n���z���;��w��{�YT�0��~�=b%�;&VtM����_M���g�ws�Վ2��I����;�C}�м�#����rE�tfu�]�%�`��7#�ާCz�a����$�m�FYy���u���+��;�o�j5^�h�Hh�g���f���'}�w��n��Y2�
c:u)<��:j���d�Y�_'��v�/��7F����n��q�x�+��{�a#xQ�{SF�SAȝo:֮�\]�o�XLl���x���$7{�n=3or;���%�e~�Oo����s�B�4�փ���Zq;��Ϲ�Ot��|E5C6:L�EhC���4s8ɁgGIA�};�_�r���j�=4��f�2�������A�k�o�:"V�آ3�@w?�z��;�{�{�W���`�76�\��.�D=Qw)��-�u���C��Հ�ʆ��l�C��}sʭ[�=�̶ƿ|��s�7�t��������w�8v?!�I�Ǌ�kd����(��������Z�����^�r=�l*�X���AW��{��f<'��l�@��Ooh<=�3����.�]HX��	OPZ1:f{��l�18���9��w]f��/�a=����ck<�w��'W�&� �c�6��>�@���i/%�Ʉ/E���u���AL��(������-��=�N���6sӽЅ�ۼY���H��n�l�Ppt�c��;����)^�������\2t������Pɂ�0�����Yz@U�$��)Q����a[:�,��%��/�lޙ"���I��-7:�^��{Φ�$�y+岤quAs��6�t�2V�EJ�;��!+�����&t�3��Q/�Jfv�ۉaq��ISvC�sfF�:l���,��k��~��X^a�ֱ��F�o�C*ˡ����h���{�揬]�;=ن�E���^�~��\���ë}J�n;�.���e^C�u�`ozk�Z����Z��5�����NlnK��ia>R�jQ[��;�ñG�}=�8Ej>��&�`vA;8��%�ބ79*�L��q�ֵڑ�31�=�=ۚ�m���:�n��ꌲ�����P���؞	�؜H]M���H]=�(�s*g�;��Ooy���O�گE�i]j��SzJk�޹P;�ރ~�0�X��7�P�7�a+|�3�A�;Am9��:D�K�?�@Ō_�N���{�n ��<��c}�v3������u>��S �;��7��ս5�i�t7��<���RW<�BW[���NC����p��p9tuǷx{��9��I�OG{|��)>�_�仯e�e�g�̟;��`��c{-���c�|�!/�������Τ��y��%]$9�#�e�*���܁*Q�{{þ�*�O��H�׻X��|Y�L�a���ή�÷��E���ƟL��#F���ˈm嚗
�|6��Ꙋ�WӞ7��7Yfw@���%��ШL�TPq������_QPA�����{_g#�15��o�}Y�_��"y>����������Ø�˕���5&^+����^�=��{�n/��~���L{:g�<\9�\eh�Ɗ�����:~2�7�揟��W�VL�Uu���g��Q˅|�!K���߱񲽴P<����>�	�UX��`������qb��[��>���ay�A�B�O�+=n��|�|o�4<.L@P���睡�
���}�[~�[�ٺX~���*�ӧm��������/�U��-���_�*��?pY���3¾��W����a��~�irǝ��<��e{��&{Ԛ=��c�����*���.��0���$^�����vn�����-S���M��a7nĮW`�޲�1
1.FP�A�Խ�NE8�����S_�~މ�k>����/~�� �u�+G�0ǏnZǞ���'��(��9��%�IU��R���%_���4NG��ۻ6�} ���%��e�gr�w,;��Y���>�f���8?#/�����]\g�,lq9�}ˏ�t��7 I5��v�ܑL��^X�_�Xu!۩��r4�;)dĜk�Uw�f�*J��V�n��T1~.��7�ܮ�za���:�{ѱ�zx@�~�J f�Dr��,r��,r��MZ����n��Bշ7�}�5z�71��i�[��/oU_�{���mL�o������P�+ù�8�ܦ�U}\�Go��]p}�1�a�@���޸�GW{�j�`�����-�n/�}�L+��7;ܱ.�-'�5+��>��'�#�_ޠ�3#*����.�V����)���o&�Q��ޝ�V����ࠏ�LFe{&��̅��G����tm��\�
����
���0���Dz�
s�J _h��g���y�ó؄�.6��\��8����UdF�z=b�|��1Dݷ«=}�v���lM,aW�bΊ�7���w�V��l^d�c��*�T	O��{Խ�׫�&	�w�^��g67Vlg}Y���ۍӠ�U�2` ��t{]���u��*�X���a���v�P�T�$d�����:�Z�m��-���EO��㝍*w��X�=���#��H���8��R���`�`��f�gw��6I�q��#T�,y�b�S�1��(̸#r�;G�Ӌڒ+�o掎?3��X�*Aήkheǫ��-}fLk���8W��j�����T�K��-��*ʡy0�_�9~��pr�W�}�^w�o�^������8�Վ2��I��Zwgs(o�����;�O��E�񋬽��C�`���
�!���-�����%���΃��ܿ�~�2,��g>��S������K��8��)'�s��4�a�J���h�,�&�O��תl��A�Oǂ�W`^X�Է�f�֞�=���N��amx樎�{�Pr}s��rt�|z��%liFw�o��ݳ)�{&�ϟ�ڋo*��_�p-ސ�����|��~l9\R{޿h�7Gǔ��]{||o'W��j�<��ܹ���)꼥�S����J�:� ���Hk���8�DW5!{�}����k�|���<}�q#���;��;���Ո���/P^���w���Z٧&�Y`���%�!�OU�ϰ�-,�6d{�r�[B�]/�$��d��mP}��ͬ��v���v�f5u�p+��kU6r=@v+Y$u����9>�"H.a��Y�IJ���)�e[���i�r�~���V+i,����̥�g6����z�>S��ۉ�m��w�%��T�ǵe��كÜ�S�2�lߛ�p��=���o�i�2s�=4<|��|�NxP[�d{�ޚ+=0B
XŀX��m��S�{i�����O{����+�j�~�!�bo���Y�`韘n~�̴b�/[P({OoEw�$�3�k����1��aZ��5�m�ʲ��8{|&ݬ����_����d{X5ތ{��us�l:����vK��>�;�����N~g�{�<�M���LWa�K݆�TՆ�;�e]���8]���K�t{xZ����Q;c2KN���l�`�ؾ��l1׷���hE���6���ꌲ�j HC$�6�x:�:���p��v
��V{������5ꀿ{�����M�J����Cd ���G**�O~�I�@9)	P/�Ŀ1�faܬy�5�%(�k�[;�JHM�gR{Pb���ĤxwB��N��e�lfa��6�}�7[�5TaW�v��ky`�ʸ#8p��*�ف[�J��(��{�*
��i��%�d�t�fL�m�����)Z�&u���Q+p�������֛鰩�wh-���sAtw�W�|��V�k��g�̟=�x�k�!�����=�}�>}�%_�f�G�r,��.8�����o��_�hݴ6�U�42/�]�7���z��t<�W���A��b+j�{�a�;�3�4w�֏Gg�S@���k���{�h��F�|(�+)����'�X�`k������H+|�h=��v�5��]e�%w�
�,�j����x���'*��u�X��4w�|���R��r�/r�[����Aw���x���S�$.�u���ηƦY����tg0��eY��u3dc�?��׊�\��xL��'c{B��������,؇՜O~�{�zU��rсz��rfkʬ���=l.�y�M�}�Y�r��o��ھ�#1�mC~����z��khN���X~��AU�N"6 ��md/KSH�G�~���O�$B���G�c���w��u��*	,oi�u_R�KmC(��z�rn�v��{g?�4��՝A��.6e$�z6ֹ7��[zj�Cs�#�SЪZ�Xk3f�g; �{#zkkLwOv�˳�t	�z!�T�7�:u.�Wm>F�UYo��N.��	�_������(�����jǩ��a��!��������DJ���*����Z�wos��U�_�2O��a�/l�}�ڸ�}�t�9+��ችX��6�ؕ��m����{��= �\�S��?�s�$�O������\��r�v�YŴ�q�A�]}�eV�}�T��"L[���X����C�ë����7������`���;�mw���=���W\E�i�>��1�0N�;��j�ewy����RR����Ê=00!8k�h�w7;��#wP����Lw�c�-�֕e�w���8��R�`X#+=�K��g��U��vXި7��o}�d&�N����[�*��Ʌ���=q�o�gv���.�r��u+��ТXߺ����/]�T���͇�.f����7~M��C���.��{��X!J�?pQ��f�s!��%3��d��eR�*s��CM5B	���LV�)�W�cN���W �U���W��m���e���C��us�}g\����ͩ	ɭNGxmM�3��;�Z�����ۜ��]B_i�;���,�{Ҥ�(���P<BC%���<}@�h��zwxM���a�_ۣs��)�}�ü/�j«p[
f�P�Z����np͍P��
cћY�w�b��m�{=���ɺ��'1D^�B;���M����̆1I������׾�������A���ܴ/<de�3o��ˡ��	`n=�K~��u�NE�A����kx��x��T�t������ܤ�#��ۡ�eV�O�%Iή�M_nAk;Ϯg+�퓪;���m�Ʃؗ�v��4V}y��R�j����{^՜K`�"W�,�Ϸ��`�//�v����V�nB��Ñ1�^{���b�Bü���}���BoyV�6����h	$���\�T(A�~��Pl�!g�N�ϬW ��i�\��;i�VG����>�0�y�{�GgR�z�k�}7�c������nRY�y���hR�r��sl v+y�4s2�V]g�e��E��^骐c8��*al��N�WD_�wL!k�1�褽����ܕ��7�]Nս8j:V$�`��T�.ۓ���xOTsFwj6�ǃy��>;��*s�cgWP��-�j����7q�=0]��۔�0źeel:v�d�\��ΐ�L/mK�ˢ��!֑�4���1^Ψ���R�9df�*��E0��J��|�v�<Q>{�O��t�����Nv�U
c4!�%^�yY�j�$Vv�\P��f0ٕ��E��Ou��Ǡ�Z54E���B����\�e��tT�3';d������c+�
�W��>��Ba����5K�.�j�֓�jWk�;^Y��$&�5���4)����ͬ5N.�W;:KZ�}�����v��<�܆��.�)����<�L"E:qpG�WG`�̈́��.�"��5o6J�/E뗰�M.��osD*`�{Z�d4o���L�§׭���s�����q_^]:D�EHry�G�r���]�ۧ.��Ga�`�:J�̗P�L�wf�ҹ��x�b��Q�|���l��	����s��M�0k|�x��x�f�f�v��̍7������\ ���4%���T��3H͛bZ�75rЂ��[��0�:L�Tۤ�Uuٝ8ǿiǩ[�"����s�܇�ʷ��(d����e>�p�,�uh�\Ռ�����!ڝup��ش[���D�w׿c�獮���A�Z�|�q]�cw��`��u�B�B��������M�]9����db�Z�sT�goyw��<@�W�������v3��$z��{7f7͝�ŵr�M�Q�9j��u�m�:�v�o��ʾ��'��J�4��` �2r�\8B��ܮѼWDk��=��VOC���;ʉi�Or�8�c5�WDo ��.u-�b,�3�-4���9��ܻӶ:���&z��V�T��KV������	��˺�kk&s0�����5ƹf��z%�M�"�]��ʈ��_����vs� LSE)YN�Dzm�|��F��|�Y��涬Ms/G���f�
r_AP���n��C�V�L���H�W^^�r�#Y,���.fW�e�V47��l�h�+����/:�wӬ�;�-b��v�P��Q��I]��ݩ&���]K���r}U����v�+�C�{�w
7LM���C��N�M��xZ�/.���Qh��[�`��|�z��=��vH��e��a�$���i�X�8(��{�jM�GL�����`5&���5w�Z&l��ؔ��N�� �C/o��Z�X��SZb�T�̝ۡ-ݼ]C��V����v�0\*�c�*����$^E&�k��y���ꦎͩń���L+�9:o��
YEѳB�&�k�*rJ�c��bRX:b!���wM�y�����X*��z-Κ�_Ƿ����:�-�&�k�ճҞ��'9�ꩶݶ�*�eAК *��A�F�_�r!�л̋��'�UVw��6�y%,���?���~����"�E*�PTWT�"�ws�+Xzܜ�.^n�]Q�1k��\�|||||�0��	'D*�NG�q��A�%u���
s!\�C��%=�=�=�/D=�W�&�Ukz�YͨV�
*\��M�	oD�2�nr7���N�t���3�����į:(�
�G2y$z��F[4F���^w*C�)��ȉ��1:�������2I9k1E�b�^���5Z�I�S�QQuK��Mɮ��2;�'�TO2������[�J�))QZ�d]�%.�W"�qD�>�8��\��]Ī-Ny>g�"��L9��9!�'�[���PUG"�"��s�V��E*]�u�B�ݚ�v�V�d�t1�z� �ʺxY!���;��xU�z8�J�jF����YBr*.�r�T滱���Ră�p�[-H���E���]�}�ɗ^��茎k��t��E���5�7z�֯�����9��lp����o90�}WWR�M[�I����Y���/(�0݃zOM�����C��F?������T�z�j�������:`=��{�?YF�����\*�ln��ߓ���h���g���Z�v�!�R j���<�rSF<�f�n!����g�Ou�)c�\��m+�z�v<v����Wm#��!:#s���P��<��~����n�Mu���νr�����Ev���X� j}��Uz#W����Brgq\���Q���X�ԂC��蛓��^��u[�쓻-�ኆ؇#��%���V6���p��bt�d&�b���������=�g�-�͞��1a����{;�p���X*�N�Y�f{�&�sj���OߚF$_��͕[PF����Ŋ���+��Z�-���~���}��¿~��>\���9/y��ў��*˭��>�n��:-E����s�<����~>��W��ީ��?h����+�����'��ў8�I�W�E\�BK?=T4�X^>:���T!��Q��uLk�5Yr�N�yV-W,���(P9ԧO�!����Z�7��Rub���t�ri��=�Nv��\�S�:�(G����b[,5�{���d�Q��n"��BgU����d��.�ڟG�kE*$RP���;�xn^	o�[��+%����r��6��^�ps�:���(�d{2<��VMZ>�����$,e�Zp;І�%�[P��팟H�F�+�U+HG�}k���M;����e��>��Iln�ﳂfU��~~S��G��3��K�܏������{_.ű��,0�H(=�O�1ζh�Quw���s>�bvWo��o��J�<NR�z����P�@�0�Q��ϩdF���x=5�gS��+��տg>6�����>��a��:�ٽQ���&��$g���v�T窻Ǖ-)e�7��4�pV35ݱJ��37��_�7>��361��S����X�$kG����e'�_��`/E]���h'�<9��;�y��v��u�����a�o����r:ߤ��t�;y�1]�}\o�ի�;M�asex=�C��`���j̼C�lM�ߧ�xl��;P�"�ⰵ��]�}��?e�������17|�gR���j+�z!�ީ����Ը��2��5#)���M�.(;e�dr����W3��嵶��F��K����Ʒa��ɚ��1Zu	݅����1�;qW\Z�y��;�~����ɜ��AHŊhj�Ö��-��ʯL�����0�����UW��[���[��^��1���؄�yp��
�w��wӅA:=7\��G�����p�^�F$��N��퉓���wϛ��m�>�;vϫèG��	m`�G��ߖ<+f/����������ONP�s�;�$s��~���w}�j�^s���Gϻ2����0�@�+(I���S]	�+̛7>�y{]i�p�K�U��V�v��ê˫�?H].P�[���(w�Ge�;ݑ9��������|��a�n�r���:�au���CÎ}/����ɯ���o/3*,�f�����z���M.��|i�|���P���^���x\;O�p<�t�P�Q�P�8i�T����}Mͅ��`����v��mN`{�j���4}��Q�?hkh;����Y]�n�=5Ԕ�Ts,F1�+630(���L���ފY-�ʻ��X�;5���W�H;�ӳM�V�#�)\�q�Y��l �W�qU�i�xbӗlf�����b�vf��4%�}3guv����g]�Ee�&\U�{��\)Ԗ�7�Lg:�W""eg*��nJ������3.���t�ߝ���3�|�-B�,%p`��U�����ވ��6��ا�Ae��c}끽 ��Ʊ�5������;���z_JLk�qK��仩�M*j�*��}�Ac{h��+
���h]��v��~w�*[�f�5��<�V!�e���;]���a�&+2Oh]���g�\!�~����̃��n����c�T�Q�ILOx__�f�;K,pW(e���||�`�s#Ft�x�mg���Ӟ�&��B�m��*�������M?.��@^��+ ��C��o��md��w���њ�����j��w�/.�,Y�������}�����k&�]N�����dǹ>���u!�Ϲk��0�z+�o&���0����fIY��W��g
�|ڗ����Sn��[�9�v��2�z
�dpo��ps�������q͌F��W�8�a�xU��۴	D����L����P]I|�!u<���C �ˬ�H���f+3�\�@b{�b=���Tx܎f���S�5�����u7�)�d����0��f���c���r��h�u��E��u���������6D�n��'���g��3�W�2��I�ӻs,����3�S�Bkp���$>���(<���{ʷ������6�fa��F�X){=��*���o���]��C?�O ��@Zq#��sL���Wb�|s՞���v�/lڱ�Ǩv�T8فl1�<��5-�[� �N���|�Y�p�.���3��*�ּ	�A�<Ԑ�=�3�@{7���!������X��}5s�O��r��ɣV�zlR�X�d;~�X�ې��}��W(ݯ-@ȈlKiU%c��n�K�\��J��쫡��g��l{(�b���>���A3 n����Z���5|��{'�]��b�c�U�q�����#�󂂃�� ��P��uGv&��>�p庪H�5@�˱��_���载-�ю���D�a\���L�W��y���K|��
2oǨs
�7��.�kl�>�r����kubj��
1R��7�u�=Ekh�I������.��Ӟ�9z�����ؤt[z/�E�݌�M��ޢ.u%Y/x�)I���gs$��|��jN�6���՞���.ѝ4]���L��3�;��ɜڑ9�y%��k;;�7����l1?>� w��ٳ�=0C
g�yPמ�W�� �������g*���ޑ���^�ݵ�(4�H�[�Ef�1�D��vT��e�N5o��M��}4��ΟR����0�[[�kb��ۡ�e���V�fn�;~��=�M�O���޷������{|�v��Kq��.�x����yDǎϽ�����eYUb>��6%�_�M�{��a������}:����fo;���i����c����Z��^A�B!�.�����p��Օ}�R1��~�oV�ow ��_'j�N�e�CT�2�bG���b�m
��ZP���}��WRoË�cM$�����{�~0�̪��̠�Ya�{</�]�7:1w������V����q��9���gؽC����+эb9`����e������*����)��=�� �^����aY�w�yKV>��Qw.�1�Q�~.��3;J��n5E��3j�
/��t�̼�H=��؛et�=�1�o��&ι�*j�M\;Zr�_&>���0�5���I���V���7�s�rI�:r��W��ݘo5fl��}W�n?B����UH�@�5�����PC�j���e,�����I5��%iF�Ew���������{���l�7�6�Ow�|���'޻�]^�L�1{{>p��s����.���X���@ߣ�I�5��V���܌�{�f�uo%a��`l.o��}쮱
z`��#���d��=��7����Z'��U���p�Ŋ���C�j�\V�]P�zco��'ޣN�賯��D �EsR�X���S��'ypߛBB�3�?c���4��v"��K"�|q��x[�Y�g�Y뱾^�������X�½�Ȓ�w'1���B��+��;+�Pp",7 �e�֐�����_�rs(;.�Wiyz�GN��Oǯ�]�d��^Q���0J�r�p��Fw���'{Vɬ�Өp�w!C޽��R�Z�u�M��]?9C"L�b"6O�����.���_�����uؘ$
��M�Ż��r�斎f1Pk7q8;]�x�Yβ�I��c5Utn�����:�T����d��<��V�����zX�7����{��'c��-R֓�Ϟ�}:�]�a"g*�V���IC�V�T�oEn�����������7�]w�7X�e�~�F{s<��P��\R
����)ݖ�qm>�z�=[�Վ��<�E^��w	���k= ��6������'��7k���-z�Տ*�CjY�x�M\�^��0(���Wǃ�MP^�����>1��I�#�����Ϯ��^]�;�遤qc�-W����E^��f��`���;�[��3����j�u�_R���ޘ`7Ӿ�|�����ot�N\��j��~�z�a.�yM*j�PW�@�
=�"�{��USPv9��{������;({5��ɵbMa�����p��+
0�&M̰���m�j�7�A^єC��X��c0b��ʐ�Q�A)�9[}x+�H���מ�9cڇ��, �ъ@2�_�<���r�<���~�<�?�K�H��`�}2e��Z9j<�1�X�ww4ÙQ�j�K�)��6g(����Eun�kj���ϋmY��
�Mь���Yp`�8T�K�I��{�����t<��b�x�l�w@�a�T�tq^oF�qu5wnf��9#�v+�o���Λ�����:ᚢwEΚ*�t�c��|�-��G��ۧ<�R�_�=�ި����[X��q�6�7��0%?1�'���Q�=8K���ow�3��C�r������_[�A>ȯ���*ʭ�,^�S1oӗ_@���\�[�����X/�S�T��h0���P��R��vP{�B�ʃ5`A��T+�z�w�$��/:^���g����Ň_j�֒n�����&�ﰙ�3Q~�9(f�;y!�W�X�}�vB���M��]U���E��N�c��.��{����FYT6�2}��:Ñi�e)�U��D���}3[]���ot��C�:�Fȁl1B8?T��O���L7	���/�~v�#�i16v�z���������3�@�c������n���Vz�dA��5��ۏ�Z�<�t,y���_��TE*}�]�j��oNo�W�o;���AAJ�-ei�0T�xpX���9v��_m�������d���lטV�cm��
��2�R'�g9.�[���/4����|e
�O��x�xy�L�{t��TWCJu������e1G��PK��W����L�}+�w����}T��OR�{�o7����0�Fmo�nZ�(���(���:�	����S��R���4��}����@���yײ�<�¹/+u,�͜Y�$z�l�������!����mg5�9{1Wf�Ƒx���1���p^�{�h�C�AL����b����='���x�[z)�<]�{���i6(6��L��Cf�W�`�/�D(�|;ڻ=��޲������߯-	��\�#�d[�E`�d�0{��\X9���F��w�e�ѝ>��6+����cW�kc�N��ޯ5Y�Mv���c=���y?`�?z}�X�wꝡ���l>�ܯm��S�o0x����j��=y2�����Y�  �E���hWݚ���K	��:��"*�\����\"��ޞr��ne}��yHN�Zv�8{�|�ʪ!Wx�9���]~��K���BoZ���^����3P��G���x��֭bKr�n����/���Ui��Y��o{�mJ��ހ]Ы�:X3�����'n݋wX8�� l�ʽ�gCK����kVd��i�\�	݃f�ݚ�0fнf�H�o5���)�����jf���YKt���ZDӔ��meZFc�"�j�����] ��r-P�lkte\��Fi
V>�A:�G�Yu��r>�w��1�p7k�YcW*Q�I��oZl9���E�E��y
�̙v,5Ek˜EU����˃���w��T�7��������6�z'�y�/y�De�������>����M(<2o׬!~�v�I�#Vh�^\V�^�����h���Ȳt����Kz�X��65�]�9Z�vʌ��acE��34�Yy��&��1NF��;xFY����[�f�&�OfX�Z�oNf�T-�"�1��K;2#�"�8�+J�;�ye��F��9�M�3��6&D4�xgb|7�+fJ
*�̻�+(�6C��bi�}_b�.��a����FӶ����w����N�nꭠ̣N�9�xZ�����st�Q�I��Y%5Ox�y�p���ΰ$����r�!�2&�V�ݶM�v�4�:��v��q������EJFo���3p�Y}Bgg�Yy3��w�\����{�U����5Z���e1[�[X���X���kY8�V[��!�;� �oc����(�\j�Ԙw���kL���9;e7�p�}��t�-˝��S/��B:�j�h�`o��d�Cp��u�پ=���5>�[�q��v1� cR��-T�^]��($��'
܌);�t���Ś5n�<ʝP!t:SZ^��&5�-ו�*����i��j�e�훭�V7��9����̃�
�A�/����8�N��ʆ�j��Dƪ>��M��{S�2Б����ɂ��v�U��䧧��b�^�Y.������zk{�`�|��j�\�x�1sY=b�s���N
�x��^�W�V�Z��r�(
Pk7h���Yӭ;����`�P�M(T7PT�"Ȫ
��n ��0vc��-�����9���}�S{�6��X�I3�{�,6��|e��6I|]6`��w0U���l���S
����,)Y�k`�g+u^͙����2c�����a�ff:�����:���5ֱFݼ<����n�����T�;�uk�T}A���ϳv��Y���'�*Vt��Qb�:��=Rs_-�����]�4WL�QS��PJر݊�of#˩�sJٷ�qV��1B�����܊�vF�h=��!���'����n2�F�0�d�º�J=qR��Cq`�n���/� ��$AWN�X���kt���{2̨�.���&�]+�|"W}c.�,3u�<[]}��J�S݆/��}<{7��K�֝��v�'FoY{�˥�S��A#@���?�K��i&e�}׏r�C�\eV�b��8�	�=Dq�?������pԪ�DE�3V��NW��һ޷&}H��R�ʯ�����|||}���~IUy��<����/S�U&�.DGΜ3������r��y���QU�DkY'H**�QJ�"�ȮG+ͅ*��ΐo[��8_2�ҹ%YW	X�.�9��ZAsZp��RQ��r"�һ#ҍ��<��s%��k�ܪ�*���rQy��c�Yn���TEUQO1E���D�r��2>�ܜ��J��es[�\��� �P)�G"""���P����s$�UE�(�
� �%�����)���ҹy!TwZ:�^aTQ�gY��
�����ET�ӗ"�K��E�����V�S�G+�UNI�+�����!�E^K".T��$ ����K�d+��/�<�^~��.���1�YNs��ݞ�Zf��z��G�v�e@���s:����v1�7��y�*S�����)��WXK�����:�vYt5$!�[�8��T�̽��y̟`����r�����/��ů���T#�24`���Z�e��WA8}�sNp�A�c��:v?�݌޶�R��>ge������
�{Ԅ�g����W��7�|��������ί��͹Oq��NR�q��O��ӁPƘ��4{����T6�Y�J���n�2O�o�}3���g��zUy���� ��7��RBj���P���&MvP��аqT����OΓ|�]�J�]C}�#���~�I�5�/�E�j������flC�*��-6;XnS�}B}�GE4 ���d�P�W��ޱ"��M4�w�Y�S¾�����D��ңo=߽K����ޚ��gN��9��
{���Y��}#=�M�h/��n�g9_b����u�m5�/'2�����#���$�,=�Kmb}�Qyt�u->Hym�ۂ��]�oЎlAvom���v�9c��w	�"emٛ��@�b�:yWE��@ҷwF��j����O'.���q�ޒn@���-l����.�)%�L<�Ҏ�R����l���h�g�ũ5��Ug�|�C�µ�I9PP���t̊�w���^x�Cs��~��e�����7?̾~z��IώuxWs�T�5�/ݻ���ۃ���B�����u๢��$`�?���5g�R��\�{�s3�����J����&�l�O�;b{=�F���]�4�Oɿ�������m�1��H���iA|�m��^��}�����f`S��ﻵwU��=M༒�͔d!Z�����\��6�f\�I��>Q#�goA���,�h�S�Hu}�T�8߯��]L�Y��,F�:�v�j������k����@�}_u5K�]}��s[�VwcR��ö�_l�;}�e�˻ˣ���P'�="��?H:��N�c�>�̪9=��lr�'w�弲�r�cr���K/h��!xo0A���<��V����K5�z����j����ns)��p��j��U�Ӟ�͹n �_v�����E��r,q��^�{�J�ˤ�� �S.�R�y6��rĭ<MȓӴk������o�C��D�&�v_s�M����L�h�il�	W��	�2����A�y��֫p�{V�Z]����_+� w����ūʁ��5f��
�rGt䅕�|��JVX]9_oN��X����I�ݶ�X�;s�M�\#�
<9ٟgzB{�H�|��T��;�u���3���(�眻���[��=��x|L`b�ъ~2�_�<�}�:F{�3>N"��aR�b���Te܅��ˡh�kD������Y�n��z��ƬT�r#�{Ք��F��P�v��;��!K��fۡ�fv`��7�]8ߕ��G�jY�هE�x�򽜮��-a��⠟dP�[��*��\s������k<�@xW��q�������Sn�5N��W�s�2����Ug4���o�ó�:�Sb�Y�V%�8��j��M���mT)�{깫_fz�r��ߨ�=Q-�B��[��d��$�7-�n��x�~��k��4]�M�r��}f���e��r���ְ��[�R�З�z�$��Vދ�Ǫc}�&�7C!&s����Ō�5���=�z�;�����k0���
7��z��i�to:�i�W*#��o$CF���	�z��N�j����p�i���%��J'�g���#׾��J�����{:����`��-=��� ��Hy�QDN������Q��W�Z����}�{��nuQ�]0���3qx�6��ק�\�����Xw�}�ԭ{���z���5�#��cd@�ێ#�k���f�`Z�[��@����v�g<�94j߸��б�XY��/_z�_v�h�$�r������]�>��ڭV�:�Ս���J��ǣ��=A�r��Q�Z��s��z�{���)��}�cs7:�>�t�Y�r�<,�@�G�В�$N�=�_t�u��z�:�5'qP���Gxu�tFD�uJ��r�VgV���C�_%=KF��A�L�t��x��1�����0�o����ϭS�PS�,����b�͇/��x[��i���!���/������o;p^�Y���Bs��Z~a�|��}��*��|/_���Y�����h��]jkr��z��;���� $�J]ne��d��F�j�P��H�:Wqԭ[�si��s$}wn_e,�R_w���O�M���\�[���*���Ϲ�r.����d?��k�0��f����+GLܐ��ӲD�(:�Jг7S��I��?�o�u�n������W݌urƓ^�bf%ڟOed��ˌ�<'��>�6N���Z�zߤﻘ{Ɇ���]�H����wmb�FU�q���VU�_Xa�}by��;5�K��'ݍq	w��ޭ9�9���v��`Kꥹ��ׅм�!B�KLP�ZTh� ؾ
߳�����؎yu �J���Iڿ�N㯮��FB�Ix0H�Y��M��Y�w��<=__�9Ď�m��_+�M$���U�{��9���g�U�ob9X��9��@w��݌�׭�J�4��8dO��}W\5�w}���ϟ߻㌌��cUmS�����U�zh_6�[�z�"���6s�����^hΘ�����_*ڭ}*������8�޺��G��4�F�yϷT�'!�Pۀ~��<3W��{��wb��jC�^��IG��c}�7��ꨝ�����ӺT/%=���U~r��ީ1`�3��{���7r�n�۔�k\FX��ܩi�-l�����'KGkT��vvc�n#m��b3�̨��@<�΄�ɿ���q37����Fs��j2�IqZf�k=��4%�e}ܶ���Gw���  ��K���y�A�c�����-��(��a������c�C����<R2i����5;�0��C���%�[�o���<+�j�\V�Y�y;G��42�31�Z��G�LXg�;�S�X֏j���rhP�Ͻ;'�.�<M������R��+�h�����cX*��c|�@=l,�h�{ж!q��xV]������+>ׅ�T
�vd��քw��;Ã�'�EU���=]H-�cqkߥ�}�]y��^PXy���}2����3|�yd^7��7�_�#�x�&��RS��vz��JQ<%�>�X$��n���?|9�\��P�b~�}_iM��m�\��c�,9��[l����DuWOw!7�ev9���W�1��w�	�T+�M!��`GS��W�����W��������[�',qhE$��y�`�6���3s�zx��<��
;+Ƚ�Ra֍v��?�D�K@�7��[̼/M�c�Ŷ�l�8����8l�e��;0.<�h��i��
T|�8r�\z��oN�"�#V⬺;GjG��t�^��%r�W�|��j.˯���= ���!�ک�=���}�˞'U��g3��/�o{R�*���{����b�����쮽�qf.A�wڡw��t���_Z�����.�N`w���0�^�+�#��M׹�>���>����Wܹ��R���K/z���j�z�2�Fo�˫�Z�6�"T
��KU��[��~��k���o)�MX�W
�>��p6�$P�n�ߴ8b�d�7p�0{����f���zv��o�7�~ʉ���f�q�~����:  ���3�������_.R��U��T8Q��-��y;�z��}�j��.�`�1H2�_�<�w}1F1!�j�|���7L`���j��ءϢV�����������J0��+y_Gf)�%��W=����&�X��
��fۡ�I�+�#�=�p������M���Y���
�-FN֬��`��[�J�
���T7����٧.�������B����e��V�l�,�s����0�V��Ж�{#��9Ԏ��s+��<ͭy�w�;TvJ��o�,,�&�8�wvwcP�g�l{�Xz����-aӾi�E��VU@��9g��X�<}���|<~�c�v���-��g�+Xy�6�e�ğ��^�>��ĥ�o����U����_�Kb�<���8��Ƕm�=�:��NEw_-�C���<��L�e��M\$s�ǁo;!	������P�{Q��{��޽;���8Ϋk������e��B%���o�}���0�{�*���C{"Gmry��yƝ���ΨQ�a��.ks{�j#���_��xL�ƶ��%�tZzhoZׁ4��=A�2�7��-���]Pqb�����6�?ze;��{���G���[��� ����\VL��=W�j�c6`s��mV���Խ���i]L�%
�~��Bb��f�R]q9�/�*-���c��F��}�����Z��׹B��� �/1��ˈ��
�P��Z;�	�oz⊯���'E�e���Wk�ШR�2�1��9s �M���]Qú�<2�o7��9��OhL49���e����	��+��.��b�6��SQf��k�}B�<�wc�]��i���WJ�Î��X�W�q#�u����:)��<����rW���������ӛ���y�v!�+	�|��1WX�4�;�5�.t��D�;O���q�k�ܯtl�ch^-����2x[���׳]o�g=b�`xg��YK�q���] �I�W��-7��׷����i�muލ���F�v�"+���&����c�B}&�]]�s��b����	�]�Hh[��d���ƕy���:�U`1�  ��9��)�w��N�suݏyX�̧=a�Dvo����t�on5ٞVUXa�X�~�����B��ח���-'�HjЄ�r(y�ܩ�mӱ/��nek�����!f�${n�4�^{ܫ����<��x-�A\��6�����]��ہBz�n	�=	��7��`�	������'���q|�i�_%��w��}`ꌳ�q�0*M>�U����b)h��P),�,�KU�X��[�s.T^�K�c!L_J�}{�/�+(M�8ɾݰΠ,�L˖�sv5��륄\��0�&b�ރ�h"��J���;K�;�j�#�9� �*l��5��rʴh��&��
Ǖ�cd
IC��)j����~d�]�U�c2/[sa+|�n��{�j�z�bvj�w�Jk}�>sx��F/���~y���x͋�5��v��c̷Vַ��6=�},���^��� 1����[U��R�h觞�QTsbd��	�n!�n��Hn��ø��9wC���}!l��$&���w�'3�Nn�k����V��O��Z]�Wv��6��t���WQ�דV#ތс]���E�;���9N�&�F�\arex=�[�!�?/�O���x���V��v�sEa�ц����2�o�wX�h���[�Wd�C"��M����_z��Lpf��Ο��@l�5�� g�	�\�	P���	䷻:R�C�8�����h����Ƴʬ��������{��@��9����[��_�7+��hX�A)��wZ����t��9R�sUEi�Q}ϰ�>tQg��jT��HP@ 8� El ���"� ��;m�E����""�~{�x=��D1�A 1�4y�1ñ�p&�l�� m�Cm�m�A  A��n�#��1�m��U�U�U�U�U�U�U�U�U�[�Gm�A6�d�� ��  @���������  !�ڱ��m�2�
�����*�*�
�*�*��P*����*���
���*�*�����-�������L`��@�OlE!EH�ףL�v��g[�_��>_�����>߫��ʔ�+�Y��N����r��PTV�q������*
��<QQ_������H�r����`�*+�vN�C�nP"n��=������Q���s�(�QDE .�  ��&0�DE@"� M� L8��� D�
�"*� *�D�*�"�@�(�B
�Z��%����?�"�+ 
H���Τ�{�p��í���� ����lS�r�B�[?���~�0��X��UE}G���_ �ñna�EExE|��@�:���*�
���8�"��4y�B���q�
:я���p�o��c�b��uPTWr���s_�>�PTWR��%j:��?�<ξ���+����L+�t
*����Нj����k��V@�>�PP�G@�N��[Q��q�`c������Y!a��G`���vnuv�PTW�ٹF��Ei?��U߇F����e5���� .��� ?�s2}p$���}J_FM�l�5���f����mH���UM5��҂���#M%-��4���T�m��Fت��*�@�KfƬ`��06��*�ծ�ۍ����r�w[��l��ݶ,���ݤ�Fl��}4+������e�:ݭh��;i�5�A�l���f��6�M-a[f�nd[=�
��ݻZM�[k+Z��vVU��sn�[�m��Z�h+��֤�6�V��۝T�����Y��5�m�fM��l.�"�Y�N1��i&�;;���l�v�Q�Z�f�   ^/�|�w���$g���j�nնsv��A^�u��-���aw���O]�g��{�M[m��[����A�����{n�N�^��ݞԝt��F����TvÙ��e[/�  �r}��H�aFC�W�x�K�6�I[�������F�t7cZn}=���66�*�K��������íLVm��nԧz{s(K�sT������
i���]ڻR�aJ�yΚ�����V�ͭU������[�y�w	�o�   ����:�wn���ީ����M�vm���{�[ݦ�u�uݥ��%(�A���+�{v�^t���p�Z�ދ<�{gWc��[�ז�v�3ܜ�w�T+���Q��kgpm�F��n��  ���b���ފ�=�5����k�T��U�f�z�y^�U{ǯM빶wj�{�փ�gs��-� ��z�קMWM��c]z�*\�w�����@B�K-0���uUZ�ݜi��   s�kֺ}�ܭV�u�颩.��m Ӹ�]�4�-<s� .S
T�kTz�^l��f�%mK1$��h�fͱ�|   ��(�De� ��S}�h=z�*�U�5��5�q� �&�\  ��ᦊ�yP�P:ow���A��fSL�lZ����fvݭ��  ^��v�R�UOvyyGZ��]�X�=R�^��������Th�;�v2�Y=������@�� ��VZ2��wmӻJWZauw�  �� ��r�� ��ڀi` ��{׀ �����B�Л����[8 hX=���\Vֲڨ�WU����J��  �� ��w�hР�{p Oz]p h,  3.������  {e@  f�ptI� An.�v�黶�f�j�Rm�CV�   ]��( >nӀ4 ��  Y� h �z�  ^�� �myp� �  ��� E{]��� /�"��JT� S�0��� �a ���ʪD   E?� �����&�4  $�T	�I  O���4���o��ٯ��M�����n����,�������}���<=�<=�v�E����oa��6?��1��pc`����6�6���ǯ�����Oy������q�+�M�=��AdC��Z�Y����Rl���R]X��5� ˂7 t1�G�i)� �O6���l;Ӫ���23����bYB62;�,� 3�-��w�C��A�vɓhe@�"�����%
�/�*�AKT�a-���-����	�Xt��9����t�:�æ��*�������}���J�JU.���m\�l�J�����Yr�\N����6v�)$�dN�'�B�����m����<}�T�Y�PCL�ҽ�Q�IS���EVV�
A娊EZR�˼ң���˟Y��4�[�i��1�˒�����D��kY��)����SeI���XX�fXh�Ak^�5��*��s^���/,B�;9�tL2�/A������L���F%�-��>v��%���t�B�0.�s3w�z���ab�����M�T,gƃ�J�-;���{�6d/D(D��cU�����l*��\�el�������А.Z�W&ѐ�K����zR�[�f+P*o�ɹ�����/)*� ��6T���L����Հfw-�9��tI�&48�������7,6���{�#@��
�UƶS%Qz�.�\�mVR�qK���	�0�i��X���:6��@�����t P��5f�J]KD��eK�Gb�)A;Z��3�W��"qc�G�/���8��˽��hM"�h7�F�I��/*Ƈ���.�r��4�W�"I��	
�"�+H��A"�����j��9pڛnk���3%�0ޒ](��9s.'0z&�S�c���9lnPZ�D,����;�����d�/1!B�Ga�C��8[r�	��`�Ʈ�-�[Mf�z� ���ŭf7���B�-<l��9�$���}e�y��+0sa7t-°�>�yͳ�N��BF3�{
�GJ������ m\i�IPŀ��g����\�ۚFv��.���h�W�r�`+��v�;�N����c8ygN��I��7�1�z�h�I��6Hr-������'�Y�9�B�R��M�����ڏ�J*��fcO66m��۷/j�P��$qe�ܴD�в�ڸ�ۈ�{x�������>Vم��k	5��)a
jk�,f+_#Cb���X��֜��X�R��P�en�;�Ʋ2�R�oK.P�d�iVm�y�l��lڶбv�5)�)�dÔ�)QDލ)[�ٗ�H�ܖ�4J��mbc
0�Ӷ�J&Xm�Ǥ^^巉I((�Œb�5Pܔ/41W@VI�6�(Ҹpm�5���=O&e�vqM��ƭN�ɩ�颦f-�ʕ)�X'���
�®�Cl���H��ڂ��7h������P�M�٘E�I�U.�իV0�cP̛�������MZ�l�-�՚V�jۂ\ߎ�%cb�"F�ŀAM�CFe�7!�$��Ӱ)t�-�:�{P�����7[�ػ�0�6��ˬ��ra7�%
}c4Y��o�ns$�2c���|���r%��H�0-e�.Yj�kwI��"�[b�&w�S����^����I�a�l�TP����;�k%	��T��/�nfMWr�Q!��uB��Ŋ�t5cn�����& IlJ��v%˺+`�����X�[@5�v��껺9b�����E�{��ӣW����1�.�L��p����j�gE��B�7���r��#R:����sYy�F���-T�X"p;�tҰn�{D|&Ѹ̔Ƒ�Z�L*�x!-�3D�����
)���=Uq�n-W��h+̷���d`�p�2�I�K������b��M����`ǽӴ,�Wi���k�
͢�F.(���G]�Ҥ$?ӕ�je�"�$A��\V���8�͊ީaP�>�յ������<�2ȸ�Kua���5��p��m��S1�F!��sĈ�OO7f�Z%�)J�Ct%^�Œ�BǙ���i�S&]IjmI�(ljD Y�mD��	�Vn��L�ZƙR�I��T!�X�^Ɗ+�p�:�pK���1����X�m;4�2�v�5��٬,E`���h�hԌ��Q���H���V�`{H�bc7�	�Ѷ�������H�ď�0�7n�3Kwl�a��"�7*Q�����D2�Y�C�\xi�l�yu�d�!��	eDV[0�� j�%
�B��yte'�v�ܞ��.����y������ �J���V�8��0���t�`L�%��f�a���!Wn�h��J�C!�� ���L�F��e�%�׉�7	h��&��.�q��M%Ѹ4�Lq,	eM�,��hµl�3C����	��f���F�^N��k��CYY��͇aث2�JA8�+k�d�vNKSk2�VLץ�Ś�X1�Q�$���.��*�-��os3�+jVa�P��lޤ��.��-�4#A,Ƀt�+I���ӹ���]�,��Q��pb�啀�30�Q.�hٙ�!Cja�)�Tqa�3�k\&t�	����,[Ŏ	oɴ)�Ӕ�4�IeBw&Vb���J�cR��|k�KnȼV��Zl�4Y���?µ�01��z݇����]�֞�7wEin��X��2naA�`3H�[���K|��&N�DBp����x��XM6�n�o��K>ImzD��f��ˣ��9	ғ6fI��YUp�w�X{3*��@������ɵ�2�I�����P���n��M�3iCG3B[fԼ�×lMvձ�l���KEaP[���ۂʺY�Z�f��r'չ�S��ʬѯ�oF �#��*�EP(�$��Y /���cx���K
ot�Tƙ��۰���Cbv�ۺÔ��]f�t\QTN�"6soq�Ӗ�0�F��
��!1�^�SE�w�uGBn*�QKh8��`ay�[ջ���q�&K��c*��.X2��[x*7�m�u�0��i=8���Z���l'Q�m��˼��њM��E��+	��e���^:I�8�X���Ix����Y��M�� ,9�lc1:����՛�T������6Zk�ߵ۔7p+PHU�t�d۬��n�"��l��ܻH彆�8)Q��I���֐pfe����MV�QMp�`�M���B�9�km*�%�{*�Kf�bk`�`�ڗ�9I�h&ʧ�Mb0/N�m�Y��8Ջ�d"�d.�e���4��`*}#��h�4r�Qe]Z��=Ұ�e2�\t��l�Ae�v�uݸ�J!C4;@Ф��̔t�oL�&T�֭��TsC勐�<���P�$z0��":3_i�Z�n��c:-a�%�Q-���4m�3q�$��Ϛӫ�y���WVb���0W4��1Kv��_
;Xr6w�E�� q���I
d��@e�KU����Z#�36�غ[�nVHpf-X
ڕ���L��$�;A��ŏ,�vXM��T���4N��m]l�g�~>�^E�o#������>yy�,G��V)��֩�a�eK� ��/V^
/�en��p
x�G�'��"���].�"�Sq�0�
��8pY�ث����]4fbC]��kL�YZ�:2atͺL��S~ ����"P]ƭ"ۙ*��3�[C!�U��Z�VI�(��C4AJ��d�D=��!|:F������&�.�dKY�B��fd��Rb��:��O"�bf�4�Fol�*�N�Fǖ�^Q��>?m�E%
b���~:����.쉖�qH'lڎ�@�j��6���{�� ��)�2n��BSU�ɒ�3e��\�9b:d�r��C2rS1-���
����Hs3-��V�PV8ųs
��D�U�I�wY��m�-��g��3\Q/<��~������C�p��b[��K��d�z�`�ٗ�������/��ې3vJU)&([ �z]K�2�ZD桁��vR�lG/h�x�L
�˸�5P�D��2�Q&�LT0��L��\���Y�ƦTq�d�[��Q�{e�QBT�K1D��Ը)fec�6�Х0�Bf�\śoo:^EftD��IU֚��?%��i5�,*�o�ekB�-�Z� ˄�Ob&�0t�K�`�"��
�m��[H�4�Zxf����c��1*͜�)(]�Mm�z�!�zȁ�J�u�նC�fe"[�I7E2��i9�&S�?n��}u��D):?�qiu��^i��Il��s�U�X^�%�{�Xg!�����g�	Ҏ��`�;6w)��̊�?O&��a�Ք�t�S�Uj��YiD�D��r1z-����d$��������ieژ�#\cB�f�s
�g�
q��*��Wvv�A����
��a[f�cn,�!i;A܆�kL���b��1�3��׊������fˤ�M��Y��6J;��C�wI�Kzv[Re<5.�54��v�0.�#;&&]���3�*���F��(��Z�NΚ!��O��;���˶1���df��W�NlyV��#�@�s1d�*�x�%��`#bCsub��zt(��פ�հT5.��Qj�9�j*X,����"LAn�2�T�`��i����j�`!D��w`0�T�Vң�#o@�D<vJ��1������!<�����dG�H얷W�kY�Y���;%6�Ou�ޑ��U���7��WV�dD;��̈���e
�F��Ԓ�)��zm��2�qRi�^�7��$U���\҈�jb��l�؁�u.�\�h�p��(fu�`!��^Tb�XC#6�R
��`.|>�d��ӎLǶԱh��N�N�E!r��3!8O�3��^����e�>Y�C�#za��r���w�-ĉ���@��hLі�V��<-5�%B�-��r\U�J�B_���-�ڍma�g �QcR��7T��
��[V��t �B�R����L2��V�BX�rPWA��g��$Z��F;�pAf±��(pF�uLPo�3vm<,5�[��j�f6����Y��-��6�����h�U�p��T�Z�)��%�`�5Z5�[�7e��YO��l�[�'�+{��%�����Ov��ڈ����0-V_�>�z�AƵ�@M��vQ��S��Շ��K���`���3�8�B	�<_YXd���k���IC%��5���M�h-�( ��M�#j�T�^&�{�PP:�����(e<xּC2 �[KH�	B�;��d�*,�7�,�V�Ǵ�]�:id�Q�!�Y�;�ڑ��( m�R]�K�^M�+�u�f�0#����m�5�U˿�)�����&^e�7Q�v��t��������H�2�z,����{��GVD�m�Y#RX.-ù�-��ZH˥��5m��LςD�x�^It�kbJ���U�TV�Y#h
�Q
I��{�[�C6b	d�2XV�,�m�8e����,�!r��+N�A�6N',жX�&���#��*�΍�����´�dI��8C���q�_��{eZ��jUҗ��ݎѡ5�ѻƛ[Jkd�#Ĉ�^wYZ�\j��5��@8�,�7��D�(�u��Z�梯*ʳG$	�1�.�I3._��GV�Q<`��e���$6&^��rk�,46|i�)��� �����KrF��]���&Y�MEJE��b��`݁w�GhQ0��yN妵2�fbU/C�N���J"Y���@◀�����%+0d��|Xt�f�o��dJ�L��e�U�K���y�hCf���d�j�)X�YC.ڲpbi�/u;�d�^��5��P�>ǨRB��h�$o��/0�5���
0��yaSl�e��ۃo�7h:.�����zj��Kd���n�i�m��*Ve\6����,3Hyq;ƷG��m�ZEgp��m�V7���l@������Sl�&���ek33N�U�s��Rњ!���]�Y��m���6MɆ�pR`-M��*�'*^iM,שC�I���t�٢��\U���CԦ�w��K:4�ڔ��Ԙ6F��m%܌�/&whڽ�l���b�-^�[FVu�Z/.�\1��Jy�LÊv�;�F�q$K��}�����.�b�Z���)Dq��W���U������hk-"��mP&����sq����,M��`*����{u-�
-�+Xզ,��E1��7<���`�ڻ7L�v�m�y���*U(�)�(X�"�X�]-ϊ��[h_۠
�ý�(��G7��軕��F4m��J�F�\��E�[t����Q��0�����ɱ%�1hL�x��qJLн'-�ϔ����,W�@�PF�W]�;G^��9�1#f�Z�Kl�Im%E]Cu�I�SI��\���u��e3lnޫ�0�x�CK�r�࢞d�P#.�N`33N���H�s#�y;2K;��E�-��1���<�9݄v���*-�<��j�x,��c�jS��;�v*��q N�ȣ�Q��!�>!�$��|�eԤj\r��0(m�R����:[nƍ5*өu��A�[�Z�mU��n��-q�`�E���0�zE���l�v5��[���AE|���:a$�[:��6�X�b�Bm���B�X�W{n��h�Ҕ�=�jP�q�`	&ne��u@��>`�j-��ܸ����Y!�y��(eK���{Cm���%S%�,h�Em���F�h���[n*R�ZK�Y,�c͠�~X/���t��M٣4Z�u%U�ieY�
Ĵ43��35ȷ7b�ף�������d9�p��X��w��ظ�nR�8�'W}���T:��<qT���GPz��.���S �%N��{w�U��s߇L]}R�!�#����N]y(�7>������.42�r�x7�z&)� �[���KĈ#�d�������_����v��,�W:�4�̶gJ{L��'�
ϼ`x�ِ�S2^<��t�,�P<�J_����ف{�%��	�B��Z��=�嫋�{��.ޞ�yxoMؗV ���y	״�(>
@F��ԯ9Z۝�����B�*5+��R�e�%�D(�������hd����
�,���XF&�|-Иߵ���$�
�����+�O��[�(kR���c�c+e�u{�����*ũ����2�Z���$��J��cN7o-f�kV��T��L`\$Pݕ��s�->x���U�M���Y�Sg>O��L7�R�x�@�]vG���Y.��o	*k�l�c
!����1�@o˝ݺA��]s�Y׀" K��{(f:1�Vym�Ż�Q��4�
�E3�����ר)��e�E���D�4������aoS������J"V�ۢUZR��՗��a�<OUb��A�]�_g<M��4��z`4`웽��&�{�jg�t�jG9�݆1�a��b�Z4�ub2�T�2}�)�uݻ|!�iV�+����E�9���|7���,��/T��G��{��n��/NO�d��^'����GSƅ��Zp�m���}ˍb�T��l�R�s $���%d�6��.��B\.���8c+f�e���`�w4��Q庰�cy�%�n��-�9ȸ���=��!�#�-Nʝ���&-�RVt����޲4���y%"l+�ۨd��],��d^��&��$�|d�)!]�shv�!/��S��H�{K%�{B]|O&��[t��N	�kGF�̜�l�L�+o��b˗{����D/p����ÞÍQ�M��\ɷs4�ݹ���X�L�#�U]��H�)��ޠz3��ǡ=Xt��֝�J'�@��|�gRWϞp�V�9�Z�p?���nT]�.������;Z�G���f����ٗ4���5�gjXd_l�8���5�i!Ѩdޜ%m-˫�-��9��*m�K��$M�V���%Q�0�i���
���7�xy1�������9���cM�^6��������,�3ךDC�B�13b�'����iDeLɹ�^�L�އ���ؙ89���(N�{�R3I���� �
η�@���	1�:ʼ\^,W�ۉ��ީ#)N��E��.�f���e^��D9
���֊F����ι���1���}���:
��G�{�u�3���sr۞��b~]�*�n����!4.�]�+��=ɕ����4���
��|9k׌h[��)�2}q���V�YՆYL�P�v-�;�R�%�����Vё�c=�oG+�<;5�p��f�Y��R��ܦ2C���H�7X�3���vv`�Z�l5���5�v��f
C�7��z���E�a��2<C���1���:D�p_i�uӻ��ޙT��N>�^��煹��7C�f��p�.�J*�G�z��,�;�T|���H2X�V�oue&�ɓ9n�����ʷ�C��kU=���_>�:�e�e����+�����2���ꖝY�z�&B���g'�j�������a4�ʡ�����HɅ�w.&�k��E����w@�4��v��W2��ChU�*�z�FB�9�z�*媳r��8�	�H)�ɢ���mmF�+Ky������;Q�,����J��"�[�v�r�G�2Y�)A]F�MM�޸-�-dو�y�K�YY����s!���{7�40]5���6�2�%���^V�8E�vm�|d�R����,E	���&u!�bb�|ڱ8K�����Z�A�Ugd��l���sL���V4,�aQPF���q����3���L�h±�:�4YU/���K;�{�wّ��<�x�E)��X�*�X�a��q=2\j�x���!��j��WXc�w�Ix1���l'V�-pB#+#�ks6���}���.sܛ�6M����������`M�-���	�#)b=�\N.hPK@]�M��~�}�Ƚ��۽O��S%b�������r���9�C_�'��w_;6��7�7���b����!Ζ���(��nl�i��(*í���Au�%=�[sOM�f64�o"�(�|�S���k�[��һD��U��.R�C�X���\!���j�`[��L[���� �"�sͺt�mEB�)ա�oQ�c�;A��S.l���˭�_,r�7I���ާ�x8�����{�>\{�F�t�#v\��e����+��rN�F��b���F��p��B4ʴ̰��`��l�ʄ��{���Ec��#��&��h��W�^���/:������7G{x�ÜRw�p,=��i�0N���j+�E��9��a�}1NR�+�lwr&c�=x����c�j/6֎���>�s�oC�H���HН(��Y`zzcX,:��:�v4���K!t�2�^�8s�t��kr��gJ�Ncն�*����{-)-���E`�����	��k���Rw����r�](b�R۬.�w��vB2�G����;�搱30VE�XU�h��*���w���2��� �����.��ZzȊ���%9/b>�U�Mı �漍�.�\��4A�\���c<�Y���Pz���-�NbH�����P{[3�g���V�5�q�O��D�����7��|2~���|����õ�kQS��s�.Ý��G�)�Yư���y�L"C���8�l��Zdٝwu�F4�A���̼y������J~��61�=Jdz����3n����ƈ����RYW����Ҳ�{�� �Wpy�*�q�.�&�O<��Z^@�e��D�� ��N.X��� ���hPK�E���p��$�=�2x���8S@����Ժ;���=��ft!�|kk1�/�r�̹���p}J��fH�ǻH�Ӥn��=��{s��,�����4��<�aZ� ��;��{�Y<��.{�[�#*A��W��^�8�Q��f��w��&F���k����imÜbwn͛�3B{�˵�ӻ����G=�	���ٲW��FXi˶���vOe�>o�s5�X�u�Z�8į�;A��U:�d�,4�u�M���ke[ìf���*������b���L1���w�������\^��X�*�������9��}��e�m�8M���Dj���k��M��p�W�: �n��Fv�|�l݁�a�G�wy��s1FG-3���2g�mr��/��tR���_gv޻�֣�-ή����X���s#��L��h^��b�92�+f�4�fF��'Jˡ���75(�Mh���ث*�V0���BΖ�8��|jj�..�S�`�,$��,
�K{���J�[ܺ|;R�Yy)�H)@n�l��m�g[�o�@��`���0�r�'WnA���/�(�g0�Y{�� N�W����4�F��O��񨙝Wb�<�t�b3
���f;y�/L�N�h��<�c���3J���ײ��l�d�`I-�m}�9n,��f
t��5��r��#j1���ه�(!�C�B��n�b<�/�8�-���u�2$��A[OY[�|����\�`�&���$p�!�˞�^L��u��>���Tw�s�s�ϩ,�1�⁬Kx��:lC�{Ϣ���A�m�]���G9�����R��v8�1�ú%֚��>H��l���aA�ܣZ+0��q>�+3P��9V�;�y�Jn���=F[���P��øB�����9��y��p����v��h�  B�2������,��΁|/;�ȁ���T;rv+��agd���+h�Vj���	����/"�c9�XwF��╛�21�su��#��Þ*�Rnm��_sď�2�ܼ��vb���L�z�u�ي,q%tm��z�HŃN���ύݺ��bzAw.�Z���:foR�m]r����=5*\�qo�fW��̲
M�}��|����ﶾ��'ikw�vq���(О����`ù5��԰�H�\}��M�q��;��[��s�Ux=/Kn9�[�r#>�w��G���'�p�[Yel8�=�M���G�6_�}n��N��z���zo�d��#{�ứ�OA�7^o^XeW-�8�<��C�j:��%od��v�1�(�a��uת�"���C�DUq.�܄9��	]�}L�����>��%���z*{Nd�s!P�<�t��Ů5�wP�Ç����ֻ�Gk��ϵ��E#5Q��;�db_O��3�xwUr���e}��4^#��J�5�K-n���)�듊ҳ-���T�ퟘ���'<~�+i�:��&��V�Bťtm�Xr5��w��& D Bʏ����_a�����Ӄ�,<Es��8E�S�8��I��V�����\:F�pL��=�(�3!&A�1���
�0�fMg(�����P>�hp�V�vG�u�q�:��js�-�<�;jN%gH�X�x@#��o�E�P��rU�xQ���7B�SZ&��̢6vm@Rl!e���g���r&���[4��4�(,�a�v,�˻3��&T^�����K�x�kL�<ʭb���`�r�&)P�a��v1[6��pj���	}���a���Q��gfݲ�!0�$=�,[{ٖ�*֮�Z<AN 7nf4Nb���t��܂�cZLѐv2Jbu�Ҝ��,0�J��l���,2�^t\e��G�x!W O
v�.�ɇ�vخ��΄�\���A%���yw�
Ï�����n{b��;�"�Ҥ�k(�6Mk.�:r��p&nd5�:j�3�b	�PT���m�]q��k������/5�Lq17��3�Wb*-wk@!�nm�]١��mr�(����9�;��P�<YRri�Dd{�_��Y���I+��,e��R��_);�'Te�u�a�c*���-�W�eS���j � 3��]=�[�ܔ�1�go��t���䷖�,5�xg)�F�ۮWʲt�8�K���d�o[����&�TsGHq���/ud��q����(#烞�㳮��}�Sw��E��Q�.����h�C߰I}W�q��}.�*�'�\��t����|N��.{���m��L+7��R�uH���8D3y�V����{fEg�K,T������h" �/�5�*��T:m:y*�޼`#��h)y�ݽ�g`���T<f.�5ḥ<�ըp���B�{5K��.E�V㤛����n�ְ��w}���M�w�i��&��Q��a+v!]�� 7������K�j�OQ:f?r�����+�R�	������Y��y�6�)�,�hP3�.��-^��x�P6*=z�=�O����n(#뽙��G/�.M�.qbu��Y��F�fc7�s�
�&�k���M���W�_!���|9�۴��WmW	�l^GgI����~��V��#v�v��W�NJ}�Aj������l�6�a�{J�F���涰77����8�֒�w�:=H��h7�_��<agU�[u]�Bh)|���p�ӛ��q�|8^�,��s=н�mK��b'�Efn�k�����b�ݐp��\S�
���s��C-v�
c}+�}K諉�r�e�H�}��I:$z�;Zo���)lp��:l��F�qu1��h�%�z��&1#*oP�:��;�%��<3W�\YK�<�G�,�DVVj��8F(�Vm�YC:!c\����ݬ��~j�jm���I�!�ŧ٭�^�U�Km�����ӭ#Y�W�S�q?B�L�H�VT��q.��"�k3+*����LV�Љ��qۦ-d��`N�Z�T�}V�v������N�t�<�1N�������u��u���԰̾緛5��wP��|a�v��%&�5}/`�.�E�)m!b:'�@�vb��R?Ws�V}�����T�a#�(�EV��!&=�"��v��
<8��E;1��9����W]J���1�.��U��V�,���өM�������"���3���=1g��a�:u.�� �ZE�n2O�؝r� /�zDa[P	�F�_=�1H�3{���� rj�3LѪml�+���a��v�;��|{z�n��B�y:��������̜�-罶b�#"��#	���==H�1���S�E�inp��ק��P�������6�R°G�MX�*��F�eP�?
dE���6�r��U��v���$���c�9��c�t#2��gLe����Wt�{�8x<�w��2+�b���Y��3`h�70�#]2�x]�//we��a���g��m��M��(�O�$�<��<L��M�{�%8|`8�r��6��b�'��,_:�������ţ1Sf�����AMC���@- ��xw{�*4���z_PX7I�������Pr��}�糷��еq���eJ
�/b6v��^�]��.��C���C5s���A��B/�-�gף܍ң�F����])[q����z=z�ef,I7:���h:�P	��x]9�m�s(�Er&4wZ<{[�1�U������"_-��s�l`(ë��ގ��6����gm�ιC8O�ޝ0>�FⱲ�D��t�V;�@�.�֞)ԟU��d9�wgG|C't���+Gy�:�q��T���l ��!��u��v��۹]Iנ�i���������sc�dk��ui�tɹ��c�����\0�x��/<��v��m���5ޔ�6�����6��~|���?߾�8������ ��uʘ2J���l�Y�,g��+P�h0Kr��)�݋T۝yԏo	��1���EĊ���P]��pghFʺ{P��!;7�0c��)�p	yk���Qp�k1F7�w��5p�gBݪ���\�;u�ӌj"Z�X����q4�}jɂ��339�6�Q�'^���s+�`H@�pv�Yl�,C��Co���3ؠ�DO��:��x� k��3u�05��-r֮+��:ݮAaZ~{@�����׆����$cɷ���Ӱ��#x�Nu]ܢ/�U��6
�d�KZ�W�dbU}�a��pę����JT6�YB('�l�]ZB/SY
y�m$	���7�s	Qa�C�������x�����uD_��ův�q�}��)�敕�pr�V�m@�	[�
bd�������F��mj.���IY�j�)](e#;/d�J��P��?�\V�V$�q��!1��Ӫ�&v�f�=jfϞ�%��	�C��\v��|`�N��.�i�F:����wi�/�U��j{D�Y��иow0�B<=�3~Ȝ���`����Fd�{���O��İ��ޞ���۶����`���C��8^�k3��Es|L/'؍�ɱg37gN
��M��DC`cSi��6�M��^�$%���y�esunMZLo,�j���I�w_G��6��"���yP��@����0�~�/�MY��D3����Lw�f�9���N^qŹW$*�D��V�(�๩���^�=�n��kr*ڊ�Tꦧ�6���]:a����g3APx�f�2ep��"z����	|�|"��WL������.ك͉%���ω�����Of���(]t�Ѝ���3[gu7{c�'������/n�X�Y�s��[����RagE8��&�;�Y{�o{�y�}i��!Y�"�3}j嚽ܛR쏝6�j��{̳�c�����C�hF씲�I�:�v��. ����Th<�@�(ئB
!����T�*-�&���6����M�ϰ]k/Yk5b좫2�fe�j��B}�"�(���z����Ô�
�	�jp�㨣�x���Dn����g50���1B�V�i�S6lP�
��r�(D�n�1�#��BWYz*(�x��W4طx��yQ;a�cݫƝ`�ļ�M�y J�ofu�A��;;Eb�H �c���V{���O9���^�r�ƔXބ� ��+�&����]��K���������h�	cm&@#%L[��̅[|P�4�]��[����¾�A��#&fE��P�t��S�.�:�<�f؆Ś$���z>�����8�L�[Xt
�ճ#���hpR���Tu�ȱ{�VƇ�O,b��t-��cT\)h��ʠ_�u�7�ԩ�d�v �^��L�{�V�v��/@�a�Y,�[۷��y�Q���+a�[����ik�P�L{�3���l
�Z^i��s�1�x��cWv��)�Q�GC�wn�)�V.@��!��ܠu�B�A�}j�*!�A�f��]�D���&���G�J��sq!h���`�#�鈧!����]�#3^��{}�T��2�{dh��lk���Vf 
¶ ��f��Wm�R�K�p�u�ƺ�]v�P}��@2�\FJ�����{l��4�Ij�Fe7�Fr�+��z�y������iD�� �kT�L�0��f�F�gfԲ�m*W*kC6�"�t_�9��R�yث�׻�9A����	�j��NqGka؉ۺ��gKc	;��5�ebT��e�@ $�γ�w�f���$�Jd�G��v���c��t�kgl@��is��+s70"��pۭ��jS���;�	b!Pv!@�����Unۚ�cX3����# ��X�.f7ǚ2�Wr��܋��'p5{��Xc5�����h�EP�}cT�me���M�y�PS[Ȥ�B][gd�^��i7�vq��*��O��5��QN����a [T�UCF��Ȕm%Y��KÝ��u�9�@[$5S4��'%=t/�46C^��jh��Ũ�����9[b[�΁��E
��:m��r����7w=C�����dS��ܪh�4%ֹ,i<=M�>���<�� �V-�[�Z�Q����QYN�]BuHT�/;	��d��o����փ�n���w��I�5�i8t�̽���4���^|��o&!/:(8k��.ݙ��5]д�;�H���h��a^X\4�;��.̯v䌽gf���9��_�4�g|��`d������-[22��r��\��^���ӿ4��w�ή G�k��֮w�²U�d��$��9���~\yg��N�t�=B%�E"޽�Ej�v,dS�c�F?uٻ�k�/����7�y&����1ies�̥z���T΅������<S�5 �1o>-o)ό쳷�`�
��4��|L�ek�ύ�Fw��1w
��:��O���K6u�I�e}���yt����0�GNqE�KeJ�b���w�AܢHgN;c1��H����E	i<�[E1%�xbdpE1dU藩�l��^�#\�A}���q�Tp���:���C�]�Mn�j�\�Vk%���E-#�S���c�2��ޞ��JzF�{&,r�;����$՚�F���;B������$�1��DMf��/-'�[����va��pb�m�A�SI�����,��� ����>*�K96����K���ʲ���lѠ�UzM��-'������bC=�����x�ٔ*�z^g��1LjB]��n�{u�cuy�s��J���ڞ]�\Hwu�^��R�� �\G:��:B;��4��Gt�(��2li˧ˉ����Tέ����bS��0/�.��>���H�+�Y.�����v����T��ǂJg5{��v ����L�"�vy��*��(4v��N,P�w^�v��(׻C#�tX��f�T�Pdwї�r�}!��b	u��n���B-+D��iM�2��s`+q��'�*�s4l\F�3���&+�d[�Q�XTG�hc:f���K��8m�M�u���ebV�p,�'K<j
�,�n�'8�ݚo;��h�9ֆ�t[���ĵ�`�}���/��6��]����)o	o�x>׆��A9���Dw��f3�M�ĩቲΔ�\�X�;�y��l��� fa�wٺ(Ze1ƇU��ND��vd*�
�X-��\ޠ�u��V��7���<+��4��,��C���V�W��hU�qdU�ƀ��$�i��c�>W�u�sx���v����	�����H�=��ێ�aw�E:�w�N��s;#��/��k���-gMvP2ĳ��Sa1���-+�0H3�R���诪�Z����}MJ�B�<ytB0f��P�eݎo(2�v�Ժ��vi�gFA�ʆ��{�ɫ8Y۷�^S��̓IH��B�S� ڕ��|��\�qɽW'&$[�z��{25�h���1����*>F�3<yv�v����s���)� %��3���r�|q(e`��m�`V��n�<�enjs����=0%7<<��eMoŞw|�[�S�.�􋑾�#�hu���t���7(�����Г��ܮ��҄����4ݛ�[�MÊ�'m����Q;��05Y�J��e�2�R��8��4�.P�G���f��	/�n��f����F��ﻗbӸ���i�g�	�x�����teyU�L~��e�Y���F���v=����P��Fr���S�0�e�wX%(���d��Z�K�e�/Eh���p�ܗ��5�wT1лX��w�ɵ-�v�=Z����#�{�2�{Α��x�>�貗�	��+w�c�")�Z�˰^2����7����v�)A�k2uCQ1V��O-sU���ɷh��M��]����;�����|"TUv���w�L5��Mʃ��GoYP����5������t�<v�B�����B�:�~��x1���]20ur	�f�u�Dt��M��GAʹ���,%�^<��,'5�v��[ڷa�����&@kU/��+����i�GD�XM�WW�(μ[A����=�4����)�h�����ܫ�[���%mw���,U���:m�� �@��<�2���v���šdX5�[�h@h�$)˹L+{C4�E�o�֣puǤ�듹S���:Y�ֵ�ppS�v�0�X��!LJa��c���5�2_���FSºcܟ\gn*�۩�g-�(Kp�.�O��5,���%�J�i+��y�a��/�v[w�B4�nK0���6)�&�
��)����t4R9zͪl����eryq�
�S}#-���:�C�b��]Aګ<:���)k�TF���z;�����>�}����L +��1k�lelٝl$%Q<�т�~у"ټt�5�[N])KF��G��ꮅ�N2m�Q�9o�U*�d�0ib�9^i9�E�����=ݕFX�/a�\�VF��$�l<zo���<N�e������q���69"��M�x� [�gE�0���pXnD�������{Αl�F�o���Β�z�]���Ӷ��|t$��b�'�w���5_9�*3���Ah�+����'����f��q*�%�4���ΛT�I,Kq��,�[N�T�<9j&�u�:9����! �ĩ3�֯B��}�AuiŪ^̋4�˅��e��X�<�<Gc	��YpF|'n�\����3sP���3w�/b�Pݹr�R;�\I���^U��D���̭u�K�u�k�(w����\S��`ʴ��O�R��þɺ��i���Y���//!���0=��֬Fmv��rQ��8�uӐS륳ݮ�Ԗ6���=]x�c����՜�:�ɳ)���r�y��:�(��-��,'\���	ӫtA�
�hҨ��\��N���n�;$-(
�ѬuɄa�koUٙ��εku79��c0��z3Sw��|��������Ʋ#�2�1��.�Ϯ	�_.��,�:AO:��,�[��V�
��!VpU3�eES`3
��#�}l��G�O\2�(&���N�8�h��j�Bs�-/���6�K��b�D�BQ^K]��X���\��cǮ�x����� Cލs�۽�y�	�Ȉ)��ܪ�f\�)0��3.�&'[T��1FV%���J�3w��9*y�E�h��X����m����"��E'IOin$1��p<j�m�{,>a_S{qCoEr��>y��})�g�5֓����:X�����Or�����w�+ʋŞ�v��=�J�!O�Ib��W?�-��s)�"��E��E%�]�{K��L�9h�'�g^�ˈx����)x�]���Su���/�ܭD���û���i����xGgX�Q;���E�I�ū��\��	�z�_5�M��ld�`�-��Θ9���au�S�Wg��ΥmPL7)�yg��7X ��ꡎ�7����zTB��)�%M�X�jN�bh^_L�q�&]<pI�*�b���!�*���I�V��F�:u��N��b�:�X�j��Z�AQ���Kב���پkGI�oj�|m<f�q�%J��֖E�5��j"1b���caL�:�N�'P;��8<r�[���o���1Y��ﯨ�(�⎻]�7+#�ր]�o��i�Yj���9�4�A@��T���Һ5�G2^%R�~�P�:g:�s�P�� ���Q�55L�[�N�.Ô�"�p�e9z��4c��w3-����%VXǕ�{(@�
�0�ɘ�8-�ξC_��ڕ�[�W���6Y���;���!\����m*6e 	��Ⱥ��*�t�2m$mN�A�V	4w�7wP)M�@����������W�o�Z�0K M'���o},���P��Vor���k���.�@�c;�� ��(��ur��Y�+{
�\KSa�r�w��r��1ܙW�ڃ�eS�͛lqr�6KiX�,�Ӆ|\۷y�쯦��R����cݭ&n����^��QŗD��;w���@ ֈ��}Kc��Û,`�R����U�%ۻ���QoY�B�:f�A>nT)З#@X���F����t7m��K
�O��ȟ<���G^��-S�,�J���]�[�sB/j�@�e,ng K��2	��1��C���Gw�e��v
ƀ�Y9��T���۵�Uy��Q2�B��
w��FW��S<5e�:#���,5m�c˯}��p{wQ����:efWvXVpg���J�t�B뛬7 y��,k齨�능�婜��%;�0e���!�OUn+Sa�
�X�9B�����{mZގ��]r4�79'Y������a$�]��X�Vn��U�x��j"4����Sp���u�J�ں���)�X�O��qg���`�w\�t��DV�ewstn���H��ε�C��,x��B����ŵb[�lȐ&6�$�
W�,�w�-q���h�
r,�	^�U���wrVƲ��ّ\`�X��w��Ե��Skxq.H��6�+U9�ckj#Y�k%3V����7d[I�,�'_|�	V�`�nލg"�6�n�(j7%��w���0;7V��	�op ��m¬vhx��K���3��u�|.m ^��}<i�sS̝p���}�S9�@{vx���Wu�:�;�s�we���ŷ���wu��.��*S�a����,���n�:�J���N.��@�wvo�8��bn�Do=�j��3!��.��QJ�tI]�C���A-'+R�nqg������u21������%<�f��"Lh����� ��<=�<=�z������}d��@6Q��u"�ܬ)6���jS�3��KY໢�a����,(�P�=sɛ��Avk:('N��᭾m����-�_E�݀ޟ��������n�s���iՏk��U��8�ޒ�hĥ�R۾��i�Vne��7A�����=�#ږ3g 4*�dóXo�������Cf�%� 'B��%���V�p���լK�c�Qd���{�b68�G)x<{+�}S8��>�it�w�9p.}˶v�]���%#(�0�Y���� �����W�O�Ρ\y��Y0���9ϭ�PM��B��<��Cŭ�y�![�mM2�]-E(��]��`�/�Z�7Y6ڳ3L�䓜�/��5��t��k���j�g�;�+;b�y媳
��C�Ŋq���J	��f9Q>d���뜪`�m���;��#���iWA@�!n��ڱ�]ǵ�*�]�nټ��:�o�'8�kH9���v�h�����8�N P�;Phq2V[F�j w^
�y^�}�NDSӗգ���C� E��.�e�,��9��6r�ӥ�H�y7 QR�r=rs+��R�bb�uBZ�`��p�'�Y�Z�����i猴��P��;�Y�S�>�r���J�ag�����'��pcJu.���r�qu��	�cu-�s��f0B�;V��ހBӶ���yxq#~)6
d�����X���U.��;���+�G+R��p�� ���s/+s�%E]n�wu�P��r=)T�I3+B���鉭"��N�s�'��c�EQt��*�wB�β5��x��On:��B��f%���*�)eQJ���At�Y�wn��rr�T�'2�"dRF璎q�SR-%BU��3[�⸸�T:����=r��W2K,��5���L����.�)"�\<��	�32��fNHT�<(�swt�Q����t��4B6,��DD���'�4��i:��� ��F���T�*^���8������DRf���;TLR+,��p�4���z�څ���;�M�v㚙�DV���a�������SݥI�0����Qd��^���A'����W�5��G�%\T]V�0��7���K�/f�7���`3�/����qj�ۺ|��0��=
���S�Y�!w�g!$^�]�p��K�+��]������EoM�iuH�D��Y�o��״�Q��֛߮���6�}�hXn��(s�{����R�?Oq�f�,Ӛ��a6��o�|��d?c�l`�¼6�\6|-}�����p�җ�=��0;c�s�Z*Qq�j�D�'Uõ:����HŃf��c �d�M� r�=�]��V>S�:~q'C'1J-��
T����;�7V;��x�;�Ө����yō9Ü�{���[U���tְ<%�`_:L�Uξ�M��W_f�W:]��i��[�b�-�OT�qQ)��~��zX�3�@\�����l�QnSs���b;�4�����e��CBNW۵29�6�O�y^�X�k�'����B��.��彣��3�9��R�;�����9B���X?u	���:1LY� �jRʃ�����J��tK�;��C/�i���u� R+A��m< �Pվ)nzR$�3:n��r��0��p}j��SÆ��U�˵cZ��Ҏ����s�[]��P���a��օ�(/Qh���WxU�w/��F��B��S��
zv�n�}���4r�]n��>���;
o���3wv�[�{G�-����A������s9�F�V�Ȧ��P[<0[Z�#��F�pq���sB�%��u(}Y�}�H͊��7�9U"I�d�N�9腉��_ �e�븛�z�'M�%��wP�}N��S{U9|�>P,��Y1q-WQ����q�W���ɫCt����7��)�HX�F�ޚ:O�{a�B�>��h�9�����WJ��Ѩ��*�&������*Aʂ�.�4��[�;_t�VK�Q�\�^~(&h���
�C��;�i��B�bq�t�����ev}ٳ,�d�M��˱Q��'Mq�!�YC�Ʒ�S�^N���';��}O*0�N�:��<*�ھ�;=�����Xzʳ+�4���l�靊|�R��Ky�ڊ�f1��x���a��_:}������X�c}����Wmm�}��u��wJ�~����M����7z��~u�>FY�g>�:�bښ���S�0n/���k�]��;�]u"�2x��a��)W�YQ��e2Q�7��HTa�E�XxMwov#����ZN�̥m�7�q�[G��=�o2!�p��o�w�����՛:����T�;�#�Vki:�ceL{�.]�˧R���m}��� ���ݫ/0p�DV̙�&`��3�f��8[{3F�W~���i�4��M�t��If@p�9�Ef�z�Ol�5;,��xZ?frC�?B�����Fˠ���t&���,��߽4��k$���޸k�.��T�CpA��&�������T;Eܔv�+���^�e�޼�!�m|�4�`�+����^��h���N
:[�A��\Gw��7^�H���;�9o(�qJb���;c�p�ϋMT=�6�D���*5NMv���W\�8[d�̰$�d_�3��qM�	��cW-O��{*XC�V\��<�f�+Ϗ�k%�0P %8J�c�Y�}��>�ӿU���>����'�����f��sp����܉�3��RV�cS�y�Ϝ�ϽZh�7��F�{{dݝ�ƕ_]YpztCg�`75Z4 �L��2�]�@�:)��v����2���S�dqz6��FG����u�'�x�r�er|���¨�[���aOn��<<9���{�o��*^]k�z��Zu9���xT���i٣m�F��U�:�
%��tx:��K@�fO!�
�^�t�����g,��f���3Q�2�ϻ���u)5%�ɤ���l�cw�����HM���+��w0ܼʳ�s1CٗB�����DGBo\�2��#2���w��Q�+K{s�����1n�����;�Ӳ��c^��Sw26�=441����uT`t�NX�_q���
Dt��p�&���fsA��8��!�l}�;R
�g]z*�x`�v�%o���g��{z��NP̗)ћT&���
/�1"{��EFJ���pž�(nS�V����>�mb��5�*#:�6�K�]yf{f_u|���GJ����Q��6i�B��c�-D��O�p"��n�{Y�o��B5��N�HtEe�h�T�dࡈ�j�ގ��P+�Շ��7>K����{E��ߴ����M� �oR6K��r6e�q�a��r�`�l�1���Ŋ�B���V�諂���x�:������< �Hev�VF�_V��q�g�!�ph�7k��O)T⫦����t��h
��|aZ�#��y]T0}Ηt����z3�q0�^:m�rl�o��R�qO���^��8v�6�.1%7�?�~ ۤ��WpY���?W�*xl��ŉ����p�f9��M�ީr�Ҋ���2O��5Q���BE,d�����+~�s4^��;W�.��j��1��[o"��hSov;MM�Q�|�"��ܮ�ѓ/�;j�Z*��L�Hsj��v�Т^�0�z}h���u�xy��t{ؐ��0G�<��L��闐\����Nc/"IJ�g�����؉�*�6��"a�R���u�gq���9	��H�sH�$��h�:�y��s�x�*��♶rOnf�ʆM��p�5���d�m����͌"��}A��}U�f�jFZ�u/K3\w��I�=O%5Dx���ۨcqa�|~���[�@��y��B�L���k!7R�u�}%LIW��&�j��q{M9Y���V{��u��sT�y�Y3m�͍ж��neM4���`���x��༨��պv�1��F��Q��ګ�x(R���3�إ:ô�Iܖ��*�@v~��6��ƅ��g�@��;��w
W��/rm���s�z�U-�o]��Ή��K٣�5�cyhB>-[��/B��y�,O��&��_=����_ܥ�Ϗ��̯1ֻ۳Ü�4!z�ڮA���jٮ�ٔ��Y�h�(�m���	��u��$��r�Τn5�×0�'S��D7V;�s�tcʝ+;i���8y�Fyshv@nŉ�G2�u�^��t�`_:L��i����gr+����������{�"�gΣ�9�q��:��Du�E]-_iaml=�ӽ�7�o?�lw8<	(2���K�f$a^��N6Ė.�ް�:�~&M��fs!�9���e�w��ۄ^٩�pΨ�����F��m8�-�/��g�Z���8������&NEj�Ȏ.�}al�_[�����L��6���캓UJKb��Z�4m�*܍�q'���WW�=c��.,��d�bU��~[����VA���{W=��~����6aʖ/Tx6|&���ip�U�[
������B�oe�O{.�pОJ�����_��P��[ �<z߭|]�L���A�mV�o��f�c0G玫YȊn�4[<05���9Qϗ�}��^4�AU�:�/Pc&��.�z�(�)��ZH��mN�S�+�N�hϥ�\{(n']���]��!�)�<��
W}��ܟ�Q��T:�:LL�}s�1�A7�W ��1iŐw��$�[5k�e����d�j�d��^C�>~zE^Z�S_԰u�V���֍Fp��p��ǉ�lN9�}��F�&K�t�y� h�l	�T��GJ'����=?I[X*���v�Z�Z�µN:�X�CRx�iT�n�}˦$5�̚6�`o�� u��%}���tmp�C��G<ܞ�25��ʟ�F(�ww:"Y�rpv3�;v������qļ�%�����K4��1sS6�*���23�αT4�2��y�xN��_���kJ��Z��
Ag���:�4���=77Bs`�8�7Ӓ*N&���b�ʲ������z����\�c�����Ϊ�N6a��WP�wh�>���k�v�����!1W~s�wz��-1��|�9�iy�q�`�炭Ү�bS�\L^��f�9�ێ\�Y��YV6�Gm�c����Q��ǜ<��g�0�30��(�9gZ V�a�#=�s1���y]�r(�Z��<-��ScBJ���J*�˪>���n�{Į��~�i�⯺6(���0��Y����^�s�[��l�>).�a�E��veW�MxW�Ú=�=ܐR?��:M|��_k���g�foΣ���6%ND�UD���e�>��t�j?er£���ɹ^�T�u�.���1��!�ʳ�ܶV|���"t�x�) �	��0]L�9�[� �pWK�#�E�Qf�)LP5��k�(Z,v�5p�"�?R�U�f��Ɨ����H+@i�b�PO�_��Ċ�K���_<�"�T����h�>�����p���j��TV����6͵���0�$�$�I�c�Y�W�+�-�pY��������3��)#?k�t������^��tN�j�W���^��5ꏽ�2�
[���s�q��F�&(�٭eĮ�.�q
Z���[�:�ZYcr$/T�8��)@/�\��>��f�	��,Nf=��}a�j3Is=֖��t�u'�k!�ޅwK�X�wl���g��pz6��D�?!�%iV59��ڼ��B�S��Wstu?&����$r���9X��h
lA�I�pԤo�`<#�:�냯��w��J����XRٽ<LeG.�F�9�ŗ7�_d�%�F٠"QHw�2�BڅI��O/��^pssH��h�1�V�N�;s¤�4����#]������=�C�����S�ҷ�����T��. l��
�O�4dFҧ���6�]����� �S)�$5@�2dNQˢ���dhV��t-Wl0���l\+۟w[#&午�T�(7oa�m��oT���om�A���P/�4�΍
vx��g�Gu���_�`
��0��s��6R8�Ax��=��g�Űz�G3�_��h�WQ9��.�:X8b�;3���㚉b�@�����:����a����D�i+`)��%������29�Ä�yFl�[4��3�i75]򹝣��OPJsfXZ1�2����UC`��j��a�]��>U�
�S���� ��*��=}_+�܎Q'�e��yn�ĦwRlK��
P�'P���~d?.���%�s@�,6��X���K��j��#á��]������٦��}z��gc�|�M#U�L��=� �/�o15]:	�ޖ�E�]��|x��v��8�^8'���T렊�.�,���*�:B-�P�{�r����l��S��9��^�mq��#O�V�T/[���V}�DM���渘C���H	�e�����m��J87GK�ĞeW���L����IG�}��}8�t��K�"Y�� 7�Is`�#�c�t�p��F�ʫ�I뎐�(a��0�Z����q�ܬ��Wֱ.��	�U�e��e�1�q96�;��摚�L�#�<\���u��n����~#�(F7�F.�S���$����ٜ2�LV{�5���m;z�.����"d��u��7>FXa��7�]l!��e�"�+�u�O8s�>$��X�w%�1�'�o���Y[f�#�ȿ�]���|=3����뚦K��P���[\i�w�/���v8�Y^�a�D��fj?[
s�YH|q�ٮ���g�����n�ӎN=��q�nXZ���þ��OT��P���;��@�<N|v�0&��s�DD{�Q��>�y�%�]ū�x�wv
�3�x���,e"��=Nj�{�'���C^�iNP�*۫����Fa|.	H\��Nج
-n���f<��!�M9�e>�/�۸(��y0���0�Fs]W�1��BACQꍉ�	<v�GFN<c�]~S׏{������|2�ףa����^��?s>L�(c��.�W���|��ӝ�ٿ�m�ȘxPNgQ���\F�i�(�#~c���ja�d`���y�lh���\�e��$����:��n5��|��^���:��܋�
�"�yJ����*L��B��ѕ/.�{P�,*����0/�&dt+N�.�:U�Ev�B��G����H;o�G�Gd诳r�M��JB�F���(k��U[(�3ܾ�>��#3��
�&�[vs�Z��}HGZ���/��BeEĜ-�tW?�,U�U�� ���4-��e�鮎���J΋����?0���f.*cMN��l��������+ګ����BG��q�a��+�Uؐ�z`q�١5��o�s��㑧�6��\!d�*��}�@bk��\��(_Y�E=վe��8��o�b��r)����k���Y�~�aJ��Lĩ+XuՏ�S��Zp����&�*6g���tGF'\4�U{VK^�l�]}_&Vb���Q�L���I+�&���b�Λ�!L��)��S������ΰ��ǭ[��_٘%�s_n���Y�{1U]b���8OE����YLK�0|w��$D5W$f�@̣��_Q��)z.�Q"��N�v��n�IC��ov��t��&:��j��(�K�wۯ�١I�)eX}i	ִ�{%���RyB�\k�pw]���-^�}�5W#�����]�}Rj�W;�\a)ȅGǫ8�mAw�m��I),�1�W���([8�����U�]�NPu��R�[��c���j��B����G�T�k�y���Z�B��v��m���єa�, Х�q7���2+;���Wg{<�%`�'^=�'���n�;���s
�����]%n���F-�#Ȕy���S�aG��4,�����g��U��s-��(=���2o<�25����{�;H����Av��q��í����b��Q�Y�Pߕ���N���T�i�*օԬƬ8��k���A�VQ6���� i�h���M�	Q��s�*���9yx��֊�˞8�Al�������N�Z`Ţ����iC6̷wb�X��/�W�:���wk�e�O��ď���fff�׉�Ruܺ��˺α���d����3v�ۜ��>w�\ՙ�m�`��]�w��惉�Ð�6e��{�u]U���喭4��:�ƭ�q�O�th��9ݵm�5���ŦU�����F7Qj�cXF�L���|MhUR�t�iP�󼳽��N��Y%0��E�;�"�v��r�=w�el"���ףe3q���p:�վ꺻a*�Z87Y�;}�.�v��e��{�Ё�u�G��H�n���6e�}�7	vP�Ζ���6�t��/]�Х�W��)�FFf�9���1��ZW���-x�.����A�~L��.�h���,�rڛј_�np ��J98or,ڃ7Kй���+���[=�i=�X�o;O��^`8��y�igҖ�r�$ꋸ,��NGh�D�;��3gk1*Z�ٳ�ջ8��(_[lt����g*P�]��[���D����(��u�A�'����L�:t����,�i3ƣ�̰*��b	.��v��q��t�hm�"н���j��ME:� ��f9��B���	_aW���ӯs�uy��冪J��]O��GY��xo���k�V��t��/�[ݣ��z�]큲�	�Y�Yo���K����	���-�WQ������v��bgu�okk��Jk���V�wR,�{������Y�5c���>��܍��P��wQ���nU�j��سtu�b<;A��a����I�K�}�9�z�<�|� ��p����a���uגf��֍wqQU-U���k����-� ��+pQ��r��v�z*�U�n��v�]ڸ�M]���r��T�<s�k��y����,s�
�N����\�>�H$J����̌ʪ03�,�*�2�I:J!���(��4���*�6�IL3$���E���P9��&��i�Q&e��sS/A)�̹��+�IF�JVZde��Ӝ�"���B��D�e�ad��Y�F��烇(L˦f���]Br�j�(ɑ����	�IIeΨeUh��(��"�.�(�D �4�J#KE�2wwK�ۑ4���"��*��X�d�iQ%��K�20Њғ���IEI,��T#��ҳ
9�i"iJ��T�9XHU�V�R*�6����9z�J�"ʭH��H!���UBf[L٬��Z�Q�)H�*�L�H"��-Zi��gQ�) ���BR��B��TK8tD��E(�4��L�j��!b��J��(kU9ԵQ	�h����V�#D A��)M�f����nq��	��fD�v�{��1zx<'=���/F��{�x���$`RXY��M�f��#5[իt5��tr���<	�|Ns�L*���E	?!��4F'}~���nNL/������ d�=D���!���(��|}��e�}�@B"��߫������D����~��D޹�&��Οb\="4`��ʛ�����v��'��<;۵[�_��0��{�
o��ߜx(�p)����>;wF'z<}��)�7��޿�pxw����.�����®��h���C�h����3�����^�^�$DRa��<�2�'�nv�}�ߓ˿�������o�N��t�}��ސ�w��y|���w�<�[�מp�GN�o��9޷G�
�\x��|O({My����?�^���9]�o�?|��C�S�~��|w;����7��
��������������v����m�<��I��}���������r������ׄ���o��z����B�2}����tx�n�pX�G�}�Y�����~>d� s�t=��8G� +^��}��ig��+�F�O�>�ߨa���C����e?'�9����x�������y}�yNpy>\���ohr
���4Jc>��o�I�ʐ���a�)��n���x�q����{v������;rr��|���������-C�~>������aG�>���^���>'�h��d� H���;���ȼ{n��������(��8D#�'�ޓ���w�������	�]�Ǌ�ۏhra��y��e���Wp}Nw�k������k�����'�=���ϝW���C����Ug�-�
8>ʹ뻹������$} }�q��]���w��cۏ
�]�տ��yC�k�oG��w!��raw�=;�gG�}C�aWy?���)�!&���'?SuH�q8��^��]qW:�7���#�#�Dy��Կ�ߓ�s����a�}v��=~��}v������{w�|v�z~!ޭ�;����97�sɿ!{�x�xw���w��þ%��O���?g�͐���}>���d3E���2�����>� �8� 3�J��<щ�_Gw���';y���þ���ѿ������U?;_�����$��>;��<����oO������{v��\o�xyۓ�'i7���������?#����3y��-`����U2�w˺��@sEi6�(RWݗ��.�zرׯ�=�.�S�w��*e�D
�Vz�����ʃ8�B�:�le�;��+�����M{ƣ+�5�ܒ��҇eR�\^�+.e����1�֍d�'����<�݌]�{�dxL/���>�yM���Ox��aM��>_��~v���t�?8����s�~��<;�~q��=����=&?�9|8�@g�B� ��,�}�Aټ������cc�ӥ��M��Q�G�G�G�x��I�V��{Cǿxv��M����=����*0"(l��� Xߟ�#�=�`�@���(O�����#�u�~?X�|�n��Ү~���~G����G䀲M�	�������w[�ԜN<k���~|&�����p��S�3~x@�<_����ߨi�>� 
!?���>#�|G��?h���c���{z}�TΪ�y%�=�G��G�#�<�#�y�������0�����s�M�@QC�;�����Q�<u�����ۓ����˿�[w���z���aw��-��B��i	�a&�lS�V�e�ߪ��$����}g�G���E����Y�߸��	�v��[��<&�'�y?X�~�'xw��-���<�G:v�}g*�������<��ѽ|������"<#�j���+|?n�kΝ����O�#����'P�dx�߿P�_�>��������$��?;w��ǀ=��{v�=���S|Bt�\w�ě��
"��ˈ{���gޢ ��Y�4�'��ȏJ#2�OՏ���7Nu�����_��χ|�Dz��@�<�p_������9@2�H>��w�yC����	���~BOG~�<z��N'��c���I�ܞ��>� ,��Q���}����W�g��U[s�~� B<� ~	{�,�O���~����Ӽ;O�z�~C���;���ۓ}w��{���ǈ�奔~���q����~�����>P�=~���������^���$�G��)J��~��������}��<�y���� ϣ^����<&|C�[��zC��ߟ�O�oJ�ӽ��=���?;|y�S�7�#�޾�(a�|@G=�߫��2��G�=�������P���`B��}�\f���e/�~��{v�xd���zv��{���.��t�s�'8����{O	��S�ǫ���&��ɼ��{C�{��+�#��"�� �#�>�O�}�#߈��������
a���	��͋R�`�_�������6��r�G��	c���E��pn����[Z�#j��^��/i/+�^y�T�Du󛫹,�m٬tC'd����@N�����y�^n���'�X"�����G]�y��p룼��v;a��}�y�������Nߞ��?x��]�}��ߠ��;Hx���yq�Į<����rr�-�1;��������0���-��]��P�o�����p�">�N��C�>o�Br�comi�<6���G�_{��Ъ��������7��}�ǔ¿���z߾�7�<�����yw�i7���;s�yq�97�.���_��97�zy=���>�>���v"�G� ��y��|�V��'8?���~Nq��9=���xWe<z������󂭽���˾��s�ۓ���1;��n����P��U?�����|C�<���Nܮ��y�����_�;���{�ir�u�ё߯�]����ohO��¸����缿]�'|�O���o���xC��o��&��>w�w�iP<�߻�o���~v�=���yw���������90��|O��@�G��ob�G1����v��?o9��/�g�>�<�>@g��� &��Ǆ��[�&���#���8|<|��);}{�o���� }~���<�\.���z��S�yq�ā��c���xD��WR^���b�Y�����|��y����<��>�&��CӼ;ÿ��\J�BM휦��P��Ǉ���ԝ��xq�?�	�>Lo�O�ޱ_}C����{�0}���ܩ���`�dfj���� ��;��pyM!~����~�J�S~wǟ^,yC�����q�����o�N�㓜s��Ʌ]�S���~�*ǝ��c˾�Ss�����׃�a~����v��r��=7�_+�ˬ*��]��q�!ɾA�}v�w������}v������o)�!?��`�U���僟.ܝ�`�o�çj���'������C�t}|9w�iD}�微B=-gfN�b\�c��3#�=�å�}�C�������#�'�FU~�?��C�=��
�ɧ���;���x��/�����	;۽o�x�o�ܛ�}Nw;]N�XP䝿�F#�g��]5��wU�W��BH������|�\.�y���7�����'W� ��dߥ\C�B�����������ސ��w�}C����q�	Ǔ�������7���G���v䈡���o��c.=[���^������\Du�I�u	��f�J�_'��Sc���	�f�۶&eH
��˳���7����L�^���ۛ�b��b� �1qǽ N0�1�,��>u!1*�<��z��ݶ]�wl��_{�k�*�^���x||!��G���¾�)�97! z<G~��'�yv�[��m�<�ߝ;���ɿ!~��������S|w���=&���1'�߻�o�����=�݅ޜ}Nq���aGI�A��� ]���9��#� �޸<'�<�o>��;�ɹ���NL.��aN���L/��q��������;r�˾|����$����޳�>�#߈�?9^���> �W�`;��\��r�~s\�4�@Ç�d=^���xw�j���}����N�q�χ.�iP�X��zw�<����S��6?�"��'�+�!�8��|4v?
$��G����a�#��6�u���n�t����+Ї�p��G���_}~��ۓz׿��;_i�}��~BI��߯{�hyw�i:������?��7����y+���������=X��>�`�c��!Ͻ����a�&��O��1��ޜ����Dh�G�o�w���|�>!;�zC�a������_�܁���N$��M��k�c��W���zO)��&�|���ݼ'�{M�:P>�;~t��;xM���
���b�ܶ�W��ҷ����> ��)������/�B=>�����ÿ8���������=&v���4����/�U
>��f�O���<.��z��q�!�O�ʞ����jl:{�#���_����w�~��g�j��(�O�.��I�;�^N�S���P!?]�;����˾�U����zL.��}?y�oϗ.��s߭�(�o�}�~��*��G�GW�����6V���|�����#H�!�����{q�<!�w��nWI�ۏ~{��a����'� }I�q�����́��c����?�~��&eO���s�����\G1|:�t�h�������ז��>'�>+��U�����n���v���m:�,h�%�}�~k$�GT}�����/�-�*3�hո��Mwʂr����-��rd�a�=�(�1�M��{ �y�ޱw��VW�we鶜t-��X���!o��� $��OU��3�!ɹ��0���G&�xm��uet��2Ѳ�����l,�NWsܜ������K8�u�����x+��R<N����2/{�2�\����a��2k�A���}�厡�zP�7Z:�N����Gz����y�kS7�;jtF��`3P4&�R�Ǚ�/�?!�:� )�`�驛ɝ�I&c���p�a���{L�l�q��Yϩ����k���\g�7�7��*��x�Ҿ���MEZ3���BjF���G���]얮}���kδH��ki����r��1+͠�|_�� b�% ^�}�u+lq�pECe�e�t�cZ\�7<.6�;96ov��i�iU����N�B��~J���5.Xt�#��"�-h���}��9�&�zj{�W�k��.������Q��C�I��^L�
R�5(�� ����0i�8-���N��
f�gh���q��O���HXy�G�t7uCxŒx�="ℑ�3��b�*f^���������1��u���U]BI�q��~rz��P��u�c�#�ޫT���7.%=���1W}�r�X���f�x���A�a��O�2#��������fCs��Z��-�x�SH��I�ث2�E�(�\�2��SW!v�R��]�N�X��]}m��m�ޭC���*lѾ<ߨ.kwU�T3β��p��%V�.�U��vVb첝����Z�0J��;a�)n��Is��3�g1Rc��Ó�}��|�/:��L���-�7nfϴ�wl��`�������@�0ƚ��;����5�:�6xQ�ݛm��}<�V�'0�l��ڭ`ėx���]���͚����/���{�FB��ɞ__b��z*V���b�i���\����cڞ�*��b��Nv��{^U>6U ��Y5�9L�ߞ_�uÞ�p�:��Z=�
:xC�l?NZ���;y�bføwT�b�QX�|�4�`�`2��[<�v��:rcD�V56�m��W[܂�B��A`�,!�ڮ�g/��7Jb���;c�p�Ȃ�Gr���)�*
�j�w���L�<~a�O��p�]�6lsbE��_?��,�-���C�nwG-y����1�M���8�U*P��x�}�8IjJԬ#���*��ï��Yj�Gf8��Oq^+ؗ9�.
�|wa:�Ľ0E��%)j:���PRV�'������=}�f�ʆU��p'��Q��|���g$[����6؃ē��H�"^����9M]`��6���ד'k�Y�w�8���[�+*���V��ʥ+d�ed�.�U�,�M���k��|y�fgM�y�5:�j�\1��w(��{]�,n��HZXԢ�;k3�.�߱;��)v�EԊv.-�,��ɝ��.�;����M��1]��Y�>����l�p����h�݁ҙ��O˩�h�/��~�`*��$ r���y��|(#�U�U;�*ЅN;f���Zn5:���<*LW�ӳFṈ�U�1���/jX�o+�=Qd(���'΅����i�핃/Y|pxc��>�;�#�P��'cG���/S��l@"^�^?�L_�@�\O�U�>0��+���(C��u����;���6(u��X��M�ɝֺ�c��t�^�hS����1�o�kc�lu�g���%wO3�S�i��l��W�<�y>�}Ҙw�X^��7C\+&R�hL1o��0�����^�{�`�٘�橁Ъ�,�1mW��ӚhC�.�@�ji�Sd��S�u�$#gK�^��u�9O�?G�[�����P�e��S��d��3z��� 	��g[���VD>����N��7E=P٩,EN���������*�:B'{�qډ[�-Xʩ7Up�{sE>�a k��m�D����>�oյ\�x-Y����vA�{��y-X��!1�r��`���X�r#�l\z��D�R��f����cx�]�"��Yvh�'Z]%"#yY��ha#��)�h�^���c�����ݢ��x���l�����n��ܙ���b�r�[o�+۸��֝��>i=��S�7���W.b+���gg}�f9g'=&N��'�GIUc��{t�Z�P�36����Dx�qA�}�A������)eܳ�f�2W7�0Y:�Pښ<3�U�Un���v��Fqo�>�;�O��~X�!�c��@�V�E�4�ҙ}��e���z*��
 ���:~L�(F|�5���dJvٌ�oJE�7��D�jcPZ�UkS{�]֎eIY.Oξ$LI��B��Un#,;/��Q˭�0���$'ja���%���mP�K>��C_�ɠ9����}���(5�ɪ�\b���֮CL�r򣓴���]���Z��N 9`k���N`����@��e[�K���"�E3CDӎb�n����X�i�7v��MUѸ�Rr�����;?	�����?-#��vїO�9=%����x����qԦ4TneB��N�� :����;����r��
�
G~�l/^Ёҏ;�yۖ�Us>z0�k&z ĩ3�#�o��ɇ�N��\���k4ҕ��3�X�rm��5��0h߶>�ow�4O v�������X��j�O,]�x8���/ɶ~X9A��kƻq=�û�A�&5K��^�,�;�0 {�9�s�2�]N�y���-$����(�!~��N��]R�?\�yThn�Ԗؼ��<`mml��W�W�XnG����b�c��ص!���q��7���k��e�T&����c!Өb-��;.{���v�2jf�.1;]11F�=®�ѕח^��j�cb*U ��`M�̊�/*��gwt����b������0k�;L�0��}Я�Gs���t��.ī�=X��-fM����S���Ċ�)��u�Z|�xf�-�йp�wŕ���@�Z��[Ҩ;���[�'\�J�qt����o*0�*c�&�G\d��ON$���I�ΈLs�[����Z��_ئ0ّ9�[��2�柕������vZP����c"����[�r��'��_�>�ާ"�F�����D�ֻH�G9W�6x�w73�\�%�Ε�����*K5�@�H"�66g��Ч�W؝pё-���clH��w2��r���\N����+�߬=V_��D\	2��=���8=�j5%Q�̃���Y�!�.��uA8��U��[�L_�ņM58�A���^�R֋m}K�J�|���vE�j��6,wx� ������.*�C�3u����H�%����=����-�B�ÈQ���7��$�(��rE����r9�y���;Xz|��!Q �n�>�EZ�{�+l69��Sg��z�^�&�m}�|�D�}�G�}x��Qk8�{����f/a*�%7<A� h�l	�T��t�~Ϭ_x<gMkC�U�4^4����}�5��Y���7Ҹ�ܟ_�ک���M�7@swT7�Y$���kLo0MGgn��R�V)��<�p�+l�w���U]Bߒwh�>����{T'od�>�U��ʢ��WN}�'־�-��X�	�Н�c�����&;��A��\s��P����g�s{���3{p[���|/�U�{�ՙ��̅}��7f�|��a�aP��Å/g@[�\x�y5VLXhΝfq��bᩡ�sr~��wR	���6herT=���Z�!�ry��/f��n����q� ����
��|�s�%q�Ǧ�[C)D�9`71V�:�:z�w+�1��+�T�'A�T�$n6] ��Yd�s��퇗�p�6j��/(�8��a:��$x�s8����k�Na/��|�̊u}��.�!�ʳ�7-�����[�.	���SYN{4y�iB
:}O��%¸l�U3�}�Q�bA�N����p�DdK����=�d��M��p3��J�[p7ޤW {��w|�=��J��yl%v����._>�5�Z�jqo8st;�Nn�!Y�^�x��N���]b�������WIә�;�B��#'+��c��^�ڇ�m.�1q|��Yj�����4�/��/.��^�ōMWE�}����{�c��-V����|�m��mb�-�ܻ��oo�g��F��[�`G��D�6��pnM�>G�'���kϮ����%�F�]��Q�CjdU��yJݦ��BV�)s6��"���s[4*�w��d��Q�%�V�u��X�%���s[�����R{��0� �l��3$�J�o�c]x�����=ەj�ݧf��y��BV4iJT�[�"���Ѳ�aG	�gCbm�/e��[�Ƈ��M��vkX�+7ka�k%o#Z��
�7�SS��VfwKZc�/O��4�U��?F/�C������b�ͧ�ȬGY{�m:c���w�)��*!h�C��璺.�����2A��ٳV��X��wY!�[�t�P���4.�;B�j+K�~[O)ĵ;Mm\Y9��C�n��H�����S�1���J��,��1���F� �>c��N���yQ��mj�Suo�lM��P�L���Ä_l'z]>�Vv�'I�����Em˓4���2���%;�_�+B"+T���O���k��<�Y���>��ׯQ��ť{�8�7.�Z,-4m��g�VAf3�M�f��\&ur�#��NƵ���l�k��@--8��j�b������me�E�[��:Tv�v��Ƹp�y��׆�^k"���TwY���ӕ8Nb<P�a��Z/�	z9�Vq)Z��g�ؠ� �/)�9��� �2�<�NYҨ���\�}D
qImu�V�}9�x�e;�������hZ�jP<DRRh����$��5-��!�.�P���'����&
$���g9��4fA�S�f�����Q����w/����u�̼i��G%ٖԻt�h�c���7��̲[���҄�,��b�Y#�ہ�s̩mŁ\��$b=�[%:�:��yMd����LX� ��>����,k]��AZ5�P{�[��Ugw-�>��Ը;7afի����T6�v�@�"՗����(� �/;+�WK���\a���0��1Y�ǟk<4�n%7Wbh�������g{�e�B�Z}�Z��xHȮУfRU�]Ȟ�sfǤu#v��
°/���Q`�Zi4Yީ�a@�Y�M��%���ӄ\�����y��<]�0���[[r�og=�KWs�\��\(� ˍ<�K�0��b%��X�]�7B"�.kΫ:jlŔRBrXc)�pvk������t���1
b5;�X8�v��/;/��VJj{�xHF�wӮ�����0�Gm�L��K�p�;oU�����}y}Ң��
ÙbI�(**�6D����]P��*��Э�j���ST�TeZ���s�=ݫ��2��I..�faւa#3���2�[�2��%1�b��R��Y-	%�t9m3
�R$Ԭ�$,(�fZ��CNY"�R�.ua�A"Qa������)�gB��Z�r1C0���HJ���Z\��H��l�� �HL$.-�Tԉ(�Z�&�w<�2��tڅAQl�&X�DVbUer.��2ЍL�9j��Z�`�%
����	B6���X��2�4�Bՠa(�UQ�u9��S�j�2)$��w��6TQGMD��uI��ᡋ-52Cj�j�Ez�Z�tE�)�j(Z�Rґ2�B�-"�,����f���*LTLؚe�Y�c��z�F�b(��֩�e"t�J��0�B$�Q�	�V&Z�DE����i���)���_��|β`���;̝�7nK��r7öY���@�6Dw�.�c�'e�\2p�Ll��w7iM�T�����W�}T3�R2۔� U�Tn�H��P�'��`�2/�a#����ܨ������Ӯd�z�]}#����cI���8T%J͵��4�%�%jV��ͥ7}�<���_&l]Ѯ���>5����p��΄�of�uHM)���F@c�Fo�R�2��]�M�p.4�e��'��X��ԓ��As�9r�j�����3 ��\`�kx*���G��� 0��%q�������c*9u�)��(.m���Q�]2�^u��^��c��X�A���]�C]�����{L\oJ�q�Hv�I��杝:Sr��iq=<R�k}��UL8�'����@�uo�V�?i����U��ar{��V���r��&7����f�Y��t���A�:Pl|�g� �κ�1+øj\�z[�&��w�*Bud�ULE���f�!�@p��z4)��m�0o��UƷ�i|�>qP�S���q��6k��0�X�R9����C�3i�����r��^��Ln�W��Y; �KHi�Q�k�+
���<�e��!Y�"���\�HoD����cp���D�d�&f]��dxC�j�E�6�>u�\��ع`��ܾrc�p��OnVc(�ŒA�Q��s�X��yz��V
涪羓ziB�uX���Wu�������]��w�Q�å'ra�i{��Ī��t���,��P�v�W�_Ni�����r�ql��W�ק�*��I�{�[	}ؗ3�jU�>ٖ�G3̠]:l��nI���x*f�8K��������8j C��)��4��S�F)���3O��x�v��l��5jZ�Gf�Gl�=��Xf���F��~L�҅��t�ȳc�#p�n]]U�S[ϥn���+ё�&ˌt�N�zL�������_z�]��J�Nq�]7O��z���&V�T>����gc��co�ta��hg%�PD�� {T���ӽz�Ujm�s���!�1���V7�}I����;��\��"�#^:�{iQ�|
x��uM� ��"At�"�R��}�S(F@Cx�.��Jvٌ��ґ�s1���\;}��l��ቹWQ:����$�"Oˢ�s顟u��7!a����k�]l!s����a�{�G�H_�K���ɮq-��}e�!A�?5Unr~ި~�0�f}5=]mL�)�%(�^%���_�=�6������v��ʄ������*��zWeӲ�14�J�����y�9��T�r��!�������,�����vND��hD� �7����T뼯�vm��m���
�
\y	v���h��T�6�w������e���0~�;G�J�/ 9`k��d'0DO�x�`��g�}n��v8u�9�ڵ]�6�h�6\f�1�S�j��c !�Br���eX���'��� ������S�B�o��d-L�:��ټ�g*1ʤ�a�k�����=WA����Ĥnma�5&ړ;|�R���._u|f�������L�ӯ�0���3���hJ�5��E�ܢ\:���=�l���5n�ׇ/��)7p�>GG��W���Ʋ�N����C&%M����Jww����$r�����{��]�vN������ՓZw�Ta��=�N���ongz��e{���^~�������82�-�,q>�+���x�3�Qή�,Tܾ�Cǋ2�ν�;Z=v>�)�+�r���,F�:���mL�˔I�Q'��6�E�O�MT��<����SN��iUG(����?0��Cf:��J<>�a5�)�-��F3~��^*�w8W`�Ne���t�1q�`3P4&�ԭ��r�q��K6��U�LW�&@j��z�����J|&��z����u�\����4&Cw�=���>3��+� �j������j�	p�)����D_��A�����z?3��VE�9X[�b�9���A�:��q���V��4|c0����9�[tD0���������v���@���@B~%#���#���fR����x`�z�p}������5&qཱི|_@.���"�W1�5pD��6BjC	�r���E:��т�Ƃow�����]���[]5�{,nCu�M��q:`��1ux�dR��WR��8��5�������6������I�\��j�ϋt��"�%�`uuD�C��DJ.熑���u��=}�l7���|z���-h�bSJjt��E�`O��"�j�~���������[݁�g����!��{zW���mLH�̚7	����*r2(S�S���n�n��+I>j��f֊cD�=���l�wO+�mS�ww�`��L��$�nvP		��c�ӝ;y������Шo�4!�e�2���ҹ!`n�~����/=��w���-Ml��>��K��~߯�o��2��9���ʁ�5ғu�7
:N����r�*�����Z3�3q։\W�qW�{�^����_)�ГTKv�bb����!�>�8��oZ��7΀�-|���_���*X���m�|��-��)�gi��X�⹂��}�w���3��f�nbw�*ԀMH��{t�|E�D�����������Ɠ9�w+��gk�07���PyKQ|%��0Oy�׳v{z�ѥqfZ���sݻ_���|�'U����ء�gY+>�b���1\��3���R���VÃ*b�i���Z�K���*�{��x3e��f��Q�Ν#3��h�l�_Ĳɨ�)����c��ݸu)Fͬޡ�t��Z�J�4�M{�py�KJ�����y�O��?�C�A`2��r�Q;vV˽�Ʉ��:��}Y�k1HΝx�$�(	�X���n��<W@�w������H;xC�K{Dt��@gi�p��?P�82Og�Ps�L$z1]Au��\�T��#��u��V$?�'FK)�3�sX���V(�M�x�}�y8Ie*�jz�0L�!�';���K��G����Tc}q7��.��݄�q�D_�௒<��@�Fx��R�4��(nh|�u0n���?g���t���D6s�9XS�l)�MOβ���[3��{�I�\��ɀ����F��L��b�9u�)��"��/o1���k���T�7=�?�k�dV?&�K�8�Ś7j��>�<&L�v��#"��;MHs<����%���P_�$�w�X�}u
�߬m����+[�Լ��p�+�Vr��oV�~2�`��X��h
�o�ncr��JYY�SI\P<�bJ��\��mwB�O�^�z�Cb������q������ewb�}��/�� >	e���m`�F���b5_ʬ.��|Q=P2~�ي��]q�>�T��nL4[�:3�{;��5�wB�����0|������-Wl�,����;��ONP4Z�_�{m\B�o��nׄ�y�
���<^�y��AVz4)��m�0o�^��w�:[�\I[���Ɲ?*�h�A����q�}l@�s��ں�������_F>gfęq>I4T�a�|L��uX�T�Ɇ���<o���j���,�1��W���yY7`��<����9��u��b�Õg�ٟQѵ*�S���i�b+��)�Nk�ŕ��M�4��ֶ3&�pi�;w��Y��b�+���+>s����=��= ����$�999�Xq�LE�	�g��u��3|b�vT�Y�az|�}Pح����[#���1`�����G��o�ݺ����|�YHe�����M����x�I@�2�����o�kU��y�ǓӀ[S�=wpY����*xs�r��t�oz�l������Vc��{P�노�鍯�_';����OU��\���X�Q9��B-T\>�ң��۴"�̰'u���O�}i��Yϓ�)e�Wǃ���Ϸ�͉#�{��Y�{j����-�+�qE���tC00wg���h��۝�� ���Pn�}��0�j}%�=1�+L6U��")5q7,wL1�S F�x�FU�p�F���ҫ������?��Q��rW�2�B2�O��ޔ�SMIX��nn)ys�oU���5�ɭ���=�}E���D$wژ�9׆]q^����3�{6H�L;f�'��@�K��r�5�%�c��kO�Pqv�f�Oc�t`��!�Ӎ�����c��\�/�z���2^@r��?P�N`��(��d-6^Tep�T�E�<RX5*���(�.#v��Om���WF�2��4�YV(;?	�d�e��N��)�v�@Կ{�����h�<d
�������Q�8!_'w�s�t��~�S#�֘��CFq#�_<��`s3��ԿP9딇���G���gx���{2���:�e�X;*�G/"�(���w:=�w�֚������k��͎�����<9q�H
�q��.��YuP芌EU��&N`m+�V,^w�ۊ�k���c�n�&!d}�yW�=NQ?��4��(���g^nc�f:��:� �{�x�����ya��񦹨k��%��5��f�,A�87Y�*s'p����ڧC�⛕1h�V'i�@D�5���;�����(5�t�˜���w�BS���K���ttV���<=�S���G�HG�ջs�8������,�T�f����z�֢MY��I:!e8�6��zld���u{#����WT>��!ŹM�o����y��۪V��i����o�������k�ռ�,��:櫑�t |]�I]��Ã�:�ۆ�_Ε1�M֎��v���{6�m�a^"a���%��,	�.�wt�1q�5�lК�R��9�e���>�v��n�I�=��|�����Q3� 0/h���!�|T�+��-Uk2��{���v\TIƮ##��U�\n��)z�3�W�aT*J5�t{��"�R45��=is�U�\�/k{w��8��Xw���;�������`������&J�A�����վ5r�tP�߹�gy'�3�vת
���pF����2t��"�%�`uuD�C��G�+�u.ꎁ���\�Y��� �J���G��|��Z5p�C�I��}? 0p`]s|�*=�ۧ�����%N���"I��"��?I{X*�49�{Ҹ�{_t6�$W�'�4nt9�R�G�i�p�����e��u�W:�q%��/]q��@�m�)C��]�X�[��)'_'�ЂU�I𲫻^��!�P:�;R�� �:L2{�ޢ��#��A�_�gW�ٸ'��C-Mv�N了��&�Y�����������qj�{�Y �*�Y&ra�#��
���q��جه��^\$�Wє�=�:�?>�=�u��G�[����7��U����Wl
�q5�0]=��a��FL��u{�Ϋ��P�òwn.t�,�]|6�*���-��p��{,$+�ey��%y����7ܺ���<�޾ Tn*�-gQ��W|���twV��/�n�8���ŖF�Fl�l4�g�}[]=oX��m�J 0��O$b��ɸs�-���p��X�pW�0��Μ�1>�u�`@K �������b7��d�ɮr�|�cS��b�@3!&2���EVB��ND�D���Ҳ7�S�dS���q�����R��um��;ŭ�V2I�)ҟ{�_�����*�@㢸�pu��~7U6���k~���Ft��ܝ5�y���J���m&�a�g�#�I�2����s"��H�ye����;]�)r�ZƷ�����.T����h�|�N����.U�"<k�m�W jE�{�o�;OnՓ%�%�uF�ᴂچ��6���d�%�"�2�b�M�G��*���W'�,e�Q����؀�[�x��;��C4�w6i�1}�03kzv<є3�.y�ǉ��Fk�A�{&�� w���]�n ����==s���^O7�ՙd�W��>����"*�����7u���f@u�O�'���]���p�m�����<�tܒ���߮�\��h��ޭ��q{�'��Q��ܜ�Qs�9r���@���4w�Wu����2I*˃S���� 6xEuJ�tt�n4�1�˭�L�c���6���G�&ywk���>�����V&�}g���..�4o9��}L�㔞�W<
�U�$�q�&LV��E�s�M����5�OP��jv`�J���1�h'C=R���72S~�ܘ�9�]���n�2�BC�8��q]HK8R҂C�Aȸ���b�X�/��K���Bdw[,ed��e�X�#Z�E���f$k��Q9��ޣE��&��"ݢ�G\�ZG"Lh��3�[L0C�3i���j�'/��z,����5���"��b�/��W��;fr�N��2Q϶f"~�j���,��|l� �S����k-<�h��w�U�t+a����q.D����C��k��+��iC�PK��M8p�9s����Bz��nV_%mUl�L`�Ҕb��W��b�'��*�R49�ec�-倎]�<GU�4�e3pU�͠@.J��cfí|�zC�jĕ�v%I8_]�h��`��8=�>���.�ed4���CHp<�-wX��S+��"U����hn ����lK&h�u�]z3���-�G�,vY��*9�~�C[oX��{�5̲��v<q;�ȋ`;Ǉ��;T����׸Ɖ���ݣF�f�A��v��C%6+'ǭtY���`�U��#f�G}R��d��	u��Ѯ������Ǖ��qtQ��́�|�*]U���`��lݼ|�
�5�Aj�лv�,Ȝ��y�n��g�����0�;��7���e�)p�Lt������M[3r��!��sP�t�[��B/m�{S�m�{�[:8�}�ʺՠl��/�d����(m��K1-x{�j�m�3y"#ojTmI�f��!�8��a%��������ܴ�|�[t,��d����4����j���5_��ҟ���!c��Uk���X�+&ΡY���{)�{��qJ�GwJ��:%*	�$
G��Qd�m""��:]����ʅ�ۏ�iY�����0%�d�V�v3�m�.�ԁ�L��l�����ՙ�D�q�Q����,{d����;V+��s����+���O=�����9c<o�B9j`�=0�/�ᢔP�A��4x�F6�*��y&hDqd�H��@m���t�8���G�5�W&-�%����t������p����8��Eu��q�#��;�����og^	�n�p"mGp�7r�;�%��e����2�=��3p_5:�u��5rx�ӵg�شq�Rh�y�_�ݥ���̫%j^S�i�4z뉕���C��R�/hs#ψ{����8��Vܒ���q~{�tX��'P}��7��w����p�wAl�:���xy>�-��,���]L��o%v�Х��$���KB��ծ54�_V�((hU��[�_&�Eׅ)y,i"q��%(6-ϯ�uF����:�Ւ�{!b�8g��}6�f�3����7Ì1aƝ�YP�qv�Q��
���_9��C����kŵ���q�MUG>75���)���S�W:�[�A'<�=+�sg(�����ޞ��mv��s*\���M$�y��}u�"l�<�z���:��no���=��vz)8���Z��u���DtbO��M>63��'�S�B�ӻs�	��I��罯� �n2�%���Tmրv6r^sv��Ը>����&.����鎯X}���1椨����@4���09Z�#޵:��1��yk�gY����]j�1c�{��k��O.�������z=e�UI!BI��4�C�P���T��b/��r�##--N������E���U*�K�XV%DRs� �@����V"��%q$B�%0����Ф��2H43:�d	�!,��&,Ф�6YmA6�Y���q�Q
	E�'���׋��bQ��Sh(hF��3��r��OZ�U���"L��l2��Vr���1BE�fZ�Ee���\"�P�rr�"�30�����J0�,K2,EB�LK(B��#���g���H�7d�;�F����m2���\ ���N�h{��JB�5�GK���;��*n���x�(˕a*�z�ˮtt驙�ab��*���+4M$,R�w'R���Y��s��&&�@"�wwr���xOk���fJ��r8��J�!�l��:�4��z�;��Ĉ�{������G�l#�&��)���G�$`Wvk�1ĸ(gw
:��N`ۣ����5ȷs<=T�i�����n@e(��������lڀ��K���ms]�*�3c�CF++��8l���|��b\nbv�R�������?��P�n[<�x>��R�Ř6Oə�=Ho5e�fRy7x�-�6k�eٱ����-��w�\B�:ju󳩬GK�<I����vY��:��V����(
WZ��U��Qz~�)S�̆c�����HۅU���S�f`㻗��inw!���7e�Ibb�b(BE/%Y�YS�a��`|������Tv��g\���g'*�G8�f�d�G.H)O�cL�P��ы��d�m�軉)Ȼ���n㓹U�x�Gq}�la�}A�����R2צh��>�j��ϑ�QWuҡڱ�˳V�G��v�!�[VY�b�*�u�"�@��'(��]�i�8<��Yhvg��[�5��c3LSަƵr�z���S%�,y_X)����2���K5�T�jL�u�LU�3|¦r��ok�����jj�����',/!eX���;�gΔ�v,Z��������(	H#$�5��ڵ�l%tvk�K��� ��վ`�+�s^����<q?:���&���b]�����'�O(���>�}�&���1f��J��
I���G��$b�v��$�E����UWOy���Y�~��x��� > 2�JM��֠��͍����@��-�)���-�N�.t�96��=�c���
�v��L�rҸkhF&:�O�,^}]K��wJf�m�Șx:�WV�^��y��vޅ��X���f�G=��5��&�WT0vRn��#��ܽ|��]��y�⾻��n'P{�����9~�6�ךi����~s)1�r��jߪ7B�̹{=OV�'�{@hq�~��3!Ru�R��ooɎ!�Mn0H�=��������9����xT���Y�ݏ�6H�)��t�qs�������FZ�y�A|��\�]��I4�E�{^և57�	�Į�dqt����k�{pً�����ܕ�L-h�bJK��/}`�Z8w&x	���_]!^)��6dN}�[��C/�B�uV)H;ƈW��u���W���*��ty���w���~���缡���Z��k{ZK������h�9z�3�TC�B9�h�m7]2��Dķܲ���kq�[�{��S�� ��I���Jv�^1\R�:J%-`�]k����[���٥�۴������/�sx5L�jp,ڥ�':�<� ����+��I����!���(6Ֆ��wۚ4廽~d�Zxn�&[��LǣC���l˭�����ԟ�  �יt��}��F�O�m_�����w%��A���聋�&L�/R�(���oQ���w8���xv_����D`I�pq�Dų-!Z��C��91|�إ:Û!dqv��]��pzH����\�z�#��ƴf/a*�&�7\��E�6�x�TspSڗ\�4W�+'�@��~���p��8�͕��>���Q"�O2h�ʎ�ѕ�HF/�[3�����ꬹ��P��WL��N����p�1��x��^t�\|y����qr[�3'��+՚��;+��Y<�
���"��X�k�`��������"�iG,0�e7���FHO�4_*}���!#]|6�*�
�8n4�wA��9�Js�?���-e-lٍ��K/�V��a�FY�e9�a|���9��ۺ�|Q9���Q�������x�Lm�w+�91���<�� ��Hϕ�6M���JtGvN�a^j4v�m�;��rzL?��P�Ie�Ec��ͳ��U{���B||MG9L�ߞ_�vDG8�`��n�?L̀3�ٹ&O.$���Y�O�N�J���\	�%�oQB
�2t��-��b���.��2�U��=�7�:ޭ^�mx��Djƀ%���ː��ݎuղ�Rs �0���.��S�K�e�6A޸�lW�|�[�u|Y~�#��oh��k��B){��ٹ8)L��	�
����S\������^,�+k�+�}.�}�;�����xr������i�GK|�8���p�����#�k���F<Nl�پ�Հ��3��׮!���rj��|f���P��ĝ�*w�UY��3K�c��ym��H�	�z���n�8��YW�+<����V�z�`��>��>���L�cCU���:� 8-P ��� *��b}q7��.���N�q6�`��T�������G{B9.0���}PZ�����`O�Ɨu}��EAs�,��4��1 e\��a�7E��O�^p����%x�?��& !~<"��WS.4�1�˭���#%��I����f}8�0����H옜m� �6;����@���sVͭ�z~�j�f�ȼ8&L8䝚-��jh��D�(�^��_Z�:���>do�@�X|S���,o�;���������<"���z|�,�+>~�tʯc�|1	�iC�~�i]�k�Tz)�7�I�>IG�+��n�G����"�Nޕ�K֞f}�0�~c�D,Y�c��R���:��X�'�H��/|
?b�}~���v���tgc�(��1��j뜷2�+��S\:fN�<oI5;�������9j$�r��qv]Q����|>�;Ym����񝧇>W(B��cE���/��T�\B�A��Q`�f$N��ܸ��yMYQc�X����R&�j;�}β�Y�CH�@g9�ݮ���l�S9	�����p
��ى�7�wb�;8~�TDu���L�г�c����4�ģ��o��[Re��P]�}�2R�fF�-M��O�	��U}�o�F,8�+Xn�[�kRӢ���x5��_l������[�y���Md��V�}�U�f��������Gݡ8n�z��G&��)h�zZ~���{6_9��Xz�[�HE�-��w\�7�+��R�4|��Хy���`e��H����q��֬��K�&_}zs~C��������M`�d�q�X�õ�9��s������@�ۦ���U�n(�?T��Ȏr����M��z�m�4*�˱�و���Tqq�����<$ϝ�j1��BE/�*��s�A���.�1�`L�n�z���g)Ng;����^Kg98��F�!��<����a�_
�)�#�O�L��$�i�b�R��̝�J}v��:�5��=���2��X�l�f�����d��a�4����,.� a�"�F�U�����{JU��jo"<)Ը-B3@=��i|�AY+�W��szA�)�(�+�����Y=4ZU=����[�U��%��{�f��Ǉ�=���U>3~�,�ڳ&��r�����uLȥ2R�E���1F�S�l�^��۷ײ�j*�9ʹ�F���iu��Ֆs�Eĥ���z9L����lw��B�룦�E�A��f�T$t�W<�UƺA޵r�g���K%�偮~��'0DON�w,*�I",B�.����,�TT�[�6�ٽۄ"�=�3��]�c  �`a}�ʱβ�íPV�j��F��ԣ`��h�>lZq3�@������w�lB�����B�@:S��6T�J�H��v��}��m!�=i\�ׅx#�-}�0�Z;7�/���5��}�+,[~JdS��Y�}&���<Mi�c~�Fŭ1!y�!����U�����-}$�=t+��ָ$��Yc�P�\K�Gq����[�+T�B ���ԁ��Sa����3��^�湁�W�k�U5�fF+N�鳹J��7'Ef�N���1D�β�\q����Y��Mʅ(T�ސ�.�}q[$[)��銆��/�Ͻ-���r��7.D�����W��68����C�>`�zzK��ϼQ �xRw#��2ֱ���K�h�ʦK�١�0�񱺌�����Ӊ���@w��wNr��Kŧ���z�K׃��Fs*�Bm\������s_!��99#��(l�/;���}��g�(�&�Y;r+�s��jO3A9^����C��T;O�b�j��e����+!��E%R_v�}YX5��=~*��)-��%����p��d`��6hM}�[�!����Cd��]��9������u�M���x� ���q�g"4�G�UZ�:2p�'����Z�W�ã��]�v9������!
�%��uAtDɅ��.M�Ž=���|�a�ӎO��n�hȖ��lޔ7>N���z�'M�g�F=@�� �]�q��qL��iH�)℧,�s�N��<��W��I5hgźDų5NQ
���;���yq.p��JT��E��z�Qh�oW�8֍F%0��Bn��@t�(ٶ7�J�Fc1p5�SZܮ�WI���d�?4z~�+kY���ޕǓ���mTHxs��݃�1|����v�4_ݮ��]z�MBJ�\u3k��u����wS�a�=��y8��G)�]��r�p�]���'�̉�7'�J�8oL �Н���W�c�Xk���gXT�f���w��t���!�&vx<l���x#�M�n͟���On��=v���E���=�p`܄�t �蝍T�k���9�pK]��P��K�����N���%�d��-{�Kٻ�1f]�a�nm��en�@h��C��D}���[�.V�>}�]�Lz7�l����:}������V(Tsʜ7Q;�g���.o����CyDK�m��1O骆�:�R -�Pţ,�3��s0ё�wr~�wR.5�Yr�����
��&7�W�ue7�۟%3��,_4�F+�l�~���Үv�WZdlS�1�)�9~��`�� �F�9���[��u�ѿ�] �>%�O2�{�T�Z�p��P�[��A?���ݸ����|I5��%��F��J{̊w�#N�Y-ͼ
�/E�ך��]p. �^�9l��ۿ�D��D���~���{���Rܭ4P��נ���.��u�G%l}���8[_&��kE\���uq��E�wv���|;5�����u-颓�vֽ���)P��:�������Z&$�K��'�>f�Kk!gtb|j}��v�S���q+뎦��LZ�Fe-�J���,������J�ͥ�-�����z<�R,C�۳^�ϝ�\�e�7ᆷ������#: Ī��5��O,�d�U)�F���\���'?FbjN+���7�P�����x̓F�ۺ��y�Fh�9��y=FҖ��)����X�"v�܄y��w{A˴���9[�n���1{~�ﾈ���q�ʷ�m�X+7#�u�(��R��'�}K�r rx��h�]Nx�T��5�Ԓ���p��\"�o_P;�Cb��y:S�������]ݺڱ�i�y�]B}SQ�Q�~?q�������W#���ơ-�y��\�w^b��	:�X�M&���m����~��+~k�
�,������_Y�Թ�w=��+"�c�:�헾9�p�^瞷�%#�/�}�`�'j`Zu1Q�}q+FTFru�\�/����7]d�VTKTS����'���3+��`{79�'�;��i��bm���_���'~Z��w�CϏ�[S֖��V��ﵚ����x�?TO��eftMvqO�n�诹&�Ķ��&k�/Bο9C�X}k���O.���3k�U�=.s�U�T�0�*�5���!�>�5��{"�� W+�B�V%�`�c��ty��b�\Sm:� wΎ�J@׊�v6�J^L��s�@>�8�;�%p"���C!�U�h��*P�ҝ0Z�̊b�S��Y�)�~����X&�zr���𻏌�G�k���yT�5*��g�}U_DF��m�u��uWҥ=A�JT���+��F��������\�@�vk�0�l+Co@�W��6RJ1Pu-騂��p�,p�X��ٙ���Y�n挖��t���{B�LG|�J!&+�),S�ҟ/�o��=�"�{����z�ڻ�RR���Ôg�Bﻲ �`���Қ̀���r��Q�)-q5���}Ư��*�f
�����2�]_	J�h�Lf�
N7�q.w�L��3��ת��o��9����;��p�
�b~�6=�f7iF��n�6wkr����}6���x��	��i��´䇱��LK�B�+�N޻�NߎP�H����)����z!c�5��qY0�ؽ�A�u]�[�������"򓾣ΎŞJ|����r�_']���UR:�pd���`�k�[��ؕg��������w��K�[��}�U^�v�f�H}��a�����mB�������*7���(;�٬7��NܨM�F{��7�tC�j�\��N�m�{BvDc*��#���h�2E��(;[��u��%��3okh_T	���Y"�;˕E̤�ᗬ#rk\�~�S�v��jY��[I�o�ܑe�6����`�u�Qf]��I���K��v�ڷ��u!d�Β��Jܱ7v�C�}��So��r�ő���fF�$n��4+y:9���Cw�A�JಐwuO�g�0-r^��D�Y}��Βbc���������m7Z�>�i�њ�4%�`YH��vd�.q�ʷ�c�Aj=w"��B�[�sNz`SGX������~c��fNU_N+�&=�.�:��M�F�
S���$�=�TM�E�s=���q��7��p3�̘x�����7!���������!-s�)��#n���h������!�)���c�b/���xG"�QP�X�%�\C�Ǥ�)������(�'n�h�����ה��l�w������)�VK���\��n��|��\+U�s6Tam����0�~GZ��k6����I����7׹�)%ci\���Q���,V�K�X-l�.=�Q�����Ү��aƕ��Xw��d����&`}��ޥ���*&!%
�Ȭ.IQ7%_23�ȓ�*lk��_3t{&E�P�s$@�v�mu}��n��,�e'W3\�q�q:����3r��Y�#Ҍ�Ao��·B��FIQ�_�XyZ-6Q]�v��q�b4�Ђ���yp4Fk+3s_>I��n���c���u.6ٝذ�cVo9]��5ip*���i���Jd5�v��uyjC������,n+p��/"�����
����L[�����T2��z`��1⺁��g��8�Td�;��	|s_��R/<#٨��Ѯ�6vY凶�9�r2�Iٰ�PqZ�CV�|eZ��io�%��^�hx��Hˊ�&��)@��6-��XWiOA��{<���1u�HW�.��1Uop�^��v�^�H��n�z,>O��B#��f�rK�C[�vs�1�ŕDDpo�ܯ)��q�b��}�H�H����y�^xOM�ĝW.��n.-u�J�%�kC��,���v�]�x!VNix�y%�w{�"�x+:Z�T��m��-��t�35>]Z���w�=�`��D��S���v�L��ƓnV"GL�V�]2ҽ�5 �M�r��I�����f0�9�B������oZ���wŁ�k��+n���[u��,�O*�Ҙ�j�N��9��5$N�*ѽ����-�;^����o��v�$�F��"YIXbڶ�����Y�<�Ⱃ8������R;(��/�k�t���?�B����;�nƎz-�3�NDhG&/)�7�6�Eϖ�=�{�o�Xk9C8ۓ��oK�s�Vb{�ȫ�gMY�s�B�Qe���M��a��}��We�pY6>���U��a��3$n++���=D	�����ʋ�b%�,�+P9��v�2��U�k�SK��br�5N���&FWU�B�Y�T\���5"+"��;����+x�[��t�{�],,���*-���a�ZZF"�"I6�|3̺Ta�(��IHZ�L"9HZa��dWB���QeAfr��"PB,�,�ҩ�U�I�[��mH�н�m!#P�cB�MVK)g9fȪ���0Ԣ����EJ�BQ�f�Q��QrN����A���I*�l�8�
�Xe��{�{"�,Hº�'\s4QDMgsWr�:�t<P��-�g�rr��(40�AVTr���u!�":nai�wZ$�s��"u�H,�"Q֎�w*Ւ�J�3E �������fUjĄ��l2Ei%ʢ/Z(�Nf&�TAj��Ej�#��$�f
*9�K�:��J	j�QTEDDI.�%���4V$uku�AEUTz��<�飪"�neqΎ���r?��4�ذ�YU���xq=(0�d�#����kP)vs�|�i��]�m�
u���i�+7-ۻ�s,e�������7K�r��x����7<�k��Y���j�9�����:ry��0 e�"3�ڤ�������'-'jSb�%����b76~�g*9����Wif�絒E<�/�YI<��rz�.'�晸T�����͵�1{g,�IO1I�{���L������؁�<z�Y��q�ҿ��*-��)�����7L��d:��E�d�VZ�Bu�](mK�WHU�R��Kyq��1F񘧰f�i(���U�ޭ}�>���Ceo�E�e'ب:���"�!�XX��k땳���b����f�����j}�
(w3Q�$�uA�f K}Pȡ"�S�x�vZ�=���/�x�dk�ڇ��9J�P]�vAbj֮����#U�;��Ҕ��xq�`{Չ��Ҹf�n7�3��D.:�jй��B��MB��4;�;=�:!U�.:�I|��!�a����,c�mGa1{�f�!������q�i���u�S�裻'L�{��L��IV���l��Z7b�8�Iq����f�ݽ�f5���,$���|b^싶�u�����S��@U��3����=z]c�=�Y(��X��V�l�SW{[,��}�}��[4�g]7\���`���,�sһ'cy:֎%�z|���Bl;�ym�Ȉ�{�'���;�p�����T�=��zݩ'��U1[W)r��T˾hM6�_5uY�B��N�=9��s&>�&������IیZ�,�y��X�!7]-p箽��D����y	�W}�;�kY�����wr�������u�ܬw�_\B�ϓ��ZOw�֒�l��{�З�8\��r����j�mė�3�v[N�S/Q]���bKPr^o����6A
=�������uemĔ¸��~�i�)���-�������Yª��A�+O�f��J
�
�z��I�`q�0�3g�e�Q�J@��(m4�Wn�����v��^�̤�r����	Ҧ.&j{��8����YO���[������/C�ו~޻x;�N�p��8�$�x%%K�i���G;��� Z�0����R��?y>G�U���/Ԕ��A*y���շV/MaP��^�A���æT%�R��.�ݽPY�˔�L��-c�j��i}x�_I�QKG;�e��_kᣔ��˷i�JN��?���舋T�t�z����}[cj%*5��pլp��M=��5P(t����:/�Q3���Fm[�n��PԻQ-颓ˎx�d>��W�RS@�V�ٮ�ؚ�i1�S��6J�-����-����ž������v0m�u`�O��I��ϭd_-&_�H����hj��ި��*94�Y��Ø/0q��l�/�u�s}��T;fQ�JT�za�ѵW;�/Ѡ1e�W�[�����S�ޚM�w���(�Cw�y�똂�Ʌ)w(�1����Wn�ԬڼX��˦�����bjq��ƹ"������̺�Z>)WLMK�3�6y�7�Ѫ�$�U��&��G\�b�2¢h��.��/=q����57����ͬ���_\-p��� �+~c�T�5*�S�[F���@�@��+F_���������̋z�噌��<��m�DR��'S�Ӽ��w����݄�9K�Oo}C�5�,/���4"և����N9�I��]����;˴��v�a�;�E�`J[)N�� N����{e
Ӕj�#�Y�ݒ����s����ښ���������W̫�m>�T��G+���F�������Tw>G��}S���j�G�X.�9���z��:p���������!{�OZZ8ոj��^��v�o���]�ױ��㪰�)�ظ�m����]�^�ʪ|=��H)N�"ze�������	^�J�*�5����>�[1�g�{s �c���N{f�_8T����N�q�})R���c���vr�O/�nk�*���C.���QW�/�C�7�sA��F�K�Pe�!'o�p֓8��U◀�b���B�������ʎ������Q	1ZRW�z�>9S��f�֊�K�Y]4�޽��:��9NQ��Bﻰ��zSX��k+1	�QT���g.�I�v��-�p�X`��ʇ,�"AJ4n>�UP]:�rUu�s����}���.j��w�
���J1?r�pDjqw֣F�s�9�{hbXvl�Ձ@`��B��)_F��:�7�:I��+	��R�h,�,�J��B�^�����)�%w�;��0V]��ȟ!�vҬ�{ÛԞ�u��^l;�7޽P��D�ֽ��c��)����r':��~�����X��;o�5��:���M}6�j�y:֋������n1ڳ�Re�<�{GkV%�������l��M���~>�no/Wa��>\�#��{��/R:��Ig�-썧�����ǹX��wz�_\��w��G:u��z�흯������b~�m.�|��k*�ַ~�������C�;�Szp9��/�m�Ed���KG����}�{y쀉$�ֻ'�ϸ!���x�e���źŭ�f�l۳��fT�/f'-��[�9A��MV�{_*�ۓ���q7�3*M����J���f�gl�F-���%ݥY�.�N�\�:�\���it�0�*�or�|�X��|jw�L�=	O,L۞�9T����yTmK�q]!RR�X˃0��Ç=�1�X{ٸ#s=���>��oT
�
7��l��1Pw�������I`��
N���+b�A��qNF�����˰�xnH�`�����r�X 7���p�]8��8�vM������]�.vn}�n>��i0�6���,E6Xή�L�XCt,S������w���P9�́"]�E"���L�p���s�T �x\�1Ͼ�Ʃi�F��ިko-�y�o�6�
�>ϊ���*v몳yc�"�̻]+>j�9s�ޭ�o�Ao��5�k��y�o�.�A�U�n�5� ��UqOmo�j�u,�����LV���E<gi�9Q�4��V���/_�]���0K[5K��:���W�o�b�Й�˹ͱ�K�l��魏}��q0�@�J�OJ��޴r�.sf��D��e(:��kFPȵ��p�'����|�?��<4�6��g`n�ٓ,?Q]K����z��s��}���vD��O���v�{r{uN�i���IK���� ^z��_j�]��y�����{^9�. ��;=<��eE�����b�]=�vY�yr���ۭ�nV>e�-|�}���e����U�n�'�7��p�po'��o��q�&2�v�^���MV�Oa�1d�i�O�ィ�����7��!V��镍�{�1m
ZU���?G�h�vU���(�)+�v��.��s2����GA|E#��0��<bq<�BY?�m��\����s-�����G�__B��*jCn^��B�تJ*�/��ƕ=�y$�~c���Q�CǨ[ns��n�8fQw0*��+o�)�q���4�¤�c:��=�]_Mb<��gw��}3�2[�g������s^?4�b��#K�nXW�����qt=�<Fvn��|�s�M�uۮ�ol�}H��[R���怦�l�9y�-�����<�4�+�p�[m�ä����v�ꈤ��3:�v�R�X�3krJ�qNéJ�F����YF8Z�x%��P�o3C�SLq�;��
�N�i����1Pe�;�I��ƻڇ�pHǱu!//]f�c��
?F���PBZ4sW�oV'ƾ-�C��՞YF]t�r�\V��t�?"�%!����J��.7B�0�d��U4�K/��������t�"AK h?�j:�n��j�Ȩ�r����ۦy�n����o�P��\R��Cf�C�
���(��
�>�=��^Dj�{e r�\��]��˽�������3��^v�<�i�+6�EV)��dV(��¬���]dR�i('��-�ٷȴ9����4��f�����`�����v��;,8us5�7�&��'�U9��a��着��ξS�=>�&��\k[����O4��6�]��k�&9͗U"5n�#����4&��2�y���յ���i:�����o\��������ոm��j7���_eY�m)��ޞ�O=��x��}k\9�98S.�Nd^ɇsq9X���+(��u�1�/�@�Tf�\@��3�P��z��:�VyA�����Sг��Gw5mQʏד�F�9�����bϠ��_�'�Db�M��U��9�{�W�-IF�;޿a����CUϏ�[=im9V��6�
�����T�J�W��[&m����W��r��!���4�<Y�fP괡�ˁ:�OMD�CW�Ҹ�د��Yq���\�+��'p]M���$��G\Eps��gg����*�J��5�����,Q��UZ�#+#*M�R�^f�Kj��@t�_>Q��_b��zw���z/L�19�%m2`�[�h=�.�h�p�@��E��{�2_
��z���M�Q��xߒ�Cy.3Z��}w�4�oZR��7GD���۽�����b ���8����vC��5�)}G����r|l�av\z����3;D�rp��a��5v�[�UW�d����^���,��~�)T
?wϤ�cBK��[�ڵS�z���[��z5丏�5��nBq�O�r���S�wOŃ��MJޟ�f?s�}'��^�N�F5�9��FGy+�,06��g�B��JXx���8�DN.�.�54�sP鷨6��� �q�
��R�vV`)Q��%B��NP�8+zjm���'_kE�7�5��7�G)l��;5��]�6��^��ܕ��\�o��[Q�븆�N��ܪ���)���c'-FwT��/>���g��Z3^������<�&���u��$5�a}{��ㅽ]k\9紳}��6Z��~;<s% ����He��*�Im�vo%[������i?m��VOu����mJ}˞l���m�T�v�������jSb�b�������>��<�d���Yy�0�=�&;#���jf�2m pj}F��G2F�z�)�)�t;�.�z��Ee9��;x�S�尺�2�X�1����o�N������R6bc&_w�}�����u�e2��aq��<��^�ą��8�.��}�0��f���W���YFy�hv
�A���WVV�ᮌ.&/�f�&�Ķ��vn8�e�Sŕ��X˙K
S�9G���us ��u5�ꄮ4�X�z���]����uN9���)����v�ʤ�p9o�Y��[2�~]��{�f:$�s/����NNzd�u<�����sj��N�о|�#i&&�gz�n�f/2���Z[�c\�Q��놱c����J$u��>��c7AhP�q���/����Kӏ�1ֻ�[�_Ao���vF��x��9J�Qi���"�֗�۩B����բ����Y݉��Ŵ��չ�7�+���P7BYZ��R�o��]��."�yB9��O-����X��D$Ұ����ʍ,$mᶽ7��.�%{��/��w��>���s��O���yW�a�����>{ԗM�ˋ惸�;�WJ%oTy���Zq�z��;���2bG�q>�n���eE�a!���	����Ӵ�:}��F��W�i���+�[w���]�Ev�3�$�\Yq��>xN��$��wӻ���Dt>�[���]V����IY��j�l�ڙ��`5�H��d���Mg��4�N����׆�����0���S�P������fzWۉ�m�
���r���F(����֮�[�ڰ�dC1�=�`��nδ�c��6�����"<F�zs/3�.���{6z`�mďJ���E���4�W�w�^˗P�i��'�$�t2V=��T��!�2٤�G��9�tAG����zK��5lsN,�n�	�O*6��u|�B)��&.���e�۾�{ӴL51^]�K�/�W4��T.�]��j�������f�܅������N�X�)�qo���'��7�W�ܱ:��TGu�Z$(��ն��8Uc�ԇ�-��O��7�9��#'*0�dy{�
�:&�]�f�͊�ip|po����gY��z<7^��x�J!n9����V�^>88�xD�����|ƙ�ne[�ޣ�rs�D�vk6��)%� ��B��M
ż��hv��.��w�V��P��O'��^���݂t��zw�n�.`jո�%�}��3��㧦Z�yzAJ�d>�;͖���#o��q��Z�'Xɣ���j��5���]sge �a�[ъ/x��p�ܴnq�JD�u��R���YA<
%^A��X������P�ȹ��G��'\ y��D{��uL9�V�L��ٳS6C�����7R��	oP��K�����ڱP؈�g%���r�J��3O8N|�Nve\�����`�|�`���;Vl��r��
�0C��Q��8,�����HW�?{r�1�.��6ps�!]��[�G��e��5�¹`�G�o��
�Z�y��w��1	���-sHo40K�mW̧]t���E�A7Y�ٯ.м'��A!l�\<���|uN�ѽ��0ZO=�`h�n�l��	�������Q>Ob݋c�]�k�vN+Z]zt\�c�469��Q�q�|��S1q�0>���HȬǼ����v��~�������v�}�cK�Tj���y��h�/"H�䫚���YC�Z/��E�y)����ќ�$Z�O��lEV/�^r�LT�j�{6��4O�
��ۧ��;|۞Mx{�Aӹ[�gIY����̈́�w)G�gQ��eN�Ec�]'��Bz6�rJcw��E��zU9�7�\�� ��B^��]2�w�v��Z�v0ʖ��J���qz�I�m0���^��vyk7�'�E�=�"�u�A3q\]1�]��j��c��ً�K�t��x�+��V����=�E1��l���O����A���@�������e�o�l�{�)J��}�c=�i�ob,����G��~����r�����q�$uY[��͒���%^��r��;rws��beȨ��E�Eg��UV��EJ,��)�l��)iˡG(�SV����Q��d�^H��:�w+<��4�p���wK��J��H����+�N:%�Qʼ%�$�!.��듲u)�9[
'W%:V�TeD�2���ZS�H.EDW*=[���z���C�H�T�,+:��j�J��瞖!Ds:\�NIUAy	I�yN���++CWA*9G�r$��YY����r8rQr��u��+�k���M����4=ܯ$2��
%��p�Y����ER{���V:8sut�IN#rYtD��+"�*.$%�܀���Nd���f%I�8^��xg�aPP㻃�Eft�F�LL��'vRwT�k�{�QS�\�����/Z�K�W�x�绎����+*3.z�:��.��`I��x�*�Z(�iG�"�H�H�""�׸/z�%�_ok�(t߮o�����T0Y�(��^��V4j(s�zt�:Qg �ϯ&XF�B��h���c��#ﾌ���17��L����p������&�Z��vD�"����<7L�i]�
r�+[4{\esS��Ub�I�-p�S�:��[�w·�t6EU��M8
;��v�}����z���T����r��0�
w<��a���'im�W֗Q�{rV��Qіӿ���q>k`�95�7�M���F�������3����~��V���|P�a���m����q�Xx�)\8�wK���W����O(���*��Ѵ�j'T5�e�QN��z��Ŵ��Y��or���vٙ�d-�z���[�^�H8Wc��Z��������q9�k����nˆ��uކ���L�g�&ԈOjzf9|��G:�cuR�R�记��J�joo�p�^8[I��Z�o����[�hm�ʃ��),RKzj �����zZk2��0�z��G�0J��}��Ƭ�&]���Su��ֻC�K�^ۻ��)e]$�³#Đ��[u�m�ֵ�=�6����䳐��E��C�u(3
>�`�e��mp����eèؐ���:�Z}dk�2�L���}���ֶ�ů&v���PoV�6�eE5���y��N�):Xw
�G�����Z/�<�d�X���wF������*�������\bwn��X�S�P
��(��B�p�\���b9��������n3�����w��9����æq�
Y��`���V�G;���=���J���p9�|oc�9��q��\R���C`sy}E�� NIZ��ܾ��No��rm,��庙}�7�5�15��j�����]��(��dK3F�@�jOo]�[J�O��#����K������X�MD&�Ӛ���:ut��:6]NP�i��e�4)��gW�^gJ�;���c��K�V�Ĩ��6����`�k��k3:��Z�M�w̩�hˌ��B������O\$��V,ת�����g>o�����~���7Q�fTs��v�:��_��y�r�u��t�[��ӱ6�qB�طX���}�n�g1�T8��ע�<C��)iU=m
J�L7�0���:c�2Tڶ��+*c�6��	ɧ3�Ix^�[���s��ؕ�\�;�w/J=�;�6�k�QT�u^h��.�F^���ὝqEZ�s��O��͋f
�ޮ�)M���΄� �V�YG�G�>�;K[uu�ѕԮOBW��F�I����Z�Ϳ���{a; R̭���N��g}B�3OqMN�J�K�x[nˆ��uϾgy��K�5����Lզ��Sty� 6JR#����
�*W[��e-�R]4�t�˶Z{�'��q�kz��@t����m$�Rސ+�e6��u��{y���ݎ{�t<�
R�wϦ
?���wqSU�רq�~�z�jzDzz�j4[m����r���S�}�%�t_�j�
�M�H��q��̀��v��4�֤�������]}�vgn�`eA�P�4�v[�p'�Mu.{��u�>;\���w��!�1`յ�Qw����V�\�qX2����4�+�y:�h������i����wǶ-�nԸJh�v��Ԉ�4\�j�s�i�+g����?n�;;y�/>۴ʭ�#�#�����Y�f�Hĵ}�*�
ǸM��)���I�כ�V�&g��97�כ�k	�Uab	�m�ʊ)FҬ,5�Z��;�%���K	�{fp$�j".�F̂l.��^k�f6�n��}O�}��;�����g�%9�mƻWS�ȟ�����}Q��vW6���On^�a�]8�����}������[�:�ޫ7Q�9�Z��@`I���fb)�{X�Z6{���u���N��Չ�5����^Ls�u�a����a�U��T�FN]��f�~�u��iOVe�����:ũ�f����M��M�c�	���{{��=��KD9rv�Z��5a¾i�T���auP��
/���R���UϘxݯGf��̤QW0���SS����W��c#�N1Xgv^�墻u���|�V�v�ʈ��� ��.V�H[�v���x�u��Ӆ\��+)���^8k-�|�=�[�#��T��l����n��gkj�'�?���T�GRyѮ�p���/��P(t�ύ��o�I�w���4���ߒ�Z��.��Q-�}������R����g����lP}
�n�u+�ɖ+aU��EX�d�����2�v#W֝5��gu�=�2W�=����	�F9 ��1%�@իk�H��ag>̭�}�
�%��{ic���8qvb/��w��5{@Z�	���.m�=o+��H���)��!����52�Ox.��~O(�`����Y��}���|[J�f�n7�>�3}�y �����ܫ;�N ������gesĎ���i&�Uu��Vv��83BSؗ��)�"aR<p�zWd�F�g8r��F�\�Գ^�E=��M�p�Z+���u����aMǝ0]�ܜD W���u��Z�g6sbX�6�ig15�n5�Ю�]�1�t�-lr��M)ކ]n��6�es��\�u�j�V���������g�C:2&�\^@y����U�%�om.ё#Y=-���a��CU��=�]�
7���t�7=���7Y�05��JN��f�ѝO�ѿ�,��`qgQ貹�{�7Ĝo������2��W�fQW�M�lIL+�.,켵Q�Tg�jY۝u���l�]�\:ŷ.��:�UL��>�����uX�ѪBW��o,q`��䘽5�1]_o�5d:lԾ��NU����g�'DfL�)pҩkՇӚ#���/"���8Q�x�6��Ŗ�/�Kin}W��ed�u����O,ܡ��A�sD����Ҷ7���6���sz�;r�m�R��q�0���]�Uط3�u�m�;c�5��m���m�L^�ʊ@l��4��%M̳�vwf�&��R����bt�4�*�5��}p�>�[1�g���TT�6��|Eq���\�P˃��ݓ��%����k��,�Oc��-��v���r�X������;���JK��-�	;؎x���a�<��U��W�p��ʎ��B��IPBZ4sW�oTb|V�����^a=0��-y�p�k�䯏� ʸ)�%u�	�rww���x�NE�u��5ݥ'�q6���[�s6�)�2�],R�o��C.sq��kf�Vc<|ob9s���a�Td)D�܆�b���꼥�a�ȫr�%�q�ඦ��m\o-���o�v9�&���!_�����E��BUթ�ތt\滫��V��Vc߮�5�����~}��w�7�^���C��a<�Γ)�n�0�Eb��� �P�V;8s�7�;z'NK3�k�*v��)��/+��2�lZ+�6r��v���g�#��h�թ `ʞ�t=[���yeA5��&康�""�r<=��j�|�m�����[�H�Zy��4�^�����#Y-m|3:�2�:W=]�j7+�Y�5ļ�m��ڥi�]=��7��=���G���b0/�D�Fm��Z3���j]���zĺ�{kAN��"^"��5G+ם�k9�����zL�
4��c�+;���ru�q�E�N惇X��]��f�E�9Q�fp2��}4�h3�,.��j����T*U�'����6惉m����Uv�,���qY+���U��'����N�\�����DꄯK����nˆ���$�`��V��E=f�^n�>���s�z����U���P[�+��p�q\j0�z��K{Dvk͇��{f���C��%A�V�J��A�բ��Ρ��u+.�����ڇ�r��B�wϳ�I��r:v;"����X�+˟ѽ[�-��u�6�r��޹Fa�;��_#0(�	�
)�u�jE�����*b=+�G��y���Z;r�Uԭ;�T<Rc��kh����W5��56��%�~�j��^X�\��d����*��Q��W�:39Ԧ������]m�.ծ>klHNc�]�5�v�mp_P�ԾL�����S�iBUA��W̶�ެ]�pSJýJ�ߛg*�
�ݒ�����S����]�++����M}Թ�B-�㜵��p��F��WeO_.!Ԁ�*����A���z�
o�\�����u�LuD���띶��ݗ�h����
��tG!�
��ܼ��{:�?E��K/���]-�O��k�:/W9�K)��k������:E�����{�ݖS�qZn�iN����9�|���rmo/W\B�z���w3��b~�Y��)IGy���ӵ�e��՝%�߽���z����t6�/'��a'��z u����^/�&�G��S�[O�S)���rs�K����V)G([�9κ��.��Duem�IP��q1|�6�6�b
�Ӯ�����&��}9�����D�З�����+����sq�w;�r�`��0w�=��[�k}�C�����3��
8���Ƿ�͎*	8����yݕ�`�-�'M�f�މbL�{Jc&C�;��'D��m�a�D���+����vm�Z�1/��	m����mV4���d��\� 9���"]<�s,e���>�{��C�o����U��C�zy��Td-�뷂z�q��{:��#�q4y�^���<�p�=o\��kz��@hP�y ���ӝ�NW �5jS7��6�_g��2ܜ�I�놶��p���-�4�@���eٽ�n� �0��.P���/��n#Kj�k���4[��mj�\f��s�W��B�����[�n�W�. PS�'?A@�KEF�k3෪1>��J/�{ඵa�c���ݫ�����ڈ�fa�����O=����X���LΝ|z���4δ�_M?�4�ͱP�D�G�/ ���zWd�:������[W+�.�3�7N%�SZ�;WJ&c��8�qzkyĮk�Y6:��Tz]�=�k1<NU+9��M��ǥ��߭C�ND��0"�i�;"��Кp2�nd�r��׵��$�����;P�Mh*�TX�����k�f�����{�6��z
�L� }����J���&�S����Y���މ-�9N�1-�a^�q�Vq�X�M��޸TS�1Q���J�^yy�2��S��͈j	`c�Q��Ƶ�ؖK���x7Z��r�T�/
�l�j6����*��:&z�y#�N����F�c��/���%�򊋰2���*�Bq�=�j��3(�b��6ؾvL���x��cʞZ�h��"��;m��y��G��֖�9~��SV���|��V�f)�[�Rg�u��� 5ԛ�m���;6~��������w���=��8)��X��y<|�ʽ�a��e�\�{��sٚ���U 5�1֡��lј�W�	�[��ӑ;�'+�Kb��Yp�}p�>��4�Zm=�}o��4��G\W ��s�=/k�*�J�joo\5��ж�q҇���+Ndf����{{s']��w�xc��%A�D���)<zm�ܾ�&�C�y��+��7�m<㔥*�|�J�-��k0-�p����(T�7��qf+/�y�o�>OtW����2�]�X0R������|��"�njy���&خoj����9{F2�h�B�e� ��ћ� �\0L��Z|��6{7Dqg�4Z�E[sUk9�C�8�eF�<�;������/T�"�0��B��+0v&��N��ǴUm�%Ķ�Ѵ(iѪtͬ��T13��E�^�7(
.f\E˷�֞�Sy�v>/nE���s��@T4n�m��j9J;�	�JD.	gl!�8��z�9�l�<������!�B��*�;&��΁[�7
?Wo3�!��EU�wuz�J
Hf�N�(-�C:�V���r����\4McS�Y���w[��0��r�l[ǀ�`:�Ķ��	Yw��=�l8(e�i]\W�0��n� �*[�7���	�wa;01��#|��i�]I>���3"ɋ;�G�f`�o5��N���F�z�K9��ήJ�K��Tз/g�+o3g	c�p1�V����Qs*�[M��r����j��I]ֺV��*��Im'r��AQ�f�r9Q3�K� ;d���-��HՖE��*�CZ
m00.��}A��[�;A�3�S��X�Ѥl�b���
�#���tG�=/�g�O#w�����I��^6Y�˥ ��ݱI�*�-Qn��\���+�7���l���7fI�<B>���՗���%:=����8�P̥���kdw	|w;�o�K˚7��A��	�m����Y�[���x���$�{�J\�+n󡗳0�);��Ǔ�$R(�d�S����%�Zn�cᜧbB3�$�4�������ؚ��g�.���ZY�k,��lY���|��9�=��p ��c�Eca��tӛb�<�����Q�m�"v�p�=����*L(���@�|��M�!�Z����cx� o<YOEɡǲ�ظk5�r���Ҽ�������f�P&�4t;�b3ʭ��=�k#�f4f���s���n��'IQ�n�;�v*�@��=9V�:O^.�)����T���JJ�)>�[� �D#.��������,�K�p�����̰(���}���NO#
��,����x���F!�]�r)|2V$$��&��j�Ԩж����e��Y/Q�c��Y|G���oC�qi�i���3~T`Q�V�.�L��ݠ��*�[�t(e��S�]�s�2ŧ7gZ��(q�7xA�Vӣ}}�$q��f�J��t�|�`��W{'&����1�%��e��t{���lf��^n�L�^`-iԠ˱�~�w�n�бz�qc���<Ej��C�Q��A��	d�t��5�z�f��H1���j�����������2g1��ǽN�jÜ�����b���3���O��f�ӂ>��ܐk�,7�US� ���u �q�]��%�tb�S/)R�\䬑j��x	Ì/�4���;;�jE��<����v�Ia�5V�e��p+HM�@�i��t�TX��^�D���î�W(������P�y
,V�#��;t]3�۔���tI��e�'H���<�j���/$
��s�H��듞g���-��gs$����E��6�N����jrWu�{��AøY�<��I�H *�qӬ�Ņ�&�B�S���xic�q3�Ĝ��Ȋ<�(�C#$�P�����rr0r5���2�+�f���q���:z�Zy�N���"�Q!2.�k���6q[�9�<ʢ�u�e�d��4�VEE˺���Ӻ��=��y��K=��f�Y�]��W��uA��w�u$�9d��^���-K����9���^���)䋸P�QN�q�� �L�ֺ9���[�����r�$�o�������J[�`�.��bhߍ���-L�y�L���\ENw\�kJjg��k*�v�Oo����&^��*S=R���˕�����1q��Ҷo[c,l6�)�3��%%oa�b܊޺���x�9��ֹ�Mn�&�1��\�7��võpb�`l���b�ќ�%�Rm*@K�U���[ӓk��#ymje�}SQ�M��d��&k2��ٗ5ܧa�Qh9�[ڀ�.�����umDj�V���;��TՐs���@����J|�+�9�A�C�K�^.�Q�Қ3�L���T�q��1�r�ETJP���T���g�k�:�?������b?�C1T���B�v:��"ҋ���o�-����7�ܞ|�^���V���y1�F���|v�&�7T	��sU�)���=ï�*&"����5�\��n}���75�q���vhǫ�[������.�.:��*M����Z�͔� d;M�t���;3݅���+l��*��Q�.k��	hr�0�*�5�� �3�V��]bɝ�uĕ�����w��-�uii��htj�5��<p��%�<f��@�������Oh]r���-Zlx/�[��{t��[Ha�������� �n�it��˴{�$$�s��/~�::ن���b�}�U�9��1��ܩ�w�l�O��Bɀ����}7��#"n�۾�[;<]�u�R�'ev%U\e�vA֜�zdJ�����k�m^�Ϫu����|�e$t�0:��f�x3��ե��5����p�c���"��=�����_)ʄ6sJ������K�S����q>4[�m��q��ߜ�?"���E�|n����'�F�J�[����)�z��*g.��v���f�T2�뷭M�tC�<��˦�s�\=��z����~��C�Jz2�=���w�+����.l���<�m��jOG�����J=R�y��z����x�mL����q��\N��C`-���H��x����޵6ґw&2y7�53�,p��7��WS�ȟ������F���Y�˪��O!z����>��Hឝ퇟��<�'��gψ+��e{*/�<���'�h*�~�VZ�Vs��i�6�<���h]rm��Ov��"�����n]N���-�BS�6-�h�4M>��Vʶ����wc�rVV.��Ⱕi��4E�.=8����/b����_wێ�ٔ1K�����ٓLV�Q:��b���u�b��w;������>{��۔�%�����Ck/!�Z�=���M��ԧ8��h̢���Fn��֊�Y�>�����{_J+�q-��5��T�����O�f"��ry�W0*��ۉ*�.&/�fF�̻�٧v�K�v�9�n_f�͟�l�E �*�������]�y�R��OM$�N�&}[��h��W
���v��;�{1�g%�=,N�}�����߽5���Z���T�Kyq�ˇ���O���@���r{�]����ߪ��J��ݕ)�H}-�ԞtF�ko�p����4��0�j�Z.'���_G�=B��wq]Z�|x����ծ3Y���Qw�xWO7�y*Vu����Ps�wLA`�KEi��_9��ё�wZ>+�	e��<��Rw�G*ś���Yϑ�J4i�P�����J���g}x��q�����2�[�D루��0ٹ[K�hf��`F�6i�i��%F��t��d��ݿw��ৣ}{VX�s�1��"Z g�3��v�'4�L��m�;4u'�����L,��� �^6��{��ꃝqu��qEVgs��w�6�|�B�o�(���h?�i��}UU��z�s�Qw�/y��Z9P�9��|�n1ܰ�q&:eO�k�#������9��;*��\M��{�kS�6�jsI��p��5�Y����6�$����� _�s!R�����\��^֪�i:��k�5��vWw<ͦa�ݍ�Y;�VzR\�g�5����{Z����>�8�g�o
���Y�OPiv����ޣ������z��C��vZ�C�K�(��7�(��Y��VͿ���8�5p�n�n�[�u�fQW�uel9`Y\Ad�3v�=6�+U�=��k��źŭ-����9������;P{;M�ܢ�3�m�5Z�WT�J�J���alW4޺oS�ݸw���b ��\�i�U����He�y����q�~P��_�[n����>Q���;2�8��,��r�:�"byrj�/[�Q�m��kL�.�k1w����ߗ�Ǥ!`咷�K���|i��=�g�*2�8{�{8��m�F5�8 �U�]X;��=w�P����"���ѵ�]@\YW�čK.Y��.���gNjm_n��5�4���sը��޻x'˕�������"R�Z���\5��]wf*x���	縻n5:�0T�s5�%b��%�2�ș�u�/l�֠57�wC2z�E=���u]��WAwϲ �KF�j������V�s�v$�Q��u�o�<���r��!O|��:ц��T�l���cJn�<<�Cε��&��޶�X���|�D.juk�.�
��r��8]6���7�һ3�'���G.sP����Td���o��a�껮.��ub'�8-�t6#���Z�庙m�ˎi��fXs(�9�PG{�r���Qz�h��u��<����"�[�x[�O�vJYxq�y��=SV�N�S./�����\�.1"����2�/�s���$q�������<�L���5\�^�|�~�~~ ��Yfz����l��r{Z�l.������ \�E��c�i��c:�&��$�	Tb��IoCj�d^6�o���}��}�]@�R�����\�
� �f�jQʻ�R�ַ}��䃡�7�aߺ�=�)6*�"ģ��]�5◛5�uu]�}�Z�9�פN�LL����Yxۭ��)���|��ΆW޼��7Q�f,�� E�U;��r⋬�\�m�]Fn��$�:�i�)M�6�a��q��ޙ-K�a�����^��͖O�;s ��U�%CW�_alW�&��-�⧧M�e��L�{v*N:��휖iW0��j\�ꄴ9]��Q��ː�X��*���\�Gn�j��_���u��0w�obŧ���
���)����[ϥe?��ˌp�^8[I��f�cUo��Q�Iء&c샥����ڒ��\�z�W�禊O/�5��g<㈥��LG|�5�V�Rx���*����ԱNwJ|j}�����9�6�s�����]�>k4"������X�)h�)�ςެ]�I}ޥ��	���q&�_*���Vw�B��D�Ϧ��\�!��|w�4>�������輝2:��9z-_!��KD��-�/�j�����՗��&�3�¡A�Z�,n��AE�o�dcM�B�c�Q�P���X�З��c �)%hhmU�-��U��76v�j�t�נ��I^�fG��ܡ��)��s:'�wF�6��v��2N9G>9`K�Q�l�ξs�Z�&�m\F�v!�s��_t9�}KV�F�ۻSQ�0�7�\��&9�V�v勭�%���5�&I��H����%�ϗwL�Qu{7��~<w)����y��q��V�������=8�{�:/��ֵq���~����c7��gC)l#���AT{~ �[�η�����[n'����7);�2�������L��z�ڪÝ���=�辳u�2��0378G1}�r��iڙO��V�U;���;����s�j�'<K~K^_ZZ!���SV���o�u/,��S�/79�\�*�`��vm��f�\=���s��7�0�~�.X�Ĺ,��{n#�Ҽ)���܇m��粌�V���1U��4��D�//��6��Թ���u�R�-�8j�C���'���uA�5�W�Ȣ��Lz_���%7�&s��_�9K��T��٩���6�̻ν���n�Y��J����
�w��t�C�Fd�.�߃��飃Wh�����aT�0P�_V�ܼ�̡m���#�	c<i�fw7�n��i%3m�[n�f�j>�G�N��%�p`v�mJO)Pe�:��᭼p��Nc4{L݀9�!q�y�Q�F���(����RW���K|h��mc\�~���`齍H_��ޢ�(;�^�O}�?�W�y��������h�(�<��
��ws��%��Lu���<gi�3�=	H�O=��\�"�h����P��u�|����N�&҆�4ͱP�D�F~⋠R���!ښ�7�l��J�V��+��ƴ�Z9_%�k��a��p�
�L�w�E�F����������{[�;�O]��ig1)����9d@��^��a�o���l��Vc�����Sޞ�ߞ��\k��?W�^߹r�v j኶r��;�3���z��Eiv�3����o��j��/V�Ρ��q�潑x�L���S�������*�]�;�.��=�.�~cg��ΎX"�҈���lh`������$e�>��v)6H��C�m�y�n�s�G	C�+@�(>G�b� ��r����z��f�p�y�����*��m��"�5�x�I�&��n^�y[���u�~㭼������ S��y\�Y�`8�h=����=���}�暜���tk��Ү`>I)77h�^�gMP�2[U�i���|�6�6-�-���u�l�휔�Ĭ��۪�G�yx�:�`�T*U'z�-V�sM�C���v��.a]���Yz�Y:e� ��A�[R�ꀷ���N[oހ��燨���ѣ"�'���C{"8N��J������2�rR�l�������e��F��Dvk�t=���/��Q(��'���J�&�����w�?\l�����ӟ�?���Y����a}���+c�@o�������p�5��j$�%��P���U���9�Z]��ޱ�^+c�7��}�q7�ZG>>��\u������둷������,���Zߦ��+fm^8J��索�7�>���gQQ������c#ӝ~��L��q�z��Ӟ22���Q�M���j��M����2}�Ǥ��-
�.=����|�F�&��b߼���A���wѓ~쩷���Vx���K $���u_��d�&K%m=�w9gi׎ةs��D�ٛ�~�@J7۽�W���Wv��k�jJ�oX\����Z6%v�/:ʋ�g��>$��A�=�e��QS난��E�;�)�+��� �G �����'���m�$`�}�%]��]f�/k�̈�t��G*c���G����b���p��觵�����Gl�n������R��0��|}�-V��ۗ�՟w[�[w��ڋ����ew�-�>���?W�����B��yRF�'���;�
�k׺Ecn�h�^�w]��}���<��Zw+)�D'U�r!��R��vTO\{.�xܛ͖�9({�ǻ�Q�r'r�eս�P�}5��pԮ'Nj�x�vڸ�:��'_�x���;�M�C�3gʫ �[���v�V��ЯƎ�"gPS����b�S*t��+�)�޺�{=�p�g���0�����gy��F?DZʖn8�wl� �C:�U��5k�+�O���^~���99��!o�h��tw��3�E��u�r*�����v|O������1q�U�7\��z�C�S�l?��{��s�W-���؞��~�,�]��n�.��v,�O�K�*��R}��9�[�]'@D���Rh��'�?V�My}�����}#��G���~s�n�+�l�P��T�I`(�����h��`A��=}ۦ��J(�Xw���;�,��������*�z�0:b\�E��r�IWj�P\ ��n��2�vPR��Ƙ����0V��6�!����m�W���.���\mǡ�����4=�л�ܑ��=a��U�����V`Y������%c�[���߯!J,�(q{d����n�`q���i��B��b���)�����̧i��f�ƵMR�Q诗Z�$�}Z,`�a,�1���)�/0��pH�˙�,�Y���V�`;z=Pf��-�J�����˼k�4�׭��
}�ȃ� 7k W���V��͵�8uh��7��!ɩ=n��.�V�7A'�)]�7���O;�w�8��Y5�*2�(�E�! �R��{��1�
R"L|��OxtK�,ɸ��S3r�E��]e��u�W���6�d�XO����9Sq�%���u���Y�e�rw�a�m�|�2�QKD��ƜF0f�i�25�(N��	�رwmD�j�pui��R���f���q�=�v^gv��oT���v���8-��e9`,�)d��Ṉ�����+pw��
�*�M�u�~�2ճ�{W%�5s]��fK_ �f'���$s�v4 �lU��$�ݡ�elWZ�
-L<� #4ґ.��ʹm������̝Ԫ܊�
絵o�����=P>�)F;�L���`���]��>�d˶����
�mu����NԾ2���K��@��pC�ћ�eN	������ �tkjD��3z߭��B�'bn��HV1�V�0����n2z��<�9��Z���6����
�%:�
6�*�O������mk���dv͠�����i!x<}��o��h]ٗ���-�$SBB�p�}�h_)���f��(����/��&�mﳥ����\`��Q����=�-;�{82xf�8�EE�&�J۱��*ӛ�n�Uq5n�S,�ܕmK�X�O��7�3GO	J�b�J���:��c�n\�Nwۆ��/g���X�鮻�$��;)l-a��j�D�+��՗��TnK�:f���d`}UD����t�m�m��h�	��e9Gy6�tApu�Nv�i�d����op���`�\��T�f�85�	��[]b)�&.#V,��X�wǙFg��l�C�l����N+�L5��e�x�Jq2�H68i���,F����H�nB�M�(�A�չ	�`:ȕ���WU�T`����B���.��+�x�_If �B�k%�:ﻣ�5��⌏U�]Z:-gͻ*|"�k��`���I\n�񽰚��%��d蒩W�c5�O^�ڒ�8򋷽�h겋徶�y-'�G|��m��ѹҐ��W:��+],���"2bM.-7n��J[� �;8��/�wPf��0�P�5� o�93x�AǳI�ê=I�#�g{��(f�V�̴t T%"I^LA�73sg�.�T�'tH똗�������c�u��w��2�]���*"�G����t9K���a����Jw\�=�c��^xn;���!�wKZ���&;������Y����h%d�x(����QDHIUU�w\V���C��$Y�j�����벻����^F&�T뻨�7t�� ��J�R�\q���&��9�"���
����(�w;�L�
����'..�W��$UV�Q2wq��p��(�
�j^�x��*��s��W�*=q��3����R=V�`�*Q���]q"���J��	H5��*�$�L�ۺj$I��P*�*���p��s��g�\������Oi�K���f��\��tGu·/*��ܼ/A*�9N��YZԄ�q0�+���R��;��6f��q�u(�D���S����(�L'���(c�Y{	��n��]�Ѷ������4#�҄$�5;���ڡ�˧����[�+�ꕇ@�Ե)���ߺ�P����{�&����zG�����T��4˿��Q�c��W.=�N�����(���05�q�}��k��s�~�&�޴�g�=k����4����u�䝧싓~�8N��6f=t��L�\�g� ���7�Ft��;��q�Z2_�������U|m��=�پy~}^zO�9\N��^���d��T�wx���z�W-v�^�*���#��XG����;e�*��X��z�>��_G�0��J,��d/=����Q��h��Q�x����a]ػt��}�Ƽ/�yUѸ^u�}�W���`�R�d���gӃڱ+ެ�֤j����TZ�荹~=G;��~�d{���H����{"]����dҟ��Y�C�M7s�Ѫ4���B�g���GG[W�u)���ۇ�	��}�h���F�ڴOӳ�9��^��[�%��M�r2ϴ�.�d�+�l�w5Y�):D�Gu1��Ꭻݑ�~����8�o��^�]s�������K*p��|N홇��X����N}*��`
��;�mA���Y^�s�/��yD�SpsOI������,��)t����3�̦i+W��aQ5�f�0֩J��|ᣇ�g���/��(r�	+=��U,���d|1�D�gu�9<0�q�ߖ�j_<GeoA��y�xz}5sK����n�v^���c0-���e\ߴG]w��������Y�҃'3`�<5ʡ�ڮ2\��^3Bg����-&�M_7+�@}��H�r��9^�qϩ���k�gNI۹d��/A��~����ߵ_��T��u{>T}�l��GK������n3��}�ˏx���+��V�>�h��<�:�~��7��<�~���h�|'���S�O��n�>�a���#�>�Y���yg�o�ח��m�eu�O��7� ��>�$Q�0G�����b���zhO7^=ޏS㑾��j�����ݟ!�d)	�|��;�o�:��F��2��R�ȿ�e�9�뇲+޴$\���-��0�����֣ۮ������*����q�u�\�i |L\�\M�2�^���r ��z:k��C��2�����N�0�+�����~�T����v�sH��H+��e�tL�F�珜�9������j9h�k~����ԁ���=��h�fQ.g�`̶G'+/>�p���u�M��D�W�_���Q�R�n;��m���n�ȟ�H�6��9�iFz�x����\{���ѡ�e��&p����_�p�)�X��LT��Y7VN�gA��ݣ�B�����g������9�M���lW�\�5������ZY�i�;o�U�@Xqe����ё�ޙ�Y��8X�]������0�P��s�ĥ�╋���D�{M��O��*|n9��=���z�����f4V�V�/�@)�L���u�fI���1��,_Z��u�^5������1�߭d?"�z�v�F(�.z)��-���,N�`�[�á��0�����N�=�Lxk�2C��ʊ�7;׾�T��=��#��Az^}[��t̴�~�	b�9����f*�U-G���6�o�̺�����@zS��8�w����*7�uU�s/��/��dE��~Ł�Xa��6'0{�4Nڟ�y{yV�z���2Kd��ٟ@��yߤ�^,��|�g�n�,U�k:rN�����"MbS�}����9�2�σ�U1�ޡ�93��4����?q�d��g޵qܫ /{�q3F����5�9S�c��R��[��ρ�,\u�z��:��k�X|=>(�G����	�δ/w��'��3���4_�[�K>3|aụ�Y'�`�7c|�+�u�>����ʀ��~�1�z�_{�;�n��q쐷�?[�M�����#�J�0���x���csݘ������>��u����mN�ś-�e�y;�e�-~��a���Y)^�HT�x���r�U�l�2��3�\���+׷I��h7�kЎ�X{B����i��<f^�B�S������y_O�s7~�R��ܘIF��GRSX(��ioe�Wj�����q{k̭��P����m��
.P yJ�����c�����M��}����=Q��F�+�>�$G�����t{}r6�4���dI���1*��Ë����8Q�>=$O�ʸ�)ߠ9�o�h�m�~��x�W�\zg���{��AO�׸l�������{��d{�>�a{`u1��49Zw��=o����z�'�+>5��od́/U
�G.���T֓�ڌ�=^��P����L��f2%�z��:\o>�Lu�?\�� }1=ΏUfV����Q�l�5�!�`��]H5
Y=C&��*S�w�~=K����DT�^%�f�!��c�?z������~�=7�ɡ_kʐke���څ#��	�u9r�vC�����gˏ��x�u)���:�#��@z��G�*'��t�V����p�n��A��������w�|�y��:�k-#��q:sT���WȇS^����Ҽ^/]���Y�l���#�|�f�~�Ƨڌ����:O��8=�U�teJ�9�,
���:~��gi|b�ml����r	�qu=+J��o&Ō�L��J�8���7y�ZF��dRs�k��EO���+�����W�����%B��ljP!�r�-���m�v*ޫ|�f��f;E�H7{� �p�Pom=�Hoe���ˬ���(@rۛ5g�����fz��<�R��L��J��:֍�����~���]�
�]�:nd���X����_���K�<�4׀W}~y'/��0zw6*�A�Ӫ��%»������T��]���ʝ7Y>VfzXȎ��Q�rx�K�=��_M)�rE{D_��Ց����W��G���F����F��$�/Ơʨx���I��r�z�m��mVl�I�G��px�Swp��{NF�G���X���ɺ��l�JX%L�.�;`�S�-JF�^(�X��P��2�F���q^�\Mķ~Ӑ�#���ίj�ni��מ�t�D�nM�a8����b��g�����^㌶X��u��?Rs�ZF2=9�\}�p�ǫ��<��Hr��R�D����E}�'ơA*��"bK}$qs�q|�Wա�"_��%VJ��8]]=I^ypU���=;����'O����eX���O�J�¹h���]{5�6fTz���yf�N�Hc�����>�"}�N\�X]D�d�d/=������k�<K ���S��}*ǳ�_��q�n;�ׅ��*�6����>� 7����/��K�{�~���cmը����ݶ7B�����]��"��؇��v�mן]�~_`�m3B8<@*f��8noL��H�&�Uƻ�p|�uT��0wN�a"������~��G�����r��[�nYL�?n༠9d�����ʏݦ�tƯ�iwn�U~C�j��6��r;��~�g��p���oޠ;���Tq�L����y0��W�p���u�@��<:�l�}R�����O���T>�?]���<�ݗ�+9��{l�r��7S�>X}����<K�>
4�}5Y�S�N��=}��<1�{�/[�J;޼9�7ˌ������a~�V
���LRyS���wn �?T	�,\�U�ȩU�w5[ >���ۚw"Y;F�m�����D:����z�Y�V;�vO
�eN��E������U{�7�K,�����A����o��ν��;=ƸQ��Ht_�%׫��r���k�gNIۋ�O����&��������N����W�HUo�z6���*g:}w#O���g����u���y_�d�p��Ӓt<�8��׳�Uʹ���U�Mz&x:�=Q�uJ�.��f��n�<�����H�zr=����wWϷ���f��3����܍{�lk�RA�2�����M���׽V&㛿��>>����I^'t��F����[��/1Tv���ñrQ� X�)zd\t�ns]�g��N���S�y���ev���J���y�s�Ux�/��9�E�h�T�s9���k��u<��J)��6~5ݵ�3���,�L9�p�;/��妣��w��#q��cV��j��좛��Fev9`�q
x�����y���/k��Ky%���=�ix��<����t�ާP�g>D@J�ω��n���Ҽ^��'}3q~��y�]׉vۆϒ�|���\�o��p�}���z�q5�O���F�1[���!~OM��	�r��*��Q�ܯ�5��F��!�[g�H��x�δ
�sl�%��a��~S���W�Jz��$z}�B��G�}�_���F�m5~�p�>D��O��`Ρ�}�~�������C�Cg&�A��s�к�^�yʟ�~�����\//Y�L���m��<i��6����&��o��OfIA����}p'�b�k��m)��nφ��ކmy�3\Y�����i��z3�T�{���ǫ
�ו"����D�}bwL#>��(���,��K�#&}�د�zC�{|2��9��<V�h3�ͽ��r�:�߅���YEۑ���D�C�k={���Y���:r5���~���gb���y�F�N��NI˅,:�f���x��uٴ�{��Lu:˽9S>d���>�X������P�|�{�ړ��pg��տ����!t���ƠP���T^�y8��	bx���s���7��`���Z�[`v+h�h�.���18��C^��g5�����y9�
=���ڽY\9�|!<���s_re�k�nT)��8UY��G����,6�Va��\��=��%~DȤJ8N���ﮝ����9͙�Z=>�z������t{��uUM�4*f��r�N-�Vx�FvT鸲�P�@3Ŏ��Q؊�A�~�F�W��|��ݰ����ý�x�TǷ��xi�嵦T<����~��u[��>���Pu�^o�Eu_uWu��ҽ�=��W�#}�w>�Q��~�=�хO��=Qa@��^������B-��O�w[Wy���ܮ�q^�\Mķ~Ӌ��{7��q�U#nS�&c��7��N:eM;��ݏ:��*�73̼�Q��c�'޴�A���ӣ�=��zi����?�>��=��[O��<H-N���p�:��'�Hǽ9������@�Q���f�녋�������V��W�$鿊U��d*�V=z���#o�J؂Tk_��X�F��ĸex���g<KϝF@�N� ��0�p'��K����{MoJ���3�qF���s�פ`�Fw]ȸM׉�������`����A�,��>���պ}A��?��E3�8�u��l��ĎC�t{3�����KFS�x@n��O+��k>X؃&x_u��f�y�� ������5]\��W��i�i�����S1	>��I��g9�,-2����U���!<�Ct>�]��vL�k;f�b=ӳ�� ���N��:�ǎvFS��{���4�_�ϭ|ߪ���C��7
�}�*A��d�Ǔb7�}��-�7Y~���eu�N;��Ga)��ʍ�9z���H��m�N�#�t*8�7o�4�Us����|���*pm����k-'�N��/���Ǳ�׸��?J�y�;A=��"��IYb�������ќ7�aʙ�=P=:�VYёR��7��������0j���Z6������E~${�϶�551K�c<9��(�P���_���yk�V3�-u�����9��Զo���R�>�x�wHof+*f�O�|fzcg��>=��k�<ޱj(J�m_��޼���z�C�/�E���{��垻C�d�p���R*(�N��J��.����*�����3kн�^�����xַw>G��9�/r#}p���μ8��\���D�W�壵���.�	�$����uF��6|3�wG��ި5��ND/H�|s}!�����T/����eO�0�k�~Zk�`��e�0��2�C5]w�}OԄ��ք\y�q��^���c£�쐢�G�� �s���#02H�{�d�ֈ��-U%�@J��N���Zp����%�1c��󂪻u�NRM9����d�3��2)�4N��.A�k�~�C<=&�(H�:�E��_��	�����C�6s��˾�Mȷ���-Z��6��^�Ӝ��<��OƱڪf�B�C�E�o���#��S��z�Ј�P|r�<CT{*��im��Ǌο��t���q:o�ꉨfK*�n��<LOҽ]G��}�^b��y�FwU�m��F�^�ۑ���c�H�`��dߍ��*Xu�%��L����#�+x�=M��c�T+ʏ��W�^}޸~7�f����Q��^�=^ o�`�3҉�׾Ү��E�n^�|���5��#��O�Z2O�r�j�����=�:�)��:/ސ7�!������0o'�՛��w�,���pe�ٹ��a�A-}����k��y	��ϟz+�W{�T�8��a��w��W_��m]�+���UD��8�W�te'H�ϻ��v�G����.�����a5ʟ].}]�ޏo*^/{�`��b�~�C>��s'�W~ta�b����;{;NeI*���
�m��@����u^�|�\�ϟ��qϻ'�g�� ɻ�3uBׇ
kp�r�`m=ۜ�u�%�^�L���!�^r}^�zn#�V�ǵ³�$��r���~�n]!��<u��(�Xe0NtZ�9��-_E�%ǻ:�-V��cx�u��V��m�2|1�2q7Òc,��ߍKjL�.7��(����$]��W�!��feFb�<ɼ</u��[�h^�qg�@��n�M�ƩyK<�-��m�A��T�C�E�z��7�&�s�Rk89P<��[��OoCʬT�Enԙ�J��w!=��ɱj<��.�~�n!ˆZ������&����Q�ʽ�8�!�>��L:�u�w���5�r:��K�_]�yαH�� _*Y�n��m�n��BǍ�bP���l7��o���:]��J+;Z+SXz�&���;���NR�2��f�j<(�Ϛ�Wy*�KD���F8{܏��X)�%*@,���ES�m�n�mT���/7[x������q��go�����JT4�����Ҭ&��@��睨����d����!|��Εjt��U×J>�[ܲcJ��e�lV��5�S������+4����Jw �dG�*�Rʗ�/[Qa;JI�;��N��4T��9�+�c��n�ꡏ��'���1�g�u\�#/��;�;����Eg,���ک���:�ȘGXvF�yE�//�ݺI V��Q�	ff������o�sn,!Ex
��1�;	��@I�����]�ӷ���:9Y�r�ڏd�(�ȧr�:]9H�T�j#�^t�;p��5�ۜ��dT�c�>'�w7�{��榭�)p��<t���+K&�\5MP�pƘ�/�X����Y����i\'�����g��*׌�/��i$�ʆ㶦p�#�uk�'�i_�n��`����[}�x��s_��ͣd�50@�)���p�v�=��3fp���zbu-�z����%�{ݛ�q��Q��9+*�f.����ҩ�o5��E��k6T6[���ы�d���8+Ӳkwٷ^pJ���np�D�3X��.�g����3����F��w2i^�\���=e\x��⊰�B���kaoŎs�Ӛ�EfH��i����C
(�2����ZgdJ�y�L��o�'�f�Ů&��a�L�"�
��:��AI}mǉ[*�n��p���?@}����z�Q�#<)��Ӌ9�VUH��������M�������ͼ�Q��그IM8��Ш�DX��wU�#V��2*O0�4�,�+�]ǐ�{���/R��LnP�����o �	3���_��լ��]��{����re_f$wn�j���/�;:�ʜ�N텹`@��5����,Vh�.��@>Μ�j���;�2rLK!�*�r�����ĥ�%rxG�N�	ݺ�<U]����֖+ڽ{_;��K��/d�&�3.ܽ�{*Q����h�cӜS��G׻�__J\��C^/I�^{R�Y�L{Q:z�]��a�Vm�@6�y2�}[��6�q�'(�3#jǷ����]O�J�)Ln��i���WOmnfSX*אi%�W�!$KH��3�7q#sێ�Qq2u"rN�'��Q�/OWD���B��Bn����^y�ʊK*��]#*XN烺�]��W��"j fz4!�!�/T�P�K��:���n)T��w�E�Zy^k�]Ñ��\�:�wC.�.]n;�9��r�WtH�AP��R�̸��GwpӳB�Fynn�F��I��!i��$+�)2���9��C�	;����r�B,�.9,��"tJ�dZ!�H��wU�*#�](B��Ш;�y�G=ܜ�κE�=<�\�/qӡ9��(�t��NN��<�B�O���=�U\㺢��ۻDF���^By쐜�1+�<�
�U��"+DN*)�ܡ�uwwZx���;DNPE�@�V[���飺^�YҺIp�݃�n���Z��8�bd�I��銎�)�J;����E�V���ڹ��B�j
L�si�ȅ�4E��X��`�tZސl&i7ܜ#u;�v�Nx���q=��jS|�����]��-��+����0�3��t��<�t���i�x���}����K�w:#�O�3�v7=�Q�k�Y>�4=���}_L��	�{3>���TQ�^�>����H�xr=�����>�v,{�)3S>ǲ�Vz7�m��6
5	���,	�"��ҿ�WE�����ܽ~�4��#ׅI���rg�p�����G��}��a��䢀Ze�0
^�2ۜ�]�{R���xˠ�o��Zx$zsz�d7��V�ޡ�_���J�X�(�}�@�3�[�&W���!m�^��9j�/�r�>L��Q�ＪyZ�^g���q7��HۏU�Q��L�fs�6ma����::��}+���}��L�r:ј�o��������x���2��m��/M�T̩��2��6=f^�� �,VD+���/����m���Q����'� �|7�De^��Ҍ}靚�s��5�203�ߌ�:6*T���^�y�*|y�c��y]р�B�ˣ;x{c�+�ZX2���g�9�y����L�>']U�~�N��L���k>�� �)�g�g��[6�mp�tŤ}�c���c<^�uj:O'r�OVM3T��iQ�1Uu��dn`�E�������i06����:o�G�"/ z_�8�/������;:(�l�.�~X^b�/|ە��L��EH����Q�Fu�쥝�ey���.��������V
�*EF�O��zPHWJ��[w�����;?D��K �������߆B�W�}�<�}V��dШ^ʑ�����^+ΑWn_��LϪ�ۭ��W����|jW�>�R�F��gΪ��g_����m�֊���^�uXdOTV�����z�',���ӕZt��F�e��^w�����Q�w��w	h�]��5EL�_��j>�6K�g6&X�'�Ϻ��b�9͙�W}^�^����\2�ʽk'�΄��P��=4_�W���|j�%�*=��~`�>���=�o_�ì��O@�}s>� ���\�����������8��{� �i��ʞ7ez��x)c":�zw��A���ݝ��z���WnX�߫��O�܏u��~���h�i�']]B%^K��o=�=�yiwk*k���s�+7�p|n����r���}��j�:��d�M�o*Ċ�\__�|�xn}'�s�#������9�~Ws�ZG�<W��tuǷ�#o��Q�UE��m�{����2�����<u[����55��$ps�*ў�~U�.n"Mv�o2*������4�H^�K�F�s�1M�\�:��Ks"��;;�����+�ư�ݨ��� œ��e�	<�54vA�#�f5���l����tE��mm�[�]+��g�̂�GA�RAJt�2����9�oZ���?[f2=9��Ԭ��}t=��7�3=�y�|���Fr��9�"��jl��w�� �q�q֫�{`)c׾W#}]��f?v��1B㚦��y)���/;>9ӌ��G�2çR)OA0������F�'��x��.m+�!�P�k�٧�nԆ=��E��q�O��c��??]H5�OP0��T�J�-s;�fHg��u����r�z���EF�m��ߪ���P���q�W4+^T�],�^��{]��.�7R���da��{�>W-#�����m������rz��)��ݕ�ˡZ�nz�8܌��[�����>D�d�(��c�����"k/��K�t�~7��=��k�X~=ⷍN���u�1ٔ��wz�~��_"��7�9S,z�����QѱR��7�X��<.=�{��T���u�_5�߸F�o�*�~ڒab�㘄��7b��X�\�ٰ�K�<���X�E�헑5y�+�@z/����x^�x�C4��&&/n�O�ҫ�����ކ�լ��h�z'��ś��0������.v���Jy�s��Ȭj�*����\�_�{�xsi-��׃	JՂ��Xk3N�X���uA�7��;d�O�<�PTm�0g5ɶ'�P���(X�=
�O��)�U��U{Cdx{֍�9�*|*3� j�]؇�}�"���w=���Ͻv��ț��dg�Y'NL�>��s���{9�}�o����f��Ӓ�-T����>�i������~u��u�E���V�C���ox+�'�(f ��]P�6�"�F���W�Py��^����g[��ښU�k�dd��;ޥ���t�\`�� �,����i�����)��������N�b����}��\e'x�r�k>�Rt�{����L�C�,�( %G�A����>G2�n�^酱?T;��*O7��z'y�}�lc��q�z�t�ޯTM3%�`�t'���^���Oz�t����9�gR�9yS��9z/��ldz�>χ�&�����+������ۚ̿����~����77�����F�>g��C�}�j)��Q^s�|�� 7�� �uD ��EM�3�&h�oz�$���g0��8.Jg(��/����q�������:7ޠ;҅��=���J,c�7�?A���]b��1xex�ٲ�ǆu�~�>�F�ۇ���S|/h�67v�b��z5��f��B+R�yj㓘��,l�㽵8T"�:p��ɔ�^D��䖽����?f>��u�<������|[��
�Wb��SM*I}\:�ȸ����}�k���8$lޕ�p:�ज़���Bf��X�O��d{}���Ef���hM�:kO������a�����x��N�=��Lz}�d�xD�\�g^�R�X�����oԼ^���덬+�SgC'0^P't�7>��+�=u�}rY��Iw����
�ܭ +q��ȇU�`���̬~�Ǭ���eHA�w�a�BﶲfG���9���i8~��Wl�T�����B�w/ޓ�Ez���S�^N��9'H��:;�}<g���^�l{�U��>�{]UGk��9>�w���W����eǼVDW���p�uw���}H�7��Vy�_NIb��'�e�_	�uU^����E������<^��;�7k�Mu�f��6�3�E��n�,�7Ƒ�Q���X<��J�2��f[��o��]8M\�!�β+i�������t���v��\>�6�8�Q�@�,	�/L���m�{u��O�6�Y�u7�}���~��Om�"�^�����+�N�L-ҨW�_Gʌ�C��N���ۏFY�q���O�������[��W���.����3�ӣI_{}R6}_����<�o���ߧ�1<��瘶$�d�ahK�h��;�ȥ�:������h\����ۖ����BoU��7rё�j�w}u��y���`�}�q�t�0�8V�������\nu�K{ �[r1fU�����옦�͟W�ӻܵ���t�5ӫ�]�-��v��)b�:�F��h�m�߭�����9��+�ߝht�1�1
�o�#3�E��Z�����}&ê)o�"����������/��|�F�j�E����`L����$/wۖ����6�	���3!�31�6*T���^�yʟ�~��v�sV�r�9��q��{��>���u����7�,��0�b�Tm5��z�{�&7�o\��`�����}!gU`c�����Pu7���O)�#"5�H5��'�&X��	���"��G�N��ɛ>\gx����p�^��8��<ido��?Za��h\�^'3��+��l9O�������|y�u�5��ύO��9���vڿ��W����B��ۍ��z o��jͼ�c__���Ƨ<��Fρӷ3�4\����]��%x�n2e���^C�~>'>�\�=�o�=S�*��^�}9���z��+��������ֿ3�Z����3��>��{ѻ^�����K��x}�]���W����ʝ7e��b���>�7���C�Ճ�)�{[�PZ�"���|pg3��؋J�e0ֵJK+J3��X�i��-��n�� ۜ���:�L�Z"J�/1\�PkϘ�Z:./�]��-��ۡYl�����f@�N�<��)��pB���B��X�n�U
Bk;GT7�םW5q<�rE{E�s��c�S��W�V}�<���]�(�d��3ƾ2����~ב\"l��N緒���t��*KwB|��z7�|�?�}@>�~�=�>��
�\�iI@!�W��r|;�C��J�\A�������}^�\Mķ~ҼG���P�ǵT���S�o7����/�OtM+z��2_�� r���'μ����V9~U����"<o�iQ�4�:��ƽ*w���{ �<ڕ~�����d "�'�Dķ\�X��#kT�d�[f��|����A�\�m,j9W���:g��O����Nd�6ja���A�hg��/����C�k�`�S�غ~��jӫ����2 ��ώA��%�ި��H
Y=_	�^��b�_W����Ozx�.w����Ҭ{7��ʼ����~UR:�x�dO��:���ԃJY= �����7;>��lz�w-pU|��j��#nZ=]�J��y�Q_=� �߯�q�<��{*A;��)Dˉ�E�5�։�7O��}j��}�-#�������<�O�h��P�9�Z��ߗ����ι����iKV�᾽�����7ٴ ����Ny��Kay���MNur;.����Ou�	�HE�QPXd'�L
���}��A�Kz�e�rl�1]�t��G'�쏤~W0�:RqǮk��ѧ@Ι���Z�NС���c-qm�y[yxSY׼{��{&r�g�Da�[����k/�r)SD����v۸�C��qc�nUr�3�vK���=��7م�����Y��36u���|?P����QѱR��;�����#���S���{%mf�wW>���W�s�Z�g�V;����ӿ"���	�,_������$<m�}I=�O:��vp��ݿ���9�z��Υ��'�u����#0�@�:�x���vf�$�����W�^��wF����i����K���/����<9D�p�]�#L��uc��Lp�٥7�|�z�4H�}g�:릔��Z������q�{No�x���Ǽ�>���﷯���n�Z�1 ����Uҁ'�eL<�φF���u�U������H�|z���D��l���i����v�`�(�( yTA�"�g#��Xϵ�w��҄߯L�5~���3��]�]+[��-��<�U�"p����w�,Ê%��C�EĖ�H��^s��|�Ȼ�"g�u����M�ݴ��ڤ��7��]����\N�O�'Y�ʰ@n��1�:w����`fg������d'2>iN;�R!#]�Sދ̗}�+zpH�΄���:�=�z�ך;�c�OwU�s&��!��"��"��L�!�m�Tm�-��=Ck:�l�Vݞb����.p,���:�Y�����_F�+}�ќW^d���+�������uѷ+���Ƶ�d�	���ԉ�NO��5۸��K'Γb�	>��	G��y	�⤉�z�E�����q�3Q����J�z� �c�������^�>��tz��Q�h�����KyX/k���ߎ�{�����|�W����hڷ�i5��;C/�k�k�,���T}�dɨS����X��w�K���u{������o���W'F�Sʨ�^�i�W��G�����(�vf�id��d�WkC�����"zn�G1n��oOGrY�����j���!:��}���V\m`�_/eN�K�����0�ð3F�X��=�^���u�;,��`�:�N������/�47N������.r�9���W��Q(�L��:�Ga���j��EL���MxQ���#���Ϧ1���n�,[\DV�
K٧ޫ��Sy�#w�6/ڋ�����`Gs���3)��<��Ug�����w!�Cg�h��+�M�p��au�S4�BW��o�o£:rN��ܒz�eA<G]W�b��tY�~�>�>����%�q�~?��Yuo�4�1�6$�`��br�P�ΰD�����8s�\U(���������j��wV��o?���	��K %�f�49K��������^��%��p���i�ze-�n�	����Q�}wBd��u$�wi��5v���,ݗ|����H<�W�Ͻn����{�qnH=FX �/��׍+�ͧ�Qk�?{�H2�r�ӧ�o����޴8ds�S������3~0��rQ�GĕPe�/L����ܿF��s�����4��T��n�H��߯FG�י[Tt���HN��N����q{R*4H�S}��N�>U�G�2��qq���O��}��y�ti*=��q�&��w2�+�<O)�W�o���F���Eϝp7e��߃��n#Z5ߩ���w��wӵ���j�xD԰ೆ�����ѳ|f�d��$�gOI��)T�tj
_�����M_���z&f=��x��{4�KC�'O�;9�[�a�9��= �^��D�����T���P�{^17���b���e9�z�\Bo�h���7����d��Y=C&]^~B��襸��Lá�;���9Z�5�ޤ:��w��o�t-�:����X(V���Y>�0���_/��`��_��d��ƙ�]��Mm�L��|ҿ��ᐽU�rz��-�X:z=�B��R3~�
��z�����H�ӽCM�vZ�+���mmɧ7���WZ�ы5�(���r�A�]}N�[�e�������W0��T�ٺ��K��˛�"�9{&���L��캩5�<}�-D�D���w�2ȇ�{\�l.9{���e�Aor*Vs���npEo!tQ�����T������)�O׍A��b�~ɘ�PX�U���q��8��R�t�]I���y�~Hu��m��8�]���_���J�{�G&:�mkɶkkXJ}wJ̱���(�.��8�\�!
����w"�,v�1.���5�n/�sp��/:���T��[u"�\toiw�fR��:�#<w��L�mV���P����d�w���`x3'�4G�â6'�=���,е=KݓkW	��3�t�b�Te{���PB_	�3 ��L��F�b�^��s��!7r��®��������,Ռo�r�)���څ��qm�W]���U�Og\q1ՎXUf�o 
�F�֎>]�jC��������W̃��g-Rp�p'W�n	x�t�Yi��F�;i����!� w C0�2���.�L��fdoӅ���nG
~����n\���_v�GS�i�V1�.��3i�u�Ǉ��)v޻��I�hx	��@�]+2S�(^#N<T�J����0y��(������"\h���E�H�P���tך�k`��@j�<�8Y�*��a��]�\�֚�7�4m&�e+! YϬ�����x����;�CJ:}s��3��߄�'���<��)�|��j���� ����Kr�e�:ugks:���o�&=%Ӫ霔'I���0PS�5;kR��nb�b��̴yQ�����_,�c4C��G��7E�q��Z�9��F̸n���g�7吏\�9'��F!�MX���v�m�6P��;A^�*� ���-l�7�*i�L�nS��΂๴�T��;�^�x|l�հ�swVWP��'Y<d>�y�[��{-{6ik �#q#��\$�m�j�+�Ky}�X��gG0��wr��l}2�捼���eRj�o�M�R0(��̤u�N�̬d[�֚P�u"��/`r�J��%Ό�}Ԉ^�	,V�W�r�`Ҹdw���Ɋ
�}�V�׾��n�f���}
מא���6�4�F�,-����S�1Fp��;&nt��Ӯu�6�z �3���Hn\\��⽞ű�W����wæ4�f��m	m�_�[�^��f���R}���)ݬ[��\I}����U��y-o�m�po���#{8��Z��M:"��D�}ݬ�wr�@�r�D��x�6�V�FZup�d�f�5��P)�3�6���ά�\�<z���'�rI��!��A��1�u��-ξ�WJ�ío��v������.��������c�&H�̞��eF�W��w�Ktn�}��<3����P甚L�FUe�|��"�A"H:�P�HW��6D!���%tM�q�N�ҡ%��.��J�.��l2,DY��8����s:��B夎�8&�H�J"F"�!wPqE�����p�n��f��M�IQ%�����X��ɤy��/\tN�+�8�a(l�R�\�����9	Fq#I$S:�d�:��y;�R��t���N���RJ��p7p��]\(Q�/2Ye&[���'!Ut�D��P��g���H���]ۮ�3 ��<���N����ꖊXW�xb�\B��e��P�\�N���<I��i8���-�/*�f��j-iV�h{����tOT�0�!h�QY)HE�z#��������E\w�%�n��.{�X��dar�����y�u,�4���=�J��a�J�j.�,͑&B���2�i^zH����;�T�fIy�-3�D�J`� ��E��`�̝�b��>.�}\��`5�LQ6�"$+I��[8��8�b��w�n�g��t���Y3��d�wp4���Av��7�&�p�#2a~�&��9���Q~;����U^�3���s�;��^؝�R����͋�5;�+Mɿl�t��}�K������$��ٗ�y߀ϝS��&�!�Q�nU�ܿ7�=V_�W��[ư���k�t�̱�O�u׬�Ϫ]9�|��'�=UGŞ������H���^��j�"b1Q�S��|��@�C��G�k5ݴZ9<37�\�s�~�7��Xz�~�Jܶ{��C�>3|aụ�Y'���^�O'��c�ޠ=�ؼ�����t���>����<G޽���;����1�*nx+%#;��GZ�®Q�n5����I~�1�Z����/]T�uĖ��W���o�����n�z[��~�YlVV-V｢�Q;��Ԗ&u�n8�e����#��?+����#�Ӟ+��}����{�-�]JVo^�,a~�w#mM3,�Y�PB(�H�n��/ō�u�R[��v�蚿K�\=�Ie���x�����gt���q=q�����n�D���B�Kǻ �\Ud������2�R��C�c�V5�4��z�e�.�:�H;���P��8z�K2�e)�U�N���-u�B7ȸvt˨{;=1���8Uץ��F����}7��訒���3^��p���_&b������:%w���}����GJ�Zbf�l��Az#��G[j���+>#��/��u T)d��'��P�5u��'G�|�JU'ʏ��W�o>�S����E�����ϝ�	�~��iK'�%J� �Gh�~�C����ʃ�N�߶��=]�J�~�������y��cʰ=l����V�v՛�Q����ހp.#M��u��=E��.�q��onB~�Gz��)p��S�0<�̸��k+�}�44tJ~�_��]^>�b����.�SD��/��m��,�e5����=$�������G��*����Pw����g�>;;s>��:�5YgFDT��N���>ٯ	c��졈��U>|��@{;VB_����ֳ��U����x�g��M��ݳ0��6���=s� �m�نk/���+2T���i�/S������^��t��Ǔ£;*tݖO�����Eg���s�F���N���\�<��4��E�z_�=��������r�"2��~��^�٭����S�Tt�Ͼ��5�P�k�])�Y�n�q�{N}����7��j 1{�ڼOL�umlm]v��@ ��w\R�
[�}{H0�n^�}&�|������_w���3��,w�s19�.����y����w��Kv�9������k�AL�XxY�QvՔw�X��>fKD�g��"�뵀�AQ���Op�'M_��Շ|:��U)`��,	�yT;���>�{�bo��q���:+����wq��=W��.�|���FXJ��-�3]�x�EKIc�#� �z�}���O�so�������*�����S0��f�A*>�'�-��/G_(��
��r������*��}�CB�y���ƨ���&����~�TMC2YW ����ސ T�~71� �k3c��ɏN�z�Ǯ}���f���r4'�H�~�������Q�aIlTFG��a�^�jW�5�d,7�D��Tn)O���P�_��j6�m_��C���� 7�^�j�r�r03��*k�ϸFUt���d�}���K��W�e���9�_�~�g��;�9��n�2���u��=�h���7uC~��5�eMA�c���ꕧB��������w�����:.�3��v*��7ϕ�1���^���T'�ՔkK�8t2}��j�mhw5^Ӣ�/]Q��:������^W=%z9S�n�xd/W�F>�/�w�����Az�l�id�٘^��j�)��Ǿ�^���j.��V7�ٽ��HR�'.�a��X�ܜ+5��1�ۑp��B̴kK���䫫�a��s���8_`[�Ցc��8	0<����h�2���2��3�M��z������vA�,���J(!l奕Ԇ��ؒ��ъ�Mm���U��}���<��W������47N����R3�6G?$B��3y�/i7��Y��z�ڽ��S/Ľ�Gؼ��2������}>ntw���jML:zzg�1x����qr�cIvs�=P��]ў.�Q�������^������'*�.��������-�rtl[�OW�(z��3��]W�by�g�_��{S��t Ͼ�H+GA���[W��ݡ��r��+"=n���ٔT[�Q���}f��;�.��Gh�w�߮ܢ3��}�V&�w��;��cr7���q��3~0�G!U`[����y��V�z:�o��>�鑤���S�w�AI�G�י^Rp���HN�.a���D�`	�2TS�n�	��XO:�l����Q�޿+�>�eyߟ��{}R7��0�.z�๜Y�^����̟O :\�1-�|e����9֍F����#�8�ƕ��=~��7�*���){A���7�(�S:j[6zH�����WM�K���j��]s�&$��<=.^�c6�t�}��2�u7��e���&�l�ݷ�d:�݋nfn�8߂ΐ��X� ��1��#��&?fYI��I癹t�?!��WQ��DO#:��-b���PV�5ݭ����q��iA�6��ֺ���B�d����Y�>�FRݝޓ��?R���|G���/�`˙�h��Qf��}.{ƅ�:\mɡJT��}C�{f�R>���~Wtbן�Ѹ���;��	��Y�iOW�&A�����k��:z&*�p����5S����{�guxu�s���D7�}A����O)�#]̃���ЎVz֒=!���z*�u�w�e����4{����ȅ�#��CƖo���29X�W;���ef���ڔ�zC����pwj��#�����_��;m_�|���u��yϧ/xi�����:�͊;[��z%�e訄�$���t��^����k.��T��(�lˁ�μt����=~u�k��rZ=:x�}�;����,�[��gB�8qL��&x+�Y�T�s�N�R0X�~���-�C�g��p6�?�z��=��\wc�F3�gMO�c+�g���S�$f(�O����-Q�ժ���Շ���E�=(cr��}�<����R��d����#�*���)��c�z7��S�]9�YP}qM�h{ՁDo�|����}?[�s�q��u���a�+�����=WN�}�M��P����MR��M�pr���Y�>8�3Bn�n����v7;��ؓVi%K�j�`����_v���NT������+��ߎG�o�J�n�����)�n	����+e.��巏0�ޝ�l�ӯ�xA�� ��JT���_k���u�u��Kw�9�<����_]�F�]��œӦNfΖzG{��:��UB�SRX��x���^������q7�ZD��y|���퍮�ĸ7gY��H��}R3���2�� "�������_���F�����z�=~�n3���w������L�q��'��UxȨs%���L7c���+�h]g�1���"ßl�;�J��w�3��ʤj}^z����d�ꌁ.�H
Y=P&az�;3�1�ʍ�ɇq[9�ΎR�5��͖�oܩ�\Gy܏�U#�^u�}><�w&���5�Q'q�$�$�&I�#0���A�N�ݹL�gu��G?u�g����=� ����gw��k�+��z�Pw�N���̃���]@8��޿_q�-q%>��YP�"��#�rW�2;
�%5+�݊�=�?��T�cC�S�b�?��kå��k5��oo�$��'�i��vj�U��������3�+}U}�4������N���gC���:.n����}�������uL�|-_c�i�7-�|8�$^_A�;�Xw���S�������n,�թ��Λ�X[�5�ZZ�矍���G˨���/\�q�����Y��O�9�#�S�0m㰏h��Y�;��S.�7�,h�c���Jε�˫�}įr�n7�����Dz�Y�zhn�uo��T�E��fa���� ��tP�7W�ʯ֋�Ul�T���5�*1zߌ��o��r+��	�δ���{J-�"����,�O���y�������3�Ԫ��z@i��؇�ޢFz_�=����ȯZ	��;����5~,��EV6={�!��$񯤶AS"�k�^Z��������
�H�{N	�N�_q�K��{pz&���C����U)`��2���yT;���>׽V'�V����qI�{�_{Q�t�}�7��j�z��2�P@򯌰&��7e��пa�>��viޥ��˻-�g�P��p��:\}�UǷ���fQ,�B�C�F�Lצ��kglW����^gI�ٝ�	F�Z2}�la�u����M����鸏W�&���޻+|.�v���(�Rf:�����~���*�=E#�_3Q�Z�;���>�"}�Ӂ��lF��4J��Ln��w�Ϣh�9�dw���&_W��-�U���f�[U�)�ԁ�qy�{�/	����eȮ�����/��3��÷H"��Յܝ�y���	+��{r�1����;d�W,�WI�87��B�',���8�5t��HеD��whi��"�E]ɫG5��}��[@c,ү#Ĵm���,���9ڵܡ��u������2Ē��w?`���խ�E5>'�%���N
�}Z*�.��Q�R��s�\x���jA`�NtR���q���O�4o���Ǘb���4�SPrX����iУ�����>�ޏQo6I�F���h����{q���v�c�Ez��uP��ܝ��ﴲ}C&���oүe���v�xju�zѿJ(Nl�w����۽�^Y�=�z����B�{*p�d�%=���SdT���г�	�c��.=>�r5_���~gլ�~���άw�RMFM_���ڶ��;��g����a��G�����~%�����F;��I�Lcٮ���do��m����a��?�k�}�9'n�����Fz�__������y���PG������='��߀N����G���p�VG�\wd{-
�3�$�I=�(z�L�}S>����E��+����{�Eu��n��SJ2��h�h�xrX[-����yg�o�fQط$�,	ȱ��٨�VH����=T�qjJ�Ju���G��7V&���8g���1������a��~�������#߼o���%���en���V��p�yq%�U�'hp�iF;��!gNL���s_ك�G��M��
G�¦���Y�;�ݜ�Y&U��[�m�(�*�SD���=�<�uι�u��+	qq�r������_�>Y��52�[k�������v��2<ܨ�u��{��E�~�{^eo�Tt��=���t�-�>M����Q5w��1x��a7���n��=+��Q�޿+���yb�>G_�F��{��H�����7'hI|1�*�#��LM}�'�H�٣�"b[�㌴}��r:ј�o����M�$���Y��z^5���q�t�h+Ӏ3L��L��nKdq#"_�
���G�o�K�{��tN��L�2�vo��>����|�>D���Ӟ'��	��9��=4faz¬�hz�}B�MWM�{{�j�{���^�������Tc�/?Y�{���6��̓Q�z0��+�\�5�V.,׷/x:��mb�p޷O�dwW�\s���C~��o}A����O\*�C]̂�	�*�"�����r�h��1���fUn�R��ԯÅ��߆/Uy���x�Ͻׂx�V�mz�����FnCӲ~W�rܴ~y {V��!��sY~G>5/�ӑ�_���j�3�U{�Ϝ�f�F���_����>��Q;{����7�>N�g �t39U�I^'�ٗ��/B�p�ƿ��v�Kŗ���D�UWH`E�6#�U<�F%�ζ�l�F9�֓�C�&%�mU�;G��3g)rd��]}����˱�c4ʹ|���J�%�Rΰ���w:W�(�p�X��UҒ����ž����%�i�3��2I�S����n�+�Z�r��w��nWVn%us����9�g�=�p�-p+�s���`zʫ̗��,�ϴ,�.B��ӽX����^�vO�L�w�ׁ��~>�>��]Q��b1�s:v�'���bȊ�D�'=�gk/���~��aѕ2�����Ȏ>�"4����z��z}�ީ���o�W˲���ig�`��{5��y?t�����"��z�8��A}qM�h{Ձ}���;���ROs'��'��S1M�3sT��!^�rQ��>�3�*`\u�
�;��>�TOKw�9�<罖;���ü�5�Ju*�q�Ϣ3]HۅU��Q+!H�j$�0[�q�[/>�V9~U�cO9�觨cͺ�k/{�S�h�7��h�:�Ԍ����H,�(!}$\Ku��q��ƚ��0b��On���vϛ>�����Sf�u�w�L�{޸���UxȨs%���L7q����z�ƍ���Czw��ٝ4=j��lxχ�#|�G_ɫ�c����N2^}ꌁ0�Ԁ�?D�>g���/�:�p]�6�������VJ]7�ʡ�F�l�n}T�}�}��v1G���������`���1�cm�P�����1��\c`���6��l��c`������g����o��6m��1�cm�1�cm6m�`������6m��1�cm�a��o�l��c`���������c`����(+$�k+T5��60
 ��d��H�|s�E	@TU!$$IPTE$�JIQDU$*���E U
	IRQD%AH�@�T *��JH�U=W֒�I%)��EH����R��5Um�IH�IU $I)IJ$��D
E	V�*J�ԫ��@�IU.�AU]�DI(+�� �wI� *��B�
�J�����IUJ�B$**Kmh�PJ(��ʐ�UIV̀���U*�ER�)E$� �R<  vs�t��@F,ӡ��b[�I@�3Z���:�5������l�l�Բ�CdL+A���P��Z��h�bU*�D%%+�
���� �T.�j5-�Th6�T� L��5� -Q�:�
(��L  @�[�(  C:0 �  ��n8h � �;��:���B��vԑF�2�� � E�י[f+Zm����6�@ ιuH:�ekZ�L��	(6Z mf4�֦R�@���
(BR�E
�*S�  �z� 7��ڠ���QU+*m�цj�dEZL��@�)����Gt6�v�U��l�V��D�%*�)� �Rk/  ۙ�F��C���C��Uh�R�vك�+��:p��*ݷI���-�Q�SJkC�v�5Z[�aѶ�8n�Aȵ"��! �)P��  ��렪cc�(҃wh�فE����� ٭`A����a%t0��֚P�GN���P�;�aJ-��M��
D��������  {��P�X�F���*�ĥ�4�u��a�]P40;5������t%v��� ���-e�v���-f%"h�D�J�I'�  g 	�R�
�Z��
M��@W`�룭��5@ �]pZbv�M�
��u�l��m����:rh!��(��% �
!v�J�"<   lw��N�j*n�UTv�N n���]vРQ��樫S���@t�Ʃ���U6�m���C�&�[4�Z�����	!!B�� �T��  �[ZS[`�kB�l�-�����iJ4)���v�Z�wv�t&�5N�J:CX���,K��]kV��F)�hUr�T��̪J�L���$�%2�T�<#P��  S�A)U4��E?j4���� $�SI�U4� h��\�0H@D�o8MHR�%!{��r����}�o�?_}��=�_�B����	!I���HHd$�	'�IO�BH@�0��HH?v����|���k=����ْL�IJv���bm�vQ�Ih�y��H�uc9B��5��MĘOe'�aͰ�����[���8��Y���e���䫺�vJB���&�Ei�GQO[�B�!Ź��w��� ,�a������(�,cCm�U�����"M7e�Z�Q��V&}yr��J6��̙��3h�΀���ո�dci��-́b�,�ʻ����,N�(�CI�9F��4���j�-rՊ��ݡz�V)�Թ����-��m�a�n�i� ܵ���b� �
� ^^�-������1ՃQ^e%�V�K�+q)|�6VTȎ\ٲ�7�V�
_�4��F��; ^�Y�fɕ ��q��M�(,k`�+��|ིt5�DlK��U�|�m��aV8�5�\ m���j׮�$�l�2�Ȭԕ
�Z
�����PT��NI�ޭ����FV�$��Z`��˨�J��(7�t֜uz��i/�Y�����_#�Ez��3k�&�h�
sLOQ7O5F4맘����N]�57�yfh*�E��B�vh����e��l�o.�1�4���v�dQ�un8���X�.��Z��һx�����]�#]���ʖ�M���7m��MU�2�$���/1�,B�0��c� ��,*�m�¤�c���L�w�;�V/CU�������.@�N�z3i�0��R����r���ջ%���&��"�[��B=kYbm�$1z�[�����p%,-�6���;sK~�u��2���6��ķNd`Z���~�����L��c6r����J�m͉��atZ-��̡�:�hi��՜����ڶ�'�2a�Y�2�U�r�g4����SB��]�m�Z��wj�qH�6���*V�jj���$���ͦ��ef[�X��dZ`ق�+�O0�Da�Z�Z�u〜X �3p�v��۫sI��bZ��`ې�t쉺��6SwP�$&2n��O+	U5��uv.�ŉe1�IG��j�e��wi-8-H%�F�;[u��Z,]jk��ڀ�/�6h�i�X���Ud��ZG@�`9q�YF�6)�����8Y�F�-
�4)g*ޒ�{\ٙ���;ԘI�}�D@���K��G�nQXO�ú(]R�U
&�bR�
x�;O�J��L��R�n�wR)cRء�(SòɏE-�4�X�M崊܎���F���Ѻmͦ�hX/)�̡+,c����؄I��Rtݶ%�5X�b�1�Ո̺l˽
�� �B�LӺ�:��ul�����+7iӴ�ź�z�]�Ă���L��c>ƻ��͎�w[Q���\�:�� �&�.ic�JH�����;��cu��MT֎۸�� �Y�Wre�:�`YH����-�pm*�(�r�fmFtQYF���?d5>I���O� ����Rk+e^o۴�Y��Qˠ5; ��{C%d�iܽ�2R��	��ʊJ9jV�^*ݙ���R�݁�N]/��F�Z-*����-�[�X�lش����7y�ݻ�d6@#]K�Al"ֳ�C"+�S��f�W��L#R�J�	���ۘu��)d�/R�d����I2���ݼ G(L�f]�-X`�7e0=���s 7J�R�l���)ey�	��WN���;�ˋ��:�ɼoC���օDq��5�����Ef�����12�����6��,mL����,fk����m�=
!VeK�І�]��l�Q����ej6,�Q���B���T����D;k+\�$E����ZI�XM.�y-�+�3L���f���:���$]�b�#�@6Z�X���4�1 f�ߞ���whc����9��f�f�'NE ��x`WP"���Ѭ����n�
*�Y�f�d(��8���i�Kq�zN�Y��wq$��ݲM�ۙ���Q�5[�x���f�r^��$�ë��
���<��m]���U�`��d�������� �rҒn���m���k��Lb!n���>��b�q#%nƝ児�r���y���M�u�i7�j��׃E@o�JKC�n����v�$�\�6���j"�X�r�L#�W�)�������pb��)�m�U������{���!h9��M��x���58�㵊���̩tͬ�1c�x%�ݙf�[i�ɻ(MC1�!H��L��`^���y��/6m�j���enj��\0�	�(r�kO7TV�wi�#�����j�3�\ԥ�;@�AV���Z��[�,���$�����f(��B�?Z���Q�v�4Y�Lyf���J�đtf��.˽�u���v�\d����0ވ���ٻZ�ih@�Ӷ�����dJ�GNh���cI�G���:���f2��V�lty:A�s&r�osCwk�Z0�Z)eh��K2n2�З�q1��k0hW7Xڢ]mc���`P��(�fLzų��w��j�X�c��տ���[u�2�Ђ�lV�F�x�
��Mn��mM�ͩ1�Y�6��C�ٗF�j�J�*��#w���P�n����Z4.��_Y���j .n�c�ph_+�/lG���,7&,�	d�j��sr��5���̪T���d+y��Ld��2 ten1�T6�˨��/�X�Ţ��τbj�m�"��]�3�5���B�l�ʆm�������%�L���A�w������.X0ޫ
`����f!�]�����:�V,���	�E���:�@Z��^�ĬjAhJɳ�$!b=j���D��<OD�#2�b�f�U�}n�i{[�
�c7k�e�%�0��Sm���6��U�5b0Bk���4&G3s&R&�	�բź���n%f��ն��]dە&�S�W�
[�h^��5�-��
*���s,-`b%�:�����YYy+NK����	�X�������R�2l��l!u-�*ͺ	[�Ɗr�T��jȘ�.��D�Hm�uhއl�ACm��ZV��Me�t
p�9^
u"���æ(��ژ���X��aح;Ck1|�*���Rںѿf�w2�I�ͭE�Iߤs]̄n�fa�����O[f��0���Yh�	n(�Z���-7@����Zh�ۧ��L�U���#x�y�]�g(�/#�hu/B=�j�:��N���XR�|3Yn��W�yg%��n*,��lU�h%hDEjܭ�A �U���kՒ�|�h|�츮��!�ǁ�.�.q ��NX��ʹv=Su�����*�xF ��z�f*0\�[`��V��[�7r���!Ӽ�)�oD�F��r#�`���On�˕�)��D�U���h�]�̡!p�.��J��t,Sn�6�hϯlF���3S\L7*<ur�����{h�c-�Y�	Z��M�0L�vP�[�M8㦩i�1�bhl��M�W���)�w5U�h8�9���k�H��u*P�+/ZԴނ�FWB[�U%�gi��ˬt�-#@t�KAb��7C��^��ef"b�a�3��f;�[��сh�4]k�Eګ9LM��M��M%�64+{��pT�7����ӹ���d�D�,^Is��nُ��2��r�A2�=���x�JBc���ƀ,�6��U#-�6�E&~�VjZК���oR�=�Q�Y�J-9���p�D��(l��0N�m	�N�E��em��5�wQ�d�k*��U�Բ���g2�l%��P͌}/F�� EtM�`h љ�=�[�O!��U �QAKM�ǣJ�&�WH����qP�,�ݰ��4��t�If3X�-���q���gL��Šw.�;#��P:�T�9�#J���xk�4� +G0d��둂�"��n]�ɗi�u���va�kKXN�-�Nf��-R' l�+��^�wL/1�;I�N�2�Q��D���e�A�lP�Z�RHK����U�����b�����^�A�;qi�u��A[$*�0[� ��km'�7���j�G����u�on-Xɴ)b� �4�m�v��Y�j��3w�mX�Q˥ y4����#��q���ؒG0h��qj�h���|����4fJ��1�zH&����E��`�e�o&V
֫~>Q4���-:�gn:Y�����N�t�0�Xa�5"9������,.�Y��xX���h�˛�,z�55^$V�V���؅*֟�VnU�R��L�vx���8C�>{f�,Vh6����gU5yDf�v�n�;kn�N����̌�.���3죥mK[�5Oz�a���okfk`&�ƕc+l�%� �$R��U�����:Q�i`�#��0������3����6�!�m�NӋt���(�ܠ%*H��`��QJ#v/�������Q�tbfL{k5,Z�U�m��!	����b9�嘋�-��]��.��Z��t�j&Q�SKX�Si�5Iy�L�3m��59�%��@Vq�P��ܡN����`'
B���P�ϖ�ف��:�<.['T��jM��P�:f���ľc�k �/Dlj��c:���ܱ��m#��˄�y�RDL�k�4���w��C�ʲ�id!u�F'u��p4�Y�1]aOp�8N�*R��+]:�c~N�C��60�޶���A[%�3�{�)�Gco*ʕ�M�Nܛu���^�&�è���c��V
��㔦Y�!��ldڷ�;��wM�#��ܻ.e�֞R#K�P�hcԙ�Y���-��b�we��2G�)���Y�
��f�O������+����*F)�٦�Ы�t�m�tZ�1=)��L�u� 2m\&��i�D9��M͂�]-�SD)�@�f�H�h	Ǩm�C֭�U����ĴQʸd�\L�:�)^���V2��`U�����RRVV
a���M�΅j��v�n1�l�j]$.��	�s��2ŕ��X5�3��:q�(�Y� �;N�Fp%t2n��Z;ߕز.��(�Ux���[bX�͈7b����ک;P��NH��@L�CV)�3]�ҋ��8�;b�؛�7b�ԩa�c#n��Ƶ�*Ȍ:�X،�p�HX�m���j+NS���)�.�ͺ��N��yJ�!>(���6e��f�֜L�fjiP��C+nlV���]��Vt�4��r�Ш���v(���!�P!Y����q"5G�\��N�ݧm�ܺ�$_kM��k�iȆ�#�!�F�/H��U��f9�Wb��VЄh��W�ʷb�H��B	�d�Sd��~�te-[Z[$�{.lB+s(hF �0V�n��VZ/r	��ٯ(�JVQ�5+4j-=z�f%{���P�� "��e	b��� �a�0��_�v�#R��f����u֋5R��mӒ��'4�e������`2�;��j�&fi[I�k[M�rⶰ����`�E�ǚ4JѨQ��AǊ�T�
i*�Z�(p9���5�V�;�72���B1X���q�hXMn��I�PV��GTHE������9`ެ��I�.R�%YLe��+h����t�p�l���f�[�c��>�ȅ^^;jæt�,8���݅��1�Yt!n=0*�c6��a=R�1�I��@h��5z-��j*K4��oVL��3����δ
V�]&���i���5���� y����A!̼�	&X�n�]����)��`�֚V�J�6)��
�V��ؓ"�ۧbV`hS@0�O��L�+7S5���3B�����:{����iO�����X-�0ԫ�Zx�삲]�R�E������m7O)�R��ܺ���ܢ�p�AbҜ.����*�6�-�D����fP!f�d�iV���[Zr��r�^.�7��F�������e
35���\r�eu��j�w�Km�k�̩B�4�&w5֯�!MvmhU{u�r�\��]�s%M�U0��̖
���7s`�Me�:��2��+q��,g���T��!V�M3v�K�YZ���"��iV,���&Z��i���z�)���f\��5b��5Z�b��7J�r�J��SȜ�k&��)���|���5`��IZ�Iǡ=�1��%]n��,���E�K�E�@2�4!�����m�4d��M����+/]k�I˵K
�so`�p�Cup�w��c5{��O��)sa�^�7�kp�;�����c"؍J��'jX��$Ƴ
���mk��&TrE���ǚ�c7r��V�v1��.�L9�P�r��9��Eݫ,�Zރ��B7u�H���6�)�V�
�8&J����
¶\o9��jel��Dv�j�۷! P�54������s#%췍��֪w��u�e�Ʊ͂<C�Y��Z�=���3+l1>2
�q�:��C���\ ;f��8���[W��6�l�l�� *pH����j��qk�
^�#Y��4��X�A�n�e1�Q�.�%w�Y$��&m�o��j��Ղӧ����fV�jhCҰ�Y��]�L��5)��V�5��B�=����	�����hR{���مM�I�4C(kL��.�5G.%X���.�[�`�t!�i]��ocf��el �Y�A��M]P�D\ܦΘs#��m�� qJ���à���YCL�{.�3X溇-�Z�Cy�6`�e��rњ�������0KV�[�.�(��4mT�Kwyy/)c���e&�a�,�`*Ǹ��i���vA��š�.��h���὎�9��da�0*(I��#��#[9���1�푌V:Y��:n��է�z��_��swg8K^���=�XC��������YP�o�R��
�,:Է�:�X��;�2�F�#;;�!��R���{�:�iC�/��֐�s7r��h7ܓ���\Y�:�sṥu6w@�2���� �ŵ�v�ug%;T�`�\����s�׵�2�J��Sa����'}�wTv�o)`��I�WP}�(+}��ƥ1u̙	��AO2j���'����qi��[C,�!lX��0�J�'/R��sT&�C;{�'����N���D��s�=D�\���U�#%�s>xh�87��%�L��BZy�Zw�b��M�c��sz��ȶ���Ҧ�a��ˠ(�ƻ*ب��n��Z����J�]���e�u��+��\��G`u��Q�wN��T�6�Q��A��\z1�7��.���w�+V#�{�����;o�������ya,�Z�k�䐛��"��p7���W>z3�f|5]>�U��L��w>2j�WvތB�j��K�-Ez�kIS��A�tW0��z��C4-4�gmn�p�;ՙ�guٕn	�R��q�滺��u%0Y���b�n�SB�������Jz�i��~��!j��b|����V��qb��uL�ۭP��ܞ��� �D���Q'��=X��^��k>��5g}ԛ��*�o`b�3�#cS5�2W
�w��+��F�F/�m��Pk�:�Xe

OtY��vvf'R��I���w]�V���G���e8Ou�Ҝ��F���.�:�+��:�N���d��_]��ik}����л9��Tba�I���rp���:���0x��N�о.kܦ�je���$]i�a7y^���UT��5��:��K�5坍�#���r[Ss�x%�t�_�Ky!���1Ж6���k!�R��xOe�EWs���u��!h�j[xμS*1�i�;WX���Sm���h���B�I\I���,��	vPŵ�`Ƕ�[[Ɨp���aÛ�sܰ�
�	��V)�������s���y�TŮ���
 �k2��b�]1��YK�4o;�kMG�Zc;Js��M��95��^�N�^���~��_lm�G@qX�����7��-b�9>�]���7FY=��w�dhW����11�ƃfv�	b؁�p�[��/x��5u�GCwO(�o 7S�Z�./*8A����i�P��cMbC���>6���w`��+�;�����_kOGݫ*0#KNYBt��_-�x���K��ѽ]ZML�{2����Ac�6%n�9������ԋx�XS�R��}�h�d��sU��{��WN�q�/����{]�9��Q�	�ʷǀ�cͷ�ov�ۋgN\���q>	�j	���wR��յmmC���S%�×\;nͥ��ޖ9��[V���f�&�P��s���r��K%�%o:�ׯx�R��e�W��Dq���m;��H.���ˮښl=x�7W%a�]m�k��������`lVrf]"Ɵ��T7(�p�fރ�!��0"��K�J�u%벬Fڸ�(x�ӧܤ�����=>��e0ǽ2���6n��>���y��L��Y5�m�Ζ%#1��GM 
�g-��u	I�w��n�o15_9F�'�k�O˽ʁ� C�Y-\I�v�Яq����԰�̮��'����Ft�؝�N�YŲ�ʕr<��,�V���гu�r�Ӯtޙڑ[}��x�W*	�lMu�3���y[B�2�'��ߺ�'�6{o���9Ɉ_`;p�'���Vʛ����;@f��P�lO&�h��۴�K�V\q�� �45��W�|̫��JWRV�!M\���ȃ�H���.���5)��G�I7���W�e!� ��.��m�g���P��)�+v���G���ι���lN��I1����EgH]���{��hQ»o�x��Q�NI�V�2�����[�f<�bC��]�w��bI��|�M����	�B��ϬI[�̞�@�a�6�s�Vc��+>�TǠص@�a��[�ot$���V���v�B-���s�	4�Z��ꂃ��H��[�t�N�_wy;c=���S"x�p����T�Zc��5�q�:�\�sM(����t�g E-� ��޵�@a i�tXU�ԯu%��|�ގ�����7���7��KEeYI�]l1˴ ��2��Nj���r�/:�Er����R6J{��f�?����ֱ�G H1��d�)aa}�|�α{+^#��HB �M���o��w}x�R�Dz��l��V�ӡz���C�1bؾwn���͙�]�U���҃��^-{��^�Y��2�أ�����v�˻�%�ڱ+.P�=��NΞ���dG9OoK�S���9ݼ�aU��R%�&�W+�r�9��Y�u>���DP�O�n_ºs��	ޜ*�P�G2�ܳY�`>Јv�Ό<R��6;�#�3�ޥ�uڜ����J냆o,�����lr���Us�Ժ�����y����	��ֺ_Z8�.�[Lֻ͕E��Y%0�U�k�s�&P�pԚ�g�����%ʝ�c=gۃ�V�ڝ]W��"�����L�g����ύ��]�G�����R���g;�ܠ��Sb����ü�qxkF��kU徬S�М/i�.�D,
��Nt�'���?nXD5e��s��]@*6�c�q޴���}��nk	D��p�V��JH�]Do9�Y]�&jJ�D�N
3׋.�>xӖR����	T`��F�1�)\�����X�I�؊�����f�KA4[޻CP]Ö�Ŝ2�`�(=�������K(��F�_�wM2��Db��bU�(6��@f<8�;�{�<ݑ	ٓ`̥�VPf�8�m��]Y:�rq��ԡÊ͑e�m#���ɽ]��Ϡ9�9v��9�����aڦ�=%̷�+cx74�Ę=���لٔwv&��N.y�r����,�L�S�R.��4����A)�z�{�f]78�']�6tҶw]@8��V��H��&�])C\!il�)����+�+
+�P��(٬+�+̜�K
�ە��	�����F���d0/!�)�k�)�`: ֮�zv��i;|�l�D�W�ÀO��ob�:Wj��3�d��vV���� s��	hs;Z���|ʴ� �ޡ�R}g�)}�9ͥ��]��QXૢY���}���G}�νq�܅1]@�VS6�"�m���љ���s}*�,p���v����s�֒�B�L|>Պ�̚��V�h�b�[|c�i��j���wM<moG��_^�Ŝ-;�B�9ܫK�oWT�oa`����E����0��Q�$8�k[U�#��l�
*�TWx3~a�B�6*�7+��퍘ʰ"9Y)�T��}v�^F�G�CX���6�h�WW��D���Ѧ�k���[��ne�V��ل�]�o<�\���=	�#��VA��<P�nf�A�̃.AD��jaVn�0��wCN�m�4��z�R�fG`�5��tц��pP�'�؆�-�9r��j|�j�wu*ܻ�h�;����6�N�C拓)g2i���][@��\}XG^G{���ʵ�Ω�m�n�sv[hʕ�`���%5['��Ď��t�:��>����8��.�q�{V��X]��·���l��FI�漋�t�.KU{
��fX�kM�Q���]�U�ܷmJ�MZ�N:�X���'C�}u�Ճ[K���J���ƐV�3�3��+ޏEbP�I__D���y}{�o�CC���u��3O�
��8�.�tA�F�v`ӝ�5׋�5[��a���{����uY{��^'Yj o�qƪ�ƶ�`�MN������q[��S�A��$�] q9�ܼgm�m*u�S[#j���䊮���4G��՗V�v
��,�-�&�!�-bnʛZ{�����oc�ַ���`.yk+ZH��x2�՘�.WH�ﻰW+�;q.u��~�. 0�f9�ڬ����)��B��.;˓����T��*���峏t���u�&�nn�u��q���va�)��9������O���1so�z��gn����_Ò�i����4b�4ʆpg��H�m��'n��T/2:�v�so1lݶb�4W�#I�`̤5�ɔ��[v�uG[k��.m�U%ީ� �������5�n7CC/[L�ر�*�ܫ��@L�b����@^t��3Zq>�n<�����I39�[�a=�rnڢ���(^��Y�'frG���m�5�w���B�8n%��j�� u(^�K�X*�(�ht�K=�]l>*��᭿����@׻ݚ��*�α����ً����)��_��z�gܶTϺ�TWJ���dj����;#���QB�����Z�qSu�%�����v�F�|�w
�b໰�P�Zyt�79].�!u��(�t݁�&E����)݅P����+^u����b��h�AaWj�o|÷(hoaۂ5fҥV� mj
���7DJ��E�-v/�K��ܴ{�C�FŴ�bb»��w.MeJs����uy1��w�1
�ɚ`=��}��������G)�"=t�����W�K�&7�zm��t���u�G��:�.�ͨ�Z]a��f�,�.��U@�pS�ǶV!�bX�^��׶�ʇ�vgE��C]e��n��0Z�--���!�-��;{��S���������I�Iٛ�)9���u�T}�[n�V�V�y\2"�i2,�͉S=�� םu��<2��(9K�J9�Txh	�����lr��>��4{N���u݈����v�o����L69��t/�E	����:���������w��aA����,��晝����XmsSR3`���U<+-�&�t�uг�v-��b����t�@�]
��]�0�R,'�m�|��Ty�5%a�S�(�i���[���v�V&sš��%��b�:T#0S��IW]3a-P�^��:��+�������xn�1j��[��_×�eK໊�&�9[� ����\hݧ���q�0E[X�agZ���{�W-]�ve�Ϋ�&Q3���kw�ҙ�@Fe�M�w܉�̃o�&��N�Y	;Һ�Tֶx�����v�W,]%��4f�X�9OQ�I�[s{ �+y���m㡤��5i�_F.���+ԮG^�F�z��\0�N�u&��n�A�l�k;f�����3����2e_f>��1�ʱ�\����^::4r[�����菺q�V
�]vVij���u�8����T�(ݛ���0�e3�CD=BJ-Wfv�-�:-%e���&�(�R�mX�<F�V����.|���.��<c�y­A�m���d���QU՗�i�E�X���}�+����#�EP����Ե��iMn������V�����ԕ��"=��9�l� ���De��A�7�%�\b��r�A��?4�~j��i[˱Rq[c�%������{k5hKk�Jm�t�y�1�Ku��ٹ��u.�f2�.݋;B�Xa�Rp�Rv�%Җ~m+#'
����6�u�UN��j��oO�q����۟Cf�����R� b��nLܻ��;3�fŝ�Кmn�`�*.�
c���3.�WD�a�2�0fc\�ut\��Ww8�U2�j��q��9�����v��cD����ۡ�y+� <�>k�\��]ԩ�F�vPjVh�A�(u+�.��ԯ��׺�]gL�Y�Ne���	�wr,�¥�։�S؇]�tN�k��c"�|zGt��B�p�[]��]\�Mrd���ص�U4�f���^c�����[G k8���dTU�q4�Y�6���X<@Ӹ�ڀN�
���w�����
[F�5aC�v���kl�FI2�J2}���-�x#�NT�J���n��+lɺ;n�l[=u�A�>1Jj�� ���%4#�Ti6����˼�`]wA�YT�����p�]��:�Ώ�ii���1��,j��)a�t���^�0\r�i��^*,vf �!��x�����&&�p8��՜�S��q���j�j�0V���:��$�(��.�б�jҥl�8=��Q���H����W�xX�U����)p<�lGV�i����/��8��N�J��W�K��.^��b�|�ެ'DP�n�+Y�U,(�,���M�T>(��WW�\��*��o�U{L��]��yV;[O��AeJ��9�t���YZ6��Y\���P��%�z�������Vࢡ��լ{R��t˗f���E] �U�&3��8�뮮�0\��E��m�H� �mE�,���+0�֟vo(+����V�.n}k��ӁqVz�!�XՆ�����y�����S3��/�����;#Z4f�)�=^���}]>��e-��MŲ�G���YJY�lQ���S��ty����}��Kɏ}p�Azhbu}������M��SV`[ܺ0����w�g������+W�Lp隻�]j�ðN)Q-�2���+ˋ��AWG�l;mh�v��o#��!��B�ܺ�0�];��rmӒ���3�i�t�;��8���u1\ټ�	����=��ʥ�^�ҝN�(�R��GH�o}x+;T��p�k��7�'��mP��i�Ky�ٚ��qp�6iPý\��xU�t;6���vi6�t�:�i��3m}�
0�E;
M�-an� E��l�����3�n_v�ۑ��"��F�8z+��6�RF��]�2nԝ��}�i��6>���)�EY����`�������Y�䃳 �͆��=�֔���en"��X.���am�]A��T��b�����o��׭�1;�6�z������ ��!l ����$�y������T[B��_��A.v�Eګ2�ot�{��o���0�f�Ԕ��=�z��Vw\]���f��L�Wض��>a��$��b׹����S�����Z�v*�PEJ�Sc��S��O �Wk�'�y�A��>��޷�H�U���[p�7��\o��($h�V��Q.j��_���S���;x"ѯHm���.��e3�c偛8����wu��E04�߳/��<��V�1��S.4ff8�	��I�*�lMB@pi��&��ң4TB�Q���ZMC��;r��n`�طi�ңq2x+v�$�������,ٴ����u���C��#r���;�yJ�IoM�2p�{��4�Y��J�r�^r���Z��2ˊ.=mH�y%ޅ�L�z�m_}����0�����䆕��-���Ѵe&�5�i�}�헫�2\I�w��8�Du:�5�]�+-Z�]u��y׸�ἇC�g�����e]q-�f�T�� ���Jvh�
�cf���WM���*�CY5�C]�o���[nk�S�ʂ��Eir�����GlQ�ʚ/�Bܠo��H#�4�Y�S�>
�:������,Il�d�n������3E���,|�+�.���`�Ů���^%mm��S��b�۷Y���+wi.Z{�F�ӖkJ���J�EŔ#�{�)b���5���[6[���A��H&в��"��^���T!�T�╬�R�QQpũ7�s4L�r��ngJ#P����r��3_\�EW
 ��c�'���r��)�W�H��P��GJ��Y;���٩��W�˻i��}�Ty�����3(#�������:�[�yH�}��o5j�����F
�7� �}���sV�>t\��Ԍ?�'$ZBf�c��{Hn6�d�:����LJ�BU�P(+f�μ��]�7��@�� �ݺ�<��+P�y�۸��]��'Bd�\�i�	���݁���ъ�>A�5�#ٚ��WLٲ��&Y�s�^2ohл�Oz�!�� $�{\�چ�̌Nt�8�=��\v�a�;w[ǝO���I�+��cggqP8 �f}��E�Yu�M���{�s��y���n�/x�Y��|>����y+ ��Iȣ�+���h�!D�WޛJ����uA;��� ��A�)�e�ʙ
B��y����\��i��P4�#Shvd�ݤ���Ҩ��Ff* H�0����ً���Y��]'��G��r9�\K�@��h5�c>�g�>�N�r�)7oy^GӁV9�%��#��O�gT4���7V�	�Ą�҄f�\��nu	�]k�A�Vz;[�ϳ�st��{�����^�Y�|�c\��L]$�]:"6qt�H��zv�V:��.7z���V�Վ����`ꕏ����D�M)6r ��U����%�m��f�q�z�^�gI	<	U�@M�Y�#����y�U����t) �ʠ(V���\�\j^��-8�r�1��Z*�
�n���Uݞ�yPb�G�Ea��R�,��mM���V��w+DC�/2��U��¶ D�����k%m�Y���>k�P@��$xe<Ș��H�E{,P�r.��eMǙ�E��e5ϳ^Mv���*�sW݂���b���=	�c*�Ԃf�x�W7k���oC����-j�ƣ|����^�鵳q
k/���M!�-ڃ뻚��A�U�B�9��n�a5�O�)�{3B�iֶ��ldЩh1����/erw�-|����<{��H��M��W^c�]Ho-�Fmv��4Y�
�8�k��=�-�X��U�x;u7t���q�c�&m��^ ��\;��U]�5�y՞�sX�+�v6�h[����n��t��|��[�
��'�Xn��P@�n��<ژ��_N!c���k*�b5���:\h��c���ܸov�iᖍ��>F��)���S���t�.t ���8�v鲲�3�Xm�z�Z��.��)%]����r�:ôN��;zR�lu
?y��&|Y����T�-�2��5[� |�]�� �!���V��_�N=��Y�����v5��4����h�a�)�u`n8ڣ�i��볶�`�������3�^�B��@�u�#O:vT�l�<�o	���۬q]�+� ��]5���Te��ZUK�9�'��v��m�f�=w���(�#A�ЩFi3��g2k�03�F�`�]Rbٛ���yL�M�F�۵Ru4]�U���y�������7�P"K��+�d����@>���r���͠�~��v�2�U�S�m8�Eaf�k�7iһ�����Ua3m`DԐ��4�ʀm��d[�G+�mC/&ZT�\�#�iT"۱P�k!�;4������Vu�V�F�Ѷk9=����D�C�}����S9?��s5c����g��q���a�]��<����`��a-\�]@K[��s��J����\f��g�M�Y���p/��Vf���[ʞaY�T鴅={��Wn�H���P�}�`��x9���,�-���-]X'X��-�ĳ ���e����)�GB�����_]��=���=�)�{��\o��\(e�m�@X�J�us��oN�e��⛣�j��J{���
�:����n�9�����ƋÙts+��@�X�B ���%7�7��FQ�)Z�lN��E�.��	%@�x�3}V�Xz���,���j�Ӳ�u[�`�\�[��A���ȧh0�;�wRh�����^�{���+j�T�Wg�̭���Z�)��=�@�JU�Y�d���hm]�h�˫P���{-�@�Yp���j���7b����x;��m���fA�f���r��W�,+@�5�I �*DC�����l��PI��m`N���f�Vy�\�:�m<*�j>[U�3��ͽ��t*��ЗP���ϕv[�s[����κΏ8�� �0gD{���3WD�ғ������mk&�.cxgG��
[k&I]�9N�n�aY�}���)Jh��tO��۱�����o�=��q�"�;DD�V�W ݒNX����A�'�7�]u�A`��O�7�q��`���u��q�n� v��#R�l^1SQ-.�[s��CVq.�����(3�h�6U�;�x&�>�>u��0Rھ��7��ܾ��Q�����{6��K0;tx���ې&�K�fh�mg����Eec������͂����j�K,�%�"^}&Ю�G�� ��v.c�
�����%�wad*)N
/rv���Uá\&a�;$��A�����		P��N�R��3��Ia("��b4�!�gx��}b�,eu-W8�e�Y�cW�eR��(O2M���_f�ɳY�n�K��s:�7�̝M��\.Y�:K��᜺�����f.Gs�u��.�ѐ�h�hR������jӊuKR,�]�Pq�kE/x8^�Ӵ :�|7 �ல�J�	�M$\Y���6��������3VWt��r�'���+a�w��e�ś3c-<ܶ���3�F�inu���
���K���&,���Aۛd5]l�C@�Br½��kCv�j��z7|@�Y���q.k������(���r�wjط�T�\�C�R�-��Pcr��9RTU[��V$8aFt�Q�/X7���	Іj�S ������]R(�n�=�VCH6�h'��u0�]�[�F�wxG�-�2l�6�l�i����=�J�eov�hC�%
���t�䵥�I|x���f�bj� �P�44L�䕫R�^��|�E{�c��5�̢�ɰ��v�6�y����	R����
�Kwf�`0�C��F�í�5m�G:�;�	^�,�Ѝl��Q\A�{˟%%vVG�mI(�͋�@��B����G��}�3�ʛ��h�jל��R�9��vd7�T߄9׎C}�wX
��j�v1Յ�ׯ��WN�D4�'ܵ��E�n�@���y"�t�r��K	M2�pQf� �e���c��ɹ@�F���]�س�+w�,l��o�G�E�m�knP�A�!G�O�a$0gM��%\dol��7� jj�Cv�C�s(j��c�����,��'{[n�����=R=�S�h�U�[�/n�Bi� o~WF��l�J��=�d|@x�eɔև!�=Z���]ʜ9�iA���1b��f
���IU��+x���%�`�tᛉ��co��y�΀��gQ�,#/�n�r�rWkq�u� �;��1e���s�^��Җ�f�2�S �����Vo�lޱu��3/~1�`Y(Q�mg,7��7z�G�i�=#�Mv.\/_TnJ��p|E��c�W^�%V-�ƳVs���ّsW_R�$�0�heiL�t�������4�܏Y�,%]���fznc�m��\�*�T�q��~|1��X����e���	�=��
�RT�t�6���W�Y �E�5ӛJJ�/Y��rjm�;Tr6i�7&��H��n�k�A�
!�+v�.ju-��]�d����?)��X�_��p�������]�@ޖ����g���1�d/{��[�6
��Ŕ�8��C�q<tiTˡB�X�Us�;�H�6
�uY�L��#d*�y���g׮���nJ(��v*ʚDv��{j�O��M0F�kk"n�EkKkľ�Un��vH�W�̱[��#X��hD��m����8�ocT����!�YW[�`x��iބwE���Gή�[�(���m_h�n+8�Շ�U��٢�h�=3�,Z�n��\�n�RW!P1��V�}�s)���MՅ,��+;�&��>���YF=��(J��]y�H�)`�|'hַF}�!�fb	�]�i���nCP���]�	Χ6��s�cw�n��)�a������pv鷶z�IV����p��5|��1s����	�[ǝ�Q�]��	� +kAO�Yt���Yת�'f:cؼ�m1؃ҝ
�{}��S&���0Ҵ.�Wx�٦�I��q��K-`�c
HZ����z��#2W8i'X��FŊ	]�P�X�6f��9ۼ{w�O29�8OG�+�׀;��J���T��Z�S�tV��]�yLv��Ү�t���;Kv����K���qN�"V��56�����Y�9�]�oA��3c�r7�v��(���h�$S��UsvfZ��]��J�NF5���iX����[���)�/�֞�K����[���ĸP���f�6;d����]�.lfK@f��}�D��h�k/9/�����g���w���*p'��;5ǜQ'j	�ܬ��rǕU��w-�d�v���9�A��,������I.���Ң�\#E���ηѱ;3����u��9��I��\vj�#L{���y�>X�s#���7qZ���XV.�*�T�m�SOj���E�m�Q���D9���ɗž�r�G�����@N�#aw�Vp�� 4�t�7eƵn���ʫ��Y9[�����>���j���*�;��ҁB/{0b����������R"�=զ�j� ��3�|�Ԝ�u/w���c�%#n�g*!v�/{IΩ�u�W$6�Pcw������ ���]��@{,�P��ʽ��GS��k<7�kkq3�f۷(�"G�F�����v�ұh�H�gJUXe]�4���kM���NSFgգ~ǃ85��s�E��3S��D���Zy��Ɖ�zu��Ƈ[7���8&�*d�!H�x�{��y�3SVz�q�2�:��fr��9i�WIM��e�c���Cj�w
�k���6	�7� ow+-� N�
fb��:��Bg)X�Ri��A�Z�&=��ui�7�t;��.�:�N�xWQ�%mΜ:Q�U;��#U`N�y�Qnf�5���G��,�.*����#�rֈ�'V�ڝR���J:t6�))��|��43�ӽи9�4nw�n�sT���_�<��v�KHx�Nć-�/���K<�8�PKMQ�����C	�9�A�d��fd��q�eJT��J�址R�0۫q�E��i�ɱ[J��݅� ՚S�.��Ѵ�٣�W�v�9���֧ٽ�H�G��G;T0P�P�Q���{ϓ*i����*fW(^f�q:�F�R[�#OS�7�iq[��*���T�vt���q���C���,᫄�z����8:;�")R��D��"�ώ4���ݢ.���:�ʇK�u��j�+6:�����g^n>��)sA��p�wR��oLЃ�ܩ���`-{,�գ��ٍL���q*�W��Cx�s�]8+N�EF�(��oM�(+��)�U��܅��H���Z��h�:�
U��R�خ�v����E��\qL��T��U�e��A_p��%d��n���]�-����'��Zf+�J�,��i�C@mwv�V��ҎeFF_S
���f��y�+�l��㉁,�j���ݵ(�9Zr�s�ޒ�0��!�w���Pd���]�®号��m���w�C��m��G�����
�)�*S�����n��C��z<C@©n2+�#�r0����zwt���"�-�?GB�Kc
����!��j]��s&u� ��9{�u.k76Sw#?wBC�1���\�OF���8	�gdyʜE���s^N�n捊nvX�wQJ<��1[��C7D�|yvuA��-D��yYӕ�w��X7��;vћ �����I��Tz��4�1e P��w�^��J��լ���bJ5�ԝvu��X�;JK�}`�:e��V6�j�1�Lc��EfGW�8�앭s��c�i��6��;�Ⱦ�
�=�ԝp0��:�v�ڹ2���%Zz�Y�B�p��y�ai�!<�!��	�s�����W�_}�}��@=Y��=�\�H�Joo.îr���z�D#��ԩ�q�W��s�eg.�ȹ����^�ǳ�nR�6���t����J�]��Y�3(7Ց����m�ޥ,,��i��Ms�V�A��c�u{��g���B��U1Q!��Eb(U�9oN�y]Lέ͠o�u�:�C���7T3�$o��1��T�r���֎���|����ڮ�����"H��֖ʁ��*_59�Ew:��1-rg-h��=���/��jJr�ٖ��?ɮĝC3���y����l���Y�y�Xf�����يު������6�3���}%v\]��i�Q����s�}Ԩ�tB�e��q��y��;��6��C3������[�3��]a���s.�6_��A㹴E6C�,U���m�"A�oj�����[��[��tuI:Ï�m�7C/:�E��Wr.��>�5*<��i�[�25��o.�#����ǏF�jr�O����v��a\�������W��������״�IҸ�ٴ���3x�[��j��s7e(���8[�;Q�%���Qr<+Y1]e�V����L�إ,ȩ;'Χor!����],{H�6�i�Oo+���A�]Y,n�;΂3�6����x4�9̒�A�˝t���|�Jy�`᝟rh���gR���b�R�+��$�fl����ռ�8����`,Qm��("(Ѝ�`�*�6�UDX�#Z�ʊUKi2�r�\@�E"��,PR�QYY��J� ��dTTX��ƌXV�4�@X��,@**Teh)��b����QdFLeAVT*k
�
�Y*
,�"��r�ed1��P�V+-�A�X���
b ��E�Z�[d�&Z,��m*L�!YX��[d��*J��\Ƙ��`�Bc!\���+����
VLHb���!id2���d�1�Z��)
�(IQT�ZVc$�RcJ�̤F�LaRLKh�(VE��̧�9����]��������L�tݶ��We�^$<�����a�X�R�m��*W-�FӌHk�*��`O`��/ �Uβk��T�!��rx\5����\{��}k��/�*�hЙ��V��ᛴ�,�<-����&{-��}�K_1���uu����Mj�)xa�b����B�5�z�ݹ�-�nػ�V	͸Il�˽�`=�r���{�љ+,EM�]�H����m����d�F�����Ϻ�7n��k=�W��Bǟ�=k��7�
W�ܑY�~pSԼ�f��C���bq8s�XCE��n�^�\/����<s�<C ޖ5'�P���>�n��5�ߪN�P��0�����c�P���%�������'��Fk#�j�����$���:u��|�O��iz/5�t�iu������Kir��V���w{��\}��B�3��z�eq֌��9vF��n2�I3�i�{꨼<�WR�-�Fx��e�u7����u�dr�W�,��*��)ۦg;��}���0M�;��3���^����{�j	0�V�JZ�t9-0��zT1:�̷w9C�K��������&󬋞�F�m�}���}}��n�������y�)lO�Rɮe;GRź)�@�}4�Os���������鲴��{��c�:�`��#&e�	$�J��;~���ݾ|�s��,��CgLt�Zq'i�Ǆ�Έ�Ǘ��;۬E��x�����<�"���^)Vژ)P�/�ZŅk��_��(��L&���Ň�U�g��J�&�����˚�ۓ1�9Xk����D2-U�ge�c��)��O%ˠ}F֮ov�ne��f�{�&}�:І5sM"K46�g������?��5��
��'��׋�ϵ:kxu��^ͭ(Y������z�!����O%�S:�P"�.�nJC��n#MY�ylg�n�{�{~=�NgGXt�zfq�}��!@���@���p���}�4��tۘ������v����7YU呩��"���ݾ�}`V���52�'�$�=���[]uA��7"�r�Y��ܕ��e���
^I[��,L�lN�g�C��˲��dt$p�4���1�[�x�Y���ޞ��Њ��b�����Rvf��-xwΡ�cѿ����P0�.矃���c�^��i���/#b/^0فY�>*9a��Ƽ���r��w�^[<�&+~�U'�ѥ���o�V�E��0�K�l8��;J��e�ꩭ�F,`4� �����h�C�W���G\'^�����vO7��^��M�-l�A���]Qe>��7�K�&��j���i��{
�õ�X9��r]	�x��q�R��m���Nr:+ZݮNZ�OZـ����!WL~�����8���dև�	"�s���r�����h�^^p�,-ڨ�]�G8�Y��<�%��Ք8��k�0x__���>8�<G=6����63�¤u��5zʗ���sBǯ�1�y�ږ5_�V3��9�
�fu7�l_�|;�W}Y�Ah�/��7��W
�S�ŉ�X\^ǧ�c>�x�V2�y�z�Q`�&�p�����U�p]�=�^3T���"Ѻ�X��p�{),�Ih����9�P��P��5��b�7��Nyj;�M�b�'P�u�[�b�k����uP	y)
��R�-�g^m�[���uu����H�(L]�D��;�߾�5�q]���hqDiϒ�>..��3(�w�kd���)S=��⣎��^���2�����do<o�B�X)M�xK=��k_W�c�}���%9vP����=i�۹���5��*Ƒ`9�������:6�_��/a��E��֯�ƀ�� ��" _
���4��_�4��A[Cƻx׹P��+�#ԐOk3<2W��k�j�0^(�6C�u�u��&���|7g��'z��I�SF���$k�$��K���N:��U�2��o�AK �%]���ӭE���<�9W�שs.N�ٱ��G���W���� 'I��S��OZ��ص�o���1nz\6e����)4���Ԭ�v�b�/������$���Ҽ���K�4[>�6WX���y|1�z�<ͼ��%"���qb��I���`�۞��+M)�`��V�I:�X{�$�/�`�H�6��wT�֒f�<�Fh����W*����Ƒ���z�5�̬�����Kŝ��O��M	Ȗ��&�(}a�X����{��WG��{��Pؓ[Z�����]�ݏn�Ȇ{h[]��<C�_ϮF�{"&'��M�@��ۥd�w�[��=��N�SV��,���|��E�Mz�״�A�lz,.���N,��;��8���L`{�޹e+v�֒��㙺�S:�T�q����"ͼ=��#�Kai���8��#Է��Bp�6����s�x�'�
ࡲ�D�zK�e�'��m�+��ռ���nIͺfc�x���x�;��L���_j���8�N�e,Yc2+����NԽJ|2��OtH�MH�z\"é�'�e{�hϽ�f�^��e(Κ5kvʧ�ܐ
�Q�\��=��bD+e��W��x-B��Ծ�#1�6J�X�44�{-�/�ݫ	�/����"�#
�����)�����u��7��rJ�����-��#=�_Y�,��aF.A�%���xrt��Urac*;@A�j"�ȸ1���Z��,R�]{�N`��
8Yik�P���0��5�L�z��3M��S����d�X���ѪF��ʀ��>	�_�rf����fo�ّ!d炏uۥ�g�� m�c�W�1�E�GFsD`��@-�|����a8�k���ɫҫOy|�Ogjױx�=&�Q3���W,���𹃱g�3;�s���cHG�x�mB��l�.��Ό9�{�6�qy�*e�e�~\'�bp�1d�A�yhi��:��n�9u~�@���華�n�����[L�,w��l���Z�r(E},P��$0���Vue��]{�(����qw�]�Vm{�g��yY��f+/�h�pS�Hg���S�<q8�������+9�P���C|��赺df邓ۑY�c=A�"�ұ.��&N��9mz�����4��(X�Ed:��]���2=t��3�o���0oK���L����z�Bˉ���;t`���Å�-p�u���AS��
�2�����O[#�]�t��V���B륋����|�+�&���Uh�3��۸�Ki�T�u�d�|qչ�R�1���� +PB _����x��\E���
��NKw[=�WGܥ]j�Q��㌷�tE�+�I���7)*���ƕ�g"l5t6rY��"�]�����A�+H��Xײ�Oҵ�K�զ��ۯMv���.V=�{ �����9t���5�xz��zDv�{������ج���(`��;�����Qg�M+�S�;�LļT�����1xG��س�p�,�N$�m���a��KP�&˝գ=L�������l��������Gi��X"�J`��e�+K2����_v{i1�d��?R:�n�$h�{�Y�	�v�x�F���p�K��U����y����Y�����Ṿ�r�h��\��ڹ��6�}8��ɘ���g�:=�Z=+cb����������r��.]zD�NAyf��J&���v�1��8�dX�hm��֫�����A30�/e:�+6�#����5�C؇,��S�"f�Ny�~/���D���%RƮJ�
��w������dE�iv��3�֥z��
s8��GXt�	��=��,6}=�y��R����Vuu����4��S�`�P��;��'QhX�Xoҳ4�jZ��Cz�=���ܱ{-��{gg��ņ�u��z��6OT2Ln�#��e^���u6����V�hi9���hѾ��R!�<���דRR�c=����:М��N<�
��{��{�z;6�Je�=w7^`��V:��܃�r��Y�*���v�&o.��&&'{x��(#h<�٨�-x�����pQk29�VD\��������ܬ��/y���|�Ƭ��P퉍�	�XD!¶�<3�,<*;O��k����>i#����W*�M:/�C�7�ؿ�æ{�Î�L���!W��+��hT�s�����k�S��`{�}���O<��鷫�+��$�4My}�s��='=|1��S<�ַ��E�{��y[���v��{dv�K����{KvG,7�{�j�gm��z��:J����L~���[,h^�7�o_���R��N��v��]Gy��H�\�ӂ��HХN�!��夳�^�V�z�Y�N�^�i���L^���������چ��~�kry�t��wi��}��{+�3i�az�;=�k"9B����R�n�=s<Ƴ���:p�\��k����X��\'o$�������)�,�n̆� `n;kO'G��=�{�4tTJ��.7za�lE���3V�q���o��W|N���KX[�����^<�:�ǫyR<�=`�[Y[8kCa�1��Y�ss��$�g�a�V�ݘJ�ٜ�t��JKS��|s���8�6�r��'�~�~���=����Ǻ�h�z�-vD'���ɰq����]oZ����8�t����}�}#���Ay�Ƿ�,;N��]�q����۝o9����^{�{�sJ�����Q�B=���NՎ�_m۰��x�y��r�������˽�%>��zشK��2on5~�s������Pl�uX���l\�v��"�wYy���Co�\�{d���e=�!����C���^'��"����V��^}����aݍ�M|܏>2����;��\u������+��y">�i�q�E�:��H�\��ԫ�b�p?������1r{���:a�=D��[γ�9�J��k=:y�OPuOў��E{r�l��T�ћ"����x�{~���@�����y�v��Q�gʴsP�v�{z]������w)䏖�iz��K�j9s�I��A����uF�b����2mJ�,pq�t�pu���w���`�f7Ħ�fH/R�B_B���J��S��Ҏ1�幧 �f=$*�SNZ�F��*�`YF�_;I|bk�{����]/�����/Ww��(�ޡ��%~��Kv�w�������[ބ\=�N��z1�&_T�{�[�ĩy�s������޾���r۴9Y+s������-7�Ա��ؚ/����n5)��
Ά���iޓ��ff��V�^]J�#��z�+��_�����S�5��N>�OD��OGA�c���~�g�Ԯ��ض��͇�OgނP�5�Ϭ�/u�<4��у<��WY�Gh���\�n]_Sf�����rm�$�6�\0�/�z��y��ْ���:!����^�mԞu��2��O���佰G:��T�.�\�e�E�O>��B��!�Gdמ��6�`L�]�g�����73|�{x.K�a�#Y�޽�UQ��$���/���x�t����݁�ǆS�%xI�%����Y��^��Y���7pJ�S��4�ӗ<װ�GF��>f���YN�U�`���{�<r��N,z6���x�wb��׏�D��;�S�t�w�����{;��[�s�A�\|e����[l�&��u�SE�z����^���2V˒�z_p��I��i]�f���I�����c�a��3���Lo��c;�*w��V�z_���۹6��y*�x��U�E��v���{%cQP7�l�s�%��;�t@;�|nOPwO���/�)�7�I��$�m�ޫU���[�����`΁?>�ӝ6���X�9�z_�g��~�Ɨ�9<836�rC���ݛ ����'�m���'�N<�_���~������
<(��<&g|sV��
�86�h�/s籜�{�/����6)_U0xx��;~>���MI��{�9�k�K����'h������J�ף�JW��+2�ƴ�?|��b��[�ؚ��t��0�fW�q�B%���{Cm�֯�hr�eְh���C��vr��~��γ�f��� ̓����8�ܷ֬��c>;���r����Y�;=����^H�*o%^�K�Xk�궨�ݩc^t,_ťɫ��9]2\�LY��R�%Kś�B�hc�)yZd�"�ǗC�m����pJN�{��WDs��8Ք�=�kz��E�7b�
�Or��v �5r'C��U�r�]e�Ի�"�q�,�s��
.WVcq�y|H/v�t�;+��8m�7]I�Ȟ;K^��|�%͐�ڍ�˭�u}�+v�)�ʡ]o��g���*���L#W�}fuǱ.v�$��΋��J�cJܴ).�љ�BsLu=�����,2�tO]��E��(����"MI�N�N�NCDtrsAVmǹ˜��4>Ǿ������ȕy���\*�����'wY}7�Hp�R����r��|09��h�O�6�53H�c�O 9�3��s��u��A]h�D��\�c]ƙUc��J�dzfV �b��V�ۥ�HP��w;�ZY *6�<����&�=��4��D�"ҡ4ɽס�3/�� NL��a���P\ѧ׌��N��%�S<:m=T���=���9���r�i\!�+���2�م�T9�+���S��q6��U�u�����r�_~��o�Ec.U�d_I;�[p��c��F[�Av���릚U)'�m��&�a�<V�MBj��뻂�uNד�jǕ��b��/kN���b�:Q����𵖚;��,��+eHjशR�컎�;ߣA���{<��|��¾�dT��E1%�ɛ��oV�7w�I������ �t`!���냆��ݣ#��<`�w��G��&PB�)�|y�k�
��dj��s��򢦮�r�e�e-��iYm�X�����`�(U�,'T�Tt���5ݚ�7-D�b�z�Z���5/g�ݶ�5Dڴ��z���r8Tc��30��y]Nf�뮲P��n�^V�T-�p����+uקWT�ۭ��׹:��@�<R����,GK�e��β����[��D�ڐ���3�C�����:�����)W�ʈ.$]n���ts:����ZZo�ㆥTݻy��ʒ�=�䬚4W��9���e$��:.s�� 7k���l�s��^���
�r��*���R�F]�	�ZƋ�u�!J�YY��f*Vɻ-aT�@��`̶�R{G)&.vk��������0S�;d���3��H�yE�z���`��}FU��u:FI&�m\�9uv��� ���;���t������=SJ�'q��j��-�����c������V�����7".�En&��sG|\��������q��J&Ͳ�wF����nL8����)d�Mn!uA�F�� o(FX�t�����9�Q׳J�V��;�T�.d��T�����b}.��&��Wrer�����⩒q6�%����tּ������������USeC�(���X,����`���J��$�X����RT&%��&1-��l�e@�Y-����,*�m%ADk-�RE%B�*J��6�-T���+���eE��@��!XT�f2�r�2�c+����RVJ2�1Y��0�A@���(VE� �̀,X6��)S1&2���YY*#+��!FH-d��
�
�1�e�E	r�HcP[l�`Эd��2�(bE R��*�V*�F�+��B��"����̢�c
�V-Z��J�%B�c1�U��k@>) H� yo��y�Ab>�&/ξs��b��a`Ӌ�*��t�6����i�dmR��Rc�_p��x�Ep��Nt��j�]o�����7/���7�l�{�M�nq}K;N����y�<k�,��}���}�z7铽�y�l�sz�|.oeH륙�sSˆ�EA����K_(�)�|̾�]��;��nG��2^�N�^5�+����=���K���_(��A�nC���#���ar��3|��6��Z����9��<h':�S�xǣ�뿟31PAw=4�L�W(��J1��o>��]־�k�l ���{<��U�2tW����=�m������c��#F��[����]t��Z���Ny^�y��z�o( ��W�n�s)Ty�'w�����*�c�ޛ�S;y��sY)��'s"뎽/E����3<�V�1�>���*~��Ǖ�T ��M��0;�=����ق��o��k�O�;nJ�P1[������vWZ(e��[\��Z�i��L��;���wKv**�Iά������N�U��˘mNW�jq��+�7��d`CC0i��W;�����ŵ6������2�� ��P�)r�@}R�^�E���w{�Բ3x3E%�ZkV��R�qp�w�>�w�\_���+��ۣ����N)�VV�����"�2T������;q��=�r�������ki<��7n��O��+�>��:�G,���ĩs9N��ɽ��mY��i�az����������<��hAlM3��� �:N�_b+��{{��ۥ~�zľi�d�6��_�}� Jm�u�S�w�~�0���Y'<�K�}��6�	�:�vNfW���U�����%��z��G��9�}:*���;��Yu���1���u\�ޮ�2�WΈ[����η�Ӟ~�݁��v��{�rrք�p{��3l�%;��ݻ����'�x ��'���T�,�mV͛�V�駧��ފ_����\�K�-�:�uX���F�k����{N���ɾx�I����*}��$5�`7�vQ7�g���-o��9�/�|�P)V���7�0��k����}�O�����/�-3�f�O��,\�E���zA����i2K�de������|�vq�avZ����f�y��Q#\ŗ��_0P*��ں$���ҹTR�']��k���i}���ӭr�q޿$��ws$��
���f���w{���)�p? 9�wO�i5�]�~���q�Γ���綑[��=�$��G�\���{�b�p?�\{z���ݥ�+����+0#e�FnqG9i^<�����}=@<��p��G^{c�s<]�%��/�ߝl:|e�G���Υ���r��ǅ-��E���t猝��R��p�F�'��ԯ޴�|9^}[��#�sq��l'�=�����s�y��3�{�y��]�k��-�쏶Y�ˮ�f��/����p�ۖ�o��q��4_�N��l���4i9EɌQ^����4��\/�C�dr�N��Q�}8�|=-+����ꮛ!���F�fq�<����B��`=2{���ɮ�O])+\[�c�=�����{���u�gk�Gh��@��~n]rl��9��c}�0:�*R��yV�a��*a�9��1�94��|���=c��#(�Yn�s��}�f��E���JՏl�[�.t�F�ξ�،��`V`Y�����=\@Ֆ%ɕ����P�B�����k�gR�)m���^�����H��܋}ύ����kzBkާ�%�����,W�\�9н�~�/kݔ�����,~p림�z��zdٽ�<��Oz8�����+4x�wV�
YmZ��R�v�{T��_��k�<�K��s7�d����K�vBڵ^��t����lς��O|3b�=/��x%\x����d�E��`�uMt2�{����Ux�5����6?6��2ę��u�(h��]S�R��	�Ea؏�+ۓa��T����Ϣ,���<.������$��<����}��Iz/� ~�}|�M�s��ƺ[�>UNON�� CG�*��eiC���z+�zz�r��&���:>��=����joܒ�����fd'��N����I����翾�yO<�7���}����c0��m�d��Ry���x��s�a'�:��7�PXO��>ì�J�׽��&�|ʇ�,Y?2x~�~I�@����Y:����4�ә�7��sm?y���/�;	��&ӳ,?0���j{��u	����4��(�?d�C��A}�XI�CS}���$����:�ĨM{��Y>���ԑ�����z�����t�X8�Ʀ���a�U��ʅ��V�����<��j�U֬��F_>2��^x��͞6�ι�I��>�t3qL]�t�Do�S�<�'�(��9����i���w7Ks-e������ӡ�����ƹO$k��N��3��gL#8�����_e���N5&2|�2�|�2i4e�d����^`u'P��c'Y>7�$�d�Vz}�8��js̝M2OY�)�N[���:��g��N�[}�����<�N2k�N�{�q�~tf�J����?5'�:ʄ������q��
�k� �O5���Ad���J��:ʌ��Џ����ӓ�C����U��k�߬��;�ì�$�������l��{�q$���d��̇���VN���!�<d�h�c$����`q����q��XZ��2�Ú����}�oIR~I�T�����<��v��a��`xɶN�M��7;���&�Fk$�>Hy-̬�b�`|�Y8��QG�� �?7Y3����w�������x�~`u����Y;��w$'����d�'9`u�M2t�܄�6ɩ�d+$�<9�IR|��[6�d��~�i���ί|�]�6����6��I�O��[�m4�1����'̇��������C���u��&�{�x��'�����z��ӽ�N&�;�a:��z��y��}��;��~���(N�Y��h,<�$�M��&�u>Ն�q����:�I���O_���d�'�&�;�x�������'�4w�w�y)�������d��e~}��X$���k	PP���J�Ĭ�ei8�l���'��u�>@�9��_�:çy�Y'!�;�M2~a���߭�g�h���w����G�@�}�'�,��	�>d��Y'��*V���iY*N u�~S~XN00?{��ԝd���H.�i��;��c�߻}+����3}�?����������$��<d�O�;�
�2z�σ�C�~d��IĞ�ܒ�I3��+&�P5�N2|��)���8���=��� ~��"���GU;��Nngp��輸�z4�ՊEum���r�b�njʿ�K.�U!-u�ش6����c+�Ξ�Q��5�2����R��ͫD�ɩ��K�:��x:tBu>g���p5�䚹��8u�f�<���������|6f�������&�6����M0����$Ĭ<��a�\�M$�
C��P�'�,�t�R~I��d�$�M��ud�}H�u�'ɘs��<ɟ����}���+	���a�'��O_̞��O��@��d����$Ĭ<��u�c�d�N �5������%a����'��d��'���}��o]�g��}������'�{�'��>Ma�I��4{a�N�����'�8���i��_g7����n�Ad����d�VC����Ì�%`��{�2���z����ٿ8 z�٭s�'�M~�.�m���,'��f�P�	�:��̆�q��t�<d�N���8��:��xI�a�ө�$���޽�������g/�����Z��'䬇y��d��'�~d��~����R~k'��J�z�'���q�~J�k̇Xq��e�$�
��|�Y:��������{����޳߻	ĚB�g�&����&�XN��2u�o�?k܁����䕓�{I���0��!��2u5�q�~J�k̂	}������]���������5o<�(|�h(��I�N%f����I�4��L'XnӬ�}I��g;�a>v���d�:�IY:��7C䬞$�+!�������茶sǷ��_~p��~���~ϼ�d�!�g(~AI<�P���X9�	Xu��Y�{������'Xl/2�R~d���u�MNk$�	�h3Y%a�!��u������?�}��߿t�x��ğ�RC?'r��|�٩��M2Lu�2d�V>��:���6~�H,�C�\�ߩ8��'{@ه��������Gޞ���}���8,�����%d�N�y�V�Z|¤�-!�d�h2��m'^}��i$�F��u������`~d�'_�~��`b�]ϝ�u�ė�����y��|c�O
����nTE&���۫>�A�{t�C���,����T,�u��n�3_Hl֧�S�1Ը}�����/�`̭����qK:��BVwU���H\��K*��Wr�Ѹ/��Ou-����
_פ�Rj��e����)�ӽ�����{)��&�� ���0�����f�5�d+$�<9�IPP�Y�*N ���6���ML,�i8�O���4�q�����$����'�l	{5UO
w����������Y}�n��z��Ou̓��ORx�5܄�4ɩ�dY'��*
>�hVN�d�a�M��	�����Y'������_�n�A�9��5s8�}�f����2|�:�fw2~a6��Y<a��;�u4��M>�НC�N�AI8���IR���ĕ�iY<��u�o�~?>��~��o�~������|��w]�s)>d�N}�l�C\�N2M�C�Ou�p�1�l?0;��$���	�?2y9���O7�%ea==��s�w����w����+&j�锜d�����(|���i����Cg9���a���%eC�s'Xu�s׸x����w �ğ�Y��!ԟ�9�?l�ɟc�x~ߺ���ݽ�ּ��$�'}�	YXM�Ȳq�O���N�������Y8�y���=d����>N�z�߷�I1�}gX�LO��d�
C��W�����gq��������AC��J�yd6��'<�0�@ެ�VIߧ�I��'S^Xq�z�M��'5���OXq'�_d�L�a�7�a>B���<7����'������߼����'�)&'y�:��T'{g�8��+�Hu�̞~�~d�dѿrK�'̜g�P���4�2Ì�ש���=I�^����'Xu&��~������q��~�����>�d������I�6Ü�XOY��q&�Y��'�d��'�̟2x}���d��O�d�'SFP�N���0R���Oȍ�Z׽x������浬��xÌ'}�M2m����hu'P_g�`N$�s�:�d���o�:�������u��䟵�����߹%d���O�d񓉺�������������ꊏP]ֶ�}w�k^�n�	Ɓb�^��R�1;�T��ܟ���x:N��065y����ns�;/���O��G6�Wf΀�gM���N���@����f$�]���������k��w��=��3wV�e/�jr��^	s�ku��W{����=d�2���*xk̇�Y&�(u��,�o��8�ԩ����:�G<é��=�d�&�XOa��ԓ��O|�$�$����f�wg~��~��������Ohq���CYd?'��3YgM�S�}��
I�Zd�T�=��:�ԩ�{��a��u�$�Nfd��O�{�־�y���>~���p�����RO?�sY&�']�%I�C�a�+'Hk,��'�.2O��g�Aa+�ky$�+�XT�d�7?w$N�{���{��2$�K���7o���>��!�~������ON�*I��N�aY'��Y+���䬜Aa�ZC�:���\a6������i�x�7��N2�.���y�ϻ�x�v�{O�y�3�r�s^�2~d����ru�<�s�l�d�ٮ�v��N��'�'|��'�rs̒�a3�m
��
C�8�ԣ$�3zן{�s�{�s����o��}'�'��2d��!�����|����2m�׼ïz��'uI�u�L4��ri�M���CÞd�	�����Y6g=�7�h����=�;��$�ɴ�I��٭�ی���l8��ԛa���Y'�=��O�&��8�'�>@�wܓ��O�i=�rC�4�]��8��u�g��^�o�\7u���y��Ͽ}����J��*M����Rm�~SS�	�O����q&�Oy�H.�:��̝I8��0�$��O8��yܓ��O�Y���|Sv�(5��:���?������ ���'���J�$ɻĕ&�Y<�N�|���S��Hy�잿2u��?s�Axɤ5>�'J�a���ԝI8�}��X�nN�������~pq��?>�m|>d���r���<��q���IR��|�d߶�Rq$���d�!���_�z����:ɤ?]]����?]?d*=��G	�iV~^��5��6 n�P]��q��]�U�k=o'�*:z����E���mlu/��W�L��X'e����:l�|'�,��vT�"W�f_K��w)��@�v��׽�&.�6���#��pR�C5e�_PI�z���s���濭2LJ��5�:����9��8���s�2~J�[�:��'�5����57�I_Y'5�H�w�O��(q�z�OXx��C7߾��+�7��;��ٗS�������#���8�?}:}��	�
�7N��LO����&�X�p?$�O�P�C�?2{�$�&ɿrJ���-�������_9y�M����y�]��ē��t=���O}��x��I����/'��O�u�Aa>C\��q*G���&�|ʇ��=d����g䘁���zky�9�q����y߿^�ǰ�Y1���XO]�i52Ì'��5=�I8������d�O?d�C��A}�XI�CS}���$�����q*A�s�d��K��߭������7��������}G��;�&ړ�N%d>g<O�g'��P�N�?�<d�&��M��N�g��`N$���'SL��:��[���zw_��]~����z���	��Ì�d�ԟ��I�I��k$��`y�O�I�N2�?&2u+8�m�O?P�$�`u��,���%IԝeN���5��>�k���}�������6�L:{��q�m:��ԟ�7����l��{�q$��k$�>d?2�u���C�x���S'�u4y�XJ���6�̿<���~��g�;�w���iX����N2�O{�'Xy7�:�$�Z��?2o�9$��&��$�	�њ�*O���VN1I�l��'���s�]�s����Ϸ�g��Y'�i:wY�L��S�`m��X���:�ߨ}� �3����l�$���I�N�nBq�d�wY
~��"��_|����I��t<n��O�����͡Y4�ö��d�jad�$�}���I㼡�N>�9��8���>�:ɴ���so=d�ٮ�;������W�xT}�[k�����Zc��/KKQs=K�j���x�1�: �����v5KYw�s�����E_g�|�ѽ�/�2���2�*�e3<,f�oJ�4x��.X��oD�=B*#��d�ATmEh�3���U��MB�X��nծ��s��ӢN[GCgM[�p�s�y��}��3� �.U��XO�?�^a*
�6�d�-�8�lх$�N����7l����d��'p�0����s'Y>a5����x�8��1�\��p��5��}?^~�q�L4��$��2o�$�氕	��ĕ��Y<��q&٬,'>O>�!֤�f�~��'Xh���$��;_}���߾���}�~��'�'ݏ�:ɤ� zo�N�L�1g�hN��'|��N!�sY%J�a�q�d�VO2��dߔ���q���r����@�,���׽��w �o}�%�������0��a�����Nz=��N$����c'�,��C�~d�sXx�8�F��*T�'oVM��VN2|��)�y�l��uOD:��s��²�Gﬁ���2i��7��^$�~�:�1+9�:ì&&�w&�q!���8���7Hu'��ON$ެ�VI����㥅/����3?~�ܷ��_��i'���'O]��>d�!��ܞ��=aԛ݁��2uo:�1+}�PY&>���8���;��N2|���I�&���w�?-|����{��wZ�Ͱ�2kVJ�$�Ӕ'��N&�Ì���k�2q���~N�i'nk���d�ӛ�O�u���è,����N%g�~��O�O�M{D�Qs�~�w�z��]V9@��'��~�I�M~�.�u��XO��<g���u=�q����L�IԞ}d�2u��xI�`��?��C�L3�S|U�9~F��H��M�d9�Xm���'gl�>d���Ld�Ԟ��8�e���M2����T�k̇Xq��e�$�
y�7���^���{��ṿ�Ԝ�}� q��nB|�hw;�Y���=�0�'>����2u�o�?� ~a?:�%d���~k'�8��Y�񓩩�q�~J��eM�Z�lJ���)��ə��"���`"���y�M�\�<�7�1u(Ui�O�ȣz�sT��L�s��nd�ptЧ���R��A;�B���p<�s�F3iL'J��=�ͺ94滉��4b����B*,�W��}�\.a�+,*r��� �����z�9���[���e �d%r�(�o;��5�]y�n��mn���6�V.��7�����TS@�����gj�;yvyW�����[ϊt2�0X���{0��G���s:j>�\P���K��v�.<�:A;8tѴe���x���|r�'X�n�:t����ASuxr�k���Y�(��V�+}��pC{���/�:���+�:��-����"��eԼw���
*�N�w�@�ǩ���0[����0.��[Q�Z��il�2�	��c(h`�h˳�0h���8�@5��
qR�wg�T�@3����9�g���gA�~�1��F�5GB���_�_r����B�Gm9okh�B�L���R��I=A�ʻ��*��Η]�JƸ�[d�&ml,/�(+f�Ҍ�3[w��zVGj�S!��Y7y5:�\�\9��k`�mɂ,�o���hܨS����5�P��;�Fέ��=]tt�h,���F���E��+� �ew�f"�bT�}]�wkKf]+�±,��� I7G��f�������u�o��7R�Ι�ŭϜY���e�г-�X���#2Y��z��������J:aU�岦_J�}$�)u3��Ԅ�L���Z�����m���̾���t4����[�"�l#���H�v��M�v1�x��Q�!�oغLjmt�
�o|mb�)�hQ}�غve�[�z�Y�m�F�p`��Un��˅���q��-k:�0hn�<�`�͒�4��V��"� ���.���}m�Rb�S	��vfL}����.纸�J9X�3s�=t�o�����VQ55�;�B���MĠ�1���;�ǻ��v��IL���4��w��6���r��k���c��1+��! �*վ��+g)C���mH��i��֬y]u�q����R��eL��ϵ�ˤ��Ӯ�[H��ݷ��@�gf=n�&4R��v�T�Z/LV���<������
�oP,nawAu\�x�vA`���u(U�}[;�5��+�����UvDP7n�*��ъT�\&�콱��Ǔ�u�"R��߲sW�c����YA���H,��A�C��8u�.�4����C2g�_��6��ɚo�����[wi@yn.+S�k�Q��t"�62�Wd�%F�v>��Z���X�c��&E�5��(������3ػ%WU�p���;S�vۍ�����=����-;rP%t�(B���-%�hN�}3Iv��@VQ��<\(\��Ɯ3J秠�5�ys96p��\�rMك��уr�8M>��;����7��o^{�σlZ2��X��J�Y
���&8�	Y�B�HT
ʬZ�VFؤ�H���Y
���LaU�*T%J�aQ@m�
�T�*Im�clV,"�P��*DeIY*��VE�h!X,���eH,�(��Qd�E
��(�)IF��k�EĊ��J��Z�-�X,�)m �V�V)R�b�ekIQ@�X�%`��#��U�)P�Ң�BV��Z�3)0T
�V�UH((LqY�bQ��H#�Z�� ��J0QdP*5���bԂ�V
aD�1�0��(�R�+*H��`T
�*��D"���{�ue���%��k������J[D,�}�x��ɩ{҃TM��1b�voCPfդ;,tmN퇷��Ǆ���}_U����ږ?��۪RO7T8��
���I�N�f����I�5�0�4�u��:ɷ�s�ΰ���3VM�N��%d�st>J��N3�^{�w��^�<��3�s�xvC�z��;2�$�f����
I��2u+���%a�N�f�{������'Xl��}I���$��M�k$�	�~��}�}����w�����}��Vd:ZJɴ�3YHq6��bI�f�>��i�c�~d8�Ĭ}IXu���l�ܐY:��g~��'���p�d��W9���Nuu�����^}ϟ^�<t���	Y'��2J��AN��8����!�N����m'^}��i$�F��u������̜d����`b�����C}��������?}�Y~�P�d�����!8�2jwY
�>Ne���5��B��
O-�i8�����6�����f�N3�y��N��~�����Wz��Gt��;��~x��~���|�w��4��M��I��'�<}5܄�4ɩ�dY'��*
�m
�Ԭ�̠m�6���q��O�u��ߢ���뭽����t���?~{@}�H�S�~�<~�`���(<�>mj�f
�Q��[� �����{�n���<z:���UǆSܐׅ��Û�59���C�6P��H��&S>��բ��ý�'����Kr>S�Z�ʤ~Nu{Uj�ҽ-,���#v��a����ݳ3z#A��F��o��X7 �S�v�߷�	}`(����p�6	S���%5��+ޑ���Ō�Gv�	ł�5�zt�6���ʔ����q�����~�/0nm���SĲ;;�&+��er �}��eV�5�����)6m��WrK���u'M��������޷4d�6N���w��Ɏ���':˞t�[��S���T����;���G̣��g�r��\��5���l� ���*0���A���wmVr��==��l�w[��A��f�{�|��6����-{�\]|O���Y&�
��]J۶e׽cۃ+���Z�R���3��XvT��0��S(�b����u��;��4��1ٮ��R�r�����:Tz����k�o�'&x��~E���b��.��l�:Cڇ���zo����lu(g:��;�D��^���:<c�]N�[/�[��ͽ2x��(Z���s��g���ə'?Eϧ���T,u*���D�:�� ��Y���E�k���r����~��r}�ޛ$o�,�Do4뚲z�ፌ���T��y^��͹���9��=}c�+&I��:��eӢ��_�4d}�_j�׾F_TZ�۶n�S%j}�[X;˾���2�z;��u�����izŻ�2v0j
��՗Hl�S;y�k�Rݝs�L�BgEQ�Ⱚ'l	��?�^EC{��v^�dv	���=�Q69)|��Zu�.Z;��^u��UW�W����G�8������y7�{���_�����d��%�֯���}x�<���!{L4����ع�GK���q�d~���
�zI(ʇt9e�vmu>�&]�n�.����iʛ�K��ょVo��\��{��;Z,8���_=�ߡ��T�8���ȋ=]���W&/{q��3��F��V���Γ�6�h��O<�K8��]B��qÙJ���<���O}��8[�zpt�W���%��K�|��g�����C�%�Q�e���[��K��3�'�N�K���}*MT�12����]��/�n��Ŋ͌m[�+��f�~�bZ�ї+�-w�yr�F��l�_:��gw��v�u&pLvk�{�Q�E�Q݆m5�������@&����Y�⟂�K	��/��z��P=r�,����%����UG�:��w�mvk��V.gn]ʷ����v�3JEA��F\�+우�ZO�A/>w�h�m/O�m��4���#�V��y�L��l����`���
�2�\�uX�з�S@�$�t�.JP��ϸ�kk�˙�|L�׶�� &��/���9��o;�:cR{}9�`�zh��/S���R��x�����I�߽[@�-�6�!�&��tƷ��6S�Vv���Q嬚�˂N���f��lJm���(·��}�����u�Ǚ8��w�mCx6��[�6����C��ް�:�s�����y�xl�';�����h�SLX�]8���r�ӽ]���tBab�>��J���?9�ҷ݁9�4�<v_�z�:����VG�����/?O�%���;����a<�� �r�z6o�"י0����y����U��{�Kђl��;%6x�:���]�G;S�֣�9O=��	���g}&G��{�Hk���w��&3֯���v2%���{�$�
����������Z�a��/���5qS�~"��E?Q����aB߾���e��U$�۾���4�\�瞛>�ĺT4o
�C=�_xK��]7������9��q�~sث����� �+K��v��bʺ|��1�4�i<,�<Y��P�.���i�1���u�;f�*i�`̽A7�*��_v��mf�^���ѷxᇭ+IIg�ئ�q�N�e�rr�:�}��}�S�T;W{����۸�;{���)���Y���r��ޖ@�1��ƧY�y��|����v�j��,\��\v��ٹV�w���9CR������y�w���~��{乿$���^u�b���{���WL~MYM�էy>�+�]ެ���N^g����k������P�v�Sw|��6=���-�r?W]3.�(_��x�}�R�S����W�у:�+�C�*ήF]e瘢�>N��Kz��b�8u��o �'N�{�Mv����'>$�_|R���mA��1��P���L���%�]x@�
�k�U���uI����s��_�δtqcN�%�oR�T~����%pg��C<���=�����j<���#��u�/x���9�۝o�^�0<��Fg�����e5���^ɟJ�|���rL���]�a���[��N���]�V�їm�n(���*�K����n1���N�|��+q)l�M�d�����I�ff�GSt�.�5���BO,U�	��y�{�䃍�g:X0��YO�y�k�V�!�|�-w�s��øu��ת��ɹ�u�׳�kx�y�~ ��hkr7%W������o�gΟ�_�>��|$��yw��L)�MeD��2�w����9�͋�|�u�}"��Os�x[~�w��f@nv��7OS�B��'<z�)��
�޽���{��nG�Ly/q�6j�8,��ù�+�����u��K�)s��ܪIs�w='پ!����2�Kܸ�n�᷍�h]��H���u/��h�~�+N�V��������m]�m�gzNzlN�P~�۞zpt�W��oC-�=<�%������	���o&է2;���p-�����3y=۾�h�;R�zr�39;�!�)����-�����le{�\��^`���7k.���������<���,����M1_^�Ŏ�8pm�aԷ���A�={����~C��5_�S|�_n��mx{E��;���28&��C[9�2��م|��"�(��Zs{����v�5O�.�N=ܱ�g��}�+6�T���w�0��f(�sw| �[�˼�v5)�O��(���k��E䓉&���$F�s[׺�G2��&@W}����i\6�/���r�������O_)�৒V�_�N�xN>�v��Vv��n���k=A�pe�V�;f��(�貤�>����.Ms�.}�N=���|2��[�m9ճ��-r�~�'��e��޶����];�} }	gi�o.y��{Ԕ�;�>�ϐ���[jL�=o篯�q�K��u�/�Ԩp����%l�΃�"��_'�GOnqv��L������j������VQo�.�~<����t!��=�9r�OL�Vl\ގ�8�	W�u]V�J��Wfk�?n� ݗ�$�Ġ��	��#�ܾ�]���c����;sy����O�p?��:O�����l}ud-���6�{�����Nٙ���J��n�}=N���~�D�<Ĺ���7y��ޟeʼ��ݴ���o�T�8_�y���h_��R�S�0�K�$�8|�yWV2��T~1���tX���j���r�]Hi�M���CI���ck�ya�vwv3fv��l�b����H���ԱO{";ٳ;���kq��ɜ��5.��^��^�˦j�39{�[��_����=�3���|f��mvIo�o-�L����c���o��>̦>X�����s�˴���W�qb^ӛ�F=�5�{�i�����1T���u�%vo'癞1�{��C���L��j�L����
��Eˡ޵�3^w�����^�qd���9�vռ4g�`/T���a������J�-���I����ky�bO��réљ3�{گ�³��>1�'Y�H�޲�U����=���B�Ca��A+������b[�Vvz�6�[Og{ٵ6�L�\���4 1����l�ɳ���lS�:σq�}8��T��g�~����ɣ|��!�w��nu������Ny9�<��iݾ,K�-�/9��u9�ؖe}(��`�ϭ��o�k��ܛ>�ԋ� v���ܽޝ�S|�o�y/o.u�çd-fψ~��_�\�����U;�J���ws�w���ec�͜��;'�+E�;)E�1U��*n/u	�1fs����L���b�e�9�[���3{5(}&���w��ʹ�|ktxt��'ɾ��ݯ�:��3woo_9���%�o�;��M������Ɏ��4o��_}�W��g��ې����{d����z��jXu�Sg�':��yk�aek|�9�u��w��d����5�m��Ӿ�}g\����=�k>���W�WZ���n?�.���h7"���/��~��Ӯ:1v�����c�"��^�L>wy%��?}ݷ3�A�
����󝗺��*���mg��e';Ks��ⶎ�U�{Ω�z�o��}�9�@�<��/��<����Ӄ������.;[밞��*݌�=4��~Y5���G���C�ש�������#伔��󫰹���X�}J�YvE��.7���O{մ�AZ-��\��8�>��mY+��(��򝌫�����%��'�{ƅ֊�1}��G/�R�}�w�9��Jo�qJ8i�
gZڞB^o�����-'_V�B�8o��!�&����>�x	<��֑�90XΝ��҇t�O@+�]�~9�4]<�	���)�ʝu!@�����雍=:W�j�Y�f+Is�����S�h,N�{�-��k���TCX��U�,�q���1^]FᩓrtKz����%[�.������W�}UU�7z��Ձ-Y����us'9��.���d���6�vS��8|���%#��S�5��Ǻ坧Gh�l�K�ޥ����5ޮ�M�lS��lK佛qW�7�`�ݗ�H�Q�|腼X�y�C��9\���d?��~��o�-���~���s9����eT�ߝ�_;!oL^�P�!h�v�\E��վR�~�F�mK�+��IU,;j��m��Z���{oc�%3�;�M�͋�|�u����UǟOd+�y��A�k����s����̪>����{-M�b���d|:��&����;�8��I��g������W����.���[ ��W���?�ܤ�;v���r�����:��}�����P��uW5�a�G�]-���'[��U�yə����u�Sz�g��
��f���3�b�l� ��}����d�i�ͧ��(�v���سzϯ�����Re�#�m�^1�),�X�u�սܩ5�yCƲ��ںsb;�܈:EۢB�\������ǃ����Y�P�Cx�>㨧��cu@�h�y8X���|��4��ԧN�P+��2��Y����D �9��ۜE��["ǯ9]u0����3#��y׷|frEߐ鏶�oE���x7-RMZ-g"A�})6�2;kG:�H��|�T�Vk�L:�'q��:ͻE��Ǜ���/4$��壖�������`c����E>j���g�*�*D�umʰ�F���CB��t//\δ���=�� 1�%��R�v���Gt*�]�n}���D�%y���Z�K	W��p�"�(�4-��(�ˇpN	Nf�&;���QOa���7W�ǅ&A�p�8���X��.��#޹63��Ѷ�*n�V.��	�v�����DZ�%�wd8��z3yy;���i��tfz�����S;���SC��ʄ����6:��B�a�^VRDS�x`��9.�i�V�|�-n�N=�{(̫1v��	uT��9i��W�A@���o��.���at�E
���ڂ�9ٔ��5MZ]�`a�ҹR�:#P�i�N�;��l�2�X1d��֝w�ݼ�Ȭ@tR&���@ھ��n��*�n�F��xݚ���d���W���{�#K���Y��?�-۽x�Dd)�}[�Ǹ,*����[7��^��sIW�S�X]��B����3z�#{����|Մ9噡������3�Y����{{1Y�bK�u^�ӓ6��*����:s��yohxw'>��2����Wp'-V�YW:��P��<���[�յċO��m����{i���ޔ��ni��`�x���H�S:=�� 1i��+�-A�wW����8��1:�څJ��ʔ#�3�_!J���-꼔V�μ�n�5��F5Ϻ�Q�rѢ�UkvQy,���znk:�p��O�rs+#f��^��4�̝�׮�K�95|��1�3q�����ޮ���M���U�o�atPpC���;/I��JB�,�@��xܧ\f�9D�}{Lw:v���R�Z�;�i��e%L���9�-��N����R�Rn�ZMu�3h�l�hwc`j���"��	ڻ�����E�nl��T���μs2��#�2�[ꐇ3mռV5���c�荤-l� 嫑����82>�q�o^����!b�օ"ݯ�����$�d�.�v���o��fu�
x�wY��ww�9}�U�1|�>Zc����v���]h�U�]�G6�dD@��ۢՑ�e�w-Ԯ���U�����v���*s�xܮx.�!˳G���̾b���,Y
�Dɮ��F�t6��Z����g~�(��
��J���6�A�8���y�C��r�����+S��s�Y��]maU�#G��;��m�7~�����!��PTH*��E"� �`V��P��Z!Qk��Z�YX`�DR��H�bdE����+���"�*�V�A`ҕ�U(�"��Z�YFT��Z��)�X��ʋU����[D�[j�ʩ*,P�%IQEZR�AC)Z�G)b0�(�T���[+"�ʨ�ed�T�jJ��U�*��"KZBڰF �T�m�X�l%E��P-�J5���FH��j�
�Y*AJ��V0�2Vƪ`�k
�2#-�#��
���,jV�0���eb�b�`"��(��)[A������J��*[V���(���***��U��j�@�̢¢�3(�	G�)S{�h�켖��u�f5��9ru{���pG
��<u:eЈD-^e����u ����z+�$������v��ח�>���M�W���N�s�d/J{�-}��Xϧ�E��Y�:�����Գ�T�H|�:+�ڣ<���Y��qԼ�q��n纄��;��fݭz:��u�����8ӵ�e��]1W�1���r�K|=q{l<�/��#�|���ܓ^�g3F`�4ϔ3�z��῟��\���O�j����ϻ��sہd�Q��8�o�ol+:<c�]N�[.�S*dŒY�\�j���o<����z	�&�=�w�K;N��>/�a�X�.%�����WaˀK۫�{�o��O��C�� {������E\���-x���q���!����xI�ۘ���<��&^}s�8���Y���g׾�uQ�腜a���:y�}�r�>����;���^X��&�Tv�>�׼���j��yss��wڝ.�6.x�t�n�����or���e��{}�
Z�\(n]Gv�Q:n0��w���Jz�Q�Rm�}�KSqn�-<jș�
�n��y���Kr�FLYՈ�;I�l�]�U݆�P!+ܢbqY���R�G� á���Yt��C�6�\�8:�复�e�{بMp'�M~�����K]99sk���~kwIz2M�bS�WpЪ�g��Ʈ;�?']���]�x�]%M���<z|�F"a��~�ӱ�^���>��֍YRf���W�y�7���7�/d���b���OPwN�<���Q-�K�M�������ͼ���s@��7���T�89��zm��U��z��_�gO1e=�0�3~e�p�y���^���~�������ce�ܪ{Z�gpK��'}=��o�����l`�t�6�oo�1�Q�W3Y<V6�z�>n3d�v��X��gex'�_]I�˔}Y>�KY��el�ӓ��褼�q�Ms�׏��@w�;�z���߻=���&�;��hKbh��!��[��R{g?k�zh��9W���G�K^�u.tts<K�+��p�zd6>�%t�05���͹o��
C��+�[��Q���jTwuo]&P���a�xX�������ɼ���<t�e@A���[���ŗI����Ap��ln�l.Bw,M��ۥ�������c�u����f�__rދ�g�9ח�)��+I{C*	�7��H�/�[�_���>��:��o��Y��0�_u���e��l�����}O|��o}�x�nA7TE�8��A�z���\#���\��q̛#�ߎ�٥3��w���9�{�Vn�I�3҈�0a���_�-��6W��;�\&iV&]�p:��Vx��y��/kλ��t���|'K�|M�J�ծQ@u�=E��^����7*���r���`�k�a�vJ���U��R�)���'��r�3���u���$���{!X47���:u2�g.[�)��N^���K;�<����nE��b��K�֜�-x�^�W��ɴ�����Vx�>�Q�ީ�	��b�V�E=+5�;�UM&<�E��%����nzm�*e{Gs�į�s���X��=����N���3�0�͹�;=@z��������O���J��Q~���7G-�KTDz�z>�ˮ��3��nu��ӫb�M�h6R�e�*]kG�R��S�؝)���6��kV���V�6,�k�c��V��i����َ�w���2���:S=��}f�w�r�:]YD��5��N���I2��꯾���ڽ=���O���1��y.9{��f�����^O��4�ds���{� 2��y˖���]��u/U�����*���\���`<1��T���#�Y��;yg.��������u�h��8ԩ��{���ܭp��o�B�l���_���ii�9���lc��!h���8�q]���L�y�~�'�M곣�O˙9�g�Q������I�z�gD���~����m�O��>�{�K;N��<X���·�Z��U�5	Kn{}�f=޹�{�tT.oJ�3�/$w(��X��m�I�K��_���ݒ��2�͹���E���{|�ʩ%�\�a�����Σ���l�Z�c����M�	(^�ۓ��|����~Ϝ���\���왻�V\�94FM�P��4��Ohf�����Ϧ	W�����z�W�1J����YR��#��]#����_���==t+S+�i�:��՜=ک�U�]Zu��ǳ+u���,�Gp\��\;8�C��+�x���W����2����g��XƳ���t����M}�y��<���_��꯾ m��q��2˱��T��D�g��M��~����vu�C�I�=K�k�ɢ��������v�'�v�D�;ͧ�'V��5��ݻK��@�>�0���0M�W8Ň񾞧u:Ϳ}��t�����~=@���x��������Ӷi��*~���y���k��c��g��+L�+��C�%�g�E=�-}����ޣK�(����j�����-6X�7�<��ƶ}��}��Sƾ�����c+� ��,:���8�i���}=��짗�u��w���@gv�,�]1B�F/���p��Ʒ���y^�}5e�/r&�+:Z�+��NתZ�h^�]��{��R���u�"=������0zs���G��ӏ��ޚ;��&N�6x��}�Dw���2����K�&w��&�����^Ѹ��.C]Vv8�m��W�-*1
qi:���'4н�ӕk�dن�t�LE�ӣ��,PÉ¬���v}���g>���UŠ1H�\ܣT�X|�^���k���,�vQz9=И��YQ�dA "�>�����Ϣ,�qq�+]ǔo��j�ݔ0m�����oﾪ����2�܅�z��.�}uasf�{�o��?k����7=����j�3k�8�{Wu�u��}$�ν�۩=�E������V�e\��=����r삜�w�OF-}�Q��f���+s���5�J�fVOA=g�4Rk����ú[m�y��/o�w������N���l\�����G)�Evv��߼�ޒ��Os�%�Ϥږ%d�x�OeX����ֺ�k|91��N���eɑ�2�p<���;�%Ѓ�)!iCh�;����BO���+����wk�ވ�{%[�Ň�{�\�+�����ìe^�7��P�ჳo�y�.^\����g��M��W�Ӆ�����^>7^z�B�s�@�=��f˄�T<V���������E��OR9��,oKY����ߣQ�ⲩj�H�aw��MV��+� ܝ��t�y|��}�bq���s�5.��X�d� �<�S��C�����ե�>��=5xA�WF��=sZ�V6$
�f���Ż�L�v�mL�#�L���-��Og����k�z9Y���ڹ0��(g#����S�}{Z�od7��\4w�M@������|>�eI���6�ۯ~zٱ�M��Չ�q�ke����ԏ9�Q�ٱ��y�o	=+\������;酏-��Y���/�{��y	��fo�\�u֘.h�lt�C�k�N���9�X�{aYܙ:�	ޞ�9J��<x��G���m��b��|����ld�I�[۟=3ipb�/X۲r���F� Vr�f
;��ֶR�Sf��M���=󮮵��Ч/:�����s���,�Gk�x�_r��{ԹG���3��o�옑���>�ۤ�����۾�""������Cs����Yj�l:�>}�y%o�|%M�#Ω+�Si�����h.}@�yv���t1Vg����jL�'����%_�9^�%�Ϥ�Xu�vL!��
J��3�7�T��=uT_{<c��u�ϙ�&G��{�x+��b�T�^���=4)��(�o�����ܼ��ѝW���j	9����_:k1;�%&Jx���{t�eoFħ���B���\�y�ƛ�J��(Kg���aSyh�>ɴ���6��L�ӝk�������{��}hs�K��4�j��;���c�w�K�:�3�����m~�����K��n*������}��)��V��f�����9Lw������(�x��G���׶�W�g�ܓo|������ڣ�a%R=��w��y�6����NyϷB��c���'a�2��8�;�D��W?u��͑�3�= �q^�{�w��q�����K/�?s9m����=b{���JIݾm�����w��r�>{��M�������h��}3�y�cw��0wV�a��fpLo{��k����9ǳ\�NA�_�H�_%�on�7b-9�=�U�&�xԈ��a'��31ܼ�Kz���¼SdMR��{E�4q�R�L��O�AǤ��I��Sl�g�ȖK$qQCS!#u�)���o���w��ƣY�ʆee�B֚�#�6����z"<8�z�K�z��QƹŔ�"�o`0�d��Q�'[��f�/�E�T-I��x5GP(���Z�l�W�t�b+��Q]�����ە�Kֳ:�m�H������x],�}jQ����^�����X-z����5<��Z/i�]ֹ��t	�5�Q��,ɺމRsy��|;]$��v��}c't�Hc����t�n]��'O-��W���]d���qd�U��o�aW�<���씅���Q�&Ww�<$�r]#�:��1�N�5,��aǅ�y���t��=c��	��M^�Z}����㼵�*�R�Zv4ϗe+�#�	���[�1�r}�I�uP����U�+��1�|*e�~C~X�LB��Ga�V��/hȨ�l���)��ƹ
�<�\Ur���;yIm�kb�u�^����ݙ�&�~��A�/a�E;]$�Fk��\e����A^�ݗ��1~Xk菰d��̞���PuC����\��BS�!��!W<��-�x���F�����ȫ�2��^�̥ �{�]�`��}F��\LpSԹC�
�lr8����(��4]�Bh��6HZ�;�=������5|����ƥ���V̉d^,�ο�x2��g�%u9���ۣ�B��J��r�����5�>�t�Y ���ٍ/E�Ug�躬g���S�����5�='5�V&����K����g�M4k+L���fg����n���;�ʄJ���(R�լ���c@y=���2��#֛�9��+e���.���R�Ԅ��m�����] ����]�w�4bO�[Y�M��z�屑"�ؗ5 8Cۅ�K�݋e���"̓�2��]a�Tw	��-�ݷ{����{y,��a�Y��ͼ�[�O�娬&�ł��v�T��e/�W��K��ėu���[�5ou99d{�|���^Q
�{VK�è�m����C�P�V����W]�ҧ��ƪ{�G-�ӸғMCW�2�m�O��/:�7U�
�O�>dhg�T�EFN�\�WpTٺK���+���%M��$�(��l�a��MN(�4Ӎ�1.��v����c�5�O�{��X�*�I��TEp��X�Ʀ��M{��x3�d��#��]��Kڕ�`�y�x6���A}z��0����fX�y�J�1�W�|�g���{�iԁ��,wS���/x��)G�Ԕo|�X�8=����a�	�ּ%��uu�k��P~�ʻީ׻Ӷ�f9Xt���38�ʖ��!�΁
ƧB��6�ꦶ��]#���h��|ϴ�rr�p��<���{�Y��|e\\|Pޣ���tL>�$��ⲓ�.�����$�n^����]۽j	(ř�t���Y~]�\
��i��m}^�U���bIm{�]������)a�ș����7ܤ��s:�D����v뭏�Ꮊ��yC��q�/ Num����b]�s���}���nv��F��r�W7�(6��]k��up+�$��;Fe\�{չ�VJLe*�6��^Wa�!\��j�()L]sHf����4�%ڜtK�22�ci�8�U�ˁR*�Dq�멸�$1�Qٸ���%�:-���zmoaֵ�/��&r#9��E{�.Q贷P�\�!r���k�Ġ|t�
�L��}�|����rIn�ȹ����o#]C"R�R�\�ޥ��o\q�H}�{Җ�_��h��.�uo`�#�L;�W�w�<�-�z)A>���>�V�W2�E>\5���N�gF�>v!�a�Ǽ�5Eނc�\�QNxv��IѷEgCMN�T+D�92�.be��vVqsx�K`�5\:vv8���V�{�E�,Tڽ������r��ˡ�-�S��k�ƧU�緼�����	�����D��(o�_2M��bo��%J������-K�ݑY�\�fl]���"j���;���z̀��c�I��J�*�ʕ��ӼW������7��r��c.n<���إ�u��7��u�'�l!ݹ���n��9�e�B�50����}N+m�lL��)�S�g<0ܰ�V�VyLn���������2��C4Χ{��������G�@��缽��oT�����+��J���[���M>�jR�ס�M�f<k{�p�6r7��,����Pw^�*wh�F�ɰ��'�u'iI;��^�R�ݢ�}��]=���h��5gC������ܝ��Zy�&��$�h6�nA&�G:�6�Smtwp�Fqn�D� ��O�w��}�=tL@ˡ(���sd�+���<�7h&���H;��t�|Y}	q�ۺxWs@巚뤬E�g��9�N��]��.
m`y-Ip*ζ�n.M Y캓^��]�k�Sn����^d�Y�Z����NB��;�l-2��귻����S��Z���d�)WQѱ�����<��_e�U�d���E�ފ����K	�;J9�Z;4s�:�3-Z;%�fo�g^��"�/��́E�`x�b��V�Lcf�\��d1i������j����o��@|M��%�a�mu���=�S�j[MF>�m�C,��o�u���ڹ]X�'�����yƘX{*�ZB`����R���1�5�%ۤ0%\��SԘ3m�B���Bo9N�:�i�L��7B�,�
�qP�!jKe��]��Nv ��B���Q=K�vu)+����Zj#x��Dj���`������|1]� �=</O;h?PI��wE��b�]\du��Gͤ�pFѭ��{*r������Om%I_+�����Y�ǀ��I�p��6S�j۠zpTFٸͬ���:�����m^���H(-jVT(V���b��[%Ls(*�h�Y*���EDS-��T\B�4���Q*)Z�eAYRڕ��H@QH����kV�,ET�ֶ�b�b�bb�QJ�HҊ��mh��VB��Jȣi���
�[B�"�Tc
�Ƹ��dZ�+TDQ���c!TU*#�*�(�el*@Z�,2�(V�YX��h�E0�
*-�aP�P�Lʡ�2b�˔�����[j2�,*3AAC2�d�c���XQKj+�LJ�`��
"�.P�����U����*��E(V�Z�m���E�J�-�IZƶ��X�

Ea�`���`%��X�Z�B���0P��k#hUHTRQPA�	 �B ߼��]�k|�k��7��j�\�[ǚ6*�jﴦ��ti�<�;��#�aK_ts�]��P�U˼���2�y��磌�H���(��)3ԻS:}�X_���
J�T"��� ��g��ҥztt�R�7?zuo�[�=v�������8An�|lg�3���Z�7��M�B�M���8�^���Y������ח�Ġi��څ�X�0�{P1�΁��ș��o꩔�҄�T�$k'p~6�MYv���D�'�������� �ԤYI�̩cN%M>���aq0�	f�T�߲�c�	�~/ ��/c�r:��3�v��/Bc�R[�'�ΰ·=N$�Q�odޙ���șރ�!�E����N�/P�Y5�#j�;Xj�P�
V��]vEb%y�{������g1B�B��(��/�����Թ��.hoUF�� �Fe�f��s�~�X�<|���`zbKG�S�@��v"d+>���:���o.Iת����3ج�q��h�iS0���l*2Zv)W��0Ӫ�#�N�W�(���%K���[�������~�f�tXrq��YC��Di'�`�	kS
��ڣ�ܹ�]�SZ�i.�D�5��3�cW�&YT�-j����V�$0z��w�p��K�N�]N
�����C�ݮ�T���y���
�(���Dޠ�B��5Z�>��h{��^��g�Ap�>�}�w7�Ma��ك�RLͭ؆���u2�R�K�t�:�k�?|>4{�0_�佄n�|}�����d�7��-#=��@�����w��U<��������b��]����
��^��6_`��*ƑnG�qђ^r����Ir��R��H�ǡS���2��c|�C=�
��1�1x�Q��5�e�▼8J���0T6f�`�Y���o�m.R��:����x�/�s��`���	=0?v4䔭xx�w{��G�˨��ǜ��T��T��e�N�#��墓�X�hc��c�	Y�h�.(h=C�Yz�Q~�3�v�~{~�$xO+yv޵��}�O.ϯ�I��ׯ	u������y���$���n�l�j��.e2N�P폽�b`�Z�W�L�c۞��N)10�b�#���]�>l>R���}(x��>���"b�%�`z�a���*�VF�v��n�WH)=^�&�/R�,N���x��ܱ�)kN=��ɻp����n�^���� ֫_�;~v�T�,�ii�S�p��p��2 +�%gx�W���θ°`X]�����C��=c���ʍ�����5�N.��dV{r��O-U�o�}a�i�P{�^G�.�q:X�uǠ�W2�,��p
�!�^���!�� ��l<O��=���aj������\ؽ���]_磌��S��z�6��+�Ce�������Z����H�NE�@�^�;���x4_�H�[��x���])F|]
�K��g��L�5�8�a��꟪��I{��r{fot�;$V7c���Z_99���顀ׅЭG�ȪΟ<����vw_��]����<�����<+��0����G��o��Fi��e#�.��a3Px��B�l�]rCҷ�|�	j��+���p+ə�};%!d炎L��VIL��e���'Y� �f>|/3��o�u�F��h!���A��۞�~K鰻:��Kf病D��Y�HRg�O��&��|���*��x��PP���a�7u\g)�L�/�C~/��n�ᙐ�a����QN4ǫb�z���tƹ��eW-�mA���R[e����f*��2���woZɼ�˟�����ҁ��m�Eb���I
��yg�댺��~{^�!��uS]�5ة���	o�{��h��/%[Dۂ���C����A�S���{�ow���<T�u��4w�NW����7�b�u-�N��^MӌGS�uG&\��%�E衽姼���Pa�4m��y����u�؇Lk{D�W��V�F������K��[nyT}W,<�T���+��Y1Rݍ�q���X{Gh�Ǖ�  	�S��p�Vա��3ܵ��3zX��=����=K�>4Q��#�:�fz�r�}=ޕ���Gո�0�KuE>+�љ���L���~��g)���9	Y�b�Γ4VHVof�P����%�Eh�2����2}N�_W���Ac��cH,3�r�2�w�͕��W�Aߪ�{�80�������`��8X���v�{�X��͹u�2���j�̙JG�쌍�e	�^��t��M+�-"�#ʕ0w��P�c\5]��j�w)��i6�^Ġܾ/ �3e�;�%�_��WH��U���ʬ-�+35��1����y�V�u�^J	���+ř;��|K��8׎��g���G�C���߸�K5r~�ގ�'e�!��E���Z��S}�	��)���W42q�۟L�t��naQ����2C�9�)r6
e�����;.ȫ����S;��JSO6�K��yw[���9���_};�,qe�aݠk플W��g<�<��d�^�x��>����|j�0kM�3Z�ϴ�Yb�k�#��k����!~��C�بH�*&fu1`3-�C�/�;�GՒk�y��ۭ�|:��jÏ_=��p�V�'o#X�^����|��y c_0�15�5��nmC3z��V^_3�oJў�y�En������Ӳv�ކ��S��7�CZˮ W*���&%u��A34w��&�#�/Uҙ�`�=��ݸrOmwx�w~0�������*ZmCY�I��~l��np��.VK�e�����D�B��%fB�e\\}7���T;L�a�l�]KF{�?a�о��*�����ˮ]�_�n5�Q�3�`F��� ��`�
�FJ�lL�0�|��`5�<�ޫ,Q��,0��pt$��/\�XA�US�U���3[��R*~^R�/���-���]�cj�ͧ􏄹�����ԩ�S���/'��سއ�:�Aa�����	]h��YUxi�*�>LpU%����ȃ=%L�^}���4IӮ�a�3����i(���3�{��y8���u��|k���>�v�/}/8w��ib|7-��4|u�x����.����u}eK;5�<Lz����j��/Ju�v�*ǈ�����D��3�k�P�S]B<���V�`ֲx�P�L���y�C�B��/-���Fdd�n��א����F��s]�P9㒆\���``13#k;�y���������y ��ݰ��ъ�{ا%�y[��i|�M7��e�C:n�k'U�4�o�9D�H�sa�|x��� >NZ�F�7GUK]�L���,_���QE��q[���K���C�hY��طtqŸ�X﷨�PV{�Á�y�`~2�Z=>{�s�������b���B\�j�0ߑ�����X���*_o5����|��C�U��^I�-�^}J����f�w"G'm��w���ж��\�=��~�������M�B2��j��R#p��A¯������3�e��t�m+N��
�D;8�� ���{�&3�zu�+>��<o�j�R2��P<D�滺���ܸ�^]{��װ1�VJ�SS��=�U�"܏��%�+�Kg%�0�h���}�ҟ&�h����I�q�!���lC�uN��*�P~P�X�LZ<�x�@���[^����V= D/��ZL��d2��7�;-f}�Q\���2�i�z���71A���y�K�M`�W����:�%{Ȏ���Mc����r�6������f^Ч�d�V��L��4#�10]���^L����~uy*�x*�K��Q�%H�^x�n���{{;W_}}�*n:4jv�[�]{���Y��n;3kz��.���je�J�q=c��T|��C^V]�N�`]�Zڕ/H�|z�z�j��2��nN<�+zi���@��4 ��w�Ε�h�\�ى�۲���7����z���� �ه����O]�_�t#D��z�&_�4skƢЅq�����m�ϱU�{�l��Ӛ��V��Ou�������C�[�Ѱ�<DLO�o�^"�����]����c�zu��8�A�R�W��z�"<�0C�{Oܱ�襭/e4��u��n�/KZ�+�޲�f��ÎK�d�k���bP�WR�~b��=�Dh8��s0{�'��\#K.�;�c�=�չ�ir�Xb�z�-z|���x�[����{h�M��L�lS�g����o/l�9�/C�5-��Bj��~Q�B�R��F��H��WP{G�H���X�γӽUϑ�Ġ�d�'X��u�Z|��jZ�ue�B֚�u'`P�}�R�>o��Ŝ�.NƲMїA�%��o�a2�X֨����x�6��#_�#C<�T��xg��l�,��Nq#�X���]Nߗ|W�3ӮRd炎	����Il�G�ocTײ]��y��k�þ(��K��T<H#��ԃa�ɪ%㜻�Oh_�s�=k�*��O9R�����F��G"�\�m����!�Ӗ�Je�WQ�$� ��nr7Cz���ڊ����Tܽ�O�]��x<�����nt1V�{��4Z���-��W^>w�J�ԭA��sJ�k�W;�N��F��)���I��������9}6P=;��C����+M��4:R�$�kh(E�V �o�ϝ�1�T����o�R�m�m�{س�m��|��18ʘ�z&;�'�r&9:ʮ[^ڃG<���k0{���78a���y%���7����{�P4�,�|�Pw�i!C���3��G����G���F3�w��ӳ���u>ݖ���\T�.�D�r�Q�a4�<��}m�q��E�I�o�_�o�&W�vK�綰Ng�xC����OR��+4a������}��x1��o��A��,4sץ?���@ϟK�>��_�fD��ϐ���?6�������a�V< ���b��W���o=����v�2��E�ǖ���l�x�=��ǩ@����k��ٷQea�k��v��r�\~�%���ޏx�W�J�p�X�2_���gԷv��m�2l�ܴb��-E�Ҩ���2<�SxOjT=R���{��w������E"Y��K�;�w�Ϝ��n���2<pO�#�Ҳ�W"��ս�e3P�H�^��#-�V(�ÕC����8�����䊖��2�tކї�[��rd[�v!n�z�g�@`tE��C��,x4�����\�����fY�SFg,��"�y-�����'ݎ+F�
�<Ý�1V��:��嶇:���*^�f'��U_y�Y��ɸ)��A��=5Y�x�-��P�:�=�Ӎx�g��Yh�Y�l�&G�Q�>�UK]��!k�L=��}�	���J�h`��iXg��}��*.=6��xV�Qk��*F����Se�b��+�ձ�������4+}B�m}���Wl�j�1a�r����5�H�eqqe̱���Bb�kCg��/wX~�gB�>�6�����[���R������	���}=L�)�ަ�p� ����i�����/���<*fiʳ���3�xd��P!�:��K>��u��Řm����d���xN�и�⻅���,�^FJ�e�0�$�����{ڬ�I�zUM�j����uB�nH�F+����Jȃ�2��P�E����]��*Oi��X��a��Ф|%-��>ͬ/���{Ü�IX�P���`��V/���Ck�ܑ���(%���7�u�g�P0� �#��ߥ�ãY����
R{o/m W�����)�.-��o�Q�Z��ӷ��t�om��:���m�çm`J��&Z؞	[��Q˸�^�'wY|�jIZ��m7�A����ӫ��Vp�}}�&\Ѕ�#�B��t�Ô�{kq]xgZZ�B�(��d�����)��n�^��	ǫ���;t1_�IcA�[<��^W+��Oȋ�W�M&��0������&����X}�7�Ϻ���:a;��FL��Z׵m��kR�gԞ��*X�.���2�aڏ���.�U5.��������Cg��v���7W����_��9�����43ٶᗈ��i���J��eX�^p�`��L^�3)������>���t�Zq��vȊ���]^�'O]����j�KirP��t/���J(�_�+����:�5w_Ow-/g���_��{՚i�7Z+�0�3h����>2�Z&_L%^;��{H�VzQ��%(�~���1Z��u���h<+ul���SC��T��`�j�R�.�]�uR$vXG�U��޺sRΜ��j�t�h[��o�:�9��O���hTF�y& ��B_R~ms�����c��������}�����I?x�����k���^��L�e�.�"��X���:UW�3H�����M?.���<�6��Oe�~�cH��~��/9_�[9�e�����jym)��2�1��CqBY�t9���+9���"�N�}k���3@Ϝ�[اD�����m�W��p-q5FPt���j��0u���.���=�yƶ�2Z���I�ivŰpmgc6���.m�f����b���x���b�X�9��@���L�� e�$"<�*"��Z�����.�[� .޾7���yu��j�D��|qM��=�}ӕ��Y��1wp��K���!z+qr�6�Nb=��!�xlN:���0��A.��FJۘd
�fV�D����aCOv$��.��˻ɵ �0J�er.��yMnq��E'!	٥S.��&� �Va���ę���W����9�R�q���\���<�#����/`g���P�ܫ��羙#F��3$��]�#�Ε��q9LW*��ҭ��u�����2�_)S�]hZ��s����9�CC��1�o����;��rM��Yb��z@� ���K�YE�+�c�n;sMLX�S�iX���$
H���{�����w0=P����)��ndP��ş��������GiZ�[�qU��Qו7,�r�X��ڻ��S1��)���}d`ۺ��[�6�=S�@�
7ؒ��#iv��qyJCc$�z1K}.uku�Z�r9��D�ۇ���q���.�7��Zn�}�'���3���]�t��
���W�O�)��AX_
����p�%Op�u�X/�8��n�P׃#m�͂�g`W,[�G&C�I���x;G��z���a���Mޜ�t�T��MXgm��R�� �}�RDq�i���S/�������g{=O�����������-�Yw;v�|9ޡ,��ddZ�3�Lõ}@G�����cs�����@��0��8(ⳝ����r�:���Rgm��8,X�ĭ�Gf�@�z�o85u����GX�0��ͦ �����\����2��](����zqyj�.�#�:�k�wn�X)9���meXs*o	���{�������֋�f�H��9��7s���\��x����b@�Hr�=s�(P[�Ē����HعR�Y"��2EDVu:ysX5k�ÓI��lS]ѳ���ᣚ�,o\���0��>��|(༊^o$Ѳݙ,L������
P�'�[)W�pƳ&
$�*�A^�j���(�2+�{��溉�N��u)Q:W��I2���u�;�u�K W��F��w*kwΉ��լl�"�7��[꛷��bDq%\��Е��W� xT�3�N���K̮�}�؆� �:�������Y̌��wu'8�Vq�{���ێƅ��n���r:4-7�y�6ڳ��s�U��`�g8�1R���S �u$4�ϰѬ]�6n�H#�ͮæ_2d��l���^m�֯�����5�"�jic %['/�gQ�r��T��
�9��xz]����D5 @�TA`,�¤�Ъ�T+m��Y
�*���AEDP"�Q������U�DcX��(���f%Qb������P��ʢ,q�J��fYr�.5EEEH��#+QEPQT�+YZ�m��0q�eDX�Q�8�X,�TY"����J�,�2�lX
���-�k(��UC�D�Q"��U���DEB����m*��FC��(�ALV���X�R((��`�
��¥�X#%aP(��
�(Ԡ�
�Ŋ*Ȱ��X*���E�Y*����*����1��["�*�-j�kPQ���1����Y}q$9�z/��:&�;m�oU�޲�IÉx:���Hq�E��Τ�$�[Nq8�9��1�sh���_�|�oW��A���$I���{�
V����-�����A�B�8���z���ˮ꧆l���>30W�e�둀r���#��\���I�p:�*+z`dŢ���rI�^��{y�Q�|�
�W ��Y����|���qu�͎Xw��u�&�N�V���Vr�u7�+i(r-5`7����<��y[˰�kɞb�cۀz�3٧�qT������iy��զ��]ґ\L&��\��K���	�Ѕq���t�@���8i�޾���׍{h[U喘n�����{+?_���-[]~v�j�L"c3lʻ�r�G:>Kܮ}U<�Ȇ}�ق�i��rǢ�R���[Jo��y���e�d�o{�	�(ᣩ3=�V�}U�*�ԯ.\9�.�9��dA��X+�M �#�o�/X�0���Hz=K��v��x�%+�T6Z蕇�*�,��`w�H�=�a&�{��=�.ps�Wo��=r�8e?&"�V}y�&Yj+i������L�.���/���"[�����[�}h��U�^Q�)q�����6׳9J��4s�ƫ��� �]�c�XW\��LWX"M�6^0�hco*S�.5o��'�Nk����H��xݬ)�4f'�P�`����4����Jin�-�/��l�{7�?}��Ny�\�1Z�?��R%��H���@�b���KP����W�U��ҹ�B�mQ������ڦi�ڣ 5�%=5ݖLy,kTpI�����	��X�h��'=g>�gݘ�'�v�ǰ�!�F��{ق��c�⼙��q �Nx(��]ެ���X�[��'\��ռ$��y�Y�h{�Dl�a�����|����*������,s�=kc˺�+�x��ۖy�^n��E����ǂ���R��D�f5�"���<t7�`wlƕr9B�?:��^��כv|5��19�SO
�"eo"8�K��9M�k��GOb�MP���/3]�s8�֙�mA/.g�,~i�N�vZHTf��)�p�@����b��M!������Y�q��4�V�WP��V�.��|�>i�vA�,�;-IK��j�O:��:�(q�w���=���ޘ)_��@h�������.P��(���d���u�g�(��>�q`:�����ν�����]=��==[Y�ϯ�o�/z7���*�m��7�t+u��`q�S{܅�<�o�EV������ugG�^Qǭ�9���խ��܄�+u�v`�[��gE��A�P�;S2抶�s��@R��괂�W�k�S��g}�ky���掩��� <��g_ﾥ).ۛ�=�
�uh��&? ���%�W�fl��C4g[��XC1�r�� �o�J����[K����/��>��{P�^2��5�~�i�V�?N��|Fqr^�Ev�WY��v��a��t�ͱW>�q�2l�ܴb��yj+�i\X-"����DY{]�l�c�2�{;�\��n�3�x�R$�-��;��{�w��%��q�Yh�a�W<|��p��Zz�Ke�_.�����^:�=M)��Pŕ�̷w9C��X��N5�[��;��A[r�>�xf��u��!��`���
T8���
�\�J�iE7�0�o�SS�%�}MT�}S=��>l�ǋs�f#��\N���
�"ʪfJ���GWp9\jq�� -76e����o�C�;�{��8{�`p�dX����;�<W
	�c9��v'��̃x?!�t��N+=��t�1ǞUﯫ���#hi(~uD,Z����*\=�Μ���N����L�L��ݷؼ%��~���nV>�3�\�hP!��B�Y�K/���g�]|&"�n�*��g�[��ol�;��Z��ft�:�<�]h�'b�|��b�m����.���[m=�X��I�{�Y�%�<S�?u�i���z�B(�L�;��#��]m��)ȸ���������H�%���V�MVڧf�5�No�?V=�� ;�}Mn�	O����c��'�Z��%fB��qq��=��v�Y0�}�]�u\[�y�ry���"T���]z.�5�����s�`Fĕ��.�8�tej��t�݉��s��p_�lh�a���
G�"��͟f���}��9���:�Ժ7�y�y�1����{��yj�.7#~	��Z����1w􏃪�~�;(����Z�MZoO��>oNi�Jz�U��8r�֥��r�ڇ_�yt(f�b�VY�HG����2�c�珗3��#��-��w넑y=}�{�״m2�����4d��w���Q�S�]Ua�J�@;j��`��������x�IcuxZ�C��E����y�{ґ�}�v��9 ��fS���U�Fp�`��9��^�1:��񇼜�p�s=��@�1��t��ʫ���+Cv���VڙUJ�΂Ł�P���(��󋃹�_L�XMP��#샵̻�}�`\��˰���U��az�O>Zm����O} .s��"=�_�Z6�˖xCy�|j2`��v�c�V�_<��U��t��eh�K��� �E&�pm�/2�9	ȕcr*W�[X:wnjt�+�OIJ�l@�DE>:��`�qr�3�媹�V��SX�G� T�Z����׻�|�֬6Iȭ�;�SέZ�{+�>-��&n�z����U���50�:�P:��L���ؾ���{�k����1�h���7�2nؚ�6Q5���f��Âq��YC�#�B\��֠��P�U�oL���9K�Tp;w5{�+n�}�c8=:ߕ�����s)r�$������-���k��G��k]�(kXy&t?;�����%X�,9��FIy���ؗ=���s^�ZB�vP��x�� 3�$�B�Р�X͊���N�a�����A�B��x�9<=۪���풱cX'�L񹂡����$�Һ�GR��p7,?��8�Z����pW�sw�����yl�[��۱�#�k���S�Z$�y�b��I�|�2t:�!�KΆv������IO����c>r��O+yve,L���c��9�[�0��޲�� �hQ�+'�>4���O��M	Ȟ�\I�Ϡ�U���^A���['�%<o}��%���[-�o
t��>
��#�vR�oϷ�b�c�x�'�`^"���n���jz�F�4�^'=/r��c��:�c�F���ۙ8A�����Oy_���;�,���$�C#�q��ȹ��:e�\���j��=R	ۙ�
�������ǇvW��Wv����i	f�;��C�\�;�v+�:=hc�"����J��wWwgC�:'%���R�J�u�̌:��>~{ق�x��ܱ谹u�>{-�~���nWM�i��~���7����)Z�0��x$y3�,�ˮ�W��OB���t`�aūݦ�R�iM�c3r�s;w��>���/�Q�Z�S�Y⥇�����>�
OC��<S|/2����T�g�qr�X�Է��}�>��e���"��K֚+L�Z!���!�o7���z�P2ة��8���E}�v	�뼴��Եﲯ���Ї٥˶��m�1�����9Vqc(_�q�]}��@v�u��Uݏl��Gt���޶���ʝ��$l���K��H�j���{�c��W�3�ّ!y9�Bz-�Q�d�[���Ϗ��ih��:g��_t�����C�����q	^�v���+yc�+��>���ߧ������ʩc�k�L��@�J%�T�k((E�*]�>�WW���Z	e�����yO�e逳X�9S��eLY������U�:E�t�x�=�m7����<&n��{�W���f���Jn�B���;�.��^����Cg�9�n���k5���Gr��r�aH�<�|��|�q�g�^���_�(t��$yPf��;l�p��]���
����+w��b	PNN�!t�k�N�Z�Ro=�|��C����¡g��t�O��g�(^�G���-$(Fk��^��-��HG��ȧ�:6Il�˽�`=�r���vZ*èax�h�~D�q�TC6�|�uAG���˝��ۭ�hm`�Q����eE�����.{�6q0\	� _���Z��E�s�:��A�,!a�dCX�B�:���)����~�@z�z�V�{uq̾泯���yZ����T�|2�&?	����IArQ\/����c�:�(	��wn��x�V��|��h�l��^�ǀ+��H<��P��L0*X_{�W�:�YR��vf����rda_<��^�/��Dz�*����2����X�utg�՞%����Y�v���^ݗ=�1OooS��!�.���1Z`8�8�n[3��c(v �yA~�1]�w��S�v ñ�N��F� ]C�֖�.�Z��,�e���(|�X��N5�kz6�O�5w�����;+-ʅ�S�2�"�`��4�״���	��)������¨�)��n��'�|��q�pB�Bꂺ��I.���
B�Yr�;�ݡ�[���>��t_ܮ���o��v�w qK�x�^��B񈑋)S��)��'����]9�8mmXBG�(�F��	�+,W���LÊ,gk,��w&��=r�sC�ύ�f#�ݚ�am&��
�"υU33�˲*������xy�����$��ȷ�q]��g�Ё��c��"QC�ݠkz�b�\\YA3,g<�.�bU����b��5u5��:�k)�(x�8���2\�֬���!�uD)�C��vZq�^�37���n8��9��񷕩96�ׄ�~/�34��Xt����=�K��:� �����t���R�Vd��wN���^I���-�Xo�J̅��-=7���q�d�|_����)�$Ml�z�b����f�ٹ"ߜ�`��\A�lkO=ǒq+�փ�7���J����:�l	�e�~4���݊�3��e3`�6��w_E�s�).��3���.o��f7ݬ��I���r�Z�C�.�u�gҵS��u#��ߥ������jH"��0+��l ��[UM��ە�/�r����^]<�{P�(g��{�8؇����kj�f|&u�w;o>C�[���	"�z��{
�ʇy8�$o5J��������VU�U��~ܺ��tҳ�.�-{��W�����(ά�5N���r7Ôm�)h'�7����iQ�Y��ξ
�����kջ�D�}:�V�3&;S��rmv�҆f��gJ�X��'Vd�tWͷ9pr-�f����w�厰8���P���z���3 u�c�pzK��Z� `�ٷ��x��fޞjsB��P�%�d��X�*�"����w���w1x�P�B����[O2�ީ���]L���ώVf�MY��VژT-,�(h�(@m��Qd��A{&t�uYb�@��_
�׷Y�뼶 ����]�Fث7��^��U��ʪ�+����I��^�I3��y�����w
�t��'P��f�窣���L���aa?�¯��N�d��4@�Τ���͏�ɓo&gjFN�W��&���f���8���*#I<��J�{����M��v��ާ
���;x�����Qz��d�s�N��g�9��B�X�Hϯ��ql��5=zA�ez�#;� DH�h$�vP����<�6��rr�ǜT<Dr?{�䗜���)���z_�S�:���{-,U�ڔ��J�Q����g��_�>x#�y�1w&o^�j9�v����o��1h��x��Pؘi�JM+�/
�X���^�b���yYZ'U�+�!���J��ق�f[����L�9�{����h���������rzΗc�H9P��ආ�Uj1��)P;���tW,ޝ\�=M�8�͡�:ɺ+e����lE�� ��|26g,�eʅ�L̡ʜu���H���>��Ê�{�? ]�ӒR�ᎃ�o.���IP�JE�eJ�)m2�,E,{}�·��pX�t�Ň��J�qCV�c�G��S��yvw�y3�����tz�,�=����kׄ�K:���k;���K&�Ѝa�[$�(v��U���Zf|nc٣��t^U�P$�E�J��=��Du*�~�}�m�x���'9nE�Jn`���ZX�W7baߨ�.ݏ\Z]���zyU���B�����c�ar�N�#|�j�yÎ��w��K`{�z�j�`Xl�Wh��ߋĸa.??	W���2 �難�C]�>󶊭�i��U�{����0|�}})�3@�zȲ�_�X~2�,�} h���*1�m��hݼ����"�0zS3�x'���xD!���bee���"��^��wn��Z+��&�Y|r��3�b�$q���d���N.��O��`�P��+�׹d�0E����r�����#���P���x�ᦚV��o�ل�,kTs�:ߗ�4ڡ�(�����٬��>8�v;��!��C�Ģ�u6e�Q��F��S�����vZYɘa]}�yGn�%�Sk)��IR��֗�V��`�&^�K�����[�����мڜ�V��Bm�<�ǵ�L�v8v�0�nRy���K�p.�.�.��C\.��;m]ޢ*Ԓ���v#Cu�����4�0���:�,��15��6�Z��r:�6؁ay(U�Pj���P�	t��!gf�)"���>�2E@8Oa���a)�Oi끝�u���h
q����s��1�dW���[/r"�EBw�J�ӌ�KV���D�7h�d1 XVk�WVo��t�*�^+�M�oN�y L�[=�\�]J��RfӉؾ�͕��X�ċjkaX-R�r�*V�Ԩ�� #ל�Yح^�c����]B��b��hع\� ѝ�A�]oQW.Ng]���.�'
��ܷz��u��9n;����|Nm%|,�;[. yvn>���&�a,�UNJ������^��5�<{'60۲-Nu��6�RýZM��Nf�y4��XZ�!�BS�WŊ�6܂<�����3D�a� t^K]]�[���ӄ٭m�I�.�Y։bP1� p���]�+����]�V6�w�a@�Z�;;WRof��Ym ko��Gf�СUڸX 4͵(��
�n��5Ӓf��,���k�fY���n@D��q�&$ha�3,��鸞c��et�l��l��T5�m��0���цy�o���ʺ�.��[zp�1P��.�$���m�����Pyn.�X�'��p)܅�YXNDT͔Ρ���p\���C�0V=tڋ�3����H��.��yns"B���m�q.Ȗ�	u�c��vT[Z�]��|�͓6A�|��p-���ʛu�q�Ծ��֫��u�Q�p��)�A����3(�H\�L�\!�e�m��<���S�:��Q��B,-� 7�b���i7�C82�Yu�b6#Rk$�[M�o��q��Z8Ax�A,Ǚf��g�ԙi%�ƺYw���^��G{k���<����m�!�����C�K�X�9������w��mT�����љlʝ�ɐ	B�h�p�c��7	�%��R+3d(�.��.�� M�q����QnQ�e#6�n�}b�G�����}e����,k������dwtxo-	�S=Xuv$�&;9�i�D ��;�B��(n����pk�`�#J�N�`>���*�����N+��
R|�}�2�m����N�r��6�����҉�인�yΏgv��k�1ە��`ܱZ6�M^����-�8Q�+3.���S2�Y�J��3������S{;�y�v�ot���s��]�X�⺥'Ǻ@K��!�.�5��� �!��}2v�ɇ���������
g����QDT���Xb���F,6���)`(�X��eBT�`�Q°F�V
Ŷ��3-TH�(���A��#E����*1X ���q�c+"�R1U�EX���V8��U֤Pb,Qb��Q-
�,Y3-�PU���*�%j"��m�AeaV"��1���X� ���QQ��*#R�,�DUTc"��V*��j�UAF �����b*(�	.6"-k������""�QQ1*b*D�`�EX����-U���-QTE,D�"�DV
�B�Uk(*�( �,\���)h�VR��T��S)T��*�)kq*�kb(�H!$��B���3ՙ�No��˂��ٰݬ��ek�
���7oq9��N{#���m,�]�o9GN쇢��:kv�1a���x�N�kY~����6��E��>6���.!�DsV�f
����&g�\H02s�E�u�{����^��o�����+ �l�2��r�\�Dl�a���u �;�RUi�-�S�;��N����������d]Asbǂ�����t�I3߅��V�²��g#�Y{�j�q��W>�zd^��^��T7�ʘ��eLY<(;�偬K�N���~��u�W~����7�G��7KW`l���=���l���ixi�@;��i �r�} ��ݽR��Q�b㧲w�[��!���vZ*�Cό�h�
z�!�G�edת�qy��a�fC�p��R�=�"����D��-��0R��{�7�q0j�]{j���������y�P:go�f�69Bj�)�L�Ve3g�g�ѝ]�g����X����m�^�%���s�F
����|"�gWT>>v�4ASJJ���~2�����<<���_2W�u�����ϖ�����X�f4��Jֻ��ӷꨘթ��m5���U�7\��ޝ���� ����1X�z^�\�;Vr��7O#ho��a^��ܯ�����d�^�B�=�~5)��s��K
�W�o����M׷Σ�Z�m	;.n����.�U�}�(�Vk����3w�Lh�wM�O\������rz�o7�����H�ޏx�����y�G�wC�3�hŧ���V�J�'����������MM8/贏*�����`�>��Y�l�w3e���VK��c�|6�t�������������KmN�+��*�;�c�PşW�1�NP�cڽQ��{��'�X����߫a�X;��������G���°������l�a�F�h���ރR��o}~��@6��';������� �h��fv]�Bgu���Mî��}�"��,{��&��c��p�Y��a�bY���@��"ŕ�ł�fiW+z��z�F���nϠ�w��^���L�q�ܩZqdmġ˪!La���؟�� ���q�{���+K��iL�m�5�}��~/�34�ŹXt����=�K��>[]�T���%�Z������Iˮ��u�N/	�Z��Wc�Q�2(oQp���f�����o:��Xr��G�/)�a����s]�=�)�\\6e;l>i��FX�v�]�hm��%���_S(���P�x�̕x���o;�
הu�׹�eG���S�Kh�Cum V�Q���$�vp��%�0�K-RN�Įb�7K�l՝b�8��z�����q�Lr���� �
��R�\�""z�n������k�;EqџJ�neه�h��R�)X�L�>ͬ/����3�/�"���$�}ylRSi7������t˪��?R���$f�u�s�����%64q�[��s��|�EǭC��ɰ�a���5�z�A��x�!��)n�3���"O�!浚�$���P}Uu�5�{�lZE���a6�$�z�J�kگsl=�<�o�4�֪�}�7� >Fa�����OL1��_��޻�r�b������We�����1t�������!��lՙ�P�Ա劃#٢���tS/m���b���q�뫈��l���ŏV��U8�`�^�LtK�K�����p����&�R���W}�s���/�|����
47���۫6+��(zRXI-���	��ש��[����7ę��#!Y�F+2u	�W��ؚ�r��U�^J[P��w�r����ϧL�Úr�ݚ��Č�&,��|��:�8'�(��TG��}o���9秙�j?$u���:T���\��OL�^ק�[��ESs�=�(����a�+l�I�P*�	H�/�)�n.��7���j�=CF�쾳Im�,i!vm'^�^�%���c��_j���P�ȩ��B�L�i�Z$|-l��g�c���BI���vJ�u�ؽ+n�l�,d���d�7�.�M��ת(v�ù�UH�H� 4��2��+m����m�8�x��~�ޝ�3�Ë�&ݚ��{��s�s��tL;0�5�"I�On!C���b��/1�:Oi%����\��S����������T<n`�e��II�U}�P#��އ!a���#�r��f�2�A�Y�Ɂ�˱�>����z��˴��)��(<�y�$�tv���ZB5fyo�u�����Jˊ*�."FڞW]�؈���m����Z�2�r�[��}����mu�Q8R�L+����bt�M�:�2M�P�֑2�e����܁���]�KB��w���G�µ'�`�Yjpt<e�
/c�}~N�U�ò���^k=��w�~.n��Z����P5�1�D1�f|/i�n�E��';�����z��o��W����/=�����>Hgٔ�yU�&u-.\9�wӅ���:�-6[��~�&���W�ge�oˢ�\��I6�
,��h��.��������e:Kw3m)�l�����AcB�^c�-���d]�"����QS��Z]8SE�9*��^�d@L�5#��#ϑ�nEP����]{g�����t����m�k*L���e�;��n{ln|��hb�'�~�ZVN��4�O|�y߽[XM�OQ�lBO�fs�x�RޯD!ҫ�O}Yj+�R��@���}�n5�{��d7��H�zjD�z_�:N�<]G��2��̨fZ+��ܻ${4�{�~�{����(�4DgNW!j�0��x���&^K��'[��g.��9�{��"�H�J��G���r����KHv#y_׳0Vu�dn&fpّ!{/��F��^�]<�!ue��d�IL�|&Z<lK4O4�>(CH!��z�����d�k�����B�����S���hX�<���u�\�؝�w甁�ΔJꙍg�ɞ�����{��-�S�Cڃ�S��k�2��Pߓ�ZzeLS^Z5�:E�9��t����@t?v��5muSO�`�>�JX���lY/.%S;҅a�C���'��+��-��V�V�y���1�ƒ놴�L�˽��k܃>��/+>ݢe��^*�'���w��zT����^�k���jYK1��"W��*�˖� �᭡���t���G���v��+>�Η7�&1���M�_0R�6��Z/%u�\�<�x�.B	X��M_n�u���ը�����܀S���SH����)�[�����!ZH�u���G�ޯx����z-����I��GcQl�9�3�f��z���䤨v³Di4�y�:�0�u�+�|t�E]:�ݚ�T���mv��ep�S�sfC��YՃ�/�� ������~2���j|����o�����Ǡλ0+�t�����x�;������X`Wh�-ΗB�<��U i�X7���ɏ�z��졦�5���/�Ŀ��#��;���d��g�~�DL���l�����x�L^iV)Jv�_]\63EB��}�ĳ��fc��pt��C��u����=��ȉ��5������|�#���V��6д�jZx��.�=5Y�ifXws�+��b�7sS����yw���Rux��g����t�f��2�*Eט���h{J)D��Tkvԕ��7g��'�"�%W40N4;rf6�am&��5w G{*�D����v*�c�u�kx�9�j��Dз��gř�1�a�r�uH��"��W����p|�;��*��ƺ�1D������#�c�5 -�4���0<��ޗLS_;��u�1,z���DN�rl�zc�(]5�s_,��N�ŀ�I�v�z�e�¯#8��n���uꝒp�`[Z����㜪�I��o}=�	�WCR�[�b�������?=��*�9�TB�=8���[��i��KL]L��\e���3�ּ)Y��!�[��O�����vk�	�wG�e�`ǩ=.�!�5�J5�*��ꔺ':�B��ҳg���qOǎzf���2�s/c���:��,�F�#�-+)sR�>�}�"��Qk3��(_��6Ar�~�)����»�\��8*C��eه�#G�K�������YTڽ�ޘ�Ǖ�'��IH���ܢ��Ρ�`L�� ~��3����,��Q�2�Gn�����*��]n�	q>۷�)T�W��@�__1��\�-u��z�o̔�A��]J���VB��mC��x��0ǲɏj]�oylv�m���4�~�vA���������_���>\��=0h�|r��Ն50��;~DPGsSS��q���vx1=]2!�f&:RPڔ5xeXd^h��s���f!�焽6���W6�b9)N�ef\�:3F<��a�4�5��OT�G�]�3��H{Ɉ!{�mf詙W����ȩ�LV5��g$2��i����%hcv�]3\�)�����P�a�s���lӨ�	�<�ڥe�q�tܣ3�WV9�����n�.�rx\Mwں|��i�/>��S*�&�
��`�p�;�^��]9ZŊT#��.\9�-�n��C{.�#lU����U��ʪ�7�S{}�:Ɉc�5���jɘ�l	�FB�ҌW�2u	����V�:��A/%�Ǖ����K^�G�㨦v[y��;�9��� ��e��o�P���i�f�֎7�N�<n4�{���g|E�Ը	w.ʮ.�η��;�5E�gl�/&���Gӊ�����i7o;xp=�.3)�(�$�'�:,<Yߟ��Oe�~�U�"�����R������/=��o����d�&�h��I?i��(tW���/0�e?/	�ݕc7��~�u�zJ��'�t/V*b�*7�*#RRi_�_j_q�^��W{��+k}�#�^��='Y�0ua�2`~2�i�)Z��A�v���IW�R/��{�z_����n��0R���*�Ϣ��-aϷ��V\PۗlQ#����/�uޝW'��=�:��,vY8\�̙7��T�V�����CF��L.���Yi����V�'*9%ޅ� �{p�Z�Iǅ.�u0R��䇹]s���L�\�-�B����׷�-�s��r��1���wb���� U���g�dݕ���V-�	0�%��uk���U��t-�X�_�ׂ��CڼdX;����	��h�r�'�Ľ�[җ+ng@���3*����^C�j��ʝ�[�4���SJ���y���s��4%f"=�v�{�'3űtHh�Ur��p�e�~i^��S��������(=c�1�V�y/{����hs^0=v����v�:k�^HP����ȗ%�~~
n}~��A3���:���p3�ȃm�}Nfx'7<�գ=�7���TM���kM�V{=�2��YS/p�atG���虜�^楽^t�_X�+-EW]�qԛti^Q�2}D/)�'kr�OX���G��,������O�=�;�kc��dů,�۳�S�"��� �,�9Lb���{Y|�i���<��l�e��5�yr�x�X�����;}����F�6�L�z��<m����Ef�T��R��8A�xz�}������=Fr~O�O��h䧍e���*���ϦZ<nY�ht�6P��!��c�R�����G��C�Q�Y�tȔ���B�1z��6�@�s����k__ϐބ�Z�[�B4���2�z�7�\Ʒ@v[�>���	}N�P�[(uj�Wݝ�Q�+���0������o2m�h�:rm��T-���b���xЮ���o�-MQ=I림�}ؚ^,ώ͡�;�]�J�ee��>yL�yHiD�T�k8M's��E~��`_~�U�����˸u�}S/N|�7�9S��*b�{��E���ٲ��J���֯pzU�1�JS�.�]������}�'Ze���˅�˶{҅4��W�;"=S�GT�C��e��i�6\fg�{��� σt^V�&wΡ��2��}��^��Z�:�}�5c^#��#M�C���W�&}}R
�I���%�?9�XK�2:��������;��\Z�)�X:���0�`��Cּ�	�>��:��<xܼ�~0�qOvp��y�M�ƥ���Oe��x��\:lnmÀ��ҳ��}G6aǏ�RG�ʙ��U�z�0dy�f�]�}��E��X�{1����q�7���a�k�v1��-�c���C*��{����������*��GoG�E�u/�.����(d�3�oش�g�j䲮M�9o���v�AQ�k��cʮ��С`���Pn[3����=���z�+�u��P�ڰIn��Y@d�Y�2��{`!��ToL�cgʍ��@���v;.T�hf�G:�1{dL�v�V��)t�n�=�븱v�cb�)z���ʌ����mmu����S*N΍��\��컦ÒX�k��$�P=�΋n���*屔��K����U�
���ɲ��:P��}D��;�ʔs�[Q�9�
�:ۻ�2�gdS����̮�q�sUw;��^/� y�Wt�t�ȍLL"]O4ei�V�~{���[��U��׾dms��_� ���Џ�3]�(N�c(of��-1w&ҽ��qUQU�7�Rn%k��Ꙏ�
l�:z}����
�i+9ޤ��»�I �C���d���-Fe<��b+��dLpyJ�t�'xV�<�t>�b��q�'��qF�,Y�v̲�5��Q�J���{׬=������{�9���V��ks��]^��Yy�o-$�vٜ��$�f}�7	ʆH7].}��%�Y.�@����V�ط�S��wAE�u�9x�-�v���De� B8R�����٠������uYʜ1�˥��v�,`��o03aP�������v�Sf�\�j�ͷ�ʖ�KxS�0s9��_h�pm��=�m��^cp��sVtK
,.)#2�]v�x/�5���U�����}�ݎg��D�dR�Q䒭�����x<fHw=���e��%�'���t&�����t�c��FE��t\5�w]&DVM��;�:�A,�3:��ro+ޙJd]Xj�0I쫘�viQ*g�$66�'�b�g�n��1 �y�.K�R�B�o��wb���5)��N[�� ��u"ַ�f�X
}4�0�6<�P�}�WrܝK��֨@ʭ�<��)\��õ�Kn���7Eu4�h�;ñN[��2P�*��)Z�좺b㲠�/F5Kz3&WHz�����H�*��K<��:��9R�]���j�B�]�i&Nk��т�N�Ok�"�1����r^��Q��VW���|�ݴvn_rt�B�0]h��[�M�iN<���/����Cu��V�[�pȢ��v3Gu�)�s]h��I]|�,�`�ۥY�������s�31T8V6x�ǭb]�h�k7�.xEWEP�ڱ;y�#T���I�D���=V;޾�Ͷo�GZF����ʜ���E�:��r�u�����w�B�up�Bl�21;��c�;�i��	]:tODu�����|�V]mfw���A%TN��S2̬�Q��͔��>v��k�+役�f����[���0.�����+� �y�8wg1��plo�TɑVݕ�>Ycn�sb�w��)���0v;C�4�J�%k���h��t\/5,���Lv;��\��r�,`��o|��]���
L�h�9���o�g't��e�;2�Z�
�ec}:H�l�k��*����ϖ:F
�EUb�;J�J�4�i��U*1�� ��Q��
���"*��U%���)l� �"6�T����#�1
0E\eAq3*�����#"����((�X�D����b�#Eb���Qh�X0U3"��*#T�f5Q2�(�����E�Z�Ĵ)���QDQq���J�E1��&P��B�-��JV**��"¶1F"����,�j[-��(*���l�" �-b+**���KE�"��`�B�J"ʔYD����E(V�P+Tb��U��b�2��q,�QU�b��+c2�2QV1E"*"��q%Ɩ�DF(�E�6�X�ګmP[mJ���F0X��T��QUUPUb� �mC-UJ�E�ʗ"bS���UF*�X�A�KlYV�1��QV,Z�K,QDˆQKs
9jFb\��&Y`� R$}�6u��VӾ���tX��ݡ�5����e-ͥC��Ҋ��xu5�R:�Aۚ��o��i�7����q�����7����l��|lEb����������Ǧ��if!�W\��ke%�/���ע�\�^���=��N���l�G����$��U`�}J��sO���w'X����ز��Z�ɲɆ⚜^UsBqC�.ǋxk������EU	߶��ԎJysz/{�����4���j��(�}N������"��hm��kz�`��~=8�u6iK~��w�����y�Px� ���ֈ�f���<o�d�r�D:Ն�V6=�;��w:�<�o� թq�閂fh�[Jdۄk^�X{)�Ӏ�+��3��+�hȳ�������{ϲ���4��#�W%�R�*���t^�u��,7�+0q{<=L��nϵ�����,>,ב�T;be�+�D�ܖ���)x.�5��nE�(�tbMz��Kq��
�/sB->����t��5�]�9�тT;beم�H���R��u�)�o'ط���b�c�z���p�oL��Z�`�Z��:e�C��/)�D��滛P��m� {�N���ʵy�b��95���:W�W	�>\�U%���ɦ�dL�Kʻ�`�{z�w���ji��顭�&*��[֒�'\W�N��I�X�E\��R�jm�h8�c�k���W�b�.Ș��NL}}����ܬ���x����g����q�L�J%�*9c�qc^KG)��*E�+��=�&���+)�.{��ӣʥ�*7x�ɸ�#��/��a6ڄ��Wx���.��Th�т��K��V)�c��6�mX��d��X!+M�ь�Gz�=V����ᶭ��21N��oz_/R���RF}�lȇ�`(v�%��/:��'\+4Up<F�o>!g�a��g�x�����^�g%z�/�z���y��l<5����ꭵ���,�I�L�a߼�8���cCOR��qXw.���@Q���a��Vlo���V�k�����b����E�f��~���%�#!]�F+���&���zlMYA�iP�.F����s^|КݿuF����`�\^_L�Y�wr$ru	垔L�;!����a�8֘5޶��}΅��6M�0��@I�O�Wg[�G w.j���L�o������Y�ҥ;�56����y�{��ɞ�L�i� E�0I�Q:p�<Y���jyU粳�'X�:M��/��7��ǋ�c�e�1Ic� ]���'���F<��<�_vM`��^@f�����U��Z�tV���u�1T�wNk6<9K	kE㐒{�Ǵ��)ǝ���e�h^�-��SN�0EY:�e9Vxn=]�r��{�e�}jm���k�9�wo2��Dfs�ܹ���Kg2e�����D��#Om�C��������q�i��6�|x��Xn	W���2��Ϝ��}*7��Cs#_II��ڕdOq-\*Y�	�=�dӼ�x��qWM����ɓ�x씭xc��XyL��IyE���mU�]yΧg�Z�b��u�U�[b������f,=ҒA��:�(��m��:����3^*�M�&em��Ih�r��7[��-��F���W�$�U��M_΄h�_m�Ozj�N�e�gtYL�����X�zא�զX�tQ���
Ԟсk�G�e+���j��zvƷIf̝��ڧl*�\��_��s}��QG\'Ֆ-�q3ĸy�sƻ5؇:���o�Zw.p��Ooy\��։�c�a�i���m,�zm�ݢ���W�w'�g�]�2��Pǚ��
η��쭭fz]�96�`���ϩ�����߼�}q�S�d��hfoy��]��Y.�[���A�>� ��*�_a9�H��IƸ��x�Rޯ}�J��%{3��|j�І��Y��*5�j��{�{�f�ke����+� S���h�.��fE�Sbu���暈��]��c�& t�� w91���'�;M��5�zr��r97�NΠ,Œ�}7�ɳj���]����%e�go%/09�����v󩹎�m��>ի��"�X�kpUivP`��8����{�k��ۗ�i��;D�s�l��-���l*���V#��U�>��Q�L��=5�}�	�uY7�o�Z��~'��ПMv�FS���H��.��h(	:CĈ�W����s���)��!�]�Oږ7�/�L�9ࣗ+���%3��:%�&�҈�!ϐCLh����n~��׿���®�w.����Z�*�R�Z��v�9ΔK���XW�YV����/ގ#l���>��bg�C�����Z�L�,�X�Rг.Tœ������泒�A��E9�OKN�*�mG���|%�k�^\/�˶{�J|[5+ꏩ)���}�q�v�_hpQ�[�d�U�R���w�X�r��/+7h��0�T*tⲧz�ٛ�0�=��v�gh��q}�uQlnC�
�WI�_T�Xɕ���]9�M>R�R]~����
W��i�a�OR��+4EF�k�Cֽ�xm�</�{�y偊a����d�-Ĵ��ҋ<���M��ԕ�DP�w��Ru+�ɣ���\/y��}PU��2I�5���{�`���7E��1?;���E���A�0�5f��Y��]��s�N�C��՛�l�1p�75�����.�GL%��t's�����0l�5,}���ȼY՝p��ڄY�M�
��EFԚYU��&���Xt��nd2���X+�_� ���ٍ,��q��}yUH��k��l��}̎&��?Mi�#?���Y�m��|dG�vX��d{ �q�3�6I�ky�οY9�'\�}�㭡���u%|�R�.��j��3EB���Orَ�ٽ�'ܫ��F�.觯�7�k��W�ϸVZ0�*�R��kO/��t=5^��}mj�6o�{��t�˹>T��^�^:�x�Zj�Teҡ�/1A?TS,�o�ȷ�h�ng��J}=I���Ɇښ�^��8��cN���[I�`�D7xzoL��8G���2���K�"�W^°�Ʀ�l�m�:Z3�c��"�aݢ����b^�,��׬w��ŗ�
���p:�����tP�y9�ܦn��Z�e탦�
��h��*$z]����CaJe�)�ަ���G�Iu��S�w]�͵v/}�3u&'��S�e�����3Kȡ��`���]ﻫ***��$����w0����&^̳�C=�Xu���t\վ�uͼ|(Ip��\l�q@Y|ކ��M�K��P�8;�b�=�N�Ug�^7Q���X��Ĕ���3�u�}�oz9�a���̓@�]@���Q+��vT�_z�]�QhG(7�_{�|I=*�Z�����{��@v�.>j�rT;be�+�D��X��E/.�5�ۑx�������7kw��Ǘ��{.+�>v�}!�tE�L�0��h����\}.���K}�N��u^�T܎
�]f|s%a��g3z`��ʄS�lr�Z�>;2�~��^���^��=���M����go���=�0��P��d���9CA9^kR�)�����rݪ�� �1;�so����N�7�xeM�>�2�L&��$��luCh";kW�En�޷�s=�VLw���e�����a<��~�__�����FK�2�g��j?��^6|{�Z0J��s�����藃t��˨�p�2����q�"eúu���wi��<�����`ϸ�v���Yt�@�n�D���P�e���څ$����մ��2z�QeBVˇ>���B�����m`��e�xo����<2,��[#y��x�o��M<����KO�QB�Km_�^���vK���U3����Ԙ�q��]֌sip\���~^m{���5�4���Y5�3K:֝g�ث:.չ#s��n��JX�^�X��-|[]��淕w�/�+L~�������q�I��FB�zQ�I�#+O���a���<�$��<�o4Z��Jvy���B��85WÝZ#WdV�ڛ��H��:��Ͻ(�c�C~�5�xZ�*�Y|��¶N>;�e�*#ƾJ$����2����x���<��B3���OGd�����>Oob�j��ߕx�讹9�Z��� �e.���۹���r^dܲ�d;wY��{�\=�U�"��?z��S����,�lL4Ms�I�8��(8�8
�����Զ�w-p�Go~�5z�9S��f�
���H��RiU�mnz)v���Нdu(C=_?q�/�����g�r�`~2�i�%+^��;	��k�팱���9������Z@��uKi�rñO7e�8t���\P�]�p9D�[���lO)�_vk�Lx���Mh^�J�;��R���&oޖ�L]e����iO/_$Q�{�ms �E�躓~����xz��ͯ�!]#�}��Z|+i'�x*�x����]F,�Lc�l�O��J��Z6�&��U�f;��T{y��;�k�&m^ z��:��uBc��L�/���l��Qwd����JJ=崛�]->�r�}u"��F\���ؗw�kr�o*���Y:�,@o!�E_l���Yh=�lv#������B��~�C���D��=��^�ۯ	�-��J�ȗZ�\W�xf�5ةؚ�v�<Þ�Ӹ�2��(<7,z,��oe��M�{�R�a�x;�|}),� �E�O�w&�,����AĵjǪ�d�x�W��.�3���s���Z3�cM�φ���mG/����|o�=|@��g|I��R"����6陎��`����A�|���j�}=���j{o�'"�-P�ErGԢ��Z�a�9�R%�����&0�[��]��^����6�֙�f��*�Yk����f�I�*+n��L��禡��+ޣ��p��n�=�����2}���>S�����k>�H�˴x��M@m.!�H�j��&�}�6Z����ZN<��\1Hn�}�8�u3_Η,�+����0��ȴA���e�(�u{=/<���d�����rU-�d�ҫOyx��1Ǟ��=P���ŏ3n�݆��=j��� ź�GViP��>�~�u�T�Ӏ4��^���YϮT�\B�si:;&oI]��Ļ����_+|aC���ʌ��nM�W��9g���C�&幼���&��p������n�i��e��5:�֢�X��9g���e[����3*�j��z4�u�g�l��y�rCw�v���d��,n�h�����wܟ�m=}m�[�CF��Af�a�����m{j�Kxqɲ���Īgm���ou?qn�6�����,cX��"�:�ZHSf�+S�2�뽊�k܃>��/+u�1u��6��;k�Z�d���e�*�&8)�$3�uD3c�������&}W�\�[�vz ���l�=��������n@��x�A��R�r+"R�z�KS>�+4Y�Gw�g�p5��R���`����D[g9�t����>��p{1��/ug\:o�͸E�z��Eo�׭�˄^�g�:����+L@߯h�O_���U��w]=YI�������X�µ2���2I��e��j�yD������k�h��3㦚5��Dv��9vF��n2����K]@P���nc��x��^�Ca}�mE�Ҩ�
\E�dyZ�pTX<�8�}�l��
�&�X2�����jǇ��P��.wU�3a���W
[hZt9-,��."����Q�a�!�����Nr/��<\����Rǵzs�=uN��24:8��Xϥ"�E�ղ�K�P��J�H���C}����l�.H�Ae��=m�a�t�r��[�I\���~�~��԰Y阧k˳$�l(��?d��}G��H��U_)��yp��1!�KDQ񗺆ڛf���;!g���Duf�۩'F�urn>�{r�s\�<�5Q8��KV��ԬM�Y��a����U�ЫrW��(����n��4�ޡvϚə� �0��^+cb�Z��n)��eo�ݮ,Ƴ�a�(���<.�
͊�N�t�6w�y@R,YL���f_��0Ӫ������,��7�����g�׾n�"ق���ɞ��;�H�@��`��e�L��4�M�F��/oǽ�9�g�Dqq��7��������3�3fg��o:��(PcS�Rk4����po�d\���}�j�;z�qY%7�a.����/�E�8%C�&Y,�6I	�\U�N.���[s�bw�L+e���L{��):�Y�G0#rVD��o���՝%C��˳?D2:�Ѧ�UlP�H������n��Cgٵ����oz`��*V�c�֌��be�*�޿T��������ի'ޢFj�>�w���<^����sz]%o��V�7���ʜ��|�P�S���i�Q;���`A�X���QG6��[�:���Aq��a5�rĬu����<�<hSM%o���cS�S�)vx����GF�X��Z�b虫ojLHjb���u3�#G��UM��*'��Ss��Z�ujP�z\�s8����B��O�i2t�Yx��z��J����G9LIr��9�ؾ�'�p�!�?*0.�{�W���u�諫�z�T�>���:=]�����U�R���b�)6:˪twt����hf4�T�Md��2k��
��/��8���u�X>KMA����x빗��k�\��Ɋ/\�u� ���.����(�)>�ʸ��Y�gpm����S��Qk6�/xR�:J���Z�LDyQ�ki�r�fr� �sln'.�Ν�4(�����4��s��d�a��%��]n��Ň��}O 8(u��4O!�).ճ�^����5um���;w*M�Ly2>�,R|�Q�]3ul�8,�c{��xҢ���:=&L�v���Q��P���aǜd|�9g��P��Q�s2^h���S��n,'�u��̹��<ݕ�3&8r�ױ@��_� �n�_W]���r�9V�*"�U�r�*�c�׆t�-��"�/�}
�6����������TH,BIʙH�JTT��rh"��r���ǿi�v^n2�ǁ�F��ǣJ�k)�b��V�\���Яd�}���1I�˸l�Ա�Kr�*
���4���c������l��3�n]([�n� �R	��К��V��S6��#�N�YT7gP�t�J긖���Ys��kW.U�r˦�N�{(�T;@��� �齼�'t+�Z��y>�{�n�!��_:=z����|�a��fBw;804V����F�rc,���n�xRĒ[4�vYӻ� �|wǏ��k-IFr�nVV��ie��u�7x�Ǜ3��L�����1�Da��ru���c�X�v�(��5��2t�:��q�$����v��}�����]c�\��q�6�
���Zo@c�MS$k��,�7�Hs����۽�mN�eh=�Qv�E]:�V���"n����'ؘ�_Z�ogZw��)'Bm��ME	��>�h�%|l�=��Y7�R��B����̢85��.`ͮq�Ճ�ONAgPN��+o�k-F0e;�G���u1�4H^�h��cr>R��p�e����;x:������(?	=�׋ɘt�kJ�6��13ǐ�����͗ك3���I#�[Gb6/O
OT��ZԷfL�T6PmA�ߘ��X|/:�m�0���T����ֱn�6�T^�ݫ`���-F�P�T����%��ܨX"�24�X��wa�z��� N&v��� �3��kHp�0J�r��#E2�PA�`ּ,b�l7�^��ա��m�r:�Ղ5����u�JC6��W���A��X�]�4�{�l���U�����e�j2���i�o��r��N�	F�y����m
�`8���l�3���6H�����/���X��*$Ucl�bLh�EUj�""�b����(*�U��J��!��LblA3,�%�X�[ls\B���j��\JF�QUE��D-Zո��[j��h�R؈�Q"
���U32d�+Tq,�(�[mX�j���E��Lr���(����-
�kX��Ң�h�-*�A2�DUa�Qc���KC*�1E��T������¥�l*���5��R�����-j	2�ƱQJ�e,��Ur�X�"1E��Z���b\̉�,�V+�(�R�X������mq�"��%�ʈ�1\lF*8�D�%Am�l��,lm�V1���*R,U�s1)r����,��*��E��B�\�YX墊�TEr�fe��G-U��\���AdUQk��"�\�1Jĭ�1[d�������*s1�j�J�q�jT��_)ӝ�zR�&��mF�9CrY�1=H��sǧ�L��y�й��)8�=ʓ�雞���DY3'� ݷ�Q�OD=���cWw_��[�\�a�TwM�ΘՑs4��j�;��4`�:����
Tw�Vlp��[�13Gz�#��ln�����gF�/W�	�m1�sk��OG+v�K�?ID疱���&'׶�ϩ����P�Y5��N;:�x�|w�ڲ:oh���oo?WZ�Һ�B|3�y&���s2R���"�A��*��܆���'vn��;=}K�9��I.//��(Ix����F+2u��^��؜�R��g.[xš8N׶t�+���d�;K�٤�js�T�����ő'��y�F�ӫݭ���䞘jK�[ۙ;Ú�q��a�֨�Sq�����m;%[��ÏO]�ʔ"��a�fv�&aO���~i�j�����v�L�vû@��0I�=>�ʝ�nh�ٞU�|o��ֺ<�^���}*ƑnG�Y��.y_�[9�L�a�0�49�$�#���+۪y+=*���y�U�j�*���L�����y�?(^�TŹ�pٹ����F���ܞźn�:����^��V�y��+�(�o��ܘj,�s�n61ԃ]L�\��q�o��!J�R�$��1��@�}G�qFe�<��+�Vl�l�j��0/f��·�:h�ۓ9����4ZF#�.�<X�l��|��7�>����F������^�׍�oh򶸳�d����rJV�1�x*ѭZh�^����6O]���/�=�
��U�[l��b��j���ZJˊ�˶֫ݷy,�K���0��߿d$X?���\˱�޴�7���jP�ߖ�^|N����A�Oh��[>*��A���n�QК��&I�P��Uס�Es���{(���V�$��C�{�Bu�{_����^k���.���\�����Mj����k�Y��~��^�{���&bv��l�U��uw^�h?u�f�x���D��W%���vP�ӧ�3�z�SE��\ٷ�QA�o�s��->J}���ِ^�"�]�9�<\M)�L�{lo_;�y�W5��w� �3Ŭ����R倸� ��������N�L�w/�Kz��R�V��9l��<C��V�g�k�JQ�.�V�^W�/Z�W�A�C�ӉMH��p��[:�F�U}~'�߷�ϏT{\v3Z�L�{+-rJ��>�Cf^_B}cL8��Zk��=>�*m#����2M��#����b�^�6�<.���m��Ɯ�z;8�V�����5e�0e	��r�\�B�W<8 �-�CTU�(Ҍ��V�����Bw���@�u����5n���s�6��e�gk4��}KOA��z�i-�SEu�����e7���vK�%�j:��#4��2���6���K�v#�w�˩E嫽ގ,�uW�N����o�ّ!c'<r�wz�$�K�x�D��J#�5���=�c��Q�m�wN�ó����ɫҫOyx��㼵�z�y����LϮ�W�5�w����{i4�UB�@�={��ϝ6���:ׅL�,��˧�bJ��[�c��lf���v�O`���h�Lru�U�}��~yIo��.#�w��R�+��
�'۶ܮ��-6}T�KL�R�	a夃er^�\e�l[�^�mtw]��~V�/ڽ.xI]71�7a�𺶉�=D�sΨ�lvA���&}]R!��ޭ���qg��z8W�=��ܧ����0R��$VD���৩`�l+4Y�Gw�g�_z;�㌷v7�P]A�Q�_�h�R�浺x��cR��of0a�ϖ����p�zq<����J�V�Tϵx�f��pǝ}�>���s�����@�qݽ.�n��1�s	��)noi7
l�x�s	�a���^�6k�m��,�'B��Wp�<��xf>��N�M[(=u�9W)��+x��Ƿ�6�;{/���������v"��Ȳ��o����B�f[=G�Tb��zN���o�F��7U��֝��fp��D]��yX��'	g�%S���"�;���}o����m�K���阳J�st�6;k�}g�~1�e4�����j���/u�;�%��qɶ�O\�;���;����F����4��-`�u���f�b�V/��m��cq�&��,���/�w9C��X��Nw��)��Yh���PĶ�Z�f�vt�U^���vD��°�����=0�m����U��q��.�㴠Z5��e���kԏ�A,��u=6�,�I-/n�����+9�Ᲊ�}��x�̜l2!��Xv��:�Uۄ�c�̚<3��#�'��.$2�ݚn�?!��nmh�ld�7���ǣ��n�'EU���^��5��C�BH��]�k�\��S-�즔~�G�A/n���+L���g�����lx_yA��9���2[�(��Aﵚ�].k��B���tG.�n�޼���='�>��<�ڻ��]L\|"���T;.Rj%%�#d|mT;���^iC^�r���E*ޠu�U�
�m���6jtթ!���gc=2��u�����ޝ��E��۷�GtC�v�amkΩ78A7�;�d��x!A���b����]LL�e�4��)�o�OV])��ֺw։ݴDuM\s�9����g�!�k�IE�ϣ��%dA�T�t����P�2�ß?FTE]R�$��[����ϫ�xf�.\Ņ���f,��0RV�B)˶���a׆�J�Xx�"[�d�vǮѳ�@�Cg8d�o���<Y㴡{��+}�����8�bu0g]��b��E��bS�+r�Լ�yP��i��`�,��߬�ɸ�4A�K[�6|�-��aS�u����I'��^�����V!�g��)yև|eϼgAt<��7��Tjy�yKU�j�5���5\��Y���^
޲�_Y�n�o�f/s�L	������	97�Ec�� �.��tPg׶��w1x��^���w����s�Qj+��Խ�4�W����j�4\c}�UiԲ�P�0xw�5T!��]ã�[������7<�hS	[e�g��]�⊾Vx/Ԓ����	��1P�a����zQ����L���-�ה0Q^5�~d�*�U�`B�����٤�jy�v���ȑ�P��҉�oJ�{Bxe����s�l���1���&���l`%>�z��m��)��|�h��x�c�Fvs}��{1�+���S}˯�N������fE��Dvʔ&f鵛F2^cZ4��8o�V��Ƀ���C��z�C˻�ls�u�K�m��)���P��w��'׬�s}םl�tXpN5ܲa����I��-�`�\^�x��w.jٛ�X\��1������K<F��62m�V}���|�v�L�v��W��@��T�{��wMn5���:�F�S��r_`��*Ƒ`9�g�d�<��%���e�N��&��NE��9��h�w�B�5c+��Lv�Fe_�|e��*b����*�����{�{4�{�:�F�Z���u+��v�͋8�>��`\Y��y0? e�ӒR����ne�\;2ϥ�Ɔb�0S7�H&5ȟ��Q9��ik8��2��ޡ+����.��{��������<�<��������O-�.X�����'
Y��w�r��[�+7�*����V"�l�j��6�I��[ʱ3�Z�3?o��+O��3_Y�k
�o+-�[�ڂ����ҵ�c�g���3=u��mz�V��*�L�Qޗ�yL�h��a��u����r��f|/i���Ǣϋ�x�{-���m��c�d�7{���b�
eb���;�V\�A�ڎW:�����]	�g"��$Uj[&h��F�ߨV���,�=�wdЁx��;���B��I�=�s|���o���������Pt_=x�xv�87su����V�)�էx�ՊU�A�u˥FJG6-�;��#y�f`��{�3�%|dKF���_l�^�"�\����i9�p�*&{~���6|ܧ�)���eu�Pذ�p�K�+\�@M��>�|< ę�������Q������������ �3�Yy�
�QYE5t�j`�z�����w������Sy��m��=��<�^"�v:Q�q��rbeA�Ftӣ�W���Ug�����b���O3�=����<+��0�y,kP�)��{��6��{G��7��P�.!�+=���Y����	j���@:�"X�37�lȐ���
5vWH)�ɖ��h�V���`����c�b3�T0�i��Z>w2j�x�!�8�ֽ=P�����G	�L� �7~�,�_�}u$/hp.c���&C��b��~��z<�=�0��_>z��i�Y�y��ƅ��<Y��B;�}Αi]:��]�������=�z,�׋�"����K�Nj��~��zU�p	BZ��P�A	�夅6k��N��˽��q^��8���ީ����3�N�G%��%��)��L;)�E�������[����X���Nx"�i6zM����j��8G�C)���eU��em]L4yY��)��3���Vsb����\���Z���
��3.v�S[sp�#%u�ejU}·�D��΢��l�/g����i�T�oZ3%a��m�R�"Q���p{ U���-�GWp'��X�2{��y���ǻ����=�����-0l=K �o�f���v{6$�"��y�W�:�MOn+Lr^�K��}��Q�s�LU�բ��`�^,�����/�l]��*����"��P����A}(��\\T���:���`���H����g�"u�Jӄ-����}��y��`W�ҵ�ǥ�8K8��[�N�]����#�o���\�+�27q�=$����i߮�ϼ�W<Ex&G���g�U�
�*�2��2�-GɯbP���\�;����3�\��g��{Ȟ:"L�*1�x���c�Ǎ׽8� �%�8�Pŕ��n�r�Υ�j�����T��أ#C8����t-�јFl��wJ5�� �Bb���asQ'�Eza0�jrq{�*���q�ۂf3ǈ��h��}�W�'�y���0)K����W�v]�W�u�V|YȦ��o7�=�U�����a�m�?O#5�2�+L�5�pn�ݘ36Ur{(KF��tf�	�:f�,Æ�q�e�Wr���L�o�rk�7c�j+�_6��b�^>��k/;G1'��I��[ n��p �q]�Xe^s�wJ���cS�6�����/��u���S�p�ҏorgG�����/Df�[�Z��),�.,��f_��0�;���|���ֈ�e>�Н��z�0���/k73m��^�;W"P�CW%���yB��;�ҘۄkZ²֩���Ӿh�����޽K �{�C�P`����%�7���� ���J���vP�{��3���_Oe[�1�~�Iꓨ�,G,7�fi��b��7�����e�͛$��.+�û`�~�Ep��!:�uϮ�4���^r�Y�G0#bJȃ�o��5gDP�]Q�M�G]�n��<�xz����V8	*�#F�X�x:�su�ǎ`ޘ)'"���[�Z���-|fˋ6�uj�ut�6����4�!��tX�8}c%Þͼ/�\z�;ҩ.},P���>7�=WWt���<���ӫdR)��.���K�g�j�~TY��\��+q>#k�o�cA$��C��6�����ޢ���ǵY��XL&6����#�h��j�����B-T����+��k-����]Xg|�>/c�z���a}��S,���c/�b�2r�?P.2�-�l�G%a�<to؈��⾥���į�4�p-t�ؑ��i����o��&��X��*�d�z�0c�����K)k�`V��%N��s�_Ry�����U��(��J�1���3~�dEX�(�#i��.=��49T� ���/��1��;%݆��*ǈ�*�;�!�A�^�1:���P�X&��o�ח��ơ��������b����9GgªZ�L�W���6z�QeBV�fC�oWo�D3|��T�߅�ɻ�\�+=I���ȳ��MşUW��	�1���䌅w���B>��?z�ݶ9����?sX���u�K�ԫ���k��#�N4'�rp���K�����{�O���<��P��Ӎw,�a���\���q�57[N�S�U)�w�G�K�8i�=�{.��O��>{<6���jj��G]R�!�O5<7u���}��\1g6ۺ�=�ϩ3�sS�}�_��cH��~����+d�s&Y0�������
j챎�%+��|�?i݁
+��bb��)����R�P~2��8��gK���S�.��xF��u�JǪ@�W��-/
�X��g����Z�z,���cM�J�vw�qm��J�7}���\i�uĵN��/�WV+m��b��-a��i">�����]�=�*Z�
��bX.�T_P�8�� �/�ʋDWz�i���];H3}�fQ�Z�8�L�B���-wd��x�IKą�ӏ�m4�[��牺x�;�1LJ`ѡ�M�LVia
����R�zK��Ld�N�'^X=U+���`�aZj�9��+�9XVܫȖ+�d��.k��*��u� ���.�wm�'�hI��9���.¬໦��%��ê�ުC9_�M�)����_]G�6�u,YX��F&�o�J��çw�^c���*�g"�2�+)�gek�}f���๩F��VM��^���94xi�of�۴PS�K�« �t���k�}Y�TZ�qo w�
����"DҮ����U�O}$��L)z.��*��)!�J;.��;u�%�U��v6�]����B��-�5j���wh`�3��'T�]�U��h�V�{��ѲQ�,С}�:&m�P����d.�5� �C�\b�e�GP� �r��9Wmw_J|���T��!q��G[�|�2fH��֗m�otΥۧ@�����[�6�/�!t�65 ��=�
ኆH�@�B�gff���:��7��h��2���VA.^��1��Kh���mrpܩl=zf���ϟ'�7��ybg67���C�bLC|�n�5Ʋr�r��A<c�7�Z�-���V��8�B-�a$ҙ�hA���T嚵]���a��Jz�[��VG[�,�@+eu��*�(�eb�/�(�V���BNI9]S��[�Ƽ�H<����J��@ڭ(Mzk��f���p�|/d�$�����w�����Y��q���N�7��;b���ՆQ]�Q�=lpD��\�Jwt�7V�i..1�X��l;6�N��]ON���ۦ�fV,�B�[o�ª��A�V"8]�AV�ة�쫾�2�n*�h�a�	��To��{6����;�$���A�
1]�ܫᦀ�U!�v������<VC�I�׏����9���7+�\!o��v��9��5zVR<�rl�]y�^sז�	��h�X;��f��#|�ӯ��T��5im�R���C��p���H���s*�\D}��>lfw&Xu����y�E�1�ys�ۯ�7mA��j^��m@¯;v����[�uX�J����K��4X�Lb�w�vN(#{�Z���ٜP�]VJ�夨E��T�K��q�HA0M��z.��ؙ�)6�Lبa�V�p�^������m�8��KnbScT��zL�N�Q�4�[�ӤR�k1����\;Zh�N���#�V���{1v�[}�!M#��q��AIfP��^h��'���p� NLQ���lC7s;�u.��<����<��/�	��V�Z�6�.ݘe�
��*Nw���b˻N�ѵwYRdR��KΔ��j�����y++!o+���w	��)w+Z56ފ)h�w�Y��곣�2ަ�̥�����Ɗ�s��XKs����]K�y"ȯxc����=X��F�7ϣ'�t��Ov8I��u����P�
)QT��5�+q�R��Y���m�"ʆ81�,k
��-�ī��1��*�B�Q̦1�XcY\f ��qĘԶ�\jQm�J��qS1�LFق�BաQE�1�֡fY1�&QV�[L`Tr�,b��̲��(���qq��PDUX����X�*
��G1��+�aP�Q*U�
����
5�S�Y���F�b�YEE"�����(� b�H�*���E�LaYm
��£h��h�
�*,�6�-Y*
�11��rZ�����73�W�TE�Q��P���(�L̘��9sT\h�Vb���\d+EF"����(��L�EV2"����Z*5�mEAaR�DL�a�UH(��).2�*���B�Z9�����
�Fe
��R.V��5+F�AE-k��dQ���Z� �	 �E��{����6��S��%p9I֭1I�m��&��Wqf���"K��N�xI�܄=�|��k�X]�JMp;�ɦ���Sz�Ws�u��^�r��jy;���I3��[QT��\�]�
�7L�N� ���;'���;0����s�W�&Â��ڃַ�mx�Z�3;��u=q�׬_�8x��+o\qVS�Bd���n'�C�X�pl=��[�����Y��ֻ��~t�;���Ԗ*�}���D7z�B��<Pz�Ǣ�C�m/OS;�a���]��Z�g\v4Y�eK�^�q8=<��%�dK�	u��>̀���dA�V�q`�`��q4��5��nj��Ō��zd}f���\6Z蕏C*�,�} si{�N��$��n�����`�H"m��RMY~��^w��X��E�8�iR����X��vq"�N�@����Ew�_Us�wؔ�e�,J��y��k�e{S�eC�+-r���4P�쥝n�����Ǔd�z��`�ԯ禡��ɗ({�%�v�f�R�=*���M@{�eu=<���ɾ#�Dv����Y�[Ɩ|wə�fD����
9r��R�w�#F��%�BR���o+�V���<:�<d
D�6��y{��8/(z����L����d9�� ����aǉކ�2��u�7,�96Y����M���#�6��M�x��Yg�I�3����;̭�1m']0|��ʙ�qId�r��S��@���u�Q3�m.F��Ă8�]H6̚�*������c�=k�OT#/{��R���߾���E����>������a� k�(��3@�=��+6����0*e�)�Ǽ�o�[�����͝�p�4���A0Pv>yh�H��P�۸{�Ar���l��Jty`���%�������wl�R�0�'��	o-$+�ٮI���Sy��
\���οh&z={�q�N�2�]#"��@e[Dゞ�C9�TC7�M�\��q�ò��/`|�#�}WXО~��M�"���I�Ȭ�2��pSԹC�Ed���������l���Mp�2�/.�/�[��oJK�Ab��0�g˅��雙������W#��X�)��|�ҍC�Y�o���f��{��x�����/)�����)������(V��zz���c^3\�?]�x��}nN��O�l�x_�.�xۤ�*�ls��w,.3��{M�27{�}�ƾ�uy4�,��]��򯮮E�U�ۡnl�I���}3mn��W�]
V),��j��y*+������eo��qu��<���6;S��
���N�=�z�j�L3��k7��W��<�� ��d�w��)��G�*���;��gf�7�<�Ϸ-�\�.�v'\�;��H���{ә��������'ۦg|�f��a����L\2(��u���5�nu(�U7=�������y���I�'�����Pł��T�:�=�ӝ�����+-?Fk�����{E�(���(�O����J�b��
�5�������'K�q��ۃ��w�+�v�p��ָU�^]j|�'
����߻.ȫ��X9��M}��'�5
T����ѹ����Om���B�!�C�;���R,X+����wf�;���:�����ʏ+�Ξܞ���͙�9�7�w�z׾�;P�$�@�ڹ(��Z	���iK����!�3��iU�t�l��q�	{~3�&q:���zfq���
?:��Q+��wB=���{�9s��%�����K��E���Vf�������(oQ�P�̲YI�u����*��Wo��TT��;������y�-f�nJȃ�2�����%C�
k3���ֹZ�����b}v���H�g��<\�����f,��0RV�E[�����_�����Y��˫�&��H6��:VsOݔ D�����<��8
��6�WB���U���;�b[H�@����h�yԧ��-�d���]�9���]�s�+ ��Vt����	�n�u,��-e�����w%̮0��<�]���ѕ����j���JgM�2�����j�����~��c���g�fˤ�w���HM�ĕ���m䝺�$��ȱ�%�r����~���*�,&�\LpR[��g+��c�ܳ����7��>=�����$Xs���^�csl=Fԋ��ڳKY���]L�]�#zv��mY\g|o���t�����6|^�h��7W�^;��E����Xa��L�+o�Zl-�ҶƬT!�탃����fe;��|�/V5�!�:�^�}a��p��lnN[��\!�--���T:���b�y&��8�;���uKz�%�U��g���<�E��]Ϯ�.����D��I.1����*o��FB��J1{��=׻��b���o��AϏ�|��k#.!S!�,,<����$�s�T�!�ȑ�
��^{�_L�#�׹���>�t�e��o�P��+�t�C��F1Hh8T�_�N��P{�T���]�ez�2�:���[p�zt�7�o������-#�ݠE�0K��TKł-�
ˬhP��n�_d�\�}e��n�T�
M��W��p{��Cit���rc�� �������>G�{��7�:���I�f��EuP4�Uf_c�V���EP���Y����P�D�j�]۲d/m��_m���KM��}�jv[�f���Oˠ�Cz�Z�ө�ؗ�5�J��_�G�Y��d�<��d�s&Y0�㯈�[����/m�c}��{H�@�{�
+��a��8;x#�R�P~P�#]���DA�aS5�j�����j�h�@��r0��Z���P�^qZ���L��=KɁ��BqU�^Wi�=�߻|0χ���t�a3甒�$�_�/-�,|�3���s`>��:�Z��*q��zV��Z�׏O��`�H�,�^yv}޴�68)�rǷ�3��!�LS��~�iy�՞��Zf,��O��M	Ȗ�7�[ʱ3�k�<��|��e	�k��+}�e�����hg���׵���u�a��h����~C�鞺ϖ��[dt��[X�����!�����2R^��_�L͒�j{c�ap/��Y=\wr�6��ee8�8ڃ�2��ΐ��t���RY�`�gRʕ��d�2 ^��@�fu����a���]엘�(=�ܯ=Cڰ�k���U�1&���-�9�H����<ѿ+�Q莦�4�]������!��cÝ\7�2�-�1B��F��[��4�~:>�򦽵�fA:9A.�u	�Tz4�,�ȹ�%dW`��u����:�O8E�ƻpGN�WL�2�=i̓6���E�`ŮOj3�^�0�:&��ư6�>��o�>{]�g'�^襽^w�9��g��x�6ϧ��Auu�}��&T����5�t��`���tG���u;�U��3[�&T<��!妃6�M߽a�χ?NdWU����d3�F�.1+zj�0�c%�j:����	��X�8Iu�bw!�����;��f�,�P�$�j�]�!����9أ�+���3���~��J�7gk�̕�|f٢}�D|
�͠�`mu���ɫ�Ui�/}U���h�uq�P�(1���/�/r\����ی��v���RB� �0��V���si�K�u���r���P�uI���}Ӷ���Y��?T�,�ʘ�L����t�J��.���=�&xU/����-���� ���c��q�u�%�<a���%��$�|ٮJ�<����T�^Y�]1t����C�W�/
g��yX7]�0	Xaxe[D��
z��:���h<+�>gVl�O���R�.��D<�"��237�
V��i�n
z�(|ͺ��a�6�*�5N�7�#��]��o��jI2�;��>���{s�؜$X� ���!ѫ�\�s��B��6��u�WK����ן��ꜴH'i�oᘧI����������Q�C��d��6^�)�.���G�2]�\�+�irw`]+���]ݝ�{�kzD4A�ֿ�P�X�	�4�g�3�6����J�X����i�=��;�g���/x������p�8Fh��0�񡞴�G:��>�35���?Og���Ә;�7x��T�:�,z|�<�\�,w���l
�C�7;�=y�疛h�w�b5SI���<�֙�Fn_��.��{q�3�L�Z1xӿ]B��
�Z�|56�����
Yu٘�g�vڃ�U�{��?�-���a����0	��u^&}²ц�zj��/||��k���K��$����"������8��1eif_��r�Υ�j���_���P*�֓�}�we��r��<x.�\�G��b�<�K~{J(�za0��NN/*��P��bYuoI;�:�̉�Ճ�?\�8JP-�<C��$�κ�+���L��yp�D�U��>�2���p�G;�ݮ�Kk0N6��Co�v�H�⸸�,�9�uA��������U~S���}r�Gӊ7���Z�:\"$J�h��@l.�^P�g!y[^ü�ϫC���ϻĪt�r��չ���a|�����v�

����us ��%�2���Q�bĘ�ۀǰ���k�q���Y��nǝC2��6��v�� ��_r8�f����`��up�fr�=��;壣Y�s�Μ�.�iv���\M�Nr���KӶ�����3�#�:}=38�Kx�:t!k5��,�==�/��b���O��ſSK�s��/���+3Ox����(oQ�P�̲Y6GfR�^��5�s���D)x���]Pg�o�܋�9E���s6��%S�!T|�����2���%N>�뺣�o�#@GbF�Z�3`�6���1f邒���EI��~M�kw+{X�cӟy��mZ3�P鹗p�~��&�*a[�~s0Z>�<f��K�ә��3�n�U�P�,U�݆�+�j^�+�p��Լ�yP���E�����|RO|�R:���o.�{�3��#���_ϦV��$9��V����t�Bx�Gp��S���㮴����]Ua��W倳��W�����c�l��������E����\��lU�En_�=�3�P�����]aq:�/��v��9����)����/��5�#A�bW�[��n�Xڝ�����j����U��P�Z2౜`��ME�q[����MY���FZ�y��W'�J�9���2�H��gb��#{kn��(�N��y�j�o���F8��$k;��n?Q"v��N��y��{{؅dj�7�j�ݸ��}HwYgU�Fs�4�Yϲ�5���ank�q\��W�m0�{��Zu���o.��j�47��26��7�Ҵ�
�6�}U\f����BM�R2z��GyX��j+�o�>�"��*z���&;G
��aa!��.vi;�u;����z�������q$�uoe�/�Px�ޔL�;�(sXrq��(�	TN��9���cy�G�eD���v��r�N��Jۄ{�t�62m�V|F����ږ��;�����P*�MZ���.�]ځ������{]�Oe�~�cH���޳�2K�W��W��J$Fg,�Ɩ��.�R��p�_ZY��>�x������K�ʯ�Z����v�{2hcD���a�3�l��P��#"M/
�GR���^��{I�pjkx3w��촰�
�=w��_��u�۱�4�`��=W��MS����TN�9MTF��������;fXH���Q��<����y��7�"��2��$`:S��˰�}޴�68)�rǶ��s{�rQ+o.+'8�̤(Ǖ��Ǐ������K&��B4M�2M�P��ʱ3��� �>=��.P�R��/���e���O���X�`��:s�*�jZ�eu��a��[���3e�6T�;\����Tg��/;'��Y)؞K��ൺ�&�d���o�Y���^��)�}�4�&��j[S�:��Q�Y�3��p�N��	TB�|��mC�ċ9[I<�j�C�ڶ�?-<+J{G�}���V9��c�D����B7|�Gu]S�U�|���lq��>�_����n{�y��]�k˭A^��aa�e��,N�Q����'�Z���n��i,5������J��Ãϳ >�ȃm������ʴ^{,���S����8�N�~~�>���Q��(l��+�R倨�v����	Տ#~��cqY;�ke3�L�m����~�oW��_P�T�>.�h�ċGּ��{лݙSϽ����E�xjjG&��,�T"�u7�ܩ��;��Cʩr���9^�7���.����Q�`�Bn}}�
8aihzj�,�r��3>S���ZG'�͉g4'ҭ�'�����[@#�#�ۗb�:�4��3}�̉��!�?-�W���[еX�5�-�[���� �Z<m٢z%��q��A/i��\j�||¯f;�*��)W�yh����V:��d#4sY��e<�o%�u��$�|���/J��9�w������섐�$�ԁ$ I?�BH@�RB��@�$�䄐�$�bB��@�$��!$ I?܄��$��	!I�HIN�$����$�@�$�����$�D$�	'�!$ I?�	!I��IO���$�H@���d�Mf�{���_~�Ad����vB������}�EI�z *@��)J��Ia�uT�������@* B\fQ٘Ƒ�EJ(j�]��릤ֵ��[eL���nκ97`��j�]�MIEM��u�	PBؘ��E��˹�9�:j�z<� @  t���M۹ԛj�ŵ
5����q���F�KL��U����{(�Z4*Mmj�d՝wU�����9{kMV�ЋV	caj����y�s��+l՚�)m�V�[f*Ȋ��o��yj��iae����b͛kB���=���[5%j�jj�қ5aP���[ʉ顚f63Ti���mm�z T��EP�jz%%%@��  � �O���@       ���a2dɑ��4�# C�JR�40�M4��b�U)��c� '�ѣ@ h $�@�#D�Ѥ�<��4��f����W�5��i�},�Z.��I$��4}�� �񱍶�����������@�I.��O���L$$�P�ǃ�r��������rr���"x�%��������82A�Bw�ID�����>��I'���!��䌄R�$��a���Y�4}� ���}���~�*�*�����*����(��������I!HIR�ӱ�i����m�1�����*�����*��-W;��$ǆ���10�W֔<A��.|h��'��_^�?٭���D������/�
��Z')ym�bm����W���!v����#U�0C*��l�Z^Y5����#��`Ӊ]��^[S�	7R��n����3]�fPu�%l2#�[TKOq<��+6�(�ӫ�Q�̡ɯ�����}�>9Dǖ>8M*��E�
��7wn���ҵ����Qf�{wE�7�ј�]�K
z ��Ƙͱ�A�e�L��ܿ��j�i�EԚ��3�&��Ht��kR�Q�l�@9��j� ˱��75�������&���*ݝ�op�,U���h`���4�n��M�a���W��v����raS���[A��{�&Zа�Ǖ�܇a�]�C��h3���9b��V1�b���NJ�	f:A�(]�+x�L�f�0K�b��n+�#6�p(���t���x��4�Y9��P�vK�m��&az,�
�b[B��+NdJ������+iP��1 �X0��(�YYx�Y�,��]�wDc�����:�]b���u(�K`/x��Y�N����;X�/���$"U9��O-Y�1WTs	7!����=/���;�b45j������m��"(�F�X��� ��x�WeQ�t�x�n���cN��+]2��:1U��je���~�l'Ȃ�B��M���oT۬t�n�-1�d�+��*!�Cȓ�a`B��a���9+l'7�)�i��T���d��^\[���V��ud�A�.�vn�'7���27���*��y�]u.�H�+Dm��H��)?����m���M�dn-U"��E��-^�Y{�#5��׶�ѷCn�-�Mj�k�i�˂�9�Gʽ�s:�3��h�F��õ��4�gβV@wj2��V�B��i�֯�'G\4�CI����-��Un��C�vc�T[SD �ݪ�A>�k�1@ko2��\�"�=��� n; e��R7���b�Fne���Y�����U�҅�֫�;�2����05*�AS�ģ:��ݑ�T��:��N�*�6�`Cmݐ3��xR�5��/,�!q�躸��e˰6k`Ԫ���SN�=�Ҳ�e��5LѪ��Q����b�5er=��XEkEe���j�/PB�4lB�R���Z�
����J0,T(%��%9�h/㘳ڐ2����YLn,a�:i�H�{�VV_-���7f���j�-5�ihV�h eMy�F�6inA���Pҝ�����D=�ƪ
A	*+X���7��� ��nxv�
����/(�Ua�QR��M��ώi!C�U����9L&;f��2�6^�!Q⣽7N\��9#��,��3 3,��Q���c*�c�Vo���[Z��ӊT:&ۻ8ݵ�aR�
��b�--hv�)�bU˳M�Md^�k@ʳO5����V�]X��wn]iP�5�a��U�u_جEA�X�E������ۢ� ݩ�A�V^P+^z���\ݧX��!*�Z'�u�����fZcG7B�>۷*�Ff|4֠�l'����)�J�҉
pܽ˿�` i��#��7��_8�sZ�Ɲz���M��F�eg�~l9D3GAtln�����4�GR夐��n>%�ոD���^�qX��Zce�n�\��.�:�5y6�Eu�1U�����Yn�\�WY��X�R9�>�HH���R`�I|�a嗥Ы��[���[�T�j�╘%�O6�dY��/VW�����Η�2�*N�0:�	��L6�&:(�c��ݛE&t�(�yvS�˟=,��~�ؔ��%���������
�1>�<����/�=k��,�Ph��o��v�"@��/qn�����ߡj��I�q���]����J���55��p>y��0�ƒ�{��]�bv�޷�o	z�7̪f+�7��/tK�ka�q)MΠ��k����װ�U$�h���ի03/���ypf��q<e���3T�&� �μ���-b&�;�.�c�z�<}�7ӂg;rl��_M6��#lc��Q�ɗ��^-ǹ�p�iջ�T��e�@[�Y�ξ�}��\ۖ{������큾.�Uu��/@��}('���F���taފ_%��C�0�?�-Wv�Ӈh�;�_5�眈6����UlT;Z�e94���`p�-n�FЧ-F2�9�>зlN^����.jzjM��*T,���:!�A�̜I��p�Lި�)�K�Ν%��8�a������.h���{��.q}58݉�yǺ�p5�1�h��Lm�+yyǍ�	��E�I�p�r��D�o���h�poT�x�ܥ\MH�,⓻�i��?A9]�k6l��B�3�ng�76�����5��Bĥk'��q�������|����Jr�J���S{����E��ֺ��q�˄��}N�B{��<"��T˲p�k:۵���1JmT�Y���jxc����>`DV���5�^�c23��:��re��歮�(B(�P��Ȉ�;��Kx��nӰ��3> *˖��\�KYB��K�*^mw`WOT롄��k��Q;amۄ�e^��HX8U�I[/SǮj�x�����5�1iGM%Q�5�v�z���r�2��mrYoi�y�V�i\w�0��s�U�f靡�dN���Gfĥ��]�<�oV�����t�BS���u�\$|����8�u��l��-�s��
v�`���Z�(��q�WG���'�,�Q�JNC�:JK�Z�7�ސA63��/�E�v��	����qv��.�������-�qo��)Z���W�Ղ�(��y�uTғ����dKyc�4�PR���{te;�[�xp�rv���m�2{����W�R��9�s�f�U1�t�,�qí>�.�h��=��J�d�v�FiĨ'#�T���*�탵�¹���p���|dF��;�at��]���.�.򑭳��8;�J*m�08���J���0�Cy�n�6'X��^�o����Xu|��Ysa5�3Db^�D;��M�!�{Y0�B�����&μ�5k���;�Ƭ�W��جjE��f�#�c�����o�V9u�)n:��vQ�
BG��U�BR���n�]��ѳ���-��V���d��I�%c����"�(�Ӹ�!�5։I�;��!�(�+wM]�'%�b����h���xCP=MJF�����Eg^q�ܝ�@��"��sNc��Cцfր�f�ԙ�[6Ӏڠ��:�H�Y`Q/J��-���f����S��
0�uJڱI�ˬ���qi�u}�<�{A�u�+,�ۤ�dΚEYQ� �])du�wij���raݤ�ܠĝS,d���3�P�y�2��^��.wr��zDB:�rF�tc�L��(�o����q�ň0kkw�)�CF��3�N�g]*(�`����fG{��J�M�{�\��$����C���(�5�D�F���P^+�d��5���ͭ�97@�/;f�.�Kr;!PD'�1��qy�Y�3v��=�\�c�$�Τ�O�����ny��<{�����M{���v�$�	&/����s�H���z5� QO=��H}�9��	'�8$��޽<��ξi�cy�?ћ8d���l輻�âU�DM�-;�[Sys�yW&;"�va&f��b"]Y�@a4��ܺ�Ӄ�8���x�i�[݃�Z{xvX���j��tY��ň���"l�C�d!�ю���u&V�&"�ʫIהz=닞�ZV�����4^KxQ�O�eZ*����1�<p���#V̑���v&Z�#I:I �)�d�ʒfd�M�I�l�Hq�k �#ۡb�i�d�,nn'a�Yô�����9�5��W��E���A6��.�Í��;Nj���x�,�&�A�p�H�u��0��O�y��zmM�& �;YQmBaN�J/5��1�4b�#H��Oˢ$B�Jw�s�wy:�{r��Rj�ZN��[�f�27�,����O�Sޕ$�I$�$�&�&��$�H��$�G/j��=�%�{��J��O*&p�I��ɷ'bN���Q	jD11%�UP�S��Y�݁g0@A��לD��W��I�VJ��b�����L�fcm�WAVu��wkM���O�3n����N�����zM�c+)�1 JXCn�"w'I��Q�}aʌ=�D�c��y��#JgQ��]�6���ɫ�<T�xC���\�at3aH����r�Ӹ�,�J��/�T:��8��LZ�e��ye3�d���ش���G
�!Ϋbg���������d�[cQÌ�W]u��R;��,;�bh��I�p�"e��Um"���d�;�(\�8y;3f�
e��7n�U�+B4��ƫ�:;
�9lwck�\��%���TzĥQ���Jtѽ�vΝ\-�o
V,��pv�`��8ͤ�s��$v���e�Cz��4��]�T^�C�|m�	hf�d���i����~ib�ȹL��P�e5��b�:�Łv�K���V�FV�I)�$�<pÛ�e5�u���<�@�
6(m's{�0)�ag�4e��Ձwt�b�b{hAU�"]I�Ԫ ҹgo)aw���Ev�m�nB�TdBt�[
���kl���*�Wɩ�)S�Vi���m��$�gH�a��W%4�n�i�y�ռ�r��#@e_hdĈ�Ō���9��	V����.�5��Q�5`�*(WZ��u�Mk��̦�:�
8xa�tL�L�&�@u�p՗`�t�s�a���F����f�B��*�2-�u�`�[R�Y�G��	u�����i�a�,r�M�n�.���g-������s�L��
�'c���nЫni���j�d.�kU�{����R���e�h�ʜ�zB=vjM]�c,�r�(�Pf���bwi��0��=5�Z���Ȍ�J>\�-sh��l�I��6,�̆uԜ�c�`�!���c&�HI*B�*�G�V�|�k��6Lm�l�oW:�v��;w�Д�Z�;��s�LyQ�p9xtH񙺹&֮�#E�����+.�MX����A2�u�����=٧n�Y�zb���8ڜ�ã7`"���˾kv��i�3	��TLX2��e�ԳOY��ɨ��f
f�fB;���.��s���WD��7��`�j��Ȳ��l�ܹ�U���.���:��h��m���pw��s������D=0�ْ�\�{uuu�V��k�5}j�
���X�ݵL�ea�U�
�/U�����[�8��mkZ�Ԯ?�F%OmЬ�DIwW9�,P]�<�&�`ڵ���)�rb��Z70C�_@��>�k��۲��Z�+�|gg@�v%ٹ��%I�\�Կ�U��� |{�����]unq�r����$�$�I��=�p@NP]�b�
Oew^�ԣ��Ut(��Ѧ�F�b�/�A�A"Z�[4ꪪS�Axdm
ƎU'xMwk�f��ܞP[#��v�xݮQ�q���v���]��*D��|�Ty�e�$]@�V�{��s�H��E���]`�JOh�.'��,�ԥ%�D���>�����c�]�t�����/���%AIfs��)ni�X����Z��*�c*��s,zZ����5z��y�d��dUMU
r�����4Ұ.�iP*��ka�"(��QQ\4 ��#MEb�DQETX,
f
����[uQUcl�L��Ћ)��Pԡe�QAm�&�h��	wWT���܆�U�p�>ksi{���n~��&d�m@~��4����� ~"�;��ӿ~L)_�n#K;����}�߳���ū'Gb�e����+��BVw3������!W�O�KLR�܈-���Y2X���|�@P���w���,�I3О�;�?�ׇ�xv�B��h��B���i�d*�����a�*B�)_�C����@k[�zt�ޝ�[�Գ`(��v��̴*`:�գ���o!G��Q�T��!�4#�Bw��)�:����t3�"�@��vH"�tߠ�9�o�٭�

�u�3G��}���6bZ�.��4q��.�Տ��r��]��6�o����L_wVu��2tӋ�xm��p)m*NgB'e�յ�Qo��ޚ�]��W��~�2�c[�7��r��+�2��{���Uխ0�zG��p9���]k�K�=�= ��I�a*͉���G��iz���hV�˕���nDWz���{x�F$.�V6�h�]@�g]�G�t��վiN%
�_J*r/}��/#�[u3��l>�����S8Х4����^]<+S>�$�Z�sz8��Cw`����E��{u��7�k�{���ִ�I���A��inG�)6�5R%z�p�3v%�?p{W"tS���Y"o%B��!4pӵ�=u��'3���J��?����]M���^�>Ԙ]�.+I�ӿe��}J5�l;pw�T�+e���[�4��N��<}H���ٱ����o~"�ຠ�8�D0�#g�cK^;��p[�0F�r�@�>V�,���,�|�i��
�Tt�Nauomhf�+��M��m��y�Ϲ��}�Zn��Z�9P�ɮ��㺂`���%[��̼���$�hsed��1����hA�;�[���Q�}�x{���T]&�Gˌ譻�-M�XXiJ�Gȭ�H�1ꭙ�[K�g��������U`�,����8xp���>�!�d�;d���`x�4�ˬ��M�=2t]L�������]vuyu�8�ӭԤ0̡�a�f��\^7����KL+��Jm�T[�:�}����[�[a�m-JJ6V�
A���!U��V�AY�lұN�
>�&H�Df����R�]����U�n�_5W�-�G/�)�	/�����Mb�s�
>���'�R��r`�Ψ����L9e9B�g���9�|�d@�d"����ǫ}SV��w*��}���[~���V1�N�<f�ZM�X��ra4�b�T-�,�I���b�����w���AB���q�.��9Y�ͳI��H��Bq�_T=�/]���Q��YT���e��YGX�ۄ�	��d�5Q8��9�u��݈�=�"���|��i�!dҟJ�D�RNE��S���ۯq�&��ƛ��4��'[�<�Y��3ޯ��z*�����Ħtͳ�����_p��
�#��������MuQ�L!�9��F����M�L���P}��#Ǫ_s�@��<Cس�h[1N/��x4��.˙�7���I���{�Z1OI�T�'�(���V�of:��3�j��)UB�S-4�y��6��/�Fyզ�i������n5G��s��"ێ�r��ٽ�r���%%4����mm���h�l�4c��b�-<���XC)��Ӈnz�HqG���zH���;�K7&E��~�V>�AL=5��+���ny쯼&�nt���K�r�\��ލi�q���Zi�����ުj��Q]�a�+yR��\�}��Ue�EչI�a1�9�='(�i�Y��ٛ��6��g�� ��ּ�*��sI�>�V����ys3�M��� ���7�fc��9 i�fn��!��8����"m��&�ΰ�Ń]�kLR��(��[S;JV^'�a
]��nc��,�n�� �Vj\f�T�wp��-�xA���b�W�2����ں�ݾ�{� n:O����Y
r��:��ϵu�w(K�6l�Z|z�37��f����ҳ��7�����˫������~5tnϫvh�![���yIP�@J�%cWs����g*��=�X�X³����AG��&4řܯ���gWZɲu��}1t���pZ��֐<��Ȉ�F2^��K�e��i��woP�V�oGL���Y���-�t���9�y;��3j.�W
d�$@^��{�ӱ��k�îo<Ƽ='e����D�Wr�`�o]kb�WJ�Ce]{�����!BS)�P��e�P�
�B�T�IL��uiB4e�$-(@Yl���[��H���U*E�������4��I(�  �R_	_��Rn�~势^�����IM��|w~�>��H��}(���/~��&�UIGTe)��eW��~.�� i�|���}�����7�8ͺN=�<��<f�����Jl�����W�X�xR����}R��oil���4!ˬ�[g�)�u1����ti�[��u���@Ӷ�3���ۇê���^�J>�Ly���'�Rbk�ǝS�Q�L3Ta����b�X����;�B��]�d�u�Rw��v��7�J�:��V%�M��	%X �}$WU=�S�W(�y�R�g��v�x��H/z���3��u�C��;���6�뮸(�P�jb��=6�����x�f��+��c�����uF]2�F]!�ّ
e�e�Tm/��e�u9gO��2؎��V�Si��|���ʞ3oI�	��F|�" Q1��(ڏY�)9�!�ɶm�%Pn������&j�u���[�H��b4p��fo&�B�w��i4Խ�����8��H�@"O�@g�w�)s3�*��U!�
������E�yY��]r��Q�3�sN�a��b�D�P0���F*�k�#Ѱϴ�:��I�dO�:Q��N]$�Q��\���9��>��5E
�*�����{�1�kTV�e�|lM2�.�<�|����|�gZ���c�
�7�&2��"O����i�H�d:�?Y��9D-ϐOT#I ����J~� �F]�|�'��MpZ�G�tzP�H�^�ǜ3}v�OB(�6��<�.Vu�kAQ��@�S 
��C1���z^�)�qzQ��%"�C��s�)�:v��j�b��*�<ֵ�m�B9y��,�Cy�k�)���<�W�le!�x�6��u'����[��^g�mwS�ktZg���1����&�
0֨����k��Uz�]��4�6�3<���k����z Fp��t�&}�U��/)�������y��,:��A0�>�� i#�u��g�鞈���+U)�SX�z�ۉ_M1@�c�E@��3�f��W~lӶE��N��εS�*���&<s�w��Y��g������Z����®�<d�	I�oX���h9���F��~Sʙx��k��˾T�6��3}׌<M�/7<���x�۷o����v�%&Ng,|| �O�d:�\�r@d���J�*Ŋ"�TX�Q�������Ӳ9���`�z�*z���g= A�D}ޏIE>[��S�>���+�b]L��wx�٪��2�2ٷ	����g���R�KǗ,C-D��c�_]��sU0�L+�:M��i�w��2�!��J�"�*��Y;v̦�6��޿�7̲0�聤A����w%Ս�uS��Vh��BE�ќ���]ܮQ����c�X��~bo���^����-p�B�}�Fv��*���6���B�j�l��7��m����:�8�WHg�Y }�+� ��~#N�#�>��~{��`V�UH��?*�������WD��L}��"�|�tW���V0WV$
��TW5���N\�i0�r���t���}�=y��2�.�ݹsTi%���y���66�M�_��N&.�$�w��Nu��T�
�X��L5@|�y�j��*�=���|��S<OZ���׬���mo�R���
Jc��O�tu�ڄ���%� 8�#HB:D�_b�����~���^Ȝ���,�I�]r��y��3�ǭեn�^��b�z�E"���S)�Q�m��ѮgU�kL4�Ψ-f�����x��q^'�D�G���D��5��/o��Dq���� H?�J��(��8\x���M�O�`44����l��鞝����;v��a���S����a��hz��e�^b��Y$��q���s9��ǈ[.��-t���ַ+�Ǐ� Y���{����Q��Z�G���I�������^r�g��:L�'L�}�=�g��T>��a��+\�W\���Ȟ�����fn��^�$�g���ƨ0�����v�0�q��;�[�M<�~�CnQ���>B�Y������S��64p�H��E����2��E9�k���g�
C��5��e�Wy�9�`��_u� �⑉�NYEs�Ve��O�Բ����!��@�>�����4c#ԣ̲�N~2C"��}��'��9{{f3A�Zw�ou�v����6D�"�H{ u�QڧP@�H ������#������7?q� Q���������UC#�j(�����P(�i;^g�n��ʩ�m�x��l�<�:s�g��(�<f.�+�a��u[7y�u��!�e(gǷ(�&d�YW��\��y�������3�t�ɂ�EZ�%u��[�Ŀ�s������Q��w��+]"
��#��L,����2�7l�M�Iw�R�u�O�.���W�5ɓ:�}��qv)�h�����5�ǖņ��]��*��^4u$�<T6R|�>�-�W͓K����d��)���j��n�\WAMهj�p�:��vG�1�v�W��͂t��fha@D���J+;���X��-voYJ���3ew]��}P��޾��
	`��{\��S���oBv�	BU�TIEj�d`W���|'�.��1�u	�=�s�#�������ұ��Z�Gk���x��ų�s�#�Q�H87�s��s�zO=���꼤�B��A[��d��]�R--�ZїK����-bDrʙq*�2�%D�SMԻ��(�**�b�*��b���m��)j�P))��h�]�YE��%(�*�h�۹���ۛ?��V.j�k�aWK���m�i=�m��˲��O�h�#�AН:A�k�u��Sn�)Ķx��O�D9ޡn�/�����륭e��r��Ol�*e:��]��։�ۄ�*c��r����OOI�+%�y.���0���Y�(<p��޼�9t� �T�AH) ��KH)�N��Y�Jd�)&Ф�Ȧ{Ǖz�9ƶæ�_mH(
) ���Xa�$������R
B�)�Ka�T���9�1|�Ì����- �:i�U�
IL8
AH(
)2�I
II����
AH(
)��o�:i�<�Zv�HJa��[Ő����ah���III��RAd����R�٧;���s�Q�|�x��o7ԇ��)��|��e���o�8�:볛�� ��
O��P�%$LU(�����Q�2Rx�L2S
H(% (��B�
AH,0���g�$� e)E�2m�����ȱa���!I�)��) �h�KH,4 ���Ĕ���R
SD�ytAH,��"R)�ƒ
Ao��l6�JH,������;ם��
a�
Aa��R
A@QM�RAH)�
H,0�Y풑H,�%$���V{��)�Hx�AH*�PR
Ad�jZAa��,) ����Xt�E$���Y�%$}�{�I���hR���
Ap����oL- �% (�L��
AdX��
H)<B���:�z�
)���Xi�b�$���x�I&���bSa���04��"�Ru}󷗩�Ă��I�l$S
���0�:�aH)�a���i����
AN S<��y[̚a�
{a�-0�I<��)�0�\e�$�H(
)h�Xt�[���r8�9�u�A�JH,�C���R6�I�����Y���R
AH-�) �B�ZAC�ZҙG��3�[�mZm@�G���b��Ll�wH���d�y�x➨�4�ݤNӶ�
AN0�,2
M�I �<i �
AH,0
AH) �o���O+��\��)8�0�����Ɯ�) ��6�R
Aa�;m ���R
AH) ����k�j
-���L��7�$0��I&I2��y�$��R
m(����a�b��+0�v���2�l,?}z�?���F��G���o�VCYg�y֏�W�(�G�)��_,k؅�l�\�p��{��o��s4[:�[��#�_:��S�M�FS��7Z�����rZ�pc��MAR5���/�x��}^�ل.�wf�6�-���Ci�2�Ov��k�)�M���0�U���Yr�/lZ"	��̗NE�Z������I�7kw�/~H���L�"ޔ|��|1=���vb�ST�̊u[LrG%R �r�;Z�c���q>��}@fot>u�]��������^��z�0qZ�a���В��lM����}+�ރ�/X����B�F>wlb����k�y�;�3���ݮ��,�����;�l?X@`��ڍ]�D���89d���x���W�Ԅ]Z���V_bm%�}X���}�*���di�`d0o(M���h��qq��Qk�O�����o����l@r��SJ�/ݷ1������8OW�e�:�.�Z��A=����ч]�Ǫ��=P俳���զ��T}���g��<����qq��U����Υ���a�I^�[m��G��B��4^Q�t���ʒB�d�؜� ����w?Y}S�Up+a���M��тg:{�2kh?G��ӓHSO۱����؂��-߮.��MQC{�'q�Ð�H�*p�s��lʍno��P�4L×~��3���>�BW3Q���.h[��xh�TvR�y��e=O�KT�WB~�u�Z����e˟���T���I⫴��}dns�y
V;�R��op^�]���G����h9$}�B,̥�ۭwog�L%Z�9����OS�||���/^��WMc��o�\�竇i�?<x��n�țz�R~�ΏӇ(!�A������oM�9h8geC�`�D�g<����U�C_�fAE<���0���U�:l���2a5�H�b]�J:'}ج�o��Irt�kC�e�=V ��p&T�SMb�G�U���ɭ(�y-;����W"k���y��~����ȸC��u̥	S��W;�a�b��l&刵ʽS:񤏬��c���ށ��ڔ�S�f�L�:`�$鷵g+K�|���x�=��Z�dTczYy�7��k���%���?��|�j#z��W��(��G>Y.�.U�r��|k�u�E�Y:��aׅY�����Wθd"}9�#"kAnՏ��6/V���;��TYl�+��Y(>Ŗ{�-�e�O[�vq�k^��
t��v��H��)��1�3,Jg��Ұx���bhe�8���f�)�he����1��it���v6`�`�1t(j;�f_�gM���Z��7 ~7w.�+s�������kQ����I����;Y�����!d�M�,�z�.���yYH"��w��Y����ݙ}�I�Ӽ�;���j��(�.�ծ���J��[௲�b����R8��Y��\C�m�� ��3�^��G&rue��]�r!����5^��H��x�JJ���uE����iUE�4�QDQ+Zֵ��j�7U�����2���UrJ�
n�4��ԥ�1JiQDE����DIHR,A-�DQ� ��|bu������!�6�MN<m�c�O���o��+�������OP�����}V���k���mRfo`2�Ē I�R�ïHE��^�wJ�ܣ3Q�'�,@=qܭ��==8{�����o79���տ/�� }Uk>�����ުSΪV�[_l�8E����7����0�ja3P��y����A#�i��߿����.M0���w����Z	(����H�-��@�����'S�,譺Oԣ��3�=;3h_��$���Y�_�� �=����'�[��'�l�:�v��p>�z�X}��^�������!q�Ν�A�KZ-����|O� s�J���쁋�L꬟���D�d�n[[�����f�P���铽���'����*�|��Z�)7;����C�%�����D��=���7�2�䒷"�i�<�{K1�OLk� ���5!Y���(����ܕ��V"��M[R&�cԖ�o���<>���O�*��,�f�O��$?E"�0MԻ�3�`eG���O����U��>�k'g)�\Ү/w��:�+�t����Kt�\5�g�����"��h��^����ly�xx���{4K����7d�X�oټ���̈z٧	hE*ղ�$�����$x{�~�DG��~�ܿ�P���FN'�O?��y�����($x��)�V����e��m�!=���?r�d__>�I���Rm�p���OH�w�P�vJ�s��y��/vnmAv�s�)�l�Б�i��]�/v�����6�4��x~ x���j�~=p��H�]�q?�L�?���ӆȼ��2Q�}Q�?�Cn{�xY�Rd���ő�VV�8���:�/"������)^�SX��܅�n�y�QuQ���J]s=7$lyk[k̺�Υ� ��qQf2[�%�[M~ �����{5�t�`Y�ﾸ����yM�AQ�&U�w�Q��[�X#�,V>����h�d2��:�^+M5��4��÷>�E�!=��� �~1]��L[��������՚_-�fQ�$�T퍵�ӡ�qե�
����fҖ �ŭ�� ~ x��<M�����X���GNu����w�O,�:���o��p��ʇB×�+��&h���U�5~������=^�H��9g��p=��}4����[{�w���Z8����/�Wz��rvx��lmn�����~> �����n��3�|����+�Mܨ��4˦�_U� �'P/��+zA����sִY��ǃ�8u�t/��%r7N�-r;���x����Sr	����?�����A�j�d�����R0K���n�t-*��|�j^�ͩ\�o�<?<O�� i�O�Q���D^���ȓ�3���/����\	R|'Nǚ��K�������(z<=u�UN��zrqoգO��ƶ���o����+��U�9�r՝�s�x	Z�r��;�=e-�u+��j�*��f-]�B.�9��4�-�d�a�CRk�D{p�`�p�9��/ݵ��7yJvՐ�V��%��y�o:����s�h	X[ M|�/�+���"����o9���;Z�;KY���+�)E"+5�tDԇ�^'B/��Ov�gW�ۨ]k����TG6��z^�=.2���&fM���9Zˑi/r�/{g)�j���&����'�>�F͋#��]r#j�iRq:3��w��O��Ų�ohmw�Nٹm��gg+|2F��I��U�I4z��B-��a���A��p���Ѱ�E����f�kj�sٳJ8�v�m��X2��[��|�3js�\��b"��g�}��eb���MU�Z�X�X����@ar$VA�9G*����RJ�]3$9Xl��U�Ur!%RC�΅epC����Di�i�**g�k���eo�}kx�rHu����Q��ԛP���{��{�'��,YN��cc��S�S�����E{F��V��V�غl��A}���(}j`Ɠ��r����z�2ru����вJ�;UK�r3yW{]{5B5��k���b��ob��g����DV@κչ��v�ΧF������%�e��i-�k[���������ͽ���>�����j=�wƅ,��J�NV�~�V���TEM|����RNE؄����c�a��ݢ/{[�<� �w�w��S��̒�u�T�57��P�)]]$���d*�yÙ�c����.+��q��q���Ò��*d˲�JT�O慎�=�}��w>��dO���'=(F���'���;^k�C�t�643/�>B�=��n���ٸ3�v*Y�@Q����י�+iޫu�.ζ�8��ز��5�����N�1�zV�D����]ª1̾�$��SNk�5�x��'������>�ݽۿ���ۺ)�}�ʅ�哀<��\#gU��яѮ���I�Qr'#����6s^�ḩh	~���.=�0ɮ}�Դ�L�ʓ{��q��NL�/}��7�a#�bWts���E/(����W1X�6��\ΰ�9ЍX�˔97�\����ā����?��~�Ζ��ߚ������?��nz�uH������x�ӻ�h��kz^�<�X~���y%�ا�����D��e��EȠp�Eu�+�jdjnص�,��`��s�Q�񬮝{N�:�h�΁J:��~��"2��A^ڎ��$ڄ�������x�xy��~�B5������#^�!��Ky�h��<]a�QM��z@e�c�Y[
ڭL2T�iTr}%{}���=-����3��jt��;�l���Y+W4��e�7\b�_麬Mu��2R�a[�a�B����/	�Pq�K�;}�� �<	����r
���=�������N�G�P0�<�]��v$�v�
�Y^ܹ-�����g��Z�_\mx�e�dDIه�C�T��'V�.�����`~)�wB��=���WE��s����ʮS���P闁�I��ى-��"-���kE����ߏ���o*�S�=������:X4�T7��x5��Xo�C}�m�#���9K����\��
;��tv��(��)��R�^�EZ����幸�]���s�
�_������ܺmeq����BZ���f	�wy�T��@�}�L0M��6dgcRmz=�` o�<��:�w�Rm2b��@����Z�K�~G}��xK����t� ��٢��rrPr�Wr���7�w�"�T7R��&�1De��t������X/3�S>��I2{���vK��r�7�$��ɀz�	X��W`��j��-���闰�j�&SoZ�m ��>���Op�Mѿ���/�m{D��}��qڄٹ��9�^BD��ӽC=��v�y��֬���ZGB�b��[����oמY��Z��i_e��6����D=�d��w�����늕[�+�@�6�a�'LL��qCru�.��K{�`3c���io���ݺ����z���o��|T'U�*���4�˵�N�S�:]��)��wVuv.c0��̚��e1�/Sc�"T�y���#كhRSf������T��B!:�UT9�͜T�Ӏ�^�6�n�[w���Vݱ*�0Q�+�]g�5�í�.$ƸBdV���p]PۭQ��ُxQ�[:�h�hl��+F�JB:��v�쥃1� V�0+bݱ��Ɂ0nT��C���Yn�-�V�)"!�bWyhi�&�F,,N.�)�b�3�G7"�.�_T�էvl[o��bt�)�p�1�m���V1�of������*�.Ґ����}gH��QTRUP��CMj��^�(mR��-DҸha��I%Yց��*P�*5)2�EK��&(�uh�S29V��-�����)%"�*+0�C��Ǆb @�{�����F;;�*xA�I4[I�����Ϻ�����F�z�R5ϟ"�:D���燙$zBo{5{�/�y����<�����ڒe4�bk�C��Bz2�̚��*�rk`�� �i���ΚWF�{���fwIp�k2�ÆR�p:m���CA$��O,K��m��9������}_}��/'�����~⹯�q�#G<X�V{���E��iw��|��$��_u�����O�{v�M��H����)}���#\��fD'�����GbN�GU�Ĳ�<������mw{�W�kG�ߓ�N���Ě�㒶����m�KV����߈�#��������S�B���9�,��;i�N�	5��ή؊�QU�.��0G-��⯷�U*v t��m4��q\z��A^������ˮ�^a���u�]�|�5b��P���E�-+,`��s�N���]չdQ�`IS<I	�*�Zڇ�����$�y�G%_��\����7�7a�?��A^���0��y�%q1��e�� գ~�����W�h�T�ӻ�k!��O׶�R�G��Dd�[����Ⱦ�?W�)j.��q�xG���Ԏ��A�<9�Qa��<����]?!ĸ�Kc���i�߉  3��M��ܩ�G��f}��b�D�{�ΓB�S�h��Q�����Z���Y.���DFp��y��A���)�j�����5�ӕ8���H���K:����.A���d����Tt�'���#�2�����+#6��#m-h���?�|<<5����Z�?\N:�d2,�j�����'�]��K��=�q�Ր#سpYgܥHcY�WL_z�*�7��z���cƴ��hs�Edly)س%�n��Ѭ��v+��k�8�F_���w�j�F�ڧ�ӰMK���jn�O�������v��4�s:�;?j0�su�Ƹb}��"`���b��R�ЕO%W�og�k�������Et�]}4��R�u(�5鞘،��ј�]��-��o�mn�7v!c�{�ϩu9Zǫ'<܍��c8��n����o�+:�ڭZ�M� ~>�'����TWG~�G�wB��{��1Мy��؍	7�����[��)9#^ݪ�j�Ȭ��R�/RiC��n��)Z��1����z,�x��J��s���{�0���ND	�O8hҞ�.�3�*���
�3v��?d��P��� ?��'� �n-������:1�j�~;P�9U�vT@1�"r�^��!�l�P���5jc���G,n	k<o�_������ٯ/�[.�Gڮ��4S�q�^���О�O��!��S�܎��]�}���e��\���a�P�2P���4d��?<O� �O?�����r����nP$ێ�ܷL�b��xW:�J�Yn��g�ٞ'*�:��"l̮���:����!��!�r��l�v�n�:}ާ�d���!�	��髹}��Ã�+�V=7��
�>�r���rn� �^{�fF��'{�V^�4��ÏU�vE ��ג���9�=���f������6`���I�#g˘�l��e:
�%�f ��}�� �[z4Q[��j�C5R������n1�tu}�:����F��ş�2%ko�VH�g�4^Jƃ��a������*-��P֦gN�2; iVo
��d�*k��s�=g�����w��If�4��GfA�8y��� �k�u-&��������p�P�7��p�m���3�
M�}2e�R�}�e�0�1�v!_Iׯ���l�ԋ�<�}Satܺ��b�i	�.ßmd���s�9��j���nجV���� �H��R�J�V�9��K���UU���J��TZ*��kS"�*:��R*V���� �R2T�Q:��j��auDҕCT2YRkJ�9�#�hJJ��+B"4-E�Υe�j��t)D+�mVi�H"��uftq�52����U�2u˃��n��'�#� 4ޫt�?�qE4��w�݃aV{N]'�b?�nr��b������v3��WY��9�6C#��[����΋>
�Ņ��Α�)Vt�Z�Z\~�^�^5£4��v��ҵs3/U�0zQ{Q���b�����\7b<i=�m�?	 {�����y~��ً[Uu��Cލ�į^��J.�R������-�֊�&����v��/y9u�������n�pEGluʮn���!?�]����<��L�gU�+��
h��b����F�ۣׯ9�3I�B��\����M�� \���}53[߲�Nm�Wu�M���q׮�lL:Y]Pst0^�S��^iQ�E�=���W�����Qb�jo�*��R}_`���&#㎄�"o.�ۂ+Ii�wxמ=8��1��Ay�׋ۺ�Sr��w����$�wx��~N��Q��U4�D �|u7#�����M>쇓_���¥o�J?o4�I�0���i���\{���#s|��|Ǽd6�.�q�s���������%s����5k�%����-��.ύS���յAE_�F����ʽi֣�vz���;�@a�,6�-����x��fWIol@�y�)?S����|a�i����Re�Ӑy��W����ݻ~K��|�'Vs�z�>���5�ol��Aܚ��<��O�����3�������ϭS	�s��6���ab�fQ��r�d��ZhA�2N���f8v��]Z7��h�G���eYa�*I�9�)KM��~x�8����?������>�u,�神7�K�7;��uN�Y�d���ܙ6��T/5���m����Y�v�`3�G,y�����h��'����-����t<��#�ͼ� b�&]Sڲ���;غ��,7;3�-LPM��6dgc�TQ�L����l�7���7rO�>t��?z�Rn��#�O�7"y�ֶ���W]3���������]���:.T�?��+˪
ј�r}���T���xfP��g��6��+l\*��9`[�Vt���upV^��mu.����9 �vD�Kގ4�jo�]��f�@�4I����e\�9�=a懻�`!x��X�3�fH�������<4^�;�Y�����!��ݼ}"��y�B%�nބ��/�N%�#
���Y�7��܇0ż�'�b1�ߜd���g
�+��Sh�=}�d1�����7M����A���_���Qz2�T=��+J���L��OF�:J����V�ɑA��otVq��[�p) R��c}��y� D�;����L�o�������r��Ö��כ2�̠G���d#�y坳��%u�oQ�x/,�!����
'2b�\w��#m·���]�ߠ���ZuG���TC�cM����&���j B{���Wda=[���ț:��!��v�9.��j[�f�d��R�C��1]D�֎��7o��UꖧfOG)�������[�oUn_!��-{S�N�����=m�/��̏H�=Y�\�j���X����V�� ��%��-���;)v7t+s�2ъ���o#ڵj죄�^@�&�0Q�����I���]��  �/;�Ԙ2��u�����i���iCz�.���at�O=|�5�������c�7(��y%A�;ȋѺK��i;b,���Ҳ��Sj�:�yqR�ZbN'��%���1/�k7�kJ�%���ɔu��#�f���*��&�Pv>➰��R.��|+�$��{Dp�m�a�s!,��e<��bs��$�r�̉�M��b�Ve���M.mm�IM�;Q�Eխ*^�)����Cx�N�b���{��J�*�kh�镨:�Ii�&����7��ES)b�,UA��q��Q�Thj�J(i�*��ֵ�tU5J�(i*�R�
��4�����jh�hEi�!I�4�#A*�3�TAVWS5!T�#DB�:F��5R�U,�EF�iJ�4"�j�(�TJRڴ��9�M�/^KN�:�!��$�4��Wmι��6����8��T����2g�FHQ<V����7*\��L1&������K���=����O�{���5�u�_J;6���#.�J�2��T���!s씻xe`G6�5BJ�.(9�/)t`\a�)M����N���[�j����H�ȡ}yU�r��\��~�o{#9�%N��5yy��l8����;�qvM��V_�u.�O���֦�*�sX�&PKv�%9��2rdU����L��G@P�dr���G�j6]w\0�q�5�S� ���\5U����&�S-��q5R:�P�V�G���⏮ό��38�U�>ux/��ᗷ,vk#����+*�޸��(m	3��;�ܭ&�Q���G;n��?y��u-{��
���a;ԯi�|+�y�<��l�Wp+w�{�U�B���FU��U0]${.�mGr9HR�����^�5�ڳ�A����JV&jZ g&9Sû�c{TePʰQ��g�3��Ƚ��Q@ѫ��E.\�u�y"�b	4ޜ��ď���S��c���K���������YSv���	�����]����jG�(��k�Rg2{�����4���uEuv�iW+��wf󽬨��Z�uO��?��Z~�z���eʎ������Ü�Gm6�8-��wu��mu�z��Ó��+�I��7s{���9߶�V ����{
��S3�,��
� ����[4�!m�Z�X�������_�=)�;����nmr:�%�ٹ�\3�O<d/��˳��8�-��k�؂�Ҽ/]�r�P���_v-�A��7����KLZ宓��1�����<���{B�>���"���F%p#w������ok	ׇbHr�2���x�A'{��יnv5�������3��Ww�Nc�U��4_6���w�R���s��u��޵�]�J�
;r{rb���v|_�ٙ���S��q&�9�R�8��LMY��%���*DF����y�ʼW�fbv->�����[�m0�.�їrP��|�M=ڬt�u=`�aKU�֋\)Zc?�?PYw�2�>�?�E�Y��7��ǩk�jl�{��/��|�����^��K�-�`os�"Q��c@B�.���Jie�w4�%FAY����Y���ї��e��Be�|��粲�-Gr
X���=%n���L۱��"�;�ڢR�c>����wi�#v�c�:��VT���q�4�b�Gnwo}{��^��g�4�N�4��ź�Cթnn�W��e��5��X�O*����w�(J�#MČ���hHVOmt`Ne:���\@�1^�5����qILRP`*�dm��������2������޿�>g.�cٻ��d���*ζ�X��j��.н�9ɹ^o���E�$����g|�p=�VO�@R����j����gF�ʅ[4Ȋ�a#H(KJ
2���\��Z�&�k�"��p�.���"C����]�6��EUྻ��]l�+D=	�
z�Pk��zE��g	& �g��Iε�_ˊ����+ygAt{��ܚ]�i������>���+�Lk��-�+��uw�����Z����O1�n�'�F�۝sU�}bp��\��2�:�]en�/!��o����'s]���:'_l��ئ���/�ᱤ�
��h\ؕ�-[j]�9�vP8ZzS�pnXB�BbQ&5	m�7cT���6$�K�Yr �0�%s�p�ނwWkK(��ȸ�u�v��`C�����+ẍZ4ne�pJ�մA���p�Y���q���Yb�,�"Sf����fj4�T�U@�SCTj��kZѡM	EUR��4�B�T*�RH�"i&�b����hEq$-ZsM"�+�QE��֢aXd����+�ш1&� ?�����v�cSk���K���+�9%�������B���(�9�Y,$�=}}��zчw*5��|yF�R�D���~��ƛ�:�ݑ<Su�L�d�}-�NR�{o<��Mdt�9Hpw�f3vj�޻��(T�������nơK|$�^\&�|���^]�q�H/T�%����܏Rj+Sq?�Yn�G7�����X��~İ<վ	٬e]�W�"�@�Ef7C�钊�����tU�=��.
�NP�k=�>��V�a��vߋ�b��7���w���܎�-#�^?/�~���-�L�߇�AEح3����tõ�E:��y��.#(I��@�[�)Do����{�eh�v�]�{��`�YC��}5c��l�����f��4��{�ݫ8z��?��?��R*�:ߌTt�An�D~�9�S�^�8��G��7��@׏��7R�-g���+�lO�;��^�{x	���P����q:�VXiJ�(�Z7���읓.���fu�Ev��1Y��؂{�~y��������H��'�]U�zu�|CQ/b��Y�����&k���C��Ne�d��V��G�z�������tZ��kG�og(��u�Z�pU	�қI9��徙X�����,��r�79wK;�ZLܬ��g��5�{V�xl�)�YR����y)��0��ҨV
Q���kP�t�MQ��R
��ڎ"��v�J��W�m�R��$ٷvk+��M����t��p�G���pf��3�yؒb6��[6��BWdK&Y��x�r"�yk��k:D�ÛY�@vY-��{���(�{ff�θ���8&(������O����M���N|YG/g��rf�)�����w��$��#���>��:���E�ⲻe��	TM�����.VH ���"܎��ի�Y�j��wܞc��qU��[>�o�N"I��o�o���>𠗜͸�#����v���w�Dk�}����G����U��>����9����%n6��>��=�{X7,��	%__.��B�_+ی?�;/:P&�E��å�.;��Y�6��H<��7��e�IsV�G��o{�Օ�u��O-�S���|�y�Qng�6�;��{�w�Rv�hT��]�;��O���
��6>��Ls��=G:���)h�~��yh�*�f�e^�Q�6!1�:�x=}�|��s��#"��^Gw�����ԯ�"�]��?}�[��b2I��x���ϵG�l�ֿ�M+=7{?'r������#������|3�D��r��[Sk-K�����3+:����d@KpL9mua��v���	��j.�����6�N)^s�.��]��#t�ڸ`{Xn(�C$e��C�w���-�Mn���][\�@�2H'��~�����_�L�ʕ���;ݯ�"c}�q��q�25;����/ݓO�{;^x�E2ѥ�i���>coa�R��q6�+��۰������?�=�HMk*��=Q�52�,��@�@ �ٵd�`��k�)`�27��+.T0���هv���%-!z�}����N��庺N�V�Z�]���`x:
�4&��%Jy�θ�M�Z�o��~YB�byN	36��aZ��N�z���8t"%�����(���*��$7��
MbҡyEL�HUf;��LLp�����!�[���Q�#U��SP�c<����ѽZ�J���ypTm�;h�fLw�pd#ՙ,f��؎4��**AW�hn��d���Y�-i͵x���)�7R˸5� ����͘hkWK�A����ٓx)n>�Z��얲��JQ��B��2�z�h�+������ߍt��������ij������R��Zi
*��V��h5�F*�,2�T��51RC#1%E��J�*�%�T�uw*���U*�$���Y�I7�T����(`FD�bP����m����TURP�TAQUj���~��<Q���\�DT�&~�W��`Su�^�?J'�:�\ձQy�n�����vh����|�v�t*���V"��/
&���6l9gUK�p�-�k�d�x�VXjk�Ú:�2}��{���r#şC�.;��m��~����KG3*�ɽ��]a:�J�-Z%e�ڎ�n"�	�/kn��ow�J�B�s�"���r���;���ʮr�C�A5׶o/rD�%�[��=�U�,�L�S|s���9bE�/x�^�~6�`פ�d�~]��츟{����g%��?<������^1]:6�7okV�[z��\s,K��m�"�4�wn����]�)�y�.�n��e��j��A.)��n�E^}g�׀s��ʿ��w���j'�жy��v���V�^g��^��~^�oZ��m��󪊗r��+�.8䞞�z���F�Ճp�G�	�Qy+m\-��J�u��5ҹ�]��k���v��y#,9��yy�uÝl7��N���2V�/lEl��Z��P��Jf��2��|�k�0�!��vK���c�oy[��=�MþO�m�}�{.9�ϠB�e>?�뾵�/RJ�?��ؚd�K�n��K�)s*�jG�7=��;L_������H&�pS�:�=~-Al��ݾpZI	��w�0v�=�+�7 �'7�]�n�.\�׃g%#��UmnZ�`^V���ڙ�f�\���Ѡ3���+�r�N�VD���
�6����8���K����H�0˹(�ͨ�q���W�r� W���͚������2av:��ol-y�>�ٵ8;Qz!���n
�|�{#���I/������Y_:�>J�WЦ.0�gf~���)�Y������r�!i�o�7��Z}u����R�d�@n�����ҡ����Yi�����m�|���UaP5�o��S�+X"ҿ�R�^�H����|1,9�-��9l�����n�J2�����u�'�b�s��G\mTBo̥k�r�����(	�]�J"B����M�LjO�����6(]g���wYR��������9$�ֹb�8�Z��m��ؠ�?�_m۶�y��O�q]lp��3��:�#�'1��G�b�Kw%��W�ǲ�g<�"�鎼�Y~Y!|�j���q�7g��.����T�ڭ�x6E����w^�l��Ҥk���W�����gr1�{o-|,�����f^�ɩ\������c�a���'�Y���=Zq{���&���0o�q��}El��R`]��[3�ه�y�⑊�j�������Mо�&�ݮ^F��짯�f�x��;�0wr^�0~z�%}��,֙�.���󧻪��#�*%����I�	�{�����C��f(�gX@��%t�F�ҝs5i�{���_
��܏�����N���ig��ۿ��/[��c"�����+��]Ć�� ���%��n�#�u&l�8�]^5_���I���	��AD��
iUQp��0��cm�$y�1��|>S�� O@�C�F4��f� �j�g��=��F�0�����V	���z	c��T
(�*���Q���*���U�L610%��d9�$		�������m��vR(((�0PQEX��(0�((�PQH����((
�͗%�Z표H��aR���0jRײ�ϔID�*J��t��?! �E��E=��#�^ߦ��k۫߁�Hy��A_��2d?l|	����(:0C�����CFl.Q��M��H�Ͳ'�T�a����{6!�`��O�!��~~���}@=���$�Ow��;�|�$I�Pd�!�@m��l)�ۀx�w�O����,�?����>��3'��S��t�Y=�G��� �F�$�. ��u����a��$D@��h&���!`�n!c ��J_���2�0�l��?����	��8�6hawу�|��}���`�u���ۇ��R�W���'�蠄H��*yhh��Q�IO�cb`��>�2� @�_��$�.I-�C��Ш�I+D�r�!�Q�B�*�?qG�0b�?,���O�d�5� n��aCt�؄ؓb�4dA,��~����ٙ��O`Oq��C*ї_��:D���V��"A�4y'� '�R�z0��`?_��ʺ��C_��%�aDIAI���@3��{�W�	�4|H(N��z��`ဣ�OP׾�'��r$?�}eO��>�A� ��9'�L��eFO��<�N�~A�=��6}�������s 6����w����ӥ�2�xzd��O�	@x|�p<!@�-���8�m�A �`m��?PA�@���O�Qh���0�(C��CT{:
���@O�F�fB�p7��aX0Bz�V{�!�a�;��H@�IDL�&I�=����l@`�{���46"RJ	���	��A4�́x�>���EBw79r �NQ�:4@!$�(�_������d	��� I"`���z�6�u��Ɍw�w >�y���q�=~��d�A= ����������C�>��$����>�B�>G��}G�?t<>ԇ�C�T�c�.z�?���>Н��G� �n���s���9�q 6|& �!����>�ID�V ����#�?���;�~!�A�;@v�s�$��C��o@ql�˃��1b$����?�غ�|�2����OjĆÇ�!��A���b�|�c���?��P�<5�g�_�=NN �D��O�P�i=ag�#�=Pd=j|L�6!�l(Opv�~읧�$���2}&�=�FH`����[��%��{�D�@$���?Ys����u�	��"}���}#��$�	'�O�}@{��D�{D�~�&�9���?�R�k��Y�]�C� ��
	�Ac� �p n��v��c�nSNb�H�
����