BZh91AY&SYc��hָ_�`q���#� ?���b?^ � ���
��V�Umf��m�D�%��@&ƩP���ԶZ[l�h�[6ĩ@͚��T��Tж[a���Ͷ���`R���TӰ�N�a�l�
э�U2meP�M��5l�l,�L�2�Z�cfjSd�i�eI�mf��m5���b�k5j٦ֶ�R�kb�M2�2 ��3����[mj����Q��4��hK+%���l�����V�f�1�JF��)�K4�V�D�#X2�[K6%���iem%T��LV�5��7}��B^�m4O�  l�ް
:ꎶ5]���t�U��N�ڬ���Y�:t*���J� �Uv��t��j��l�k�+����KJ�K5�[j�V�H   �� h�ƀ ���  f@�v��wQ�( c������4t.��  �v� �n�+���+M�f�aZ��Y�  ��  ;��   ۓ�t wZp� �@ �s� ��p� X�  in�(  'q� �ht��֓m�fke�kl6�׀  ��|  y�  1�pt �(� f,: h�8m��: ��N�����P �k� :�.���-Z��E��l�%�  <A@^��l  6��P t��p�(1θA�q�p 
4� ��� �8 ��F �p���-Z��m�m[(El׀  ��@�9  n�  �nkp@�0 ��ˀ4v���  ���à ut�]��\ �ԳIFٚ5dU��[f��   �����g  ��Q�  v���-:p  6]� h���SZ��6p;�k��@��+� ���VcmEE�l��j�mdx    р���p ������θ� 	݇ 
V�i��j�gQ@]��.(���P��[Z��lX[m�m�[d�x   ���mڝ��e3Z �iʠ۶n ݶpZ�� ���  f]p (�˨ WL��LI�ƫ����   1� {\ �B�@7\
 .�� 
9� ���t4t9X
 ��ۅ +t��J
|� 
 �{A3*���bd� �`�d�S�h�)ET4 41  @���%*�  h    S��T�P      ���i12�)���=O��Q�42��j	2���J(� �A�@#|���³�8�iZi�s�Z�[KV��v�:L�]0�V�3�*WLa����S�**+n����PTܢ*��q"�*+��Xz�S�~ǜ�}ǿ�C �!��
�����I'C TTW�G��@�EATW/�u�����@=$A{�*�" w�P;Ȫ" �H��"B"�Ȫ �\�!rȠ"�\��r"�6И��@�!�?B��v\�	r*%Ƞ7"�܈�d� B��1 �\�	r"Ȩ7"�APS"�8�@Ā��*� 
r(*7 �r�7"r 
�  r 7"��r"b ܈���)r �Ȫ܂!r(Ȫ܀�r �� � X�Ȫ �	���e�c�O�`ҿ+���+��G�QF[432��Ւ��zচ���flEյ1�V�GX%
�onF^��u�Qz��Lx��Z�X�0���{�ҦE7�*$�bIbʳ����)�s4����-%�1^8�j&��[ǉJ˷)m@r���j�^�i4)h��i�*VL�॥B��m۱I�ޱh^'R�ω�U!������һf�$�Ml�U�����s*��G	��(�&^�w��e�˽��ۏHv�1��R���N^�$y�ݪ�����cX�Vim�]1�S%���VӶ��Hm�d`m!xn�J��׿�Yt�;��4b���-�dYN�R�׺��ܣ���$�D� k+ZXX���?�����xۣ2e�,�4itA�Z�˘1��	7lF�9�JI���ͧ������Z�R��֗*3r��A���\r��Xl�I9lӬ�p�C�;w�W{K������c6� �K#*,�b�G�2
�����ݹ��lZa�;��%<!��᠝��H������Hʈڭ���qJ��chjHC�[���� �btb|���WGqҭSݫan�e\åգRT=\a�p�m�Vs���cJ�cn½��j�u
�����w��xt��&v6aˊ��Q��C5gAEZ� 	*+�ǲ�
'ok^ㆱ��$j�E�W3/F'j�7��g�f5V%U�VV���XiʋBʶ-n��$z(�v� Q���h.��G����Kj�Ɛ�*%������8zN
�7-ѹD�j�nT��&�i�	���y����n��U���� 0q��F�q�:�gUCu����p���Sȩ^b˷���[b�S X�m1r��oC���ң#.�]�v��%P�43�x�5��F���*P�mԠ�6����v�^<�U6�
���ha��G2c>�V�4�hI21���ۻ�I��b�ܒ�R�G1L��O^���X���]�ݼ�`�+�h��5d�uyj!�i�V��v��C����J�]n�}���K����!J"��a7��Tk��iHemi�<��Տz��=��I>�6�5�k��H�����10c��h��m�)DF�m��k�>�x�N1pJR�Ks�U[1�ii��T��zs�FU�j�ݬG)E0*P�FT�n�]���c�4�n:x6�T�`��6S��%,�U�:К^]�˭�4;���s;�PL�"��s10�x�����u��V]C2�j��ɭ�,��mJ�(Ć]�v'0R��V�նjd�Uc�����w�K%��-�0��J�JR���ݝ����m^��jwe�OKT�W	qh5lv x�6%6�Y{�����S�;gF�sZL,BƼxʽc���A����cN^�I/I�V�ߒF�R!Y3u@V��^��{��ւ�̴m���ݗ������+�y��y��f��(Ҧ���CLM�H�k7f]㌪M�RF2�fŤ7.��Ƶ����
���-�Ђ�I-M��j�%�&�dҥQ:Vc��,��E�\�{�7�����fc�.K��n��j`����XF��2�8^l�����B�4X4���TS�J�)��xEYnۻ?,ڴZzU��ʚ3]�y
�'v�D;[cr�+pnV23����� �� �Y��݄�+n�`QE��t2RV �Z�^���]j�H��y����@"���h���2�e����kӅ�4��>��:��9�IѸ�V��z������a����3�,��դ��l޻�K�(wM&ܥ�PCU�A�7Z�! eG�s"���̧Q*b=Ûѫ�k`J1�8��=�|�z�]���ϧ�TG����[5�B��bIi�N����_��
�� FB����Շ(AOv��{�QX�CEx��G+��KԬ�6��>��(,Z�e0��%m(ޝ�yՙ6�j+(c�� 횼c /���F�;�^h� j�S�g6���
��Ɲ.P�jvBr�$� n�B»�;|v8�Y$T���n�w�^n����,�YԗOOv��L��:����4H�d�fa�zsEm^GX)
�7h�*�y���6�7�)Y�Ė���W�f�N;P�]��{!dd8�X7���X
7V��]3F��Juik�����A��WeA�e]M��w(Z�`U���+I%�x�9��)&��X�^�v��ȶ2��aaP�wPUL*��F)FS�n�A�#!�!H��w�؞��TV�f�.��q�x�㶳�����Ҭ�������r�@h��A����x���ӽK5��&�2qZ��P��ҵm���InZ�eJ�s3Iʽ��dN�z�����,�0�-�n�6�J�*t�T�b R�J���-%�\5a�׬�Ԇ�T��W�q�	��������6It��C^�xC(�[�o�q]m-֋�4�4���sekZrP�V%�]�vʤ��"ձ7*���Cq
1'e�*�
�[���pi�õ�*��;Yk\����20��#��v�j,"Q���U�9l����b.��a�G)�ݖ���q��^:#���X��V�V2���t2s��6n ����̄�j�Ճ%��r�e��w[+`u��Fwf��B�p3ZH�<��MB���j��c�x�`����m�$��[pA����oq�U}dmاO�Q�[���YX6��L ��o#��Ezm��֤�]my����Ln%�Β��3b���,)���a�Y`lS\�wM¢�5�[ķ���0sq�� g��%bՓ�A��ʛڈ_G�CV<eh
�(	����g��J8�&ǘl�i�:���e��Q�gj��f����YoR���a�-8jͽǣkJE'
ɔF�TV���M�xY%����G�{J�fT��ь�ֳ�����hh�*�n��+fF�eL���s�p�\�qH�eTOd�Y�� ];ʲO­�%��/e7EeǏ'��U��@�v��ƒ��(b�C]�Y۵����$���-9��Qoh���L�����jda3ig�).J�1�Vs�[xA��%�x���z6��&�����p*��F��o��*8U۬Շ{j��uov��+��r��V�ͦ�ST� ��v-7B���.���H �g"��4�=T�6�y���&��b�bm��
�a���;ĵ%�	V��O7d����c̣�{z�8kF�U����)����Hq�P%F�n���,LA]f,�-�Ev�`�ٯ��M՚�*�O.���>�㻻�H�.�m�������*�@��5g�	"��IƲJI�gvT�0�,eA�kul��Ea"M�2}���J[�^�p+t�E|>E��5�M,��:>[1]Ղf���a��c1�0pҘM��7uY��sO�b����B�Ĳ�]f��
��K3s%<9G���AV�� u��D�j��P�����Eђ�R���v|�U4�k@�.-�Yl�,@Ҥ�![��b���Ǩ*��Dd�cN��]�2�Z�T��im�^mc��u��5@�lJ^2,p�`�y��σ���ƒ̧�x$��mSKfU���-���ݦ�m^k��ФV�A�Tt�g�!?�sq�C\XTVd*cz퓬n+&��y���bθ�ͣ���0��uM��ؒ+/s�ڷ��4�Q�ݍ�'{�j�^�x����LU�"��ô�,E.Dv�Q�Hh5�C]����]�9�����vt��U�V��NZ����5�B�b�4�aZ�1�lH���7k"lV<�[��y0���JB�X��E�`0+6���6�M��:�(�tW^�g���C5=���i����U�c��4�C� Z���X�j5Ksj��=�"m")K��X�<ثj�09�y7Y��&��X��2@�=���Œ��u:��.�ƶ�2Al� jQ�i��@X�A��ֵ]��	�����T[�Z��q[qK;MGH�YCm���U
5�p�)�;B�x�g6�Ԯ�@ �!����訶���Cc��#�d9t�+����1V��1���/��Tߎ!��Z�m�`�-�?:�U��$d
�X�pԙ6��:%�S�H4�N�i���e��7\�[��Z*��e�(߈c�*˴�j&��s0A�����v��zn���f�kH��blݻ{�2�7SߑV̩�,�a���n�Ѩ5�x9�N�4�W%��m'���F�Ɛ<)5k���aZ���.(𴆄m]jǷ�eG
7�3�2]kGh�IAffS�L�VlT�[4��5�"���F�yWqE��l��#�TE`�I�٘�9٨��UG,a�Q�^hts��޸,+���V�j:f���l��������ne])F�I%XM�y�/����͘pG�/w7[Q�xja�by��
+nP6� �qc �i|�u԰��E��Z��*mi5���m�5��z�sN�<׳1A��S]w���au&��r���)�O����ަ��q��,h��uu�UK�7�m�egAt�]Z�bƍȎ0�f��������K��3o-�L�t�n�m��wm�~�F��ek̨�bZjµ�𼄸n�%�*�%,Ѣ0��q�����Ƭ��/w�G�$�?fm��[BEOr�4�fҬ�o[Y�h&;ݣ����uRۏ �c�f���L��_YV��v���]�H��u'k:�V�,��o[T�쫖��B�bQ94�{�����Ɩ�2�aJ1�K�%�Řv�D�l�ܧ&��ctQƊyR�(RЀņ"�^��a�$�O�溛#^i���t0�ҋM�w�V'�f%#�(�ق��ݜ8l�t�'c�wwuLx~vC �7I1nCg-\6�u28S�C��kÂv9d2�ȦYD�a������\wv����swj��W�2W1�PI}Ăxm+v�c����[��n7Gr��wV���i�mK��e1��]^8�0�o�ۺ%ʽaJ�c���:�5��k*^�)M�������@��D4:���:��5fmj�#�I.��m��C�M�X*�lJIĐ7X�t�m��P��E �"nY��m9�����Y�áQ�m�G7�0m-٧�B����ʼaP��^�R���ż��n;��h��#X���/�YY,ձb[� �N	M�̔ ȁ-ʎ@��_�t>��^I3,:�p���u��"c��f���q�R42��Yۡ�'4YA���u�i���YW`�֑uՅ��Fv��!��	X�.jpJ3A��B��X�0�hk�^��IV�,�\�@��Ӽ��o2���
�4������n�1m��AU����wb��n����t���K�0��&�rh�[{2����YYWJnC�XТ�'�jd�ʷ����Kp)Ֆ��P�Y02��Coc7A�<t)�)a��k��7jN�rvC^W��qU���MV����1�	�S	��ё�Wf��E�kf�0BN�a6^�db���V4^�
`XXL�Z�x+=�t�����^�j��.�1���z�e�u������j�\���c�QϲMd�8�c�[��5v[:^`is94��j��6Ry�e����pa�w	5>0+�AC]�cET�&ō��ۣ���	P]�Ս�.�/(�`�a��sY�6�*��I�,ܙy�6H'M�1V�����\2�P�cjS�7h�u�R:��S.R�h�t�l ���]�m����] χ ��j/4�R��V���*͍�8�+hJ�qn�Ωp��cN��E݊q2�9��F�GR���*Cb ��M#j���ј�G֘�L�G�-P�h�8/�����a�#bYYB����c���퇪�H�#�2ӗB�%��/������O\�W����s)Vyk��}��*��[�"������D4-���%2��LW�F����[(]���:�kF5��-Zm�)�0kP"�%`�{eL[v)��ɱ[NmYH!	�eK~&7rfS��Ѩn�AL�`lT���:Ԣn�n�APl��z��F]k9b�(:x��էb�7�Pjm%oB'K����g]!�,�i2��Y�3�B*ŃNM��>�_m�q����٥Z��aYV�И6���y�؞f7�A՗�yV��ԭ���K�B���^k�#pCY�V����P�m3[����c�wH#i�o@���ݍ�XK�����K�'uo׵H���H�l���!R��e�:�̄di 5f����$�������������)�*;���V!��5Ty6dÚu�B�ˑm�"�Ո����B�����a��Fa��`hD"�Al�x�F���"h�n�\�Zt!�Gn���K8F�yz��5�ŉ�#l��MI�n��ӗ�3X�D��C3y6��(�^^֬l3t���قI�,�I��Lx�eh��[�M���CV�̂��kh$�8&�RkwZ�2��4m��ͩn��0@��9�����e�R�vME&�e�t��Yl�1��.^	��#&�rX�D�㔝õ�H�&�VG�w�S����W��T̺��
@�/5:�
9EL��ق�ǫua�u�/PC2ӡ���յϓDͺe��X[��]
�X�,3����)��V���u�������l�`�SЮk�I�Y*4�jy�K��x(e(U��6T�{ViG(���U,d�]��IQ:.����l�Rٴ��@�h;@`7q�2d���m5�B�!YliٱP����Ѡ�̷O��o�k1Y>�L^#*�%��֝M�L��hQ˚m(S
YlU���"٤�,c5����iҾ�bVTy()�b�I�r���y���n�	������w�6��oZ/�6�E��饴Ry2�v�EKq�ف�0C��O�A�5R�g3���F�;3���ӭ���)��5�_]u�\3��;�E8�̼��9�l}�J���MXSg:)-��N��X�c�	P��q-�yM��;�m�����ܬ�m\D!WF�=�۸��}��']7:��0��R�L;��]��s�k�N���dn��Z�j0�´���z��'��}X0�����c��!�ι�n���pm�LN����N_M�E'���*iڐ63v��P��*뭡��'7M(k`�3n�#|2R{g-^��\�t9&��M���]��3��*��\+�L���].��k�Z�ɻ.�SCt��A�(u�M�'�d.n��r~���[��s]���ԝ�.�sYW��!ɴ�C����-ӑéNy8�Mh�i��y�k���`�쬕�WVJ5���l#5���u���̈��f���H+�I��R+!lWar�%����ְ�M�C�0ǯ�&2�u�u���3�r��Nu�f�Yl��)9�^g<��2j+:V���8%V:^�un$p��O_.�G�pU�U�:�'E���]Oc���=����I��W16-#eܳ��S�k`v�׃Wq���W��S�K+	�N�5"�g]D��FH�$�ܕ=PFE�_R���O6w�C��*�3��9G�]��գ��<z$6���,]m^�J�H=�����7�F]�g1�5Al���C�Y8��.�tT�pK��c���Λ7f=��7D_hϴ��!�A�p���5h�cUe�|�Y.`�o�X��X����N���}������ܲn]'	��8��p��m�E�&�i=��ⱽW�Ii߲� �8'l(VT�-����fNIk"��hܭ��ZW;�[���qr2�W �^Φ:f��nT���C�cH܅���5U���깯��=��Ma&V"��4��L�{V�wW�tv��R��$�9kt��l�{�h��@��gHlᤝk��!�p�nV+��m㵮��ۓ[���[C���TVv�t��QC�����R��Q�\�Lla�5�[�L��8W*�T��g�:���r͡.���=�uR��>?:k*mK$1�v;ene�1���oO��J�p���-ǃ{���u0ɣp��!m��tґ�3�B���2��㐫A7zn��ӛ�;ֻ6-��	��2����znŕaH�t���l��}�k�fP�̮�6V�x�y�}�\��xr��x�{��[SM���U�������5"5r5p���X�XE����ƨ�kE�b�e.fm= ]�o�K`J˝J�7m�t^��o��PN���^�|qy&n�y��B����#[�pA!VlM1�����A� ��S�����Ļ��<ސLu1-��|k�Ȧ�}z7%J��h󝹑��n��OC yws�e=�T��B|����L~��ԫ%��Y,wެZ�<��,�Y�{��1�@���X�s��23|i��W&3�wݸq��R�1�W����4�[l�6.1g��U�7,�n��M��}�7��ڵ�.��ޠz�F��QtE�Pw�1�Ƭ�XE^��Y�qb�&c�si�C��.G�6�FE�Kz�6����TZ�}�����eu�y��t���YNJc6���Ѣ~p�3:jQBw�4ں�bc��ި`��̚"����%Lg�1���w����@�r��[���Β�֌�끍��4I�4�j-[���o�R�����>�+9VG�Q!��T6re�V&�oc�����gAưP8w%1)��1GG�F=�G��w���N��xt�vFۆ�^nË��z� �Z�8V�.��� �٪�]}��o_^�6�)ʄ;4��V�׬f��t��>�ޖ0ك;';n���NjR�%�uE1-"f%ege�ʔ+j�ï��R����n�����ks��dr��� ����Ίm�ku2��Y��\i+�k��e�Z�^��s1m@�7V�qS�T���jX�k_q]*�LɎ �ڝYY��
��NN����Zص���X,�:6���w� � +.��z,��*��a&�=�Йn���Т:����W�gE/����%W�OzK톱�p�n��w,B�w^�l�x���L9���
�Mu�-i^�a�yj� �W8�5�Ab�ԧv� ��Z(��l�ԙ5eE橴����sT��R���]2�CZz��av�n� A��,�8�۾���x�m���%5����7t����w�+b�qme���tu}ܹ����Ab�J�m{�3_���e9q�a�B�<ͣ��ZБ���}C/-C�l����Q�i[]x�b,I�Zf
j�bC�)������]S$���}������o���Ǧ���قLy�z%1��znZ��u�05xY��ޣc�|4=�����^�`  L�7� ��lӀ�+9����B�B��ۛd^+	7L��nYژj:͛�鶸��C����х�nay��,T3(��@�	�JOv�S��'!��]f�I�Fӥ�	WՀ�N��\`���,��LSV��2�|�*�e&����0��g�%s�wR\��tT+)h�0�U��"�q`��P�[�X�.��`���{Ʊx&�v[��U�KI{�l��s�q�0Fd&�������Cj�Jܩ���@�J"�XO&�d���.�e� �֥�K���ǥ_[�j���`��`%�8�cW���+���4�.�`��X6��CO�u�@��"������Ș�7{f��`uG�ݭZ�wa��,�]��ۓ��Vp2V�x�Bd��4�e�W�]�_}�ȆS�'%��~0��J�J������lš����5�$�t*i�X�]�����wCs6�F(��|3���=�(U'��2�^(vR]������{��;�@G��B� ��I��WPU�@]���^t���f.<�
��cy:��1t�Od�����yzb퀥!2_k��r��b�q�(c�AW=W���i��:���Tf�c�t�*�������q�G+��o���{v����雷��db�İs�9�p�Ac��z��J�ݸ��S�w����Ѯ��YXn���~�Ox"85�h�����\��/��h0�EW�ҟ}�uMܡ��c8����=4h{�L��fF�t
캰�������YԻ�Z�m$N6gS¯�R�Kb^.�}��mr���7u�ژM��ʜ�(`�K��N��GR�9>���
 R� a�d �\�5�d�Jve;�z�;�m�Skh�=$�W�b��dF��u���p��;R��g�lL�����=�e@�v_95��L[6nH.��qj��fj����ՐpAu��
]��rдM���@��V��,9��Ո��Ԙ�����n;u�{Rt�ɐgL���`�x�3WQ%V	r5�U&^����z����r'͐��M�m��}�T�G4Z$a��:P��Tة��G]�f*��@�Jj�.�i�Y��qo�a ��h���@O��^{G\�6;�]th��r<���%vt�����IvWo��3p��8*��׮V���Ju�j�+5�tI�È���]�^��}>i�ÇXBѐ��nM\������ԁ��V6��f5��A*���-E���f-e�M`ӆ����x���#�(�M�f�eY15��]/&����z�
c>���@�\ղ�M<�M4B��6��D�[�|���Q��\k�EeA�U�Y�2[X��Ѽ{�R���WS�c�����A&I�?��)�4&q������FM�[�=4�71CC�U�n�r�V/�(]*B��ኮ�j�6�	H�6������<�~�x	3�ХL�י�t�u��3�qT��"�g��s�18eo��sIf�5���h�@!��ވ��p#V� c� 2�Mc�(A���=&fe���Q�\u��r�Wԕ��z�Xh�I	8�(�x�bqi�'�PWɡ@P�-��ǣ\ɲ������)����PcMR:�˕|M^J98,��}�̼Ē[O�fVJV�U�a��(f������甩h+�˶�ή�8����cC��7�ޣ�Ʋo������C@�+���\�����m�O��
+�N/6�i�c���**.p9���7Hp��L��ч�Ka�y��f�Ri-��en�{�K��f�r7���;Xh7��s��-�x�͔�;��\wY�s��m�;9�9��������esp	n������(R�=�C���l�u�:.���2�C\�V�n��-��s�����,��J����	D���2��	;(�s�}��s��ySn ���s��X6����N�6��0�Df�8qc����ɜ�'زC�@k���V��d|lν�����|+�,�yv���zI�#/�5$��t
�Ts��4f}zb[Z�r�H�3%�SLm�!J��9�~\��IɎ��$�べe�Z�.�/�w	o�,��0)@U���Oo �QC�=��u#U��-e��.���2��$���ݽ''l��L#~�X�<R۴�uv�w���z6��¹Љ�b��*�`^h`���/q�u`���:���Or>i!����)lh��-u��/2�*|JϬ[�nP�c��Un�����ٙjBUey���.� �o� ��5�i#��A.'�޹�ru�WX�:�ol����� �x�x�ut��֗�qF���[ڱ6�Ђ�k���bgw0�_A�M��uQ�jV���4��x0���b�w�E�p��ڇ�۸�W_C�֑���Y|tWP��[u�N�{5��Iwk���;���PI\�ܱ)ȥ��f�Z(v��6	�&�-[�f%�:/��)�mh�.��J��:�������.G�wȧ�C��o�X�NҨ�s3iY{oY��4�x4�W������S#�P:�R��s��kq3�o7��Pu�Qd�^p_h�4�/jҷ5V�9��!�zV�R��3�����"���ݵ�rݛ�]ύ�V�Z�[���-D6e�Kmn��Z%䭵A'B£ ��o�S�-tֲ����_5#S�j,5�.V�N����\����k��ǭ�zS�������Mn|w�F��g�,v�s�L�,�Ǖ
��9 �^��9�žz�ʴ#�h9�}u����WR�6+�(9��7�Ѝ��Q������V,���*,��ƀ��	Le^���j�	K'ee+J�Hn�][b�LG>tp�+H��Oxi����'��kt띓��t����k7��bμdG��"�Sm^���ʍ�;�F�ڹs.�ĭ�iL��Ps�ݵk�.�揺^m��[�TU3tM�@Y �J����M�Hj�nN��=8L���D8����X'G�;�]+]2��:���,�1�"�$�E��?9��S��#	�@a��U�;���lK��*0��Q4u�(�Ie�0�`p��B0"�@�}qh��2$i+��-R��~O+���ak�ȶ1�r�m�1�,�X"�9Vm�u����D��m�3*��dn�{6��Ʌ*�!6�wdR>�+;;Jsp�@�\�T���r�o� 0-�����ڎS� ��̝?ﺐev��[]-��4Il��,N�[�]b"��jf�nj�l�i|B�WC��#1�Ԥ�7��kBڍT��bal̋y�;"l䲮�|��I�yj�w�D�]n4�\g��S��$%�4�!���;��as��;GF�5�]y/��z�܌��$�%l�ꩵ��G^�e:�[-f!��Gd۩�4�T�Oa���m���W|p��e�-Lz���q�-��Q�0���c�ӵ���)yh�kQ�PdT�T��PM�JwG�\Q�tM�sw\z�v�o�n��4b����'3[ϵ��8��r�x���G(!h��iܱgV1֭�]Ք�;�P�K8H�r(ô�`b���]e4Lug/�a����龴�k��X����e�4����}q���-���h�B�[.9�U�j�1��*�t�f�F��5{�/�:j��sg�L�˭���`ʉR��p}5%Y�	r�__>Ǌ�H��a�B�ܜT���l�@4�Or���o[[�9p
�Ғ�����=��Z5�si;��t0�Eb�=C�ʴz���#RS ��p�pū�:=Pc;�Y�l@�;ou�:�C2ܥ��}R��� +lހ�`
�B�z��鎺��+��&�4�řVf��y{V�]�n��t���^6���[A*��D��ի^���a�u
�2b�6��v>��V�ó\6�ͣ�P�ݮ��Z0�V��Qo�2`b�ñv�����..yv���n�OEA!6�{���l"�6�9v��6x���`6�αЅ��7q��/T��ø�1�q�yJN��a���7��6�1�FU�X�zw�h �=���Kr�1�A�q]Z-�f�Z��5�g���!w�bR��+q�.�_7�Ů�Xw���Z:��cEp�����3T����\�[��܂إ墳���rQ�	���������:���K�-�dP�җ����L���� ,��Y'b��݁��>���c�ѣlSS�̕��4�s�F9�8����%ո ���XމnFL��mۥ�i�ҷ��J��x�h�O����h�C�}��ۚ"�le.8V�em����f)zl34���ΧT\�
PGy�\��kO+�d�k�h����3^+�:57���۔u˲���ri �*�������i�%u�7g)��%.��щ�;b���S1��qtM�U{�\��+S����\Le��hh�-�u锢���L��Je[�m���;7D�L=�P�ҋ�2�e�).����ԗ��1"a���+�p�Cbfܥۥ2��kMF��sV�2��Sr�EI�9b�{�����9��W�D}^�-*���p#��es_xV���������՗�Q����ПO�� i�&v��]O]]�k���p<��DW�������^�|��)�*s�������g-8�Ƌ���J��0Umu�·��]hL�ʂR�U����[]	��(�!�ܱî Ƃ�NA`}76̖�.Ok���.��C�e.�NM���Q��hԲ�1���	�v���L��׍i��@�.Ns9N2�#z��V��ɴ[WʺƗ�o��K4N31K�/�Qٟ^����.�x����^�
dUyۗS�-P��,t��]��m�PWFU�/s��ɕ����2@f5VR�:�,}��0r�vP�{�Td�������Y�{A����a�����ZQ�S.�u�^J��P�������k�>Ű��+n�u�u�^P`(�C}�ӊaT uܦeE��	��a̷Bz0etp�[�;I�2�����n�$'�܂՞q�N}���V��˺e��<\l�y(i��V�e��Nilt`9�q�Џ��u�\�چ�%�V���1�!�h��ʃ��ڵ�o8B7�Z0P��#CG'�wd�<��6�3��7�G���\o�{0�t�2ĥ@ǂ5Ɲ23�O~�� �\,��|��H'ū�z�M|�+��
�b$���	��+��laql��F
����i��w����1G���໙��Xkw����D�brZ�2'W�����ݗLԘ��'哕�v�v�h����t�ͧ���\����ܮw��Fg�o)����x_��R�TT����|pa,���Sz�
�����Wuڋ�D��lb�.�T�B+x,f=-�}�V���8���Q�vn��9L�ŐV�9�w]�	0F�֜�I�k/��S%��Dh
�tB�]��%a�g�]&�Nխ���&5EK�{Z�%wC���:eZw�Y��cLT��}M@e����Ff���4Mt���t�8�N��s��:}��hs ��{���	��rv�F�e�n���9�������G\���2ƖL��j�-M]��[w)��eV)M�'�F.�C蓩�*ea�Nk�%��a���|�<���l<`D5d�X9��nK���"�	��4��L��ڶP�DεMI1��y��Elߗ-(���T�ꭝ3��\�:�.d��_n��\�6&ԕz%�ޠ���� �(8�az�-y&Ҏ�y
[I��`�2�#`=|�ǭ�U�o��^�f�D�O��\Z�]1ç�dm/T��w�mo��_q�*�sTiv��,�)�^��nމɫ�dN1u*M�ѣϦ�S�=,''9�ҳ�'҈w�旚ބ6X�Jʛ�f�5dR��H���Л�.{a���Y�F�����ی��)[N.��������_:t-fg	�8��W.��'��AV�N��x�+�v��J��9�wz�]�N���Nh�wq�),�Ğ�\�eꡌK�Wuڳ��djי��my�ilк��y����:�W�i�[����ڪ��*q�l
�Z���{��jKg%:\Զ�+@-4�yՒfB�WK�Rոe��.���{h���Z� J���J��c�މ&e�\�D���s{PZ�7k'R2�VjZ�j�>Ǧ��J�	��ҠX����&n5\�N+	N��'�0o
SU�q�Ns������z����-}�-+�3VX�:��*��}/aȯl:�C�f)v��ۦ���2|�LI���^5�Z'XS���;G�)���ugy�M���m�b}�lu�wkn �>]wXn�s�V�
��m�9v�|�JX�P-"��cd�܉2��]�T��7�$�����$2c���|�_Y�ԸE����n��M�)8��a�;j�ʻ�68؈ d�1�ͧ%9�7k\s�^ox0âޭѺ�	����Z�o��B�}1���AF�p�t�飥�:k(��L^Q���k��hV�W;���X���1n�
�݉�>���%3R;H�uY�ݶ���/�Q���y�{Q!������������ ��������2�F�Z*l��֚�镂6�4+�Rt��K���hY� [����u��02���c)#���5�6T7�U�^q�O�5��=�Mr�ڒ��@���m�̸7�c���+Y�{��.���m��9P8F�Y@:��<�����F��u��9"�>����tv�1��۩#<#�^5��ݬ
���&j)��J�mbY�q�L9K�t��p���>"s\�om=��^�T�.Q@1]-�
������P����]��l�%]�8�7�ᗷ�� *�w�re�1�vѱJ��w��ۛ�\�wj����j��@8����a䙖+�p�6�)�lᗉ�6�ޝ@wr��vAv�t[XtB%.��#0U�CqmA��+@MSà�ܸ򛝺��Xϯ��EJm�;]E��Gs10.�:�K����֫P7�d)ի+���4]��nhԨ��a�:Or��zEjO!䁱D�,3CP��J�*{�s���O���j_^�ј�<17���"E(*N�D��X�:��w��هgP;�xP���䴺��+�vf@�h�=�c�K��ǯ��u5�B.ա�#E�跈3me� <ݥ���+����M&9���*��ĮI<Hs��͙N�j]K�Y�C��7&�����Qù�OGw�&�]��q����oiN��o�/�ww)�Z�sB� �KXX� �)tz���\l��Df���ۼ۲���f����)Ϯ�+L ��[��a�\�t�&B �x�|26��NϹ�q�)��r���:e��1��A�˼�c�i'(Kq
Fhela�WhKA*Lܮ������W`�xFzWW)&�L���e==O�����5�-��Z(qco����(�I��;ǫL��V6�zR4�(]���_l�#���\�0�v��E�����)���%B����V�yy�&��7t[�3�� �;A�:0�XF�s\lKP����p㣫y��3a�y%�$%Adk/]�{�vwD���F�VM��F�Û��o['�Ɛ.Xo�mQ�U�WNb�dޓ:�
<EZ�$��4-j�MӦ�穳���ݾU`4��6�Yc c��t����t�	��JL��V�3���uv�l�����v9nN�v+M,�e�y�vky���]�F�8cu����6��&nS NO�w.]o�]�R5��)!a���%V�	<���ջZ2ڱKS%H!�|���J.(�<yދԋ7u���y�<'�����*�Ʀ�eY|� �m{�l�&�=j2�#k��R�F��Z�ղxΡ@�f��ܩ� G�n����]3��O�@���t�A]�E�^��+zI��9T�,EѾ蒀֋w|{B�!-uj
еz:�q�bfB��}� `�*L�ON�[�h=t8�����;L�u
���7-U��buj[�8e^Q��Уm��q����khL��w�A�3kb��i*\+pW-&��$�\MQ��U��H��K~���\ҧM���[��8��#�ޝqHٟp
��U�.���P#�U��n�1���I��8��Um��DC`eYk���ĭ�-e��/l�0Q�M���T���ږA�y�p�)�����iv𼴵�σi[�v�+Q�9��4��80��c8���"�uV�%wB�0�@Yʶ�TiW*
�_;un� �P���Nf�E�.�����ܥ��\�'Wt�q@{;�-K�5�{%ػ5uiKv������*���JEu@g31�V�eIآsd0J�o1���I]KY��Lcwv��ZHJV)�U�I^v�a4��u{q��jR�E�*H�<ʏqZ�8���I۩]%�keѡ�t'�5���P8�1�V́���*�Lr��4D�p%Y��G�X�v�
���:.��ժ��M�T)ċ��ʾ��%ꍞ1��y�3���#��B�[�2�>M�Ub�:���XJ�Оޢ*>����]�f�li�g�E]4�n8�a:���;��О8�[�V>*13�v��t���!
�
�+fL��>G��GbFL��Q��IWQ���Xnۣ˚�-Y|]�C
��A��,m��ݍ�M��n�eK��x�]i��;��s�.�f���L�I��dG �ђjTy,��3A[��%�����%�h�f����Q�T|��Žpuj�i� ;�$�N��)�T�Yww�3n�0�����ڕ9 �P�����Z�	]P��pA7ZȴUJ��j����ǫ0iǽ�tB��D֩�Ce�GµPzc������� [ o+�i���v�u7��n�z���,��ŹT��-��U�`إlVԖY�����O7@�F��'&�D6�Ǖִ-rKd"5,
�����[`�Y�v�ҡXjo^Q�ONdH.5u�j�&T�a-��yv��8�J2���v����ltUȘ�u��(�|�R,���[�ս��ۇ�N�nw����0n��U�q�H1vt�s�Hh]��������g$u�]F��!�
HY��zZg�{._'Z�����"F�Uj�����(I+�T�}���ɇ;�h�1��j����'�$Es�N �Y��
�y�.Ą͢�y69�b�qh�4kq��Y�n>�u�|u4�uu�R�&;\�,��|soi�D�!��
���d� ��(�U�Θ�KV��n�� )t�'�@�n�PR�u�b+��`˾���T�_T��r��f�Gf��4"�(R�Ic`�2����c���ō[٘��.ѱ�m,"���`��Yٶ�I��������]�v+�c}�J��]��v���Fp����q�s�F2]��� �^��R�\Z�*�`H��b��Z��3(��i�	�)�`Z.C �"�Ҫ��_v��S�S�Ǳ
��K:�4E��0��+�MU|Ĝ�*�d%�BQ��{I�gnQvr�3;�����bj�F֨�4V��|�']%"䶆F�;^�(���..vD2R�*p������t#i��t%��<�����Ce-��7H.�ёcV�K��]Hwȋ�ЦmGN����'���$�Bi���&�Sr�1W֒n"@Mm�O#��d�O
�m}bLݭ�U��z�
���4�tZ0V�*������
��j]�F��t����z&�:냬X��U�w�î ����� i�C����b=;�;�xͺj��19��Er���uʑ�Ox��	�Fܝ��sCҧM4f���t�Y��NT�σLJ�A�mslb���)#��M�i�ɂ��έ�Z�����&�lˮ�\��ǥ��v��]�}��Jƅı�청��		*3h�Bč6�;�yI��]�E�46��-��F�l�M��tܶ8�1L�5��7�٧rc�WQ������c�Iw@�1�m��Ӓ�
��M)��i���QE��V�&ed9ۖw������ԝ־)���=�?�*T��� ��1�bgmm!ϵ�=�j<�G2V �w�H�A7+�:@�D"�ᷖq�N�`e��}��_<e�,�o�УGX�55h;�����>���ҡ�Z�����h�
�
TYl$eoU�7p���ٔ��'�)�N����NY�f�סPV��Ɛ�$WU�j��U/yR�N�ضS��˵e.�9��1�t�S�d[�v0a�oEM��
P��y�Y����� �u���n�
N|\Bd��q�C���6j��l
�t�j�m���/��� U'���c�+a�����VsKȠ]#��*oY�7ue�o:�%u3�6,6;{��ʒi�++;.�i,�e���죑2Ҥ��(���:��n��NY/LN�T\�-[OV��u�����qu�+1a�2�YqiJ���C��S�Zs�`�y��C,�P����wD���=�Y�[Z��_t��5Wfk	tH֢�Ƌm�v��V��N��j�`��$?����+g��δN�ԷuǨUūLY5A�U�G[��ܮ	��s�Ԟ`˫Y�L��X�ăNd��� )��3��A����7L��N�qC۬M�HV��&o={ut� �]ц*�[2;�k̬��=���v�nM�������3gy�ٝf�U����ˋ�KwkMF���+^���,���r�ꮆ��{i�*U��L.�vaDb�Ј.�6�����3q�eA1�*lM�C�ͥ��o2�L���Ԗá��3H�f:�U�b��\�	�o�ă���:��� ���N]o%6+3#�{z���pҹF�Q�����Ԇ���˙ư\/'PZ�c���.\Y,P�v�Z/��|����Lg�32��]�X���Xr�@�4ֱS^v���;���
9kx����.S����Xj�����#Gb����z�U�+���qX�O���樷sRߟa��]F$�͹j�ܵ���^�k����@%�����ir�����5}��0v<�е�V�	�gS.�XwڍE��V	e�vӾ=9<k5����f��P�6}	�]�<Nr=bZ���z���6��Q�I�jJ�X�{�j��n^rmt�4΍{��d���`����@���ԯL˽��.*��Td�R��}/4�l����kVgc�J��C�?��p�Qh��o�Wem+���9�6H�"��t�1��ג�'<��q6r�{3&��]r�^����wG)l�mV���O��{��(����^J�#��6¤�L�fgr�o�=Vs�˶W>���|I����b;�Բr9���g#�n=���SU)��rZe�j� �!؞�2�fono�g5j��v_�VR'vk�5�N&����{҄dƫ����x��1E����˼T��.�b�_Tն��OMm�4E�6�T��|+���Ί�,W�f�`}�!v	���J|��)n�+�Aa��ee@�G�Խ�gc�G�M�5���W��L��d.����Im�6x���e��űViB6�;�J�����1G���_�1�JU�[���Q9Lǔ�b[�E-e�n�ȕ���w��WJ��e�����ct([3M�����qQEEx�������<}iؼ�gi��q�������ց�YS�ݻ�n���u���wyV;pfJJ���&�z�k�Me	����m�ph}�	4v���L��)gU�sS�ȡuY�0��8T�-��[��Mz��^�`�!��7�cf�YՔ���\Wr��l�ح���%�[j�緯j�Rۮ�{�&�����V%��LY�В�WBWx7hVM��Y��1CS��w{���s�/A4�����Ni�`��3h���Q�ꃒ��FcQx������Ll�f�M�[�;_eDͪ,NG�h������l�)E y������*_��"�@�A��"�I�r琲��|w6A�gT���R���x�u	���� ێ�����ƶ�����}Y˂��u��X�r�n+���ׅ��^�a[�Ԇ�쨟4�uU�,4P��Y�,�W�mh����R��e=��
���;A���(�Ҟ;%��w¸!ZV��n�
�D.���Zt&Sʒ��#�3f+e�'fV�[G��M�z���;@8��{t�j�}a�0p�vJRf�t"R9��$HQ�j�#�v�*ݫp�*m���0�x�k&Gq�\�%��q1ύ�B���Tޭ��U��F�*���<�ֶ�>����B�+�D�W���Y��!2f�ܝrY��;��bI][�9Q�j�.�;Qnj�	ߖ0�� "|�(T<�rۼ�����5ͱr�V���z{�;D!z�*B�%�� 6m+4/�>5�!h�G�`i#��}��Ћ�M��e�й�P�_UBN�OR9�����G"�
���ɐJJU�L9E(�}0��(��I×�ϝ̗ğ����#�Y���g.UZ�vd'(�rC�-eBg#R"((���I��NE�w*��U�ZDs�8�#�m9E2�Ȩ�@ќ���QZ%Ur�D��¨��U~?<Gwr���(�4 ���"�H*�2E�\�xC��ź!�UtȽ�����B|m޻�QPӜ��TD9�H���zV{�Z��Rg�L ��
��"$���r��j�H��R4J*jEw���^�X겨-H���8r��!T���t��Bh'y�ʈ��ԋR(����R�G;9<�D*��Hp��ET}aH�[��/B������0F��5���[�$y�2;oz�=+@�6SZ�FP=�����7�>�Q�����}V9\&�Kr�O5���^b��u$�Y��Mo��T5[8��#�o�+p�Q�6f�����~��:^�O}YǨ��Om#���yo�{ƫ}��_n�˰��h��);��qպ���_�j>���=O�+[ x��cL򴒅ʪtM{d�����=X��G�^�Q�/I?����T��P܎/{t���4�b�B~�#�P�oO(}Ҏ�}Ny���"r�+*W_���P�W�;=|p#K6tަ|&��^~�f=1��~�0a򁚌�"�۔�^�hJ�5P��d���j�tn�����s�Ow�ca�sƤ�˯eו���.��{r[�}Pŋ����'��Q�d~���J��@w�����{����
j�A���}��)�a��伽F�{�*o���+�^��	g/v$���
]��˦ks���xu	�%����iXT�
^��]��������{�G|\�롵���b�r{YjMUɗ3H����^���O��2�V.��͵K4H` s�kS�ޮ��0��Ɏ*wý7�FsCwT	4&�gF&ξYڋՊⒼ̶J2��ɜi�&��Չ�*tv�K{�Ak��+9b�N,��Co��o�7ɔz�+0��`��mC�ڹ(өaW�WaJuS5�R���{Ul�j�DourvG&�p=�^}s��fTU����<G�t�����j]��R:q|r�˰���X�����{��Wz����r�g\@����8ߧ�����d��c>�9~Ck:�v����Bhv$���q���j�ٳ#�oU\]b��6H\��Ľ�4G��:@5�k|*�gϽ�p�ϧ�*��I鶫����t�!����V�=�{���j�E����V�U��2jש
��>�|��@�mߌ���R�����Vz� �Y#�!��7%m}�j'k%^[S��Ow�K����Ϊ��n���ly|��]�b}Yh�Ϡ�M�AgM��nѣ��Du�*.�9��3�k�]A.W`ͯ��d��D������ݝ��\�]NyL+:��Tϵ�Ϫ3�{�>�w�y7���u�hൡ�����b�{i���671E�;��!dI�k���l)��s�����<�U�3�X��]$*�n���㋍`���yh{�����B���o���z4'Vhs{�6hc`�+���|?���׊B��"���7���$��aꊜ�D�hB�v�M��4e_꽯#X�z#�|��5��9�~�$󁿽���촵�u�@=��z�S���-ˤ�Jx�<���{�?-��������Z[��ɻ�����^,����eәt�
��&D$��O�|�6�/e�?Di5~nJOݣ�}�Q�R��7��S^�3�K���4i��\�w3�1��d>uùr��|����l��Ɍǵ�ռ��*v*�zeJ8�c��E��O�-PM�w���]B�I�Jz�ы�E�ᰰ+�bRU[1�u��o^�"�uz��[�tn��9W*CR
Wi�#�f��+��V�	[���=6Iޮw�@� �K׶�7V{�� �!K���{z�)��Q~�jv�R�Wf�Q�]^�Tv[�KMl�==��t�r�^�qQ�	�>����lC+��+5�Y��g�ۮ�W�yy�Ғ�y�^[���y���=���2Ⱦ�fQU��?<z��V��s�A����\�7mY���+<��z���E=��9��u˩_ p�Xe�)��� =Z��Ejϋ�ANM�69^%�����=�V����o`qۅJ�oo��z��h�gc��P�9_��;8�=�g[�.�b;m���Kxw�|9�R�ۏ|;s2h�X��<��ϱ�kh�ռo�sN����I�d�����)v%H����jʼ��G(� �;9��9f��o�]�]�b�n\hW��iIX�+�T�ޤw'��*��:/0w���Z�C�BEF�/OW���{�;���\��|}�&dh�<9u^�F[˻*�/I�w{����S��+̳*�Ӽk>�l���.�U�a���^7�z�����v,�v��y�P����>�_C�mE�YG��r����;�1�>�z�j�l�}�?!G����f��G��[�[R6iz����%hO��������P�{6�|=�K����QL]&�{Xy��L�JQ�^�S�W��`��Z�a.�+��M�f�̟?sή�uJ\��z��U���v�����%ؽڂ;Yؐ��S�iV��R����I����o��Wq �5Ue��P����Ot�%l���Sz\E�Z}����Q�K�8��:��F�ջ��
Ւ���dV;6�u�}�^l���V�Vh�mAO�Tk��u|�Y-#��m9Y;�$��R�M[���%�QA�&��y4!.�Ո���aA��"�}����^����V#�?{�9jw^K���/I�X
��Koز�z�b��	�!��'{�++Mw��v�XE�[nzT7۹^���H��>��+��O�*OzRSc�{\;�sW�9��zD�0�H��W�{��>��R��}>��4��o��j���CB����L�Sz��W��Wo��������z+5I�}�D(߶]��޿m�A1�Rg��A�s�'Bs�_ީ��/^�U��>���ߣK�9��9J��^���fp��c܁��W�%!Cs���iAu�2����ݯ��[<�k՚�����fC�FHY%!���}���ݔ�������`]�zwo��7z�s��]�yP�׺"��eJ��,ʆ����.|7�%�ᇥ�W��K�ˏ�ԇ��Lk�j:�<D(!�:�Rb����*}���G���בwA*ʊ�P朑�����~ݮ����*��|A�f��}�X�}�r�8"x����Hԭ��l�ˬ�D��p8�d\W�w�͑�+]�a2vN��7�^���6p�%[�㉃�nԲr�[���:���fNݫU�r ���\f�P�����=!�8�]Ek�hu�|W��te�\q���ב�g�1t��z�z���[�T��,��7�{Y�YW���VQx�%@���qq�m{�i�Iy�:nƪ,�䫜�=K�Ko��N������`�{6�r���Z���#�5�RS�ԧ��|�2�ס���S�j�zr�ms5�i*Om�v���ޛ�=��1��O��ə��[���=P*�8��u+�7��
��ݷ��f#�T���9�HjA[� x��ɂ��{�:��쎲�%i{Օ�d��<�w���ׄ���*�,CWDx��f�R�]Ub����c�WI��/�[H���]�a��g=�qz�7���~\�7Sf�.><w�x\�bg�b�L��̋k|W��#�Q���������@��{�B�su/6�s4�F[Θ+6'v�������ti9w�l{:[,GR���z�N� >˽�`^"�^˘�N<0bB+�f�N}��4:���>Њ�(�Qq9�wB��ͮq^�û���tų����0����)�̙Y�sټ�VMQ���ݑ4ϕ8ޯK�~��~��Q����{mf� *[��N9�;�� �*Er���em�29z��ʒ�j�^�n�����C��͍����y,������.U�ͨ�*�@un?=��mb����=9��gJF��L������������M������U��l��Ç�bDr������!�����x=�`��~�������L�A^�V@/�t��U�>��5P���^��3r/���O@}�k+�A��'�ȏzU���){��7A��s.���%�L��&���}x�����W����E'6s��=�����ϟާ�s�/G������sڮnwuIggS�$5�9\^�[U�f����?!V�W�A�׷ެ���'aN�w��Hz0�t��ߡ�׽Q{�yV�uc�-� �^��p��z��Mb��L���+�;�V��\�y�u첼�x�6K��+y#8��&i�kW7��a�Q�(Q�(�zIMڬ�����zTV�[t�|�8"��ʹ�iu<�ƙ�fc5���`�Z(j#���w7��n(��r]����j)ʺ���!�s/�����x���U�W�ݦ벟{��<]^`cs7�s^��@:��g���{���z��z��9u�1٧Ew���s��vU={�L@��T�߻*�Z��x���}��$�3=������h���RN�S����N�J��Ƚw=���u9��}R{�I+�ч�y�j/W�������dU<�
�y�=�V�k�����ZY��\(k�WEvHj������o��>�LU�jg��"o�vg��u=��n?	��ԝ�^�BoWl$�q��V��g�=��v��Wo=�RJ�|3�8H��l�6P�^�{�;���\��*_��T̿e�a��~�4��;1|%��`�[@mp��^�F�R�.����-_��]����;��gw��ʊj"��o*�^��Sf�>{P�2����� ��{03}t*�V�4�q����8�7��Q��[��l��*R��{�}fz�픫p�M4���%�b@sBh� ڵS_��s�9;_&. �� �r�i�^�ص���z�s����Iz(^��:Kt�&>�~{v����u��#�#��uh��b���/0kf�ٳ�~W���]���I�Uמ?��w�c��Iq�ӂø���6��u�C[��o��۔����Ԥ� H���#r.҅�T�ީ���Z��'���^���g��4᫋��{[Y[�9�S��O���sr�o+��H�O{��uΟW�O_yw!�C�$\o����?/Լ���T��J�)W�h�ϾD$�tl���ვ�Ss10{��hFs��}QM��	��{lyb��*t-�a���Iۻ��:�]����L���mM��y��]�ðZ��l��@������K����{2#cd��yfb&z���)��ޯ{��_�`ٲ�j����R�1o�D,�/(3��ޭ)z�^�qf��s��^�nyW�����"��3�w���,��M�����;�҆ny/I�,Cy+]+~����+�M^�\b�zc�����1�X�]�u��b4����d#����bo��,/bRƌ5ձu8���;�qG���	���3%���y�Pe 6�AUs;��(��ԂW�>V#�v�]�"gO���-�R�&꫘�Ab�eY��;���jH�#]ܐuF�a�C*���h���7��z�a���z?��A��szOV>k�w���I���8]zY��Q���:�����|C��%:�4z7��4Ϥ^����g����[�ZG�RR����T�X[ܷ:uLO�����rq��/}M�����}<�#�ɆjeS��K~���z�HT�|����M�ޚ3�f{�E�2/u���o��I�{.��ZhwZ�����qc}��>���)��#=�6�;w�=�73Jݠ���)#���3�QJ��#d!=t�ͺ��=D�o���~�q�o���nl/��c�V��=�@�)��^{c���
t���^ϻ)q\��=���j�+k�	�t5F�G�6�;�PJz��U�#�u[�aW��%��zyy�/ݵ��߹��B�����m�%�r��ȨΧ�q�4�<3��4#�Ⴥ|LD<=O�x^����Ak��"!��'�fe�ⷱt�`��5��8��j��b�k��n6<r�����s�)�s����&j�槮nHx'��C% �S�������>��ßYÀ��c���sw@�)����3I�t��f����9�Q�q�%>�Y���z�Ȩ�7���T[o�����n^f&��tfL\��p;�D���5'Jܘ�(ݛa��l�~�W�i�W\ �Z��������Zm�fޢ�O(��h��`��j��+��|-�LN������]I��ӫ�}->&0���;N2s.I���)�4 >yte�h�N�d��m`6�����'=y�ۤ%DZ�+Ir���u���ǩ!C���PV_D3��C9%h^�%����o.�2:�:�¡�����V)���y�[B��#j*�U�ܛK0��ވ:���]�ûG�oZ�L�\m�[E(&W!�/Y���1+��u;��f7���WT�����P�ȕ��;��Zݸ(�Ւ��I��Vg�D��ʗ�+�s[N�ˉD��A��r����N�U��Ҡ����3���b�:�.�+r�b��юJL�M��-u�"�!h����D�d�� %����7�����K�<��+V����8�z�kANǨd�杤��0lF
�kN���D�Qn�F�J08s�H�K�o��]�^TQJ�]�}��5�ҷW)oi��
�+F�WlY�d��c���n�z�ᗖF�J�q�˧MS5�mGiɂVS�{�ͧ�i�tJ:Ջ����o�������J'�AFIX�n��S+�Ԕ�[;��ƬԹn�&��9��{#�{�Ǧ�ۃg^�[d�VܽE�{#����f[��=n�ݺS�k����f��4\�����܂_er��������,�坿IX��ȉ�~��^]�i��m�[M-&��Å�?��@�kb'�)��a,c�Q�Λ(�����ۜ�׆�����b�;4ٌͰu^v^�q�y�FF�3��%�B����[��+������ħC���sQ*�L7\�2����˲�-�DTY������w�����;n�&���D�a=H��uqZ���l���Q݋�Jۣ�us��cS�ܬHb�"Y����=��2�BX���f��,���W�
����Պ�|:!RP�I�eK
ZNd���n/�R��r}p��/,������������,Q=�U�˧�>skD�P^�
u��,f��R�� ����rb��ᓵ	X�&c��^�n� �Ӆֺ��ظ�	�6.��GUi��q�o�&��yL��*���v��&�*�Д�@��e�y�g���e���Ytjf�!�ڟ]���9G#�v�v��eԛFaܷ�̸�)�+Xȁe��p�>P�`�'�Mn��{�e�O$}�o��e�t�C}Z��h�<T�Ų�Ѯ2t�yzl[��5�L�3�?_~?`�
���;촣��Y$&Zb4
��B��Dr���"�yĊ�tFU�rzT�'I�g�\�)��UE���E�J�H(*����s�ThAp���Fq8���r�^d®��E��"�����"��֑"<��8�C�p���WH
"��>�
q\+Ԣ����C�S�&�e|�**&QO��\��Az�UQ��
���D��ӈ�Z�^r�.QE˗z;�̢��ނ§ø�D�����,�#H�.�j�
t�TEv��.f˲��@Qqi��Gee2%^�*��*g�J��Igw[�Q3�U\�������EDW)���P�yУ�\��Y?�������kn;I���񃷌B)��*�5�׬�r�yl�0��<:S��f�s�XaTe��5+�}��M��ї䫄��q^�nu���U�@to�R�7�bCϬ� ��?Pٛ��=5�VmD��U�X3m�.�`<���%E}79	��i�������jש�m�9O_f�3�}9U�=;�
כ�x�L��Y�8
��AK���{
z//�G�g#Su�-�!��^�����'����8�����/.e��ͬ�~7�WH�px�8F��z����!��_.b\zc�{�(E�����8U��ޚ������a��(��#������*�l��A��p|�Y�i�trF+9�l�E򚆎6����ո̙�E�9����.6���b=��qA{j�~� ��;hץ�c�(!�)3L�|�2���ڧ�����>���p����:R7�ie	��g�z�g���Q��!o�UT�[�ǾS6�~�v��E��|���>R;Fx�Ew�}�`濏8;��|P�u��:�vߣ��s��e�I߹N3�Ą�`�+���ᑥzK��5%��;�{���z0IC����|pu��; �;��Z9徭Ai�_�c/d�ՄV�eAu�>Ka����q��^[EӀÐb4ß>�GTxU�,���f#[���&=C!��MѝgZ��o31be�[�Y��2L�c��v�Ж�93/R�me��Y�.q��6���1G���)Pd\vZƤ�V[TX��l��$��yﳄ%���^��C��,vˀ��G��u��ɉ��0����a�W�b��R*�u��=͇��0��3�}y��n�q�\y���^���[{b��u�;�}f4��B�H�Q��}�/�͸��y��
\�S��R��W��S}���c����z��~��^=��+��''#�ϝ�3���X��+l�����Am�6��g����${_�GG�
ګ�+���CA�z<.+������C���Ǿ���:�b�n�>qA��"4r�W(dl{0�<�g�Y�M��6�? D��OA����:�c��u���EoJf�lR��J�.��j�%�9�1B��U�����^�ud�����԰Rj<�������3��yИ�~ȫEw�UF�^->��OԄ&��tmd;���f��20)�-�	��9��������{Q���^��y��)M�XJPgc [,3x�T;��
=�#��9%X�0�g�|f�鎨Uw"A�H�>�u�r2��az�_�Z6�b�F�h=V-��v�d[�Ȯ��.̦�V{B��O?^��޾"�>�z7��z���ED<��f$���#0�0jV2���kx�RM��Wm��R�R������+đ���W9*g��5Nn�r��xLŘ�Ւ�v<W7�6��m$wY��7,�{7�x����.��n�s&�rS����CY]KN:�J�_���Ջ��UDeє�^��}³�B�2᳊f�Y�n�<�i��棞MF��K��N�`�s�e���O��^��P�>�SPڔ!�uD!r�u�p�2'4=������"�cgsUα]�+/S�'��������zō1JPe�����ם�v�F��Įcыj�x�v�4��#�~FGC�dn����UJ
?_���!�=Ƥ�`��e(cئ�4^T�Vǹ�O�Ð�%n����"N*��rt�_=��-�&#��8A���`��*�����k!u�{�����#�ij�cKH����>��T�`hg,�,q��#�s*��l�36���y�c��pC*;�WP�����ǀOH��SӁ�H�e9H��OBh^���B�O�]>�V�9�*D�~�#åG�G�^u��JG&�'5�71�j��Wk�(T�>�y/I�u�<�b7�@*L�R�����ۨ��������D?2�%�rN��:�z��yf*�^6�T� �NB��2
5��a7�|�Mͳ����h�T�m|M|z��,�/ z�t(����z�?�f�/�V��5h��hgE�R�m:��/<{j˘��[,����D�t�ɷ�54�(�;��uM�.R�����Xw�P����5l6�IX6P`���0Ȩ��V���S*7����U��qIg�{�;����7!���u�-!��0�����c"
J��2r_��q����+�o���p�핦���`�Z��ͷ�_�+�+읲��꜒�t����!xT�3����w{��zA�z��W;�m�z-s����b�~�ov��{��P�{w}�����b�v����>��?xOG���Jf���hŎ�l7�wP�9�q��A�ƨT	DM,��i�&y�����S�j�.��l1 �}��E|Ȥ���쯐�κ8�.8s{�F�s��b=-x���c0O��7�|e�|M�>��>B�w�B�>�.zP���X4o(�G?�Z��/a�G"�7	�N��,�T�cAؑALG�e�|jw��a17�.�~|͟?�1EK�JM�\U+�`q��a�\�Z���ؒ#L�B�段�,Fяo�F����%�(sbTz����(Rն䋿�;�8����'*��'��A�/��õ�E?�EJ��������G���
ڶ^
U�X�^���'jM��{���[��~=/S��MC����X�`��*ম��A�� �^K����M�����˯רνʔvA
5t��QDL��vkn��/`��t�{9^��ͫ�{ �m>O
��ѻK�4+G	�r_7zqۍ������2���v&mKm�'�J���N������y/�.:�>�W1��A1B�t��������k��Q��[�@˩�B�۽�Y3�=��y`�������T�z�#�9 �T G ��O#BLiq^����}Րα�ʣ2"׷5ܿg������|���Js*5�TC�8 ¥" ��P�Y���GX~;�k�gbX|�]_�W��a��S��T"b�Jz�Oԁ��D���7��r}�	��&~`�;I��bYr�y۸ǅ@�� ����w�iP����ѾR�6������ч�ٛ�Ԗ�uE��z���]x�p��x�����M�Cg_
�>Z3��E�k����p��X�H�gk�ce���H/��oLΕ�/ư�P�8�� 8q�o���)�W���5�q�X��3��s��*��f��/9�
��^�l{k8ߍ�c�Y3�FD�-�O���zi�o���~�.o����~��k%'+��zf�P�r�W�X]>�7��L���a��xM@~�"�6\p���y���]�}�g�`pj����Pdr3��'M[�ɞ��t\|�&h)q�<�s�cJ���Fµ+�L�[�v���G5.+\N	+b�q�8c���U�u����S*i��m-�o�.��\��.��?'k|��J.��-�GsRS�#�c���J̵!.��_on��2��5�}���Р*g*w܁K���O����t�v \�5ڨ�a���Rw���P6��E(�h��e���2���m�q��Oz�,NIwJ��V$xvT�������b�LE�J������~Ub�H]N�(���N�зoo�tyb����ӝ�-����TM����' H��~�P�b��G_ݵ�h�s1h��;���`�f���7T�T��B��c�X�F���p&�P=_@�@U�@�T���w�Qۊ~.���O���E��֡׌�;(z��=���9aM�:v	�1�@=���g�U
����4ϋ�3�h{�����y��3у�R�X-���˨��ӄ�u}��H`�1���>�LU�]ؼJ����4�/�s��j��t�pGa�ЗW׹�)��G���&:�`G�Pu=2��0��%���yO
���7+�r�Q��0�yu	����6BM@|�sj-�.�c{��H_�g�xC5pK�Q��ҽ�C���hy�[����n�@k�rt��w��t�����o��Xe��L�Dƌ=&�/�}e!����;���"4��V���E��~�j�m�q�cY��D���/؆���~>�&��U�tD��N��k�h� Õ-c���S=ٖ�W0n��]�����x�Du�^QR�I`gT�� pd6���[��슞�������m1w61S�1��0I�J���yf�ν"�U1��l��a�mdς�T�@��r�>��<���\;���o�[�}Zgy�05��n!ze��~	����5[���~"���ɟ�)�	l�Y�����r2��~�O!珠s�l��ټ�ņ}�Xf�Ȩv}~�j{���>K�k���r�韬Pb_	�*7>�6�_�naǤ�t��O#L��X�>�J�ܜ����������=����i��A�B{��e�FL�nI��Nq.<�i�����<|���'QY���*�xW~�U�Co<�Q��b}��%~��Vr��u�p�<��o-��'鞵���}Lz/ύf�r��N#��3���b}��렂6�EC��I�)T	x��1y�aﮟī!���2:>���CV�q�z����J�|xb�I���Uu����O(����X;m@��>31e6k>N�+�ψq$�v��v;D�/Nc�fUG�cn�K���M���/>W�1B��/y;P1���WN����a��N��G���L�U��E��U�-���$�8;����Ds.�/��KIΩ��=X�b���XT�NRA&����A�t(b�=��m���us��^�����z�N:M�p�b�[�4�x����3�sdoU��6����̹��{f�s}\7Y��JE2��u����@������$l�w]C�o��c9~#������#����F߱�#�~�~���㕁t=8	u� �����bA�*�]D=�R���M�� 3�~)�[*C�ڋs�F��N�K����[u�*����Q<Ɖp$d�Ќ�����yv�K�b����/l��e��XB�H�n��s3�h��}# �_i�g����hMͳ�g�ӽ5#~�bNwtw<������]fx���.|܆Pk�ax���0����R+˓���[���`�����s�ָ����������`�Z�����Ň�F��ܖ��&Q1�ZVT�k��g��ү�]J;ƕ�c�}�.�kC�΃Ӌe�w��-�v���n�X�H�a�W��i��@�ꛒ�z~�2���W�J�gH�c���o��(�y�q��1���R]��!�l�v�Փ_�!�O��RwV��xf.2`ANE2)�R޿���uѹ��QGW1n�,SY��N�o�0�֗��p��>�xޝ�r<O��h	-���EHA���'��eT~�_�:ݯ"{�+%_hN��d�
mdUt���ti&cҰ�V�r;�Ⱥ�v��E�����;������@p)5me���G%Gҝ��:��)H�XpJ�d���AZvT܍�����ˮ��lTeVj)]��ZIǺ]:�72�d��Ի-��|�kEu%�r�*��p{�����/Ц���#��6���7���e}���"���v������@�۽q~��[�=r�m���/[�Y�l����8�°��c�OYTo�2#N��M��BT��~�W�=��<.b=%��v+�8V�,Z��ܑv1;�7�)�z0'*�RzUr3�r}���Q}䪭� �rP�?wУbı;u�l��YD�)�|�t�1�qU����|l���w��w�o����#���Gl�$1=P����OmMF�֣!�� _tA��֌u���;�j���<壖p}mR�똎Ч AP� �O#RcK�I��:�[.���/B�����%]�x!�Y��w�鿓�Qo��6 �DDpD�Z5/,f�9^`�Fu�Z�C�7���"�nЈ�R������Q#�a)���r_`���ʎ{�=+���~��/��P���o���Z�q�>���+����������c����<�/���o��݈�Irȼ��}fc���x�𛜆�Q�6�Ӎ�o�DS��;��Xb����y�MS����WN�#,��N����xz��ņ���p93���������]��{�Q�X�s�LGJ�J���|j�61ʲ��篃X����{�uEYcvp�~ȣ�;��Ϻ��]��\t?q���v�a�o/�j/���������T�Y�'����6f������#�TR\P��{
uu�#�ʫ�cSwԺ��Ċѕ裏����-��^��i/X6=#c��.��� x�#h�����u[�[�ײ�8U&=^���B}����+cs䩈qcU����W�X]>���9'�9�3��>J*x�����Ap,<�ʶ��	��X��R���Xd_ܦ��ۚ���q���9�p�s��|�q��dz�歾=�`L�1�=vD�8�H��e��3L��M�-�q��Oz�^	sA�EZ��s��&�� Hو�)�F�V�v���Y!u:h��m��8зZW������ݣwj�HU[����>��Ё9@A��~(K�����mdZ8>[��.:Ovd����'��8��U�c�͏�#C��\	���������q��1����c��bԣk-/����>�r�9�[�p:&����`r��a��֦ɉ�t��
��{��g���w�JL�'�7aV+J����������l�`�T��j��]Dm�ӄ�ut������<(`�x�9#��,{�v!�G�v<�9�=EL�Z��"W��m�KE��������$FS�����+� �_���(�Gx�f�3��YH��ꜙVm��:�F�흘"��b>ÅC��(V����.`����2�IX�w���kE.#�=��@�os7��l|l� �Pz�9��d�֝���72k�Mِ�$eN��ɹë���6Ckj��6+���T�s��kR��#X0�L�Y�����cGf]rt:V�Q�d����3� )d��E[,�׎�A��F�䪘g��,�*R��<-�[h�+�j�cՍ�� ��I!޷�,�-oc2�s^��i���U�ژ�ۜ�E�!5�DTU.�SaЦ_E�Qe�ovJ����L����T���QЁ��efb�٧y𳶐�F��g%	"��#��k��s��d������X�5���#q�|Ufl�����j,b�E��c��K�܋�Uʂ�^]���쳝�,Ř妵���w,��x6ul���,Ѥ+��1p-��X����D�|�E�=�Oea1�4�l2� ##�e��i����:��յ�Jͮy��ְ�\(Cn�D�7xf��L�k6��֣k�����_ �ad��{�)51-uI�_dӽ��_^Z�7Y��ρ�QY�]�@��sQ\�(�vB%�]ug�f�{�wn*}3%|��bw�JX*�;׎D��B]9��dL�����_\�MBEq7O/��8��M-˹���9T�2D'RR��;��&j7�7㲛��ʅ���s=�X�ʔCfM�j7��s��M��ѱ[�p��W�Ө��構�k�f�ܞ��r��4�X�)��l��O�',ԽT]*:	7%Du�vdz��q��T��C����:%*OEF�-%55���[twG+^1���鳲��2�����PT*��T����[vn���)6�YDl�����1o\\�](ƙP�V�o�sE:B�aɱ՛��R�2J�9�zk`��U���st*4fΒ������m'��B�+�K�-��V񭐦���0�{����CSEs������{�ښ�d�(.��]ۗ��	��e3Q����m�B�K�wu^6#��wIq�%I����P'���TM��F.��jI�����\*'U���8)r�n|
�b��}�K\��Hx�RP@�0-�I�1Y���g, �nu�Þ�
�j���b�u�������־��3�4�9S��
}�Ը��)���������7u��+�ǹБu��ǈ�{qF*��6�i=1�n�.��Ȣ�4Q̦�E��+E�=�9	�䫷7$��:0֑�byw���skC��"��z�C!D;�j���V_)�c��ppwl��3e8����&؏2�7
�Y��4�cf�=I�.����H�e�)kd��-�:Tmuj{:U�Zm�Ai�&�t|嫿��}�����˗.U���%�.�
	QQvG=I�ʎE���h'"
.�H��vP�y48U��At�*���P�vTE(��`PkB�#�Q�r���S��
c)*�����%q8��
aDAʋ��dXE�X��P)+�$�"�Y�:�+$�Γ�r�U���*��;�=�2�U6PY�v�Yd\��t�"�r�!�ȡEP(�\�u.��H-YT]�Q2��j��$�٠�ӂ�P��gC�Qw2�'��;*����T(*�.5�t������S��F���JX'�L���r�^BT�$�$�� ���8�Ȋ��Z�8p*�E� ��]'Α���>g�pM޺�R�Ƭ�vXaS4B��\�5d�Ni�(��/�/i�kQ[���[� Z"Z$dv�X��pF�� 
ݯ�ꯕOQb��;P�a�I�+����v�j�����*��K��ܥ7�a�~��$��|�=��^�P��C�0���>�A���:\�~]bz���j���b��nmBڿj&R�3Δ��Y×������8	�0d�bG������^�u��o��q���n/�f
��D+����96��8d渋�ޕ$P�q��Xe��L�D����7R�}S��+u��qY���7�>�j�ݡТ)�����E�4�b����l#Xe^вdx)�b�譁g��~,��� ��Tc��?Lϩ��iM�-l���b'��'��2��d?pY���j����m_���-������q���������ls�5q�Xgc>e�o��m��
=�#(��W��c"��	�����!W���Y�f/�[=%����zs��/�b�;� \f	p�u����&��x6�޹�;y>�@�?g�]Deі�o��:�(�\6yL�+��\��Q��}�s��ad�ZE���z}ޜ�W�W���EIl[R�;�0�P�Tc��^svMԃ��г&�޺@n�o0-�'0#���]E��(�]�N�n�e-��C��>خ�w2���4��oj��g����Z�˔���M� ��|؇�y�vROi9z7CE\�eO�����Nw��۷R%�%:wՆV�S�c}.T}j��	J���Nn�jG��^>�}�w*����~�����o8ж[�A��>�0+��?0��+�(3�]~��w��{kј�y��t}�Lk��+�f����a�Cmm_���Ɓ�,���i���<v|뼴EQ~��w>���Z[Ngة񘱋)�X��с��&"{�|c�kZ�N;cUv�cq�
s|Z��kJ��g'J�WB��{�g,��67{��:���ލ�V���lG�c��D)p�+�tm�r�� .����S��H�<�]�v(D�W��3�u��X)��8�%PR p?DK=$2��{~�P:,y7aX��]�*�(��OTV��>������C���eUB���H:�y5[��n�,k�'� ��(�Vm1���{>��y[�#�摋	TGx��U1KD�."���,"&�O������
��P��C��֪;l���mz�'���zqW�A l7!�k�c��r���0�dD`ޏ7�Q�<&�^g�xH�9��qoޤ����r0v��c�-�QazXf��/�ҿ��vˍ��5�(wS�>�p��zsM�ϖ����J�͛x*E�sΒ����ir�jj�Ss�˕�Zw�̳�������c�2�K�V�B����)�[Պ�#�RR�9�YYI�B��Z�$��&��2�pH��=���e�[�!�4�F�-��WQ��W�_W�h�߼�B���i�?�%��0�>���|/+��Y[u�\�=8���[���2�3��Vyn��O�?��,�>�m�d!.=Td�Eq��a�wP�9�q���I��;���&����H��e�'���
��B����O��#^����� ���.�q��ъ�}�>�c��L�}ʜ�B�O��7�|e�x�d@xw�-���k�j��[��	Y��gT�1����Pުl�#5�7
�j����g2������dr�˓q�F��y���n#\��^66�V�
v�ɯ���p9Դ[f�=��
zʂ.i��Dv�
�&�ց�#Lȡ�#!�	q��u
��Ki�؝������B1�6}�b9��bJ���a��P�� ���;P'�0�����SH�S�/%��9;Rr�{�M���ox�Y�=Ӵ���ٿ��gA� �bz��t� �����ƼJ.^�ى�����dL<���g5��KN7)�MJ���*#��yP�p���2��?������,�O�Oo�Φ�)�B��4�H�[B�]<(��Wiap�9B�&��3lli<���)]2���Sl�2[�/Wf#"k�sf�/Ru�z�����7o;(�r���x]�Q�$z��Ȁu-B���9,a'.j���{��c�������q���x+�n"x��y�C)ӄ�9�>��}^7�*��]���8 ¯���� 㻡C4�Q|����R�N����NM��|�"���_b��d)��69D�������ru�aW�C��WWO�ⅼ�z�~2�7F̊�}n�χ\�ҡ	{o�)��)nDM�$1C�َ޺�5��^�ڎ:�i��Lܞ��3�\T1��nr9�>Ӌ�.�7��EX^���q�^қ&��,��/Z�,P{�RAuS\�qp���e~���ߩ^<��t�`ބ����Ĝ����1������(�`5\!㜀�~Mz���f��2�u'�E��>���K�W4�y_:�"��N
�؍�ū�g��kW7����X��i�>�@�����(�a>a��[#re�.;��H;�V՝���[T�����w�İ��SP��up�
j�a=�#�r8$5�w���2&s�]�<��0)����F#�@~�w��,u/&Yl�
f�Y��
�j�dE4Hר��DU
cyt8����;{?1-�F����0�H�[�ϔͲ�.��ʇ��t6�ol���q��}��D������y�M�l�p�j͎��f��*,|f�W���y�1xt�z���"�w+v��2�+w^I�Ύ�q�M��s.���5�؃}uw���A���B�Ml�mE*�+X�NK��{PgK�sS�6��ܑ#<�u�R,++ﾪ��뙽���~?s����]>F�>����0�� �.:�m!c��-�]LK�D*&k&#�k1�3㶔l��9ſh$l>F�>��>]@�@�@_3ђP�+�a��ϡ�a�c�Ѽ�'�Σ��;�����Caɴ��g��u���&'~c�*q��u�����<���q0�Ų��T.�)^F`ަ�F5J�/���_ڡ k�(lR{Z��ۧ��}���A�NY�;Y'��k������].��r��E�+���wy_�u˼�O�/��C1�L8�?h�(O�cQ�0�p������B�j����c���<�-<}~����;��0�>8	��:'�ď**}t�����k�?+q{�{�W0���WꈜpsϺ���Y���PJzH��q��a�m
&X"btd�T��e�u��a[�e��O��p�
4ҟ.�>�����"��#�z��S�c�2�6��>
ES蘺�l�Jʾ�l�V^>��]�G��������k#V�`�^�!E�������~��v=# �\l��	A�z�ߦ�����f��g��ޚb2I �CF����
�n��=w�y:�<�0V�+�BZ��i,z�Vu���^(:�]�1U��]������A5��s\8TXF<7W���pw6��|n�U'Jٙs9�D�ȝ?�]�eq�;�����_߫꯾u��_�������΀�Llt뽰�V��X],3��l�NH�"�������CR}u�Ϻ<V�O�\��}'�DC�äe�i�fы�VÏIh��b���y�z��1��N�Us����G=�Z�7-����+�cnrOa�BT}!ʨ��2ً�}F8PΧ
,�q��7.��x�߶U���FJ�yShZS��̞�@���K�:�H���6�(CܓD5�^`�����3�n��&��|�#��b2��CG�KO��������}��:�s��ҦϘ�ŌR*���Vu�f�%Y��������5�	��ƈ>��M�*G�'W�۬Hb�1B;ۛ��_�Z[Np�O����l�}	҅��`k2LFe��˺�M��\>�G�x��������������
�cKH�N�c��U���*1`o=>R���=Ì��}q����6ѱ��\+�:6���<��K񋞏k�	`f���Yfu�í����]�U)	� ���E	̭��{��jGτ����^EC̩Y��r�pꏹ��M�B�*$:	ոv��·��lv�n8e3��ٝs�{ߜ悪�j���μ���8P�o��@Ů��Fm���J� � c�{if�mI�s�]�q�Ws�H�ѩ�N�(ˮwew]���.5'+����UUOUȼ�;=���?�A�����	�B��c*,AJD���?h�FMV�����Dn�`��38�%�LG?/Z���1�%Q�|��)h��c�dkM!�"�{�{Z����{���O���9;�j !��8���	�7!����)xNC�6fEt����f+����<D���~�$x]ϴ�gݲ��K`�p^����-�G�5L[/�{�k�w^�>���:"6�x��.�.H>̫E𼮌Y[u�\�=9��bp�k����c�d���U��ǭ��ZA��� VTܗ{7X��Ts�i����w��=�r�x<��Є^��>�v�Ui���cj�C�jų���3 ][��o�Y�1,)�p%�!���=^}r�qȣ�z�A�?�Cʔ_�P�	A�W'N��Zv3���i�f��������S:�ݟw{C�R�w�B3���2�|����t�&�8zs����s+�R���p��g��1S.F��!X[)���5�6ˁΥ��G?���t)�7�M��xѾ�{3H4_���ZJ��!�80�6��$�#�+Բ�z(�+;����|.'�D�E�,U�ܺS�v�����lh�O���^�벉}�W=[�(�Xxw��X�(�"�>�JtY2Wg�q뗢o9t̣�-���qu	����X�� >}��B���r���Ƣ E������B\u�Pp�nX���$]�N�M�g�t�Y�B�9P��b�{��o�?E�g��4Ed-�v�'� �𝎽��^
U�
<�P��)�}���y�B���kTF���'���n�q~"���v�"~bz� t����W���D���S���������uLds�W��_��#�p[T��~ʈ�S�1*B����<�+��dl���v'�i�}S���VB�N�,�=g�����*���1B�aPR"*�:�}=��Qo=]|$K�M�R���z�2�ݡ���=��H�;�SPZ'!E�ܤ�!^8۹�ǘ4L�.�>�*}n�����ߒ��^���$)�o�ؐ��ʅ�݉���J��{����Q��~zf���J��<Tznr9�\�N%��a}���(�链M�d�2�����yk [���8%*H:3k�5���
��0��~���a�����_���$��ȟI��{��L����k]q�-�!㜀�S^�l{k��xe�'�R�����:;l*Ϧe!2~ɹ��to�?[�C���՛i	S��7[�ߧT�^u,�+���;׏5+S7�̍OoV����A�M�κ+���f�_.�n+"�f�a�6�ruϷ5U� /�]�j��;=˖B�E�n��o�1���{ގ��3���  ���r��4����#j}�����1N7:bO�O�/ܰS�u�7���LGs��`ҊB���{<�1,P������X�;辙a�c��4q�W ���`����%��\i�~�<"}◵	��d���3�����f#�F\މnu$o[>S4���.u��{2/}#3���լz�^FC�wձgӒ]���d�	n�6��Wvр�b�H��ݶv�GDv�}꺙�Z�u�>�~9�8ж��G �|��O�h@����@�ݭ���Y����q���N��fM�9���'��y���������\	] �@9l=$��<Zc������5��Y��>��<_�*�`��3<��61��rl'=��>'#�)�c���1�ĝ֜���Hn���!R.LY};�l��\"�\_���ўj�����~wU��g	���e)��8p^rc�?�.��5&4�7��o�XǅӁ���~K�����!v��=�If��w�ڽ�=bL:����k���QC�;�u�3�<���*l����{oԓ�(ӛG��z����t���+�1�帝o =6׹�B0\eJsYY^������3o��N[�'�J��`?j�J0ޥ���N����;�3彆�Tc����`k���ˬ�������`PY3��n���,w����MO\F_�����| <��������ƶ?���GA������EO������p��(NNܗ��u�V{;�7�/"�ϫ��C�jzH��q�Xel�'"btd�P��l����7�dgD{=���38�/�?�WӞ�qcz�1a:�1ҩ�v1��Xel�'<��~H���:w
�_dn� 1�Ր���+�}��4-���,C��?R&�`�f��ޑ�Y���'V)θ�/Q�%R��<���xJD��7�P���\�E���ϖ��"a�}~�.�!�E��1���5F䧒"�e`�E�噴c�;;�e� �!��Sl�Hzo�p�NN�T���������ݱ`�7%{'�hXr�#&f=���p��Ni޺�r}#oy�N�jP�nf�ۄ݌y�;L����
�ND���}4�A���ԡ�'�b{�7H�V������8G��F�_��FC���4-�o��zq'�fh�1>�Y�#*'}X9�,�����c�F���o�*��:�X�d4_�FGC�dn���D�;��`�c���bb�QH�^e�h��;F�^M��� �G1NÝr�,�^ë�����7:��fFd�O��xJvM��E̊�n��Ί����[Ĳ�m�J�(X�r2��8�vt�x�9ۙu/�@hs����9[�5Ģ��HF�R��W(*��e���+YA�<)���uz�R�Y��Wt�w6TB�#���-�����Ȫ���M=Z���U��\T>���e\�[���c~:�@$�V�t��ś��͔�x�v�.U��ѕ�Ao��bu�v�唪���L���ϒ��G�漛����6偳���������ԍ��"�P3#N��c&;n�a��2B��m��F�i��X��M�[��ur�@-��b����u�U�m9з��0 �{���+�V)�7��^�	
W�p�bv������k����i�6�e-�n�R���Q�ֲv�eQ���z����㬲�	�jwU�������::]rlAX����]j��L���Jq�t�ᑕ�N���;ۥV��Y(���Xf\"S�<�V嶴�� �N�a�{Gd%��z�Ӝ�wG/ǠA�7	5zk�=�˽'�!Yҕ�1�c���u�Q��l�i���ܣ�\�eN�Ws�I��u��i��Z���̺��WV���t*����y4���+�����dz΅۴��X�F��Iޤ9f�˶VM��3@ps��D�#ι�C���S���ܢvT��� �yC�8��H�Y��-�1��05�6
���r�w������6���m�S
���Z{���Gb{�漐��
��	��i�!�oZ�Ogwa�ؗfF��(٭=G7�t7��-���q�懲��1u3h]�w�B1���L?�1�ijx�ȱ��7��T�Y��������%˛R�fH!�FdlW5�s����ŕ�.
�����5�50-x{�ʍ����:��]�f:1�g-9D�˰uU�T�E⇅I+� rC�>����F���E)�'nK��-���vv���ڏt�ʼvvom,]����4�s0k�^M���������"=P^�v����FK�Ӎ�ɝAlMuK�S^e�h�B�;�%�#e��Y���%*oS�]�t�"Eɛ������V�M�.�otN��K��MZ�����I���!��-/SW�^��^{@h���;�>ͽ���7Z
f���w.i��jL^t�3�Ts�f�d���p�]��Ѧ�l�o �G�(�|�ݠ���iOxb��T��p>���m=iꥰ^�p����uks�\�E�8c�v��	Ա^����^�fM�HΎ��n���GY���&���6Cm�����З|󻀥7�\�����V�͸� d�7s�!"��*�@��8���H'��,��J	R\-���ƏR�ݨ1�tWs�"�b����s`y�:�n2��*+o���W��$�$�\���y}9��v��qd�.�Z۩�%��y����~���<���{.�'�G(����A������ΐ�:v�JƝ��LEY�Nq&�@VI��y���[�"��C��H�e�W���*(���Rd�H��ʈ·dU�ӧ
+I�!9�dQgԣ��"*�@5|�����*:ABe�L�[.�	Ҳ�MQWI:mS��i�L5bd�(��QB(P!'9�)��2��$��M�3���+T�M 5��r�92���g�̔HȡL��P�-9�:�*#J�A��U���tML.\�ZIQqP�*?)e]��P�3RX�E�gI>�UEd�*��"UB�t*ΦW,�Yu�\�!!!;��)��*(����,�fQu�&��(�G�q������w�q��T�7}�N���gU��:^����O�}O���	e�4���3"B��ք��bj��fg�M/-kes#m�e
�hIb9�m���b���]��c�f�:P�s�0#r��h����"�#�]�UkI�c��4A��G`�9�����1aT���9;P/WB��p<�1o�\������V�ӄ�H�����v:+�\+�:6���<��>s ���q5��nr�q��NR"�X+���JE#��**A�*�ۨ��G�f���_�(M����ٿ`U���a��+���#c����uR�$��:%�wz�GP��S
���{b��8��D$_t�w/Z�|���	TGx��U1_-���dk�4O�n�����4�:�z 9�8N#Bnm@���m}�q@�N j��$�!���^����p}#�UD.�ֲ/i����4"&Пx�����TsM����`{e�j,/K����7N�Oxv�-�/!Yr��Ga�NIW�pdxJ��#'���.�z-O�h�:�W�|"�����ka��x"�k�+ZA����V���V
�Կ)�X�>"���l��wB��^.,�oG~���y��� sI�x�D0��Ж�1�%�/�r��b���8{X^�*���I����8Z�v�Vw+��C���k�?������ ْ�]���է��0V㛫�c����,�ή;u��	��w����1��#���������A
��
?��V��*�jų���3V�<o�g İ�p���Z��6=��Ѷ��ٞ�v�1�򿐊ʺ/��p�f�X�8.Zv31���C?�[���Cb����0Zw}���C��&�>�#�6;�!�����T�~��h�GM�mS�ǧ8�M�����Qy�����sE�z$P��L����Bؑ/W�ɡ�6ˁΥ���7
�Mǳ��PU,��HM\��cg��DӀn'����EO	q�+�8Kn�-[nH������s�Fj�9�"z��Q�>�~>��.�Ԥ�["�2�A�'<'c���r� (���"����|�8ۼ�b��v��=�R�w�3��p�=��'�/��`����5�^�{�����W1[n2N���zp7)���(���9�W�T G �a��b�z�o��P���1eE|�b���VC�)ۅ�������Ut.��Z��	U��;���h?\p���Dp�'�4'�zw��\�*�hDmb��d)��7�$w�%7�FX�gI��:O<W%�ѯ�L<��w�_��ȡ���LMntY3D��;���D�}-G�yw���#o����l]W�Nz�{%wZͨb��9t`j�ٷ���7��NɵwA�v�'
��M�8^h�f�ܵ&KK��=5��^�S�>�ȸ����tF~��<�6�)J9c��*ۂL*�f�BA�7{�G���m+�����R�7�QꈂjBr������Ȝ�b���lh���RV�j����6r;�t�N/.�
�	��>��?wt��Q��q���	��ƵJH43k����MA��� ï��~�x�d�H��5�/o�~�K)��,%U��;���m1�:�k΋�5O��p��Uʙ7�j=7�y��ҹ���~�O���=���*��6�`sCno�\�8��LC�ji���W�Z����7�QF�7~���w��D��5�	��A0{�!�[K�9MCGup�����)��Ƀ�|j�A�Vp����nf����9���蠆t�x�e���2�j���v^�Ƴ8]�
-���#>��t_�ӒW�B����Ń���C�m�S$]�{<R1��#|}�����^]�3[\�Ņ3|[��=���.�#g�����	a��.7mp���v��6��"!{}{�J��Z���I��r��)�y�3A"��>��+���S�EЯ˄��Nǯ9߽�b�!�R�q<�Tއh�$}�����`,��2oS)g_�@%^��3�),��6A]}Qo?,�O%�09	�;�.>����qCV�v�f\�F縆�������\�Ƅw�Tl����{��AQ��'rm�4�իo����|>|ncw9g�R��G�Zs��p���Fg�4f���ro���g��r4Lq�0e(���*���c<�1 ߉�Ew�]���R�p��J�3>ަ�F5K����>��ݢy�~�/�4�t��z���L8�����cKF����V1�,Ӂ�>�;�]_n}�ܑ��g1�>/՛�M�^B����bF�>�A��Y떰R�S�k��ǵJo�)S�;TH��ef�ꍾ^���P{��(�P�شp$3A�1c�ʃꗥuH�m���n"=m{ϲcOf����1_���E��3�����_-��M�^�L�D���'��Q�{yH�F�羣޲_��u����_O�TF��$bۯCa�S�ь�k��O�B�"��"{�`[�	�Y9��.�_+��k"ߥ�E��bZ~�!5>���Y�K�(�A���~H�1�|_&G�����S5���w��5q�Xgc���"����"�z���LD�3=]�z�]A`d�nJ�H�(9X&�q�fm#�[.K�X���j�1'��[e �h�Q���kFl7�px(S0b{���@2�c޿�lჃ�x.%�U�>�K6:���Mqv\y��'7e�f��)�o����T�)dH����D��Q5;YN�N����V�5[m�h���[���{�1����4�4&*����z&v'����� ���Y��'�S����-c�P.��xu�Ix}�%G���ˣ-��I�ݞ��ұJ[�o�������.5S4�mж�[��f,x)�(����԰G��4"5�-���}�����cB3�������2'��f��ad�y'�f��̥8"��f:���;����P�n��"a�u0�u�t&0%Y���Q��f��mE�zk��],�VVIƠ�d����|:��X�X��m���O�ŌYM��iڄ;s���옹�>w�q��`04�13�|h���
���㑿����+��XU-#0$�@>�G�ȹ7ÄJ�y��Y�y�m0�����ô,������X��ѷ��X��Bj�WqN��"(���w=�"9�*Zp�#��S����WB��D�?D6z(	̤���X�k����j�36�'�]n�m�X���D_'S
5�f��)M�
A�+r���;�����-��$[��<�j�F��àr����rpQ��O0����W�g�*�*�eԩ�]�s�]$}&r��g ��J31.*�Fq�ߍ�4�G!\yJ*�g<u��`{��ڹ�I:.J���J��������5��l��w���vT$�×����ע:�s��w$�O"�Z$�CF�(�����\��b����諭�|�x]���C?�O�"�̛4Ϡxmz�xmKz�@�r���Q��^{4��Vߏ�c��"��q�c���1�6DAEW���E}7�[g�s�9;e�l�B��a����
^LX��Ė[�,Pw��2v�E�NI|jxJ��# �{׈����Y[u�v2�.��[UuU��owO�c����<yB����4n���5h��X*�R�0<��cT�[�?:@��߻7�݄��nfw����n�Q		q�R&1��|)��b�����a3��pt�S�����r����6gq�`4�/�|�o�κ/�)�ϑ�eg�Ӏ��c3��{�cp�8�̏]������Z�C��c����*B��虄3�}{�M����4_����a�n��pz�y�" �`{��h�x�˙�h;����>=EH-��b�Mw��p9Դ[�ĉ�2��=n�_�j-�w0�OYQd��.)�1��'�q~����krŬ[nH�-�Gu�Ujss��R;|�K^����
�R��a�D[ ��}6.xN�^�Z.�>9�{�ȫ�a�J��y���j�Nt�~gƷ)ɕӅ�5t�ƴ��V->��f�O��K���w�ʧ;7	UnAlaMmͮ���[W(� 5]PXbm�5Լr �둻�#�L.���L�di���R�;����6nj���|9Q�f�Oy��W���ﾪ���v^��	��w��{��&�I��{���c��~��o�p�=����_@��T7�(@wC���b����c�{⺦�'�+Q��u�9l�ܤr�5*;�쨎~�(�}�B�&���,Q�
��ww��C��m�a��1�o�d<��A�������*����{e@��tx.�>�����
DA���:%3B}7�Q�\�*�hDm}��<�P<���AS���uZ��N쿯A��{�L:4L��P'�Ȋ�w�}�t�ҡ	m���!q�ݏx�d24(��=�]}o(@��FGF�fnOX��
��zTP����WO����[s֩ϒ��ں�K�Ѿ���#R눫�z�m���) �ͬf��Xf6&����q�K+�u�/�[]��q��ut�G�Vŵ��;�b�@Qi�X6=��ߍ�c�Y8b�R��]�||��<�^/����C>W{��no�����qc����S��t�����P*�N�4QIC|`��S���ʰ�~U�M���w��E��,2/�SP���\8^{��]Y�j���W�v�L�\���Jr�&T���c�%�I�J�2īК����a/�*�a]�>��2)���&v�L�NpW6Z�᯷w+c��j�':+ܜ��n�T��vk��ݣc��3`�遑��RJN����Y�   �EϹBX�VO��3�>�Ӑxг��E��f����2�;蠆t�w�i��d�_�����l6=����W���ӌT.�ռ#'�]}9%�O��ȱ-�Fح��-����Nm�X��1��~��o����>S6�})��o�t_˧����v�N@a���%Ə<+�-1 �r������C�g�㝪�1'~	N3��3A#o�����Au����ogfH�������&�"���&s�U�gk��ϼ��7�:M�=���9`)�b�g@�;2p�3Y�;�=��"�����a}T+�ߩP�W��y�z�=<�,5N~�(��%z�s����W�p������t�1�ف�$0ycKF����_�y�N����ޘΔ��#"J��_������oh}��us~�u����EꝍG:���V'���C�C+"=Ԟ��Ef5ds{� 6č�f�h��*	"x��ŏ**}t����؊��EU�M��;3;�oڡ���:�_)�a��D8h���qk����B�����Ş���ħ���]�)-�ٚ�Q�|6�4g[;O�Z��]��Ԭ�B{�
��.��C��*ZS�ѱ�ԙiH~pc��<���M��93���#l�㮭u2n�xe<�z�N"�T%�=�q�m�5��)��J�hLQ�+�#G	F�������*�5'�eo�����j�������>�b����K�[u�b/�LW�}́ưʘ�n�D3n%�n[w�s���X6EV	�k+#������v��/��"ץ�qa?R&�`ը��ps�o����<'��y�=# �CM�8�P��N�����l7��o"��a��[,3�v�Q8���I��[�ԯy��?L�+��l�y" �Ñ��i�fю��8�T�sf>�J��C�7��:-j��U����ŷ6�z�SN�@���^��rK��A���UDe�F[03�!vO��G�zw�Vk1���Q�aL�l�
f�Xv1�;L���^�{ӑ.���}?PB}C5��6�q�7��=��}�0�Vs��u�p��7�̀�+'����3�3��8�ջ�m1ټ�{Vp��,NEIc���#kdT;^w1C:�X����P�P�|�ԋ���8Ky�>����˸͗�i�2��� �'��Ib;�Q�V���-g�m���񘱋)�]�������U���Tw����[�V`W&#�O�|A�m@.:�!�#}s|^
�M��Y��T-�A�ߗ�L�y���#Tr���9����y\�𕭺�n����+��O��H
���K�l���)wJw�%y����K��r(�l�����V�Xb�R�:F�ξ������!��p`�����S�p"��Β��"ތE��*�����W��$�r���? ������
2��� ޚ=CG|4p˯_��W>Zi����5�Y�Tw�t����^!gк���G#9H����a�R �O�1�иT8� �'�}���]��Z��~M�Y��W�����;�Qa�f��)Mz���'#�y<�����	����w�{n�/>�/�ځc�	�b�Q��|���p����5O�@�!n��F񎃥�4NDމ���g�0mz��u�	�N j��$��1����o��d�滶j�Y��n5���0�
E0q�7�[g��f�%v��o����2cW4���5�|�
�x,�?P����FN�q�nK�M���%@���O���^�y]�<�hF�L��Q�պ�O���`>T;J��41�żN֐w��{*nJ�PrX��*;)I����w�"D���.��_{հ��u��)��*�V-�}�/W-���¦`!R[�fM�.����y�=�������xw��"�s��,S��#4����pZt/g��>�jV�ԫg?h���p�+��=�1a�LәG���x���lv)�s���y��z��f�SΕ(锟��6#�y{tB��^(��w�l��|(���$�d�ݚ���z�oA�b��:u4SȲ��z����':�[��ߐ�H�P�+tV�[�(9��#gh,�Ih���=���a�:�7��VJ	��4].���}��IhgR��qn�:�̹ �+{��¢#켛�T:����)�Q	���ntH�6�g=�}��Hݴ2�	�ȗ,�h�R�|.��.����+��u��*�#O`{��n.�����t����I��>@t�\�&�I�ޭ�zz6ś��Q�����PY��Sڛܙb��̕��&H�@�^�mXq���²�h�nZ+��Z�B��Ͱƺ�ً��ø6�.卫���a¦�6
������*�CnkYd,����nT�|�G��r��b ^��:sou$S���aX���s��ٯ>V��*�"~��ޘH����H+��vt����Uv��耙��=����/�LP�?qu��)�Cx*���YJ�X��楗��-�:�i�ec���Z]+�bgJd�{X�N`�8�v�ּN�bL��7� "���q'���p����WɊW��}�ޘ&J9�*g��vf���;�f��̌�ѿm,�a���43�K��Y��ܿ�Sz��ŭ�ݨ��uҫ{/�b�+2��7��'c7z�����A͒���\W��j�+���u�ڒK�Km���Ns�0'`����qU;� ��E7������n�Ã ]`����������F��g�spv�]�+ۈ{{\r��̥���ͽ�̅�1F�4��]�� =U:��+5�3G� ��6�umr���A��J.˭Y}�F�][P��C�EG� ���f���P��e�@�Kl�)��;u�	�&���-�2��`�U�M>�j�)� f=\MѦ����n��=z��.R��6$�؈��Ժ�pTb�}3q�1��{������0k��>��GL����G�����	�;F^�ZjL�G:6�.0t��3r]` S���؁�7x"�6�Aw�sf#Ö\{M>o�U�v0�ef����h�}���+���æ\���!�n�S�O7�g]��{o� ��]y�E����
�������owP� ��V+��=��2_[��^�Md��}�)������*�	N>W���,�7ٿ�G�x�C[-�N*++��[�G�-<���%�$�Tڹv!)_r�%8^(][�����Ν�6v�1n�}6U�rQ���fVV[���
w1� �m�QQu��vR�f�E̚2��.e���T�Gٌ��5�K���&;�7-�{8-..�R]Ө�ɷݲ�s5�;�6��L�c��.�v���sJ�]���BElE=X�����r�@������27��m�J�Z�Ӥ�n�j-b��:�t�����n�̊&�q�k�P�ծ���Իȟs;�]�;�8�\� �_KM��ª�"e�~I�G�eUd*1"����
�+9R�˴�����Z�.�e�K���jg[4H�TTt��:YE$TR�.�yҥD9C��Al�$�$�t԰������ıs��L�9ܒ]�
bT%E�Z+rB*�p���B���vS������뵅�tI���t�e�U���̄�p��
s�:�DHp%N��s�嬸P�'
�V�H��M-e$���9�9#��f�M=ю�ª'3��l����)�#;�e9S��P�R�
<4�U$�!eNyEW/ ��XPU]'9z��:E�
�K,���39q+C	�R:	T�g
b-6'�
�wR�XH�
�9�C��I\ԩws����]Z���W_o?RA۹�y�-����Y�m:��+#V��gvq�(�-v33jgh����5��Lq&�S��úv���Z��_UU}\���I	���f����S�!l�HC9W��-��f��|p�✏k�wgz�U��\�O���R͍bE1�2�>7�(B���
v1[&��M��EE�kL	��Oe]�5��S�>|f���z�:�S�TY"4� �Ha�G���=!�ߖ�C�=�F�9�n�,��y�����5$S�;�8����ʅa�)=�"�2�Aځ?t� �ء<'c���dhʎW���'��Dŝu/�)���ړ��H[��l?H�6�iXO@W�r{^�@�)֭�D��D��T�wN�E�b[�p#]ON|ܤr�5*8쨎F�~g�G��3e����` ��9����^������X#�M��?7��e��rKXN~߉�;��Q�F�F���:�dDR�ѡ>�Ө�u�2�dDm�|u}
~���n}�A?p96���66!��<����ǻ�u�Dئ%@��;N��WN�o�X��̨�CʡD����Jc|���N�l6$1_s�0�E��fnO_���bTTW�zTP�����5yJ���lT)�>���=�I�9oj�~�?sJ��gQd���AY�9��9�� u/o3�Js��N��'��q�V?d�Pq�D0��&`�57\�)!�������>�Yvg�|����^�V� wܑZي��kr��L���UUW�)w��?Ozg����+߂v�E�k������w�o�_߼����?����e,j@~ҡ�(��O�O��82����#
�0�����G|����i�w��E����{k��xe�UΦ�d���{�om1$�(���5>�}l`w{��no้q��LC���g>�@z�|���7�E�'�s�,�,�����qT��h!?z��X��j,�o�)yd���&�ߕb����ޭ�'p�?��j�?

\m��1�2�;蠅�H���%���Eio�Ui��E"��qxP�Vڷ'�]���}?
b2*[������^0�ƽ��ӷ���Uڌ{ԉ�m�3l��4-������6�� N@����c�a	����ig����#l-�E����(R��Jq�~��	���p&���-׶�ԣ`͋�ֱ@���E	,q&a��_��v���Tћ�Caɿ���a�����n��	⿑w�~_�T���Ɨ���B�b��v/��J�±��y�z�=�a����b�u�O�WY Y��g`[��ce^��!��T��u��i2�%�7�,)9����Nw4��5S�H����9.�l�vD�V�S��u��b��J->lB��Өe�pj�xIz1�s����eL:�rH6�g	�FD���}�}_lG�f�J�}��߱UD;�&#�l��#�1��Ɩ��<w{U�x]83�}U�@���*�χ8�ƣQc��׸)��Z=��C�!S	��E|=S����g�v�9T1ۃ�Tz�8�N���=�D&ʫ�����Ql��p��
����%�U�z�~����E�̵�!+l��8��(O;�G~V��'X�Xn�SS�E-��M�^�Ndqy��dEF{�� !Ѣ�C��H����+�oW��{�U�R��Ca�S0�1���:gv��xC��޸�u�|����B}Med4j�~�����!x�9?Rڅ��]o��
�1���1Yr�ά���#(F��3���z���Ӻn߮��xl�E��ؓ���n/��#^wBt�Yc�EG_$l��}>��IV2DAa��&�q�>�6�X�VÍScb0\�����ۏw�"��b7Nr�e�T)��ځqa�W��\�\X
����~^`N����zdX�S����T�^q��1��R��.9��M�Чi��� {���K��G#�E�@��O�OZ+q���Øǿ�X����z����X�GC�h-4-�#5�&hR'�_<��=հ�Hԉ#sSD<q_wr���w{RҽYl|vȶ^�(:�����Fj�C�.����B9�ᒉj��z7�e����諭�ۏf^��07��Pڔ!X�Q�"����v��#!�})�o�����u�Z�wG��1ۓ��N>��#Ä�(IA���#kdT5�S�-��4dtu����J��	2�6�P5rX�W��	�x��? C�RP��uͲ�e
[��p.�S�1��\�:4�Ū�����g�K�4��ÿ��2LG{DΟ|Aؿ��d�q�����_�b��V�Uܑ'^y��n�E���@���(�=�c���4ei�@ר��(��!
hﰿ��!S��ugN\�1�w;�K�;�>��>nR9O�H�`����Q>u�B��K��cX�&�g������pDW�b����M�Y���~+�7Q��wP���O�ϭ�C��o���8��pN��3�+�u��>��<�_�_��I�]�Ga��6�1w���V?z�3*z�m{O��9쌂�ēh)Z'����>��^���;� H�N j���O}<�$}�6<k��|�'�b�1����"r:�k¿�DA
E0qk2�<.��r3�^�r\[M���L�јU�H�n��9��H�4�������Y�q��,����h	3�dH���U�����ra�F��M�
؊�A�M��fV�2�
�}y1]9cS�xS�ݮ)�d���,�	ewvt�Ώ-h��Z�3D�.ێ>��U�+�����5L�����yP1���E��ƀҿ��N�q�nK��3�*�-�S�z���Q�BD/ڬ���ϩ|6;]+��ZJ�ӟ-�!���b�'kH7��d
ʛ�{5X�f�*؏��T�A
��J�)��ʑXb���y���tG1.=�r���T)���3��6<o�_De����UM�a�����E }qRb�z�B+9�E��)���e'.�-;��l��(;�'`Ǡ�yG�a�(:�	B�
��t����W�{fR(#1��Ҭ�n� NOG�t߫q�j/yV�g�8�2���ALG�	���(B�Kbż���/�:2�D����+��]���v�@kn��>){ja�
U��"4���u�r��u�a�����O�Q����ԭ�!9���I[�.����)�z19P��Ԥ�8AŲ�	��@.6"���!�_QYi�k���ul���4y/X����&��=�V}n�q~"��8A�� ���}3dYlO�w�������>{uq� ��u�.���IY�E�eDu�b���������(R�t�S~>/�LV�}��R�h��Q���uI���Z%>pb�|%s2n⩮�<P��)�����IUאb_�����&\yJ�����\����V�n�l�Kr�c�-�G#ڌ�1k�nx�N��T;�W+h3��פ�P�ɇ����	��r���~T	��d�D�4$Ɨ=S�7���y)ۅ���g�W��Y~rb#.�پ����˖I͗�ι��:pA�_)��gD�j}7�Q��s�ݡ�1SG�ǥg��W<����e��v>SR�9
/�I�]��2�P'A�"�����WN�n������Y�F�ef�����{֠m�`�bC�>�
4Y��ܞ�8���h�z��
�d�.�{���/�_�4���ZϽ�[�7��EZ�8�~�ŵJH43k�3={Z/^L�@�YǾ���6�2z(]z���OҎ�Uz,>n�;�b���E��`߶��z�m7�9nԘ}�	�}��[�3��,��A#�������k����S�Ϲ���N΁�%K�KҧJ��O̾�����\�x��o�c���W���T�{h!c���e�DW�MCRXZLDX�ݏ$#%��7���N/���E��B\���f��Fؙ�b=`Q��z(!�y��&��;��G�en�X����:��S4�����mS���{��`�rK��HS�R�Dl-�T���v<�6&*�_\U�fj�<�"�)�Y�	���j�4VQ��.������ڈ����ҹ�T(g
�V��d�]f7���]EE7�]IXZB��Q�:�	'b���}��9c��w �A�r� OuS�#.��Y�s�Z�p����磌�z/@���߼��T3�(.�m�)�e?4-�����6��v�	�����1!U5���
�hJ��N�Z;k�l��]LT�'S����N�_Ϫ�L�������Y�5�s�@�gb���V��>=Y5�;]�^}�M�#a��,MԟT�mu�L)�W��i�7aM���08q>�{�	0�+��F��WB����7���Ӌ0Ӳ+�do��
��Frg�ҿ=UcZ�3j��m|6`G���hI�-�x��cݎ��^��ӹ�t�w=�h���,%���]�`?PbLu�`AA@�Q�z�cQf#b�����Z�v�36�J�T%1�m���W������<<\(�H�3tOA����r�.j�	�C���/�����G����^'X�_��C��IZ'�5�SX�׋1�y{^�	Yy�8cO(x�5Sȧ�[�x��~�b����K�_�ס��ҩ�̻� ��9���W�8��q�>��:��L�9_1>�����w���;f��[X^�!��J!��<}7g�l��Л�;�>Yꎻ�u؞��u��!����|� �K�.k�[�[�v;]���q��B�g&闒�"�er��\2v�{ΦѬ�K��įM�GKn��szH�u���x�x��8�8�i_Iɖ���CY������W��\�н��B?�~�����q�d`R=^٩��9�]��o!�j���*���ڵo�P�h#���F�	���6��}��rJ���#,H�ڃH�[AYNZ��#o}6�"���U�Ϟ�C
�#eJ��4�OU�x���r�_�j#��,S����`�՜*�^,��9�6�F1+L_z�!Y�㣉p�D�<�m�ǔ�20��ޜ�x7Լiz�vH�;�V�8y�}b��r~H[R�>��B79S������	�͆�XC��M��'ވ�B��]���FY��H���2J���AdE�:�ѝt٬VCE�j����W��o�B�7��c���X��<h��|k�(Gq��6��~��m��ߗE�cޅ��;|�Zf٢���B�`8$�wzO�|A�m�_L��Q�,tL3��-ӭcq���hO���?���f4�@�}]
�[��_r�ذ8�~� A@�u@;�dA,��eϭ���?B���guP�a�����R7S����X+�єO��T(Wx{2���a~�$$+)\��=��Ļ��F��2�d�b��6F�&��q�)�B�t����S��o0��ͣE$���v|���e"f�T���{*S�Iڏy��m<�{z0@7i5C1ko	�ҳ.�Gy-�X�9�{��uʜ^�nJ�/S��v��k�U_}_R����(?�?}���} ����[����v}5�p�E�u0�_H�L���u���T|�Ee���\ �H�^ ΉP0�U�WT�?�uDuyz�FQ��F;��`���'wU���϶\����ddv$���"�h�#Ssl��V�^#=8���q�בÉ1j=����c(��9u���;5�aX���'7�[g�s�9fQ���D��Gy5خ��z7i�>��C�zXf�~���ҿ��vˋ꜒���T	dW1X|Q/_�e?Ssr�?f����[u�\�=9�[,C�~�o'�H9�Y���ٸ3�7���H��>���u@f&<$��H�bƪ�9�����1N;>�Aüjų��z�`�t��y��x�C,�gj�x�ld�����S�!�w��"��tX,S���V��q׽��R�:�ibv�㱸e�'E�O�[�!lw�B���ުl����(�T6���{3Ϸ�]^}�_Ц����ӜDe̳�D�P��#(L�����lP�C���6/��pmV֍)ҶD��g2L����0���	�
���ԗY�rV�t��.�ι���5e
��e/���r���$W��F�j�#����ҭԻsP��	] �ٮ�A��m3RIc�$��m��B�f8��՗V\���7����8���'�}�چ�7�)��ȟٳl��r�h�q��E����OYQ`�g�İ�#��p��������k_�����=�b��RE�؝���b�g��	��=Ȣ��Ё?pՍ��]�'��C�Ph�ښ☥^�����frv���=�Vv;������uP��i��L'C3(��=��Tc���B��m�Ƭ��>���9t���H�d�R�}})ˡw,]��Y���l��������⇪b7���ud<S�9�>|rPɠ�ģ}����oG�}�q�KF�=��߫ʀ?uyQ[I�S�:��\�*�hDo���ĩ�����*��<�f5g�������H��-����aWM,F��A�:�5��8�Y>�U���Gog�}N����:�ߠ~�c���ؐ�s�1@#��MI��Pd%EE�*�5�>R"���btF;�>�O�qϫ��qx.�
/{]�U��p��5*H;�X��3��L�	�N���K�c�:�f�S�f���L9�@�Ϊ�X|��v|���`c�@Qa5�O�xH�B�e׍´�1���Ϭ
5��8��w����/e��g`�Տ�:	��CGB�ڄ^U��B��y�Ղ�4��R��h2���N�:�a5!5�V��_%��P�tQ޶��]b��m��O�R� #-o/�X�C�݁7�ݽGcu�2�k�5��0ZpU�|Wu�Y|�ʂ��4�k�\��7A˒dhVr��B��JM�NT��/x=�l���D��lSN������QpX)qd��G���8�n; "L�ښ�ytv�����ԻI�e[j̥v�_r�թ�bo7��s)��+��˟n۝)Vo�Z�ʏ��#gX���[���:f��h��sSQ1��U���`!�D��J��o�E�]��cYeAib(��(&Q����@�.�(�e5B��Ӕ�gsw�Н ����e�Εƭ۠�Z��)tjsR�ltgr[�Ѻƞ��)2^�vE��wӪ��k�z�n��SE
Ê�Չݽ�Q�!R`�r���B�p��e��^��c�ȡ��8��{Z�;���F1���K`��W�Ͳ���ڬ.>ղ��]��W:���͎��[!���q�Mӏ3YL�b�F_�on�"OI��QmGA%�=���S{oC�����Uv�&H�E���i�f������o�3�_PM�VSv�;�qV42��&�k�ڒS9͔��]�0WT�ƐÅuu1��8�U�軖��6���Y�^����ٜr�4���U�䯫h�hؼ�8BFua�n�1.�M�t�K�{g^4+�a'��U�9n�w9Pf<ߊ��m8����/��~(����	�Ҥ���;ruw>]��2&j�[���Sx���r�m�������!�����g�A��6�
}��$TC����!}��or.;�:F�8�jBu^�G�Wv):�Ix%��R'��s07���͖���n�%�%�TBо�u�c��jp�O7��&��H��o�Ex�����(�W83C_�ux�^>1a��w��L���b4���;W�9WZ�+���СoA�\�F��Í�H�8�Rj�ǳ�Ou\��G����4�D�p���i�CQ�St�>�qbƹ9ʻ�L,�oF%��=�t뢀fݦu3�:h�(�3�����U��pǼ��E�Tᗵ���-f�*�;N�����-�f$��i|{���v�>F��m��A�b���ެ\�-n���,�n��΄5?���I*��J��Bӊ��@�w3+/sJP�#rv��Hm�{�yOr$�����E�jU���
��X���C-y����ha�d�"tԍdk���r�I�j��'�MΫlGzm7х�~�FV�Oq���R\��Yx�2��h������=i���]b� ����b �t�/���u�"I���6ZN���7,�Օ������f�a1ё��Z�Q��n����-�j�����9۬�e��J��v��rR��aR9�g7c�*n������g���
�dt�����#:Q18�BAfAT�%S r���-*첢�8RY���d��=y12����aL��94��e®�"J �V�cղ�T�C�.��h�)T$�0��3
.2�9����t&\C�HS+0r\�H�J�$�VQDEˡ���(��"����(��tV�L�Μ��rȢ�H���p� .Bq&QLC$�
��%G�r��rI�$\(L�N8�kO%�8S��('\��p��0�
�U3�sK��Fp�w-9q:L5z�5i�76+�r�.:Ewʻv�8E	34�5B�M<��;�$&E�p��i�z�'B!;��6��*���+������Eg��
� �Np'��y�w5�!&	�LL�H�E�p���E*�I�V2�VUw��e��C)����IRR�e�Mj��4�΄^ؔV<R��q]��H��۠�z��,[Y"�������}��tgJZR�&���g�xefвdx�8
F�ޯ�� ��x6����S��t�8�Yp���g;"�]�b�O�gzr��,a�2͌>&CG�O��d6��m,z��C����c2.��x��է5 ܂��gn�S��$��880.��y~ݯ1�6�?v{UI�B���V�BᕛpoR≔[<�2���ڧ���0�?��ƕy���2~������ǫ�ϒͷS��<�[F���"�[�ς��S����:-t���~;>==
(�� .�8s�!���'���=����g"�ծ�(aq���N3���H�|��lO�{�2h�\�<kQ�/`N�	�����[SP��d�w�]�b�ћ�l93^��)���kr�\#|�e�(��c�ɉ���
c�*���yxuؾ.T�����`=���:�xQG;��J#q�*�z�;u�������&#h��t#��Z3��һ�TL�Y`�Ղ�ϴj����3��P��v�����Jo��=���	��=��B\z�Yw��㟕�Z���d�.7����Ӊ�c]��
�ѨϮ���-榚��h�=�G]o'��nL�̊@��LT�Ҭr��k�؀w��U�6��xLӼY�k�82αA�{F�sd�C�U�/$��
��s��;/�j�!3��n�>���/��?X^��8�?��E_��=~V�*��ؠ�ۛP��H��`�1j
9%������
`���*�i[�C���#�?+qx�f-��p��!xEv�k���u�Ոǹ�-��ZoeՓ�(Ջ��|[������7��S'�	�R�u�bf�'�����&�n��fJ�xz3��5�]��dς�T���YY�W�ݦ�5�Ց�D�*�T�&��G�]<pǟ��XIW��f��dk��ɑ�H�	l������.	K��\l�V�ʭ� ��w҇�l�͌r*���S�>���9%^H�,9C�.7${rڻjؕ^/8��[
/�)��?��x�X��
�r��9%��O���Ѣ��`��{��$31Ҫ#ОF7�a��S�z%�g��2��۱�;L�ϧ��)�1R�ä��}r��&��&�ʽO�4O���*D}�(C���a�Rc��8Mϸж}XE=��dr������h��c���'�f�!�+b�ʰ���V�0�:�Y�M����vh�-
 �Ș�Nc�Eb�u���I,�^n���wv��w�z_/��֋� B:�j)j�.Q[|��A(l���,�+��|���.��n�<r!��%bX��sǷݪ��˶̍�|�R�R���V�z���{7�Qm���[�E+�	+2^>�1BS~��ZMo���~Z�����\�J%���=Ƅ�#���e`W��ָ�~�[����b��H�ƠSݧ�b���5�҅c�فL�1ޓ�@��ڀ\u}2r8�������&2�w��i�m��(�^"�'j���U�[��@#����3�@���甽g�Y�^`�u�=�wEʍ�J���*�O�vC�zp|ܤr2��CV'�Q�J�w�H]��~�xw�����X�������BA�={u��֠t_�vC���D^�N�>j�{ƅ=�5���7K�N.��L���gD��U�=�l����P,r�F�y�ܣկk�9;����������H�,��5&PR*���&�3���l5��q�����ȯC�{�����`>���9E}F)xNC��Xf��
ES��~��zE[u=h�[~�����w�g��c��6=��5�,3a�Pb�i_�_K����P3*�*+�k�s�`��E�߈�xe~PW�E�o}����j,.t���k�[ϓ��Ր+쩴|(�����M�*�������b��#$K/rW	��F����һ7{۠���]N�jL!1���;Z����Pɴ���^v�䬦����7pr|TZz���	8�%�E��Y̛Gl�̗8M�<̧�np ��z��;}0��96ΧQA\�}���wm�Zy��`��$�`�H�b��[���tY�)���8w�X�e�P���i�G�<���`�yE���rN���X>�����W�F�:���8J�����L��^>�cݎ�\?���������;�B�0�9�Rf��D�(g+�V���l�FT�����ӻI#��Ƣ����ۧ4ޑ�2���v$PS�p�!^bL�e�����������oZ%x�.�wM��÷�sj�S�n��b�W�w0�Mղ�h���*��u��PQ��Y��rE�u�mga��B�Ԥ�8AŲ�Uw���^�ߢ�+���&.�'�on���z��^���ړ��T�n��g�4�u]0s}��Z��8'�6��������^�]j2	n��u=-��ٌf�ϫ�`��}�>\�'=/���ʈwӐ
��@�8t�,O#@O	<\l��ӣ��!�ҝ�����5D<,����<��1�׊y�����F��Q
aP
DA�:%�@O���>�a�]?+֍{؏@�ۻ�����`�'�خ�j�*�y���Y�`���j+|L0va��_U�o�s��`&�?��B0z
�DZ%eYYy{��H_#gys�a��pu��r�wPȔ��.�t��Ԙ��6���r�-���#YЧ�!D�f+�hѨ��;\�h��+���77���걱����?ņ~���$w�5���9
:�0��;��P�|�J{k�*�*�|�p;ѻk��V�8���u��V!W��ѱ�[��}fh��l������Nx�o�ƽ�y���|2TT��&r�}���p����EX^��~��R�������c�5{��Z��o�b�A��J���.(�W��U�������඘�x��j�!R�Q��o�^\����6<o��D�@��ѡ>�}|0w��5���)��E�0�Wג{���1�-�U���j���������2��>&Xr=�f��U��l�=�.3�PEf��=p��jٖ4�Fa���W ����r=�������s4�G�y�X����`�ޯg��5�y��W�ԑ���[(�~�T22�V�#������}?.�m^�Ms$�=;�T�����^��-���L�K��g�f�O�h[{]�i�<��^7�5@��x��p9���@c��AB\n�����^�Ek����Y����BF>m�¬�uy�^ʷ��/Z*��d�hqՓ-L�6�%��$gU���r��]i�|��N���Y������xK��Ƙ�w:�R�J�:�U�zI��Ꮜ-e��.�� Ϯ���\!���L�ݾ{P�Lv39ۈ��w���P�']���,���g�2�$ܟÿ�� ���'�}�A� _�z������3ʚ3X�J����ځ��������zKv�f��9aM�:v	t�B�&!�]T+�T�\,����,j�K������sQo��=jU�V��s1����ml��=~@�4$Ɩ�?(�+�p���#����]Wr̞����@�!N����W׹�)��G��u�1�:`A�z�zk����e�7���4��(J�u���sд�w0�X�V'���!c*���͚Q�3���y�'p-Ws*�3�i�c�	�1"ǥE>��+�BC��q���J*��X�%1
7���7a��wSV��5��^��*��:P�!VԾ�m~�g��h�}�������A~ԽJb��X?9ߢ�x��W��48'���{U2g�^T�ߩ`�\p~��oϥv���}��U~@���٧�ۮ�q�}:!E�ߩ��U�7�c�248�3�H�	l������l�J��"�����g�c�x��	J�`[,ER;���A����>���IW�KG�_=�W��2��|AؽB�0�%� �B�%U��}��c�w9q��'b|����e̤{I��T�{�`�׽`Ef6�m�!���Z�g�g`ʜ���ӡ0;��9b��\�$��^dYH�Z��q.�����֊��&���I��f�ß-q��9�u�����3ڇ���#?}fo�,/V��-=,Cӟr�e�z�[�v�\X{�迺�$��~�f39En�]��<���FJ���"����1�:Ttq�.-L�>ϛv1ˤȹTW���Z�Z�c�<}��v����"v�ף�F|$����w�z�!����v��#!�u� fJ��P��oX�������OW��}�`V�H��E}%z�� ���*���b)��2��dJU|��};r֚cʲ9�����z�����=��'b�!�BhO�w�ey\lA畆o>�l=���+�%.�:|f,YM���B����b$���������q�zKW\�����[�٥�6-�6����<��ZF`Iځc��U�[���(����EV�:+�_��ʥ���u��{�P{pÂQޮ�Ѷ=��<.���SӍ�G#9H��OC�Δ]��`���ڪ�y��@�~���>�|ʽ��{}��ty7A!��_�u{=��gڹ�~�Z].]�9���ǔ�F����B���)Ap,d�o�{n�/�n�徺�Opp�g}I�ߎ&;�u��/�Z��8W>�·p?��#�ξÓI�@��j�ld�6��)D��Ԕ1��PƁ��>����zZ�gs�h��Ԝ��S��K]��y�/,���p�W�5��N����=��g0��s�/���2�Nb�	��4f���x��T���Y��z�/��-�{�dkM,)Z$�L�ͳ������ٱ����܏.�[��=�k�C@�nC\��P^����0��+Ɠ�J򠄛��=��쬂Oݻ��Y�^����#���V��l���6�U�nN�q}S�]����}�gq��d����'�����A�"����^�WF9ژ�\�?��c��x�� �M�����=h�����}'Ϧ�Ή��xIQ��"�ōu�����b]��R&3�ųg��Q�O��Q�>�����ɖ1�mn��3g ��s�_|Ȥ�*Cb�z�B+9�E��N^��F-�E�#��n��K^8���8-:�}^���2���3@��@Il	!}�z$!�c�c�p�zb\��"���=�O���5�7
�mہg�s�Fd�9���A�`D��4�6"#y����
b�G�{����u�H�c:�5ޛe�χ;����f����\�Z����$F�q�Y��.!��Т�����B\B�@����ܱkے.�Γ�S��L�H|����� �ul���zh�2��\�N�^�`��[Os��c$6��{<3�������5���'<�/;$�m���ܧ�ҳ���lP(���l��]��*�VZ�{�p�vS�=�n,��b���EX�!�(�e��z���2A 'f��܀'���rE�ϫꪵW����C7�=�@��`G���;
��[/)W�(�%����&�:�U�ݎ�u�͈�U�/ѓ
�ޡƾ�/ţ���"G	�
�t� �����W�E��%�W[=�4Y�������RNы��ުQk�Q��+ʄ?p��������/s�����{)J�y������r���q�_W����Q
���
�R"��D�O�i�wgB��f��׆f�IOU��R=�B��c�H�$k�/�Q��L*�g��P�Y�v�5���@������*�Q�}��J�z���l��!�}F=*ta��ʴy' U���ʟ��t��z�J����l��W��j�p����EX^��~�ŵJH7*g�(�"�����z/{zft�i~5�c�0l`�2�����+�U���������3���g�G�����B���c��`�f���2�u&G�!��O�__�`7�so-d׌��w�j6�������k���/�g>����a��2�����G�xM@~���7G�{?pʞC+��%)��˩[�r�38o\�����3gk�n�c0��s$���%������KJܰM��{�I��:�m���;{m�ht��&����P1����ӜlY��V��l�1N��$7��[���(գԇP��k��<-��|�kG�U��9ݿ�=٘����T�E��9MCGn�
j�f	���_�r4,�3�.7��n\�ZY޻>���b1ѕlOz,!`_SF�f�l��3L��>�p�6��F}=����7f|˩y��<|�9�*�s����LE�	]QV��m�B�t�)�e>�߫`lw��`�X���b;��ƺ�}?P' H��~�
�sn�Gp�6��-u1X\k)g����e�8��Q��o���7���.��4P=���=%"�����ɨ�󭋩��㟡��85��JkxF�Ze��M�=��>'#�M�Ӱ`K!W��Ƥ�<����e�Qf��?m�͢|b�핍���7��I��5*�/����s1�6p����@�	@�0�ޙ�艔��w�1�ƜFx�SU�p�����?�.��e�߂=��@u�1��ˎN��01:��<*�;�Ɖ�p��;�0�y*�<��|ʫ��Au�6��.�g�d{�?
����z�p$1�0l/����}t����;�G?*q|�c1m�C� EH���c��؋܎�>��1q�َ?>��/�8x˥�97�VW4Yd���-k]�n�zA��ז�3i1�~�5/m¬$�-�ƃ��#�ņ��)<=I���Rq�V�"Ղ-}K/�&vV�)�<.�%�v:��2k��[�A}�@8oP-:!�q���4��n���,��vM=˚;q9���tzeL��2n�ǒ�����$�9]K�� 86����b
��5բ����Y�6�m�f�J�]X�秴@�c+��'Gf�Y�0���[dݐ�:�:wtNs��y���0D����c^*[��i��P����]P��!��f�cɮ�f�Z0JA=��ֲ��utES��,�׀�l�嵏� S��q.�3�9B��n�7�����Y�_h,���3d�N��T�AV�Bͫl\,�����嵐�u�=z�fh��](��CM�z6�bV�����\��i�n����(*�T��]!���]M�P�&ӿ��t�Yէ��q�3f�}��B0��"}�ʽո�
�6�)*vp��qS�iu��7ԁ�V/W(�4�g���e1����ݟ������8�k�,������kAN�����WL��w���q���.p�'^��-.xce�^�H�۫�|��j���q�:7��^3e�1��;�2���%�w#����[��m���s�����3��z�=t�Iu�Q���fQ��A�|�;�b݁�'"37w/)q�2r�t���"�Gk����K�O:�r]9�6t�N��,.{j#\�a�Hnp�q�-�ز��,�u�#�[b�e����,�v]�1|��L@�.f����4#�1B3kWoc���(S�y0��4hN��A#�m��99O����7b2�F[WN�HumC�q��7I
�6��BN�y)K��-��d:� w$c���-�@��p���V���`�ghɉ���`��@a���@5�{6��b���[y[�:m�J1h��p���8�� &C��m`�#b�i���]��*�lMq^z���x��y��ufg;��� ����R^�n�k8��W��ŷ���
=R��ư����x}3�ދ��t!j��5xjŤ��ԫT�nm��U+��p;�-Z�Z�R���@m�[e���\��2-g�JY]R�l3t���qۡr�0�\�TB�u1�����w�2��S6
Wy�{5te0!tNL�U+w��u�[]H����/1Vef�:	�ۢv3ԧ�E�;,\l=����0��1���^���l�̙��[�[Y��c�X�{���\��Y~�"_e�L���q3#�
�����}����hkI����os�o.�-Y�29��̋�9���kVImr�g�:pط�خBBv�2�i���Vgi�Qs���r�IE�3�q����`%�'�v5�����?`�|E0p@���HP&�
Ps�j���i�δ׭&�IڭȦ99��MD�)�ejI��]ȳ,�t�Q��.D��vҫ���K��g���9=��y�T'�^�>q�S��P�)$��Q4��HՊlI�v'B��I:e"��8��L���� ��;����
e	4DH�Ty��r�R�y���H���J�'94�!3&�99�Ԥ�W�pK�v]���v�NU$�d�$���{��t
��Q�JbO'��i��yǫN����듪�T�s��L�8�.P�ZlNP$�*�d�N&A�8\Ҩ���SbIǓù<��;Ϟr��'ɹ.�r+��z�kH�B�{�I;���:���q+VQ��==N$�[�r�{��#"���%z:�\y	�� ||�b����f�t�ܿn!7ϷGhޭFp�)�d�O��`���E�ŀ�����7R�t�3����i�)nv|�l��T�	h�"ɔ���U_AuGUv��9�RG�g	�oMa�`m
&CLHѓ�Bn��:�c��}�_H�b��{�K޻�yϽ�:e���
�yf�k��S1�}͎5�VȢpx)������VO��z��N��ǪўڼIf�����p"ץ�Qa�Ra5^�~��w�����8�W��c����'��E&6M���?L8+�|޺���p?�K�`e�lc�P�A������nJ��V��V#��=���O���T�w�a��ꖍ���=89M���o wjŀ�+�2�����y�{o F�<�����}>�C�z>���#�K���_�q�}2᳊f�X۱����t����\o�p�XF1;^�C}9��G�A��P[Vԡ��Q�"��Tb��ۆ�>���<��Y����1�>4-����=8��}�`h��O����_]��EC�_?t�&-��;���=��/9L1��|i)�h��6z���|j����A�H`�ƀ��w~	.j�/���J��Aa�?|�mo�=����S�@����\�
��`S2LD�Y�(`�Cֻ��띍��>7�	��wg}��`�@������k���.<L�+�� i���c���
d�����[����Ť>�9~��ƺ޵�K���*��ֻe�~$ޤ����J[��A2�^���T������Q�0�Ie�''m��j�,Fw�ﾬu��kX#�P��h��
�cKH�Iځx��e���b��F���j����y�������R:T;�:6ǹXǅ������7*�����E��]a�%��/`(>�>�J.�=�������A	� �.z�2��!��m@��݄Mas}2��?f*��{�/�k\Fwz�6t�f�GAP�g��t�MV����D6^�Q�k|*�a��!z3/o���c�Π0�i��tc�o䪌R�9
�H�(�I7�
EV��4&����������1%{��ə�W�U�	��_��ې�s�1��9�Ma�W�Ȉ>
EN�=�<�Ǽ�LyD��Ts�����~�l�^���A�+�+'l����.g�՝��0EcQ�,Fw�o�~����u�A�A$vM�#�Ldys���,CC�[��� ��7�q�ܸ�̊Υ��\����?TܗM�@��xIQ���/V�y�u1N�O���W�1u��e�j���Թ�Ը����fwV�<o�9G!��	!���_�E}����a�e͋=y���ܞq�"�l!̫�}�P9��ΡEN��[��Nh�p�`����VCҥ`���CK��a�������:�*CS�n����JhJʼ��k-��^�'K�n�R�8�z����v��qTwr��]*������Fs��jg^D�M�^Z�MdG����֗�Ӏ�������{����d@xL6(�33N:��9NWwEݜ��=�$.����򿒙L�����#���p,8��s*Q���PF#ƞ��D���N��_�,{��#VĉZ1[&��M�l�w-���;z�9��A"4�ٞ�/��ɑ��V�1��x.b=��=zC��rŬ[nH����S��br�>�'�{ϟuT1��f3�ǯܲ"n#s˸��Ɛ_����L�b����ul��R�@Qc�z�rt���{����r���}���=�#|����H�~�8A��K�@��~ �5�6��^]j2Kw������95���oY�ns�X�Y�j�[�TGZ��R�,p�C�Ԙ��S�-m��q>���؝��ѩ>�y��V��9�>ī��U]�b��|�D
A��ˊ�lvk$gҢ�c����s�������C4{)��7�$w�����r_`�
�h����dN���_t%����ZA���.�w�~J�*�ߠ:<�`�bCϬ�|��?�,Ě�T��OKbv"|6=����/�oh˿Re�E�����)��TZ����~�Y�ۡn,�
}|�J���e��vl=3k�2JY�FƠ�b�R�6�2����{F+���٨��~py���beZ7��"�9��>��H:�Q�.� �=������L��u^�J(	��l����8�[�7��E/K���w������C���o��b�I��O9����CB�R�ïW��:��!�����y�Y���#�o��d׸MKj�N���ݻVS���@�Ie��g����(�� �=�.MO�__�c���a��1/��Az'��Z��<�T�8��U���W�X]>�ȫ2����e�#���� �toE�"�V�G�1���p���`t����4y�W5n3>��8�`?�f�$y�s�^H���~��1��1�3��ފVu$lt�2��S4���.j�\t������*!.��1���p�ߟ����6b2+�N�6vxCմ`:�L���6x3l��ж��Ð�5����Q;�t��9���,�o� XA��AB\l�}���Ek����I]��XȾ�+w��y&�ߎy񠙰���p&�P=P'���`���ښ��_���2LsL� �����]�>�c��3�FÓ�9��ω��
l��`_�t�@@=��3Ȋ5�0x���:��k�/]�9�vݪ��zu[�L�d��>��؃�mu�'%»\4Ҥ�[�m�Z�[N#X��:�L�{~bV[�"�%��z�Y�@�9q�
xڵ}�viEB��
Q�ڑP�!˳�K�sㆲ�R+o�f�ԭh��J�|�]@S+����Ǩ��EG9�y�����<�,5�u������&#}�
�)y.8\� r71��+�b(���<}���Ӂ�!N������smVT(���&;�!�~��+��mp!���'��ꝍ���z�������!c*�ϛ6k�7���܊����w������$H�3�	�1>
TT�+z�t7�B8�~V��'X�lQ�cI�w0w�� fo�یd渋�zT�CtN3�6e�'CLh�ѓwM��>���ޯ�'%��+�ֵ>�.���q��Q��!�֕LW�}͎5�U��d��R*��@�YY��n��N�v
�ޙ�S�y��o�ke0E�K��~�!59}����248�3�#ҽ޾R��'k^T��2�8w��W�j
ټ���v0��61Ȩv�_���Ox�=F��+��M�~w�|0k
���Pi��ý[/�ꖍ���=89M���m�(�ӕ����s�$ϰ���pۨc�9'p��'��\�fEKf,o��
�:�tq.=^I�> ��+��2�9�s��Ԟ��BM%ߓq�?N��d�|�T�Im��[x�ޛM��)�V�Ę�k�e#,A(������G�S�+��_׉K���k6�Na���{.�]������;awHF��WSGpf&��YӰ��W>��qr/-�y�T�'�M�D�{;�8z����v�����]�ȕuz>�O����"����z�!ȉ�8�$3�}�z��{�{<�k��o>�Bٶ�XY��y'�f��1>�Pg�u�A}���^����G�彎WG��ƾ�s�+��`	VCE��dtPQ��f����5��?0C��Up���Yk�}�شEQ~��w_�Z����/��}�)�X�
�=���b;���]eb9��b�.�,��c�n=S!B��k��~��>R�3N���Ъ��^Q����oc��K4�$� ��3���`@���@;�.���T-�.����SӀ7)�ˮ�U{Â}s�{"dg����8��U|�@�~����� ��{u�����ɻ�Z}K,�L^'�7C�Զz�o����Q��wP��΄pAT�D� ��%������}{��o���Cތ�ƫ�k��9�����摎Rc��2a-���d�3�{(�u���)�\�6b��*��{�LWm�>7�z�'�Q���ޠ�6��W>���?t��{"#�B}������ֈ5�[�:��h���.���1:P���2���x�\�y28U�;� �ij8��0+��\F7�����m�cUk��i������Hɮ�J�"�l�5�7i��,5�J�����E�&��K7�t7#U$�V���S`���?}+;�I�������zl{e�j-zXf��/��o�{�֚>�5`�Q��ܤ���x�3��p�>���us�iV�G���A�ZX�o(R�[���n����}��s����5AJ+v|�m�W���
�'�+�k���U1Ї1.7+;މm�⩗�ytbQ�����k`���/O���e���dR>Cc��B<�i��0��V�����x�>�#4����qbZv3'��Ӿ2͌>&h�hIl\g���Ʉ��@���o+��4q��81����z����)�h�ơpmہ��,ʖlh; �Y�gԺ*�δ	�&�~�S��+a���*�^O�ZiUJ��f�_�����LM�\��x���q�� �&Ǧ#�x����,Zϖے.����ا����DT,WE��%D+�;䁛u%C��g� �@����b����6��r� (��c0NԚ���`�����Y��Ӵ�l6l/H�6�����O�Azy�Lo�����W��Ž�=5ީVZ�v�X�ua���R��(l�Y��,�Uw�h��@��h�7,w�W7�.|}�+��s�J�D�'Pc���s'ஓo�����k�٣� :l���3j^-N[Ż�18*������9���7�[K{��ީ�8�F�6�	;�{��k=ߔ�w*Zs��#�rڥ�����P� ��Ԙ��ٿd8��:#�y�ٷ<X�u��U����Y�r�����Uж�!h
pA�_)�3<j7+�����@�v\��g��W�B#hT���ҁ�n/������Qc�I�����8b��iw|K@�����[�3�:�z��+��m��R�6ؘ�s�1�}�YZ��G��6A{�K��t����,62	qQ_1�Q_M�Cfx�Ki�G�ʢ)��pu��C}X\B�߯yz'<X���~F������A����R�ï��~�d>��ˋ��@��������wt��׻��;�!6���^���k��=����2�Y>2,`-�}���r�fceJ�N�}��>��;_�����B�nt�8�j����W�X]>�7�Q����G�ۛ�˵�}9���||�=�v�/k�A�}K�Fa�IMBtո�{G�����2`�p*���v1���9��F#��P�ފgJGGL�-�)�e>�P��Qq�(vy95��uT����,��m��}��0���2W3]��!V�}�8��<���l�8pUz�*8�����*�V�;����}�,�k�ȫ�I��R��̾�)\[ݤ7YX.=��F�X�dŷ��]}��Z9o��Uk���彲����E����dY��������D������o�mp�cʢ���"��v��S���+aL�#��Mꢗ�·��pZ��6}?��N@���,T�j�����=���7]?��J�	�
��^���m��/�s�~�	��Ϧ�O�]@���}�E	(q�5�=OT�����z����}��;�V���X��&�N{��ω��Q7&'�`���HUDOq�y#��� lQ�.�?GWyƜM]�eJ�P�JW�����^j�*?��� 1��@ն(~?���kެ��k��86��!A���m���6+�����<Ӂ�!N�~)_W״)M�(��~���F��E�ӻ<�^�c��`A�\C����p��{�P���m��2��<���ݧt'����y'v_��<T_�p'����zH�r�����DuP�m�؎4���93�����NN�l���7�A�ca�?��!�7=$W�h�F��*���0�zn���]lv?*�;�(�욫b.���Y�^?oz�*�u.17^�"�����Ql�M�\6�����b} 1��=Ե����U�H�ەy�}y.Q����7�|6�q�����fC޹`Ă�����ds]wZ5$��샶����W���%Yѹ�YU����7/-|Z��uӳ,��i��2�s�E���u5Z�Xd�i�;k"W(�\2v�,�}��Q�o��5Y?V�;f�K`���P��!�j��7G�dk�6O�[��r�o�Ǽ�z^�#�S'4��Ӻr��Κ���a����W��T;���A�1y�j����O�*���=CUЇ���$���Cs�w���<�*i{�w,�yr��^] ��Ez#��m��x���ڳב�K�2��+���7��o�Yw1�P�cDz챏�d���W��Wgq��a}�xPC�c+i]�C� lE��?Aj�D$�3���R�ϸ��4�]gs���*�����N�dd��}�*l�ōYΕ�i�������|�?q�zvP;"iyǯ�ulG�}���I�յ\��Y]�n���-[s'�Z���W������lj��=�k���jn��+�w�s�x����������u�4z�qu��!�f�!� �D��@ހ����~�n�y�_�����|��TĶ�td�I��.�Mؒ��E<�S:t�ҙLV��n�[TR�D��q��r�޼q�r}�tj���D�6(�iU��J��W���IQ>;+�DDG&��u7.�M�L��}�"�]ڹ�ɫD��I���»gp� �,-o�!*��@����v����`Q�V���L�괤�.�=�{K�UJѨ��GuG]����w�躥�`&�Ԡs��P�X���j��V�f�⭷������w�vh�4� ��<�,���f��hM������7:���Q#h!���|���}�T��[%��;J��'&o
&�ظ�7���ƻ�m\��E=s�m^k�/a=���:��S��a�Wl��{����e�Mѝ|0��&N�,땜]����Tu�楚���B��M��
�Rl]��� �T!�2����/(�M:s(�V�%h.�QX>�c���φ�'��-ڋ��{����p��7,�39�ft;��y�9(m\�-�*Q(�.�Z�3E�樍��_*B�u:Gu�8Q�Ԗx������	:BXձ\��+ws9WC���촮]�F����L�nS��_�[�2��5�O<�;���Y��JtKk��="@���ֈ���XyG���6�������wm�T:ľ_)c���5�h��S�tx�Xo/srJp��Q������r�a�J�>y��.�]��jW)K���p8`��KX�Yy>T�*�[z����5�v^�w��▾�w�M\5��*��aFeCp��Po��Ӭ{��X@�ʺV!)36������R��nk�~���J�NU1^+��P��@ܧ��"� ��'FR�ڟJ���YX[5�l<%#�=9(H�����N��Y�iԠ� $�R�DeMJ)�D��Tճ��g�ԓT���f��Dn���Z�)f�b����ҷdKW+
���U,X�j��+,��a,��ٲ��.��bS�#�li�ˣ���EP���]��]k޾D�m"�ԥ�W�&�����%h�۟L��Æ�nwb��k-a���-"�H�A���gu=�y��J٫^]����d��Q�p��v={�7i[օ�Lm&7����ڛ��|:LS��o��C^��d��#I�.����C��:t�]�k��l�:����i"�ʩu%:�j�˕!*qf�tt��*���oi���ʬ
���t�:M�lj�Z�}ژ����UX}&M%T���]�l�i��b�5P�](	�s��jiЊ�
Khv�	q%R�����b\��;�eޯ�t��Q�)r`�v3����ؼ;T� ����J������
�V����hȷ�>�p$�vKJt�:ⶐ68���7s7�#fX��j�*S�^e����eXE=�݆�=j���;�Ã��囨��@�}n�ťɼ��ܝ4��\�t�_�^
�Ů]%S}�st�����:��(�����y;�q�E�j�
��r�l3���N�)R+T���2t��N������zP\)&�q2P<2����8Vh����f�43�i	\���'^eN�,��Q��y�y��Ey���Q(�,а�aE*Й�����׽a�^�G�Ea$�$Aih��^��LȠ.D�e=NU\r���0�*(��y;�r�%�.\�pCϝ��'�κ9�*p�\�K y����Q���]/D:g�!
����Ӛ�Xgtq�� �r�a��tnG�6gHy��5bJ�'�U9R*3���*��h��ȵ�+��uݱ:�r����2�+���EQeUe�fkZ)�#JY&E&G"�%�9-���i'*�E��"���\�E2++e��!+0�'iU<��J"�
����B(����,'�L��Dz'"5���\��UW�E����h�RH �m�o.���r���3((�IKh����5���_ِ��eT,f�B����,��	#�\n��&]��%fK�Z�w�9�g}�S���%c��b��4(?1�?���|�c=�6(��z�b��</3�գޛ�B�C������
3��d��������r#�gr�3�D��x�+�HWܣ�#�x_V�*���SD:��[�s�B{5v�D�T�6{R���{���9�H^��O&�-{uG
�r�1��65�Ƴ�*��ݫ�=��X�Ж ��'j7�US����1:o�h��������i�U�����Ŭ=�βY�\�:*�^�u[�r����P�u�e�ڂ���*Nup����癡�	n��d.*�_O&��r�G�����;��.��{�YT�0��~�=b%�;&VtM�����4����w0�X�/�$��i݃��7�]�29�Z�jW$Z�FgZ���^��Cr8M�t7��i�߫�I���>��o?3��������v��U�����fx�j�w�7{��Nu��,p�1c�R��=�Rh�ld�h�[�{}��|��j�jL���n4O�q���턎B�;ښ7��D�yֵtb��}R�cd�.���<�!�݃q�{��N)�(��{�|}{��Õ�	��/D���w)'�s��D�~Ӿ"���3��woD��P�&�=%���5-�V�����ֵ���ΧWPCs~ʍ�#|FR��ǫΈ���(�����ޭ�N��į�z����O4�9�6'�ݙƷ�$nw���7�Acο�@=�v#�ڰ�Pڭw����J9lzU^����z�;��s�}�O�}Բ��2���à��/�ku�������(��������Z�����^�r=�l*�X���AW��{�K`Nw�_�t���>Δ�{�g��5����A)�F"�L�x���&'�#���z�4F!s�z=���?,^��t籺��6(��5�X����Pۊ4���M�½��e�ޘ()����k���u�-}_{|���\���ѣ���/.���$bE��t6l�Ppt�a�9���WWE�*r������g����)��ɔ:���ɬ�ޒ���}�wR�%GW�¶u�Y�KKk�f��V\	\���\���8_=���ι��(�"T�S:�ci�J0�'W
��ܧu ��:���;�X�rgK�9���^d�ga�ݸ��h�7d;'6dlbX F7!`W��^�ͤ:�����&�7�n�U�Cj����M�����X��gg��i�[�u�Wꝥ�=�l:�ԮV㿂�{&����u�l��uY�w�[՞Se
׮+���7%�|4��)i�(����أ�>��"�ojO�; �ނ�d��z���2���WZ�jFt��X�8�nj9���깻@g�2�ןH|#�[By����8���qOސ�z�QF�Tϯ�r�}U��M*�����U���%����\���A�Ss,v�D��({鰕�x������]"�ߥ���U�b�/��']���[q�q����۱��է�o�����u��~��r{V��F:c����'����J睨J�y�<}�7I�wCշUW��W..����|�'6=�#S���o�='�!k���u�� ����'b��x����q�Qc�f�o�v(�ƅ��g��=w�Iq�zV:Tk^��I/��ޮ���5A�{���\���%t3���x6iS���3W|��T+kH�0�ȍl���V�}����b;]9�yh[c�ҩ˺÷�:�B�3�EQAǫ��[W�|ew�A���X:���;C]a��7Ցq�%�ޑ�o�t��ދ���x_?�X�=0F���Ԝ��is}ï���z����y�mbSΛ��pA �5�V�\h�a3��T�9�掿q�U}��d��V��F{�˅|�!K���߱��͊��a�_οQ��{Fa��u�*N80S`���U����}K[
���x�})��g��</�O����é�Y>���<aXޑ��O��o�]�w;7Ak��y_Zt��w8���E�g�*[1ˁ�_�*��?pY���]͡o����j�������K�<�9��#+ޏy3ޤ�����w۞��eP������7#����`�;=���[ݙ�t�ZI�:�&�ؕ�����_f!B ���H?z��	ȡ�?N_��U5��C��OusY��>�{�o�Xs�FYZ=��<{r�<�o��x e���n�R�%Ř�(C1���>Ӹ��F #� C;vw���=�Ay�_�JP�hG��q��𢺑^A΄�K�n+���p�w,ѵt��7 I[B5@.ݡ{�)��K�Bk�b�#�u:��F�;�e,���wj��3��EIZ���3�e#�V����uX{�_��˥N�������
Q7r#��!c�����c��j�eu��wx������������N"�G�{z����m�j`v�|��\�VZ��^ϝ��SO*���&b7ؕo;��cc��ځo�1�p7�6����n�o��M,[��_���aU��hCs���r�}CR�
@�}�xbzAj���T_ר��w����69N�x�cy7p���К��yk��,�0Gx4�b3+�7(z�סn��0���ܷF�^�ʐ�Q�A)��ϵaT6a��؈�F�|�@:��} �v<�����v{����p+�B�V�<*�,���Բ/'���EQ7m��_gݯh{[KU�X����M�G�G�������.�}Cfʮ�8��7��=��m_�AN~��K��~S2�	���H����3r�9W$ɀ����vf�q��\�,E������I�%�����	�|����ו���RXv̝��5)�"8�N��g��3��ӨT)puv�����7#;��̡�N��`���c̳����	Y��(��>��^ԑZg����o�~�Rup��[C.=^1k�ɣ��e����cy�x�;�.�[�VU�B�ac���/������_�/�w�o�^������8�Վ2��I��Zwgs(o�����;�O��E�심���C�`���
�!���-�����%����q[�o3̙������2�i��$�}<�߱	u���e$��v��ƞl;"i^#ʦ�Om�bBj��}�P�?@�c�����X�nR^fw�OK���'m�0����1��4����1������5DJ��$���Ǉ�fS��$4Mw�7"�ʶ���\w�)F=�nf�6}ߺo���+��A{��c&������u���@O�����r��WW�ܲ���o��ﮪT������w\r_�(��DW5!{���k���o:�NU|����C���=�7�I�<�`<v�� ���D�Q�w���5�NMF^3tP�F0M֚��z�)�}�����/yni�ܺ6'l.�RSkᵍ�,�[S��cE�mØ�{�h]�a���і�d��">����8� ��N!f$Q*G�;��)�o�����ʥ��W�X=�+}�;��Q��&��.�/�w�)�j���6�፻�S��*Wcڲ�t����tyO����Nkk��:~�cu|�����9L�i�^��TkϠ�J��{��AK�K�����ޯ{����O{����+�j�~b�F&�oM�PF������F.B��U����'�i.�ϩ���O��co�µmjk�^�u�e��Pp,��M�Y	o��mO�����k�6����0���áo�\��k����쳻�)~�T��{W�S�4ߺ��\Rb�5
�{��{ʚ�ۧr�]Lt�vO-!/����]�~�W�W\���-;� `g%�[��b�/=�t�^߷�8]H���6�����]D	d����C8'_bq:��6���9���q^�SX^F�P�u0||�龋ƾ�x�@�c!�6�r 1�z�N;�&q������/�@k٘w+k���R�$��K��H	V3z��lGPY���˶4�f�7Y�`u��O���ݗ-��>���$��ʋ���mWW�)÷h�Z�;t��uM�
��i��%�d�t�fL�m�����)Z�&u���SR�4��?}܌�i��
��Gv��;_=�4G}�p?L�ĳ���������%Y��'�j>�ސ��s�i��>�>�ο��.���as��⻸z���=M�;���j��E�R˽��uORrj�v�����a��;^�U��T��i~�uh�v{4
O��%�^��FǣT>p��^y����N 3l:lGH�����VuՉ�Mq�WYv�]����7���+{?���	ʧ�}��>1CG}���~^�isx9�J-�z,֤���}�W�����]�6��h�C�ʡ�ќ�w��fb%�͑���%���e���X�r��W.���u���1���~{p��/Uħ�ƫ�At����-ɬ�yU����筅�/0�B�O�+=nR�ڡ�@�W��b�=3�x<��{�Ϋ[Bvn�Z����
�:` �O�=������f<��<r�:Hա[�A�#�����&�#��`.�u��E��[akP�U�{{9]����k��-b��
F���]4�ml/{����4ծ��"Gb��T�2��f�V�v4�F��֘��K�f!>���\!�0���>���e���s��.�UB���*�P� �pJ~��3s����9��T�w��[��$""���W=��v��s�{������^A��~P��܎ߢp�M/n�FV�n���x�����ݻ�\m�w���z~����x������H'��`[O�.VV�x��YŴ�q�A�]}�eV�}�T��"L[���X����]�Nי����b�t�q|�ж�}6B��\W���]�{Ŏ_�_K~��T4�$!T��O�o��7V���JZ}���qG�'u�r.��v�n�ـs����ls�:Ҭ�`���s�:�W,�FN{^��>�{ҫ��챽P,o����z�MP�]��~���{yP�~���H3jO@�t��nw����K��ԬB��B�cz����/]�T�����|��l_{�w�ڿ�>�y�hW�^v��	��(��]���}��}�Oe%� QR���Dl�XT�sT �k���j���}�4�-�r���n@��({�\5�GdhP�vGboR��n�����y*NQu6�߄�h^2f�[��nr�u	}�t�{����J�0�[S1@�	tz��<}@�h��zwxM�������n���|���m�_𾡫
��l)�uB��p�z�p͍P��*V?m{Z��;=�O��	�1ϣ��P�ɺ��'1D^�B;��C�ghy��s!�Rk1���=}��ﵱ:��^U�QF��{rм񑗮;��.�T�%���e'�U��ν�cs��U��.`��ǩ���߽�r�܎��n�U�[PXy?`�':�B�T	5c�"Y�}s9^�l�Q��Sn�5Nľ˰��ɢ���,,J��T_g�o��v�՜K`�"W�,�Ϸ��`�//�v����V�nB��Ñ1�^{���b�Bü���}���BoyV�6����h	$���\��b�q�j��tq�Hї�M���b�8딛�m>�����t�Ұ�L�:�w��C܏Wmu���tz~<��խ�K�Ͼ���P���V�"<�P&,��31��qli˨�U�� IX�^:pL-�}W8+@�����;��)j����s+��rW����qu;V���YX�����S�nN����R�y����V�m���Yf���P�P������K��Sw-�ҥd�o/�T���-��t�4�>����t�qQ&���Z��bl�H�{�:���R���:Wo #�Z��4(R�al�)Cof�N���͚�1�J��
j�\�X�Ȩykz�һ(�G�d���U��
q�,�;������j����Ckm٥�6D*�e�ۜt��Tݡ:c����GzÍVwE�g���% ��v�l�su��ɵO�ۮ]��oΒ��i�¹�"�)+F����� \\ ɤ07Pآ�S��v����q�H�R��\���1M�υh�kz匸����(󼼇H��M[͒���B���9�hξA�<���i�9�:_*ai['ݚփ�o�jԶc���3�lI˪3:d�d=�k��0�6N��gc2�lmo
�I�����t���21�̇vk}Y�O�kӥ� G>�Zr>�k2��N�v���fo�o�o����ȴ�nn��4�l=2WR��\]>�{�IH�4�ٶ%��sW-*�ջ��s�͵M�M�W]�ӏk��ט6DA�L2�d!�)P�39�Ik�(�y�$ꊖoXh�]i�s�T`��W}��u��n�b�nBOTE.7�'i�&��Ƿ'^�N���õTٳ#�i��"3k ��(g�jHso�څ`�\�`K:P��D���V�V��{;5�p��CY�0K���ݘܳ�:���E���+e S�����vbx۫b5�t$<�k��hiT:!��rd��d
�p�]�9�]�x��,׶�{Q�J��c��Y��yQ-4��8�c5v��f�f2��j��B,s3�-4��=�=���2Q��1<"��M'0���aX���J6�Y��s���Jg3=A� �{�Y{/`J���X���v4T �4F��ڋp���k���h�+)��H�����l7]�.��|E�c�7�缊�����n�]�HΫ���Sq�ʕc*�)�Z�����OwT�΍v��̣��%Q�B�-�q�6�f���,�����h��g^;�y��먓Y�ēvm�ju����v��)A�K����f3��H���V�M����C��N�M�+��� |lʹ�u�v���Z�v�t�s\qҫ �ݔ�G�!˻�� �v�#�(�=�"M�k�P��H�u6��$޵*��
�r��|�L ���-RNY�8�ܬX�tr��@)Y��t�]�Y(��xы�Z2/y�Z,�� *c-�V	֕�%1�lngjqa9j��S
�oNN��z���QtH�F.tF�ˮRA��ju�WL�M:`wN�K3_�IFP�b�C�z7�zu��ˑ�m�[�����z�g^���V�����?J���O�z *���A�F�ZD$h]�EuJ���M��IAE� �0��"�y�E*�PTWT�\ ����r�k[��e��á�K�:�-ww"��=��z!�8���{w��T��wL
J�M��
s�p�]�$��M�=�=�/D<*J*���YͨV�
*\��M�	dW8�"�����<G�����]s�����į:(�
�G>�z��F[4F���}y�T��)��ȉ��1:�����x=id�r�b�R�P����5Z����
����͎��]{��r�̪'�]�]޸��r�EV����N�h]�%/w+�<���Uqdx�HT��U�d,�<!���Ü�]Ǔ�`T�w��AU�
�$LN�]�YZ���;�/q�iP��T�H+D�E:�z��pv�WC煽G9w���=H�q�V�$ԍ#w{��:���T]�r�T滱y���zY��[-H��I�E��\��e����,���7��ӥ�N��[�.����Ω�T�VUu��R��90�}WWR�M[�I����Y� Wy��%�Jsd�:�F?�����	�@>G���[?��<7�2�A��Vo�u�;7��kpn�����O�ͣO�ٞ��ǝk � �9H������M;���1b��r��=֬���s�[K*_y]w[*���/���N����\(l`�Dv�H�x�`�����ӟ�ߧ�=�/4�ǚ���k�[>�W�O����Brr��'a���w]bR	�c�nO��:�{��-�o��N�3�*b��?0��,>�僫��w��7OFABjV(�x=�>���ݦ{�ޚ=���,b�KC���2�1��"3݌N]t���>����_v&��7摉�t����G���Cu��VNPz}��U�;���3�4eɅ~YzgjCۈsY�&��|2��ڏ�F���Z��ڏ�;sʠ9z/g��z��z���\���0��R�+q��1�n�[�2�6f���W!Ї���U<V���w��_E���k�Z஝-̥�l����4U�Ν�V��uD�>��Z�"�iM�r��q��݃�T����1'-�Q�v��]�T�97���&���pŃq��:�m�p��&�qw&��<�P2I%�,w�W�x%�	l{�P�����ʚ�ۦ��:�\��<󊋡y�pg�W)i��3��{�Ȑ���~KNz��j�W�����Ewj�i�o�{��	�W����/V}!��ݞ�g̫��|�{����|;��t 3Է�%rZiR��]�c�;�Xa�����C�f���*�}���}��,��q�|�M���x�u���]nh5
D;���^���Dm<w��#_�u?�����[�s�i�O����0��Qhި�>���ۥ�6�Ɂ�sͪ�yRҖ^�~�}�6)35ݱJ��37����ka����)��G�,r�5�����[��녯��0���͵΀�UO����?�CMTڎ��h����V}�V$u�I�x��v�p�Y�_W�uj�N�x�]���z1�X�?t����՜��;�D�M���FӜ�ZP�i�w0�)�m ��+"�z��Ř��g��\
Y�ŵ�=�oT���M�j\t�z~��R��9�cs�|/5���mT�9>��Tkm�}.���݆:�&k0n��i�'v.�'�`Ǡ��]qkp^��q�_�Wn�v�L�:V�#'V9�	����h�]6Uz`���tT���[�1���7=�}WI��ܜ�_J��s'����M���3o��
�tzn��=��q�+z>����K2�i~��#��[#���~
טm�>�;vϫèG��HS��y�~X𭘼07�{���z�����k�;�$s��~���w}�j�^s���C�̬�.�A<�0J~�F���5`z��N1^dٹ�������N��Z]Z�R��s�מV]^A�B�r�P�؅$�9C���8�;ݑ9��ouqi��j�n���w��u���頇�G�g���1�2��{=�].��y<<��B|�wi���o�:o�Y���V�����#co�f��8xu	�(oP�C���3�_Ssau�X8�����[S���Z�s�tMd���� a�C]@��]Tժ������i\����	L�1MY���p12�S#z)d�c*�0Gu��h޼����ԓ7:�3�+K���m�MbZ6_2�0K� Kъ�����zglf�����V@N������o���N�����`Z����l��#���&��Q
�DL��Q�\m�V�|ܿ�e�V������y�?��VZ��RXJ�����#2={�5�{�l/w9�Ov������zA	��5������1+��R�K�I�~)�q��wSB�TՎT,��~Р���xC�MzW���v~�z�Z�;�-�3R�~�^M����B�\��kƬB�r�	������D��y��0��"����{h&�tl�g;r�(r��Jb{���4��Yc��BE��x�>>w0p9��:MSŃk��w��!47�l]h�T�]]XwO˻jo&�>4V��L�1H5��
�ܞ����ؚ3P���#;Tp�����yv)b��w8ͧƋ����nO��O�{j������dǹ>���u!�Ϲk��0�z+�o&���0�Y�%df�l��Sz�g
�|ڗ����Sn�v%�]����*��u�WR_~5ԟ�[��9�M�5�ۓJ���l��<*�P���)�s�����WPj�����f���e:˘W� w�6z�b�>�X�0��p�]ݪ<nGS6��f�ѭ5l�p�{��yM ��D	��;6�v�6(�CNRGE�=��r�O�m>�~��t�����"y
�vy�9�qa��/�$��-;�w0B˟-���)�!5�e}�{Lx�B~��[���R��\30�ԣ@�������=W6��s�#,�<~��Oŧ��-�%��Oq��a�&#��p^������'��0U����]P�f�Ǭ�{S����)n8��:���,�g�L����}k^Ҡ�jH[�� =��e��L����Ջ{��W:���,��5ow��-�X�d;~�X�ې��}��Q�^Z���"����>�V�����m����u,����H�c�F�~8=�����
��u�o�o�Ք��~ν|��y�>������>�w��`�P�C�

����Y�0>�Q݉���[���c�]�����+�oE��Ln�u�X��)���R}O�>����w�#=Qtiw?��4�{u�g%���g3��ۄwm�Պ�uS����疴��Г[m��͘-��pG=ۇ�S����#KpX�5��"z�<R�{���������7�Ue�!��� 
�����jN�6���՞���.ѝ4]���L��3�;��ɜڑ9�y%����&F��R�pm�'��d�Cf�P��)�1H�6�^���r�7����=��39U���mm$"�-��5�(4�H�[�Ef�1�D��vT��e�N5o�����iӱ�>�͍��a,�����}�C*ˍ�����ܸ����_+C�$�t�.����c�v=S�0����������V<KVNo��c�g������2��������-���lvj��a��U����o�?]����5N�����k̭xU|/ �!?P2�T����!9�g�л��������p���z�1�w��{}z{'�2ˡ�Be����G��*�T��%
��C���wM��|�i�����/��;_CfU|E�Ps�W������3s�{+����}:��y�=������]�g��C����+эb:�
����f_{�+��ۼ����)���C�_��=�����K�5^<[:[ �n�o+�o[]1��<��؍@��ʰ��Z���ˠ(v^�+H���{�u�������]s�Q�o\�f01�V氡��`�u�*M�}"�&��i�,���N�Ӕ�r�p����o��_&;�������WO ~���`�
�>X6�]�+VR��oݏ���b���r"���wu����B`z�t��>czC�kX'��[�n�)>�ߌc��ze�ً���c��{�ĝ�
s�X��GH�h�? ����k�sr�nFg=�S�~'P��V�n���J���]b����G�^��.#�1\�p�ﯢs��D��d��%�&;�N<N�s�($�����[鍿G�O�F���g_+����RO�6�}�S��'ypߛ�(.�6���@�boD�Fw�Ցy>8��3���k>��_`�S��^a�o�½�Ȓ�w�^6cۍ{�e�½��e{��07 �޾uZ��kXy-�̣6��A]����;G�?a��謀�2���Q���0J~�G�c}�Fw���'sL���:�
�r�=�ޤ�RSΞ�l�j���~r�D�T�DncN��o/�c������rU2��N��}�G�����h��e��mf�G��u�ӊm*�x� U�T�J�Y�o@��H���fm�1��0:�w-^8�ࠓ�RfD�^���V=��f�D�pĺeu,r��eg)�����z+cB�^�P��j\۷bW+�����������.���3ۙ���\}�AWz���M,��}�7ˣo�Z��`����A��������<8zAA��:��*w���}Mͮ��8���UX�Գ��p��:���v6`a�}_;�uSVeu��wx���$�\`����,��2V�Z��;����s���\ʺQ90�����z�Y�v����v�[�.��,��� ���B�zHMOl��g+�2�7�s�.\��Re?m���	w[�iSV:���@�
=�"�{��USPv9��{����T��}y6�C�ǟ4+܏x-x�,��ɹ���6c=;��3��`��&���m�� gg;�
���؜����ك$V\z��O��C�
�S"4b�Sś^ֳ��Ӟ�&���t[��?C�l��H�qc��ʛIZњI�8%}��Ѯ��ѯ3fr�K�t#�Ԧ����6-+�N�Rr�wz��NVV��&�}�7�Oq�Z��p���b�x�o��2kb�/pSX�������nS6�T�y�^d�uJ�Bۊu��~�����fYT<��)��(������v���_\�G���[}=�ި�v	_-���%�.�3m�������>��9���6p�EdX�޷�ޙ�f�������}o)XO����eYU���uLſN]} ��$�o��{W�`�-N�R����6�}k�_һ.��z�U�j��moT+�z�wي厐�Ħ'��o��E���2��M��ӸZ�ܽ>�^���`��C3G�s����:ǫ�vB���M��M]�w#ٱq=��ۘ��u/r�`�u�*��!h�CMm&b]Zq�R�5XMT@;��Z��5������q�O�v�muB���c��;�/��wz�;�+����	&2l����l���	Qcrt�q��y��)ˇw��N�{�y�Zz��vUo>5kṷ�u��ݰ�>�J��"��|/ �vnȘ��C��|Q��()R��4�
�Z� ���K9�ثwp��2� wV\e�V���>��s=bAR'����71ʓ��M%�
��N�f�_ý�x,�:�C�v==�[� �B.V;U ��q�ћV'5,%�K���Mq�sۜ0{
�v�U���`���?7М��ݴ�}6���}{��E`��S<��������P�W��&������e�y�&2�r^V�Y3�8��u�<���F���o��}���6�5�9{1Wf�Ƒlo�4�SN�<����ъ�X� t���h򟏩�t��zw��%y5��,�{��͟f�N�SI�A����L��Cf�W�aL��TC����<�oz�z��k��������M�o�摏_�颰mA=����"5ާh���/�*s-r�gO��͍��
�Y�_ɭ�m;s�z��a�z�����2|qmA�y?`�?z}��޷~���=�l3����p>�'%M�˽Ȕ3�K{3���M��A���د�5/}���c[���~���[�=��k���ߗ�]�̯��t/ �	�
�KN��B}�	�A8�b ��f��wE�T*��^��&��ɜ���qi�s5
}tyN,G�<}j�$�*���Y����SA�%e���k��%��Vt�Hh<����m����h�̳ظ��n�21���#�E�Z1����#�a;�l�`�{�^TՆ���")������-Έn�����6��qR�8��V�4�< g�YV���H�Z��;j��qW@57\�T;�[�z�r��f�Pe��D��H�c>NM��E[*��n�[��4�e�l��}ՑÛ�����p�s�T���+��F��z�N4u�گ�.WC���nE[ڦ�a��#�iR��{K�y�M�T�dCg.��{<|�c	�wr�O+��
���n���B5f����m��m�V����'K:�9������r�EN���FH�X]m']v�Ӝ��\�	�������l�Y�۽f�fjj�e�%�V��k�B��.�QS_)zd��";�*Ê´�s���^��N��B�]ͱҌ�k�ei�xge���&PِU�lĩk��ԭ��^l������si.":e��0U�hi���s���r���	�J���� :���k����V%�J�� �/z��&���siͺ��g=j�!�2&�V�ݶM�v�4�:���උ[���o�egv����i�����.�ƺZ/&u���Z��=�X/~����� m�I*�:�4eY�oG*M����^g`[�Ж�!\�ϲ�ǉ�A�XF�=͌�[^��Vs�w��	9��ˍ
�cu.�(8R�E�}�)��A!c5K4a07�ʍwCGpo��]؜;y0`j�}ާ�BC��iR��'E�^������AI%{Ru�t��9��Gw�6�!�]y�p����-i����-tKv�Tk��'zɛ�����>ot��*�_b}ßhZen���j��� <c�����'vg=�`�l�VA1؏�֋H���K��4VӠ/�,��*��f� ���9g%���ļ����vQ��ΏH�kT��Q������R��0^��CW:o`{i8*\Q��$=ze^�[�9j�m�|�)A�ݢ*��,�֝��t��E(G&�*�*J�dUƈ�ZNӼ;���q��ow���mo8��,��s�[�V�b$���D�@����+��!�otuv�yU���ي�� up�,Y���L	ê��Ǻf�Y���c�qó2��t;���4ek.۳�Tf���M<=tD޹{�1�����6�s���3�4y�n��r̵��LDwv^D�gJ=�,]S�u	���]e]��<��gcY�T�9�H2,��و��w�2���5���ͫ����m������{OxB;M�O	p�e.��a�8�υu�z�1^���v�7��_\8J2�G�
ڏOM�}D��mz����$���mrz����� ��-�8�Tx���y��֧�_9��b��޼�[M3��d���oA{Ϛ X����˧K�n�I3~����>��!®2���V;�{�q��z��pԪ�DE��ZBQ9\B
SJ�t��EG
�NUU�,]]�g��%U�eDy�^D��(�M:\���8f3�/����}C�|�8s�W՜������**�QN���;"���
U1�ΐgXQ/2�rJ���{�w��QM֐\֜*���ge\���]��F�^�d�Qy-sەY%TU\�J/�'3��w��"�(���y�,���'3�.y�����Uz����ݼ'���s�3P��@�><�DDE�tG�Y�]ә$r�(��G(T���,]ĝU�w�q�*�G|�{��/�UG�YŖeDE5B��"�2�P.E�\��(�8�h��T\������9\���rH��8���S����h�W�ȋ�VE 資����Ͽ�׿w���F��N�i���/��g�eԶ1n;)�u�["�s�'^Ϧ	��՗z��S�0[���wc#}w�^��otEgo��+݃��������:��2ˡ��!�[hC��:�����w���]���g(��M���/�����|�ʾ��5u�j���ٵ�/̴�J�(8���Z:��N��3|�N�o�|�u=GV˛�.A�S�1�r!o����3�P��ޓ�]�}ueu���s����)��7X��R.:=�����to��퍱Ô�|�mV�ʔ%u�k��G��f��W��~�rK<W�zi��<��u)��S�)���q���Ǯ��Z����/���/�,�zM}��OCMM����GAA��[��^���z|�<��̓�v��bK�t���a�T�c���::)�,W�&:���o���qS^�>O;�N<N���_$�������Mߗ5���tvc��g�\��)����k>���Bho.�+��jø�b��,č�1��k�N���c����T���� �Z�^3�6B(��g���$<��ym�P��7�G63&Ǐ��\i�X�}��ܑ2������i�ʺ-b���5�X�nRP����|p8�ޒnJ��Kq���Fn�)%�L<�Ҏ�R����<��͎d1I�Ʋ�=}�sC�µ�I9PP���t̉��������B��_g�q�}1�`Y?`n~>����޶t�s�^���$T���������ڂ�
ӗ�7ޅ�x2�����0J~���.l՝����q�߻�fs���IP�~�-Z��t���M��D��cM=�o���9��b�m��$^��m���er�q�{��GX���'{�wj�[�z��c$�3e�V����?���q��w�24A~l*����'���+6�f�P�C�����}Mͮ�G,�B'xy��+��fߥ\�����C��'�
��U5j�������Z���
�ö���y���C��M�˻W��N�J��7���>V'���ϳ3*�F�h��[�	���ye����>�7Ov�Xf�mЦ���̫�:,��Y��a���$�p��)g|2�4��ޚ�_���]�^V�[[��zs�ٷ-�����[nE�!�z+���V����@�L�B)n<�a�bV��ۑ�Ӵk�Ƀ �W�2�f��oH���'u��-<z���3�[3BU�n�j�o��{:hG����omj���-~����K�V:�V!H����1j�rFY�������9!e{?&҇ՏU�����Tq2)2{�ձ�#6,璛��G�xs����d'�������HP��?M��S��o�H�UuY�d��/E�}���Tő��r�,����w���9�ϓ��5�T�f�Gf��w!b|(r�Z*ƚ�=~�,)c|j۱�����r��U�ȏ����fz����N��K���m��;0E���g.�o��~#ö���Y�횝Yӕ�M����*	�E��ʲ�mE�;��ʄ���5�U �<+��H.��JX~�M��;��_-�����
1U���ž����{�M��f�X�P�á�_XI7�w�P�8=�c��|}��ʸ"C~���D��{r9V�6�&�I6�M��������_�s�{�g�@ᛆ�	\ tD\1vJ������F� �f̮@^��wS$�}�[KǷ1�K�1ٺ�	3��lNn�,g���[:oZGs��K-H�aۆ�F�d޼TZA�0�)�2�I�mԶ�1)Ӯ�\�����t|.����н�����w����95�U�k8|j�������s�h�B ���x:�;u!�ME:dx��o:����r��D���}۝Bo�L0c�����^>���4}1�\�����:�>��W�F�ӽK���U��z��!ll��q�r�wP ��.�`Z�Kx<���=3���yHrhտq廡cκ�]'K�޿�ݪ�;I2�%%n���9�����j�'��ǺՍ���J�������� ��+��tsmlq���=l���c��G���o��'�#��2��"8dVc�o�BK,�;���}ӽ�:Dn��?h�?0Ԝ�+A�g#�u�tFD���W�|+3�X�t�ޯ����u�?i���ԃ�~Yc��\�ۊ獘�k}���}}O�AOس��M�6��=�n�͞��0C\WLY
'4X��;�bE�6� U�-y�b}�����H���f����,�V�+��ޒ�NrD�p�֦�(=W�����X Nĥե@ₐ�nR���ۋ.�uYW;�p`�j�bݑI�_��R���3��{J�i�|�ޗ�'$��e�9��&-��r�����3�\��Y���u
��7$=�t�-��Ҵ,���JN�������c읇�f��O߅}��W,i5�p�&b]���VHٜ����|oq��a��J}>�����N�����o����\]��v�!y�W��w�YV]}a�u����hP��Y/{p�vv��{���ӛÛ���i�v%�R���k��^A����-1B%iQ��b�#o���ep�G���E%|eu��_ͧq��E�!�;J��e�D��>��OW����q#��y����I-}�w�}�p�f.��^9��`�b��X�[Luޗ_v3?^��*|�g_��*��3�μ�1�7V���/�q���T���������y�|/��͹V�^��
!+�%sΌ��U������MZ��ޘ��U�Z�U-/^&ۻ���^Yƒ���!ٺ��9�z�������PސBj����͙6�+�fAq��b]��3���6��i�����L��ӷh��=�&,�+;�z*��p'���{)���Ojq��S���&�[��ZC���襽������ݝ����q<X���*3�P/��"�o����\L���{Q��5Z��R\V�ޱS���8r���u����ߠ>�s��@�B����1���Kq5�=/�l.l��1���*|+O��g�,{�N�/�WA��KM�Ls4�Hs����&�v�12heDfc�7��*��φw�Rzo�p���b_o.Bgޝ��zB�&�{{MfIV�:����`G��Rk1�Y뱾^��t�4c��[�8��<+.�__���~��k��a�3/�V�#P�\s�8=2���KGlz��[�����K��к��*����N�S�*ϫ�X�}��
����U�͵C�y�ɪ�Ԕ�]����l��c՛�JG����h~�](eI�(n1?^����MfZ-��x�xE�1�+m�7GN��r{�Wc��w���m �M�촇6�:�g�y���30Y
%�n�?(��H�-������T���a�g,��]���G8Q�XnE���j��k��q�2%J��h�O��ܼצ�2Dbљo��GXi�c+y��N�}g"���F���G��)�Ǭ����(�5n*ˣ�v�pn^�Ͳ�l��\}��(�ڋ���~�l�SU��Wyӹ��}|�~��/�C3�(�s�o{I{Wy�k���mt���XOh�}_��/eu�K�1s蛱�w�q���Ln�5��n�O����t�z=@��5��9b��sX}Us�}}C7���;{�/�{�����M]S�Uh���uu���R��H�P+�{�KGj��@j��K��SJ��Ԯ
}n�m�H����hp��n�0{;��h=�M���y`^�����_W�BJ��-������Dx5y5�vm����_>R��U��T8Q��-��y;�z��}�j��.�`�1H9Om{Z��Ϧ(��$!��X!��*�:�qt��ò�]�W�Sb�>�Z.~�G��S,b�j��(����|#���������y�S_,j�X���m��;0~��9�x)sc��2�����9B���d��l�������J@�ݠ+{�f\��q�O#IC��\0e�X�N��V�j�,�s����0�V���鄷{���Τu4��z+R��Q;���w�S�i� q!&�8��N��o�88�����>׾��C:r��7�Xt�}�C=n�U�P!-�Y��V,�ge�_V:�m�:b�kwꕬ<�ѩ�mK/n$�������Ʈ%/x7+�.�����_�Kb�<���8��Ƕm�=�:��NEw_-�C���<��̭�髂�~���-�d!?^�^���*�c�*0���Q(�ّz���3=����:��E���i��[��y�A|n�s����tjމ�O/�4��:���]��
6@�l1]\ �����\/�K<&T�[kr��:-=47�k��T���[�����.�;S��ϖp���
?ze;��{���G���[����",��~���L���5A��09�z��]�S��^�om���\��A�\M!1Có}).����}AP�z��9�Yr<�r�T���Cߚ���ݽ{�+�nr��ls""�9Y(�{�������hH89EW�Pݓ����ǥ;��x������l47�!ˍcvlҭ�����p�9�kWh�e=�a��*�e���[�s�������f,<-E�Y��|)]���[}�H������:�0�/S� �������k!�x店H5?�+�m����O{���P��y���}9���7��bR���W�O!q�u�#L1���L�k�Vd�(i�|�h��'*׫�^��ōՎM����2x[��<VX�)�g-�̺^���ޑ��t�T��M'�^�X��{��M�o�4�e6��F���X�B����x|]L1�L���n��5���<6+�������$���������W�f���ˎي��^>�/
z��=S����wc�V's)��w�x����t�on5ٞVUXa�X�~�����B��ח���-'�HjЄ�r(y�ܩ�mӱ/���V�.� �	�B��H��Fi����*�F�6��(C9/���W$�ͧᇳýe�s�{tk!Ƕ/ߣ�-��U��X�T"�7C9D�So>��X�J�K_Z�&��Fso�)Y_�?.ޡN^h�P�{ҷ�2�-Mr�I�w��8"��l7Y�]+���'8Fp,)���z�����!J��,������W���z�=b�ӓz�v��\�^-��ㆈY�D&�QJ��WRnծG�s:,A2T�k�k���h�ObM7�+�����?Ǉ����������������n7d��5t�"�a���@����5�?@�A􂆭�}�Օ��uB��>�ņvf��^�Az͏c�K���_)�~����>�_*ڭ}*��GE<��<G;�O�_z�纤>��7�̕�N]��}��HC�(oI	�F�=]��8ŏMn�k����V��֗u�ݡM�f�̟]S�zjoaڴ�yүwO�ٹy����Ķ�5�6Z��+�������L�V�t�F֋����h�B=2����ԓ}øb����᮹q|<�8Tm���6�w�}뎟�1����:~5M�9�ڤ�!;˃�u�<������N�K+ˠ��tߦp��D
e�S�Ʋ�=w��y����'`�8s1�j7,4�Ò��nW,(Щjb^�%+\1��ci�{�{��R�pEEi�EE}���}h*��G�����?���� BN0	��; ; !�L � � >G���� q����`��1ñ�Ȁ "m�1�Ȇ�d@ ��d�cm�8�l���#��dM����D6�#��dv6��m�����m�Gm���dp ��dM���l�m�D6�$��m�;l�m�Gm���dCm�&�l�m�D6�"m�����Gm�6�dq���l��m��țm�!���;����!���V���� **B����&�\}��p;5����U�(|���������?<_���\M�gr�*+���}/���
���;�Q_��:;"�nG3P���v<�E�;Yԇ��@����x��S�9�y���� ""��  !E@AR�@T �L � �!�0� �̈́�r��?�PDV@R@R@F|�q��GN��(d=�8zF�TTW�֎%=��(aU������"����
���cc�z�-��x�*+�E��Υ�����{�A� U�`���
?,R��
9я���Cّ���W���Cy�8�È**+�V��|��nf绐ak�_�u`y�c�P��	�
����8���{���r����9��GO[MrEEj�CG�Dy8�`ݩ����EEx-J8;\�
���~f�\����(+$�k ~�q��0
 ��d��I{�R����T�J��"�H����$U�
�RHQH�H�D��)
*�B��T�$$�����B��EB��*T)T$��UQ)$)V��h�B�"�I	A�IT)Q	�*��J��t5"��� ��U
�U*�B��OF��U*RT("��IJ��
��"*�*IR��TBU��J��B	  ����$'�*DF�	/   ;i�=ip0���N����C���l��u���wT��p�[�;��WGwp��u7n��hI��)�U��L�s�T�۹��AC��Q*Cl"$(P*x   �뇡#��C�СCާ8z�
$H���
�(�dHQ�Pȡw��B�
(z��27:��m�+w[�P�ӭ���9&��v���;�
��VV�j��d�*TZ2�El¨�^   k� ����V��u�:�Ki���n�����T�Ս�w]��SM5��-:�n�,3MMm�@av
ӡ�ܗ-��S��w9\�km�n��jr��IBEH��T�/   ״z�i�6�r�h���l�&Z�uΩ�f�i�b�:�Xi���kmݜ�s��P�]wt���v�K��E�j��Q�J�UB�H�   ���W@lVP��V�j�m��bIh66 *�X� Pl�J��
�QQvak T����H���TJ�   k��*��� �*j�5@CV�T(S�����A ]` ��6���Y�kE�f�Z(m�!AT)$����  �Q�ZUZACoZ�
ִ�l	R�ch�["(�U6ԨF�UF�PmQ�i� �1 $��(�)Dx  �<� ޔ�@ 9`   �r�������:R�7T�: �Ai���X t�;�`��nR�%*" �eET��   v�  �ހ@���@�s�l4�`� K��vq�B�[� n���] ҳF  ��Z�)T��R�D��	^   �:�@k:0 ;a��  +�$� Z+S��;I��K�`  A� ���`@t��:�@ x)���J�� E=�	))P  *~��z��@ �JR��  &�R� 0 �)P�U$ hM*�[���H�H��Ƹ�L��J�LP����U�)�r�e������7���\F�������m����6m��`�1��C����`�cc�����w������;�#�9XfP�o0�i�M�2"�j�2���Z�e�t ����P���\���Z?IM�
y�^��w�U�+-�dgocvĲ�ldw�rX 3�-��w�C��A�vɓhe@�"�����%
�/�*��R�4�Kf�u�e�5�hV]-2�c8 �=�p�p��&���cf��Akn���K��k�ǛW0�93*!om<̥�*���ygoB�K�p�B-�Lۧ��$b�)KK�EJ�R�fIA2�kJ�EG�%N�6�YX^�)��)iK�7.�cJ���[.}dK�h`�!n�Q����3.J��F.P�%�L�Z��N��DF��*Mմ(
�ī2�GmZ�Ѭ� VF+��\��yb	��0=�۩4��S��϶�i�uyb�,�۱)�"#hҬ�N��X^]��[J�6��y)ݩ�n��j��m���u��(Xύ���Zw)_��l�^�P�R	�ƫU�ux�U3�d<��k�R��SB@�kq\�FB�,^b�W��KinQ��@� m�w&��[�~h���7�dVL�R��(P	3�osR4c�R�q��j[b۱�j���7,6���{�#@��
�UƶS%Qz�.�\�mVR�qK���	���D4�a�I�l�B� E��MHٳ,�W�ҋE^��r)���J��P҂:v���g2�7bD�
��0��_��1q��1�{&КEn�n=��	n�%�<(^U�'3T9v]^�fi��D�͘6jE�V�Y��D;��)n��/,r��6��	��f *K�a�$�Q��r�\N`�M��F�-Q�W�r�ܠ(�(�Y���w��72-jɖ^bB�<&��n�kp4���+(��\9�[������AKIQ�Z�oV7)�0�tZx�E s�IS/Z�˼2�e�P�S[WwN�adF�k�$��Օt�c�ͽ�h��`YI�[h�6���)*��`l�ۻ˕�sH���مм�M���PLb3.��Mf+�E�ѫt6�u{��Fk����W�&�t��d�"�9j�`@n�n|by��Q����!o�)�����)-��nԢ��f4�cf��r��)
U�BGX��@�Lm)�Cr�f܈�½�`ː0*o�תen��f��Zob�����b�E�)b46*��M����iʹ�u+&V�Ic�k �*��U)�F�$��p&N��f���JVͫmn��R�2�&L9LM�ҕ���o�9f w%�z�=�X�,4���uq���m�RJ
+�d���T7%�U��f��J4�wMD�eg�Səd]�S`�1�S�2jyzh���sC��Jq�塵�pbJ^�ݵ����[��nm�CR��h��T�-��^��I�R�Z�c�5ɻ*1J:i<͐Tծ`��0f]Y�m&���%����V6)�$`!!��)��h̼#B��6��=v.����[/j��[f�su����Yu��nL&�$�B�f�2���j����K3%&�{��M�a�6I���cF�Pܧ*H���7�nں�w�S����^����I�a�l,��h7=�wV�J3�Gn_��ź��f�C+.�;u��.�j����׷����%m��{>J�)P�l���33%cm 0�TC����NǪ���
�BY-�{N�^�WCj���Zӥ�*�2�t¨�i�sJ׎�R���DZ�SC��Z��x5\�V^E.Q��,bKU8��]4��^���n3%1�b־�
��KmL�Q-:E�CefB�mn\F�ۋU��Z
�-�F��:\&̸�u����-�{�X��{��OF�З��t�H�yj�*�m���E،\P����:���HH~-��52�q� � �ٮ+Wv�����oT��Z�j��I�MU��]d\N������^��8L�6�ū&�J���r�bwZtɯȣJlَR����W�qd�б�dE7@�P^��.��6�ܔ65" ,�6��M�$�+7`{�	q�cL�c$�t�ħ��cE�˸V�E�%�Z̘Ç	Qel,C����qE�Y����ҌE`���h�hԌ��Q���H���V�`{H�bc7�	�Ѷ�����r��b��]�[;v�.�\��襻��0�ii�(�B|�Aj��R,�!Ӯ<4�6f���2n��拼���f[�ZD�X�^�O.���F�[ҩC5��;{��]�(�����X�+[�(lr�[`ⷶ���Ά�U��uIhS��X���@`��̙f��dC�˚f@d�AKp9��%-k��>ןn!X��N��SJ����Tѻ�������+Vˣ4:n�mЛOvhq�J�i���]V�qD5�e�{i��v�� H9vo6�����7@�h�t�f���`�Y�5�5�Ik��`P2�]�{��<�[R�vࢄ�f�$��K�� ��#B4̘7Kr���
��;�JI����M�-nYXsR��L%ʂjp٢�T���f�*�m��X4����u�;�*m�xiѕ-��6�!�b�r����,�N���T1�xP�QlbJCQ�/�b�)m����kM����5�[g�B�V�f6<nk����?K�Z�І��!�Ґ�i���:��/im��r�)1�'�S'D	�!8YyxwL�ʍ<_M�&�WY����ރ�N1�sG3��Y�q�Be1�N���2LF�ʫ�[�z�ٙW�к�of��&�M�Y�rL���Z�w%cwN�h���J9��6��H\9v��a-[F�)���Vu��:X�"X�Ol[3Z
�ŷ�E��8L�����`	�0i��[�ѵ ҉bL�Ւ�*�F7�l��c{�R��4�ߖ݅'5���؆���wR�5;�⊢t���{�p���a�wR7�XU�	���-��-3�-��*:qV�Xx�A�hm8,c�Zޭݘp�ˌI2]dkT.��b�*Ze���z��7\�	�����o-j�chM��DI��cO.�cWFi7[4�&)�
zx�Өqر��9,�����n�	#��� Xsb��bu��%U��7`�G.�jjw�-5��oڎ����$*�:N�m��g�7h�V۶cdn]��$r��r���a�ƍh�ˎkH832�}f��C���m0s��~M!f��5��Z�=�t��u�5�@�n�KՂ����eSئ���S6Ӭ��jō�O��@��5e�i���T�G���"h�E�tkK��J�� �5q�b�E��i���v�U(�i��B�W�2Q��3X�P"�Z���Q̋Qa㫵��4�mn�	���] ���ek��y�赆���DP�^Z�Z4���8�܂gڙͽ�$9J���/�#,`8�inb��Yt�*v��l��J �����WN�V�-V2�C��h���ڻb�n��Y!���`+jT6�c2��H�O<���!a6ˉS֋��:�y�u�>2��
9��b��W���t��u��,��1X���Z����.��,�Yxl(�]��tj]�)��:���"�Ɲt�BȊ�M��xT�TlYÂ���]�Ͷ��3�kZe��ׁб��mР�ddڛ��:/wp�Aw��knd�0���m��yV�	k�[���$6T��f
W��%!�hmi�i�4�Ŵmj"o��D��h�.�FfKn�&,]ëX��+�&nRУB�i��2dy�L�IJv���bm�vQ�Ih�y��H�uc9B��5��MĘO6�fl%��Qo�J^������� ��)�2n��BSU�ɒ�3e��\�;J�q���t��tv:q�zw�%�:=!��B��f[w,�10��{�ٹ�Au�"v*�$�;���ֶ؂�*�9��e:��ٺ�y�\8��B�	[��
A;�Z��JkL�;.R���e�/i�@���v� �ݒ�JI���6��R�̰�9�`v�ݛ�f�r��Ǎ������P5�H�]�!c$�I���	�˗ ���7X�ʃn=T��Y�r�*1�l��TP�2��AQ"��.JY�YX�ͻt)L)����1f���Η�Y�]~�e*��l}�k3p���,	�՝��hB�e�KA�p�)��D֦#4R�wX3� ����sD��V�j$EV���i�쳌J�g!
Jx��[p^���k� t��n�m��Y�H�V�RM�L�u�Nhɔ�ۤ�]f�Q
N��fD�Z]f���DyQ	-�WN`��j���$��op��s*P��]h���4��[�ǹ���Ȩ���Q��`(���YA�N�;EV��u��OtK('#��ڽ܆BA���
��V�]��"5��4/l�0�A�qKp�.¬_D �=��Ɏ�my�)l@2�ݬ��Zd-#Gh"A����i��b��Y��<a�u�Z�T2��u�4l�Yt�i��K3tf�Gq�(}n�6IoN�jL�����SL'n�B�Jb0S�a�eۋY#>©Y*�h�b��5�h���zw<H86�0�4[��.�ƫs��ˁ^�9��Z�f�H���m�Œ���㨔OI��y��Պc��Ў-�6�d7DQT�J�K?Ô�YgSz/D����eЩ��x#��E�i��h�B�����a2�P����#o@�D<vJ��1������!-bi6�������<��t[P�u)��Y���;%6�Ou�ޑ��U���7��WV�dD;��̈���yB��{5$��k.^�wCE?��CT��E���ᦉa���W4�&���*� g]K�A�5$�'_ěα7�ʌZCdf�P�a
AU�LχӬ��Zqɘ�ږ-u�IЉԈ�.T��d'	�d ,�R򂖐�cF�Ř�Uy�J���EEܹz�p]��q"t�x2�-GhLі�V��<-5�%B�-��r\U�J�B_���-�ڍma�g �QcR��7T��
��[V���8$E\W� N��ͭ�N��b�A\e7%�WK��jBY�kn�X�t��b�z�l��+zՙY7f���X%�[ƨ��cm )	[��à�x�u7p66�m;��U1�Jok	Dm-�B�a���eæ)�Y-�K{C�ec��t��^�R_:i�#N��Q���"�����gُYH8ֽ(	��.�5p�u:-�8%7���b��i-7X�]mh�T�+�����tRi(d�{����ocAhwqA�l9U�����7X��r�����m�`�h�C)�Ƶ��J�XF�J��][&�Q`���"�Uk�{K�s��A�2՛C48�ojGwL���IIv�,.y7@�^k�K6�h����Ϸ�l��l7W.��D�@j3���y��Fu(����e�5v_�@`Y��k�d� ��ش��:��'�m"���qn�!m5��F],M[��n���f|%S�r�K�[[T�ϛ��⢶���@V��RL���j��g���X�ɒ¶i`�cn��,�4E`d��;��)Zt�ٰ
q9f���Y5�!�	U�tm�'OuU���ʒ�u09�K$�y2�LD<f��j*ͩWJ^3�v;F�֠;F�LGmm)����K"x]�ejuq�ˤ�2��E �0���ދ�(��;��ק5yVU�9 H(%I��V�I��r�FR:�ډ��.n�!�2����]a`ᡳ�L�Ld�n�֪[�4�2�ַA2�xa�j*P
,n������;B�����ZkS,�f%R�9t�۸�%�V���]0����)Y�%ŋ��i�����b*&3�ȕ��i��:�
�{��f�rІ�Mo�ɶ�BR����j����
ܽ���-znT���L}�P����:Hߣ�^azke��a�7N$�¦�.�	����Fnպ.�����zj��Kd���n�i�m��*Ve\6����,3Hyq;ƷG��m�ZEgp��m�V7���l@������Sl�&���ek33c�u�Y��#mݲ��XnZ@�ik���A��l�����Z��P���y�4�^��&����f�ct8��4��MR�-b�tiٵ)e]��l�ю�J��&^:L�ѵz,�O4ŀZ��"6���"�r�^]ظcCp��2��*�w����H�KZ�51[��]��D�i#`R��q軫��f��B�fd�45��F�6�HF/�@�tlnYҊ��*�u��i�@_�U=����q�,j�<;��i��TW��]��Z�,�T�x���11�C�J�e�<��$Y+K���T�m�t[�Xw��Mx����]r�] �hƍ��	[Hӫ�����n�R1�J5t &�����6$�F-	���)I��a����ŷ��"y��Ń)1��6T;3z�����@�Q�)���W�K%�vӤ�������$ݩ��wW1<4Gb�YL�����:9@D���\��(��1�ˢӘ�ӣh�bR;*���^EN̆R���Qqu�vN؛̣���3jb�٩�YA�[O E�1L{�JzއyN�ZaMn����aOa#uT: ��m��~T��R5.9J��6֍�Z�b���D�\if�TA%嚫�y����e�gs�ݰC��^Ĉ�[�!��l�v5��[���AE|���:a$�[:��6�X�b�GXN�̕��K0�`��\��^ո�i�@m�y�$�����3 �U���`�{{r�.G%d����vXʗ�����idJ�K�X�N��ɻ�����5Y̶�T����)˲X$=(ǛA�(��_�Z;wD�Y.�;�Fh��r�J���ʳp-�hhf	E*fk�nnŭ�GՑ�'U�:�s�Ṋ�9��ٱq*ܥ`q"ot㙀��󛢃�;��j�Kx�m�h۹�1�A�T�8
w�|E[��l�t�u��-��=0.|d�ג��s���p_2�C)(�{�w�b���%0�ݹ���mlo[ŪfwlTx���-I����c�%�'A�����cY��S�8J6wT��{.�<qV�����,���)��/E3���;	��R�JKc����)�//43{CE'wt�|jW-�ۣj>k+k�)��R��knv.�"�;(��+��R�e�%�D(������nhd����
�,���XF&�|-И�����N�]Zj��r�v\����8Q���|6�VS©�[��9h<��T�SӨeε�N��IAԕ��Ɯn�Z��֬:5�	�[<��2�H��+9Z��Z|(�7�j)��t6���s�>�ۓˉ%��-�){E
�8�ov�m���p��xIS\'fcQ�ư)�Z~\���7�랪μ q]t��C1э��l�-��>��T�)�����ǝ��=ALS.��-���� D9��l!�ی-�r����IDJ�;tJ�Xi��}Yx�v:���V)d�E�%�f��Wǌ�:jVJΫ�q&�����a��z�*Y\�E����w����]&)�KV#/EK3'�B�']۷�Wb�E�|0��Ԇn�ֈY��Ư��,��/T��G��{��n���)hiOn��]�Z ���\hZm��������ܸ�*�Lݠ�'����	=��5�Y1M�%K�냐�����٤E�f�m��;B�8l�W��rW��ެ�2Vr9� {Wq➣,��Ȇď�p�8[*v�xbbۀ5%gJ�9�-�#A�]�W�"p���뙤FE�V �ԏ�8���]���$+�.m�$%�}V�vu�/id��hC�����n��9
��F���D�����y��q�;��y�Z˺U�XQ?�NJ�B�˶�w+����n��Gx�r���V�� jF)N6��ј�p4�=	��(^�i���z � ���ʦu%|��	�a*Ø��7��*��Eܐ����x�=Z(h�]͇"a�4i����+�kr+�N�E\onV +\�趭��G�m\N:;�����Z��Z���;�c��֓�R We�n�ٮ����f-Rw-��m'���x/�h�Er�lV��r�2�982����Cp�Z���c:�H�p^�&lW$�1<I�ܫ�%�w���r�l��&��S�LgO���Or���ܺ
���{�]npГ�������p��1;���!�e)ռ������,���vS�ڽ՘/I\�|�f
I!���g x=kZ�����)�f:�]'���F�x����ױ�;�����5��ᛨ��HM�WcJ�{ren��[�W��:�f<+%@���t�Y�+�n��	^U���t��q�^��ݷ�sll��o���â,o+1
�\WY�V�b�1s3y3�w|9BHwR�`����r��b���P�a��Mtݬ�������_�X4P����C#�8xp�P�s�Jw���bC�GW�W9}����3y�Ɓ���}Y������pUq�2�n��M�0�B�G�G{y��	V��1� �Tx�׼�j�oo/㒚T3�.�A�T��[�|�d�M��Cg���6���O�do{��Wg���>6\CJ�����ot�*:J����HɅ�w.&�k��E����Vi���eƆЫ�Ur�:���s0��U�Uf��#Hq�:6�S[�E�����"��V�����xn�c�!R����%Ѿ�=��Th�fK2��(+��Щ�������hV|�?"�|r5]�f�m��of�;����������^$���9" ���'��Ͷ/����W��#刡6pU�Τ=�LT`ϛV'�y;�4��i�[M=�r2a9�7�k$����qf�
��7��s�f�]! a݇�;O�d���+3�sE�Q�1��l`����œ�Pu^,��)L�ƙW��-�ˉ��sU�� w��^�W r��3�JK���6Փa:��k�b�Y{[����o��}G5ጫ��'3��Ybx�b�2ޚu�7X��8&0�����hZ�NΖ;��(2�q���l�ʬO���a�܉ڔ��ﳻn��&������ٴw)�齤��������t� Ǘ��	G��sfCL�yB�l�t��rWr�y�T��8���j��ƛ�Щ�󙦎��Z�q�-<��۝VGT8�JP5�c[�Ep��6�#N�召9jT���Z�����f�:QP�
uha[�`X���u3�K���<��c�����i�ᷩ��.��DE5���ϗ��]$�#v\��e����+��rN�F�;euB2=͓X�;��c��-�O5�v��*���k����D3��U�,9�غ�#o�r�c���3�#;'
�,6��⧕�^��i����4��'v���̢���vd��V>���F�Q6;�3�ط�^.�h���5b�a�h�n_nT^�y�oC�H���HН(��v( 8�Lk�Q_q�}��X�,�����w�8R�\��u_�t��Tf�uV������+�-���E`�����	��k��s-u'y�p�� �u�JӴ�\���u���n�F^����`�'t�{��3�f�We�
�heqٛ0�"���!Yxg]�PɅ��\]��"�`��'7{GCc���M��E��>�n��zƈ0+��brə��@�{�t��m,Ƒ;b�sOV�����v*c�c4��j���R�Ԩ��4�F�W���®fV�si���4���6�w�3���R��e�`�X�۳���f�_hgC��u�c]����V�K�;s���qw;i��=���w�� ������e<�\�����%�KeT�cc��C��ؤ�����ev�- Ҳ+�
�u|��K�į���e��Xo���K5��7�8�b6#\��QA@I.=�p�8Pp�WǱȽ��z�h�Z�)�5tЭ�@����h��ǈ�Qf�A%�>*=���WSrI���)�]$�-Y���֛ݶX���YKZ��8j�"�wuBN�9�59�r�Ϯ�9��Qz�O��l��ά��Zm�3y�����dI��=���q.�-Lr�eF��(�����yl�Wh�����q��Ŏ�l5��Մ�h� MVA��U:�VN=,4�	�$	���s�X5U�� ��r��Q}��p����꘻��})Omz�/�g�X��fŚJIĎb-�K����Gզfs'l�4e��O�h�R�(�e�M+ӝ }���o���P8):�,lϳE+4��kܵ�"�wB�djƍ����d�+����m,�֣�-ή����X�=`���]��h���|�˭3a��A�#ckV]���79L<k�_.��YW�����C(�Ә�|jj� �
�	({��*�.�����u�˧�	u��N�AF<V/T6ث}�s��X�r�*qFiB�1Kܝ]b�RFwX��dҜ�Y�E�tZI�Z��b�gb��<(�c��+~�.����_RV�Y�Іwt��B
�' ���*]����F�����1͋,sL�8_�]��۟=�;������"�o�z�����7Cse�8��Y�
��P9P]���{c�G�J�6C�ʅ�"����,��N%�oC鼝`Y/xK+f�O\J>JɃ�x�c0U�`f�͓�HL�αˍ˺k(Z:���gsxb鹺>�x�]��z�q�6�)��sF�Wmm!Ğ8{k�#qVM��2�g���-T�!FΊr��/��k
&��aA�ܣZ)�j�<ޘi��V���oi�} � ��"c��酔�X(�j�wJqS���W�e..m�;ݣ}�$��e��ƀr�2�i�ӑ�8��%�e_fq�<��}V�*W�7k��'}CS�H���[�W_E��
�1��b,;�`G90�U�:�=Gs)�0X��l��Zy��z��2�ܼ��vb����oQZi =bk]u:�X�Pb����>�wcyX0q7�;4�M�gc��]�����TE�{uר�۾*»�+�:8t��K�\PH./���]�R��:]J9���U�Q�_�W��)�vjX{�X.>��&�8����-�����*�����魌o���g���ںӬ+���V��Q;���W&tj*�ႵR��=�{h��}�sޱβ�+����䴪� ��n�޼�.ʮ0[Bq
yV�X�u/JJ��k��\�p�����u�^� ����n�UĻ�#r泈%v��3{\�zWp�Ě��}g�ocYw"˸T#O�]'��k�k�:����f��Ob�4a5�5���*��&�+Ż+TS4�����Y��tL�"�x��!+\�w9,���c0���N+J̶�uS�~b�۴������lh���G9[��ѷa��S�ߋ�p���*>�v��}�vW�e�G�)�7_E�v�9��f���7{*�r�3�+�H�.	���e�d$�#u�2�[�R��ɬ����J�0�*��򮹎2'Y�Nye����mIĬ�� ot�m㗡��]�Cj��
#vb����V�kD���F�ͨ
M��,��17�����1a�9�D�T4a�b��׆�e�r�0.Śywfw{!ʋ��|�^��u��_mi���U�T[�4�NB���*,5;��+f�]nZ�[�����/2g(M�S�W�k�N�+Ob��-���l�kW|� �	uݝ̻�cL�$�W7G�ՙ)��c$� W\��)�ق�S���J�����-�ή�{�QQJ
��m8�ۻְhAZ��,���:���s)R�W��:�v{/��J�j��3V�d�]����A�k��=��.Dv�fS�h��]fEw3��P�v����ޠ�����.��h�[���/z^k.��bo��gR��T Z���C ��r��C2��Q=ma�s �Ki:9��k]��D���X2��I+��,e��R��_);�'Te�u�a�c*���-�W�eS���j � 3��]=�[�ܔ�07#B#9`5۴�Sյ:g�[�k�f��5tﶺ��S��}�^c��c��&�TsGHq���/ud��q����(#烞�㳮��}�Sw��E��Q�.����h�C߰I}W�q��}.�*�'�\��t����|N��.{���m��L+1����{d��]���S"f��d�Yos�=�"�%�*V��bt{�	�
��i��oy*6�<�p��%e;�uy՛���`[������\��v۷Y]P�j��`���h�\���3�I7KML�խ`'�����.p\dp+��O4OIM�^�]�� 7������K�j�Vul�kD8�k���ݹ�y:����o.g.����q��Md�B��)uw+M�=rt[����gwi!�g�5A]�͗9|�rm	s��`+��R�w]273�[� U090d]��.����暘�5ݪ�̬�ﯗLq��p�6��vt���,ᫀeazn��7mQGj�z��ہ�6�:��O���i
!��D�Q�j��wZ'n����h1��ݘM��z�����4�/�YZ�0���-��.�4�Y�`8d���g�ܾ/CM�YL�s
틷[�/s.�F����-.=����ut8�f�r�;�������D��X���F�1��Ѿ��U��9V2٤{������=[�7��㔶	�nn	6l�#\����]M4׃�̽n����7�U�R������+֮,�֞I#�]�++5GN�#t�6�,����Mԃvi��w�� �*;$��enem�j�h��tv�ʅ����������H��X�`�*^n8�vjC5��� �K{q�+FhD�j�����V|�'o�p*f��i�}��Wsm't:}옧^�ւ[a|f�:����F��Xf_s�͚��;�Np�0��;A�f�t���Rn�����٠�;1�Χ�N���墣��IM����EV��!&=�"��v��
<8��E;1��9����W]J���1�.��U��V�,���өM������Ր��5&F��fN{ed�t���fVV���3bq�H���9 6�TU�j�	�D)�rTBᱼ�Wөf�ݦ�����ˋQ�Y-��R�����(Ѵi�����,�w�9i=�*,�|�ӟi����h��r��+����t��2��$v�W\��#x�`��O�	���^�^��@3�[�ה�9K
�5b����B��ѵ+XuP9�r��u�ݑ�ݕ�$���'�f^��3�l���p�{�"�w>:���,^�1��̊�؀f`t�E���L�=�$��L��b���`�Xm�e����b��Sb�oP�D��.�Ymb[w��`�I9��4�������X���!�Σ/��Ĩ���h�Tٮnf`jPSP��.�v�@!�^�ꊍ*p�ޗŔ�l,��t����T�4m�������-\er��R���K؍��{W��ij����9yP�\�`1�}�P��f���p�ͅ��`�r����u�_oG��Y���ŉ&�W|�s�[J �Ö��7���eȮDƎ��G�kr�=�|�������K强ntM�ut��Ҟf�v72l���:�]>@G.�����	��7w����ƠS	akO�O���2û�U�p��9�e���7��5�����J��7-�58_�����w+�!��Z�1pvt�Z]_ �Vltl�cV|��1Ι74�lu� �ؘ�� ��+�f���%�RI%�l*���P��6?ـ�1���߿��y����_�ʅ�=��K�T��T'�KgJ�x�ʔr/��s�[[�:mΓ�7C<]�/:��-�6@�&!��h��Zݾ��u���WOa7VBvn	�`���s�/-s�ݪ.�f(����r�b��������[�گ��jr�\��S+��6�N&�Lľ�d�ck���r�(�J�j�x9��Ӱ$ R8;_,�n�!������t���PL�'ήum�8�}y&n���W��Z��vV!�[��,+O�h���x:�=ɛFʳqpd�\�y��Rx�L}��D_f�]�����,�)k]����J��,3Un�5t�A�	J��+(B%
Nj2�����^����'wi��R�b�(���T����Z��w�c�y+����u��)qFe��E�g9�eS�.]�n�&�����S �wW�,v7���6�E[hQv�B*t!$Eg���WJH���3R��l̴���Q�M�:�Sd̄v���ٛˁYjfϞ�%���8Pݭr�+fq��;�4�!���{���B��YO���J�����sd\�6�o�nSUt���v��-PI��t�ݼɸ��&d�Ɍ#�][�z��������,���J)���owD�Z��{���1t�n��ƫU��M�k��56t7�zt��K։�w|bZ��H	��'����KN}|����\��դV\=o"��H_R{4*v�����/3�V�V*l࣎VY��i�ŦS��qnA��� ��q[��qg�C#��.�*���h���|z��*-7�V_c�p�oXb���z-��A��HɕÃ܉�xn1���_�7�$h��GmnH�����S��ݜ1̔�G�D��8�u�gB6j���m�Q�`�펔���c�{L��qc}g��nr�5}{C3t��j��Ȓ�o�N`��u��s�8�dL�T����j�rl}K�|�cT����̳�c�����C�hF씲�I�:�v��. ��kf�4o Vj�2��t��ǫl�qn��7/6ͮl�y�ן`��^��j��EVe������Ą������Z�t��j�S�Ըǹ@���k5Cd����d�3rv�z[���*��@K"�	�ڽ�j�|�jy��N��y�C��1�D�s)��*����j�2,�Abܺ�����^4�%���,�H�[� ٝz��kzvv.�ž�A`Ǘ�$�4��R�3r��쳍��$�oiVN5ٮ�բ��4�)��־2�f}�Z4u�����C�y�˼�P5���Ѧ2��&��}��)_r����մ�b,�^�>��W�� Kw"��jA�;�.�e������b)T#����n͏�V�U�1�K��y>1K�g�(�YJ�w��dD(� ���.�KX�P/��S��_R�0^��؂Uz�Hq2I�Ub᜶�/@,��a�Y,�[۷��y�Q���+ccO/�:�:��4���;B<[�֗�x����L|*^*p�ݺ6�u�4��t��Mޤ�\�ݴB1�z�����*Dw֮R���`������9Dޝ<h��S�wFrB�wVG<5c��^nW���{u���ˤ�E:�d�j=��ݗ�}����s���� V��V�5���oZ����\`+�ˮ&5ֿ�픠�1܀e^����Wmҵ*\C"��B�du���b�]M�s^�%�����V�B��L�5�g&K�iسq�j��r�����ʚ�Ͳ���2�h�5h��j����NPE��x��l[J�=c8`�� �WgP<V� I�V)�:y��t�!�yvfX|����WM�y�n�N����f��v�B�G:�l��,]�mg]���7-��
A�nU��WJT)�����B��B�5�~�����qmpgGR��u���c�Ĺ��h��]�5�"�5I�^�8��0�;W��S�9�eCm���+�YF�}���q^}��r)8�-um��^�ڳ�O�>�|��c�\_MM#s�܋��S�>�;�@�>�P�Z܊$Ҭ�¥��эV�h�)l��L�Se!�L�є���*�kN�Z��6�Q�ro�����l�R��9'p�ʾ�]��k�2�K��J�Q�����%["��_>�Q�T%��,i<=M�>���؃!�b�e��eX���U��%�'T�JB�5w��̀������}܌����2D�κP�p`u�75Ne��ԉ���x2��*�zjnJTu0��)o������X��K2���*V�Lѷ�gg+\.Ç��K�lR� [�G��utiH]��v|�ozQ��l���R�ʢ�g_T�}rwygvn��_9n�
���t:5����p��}Y:q�3�ˏ.k�, *�w��u:Z�]"1b�X8_��[�t���Ϭp��]�&qR�<�|�U��rcT����Ԭ"�Wb���� Z�е*u��l��ŃcM)�Z��|Z�S��goR�f�Yr�l��-��D�o��$VM��]]��߭�:�/xT���V-���(!����u�9��!췈��l�S�O@�{�n�2E�
�F�8�͚�K��:"
���X��%�ʊd�̽OCe6�����{�W����U�٪K�s�G[���Ul��Ng��+*�$r������R�Ծy�;/T{�L[�O;��gl��5tb�Cv���uì���[�L���o{����KroT:���!w�I�$�+��mpb�m�A�SI������{ٴ�n�6�^���d!,4�p����..ƸEڄX3��F�W��;��v��yR+�\��(7@�SThehwP]C�:�D���N��=�;{�����ī�]_*��[�o�f�9� ������c��ѿe���ζ����6�iȰH+	}�[0������m�t*gV��m�ͱ)�V�ϗBD���{$k�䬗C\AZʻJ�];ֹ��1䰔�j�C�Ay[�JEf��e�����h��P�$z�θ)Aӵ�Y��R)u�#�{�t���w[���k/��I�<��p�[�$'�ԨE�h��>�)�B�s�}JԬ�dҭ�:�e+�Jk�O�1���6^.�r1te�!�Θ�+�㷡f̓;���M�VU+�g8Н,�+8�a� ��o��vi��-�@�Z��nb���d-���q�ֳGωu���eu��xR����Z77�C%F{ճ���u�n��3�&�:P;-v���<_jq �`���K�H��V�8a��ʲT�¨��W�\|y͡[6��'5-��3�T��t�IR�A�m;8K�*X���r�7Zt�m��Y9A�ߝ<�@�P���8=<(澚�qkj�p��9y��R�${;q�Z��y��,>��������,��SoV�T�N(;79Ղ����F�>a����)qή��2[�F�}MJ�B�<ytB0f��P�eݎo(2�v�Ժ��vi�gFA�ʃ!<}�yb%0�1ܼ�}9���_8�����+9��84�b�z�NN��Ύ��\:�R�9�F�ug,�
��pnt��Y�|��X�S�7ŽL��A�݃V�ճ��屖��\�Ӫ�<W�ۖ�s��V�:����Ol2�ٵڷ��7}�!�w7G��Z����ȃ���on���	�n �]�@�����3�]m�5�������E��|��ݰ��[�|Y�]E�'xa����)�	!�v��mVVӲ�Y�,]%��m�x�����Z�$8�Żцhd�Q�8���ش�Z�{�VӾ�ɓ��m���_@[�w�a���[�)v��|徥\O�[����r�\B\޳�\�$�P҉!��)E�וK%�:�v�_k.�z+Eů^l�7C<{/�n�nQ�3�	��H�eu���#5�ګ�(�5��5��a����K��`DM���2&k{�	��tM��6��kѸ���	��i�j���F�:��(U�lǫOZ�"�iG�3ɻcV�+���ݮ�b^QY��%EWk��Yw}��[*�ܨ;P΄v��i˻AC[ܟp�܌�0b�0wS�1Na|���s�;�[��伵R�����M�7����נZ8{O*�2�4��qf����
Mwݮ6��(6�PLs�/��G��;K�m��k&�sI��δ�0�pQ�x������{ka:�:]m�����E�r�y{�%�u����,U���:{�L&����\�i��v�v"�T��#�̋f��`�mą9w++df���M���n��
���լm������ヂ���������
bS� �+�=I�������t(����e���+ܰ�����t���n�� C��Eө�b����7{��+���V2������Ҵgs�m�܄ir�4�a�>�cb���nY���r��ʽwCE#��ڦ��2��!s�vkGi��S}#-���:�W˪��J�Y��ԑ|�H�pf�u�!��U�`h���P�+��V�d������j�[���ř�Pi�WjO��g!�%���-�.�����b���b�WB�'��j���x6��V��77EZ��&��
�2�k �0s�������Bk�n���ٓ��݅'~���qx�d8�ډP���ދuf��o'4%�%��y#j�I�)�:�`S�nMQ�R]˸L��v���|�Z�ñb�[���m�Ls��30�&^�|�۠��=��mwU\���:V�V�cEu�����v}�[�V�a��ķI��{H��q����ନ�!����@-1*L��C��Z�隶sX��8)�;ki�R��X%m5ڗwPc�lF�.�T��E�Nһ �{{��cF��	����ğ��u�E[ytK ;�<��\�{�:1��^�Έ��KO�k0P�j�+�T���BB�G���{4_E��4hڹ1]��ETv�7"�1��r�SG+,�|��r=jE�s�s��}Yu5����m��Y��j�I��0r��^��\\��5J�˕Jts0WX��v��`4�+wu��_R|�է�b+�[�x ���2�Ni�����uB��� C� P;�KI����rd�Z!��y��E�ܺ�ά;`F5����Y�2E��8��v�&�[�O:��,�[��V�
��!VpU3�eES`3
��#�}l��G�O\2�(&���qO��W�ocԀ��ݨ�;q���P�\k�?�s�7B�f+����	s����C�3���:��f�u�a�!&��i.��f��殾޽��\�)0��������w�]dX·�0��uD�έG�չZ\�ˣa�UŠl����Y}M�롈��p���汜�j�.�E�
v,�s����_4����Cx�<�I���3���I�dss�,NF�\�
'�M��9�엄:�9�;�5}����}J�R�r�{Y��Y����N�d.f���+��YotRX�U�W�����.��Ա&m���Ӄ��G}�ʱנN�{w) �T#1�4��M�Y������(r<�;:�Z���u��-RL�-]M��]��H=[�*���k���ld���
�����6��.��x��ⶵ���өu�T�w�qAI��u�]	�n��Sp�Yu�;q�:�(�ҙ�%M�X�jN�bh^_L�q�&]<pI�*�bW;|2�C[�{�� Իc��S9�҉��0]���^�bQ�K�j G�b��,k^G7�;f��&�����=����d�+�ZY��sq��Ŋ�7E��2x���
3�I��ؕ�h�ε^w]�p�\rs����pQ��v�3 nVG˭ �&�-FӰ���ps�i���xRªU���]ף�y�N�������mΉB���\�Э�-�;��+si�r!�\G�S���SAv0+�Ws2ݧ٠
*J�
�o+��P���a��@��j��v��Q-v�u"o�A�6�sv�)�+���N�_-t˓5��q���]����<9�]nq��%��i"��T�u`��GqM�wu��4	��|�e���]��Y����s���y�]���kk5��f�+�[(����b���B�w]�A�P'����c�V�P����,�4:�c,�1Jc��*�Ps̪|��m�.]��m+2t�9\]�\�2�.,���Y��z��{��
�I�D��u��wEe9]L�蜾S�n���h5�;��_R�㺰��:Ԣ�+�s	v��'�G�[�p�жΙ�O��
t%��.,��Q�pe���g~�¹���2'�(B��F�o�[/�N�8�Ԗ�ro����YŔ���{�f�vs�ƧuH�^��]�9�r4�����D��܅��Hv)�)]��}�	V�"�T:g5PW-5u�+5��t�v�\�	Vo�B�̭�Er[�p�d����,Qê}�R�;����O8 5���ou�R�r��Xr)�1�(,V�A�z�qZ��P�Ƹ!���\罶�-oG[s����c���:�|�V+	 � 'u�(	ۯ	�J���t����Ǆ��{Q�͞N
���Ŗ�եnm]��M"��}���;ـ�sx%��&�=>�����ѻ�mRKys�iP���.��ڽu9+��w@rF���m\�3]�S\���v�wM��4�2�v�DHJ���^�˻��5��.̊����㿖V��n�[ÉrG�9�aZ��D���ڈ�u��Lխ��ž����uK6���%ZE�	�z˚�wZoW5øa�3�-mN���S��f�
�v�|*�f��oq��!��;��X��6�/��>�4gu�678.d��Mq�԰M��>�9��|j���d��9�,Y��pw#1�@=�wZ�.����9�(J�]�ПM�q�[C�Z�]J�]�7l�*�(�V�e�����#�	�t5�K��V�8��mУ�J�`�n�	ii�-��{,0�^��mGQc#Y�jά�rS�6h��$Ƌ/Xϛ 믪��#����U�;�F2�ط ]B��C���"�ܬ)6���jS�3��KK�����We���x�x�N�o�/[�|�Fh�Vlہ5)��Ά�b\m+��V��۰���|�y=?]\ �� ����--�uc���<h4$����o�
[w�p�9���̲U��:x�<'�${R�l���[L�v`���|�aw}V��c(l�$�@�T���m[���#�:��륚4�����e%��V�X��c�ʂ^��8��;}�rw8R�J�U^��T}�t����!N��w-Yʮ�Ԓn��
�w9�R�J���O4���P�<�C���r�X�>��fJ	�u
�س��\��
:�,���­ܳ�a�3P[BW��Y*13�9�"ͧ	�ݸ6_S�k�@�D.��.�(��{c���^֓a*W=4�}�3fૅk��+y$v���2BY}��U0O���^��kGe��Ү��B�-y�c���җt�vŻf���#q��|�٭ ��b��a�{�J���8�B�A���XUm���x+��XYzU��9ON_V��]���:�痺���/N�5#5��EY��rs+��R�bb�uBZ�`��es�2�n7�/֬��Z�"�l�}��S�՞�:S�G+��	Rl,���\��{��iN��=��T�.�_K1+�-�s��f0B�;V��ހB����޼�}S�5ݛ�b�����X�yG�EQ��8��/D�E�D]K�Wq"�ڵ̼��p�u�!���U���DʵJ��2�t(��^����N�;��䞋�9�%E�$����:��;�����'���t%Y�J&+43�VUJ�����Gwp�
 �r,ٻ�ZS�99]*s�r�2)#s�G8�)����*��fkt�W2��S=�;��S���Ij��9����*e'�yvII*����N��E�2rB�y�G����r����맮y���Q#<�C0��r=�e�I�D����7]r\B��%B���]G���г�U*)3SC����VY��zi��9�wj��^T�Jn���9(�Q�r0�]����$��YRgM�ba
N;��E��^���9$W�z�^��|��G�~L&��SS�Y���\�Y�W��e0r�����W�"�Ӻ��[�u,s5���+J{w��}ojI�{zT�.��B����F[u�r$j���T��@��\5��񛋽{I�0p�e��a�-^']�af�>��(s�{����R�?Oq�f�,Ӛ���Ǉ�|���uC!��cD���b��k��v�V��m)�m΋�YC�s�Z*Qq�j�D�'Uõ:����HŃf��c �d�M��q���ثZ�ɝ?8��������J�B:�Gs���vuo�s:u1��o8��PUzڪ�u��*��T� ��/��d*�_�K���+��M����z4�y��:���Y*�����N�3��4C��ɜR��ݏ�d��r��߭��0y��q��Oe��CBNW��'���YFp�J����^��p�����B��\����-�p�q�+|jy����,�&�i�I�Ip
���R�1ъ`2���R�T��ZWؕ#�\nm��R|sO�m|������@���:��-�JD�|dY��m0a��J���z����%�jƵy�ӧ�Ӻ��}kk���z]�2#xQ��л��-�݊�
�N��{��N�*����a���QU�*�	lܠ4��z7z�
X�|�-�fօ�r����]O���=
�ꞥKeb��s9�F�V�Ȧ��P[<0[Z�#��F�pX���0�u@�<j;�C����XBح�s�r�D8���Jr��j�A����q7�A�_	g앨M��S{�����|(m��,������G\���F��pF��ա��D��H�نx�� 5w(���G@y{rA�!�����"~�}F��#�ʾaF�j2�J�ɮws7���Dʐr��G�-��L�ѱ*�I��A��x��ۋx�8�/M��3m�ӎC��_n3+��͘��d�&�n@�޹�5	:k��
�s���W�D5�5�NwD%���Ta���m��:57b�#'�!��tT�m
�oX�8���*zgb�1Ԧr����j(K���pJ��c�7e�{401|��0����?�;p1��Bz�o�+"��#��ZC�8���1�U��gA��@�u_ȱ����ֳ���<�2�,��JR��{�e��'��w,�Y n�x���}QՕ.fS%~�i�F$O`�RWs�G���kώe���`���\{����`���dA�g��I�;�nwf,AN����J�'��kU��1��vd;.�H�z|]�����e�V��Hkw��X.�e�v��j��īGk��뻝ڤ^��0���SN�$ݗO���d	#�tW�F�f���il�o6J�����[D0����wFx�4z6] ��7��NrtݖC��o���ܞ��a���\9��c��у'"M��%������J;BL�T\���{ךD>�ƕL��f�=˸�n��c���v0��9q�k�I�ٱ#��;�#+h{N�M�c�,�R��j#S�>��������C�3l�H�b�M�ܼӑ�\�8[d�̰$�d_�3��qM�	��cW-
�LC^�aYr�n8g�l�W�����F>L 	N���Vd_p�鵃��w�㾁��ק�17^D�^��0�U�j\Ԏ��
C��{�i��<����gޭ4T���Z���n�Gy�W�V\���9X��V��3P���a4g�tT�Z�81�y�<Z&�)Nّ���;���w��W�>S���+��uƆE*�O��x}4�M\"8��p����R�貰È�+N�2��
��;4m���>� X�
%��tx:��K@�fO!�
�^�tm�.[��]kC����	N�Y0�s>��ǲ
ƺ�����d�@�}�p���uqr�d$&�q�qL��w;�n^eY칉���ˡL�T�e�"#�7�v뺰orYWou@==S��㺚������]W�20b��^R�:�!?T���4dm:zhhc;U��$� ��i�	���GI�Qw�|�q��,x���T�����H*ޔ!�Gu���Y,\s�b/官�Ι���D���o�A�i�����v�����|�K�mGi�Bkv��7�����˪m��έ�SD���<�B��ٗ�_4n����^���0E�KPvQ��t��L(��OiWk~�<���3�K��ZC�+/k@*��'G[U�mj�.�z���#f��p��boh��w�N���wY��:ޤl:�C��l�\i�b+��X8�<'�f)�1b�����*��O��
.U��tc�f�����,.�������*�:B.!�l�D;�\a���`�	�*�Ut�1ֺ�UC@W���
��7��ꡃ�q)]�YŻџk��2��n;�`��y�[=cd#.��ɯM��k���c�~ay�3��s����O��=7c�8��K�u�/�ޤ�%�Y�*y���2�Q������\���\�G�xS�]Í.�n9��
V���h��v����x���1��[o"��hSov;MZ0!��B��ܮ�ѓ/�;j�Z*��L�I��dc��f�W9.�>�q�N�K(�i���Hn��
��JX�KZ�Z����Ƕ�q���m�\�]���@Q�f�n�`_V��/��n,�u�gq���9	������ E*�:5��!.���UŹ�4-�i?zv�����pj������,�7�jv��LTy�#D����4�D��;���$�t�qBSTA�h?���7����u��mQe��V��1
UHF2��LS�&��y�K	4�L��.�deN��u�ъ��H;�֮C��9�d��偬���f��[�[�Q��ƀ��a�M�yQQ����Q�2Wѻp�Tj{ld6���
�c�Lų��)N��,@��%�:����/�x�`��Y�̞���ػ�E#:�=hĩ{�m����׊�h�kz�.t�1�~͇uB����0�1 �\�>�=e9Y����W=�c��*��Qr���ۿ��3J�W2���^�6��k-���i6�^v�ҀZ�����Roa�R:4��_R�� r���qȆ��wNq��yS�gm4kS�8y�Fyshv@nŉ�G2�u�^��t�b��fGD+ޟ<����f=Vw\!lTe��*N�"*�|�=���k��N�VW'��{�����Eٗ����4(�I�RJǽ۵��G��֪[ٽ37j��tM:V!؈�$Rk�{V`�@mګ�X%sW�β�(�����yu=�h�;�tY�5�)�C�&pw�R�% ~��腥���Z��#��O���O-�Yuw�E�wh�ʘE���weZB��_���o�[��r.$�R;���󥊼OO��@�u}�W8�>�p�'�i#NO=9 ������w�r������6LO	;S(}(��B�w�FP{�D[�G7�ݧ��K��hO%OO}�C/�i��y�H����־��eU��|�j�z�k*jsL�8��V���|h�x`kn���k��+ܛ]�<����Q��e����oZ�!�C�I�-��
xE}�������e�븛��������\��=���ʓ�0ʀ@�P'	����6*������3}�@�ZM�a��d���8�[=�]h���;ǆ�n^g=�G�C���
l��ugܯ�+�h�g���x������ݤo�d��H�0�F�©Rf����L����m謃C��-�kK
�8��Ab�I�Y�R9���.���NpA;����2��4�����R�hg���{K[rz���_*~u�1���g�����Nՙn�0h�V^����e7�p�Y���i��b�m�U�S��tM���Y%l��2��!:��gGR�J�����ȮT��f��>L��A꾮i��o�ovuۙ:c�]���mǼsN�Ȫ5�Bs鬑Ƞ�R�\��O�uW
q�N�����'�/L��!�=��kڴ;�0��]��t��7���l��P;��][G����&8mL�Â���(;١��r��MU!]y���n-K���aY�����S�i�`]Ƚ��Ch�u��O�']�7C1��D'Z�h��Wh��4ְ��TY�Q�rɩ�f�W!�Cݿl���IL��C O��<��U�F��|i3���6Y���uv�ł�G�F�9*(|N����%&�+�e��i$�O�'N�_%)����c��Wy��hSFĩȓJ��t�������%��\��禦2n;���%_+�.�!�ʳ�ܶV|���"t�t�ȃ��<&�d�u3�8�eo��z��)S(�ѝ�Y��Sjv������M\>ȃ6�ԧUkټuq���sx�
Ѝ0�'*�'�{�Ⱦ����+�.��.%K-���c�8zjkW0)�Ι��ҥ���i�m������� ��U��1̬�����Ė�8,صa�%�5%�f++�rRF~���c�MW�z0S��;��rL]^��n��'����{�n���yG��;�h�+40Q}�]�3��w���oE�Ǎ���[h^�7.q���->]}n�˧> qa��B�5æR��.��vv��ҥԞ嬆�z�/�c�ݼ8� 
�T��}�'�X !��|R��i��<�^|���� �������gQ_;ݤ�:!��r��j�
�2�`�Qt�;�o퉦^��N��tΣ߯���-�t>�i9�ŗ6�x� ��4�dTB04�c��B�Bd���c�r�9����H����1��=�Hv�I�iѣ��F��i�c�0	9ߵ�Ou�پ�|��N*TI�6~�Y����2#iS�YCZ��B�wt`)�NdHj�x"d�V�#��Z>�L���΅��f�s�s�Bg��ƈɹcb9U1
��}�c��Pott�˰dФ����_q�thS����7�f*��{���X�z���l�q�����{���7�`p&N���捵u��ѱޘ"�#����B�?���ܘFݘM���Vl�߻Z��;��{3?ZJ�
e2�p(b,��~�bc�h�j�� ��*��"C�\/BY�|�����,gG��c�^/0;�#c��X8�=�����1Xl!]w��,U�����9�V7����_v�r�<�,� c�v2�75�&��;�uu��m>�b�^	�KvUٛY$�Ϙ�skq�'}����2�f���c�%hѱ�VY5�w���٫�.�+H�yO+�s�g�����&��A<{��ȶ�A��p�B���}N��:)�,迅IB*u�#K�4��
����gT;� �q��]wU75{�N�^�mq�����
��bZ��>�ʨB�����q0�3y)"�`�Es�{w��˟e�-��Q�a�l	��k���Ó�hx�y���iydK0���I#.l	������5���ۿJN�) >�� a��0�Z����q�ܬ��Wֱ.��	�U�e��e�1�q96��.��3_t�"\���v�~�ڴf�L�a�����t����[����w�f.ۃ�`���T-M���Ğ�Fҵ�B����&O.��Z�cs�e��~���[VY)�!��<�SI�$d+��J����\�8�%[�٧V�#>v��9��zg�Hbឣ�G5L�#r��¶�����3`m��@�5Q��8�C��ERWV��0�J�ۄ"�=�I��E���]\�r��UU���7,hj�:?�&x	�c�cB�p�� P�p���ώ����;� ܩ��6��}�̩�[y�>�<y];�����m�%�u�l�:���{�'���C^�iNP�*۫���rau�S���m�b�)�8���<��!�M9�e>�s�|ں\,3��u�r����&��e��c���1sy�:�'����ǌv+�Μ�7w�:Ҝ�m����P�ҲU�\+�|b�g�gɛet��ٚ�כ��>tT_�q�˞�h7Q����=<Mj��7�o�p�ML<���1�#O=�f�������`������n5��:uC�h��uc�>��5�E����y���f�Rv���yu�P��ʽ9*�b��_9L��V��.]6t�2�햅G.�9}��5��v�֏��J�=WP��I�����n�k���K>����$fs��^D��`.�}�:v���¶/=b�m�&T\I���j���va��	枩�l[/Mtu>�jVt^=������1p�Sjtwd��	;Q2��Ҁ}�c����ݿ�*���r�o%]�����_jV��9�9~Cju�M����m<ߚ.{U/��u'����4��fўG��U��Su��6�i�#J����!���J���]X�E;k�ŧ�`���rai"�g���tGF'\4�D:��:�$G��m����Q�L���I+�&���b�Λ�!L��l��m�c�wems���Ɖx��M�8���u9�Z-,�Z���РsU�,O�(��X�� Քľ#�y�bA�CUrFl��y��	�Y/E�
$S�֎ҹ�	(u�-�ݑ�٩mK=��ڸ��n�}��Dt�B�2Rʰ���i��Kk������B���e��Z����w]q&�>Ȁ�[���z���s�ND*>O� ��R�W� f:�Qu}�Z�d�{�?ak�K�q��_)1�u�us�r`cQ<��o�)�e���ΒAj�
��ۗ)���FPu�X��B�i���d�p��.Ɖ|��Nmb���Ŗ���K�ݼWo�$}�luY��
��M�h8�[�F�l6�E�������U��Tn�n���T6��C�h��K��<��N��2���̏�I\��*ɍ:}ݹ�a���Z�K��	��b��<�:���T�i�*օԬƬ8��k���A�Ӡb�[��ww���\�j�y٨��ϕNr���T{kEK��a �TL��cw�'g-0b�n��I���"�}�)�q�㷣��G�s2�ս���kk(nL�  K��2�u������ )p(�����ٓ��} n��.8ղ�f�o]nv݁Y��P����{�d㡹��i��(��ic���WF�m&+ye�M&f���`l��"wNwm[n�nb+s*� �,]�cqU��5�j��7ļڜU�S��A���PacInb�.�IL(�{�Ȫ]�;�ܹ�]��[��2u���L�uw���o����J����w��m�ݦoYd#�t A�]`����9`���yu5���&�.��ѽX��N�ue�t ����uE5(���5����2��t�	��,w��f]uԋ���.�)޹˪��+�e=]�����j� ��J98or,ڃ7Kй���+���[=�i=�X�o9�����/;M,�R�.Xd�Qw����b����'s��`Fl�ffVL���m&�ٛ�D�x.IWt$nc3��VI� �v�O|�=e	Q;Z됃HN��N�Mc�2�P��'�cQ�3)��bf9Np�j�M��Ye��Cd�0��.�ܹ;_>?<q��s9��]v��i���V�{��S��ů,5RTu��}�:�39��;Yg++�i]�Wgu�N��:�iާ{`l�{/�t�[Ʀ>q��5p�34Ve���1V���#�w
X�;;�[{[]�jS\U0�"�����m�t<z���\nt��4�t}��5\'���JU��U��_k���x�]1wGX�#ô\6���Yt���`D1��9�=�^���n�2�yu�2f�k���0�D�.�k����j��3��ob�$�L떔��F=Ǧ�gF��۵�ew.�qw^����f�:�p����ڶ�3�Y�"@]�zP�t��9Q�n���c�$�0�绂���̌ʪ6�ȖH�D�y�t�C��c�Q�V���Vf�i)��KJH�����s�ݦ�I�3�2�,�z	NZ�-�R�����a��7Nr���D$Т�R�fY%%j��<p�@���Ij*�UmMZ����F&��p�S�,������s"�.�*%�P�.F*��t��+'nD�##�V��a�V&)�rH�R���H�D�UiI�Y�J*If"�-+0�%D�M)T�)ZAXHU�V�R*�f�T.�-�]%R貫R+�D�XZQ�&e�͚�ZTSJ �H�(�D�-�%KD�l�NgQ�) ���BR����Z�Yâ$V����j)D����\�Wu�,2�ZUmP�CZ��-C�Bf��2�<000��K)͊+*�����c�'��Ѯ˫���pGuC��CA/%5s�:g���ve�a�䭓�E�ˉZK+�o5�̥�/w�������p��90����}C��<�u�����<>ݹ90�<G���~F�!��7�O������xL?���翾�.�i�I�}����_N��DF�{��S8��s�M�ѝ>ĸz4Dk�ۓ�7���)�!?��;������V����yC�i�u�7�r��<r��~�̞ݻ����n<'��S�z��þ��������zM ��|A�
�t9��o\]1y�O{5���DE�1�B(}􏾸~����[�g��7�'N��?>�roHN<}����os�!�� }y��t�&�����t|q�\��w��Һ�u�"��r�����>���;b��>���r���X9�P��wx���U���x<&������w���!�ϗn}vߓˉğ���Ϥސ����/�nNM����~���<'��}��b�S>�|��:=��;}�c��N��&���]�����W�{���]�����{�eߓ<�����=&}q�������ra|��E��}���o#�?�������s����}���h��"$@66@��>}��}�~�����NW;HS�����o���'��~C��ۓ���}�	��?��{���F'~v�|���ߟ����ӽ�����Y˾��=���1�.������it���/�����bG��q�<&�NC�i��r!���	�]�Ǌ�����~ǯx�'�nC��S����!���S}Bt�|=�~���������m�����?P��MX�Pp}�s�ws���=�1�O8]�|�Ǉyv�{Oi�Ǿ��
�]�վ'��רޏ�xw�9܇�=�Ʌ�P��������®�|���S{BM�}��N~��?0G�G�DLx�.���U���W���!!��7��m�97>�x��뷴����뷔�	���xw�iǧ���ù]��1ɾ��M�������S<�'G�{O)����~O.<�P��.�N��"E	ɽ��-<�� >�#���>x���1;�������v��o??v�￭��o�����&O�������$��=���<��;Nޟi������v���7�<<��ʓ���������i�?@5c�Fo8Q2ӢŬ!B�������|���J�4V��$;�v���r=lX��Ş�}��;��茻��"w+=pf`}��A�]�k\6	2�S�޽7�'����1nJ��g$;�1L�ɨЫ��(�� %���OJݒ��I`��Ap�?{�ǟ6�_)�������.�Ss9w����yL)��ǻ������X=w�'��S'>��݃ÿ'��S���?!�0��ӗÏhs��A&^O�܋y�{x�:K��$�\(>������?�zw�����nս��x���=����VJ��>�{#S3C��;C^�{������S|M�ޏ��������>;o�{Fn��~;���k۽/<G�}�"D|)���ohHx=�N!�u� }I��ƻ���ߟ	�!'��8�o��=}�HyL=~v������w�i�]��:w�i��}������]ɻ�{z}�TΪ�x���(G�>�">b0D���M�����~O)��_E��㟨ro4
���n�?\��__���ݹ9[�����n���ӟ�G��}��ꏐ��@�, �3>��e�]\��$���}@�}�G�T��-=�~y��{?~��o�O�nN���&��I��c�y����w�<x���xC���N�o��S�P�t}�b,}��:f"��BD�����B�<��0��u�9wo�G��CD��]Q �P�~�����\}C�����Ǹ$��?;w���������G�����ohN����rz�|��|�G�j�>�1#��>���P��8�Y>����z��y��S?�
C����W쉊��~NC�k��v���r�}��rraw�~}��zw�yC����	�!&������x����O��c��N$��O��	�!z��9���;��o��U9X� �ö�	/|�B�:"=A?}O.�v�<��x<��];ô���c���۹���ro��y7���<F'}M����']�90�w��}q�=8����߸�P���[��`�����
�ʘ�L�׍G�|��}"$G��s�u�|�濐�]�%n���|��~�>;zW{v�����}O)�����۽�$ߐ�n�}�����S}B}o�x��z����{������<!�?i__e��q���͔��Ch��#�G����L/��c�<�õ�&�~Nq��Ǻ�O	��S�W�=��L)�;��y�!�?�z�x��'��>q��N���;zv�����~>|�쩉��\[{�`���<�������.����j�ô�M6�(�2n���tr��kPdm@�"��ף�b��%�{k��9J�(���n��Yv�T9#��&wS��w#�{ΈL�M�΂����G�:�{������G�����V������u�>�>��Dx1�'��˴���Ͻ�p�ô��q�='�J��?���S���p����~w'��h{O)��^�o�yw�}C��緅q�	7��G�ߏ���߾��3{kG���1�#ڲ����8�/<c���7��o	�}�ǔ¿���z߾�7�<��zq�<���M�?'���\{NM���;��vM�ނQ�*�������؈?Q�D<e��������ϗ��9��<�����s�~������]�P�����=?�m���o.��M��nN�<bw��n�����zL*���?�{C�<���Nܣ�|o�1�"G�h����F�1c��n/��^)�^��#�`�=�1B(�
o�y>��/�oI���㷊���<!�ߏ��Ӵ�����<eߝ�@�|��}�;������ߓ�O��;�o�">�>�!��F�"$G�6nuP̒<7�6�B�����|��P����E���	2�O���x@���8R�{v��P��s�~��g�}��������~���.�����˅���|��݅?'�\J�ߣro��9n���ϟ���6,՚����}l��G�"�$DX��raOo�=;ü;��ˉ\HI���a��G>ݼ |I�?�Ï	������]ސ�
���x����7�a���^����ڟ����%j�E���U����������S�����������4����z���+�M���}x����+�/8�|Nv���\rs�~�y0���}��|C��
��{�������}��uCS������R�fj,��	��W�{��ߏ�M�L*��]���ސ���A�}v�w��߸�$�]���?{�㷔��n�o�yO*�S}��ϗnN�`󏗇N�m���ψ��çi&��x}� Gݾ[��#��vd�v%��?���1>C��.>�>�}#oި��zL.�x��|C�����xW~M?{C����c��}�������;Ӽ��x�o�ܛ�|Nw;]N�}?@>�@��3��[���~�;��p�x�yC��M��~~�\.I�����~Nq�į����{O��y�������N��}�������u������r~��xW�N<���xL=�<�b�Xc�DE4�c�yꌋ����pZ	�Z��K��6����u��9�(�%¾O9Z���#��͡�lLʐ"�.��o�;�Mv>��g2u]_>����c5�{��Kw��42�vQ�Τ&%]��3�_;�ˠS�	9z���}�	�"�������]g?ɿ����	��)�97! z<G~��|O��>��]���;~t�o�7&�������<nW�ۼ���Ǥߐ��$����&��q�������.���D�)���猗�`��{�}��vQ���{C���V���þ����.����l)�#zC��������������>�r�˾{����I�������ߐ�����o)��P����7�-wxe�zVʴ�z4D`������{��ߝ������(zM:v���~|9w;J���M���{C�n���=��[����<�y?���|q�>!�q����]�4�q�={�Ǥ�� �����f�c������L�B}�"9'~�~}�V��ɽk����N��@�w�ߐ�������C˽;Hy��O8\.����~NNq�%r��S�ry:?�x���=�q�ސ��!>�T���dri{����]���h��w;㾡��|��ǅq�	����	��o�����v�������O����{�zC�
����I�7�$�Opw����xw�oAҁ�!���u�����dU�^n�ƞ�s3]}��_߷�xW��tzy7�/Q�ǟ�|o��<��9?�|�<;���=o��x���®�{�P���s��}������M���|�������{���ohr��r`��&>�"����)�NK�����������o�(�Oh.�y���on��缿�ޓ���P|B~�rw�=��o.��V���w���ӧk��>���ߝ�}�<���`�{O߬D������u�����r�7��Y��s�~<�����]�'�)��s�|��t��y�	�������O�����}[۷!�����];_�ǯ��S~Bpx����?c~C���O�c�<,} } |Dn����e��!ˣ���?���X�CH�@� ��E�,�������.V�>�|/K��ҫ��o9�ݣ͏�]C�YOֲ�ôcM�������Q����l�\X�쬹��-+@��Ccֆ�o��T�8hZ�=�(�1�M��{ �y�ޱw��q�[�qwe��k�h��e�N�uHk��L r姪�ٙڐ�d���cr죓J<6��:��bS�h���n�<���yn>IJB��i��T��h'���)V˷|3�k�U��}�S(�����V�#&�T�ez�s�WCw��r���x�5������ޥΖ´=-kS7ˀڝ����	�ԭ��C/K�O�mCθ����0:�R�ϑ$��{��WW%��i��-��1Uk9�7_����v��r4����:2{,Q�TYxi��J��
��l�����L-$Tl�5;�<#�;�m\C��2��RPԍ�xSFznr ��G�<>�*�� w:���T��Y��V�e�Y���D`aI�+�z苍���A͛ݩ�Zw�U}=a�S�L_�ņMCS�R�rB����q��y�[q׹�1��p5�ճ����?py�j2Ҩri7\��4!CJ�5(�� ����0i�87x������ѿ���q�_�����&�&�n��$�zE�	#w��7(ԮT̽��bu[a�m.�+#f�Uu	'U�C���뇵BY�j�S;���Z�t�1����p��8{�4!v���:J�f��ZMnb��(Xcy��cb�B૭�*g�������@m^.��/iRz6*̱�QyKIz�{&pr�����"�}wI;�<5c�Mu��`Ra��z������F��~���U�V�P�:ˎc��h;����R�K+��Y5��r���ιj���W�pa� �-�>).w��u,� ��hg؆��G�}��"�:�˭�١#ݕ
����E�L�P�$�c>���'^�ez�أ�;����5��lg���O�T=�WK�ГĶ-�d��=������Oy02�f�&�uK�����B뢯x����)�碥m��Ѧ��F�9�cڞ쩝�1Ioy'a{�����F�eP
�e�_s��퇗�u�M��Բ��V�`���[ӆ�m[qʖ�bføwT�P�UDEbu���e����l��ۿ�D�ɍ�����9��U]or:\WI���P�+k�Y�좍Ҙ�k�N���\:C2 �8�,^�x���b����t�S=EO�cB�ĝtW ����BV�]���>Mމ%K:[�0(M�;F�trט�9,������J�B�%�}�� IJ���c�Y�_pxu�Ѓ��*�Gf8��Oq^+ؓyQ��WO��'\8� 
s(Ot��V|��*�a;b��C����ԹPʽ;���j1q��r����s���8x���H�"^�����5u������^L���g��2�y(��;l��x�gl��'r9���u�ڭ�djm�X��|���3:nS�	�ՠ�T����D��۫n�����m�Æ_Jo�U_)�}�O]5�Wb�𓳧=N/�^ur%��=�%��)���_W�}���c���'
�R�ѻJf��<Lg.�G����f�/�U�L)�3"�J�ʸj�La��y𠏾)V�T<�:�U$F"��}�V��N�;��
��4�Ѹnb5�C�T:V��|t��9�8��(#�ht3��Ý#EF䵽�]Dio�q��B�wt;��x��бu���R�>� �w�?�L_�@�\O�U�>
��x]FA��{����g�K��X;͊]C�v{�V*��c�gD5����U��DL�hS����1�o�k2��õ����%wO3�S�i��̛<,$}�������j�ʎ��*":��٠9���}��Ӕsu�=x�
�0A�w�&i���|m��8)��K����Z��jĚ�fr~��ؼՙ�ܐX��q2�A?+�ڮ��*]�#e�
��1�2�ϩ�g�q���B	Rf ��3���*�FY�Q���+�`�< h�SYχ^8:���;p���a�j%o�c*��U�M�e�{��p/MvD��@_������z�����uK�A\��g���]�Wc\	�{��[ME��e��5Mx��&����ۺ�\ܖ�^�K�Z{��kB��Do)q������~����R��ߤO������ݢ��x���iw/�ܶ�-�|;�4S7LA�n\�m��{w���v�z�`��cS�U_G�V���k絝�=�tL1������o��6�	��k�������ZO|U�l��<g8��ǾР�Gv�2�� v��F�*��D�GH�����|UZ���g�)+X��=W�cx�Rj�o�c��a�1)"��Fk�AfdYb��힊�y�B�!�t���P��!�kWȔ�ޔ�&,o�L��7��KZ���:�w>3YA�zר���P�B�w�1>�μ7�������[VY��0�b�F�3�Sݰ�A]Q��Bw�l\���'��FT�rn�R1Z��֮CL�r򣓴���]���Z��N 9`kʋ �)V�'�a�}n�[훧>ث��f��f�Z���{~s�rbV�y6팄�]����',hj������ț����CnMO;h˧����{϶z;�\m�e��Lh��ʅq���@oW���Ѱ�ZW*�p� �w�F��f����	�ܵ꫙�фKY3�$wJg��}�)�zP�깕Ϊ���4��-����)��8eA�� o�'�;n	ر����X6ܚ�=���V�q3��J^#�l��r�.�׍v�{��w���Lj�G2,�Y�v"��wY���e�����EQ���3������G<�B��:���#0vQܹ3z�"�ͬO[['�����������T�査�X5C���S�A��1�9yԀ��� �t��u8�˞�n{|}����/�'k�&(Ø��U�Z2���Y5�b*U ��bo�&dU�yVH��8�.���]����}N��7
�Ȗ���B��U��E��`wx�yj�V�
p�PSVvgi����7���ܩ��Z|�xf�-�йpԞf�����"V������mV��I�D�����]=:>a[ʄ�7J���&��xq&�=)#]��	�>�u4��HW\!��f2'5+|y�������θBɴQʻeH���� Mv�k{��@�FA��Kzy�2���3�Su�����i��#J�5��t�w73�T�/0�uC�q��dI(ۂprA����<��<"��놌�m_�KbD��;�uPm9U��.
�B}��M��A�BY�c�* 	A�`󝢣�c��F�RU��UP��Y�!�.��uA8��U��[�L_�ņM58�RB��F��Vˣh�&u�۞�t{n��r�
�^���`s���lrx� NM::rf�4��!Y�&�w�Q�s[��c��L`A�P�4��I*��#��E�6��n�E�i�;Xz|��!Q�7��D�ȫX�m��2�
l�ռ�Z����A��J�ﾈ��Ӗ�}*-g�r��֌��%P��h:`��\�"��'��#�qdr�YV+�
J,����gޣ�^�����:��C���EB��M�7@swT7�Y$���y�s��ROl�3�+���7���~��]lVl�Ӫ��o�;�cO�O\=�LG�|���:�
�����+a��rʳ+�v�Uc�%^�ao-&�����f�.9��c&+��F��B/�����]��׋�~����޶��<Nd+�/����ݯ0j�aP��Å/g@[�JѴ\����U�:5���Y����鼵򪞍	*�q9����ꏹ�����C�\�wtG�:��8��-��U��H�W0�,�k'ZU�/���znLH@z̪��7i
�C=o�����\�����7�)�H�l�_Ĳɯ��e��?z�d�l�{j^Qxp+#��u/�M�a��L�{�4I�Q85��2do��U�|�9`�=e�ܶV;w�me^P�Kə�kN{4y�iB
:}O��.B��v3��2�H9��_Ѯ��k�U*�����{��El ����g�������c���E*4� T*�wf�mǬn�Wk}mmA1����_U�2��b����z�8u��f�{��2�:�uu��ZzC��m\!'Nfu�]\U�q��"1��ݣ��hK]Y|�V�\_#tZ�f��)C/%��;Ѕ9���>�]�́خ�_c4j�>7*�q�{7�[i�X�C[��9���h��{����ҷKZ���!�5Ãrh��=1>��+^}t��!�E����[�X���\��x���TX�2���K��)t8=��١VB�,��J���=]��Ak�u���w�"Z�L;�V�@��SPOk�R�Z%$��זt	]]f�kV�;���vJ�(�Ge��t]Y�����w�åpW]���t(�t�MX"�b��J콖Z�n��	7�p۔�E�+: O��F�E�f<ǄSS��VfwKZc�/O��4�U�4CMP�S9W]C�YLC������.���V#��ඝ1��r^����� vP�t�䮋��b��L�~-vl՗1�k�#z��$!�a�.�=JS<���кZ���_���q-N�[Wŀ�Nw9P图�<7u4����tVv��n�m�9g)��nu�V[,��Νo8�=���;0���!z؛D9���q��˵\oR�޴we�ٝ��b�����-f�r<���t��5�UC]kU����#�j�^ұ�-�Wh�ֱ\�mm�Z�:�1rѹw��qai�m��?Xb�1�zo�����gQW.":���kZ�ݦ������ӈ*Ʈ�+JZ��/��]�Y5�_�@�nI�jܬk�י̀m
M�9���,-l<�V3�3�� .��k����o��V��z*�A��!�ګ�Jx��+!\�z���)s���*���E��'�@����=��f��Ν�[�ͺܭ(�U�v��CEu7��#���%�/	�e����
���@2z��:�`�L�̦3���Fd�=�iJ��Zu�\-�|�r��	Z�\L�Ƙ�r]�cY�c*�1�c�L������S��	A�~.�c{,UL$`�����+�-�n�`��{ڶ����)B�W��C�<yZ��Yn�Vv���P��;̡edT�|y^�hi�u
������~�֍��̂ŀo�ځmlk�����`j-��Ө`&���q�\R�u�Z���y���H��2Suv&��o��Nm�w��](%���ާ����
6e%P�܉�w6lp���n��XV���*,+M&�;�:`�(�7I���Sw�p��x9Y��-�xz�+5�Υ��3�K���t�w1�u�X%0���4�a3�"^`�E�eؓt"/��곦��YE d'%�2��f�nled�B��M�U�j�
�k,�LVw�3�������Re)܄|��v6��a�ʵ2�,r�Ú$�W�ח��TV��"��X�X(**�6D��'���ͪ���Sf��0��T�9UV�.��*=ݨ�{����K��Y�u��F���*4�����**�S�(��u)(��"p�%�t9bf��I�Y"HXQJ̵����2�	R�e:��ܠ�(��ΊQDRr��3�Hd�H9��ETQ$%Xdm�4�2�)V�[%DD+H*�I�KA-5"J-V�I���2L��:mB����&X�G+1*�2�.��2ЍL�9j��Z�`�%
����	B6���X��2�4�Bլ�Q*���s����5V��uT���FH����:j$�êHYi��mDKU*+�rԃ�D�-��juKJDʕ
��Ȳ�,�6jYR%I���L�R�#��J4�D�V�N�)��U���D�J*��C+-K""2�$��}���y=�K����{�2����	 KISvgf�d��(e���5i�#��t�y;(]ZᓅJcg.빸{Jo��^諭�ꡜ��ܧ� ����tG�p��=�P �9�}3	U0_E7�$f�Dݽ��D��s&�����nW3�N�<�J�X�(����@	)V�pLs+6��}�<���_&l]Ѯ���>5����@K�	�&ـ.]R]2zT ���ʌ�P�ne�f�K�m)��ƙL�߄��k��t��.tCg!�VmV�JlA���:n��;��*����� :-�}R�ѻ�)����Tr�tS1�P\�%�����eEgT��x�l�iD�Lȡ�30����YN����V���+M�ju!۞&*#�vht�M�[]�a��,�AK�y���UTE0,�(�NxZ��iվ�X/�|����3W�h7�5��P{[O���9[`�z���L+��6x�eU҃c�C=�uס�^�R��ݙ7wc��Rc�'E�b/官��u^4��F�;<M��1��cK���"�E>�Z�5�D�B,Z)��A�!ꙴ���WQ9q�/Ew���W��Y; �KHi�Q�k�+
��y,�mLB� *EE��ܐވ%-�(?kg�]z'�$��32�T`3#��T�.9����v����b�:j��\�K��ܷv�f���gQ�mpҴ����8�k:�z�YBG��r��R�{�����UUO<�{~~����=(+���ӑS-��F��M�V���pW������N*��S���5��̝����*��I�{�[	}ؗ3�jU�"6] �b9�e��g��rNF��S5��]��'Ռ�}���Q��e�gJ*KS��+4���9��n��R4m�|�KV�����g��pk�]s(Ѐ#6ɐzP�ڮ�9l|�n�s��)=�ҷD[ҕ���e�:m�=&N��rx�D���]���W�G�8�.�����6���&V�T>����gc��cn1��{5����A���Ss��N��	TN��s��0�8f5x���ϩ5q72�q���c��BrkrEd9�g�U�)�9�4[ă�@�yY�䋉J���L��X��v})�f3�oJG!���Yp��>	����1750y�V�I�"Oˢ�s顟u��7!a����k�]l!s����a�{�Gxx6[c�{V�w�Zt�:]eU:����U���y�B��BkL�뒳�����x�f�z�~P���G�>O9�7�*2��ޫ̫oJY��)���FD���̜�Q�N�^F��I�Z
�	��wۖGtwX���W}��,��3H!M��;z)�+�����,�`�o�x�PT@R��K�֮�k@�1���>�}S������X�R�G�xR0~�;G�J�/ 9`k��'0DO�x�`��g�}n��ك�g�ӑ�=�U��k��1�e�m���1�6���2�',/U���zY=P�O}�v���_���^��|�o0�ʌr��L8`�y� �[����1��!�ؔ�ͣ�4F��;Rgo�V�C�Q��k����v��������u��^��<M	Y�贛�A�t?wa�{�*��պ�^��t�����&�gR�� �N����C&%M����Jd�~���#�Ͷ�&+�.Z��v�R:�kN�*�b�0P��c�s�Z�ս���S��9�y��/���d����VC�v�.��k�=m5j�\�Sr��G,�K:���h����H��)��r�is�q9_v��̵�Y�᠝�y���B�����|�ژrt@�J�9GONi���j1����n�x6U	�Min_j1��)eZ��
�ḭ#�x�!��S��١5��o�s�΋�?p�Y� ����	����C���Vv�6�O��()�m��1m>�Я�t��B\sd>>C�8�2�֮�p��q^���p�#k4�z��\(�N��FOg�AĜ�\(��ʺ�ڵ�O���*�-��V��4|c0����9�[tD!�UU��U�1
������?� ��@H��gAH�jg����-�.y���oP=0�`� �ǂ��I�}��{�E��V�/���<��H�a#	�r���E:��т�Ƃow���Oi]���[]5�{,nCu�M�u=,�3���X�i�Ό�rSc��Z{�ꑙ���1�j�+k�i��u�)6���H�b(2Z6WT��!`�,�"Qw<4���u����{�YkY��s��s��ZѨĦ���)�0�F ����W�?U�VU?n� �M��U���)V
9E���>��S9d�&��n���J������뫭Y�׺�pە�%�ܳ}��c��ޖ�dl��Q�.N��(}?9=уyL����}�����W��D�#_1V9��V9��z͉Oy�5*�J��_���������OM�K�2]OVy�1ہ���ڳ+�(����])UC�q �����ڎG*2�*�M���8 �;j8\#,�3��3�cr~�wR.�Q;�aa�-TC�C�cUi�̈́Vm����2��/�U����}%h$7��f�&a�fJ�62�\W3��̱�s��f�ެ� )�xJ� R9�^�*�s�2�g��&d��n�hON�i3��r�j�v�mcq�]X��/�����p���� {N�J{�5�ԟd�Z�en+���3y���˃<�O��}3:�Y����<��Sw��m�n݌v�-��!�zW�r��eS�y�/l�]��>*:�Ӥ�q]1��@+��Y5�2�^_�u�����(�ٵ��7!�ΕVZ�O$XzI5���A,*�7�\�ȧ�󯖇,��ea�岢v쭗{��	��
��odUz�h�Yn�Aˡk��X�+j�霋좌�jv���&{�I����<䷴GNptv�W�ͳ��폏�exZ����Ljن:*_`��j�c8�v�ηԪć����idv�^�E>�Q�Sm��H���xZ�IJ������6v���+7�xc��c���\Mķq�˺|wa:��ʯy.
jGWO��1��KP���74>q��7�2�{���b�_RN�8\��|�+jp�6 ����Y�3o����t�aۺG1��gq��8E�T�tn�)�L^�.�E3!�\�%��41ӭy �YFy���Mt̊�C�|R��C]�o�x!WǬ��Y˰���Cg�ɂ]N�=��ddX'i�fs����a�~g��&��c�]B���`�<�":�kp���YN%t��W�m��o�S�b�+�[m^��#�-�nY\�K+6�i+��Lwur�no^��M
�>5{��J���CP�| ��ݴ5u��ʻ�&~������At[���H��v�F��U��ђo�'�O�@�1QK�4dm*zk�7&-܃�ӽ��ew�޻�p�L��6i����hV��1j�g�f��yݔjzr���z���j��x�X�v���U1]k�E�����1��DVmX7<zxO\��Ɯ̌���u5��9���q�}l@�s��ں�������_F>gfęq>[���9#w�d���Y�T͔ބ�CL٘��歁��2��C���q�[76j\#���^���:�!Q�N��C*�ݳ>��jU�K��3E}�2���z���	����z��d�N3W�]�V`6X�
���F
�����|:|Ǵ�g���>�D��T''':�����\Br����pk��]�(ϡ�+�����������Oe�X0�!����p���wn���x�__2mz��w۟oO��e
�
�@�=B��7�-��4֫gb�����.��׮�2���O}�C1���Zm�2suN�s�+1����\���nt���远����j�g,�p� P3"�-�r2���]ϫ�7����L��j��]�	�h��S�C�Z}��s��
YC�L7�eN��Q�B������M<y���5d�3����Lׯ{�Z�T�J
g��[�F��ꪪ���`�og�z -O��zcDV�l��V7�DRj�n&X�,�c��@�p�{r�*ѹ9���4��ާz�ˋ�D�l�*H�J�e2�d7�.��)�f2	�)��"��`�8�R��rޫ寧6�jGyO���1����Sg:�ˮ+���>Q|p�f�wwi�l߄��tMN'���ys@=\N:	V���Wm`�2���L���r.��T��N63��ݚv�=�_���9�d��偮b�]�DR�����ս��`�}b\��r�U9�v�!��7n����ϛUtlc !I�Kŕb���OY��/���j���f�|F�� U.R-��4TnNW���\�],m���!��M��vY]!�������%¬T�P9딇���G���gx�����=(g��s(����V�S��}�NVs��
}Y���X6kK&2� �i���H��7*���u�&{\U�/)p�2����J�Ջ�]�6⪚���%��&�U�
���[�n���r�gX��aD�f�8*�s��1�����z�pQA��s�WC���.^�y��(�Iv��|���vKl��jʜ��'��*v���x��G�CZ:��c�d��q�����"�\ͬ����jqORr��m����j9D��ވ���>ʥ�5��|���V�22!Zw�.[9�R��M���Y�S����j��bI�)��Kzއ���Զ�dt��@jઇ�$8�)�����/=uJ�ۍ!wp����6���ۑ5��tp�=��Q�c�Y�J�/��on1:T�d}7Z:���P[��}Ϧ�ͽl+�L?��$��e�?����!���0��f��ڕ�9�2��ѧ�4k[�6�-��r��W:Y���6��6� !$�$t�
Zźzkb/�ܼg����sC"�e�#��U�\n��)z�\���a���u7]Q�!}H�a!�%��9p�jj*�k��E�on�Y�����P��t���8j���UUt
̞٠��|X���W�sN.��O�b��Ѹ�F��#EBMZ�D�A�Ѱ:��ap>H�et��Q�6V8�t�gCsd�3���r���_0�֍F\%P��n��� hB��UJL����h�h���6L��6�64��<�\�7/oEgƇ#�oT�<�����pA-���<1�4P�,�̎�Y@�{E�F��NP������HyCB��e a[[gP�;k� ��I���t �v�|,��ש=Hq��c��`����*E�KV��K�:�y�U���V�_���'���h�z����]C[ՙ�i׻��������\�fy9��0Œg&r0���n�O�K���ه��^\$�Wє�=�:��2\�[;�����G�x�	�!�(*�v���^����a��F$Mt�R�;ȹ�z��8vN�ڪA��}{������D����9T6�+�u�+̔���zN�����w{M*�-gQ�N��������ܟ�-�H���f�W �ӝKo�@��`������/�vc���H�@`��H�W0�7>\�׻�]��
�s<�әf��]���z�*a>�wF������Y,�k��_;����n����I��◜y�p���>��4���%��e�:�2-U�|�4�`�`2��R��6�k4ex�y��iwr�����<~��<+N
:]S�A�Ep
����n�ţ�p��*|��W���@�rt�����S�X�&�a�g�#�I�2����s"�:f#�Yb�v.|�wl�9�yk�˨:�w8H�R�k)���Q��X��6��4ovW�����2�6ߔv�ݫ&KK��A�i���m�=���[������n��b���I�m�rz��_���ym�ż7�IYc��t3LWsf����:}��2����ұ-�u��\��;��;`u)1Ϫ���{[�ܫnl�*����ҹ^����菢*�}I֖�@#�����D��q�˺��ʮ�Ѥ�*�7�:Ԏ���rK�H�:�|��Weٺ���Ps]��H<�	�x�F.5�')͈H�s���5Z
2�\�$�m�=�|
(�zQkY���E���H��
S7����]~��.�s��Sh�dxBg��v� ~�`/�?$�
l�[�5�uo�x!W�a��T�7�ԇ<r�Ú��V�ʽ��w
�Hh�� ��L�ڡޚ�H�=��X��:�ծ�V3?aeѼ��[H[�c��uv5�A��b�7wA�L��6�U�	�jZ�6�G�����ۃW��|g�#�S9�]H}nͪ�c����F���M|�H�S"/�(��+n��� !E�ӣ��t6J���D��3�g2��`��fӯ�7��b?"��x���^���!��b��k�7��T�*���,�ҽi3/N5l�T�dċG���^͸��F�d����z�&6�J��`Aε@}.6��џT�NF̰�bDeB���s�jôyS��\�|�wu�;�ݽ�SrK5�,�;t7��)�'j�"݌�S)��2��B��G.�#���u2��*��	��@���z�6�
u=!صbJw!�"�=k�+pL�`��8=�>�9{�H��Ked9�/��Zi�JW�)�֭�
�x/�ov�7 Q�J�zT�&�q@{+�u���f�h��D2���5gԨ����m�c+��Cd�2˛}����\#	��NƤuʬe�N�WZx氹�]J��7+�v��C%6+'ǭtY���`�U�r=<N�WGWQZ��WP�;���]a�A[-!�+r�裠=g�6�<�/EP�ܮ�K�^��>v�s�� �Zh]�]dNv�n��KJ�����4�V�s���o��z�S��R���I��I��X�{c�`��z�[�[mj;l�Qm^�=���ִK�5�G*�V��� �E��G;����� +�����+�]��]2����� ���E����NW�U��Q�ފnZf>@��a���tk{��1�z�=���C����W٘�ݮ��lTi��[-c���:�T5f��5�2�e���+]�*�蔨'`�)�D�M����{@Q��U��pcs��.�A��'w`K��̭@�g.��]M����	���4��4Ȟ. Њ#b�}�傯l�vּc-�ד,c������/��WK*�T��u婃X�,������QC��4��i�쫠NQ䙡Œ�":9 U��;y�ڜY3�4Ues����:��b�v��crнZ�r�=���]���ǝ�u�j�J�Y��u�m�;�0"ڎ�Zn峊�n�'�n�Lά�Lz5_�^<�X�1�vl�45s��x�kr�j���v�*��F�#k*�ڞ�Hcz=�S�i�4z뉕���C��R�/hs �U,�52����\�]�{�^�g�[������u#�G��J�ژu�:�`%]�P[0N�b�ם�����`P� yj�V%��[Yʔ
W4�ն��#k�f&��\jE����O*�p-�/�yC"��Knq5�m6c�'��pXluj׺��Zມ������X���.]�2[�i��S�S#xӲ�*�.옆2����rg<ݮ�.���Oo��j\��-�G>75���)���S�W:�
�=Z�T�薞}5G�Y9��;�4���3tQ��F�Il�	3�oV�tYY�f�Qg���Z�l���vz)8���Z��u���DtbO��M>63��'�S�B�ӻs�	��I��罯� �n2�%���Tmրv6r^sv��Ը>����&.����鎯X}���1椨����@4���09Z�#޵:��1��yk�gY����]j�1c�m�x��
���.��� �@ (��r�I5di�ըdaG*Cm1^{�ʈ��4�-N���E�aa�bUJ�D��i�%DR��Y�h��Y���H���!X�U
Zաf',�� ��*U��6�R��C@��B��e��fê�;�!A(�$�UK�W^.rx��̐悛ACB4Na�>;���x ���ڭgNif�C��!al�iY(b���-C"��N�.D�{�9i�Ze�KDBRӥe�%�"�R&��Ҋ4�Q`����8�5��;���<�f��+0�ZvA"�R��w��k$�����<w]�T�\%U��4#F\���T��<.]s��ML���U�qY�i!b�����^Z�2K=�p�tSD�ب\����NV<pxO	��u�=L�U�Gb[IQD2,2�N��9G����N�*q" ԏ����(L&�/.,JN�q�H����8;�s3��+1[��4��7�5�yt�w`;Z�^Z�S��|���}O�������_��wKf	c�^�����o�la�pЄ!�B�(D��R8��s���n���%�_ ��h�ܶy��|i����0l��3z��j�%�̤�n�+�[�Vl�N˳c�)U[��F�0��t��燦�GX�<j8�J4�����n�d��V����(
WZ��U��Qz~�)S�̆iw��w�9�l�n��EبfP^'<�ѥ�܆J� ݗ%��.a���0�W��o��������1�q99ʎ���d������({�(��v\�გ
S���)�>C8�b���)�f:.�Oy	]ؤ��E�6_�G3�}�%V)�*7�qB�R;���b!R;�LJ�μ7>FXiE\M�J�j�W.�Zu��ݾ��v��N�Ϻ<�jN�B�:��![Kq߰5�7-����7'��m&b��0�5��ų�~�j�/ 9`k����L;,4.<�}��pxQWM���99mW�k:����6wj����mMQP1��健�,���uMQ7��X��#9�ˡ���P�Fn�)Vlڵ�l%tvk�K��v��\f�k:N<��Jy}ݐe��C��6ɇg�eؗkpeutI�S�$�o�E8�e	�*��Y��R�wDB�z��4-�d6�+F�-�:IZ�S�5ok�)�c)J��UR�s�{����X��j���j��|�а���d
������muΧx�Om߷�U[#��^�Y^���:`�C���X+B1xl���d��dn�żN\��A��xZ%Wq��ĻoB�Ӭwtv�C�ݠ��0��Xx��\=P��I��莏r�� /t��3���/���A�z��G��.{�m���m/-��®�ѐ��!�C�&��3m	y��g�����h�1�O֕�d*N�
]6w)W٥�$p��ύ�6&�����UX#�O
�T��K8�����7=�n��.x1���mL��p�jIF:"�*�5y����8W�6#o�1ӚTF%w#���G�+_Cۆ�_Ε1ɪ�Q���֎bJK�󗾰@�r�f@&�}t�1x�0ّ9��o�G9�5I�X� �!^��׏�_Thl��l5�@`q�gcL�~ĕ�����7=�5��Ѝo�s�ݳL����h�9z�\�9�#�I�_( wTDI�<��,�����m��E�4Ҟ"��1bS���?�m(6��t�JZ����Cu=��h͓���_����X�w�
�\O������g5�':�<� ����'�� K�*��ı[���!��ܻ�c�)��H�Lt����|�˲�Q�qa��`�F�yF�Q����>�ﾻ�y�I�7�|�n������p졹	�q-�0Y���COP������t��^m�0�o=�ҫ��/��5�T�'�����Xd�l�j�D!w����Q�S�9�GoZ��M����-�Q��H�dG+��h�^�UMBn��0��l��íݜ���󴣮�ˋ�'�F�8�w+oEa����+��}[i��o�g��g<6�ۤ�V/�[3�����ꬹ��P��WL��N�������|^�>�O+�k�q���徥�gg\�BfN=�G�W����!�=�Y<�
���"��X�k�`��ʸ���eɥ|F��'�a��w�2Bbb�	���W��º�<���=��d�v>򰐮��b���v�,.g���E�:X9b� �sr2Σ)γ榆��ܟ��ԋ��udB�	��%��6�:�Se���NLh$�O)!�&���3�s�n~Ųҝݓ�XW��W���WS����Cw��שd��a\2�UTv+�!�{.�VK,��r�}�<��6�}L);��~I ��7$��ĕ�ºk8������\|=W�OMm���0AZ�!Oo�ހY��tE��8�CcWJ�ǽ���[իʳ/�Q�u�hP.z\��O���T0uf�b��G��z��RwM�w�>[��!���_�O�_}_}�<�M5��!��M�ܜ�& ��΅VF��G�ȫ�/�Ǘ�Z�i�+�t�q�8��ǣ������0�t!o��P���^�x�"g���b��__J�jTh.#3��׮!���rj��A�g�B8OI�(	�{�e�U7��~�*;�Y�"�!�Q��(_>�Є�i�v��R�Q��z�\�#�[�Zk�g׮���*���s����P�<���V'�q-�p����l�.�	���Ҋg�{�M�h-��1�Aj��+�݁?o]��')�l�s`��Lā�s�;��f�t^������g&I�D�#��A��9t���x��3rz��xޡ��P�_2��#96��P+�CE=E*�J�:�μ�CZb�JӀt���@��:ո�)�xpL�q�;4[1��e���z4����[T���u���˧ꃐ<��цoM8:8m}���uT:`)��9a���Ѡ_ָ�U��J+��J�]J��O9�RH��Ks�ا� w�����"�!'%�Η�5��~m�O��K#m	����F�.o��ŏRq�ԋ�r����-���>+ΤGx� 	y���
9�F�b���ۗ���4m��MN��m+�3��;�2'1 �DvͮY]����� [�s׹m�����<9
�]��lh���������k��vC��t�3']Ԉn\\�<����ά���S�NC4�ه�Yi��h��)���a|&K�3��|Ѹj�' �h����};�t���gLu��� �O���-�,�4�f�Nv�Re��P]�}��}fF.���yw��L��fg�f��o��r��n�_n%�pe5�{��%�����F;�3��y�Һ�5�XU[���T6
L�v�+j���+۔W�XxJ��𥉫�Jd�5Ʀ�c�oz�:�G�����:�:B-�l�C����1_.ʔh@�~L�t)]�������Hͭ�;2�e�f�΢R��8�z3\L!���[i��M�n;��@R:v�f1+��W��w�8��Q�M�����,�Qz~�)SÑ�3c����H���0��)+��c�;�/��X�����*���L$U���oMTI,n�f�0&b�l=
���3��3���`BZ�/��7�j@�_u�]/2.��xWx�3B��=�}�`�a�D�R����C��5l�{���%�ݾgX��_��\f1��t���;��� �&
ER����]7.G�ڌ�Vn�G�:��Fh�a��/�H+#�`�6e���OQ��f.��Ѽ�T�ۮ��f�3��ݪ�P���f���DDG�}��T�Z�Y}�f<M�l�*�Oܨ���A�G|�����A�kꇶ�o�W�O)�~���ؙ���tp�?cK��0�����V��?)U =\N?�U��٧�8c���罛�����'����H;֮C���d��5��3�����n�R�$E�Y`e�В���ʊ�n��Q�2V��Z���j���1�L�0��eX�Y_a֨+x5^o+kw�G�&��ۤaۉ�2P�p��vS����S�L
���>W=������v��}��m!�m%S�۝��Y�{`Rs��F�a_I��j3���dVX���ȧ���~�M���x�������Wº��jp+����7*dIiM��B�>]k�@8�Ր�:uEĹ�w��ռb��N� �a��]H�Q}gSz�w*�β�U ���a1|�3#��t�ܥ_f�����r�MKT��f��]��Oj�� ��
P�3� 5�]���0�H�Ss�-���n~|7���ɹr �� �l:ȩ<�{��f�a���tr���.��>�R?��"����ɶ�,+�HY�O*�/Wf���7���2jLv�OCSN'�P{]��I�9˴�/��)�5ׯ��;�vw\h롢�����빯����:��v�jJ.�L9�7��{��,ʈ����[)��`q�!���k�܍|q�6�Tv�+��.�6cp�8�<�:V�D#�-wdTS�)�|�9 �p.e!�B�!��0�١5��o�܇͙�kmy*H�K��}�{�(k��h���� c#�PǙ���)�1Uk(��˙B���o�����:0\r�i�r4�c��0�u|*O��艓I
\�;��z{)��P�˧ç�TF7\4dKj��oJ�']��7PpЖ~�08�����ۍw{�g^�JF�N1BS�L9�EцwЍF��Wh���3��"bً��� ��{,�.���՛�ʊ��լ�˼�H.H��=G��v���kF��rz!7\Ϡ:`l�ř]:3���Fo�n;�Db3R����A�ɥmͼQC��7�WOk���Q!��۳v!�_*⭬�M�k�9�<��,�=0�M�>b�϶�������I藬S��8.z9N��U+�k����}?9<�e�r�cY�*&�w摷)�5>Ǚ&�)�ދ,�++-��+�vM)�60¸��HpI��-�i�'@�S���\j�]7�5ՒC�php,�m�샃U����:}��/����{y����;�q�6���jq�e:ʁ7۷�;����iB�P�w�񴻘�r�m�Y���>����}߼��y���'-��ϳ+�I�F������O�9�՞uno��2��9����{QM&��v���'�����?��08�7}H �C����Bu��FFa����L��z�\��s��|�+�o��Py��YQ����L��I1|��
�%��d�4���֙�����o�ѦΓ��%�YX�g�=#1���K��Ĳ��S/wj�R��uJ��9�}�6.v���lu�(�� j�`t&t+۪u1q\���N�F�N�[�x^���5�ں�\A�4�7�r�Y�p�ӜtA�(�t!U�L��-��E�z	k��p�{^V�ډ[k�(Z����5p�g�#�I�+�O7t�ݵ��.׼�8�1!�J�u�7�$\�c;��=&�7<
��\l���ިP�bC�\���3ͨ_E P��ZM�+!O�:1>���n��]��΍%|�i.��o,�ŭ�e-�J��s%O �|b
U�߬[�]���[�z3z7G�]����,C������l�N`�Q��i��8���Q�ͭ���oG�,BI5���r�k���d���MI�xZ>EF2��8f�b��^��JT�����A��Y[��<�K�9qw&���WY����F�g&P5�5��/�b����u֤���]vY���}U_Q���菽����V�AEjD�E��	��z�GF�@R����Ɗ���P�J��[�I)�UE�)�!����/`ʙ�#C
��U��5�[�^Jǰ����+Q�M��/D��<�ܿ�K��goI�w&k��Ļ�� �41��ӝ*�N
����x��'A��z��<o�v_(I���
i6v�뙌VD��0p�H����B�h%�i�����\�;��ە��z�p��ӹ�S{p��+���Qwa��N�U��ե�0��v�#9:ܮh���|����
ȫ*%�)���?ד܍�s�]�b�2$O��3=��Q��/(��������a;���k���||Bڞ�����}���u6Cǉ����f��f�zrn�诹&��o�vm¾����ނ�8_z��X�!��%N)���w�W��j�*���[����D:�����dRZ�
�whS jĥ�gb�U��廆�]k��O|��)�V�^+i��)y2h/Π ����������syVȚ1>�/�om*�:r�a�˾=g�4� o��W]dY��6�|��0ҳxz����k���yT�k2��^�~��#��u#v��n����R����%*Wż�p�\c���z%�\�@�vk�0��_�]����x�Q���oMD�s��c���_v��^_\J�w4e�:�,)콡C�#�]%����)��O�����s�=�b�T�B�׍G*��;�91YQ���_wdA`P�w�1���Ϋ^�',R��L��jWޥ�`�h\���9��R�>��B��hvb����.]*.�q�qj���ysK��p���R�O܆��u���(:�^:��5�9M��7��[Z���8O��sL;�7��$=��X�e�^�`��T�,��.^��mr��Yѩ�mL�B�
j!7�a�{�F��7*�FSjz�^�I�Q�Gb�%>{��O.kW�ظ>h�u/,Z�}�m�Mw�r{��1����E��������}�U^�v�f�H|��P�ٔ+5�̨ �85[���*N�l��zGDG�M�/-�z�r��+�eq�Zۇ�'dF1Ҭ�;�&�$[�򃵻��\OZ8�6����@����E�R(���T\�H�z�7&��ˇ�e<�i޶����������X�k��hf
�Y�aU�`��D�n�t�Z�o��{�nGRBmj��w�m4���� ��fp r�ő���fF�'u�U�����7Mh��%�r��e ��2��)8`Z�-ʉ��N#m�$����=m%��Kl�n�
}`�գ5�hK@�X&��|�\�ŕo@�N��z�E�����V��b��o���V�>44�wuv�qۺ�e��j��v��tF�
S���$�M��i�܋R�A�r�ӭ�d���& o5�����e��1>�7v��K\���7�}M6���:ĮT�v�E�tl]���=6�� ���9����ř/��='%��Ll�V/5W)F�;w�.l���Hd2��!ºE7�7A�ʺ�f�o!I��x�R�h�3w��^�Z����S�*��U�⮖�n#��v��}�rJ�[���C�)쓍^Z�{�����,V�K�X-l�.=�Q�����Ү��aƕɪR30i���JH�Z� s��Ɩ"x�����+7"��%Dܕ|��"N�\������s��6�ukWrm.9x�y�-crtoZ���J�S�sm𗘕Ʈ���U�c
��@ӧg�Q�'�e1�rv�<xG
���i���>k���ƅ[Y����ܫF��Ȯ���AM*I���9��i���R�m�݋�5f��-�V��
�v���)ԦCX'o��t�;�ݫK+i��T��mt�4���WZaR���)�t��s��=��#h讑�qM�P:��Y��v�Q�Yl�ayh��m�Z�
����J��e�!:��.�V�2�Iٳ�e�v��Z�pd�F�;�efs+�xƁW������n>�ݽ��@FoXO-9t���.^�kv�ڜ������
�/�t�U/U�E�˻L
>�s9����òEнݺ��ģ�3�m�EQ�mwXU���a;�9��[2���X=+A����*tjG���M1��S3���nqn���^�ԩLnF��ݼm��l�W+m�j�Wn;�K�t�v�M6ښS�)Kj��r�+�f�n�����-��́T�I�+	�i0;Q[t�J�MB�nr =�U�y�]��
�T��72��%��֩��n�Dk�y{"]��I[t_0��bۭw(�e�yW��ŻV�wg�O�"�:�˖\/�z+.^PP�A3��o��K���䨰��;碲�f
��&\jKq��!�l�jm^�w���/.mY�EQzE(�}�i��;"W/�E��w	ȍ�^��2;f:8ܙ���YX�n.�6�k�z�˶�JDno3-Ź�s�B�Qe���M��a��}��We�pY6>���U��a��_rBW�j��ϫ��"|�'I����B��r�嘉s"J�ruݥL� �fF��ȩSK��br�5N���&FWU�B�Y�T\���5"+"�˼w#��V��'���"�XYY!jT[����l���EhD�mR�g�t��HQ���fZa�B�"�%R�*3���Y�eff�Nxr�2L�ܗ������$j�hQ	��e!���,�B��F�]R��3��)P�J9H�J��L��'Z�H� �QN��r6X�R�T,2��=�=�V�$a]E��9�(�&����R���x��%�[J�R��)Y�PhaX��*��]3��C�Dt������$���Q{��Ae����t��V���TA�)B�exxw3
�*�bBT�6"����Q��s֊'3T� �TQ"�j��U�L�QQ�^�յ�PH��T����*" �IwA,�N��Ď�n�((���R:g�=4uDZ�̠�9°���;�T���C)���u�j���`7Q����j��R�V�Q���
�Ok$�.Vn[�w��8�oL־o{��3�Tv��tF���_��k5�ܬ�vn�ʂ���Tf�9<�S�2ӑ��R\�u�v�{����)�q�ksy��?[���`UF�@���s^<�)�H�������WR�=	^��L�*M����Wf�͘���Fwr���7��֙[��ì7��{]SS����_�[�{���|���
��0�U�Sw�����<��� �ڗ*�����F���5�b�ҩ�(���QH;��+�Z�v}�y��\rB���I�TKtxW���acb��\��.N��7S���s�=Ճ�;��E�j4��n�2L�	���BF,���.��{Q�-�_�������+�_wd&�j� ��5Yӱ�ԝiJn�<8�0=���ni\3z���ȇ,���I+��(�*���(�cA�������_b�4������ ^��0^f�v�`FmR��f� �0F�LH�W[�j�GC��|���{g]cϞ�ڻ>���Z�)�j��t�yi	&m��ٖcY�2��/(�����ֻ3���ꛣ����0�֛�#s�w���u�0��}K{��m��Jj�ke��ﾯ����u�<�I�`���.�k���z5'Z�Ĺ�Bo��v���(M�w�-�Y�P��d�1��)�뛕�9<�z#R��5=nԓ��*�����Z�e�4&�q�T�F�"y����_mv��.sUy�%�v����Y����q	���?W�������]~�=).:�����Eu�:�I4l��s|6��n�+������O�mh5<AߗZK�G���B
�����)_[�����Iz39�e���2�O�js2��p�p.�����׎Ӿ��O����VV�IL+�.'��R�
bڹ�@A*9[�ᵜ*���r��6ol䠯 ��w�iԝP��c6{�Zu�D�L‶�K�v덾}p�n���@l�� ��.N��*b�f��nlӍ�]����/��j�o��}َ�=_Rd��'�zU�Y7	IR��w��Q��~���(��x���~��O��Un��K��mo��Ԃ}a�NؠBͼ�/a9�?^��l2�c��n;�iR�62j,��ԗiKk�<�-L�ե��7q�r�}L���e��_kᣔ��˷i�Jr�Q?���舋T�t�z����}[cj%*5��pլp��M=��5P(t����:/�Q3���Fm[�n��PԻQ-颓ˎx�d>��\��wMha��כu����k�}G��w���ܗ�oV'ƾ-�\o�>OtK��mӫjt�IqYS7S�V��>��T<Q��Q�s�z����f&`�H�q�6Q�ܼk����i��<��H�΄�CE�s�-܀���	��n��ך��)��M&�;��j�O!��=�6*��<�r��Ԃ��΍s��v��������]7�5���Pۍv�5���<��k2��菓t�׈�_i���y���w^tj�I9�n:_ɳ��3����C˰h���r��߭.ё#SzzdGs�ɷ��_\-p��� �+~c��5sɞ~�-�r��	�t.�������kg�fy���E�a����WcQ�6�l")]{��i�de���Rh�	V'QD�g�61CQn�������ݕ3M�_)�q��>��|R��tƽ2|]�v���QkX��S��*ā8q�[|/l�Zr�^��v�8{�U���U4Nr��w{SV]>67=��D}J�y�u-��*��h�~��H�}�����*3u�����
1E�].�`+��ڭc�q�xަ���5}~�j�~��H^�A�֖�5n��צ;杧[�K�sν���U�1M&��Ko�Wf���d-�޿Ml���&�HZ^X�z&�.OK�Е�t�b��X�z�s�5��x��26Dc���N{f�_8T����N�WXU��J�y��q�˖n����#�~}h�!��ÏL�^�����).�A�􄝿��ZL�{9W�]�֥�m�!_Y}׏LZw��GKU�O���(���)+�U�r���ɳI�kEm��,��zo^�q�Pعr��q����KE�M`2g����'�EESٜۧ�i'ڶඕ�w�`y��0��#��F��EP�
]Z�bUu�s����}���.j��w�
���J1?r�pDjqw֣F�s�9�y��Y����Wʅ%pR��V9�u�zt���5;c|p�E��u��,��녚��U/��S�J�w5�`��=\
�>C2�YV��6�=�v;�+TH-'s��c�v�t��&�7c�_P-;9x�p��}�UW���L3��k�� u��-��Ӊm\jN��龩�i�p�v��/��R.8+�N��ZP�c�P:��߶���n��O]��ic�ì%4|�9��L���v���G\�~�,�S�6�~^kWz�/�w�����H�N��7��\=��󹟵Y��A�]C1T�������2��|��k���v'|���s��_>�z����֖�;�g������I�h,V�qô��x�e���źŭ�f�➆��i��T�z����l{���<�u�|�+nOCW���4���6.[{q+�o囕������;o�����(ˤ�=s ��s'T.Q�Ҽ-���ܦ�-V9����S;�BS�6��U 6~<�UR�\WHT��������8���g�d� ��n��y��O��[��rB��>[)>�T��*vFX>n����F�g7F{k!�����kq�*�(l����Wp�W)Š�� oa���(�qf%�qh�1uI��v��ٹ�x}�`��_٤��']cH����	��n��a�2���b�]�i#Էj�$�m0H=�.��
UF�К�����o���ꝴ�,�x���c�SN2��̯W=�)��BҡC����P`w3EN�uVj��h�2�t�X�����#z��%�5�ˎx�d}�3i�s���L/��T�,@ᢦ2�a��T���Y�oV'�e���Y���ld�eTl��b��o�jr�pZ���n��Q���#��q�I��6)�	�Qܻ��T���t�~��Ǿ��8��ʠh5+}=)d�����	s�7Xp��&6�c)Aե�Z2�E��+�Q<����TV���\�n5-��+�����/.�fWc��Y�Jn1�B����y�N��Y���#Y�~��x�N̛�]<M�����U��']k\9�{%�x�|�������~Y�S��۳��7mm󝪖g\����u���{�_5�k��s?G;7�p�} ��s�q���Jm1�v�R�YH��{3χy�w�[����<b�^�32���G+QǓ�oc�B�Z����ձ���uw�2�`tS�g$�z�l�왌��F��P����oR:�)L9�쨙���O[�ﺔf���f��:p�]�e	��t��uD�۫�K3b�v��o_N���o�d��x���}�WR2c�g��I��v���x�_Nߦ�w��¸��o�f�Rl1�cwܮ���	�'w���/�ej�}��-s�k�SQ:�����[��v0i��]kO����_����z�v���9_RG;�uVԹ15y�)���%N^b�oz�n�O8�)���5��}p�>�5��z�)�D��ά���T�V�đ�[�T�vJTj57����1����/�y�J�c����m�8Tp\�M}��q��-�ߊO/�5��f�>4cغ����u����K�P��7��
�ѣ��|������o��D�OV���Jqk���й�F~�:T%!����J��.7B�1z Y5}�M����:���s5���9�K>�)��u%�������Qp���勷L��9Is���;aڸ0�<��·\3q�QOs8�����y�E��Ms�w�5�*.��o+8���W��O(�v�ͼQU�k8��1�0�;����Y�ڻ�>w�hD�;E����!���c03D����`r�Ֆ��m��`�ë��a�97'Y8�j��@'N���}UU^r�I[�ύT����q�n�_7�<��ۍw�1����76]T�t�� ����К@˘�ot�yKu�}��ZN��c�)���.jb�9E2��	�չm"���_�U�U��қ��H�����j��r�ֵÞK���"]윸����r��}zVQq�f��c$_:���;��+Fg&�r��"쨣󋅸���{=��g#�'���-��~�v��-�x����u�O�&��қ4�w�s��\�|^wE�sk7��u�vl�n�W1�PU�Xp8Jp'VԿ���y�������J�-��aD���vm���9T���TЗa�͛2�U��\	֪zj'z��.���}nˈm��\����]U	;��hͥwI$J:�+�c�{;<]�]aTJT�7}ᬼp��Ib��+-^����&�)o�3Y���LG :`��(�I/�Pe�;�I��=�@��狱��#�V�iK����.P#!hu�{�2_
��z���M�Q�u�cG��M!���N���ݚy��)In������������W�P�R���݌�R�u�!틶`T~|��=c���ύ�1,.ˏU>|9 �gh�NN�0�Ʈ�+�UW�{��y{���ِ��M��P(t��>��I�	)��r{�j�T�'�O���K��k�qW��Oe�o5dw<�Z/`��ً�9�5h���?V�V�ڭ�9Y���C/�÷�v�M+�,04+�?q��)a�C��⯍����q�sA��5�z�j1��\��w����(�ef���T*���0:�S���78���N�֋�o�j9��n1��4.R�oN�s��V�����_��ڧ����=�O]�6�u�^�T�p8=�S�+k�J=JM�?y��̫<��я<�{��T�bz�� �7�H(k������-�z�ָs�h���f5Y��Z��f*�3o(CXw��%���9���nRv�[����O�oi��}ih�[R�MSn>�%���U�)���r{�g(�|ڔݟj��bN�x|BB�|�4�퓢�-e�������.Y��ɴ���V-Y�9=u����Һ�ױ4��:+)̮�سŪ�G-������}��Y��g ӹ�ʯC�4qI&(�G|�#��
V�(�{CWaY\����@�g��9���&zLø����}*VQ�|������uei���b��mRl\KonWfᣋ6[Q5!���X�)aJ{�(���.��`UN���P��t�6:-��M���맷���OO:C;Փ���w���U�ϱ�.�=C������ެ�!y�{po�$ذ�rs�'�����>�����m^��@h_>[��s��S��zc7hI�ز�޻�r�G$�\5�-������Q#������B�����ܧOQSY�����]�-񯠷�sƻ#\f�+��C�/�ɺ�����B����բ����Y݉��Ŵ��չ�7�+��d��qd%���@b�}}���."�yB9��O-����X��D$Ұ����\]L�#�NT���R�[p���a���$�s�u%�z���h�]�ف0���+OS�It�L��h;��c��pT�+xb�{�lQvb��ؽT��;p��0��'����,��,#�1�T!4upoNWʱZ6�ƹ�&�C���b�n��ū�C+[����8�䏌��b|�{t
H���w��� ��}Z�<��o=s�����/�4_ʆ0�$E��`���X��ˇGO�X�H���[���s
�V�J��u1H��[͠vj=2Ô���wv��'0�EuL�v�ކՀ�p�"���+��vu��Uϙ�}�0�)�*��Z�+�G�y��^�+n$zT�8�,��Q�@�ھ���t��\��#MP�=y&K�����D�oIqT��ݶ��Q7M:�k��u���h��b�4I�eZ�Y{h�.>�yQ�[��:O1u��E�/��$LF�^v��|�N8U��gh��ݕj�j�qa�����4��)���0;XM��F��:�cP��żn�XC�#�o��B9H�w����P���`�a��lQ�p&�Ǚ��['0�o,ops��FNT(a�����\;{m��`����b��\\��(e�#o�u��8o9�3{SvmwY�ϻ���]ϣ��E
�`ֹ��1q�k[μ�{��{�Nwȃn�f�[��$��(^�I�X��0m�|E�>N�b*ќ���i����۰N�.�n��8
�T��M���ہV��G����4I]�"�C�'ҩ6���[�E9k0av�I��2h�)}Z�vÍf���\��H"�XkV��S�f�Y��� �6�r���9��sIe&��u8`a����KB�2.l�Q�y�� u�Q�c.�p�Dfվ�6�n�l��͐�5p�{�Ե8BA��/o��6�/y�*��T6"7�j�r��������ӟ9�n����W�o�x+�u+��37��������1To5N ���wԕ>�!���G�%]s�^��aHWm5����m*�p�X6����
�Z�y��w��1	���-s̹����[@U�)�]:�i�rPM�e�k˴/��`�H[*72��S�tou�����G{���b�D�2���ϳ�(�w;��Sһ��	WOz�
��̝g���+ա��1�`橐xl%��Bw	ɗ�7�l��)7����TR�+1���$L�t�!u
�)oWqk&s�ͫ�����j!���SʧPԼ�#�\c��j�B�)������t^������ќ�$Z�O�����#���֫�N�]t�8��C[�˖=�p�ˬi�A�7(,C��gIY����̈́�w)G�gP��eN�Ec�]'��Bz6�rJcw��E��zU9�7�\�� ��B^��]2�w�v��Z�v0ʖ��J���tϏR�u:���1��Wz]�آF]v���ќi�]����D��:AlT�f�w�l���8woW_N%��CY��]r�k�fȚ��*V���b)�
r��l�̃^HGp{��7�6sV�=؞���(�[��a�;�}x��#<w�ޯ���r������S���T��en�/6J&[X�z�(hU�
�������k.EE�B(tV{�EU���E�*8�ÒP�-"�QR����S�k���K'J�uh���'\��g�����8��wq!�U����9Ez"�§D�tJ9W�����%���rvN�8c�G+aD��B�Ҫ����Xbs�Js�Ȩ��G�r�t/]\t\�s�J�#e�gB7q�]iQ�\���(�gK�)�*�/!)<�)�2\�ehj�%G(�D�Y�+3��3�GJ!�T�x�z-wqP�V�������U`RaD�y]n+1S����Os��u*�Gn��I)�nK"n����dREEĄ�]ېW�)̔�q=lĩ<�Ԃ3"�L*
wprH�,Ι�֩������N�matOtJ*rK�QS��E�[�p��/��q�Rwv�eFe�UGW"����L	5��R�E-(�^�IDDY:��|��qoq���:�R�]p��q0D^Q�[ް3ש_���{QB=��O�p\��e�a�T(Ƌ���F=��W�}qK�bof��ٻ��5SK9��MƵS��C�Z��;G���-+������>4{\esS��Ub�I�-p�S�:��[�w·:X��*�8��i���y<�F��a���5��ܩ�m���-�ά(�|󱩴S�3FeANcᘨͽ�+Fg(��i��e�8�5�_���\���u�y{��Cޅ��J�qʿN٫Y�޾(z��w�O6�G�����J�ǻ�^7~Z��Ot��yE�����@���u5��c�Ө�^�=zEk��Ht[��I7���]�n�~�!o��n��*��@a¯��U��x\muf�K��X�-��p�\6�[���k�DλVp�mH����}�N[z}+�T1��T�W�WXu��F�7���k/-���-a��Eo���L�䂴6�eA�܍F��)��5��_��h���٪%�o��6Q���~]�Ƭ�&]���Su��ֻC�K�^۰�"�5-ܴ�ݟb����b�֠�L�.�׫��Cý�a�Ԡ�(�4 l�*�+r��jz��:�"a�!���u�u����wpT˔��v�[��EZTeb[�{�.u%�fI���Mo��!^t�xRuc���>��I_%����f@[Չ�-�ti��	i�*�������\bwn��L\�G��P�1E-;���d�[͍L%p��u&�q�E8�Ԯ�o��5���9�K>T���Ww^#���c���o�E��8�>7�˜�o����p�)D�G!�9�����0�՘�6����No���etj[���C}S\�Pۍv��荕�-�+K3F�D����� X��Uq��w'S��y�o�$�j8SQ	���c��Ν]3�N��Y#)�=Z�_�;��j�)��FoOERy�Z�~�/�Z�W�rD�c�hj}�"�>�.h/�;K�g�g��.ч���;F��WB�����|VE��*�f�U]4���9�|��5G+������c2�����Tf�/�/�	ռ��o�:��:l-��0�$���)�n�m�k��6��c2��i;�J�!�ה�����%s&����_����1*m[V�VTǘ�|�NM8���K��z��˝��d��|x����]��G�wa�篞n�F�*A3�h�0���:��6=�5��Z�������X
tΞਭU%l�BB K+U��ߣ�W	������^���rz�/�0�M�����vm�����9��3�G�7I�Ah�pz�=�ڕ5:�+�.��lU�k.o��>����/���V�ܩ�MIM��� 6JR#����
�*W[��e-�R]4�t�˶Z{�'��q�kz��@t����m$��n{�]�Z:��X��G�0�7�,�y�*�:��L~	1_iI5_�z��-'���G��#�ޝq��N/y�sQ�������XAV�a)Nռ�I�ԍއy��z�wm�SJjH<�PдQ�#��ٝ��9���C�X҅�o���]5Թ�B-����r�7��@v���pŃmeTm�E�5iSQ�a�`�]@۲�ɴ��jN�Z.�o�j#�a���6���i^���x���U�Nh���X�^�s�i����=}���'gbo1���v�U�D{�~��q���!���������e^�]G�M�$�)���I�כ�V�&`����12�+})�N$��l��N�Ѵ�e��uN���Ƚ4q7=`mDE�h¹�M��0��}B�Y�Z�ѻ2oTo��͋�R�v����C���?;��^}=s*�=�ћO|�Ξh��+{�H��v�+v�{6�ɺ�Z��[�:��j�u�������錙�؊afm��|l��1��u���)��!{'�S���VT�i��0u�zl����F̥�Z����񛬸��ˌ��Ӹ��z�W�s�bO�^.�1�<����s�t��2��3(��rά�!CV+晵I�q-��U
ذ����R���UϘxݯGf��̤QW0���SS����W��c#�J�/L�N`�>N�7�g����j�!mV���=�'<����䝥)�i�#�$��*�ܑYO�/���Yo[�)�މ�Ҡ�+f�`m�v�{;[U�˟ѽC�[��<��n8X�{�Ҩ:{�����wH�ƙ��P�Wٜxgs�k��o�|[��vF�ͨl[+�L�Գ��9ו�B�[�J�re��UC~�J��'�����
ѩ֝5��f�kY�R�L�#�JG{�9��Mݮw�%V���#w����2���*<�ϝ�v��3�gl�lV�����L��-
����6�����g�H^Y2��ub��~�$�t��|��/���0X0R�Zy��z���n>-�3z��]��ȼ�A��tKcsC��98���9��x��X��$�ꮵ�J��1hJ{�2� �9�L*G�pT�sҖODjL�nB"u�8#�Ĺ�u�f�:�{�қ�ᨴ�W�(��6`���9�㜨�椺����{S~~X,��b�K��SK9���q���u:쉎C��kc��iN�<�s��,ͧ\���)�yګ��k�=od�;��f�R�a�!�����������7��h�̸�|6�Sܛ{�__�_5��n�pP�4[�͙��Ƚ�Nҿr�K�a��˥:���x�ٞ|jB�u����{�7Ĝo������2�Ѧz��ƽ��U[#y�Z�i-uN�S��P��WК�:p�v��5�\�{�C�D���y_AW0�Dm:�"�y[��*S���+��-㰦��M����t��Z���޷�f3L��3��K^�>��wG�y-�i�ǡ���,��y�V��h���r��YK�Q� cj�C��_w�Z|��V�������y�oWnQm�C*]���]�W;�4��ng,���|v�>k�����n�N/M�PѮ���Q˼�⇼�*��n��T���pU�Ҹ�ثp�\Cm�î�#^TdM����g��2�k`J:z,�?��=.z�Q)Q�M�Ƹk1���4�;�ڍwkNf�v�X������;���JJ�Puސ����q�}`��yY�6����X�i�1��$u����%�G5}oTb|LEF��5v���g��k���_W%}ק��b�I��(H�X����ĭ�+Պ�P��5ݥ'�q6���[�s5�0��9�K���:J��n���nuf0����#�9�M�v��FB�L��k�)���X�l��G/:]7N.[Ss�m\j[Q���L�sLMCn5�B����랋}@���Sݽ�ym�	�]̫1��U,�ڬ}祿=���=�����r����n�:�]���|zN+������=A��Nn#t�`�it�f>!��(T�s^S}F0^W�e�شWJl�c��o�1
ϘG=�dgS��4�����f7��2�7�e�ˊ����ܮ�:g+����� //h���$�u����H�ԎeR�Z���~���3�L���y�5���T��%�chE$��+N���y�y�tz>�f�Ɂ|� f*3o�Jѝ�KR��;�%�oS�Z
w����s��9^��#Y�fW=��`�XQ�md7�f֥Ӈi����8G�bۈmw_ݛ1��G1����U��E������YP�Vܞ�������[}*��]�'k{U�	]���e���F_�H'G�A�[R�uBW�����e�m��d�sh�h�S�je����X��1�g��@l�NA�Q;<\��)R�-�7ƣ�@�Է�Gf��{M��kz��@t�>Q[I+�'Vٰ����.��z�M��ez��y@�JT(w|�>*c�����슫�kec�|�g.qսr�-�\3o�!8�lV9Fc���u/��i���6b�w�3jE�����*b=+�G��9����;r�U����,6Rc�q��7 ����e-�M�=If߽��D���������}B�_]�7���.��ˬ�{�<+�HF�xb�ֶ��sr������k�r�ڀ�&��d��UvRR�(J�2�����`[Ջ�n
iXw�W���E�.5�)	���n&�vx�8KbVW������s܄[��9k���;Af����<�h�RUr��S���LLZ(�ȹZ��Y]������ʛX˼�a�}cҦ7�^�kmQ�3�W]�:ڱ�oĎm:{<�O�xyR���W��Ʃ]ی��p��ic�4���;�S���2�:[=�y"#�Oծ�n�iN����9�|���rmo/W\B~�d>d?h4�����������R���2�ڮU�2�q+�m�Q�I�)��>Ny��Cj2�a'��/h�ثԐ\'����7YI�2�9F[O�R���9�����V)YB�9�u�V�w���|�#�+n"J����晵I�赾zL9�C�Wa#9��VWyk͸���9�S�
����Q��juBZ�`��0w�=��[�klWQ�u+��{X�F�uհ�Xݻ+�u�f�feˍV���:�1V]��kD�1�L�{Jc&C�;��'2�z������ƕ��uК-��1r�=ã���ퟻ�cN/�A>5�h���͢%��W2�[���w�4:&���~jO5^>�?g���^UFB�޻x'���糨%�B���p�m��c�^8k��yk5�B�O 4(}��Y}p�΋�+���V�3}�#k__��2ܜ�I�놶��p���-�4�@���eٽ�n� �0��.P���/��n#Kj�k���4[��mj�\f�b��{�+�0�u��7]�Y. PS�'?A@�KEF�k3෪1>��J�[{L�Ed��u��J�����d�l�1�r��we[�'�<��֧.���M��т�4δ�_M?�4�ͱP�D�G�y �:|�g���R���ju:�]���L��Ӊs�M�v�v�
�L�!�c�Svz��:{�� ۉ��zܙ�{:�bx�6�VsЛ�w+��5��s\@�3 ���w�F��hM8yҷ2V�_F�ڍU��u���z�엵�]�>������o+�Ms�;��t��O�r��|�i�ë��7�&z�"�VYm��"�8Ѝ�=���@Zh�j� 郧,�z:>׏oC�x'�p�}W:���{L����W:�u�[b�Z�o�)W�bY.�Xz �d�Ꚋ�E���ml�j6��gp|8�������:[5M�����\���|�Ĳ~QW`d)�)�Uv��o$ѧ��KD�}iv�0���dή�w�[&<��V�^�(�����N���yT|Aڝih���U5k8;��o�l�ft��y�/��{�¤ظu�m��q׊�Ck���z sj{=��8)����x������q�B�-��܇m��Yw���/k�{J�@F����Нe�i)=9�'+�Kb��Yp�}p�>��4�Zm=�}o��4��G\W ��s�=/k�*�J�joo\5����K^ޯC~w��XJ�����z(t����f�JJ�_Kzk�ǦњM��Bo�=ט���N#xf��r�u
0�}%A����O5��8T�V�*j�縳���۟'�+����qZF�wX�4{�{�6I���2E�f�wS�1]u���vX};�/h�uVs<a�2e�2-Y�q�I��+@���]}��Xq��8h������s���q`���y�wa����^�(Z8<�Z����M7v����h��NJ�m��hPӣT�Y�bg�����nP �[G���76j�;^�j�����sj��Z�*"�11iw^�)���^푧D`�`���
(�5�sR��Y��̴�[�7+^�;Z�n���Cm��ꛅ����ڐ�t��ٻ��y%�3c�}�𡏝I�
����@R���*��Y���w[��0��r�l[ǀ�`:�Ķ��	Ya�wpÚh�J�����v�IRި��%�xMk�	ف�Gy�w�N��I�g��x��LY��wb5}.�S����]/�\+RÖ!�}\�
�ռ(��jS��&/��:^�4;y}2��j���7�J(m�Һ����U%wZ�[� �w�$Q���#�GY�K��\�D�u.� �Ϯ�t��`�4Zk�QB�%��mۼ�Ю/� ���-ʝ� ��)�g,\h�7�:m����DVf�&*x�o��i�n��y�]��O��+��&�ͫ��d�AʺgT[�6'�F�������";�Ţ�����\�a��\M�����}�vF8WwQ�x�Z�fR���5�;��;��L6)a��I���Z[]j�\�ج'�n�DD��4�{�*��G�;�ۼ�e�l35V��ټr��EL�jq�{���kM��|3��Vp�}o3��lu����v&����&V
k��Z�	75�]�h�L}X-�CH��B9�N�������I��#��up���,L�����ДC�sF<z9��
45:�Vwj]���˲n�4��u��X/��K�V�48�C��f���T�W�>�7׼�L��j�F�Q��C�{Uf&0cVέV�F%���CE�@�H� N��4ݚwŖ��3��qPƝ'�v��R�*|�f�%K�T-Ґtzi��u��/�t�����Oz���O�$�*u�ǀ���E�����֧�-Tu���U�F��9ݓ�'��v�ŝ|M	2��Q�m�:�՜�yCK%��b+��\P�\�Poj�r����*0(�+\���wKLk��;�!C-dB�컎-B�{�֦��!�:��u+h.\�H���ƕ�gL�tEt�����zL�O3�^�k3]��
�Z�wٸ[�ĺכ��!�Zu(2�jߟ�����/T�RN#,q�����_`��z�4h6���:kt	��{r�gqv3��B9�vgm�qs�}\D�膛�*����**Ň�C�[e)��>�]�z����V<G0��Di�[�����k!t��JxD���@v����U��%�6�����e.rVH��]�<����\�(ڥ���:^cT��c,F݌��Vnm�߶��]42'SZ�]Qb�yz%s�"���U\�&��$[���By�(�[������t�GnS�b�*�I�'#ٖ�"��<�U�{����+�=�q"��Ny�f�4�DvY�̓ւe.����xI:ӸBBI��]�y�[�ig(�'u',u ����N���Q
iN���᥎���;r�3s"(󬢽H��B��������HJ���.�雨Nf��8z�T��i�:N�x��D�Ⱥ����<��-n��p�*�=�%�����ҽY.뻓�N�S������[�E,�JK��]g-ws�^b��wq�R���<哞+�z绘�/wWG$T�N{��z�"T��.�C�E;���w��2�Z��s��nn�{��y��� ��տ�z8"�[��/��OP�g�<қx9}�����}����U6�ެ3��ɣ����Ժ���]r�͝��n�w%ӧm�����m.�+�Jٽm����D�Fc��BRV��-ȭ��u�8�9��f�ͺkvj#��z|�l;W!J&�z�.-β\U&Ҥ�]|�[�m,��j[Z�t�T�G4��n5�#5ɚ̩�r��=�v�1h9�[ڀ�
�͝Oj���S�\{��p7�kf����{Ͱj
�Ht�j��&.^�;Q�3��Z܁�h�%3��}Ry��T���n�wW�x���m���r�u�;��]���2~Άb�3o���)waP�Qū����o�-����7�ܞ|�^���V���y1���]�?�NK�%fu���z�x�{"Op��
���i���6.b���}ٳn�V�[[��D�)�/W$
��[=9�\5x_V�CI�q��Uٲ��@�i���؃w�Ov�������૾UFԹ��T%����ثp�bh@W�y��;�K!����k��n�KLm�C�Wٻ[��/gq"��W�Uǡt��E����.�~M��6<έ��=�e{�.ʂ��Hg&�ƛ_�9�եӛs��2�,���h^�>tu�Ic4Ćv�������cgs�SN������5�9�+���n��nC��;�7�b����9����wn���ċ���D��=Q4�ۏ�oT
?G :J�򍔑���͢s7��=�#o����=^�Խ\��ù�����|:�_)ʄ6sJ�.�r��C�8��o\�Ƌ}�;�N3��9F~�9����`���]�o8_RpP�h��Q��o�W�w�d�*L�wa<l|n�C/o��OItC�<�h�n:�=�E���\��=�~�z��e�
{57�r�ݱZ�4#e��7�Cnb�k��Kj�'Q��~���+U����N�6�_��a��p��tD�m�w7+wsk�ξȫxw���C:�gv%�g�n�ML��)�M�z}]�B�᪄�P��e@��������l�Fq�m�G��l<�^�낯�)z�I�~i���\��^�d��"��?w0��aL+�;�ґ�`9幹j�6�k$�Wz�vf�ޮ��FpBS�6-�h�4M>��Vʶ��\�,X7iR�G-��M� (�3WZ���0���W;�՜H�X͈+<�K�5�]zNH�oU�'S��P�x.�ڊZ:�մf�.y���N�ܤ�/'<�F�Yyj��M��Oz��bS���h̢���Fn��O1���~�i�)M�u�b��̨�٨l�j���V�p��0�:�_9W��5k5���P�e�26�e�f�8��\+�8��{r�6���d6����s�s�?4s���1�Va�4��U��sEm8¸U����zyO�yQ�����K�3y�{��8k7[�ݞ�q[#k�z[ˌp�\=o�����]5}[�f�N��v�VC<�p�T1��V��C�n���5�[c��o�٤���Ge=�g(���h��>�.�F���k-��-�s��k��i��]��U��o��UC�d���/��,)h�<�`[��m��n~�PO�r���*��j9V,���Lc,��\ﻩ��6���\IV�l�yY�U9[�H�ٔ�޲']E�i��\tJ����|����hӂ�<��6J������y4�|�)(M��Yт��:�c��D���Y=���u�;��[��۬�`}��S-k��eZ{�3���o�ms�\Ԥ�@o����+��r~*�+\�5�UToP-N���Ң�v^�U��r�.s_&�;�;W�f9�S����2FS�F�9�9U��.'ڽKkS�6�jsI��p��5�Y���C �I���n��72,��ݽޞ�ߞ��ǻ���^�~���V�<��_j���&���
wά�����$k"᷺�nV;����8�g�o
���Y��6���{�m�G3��]i\�Ά[���PQcK�(��7�(��Y��VͿ���8�5p�n�n�[�u�fQW���u���E��Ms7a^s�an���f�Rl[�Z���ͽ��H<}�Ћc�mh�X�i{}ٺ��f�D����.alW4޺oS�ݸw���b ��2�,M
�Μ*�4��%�ސ^�mJ���aTbt��-���5����|�Wmve�2p�D��Rγ�g-,=u1+�ˌK�k��ȧ�`4f}�s7�F/�W�7PX9d��R�g h/l�
����;R{7&v�dT&��[D��K{m�5IC���մ�9hL���Zu.ھ��ŕyH԰b噌��i��t����,�[�zu���;��>߻zV5����s/;�o�p�C9t'�<pV�kc��]���q��*ù��Ғ��Pu�ȋ�<uz�"�Z��߽����c��VD)]P(r��D�Z4sV���8��[���'ڍ��;}�����9Fc��P��:ц��T�l�������E�]p�o���ҿ������D���9�:�4쀩�*�S��o�(�ӝIn�I��{˜�&�8tǹթf*D��C?U�s���Z����y���Z��q-��Ku2�ٗ����g^ɝw�g-��U�h��u��<����?���������K��u���.:��N�S./���lu��D���'cz������VB�3���d6�����uf�r���Þ��uѿ��:��Y������keܞ֯[��unb�F��鎯�gz�E(/c�<���Gs��5v�f�;�!3
�O�����u�	u.k�X�,m���2�i�����z��:�{îJs!�l=O��v_>;��)]V'a��Y�yغ'��;�|��gc���*��\l�A�-�n�+���^���W�:_z�c���s�0�HUF������1�*�qWQ����-�./�qХ6�͆�u�f�'��/.�9��en>�O.�|S�'�9��<��{��_W�[�I�Ko�x���sA�)�S4��]����1{g%��U���ڗ5:�-WalTe��]�X��*���S��m�����~�"mo]��U�x�u��'��	M�dur�}+)���\c�����M=���Lr�
�(��ugKg��+H����Z�?S�s~���E'���p��q�R�C���f��ݪ�,�;ΰ�J���ԱNwJ|j}�����9�L����Q�1M���Њ���'�=b�w;�;ܗ��j�����K���&�M>�*Tj��g�#�	J�����_u.{��u�z:{���#�P��輝2:��9z-_!��KD&��׃|�-�Wtfz���-&L����E%j|������!��6�َ�D2qB�w�b�B\b�9�<�������W��z��t��y���y(2�ҟ^��-%{��/r�oX�]��2Sn�.��.e�|�b\2�1�¸�p�1Q�l�ξs��~�U���}�7s��%o2i���ə��N#o�ݩ��v�w
�����<��H�խJ�=~���5�&I��H��Û9��It��b�4��v��5��J<�r8�u+ii������|�ӏ��{Ӣ�O=kW���~�d�П�9�> ��G�˘����ʿo��4*�*M帞|6�S�ܤ�������ks�&O+/���}����'��;I�[Cݕiu��#���9D��Jl/�T��rNg�ܻ����s�j�'<K~K^_ZZ!���SV���o�u/,\W����jyi�_ʻ�-��]�,ٽ���૾Um:�\����(�Ol<�ܑ��tϪ�z�0�*�or��/��ٌ�ʤ�A��_�d�-�W�q�f�8ڗ;S���z[�pը����O�oT@���=ԙ3f�w��g9��m��!ֻӔ���eL�횞���1L�ν���n�Y��J�����5A�U�D���A.���^��sPw3��ǁїİ�a�(X/�In^t��z��K
�:�<�.ۥ��s~4������b��w;QgZ]�.��ki'x�2ܝI�p��8[Q�i�.�����׽�{뵋e�;�0��w3_iI^*�q-��e��v���R�⺔�w^�1iš|Wd
+����`�����b�sWz5�Q�sAެ�9ͻ�7�8�'%��Lu���62\�1�r�	H�O=�{��V�w��+ڮ����|u�:KԜwiڄ�P���*ȕH�܃�R���.#S[�f��]��
5����q�:֎W�s��7��n1�+��<���.�pAѧ-�4���:췳���jY�jz�SK9�M�>WU��Oa��[�]�8_�e̪�M��6j���׵�������
bǑ�\M�]���r��;�3���z��Eiv�3����o��֯m��k���6 �x���L���=��m�����4����]�*{ ]����ES�7�x���>+cC%/F���#.�z5�QKRES�V�jIһ�S$�IC�+]@�(>G�b� �[�^�kp�x3g8W<���d�W�o"T�!Q*�E$IQ��6 (_^���9�Y����Z�^"�N�Y��I��bf�K�hP�s����s����3v���.����JM��={��y5B�,ݖ���9:¸¢b/�f�&źŷ��͘��������8_n�nuA���-�YP�T��k��U��\�{��]��˘Wz�g;*�� �Q�\���UmK��-��hlS���o��{6�خ'F��<�����l��v��~��=Z�)��s/��{',_Z�j�8���V�����{M��Z��
s5��iv߫��"F���%����x���ˎX�dk�ڈ|.aJ�C�!|�hu�w,b^��ڊ�Jkx��S�V�������ۉ��?9F~�#�$k�'6t�1[0;k0(J�?��)��B����+�M+�o[�wCY�nG�f�N�{�ͩ;<{xI���#\�n:���	:��\�|�l0�j)춧z�d�t��H�@I+-��]|�o�@�P���4�ӽ�ةs���lؾ�<��%�i�$�H�d�U���(ԕ�ް�-��WĴlJ��l^u����A�u���A��4���*}pS�q7���'v�8�r�� ���33��)�%����s+\�D�[W�֦[}3BS7�`9�=#�)m2��.7jU����CdZڏ����]��������'4�V´3j-�yئWgf�uQ�=� ���'OBɡQ����e���څq5��"��T4t/i����>��NGx�;��Ǣ��9���NG�*'��e���y���G%z��}j1�D�T�ۼu�[^�^�ko��\N��>��q�u5�.N�J�y�pw��҇�fϕV>�q;��\Ok��
�h�&pe:��:6*U2�I`Z� �Lz�Y����U�C��pxç�q~�s���-eK7œ�fX������� y��^
����"ן���NNod[��0���-���~�]xo�����;*tݟ�fa�=L\u�z��:������o�������j��{v'�w���#�hx,���e�,�ƾ��hʨ�A���D7�*�Y��UF��D���Rh�o]�Ev��ϙu�9��G�܏������T�pW �*�K����Q���H���hQ�Al��2Τ�B���z��ü"�m`H�9m'�,��f��:4u��&�^�a��J]�*�	���
T�8�w>Y&
ޒ��$;��w��}�M�j�q�#��;�k���4�^�}�����r��<����2@;J��e�OhM6��Np�y	Dī�f8�w��R�*
 pf�O9B��S��+�9԰h����nf���f�o��f�`a3�L�}��Q�f�ƵMR�Q诗Z�$�}Z,`�a,�1���)�/0��pH^N����m͎�U�t^�X�¶U�E�؄��Jܻƻ�N�z�.��ܐ�}/.�oZrȇ5ŏ���_n��ќX,�fc��^�뱕i3t⭫��-łV.�`�]'�v��f��X�/Xm��p�F.����[&ul�D�������V>Y�q1�`�U�9F���9c__tr��('�,�b��fuu�f��8p��ؠi+�rw�a�m�|�2�QKD��ƜF0f�i�25�(N��	�رwmE��t7�P����]H,;5��Î����<�����)� �}�v;YNX-JY0���,v�}5B����Xh�����K�є!ѣ�ފA������<��{�:� r�Wd����r5Ն*lP�k��17���|VZ�
-L<� #4ґ.��ʹm������̝Ԫ܊�
絵o�����Lن��5�tc��4�L�Ix��!��Y:����O)wN��w7��R����H��bs�yz3wӣ�M�n`�7[��A��ԉ�fX��	lԻ�ܶ��j���c�[�ڭ�OTUǝ�#|��Wf֒0��X�ZaF��Z��S83�}m�}]8SV����p��̈ۮ�S��a�/�z���9ST�g��M	
5�y�q�]�mB�s�aDEu�x�|y4�e�/.ѽ���\`��Q����=�-;�{82xf�8�EE�&�Jޫ:f����M*���V)�H�J�h�k��������R�����R�E�;&ε�j��ۗ/�{nC���R*�]c����p��q�+�X�SH�vAFu!ۙT��ڜ׿rq��ʖ�^]�S9��O��9(�y�&���랜�H�e����K�X�o�C�&��&X��/�P��u��"�@!2b�5b���C��`��҉sh�A̭�t����Z�v]��d�-ăc����n��{teL�U��Y�`f8'Vjk]w]u�%q����*����51g]+�n�n�O�i��՝w���ݣװ��Ӗ�sQ�I��]Ma��a�N���ֺ��z�:7M�4n����)B��c�|����G��i�>���E��]�uf5P��Aw�¥})�I�s������M]�#& T���@����`̎�Gg�E�6���Xnu��^�j�0w�^��v�=�
H]�Q�N!��;ش^7t����p�!�-*��ʎ73sg�.�T�'tH똗�������c�u��w��2�]���*"�G����t9K���a����Jw\�=�c��^xn;���!�wKZ���&;������Y����h%d�x(����QDHIUU�w\V���C��$Y�j�����벻����^F&�T뻨�7t�� ��J�R�\q���&��9�"���
����(�w;�L�
����'..�W��$UV�Q2wq��p��(�
�j^�x��*��s��W�*=q��3����R=V�`�*Q���]q"���J��	H5��*�$�L�ۺj$I��P*�*���p��s��g�\������Oi�K���f��\��tGu·/*��ܼ/A*�9N��YZԄ�q0�+���R��;��'�q$�L0���U2&��kƊ��c��[w�1�'
��c�9a��r�;:��}ո۝[R%���\˶gP�����qjnrڔ�w��]w���>7�u�ܷ~ӟ/H�|s}!������w�6
7La����ǰ���W��߾3�0u�q�}��k��s�~�&�޴�g�=k����4���;�'i�"��ߣ�o͚�z�ߞ����@�K�o���u�wC�
�Z�8d�;c������N1Sez�m{-�G�a�V�Cd}��F�/	���`2���Tm\�}��x{|�F�Ԏ�.aa>�������}c��d�<l2�}8çr,��d/=��S�����^�����n�݋�K�G��k����]��^���x�ϡ��ԲxW�e����X��VL�R;�vtr�U-i�G\������?uǲ=�wE�E|����.�}��2iO�D���&����Q��mp䃡~���UK㣣���:����m��Ȅ�v�>�O���ݗ���=�S8}�^�+��Y��>�e�i�]@��W����j��FRt���c��o#�W��z�x��,N/`��yn�ez�uϋ���oz!,��q�;�f�N�b��ʽ9�T��;���*7<����ñf���WB���Z }��b`��HHe��>"YtR�C�_8w��~��W���f�i�T�5�wh�8h��Y�.i���
�\�@BN�fa];w���k0l���-������g�]]ۿ�S�U���h
髚]}fhG�t����S�l��9h����f�ǽ顺{�xV{*t����3A�j���� ylW�Й��o�o�I�W��䇐�E�5�1ܿzNW���s�j�vG\c�b�\���Idu��n��{��W��+)g�=����e@�r:]�<�>�q������\{�dEy_�dD�p�Ӓt\[�OT_�jh����ޯh�|'���R�)���[����s�x�>��O�V}�wY�����o"��2}���i~`��� ���	�Z>�[wᑮ��Ͻ4'����G����Hg�y�q���y�ϐ�2��J�ѝ�7�b�JT`L��E��-�ȍw\=�^��"��W�lgq���fO���w�G/^��iW�A�Q�u
�\�i� |L\�\M�2�^���r ��z:k��C��2�����N�0�+�����~����TNB�*]�dq �OQ���3W�>s���Tg��o���u�1���>��R������u�W�m�E�������;�o�.+x�l57�=W��Y�3�s���3Q�ڿQ�~�"|G� g���4�dU������q���F���8)Eޠ�ɪ|>���b3��SX��ud�(&t��=�/ ���(�n���-�S�S�%��7�}����7X�κ��#OQ����(H��cjΫ|��sw�A{�gr9�c(� y8�'f�bJ�����g_�ӂ�+��hdV�|o9��q��q�������h�?O�w�1����|�Mx��>�62̓�>'�2c�p'�X����>�t�k;�î9��c!�Z�~E�T����s��E4��u/�dN�`�[�á��0�����N�=�Lxk�2E�S쨮�s�{�UK=��Cꤎ>�/�Gz�7�4�d^}��ݳ0�F��؉��q��Ψ�^"&�ȨWd�^ow��|��}�Q���c��s�~��)~w\;#��VzrNZ��%ٮ��/���w�MW���mw��m]�$�K+��
���L���N���}���[Ƴ�$�۟lq�$�%<g٫�,񳞙C(L�>�US]�s����i�x��~>����Ͻj�V@^���*l�zx�h�M3�ʖn"ܐx|�b㮫�n��f�5��>�g����o���Z��t���W�lc�/Э�%��0��Q�,��� �;��W�>���SybE:S X͟e��[�O^��ugy�<�=����c�s�T;�rQ�|ITf ��O�x�n{�d`��9���N��ڻm�iգسe��̡��'c����݂��VLa���Y)^�HT�x���r�U��s�w�	j)�yD&{.�/9u.=��J㪰�]:�����+˔��o���n�3fo�'�]��1��L��Z��84qE%5����V��_���v���n�����؎��o�H�uL(T� �.@��,z��k]i����3�+v z����~W}�H���)��>����M1G�'4�W�o��,�.|�sD^W�ͭ�I�u���O�����I����-��ُ����L��q�ZL�~%m���Q�7�v���JG֝�[>@�k��h*r��X���W#SU�0�����O����6�T*����ISZN�j2�}	�|t�~cdjj���
���&�Θ�~�:@�bz��̭�k�)t/��R�`k�C� Lw���,�����}�-Wi����&}�;��*j3ubY��C�׷�?z������~�	�u���h���`�����u�k�aL�N\����en�s�gˏ��x�u)���:�#��@z��G�*'��t+�9'.6X:rj�ULɟM�;>\�SY�����,u��ZG>5>�t�~7��=�����ߟ�x�^�����J����F ��f������Y�}���I�g�j�Ό�U�6e�X�������T�;I�zE��t�g$�4Q��Z��xr��M�6��-@�tq�;S`n󺴍��ȥK�n{آ���g���Bku+��p��˒�zK65(͹G���G��;oU�T3]F���$�� ��h��Oz��{m�^]g5� 7+��v�u�)�yqW�U��r[V8����54�PV���o�ŕ:nd���X����_���K�<�4ׂ����#�9~�Q��ӹ�U*��P=��.��}�mw�z���vT鸲��0����Du�z����_-��Mz�iH仒+�"�����p|�(�z�<�=v��HX�ەIi8!�-��ڔ:���9N�x6�v��6|�����<n)��y���#}#��o����ׇd�pW�6J�,�nB��|��bRU�*������w\��{�q7��NB��|C:���m��^O^zҩ�6���כ����d�p|���q�����Bn}�H�G�=k��N��w���ǟ��S��Uz{j��_l�f��@J������I\��_<�V��~v��Y(�0�ut�%y��W�O��	ކ(�ɕh�>������-�6¹h���]{5�6fTz���yf�N�Hc�����>�"}�N\�X]HY:���eFK��5�߂�%�i�y)�w>�c�ǯ�r��7�k����]^u�}�W��X�d�,�e���[���V����v����vS9óP�[��/�t����%o�s�<�O�b��m�h@�g�Lg���5���d�o�\k��ɧP��[wM�ٷ��6fa�-�]t���#J�y�L�uq �:v@�J����' $U�
���V�O]#����*��{k����g��wK�|��Ͻ�wF��F߽@w�]��>ɓW���&z*��Nv6�N��>���\��W����)��ʇ�'�cz+�VG�.'�Vsgf����!u�tyZG����q��u'�F��&�<tJr���ǯ��G�:�v1�/i(�z��L�.2��O�s�G}��Ϯ*ƍ�D��w,�n���b沯NEJ�����n���ӹ��7;o/�VO�z!�W�r=u��D?U�²�<W�
�fӂ�|&�!���.#	�4}�2+��vl��[�Vu��D��co�!�~��^�q�j�vD=��9&�p}��An_(��e�fR����B�}Ѷ���9P9��y}^&�=/�����?���;'+�D.�����L����r�Uͥ悯k�3��	ꎸ�U,e�����Xy���9�����{��+#��<��o��ys9��z�ѯ@65�) �D@O�E��n�2>�t|n��7��p��G���g�Xf�jW��&'�{�Kp1e�*���v.J4����/L���m�k������B@���W���o4��uҔسY�k���lU^!��=��T��u���X��c�9�7&WS�䢘g�]�P~[E���Zg�1����9i��4�w��p��j�ҳY�vQM�ѣ2��yŸ�<uk
�x�Af<��>�e� j[�.��!��K�w�a���Pp�G��&�ҽó���d˺0%�[�׶�/雋��tc̺�K��6|�;�}�L8>��{~����3~�z�j!L�.��8������zm��O��pO������+��ǍG3zѨ���[g�H��x�δ
�sl�,�9[/�u*��B�Vď]{օd+��QϹ����m���n�ȟ��P�u�K:�B4!7��޿(��8vA<=�N
�)�q������>7���y�ы���h�>��k#O~�2ͨ���I��@[�\V%J؁���k��S��[���w��[^f��G�h�w?ZGzo����?5�_���W�a�U���ϰ��ΨZ��N�gոe9�u��f_z\�3����}�����ᐝW�ȇޥ���@�Mf���i� ��]�[y^��.܍�^�'�=zqo��>�>�S�'NF�@V��d:��9��~�^s��uú�g�$��I3Hs�m���ٴ�{��eG[���3�K93����&B�d�w>g��Gr�V��ex����Dg�����P���T^�y8��	bx����������;x��Uk���VѮ��r��+*���OvFu�Ó�4ɉ�����%>�fX�3�T�鬥HTW\�_V[�S�5��(C�9r�ѳ��^X7xp��y��d[s����y���?�-��U>�t<�:}@=�нO��}g�=�{�f���a���[�}����u{ma�=$d<X����tY���q�x���8 0H��n�oh�|;к���:�r�3|b�vT�qe��� R�Du�*�ҹ��Pu�^o�Eu_uWu��ҽ�G��J�dw�|����!���Ǹ����rQ�|IUf	)W��_3�G3�� b�>��m]�+�r����{�q7��N/my���x�yIP�W �SP��s|�Nz���S^���-�;u^�ʼǌ�/t:�G}�Q>��r�<W~��n=�#+�M33�<��5%��4{3���l�x�|��_p�:ј��I��:���~��:<���D�սMWa���'��?V)�$���*�҆2&"�W����T���X��m��[�*5��%��uZ6��4V%�+�O�;9�^|�2�u2Pd���^���e>�Qϫ]>7�X��`Z�<7nn߷<mzFDgu܋��x������|� �w��R��B�{L?��������ݢ��v��*9$+t�<���Ժ=����A�e��)�< 7]p'��
G�5*��n�N�S�3�wR�.gm�x'MWW%a�Pr�Vԁ܎6�[����{����rh�aGOE����{+*BS��	4bj�����.V�&m����ҐXV���^�C�p��;#)�Nюp�z7����ϛ�]��(~�	�p�hW����O�`|y6#z���-����^�,��_�����E�����mexwНW�}�����D{.�GzrNGg�5UD��s�:� h�
�p6t;��H�>�p�F�~7��=��k�\���W��^����@�+�yT��[���g�ah��'N���ӡ��e�*�92���~ 9^�S���E�٬��I�����ڽp�B���gJ'0-�3���U�Ϫ]瑦��:v�k���o����[��l߰~}>����:�nR����	��1s�%�u�k�<�,ℱ�vݬ���<o���K��y�3��W��z��u¢eN��pG��Q���S��
6Ϩ�ϑ�^�讚��ϯ�p|n����#����������ׇ���U�蚊�<�v�8]�ܡ;�!��U�_]{Ō�]�����n%����^�����C=q�W#U����T�wX��=5x���2��n��l������	���#���3�Kܾ��xTc�}�^�a�R���mh������Gu��r�R\���뚰�n�*�`�Iu����ɵϞ]�)����,��;`\��X�2�l��F6�)U�:�)g�z��:"�jC]����ґ ʖ.����B���<��u��5Y��a���JlO��705�9>/�x!�Խ�r�S2%������I������Z�!�0���x���U\5�������~����&��t�&�(��T�w�	�b~��TU����R���W9����/wu��p����ޤO�zp2�<p	�ӹ��z����T*P�N�ϸ�����nr�F���+ex�����}�k���Utmyׁ�DW����	~��iK'���*�q�]V��q��o�8s[��8��W�}Ǩ��h��|o����󪢞��t_� o�C˰iy�F}S�}]�Bdk�W��꣊�Ad�m�w��Ϻڿ"�����!?]���Ez��xj��"l9خ��*��D�ue�^�q�ĺ�,+:�Vx��N�=�wS�q�O׽5e������&�S�ϫ�{�=ʩx��U��k4�/eN��'v|&]��\-����q�k�����P���Z�� �ή�O��s�]k=�?U��vO
�eN�9�a��P��qq0��`ۗ�v�z�'�fK�9{M0/?\�Ey��Ez�=�")�����Vt�>��������o�_E��b��L�\�2�':-
��ɖ���F�ݝC�vXXW���n����1#B[[�����
��m��sF�p�N�3��(?"�x���۔An����hK�c�:��Z�Y��5���b1�^R�$�j��n�|u3� D�r��fZ�J�%�S�Rk89P<��%�J�b}�����ݩ3��k�B{;e�b��y��]-���u�(w3��:=���Q��)qQ�ʽ�8�!�>��L:�u�w���#H��ʙ��j�"�!H�<k��5wk����t��̠��ǯv��ո4:S9�K�8Y�=���m6V.2��8��M=`w��e;N0�r�xP��5���U斉ӓ��� �
t���uެr���Z`��X� ��7*��{w�i�P�֓�����q��go�����JT4��u��y�s)�[>~�}��tzoz��^��ȞqS(wv��X؅^�,��nY1�Sղ�6+[L�)҇���/3c&E�]u�;�E��#�r��eK͗�����$��g�@�*h����0�Vv���Y��w�@�Z���:�V�]����}j�m��r����t�^�U23�'Z���"h�g��;�j̶�Uvv�d�ן3F���9�����d����i�w���.�go>��>%v����8/q�fԼ뗃F�#�:��W\����Y��w,%�8��fe-����2i�ʟf3ZA��Ū��דf��(ې=n���X:�2�k8cLM��P[zu�,�y�����9�G-a��p�<�W;�)�ؖ"�$fT7�3����]�A=�J����[�魮&���s�7��b`��
���6O cQټN�9�Yֵ,�����t{��%����^8fud2p%7j��բ�7�4,rVT.�])5/�S\�k���l�l���ţp�(���̮+���-r6�vVn�\u[�2��������B,v�%��8:�v�S5w�g��ռ.�Y�<X�wJg�烤����ߋ�K�5̑c&OF��V$aEFQ �3��@=3�ҥ,]��ЭZu�*	'd��ӽ�3�V̮r.���E���)/���+c����H;0k�FD�˔Q7����*��o��Z2snoeO�]��a����.�jc,��!�����.�x�^:y�P|W3u4� �5�{�<�_:{����"WTP�d�l�c�w�W�����.���X�t�7�S��ڒ���Qf���s�����Nu��n�"j�t�(�����������2F��gJ�Lٚ�HJA��� b�'��ٛ�7�pG��䘖C�Up�w���!ÉN�S���O�;��[�o{y
��Gv�o5��,�Z���|Pdm`���h��Iʶ�i�.38�t��!������ױsڼ|��Xl-�uӦ�1�D��5w����Y�Q �1�di��S�m���NQ�f>F�/�oT=Z��߀�`R���>�s�"��"�g%��|�<Ј���*^�ٞA����tr�����wA8縅:�^�zz�$\��"u�����.TP:YWf���R�w<Ԋ�W���1Q3ѡaaz���^na��܋qJ�۸Dr.����]r��G���+�w9r�q��ͮ�R��Eb
�Tz�Ne�V�;�����3�p�wr0�]2M$	LD�!\�I�����"0I�ܼ]s��a�d\=z�z�:%z�-�$I�i�N껅Duk�@U^�A�s�:9���^u��.y����9{��	�ĩDˤ��rp���ꐅJ�-ۻ�{����uE���v�F���^By쐜�1+�<�
�U��"+DN*)��(q�Wwu�G��C�D�^�	P�e���*����{�gJ�%�WvỗGUjtV�㑉�&:��*;�)�J;����E�V�����ZP��HN0R�Ll���H�2����3B�V�s���*�2]%����\�Yfw ��͑�./yĥ|�"�Fpg^)J�n�f�6ݻ�7]*�Ο]�����9��}��q���~nx
g�>������UMr'�M}}$�W�<=BUC��Kj��z�Xy�W��o�x�9�����>�v,{�)3S>ǲ�Vz7�f��lj�W�X�>E��n�25��z�M��߇r:�����Rnlb܃����#������j��|fه�����`L��E�L��>�u��*w¦c��.���]i�����ѐ�י[�z��~�A�^�P�\�j>d@J�ω��뉕����^��;��9j�/�r�>L��Q�ＫB�����}����W&��#*=^���L�.�'1K��2d�>�gG)�G����>��jf��֌��~��z�>9���7�Z9�ey.����*fT��K�MD����H�]HV�+�3�s���3Q��j�F��ȟ��P�2�f{iF���>n}�{&�fF};����8+)�q��Z��o>�O�?mG������V��!t+��V��>��}�C����d��Y*�d���,\u����x�}�^�R8S�j��=�=�v�n����,r�\wlg��N�GI��X ׯ��uV�����:V���]�H��X�ف�M&��?'QPw6��j�j�z�+V��O7;p⮺��n*�
 ���,�g�%� (/r�L���P�yܦ)��4z+Y�C�+>�U	�V
��Q-g�Cv�T7c(�n�1�;�r̿��vos���h+���b�oo�!z�Ⱦ���qޫ���Ш^ʑ���ݿ���:E]�~��3=��Su�>���ߙύJ�t�ѩ��W�:��9�~�^s�w\;;+�FzrN/w��2'�+L�Nj�	=��|W����Ŀ��ϠV/;���w/����3�n�-���ƨ��~n|��^�Ib�,����Y�]z�b�9ΟP�O������}��<2�ʽk'�΄��P��=4_�W��U��u��ط$����x��3�;\�z�Vg0_Bz똙���j�~@�n�W��O�yǭ�ydA���*Q�,��X yKU�o�q�B"��zE��>�?lh�	�V��3��!��1�*o��\�k�|IUa�����.��=��q*�eMw�O�g|Vo����{�q7-ߴ�/my��Gz��7�$e|�V�#�g<�H�E���w����� s�#�����G#q���n}�H����?up7�[�~[^��Dt@��EytdYFB���A��`'��+~�}������~eZ3�%�m0�7&��̊��<��;��5��R�/�\�ؓ׳�m
��w6��{1Gu�z���T�V�"t�o+h��2q��@<�54vA�#�f5���l����tE�Y��̍i����s �Q�S4\�[�#��|7~y֍F����1��οx�VSY>���Ꙟڼ�s�zO�h7�"��ND�o~D\��46�|{`9c׾W#}]��f1g޻��sT��ޯ%7ު1�^v|r�<O��uaө�H�z	�믂�4�߶~f�y�L�w5�с^zǳ^.�>��v�1�~Wr.�x��{��;�� �z�A���z�L>#�0-W��q����d���w?s���&��jx�c!�Uѷ��\?_��Y4+^T�[,�^��{]��.�7R���dgLo����\�|��S�7���'U�rz��)��ݕ�ˡZ�nz�8܌��[����)�9/�<�9,z�:�Me�5/�Ӛ���vڸ�C��qr_�x��S�E9�^��@��A�w��G��5�)��p�'N�φP�:��:6*U~*sfX����w^�=J�\8�5מu|փ~�}u�=���%9�/�3�#�wAb� �W���K�<���X�E�헑5y�+�C}z���x^�x�C4��&&/n��f0�h�d4�y�3�,���D��i?� �Ł��j+qM�u�.�,�ޘ+��m�'�3��Z@0�e���g���W6��~}x0��X)�冱34��� 4D�ə;Xҷ��1n��nQ��ƹ6�ᒡ��P��z�xuv!ڶ�q[�B�t���]�s�j�*3� j�]؇�}�"���w=���Ͻv��ț��dg�Y'NL�>��s���{9�}�o����f��Ӓ�-T����>�i������~u��u�E��¶��:�f�{�_�=��@�?����q�I25�����װ���|C:��Ҭ{^s#'���g�z:sǮ�QP h:
�Q�R(dj����Bn'޴"��;}����A���q���Qʽ��9Iҭ���}�b�\�j�� ��H��#�N�7e/t�؟��G�'����=��>ζ1���[�(�tt2����wC�L����_��uq'?L�^PG/*~^����[ޤO����ɸ�'�J�(�o��^=����8ٽW���Y�no��o��r+��z��?�f�����>����}��L:�
�{Т����4s���'��UC�K��"ޑ�T�˰�g}��y�ѿ�σ�p���([ܣ���L%7��9�X�a�50����N�����&~`�OŚ��~'�ve�lln�N�'��k����\�(V���b㓘��,l�㽵8T"�:p�tre-W�<�r�%�h��xُ���{m%� ��G���A�"��)��ز��Aʒ_WբE�Nx쾁`��|j�6oJ�8s�R��ft�3x�,k���=��[Ӣ�_��~�&�L�}B�Y����l��O�_|S�oF��;��O����⋞���b�^�{]���U/��z�kJ�������	�0ϴ��]z�\�nk�]���+@
�n�2!ש�?V���V;�ãj�[C���ʯY����v����V�*�N�6��92�y�� ��됢����}^�z|��ד�gNI��Ύ��O�������f�3ꇵ�Tv�}����z}^%x�k�\{�dEy\mW�W{ېd�:�sy�Uw����.ܒu����J����s[<fw��O��K������]{険�M����~�[�K ��li9 �A�"�u��WE�nhNپ�Yt�5s܇�:ȭ���W{���ǳ�ۇ�p��0�Gʌ�& �2.:e�9���>�ڠg���e�/oe�;�=�����z2#�k̯)8{��Tu��<k�D@�3�*;�ϧn=fM��ui�q>���+c���_�������}��y�ti+�yo���Z���}��ߧ�1<��瘶$�d�ahK�h��;����1��:�;�#��yT�y;�����A�~黖���P�k�묝��_s!�'�L##�j�؝�>��sf�幕�ru�]/�L�1�g���Gl�>V's@�׽��v2�qr��2��G��p�)b�:�F�5�Q��~��Ox�ޜ�~u�9ӤǼ�*��\�έV^���>��f{���M߅d+����/��|�F�j�E����`L����$/wۖ����6�	��L�CǧL�z�M��U�42+U{��:|n9���	ۦ�[����s��S�1�^vh���7�!��$�Ȳz0���1Q��z3mW�i1�#z����C}��,��:���]����Og��B{�bFDkʑ_id��\���a>�<�]^��ޮ��4l�q�>����ö��9z����W���U��~����йX�Ng�hW�N����z��~m����>QS�W�_`YMz�x���~�s����9�uq�Z/�Tb�Yƾ�[W��眗���:v�}����GV]��%x�n2e���^
K��9�z�Y�P;|h�!U5o|��c��>������v�e��3�uO���:s�l��W��W�R=�ݯ�gnz�%��<=����g��;��#��:n�������,J���V�x{�oFSH��3�Q�cn^^�o��y��iT,����{X�򜭭�}�.�������W��@�V-%g��.|��&��Щ|W�.�q�����Ь�D�P��C�z�c�,]��֭��4њ�B��X�n�U
Bk;GT7ղ���.K�"���9�G�ǩ�����+>��{��XїP���2�M�ls��)���6K���uӹ��d�]>�ʃ��Ѝ���z7�|�?�}@>�~�=�>��U��,��p�>>��wT��y��8���L_��y�����u��Kw�+����P�ǔ���a{-f�sCۗ�'�&��lg�>��zj\�%�`�^/#]G#�ʢW�>��G���*!�tw:��xW�N�z�/dx1�5�7�4���2>��A��1)V���P�7��Q����N[�@N�����O��5����3�M�S\7)�<jF�����ϐ<��ײv7�9c�C�k�`�S�غ~��jӫ�������+>9ӌ��z� L:u"�OW�f����}~�ϴ�t}@�"�}.�o>�c�ƽ�^
�޹ʪGB�q�O��:���u ҖOP0��P��\���:���G������q��s�=]�;W��o�TW�}@:����j�}�*A>ȃ>%(�q6ȿf�Z�5���ه]J�N|�Z>Ga)����^�#��@z��{��z��>����NY{q���+r!r\�9�3+�՛�v�����qH7=�\�/2�ЫK+z���EP���Gv]�2͊��֢���O�D�����'����9����٬b2�F�T��DeaQ�\�Qi���;v�� ��J���K_I�7��e�-�uO4>3��W�� �,v8Z���s���_�ĩ|N��R�o��w�u5�,vmê�Sf|��u5Շ��G������՚Pl͝Da��e��?N�fr����_��R��~�v�I���=���q���`��ݟ���/����̟dU�_JV_��r*�qB���_OH�����ϩ'���^�����x/?_�ϫ��u(f�y1{S8h2}�fh���ףj����Y�9�q5~�FWS�t� �Uj4��E���G�^^�CÔM�
��R���N&�1�'f�����$�#Y�A��뮚R^}j�3Q����G��9����7�����þ޼8Hg֮=��jUf$&�z�Ut�I�P�P�I�wG��ި5�7~Ӌ�<_��j;�B�$j�=���|,�Fk��S�.��Q�P@�,|ƙH��j��~�&�zd)��u߰ᜬ��B�X��.Imw�G�s��_���ި9�aQ(��	I[�"�g���;yrL����~����CAmR�����&��8\���d��߯ ���~6���%�a��`�#$�fF���6�pi��b��OWIyu&�����:bg����ƍ�4$Î�=�V̚P����8���t�\*C����d[���z��ub��:��<Ś']���y�������pec��j}��3��G���ɝ:dZ:��h����G�m��}�0�>�9{��>�"}�Ӂ��@b�r}҉�� ^���<��q�^Pא�>*bn}�Te2�5\/�y�����Eyρ�� 7�����1KUz�l�c)�W;J;�EN�0�|I��=Q�8�p�����Kg}�Ϛ����ڷʓY/Ҩe�mwMx�߮@��=i\�iF.�c���N�����O����nF�z��\��eO*�Q}Ǹ)�`��g�OߦЛ��:��!id��d�T�
��:2):D��h�b8�/Xޞ����=!���w.�v0�3�)�z�������ٿ���/h��ð3F�X���۷�j��'e���l��^	ש�p�Z�?M���<+=�"�d�uk��b�����5A��:�vAYQζ��DT�y�� ���쑎���g�}�Gc���"��fe�3��Z�7{�b�ȿ}��F�s���3)��/\¨�.�7�S;��4xk��&�@��G�������^���P�Z8'�ȓ������J���_�[<fw��ϣ����Q�3�M]��1�Vzw#+�ky��
ɾ�ݵ�z�mwƲ�Θ��/-�<d�=�+K@*ZV�k Pͨql�)�|"�Bm����a���¬nd�Z��:u���(�b��=�k7�K�ze�n�	����Q�}wBd��u$�wi��5c)F�d�ps����>]+�g޷q�o�B6
5	���`"�����RY���-{��z	\N[�t���T��}�և�q�b����P�A�f�.J5��Pe�/L����ܿF��s�����4��T��D�}-��dy�y���GJ��0,�:UO(��$t�.�>�T�G��x��̼�1�\k���W���Ѥ������T[��.*��zc��x������@ =#ċ�:�q�-n�G#qѨ��M����9���7t��1�r�7�0׿~���~���5��'�6vH�_��R������#Q�	����D�ǣҵ� 72f��h{d���g�[�a�9��= ����J�ƆEj�q��O�������'�3:����=�o]ы�Mz�����Q�n�mez��V��2�4V�g�Cxw�ߗ,}�kѽHu���C߮�������=~�+^T����@�����}/;��:��;&��SL��W����Y�w_���m��d/Uy�ޯ��G�hR�T���B��3ޥ�}}yA#���<%v9�ŪvZ�+���mmɧ7���WO'�,�4�Ϧ[��
M�(]�u�;=o���3�jN�o%N�ݼlRB��/$�kkY�u���6���S�S��g�07;�33�:r�}������6�+aq��Uգ-�{�iR��������B���m)Z�]a*	�7�~�j��k{�vL�b�ł�C��Ën�)�A��Ԝ���7�_A����ӊ��]Ne���|�g�qdrc�QA�Vּ�f��5���t���i�/��Pb﹃�e���7S�ᮅ�+-���؁U�]���,%�C����B�(�Zۨ��{K�)#u�c�v����
VM�.� �Jghj��5�`�)WF��
�ꅐ��J�����.����{���H��E4��P��Su�i�%�Ψ�K�IR\�]mʽ�2�u��Y�S��)J�S5�6s�ʙ[�v.-�bR�����H�mB�W�������R�\q1ՎXUf�o 
�F�֎>]�j5�>ɔ�r�_n9Ʈ����j�:{ӆ��:��[pK��x[��x�-�Y�O6��9x��Y�rK�$o �[�.��":�r�l4L�f�\���n\���_v�GS�i�V1�:��2ܭ���~0�親�8�O�C�L=�"�Y��	B�:q�ZW�C�+�y��BEuv��b�V^���ĄJ9{��G�>���3z�S�/&�6�;�x=Lp�lU���纻T���5�oDh�Mt��	B8c ]te�tiLt6�|����Gv����[���o�D��ziWN���:����c }c�쥹�2�:�M���yf�ї�����0� =7��)Ś����[�71j�Kr�:�bg6*�0k����d]���ZU�<j�|2�k,�"A2�戾��N=!cUt����^A�՘���d��f��(f����j] {\p��E�4ݦk�)��gAp\ڱu��*��L��۴�ޤл�)-}[H�돤&�	��_B�qQLGu�쑸��b�b���5v�ϥ��ͬt��Y3���4J�ܷܶ�%�3�j�,.�7Ky�m�)_V�}u�-�o�Cj�;Ò�����y6��,��c�,��!�ӕl�G���^�	�Ӯ�w��)rx6q�H!��s(���f��SJԥڋ��!3Q���
=�ըn����n�=@Cg�s���rܹF�oD3fc�:���[��`!��ɛU�m��Y�7�.���������W;{�-��c��ɴ��l��-�u�$�����*�O?����6�ef,�����R��d�����p�+��,�4�wk1�ܮ�+\�@�*u�'ͬջі�\9Y%���Mf�T
o荰-*Fs�9W#�F�p!��ܒj�b�Pi��vl����҅X�Y�&.��ˤ����Ke��	Oi=.ҵ"��ͳy!�쓟�eF�s�~�Ty���I8Z�Q�
�z���K��j�Q*��#��jt�+�,1J�Z��
��fȄ6W��.8I��R���T �ܓE�)WE��z�E�ȱfG��jTr����]��;���E"U(��Є]�A�$:z��I�㙚M6E$iGKG;�x�����#�ȶz�t�]��	Ce
�:��EwT�r���JF�$�g]L�G\��'v�W����wIԓ�jIR���x+��
:��K,��r]<99
���R'�:��+=��"F��j�ww0���s�$��Ӧ��t����y��.��-��Y�pu
�d��̃ę���:Gs0�wȩ�жnK���	V�h{�C���Du]�+�:Hd�QY)HE�z#����qَ��M��U�q*R]v�{���bF��ʗ;����������kO �,u*���*y��$�6D����2�4�=$]�E͝�ꘌ�I/:����� �A$Q	�n��T�\h���\��`5�LQ6�"$+I���u��6���HK���1({!}Ĭ����2c;�J�\ ��]ݏ��ں�"�a~�&���A���Qc/�^uU�s:�P��>�^؜���A7��~��^,�Oֵ�.|}B97G�"�pA��f\
��~�~>$��<��7*��_���/ѫ�	b��Xl�ޓ�2�A<}�^����9��wni򽜪>,�f�t߸Dv�G�>�ϼ{!�\wdC�F�U�B�ep��Z|%lo�>v��J��.y���b�Kz��<�U��ρ��k�r�3�o��
,l�K�@�a7Þ
^�3ю�z��q�^Fmyu�z�s��T\Syb/��z3}�w7���c�R�����Gn�{[;�=���2��7��z�/�f=KU����/]T�uĖ��W���F��|o�H�����S��|��eb�n״T
'�@�R�	��x�2�^F��F��~Ws�ZG�<WZ�gO~�l,[ƺ��޽\^�tFR�fQ ���<H�J��+��a�EkU9��*���p��%�ޫ1⳯�;靰���O	��[��|��>�=7Z��݅�\�1���DV��"o:�v����E��2�/��r��ΣCR���{83�m"��ˡYyG^���]bU��p�Q��-ؖi�K2�떚���i��:�гyN���(qK[pC��"PS������ذ�0��o��H_T;՛ԭ�GJ��R��F���r:�W���g�x�%�b�7N�T"��&�Oa��fj�+N��W��]5S�G�[>�W���w��#���]ȸ^u�n#ޟ�ϝ�b��R��ITW_n5����9�EY�Ǯ�O�]���x�wT`�������y��8Z���=��[8�.��՛�Q��'� �\F�[�S�ӊ��v�q��on.9z��>��R�}ԧ6`y��q9^�W^�%�ԎMz2|5%_����.%K�t�/��m��,�e5����=$�������G��)^/�U?M�H�fp�"0�L�����t;�j�Ό��U��V<��h���o�b*}O�>����Ո ��>s���+'�cE}P��8.�M(�x\�3������^U�S/���k�̕ j��i�^�:��������d;�7�<�����7e���^�<(������u��>3u\�;�r�<��<��Y��;��W��W�����E��d��E�����io'O`q����d7Lb�I�)��kwp�W����/s}p���R��3*Mz��������}|���a�&D{-RԚ��J%�3�GZ�g�<������� �R�{Y���co4�W��E�ڼ���V����륻L#m�}�w7��_Y�B��w:�ؿ�>fKD�g��"��-n�Ԯh��2��;qok��7�(�6	����0K~�@_�t����t|n+ި5�ߴ��x���������#�C;���A�e��Qϔ<��J��-�3]�x�EKIc�#� �z�}���O�so�������*�ި9^�f��(�8 %G�D�%��%�����X�[}W]���C<���S�o�Hh>���7���MǽPp׫�P��]� 7w�w�+��M�iH)�����Lzw��n=s�v�5����?*@7<K���d�G���܀��^ب��)���f��ԯk��Xn���}j�E)�=|�����F�ͫ��~� }����+��m]�Q�Fw��>n}�ѕ=&j2Y> �x�lo�O��gѷKǨ�9|n9��=�G�����[�����C�,l�>����P߸�&M|�SPrX����iо�j�+>�qŝ��#�؎��wQ�.��T�q�|�ь�ފ���=~��Z^á��~��(c�����ߣf�;Ch�F-��r��礯G*a�mޏ�����_~Ϣ\ɸ��ߥ))�໑6��9���������]��΃��$�i��q�ĢAVpʻ�R���َ��³_mc+��'
�$,�F��>-�y��shdi��`3���5dX�L-� ��.̆orށ�h��+�Fsಊ'��t+F��G(@����WR�J�[IWz��z&���T��w>�l[�wᎽ\̿N�����;gC�=�#;3ds�B@�+��7�J��xe�|W��۾92�K�> t}���#!ܿzN}^�����Gz��A�D�t����^=�=}9%�\�X�]���T+���tg���Tt��z=>%x��w5����Iʧ���Y�n�u��Z8%O"N������-㮫�,R�,�k�Xojqێ��܉h�=���j���۴8�NC���dG��y\P�2��$�,	ȱq֪|mtfN�����K;/��w���]�bm7~3��7#}A��~w�7�(�r�%Q��[��}v,��ЏE�R�k*}{�#I�ӎ���D����=�2�������˘[䣑1�&}2TS�n�	��� �θ�=>�{��j7���O���^G����������gٜg�X2�^�Y�^���>��gK�&%��o��}�G#zѨ���[dx�xҽ��G������]^<��/h7Ӏz#��e:j[6zH����
�t������.����ز�H�k:?V,��,"~�Z1�nL]�+��U�ރi�;w4�2M�c���s����$�Zc7U�=zút�)��[Tz^�����h��c���qry�"�㷋r;6�2�)�Nu<�&��0+�ݤEd�o���k��k��)%kރ2�9�6��Ur��]�}���>d���>_7`x�$������J����ߞ�,[�O��4 IB��\���y/c���Gѽ�#���Z���7��{!�1��2Li���݌}#J�K�����40��ժKk�ƪ{�=�Z�q����wzȆ�wB��:���ByM��d,�l�r�ִ����%��W���\ӽ�(�}����v�߆|�U�q��o���29X�W;���ef����Ħפ?l�;@��b��Q���`Yzw�y��g�:��9�~�^s���i���9��sb����މ~Yz*!)�9},;�`�t;�˾92�J92�b�=�h O_�b���7ܖ�N�'�m���B�K!V���мNS,e	�
���xg�.���ӼԌ�)_�k|�|�������t�|Dz��=��\wc�F3�gMO�c+�g���S�$f(]6֥՛-Q�ժ�<�.�=�/��C��{�]!�eM4���!�'V��F��oN����U��>�=L:�t�eA��7�!��V���;�����l{�M��JVǬ��2�_;���c�p��h�ӫ���V�ͥ�� �VS�»YZ^l��+���hMҭ��r����c�|[j�$��}�YL�}�k�О��ʟQ�[��	y������ז��GF��OCpO��W�|a[)tƵŉKg%�`.p��R�����0���M��ݦT�Z�]��{�&�[�i�^��=����2�Z틹+.�Y����9�_:���Lm�d�G� �ԹKu�o�2�z憢�����O�i�a�q��_�6���ݝg�%#O?I�zi�D����S�"b[��~,byc��dW�}���ٸ�/`~�޶�dg[g}3�M�{Ύ?�ߊ�#ߔ��^��T�~��w�Ll�uH���9���Ң���|��=��W���+>#��-z� K�RB�OC:M�AŲJ��kQI�Z/�+5u#7����o��\Gy܏�U#�^u�}><�w�	��:yTI�oI7��%I�g���7�yQ����r�������~���y�Ѹ{���xh�wxzv�������Hu�Oz��̃�%���l-�������S�=���!?]�=�%{s#��R������w�h�t��lh`�J~�^�tmxt���'s�˪T�<{���E��]�sFr��V:���u5�|=��[�;��Y���͔<rp�߆,���R�������D-�Eǽk=X+Y@ƶ���y}��ia�K�n����#p^���թ��Λ�X[�5��(Ěa]����n�(��p.k�2�l�ɶ�,��N���s�K�#��t���m�9aik�wx�]Ծ2�:�ݸ9u��]][�%{� +q��!�����ֳ�������1Y��p�'v���Y�����&s/6�U��c�j����@7���*1z����o��r+��u(f���£;*t�rޓ2͹��,�g�A{���Xk�>�}J�����]�z=�!Dg����~�,�����_���;��W��U�"���ʐ��x��[ ���]5�/-U��wp�z}�o�x����'j��ϥ�\��=J}
�!���pW �*��I��e�?@���M��wG��ޫë}~�^ظ��=ϯ����B>����T=Pgv��( yTA�&
��7e��пa�>��viޥ��˻-�g�P��p��:\}�UǽPr��L%�p@HzH�ɚ��_ml튿Wuh�Β=�;�;:�~�8d����>ζ;a�����ꃆ�=^��FJ/z��Q۠��L�������x�	�bg�u�������\��~v�z�>�����6�~�Urf;�1�3�}=�����Gx��"n�_��-��u���f�[U�)������%֮E���韑�]v7	+M�_E6f7q]�n�EWM��;6�1�6Cu֫f�bcf&V�퓅\�}]'L�޷,��Np"�x���י#B���ݡ����qH���r�}��[@c,v�y%�n�vL�b�
x��g�Q��3_m],E��=l#��B��e���nM�}S�3J|O K�ϊ�O��dm���9�_�~�<8mC�,���ΊU��ծ:�T}�)�&��ޠ;���W�}�&��*jK6T�:u�~_3ѻ��-��;�Ժݭ�}�n=�޻F1���Eg��OznN�fl��Y>��F·q7�W�� �xg�o�+S�����(�9���wW��;n�xb�yg���x�ޫ�6�P�^ʜ:9�OG���>�9z���,��y��9K�EO��܍W�ny߃�N�)���g�X�9�<6�(ɨɫ�Ӹ�ڲ���?Fωݸ3�E��\+۾9S/ļ�^ Tb��H�r��3�{5�ػ|��
��|?UW6���`��
�:rN��%������B��]ѿ����9>��O�㣽�zN9ۙ� ���֏w���x��Z����_�^�G�$�%�󠖏kK�^S�,�\%L�t�ٜ�}U5є�sE{E�s�ې���l��n��>3|i�(�[�Q���X����N�+$_x`�S��%K�>��<n)��7����>�G����Pg��ǻߌ;�\�k�|IQ���7���F��k2�7P_�u�9�6��H���q��9��!�2iɕ���k��;0u(�1)����H�F��àY����)[X 
�A(�'8Eʘ��P=���\o���g�Fu���5�����wLf�Dr#���ъUu�N�%}{���eZP�;�s��nTk�������"�^��=�2��*:U���N�5�gɣu7��&����/>�"�A� �-�g�x���5��q7�,@z������T�{ީw�{���	|1�5���	���.}`�٣�"b[�㌴}��r7����m��Dޢ`&ra����p��};Z
���2�R�5-�Č���B��t����r�D��}��,=�q��]��:����u?O�>9����C�~sNfEq���Uߠ�aտ=�X�Gf�Φ�G~��Z�^�oW���2=�uU����h����ý�>�$�B,��0�J�+�!q~�;��{xǣk����|k#��:�ކ2��{��c�P��U����@U�Em�x����Z�5cw�	�0̪�;���_��^��9��W�,��x'��hv������O_\��\�}O�mBz�Z��g)��K�n�?i^!>'NF�~7�m��ϾuU�s>p>]��S���~k�z.��]D��^�F��t�;'P��[�#�a��3�z���c���C���e��pQ<;hgL�]���v�[I�eЕ�n\�h�d%J�Ķ캤	���,�p��&75����D��]��U�秮�� �u���,�Ε��J-\,V �9殦ӻW���9Fi֫��� ��K�$թ��BZ�c�C-t�a�;̖�t��qӟ�C�C��u��y�%���\΍��:���%�����K!���+����C��V?ncy׾��S�������?�x뮨�n�ι�;e��pe��dE_�\�zv�������fS*���a�GU��}^^z=Lo�>��T�}�7ţەN�Ϋ8�\�}V�Z�߳[~�(�A��;3ҧ�k*����4=����D���H_�����z�F:��zn����.א�@�(�qD�T�O�0.:�x���{�'������s���UFX
Ѭ��֫}��c>��$eB��P(��r �r�n��l��]X�e�TO�<�O����6둬��IO9�4���0�rE��L�$r��q-�q�_�j���J5=�[�}�>l��c��M�g���߽3�M��Pv�S2*�^����w:�g��h�{;�*�R�ft��m��=��>���&���>��}8�y��2çR,t�������f<�6����w�ۈ�b�[��qY)t�G*�Q��bӪ#��KA�_��_�`�1��Ƀ`����`����6����o��l�X�o�6m���cm�������6��`�1���`���`��0l�z06��`�1��S����6m��`�1��S����06���o�����)��(���o��0(���1"]�窐�R����Jk6�QB�Il�+mQD�U
#c�+j6�B�Z�F�$��3lU"��P�Kmm�5�TP���VZM�6��:e[[fjD՚�ii[M��l���n���L�6
�6�ՠ��+fi���66b�j�Ԫͧq��mT�k�ѩ��mekTm���E�Ӑ͋0$b�R��[2��m�H��5XRٌ�T�����j5�a�+Z�XͲ�F4�ک&Ƶ�1o����;kmV�f�kj4[hV��-��  ;��}�u�=����^��޽�ΪJ�����;o]�mjʍ�å��i���N�(��C��m���àV[��� �n�[AUg7�4r�.��]��m��Զ�_  -y!U�U5����U�j�`��P����� �����QE� xwۏE 4QE�� tQ@QF��͸������pѣ� :�PԳV��Wi2�#�4�� >� 
�^Ê�Er��(	��  u��N+T=�+�S���wtB�ι���ǜ�Z�wK�%�k5��h�)�Q�Xk|  �Ez�M6��8�CtsGvj�l��V�F��Pu\�Zh�T�4�2,)��@�.���hՁE��6��f��  (�MiE���:�T�lZ�B�Z�����h�s�ݻMQ�e�� ky�uٯ\�:�ݻ2�5V�'w�w���ݶ��
t��i�R�m�m��V�ڒ�m�W� ���kl4Ҕm�p��u���څ��=��קT��,��.���B]��h�*[{�tv�U�tm�MǍ�A�`��]���-���aK�����H�j����J�  ��֍�֟w��/N��
�ƕv�!�0 h�{����A���v�:P3& �ݮ�j6��u�޽�{(m��N U��9OoG	�kMh��V2�,�   -w��z�x�:bhU���$ztװ �7s=ۻ �V 5��m�� �];�WT)��ՍF�cW]�CF�WK��5b�-%M�ږ���  q��3�x��U\�=m���a�J��P*�U�u׻]��-gK�t ����Q� �g:���Һ�]\ u������a�P{�=�f�ljR�&�F����  ƕ(th3W� u���h�hs��کCF�^���^���m��t(�k��^n���E)���t���Msg[h4�jN^�:SZ6�| j����IR&  4"�ф���H�4`��zl�����20�~%*��@ ��{ԘiUS@22 I���b�)#l��O�����'��;��&��N��8�1�z��<�Z��{~������BH@�s_�BH@�a$ �BH@�脐�$��$�	"BH@�(BH@�p�����?������,��d�g/l@�����ՐŊ����M�:�z�ĒMб-͑�e�����-i�(�r�;�=�,`۬��4i�(�Zր���ӊ��4k-<û�$,�ueX1i�����u�̌m8��,Z
�xa���n���� P�j�Q�@e�/ n,J�ɥb�Qԕg̙{J�Թ����-��m�a�n�i� ܵ���b� �
� ^^�-������1ՃQ^e%�V�K�+q)|�6VV����{I5w[B�"g�\�"�;��0v@>�x�#N͓*W.�Ɍȳe�d
�#���8/l�>g��ɕu�2�F���5�U��6MjWbC�`���I:��2��+r+5%EF­��x#�*�%�Ӓa��m%�!ѕ��-<V�)��2�-[Z�7���+-ŔMRU�3�kMӫ���_#�Ez��3k�&�h�
sLOQ7O5F4맘����N]�5��!5���ZZ�(Gf��lщo[Y.���vU��SUh�q�(���6j���,�{�l��� ���e��Wj��h��y���Sf�h�v2SUe��!�=��K�u��Э �fC� �Ņ^�T��tZ�9�(M��wB�^��QCkoE�"\�8Ɲ�S��T.��Ӡ�[�3ha;ot,$%��M/v,E�5�M��z6���۠60Hb��!{S1Q�JX8[�6l=-v�����,c67'�qw�9ѯo����A���ȯv3g*���OqĨ�ؙ
�E����c�Ɔ��� ��#>�e-ݬ߅@Mͼ���O�h�Z�-vsH�84.�U݆�5�L"JR<&ȉ6���*V�jj����ǖ'Yx�*Hb��U�j<�0)��$�	�F�e�g^8	ł
S7 ��nk,���4��%�	�`�ٻ%�t7*�l�6HLd�-��V�k����]k��c:���S2ևD;�����l�s�)���S���[XX�2f���,��j�[�U��5i1��ǩe�ا�ҎN��g��h*hХ��zJ	�]sffK�p�Ra�&	����.�5��DYa?��tK�T(�e�H�+�`��I`=���m�*n�,R���CFP��e��[Bh%��@�Z+r:Zc���r��F鶠$A���.&1�����E��KN�!GM�bQosU���*��X�˭�R���_2	�/T�;�S���Vˍ|�ϲ�v�;Ol[�w���Q�lH+h�iH����y<�=�x@���5�yL�uz�4�ѥ�j�qh�ު+�e�h��kG��r��[��������������٧ҥ
ˠЬͨΊ+(�z[솧�5c0R���U�2!�@-el���v��2<w
9t�`�`W�hd��� [�ŕ�tZ2ie��ݣg4^Ӥ�z������`Fe��K�h����J��`z�d�㧹��Zʹ��źp;���.��{h-�Z�c4�dEv
e=I�X��b���L�Y����j�,M.P�f��e����� �f�"b��,�ZI����ð���w�����¥{�n�`�G���Ʉԏu+�xV|V���ŏR�EGd�7� �)�ۭ����nR�-H�3I�F���127�*�s3B�%ڹE�v�,fk��%�e,f��	��Q��ʵv�ٲ�mF���ѕ�س�F6�m6�*��wV���r�����i&�a4����lԮ �0j�ZUz����:���$]�b�#�@6Z�X���4�1 f�ߞ�2i���)�[e��X�`�G�'��_K�0+�M�mh�em�M�7m�JТ&�d(��8���i�H���I���̝�$�1���L��JJQmTj�X�d �;Z���Hi�WSb���yKPڻuf���Sj��P�m�?[n@'��$�c7r�A��ׂ3.��B�5w}y
Ŕ�4J�h���,,��%ȥ��ͽ�<0�l#�n�w���"
,x�5��?����(�9B#Wp�Iڹ�m[j�Eֱ��\.�WI�Z�7N��e�Ӄ�O+lҬ��Mח�k�%�0^K
W6� q�"��@��ώ�*w�F����
M�z�}3�3qgn7������9�Q
F�d�[�LmS�~��1e�@��[��㈂]�F�(��$�q�Elv��0 ��� �X�9.jR��栫uV�w���z�wt�咒�@$��BPVl��(T'�X��?��&�?i�,ֲ�V�Yx�.����%�w���N��6�z��Q��Ge � �f��x�[6c�;i*j�D�t�ɯ14�i�{i�;ê�mfc(�m��G���2a�Q�,�47v�^�-�����K+E��:Y�p�a���� ]���^#&ܪc~U)�C;�
Y�,ɏX�wn�\�ZKb��������n��R�P�����:�E�;5��4�o6��Qd0鈶<4T��%�45J[����*[�,d����z��ef8������t/�ܗ�#�M��[��r�����'&k$3cY�T�3�!��V)��ɭ�d ���b��r�d*��;j^t�=�E�����(DY��8f	Pk5ch�%n�7��Y3S���K0�7�������z��Ռ(�)��jU�� 2��%��s)`R<�JӣY� L�-h�����'��0�%cRBVM��q!�W��%����z$i��6��s�w�K�܀T	d��(��Kaь�����m3�$�@j�`4��Ye hL�f�L�&M���E��.�-j^�&s(X���
Zr	
�(���IC�Q��sM\˹��1�mj�Kˬ����%�j�`����,ZBx��iav)R��(\�m�9Y$�ڼũ��U �d̈́�S��W�p��w$���9A�횈"(m��+J�Vb�I���6Mf�Ql��en�",G�3jnmLYq�Q���V�����I�Z�e�m]h߳Z;�L$��֢�$��9��B7h�0ÆR�E�ݧ��y�A�[ܬ�^��U-\B�̖��ɨ�V�-4wm�ԋU&U��`��i�V�f�m���L�hfԼ�l���ee��)w�~)�:[6�W�yg%��n*,��lU�h%hDEjܭ�A �U���kՒ�|�h|�츮��!�ǁ�.�.q ��N+3,8�C���ڋZw��U�o/^�z�f*0\�[`��V��[�7r���!Ӽ�)�oD�F��r �;�KkbU��cFj�E��SQ`Ar�MVH��R��[{zj�۬͸�3�ě�-c�� Sʏ\�u�44��7��u�h�V��Sy�(]�,�@V�N8�ZeLf��MAU��2nL����U�h8�9���k�H��u*P�+�wnfQ�te��7#�8�0k7�����nkލ)0���	�� r=�`�.����Qn^[Fm�	���-ОlC3q ���Y��߉�`�*L
���YZi���y2D�U�/$�9�`߷lǂ�nRӹ࠙x�MҼy%!1�ff�@UJ6�:&�M�v����e	Z-�|!/R��0y���
���/D�"�'"� �L���BbF��+�4;�N��²�6�;'rM"�t�^��R%�g2�l%��P͌}/F�� Eu +	fSS��H0ՙx�nf������9�F�5PL1�����w�T K7wl=496�0RY��;~B�A,�m�œ&�h˲��E����0��|�Ҩ!�Z��1@H
��-�u��`����hKP�m�0�u�����t�.,�nV�6X�Y�/`;�&��"9��4�d!&'1�����<=���B]m�Mb��F���K��1�*3���`�$�2EقyOc� ��km'�7���j�G����t��6ݬ&Х��8�8Ӳ��3uڡG1��u�'�R�с��n�ft�����k/�=���i��n��ʴYߖP8f��B2�63/I�WY�C�H��,��M���Z�o���&�Ҿ3/+@�nU�N�S�k)�1,�mMG�mnf�á'DK0��Vd��h�ö���ѓs�ܐQ��`�IZ�wcb�ZiY�WyKh,�y�e<r�PM!�=�j� �+4@��Y�����3pٻM�v���A'N�;������"��ٿhEq8�G��6Y1�����7Kd�a+.�1B��0�Q�"	�E*̡G�`X҈x-KK!���0�WH̤Tq�e�����[l�v�[��f�YFf�)P�F��T�Q�x�l�1鬹zUF&dǶ�RŪ�X��yB��0���jy�m�9WV�2U]��.��Z��t�j&Q�SKX�Si�5Iy�L�3m��59�%��DҚ7����B�'���<�N�]�@�/#�-�U��1�u x\Z��b���B6-�g�o	�%荍T֬gU�0�0P��t��%�f�0Yv69��nd:���N��Ph�.�qh��V��K7+�\ά$sxt�h,1��?sA@TP�2�=��ot^����u�	����c��poɸXJ/y�ݎ�=OJ�h�F��nm^�OvT��
�C�
Z�pC��hӍ3PV��U��̨M5off�����	�Cut�Hmg͛x>[c`RK�S{��*�n�����-�vNJ�G��G��1�'
49�W[m#�թ��N�
`]ˬ
�ٔ�,�N!ͤ�nl��mZ�!O6
F 3@N=Cmj��n�B��t�u�e�%��U�%��e��hЩv`��ULP@�Cm�w{��a���M�΅j��v�n1�={+E]��n�g\�74�eE��S���}i�8�t��d��C#8�7CV�����YEĔQ��X�b����d�����Nt�r�T��k�$Uɠ&p!��i��.�iE�vx���vlM՛��VjT��������΄�ט�"0�qcb2E!b5�n�B,�ZEX��صG\Uk41[Q^��Y�Pg䁛2�u3^kN&R3�4�w]��v���6+N��.��A�:L�ou9e�THUr;D�������n�����Gn'{�nӶ��]G�/��Ԇe���Cm��N��#R�kk*���f�,Y`+�B4L݉��e[�P�P�!쵪V��ʧ�ʫv���%YA��@m�Enb� U
��r^�t�/r	��ٯ(�JVQ�5+4j-=z�f%{���P��	��L�gA�z�2lسTc3�&�F�23G0ͻ����*�j�,Bۧ%	�Ni��i%Ch=�e�w���JL�Ҷ��ֶ�6��ma�7CQ����2b&瞢CC
/{Y�(1@���5���l����^�hc��s.�@�M�#�ɹGƅ����t��i�4uD�[��jYzˣ��Ȝ��I�V��j���۰f�&��̓ ���L`E�0f96��^�8*���V3�aĔ�����bl�4���;bB�z`Uv�m]�lm�QI��@h��5z-��j*K4��oVL��3����δ
V�]&���i���5���� y����A!̼�	&X�n�]�������p��J�)Y���7�AXJ�:[d^Q��t�J�
h����b�f�Jf�B�ۦhSÐS�s�OuP��)�W\�K %��p�O=�VK�
Y��>�Y������7jU�{�T��{�Yn�H,ZS������S�%�r���8,�,�,�m*ח��ӊ���*̘���ֆ��F�ȅ��!4�� �=�
:T�V.���mZn���m��-c0���t�V�ę��Z��hT�4-ٵ�GN�s�$wg�Q �
k���L͸dp� SYw�%�.x] ��cMjX.��֦-��Ct�k#Scv��YZ���"��iV,���&Z�)4�5/Bx�qcwr�����߲��hڦ�\�QiV�*`9�Mb Sbc��z�ۏb�{��bM�Z�RV�Rq�x�J̶�Ц�ӢlͶ�#Iyc(��fVf�0ῶ�5m����XA�G��jmM�y-fiK+Pn`M���n��݌f�O`x[��we �a2��Tf�ngq������`�[�V���Kb���?h�s� �ѩA�����{��d�t ��݌s@v�A@�A�%��oNA�ym�wj�K5V���F5P��ٍݒ�C�+̢v�&Ĩ�.%I�oq�a[.���v�52����N�mmې�(U��ZwIm}�S9����[��ykU;�E���2�cX��#�RwJ���ѷ�jT�ÿM�N��q�yP�e:�ټz&�u��b��6,1�
�%�VFL�Z������l�M $V6�x���LC��eK�I]��VI;���gp���xh�ݻWXf��</7�#2�;SB���B̧r��Zg�Lժ�	���1����H���򔦅'���M�Q��D��D1b���̼���Qdr�U�+r�5��!��E���z�-��{�K���-:$���2���M�0�G/ ���vf�@�sIq�A�4���Bi�U<�M�u[ֵ���6l6��a��&l�̀��eb�k]�Yc �
*d���<�����h�2�o0�eZ���c�g�4�AF; ��[b��5Ic��+���{Rs��4Ø`TP�A.GaF
�sh!He�Db��ֹ��Z�dȷ���ܕ����$j͚�&�۪���V�mh�ր�N�)x%݇J�i�Hϱ5�s5a *�/�+�o����k��(�~����od�u�=�XC��������YP�x���U�Hصj<���N�ݵ!X�|=�]�lP\]��[�j�y�t:���]0yf_hnGMIW|vf�8-q�K�#wgS�|74����FX}�����"��w�m�����
�)iwީ\!�O��;���ɚ'���i�Ҵ#�A�3����(� �c���,�����n�G)P�ـ�ى���ڴ���մ2΢�������;���j��(gou���5�b��VT�f�Y�X�yrJ�QV���1��)P�E�n��W�u���/��{t- ��|������J۬׃N�%������7±�4�/��?-�a����|0�f�s�g�����h�z��Z(�;�\d*U�G��O �i�=�QO�_T���v�"�M�;[�1�*v�q3��9����YԶ�y�o�&�)ƈ�En��cd�ƙ����7��f�<�=��䦥����c��N�v��U�wAO��MѾ�yk���S2ȼ��\鼇S�Y�vw]�V��e.�l'� 9� �$��ԔhX�f�6�5�}Mg��xw[΀)ꡧ��8a�[ĂėC��t����+��[�e��j������=�4�"$m�>^Y���f��彔����i4^���^��FƦkzd����0W���k���A���oua�(d(i=�dް�ww�C:Ԧ�l��Á�����鉭`�z�{��U�n���T��"�p^�H�E��l���t�qn��A�ـ��h"�Q���'_oQ�ç7֘���5�+Q2��lu���_�y#�}�xU���z:��UPkc���bĔ��d9�wf����fJ;��,S���^�[�Ʒ������V�YJ���{-�*����?qFR��u�Q��O!ں�%F�:�j�%&�5�BS�+�6�wa啽A.����ob��*T�Y�ux3��a�1N{�S9�
�6��br<��uX�4*���U�aA�MfV�Px��A���9��k�xf�Rvf�s�9���f���/W�h/Cr��f��/�6�Q��`�ٍ839��Ϩ�b�9>�]���7FY=��w�dhW����11�ƃfv�	b؁�p�[���u�$�5u�GCwO(�o�2f�Ȇ./*8A����i�ޒ�2���X��o��ύ��`�F9�[^��0�;��Xt���ayc��0)��N����Bo\۩t{Z7��I��/o�Y"U\W�"lcYFĭ�g 1�]A�|z�ob�
s�[�M�,�4�Q��.x�t`��G+�|k���w��XTݭ@���ko�b�2�2��f��e��YP����M��&��&�7�A�J��Vյ��[~��q~|.W�E��e]���-�VCQ'Zx��zH�{w���.�K�J��nl��n�Aͭx��',iD��ݯu,��o��X�0��w{
�q�j�.:��Bm�����j0��n]�m����s_iD,�2?���f��;t�u%벬Fڸ�(i�a}Ɲ>� u��vS���^K)�=�TT̷["~´��ն%sZ���K���l��� u���)T�&�|U�04Zɸ_���|�����b�@5ZrY�g�C�6KuΣ6���Y:���������HΝt��>�YŲ�ʕr<��,�V��ֲ�T�5���j�(��w��׆���b�&����
�d���W�f�%R~��+<�S�������;�G U��ıҥ�g^D^�(l��6�9Fs�sO��s9�18�%��Vvfy����꿭p�3H,a)]IZ�5r��W"�"� B˾k\Ե_+��$��uھ�)�MytO+n懫�Ρ��S|V��Kj�2Yà8qV,;2�[��c��e�� k���"{�M
8Wm���WJ8��6j��Q"�q=��[�f>�f�ԡ���F8��]y��ӻ1U��s�V��'��7Xf�����#�.Jx��%3Ν$t�N��x�]��;b�5YӢ�!��$�Qo~^�F�w�U��~4���P2N�4.$��9�=��϶Na�;/=[饭q�ך�r҄���]�7.�T�2d�zPjۏZ�0�-^WwR�ԗS��r�����ct��l��7���7��:+*��[�`��d��U3]������(�[���p 3d�&X���3�N�cآ&��s�ZE����r��o�)7��n/fcM7��5O����zB5�b�iT.����]�7���Q��_)i+�� �r�6�x=���C�0�X����Ƀ��k�5�|-v**�ʘ�e�b���+2��Ch�=��NΞ���dG9OoK�S�����K���}��_yyQw�Wh�nf�a��rW\BS�G/�]��(��p��C�Q�k��r�gU��B!�1Tp�KW�G��2y_d�VE�,�1��������ۖoU�՞�H�.}��]��O2��S�t��q�]�����wh��$�V���9�N��"=���KOGvdңW��}o��D��ިru��-�<׫UgL��un|h`o�J�j<0�ܬO�w*�F�9ݮ����8f�e�n�[CQ�����dHg�/<�����_��3#�`����5m7K�م��*(����s9����zXama/^�����-�F6��P�$�IZ�n���ŗq>xӖR��{{�%Q��9��p�sDO�ܠ�7�i#���]y��>�
�KA4Y�L=�2nm�v?=w!�tf���'a{��f�T>,+���_v�Y��xZ!�{�a:)��l�3�r����7"�e.r��5�ċn��T����''N�J8液��6�u�#}Hů����5c�.�';X���M�;tj�Ҝ������I���gi` hIn������bkoM"��C ��x�p�g����� S0�l����J��M+gu���V�H��&�](1����2�/l|����+��P��w77�T�j��S�rB-h>:�pѸ�u`^C0S���SH�t�)�k�6��13!�t����JD�O�j�943�d��vV����wa�� n_m	S-��@�ZQ�U�P�:��R�8s�Kq+��f	�a�9n��=�6+ń{���iݨ��+���BE�}�h�h��p`���k�8wv��}jZy�JZKE
ӛ_�PE��9��m��B<c�h���U����xM�kF`�ޝ��皇�-�S��.9�P�u�u?'rta��G��^��У�o�2yh��ӷI9�|�oY�{�9��.`�:g	a��m�cjy3ޜ�l�iw3�͍��!�)�y��� Р��.��F4�I5�^ح��lo�۽���O1g�m�B���B{ƈ�/�{{O9ۙ��zs ˒�c����%=������B6��qr�L�J�#�]��+��5wt�8(	T���A�3,E���^Ӽ�b�wU�@RˆN�:.!������3�.9��4��JLմ�e�C�VuI�G��^��!��ky�I��2�i:�=WY��3��է0NxN��˹[
еF���.�q�j��`�aj�� �[=mQ�>5�\h���0���t�]l��Ea�Dg�<]J�;�,t,�w{�+�Չ[P"q �<�*��T���u\�oV+(�<��wc��ޕ�uxnb��/p�\弶�D4:�n:��n���ҧ�Һ���bW(7��W��������}��Ul=�W	B�8���v�au���wj�ƶر
�&^��<G��)Ѭ5�'�b.�Ё�$�a���v���u���tN�s��\+�<���]Z�	��v����t�@؛�u}\g]+V�i�P����t�����fs�5e��~��7pJ�]me�v�S�ܸ��ј�sk$���S�#P��;�ۅ��b�J��<���""�[F�,Q4�:M�����׺�����vt@�]����֐
���1V:}g`Y��>'����vҭ��_Òs�f*����[3�<�D{n��:)qHՕi���-��c�ք�o/m>�W�#��(�V^JZ���V�Fv��q/L� �%>�����P��5�n7CC/[L�ر�*�'j��+��`�)�Q��٭8�t�-����/wR쒛7Ǳ�l]K����_m��y.��"L,��1�B3;0��ǝ���.��,��ԡ{5-dp.,����߉�2s�:f%��qy���{�B^7�n,�ʩ��li1�b�����ZY�7ࣗ�s3�[4^��J�e*'��ˎ�d#k��|�����l�]k<0ɵّ�o�=S���*V��lC���[sM�9���Y��0=�`bnj�uH���[�h�I�� ���)\�d6�ޣ�{�r ���|7��a۔47�����iR�e 6�5we�
�%hr!=�V	��;*�XE`�s!�у�m<��X�����˓YR���r8
��c��p�6B�sF�X@��X�� oz��0\E&n-���km~%���������k��ϕ�Y\G��:�.�ͨ�Z���vnRʋ.Td�%�56���]�kS�:v���d�[9�,t�`B�/��s�γ�.����N���7�;��9�����d����c���$В3N���[l��aT}�[n�V�V�y\2"�i2,�͉S=�� םu��<2��(9K�Dr�o4��T��W�:��>ůP|�G�<�b���	�d�-#>�S͎`m]��Bp"�m@wΌ�ݘ��u,�'z��l�
9����i��Y����55#6�[eS²�X�#��w���{�5�e�D�F�F��M�2�IT)�6Xm��|��W���G�ڹV�\Lyݸu�竃;lKr#��pt�$CwO�4	%]t���B�zT��bP��dˈ�>�{֞o&%��k�߽v��s�.�ɪNG��-�u�{7i��{=V���k,�Q#�;opnvE�0�f^�긲e8�;F�{�)�/A�16�r&[2�ě�U�ϖBN������+5Js��:)�YV��tћq`���Q�I�[s{ ��}�*�x�i :�ZFo�ы�oMu�˙z��:A��w;�)5����Dv�N7{+dؚ��֋�V�`�>�[6�l��Ŏȡ]�j̃��!>�+0�+�L�'��*�V
�\���P�Q�ͽz��Q��q�	✰���^N���L��%(���kR�Ӣ�VZj���k��iJU�b�B�TSna�yظwJ�-ᦣX�Ɯd�E��˿D���r_N�0bt�3Â�����3�&���
1���Q��k�X��|�g�M⦬ܽ�������U���=h��R��h|�y�%�n-�Q�s�PC,��	v����\��F��!Äߚ��%X��ޖ�Xkwh��������sfn���n��A�%׌��!^�Y���u.�f2�%�ݏ]���î��J��K�,�(��dd�Yz�8x�G��z	�q�i�n[I������J��'�n��H��>��h��6��,cu4���y]�����p�M6�v�0Wu1�qm���]+�0��+=�^m�TU��{�_)�1a��xܽ��WϦS�b8����y��<z�s*<�؏��g�s���z-wR���9��jVh�A�(u+�.��Ԃ���#Y,��}�{��Ź|'W�4�wr,�¥�։�S؇]�tNc.×Z�a�+x<������R{'���L��6�`kb׽T�H�S�^~�,��b;�y�wϜL���6�8���S\�}�*}�[-[�O{і��]�כ�y�P쀥�n#V>w{�KM���$�m(���,t�6���hp}ɜ�����WV�V��t�zQ�SV���$!��vw*4�r����e�J�*�[���-���j�qt8:u^�7V曅���[ ���|����h>�Uz��q�U�tK9x���	�|��X5�[k��k ��q�,⢟Vr�NJ��������x#�>�8ɉv!�Z���Z;�ZT��G�*4V�U���X���/�4�O�V��yS`;�2�a�L�����9�#�|��ԬԻ �ǥ���Qo�[Մ�-�m�MUh3JuK)c��z�O�"�R��3��օ�)U�2w5v[�X�m<|C�/d��x�|f�"��j�Y.X�	�ݹ*�tM��z^��>C݃;Yu��lܙ�H_mt�:�VD���X⫮����r�c"������N���3l�����-��f�}�lUi���ָ��8j�מ���B���5�D��X��v).l�62�s �hћ4�xW4�4��-�Qg՚���^�,�d��}|����q�)K=��1#tr��jv7��=^�ՠ����@)b�1��t�/H��O��˼��	� Ц��-ڎ�«lO�t�"���+ܮƐK�t�]����La�'���z����M0�9�g����6��D�k�I7���b6��wɪ^��0�d�����3��Sk6�jŢx]p�T^#��Fi>���B;=t!�M��5'A�L7�:Ek{��YڧW�;]��I=�v�j���Lr[�n��ˋ��J�����Z�,{W�V�|��E�b��3�g�b��&��8{oyN�ԙڛ{��I�j��k!R�w-4��chȦ�AA����淚�ԑ��fP���.�^v�:UC�e���7<�m���ꨢ:�b���AـQ��S��36n�n���4����#�N��Z����8����Ԭb�R�`=��h^�u����m������В		䄐�$�7��|�s�T[B��_��A.v�Eګ2�ot�{� �o>a����)E${>�^�Vw\]���f��L�Wض��>��2�����cb��n�0}��^,�v*�R*U�0v:��e�S�
]3��U��qU��l���[��[Z�f�]+��إ��Jڼ�%�B����v�*s�r#�oZ5��ó\B%�u̦xl}K*��i�m�k�nx!�e�&ܞ�0{S1��&Zљ�ֈ���&i�V�P�;���`{I�c�����ֱ�7;�E��C�̡ӻ�x��l���L����l�\���;Y��Vm,&oe�t�u7P�y�������3�T$����8U��ŚR��q�]�9|�9 ���Z�e���E�2�B��v=t+hX����؜G����D�rD�Q*�B�;OFRl���U�(\W�^���q&]�W`�I��JyY|��4��^L�]��n������+�x�I��vhj	�}��NhXg����h�r)�B!T��BɯB�г|e���s]��T���u�{��pj�m�G�k��]��P7�Q��
N,ȩ�F�X��]�s$�F@��nku���_Ė>B�ٗs�t�Mtܬ�=�%ױ�#'�ؽ�I׊���Bq[��眯�y9�=EE,���+��SHGul�nޞ[Y �B�'��zeI�	v�;e__�f2��0����-I�8e���d�0e73��h�ZKg9Wޙ�/�V"�x�/N@b`�z��-�L���%T�Ռ��^�w�!��'�S��L���`>���֏���lf��=ف/A��,wG���n6B�{VN��:��\����������|�[�tNH��͌�a:���D���C�=c���m��1+9	TwQC,-
����)s���w���رg�=Ѣ�W�ݻ����"t&N[��v�ИJ;]���zs]p��9|�[e��]]>X��q	�x���ZXB�*��E�ƿO$�̊��؆��)�C��ٱ^��`�VS�Ǐ:�J�f�VgT"���@��	��G�]�ed�e6�g=�/a�*R���8����;;إ`̍�)ȣ�+���h�"r�^Ǵ�4$��PN�$��>��nG	�e�p�+^���X�^\�^(i��P4�#Shvd�ݤ����*��Z31PFy�v��;�E'X.�A�O	��GD�r7¸���1"�k��}L(��4��r	��<�dS�3�z�+�%��#��.j�l�:e+o�Mժ�i�!1�����W��۝BqWZ�P�^��3,&m5Ӹ9I���>Rtۇ��oE`�V|����3b��H<ֺtDl�]0���X�r������z۽��eH�wf��i<�g�k-4���/5WVr�̠ؕ�Ѡ�Ԯ;��U��՜�'�A*�H	�5i�irl~�X�'���LԖ� (V���\�\j^��-8��Q�72kEP!_-�7�J����*P��ڣP�Ǿ��w]ZD;?f��7�<}�͍�s��n{'y��_�d��;:B��p�������i�e�nE�BwL���[�ŭS��i���q{���s�j��Vv3�T���!�[�e^����.m�R
w��������]ncQ�շz�,����)��Z��4���j��k[�T	VQ���n��Ԕ�	������3z%e<��
�n�����YH#&����Z�{CV6���ݰ�jvlϮ��7YΣ�o��m�]S;�3{���f�.5�A0�X�v�n�)GS���>�3o�U��θws����k,�=�H汏�n���}ē�������n���s�u��7v�u���Ojb�e��D��Ŕ}�8o!�q�c�	౶9|��\7�Y4��F��#x�� Y�=�'b+GV=�-�W
J�ky�U�^�L�>[���K�%ܡΰ��S�#�ޔ��(�|g:J�9(��.w��2��M��B�о 
���͵j�u�T��c�x��1%'-��:s����{}ۨg7�ՀA��j�U�2�����태]e,���A�@���8* ۬�2�YtnˍpW�7Ҭ�J|�'���N�� -v�.���v*2��-*����B��E�o;0�i�e�)o#BX�T�4���3�5�Ϙ�W#w�h��7��v�q��W�����7�P���U��շ�X�Q��[�z��ĜMH*m&)�/�y�ڗV�Ʌ8���f;���Kcy��Y��0_�8nӥwZ&�.7YB,�	�;k&��F���Tn�8s"�b9Xkj�ZT�\�#�iT"۱P�ke��B�_K{݊���e,�wNˈS�p�"@
�q�N:���S9?��s5c����g��q���a�]��<����e��a-I�����s�-���V�A�2��3��(��6);P@ž�(l=Zx���L�v*���'�k��nݽ7�lO��`�d���)��_f��Z�nM��V^�|W^�y�y��}�Qy2�$t*	(+lU�݅�{q��{v
Sp�;��pA���p�Y�Ŷ�cA=;���e�髛
�=����0n&�������W]ɱ��g2��.W�u��:���A�>/+8Jn.n�،��jR�t�:�',�<3�]+�J�(��f�<������0Y5���M�d)��X�V�\v(#�pw��'v�M#�}���d+��RY݂�b�h ��3��h�.�p|��SE�p���J�I76��3�V�����[t��p���úqT!Sv(pKh[W��Z���f88�ߺ�S�j�%��h���$�J��9.�s[*�Tp{�X�6�,���=�؛�Y�ZG�j�&wc�69���.�S����p�g�賍���0��{C�E���"�c �0gD{���3WD�ғ������ ��_����xqΞ�;���Ӵۡ�Vv�j��j
R�8~�|v�@l�v����_�gv��'tt) ��"& *�ҹ�r��𬼺�=���Z(�f*|�����#�5��n���t���!�Cb�)it�Z۝����tu�.��Ltni��~J��v������<)�zw��ֹ��	غ)\�<VZ�m�D%�34c6��WW!�Eec������͂����j����|ܣ3>�hWb��� r�p�1�YA�pqޅv;!QJpQ{����:�á\&���&g*h����`HJ�M���0��I�0��m%�����Ҡ�u��[����L��Ե\㕗IgM�_�J� �<�6�+U}��shm\M�7�ɷ��n졵<���,˝���sp�]{�����r<nK���T��ȏc�̎�=����ӊuKR,�]�Pq�kE/D-�Κ��72���y���kB��F��\Y��ǵ;`:��9 �Ys���P�ةA�N�H3r�k�s�.�����6�N�O�cy>�z�]*�)�ԗiatLY�ɀ��6�&j�k�o�XW��Mhn���T�oF��hw�C�_v��J�����{-�v��zQeKU�D;E,��f�Pcr��9RTU[��V$8aFt�Q�/YgI�::��k���Q�c�6���:wp3Q��iՍ�v�k��x�����=ana�`d�],�c)u=��	+����<���019������MG���C�15Vr�+&��,�%jԅo���7�^����3c�2��%��Ƌ�����e�!�Z��������&�k��v��uO�ȳ�f���y�A���T$u�*�c�\��(@�+��>#jIN-�U��t���a9Q�9�[�XQ�S;.9d���3�B'n��罜������p����c#�\����F��N�}�Y+T]w\;�2�q�d�5��t-�A,%4���E�� /!��>�n���n'�V�E%�b�̀�}�X�cf�+ʏ��ی�ܠ5��M��O�a$0b�Mp�W�&-���M[�L��n�B�!�<$ˏR������q��H+>�dgn��F⮒��xkp>�L@ {x���4#d�W���#>Yre5��{��V���DWr�`ZFЈ��1b��f
���IU��+x���%�`���)�$�2�9�󂑘���)��2�Q��lr���+�ӍӬ�	h��۝����vN�,���s1a�=m�5U���z�ֳ�̽�n�)���<|F�Օ�ξ0���x���9Rz��DnA�E<����W�a���R��}P��\�yz]��j��]D�f�aiL�t����LAZi��z��a(��O/,�0+�s�hE��W!
��&\s��zu�C9��d7Yc�Bb�o>»T�.g�i�"��`.�~�xE�²� ��Z�g�{<f��@[A���[�L޷�w�peh
ݼ��V��qWp�)�q��)��X�_���-ᾷ��3\zfJ�_�;�r�*�k\�Lږo�8g���;c��:7�F�L�/��W8������/�U�9U�	Dkヨj�o���z�t7%���YoH��2�omQ����i��mm`�M�h�imc��*��l���@�y�u+�K7x�&��wd'pN��;�'�ք�,Î�:D�M�Gn�/7 ����έ���c9�",]-����=�{2b��s9���J�W�^(vBA�לO*��
�����b��쫙L�Ɍn�hA�7I�o9�{<�3�/�w���]y�H�)`�|'j��џchoY���v�obc�3��C���c��V���G�{fN��A"3v]6	�s�VD8Kt��=J$�t�`�w8\L�}P����yu�r�<�5��*��L[Z
|˧}�]��νV18���r�X��y�vVcqg��fgA�8�Jлm]��f��'7\1��v�,����8��c"�����̀U�.H�&(%v�C�ecT٘j�,�n���a<��2H�=h�+^ ��Lʁ(4��&�{0U��Ⴗ���G�(x8o"8�yd������BŪ魨jmc��p]%�Ü%�L�1�I^f�uz�oz�#vP=J���,����UsvfZ��]��J�NF^��iX�o�AQ��eZS�_-�<-�+�;���ҳװ1o��t
|��(Vb�z�����*� hB �����5��@�GQ/9Z=���J���7�+�<���%ʜ
r���q�G	ڂj�+ �����Uu��]�r�ݶC;��}�gvK7�;|tFcK��k(gM"�Dև�Gmt}�6�l�.t=��;�w����Z�Tg}r���;+xV���Y�����uM�II��4�yx��Qf�$qW�p���y����g9d5���_q��	�4����9
�W]@�n����5�u���]
:zq��&�ve���ܞ�-X0y0q���5{:V���4�A�{솊C]�����Z��&u��:��ݢ��+o���K/Pt{Cy�pm��:̼W����F�����1p�{\�@c}�e����W�6��{>�g���mn&yl�v�$H��k���ϥb�v��Δ��� �lf-Z�c(�S�љ�uh߱��r|49DXY���N�q[޻�k��r"E.�:�΁�C��ہVf�{����#��
�����|�LY��a��ˡ��|v0Wi��p�Q��Y͠x{��������ݔ�;�d$+e��LɜZ�*�q8(u}�s9J����J�惢�bL{;(P�BH�rͤ��������HK/���wu�|3ޖ�"oj<���f�-굋.���D�%���Y��	զ��T�EhG{����L���!���n����9�s�uu��*f�㿈�P��	�0�GO&aΦ_U���y�qĠ����q�01�^^��~�l��$'����',��G4!���^�uט5~�8�̙3�x�1�6+iT�۰��`�Jr��9�6��r
�Y�.�' y�޺��7�	^���[OE<=|"��sM����^��O"T̮2P��۠�u� ����AGj�[s��3�F�] ��]��֑U�g��a��ik�P�5�eK�\Y��0gw�D,R����(���\��}��s�B�@ْ��")�E�h��È�3��A]����r�4��i^�x er�3p穌�v�g3K3'��vr������NN�(��Cx�>�SR��.�Tnb�������\���[�]�\t�.]e��,�6���p�X�*͊�7in^�(�X�zh������4,P�e�������\d�H�q���#�؇%���%C�e�4�!�6��Z�V�iY�ƨ9���Ms��ׯ�op,´�<�] 3M�j8Q�r��`�Y�%�g�s�wWm��0�˚4�֬Ю�,�ۍ���y�q�0�s�jR���utS�T�o	w>�sZ���j�x���R�dWlV��#`Im�Q��wIlf19oh��:[V�o9ݫQ!f�AM;ٸ�����_>��6�q�	��ؗ��}���D<9���R�%�ʴo���x-��Ԩ_��6G2-Q��`���W�(}����b��hu^��K��/o(�K����`̤Z!X�I۰����0�O��������Y@9���W�7���uk �����B��G1v�n�g��:L��9N�r��������b��$G����Q;Z�/���_�p�f��/���g5'\:6N�G��v�L��n�	V���VeЫ37�|�Zu@�O:�Hq�D�r�\���}���W�}�|�<(�<='��)�M���uι��M�B1αHMJ�gu{0l�8fVr�|���)�K�{;6�+ˋ�k
��.�f,�n�8�u{�L��0X�޽�R�ȏ
v�N��:uj�'����v�Q/���˃�޲�Eb(U�9oN�y]Lέ͠o�u�:�C���7T0.#x��et�'\�N�;�<_*�2�o6���j��Ȓ�79*��Ny�]Υ�LK\��Z%��h ��K�ڒ���e�6���k�'P���v�{Ai4�|�W6�b��� ���'%c�;Lz�N�3���T��qw�ݧ�DJ6.�v�FZ8#�o�Ś��5��R�!�x������m1��Ɏ���[�3��]a���s.�6_��A㹴Et�L����l��=���Dз<{�իC�����I�}�p�n�q�xX	��.��H��;���
4u��,�Y#��k*[˅l�'c�+���ѫ�]�s�j</+u��¹H(m��.��4汫f�P�9����U�'�;�{�U\~/��EZ�]���\����yh�B��wT\�
�D�t��eYO,��ݭ�R̊��2O�N��l���w�k0o�$���ё�3��3���N����7h���Aʛ]H�e<�[ZK�O�ˁ�n�=�s}}��rh���gR���b�R�+��$�fl����ռ�8����@X�
�ATPDP-��AdU�m����dF�U���a�����&*()b��R�ʑ`[d�X
�EEE�)hŅh�JVE�,������FV��k
�,
ȡ��DI��*ʅd���������AIR(Q-VVCAj
%`���dE�ی��� ��� �,�-��LaXe�1��,Ҥ̠b��
�e�J�¤����i�
�`VXT&2˙	R�1��T@R�Ć.Z�\�K!��ĕ�%H)��Ԭ�HTBJ��rҳ%2��V.e"2)�+	�m
��>�ꤍ_��I.�ZV'k^r�^�i���b"{�[k���.��b���)\��N1!��fv!�e=�k�yW:ɯ/��R\�K=���+�+��\{��}k��8|�V�F��D ����T�ݧQgI�o$�v��.7��&�>��_�3ܳ�yp�|e�<a��0���BXyi!M��y����ŷl]�+�ۄ��\�֬��A��wOu�3%a����\��q����8�8��)Q���i3�ۭ�Ā�>�w��0kמ�5�[�+��H��#Q�>R�-���!:ˮ�k�"�9h��ð��\/�\%�9���j�,jO��_C"}�ݙ�k�T��+A��x��.7��|��}U�� U�xl1�.�OeMy�]�Xx)!I�O��u��Ք��><�\��3�x��k��%��X��rp{�܆n�/o��ng�����;/�g�]���e�gr����Qxy4�,��[�g��Fi�f�R;�o�,lV�4����ܤKn���f�KP�6^�\gVX�ރuY��/N���=���g+T�-�:�����K��*�if[������j��zy^�x���>���ఒ���̹�^���G^V�<��;%-��*Y5̧h�X�E:H��S��1��m��F��>�!=\�զI��ξ�/gəhBI:����m?f��u��_�8#Լ<e���ӊ���$=�k�v)\���oy�җ��Spg�dXå%���q�bµ�D����Qg�������K=|�U�7����/�4#�U�='@�?�#�P�����M��V:��PL��mj��h��_k�n���g��3�cW4��$�CmݭWGQL�M�ku�c�z���w�jt�>��B	^���"��8���|׭}�kD�N�%�]L�f]�ܔ�G��SV}^[ ���}cZ����{�8��������S�)Bt��P��z��)�֌��� ��7N��_z�]�Z���trv�ȡ�G%C�|2)����)�pje$O�6I{iqH���<7�nE���#��+"�˷������e��2�1;\�8����]�^��dv$Y��ɑ����`ޘ).y2���U�~�ݬ���4kþu�.�x�L���u�W���n|3�C0Z�����v��L�3��/}T��(Tr�P��Xg�v��+���K3��x/|9E'�ѥ���o�V�E��0�K�l8�2R����x�[@��c�{|����;��P���g���4�6e��	u�vO7��^��M�-l�A�)�x���nu�.�����8wUf-�'������fVo�0%Йg�}G�-��m���Nr:+ZݮNZ�O,�ؖ7{���R��\���q����ɭnE���^��[{A���"����3�t��1�u;�M���\}�ь���5�</��`u�{#��cu{�gxT��}f�YR����NhX��&4���W�U�E��v��C�����N�/}�ð�w՛ф�1]t/ɩc{ڵp��8�X�u����LzRXϢ^K�pX��A�c�I��P�]�X�A�{�͸.��ׯ��[�����i��J=���$�zS�@�^ i��a���	�ު��Q�*l��:����ٗ�ys)G���Ta)�qJvX�H�kj�y��o_{�,��X^�nrE�Bb�J&�����Ѝa�Wj�&Qs�&���x��1]���-�p
T�e�x��sW���G�'L�y6�+>���X)M�xK=��k_W�c�}���%9vP����=i�۹���5��*Ƒ`9�g�%�.�Q��~������gw���l4M}ґ&�#���
+�7���x������K�A����UQT��;M��=�ڦ��2M��l�q�m�ɶ�����@���^�9�hTѷ|�eG��7wR:��t+�m��1������r�<;}�Ի3�,������zql!^�^�̹8�Ȼs��(3�\z�pDu����p��mֻ�B;���|�ݩ�s��,(e���I�uL��d2��^����Y�]��C�꽳���z�Z��?v4����t���"J���f/-�,|��������P��ZiN�ǚ��{�o�ܞ���lr�ڞN��z�L�#����sv{�H��c|�%U���q���^�S;�Zf,},�hND���Z|-�D��L�B�}zV��k7~��^׼��C|�!om&j�+�V��^���ү���=��[�{<�	��"�M����v+���*'|s#Y�\W��5�_k�#Ծ״���^3��'�o�n��͗�ڔq�\����v��I`���lY�l��	�ߨs�½Nc�eo,rK�X6���q��q��&���^^�\��S���(l��+�R倿���������+V��^�0M�a'6陎��~j[��"�α3��Q}�&��Qf���29O�כ˱�]��ꊲ��Ď �ԉg��,:��x5]��>59J�^)Ftѵ�eS�nHg��V���"�2��+�	��<�C�j_N���%_�x��Y��cyS8��֗�D�m�l�a�oy�d���6�Cgo�.6��@P�Gc��:]b���f.{
1p�,T��cÓ�nR��j�':;@pݵȣr.l���K��P�J[t�o`��
8Yik�P���0��5�L�z��3M��S����d�X���ѪF��ʀ��>	�_�rf����fo��<M?���!��#��Wd!Z�.�7�_<���GL�h��Dl�!���]h<�M^�Z{���]*�{6�fK���ҩ7�g�]k£�W�k/�pu��t�WT�i���+�q_��׊�[}�j���ԮK�2/
�zYq_�	ꘅ�)j�
��@��ixS�[��7�F��[���F��o�=��m3ܱ�\/�]��
kAȡ��B;��tã�5YՖ��mu�J
u��}w�_ö��3�輬�u�3 ���U�N8)�$3�oW��{=��:$�ei`���)�X���r!����鑘7�
OnEg���)eӄ�T�_�7U���[�����Ɗ.��]�O<���Xt�޲��^�vqC���OM��jm筴!̸�yӷF
���8Y�����p���L��3֘5H�ԙ>�q��T�
�g��(�Fy�ߨ)��r�rjZޥW��jv���N�x�:�Ipmğ��t3[��}��ԊɜIV��6@�/g��pp��3b���u��etv�:h�3:���p{ˊf��۾��W�!^as���Ҽ���M��Ά�A6zPk�^��u~��u�����y���f���G���O	��ߓ�r��$���}���z���ż=^L�#���?#����dn�C���e����}cq���.������r�/��1Au{}�e�=�ĝ�1��>��a��{������)א������~H�_$v�-Kł+D�x�Z���-��P��RǵVL�Z��G]��$�s�;�Ngիe�]#��i�fUm��G��b�<�K^Ҋ,��at������k9F�r������>�Ļ�O��V���4E��#�Y\dYU\f˲*��{ˮl�*L�פK$��j�t�h[��k�����E�f����j���.-3���ʷW��~��k��Wa�a�ŵ��8���2_5�^#�SD��7%\�A�;�ih��ײ"�OAB���ҘۄkR�X{�9�s�#�:|�I�_�2á]���g��5�Z�!շ$�"S4ҿ�N]��C���\K��E�b9a�J����kOE�:���|o&X���M�=���rV�jߥׯ���I���$pR̫�b�<n�ݳ���)j2�3L���i`-�}9�B&y�Y��ŷ�+��Mְ��U���:���L�)l�=�o%2򞻎�� �u��`幔�nU����2I�����ë3ov�m6I��\Uґu��g}��\�Z̎`Fĕ�2�9��*�]�M��>����k�(�:2T;beه>~4�Gb#����;ku��խ�ۻ�>���wW�^[�����m�0s�(���|w�2�Լ�u3U��g�¯�}r���I';YO^�x��&}��(Ab����+�j^�+�p�K�%^	����U.���MK��-^oC$�����yC�gm�G�q񏥓Z��wu�9�����/k���삡��iS�"��;�CJ����s���ƌfE��Ն53��>���+��X཮o�޾'_Y���s�ՙ���fT���2/8]�s�蠭�bu-e����$hR�@����#Խ��N��b�����O��}��_���M0w�I������j�M�����]ӫ��j���:v�v��˰��F`�4�/S'g��bdG(Y ��Y�S����g��`�2 �'N ��g��a�l����y���}�2���𗵆h���2, ��v��N�{`��h訕j	\n��@؋Wu#����[��k�9���+����e��௰�{�u�V�x�z�eZ���Z=яf�̣���$��IN�58ˣ��Ի	�\�X{��;�<{}�շ��8�V�r��O^�;���	�䞛'�u��Z�-oD'���ɰq����]oZ����3�EW7�K���s3�^u1��a�pt����3�c�s��[�Ny���������=+��=~��PvҴ"���w9�n%ιs�O>�W�������8��3�:3�}I_��^ns��>���/nE�à�<h.�V)���k��v�"�wYy���Co�\�{d���e=�!����C���^'��"����VY�ϳ�|�wcv_7#ό�-��,9��?�`�V�*_�tV���[�=�s˳�g��ٶ�>ٛ�{�q���o�kF�ܿ9�����x���M���8���OǱ����}=A�r�\U��<5��70S��G�E�<3��ׯ���z�-��O?�Η����S��olt1_�nfK�5�����;�{�Jg�����9s�I��A����uF�b����)�;���#���[�R]�3��=3l2�x������X�K�R��IZ�v�wZQ�1��4�y�$*�4�k���k�-���:k�{����]/�����/Ww��(�ޡ�T���A-ڡ��{��{�a�뫇�I�<�F;$��Op@+yؕ/0	���/y�U�-������VJ������Ks}�c�z����Ot�>�q�O�����Vt4f�N���37v
�*��V����н�]���d<G�9��g�L�OD��OF�)�9�����{mJ��-�`>�l�zd�}�%�\����B�[��t�����ĿTcj���3��������>��e�&�x�K�l�;��p篻�A{ݙ {(�/�p�u��<���������|���_��ʗ%�	�N�h�|a<��t^����Ա:�ڗ�'�q��糠�x�X��o��/o�R�tCg�{�er}UG�����kd�ꂹ�����vWO\��'��&wB�n�����Q��W� �����j�K�/L�z��:���	��4��~T�6�wP��V�-��</�5{h;Ď^�{Y5�z�Z]�w8���1��.�f[C[&���=Yݞ�c��𛷑�.��ۘe�[72+=��Fi:|���l�}=�w;�>�W3�wR���f��ý�gI���߻��N����yI뻝���ͭup[]��#��o��l���V1�~��w?"^H1�͓��D�7����k����Kr�9w��ۯ�]��]6�	o��z/7����])�ys�<���[Ά_���澩�p�8�Y����͡ws�1<�|����̜A��n��Gg��Z�m%~������
<(���uS��U���������:K���g$���:�;��G*���f#����e\Qݮ�3�c~�s�>�réy���f����v'T6��R�́Y��5������/��ߌ���,^��P`x�
ʎo���Ӝ8y�Vv�>1�'��u���a��u���>�7�yv<[��(���zr���o�Y���|v;-v6��]R>�U�Vr>l��^H�*o%^�K�X<�wmQ�RƼ�X��K�W3�r�d� ���5R���J��7���9F��'��e�˂G�a���su+���@=g-�I�{���k��s�Q}ط­��EE�:�=M\���ڔbuk.)�l�ܒ=�Y���6��{(�a=ʗ�':�&ݥ0���u�䛬�㴰eg�r\��^�hB�������¯zĴ'���U�i��9�vM��������gNW|�2I��X��Ɣ5�hR\!��O���e��ǽ��Ejhw�x�B�E��(����"MI�N�X{���h��nNc�*�͸�9s�צ�Ç��Ѵ��W���5B��˅P��H���)���b�FK�x��<�v�!�7S�M�ML�>��z��ӵ�(�+�o�
�E�$�؂���wUc��J�dzfV �b���E���B��k��*��Q���啸��i7a�I�G:&��	�M���}�preL�E�R��>��x���%�S<:m=T���=��m[��91���(|-��j.R+��sXV5W3&�i��mAl���ܘ�)G�o���u�{=Z�<
G�Ww�r��+���2�����AD1��M4

�RO,�ŴM"�4x�ꚁ�������
��;^N�W��1ӏ*�=��0iF7t_�k[��^n�}��]W�F)��maX�H����ٖ\3����޹$�jQ=]�"���Gd"�#�.MoN}Nt��G;�:(Ƿ���s7"1c��V\��K;ʷ��8��u��9HL���S���@�w��st�5YC�EM�&g����Z��5��4m����1Wca��!�%�k�5� nZ��ň�\��˯:c�;�=�	u�Su�^i˾��ϼ���x%h\��]�cc[;���9�m��ӷx���j\IF�ge�s��u�9����_qA���'m�i����&s��x9�c;:J������A	Y}���z�;�R�[���Z�zݩ�ݸ.�8jUM۷�LAL�v}}���3��u��qQ6�ꓢ�8k��`=��|��U�!_nR�s�F��r2�NR�4vp��R�d6�o�
��n�XU.�������"�T�sr����*�\�q��s���A��J$�(��OP۽��&�!�^����"��HW��C%�)S���N����Ĩ�v8���mU���u��'q��j��-���zL&�2=��[ů\�M�7r5��iYn�k;K��ty�kU�Ò�P�Q6n�E��ieMͷ&Z^�d��{��i��{�։���nH kyT#�e�L�
Jv��ՃB,º`�p�y��d�L2�7�v`��wx��a�����zk#�+��d�Bͼ�}a���5�!�;�s��_<ߏ��^{�@��B��Y
ł�bV X9L�%[A
J�FH�*,
�*�J���A��e@�Y-����,*�m%ADk-�RE%B�*J��6�-T���+���ʊJ���aR(E���ʰ�a��RV��IY(�h�f2L�����YT30b����J�ɉ1!��@Q�+%Deq#�d(�Y*J�jV�2֢�	r�cP[i"�-�Z�R*e�P�
 �e@U"�`�P��E�!Z�R([J��,�0���h��KH)*��`���-VAHցAB�_ޞ�o_�E��V�χ\쨭��(�*��t���m����������ч��d5}�&���98!��E�-u�=��[ǻ�	�9��`_S�:n;s���Y�tv�<X�uɾ8�W�s�X��v�y�Q�V��ߦNG��]�{�s�V�Ç�gm��a89�����-|�����.ߜ���9��y�%��V�k�V�׍�{����d/i��Q����܇^=,G�W����Bf���m�T�/��ǂ{(GD���	Ϋ��1�Sw�~#)���2\���(��y���Hk��~���v;	Q��N*�yQx�����z<��fW�*��܍9"�-����/t��Î�L���eꑼ��� 7�}�Ei���=�k�oDi�
�8Ø�w����Þw\�GXE�>{�z�^�,ͤ�c9�N���*~����{=�,��n��Vw�"}���ƶMn����F=��u�:J���e��C�?*0R;缸���f`�:6N��{��݊��Rs�)e�b뻓��l0���DS��u�Y����A+ƙ���&��;��U9X�����ߘ0�8&Y;ܒ�@��y�&��l�[�l1�_c=��5��x�ې�ކiZ`�j��6��7x��ΐ����Ό�g�'Q����A��x|��3H��ѩS�-w*��7���� ҳ�}崏N����(ݻ�v��kE�O��r�����bT���{|���Ƕ����Ӱ�N��C�pq�~�o�g�{Bbi��P�:a}��1:ݷaY��"����w�+�����<�$�~���r+�d�{���\��Y�Opa�K�s0M��oXK������^s��tT��X&we���!�5�3�wX=.s������	�|y�9�s��t矇��k�Β�J���4����o�~��	�c۩:��t���y��^�z���ys��2��X�D���%��^5s��J�Ȥ���㫧U�u�GVk����{N���ɾx�I����*}��$5�`7�vQ7�g�5z�����վbeX��h���L2í��鹱vS�t��+����	A��E�׏; �����!��
ݭq�$��FZN�������	���؝c6�ͼW3��U�Y|��%���I��~+�	�u�.���������IE�\p�;ڀl�']�y��2�/ܫ��ov@7#�e1n�`=N��M&��G99G��=Lm�{i��һڒ�~}�3z"��q����Rq����^b#���:������1��k�ݾr�����}4��-������_�����{��%��ϖ�mJ���kv�i���{�c���_�-��E���t猝��R��p�F�'��ԯ޴�|9^}[��7��-�����񷫦��1�����3='�W�݅��v�.���^��`��#�]t�]x_�{��ͷ,R����+�h�=n�e�����h�r�������h�+��_�����S�|�g����i]O0�g=Ut�U�73�)�_հ͛��=��Mp,��z�IZ������;��;����Ύ��b�;<�ܺ��׾~qN���W�JQb��O*��#�EL5� ��f#z�&������^ua�齊`e�-�.p4ﳬ������Z��qH�ҝW:�Cb2xv8o7������=\@B̹2��bx�E�ܡ����9��|�����N!z:&���]#��r-�>7�FzV}ق@�ĳ���Ŋ 떇:�y+���P�)����<���8.�o��S&��q�`�&^N�v]|��ϯ��1Uo��A�)g�\�W�T��X�݁ӏ�_73|&Kۑh� ���{��l�[s�i�>��=�͋�|�t�����q�2���Kђhml�X&�S]���)�!UD��<iMt���͏͇w�̱&F"`�C5+�~�Aѫ��b9�믰�Yv���w�o��l�ވ���x[X䞜ǝ\=yϻ]I-��^�r��yv0��~/s��(���zn໸h��]Xl�"(}^0��E~�H?N�zpt��K����g��3�ڗ�3M�����&ծ����d^��o�$�������5ϰ�'�5��=I��2������Ou��� 5|4��ߏ�B7kxJ������o߼�p�'��6��a�	�|�O�`i'P�?o��N1@�<�$�d���a'�:������I�?s�:�ĨM~�u��}I��I}����h�����'��:���`��on�2�r����7��*v"�i����iCLgV�e��.a���׋}���n��Pꔝ��;�2Ջ1��=�Ro�\�~�{��7'6 }� �l|rNp�2�\�?:�pY�,k�O$k��N�����O�<��N�?B>���~�D�O��Y��M&����Ԭ�טI�'��d�'���6�:���ϰ'uNy���I��r�d��	���_����̺�Yw��u�M��k�d}����d�d�tf�J����=jOu�	�c'Sܳ�&�T�_`q�y��d�&�{��:�����`N$���{�Zry�q_z�
��m~�ﾇ����m�'̞��a>v����Iē�S5�V2Z��u��YS�N&��2O��jy�XJ��:���Oޙq���y�;u�w��*ORi�;�rAd�'{�]��X{��6�l��d�}d��N0�M����!�=ed���:���e1�|��:Ɔ���R&��y���{�b�����Q�O��4o�P:�ߨ{�rABy�|����$�,�I�N���N3l���B�O�Þd�'�%�hVN ��3�s�}��<��<�wͯ`|���N�$�'���6�d��~`q��������$����Ì�I4~�u�'�O?k���~I���$�x��,+	�w�}��M�ߵ�gu�t�	��>B�m���ěI�Q$�N�ڰݲN3�m���6ÙC����̝d����s�?0���a:�2|�O�g����o8z���������s�o^�q4��kX$����	PP���J�Ĭ�ei8�l���'߬:ԟ q���_�:çy�Y'!��&�=a6~�7�|�/�ߏ������}��'�=@��N3�OX���'P����d�C�k$�XN'VM�d�8��M�M�a8����C֤�'<���>��b�@dc�߻}+�����{�Λa+<a������'?0�>@�l*���NY!�'<�2N$���%J�a���o�e��'r�M����M��8?Wǩ��k�k����;����y���)=E�fO�}���F`9
n1t�v�|kD�7��Y��}����r��l薱�{Yw�.��`�!�WP���kV���R9��t�����Eﬖ�Rj�Dm�\����L���_�����w�����}��M�m���M0׿gY&%a��0�����ri'R킇? ���I�Ok'�'oVK�$��ԋ'_�>Lßw��L�+��=����IXOϩ��z��C�����O�:��o |�2u�o:�1+9�Ad��o�:��)s�=I�O����C�>I��x�t����TG<�0�4s��W�~��x����ܡ?;d�4e�'��ѿr�:�h��>N�~I��� z�2u�����:Û�PY&'?S��J�rs��C��B?s=r�:�W�{&�̝��<�zɯl���d�h�	��M3S(u���M~�!�a?n�'��IԜ5�I�4���}�'�:�}�S�I��{��r~��_�E���<���ﴄ~�y��6���N0?$�{��	��`k�&���'������d��O5�C�8�k�̇�8���l�C��A���M��߈��nߺ+��W��F���M!���M�a:w�8��M�$�_��'���$��@��'�d��YY�'SYg'�S�y��
I������^y���23�����[�?ā�|��?~��"N�q+4{�	ĝCA�0�4�u��:ɷ�OY6s���l����q�|�3Y%d�����x������N'�8''�z�˿fv��?v�M������@��r��)'�U�8��Ӟ�+�u+5��A@��ݒu��� m���O���']���N0�f�5�V2���}�0ޙ����ow���x��T��OS�LI>Cl�����&:ߙ2q+�RVd����$C7���m��Nr�׌�d�ݹ$۴�ׇ�Y����������O���VI���%a�����'PXyi��'A��i8����I&:7�C����~�3�N2u�gw�X���s�l�d�'�w�o�՗�+¬`m��I�x����G6�Ϸ�j�����P+�>��FV�)��7�~}�5���u.c�s~��3+j��w S�q�,�Z�]	K��*��^ʣ���ܢ��n苠mN�[�,������X;�E���)��׽��W�/�/g�y���d�'��	�<d��VI�xo̒��0;fЩ8���d�N2u4ad�I��}�l�	�~9�:���7��~igᰗ�UT�y�/;�no~�i�ē����~d�'�s$�u��OӶl���dY'��*
9fЬ�J�P6Ì�OL,':���������y��_�n�A�9��5s8�Hm�&���2|�:��;��=a6��Y<a���:�d�&�Ӵ'P�PRN!���*T�9x��m+'�P6ì�|{������|;|��������'��܇2��N0�s�Avɤ5���$��;��'Y'�6��yB�ğ�Y�P�C�O'5���I�����'����=��|�����|������f��I�O�8�����7�?2u��l�0��L>��$��}�d��N~{���AHh�r
I�4�:��Ov��7�y��O���?'T���]}�,%ea7�"��I=O|��	�����u�������O̜Cӛ�'Y?0���&2�Ϭ�I����Y8����~���:�QX.�o����!��!?K!��s�c	���ud��}����u5�'�����8�k��|β~aĞ�� |�d���u��
��xo�Ϭ�Q����v�Ͻ>�#﨏�P�~�%Bw�~I�OR��t�X|���Y'Y4n���N3FP�>�i4e�'穩�x�q���p�4��I���ߛ�V9��c}����gﾇ���H֡�؆�s��	����$�+!��rz�l�}d���O�<>�z�d״�����MBz�ɤіq�zʞ��/���į`(׮~�s3+|,�!�}�ߨB0��Ad�<� �I����	ĝa�y�SL��?C|�Ԝed5�p�'Y>~I�`���7�$��`x~����2q7o��翚����������klG�y6��F鐜h+5���+�û@��M����g�k6�g���ߧ�ɪ��
��Ξ[�N̯��O]2�y_y�Λ�{ܜ��e+��sf�H	��7���g��n�9�̣0�~Tż�'��R���(E��}�}^�X*A}ޯ��]&M��=I=eOy���$���q����m2u*~>�Bq�Xh�u4�q���N�o�	��I>}I���&�'_���~��������{�w��?t�����ed��іC���k,�	�*y��AI7���N�Hs��I�N�N��Bq�Xk�a�l��?́�Ԟ�>k��Z�>��o������9��w���$���'5�m�uњ�T�$<��d��e��$�4e�I�L�è,%}��C�8����'Y;��������ـ�u�]�K%��c���x�C��gـq�&�~;��&ߙ;�d�3�d�=H}l=J���>C�8�e�i8��Y��'��y$�+ M�X/�z����g�箿=K#��
d����;���By����:��'�]�6��N��'�N�IROY��2Jńϩ�+'X)��'R��o��e����g��j=��c�g�������&���f�'��?s�8ɶ_��^$���'uI�u�L4���x���a+	�<9�IPP�r�B�u+&����~��W��|�+�8��M�p�OXm����:��Bw�'�9�0�$����i��[�z��O�=;�$�i��Oݲa�O;��q�����^��ƃY�������o߾�	�֡%I�T�@�M�o�jya:��<?}��m���ϲAv��5�d�Iǌ?w�4ì���ܞ2q���ܓ��O���}d���@Ѭ�N�w���>��N�X	ĞOu�T�&M�$�6���Ru��N�:�Xz�ć�{���'Y8��s/4���d�	S�4w�~I���_�K�&�_��}��w�]��������=Af�BqY<��q���$�XN>vȲo��ᔜI?8��ì�d>7���~d�n��:�n�_C�t�U�da��݁��s)���֖�؁�eAwS���iwhWQ����I:2�����k�����ԿoLԽG�hX'e����:l�|'�,��vT�r%|Fe�����*��2Y��`��=Z��	��]���||;:�G�| ��s��Kٷ��~��!���ԟ0�&��4�����(q�Ԭ5�C�=d���q���d���9�����>f���I��?{a�N2o��C�#���N��ve����a�>d|��r��x��:}��	�
�7N��LO����M��5��z��>eCi������I�M��J�I���i�����r��6��n�y�]��ē��:�����'���x��I���/g��OP�9�:��|���d�T&����M���ܰ?2z���Rb=7�������m�~���=�Ɍ���a?;d�je�OSl����q	�����d�Ǟ�C��A}�$��P��ru4�>g�a�N%Bh?w:����A_.��ڄ����]���}U�_L��Ld���6Ԟ2q+!�8��{�q�z���I�'��⇌�Ad�oܓhq��Y���	ĝCS�d�i�}c��/p�_�Ր�L�?u���}����$�{I��d�d�u��+'Xn�֤�'P��2u+8�m�O=��I�l��'PY5�p�'Ru�:s��(qz\��I��&�wz���W귇{d�a�N�u���M�xq���'���'O�f�J��AC�VN����<d�k)���:�<��,%M��~y����|�o��&Ұ9����N2�O����<��v��a�@��O�9ݹ$��&��$�	���d�'�C�VN1I�l��'�o�=�{vs��}�����G��+��i�x�o��u+\���w�v�(M��>}I�Os�^$�';�!8ͲjwY
�>O'<�*O����v�����o;y���}�͡Y4�ö��d�jad�$�}��i�$��P�'̇f�'P���'�&��3�?2xϽ�~�G�#�>�}�"��j�W_��jo�Lt6�ibj.g�p��A��>��5^܇�Z�N<�cT��}G?zy�}tU�x�μwee�"�\������u�qf�+0���<�bAb�q1��P���$0�UQZ.��0nUm6�P��rŒ�k��Ü�}@�蓖������##�ʶl)Ǯp�}�}�˧[�p��~��B����y��(L�m
��ZRq&٣
I��O�d7l���8��Ԝaþ`|�z��̝d���;�x����1y�����|\���_��5�~g4�O�'�����6�y�%ABd��J�Ԭ�ei8�l���'�~�u�>@�?�.�:�Gy�Y'!����%�m����{����&�<a>�}ì�I��}�u�d��?�:�̝��8���J��Ô�
ɴ��e':ɿ)����|4�>�~�%�3�~��~���?[��|���t;�0��a��p�ì����x�ğ w�d��Ϲd8���Nk'h�쒥I2v�d����]}������lr��l���L�Zw���z�O4��7��^$�{�u�bVs�u�XLM�M$�
CS��(q��h�!Ԟ���x�q'C�������:XQ��+P����3��g���H�c�����N0����l>d�!��=~d�é=����'P�}��$Ĭ<9�Ad���N��
CG;�Ԝd�+�:�Ԛ��9�t�j���s�k�ֳ�l'̚Ւ�I�ޙB~}d�k,8�?>���C�'}���M$�M}�=f�:��sxI�a����$���'�k}��y��߽�~:������~�����?%aӔ��x{�|�u�^�I:�Ĭ'ϩ<eC�'��k,<a���x|�d�N���'�<<��O�u��5^���;�4���|�����i�z��N2m+!��?0�'��;;`|�{������m�����,'�4��2OR����u�O�,GЀH��o�P��4կv|77�Z�>���|��=�O�m�p�4�~C���Y9���w�8��M�$����	�~�+'P<�I�Y<a�52�z�:��g'�S������3[������>p�����(���-h.����A�x���B�O*>E�K��MJe�dm�L�q�^Y�uu1�{)�.��DS���Ý�1�H�a:W�A�vaNZ}��tb���g���-nj�q�n��
��!%��*���2���p<h��f��aH&	\��&���fW^f�q[[�5�͢���)Mg-�Ao"�g��:�����+���cj����:�v;1K�(56�a;��+� �t�Ϋ��9w�E����*N�N�4mds��=m�_�	�>ۧ��W*7�����9rK5�Th,۔{S�v:c�t�A�E������uv��.$��� �`���_���H� ��[�`�d��Յk�����a�qE=�סǈ�Wn^^�u"-~TJ�8��2���81��*���fT7W*U���*�ha��Wݕ�>�������y_���}ƻ��=�Q�У�	������1F��f�J�R�������E:I�^U�|�U�t��ZV<�D�.T7-]�����w0�Lf�&�P#����Յ'�,C]��"n�jub�\�s��2���ۓ};q���3��gY����1e4�S"�
'��G��T����16`�C7Y�[�"���W|�b)F%N���7v��eҽ�+�o �tz����#j���!y`�w�Y���qn|V��fk||C��M�ȯ���D�B��dg������8z�A>�]����Rd	{�*�5fv�חC��e[v�T�e<�N����S��D�?\w#�yo�]C��6!�����n�q�}�������/,�s�I�M���A�b����S�?�
;�͊�2�ͩK^�����wGu훾j�ޖ�p�WЎ5|��`�\&�ǔl���Q���m�*>C��,S��wa��o_[D�T��T�E󳝙�D�l�-�|³@s�C%�T�;�p`x2�1�������'Hw�z�k�y�<��~:���쁫(<4���+��C�3��P�^����`�����K`��S,e�>z���~����������.=�S&h�fY�Y�2j>�.�*�N��#''w{J�qvLǭ٤�ܥ,'Z�����Tw
��<������7Z�Q�ZS 귚����8q;�R�^ǵ�;j5��+�����UvDP7n�*��щJ����]��40��p�i�L���)���;�Ruh�@���
n��TY�ug�`�'eދ�uX���{��;'gd�V_90Bs-(-ŽkS�n���Ug<v��Ĩ�N��pG�Ǩl��.��6X뷹yjֳ(���芩�W�~�Ֆʁ�vgY�N8ߎ���������iېb�+���aB��ii.+Bw@���K��R��gy��B�,�4�`��8�b�gghfN|��nI�0t!�o��$L��Mܮ���.|�YZ��Z�T��g�B�11	�"���E!X�*eV-H�#lXV�QJ�,�F�c&0��*��¢��h�T��"�lV,"�P��"2���
�c
��"��
�V
��BbA�YRE��((TY*B�6�"��(µ	Z�Qq"���R
VV-B��ЬT��T�+D+�X�J2��)*,
ŋ	+3"1L��X��	m*)%jJ��Q2�@�kUVAb����J0U��T�0Xe�Y*�RQ��"�Q��
�-H(U`��LC#�"���+R����@���"֥B�g����٨ϯve�u�tvS��z��.��EvyLU,�2x�<�$�B��!0��Oi����i���:���������=��\�z��|,�H��h�!i �?���*N�u+4{�	ĝC\��L'XnӬ�$��s�ΰ�;d��쓌���d��`~���VOq������7]~8y�|���m������ve�I�6�O7���[�d�V��p��Y:��?w(C}���N��y�6�I�'�,���6sY'N3�{��￞��������\��vJ�L�KC�Y6��k)!�&�YLI>C����M2Ltȯ8��ϩ+�u���{�!��紛d��s ��O̚�ͿgZs��K^��ןs���'��w����|��$�>d�
��,?���u5��i8����I&:7�C����~�`z��N���w�X���{������wz~7�{�����d�'}��m�'�O�,&��'�5�����Y*
]�hT�AI�m':��Y&�q<>���i��~����t���7���Wz��X�ߙ�����gC������|�w��4��M��I��'�?��M��O'5�d�C�k$�(N3hVN�d�2��d�k	��M>y����_w�}{�o��{�/4���e�z��ܐ��'�Y�I׈p��OXM���:ɦ�~9ܓ��O�i���x��()'�sY"!��#{��,~����,���/��A}�{9��|�`�q��$5�m�����MN{v�kP�C��-��9�s	�ϰ�uh�u��f��û�v܏��Ŏ�r�X�T��ίj�ǥzZY���F��P��>�J��Ĺ�y\�B��uk��pnA^� 홿oR��Qg����8l���RJk_V+�".= [�X�Twj �X*�^w�Hcm^��,�OL�_��oM�����J�n]<K#��/bb�;W"
�ٝ�V�!��U9�9�'J���Ǚl�zo���t؉����s{Ώ�e��su��*j���=*=����q[Iߊ~<������K��D���(������;3�b�Z�C[}�Ta�s����ڬ���YR{[~�z��%������n��hm�;��2Z��&����K�ƲMD���R��u�_��pe{�+\jU���~^�Y�ʆ���Æ���&ش�s�&U��������réo4�n}��_*=Hz]�5ݷ��<X�k���S�^�_v��d6G�!�R�V��3���qԡ��ɾ��w�omY����v�
�_6m�ƎiB�u�9���3��xd̓���ӏ{���Gh(��K���u���sZ�/�����㯗��ןo��T=�����XӮj��.��63����~mG����͹���9��=}c�+&I����v]:#�;_�sS/�F_TZ�۶n�S%j}�[X,�e��U�pd=�a����a
��aB��b��;5R��ˤ�V���}��tl������e�~��N�N\O�������p�׮�Sȭ&�¹��\�.:�-��/:��|%��yt~���{�!���y3[��#ڶwx�����{#�uk��Ҍ�Hz]���G�t��l\����'��?}J(W��IFV��?nͮ�}tI��c̝v�]��H!=�+{�y՛����5E=��7֋�a�ϻs��n��4�#)�vơꙨ�Erԫ��ی<y��=56J��n�t��ͽ3n�y��q�p��{͘�̯U�~�=;�oO}��8[�zpt�b��/���|���������C�%�Qy,{�nx^��϶zX�ױ�=�p<�X_N��Rj�5����m�����~��ʷy�b�f�6����3E�{1-Hh˕���u4�k�����N�q�-�a?Rg�f�W����4\��uE�h�n�y��^�>��j����XO�^�|$`��@�Z������s�^N挣��+��s�O�x�ۗr��;q1��LґPozB���MXN-'�}�����;�4�%g��.r�ր6ӫ���ZR��]t;֌�rD-�Bג���֠��<f�Mǎh����J���mu9}Ue�u.�����4<�|��I���yܩ�����{c�Gp��az����g�",�?A�ku~�� �4��C�M���=>�8��}����cЪ<��W�pI���ݑ͉M�������o���α��'Ҏ�ͨo��~[K|f�w�=��t����_nu�����L���w]s{+_�i�����ۓ�.����tB��}a����~s_�o�snizx�j�Zu7W���q���^~�nK��:��aӲ͘O>�=܇[��!�6E�2aU;kt�����:����$�A�vJl�.u'����v�U�G8r>�{��C����L���>�׃y�t���Lg�_^:9U�dKEw���	>Pw�w�s�;����[�k�Ň𾞧t��N��R�DS�~J��V-��Y1��[��u~��}ꏺO`U�1ny��,K�CC�������\Z���hnpwO����ܻ����\\��oHyZ]�������N�[�N�N5��Q�=;�Y������.�_������a����mL���˃)�k�=�,sll�g�m�8a�J�R_�è�)�n�����NN]_��ﾪ}�v��Wa_�qj6S ��P�[�I���T轵�ԋ1�����{W{w=�z[�;���ޯ?�q�[�/f�[�ڑ޻��J⯷�F��n�I{�=l�����+O��u�b���{���WL~MYM�էy>��n���N^g����k������P����̳� ��������u�k���B�l;����:�0r���ro+zhʚ�-߄�*j�<�C���@߾<��Nu�Z��p���A:N�������%ѥ�Ǖk�+�O���Y�au;K]��G�:����
o�P@�
�k�U���)=�w���=�%�h��Ɲ��K�ݒ�y�$�}{�VwWN��hUi�=u�y3��Y|�������r"��8G>�s����������~[{8즼�z�	[�J�nG���Y���:��	�\�e�;B�-Q.%��ޛzG���\2kq����.jt��N�[�K>�zbN�U��{����#�(_��5���BO,U�����F�����t,m��)��=1q��s$9]y7��w�X��Q�p�����20�ntV��)�r�\s�UU}�y�}�&]�xutjOo�gΟ�_�>��|$��tM�~��o0P�{�{���i� ]�W�4/�kϹ��ϤT�)�}!�o�������r������AvJ��
l����d|:��&����SK�g���8������qXv'ϽN��˾�^+k8����I&yt~'�</k\w���F��n�᷍�h]��H���Wn{a��Mo��jG��~=�J*��FѐE�W�	�ޜ�k��2�{�{˝��e���<�rۣ�˒[^�O�� ��)��s���9��O^��m� �����(ڪ����_�9w��А˔���H=|}�����c+� Z�R�8��{ͭ)^�x5o71�<�n�>��Ϳ���'�B���F,w�Ãm����z�����}���R��W�՝���Rת������xd0�z�O:�=�����+�\�)@6��Ә��Tœ���}9u
q����<���K�+Vw����4û!�������Mn�#��'�JGB�S�
+h+��=�y$�I���1���4ͥ�Lxt��էY�X����*�뚪�u���������t<����I[��幸���c�,b=Ύ��k=A=���j�b�!t<�f����>����.Ms�.}�N=���|0���v��1���ꭗ�Ϋ=�UG_����!��ҥ�_H_�Y�tBŋ��hj��%-��O���=�}�ړ!�[����yR�����xp����%l�΃�"��_'�GOnqv�=���eg���o��/n�OĢ�b]��yk���۴s�C�/�.�I�͋�����*��Ϋ��I]�����bv���d��d�BX����=���7ٱ��ûч56�K٧z��ٮ��@]1n�7�I���A�Y}�<�нJWm=�ua��)=���f�F��*ÖŸ���;��m�홧��!��#�	��Z�z}�%��mG�4��?N�zpt���gO�Õ/����xY��]X��xo��iQ�DƻlKE�bN߰˔y����]V\y��ǡ���d���	�������㯧c6gk���ʖ-Qx���t���2�xt�9�m���^��{�'�)�E�VON�ݝμ�Iभ���?W������h�_�v�~����ܞ����=-����'�O�)�O�?oc�-�I�=Ù�7�]��v����|�n60W�A�o%���1T���u�%vo'癞1�{��C���L��j�L����
��Eˡ޵�3^w�����^�qd���9�|���8w�;z��Ưj��\w>�$�Q�m��H̻}�M:�Ğ1���S�2g���_y�gk�|c>N���eB*�9�T���*h4/�L��	]'9=s�m�o��u�����mM��4�=�b�}a-w[-rl�{�7��γ��y�N/�Owk>��ء*I�ѾFǋ�;�t����r5\��p���̿	I�{/��-�\�{��{T%�_:!N0Q�ևJ�s���5�	[�M�Z�E�;U���^�N멾s7�<�����v;!6a<���܇X��8T㺷�RG��]�ҭ��R9P��s�97>vOvV��r��E+�C�T�^��b��q-{����-��ʏ�ov��O]Lل�_�������!�2�l�/�N�}��'l?E��'U[v�38�9���p��%c�V`�K����.�|�����Mf{���>��H�;K��J��6��A�)�Ɠ�Wt<������r���>��뿟3$��]�!�o���^�%���Ov�Ǐ�vzU�ڮ�_w�q�w	w��#A����{�[�qы���^0�����} �|j��g���{q���s;�4���`�9(�͌�@m	�]�
�r#����T
��+j#�T���3���z�o��7�����t���2�ϳ�@�nO=9P��j�U��n������я}��}��&��7F?o{)�>��;K�c3��~��P�s3͞�t�����]S^nM�=�Vәh��-s�N^g��3��z<�W�QW��;W��{�:��lfz/xк�B�F/�\7����\ϹN��97���7��j(�]u�%��ٞ���>ZN��b��p���C�M�:ג�VB��^�ں�t�幧�^=�G���*��ȗ^	oz-`��>�^X�����������f�|ٴn3{c��UhC�ڑ1,��
Y�ny3�=,'s^��ɯ���G��AnC�<�fy4-TQ'f���&ò˷��9��ڇ�s����������v�7�@�MWV��|y��v�����.l��'�Kv;)���>N�����^s���d��r�ӣ�x��O%�oIkg����;�6/5.�5��B� �*����;������>�!N,P<劜���7s���������[��L��=�Φۑ�g�$ʜ��a�vB|a1{�C� ����q�7V�K�}q�/��rW�}%T���շ\j�j��a�nx�Θ�7�6.y���Ϧ	W|e=��Y�ʯ����Wo����9�C�޲P�e���V��쏇S݄�nGM�e{�O����'�����U橪�U۝��gμV�q[�^�I3��/tghC�=fe�ޏN��Pʮm����u�{�;�y��������n��t:o932ߵ�n��o_��>�P~�^��;3�b�l� ���g�>=DT���<'0�O�tE�w��$`�	��9׃^vw�7�z�mѧJ7��n}��Ȟ��y{��'R}"d�c۶�:b�'�
�K�0w9f�DY,��������5a�`�����w߉^�L�=Jt�e��C,�U�
���@�����_>�,z��PP
�'��{�����<����|^�A�E���x7-RMZ-g"A�}�y��שՃ����!��,QzվF�u�v�s��7 ��^*hI[�G-QUQ��:��'M�K��|�e��}U��-�Z'!ٹQ<�v���ZYD �W7
�D);�˺�%b�[��+�a��k��wAҬ%�&�ګ�I�Pǚ1��䰕{Yw
� Ωr�cB��p"���w���hc��ZE�J˸u}\xRd�C�o:�#K�6{c��!�����^�o9�{ǋ��A�T�I�-滲YW��������I��g�3={S޻���4vQ��o�[;T$t��͎�����uו���C�yK��q���;KA۳��v���6��	�+s.��q��P�Y��^M����X4l!c��(�PY9�P]'9��`o9�d�U������5	ƞ�z�R���.����OP(�l�9͑X��ME%��}i��Ts폸�{�s�q�l��eM��	����9G�"`�%���o�	�Eϵ�u�Z��=�,�/\k
�a�˚J�z����}� 0F�3�3�A�a��3�V��	��r�W
���#/'$��5M�qe	ֱ�3{c����Q�q[4���7�^�+����Ɵ=Get��O��F�p[�8��%J���K�W1��4A}��/ݼ8�5��5Hw�+�)B����׉]��%3���P�<r���s����[����=���7D��o���w�b���[ƌ���²ٹH�k�L�n@:4SUovQy.��罃�Yo~#��Bedl�~�`���`FQ�;X9�]�Z0rj�44�k]�:��P.km��E��9�X����q�]��76G��zOARvnyK����Rܞ�n�W@}k8�c�3�{e��b���̱m|�vvC��тL:��;E���>��n��2���q��E[;Wr�����TB돦�no&H��#��u���s6�[�c^ax�;ވڶJْ�W#�״#�pd}��#:޽��&chX��u�H�wk�$��8	'�*K��]�8�5|V�g\@�׍���sOwA��|վ����@ݘ|r�[h>۵��*|!օw��ՑH�Ik�p�&뻲L�[��lʦ8-�)7m��;G���X.�!˳G;n�e��$�b�Vb&MvOj4s(�*�˻5��X�w�r�>���q�L�Q�"������6k�̝|u<>�<O=]cvgj�d������������LC��PT`*��E"� �`V���Q�ԭ����Z�YP(���FJȲbH).Z6�PR��d��P�R�*����DR(�Uje��j�"ł�����Qj��-��%��TUIP����
�bVQU�
��kEG)b0�(�T���[+�ŕQJ��P�
ԕ�,+*�UKlD��+�Ղ1R�Kmeb��J�,�`�[T�jE+*��Ab�(#l���T����V0�2Vƫ�Z���e����Jʅ[Ad��aD+SQ�H��J1`�Z�U
�i�����+b%,��Ҭ��KjѢ���TX�ũP�QTm�Q��j�@�̢¢�RF�4| AU���_t3y��L�ϓ�ݵ]3�8�V��i��.�B!V�2�Z�v:�[���=�D��U���]�k�����&���:D�?�L��m���p`���ױ������UX�����`q�'���3����񯮛��af���R�9�lOI����L�~=�v��ꞐEו�f_g�;^v_���z#�p��-Է����ɢ��"=�7ν~��5�Vs4f�L�C8��P�.���e�\��֨�O�<����=�H�E�ӏ��v�³��?��%��`52�LY%�%���Iu�鷞{�	���rk��٧}c!����=ށ�Gk=�6�����>���%�Յ���7�d77�p�ݒ�,�|�UȈ��A�o�q��a��[��Od^�����q�d�1Ͻ��^���qp���ܵ!~�hQ�!���:{s������Կsr���OW����C¼iL/��c��RX����K�U�{Y�sǣ���wp;�v�ܯ��ٗ��?>��39���ee;x���
n�OV�7JM��	jn-�6姍Y3aQ��� ����nQ�ɋ:��i<���������%{�LN+9�����ס��N�z�����}Z9B�9QA�{)��ri��}����NN\���߁����^��jX����@'��W��lw*�ݾ�W�n��S�Sq�oGc��9���pv�j���[ ��؏C�L�=h��E&�p^V�ϟ�1������+~rط���ӾÏ$�;�Ku��lS{���a/J0���U�o�9�{]=C9{���w��\p�X�ǫ�U�Vt��S�3s7�]��~�Ԍ^��͞�����pP:�9k�u�B)W����"��=�Ko�����Sޢ��#���e�
��O��^�O����$ݫ�V'yƙ�^	���Rgǲ�VO���gh�[,����{z)/3\{�\�����fP��߂�h�{��_�gΜ�KW��ζx�nk��t�Ԟ�����;��?b��֏��=��\���x��Wp5|���l}�J�9���N=�-��R��z-�Vr�Q���jTwuo]&P���a�jaV��"7^b4oiV�f�:V�� �[�r����m�ˤ�pv� �]ζ7j�6!;�&�J���^y�o҈��t��Cr�>L��RYV���s�<���o�
�R^��ʅL&��˅#ȹSz�����}_}�T��ƚ�b�����-�[-_Sf�}&�l�{�M�{{�[�Kr	��{q�>=�e��Gh�>���nu�(�s&�����.�Z.��o�ӓ�.�-�{�v_�'0��t�����9�'_��/J������ſH����{X'U|�vv���ן	��`��5k�Pn3_�����mʿv|\���$��Xt��l���|��R+�?oBOmJ��g���sv�e�2<2��V��wN�L�۔x��2s�xJ�>]�Kg�{7����nE��b��I�d��\�K+�n��F��u߫<U礿{ۍ��n�`{�շ�OJ�bI����踺d�~��-�M�\��T[�䟏����wL,ym�����:t,�񞡕\��{˝�VU-]�*�u��s���6o�E������5-Q��1�*�S�w	��n�Uj����l����T�֎9��q��ñ:Q����'�@�rry\V{���q����A�ʮrD�|zm�5�S�P����ŉG�����bb�	,�/G5]�ˠ�ffq�� >���:U[��m��L~��q��c6�����g����g���r����fp��\��2�ޱ�p�/���p�W�w���o�=��r�]��g���8�pnOV��m����7cGx�o�ƥM��5���|���_=���X��W�{7%sa��{�C�[�*-s�B�W5Dq��o`�M��	ǹ�z����u;K]��W�\ٿ��U�٘tw�'��5����=�zq5��α,�:;@�b��O?
޵jz�V��&�ML�no��U�ᕾs�k�C��:>΢'0�j�1'\5.�~4CW�v����\��1Ӟ~���u6܏*��o�.u��b�'�Q^f:���g�'��@�w_�IB��~ܜ8��/݅��|佼�J�ƺ,;&n�C՗5�M�l�=��(��S��sz:���U�<z������R�æ�}T�6��G{WH��nGF������=OO]
�Ǌ��vΡ:�gv�f�h�V�]y�� {2�Q�X<��TwΠ,�ó�T>[�R�毪�+�}�eVt)�{���5��w�5'�������j�|  |�F�<��.��=BX�n3�`'���w�d�a��'/Q�c�n�R�Z��:�(��S��yv?B,�KuK����ǥ.w��Z�Dѭ��;3����l
��,8���6��>����~l����|��+�sL��ۙ:i��*~���y���kڽ���l���J�6�����	z^K�=z��:A������|��0	����-6X�^]\t�~����,T<�}u����W�A��Xu/0s��<,wo�����p��[���*�as7�;��LP���s�6�0gq��{�U�Y5_�>�����}��-Y��q�k�-M
�u-����Q�jЯvS��/{��0zs���G��ӏ��ޚ;��&N�6x��}�Dw���f^�2���2gz	rk���	Ƕ坧GhPc��m��W�-*1
qi:���'4н�ӕk�dن�t�LE�ӣ��,PÉ��U�OV���v2�;�V��-�G������/��D�75W��yF7��Ϯ�ϯk���cc�^� �j�r`�����u�2��y@����M�C�k��<��������r��_�#ڛ74N�߹��O���7�g�;�@�����+��V&�5<����j����Iu;���y�'�}4�����s}䇉�ׇ�X�4���)I�N�����t,�\��C�nqv��	S����'���C�{�z:�wKm�/?@7%�����aӲ��ƾ]:�S��6.x��F{#��ݢ�;V�o�]�IW�����g�mK��[<p'��W�T�溷k|91��N���eɑ�2�p<���;�%Ѓ�)!iCbё�&�8��c�o?o��<�?��{%[�Ň񾞧t��|z^z��t����������/~�+j�>(�zWI�?9�{��3�^�����\��j�1�n��Wa^��z͗+��x�0����y}�o��/t�#��R�����_�.�]�5�+*��ڕ���[|����:�R����j�? �|��q0.\�MK�򧢙�v;���)�q�!��	Z�^m��{����w��]�i�j�Xٙc�t�[��;q݄F�A'��6wl�U�����mw���c�Jzv���OA���}x�� �pȍ׼�`�g�~G7�,���}:ʓ[2u�����;���{2�êsB�s��_�]I}����d�lg2�k�OG
�8'/5��5�ڷ����g�f���U���̣�G�o�랮���/�@�d<&�a�適=����Ƕ��;�	��r����Yy��Ֆ�c����o�:���P�9���}8����ly�6@-M�>A��b/�R���9��ٷ��}�!O|뫭f�E�)��}�s���q}bY�����b�:����A�=U�w��%$�K�1#�ǒ}ϷI�u-�ec�e�E�0WǟXC��/��W�qe�������䕾��6܏:��T�݇N�M�h.}E�˴�o�ۡ��=˯xmI��z:?����+����@K�Ʉ9ޡI\b�@fa�f����Q�'����g�x9����2���OpHk�����W�t��q;�B�z����|ΞlM��x��{������z�e󡶳�Rd���+��	lJ��������^�.o��Y����t�/T��;�}l��-u��6��L�ӝk�������{����K��4�j��;���c�w�5�v���2�掾�~e��| �\T�qT�^��f�.�M�b��{7p����܉�c(�y�mQ�g��s���X�',�ےm�:�^�q[TW��&yt{�'�5��Ұ��L>Ǫp��}�nh��y�6W�^��lG��~>�"�~���#�g�zA���&*���OP��rgx���W����o��{8ٞ9�݉|��������8>�暈�3�r�>{��M�7ko����;W��u<���t�Y�z�co���u�8&7���Zr� ��s}W�[W̱���ݒ��+�Ӌ`OƮ���c����店3��k�~V����W����7��gKV{����v�u�_��d62	�EL��Q�p�������`zg_�۴�!c�tus'9��,�p����G�P��^]7S���`��Mu�Ny��u�;A��Ō;%��ZDFa��$k�E{|�+�rW|��[r��z�gR����"�v6�sO����J"±{;�+�W~�|�".Iխ�G)��b�����Yܳ�gM� ��qu5��7[�*No3W�p��os�g.#�'\�Hc����t�n]��'O-�W�W�Ut}�k��[7��}������9�?	��xS���!	ŋ�W��lOiE�z�w�/���s9��+}�Mr;��&T��4�/]+�'k�疻������JwZU�'o��ӏ>
_� �;��<�2�=���2hE2��s��g�%*�h�+yĵ�Ü��5޺:�=�{��]B�W���ŵ��f�7���x��ix2)ؠ��$23]��/��E=�r��/+��=X+5��R��ѽ];1Z*�t��4K�w�hC�uD3}��w�����>���e�`]�J�y��t
�M����R�z���ޘ)X{�6��n
z�(}�Y��Gv6��צ�k��M�X�!j���zz�Ͻ���_-�:t��c�,U��"Y�:��;{Pڢ��GU^���W����RPl�Ӗ`��2���@|/��t��o�f4���Y�=U������L�w\�j�k���t�X.?N0.!E��#�_���G{4ߦP������j�v���k;=�X� ^OGmmz�������a<���db9ˮ�0�Au!#�[~+=ho�H<��܇oq�x_e�����u�q���ldH��%�@�:1�m��<����d����J|2�ٌ;�xL�Ո5m�k5����o%��l<��4��y���sէq��V��q`��]�G�][�EB���W���R��M<�.d�',�zϖ���y%{˯��ee��j�Gi)C��ZX#,Og�]v�J�^s��q��N�JM5Y^,���P�:�=��N5���g����kMC0U;QQ���;U�6n��z���L���J�,+�D����L7�)����q�ۂf#��\S��4��q&�	��t��CI3:ꈮ��+���Z62sɡU���V�]%Nz�^袥~�acL�&��v���ԌWPL��0�ٕ�*}�Z�Uî^��z��U>�)��Fob�3��Yk�%đ��v�g��{��e����Ґ	�ּ%��uu��)+���g��=��Z�a�k����9����t!�rWK��Ϯ��딜O�#+("y�>����qÏ��{lI�fB��qq�Cz�J�e�0��l�K��OT���ޗD��x;�o�DVf����PIF,ϻ�nJȃ�2��P�E��c�g���K���\RÏ�3����o�I�ynл�D�y�^9�ی�<�,c3����s�lݦ�c�˜f(��p�7�G+s��ժ6ӗ���A�v��^�+��_5�$���3*��t�9�����Xq��_��W ���
S\� ��F����`j��XԸ�S#*V6������[ܸu"��G0.���RCAE]���Q�r,��f�8&��srh�\6I3�φ�(�Xyr�E��(B���G-�-�o��q�*�2���oq�Ffn��%��"���Ox	��u�HxwqJs�z�.5�p	�M#90�j܅����։N�"�GV�R<ðM�ygxC͂�q����g��i����V��k��u��݌�ˀ/��L;��������Lx���)���[�:6��i���\ʅh�Ŗ��m��c�+8��y%�0I��F]s��4��F]����'z>�1"y�J#.�$�N���#�V���a�ٮ���	�����D��(o�_2M��bo��%J�l�f���L�����vc�?oW��G =��lG��"O�oøf�y����wL����w%oH<�k(˾Y�=���u���Kn��4���屽C$n4����c50��o��Y�1fes`�/�Wt*����/&?r�ք�{�S$�{�������2��C4��G{]}�M�;�ҏR��'Y�yz7w�$ީ�gsWQ��miķ�12�|�ԥ�F�͑7�;�YY�9l�=�C���wD���ho�JyZ�T���a:Ȥ���)'`9K�jZ#��CV�+�g���Y�S	N�lR��֬�N��<֒�4 �{��&ɝ�(��F��"C��[�:�'?�����`�]2�J/��$��7�h���Xd�������o>,������x)}�fn7�� �\���h�ڤ���R�=;�.3�m��\�@�:�סr�b���42�+�י>Vn�� 7x�ӑ3����*E}�]�c'M츴9��mj�	-JU�tl@�)C;�}�P�oޛ;��'�}4�N����W�����FL	�j���8Q[u4q՝��%�`��x("�U�BIV@:�v]�_���tzY[���䯝�ϕ��6�Wp���-��"h�A��.��{�&����b�gW�E��0eE�2\���2�˞`�7��4�F&VӋ�d�kO�]盘�������^�+uQL7��S�ͽ-���W�����nSkt����R[-b�K3y���P��,�mE�4�YWaWPRWM9δ�F�](��O���'wF�fը��H��#���x\���:#'�,���GZ�D|�Jgm{�ǟ*޻�� ����T��/뾅�<x�T�'�e=����^P��:9�NC�Z|o_�v�������
� ��6P�++30�+Fkd��e����E����1L�#YQq
�յ��Q*)Z�e ��mJ�F�
 (�m%�m�Hڊ�j�E�����Z��¢�X�\LLV
)R)QA`�Ym�6ʄ�l��(�C2�B*��Vжȵ�°��,�Qeb*���TX�ȳ
���Q�!VءGC+aR�`1��(1B�
��@�E�,´(���PU�B�aD��Cd�E�)�YX��[j2�,*3AAC2�d�c���XQKj+�LJ�`��j(`����YD*�Z�*��-E��j�V�A��)R�����kij�b$R,�6�-`�YZ�KQ���b�j��0P��k#hUHTRQQ�P�DPwg���9�mwf7��gnrn\�P]�ĺ�ЦЭm�1ؘOI�
Z�������ĸ�U�e�ZWI�r<�}��U����藪����R�m3�}Յ����{Ü�I\�U�����֬��:T�N��
[�؝���rE~K{.豿_Y��R=f�ٞ/@\z�9�/�n
�m�!ǂ���:ͬ,n��ѻ��X�>[{P�K�j!~]i���ȡ��\W�S)_����$�d���>�.ԙ�w^��lvpLo̽��T����NzƜJ�}I�X��a�"͜�'y�e>��>��^*:^�h�t=��k��	z*��>^u�t9�~'�Q�od�3մ ��pD:(���)������&��m]3�kC�U_3{CU�Ⳙ���i��~ Ϊ��E	8���Υ�]�s5��p��z1L=5<��۝w,s1J\�Ui�YU\f}0���'^�2�zQ�̝L���iJ�]��^Q���!�u`�����iP�v�8�t�W��0Ӫ�#�N�W�(�o�^X�e���'��'�>��[7��Ó�>R��*#I<� KZ�(W�N����|�3=Ğ\�{S��GN��ݛ���=�5:U��1�E/?+��i\!����S����ftP�wy�M��'������_Z��!&�0G+[g޾mrv��՝L�B�/�U����g���y{����F���u2�R�K�t�:�k�?}_W�M�u��9/a���zu�+>9��S�-#=��@�����w��C��3I7�wD�7<��/_+��轲9}�_��E���FIy��f�L�a�0�5%"N�J�t��m��i��!�؅j��_�����^j����-xp��`�l$�Z���=s��x�0\��%�u/����_�;-f�ʊ����cN	)Z����*�c�e�\�<��
�>��oD�-w��WW�m����{�f,87��V\R򹊀�ï����o��{�=U~���lE<���xzד9�<�>�c۟&kשbk:�pw��y�±��o޷X��6a5n�h�2�'G(v����� �f&<s�I�exV��Ʈ.�4G��̻~|�|��{�P��}p/c�D��KV����9��T/>���;��7A��I���6�z�ib�������"����m,��s�����z:r�tT�Z۷��ߺ�j�%��->J}�.b��=�Dh8�S���������@�,��O���ni��c���WneF�P�@���bwN.��dV{r��O-U�o�}a�i�P{�]Y��o�@N� ]q�9̥�"6�o�j״�+��n';���K�ۀ8���)���Z�Ǟ�6s�M��g�����6���*�WY��ࡲ�JJ��x�-sv����a'"� w/o��g�/�$s-�Y�ʸf��:�J3��V
\_��=�R�3.��';��R%��?U�֒���������vH�n�C+���*rs���顀ׅЭG�ȪΟ<�����w_��]����<�����<+��0����G��o��Fi��e#�.��a3Px��B�l�]v��ۭ���=j��+���p+ə�};%!d炄�[��~��������Vk�H�����Aֱ
�͠������o&���ShXr<��d�FT�Ԯԑ&X���I��k�z
�=�QXe�"�yXm�W�}S/K�P;.�5���fB� F�/w�S�1���KO<����j{w_�����Obƙ�u����U1wvs;Y�������]��}(^�dPv(;촐��w�}N�˪���B���U5�]��M�p����PM���P��U�M�)�8�>�Q�a4�1n�tϷ3���T�t՞�4w�NW����o�ž�[�i�����6�L�Q�K�-�C{�Oyc�Ҡ�Rh�E��[;��Q�tƷ�L|�/N֮��ô\�Iw<�c�*R��Xy�0�W�1�v)7�x[��8���#ڞ��׏+�  x���\9��C�=ٞ�c�#7��]�܀Ѱ\LpSԹC�Exr8��vg��!-A����Y/�X�}[��	��*��W��2G��L�P��m&p��p�9����V.��3iOB�{0w�\�z�4��(.J+E��7���e�;P}^"���cٍ$o�+���[�yJ��W�Aߪ�z�pa5���O���q�p��q�������ڕ]c�_J&��ɔ�|�����Pɲgr�^>yJ'�\X)iYT���f����y����TPk�M��I���%��x��c(v!�9/uz�\b�Fʨ��а�V앙�~�BF3/܌�by�V�u�^J�Pŕ�̿������j�k�q���f����z���l���?�SoGj���b�J�"�w�M-{J)�ل�c���ҫ�8��Ϧb:{y�0��z�\~�!������[X*����슺�l�E�<�d�o'<����|�2�h�X9���u��ޡc��,���_l�`����,��9��%؞C%z���q�}�+C����`֛�0*f�e�i&�Š�G��״���B���/;�P�!TL��$b�f[L��_L}wr�CJ>���6a0ܢ�ٯ��L�t�l}����l��{�k��&�k"*�چ޺B�����[g�ўw\���?�}��	�d�09=��������|�T$:�_3C�Ӳ�qض�û'�[�I�wC`�AUn�9'���u;�IXt�zfqȥ!@��`�5�#�u��힑{���W�\��\���e.��<���J̅�ʸ��(oQ���v��d�`�$6��纃��*"�=͓��\�����9(ř�0#`IY~]�pC�%C�&]�|>ya0�眯xm��Y`����a�W5�.�A�[=���������Q��(̹�&E��H����K�n�D��d#��tXھ[�]������,'w�R-�X������ޜ���NǃA�Y��Aᬽ���	�2���E�״������ �IS<W�wi��t�n����#&Vrߚ����/F֥"�s�ΰ?�O�z:�p�����-�\��>��j>:�<G�P��Y�k��	z)-�V;ߥ�2u���zJu�v�*ǈ������b��Ե�G(^���b���ϫC��Ogz�}V�iإ�	�v{غ}���)��]���^B�2Z����s�F/�2�Ŕ�{��YY��sf���6s0.��:@##7l.ptb�x)�fF^V��_(�M�wPΛ�D�R��w	��4��O%�����p���7<Y�;��Z�e�`gAb��(@_��.�����|�\b\�I����[kU��#��z�u�g�L8Ǒ�ؖ�)%��羀�M��d+���'S3*ի\�~F���K�c?~�/����Fl>Xm��*��A/$����/>�\^}}3c��#��ǘg>�.��k�/��5�܋~����f�ßN4�K(v�#M�&�����VK�3�e��t�m+N��
�D;8��=^ǲ�'�����CmN*�{;Ṳe˴�x�%�wuM+=�q�,����������aԡ~u59[c�%X�-���;�^r�Jf��0�L4Og��xt�ɇ{.��ǵa{�A������1�ߥ^j�����G���4}6�����4��i��K���GR�^������>���OL�v4ٽ~������tks���X#�5_�.���IT���ʕ�U��/L]n��o�$I���c��M����j	ٚ����.����'g�C�CU��L�f�{Ibk:��4N�~����g��_������BR.=�p�-w�`��44\̶����\n'�{~���k���8��FL����o��W�*��Eq���e�Lܜy^}�4����T���Vc�Ft��F�� ߸n�NݔuY��P�z��ޙ��=��Ԋz���'~�-뻗�M�� �bcƳ�I�����y���Ҧ�x�o�5��Χ����(<o�F���1?%�ux��Xg<2�wcg[�����8�A�`~��V�Y�.�׭V��=I���~�Z��SJ{��졧O��^�zl�l��޶:�aq��xڙ�Pt`zzz�wϞ�"�]�9�=�v�ή�q1�<�Rǽڷ8M.Z�V�UCe�O���O#���"v2< _�	͊r��49m���5e�s楽]�W�iO�f|�>.�`�����ґX=��H���b��zw���=��,�$��.��O��KPά��Z�B ���
T5ݎ�Fkݯd���?.��j���v��ג�����L��5�8$�~^3M��H�˴x�f�#���_�����{��̺��1��Y3����fzu�A���Qɕ���:�n�*�i^7<�U7���ų�2�و����q���l;y59U��?�M�|�y�^�P��y�xq��)�N�!۹�{{���痸�j&�3��^*�����B>�	)@.⛜��ޮ6�5��/*߅����{�b�U�y�d���Y;��f�0���CB�s4�s
�{��M�Hu+Pl1��*��Y���֧�o�tvv�K�I0�u�>������c�9hx����<���I3�
B����:�3�v�k�2��#����W�\��J��䭡���U�)j�
�ZJ�n�i&�w�p���=>�`l;��z���k��9�Y������8�u�o��yPF�p�W�:U�c$ү��m����S{���1�����׺������U�P�⦉p.�$C�|�f�	��h���ǘ�����^��-?.3͸W��ݒ�,R��L
z�(}�Y�οj���<�H�hV��D��Mo��zg����C>�,jX�=��>�)�r�2֥!�����W�7E��w�^�,����<<�s>���=���-�;ٮ�{�y�R��k]�f-�׌�8My���.V�ӄ���r�|dF���»�OO;��+�����=���Pɲgrў�;���^:�D���	��j�3�{R�ꗷ\w��@G3��V�g�|X0�)Ϸ-��]��qU�j}���7N֏E�'��h�W"��彅e3P�H�^��#-�V+��s��q;��ʹAl��lx�i؛[��F^oɑo]؅���*]9�yn��^9�fA���K�K�����~���۞�'T�"�A�@��rͱu&���1E̥t��Bg��C�P`X�/o��ʪ���,�ޕ6�)_��(v��=5Y�x�7�>\���ߴ+�p���dh]"�hl�&I�Q�>�UK]��!k�L=��}�	���J�h`��m�}з��Z��<C� ���>&���ʪf`�"�W[ecC��JG��hZ���ed����8�9�p�F,2.Y�����,�.,���3�a��LC����+�V{M�ձvΧٽ��k}�l��9�7�w"���&I��/�hp{��p�J��,9��&罧Sgϻ��R__�𩙤7*ϏOL�9�*Zxl�K>��u���Y��9�ʯfq�Kt�/	�Z��Wp�5��k��P�&D�6��_O{U��<�J����QR���L:;}�"����o�+"�˶�C�����]��*Oi��X��a4}�fY�׳�[S���*��X��U��c1P�7��_���,gzH^�0���`~��h���L.�-ďY�M���%��N{`�7XO�{w"��z+;mb� b�B�^�&�����;x��M���
ө~qq�یA;̯nI��'�V�u�r�;׆^�mW�/d=��x�!�G�q��N��XI����$�sB���:va�GoƷ[���:��z�G�$f��<���
�޼���WA��v�b���45��O�͸s��^]
���}]�����(QR�z�e\�
�Jy��Oo1�F}�<]��	�}p�2fEa�L=y�Ξ0=�~��&�=��:��2�a��}�߲�SP��p8/�p�����6|^�h�IcuxXk��E��^��p�*�1�������ޣ�,���U�E���D��32��^>�z���WL�8��;dE~m���s����{�d5e���(ZO:�P��~�Y/���vC�K�����;����MR�u��o!w.�.�ޛ^���U���U\f_L%^;��{H�VzQ�C�9=xؿ�o�֧��X�OW8�z)bܙQ���Q䌞�II;v]�uR$vXG�U��(Wz��K:r^�}҉�ow�|�F��Ӎ>R���YE$����f[�/���~���u���}7�]�}t���Y�ӭ�Y��9��S�L�e�.�"� �P�<�Ȥ�I;�Č���p��U�<�6��Oe�~�cH��~��/9_�3v&Y0��iJ�V�6����L��C��r����B*��7ֺ)𿛀g�\��S�[x�BV¶頋Wix���(:TMj�CA�:�b�bgUv��[c-p	gѤĴ��pmgc6���.m�f����b���x���b�X�9��@���L�� e�$"<�*"��Z����]ڵq�q�f�z����s�0�v�,��|qM��=�}ӕ��Y��1wp�YK���!z+qr�6�Nb=Ŵp@����q��)�o�K��B����Y���%�o!�P�݉%���u�wy6���Q̮E�C�o(��tf���;#�.���XT��(X�EE�0�1&h,gU�+=�p���t{�< ���(���5@v�����vCj��A��V�\%�w~����@^��`��vuKC�0��s-/�b���5|�iLc	u�j�Φ����hMd7t�پ��p�#]�<�β����\�N��1�W��{x�Boo$;<[�'��6���w;�-�;#wlu,���v�3܍̃��`:��� �v�n�z��\|��y8c��E�]��9�g�|#2�7Z��=�>�0m�K��t�� S��IRjW��6�
�v�B�U� v�A$E�R)��<J���������ǲ�z�=��Sff���E�E�{�;���J�^��R"%{�$��4�ӓ��6��J��v�:�^-�q�*9j;�w��r3�I�W#cA�m�e_g�yļ���KO��������<��/(�Bl����{T�7�ߵ)�ܥ*��,���:tף�~f"����m�$3	���.�/n<]�ݤ�w�D���ə��alJ]@G�����cs�����@��0�
S��{�v����P�W*��t�N#1!�w��a���٥�
��wSJ���`Y�!WC+�����)�<�j�!�l�7��vU�As3����R<s�)aL�ʰ*�R��r�Pn��i�f�.�s�)AƑO^sO��p�]#���_݌H�ث=�]BjyX�\��8l\�Y,�u݆�wj���t��j
�l�S)�MLR�����G5X޹�Ӯa���*	�
8/���ǋ��	t�f`K�(I� �����z��e�
$�*6�
�(�V��Q�6dW�����u���'R�EU��I��\����뵦��̣v�t;�
����D�R�ceY+1�gV�!�}�CȎ$���������/ng�	��QM)�:�E�-�܀^ �
&U�մ8�z-��]�Y��Z�Eg�[���ێƅ��n����6{�vҵN��oI^��X6Y�/T�8���)I9��4kl������sk��̙��)S�9;4��V�5z�.�Ox��������3��/T��э������5�������V* �AIRKhUE*��E���E�QUEPQQ��Tb��-(|�r��V"��**�,Ģ��
,UTb#`��WTE�4�V5��.YEƠ��(��� �`�D�
1���EEAER(,�ej-�"����b�F�`�1Qd���d�F,YeV
ذk�,[h�Q%J��!X*��Q"��U���DEB����m*��FC��(�ALV���X�R((��`�
��¥�X#%aPQTr�jPq�EX�EYQ�Q�X咪)Y\���h�#��.R��֬�%�>J!(�������V8ۻ�h��g��z�w9�qޝ�)�d�=&#�f�*�N�.�fu&i&J�s�,�q�$���(.W8*������7<t��?�u�Bj�C\[ZO)q��J����/S�Z��W�΋�<���s<��7�IJ��y$�
�l�P�x�/�s��`A��=01��o��,���;�w(����Ы�r�7�u�J��Du����I�|i�!��1a�s�q�H��+9{�:�ו��9���`�r���<���y޵��1w\���=�!��;�u�dl��;K�,ޭ0E����a4Ќ]��K��=mh���-;嘘�t�E���V���B�P�����n�����������oc�s�<�������7������������Bɽ.}U<�Ȇ}�ق�i��rǢ�R���[Jo��̆��c-3%C{�8{]!O]��J����p�\~~�]�s�ȃ+l8�S���r�l�F�'�-Z�!엘����|�g���XD5P�k�V��\�@V�^����M����{�2\��>��3�z��p�~Zġ�ϯ��+-E`�"�Gԟ�V�H0Uh2��*T.���Q�E���z�*�(����;H����L���cU��K m��1�+�*�8/g�(/�Ŝ!L99�O�<�5o��'�N�Q+DO��-v���_7�����ϩ)��|��rSKv�o%y}���u��T}�R�w�1\�1Z�?��R%��H���@�b���KP����|�O��k�p�gx%<�uL����N���Q+��f�c�cZ��N����6�L�zĻG�Ey9�9�k>���=3��=�ġ�6/���s����ˉ2s�G���g�q�=V��	�&���$<���ϲ�C�J#eC��`mu���o&��]�ּM�a��ֶ<��R�7���y�\������X�V�S7��@���Q$��m���+��1�ZDT���?Z7��:e�b�pP���؅��E-\�A������u�pk��GOb�MP��ݞC��y7�� kL�������]����4�ty�e��Fk���q�����֮�<GE��d��ʯ.ō1��e"�:��ʶ�p'�{�!�H�s��]���hM����sE���[�y[¡����Du�foL��� 4o��`�pSԹC�G8����K����#̫�/�dWmWbC�u�kz����̮�3��ƥ���V̉�nt-��'�mὅ�k�V�v(�B�wP�m����g8��	�_M����=���i�ꗔq�B�Np"�L���ډ`�)Q����k����Y�˰2����`�)���7��v���z�Ph�׏�Y;H#c�,=SQa݄��,���ԥ.˙���������e��0����(��*�T����S_C�XC1�r�� �\Y�|�W��@�S�٘oݓ�嵞�)a����~�O+��	Vp>#�neDW��6�/&�>��b3r�����}��(d�3�h�X2u����/�U#����$S�w����9c!/���ƹy�ݰf1P�#ܤI�[3>w3��P�!�K�^��2�ц�f�,x��p��޴�`�ˬ�\A�y�4�t�z�S禡�+ř|ߴ�]r��~Ьd����?N��V� ߦý���~��f&i��U-<�q�l�����Ҋo�a0�ئ�K��KW�3ܔ7t|�Όx�W>�b<]��M �2,��f�vE.����G��O��oN�1u��uS�?zB��p�,��Ȱ%�aݠw�,x�.,2�s�3��O!ٙ�~B*7���=�V{S,�c�<o�d��xԙ$<why(�����P�d�b��Wx1��_w(3_��������~/�34�-�ç�zfqȥ!@�àA�കc��ᶵ�zQh7SaF\݃�&T�X�Bx�!����&x��6]h�'b�|��b�m�6=�X<�Ӎ�f��cm;"��s��Exm	~��l��n��>���P�hE���=����w���R��?e���
��R��d1�I���V�MVڧf�5�l�ǖg�Uר���n�-��.ǝ�N)ȴ':�J̅�*��5�{�P�̲a��v��긷��	�:���D�K�#ܺ�]�f�}�"��u�F	+"�[��K�*,1��{�F��v���#cD��t~�R>���(:�u���s%buB)�t*n�&^y�z=�w��mZ�K�M̻��X���F1]{i|R=f�7⯝	sG���ֻ�U�y�2dݼ�Ġ�,U��8r�օ�;L�OF;���`�����_D ���xo�9�+�<|�����uo��\$����+�������R��vZڹm���څ�gVwI�J��;j��`��������x�H�0�3�v��~���^mO4�{��z�@*�Y��j��b�*�:9j,��N��<a�'5�#\�t�P<���=��{7<��cG����*��fUBҿ���`c 6�J(�|���vC��/�T"�� �s.��j�47�u±�I��Ѵ|z}I`|bKG�=� ���؈���	fיr��!=+r��E����bU���$���s2�X����W��ot�w���ƈ�xO<J�Փ��b���� ��Ҽb�Z�nՍ�h����Q�CoW)��vL��k6�=����H���u]���|��2b�H��Ώ(��������t��ܙ�1룈[u��sN3A�`hu��u�'T-����o�r�<��^t�o�2��7bj��D���q��΄k	Ɵ,�hqDi��$����:t�3�}ںe��x�/�Q�����G��Ɍ���~Vns�6�;W2��.�"NHn�\�"ߠ��Q:ݵ��G3jT�eF��N߻G���	V4�G�qђ^r�Jf�g;�1�z�i}�C�I�0z�@��$>օ��lW��-'���߄��A�B��x�9<=�iR��+5�}���*�iJM+��u+��W���~�e���Qvc5�^��|&�`�:�z������"���]��\/�I^�#��墓X�=0d<�u^C4��o���?a�㏪��5a��|�^��7��t8�uR���}��ӨF\��{�K�o�,����BύD�t�S�d�Br'�Wt��=�bgzז�b�3�l�����ܗ�;)l���Ƈޱ�x^ױA�C�_�����3��XW����5����Y���k�ڽL7fP��z�i��v_Oh�}���^W����9�9�2���\j�r.}1 N�d,d��^:��'�;�E��ܡ�yʫ�wǳ���Z�1�W���D�v-�z�xQ�+���t�ܫ���Z-�b>�9ɏ/`��e�Wję�ޫȆ|��>��A����Zs��W�Z��<X��XҖ;����=���vJ=�^�gRܹp��b�6��`�aūݦ�R�iM�c3r�s;w��8��y�v����+�}P�k���qr�\} ��!�I�x��-�t�n�^Ԉ���\\�V'5-��!�Y�㱹Yj+#H��R����<|!�#�\v�l��=��@�b��{Jq'�d������yi��Q�j�*�Mp}�^{�zOT6��}�VÜ��8��.�.:K���w�ڜ�A��{f��;��De�-������r�nA7�0-���:�"p�7k�aXC��?Z}8�Y��-G<o���|5�ӷ���E�}�"k�)Dl�a���k����lK�;�V��]�����6�<�!��;P���:ռͼ�iD�*��e'�]t�Yg�-�i�f���h���X�{iq����^�5�C�18"��邇?��$���K\�9ʦ�7ϣi��Ѣ�yY�&��K���P��VMՠ�[�_c4�k�>Y�}�l���#�Mޕ�-f�ܗ�H�\��Yl)%<u|��|�q�g�^���Z=�p��*�:�m����R�t;w�@|+T�1_���1�''S��m�٧O-e)7��Mq��{�n����*鞟v�zP4�,�;�ZHP��y*��$[�ꐏ]W�O�.��[=r�Z�׹|�yY�-a�0�U�K�?"D8ê!�U�Ϻ����/8���S����4��i��xQ��+������b�=� ��.��/������Kc>��������W�!dS�x���δ�MoY�������R��յ�c۫�e�5�}��c�ԧ/:�C�d��>T�ҩ(.J+���c��߇��7��[ڝ{�Qf��oN�Ӟ��u��W�0���n��;[Y��������x��l��=��p�rda_<��^�/��Dz�*����2������Z���i�wYx�Ȗ��I�����v�������
��}�Ķ����1�;q׼��W���:�;�4���A�b�H5d�F�G�r�����KC�Pŕ�̰���K��Ƽv��w�'ꚋ;���f�U�����eB��ڙJ�u�XG��I�e����|E9��255�0�-DO���:�/����զ�K��I.���
B�Yr�;�ݷ��f�Zmϑ7$b�p�x��"��d�qK�x�^��B񈑋)S��)�5+��5�%�/�Ś;�G{B�������u�3(�5�������h�2K���>4;p	���vk����7�+��>T�ϻ.ȫ��(3mO%��gq�͒tE�s���OЪ����"QC�ݠkz�b�\\YA3,g9�ʄ��B��=�a��v�k5�.���x����r/Z��d����MrQ+����ȕ���N]�*������t��Ԝ�p�k�\�Ꙛpܬ:}�����T�`�!��->�=��t]�a�k�W��R�]yv�{�Rq1:�B��ҳ!b*�OE�1C��l� ��u3�JyIF$����X�5;�w����d�~��Y��`FEq�]�a�u<�Iį{ZF�f��c�r��U���:�#Ώ�
G�E�B��|������&��(�޺��5�H�}�Ȩ��(���>;2�������
�][�w8K�����l%�o.?Q��~���Ü�g��K#��_�lj�>�f��i啞��K7��x/C<�h�h�6!��Z'��w^���O;�P�v�D|:����	�}p�/'���q�/&4:b�}��x0�����ր��J�eZ]K}���
�=v���Y�{}���f�yS��9�a�^�'w�(۾R�O�ox�]��=���;k<�)r��˾p�R��Le�fئ�y��5�LVn�/���R�H���wͷ/_98׈><����;�:��O�|4c=B;���z�zUuCg�������ְ�#6m���YW3oO59�c���ؖ񒗝aq1��v��9���32��^>�/P���z?�.�s�y5�3��W
�8�X�
f�i�3>��S ������R�,��/dΗ��,^�W�|*�{^�g������vb�ޛ�z�OV�k*����J�w	&��xB]$�D�ںo�Q�*}ҌV�L�E\�|���IG���L��~��=��}�h<��)�I��͛{1-�6�fsH��bj��Dз��߀t#Xg�t�C��Di'�`�iWOpݶ=!�)�|���B[��\z��o�ܹ�/T#8l�������'<�Jv�L�g��~8�T蚞� �2�[����"�p4|�:oՇ�fߝ�NV�󊇈�G�qܒ󕱢��3�o�w~�s�/3�2���"N|G� �{�د���yK����%^j]ɛ�ײ��b���7���LZ=*70T6&F���J���u+!�����~�e���*"��]��V�y�2wA��w}���޳(�4�S��y�ۚ(^�,]���x�'�A��䃕�hm5J܃H;Ҡw��7�z��UE٦i3{2筎c��]���]�|�E�� ��|26g,g� ��7tz�q�n^尷|�OxqT��v��rJV�1�z���8�@J��HvT��)2\9E&��+�ص9|�pX�t�Ň��J�qCV�N�;�
�O���7]6ٳ�mY۬G�tz�,���^Q^�q�^�������Y�-�Y5��h�z�'9C����Op�:�0��s�s��Z��L���y[��k�G�We+��뀣oc�p�'�9�r/:Ss�ݗ(���U�ؘw�"�c��W�j����Uq���i��nX�X\�ӻ���>��^p�{�������޹�'���,�7��.K���U�;��L�!{���P�l��}�z<��q��i/���>�_@�{L�7^�,���V���u@7��:�ʌy�}��7o<��"�H�L����^	楽]�P�y`�v7+-Edi����˻t���]��So��9Hx��zjD�zY#�������ƣX&T3*�gMvǍ	<p��C�恛�ԁ0�Kn��Ǌ�i�a�f��L��ƵG>���z3M�D3ުJ)���d�(�[� ��4N�&̡��1S(�!��u�Zx�K93=r���s����Zq��.Y���ī�1�>����8�1�r��~���S���7��M�)Y�͠�St4	�y�d��s��6{n<b���]�\/,.]�І.�]�21� vEZ�R�"�.�hn�x���f����'S��F&��F�+@T_nGP��,/%
��[�J!.�}�,���$[z�&H�	�7�R�m�=��v���b��)�2�vSH��
�[��E|��u��! b,dT'|�=8�t�kz�K��q�j�]�r�aY�}]Y�^����(ax�]7ș�4�O���8R_ѽNMI�V��t�g=��)Y9(�aX-R�r�*V�Ԩ�� #ל�Yح^�c����]B��b�G.�F��Fw-Ita�E\�9�t����Q��w���#�o)��ז^���>7���W�ʃ����f���k;Rh?�^��s۬:���B�Vr�*2l!�z;�RZ�]Z���:�T}�����Z���k�KM	O�e_*L�r�jj�n�+L ��6n���Y�ݘ�9Vv�7w�NQuZδK����7|��v����o�&�񋼏Iٰ�vmL2���X��e�4t��T�СUڸX 4͵(��
�n��5Ӓf��,���k�fY���n@D��q�n����;�����ɹL�;�Mjʝ�.�erً��kx��a�3��� �}��u�]o����x,b�W2]�IwW4�wY�̠��]F�OV�S��X������()�C5e2๓�̇8`�z�PfE��R �W4
]�����D"��
!|%<���0C��:)��8���-ӷ`d7����i�L�;�����NTÂrw��Ծ��֫��u�T��b����t���" SZ�o�7ݶ���Yʹ��CN��j�P�n���̓]X���I�����ˬ덈�/@�`)�m�]s�5R�G/h$�$'>l᛺�-$��t��-1*����}���3fj�^գn�(�\)en�y���{8�'��|��m�a�v�TY�G9��n�R�c�dP��#(�z����`�;Y+7	�Qi@r 4a�Z�ǻ��j�+�t&�+u�F��#�����x�4��q�d��y���[�;�C�ۊ,�&�u(�O�c�����B���d/�b��laݎk���F�0����V�]N�ү,�o���2"����`̾o*�t������qFm��+=��X��t�*�0w�ׇ,bm�y`>����Bí�ۃ�2�1��b�O�)Q�3 �ՙ�Ԭn�;ɹ�XE6e�OJ�H��J�F�>ͽM�T��'Ǻ@K��!�.�5��� �!��}2v�ɇ���������
g����QDT����,1
�DX�#IPD���Q@R*�V�+	S-��Dk
��X+�Vbf$Z��DQ*QX�b*�őm��,��VX1���2�,U#PU�lEc�(�X��"��,Qb��X��d�������U�,b��ʪ�Z���[jDPYXU����$�Qb(��"1EF.$��"�ZY����EX�U
�1(���A1b�TQ,\lDZ�%eAc�DE���bTU��2�#DV ��e�EF �*,�TUEQF"�Q��P�UDZ�(��( �,\���)h�VR��T��S)T��*,�Z�E��Z؋[�lUb��;���߾���r4<��a�3�y��,t]O�4��gy�ׄ���7�Gnx[��(�Ect���ȳyٰ�Y;z��p�?6Z5H��v���Ơ6>K�v�Ձ{ق���.+ə���QF��J7����ؽkb��-�E=\�7U���n�Q҈�L�h!���A�w<�K�o�5�	n����o��˝&�Q3�ھL��%��o2� q�Q$��o�U�+��Yg\���,��5t8�u+�K�2/
�z_�Pߖ*bp���J��ђ{�M�^��\��zi��J1����E;�Q��c�W=��u��9yp�v�xJ�����A����4����j�g�����Kw���+{^�!�t^Vn�E[�ay�m��OQ��>�}&�Mz�G�ZF�a4:�
~[�]C��܈?�w��F��`n�R/�'� ���^j�4��Y^=ah�\�jǞ%�v�Vh�c��&�b�s�0i5�g���tfB(�^��`mg,粛v��n��o�т�ng%��pë�Ż^ ���%�Ep�V`f�ۙ��篙+���v1�?+�<�h;k�I���cK>��k�O-;w3�X`.��ߧ���5��h�T@�n�]���/���Tͮ��b�h$�}��K�QT��U��W��71��'L���!���Ofӝ�XT�g/s��\�Z�����Hݿnv��l�K��t_o�:� Y�����0���Lh�wM�O\������aw3c�8��'_���,��~�]���.�`�2�	�grў�:�X���#S�T��E�EzH&�>^�:-#ʾ���h�X8�8�n[3��C�{�}~�3Գ�ϕ��w4s�{s��$A��=2��i�U����)_q,zj���f:��u,{W�1Yg3�/�?-��߫a�X;���g�
�j"��+`��.i�oiE7�0�a(߆������~`�{���j�M�8�ޗh��������EUp���#��p��dy^�}ֶ���4/,�>�-��%���f�E�f����[ԋW
	��\�A����7~ηg`�w��^���L�q�ܩZ`��M;��(�����$k+�q�{���+K��iL�m�5�}��~/�34�ŹXt����=��j��C<�-Sљ,���m�D�rH�]uP�{�RqxN�и�⻅���2(oQp���f�����z��u'm���I�}H����pu�{=��s�`F䬈3[�^X/��ͻ��{j`*�Ս]�hm��%���_S(���P�x�̕x���o;�
/B-��Ӌ�,\S��q,X1�yqV�;W|	:�� <��GIk�,R�T��1+����5gX�N.m��;W1Ǳ1�	���9��Э��2�@W�%s���[��z:�~F6c�P�̻0�~4����UI��ce3`�6��w_E����1�R�o"+_�J�ז�%1֑W�y�QkVp�U
��<~��tXګ�6����Jlh:{P���ز��޶z.=jޗ�`nbm��W�Լ)��6���^]<���c�Y�bD�>���[�|0R>������(tgm�G��8>�N�}p�.���aWƲ�/���6�f�%�Ş����7�J\��>0h�z�w����:�ώ|�<G=%�Ֆ<+:��F.���z�^���8z��c�-񒥍X�B=�.�89j,��fS���+щǃ��",^Q��טw>�#��g�YP��՗�[jeT-+΂Ōb�ߩE�@�o����;�o|�L�1�����w(�͟7\+a�GǢXI-���1C8Z�6�]�v��X�<�g�Ԍ�g������U�?͇�SC�U��K�0mmB��1߉˗Z-�[�Ӫe����=�5ۉޡ<�.��3~t#XpN4�K(v�#M�����zy��~Z��GĤja�7q7�+-�3G׵���=�T��:��z
6���e��7�v�
�BR$[7��\;ԚD���NU��j�%E�~�0e0z'�����̢��*m ��/ޥ�V�!<<3�v��q��8�K~[�u�k��ImjK���Q��\��+n�l��N��g�'<�})�ɹ^�:�E�xw5ʩ]R@x�%�C����3o��'+ly�C�G#�����f�fA*����/3�+��ܺ&L4M}%"O�_y
U���~I�.9����f�UK�Ǻ�o�����Ճ�LZ=��x��P�)��J���u+2��7�򘏶J���|�Y�iMXz`~2�iϤ�k� t���/K�R/�E�P��BI���I�u�J�k���ZÛ��+.(i˶����S��˰�)bg�4���^���&
/��o}cA��҇��u�RX��[����	��h�s��89C��"e��{�Wy����8=�^L�U{T�RǷ>{��f�XȫVZ����/]�Q{9���Vv�!�uy�n�B}�+�݈|-B��+I��z�"��>��J{�|5*��r'ɣ�/R���zb�Wɾ�
W����U�FE����O�o�'��Q��K�o�1�O�I�-��S0���s�'|�v^����/@%�x�wXzjd_1q��wg������kk2F��3ۣ�`{ �*�*��mw��"�y��.�\4���N�QvZ�W��x�csP �E��'��_j�g�{H�M�,��F�̌V�沤�.'�滅������a���t���u���y�i�����w�V�|�d�F}3���<��v��*�Cw��QX#H���q,�w���q�;��!�|���kh[�]�N��K��(t��x��-/���ʆ�WA�vH�iL�?F�^���x��>"R�P�[r�4�Jޚ�o�a2�X|2�{�y�Y�B�yOz�El*E�6�P{)�v�
��K��#���{0Vu�z����2$/x�y�A�K�7+���.��V��f�엻U�A�a٢cJ#♆�C���փϝ���W��w��A!N]o�������M�b8�֮(E�},u�a3�R�t�WT�k>���B�Z��W[ئ�J��P�'��תe�~*��*br)gy	ۯ?7$0Z랹2S��3�r~��-q�l�:���=�>i��%��ĪgzP4����ܞft�f��GY�}���q����{���@��~˾��׹}�t^V}�-:��ʶ��২������yu��5�@���,�.,2��c�EJD���U��-�A�9�[C��	T�!Q���Gi���9�V}��.����>Z"}����
Y��+E䮷�+�G�oe�A+���׎�����Ӱ��x1�z�r[/Y��g+E�:׾�˩{H��=�Ygs֙L�͹��Du�f}�0R{p;�g��e��c6>�ՠ��%%C��0�6�՘�nu�9�)9����usݚ�y�];�{/e���|��ݝ\������`d��0�,[���~2���jИ},n�}������=u�P��[ܥ^|��l�5vNǶ���a����=.��yw�� ��Aۓ��&j�Pe�i�-7�W}��ϥݑ����Pɲgr�^>߃����ڥ��t`��Z>���*�)B.��<�뫀���'Ϸ-���a�P�!��{���gK�jDO��@��߼�c=��a�k>����C�����Y�zj���f[�����V�M��pP\��v������+�p�Q����Ғ�})8����<�KC�QM�V�Tkvԕ��7g��'�"�%W40N4;rf#�ó\l-�ѰWI���dWr���S�-�o=�zQy淊�Ü���ѱ��K^���Y���hk�@��"��W������i~�F+��2*�J����h�L�0��0�>cP�3IY��Ƚ�t�1�󺾷[��ɂ��T;�f��t�CluUZŇ���_k'sb�f��;R���Z�*�3�s�mr�-Q�0�K�е]���P$z	�R�o||ɿ.ݯ!F��Z4��/`�m�Z�����@�/S~=zq���W����Ԡ��^P�2��Ҙ&�#Z�X{<�p�a��=38�K[��߻��2�0cԁ�@����X���v�{�Rq9�Z�߾����ʸ����=3
j�����B�:�/����2�f͒CiqYI�U����ݒ-Q�0wL�=��Y�kV{ɮ�{��>=w���
�DP�}���a�~�H���X�j*m^��La���^�
Jr�S�|r�Z��p�&]À?R��H�Vg��:,-[Qۢ���뵕a�y�gO�q���б;��=�oL�����}h��k7�fJa��v.�Kz��/+q3~��5�m�G���'���H����/�&�w�=�iz��!qJ�;po�x�x�G0���$������+�j8`c�v�:���櫬����=�;�S
z��C��Lt���)C�����l�9��^�1{|�3\�Y�c]2�����P�I�<a��q�ܫy�0��]�z�J>2�9�7x��^L@hi�[k7ELʸ^��]�"�Mbc�c�v3�CH4�\I
B��1�{���j����dcKc�S�Ly�N�:�$>�z\T��O����u�|u�/<I�w��B�`��±5���u�>K�KÉ��B�B{����z�}K�+X�J�sV%��|�\�����]�Fث7�שD�Ui��������w��b��n�޽�%Lw	6m#!Y�F+�:��W4�#6,6��U��������]�%�d�#���S;-��X܉�vؚ��&���7��F���>Y0����>,����{���`KR�l%ܻ(Wg[�G˚��B3�Lg=:ߕ�d�6_=É����vy㏗�̤}aݠEC�k�B�E��g~~w9=��5��V4��W��ZH#�L>�ӷ���L�:^r�)���L70�5%"O�_y
U��|_�ZO(�~ʈ*��ݱ�\��d�K��,W�_ek���G���L����)4�UB9�}�<[�	E�/�����/���ǎ`���OL�]�9%+^�=N��Wt��L��3�}^����wz"/H��z�XwxwYk}�.��↭�:������O����m4�ݩݶ��gY����e���|ɓz��Nm<SdO^�5X3"�+�XJ� �Y���zx]�Íj�'��|�{
������u��#mv����[i~v�Yϧ��������*�w���� U���g�dݕ���'�x�K�ުr��k}EͶ��M*)FQ����6=����ִ�X;����	��h�s��:���%h�z�O�`'6���;��=�[��xQ���|+VZ��z�����ֽ��Q�;�{�'3űtHhUv+�Z���ʎz��v�ʦzgޫȆ|��>���X�Ll&��vt�v��`���3q���
W��7r�X���d�uv�=)+�.K��p�v��zTch՝���՗=�vp3�ȃm�}Nfx'Փ]��h�m�J0W�R�`^5�^����\����YS/p��#��I�L�w/�Rޮ�(C��ݏ`��-]v��RmѥyFl����ԝ�ʭ=c(0j�S�zjD��K��N�<����ƣQ�I�-G�sm�ک�U[�],B�44��4P�׹
8Yio�MC7�f,d��˕��zŮ��a�����x�f�X&R=r�6����i�Do+�f
ι�ʹ:��ǽh�Y�a��9?'ȧ��2k�{�HJ|�m]qя�@*�:Q(C_���mO����iE����@�MMΤ.��n�o��r?[i|]ϝ���s�H�}�x6f�[�}��j�l�Ż���#��%�:%B(l�ժ�_vweF��|q]ڤ�灷ۏvʽ���zqL<��
���p�P�3�W9\��%��'��#���tj�1�_���nG���T#+%��<�l<�iD�T�k8M's��E~��������ܬ~h~����?���2���C~Y�19�, ���G�����Wۥ@�{�W�=*�֎%)�x.����ar���2�D����e�=�B����dq
�ٝ��ݣ�e!�s2�B���.33뽊�m{�g��y[���:��ʶ��Y{בk��]�r5c^#��#M�C���[�]3���ǻ��G\Fg��+ ��du�#�#�Mnǒ����^_����S԰uC��Di4�g�yJL��5�f���S��X��yC+}�*lv5,��{-��ŝX:��csn�V���3�9�<~�>VT���U�z�0dy�f�]�}��E��X�{1����q�7�먳�Z�n�م��=��r���Y��#:�'�-6����vX��d{ �q�2l�?��t�ӛ�m��}[�1�#�l��=�)2�8VO��+��*��Pn[3����=��T]֓C3lNƱe��g�:�퀄37YQ�0e��*�-Og.���Z䢞ʋ�s�D��j�a;�2�GOQ�����I��m�6/���xo,��,�#-�� ����c%C���Ѵv�k��'�*ݽ$�(WDfCV9�����6�屔��K����U�
���z�3.yص�3	���?�=��0��f�qmG��|+��n��坑OGɖf'�2˭�߯7ǜ�Gz�
�JN�Y���K�ㆌ�=J���w���su��z��̍�c�z+��Q�Z��k���	�Le�À1���i+���Q�T��wY�srк�c�2���h��ZJ�F��;u���RAG7���9Y4xEbCѓZ�{v�%�so�]b���	�Q�ȇC�[�!�n��ql�jQ2Ş�l�-#P�n����}�7�zÜ�����{�9���V��ks��]^��Yy�o-$�vٜ��$�f}�7	ʆH7].}��%�Y.�@����V�ط�S��wAE�u�9x�-�v���De� B8R�����٠������uYʜ1�˥��\���Ѽ�TL̈́QB���lTQ�^c�A{��xJ�{���ŔH��o
�_eN��B�o����K������X\RFe�.���e����:#�X�v�u;[��^9|��\��%[#y��AS�n�x̒5�x+ݖ�����B�AИvb"��ͧ�|��2.��s�����2"��ow��Y�"��x��,�+��n�q�!���6u�:���W1N�ҢT�`<HlE}��Z���r5�bA��\�z���>6���W���Ԧm9oP�`kԋZ޵��`)�Ӥæ���qC9�a\	�ru/֏Z�*����0�s��h"S`m��	��StWQ�I��;� �	�N�7�������	���ǣ2et�����t@c)��wz9�	Y�;�{��{�ۏ�Q��t��N	n��mt5+@FP�Ź/ag(�P��'TWr�d��[x8��w}���o17��8� ��n���Zp�6�����=v*�����X1n4��k�n�9�����&\��,�u�)ݶ�c1���(�=k�B2��wء�hQC�j��ށ�*z& ��ı�A#��x�F�p	��\}�r�������'E�F������썎��->�h������k��_�X�eљٕ�g3��Z�=���y�`j��IwLP��A%TN��V������z�&�H��ײ��\�C���W���w��uC������k��$�;.���c���L:��"��+`��,a���l]n��E:���/���H1�V��F���@���R�T�c�j��ːM7)U�3j}��Y\�_���L�h�;rwAa7[�ԭI^��=㹰�Kڎ0ɪ�=�7���z,�號b��AX����VZUq�+L�b��Q��DAE�P@UUAEIkj"
[*�(ȃ��Ub0c"��AkLB�WQE�̪��1Q�FEkYPQ��b"(�mEU��U��X��(�`�Z1DE��$UQD`�1R���D�(�**�����U�hR*("#QDq0mR�Lh���-�EDEAFбD�m-�U���"���Q��(؈��V���X���*���""R�"�Qb���iD�[E��
�(�*QdU��b�-�[@�Q���U��b�2��q,�,UG)DX�(��3+s%cR"�,@PQ�P�\ikQTDb� �(�1�
��j��`�ڕm��`�����������X�m��e��Z"cH�R�DLJcQT[J��TE���b[bʶ�f"��b�
U,QDˆQKs
9jFb\��&Ya�`�}���Tg�cb�uk�:z�heMb�#�KsiP��4���{���n	��������'Ǳ���PH�u��ǹ�����C�ڲ_�e�̀¨�R��Z�ZxW�\8��1`�,�;*뙙-l����Y:�U�Kڙ�Rǵ{�����WH���P�#�IY���pB�n�,���l���es��e��58����z]���[I���m�j)�H䧗7�W��TEJ�V�"����h�u)p0�,Ϝ6��Cmݣ[ԋV����멳J[�p�Ӽ����3����W+~�uǆ���t�����#m*��;��7~!cю�T�����`�.6�2�L��iL�p�k��e9�p�a��fq�yv_���y�{ϑ�>�@e��`�.ʦz�z�]��E�q��J�^�S9���۳�a������5�`�ؙd���$w%�e.�^�,�ݽr/GG�щ5�y-�6 +P�������t��5�]�9�тT;beم�H���R�)^�dUϭ{������ޮ='\9��$�V�38�� u�uP���K�gQ#5f���鵶r< �НOD;ٕj��3�rk%��t�z�;װ����J��7g4D�����:oǙ��H;N�C���mX��3�_��vnU�x>Y0��ݍm�x��*Ʀ� �q�ǔ�X=�گ�ł]�1e2����)};!�n��<}]�f}�����Z�zQ/`�Q���Z9NW�P�-�]��n�14�>�!���R���e&�D��[1�D}�<e�L&�jC�]�J�D���Q��s��-���V)�c�;�h�Ӥn̔��%i�1��_��޻�����j�5�E�_{G_��dz��Uvg�`_k����(v�%��/:��'\Fh��w���8���fb��~.�c��W��^����&^���b��C}�����mD�'����n���w�*�>F�g����ԢkBVˇ:��-ߔhoe�dm՛�{U�ڍ�8�o��;v���G�3�a�,���ټt�/�
�J1_�N�g�T�`�lnA�iP�.F����s^|Кݿ1�����`�\^_L�Y�wr$ru	垔M��f��B5��Z`�z�oy�:���4xd�QIԠ$�'«����⣀;�5xJۄ{�&�]�zޑ�T��|�������z^�@��-e�葧T���'yD�°�f���W���.�lt���_]�oݛ�"�R˘b��h@�w��Oo{(�y�#�5}�5��uy�z�/��T6�Uk�ǅ\�&����6�=Z;R}㐒{�Ǵ��)ǝ���e�hn��M:��5Vε�Q՞��WMZ�����]�����|��-�ʹ֜}�(��y�[�9_�����&QJ �=����lW��C�ު�r�E����6���U���z��*b�J�����P��H��Ri%��G�����8){w�%�4�-�����gˋ0ܙ01*���J׆:U��ͼ������mU�]yΧg�Z�b�
u�U�[b������f,=ҒA��:�(��m��:����3^*�M�&em����r�_hn��I�L�Z@���W�$�U��M_΄h�_m�OzmQ�]b}�e2Lk���b`�^Zg���6�?R�xQnm^"<����b��������%�2vr�j����rs�~�!ږ}��Ya��hʅ�گj���� ���<�/_{�;�Wlz{���g6�N���M��ig��m��<t��
j��ҙ�*��q��a1���a�η|�쭭fz]�96�`���ϩ����f��wj����XC8|��ͿV�[�}��%�����P
�Ҭe����P��k��;���5-���P���C�yطx�Ѡ�'笍���O
���ҳq�����W�ʐ)��i�`d�e3"�:�W�����v®�j��:U��g ;�ɬ(���8e��s͝/�Yz�yl4�v�y^��s��,�6�)\�e�>��V]�pf�R�5�9�����v󩹎�m��>ի��Er�)z��������N$p=5<�}=��!]�yW�e�i��Nu`��WE�"p����\�
�u�*���ro-+MC7�l�g]VM�򖧪߉�;�4'�]�Q��?�R=K�x�
N��"7��{3g\�j���ah�lWu�����K�6�"B�Nx(�]ޯ��GO��D�t� �s��������u�s�����Cߺ�gj�%�GOP��y�^%B2����2� q�Q/o�V�a^yeZFF��z8���H���U��u	�1ݳ�L�,�X�Rг"��`��mJ+�=��g%�s،�H�WR�w���w�;4�E���~]��P��r٩_T}IN�>9��F�wo������I�[�hg��^���m{�g��yY�Dơ����eG�fol����~}ډ���Q��5�
�� 
�����k�9o�5*�3eű��*g���+|ǔ�0>�{y~�m�0�Â���hVh����K<���Za3�c�Ĺ'kWo!r�,�=n�M���+;�kK;�s���OjJ�(o���:��dь��yp_.�<�Q��*�U�$�ׄ箞��X^�ꒋ7�b~v1�ݮ�	U�ʝPMY�<�gvn�wǅǖ���LL��9�pλʹ@9��wv���e���q�����Rzgb6K�>��[ٌ�^,�θt��B,��&�̅@�Ţ�#jM,�Þ�i��)�M���C/�����E��Y_<�aJ�q�E���x��ڢ��XM�s���������:�`��}8K8m��_�������r�`�2�|&�d���{��]�zW��v�N�,=�)2�l+<K�J�OCP�G���u.��q8n�]�51wE=~���]����a�U>�CV֞_	P�zj�g����nl�n��;l鹗r&|�cڽ:�u�3�Yh��3*�˥CH^b�~��X7�ߑ�ot�4��=\��z�S���58�%W42q��.Ɲ�6��F�+��n��ޙVp�����_xع���*�m�+jj��h�u)p0�,��E�46ûE��+��8��Y��X�#�/�y�0�uA�eLZ�<oy�w)�����\��僦�
��h��*$z]����CaJe�)�ަ���G�A.��
�u���W{�)��	1<E��s/��.�4�,�n0-��������n1%��v��w@_Y2�e���b��k�൵+�.j�b���>$�_}��6G8�,�oCnu&�%��y��;��vWI���j@�����ōn$����]>ћ���W*4u_w�].��
�z���"М�wv��j�OJ�ֿ/m�������ˏ����ؙd���$/��iV>��K�����ȼE�`}f�r]����K{���齁���g>��:"���˳�H��mWԸ�^o���kӺ:�W��7#�/-u��̕��;���邒�*N]�u�-kP��˸q���	z{�={o ���7�$^(E������מ0��P��d���9CA9^kR�)��;�ނ܀�j���$̫���8�I��+P�)�J�xz���uo�ojD�:���r���]Ӹ9��{&c����<���Ƞ�<�~�__�����FK�2�e݌L�����X��dz�����1�$8m^��D���V]D�9��д����.�㬞~c�Mv�G/3��/VMw��m�lv���mL����}=B�P���4k��V�b�C���QE�qXw.��[��
47��#F^Sk�c/��|].�I�f�:�^"���n�%��y1��%���z��>%���z�\�%��ȿ���b�r�I��yK`a5�h�g6�˨Q�w��kؼ�s����Y5�3K:֝g�3�Y���r�=��k��1��}�_�tx���D�ǲK���3=|~��j^$d*J1	:���;>�lFװT�sٙ�v�r�(�a�d^�6�J%��N��+��}3g��D�	�'�}�Dо{�߃��<-[�xV��
p\u���8���hu����(��[ʮ.���T���7c�=�nC�_�0�9=����0f��7�N�̤ZHgH`��o(��,����M�ܗ�7,�Y��h:��Wl�cH����%MVĦn��&QJ#Om�C�,�)���z�Rۊa�t��>:\��J���2����L[�P񹂡�0�5���Uy[[��]��'y�'~ԡWݞ7xs��,��d��e�ӂJV�3�A�v��[�%��+�;��8 ��H�.�<�����&�����VqCa˶(��kxa�T�� �_vk�{T̻���uR���i3T�����5��W�'�Xޞ7y�G�cG�/w�� �E�躓D�ޭ$؊[ʱ3�k�KKL�3��W�nm
�^"<*�ب�m���y������a���q0D�J��1ߞVe�:q]���e�VhX���:�勝ۨ*7Xre)}�\�%���t�F����%��M⮖�r9xѾ��r幒6ﶄ{b]�#̏r�oj��]�%�O��6,�]��:,�ۆC�+��������}pl=o�g�Գ��u�eE��-�"\<�9�^)���Һ�'s�U��7�L�����>Ŧ��m,�m���������Q9I_� n��>�ܚ���r�� �]z�`�]�q�2 [A���`��q3s�}q�E=�{u֨��LZ6�������-mD�z�-+r�y¤E�I�Jf�چ��ײ�r�iR����c�7Y;͚����P�ErGԢZe��vq#�u"X=/����C-��.��wGoٯV��f�X&T6��,/�#iuҡ���GF&ZW��P�f�,���_���s�&��u��|�נ�[����}2��h�PKHv#yX�����V�o�2��Rޚq�E:L��*��!8~#n��'�q���}f���h��u)(�6��w���˲N��~�#�TD�}�'��8zmG���=P��X�V򙷔��a�=og��v�i���������S�1�T�Ӏ5�c�19�R�XV��N�ɛ�Wbz(q.�+s=W���(q���Q����mɾ����,���@x�ܷ7���d׹�S�8>[-ݐ�9:�WƧY�d���<!�=��7�c�8�Pa#-���⦺U��5`c����s�G&�%�cx�o���ma2z��}X�h�{�?ď��E�������ar�"v.��z,������빽��Ż����,3`ϹB(PCke��Fk����2�뽊��u�����b���M�<==N�ăZ2l�x�Ǖy���U���4:������;g�D1��z ���l�=��������n@��x�A��R�p�.�]�3��DV�hu����tϵQI_o���_M9�dV�y>=��V{�jO��\�g>�ŝY���snd^��~�n�\"��=���+l�W��`�����34g]�l��
׳�pw<��6�c&\�;{�k�㧖j�yD������8g�\�|t�F��Ȏ�>r�g��2���zZ`�|%fi�K�W^�]���ͭ7��Qa�U�KH�\G����(X<�8�}�l��
�&�X2�����jǆ9C��%���ue��U�^�-:��z�K��}�jp��)N�s�~8�i��T�:�=�ӫ�p�g����ai�dI:EV
<k�Z%�(_Z�M��@�!����Jz6O�$s ��o���Y9Ji-�$�L��?d�T��jX,�oZ��sy�	v���g�����ɧ�}������O.�!9�KDP�*L���+��\2���e�woK6��5�黤{���q�=U;����-\�5Q8��Ե�e�C�Q���^�0�jjqzUsC�C��m�'Rd@Lb��:����z��>k&gpD��UC�6�ȫ���6���Z9J\a�Y��a�(��fb�f�[�r�_�;�z�b�e��2��y����տY�����������z���dC�0�Wnl��Z���69D�����B���iI�{��g��iv�0��:�U�>~�����^�|fl��~�ѠGW�@�q����&{{��"��&���T����7s��)������\|Pޣ�T;be�($��KJ�K���zY����ܘV�����-򓨵����� ��g ��:%yxc�ѱ�+�"*�uaĞҤ�n�s&��S��������ͽ邒��E[��r�[��:lL��V;��;���:�V��z���"�U��p{vg�ߗ�oK&�Ab�,p7����NOY�ְn���v4Ǩ�w�3��,Qb���E�VQ+}��tc��j���-��`����B��哅�������ѩ܀��<Y�����C�Yz-gg�%"M��Y��Ad�`�z���UM��*'��Ss��Z�ujP�z\�s8����B��O�i2t�Yx���4k��!����{�w�~l�`���#�tOʌ���C輼]r�h��B��F��X¢�)��a�1"��fڠ��q0D���n�y�Ɩ��i���Mp��Us%�b^m�#�B��'W�nV��uN��]T��Z��~	�&`���)�`��w��]:����G�����d��a����!݃��ȡN����QN�+6�K��r'Jaͱ��8��c8�[��2[��L�*���s��d�(7ݮB�`�OmN��Ŧ#G��v`�9<����V��z�/8�ն��s ��zkٱ�=��<�X҄��5b�bѭ�m�}�q�x�F�f�DPFpB^����݅|�����ze[�2��V��z[7�#;���'���(Oq����|��*�ٮ{���(>��{$�ӫ��p��C�Z�*��%C�^���Pє���X<j�Ǭ�]�����1锻Aڜ�ww
ju��I!��S)�J��Õu�MS��.P��8��=n���RX�5�ѹ˃�u�6��w�R�2�=lV���̮�O?)�l�з���c�w# l�9E���;:�MH����;.0k�Z׋U��q,����5Wh�T�M8F{���x�G�s`�'q�N���Gݜz��FH��	BWBP��(�G���y��c=Wsc�L�]6��'����F-�¸{؆�Q�Q�vE�]��`���Z��s��Ɍ�B�1���KIl��`#��6nw�3N�#Y��jJ3��(1=���As��/�gL��D�.��d鏂#�6�������ʻK�(�G����铦��=	�f����~Y�w67��,M��&/hb�ڱ�G�w%��:���;�:��v�^j�iS;H�`�[<�2p��B��t��G+4�V^ծU�l��5E�����r��f�+�+W�S��w��ol:���X������C�-V��'�u٭.�Ӗ,�	��em�b� ������i#L}MW�7{X�܏��|.n\9�s3O��!��.j��s�+T���C��y��DA�ܬ8L��&����3���0a�`����I$~U��zxR��4��֥�2`޲����^i��&߫"4�vݬ:�p�B�u5]�b��m�>�$��V�	8Z�����=;A��K;�P. �E^di`��U��� ��^�t�	���tt`ٜ�ZC��af僴F.�e<��v��xX8�P��I{�V���:N�oS��z��t1�gX��3j�y;�d���ړH����E[y�j�_H;��(	�����o�'0�r�̞�	�w������Rӻ�jT_��$�nc�_sL�fdE�r�����,�"�QUQ���",V(��*"��mPA�K��*��L�� ��c2ʲ[E�ն�1e�-lQ�ƪ�ĤjUTX�DBխ[�q�U�����-��% �+l�ES3&H��G�B��Չ��
�PPYl��)�1�������ЪV��,m*(֌Rҫ-DEQF�V8�a�T�0¨�X�Jʪ
+1(�*QX�ª�(�Z�5(���"�j	2�ƱQJ�(�Y����*�DDb�#m�A�"Ĺ�(Y�*�W
Q�`�1G)F*r���"(8�c*"��q����d�-��m��������0q�EA�E��.f#�.P�"�9K-�[J
�"�X�S.G,�r�Ek*
��L32�֩�V�!s3�UE�& ��s�+�Kh�m��+�6� �k��cV"T+��R��������{�다����T��d^��+~�X�,����;�r<+wc�''�Rr��N_�YO�Md̝h�:�Zz!�ƸE����U��*��z�/����`H(iܪ�X�{�5�yw9����.?V���L��������,�V��uz)/םYu�վ��:|��l��=�mp,��ϯm��S�����z�k�F�^X��|;MYq,g�gz�#��T{u�{4f��e �B�(@{�5}P���)O�F��Pdn��c��	Y�{��iݨ���)�[*��X*�����P��#!SҌVd�fB�����M�ǋ�Ş1m�p����T�P�T*�&�6����٦��H�Bbȉ_=�lv��ϫݭ���䞘jK�����՘;�`u�c(U�TN�9���Z9�}
����=tD�N��0l"u�����>��މ�w�s��%;V&R4R�!�N��
.��d�]�S²��n��������/�l�Ҭi�~���%�W�L��2Ɇ��DЈ�P#Oo��wT�VzT;����o.��cm[�Z\-<e��߾�y�?(^�Tž��*�@�����+n �dØ|r򞜉�p�׫4U��b=��
/��(�&�1��%����"����x��w�:�D��hy�+]��YBƩ�uu����5�~��H ��{5`��<㷋x�2�v��}�*��<�軮x�jُ��żo�}s!]H��f} ˯�jΏ+k�0ܙ0?v4䔭xg*�!��N�����w���gXl�s��J�*���CU�D���e��-%e��.�3Z�v�e��.��,��߿d$X?���\˱�޴a��/ض�����^��&��@���=��wEl4 <�W���o�t����L��w�>��bC��}3�{+RP�
5Mͣ�����_y1	׾]�~7;+9y���ˀ��;FU�`A�8v�ˣ��5�'�ο?)M��3�gSf���uw^�h?u�fd�9^W���t+�v3:U�FE���8v�v�<y�0'<�ɭfQ��b�e�Ày��q�2 [A��S�����Φw�������eU�oi���0Ze�D��e.X��m/x�]�� uW)����~�oW=R���i�֮��̶Ύ4e_X�+-r��*+���4�����H�zjD�K��1��a�Y���/z���{�l�н�&T6���|Pg�K���{��be�&;7�2W�Z�s[C$���<A�~���.E��ns�b뫆�.Yy���������	��a��c��riy\�� 4�v���	4�hW+[g޾gK/����*�%�o+7�[�d���$����/�C��ྥ����ؽC���)�k�:��7�Sz���d�2Xք�OS�m`�H��v�(��a"7�Ӿ.�X�����{0�����|e�hz�����9ࣗ+����wH��DЎ�G3_Yۓ�f;����'G�Y���A��5=�|Y��h9���ϥ��a�3>��\i֍~���9�y�g��J�T-��^�c��<�;�c^2��b�*bJ��[�c��o6�6{qL�C׹h��H��P��w{�.[�Z<g�xo���õݷ/ݒ$�cw��o޼9 �
<�ȧb���i!:.�-ig�n+�\;��g4�u��/ڽ.xI]72ɩ���մN8)�'�5!ZdV���̦�d���q�����߱eI�ҥb��% ���D��T�=�h�C����������~��7'V��*�/0�5ޅ���,yL�k��ӫ�%�K�,U���8Y�ߺ��csn�W�ON"ǃ�|\V#�X܅p�6�����P��;�����������.�z,<]��7)���� 5����΀"2��ݯhe9��0�yk/y�5�6��Bb�����y����}喝N��U�>U8rw���1򷏪l{}�o#��2��N /:��+�\��!͒Q����+��ˎ��̶z�R�� �C��PK;�Aֻd�c���#�٘ǩ�&����t��z[�����������~5�ݺv������`�9J��A҄z�w-ͭ6�n�ϼ�+�)qa2,���e�&:���H�u�n�[��W�s��rz�a�}��g���X��t�-髋)m�a:���G�#ռԪ�����m��cq�&��,���/�w9C��X��Nw��)��Yh���PĶ�Z�f�vwMu��*ew�"T�aX�D��(��L&jrqzUsC �ny�6�F��݌�y�z���%���l_+D_$���TEA]m����j��-��%�[Y���D9]k��Y�p��z9�G�uR�u"���Ŕ39ݚ�v��^����<lc�<o%Om�GC|�(|�^Q�1s��sYj��$<�ݠk�(��Z	��M(�\*�����ؽ�Ei�X���י���9Xt�c��o�S�(��@��6j"��;>�K���~'|Dj�[v�n��='�>��<�ڻ��]L\|"���T;.�dQ$6��Ԝ]vG G|\:��gc��z�Y�"�W�*I�����MZ��Yv3�-��\�.�B8vq��㎞�{%�A<]׫��b��k��|�M�vnb'��k��������bgd3,	�fL������}_�_��'9z1��S�ޭ~�tVf��>���/�s6$��1*���՝*�&]�s��Hʈ�������ή���j�3����������X�})��y����a�:}���kSN��^��&etW�!�.�X�^ٔW�����_\����K���*�r�0������v9P.�=�e|ǧ����);���%^�*�����?Y�ɸ� �L���`=�P�\O���:�D��$�2��Ѧ𺬘��X��xϑ�2R�$�ʹoG�;l���1�EQ��s��-W��~/�l��c�pzm���k���
R�o�f/s�L	��������5����2�"��2��^>j�k�G�����*�TZ��xu�Y�p^S]�ɚ�C���S9\(_<;Ԛ�*�u.���-����Ƴcu²�5�v��ؘ�{���g��bq(�6N��} T�^ :�R2��J1X2u3<���;�(�sj����>:=��Q�$ʝ�C!q{���5��ȑ�P��zQ7]k]`�*��g�_�pM��8f=�#��X?-����Mߝ�����:����[��,z��o���a�5%q�
o�u�$Ҥ~��:#�~ޭ���p���:�pZu7$Ĳ�s{�(8]3xŨ��]��܀�����]��c�v
�*a7����G���������Kd*���a�8�rɆ�F�y&��)��qx/�⣁ܹ�foUas��D~�����,�s(�ɷ�Y�F�����j��C6hR���� oZ�[���[�kq�ݑ��t�v�o�u�=�J��XG�Y��%�+��ˢa�Q1�I4&�r.����#D3�9��X��w�c��3*���(_�*b����*�����{�{4�{�:�F�Z���u+��W��K�;-fŞ�>���]�9%+^+��^Eò���T�C1A�)�ܤ�t��Qq��پXv(����-%`��~�!s�؞Oa�{�?=�>ݢG�������޴�7�O-ʭ��f�5שbk:�W~!�*�����ߟ�k���X���	�tDۂ�&�Z�9���Z�3?o��)��Jxv_qØ+=�^V[�����n)�%C�k�
:ǈ��y=K:�=~�p���Uv�̓��~הͦ����q:�=���3����^����E���[&U��Uc�d�R��E1D2�Jvw}�K�h�,xJ:k���d$`.��3�@J�*��-�4r�#Zn;���Kj6Oo�0.^���ڒhW�ZO���籛��������\Y���2�3�wl!�?_7��_�8֞Ǿ�Vvs�T�C��YZcG�]Ԋ�f���q̓3w3�Q��+�"Z0�.\9��f@}{L��qpw3�����܅Oo��^�ϛ���7BWt������ ��ZV6�`.>�:�K�"|�ل�����^��,���d=��ߕn(A���ΰ�VZ���)���SK�(0hvq#��ʡv�	�y'��2{��WZ;����w����ʇ���!ai��ܓ�*2� (��m�7�n8�)z���p6%��?e䱭C�[��4ږ��K�x��M@o万�����drs�e<��#֩��T��%��3}�̉9�Qwes���GM�4K�PRĶ]�;�u�F|
�A2���A���MQ/�<���zק����Z�<���I/M߷KS��e�ܔI(cN�d^��:˱ݳ𩗧N,�w˭۾��	�W�k���0N��0P���7H���B�.����arx�=Eh8�'���y�r�W'5s�^3��;�J�"�JL-$)�\��u�^[�[���=���5��q��(�T:�n+�o#���g�~�h�~��V�km�i�Sc�<X4�=&��}ŵr�-<wQU��"%л�*�
�*u�����������t���WB�3xKR�Wj7�f\�0�	9�P�����*��[��T�	�QX�'/g����i�T�oZ3%a��m�
z��|�f�	���w�,���m�}ݶ
st{����So���r�S��J�rEg��6����uC��a�"��l>I�E�2�د�u5��qZ`��Y������Q���� �>��=���YՃ�6Eym���R��~��}B
�z%���^f�=����ؠ=�{w��D]d�+�zV���M��+��r�o^g��p����V�X��'	g�#���"�c��+��5�q��K��vFF�8�w���_���+{�6�+T.�E��VX+�������&��@7/��s0�KP�I{��q��pO���yV�g�l�����զ�b^��v��,�,�ws�>u6�
�;]�U�z�â��w��?j�^IwK0��i��k1zJ�"�w
��OR�.��a������UsC�C��g�6@�ɬ��^ON�Y�`R�"-���3>�"���l����M^�����hU}~�~�N��~�Fk:ex+L�5�pn�ݘ36Ur{(KF��{���P��:�Qj����[���^{V�[|���]i��P�]j�����.��/�{���H/|O�$lJ����ՆU�=t����:�O�ma3�[=���-�+Y\y�:�)�Ԛ�@�j]z��T��o�ԌW}A3/��k�~C>u�^3�t�Н��z�0���/k73m��^#�SD�@;��(����̱޶��&�#Z���Mܝ���DUW�|9��;$�6\u�O���㞔�Y�:�5��s]�)�Źx��쫗��V�{_�z��-���Y�{�����E�8%C��d�f�!7K��p��-߻\<��	�ˮ}v����y�-f���+"�]�^�՝C�uF6�wi�@��:7,���V8	*�#F#{�������<f邒qB)˾�E�n��w�l�Y�ӵH��^W�we�k�˺,mX�L���-����w�R\�X�}��>7�=WWt���<���ӫd;���^�E'rY�d��C��6�=�|2��_.�����I(,P�M����	ՙ�2�*3������<�:��h_
v����́�Gt�g�絖�yL�x`��3�u���,/=����^U-[�֥������2���K}����7@⧎��[�ֹX�WԵ����� ��f�N����͙��ӽ������Vq�¸g=�yv&���Օ�mߵ+�b��o�P��0�J���*��lb��;�n|]��X1]��C��7�\{]�hr��i\=�_�Dc��gd�����U��*�;�!�A�^�1:���P�X&��o�ח����8��z8:�Y\�;\�g(��UK]���J��y��Rj,�C����}�-���H����j���y7|�g�0��v%��g�U�e��lb�&ߩ
�J1	:�|3��~���l>�7<�g�b�k>6�v*��O��.T_R�//�a��D�}8ОPi��6��/_K�{ۭ�i0d���(F��Ӎw,�a�֨�4�$珈:;�����Rt����D/e宦�ﷱI[|G�'L�`d���n�۔�X�H�@��0I槆|O�s+�,��7��=�ϩ3�sS�}�_��cH��~����+Jf�e��0�9�oӽ�Cm]�1�ĥt��'�;�!BEy��L�|�o~�K�A���▽�.4;��OL�Y���4�HU�T���Z^��\;�x;y/���E��`~2�i��_n���-��F���wv���?)0S6�R$^/T�"�V�7��<vZÝ��G�<%��:�軒Q�B��T����	[~"��;MD8����A��2�����m佣C(8Z��}l� ,��'�Zz����+s&[��牺x�;�1LJ`ѡ�M�LVia
����R�zK��Ld�N�'^X=U+���`�aZj�9��+�9XVܫȖ+�d��.k��*��u� ���.�wm�'�hI��9��v�W�������^�:���3��4�����%�m@��V<u�_Tbof�ī�l:w|��0�m®vr*�.Z"�⚶]�����P�2�jc���urrh��P>��q�h��h���V2"@2Nb�J��n96���bw���H�U�!���ʻ�	�/��؋o
���c)&�!�J;.��;u�%�U��v6�]����B��-�5j���wh`�3��'T�]�U��h����M>�X� �x`η�Z}�Q�N�d.�5� �C�\b�e�GP�>Ej��+�w.��WI��e�B�EZ����`d
̑+��.8���,�:���c����c/V3�L�`�AC�pB�p�V��r�h�96�;�	�xyƋC-}%d��s����.zv�+܂��/�*�ছ����<���1�zn=Ӌ�wjHp�{8�F� �1�­}�x�S1��;{��I�38Ђ733d��5j.�Y00:�Ol��ַ������ỲV��}�U�Q���h^�=w{O�XĮ�(U՛.vB��;v�d�ҳD��`�rμr�x։I����/��BKc�vyC�j���<�����:���e��uQ�٢Ⱥr<�����M�}��!8a�r�����3�'�':��v�t��"�8d��=y�/���P�w6���*�����`�
�6�O�*�
N�!�۫7��r��+�0�/z�;�$���A�
1]�ܫᦀ�U!�v������<VB��/;]P�܇|�8Y%�Y�-�w�;��Y:�k�+�w�{�n�5�\��me�+%���h�[��ON{�+�Qt��J��V���(�9k�	O[Ԉ���2�6��X�l���v��8�T�ss^!�X2�bN��滿'�
���d>�~2�j3��ʗ�`o��,S�1X;һ'aX��N�k9�۵w�b\v�K��=t<��Ƶ�HA0M��z.���4=���"�Nܫb���u�r��������������!vN)��G��l"O<JW��1˻v���k#'�8�(!�b�=_w���W05wz�I�\k�w}I�ܻt�RW�/g�,�	í*3\7Y��OQͺ]�q�٧�"f)u^�V�S���t�Ǝ�ԧQ�g��9v���էv2���a=�7����+N�ѵwZrC̃6f�9�9�x�-nۺ��!o(�e�������r��S�K��2�4����(��2���'5�����<|+�T��r��-�bf��ַ�Ƨ-`��V-cQ�M���W�������̒�Ou�� ��I!�ְ�1ƴAJ2�U��XF�,�c��ư�[B�J�ʓ���T*9��#�k+���8���k��J-��PW.*f6���0VahZ�*(��0���,�&8��ª*�+i��),b"�2ʋ���kU�1ƦaAUb�,�ұb��*ʅs9eq�*J%J�¡Q�rҡF��cq�2�V+l�Z����E��T�A1J$PB���Ȧ0���A[aV�*��*TYPm
Z��+l��\J��jTr�R�����XDA\�Q�F�
�LeDD�ɌcS��*.4E*b���\d+EF"����(��L����TTr�Q�Kj(�
,dD�V�P�*ŋ��
�*���B�Z9�����
�Fe
��X.V�*+jV���!L��
�"���D@U���Q�5�V�<v��<KiVT�	\Ru�LRm�j�I�1�œb������\�X�t�{(.��V��_T�����������ߛ����z�A��<����̮Qh�U����*&k�R��u��R�Pc1ӗ��r�+�qy��:a5:�l8)�lr���L�^C�Ƈ��i:O\F�mo��V-���*��Bz;��n)�%C�X�pl=��[���~�}�+K���n��2��z�����B�^�ݯ[��A���8e��=L�ޕvr�kٝq��g���<�+ZfJM<��uf
�u+r���ِ}{L�3��,���N&�]{�^�_���V��{ڷ8M>���|`�
-tJǡ�T�J����"8�ل��m�3޷�,�M�|*I�/��Է��!�`��](��)�}J{��b�i�/���ʫ��^5u�V��2t��?k"ĩ�'��������2����M~�(l�RηNWr��ɲ*����F�J��5ݖL�Cܙ/k�@#4ږ��T��Zj��k(xu=<���ɾ#�Dv����Y�[Ɩ|wə�fx�uS�Ґ��v�P�{ё�/I]%�BR���o+�V���<:�<d
D�/;SQ���ӫ���g�O�w$.�4s��kÍ^p�Җϯi��G��\��,���[&��rLr�nHmz�]���l�s����#Y[Pb�N�`�1s�t��@�a<��z�칐%��mX������Ĺv��u �w2j����^:����<��}=P���sJ�;��~���ew���C�a��NR�]S1�#�^��О\ꙍ0*e�w=fK��U�f/3#o�˼���Yt��(;<�7J�����}qL�E�o�dRS��_ml~����Iy|_�.�0�^D�	o-$+�ٮJ�:�/�����u���az�8����8ϧQ�[���Yg�2��q�OQ!��!��&��v.Uո���ti�'Ϣ:�����6k�E�-�L�܊�-0o�=K�>4Qf@n꾸���&ۋU!v���gڰ{}p�fz-��!�(y.}����`Å�.;Ӧ��v��ӲK�z�S��J�Ex^f�$��}:���AcW�^S�僋�S/Yo��0=]1��/,w�2�<
��|���Ζ��Pw�,��e���iu���'�3
{ݥ����9����(dn�T�|��,�i\YK��	��_]\�lo�t~d�#g�..,�弸��it)X��{��'ͭ���*=�`(X�}%�s��Q����!ڜ�SJ��q������&�o���x+�Z��M��!��@�� _J�Ad�=N�Yr�\���[4Ӹ�u���[��{���s�)���%�v�E�F~�Kn���wå��zJ��_����C��`O�#�ו�ԡXWw�}���g&M\�}t��ρ�|:�8��1`�,�U9CΥ�j��z{��l�
�G�њ��08%�}�#'y�9G��k�R��X�bµ�D��(����a���惜hv���x���铩`.�s1�+x�N�F���Iq��e�b��+g"�����o��*��(Y���k�S)��<��C���wkU��X�W
	����hwa�u�\G���6�3ɟ$��m��.�W���B����!��������e���޶���)_���x3Sv�u��]i�k��8�Y��=38焧hP!�A6j%t���G���oc�PX�ϧ9�^��7���/	�Z��%fi�|]L\|"�����%�D����5�ŦtJ�sU��2�)=N�>�}��^r�Y�9��� ��|�!�:0	P�q�v�#Y�-P��x��X��]�E`�fR>E���?��Pu��2Vo�"]w��Y��z������7Ƨ�Jj�"n�M��j�s�g4��A�Hk��os�l#��	�j�t)�K%Z�]���%�t��
9z�f�rvV֧g�����' _n��`�onV6wʬ�k;a�/z�Z
�X]���Ѩǒd�T�ޛ�#=�z����)�$�3/����L�g ~��0u3U�Y��鞳�n|�Kz=e�n ۉƀ�?d�����m䝺�$��ȱ�%�r���Zw%�֑*�^C�WS�8��{��Er�M�!>%K9~��N� `���o�
�{p�,9�zW�/j����jE�R�2R�/�k��잌ꝿ��VW�k���5�����3�P��{�Ǧ��7�bդ8]^���d��H8��am���5b���l�E^�3)����z�	��������+X^�Z'{���ݎ�����qϒ�į.�(0{�5T!�a�̇ê[���~������R�o!w>�D��|lvҵ�M$��/�c�I���
Ͻ(�l�����`U�Q7�vM��J|��,�K��RQ�&
0���T^�U��K�Z܉�����v��D~��4��G�5N�M[{�o�Ѝa�Wj醇_ʈ�IrLKb��*�� M�Q��<����Q�ی����n�m�=��(�M��φF����jZG|�@��`�|�ʨ������ۢ@��}���s��֬-��S(Jݭ{J&��v����qs����N��tv��X���X�R�;Wyۮjy��y�7ѷ8b�u���;�_-�<;��Y����P�D�j�u����]��q��Y�w�_�������[؁v):�9	���sp������lK��%X�/�#���}�\�})���L(x��u����/q���o�t�/ihu�A�y��3㸧l׹P��+�_��]���DA�aS5��/_{�`��-�G��G�%µ�ߢ�/G;-fŞ�%���q!8��(f��۸�r�Q�}I�Ш�W1�A�<��%"���qb�پXv)ʃ���ӛ�<8;c:��=�{T`
����wlr����.�ϻ֒f�<�.X����g�<C^���9��/Lz��\`�LŃ�Z)��i�9Â�&�C�yV&w�y�uo�����<�L��_����Iyx�
)ͣ��#��P�V\���y=K>�W޿X�2��e�X�������RY�JJ?;ȇn�`��;P;���x��ў��291�]�	������t��3��wh�����2R\0���2�d�����s0{�7��{��]Z���9�s�\�W�
�P�k�%c�&���-�9�H���$�~���)k�7,
�iT/�ۇ���M�up���.�f.�F���0��|�"��uL�ʶ����B�p�;�W'E*a`�`�7Zl�c1eE���F�2�[�ߤk���Y�k�'t��pL�2�=i̎i�r;�������΁{��/u�%�������,�P�%��}qO\��Kz�"�^u������Mz������]E]C5v;�dik���/��o�֑~)�������'�������eC��rZh3`�����L�s��Eu\ݔ���d3�F�.1+zj�0�c%�j:����	��X�4@+.��k'��`�l�z��B�I�l��oCq3=�2$2s�G�Ww��
g�٬0�w��K����J�>3l�>�>qf�C��6������{1�A[镧��h�uq�P�ޫ�sf''��E���m���l;�iD�f4����a�<��f5T���[��*N�1���v�كS�5{�ꘅ��Z�0PvZ��ZWN�w��Uz��ᴒ��Y�b�^<��0���x���\/�v�e/�(E	b�?H
�n'C�\�w��ke�\�.�����h�ʯ)�D�t^V�h�V^V�9󂞣�}N��o���⏙՛&��y����~Έk󼉈鑙�0R��$Vp�LpSԹC�]����V.�Q�+vc��H�������L���+ϣ�x;�����v'	3��)�(tj�a���We�9��w�Vv.�MV�<k�a��ܴH'i�B���n��d,Ǥr�`�i��9���>I��,�u'����٘�W�5ǝ�9-�u��=x[v�^�5�nLY��EM��rY`��q7�=�h����@�=���9Ƕ�e��{Ǆ:�X�d��(AS��A~�W��`�ߒd����U��;�~Ey5jN�nͳw�;�Ls��ǧ��iz/5�w�զ�1�Mv���X��'	g�=��1���bo�vT�L�#7/��dn=�p*����~�)X�����
�*�I�y�ݥc{�ԽY�*�E"O��fc��w�t��l��V����7��W!{��w,�]_T�*\� ���^�֞U�wǦ��+K2�m�O�*�}��g|���
����x�����ڍ���^Um��J�`V�aj%�=�X=0�o�'��\ШUQ�,����͇�Zl�lib�{1�pTC8��G�e$�{ZB��}���<�l�q���	�G���eۄ�9�~�v�:[Y�q�ȿ��;���E����=�Sz@�*�i����FS��kn��>K=��t��<���z�ܖ������6S/(S0����"���v�:�|���YT��1{�r	������9�����Y���A�>KRd-��m��$ŉ1[��a �p�WZ��t�qs{���R�A}E�����R�guŔNhk�XV
�WO��ް;�=veGw{����`|��t��&�'9}Z�f�����*��W��q�du�O��g��X6t�Bl�K+<����T�#��v�%>[(W�M.�΢п�����=��b�衽G%C�2�d��J)z���aΏ�o�IT��R�]uA���r/|�����VD�OT�Q�k�:m�J��gO/h�-��e�B�+a#�R��̓����;�Ř7�
J�r�&=�6��т����=9���A�v��>�����֍�M@T�� �/���4�[��ו�����]�n�.+�>ݼ����X���W�Լ9NV77}g�X~C)1[��(�#��y�Im�=���ʷ��\`��ȏ�>�M[ۄ��S�[�گsl<G�.��mN�O+���u.�7�Ru��'f�ڑ^��������c�s�ln�}�}���e��tb�˵J�RW!�Zg��^k2�ƫʰȿ��� �:(2�٘;��Y��?���h;�J��x��b���sX������ı���.��ޤ�YP������<X��|*3����m\�n�*|��t��"4F��9� �Y�3Bj��V�2���m��T��z�ɷ֟{�K<1����bO�a�+�IH� ���c��<��n&�f.R�<V�ŷ��P:����R�e��6���i���zӨ/yS��u�?P�+67\+ɇ��g�RX�KG�=��:����5��z���u��ۛ��8��C���[�P��6�wT�M���1����} ^�5�����sUē�ռy� �V+��/e��{/c�Ó�w,�hqDiϒ�6��U1��#ղ�Ssǽ����aC�/Y�[p�xN�F�M��π��x߾��KH��M�����{�O��}z����Z��Xz�8����_`��V4�����>$��~���K4��$R+v���|�'L�4O�D�"օo*�
�5�ƽʇ��\����nl�h7�T|�l2t�X�dlٹ����FD�^L��d2��+��9�k0.,�Kzy��f�(o�!�>S{jz��ӿ0��')��)q�RpC��aN�9������<�;fXH���Q����yxϦ�I_�E�e��H�t<����_E���C�3��OQ���D��8���!l�W�Y����e�i�KE>�Mht#D�pS$���<���+��[N,��/jTe�V�l��[�)���á�)c�n�=�=���(�-I2��o0��-���X��қ*e����G[v*3ʹ�}wGNZ��wָ����1�ls0��wz�t��1����#��w'���Q�z[_tr�aL�>y���_������%t�P�1"�V�O!��������Sep���d^���j��4`{"&'䷪��;���c��fcc�L��Q,�k�D7z�C^]j
�hs{-��bp>ڈ�U�k=�o��t<t�V'���>>��a��a.??	W�'��D+l8��|�&�U���eXoR�5]��	�ұ=.�g���XC
-tJǡ��`.���>�	Z3�w��q6/k�.mS>$φ�qy.^���z!�U�	�VZ��E4��OW�XG��F�9J^�5݅-u�~��y���R%�J�P��~��w��N59d^R:j|l*�B+��>�Ms8�}�+�l�Mϯ��G--MC7e�.P�&g�u�Q��KH�K;�U��q�x=}=��$l�p$�;�":-�v/í� m���~>��meϷ�"�3˅���X�5�-�]�}�K�\dh|��Q|Wo���mu��s&�	U� ��L��Q��֢�U��R��&B1��_5ʱ�`ZkF������>�}��_zBH@��	!I��	!I��B���$��	!I��IO�!$ I?�B���IO�!$ I?���$��$�	'IJBH@�~!$ I��$��$�	'�BH@�bB����$��	!I�$�	'�$�	'����)���ZQ ����9,�������_���0K�}m�� 
J�(J(�(P7{�ATQUB����D@+�1T�RER�UU	*C�`oN�����4�3�P&e-��h]��Q�]�
uU�t4�p��۠�ʫe�*C@ (   ��n�͍�Գ��FƇ�f��[h�K[I�ZXl1���5�i���� �m2�2�.ڂCcL�h�M�f�!�!�.ڡY5VMkimM��c%.��mmdխ,��͐jF�cj��� ��]�-P�m��&�k( 8ݴ�,چ�CF�U�՛S��J �     ����R���4��  L��4�S�R���M20F�2F9�14L�2da0M4����E?�R        *HB	�2a'��S�z� i�7��5 �J%(��i�� � :�녹ߙ�X��S��T�*��r	"J��mt\��H����%���		�Ix�})�J����DH�4������ߟ��>��Y4���_������G2���EDM�H$�]Ci��wdA"O�D:�$h��5IPgH�!e$B$�R<c=<rf��dS�w�c���z�0}��	$�I(I$�$�}��>|���D�I�!'�	$�(B3��}��|�\�$�Ir�d��Gρ����(�?�#��Fh��K��iG¨�Zj�Q�W%��������f�]��<�1�y�;��N����܏-�%�����Hĕ�w@�uyض��"��+�5��?��AOH�ݡ���ev}��He_hC�l�
��k�cI$0h�5��C-R����*��AWY�1�cn��&˘�Z%��=t�J�D��5����<l��I!��S��KeF��I �:Y���.�KH���C��XFZȘb�V��vv]�t¤�W�h%��
�;�,�U�7a7u��v�\b6���f�;{%�M�N�!mwe�`�kBV;ru�v��tnŠ�V��R�X�y���wQ9*,%��H�t>�
i�3-��.9��5��l�ہ�j���Q�+rJն%[�.͕ �{vIHP�vK�m��&az,�
�b[B��+NdJ������+iP��1 �X0��(�YYx�Y�,��]�wDc�����:�]b���u(`�}a�l%�Vhӧ{���PZ/r�X�eڧ2XI�2F*⊎a&�1VSܧ�]�P���Yop@>���!�)�G�����da�X3���ʣj�Q��t���xm�����ѯq1U��je���~�l'Ȃ�B��Fs���/9�[Zm�X�k��)w׆�2��<�<�+^������qCx2��ƛ��L��FH��U�źI�n���VItr�f�bs~Mޣ8 ^4z���7�����h�&��b��k���mL�ѻ��0˄݀VF��R!��^<��酗��3[i�{oMt6�ܤ֫��v��-�������@��dU��ʍh@���o&�o�󬕐ځ�i��P���s���	��W!P�bf}3�sv�[���������� 5wj�PO��y[*E��$dr����Է��Z�&�_͕#pZON�+tf�X�.;��[XoL%Y�(]�j�̣�\�*nR��:�J3�~���H����u�v0a��.B⳦�Ź�?��ɲ�N����YF\�f��J���%4��m+-�X�3s����(�|l}�����Ɗ"ȡ.�2�+CF�*�5-m�լЪZ�i��B�[{2S����9�1��,uͫ)�;�M7ԏך
/R��Ŋ�3]�l�Q	��4�+u� 2��ۣvM�4� �Zc(iN��Pڎj���cU ���uwt^ަ��G+�����_]sy�m�T,���*�,����U�:�}��G�ܜ��c�oc,��e��*;�t�U�L3�<�92�H+1�2��(^�3��ʾ��EU���F鍥KlN)P�n��v֡�H4�(^�E�t���M�ܧ��W.�4C�5�-gڢ+S�to�u�V��ѻ���ݹtQ�B�עU���V��b�1b�j�S[Ǉn��v�7��Yy@c�+]�KI�kv����WU��H��iF��*e��4st/��r�fg�!�Mj��yx*[��4��(����,���9B8~�{���G5��i�w�
�$��A�TlVV}���¨^�ˣ}����XF�Qĵa'��H��h[�O�YE�g���6Z��1���_��3�W�oDWY�[�ٌ
8F��{sʔs]e���ws2�h͗������jP�j�Ć��.�Z��Uw��-�y��"��L�z�k� ���y��+��_z�/W�}�l��6��������I����p����l�Y�\Z*bvѷ��,/���6�}���ť|�Љt����F��l\hA��H��,����!c��nT�Kz�n�*�n�%��Q�77��%D�eqћ��x��ۛ6�]L�5�ݲV�62��;�B��`�l�NH�0�i�N������pYS����Ҟ"��ղS{5>�dI���m�Ƌֶ�F#%XSl, �{"\���&��0���懵x��w�G��$��HC���7&�j�Y���ޛ�&�c�lR��X� ��!��t�H�J�K���88ӹ�%�Cj�+������k"[�Qg>̜�ԇ�=<X��!׻%�{���U��<��TjW0�ܑ�C�WXa2L����ʢ�]Ӥ�6�l5w#cxZ�u����E��%K��]�f'���'Q����,KOn���p�sv� 8,p�	9N�\#Q5���-�ru�o�������Rwxm=���'#�!���31�B��`��Nq��\�����5��Bĥk'��q�ղ��]��KSv�(��*�J��rl6pm�����-����Du�q��D�N�ß��mwP]�m����n�&��W)�RfM/�����$O_tEf����C�����=g�� ���<��wu|.��lA��.��Gm-�[}�N·�� �.Z
ms�-e��y%K[���U:�a!X�ku���-�p� �����
��+e��ծf�o��*��F�n��kz	�#9r<ĵs�L�|\6֤!��;�\un��`�^�mMvj��f���.sV���'V5�@V[�N����u�0]>P��������gW	=$�ނIA�m��v쪃w4(E팽����+x��k����{�WG\��O_!#����t���b���l�:dg�,��W^>��rOiv�å��Z�z�E��8��唭]y�+�ٴx��c���aI�v�ig��|�i!\�ay2��e;�Y�`��ɹY��o)����e��
��.�3���sw&l�UT�7���4��]lθ�:5VS�ӵY�J�95�j���	j�9OE�},���p'�Dk	�t��f��9n�q_-�R]�F��è��p	EL�W8s�nW�Q�M�ho<����+�M�7�����n
B�t	��gG����zް�E3�r���L!о?k�gI��:MZ������q�*����v+�c������ã �i����Վ]oJMmv:m��u�K�b�ڱ���"�s,]���ه/1�j�h�V%9���`�I�%%v)��u��[ٺ{5&:Δ��ve>h���-�V�rM]��'%�+�#��bν��`�S�&�#Z�	-7>� 6ƚ�ɹ��(���NL@s3�;32�����d�e�8ڮ}{�R;�/��xT���ǒ��Sч���4|���Ԭ��N�y���,�B�{�z��*����.na;B�z�����u����[�Z��/�@s)>8+�I��I,��Y��ݪ�0k].�I0�w`�:L�Y�9dHwm7����q���p�mfle5+��5�@n&�[*)ϳGof����$����
��uj&T�39�n��V��s�L�it�k��.��M�0\po:k�ct��mr�T�#�Bc�ڵg�D5�PfXڹ�CW$A�b�RNׯӇ�<p��16�p�G���§ޒI{n�wҕ��-�j"$�i�3�܍�w�U��y��Y"Nè��v����ۿ�g�e������[�&�&��yw]�D�b�ڱi����gT�\�Uɇ�ȧ�d�x�p��.����z�գ�u>sLQ���NJS��<�H�@��*f,}�)g��"�-��4�ؖ��-���VL���d�Du
��I�(�y���}g0�[��fP����R�f�G
��㐚��4�ٺؐ�ۋ��F��@wR�3�%>*��ɰ:i<����5+4v�X�b�3yW-i;��!�\��I��GK��y�-9�wrk:m��e1v�]�}1� m�ھ�V�3�b����GF���1\T�C�4iEe2itD�]�W��d��hԿ�+7K9��y1β�jCo�طk?���z��>��g��R5��;+�7LU�MǘAhe�m-��Ԭs��`�nd�I
�&�:��]E�_8^l��:���/4Tʹe�`�����v���<���Й�]W�ħV���|˽����ā)a���ܝ$c-F5v�k�r�{6f�+wK6���9�*LN�wwi`M3�C���\�at1��fv�[�V�J��f4:��ڇ�D)� X���Ŕ�c�i���g*]q��:ˡ�Y�0��γ3)�tCW���H��v���'���VD�*v;��r�+�YH�kjE<��Eu�F�;FM;�2�䛷]*���6�ۘ�u�GaS���T��{�{��Օ���+'M��l�����a2�	�]�����3OM����F�[���bD�T^�C�|m�	hf�d��+���]�,!b-Pf��{A��ψtqs�v�K���V�FV�I)�$�<C��3)�k�n�U�r�a�~��y�ޚά��6�|��$N��$��+�@B
ő.��jU�70p�a.ղá�K/w<�)m��w:��b���K"ÏWp��
Tk�V:����\	W�D<��O�D�L��bf �4�V���-�����.�2�Hsǒ�F�X%Z.>W�H����5]`nR�(�2��o�5��7[��wҰ�e� �9ɾi$���Es���^�X�6Ӛ�y۝w7�ћE�4��ȷ�q��mJMd2�	�K̄��Y�a�h�/�o[vkm�f����np���Q�]$��jM9k�h7x�1�[z(��5��`ʻ/cTt3jQ�T���S�OHG��I��V��MƜ��'����r��L<�C�0��nr#*��.Y���M�6r��q˩jnY��V��KK���)����*0*�sX�z���H{͝��'��v��A۽��:�1ܬs�zcʛ�zn��[���-��޶�[l)0X������DՌ���}L��bk�X�;�_Q���Cjj(Ꮼ]8�L�l��u/�6����ʢb)��2�aVŸ��Κ���2��Y����h�,*q�,ۺKElK�Q�y�V
��PI,�(K���]���]QJĥ\#�'`z��/8�MN��m�g|Ӣ�`l�W.vGm,u�3���խ���R��d-Pl�Z�t
1V%��Tr�ʥ��F��Bj��k��M̽�:P�E�E%�\�3i��:Ʌc�6�-���Sz��C�!ٯ�E�l5��Mm�PE-h��>3��x���Ì���.Z�_�68T�� Y������<��g���i $$@AE���6�?�����p��(k�%�,��r9`�Q�o�d@�~�uU�T&���|1���b���1�jҳ���&�7��6S��#�T�r
��=j*:�Ys	��򷙺6��ďw���i�t;�)<�'\L=�,��jR��Ԣ{b��zE����-�6^ؤ��G�K�tU��R@k�����Q��h喧jJ���ʺC%�����1��W��{�+�[���ª��E'Z�R����(�*(���h��J�lP(�EUE����q�Q�.qf[V1�`���%h�*-b���Y�X��aS&,�,�D�.-Y��l��5o��׵�g�`��]w��smN|����L���W��_�/�]�}�r�f��ۦ�eN���
�7����^w3t�d�Z�|����U�,\�Q�{�LӗGӳ��|sn��ܹ����<'�[��Q�i7��>]0��<Ą�i����R�j�(i�w�GY������TY�R�."����g�wa�kݭxp�^�CG���LfF6OUC��0��B卆؉G��%�H����|�w1b)��A�'�Py}b���f�E�t}��<z�r�oӵ$�x�Y��K��S���X�|�̈́X���OcB���^lO����HcqlqP�ODŽ�E�1���/d*8�OO&kxV��86�.����5��:"BI~���!j����`���yj��2��8�˛���Wע\�v��8"��E���\����[��w/��(a���<׫�<�r���Y͸�kr"��@�{7�zvQ�u�P6mth���t0*� o�Җ��6��좦����u�����
�i+�\y�:כF��֌�ס3j;�ޓ;fU��{W��_�g�@���,���{����=��oS��\�s兹qIaQ%z���dK$~��{�s�iʳ�ݢ��bryތ���DY��S���|.��z�����͞�W_�e���͊a�.��Q����v�h�*ӎ3�ۂ�,ԙ��t�c�j��^m��x��:47=O�,~�k���� �|�Nu�ftm��]Z���]3쏆4
��=���`~��������ش��z��w��̂���C ���=��X�,����a*���e��失hsed�rc,�Qjf�󾵽�,0r���yP�$[����.�Z�է����2���*I)f���x<U�-��h �p��V�ʑM��Ț�V�]�G,�E��̄E�3}��BK�+�b�]�,��t�aU�ϳ�u���b�D�+|�ЅV
�[��fU�Ki���>p��S��.�>Ϲs�}����i�*�n�^�V:	5�z"�N�_6dg#�r=3�W�{�YuY}u�k{��d��R���*e�+�(Ú��ES©_��(W��v�꺬�g��t���{��O:gR��s������ǌޮ�ݦ���֌��X�Z..pWi���f��8ƾ�_"���M�8t�s�w�\��L5<�8�1�?}��w<��ӎ7t��f^���`�r�A;L&�2��Ω��{��&s�ZM�QOD�:�0_�t���aOen�"l�"+���uN�wח^��w�m��v^ł �S�S��UOZ�|H�X4R�T��(��}��Q'|�{��*���Z��S{�w;�f�<�ՙC�9��.<��Sf�gg��|�:v�#�q�{�V٤*������R2��uc�F,�&�\f���&_{����5�E;l��O�i���'��Xާo��( E�aҼj	��^�������e�����i���u�V�>������jmۇ{�|�(0�R�g\�^��M8gڦY�(��ǖ㻹CI�Y�/�zʓI3���a6߬ƨ{�Ǌsx��Mvͦ�y�L��<ʜg�͔����<?x0������U�Θ���|�gY�8�	�>޴=}�n��c4����=��M���G=a�`�)�ä�fS;5�k�ъ,�y0nϰk��'�j :���߿h�����_���> x��nI��;��ϳ�� `n�;�i�47/nQ�51|��啛��XGb�����)RR��Om-����(XLQ�����`M<����wq���i��S�h���bۖA�еՁ���ں�ݽ�x.7'�O2v�P�99��6��b��w+��6k->=C����g�\�ph�iY�R�ѳ����5��z'��#ѹ��ve��ZGq1�HѮ�Z��6�/���^P��_
�/�CR���.Q��}� 7U�9C>Ckm	�m����Ŧ�ycss\u#SQ�����q�F�@V����G9�[`�7P�x+�:rKe�-{��\�&죻��vJW��K�o��e�uqkw���ρgl��O������V ���p��X�UZ0\[�
�B�YX�T���*�!QT�IYm!�\%+XW�"C	D�e[����*EEVKe�kFIpЬQ.)qEU���P�5ߖ���P26�΋��~�F�����*���SܡWx��j2�dŵ/��W.�g���߽�G�ܧ=C��:ÌFW���5�~g�i�s��O3-���i��
�`�Ã���W�X�~�|�6�Bv�3�Ɇk�����.�x����͘x��ۃ|�ӛ�ځ��??��΋󛪛�~>w�����EK�ˮe'Y�oޯʝ7L�e�=C�3?}������~cފ�S,�e�����G�t-����S�yX�ڊ�96�Kz�����u�w/��/)g��}�~�kha��� ��:��|����gwHc�;�6�8�k��(#>k�K��tˬw�Z���A5N0/�i�{z��逸l��������kt�c42��s_�^�f��ݤ��^w����?3���j�����m��O]v�;L��)�bM�lQ-��������[�{K���Z/����<ix��|�q�FH
Y+���Ԣa���|��}�o\�56�Y�?3���8�~��q�)�N�ZAg��:���c0RZ+�5b�EX���kݿ;����e�Ӕ�f�=�^��l5Ȃ�Xjq�����9�$9�p�L�b�*�<����s�ot��;8l4�?}�{Z���|�nڤ��c�
�7�&3VJ�w8�&Ӭ�i�~�����q�����⇰��Z��}��)��/^D��h���꺃�M
��j�K��~�9f_��M�@�)���}Ĺw�m�V�]P�� ����N��Nd]��u[�S��T?���qݕ�<����7��?=����5�t�wɃT��1�N�o�{�P�|̸v����ɲ0>��V�@��EU�*q����q�'��Je����K�~�ƼϱN��6�8�f�L~M{�s�2��������l���P31�:�S~����[��Ci�m�C�~r�~�z�w~g�ًLr�vW)[�6Ͻq����+>e�.�z�M55��{>���0�,�i?g�On�~�~�M��kC,�T'	��c�7�U{k�(�>�(���r>�uy9Jo�L?�f��1���t�q�rn��ϯ�M�.���4O��x���3��p�)�{����>�>C�+��q�����;�}�ה��
1C�GQQf����z&��ҬȚob�2|~UW�C��}f�g��k�<�O����]�ߵ�cx���N��͡�m�r� �k�����i1�(�Z'�u3��8�6�ݙeL��?&ܱ�Ӊ�������C�1�/��\2�kڛfSo�\!�=�gﵹש�+�8�C�}NW�ǳ��P峯]R�H�]��{����y�콯�1L�3S�4��㊣�(��TI�a�/lM�` ���/���G��ڎ<�wq��Q¢���.T���y�́I��q۽ӻ��q����6��-�6`���4�4�񛏳`e�aS�3�����{8��6�<r�@��Խ��� ����*�"����gc��fb�<t��*T�s��~g���?c�L�I���/��M3W�<C�۷	�8̮y�]f�e|�8r�Ǳ+��9���2�1�p�����퓷4J�u*oA��O���nFRRH�UR�O�&���}�k���S��8��؛CL0+G��L����c��~~c��)��R)���l�k��8�v�}��w������|���>�ߟ'��f���VSx��ݸ͟��xkz�i��a��i��;��s�����=���dZ�_��>��)�6���S��?��q�,�.��b���L|����U���_�E����(3�rܸ������ew�	]6��Et�֯�u]u��o/��������o�T�P�^�HU��/r-�p��J�,�e�u���׹��o�<��6�<�c��{&~�:w��hi1��&��4G�*=�WLW�}<�xS�T���*e�?8fP�������c?��]��}�!F�?d?^z˖���©#��aI���c���u��������4�HUM5V���{F�/��˖�y�/_����Q܅�R��ۺ�cI�P�O�0���M��3��>O3��?8AC}��o�R~r��v������˯-Hw�F�w�^�e��YL��i2�:c8�������v����_���}�c�;�?'�{���rn��f3f�0z�z���\�/7;i��<�d�6�s�u��?'٧Y���2���?�xs�w�O�~r�%�u2�Bg�����5���u�}�̺�ܘ(�U�BW��
��%��̳�(Wj�d��;�̬t�+gG�r�\�������&R�핽�lHggb�Ѕu`d�v:��e:�٨�L��+�;�4�j�x"�{2�GmiՑs{+V�q�eT�8�T�U�)s>P=���W��KOt�o;Ђ���/����q"Gdu������Զ��^����Z$�a)������V�^�Ļj�]59�b؊��b�+v���a������-�}a��J2�eݺ�sfcy����v�J��QZ�ٵxTZ�wY��.l�l<�r��命s�w���]��{(9�+�]E�\�@7l,|��4)����9�k������?��oߒ�%E2���j�!�K.,*#
ª`(T�k�1�Eb0X�e�F�AÌ\4��0Uj(�DiI�b�%��,|������0������e�W�	Jɒ�.���=�`������/�6(�Oΐy����͜v�N��T<����^���a��Ì�{�wzv��M>e��!�c4�o�{d��)~�?Y������>|��~��4�ϓo�_sܡ��<��WN�P-���?���� �)����kY�y�H/�C	E ���R�� �� (���Ť�̦w6AI�k[�q��:��P������\���AC�+�� ���@�
��L3	 ���9�]�Ăÿ�0� T%a���8!��Ͱ����P2� ��
�R
A@QH)!ϰm��]�2:��t�:;7�Dc�F�G�e�Qܟh;/v�Y�������7ϴ�Xe�O��$<��Lڢ�RT�m ��%O���V�H)E  �}��:����P4�E��q�$��b�l+�Ry
�QH��X~aR&�ل��l*Adc�d�
) �i3�AH,+ؤ���RhJ�A`u��\z��0�i%H,��(
,ܜ�﹄��R
Aa� �����@� ��*Aa���� �(�q������{�I���� �`(
) �sVa ��
�L*ACi*Aa�TP�J�R<�R0����>�rq ��EiR
Ar���0�AH(J���Y4ʐR"ņXT���!�����|E ���R��i���}HT~d�'�)�Va�R�`m�a
�AI~�cS�Ă��R0� �JʐR� ��2�	��Xa �c�0)�
�R
u���_ך�l>a_�q$
�E ���R������H,<¤���0���9�w��T��0��ԕ �q��aR
AfFJ���R
AH)�a���{I�%d`G���=��κa�i�w�lA�47t<���+�=d�Ȼ��9��ݽ�=�[���$O'�$��aX��
�Rq
�R
C�R ���,*AH) ���w�ϫ��_vGԂ��Va�XjA`~k�H(~a�	 �C�	 ���R
AH)��:�gpP!�@�>I4�l��!� jH}��}��AH) �O�?��.P�i��q��f{M3Ns~q�&���ɮҌ+��>�7�o׹��:ΰ�T^���ɞ��ƽ�b���/��c��za�粀����}O3lÔ�/;��S�Xsr�I�쿯��������~�a�J˹1r�h_���F����];��-Mt��c9%�A8�Ci��f�f;��+6�|���*
��Ws����Cu�3%�Sȱ������߹+Y��<�x;d�d)y{ѽ�{=�3��J怲��39z]L�ey�]y��w��,�j/��w�zUR���R� ��黋���������	V_4�I��H~�#=�ݷ�u,Z� ���١�7��Fx֨��r�V{�v;Q��*ew��@я۩���d�
��v��OH�ڰ��8z.����\�RujjS���v�:���H�}��ȿ��{O����x��c��-�j�EN�_6dfk�j=��)�6�|R����;�.�oB�O�y�6v�k�)}�e��>��lݤU۩wR(�l���j���0�˭�{�N��E��N�d����Y�B4_����I^�_��tA�߉��!n,��B
4Nܨ�g�����'#��Ȋ�����f�J����y|ǟM�xT��4��⻃xʱ*.`X}����o -�u���^��ݺ��D��ز���&�j�P�Bʞ�� �"�"�_��GN9��u{��pq�|���g��k�)r��{��n;q9��ő��`隼�ܸ�{�h����v��<*�����B���T�t���D�t��������l�ٶ%r��-xN�]E�����g0G=ᏹ67Y��s�].�sGlӀE��yYY,��u�D���H�~��{T?�e+8���y��gs��f
���g^�t�4�<q�n�S��Q�}.>�a��T���E�Y�@Nm"�vҎ�g�+%�n7toG^����k{d�nW��]����uW���jc�<B\w�Ղ�Q\�?��|�k�o�	{�~���{8�}��Q#�ܾ���yaO��=��{�f��/�t��I�oj�V6�����.���^W�*�ڒ�k9��7�{��ޜ��T��}�g���Rc���h��%�5�:��.d��Z3T^rkF`�4t6�����O���dMg�_}f}x���&�u��-����W%sш���[�������::ּ��/O����Snc�fX�.�g�`�Wu���˘p+S��8͎S���0��fM��v��K%m	�l�Ȁ�������ߪ��ra�
��5r�'7a�]Fo��r>�9��:��)�jX;�RʛG��a515�nd�/�; k)ST���(��1ڗ��]f��7��7h��b��QjZCV��(ĭ��Ş�z._[�s3����Rv���E�.ۙg���t�0��s�I�V^����0E�6�#�����������L6�b����d�QQF1dcq�L4DX�X�R*ȵ
�m�qh��-k�\R�Q�E�jE%eE�(8j��J�Qc�o���:�����:���<0�?��Ԛ=��V�ͅ=��H[�z:����d��8��}[�I��8˄$��J�c�C�g����aҲ��{/}'�Q�wz������L�<h}^��w�mTx�����ĥ׼�B�ߨ��o������Q|�ќv����q�r�8����UT�?߿~��̙ں}�����q�� ��W����z:(X�&�*���}�.��)�49�W�#�'w�|BCٚ}�3�>��Ax{!#b�����g]nɑ��g=�^���
=��
M��9nV��ծbP�[Q܎O꯫�'?���z�"��sӆg���U�6ܠ����b.5�AL��:"���͘9mr�Z�%�=��u����m����;��j�.%���Z�7$�k��\\L+o��ؙ���ּ�Ta:�bP��
��Xr�M;�\M�z)?�����?b�훎������6�,��3�5+�_`�'�a��_j)h������Q���;�}� }C��A:�4�X�=� 1tou�#�yw��!��	�1���Kr�w�J� Ż�@�N`g����)]z��Zܟ�W��zH��z�{Nቸ�$��e��Gr�;�x�|�Y���w�(��+��������k]�P��j,99pOa@�6 �n6u<똩����v��6��nuA֢sՔݶ �z3M4!��ź�0$�T�*�nFn}_W�4�[��t%ފЮc���)����s��d^|���N��1���$��p&)ڹ�;W�;u��{0�M�˝\;K���|�6{�\��i[]}DR�A����
���ڧ̉�]��Ί��$w�;���w%s�ڏ����������ۂ{o?W*��Ӵ[>�V���2<b�a�Ǟ�c?
��Ph�׳�:�^+M��������(��_�\w[��MsG`Y���G���VR���Q�Iҩ�쵹��o\\Z�����B��y(Ye��C'�W��SM��~��uQ��~#�}�r���!w;�G���Ly���5��V�33S����FX��f9�X:=w\�>�G����\p5޿ ydc߇*�V+�v��Q�z�U��w�M��WJ����QI�U��U5��xx���M�ş�����њ��.��{V_#�I�����2/0)��vG<�<���3[7�V�t푘��=�7U�Fa��c�u]"�pXWK��xW��I_������N1Zi
}r�Q��qZ����+WI?��ꯩ�F~�{�c����޳�n�gY����\��sw}���z�1��Ƽ��=ko��>�h�[���-{U+�Q�k�/���q�0F��z�j=�y[$A^�᜞�@T�~���R���4j{]��Ώ᠅�m�%[$j�]��#ۅ[��	x�i��S���ʴm �.fSȨoy״�ύ��C�����y���bUN`�κcP�*e����Jˏr ����Ϡ��1�؉��a:��)<�+��Mgu�G��[*���B�����|��sQr瓮���0��GDf�7Rx;�(پ���"3�3J��mHIͫ 7�\�G����:Sr`��v���U��p����D�lJ�)&��y+����^��/:���p�8؍Ѿf�����'_54d6��
ǫ�+�:�Ycv��P�#��� +��db0Xe(�X�+E+DQ��V�R؃+X��T��k-�)[m��J1Qh�T��R«
�،�eJ�
2)-h"�P�X%�����h���u�T�d�ȱ�&�a�'�}��_}�<s��h�#�����㪠꼛
���F���g�H/����}j+�yK��{L,��d��*W^�]Ԫ���8U�	�f��Y���휬��d���a��x����1{t6{w��F���WRf�B����]9�h�#c�GȈ��?~)�m�^gtW��;0��F�
�r=B�X�o�n3�$��3L��W�U^{��%Wku\�i�^]�":�����������\*r�s<Y�37�]��=�r��4�^&v�==j_	F*.�=��%��|����%�n��އ~�~蝤Y'��	/v��!���\��{i�o��r�a��9�V��3�<|��`e��G3j�aKyy�Wk���#��x':�l�^)��;����\�����ªr���=�{�p���_Hcqkr}U�}\��@;�f?������D��7��;&����vQ��~����e�Z���H���ʳU:V9&��`b�V)�|:�Xr��ʓ7�3f�yt�@%`W�S1�ھ����_OwΪ�ø��i����a�j6{��ڛ��g%�>D|��rϲ_���;~���wˎ�����@+���nT�?�����)�1��q��b� �?=��jK�mm4���zOo]^�:���� �KC�#�{�;y9�qeNC�9Y�Bj9��N�˗
f��{�/Q�D�~��'JM˗1��a�'�_}_U4������{Bo��z���{�^��F�1�,�"���{YP}�*��Vҩ�o{��L��}!=Ɣ~ܿ�ې�>oz<U}�����E�;������e�n���fu���x~%!��J��2h�Nu�fB������+ﾪ������;���p��8���ˌ9�w�O���8�����n\����4o�>�n��6�1u�$��B�A{�	��A��:���3��oG��>���.=���|:��ߎ��S���+�~��8�=���N����2����I�W�}�4�n�k�����Y�&�J�{K�(�,��ͻ{c*j]S5Nʳ�{��G�K�[H�_Wg��:���{Z��fx�� jw��nYz��j�W�om�a��B�c�kӗ+���D�>g��y�{�V�`8�R�X���|ّ��I��UW�Q{��Y����_V�S�v�<qqKq~G&sH�T�/'OGv�n؞Z����xE�|7Svr_��\�a>��d�f(��5�N��D���K�/�%�T�(H�����m���[�3>?�[nv`F�8Wv���qs�#��Vc�(ʑ��U}_4�U�gg�ߙ����kǟ_Z>�Y�2��܂�g��'���]��������6�W�f%۩��>��i���s���R�"�u�/=�S�R��X}��o�~Rf/��yߡ7�w��dX.(nM��뺇I/��NfG9�halp7��1'�ucGJh;��� ��h���WM���*���4� c�h>��K2���GugWb�30٬�ɩϖS��68R eL��P��[Z�nu�J��I�=�側h�<�P�C����Hm8+��o���d�j��ȕA~�ȋ�8ｯ��x��rv�J3�n.L�+e��B�&���'P�gy�d��gJ�KN��R*�ii뻧�|���:vЎ��;z��u2T�f>�6�`K����ȕص�qɊQ��K��>�3�G0E�]�=���Nv���Yz����i5���9C��\��-��9�8��C����T-�2,b�KJ��j�R�h�mR�Z�҃ikj��Ѣ�ZT�Uk,����YR�,m�V�R�ՕQ+KJ�-��[Z�b��mb�Q(�F���Ԫ[milh��eb�T����=����s�N�}֗c��-�w#s����#�[��0�
��~J��}����6�s�̓ސ����^�
tJ�y��Q��/f+ژO��g��0/��`�4I��xoL9���@����%˝4���S�,��}�f-k���g����f��\��B����h�N}U�S%�k��b���vtwzO!�%۔�t�bl-{ػuթ��}��)�W�m��wq���7N���B��YJ�kf�T��9v^{�(��1� {�f3�:���[{��n݀k;z�o��'K��t�X|F;p��*;��i�����_}�6��&N��U����
X(��c/dY����OL����ެv%Pz�!��v��2GA�w�?s����G�.�%�}��[g��x��j	��U��Y�Ku�����J���B:���[��G'E��1	.�
�mH�F9�}�S�D��.���o@��q�c�ᚂ��?5�y�.��J�����囆Fm}���8T/.�l֑5�nrz5�=)n$�n���+XP���\��\�V^mJ��@t's�L F~Q��w�b�4a�e��(����8��ꪑ�?Eٟ��TwMh���&tgt��i�~[��x��7W��n,�9���a465���m	Jb�^��kZ��7p��i��gڼP������[3�ߣ�=N��>��^-���̦�G�o'�Ek�.�6����W�}E�mW�`�k�~��/*]u�Ϗ�/��_:h*�|��5��¥�dh�E6�dj�V�TE�{Z���g�@��3N���蟛X��f��y)���&�poO
9���{-��pH����U�ܸ��s���Q7���fDӓ�s��������NK��j&6��5�nÌ��*�T�Uc��ީJ�3+@�ƻu�O��=�y�����^qT�#�� �w ��v-�����y"pR�Ry��w"�d���M��[�a	�ic{H���6��ޣ"��	֥�=MM��Oꪪ���hl�{}~�����>��d�\E�<z����?�vW/�Q=�g�-S��_�����i��grR��������w���)A��{mBkw��?���թ�ԩ[�l���1T��.b|q�#)?�����i�� K��~�4��ٰj��+lQX&�����Co[�� �r=;����!�r������5���^���q����y��虗傭,�9�tc:�@}�$�v1��ў�����=ץ==��"P� �Z�%x�FWH�����d����}�c߇��x��[@P�n:Wr��Y@!±ՂU��w%�4���;�&�,�r)g i������޴"��l�������r�����Yt�ܽ���/��{u����q
xcũ�'��[��'<�a�l�sv��$�+��):N%��Kw�{���t�ܾۣ�LJl�l�0ӊ�k..��coUI� �ڙBf|ـ$�_D�7H=VލVŽ����P�T��-�(����Gn�_qΥr�3|9�@�>��J�^�VO[��n]WPU��gT��n��5��l�+GS�����!Q��\�6hg%n�ZV�RY���b�ِw�`+���5�KI���2df,9�,�!��h8&���	�m�&޽�
3�]r��e��1�wп�d�Ǩqf�rIjE�X�{S!t����+y��*Ǔ�g�NW�ݾ���&��h[�7Kc���VյiUAVKkj�ť���������AT�b�QR҉J4�(�Тڵ-�YF��Ѷ�
�e�"ҔB��5,T���m�Dj�`��-Km��[DD����le�j���F��E-(��lXڊ[kB��~���1�������Q���|ҕ!s������+����m�^���k�PNWۜ.��~�sUg���Z��3�i�u] �G�̑�����:��W6��L\p�n�0̩x��UR����<ɪ�P���[��9~13�8^+�ߥ�r	�0���p̔�w-��>|=�}�1�҂Sg�<��&���;Cל=iӗ'Wn�([w�;Y9���O�Z�G�;�.������r@gU~+W����gg�;��&�Ր�~���Ku�ݨk��SS�A/ҹ8�r���Y͸�kr�}I;�3-��z�z�e�HV�!S6`Ҥ6b�Ҿ�\��y#o��BCȢ���B����/��Z�dl��.}8���Y�a ��[�����YƇ�bC�j���u�(H��%c�	���U��&MFAG�1>8�����T�NB���u�_�C�r����}�-)�)vyr��o�����W��[7���K�{2&z!���>NU�`����΅�d*��t��Ԍ~���qU��c�A���+$6\��Ĝ�v1�:o���}�P�lj�D�������}�]a���m󅥸<��L�N�ѽ�맑:�WĜ����2��I=o{���;�-NM5k�[]�{����g��(^dVð{;3�2�e�n%�f=^�\9�G��)V��Z3V3q]9i�J���*$����5g�$������.��e����b�-^��蕡�H���.�� >�v�t�ݦ�c��Ş)�S�D�󻰮S;&ݧ�'�R��R�p}}]L!���X�e��6�֋��t������
t�j��#9s��jH�'����.0r?�}-j��.f�Z~��n����Z/=u�9+�^�/+8�V	�u,���y�U���y�t�ݓ6e����Ln�O���C������~]\����u' �15R���$$���m��En�n�
J�֗��ܾ>ڝ���<;ϭ�����h:�xL��-5Eկl�����Z1�b�]^4��n��,"c6Ϋ�<�&���y�7���uu�6C@*�{��o�e��§'��z:���-A�to1>��#������s�<G�[��K9Qg&��̥D��G6o�J�R�4�uҞ|��5����)�k7$<w30��0�{9O 	���v]������n1��Q W�j�|L��=��~�מ�;�c?'W�/���4ڝy�	�Sw:�#m��H�O޺�0s[�s|J������<�ۚ@Xr"a?n��'����6�pghIG|��Վ����]du�R�C��̠��;+.��J�TT8��,� չ��=��P#6���i�߰eLm����2��h��Gh�Y�MVC�����^��b����_ �ʘѽ�E-M]+��h�\�{���Z�vQ�	Y/ V�}�(���fd$��Ю�c  X������l��;�L��;����)Cx�-�I�|�_��&���|#�7(��y%A�;ȋؕ����󴌛��bh��Ҳ��T�3��7�<7�X�.��'�̞N��7�]���H(�r9�gL�%4����-�f��@��;��a�����|oh�+�tM��yp�d&��4��f.�]r@nW0"l�zv+�L��2�y�&����$�T�]�8�j�nE�0��hH]78h���|�k�v5U���h�镨:�IX���G��wTB�U�+A�lhڊR�h�X���k(��V�V�i[Qm��KZ�JUV������V�FЪ�V�X-VZѣm���5JX�eFƵmTleQQ�Q+j(����R�m�*Z[h�D�j�l�,S߯=~���_?;�����Vd�o��-��È����(�c�7�}�{�W˟~6��>����/�%��'�V^�K�5|��H��}ܜ>�~`g��p���re�]���Skn�]��<�l�L�4����6cg�k�Hr�֨B��h\L�=i
Ԕ,���țW��d�]�
啴x�[���`C89m�(-�0��v���Ì �	
�A��3��X9QU�Ҷ5ֽ���}=�`:H�����1bT�����/&�YjH+��ӱ� �B�]ժ��sj�[[�7��%�7яJ3Ǽm�ܽ&�jGh��V���k���s��cr�&�4�s�`>�>�!�2�d����?`&�V���hy�2wj3K9uԙ�2RJ�4En}��iܨFٻg�[�y�e�ٸ�!�j�s�
MBSk�	��ɗ�7����*xU�yǕj3���<.�6������gO{t��7�y1�gs��[Yq8.z�})_A��4{��ڪ�<A��<�y�%��{c9�̋�n��~yy�M�!�B���a� ���Ι�gX�ђ���|i�ld���-9��jc�����L9I��WT��i�1H�q���S
,z-����>�gYo5��77�猳��l��1jr�GL����\9��v�h#��J'u6�em�GпFӻ�wړ'�s$A{r�>�;3hK� �o�Y�ڜF7먭wTl�,�z��ש����n�ou���9��Gv�˵��b�"�s��=z���X Y�lv%�Š���ҳ"�V�f�E�߻�-u�\=g�~m�HD��9j�E��nl����4�T��<��"���F%p����"G-
i�ͯk9�p�B�w�9g�7�@ټ�����B��GL�9Ҹ��+���Jit�^�}�:��:�7����N[ݺ��]�� ��9��M"@��Y�9Y�{�=�r�b�Pʥ�}�������s��u8��)N�U%�Qteܕ�/Qi��ۊ�g����8;�-V]�9�l����TB�����h�-JUef�!�Wk7b�۸�]�\:�&Y�hSg�� K����s�rlb���1�!�w�� ��Fwvܻ��0�y�䙺*��,(G��X/H���83����e���� �Ͳ����]��i���-�<�K�-cO^�ĈY��zxv5��,�����＿��HS�o_��B��T�(�%�r;w��Ӊ`Sc���^��,2.;[+,�a��=�*��8D��\��}#MČ�jC4��<�Nf9�Թ��֖m���E1IA������ɈW��寣��c|���b�0+0�է+շ�
�W�vN�Ƌ.i.J�p��,�Y�ʪ��7ж-l��t��uFd;5a>�ԮVo���Xn���t��G�\��Z�&�k�"��p�.���0�v�62��7��YH��׷q[���[�{+y:}���
ʘ*͂� ���l/or�]b�_�J��F\��Ce����M.���{MlxQR�ӧ��;T[xV�\��Q�+�Z���v�v�i�u;v�c�	�l� �vp�[�Lk��=T��O�Д�N��3n�5E��vr���/�ᱤ�
��h\ؕ�-[k��eU��f]�i޹�/�_LJ$�:�$��bԚ���ܽ�=�
<��p��@@�ݨ˂�M��!�9-�������n���Q�@�5���vS�Ӛ��)�s�k�V�ūJ4Z����ԶX�-�m��V�Q�QJ4JP��+Q�h��U�ڕJP�mJѶ�ikm���hմEaR�m�����)h�mQE��[J1�ZP+EhԪUE��lV5����jR��tq����9���W�j^s�ԭ��J�����T=�]y̯x����'����^}�֌"Һ�����}ےg��wj�E���GvnȜSu�Lɬ�[0�����ymV�y�{=�תr����F_+�@kՇ�98b-g	6�-��<�6�{(�Z}RY(�,O�&�a�&"�7�mݧr"o��ᘂ_��f+����H��H~B���`ÙW�2���׻�s�i�F�i�&�B�C޿�Vekn4=z��+%ʑ>���0]6�܎�-]*��_�<��9A���UB=D�ټ���^a�	��m��y����]9��TR#۞p`�3|�Vu��,�K<�_�I�����g����V}Lc�YG4��C=��,$�gk��L�|�x�W�m��j��;stV���l"�^�ه�Q䬏�5�����Ze��p�[�<���ll�Ń<0 e�X~��Y+�m^���J���*H�Igg�I��4Aw�u��
�,3���kۛ���k狊Vm�uy�ߧK<߇_ׂ=��5�\*�&�&x�-��ٿE�fT�ٙ0�jV��{�z������-�f�4w�Έe;��{�e֚�5�X8IXG�l��f7�&��w���ʐ�~XL�B�n��!.�;YS=�Tp��8	����8/�b������L�a�hK̛�ѱ��9�}$�RjV^���Q����l�#B���ɽزxq�����y��K>�ue�T���=~M��D�u9\\���,{��n3����T��n-����]qr^�폎��0EXZ����w~ꁊ���|v���Q-/f�s4y��>z}n�VfA4_(�į�ouM�1�g�q��c<�{��7�Yu��3]�:�2�r��O�-�É��O�(ܼ�{(zw��3;��ﯲ��>�o�N"I�����{��;���wSD�ÈW��0!��O=��u��k�R뮁��Y���Pe�t��+�o6����四��<|�HZ��{q���e�@*^n�&r�7s��2&�.�D����q1��dŘ1Z������&��S.\����-�yy�F:fy��{�x�v��]���0_E�7�5�����N��pU癱�������0Ԙ�-��9,�Z5�O��W]L �@dBc�}�4��Lȶ$g�Wo����P�]ݽŜ���U�/�x6�쨬��+��J��z~W�2�$5}���]�^�/�ܷ�Ga�.f�S�~����>P*���SnjV�}���:�r�Sϖ՛�[]���4OWZ�[ԹJ�N�R�+�Kfh�΋ZT��g<�W���d��fV�MJ��
(k2�vj��Ԛ㡒{������bfj{�j&W䭿j���Ө�����k��+u�<g��t�ԨZ/W�u0(^F�+����ݗ�ÉV[!6�+��~�����+��x��YW(G��Q�52�,��@�@ �ٵd�`��k�)`�27��+.T0V(>A���38�Y{cdP�W}wN��庺N�V�Z�]���`x:
�4&��%Jy�θ�M�Z�o��~YB�byN	36��aZ��N�z���8t"%�����(���*��$7��
Mu7]KcRv���Y���<����r���-h��{������g'ג�n:�*WBf��ռ��&nQŕ�m��g��_�Y�l��aQRuX�]��nc'�@��	ٛӭpi̵a�R0H���K.�c�;� ���Ʈ����E�A3yKq����Y�-
x�)F�]uh]�e�V���o�k�u�k����E�+YZ��R��֡KK���R�-��kh�kKjQ�֔�����aU������n.1-���Ų�J$���Z�C[���Ub��jZ4��m�iA��e�*6[KjQ�QETQ~Ǳ�����0�>y6��EH�]�T�q��_X��#M+�ܫwA��.��f3�Fc��� h����sد�Hx�2d"�)tnx���=~]2�5c�Fś���C�����Lc/;��nh»�W=kQܭ����Lܭ����Z��V��B�mGr7KI�=Sz�W��߶f�����Ĉ�mw\�8[�i��=0��zA��B�(�ݛY�ٵ㧸y��4�l{2���d���*� !�"n	�T��7A�H�P�"����v��ޠ9b��� ��iQ`u�kh�T̼�0�p�x�ྗe��W;;��db3��qú��;����1������PK�d��[��W�Y�� �b�^{��]��fǲ�!r���t�^�@���x{h���{����Ƽ��j�w$'�z��s�4��{E�Z�3H�h�β�d��kW;h��ڕ���i���Ȓݽs��>7Ct�<ݏd��sz��PJ:���+r����x���^��6��D�sy����
5c���Z7d��Z�=F���y��&�~��c8�-�#ܥ��<�S�s,�e$���6�&�8��*�Z�K����a��Q]�/e�5�WD�5�O�n��ŭ����N���.6�`��	� baH�z=3�xMW�Ǘ�W�R9�mX���\��Y��D���7"�Ug���|R�:\���$����u��7O����}I�X2�J.kj>�5ȯV��sT��Y�u�1޼{��7���fX~3s3d/�5	���5���G��:�-�	�4�������M�to�!U^�/{��F�P����J�z�
�ɇ{�x��T,��O3����y���#k�^�Bh\Mk3��璅�Z��2w��f�O.�Pkj=gh,OT�M�~;t����w��0��@��m<��ju�n]e��#m�R8"f-�I��7�4�f�I�T�3�����}r�J�V~;��l$_��v������i�+����wB�wv�OSJ�R���O%t�2wo$u%�e�TE}�N��v`�%�$Uxga����$,P��7��3��u�����6�c��J���b�(;gqZ� ��kC�~���(�ⵌ[��Ժۂ��Tc\��S�@EE��!�f��trB�Y}�5c�D�m)���f^s�ԭ\��>^��_3� �Č�QU��l�l]\")��7�D��O`C�â��W�:mf.�Z����t��y��q�3v�|�(���ak�Q���*��);+��ɕ>f.���<�sۃ�å4%�iz���n,O�&�a�"(�R�S+�xڼ\.���>BWN�mM)�3V�}�w��-���p�y���=4��F̤)q��(ik��k�ȿ�,jn��s�Wq!�f.3rK׾�pH�R�g���2���y�o{܉���Ju,Z�J��*����K$$��g��$��TZM�$���ţ�**�fߊc��"�.��w���=�f��ժ߼����	�l�n�����m�ж��q1��m���Y��1.��gH�`BB
HI	i`m$	��PX�,U��0�,�,PUP�-���K	�dgR,/�,����P�a�r���}I)7%���?��Y!!	A��S�����_�rݎ���}��Ě���n�Kg&L��:S��]�ƶ�Gɻc���T���M:�������D��P�U�24��4Qֵ��!"O�~O^�ۇk�V�]�$�N?F�;d���/$uQ�?�,�T�$��N����:����;ȟ᠝h��!���5��t���%L��y�$���� �&��G�W��w))J]9��ԩ	��T]Pi4%�����*1Q�w�ڏ��me���B{�ؚ4f7/}l6HQ�7��9��J4�^�Ƿ8�r����`��l��H'���g�Cg�KK^�4SR�����H��:44��p�<�)%�,���гUH��\��gՉ�8�7}�GB~l��"I!&�hZ�#5�����Z�kDUT�UR�s��C�;[L�&t�N/��#��R��;妱�r>5Uz���f�'����~�C&'�������{i;�{$�ܲRZ!�R�3��XQ�ts��7�w#�S���G��S�u8���Џ��.jH�]�O>����x�J�9I��RҤ�GY��؏Syv�9����o}����@�%�y#��RV�[�E��ѐ��dj.�?�,6���ԋ�ZE7�B$�(���	|�D�Tk+'Ɖ�V�VG%�sޖ$��3�v��E.�O�L�7bB&���qb�UEE�bZ�e�Q�Mq�S;RH�$�)&KI�h9XNn�@�a�ت\�6�3Uԥ�,O���ST3&t�FRĴ�EIu-d�daf�EV���l�	TY�}��w{#���	��@�%0W[o�'�)$�o��#�wq�~ϟ�-�?:��:Ӡwo���1֌:�\�ذ���J.S���,N���^4�4z�)$Ǌ�QQ�I����w�db�Z@�'[�sdϋ���
��U{V� ��'܍h��A"K$�`f�)�ka�g?��G�7G>'�<^����%ܑ�=lF��TRQ�/�.�"�,�uw����Ufa�CS>�eC��o���O�,{��Utw���v���-&�ne2���pj��	S���&Y�ejp��rWK�E����&�h��B�q6���~��N�%�]f�����Ml��6�OW����K���R@�?�*#�/=��5�bGJ����r����%v�I�N��q�L��4��fe����\�3��ڽ�;�P�N%QOu�DvE��	����n�M��ܑN$9_F@