BZh91AY&SY��u. �(ߔryg����߰����  ``�zP �B�tѳS��ZjR�M�6)X�>�6Cs�$(1� ͋Kf�j(e�}�t\�#E(�r3�l �#@7N���`(P�(`� z]kT.����� C��� �73�-
 ��T�42�<�h{��H+6+�    @    P T��U"mF�dFC&FLF�	�5O�z�IJ0        O4�R@��`#MF�F�3H�5EU=LF�&#	� � �QDA1 	=OL���&�����i�&eD��*P=M�CC    =��c����<�3�q�D��0�z�!!��*b$�DI!'RDI�i�+�.*�h�	&�$cf^���;�{����~�?�j�jW9Ա����(�UR&�&ؐHTeF�E��0�-�1����C�6�'���8X��$kV-��m�
N�$sQ$I£�G�����z��rzU����5��v�F�'������"Uϰs��>�92�""i4�����-r�N���2���r9,o*��'w=��ʓ��ݺ����/��y1�g�{'��NG'=9Tn9��� @��a�7Ni�{�&�$^��E������}1�%Dy.x�$G"c:[8BS(����J샤dD�:y))���)��&z#��2�U���,��DY^.Dj:�n#؏�D3�ĿJN,��+��2:G*W��ؒ����Rs7)��Lg�g
�N,�Bk΢;���eAD�\�n'����e���/l��]�N�(d�Dy�%�i:�Ra�H&2DS�śepa���+�gx�x�p�|eX�|e2B�j̆w!�&3bw�b΁��V�
F��j���j���R��%&=����z�,�2��I�fY;t��"Ҵ��/KҴ�l�
��i�tvG�:�6K����g��5]Z�})���H�xn�k.k�7	�+t��|f�{$��=�'�$��}/rI��C+�~=�qs�&n�ռ=�a����h�h,[F�Xt4f����L9o�g.gZ��T�j�;<�2س4�1�>]�tF<}��7^�z��U�NtNa�-�Q�M��O��H��ҕ��'�wg���;��-!�0�H�$9P��u�%��L�0�5���dxA��g*L�GdFz�Q��OTD�ˍK�*FFF_&�#2��+�-J�JĤ��%cN/a��d5n��;�|�ǅ���X����M�1��fj���	XM���n�Kdg����r�������fy��'rE�=3E�:.�����m�]�{+��G�2V� ���U��O,�7���dH��G�N��]����%%c+�:���2��޷=Ϡ莥��E���y$GA�I��l��=KA{0R��xo��.�z�敦�N��<�|V¸n�	�m�S��v�����#�M��%ɵd�j׶#z4C^��"ZK�����"q��2$���o�\�;��Axx(�q�4����eK̈́��ۙ��`�ctr�+9�ϖM�4S�BaL&�B����Xs��L���vR���#{��&����**�$�	�]m�Q9e�F�}m�!�����y��9��znE�Erf)��=� p�.;-_`Z6'k{w�S�R�Y*�Eb�9�U�˾�g�nz��_!SwXM�}Y+\��:�Lc]۩�D�����p�זdΫ��nr<;F܏�Vm������~5w5��|�ja�Lz�m�L��ԑlou\QG׵�z��7K�v��[���	Q��)ޘ�:���`��EJo�g�gd��ڗ����ݮ�����4[��5T�����S���C�c���vD�1X��ܹ�TfS�:ٗ�/���y�y,�F�V�N�`WYd��^8��[@����'�7y�sW,���,�)�2���ܹ
[��Y�#ڠ�n<i��`�S���\,醗�����v���!<�VmIFߛ_$}��J�/|���q�e�|1��-�|��d�B?}�s<���}���K3!lIQ
y�+���2��U�q�]Z5aY�[\�(�� Y� �Q_-ie��Q�S.��+�r���q֪�s׽�q��/p���~|w��O���*}�C�VD�RaWd�T��1AY|��rѾ[��;�.����ڈ۫�@C�����L(�9��_39�!I>]Yft����g�����}Ӹ��ӯ3׏`{��7��k�@��I���|����as�����O�S������eB��B�Pa��n?�"��+������eeg���T�c�I��
��e�1X����|�N�~�-衜���#�f�y������;ݭ�����Y!]���Hzԣ�ޢ���o�a3��A�:�ܐh�M�;w���fd��׬�OJ�qC��6ܸu� �Yײ��'j�*���cH�Oh����6�p�R���SW9L+����c/'2�����2��9y&d�t�r��[z\,(9Z���qO+ˋE�i�oJ����hnVmb��5��R�J��_��Qs�k��I�<~<�2�2��O"9 QǛ��}ދಞ��*��y�խ��&T]<��6�o�C��q��w����������viӇѳ�Y��wc2\��/�v�:�p�j�n䙙{
n�̀�v���1/>��i{�bx���\3�ע���mq��9�Agd���m��::؎i��z�t�q�q\q&#}竍�h�H�?L�_�;Q�\���>��}D3X�%{�ߍTӱr���P�|�zD�iA(`ˏKfE�
�ׄ�����Y�x�<8P��,]�Y%�|�����j 	j�F�����p���/�OE��F��X��^:w.��4TK�G��)H�v6���v�g��x���Ϛ�Gz,]�mj���*�8G1��!��s�Ά�b��d�<�A,�y1	�[�4(�q�JY�\����=�sSo��f)�5��	k���G����ug[Rsc:�8��� 8�T�t�GP����Anb9F���E*3g�]�����l^���]sc}4�8�Ij��N�i��̫�ޙ��=,�9"�g�vɓ���p��ltMN�����79�]�'��=w&��pu��?���]�EG� O��ӓ�g�Mx�t��$q��ių�[9�HC�|ݿ��D��a�Owl�l�+��h�wWY��́P?��(�&�UC���r����|���UU^s��*��U_-*��;�:��6�a,�3������}��7�U�o��W�����n���F�<,T�<P�jЖ�D�MCR�֍2�}��iUUU�^���U^��UUX����5�?TLlm�l��41!4��*(4�j�`�	z�H���Z⪢����m�n����UUU�ᬚ!MNQD	2��Z��ʪ���D���8���Ҫ�Uxݽ��UUQUUUw|��Fm(�0@�	PPm:7|�UUUx�ڪ���ت��Ҫ�U^氚	5�5��5Pֽ4��&� kZ���:������Un���UUU^*���A����zkZ��$Ԛ�ŞUWU\b���ݬUU�Uz��_�k�D��©d�9M��86��b��t�9;$�HYR�Ul�,~�;~ϯ��C����Ut&�S��Q� ��0K ��"bp؉�,��,�Λ�,K�xJ�<"aӥ�bP�%�g�ԗ�DY=��F�sI�N�˩;�wٸ��]��&����$CvWEc,vʪ{k(�ɸ[̵�Z�	��s�p(J�;`E1˂`�N,�u���#n)�X�!X�Tg�6	�4!�5�r�V��dXZ��b��rUbm�9�:�4̯Z���'c�@�LPT��������W�/�/ju<�Ԕ�T��Jڀ�D��W�-j�ݰ�r�V�Ӵ%Q4�E"�:�q���b�VF�R�[��
܊)_*��NŖZ![tpRX��T�j֢��Usr�X��ÍAl�/uT֬��2RV�n:���Ȧ9:ѕ�z_;g/{�����M��333i������Iffff6�����m&�333I<�9�s�|��N�$��o��L>�"[}�\V���NAHUlR�4�!ɋ�f#�87�U�jU$��\8�b��	xB�$'���~��J�����nQ�b�����O�����F ��;�Mb㣋E� �ĖW"p6|��˪��Qב��N�J�GQ���ۏ_�S[Ç��TgW���>u�x��$�UE�J�"B(�_5�!A�*��Hk(�B����q Ɔh�o���Rj�`��FI�D�։�1ήđ)
 ��kN�,ז��o��/�Gf:����|�����$��%9x��§/�\LK+j컨¡4��4�o1���Uh�\����� j��V>�rM�
0��-ί��ʆj �|��z
�|�((�Z�-�%?�����L
7���nľD6��Z�<�����kWQ�L6���M��F�_`JӚ|�F�Y�PQ�i�꓁����k��T��l$�����?��}1BE.O�,%h��è�8a��s>��#���.Q�j��
�ɺ���ė_}j���|�G٩Z�8B�`|{��&GW��ӇN�p(���s���o�rdL�]{��%u�@����X+j�2��r<��0ᲜU<&ѥ��%�|�.��L� |���{�P�t��ԖTMTL�5� &�jN����AУ曁�!���+g��:5'�uU���j�w�_xD2IP�5�"��ӎ�*�w��b�_�;��l��> c0�M#����'G�H��Hf��#H���F�#�H��i;�����p�(�����盃��}#���,�4�G����8p�4��B��I#[�D��Y�/�h9�c��۝���
ꮨ�������xk��#�U*,��j�l�ع%��Q�O")�4\V_}��MW!�j%�o>f��233)$��%/<@��H�@H�@HA	(P�(V�5d 3 P����nq4���Q(�ŌM,�7��j`p���զ�i~~(4�r�5ϡm�ψ��J�⦣��n�&����d0��do�RO]X���u�؈\MyQ�F�m�R
LLG<����S����B�B1��ſZ�b\�&�$&���U_Qubk��0�Z�WҊ4���#�!�q��Ld�&'e������M�Ek�CcM&�s���t��� P�3F���T�GS�Pզ�e қp�:�"�M�8q|�G:� ��b
4�H0(�m�y�$����3~P�l0h��R}�W�����+CH�9����Y�i12�	��T�L���3�;+P�M�lrH���A��4,�y��� ��{�	Y�P�mC ��u�	!�5�>1%0�HSi�ZO�o�@��:46�)1/�JcD�"����IbG�3I ��N�����#(!#�U� ��d�H�g��Z�����h�5 r��t�JA��Z5/5jS6�b���^[�өF-i������FQ�^%����'��兎1FD�۴.E<�c���Po��QfM���uW1e��Q#������ 7�ȑB$�jT����i�Mq4��&��y5�5�6�$�8�N��-9(����^r6�-�R��\���iш8���J>m�ԯ�� $�'�d�b��X.�#A�pm�1���q[!kCM|�@h�14��b��:����6�t�Ȥ�ʄ�ޫXZ�d$À4P����]hᄒ$�Y�ɈZ�1��	,P�c�j����&��O)	�q�t�ʒ4a3u,l���<�>;���5Z(�V�g�PW���-,<I'IгU���ah檪!�����R�q���'���B��sƩ%PB1@u�a_w�Pub�܀�ӹ�tl�d��0�����H�F��4�tz?g�g�?��!��4x���ai�ǣ���8<��pvp�<I㧉�~�H��>4�G���߇8FE�I��#�a�9#I#������I��sﺭ��I��O�\:�a���'rE����؇���InB�Eݵ�s���G"D[�.���=2�g����q0��Ű}��z�wZ޴��ڲ��8M�cS��wlЭWd]�����W�s��kr?%�P�ȩ-���͘�1�Y2��(�mv[Ɩ8�mUj�I��'���RO�G�׭��(#�A	 PG� �� X� ,~ ��R�*%�ˊ)^�زq�4:F����n�	�6:8JV"(� 6��D���������U(��&]�*f&%�2	?%��g�:�ȶp"[j��ը�|�p�P|�R�(>�|ؖ/��BIyy�KK���������
$e�����O� ��vχ��r��cE�ь��ռA奒���,$_46��AK��m������:4aH��y饒3�e�~tKq66
��&^P�T6�qPw��{Q����Bs�9�����*��:�B���G׫>4����xa �V-��T0����|����"Y�Z����@qU#Wͦ�����<A��BO��P�m�:yM�F ��Y9�_K�;UEEӪ��l��'+�7�O�N���
(�.�li���
�
�. �*����DF�PZ"��TuXr[l)uj5�,��!妬��6�FD@�̳���`}��B��}\G�Y� �,-z2�,��[>(8^/�e�Z}G�T%a��_
1��R�,}�q6�����%ģ删���p�e �XYr$ ���i��PZ�����p��`Y@��
%B��/����,/h>R��Ł�;�b�GQ�����ƪN8AAb�o{\��&UM�i�_:K����G��ߐکC���2|��ja�CG	^P����?b3N�si�(8F�������uqe��1�O]6j�5f&�	�euu.TY�h�+�0yJՋ�:�g��"�9ߑ]vk��O�1�-M�*�XwY�������>\9���#���ύ>:AA�jj��XT��r��*�JM�ůY�|}A��XPGԚ����1�,������hP`��tw�+����*��̼&H3��1����<���#�I��N��ӤQ�3Hf��#H���F�P��(�$�,f����:GC��tvt�<G���Ğ4�A�z��i��ӄp�,z9���L=�$i$s�+>��"Ϸ{z�De:���7��~I�7kGgs��_GM��+wz�3.�U�M�q^���*�<�WEM�W��{�Q�X{����      @`~B�!B��+Q��r�|�1XB��e����c-G(V�������!��C�_�G0��E�.�a���`�)�t0��וj5c8||AA�e���-�J֩4��5�a!��\p�����,�X����2��5�_+P�E�~���K��a��Ah�O�:i����߯܇��v,i������1�i}F-ѯW��u.��2)ƚ�)8�!��0��J��d��aJT���
Ԣ�$�YE�{�P�� vծ.r�ŀQ�T�����E b<::-�܌`�v�(�a}\a�PqO:+G�S��D��^ZQw�
Y�/�u��]�J<f��u`a&�����-Pt��	08|����ksЪS��+t�T���z����QA�� �GԌ�A�Ġ<����N��V�V���с�-|�D�>$�����+�PE,,2-�gL���RM�H�I��Ϯ%�ՍRP�%(�A��U�7	�GV���x�VJ�4�gN�>$�>9V7�by����ҲY+mn��X�"U�MKVp�U�P
�a�{�O	���Q��G�m�)��a'�~EWiZ�ב��'��q*�5��n�f��5��a�t��L7�� �0�m���Q�_+-Z�a�/p9E�̦��{��r�\<�Q'�P�߰��L,]낉	�m��0�.(c$vA$4q2�I��f8�I<Q�*�T��DF�h�V�o���ns������"Xt����8V��D���#�/�MX�)o��a�K���{��%. VUe\�\���_"q��0є�q5�:%c�� ��
�q��E�>D���+�E|���^�����GI5^��A%�q}����Y/�R��:zZd�D��'��F���N���}�f��#H���F�P��(�4tY5��Dxx>��tvt�<G���O��h�����4�?�K��#��g�#�a��8�h�(ߙ=�P�]`���,�
��"������Vt��|�<O�]���S�+�;��*�f��+˒v��Z4�Ԋ&��1�Y��Z���sr��j�y=��[:�r-B�}��
�aefU��(m˽�˽�oW��"Zen�U�t��L��s jͿ>M�&��m#x�D���ƏSQ^g15'+�چ߭0R6�b�mYlҴM�!D���������^����@    P@  �P�jKĽ����Դ��H5%����9-�u�`�Ր� x��s��b��Y+�T)@D�qђ�X��,���1I7��|�>9z�W$�*��D�Ⳬ/�;/��'�S��GZ:1�;��$�2���\2>��N�"
�)t�>�a��>$��Y��e�����=�ID�$f�dIǨ�c09�����^��)	$RF��k��\l�J����^ç$�`YF��jF?����E,zI�\e*5A'��k���2�0��TuB����3Q��,��Tx
D+g�x���g�7�>�"��TUC���X���S�e5$�&�φC����pՂ�e��D�W�X��0h� �$U�g2�V�R�t�J�Y'C�e,�Ey�����hKd��iw0���G�.,@���䌑�!@dr#��H�ԗ�E��u+W�I|���B�!*%\\���
HF�Q�J����4�Y��K�x��i����h�I�$���H�Џ0���c�V)��II�8��D����t:��s�"�����kIPUR�IVaԌ��e�5��a%�����C�d$!��
�=�l����n��˭5�)����Ku@F��������]��E+D��Vt�I(0,|����CD��<n>I �t�EIT�e�U�J+�B;H���:�+Zqx�D�=�}T�K��6-IWR��yEda3w�;�nM�����r"׫�\��[c��c%j�r:�p�w�~�N���2O��D�ܯ/�c�����^��K�)q�W��_$�#&l�G��!Ei�K*��c�!4ymy��L�ג�("uq9�Х�kh�I��t,���_"��Dעօ�<b��Cֹ�����Ń��x���qQ�>U�v���/��LZ֧��_Q�)#�������?F�#M:N�F�4l��h��I�a�EF����|$�������y�$��=�G�џG�#�����?G��G�ɰ�$����D�?s��)����'�?7�og2s��^S	��77:\\�	�����f�fO�H       ��B�J����˓|����X�� �"����ώ8m�pľ�-��A���H/��Xt��$�#�˧8t�'C�gŵ�%��IəQ�O��V��!�?D^�3��(F�B�Ф��_+5��S������d��_V�i�L��H��u1�Nʆ�EB�EP�Q�$""��N�Wb�t��RJ����#_\�/���Vխ���'�Q/,!5��b�Σ�U�E�,ıp�W�1�^�
�h�a����➢� �NBϷ"c�&!u��p�D����j�Q�8ן9MR<E"sU��
��]�ڸe�bՄ�k�o��IEto)�,E�_,�Y*J8* )nQHk
 ��؏Ob��t�xph�֢Q�	J$�p$���"M	i��c�h��/I%����K��A�I���ljH��		$�A}k]������}K�h��.џY�F+��G�4�Z8�n�b-Z:��M>�ψ�\D��C;2A�<�z7��r�EVӌ�.(n	��L�3$�E�� ��ca'pv�pV�/�N�+񍖸�������ZϦ��
E> ���l\���^�@������"L��G���p�AkР�-|��D���5+>���"[��}��>D#�|�Q�^T2�_��41��Kk�#���N�5�^��X�m��֩/CIHT"T���-��C��m���w����և
1yj����k�%�R���R�aԭ�b��8"��8�i�R����Ӕj�G�}�mǖ����֧ܓ��oO#iu�O�I�I��g�Α��zAF���i�e�>4���z�1���ri4l7c�H�H���x=�H��o�H���G㇉<|G�����z?� �|8l�'��d$�Ñ�rz��r_�;��Qbx,q�	$'��Y�i�t�{�г�.�/�5U�S��9�1�y8o�s;�?��Wޯ�}����H�����2��,�l�����Or6��.�d��w��U��U\E�"jj��2��{�s�ߧ��8Ckq�c�Ԭ����g �H�����qu��`V�r�h䨴jv[�XjϘ�6NE�A4��U8�>��+fmCM�W��=�            ��T��J��5 P��'��QZ>�"&)Xղ��P��)�V��X�j�e�[Ƙ@M؝�Q�njJ��Sq�;`��]�^�9{�z`!w����I�5��G.��t�D��(�|]ѵN�n�y�V�#�,�C�ˈ�f%�%q�_��p��:�x����@H:�Alb����#�7��?.�ۥ���KN�r�E�������>D��"
O�>@���c���GV�>^���k�1b�o���M|��p�'�G���.G�8��ů��g�T��^>^M���Q_l\���:�Z�<L��b�4�(F�O�z�(���aF�#�}q,��ݺ����Dqd��lSz��n]��mnnBY�JVY�q�+�g#��V"��QV�??�� �-jTQ�>�Q��ET-J)#�@�ǭSX.��N�QH�X���6L�b;\~���j�R�I�1�?N�Ο1�׆C�V�.,F��]\G�P��- ����9�ȇ��gR+�(�(j�Xx��8�.,�m=xD���&%��q$��-y(E#�j5�8-B1M.Ғ�`XIm�G!M��jϊ*����a���l��G���Z:�T/��vQ{��8���q��VZ� ��(�ώ�w�<}���&�.�E�\ٜo̲d����|�$����L �&*��Ig)���APR�K��X_�|����x���8��:�JD����y��|�6�U[oG�
���Ji�4�ч|�]Q�-���qG� �A���i�UO���m\�U��>^�� ��Z���G�W�O�h��:���g�TA>$eE9R�
��R�"��?,i�O���}Xi&T��!�?\�!���G�L'N�MM4���f��#M �H�a�F�F���0�$�G��<:G���t�oH��z=�G�|> ӄp~<Y'� ��~��$A��Ko;2��;/��߷D����;���|M��g��f����ۋ˪��FKtc6`�V�ňřx��,Z)�%{]�   J@       �P�iZR��~�E�~Z<.C��kƍ�(G�6|�Q��~LBqGh��{�¸|�T�V�>Zp�<Y�t�aX�}61���]#�oZ/�,�#�V�4��Ҿ���e��"A���M%jW�UK��7�%=���T֧�b�ܱ�����X�Ε��mX��[��$��B����dU��/���<\qr��M��|��J9����%��n!�U�DOp�m�Q�Á&p��Df����#�%�ɴ�G*���Zs�~Rum��hҎS>�|�(�����pD'�����7T�u3��F|5O�� w���O�K*�l�څ�C5�7靣���Z�k�/�����A%`t$g��_2U���^�ϒ�;�Y_�5ut�j[����>Rz�l�Ś��J���(����|mD�ޘkӘ��Rxgze��1�l��w���S�iF����:�K��$n���b<�_agS�guJ��A�O������ֱ��}�QBT�1���ţ��e˗23�Ĝ���k���h������������ڡZ:��E�3�h��~"�>G�#�^jK$��a'�����;�ǋuu�u�{�H)PZ%���m��\G�Re�T�>�5�%�t0$v&<��,�	�iJ��Q�5+�0�N��"�|�%@g��k�D"Wh�r�T7�6�i�C��ē���4���tu��K:6iGai���#K#FQ�2�"����٤<GO��xz?��4z=Ƒ��p���-�I�I��OC� �ð!��:F�VW�'�$S�h�YN�"���Z�h��5T�kv.v�<�خ���=�]�t�?�EW��:¼�]^�m-m֎�<��WF�y�ڮI���eX���oW���^�W<��9\�+$]�)��q�Q5��<˙���\O\s�f�(fLdT3��fݪA�e��mũjkt�]�������b�|nj�M��+kV��5�[���F%#!`�ԯ���O%�MښM˚P�9����(�m�`          �RV��ί��ph*�� ;l�(�$���!F����dv
�rT�r���"Z8Ӳ�,���*�Dhu��
���KH�ND�c���da�����	T�2�~���X��(�Ж����w�﾿c�5H�I'&bf��1Z��0:X`{ol.������Y���^�O��(\���<�8���ުJ��A���!Õߑ�lqa=�)�Z���:k�E� �Bz�>����}|�t�8�b����	0, ��}��"��1�5�W˒{
���b~��2�Z�����lc>X�yb�M��*����������:`X�5:Ӂ����1<̏H�n���e��E�#��Ф�m�hQ�"Ĺ�z�A娓��w�Cr�x��jU�8�:�pLI�*Z�+\���OˉOa�AgH,�t+i�����U�+�-�8�'z�13,zKn�;���㦾F��GC[�� ��%�Wv"%f���E���>��||X��=�lld.AK�{4�pk�w�H0��F�w�.&#mPyZ���; |>W�i=I��*��1u5��������T�i%�8(g=��p�ɇ�6L�B
��X�5�q��%C�ʨ�F�TB���P�o�x<Z$){��m8D}���V�x�=j��U.	�עHO�5���֯�_�wW��;&��Yi��=E�Fk�+S��XSli�cdCm�����G���,��π|��>"���� ��ٱ(ؔlD����f�,����8i�Ɵi��0�ϋ> ��M$� eG����ϥ�de��^��9���y�Z:��p�S�U��sg5��r��l&w̺s���GU���Gd7<�;k+��Cű�{��B�iwJ|�{&�"b|�v�[��S��8�a��"lB'���n�s�7f<=]ߠU�>:�3K���p�       #�
    �
U%K�6���X������ƼؕF��Ǎ!}Y�N���e�ϛ��Y�|E��ojïDb<q�\G�~}���t�>�7G��B:����|1�j�K���C�(�?i��IAG��"���'�7T��l�9�)�h)�eV
Z�Q�X8���x�Q�s5�61q�Ǹ�Q��պj����LB�N(�\G�[��C�Ēp)���3�	u��yr:珔^UKϫ�����O�\�I ��B 9�voWFg�۵P)�u�t҉0(����&lY���6�$�D�cxj'��t�ɞjcjO.g:�l�d��O��E�#��8gÃ(�	>
+���}-Ѿ�D��Toݾ7��� �*��^gƼ?�[��CU��zx>C-I��I$�L
"M���(�]cmr�ʥ�&Y����8�ٖR���j>Vƣ�R�B(���@�<�w�ΒH�^��(�c\%��Qt��W�/\4�oPΚ:G�p�����&[rV�\F��6� �^->8IХ�]�E��W���E���Q�~m�+�H��>�l��FRV�R�P�kb�^��wV�h|qUI��g����Cj���-ǥ��W�R�);�=#i�Ww�4,��I�F�UO���O�Q(��y����M0���i1�[�"""�)q|�p<"�J���Q�K���s>�v��}D����YR&a�d/�GLQ�_&�g�S���x�J%�Ե+�T�l��m�����!!����O��{��F�s,|e������,�a��k,��$$�`��HM'q�PҎR%2k��s�&(��������E76`��&�&!JJX��RȥIK
XS*LAJ����K�%,)aK
X��&�)R�%*E(��R�R�J%1I�
X�Y
Q)Q)b)RR�)a)R)�L$R�K%,�*E*IJ�,E)�S�d0Y�R��%,�JE,�T�Jf�)aK"�
RR�R�JE)�)�LI)d��)d��*JT�JU(���*R0����)�ZLJl��s��Uf)lZ[�e�lPҌJRU(X�b��F"���)�8&e),�1P�P�B�0�aK),��p�,�e�T1)eE�����*�),X1Rb(YB�,-��j�Vpf�b��%��T1(��KJ�R�0��J��U-*�)1U-*���UJ��KJ����T���YRX�YR�UUUe,��VUR�*����p�m�-R��1QK)jK,T���b��T������)eB��J�,U���X�eK**X��"�T,�eK*YRYK)Ub��,��~#B�*�����b�*ʵb�U���ʪX�b�eJ�,�e"ʖT��h��ijZ�VT-*�f�*Rʪ�Rʒ�RZJ�
K��Ib),)*JK"RQ),���K�TJTJQK"�B�IK�E3�4���K
XR�J�XR�`�*fɆ����K�
X���JX�X�R��q�1Gf��ȃ�1u1�Y	�@��6jC��E3�1"%�!*Ȳ�ʓu��xَߏ�ͷſoOӹ�:f~�1�ق�5<?v����?��lUi��f��4y%7��u�خv�Z���=n�~��ڮu~?ǖ���<M'�O������	���oZ�i�����lca��;y�i6�LtA	䎏���{}ĳ}����)?z:$��pGm� ���T��Z`29�$�Om�����:Z���Gj,bH�̟=G_�'N��g(ɇ����~OY���G3��W��n|"A!M��'���ч�z��-��a��}�#kD��۔4';�,lZL�B�e�(Ͻ����f4qid5�H�s�ֻ�Vެ��페m�G��2kV�8,�-��71�mr���X9��H�YkX�F��6$4��a$Ls2��4�M�I#%#�Ɗ���H�"ԌT�M��&6�D��`�Ë�F2bd�y�Oիq�6'.���'),8R lQ"b�D��RҨIiUH�$"�!)e	r�{�i�e�Nwa*qF��;]M�$���}�O�S��؛U,}Vq��S^�a=���|���-�g����0�6���	f ��c�&	[Y�Ja�$�[��>�k���aչ���F�����6���� {|X>�;�;t<ǁ��b��§�}΂��#��:Lg�G�n�=���+�<bA!��gL��b).g��\{<$�{�=�N���w=eڌ1dU{:ӣf"$HUj����O�"�;��v>�Q�p�̎�MQ���2s��M��&�{b��b�r�$�5Mbt�lR��ۉ�z$ᄣG	�1bI"�2=�n��x�M���7%��jSD�*c���8�0��m���G�-#��b��K	e��\�Tn�n��47��7�BC�`�W*��y4y4zܐ_ԚlwD�C�4��D��IN�<��OK�k�;�O�������9��͎�x�@�|#�h�FDvu����	|���Ki�z&�����,'�4�{��~sr~���I�?=O���[Dfξ�u�1j��da*I�����$���]�~������zDr>�����:��':9�����r��%m�,���l�Mu��J�Ֆ�цP�^��M:Tݧ�Ň������e��L�f������nFƮ���܍SM�t/��˟i�n��ֳ��d��41�=gJ:S��2��s�N��lP�ߖ����s�0�j?V_���H�9���T��*7al�S��=��4I���|uǅB�"M	Rg�4�0�w#{�DxE��^��#�̄�:O���$Чa��6<��XI�7�w�z�����yE����i��,I��t�p��g���"�(H~�:� 