BZh91AY&SY�;J:��_�`q���'� ����bG>��      y�Z5V�J�6����44�l�T
*�)ZFڋ`��h*R(%���I�*�T�m��e
�J�j��FU���`aY�}��ք���*MkkE�͙aM*UT�5�I�F�VRhm��l�����U*T�i+f�&a���խk# �>w��5Uj�x�K)��X�;5�٫jmkf�کV٪Ԙ�[15U�T�lB(�Y6(����[�IKj��*�*��VA44Uk*�qR@٤�`   bO��:n��j���U�AUU�K��X���m�WkZ֓u�W;���"ӧM�k���˷kk��ի��:)�#��S�ҪAUIT�Z�ֱ
o�  �ǪZ n+uAJ[���&΅���N�@*����Ն���; � ��\�J\�p�P&�4(5������4�U)�x   �z�^� [���=.Ƅ��5�d([�`u��Х)Tm9�  ���ST��{ǡJR����� �-�{ǥziK<)$�d�-m �T����   \�ݵE)y��t�OB��t��GE�x�t�

3�p �M�_x����nֽxW��u{Ǡ)J��  ��t{�P�z��S�Z2JRlj�63F6��  ݞ�(R��� �F�J�7rp�%��
���� ��J�)B�r� R�Uuت t`Pr�tZhmJ���&�Zʙh�׀  �@�g���P�Fu:� �ݣ�҅�`:����
u]6ۻM�@:�gu@tV���ݪ@Ӻ�s��
�tYa�U%)��KCm��x  .���P �-y�tUW]n ���t����tgJ��` �� �Ƙw`��h c��q�U&�*٪��"�Vo  ܼ �0( �F  L0�;]\ �qX�4뫅 �� 9tۙ��7gh�A;�mJ��SM$�RB�� �/ :oS�j��L  [�� hsQ� .�:��;��P
��
�5u��ڌt���e������D�+�  <B���Pn�\h����  w� tgF�@�.r����5�@4���wqT
��    ) �50T�T�1&400L)�4b��)d�M0ɣ�2S�2�E  �    ���J��`  C  L "�d�hhhT~���S�Q�CA�z���!�%$�$�D���@  �[�F�7R��wo�|�0�	�`�-�:.�F��\=��m�2ڶX^����{����=�_�XT UȂ�*yD U��TW��	���u������jT�"*�����C�TW�����TҢ�+�����/���S��2��̦d3)��3)��f0���&a3	�	���S09��.`s#��2��.es#���	�́�29�̦a3	���fC2���&a3	�LØ&0���&a3�L�f10��&a3!�L�fS2��̹�e3	�L�fS2��3)�3,�f�a3)�L�f0�I��&a3	�L�f09�2L�d3	�\�f2���&a�3)�L��S0��̦e33�L��29�3!��f	�2�̆a3!��f\�fC0��&d3!�L�fC0��̆d3.f`s!��f0��`3!�2��d3!���G0.eÂ9�ę9�2��+��+�s �`Q�9�2�����s*.d̨��� s
a̠9�W0"�P�#� s"e� L9�0��@�#�s*`Å9�d��s `̊��0��UL��3
�*��2��D���@f\«�&P��f\� fD\�fA\� L��W2 �2��̪dU̠��W2�0��T\� f�)2.a̂`U�
�� ̈d 3*��`3
���+�s�eD3̊��G0��L��W0afC0��̆d3!��fC0���0�̦d3!�s	��fC2�`̆d3!�L�f0���`̓	��fC2�����f���S2���a3!�s$�fS2��&d3)��ff09�̎`s���33�I�3+���3�	���)�߯�Ly����������pKR*£F�T�@�̛���0b���Ѵ�Y�N,`���=Hc����/�QИ�Y��k;���B��c�Zj7D�hY�:�hԐ��T�*Z4^��%�Y0�+�	�n=�.�-�s!�zz�y����&���A�,L�2)���J��6��v��*��4_��f�ƁJ��lMK4��x�k����wBm��p"��N�됩𵴞&��O���%d�:���[�Sm#��2�P	�E~8�T���V2�A����X��4�H
�1���5��N�b��EX���@��yrŐ���Ǖ�̦-YI�Hn���KF)��^��q!Lb�'l�.�A��1�ma�֝��*���T��ulE���%!VmAz������� 27vl���s� �M9����u[o�������^,M˧V�h��0NIH��ʖ���cY�k D�*[p%�FȞ��NR.+r���φaU�V�Suɚy��̙�l��R�� HJ(��s5������z'�2��#;�b�\�A��F��t�N��*��Y���n�A�\�K�j�A�gݨ��{�s6�r!.Rs(���?�!%�a��^a^�6ܫB$�b�gp�R������h{�M�<���A���/jن�x�y�tRtU�ctO�C�#��<����8�D���k��e��k�,ðh�ئ{]���,���#��2�-�_wkS��f���2]��S�'i�Űd�%ӧ`�16Q�r��n1�2	�^�_�+u(��bRQ債���:42��%n<��e�z�3i�4fm�#x��(E�։M
��C�x��W��[�6V�ebe�E���Q�x1�v�,�F֍�c�XȠ��#�M�J�"�	���K)��[F��	13f�(]�ś��GI�d��E�����W�P�N��!���Z���c\I�9E��j�ջ0LB7���7r+� �:���D��z>��Ej��������V������/X,A�)dӺ��%W��H���W�+�� �E�C>8PU�����2޸0*��^ڽ�Z��J��j�n��˧M�Rm̸�N���ܖ,�S��8r��i�#p8mC�	-��ޥ��@15E����[��!seD��׋l[x7�Mix6�@-^l�tV]Z��cX{Q���t��5;�u��m;��*�';������QI��H�y�6lfoE��\Y�*f�Uh�i;�!&��fء�Ȅ�v��cFnG��`�˹��W2��*'��N sFlM�65vi��h�l�f�T������)n)��fl��c��,q��������!�u��e��
��Ƕ/i�ч �(L��5�Wf�2�Q�6�ǷI��!��-^�pUc�zNm��&�8&��+i��Q�>4��*�Ȱ^���E;u����]JYTĚM""��Z�����c+ic�2�8^P�"��6˛��]�C�VnM�2d��x����	Qr�X�Yl3.����l��Y͇p�Ee�f�Uz+�6)���[�,]
j=u��h�e��j��Xݬ�lx,��oU�NՆ�*�z�J�|t��
D�wǫ��_e�W�bR��#����6�%^Lۀ�.�����k
�X��t�f�[qʰ�ʃЖռ�VR�-��6*Yi������"�U��7%�M'.�h(�FR�[�,�!���'�e�x�kMRz���Ȭ�Cs3Rt>�& ���t�f�*�b+�q��h3)���!0���$��Z)���Z�j�en�ӵ�&�����8-�NF�8��z�#���y��,X�vΪ�����˨�$�h2�Ż4�*a&��,=�b,76���2ea&�u����f��o5�=č��z�X�Fc��Ml+��jfc03����o>�fQ���ӷO$�[��>���N��I���Ֆ0h��kF#W�o^��V�m-o5��f��ͦ+q�0ˌ����#�r3t�`�Ч�&	U�oq梯�%B�s����	"�vJ˶3l�v�(�wv��FKͤ�-��qm2��Z7���lc�H:�!\����gLׁ�q*c�l�v
Æ��a��"�@#�0�Z�h'$)��w����SS1P:���1���Ulz
;0�*�h�S%ҹ+R��
�9�Z��el�Re:iɷ��d]
Q�)��&m�uJca�� L��CA�t��5Q�UlF��9
WD�HPp�gF[`bDO���Hػ��c�&0�Q��-�a�޲���3��Y��T"�􄤺!9�]'��K��źik��6����J�J�X1,-�M�o\�.,���M���X�f��RZ�&�WF�S2��X�(3wn��ƥ��KN�,�n`�Rf���V���e�ؖ�[;�$��"�Si맚K�vu�#�6���*y��YNr�o��^h̙%��`��u���fR��G7inf��-V\t�b��M+.��f^���?ʔU�*�F7?mJZo6Y���c��ޡ�hdB�[X�V�dDǰ��T˽Pҭ6�Q�u*`���e�D�<	Yے���[a���vƮy>�)a=��K�Z���-���<�>`�N�� �\�}�y��,@����{e�4��N9��A���T�@��6�ӯ�n�H���J"LƙUr�bqe!�u2�+9�����>�-U��	�h��X�(3�m
-f��X�vl02*ªӶk5���#Ӡ;Xtl�@h�&��J� ��i���w���Sߔ��R���I��2^���!X��������;xAE��\��6���M�N���kbm��ƾ�3Y�īe朹�nL�)��'���Gc�r2tU렮������?l(2wa��Tnj������%��[X^�j��W�q'�{��N`���) �~���fɓw]"/bYz�۩�nAx�%�5�f�%��i�oN�w�[�{cqm^=N�?�2`o(ҩ�Z���@)X�v���u��\.�lh�6��J�G�]����5/A�r2U�KUv.�:�z�r]�|���r�x5Z��� �9b�C ű{�]ҦAT��BnQRYKw.��*����t��M\m�-7U��u5P���ۉ��k���(��FJF�;�k�ŵ0f�V�f��h�YKL� �Jn|坦V��r��a�]�)�m����d�E5���Uf�.[Ɍ��;
��{�Cn�u x�|Z.�����	��wjM���6LN�%�i���g�y���D;��*�ZC�qK�,�1�On��J���ۻ����cQ@��J�;㜷�V�d���|@�C���"���Ĵ�|V��A5�Vn��F���+D��6��d�t#q�.�H��ŹY�TH��Jv���7�U2�.��Lǡ�;�6c�VT������2L��Lۙ�	m]جKZ����B@7.kb�v(Ip��5Y��)�R$�j�>GrQ���l�V�KNHs1휳 d6����ۭ	�N~�ص)j!a�x��̽��y�� ��%��R��к2��Z���Kl-�+�si��Df�/x�w1���FS7[af���$L�0�ce��㺊x�ɧV����7&D���L�8��4{���E0$Q��Y�;0K؈�4���2R�(�5OJ����ѭɶ��X�;z��[�E�v3��W�����x�t�.��0�5u� ��zr<آ3fS�z����u��1��t4n��2e.�Qj�&^[4iU�m3�ӊ�X���ޱ��p� &"�U�a�5��v����9 �Ӄn�*�0�yM%r�dm#��%xւ�,�����72�M������ų�3�~�]-�A�H��>)=gt5�<���\�#i����r��tN���h��F�fK�e�T��2��2ܵLY$x��B��|vj5�%��!ݾ{ϋ����QG��v��n��";+N��e�3.�B�P g7�)�{�'(���]ݠ5�t,ԧ�DC$9�~�g���)�k�ݥ�h6Ry��[�����k����1����Kd-��Y�wH�/\�3Y��c��#`�a�Vl!�wDة��k�]�MDT��^=�$7$K2� B�D	�v��(�zP{Ki%Z���X���+$���q\g5+fZZ#K;+n�H��(�i
�t�Y�8�����$Ʌ��D����c�Ŧ�y�k�V��u	Q���ˡ%2J٥�r�� ��MOv��x�`��-ؖqH�3v�e �ٸ5'���C�pJR�G2�:9$ �rYٗ�̸�,
�ُ�zAN�휷%�xX��-�,`��m��m�2�ц�K��%@\���MP��U3P��Y�Xali�Z����4Ƣ�B�VY�0��챘��Q׍�-�s�ߙgQ�KT�� b��ճ����^@��p^�c�P��zj��@a����6�:v-n�[LQh*�T��V�'�d�X��[�jM���ֵ�cB�(jdd&L_�0Q�״^ЦEjM�CE2A��Fnհo��,a��hk�-�a�q��a���V�^�(�{R��գ.½h$kSj	N�ڎ�䔞����4��J�;I�ִu��9�EZv���2�3D���=_k�HwYk.�6l�����~1fhU�`ݣ�ZV��{y�)�Ɏ��H�7�W��C* 6�G�	j�i�0թ*��׋Lm�ĩ�`ދ��q��y(�&���~,jT�v�[OYW��i�\Y{F�^��=#�q�yOp7Qݬɉ�{��GK`Es6L7�ڨ�%F���F�J���J*]�ǚ�\��T�Jl���o�AE��Z~0Y!�6��l�p�j��fEws~��A�֋³�e
ch#����n<,TR����E����Y���%\�����[p5u�Oku�BitR��Ue�uu�ձ36Uͻ���A�U~dbF1ֈ�^�qV64���^[e�ԟ��܃�gHE�ռN���pf���r��{D�m�D�h�N:�5��[Yo.�� �4�0�!+,S&�Fb���)X�Pd�n��%F�Ûםi�x- �J�&�~j`�j��Ϯ�Jnm���mVZ�ϖ	�蕻��0�Ch��:�*�xU�h�n����qsko&쫰Ƃ#	���7�҉�Wz%k
�����1�()�n�lȤ׷O2k�d਍f�tta��5҇˄C0�6ʎ0n�MFA�A�̎�E�G�]��yH�d�`�o�Nk�hf�K�k.�ݽ���Ѻm��R��7d�X�B�
��{N���Z�q\pnh��Y���kaF"cj�J�{5�"���Ӓ�ٻ����L�O��hX��cP�bD���D L�R���IA
I��7i��b��K��a���1;�1��OBm�Y��-CW�+�c.d�P3v��-
%U��M�ʉ\�ɱdL�*N�Ksr��`����1�b�:֐h�I�������i�J�h��ifL�O��>�f�h�D��4�����8汚a�,Tɼj�2Me���x0�FL�S̃JI�h�D6-ӯ.�
]謬�caV��؋��60�^�5�kJ����`���|��UJ���\�ɸ7K�mB��F���*�dD��//"�Z�s$Wg���Ҵ5Kpo[�[�[��ɲ�ڼ����ځ\v� L���d*yZ��E9�^�ZR݅B�v�Y�[khk�E�)�[u�ժʿ����ku��,>��ߌ����	�*Q���;�`6\T�Q-7rY�ϋ��ҵVVA����5�]�råɏc����X�1ez\�-AZ�I�Z̲��ZJ��ABv��u�ɰ�*^V��V�� �v��-��h�c�;m+�W�-�RJe�I̫�S0��X��:����oAmV�EBM��e!�>=u�v�������r��sNS�D�a3r�8�ˆܬ:ʦG�w
C'�TIƙuu��%m�n�ASc5km[��X�_�n�^!N�"�;�z�Zz�m Mpϕ^����E6Y'��C� "):�ۦ0=Ɠ1�I�<�	N��6VQ{����D�w���[G#��Y*XY�dn4�dg^<���^�]��]m��0��w�df��ŉ�Ӷ	��4�oT�W��<�ˑ4�\���E��%d�2l��eCa!r��6�-:%��%�n�>���b��Au�3q�ܡw(e�|��I㳯�2됣�2����A�ӗ�.��ۂ����V-�r����TB��4�8Q�hAu"&��1�npe�s@ԵAJV�V�K��H��r:0f)`"S����5ZӷO�V&��C �ҷK��Z��BY������r��X;� �ul�l�ĳu�vڥn ���+H�L�y����{V��������Yt� 6� �~�>��o�$nQ8&ɯWn^,�^K���:�]�50Y	b$�C�V'w�ޫ�9޶�m�J2�#`PgS�{�)6�_cnT�u�	����v��st@`Un�elN.���1P�J^3�gJ.w-L�����u�`[TO@PZBX��FN���nP�2�i�)��;8��l��ķ ����f$���I��*��F�KZ�u�1ep�&!]�>��-�}:%h�Ĳeҋ1H�Nq]�QŊ�NGS`�Y���\�-.�ov��A6�_qE��������_�`$F�A��p���P�XƸɃ��򜏼��粮�M$o��#��8��v,2��8ˠ�T'DP�)�G	��	ӭ:��ц����6i�W�ٟ��LO�4�L�D3|��3�/l�w�A���s.�@x�N�⶝���;��]��5�C^��5�
w��[�Z�9�70tڇ���ԊH��0��*�A*��Bxo����?�a��~~7���_�X}��L�����_���曍�R��\褡37�w��+�����{4G�%�F���N��,�ٷҦtN㹑��q�jkɔ�(�hK�cT]�c]j��3m�ܫ|�e
��ɏ^*���a�;�׉��dA�zd�}�SVz���u4��NyC�s�YS�^�
����U}�PTׄƆ��4�]i�ՌU�jl��0;+'v�ةj��\��PB�[�6��v�R�k{��e��W�1� b��[b���#'Ne[c�;�:�<�f�!�pʲS�������֡�\݇���N�q[��_����F5&GN];8\����5VL����WuRqv&n�ӱ�
�4e]���)�W�L�����-��A=�l��v�mN�L���w%�c}���U���R�=֦r;��o���]���լ�h�{��y�z�ka �B���+�'��WWN�%Q�w�qU�M�6��l�0ru��z�o^�%�m53�(� ����4:�a��C0�G��(��w8�A��m��k��oq��גCn�l��wy(ӓ�6����'�
�:̫�#���w%��z�z欷:L�� &[����I:\�]����\�qN���f֮��er�����l:N�砍��+CX{N厌�Z(}��u��Z��-�iP���Ȅo5`F�J]!kr3�VE��G�u���L�p� �j�9X��[�Y��3}��-9�b�c���E9Sk7Y5�"޴
����T�|o�^�*���o[6�1sܘي
{�b��V�matE��:���vfɼ�m�'�v�;�c�:�Γ�2L��.&K0�`���n�͂�:W�![�S,�I�\%�\)��w�^�퓲�f^�Y	7Hn��\ޣ�%w(��b_ps!be��*& s���Z��ѵ�Lu�����4���/c�v�b�3���5*3cȠ�����M�rfU�N�}��L|�\��EG�)A��,V�� ������v���HC�a��tഇ��<�bV�Uv+W:���lᑣN@��VJ#�*����c� h��ZA� m���w_+��s��}��:\�����JUxJS5_M�Rɱ�ҥ��|�[�8��\���g�fs��9f����I�{3�P�|&��W�di]+���k�&��x���4�oN�Q+D���H�!�{4(H�uÍO��ŞE�T%��]���A��5�Ƞ�\S]�/v��b�
:��Xn��}0V�:Ň;�m:�V6��*�n�U*����yt֞���cl�M�c����O]i]f5:u`36�"P�T��#��7��X%�G^�q��s�qR=f�fƚ�{�15[�̷OSW]}}�[�/$�P�r.l!	%��мPNG���Un��������GIvL5�O7-.�b��o~�6p�j���b�\N�V��ebH�iPr&R�Vs���5�C��=��sp�;/�M$�9P^{��FW�n�V uU܃̧e��Q��.K<Q��:ڗ,���Yr��&��v7-��x��֦��<�ˍR%X�=.�G��)Y�.8y�QJ���-�Ap�%q�WX�Gy2��9f3Ft���>s��3Y�����nVo�h�i�3�w��: �v,��
�l1���q&9ہVt��Ί�©��Ո�J$N*n����N��N�����,��)6V-�O���b.�����չ���7|��=��3�m��;�:5r�`
q������z늝W�����n� �tDҀ�e/�%�r�|cD2l��Y��K��m��F
�\��|K����*_멂��~�+F<�اɡ���s��K28�gv�!2����c��3꺲��ըwgfc��gKU7����\)=SO3p�>�:���i`��0$\�d������w���E��3�:�(�g����m�d�\u�J�1�,K/���9��w�r����{9!-������Tp��E��س���@u,�8Yk'{U���*�d���c}��^�2LnDAݣZ^$��@ ���Y�����_���]YÛo��㻇q�ҨK�s[�xZ��{MEr�{Q����aiBu�Bkg.��N�Q�d ��Gw�6��ПF#��<y��񮥅��tfm>��t�d�k�aۨJ1A�����vУ>:�3g%�U��E�i#GO��ySe�	\UI���J���;�v�'wj�}���M\���@�]�j�q��*mr�j;�X��ǥ��w�|��r�[��{Z���IRB}x ��t;�X�02��u���k��@6��e���vA�Rs�GZ%�>�X]���9�K��]��^��b΂΄��p�,�؂@��U̺��+&�}ko�h�廅�@e.�d[�WZ�Ũ��w,ik�Zxn���\�x*u��ǋ+�:����,B+�"��8��n5����{���+ku�tv�<V�UֻL,B*V3��"&Da�efN�ӝ��#�.ٛJ�f����a�g���.|��Rw�*񋛖�6�-Ħ�	��n�&]@�N;�^��7���:�]U�h���C�(�.t�0�dt�׈N���*��w)�IM��3�u�EM���o!9Ǝ��9ֶ��:u���pK{L�SX����vo\J�[fvX=Lt\+,� �f����g�m�N�'Q�K8:���|�M��{���+L��4�V5,�uC�.[��l�u�A�V
z�2�k�v�a,X�r�t§
6���у�lW�K�]n�
��0}\��
S�ۢ\+�;}ǃ�9�+0-2*���W�oF
oA��O@L�����+�&$��*&:�w��|�_B�6v9�F�d�b�Yzi}f+"������&<׊���y�/~�1Fr����EX��3��c&v���˧/w��Wc(�_$R����ojm�:�$���Pp����i���q�X�V�x1�)I�Ab��C�+�
+8}A��Z=�F��Bw��d��-��ϵ��`:l-|���@S���)t˔��\^�%�Xv<��)���a��؝��4p�vZ�YrL(��ܤl�Θ=�b�	���G_/���4D�c5K��	I�YRDʭO#�YW���A��91:�6���Ƞ�J��:�x��y�[���T2��s��hO���m���m�]g��[��<��)�x�n�jbUI�:��x]��jI,)(��cz#���2rs`��EBT��V���?�-ƃYaC��A�sF�>]�g겞�β�H�g�)�lٹ%ЎY}�c�l��4�����%�a�z�!t�NcCu��nmol��.���I*I��2���/���7b֨�5���* �]:7�I���.[����g�� �Jh��BƉY�7x����]��&,�0qf�����	�kd�0Y�GL�m�<�ŉF��k��6��9�F�šÂUN���^a.��pn,��cPl=\�ּz��ɣ���9Lk��_SF<�*�۔�zq����E�{���e�}�	Au)�a׹���'%���媺*���vn���=}��k�-��ꖭLq�F�p��� ��TR�T���
}��5o�Q���so����Ȍ�]\���&*�F�ѽ3p>3������Y-��4�gtZ%5�\B�X�j7��tm��AV<���s�Wǜ}�a�C��3���gQ�]4rI78����
�W-H9cG��X��i���	M֗�������;����W-TQ��:��f�Z��}Q�Um��)�B؁|�bɥ���Mފ�����ޫ����K�4yù���恶�iv;�����ˋJz��e����;G
;|�»���;��[t:�����Ù�+�Ko�or?���gf��'+c�p�x�-Q`|
����)y��V� |;SP67j�'v.#or�q*��#-��R�ngZr����"7��2�wF�:��_'#Ѓ۶��,3KDf�9��� �nݕ+	ˎ) �\�6�ō<�dY�R��f��W���m;�O8�;���*�ʹ�x��8�j.Wh�/�t}-�z�ţ��Z1�[W�,���u�gk�Ù:G��RƱ�����jF�k��JDf���]�'r�����)T�,���Q��]�tX����m���c^f�呙7pN���7,�JΝ���ÉJ�C_:����9�\�c�G���gny�[v)[K�"Cn�s�a�6S���s�m�fkl>���ƻ�h���Pefekj�I
��[p]c6V3pm���Pn�5J���ݼU)9d�3�f���x���P�f//^=aN�V�֪�Xd�o�K��a�GaʧA�w+U�+.ˈ��dd;-�%4�u����K�7��>ڸr�C 8ZZ�EO!�{�'|V	)*�H�9H���:>�N���m���A�@��v���f3�Ԥ��L	�p�X�\j]u�x��,s\N�waÐ�Y��q�\�J��ž�kdr[�����{�%�Jt"�}�y�wY{Ռ�a=���z�ܽd�I�O���`�z�(YY,��.�ֆ�*$��mq �G]8{{b�gg�U��G&��-2fJ�[���rq��,�V%0p��Eq��䜱3*�t�:j�B�v���Z&��܆]�s�-�+(̼&;V�1}��mw�wc��Z�,;�@Pr�h�Y2��C��*rs.�3�'s�}�˙"mZ63�EJy�*�$���:�d}�f���d=N��d�ƥ���{��X'2l�Z�]9Zv�V��K;Ճ,,6K���}:H4�R�%c@��A_BƋ�J�x�B�+��P�Nt4�<Y��õt�<�7�t�k�N��6���S,��V���sV��8l��-Se�M�4g��X�����h�������t�8�႖�	2M�}3-V��m��H��0���6�]�tؓ�ܦ�nԭ}��fm]o!D=��`rܶ�gkC��{@=j����n.pJV����=�^.j�k���kR��Y}��%�G>I����PN��˙)�e\�'�+^.��'���B��7��t��p������K��Zp�� 4�Y�v��9���W	��)��]���6-.����+���۳Y]E���aÙ7�-d��Hm= T������g���J��v��6��_��B1՝�/�+$��/���%����K� 01Y��Q�.�|��n,\i��w'|Û�r]�\�PC[�q>���%���q�`��_giök.���P��q��Z�u��5ݚ+�]����02ݵ�qٻ��V���vo)�L7�%�w�}��uv+�L��+�u�S�S>�t��ܖ4Ɇs���}X�{p'o�XK^T�ښ�a���Y�Ѷ��KH�u��gJ�(r.B��Qλ�/�	�4��g����3c�{q����Y��o2FY���v�U��m�i�I(	���`��(_gK�Ùx ���<q��
6��y�>���3�XS��+F��f����e h�p�a�b��8t/�+f��[���5ԳFlԭV�1����Cނ�;����9ck�"�vLC���2�o�
�s ]�:�ѫp�jИ�Ƅs�!�&�#YҌcHg��uhl��_�d�t�F�6_/R�I��NW��W�l��U6^g�Z����mI�EXҟj�����1մ���懽��N��	����\�8��q�o��n�@gWtɪ��3\L�]B�̵y�&�2UY<[����Ii`���҃���>ede*���ʎ�u6-Äm��\��鲀��p=��L���Ǝ�M\ͮW9.̷Zc��:���/f�9"o��ٻΈw0�2�펥o��T_4X����Ll���C7.�K��o\�Ԑ]��V�1W-X�)�-8Q�=�3�3(׾�qc�����tK!�ꧥ��73.��,Ċ�S��P+��|�:V!{�h<<n��U�g����U��(��T��-�>�!�̈��؝��++�u�:m%��V����"M���	lޘlԕ+q�AޜD�1�-a�tIS����S�{6>bN�m+P���3�cA�nl;2�^��>��:��=����8GY�]�WhT�i �Ԅ{y���AJ������Z���p6>֦��R5WA[W�����	N�}p����S�*f[�}�o�Y�FL�ͼ4�\�,�C�s�Gb�f�S������Y�͔����Vvm�D�.G,v�`�U:=9�B��]ܤλ���A|k2��v��K�w.n�*$�9u@�3Y�Ul�`��\��i�t�>���cO]�и:�Z���%���ו�����b�H�4#��ۙ4����u�9�o��]�aJk��1�d�耹^�r��ܙO��mPW�����T,Y�WG#]��� ;��T�a��J�(U�r���FKΫ�߹���8D��Y�Q#��D#����� f�:F�6�s��� ��0@�l��)#�
�����?��_�e������")��kb�@�0��)?~�n:?�!q����
0�Ѣ!�T��@@���ļ��Ȍ?��M��?Y���H����5^�"Ȗ1���G���������o2w�9��r +R?�<�X�����4���ѣ�CUM��B|��?	M�f�!��sۖG���(����2�~D�L�!<`~���lVM'Q����� � ��=��PU2�(#-z��T�Q�|���`_���)�+��m���%?��)��x����浻��Y�Q&�:��*���'��S�m�V��F���.�yY��k"�V��6��)u�N��3�]LF�1aM��u�$�z��t�u�q��vS\��"���Yr��m��ĮPV��]�R�6�d�_BZ�F�A�wCt>]t	��.��4�
����n�����t����Y��u�[���{�j�S}�{a��}I�9FRm�pe���I�qz�X���#���R`wkB�-BU��w1C𺾎U�ؤ��5/C��m�V~�|�ТQ�.��ׯ���-��,��W�Ǳ��ںY����_S�>BI��u�\��˝]Q�7��S��u�0@�S�p��R���Y4��gNl���c��VQ߹�!m�
�x���*fTU%��)����.v��0��	��l�t,�X�%@][w�%��n�m)���8�.?�1tz�Bpa��x�=Nf���݆x�\PPŵut��:��s�h�1@�_m�XQ���l�-\��n]>�p����&�2
�@�+����b�t��N�rņR�N�ծ�IiV0ԝF�M7�=S�]�}��+S�İ�Q��Z�ݗ��,U��q��pv��+Euib%2�=�sm�Z��5n|����_���������ׯ^�}�z��ׯ^�z��ׯ_o^�sׯ^�z���z��ׯ^�z����ׯ^�z�z��^�z��ׯǯ\��ׯ^�}������}�z����=z��ׯ^�~�g�^�z����׮z��׏^�z������ׯ^�z�z��^�z��ׯǯ\��ׯ^���z���ׯ^=z�����������n�竚���e���"Q���j��N���uy�eYS C�j�Z9K.��[˪0��6�%,�/����:��yV7���'(�<s�<u��ut�!;lu4s��+.W�̂�(��tP��SU�[B'f�u8wf�����ǚH�c!�����޷�7�^�/n�i��`Ǯ�sS�2���Gk0�E��<��W��/y��wh��V>�nc��R�@���TI�W�i�@���I�*[}TN�9�T�ܦLZ���*����d#�K�^�Aj'�% �z��qG��L�ܹ�3rμ��@���r���q��_ u��@�w��(L1��G���E]C����l����V_.�m,��i�_h�\3�ʧP�<�aA�w1������67&�u�u��f�哤V�����Gc;�yp�NZw����f��>э�2�
t2_K�չ
в��3k�ra�S�+@k��8�_��y�T������Р�����I�;��BU����N�M�+w�wX�J֮$�ks!���¡W�>w!�Y[F�Ut0Xz����])����Ó\O��"¶E;�iL��;�s;ـֶ\�̄����!��n°rLSS�6 (1|��ͮK�+�;q�F�!ۇ\DƁ-�Wt��ҭ*�B��۲�c愋(UN�3o���ǹ @�W^�}H�׹�GY���������χ������������ׯ^�z��ׯ_oG�^�z��ׯ׬��ׯ^�}�x���ׯ^��z����ׯ^=z��ׯ��^��ׯ^�z�z�랽z�����}��o���^�}=z��ǯ^�z�����=z��ׯ_�G�^�z����׮z��ׯ�^�z����=z��ׯ^�^�g�^�z������ׯ^�z����>�Nţp����:�wTi�׬�v(o[�okf�����ۊ�o60jЙ�SHeV	�\׊�1X��1�Ço����%k���5�A3���6d�>�]Q�k��1j9w ��G� �t�⣤�1Vgfe���]6vv�f2��T��ݜI�ʦ[ܦ���4ľ�}Z�__/��f���TX;ŵ籮��]y���$�� �dZN�r�c:uc1_^�ѴcT�Ըk�k1Z��>��qd�G��tZ�����Ѭ�H�n��&��6^;GN�TMMr�KMc(.��<��փ�U�n��w���f,�g���S�$�t��t��f*���T+2Lou=q��c(�?�<���uq� |F��e��w��!���=�1�<�C�T-3��\J��0�-9�sR��#��tX�P�wzS�j[��<��ïci��J������Q
i�ׇ��e��Ȇ`vQѧzT͊�o$d
X���EB�������?�s�y��b�87%�F:����]����r�s�"f�θ/R����#�x0�nD�n��u[)`���2�8ؽW��-��%.�D�߱� �v����Y��{9�ŐnQ��Ky�<��B�;�s��������i*�Ȼ8j�MJ$i�f3�a�ΐ>�%�7��u�9���d�k��Vg4��
6"c;q%�Q�O�^\p;��P���A_Vlvr���q�j��b�9�5g��V��:�Č��̊�����f�U����ۉT��,!�jJg�<ƘD��[�r�Ģ�I:�܄h�alx�et�`]��Q�+*gIPd�w��]]��.�:g*�X�z�9�hI�3Z�s��9Zw�q|K֯.]�Ր��tfP�/�J$>·-��敟L��S��t��/&a�S鏒b���3� ''j+��R�u��[iu��t�1� �t��h����=--K�ʺ��Ȥ�K�2��A�cr�q��e�t���&�j �����v%��f�Ϻc2��uojp��͘�w]�v�$Ͷ54���V�|֌�U���D��ʽ�X����[��\v����\�\2�Κ6�WU%��l�kfL\M��+��Ծ��"�H7��ZWP7�KG�I��Lgr�u�`�@%��eӁ�Bm�&�i��tKȰm���n��evn���'u.�b�
5��f��6�V�6p
A����1����bU���M�c�o!:��6$��T5�����)7u��.���tB�y���t�M"W,$@���"ړx�ܢ����g,����5��0(��1ZK}�6txť�|�N0%kf�d��r�2��˶�i!$+��Ed��7���I�������p:2�Ch.V����]"4��,�X�X��U�0%�;[SF
�.�"����ʖ����O���Oj�XB)P��S���NJŵ����pI7�܇\�U�㣄�|���k���n\s�h:kkS���N�Kj��q��U�3����@�)�f����\���V�2�����R�>�/R`�b�U)^��0��΍Js�ӺrST�s����'6��'ս�3s��-^:nr?w+g�dH\�����O���%��:N�ï .�9	��l睲�P���j�J��; ��Z���є���ҷ��H&`gV=�T�B��MJUv�)��$/����w�`X��D�|dhb{�+�P�G)���O�X����=u����.e���[�Ϧc�l�-�8JB�@���d��:�"��m.��|��B�tݩ�����^��+����&.PRŉ=��)�]J��νX)�oiWt�g�hU�q�i��c_r�~]��Sq���幕���-;Է�^*�֨s��BAȡ,RW̽q���$�λtZM]$�V����7�B���f��ݪ廊�Y��*N�&���1T��U�"��.c <����c�@5p\])�r����ti�dHS�cp��و�]�]Z��}[&�&
{���X�u)�ǭ�`���\�R����)�׸sq!1�p�t�盗S�ϱ%)���ر[���*[Պ��e&+�jǻ)of� ���E�@[ڌ�]�v���3��ש�f94�b5jc�޹����)�㙥����U��#]���q�����z��9Y�Q���ob+6	Wn�]�.����2c��7���D��}enct����u�[[�̨[][�ި�N�]Q�K�Ga,v�
.�ZS.����!c�Q����K�0�2���f�|��[Y�]��-\`V��V����U��d��/�:@���m��C.>��Hn>�g��� S=�ݸ0�W�+���v�+-�%��+�Y� }�*�XKS���Ix`����[��a2ا���C+�	Du�!����"º{��ͭ�j��h���1���W�4�n�I�]؜�Pݦ���,���U�V��{�Zn��V�V�Ehe�^�_b!���dt��i���]��!h���U�5n�7`/Ꮫd�Yh��r�b|M:;�h`�k���+�!��>2�S�UuZߠ�;uU��hl�Ru$v�1�5��9���w�*Ѩ۵g��i%�t[dd�Վ���e+�r�����~��V�r##F�$�����"�1��!6�n�d�ֽ�;�\�㲗W�X�m����V�WO��g2w��Wٱ�vim#S������}�MX�ذ M���9(�T� 7Z*J�0c�Z�C����{�V�e	��@�+�uΰf��.7�uvfHk��L�Be���Q�~XK�G�K��
��uv%ON����%��W6�mЌ1ռ�9��X�-��ó,�ò8+x��;���o���2IL�f_�>}��T�	�fm���V	�Tw��<��Ӕ�.V�S�F�bY�n�i��,m�V�vLl��>�շhG�J�w$6-[e�[�fP3�P<�d}%�7����x
�*��|j�H�x���E@���$�=��S�20��=4u��q��j�`T�����ZJ¯H&��k��.��f<f��+8�5�q�Zy0V��P���A�Mmɳ)+�ST�y������#�qTwV]�d`�V��^��<������X��x�Ϻ�-4Q�䇻D�//j�U�˟N祭�f'��.Yږ�&e=J���+�կ;J�\$94V��#�+��Ir���/\��Du�m
ꛇ�5��f�W�j-u�Ys�쮨�9�+d��æ���m�*�ޘ�X������T���<tYQDD��2(wCO�^ӏ�T7�lGI���B7to:��vK؎�v-�4�����ӽ�X�/��0�)��r�[�;�t��b��|�
��ݽ��΍B��<Z"�dӫ2-e*�"7i(%ԃ��c����6V���+�q����Iۦ�*�E�
���y�����sk��O� ǜ(��㒇�bl�0�C]��utҪc�.)Iv��Sj�5{r�;IH��x�m*��U�|T�{]���6�Nn�>��YWz���v"��K���!�L����]�Su�뙍G"}vM����b���8z7���z̼P=�{IKl�wD���js�C��.��n$�mҖ�<=�kiMt�ɂ�aԱ ���Y�-����G2U��l=�]��	��m�%�ׄ|{����s�%�!�7��ǲ��%)�d7�;���m����h�{ɑs��ί�4{�ޙ3q�n�gT����x&k�v����hb���C��ʹ�;�3@ò��OS�K泖X��C����B#ϯ��M��2=�v�hrfIXg&:�9�pV�e����ɲ�5�xv�u��yʈ��\�N�έ�U���s��|t]�aВ�YR�Nm��i�+vdDyU�&�M��6��`��	r�̮!e��G��ck�콥%��[��]"ԂF��}���8���u
x�^��(v�|�F���^ښms�V?�p3ovc|^�yPsM]fC(+B�ńH�Ƙ���V�XֹN�48�t�Y����q���/��FE8�<$-he��؊�éU.Q��a�8�9�Pf��p:�;Z7�,�ڼ�pB�;���v&�f�c��_w�ֻ��@�kp"o�����2�xщXĬ(�z�f�wВvޙ��x(��O]��';���:���B����s{lWs��k�W�ʋ�U([��<��Ct��e'���y�d���kt��Xu����|	���	��9aX�¹�=g92�,�N�sqQ�Ĩ��A�gʦ+�[��,�b����x�*`	�n_��6���&�V<쥝��#%�5�}P��mĲ�U�n>��tͣxi��VӎUi��p�I��e�z2$솠ִeٝe�K���#m��I��&��;���Yj�]m,SB��^s��b�Ɗ�[�������ֹ]ԧ�L5a��<ܸD;�ϛ��y5ֈ�-��֜�Wo�;sG6��݌��6�.d�\�;ԸSMZ� ��E��k�g	�7�+�Kl=����kWCz)�6���!��?��n^�^@4*`�3�U��Sc�cx�L4���LL#2~U���%���3^6�Z�:���TGnVTUleg�74h�@Dw�\N�1��r�c�8��:���oWS�6	R��c�q7x��7�5���S4�hn2�b��q�Dj�x#�Ŷs����:�5 ��L��
@�r^�d�ov�;�mw	�ޫ��"վ���0��Xq���P��`��6aJڻ�� �]cuHL���6�]�8D�hP�Z�� }o��?���^�����6�nb�2Գ��}J�Bh�f�ܻ���-���r�Ip�p囉�r�ֳ hT�9�x*�a��C�u�t�����%^d�� �W�d��J�7[>�5���c�f�#�Ve:��'>�O��[��|��<u֖�؛��[Y1�؃�:%G�BS}o05�E]|*�G+��hi;@Q��o<+Ṁ���V�=�z�X�ܑ��Tnu�c���w�N�ޫR⡸YV2F{3)h%v��*Q��5�Ax�XΝgJ/	�O2T��c0�RR�kU��:����?K宭�|Iu����n�c�<8��+� ȆT뫍���=��k�v����ᶻ^��3B��`����J�+`!s1̦3�u8�WZt���HG����w�՛����u��m�J� G)u���sO7�K0Wq/9ɛӔje�:u�@Z�u��k+UtIi9Ɠ�z�^�ݾVB9lPܕaȷ�y��9vqt�ۣ�(�R$徨)�q�o\&^ǇB16�I5f�{���Sn5t��;scڪ�t����Ψtl�� l�
Ζ
$7�EwmL�.�əQ�ߌ�����B��J��@����iIGĖ��[��k�Ca�����HZi=�i6{O`�ݛ/t	s�rK8�ʹa�ws])fŖ���ƞ-����RP�s�zK��MJo`��p}���W�}_R�+� ;;��s���v�q�1��x��uI��#���	��-"$Ii�N�2)�T��q������$�B9�n�i2�"4I�Dd"������p�,���p���6du7�*B�1������5�ɲ�����ţ׹ׇ��i����7��T͸�����gK��#JY�C2��az����k$�27��M�J]�gp�����bf�Ȩ�V�م��\���ZC�n���s����9�J��5@�B(�<����;>ޑZd�k-n's�\���el�X���E�8xeX]d,K ��P�j�s׭J�ZN���P4�e$�e�ܤ����x�7��k ao^P��L	�Ƿ���Lh�,e�:��"6���qgmw m�a�׏K�]Ҽ�>[���c
'gN�>EgJ���@v0dP���m
]vm	�C�֋[�7U�F�c�/3��vx���3�q@\w��nR�h��HfN����gF�6�9�G�T���el)�:z����!W��@��f�����.|f�X�)�}��j;ފ�g#��jv)l%|���������,Ie^
�rǲԡ�%���[��XP���6��ww��!�j� )�н���o٦>dQ�˕0���ea؞��<��R�������]�T��nʜ��ۘ*��1,�;�)6��i�'������0�)��\�z�B[7A���j\�Y�zN*�W�\Oy.s�McTSaL�+0���t8gv�.n5{���뷵�Z�k1T���6^�Q��}w��`��X��H$UQ�ډ""b��$2�^U�U!�1����E�c���鎈��%�h�ۍ�PE�p�6���B2dLĤ	@��lmT1PD#"a]~�Pa��m
���m0$2�ڈ�ˈ�O�a$4d)0Rem�D$�!6��0u��b8�n8P
�m0�($C���]��ׯ~y{7���~��4>��k�bb�ն�*�m�����c%�+9�����}��������}����(�bR8X��I��`��d�����4I�ш���l��+X*(�Z�9r�D���>�o_������~?�Y�J�J��i�C�s$F�UF�c�ED_y�1CZ4m�h�(��]* �X���F-�1�b���8��m���$�gTDQNΫN*��� ����19��'mSí��&���mN�� �j����t��Q�lU6�"
���l�[m���M�L[m��\�LE�����"�(�ήz�"*���y�p�Z"j�v�SO�s�ًZ��mX�/��cy���[b�lz�<\��9m���E|��n6�\-mˇ��^r����"�mcA������9��1�ܞp�+��ڢ�ع��ÉF���l��ƚb3��q1z�rة��l�IF���6ǖ!9mX���s��k!c[W7:[\���Dj٣Z)*�m���[�q��9��Mr��5��nb(���M��ŧnQ��j�1�F���YP&I����d/��f~@��/�΋6�=ѝ��@��N؝�
:X�hmI��q7%�z�>O]���/g:��K�N[Ӯ`�u�W#��]]��L��H�D�0Y �q��E�!l���e0K'�� PU9�ڏ��U�la_b��l�j�J�uW��v~Ot`�/��i�2�-h��)=��hn.�n��� k�n�� � ����[ώ���U�z;Cg�W�9�`�R �ܘ�"��G c�ݬ�w�2<��ݡ����]Mv�L�xx��dyyO�U��?q0|C@��of�<G<����/,��V@���[<9�Rƪ�G�%YR�E��2Sϵ�x����Ͳi{�zLמ�sb��������4�܀�㢼 �����j���W���K��˝�R����g��zY;�0>5��?zO&��)�Yt�]yl/ko�Er��l+H�;�ݞ��(��>wz �隫�V�L������o�yAB/}tG�S��Fo�H�8��zMͪ>y�5��y�"�
��&��>^��J>Kռ���֮st���c�q�z{\7u�,8׋P��.Rڸ���{ ���!	��9�@��)�=��p�>�o/�4����~���ΛP�We�`����[/�ݵN 7*�"���2gv��ہ,)5�=��֝|Ӯ��_`$�|��r�� &so	
q�ݙ_�K�M�H��&jۥN��gΌ����ʶ�����c�]�wD5���q����:H�>��2ǫ�WzǷ�s������=��x�/ϫ�v;���8g�J\��EW��}Z�{2�T��5���+~����o��R��ҳ��f��zl�4�4Uё�O!�ϞB��N�x��Ŀw=ߜ~�o����[�wC����>�{�g=eMa��^�n��]?�}CK펛&�����d�4L���/��^A��{n��TJ�Rsnz���N�辔�_˸�)�1�8z�Ы����q�`�n���F��T*�Xĵ��.`��8�=�	��zn��<؋�{�����N��鞞�E�����T��]&��W },_{�t��r��)ek����t����ɳCWֲ�i4���ufmZ��m�G@Uu�XB��������$�Pq:�!��&��Cv��S]?^Q��yI̶�� (���m�mB�e��@3������ǋ��ѝ�^���~EQQ�,������ӵM5z6v����[�2��}��wsZ"U��Jج6D��5�o�lVl��-�Wy�GM�� ݙ���C�5|���X��_zm	N��Qe��;<Ƿ�y��ͩ�]t����	G7�-Kgc�az�
?T��f�"��F��t�z�����۬�_ޟk���^}竐+w�x��5��0#�V�,���c��P��r�f���kP�\��~��S�����+aqϵ�[ϗ��]R�ezZ�uv���W�Rh�$�s��]��^y�����ջ�N��y���=�2��Nm��^��{��멃M����r�H�TeSA���C�1ʏ�}�|o�*2�̭������t}��~�	O��R'0��;=%x��`��l�m�^�+����3y{�j�z�!8;��⬼^�ۚ�{<����࿦N��{P�^�YO��wE>���O0�;�������0��H��W=��
��Ս�d�g�9ry5�����،���w�f��>?e+�ܢ��6k�͇�h��k]��"H�qVG[����u���SP�E\?��3Ӹ_x��;���]�*�	ѷ:sE�E�+\ލ4�����pȲ��$j�1�lr�~�y������z�z��d�xz��`h��W����4m���[�r�n����(�x4�4,�&:0�\��}n���Nr{�}�-{�Eo�3Խ�+GݲI1�x=�v��T�P�?�f�EDe?u�����K�K��纝��!�Dy��"�Z3d�`s�4g���d��
��kC�^���Vή��z쾌��l�h�8��L��Y�_��'���_�b���ϴ��Ͻ��73Y�ޞ<��<o��f�3z��L�/臻��o�!~�2�-}�}u�ux� {R����4�A�w#+�Ճ�.�gVq��$�Q��1��,3���n���y�h���$�w&�=�s+g�m	9�\~S�^/~5��Kڷ��=b4g1�G9+1�����=�����Q~�߯����T�3�{7��$z��ۆ��*ʨbF���#i�8����M���R��v�h��%��Z
���*���ZW����HӪΊ��������ioc������S(�.����z됮�9��N~��36�8��y'v�z�
u�Nମ�+	��=F`����$JIJRjf�a}'JOZNq������S��-j��������fη�Q����6��ǵ;�^��)�������rU�9Q^��~�S������G-���ތ�8�)�3蠟���^ >R�k��Ֆ$���y��<r$�m5���Fm�������U�ח<͎�+k��{�q�Րךl��w��0�����oV<w�P��z����j��Z�Yc����2�<�G��;��*��͓�r��~�I2l�1�*>DՉ�����=�5���=E�t�=Q�1^$H��\{ ��O3����ck�������^�o�c�r���y�3�.|��֎[ٮI۷����--<N�j�|��P��<睢��v�u.Y�HOL��=�|v�/9��ݱf绘�3��<N��g[gözC ׫�מ�/r�U�1���V�u�-��j�^x'B�0hȨ��z`�9N���农�x�C:�ͣ@��ٙ�Q��T\uV<�qF��+�	��YIo%�b滰v��ڎ�쩴�м����˖p�c2v����1�>�˘\�<*�,�EW_Lfr�-�'�����{<��Uo���y�߰�Ì���4Ʒ�}t�"�\�����z��{�u�u3!��9�7�̇͟s�Ћ�no�.�S���󝈏1�a��WM3Y�Ƒ��"��?l�����yw�t?9箋��}�̊�D���7��#z��8ʏM�}'���{:m����'��7O۱y�>=������88�k�g�*�_8�3����OI�۱3�}��,c'�m�tO��3��9��g�tYg��x�:���s*ܔI��gw��k�ǅoic�S�@1l��ʹ+�	.�{}����ՏP^o��i8n���;}���E<�����t�z���ũ&��j{,�1���w��7X�FP�#���x�^q�A�a�~�9��`�����A�)�[ȵ��6M���oIW2+{+c:�3D`m�Z���P��wp�D�*{�FE�z�B�Re^�z)�����t*P8P�Zu�k�`��*S��y�.�=�3:��J�ڰ���,���t�ٷnu.���57/vK+�Ba��l��vD5�H�W+�an7Wu�N��og5=/%��^�8=^�Rj�u*��U��؊ d_�nr�'oV�=\�n��5Z>��|����׬y[WEU��=��8RY/��Z�>�h�%�=�:X�c���2x����Nd>��j%�}yC˪����m���y����g�5��=������}_Z�����z���ν�G1����:Pͮ���aS�����T������\{;T��l�%�}r�����?�f7{o��Vo������e��C�^j��sɔ������iu����B�������{�Ut�œyo]��Y�8�H����w�����X���te��g��v��g��a���̫/.9�Kݴ���\F���n�κ�W�c/_�3s�W!��`�Ï�+ݟV�����\��Lf:�@�#���9=�6FG�v휙���8��ƈiu�N�137W)�2��L\��h޾{�r�F뫆�&�Q�R3���ł���h�82C����s�\��U�FR�)�<Es���q�)?�q[VE�y%{�W_t:b��a���=�:n����;|�c��9rF��Uv�2���U��1�y��y�WD_�he�F�ԹU��&q�)�F����|��&k�H�6u{�جr/�5�͌�{�Tz�jv��$E{�o;}*��Z෇�j<���9Q�Ȁ<�Ɩ߱��W�yP�&�j�?�CYN�BM���y^靏����Z�����������*��](y�=H.�'�(5�-�Μ䓫����UJ��ɳ���2MY2k��L��Ͱ:�́V�x�C^v璾��OX� תz`�b���i&�����Lq�|���;�]�
�6�y߹2����+~��Puz��
{�z�'�V���g
f�r���\9\�Ht�Ńt?;:�[}[���!4����!�0fٹ�ئ�w)���L�v�������<Ù=��Q�-8s.��g��yV&gt�0:C��Ldtxo<(KYCt˔ȅ%4e�S~�������^�%���㭣��>ei�>���\9��u���sMJÖS�[�A�:�LQ��
��]��ӘV�T�3"\���������bf�L��d���*S=�<��^����[u�~p�N��={�*У�2yj�{��=���|����b�g�����耭��n�d��ۺt$�d�.d�|$����jzMߠ����m��ÃHf/�V����������~g����=��c8|/u������+ɵr�I*�7U�x���"����W�8����s/���vܡ�Įh3������y�U�5O@��_�ZS�F�~���hS yZ�n����{�&w7������0���}�,��}�2�U>�Oz����w��+�6���=[ϻ����}W�D��� �,��0 Uѝt��Վ�ܝA���W\5>}���P�X��*��1�-��^�nES��Ow��^1�н����9����gʱg���v26u�O��$�,ɣ;�ѴNA�V2�e�%�GU����Y�����	�T	9���n;�R�7U��{-�a��ryd��#��c����:F/sL�)c.��:.Wp�Gt���@nk�|�ll��zL�	��v[�q�r
���fK9����*
��h���J�8�0)����Zta��o��{������{�ǥ�xb\��۔T����{�f�c��d=t�?*g�=R�W�=���k�q�y�S7��\��!���^}<�f{�������G�!YR�>�[����ͳ���{8o�g�Z=F�\t�8X3���5t�Yz�]]Mi���rg7}C�;�����ϫ���4v�L��|�#)�r�K�7C�I q���u�*e�s9�xS2�E�Nz�nf��ro{�irn��0fv�������<����0>1�zDF\���9�{Nߤ�TN��bAw{2K���D����ww�i��y����%�z���-u_����{��;�q�)�XW�ڈԀu�h�������-����{H�YjIc�{Ɍt�6��Dv
���n@�m!��3��<���
=N��qw7��Lv-g|q���p���S��ʞS��ѷ~�Bb��Y���rgN�s}P�w�9����2[2 �����]�z%PCWǁI!�.��ʵ����r��Lk�����j���i��{+y�cJ��f�1ެqё�P�w&G|�R�'m�Z6@�v�ƕ���J�P��y�j�̭�
t偘Jõ�~=ekU�aL��L����m{��k،ݽ���9y�,��Tx�ٻ��r�k*X���j�Qݻ�����o"�:��ʩ9(a޽���)pm��y�v�t���L4u�>����+e]�� �����ؕ]���w�9�fHWdk��:�.=�����}O�V�-�5���:�(����i��h+����w`���:�;���l��V������ꘚ�w-9�u��%�q*�!d{V�)�{�p���:�B�irtZ/k;�N�MV��w��S���M��#n������!����:��b脙�]^sӐ����l��+�u񚱫u����"�P	QN��W�r���6�e.]��X��l�$�=��*_��MRZ�9{A�б�����ʝ�QU�a��CF�iT�V��%)`yW��V�#64�lz닮���5����9���R�k�[�ޭw���ULO�ɴ�7�Ƀbo�룳�*!�E2��&��
�4�2�e�F��Y�:P6��*E�!w�Ů9�n2��Hy��Y��D��`��l��&ud-�ݘH�̚�WG)C�Ë���JO��?�P�3c=�U׹�$�s8�9Wj��A]Jژ�U��U̖��m�O]��ʎE�3��r^Q�����Ӆwl�[D��p�V�ƫ�
�gw�luK�x���ec�t:ý� 爌.l8g��uwu�p�P;&�9J#Ϸ��KT+ }�Y��jڏ��N��]q.��\�R���.�&��?��}�C��pŚ�)��0%�vt�t��6��3 R�qb��2����\1m!��[2鍶y^lWa�#I|�o*d����&=8;�E�^S�4հ��u��W3�K*T�2�hP c��#����)����b���B΃\��J냖<�����-�;�-�=�F��;6�q_��a��@*3oZv�z��|��r����Q��z�<w�q_f���{�F��S�<��*<��
�ٮ��9�uj���:(��e�{�X~"�D��]޷V�wk���P���j�	\�O�ޠ��i�c`i�)g^:X�Xǣt4���3ae,��CD��t����vY���p� ���:���|�@J��O1u��3N<�����ʊ�ݶu���h��\z�0���N��4;0�:�,g���L�!r�{6��ʂ�R"��/n�_,�o ��<b<81���ҵk܈�Ʃ��ځ$���cm��c*�Ϸg&��s^���R�����/��-�� �j�Nsujۜ8�\�&�i�Tk��m~܊��m�8�Q4��V�� �?������~?�����?��?���rڌU:��<.D�v���G�9���1��fu۞`�W��k�v�Z9��j���4M{܎3������x�}��o����x��X�f����Km�Z��v�\����`�T�x�3�>F�/6����n\�ִW9�Fϛǘ51���h�Ey�sZƏ.[j�����j���� ���E~�������gEQ�\�`���`򉼱U^l�i��i��HH���X�^���)����'UU<�G'y�1��Z.mPI�\�Ey�E^l�>cTr~�8-�UTE6�k�5��lh�#g�؋m:rT�m����6F�ѵ�*"��mmTyi��ѣ�ry��sMRV��6kh������8p���U4�%h4�j�F��a�PPE�kl�F�DkQV�2s�գ˄�6�IAL��A���ۛ�D�G,E4�T�1D4L�탖�~�=��,�U��+�������x�
��Y���V���%]�L������+��16��9�<T˫�k�g
����x���և�H��zb��=.�ս!��ͬa;�HzZ<�	�-��ױՑ,�������<V^a�����C!C
�|�s�W��8� ��Q2�!aԖPB��Nz#�(���9f���h�4����Wq��W����,R�1���Й��\���y�ױ���S6�����_p)K?O,���]�.3q!���0��t��Ӂ�o0�p�����^bఢ�u��QCӼD���7�Pn�����C��!��q�5�g����y�����������{C�ȃ�m�3^��]��f�AB):��h������J �qID�/e)�VMm��o��E�C����<���<��ٛ�����6us�=�邁dH�"�O8�]'�b%9�R)��&��ny�ϑp���e_"�fM(��{5�n__���q��mBc����"�@.�w��]'�b)9Y�h[�[\�y�>�^��#{զ����q��XAG�9ͷ~���l�.y�=�
�i��M���-?,O ��tgne�7�n}�!��xSL$��4w�&���/B�C�N�xmt�u�8�YlOE�}�Ó�.�BE�O�=]�U��vV��7����r�ĩ�dQۦ�ǐ�����g� ��o����i�9��:���歋c��;f��qF5���Z[�WT\ ܷ��t0�x�[u7m����@�.���o`r�,�>*�}>�Ž��oޯw8��tzz/���%ݠlc �#�c��O��y��}�t�(���<՝_t�̊�M��{;����=��|	�O4+ ��@H2��1����'����E�Cm���&�W!���P����K��5�=���i��K����C�H�`�4?3�fY��wP�:�,�==.C��ӷ�8ȽK��H�4#j�Z�qV�Y�:���sP/�����E�b��G=���ػ��P\2
?X��"c�́01��f�}y���Bk��Eڇv-���!s[�$���z�<��{e�����g�c�@cm�N?�_O�a�u��WF��͔��|��m��f�j�]�Q1�{z=�=.���_y��@l�w���P|aoql�ؚ��u��ֱ\M���5�?)�LN��=�͇���nb�mHγ�͜eY��Ϲ������y��zaL��j��3+*��-�jv*�'!>7�%C�d	b�+���|l��s��3 ��Un�;2�O+��o{����|#��k��FF�� �@��^%B��U yŵ���>r������2��yl/���Z�
�z����)|�����*��Y��z^�ء�U�t�a��w�b�㚺�p��0i�x��οQ�/a��zlܭ[�c�G�"SMt��[��]����n�o1���Gu}s��;��DmM8�p������9��pƊJ�)���6�S�M3��i�<}��= t^��� ^�77��s7:d]�Nl�Bҙ-�¦i�k�4������/@��Cۏll[A1��� cH�(8�rMl�pk��3�oR��<�LW>�[w9W�*u��E�]Ryo8<�{��b�z�o'�Gm
�����!�O���z�˽|hfG���p�r'aU��7^t�77���ع��t��=;�?<�m?�בCw=/)�����{4��T��T<g��W�J熵P�����W��g�&�w�b ��!|@�H?��gVu�{;_<4�_��8��<ه�[
���f�J�������k�[��@��A��/�o�[���;��!a�2oK0����[/zE-d�d�t�=+��A/mr���+�hN��ٞ�a7��nk�<ZC��y�~�8$<'0�~t�{E���e�{�ӛ��x�s-+�7�v��C�^Yi�|��+z~�'���)�����Z�]q�$�6��;d�?��hf"6�57��=U�x��:a�q�˱��Ž�rW��O���Ht��ʚ� 0���������K�Ef��5кF�[�q�*�w�r�\�JL;�X4�ʕz�:���o\��0��^���V�Z���p�������4 �4ȸe@����mN�o��d�w]��κwk���6̂�����;�t����oA�Do7fI#�]�!��'������HG�A�ʄ�չ�zY�`���I�w���O}v���ىV��{p�d�^��Ƕ�3�Zo ��4�vA�W�-��J|�.2ߩ�t�ê��#�x�m����Mz�!�X!A�Hw4��
W9R��)^���\�O��� �r��0��Nj鰹���G+2���<q���gopmlk&L8�s���N��~{�"SoT!��b�I֬vRzv-��R�g_G�({�n|)i��ƚxk�=��x��=!@��B`$�i���G6��	L�Tc��3J���w�]�{��? �y�PS�*�3#�5�s�'ʀ�� ��c�}�[Q��)|�mg:݊yn�w՚ܢ�J�`y�{_�<2.����L �>�s�{����cZ$f��`���hJ��6�����ӻ�x�+��V�up,��*�]`�c��ۻ�9�LY�6�4���/,�&�dא]�j�|�~C�ٵ�h�l8�9��B��R�Bʮ������9o}����@h}~E��P�U�u�u��<���a	��~-�& ���C�����.��0���i��T;�8l��ڶ��#�ѹZ��^-��Ս����8D\��a5������} 5�+�U"2�D2N���t2�����V4�ʛw��:ی�b��]L}��2q��.�3�5��4���MrL��u�1fϕh�5q�m��:�3������Q��b�t�o�E7�V ����zG�s���]_���TZ�93�7�J׷�m���1����vZp������z.Yu,�^�?g�~ØLx>�4u|g�'mJΖ~;���*5�z�i��KĞ�=�bX�2���*}8�\m3�if5���@f~�>:!������w�����e7�q86�>�<Xw�/�;�jJ~�1�/\Zeb��l{�ob��K� �-ڰu�4�D���ZҦ{��pg��;*�K^9[����8�y�Ŝp�ن%�[�k����מsBj�aݭ#��R֖t xa����h=�9�+�oP�3s�L�vH�PK(!C��p��\���h]�fo�S߯>���e��Y��)�`c02��`�7����z�1�o��m�[(05����lN9\�vP���{���2ݵ���8^�������a�����˾?���*�a�e��x���*�lKVZ|\݃o��!��G{\��X-)��>��E{��j�?*ߘ��ٚA�a�"Aڧy���8U���h�0y�NRj
3�BqbTK"�R�ebT��k�Dn>5{��gO>��xe�\e�be�x��C��a���S^4A��L�3��4���D���#l����Wc[zsF�t��:���=rԸ,�):a��Ʌn-���|��1��q����$�y�쮧�̜�g095��$/��V��HM��%��og^E
�k]��뷺��qQ7��}�c�������a$=�������^��2����]'��NoڤS"������ȸu�L�o2a��e5�>�r��1� A��jc�)��`��K���F�p��+Z����ǇKۣCB[
����N4<��ba�y�4[q�k^"U??�05Ƚ�`(��]6��z/������ޚ��aB�8+J�qV���ׇ_�Q�����B>zc^�i���eQ���w��T]ß߻��%�;���_�ӭW����$;ɤk^*uА��O�����k^0���9EQ�x��sE�[R0[ɵ��d�́J}U21�Cc�p��[��#�?7�M[&����5fC�6��h|�B]��"���P�Xc�kعH�������h/�:�G���/G^f�⹹tj���!��zb�6'�K�p2}z�F�Τ��K,�dq��oP1�ܳ�蚗��gy�{��m�7���oC	gg������9遌�xf�}y��^\f��{���a��
nn_����������E������[�`B�F!�[�~���\ŶS�͟@���	Q���F�cG�J�_l�c/���v�iސG����]�����1R�s�RS
�"��7٫��=Z�#�n5Mt��ÈC�8�?T���h�f9�v��/W8�WU�e��d��c�.���(mWR<��v�̤��"��8��jtU{��xN��nf�������o�;�M+:��_X3Rzi��4���������d��R��z#-��U����C`��<�~����?��s/�К�V'�(s��A�9ԇ��2L�P972W6�gY��3cP�Ξy�����|��\��|Bʻ��״���X!r;�NE���O�q�.�@�-�1�Lu�S�ʋ�4.<��FS�ڭUg���k3�nC�-��x��'P����5FB箈N�c�(���xQ�Te�3��ƩaD�?���}˘������\s;>#����B?�F�O���x���I<�)͂�xZH���gU�2pV�ͺ}����=���|�j�>��<6� ��2��bޙv��J�L�G=Hg��B7�z�f{��k��"��k�ߠ͗����F�xBF4�r�	�H#����	ea��CA�����$x��S��hͲoY��!���E׏Ms�^�s?;��-y�!��zT�5�_4�U�c?V�,��zuP����xUY��V�Qy���X�=P���1���e~[S���C���o��y���u!�K�F�C�ׅ�s'\]���­t� f�Wդ|M��1�B8Q�<�{��5Mg|�\;\���^\��cC�^r\�j���Ӊ�s�Cs� �_A���t�F�C.�Y�[�|&L����0��[0�Xz�f�B��	�ƺ�6TO$km�i�]��s�@B-Lq��j���S������Kӥ�Q�^�����ǼC�&pĮ{�0`>���!��M"�c5��jÙ,=�8���A/m	������]����~7����D�ǰ��
B<��!�����L3,���-�^�J��Q5��1�b��xuU9c �W�K���@RőqE��c90!�Ń�:`��O�0̓���Z����(�Nj:�=v����{S���4{��9�{C���,�)�$�@������-��gm��r�ޝ�TP�/-س��E�Yy���I���f~�g���Zgլ��8���g�>R�uhB ��d<�\!���	��{l����D<�vA��{$!\�y�\kz�5���Nfʩܳ5��O����=u=�́pϿ~���8-� v��qa�;@�R�~{\�.{̈́W�e
6�<���r7�'_
�ϕd��g��V�w��E?!��!�\8�y�c+v���t)��)	��5ݿ&�齂1K�1�<z=r�2�h]�L�X��4l�~vg�O,h|�_W�i��j~�GJmkȬܧU�hx�m���u�Ҕ�2��V�ټz���Ukb,�����Wg����y�vJ���(��Y��؎��+�?َ s�Q�E�����ט����ࡹٴ��,�>�����=:��]]�u����|��Π��k�����\�V��S����]3#����+P��w�Dfe6����������?�{���;��ӜX��Ix>�}���tY�9C�)�FS/1��.|Ϸ����#a�*��l1I,������Cš�s�Cj��"z�}I�}}]0�U(��Ͼ�cz�;NZ��m~��=2�i�Tڳ���\G��)Ŧ�n�0t�/�pQ��*ʞ��Qi��$�)���1^�k�&:�j3sͶ1���}g��H���Y���20>OW����<a�_;�Jt^��F���p���vr���ٷ��x�\`&S��� ��,:=k�<6,�Z=n�&��4�C
���{=6���N�B/r�)G4���;\�Ӡ ��A��~�:�3�pͶ�<&9��̙eݍ�y�<LF�BW�ˢ���v������y��>�	�;�0DH!''CVh��StV�c�Τ=�R�n��>ȼ�헰��1�/\Ze�:"ص�Ǟ�N�tpsIU��v6���z�>0^��n$<I�/���ұ�A�}�X�w���Š�'�����OEiH5FZ-�fC�aϱ�g��qf�c�5g�Nw����i���;�ﾸ<0��9n�˜��b����&Pה������Uc�O���s����ôe�O��lR����H�B��w{�[ko,�-K�5h�p		A@��J��gz�9��Cp��LT0����t8v�Y�LL���*X�͝�Ϋ�k�������Ǉ��+�Z��aH{���=�V?޾�ǆ�k�<`|a��x�W��.���М�T��1������Cl���xy�l1��$:͜OC��P"��`qm{pZNu�1�1��%���eWn�*��#�K�g�ЌlA)A�U�4�®�1��ǯ[ռ��FC�
Έ��f�]��B�c���ѕ�{XA�G
�5���'�s���ebQ��q����t϶�%:����_:r�qy|�����NS�eLk _	O���z�N��1���SMmq�<��~<k����99Wx~�T��-�B��0�}О����K0S�}%�H�i'�b)9\�$�}ZK���';���������}l)#�C�lLpm����na1��\1���
NM�Η�Hx��p������:��=[\9����F�Ñ���k�v�y�0'��^y�2K����b�0y�l�&;��|w&%ݢ6aD|5�j?�?.���Yc�ͺ�*yD����DÕ9"�(A5mv7���FM��)� �����n�ۮ��n`��=�x �aj�G�m��g�Ͱ�V�_c;uB�WZ�F.Ͷ���$rp<p
[�����`/dN\7j�9+$��\gK Ja❇�@^�c��g-%C�/�j}�\�J��N�cV������	Э���0�p
kͽ����'t)֩4�����Lj�s�wr/��r�ب��T��*C0sv�dl-��e�O�������5l�8Vs��(H�٬wj���L�M�6�;�0ּu6�<Ii�9n��ٻ����֎Ֆ ������N��Eq��v̸nh���lx+���'���%�����m��X�����c"�Z[�:y���Ki69�6�p����H��Շ�v}��ъƼ&�ۣa-.nb�]dJ�6���a����x��Σ�{l�r��;�x�ft$*�[D��W�U��7.�f ��FҧieAnA��.���f��ͱZ!	�8�%��/�=�n�{�]u��k2�4��P��fF�;|�pNʋ�.�6湶�%{ڶ � �geT
�}�!��^b7��y��Rtm��0b�ُ%�rv��]�Lff��1d|����Z���_�����ʒA���f�]Cf��Lݹ��:Y�9�[U�f�<=.3�aCQY��v`�cW�--ř��cgoEܮ�6��\H���p��i�udMf���3�P��r��U��u,
칰0j;�$�ta�/WK��� F���Z�RNoM�J�f�ROwB�$m�L�������%V�>4�@俱�������4V��~ᢠ��o˰�~����t�t�����=(j��N�%{;U�1-D��%�ޱW	��wPe�w�Y�T�=t`\����wW)�R���Ӯ�`�ֆ��I�P��e@��,�)3>PQ�%[��vN�ݡ�E�.�$��!ڙ�.��W0�]���[+i�M��/_Sd��#mi���:��\-�c�^�޻ar}�A�jJ_:��źl��c�mNׄʳ]�G,/-��L�!n�,O:���n7X���Jab��)�ٖ_��/��wA�a��Γw%^�EV���P�42����g�� Vb*}i��	rD��B�i���g+�O����,K�1�G��moi]�6>z�����JW O�mc�v�ņ�F����Y5��ǲu��=V])���8��"�8��RPP
�Z̹	���f�Y�|c���Rg�K]�]�%zE]���{��M��}��)3��� v��Z���r��E�t���Da`Io���1���Ҿ�%+��-;Q���T؂yHc����8�y��.u���
���j;S�O1t�i�;L�ؤWs�9�:��i��k���5c��'\��8� ;��3�64�r6�=Ock����fVc�rd����tJkMhz���*h:�i���Q��X:��D-�T%vj�Y/�'Sw�!��쳏a�K���������g�=��f)��h�����S��QA�9���>�*�m
��N��9Ϗ������~�_��������_--7v��&*��&�&j���������TQ�4zg>=}�޽~?�������~�����TAv�mZ&����4�snZd�媪*��8kZ����>6�<�"�"�����I����!�1�Ӣ����ŭh���&����j�*t8�j
"
��;��j"���)�`�3MQ>Zy�*���)�"*bւb ��j������� ����Q-4�U1Q'�fi��Q�媂�h�F��|�(+�4QW-��4 ���i"����B&夂�����*
*&����(�f}h��AQmDSUUDG69&*�`�c1�
�*�tD�Us%�j
�����b*�&���"(���lsb�gm�*�(�J*"�ovH�$��k��*�� �������hh�����p�so7�o/6�l�T�3��t�Lz�?�j�wR�ę �lԹ4�[��`2�#^c�2�_<�[�a謍�`[�Ձ�}��vR��%�-�,8�6��d��.Bˀ�$5��
x���9���~s�����}�|�o;��*@R�J�>z��G�>U�e��W�`���6]cǳ��G�l�sI}����ܵu�!kﱯI�gwc�<A?�P���,Z}ͅ�>`�4#s�'�3L+�h��+�!��Lq~]�{s ���Z����� ���D��6&2U�A�*/m��5��|ɥ��g��?o�������@(�}(�ê�
�V �l.9�&u~���sy���Cr�a�w���K�q���?r�o ����4~��W)i��
K���8��E�21������S�9�����{o�#�Pq^975%�I�z����涄�9����}4�{&�Q��N]�v��	���1��� �Z�v�(���W���r�Om�eEÞ��
��а�Lҭ��&���J"q�P���>�m�{��шA��E'V�P�aU��Y���'Rs�Ѻ�zq�e��^ʋ�4�3Ĉ��R.'l��n��M�OЙ'.���ܼkP�1ϳ�h2��@�ڮ..�m���c�B��[{`Ɛ���?Md�:/z._zWx�~���?����%<��ti�bO��lݐw-�$��Q�L��ξ�I4�7.�K�yo닆�̶�*B7�Q�![q�����emꡯ7��+��	� �͏%H(m�5|��5 ̶���v&[�%��kƯ��MU���%v�ٯ��w�-�����9��}{�����R�����|�1V�Qz(��͗f�w�8��B5��O�&��֠iq&�jܥβs��b���mT��~�6\sp��#h�������m8Z�E�k������G���+X*��^S��4(�L*�.xjU�I�nH�C	O�7!�����.T��ݽ�����X�xL�� ���K�:�uX���⨰�-t��R�`����D�����H��ÿD�
�!q�y�|����"�����:���V��������ة�۶��7!��-w����L����aߠ�\���� �ߗ��d����|C��?~߫�I��kv �>h���P��vߋ�F��ʥ���e���3��p0=�w�~��d�e�aæ&Ub�3ܝ�����j!R�������v��;>��Y^STI�<Āhy�y\p��-懭�U/l��دٴ� ^E��ސ�zJ!�i��ʺ&�����z��<�U�cT2汨B��$Fd�{��Ƕ�|m��C�Wd�A,��r�~0[�_���K\�E�^U/�d\�9�:l�u�����e�!`��I�f�*�1袍��c���ǔiw���װ�Α:N��2|�&�l�/�EQ�>zճ|���it���͂ޅ̫�[��S=cX���!�Ŏ���޼�]�3�̬b��Ѓ��s�׾^����?�@��Ns�  Y���=�e��K��)��a��8�sE��j1���ʖƯ.R���PY�(�1ćyTc��&�n3��S���뎚�~�E?���`y����Z�'jX�t!)��
����Y��l�6����Yk�Ѣ�#�µL�p������׋���`��pl��:��Wp4w'{�2���n�^$�X&S��B�6o�5�վ;�amI���y��8�f�p�l����]Y6}|k�b
u��Y1��S��l�a��:��0wʵ�8��k�$��^�V�r�����v~wK��b	���[}]0�9T��9��.�n/��Os��Fs]�\B�ԌY��A��w恡C1g!�v	����У�S��𲫡���Y?5���fv�0ѱN��U�k=��!�!�D�Am�����L��;=_��_WT��	�`qTa⦃�y5V�����1��5��{�F�/@�i �8x���9��k�LKb�2Z�fR�޹WCk^�Z�}�Ϧ�3�S���9���+����P��vW�{� ��x9�p[����g�?�^�`l���]37�K&�w.4{�fF韠��R�ރz��KR��G��Z^�zK�h/K��k����DOm�#sW
`Я�y���&h�uK�V��!�R+y\P͐+���GU���[��ڈ�νp�IY2���9���+29��������x�����x(6��|���3�����\�LHeO�9O���ӷ,ƌXgc������"5q��5bY����B{u:轉�C��z�C�O�e�\w�Mz8�@�b�;�-�Pb��+MZ`#�6��U`��=;J��zڄs�e�^�ұ�A��C6���9!�@"A=Pճ�d�([U�sZq��+��{��G���D&ZH�->��I�w�x�sz�Zj��#��������5��W�e�ܝ$��7�C5�A}y/ʹKL�eU�斔&���s�|��c2��ԲZ(���z{��3���`[BGh>lZ}�z��C�S�{�h����7�4���,q��vɱYd��8E��ڊ􄈔�~�(2j���ڮ�`y�� ��x/kϰ�ǚ�d���U{K{CDrН����<��8dG�ss�	��(�E���+�i5�Gc�W=���I5�%�\j���F&;V��H0�f̘,�.PB�E˼s��b%9�X��Z�J�^Q��R�$��JYظrk��iT�u	�������K��oQ�������x8��q+��>��9%��Oz��p�=�i���,ZP���n�MD���
A���`��]�Ous,���GqN��歚v���2p��^t��em	Ŗ��:XQ\�ؽ��YB3�v�s_8����]�1�M�ԡ[�NEe��"�5F5F��?�ﾪ����<����<;87\�)v�癉�d*~ ��^�#ϡ� �z�M�1��}{<�^��K�9������D���[a���'�K�/��	(����Y�>zc^��vJ��щ�I92��1Vk;}KX��֫0y�Z��a�(�z>;��fiݧcY�B|�Έ��S̳<qG�Q����L�O�$Ȧ��wU�����،y4�Ъdek����Yj�o��>���C����
C�y쟋Իk��B���,8�V�9t���͢}�c=�d���E]=���Ns�Ǒ�S ��x��||Q����2{�z@��)8!tK8��]l&]�T�:����ۮ쵬��������p�E0|�`?�z�F0��f�F�{{M	���щKlS�|���UN�q�mi���w��-=sͼ*K��`�o�q���㳔�(����m�Ǔ&�B��:+y�yy[�&���d������k�����C`��y_�F�*qm��q^���z�Yj�К��e�ֱ�yt�(� ���O�PHγ׳gV@�����\<n� 4NU��C>S��]���G+�}S9��냙��J��Foݯ:��=�'��b:V��С�$�lS
�a�73���R�~#�*�O޽�"���$���Qj��t����{Z���Akeu�{�{V�W�g!��h8���q��;f싲am^A���"��8U3�(������}�~�^���X�����L*&�-�NEcW�A	��� �c�c���g�c��k^�9��'��Z��0����:ϬD�@LO;O���MQ���e�`r�N�Z�J�!Q�ѣ��
��wG7.aL��O�������x�	�
��&v��f�}	���$�,�1��N枡�(�,w�'7Q��˨Y�TS�}�a��m� o`cL:Añ�V+i��o�J9�Ԅμ�E�N�.���.Ȫ���e1W��^�&�� ͗���n8���"��on�'�D��K��a�$J��(^�[o��m�IO7�S��E�Nf�H�=5�Aߙ��K�(�v��"X-'�ms�l��:���t!�2/B^u�r�'}��
�,�熵P��%%�#�%<;�����)����� 9=��뢻<;�������Kκ��h[��Iq^��7}�V��}��fT����f&lMܒ�3�,�֧���}e-��9��LaƵ���ȴ���cҵ����cL)�̾v��{e�0XO�hM4+	w G��|H����̴G�&?
�/5�w��^�.���Q�ӧ�:�SL�zP�}�!t��{\��Q�ՠ�v�[��&{��ۯgcG#�<�}�c���֯���o#����#/(����3ڣ]��W#Zy����|U�	O�aV.;�齥�ջ��!�Un�k�v�mG�x?���<�?� ��JR���WV�{��.�ǲ��r�Է5�e���g�D��.���f>jzԕ�4��n��~�{��g�	3�3��l;e���{�Iza۱�2���lj�F3��yw�2���X�D �77��v��/�55|B��}yx�����J=0��ʺ&��m����{�_��)Մx#��X����|���騼{k͍i��C�WdΕ�C}�כ{"��MX�\�op��,��s�
���C���
���?Jxk�eC���!k�;2v���Sm|)��+ꈎ��"q��p��6�}!e���lS:���?B�X~O�\ڟ����>K��xWm��jﷂ���,U�i�+��vzs_i���[;B-���Qx�	k��������m�s�ڽ�������JdY�9�0MAIT.�d�=k�<'�@/�
뜧*���~��u{��8�eXU��L-�_&�W�oL��x��b�ϩܮ��>�_�e�'�{1�2�����.ͨD&�B\���%W���ϯ����t��noQ��9�/�.�{�i#�/+~OE<��Θxi�	|����^�]�+6"�OM�8�V!����!�Mf2T��[�o3Kq�[64jV0M�{��r�cSw[�]+o5�ˤ;�)@�z`)�t��*�z#�zQ��r���X4_;����7�~�������*�s�}�x�<#�*���|��<�LG;66�����l��ة;���YU��-E��g�
qqىݨ�\"�N��M}���x��������>OP�y}C�K�NH����^ u���,�J��v/��'�G�`���w=�9����B5�O�ty�-~�LKb`Y��WC��8�WOj��([X¼�J�)�z�"�t���;_�,������X^
�_�,q6��UL4�m,���+��=��[Ȯ3m�#�&7�u=o�1H�����	�����%줊�Ϗ{Wى��X�
��S�{��'��ق�q00࿠��}ŠvQ1^�tE�1�c䐎�
�.<���z�!�5J��>�,��6^�/x�^���mci}�H{��q)��i��s)�D�����9�������E��~(���*�^̓��S4�:�w�(�n�y�;�<ր�8W��.���m={�������|�<H���!К}Nnj}<�s^�L`co�^6,��G(֍匹wS6��J�,�nb�@���b�O���RL`B̓����ٻZ���w�L�_n7�HɋY�?*��Qݹ�];d�dw!��}��[(Yxïl��VL,�L���{ܺʃ�h:DV�=UÚ�j{@�ټ�Rt�b%2������2�y�Vn�ۙռ���KUp�P���S�;�;'����~�ע�Ҋq�8@s��������Wa����лQI� �gw߮���I�6�W���٣��ɨZSI�WN0{���
��=�@���}�7�ٟ-^����u���t�:!�(�E�$��B2�����ϙtu5t��
6���.o��T�۪}w�%D��&7�A/����N�ሔ���E1ͽ5M�z]������<T�x����j�ɸs}�\[P���jc�)��� _Iw7��NV�v�}=W��?TI�Ք���D��n�ן#ϡ�y#�C��ޖ�{<�^<ִLK�AD�@�v\�rv@�-���O�4�]qx�%�k����@�`m��m�	�%���n�X4�x�Iuf�}���v�u��4݇��b�^-o�3~J;��|Ht��:��+�t�tN�s�F�}��׍��>��;k�Bg�y�	��B;����I��4�iO�*��N��n��ؼ ���~�ɜ�^�ߠ_�/�F���.��7���@�é�kJȎ]>��U��0�V�=���K�̅z�evS���Єt1k�?62��>｝�#hgR[�(�`a6��kv��ǇU���6�K*]��j�YtE��m��Q������,ڝZ�V�z;^;�*s�\Y�iLHeZ�j�Űp�;�,U�����c+���%\�9�dC��8�WV�lZ�}�Tu��򡱪�VW�Qߙ�U�U�,�IU��}������?�"��.s�(Q��vu��5-�B��q���-�P/a�G��=�9��`PZbac����J��A�ȡ�N���ښz�����k�y}���	������@mP��?�V��73ä�'T��Rf{��]����9�-E�S���M2yڼ��JL� �� �Xo���~��RO�1:Yw�c��Gs��ts�Н�K�t&�}F�mkv�A��� ���HjH���/zu���[Bs2l�h��T��ui-�رD?�l��;�c���؜��\�'�㰂z�E1�kY�_+���̊R��zIǥ���l)�[��`��\�B9��rK��7���e�c�RuY.����(Em�o���O�=���L>�x5��,} 0�ޅEä��Y�M���Y�H���r��]���~w�}E*�U��� �v_��������xMFn�F�^i��ȷ�W��b�e�R�I�.��A�E(��+���0����|ݢ�>�}�A�޽+~��A����f-M�2�;_L��Y�09�b摵����;� ���x�-p-�y���RВ�#���-
�,��睠������2�q�	0<���4n!��1kc1���������sE?��]j�����9�P�3�F�v,�:��f�p�f��Kj;����}��[�`�J�L��t�mm;}�e]]>X�^�M|^b��(l�ݩ&8i�wMi��.�C3�f�p'�w+��풶�b¡�6��A_�˴B����.tvEcl+��n��Ί�`���|���4�IC����Z����������t���!�QN��8m�+��vH���}�u���2F�݂��b��m���]�<��F���H�ʮٛM]��*tR�,6�)�i��gu�ⱛY�P�������c�m�6�<|�ӎ�t���~���݅p3ŉ�ß{@��Sϕ:��}�^�փ���r����Jr��c����J�t(3&wH8��}�6�(�����G��NsUr�Y�{ĵ��:h�r�a��9���p��O>�7��-�.\�r��q��(�N�i��of��V�L�ì[6��X�{w��:KNR��ڗ�b�f��`Z+�gb�z1�kN�25M����z+])��]J�u�@N��@0pA|.��^+���]��7N^ul@MB{����n��ueiЀ�4��1��aX����n��¤�9��I�AO�a)b��1�'�{��(ۘ ���!�g9�>�5Q��$�j;Z�3+���[��67c�z�)>hGN��g.¶ʛ��.P�Mv^tw�ȥɳ5<b���h��P�4�v�u�3H�'v�X�;��E�}C���A�|D�N�����t�u����`�9��;���0-M�׬��a�� %����üt(����u�Kk�g���bI�{H�f.�b)bt��-Ñ��0��kD}̛̚8��l$4MP� �}�ϙok9�=�$����3�8�5|�9�\�2��F�\L��T��� ��>��Y��ͫ�Z+9��ۼG-F��]�sbV�;�h�/�(���7�<�N�Y���%�Ʈ���*3�ӑˇuZ��<\i����Υ��(�1\�@,tm>�8ie�U�����S�N��k�;�DI�_+�.sC���.[K_^lΙ�ќޚ����q��[C����&q8pm�FV}�O;|~�<n�9�k٭�3��o>W���pZ7ő>��ޭZb���8���\i�ޖGQ]d�Lh�6b�B�[������K��L�w�+
��픴�1(\LC,���(dP!�/�ܫ�wz�>rI�b��+ �ǹՔ���i��͕A�Gܸ�u�j��\V���'���2U�qm%�<a�Zn0gEk3�����yn���7 O#��L��\�0h�y)��m܁\�T-��0�<�����T�<<����!{�]�a���V+f��
�x���+e�ÌWl3)-�Gs4�2��gH��M:�Y'f�g��"��~u�b��cTTDM�QDƱW�1c��h��"
j�(����k���T��o����~���ǯ�����~�_�����횖��֢((����)�b"*����*"
���U53$P��k�3�>>��z�~?�������?{DQLU}�b*"&� ��h�h&��&���)>آ�ֈ&��cRӶ����
��
���o-UU4\6�**"�	*���b ��8�**�j����&`�͈����% ��������j**")��h��*�)��Q���H���ADT���UQ��ITI1ELM5Qz�U��UG�i�����E4ARD��TA3PD��MIRh�SC1IT1QTC�4�IAM4PE3T^�A5D�ASQQA$ATsj`�h��)��C��)���a�TĖ؈����L�D�2MR�ĴU�JQ�<�Qx��������TUPEM4S��PMC13UZ�3@�(dQ�47�t�6૷ĕ�-{��[ޚ��s�e��r�upi�!G�Z8��O��%�\�����Uo���r ���ϝ�~�s���[��Qy�:�����4(�L;�c"�ה})=J�n=�,1}$G1ٲ��z�;�)������� ��/:꺍7�2u��E�Z��2Y�����֧S7�N0��r�'�����`��� �c5�/MV�N8����S�4s`U�������<�u�P��B~a�m	��XK�0B�$Oȿ����ϗ��7�x�������^�!�I\3��+��ֽ+���]5�|��r��R��@���+����>a?��:��;��m�Ϗb���6�������v����,+�\�;��_����W1eyMQ/A��SD!�^�&ȍ-b���9�P�_XP��dlfӳy��,ߢ��c���28"�Dc�;"N)��=�r�xlB��k|�d��r��c5闏��c���d��o����jo3N,;���`��t=C��x�X`d�d]�%r�������;�vs��l�P�.��;�Zr�q2u���^�aC*.s�=�D&��Z�8�yc%�K�,��P\M�˼K|��O:���YK���&���z�'W���1N����=���p�^O{[�ws �6G���ڠbO*�c\(�����$ַ�ҬM升��X�ѝ���x#�x@�E垅z��R��I;_k����W���w�~�z���<;�^�J!��8E3��VJ��5�&�t���Q½\۞JAe_n~y�W�5������
P�.������a�o���f�ؼ�E�9]�BB�{CM�nr!2���%B`�G��e�:6��C�ɬ��`�S����~b����p·2�� �S�y�@"�ϰoL��x�E�s�Ɗ4�S�W8�5D~�k[�������������2X�r�p�*��N�/����t�<S��wk݊�v&�����P��/��:���̜+���F>=��Q�)�Ozʮ��Pf<��4;�Nr�Ι���)��cK���A8�x`>ϘG��!�Bnn�IZ�byј,u��-ϼުo�6�W>�I���V���إC�P��?xH'������AֿUtSwL,xL۶��TV������
��d�Sjz������%�^S�j��������8���;Y)u*¬��Z�IО�C��i��`<������*Ll2�O��}8��c�AۖcF,3��3wX�V��l�X�2*ǅ�%��"'�ߥ�>��l��_�01�/\Za/?~s;��d��!��\�n�\�)�{t��x�B�: p>��M�Fh���p��|jM��q��q���:���w`�0B���y�37�K�ӽB>��;�g�u�4�V	�vwm!jk
{4cN7H��_j�����:aNj��hjA
��@Ie� S�~N:oz��̫Vn��52��B,[�v��p>"���B9��&k�p�L����x.[wz�C>��g����ۧ��wu3 ��k�[����~0���r�l��M����kX���p��I���׈���+˧XqW!�%�<��m={�mᵡ����˙���N�ojG�ױg�mI�{���u�O���3�~l-�`Z�Kh=����z��]"���c�(��dq;ԼN^�x���D;��){�������z������(2j��I�l*�|~���5�;W�a�.��F�Lv�5�H0.F���5��d)��t��Q,��0$��FMJ,.�^K�1�8���Yol����F���2�)0X7��'ד���9w�䗘�f&��}D�}!��P-�gu|l�ۜic���9�Ly���B}!;Q�e"�Y�����kN�m��`��k��vq��]z|fc���<�4���5�/O����ǐB<�:`:����'���3b���N�T�]e�Ӧ�}���'�K���:�^5lp�|�l��}��}��l����7��R�	��#�W!��yG��dd�4>?<��D���-�˓ߦK[&��*^<8��+ Ƙ1�%n�S�~�����Ǡj���q�8jG"�\ �ˡ+�It�^){���h�*hV(R=Wq]�����eAL�3�w:�u!��[q���}�S��|�������{�����'s5@�����n��[�|��U�Z��a�}�-n�y�G�xQ����t���4�k���?�9ݘ��dN��="����V׽	g�X��}tk���ʢ��J�ΊU;E�sv7}&|>��z!�yG_���������i��+u˧���{͔��[��1�+}Gpl˭�>�K�/�(4Xe��� ��g���F����g@�3h��f��v�seZ���8����W5�-��؇�ϼ"��0(,���2]�7k��ݜ�����N�]8i5\)��C���q�wtE��|C�S��J�2�[㨟vN�0k�ۭK��w�^>O���V�cv}JF׷�s�%8�7#�lӟ�S�e{dS�����;�����m汤D���Oqm��j��6-��A���A���,��Fu��gj�������L��
�n]?�EyC�h�2`{�f*!;z~�V��E�/��a�@�9U�}A���/2�S��;���{`��P�3�����'^"K����i]:ɨFB箈A�=iT�o4n�i��%��!PAj렁������G-ڒ�sm�7b���
���Lʹ��1�IS{F��ܙI�F�Ьh�Ml����?<���%W�����;{�2K�����T&h;��7���[��AښN�Oo\�*��}^����� ?��=�<=Wsv�;�<t���.�F�QaM^[s�]Qpꀸ�x ��z��L%c�gK1�'̕3�B����[�[y�DJp��ZS%8��l;��oD���t����x�!��m8�*Uf��|e�F�L��`&(t	.Wt�0f��w�xa#r�h|٫0�V;����C�O�08�_@�U|i��`��QL��`sM�.j@����H.���kU=�u���u�Z=��O"�w=K�~��B�L'��.xlU	��)G7Q7ɘRr�-6]ݨx�8��daI��b��X}?��C��Y�<�F��s'\]�����9_P�֥;�Yc��n������"�Z�c� ��8A���[��bA��kl
�]O�QRF��;~��Tu��t�#N<}=��A/mr��J��C�ÿO@`��fr69�@|NwE!&kJ͗�=�Y��/��kW��@��k�C��5-�^=�׌�}�H�]^Tyd��y��k}j�p��Z�O���a���l�l�;�XP�\
a��׸̻O���4:��0t7LM]������f�os�������J������;�W��n���D�*��W��n!{G�Șy��b�\e�ɣ;�ڞ(lit�םk��:�Kh>:��]pn][�����eJ��lL��X�N�W3Q�paitY�>|9�~z��ʇ��9P�p�'{��ߝ�~ȕ�]�="�L�Sȇ�|aB*-���zq7���B�A!�%G�,]a�1�:��n�XF���l�țxl��|И�x<�%L��咝�c9�ڥ������&���7Æo��\��	��9N�[�:n��P�1l�0�a�8�R[��U����?l����|������]���%�7%�B�Ru��ޛa.:k�5�_����4.���}�KʇN��e�=���d�s%Jl�r��PX�R{
�h]��ס�V������m,T�O�JQ\#�P||WR	��pi�y�Єȳ�~@�LR��]�FM���o���[~c����3�)��j�Yk���By�|k��锝ax�E�s�1��&�n��yj��{-\C�7����['#~#�U��| �U� ]��(�a~�R��T�2��׵w�n�\�QnC	�nO���6�yޚ AC64�M�&n�2$�N�XG�L-�O;�{���=k� 
�Ƃ�0���I�����s�B��\����/�����w�s�7h�k�?y�9z�3��B�?i��U9|r;�_+]` �ysuFӛ[rwE������\����bj��z;�v���.��q���54���6�2�Ė=�+�̹��+5��o��p��2Z��{X�Ulmf�����栫H?ӔL�(�z�z����\��Y�OδM��A4ܺҡ��C�3Nл�F�=��s$R�X�zY�Azp���>h�t������5�����B�ڥ{��ϵ����hI���ɛa��ҵ��A/r�)G4��f��������ΈV��F�X�	��C�~gfm���O�Sr�����}8�Lsp��ly�H鞜��8q�T��:�J���$z>�$_,Ղ#��y9/b/�Ǥ�qh���������mۯ�3���Yô>�yğ�@�CB~��>��kA��4$�����m\��b�_�V��ד[ڪ��o4�
�S0yh��n��p��~0�>�c@[$��z������3�*���r�of�4�9%�RYAP_ E��'Ƌxj��a���y
��-�/�^��{݉��ｘ��К�N=^�4�	��m�vPcAd�ԑ�C6q=cռ*�H�z�\����Y5���f;�\0\�����2=&�V0�bv+ӼD��Q� ɏ�)���]9�q`���EU�I�,��6�#�ZŽ��{Uܲ^�s� ����ߔ�rB�Ed���'9D�/a% S(&��}��G��\�/=Su�	�ok�k��X�CR�f�[ϯ�9�ۣ�ɉ�������ѝۮ#j�.N��g����c2Q���=�����B�1*��>���0P���ox:��J}r�֜A����xAY;��с��<ú�|�ߛ������	�s��(H��� �#wJ��;����3��)��=!@�D�fʘL�_	O����'I�t�k�1&����ySٺ�?.R)�y#H�[O��v��������a�p��p?h��`L��'`0J�aF�qm���#*����w�r��F����5�e�>G�e��BFy���,�Ŋ��ֻ�!'O*W�G�e��J]�0���='�r)�Qz�����M0������>NF��l���6��l�he���'!���^��*q��)EⅩ����'ćO8��*v}���d�����g̢>���2/b��:�="��Gu\����'-c�o2��0��%M�p�J}�̃��}�'���~�.!�yF��/R�zhZ�9��z��2�����v-������/���׈���6��:�G��d�q|���ZsʄG�ɽ4#u���<�ZVž��g<���F\�]4��)��r+���-E�;��x�y��hPZbac���uUE�LVʱQ�)m���Aۭ��5���M3Eی#㿻ϒ��P�-?k?�J���0'ꞟ��*]F��b�'x����ȑ/��{}Z��Y����wYM�K���s�{Χ�k�4fkȀ��{W!#EA[MI�*ޗ�eG����bcӚ1鼎5��2����&�%v]JEҳ"�+����5m�͵�ҡ,�7/l-i^]]8�����]}��}_��{���(��K9�Q��7�cS���l�W�>���Aq�]�E�ˡۭ��Zt^q�2\a�P]����y�#פl	��S�i}��殱�Z�J�H8�rnjK$��Fu�WU����n]���8ϊە��r�^��
H�)�1����K=[���'�8���;�'����ٴ��P��/v���:������̂qt,D�Bby�|�z���2>�ͼb���2##�-��l��D6C�\�R%TXSW���PꋇUq��"z��b���h�niK[6�wrf����MAFzK$�*"S��J#���f�IȺ��X��	1�Un�����0:���(t'ղ͡�צ]��ԩ2��b��E�W�����w|2�F,1jM�+��H~�J�W��(�9v�ǆ�/����}�F�?|���Y����1�~�Ʒ�k�T��>8|V��Vي�ם�?<�{h^}Cw=K�~�<hQ�4�U��W<��W(��n�=��C^�G9SZ�5�Y��{rC���2nw	��	y�T:�G�͇2m�͟�������L��.���p?�q��+;���;��x�󉜢��4g�#+��^�c�>���Q��ķ�F��f����x��n��
D�Xy�֕Vs����5��M �fL����b�:��E"i���݊���ߝ�ޞ�ӛ�	����"Ҕ*}8W%&-Vv��jRX�ҭa)�Z���z�~�U�WW��01�����R4�%Bԣ�lM�t4��w+�.��S�ʏ�����Bi�A.�`��>����T�:�U)�Mov�vY�C30V���0̌�j���Z]X�U��~N��j[���^��g2�w�ƻ������1mn�w��:�� naيuٲ��%���I~.����;v��o��ѫ���a���C=>�˺	A�>C��C����&�6݄���y���C�US�f�30zJ.磵�D�����������C���	Z5�?|��'�+�%;��Z.�/z�����<E�\��`�=�e3}���ȷC�$h�g;��t��Ћ�>�E���D�eY|Q��_f�3��MՅ��+���@�#��l ʼ�(QJN�~ӌ&�*׶)���f�������dw�y�}oS�ծ��9�[N�75{��M�˽A2�R�A������y���ö]C��Y�����9���y;e��R��q%�f��y��<�Є�V^%9�T�	��J�v#&��}B��BR�aw���d�����sr��ݾ�N×]U�v�ț3�[.�u�����f���f�us-ve��p�ۼ�a�E�f	���e�fw$cެ��J���+s�\%)xF�� ��#{��./]Eڨ�-'N�m�������y�9@�؈���	�#�N2�]}�s���Ob�ՙ��
��&\2�ãn�8�J�
�9��V!w�]�Y�~[��C��X*�Q�CH��b����$����DwC??e�d�g7)��E�=z�N�ӧC�#�/471V3�r��j!nZ��,c���ű>��ڿ��-�P��a�f��3�M~��lyVj�A_���lK�g��ODl"�*�x�\�d�Ŭ�!�c�360c�`�Fi'I7Zr��0�c; ���Y�w>�=z
�fR��m�_m�}v�j]��ȩ�7���[*Z�$���Uk͎V5Wӛ7U�X��J���X��ٜZ�Ǵ��Wr���v��f-f˲��u4�]=u��vzr��X���0�"m�l��\F�ɛ&�0o0ѱ��U|�]�p9�X�����\�-@C�p�{���2z��͹���@Y�]o�F�U�6��m�#O�_}�MSi�f�d�aM*oD�w u��F�NK0���P6	�/��qA-������4�$��%��f%�6���XmS{׶/5�^#�:TF^F{�V�7���XhSb$��\�������ǭ^ù�@����1<b�z�GS^�(|�F��$Ƒ�pS�OeA�|뷶�]gz$��:9�b=���.�&�_w.�B�D,�੾Dw[�+�]��w��(��'�n�Z"�����Uؼ�k�Ln�#��J^HH \U��C狺X�mf��v�G�Mv�]�"�5�4a�rl�}Ϻ��mn��s�i�?^�DDm����3��U���jS(<�U��jP�#+�է;m`9��޾�5�V�6*�t�d����9Ӵ�uݼ�WV�W5�#Z�+d�2�����Qs]���/#���B���ǆ	�r�u�����q����N��x[Mo`k�eU�*5;ר$d��wlY���ŝy�(������b��3:�r,��,S�[�Ԥm�V��2�z%[�@�H�i3#�&�ו�C1ҧ�p�Jht9\�|��՚�k�;�kOAg�l2���t����)�*���AQ�Q���۰���P�{��]�C��k����dW��Y���;g���@��Q\f�[ ����qԭ��⩕�Y�E������5�ʗ�"�]�#�RS$� �ݵN�vV���m'��&�h vR�d���؜YցsM���|\1 mo;�&)�>٪���.��+㫜v;��e����k@N�@V���1����J(`͎�Cz�
A5�o/R�s��h����A�$i�(�bmA,��o{QCM%35TTD�4�$�U5W�3�o������������~�_�^�5EQUEMUPM5LIQ��5U_6X�j&
����+���篧�ׯ_������~�_��؈J���c�h����d���������sfd���Ա1\ڼé��츪"J��&b*j(��1����(*� �����QIMP�UP�^N�	��5KSU <��DܱSP�m�j��J*��i�]i���(���&�h"�*�"�*"bh����͚(b�|�D�i�Ĕ�PQ�4�4�T�DRU!EECo\�4�MQCD��KT�TLyh

����
h�� ��*Z���*	�yb��N�i?X�h��g�5UDTAEr�PE壖�������j"a"ith�͡��/�{��v޹��=z�SA�.D�d/�Vj=7���[�w�Z��t�e��0�㹐�������4�&̶r�WPt9� ������j��8��5n鴎�ِJȉ*�I�m#DIJ����%�."e��x/8����� x���9���_|k���A$Q�#�j�����p!m��|�0O7�'�E�^�锝ax�E�s�0�no!ϲv�ʧ�ub�/:�(+������=	Ծ"�g�K�"U��}��.�5fou���Q���<�i�����^)�z���%���h����ѻ3�I���|Ǩ�ǥ��W�l��1�8�N�l��E�j�IWCը���9bB�0���w�Gd>�a�2ng!����?T
h=B6���o����(
�L9�ږP�JL='�~�27],��#ʐO����ZG`����\3�W׹�>�����>'T&%���je�Mc=�T�/t��\�6����e�14����S��~c����"}��-JΖ���1�2����U�׻1̔�eK��.��.�Ȭ,ڶ�<2�g���=�y�<��{�o ;f�E��Ǥ��K;3����*��iPo�>�Op�d+�QB ?hL��	w �O�Cy��K/r��W�A��{#���3�%���j5���d�3C�I�$�CI}��y���-����ƴ��$�'mՆ�[-YnΗ��]�T>�7�͖BYRi=ؖ�v�u�'�կ��t��W��gm�>}@ɕ��pxj���k���.�I�;���4�b��-��ht��-�jf;�ef���)Ze��X	��%&��%a�ziH��}���
���� �0 ]j}4��R�F�w�i��#7:���e�����rK�y��O\�o:��a�������x'��Ȳq����{�;��m�������#�6->�z������ ��n���3��u�1�hs��^5X�+v+�7���~�3�5��H��t�v��#��s8ӉȬU����9��<�#K�DW�����C%Qj���z�ˡ�0���t��������{:=_Qτ��7`7ذ��g�?;8�Ald��vl�&>���<��XTh���&�e6ѻ�V_9׌D�T����Q���rZ�"��?���JY��%�Zݝc�;��Fk�:P
�.��i`		Q��<b)9\�$��\Ø��}���h� �s�n9�])ܦ�}��L��}!cr7Hd���K���&�w��)?#�P���*A��4�A��6T�^#J��+5�fM�[��\�t9�z�%�=N��vr��=vE�H�P�Tw='�q�C`˪�������w�ةݾ����#����U��ϡ�9U3�j�����M]��I��b2m�[��UƾS�UԲz3�����0b�9�K��v���dK 6��&�Rv�ǵ�ҝB�7��a�;�Έx���7׭��[��Ay������}#t������Ft�v���|��rED�����C�WJ�rS(���;s+�}U�>�������H�ORT_l@e�x�~�ٽ� P<G���4u}�B#�%�Z��K����w}l��ܭuu���S�J}[j��A}���uv���}���ŤC�az��'��d�<�Kf��o3v�dΆ� �j��+df�W�����^/�ܵx��q�H�����6��ƃ:��������M���[Uxf�>��;s�;��h�q�b��pt=�sͼٿ5C�uV#ae��	�*��F�Fc8gU�qO��L��1m��6=����47����F]���>�	l^q�j��^�S�}�<�ञ�b@>~y0��&�}F�Z{a ��A��,�BX)��~�":O#�.sp��t4�7V@�^P=�iVi#�mpyF��\�'�dT{��!?7=5�$sS<�e�b���U�r���?<�yt85�5H("�Iq��;X]:ɫ��t̑�9ӛo�9=�����{	E'V�P�~UE�5�9/B��h�uB��9oP�"���w��O'��;h���6��-ͣ�$�b%9IH�UQN.��H�v_���X�[��-��8�9��H�����H�i��nm�Ѡ��b}<��t9b������u0LD/��ڼ0j
`��\�Uدr���f�'u�[*¸���]F�$i�*��޷�v�u�P��+��y����+�z�D�f��WU�t�K|{�?���fQ���:��3���}dV�S��z8˴��m&@�LRn�E�Mb�{O����YZn�vT�Wa�x`���B1����pG>,.$S=_v�꒞o���u��5ַJ�h�m����AX��ם�?<�{h���r��K�~��B�L'�fW<3akv릜�E����e���L�R;P�Bxw��|yp���M�"n/B^u�uW�ʹ�Ӂ���cF�s�N-$h����dҭa)�[��+�(x-=Zx�<�>��Ջ~���U�я'��v*��^ۙ8��X�T�_ˈ߶��C��a����8��ϭ<jd����:[/@}Naٷ0^�oj�J��Ț�|�P�;\U���t�/~/��%�K���}�cy�}�g���AP\Gɽ�����͈�����sʻ��@��h�I�1�,����3uocX8؆1eb��D����hy�?5'�n��y��w��Jރ������?���g�[�߄s[?`v}C��ϵo��|��'�+��
͊�M���E26�X��g���#^�%z��XZ�A��LMÎ����ޙl��s�n�@�A��V���Q�Vf�/kUM�uʤ�h�wpr�{*Fi��9"����؊w�C%�o�4S����:c��/s�	Go:�	�]L�w":�z#0e�D4��y��3y��'���eL�u�D\�3�ULgc�Z���_�r�P�k�7n��b��<��, ���]�ކX��U.������j���G�e�L5�\�Ȭ�l�󇡽0�.�>�p����:y^�~�ۆ�At��k��j�Ȳ�)�vF6���nj��!I��L��kZ|��.���{��z��ˡ�Bm�N�1�2��5���	��M�x��|����BS+/��	��2%P�<�;7�r�*�>Sv�ce�Z���bfJ�dQ_�w���*#��[���q2[ŉ�-�n�=�b���h]ڋr��L^y� �s	�k�<���1	��!�/��W�]�wAS4<��I�`����i��65�[��Ӳ�NZ��k�SO�P͍>���`&�Oy�<�[����wUa��C�q4L�:���ʂƼI��L!���}��=�d��<�J�<���Y��K����������rE�R��Z��3b�8����	�b���(o{��u��� �����:�B��G�9��تv�[+ ��z>�_=���WR���&�p��׭�� ����mӯӵ9��z���������=v��#��� �j]!�S���@ˬ�Վ��iԛ�Լ^��"θ*���0�
�m��v�����slc��q��*,3%%g�]tm�M�����Gn+�]���J���K6��S�3�>���y�>�����0w�B��� �a1�~�@���D��b���\r���GS��N9�1ݍH�����
v��c+7,�9��O,K�n!@x��~�������hZ<����JGz��L�z�wp(��>�uŠnW��z|tE�J����g�9ľ�Pг�'�,^$��%����zək�ј�*{x� !Ʊ�4�D=qhI=P���^��s���ZZB������O]�u����bv�xi/:�ui���j;)0��YA����y6���.�9靼��wY��N�l}Ř-a]�R��T� �B���S6��A�,�`Z�Gh=������gؽsYT,�>���-w��H�x�-����\zz���	\�W��%6r�1����X��H�S ����;Wۘ���{Lf�4��=5��!@����	~]���\��'�ӭ�18��4Ƭ�%��ywM1�J4�k����9�<�������]�(	��p��6����T6oJ��c�ד��u�%��D�7�E1�i5����S�[zP���0,���OQ��\0�WC��'�u�a�]z��ژ�� �|,b��Z����Y���]Jh�lg8�U�b7C݀@^�o���VzZ�ySj>˜�4M�Nm�r�:�]]���Yz@��(��{N����vvd|��	���l��W���k���i:[�k��b���q"4���E'+<�5���5x�Yz|�>Ϛ-�@/��z�;��+U��://>M�&47^�4׌9P�l�n��Qi�&�K��#�D�i[m3�H������o�w��>#a?ׇ!L��S�4�~�U�w�Qx�jF������:���h�Q�/ݎ��B��21��xk��ܑ?.�~�M_T�(�>�w�~k���Hy�a=8q3r��'�ds�s��'>�W�}?0:�\�"vk �0�C�vnt�D�s���P�Q��Ґ���rWv7I���X�n=���Vǉ�w�l/Ө4zd��x/����<���\DsVL���;n�0��;����JpK#4����K�\��HqEA��G�0U|{�}��٭�u�5GOhe,�cS���P͠��ؤN�3Eڇv-<c�ĝe뗢��Rv�g�b�y��׆�Ώ
���b���s����sc6}���4��v��� ��˳kpʉX*"n�[��_:�oCdS��@��a�����*�}F�kZ@[�5��soC�
5Ҝ�sd[]�]�ĭĭǇ�d�Вu�c�C�6�����;�4~ù�>�Eߒc}P9xPV̺4�=n���Z���DP�Q���6wS�Xz��H��nW:��q�>��^�uӬYw��zTs��њ��]����;�sa�,
d��[Q~��?_��'����ߕ_�cj�*��+�|��Q�B�`|�Y������l�Xw0��� ��붻Q�J8�@@�4
��z:�/�yq��@ft�X��1����t>(��'>����۞ӹ]��E��^˗~m��	��"W*�a@5{na詫�e?������NԎ��/�;�DwkZ�0��odp�})����	�{"S�H�O�	����[Bl�޹��*�69�:�����C�!�e[���f�y������hOv �J�MY�/2un#�-\�w�xa#��gb�����}YP�4�}0S�(�E�H����g��n��.ѭ���n�G����;�׏8��|C��>��]'�OM��D��I�<�����d�,]�1�j��׆Z�{���Ɨ�	��n;��6Ȉ
���~����+�U�Q�ݻ���v�:�(��qv�����f�V���Vt�T�z�����B�6���0��+��>������M�eP�~s'PzV��������d���p{w�p��e��Tj����x^���0�b��<%�7�=�:@�u(��>W���&�[ó�pp��n���&!�M��Ŵ��a��K{�m,b���R�xպp	F�i/kbޮKHޠ���:�9�=��:ۓ��K`�L�L��������1�� G��>
���~���p^9�s<+C]��.���%X�U3�3X�,�z�\�����=��m�B~��ܽ���-�(&"�Ū�Uxo�#�0y�����M宱2O>��l��E�����.�O�������xا:�@Ym�^xw��.�0 h| ;�'���[#`f�\0�5�}C��`��^��3�هc���	A��CO��:�9����'?x;�
��+����3�+W��c��w�!�
��,q�?%��g͢�-�P鋇��,�� �89�v7�EGJ:;���1��M@�ܘkl(��u�d|�(�Ru��͜a71P�)�6��=���.���\�ڷg�-1���`�֘q�1���T��7���`��,��
OaQ��'���{��V�R�&v_sm����
~gh:-�8�������7�y��҅&��%9��0Mf�tt,�e!;am�.p��o��5��88��|�>__�{ze'Jt���"�vnq'~�9��W:E1��Ɠ}��t|Ʉ�\<�k�D_��B����H�����bv7�5`�vW�f?�=ⴶn�}�~Â�����2�9X*C}��L�%�m.���B�3��y��ɴ�4
�>B��#�=�H���:�Gs�����cu%9�73v�E+z�rW��9D��;x�k۸�P�Y�:�=T��ۑr���}]x�,��b��q.�����3��ynX��Q��,�^��L�vf�S��ڏB�4D5�󳪛�܅1�2'W��w�eOC�����PX��0���h:}";�ㇶ["b�~�]��;l��������<s�������(]�Ta�֣X��jA?��ڗ�x!@DE?s�V�}W�ݹ�]��u�Xw���?k�<6,�)��a[�V�����yN�]���/t���do2+4��`�v[����īf����.�ٛ-�՝6��r���5>V5V�-Ǭ��xl]�f4x_L�v��֯�����7ʁG�k��a?��A�y_��*�A}8�q�)>��_""]�=��=����(Q�i)�u���N���Ǩ$lji|X�B ����e�ڗ�Fh|�Qq՘-�rŻ/d>�����z^�����OL6�-�;vD}q����]P_L�闟t���]�N�P�Ys�M��ͯE��O��zW��-��P��[�x�s�<7UV�������T݄a���u�"5���1��>Fs��O���c;Ί�f�B�E�=��]A/�i�/��K�^{�O���x�4�W`0�[t��Ɇfܙ[�`�
�
�%�Y/t��\��Y�r f���e�����Ӭwk�7J3b���ER�q��,:�ۋz
h4E̾ݎ�qF�h.:sً��,��V��eXn���#݃��[Ūc��^vsu/�:Cfo;+���7�
X���_��Rw�U�b���;t5�_fX�"vf촜������sKf��9�(�M�w� �	@�[���x�F��|��xN���KLPܨ���r7��[�q�h�sK�
]���\ȫ5�'�AK��S#���rVY��&��ٱLgD��˫1��P��C���&j	6��Fy�$�u�)ND�X�ΘkjJ=J�r��T5�|1@L�,2N���X���Y(��"/t6���
��7�Z��>۽|�=l��C�<W�(�3(�]�|��� �x�����a8j�Ȯ��Z��(b��ef�"��5�b�� �u��}:eL����8=�y![�yH�镘���zh$k��Hػ��ղU��.J�^W|��k*Ld����"��+uȴ���/��.N�C�a���A�(W��V�R�FyAkM�dP�i�sN5]|��grN�J`b�K����t���u7�X�MةO�I���q��t¹`8�R\p�n���̲Edń�5�r���yj1���,������+�E4E�u�,.lh6;�:U��~����X��1�gAw���cn�4e����w�)�f��6I�Phkx��)*�� {qgtb"g�+�T�v>�����V���M�(X�I_P�1S�:R���Ʌ���F���_K0��Z<�lL�\���P��O��s��K�
7��+���	I�0�Ƭa$>���Q��(�1������ۅK��oB����7/���F���+����%����H�Z�̹��t�L�b�T�7�w2��� 8�
=�m��vgQ���вޣ��]��Q�x����� i3����y���aGl����m��09}W�Uq�Ѹ�}�������a�K����Mw�9��Q<�����]Q�
��˭�����_Yϊ��y�c�e������sf��ے�Zn�Tj�ُ�N�n��n���ѬԹ7!V�P5x�'��nۭ�N:}���i0fIN���R3��텂���xTUٷ��\����4o��3�����7C>�)�8=[}���W{���k��~u)��!���\��r��hku�y�!M�Gl���%s�����'f�cgy���ʐa�ZUj�.l\�n����:wZ��s�)�)���m�#u���U�7q��":&k��ʷX(�=H��V�ۭ�ۘ�jdΏ�EKُp,�%4iJ�y��B&�w�)t�g{-�N�ml ��ܔ�-rn�u���?��B؛.�m :�,�kI�rwn����ﾠ�4�MUUEQ�l��;?9�hH�b��⠋�j�9Ϸ����?_�ǯ�����=OS�J����%"��4��15TD@�S������ׯ_������~�_�罊���*(�"���)����"f/x�G?cG->[�qG�AET_��BQIͨ��%���.���if"���� �����j�
"��Z(�O'D�IP�޸�<%����*�+�EP�KQ-4�,TRD4�	14�U5{�D�L\Ʀ���"�����'�|�^F )����Q#K���:�hibZJ&���� �娓��ʩ�������J�}Ά�jZj�"	�J"���B�4M1Q\��	0�:tQ�D�,T4D�PRRU$( *��P���ť�Z��}�&eu��M(M� �7}����o3�n!C��E��M1���N��-,ڼ�������ɡv�;��y���f1�$�E���[�����5������\zg�L�lNEz|�|E&��M�7c9���,VIx~9�1�;�XX&/����d��|���d�D(c���lVE\�t���I�1�Y�cf�n��{�Ji��4*�v>5{gO4��A�<f��L)ى4���Ó9�O=�����҈,��1�ߊ�Lh�[���#�D�E�?����YNʚd�roq��0{L�C��"�Y�M�q>�>�p�<b|�(�U�9��Yz|�:R���I���ѱ]d��!���F���ٽ�)�;SK�=Q/�4e��1���y�6�V�������L5��q"kН���r�Vas�(	�ݚ�H��ؙ�Up�I�Un�9˸%$f;(�<1��/�#��d�j��N��W����ۙR�:�!c3�Ó�f�;\#�%)<خ�W�]H��͌����Zq�����E�6GV���U��o�}��$���S��
�F�Ǿ]>����,?�A��d��x?5��x��N��O�����������5�`F�dY�!��tW�|�ig Z��*k�Sr�t�s[�o�,l�Bc���C�5���4^v�Sq�n��x���ܧ� ��;��.+��oI��;Ĩi����-��e�B�N4ya����yy����z�:Y�R�t�	vO�_�	8$2���_�b��j/a�G<3��_!̮�j�3���6��#�!�͹ɀY*�_;����C��sI1��N����l�4
ѳ9�nm?	0�YS�D��~)�y_��9�P���^��f��ޕ��@A��պ��j�(�Ɖ�ӻ��ۚ���x>]!�4&$��j��N/�L��~����:3LWe�2��ڠ52rt7��m�8��X9RV<��7jn\�)w�C�>�D�W��+��2A�ְ�OC֢X�ӌ�c���ʘY��

�x.�pՖ3���kѵ�`�/WN�j���@tA���9BeK
V���1ڋ�DW�M@q~���z�'緓��{�J����
R���j��&�S��	�r�	�x$�%S�|�a6k2���U�޽n���Qy��?�6h|���`��~���^�ҩ2�-��LP0&�'	�*�5ܛȽ�d7*�7VB9����O� @ �Ƙt��`�|�`�4�!�U�~��e���ހ� E<��E/���,��ө�.^��ooV�_%ԡ|%D�8��c�7m�U�g�I����٪��Q&����ާ�ֳ׶�N��n5R��G��Bm���2�qr���6�wg[�ċV��m(�h�vӬ�pk=|�l���A��?�� Y۽�v{�[zxr�n�'xK�/�ᔢ�B����ʒS������@��*�o�
%��N�M��Y��Ы'�Lxej�I���4y��xw�o!Í�&�p�y�q��r�*�Dݡo�{�˕��mb��/������3~�Z�|��Z@�����vt��v����0�{Bv8�d��\�H,��̜qǡc�PK�?�T�	k`V��{w�����x3�����nΘ��8� �=�w�nZ��D;2���g% �t�幧{�ƥ���T�`���v;X�̊Cq�3����A@x��L#���*�<���x��9�I��;�NB��f?D���8�fD�l�tg/<�ꈟ�1?hY��Y���ٱ�(��&�V���Z��o�r�t�C�l=6�^)�37�"e��}��%'�-��F��V��k�~e�Q�>��A������G���-�W�b���~�h�"9�]�i"7uN���1��
+���M@�Cr����HZ��J��(	I�^͘D��/��Z��7���\��Cw�/o7ғ�7[��e�j���yk����4V7���#�W,%$���=~�Ԟ5VX��������/y�C��9���ȉEd�=s�s&mf܍��ᔺ�mXRN}>wժ����1|�L��=s4�ȶ&6������������֎�,b�i��@��5�C�O �c%~�,��Ȥ��H�[��Ĭw���Z��D~���x�����w����o>��v�6-�kw������Ij���(��1��D�[�Wot7v�!�#N=�+��P�e|��i1_��B`$�| |g���3ї3��,�=u}�N9@�Kq{������+Ѯ�
._���3�d����U���k���f��ѝ}���u�R�.�X�R���c^��8�S��p���N�i�X��y�+���^3�����^�Y6,��I�H����='�⠱��a���B��-�T9�����}g�����:� ���Dc;?:����ᜲ��F�F��P�z sm[_[<w+�؝]���u�*p�L�����8s��1-��u���㺱�ڥk�*�ŷ���By��n����x��ݨ+3,ȹ�s����{���`0~IZ�/���`�T8�E����7���n�su�����>�z��KP�Y���x��02"D�)=Ez�=z]��{6�Jԣ��uͤ���r���A�`2f~=g����8�ٝ�M����N�܈RB�m����x����9"�狺oɏ5wK46���Z
*�]�����VA㑓����/%��qT��C]6�Ԛ��U��몿����.��+�>����)�ua�zZ@�ht;������;�3���ý��pi6)/��n�hz=s
�З-�6C��V0��������떠_�?�tEC��L�&F���U.�`ݮ"��p��2���0�D�c�`ͯE��3N��J��2a��E��D[5��2��[/^�w�&~�)�xa�a�V�����?^�i��j!��ںq���DC�U�e��-���Iӳೝ��c��@t�-�â�"��*f�#`NEzB�%6or|p�=��ʝ1v^�t]����=�@ӌ=[�M<�^z� �fz��" B�S-Z},EmTv�]�;�y��A�'�E�%4�ģB�(�|j�e|��W�'�M�7^6���}��7uv`P�$`�_I��ĲN]�9�S(�kgځ����}�e4Ꙩ���۵�W˞WÏ�~�ƀ���
�H�z�y�oI���1	����(�*��5�9�i���	:���¬�N���B`��B�r#�j`����%=��mܲO^����|��f�3����5�ƝkB�gcݔz�jo
q��`���w�l���U�m���1���0�A��,;�/iB� 7`DV�.��XD���Uim��p*��N�<V�t�<��FtiǏ;�c�3��������M3u"��F�v�ݶ6x7��ߚ����T�d��tܦ���4�~�LO�p�0f�Z��ޚn�g �U2��.�e�:fz��h���I��h�ig�@�"�㸏�vǶvc������צD���n�s8�-h�g4�W<�l^Jx��]<^e@�-����vk�`�� ��"���]%L�x告]ngd�����W��P���a��X��=<δ�`�=��~8!����8p�%��59���
o�ae�mx���?��R:U�46�Δ��.�aC�@�q��_��P/a��I�v��Hn��(���!��D(��M學Ǐ���b���+�[��m�v֯o�5�u��D��͓l�ѝUׁmo�",}�Y������g�5��J�'�M���Ϣ��	�� �&�u��v�1=nD�Q�ְ_�}��f��."P�`��Θ�T���^N3�%�::*v�>,�ճ=�����Ed�ԑ��ג��9�+�9RNǟ�~���5v���Ŕ�[�ޫ^�?����]���q�
���G��8ދ�&7����q.:kլ��|�왲/
惡k��j�b�X.K�6��dq%8/�>q���@��R�{���Y��9 ����g��>*�`ͩZWb"��V�Ҧ۾�I�P`�Y�{�n��)��8qJ��a�3WA!=H�qԷ�Ea�1_'}qIx��`3��	j����#��K�=���J�'?����~?�	��8�һ���-�û,�)9YfA8��[��0�7'�� ��D ���*X�W�I�C�gb��l	����/�7�Bլ�� ��#�Y��N�3�ޑf9�<��'.�I2

d�p��ޙ=b��B�{�l(��@�7�5[�r���2�],�4���HޓI�0!.��١
���4�f�y�r�jo5�zw�xa����DcL:O�0�_@�T/�;*��ꐟen��=;�bv\��F�QLK��ZqsHӱ<��^<���8Xٟd��Q�S�M`W�����Γ��]�F3�&�xej�t�AbW� �4��k��w����C�l��þ��gQ}h;_:�����Xd닰8�,/�|}<+��'�Ιʕ�,	�^_i8S�>{̭�6�P`�������R�jÙ8���r���"Ts	[Bu�e�yZ�s5�v�g=p�����469��y�;2���`�9)��{�s���q���h�ɻf�݋[Yab�P����0M�a=�U�)�u�0̓��;d��E��&.o�=oZ�+��ǘ�s78Eu�L[��wT=6��k!�3�h�e�_dR�@c���l^A�@+{��隻�Dd�Ɣ�P2Z�P!jBp��Ǽ����l���tq�Ӻ5�垫/��m+6rhT�{G�n�+�2*�� �(�~LG��������}�$�T������;n=3 �E1�tg/ s˼:�p[j|����ݗﵖ]�U�������N�oE�q.$7�`��7�������P������'�_�X����;ʳx�=1צ��X���r-�矀K$!C��4�e�j1p��ygj:z%��w�v�-Ŭ.`��5Ĉ��O~P%V�KcR�!k��A�ːu)7�'gB��]lCT�n���j����3���	�\@�sϬ���a�M|��iP��Q̇@s��&&��-��c�~�)��.�������"�T""|����j�S�YJm������Q˻�5c�`��|CT�Ԥ��o�^�����!��y8��p�����D�@���Qߤ��e�w����x�O��-�FS��W8�y�fT'�A1�&�zGڒ��nJ;u΍X�6�FSJ�ʃ���K��酎U(��l{�?s�~]�&���/���ʑ��^|���L�����0W0Jm�&7O�z��I�M�=C�Z~k*�a��87�T���{i6�'�3)�c�8^p�6��.�7}`Ep@��σ���'�	�c��M�%�Ѥ��W���Ք�e�,���Q�%!4����[�]aV�
��H`����n���I�kzv�"��2���ָ:.}Q��8?����7��D��R�x��{q�3�渡�ΝX��a�Y�(��|-F��*�sݗ��m,}��v|��O�"��X���א��~:=p�_�J��lP��L�Gu[xP�R��(�qs�c�.j��D���u��Q9�|���פ{��c��H�_��9k/��軃�@�Ut�Ğ��@��;_
��yi���3��j��x?��Zp�Ԋ�tʹ�j����gr��;ez���W?��6����Ш��	���e`��P[NW^��}��!�sg�M���������Έ}����[E?�b*�����՜5.�aӸ6���u�!�`0�a��=z^���϶����z䲂��x�,*��ih�ٕ�uG��|�m���w�	��.9�-9������gy�T�G!���ۣ����J�]N����د��_�Ǵ��hu�<��P�,8��Xt^D\zTE�'g"���T����Q�nq��Q��୉1��<�,O����z+�\9P�W�����J(T!�
�
\1��^��^�o���f�,mib��&cf��.Ҧ������k+��PĻk�ռGq�Z�����;�5��r�\�h�A���;d5r�^f�V��S;�9����Ŏ���T���f�j"2_M���uu�#�z���?����a�f`���.��I��yع-�Q'�%�{K|��?�JV/Z�Ɗ�CIW����J!��� �d(�}xc{S�b	�^�+�k��L�ߌD��H� eW���q:2�k�:�����k[@-�v�>�s�>R*����}_��������u$��1Z��Ȫ��\�z�XT�-V�f����l�r����E���C�	���ً��_r�i�,��Z~Jx���WU�xvM]�	�;���g<�����ͅЇd?�=�3������ީ�}by@+�V���7܎�Y������� �v��g`�� ny��y�:n52']EQ�dg'
g�1�N����5�X9���j�d��8�ʏ?������%�D����I}���}U�|�w���vZ9ץ�l�*����a����t���zu������L7s�i~ژF��ѫ2#4æ��%�>^��Δ��i�{�@��+�h�r٠��V�e�ߎf��o�H|"e00?ЇO�LLu�\�,����ZuP�TJv�R��G�rj(���c��P�@�]C�Z���c-f�VȜ�X9`��7w�+X�a��
��]Աer�ݖK�Y�`���ȭ����	ė3���(ejb����8�թ��ĩr��rh|HV����&�0�X)l�8�-���Z�:4l�� R�pjjr^��W7�̭��ルh՗�ּ*�5�L�����4����A��E�Щ��;��<pG�hz���bep�*T0'c�_�g�X��kV�1����[�qu���o��,H�������҄�c�����34�3#s蟳��ɶeo��9�<�	��ɝ��0]Ǒm����	<��B�iw��RwK�%4r�S�����]FS��ߑV��{�:Ê�@2�:t4mp���������O����"��@s;j%�*��z�Zݼ�&2�J�ΌqgL)é�RX�l�1���r�o�ݛo*�2���.�\�ƋtPM7'mf	��[�|��m������|�n�r".y ����t������͖�g��X�kr'3K��{Y�(�[.�]T�n�h�>h\Ĉ�\�vZ�tշ��j4�ܲ��d���ʜ�[W���bv..[�*L��y9r�Cd��:�Ƥ���:�X�չ���.��=���^e��A)�$+
�xCK�kI���T�]nR*}�j�ٱ.3���[�N-b .�>b�j�S�{oc��t��9hj���qӊ��x��zN�cЙ)hwk:��ų�E'm̼]���kD:��w��^^Fhڷh�n ,U�1G����/�LԔ�67^�-̻b�ak��5u�;F�G�_,�)��`��N_�Z�\i�qv�َj��������	\��E��(�Qv�w��A�L�o��������9
pv�4�Iƻ6���-�5ոpj��6��1���Q��R��3��� ���=��_�A���U|��>.�c�nk*�cɄ^�v��t�xW��ld�n'R��	in�z�	��M�y�2ܩʶ�-}a��[�ŵz͠m�l�6�v��<[;:,�]n���ҝ����
ϕ�"U�t)w��m' �JuJ�7I��Z��YRe�;�67���z�V�V��oer%D��ȁdD�❽���\��%��}��S�WӺ�u��rM�/��~	�G9���gp�[�h�$NNՋ�;�7^�j�k�瑨�]>��.`��Q�-�ܜ'��X�6n�����K_U
�3�2Ws=���ټ\��Yc�/��+,u9]ûf�'Y�[s	=�$j���E������ӳ��[U�0t�Q�䓍w �O}�J������f��է�ϯom@�l����vݣ�t���Z�5ۉǋ�e�TܱD�nǏ��ow�~����+��f���2\�[.T`�s-�*^>9�ok���s]�\Eh��v�hJ�?@�l�+�*�4Ô��[�����@����}�y	E>A�����|g=x�}=~�_�������������_M���ILMV�("����"��*e�����&	��)��x����z���~�������{�}ݚ���d��3CHr���cSQC-%rMPP�RDDP�TW��>��"����bcET�ז��(�X4�ISR�DQPR�bR�D�DQCMRP6�6���P�"���A���*��j��!�hi�Vh�(�t�m�F����"�����%�"(��Y����������䂭�S(1R�W�b��*���&���������QCCC�Sr��G+�DU'�L�y��ש7��;-�c�D�F�,��S��tle>��,��k�7�Kp܆�;fM1�k�N�u5,X'7{u�`ݵj��ɇ،�C����B�bI�R6�HQu8l6)�/ۛ��z޷�����?�.rd��׶�
g�
����ڰ)��
t�5.qDy����y��++�l&<-`�ds<�O��ӫ͟^Y�;钨�L��F�����17ݪ)�q�����i�|kO��?f�Nq#�J����.�y\���SJ�z2�WnV�Λ�;ӆs�2���(�/ �	Y$5$d5�S,���=;��`Xd� �k��pֹQ�c�vqd ����ڧb���
}k;'X��]Z�@�q>���5��051S��{���?Z�5+�2��&5�V�2j�d.z�c�(L�,T)Z���v�`D>h݈"qt���t�m��B���p�o@Pd]L$�"�G	�����	�{"S�IPW�w�}g)������[+����8�m��r-�׺q���;����n{>�6�T�f[0z�q��y镛�o���U�w�b#�r��L��q����ត溣��g�01'2}͗&�����NȪ�׿#Ⱥ�� ��,yЛ�uZ
��!�)�5����np~ю�7��ʻ��/�
�2�Oz̮xj���^҂Ƽ˜��wib��j17�>�ņ�0���/�Ve��,���L�U$�W+]h�=::�h�Y��f�i�@�9x2��V	���ِ�Y�]��\���;�:�b�c��1��Q���Cl�}�M�U-���w�>��H�bt�ΆU�_����6.��}����:Уu�E�^^����y�x-�D�tZ��Dd�9�u�����j�
�y�إZ�:s� ��'�D�¥9�+.��_9��!�M�KLs�t8�[zhZ�2q�����%�J�`�2)���=n^=�y�+�T�������d9�8mO���sY\�6rR	�k�]�|mɭђn�n�9�0�ݎ(�/a��2�ƈL!�2߯�>t�1ݳ���_$H���{�1=w��X%�:�
�nǠLȐ �$�}n���b�I�<����|�7���Ɵ����;ӖƏr�코G׎��c�}�<^�Pװ<3S�ۨc���"J�#�����f�Ǉ%��|��'��Q�צ^?�5��ʼ�P�k�#2^�5xt���Qۈ��"�'
@�<�XΤF���\_��h���׳m����'aD-�II��U�>�䈇KS�F�b��}꘨sF)�-�s��q���1�k��a;�Jl�R)/o��������~��X�>�0��q�S�;G�1l�C5��4D����GV!;}^��7��iٜ��)l>�䛢�(0{�nw{ˇ���n��d�J�Z��lՂ��>g�:v�ᎈ��1 q�#��#7�3Z����V�Y���J�:�}��f�!��&Y��&���n��ج�I���w׫=���>ؐ��}�y�vf`�^�J�R��୿ ���T�	��J�w7�^׶t�On��ڼ��|�.;k���{�/m'f�r�p@�7>A)��`/Ⱦ��%t�ϱ\ᮢ��a��E�m9%M��x>�g(a��]�D���_Jw�y.�r�\�{�)�b�^1��;���Dq�~8�N��֋!���0d��`cl���R�)�vNu��9c⠱��a��2���7c(�V���2���/763�|gg.���l�r+�yWK�}n��/�]�8��wt��=�U��>0|���a1�zGB9� ���G~�/o����&��V��͘^�?����=+;x�:��E�^�@��e�+b�>϶Cp�C�wf�Mb�-�%�Ljg��Y����ٱ=u��X��*��}§ӯ@}���p�9P(��N�A`�	�[[4NK9ЖZ��g���g��	vO�,�vɳ<���zZ@�hu����{b��v�ww6���p6ϙ*��c���
����+��P͠�gV�����o� �[E?����f���(��~Ǭ��ۜ'䋤	#9u�=����jN�QV�j�&���s�
X�'��'cY�!~}������ƅ^�r�y���)��F'^�k�-l���|Pc�*�ϝ�1�xW��Ѱ��m��Ѯj�7u�,gy���|�`����~ �~����=�O��g��g-2� ������I�K�=����f��XrW!
���)H_��g�����ܳP��	�α|9LL�eX\Y��~0�>^�%O���%L˴��֫d����7L�.�e�N��eA�3�9��N�z͜OX�Χ�"��Ì�<�!�^����&m�����(+Q���Hμ9=ܽ�DcZ	J���$�]�OE�з�x =�5�|�e{K=*�h>z��]}c3�R����@]�C$�7;��o(�E��)�W(Ъ
;�e|�t�%]���|�Ϝ�K���D)xN�p��z$!"�W=�L��1��R)��&�}�
o�C���y0y�檇��z����^��f�~�WK0W�]��T��LU�ȣXo6�.j�K��V�-E�lG���1u�"=C��XགyW��0���M�ݹ�ꍗm���=/6�VK�"�I�yXZi��at;!�>zg�9L���ޔz���h�Q���j�oMd�r���A��U�ϹP�bA�&�c�C�c�ݓq@V �&�D����<�Tݖ-�4��Ր��_<tpTٴ����;m��[/��b�aN���mAy+���E
ǗZ�mŵ�GGNiN~<ෞ �c�pc���Yx��S9��b`�Me)�2�u���6w��)6�Z�iQ7+�of�{��$s6]�g������#4�5wdNF�����2!���z^��Lkк��zqKcy���~��z�"X� /�&��a%9'5������͎K�~^}��C2��a�Ʋǿr����>������L�~�r��������X~>05ǋ���>�vP�Ҕ�!tS��^y�lJ�S�!�W��y�+��nvc���^�Ƴ��";@�`G�![���W�h>���4(q�.�6��]��g���LUv?��Ú�!�y}����D�� �0\sH����Mi��ϣ�b�MW���%fgD���BP]7��f��(4��K���T9KO��l��<ă��� C�[�e�OgC��1�++#���ܼ��T�H9���h!�� �d��䌆�ٶU�-�<�zw�\p��@�;��p׎��9>�/e탈�[x����Rh�֟��o��z3t���;{`���`����fP�MǴF���D�B1t�|!e�FM��`�*���L�Q��Zg"�eB���N]�'����"t@�j���r��^���-�2:#�F�W���ua��s1�[��D���<ۖ�wSDB�U�[<�ӥ�y�"��F'���ޚ��q����8�#ġ깝a�x7%`���\�/�q���j̒`X�����ۙ��yu�rW(uS����4k]rRX��y�Q�~��|+����{ϫ�/�1P3��>�N�P}��n]z��tB��B�,V�ʝz�:+;g3-������9�a�L��lm��s9�# :]"ٸU���}r�5��7��W5(+=�W�G6�;<=��]��|�필T^K��Z���9�2��OQ0h��,�y�*�� �:���g�$�h�ɬ�w�="Ö�ڈ*@�)b8�\
�v��(�����2����u����q�X	����HqˤGj��J��s�VW�)u��8�ԴN��Yׅ�o��k���H�t��Й�ޏ8�D�r�H�*�4�حgI1w���@�Mz7jô�#�h��� %*�k�2�=�k1�=��og*	o���Lv	���s#�� _E��5�TLgc�������Ԁ^G�y�m���x���IO<��|�޹��u9~��=B�J����R����9.k���VY��"�S�M�/jޯH٥r��Of�S�e�_��5�S��kC���m����W���zt�lkW2�%j�r��F�8̭�	]�EiM��Wt��Q1\�È}Ў�D�%%f�w�������W�3a���t��}|�#j�^m�g �gQ�Ǜ�M娮��1gV���2�zH亨m��9Cݸk�Q�XZ�V�@��1��.*��r�-�;;7%�gZ�\ә�e��3�z�,\���ȁ�*����d6��^���hsw۪1x�﫯ƎO�j�TӚ�@֬��rDy^���Fާ59huv��v��0�=��J��:��s��:�>ǏH��F �M���vַ��zxX�[�FoQUe���q�W���������*y�T����/�׺k�0^�kK���:d�>�f�#saC5cKO:�4MMq�أ��jн�r�VȽ�T,����i���������5�NW�{7�Dk��};�A�oc�^��_;�}�������[���b�sL���4w^�Ps���2ï�6��o0]v"1H�����l�-e�;@��[�zu`��/�ȕ�R^k���g]�6��F���ktN�'���f6/X�wk�uQ{���K0-&(U3s5�4�U�޼����+R�6&/銖�pգ��,.ۡF;�f��)b��o�����ǚ��S�.��3���7���&�Y��>wI'�'�{�>��Ɂr2���8�4b=����_�ʶ�+R�l�{�vVM���;`�@NP'�����݊�ҝF�R��,�ᢴ�Pgq�w������P>��M� �}7E�@~�̱pxَ�U��ݗ��r$R���
��J���g8�5�:X��~����B%m�s[��-!qOs��w+�?$�E\�������z�]:��EA���ޘ;��2svFf<��اYV:!᪑�_��WVv~�%mZ�\'�~N�g!���ףt��"��ћj啁��aw*��1/�o�]
�޾��"2��YC�	[�q�T^M�9�A����b�;�6��6oD�����w�\-���(�#�)N�0�s�V�)�MvX�z�Z	����@��0�5?����r��H׹��{��^(�p�kS[��l�Т��.��j5��a]�������f6����$�����0�a��&�<��*�fc�nե�!d�S[Y;�������>�Xa٪�C{�ia
��<��ܠ�]�v��Py�۳y�	�z��t;�o0^�����h��x+2��[͘l���K'u���1X;���"���C.��Sԃ>���?��^�F�����כ�g:���o+��w�{M���.�-��NBَ�֦f-�w
/7;}3�j���Zk�_�l,������tǜ���L��Ŭ����8a��]�|x���4R1IwO���	�k�3c�i�K����l۽��~��j�"
�P�5��S��JE.�s�IP����@�"�	��ӳx�!J�iH�j�����87�M�I���˺��9L�Vr.22Nc�#g�O��/�Fm�C48�'F�w�H���亼�M�I�wWM7Pxm�>�we��{������q��7b����{۽[��]��Lښ��{jA͊x�A�FGL`d6y�.�M��j� �3�0gfA�Kyf�y�#Q�� �����{�C{�B��
��E�oZ��y]L=fX�g��m���9N�O$�j�"�Se<"�|�����y_��LJ�M����n鲆�P����%�����Պ3��;�KZevI&1-˭+w��"knV���I��0�#a���Ndn=��2ns5���J߿U_�_}�/.M������U^���Wa)[���g�)N�u#��q�9,7-����q�[�<Z[+��� �W�D�+��K9n��^��k�ۢ�{4g�W������q��߄��F.��B��3�fN�H�ٛ/c�aˮ�^)^�y=4��L�.�u��o�[(_J��V=�5!��t2��H��!O���p��ݪ	��#�2$[��\�A
h��Ecuͻ;n-������6;������|�dQN8��.[�71��v6����8�3�Z2�t��wa�lEՔ�Жj������g�OD�a��bf�)|z�7���e΄��}d�
�=^�J���T�%� �:���U�"2�k��Y[�s�K���?�e��S)wIɽ�yr�k}�^3t��'#5��5�L�����Y�NnX=&�0
�Ha����E�N}po��`_���fVD��Zuj�7m�<��L�7dTr������dqUN���͊�R���w��܊յ'����	^���Z7�FY�F�Y���3�{)b���m��-j�i��Pf��QÝ��[�1�z	nih[+-�Ó������=P�'Ã�]�dT��ᝒ�D�S�(&�4�r� ��ǋ�0AA�Z�Q[�������J��2]�����o8�źp���e����9ـ��`�2�ħ�f3����I��a�V3z��%Ǚ���s��Q]�q��'�����$*Y�]�,q�m� d�-a���:Q[a�+�[���ڰ��\���$��ss{��ưP�غ�Jt��5�����"��Е��Δ:��]�/��3V�=�R/t�Yc9��]���<ړ-��ŋ�Z��qڒ�YP���[��ǔ1#��N�ΫU!��o�+�U���jY˺�}N�&�(�U,P��[����q
��t�o�l����7|���J�ͼ镒�䅮����>+��F۠���a�mۉ�eiYb�c�*��%g�iL�'����"��&�<�9��)�Y<[��%�Tb�I�	]ܓ����Ag��H�'�j��V��{�۱`\l��Z��T����pnM���]S�֘��JQge�P�����PG�n`qJ]e]�08�9�E��.q�}\1��BN��#�TB��ݸ%s;��њM��'S[�o[g�q�c�a
� n����(���}f�:rvʆ�In˙?eK����+|;Z��T��+�����v�U�s���z��X�����ѯz-��J�ȝ���Z �l�쾖pF�V5K�����Yi҇�d�-�*��)T˹t�J�t�l��Rv�zuoN�73�+�ׂ�lq����NZ����X����fv�-(d("�����Χ�)u�Ĵf�7�N9k"��=��ڞq�e̫Ԙ��:�,7Zʾi�FB%r�{�o��ё�
�N�]s�uǋ�$��nK���M�����M�<�5���v,)db�t74+�2���E>�W+kS粴i�t�բ�@[|y7�"�ޮr��U@��A�V�F�u2���]�r�לOhիU�̛�Z ��*�c���Ž�of]���T4w�RD��c��Yեn��E�(��)I�K�
��x��6���IK[�]�/�<mulTݺ�9�e�d�����R��1��5˜WO�j������I�A�(��꠸^% ���-̥��$��L-���_]�F�#lTB�nB�Mr§���U�GU�t�F6w���[�=Jy�)���/zJ�>ר�t;Fm8j�pޙ�έ�곢�3o��C�Q��f�;:oG�fା�-+�̀�z���,�,�MFF;D�*T��z���";��;���9�G�a���>��5���M$Eg?^�>�o^�_��������?�?��b4;��[$(����<�PruAAE4PD<g>?�O^�~�_������~����?J}�G 4L�AMP4M%4�T�DIM6ƒ��b�����*��sP�U'$�m1�*bf�&��b<��������5�y��������h�9.�j�J"
�̆�$��󚪀��Q45QUQD^l��,-͹�A,CT��Br4II�Q%D��i5E�p�|#�5�CLC�ѣQ$Ei4�40�*��=�b��lu/<�ኊ
JCI����[:=\��6���9�^�1Dh�8MRO�Ah"	�K% Q��ԧ^���v����g	z!����<����&5�aV�+4�G��G�Ţ�b�����r�!��>*�x|*�¾��6z��ɬ�d�ʨ�3Snc��K���U��rH]b�sokjּOuf�rvn��ލ�ج�6�1�~�"ϵ�cޥ�����T�ݼW�Z�C��-���LA�FGu��t3���K.�Gm�ٓ����)��5����O	�$�xF��,�iL�⃊�,o�X�O=�5�z�p�z�ں����D`gd#dN�M��^+Vn*�=�������]�#&�CG�P��pn&�ȹZJ�,ע��#B�槢.�#N�^Z��,ܻ���l�_�n~��O�ٵA�N�ME��=]��o��xm��Ƽ-)U�=rv��\ߪ�k#�z ���w�`4񮐻��v��pCV)O>!V�W\JT�T�W#i��� �QZd��W ���Y����+J��IX/�ĽI0��������N�c��gV�45�	U�N\�̇2�w��"��ˢI�΅O9���}�HWQ������x�X�J�f��4�7��p�7��E�]���ٳ&��[R����w��i�Ff9�;\�G���3/!L,�s�-���+�\����I�͕��{�?/�������#��z8�@�~[�<pSŷ6y+�*EsA�,��gg����JclE�Ӎ�PY7
��ಣV��I�)����'V��X��*�\���Fw;û<�y�|T�Z�+������>wv����7Fz�Uݝ��}��l� ]&�|���t7��lW¿8s�{G�� �
ů�z���c(C��H���(���e��I�F�9~�I�&CCԍ��:ʚ�hs�a�(	���?-�݊��^�{OP��3��a���v@��Y{�ƞ�[�w�|\ّn+��=�1��m���;�_@f��+sѱt�ޮ���fЁ��vqc�y0�l����^ �����F�b��q�Y�[�j��N_��A��tS�!�pwB��Urj����L���NW�י��uK�h�^*�k˜��*j�^:9��s(4��K=Of.p�y���L���6j9@��-f�S-�;�l�O@P4��@�Zd���a��}�Zm<�߯��N��,m�AG�(+;_O�8�&k.k�R�T�;8DM�R��e$-t���ѷ�K�1�D樟d�{W����� ���|>���f{��͒��>w0�ٴ�0;��*�^�6A�q�h���ھ�:Ζ{q���.�|�3uY�b��Ge�m��S1{�@=��,����8�#�ysNdPR��fgS3�cb�ȅ��w�#�n;dk�W(E#B�v��U�#Y�pm#�����^���5��L"��p�|�F�F�<��`΅!�-dP�;+��^D��K�;-���&`�^n
��� ^�F���ɶ�Y����U��}��bNn�iם���Y����b� 9g%������s�|6{�q�&,��s+�(#K�W��1sl���n���r7��؉����u�}���Ggh_��4QJlJ�c�v|��A����[ӽs��fR�ǎ�#C�y&b4�j����T�T���R�U9;LJ��*�_ggl���pT{BP��ۊ�J��U�.�����і25�!q4���٥�ʽQo�X�s�D��m��,k������0�L���^W0�\{K������U
�c�3��E(?�)��Ϸ��lu��[7��pVDs��L��R}S2f���|�wJCa'�W�iC�j�GW
R��䳫�5�~���{�	�}~7����wyz�F�V��亼�eNS�<$�%�q��N��Ѱ��Q�iý|�=�f�-v�ë���_TbJ�[E=�� ��cTrf{��Zz��y�I��	mS�y�9�F����:#�/�Һ���Mu>��ڡ;rm���7�/,��ypH���nYK=�ng�E���h^nE���VH0�N�Y�8�5(^f�#�v��(P�d�ޚ���ι��)���w8f��e�` c��j�Oy��jW�Ñ�$���#:���#WunI&^N�5V
�F�:W?g�|=n��~����|]��+�W�$f��g^�ṃ՜4�1�v�a��Tm�����9��t���������p��p��ͧ5�}��/��Ig�2W��mԍ�u=��n<�0Bc� +'n>�ɷ����9�|�"��K��dl��\�c��!���um�!ݿ�ޝ�/=�/=�M��]��{jښi�;3��6���m����EVyC.x<�B9��v��9j�����[�-�Ts62�5�S��_��u�4l�_�_8M��	�ȥ���8ٚ�\7xs���q�>o7��i̮��ps�B��v��M3]EZ��r�����큦�cr���m��׍���.�t��3�/��+��R R]�y���� Opw7\:�.���t%6ǡ�2�ò<���"
��d=�[˥5��b�Y��g�Q�3�o�u�M��
X?���L5��#�O�M&&���p]�|��YӲr��u�6��ԬJ�[#g��7�4s8#y�*�E��d0k�&��y7]Ί+�S.����7Cz����������0��*n���A�{�b���mqXyW�ɟqn��1���6�zלZ�KC�:ۺ�z����*�J�h��m�^[���'�{��I�|���L�d|A�$��ө�����R���n{�v=xH���)���wf�ݑO�TW
��wu2odtS�a��t BQ结@D�H��Q[Ū�v�@�O���?nP~�l�I�ۼ<Le)+������ ��k<�F˲�=W0�o��xCs ���D�U�QU�4���n��^#G�J��$Զ�4^]pl*0�sVw;���aZ�<����hӚ�)��q9�Q���uW����믩��2�gw��ӛ#�Ɛ/-M�9�j��0��n$��Z��d[�lVY�U�'���ˠJJ��*����ڹ�M9�T����.8��ߒ��{	.�+׵7F?��#N����B����J
�|���&��F������,\�XZ�Pɉ����B*�φ���:=�z}Ǌ�����<��D�N�z��|4�6�ܞ
+����3g��T��q6&���yg]�p�[�1��&�u�0	�<�� �1$F��ޓVSo�1�t&{ޞo��ʾ6n,������K��2ُ1a��S{����c��Lf�P�X�W68��٨��6�WF�Mwv����$Z���lCc�>a���FY�h6`�x�ˉ㯓{�8ůVPs~����\�3)�f.r����q�<�{��-O;��_%.2��r�n�t3yVݞ��c�7;��A����NF�< FI�]�G�Im��d��G�MIۍ�CY	������97��=��ĸ[�U���|��ggg:5�E��t�Ŗ�ku8nI��ټe�[:8i9�[v�2>@�G�����[8з�P������%,Gʆqׂܳ][ ���Ns=���`'e�X^
��!�������������>�z���6�wF�,�r����!3���VY���
����GQ��1f�қ�����9�T9?m�k���g~�n28��=M������~����+���'�VI���BƧ��Sud�t��u���]^Ԝj�%�ה���>�k����EtP����V�a��5�z����@mb����>�q+���9����xlӷ�z�H�i�q!d��UuYx��CqzS�z^���W$�q�v�����뇲b�e��7�n����ؘ:���
���[�2VN�W)F�JS������ɚx��cy��q�׫U͇`g�� k�U"R/G�=!�B<�{F}�Ý�݈~!���v��IT�6:�̍/ �$*c��X5_sf�2�+N�&G]��St����ϼhk�H㫨�6��napB�@�����j��|�~���݇���q��r8�=�wr<��\Z~y��k;M�ޅ��g|��kfb3�r��o�ە�O+�:i�$��A����w'���e��X5z�]��O:�$�ʼ�2ڭ�\]8f�,��Wu�џ1y���;��7����&�[�'v�!�Z(�������:��AuT�7@as�Ao�}���t��{]�u�F ��G`�S5�^h�&\%ܻ�3'J���E��gv�'�=b܆���#�dF��~��[�V��F,��QS��5�*g��9����y�$8�(�m�a�O�z�Y\���;-�!�f�������,��o���.n�s�@�9>�K�\����2w�o'�M��b��h%>;>���.��m
Y�rJ]BQ2���5͸xpֵi����._�[ �l��*I��2S��`�@x\w���5���݁�_R��~ɓ��}������վ���Z��\���E��~��=�V�$Z����7��L p���G%Db\������<�'T7o����џ�j� j��u�i�s��+VvljJ�(�ñ�I�z����VD��c�{hT�܍b���u{8(���v���t��֒sФ���hk��w�@��Iי�8[�t�t��ಔ��I��l��{Ng7k.�ܑ�P��G2񦫜)�9w�4�GP��9������p��������w���v��J�bk���e��\xX��w���E�v�r�Z2E�c��>nGX=���yD\��K/ϑ�މl�2J�2�DZoX���gL�7N\�����;r{�Ittߓ�E%�8�=ҡ�n�vd"�B�fSڒ�OB���m9Ǥth�9���o�"��L�߯����f�tx��=S�W�~��ܿ`�`�4��:�<�d�hV\Rz���t�6�;��=QҚ��c\\Uj=�}Rp1��{#|�.��X�J��W<�T�y.�=S�љ��b"���Ca�u�a��z�AS�f�eV��z�Z���	�ȫ��;�Rk��&��0�a83a����#�M�N���~o�ʷ���:�s�H'�(q�b}�}�l�<����+�x��x�s�3�W�ul�.�����V��J4tެS{>��o�u�C˨WW�#��ء;�}���f���`_b��
�S�+��K}W�C�yQ���{���i��pN9vM�B�vk���Ǟ�6��`���4d%�y�i�ىKT�Rf�u�v��⃲Z��7������u��K<i������� �\�v�_����x5g9��Ά(<j4 i�U��"vx��\��fE[��<������.��c�7dJѲ��)�b�y�iW���m��x7�HD�y��C�;4�$o]�p.k{ l0�hɷw�17G0$Y���6���7��ެ5;Ϟ���g?��)���̙�lm�j��=��l3���A~?Z���-��Y���(U����Y�mmv�N�^WfB]�yK ���,�PG<��c#�*xNRi���J�wuvQ�$��ҒU�J����W�~��������10H���`h����1y��q�d�΂�5B�%%e>U��+ӻD��n���,���p������O|�x��5�	.��)���a����Z���ˆ:c�����@���r]sA@�pUŬf�%|��X3�ȕ,�Ѵ����q��=��v�&���A�?�#�H�2��l���
�z�]�:��
ߪ�v�ݒ��.�MѡX6�:y��6
�����aȕ��Z��2U�6��*Sx)��Ѵ�ָbW��v��)2���뛖�v'[�;�Mh��|��F���{k{*����QV(Tx��D󮱷8Ϋ�5�%
쭑:ޕ����)�������c���6E��@*-4 �,+���}��4��)ᾋo#i�QDp�JN���R�
��yS4?��Zs{+�0	Vݬ��
�EG�Q�%!��WPQP�Np;�ն6�'7��;��A��Wo-��^�<�a�7��0WG9��Mf�K N-��x�JV�=��V8�viq���>�B��^SՋ7����L���X�V�ʴ,�
W6�m�2oe��t�$n�����h:Fl�]��V�����w�;�Ee�� �s�%f��خ�?�p��%PZ!zx��p�ʟi%]m��{,f��]NcwdL�a�}��h]X�g��������{���EH�
�������mf��;(�R��*��iWE�{��oW$�(�d�6r�k����R����ؾ��W��ە�.E�(p\86)���iX���`�h�t�3�9f���u��s�Mo\�^�t��ۭ螡�5=�iV���/��GL�Ų�%|�G
����|\MU��.���d����c�Ѵ93����`mg
�IW%�sW�l��&H˵$�x]�gU�`�;Nк����92�
��0�˼�� �7G=Y���۫��v�-��tF��]�:O��=��$Be��I��;��X��Y��/-��m��QE� 5z�˷�S��ǚ�����;Sܬ�ob�ueA��Xyst�u-&F;���"g_�`�i�,(�Az���)4j��x�.7�3��<s����4�ي�Qid�Ea\�vٶ󾹯��h7��_m�L�=����\=��+y��%���f��zm�c�s�3�KV�;�d�^Z�-⹗r�EE�l�Twx��PG#5���;�ޭ��-�Ћ�J�}�(���Y[6�y{s/Y��n�:�N���;�C2��'|���E�'9�5\�+:-�{�wʭe�fャ���][�]qE��3o^݋�Eu��q-�J�پ����;��mLO03�߻E�n4qi0e��\�t
C�
':ѾU;^L]�ս,|2�ާ���?�1B+ե׾��/��}JٽđOZ]��n벮o)�#���E 9p?q�V���ǵ�J㳨��Y$S�[�Y`a����rŷǵ2E���	��[c�u��u%�T�x������.�ׂ�gY�����x��bCռ���zz����U!�[����7�jCt���\b�4i��ֵ݁om�F]Ȧ�o1ue��A��-�@��c��6V�U�(����H�=�-���B�Y��&��VA�a���y�8���x��O����@_S
ox׫CTig9��|}�޿������������U?�6ˣMF1��~^K�&!��h윔�h��9q�>�o�������~>��ǯ�����v)�r(hZ��(b����������h�:^ܐ�!��yE�&���6ƚJ-����iM!�ڹ@�6�E���EIT�%O& �M:]�6-�֝j���9)_��Hh����h�ժk��٥���4���ONA����y�IKI��MV�[cG9��*��&�9�)�����l���[k֍!�Kf��Y4�N��TP�S����mHh5e��:�cTRV�y�����^��\5�D�(F���g�c	]�z/]_!�Q�kvt�h�r�J��|���	�]����jt碥�}0��E՚���7X����e�C`Pl��B$vunFy�
��ۛ[��j��^W��o.T^O_�2xc����7y��qO>��}u@�(7�ѯݯ2m�/������F`m�0���d�ʣe��4rz0g&�G��ΤW��	"}->���l�Y�4���!�^a�����:rM^u]`5j�A�Ӳv��Y�QBS��\�'���`�;�⥮"�
�"6M�0,Ã�}//���?-�݈	��S�O����cd�enSD>�ҙ���h>��W��d���7�u1�o4�n&�P��	mEkv�wk��_Y��!��9����j|�^4��F�Pn-����ɮ2k���$����掜�K��_5��;���>�s/{|��q�q=����$"^ ��;\d��yAlu6�Tq���Un�7}�ǚ1*r�r����M�Ii6�ʆ[(�m��Z^���m�氩��/�2�[Qq��W��
U�q�Gj�6<HvR������<�=�f��K`��+��)S�b��|���Z{{<)�R��;5�W�;.��N�mr��5�-i���P�>Qw8��}5o_"����H�D��Z�M�1�� ���-�]�)5���\��^�z�w�EW��\:P�-��@�~�
����9�tG�ѵ�
�C0�M���M�R�y%^�r:�?tE��-٢�oUѭȭ��O��l�Kg	�H��0_.�Ԍ��x�hj�{;Zw�g�w}��u*4�T�=Sޅ���H7�NQt!C�V�wA�mQg'���3��\�ֆ�g\v���xo�� 9	���6G6%�x�Y{�'D��H�뮘��h�EET��kY���{�Ԗ�먯�<|`1ݵ�g�x����rQg�7��_)�Z�E#�t�v�w�+œ�(;�U"Ky��ٱV�b�aBu0[�*DGT�9Qn��*in�W����-8����z$�޼Ȭ��_�b�F�8H�����=LudNqvu9��[Hv̾v�+FL ;(f�m��o��@��`�'�Ё���qR�V���ِ4>��Y/z�z8�;(����Nў��:�s?�'�:��S�6�w��O��*ɕ�e�d>Ԥ���S=���՟�o������;����W���XYג�5O���=�^f�l
��w����ˣ9ސ�T�z�먭�h�bZ�J�s\�����P�[�Y�@b���y)fn��������y�F�9�nNp�нm�k4�O��L��h��W�]ltiC"�_Wތb�k	8ϱ=���ah�5ko/�}�xO�#N���U�nb%Q�w�\�v��{xoS����@{�O鹻��$wYR�'�pT���i��Ì�i�ZE�s �=��
�����o�ȹ\�P����aGI�-�M����i�;��3�k�سwZ{�*%��g��W X�`ϖ�S���[n��U< ͷ�ْ���o
��;�lɠꣵ}�-�� z�BA&�3)���<�2�c�{��>.�V�E$_zH{�+�nDH�� H����M]rQ������F�wA�5�%�C+G��6<����\e�v|����7��|�6�r���ףQn�б1�;��ᵪqn���B�uё��}��ǐD�������F��2�������]>�~j�=B�*����#����ۢ6��Č��[�\[�<��*`�츶��Z�;�L�wf���1�N�v�%�U�"����NY^cAӥt�=�&0���'m���-�}��v��lM=�U�&mm���Fc�'Tz���y���r����rR��WL�7�����E�<sf��:!h��d0�,�ս^�*zJU�Gh��[[�����7=Y���Hj$�	]��ޖ��3}��sͩ���Mŷ,��5D�Ok�9nN��=ԬJ�[#g���{����x�]4�q��eՎv����S��s����Qs�c�Q�l1�*�u֪�Sg^�[3s"��f����&�b̙[�|Lv	�"��kD��g;�gl�_�������ͣx٢��7�b$�7�5���ܑ5h��u��"����+��B��I�z�76�r2��jq�����x�K�OH��)ʍS����w���xa��t��rk�1�=Ys�R����]�սU㝫���B�2�i9��%���*E[�p�m���𜞻M��G]�Ќ��+�)*��R��4���������l�!���}����QU�-�bE�5���M�ON��Q�4�<((u=�y�7E|�{'J��J����r�Ϡ� QJ�u^_|��A�2s�����b���Μz�(�څ�Q.Ժ��i��S�x��U>.��^M}�BӬ���Q*�e��}_�t�R��w��(��ۊ��ϫ��.�k�	ˤs��j��ĥ^R`O�ʶ�Yl[F�e�QU����l58� +�M½�%(��������%�{��t���p��:��MӨ�x�g�:+c���W���SC�����f��f�����SOf����l� �,�F���:�!l�{�u�﹫X�e�w?��{OQ�NQ2��#㭰º%�2��z�Ue�}�]��2��|�,+�Dq%u]�M��K9���ɵ�0�iCy�an܍\���z^:N�L,��ceO�v��o%�Q5��T�;��ǟP�d$�kc0��x�.0õ\���T��[�د\�V�ё��m����{���%�1�A��gA3��}�0��϶����Fg*���L�n��=�1�MT֌�t��Y��Xhf��vm�Y�"Ҽl���	�Xc+�]�[�I�J��x��K��r��q��rohg^pƌ����X���÷�����,<2�M7I���aux�n0�\�l֍���As�>H��!��ϮLZ�c�B���+5�r�T�$�կZ�{6f}�~��oF��;�F����sD��<{^`�;�9� �t ���k�����xn˼��=ѷZr����&䬄/��#]/L���K������Vz�G��լ�j�u�ׯr=ܐ�ֆ��q+��m,�e>��Ӝ3�U��tEv[8T�k��d�M�.!_P�* ��ǲR��l��!M;��"[�B�ߍa�T�iX�s{�g��C��\�1�n�q;���3 ���q{vK����)�z�T���7��6E�l�5�S�Wy��J����>���PT�]r�N�7��u�5+Y���̎����������IJ�θ�GG���������Y�|�:b�s�nk?)��zD�]ZZu�.W�[��G?�UIr�^����:+������=YDKr5O���n�����>�H�]���d7��Mt+Z��љ![�P�k��a�.Z9�^$6b�]���ջ���S�A,�THj����{0X[���|�mow���$�	g�E�`�je�=���m�D��*�p#�1�T�9DZ���tW�����o;�zo��p_G�Ȉ�������;�w�ߣ`S�!��~��}��;�:�"#��S~v럿���+���G��&�)��H���ԆRi�z8f���%B{/T�?q��8ZF
k�TUlvVv���UR��r�H��7�7��sv#��v�ܘV`�Ju߮�A=O��o��ڟ�#�e�#�1��9�`G��6���1osZVW�=��x�wr��XP�m���3�:F�i�y�dv���w�`��M�y�m���u"�O����/���}4������-Z{�ቆ�k���_�<�뇳A�Fת��J�=�UWT��v:��#�+"z5�Cն�1=k�n�:�}���g�]���=T�Dٛ�,�_���Q�z��Qk�d<��*-���"϶��{X�ب�J�����)_~��k�r~s�C�~	}+������FY$�&��o$u��&���i��P��2zNһ�������#��ܝ�[�>��Sٹ�7j�bP��u�%�C[�{uǳZ/����ƞ������EER�][+�"5o*lt��]����7+p��n�7���+rε)i�Ӡ��Ş�"h�7����������a��Σ�!���۞�E'.��RS�Ư!�me���θvfW(���Z����ƽ�O^���![���H߹��(�y2
�>l��V��"�Y��#o���w�mB@YpBǤA����%U�h�ej��5��q��%�����ŷ�Ȳ���WHU��G$�b<�}g��*���i��$3¸ >��ci��[��5;��w�J�n6{d0Y}[�"}&<����Ŏ������g����������I�@Z�52�i^�Kl��5���+���s�I�󧷘(t/z���s�:���R�]["���C�
5Տ�/��;3ޕ�������������7���H�.�W~�5N�wF��g+Te�����t{��e�q.�(r����	E[\
�M7�48�Y/y�͙��;q���5��j�5ڀ ��,ꍈ�^#cy��n�������^n�6t�h�Y��{r��%Ӈ3��mo�a7j�{M<
��q����Z�O���V���E��ٸb���^Ď�:�4�-���v�g�)L��L���K��i��W,ott�CC�;f�ԸIC#���w=Э��	ˇ��I�:�U��@����5�����=]�8vӚq慂�k���tG�k.���ں��n�4)��6��^-�����u�u^Av���Byqi���E<kxC����=ܛ�v�I��(�l�6r��>�q���P2���.Ƽ����;HUT5@���)�v������C���ݎǌ��+�R4Lz�m]D�7����;�D�Dmr�1�Z�9:�Tܿ!'����t�P��H�)*��l��,��e}������4�n��x
��<�@�\�ZLzF�$����v.��٘L5����w��)��t�өY��[.WX�W�ׂ�z��z��}��E3
�̝�lAi�������ly�'��?�gTn���.k����7�!����޶���ޜ\wI�~�f�}p�2�*�W'�f��.Yw�;�;���FΠ:���G����O�0}�R��yi��|�|���7��ښG���o$8^�+q�]7�)	X���'J;ӜBw�*%�c�9Cl[�S��[R^қ��L�5��/A�ų)�䤦�C{;�������L[zzvK�KTR�9Q^����H9`��E��������W��C�o�Lu��R#kԩ�b��jZQ3%G�=̻u
���k�[�����!ņ#�2���A�l��o+�W�kG/��ت����\�6v���6��<4pBP�֢���2������C.�m9�fު[���Y�u��Xv����f�vt;c1���[��7�L&'MV�Ln��77�B(�Z̃��+y~���p�s���Ί�k�ly��N�� jS�|oZ�޳��%�WJ}�Ndd��I��u��������q�5��Qy�]�o�:C��h�GFk�����_�Y��\ꞌ��$" *qe���E��������*���=T��B�W�vز��P�Tj|����3\t��ف�$Xh��T��t�R����u��"^{�w�;���=�;w>�n���	�M����<��:��5���a�<��S�v��z�=ܠ���C.ux�ʉ����4_^,��_cӖ�Qv�o��Ga��<2=.�ϲbt���&�GE�5��8r�Z�h􅖔�����W��ci�AFQw�����35�ȯ�>��w�WU��n��'��DDr��!��yB�
1���И�v۪����ʊ���ɵI�7�o���ݏQ5VUN9~�Sd���D����]A��d=OX��k������eƅc!A���.ĳ'j���?����9�����3i�ҭn�0�*,ͬn��gL��.������{��� F��(v'bsX7�Α���eA��Z��ʃe��gjn�1u�ȉ����`�T�v$n�z�ઉ�!�T;���6Xf�ʵջ{�5�*�:��06���c:�Ph��]ɢ���R���O���W(����/[VNudG��|��"���[����U0���aZ�<��"��\$�$��w	���4#����@`��� �.F��WR۫t����[}�����5�VKS�u�,.�:��7o&�h��M�uf䮺,l�r﯇.*�Š��l�;�c��������pa�y��P�әrxOe���\OD;��h)y}�u��/hJ�fk����FL��[{B�.������7Xj�k�H�K�bIj�Q;��sS#n���W]pf�K:#)�fh��]-�2��	ջ��cl�{��C:�є�n�n[�72�Hv)���&��m}�X������~�N��\�[�p@x��J���1T��7;t�Ƿ��p2!}�ǹ��r�V��Z�f�3Jd��^:����M��>r���%A�GA�]����[�UN��1^l�Cy�q��)O�������zY5�5w#�lCJ��sz��̦�1�xat������y)����i�g �gnd,����� ��tlNJ�N m�ܺA�Ir"(��ͻ
[�O{@Q���s�\��-���7�+%0��iefuC״k�1.�1,�G�j�{״�;/14E�c�L7��m�j�c-hGvh8XQ�m���%���ћ3^t��[����!��Y�ǜ���mPOF\���]� l��qT��>�lu��l�z1�X�Z���:+c�6c��vs2�4��S��Ù5�j��
����;%llwX��qAN��0)�1,*f��iD4����8eŬ���]Z;��*���o���?�Imhk��tS��C�0���+��|G*�[�+39M�{�G��r,�jn���L|f���7����\r}w�5l��m�-�ŵ#��E�!=a�f��ޏ+��|*ة6�v� /'E�\�U|�J$���YC3CɌ3�[��ri��y���XjS� 6te�9�8�0�+����hB��̦�j���i

(�6�ACl���ǯ�����~?����~==���F��H�5����4�h����a4��wf��!�V�9���>޿������?��_�AIs�������,Dh�5�h4��476(�)*
�`�a�����69Tַ7�:���-Z-�1�E45�1PӶ����z�xN�y:j�I��P��Z4%U�bj�y8�5Zh�)(�]�A[8j.C�NM��ڪh�lS5�f��$Ӫ�D��r��UO'�k��N�B`����ͤ61͚��=�˘�;h��h�jd�5Ey�rv�L{�yPP���1���1�4�\�@�(��unnQW1��/�i�Q͋�kj�)n\�-��kK��Tiu�LEEi��V"��kK˜�1�
�m�6��o|�MZ���b��̍f�!7wOvH�
عk�g�[�h�kopk���s�����ks]��?�J����?�Y�/MIw����z'I9��og{���ig=�S��U7M�ө_�ä+l��m�B�)X6ӺzGF���;{zJ\�ȥ�0X�<z�6c��.}�w��%��g̗�$�Lh��5��IQ�r���-�Z���g~�v��� CT���i�,|��H�T�-��<��L��E#仐J�y�aOܽ�����w��m�#��θȈ��g����4�y-y��zhO9�Z2�ۊ�Զ��v_�����E2`8�f6�VQUI��&��~�]9܊�#p��}o��6�����+���x�"~���<E�*�ܳǹ�ĮM�|c��>�`�h�-���Z�(�jy���������}_Z�1Ӽ�����Ap�@b]��t=�	����ƭ�Y�:�S?sD������p���j�g�9w]�Dk�N�o�}���.����/��JK��&��2�'���Oh�i��v��k�� 4övo�!��l*m�e�,W�`7�k���}�|�.gaMn�����M�	�N����ۻB���9|.[h�a�����������Js5{���=z���xb*��Ѩ����XL�z�^�����λ�-L��0����lE]v�u��g�z�V��x�v2.\r͘����M��9�]�����4�jI]��=T��;���1 ���2��/�)���Ľ�@NB��$dٓFuM_�#���ϿW�~ê�p�2�W����u�ܛY��3���%������ve��:��]{J7�e�:ٽnsPt�y�x\�!@�"��6�X�*�<�qj�5�S�봺s��M�1��8�������A�u��2�-����B��:44���5�ۓ�z�⻷V�}Ͳ�KX1Q!��W�T
�f�Oߴa|��,[����`̛�D<8��np���ᶃ�y�^�a��z�AF��+���.�gWoe�bO*��W���W���������0�t�j!m�l3�#̽x0�O�浽��͖�톖a�WF���cC82*h)r9��r���')$؇��d��|��V��
��T��P�!�S�c����e�p�_tA޼Y��t\�8e��w�PՁ'�����f�mr�c�P�+��S���w��_�����/\�o,I:ݲ�c���G#�϶~����>�]i�r�%Zd���&�����n�[��4�M�[h�Ua2��[�ÃQ��@g%%�_�����;va�_\��ޒ�D����ۈ/i��=����b�nh	E[]b���5!qL�U�gZ�#��tϢ	�۳f�²}��Τt3�x,��-F��נ��n%�Ul�V�\�3�ɣjbr����ṽ��I5�yEG���@�g@�Ra���6���R�]D���U�#Y�7�b_i4B�����^Z��M��3�ЂT�����p�p�������{���f&.����Πe]�K��-H�&���gJ%I�wSwݎ�7��z��y�r�G�b3�YZRUiJ�=/��~���}�2xɫ���
�\
��/X�A��l���D��t�T.�R����*��Z�Rk%���;yR�4}��L��Dd�J+���27�%�_h��*/�5�߱�[
J���MQ���3t���69��y�Yf��ܐ6��b�9
�Kc�����dr*�G�=�1ཌ�, &P�˿��úI���85m�٪�#��KcE��	����������V�33b�Q[j�:Z�E�+����[�^�[���y�ݽى�zNn��wܨςE�Ɵ-}8���_�W�|#�#s���uE��w_�zwJ�V9����}!�l58A�b�aTř5�DQ{��&*ʞ�YM^��k���F�!q~�����*�Ш�4��f�V����>������g-����xR�gEx� ڎON#��Př��̣�[����`S�p��S�����KJ&c�l���kG��Fo���"��v�f�:a�.�y}+���O筆m��w��5;��f㥃݈�U`���=ϣ��ǟ�������ˌܞн����d��tqT�6���6}�/�CVk	���
�+Ț�Z�FCc�@���wv����r=z���7�"G'��Qח�9��:=�U�g�9��5���,:�ޚ�8��sI��Y>R�%�eXا6��+;0�s+M�wL���P[�O�N�@��;p�C�R�ֹ��#M�JX-h�s �ߎ@r� �F����%vP)���Y�n+kQ3C2�������*[���"��+�m�P��3x�l�u�Yk����}&��;L�����j����/)�n��c衯��U��K��^�R�
�4�E.�e�,0dxck����n+ů�n�ϡ����Ω�w*,�����,�H,��͹ʽ�۱<�&�\ތ���z�%�iK�����ߪ�ڊ�0x.Ղ�k�;���{���7�-��}�)oFi&l��]w#���k�9��T�}��
a*��mk��-�Ø6����x�����R�QUO�t�F�������әg�>u�A�ε��b.p-��ѽ)+�|�G��5��e�ļ�}�q[Է��W_8�����6�aV��V���*\�̶�h|�Cv
�غ��lmp�m�IRn��ap��"�sD-��<��dMrנ,��K͗r�9�^�_����=�g6	�o�^&���ћ��u�DF-�=����=�apɮ�c�����������EIJ�,���3`��pQ�F� p����WMmW�myugj��˾�N2�v��(fB�2k�j�z5s��
�T�B��l$���oי�~"�5N�����6�o2��;��r�\TS�E����W��Ry~�n����Zp>���'3&ֺK���-F�1�q4k]6�ԚЭ����9����3���~�]j�.ܡ˺�΁ 㥺�����Sk��^�!s�� ߸hlSv��Q��+��[ɟ���%Դ�+�3�]�߾�%�=�u�t�x�{������{!��Ѓ�ܨf����c��I:��E�,�ճ�P�١gG	F����B���h�j�o/�w�	*��������[&�y��9�ok��tX/Q��E��M7y�������Dc�0f5�ṋ��eg�įg,���E\�־�
<�}�US�9~�U��hjtX�3X1^,���^��{;8IԚv���SÚ�Ν�+�_���.�����Հ\��c_����:r������%��fM�U㷝Qb��9ǅ�o��;v��[�R^�W1�"��[#\���"R\q��O7Y�t�Op��Z�l����/ޱ�����
�D
ތ�(�$V�v�ͼb�>Xl��7���S��ښ'�N�"�q���n�������������kԶ�b���g�7�P�zm��I\X��Y�H:ޱ�I���&T#�D�O� w�
�N�O�Gx���I�-Ê�;����,���f��Ԃ��J�2`[[�ۆS���D��~�|>�=��Ļ���sZqIY}Z(���O[]=�c��r�}miR�ŸWIM�"�G����H�o���}��P~�����m���.��ࣚ@�3�3��5�/���u�:�XwrԒ/4�K�����l����!�o!�'XE��*з��� d���9���<��q��[������3tZ	]�v���f#��7���}+`��4�99#N��Ǻ����T����8��:��@��l��Vۆ`�&C,:��\zs�P�"Ejz�omtWd��d�w�����Kq��vO��g��	M5X���K�s˛8��T��F���(��ng���E��Q��G5��m��ymy��SR�۷hc�MXi@���D��pV�?P�g�zg�,�v��_ی�z�Gz�v�nOWo^��[�}�Oa�F���Xri����6�w�w�!8\���*�t�U=iiݣN^�YN ��-=ʥ�k{t���͑��]m�y�?x7W�D�ҵR�h>񠋵��F��w"�������M�I�cɎ���5��j9u���y}�Z�rG;�R�<}�Ҵ#��={���;�Ī>������yo�*���vm��r�t��u!]��O��yj�@s��D�v�ڼcK-��S��d���I��3�YZRV�%J��:�6������ʠ����+O�i����<���Y�ȇ]�M�� �5Q�FT�X��hW�Eׂ:�����H��'ϔ��M3�7q�X�EoR�ّ=Vg4��Uy�����;�,ɐ8�L}�u��O��*��q[3�,�l���>?g_h� &x�R�\�Vn�o�1m�5:sF㙻�ۼ��Y�M���za��vMz�h��a��ԓB��>F`�kI.A�J�r"���:z�t_1ZDr���&����^E,�'w|m�mZ�,��:���޳��C��;̍����y�֯ϯ�Ѽ��(������[q�Zjr����οjQ����P+��43^���`e�}Aw�~i���k�ϡ}��Y�/n��8n�2�:�Uǥ�G�Z�V��Y���R���Ս�:©Z.���N׎@�ᦒ��1HF��uF�^��}��}>�G0�mT�bƋV�y�Gs�]� �6I�]�ޘ��Xd�b'H,�S*J�+��o��kx�su������9Etx��/�3�Ǝg!}�0�������������ϧ�1o�}�[ʃ.�������L��k������uQR+#�eE]�G�b��;����Q�x�>���x���~��K��Y�5�K��:� ���&�v�rog��sI�K�K�]*��`��|�yܻqW�H9��z9�w���%̚��Jֆ�6��Dn�NB�vvn�{Y�����x�H7j��&��%q	�:&���1���Vs������� ��^=y"��*�B:�(�uܭ����s7jn�u���%�b�%(�IJ��ώ���n��*�<����z�I�૪��ٴkB5�w�6�hs��.�Z'ـN�ٻ��**t�[I����1;������||8�{ͽ	-�\u��q��YCƘ������x�{����+��Hrkj�!��2�VN��A\�[�@��[�El�����v�7E�ۘ�ܾ5u�0���j��fS;��6"�~8v;��.w���U	�N�f�^l�ݜ�K'J�Jt��[�S�]�Q�s��oT�Q�/�r;dG�[
kSV����)���ֆ�3Kun�oV�f�7a�$�@anX���B��=�t�N��?V�q=�����w!����֩��:�=��a�״��`�q��R϶2-#W�gW���[�?��)�{�EފSyS��i��a��@��U��;qM6)Rx��ط�������i���˺�n�;cdu��7y�I��	�33x�=ohj!֣Q�f�ә|�V��V<S�To��������X�6[ѧU͝��-���,�5�ϕ��]��}d�i���;�UY�d�{��a����]�:c[��.�Z���/��	4R9x@3�{}<�v��6s7��֗�ny���,��NsCX0�v����x���2tZ����]_=��m��Dv���|��1�0��ƷBT�hc��Z��]>��3(�QU��DA�������" ����6 ���=� \�ʄ+ C Ȅ2�0�� C(°2 C� ʰ�2,0�C0� C�2�C�2�� ��0�� C
°�0�*�ʰ2�2�2C*� 2�2����C"�0� C"0�C(�2�C(Ȅ0�2�
x�a�a�a�a�a�a�ĎFQ��A��E�A���E���a�a�a�a�a�a�a�fP}���ߠp�0�>� P@@�G  C
 C C( C" C C �A0ȀȀʀ���� ȀȀ� ��L�10�02 ˘d@`Pa	�Q �e`	��@!�@!�@!�@9��@	��&�Ti�P&&FfdFbe ��A�ei�M���L�LL�C ��$2�4��0	10�s�C�"Ly*�a�eXeV@�!�y�ʰ�2�2�2�2� C
�*������׸1�����AhX`D ���8��zm� �a���~��Ǘ�\rn��P��$�/��
e#Lu�*���������"���������|��$;��O�kv!܈���q��;ܐ������0�ǐ�?�b���QX� ��)@@� " �D �@% 
 ��I ��@Y 	@@@I@X@F@ �� !$@X@B �� $$@	$ 	  �� %HFP��`IVP a !FP �@�� 	@�@&&P&A<��0�������'��ZPE(
����~�[r��մ(�8��QU��!��Jw��]a=�J�0=l�c�jT؟�U��!�T����'�EU�"*�����?O�����E_?��y�!TW�?���`�_��x��?���xa�����xQX���j�mDUEsa2��0�!ՙ�R����PB|��a�ETV���b"�+�
T(o�
�Bf���fHY;d:���� b�`�ʨ���R����czJPP���=l�������"���G����@Vc��tj���	Cz�(+$�k<M�S@Ɵ�0
 ��d��Hso��	�B�B��I$�B��%�T��R�T
Q��(T@R�PT*J���IQI!
���D���uҍ�B��j
��45@J-�J��
�Q��I�$kC&�*�� RD%�Z��THF�*�6���������B)� �b�A
���hb�ZҨ���*�Tlj%R(J�j��T��Im�!RU%JH���UP���QPR*�R���   ;���T�k���T�u¦7vݻ�������u�ݴ:j���w]�e�Of�
�E��=��M[��+�s��wiz�齄�.�ے��˻T�u��	T�����+�   ��:
$(P�B��"E������=oxP�B�(P�����U�V��V���v�
k��j빬��݂���T��sv�n�m��j�wj���&�[e�]NU��M6�*J")$���   ��h�����[��Wm�Y����wu�ՙ�1��Y�*֒˵5*�e[J�Ym˩S��j�t�h�h��d���cf�d&���;��N�n��N�R$@��:�I!�|   k�45[eK����n��\�ҵim-�dl�n�I��V��ۮ٫Dխj)k(�Q��7�WKF�UXզ�R�M���QP�)�����E
EI�   ^֊kU��4�Z�^���lљl�ZQ2f����be�wj��-��6�ai�Qn�+�bh��j�VL�f��M�)@��f�   0�T"�2���XKG���h>�q5H�����z�������ZR0��a��	l��WUjڂ�jj����XM�B��U|  ����U}ڜ���U�֕�i��L��A�NrXt� ��4waM��  1��=  ����z���"�"H�*�%T> ��@(H�����O/=N�S:��+�@3��@: 7(�SCN��l� 4
f�=: h;���Aր<uYGN��a�W�4�J���(��� g� |�ӎ����â�t�7@ :}k� )�� 9�x�� +����:Q��wJ�u��d� 3��H(T��Y�">   �@��� o�N��+L��V�)�v��(����B�;��zz �:���
�L4����� �h��@4@��a%%* @M�FUT46�  �~%)P  ��%U  BR"l��  �?�����|��߷���F2��,M�\�s�d}�;���v)��������4O��TS�������_�E`PUE?~���/O�9���
�U�t�U)X�&��Ջ�KSٲi�{����6Ηs��S�AܬƩ�9�X�{t&2���[���E{����&�dQ�6ΓVw�`T"��(��f�٘�%Լ�%\{R�m�_�u�x�v�r<������E׊��M 5�2�a�(<9�u*�2�R?>�mjF,���QY��e��ܕ�κW�	i`]5�����+8u�4�Yu7B�h֜gB�O-P�%Ӥ�R�[X�\�ŵza�{�jV��@V�-4v�GLYm��!yH�1�
����)G2d/7]kߚ��
�1�e�)ؕ��d{�V<N]�KT@�{��T�=�a��ѽ�Q��U�*>L�VX��Q�n҉�{�$U���0���kc���f�XFTk�m�[�dk�gwr��G�%�ϕ�xq�UҋA�N�ҵp��Z���ծn�GC(g�U�ݟX����T���

��m=���8V֪XƄR9r!�X?h�o�1R܃w$�·�=�/ܣ7^ǹoŦPP��t�Մ��*�m�!!E��,%A^�Z)�%C!gL��E맷Iiliˡ�-ed�3XI :�YY/a�u��p�A�X�kh;��-��8sB)6�$M)@и�m��v0�U�8��zD��}}T��[��@��s� /*A�\�9U�B�]F�٠u����T��/��&\-�����thw� �_Դ��:����j�d��/f�L�ڛ�p�9�Ql�`Ѱ�b�X�{�)��^�7L,.J��&5��f�:kOkl�֠�Į�c�%e9F���cT�a@��V �w�4H�B/v�۶��g�(ǰӿ�<��:J��s�u�/���:O�n�x�c�k
{7S$dY� ��R���t��Oa��]��T`d��y2���\���i{����t.h�d����G����6��h�Yr���)�.�b��z�ٮ��35ZeJJ+Xʍ1H*����0�y�`y"�v��q�d�(�EL�9��ګ�e�p�b��Y�CV����5ԫ�$6����#��0��G"H^fc;[�c�w`ċ1JtE��>T�L&i�Y�
_]�]�M%++v�b�3jj!�W�dR%6�ܐm�fѕ��ܱ��-z�!�Z�dKV�;H�wbf�����e�)6I`�뭫�d��2'��S�U�T-��[ h�Va�
�>�1�)�Wt�/n�����z�Jȶ�oD`�D�a8�]ɮ�Z]l/Q��t�>rk�P^P@,�iK ��6��w��鹒��ǉm'[g��4�v�mMH��
[MG�Jdi91�vJ�-嶲� f�sqi�t[�uux-K���a�3mG1��T$/֚�Z�����*7n���bn�Z������l�h�QȰbX���T˧(�Z`��SaQ�b0�&&7jV�a�V��o0!��JZJ\"���N:YVrm=��iM� �W
�(e��b-�@=�Wsc����n&�ׇ�,�|Խ���V��ITYXj�&�b�j��ʋ��oi9�j�`�>z�Se��T�5�o]�ʺW�����5T�(fs�\����-,2����	f%i勬���(<-�B[��-X��oF�`65Uܛ��kf�ƶhA4�Z������U����3��ۃ!�oo+EC�0J�\]�^˔s���J����X˼jbR�d�N�m	t+h�F���-�V]�� ��gL�s�#��P���iq��Q{N�w�4w�)렢S�I|�oe��(�j��.�8�M�S2,�mMSkT����(jI�sZz�
60��D��+6Q	]¤ߌOj�Yʱ'�l櫊Tb�6��e�5.Y�h�T�cٛ+2m�"Z5�
�n�͡X �e\�w��"f
N�VZ@��[.��F��aI ���U�׫M!����PԈak���=T�dx�HO�X�,/���՜���CF��a���2�`b�=��6k�r�ڭ-��X �5��J�0�ǹ���Qx�J�N��T�uଶ�w�aͷV���i��x�уPkh	y�.�yY�9#R���P�pH�^ж%K�I�mTR8] ۙsl�n��`��i�/SU�&�)l��xu�*X��Ce�4&]�v�YD��7KZ��4�V�l\��u��D�t�wd`ō�� ���k)��WQR���ZV��ِEIRh|dWi��ǘ��!P�k$�Reʙ-�p�wW�)�*!�e�L�!P+�T����]'@͠�l�:�LD"���,ډ�Q6I�[����$��e��2��f%���^Rwp��e��Z�7 b���nf֩y"���:66�}.��uf�HS��Y_-��.
cZ���ˤ�⅝6�l��r^8tKGVi�΄^����j��"���ؖ���5a���n�h�n&%j�opjsn��e4�a	��y2m��A�<�hm��і�4�2��ĕ+*ը "Q�*�&�c�+��[�aH��Lm�Z�h3j��Gnd�ĭΛRV4SER����R�d�[�"�����v;up��nL���{�=�}��IP�%��J˴3�v�H��Z`�-�V�KuwDDS�A�a+v����Sx���wCI`�EہS��(�N��[���hLUoFPIMd�:��n�Y%���6APU�M裤T[��(ص%��I����U�y��ޗJiY0�4�iI#�ec4ΰ�Q�{5}����ʳ�&T�dv���%
�NX�m�U$��0�4���V۠E�)^����{,��V���VA��d������d+7Y�G�](�wiX�3�����1=���î�-�." !�S�w]�;,��jآ�B��D�f�	�X"�9��n�.��.Ģi�U�o�R
ܽ���c�]i%�������pi���K[B��8ν������TE;拼��1j�J�fG�Z*���wT��͕�^��i3	kzZ�T�1V�zʻ��Z[�Ɲ$Mm֑wAcNҽUjf���
����.���V�wQ���j�vV@�b���A�A:,Rg2=��"w!,F��\&��Q���'Yqi.SlbY���������T��	�i�w$𜎃{a+ǪR[�K�SJ����0�y@A!Zܽ�`�1p
f�fv4�u+[Uz�
��÷�]�(e��R�}�M[ Ŷ�X�a�R�QF��y)҅�4B,hB�����y��9Ka�%(a��7�&������Tz�4�]D��9��v���:�X� bv�2�b�A����V�H��w,Ƌw����8�5^��2+	Sgon�m�4ѭ��	�ssG5 ̙�Sdh	A��;�6�J�k5�^�yZ�(v�z�3������۳-PJ�����VKٙ�`Ϯ� ĠVH��|�O���l\ٖ(iWM!)�:� WN��f�n6B�w��wۙ�0��Y�Fa���o*h2d�������y��V5*�v�2�lT�	R��Lm�v�5t��W�h��F-��\���еR�h����-��՚ݥRdX5(�\�Y���)��In�U�#R����H �̈=F���s7u��6�� ��G3�M1��47����Y�������c����ɬ��h����Gq�F[5)hR9�w��U�����hK���K!���0F���Tdhmf"w�# E�)Dpc[�{up��v�:,H��RՁ���:(䷚�Dy{>t&9�$�������
AVV^��u�d���B�����4�j�4�j$�*T�X�֮�����O+	�d�	<��r�gv���v����k[�z/��ɍ��M�BV�J�GN���L7��V���b��y�o&�� �@��E0�<��$X̋1�b���҂�7��;"U-��HнKbf/Kʱ�[0υٲ���@�7	�f����� qC�7Y�2�Ű͢ڼo��ck[�.�S�E�w���5v���T�k�V�xUrU�y���$L�FŃ.�%j$�5b�1yxq%��w�Z}��@'.��`*Ycueԭ�b޷B�R�j�����U3P`��^bkiǄ){���>I޺�͔BkQ�٪�F�hU��sck
W/m��WJ�m�ډM�6Ťӱ�1���`�ɇ(A��}{yQ")`�!m��%+��lÐY+p���=����r�$�y�=����Ɔl��;����j�z�4�F��î޴���a*�B[�5\4)ۅ�imH��YNP�(�T�Yj�໼���0M* :($>�\2M7CDB�.O�wQ�Z7^� `r2��q=��^�w,}�!7On��]�j�rjqԧsYwA閥dݼҥ�yb�e-��p���Ե�e��5S�/3
��i@�)a�jb:��A��K�aݧW��컳�Yǂջ	(�<z��NY��[leꄤ��	#&Lfm�6��% ��J����J�٣Da�vޭ��7N�áT|�C[�L���H���s+)��VRS�O���n�{���ŀ�Y�n�)挀%M���а�h��Jf�E��;t�;�j��D3�r��fc�^S�b&Kn�o"�z�b�4�%�z̽�q�j�u���ՠU�i��E��m8�ݷ�̻&�t�B�V�tc��jg��� XDa6�]��]�E���3���S�¦�v.#�Tյ��R5!u�%["���{�EM�m�ۤL�&���6VL�i@�G��uִ�-��v�Ĉ�%b�s)�/!ђ<8n�9nU(���ܩLݍ�X�Bь�v5C[1h�]9K7k*`�˺P:o"5��qX�զ.$�����X�����@M�`t��TZْ��VH��[����*m(5�zq�*<1	�a3z��F�q��c�e�c1e&�h�CiåR����t���VE�X����5Q�C,Fe��譨�Cx�|�9WGb�^;!��k'd��n�6ԍ��p6T��VM'�-��ݬ*�a�ţh�m!�H�3c��e�:�d.Q�N�nct��бY��eދj��!xudi�)�j�H�eԱV�bKJvk)�΀ӈ ^e���T�r�7P����L���+hՈ�5`�t1P(������M@S�
3UGz+,+�T�����Q-5�T:�MWwS�*�VTU( Ѕ
��(Kbd�Ե�i
���6�k�1��(uk"W�E�ܸ�?hH4�V��-k�V,���ֳ[�؁��Rƥya"Nm%�T����f
]XZ[0�7.��P�'��T�U�oY���Ӗ	0�U\nӥ���M��m���r��v@�N浕��Z��&�n��{��J��!�؂�c@�0�J�2��ޙ!��QT�ͬw/�i���Uk���B�5K��jY���-C�Mջ�ʺR��C쫬,ÐTW����R�;��qPC.73we=���&�,��=���l���B�0�2 p�_�KR�&�_�R������N��i]7�o��F�!��7�q�cw���bp$td�w�������JH��W5�
#v-����Ӷ�F�U&�ܫ�q1���h
�N����%f	� dPB�(F�dTݬ����Ma��bTǟ+W�&�^ā;4N?�mb��Ʈkz	�m�AՊ�U��	��E5Zh���z�,�]�u@����L�5x����=V��{R���A�X�K���٢��XF��fQ(�(f��j�rIj��o���Yk-�$)P��n�Ur�vݲ�wY�i�ӎ��j;hj��kZL��22�E(�vs��У6��e*(5F���08%<�������4<Z/cM��M��A���In�ٶ��jЏ%Jڻř�͠��sqe�(Mk� �:71!N[���3�vN�ZK�&3P�Sf��dƫjۅ��-�'Fb�]+X����F��ѫ����2�[WN�Ծ�F�d".��y�%]�AjL�)��p�T��yTѧ��[�����q���m�Ue�`�&�=�ة"wt�jk%Յ���CnW�V��n�j��g,nLf��L��<�[�`i�kb5�݄pL�!�(Z�*)I���,�Lּ���f�P�ї�g�DB��e;a��7B� \yFaˌ:���#���b��p��-�jܔ���e��3oa�S�B�9�� /c �Q�
��^ذ��&��"]�3tm=����XTѺ������sj���eɱ��fظ����j:ުÍ������6�\�5|m}���V��-�+Y���*ҹy�R����׻�Vh�u�&Kji iYv�cf��m	���Xa��fmeHɮ�$?eJB����K�%C�l��hgR�6�^<J�/B5�Z^�	S���(�u���!�9H]L9I�ER�w\kaV�u�P��@KE0����)�1��]�x���h$R��ɦ���޴U��Elh֍�f"�!)W��Y{��S/%���`��X��I�ni/Hh�A#t*�-ɩ^���VF/W��Bܽ�e�r��pm��2rE0`;A۳�����
������fQ��q�_+�pjV'�aS�D�,�.��)CI�yX�P��<T�-L��i���h��T�h�U)F��6��7��Ќ�ܶ
��f�m�n�9a�Y�11�+�l*Vj�q���0�����4-���z�5����ũ���J�C���������RJ]�h:z75���-�Qe)h1�Xn����ȴ���ll),!f����5��,Z�2<����� ��F<mF#��p���0:�۩�0^'�t�@�d"�iN�&ZT;\�?���u�f��{�whv�5r�����S]��U���RF�v���b�Y6��(7�1u�e�rv䋀�-Q
}p�l�J��h��^��+&����&�۠ŭU��)4���z7s�:�\*wc���9M���3�y��I;x|]^`�;��LB�:⸫�յ�F,EV\t-=�2��wB�yS��ZQp�e��ee_S���Z�t�vy��rɈ��5^"�<�C\@���w+U�� ��-٠Z�v��N��f��69�TVK�@e^�cS���-���b>���J���F6�Jۖ��I�W\���	���G���JL��o��򜙆�s��a�p�t�G���;�<����h��e�e�lE�u����m^%\��[hcB�\�u�Z�֜����[f�4�Ҭh�X��u�;yS�g���]��Aݙ���y���:�u'K)B$�v�Q�ӕ�����+�����Z�O��a�����b��\������s��Q�v�3b�b��r�\��ă�&gf6rMߋ �%8�����N��m��g����B�q�.����J@a}���ٍ�Gy��FF0�
<o�`/��=�;2���38��bQ�ղ��i���dʈ;�֌Ի��I����\�����3�\���t���r�@���r���`'t�m�>W�N�m��Kw�{��g��jJ���>�iC3x]Xw�'tz��Iz��� B.vW��/+�l����$uϏtR��%S�Q�ZC��z�o�%K93��b��+�$�f��J�ܴ��>�\�+vu
&᧳n�r���x�vp��ܪ(]����nt�#�R��e��$E�h�w���<+�V����՛�
����$+z(i�]g�T����d�Dp�<IVڻ�kw~5wC/��(��K}��޺��Ĺ��T��}G����o,�Xu6�������j�}hwc�����RI*�AԷ�����&��,�ԗTk������=�hxW�wT�Y��	�Yxn�=�I�w�O�3
n:���R�C m�f�v�Η��(�K:3�R��g��]�:�̭�h��F�vh�]�űWٔ/w�i/��o�� ����Vq�[C]�����
����9�M<�{#Ԥt9�d�C��h�̾�z3{�����n����v��8���V:
c��{Y�)����V���<:���Y��r0��r�W\޾�cl�
۽��F^����g\��E5u�6(-R4�+E���D� ��KB�"�s��\�Kr�f�1Ĳ%�0g+d�hNa�j��J�-X�w�.hLɗ6k��0��~���"��z�FiV��o.*��Y�X�g+�;��P}�uJ�����IY��.�\��nk���M��*���nR8�����u9gv2�8h�ҷ��k�Y�Du�,`�\����QeΌ����ַI�����/uc�j�WA$���PҮ�_R!���A�M�4���|�KnR���o��Vk��+��ۢ��(u�CZy��)�:Շ�uD���e>ӝ���dY�w7�3;eM�zB�5sŘ�\�gL��2�<�Ǵ�XJ+��r�o�呇�I�c���4����	l쏕ɹ��\��WS������R8�k�	�ԟb׊�Y��˥B����x�1YjAM�K�Mm��aDV�Yu��	8m<�u�t8Ζ^�D������5{���;���F9.�q�kI�ui��}K?�"�y�}\�r��o/}Q�O����cS����\Y���G\�>V��;�,�ǖ�	f��MkL�մQG �5z"�{vZ�բ��[J� �и����}HoIϤ���O�#��ìՃ�[�}�
�Ck.$:c·� ��*���vf�WN��=׻���5�imҺ�eҽ&@0բ^�HV�G�����a��So4��YY{�²�RJʚ%��>Xy��A ���r:�E�m�i�6p2��q�j��jS;�h�����K�soq;���X銃z�w2���� �W�`:!]��֎�r[H��/���au< �A�&`R�[�ve���o�X��*�Ev�َj`�
�K�;]�J��L���2���3(�O7�n}��ty�Cv�B9O�WT�x��;eF���*�%e��p��8+R���I��SN�hPb��R�5�Q�Ω+�^���L�z!���ٲ�<�uD���x�v�M6�B-St���q��%�٭ӛ�V�I�H�}{os9�|�mI�X`��f7���'X�RZ�,c��Q��\���R�rhJe���֋�%�Yj��è��8y�'#�7r9����
�Վ��7x[����ֱw`\�}�1�*ﱼV�_G$�5��J�3wb��e�!���<�7<�yK5�ԙ[4B7��1��R��o;�ä���;��4�-�f�4��l�XqU���ض���|,�y|-E7�l�7S���7��ob�۱�h��9���b�2�Q��:JYN���T�k�[���G���ivVҴ�V3N�:uC�uu�]���Ҏb����:�.��`�ގ�hM�F�X���bڥԥu2Nd��XΡ�qWC��d��}�mc;}yi��ڽ۱*���Xa{���𷶽eyn�4z�!�e�C%��x�䳍���ǝ�לV,������wYٶ�IM����ҵ-T�h9��������t�
;��G�@0f�Y�ݠb��;lEQ�㱄E�E��<4ͺ�/u�j�/�jj��U�L�AK�t���Ʊ��,���!e�6��}��e7���Ҿ�p�ϛǭ��|fM� �(�iĈ|��_.�N����3i�]w����P��l!��3�F��՜
��+���}�z��]Ա�8%�kN�Y���i+�ڝS�v�J�+�T,8C� � ��oxr[9���*�v��mΡl�Ur�J�㛘4����f��*�+hSϱÔy��q�/_70:�AV�)f�,
���e�)�s`�
�wa�t��#"��W�ц_�5w���.rt��[����e�]���6��k��+�;y���(��}��tfP��"C����`c���%��"�R�x�D̓F�B�Пm��n�����'�쨼�]�ֶ#�E�i���w������mt��Tީ��zx��t��8��ɱ@)E���.��C����=O8ށ{�+K�S���x����zV�]2
LM���^�W@<�3ݎ-�4e�L>ۮ�1k�S_<��yL�l5�|1f�}�f�eD��Րb��F������6A�������]���-ɻ� k�^�me�k@ѐ�$?
{F^�K]o���	k���R����"�������.p��-���6���1`/�Pdv� �������8Zĭh���)ܶNf�i8nq ��v��i4��J�:�i��t㻈 ��S���rQ�� @WKY�=�_�x�H��$$+-F��՛S�,+��V�$Ñm��wBl���Ƃ��mWIa=��ԛ�)�2���ٷ�Nf:Q@�X�8��&f��Ua��l ���52M�n��d[t��w%�O�V��꒍JA槩���z^����O��׮��e�n�����Lׄ-�k3��,s����4�^��}jv����e)+kX,#*��;ǥ)�3I�(1�2���z�Iâbmq���
�U��7.�:�V'd�jΗb��!�����Bc<�O�T����,0�bH%>�����՟Z՗��2�Xl��c*�ͩ[+R�+���oK�RQ��-�V7���2 f��Um���paӒ���B�^�d.�S�w�]��)[�u���ep��Q�:�rx��*��R���.N���C�{��ڶ/x�nL�m/ vT7��ӆ��쾇1w.��Ʈ�j��7��ﱫ�d�{q�[�����guD���
sN+��>�MB����l��V9���6U��f�)�'�M��c�]q��e8�[�Vk��H�*�P[{�nDȚNM跄?	G���wR�%H��G�8>�@�3E���6��c�ז:�AN�u4�F���TX�fi��K�|﫸ҷ`l���*���7hd�U����x�DJ�n�VJ�1@mF�u�vͷ�}r�hd<d4yu���X'uqt�uV�Ku�+`ْ���鲯���p����7�������(�f�����[���e����ޥ|�fhBֽa�fW.���8ޮ����'�b���;��#������{��wP���hk��3C�\��SuԬ��v	� Σ�4��Cf�b�}%��
@8o��[V�#d �n�إ���E�[�ˋ~*�Ժ6�=�B�b<�{��$ڰ�������Wc�
V��g(G²�ƨ���9�#��.ݖ��\���U)���۹�n�V%�lc:)�9��Z���j�[�����R�qǕzM���k�ܶ�`���"g�����6X~�d�	P�U�7�2����Bf��&�$���q������pj�e��o�����6uM�6���;�uX�rk�Y8����4�u�l��F����@����gK����Vm
��]ސ���U��GX�B�%�+z��5m�A+�V�	p�oF�z��r��'[ݙ ���ͷB8\t���N�V���8:+Y��J�L�)%��n���A��{�,�:bin⹩�B�et��`Y��3M�ٝ�e��7��Y��_rC�f�6��.��q,�Kj*��6��v�;��TN�
��R$���[Y���n-������_1�+���.M-論D�2�E�d�Q�kx�7�3�6�U#�ٸ�|S�d`^�8`���}[��el폯/j[��5�s��q���+w���2�N�D�$2�&d�/ga�)�5\�x��Q3�	 rE�K��ڏ�5�%��6� ���u�|�=j�:|��3m�Nӻ�����t8�E��V�	`-��ۍ��5���
H������t����c3�a�@4�"��L��v�A��avdWO��g@�mM�@]\��S�z�з)Kt�j���@VWzyfm��62���[BeJ�jz�f7�TfdXj��cN�Z㗛z�iV� �G���)wL���]�9\��3s� ]�KV�V"���Aк �J�κ�;��p��yY�o�iE��Z���JV�.F���h�;]w\���D�
���v[aY����讂w���ݙ�6M�w�ɔqb��/�W3��Q ��YnQsM��Ӷئ�i�u��+-������3+����&���{9�y��w����N���5Ƣ�Ȳ��t��(���l��5
{Y���gC�b��|�m@]��V�Gf��,Ǘd�:���\g��rFαcy.�q�W۴o8:Z�qJ�2�o��{��K�Y!������4���Q:���G�Xs�y�wy㥴���ut���0t��Е)5w�R�#4ե�r�|/X�T�yv�t�J�qI�3"[# �Z����>݂;�c��h����ʖ�4d��N��E�4^���
�:��f��A��j�$��v7�r�9���ed��_YK;nwT�Z�g&T��R�n������,g�k��#���՚g t�{�/(���7�ճ�ho�R��(#æ|�,kc����u1W�ښ��]����Gjܧ]�f��iPG��CǪ�՝�ԮY`Q��w}X����_~���o��zҚ�y���	f�!�u���^C#9�*]\i��ge�v��_p�m�:<rH��;�Y����:[Ki�R�[��=|�^���7�];������-mYx��u���q�m����4�4��tG5����Nr�ky�bJx���%E)l\�������풰�f�]ge%X�E]�cR��p�fu�-q�U�v+ŉ*�]Fi�]'�)��5+4d�/+��Z-��;���X�����O0�������B�NnU��hm�aHgw��vó���F�\Y�fK$�����Ib%ʚ�<����O���j�e�iE5WY��Y2�Q��FU�^�����6&%���,��[}��U���7�tCz���|/

��9i~��@E��jT<�w���-D2�]^��q�39�)��������0���2��"U���ʫ.�.�ĳ�s���敫W��s]|���Эb,ɃE�@)��־{�����u�+{���.*?#�І�t9z=�l��]�	E퓖��Ϲ��ٺ�u
R1V�Lƭ�d��2e�*�Uai���t��y���>bc�}�f�����V�<��U�cqn'���n��V.o�NA}�#9�9�he:�Hl�a��Xi��;뭾r�L� ���Pi��= WnfG]yp�:�u2jtٷ���J��]ό���/).S����'V�_!TRS��K��5��d��3��
׽G0��xz�e��i�u�t�1�fΆ:2�|��bڅ��9o�A�v��U���
����g,(*�㨻;!��r�_F	�7DΧ��vr�`�-Tݓ����tGWQ�3���u��:�/�D�����jہ0J�J�����6pq|�`F��\��}��4%��ˮ�t
V+c�4�>����&��p����r=z���G7F�oV^��͇��=E]%�JQvh��j-ܦ�R��[��%�'|���5�o��k}ZW( ��_n��m
��b�{��
&�����}���P�����Bl�m�k�s�]Y3@5|��S���Z�5/2�kPQu�Yι�׫�l��\\)gV���L���ee,�)DG����!O�zM�@�]��Ԃ�t�J���L;��qr����xm��`dL	M�W�9���� ��07t	Fr�ѓ�q�����ec�h�n	<grpݪ/�lfcR�:�	�Owr���*r�*N��W�U}��)��@DW�}�Ͼ[�n���ߜ�����ܨL���`Pu��o];* L��w.���%�x���%�O]X�A+Vo�V_^�}�idT�Q��%ʻ-�oo�e���ޚ��U��Iq��΁�öQ4.���*[������
%�]vw�3Vj���`�P���˥0Ӯ��W]�lTBK}��j�◖�um�bڊw;:t��(�[�!;�%Z��5,�Z��*r^fk�J#uA@�����F��_1H7}�2��|�vF��G[��u2KEҳ��nhf�5�3�Z�%�"B�*��
�C�Rv<���U{�)*�Ѓ�a�����պo(l�]堕�br��MX�V�KԦ�����%e*\O|VӠE�c�լ�*�,P�Iզ�z(lՋ�pu������W�`�/!	5]�*Ἳ�.��z��t���Z���V,.�sV4��م���ci�@,�p�K1#��ʽ�]tr� M�rAmf(���f��jS��+�3�,
���fS `��h��wj�+U�YA��#V��Nb�]��Z�YKRh�HZ�7l3z�4�v&,Ι�p1�EG
u`hi�=�,{8����Vճw�H�K��:7|���u)��c"�Ί��g/�<�;���Q�\��l��t�E�ݝ��BU��Auյ�.2>�1բxQ ����#V�����m�4f�YՃ済�)��yg� ��)	����RMo!�:�&��y,Xx� j�<�v3r��:�(�'p�+�a_a�К�����;\��e��˱z��[����6s �~k�m@B�ST��+��vDi=p�x�����l�Kv�^S*ⱝ�ɒ�p�èiT��X���˘���U��@5���䧳Ht�T�9�b ��m9��P闃��Χ8�� �i�z)(U*4[Bܻv�f*&���D��K��`J���y�����QPa]���k!u������K �H���A��J
��LD(^���+��
��Zu�r`�8j4oZ����G9\�u����8�[���̐B�V�C;�菒�KMY�w/M���˾/���.*zvW*WR���%�HY
���u�N�6�8]jfY��ϛaק�ջ}�����Z�ʔ*vmmH�����^8��R��b�v$]yh�C��^�����wxzq�D�.�� 맏�DN'9�ړ�=	�αg/�v�ׯ(Y��p�M�;��F�鷄ƀ�\̉1�EX��ij쬲�N�TBXRÛc碲�KkH�YDI6�A,��&W[W5�}nZCC9:;�C봟e���� Kw���]�uN9Ob��e�n���*Y���n?�r��uv-�4�t�m��R�b��}�a:m�D��,1fj�t#��'ۨ��g�M@�}ۙ�`�y+�4k�]"ܽ6��k���jR w 03�R��ge�y��Emu���F��F�8�qt�J��C�^�9t�@�Q�0:�N�Sct4� ��Al_
�ɋ��4]`�j��\n����4H�mQ�py�5������֎�~�J�
�������5��C�/a�9�]���sZ�ʔ��C%eTgw�Ӆ�Q(�wiI/i���w`>��s�N�>�S��D�#C�i���MA�m�c����S̓ZF���ж�h�׮�ڽ�Ɂ��p�W7op^��G�0���[�+{o+�wC���@�c-�I��cT��ub��r�����5��B�[a���Dv���{F�a�6�p��V*�\�Cz������$�UL�ܭ �_�7�a��u��HP����]O�L��m�H!Wκ��K�/2nQeͭ�`�nEr�n�-g�_r��9ێ�=�� �k��)�(֖�I]Gz�i*�%��H�p�_�Y�c�ԟ;��.���]���x�1B�V�P����+x�����Q��4.r6*�C���tO�ǔ�j*Ψ��W�^�*h��[�h�r��Ri]wr
��ɭ�[hZp�*l�3U���X����N�5R�'�S!�-��N��I<��P��v+��|$|:r� �Z��ZӮ�"�L�N�.�}O���x�]S]��CLcӚQ5�F9b�Ҕ�d��K�����{��oG�3��(]�[�iȫu�F��r��[ܠj�̴��wUi��.�pQ���7�]r'w@�-|��K�<4�f��f����`L�Qn���H(uY��]*��M�Gw':��c����Eu���"�V*FȴkrKP�;#9^Pj\�v*�`|[�yP�!5w�.�N�|%�R���C4-!��a��nݟ���k\�1���]�У�-�\�;U��Y��^1�(Y���r���gC\�C1D��tO$WV����Ų,F��Fo1puD�7n��9�`w�2�k>w�t����ĩ�bVu7��u�b�ŻW���QZ�̼7̋"���u��}ͤ�)֝�mJ�t�� (`u��'��}K��� 8knA��fũ�0�*I���U����c�Q�F�a��@�cʹ�WUJ���7}#ԕ�#�Vs�w�ڢ��pV]�ߣ�̪U���#i�w�pOͱ��\u��@��G��Ǆ�U���\g���ݓᕼ�(�VЩ{z�[��T����/qѸ��݌Ώ��lX�He��tN(���!�h5�R'[ov�`Y�Q���ޚHV�b�<E)i�1m��v`�̒ܮ�qE��4��1J�f��9��T�0�`�̘+���
�k2���p�t7�
�	��)�z� �wZ�=��ۉ�*�=&tA�0^v�q��S�1*��Q�K�>LN������%¹��c�F�� �Y��D���u�J�}����A��$�y��o⎤;qHMg>�a�
ٲ�wN1l�uoT��nގϷ[o5��i���lƅ20���|(!�m�a��2�:;H�RƎv���Թ��D� �8�wC�𖒻�a���L�D�{�#�����A��7iݡ�ǃW���z1n}e�j��b�wyd�x�_,��C��z�S[quf�m޵�{}VݻT9���<�wN�h"��#I����[��G}�.��]�ɋ'��t���E�f�\��˾��1YM�6(,�B�Tb���{e��WV��;W*U�;��J����ȃ{�}�EC�+
`�پ7q��+�L�P�֭|�S���<�b����s*:��G�v����R��"�QT������VJ\/x9v)�	�δS�&�\���g�+\�ѫ]�=���p|����!˩;�n�Vcr]�j"5&��.M����M��e$�]�y����6���G��\,��]Y���q�0��T�.�E]�j9�[����P �� w �Xz�WS� �E{d���٫t�ad��5,ێQ}>�:lPչJ�O�7��+�3Ks�e �2�.��oa��K��)L�ʹ�-I���f��ob���9oJQ�j[v���U�+��y��p�iW%iyw �B��>��mWK�A��VWra���i-���P�A`�*s ���c�y4A�s�۲���Q����40���b�*J�
JZ�Wd���8p��u�'bf�kC�np���R��own�)�wn�H����A��-@�B�Cmh����ܖV˒uY��y��|��jƉ�N+���m�4�o;ro'��2K����Wf���wJ �N'gL�K����P|�>��
X���
 XqҲd*�:[��ż:��rW�z�M��Y��{\ڴ�
�h�6R%6 [� �8Z8��L*�W[��\:�$�٘qS[�G!��Ҥ��N�a���X�B���R��1s�S�}{V�t")C�yN�P���o�X�+�a�>s��I.��4S<ki^�[��O��u.	L+��?tTwꗪ��2����I6���Ob[D��q@��P�l����ԥX�
V1cu2���X��n;Z!��`J�=��y�s-�<�[�CY��n�VL��S�.����wAܫFU���g;:	�i�q'����u�Ԝ�����g;.@m�ZT�'g6�2Ӯ��Z�6��;N�p��4ms���+v�6k�X
�(��D��Emܬ�4e⚔�.,ɢuЭ�5�P�ׂ����E��x���᢬��.�*n�ϊ��iH���%�E;�,��]\��t
�﵃��� k��r��Q�ʂ��վ	̥5��h��:��z0�݌6��T5�Ԩ_�e�h�B���v��X8=V$ʐ|�_?�Ny�n�I���x�t�0 ����X
{���zn�b�wp<uh���������(►����hX��0��vV�� �*�t�ӊ����T�ަ��b�gp�A����Y�������m#�N[5��t��z�s-�pX�X7>I*R��Xb�h2��|�t�;N*k�ZO+�\n.�lZ��W��	��Y3_�M=��e	%��
�����U��O�p�xX,kqӗ���n����WQ��e�����:�զ�b�\U)�+5��
6��l���6Q�l�SA�jޝݣt�\��p��<wx�Y:#��ړ2�<�'L����-fq��t1[yWo:�i�4-l㝑$Y��m�9�(]���["�T�M9��_n��	$�� �f�h�;��PͳL���B�vDU�tٱ+t&mL Q٩ �7G-M@EKU�c�N�4r"xr�7:�K5��x�'�0%�x��w/����b�3��r�%���cᵗ�]s�WȊY1����a�Mu**`�f���)���[�D�`�ZGcV5j?�q�)GM+�ZFa�rV��]nek���;0��sn�rC"�Rvdh�.�tU>�S�X�s7���.���`���� N��������9�	��R�\q�<���Ŗ+���&����Nǔ��/��4��VhLGκ�켜�U�b=�ھ��s�M��}:��A� U�H9M�t�������P����5��S�ō� �nP��=��rս�>���*ê���x ��s��3{B�����|��"�=�ydM���y���mT\�
Q[[��H�N�Rxj�kf�j�hQ:H���6m!�x>Nky�.��.���z��.��KI�e������n�ի�$�8��r�u/;'e]�0i��G��Y�)2j��ZpYܺ!�	�W�;፷5�Ƃ��=�V�S�Ф�k�%d4;%p��G�r�N�f
�U��m�+��9#��JҨ+f�6..u�]fL��V6ӗ�=�-L/C�3]]ZsT�ۿ�%D4�Ԯ`[�J���O'��[4J�y��nr{F�n'"6(9cw�*�fn����Z��{q+(D��CFt�OOV�� P�*E���K�e�%ݬ�2J��L0ѱS:�pj@c%�Tm���0�*u�zsx�)�(�ݢ�Jܾ��N�̶'{Wc�H���9s� m��ꏱ�l�kɲ��:�_ch�Λ��ŗ/��'o����u�������s�����u�9�~�D!��V�J�iI�%cx������ `�9rd]�A�v&Ppæ�sM�����HQ=2L����Q�a�R�v�h��)P�kin�+	5n�dY�+"ywd>� "������P�j�aį���t��T��P������:�����R@Z��=d�`��νè^$�=�ez4mC�1ڒ�(]r;j�\���)՚4/�����:�#�4�M�"iNV&u\OU��(�?O���͝Z�LW"9���Woo�+`���\����2�o=�v:*f`@YhDUݡx+�ʱu�4�Zȷ3[�X�W
}��<%���*bi]��R�tto�S�$��N��闟 x����.3d�K��u��]yk)h��F�_Q�d7������}z9Q�i�c�M��r�����ݕ.�7�����[��ʤ����箯�ƥԱªcuM��s�XRi4ԭk1^j&b�C x�6�l�!�4��e�U4��M�nu��a\�X�����ֹ��=ā�@��V.�4�R�ü����K|�^t����SYM,N��D�0M�V�p|zn�D��[4e���ol��ʱ�%m�ĞU�#��D�oQ�oo��NkΈc�S"����7)J�m46��\g_:�F�s���x.�O\gqD�j�w�w�e$Xq�Z��j�0T��dYRۡ�z�4�ۏ�����^�GZ�RΞԲ�N�[,�ز���Jn�%���\�9u,4Z%ӓ:n�P�6��\���\Z�ek1��H֍2k��u��3d{gf
��FӁ���M�� ����PͩXr��g5����#�?�I��@�v�$*\W�$F#�9�}z*P�O쵃���O*�n�j�Ayuz��4����{9�*�� ��b���И9��zf�B��Փ�"�K�i7�S�7�I�<���ΡX�V:���y�^:T�#�R˦�����D�+r��CKfj��*ZHݪ"��b�5��7	�N��}-Ō�T��x^o1YA���o]�I2��?XԬ�+�jE���z3��.
��̱�2Eׇ��ӝh:
��z2���"D�m�%d8f�2�e�r�ڑ��7ͮ�r�s��7�:�#���5�ș�Z]DB���&��N�u�W����#�D�TѠ"�{@�&�W�q��i�`̤`��6�!!��
$�f0����o����\5+QVU�����<���N^�Oi��	�8������*R�J�xj��Ԇ�tA�9W*ͥ��V�`V��m��i���HЧ��
�{+�].����-ݬ��细�t0�W{�Et��Wt*7��9)P��-�(�:�K�K�̧��"лD<��Ih�����p	P�Gt�+7iɆD���ĄJ�o��\f��쮀U����;�O��Y靮��:+X��-Q�]�wT�n�:�1\����`�͐�������_UW��}�ξ���~�g����mH���dp��B;5x8�\���1�r	��n]K�[�>��Q�t��cɽ:.�%I�:*��l������âО��F�v��e�yu9������s8.^eB�oR��`w�	�7�����2+c�8�6+�[����x�<)�1Qء��O��0�uJ�c{�~4D�M�&I��]���� Is��
b{��:"��m�Dy�Q��7��X9��ۼ�e�l�Im��X�u]��oWZ+��7��sV4-�y8M�zU����e��m�X�5%�B�=�k��V�h[s9l{���u��:�(�j��ե��c�R�Q�;�"k�=���h�J�����X��e��y|Ir��.�4� ��w��7Z���~k��1)�U�P�r���3�MbD�3%�iLT.0w�Gj��k4$cӎ��Qz(E���7�|��	l*�'	�7R�[�d r�5�j��ڙ���,h�r����ٙ���PY˞oc�5ags�7�1dZ)e�����}>��ow���+���v�ǝ�z�s"����7*�V�6�Z1H�T��V �w�:ռ���03�Y.�X�dIM�ii�͢.<�����(tU���n�h�+.��|'i�iwG�ծ%�W2a�%vh7��a�0]5�:�,]�(:+�.�ot�&/Y�;�W/e� ���tKL&j�7�#� *[x���N_���߿~���x�U�s' �%j�km�֗Im���q5C�&��,�F��QNmV�ւ�VɈ)�Z�Z�AZѢ�mi5����Z*����kQ[m�l؍8ؤ�gb��í�Th�
v�mAN�l�PTim�(
8��F�f��:�tV�F45F�b�gK��hѪh�`�X��"-��.�5�5�@h��h��44SZv�h��ƬKT�A���A�i�SA���-�`�A��q6��kZb��m�T�

SE*6]����6������I�����;[N-#Y�Ĕ�!�"b�5�6���� �!�9�KX�̅QQ4�L�e�N�
�4ꪀ��&���T4S��Z�1I�m��"�mDh(�m5b[����
��˝�&؈�I1LMMM�V���
�C���b����*�љ���gh�
�(UR�n݋�@s�Iq��ƴ��-!�C�6�9�B.���٨E3��N,����Ԙ

�&G���rܜE
FD�����k�#�57&$j��v�4&Vz�U���o��[Rs4{���}{u��KU�{<�����[Źv��S��!���Ec�cB�|k}���:pu�#�����ݏ@�3��(��!�'���
}t��n<�MxV�b�ڳ�e(�.S��N��q�BiU��f��i���[^�Q�6�я���Kg����P]a�jٮUBՎ��Y�a� gl���V�{��-����*��n�=��s�m�ڠ��V�uvK^�'�#�u�3�hyJ�lK�S�ٔ_� ��M頉����_�o�;~iS��Id끪�w�O�q+#k3t�ٽ�!\���'x���g�it�[b;kXH�Q�F���u5���1��;��/b�Z�|�ݍ�p���,�:F���@���+�����P�֢ڮX��$���l�m!���O�ntu&��N?�����O�劆�r{�=l��	\�'���%��*����7X~Ꮍ{+��W��Ǩ������j)Q��rwl�=��e-h�}v��+h��|�D�,_��Y��k1�}7L�Gy�b
���g����.TLl�r���,f���6
G:�r�ٿr����ȷ���j�7���X7�$��w��f�1��R#�;v��l�|��.]�V�Ҹv�u��b��"Ҧ}�N��Ɣ�'�	{zՊ��P�6�-��W]s���jP�rqx]*GU;��{$^
n�y���bQv���|qN�=�F���'��S�,Tт��T3ba�"���"��sl���"����ҥ�z���(k��]����{�8Y��ԃS�)�6S�
��z�VKɚ˷~k�M0��}�%���rzJ�MFM6*��X�yk�&Y@M�wn��L�ʯMK.��<꾹������|<,��:_%��;�i��aƻ��f��ԃ��'E���P�a9s[뽆�J�$W�R�}����Ud�Z���F�
t< �ϲ!(l�YP��%��])]��'-�C�v���*�C_�ǔ	��e2U�5��ૹDWOK�n��ʵH�nser!�˱�N��� jl�N��d�t��em���j����Vl�
�C=�0���a]�oH�3��W1w�6
�Z��}ξ�8�)�t��k]����i�k=���d�,���iܲ� ��em�}�梫�]�v® )�Љ�ν�]l����&��4��I��3_��X{�����BPy�f�t4j�}	T���� JhYLU��`�j��n��c�ɇ�wm��(,��+��>FDcCU�ב����95u/��W0�V�����k2�[��W�㒜�ƻ���>����Զ�Z�~\�)����}j2��OA�9p�4�Δ��J29�[�M�� �֌�J���uT�E�g7]}Ω�Cfv�k��=|ՐC0h�	`�M/j��Φ��ۛ�*�y�noA��pz�=���]�47�B@ܥ^g���	t8n��3��fSH����w<�B�y,z1���z�0�������KݰN�d�F�m��C��b���1yd;�Z8������, ��W�͑���ס�T�xX��~�WY��T��%|��	�v9�,+�/U]@�/��!�<x8��3�yc�j��jY;�]��׍+LIuo"��X�}��-�1��ܑ��8ҡU��ρ�>����4?�wq=Q*��̵s���U��d[�B¹��*�zS6):���Z=�Q4��:)�=���ӡD6�3a�NJ[�'iMA>'���b��"�
؉�y1D�P��ڕU�W�m0q�����9���y~�\���7
Kd~���.ޒD��͝ZK]a�(�����ܾMb!,MH�y��
���Ų���JJ�{���IՎ��tڋ�k&()qS:ΕݼѮ*{g]�c�X�,i�3�o�a���#6��=\�*US&xP�{#4D7tM�'���cM����n^���-|���6�2S�χ!�l��J|}Ve<Fς���M��rT̾���D�	�	��f��
6a����Y�`>m�8NT5��0��+�6.���P�k�o7�R�<ǋ��	��5����f;Z�`啃�^�Tîq�N�n���e�]�q�*�V%)������p(�ܳ�%\#��o�{V
��5�#�]R�S{�i�z�rƗ�!�E���a���ia}���锖;H\�+��ejbu3��I�֩�0S��:�#f�\-��K�Y΋��	H�,�ӯ���q�!ؽG���8�8�p���tٮ�|(��1������~�t=���3��Pax�����������`U�{L�;o����#��e�*��O��v��#�x���Bi�C@V���QZ�;�gºWN�Q�	V=�&�Ouj]�=��WljIt�/����랠�[D��7܆�stI�d��K�}���9ʬ/#� ������ȳF��V们6!�Y*�*gq f��P�T��q�\��s����}��4*#�6��^v��<�ʼ���nxtÑLv��ì�_-��ǯ���+n�&�=��G���#�]73엍Eo��K]�>S>�tt���;�Kj��p��<<��kw�#�g��Z*V�)�ZX,:���l�{�h�-;ZՍ$���J�Ar�00���w��������r@�_V�t�yɟ8y�ʝ)l0*��9�h�Xj��er�n���%��Vѽ]�;������))h�S(C�I��(S�VB�tn�h�ڋ+1Ny�Rȗ�=f�Nk�5���;I˺FB�:�'�d�E^y�Ѝ�����ꔺ6x)<p�0^e,�٦�"�i�uz�zv�#½�}�ol�u���Ͻ��+B`i:�VU��;M��x�H)��~uK��7G���t���^��mu�~[�%�k*w�%�)b�-5�58˪��|	8��`�|�3��YqO��������������J8�������;jl�U���T��2��²W��	��bW(ׅhTb��B�ݸwֺ�Oye7\�ו=�xd�2���b�@��`�L۔���!��Ԛu�t����|j���Պ���޶��]6��Kx�@m�;G�y��#���^�^���5G�vm�>�_
,��;�3�]O{q���oE3�WB�O�q;!wN���p�8s�U��BC��`vBp�U�j���ɸ+�ɕ�1���95��r��Z��0>i��"3g��,��&��s�����^��n=�19S7F�͛
���
��j���WV�sZFҷ���o��A O+j�qeD�S	3�7�O��$$�9��=d<�'w<U�;s����f�\eC�{�_@��Ώ���s��!�P{ďW���B��}j`�:����)�!ļO`��磆]y�����p���<���{K�`����+���H'4��_��gn����':�5�W�;�:�&��N:K�C��<~�Z�^��t��S�=��ĝT�_�C��_��⽖.��<�мX;����X�����'�X5e)Ѹ�8;��iْ���HcӭX�����mC�0�����U-�2��~����.{]~ʀ7�(����.�ϰ]��)��	�gU��;���Ʊ���;���Q�{���wV}B]��A�O읳A�E;�76��C@Xu��.�����ϕ^�wϫ^�o�Ūf̞�YpQ^�vk�͡C²��8�K����=�k��~����"�@���{5o�~m�#�~�^/�p�9.j��΁����v+���L-��o>˺�j�v��qF=I��$e�����;�,��憠�1��
t< �(h|�(��Ʒ��Ь۱u��g��_��
o�ėx�Ѣ�¶�-��I���\��g%컬��ქ��s�����}FC4�}5���U�oy>�9��yA�dq��� �rnVf.4-������8��n��<�09���r�*N
ŧ:���^���t>���W���Q����ޑ�A,�Ѭ�wMɌ��,�3�똤�'�ִ߲{%rF�У}�^A\��6����+����WOm�1�.��Vnny��~%ǲ�p��c�6hgݕaY�F��]�������	U�x�3���{>ix�'�n��������:�q�%j�9�����>��QU�Ox�B�����o	��y?u�NQ^��;�W1H#�v)#:�Z�u��{�BEϒ�,�u�����ت���Fy��CmU\ʬփ����#��W^N���6gl��kQpc� 5�	�^#i�,�;�)]����0љe�b�d��܃b��$�U�0עX�vKN"Oc4����'B�{8���E`$���T��cp��-eRSbe%��w#�ҽ����8פx�Rnn;��0��P$c�|� w�
f;[km<���Z�S�}?e��>�9�s��vbu���r��ӰG�,�_Y��k����]A��xL�wǮ�?�>�l��+CO������fkdb�W��'n��T��>����pҫ��l���*(��zt��߭=sv��w؆C�{�g��KB�6���IeZf��)\����7����	��$��&��ʚzգ���"+�um0��4�q�4fH2x�d۵;����.���;��Ѥ�b�-�1�>H�z@k����>�ǒ���H�X^^u���I���f���2P�
-�!a\ۄ�۾���h  ^���+�gq�xN�ZRޤ�&3/�Mv�3q{޸����A��m��t>�~�*�^�O����q!�EG��[㞯1~nX9A����^�C�K�hB�z��b��2�y�Ө�(�f�DK[O�y,0x�o�Jz��:󓝸y�}B���a�K�Ո��e�68c�vO�J⪥��	���.�F��3���@�C��]W���y��������gb@��½�[����xo%�Si��/G�|�9��~}��1���TƬS��*cSHU�&`0w�9��|�����V*Ľ]�}.f
���^{p{�޷��	�c22��ڪXewe��*�S��,4��G����NqC�y�<vw�ʞ��H(�!����l�hs�拻g�L�q�H�{=�j�:�>!�e�|�������T��b�=����:VU�s���{��.�u]��Q��a�_l�0Gyx[n�xkh�Vun���s��4ōpF�ڍeR�Ý��@+�idt8(0&K�fKF��.b�vߔA2��N�
��[��s:�y͌8�Ӿ�p�V�������T���&vq�Ya,=E9���,��m�s2�p�Qt�;#:.����=+��u�½�+�ixSY�q롉�u����_�����BCmT�j���ƴ�SP����f�-��k���T~����|%4�L����͊����R���[��G3Q��e/3�|���������88kh��f#���-$n�ڕSS��|�w�c���͟v��un�I��ۨq��~`v�ֆ{�����@�)UJ�V�̈�"�/<^�t���o�P]�VM�N%�a��u�@V?�~�\�G8�؇�0�)h�~�[��;g9��.�il/��Y����ۊS�����
��t���%-�e	|cɲJWٞ�ol�{݋S�D$w��^4���!9���m;I˺FB	�� �2�ۑ.�t�s�:����q%�y�B�����4���[=���|=;z�^��:�����}��[ӌ�<eE��vZ��:�Z|N0P�#�U��y�꙯Z�H�]l�g֗+!�j��q8��f,�U����	���"_P��lp)���p��c�,���v���N�|�u��zT�č�j�Qy���#܂%o!��E,Ӎ�˲�k�i�5�4�v��*���ؓ�R�
����]{�wWӳC��f,u��\���Ŵ�,H���T]8),S�ו��&�U�L��u����Ķ��Jh%f]�]n1)�ˮ�O�:�$pڹ�~�k�>������T��]3^�%��t7;'���5�j'_��;�������ܖc��#� �T�����fR�ړF!����l���58��@j*�sLb1�[v��g�V��5l��� �{�{M{�z�{w�Q����m��]�W�I�pz��8��d~Nd{ȧj͊O^
�{O�vB��[)��S����t�p���te��8���Kz�U�'�ܘ�MC�&�G��v.�ഺy�롭�
�Y���)�uu�gJA{��uq�5{nK�הκ|1S���42E��-�����0u���:1-�73��l�O�i�6+�����L�jRe>[��,�[�Ɨ ���"xz֦/��e{G��a�ѐ΄����(�Z/T:E��e{LD��_����QD���V�Ժ��0�T�d�:��wm�3�*=P�J}��׷�jN���C�0���w�AJy��y.�$1�t.�h˾ʰ� y`5l[h.��8�_�5�fuYe�y�>���T~�v7�	ư*�]�vͬ
�u�G�FV��K�~�]ìY���s�ˡ
S1ִw�[�*��_H����e�H@A�C�R/
F�J�`�ƌ�wd�x�Őp��+:�n��9;o$�wL ���ei*ྵ)Ij�cx ��s��P����"�̾mރ��L��vgv@�ϖx�젨�b<5��m�Ϲ�t�k�vZa.t��7�.�]�ۚ�7�C%�s����}HS���^;}f��q�V��T�A�u⊯��a���߰�I�g!{/��S�E�e>�@�'ll�X�wv�/�̜󝳗]�'l۷��zJ��|�9�O��r��-_f�:@����ݹ�t�ʹ��y��ͱ��V6b`.�d< 8R&E��gm
 t�{��$j�nwi5�5��2�%ˀ�@{�P7�
��'�.��YȮբ��5�x�%ㄚA�/^�]G/yJ�:�V�1�ZҺWxQ�y���t��8��;���o\ k���2/���'{J=�̡��ľ��H���H���K��e�_�$��d/3a�)�G ܚ��$�8^(�F�/���HdMTə��V.6���(+�V�w	N�>��8�k7[�	�!��0eM�{���`�M�c�K���v��i+m�Dm�isL���:�9� ��T��u�SΛ9��J�頛�pky�;r;����=G�k�6j�U�&��)���h7�3'jvr�W>�2욕#�)J]7jn^�U���חf5��ۣ�=kU$�T�Z�md�{��T��J�iTFQ�F3��Z��IU�]�K��9-�]-B�9�V��]9�b�f+�诫X��_
pwP1챘���s�)�H[b���u�Һd��o�ޢ�1q�E�;r�f��F8h�8��0��X��uk��uIMH^�h�ޞ{\���v~��5�� �:�#n	q��+Y��p�X Ù
�;��Y�wy�o&��AF{7���c���kl�7b��ŵ�U�Lmө.��_u˕ˎv��GV��ym]�)ӲF07l���q���B������7�k^�MO��8��J� �����A��ם����V��s���� ,M�:�庆���>T8��e^&
�tכ���x��������3_M��[�P����ƳѳU��I��s�� 픲�n,�ʃ����WT�k2�4�Ki��M��iv�Bkzt�v��R��eJ(N�zۙ��#&�
3��\<
��a��	1��bT+_q��c�&�V}�9�U轾���o`]{�r��V���23���A�F|�[\��W�\N��Y�Jc�]WWy�S��yx4_ٮA�
bU�r-Չ䮮��	�y�$�⬣�y�ASwD uz�"��*��C�pK&�E���ѮO�F�4L�r��i��6%鷏m	P!T���钰NV��R��n�b]��
dgVUc1�V�]�M�������2��Ƴ�j�S�>[b�M�(h�����N��5E%RD���E$�)-�@UQ��Qb����h�������lglE�I���Z4�Nک��5TDKA�DI��D�1P�PD��:����i5�$���6*""�6�MMR�A1I�QD�V��V&*i(���
�3�m�*�-�:�Hb��"�����DDD��Âh�Ӷk[j
(֒!�*��ւ"�"�	��6�4MTD[bh��Ր�T�DIQCkU1�[h�-��(�mb
%��*�j����v�EZ�IU0�b*��PPUƂ���F")���ժ���V�i1:6ư[51Q�SMM1�m��EM�4DDQ�EK�"(��+N�8*��T:b��bf�5��J�:��)������|�z�����~K�P�j��=42>��a��E�gV%D)���90%cZ뫻��vݍ���#N����궗k3�u��H���u����#�Jz��s�7|N��u	Tw�'"�G�r�`��N�o�Q��^G!+��ܽ~����xyQ�.����/1俏?|�.��;?y��'��x;7^������b�8٣����������^G*~��5�^G;<������?p}�����Ka����T��`������a4�u��;�a�9Pi�?I��s����}@��_?O��?L�/<�����󞦃�%����\�K�}��{��w3�?}�;��4�w���y�4?`ѧ�0ww�O ��z���uu%%�g��|�c�����
O��;k�;6;xPfh�!`��M�/:3d�E��ڶ/��ٓ�������4������=���J��{�p���ϼ��>���ܼ�{���M&�׷��p{��4������^G!���	y�/��5�^@y���g޿���淪�����tbi�?����������Rg�����C�������?�$���Ο���$�y�$�~�����qh��:���|��יi���>{��_޷h3_���h��C{���惭�Ƀ�ge�U��W36;���n�٥�/q�'�c������<����.��|�yw���T����>A�e��p��&�e�����_o�������{�|�4?�T�>��|7���:��ҁ���i�݈W<��������jv��K�P��A�>G$�}���u	T�'Fܾ��B^c��5�K�?�����.�~����?!�:]�}���(}�G�9�K���&�G�ί���y��d�v ��X�k9}�kv�:y3��W��t?��s��'��T�?���>Gpu����S��A���!)����1��p�OgX�P��C��\����_���#I����nl��Յ7ڕ�w����Nއfǯ����̾G!��޸З��_����ޟ%��b>~���{���>}ߠ��/Sʗ���}�\�����C���'G'�:�����Ruy$>���e�߆]������WS�Ȗ�.��;��7Q��9��u�Zt���/e�r^��q�{����?����J��w�|9������>����%����GQ�^�O���?�r伎T}y����^�3yo�Cb�<�<���\��Ϛ(�%n;K�ol��n�44�
���voYPY�$�������u��k�m.�F�>8�'^]<�+��L}2�D���$��5��2�f+�*��q��&(Qw7�c��EUԿ���"���4��4Z�(�ͪ3}�vZ����@묿�#�J������˓Oa���J���tϒ�d>�ty'#�~�/}�r}�d�~����!(?��q��~��[�r<�� ������~������������C�hi� ~�ט�_�=�ﾐ�W�~��G��q|�>y��!����<�P~��t~��_ ���z��|��=�ۯ;������{�O��BQ�l����A��<���9���g�cI��?_��<�GØ��%�����p�[�~y�Ώ��]�ny��Ο������vj��'�;y���T��Q��{�J�m]�d�6;x?�÷�ۙ�a�Cy��!�r��x'��	O�݃�u'/`�=�E�~��n�/2ӣ����{���r�0�{��a�}�q���2ަ�vkv�=��r,����m��nr�Z���������w�#��N����'�O}�P�A��y����A����\N�y�����������i��˓_vB�����0w?��c��3C�;k��۝��i�,2g�k��mkR�&���~����U��
���QP	A��z���9/�=����=��N{�c��.�>{�=��?�i��x���hy�c��^\�	��c�z�C���~�$�K����~󫗻��>G߼V��b���{�b���}D}T��
�HU|�|��s�u?��y�~�4r��;y����=�����A��z�|���^���q;���&�'��伇�o���=\��9;��s�nu���۵3�8�Fw��k����f���O�u��p���Ժ�d��/�������'��?߽�;�O�����u=G!+���$�>I˸9�=�� ������j#���|�eg7>k�)4T�ß�K>������A��B��*������Ov�P��A��<��B]�{��^�~˧�Y<���~ܞ�}ɡ�}���|;���~����&���> {���]��)��u��z2jkam������.�yr=~~�P�%ty�ߘ;������S�rNG���}��)�����?��%�X���}��||�u�{��~������]��>����#�N����B���>R�u�j��pa�
U��A�u���9B�H�i��&���x���b���^g*`��2�s��V-j���VvJ�sq��2��dQ��t�l�s�b�L�l�ЀϚD�Ǩh&�r�[�Q9��ڰk��W��d���U�ҫ���0n�N����%S�Ss��h�gv�۽,��ϗ;�|}�=ˣ�z������:����~����N��'ϸ9���d��	��=�F��}��)�����>ϐr^��T�`���w߿߿���O�PW�Xӱ0N9�����j�vhv�;�����4�M�]'#��^C������:���s��އ��\����'��?��{�#�^N��v�c�}�s/��l�����9�`��O�׿�}����vT��N��MZ��1k�?���|�}��䜿A�����T�Pt|��G�>B^��q�^���y:�i��/?��� �	T~������r���>Kʟ���pc��nO�q�A�]њ�u��d�I.E��n��fO�ݎ�����yr�^��p����{/{/������S�a�����hJ�:��Ρ��'�w1�Ϝ��<���~��ѡ)�����~G�A�K����BsV�ӵ�8�қ�K�����١���=������^d����N�9���>����z�i
y�� �4�\�����{�G��}?��_$��K�����Od�>{���G ����]��}n7u3n�/��u�t�{(7�?�ٱۦy����%���>�s��$�MRh4?��f�����:�K�����:���~��|7|�A�:�ϭZ��o[�o3�����jc���/,�=Q q=��e�Y�d���;����������t̿�ﻺ���~ܼ�'pu������>]I��9/g������9y=��BU-Q�~����:�<�/!��_���:>BS�r��|���r����"������oS�K���ݹ��Kߘ~��~����e�O��>�ø<�������������㺐�����r�9�C����v��~����'�v��lyu4%P�ww�����.�;�e���G�yݽ�3C����_;O�{'#�=�|�����M�� 7��O���O�s�����ǯ�}�~@u~��ߜ�g�yq�<�SԻ�HW_�Pr4��?`�~��՘8���޶��ٺ&�ͦ�?���ۨ=��yw%%:�nC�=�I욯���4>G��������O�>��? �c�������|����xU'�4����`�������>^��B���������1/�?M��2�h�����}7.��/��M�y�Q�e���+"���>�/��s�^
vj�sgq��*��e�c�[&��kJ�u:�f�_J�[�)���r�֯��}\s>�ƶm�������W�¢΅��;�)�{��9q�>��}u�rNG/����=���WܔG!��X��GSܺ��_#�_gO����}�y���_�uHP�Og�?u�`�a4}��/�r}�I�%�������>�R�;��SK}Y>}�����{��Z/{�wA�%�{?�rz��yA���:���r|v:��������w�z���yy�?Kʞ���@y=�����y.��5��>�;K���ݚ;'1����D��Z��֖��}�~���/#�������l�o/N��	O�v�^`��hJ���NC�0r����XM>G�9��a��S�ל?I�A�$�w��>ï�u��+���*���mCGg{����2�	�%ק�|��4����/3ܼ���������y�>��K�s���C��]��=�ܒ����>�#�~��*B����Gg1��a4y�{���|�K5p!���M$��uڛ�$]�b���Kj�&��w��6��y�f���DW���9�`�:��9�s���G�ݛ�~)���{*V���v�F�Lb`mI�ҍSF�6K^�.$I�%����g<�l�����]s-b�ţ��.�$��Z6��ɦj�l��nF���y���eq�.��2)i̇�ƀ�eW�i�����/��c��V��M���:��*)�b��/��/�5�����a��z&n5�C�{�_@�*�|���C[��秧��]Z�V�ak�U6�ی&7\�m�3��.����ƆJ�	8]#� ��������՚��|��7��|��ٝ��� �1g��;�M��M�٨�(2�Ȫ��oo.�t��J� jr��ʇűZŢ����N���^{/3��x�&\.�%[�]��u��}��3��m��y�j�3)��̳ի�L�G�RĹ���+I6��[vrn�d���W�I���Յ{�%n��,U���m
V'TZ�2A�>~�=A�]�'	�13�wyxo��@���Ma�M����:�^^2�b������|�i��2����9�g6d�^�8��/h�)�Έ ��}�q,�j�T��AJ�C�1��j�D��Oe��x|��*���}�&�v��6�T��6]m3���@�a ��ZxWW?l�k=�?�y�u���F_I�ٷ�V��^�R�|�uƇ�P�tJ���(VL����v��������e'[wՂ�ڹŏ�f�Sp�����'�Ґ��Z>�:q�v?3)�ӎ��m��q���m*���j��֌2�����}~/����U��.�NK�@�A�{^#��!�!\J[	�{y�*a�+ٰ�Q+k��45!$��U�	�pQ /�ep��w5V�j`�ױ�r�W��<�Y���Ox����(ߘ�U���ǔ	��e%Y@�EmM�#��z7�y!\}f��B*ݟV9ѯ �a�`Q���=
�f�o����|*a{��E�`�<�猞2�]]27@��gdB�;{b\��1QA��*?��J��6�꺕a�����Jݒ�և��ҳi����;8�m�b@���ݢz��n"��Z5�3�m��V�l�g{��Y�Y��EE|�[�Y��J�b���0rJ��
���ki/�d�3�J�NJ�Sy�3�O/�W1b���7c�V�r��_`�P���^��OQt"oy8�}��g�-6���^�1�o=����В�x��k���?�V	=�w-OA+�������/l�u��ܠ�2@Q�;�lU���1�>'E�K�����9-�����̃6z�+&�'h\�c�0�L�A-�5��޷�=6j�ƺ��LX���Xgj�/�ܿeh�3ta{�10��KF���T�'#�/fK�.��%>���P^��ߔ�|��\֮<�e���8�C�p�Ԗ��G����T¾����e%�ӹt����Ln�*�[bu��ۧ~�S�?Jx*ㄝ� wIࡎ���KB�4o^^��{si>�Ú��q�Ft���9]tE�іE�C',��S&��?�61g�`L��nٜ���o����y�̔��7�Q�[�q�z?i��=L�*"�y1�>H�� �V*�{��-?+}Y-c��~��2o�n�Fbg�b�5���T�-��vH[sng��J^v(�����ڈ�W�#3S
v#˵�acy�f]�,eG���P_؟���C�(q�z���3�E/�H4�}��Cԩ�$���}bA�[�*n���@�+���R��Mm�����×rӺuY�m����l��Ps/�fL�T��huaJ�-�r.׳{�}�ze�B:t~�*�-���ov�GqL��l���J�z?<�S�����)āW��&�īgv��y�E�dNz�;j��N�Q���:-���ڊ� ��h��ySR�z��ȋ/�q2�x��6�>u~f�v��)r��*�����;���̞K,3�s"�/+�z,����K���4��k���vPY�漮γ½�U�<0s��`��vloSY��Y��!����T�y�<��X���k�
hp
��x:�q�վ�Y�uK\hzZqVm�v�6=:��3$�r�M�S�il����}�����!�sf��پ<�Ӷv]��vcϛ�]�x��K�7^�J�_4T��_*]8�vpՍ��z1V���v�(Q�=Ih����6.��=��8��]R�Yǁ滃�ܗM澓��c�)�WC�1-�K�\+t(�����N�sz�dK������i���|����k�7g5l�~�W�W����]�.,P�~��Z�Jin�>���]~�=YX�5;�JQl�p����d�r���o�juk��;
�Կ,���&��r� ����K�}�k]ӫBu���Z)�^ІKp�L���y���Vi5+Fmu7v�$��k��U�9.�U�΄���E�90�Am�Z�X� ���D��{�s��v�UNi~Z�\.U���;��a��=��$�*�����%����`?��f�(�I�H�*��A��;�
�!�U�L�����w�mь�P�U�-�LUe��T��P)lӝQ���t:�l���c��!s��s���"�����ȭ�u�+C/Ԑ����:*P��N��٣z����;K:�{�Z,�kP9�Ā�؛]�V�:J~y������#}���|������{�<�FBFn��PZhQ�3���ᛅ$o����}e�K�z�h<�`J��v����Z:
�3�ӧ~��(�U��E��n�♜�/e��	��Hv�xb���>�rƨ�2F�MP�k�i't^N����N��y�����tR���%	���^`�y� 5���0��(v���՗�K�1�2ܖ�ճ;��>�zZچ�x��=�~�P��}�K�;"-۝��ћmH���u��J�p�]�<�}�)�T���:m�(V��vey���c��&�<��叭-�^o�=n����$��.�s��N�R�a�q5�h�����=�0G� �[��S]�_1��꘲b��k
ά[Di9�7f��{����ͬ�JE�	�\��Z���2��8��-t4����1sPId���W?�x'�����b����欋�V�S��iq���`��3�[����nIw�F�9n��fФ[����U"wPV�,|�gL���>�@]�������N̢���(X�M頊�8�_�ܹX����gF#s0O�dΑ�*}����f�ƙU��}�8�����`wv�Zһ�ZңS�׷e��Z�jQ��P����xe���λcC$XI���Es��3g�^Z��Rƻ�~ar��)Z�-�T��)X/���Z�H52�)���'����1��7��~I���D�@<;�liq��T8���a{����Z/�⽖/�"�[�W�t����I��z��Q�J XTN^:���O[()Q��	{zՊ���Ms����w�mU�3��|埡j
�|<_�D�Eʁ��C'}��j�]�Z,{_�UK���AOJ宵gC�"T'�nR�vs�f������ⴊ�,&��=fS5�ʦWv�S|{�b'��\��ڿS]��l�'ir2Jq޼��4K46�,�!R�~f�j�5�EIR<�?t�k*�p�U����$�6���	��VT���P<��Y�V���A+Aĭ��[���;� aJ���#p���κ}wj���Mm(�o:�U�q�O�Qa�}ݗF�7�d�U�ħR�0�Sۭ�Z�&����:�����7�>�ܘ�V��h�͟�官�e�{�A��� 0J,K���%Tx���4��/Y8�"�9�Y;���������H����L��y7"�R���v٩����ơ�[^u��q';DUf!
������߲x;�]��l�cd���y@,�J8ʑ{�����,�#��\�{8�P{�<� j�U�ʳ��B��׈7!�`Q�����+���蚍:SM�4�Z�U�r��,��|��G���bq(o��(��P7f�SU�,��a]��c����jQK���[�Yc����ں%�/9O�sSH�I��CG�~߰�-N+Ի�����C*�o1�S.�E��� ���(�3�e��1୭Z���f����`
�(ѫ[��+j��3�`@O�Ơ�T�>CfW��/>��G0�\�A
�뼖5L���d��8.���i{UG��4�����e�X�%r�{)�ɫ7y*��%'uڈ���G�������p�RZ�L�T��7/eRbe�y��;C��I_i�=V]�Xn4CT�c&ih�9���Ns��5���%�Y}�DY$[���Ƣ8�>���rbegAn����ΓigMN��`V�#����S��M��������G�j��SQɛkP�4$���\�=-rبQ҆��s��lҭ�9�iP�76�uo>��?���J���jp�*�충�ӥ��5�|�]bpj�gƌ��bهk�]eع�y%ʽ�V��j�����ˮ���ޕ��}J�j�o~=hR�*�cw��[����6��[i&Dハ ^�b�>ȋ�=]�� ����3�b�Ĭ<��I�C�
�5��!���b�iv�mDAC���ۃx�J�BfG�����ɗ� ��bY܅�0� ��nWju�9wq	�����Z{>e�a�������l�;�yvH�n�Սx������{��p���W�n#��Q{%:Z�~�+XKɸ�w�jDT�ڦ'�U��s	��Έ�YM@m�
�Xn��ڻ���+e��a_Q���X�|.�3�ժ����=R�2Wr�Mc���ЂR��G���)J��6���R.%a���{P��ۼ-!�S�j����{|B�n�����_Ol����B�X�׼�rs���ʷ���Д˦݅��Ħ|�k65�yi*�_k��{�un�J�%xD��k6����o��=p^�5�at��y0q���&�d�����c/ 9\�r�N�/�[�b̐��S�j�����ͫ"b����|6�!��LެF��H���$,����ܳ`T5m]wt_"�e��x2�E��p-���c���mwl�U�^gT-�u4vy�ZAYV�1�9i}��ťk�D_'�mᮛĊ)����Ef��t �K�T�	}a�ś��m���[�#8��4(�u�A�b�3e�����-\T�w�oP]��4hu�2Xx��F���ZD�PY��6�:�q��HK4�41�p����X���kV��f�M֝�WJbu����B�!e��Z�����N�63��Ï5&)9�÷)D��۵�q��mki�a+[�{�(�Y��������gu���X:�f�Om*��Q9���n%��R���M�q)��FgP�7kC�E��ؙVp����E���a
L�Zɂ���J�k4�6�X�,�Z�>*\�;nY��7������۠��vM8�Qa#]�򙄌�(�V¦F�j���e9�9��;X<�y5[ٽ(��Ζ�W�K$`���!��v�3�])�Pܽ�ƚ�e��hvP�y������� �Y�ф �Aז"�-&WJO��g<�ns[�c��)?��vn��%��D�.$J�	�շϗ��mhRp0t�[��ffr��:�3zZ�=x�NIom��ְ���/�٤p�Z�� ��5;����%H���6��V�T�%��N'[�����qu���t+3�����@T�0S33I[`��"a�
��Nh����Պ-��ckV�5Q���E6�UMN�k&	����&q��Ech�*�`����D֌QQUST�LkTV�U�Fզf�-��&)��؊&�h#m�DZt�F�kUQ�[j�j���c�1U3A;��f*	���AZ5M4ET�ӣuP���l覩%��j&����K���mg5��EE�j�kAlTF�TQD�k�*�"*��h����5D�1S1S51A[��(������UUTk[��J
���j��5M1���h��������8-�Ɗ��ի*f��l�	�ъ�m�h�V�E2P�ASTT��ET��h5�����&�(�)����5���"�֚"����uF"
��6UTF�bDmIm�5�jnY�
��堈�
�j��]X�F�M��Ǖ1��� >&�41��%���}�\�7R<Zz)�Y�I�j,�*�U�^�w5�,S���U�ǣ�X���7ə�,Ȫi*��\��ꪪ������=l��mȿ��S�h3C�r� �a��7@�Wi�#��ӯC��r|�{�;-��36���D5�b�����ŉ�%J�[P����f�]A��ω��l:��C���J�F��tՈ�Mz
�צ
�h£ +!�����������Zɴ���ppa.yr}�,z�1侼��mןN�$�B��+�qL��w
)�Y� �f& ��6*0�ȷ�j�gp�Bv���`��f�k�i�R+�T6�'�\������褲���WZ�먣Ŕ�zP�a�*�A��N�v��]	���v�q�<����W��9������~G�g���F5CS�˗��lpǻ'�	�a����Y��ݘR���u�;���P����تa��� ��eHoB�s���N�߯��q�[U¢�onė�V&�zFe;W��c����e{ʘk�
vx�`��0�:��q����&��E{�v�l��\*ī�(fI���`�R��ڪXg�u���EDGZ�f��i��?�g�ր��Rس�L�*u�5ܞ�,�h�Y!��3Zi0�A9Xr��nm��sEt�C���\��/F���M���J��z��|r�db*Wwth�����tx��vFI�C�\̢C۸V�;o����
��S�<;�چ�����n�e�޶?{���3�%4U����6-�\F��4���h��M׳���y|�S}�q������5�èw�4�M�|�-�a���]�ϩ/3bU�{U�qp�4��g�c��W���l�I�C����&8��|�]i�ɗ�Vں멬������Mg1Ǭbc�a�������Wv7m�i���y8E��������k��h
�~�Ek�[���]9��,ᣘ��2�`��W]h*��C'�kR�r��,f�\��%�����C4KW�p�L�b�L������a92�y�KeX�j�A��0;�kC%{�}�'�r f�W���H|2�FǪ9O�L��Zʬ�~ߺis��#M5�tS�p��Z�{�S8��a��Y#���gN{~�oP"�WE�@z~ysxN�ΟQ;�S�z{�L`D_���i�5���]ƭ��kiS/�_�I��䏏"Ema#>G}��O�'���NH���i�N\i}�霦1�F�j������= �����ca��Dl�˘T2f����4]�����a5�\���Q���#Fe-vl����e*��V>��n{C�s�f��߷޺����7��Y����:@v�����5�H+K��O���Ӻ���hF^��nH���ݣCM5�بo3q+ѐڢ�<�ħ�m�돁=�2�wz��л����<c]�����}_>�7o�jۉ�ձ;�@?!	�;�;�۠���7G����<�{�3��v�u��%l��e��&;L]��VR{d�Ԋf{A�<�P��+b"_)����@l���|͞���
��~n�OA2'1��2=�+���[��p�X�zA��g��*�sa��������.K�}��U��h;tG��Xw֌;����oӳ+��ړN�q��h�4�u�(�SRu��i����(��j���|����#�6�������Ux�w�4F{!Xg5�Լ�.�t�r*�/�V���\3�^��B���
��5���M�b�d��Y��j\:f��7�2��Q����`��ƴ�|Ot+������F¢|U{=H�X}��vr��d���jk	 �֣R�U	�F9{ة�f;S�� cpO��v������`��X��hx<Y�8j��6�+��ut��^�.^��h����΀���k�וM����&���族���yx��}���vP�Z�LԹ��E�}O=|R��G+�6��Ҕ%���WN�����K��`Nh`v1���"/�I��w@K�����6�����X�i��>[Wˢum	A�U��Z��	�w��5���ǧ�,p�	~k�ű���A4%��ə���}SxR�_ftgI���{���l��I��"��q�K}x`�3�k��8Dǩ�fJʔ�%�$5��ڱQ!ޒ�1��6�Uݬ��R�����
��h�u[D�E�v4	�U�����o�����X�+Uq���t�_-)��b���2���Ⱥ�(v���iR�=f3X=t���Ǝ��S	�/�q�L��vo�w{�Z�{��Rv� g�S��Э[E46��;UFz�q�e�s�1�jf��D��p��ڮ��w:�.��z��7���U\��T��9"�ã5��O1��f�4��ًy��C$Vlĭ�$a����IK���!2�Ow`�ٳJ�m���$�櫎�m`�C���?;}���b������I���ھ�.�t��� 9q+5��7�V�2�5��b���DWEyJ�~��C����y��A�W�~�M�z��pk=q���3\�+�n��|���Vl·?1 l����	
�MW����`�H��oo�Ş���rn"]�z�K'�!q�(bڢ_t[b��V��>*�ˣ�e��I�u*^j�eλۙ�\cR֝�2k}�'�3gl��=��=�-�|;��bXW�ʟ��â{3s3�Ηc��@|G�酉��:��o8ڴ�خޠ��9�n�X�f�=/B�i�`�4`M�m��Oqu�N��Zp+�
����SzH�W��������YdF�1��"-�ᓻ֣!�T�@Z�aدgEJ�[�*�b4������z?R��*�Rn+T��)n��F*�m���}��An+�'�CfR4��7�ٽѕ�h]j�lɂ߾jP@s�F?W�!l4i���f��.(r�d��N�֊�!*I�j�`�ǭ6�YF��g��WIk�2G����0����s[e��i����&��e�1܌~�J��rw��W�	:���Ht|��͑����x�OjM���y��Qp^޼��!��C��P��ĥJ�[3�C�����XL���^㠰�����m�bg��yc�i��	Sk��Z/{�F�+ب�g��O�<�i q�`�l�L�X��/����f�����}y�|s^}>Ҥ�~
-�!l͸�$���G|��{��f�����N�U�o㢝#�l]��0f�X�{g��1P��(״�*2�Zt�+�Wx^UD�e�"٣g���>�k��r���7�pn���y���ц�#�A���?X�}�C�u>7dY��sT����e �0ocB�h������I�w���XFl���iΆ�F�ÜUZ�kPi��T�j.W/6��M�׊���a���nJ�	u񕨮6�"�iq����S��6���A2�Lc�㓻���o3y�a,��rSZ�ݱ#���'�����(�N�_c���v��/Yp�����+5��k|�o��;)�܎����%�^>�?yx]o�R��hk��Y��x��Qv'aeiZ�T��&&�V%:�ّz]���O�L�&�zm3)ژ�BPd9Z��!ծ4)��m�0w�A�+A��Uw��iyhN�����WJ�Ԧ{³(�{p� �R��ڪXey��u!��)���W��S�[qJ\����O�ſT����v��d3R����Ǘ�2F���4����6yFDMgi���q/�֗��(�cڬ��:`�hl���#S�:I����D�y�ʴe��\s�Mh��ޙư@p�
��W�a�^�g1Ǭbcݸ����=CB�ꚛ��c%ڙ(Hm��u���"\z���\%4�O?L��*�i:u�����k�3.ذ%X��2z6���^X)��N�i �� $G�M��fOa�s�����щ�FCNG�*Ŷ�t-C���Y���W��OW��>s���t�+�~ܫw��������/!(9��5r^N�_yx��x��X(��Z�=L�a}S����՗ݗgJ�J�u��5�k�]M�>MQ������cf���Z�fW! 7��*�+���y����*��N]�������5�8���+U��C�UK�Y�=��ӽ=Ҝ��7L`����P��,�T=�S��̽Є�,~ξ�n��3���+մF:�����g7��L����:�����+��/ ����w;z����^�~t�t���<]W4Ek�H�0�ׄ�+�ƻ%���fyje#Hy���\uqG]���'Ҽ_Թ���G(��e�i�8<��{M,Hn�t���;.m��a�U����Pt�ζc�ڌ��	��"��uKO��P�0���_,���%�}2{�%q�EKY���Ng֙#5"���wO>J�~"%��<{c�K=��=٦0ϏL�+����V�[Ǡ�]�N���uT������Hm��>�&�6��ة�V/s�Ɉ�<�ip���Q��`���^�����7��)�(ש�C,^Ԛu�*��N(��!�!Nf4]CQ	�jqC��l�_V:5l����nn>����3�o���jYVwV�ݜ��s%W�f(��nT�kK
@k�
�����4U��Ww@���:u�.sU�vm�4�����!�.���t��3��þ�V����>�ԅ�f�'��0`��C�3�����)&��(wv�+ ��ge�\뮭���jt�7T��nFk:�"V�� �� `Ժ��),�����߫������o��;����;������E_�D$0���`J�\�ǹ#�w��w]��ԖLnu�F�̞��혆������g�$?��}�^��[�x^�;�:��p��7vgSTe컢m1�����l�Z,��,p�1�
V�'WMj� �x^󹣹���5�
ח��\��0u��!�u����j���C���wT:F?�ۑ��1`�-�8�2[*jW�l�� hTOZt@��}^��(Z�>�	{x��]�>���ˡ5��,�B,�!20�5�VB�.ƙ����~N6�<��n�]��'�OI�Ԥ�aUѷ�Q�W��VB|*3 �g�,2�~_:�48��(v��j-��S�<o�yp�Φ��t��QJ�׮m?W��;��iF��JHL�S�'�)�z���.�A�A�"�E~1s��-�^&G�g=f3�8�fϼoWܫ���`=��8X
���I�{H,�]K���3&���Z����G����ج;i��H��:(���4>����^IK�����3��\m��7������v��^��\��M�p^y���͠J�ڄd0���Ee>i�S��Ɨr��J�"���ymBL���F}׍+0фغ��lW��o]<\_^�Xs�ut]X�V��;:�����'b��I����
>9h|jvk�����}_U|��JR������X6Fİ�N�����m�\��a���j鍷�UZ�TŜ?��v����9l����x̕a��dK�C���}g+�
W��^A^�=�
?Sy��x�؊�v�^�$�����^���G�>Of�B�w I�����q�t�یgcr��A�7�	k�%z��Z�OLD!�)�T�P�ڢ_t[b���n4$��s'�WYeI�=Ъ�l���dĕv.�45:������'w��h=5M�׼�|�a�vˣU<�YS
1k�;�nw��Ϭ�`�R[e���S�|R�f�)��g�8���n���S�o���[W���k�:xM5���_D�D�y��ȟj����4�}�����]��'\��ޘRo\ܘ�<��9��>��s��<_�� |+�K^�U�?>W�Z����y3J܏�;�v����m�k�	܌�(�-����������@�t6�^Zl*,<���г��Z�Ҵ���a=�{U�!����S(mqb|�*eoP�?�7(eu]���K>�i�<�Z�yE�J.�Y�^���g���<��碲�^��Ub�L�p}rщ���n�+*��|yS��MjڙXkT�>S$�,^�,�]�JҬ�sʺǻ�%X��L��pe��wm�ۃ4(1�����q��j���$��n�
��<��foyn��pi�S�/@w����<�r���Y::����)�SvCs�/�� .J����PR�Z�wr�{��ݼx�c���m*I[�B�+�}�z`	8R�^�&f�{k�\��\@[��>w�xN������^W�V��3�5���ug;b�k���z=m����w�v���4D2�fu6��?:���n̗H��D1R���%x�M����ٙ���������͝M����u��4Y�3􍑫iY���!���W'�׏<���^���]3/�BwQ�'p'T3F*�qa�ֲ�5x��9��gAwپ��JM����	���-ݔ��M��b��D�P�9b��54�K<M����V�{}�U���N���Z���qץ;~≫��(VeN�����)�z�Xe7ݗ��k��o�d�P늖��Xgu"��sSs8S4�.-��j]�ܾى\pc��$5q�����g��P^g��k�7[Xu�F�ϒ�tO��6!|ǵY��t��U����^�xNG�F���u�Mj%h�\�9����:�ڻ�����[K��g�3��S��5�mLX�;��.��ʍAֱǨsA(���c�)���x��r����ӵ\�R��gf��0��0��K�M�V����L�� �N��B�rjp��G&��0nK�2��u�� ��u�Nιc���β��1�N���2�_u��p�uՁohD�//4���0*Z&U�	%��_FA镚f*tÎ��+�����2��0L�e��,��?&W/F@}����f;�Pʀ���³�o�>�ssQW�8o(�r7��@��X�T���nK���=�;n���1#���PQ$j�G`�pSCM�9�>��<Y6�ܰ�j�<��Gsۖ�.Tvw`,���Ml�tu�}im�\�m��![��仅Mv.���J	}��+B�G�R2�b����\�� /�	��֑��+o^���Y=�g��5�����53w pj��Ea�K�X�-ŊoT���0�Y.pgzÆTܕ�����
�Rv�c�}��;qZ���g)5}bWZ�����v"դ��F`'��P��;jH��일�
�j�╅�t��eǔJA��s\�]�I`�[&��(���P�\3�3���V�,;C�zVGj;l��� ��!�\�u�[�@�آd��@��c�k����Q����r���z��Yi���GS,`���D�M���U^�u�&s��j!,�\�KL�Va�pQ��\Z�j�J�}�,J������#S�9�Jҝ���x=��$:�r��/*��]5�%��ҥKC�gi8�W�c��D�ʮ��P�-���zwTE(̧眜�t�2-U�hݙKj�gi-���@G__��fG4,W��\��gu�ކ���]�2��N�	@զ1�(WU�z�n�\Y��>YA�j�v��Z�+�ّ��n�����-�j0ķ,�,��I�����>�4o�Y{H1�����w��z���o#����NkL�uƣ�o���F�*��ܼ�cS��k�WR3��׀�D����U�ŸDmgt"�Z_c�/�K�N�>��z�&:���"��Z�ƻ^L�������鍅���j��[���Ռ;R�+�v�V�F(KI�u��j��m.N���[���LJ*%�5b���Q�3�E^�/[c��ɽ[�ɩ��� ٺCTT�X����y0��i6�xGpU��eK%�W
���)�g��vI�@�	�L[غ�Z.&���ϊ�G�Q}�r��:up���i���IG'��1�A��@�
<2�p�A4��l>Ru`����.�<��lk�}$
\�7i淽��55b��ޥ�ҙɴz���W�oٵ�nAF����u��80]2��YTw82S�!]IA;� }H�����u��ꮭlu�\ųQ4�EDQMDDEPLM[S���4�[`�Չ��DLQ4-S�LE��ULL%Qh��Π*@��$�*j�jk��*��&���&j&��EO79����đPHEDB�(�&����4�3�i ѝj((�*т����*��m�MZ�!��I�%�������clm�U���D�LFΪ��""�(��cF��-b"H��i��4QIDM�h)�U�����)�kQW6��Ù�ԒQPATEDh�E�QF�V؈�i�l�6�QLT5��QV��Um�tִd�te���AQEQAM�T�RU���(���iX"�N"�i����5LֱZ�G1�i9�m��"����4LQUT4��EPF�1ALTM�M%CUETD��c5Q�h��������j$��Z�jkZ"&�N� �b*���tQQDIT5MLMn|�Ώ����߻8v�Nx��N"�:�Z8� ���a#�� ]֕��)����;�[�YOu�w�ܠ.����_U}��T�s8�J� ���ʒ��	�مM�ۂ���·p�����^�g1ǁC�f��^���۪�ңKޗ�M�W�嬲��^*~U:�m��1ڈ#�;�C,L��q�#�0.W�G����jv7�*ǼM��Ի��*��Q��r�� qɷ�����M�����/>�l����jڦS<��K0&U�A�k��`�D=����2�a-v��"�-J��J�� /Q��P�ӎ���u�i�����2}�eC�d�#v�45�{�k��^�>��/P�}q�.V���`�6Z!�Ó>vr������|-RB�L�=��؎�v��ٺă�U�}�:W+�O%rG�戭c	�ĽzL2{�h��}Z\�Ͳ�n-�)ET�m�W����E��H�B�=
x�[3I֕��	V��h�E/;���نcUP/غ�ٲ]W����ֵ��s�>��3�
�_y�-<N0P�3ntJ�Z��y�u-�9ws�Uz�s�(2z�k�b�;�):F&A{A�<�P��+�l��[�!~��Q]�l���ŕ�&C��[.S�Ma2��hf]e*hL�H�ש����ε���l�k�����^��wת�*���(|�:M>�����\�&�.�l�ok�Ze�j\�cy�lҮ�8XsM��Q�ݒ�k��d�9��tp��������jb��!&P����ڃ#�c��>�ܫ�nV��������X�X�H�;�=X�<�.��<�~�^���u�k>�Q�W��H�9em}��g��E����/��4�U	��Y=����^&�ѮUBՎ�[??�->&�n>U�7�˗���m���ٞ�VV��T}��k�Mȧ+q��p���*��{ON'e���d���>����>�MZIk�w�On�⊭p��(�󨄆G��r�i��=Dx�3�t���`�x�{:Y�W꣡io9��
�}�^mF���S�סN�|���و|�n����zݜ��M�{@a�@��6~����pD�5LoB���y:���d�W�?����{o�	�0��Kdbz����N4�C���.??��:thA_�&�����K37e�^�-U�I�.��{��ܕ�Uy+����먁��ՠ���r�S����<�]O=�.d�7ܢ�tZ��N]3�D���hZ�hR�WJ���������k������P��<,h����D��c��ٗ9���U��x����6$'F�&�nVL��b�{���I.�gK~�g:�.���e��핽/�8���#3�/�AC/)}ϫk7�w:���wV��bzF�����qg*{��"q��&�lF܌q��>n��3y��U#-��N�M�׷v}�uY	�ʝ�)�*h�~_>48����p�U)J>�^�k�%+!f͐��6:�}�F��;�Δh����ԃS�%%8�P�[Ex0A������1oIJ{�}�����!+��eSFM6my<��yk�,�IJu¶BS��?_Z����[#=;ρg����,=��p�D��:ȷ�i��H��+k�l�"x���������'9Ǩ7�ϵ�������VIZ��S������kl��Ky�^���tӵ���Z���g�b��B3�gD+�g݃h�:�3^�d=�Y�hT"��X�F�fê��	�om�Ba9���w��2E�zFV��\�y�G��څn j��6F}�i
��1
�� �.�@��Q���m������'w�e�d�D!�+ڥj��Q/�?M�iiܲjg�o������)D�ݝ���md>���0Ջ�Io��
� ��C�l�d��Q�;��mU��6'_��s����p��z��p\��e����*d��̈���h�5�����W�똹e�����to(���T��*�QevyJL�vO:Wo�����vߛr��ntIЬ5}���_b��S�b澕Nas2�/���>���;H:�����ݯ&���@�.����ˋ��\���u0k�5\]���'u��mRkN��y�����j���<�ӟ����#�&"M��KJi{UG��4�}����^�=3��j��'m۾�3fB�n{�쭆�N���0�x¸:K^�Y#���Y�,ŕ{�����b��'�6R^�w#%������7�4;k�6�s]�H٩+�~��z g_K4��N�t�2��F����kk9o�`0��Һ�D/��y-�$�(b�^��{;hz��a���3�y�Ŵ����`�V��*ti2����^LpK�E���N{����'=�tm#��V@k��������K1ݟiPH!E�$-�������P����W���L��Eͻ	m� ������'a�
z��7���Zܞ��j��W�ٝ���ݞ��K�~�f�����G3G��}(k��*�A�<6�^�Co��M�ht�i��E�./ 2dJ� ��kH���d+��l˱�6�:j�<x�Y<�f��=}���3���G�1,m2��I�%�Db��b�Mɡ[��y�J�{x���iY�k����!�R�9H�˧��3CO��l>̊��/�t템�g���qo�s2���z�Y�KAJ����D�yъѦ�澃gh#�y�nl�Ă��5���B�D�hkۼ��	g��έ�!�J�ɉ3o&�M�諭���u��9��՞�^�����x��3�be̮Le%��"U���1��9dw{�V}nM�I��8ٕJw���ٞwM�j6����P:E���I:�c���Rڞ�Y���7訹���L�Z�QU��=���Hh}�M���YqI�]ٴ��!�siig�-rÛY�[��W�.�Qx��]����}#�ߖmz���˳.�R���yғj>s4~Z!�_�
&���9�`��]/3�-����Zd���F�)��a�O ��2�� ;���ǣ�Ub5@̖l�0�ѓ^���Zd�����y��8��W,��xz_�+43�6�>���3<��lzǝW>��w�jdr��W��%��xW�u�E��ɜr\���I�_7�l&O�r��N�[����ѽL���ʬO[.̭��y�T�ݬ�4��fS*%�s��vLM�g+h���x�	ؽ�I>�i�g�^��YӒ�(��������b�a,B�FG7z��]�Z]3A  v�w ʭ*U(a�\��Ǔ+2�l�Z�4;����3��]E��Wq�G�֌�F���f���6��ze�Yv��#dP� ��W+:����W��fi�Wi\�I�W]�Z�U>2H\�~O��v��wښ��֟;5��D�M���]���3F��䣨�:Zꐢ澯]�Չ�Na�]_�X)������r�o5I��RٍE:>A5�"�WzR�xb�#�9����O<��b�?P��n��U�ټ�X�#1&�(�$�x���c%b�<������~�r�j�,�n�,���f�ot��8�F('bKjk�x�Z�>�;˞�y��2Ϧեۇ�jo;g����[=�%�׬�T������67���C�^Oj�H:��ڠTy�̳EE�<j{ �8��+�)Z
s|ש~5����buݭ�P�*�ZW�j�ӳ,��t/�^1L��VE����45j/-텩=�Kj�%{��2����-8�o3���׋��s�厖z��|�k�{Z��'-YF/p��w��J��A&�Ĩ�[����r�������U�l��E�r��\�u�_r�7[�Sٻmň�D�H-d��\�ƻ�P��n�����@C}2ى>���L�G����^��v��r�ѧi��P�2i<����1cowٛ���*�$�����3���
�ҫ/��<���h��e�5�+���]ZKv�荧Ԏ܈��5��5�i�(�g�G �=F���=�:�׭{��!,>���Yu�#��ݶ����'�������W}����wl���p�½���C�"��[�K�7S;���v���%Z�.c}�18��%�MC��:f�l���ce���0H�uX���uhV3)���}�׶}h�t���-q�j꡼�D�I���-��k��uE�%m,!W��7�'����j�8x�����G��9q-y�N���:�X����&�ױmS�������>qש����;�6#�q-\M��mՊ�#1��vvɳ�(�����%?�ů�^}:�j��}��%�����CM\ɯ��~K_�H4�#�%1z��^�>��~#c��'k|�z�FO����s�´I�UA�"Վ������vn��TQϏl�gr����
}�<�#N��!5p+7�,WԯlXt�JX�nWmu)ö1W,���u� &Cp]y�D�Y�c{w���v���Un1��2�Qɼ���{�sc����R�~����c��tҳ"�^{ץVE,�+�j�Y�m[�H:��s�u*[���*�\�� {����yZ4�V}H��k�<��Z����b͖��[x��*��3{Jyg��D&z�E���Q[G�(_R����-I��Ҏ`���
�/
�Z�8�"i5퍟I}�f
��l�d�F�ω��O�u,!�*-2͛I���3@�h;�U�Q��=V��M��}�s�{����_M!S�u�M�j�m�7L�ZW�qM�Gc�j�P�N!q�۲����xHRu�'���kd�_7��bY��e6&F�1��VQ�J���w�`X[�2B����zn������S������$�U#��5��s�*yt�ύ�A���s�����g�B���\�&�v�[���)[{�U�xv!U�����-v��$.G7�ԅ��I�]ws�|�6�Ӛ�:Q4� ����\��8�.u�k�9�*�\���.��[�*��sB���J�<S�17ʶ�k<�]��e]v��l��Knɨ/r�� hAR�e8���:Zv �m�1T閬XpL&Ev��mT�U���|��LY�|7�iٵ��d��A��y�L������V�Z�Q��k�g���C�ҝ��Y�'}��[*�u{&v�e���s_�2�ux���ޯ���9�_V�8��:�'T���|3���ڇ�xY�q���v׫�d�b}���f)3�Y�T�Eζ���o��\QX�p;"�҂�Mٽ�ж�}vr}�6��1,m2�d�>j��A�>8�me�0#na�|�����U���%3�Ϳ.��x��3\�(�+�^d�E�l���S�E��5 �Q{�zE��E-��ow�n\����ޞ�m�;�S�39�q]㓢�H|o�6ͼ�r�7Y�������Z<ը��ǜ�ƙ4�Q�q+M�F�M��w�I�h2z���,9��[W�^�y��À��r��FΧ�h��Gp�0M�cf���TA����r�;<<���ٌ,��*�)�1��>B5�	<�J�Ki�j�1{,v�E��61�!�)M�Ms���O<
к�K�^����:Ft�Q֢.�9��T�K�~�霞_���(�-S֋��6p*�e>(X�ūb5f�;���.!V����r���}�B�]B����!w'4��+ƺ'lHs8eDkJ�g5\���P�\�y/V�����U_}T�/U�:���q�>��rP2pɬ	]Zd�����Ea� ��OTm4Q�K&��p���ߖ ��Y�eԳ"0�z�-i�X�[{Z�J��/�٪Ti�{~�����˶Y:�-�`��r�Ϋ3P���I%-k�eh\��,Ɯ�o�a�7���y�y$�Ƿ)^xoe�u:3<n�޷JfuX����������;����1��%���o{q9��;�W'k~�Hӥ��
.�5��5��}XUE�FS"�lށx�a���}; ��ĉ����S�A5�"�ǆɨ}��',k�3z�Z��^�Ǟ�89���9�sک<�L��iF�I�<<�6��8�������`�(��/*�1{�j�Ƿ<�����.xc���]}II�����Y=myc��-�yn��j��e��dͬ���v�����B���}E˘2�j=yh�lU��RS���:��w���v�.\�%�Rʫ�K�k�2�$��f�U݉ P˺�Y�/n������˞���挘 ��ڻV�oLnj�ź0��I˚��j��(���{DE5�q.�|��1q^o8�u_�c�f��gPɺzGJ_ ���6��C ��+��gZ[K��[�\�X��E���;3+�t��]M��g]lV�9�3�%��Y�]mpSM6S\$�"޺(�*c��.�y��`�/mL��[�LK�j�w7_���K�/\�j�$�_%�h��9�0A{�v�vQ�n��4	��Y�{�e
��M�������gh.�Ʌ�W8R�XHO�j}cB6ԡ�H{��̡bU��^r�6-�h���([���7L�+/;�뺀��;�=���,�Y��\�0CK�ݖ�	�
���\�
V(uh^�n�4�e��w��l��_%X�}k��R���R8�*�]Ze�؝mu�A�z�jy����R�����$���u�P�iV^i�ƖJ�f8��ػ�ݰ�`҄S��ע��˨�굎������!ίp���%�U���`!g;f�&4�eI'4M��q#�������V�X��_R	���w]��]$(vm���,���6˳�53��b�7�o�����1���j��ő�gg-ݑ�1[O�lN�XL���m+Ũ�NP睎L]���pR���
������)�3�"VD�}��f���9������D�./�w�`�hq�˫���v\�ۆ9C��
���kK.()[�[�.X����b�
�'H����}1�u�S.}a�
��s;\��״s�Ԛƻ������Mn\Ӟ��8�h��%��r�%	3+1ɬNfʔ.��h6��ƅh�z:�����348tYKh&�+@��n�y��E"����0��L����9ƻzѕ���c;X2	��d,����9�I'f����5Յ(qW7��Wv��'5*��4@�WňV*�^��EY�-7�M*�m��1xF�����K�{w��(H@Ũ��z���ݼ/��1�n����J\�uso��d:bo6.��z����џ	�$gB́������Q[N�m�Y|	�T��ct붅n]w=J����f��.H^�v�Z��f.�h�w�Y���`�V(.J�����eve�ѣI}�6&V.�A&v!���n�m[�b�CK4<U�HEX�]r���T�rp]�������c �:�s*�]�Ou�9�\�y��a�\�9�]6��6M��S@�ݠ.�}܍C��a8���AQ�=�뫼��f+��Ep۰�0�k���
iwN��3��Ӵ��4-�;�n�:��b
��:�
*[�Y�-���]��r�]ZX@K�α�n�/���O��ǳ9�wW@	��-�Q3cz�����ǧQ�"����"�{��G����YC�Q�c�/��r�*�oE���n��~��|�����ҴDif5����$�� ��i���Z��	��F��
���*�J��*��J(�ֱ�ET�LD��DPD1j΢b�R�UHl�#mTEMTUl�((����+cA@UD��PD�6��Q5E�DIM�UUPD�-;h�	�
�
j(�j����Z(�*��QSAU[j����8IMLU$W#UEM5LEIm�
fJ"��� ���%�(h�����"(��hj*J")h-f*
j�������PU-TAA1m�b�"�����hf(a���Z�����%�NӘ������*���UQPT��&�STP�QZq%E5F�hbJRcmCDCT��+F����kL�6h*�b(����h����6A4SED�Sm�����Jb������P�RUSMi�����J$��B�"&H)Ӥ�h���(b��K"�]������5��n��>��tj r�7O�1��傕^և��8K!U��#��YW)]���=s�}�{��aSeh�ʴ�j����Sj6�dc�Z��u|.���ڢ�f[�e�����Z�%A4�L�1��IàM��)��o��R�2�Y7�]9�]�W;KovJ�c&��מ�Ei/;R{o)9,��RY�׶2|�n��$��[0mޚ�3�2У'њ���3a'�թb���BۍZ�Y�/|�^���"o���U{,tx��zϳ��㥴�*O:L�A6A����Y`�f3��0���@,��uU�q�ƪr;�:�`7��f͑�j"p��I�ϒӈRZ��f�>�}�wA���5LQa,"8�gg�>�&'�R���Goؚ�Y��C%$�<���畘ߕ�+�-ݰ�q�l���K��c�e�ݦuIe����2#�i���Ig}8cr}���t�`��:���Zw|s^��Q,�"Ψ����@)ķƾ�yv���^;vkB���B*󀺛��hN ��������ΧQ��y���y�)�A�v��㡡M�K���I��6&V3�2�4�a�S���f�5�þ����n��)>�j=vW���s9v�*��ph��y����s��e(Q749�8���{p�(�h9rך�����-t-�Dv�`��r9:��p�U�PK3xd���06�KAWק'u(�N��lb���l9�x����,�ORlTE��]:��o�*�'k�����r{*���x�8�U�z��I�$�>K2W3��6'�g���ا�lRn]��,�����2;';)�
���U�SL�\
�#s��*�\A�?G��ջ�s�E~�xfB}�1K%�m��醺ES��Z�����������#6.���b��}��2/C�{ǽh�V�-�jOjp鉼��۾"�v"<����xO�^�F��g�
"��{-��<�*��:����]�yd�׼�>����y��]>Q���a��`��}]]R���U3mNc	k�ZZv5=�L�SϫY�2EmBW>ج����������9�3=
=�S�+键��G���w�޻�^�#X��`.���t�\��j�4�n�LJ�Ơ�<7C1t ��a��s�\qńt	��Λ�)��s��eD���lV�v7p���Ńu-�EK� ށ#�QG{{4f���`��W�_}�Uj��,lw�g!Vҙ���Zd��>���z��U��c.N�v��;�o�-�ڷ\�f=�+jB�9	WM����%^���*�N6 ��>Z���Ҵb�:f�VC���u�Nώ-�`��:�F���_4���eo{9W���i@��9��>b��"�W=�nt����w8����^�rnooN���w\���W��-�x�u�*�}7�w~cr/#Lw�5�E}�9"�c�s%�6Y2�-t�K�B����,�T�T��L��6؜��ӫb����-��%���)5-b-������P
h��э��������tъ�Z��1Y�%LK1��%$�>����))�;C�*�A{�s}ǪA=��A<���=��U'=/V��3�?W�O���w��Do'|���?S�?nr:�M�S��z�,�dR}4���*}�%Q�XCT�"ҫ	@~�=��hf�J�WYe�Dp����h�'4-r(�k�|�ˍ�o�Qg�ֈu���,�ޱR��ܙ/5���q��!�y�2�c�Y}�t5}) ��t��q�����8�7����6�n^`�L��{�gVV��/k*������%I-�U����En�����h�7<��vk�b���m��7�c�^���I�螢BߟZZ$3�Ѕ��(!�c��D\f��T�׭��G�Sf�/�2NS1��*�Ք.ZU��!S��슆?A��x����}^�y׬$�i+������^ώ�7��+j��I�Y��u��Ի��/8�m�IX�M�	]5�J�֎O�+Wx��T醴��繞3y����Z� ��=���U;.���J�mL�$*ֳĦ�[�z�Iy������*��;�2�P��6�,�U�+cu^�MKZ�[pwj����]�I�%Z��sm�k�bq�βu/K�nz�%W,4�X�9�rv�}T_�+��i�V"��B�L��b���ȘQ6u�Ҁ�^L���1��״l6�=ϳJ,��,�Qy�V��2F�^i
�%n�C4߭3�Egk�( �郅�9:㙚��~�WVlְx�`��!��9zdX���\�~��P?Y�CC.�>�ܵ����1IzF� DR��k�`�01�̒[Z�	޳�Z�3r�Q�H��\Un1�����X�P3g�o7�%�9�3�YPTc^j��������S ��zgg#e�}|����9݇�*Z7�@޺�[����7�wV*�F`�Q-�aM�B�[1�jK��Kx�I�[]�/#{����[���f9����\��ÖR���ى�u=�=�=f:�_	���}髬[���6{��:�wa�rS[�]ض�u>�0#ǻ4j�%P���f�i�At<|7��d>���E�R>��]����3]��|�����u��M.ľR���Z��ݡ���E��3�h�%彰�'�)9,�ne%zބC���^�뾸Y~�����_z�
2c5�lGY�$�ڵ,�Im�k��OI�����|қ�=�]۹�|���zϳ��XE��mI>ɉ�/��*US^ٵ�k�J�1Za���9i�2���#���͚�e����|"��]��.�eA�^��m���"����(-f�<v�}7��5��'��@Ռ�ĳ+�X$ʎ����K����hVP�t�wK�9��Oj�\--�v:���_S�W��&DgA#���`��4s����J�7�r���vVadO�1�fKNS(��ߋf�,�\���� ޗ/%���{���ι{"Y�*�M����|���Z�o�}�^���7�4�u6<�y��UL�t��t�i�%��Vc�B��ȳ8�_2A��P�9#���s��݁�{C����~�-B�.�*uE�,P�.�~���^zk)�e�0�Kی-�ܻ��q=��WD�}u �ʷ�)-��\����xߕg._`�|1��+]�N�{ {j�C��A�k-�����lB�%<JI�Sq��ʝo*�=����'����\�&��UfE�Q�m�4ĩ�L�Y"ωO�c������
���w�p��͕�E��[s�k)���Y�0��&R�#Qz�%�N ?V�׷=��K꡸�\�)d�@�{�[t��1RŧT�!o��o�Eq��={� ��Ƞ�0)��-��{+n����,ɇ(�H���h�����k�'B��+��L�'{_vCi�Gwiuwz��+��Ҝ�(]=�f)[J�q��q+�cX�}�c���2��&�wW�U�맾��+N�[�<�v��=ȵ��խ��F|���f����)���+^Er�>��)����G���)gW�.�C��Zkh��y��KS���o	�)ey��aVk(^�fCP��[S�-�5"^"�������^O�d��,Mי"��+�ج��3��餱�2.tb#Y	J
mU�����d¦4fZ�WV�+�����I�<>���{�[4]D:��y3.����jݘ<d�9*��#�֘�+�p���D�V&��U`S}�n���{������������[V��[���:���A-2!F��˚�֓ug$�f�B�ʉb����-�u=�w:o���:f�Ζ�NvM��[͕�f�)=�*�����+�
���l9�f|q�CFڳ�4�u͂h�ڝ�SF���GT�K]R\���1�FK8��Oo#7<�M׬��:gf�\��ۺ�r{s��+
g���ط�a)�~�I���5��<2\6�-2�Y%��$�ŭr��b�=;b�U�vhK�R�w*K�;�ws�Iu�[q�V9>Kp1o�V=YۉKUםb�[0 ���6Р�Ɣ�֬'?}Tɮe �,�3��t"�T��u)l��)�֩���b�>���!��I���l�0Z�S��7u�W뻌�f��0m2�fI6N�Ƿ��7�vA�:XsE���t_�e̫-�س�Y�;Z�Ω�y>��yة����=�k�t�8|��x�~�*��R\����l��ַ���3�O#��f�'�l>o�;�?m��Y�����VCݑB��=>B�i� nJ9���,��Rr�p�Qw���i�%|8�_�P�{0�v����L绊�}y+Η�g����g����cf���^��iO�� ǇH�%�ys9�D\'�d�bb[:�{Z��ImBՔ�إ{�iyH��T��[��D`^�]��c�5O�-�����&��+���]ZKm�͟H�ӆ2�ԓ�U�Kb���Pq�!�-4�	U;.g�L��+0�C�um=-�K�$����1�s4�)�-���	�}��b>���M�R=p�v]K�ɕ�L�n��E&��Л�N���.�3}���^CU��2ad�
8��M��ؚ�����U󰜻�����]�e
�dG\�
,0��v�I���e�6��J崜�7���s��O/��b�Xt����;֪��Q*z13�&�փLs-责73�i,ؚ�YZ>�$�˘�f�d�xw��e�[Xy�n���'ܺ�L�\~ڮ~��{���b��Y�*йS*'�9���iT�f	�t��YL�l��g�	7�Ԯ��>9���Q5�K]S!E�%�>T���7J-u<�=�A���V�n�?a�k58��Kܓ�
Z�9j/z�[1VCfk�+ɑ��>�כ�P�O�D{-5�����n�T��9e\�@|5�!,�9(]"'��	�U��U����xj�;O5�es��o��~���s���m��&y��K(�E�%�+��+����ݙ�+��V�D>��k�z�T��6�^S^�9skHY�j6�de��c4*l�ܰԷD���b��n��=�<�<9/^yZ1�#��]��f�>��ke�4nd���U��#a���_�td�=�sU�9��uZ/1vv�qՒ�S�H��צ�f7�q�.�{^�0Fk�+a4��ĥ����J�c��z�BLV�V�}��,�o�f���1���4[��V�\��Q����ѓf��tM�v�u�tUJN�h·��T'��<�O9e��ƻU�*.ZO��Z��б1{��Qݧk|g���3O�4&u�UXsaF�,���1�I�V��VEĜ���7M�||�6:�9{����>ڥ{����j�q�`-�Fs,qI}�g�VcP{����6⚌u���2Im)+(�l��]<S�t��D&^SF�*���q�E/T��:�Sbdn���H��1kҨ1˰G�k��he˥/��a�d��L��v`#�%]j�v�5��i/{h1�k}��"׵��� ��/xV�[�ӟ�O��!�F���vπ�կs�&u�y�^��(����p�+��\��Z���5W����C&Q7�5�c�޲�9ҽ\�'\G*���`�G�J�D潴 �UE��L,Yf�rm�t�S�g6�����5K>�08�am�}N�d]x�R��VA󶯔,VQ�~�ޞ�Om0΁�PI�=��o�k/o��T����ma��⌳�]��Z�π;;yu��fop�sjI���링��r�ƾj�[�+sy�=��*&[��]��ֽ[�ЭB
9�إ�$E 4p��)D<��m*�[)2mJ��}�V��n�o�͎ĝ���H�`�9i��s�6k3�aA��s�`�k�=[4��d!W�ypvp���z�N�34���P��X��
��#�-�C�R�EkE^̣BCK2=���c�+c���]+-i�"^٦U�k�G�I���B���3w�D��ݽ!w[(�[{>�)l�k�"��0�����EK�j���`n͌�6�oY:�J�Xo0<CˬI
��%M�هu&%���fK��dc"�˰~����
�+�f��鳍I]y�2m�@>�TJ�v�^�_ �Ճ�F�c���ފ�^^�z^�"$Z�R�;5oe���	�E��A��S�F�E�hۼ�1��V2(��p@n.F�7z�p9X��.�-�C0�!�����\V�Tc�헓2�<JS���B��ѝB#�4���)wX�&a`x[�,5Ԡ൸�}�L����\�շ�N��)gM�WwP+@����^9Zy�
C�fZ�+��Ȳ��k3�fڻ�{���A���d��ǫioQ�7uv�RY��F�R�f�=UՈv�4_a%��k�ki��n��5��K ��B
Vȥ���0��/���
�������2�)5�&ov�Pvd�.$9+�u!����g�V\zF��n�;ۥ`#��k�D��ŉQ%�-�p���=�ѵb��qu�!
ǉ%�����L��TU�N���e.�nPڀ�q#�Ȥ�xC%�%��(��M�x���6��Ye�&�]�C�Ħ,mV��{8�R�v"c���D���c��VV�j�v�c�wr̽��sw�cO��En�;�S/z��6sxR�.���������;A�� ��p`�ne��V�x���/5wUMk�
��en@.�k|3n�XYz����S{q�OJAZjr�*5|z�^h껴0;��d]ڐ��)�-��9e'�sɻ<�:��S���{���:��G����qlܢ�^�%�ʔ����!���=R��+v��.�T_;�з{�`�ى�vbt�cz�l��*	�E�r�wu�aY0*M�T���a�]��pT�㻊�%�%˧�}F�*�\��YgK��]�jGO�yD�C��+���͖ue��íuZh#�)G�{���=��F�+o����j.��/2��w֙���ǖ���[���1rE�˕��lś��T9Ĭ��lb���
<�N���x������vB'�Pb
=�/imZ�I���z��B:�+��%L�Zd��}�����R*�u٪�R���.�dw5�1�_Ӝ��U��&�t��e��%)��
"(��(���+�i��RSZAD4MP�T�D��EZP�TLM�h*���)4j�%*�6ε�I� UDUEA@M[64�$MMZ�#IKL�EG1���������I4Ek���5ATTEKDͱX���������H���KZ��(b�J���j*!"*��Zt��LR�54�Q1CT�$�Q4ST���������4UQAE1T@L�j�&�
J����T�4V�1:AA�\آ�i��**�i�9�����H���f�5��F�j!�*��(��"*b.l,�DAED�sf)�$4i���"����J!��b)�� ���
���* �b�*����h���P9!k�f�3OM#���',Q�ڗ��wh����DS�Ρ��d�K��;0j[^�M� ��R�b��^�3����)��g-��v���l��QO&�^�ԇM���)�>w��3_x�$�\;��r��v��md��4ĩ���%�L������O���EK�;���I窭�ny)�~r�YY�L,8�AfW"��;`'��F��8ɺ̋�U5 ���ԋU!+5�����R�rQ[�Xt*�*Ll=��L�ᕇ��%U[�j�Rf�Kb{�f�ί�-��O\6���=�P�1��s�s����<�2u�����7*yM��)�&�j���5���3��}�i�v�Z5��t��������V�	��q�T���Ƞ�lK��^Q�叝��7^����=��X���е^��ӲN;��6%�K-Z�	�"r�8ܖ��"f4d�>%ui��kL�J+)�V��T�o��:vv�;����S���ۛ��؝�\��{��]a��5�K��QKyZ�u+u�jI�[�a]��N�,�hcciAۻ�ؽ�t����w`��#/��nV�����ѓy�Jm���T���V�+����ks�+�����7��嗓TCXΠrI��;�< M�
T-eҫ#z�w�XK��u��Ք�Aw����vw I������Z����1�l0,���'e��Nѕ�,�)">^�7˜o'���oN�Eq�J�,C���6?�8��V�>����E�;Pjl��5uV�����uv�䐹�)BY�s��e�ǆ��r��mD:�]������S���t��-uHQsL��1�#A,�5S��/4%�����k�M��4�KAWשI��Y-��E:N����h*��:,,]@W��6�_+z���jX~�c��˹�/����mՊ�3��(�$���R��������h�S����h�ȯ�������ӽ�W��Q�y[�{K}���X��l������eY�����߲s��{�^�{}��z��z@�+�Zq6בM��)|���%��S�Ow,Cݙh���T�{w���Pr�:Dی{Mx�=g��ٓ޵�}{[?z(�BU:��ƉFgʋ~wy�����9FT�|�g\�Q���նv���>�r�fv���6� 7~���sl�g]L��������6q�!vf��!�^V�.k��բv�Dn1�ǵpr{XRU-�(�r%(v���U8s)�c�eC�ގ�g�ų�{&*�GV�XgKُ��;���6k�����D!��,��';�s�T�eG�a�Q��|�i�$�ֵ,����:듭�bb�1]�Y���l��@JƐ�rN4��kL��so|%�	��;G̎^���>�8�9W`�}��w�=c�>h�79T�U,�ET�nو�)�29V�䲽9J-*}����B云��u��8||f�Cf�\�fm�r�U�h\�����ٰ���o�M��I����W�N�[�&�V,*��̭Q
,�-���lV��f8��j�iK#<i3ۆTL,W^��e��KiDӥ���|IcRy�x�e������4����6Yų��vtL���Rt�ω��-t�d���݊Q��:ܢ����ӭ�X�m��C���'�)������[���Ǔp�����*�m���L��gk�C/��n�]r��*�vyB�v�d`�ծ:l��4Tڕpu��J��t�����)�u"WM�bkW���m�D��`qR毹hv1�	�f�b[�ww�XmغWw@W9�ɴ�ww���q�'y�����zW[O�^N��Vy�_���n.~՚/��f�]#���\G\�V1k�(�E�%���V*q>Ǟ��֗fi/�wc�����rX��v��y�R��h�mF�l��W2f�M�����m��Ѯ6�"8����z��>n�+F���}<{3��ӟCO����3 ��_X1:	b6v7%]\��z�G�i����S�Yl�i/;R{�)ö	ɫ	�DV�	r\�*���Z��KO>���q�-1���߫�z�����n����y�Og"?3:�l��j�=�v��U�ۃ�c9dBR�T�V�f�d����SϨ�WE%�����d�{����LI
����ە䧰/z	���_4;=T�B�l�1,ĥ�ؙ�LrY"��ZT�.a�;�	�Ԩbi�}��L��3a�>�ǟ5-���%V3j�v���%^�����1U݊�s׃]K��:񕕴���S�W[��>M�㎰�����Xr1�餄�}C�:����=T������}�$\�Q%j�s�&s�\�#�ݾ���r��ftR��jQ��uw�R8}Y��{!Փ\d�vdv�[w�<��Z]�ٚs|�f�ES��s�/��>�;���M��=�:��~+1�cZ�B���ؚLU�U3q����a�8��9�T�vNkܶ�N`�iS/�p }�~(�'����W{ʷ�a�mp���;c�3~�iS��z���*jǚ�m�;���ɉ�$��y
N��ʹ{c^N�?8�Y�A����<k�r�cZZ���bɸGNO�S��#5�%&�LB��g[�<��sB�O���L���b���Y>;6kĩ�6�D���UE��15K
&��(-V���c]�4�f�X��VMdڭ0��&Q*�Zp�7v#d=�h:�!\�*�-��<��^��R�h����ޜ��>a�s,�Ly7./U����͆_'�j�Y�ЩlOw,��yՙËk��V��2�w�����^��&���,%����{��<�������Tk^V~����cL�}�ѐ�7���[���"��g���)�p��e'��L�7�����{h�!f͵	@B��8P�'b|��my���iOxն�H ��Z2tT��\F�V�����ٔ��ɗ��79dg_[�v�8GcJ�7A�v*����x9��3��AQ�΋�:Ē׭���g�y��I�JYM=��J ���%��t�[WJ��|h�c�{POՁ����#�=״z��3$V����^��m��ৡ{*h�M�2�i�eÍA��L�4h�lJ��%k��;���.��3\��yks�^��mC�۾ X:�- ��ڐ������L�W�P����E��\�DR�k��ak%)49�f��)؜>j�;^2��o�T��X�'T*jֽh�}Z]Wk;`߮�x*������si�wq�6��
gj�͹39S{��wS��m�]��H�f��'G�e��Ĭ�a-��5nD�k,���4���c��>Ө�:Z�<�:�*ʮ�o�SoȲ�]gw����i3�C*'ж���:]K%��E:N����U[Jъ*��9;�Vd)����3��g5�e�F��k��۫3$f'��(A��)j����!J3�>�[�,5j��e*���e!��w�0��H�qtv��|�tc���]E��b�R=�ەh���;:�O��>��9�es�̩$���rOV��1E��Ɨ`���f�0H�8������n�P�[듷��q��G������E�>��Y�jуȪ���T���Sk�TteH9�i�t�3�q�7���>���v�X���Զ���R��i��ySI�C�Jj0��ɸ4��^��v�=���M�{�f��vc�qP���"�kB�j�-@%�15�+LF���p�x�̥��2.�z�l:��u>=�]ڻ�����gpm7�E&xLv��5i����^��9^3��┫~�^O<{x�g��C�C�i�x�!����>B5a'��Y�k�i��Iv��p�ʽ����mHCߧ�i�q�}l�|p��J��c���F8��y�7g����·��f��A�U�*��~�#������g�X�	 V^�.�e���k����9i��9L�Ҧysٰg�s3gm�D'˻3zV��M�8��؟0Kn����MW��
	�<���n��H�D���V�FV�V�����8�����5�Jh!&�9�"���pl�]��1f�8�V8&�鸞�;&ʻvn�������ĳ1�'�E1c��
N镯�k��V�����v H!�q���K��_jǖ�;�v��P>�Z<�Բ�in<ȷ���\V��qgj���W�V��S���)�D�:�XU��.YL���f�u�/'e��XUL������dLWZ	���҉�t��2]�eYXT-�B����\��{�Y�Q<%�*���v(s�mg;�k�GK�8�a�,֗�e�WqX��2[�R��ƕWg^N��;��k7'�j�˿���.���sZg����YO�lE�^+����交6�sM�-L�t�0��Q���+$�٦bT�1��){J��	M����oB�a���J�܋)�m�J��f�K.)g�L-��������v�H*������K=�3Ӗjz�tʴ�������ѩ����1M��3��u�և��ΪV����[��U[�<�v��=��V�G�r�VΗ�==���K�D�mr]Խ�K�[]Mq+�Q�}<���߷��9a��0�:���!)�:��(]������ث�,�����8�P᝵{W&�:�&��+�Z�gYR�w㾿���+�u�	s����.�y�ʷǖ=�]��H7�%C(LG_m�Wm��2��p�c��C��5��te:n�N�}�����}Jq:��ݴ�-n�̎���ӎ���ך���A���G+ͷc�ݑ[�Ev?S`I�2VRXT��b�X�-8���3��hrL}�������<��6lJ)e{#t֘�Ee���X�.m�X�g�q�s�'6
�T7���϶0��%R��Goؚ�|�E��*����
�^Y=i�O-o��}F�v��l�zms�͡�Hj�}�1>����\N���Ȃ��S*'�9�m��O �ys���M�r֡�V���\թr�w�V�Ot��uv�䕴���C�m��ώ�-.�+�2�M\�+.qR�76^�#�
Z�I�9���H��S��sA�j�vu�Kw.��-��^���|��N��$�ب�lR������l`�^o�yo�pJo���������N����'��(��>N����1C�u�m�x��F��*L0.p�8�v襔FǬV A��d�ę=��w�����=�=�wU8��P���
��fz�lk�p�׳B��	�web�&]���je�Q<��[��;k�;��bokV<˔��Q�]
|�*�.���k���gsfl�{�m��_�L��ֺ�`���gՓj���c��D���Ų��H�h�k�߱���1n������0�ݙ�E-�@6�W�N\�{�L�ɓ��@�Eб�^+!�������i~~����xh.�O\d\>]�ȕ��ǳ͌��F�H�����Z����Hg��ZBڞ��q�l�����<[*,�n�|�R&�6��1�W��l�I��N|�,�������T�=rd:k���:�l��uxT���h&115�|��%��)%�}���gmj2nz;��� �}���-v[&T4dן�kL�զY�a�<�N�s}[�:MSڧtyW`u�`��!I�� �j��ˬ2� LP��q���I^�e��E�%)S˘��l0,���N��ל;��Q˴�%��]u/���
%W��ܲ��Z����~�F�W��_����&I�/2P�S1���&���x���������U�Z�ֶ�n�w)�->��g�!:qeZv.�+�Y�yi!�U��Ϊ
*�L��;����u��-�Ik�C�Z��d��\u��bY25[���)�{)ոDq_'/�������M �"q\�W�;@�z�ql-o/	�4��\w���)>��?���aQ���!�lbZ�r�奕��K�r%ba�&v��%�B���`!�PN7t_V�T�CGm��jX�(�y���F�+�4�h-��G[7� �5I�Ѯέ�a�K��5��U�҃	���9]հ�x%D��^�
�+9ʢ�����ϐpQ��8� M��z�p�z���Z�7iA�)(YШ�*sa�os�^����]X^ޙ�i'2�,������T��vF�$e�C�S�K�4Z��`.����4l�r�Z�2�|�e���jub�08 6��E�5`n�1l�!�(��DRyf�Խ����_F�O��Wq�H/��m-<�2�V��=��t���O�w�^փ�VE�c$�[�;�u�u��a:�kB���O��γ
�*Ž����g����I!�L:r���r�x�3�9�!qgδ+p�md���G���1B��r���IӤM0n����3\Δ��7V�L��Q4�1R�e��]���i���)>X��=]�V��C
���k� �.woX�����1��$�B�u�V�3�^�`��/I��MT�T-!��H͞���	ou��]�w2��6�bP�fk��'�qc���-��8;�)�(��:��o3�v\�i�]b��Y-˶p��e.ŐN�):�΋	��U�4<W���g:�MJ󿡭��{�&m�貦͡�9��wf9�X��� �h�Y\���nu����Gnv�кb��<�ki��Ofh
�rF��@fm�r��h�Nc���P����M@�ۣ͑��k�x�����Ӯ��^Dif��aLm�Qޜ;�n\(���Q������c�v`���f'�꾳�w�j�%�\����U���ӱ���Y�ˢ�3j6+�A��k�B�`Vu�SO7�5.v����λ* x *��p��f�d��qB�����-X+���o`2_e�G1��۹�|�!����VkZ��A��VSH
=���`��U�f�L�l��px�u��a�L*M��>��ʱ�$m�4�iE�}t�xm^��뫭��kղ�m�u�+Mp�l��r������*��Ϧ�wh.ְ�V��ܤ��Q	�"��k4r��t|^��%��WU�Lb�v함dha��(��n�'�Y�VE�P�ܮ��ڼVv���A�A��ڜ�{��[�L����"W��ֺ�_J�N*��n��B֍��u�L�����]�(Qu)_F���VR��^.��r�(�S��a3Fk7ۢ.�� ���(�m%SU;f��M%�PDR�2R�E1MQD%%IEh4DDS3TG�h��QS���"-h�&i����9�ţUM4r]SDI�D�QQD�EAIQ4�TAU	0m����DRU٢f��5F*��klR�QDMU��PU%�&�RDF�j"6\l8�F���gU�"!�v�`��M%�SMQ�b(
�kk&���ؠ�A��F�җ6�(��QUQNٮZ)��jcI��*&���LE%A\ڪ�����l[%CM4�m��sY9a%�d������z/9�7�}5_!'�cj�i�&��$�(V�@ӕ��K9��u�+.�/�nE�t�%���4�_.��+���9����Ҹ��y!aB�Ƕ�]ɕ"酫��9�p;��/AJ��o׽:�gK]R\�ѳ�UX�m�˺r�ee"�z��O|�\��>��Aۉ��S�Գ%�ڊuL�kR������F+h�(
�YJ���Տ:���#�����U�v�˚�V']�''Zu��]���OƼ3>~"���yf=�Fmg��\�$�n/.���9#�q���Ujf�3�(�-2Y:�M��B{j�OY�2��-��a�d����F�+ҧ�rU��ړj7�_'��Y��S���.��3��gZ�NWs�n�ʃ- �����H�c�=��;LT�W���B�"���-�sQ�'��'9e��:���<Z�[�N��%��9^3��)�;a�zz��qS���O��Bg\��U��F%�#�{Z���Az{�w�T��{�0�Xi����ո��W��hk��S�����l�SY�˂	u���r���=W��3�v�p�j�R�ئM�(��^n�&�b�>�H�iui�CTMYѳ��k��wW"g�(�,9M"+Z)"�c��*���)�����섥Ď^�:s�1����|��ƙhg�%��2bL�+�l��r��øT�G�Ij������� �G��o4{��k�]��H�d����&bX�YLؙ�LrY���Qi49����-m�&}x��#6�N�u�2�d�R�%�[u����&�V�d)&�\�W�EN��!�X4�6q���B`������gӧްH�S���ǕhYh�l�h�J �	��V��º���zL����で"`�f�L��|�(�gK]6yǙ����^�w���Z=R���q_��3�e�ǁ� �E�j�/y4u�ԗ�ߡߒ:�����w^y���R��J�p[��c"=��-��'���d�ٻ�)��h�����U�5�ě)�RM����a�K�y�交��.YB�p�:cj���:����X�٦%NL��,�,��*m��E[��4��XP��>�7��yۜ�ծ��ڕ�R���vd`�߹�~�7�b��#O)\]!�Vv�,�z�K���Uێ��A�M����
��`��桰��pC�e�e�ї���.t�=�pt$ ��a(��q�O�>�y����B|�-
�[d��f>˛U�0��q4�/Mx�I*�5���������<���c�v�)d������+�m֜:�{��BO1=;�������=i3�|=��En���/�}S{��W�BOa&VV��nf	{��'s0�&����e��3g��Nu{��⤦��M�z��颟�u,�Ih[w���-8��a>7�4�;�m�m��1�NⓎ��di�Ғ��Vώ�3��|Ƕ��d���J�^�A�k�r=���Dߦɉ�"�Sbdn���$VW�ZM{�XNI��5Ӥ�d�~��L^о�ٱ�&ND�%]6�Goؚ�-�v��>�ٔe�����g���w�e���;��8ϧe�-�`��dk�C%eڸa�֣�HD�)nc�B���LIw�m�8��?mNr��+"�G3n�,�۔�I=ȜD��a�L�4k+L���ؒҭ���{��Zvr���1�C��:�"6b����K�=dt���k�r\�G鶒J��n���U�N�G�nJgld�s`�b*t��l���e(�J��Lc�(Ju ��(�����k4k)�{,�N��3������D�|G-]�`4{څg$���eߵ�����lҖk��N��)k��k9��0o&�usս�%^��9Pi��ܦ4��+M��u,�l��)�X�ة���Y�Efr5o����]��İ�B{�jۻ��5�0�ٳLJ��i�O�L�mNՃ.�M�R�����V*65>�='IG�Jg?9U'��^���vg*�6�zy��=u��-�-פ�KYfv�iv���ʥ;݄����Ч�=jQ*rӋ�3���w��T��������Z[��^\���C��!�.y����w+��Yy����jOjp�1Gv��YԨ-��K~hq'����+{��}�������i�۔�q^R�T̦+�����sE7F�C�9(g�ٌ,K`�r\�&�Kj��Y
:T��Y�;r�������X��ߗ��@v��]xm�&���y����n�;� 9�u�ԽX�y�b�#Û �qh�W��LK�2��rz9���=ÎֱA��)X7����.��l�u*v�LrŸ�H�����u���c��X|3�3�E)� ��y�<Ք2g��gӍw"4d�3�W^���^����4��K��/r|���8޹������N�ԅ-�'#eZk�P�7*�M�f&�8��Zc���ZP����f�irSϜ��*Ծ���;[�b4Ы�rLK�YJ��)�%�Z0���o��0}�G=~Yn��MԞq�)�.����ӛ���i�b6ή�|�!aB��L*�uU�ct�[���|�б]>�s^���5�K]S!E�2֢m�PFn�m��B₠A�8��4(j+J,�K��[1-��S8klN�R�+2�}�15gYm��!�m��!�z奣��s��[2�h�{k���U�Um�Vw�:�n>�u�;۝.�k˫��u����������}E�S��+���{H�t�ke[męx��j=��fܫ�X:�����oK�H�_T���n�z#�"�s�t��:UX=c;�p8ǿI�áY�8^�:��_�����~|���ix�w.hn�Ց\��L�.޳���FJ�S���
9٘�g4Z��e��A���;�S�]�%��hi^�w��VQ�[��3}�d��J��B�%u�q�j�2�˗I�j��`�'^��L̝�q��Ӓ�/v
m�T�jb{C[��coU0�o���M�G���A�D�F���y*V�����-�L\�z����㲝�͗�۞����1�j���5�2���Ap���['�W>�=�3)�n�Bx�;���N��*���3���U)�ָTM��L��DT�͵J����b���nL"��n��E�����:SJ�wJ��2���C�hZ�9�sw��1�'��F�ܨ�;
u��2����>���h���,��G[P��%� &܇ڇ�]��1Z�(i|��\�Ч�bí6u7q���T�W��(� h	ޟ��m�(��ܦ."{.��G>�P_�R>
~�y�ԫ�o�&·Ci�2��tNp�yp�gw������)���ۻ�b����pxs�q�\/���ף����ΤF�{[���*z�E�������̭5zj�p#�����l� x��9�����S�׵ϸ�w@�s���m�ɫ���O��b��,w�U��ZA�����X@��RT��e�9�J��M�Ǣ�Rq�tV��
G�DFk��*>���qd7�����у |o==������:�7�-b��8Њ,)2����T��(�d|�g;�5L�:��x�_G>�q�w��nw�<���,x��rͤt������J�]��u@��cݙIC�u��	A�11Pwq�r����k7;�n)�]Ӯ�]-�#�y�:B�l�[="h��ͦ<'���܃�US�Y��ۇM�͸iH���.;�9��3��y�N%� 5�D.�o-gg=%<,��4�n�'f�B�w�����[��5R)�Gp;��c%j���*��ͯ��`m��ǘ�P�h��u���=Nn�=n�`[7,S2]U��o4􊾄�i��(S6��e�e?E�����t�j��-������fB~�ܪ��*;i�-�sг�f�7D�f��͔iSN����j"�|�e����0n�i��(��s-��wy��\��z����9���O�ޢ�?,\�Xe$.
������_�+5������1���k��׿�t��a�v�PxpLp~2gR���`�R\����2�G _ T-�l��OL��aFX.�
��WS��~,�C�ls�f����b���x�n�r�BWӢT�I�Ip�˫U{����N�9&�Յ�zb4�F�qѬ���^��qM}/ð_�Gp7ԩ�P�!>Є.�y�����g�J�۹%���x��{�TS��uti@Z�{��VX�/	>���fG��TH��_u�nݺ7wu(�� |l<�݄���'�FU��7n'�1ԛS�۴�ִ��P��P����U_5K\��K�[W�r���wHx�W;嗮����ˡ�J��ۻ�Xv��G=Lt����"�њy�����y�S��:]��M�"�C�[���I<ᡝh5���4 �s�9 >0�Hś�h�fT�^^�.�{c�<��A\�xw�گ�[j��O:޳:��]M��P8O�g��=0Jts���̲"�oi���'SUD��n\�u٫��w����|��:a�e<�(��HwtbG@x��\W�-sv�^Հ�^�lT�V��U<�C��<�R]I��?\[�n�w��8� O,f�<Mܭ�������w�^�����p[�y�
Z^[)�5�+ˣ�/�/���n���&�F��=��.�n�v�s�ó3�sL�~c|ϓo1��KԨ8',����3!��#��9�y<5��݉�)�n'�x Ҫ5k��g�a�8�c�R��7�)����OiuT�ygK����ajy��4�+ZM�N����==.ɇ�k��:.�����3ώ������̬W\#��M�p��Ss��{w�К�d��W�5���@��r��C-��"�!`�����~KW��z�'�K��e��+'N§:���]�(c �J�=�}#�ӿ@}��+e��������í��S�֡�.�z��.T�{_mѰf��9�:�]�-7�Y�V�@�t�򯲚�ڔR�{J�+�]ڃ,�!H���3��*M�+���羙��-�O9�ǪXm{;/^�T\�ls�^�V'ã6���b�ܹ����e���ޘ�@h��g��ʛ�LI��cuF�o˕1&+F����zc�0e�X��n��0��3W8\�Z��c���L'�ыa���*������m(�n��ᥭ֡�{�g��Z��#�g��Z瞭�F�x���.��ؗ4��V�J|����b�5ȳ�0.�]T��Z����y�؜!���� ��&e=LA"��U<���Ӳm�{7t8�y/Ky��dNѻn�/�v]��u'��亶z��� 2�3�2ʙ�B@ߘ�SGa[�S��;=b&��[���n��El���m�t���!�[�����(,��LL�Δ�vSK�KB�Ȗô��[�o�؅�4��Oi1�D��\��g7gT>S4��L�!,Ń�3�1ʫj#�N��W+�7���Jq�9��Z�a^Zd��Ґd�{\���+��MM=U�/{2`��M�m�L�����F�G:��W�d<@\b^�Tob9�e���k�=��C��E��wL{.{�Â���蛖��Fў�w<�����>�+Ū�KZ䱜��Q�Ӡ����e�/�뮹�7��(��� �#�eo35:FT)>][�/��*�N�B!�K��v3rֻ��bV*&k[����|����Zy`4�{�y}���7ke���~�C�IΓҵ�*���X-���Țl2��R���{Y�d�C�t�/l]֪�����:�תa�813�������,�7�MfSr���dT�Jl�T�e櫩�/�bd+�w���^wG���^��-�x����2-�zzsMj�c�v��ci��vsMٛ�H]�!`����+��Zޗ~�L��)�o��t��GdE��8"E�9�����������̳r;w��_+ӳ����w
ܥM֦'�5��sI౷��m~>��\)���5�P"������A�D'-���.F=3Lt�2��e;�_+n{S'��gT�ٗM>��Au����۬J��*�Xo�.�.��pʵ�O#0�.�m�%;�R\>��I�?mX�\�n&7�,�(C9T��˲Kװ�Ɗ���a,���H��.�_�f_�f�@B��rk��y�zf��}���w\���/ί�+^���UB��#e���hF
n[ ��y�aQ�}���L��h����u�K%���|�7Eճ8���p�Bw>�����uܦ/�Z[X5ؗƧ��`�"���C�՛Y�p���GQ[!YbP�z�gb�ch&7�YYCC�#��V*�Dp�x�g^l��4.$r0����Vބ�E��W0��m�jJ�S�­#�BT�D[ˠ\��;�*Tkyp�opv^�n�����c�*'��w��A�&���pn���UH~r��X��+*��Tf����ՀZ9����I�&] _g,0k��ҕb,ȹ�Iw!���%�dqZJ�����P��[��M���%�fJv��ܴ�ゲ�s�6l������E͜Y�ݠ���坈��5om^��j�����:��ʝ����b
��Sj(�2�ͦ4V�{YQ72�p.jC_d�n��iL,�I�[�z�}���D္�\sJ�n�E��C�II�V<R�? ��Azl�� ���Z�G�μ�1�]� ���li�I�H�[/6�+�P�Fݹ[�	��M���J�R�OF��)�ؖ>/��ޫ�3m�m����-Z���^�KuJR��Y���+��P�/ Hr�m	q��̹J��W�_��1Kz~�Wzy�8���#���]́a�)c�0�Sdؐ�M��qڬ�{�$Z�n�r���nd�d�Y:�v����읚�0�s�r�ztNL��MQ���QZf������YH���A���VHtP���)Lѻ�Ƕ ^�Ri&�q3OQ{�ˍ��͗tLT���c9���{fT�nkR�p	���;z����ũ�����ZGy%j=r�.
�Crb�>��5xYx��ukEKX-Û��لf��4��8Fhy�)\�,8SWz�٦�����/u|�'n�]֎6@2]����31ݫw�����,\�.M��z�"��D�y;].�),P������nP����tn�׿��k¼����.>Y=�!u״᱿1�qꁨ�Ǹ�KP��� �
���M�}����D�f�!��iޏ$GOH�)��6�i��J��K{���&�n��>����O��A�_r�����w�2�Vΐ{�lnŮ�|���9O�^ޛ�V�&�=#m�{�K�Mn0S������*IA�{9�>ak'^gZS.��Ws��"�݁t�O`��efN�+��U�ڰ�23P-k����IX{�����{��T���B����{Π���X3����·�l���[�U$��[y��:;�Nr趄��� �!���pֵ#.�oe-����V6Ǝ6mrS_�
��mJ�aA��8�K�9��&��;՝�ǰ�oj�h��,��X��>�j�������e������N���Z;N�j,��+V�̂����Z.�m�� v��i�D֚2fh�q)C�K�rV9j��d<�j�=6�^v�vڐ+�nr���b�4/mv{��Xuj��n�V��`5��3T�˭�Zo��:3'	{����gҌ� ��w�]�>Ρ�q���C��F�U]�ݧ��\���&�I��h"���r��
-�#70��LKV�!�huD�S\�U[(����傆clSE�����RQJZ3ES0�PD�ӠqE�1MPP1�4�\�F�-f"��h))����6���M,�USBU�h)+�D4r4�TC�s������f�4�E�ڙ-ry4\�Z��41`��Ѫ�<�C\���� U �=�wh�
�%Sv�	{��[/hD����{�ڶV���(���/�����r�Գn�<��ض�b�i�}f=�Mf�!��P_�?�s�Z&�p�*SO4ڕv���?��:��M���9���9�5'MR�>��y+U4u�k�Ss�K�wm�j�ƥp�ut��oGuǳ�Ԉ�c�:�0�k��R͓�q<�+��A��X;�Kw����[���E��r��Ւ�%��*Y��IYf^v��R��^u4`�T�����:8��44��^��v[�d��M���+�-BL�4�Yg/j�U�����x���
n�w���h�(��4�"�P<}��T���Զ���w�ˌl	��sXiUs{�-�܍t�]�\u�	�wο:�w�S)Ę@k��ż�f����_&����\MَD�������+6�%m7_��T��p;�;�/��\@�c���z{�eP�O]Ka
�/M��w�c�c�v�=�Z��It����)��3��������r�{��*M�q㧪�!�a g�p��3�㪘���Jt��OչU��Tv�-�sЗ>b*�t��h���_�x�|��6~�+qLp��x���s�(J�q��v���6_���r�=F1 n�x [a'8�{�:am���Lѝ,��A�4*һ�&19���l�cK+s{z���[n�击�����%6NU����-���7�mcθ�u^:J���]p oq�*�+�[q������*����t���0&^�����.vs�#����V�.�t����szp]�1�K�eM73��1�9z��S-�٫�xݤ/���,�Q�{�t�a��\����E��@�j� �SD+#e�2�,��//z�z6Ѭ�4:v5��}έ�8CPY�t���Om�n[i��@צ���]�w�K�<ܗ�K]o,>w�#��;��E2ޚum���S_K���;���MڄQl�*&{���o\�ҺQ"$w���Z��|�>�dk�>L<���\����ҟ/:]���Qw�C�j���oK�W�؜Cm��'��1�i�t$b��KGS*W�/M	uc��+��D��y�nQ��H.�2�6��K�
����;>�ɞS�;���-'p���o�01��V�j�SOE�|��\��]:�{��)���<�2�
%��=��ȅK�z굟����
�U�k������F�3�m�^Z^[)�������vN8�{���o��(���d�r�sA��}�A�8g�����Ꮦ�����ˣ�/�/�����~'��U�z�^�&�b�U.AffnZ��[�]1���l%#\Gf�V���K�坙R�e�J�� ibu-ӫ���(�٭���N����z-k��eVt�K���S0��+gv�f��u�x�ms�:����=c����[�D�4e���dJ�ks�����C�ܔ�Ў�s�r��tP��_�UyL�6��cxK�bs�eh'�?�U!���)�G3�Q�:�-`Dռ�od�G`گ57���@'@��Ἐ�qە�e)��	�#U��.����0���v�Ϡ��^�>R��u1�f��e׏OM��%�8,�p�i�01�i���j�8Ms뎂�$L�zfa骮��ٔE���	�ɧS�}�4�j��>qn�>d2�i��?k�͙��댵b�˺���h;.�J��Dv�zy�(=0�_���J��G��+莳�ݮ��Kj��캙�v:^�ҦpSLB��������x *�@�r�$���U�c��KQ��^m��q(rH{�B~�ε�y�:F=0�/�-�Bw8�yƕ'�8���(�n��X��=<t?I�h�ǮF���Қ��#�r�#��B�~53>Ŀ+��p���<�)�\�AD�����4mU٪�C9�Iu���5270�P�N7xsc�4�n�ʪ|����Nݰ�s�_6�B��˃ۻr��99����t��חR~�jnK���'�h ȆL���F{ú*��sܤ!yX^��v�S-䐮��kE`ַ�V[CT��-G�gx%ՙ�d����e��J�������k��5i+҅6��Ɯ��:�ٱ�4k�2��4G��k��O�J�Q�R92Nw�v����;7]��]v5-�#��t��S�4Y����,u�T�OX����o:]֊�3���\�� $�	��\u������K���<6L��\3��f�~Uƚj;���+��|��vuC�OM!�!�HXd���\�W���'�!ޡ���p/v���}� ɇ^� �.���h�����M.�۪^w�^��W�eؑ�깢;��B��b^�F��s�i�����Ol;�]�P5�]'���qӢ׿N��	lg��h�"`���dt��Ț�O�̊���|H�k�oɾ���|��N��B��TËc�q�S�i�S�[I�2}QJ�fe���SW�=Bm��y�I�MH��Η~��w�քK�oeC�8���h�0ȷKKT�{K���{G;%U�w�;�&A#�VM�j+��_�oK�H���O~�ۧ�;".�9�g���'�ct���?T���zL�E��.�J���b{C_�sI���L6���D6$��oW��f���9�WB�"����S���U1r1�`��㲝�/��=������g����1�@��B`:�Lʺ�Y�f4�򝊏G�=V��,��r���z��9���pif�3�G��c,:��c�ha�[
��BN��ȩB�T���O;Kv�rS6��;��l���X-�cr%�2����7�2���gZ��˔��9�s��ݚ��qfo��9��pl���_��"\���>�i�_���?}�����Y���L�N�n8�F�`��jJ۪K���/^Ó)�p�eB�#e�4��Ӫ]�u���Fv�WcOF��/�\�Pz�(=ѹ�<�nz����/H���5F�4L�XA�K2�����0���9`�o�G6�k<p��T�_���~�����-��������(>Q� ���&�U[X;��8�ݷa�� �s�Q�)R�y�ԫ�k��9���W�i�_�sǆ�eq������9fz�����5ޟ��g䠾��J�}]%�wI{}=�H�m�|����\E;�eP�a�W��uXm��!,X;���[��.��'4�z���w*O�������y���P����D�qu�gt
��h�]U�Ҝ�:��0="�-��2�R�J/��˘UY��f�x>?6�U�l;����n����}��h���:A�օ��)=Ji~ר���#g�M2�^E<�RF�E.�.;�9��ye2�*#_D.��F��qg�M�We���9����.~���q��Ɲ����o�Z�jv�G�A}�^�'�̤|�3�Aj��X2�,^�''@�-����@��};)bmZ�w\积j�qγ7$���&�D%'r��RE�u�ͭ����\)�ڷZ�-�٫���8J��y;�g�՝�O5��+�ah��M��fB�x	����~Be�G\@���ګr�c��t��l.9��Ź�p[��O=n�Ќܲ�%�Z��OH�	�c�z��v��h��`�u�6"�x� ϙ��3>N:�Lvs*4̄��r��ʞ6�iXb��9�+�"�'9�F�#4�͝X��ȭ����+�m^6+��[�7��4��w���B����i��������ȍ�qܧ�B��rE�{d�e\���oY�W����1�/��-��P�~>�֭�m�4
�>O;���*Lg��@�ŰW).m�e�1�6�Q���B�ے)�Ҟqo�+�ՊM�&d���&~B��3�f���Q�<;s�t����ݶ嶞��<��o��t,�`3=_�o�����������T�P��]���*�_�`����*n�mɗ�zi�m'���D���O|�+!J����Ӟ�}m�������3b��׽��O�sjB�k�SZ��>U���C:��-�����P�C@XBw�pH�1��Z:�R�v1g)�����deN�yG��_�V=hsW�5�2鉌�ަ��*�m�f�KK�Z죋��F���.����vM�c[�N�\�gs�r��م�^m	"#�E.��ʒ�9k���b;��*��Y�!P굻0V3ia��0��E����"r����珜�Wۢ���'�-��3oK���񂻫��ޠp�A��τ2g��@� �7��Y�e|r='�n#����s׼���q���Fӯ�WgL>SuU'�ewtctp��}�L�!;��@�܍�7�q���s-�S-/-��u$-�E��òq�wM��t��ep��&2��y���;zſp��b�y���B�^�F�E.� p�tE�l��M穯���/ҩ/� ~f��
+͸�%����+A=���Lyu	O3�9��'�.M΃��]9ş7��[YGX�'�p/p�k�a���{�S�6L������Kkc3���i���Q�_-C��e���i����׷�a��p�2���`c^���F�h�C�d�mU̴�]�r��$������S<E�ޗ�5�4�v-��i�Ʈa��n�`̖R���@
i�5^T́��8��H��\)�)W=�)���O9�z��׳���X���0�y���;J�9��?�C���b�SM�ੈ� ���L�g�7[@����Q��T�ߏV�>�;j7[��&�-����_n��<]D_8����uaTv��$��\;����w��:��R{%�k��k
�W9��*�]�����N��dॺ5���!�yC&�ރk�5mp��M�dv�}/��f1m�VI�@rيwܟ�,��U����_�u>�m�}ۑr?��W����5����F�����^��Ō��i�*�T�����mXO�$�1
.�@���}��Z6m�!Q��Ds�8�xh�t�ȇ�[W8t*oLV�uH6� ��f���9>��d�c��bz3#sW�k�uEW��\�#K��k�~��AK�AX����X�H��I;W3��ǼM�/:]�iu'�
*��P�4 dC&xe�����L=�]��j�������`����ބ��Y�~Q���u�C�n�~�q@)e�3eF◥��>kv�V9��w�8����1.�-=��^��$X�F3.����0��=4�n�c#r��0�ǫ%Z53���g{��Ytk�u��0�Z`�]I�{\��w�{J~�@�
�?$f�4�����n��zc@�l�#��.!�c8�G>�)�n�?=m�&�.�Bd�����kW{��dE�:�Kc<��-D(L�z��l0["�>�)��çb�V�6�/�x+�m�/ي�_����G;�Z��>]u%� 6|�h��i�-��:9�6/��r�Y�Ó�[�������K봏ݎ�lY��8+����>�:]��0-34k�6��ηY�l������N������b�|o�֋��ݙ���Q$��S8v,,Zu����yw�47��3���R����Ͱ�X�ڥG�6M"(��,ܓ$��$.ye������Q22Η~��w��̄K���8�1������/r�n�h����Kڕ%��V:szzw3NF��1����{YLJ��������R��q��j{Vgff]�ҽ�X�'^��1�Mϟ)�g�"�v
m�T�~S��4o�Ʃ�p����u�=��R��?GՂ�tE���FSD'�_#T��ǯL�����/��=�L��qtWJ����"-S�����k/��-�}�����ct�er�By�������1�	;���]�%�y	�������V�gT�m�%�E�d���ɄU�!��b�T�gG�Y�k�h��5�;����;�D:}�`���΃����z������C��hD�<2ʆ��3H_h�ꮫ�y�Df�m�L�j�em���[gC��Ζ��^n�<����>q@,=WQJ]��_0���3*��S�92�^����tjB�Ji�*���,���m7a�[/x#"�XF�~:q�i&��жyq��}N9ޜ�q,㒂��F�p����Q�E���{:�3���G���*Q��=�C�Ғ����ꈜ�p��[��n9w.+����є�Yc2���y@�)�z�z���Uуc�Z�E�1���\�(ᩫf/fM���GZ����R:u�r��ѕ+�x�8�N���$�r��ʺ����7Ys��n
�!���f�\Y�j���-�	�Ɠwg'��^�4ezz��+g�I`�|!ߙ��`1v���ޢ����p��`ܽ4���-f%�c������wN���т����k�@BHvte��@h�Ӳ*B���]���,��)V^R��S͕ת���\�=��_�@WwJw�zZ8=���;�@�+c�-��Fv�mV�^��	5�LxS"�[)#]"�t�|'��9�[��N	�Q�ʢ��u=�*8�s��ŏ޳���g�&��,�{i���T��,��H��}�d&_Q����]7��<uuT@��lp���u�0pc�-�z,۲�R5����l��zDm��&*�wr�;�\N&��ɜ]d܎C�E�m/p�ן'SLvz�:�n�~ܙ������~����>��E��7n��P���<m6ucө���x����xدտ�#}��\�#�M��As�A�xܛ��w�e��=��V���ǡ�}ѝ����a�p�P�e�U�LK;��W�7B����WpsLG 6��y���*^3�{�c7T���k�?�p�����U{��I57-�~dԳ2���}j�-GF�|���Uc(�ì�r����������kB�Y�ř�rŌ��s�������j�6�V�6M]B��k]f���Y��/�y�++K��%��ѽoH|��3��4s%�F�:�}QW@P�{�S;�khuf$n��S�Y2R�u��V����v쬍Z�t�eBĝ:�VXt&�A�޽�5�mJ���yn(f]w:�f�n�R@�VޤKo�x��o���f�v��{�R@l�*��'����S;���U�OwRw��]��Β�
����V �+�����t7TR^��_Wk�91����c��V��5���pNp���F
#��x'i��YM;8.��e��@Q����CQT!�ZH����Xa;�]�,��BUm`�L��)�޻��%Zζ���s�_JI�ǻtl�����$�5��n8)w;C�C���랛]2��u���qv�E3O^h��7��]1���*״!�t�x;Q��C9�=�S�Õ�P�ec�\J5]d۫X��f�)k��ƺ����h�I�j]Hi����ņ��E����}��#�|M�*�ft<�7M��P��]�P�9��	��*ʻx�?��s[�:���׳/��D�.�4I'C�/wh���U5F���`+���&�g��^��X�n�֢��k(���D�w0��B�u*Q	V��r2^�����[h�g	�ʤ���)��V�Rb���D|I�@�;~�ꮥ%e@�Λ��:��u��OMp�]�����5i����}W K��Ķ(Sh�}���f��tT.X�j�������MOBE%��8���=]M��5D.�f��F"Q4t-��.�j��m[��5cq	�N�D�T�ޓg�O;ψC�Z��%Y�x(�b��<q蒁�#���y�١�ã�A����;���߻v�f`��~[c�9D�������G]}s^V��(���l�XO\��V�|�@ah@��ˁ\0�<�A�J�f���-to3w:����m1��b]�#�;u����!u�ϸ�R�R���h�ϣ��ԍ���$^�G �b���<��o'=x 5Npߕh�פ,���Jub������&H�`#�^/f�s��b9o�N�\�D6�h�]x�=QM��`�r騴CM�3]MV�t�6H�o-��4d�
�mϡZ��.R|Ga��.�pfޅ��={kq�;�"5���[,�3(.��Xm�CaȊ�O�.��⑩��w`Ď��k/=v���T�V]���JX���*|�	m(3%�3Du���ӥcw����sq���N�;Y�u� r�4��r�9%��{�-�V��T��y8gWh�<C�vKw�z�{\�A7�Y����v���mu�����E�
*8;�|sm�;֖�'�� �mgV�Jl�Y�U�r�� ��<SzS�+��r�`�k�N�|��uh9&�)0���^I�ncE\���f��������Z�4Jry&nVδ5�C@UTKI�CA�@j��Zt��6ɣ�%"��%��C�mˇ#�S�#���DDh4h�U�ITET5���"���(���D�h
(�9��1��A����[1̚.Y�(h
#e�ƪ�(�M:�l�la�SN�և�.N�h�PPm��
"bi����ME+F��֒��lQ%͠�mM���f4D��f��Pm�E�T�QF#N�np��@P�Q���a|(m���TAC8K��E0��B�(k�v�̽���q�E�`aǵٸǴgN�f�{�4[�K�BVKGzS�ꓓ/u�p����l���3�4s:@�ls:�<1�<;z�����M��)<l\A���,��{Flt��歀�Ds�g��꘎0�Ӫ\(�-�W���S_K���;��y� *�#�w#^:�5�S{�9�bm
d��U�l�N��B{�2^�j��B����ϯ;��;�5��ٙ�]�r{��t6��Svډ���	� 2!;����7R�Ʃ����U1Wx�Yo�#��*y~�ZU�m�'�9��|M�%�t��4��y�v}.3�Q�f�%r��v�$���-�٢��̶�i��;���s�n2���+ݝ0�^�O( �wtc���b�rM���a����3c��E)��V��DS-/-��+� �+Gp~����X�^��%����Y��U��ʦz /P\> �����я�ϰ�R���Q���-n���]cE�X���:�r�t?�~�~�q!��j�
U����忌�p6'��OH~��U!��}�ݓϱQ��{kr��tKQ�;�Eh�|\�%���G���8Xܱ���4��X�͕��M�<�;|�*���]Қ>���YΖ�y�@�p��VeCڣ��[�NuГ0X"�\��6o���9N�ur��e\T.�{����is
ۼ�P�E�R�_Ϲ�3k����˒C�@�=C��q�n���emd?w;,NX\�m%���{@
��%-2�ܥw�E���HO#����+��'��5���LS7ts��c׏O[�0�v8,�����FX
��%��b�l'���fE�B�W>�6�esߊ��-���	��~��)�٨��8-|�x��ĕ�JY�Ob�Wf�W2枝�S��r�s�)���O9�ǪXmge��x����
�dα޸��K��?,?���
İQ���s8+�r �ap����e1'��1=ʘ�ϑn2�j�WOd�N���͂� �3W�9��6�#���~1l2������8��hA�;�=����Tq�te��Be�9uo�J�ƴʇ�=Ҋ��+O�i~���h��T����X�A���y�{�S����)O�����zK��(�!���5�hdC. �zf��DFX��ꇮhi<m����?���c�y��9�p�����K�?h�7%ս@B|���C&{�\����m��QW7k�m��_��0�J��Mz��g��F�t���f)�����'�~�D�E������ko�� ��N��g�W���:"�Wi��E�t_�p{��t�5��i�������\d�6�|���v�m�K��Ȯ}������U�WM�����������2�/�����3�[#�U6�ҧX��qj�n�窝.�ՀZ�{��ԋ����tRs�}ɯ7���vXZ\������Y�6Jc���܈���z�
�Ћŏ����~�t�\S8\ݹ�E-2_m�u$�u�rK�� �������tN���Z���J�B ����>�xh�KԨ�nc�S-47d5O��T�=1�IJ�U7�u�����/�- ��Kc:��B���x�0�zD:7o�2`�k��9Ӫ�/h��|�ޠ�黍T�1�<_�|����>]ui���r�LǮ[U�yT�5�Ͻ~!��&�ƒn�o�f��d�e2�J��-ܦ�W�t���us���B%�{*K����X�6K⻙~�4z����6-���0SNGh�0�Z*�����Z/̷�ߤU�Jx��ۧ�Q�dY]Z�k�n�8𧪢�G�sLϑ���7<���wapܕ-�v���2�W�Z8Q�I�v�����V|+�!8~6�)/���b��M[8#\����k��V��[��>�C�]�qGz�#y8��tK�kq�!���c1�a�^8���q8)��w㧝2enǮ��n<n����f�è���:a!��/�;��91���8i�2�"6Y�\�"��K��]D�'E�R�J��ZW�+_L;�h@,n^�A\|�!IR�:P�0J���?� gkB�o<���%�V��Q��	���L|��8�xpP�p_SIA��ѽ�I��h����M��ջg��3��ᓜ��$���p�k�b�Eм��?��M������~�[:tn3u�?i�/Ϸ�9EѨ�K�����몈���~^�~���q���#�SmG3�T�,~�����;/:����)��%���]�*:�5�l��4��@���w�~2�L��s�Q�R�4�O`;���f·Cgf �鞬~��E��ji�JNYD��U����p�L�Ȅ�`�����R�[ut��f��/�i�0=�S�2$uu�<f�G����gSFT�R�@C}2!ߡ�[���na9���N	Ts^�{���R�W]o�щW=���}]�Φ�3�ӈ@BHvtg�Ѳ��?L��hݳ�'�(�m��7a�r�a���W*Oc�H�)���w����e��C�/
��꠷�`�aF�8?ARdT��'6[�S�e$k�S.�.:ۄ��[:�w�2�i�O#������积����S���TR��q�׵�r�w�M���=��}ʪE,��H��}|�1�������Wc�\�a�1,.9��S�L�Ӌk��۲�#7,���|�̲�7��|�y�A�PYPu�⩙�z^�+�m��^���\�e����WQ��ܢ�܂+\�i#V�"��u�;u6�Ifa8���pڳ9������[+'wQ[��O�&ΡZ�� 6V�D=�>�Ӓ=�v���`�pAv�w�q4�l�`�_(�cr��k0Y��.��Z;�?�S�7m>N?SL{z�k��������-�喾��8�+/��u�?3n��k��sб��i�k͝X��̪�,S`@fS0�=/��4�����1ۺ��+�,�%�v��l��w��5�jg�\[�=M9#{ �ʹ��8���V�jn���LN�ش�ޓ3��!pٟ'��l�A��I���aq�}�1���2�p��P�����;�
�o�lO�F�(�1�a3�69�W�t���؛����4ۭۨEWfr:��2�Nk��6iK�Z��^�� ��<�`O��1�jf����ޚul�:y�_K��u]�h)�gd�]�W++��U��o�dR�!U���^U���k�	�?�������q�E�E�.�	����[�[f�{]?ykt��ΗCi��7m����oPO���8$�Б���!��馓�l�^]��P��y���Zyzf��X�9M�/�kݒ^0Wuu7[�	ݟK�L�&�.�9���8�[�L� s�:��")oi��6^�\���u�Έ{�uU'� X�]ĺ�.����G��)���]��#r���M�/���� {_]i��(�Sv�YGf�X���C���N��Pn[��2��\/a
(�&i��	���B�+�\�́��*���hf�M�R���ڹab�y����2�4d�˗r�C�ֹ���������)�v�w�s,���岊�H[���0vN8��w��I�SY�l�a{���,�Չ��G�J:�_/~|k�pe��¼�K�e1F�B��Y��j�뻋}�g����/ u�q!�^Z�4{<�m��
7��OA�4�eh�'�?.��,��Z[r�K8ۛ7�3�Cw�P��s>qB[[c�@�/p�i�4�9X�͔��Oz�m�s��l�ŏO�yU�^ۗUK��~��	�f�����q>����2�x�M�']���o�����d|�P��牮}zm���*g��[��'�%��wdK����l�v\Ww]	��ʭO}o�8��i�� �X�����*f{@=���T����׺��1Eѕ�7k6�\_T͑�0eDu�aю��0c0�"�\&yk<���LI��c7Tj��)<*^���t�3�)eG5����e��w�p�K��KG#�FT��	��`U�:h��G-o�����8�=sЂqsFt�ݿ.�A��raG�u�z�r�M1ҚWK�����ޡ�J�D:1d�T�f5�8�Ei�]p��%V�V�
�Wi]�J��^�ĵ

�yL�΅�Qf�[}3#��2�W��А�f�V�����ė|,	5N�Ҷ:����]v����� ��W {}PAk�e����y���j�ŵJ;��W�����v�T�1��'��2�?bn�|�]=�ߧ��m��ѻj#��$7xsc����]ҚO�u��"տ�S�<k�]�gt��g4w�gK�myu'��7%ճ�% v�1|�4-�:�WX�;5tNy��҆�qp�fX!̩m4���o�C�Ηu����t�?.��]e��h�QV���',�]�P���>���z9�:@�ĺ�g�Z{��D���\�x�!�=ҥ�#/�03W���SX'@p���C��t�\S��������к��]]m����U8�w"�fq�˺�2���C�(������쇆h�KԨ�nc���V�1��N�nGl��۸�'��n*O�~Ƈ�@+�	lg�JZ%�D(�m�<+Z9O���v�\Ct��6�-��;�v'���H��]ƪ^��)�:�G���V ����/�=������F����j�!;��T�#xd�e2�^'���MH��.�4��\�{��pm(��ܦ�ͽ��]MJSk�^��|�h��R�0SNGh�0�Z*�����Z�;�����R��4�ݸ�ڿCvn~�{7�(��<����e���.+`��A�1*"�=}�©�^��H��L���ׂ��Vq�G-J��	R�'N�V�9� �ꗴ쾬��p��>��`���o�����M9QwvRo��j�>Uݚ���C]��?�˛���c�,.�|�uSsϕ�+@Ѻ�J������Q[n�� �t�]5}yG(_e[v!�fZ3���p�"��#+��O��1�L\�zi�?�a;���-
;L���Ǵ�3��l~ٝV�gT�tK�v��c�s)�@fS0�W/Bz����i֜4W5j%�y�k�'��t��g�_8�n��:�n��n#F��ݢ�� 5J� ٳSm��q�*��_6F�h�R���f_�^�Y�{�q�矍�OQ~}Qr]mD>ob�,���±Z�O�~�0�@��#e�{L��G3��Z��^���y��;/����:Ts������~�1]/\���Ƹf!;�3�T��s���*SO:����0�A���Px�Ⓦ�i.g��Y�e���n)�Ƀ�����`��q�A{j5+��t��vE;���J��Uʂ�ص3=��rԝ���nΦ��4�R��u7���}�D߹B�9·t�J��qf#p��Ʃ^���/�{\���w@�Φ�3�Ҝ	Ό� kfe�`�*�#̨gQ��I/;�R�ރ������wy):���Ɩ���6��a�[^oj�1
؋�ܣG��d�[��l�Op�*��E�t���B[��K�V%[ݏ�����X��QÏ1�{�f�{a�a��ot9�_�Ex�������5:�t������k��"�W�y̷*��a���I�wI��"�]�:�^��h�QV1��榬ŗ1�;�Fpuc�@x�b��R9�&��)<5�F�E.�.:ۄ��_����^S*/�@����A
��qJ!=xDj�ż�v�<�\.F{-���u�3B�$Ju�n܄z�=��|^�]M��=�e�vD	c���O���o�0pcק�=\��=ڶ������	���Y���49���V7��OI~9��znN��,�G�Z���|�~��a�M�ҁ{ړ��g�R�;���7
��z����Om��ޗ=8�<mgV=:������|!�0��I�v�Mm.3�}b
7q��	R�e��;��/�s���q�zx�,=4�m���st�8ƍ�آ=tg(�%#9����i��1�6�<���R���='�uKj1l�Irz�34Ŝ�13�Ng5:3�#=-�^
��o���u=6�m� 3T2�K$6n��Os����e���������x%�3 i.t��M/ܪ=��W�1Ұ���8	�
��0J1��#7�y�]܂�WA��Z�ʋ��@Mv�p�S���N�+&ZC1WsǙaT�CJ�ɟ��催2�u�ͩ�޹�\O$�5�!�]%a=@Kc3U�l�����o^-�L�XJ�py���nliF��t�Τ�0J�.wu�q���=�~tr<�os��'4�6��jP8�Bw�q�'��2^��zT-�\�(#�W�9���y�s��jn��m�.�׽��W�9�l��\�zste&}��}w��_Z�۫����c��ԴuyW^��K��|{'�9�ޗ����%�t��4��yg�-L�g-�;$3��#c��hg�
S�W���2Ȋ��4�M��߇\���u�Έ{�uU'�iq�F�`���]A�ޙ��c�;��K0��5ų����̲"����+�!lâ�wa�8᫮�֞�t7��}��ʳ�&k>�~��BH '����t��i��-�
Z^[+��m;W�Ҳ������)��.��N���$숲_	�yfJx��/-P�]�|9�k�#�����+9ݹ�{I��Y�m१.89��UR���)ts>��-�;b .��g�e�现��{%�� z9�K�^�<�Y�<�O2Sϴ��c����^�t�LW���­����\Ò��6�Y�:��T1,�b��j�(Q�2F�[��>�nVW=�S<E��~]�N�bۻf��\��y��~=kצ����IW)4��|�n��ޭ���Pǎ�&�
.�֣L�3����+�3���ͬ@s}A�9ܾ]�4���X�Z\�o��k{qْ����*�vEzy\98��ك)U���5�oFb�,Y���Ԩ��W;��r��rP�y��т�Wm\�-��d�{�Mep�����z1ʓ$a��;�uk���Q���	����N��Z�]�6�ݨ����+@�����rQ3��c���*a�v�8�G�)jˆ�)�*}���h�:g(�޺��؍��IsjnFq�}�p	�<��J+���9���p_1�+��~Տ���D;��[_���z!�WYA���H̿	���+@ml8�̉a���;�1���*����t���*n��wF��woN4	�;�B��Ǆ�'��)t�R�Z�>U�%g[g��<Q�5PS4+�r�́���.�l}����V򣀊kyw��S�|j���hm��s�CHغT��.ό�e�K��ZD��Iºm�ݮ��U>c����K�,�;�.k�'LU�\��UJ�Ȯ�ytf�w!�Ծ���9�Q�\떏u����.����_���F3����x�ױ]̥Q��d��n]!3���]�6w�0
V���U��+�]XWWt!v�횪�ٜ\�� ��#'/d���
��y����Y!���t[;�v�R����i��#v��-��J��荻�z�L1��%3[�)���U���2n��7�<�ܲ	ܲˏ����gbd�T��|�ޱP�u��w-0ľdhj�8�2᩵�m�=�`gf9'FeN� ��F#ΌeɈ<��fV,*p�]r�9Զ�.�e�|�5��u��Ye�J��I���"�R�-f�S�u�'}$�Wb�����۵l3Յ���p�@��V�R� �^��ȱ��|qk3h�@Xϋ��r�@�(�n����L�X�������ظ��&kӕ(J��:��	����-҂����3f*�v�@��߳og��z��ĝ��S!�}�M��8��u�4����RTlV�"���C��d����Sr����x>v4k����)�:�Q� o�[(�����+�C����Qs�۫�D�7�0�f��&ʹe%�W7tH��*�<k7e��#���.�Y���o��KӺ+���h�����q����8�7ϟ%��$y��c%���2j/���vػ��n��,�b��rIڣY�ڻ2#�V.hgH�t���*V�ƊZQ'�\������p]�g-���u*T%`�&܇�;�{e��Κ�D����K�B�Q�ڷ'�Q�6bݥ�O5�w�8�*����3l�&����3��y:_\߸ ����`��S��&���6�xl��1¥
��m;b|;,�А�ر.�z�3ӻ1�̝o�`ѻD�Aސ^�����v�񫢲RW���dquy�ƹT���!�+�L`pe�:-gi�mV�]������[}9��w矼����i�������o�8U�UE�&+mV1��4QEr�� ��4cQ��\�s.�"	�����l-���ŉ�Zj!��SK�Ѷ��
kl�Z���R�4U�i��ՍMQ��A�c�ƍi-�U�9�k<�ki��<��J�SA�)ʨ)ѧCBN�S��CNb��Ѧ�f���("Zm��[KM4jb�V�j��Ά���Z�rSE/�Vmcc�X"�`���k;jq�b�����5��[Dъ�F�iѵ�����y;��X��3��hĆ��CDQE&�T�c@[�Ei�֧;8��îCZ���F��R��V�шō��kk4V�G	���N��N�QDA[m�D��j-Q��b)5V1M:�G��|�����.�-�e���!��m����� n��2��0��2b+!���%�ĭ>�ɶ{6���J��z3��ɻ���_`��k�(fKmznx����`���6�*�e3=�Y��<�T���Aw�⺱��}1q+�*.�N,[��ю�ngE4� �	�}g�7(x�[K�j�M��Ks���g{��{}KJl*�1��a��L	�LzLzbz_�[��vs	�[���X*J�R�xng����ųuJCnQ�ݶ]Z�a��C�&��'�q�4�q�>;.TxԽ�v�����|�}�~6�:���st��.��o�K��Cj70���72�V_)ʍ����c�����_�̜Bw�<�T�,~���h�y�u'��亶z���Qf�砠�h�ɞ��jgs��Z�Sʖ�MBU��������rْ/z˧��=?fGj_�J���8�6Xû�D�;�:R�.	L�f������C��ifgw����n���\׽P�]S\% �b���w�gJu�y�.����K�[��[3.Xe��̬�7�q�a��IC�tfL��M^���J !>3ѧ�!R=����^�N6�ȧ���.���d�w�?I#�s�w77<�ݣ1s~���iΜ8�t�j=h#�o�x��[1f���6Y���ʈ�#��D̤��u���R�,X�����;{M_:Wep��v�E�:�\-��{o5@C�X���b��������ױ�ɪ���{�)��Oc���}h�l��KD�
��1����`�>M�"��m�z��t嬳dC�\O{6K�yA���K�S�u�p�w�O-n�ˮ���S�����;2'nw���sA��i�MfS-�{k���Ԋe�.�4����:Љ|Ҙ����h�����z�}{��r�"��}���#G��ah���ceuV��ޗ~�2�]�L5��P��9ԩ�^rx�l[t��vD^�pF��sO���ny���4[n��[����J�hg�COmԊH���(��a��w�J��F���M��p�ʈ��|��b�cצ���eݫ-�k��{)v���~�e������|�p��*i�o��՗s(�eel8�����.�'�y#/���88I�~�|�w��\>��=|�=�=��A|��ݲ^��Ɗj7u�mU���n�$�!�#�l�B����gٗ�V�;�>p=ѝP�l)�O��r���c*���}G3"�ѻ��P��Zq,F�z�H��ʣ����M��`�t?�l�n�7ip�|�u�m���z.WS��_9Z]p޼]q�:��!��eJܾT���G�&U�X�"6�ً1s��q�ڡm��X��oEos2D�m>��M��7˳^,���Q!���Ϩ��Մ��`��B��S�Zy01Vu�z�"C�ͣ궋5�d���ث%�3[����n��qD�~Z	:��~�^����O��xʮ��曒���;FgEˆ�l�X.v��rv��ve��9í�S�%0w�,!;�9��Y�%�J�ֶ)�ŀ�v��i*nz�z-R|{�H�އ����ѕ��W�!�}�;���w�39ܠr��!=4��u�W4��m�mƶ�u�z���4w*N�[<�}�Ӻvu4`���i� !$;:5��}w.C7Y{;Us�,�(��)NH��cd��a���I��;�����ю���ѬWqZjr]�(��Vܮ�D�:#�C��5O��95�*c��ש���^�<���iً��K�,]6o����F���5-��L[���8��H�'�����T���h�XIN��׮��@��d˾��|G� ѸQ�����p���U�d��*�C�:�h��2��u5��%�Hkn�i�}	�m7ue~�5�,�pȶF:َ��ҋ'š���dv]V��kzU�@��.����ة�e�.z/�m�+�ٳ\V������]~�}�3?c>Z3
oG��`A.��2}��v�pZU���ln�� 
fӰC�re�?8��U���S���>�n�x���F�B!z�������9H�d�����NM�$�W��zbIhȸ�	�#�++��M%b��J
���Wc5��	6���z����\SyS+�˭�7}t��qy����_�)��pz;z
��$[{{d�e\��5MD\���qf.7t�R�/y�2�!n����� ߟ%;����=�=�3�[Q�]�à���=x��&���g�^r��X�\�Q���������!��7�G3�l<�ön��O]�3��J���j���y�{i���+����R�6}_��5�LGj�R�B�g��M4�醧������:j;\mÐlswGp6�ʛ�ٺ'4��l�)�@�9�����0d��֗���ɞ׈9�8,k�����駚��ϯ��	�{:]�R݈E�e�H��i'��;����֟�o4���Ό������Z:�R�yp�M����{z_�vIx�]���oP8N�^1�xx�����Jn����<���@P��s,���i����l����5tc������੼}��B��O'�ȁ�]�Ɍ`�$�\3�Z�Y��5�]I�Z;�n�_혫�7n%&��J�V#���6�̦m	�y��0���^k�F>[>��KK�d�ޑ9�ǨL�Χ���Bq�B��(�ҹX�xj]�#nvZ��Q��r�&ܢmn�ĳ�e[vu,=�+�N����ǀW$uu�d��}:��y"����ٛ���I��]X%%J��+�����k���xl��)���.���4��-݂3kcr�M��yH�\{��rx�|e�y�Q�B!�1�p��3�pM]�:��ԀMw*���S�b���j�51��$R��}��!-�;bt�R�pܩ��6(���D�f���!�6��voU?3OA�5�)���~}fK���t�LW������iym�q-��kThk=5ђ1�iR��wʹ�,2���j;Gf&���++����V��	�vM:��n�}�}�P5��՘�i��u�p���8��(fKt\q�,a��rT���O9�Pr�i����W�������_Y��R*^�8���X��.#FLA�|	�Z�*nW�,�"J�2l;��9�%i�����\��K�&a��	ߑÒ���KGO�����_����S����3Qs�7w�;�j���tcPN*��ܣM�k�Pj���/���8П���<�&�5����7qёޝ�~��%�^�p���<�k��m��_ˈ�7m�qMBc�y&^�ڍ���$��g5��u�#�SmT�ʵj��^����a�-{:]���O�-�����D�:s������Q���[c6G��߱�N���,�eo�͎��k�bK7�A�_�ͤ7�R�d�t�����ʇ�f-���$gBgXwyD߫�{pv�L�ѱs�:�}��OT}�RJ�0dNS��8�b�L{1�`j�n�e7{�{[u �q�;�a��"��0�^T��i�*�z�m�K��؅�y�g���-���17��&q�����w�ӽ3�,������i�ʸ�M4wQ"��C��s�sa�k�*@����gT>tġ9��	,A��~d�\3�蹄EnI{��,u��2���«���h�K�?V� �tf^��hʞ��^Q	3Ѧ}����K�!^�c���X���ěɋ�-�����]wi��E�N��G��W�[�)h�!@���1��[�Xg\"u2k�#7�0���2!�\Na�~�EP~zn�U/LyO��9�:�
lw�]tϖ]�ب3iz��{�!��6奣���{��̦Z	�sܦ�,�w���Q]/�jg�ܘ������eC�� ˋ~�^�:2�zr�#<L-͹YLJ��$��[Ȣ�od�9q��H��R^6��n��OdEҏ9��}���ꛟ>Wӳ���fr�j���5�2���ʽ75��ɉZ�sI�̴ao����(E#�F��X�Z�#��t�qq�Ӭ�����`̿��d񺒲�u�F2��vmۛfL����8�&sN���j���#�@�a��P#�ϯ�P��W�h�e��WÇU�\����\R���m��ɃZ��sc��"Lb�޸��I֍�u�VM���':,^}�
ö�Ik�gn�;�_nuz��-��.���ݫ�u4���	:^T�:���kVE����&'�C����%��=|�:������� �Ó"[�lkc��=Y8!_ .�6P��ʧ�H�P�}�~ux;�=6t���~6��_�vZk�a�?r8�mz^��y�����b6[���iM*9�!L�U2�h���ñM��U���mያ���#�l���.���Q� ٤��ק�/yT���3�8��9��ܼ�]O�f"{�-��gCa�[�/�8�K&�dBw�s�?%���E7TC�kv_Ul��i�eO5��=�ΤF6�>�Φ����A��=@BX�w�"�]���UJ������\-���S���w|����:��ʓ������������L���}�-s�[ѻYC'{�3��_3� �ѪzD?h��9�J���LW*Ol;����n����rQԻ��7M.'��>��a@��S�)�BѓM�LxR)岼���K�K��W�턽g��񍞼�iA���D�ܽҲk�ͻ'�ntD��u�%��.�XɌ�����v��I�}��0�:*}{����;W�S�YR|��4(r��Lj��m�D�
T��Σl�wG�Q�9��B^1���y���B+޸�z�N-�Fu��wi��o y���y-���V/k����r3-Om7MK"W7U������S��{dw� �t;�&_+��L2%��}�g������M8����rq+��5-;�S�l��^�Sf��Z�o4􊾄�6��YB�v�^�����3�㬱�D�o\�ϑ��n�tK�et�7v��粧������ؗ��Z�zz5sV��y���R�Q�T���S�<�q�[�>�I����9fS=Z��O�����{�%�k��eWsʎ�ʓqr����@̡��2ƛ��L��o���}e*c��@L�RڌD�����G�|�\�>��������^���Q
Í�7��d�����c��`��:��v�:�x�� ����%\�h[�-�o4�i��es�.}jP[<B~��#��uK��M��b)��4�ުX���6<���X/�;��R݅D���SV�q��	���'y��7w5��$	��|�;,����Q�o��i�us��o7J|·Cr��Q9��ޠ �@G�(���w�iP�Rm�͏*E�rlFk�-��#�(:
�6r�r�T2��S�^Wcĩ�?CYe3����$�]�����Ǽ䒑��Q)�

��]��ۚJ��� ++M]�;b���y2W<&\:;h�zcc��s�K4lo�4�nx>Τ�ۤ�_j�]���w ��F�����T�^^�.�{=���{}�%�3wWSrww�ޣ�
��]������dCx`�t
 �7l�YL��4�w/l:��я�e�e����N��s�Χ�K�����`sR>O��'D���p�uۙdE2���LWRAd�g����J&w"��V�G0ܜqL���7����|��(u��>U5�82�B�@�������R*���̇���T�w pM��rx�|�@<���!�S���B��/s��k�8�ݮ����2���<�O12�Q=!����T��˨H\9�8�-�-�� ��{�Z��d�p����u��#z`7z5*ǹ��^̞}�&�=�.���Y��1]���i�����D8���Y)�+�U�AkX�3�7m3�`m��9��Gh�Ms��M�>���"���	��u;
7N��
�
0y�t�������W0�M��d�Ź�L3%�M�S��ap��U�l�g��WB쭟Ц�m�k�ߦ~�;B���_L�fL�Y�~���E11�gϙ��X�/ԥz��,�g�, m�>aR��F��t�1FP~6�;�u��̂�Y�����y^��׼wq�9\��}d-�Ye9���df�iL����o&j��.��9Y)��-�'�P*;���7�	�s���]V�˅-�V�(8'�s2n�C�����Ԟw8~�rx�T���#j#�,�!=�3�k����/\�T��������Z�<�=������:gPN-�T�6�m�eը5{Lh�4!=��+���Φ�U��3}5��1Dj���?~���2��˧�����d5#sW\��M�Gu��3]@��$A�z��"�j�<�V�����{l����R~�R�YL�z���L��֮+=1��zi<�@�ߌ2�	�N�a-�����_�C�j�|6]��Ye���es��޳����U����P��b`'vJ�6��i���4����g��D�W�V�;ls�Ctgt>�Ψ|��BiD8@�����̔k�p���*	��]��L[�+eLv���O�� ��׵�`������#�xC�I��>�y�L)>��Bwl̝���LK���\'Ei��E�O~Ƈ�@+n��>T��X�O��l���Uլ�ؼ"�����i�Y�"�#�5�2����)�y�e ��s������� DW�@���� @DW�����E��@@DW� �����"��E�����@@DW�@DW"� @DW��_� �)UAW��_�E��h "+�����d�Mei�k�	�~�Ad����v@������w����>�EI
�6ҭ�QAkQ
�&���k �P�&�S3B�KM�m����J���m��3E����j"��mQkf�l�-������ٛmm��[fh�wlM��y�UJR�3F�hŖf�M5���[lT �I�Si�6��5�����R�6T��_m\Y�� '�WfP�h^��9� �5�Z��(������ݎ�Pt�Υ)��  �(�"���`5  �up   �   ;]�  ��  #vҍ���6�B��e��ζ��  ��ٸڲm�;jӡ�t��ܝ�t��F�
�t깚l���fѳm����l�  �Ŋos��i�i��
�\�uJ���9��;�U�T�n��J�;�AU+rV�d�[QZH/  �u��5�n�l�7Ct�lm�t��%m�wj[��F�ZiGq�)T�tΥv�h�--�R;n�U����QE��o ^�j��N������Um���ӧY����wVګv�)ۦ�ɥ*m��U:j�v;��.Ң�1k6�F� /x����6T�֛V������ht�l�U�n�d��em���M�4�t�v��\�iB��+l2�m�-���޶�^҅,�(ԙ[jG.��4t�W֢�2���ѝ��+V��뫝8��k�\�
ٚ�w9A���n� ����`�c9��I�Ymj�����k�γWX��t��4LP7q� ڭ��c��5���H;�
(  
  ���U)IF��h422d�1���)�  �   ����T�#LLC@��M2dh T� J��4�T  ��`�"h�M	����4�5�Q�M�d�M(�I LM=O@C��?_�����_���Ջ�.�f����j��}��0,�܉	"��Ŝ�$�u?*KH2H� ��$�\��4�*Լ�IđYl���)���_������JH�TRH�$�����5�$�!�!�0���%`�@�3�t����`dS��n]�o��I!��&�.Z_;ܿ��ZQ��F�Y/:�ҞE9���<�(R�"���z�3����?���������F�,h"˼j`��VH��٧%M�,�v��Sp�WZ"�V�9��FK��;� ඌ�����"�"]��X� �&*S��VhMxƉ�,�1�%���ip�e*�&fWЍ�kzҐD�'cA1�ݚ��ۺ4ݻ#^#N�B�\b�I�R�� �4��Fq�T��l��UH�Mˎ4Q��I0�2,@�A�V��Lʺ��ib2c1���j֎W�@��6�X|�XF����+�������ˬ$ͣ��n�o�-��r*���Gr��n�j�]he�q\�� ��V8h�)\ݦ�pڒ����̛����/&�M�06�ͷ�r�ϓ!AwF�P���46�l��iûLOE�3JT�d�R3�F�c�qMtJ�����L�Eaƍ�߭=������.9V/wtF W���r�+�\�*f�͈+D#��O~DQ�6�q2a��q��9Cm�cq}Z�f�DޓB�̺(	%*��V�fڊ�Rƪ��`��-���u�V(�p֢�M2��Sɏ*��Ǜ&6ffX�Sp?� bx(�-�\%J65��ݲ�Q���r�F�N�A���P �i0�l{�IaD�)�an�M3*��c ����n���ɫIZ���^��U�0����2��G��r��T�v�4Z�14*^&�ܢ�u��;��Ue*t������65b��"���V��%������e�i����r<T��%j��2��ó�ִ���D�Llwo�qV��$Uh�
�{V��2��ID6�3���n#��x�2Q�R��:�UU��)��,v�^��j��3q\YZ&0�?�{�*�c�J�����w�i�'X�;6MۧM�:��b�KC"V���H�9R��pX�&aϣ��J4n�D2�B�[���$=n9�BHe��j�h(�G\�	@I�*�e�g8�����10�h��/l� ��E�ѫH��v�$��cjeb�Yճ05a7(%��2��R�#����2�估ýl��Y�XI�,SG)Rb�h�Vp�wukL�N��p4���1�I�A�t��@�Yk)�ѣL�\**Lm-E9aX���<�cbh��ʯ�U�_H�R�&mxT���f2�S�okBP�".�X�Ye���w�C����p�gk-3��R%���UY�.���.�(��$�t+\V��[�7[���%�Q��fªn�i�m�g���Z7��j���Q��3)�f슺:X�Ø4�d9�Y��Q�iM�pe�2'h,�:%wG@�w��i����Z�t�NZ6h}i�o76�ch�x�t�kU���#iѨ����@(��ll*��l��-�Uvȫڲ��I�
���A����?P�,*�A?�o�\n)N�������:��+-��6U�D�H�_v?�kU��n��±�«aB�5T/p*�p�6�����;[P�v���Hu0m�Ʊ���uh��"�f
hU�kh\GF�co~�q�����Yuf�3%܋a)���*�ϝ�L��#�.�M���]A��k(e%��I������yy1᪺�3-�k�o.L��Uc���$Ӣ:��n��d:��'�]�8'ԎGq]S�h1'����of�N��r|��!�	Zj�w/\�&lR�&��ۗ�2ּ�J04��(!��8��k����lǪ���!�A0��n�ǔ{�K�m'.֍��̫|aثaLC3�m��� jn�af����:Txhe�������os��, �G2���M�Fxu̻'uO���!w�1ٲ�1[�)�`uYX�V�5������Rذ����L)o����4K�W�����J����³,�ݽ5%m�Qfb��E��n7���:���t��ܸ�S��d�j���i�F�5���ʳ���&lrP�@f�4e��8�PtZG��9Pd8n�B�.�Q)��H,ݫ�ag1�6]K�!����A���l �Ӿ�x�g�XJ�q��K��p���h�oe^*��zof��+#�(\#�oA��������A[�B)X�c.]��s[*�
&*�r��F�)�&j34��7J��Zt���=����/*ni	B��$�	�o�ڢ2�y[��B�Ԣ����S#����VbbQj�~���M��Ԁb2���b�T��in�6ɼZ�H�U�����UM�c�1;vZ�7K4����;Y�Td�0nÒb�V�G,jLYH�f�� ��A�y�+f��"�V%��F��v����R����U���B��D��ϳm��j��y�I�MK;�L�1U���y�Z͎��B=QO�����	�'�e�@�72���^�	�۟�J� �{��^J�zoe;v⽗w�D� ��[(����w[T��~�.JyOeu+e��nhj��V](��A��i#sI�2B1��2fVYҝy�H*&�+�h�;X�J�U�7k�`֜̔���P���ʘ�����Fa�E�� ���E�i�R��kl��nޢo)��V4��yN����;���x�6f���n,ݚ-�+4��`�MTe3QHmP��A���]�	hp];��RZ���ѡ���/}u�G�Iʃ]PPkt�x���{��q���*F�{4�z�*o�bNGx�{�ksfh�E:���w��(��6��W��O.54.+����a^��Y�r���J�ua�r��mm�Ù1i��	�k�$�pA$Fʡ3�7�m�n��2����/���q�B3Y�I��w���{�I`q-��8b�*h�	�FmV�$Sۡ{�.����I��5����B,Bf݅���!�K�J�غ5�!OU�5Uy��o��HV�4�c����y�[���i�cb�%+;�E���2����nd�h���U�j��j��y�����ZM;��PˢAiē$�V�{�֖^�3�`]�@^����GU��$([r�*wd�GZ�w�7�����gY+��*�5.�n,J�L��f�����J�9��,�
y��*��Ǹ���kl��K���&8�4w1ˋ㛣0���Q�E�ibl4�`�ZM��$3�#v�|ur5y�*�՘�pі�bE��-$����{M��.�EYkq�����R�'ue��IE�܆��T��$U*����xt)���1�J�ݼe*ͽ�15��S6�C�-�6�̴�(!/Rwk)�k�]g��+Kekw�Y�v��v�U�ęwhm֗C���,��L���tjF����#iú$�,N}�����vS���2� ��ji�ц-L�ܥ�0KR�Wd`�M �mޣ�4@?Z�%�H��,b*�Sr��U�m���;2�"��VN��+�u5��UXE-�n����eSXYT�{V�~L[�)����ws��~^|�e>����@ƅm,���b\9,ū��qe5�r#���
4��n�aAk���h�W�h�.M9���2���*�f��Z��d������[���,%�z��%?����k��ѡkl�$�x�j�6�,U���V��*�O�ǥ喵�+v�v5��g��B�(呶���:�3��,�Ȉ'/V-�`����E��)�yY����F��vBu�|	��섐f� R�#�[lV�j���l���L`ݛ*V5�̽��-�j%��*h�
���$�{�v����X �̀5ai���JU�&���ʠo������ӎ�UV�/�s�����:آ]W�/�*�0�� �P]�����Ǵ�`iz�8�����#m�k�ٛz�X�W��xq����`Ѭ�(���Q�+qgUlx�X+�F+[�
E�M�:M�Lr�����R��:�Zu��m�r�aO�&M=͓F�*]��|�̤����ݢ�*��b��I�՗{�Zl���!Pa��n<Fn�@)H�vc�tժ�.-��ٗ	l=�a��RM�j���C1��^��ЀP?8�Kgpla�J����LQ���#+��:�كml`�`*�v�` qQ{qB	�Z�eC%MB�u���i��
;�@��x�[�r�Õ{T�V�-�ٚѦ�5����#z�^�wuCNl�SQa^�鬩���e�{p�U��v*��6��r2�gn���ڴ�ݔi��O4rT��<Wc�6լ�y��;8�V9@�EYDd�W0���&�t�˻�����|˦H�E��Д/5�&�s[Z$*ΌZ�C��Ƽq�w�?���R��9DΟ�Ʊ)�T�죡�}�eR�4���U�L8tq��-mѹ%���9YN��}-�P.]�펮lX� DDK���Tp��E�+:����SY^� �KLC�VZ�o*p=o%NxӨ��C�O��Ad`�j�W}4�9�F�tcv��}XM\�����`�E�J�sJl޺ܮ�Y�n�nN��%cY��fW\�?N�*�h�<"��d�61����R^���dy����0V��l���{�l���F��銂��+)��tg:^cU�pC�oV,�;�0-��I�t��E\�|��YV������@�2�Ү����b۳��]]Y��S�nPp/M�����gS�M�21����|k/!7~��B��\;A�������OQA1Q�U���m "�G#�)ϚUٺr�kY��ټ��ܘ�׸F��ծ5,����@G"���.�9�R��s�@%�c����+n�k&ҷ�lY��W�a8��GP�0�n-�Y�z��K���)�}��[�jD.0���5Y�����xm�&V�s=5K�R��5���u��B]�����/��K�]V�yD_"F7�s��s�DjO\3㡐�!��D�{ck��i�4�q!sL{�N�9�WT��Aǥ��X�YS��4�ۃ,�3VP͏%�.�v�̶,�5�^�A=u�ө����2G.FJ��{��h��w;��Yi,���>PM��]5�K�t�Dus.��d���`�R��s�r�vk��b�� �P����uB�Ī;J�aQ�T��Ȱ!n5�d�QՆ��Mp�r�4�Ҿ�}ә��V:�ð �Yݬ2ں!t}L身Ba3y޷�<���LT��d�ٱ}��FawfN�H5����^�ˮ�&XxP��	.>	�8�]G��̗�EJCW�Y�`���j�t�uXu��x'gX���3��$�%.����͢�S�[��u�җ'��Vomъ�k;���Pc3��{&[<��c��W��ɧ�@r9ʏ=��N�e�8�mF��G��\��F����M���h������p��-�.���!���$4+j;P	��pN��ټp+�Q{������U�Hewr�d��1L��ì���B�<��ۮ�A���K�q��++h���$m���'�gq�Y�)F�������� b�v�&�o:��ǟ,���:�����1��D鸲���t76Y��9�E�[Wv҆�ɛ��'0R���/��Jಶ6}X^b�,�e�efr����.���y+X���<�Ap.u�3͎�*�d����n!ׄ���
�N��YL�U�{A`,_T��C�����GTN�@r	u[�5����NS)���K�oPy�h�v5���	�� �@%���8�)sYS�[Lm\�� ��n��G$�z�vr��B�s�+��GM�[��+mG7;�ݰ�A|jۮ��vQ&�{b��!��AƟ	8$%���K�y���GFY�Y���������,m��S��o] �a�t�	��1�Ik�.�YI$��O9]�����v`�c��K6�Z�k&$!/i�������;���JY�"����d�k��\��!Eb��Ӷ���65yKz��g.��(U��;��+5�{v��74��3[C����*�<�2��&��:2tw�]7)L̵���-�d�j�7�e��2�j1�4��즆�����k-q�~d�9���v��Ev5�G�����&vmM(V�oO��X����㠳��_m�w>�&d�����Y���N�/�cj�Z���k�,��%Jz閦��!}��7��P��6�_P�g6�j�l鑄�R�}��|����|y-I%\5�R�ܭ�a엍�Xx�s$LV���{��λ�"ԏ	i����;&�`X�E*q���{g��Z9|�E�Dl+Bʇ�_n�u�%\Ȳ���������ۖ,]��g@�]�������f�wG˷f�;���ʵ}����;�:��8����j���;���1���I{w�(v��0�(�v/0q�֛y/�LNT������*X|Z�[ӈ��Rknv�_r��������ʯ1��E�V*�w�s�k�qR�7/5�i+{��	2«T�84e�Ş�(�l�Vj��D�o�G?�H�*W�V�6����Ӂ��2��K��J�'��˲���%M�v�!�v=Z%81���F6d둟���ِC���<��פ+���\,B�)�����UբܚK�[�o��˴k�vP&��R��k^Z���Ǘ�!?��� n��L���5͔n�*�;AL�B���H�ޖ}�oX����Uywla=���`��ټ�=r�[���L�c�	cn���֌�*�u�g.4��5�ٕ��e�foh�/�W��LQ�1�~��\�]gvPU�q�"�ɏ���
:k79�"s(��i�3�\�t�a�5�FCM��a�W�k6	�����r$�^� ���m\����r�J����7]��*L�/d��#����M�c*���	�pG�V��4ӏc�S�u�{����+V���1��0�4�ʶ7{'�4;��i�E�1��_T�$���sz���������."�S�AuޞV�\,�{�-�Л�iTT(uK��L��������`|&��b�8]�_Y�l�JfN-y'Yω���\ ����T�J׊�,�}v�����e,L5������� ( �{:0��4i�x�d�q��kg
ٹ��Y��Ӭs���T�5�TT�Na>��s��eer�G�nuuv��_U�l���g\{՛wpb&�7	rk\e����Ș�v��VƖ1RS�ۃK����K%f���]*�o^��k�o�0�x1PTj�JNn!c�dih/(���~bd��x�ͫ��;ȥB��Jj+�n�.L��-��XIs�q�w��Yũ˲\�+=�F��%)��0�z\�*��u0��&Y��J�`!VG�.�C1rH?�Cݝ��3/�:�_jg ��c�)�MB��Ѭ�4�1�ڽ�ﶚc�HV
��r�(He�ػ]j�2h]����7�=�	����{��P�i$�[칓��ol������%���=F�{w�>���)�Ã����F�CuT�HSj.�HR�t�v_V�M�xo�@+c\��P�9��S�)uN�y��Qm[�ޜ�Em^^VF��{H��3m�S3;m�(s�Ko���v���崍�w�q�ն�j��y(��TG2k ;\�C'6�fnb;a)�������%���sz�3�E-�#�٣s��,�T|j�(Fd�JB|0S{��{I����`�A��g=��Yu+q��>�u%��\\w�bJ���,��亠w���)uWr�`�˩ȃ'c��<S�x�K5�N�楥T]�Ai��C9�	.�x�����q+��ٵ4��1ۥ�_��`�Rui(�%ol���͓1��M��%�.�k��,V逝���b���H;ⲷ���2N�&��8m�����\�wbC\����2���:W^\=p��=���p�N�8�,Y���8��"S/�Q����� ��wU�i_!��ʒ�6��ga��5�W(�>'�	����s�eg3q�-f�ìY�¡A�3,����Ki쮂�����,���Xǭf'�L���G��L������\��͉bY[=����Y�������AX_?�l#�31��Y�8�vH�cUZ��,�3ɋ]P�����{��6')ś��Ȼ?`����;�x:<��Lv
�D�:j��j�d�Ek���*��Κ��H���c�����oF7%��ϛ�R�Q ���DW*�sH��w�Km��m��m��m��m��m�ܒI$����ۈ�p���1>�Y����X�!,���<XmG�L�,��0�/1>l$p���Fǟ0z�K��ϲ��碭
���,��4��:I���9E�⦾M�N᣺�bvX�EG��G02���=�TS|F�������+݉���O#�Ys-c�(�U��bݧ#��=T��y��6�YNOeKTN`��$;���Y��@�a��P�Ml!��	n��F��j��m��rXG�n�Ǯ��(m���x�a��Kj��u��8��ç���j�B��*�Y{���O9��J��yw�GM�Ȝ�*�qd��T��p��{�3 ���SRO��X&���z%L�ŗ�;4���)�NY�EF�����w$��,�5<��ʘ��]:�I��cgv;u���<oX9�m��	's���ػ'v�u�	j
_�)�y�)���΍�����젱V�?��W��_��~������S/r �!}�L�}y`��"v#^��Z�z2@�!�x*km�Z���"�eU����G��e�ڑ~�r��'e3��9�����	�Q��E�JHlxte�`h�g��w�F��]>�HTL�� ԣC���6﷟Vγ-7�RF+�R�'�����̅K��wq�{c;^ܔ�3h��]
sfm�
�������D�	�ӥQ{�,��p++�"^����8��q�
�eU�����6����mE��Zgȡ4#�{�v�`/*�
��ΰ�.�D »*K�/�&9�i�E�A�V7�>,e��r����dU]0�C�i��m,ܚ�V��~�����]"�9F�XVfC�a2ͪ��D���V�՝��fTe���^�����ʒ�6� ���&Wg�m��e��,-��b��,���ѣDU�֔\M趞������f|ީ�>jWn�ڸ��"è���ې�݄�i}�M���T �e�Z�]������{����K�R�Q����8�1�1K6N4eT���ǉ��>��Q*�����P�䶍�����k�[��ż���dЭ�Hm7�[�K.׆Q�9�:�N��K�^u`7{+QͺJD^��e�����E�qb.�M�3�W)��B��1����<t2�Z	�����t��:̣�V��\���b�-FS77k�Ws6�*Y�T,���K��������5޺TM��j��I�W��L�_e-|d��o롴C�N`��Q
��$=����D���:�e!�є"$�(ko��u۫�蜝�h�^�<tkͮx�ܻH�t�H�y�,#D�Њ�t�Bi-�$�<)ǅ�U]��N��^4��<�()4ik��9��y]B�����U.q<��W�@������\y��K�C��Ӷ\�E�p ���[�c���]_�r�I�D�	W�L������h�^u�a���}�kR�Ն<����3�f�p��QSV�!5a����C��	�sB����X�V`'I,U��hA+`$7-�\G�5�%sHf�k�3筟�,D�z��IM+,pK��M��<em�����I�lY0>]!�{�up�X�qX��;�M�uhΗ7�YL��wWu(r1��7j�J�LIZθ�0����*����zq�'&�K�;	�,I��w�疭��]w��3q�lϱ^_*�l��f���XRא�gmf���ܗEV��PiCq�����ro�a;6�i�ڑtDWT�"��V1��y|����U�S��/�,����(R0��D^�+�O�X��IdC{w���]k��]�B�$���i�m�6����%[�*��;]��'d���R3T�L[��i�$S�����5ލ����üh�K��|�%��p�Aݬf+�]�4��X�.�1��|V�eЄ.}�@9Eʬ�y0v�j�*�̽�v$�X]�J��fgB�� I����j����bs���A�!.Ë�[�����F�����f
&�YӪ�evE?�ٽ����`h��$�ͽ ��2ڹ@�Ŋ]�0��P������p�e|ƁK��B��y����۸�j�	HY���]�>�U���Lh�r�D���ޒ�`ܤ�g�a��ɑR`�wwL�,���Y�YlP�����sq�׆`�Ӫ�)��T��`��Њja|`�f��p�� ���mf7���Lzv��i�0�t�6�c��Q
R��4�n�wԶC���m��e,S� �ފGH�ar�[0����ʆ��Y&&��I�	�5ӨWVe❵�C0.kW8-,���	ܧ��fk�xT�(^���0ٸ�mu6��F��TL�8�1mv�`��ō�B�W��|G�`�عK�q뤖�X�{(2�R��j���r�;@��);n�6�q�E�A�M��	��-��4�<,�VSIf �+�+,;�ٹ�7:M�CP��f�� �ʸ���d�Xu��<��3���C`۪�'�c�4v[W�ٽ	杴VB�AV�ӋP�l%�s�:��o2�q$�pcKXLeu��\4��w��F���sXP����-UH�k�]�VU<��XC�d˼r�k�/��Lj���A;�ޤ��%�v��I
��� h9�E1���W�f"��ud�.$X�+�4+���J"�iGOC���sY���1M��-�P�޲�
u�O*���t
F�d�i�E����3P=n�O��!��I(bN+��}V�r�57w0\�V(�T�C����l`��[��o�fq����U�7�͏/�5{�u3F���E��0�������I��Ժ��y�ۋ&f�ð:HQ��c���z2�*���W
x��n��.�٦-=�6ƃ�з4����m�V��ڦGuJ�ʙJ��+����H�ڮZOR�ԇtw�;D�pϲ�a��Z�ûC�4�V[\ˌQ��E؜����v���mc�����7eV����I(�jcv��@�i���\:�}@���}��2��!i&��Ueb�SQ��e��f��ӽZa�ѹ��{`����ZJҗ>�cѲ+Ϙ�Fj8�s����Q�NJ�/�_@�rw'p�Κ�g,|Wp�+2ÙKh��J\B��,Qi����	L��@��e�ɣ2�t]-��9��#�+�m���� �Y+�YY�OwǔR�D���[�ur��-gE�`�v��ĭ<��<+��H�4d�*���JҞXU�![HQj5���޺�o��g�^<x�p3x4�{�!H�(��उ�i��c�f�)��8	�5d�^0/s0ʄ�A��78lڡ�6�I^C8I2�<0���i	��������.j�c�o�Ea�>�Zmĵ:��F�r�"���kKT������ŷ�����WC��򝾱�b����{&@��s�����&�iKn����d�2�b>q�da�O,�o1FWr��R�m%�����bir��I� &Q��\q����6.�b���I��')�P�Ļb2�v��f]2�X3��''����&h��+���vZ.���	�L\'`�A�op��-;���%O5\�2D��Ԣ�*�`�+���ӎ[�yY �W��vd�b�����'}U��·[����V�N�p˷8��%t�.a�/x�D��N�-QƍV������Q^�{B���mt��������u>:��>[��t�`{�j�h
:4~���t�X�C�ְAN���ď`:h�f��l��K��$@Z�4��ޝȡ�N3����^��unɮ凛�w���z=q���ij-Z&�]�Z5�v:h���rN�U�1J]2�����S��If ,�@��0S��fw#j�yR�Xɽ��ׇ��Z��.���=�k�n��D�Ǵ�sX�;g�'Σ�Kշ��~.c�+xh���*7��p.����^��t�KD�A�]��p���j<��n���wvim��Q�E�Q���J���!�n��w}����^[�Iݒ�]�Z�����(�$3,��"��v�}�AE����e��n�0.�3$�n(���b<�h�H1/^�mn�i��4�|q�X�Th7�>$fk�c��{)�FSN�N�|�<�R�xb�N��k!�R��-AI�:�8\x*^(�@�^�����m�Xq��̫X�si���zu�ЕJ��o�WFrPre���awW����S���bY��ۤ!��Gu)�WϮ[�I�}.i��oL̢�9l'm|4��\�}�����%�#��nU���';|�^�5\��n�i���yMfiڷ��X���K���]��)��y��rc_uk@��&G32���P�Wi�X�<-%�V�}{��_=-����aŖ�>��Z��9�a�a�����9ːX8�$���J���/���p̙��%��b���Y�i��pis���8�U�
�|�;�B�uR��5���e
�t哛�.0)O���=�7��c*�s����bʺ���L�ȵ:s�>��ݙ���b΀�6�E�8�[P����?i;H�6s�� ���@�r��-&��{�e9 ���\)�A=���m�&�6�VD��E��T�:λn*C^�XőS܍�@:��$w0e�DR=�W��s7�:Ei�l�/��p����ުӪ��ۻ����y��Ro1�6�����e�?�
��"�W/a�{qfk�&�ә>���aJ�,�n
L�Ѫ�����/�����Z`��d��+��ݵ+�;�|+��D��:���l���]��c���>*��6"-7b�XM�ݳ�sy�j@&��_���}�}����� ���`~$)<�0C�0AW�Ղד�&�S˸U-_�Xܚ ��2��{k��dhEh����k�p
륊2�o�T����T�R�v�a�e�[G�9��='�wP���ݺ	f�G{S兝C;8�%p��]�*�wg2v����w�ާ�0���eu�ѹ���8ֻ9t͒FPN���AJ���V��eä�������yg��W}��9,j�s9�V�=f�u���W�x0��^ C��U�E�Q�uܸ4p�ve�3+��(���6 �7�{z�΋fP!ʾ��Ᏺ8��d��=���%�oNze�q�K#�aq{�nv�;�qI���(�}�]ۚ5y��b�:E�9�p��{�d���W�W����-�9&?ty���r��Q�9(�R�j��L�q&��"�$��,���WAˢ�P����Fum�k��9q������\{��;���qg�_��"�b�X#UUAJ�R1(�AD`�YhږĵTTQPy|&|1qcEF��m��m�X�Ŷ�U)A�
���Ԫ��.j4�V��Z3�qk
"Ų���*T�Ҩ*x[�����7
�qL+���VV���*�ƶm�B��iD*Q��Ҫ����b�(�-AA�kj�-n.yn+KJUkR��JQ��Z��m����F�Q�☭��V�Z6ҵTT�bZ�Q��)*�ѵj�p��eTiE�֔Rg[B�XV��6����l��[���]�M�݇^�u~|ߎ����l]���@�#޹cMjs)�㭧}BN�*Jk���������`�[�����lj�v��۔,�<f� ��
���LY����������Tl���Kn���z.���OmzS��/H6�{K�tٞ��0�x\�s�^�9�� =�A�3�Z�*3&f��K�G�Oz��pBƭ5���T�^�.=��&[�Ş��?�����v���Y�`�E�Ok�Q�d����OX�
Z�p�ݦW��㊬Iж�z�uw�Y�);�m=�{��dΞ�_�u+U���s�G7�NS��������s�߶���]|u?Z��]9k�W�Eҽj�+6�F��i�b�i>�+��ꋑ��Y��c�J�H���r4_%#ڔ�(�X�Њ�P(Ғ	��'s��/��Z���g��H���㼢Pe����mX�tJ�u���Nk#�[�R��ڞw�U�R{��]�\H]8$z�b�)�9��Z֫7c�h7C<+n�x����wz�`|��w���"�UoCP����ϧq�q����>R�s�D [wŮ���?�i=�m�b/7i�g$/����3.��ng܆��cŝ~Ӄ�X�{��pk�<�LT�G&�Wq���BՌ�iǺ�^������z.��x�=�_�y�Tt���V�6��0��Y�Y�Iň�:9J���r�-*�;#2;|��f8�m����d��&���"�l��M�7��C2�+o�jB�+;�� �d���RW,���'����U��L@��&��~+w}���j1�7%���>ɳ�6��%�RV'
m%������؞kO	y��?@�����4�+ڽ 3sv������>�ܦn{�]�Y3��sº��	���	�ivnS���eoR$:I��{�XT�a-S�=k(�i8�>�z9Bt��.N�yy�>-m�W��*W�"lj���z�g�O{R�|�'~[ԧ�P�z���>��,�Z�]Ԍ#w��H��In�\`%��8������r�PMc�ڭo�5J^hx�X²Ⱥ��+cdeO�8�������As����{�b�L�a�!������Ψ�l򺸎��)����
���V��H�Bdr����N_YQhs7�>�ٔF�;�>�⟥�}m�⊮B���J^b����2&.���ݫ!-*�q&sL�g�1����Nx�·�A��l����:�a����y.d�<��~�D{L��<�_l�����B~�1`��{].�#�&8I�&�M���R���Y�\܍��q�X�$~\�����mo���^�%Ͻލ8��3y��缼q��|E�����RLh��ȳ҆tȖ);k�g����?u,2�ZW��^���*�d!��|��M��,I�w�Sz��{��'W���"�>:������:hJ��Ƣ��UL�D���8�s~+:$!9�� 'aN+&�ng��b��j*k΅�����HG7+��<����#�ǩL�wq���[N���+�ŁWR�r5���{��M�#n��0�V��_*��)ə�8 �A?jm1x�>ս�/���U�y�^���UH��n�i�ܧ����<���nc�X���B�RC�����=c��VF�/��)��z��Ab�,��Y~�8x;�=���~��&}L9u,i����v��ɏ���36\�o���L�G��Ђ��U�:���X����yך��aw86Ȭ�:��m���[mZV�9�Ξ-�떃qH*��� �����-���N�M�-.�g��-�LV�i����-�s���Y�1�Щ+4����d�P9�Y������.a����j��������8����V�-��;�!�����KϮ�M�4�^yt���#y:a�	�D��{���/b�f�Ǜ�3����7Vr~�����P�F���\�<��;3��y�����%���3s_��ڬQ+�q}z����{ң��P�'S�����VQ�=�]s��;����J�����e)��#��-�����?L��U���;�m`[�ob�q^E��?T����{�\�1n�Y[��}m��=It�SE����~}���򳅪6�pbt!� {��;v��Hg"[��I� H]%��m	�Ճ&�Ų�������M?���w�qdQ�(Ȭ��\�-w�h�����D�/ٓR��F�jrk�Ow���w��P���Yv�iM�O����11VAV:�Z2�m-\��$�fN�1UX���d"+Ƒ�o{t*�{��㾃����|���bbU����l[ꋴ����j�~k������u~ ��m���o��{Z��h�xi�xD6,�R�m��=I�wj�]VK�c���t�v� N.y�<ǹ���{2��d?=%?(�l-�>� ���9pK��Up��~�*یW�·�a�^�ݨ{�v+%i�a&�^��C�n%eq�Z��<]��6��jM�ĭ㓂�Y���t�#z�E8u��7E8���:f%�d�Mc��(�#����)�*|p�l��\��v���o&h��ƴ�܄�J���N�_�_'{��@�=]�<��f�ff-%
���C�t�ooӶi~T`��3������Q������O���Y���R����EE��\�q���~o�MI&+'q��77j섰�����9{9�-�^dXxv=g�}+��؂ ��Zl��[��6�<�<��և����lܷ�y���b�1ؤq�*��bA��=��^�mmO|�k	U8�YO�AwLݏn��Ύ�	m�DN��vS�ˡ4.}�.���:&�.���]r/턼�`�P{l�[g��a��m6�5�'��f�x�e�ҋJ�+͂��ߞ�Oާ�/Pyy�;�fZb��o,7z�	��ŸA}=��3�r�^_"�'{�-g�f�[��HJ�*��d��g3�d��T���m��R��Â��ͥ+�0��8�����d�k�sL-F4�W;J�R��}|�o0����}��)�gV���_Õi�]�~�d��2�$�{�_ݯ�^˸�W�}��.�}��<���c����t]t~#�)�N������o�mOw���Ӥ��D��C#��O�{��a5�*u5��#��&�U*Yje���[�]��bW5�\\"��V3wX�� �[��rũ%��޶���.FlI�[u�`�k���G�Wq�Av�
ܐE�1ôQ�u����`���ȚP+�+$v4s��}�,�d����"��ѐ0�ؤW��Vx0��9��\�9(>������钱@��n������FN%�}����{��RXI]�����k/�k!V+�>ӔW�i���˻�[�|<7��[<����k�D=ψ�d�ZsJLm�R<�p�{��Z���y�T���Ӓe���-���\z��Q��?��?~����|��i�֑~��������ؔ�u4e"�<\�L&��V����=�9�7��֍�1S��8x<\�\y{�1.�����)r�:�<7��ܡ��czC���.JMڼ̠f&�h!Gq���/S�p���>�3J�CS�דd�Eh
���;��BG��E��n*�.�lZ�h��[�6�F��d��*[b�ڰ�������_O�0�oE�(X�"[�f�A�M󋝺v�]��f��]|�Ա.T��f�Z3yG����ֳ$B�9�!���=X��9���>�w�f��=���Q�g;3�RB�w��U��.i�LB3����U�l���ر'��䭚n�����t�W]����)T��]�븛P�P�rG�J��*}qSW[����IvsۣtK��'�U�z�{�͝�u`;��b��(����,��]mg��2�"֎��TYQ֦����un���J=|$�s�4u��X+�ɻ�v����+�W���˩'c�X��e~��Wo��3W�G>�u�&N
��=�q�Ȗ˩���S/.]*ٜ����%nX�	q����­XȭV�9�!j�";r��]�֠Х%��t�3_�g���k�x��,�wb�O�8w]��m���8L*ݾ��n���9Vz^�h�N3B�#����n��ie���
��J�wL]EE�"WP�P�ʉ �\��˵���4�\��i$&n� �DH:�]�J3�.匤T*�Ԗ��J��r�=֔��d��0Tbɔ�V�=�M�b<�@��T��R��]J�_2+�j,�����:�wԔl����gjo,7�t$`*�<��W�e�7�u3d��@dYN�tf�u�zn��[ӫR�SuXe�|a[S�b�w�;k�.�u�:U�k��t,�5�+�%�;���R�'� �YZ#-,+m���ZV��Z�bʕ�*�U�
ZT-*��H��b�Pr�0����$V���߰SUdZ�JU��`�*�4Z%���ĭX"V�me��j��J�-��TVҶ1E�FUE(Դ����Ԗ�Z9i�RQEJ2�Z��E��%il�Z13fV�l�V�)inqG���U�JVZ�D���ҍTkd�h�*�+���ʕ�¡KH��(�mKj�h�)ZѶ��j`��QU)h��X��*V��p�����&�օbR��D��!J�jc�%jЪ���j�FVĵ������Z��EiZV�Ÿ�Vƴ����(��.�F�Ȳ�Z��Ym+mmQ�eqJ∔YT�`���1��qb%��v�s�^��ʛ��u�}�Uҹ�-�U)��Y�#%�N�M���'�iiě��_���/��{<V��9CA\r�$�k]�׸-v��+�Xu��v����x]o�K�b�J����u5��츱nu+���#���WޟO)K�;�h�[��ׄF�+�DD�Uԋ�3����.�S��:�$)8�<r��(����Y��;OR?�����H�]|jƉ�,�,��Ⱥ�F&	�;:�=h��F�����};^��y�u�)��yU�r��u���q��F٧����A[��E�����J���+B�+R�a�g��hW�39ǽ�[�e#1f=�EA=�{j��@�]��~Qȃt}�� �E�Z���)��}c��Ρpf�9���+$�W�¤��J�>�����~Y+|��>Y��]a�"*'�9-G绶'Y��j����7S�t�n�뽉�B��yo}��^һ���Zq�J~�=�K�^���.�*ȖNx�_(c�*v�e_���=�SZ�g���ܷ77�)菾��Hj��\��y,���$h`w�N�H\��r��ԮF
�����p����d�m���P.��g*�:(&Vt��m�=����9O���m�.�?P��'�.�/ֽ�7Q�]�Jݦ���X���^��i�]�>��슻Y�B}��_��t���70
\���K�-j����?�T�?��H)n���n�|�5��ف.R��sŭ�of�)%$������=�=�\>�*NʫSi��y���4�W�=�̽�Rwb�{:�C���ܼ��8V�b�B����8+��Z�L��Ŧ�e��Z|�8{h��{��9\a��l�y6����f'o�*k<"�M�he�;��tRf��sP�m�=Y�w�S��j�i1�ݭ��X7� n��rqz��z��)Es��bn�
c�����.����������e�*��d`�pi��݁\���/9�w&��^ֹ%�2�ܐ2����fRmZx�{��b�4G�]��^gp�W����_9��TovЪ�8�^Wp����7��N'����āq���V��b|�h[*� ���˞�}����Sm�?�m�nV]���JK�)u��lg�(c��^iԹcF� �ZU����o.�}���J=�U���.�ʶ^1�S�N��x�X�O�8s�z�Z����>T���Rv��y����@�;�!�]������p�̈́�ɟhu�2�_3f�'u�'ʕg�c���������9Bq�d`au�@RL}dY>`bZM2|��/��B�O�q��!�N0���}}�v�w?{��΁Y'{L2`g�$�� �&����X���ؑd�a>d�=�	�C42� \s���}�wg x�2�� (c�)|�Y�3�Cl$�d�Hy�%p�5�d�r�m$��>3ܯ�׹�=�|��C��>Bx��SO<��!�3�M�O����I���2m�I�j��������������>�:Ì��d�!�&S�a y��!�>RO�Bg�SL	��6���R��������^����V���M��tw�+��/���ow�}� �s��]{}�_��ה�{U�2�7���I*�&[��No�f32��7iH�i�Mߒ�-�����]|>�C�~��`)��<=�4��͆2u��8�� iO�0�2̞Sl�$��N���w���d�'�Rm �'w�x�ɺOZ�2��8�Y���Y!�{��!�O�&�
byB|��<2g{�]����!�e�nXN�2u���v�ē�8�C�E	�>d2�`,�6��m�e$<;����Ϸ��Ӥ�N0���'��a�՛Iē�I��Of�2LK�B|�͡�*�l&�
i�i��y�4_5���~����Cǽ���ƨO�6����4���q��3���!��L�Ї���&�"�x×�|Ƴ�y���{����!�e�����0�:�4��<��N�w�$�њ|�m�:�z���$�8����o1�l�GZsۏ{�������u
�m�m$���JI�M�{a���:��,���4��=Hq�����8b��o|�Ͼ�_{�zp�I�O�Hkt�BsVE ��`yJ�m��m�a�N�=`|CX�4�\��o/y{�|�u���M�wt�fXJ�i��6�6���CSL+d��I�M%a6��e�Z�>3d�C|}�����w�:a �$��i����>d4��:2C��
I����ɦM�w4�4%m����M�W�B��ׄå��F�~���me��$�Y�>��Q;���n��҉~�h�)�C�FSމ~g-�ɮ��K�n�'/�h�H�.]��nw��w���}��߾�����tݐ^� 
m���m�c�0�1��fu@6��'�>Ւ���'\�k~g_S9���}�uӲq��M�qB|�c6e� d���!�l��a�Մ�m!����8�cT��lv�w[�c�����W)&ݲ)6��!�)�'YL��	�;`x̲$0��M�J��ӈC��`,=�޵��@>d��$�&=�$���?XOX�:�q3;d��<N��I�!Y|y�O��C�yuw��>�s����C���d�'��=d�&~��$3��L��x���S��Ԇ�Lf�	l�!�Czε��ɣ��\ֶr@�9a��(d�8��3vY:��ɻ�M�o���Oi=j���-�d�%N�C���n��{����!��Bw��C?Xa bӌ�x�yۤ��'���˃�����L�6C�e�vrky�|�������z̠z�t��H$��>�����8�2M0��i���'�l���d� ���{�c�s<���gCIXOY٪I�ORM��y�HPņ�i>a�M0��!�N!��ߨC:��4�y�$�ĝ�}�;�g<����C��(OY�ȲJ{Hu03i�@�VJ�|�d���!�N�C�CL�a��u'҇��������׻�Trsç��w/�`����/�������	��Z��ٰwe��3�ʭn/_��sU-�W�l.�=��f�]Y�xƢݤ�P�]0w�������s~{�w���I?-PɓXm�z��8���!R$�l'X�I�M&yd� ��N�H(mI:�G���������6rHw��ē�`i����	�2ɓ���o	�6�@<��>a�0�Ӭ4�6��k��\k6����w��2e�AH|C��L{N��|�a6� ���ē�fk��Ց`,���q�I�:��|�}����Jɔ��֐;�d����d�x�d��4�l�l0�!4��=Cl�C���kY�>������|;ĕ��m��'�&l'>L�a���g�A}B`�:��8�=��u`���٤l���{�w����6�|����'���'>I�y�Ha
�$�d:��˴�����!�q��B�F�:�s��|��9
�m�Xu��XC�l��k�q"���
�0��d4�a�R�XN�2yx�=�|���s|����8�T�)�c�L�t��l�@6����%�g�E���L��Y!��:��K�k�S-Ɵy�kZ�О2I0�Xt��h��d<;fRq�l�n�8Ƀ��I�M��RN'ۡ<}`f�C�������>��u�u�l�N����@Ψ��Co��Xu�0�Y��{>�8�ǉ8���o�Ho�Eb��u�3�7z���&٤O��8Z�nuo8s`̼��L �h9Ӫ�o����"+�]�f��ANC=7Pͨ���*l��S��츥K��m�Ԭ:v�p����o�O��R��������U�>�eO��>d6ɓ�P�!�l'�4�3T0�1�d�	���M2q�&�C/�Ǟ^�.�ֵ���OX7dP�!��!�f���ē?`:�<�`)��OXm�SH�|j�d�z�s�k�s��^��vd���O&_��`���%B~ɪI�- ��I��&&l6�X3a�N2iRk_��s~��;��2M0��>d�	봓/̜d�ܡ>H,<J�o�CHq��v�L�8͆�9>��s^�y�=�Ӳd��4�|���a�x��d��$�'�6�|ϵ�I$YX)!���'�4Μ޽Ͼg�w]���Ì�d4�̟2m�RC����&�<��6�cV��'m�z�$*�� ��f��fw�����$񀌓l2Λ��i���s�!�d��=���?s~���.o���?�1�ꃾ��Rђ��kͯ2�d#��{f�W��`�+�9�.]��x=x^�a�~��r%c[qG��ö�L����g�0���ᇁ>�;*FV��X�t,�ahU"�˸L�f�Nx�~v���a�;�q�{�>Te޶��.��Ȩp��S�̨op��W�Dc�/��\�h]u���p~��9�k���L0�R�3q�b04,��]��^�J��{���r�^"C��fF��i�4i�PfC:sPҾ�н��g��3�qR;S<Wl�tS���xX��Ӕg��x%��Y)���ɤ�6��5�]�+X}[G�C^�}r�o~f��C��l&�[ť��^��o��Z��9y`׽��$R����g�L����emX��2�g�|Sq�}{1i��v��Y�c���Ԙ�.z��l����[�I��W���s�N�����Gw���N�ن��ڌxFPC���jf��\^��_Ƭo�����Kq�z�����<��ҜA��i��˺m��D���|Y)���|ӳй�}.�*�.��Gͤg�;;Ն��gC��vq�
���]X#x��)K�;������餦���Nx��r�WˍFr�`��MAg^�4��w}E��O��]�T˺�o�F����+h��Ou�l�,�h��%���u2�ګ�e��󛊨�#ѐ�_����*�R�8U�2�缊����}��	�ɘc�C6�T��Y�y���.�8�7�c>Z�w�,�l�7��M
v�[po%�^f�[�V'��� >��<G?~��wVb��#:J��x����˛F��,�4��]�v�"p:'�"�4�����f�����p:��\!J���d*ջ���IQ�$I��ұXgnhc��;�}�b%�Λ���Ӱz�t�)vD�_^1
��U�L]1��Wm\�
ՠ�����u��*ܒ��n�ބ�˵#�^ua-�P��q��Ⱥ��+��@܌*zΩ�^�����q,����6l����̻�l�[�ά���.VaVc0�����hn[��=��ᷛ�c22ԅ����=��E��誹��6�i���m�ݥ��s=m�^�Vs�6�6�QN�-r��N��m�/M�gH��v.��9`Q�;�&9��%��ma��,ܠy>����[�n!
�]#$���g<tn��}0g+;���%f7Q2zl/Qr�۹ʆQ�`�.�����ڙ�$�u��N��MAf��}��������޺)hq�+��T:�Y���EZ�,*']dBf������F�7қWo;+5~�X5�(�S�6'k��"0�Skq��Lv]�q��Ż���� Kd�Gv��3�������q��Q�bj��t�.g�]g}�I�(bUՆ�Air���c�7bG���?$�ಱ+TA���}��yh�>x`�3{�p=���Su^Ψ�W���x���<HM�V��ٹNGU�W�!'*�ɽs�ǝ�x�ܜ��mu��:��D�9�u���c��7�Ӎ�*}��4s�;�fDo�|�NC+T.u�׳Om͐m^������̴/CbeL�5�����Q-��7qjC9�Z�.u�(yWv�`_r��;�e��:Vވ�z48�� J�Y���ԩ@湯]��wc;;Wo	�=��b�/dC�7,��q&��V�,�ʾL%�v�&�/��+��v�e��A᪲Z�FF4����L�|�_����~�N�X6��QV��
V��X��jQIR�hUEsefQ��-m��`�)[Z���0m�-Å�Z�%�a�+ �DT)�X.-�,�Ŕ�m�T�R6�h�h���R������J�Z��\c�TZ2Z4�Z����R--�1���4���X�����&�ۆ�+U
�ŕn1��+L	�p 6�Z�R�ŵ��%�kjT�.Q�c�0����Qp%J�\)��.-L*U����1im���̲�*�+P���mhʬZ�Yhڑ5�P�j�l�n*4K`Ш�h��H���Kh�*a�KR�F)�(T�0��Z�F�DkEm��)b(��im��j�.PPGZYVѶ ȪT*UAVE�+*,�������f�TL�6ҪQj)2�L"��j$D�Ym���{�����~?�*�X7��Jĥ[2��[iӾ7�}(�lg����'Ž���|>��-7?W���D���cs��I�7�B���W��B��;��pn���c8���;��~�=؍x���I���ƃ�2ȜϹ�'aE3����v���٪����罩I8��&qNw5|�yn��k��֗^��Eמ����ơ�;���vc�U|����6�&-���[q��$�{S�c��>����M+�6�oo/?P�g�G�T���!}3�웟���i�J �Z��l����z��!��7G55���I��4�~g��j//���gW�����A����Y��g4����z�?�cw�����s�~�r98*�u���թ�`�	�T 6F�1mw��Q����t��h�L�������m�����b�k��������LZ'flE0�~��a�d+*�W���s�R�'I�g����ꙊN �k�;����Y�׳��d5�{0v���yz��o�����@nG����~����'��5�Fq~4��b,��9L�R�k�g<���7�Gj���P�H����Q�v+��b��,�9I���QBT�3���U��*�0f����J�ɕ��i[��(��/fv�k7���������op�i�#�b5Ez��oc�gn�I�a�7�]�=+5���\w5!}��eH�i�ϳwوR��f���+2��<��OMpM��󩫌Ilܫ��ܬ�5%��'�-#�!�|��| ����� ��~��K�N��u�v[�o��^ĸ�S�އn^K���b�=��� �Lx����qj7Z[�����X��o�HRz?U�X�N4	C8u����\�3�굧a�dU�����bȮV�׷��Ԙ�x����E}�V�U�����>�s�T�zU������[�[�wg�ťBoeE�	�ss����8���H�����+X~�:vڅ�zg�le��My�3G����L��	�[,�QO�yWo5��ŗ�I�=d� c�gb�\�V�,�������1���������gNf���p��PQ�m-�����+�:��zs.���mM�O�˒��|>�L�&8�|�yh���9zwG���k�[.����������nn.��z�׻o7�P�Ô�nh�-3��䝀�x��0����[����֊��z�y^���Q��m-$2p��L#���zQ�CV|���xE������w7�-���_�U�F��)It�Q���o���Jn���c��-��{�.&1tC����ם�)� �a�w�ZӞ����������v���U�pw�N������Ae.}r���Ix���#��v��j依s�^w =�b��K���oA��H�x�%��%�ȧbs!x�
N��b��U��XcR _r�L�ˑ�^�;�8�W�c*��[���}U����ln}���U�p�W��32�y�z��9~Q��;&�ٻE�u~���c�Vm�-srrQa\'�V��#�El�'�z�d,�.�ں^`�p�����ڼ��F����ڃ���'�]]��B��[�n�>��:�cgve;s��U��EMu�1hƹ�>�:K�/_�ڭ`�%xe�������#F6�p��)e
�2�Ϯ������Ϻ���މ�q�����[�O�X���ޡ��=㼃f�̅�c��/Jx�P���D�Aș���d5�}�z�%�F�G���5�y��f��-ϥ:���n�8q+��k8ٝf�S[���C'gl;����}U��U��1Ͻ�_���VnY����,u�k(iF?wUy8��exљ���S؛=��߮�4Tr>�P�n��Dס��=ʽh�
��������4L�ҏ�x|�*���u2�C��F$���
�ƻDʼ���Ӹ�y���{�4��b B+�*�b�K�Vr�ܽP@��Ws���X�ד��*x�y��M���j�^��g��Y�,�Ϳ=UV�r��1mLf�=�ۇ�^�kڎ{�xy[�p���?q��+h����+��Z��=C�B�G1��r^���.�Z�������~k�[�N�Ѝ�Ux���#���ef�n��I�4��5�V�^Վ�9P��Y:fe�@���?+����Gp.����s���/7�a������~0��ptY����j�۰^�U~ݒA�#y=K �p���߈ެ�Ʌ)=�5w���z����`�j������*M�'���^���y
=��^�滪�sGokI��)g���W;%���3N��W�5jOޤ��K,t��������'�s5�ضNʻ��S����/�+_MI1��炱�A�C�M0��X�(�e���}�#�2oì�Vk�^�kCl���*���V&:��a��i�6z�G���]�K	\f�����cgH�W*I\�n�v�$�Yq�\���6�>NO�������"��Ɓ�K<�������\����#I{n�	�J��ʏ"��ϵ�c�</ؽ��f-��A�%2���3Ezf�fk�9&t��C p;�-�'�v�-��t�WS.�cݚb�kLOt��{v�_��8Q�(�}�0�g���Ϻb�c��sWm.�2��ּ�n�w{0��d㽅w	[�������w�#�F¾�-����y�9z�a�(��s�f�W����0�0V��e�L��Ħ�Eۂ�ǹ�VF��m?[�l�Z]�(�zT�N��i׽�c��5�~���ze�kٍ�<N�Ԗ����1\��\�+K8�����C�Ar��kXvD�K*��G9ud�ơ6���>��>ӄ�n
�~��s-%�\hF@";(\�kr
��=c��訲[)�2����<�P*�+ge��W��	�섰&vOCT[���Q���l.�;M��OI���qzy�㛦!HIU�>�����C�{3�&c�N|��%8í�7KAD�v{E�~���΋\9zI�zV�T��t}H5˙d����A�u�>�����']����A��T������c�{}-蜭�4��/Icܺ���*;���{�[P�T�0�C�v?"��^�Ǽ�2��;���:���gY�T{�m,)i���Mz.A&�����z+GU���!�-r��N(��N����t�.�uon�@u����̷��ও$����w�OiA�T1Ss	��"ȋ�ח,կaQ���W�����{��ɩ�=]��wtM��b�x)���E����k��#�o���bX�0:�r�M�|�*Ǒ��C�
>��~�~�����vO��������>�Xҙ�.��z����g��������9��N]�݋�q����9�i�ڀ�Q;� �=G�UY!�]:���n8�aUG_ly��Цb�F�p��.Umv����*Jy	+�"�Vh���Wi��۽{[��U�a�HDC��:7��2�`g��S��D�ْ��L����r�^v�wL��e����]̧����E�Z9��]����J�u�,�L�kl�ͬ\���7Q�3b�J��<�G.���\�T5.����,��N�\�Cw�س�����|���F�hی*�Wn�(�܎ty;+)%u���:��K�B��Kp��k@��zq����30�xj��
��<.�fـ���o:��qr%ƺf��f�1�X��� ĪX��Ըd������K�W��Gt9�er�=Z���-£w'2��y���@�������
�U7��=B�`�U�vD29gX�Zݺ���tvo`�ˉ8�\��D۬�5�[������76;������U>�ƣb�]Eu+,;r�^7��vm*wk�.�W#��i]t���)�����պ�D]���E�����Avv�-I��Y�o�!g�'���^+�ag
�9�^���Y�vs���z�ҩ+�Ƭbh���יCW`�[#��V1w�t��PAgr�})���PY�L�90��r�i�˵cS���K%��V�MG�{20��̊W6�]�X�b�=tnҏ8,S�8���(��'L-��:����CuJ��&��r���˝��9.)8n�X ��%����>�gv˻�����+[fb&�,�L�KG#גn��`�OE��]�<���.��hfu5�z��燪눝M��e�ܯjn�|�+b�(��]W��gB칐��V�Ar:�pD�P��ʈ��IJVt��dr�s��E�v�|Q�<o��ͨ���KUR����em����;�{�T2@^�93�C}�usf�E>۬��w�}%ǒ�Y�+���6L����1^X��`����N��@8~�~X��.� �k�aZ��"�RT(0�ڵVZU�EjQG�V
�R�[e)e��()
�����J5��d����D���,+k*-E+F6�¥b�%Q �QJ�QdKqq�m�eemkiX
��2�.FVT��QYm"�D�-jT��U�J�@�نf1�TKl������F*(,�jL�0��,
Ȩ��T��0��6�`VaZ�(b�R�E�J�hT��*E��%sl�J�R�EZ�YKaU�HU�)l���U�%kE�F�8Ǉ����e�VT4��r�tt����.XC4*t�\/�e�Ts��}_UW�LjH,��:�� ݌Ǎ�D��??;�#*h�۾��%6�Uks^z����j�{R���<I�������g0����>^�5�H)�9u��SgK�Ȼ�x^@C]�s�M�9�;�zo�*�?{}�nmk^T���J�cF&,Eӵ��j�S^w:,�յ���g��z�b.I ��LBʏږC�%-]�:��Wgi�.?�
�h=-�:���|u^`�yr��eD"���l��"��hD����� C.3���}��6���~�ņA�М�"����|��]�Z��������*�W-�}��=�0�N�7���Olr�.�|t�)j�(S�9�7r�����t���ӭv��{[ۥ���M?�}�� �IrH���2�^�Ƈ�R�`�/�z֥�G�@�gNʻ�< �8p;2���g�-:��i�O
���	����NO*}���o�Á�y�^K"B����ݑ�ұ!�^p�w�آ#��֞�y�s�]�"i*ߎx'���y��7�`'�$p\��Y��v�X`��le��E%��1����ټ���bڱ��DR����}��&�Ԩiew��v�_��8҈w�s�Ȝ�vWnIcq�H���Ǳ�!]U�����X����Gz��[�
��9��z��:�݊�f��}����zH�,�E�$��Z�`='!*��z��T�6fQx�	d��?+��6x�	�*U����;���d�;���wۺO�(N�4�}��'=��цƍ�7��>n	�V��Z�E��=ޞ���)�j/�Mj��.�w�2o]�m��|�B̓��֙�1.\hWM7l���gK���m�h�xS�����JjxWO���Ӿ���d%�ǫ�b����9׵W����!�ݞ�w������qQ��P��Ux�>��1����e�qy�#a��6����{A��3i�+Xw�[���'�-+ښ��7�~���ۜF�Y`��wF]+�:�˗���Ky�9X�L�[R0�,neN_|Z}�mV�wl�v	��|�Q'����Ux�"��q~�ضq#�>�پ�rXfƚd�ʋ��zV�Q� Z��X�Z�^�NpB�����y���]M�#�sK�����uF��D�yM�*x�*c7)����5�#��3W�~u������=h�դ���R}!Ҥ�2չ��ּJ�8��?A��5U�Ɖ�|��a�[�J�G�y=�޾5�J%�)�W����5�*8���M��$��=t弐b���l�.�{�/�h��:�4߯+i��\���5UU����{pUeuQ��y"*�<Ơ��0+r��v��vK/Y]f��o��[yp-{�b҆��a���t�X��}n��|�A��+�a^�<����5����f`��BxO4�|>�|\�K��۠H�����xb\y��,[��Dڿ�@���;�=��� 4sP�|��v�#�����riPUK�����xda'S�|t���'ZD!H�lS>���(J���wo�-j����L_�di8��1i`����˪����V�|0��+�R� ��Ԉe�c��xɕ��uR���	�%#d���]C�H谸���g���b?��#=�n�̪{�S�ێ�Z�8m�ܯP����F�ۣ�ic�;����&أ^����~�w��LnAF/�S�|���aP�x�/���d�Ϊ,5�8����Xb��f7R4��O{�v}A�\�b�Ue9k����;Γ�H�+�{~?c� \LY쥎�Ǒ7�:��x�Y+e�b�[��[u�]�.>g.��g���X,*��<B���2v��k�=i֣8L�'� ��P�fw,,�?4o]��%?�}���ZRxL:N�_��8���*;�+�1��D��v��,=��L����!F�gpy�H�=�=OO�SB="VT�h����m��b|e�j�u*�i�LT��(mz��m����X�vx����;�1�k��@�`�B��Ć�~K��rQ��{ɨIl[Ո:�:𮬦çH��/���O��n#ސ���ӓn�Լ�ϲ[�ެ��;t�*�0��d�e�Է�{=���[�B*cՏ��������#�q����9��V�ޞ��{���D�|E�K�I�x�!t�����g��UA7�[ƷSpem��I��O�/1*����NJ��=>��V�zfq֛h@��W��U�L���R����K��hQ㛥T� g|"�f�CJ��EhL'�m�VNA*�vqP��fA��3�He����7n��ڹƸ��3*R��,wSX܂DY�m�
�-T\�Flc."n~}U��u�2G�nǫ�U�¥YD��۵a ��P�ث��^:�D� �u�;�l>�,�,9�����q�P��G���Vu{}�I�y�f.%���B�t[���������;Te���5��u<5�Ŝ:>:}�6f�!�8�U��{+w|7���i)iacõ��_!���罓�n�@��7�Hw�O�ȳ��$�M�/y��>x`�?]����JF87~�Qs����;͵Xs>ϩP��vj�[<hW}<�N���d�w>��v����b�kǠ�f@�ҳZ/(�r����$S�6��X&�U�3M��J9wARV��ݕWGPש����'����m��M*�����y�N�w�zRs"h��h�ص���%�NY�1GcWi�V�c��b&�8�Ϋ=N��sy8��<�
e*u�B�����t����<�VR<��o��|>��w����2o6N���m
8�>B����-���v}}���It��6��<,/D�a�7�HQ/R(��2��������1i�OW�
Թ�Đ��C��b��^ő����}�j��+�0=�5��!���j	j�D��Vz�2��D��
/uo�����q�v��v�7Yۂ��e��^���t�PmNZbC��Lay�8x�YK{3�1�����gڭ'�ֺ+�Pv�wD�+6�3V7�I~Ѱݓ��
����*=�K���"�妄��AX����3ٞn3H��}�׍��E��;k0�B'ͩ>O>�^�����ww�nq�>;9�!�5�r�/w��AZ������.{S?i&[CՃn��x�̺*�����_���Ŏ���n�N�����iR��,�����bɝݜ�n"�ݽrT���5�_s�K��)�� n-E8�'�yک��x�?7���Zh�C�kG.����s\JAà���t+�;۴mѡ��zZ#�<
�+�Q�Nt��X/��/ �����/���	I4/Xc�9qS�'m�]��X��,�������1שi�4`:g�
��xWP�������DY�4��H�*πKO9'��x�WZ�]�v3� ��\*�c���VP��-��-���;���c��M��C��%�O�<t�<p���I7*nu�<���'��D�`��������	y�&/�':o�%C�Z���{7�C8I��yi����b(C�eg�r�<IKg;�Y+�{�}�e����J���ޗ-�-Y�-��<�{g��Ո��&'�>lTa�V⫣�9�a��.����T��b��_frU�&1��0U�!C��Z�V*�Gt���,+6�#W�2������
�y�U�~S��O�Z^0j�|x�LT��������%�my.2T��z<�6��
�b�E^G�4�<Q���}��U�U����J��6��I<u���	��;׺:Va	if84*N����پ���'r�LvyP�j����+A�iv�JQˮ�F��S���lWҋ����a��
�ߵ`��OtY#��E��+��䉶
�����͝Ha徧¾�nΈ�BϚhb�ڗ��řu������Xz==K�Casӛ{LZ���^��lR�o�k�ܹA%��I�x�5�%��E#���p:χ���O��|`8Ya�<x�Ff����O�vӾ8t�_�kz�o4��r��^L�i��M�R袡g��M����aYK��T�չ�ّi4+����Y�u��|�ɖ�9ܥ`n
xt)�[</e�Yu�3����k���js���"�ׄx@�rZ���Y�2���M}^<�¬�f�Q�f��ga5e�*�E�U��걍k����J\g-��h|+{�[�	c��e�&0���Go8��2H�ċU�nl�QV�v�e��JA�y%h���p��W�8��D��^o J�ي�4���D0����j�)�NV��1���ǁْv�!�yw����ܾ5�pJ��ՎV�=D�Ab+j1��3m�� ����"�&��M�S���b]	�
�lv��w�eJ�F�yn�yj>���qp޲G>�qXV�c72ХK1\��),2�XvŘh�{&p���\ٜ֡!�H5´���n�7t�eN=.5
�̬�\녜:�Y3�����RS�2�wt�u%K]}O�$���7��q-��~6�qx:�łΞ+�����W��f�j�bdv���@��ſJ�Y�@�9�J����{�t1'�-�0�\a�1�+��QU���+�B�ŠDwX)�>��%s�{���5���]�|�TA��<�����K(�sEL={˵��ȑ�9+��t��V�NA/�{�s�P3Pߤ]x.�<���N-��ɘ��v,�V���K�\�)��ۜ3�c�j�&��{��$��Z��:�;F�-�I��,�v�$Yx3���{})Z�̂�M���Y�7j�X4^S��뻏1��w
��vao;/���ZI�f����G��|1�u��Vm�6cyn��Ӻ�5a[�%/�8S�U?�2�R������wr���ܘ�r1\�GVD���Z�%a�R�j���%q�'��K��q��Î���d��'��)�$L�^K��3G�GP��<���}�xg���c**�YX�֐����V0�T�
�V(V`aQ�Qa��E+#i+
�Ң��X+L�a%Ecl2��,(B��3
�Ղ�Ņ�J�T�AE��X��`�Z�Z���PTjDJ�T+L�QE�, T&���EG63�EW)PYm�U
�
�*TAG8�"��(�E�X,"�L2T�HT�[BT
��PDYXE�.��Hņ�RaU�..-�*T�L0�Fұ0��͛߾��f<�t�jj��n�S�7�Rlwu}1�B��N��L�Ha(���՘u��wF�iQ��ȡA��� �o�ťǉ���c�֥jE�ۤ��$j�!�8m-5
5�|)��	ug�/{�ߟ�w�Ӈ���I���=l;Ʃu��/��JC���J���{My�~�d���	��sHb��`��|��wEhMUh�����Ii}*�q��s%�;�C��F�1G<�ֆ۽���b�
]���ќ��{�B=m���vc�6a������UL7/c�dء�^�]�zP<=@u�7x�&���^6/�R�k��/����7ݎ��n:0Ĭ����KO
�ܠe���o*
o�����u�N��M%��2�<<�ƴ�؆��M��܇g9=M��b���+�-�|��G�G�v6Ε���UE~Xt��ٶ����Z��)Q�s3G��5Q��ʰ��������o9}�}JN!.�Pr΃[� K���M�S�I����G.��x�{pӥ��|�-7>�>gH��ZXA
�t.��*���cI�yاo��U4䠸���T����S��r������]
�ZPˬ���HK�����m��,j�f��z��ڢ~�޻��%	_:=�^��ݵF^��OJ�����pG�����Cqw�C|��$t���o�D,�F�hۧx%�������"�ap�ꃬ
��p� V�W �xNG�����F����wa[�6�uq����\�WT�U��V[����t3�O:�o���[����b�@t����Eט}����i��F��+���u�No�U���3��Ǯ��ϥ1^S���d�\vƻ<p��=U�Aђ��ݱ�u���a��|���Ɨ�āiğظ����&�����(�[��h��;%N[����뱔ps�#Ǣ�j��N�kZtn���S� �kf�3/RJl�R���E�0�
-����}��	5NN
J�}_�kkn׬:�{W�v:R�J]j��Ģ�g;��|&=_^���M��SR(��v��N*��������i����~���1`#7��^�B)k��f�ץ��3 �T��t��������9�����9�/B��r�#|}�/3��E$"�IY���x����c�[����7ݝ��7�W�B�D\�%��j� �ޖ~��X���{ӽѲ�A]�@^]g�j�zŪX}`�������s+΢������͍����I�^;m���	�#����>]��V���C}�\��x�#K˺*� �w�̖��\�i'9����	K�5��x�D?Ǳi�CN�B`Y@[C��f�ы�X|�V�r��T�0g���R�9|��Y�9+ng[ki�&aW��\��ܝu#�ZأLgu��˾�y��Q��:;;�FT���t��w���v>�S�I��!�t�<hb'I8`�H����V��W�xCZ�.8[�8�S�'��'~�0�'Q<S=�=$��ȏ�!�D�:\Y��w�7U42��B�Y+ѳ�l������[�᭫K�⺞�7Z>�})5�x�f�����:�zˀ{3�=��'����:Zw+]�����R����0���T��w�'i�,9>��Kc�-�|D�b�,1y@��F-�_m�0�����[]U7?��x)�k�㥯o�w��M`W_<v�3b�n�i�x�%|���_\_�����/�VT򠪙;����&I�wt�ѩsL��J�u�Po���[[L;=nh�Jo�; ��cvI&�V���l��!�)�|��e�#�w7YB��Ҽ3���P��;���Ȅ���=\Km�\Y��5s-}t�t���}v��
��zo��X��}��j�e�s���7XMo�w�}�R�8<��d�=�<���8y*6���==)��?��7�{��<x�+�)�?VV�����o���!�/�"U+Ŕc{����nW~g�Iq�\}��e�^/�kOEǋ<B�h�}�{�'y���P�l]/�È�u��<E�oO�=a<��> ���V�=0�|l�����VΧH[�ۻ�o��ɬ�%:W(�3�"C4t���'*��%z�^'�_���i���!��"�`Q`hd]:V�{l:�J�w=P��U���$�Pj���؃�K�z���^w�v|���
�{۞�Z|
5�1G5_C�.Y�nj��yR	�y��}�P�^��1��j�lk��2���\D�F[C��:s�Kw"G�U��CYB��a�4��%|����]|�6)S�F��A��P��%���DY���L��C�
���t�P���ᐬ�3��B�s��URW��6k��ܲ�(f1�\I��P��_.��\|)�
�[N�:�C�2{k�u�O^�UWS Lt���GO��!�+!��Oko����^P{X$Y�RXl�qa��q�UdX5����rF��=Mi�7�`�>�f�K�"h���\�����iw�3�o�Pj	u��}خ[+)}tbt��� �,�KO������gw�B��2!״�y��c�x��^>����p��|��S;��Z*۩���	^���؉�'�;CK�ȵ����r�����w��H�k�4��/��&�RӞ����:R��]y^����]�+	�v�%�掓��;o�D,��B��r���7�w{�"=�[Z$i㦒x�B��KU�%�����#޹��-��C
�6�.�|�Ks%�x�%�z�`���B���^���vx���}�+�r]P�o�f*��n� �����ۖ�㹊�ݲ�!�z���<2��:�D�so��<��O��.��b�n�~[�UN�A
ֹ����hJ75������]����xj^�<A������D�#Mٌx7~�g������r������w��jg���yY�����k]�;��Ah�L�l�q*ʁn]OL޿]�w��lW������؇N%��C��c�y�����Ga�w���ʴ/�o���J��T˄���|�Pv�ۉ��2��>�F4��Qc���>!�`�7o�H·U�\q>��^��ys�,�8E-c;}G���=��2;Q/����=����_:��f�x,��>1��AN��݉�>�R��;.^�{={Cd�������w=�*%˦)R5wB���uH��F�i�gG̶j��[��������|UG�;]<ˤ�^Q�-�2����Z�z�K=���KU��A�5'�Y%l�R�p鎞���1��~W�Ț�X&��e���Ҫ��@��u��߆Z���:�=�KJ,@�yi���������'5x�\}��'���uл�͹ ��s,hV���=��=B�/
ı�>pI�3�[r��o*���YgI��+�z!��!�\z}�O�1`�gl��>��� ׶}=�t�hb�r	Aӈ`���\p���Ñ���{4ɳ��;���Xk��<h�/e��*�'��d��Ru�M�u���M���q�c&��x�U����M���b>":^���F��;���O����q]O�֏E����=-�r�ސn[d2c�/"��6�*���Y*� �9r���������m��;�=9�(e��Y���y��R�1c�%֦��ܱGGx;R/5Uk91�:0����~]m��Y["�E���v8m�� U�o*��V��6���r�^�\ <�wLO��+��:��q�o��Fι�Wӊ��ߪ�ƣ���7,m�#��uY�i�T���چ�$:�g{�K��+��y�]Ds/"$i�0$�x�Ss��Ɔ���q��r�&��B��K9u�r�S�S,,�)���m�{��W-͞}�׶��^7d�k
��Vw�:��=�`�p.��U=̮�瘭�A�e0���+$��zz���^�����yq�[��Z���5�j�����D������_��[� %�ҙ\�d��J�YWJ�ۧA����m���\�v�p���K���#J�}^\E�ޙ����D����s5�;�O�rbP�GB ��3��H^���g�\��on�aJ��s�>�Hdi�Z��'*�V��م�]�z��k	Xu�����fR(eZ�1��5�]�ޢ������:�h������'�-��4��79�&ɷX��^dJc�vIňY;��;��ݽ��>~�U&����?��0�k	/�GS	
ĵm���1)6��Jׅ��O2���ن�a^�C�~j�{�=;��4�G��o���Z��Z�� �挿��~
6໐�Kw������8�oCY�QxɎT�.�k��Hq�0���Clcf���7_T�Ժ3G�1�s�E��@�`�i��|��,�~�ws�WA 
��w3���7��y��Ä����M����j�p�T�mJ�ny+�d��0�7��b�B�I��д�X��C�N�՗�u��	�S�j��:��8��!�q��H�,%��!�MJ�~-ʯI+������u�K��\�VUt��s T6�8�����@���,M��P�n];U9(.8�\�醽�:￧�j�.����˭͍��0��et⋦�hY�F��m��=B�Ԗ$��k�R��9.4필V\����|�;u^��^>T�
e��K�fIPaݲ����ܫ^��OQ�Z�[B�o)!��35��ѵF�>I�Vv���+zC;6�sof-�t�>�б�b�h�ܫN�,n\mh� (jd�*�<Mt@z�]��uZb*n�SAgnsw�NQ�S�Q'�Ѫ�Ί�<S��m�0��;���n�?<���i�v�����3��`,����(���Vט��@�֯Fa���d ����3*��Wxy�8�`dG'j��Ϯ֓��8��չb��!=�����Xy��]�]Jր���vp�������KB.�}z!��ݲ�er�[xh8�j;�G5�z�
0~���\�i���o��a_Lu�(E�7����8"ѾFm�V)ܞ�;���r�wR��¥�7I���ˮ�0|��mYݧ�V�qV��f�L��d�kc ��.;}�{S"��#\�1���b=���o�Z���O�c�����쿓�M�f3]�c ������h>9(���fg:C���Bxe��ԑ�}^�lm\��cZavCڡL���iݿ�NڈS[��#
���S]��h4���ŕ��K��/���me�&�c�z��`�r|X��$	4`�0zk�V�iۣ�nW2�&6�;;��a�| yE��ܩ�{�����.�,��GP��ǖe��������2��X-��� �\�]��%��p��BT��Y��؉�ĳ&��;�`�L�ζ��r�]�uXv�E۴֙I%�m�"ouN�&��L�g]�]�c��W��|2����!���܊��WT
������"�ZM�����ZҲ�T�Ȱ��lR��,�C��X
d�S0�`T�dX(
E�(TD�*J��E�(TDT�P��)X�X���Dd��*H(Kl&P��AL1VV����V�%�E[H��T�V6QX�HT� *$X1T`��B(�P\$*AE$Tb�QQUa �������t9�����)߸:��˖��,7�����x��w2��ж�����v/y�i���^]KYt)�ack�bB\OHb��ǖE��*���d�Q��F��0���_:<�@�F���<��k��v�f{�R�᩟McܼF�|�ë��s���Y؍
�n���q�[py�Z�*]�K(;˱���C�?]�5.�(l��7�L.1r(|G�Z+�O���qz��
�݅���w����]��6��P�5�D8�kJ8+�c��3�d�1.���,�}���
��ς�u�2�ۃe�CJʥ��d0���Jث�|9<h��h���H_)�-.\�Ǩ"7�v2�Rc����T�Z�ׯ��4i.�cŭvT��A��<���Z�<s�,L{�K��7V��
\��N�4��/��U��'���qVW�#�������!v3ծ^��D���;r�<V]���:]�%�͉��ˡlM��o>{:��ns�j�����ht��lގM��2%'���Js���~g%W��#jn/M�i�?|z�Wė2h�N�y����Z;<$���s�u��`�u��W���`�O�ԣ��+��s���5����A����r�U���ӯK��7�K��smo�&
���ǯZ9^>����H���;�Ԭ�)�(���8�����R�� � ��j���kFz2C�힤"V�w���V}�pF��Q��1龈�$��k��o��0O`��)zL���2���"'���<�!�4�z��X���s=���>� 7^�*�o^���t�K�ҟ
v���z������=��-�ߴS�^_MA)��0Q��./;��_?!�+=��x�ȑoY�h�J��,I�Aʼ��{�'~�+�5m�[����S��k7�W�n1݁�ʠs���;�䲹q��\g�{;'���w�m8�q䡇e.�	֧�9V��R�f�\��'n��A̝�Y&���1���zM�{�u�����DՕ�R� ���rǫ�4%]J�Կf�ђ�ʬ��aP�|gۭ��I��z֗I�y^~3�0y�^�p�l�7��S��Cَ^��n,[w(�ʝ������@�p���o�=�[5��?c޷�L�my:ϥg�Q��}��
���:�U^����J���n����pԓ��en�e}�P�w#�y�x��W���I�Z�^�73�犐KݝB�������Ϗ�b>�㜨���Ɋ�KM�����k�0j��0�j�+�l�$w~la���+}��(�g*�C{j`pR�fV<�j�UJ��4߲Ѿ��LQ�d���X�*ߋ�|����^#o�`��"v����ަ}la^Ҋ�HQm�k�8Վڥ8Y��W�����@C/�}N��}6T���3�c��u�k�����ZY�6��&�Y;r���	�̩ y�B���,wj�ۢf:/a�R��4��q�Nz
�
�����B2$�+<����a�i1Z�cˈ���{���\��V������a'Ntl���:r����$�U����O8�9N�[Hi'�sG��H��8m-5%A9W�SIؾ+�۾��I{�li��&�#��cZ�������?fU��n﫳=������)Q���x����^/���a
p&=k�׹W����P{�:�@KT�>����(�kctÖ/r���m�'WL��B��>�H�^O�|~�.�6м��\o%�Ng�M�g��(V���,C\���S�O�>��Z��;l�*�ﶽ���[kr�"��s���Uu9n�ܧ�ڦ+��ս)n���3�d���Jw��q�����R!��zyU��k��w�M,�1q�6'��h�݁;9���0��bR���v��h�>y����̧��p�$����{�\Ν��
�7Xi$�XhZe�xu�z-�;*��zHUT`��ڦ��47�`L{ʾ�0��I0����#]���|
�ͳf>xw��L�������!���s$W�/8�EK���x",�d�+|22��G��Z���N5�����[݊4�Z��Yu�L�bS5a:Z}�EؗI��r��\�={�O�Xe�5ay�1��<��?q��"4��Te�'�Β%�>�a�WK�	.P�"o�8O/��"Φ�U$�i������=�ڳ�vcđ��--!l^BC�-X}	����G�o��Xp�X|§4S�/5�qcQ<�K�ӷ�G�"��++3{�Z�Е��|[C�6��������`�H}�-���$�7_x���Σ�X�yI�(R������;e�T���_t��U���-u[�f�i��iD���W�tᇦ�r���.��e�ځ6���4��ժ#�������W���o��[�q}�6_�P*�e�t�Q�o:�x�V��j��!~Xtؖ��6cuJk}�.溞��bx*$�㼶��<h�T�JcŅ�ʖõ�T��Y�ݬ�Q٢��KR�
�׮Ƴ�����լ`�끾u�����Y���X=e�%�}@�����j���9ߦm���˘��"Z%�Â�����gv���c��M>����.`4k�A���[�n��_��r����
��ѻĨ��3��xΌo$r���F��>Wʒܹ������ڔgB��.����v^Ń6��h�k��ڇ~�l1�z95��H�<8��u��2�e]?��ˮ�I+5��\|��$�v^�Ğγ�Єw2?v��k�n���=ݣ�M+�m�8���33:+�i[�gl��nZ(�=X���w��I�v{y)���:�g_e����"5�=A�Hb�k��_S�y����6���n�)ey�D<m���z��M�T�ٛ�c�= b�߲ѷ��(�i���a'��2���q�X�Vywn߼0��HѲHʶz�!Ҡ-abM���_�`�N��9::����]� ��U�t�\Y�!�D��V�J���mk���������p�#��d�~D�,ә-�._١	��8�X��t�������uu*3���6�-K�	|�ŁZ� �g�wo�R�Ad��j�{]F �+|;���C���ڹ�SO�wC��X�|o��V
�s�\:�Wqj��>��o�?v�m�+c��e�M{���`�%5x��8�{ӈ�d]y��YY@�[.���U�k���N�y�m����g��~5�EeɤeW�m<�Q^h^r;+�-n���&�%��Mt��)?��A�����_�
v�o��Z�T��>��lV����<�w6�;zp{U╬
�/�I5�a�M�䎶}i�Yԉ�fAc(E2�:��}��T]�x3�ti��U*唠��gI>����z��=9k�V�W�m�qO!�X47:�E2�ZK�eW�z�bWn��R���o�+��ϲ�<5*�j��n|�C5�p�� �R�Xb#J�}���f*�퐙Q�i@��Xu(J�l����9��AGPegʈ<��Iu}]��txy�3��Cĝ9�sG�2D,��q�.J�,�|��;����=��I1�Li`yi'	�H�Ƶmd���EW6�#m��o{�~�mYՆ�
��c�c�������Z�#;w�'���&�}x�u�\�<]�#�p4?G���=~��� N�$2�Įs�YӞqY(�w�E�M=�&u���4��YN�����ܟ�Sܜg��e/���兂)�0Zg%:>��po�*�W�M�w&k|ԍ��O���D��>!���崆{0�-*�r���L��;>;��ݖUȝ6���>����k�7�Y��c�A��ޥ�����Vᡈ�b:0�g�ϋ��D�w,���	*�ߔ�6-S����y��&,�`�d�KN+;��A]�;/�ء�j��3��H�txPޱ���@�t�>��ڼ�+V���I�y\������m�]%�����>	m����D�~l����AV��5L�s#�v� rPϗ:߽r��^6��LX�lL9�����G5#Da߈��P�oֵ!;׊��I]ܡl�+>�����V��>�h�\F���9<Xd��MR�
l�Jؕ퓕��kacGI�Eb�$ݐ����|Wi�1zOL�]���]D�3m<>w
�2XX�_Bzl�Ǩ���y�����?����*@Y�H��<��&}�w�y�d�3�:b���9�6��l�һ��wȯk>A�:���		����E��$1az���e���g{xr�}�vX�R�8�9���|%�ur�1w*��<9�t)	%��J!�Z�	Sg�q,yH���(�!洗%�oٙ�o
$xy.��Uj ��z�����ަz��V��,I��v{Բ�`��
�W��_��P�f�!������7�H����Px:It�g�r���><hѤ�!�k��݃mك$�C�@o�՚uZ��x:Z��+�m��g�_WY�wCsG{Z��@b��a֓���6{�ǌńa�O���zx��W�ᆬ��R�7���rc㶴��1g���\��>�n\&�j�#O�Z�7.�P��r�F�q:�%b���Ab`�F�����.���rzg�30Ak&�BFq^$'S�����R�������e�d��;y��fTi���8���"�n��`cz�Ǚ��_L�FU��+jgk)�o����&��� ���0�׌���b�̖�|��It��OVa7r�-YGD�%-]�Q�
�|xѧ��u��n��u�$�_h� c/�ݹ�L��J+���vY�ӗ�������t����);1̥�1M�-#�#o���-#����]v�K(tZ��NE���N�+��^�4�D�����u��\D�si���ս�k7j��IH�)��:a�[�B.���Qݳ�B�ڼS1X��>�QLC�#w���������ZuSa�?	�6�h��塋Ϸ��H���aoY{I�s�����.�3ҲEe�XI���������+U��ܻ�k8[,M:[�L�ٷ*��t9��\��,\{>e4:���T�����؄��GRWK�ƻ��B�Ǉ4t�<[A���]��@�5]9�qS�<WIӡ���:���]�Ð��eէK�n�)h0���ҳ;��V3�Q��i��҃�)�]�"�ԛ�k$��g4����F��Ҟ+h��`��o�l]�f�YO�2�y�R�;{��K��qN�]4V�d��$�+��-�"�Ĝ�w{�F&�r�v �5zh�n0�:Su>����� [D�Mɖ���I��l���A�u��Zpv�V�s���8C��ڹ���8�����vOfF�O4L��e��c��KO�C�,QN`]���Q㧿]�e���[����$���d�|�U��A:�y��/53�
fK�YӤ��	�Cݎ�),jm-�{�t�:���̚�^਌�tv����KF�.t�ͮF�����������Ŋ�ȦXTD�!U �QQ"�PRA��( ��2	(��V(��"(
�\�E0 �,EX�,X����ea1�	�,���Z��,U
b�V*,�I\V�H��0�`a"�+�-b�
)"�!"8`[B��
H��b��[@�&L���En�៍g����:nF�����2���0E�]*Ҫ���Qh�Y)����s�Z�P��N?O�x�x�,6�����ݗ8�W��:zG~��pX���oN��7�9
��F��	y�*	n/ZIY�ɰ�ƈo�e|]��",s.�����iW��T2,�.u�_4��y.Ĥ�ނ|�r�Q2ǼǦ�"�J�=q���k�''��z���]�UG���閠hS�o�4�4���������|8�>>5�N9�<h��ׂP��W�0!n��*b�KWyI�:}��{�hWJ5�](I򎦟���c���U��㼺�[���F�]O}h��$u���Tl��8�/
��mP�I��6�~���5P<�u��C)�V
�)q
�Ʈ����p\����\C�U��_�>/�4G7���辔��<)17�.�u��(�@�X�0��"*"�ԫX�PV�*Pӯ{�%G���ی�����r��L].-�b���M�jW����������̵ſ�| �
�{�8/��L��4�gT�b�p#|�˼���Z��Ot�i�E�^�p�x�5>�\L鞷�g�Fh�2�C��s���fy����C�3X=Zn��!~�l�9Obӧy^{e����� �+����>�kW�u@�"<N����n�t��U���L"��U�K�yy�[E�-i�<�� �l\*��{�bvd����+&�5�\l�`:�/�i`��M��Ӵ�y�{������jTB=�4�*�1$l�TDԌә���T|��S_�����%��#��6�n�f���^S�	��CZ�!�^K��X�g��+)>��J��7ɿs�a�>�N���2�#���_��T+_�<E�=��?��*��"�b�ٕQ@S�2��MY���n��쬥�V��G��XX�
��&���[�x!��3I������_r2������	P'�぀�SZ��2���� W�*87ο;ʞ�)�j��F���9��A}A���M�=�+�U�N
�0uܭ�R�	UJ�˦n�3GN��%?z���:����<-W��I/pS_-$���$V%�s>8�髊�k��go��1y�,�Ǎ��G�ǥ1��~���^/��;T{�Z�f�|�3��>"���r
tzLXVU,�������yv��{&�]����ǵo�"�o����ֆ�U��nH�m��N��yK�P�:�{泌e�y���1���ķ�S�X*$�`'n�l�kIr����ژ�ب�M��>#��^����t��}KŜ�6f�b�B�M�B��*K��������Ebˣ=���UkXxhv�Һ�+Pp����K�{�#��k�ȝ#�F�`���	F�:�SR�-d��ڰ#'?���/qU��6�2Q}�${�p�N-ҹLˋ@c�ٓ�د�t�ؐΙ��?+꯾��2߽F���B�T Y���3�]�%�nu�P�gq��%�)6��FO{�x�-/�����h\���ͼ�g�|�Mx��`�H�׼�h�����E��Yq}����ب$%��{3Nh�c����g�e*U��]�h����~,X���N����E-8jךϟ}k�<��2X�h�<�C�`��u�g�R4E�њA�<�/����v����t�_��A��RO�`p���ˋO��S�)�S�h\t������q���&-m��Ƿ�y��4��q֔pW1W2Wm�sw|2}�H�0��J�Xk|��~�t��)����ͿOU���q�1�9���VxϮ�=�Z$W�Ze�ٵ��K�抱*н�'\����G�ܑ��t1��`f��3J�g{%_Y��_��V^Y�c43���3d#Od�1^[;��Z�9q��S���������䣞do��,�lC�M\{���q�����J�����}g��@�[�SB�J��w5�����c�K��6��s���R�x�d�u�����C�N*��C���s��xrt�TvZ'ވ��/�XE�3��<D�K��ia�!GO��ӷ���Gw{��\n+��Վ�AS��30w���S��:���Rpƹ�����^�=��p����Y\}
x�"����E��6�Ww=�\�knb�zq���X�..�/E�l��h-!N�-�f)yٻ�aђH��<�;u�u�L�z��U<Hl��osn���d8���Y���Z�
`���=�����w��j�c��s�����Y�7��x���sX�q�S!�.=���+��>�
�G>���՛|y���67�Y�]9dH�1⸳n��[o'J�o�d;/-R���]��Z'ly*	ؔ��B��a��_���x�����{}�q�(�g����^�'�GSy}(S�t*1V����q���Aj��g�h�t_ְ��8�!�g/R�=r���`� ��8�<N"t�t�t���x��^gN��n{�OV� JTG��_�|�"aV���D�ɂ�n�L�� ����y]A�[�S��B���׀w��8;G�ռQ&�p��?x�9��aGm�2�׍�)�!�u��Z����;��5��\��@P�~U��Vnf���(M�x��U=>��ƣ��6��Q!dv���^#Yx��>�@��4�җ+hf�����f�]��`��)�<Ӕ���{xoVu���V�.��ׄ�h:X�ߥ�LV3��������EX	�����&��)�0y���#�˳G��rpn*���o�gC�r�����
�О�[�M�;�Y�����S�X�\���M&�72��u3���}t�v8�0S�b���u)�T���w���n�,E�C�>��Z��cf����Ok�6���D��lU	�ō���&|��K�=i
�a�Q���2_����,��6h"� x��ln*�B�5z��9�G~+\��C/�ʔ%>��]e��Q�ݾ�=�ҽ��1xjӿ0Ŷ���kZXsR6I�4}��dnuv{�Gy�U���d��i��H�H竁"u׷3xq6I	��(5gL���iT-���0j�d-z��}WYy찫�D<5U�����ML�({���d�f�=�<ߨ
�u�ſ*"��G�&��a�9l��C��]���1չ샩�7�{
U�Qj�f�;�5:ι���㡹���36u��3u1���P����݅��!�9Am��e���W��G���6ݸ:����ʪU�{,gX5�;�+�y�G#P/[b����q�/��r�v�	#�5����8;�'b�m�B��(�=�C�m,_um٣�2����)��\xm�Ma%�1����DsǼ���VS$�V��$�=j�@����p����%-;�����z�њ�o�U#ޫ����V��8E���B�td5��8Lw�>d�-`KdRW5/.\`�y oZ7�"�|F����?RΩk�羽�
�i��������NjI6;^���o���g�u�փN�ک.ȱ����7����D�֎�*�u�5�{����p���8��i
<x���6��� ��`��7G{I�,�}�hk�p[}���H�՗)�F�@���m�a۠ɱ��SĠז�St�7&EVJ��?��Ql����<��7͡p������^oT${�i@���l ӋO�^�Vy�K���q�xۧ��J���I� ��Z# ���!�}�H�������}���O;�t�{y7��Tn�*ۖ�;v��<��1�˖/=�$�9Ǌ�������h��L��pZ�����LL+��^t� D�S 8���r6E�0��C��<{����!��_ׂW3Ր��p ��}b}�(�,�u�i*���:m�]������/!p�|=J�O���/������c1wS�_�{�L�߰�|�>V��Hrx�p�ʬ��.���ҩ7�BQ�hZ�Z���7��J�֐Α�o���0�A�f�&A�N��`W�~1ָ�͌i&���P����]c�#�Awj_�%�^%P\+����˄g=��Д;Gu���4�(�]�ҝ�(�B����W�}q[��y�3UJ'L%�v���V�r��6�B(S��%'(Ht�,�d)O?{�]�bH��h�CKj�dDw�;2���҈�C|�H���1�g.5,y�h�]G�b)Lz�/{�L�f���@����Ϗj4ׁK9c�Z��
��^�
���U����I� ��F�X�C��S#�w�n����{�D<w�Kqzh�����z�5��{�H�$ú���pX^��#��$e���E����]�t��|V�^{�e/m�K�
�8���'N_i�}ei��E�tp��������*u����*��򜉄q�\kw.�*�(�Y���fܹ�}0�vz��8���A�)�z�\lr�Gc�{k/�}�ǹZ^>?P?O:�aGz�#o�VS��c�(n�K���٧�x��
*��h�ү.0[�q�&�C1+{5�#K*2{M4i�)��=�[p\����y7)9
#QL�ڜnt�m��Ŋ�����6�@�n#t�7��.�Y�ɕ��պ���m�[j����F�w�9M��-aǲ�v�LU�F���>�*{��:�����r��}'M�yyf�nؔ	�-6�p{���&�\��<�;�nVQe;�0p��#cXx.�UMU������^<=OA����n�K2�6��}�X(���|XY.�.Q����	̱���ۍcZO��h�;ԋ���(~ͼM�=#�����U�1�u�仳>V�#L�#D�Ӌve�K�+z�����r,�@�|+w�"1B�T�rVt<�X��,����tE0|� ���h�S��_:��l8�+������ü�MSK�\�۹�>hM�Z�� ���<�D�e+��2j��wo�iW:an����Y���G{j���V�&�d�zTǛ,��U����]�ƪ����¯�>����Vi� &m�WCs"ۑ2^�]WO�Qwm��S �3Y}��ٖM�1�MA�&���i�5�6R��Ύ��
[W�D�<T��:�"���ZE;�=\8�X����BFm5�����e���IҐ�r���8�v936�豷�c;����J3[l�X��ά�.�+(�/1'��N���	��ʨ���� ,h�h�a>���bj��ʎ��x�C�G�c�X����Ć��X��Oa�݂�$4�<�S��ͽ9�_�	N3gUm�.N�@b<���ġũ�L��p;&��(�\�[���w�,) ���#:an�#;�.����DNٳ[�Tq�K�|���6�%`V(�aP�,���
�a��P�T�d� �B|���Y5��$X"(6�X�e�d0�
T%B�kLل3i�)XT
��*T��+`�)�Z�$� �Y0��cB��RV,�m�n0B�iX�J��# �`6ʅř`e��I��@����/9O�����Ѷ���ΔK7�+s��y]�>79�V����|�w�[m�s�*����<�*�U�-W��Co���8e���g�n��!�^=�w�����QD���g΃�/<t���7�#N�,E�u���Z����VѲ8�ק��q����br�|E�,E�����x��`1HS�H�MҾ
y���ox(l�'��䅑]�޷g�1���s��1��G�����	�.�z��
�R��Bua�."R�_1��j�%c�f�n��C��!`AR�Q9���/!�'������:|XhaӦ���������=u���Z�HLb�ƾ����<�膞k�z�E�K�:�mb�r�^��,[ѱdd*^m�w%����'�^�ť�5#B�!��ע�V�v��:Ses�m)3����ֳu����n&b���QcU����LU�]�:�|���ŭ��ꙓ���n�79��IG6vĤ��^�
�q�8G�֒��0�.!���$VR�6�O��ݪ�wZMw��Ť�x���3R�J��g��V(7۞�l�{{���\�Cت��y����b�9=��e)��P�%��ު��%*�>�w�n��ԅ��C��D徯꺱k�Yٻ�w��ό��$��yٻ�R��U�r�Q�EC��C�N�}��!+��W�������N�/����������v\��,>�8F;�ּDŸ���~������x<J��&Z���0��K�c������"�x����dhΊ0Fӭ�wT/�wth���yx�KN���^(ݺ��n�VE������O�"��FA��V=>�>�7B�Z|�e�0��la#�k"�Ӛ=�{�\#��vIe��ipa|5G{�x��YSZs"�W�o��P��i3���Α���ծK]�p��v�ť�$����W�hv��WE����������e1�}.��~RU���$%���?A�|����7�n"J��0�t��裎}U��5�׵�o�;��1ׄ��A;��YyT���<SZ��]�x����a�!T�|x�Hi$iі���geD�L]8�>s�C���<5��M8��*kE?0�qӆ�����Z:I�#�U�F�a�(Е�3������ؓ�t陛ร��'Q#�Zch�K�Xw�k^��`����pp�P���/Ș=�8�<g�r��f��	Wqi��t�R��Z�U�ǋ������=˩i��(�]^�}J�����>
=*s����>��t�W�O׋��&<<���BV3��*��#�� �?��co۷�M��t�K�F�l�Gfv�������p��G!T�+j��U��0�62nW�Ħ��&x�7꿪��U�>3���i.;!�c������VEt�k{��g�Q��벴�I"����Y>6���?y���@ѣ�jr�6�'`Ҿ�֫�A֌��9UB2���#����=^4邼��V���8f�����X�X{huI}?/���C�̔���!C8����:��@��YH�r�Z�_����.!�1�oGa!F���~E۬��A���oqN$�n�7UT������ψ��_�
�7�ڼ렲qQ4%ϰs���m���GnP>���:î;�|��94��ЀKG�?���w�lu0אp��7�����|G�<X�^/֑���H�G�DCg�ڶj�W�D)�n+�	����3&f�V�s(-ͮ��>t	�� 2���i�#5��]�A�����WK����3C.�@��%J3�t�;��/�*rri9�)+3+�X�sʻ��WN0�':f���r�>�+*��{��p��/}�>C�F�0��6��Ț'n�O��h��ZNu}�����c�-3V��_��Z�\b;�J��߷�)Z���Z��ϵ|�ӝL0��Ը��1��X}�+�~���CA�����j�37�E^GP4 ���I��6�g�{�V��Do ϺޟP��o��"�7�uC�5cNb=�j9ӗ%#�j�#1�}ώ����/�k����'��[�:���S����E��pØ���i�SPHU���I����8����� ��Ի̣v:�V������
v�uu{��K�͇��:�ص+0%��
Ϲi�"�ů�q���Gy�Fi$;,��Uְ7�ނ���nemq��8Z�s:j���d)���Ã(C�d��k4�g8n�!K�nf_V�B��b�pP�U1F�-�oo{^�9cX$,Q�TCX�����!.s�e�{���Tp���hkN���/yq��l���srrJ��ϰu��Z�WO��/��%��Y'�4&�.���x!�3�<��Ť&�˦�ń��֌�q�s�Gy��H�!�IYn1�^!�i'�La��(}��9�r���]*��G��yu|9����ig��f�%�:�aI��֮kĦ�*�������m���xU	j��ұ_G��6�����MtÕ�>�F{^y/��YC�[M���}�iXس+���n��k��o;0]�^--4��^��s\c��]]R��yك5�w�c��>�	Ҏv�
�c5�P�b��Ը��2�P�r1�sc�%����9Cr��/wsFJs@�n�ܰ�k�:��:�5l�:��K�Ī��������X��6$:�)�yk�$�l��l����uk��-],+a������Szק���1�52|���ZI�!��,=�d�Ӹ��U���Z�!�x�$��o�\���(׾ǆ�.P�ڥ(��;�Ok-1��gs#�E���f��H�����܊��m����ȧ�̖����%���F/R6�E�E�-Jᰨ_n]�z��o�󲇺C��{G�
��R��[s�0��#�l���C��q���������'����Yf�z3��g�u������6=��}�-�C�/�)<�����h�����(���x�x<�y���?x兏�ˍ
�ATie����z��ܥv1����P��Y�-]b[#P�5(s� �Q���t���fTߦ�Z�ԌYa(�P��E]<���}W��yשqA�V$��/ʳ���u�����c�quO��|UAS�:�1�6�3Kv�vx%��pw��fv��n��ߞ�O��;VRN?U�����x�7��^��1�
�o���{4^0�G9����xo-Q�u�:I�Q�]خM����
���=�)���-�w�,����Ru��Y2b�%�
��o=�J᫰呠��Y~R�c���c���>I��}�T�wr���c*l�P�V諧�g���X�2��k�[XM�d��.�C� 3�
���i����ܽ�"V�3�]}��Q��JhƨE�,E�r�bK.��w�U�X�+���o�Ķh&с(��fd2J�/����g�h�Ny�.��4)^�f�.��3�0����_<�}ۦmCUu{���~���Iѣ֏�Xy���Ӳ��A�2�6�^צ�	����`�g�M�o��`�G����Xs�w��:$���$�|�w�=遫�s���˓����MI�l�w��K73Y�y���c�X\0�[��ӳv�==���	�4ұ�밞�cn���Z�.�'Q��z՝Ky�5��[��.�6s��zM#�j���ky�� yr5�H�E�o!E�H�r͟�E��@����%in��+C�T���3!���!},��1>�!��.+JU��*�J�����lc��I;^�P�.�s)�ئN<㋁S77 ]t�+h����toT-@��A�L��rN;�W�N�J���k��o/Epw���*�[��o��li�_��Wc�nQ���sޤg�96,�<���øւ���>�����3�m����F9R�R����ƅ���k�����W{�w� ��K�sv�t����鮥3�QN��D�~9s=3��~n��KAW]�a�×��ɾ���.5'���&��_W�	��fno���>{�U�F2,��V��}�LC��H5�/t�ʮ�RX�%�i7�`�xuh1V�k7���V;�o,,T���)؆+JhϦPB�V���X��tF�����Oi����94s��I�V):�S>�2pܧ�&p�c'K���E��ۜ�(�cm��(�w��v��%m�9��6h8��q*�!9�e����.���aL	��:U �T0��XިQ�t��pk4���	Εe�+��s"���g�7 v�Xm��
�ӟl�軔s6��1�N���룽Z�ް["B�9�'�H�pŔ�����Y�Z����T�Z��ȳ6v�JZ�$�L��q�`����УA����]����WQ$]�s�l�I�o�g�ݡ�'���,�pr���������٧1U���ס0�s]�)z�^K|�6:�o7�,���V���4��R�E�0���W�G͒=J�u֬*V�Ⱥ�p],R�P�Pܶ����o�3l��㉂b���Ep��J�����F�׷[F�I'7:t��ڛn�Z��$>�*�8;�n��2�z��Mr{9 ZK��KY��o��\ S� ��e�pT!.2��xV�gpu~k+Ug�U���YxUuv����Mn�V@z�r%�f�f�r���-��v�o����)��f��j5��4z���0��Q.�2��r�d�5տ	�8��<�qo��L������rqX�j�yWSVY�s/cz�iA�R7����#ld�('z��867�k9��-GU��Cb'F�%ɬ56�<��7>{ȭȀce)D
s��|�>�*��
�O��e9L.�6��q$�F�co-t�;wnꝪ�j/eE`	[2;.ě�1���qe�-���3{Lw���q2_E��N�V��7J���N�t�i��N˫��u1�L�1|�(��H,��Z��X#QU�b
�(T�m�
V�(�P��m�Q��dUdT*T��R�J¦m"�r��!K@�2ذ�0Y�e�X�F(L��(�a+V�+�[ZE-�����TP-++-j��j
���aYP�a���h��+����x'���#\�N	ʏn��Ѫ��ɼ�� �P�)sZ������M�_�/w��1�r��`q�Om���z�Y���c�,X!>Z��#�l����Y���^� �;�{U�y�Y�߼�b{���Z���)D��O�����{�W��
��s���\.�Z����ۀ�^ �\�M]���T��}�'4���I���D�}�D�N��vx�S={��M�L��|��K
�j���dsՙ��0�_�l������U�����g��t�y�a�^8*C�;�}�b��ʰr��'��1�=�}��4�>�5�/}��pf��&�V���W��GI������Tࢌ�B7˒^�4wWx"eQ+��^��ؒ�4�,��dK�����	�U�E�r�?�J�t����Q%�?o=���U������H+J;�T}���8g&8ֆ�]�&Q���>�y߸&�r]����myW���x|�PuAt�y�"��Ea�N��Vw��cZ쒞���rVi��P�!{�V{��1�ָg�=�Ѹ�}�o.G�E��y;��m:�)Զe�Pf�����ٓY��y�X�߃����弤1mFC�v�>�k�&�ڊ��Ɠ��,��E��/�g?��5�����˛�t�W��h�W�g�u��+5�{�����y�I^�,OPgN�A��~ш����N:W������������'G������2�J�%r�Gt�\�9i$� �ҩ�����x�.ܞ���8�i�t�����Rz��nVJej(���}�{RϽ,�I]��呬b�6�~�H�=�W,����1�+O�5OL���5���i��C�W���y^����y�����4��}����t��3�~�����[J�9�[Y�X�B�N�l�7OigJ��HԂ�	�m���3��,ok�$�6���^��������M'���r�[%@��e�w��#��D,�dZ7w�z'�y*C<�GV��1\屾�eƢ{��U���-^ڭF.�e]�Ѷ�����H]{V���"k�9��}a�����������M|�`Q����b����Ҷ_rm�miLti�Ҭ�Tq_���9�h�TH�q�������˯Lo,���%گ�y�Qm@��[�d��v`.�=2���N�����b��z��e��x�I��K�7�tŕ�Y��N/�0yۑx��sp.�]�{t���8�Q�M����xE�s�䝟��Cd������y��$�w��]��'=��"ŗ�RH+��������C8�fg���4;��2I��q�dVUY���x)Ke{g���m(*������I{��YUP<uV�J�t3W:�V����%ŕ������	����ݹg���ݙ̺-4���fϜ��\F'��N�p��;@���J;�5�}�����䤳��U���V��<{u	l��"��Q�]+gg��y7�_��ݐ�nK�T�Z��@A��`gOwaV��2�w|Zun�'��{���ȯ!ϧ���z{&�)%�ɸF|�^׳�����M��f�6ۃ�|��0�>:�whG���eU�ؿ���H3jw�k�y��ſ/.OwhA&v鑏@+J�DIcܳ�ƶ�*xvhK�b{���JCe�q����y��I�6Ώ<�g�N�wK�����ZP^���V�����I�ʛ�dԪ��4^wWZo����A�A�]Ҫ�G����gS�70l����+5�Mi��\ckv�u7ʰl�E��3-�
�3�q9#��kԐ�{Q�]s�W����9��3�ϼ�-�O�z��vR���1eV���Ni��D����bK�]}ʯ�4����_�tX�j���(�.*	PР���8�*~���d#��{��gMߥn{���SY-B���J$����Έr�.ػ�o���k�3Gx�ɐ)ih�F��y����������p*��c����������u�R�53�G
b���y�!�}ʽ�������=.J�LW���yo�
*��76l����Z|h��y��3�Λ�x�7����<���!;U�o�a�`Ь_ˮ����y+���?d��ҊNW���ҺjX�s"Z���0�}�FVM���!;��
-E8�zk_}��Y���z��o3��/td�)I�[���s�:�E���,mѳ���RV��o��uV��Z��2�Q�B;�P'&�Rl��ﺎc��lX��|���X:�jj⦼���[ZX�1���S�)��{��^��J�޵JmL�E�EO�>��5�}��7~��������՞M�A����l������aS���x��/zz��`�\�O��P����������OgT	p���%�(���;�z���ae�6�Ѹ�]�M�-}��*�z��릐ɞ�Y��m���5F9�AЬ4�L����;�kD��:����v�|�����u�RM�mF�p������Q���"qL�����e���G6=��!�QR{i �*�i�w՛���sI?�K��y���w�ȅ���Wi��NSeu���P��,�Ƚ(�M�+f�>P�v������I���s>�{��G^�����^����p�ݥ�]zf��3Nj`�\�����N�{���.��@��h���p<�,{������^�?�+}p�m��+�$�W�F9"*z��M�{{�̘��4�AR�]�����Ϥ�;��z�djwlhfl����{�M����P��ۆv>����W��^�r(yU�O:�2U�8�k\���_�l��Q윅��8+w��H�L���B'G��q���R#62�fj0衷F+�[����j	�l_����N�5X7ʴ��,s��[��o%Ԡ��ܶp�%�Q�~E�q��]�Au�I�vmMh��������m����}������X�N���̧��՞��L�k��^{+���C�q���
�ߏk�&8c�Z��mX�󛊨�F�_e���
�B�^4�j�Ob��uk��vW
~�3a��]+>(�J��UZ�Cr�7�^��f.���U �֋9]��K��^��N5*���+�bXe�y��!S~m�8����ӹ<ѹ��Z%Ć&f=C��]�(T�x���54죨ӈ��պU!��Q-r�X(�$��Ԓ������F��蔘_<���o=칻n�2�pߨ��f�%N
�����?j`ro�}UY5�P)�������|�$y����=j?L�,�u�U�9����R׳J1��L�c���YB�����w��9��=�H3 O�������s��࠱��8�6�ݝwQ�U~�v�ӒF�����C����u>�?O�����uNie��s����[���r���Z~��;pj��h��^h~º(�!�q������p������
����w�k�ϰ���zicz�[W�*��4�������^g���M������R��ג!��w���V.+�)�M�/6hWtuKxJ	��^�}�鶮dڌpF��<��3t1sbɗ�
�pI�.�7��R��y���dr��H_c�s+��]�s�η��)8�v� l*c]n/8GcDٰR��21�Ь�|+i�o�Z��֚�4\R��\�їm;��y��,*f� �F�O����ؙ��A۽� 0�\i^�K����ȴ��MS�;���#˖#}jŦ����+����H�;���,�,F�k�f���ś&:g�jl��I�=G+�#��5�j/\ a��a��d�&Z��`��} �Be�Z�Qv:� �8^k��YŽWg�����1�$(���[M����m�g�Yk�vGȾ2B3A&�E�k�{/���������ص�mL�]�nf[���qЕk�P��P�����M�a�\uTglɲ�L� ���B���Z���S�Շ���1򧺸�5w9U��Ύ͛�)�*�i��0Y��3�j�u�,b��VU�X���k�%��݀�B��N8�8S�9H�b�5�.��W�C�>⭻1Vg&�l���6��y�1�e�j��\��to%d�*��M�A6������pi�V�2�N9u�{DWp*�qpb3|�>�Atv�Wՠ�Nx��1��V�&]���R�����gx�̥ɍ�X*��#��%_s٥`u˅�����e��M]�v���'q��5�Ť@p�'�`��X��l��ST{�T6$�f�.8��Ϗ膩��&���g5*���q�\�Q����a�;;����Ѓ235�bޜ�(�����D�|���G��M�r�!�t5#��ru�ܻs:DFS@X���w���u���`��[Ab�d۷+r�*�"�*��*(�U+b.)dFa�X(*�YX*�n)T+F
,A�UJ��Z#�E���-8R�f,Æa��EC6��Qp�W6�UUV��(�UUQ+k*�Ab����s�
 �F"8����*���88|+�ӥC��Z��ocj�CRt���T�fg!Ϥ �v��8[����U�Վ��0l���hGנb�,v��d�d���}��k�L�y�CӧW_{���gg��Uce�,�e_*��-���_<�>��$�{���2`o��O���_��fDM�*`���7p���iw���c�+��s[��+�r��Q7��ڿ�o�?�Ԃ��I���:0}��G�;���*���fV�_�����&�`��=�g^��D������)w�B���RhL�����TΚvZ�/�ڲ�lOh��~���nG�z��WF��֩�J�-Y�X�^����bl����.�w���h�"�8�,�>W����r�od����+�zD��y�0��9����"tw�۔�6B	�[�D�d�����Ӂ]����~��GM�Ofy(�>�U�?];=�V�:7h��%N�-��
��������֣���	}�z���Z��!��l�u2g���d��v���`m�)�|P�Ô|Z���M���r���9�g����ez�15�x����Ԡa�/���c��Bȯ%]^��)h��f�8K3�n�f{�^��zs)���V�J�炑��5�M^og�Z�T���Ũ�-I��o>R�ܺ�[+�F���y�rL4��b������:lv�o-R�W���|]��iOze��Q�x��"��&��dc��r�lU:]�U�k��wE2_&rT����#5��͇-�o�-��=/����Y��}�FK������j��V�wM�Q�W��&6wfR�U�w�Fyܑx��si�qzޒ�B`ښ��^�0�Ώ�u(]�%v.�L��H7o��}Fg�]u>��m�ʻ���\P7�Տ�j5ʼ�S������a�$�7ڡ��im�ʫ#x��mm#�ˏ�M4�}�s�h�b������Kow3ڣnBtܷ�5�=�6m�R���ʩd���x�F	ƴ/s�jV8<��޿�a�j�ne�,Vy�v/&Tg0`���R�2�u�(�B��1�:x��{_>���wt굔7t�ͬ<�yk{�Z��X߈L��N��[VϜ�wʬ(�;�I�GG1�wy��}�v�Ѩ2��	uy�X�~�W�L�L����@v�V�L@���{A�N���\�����u~��w�+�ʤ�\�=��m�n(��6	�%#�4@�TȻ�ļ�go�Z��-?H�U�{b)���{>���W��F4�{]$ ��h�Z�0d�{p����8fiU��&��wiK��)�|�gm�D�eYg��>b��20��;�(���}������h�+�2�8����z����ȞNQ���ں�jƳ�l���e9����٤��>̡\��{�~(|��j�v�_�ؒ6�s�Y�U:��R��B\):�WZ�p��������6�z�泠�)'<�I+i�\�jm;�q�G{'.�Mol�)���:L��³�7՛�oU�kòwz��ːtQ)���)��|uzz�֏KO&�P+�Z�C��Gi;�]�`�wq�T�������r쫶+��4?`���Լ��u�S�Q�̆z]�Q�+��tv�R���k|��F9N��g��ʵ���%�e�����k��+�Mp�X#�=1��%-�sw8��.!��:SY����Md�1w���ُT{�A�|��=x��z�t�Kkճ5�{�3/J����Cܩ�VD�o��X�>���$G�<�+�~�44����q;N�֣̈́ۑt�o>|kz�^��k7��x�j��NH�.bNiG$�%�=
�<?3���g��"�V��A��b���y	���3�{����?.(A���g���^*f�s�Y�m��s �$��T1g�e����R��R���6�%N�G���Wt�Fn����u���W��#�����7WүOܼ������§ce�E�M+���*﷑"Ռ�����m��\��롭d��eb�q�T�rΙ8���(�����2g<vWq�����C-�~\�l�졗�࡯p�&T�lV�0�p˘|-�@�SWoS���[�%k�9kꀊ���]��G0�u9��2��ԃ7�)Q��u�*���v���jl�jW���m��ۛ���v�=g)R���f<�`��仴��첆ae8*�{�'y�*���,��{P�.~~�y'�9ޱ���{�Ug<سm��]Ԛ�E��M1�����,���]�����B��\�=!�fч{V��}��!o[!�`[[�M�.���F7F	���^�X�L�|ߧ(��b2jHx���# >̭Q�L�1�"�M��4^ސn��(�}dsg<Nޕܜϓy��v�#�4�6��1�(�L�]��c�}��fg0�����=�˱y�G����p�9v���|�&ks�یܺ��*�x�!�;�����(����q�]���{Q=-��՛;\f�֩�]qw��]2�d/L��2�D�j��-��I=�D·�L���VF1�C;�x��ޠ}tEl�ϋ���z��I1g����������⩃�<\ݦ�2�o��EĠ���<��i�;��T<"�O��&
&W_�/�y�Ձ��s��㭬�n@ꐃb�@!]W�#��^g�t�&��Tb�e�J�����g�xү�%�)(}�63~;�H2N����[���2Q�S�CЭ�-�o�܃��f1EOMڼwKՎ���ixGo��<=���4Sd�K���٢�ñ�돭Py����ܮ(��"2h::��
�L�4�*X|�O3��:���Fi_�r��t�ƬC�Mʾm��aL�ǭ@ʞ�o}���_�+�3J�B�o;�c���齊Nک���+���}�Q+�$��7��.|�PX�#;ڞ9���|YB�jmQ�6f�}�����<��'�&v}������L9�/|�J�5CwJ?}H����ir��\�G���2��X�>�eg�o�;�잶��]����\=�$����/%A��������z1I����$�����ڞ&�;�)�w�p��O|�4T	��#4Og�zm�_�E=���Upe�8��On���~Z����O��qe��2���R��-�>��,^��6�0�����Fxь�'�`�����"Il�%	�uH���)�N�2u��NĆh3K�m���j���2���~��U��Ѩ6W�ݣ�үa5v�G�%�}�n��Rז%O>^�<4��Y���5�wNޒOP���9��+v�}y�#�������j�')�Y�</��Wא�ѣ{�g�0cfp���~��^��Ec�H�ܘ�9��`����G������;�箻���C�����#��dg�:�f֨t�>f,�44�t�Fn���VgY�o0�=7���_LͼboW�����������"�X�Q_߅�d$��m?��$��=>�k$�"L�IQJ��|b�/v���l�Bѕgoi��ْc6[�Mx��"$E(�$��H�Z�"AU$�$Q��T����EbS
K��D�!���(~#3��Hb1�ۭ�E�D�w�*��h��
�X����܍��.l6�O��R�90�Ւ�΢Q|�52F��զ�X����L
R{7տI����w��>Ɠ#M�I����wn_��&�}D��@뀒!�*M		"�:�*��]�:��e��:��O�2z�ĳ���v?i�`�7�ĕgo��D�j>r=����9))Jq"懭R.�0�jd�i.K3�k��LP�V�{VazH��QkyW�IF::\���
4�ޞ�l�g/y]�O�H�
jp��d�ƻ��R���5)�$��;���I&��UT�����7,ҡk�1��դ�Y�~���7<�$C|���R��K:fgt8��>�C���{��Z��__��Z`�=�S��mN3��ͬ=���=�s���#?�������!�䴕6/��F�nH�˜8|�͑g�N|l�l��XЏo%������N�U��&	������_t������{M�I!��������%zOSvSQ�Qu)�=f�YR֑���$�QK�bI!��R{Ȧ������iUdt�2�=�cvI5x���X����Fm�$$�ff:/J*��M����J>MI�Uh	$B�Rai0�
H�uɁ���̩�=�jJ��	�a�{��
K�Z��4�&�r��#�f�H�����w��uH�$�"�^/*Oܤ��3��II�}ۓ�76qnG�6���⋒9���72�W��Wi<�NSg:�\z�/�2�t�Q���,I"D:��t8��^�Z� ����+�I"D-'�~R�K�����q6�Y�ױ8#t�%�����b4�j�iK�=\�^)E�z��ޡ�Hsw�n�3G9x>�����Ɖ��ˊ���7�I"D/�؎�c8�(�WRU����
�Jz4,�Y��86�G]E�nY�fv���2�ǭ0���J��!����2��\xt�]:��w���~G.0D9I����27�om�3��d��C_�xy�|3��*�(�9E>$s�܉����w$S�	��s�