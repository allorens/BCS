BZh91AY&SYdM1�1߀`qc���f� ����b!           �  4    �             
               �S� =�T��=���gl��       6   �                       � z$)%$�T (��E*������H*��U$A%H�P��
E@�E��P�%*E}Ԥ�4 ��������AHgϪ�8T��J��4��Å�
�u��R+��$����B^c*��x6���Ԥ�w$   �Ҫ���Qͨ�c�Pq�{*�[Ҡ�#�����y���g�s�7�mE
�w��%/}@GvW>;�)���>[�mAO-叐iB�   �z@ނ��P�� RB��wUJ�@7c��p�۾�ϸi�Sǘ����J��k/@��ϸ��:*��t�{�gԥ�gc��pu�š�  Sv�*�����f>�t x�<T�<�{�羮A���l ����:�b�����8���gC��5Ety �  ���U
��I���T�(��JQo����ʹ��=�޸�c�����]��x��=P�O 8�{ <^��p q缅I� [^��qi�  ����J��pM��w۫�	[�BxP���4�ޏm���;����$�x dx���ө���.�@h8   ßH�J�V}@U"Q*U
������:P��좜�8�&�8����z {�*����hO�q���)�xl� �   �_( 	p{������t�,M��w1�F�@�PR�:ۇ�{9$;�@  �
���)��B�JJ��V��>|�h��Aް�Sv�ݝ\��v�v�֧�@=�H��tb݃�   ��P��#��Ѝ�eU:�C���=`�u_g���;ފ��O+�b ��@     4    i�0)T�d      <�E%J��0    ��T�L�� &   	�FOd�BU$ @    &�IT��  � T���T�'���M'����@������|>����'섅G҇����x\~�=x{��ׯ�T U�&��"
�����
�g�D� *����$~���'���~�?� *��nUU��  
�FT�,� ������=~�2v\d1�q�Ɍ���&2�2c2cq�a��q�q�1�q�d�N2c0�.2c2c'L��L`1��\e���q�`1�eƙq�q�q�q��1���ˌ8ˌ8ˌ8�L��e�\a�1��c	�=2�&2�2c&71�z`�d�d�I�e�La�Le�La�Le��0�'L8Ɍ��c.33�8ˌ2���Ɍ�$Ɍ��c2�!����c/q�q��g�8ˌ��q�l`8�c)�8ˌ�A�8Ì8Ɍ8Ì8�Ęq�q�q�q�q��N2cL8Ɍ8Ɍ�Ìq�e�N�q�q�q��Ì=0c0�.2c2c=3�e�Ld�a�La�Lld�q�1�1�1�1�c1�q�q�q�q�Ɍ20�2c.0�ˌˌ�Ɍ�Ɍ�ɍ0�2�&0�0ˌ��&0�2c&0�2c0Lc2c.2q�e�^�1�&1�1�q�1��\a�x8ˌ8ˌ8ˌ8ɌL8ˌ8Ì�Ì8�cc,ˌ�ˌ8ˌ2q��ze�d1�q�ca1��n02cLɌ����Ì�ˌ8Ì8Ì8Ï&2c'L���8Ɍ8Ɍ8�0c/1�q�Ɍ���2ccɌ8��8��8Ɍ�Ì8�(ǃ��2�2�2Ì����&2c0�&0c&0c4��8��8Ɍ�ɌɌɍ�0q�1�1�1�q�a� fAq�\e�P�Dx�2�
�"8�.Q*8��0+��c*L������.0#�
�0+�� ���eG(�C�q�E�q�\eW�	����0 c �0+���*8�Ș�.2����8Ȯ2��(��������ʁ� �.2���� �Ȯ2�J�0�®0 c
0����ʮ0�� c�`W�r�U�$@�q�C鱀C�����D"����8��eS1�� e�@q�d��Tq�aU�U1�\`�&q�eG(��q�d �Qq�fE�q�\d�q�U�Ea@�d�2�c"'L�Ȯ0+���2 c 0TJ2 q�\a � �@�`	�\a@�d�d@��	�
8���&2+���0��L�®0+� ������ �0L0�.2�2�.3�2��Cq�1���`1��\`1��`8Ɍ�2�!��0��c�8ˌ2��<a�\a�\e�\d�8�cL��c.2�Ɍ�!��02c�Ì�ÌɌÌ��2c2�0�0�0�7(�a��q�1�1�1�1��`�d�d�L`�Lg1�1�l`�`�L`�Lg1�`�Lgq��2�L���Ɍ�Ɍ�M��d�La�a��g�`�I���Ӧ2�8^����y��eO��ʹB��;��2�anm犺ɘ��j��l�U�����a5�8�f�0MTl0i��7�h��oG�g7�mu��Ejv�[�K��c^��P
c2�CWx��
�مe���TVhHը���J�C���t3���Јr�v��@��{�YjڼybՀ�]�%��L^��JPt���ېa�v���:Ɣe+�F�3�JB�	%f\�ձͣ�Z��X�\p'��=h1�[��t	��)��7�6lk+-�\{Gn�f����M+n�:�g*Ĵf��Ж�+in����5ɛ*i�U��F�w�fӭ��%��+:D�s`�v�29w��H��8�֨�w1�srF�uT�y�{�yC33X�WV�om���8&��n��6J7F�'DnJ������n�f��G&A������@8ڭ�����<��f�	'����X�,��i�y���+6J��� �6�Ɩm͕d�e��eF�4�T�n5�� 5�^]7��+q�8lGYaAA WN��T���7V,l�˫�ڳ�� �]3��Oe���wW���#S{*��� �V!���\������j���I�"a�QB�wD�fm��w	x�%+���~F��#hi�)m+�wf;yY�s�b:Z�o+�Y��8\V�i;u%`�&V+��1Z`�-:�(<�n[��А��+lѼ*���[���X�n��ҽ�MT���&�#o2`��m�T���G���s6�6m�Gi!z4&Z������sÂ�ٷV�r�X�����Og�]A]�G+^J%,ͼ�V�a����Y0��L��Vb����� *���QN' �>�l(ٺvp�f���[.,lT�U,����+v�c�kR�FNRj���A!h�'o2nz3{Cj������R<�1�n�� ��Y�{-i���6���Uw��
�J\�Z�(l;4o^FSu��r���nE���ͭ)^Z�Q[y-���\ctc�W���-�zf�h�x��h��W���kU��m�HU�[�^,VV!�-c�q�a�p�m56��VHd����w���v

��{�t���Vn�g)j�g$ن�y�u�zwC�-�Cj1[�2Μ�� �@9��ݻ��衻���Rr��L�\�d崮��9�Ycq×��!ex��f�i[t *��
2U��h`ۙg^��5L�e��x�Mq�u2ղ7=]M�;�l��Ֆ�ȷh�0��e�ǯ7F�+U����dw/ ۨpAk4����S*�`��,7Wb�R��K�"",5J5g0m�
���_�.{E�5x3(kp۶@���`���$�����w�w���R�	���[���t�1[����!�ė{�Z)l�7��۽*�b7ud����Z24^U����(��Cd�����V
��㫸���Io]6��S���5���w���w�ySwj�n��6�V��CT�b�B	uu����*�Y�l�ݧ�Uo*(���QV nܽ¦����*���{f�"��{l�Ɯ&�Z�ߙ���lV6�f��en�(��Q��H�&�VnQ�̣��H��cZ�mV�ຶd�$4*[��F1�TSKv{�s-лq6/I��(���CqT!E���e�n�&(*�<��R#q�
�Ql���w3U �I16����Jڒ;hZƬih����7-$��<u�F��ѳA􆬀C�-�щ<S�K��V�"k %��#N�Ȟ�V^��T`��W�������v��)=Gw"KzI7F���@�v�Z���єf��<�u�����2q`�Yn�̉�5$;S@1֤��d�"�z���w��މ�X��X[Rnt�f�͔昨S��y�-��T[�����ap Цf�t%(XQQ��÷� k!z!۸�L$��w7sP.����ٷ�Kb���&;�rj�um�6�U�WJ�n:��iۈ�t֕�iP�Z�ʆ����mJ�t"4�Ty���Û�iK�Ið�וb�*Ӡ:B�r���MFQ��U�	n^�3%J�8Z0�O 7��(]�Xf�˺u���&=�7j9�+�u�,���u�];���4�7A;�n�=�|��ƠpT6��Va���b���y@Ƥ������lJF�n���i�W�`ջ�5��Ä�h�J�+o�xI���E%{[4ل��Ჳf]��Bͣ�����Q �ZEɺV��)^�����d��vV̅,Xj��A6U�NLv`7�����p!�.�v4B!0���I �xsMmm:�NL�@�7�Y���Ƈ�;�2�#>�U�DVT3Fg%c��2M�����Պ)�ڸ�̢�e�J���U�`n�c4c���5j�+e�՚t��ͤN���JU�����S͹�3ۻ�K��n�R��iM�Yw�/X�,X����H��\����ӃVKOr��ku�+7J�=�hSX��[j��<�o��NV,�`V���w�֣�4����4캱y�WV�E�͒�˻�^#b�T̼f۸�Wo4Zoff7kL�{�M�[�������˫�ʕ�	B�T���c\� 9�6�.�g�+$�G]�У��T�ݫۢk̻'A4N�ܛ�n��=�Cn�"�JlRξ[�(�&��4�3�n��w7UKӎ�c+.�a�3C�-лL�d�Y={���s-X����cZܑ�d�ǰS4(��,lf{NDfR��wY.������Q�Ҵ��K���W�k��$G,�7EE�L�/f�+zK��u0ܗ�1���h@��/QʻX\ћ,���.]��Y�͛!��p��Y��Sif��LU�R�/r�������*j��`�4���&5nl��S36c^�Dτ��Z�^em�����t-�t�ĖO�Vm�b0f�ǡ;�x���HJ�w��פf�6v�0K¥�j�i��:�ס�EDڨ2����(��am�(9~�R��N��EbB��bV� m��PɒGF�L��m
�QՑ����&Vm�dx��̫V��1�<5]�$Tݫ�kXY�R��k��Xƅ,q~�yj��)���ekp�������[sUkb�*ŅL�� d�a�v)nQH �O��M��5{5j�[�歠d�1�&�K��R��y� �M%K[x�&�h�3!w���IۃUD7`���q�kT��!��q�Vh����&�o,�)ut�;�rѴ��c�8&�7X��7M����)lM��#
�2Y2P� 	P_��l�Ŝ$1c$�U�rb9R�e�ʩV�apk&%;�`���7^e5y�����.�޽�V#@O7J�v� � �1�V�g��=�s"��;Z-P�Y`ݕ�;˫����h����n�S6�[v��B���i%ͳ7�5a�$4�y�tRU��TQ�n�V���3c�~��IQ'�5�����P���j`Vu�B�oJ�YKT��lV	1[����Zܵv�U`�X.�Y̠n�c�s�7{Z'�v���M�A��.���3���J��əJ�Vݗ������;C!я����4�Zr�v��Ⱥͽ��+�*�-�yY.�4��ĵ�i���A�����[ZF9YXI�Ҭh�5/w)S�5�n�ա/KKsl�(�[�Xr֗P�0ɖݑ�ϥ䧙�;�V���6TM�6������d�x�EDo�]�y�3aj�i�o"Tv�ʊ�AE���=��!o�
��i��``Ʋ��[��T3U4R�E1�F�X�ؽn=�;�q䤊d�n�f]�Th�&Y��"��3F¬�35ޛm��ufj��:[�o�%+0���\i��fܭ�.2�`䔶�i��z/36�v�)���.A��޽���5�ӿ;�_r;��v�G{�{�=޺b���	��&Ս���ΰ��{�_�X;-c2�r��{�P�Kڶ�]j��74Եba��� ��w��Sf-Q]+ǶC��n�x0JU���4d���rSv��lxr+Wh���YI1=�f�X��[�6��6dӠ�O1b��55;��&��]9o72�P���[q��7e-��x��%�=���X�{5�"�s������l�`���������d�svk��0��~����.�����`JP�Z�X��*�.�7+JU�*y�]f[#���B���Y��F��ZLN�܍Ѣ�B�q[��@�+��w�
X�Ja3�Ɓ�R��H�TĬ��J�J6�e�(����o� f!Z�LeixB�݃�:wok˲ff1Of%�*P�E�ZV��H(�^���=���o]1���ލʭ��Pĥ�{{xkkmց����Ohn�d;PR�j,�{�	ء��Z�mjC!�M�0<�n�,��X���Y{�@dLPMZKM�����݂�=[B�Dd���w[e�n���R�`��ݼ����n�a�P
���7LS-�VxNЛ�œ"�6Z�C��ڷtM\��f�<U&�ʴc��cM���U�U���dj�cu
�:�aA^���M���z�+-����,��J�-��f��:e���w3S�Q8n��7�)V"X�i��T%���MJN��&%CUM�q�WR��m^�]n=/,*H6��,PZ���s�ؖi	b�Iyp�Lr%Zz˧Z�bS����*bo'���g��˵z�Vk�
T��@����eu#M�-�sY���ax]���4u*tRr���n�sĬ�Y��V�tF���n�x[ї�R�N;���[U/*�C�����Em�U��6�9r�	)�I��ʲη,ֻt��y�f�6'cj�|1�t�O2�j4��^��V���Dѣ��0b{aS7v�.�b8fܸ��u!xu��.�j�6hV�E-�$��Ȗޫ�b�U˳�vYxN�A�Ur�i;GN^f�t��lY�F�ܫek����E�RcY�Kf��8,6ail�G@k5�GD��"7Af-�&1r�
�����˘�"kv��Ԁ��ݣ�u^�"^j�@�\�Mv�2�]l7�����e�gT��������u�u`��W��*��4�f^Yn�9�.�"�����[~ݛtUM�-��-�G(����z�nY~���)��-
W/�Ƭ~2X���)W��;�I�݂�6���[��E��:=���Ѭfhob�*X`^f�-Co[���ݙ�����f)퇖�#���Jo��[��{Ab�5z�ͥ���)�33dZTr��x7����Yt���m�2�е�3)�@{*�a�f�Y��n�+L,P�̛dZ�gJy/��7ZV�y���Op�����NZ���z�b~�Q"�*�J�U�{����6�7w=.��ۑh 鬥��X��U������.�C�mk��v��t�h��̴]J�Yf������6=p!�T'��J7��3M��wx����؁[�(��4Lz���,:m-�.���<��ta��,�Ͱ��7�̹oP�uD���((ܬX����KrY"N	���JՆ���6��J�������q�v�f�U��ה�1��6�eR�16'u���d�S,���p�-�gtf���u�aj��9�v��X���ִj[[&��ޱt֜�x�<������oDX�Lh�c�'k^;�U����6��T��X��w@ث@�h=��Sת��v%��x�k5�ۆ�r� x���MZ�Q���rV	cf�њ�	��m˔��b�	iݱ�vf	�K��X��B.c�(�P�*R�^VV�;��8+Ea����2��cL�1`�(����wPf�����4]�8�cL�H�7F��۴w+N�7��u�Q�2<Z�`��e p�pե�6�-���$��Ly�+��=�Hd�9{v�3kf	c+h\����u(��œ.��u�Em�Xn:5�7��KMɍ��Jʺ�/S[g���z�U�ƨʳ0:�Ȇ\���Cm-F�G��H.ơF�`�с���ukDw2����r�H.9:�A"�Wͼ:�s36���n����F����2��/��fi�E����%֦/	�[WY�@���خe
f���N,�vH֤�9B�e�i��#^ٕ�>�|w;LW�ͥ���v�YE㉴$�4&�T�|��Q�]p�x��¦����s\��4�r��D����V���8O�z�Y���FwQF�"��t�rdv����(�������l�e�.�ҏ5ִ���w�N�iGcU�����z�ۣo�/��N��TqW2)���Գ���#�3�g������[�8nE�m!�p�\m�Nt/"�\O�Mq�E@��z���/�_�r�W�etzV��f_cW}@Y���HЉtG��9���_vg��9��ǭ�g��?}J��ܯ:uu7��_flg�0ҜQ.W�#l�Г(+t2vVD��tӖ��Q�?^!��Q��f4i�ŷ�.�B�/����\����!̌�wOu}������������M`EX��'��tt�;.��ګ����*Z�0��< @�J,�����f������mG��ݷ��n���H�a�mm��g&Y6oDĺ�Dѥ�uZ{���:�:pf��V�2V�{�PYTm!Gz���f�75Q� ��8�"����%>Kl����pٹe*_ �3�	�x��Hj�<�֝Kq���b��$76�;��6k`X�;x��ӓ`����)�t�'��x�=&%)��vEg՟ o�)e��#)�p��:{�#�>m\�}�[�����΅�=Q�{����]�sn'����!�J;baɧ	�S���%�����7vK9��������Xm���F�˹�U��c?B�1W�I���+�|D�8�+M?��!��pVڐ�E�oTI��|{�t�}mEEG�������sjL2a_a��{����/M�����G]K'bԜ�����K�l����V��m����{1��W��t9��U�O(	y���M�+��K>����ol���3�oY|6I����M�i��ӨFn�����D�i]��(Fvy%��wg+2���%w�O���P��$Ǔ���F������Q���(���ϴ�*��Ʈrg�;���}��z'#*1�fޒQJi�zc֒^X����o�����~P��GsD����`�3~Y 4(� *�*�4��@�B� !@�* RR�H�@���� 4
-*�
H)B�Ш�	H�B�J#J
ҋ@�R*P- �J�B�(ЁJ�#H4%(	@4(�
-% ШP��B"�-�JB��+J*��H�J�У@�J���"R ��P�J
#B!@ Ī�H%(�B�"�HJ��� �B��Ј- �AH�H�B�
�@ RР4�(� � ��?=��^\�ǯxv�}�zoo.֒�B��j�S�i��<�`qͰ��Y^����P_;J����$٫�0V�l
H08obw�^�{�:��$'�e�~�~Vz�2��T��]�@��Ӂ;-d픴�R[�C�ړ�.!��9�p�˧�P'�l�<�
���۰ƨ��hX��1N����O��g�y7�����ۯKގK��%Å�,^���&>��(nP���q�z���J��3J�s���8�ĕ�#_;�=���Φ�Q���C�^�rƷ���	7uU��3�R\I�����ھ�������,��6��%��YOzM�x�CN���6��s�m�m7�=a�N��nU߀lҺ8���!������[|=]����Y-���Vn����g�$<����^0
��x�|~=Uc1����$����Tf�/�=-9�VФe%��n��s���{�j�Z������EP\&�;Ü�y%�]r�5x��ׅªn��k6�ӪA�oN�����\�nu�6�>t��k��7>�]�M���t���i 1��I*��q*�8yA���iY֪��ti\�/��7��K�q%�g{������[�~];;[���ߗN��c��N�}�M)ӧ��a�p�W^��PG������TE>~��}��O�o_�����?�'����8}��;?����������Oj��5���2�2<"��ͽ�zݞ#:�����7p�h/3Nh[{�C�K���z��e7���FŷX���ikU�ĳrV;��u����V�$̏8��ɹ�
u9��wn��n�����W���ɚy�a("��&�(T76]������82�X�.�z
T���~嚵�0�_�PJe�n�������9�6���y�¡�,l5ܦ2�����f��KwA�Cs.��23�L��������G��1�y���0U��^s�FEB�vS6��w7
v}�r�s^�_6s�a��P.��g�em�M4��1RwF���qN+F$V�yN�y7yd�܎q��<�yH��`ր;c�P�YVk+�Z�7;d� ��F�*aB
h�(��="Ւ��v�S�������
3��o�Q�z�fd9����j����be�-��m������5foj�szl����Q�,�L��u�j��43�گbF��u�;��%2���<wj+�ҫv��fDfR��C�-��wj�̺L2xZ��� Q���e��)�E!�DelpPlm�0=<&7�@ݚ���P��y<�w�0rʺ�x�Qdlm"���f���5uι7�n�e*�7j초��&�Tf��+���6�/OOc���_�u�]u��뮺뮺��뮺믧]u�]u㮺뮺��뮺뮺뮎�뮺�n���]u�u�]}:�:뮺뮾::뮺����x�}>�u�^�u�u�]u�_u�]u�^�u㮺�Ӯ�뮾�u�]u�ۮ��뮺믧]u�u�]u���<��߯=Wy�{�+��EM� �������U�~n�u��F������ڴ�t���VSCI�]VY©�lLP	WY���Z���2@2��E���'^�����w9�f��Ү��׋��E�7u8^���Ӻ3��
���oULC:�N{����h�+�:qw�F�'<�C��3����y����7;7L��5V�R�GUU`���2�Nֺ�2pwq��kh[Y�2��r���eJvfI�y�S�6U��R�M������ ��^�C����n���3���C�9����G�@�c��������L��L,n\=��eĖ��;+5���ٔ��<�ǯv�BVS/Q�K3�ne%Zk/6T��T��`��"��!W]{�����K�r��0u�'�2E�����.�.��]�%,�\�b�;���1G�բ������{Kg۪X�$�v��ty2v�+�A5'�sPʯ$r�Wn�mo"0r��kn���W��3y='!��6����*F:�N�h�7�.T�)v�4�.3��f©Ƹ��Vk]�yٲ��{�>�f�66���cqUU,#��Z:Ź��0}�������e#�x�e���̫��U4�*�UbZ�
����^U��`§�*�5��5��dV*����������{_N��:�u�]u׷G]u�]u�뮽:뮺㮺믧]uק]u�]}��:룮�뮺κ뮺�u�]q�]u��]u�_n��N�����}>�O�]u�u�^�u�]u��뮺뮺뮎�뮺�u�]q�]x뮺믎�<u�]u�]u��-������%�!U�ʬP�����@7֫�vM�@	jep���t���u�;ʴwZSPڕ��5�R-���7d�WҸ!zl]�}�M䯭��U*��a2:�>8:�������3*ͼ�P�2�3��Z��҅X�w,�W�{:��k:wD�*�]�Mgh�w�8�-���|O�aD=UXA�ˁfº"�\t�Z;�W,Ĺޑs�ݺ+��L�V�ʇ8���<��S2v����^��K�;.H���ᒕRO�-or$p�'7}B�^Pvh0Zԧ^�sK��|��*�l���L��f��g���U�ӥ;.<�(c���ڙ��r�s��ّ��g*�9kI�t��^FFﳭ���,��^jn�o(oGm�Di ��\Z�l"�vr�u�	�y*`6z�:�1@�̏n��:{Yڮ�8�gd�+컬H��-=]s��J�rocw׆mEL���\D��Y���@�!�JV��ltu��zn*����$�~��>���Yh	�n]��|�+��#�S�dh���ɝYX�R�m�3������ќ�д�F�;�Nv'����N5�uUW�FV� ����:ҥs��L���]u{.Ռ�g2q��/��/���}u
�K
�SۙǗWj�N��c:���x�6�Z�T�q�����)<�]��E����B��U�u[}:�㏡��_u�^�u㮺�:뮺�u�u�]u�]u�u�]u�_n��Ӯ�뮾�u�\u�]zu�]u�ۣ��뮺�ۮ�u�Y�]u�뮽>:뮺����}��o�]{u׎�뮺�u�]q�]x뮺뮽��:뮺믎���]u��]u�_n��뮺뮺�뮺�u׾���փՇ��*���jY�Mee�l��2.u��V'�L�T'2�oe�S�^�뙭�%+�e��~�Z.��qv<@_ve\�t�1�]��di��L*Z�j���a�������Om;�t���T�*OZ�{]XOf���y�P<���&3�4YX�=J��q�E�ܖUn�&����V�0���k��'V�U1kr���ǅ�yCl�<;}���#�U:�j���J�B�@;���$;Y��	����Q�&Uɤ�'C#����W{j���2M.r�ʳ��;aU��Y��x�5�RƄ0op�d�Xz��v�Wԓ<����u_2:�Z�f�t���-p����K#yub�V�r�W�]v����{��$�v6 �O����{ڨ��+LH���Z�i�O �q��Ec��{��vj�a��	y�L%���;F�S5��n�;���<kj�BsqֺP���g���=�[P��~mZ-���R�^�2�o��
�)f��(��3z�$��<��v�	�\�X�a�ɭs��*]>Zj�5�o]
�ćB�~���g���ʠ��˛1�t&�j�
�v��=g�`[���h̽�n�r^#/�����B�kV�xe;Q�v)����]��򩷩�t�쫺ڵ�A�f�!�œV���O��8�|g_u�]u�Y�]u�]}��N��N�뮺�tu�]u�]u��u�]u�]{u׎�뮺�u�]q�]x뮺뮽�:뮺뮺��:뮺믱��}��o�]u�G]u�]u׷]x뮺믧]u�u׎�뮺믌뮺믧]u�u׎�뮺�ۮ��Ӯ���p��"�Æou�ۦt��ٳ{�z�d
o4{����]v� ��y���\ɵ1Y=S��k�Ŭ�	ڬ��vg���l��gv��+tL{�u��9��ޘb;1n��FT�ZÖl\}{�_,��fG�y|p��r)�1�
�gn�s�2�sV�����x�E��vc�(�K���s�ުe��:��� ݭ�fA�N�[y)�sIV8�7�������j��b�X�<i�9�6����;��Q}ٰV���r�+f����VjY��7kXۺYdX�o��۹��f��c���^��t��Y�z��KZ/1U��3�W���=��̱qP�n,v�åu�������K�оn��1B���g�=�z���r��
��@/Ai�����-*��Y��2�o線wou��Qu�v����C�!�;ATf�.�ܒ�
��U�U��<�G����z*n��b�~���Х*"���*ue<��3 T�L&�v����Õ.���ƻ5�5`��&��������1`��ڰoyՁ�����;t���2�!��SIq�l��a.�2���2V���Xf���n�N[ۧ�j�em.�v5�̨��t��;)J�xУݯ=��!��5��wS��f
�>���u�$�nne�^Dc��B�;�GK=a���;�`�����l��In��u\e��N\�cl�ʺ�G�^�T��P�W��O{ƞ��Ǯ��ۖ�<��*���z!ո1
�n�S�^�b��eZHW�����He�;C6� ���v�^���8��o�h�������?{ύs���yp��{��W;x>��ܫR˶���K{*U�7�ǚ�;k��X�9�w,J-Zw�[�֔]����1��`����W�i�Nwu�+V_�ɞN��m�H�w���k*�J�=�!�0P����
ƖR����Π��1�S�3�dٽ9Yʗ�f�/`E�5^��s.X��)��AN]Lxmֈhb�NL=Θ�V��.��v^�f+}���ԫ�*�UlP��3Eo\��w�C�M,;U�9�=���W.=u����#6.Uu��w����[��Nd5C�Y($�.�m�#����5K�e�<���v�݄�o�\�i;�l��/W��Њ)�c����b�%֡�2�V�P�:S���X����;|�K�ua�S#�򡳫�����suۚ��8м�r➪�bѬ��eܛ�\O7�����ˮ1mՊ�Oo79�lS��1�B��ntU#H�u��kh}�z��m��U®C�e+u|&e��G^Y�]#j�fu��>��[�b%g�m�̹�Y�L�gB���|������uυRӴ-VW�4n: �K�=�&�����/0����U��ֺCv�e�WwtvU�V�������.�n�N�Q��34MX�^��}&	O���+ph
��-�
�A{�¥!���ʋbM�Lu�]��TvDgm��,��f��W�|�vwn�m���Gʎ��e;�o�.���ZJ�<��э��nlu�J�,˻އ
��Yc��yB��e��������#<��uN�U�f�Ҋ�$f�i�Vw&gEδU��T1��9g����x��L])�J.ݨ7�k70�UL�T�Wo=���S4ҝ�3�Q=�^sLk�1J�T���pd�w�Vِ>�wj��ys�x%���s��p�9���@�]88�]�ucwͷ(
��gsSԎ�����ٛy73s���|䧫S�!�n���t�.wx�mpzFC���z���/"z�;Mݡ�Ԗ���,��Ϳj�V�_We�P}dܕ
�d 2�f�]�k e\WJ���v7-�72���f� ���N�0P���u�p7TN��Kf�ݽM�ӌ��V��{*��h�L=���ev�Au��s�=㧷�pyhR��d=��s��=�Y�D[��܌{gt�䪌.FWT����Xe�MeL�y�VA.�͋0�TI�t�w�;��9+-�H�x�� ua���*�){��
\�X���X1�%���|�7
�Su�Y�x6�f���� ���ٹ�Z%���;�	]��OM3L4�7��n��cE��;�pKK��a�]m_�����%E	őX����`��B��ƺ�vC7�zu�� a�p�%&k�',u�f��+l�՝�e��n��bT3.f6�x��{K&[�`ݽ@e�|"�5�|tK�4Ԛ�i��.�����c7E�����|nV��YG&P�W��2���O��7�0�*��iE�An��
�ICn�e�n�4��m\Iڼ�[�ovmn�dt�/��sp�aC�O3���<�2�ŕݘf,Ք�N���m�T���9�V`������z�,�����W�=;�̶@Vox���bj��X��ښ�E��n$���rE`�u�]��Y����֖��9�m̈�z�*C->��8���@�0첝Vխ����H�IJfVT�:��6�[���H@�ͪ��S��Et���ӌG�	����	m{U�x���d=�]�gnDy��:�����ץùz��QV0V4�^/���E: `�^�:n��Ö��O��R��k7+7�W���vV�k�MR��
e]���2b���/2���pv�Ɍ��k��p�xv��őbِ���F��� ���;�k��Ή�F����CW0b�n���Q�R�r���mS��Ε�^��36L���Rw �Yw�z��{.Q7�w�2uu��/(ڭu�x�@X�����c��_=�{�W�B�l�,^uJU7��7x�*�2�ﻮ���PW�]��ڏ;�j*��U+�(�:���lD6���t�ܼݷiaVCo��|B�A�G{Gj�]�>]�ܽ���F�#A�o8ceD9���{qT۶�.�v
�Ae;��V'������75��l�m�j���@�6+�����FmӬ�~���2WfF.oqN���ڴ�BhWv�r��vqɠ�Y�ΐ�4p�,�6]0MH ���4�Q����7Xz�h�8��_m�y�Ri���@r������4��"�Q9�ۭ�@���h࡙2�u����s���Ƿڮ��]�;}`���V�e*h���_<�ʹ�|_m�+|%^�vT�7.Ѩg$��'�|&�u�Xq���gB�����xe�K�-j�2��o`Θ�
���d᥸i�=��&�v��y�o���(�����/	N�����E6*��#�)@)[d�Q[�0n���}vo���õ��J���k�[�����v[��Vp=��|��u'�xP���x��j�!�tĩ]��m2�.�6sR5҅*T�;�Yc��<gaV��| �~�˻ܽ�Z�ĸ>�y2�w�g��I���U_���0L��j�㕐�WCo@��wR���k�o!K\���슅�X��.'$�/r�q]3�Q����5�jp�ɽ�mƫo	)��J�Q!�V�P�Hg#�4+ 螮��m�u'Y{:��ٺ�s���c*�Mh�&�{�@��c/�ha�;~�/,Շ|zk�9IvgV7CU��6g��9xn'^,�G��	qoYH�mӲ�d�%�j�;9!��U��zf�@�uի��c��m�]��!;�)>ɧR��ˠ�!��Xկ+1c+zy�ںyM�֞ub:�]t�ݝ�U)�Xi��
Ɋ&�ec-e���gP�r����-�gq9�V�K÷��f̽�	���#6��J�7[.҇
�n����R�P�z�{ȡ�wN��^t��
8e�וW]�[γ�P]w��3��^�շ�N��;��J��/+��f*�U���wGdR__���i�*]tsuv%`I�NS�.��t�S"͜hRzٮ�]fA��V4�E	�F�z�jhu���K9�ֵ���FnU��`��-�t�1%T�xs���[X-�7Rɷ�74�}\a���
x��|�r۠���|�ՋE�,n�1�Ǯ��f�WK�����)$��%�.�M�@<$3�-f��T�͔�t�j���P�*�OB�����p��]��v�뱁'k7m�A�J��m  U�M��_��?����_������OG���� �k=k�3a`·Xbv�f��m�
&�:�?Ԟ}�Ͻ������k�����{���'�r�ɹ���h����g�����k]�R�WL4	FWLeڶ̟�cо�g!��d;5R��z��v�ƨ8��d��U�.��M��L\Б�s���P2��
�uub��ٹQ�T�,�m���8
Si����LQRZG�nn���k,��u���((�\�nfq�%L[Z�1ƃa����,�uk�D��52	��8�i2�xt]�e0�l@���q���!�ۼL��1�Х�`�ɜ�cW�U,�҆��*�Aїk��V��0�h�Ͱ�����׶�gB�7�@������ؐ�Sp0�5kֺ4�9�h���Cmխv2R�4e1���s,Q!k,Y5n����)-l:��]���qa��1�p5G���m\4
�9������Q��2�zԕTbr�Q�FJ����Tٚ�:��*,�6�WcXKv���9%��6kqa����ů2�qj2��Z�1l�����й�M��FX٪E�!f�٥���*�4�gV�3-΄6��\�fE���Լne�b�0�b��!i��.K�Mj풌�e�me�Q�`�\�v�(Fؤ��
�v�u�A���.�ِ�������
Bh;jXf�3.Ъ@2MIjj�1�,G�+�Gi�퍁�w�Q�hnY�f�Gs1�:�s�t�`f��u�b[r�r�#�f��Dڪ�6���:�m��D�(�\R\�҅1��l��Ø�%���-Xr77k�8k�������&n�r�Q�y���t)+aZ�,r�al!z�)6V@.f�v�[u0E�ҕ�C��lrB���a	�W;'M�gd�#���p�5a� ]�&���`�g6[���ٍ2RКe�h�΅`�j� Dƈ��A�.� #�SU��6ś#5��K��m��kI�fP)v�fbG����ܶ۷3qK���
�d5�P%�9�Ĥٵc�5�d�74�VT���2�ܸk���\k,JSE]�b��k56����Yct!�f�:�W�,N�K�����ꐶ]�is�ݛ(�\�a��u*�H���eq �[A��Y��8)M-b �ݪ�{J-��P3)X4�V��mij\�#6����l�55��а��kL$ز��θ�Q+H6ƹ�6���Q���Saٍ�*�^SG�#C69�psu6���pG�=v��ib˨���t$�6�2�3k.�k)]�[���K��f��4M������T���х&{Xb�ŷJ�u�.�Z9B�� ��;q��+xf���L���ڜ��ҹ*WZ��)1T��*�*Ŏ(1�l�YA6 X�+.�ҙ����D�^ɥ&ɨB����[s�)�Sjʤi���Sn�LG5C:˪��K��Ѵ�L��ڛE�.'N�;���
pf�avuP6�Zmt[X�ev�Rcp��0غ�X�m�B&�7V̚���`���9�1,&s[�t���%3 ���f����M��`��z�JF��XZmc��٢�!���٦���{JV��ڶ���ݦ(\k*���EA[�i�f��\�J3<�[����X�Lk���35�n�eIHL�f�B� �6v�v�4�.�i�*'+�)\�B8L� �B��mc��&����	��@�Y�m��1�f%�]WT��M(VbT-��sM(`�[�
�!v*��WY]���РR(Z��Q���B�d�����v�!2��afy��cc�$Gd%%��Ćs*K*�]c�ۅ�Y6!���2����UE�6��D������B&��j�j�3F���UR�Q͍�k�TM��q�����h<X�����k-y�hF�(\����r%�-�hkm�T`Gc))KXfo�P�Y�\��U�]�sv��,��;�h����][ �!��m��E�u�p�����[���4ÝadV�lf��9���2�ۑa���`$$G&�#E���F�Y.d����p�2M7k�j�Y�V�@�9f*� K�f��[f�␃n��=fZ�,�f6�Q�Bam�i�9��F�]�m��6��&�$�Q�2�-cm�	��U&ÉWn^j�X��,���	3��P�u�-�(��-��]i��\�	�P�8�����0"Y�M����16+����5���J��[L�ܧ��܍��+�]��Z�LsF���,fb������pӰG!�eX��hKuq&����XH�V���1�`�r��t6�2�����Pj�ZW5��ܠ�%�gL���B��/�C%�l
�ȥa���i���n��h�Q7at� lXY�]��#�ˬ!	���P��b-R��ef��2���#2.�h���р6fC$�[ni5H�G.��hR�r��@1�x�i�X�T��9�p�,�r���Aj�� 9�9��7��-��#���5�ӂ����M���Ы\찋i��YMm�v��<\�6L�ŁŢ�tt���g*ƁV��j
v�,; �bhBܱ�W3<�iBY���h.\ʹ��[���I�mL�M� �iX1#d�^��(��#�Y��Z�+�Eг�Ƿ��7�E�l�F6QZ�mNn(h��WG̭�#]���3)0F���Ո: \���l����\��vwj#ii3j%�j�c/3LΤG#��tU1a�܊Wi���y���l�F5#[��њZ`ԯ��YI�Fm^fj������m
��;�mL:�pkr�]�%�p;�mn�kdS6*.��T�G6h�H�Ι�Y\����mQqηb,��nn%��.��5���M\��kf����=�����)�EfF�d��P�r�M�Rҭ(!
�s�a�f��ku��W4�W^mb.`$���g��[�6�7���$A�v�]m���^p�֦�kX����4HQ�p4�84�XJ��b
�v��J�3�`X6%j-&6U�V�x𫆑�-�,�f�i]�h�j��,�s!*X��-`��%�D�7����4n6�$���͚��M�16$/�٣F\PX;<"6f�.E�WAQ�a�����ƹ�Z�kH�dø���-�^����]E��Yn�h`�95q2BWF�vj�3�`��%�HJ^t�عJҖ�cY�*3�"��R�	�+��C���&S1�	hv� �=�b`L�Mt���Ld%�-3�s
�D���q�H�(�NM�S)5f��u���.qU�Gkk��&�Bͩ�t��/h�H6[��L�;c�t.mDڼ�^Č,��ؕ:����뭩ˡmHM�b��`[�B���f��m,-"�E��eS� ��iB�#b-e%&#]��Z���p-%NH��SX]b2���+SHa6r6%m�TneȺ�T�q�%�z�z��K�`˳�B��{R2��HM	��ծ�f�Zb��
�źj�L�h[B���.e�Zװ����XA��f�ˌ���a��R�����Iv��@$m�9�+]�f,,�ԭۙC�j"����rA��M 8�-f�e��ia��*���Q��zu�e��(g��J<��6�mf1�h�ˡ&W=���	Q�UusQ��vmr¹6,��,Ma��cx�l��@�sl�jA��d�J���,F\hi�f-I�&���x�M�q	eݍ��]Va1�U�j/��4n!�45v���F�5�X�+`��J2�&��@�u*�Y,D�WF
���"�@%�-ibC1�q�Z)u�B2��$W�ܚ�&f��$%�Ё,p��@R],4��L,����Ԍv�f&nK�"��ق� �ʦ��-H�L�4Ԭ%[��be���W[�Zy6���v�{,�iM+�ׇB�+�\�KS*jĻ\�:hJM�����ʽ�a�3��*ݸv�.7T��c.��[Gu6\3)iP��RlijK��h�ű�9x͵��e��-��Y���eєb2�T*$pf
���Xfm�Sh�;6-�#�d�8^Y�l(mt%sQ��qlÆ�D�n&�MniSÌW ����2��kW\��j�r�/&�*�6lFs{��a��M�j]{��9v�[�D���ց,�%�q�WSs��j[�!6�.�S][kj�c����43����قV�(���q2����M5r
Qh�\$\ئl]r����-ҫ6���$g�p�m�����9�hZ2:8Kɵq�sk�+���:�u�x�&!�SK3fv!6e�(���f�m�L�G-F�f9.���vG�i]�PaNs!��XX��v���ke�YQ���2�H2�*[�k�:�q0�eV��,�,b����f�a��&������J��C.�[ٍm� �U6������56��46ih��+�t6�%fkt(D�9�r���3Sq`��
-�A�sVkP����4�e\��c[6������^hV��E��nP���������%�$&&.��Uf���aҦ�&b��٠�@�6�����p�}��p���zՍ-�4�L�]ؕ�A��aHY\B��'��X�޽��+W�.9�La�d�5���.�!�j��Z��k &kw��/]r�F���n���҃�c�;��ź$I'�6��NDB°����P��1&�6�i�v������믷^������o��=�d
�D��a�J5��O/!z!����Ԝ����t���o�ۮ��{{{{{{}����PT)Ru\��Y�E&���r
�Nqx�<zq�뮾�{{{{{{}������U4Ww �6��X`�Q�,�r!�5��)i)mb�E����b��4MHjjjmlimjjjjjjimKZ�LΊ@��Q""�J�(c�TM7-�(�Z�B�
QUQ�Sƈ��V��Dz�!ǒa5ȡ��/`U�j�d*
-Z�R�FQ�Y&�RVJ0D��*U@��¶�+Z*
����E
E�U�m�@:� ��6�"ʫb0+FIiF"���AE�F ��W�R��`�/ 2��m�*���DB'�V �&kE��b�b�`e���"��Y,EgaCn�X���kV�r�r�,B�=|���/hT9��i�S���bKh:HSIP*q�1̸EFT�s u�(��\Q"�(��{��,Sn���EϞ�w{����v��έBh,P�%����;޸�B�\�f���9暹�ũ�Ҹ2�{�*s�Yk�[��D�ʍv+j�^*�FM�jCsK6M3��Qh���[��ĭ��fRiQ#���55f��Ԡ�����X�L��M�s�k3
P�
�L���6�4݃EL�39��2W:�9u�:��TY�f�4���hgLd��!�,͹!�����l�.��6 :���%�f��P�p�%�e�.�i�)��S%�v�61lx¤1�����Ytm�Uf�0ֶ�6YpYtD�t�)t0@��d˶��1n��%i���[���k�ʧ**BЯj������%!m38��4�;�v[�4�S�L���h��ű��m��1�+TĮ���f-&�(�jK�34i�\S����mXBeƼ.�Z��h��[��D�<[�{#ƌl��6:�N,�t�.	��ؔ�E�#�m�l�"��T�F£5!)j+iƆ� !
�!����*�x�]J���[����I��BST!f�C.���Wi1�����m5)���P�p�5�ۍ�jmݑ���A��F1�с�.�t���M���Y��j�z�Slۅ�lh�]�������#f�WB�������M5�*0�e���k+kHC�\lB���H��c؍��r��Q�7�����]�1q�%˴�͵"�@baru�����eTXF8c�"]�L����]��R3k��y��M�v]� �M� {yo���1[e��2����]5J-ɮ�1Yn	��3�ƉJ:�nVV阱��ٍFaX��R��@&ny��sD�D9�z�lɠZ�͎%k�A�UZ�8S0�(Vj�Y���\5���鮅c�����8z��FWt�CE��lݟ	�h��T�ͷL旮�绸䓜���y�)�T�^*��E��VX�Q�#�F#e	H�(�H�-D�-�-�[`��EW��2�4�+x¤e��ұ`p	Q��^�m#
�e��,m�m,�i�̹�����Ź���e#jXE�ZB8c@�m���Z�i#*,�V�y�y<�l�_�����ep�X�d��j�9��+�g�m��M����83c��oz�]��!�{gh��5�μ�Dtt���J���}�Hh}��;E\V�.�FC\�/r�#6.p�Ud����k4��<��6+g����O)�gj�����=�Z��9S,zw4]o6<gլ��٪my���a	|/��`����ٙ���q�a�7y�ϫ0�Y�6El֣Q�/0�
l��g�~K�2c�ሄ��^�}�����_�߯���7���ο_/�q���F-����a�(m)�i���M9ֶl<X��m�!�v�;�ɿq�r~�y��>�3�w����ӗ�R�Q���pn�z�L��.�>��{.����_P��y��N�|��tn�5c�f�A���HW�o2��;z��僚c�]��7��sOJ6��ښ/)7��x���'yv��v����w���م�M�K�N��K�;�r��f�5�y�.�%	�&b��^����ػ�L����]���T�N;���i=���M�˖�=���L�F¼�[�/2�V��5�Qw��]߫hlTޱ����%��~c�լLq�=�����w֎N��c�W�]��HԆ�-ʿ��E�����|`��α�������Փh�G�FR��������i �̙��v_}v�'6F�{��{����CZ��T�y����:&��T������z�yU6�zHI��i����l	���M2�L�����y
�K9R�vW7��W!z���O���7HVkb#wj�XK�b�ڮ}|���.�����z�5�PJ f�ï;��Y��w����6[>l��5�>�����sgw�a�n�b&Nnȿ_�4�tMP�~���Ȇ��`�����
g���|��y�U�k5��g�������O�S�LuOM�AD� /O~O����d6����[/5N҃�5���`�-�;b�.����=�g�r�S3(Tm��dhz������:�K�/T@�Ci4�Ɔ��MP��;zl�i�N�b4:�L٧/.^�|��I�,E˳�� ���m?����!��8����1fe�<�5�I�`���}g{�'t�ϴS&�|[@L�3L}���/d:�\�ևc^���!�����ڭ�[��r��)�D4o���Л�}SU7�//�<�K��@��76l;%���]U��H��!�n�'6'u�^�>"0�x^�&T�*d��[_tV��\��^O�#�s�:(�������W�'�]���-.�9d�rO�}���ԋ&�5#�t�D���F\�W�F3J���F�����I�ex�e�؃(d�jˈ��]fMR���k�Jw)3D��Nd�rrb��/�/,� ���i�����^���e��A���fu�o6���R���g�oT�0y�$��m_��Y���ӳ�D7���e��͟�Q�1t�Sa��Vo�o�|'�C�Y�|�[]����s����a'���vS�=)3U�~�פ�B�/
VϞ�,�����F]�d"t�ʙ^nA�6R�������]����Ι.2�N]�<)Òm'�C��ЌЕ�0�q�O��7w%���!�x)(��l�;����vi�ɹw��WyP����vsz��}����ZD_6,�j�x�z����<o�sp�Y�Q���q1�	�[���2�r�3&em¶i�rtQ����/e`]����nc�bSh��6�\kSYk��/i�`2��.�e��0Jǩf�Kf��VA,î	��X�+,A��z�Z�P%]����ѹ�څ���;:�%�6�LۍCA��Q�i��t5���;�W�߷����l���ˇ5.�jڱ�3��	����]��8+x���.�_���B��n��d�}��߫Deyr~��3��SyT�įfRQ�����S�i�Ǯ�ߣ��%����=�	���Y�63�;E8g�&PUk�O��cg��B�Ļ~��gv���dk#�ҭ��1J�@��y�g=����@���P�T��qy[[~7���}FLxH�k����l������F�4�,��eX��}��7;�����&�)
�����Ԇ�1x:�Z���?�l~�4)���c-v�meaX]J̶\��9�ƥ�Ŭ�1�=@��KN�>i.�1�R�����F�7�o`Ǳg6i�����|{Mo���n�n� OIX]gX�.K��>�������u�������Е�a!V�c��2�!]��=_5�����L��ũh����������k��ob�N囨mU���޶[��0�|Zw��#_a���6���~�32/`���V��fg����6�ڷ�w,��t�{x1�
̖v0� ��(E{o7#w�{˛�1;����X�|DA��!x�hi�j1T=��Mn�r�b�$��=������n�϶a�fpTeD�ǯ+`�g��XA2���K\h3 :4����]�.p�Rֶ������5��l�^O���3~���¾�����4���2�j33&c(��K��g���܌�z�.o Ǵ�g�1������17q��2)l�m&�*g���:֕P�Dɘ�w�>�����I=N��n��C�n���=~��X���2��ʈ����G-|���-R_^��2�ݜu�_�;���-��;_s[�o�U3�-@j��NTDDD6f9i�a���B�7+3*o�Ίi����Ǟ��$�?eB[>�g<����}q��6)V����������ض�M����g͞�ﷺ�߱�Ko�������Ȥ�xZ�qhK
.�`n�0�&��fkZ��ӥ)������㓜81g$׹UY�����]��u��|���3O6j�>��ö^�\�u�u���ܜ̩���a�"$�H�bh�~i�w�<�ݿN�U]�a|<i��d�
r�g^wN?|��>�v-�Ӹ^-CK�	��H��2D������VlKk5��Sg�Y��Y��ѭ�7�4}~�o{�~Q���Ŧ�vz��"�Y��nS� ��V>�;k�M���ʯ�b����A,=��,�`�2��+a����3!�, ����g�������.�c&\n�χ�m�=c2��^�fW�{Cz��t�f�v}wKz��X�6x����;g0�!k�X �ñ�lq�A�&R�eF��إ�p�����e1i�/۹��؛z̼Oև���{j��臙���3mT�4��G��v�MjxM��eU^�}w�3w�`kO�Cl��9{{��/G��i���6g�g��S�����'��}�sy�v�+�R�����<Z�ik�ۗ�`)��hf!��~�ϻ��{{���=�}�$R�S�|j3��5�]ǘݦ�S(c�X5��@�T�+}��o�^��y�����F���z��jTP���Q�5��>S��}�;L\G|�2Q�aՋ���CY��t�ݳ3�"�+{Y��xo�]�..��3��	_�oi�k8����T�f!�����	b����,;���a�:=ų�Ny$����?={���m�)y����ntu5�@v�kr�l��TأW
Y�Myfq��1���� �1�1���i�����pV�t��mDl�˦�,M&�X�s�Eк�%�.�9h�6�a�l�aBZ�"�5�c:�rзbݬ&��V��hⲲ.��V:#T����X��f�,��V41������j΍[���ئQn*w+��J�'c���u3���jh�MM���k{i�k��_������U!����x����W�W|���\~��u�f��߭�Z��i��y�}g�Nr�����M����W֍Rf���:{����۷[���g����3���s:����9��^�GM}Q������6o��,��Av.����_�������N�r��zc�݆��ɞ�5�kr�H�qv��ʙ;�'ז$��<y]����������~p�k}%���}�}+���8�}��O������@\���Y����.e�3m]�!Me֎d��~��I�Ӟxs�|�m^��j����eL���d�g���y&�L&|�n�)�����r�z�Dj }//N�phVk�ut{3���R�g��� Tk�T����>�{���K��Kyھ˻&�z���j5Q�J�>�~��K����>o:Q���\n�'ͻ �@L��	�����ۜ���_ד�ؾ͛�ݶ��xh�Re���8v��uK�vqx���h�!������I�k��5b"E@t5��SU�(L��e1{.��6V uz���n��u۟O�{Z�s꯽���;���a/������e���hn��K�[t5JF���c.�24���*C*� D����\��&S��}7�{��ɹݽi}V2H����ި���4�2�wl�s��*��>j�]��R��S��ʨ�7��;L�&e�E����-PH5�&�
��!��*�s֞�>w��u�r��Ih���]�=�d�72Y7݃���%1b��۱�m�f,�����J�S�"nS��n���L�bB����.����z��A'3hb����c���Bq��<67p��U��4Vj�v�iEm�5%C6���<���۵�����5f�H�'��ϩ��q��9u�[�,���KN����{$��voz�>X띎�$U�3ni >g8#|�n�\���n���ʕ��޺�j_Lӓ郻wYsNM���8���]]нԶʹM��M�]�R���ڶ�Q]��Y��a�*U��Be��g���j�ko�7��1�:�/�OC��Ӭ��U��ĢՊ\�Unl�홂Q�i4&ժxd��sݠ��9�ܦ�ט�����8��j8�e
�.T��}�e��C��%�ߝ?m`��f���έ�V2�T�[��_^�yW��omo_��;l�A˩��4�dz<e��c43����˭��\���U+!���S��r�:���8^Y��˂U����վ}�b�4��z��ʡ0�r�5fV3��VgWn�f0��_ �y�m�[=D��a��7��ч��qE��D�Q�Y��M�;xl�+��׆�{h��ǖy�׻C�^Q�b��\^��cd��������N:���I��=��37P�+��CE:Z���4�L�ٺh=,88U�n
;�A��B�	׏(�bYI�"U�̣AfX�V��9�m\5fl��&	^���RI�ܯ5�bv����
`"�7�b
5M�C�ӎ�����������;;9��ikgP+��x�r�"�M%Ab�~�K2nr{>�:�|||||{{{{;��;�u)A�ڌ�5߆����5�hLM�<q��~=�~>>>>>>>=�ot^␨���a>��ɉ
�,%E9h��ON}>���������������w"�-z�h,g��8�H� 'B��� LI)��Q�aP�2V:�ވ_�ý-
��5��C��seY�[B�B�b���m�*E���.�E�+Ɖ�H�ʕ�`����C�$D���28�k)��C�7�8b�rZ£+e��m��k�qĨ���iR�m&G��H���l|t�,I�\�Y�eA�E���.�VL?�2}+(T��� �X  �dfP�}��˟^���`A�{LN~���{���l2y�\<�s6.�4��0�L�hI�6�8cT����';9�W�2��WLy�>�R{"�o��@�혇����~�� �۱���Qc�rR@���8�`�#��o_{*by�s��A�=N�أUƩ�]���x�=:*=�����A�AI9������jR� V�U��
�&��(��1��s�f�eb���s_����G����=����ww&d썳�����_["�"�C\������	���:�����C;܆t�{�5RJ��\�����u0�6�T2�S8��{��+������(7Id�2��� �n�����Z�0�A��M��= �8v��!�nS	��'n�2�[@ y��A�{���eLN��0 Q��v�C	b)L42-&�pyЯ/�4)�� �4��D����Ȝ�����y1���p@���`"io/y�'����$p8ȔZJټyʻ
uR��8,ǈZ�V$�������k8ڥV��
Y���"�%�'�g�s�l�K�u��?�eAle�X1

�)HP��O�������2a�n6p�,f?1�EY`6}wL�`�H8��}���k�7gg�:@��L�<XJ^-$	�v������z}�E�������w������ղ�Cd]��b�m��eKMU�'xPA �d#�h����SM&�����v�r�q��86;���9S��&�F�K�����=AI�������k����q��ϧ�����;��3d��S#��)��/=�V�U���,�p*�_%��q�ֆ���	�02���G����y�yXK߃�}�&��&�^w�q3��jP,5H8 U'"[֯|�3d�j:�����t�kT��y��]�;�=����윩��8��$T��D�� 7$$1��vk�[#kX��v�,� 9�\�ܧ����0r�?xO������{����̀NՎrxAN��L�*��:������p�C��'����6��<�����,��f�-ȱWg�\x{6��*�!{�Ӕ�Ւ&ڳ�M8���4��D�)���(�R��fPO�c�_{�����d�4f������RVFYBTVX�Yd� �a�H���[�^�~ѧ���F0�hF���!�����6��R�n�Y�ےh����h�%`a��7;��cI�Fk�Ȼ+��ʫ]��#��K�X;4R���"멛�f%5��b�.(b[i�lL�˛A0:X8�au�6m6&�$�X�:�`GK.�l�ĩnxb-����bb B�lT��˴�ݮu�K�����z��=��v��:{߄����ոûA���Xͪʭ��b����1��tV�nގL5i=v��ϲN�fG��m�X���Պ&k0���"�;�P����Ǆ���D��ȁ���k�����>yW�7���HC�X`�����|�8��c��{'&fy�s��E�u�Γ����� �f�&��Rq�w�[Z���1�)�ˬ[�#��=�w
޾�����5ɯ��
4\j��q$�8{�v�ئ�'9�KY��8���p]�r��=Bn�VC���M�\�@����2�+�8�8���\NJ^�Cȋ���S��T�Ѭ���� MS�j�h6=�9�51�q0�FK��ÑT��J���臇z��KL�,u�ƀ��9,����e&���XZ&�)���3،#f1�K�쟱��~�#e�!��3���~5Ԕ�vc�^6�7�P�[��oNO��X�3�#�Z����`�U;�h�r��^� ;'p^����G+3.�#y�����Ƕ���\�õO�z��N�@n����D������}�᯳Sa�I���
�2�����/<T�4"�*4	HC��9��wm|X;T�Bn�����7x:���&%9`Z��v<s������5�����Sm�����a:����T��"x{� �f�{����vg{��G��N�u5`�?a����1t��5HGf;�'"@`=��`G�����݉��r�1W������ǈ��a��-c �����V�`�����X�.��A�>T�'�s�J�#���3��^�!���M�{�?���0f�˂=�I����J��`w����v<{%h{�Z��e�Z ��]т��l�v3s&h�m�+5L� Z��Z;����������=�h�U8|ؠo�t�2�}��p�w4M,��X�44A9�9�9���2oe��`L�j��3Խ:�3As� q�L漀q/8W_���^<D�G8 M�`�p�Ѣm��{��9�0"��j_#�Xi��3�p��:�{z�7�o�!�^{�{�w	�V�Uz���A�����g�W_.�L�w�GR
��n)�ze�kRl���wyZ������������c��@g��W��J�HǊ�Ǐ�#J Ҳ$���A�y�����s�W�k����c��4��cT�pA5IȣN�\�p�I���fZ�8�@�NX�4�v6������wv�ٕU�s��4h��%9��4�)�0�vv&�0wev��R��&j�����7�@�a��S�9u���{�"u�p0���	��=���ˑ�ya�7/��/��x@�����I�
�tkV���K��ln��z��;1��b�k��?s�y��y��NN�UM�E�}t=����"'/אB����R���4�|d�)��o1�N3K(�!c�{��w�e�ߞ/�+y�\�k0	��y�25�8��Y����.���s�Xe 1���w����\��QQ��D�L�뗋b,X87h85I��Y�}}��>ݍzG���>��~���N�Y���k!�"�Z��c�v�&p���*ˌ�fxM�y;V;� U �sFoٻ��D�����c���;ѡF�3�Ziy�DSǽ���v�����Ο�L[�i���r�e,�`��cϾ5>߹/�q}��h�ߞy�/�O�?��3�P!,����Fx�x��<�(Q
T��!"$ R�Y�_�;?�r�N����؂�N����f��������or5��M�\�s�`H�NX��7�bj��m��/�"�ՂI6rrw��>��9��І��h�h&���W�@6&f�ML�5um���v�3^܌�i���`�����a�~���OLC���1��+<���'wa�>�_#����'z���T���˹��ہ�y0pE���U������D����'�NA]��ݠ�����S�'� ��Qy-8�����Ѥ��g{���~f�|.�s�G5㶯+޽c�4��@��v�!�S��4��G;���3T�,�-�!���A�OPOYiv�b����5���e��Z���3{qw���`��n#�$�~�����;X51@� �Ӹg}ۼ��NY�gw��#�܈��{p`�{}���Ϟ��Ɂ���5(���ꎅf�\�௷��]�?ڧ�I3�6b%���:͔�{�e�>�Q�'J�PB����=��n����?�~'o�6ڗr����P=z�} ���W� �*<�x�@9"�ǀ*r A�A>��?���ߞWk��#F\��"����h0�)(�B��bGVX��6���R�'�f�A�k׍lSR�5aX�GlsapM�$J�;k�6��������]&6�c\��lʉ�G.Kl�yRfGDn�R�Ylm`�f3��� �e(�\�P�)��Wd�� ����.�M�%�4��!��M�v�v��7�����Ҟ��rO�����2����lZ�[f1Ǳi���Һ����u�Ԧ��������!���"���p���ջ�~꼿{81�#+��~�C��'7z7�v#�̋��`��	�@;�N*�v��k�lP5�U���Z���O��_m�^�9�݃�k��o;1��~#C2n��͜�b�݃�"�p.�ul���Q+��]ưk����<*"kmyq̠�Ֆ�v ���i�9���xV��q��A�v@��"��8��Ӛ���y~�s��(���\x[���[`4�á�gb[N��1A`Mڡ&=~��@�5�>��*��v"˘O�r�v(���#=�*��[�y���^����Z����@��.Xv�7�� �l���E�q	BPh����[�X�3CPf�"�Ѣ�U�s|,?k�:v����!I��v��2��xNW����ǫt�7�@�P�ｌ��A�DKy��KV�`�z���>�7��^��5�\ٟ�']���x�N;<�Bq.jʑV��Z��_:N���g;זU�!B�ү���1h�fd���C]f���]���	��[�Ta̺�,/�Q�����Y��T8���Q�< B�"*�*PJ� H,�B�s)4����g��y�7P�������o��x�pX�x6�]�oU�̂�a!+#�쮔���̦v��g�X]�7�ۘ��r',��|1u���k�Z�Ø�&g���.'{�����y��}s���	�M�q�9 ;��ң�a���g���V��f�\��qk�]%z��,�5��ˑ�n<��e+��1�i���2=zi����L�w���r����6�q�E�I��*�؊TX/u=�\�a%��Nw��֮߭��b�&6J&�H���fCeѡ�7Y�����u~I�,���`�{f=��+mG�5u]����N�Ż'�X�
���d�sxb>���2��νC���?�.��[����F�g��!�L�n{7OI�z�g2�1�2�<�Z����ݝ�_�l3Q�O������AǙ]��@�E��<�p0#��u�,���7�hE����w��f.:�o0�wݷ{w���ʳ�wW�KU~����Qsz������lL|3 0b�5!XYI YH,��A�@��V���� $33 �龿�}������ƾg�_ψhG�y�D�̘N�L����<��e�v����V�x�j�2�N�p�Mҿfr�]pGx&Ő5h;|��c�@3�@�%�#u�9 ��W0^�CF��'we�����vI���x+��z��Ճ6ep��1
��d�sv�A�V=���X��x��ç�o������4�2�cl.̓�E�`�.��- �$]�k4�q���q{�(��S=��=�'�ݰ7n��V���N���1�}����Nׇ6R�	��}G9�	����_7)�q��1z�U��A6v�wVT�ƀ�.Fr��@x)�o��=uO�`�� A�P�O8ph�����!'��� !�m;�,d��N��wcJ�
�3jyœR�C�"�oV��͓½����4˓��w	�����$�n	goua����s�,`��h�ɂn�.X�p!��ks[��=�Y�Sp-Ƌ��3�u���A�첕�I��\�ht,������/�9��r�ҰxVN-k��q`��|99�P'(�d/�Q{(�9��v�$	�3�XIX�2�!���C���	 iYY@�hP�9�?W�������;f���,i��ǽ��V��s6��yN�v��?�x�n`����y�`�4]�U;����#/<��%���2�qu8.�br��	X�8qD��㣝GE�s4�f��vy���}����R~��b©ñv���#olT^{G�Va��G@���+��0zύ����� �[��oȱh��A�����>���%p���4�8٢��7��w��33�u�̫���E��G�g1\a�ϯ7�"[�{��D=���oX
���1�X�69�⸵ �B;��߇tU<]k-L8��C��Â©9Md0��;��w�v����O���"��@�B��y�8p���<�����X,���Z� ��� )���&ngd�r��0pAnX��U)��w�x��`�L(Ome�7O�z�9���N|�=�C"k��w��I @~�{����r��V�'��ŕ�xS��r�nk ,�L��NB��IE����£�mN�_�]���5���r��V�o�Y����)��6e*g�kݲo0�6!���>�W^��s]���C+,s:�i�x��$� �cw�l��W��:`�x��/����Vo�RI�V�SVU̽ſZ��.	�69� w���d���VN��ᕷ���]u�����(g�w�t���
�j�<Û��=��X����7�ι�#:2���1w_
�Nb]��L��M�^=[�u�i�X�Q��2��T	�Р�o���Ώ4���}��|E�ɤ�,��� kk��k)��9�,2�&_&ܓ�&r��C�L����x_:51�����n�\\5�+gV��;�����+��ƭ���]��}�8>9�ΠwI��np'�4z��Y�]��V�}8ݼ�1^nN��'g��yÞ���;�e�K93�j�-ٔ^O�;LC�Նf]5�V�=�p�5:�v���m���`��C�eʝx	�!�֝��垾�- r��6x,,w\q�ͧ�Dn�,�͙��]���r�Ы�\Q��%�tq �U��[�C-�k(��bt�k��B�۩�/Z�{�Y��]Yu׷B�m �b��]�U0��'�5R�v��X����N��zYw�sG�e+���J0gveY��ӫ�g�����82�<����h jy�0A�	f��>˔��Y��]Ҁ�(j�T�X��������O1��*�Yoq:���N�&$�ʴ1��;���%��[	����W6İ ,mh��y���7Mgr�,��N��[��톂�������[�� B�׺K,�A+mH�V�l��o^>�2�=kc!b�ۛ+�wF��O4�yW;kPX�Y��ۙPEE�q��\s)X(!�L���kckkSk[[[[[[y8x>�+Q���TM1
�c�,�T�(即�74L�����g�����y<�O'���,=/���-`�mn.QTl�(
���Tz��}�:�o�N>�u�^ߏ�������y7�=E)�+�m�kjX-�eaU���wf�>��j{9=��'�����y<�O'��U8�&'��u����Me'�]��6�UJ�T�Y�C&�o)�����j�ˌJE�3*��sr�6#b�Db��*�K��TC�Tʥ2�°]Z*�-��D�Z0����c����V`�R���c-��
���,�����X�fv�8שb,�QTmkIUWv�"��V
M�咶�)ցBJ���3OC�K~��#��ó�N9�3f��ٜ�W�����	c��c�d�I��Ż2�R�t.���V6m.��&�ٳ��!z�+0Ѣ7Gm(vh┫�^l3ڽi66���b����2;`���.`�I��k�B��*KIgKZ���X�k2`�ڦ��6�iЀ�`�:�v	��-���qV�C4+H6\Ķ�m1
��fd�5��%3TK���<{�x̹m��0T,��+Q�H݉;к`iY�tm�r�J�\�"���k�b�Z�Ů
�JB�Dζ-5.ˣ�4k���3,�)[�F��!�ݡ1Eeֺ����%X�"1:,�*3Z����\�fcb�l��3V1�l�0���6��%�	�ض�	�e�r��Ѯ"A)����CK�]Un(XM0F0`4n˴�@�K��s�)!MmB�i����v��gJ�A����a��,�FrQ�����2ۣ`�\�V4���)Z,E�B9�b�v��	p@� L-R���@2W�ʋ�Um��6�e�e�	f�$�"F8�V�Z3hU�6Ú,֨��-�4�l��(I���s�]7XШ��susl*�f��ԁ�0�t����ɉ�Ih]a��s�7�Y�kfȯ (L��fL`e#e�%��jl�GD� �56Κa������n�gq,��eHr3��Tb4�����q��D	���c+���e�(��pf����u9�	mqZ��Sp�k.-,vx��hl�ۉe��PہA�p35��v4T��jܱ�s���=Cǻw6�)���h#����l�h`F!Z���J�+	Z�L��i����5f�ˋ1`��̥c,[շW]�V�ҝc�a���.j�*�غ�Zl<����X���30NK�v3��1v
�	|�t�	�x��w��͈M;a�u��-�ҽ��t�i�+�!%�ҀB�e��*�ǊǍ�hF�@�UH�?s��|�v�0��SkZ�UW-��f��6�gL�flrd�4Xۜb�q��M+�!Q�a�M�Qؙ�b�3	V����X���\їku� Ԯ��u54�D���q΢ҵ2CpC:Yz�,�-�e�1��j\�l4�b̵uС�3wR�S�e�^m�<�k��e&%�l�dk��fэ&��!���y�|�)������6��[6��Pv�/�f��i`�r�4#���y�y����@�V�C����r��v�)�W����Tepe��4�u��ӣd<z�{�Aa��j�$�f��t�����%]��A��1�0~���yÅ�Na��5F���{C~�5��c9/����7�<�0�ن^�2'{p{��:���l�o�N=fSt�vr�=����u �ѕ%�
����RpE)�稿^����4�x�z���:���qx5��FW[�8 ���D�uG�wH1�(�� j`��8,38 ��NAN�U��>wR�-��G��I�Wh�o�vep,1�����Q`*W�&�3>��.+*��O�NH(�J޿��38��F�u���H��nP�P����3�R=dpF�s�8u�\n�pu��׈�A�;o3[���˜�2�74����4�2�M�wH�dSKǘ�7i��+wc=WEZ��4�s������ّW�5��7n���Cn��>����r�=K����"k���S�6���f�v�ͬ����o�����@��,$,�T '�C�� �JPiP��������"�2�N:"��ё�m��Q��#����'�9Jp�$1���X�C��]�$n'v�ȪV�@7hyMgq''�&��P�nX��ze0�N�j���yU�1ܞ^V�زR�y��1x��n%�e��3[���˜�2�8Ԝ����c7{x9��-�ڒ9��Q���'u9�FwWGor��̧^�=���W����p��S��g%�\G�ü�ݷ5��"�����K�%�9�ԇD)��PT�(�-�I��1��L�p�|��#��O��D�l�L(��"6sQ�V`�V�es+U���Vr��9#����»ø�A@w^"��d� X�����Ƕ#bF(mh��/\FnN淺'k.s����@�p+�k/���:C�1)aRvL�;��h��^���I�p���Q�)nf.�w*=� ճf���n�Ԏ�R�}�pV��&¾'�
�y�Ͳ5P��3~����{�������H(����Yd�
A�RA�R� �
�%B�# }n��GT�epG~���b��8)�Y�"��H%Rބ�^b;�Go�����p����J�~ɥO{ĿVM������NXK
�u�K����c<��(ӯxQ�{�2<x���9�{7P���nk{�g��#�Zs���#%	W�=*!<}�W�����U�B/��c��1,�m�]�k�p۷f�,��%tƊ~L.b=(3����j����/�W���+B;�l�����C1N��E�-T�CJ[�f�U�0{�����"�<1��ks&s�'�&�zW[ԓ�)����LC��}�����_�y��N=�����t%�1���B���܁ղd��鞡��̹��W���"j}�4&�Zv:����S�]y��d%ň�k��n�ݗ�8����Ԝ�j��UGWd�Ǻ�{+�;́c������	��X�tnW~�4�i����ra���#��N��0'7�h��������`��2��φ��I6�.�?�P�~���
�x�D�ǀ�PJ
�JU�Ώ���[�d[󏘌�%��,��ÑT�rNK�Z�a����!��o�;��g'*�zW	�' Ң��A�W��Qk8uf+��<"������4ֶ��
ef,�M1y�]v���Ye���6��9-�a��Y��N_��n^�f�|��r{sd���˜�ejX���9\UF�L��`�.�������!�e4��\�lr�Μ]ힾ�&@D� ��ꪸ��݉�59\�8������S��w���w���q��!���U ���b)Q�1����%��!��o=js����|��:����1�nD^���4�V:(�83uX���'�"�n��g1����G2�rǎ�>hAE�D*{�-��L������$��k�g�؂-Y�0�����|�@�e���a�؝��s����9H�}cG ��2���g�;S���F]-�����3+)�}+/k��3���K5�圹vt��u�Ɋa��^pܰL�w��}�>|!����t��hK�1��yf�!;��\�[ۜ�'���� ��R �,
���%d"�I.�����^��y��!m�5h�*0[ÕD��Ff�ʥ�pf���˂�R�qK4�l,��	]�(�i+WK�	oi�ܵ���YfBh�8*a���L˦5[���mk���̌IL�\���3U���m�i�mz�x��e&��4��@8<5��V���k�0Eu��4֫,���.���.u�n[�f{��6m<�N�������Oϙ�鬢]�Kn����gi���5U%͵��U�B������F��B�Ŵ�r�8k6C���}���d{.�_�+����[ҵqO
����pnӐMR|d���Av��d��g2�����M�c2s{_�����T���;m8,��,��#�u�@D� �'���dʩ4R� ����^��Ui�ȝݛ����Z�� �8v"� �T��N;��6�9����E�k��vv,j�|��}����T�zW1oy1�=�5��q��=9�' �n�2qC�b���p�]��^�z�Ӡe�|�;3�#y��ݔ���6��2m8q�C����8>�;:s����BR����yhpsfé�Gs2���Rc(9��m3����s��?K/.��y~�#/������h����z���!�OO�:�I�p�]��9���	��M�F��+�8ǋ��wx�B
׌+S���3ќa���Wo1�y�W,�Uh.u�o�_h7�x�ر+l�="�Xt@�0���R�+(��fU�Y}����Xv��(�ZK�`��&YB�A�P
�e��Y	D�`	� z ht�v'���o�}طљ~�}��5I1v5K�z謬�V
l`�b{dƝ�9�;T��*���*��]>V�an��f��E����R��RPLFJ�A�m@�"�;��K�Ezf��L{{�KwZ�k�OD5�vW6v�jw�m��#��i6����^�>���h9N��F��2	��8"�ޗܿz�:�8Җ����{�ڻљ~�~�� �L��
���F�P��瀔�~�����Ů�͆66R��X])��p1aci`��2�H& �d"d�{�#YA��C[�f̂��q�����=���5��5�����>0D(	G��"ۙf*,�
d,Y�����4�7o���V��b�l  )�[��;��z���'��Nn��Y������y0)��]y��2\��n�4��^/I�A1��t5-�E��1oq�q7n�p��p���rl��&6�� �B���at�Ҍt7d3�޾�l{��M�P�����9HOx��� � �J)B'�:޽ٻ�N}37}�u����w��'oS#�܈����(�p�������o�m����p� ������ϣ'�f����_��%ה�gC������;KjDH1I��RsB�.
ʡ!O�+�!л=]�痳w�w�^�LU�pG�嶹���ٲ�
�6���bԄDxQ�x�Xa:%��k�	J�6�b2�
����I���� �����?o�~�2`�)�\9�v"��d���;�y��J�)1��=v��Գ����R�"����cv��u7���M1a��<�`Fk��e��9��a��2��Ϙ
o70d$l�i�c#�j5�N���a��C��2�P�bv��$�x��?x�]���!�>���űwLQW���\�u� �+�4^Y0���T�=�\.V� �6o �b,��*�X�����w�zipT��>���ꘁˣB(�c)� ���[f���T�g�ף�w=$�Q��6R�����8(������u�U��~�&i�-?�g��
��)!e������"��20bù�;pE��Ju^A�Y>����ٿ2U�����ң��1|�*2��wK��v�o.v6\z�*�xR�6��հ�z6�ĩ��w���A|���cCf��5t*$ڶZj)������؄\]VVk��.�	|n�. ����1qRg�8����oOW��̮4�Ɩk֛m='X���}����d~��#;����� U cNv*27`D�r"�ضk���W�Gv�Vza�қ���G�� �-��3^��a�X2鹽o �dʭ ��n��#�����r3g�r���8�9��8'1 �u8r*�Ĕ�f{(Dn��^93�m�˞��hӗ�9��]����x��w��Verbqp1�C��D����W�r�Ǳb*�w�Iqw�k��N��^��Gmq��{�<Ϋ�F�������́>���-Y�v-4�cEvlv���Va.�/P�)��ۋwͭ�.���n�s9ڭy�v��G>?�Am�}�{4�؀¾x���n6N��׻�YP�%h_T2P���<x<����<S��Y!D"�(H�!���3]��5@�uoH75е������\�J�5��HW�]�T��X�Ic[�9<O&w4 �tVؑ��۴�2ݍ\��`�!�c��8,vk���&��u:���V�h<�e��W�m�d�Tv[��1Mk��0F��E�4�.�B%+�I�V��mo�v�	b���º4%�X��2X�������Ҧ�ThA��J�6՘�v,��d�dn��ת[�O�&?	� ��t���E�5N>^�f?;�N;�7�0p�P;8�s;�8�gPZ���8��!�+e��A�NE�x���Y�Ai8"�֝����7z;���2�C:�8�r:�cf͙��zy�� $�pXd7K:(��h[HB��؉k{"�ʿn�/���^�zu��s?o��Dw���޳����nYFuT!��E�3gP#]1pl�rN�����}>�����o.g��.�9�n���7�Ր�,�'bʨ;�eK�>-�8g��zj����w�c��fV�s�0')�[���f�![�������B}ݴ����M���A�N�V�\������e�;V'4`�a�m���X��������s��WE�!��yU���|ɴ��\11*�ևT�ʅTZmx�Rx�IqF�,j1�������G�B���R���������KYX.6���-��+��2鱥��D��fa�?��V��ٿ�s��vk�����t*gw;�}��l�n���>�(	<x�&x�C�(r�i�t��g�s��n/���r4y��=1F�~��]�uF�(s�ն^!��Zh=�ȳda�R���}�i|�}��[q��z�+�9�cu��@ ���,�p��Θ��Eq��j�~� �������~���_'��=��~�&��  =�dfFy܇=�c�."����i��N�K�<�no��[�x�tZ��{���|����Cr�qMm���3��&��r�}��� ���o����R�@�����q�l��L%��`�,�� w������-���{���}������ep�|�⸿���.���s������w�'{q�ӻES�͙�6 �wL[ic7Mu�o#��(���p ���j�U"����X�g��ݮ<��A�4�9Z� �v�Y�ff������}OUUS�+T*O�k�����#z�"Sy��5���Xт�-h�p��݈��qu�Z�Onr7�.z-����D0������Ⳬlq��6=�ۧ���.��dv�s
�t.���gT:���M�z�M	[E���w�<�b��\u:��׻>���:�}��S>�OL��6����bu�����]ը�kYy�BA5�D�9��z�^�V*��/�ڗ�m��&p����{%vQ���=��`-O31�G���7�G�u��A�Ƒi��v&M�2����Ov��Mֳ�m����u��}���c�<z�mk����N�[*صܧ ̭�݅�/&j�u���,'=�Rׂ�y����V��2���F�\�^�0e���k��ȕ�N�gp`�oj�*�6B�7��n-���m��[b�ޙ��&�f��Zܡ�N�����kk)��:���S S�nuwcغ�[�@�2 z U
%d��(�e���a`�;9��h����֞��6z��F��X�>y���w*'��k:�=����)JW���������wQ���kfWR��&Vn��?�3nv+M��xa�c�4s�_Ҷ���|��ϗA`��3or����r!o^�������=栛�/u����M[�Mg�ɭЉ�;�U��z��嫛�v�Ƭw�i� �>�����vx*�S�:8w�h�g��Ň�wMx4����|���սq^j㧚����LІ��>J����	�ג� A͍��cfb�xz������`���I_�K�B�Yg�C�T�J���IYɄ�&�g�_�����{�O�r��B��Yr�����������������>�O�]|u����������[Ƹ������uB��0EV<��Qb*6��9Lcǌ����]u����������*��V}K�l����V�c��g�]\Ǐ��]u�_ߏ����y<���iz�"�y��%��� ����	�o_Ya�%�ޣl��\ZV��cUsp�Q\�X�-�Q[w��D]Z�*X�,ݢ�%ee݅T�YZۼ�-Ucm�Z�����o)r:Ɏ%��QEVң<�D��&��(�ƈ���qUkU`�)�bE+(�SXX�5��R�m���Qa�1�e)���KD%����)�5��P�B��(�*(�7�j�c`�Bd�)P�,�,��YI+!#�Mͼ�o�כ�����sJ��"�9�)��;v��ݠ�j���V�C�UI��O�e�cHq���������X��!u.3�k6���=I�5��c8��v���52���5}�c�&c�q��#dd�P��Z8=�}��D!�}H&6l�i
�8-V��r��΅���w��r��Î�]e%�қC.�Pз�Єh��Z�ʘ�M��=c�)�O���8	��B. U8w�˾S���Z�iHRȜ�*��idK���F�rRpA5I�ʊ�������Zix��|�[u"���^=s�Z�d-I�]��v�F�N�9�#and'��� �l��wb֬��OMΔ_D@S�5J�����~S���i�`��^��u����uzٖ���A͛.Aj�ɟ+��:��'2�sJ��gK��>Sޗz5*�9i��?)��9�9�i�����0\Mh�n��m_L�3F����}chU�c6�KM����h^U���{�ş����e���)�,�VY!2o�7��d��0��L�ۦ{�	db��R�f�٬b�P�VL���x���7�c�pAV��AN4\�*�Mp�<f�A��P�l���W���X|�E	�H˘Ki����W/�,��B���gR����;q�r�T���dXٯO�[���~�.�Na�WN����3���Q�n�:�
 ��Ò���|��*��FL1@U�w�m�;�;ܖ\g	bRa0����l�/�H�?���}��^�A�T+-v�A5Kj���ߪ�M?S��79��3yZ�M����ÃF�8���p�W�ĭ��΄�1xm6q��ج�G[��; �i���}�s(��q���\A%x��s<��Ʒ�Dz��jg;I�4�A�C�@����B��������]���y�����	�A� �^Ʃڰ�ʾ���]���MU�q]a"J�ʸ�s�#m���)�Q;���^�._�^<Y�v�����=����\	5���.�]�F�a�n���ͺT�U��ܨ�&$X ��3u���l�ޫ��L.�!;?�
�e��)%�R` ���g�����'����rB;S�l�4R:[D���FZ�g�e�*^ۂ�j.�%�,5͹�@��&�Yj1lÁ��Iv0�X��t˫�H5����H��*E�)� �l�����[�m�Z���%at��Ι�D����aYn����4�'L:�.fz�aYqHi���wXn���x�lڲm�ߔ���Sk����h�ۤcC� ̺����44f�`���ϼ��A�N�ɂ�q�a��pA5i�~�[��y�s7��p"�r�y<��fv�*У����p��Rb�pDg��1�B����_��G2�q1yegz�sJzdRa--M%�$D��3�rA�H� ��o�?�����d�Ôn�1]���_��N%��sp��i`��tݡ������w���Юw�S<����4���d9-8 ��Nފ���o�]�epG^&�&E�O�}�&/:Y۹��K8��pA�e�-v��۴%�P��ow~��'���9;95��xz�����})؂��� �j��0F�n?�� �,�=��p�B0�ikSl�s��Ch[K�,k�2���0�����	�@?s�4h�H{�_s�|�ᙓ��-�7�"���P=H�gm�E�TC�K�PŮ�[3 ���{��Ϸ\8c� W��/��ѩ���XU5zs$��H»kpvwm��W2����N��o��y��M2T6³}�"�CI)����*���kz��5��?�$�e��-��Ò�CH��g_#o�s��'oEO��g�*黚���r���h2���yt>n��S����ΑL|;S^xc�ū#	��~Ѳ6�:�������+;Ըb��3�#mc���p�z�8�!�����w8@xIB�R
� 
���gg�����j�궨2� ̻/ �`#G{�Sx���CLb���$0TN�c������Fgi�y��%��16X��3������
��J�sT�Dx9�T$�\mlo�z��k'�7ɳPrS�cF�=S����7��a�����Ӯ ̣kK��FXm�U4[�Z�;G��sBҘ�#�h��������Uxb)Q�U�3��\���&zt���׉�U�ud@G��a)׸^���w�����o�c�N�id��`�u��;��ˮo?>1@����T�O���F�s��˾_#���vgsh��n�j{}���BK�/I�Dg���9��&������V�G��_��V��U�;�`�㙣��7��;n������WZ�����k��s�3�ɽ����@�?��e��RdɀDiW�W���W5�̯�;%m���l`n���v�ō��
��؝8��Na�]1r7\;j�q�Uy3à����昣4��[�F�H�+�A�>�rSH
��R��γy�-;�v�\޾G��ˮo:zM�[s!L��a����	��yE{:"y�;^���8�l�A�沸�l�]�B�����j�;	6�+�_�'yS � ��9���6��;�UuY<�����lR}�Z���A�/��j�>B�S$-ӂ+ў<OO1� ��}b����Nd��)�>��. �Jv �����q29�idْ�sr���� ��߄z{��7Q'����e{��]sy�;Y���NRo
TC�*� ���)ܫ�QI,b2��ߓ8�sj$Ec��7�z�겤p���:�A���:#T�;Q��=P��G���1Io��<�cQ�f��Ub93Xg+K�QI�o6�Q+nf��Wb`x{��¤c��%��7��o�0L�JRYe �$a�߮#��1S�vpL��+���lMw���zb9�1��55�ï�ه�ޤ��S�b�:i
�B��݊�j�ϲ��D��}�1��?������E�SX�k���K6!K+5����M��,�xs�v� /Pr&�y��)�2�gGj��5�|�~q8{m�ߟ���A���X��� �8!�����m��}�#�δ!�JpA�?���vtwEM��s+Mx����U)�U8$<��	8�.�#<��k��8v�D'��=o���ٱ]�����T3� �OK[�y�p�b�[1>�֍�5��=_J�#]T+�5a�,/*�?F�����'.o���:l��x���96%�^p�Yc�63ݯ�)�-Yj�7�ޜ�؆+S�Fe��������pF��ܷ�v:Sz�X�6l��m�s��w>�7�T��fr'��.�� ��+���3�3�/4g��m���_�Ev��<՘�#٣��Һ���!�ˁ1ꘑ��g^�%B��[�L�2	�Y2`����~����,ʆծx�t��i,\��E�%! B.��m��Bga��	�\JJ����B�s15ay&��R,#Zܫ�Iu\�#ad��ҹ�8r����2 �m�,����W	F�M`lf\�rۜX-+�&2�.��6���c�����ٛg,�b��D��ZM�Yw��̉&�k�O3
�շ�Eد�Er�k�ilq[Rm��X��V��)Yi��h�v˂�;�)�_�g��.A�p�U;��D8�ʧ���]㓋�ޥlG�r������1I�i���#���6y|�E�w������:th><\��r26��F��9~�o?��Aiűq���g2i���AƱ8 ����*!�Q��$26&�5a�>O%�ϫ��9���F�1�V��A�v�GĚ���$zfur��zp�����vv�D@��*���Q�f�~�R� �>NEoN��®˟�D�/r{dR}d)�g�`Nb�-�k7,�{{������#B.?��+�z}�Yq������c����̉��no��K�I �AJg�0�'�AwrF���	fjF��l���e��v�Flf(mn������NY��9���v&��i�`U �{5�v��zk#+�7́�ApL�%����u�(�n:|ER)��+�ٺe ���F��m��b��Wa7Dx@v4v��x��=ݠ[Ǚ�WX�6�Iw��]f��J]�2��)����q��)�(P�U[��2bŒd�2�>")݈��;Gu*���Q��_�Ը��8 Ң��{aWO<��c���
	@��{�b2Б�Vl����M��$�WW��̵z<Ŀ ����8"������cia
�7��&Սd!���,a��k������[鬌��	�A�~��[��^g�缈�>0g<��vaد\�����֦E�Y4�a��rU��y�M�\���½�*�~٥��g�ȣE���>c��]��@3k��+�d��� ��O��2͝Xp&\�5�	�	�yݥ*�2S��ݰ��F��c@M�A��Ú4\�N���P5[º��R�i~<��%�z~�S�K,ɦ���2N�ܚ���Dk���޲��<��Yî-��ljӃP;i��^�GTF�Mc��F��oPru8s�T�y�/����8r7�gK���8r*�;CR�;�%�]�^]�c<}��Sn�,��{Y�OJ0l�ϴ�՗L�4�`�pgO��np�Z�$��w���{f(��%h�y.ď��d�2L�&L�T�==y&{)]϶i�d*-T�,�R�"����GL�;�Pv �;i�� ��{۶!_W���W��P�!�p�pBy#���)������ڙ�( ��pA�d9�K�K٥���X�[�������X�<�b4'��������$�G2EK����Bɫ�H-1����,���Fbh�<�2Ar��2�p�8f��.�W5}>Ƿ\d��l���Ȼw����5��q�g����f���zN��5�M^VC�NS�;��<v�P�,rPr1�x�9W:S=�����e��r_z�*��u�J���ñ�fH�;�MD{�ϔ�~�,U��xz�t7~5��!��f}�ۮ�K��T]Ltd�>Oo�k��:�x`�b�K���@P���t��.v$��k�Ga8؞	f;��d8��i�3#d�e�����@{�7�m�:��wЇr�=�ʕ�p9���lܼ�[�qnS�GgQxLrd�лۄB[%7P�-'י'9��߃,�&(��*����o�G����;�=}�,sp�cjwzո^���:�j�VÅ;�U�}�We+֗���6Y�y�!T�؈TEV]E�Q�@��w�g%rSRg�y��٬ò[�Kbm`�J��Y�v|�쟸I'%:d�hHp<ʩcy�1�5���ݍU;5����^:2����6�U���p�٢��T�Ux8&�h�b�;�+vrd�9Z,���h�o��fdl�vZ��tיی˳9 �^!�R�yG���ږ� 8Gw &�ÃF�8N5Uno<l֟E8$�{�V�o��[���]6-��T�4D�#���Ɋ�+z=ج6զs�|�y9`@1Il��G*�����Ў�<�ό|V��C7.y�[�8x�r�e�6�c�$I����Ȫ��vU5�TEI��W~���UU�\�y�\Fy|qG�.�h0rI��wߖ��*s�u���w-�;ϬU�A)��k�
���}��*�u�(�ꓲ�O��SHe\�(�w't��� ��X�fh�כ��Տx۹�G��!�nR�����4��{�mBMc�;��2�^K�s�(�Õ���B�5'"ƽ��ھ������AXV�9*>���b�Gi��Cδ�]�WVY�Ѵ����ۏ5��$���ݽo��8eXgL�l�4f�����#��+N����ՠ�7o`;���c�5V�"�mW�j ��c���Y��ha{7;Y��w��N�Z�gg�t�����iU�b5C.�ɺ��O������"9K�{K�U�F��ݢtT=/o�DT����j�jU�ф��}��;��٣z�۾��9�d�qE��Y��N�r�C��l]�92��n��w�>�����+��99D���t��D	�6&�����W#�8�nef�E"��m���z����ծ�U��=eӺ����d��fգ��i=&�}�2�� ���t�i�R�����Y��㈝9��3�z�����םCyZ���j�Z�����t�\n��^)]v:�V���eBҽ��7�ͮ%��ヶ�����tyF�ug�u��Tʞs/'^��Z��@��Y�ʺ�Ph��szb<���;�zVu��b蝕�w����̃WJ��{���R��e�0֛��%��5�u%����K}�|�7^�w�nf)�"C���-3�z�Aj�X�&++R盝nW�6�J�;�2��E}[��+T��+f�� �a�c
f\��hLO��,����|��߉Ԇm
ی,U���4��2��t�g�mHK_6��iy�����ɽ;ٯHc�帽/|�c��T��u�l^�fk맽�f�;X���|��	�-'���-Ի��v_ ���n�\����E�mU�����dJ>a]�4ҲZ��g�ǷǷ�_ߣ�������l�_32�����ٍ��V,>�eVn��-����̚���g��������������G>G���?���H�+L��A�$��8I�Acǌ�㮺믏s����y<�N��zʅ�h�un_SY7lL����ԥ�E
�*����DM!�fFc��뮾=��5���=�2£B����h4U
�P
��z��S��
"#�'���,6��Z$D�TUXu�("�h�H�
���X*�dGkQ$Z�ݒ�\�i���,$��.p�
!���D��l
��X��KX�E�,�V��U1��X�:��5թ�U�mDX(1�T�"�[,����R�1�Ae3�Jw3B|�kLu\_�9�u�se��f��+�h��:l0+��K���z�d����e[Q�,f��m]��uLۂ8j�bK.�j�p�u�K�)�408�ZB8�4	�6�ht�{a+4�?��{����E�nh[l+f�`�-&���h[4H5�u쬳l���ŭq�a��p�F�U�J�Օ�f3E��kU��FW�5VRRԆ�m����t�b 2�*j::�kn�*^[)�ј����	r��j������!��Δ�qk��j�L\�^)QY]v�e�4<�&���M	����K�	���A�����*`�mKW][�z�u�R��ؚ4�yR3���cJR5�Q�@q��,��k&e���e���p:�آЕj�Ԗ��Y5��5Į��6��8������4���mcl �F֙�`f�ãˑ�������.BĨb�&���6[��Q�sm��Z���S�,z�0Yl�E��P9Yv���e�R�@Jۢ���&�;uX�15�Ti-�CX8cx�ե�t&[m-y���$�0��յ��kU4�셎n�Ջ�cgj�74n�� �\���D0�a�LB-cM�m�5cH�WYQ.��n��Ku%)�r��Z���Z�F���ҥ
��˅ֻ3Aq�%&65�ca����J�{�#ZF��b6T�k�c�b�;v֐c2�#m6�A���i��˰��p�Xgm����.!��;M�պ �t��bblĨ�HjŴ�p�Ke�c���b�A"�kVQk.D���$!�Cs/,�)/g�����`�Լ��1��Зb؆��fԶc�[*�f��Aˮ���ֻeh�瘰��F9�i�CuQ�Wom�ٚ�\��m�$p�b�܉Smu�L��tx���I��/^,:��:��s���:�u�i\���h�V�Q����*R:�Rg:�K<��`��50��P���Ɨa�.�bB 9�39cr��x�-qak��̊��pU�-����Є��Lѕ,�Q!/Vh�)���#�[Ic��#LZ���)�Lԋ&l!H���$2�����+.�)rԎ5���9aQ.@Md%c�[�h�G�� ������(~`kn%k����������,)c6����X�����o�n���?v�"{�>6\�9� '�՜�޿Mt�i~q�g��'�[�~��^_K��hP�G�B�j�X�j3S��F����#r�,SԪj�v&��X�z�d7Ƀ�a�W�$`�M�[D����;�WB�.A�p��ƕ�}B�@��_M���ffZ��t��A�T��!�R�4<"7.��F��ew|�cQ�]�=��Z�}��:\b��?D�����zk��K�t�2�;ce�W	5|�ȼM|��bqYk�x��p� ד�%�������
_�ʾ�}y�������@���-����EȪ@��Wt�����A�|׷�D����ю��]c^,��`�Jl��р�Y�h�#�R��w!���<qT�����"�d8٥���p��S7�\C�g���wǅ$k~<���NAn�Q�	�@����=���$r�S�3�"�)ONd�n�l����v��4�!�SݦE�2!B��"����|{�wy\P#3߽�e,��YIX�����~���y���MWa�i~~hd8������q�)��g���zV�($�_����Ld�1֠�.ԐA�I��`eܴlU���o����#�vJ� �i��&�+�9N�
��4GE�F�"iÑV��Z�J�>��u�s8Gf)��M 8�'�L����z<� n�9�Oq� �h�H'1 ���!c&��r�l�+wܔ��Wd�iHp;h�p�X�L�NŤW���\/8���Y=\H|��`k�,�Ԭ+Jl�.&It#��LZ��?>}~�Y�֔�����pF��w��g>��_Mc����[]�����ѽ�X�H	n�m���ƍIut*K���,V�K3��uX"}-��@��~�y�;-zs�4���9
U�BR�s��dV��: �?uPp���n.�a�����p~�ݿW����Ev�ϔ���J�I��I^>D����t��{�]�2o��n`��u��ȣΤ{�����ý�o������I�,�>�mo�/{f��ǚW�	�d/���N�iQ�eT��8�Z6�t�Uqm�ǀA�S��U��ŧg���Y�}����ι�&�{SN!����Æ�х"���&͗,ۇB��}�����8���H��׋�e�|��8ءA#b��+CS�EP0�=y���)������t�n��8��uxF��^Kj�ê��ɛ�W���_�sޑ�Y��Ú4\u��LNet�O�eWd-i\�u��k��3�{:��(#-3ڲ5�b���������|����z�(�!��N��{�����+�+#3]��#�jvY Aenѣp���]�X����B�:t�b.�pES��iQ7HӲS�箹R�+ַf)�{f�1�&L�"ۙf* ���̆�BZGq�sÉuG��^�n<d�T��s�z:�׶�4��	�Յ�|n�'�t ���d�$��V��W�:��6�0c�[כ�������ީ5��\�j���u��O�4��|�?O�1�cd\փ\���nev��n��ڲ� 7>��a��@=	�ѳw��WdVF_t�b�X㘃�7> �ZE؃~qӵ0c�F��E(P\g�?��~�ٛxm6�b�&��1u��76L�MK�6����
#��^���1�w���Ң:n�����r=��Zh㦔������@֬i	��1p�bl�{k�����a�� d�q���7�/�*��셴�k��p�_i��5$1��'�� �W$z��yx�os��g���:�8�w"���T��n�G�ː�w�OlVdM�_
����L��׮�)g{��pGsC������?y�3��1]�� �8v"u\A�[����]g#���. �����j#m�:��l �����4ZCHT��~@t&�Z��U���I;�Δjkg�.Į<�,6\�{0 v��Eg��d���%�c�HY�Zj.���D���lɧ5苎���Ū4J#!O�q3�a�:����HY�;)~C��������I�J�.IKvk�Y��I��g���0K,�d5�����g̡���.��)e�V����1��gF\X�l�T���72�4m�]/�G��a�̛QL��#tm���GkE�� ��յ�CD,�f-p��3)��f�6��i�����*�yIe�$%ҖZmSe��F� ̉�W5n"bŵ�]\-m(:��f�iir�ʩle��)vڱv";��?;�w�'��&�=ȕh�	�G�ŧ3��g&u�`;��Wi��Pv}�ѫ��d�pG0��' ��{�_Fa�}����X����~#Q��w�;k�9ӥ��鏘�Wp,gYC��Z���f;���{���i���y��b�&|�T����	0wD�<��N9�'Hp{Pq�Rl��ݸ�zpr6��oM�T�[�z<đƍ|�����!Ų�P��{W�z8��G�!]^NAkRD��RX7|��7����7����N�ɕ�9ӂwKL>��0��c�����[�h{�5+����;�b*��A��ٌoyi�u�{����g������ϓ8�D85I�j��_W>�v�M��+����m��b��p��L��Y��Tt�"4���#�Z�^�Oɏ�԰����>��َ(s-;��I:����w���[�X��$Ǭ�%�WU�Z�Nc�$�VC�1WiǙ��9���/�60�囀�ך�*;il���ZVDw�:��c%��}�-m�=���{�
�@�]k���~:�Uཕp����Me���,X�b����pZ�;ߺ���b�ֲx#���*����ѣ���5�md=E�a�An4��@jTB݇����[B|�S�L-��}�y��v�����ٝ�L��#��"u�R��!�w��X�,5�;$�pER3}�luD�{�-iHqv�f
;��ʶ�p8W�3�O�=��^�����ɩ{۞�
��/΅��;��^��b�-d�Gy��P� ��� �;��Kf[��g���J�����nVmu�v*:��R�Ŧ�xF��P�<Ax�%�%@^����f��&��3�""�/|�=�/#=�8���6���}�NG��;@�:d(����̘u�O�����ϣ�ْ!�r�W��T�����R�v�e��n��������(�Ɓk�q�J����B��pnӒ���ѧX����~��cꑅ�*�fV
�V�_cZ0�O+��{���X ?�T�z`�1n�mfV+�]�u[r��1���,�M"y}�1z��WZ�~���,c翷��z�~�y߂֠�ږ�h�v"�k�[8ă���'�R��DS� o@r#�1p��ݼ����x^F?�؛�&e݁	�^������;j�N2ܧ��m�;]�ɂ�Ѣ⛥�R�fV�x�Bn��I�������繭s�l�p|�h�E&�DW�9�G��͝���?O��5h�%tx�i	[L.�.%�-fl���ø@��W�o���kH�5I �vz���ޏToA�����t���^m�E�^��,�NT��)T"y�@��	���Q�1t�4V�g�����y=�:�X�I�h��4�� "$as@�9+"2�f�ni�6�r�,cr��f(Y���q�{S��a��%�¸�]�{�Z���a�A�qlF��	6��&�9������K^Tf�pK6ۻX�%Wwkw�S��#x�_�ƀ� V���~^���)�%�N!��Oۊ�˘�=�#���݅���� ;��<��V�M��G�� }I�YJ��zo&gxnbŋ,[�n,�d�Q���F����o|x��9.wY�EL_����s��o!�k�=�cۼ/!r��]�(�b
�� 	y�o��O�_ߚ�'��s�O�����۔�0���PkT������)1�MvK{�r�����;��/�xfK� ����f�[���دx�wqa��V�������0\2G��ȌMF��[*k*&�8!����Z@�O�C����s�]ټ�z�w:���թ��NӇb�J�ۘp';x屔���w<\T��EQd�J��'�]nlj�~��^�_�Y��. �O�8 �*.K���� 9��d=ǫ}x��We�+p��R�Fψ�C���t�h���,����6l�"�ѡ���l{���2t��IY��vK1ܐE6> կf�Xs������L;����c$k��q+�_t�W��VGw�@�@m!�h�slUی���N�x�9�L5�^-]am>W��ol�]:mwe,�zLab�Yl %0���^�7��w�>"��?p᛽�7���1���A�5�&&1Ŏ�ˋ��ks8C�c�3�T��x�|����h�Q�s;l���Uq�i2-���4X����6�;.���9��)�*ζ�e4�˪v� (ce�H�g%E�����$�Ԅqt�(�0L]���RXXLB��Ց�!�Ԗ-�����.�RɍF�q���MA���j5� L��̃`��&�j�L���ۢ�f�1i�����ґŭ�Q�j��#K�Ir�c3h�5`�xU�3V!�Ο� g�;T��ң�0�ow6L�ۼ/!g�ڸ�S/4�/����ؔ�IӤ9�NZ�2�� &� #��W��A�J��$�4x���l�$mf��w�Ŝع��.F�1 VӢOH��a���ƶz�� ����ZՖ�^��TU�X���f�l^�&.�b�׎��B:[��L�PrIO�E�27nk!���(БÅ���m��/p�Z�{3�8L�ۼ/!_��uq�)�:pD��R^����F���pEpj������O���N��7�p�'s��������m\�Y"3�mÚ�E;�����^��H�5�����d6G+u,u��\r0n`�iZ֕��Ç�*o������ �'$��� U'uF�5����.�6&g���V�@ ��`�F�5OcZY�(؟a�m͗��.7��nn�"�����J�p���l*֟��aB��P�����\�&�*�^�����jb6ʦ��7̓&BYe#c,�B��>ق��(���ׁ�}�����w�7B�� p(�	�|���3�S�rg�U�؋�S�rf��b&�����`�����8�����O��|M�D�0��32%��f���h,|��X� <��|���ך�Ow�XθpXU����]��� �8}d.�D&!�T+�)p�.�/��]����]���ȗ��� ��g�ʆ3���R//�^�h=�ߞw����_��bDhP�cU]X�c�-�S�f���ٛ7	�>TKY����}�g�����7�D���Yͫ�b�����fj��Ռ��}�+��r��Y��uk�DH��d�܂I �]�}�5���w\�wn � �d���a��5桌�s���e9�b��*>y�D�2gbS�y� �z�Z'�v�o����)z ۬)��pl�)��h�.VJ����dAR�vt�k��o��vA\LsP�tF^�C}К��P.P͚phSK��
�cr?}��	k�9�S�����ы^>���g��~Ȇt�n<�l�.�f5/�h�Nwk�+ɳ�:	��{�Iͪ�lԇ$/���ū�����+�9�㳜k���n�D��C�F��W}N��Am�8�þ���ٹ��m�yԠףD�gqj�
�ͮV͖�����|Ns��S�\Uf���By���d��S}wB>�mQ�+���X0�l�Tܫ��o��W��2Ψ�}��30h�LQ9w�X�HuBN�q㫴�#ԃ�U;sd\oW]�YȞ��77p����V�ln�Z*eN�ʞ�˽xp,��wu��)[�֗q�+/ya,�B�W]_���9}$����.��:x�S#+8��"�+�GS�i��C�O#8﨩�a�����|-՘�b;בث֫yks����G��[�]vl��rx9�"�V��y)�`bZ���4;��Oz�5��
Yw�^��I['U�si_ ;���ˌ���%P�j�־�p�R�e���
ɣ�\e����އCa��6�U�0v�Q�*C(�4�@ZӘ�t�&[ĉ�����m��Wi��v��۳ַj�&C������yF�ӣ�d#g�>Ė�Η���Ɇ�趙__P��P�9�m���>s����*��8h���:16� �S
uV������v�\�U���;��!���݈tH�3mgR> j=k���U��ʛ���y[����ߘUTN��(,R �SUL@SE#�SXQZ�F*�*�bZ[,�%{|~����||{~>>>>>:���ʁ�
EJ[X" ,����%�x���뮺�����������$��G
AF��Q��D �+QvI�PDQ�����x���뮾:�����||||wd���ys��)�&�C�0������T�T��0X�szqǏ�ۮ�����������ɡDT_(6�dZ���`k�œ-X�^�T0T�i�UEPPU'�B�,IY[k,�ʑJ�IP*+r3��TYPD�aF*�dQ(�$��Aʔ�/$i�^�)1"���2��eLIZZ�,��XEQ$P���$���Xu+M8�<���Ă�h*�2�
2�TF�)���BPSEDO�R��Ab���}(U�P�22dD��k��gu���vJ�>�v �-2���xѤ��B_1r�����fy����  �(۰v�;ݽ�n���p��@i�*.�.���_�v��	�;t�����X�N&�̮���8�(�K٘�z:��U]F��D�;H.��d��̠�!z��շ���O���ik6bF`��Q͎q1xGa�LX�5�iM�" ����[��qDf'$be'���[�t��z{Ez[��}h�(�yֳ����"1�s=�;���_<�K#_���)���	8�}�3��'����ÝÂG, W���hd=B�`e����Ѝi<B��ؠ��r�A��?~_�˛}�B��Ϡ��:M��t�s9N���w����w9�����ug	��(�:L@[.���$H���&'7݅�ݶ�[�J�.������c���ꌬ��О��iһq�x���N�@�X���d= ���3���˅}M�}��)��3�O�l���Ye�e�,��T�<����W���na��f)��sY����簩o������=��vt���m��?4G~��fE�^���d%�����_ܕ�s̄�.������İ5lƯ-�Tn�˥2挻>�o���vdz�<���\���=�������D{��?G�_�Cb�3S�nw���/p�D��x�u?]���w~��+�ؚ":k�,y��pǉ�쮡B�G��ߍ��_7Ho��F��i5�!�UN��A3.
\^��g����[�T�;sb�Ic�"�Ñ2�T�ݩ�'�^܋��/a`L����3)�}�w�ޟu������;k��q�Vie�0Y���AK��2B��6IU�kdm����AܭՎ�s�#���\��NA�ɉ�w$�3+8Ŀm�ޮ�����8�=��@�ν��&g+�`���T;�v��Բ���"�͟����t t�T��2��|�Ƃ�6�P�uZ�y�^1�PT�zQ�]c,H��,*[ۿ�dc?�%�P,��e _<������ˈ�q���m`��\g]1�6��[�J� �Xi���sj� &�n��X��VP�A4Űm�9B�2m����lX3q-�Q��ؙɰZF�4й[FsGi`"��CAb��t��jX��5��j�ZRF�ƚ�X͆%���Kfeh;B̈́�0�[��b����-]_��#�~�;�P�ɵ�ق���&hn]Dc����(Z�<�Yt�kg'���Ds����p�a�P�l뚾{=�S�sY�l~vK��j�og��� �R����e2�T)@s%v������|]v$Tv �An�w�]��u����n:'`�� ���6FD�~ό�x|kx`�/ق>����o��Rn��U_�t	�A�z��{/�2=>��}��2e8-2�L1�.��#��a�#+�x�r�;s+!� �S����~=5;Wu�����qG�Oa �B�>��}g�U�^�g{��'i�8:�c+��cj�5�1I�y�7��y��uߟ�(�l�m�������@�T�՚�;��������G0�X�Q͖"�eu�G\���m�F!X��T���7���fF�_�9���H�/��X�>��XqNu��G���I��>�~�w���6��J��`@	��
��OS5�W���߃��`����]�m����°�$l�y�1��7�,I7�zĒ��^�+��q~]��,�4>�F����ɾd&I�,� ��qŁi�rG��u_�LT���{�lqg"����A�b��{LL�:�Y	�/�4���,��9��=�}rL�3����Ӓy�v�_��y��j�2���sDy�����C#����ƙ ��������Z	��gE���;��߸dL�}�����ͪ��{0R�$�2�	����2��d�bk��I&������z�n�/�8���v@K�AN��p�%�N|O"���N#VX6.��fWY�Vl�A]���L%�e��R�l8p�eM��	����,�p�x���J�Wr��۹}������޶�Ɨ��F�iS��N�ؽ�٪ID"5��+�t؀EZ,C�&M4{A���3����T��˹�*o;85K�x��^�-�p�A9�9}�-!HQ*�������2���.GK���Ō��
���4woH3&uP�t�&�C7����q��i?�5S�;�mН.��]��mH��w~
�'Na���,X�������j�.u���������2>G�фC�Q�n	滣������sG'�k���
7U}���'�:n�8#�95jE�l��_����DN��})���cԺ��{�uɉ����cY�O�֋]�o�k��m�@O�0:�L��U' ��-��ّƯ����َN�w�������1Z�����R�n�0b�A��4L�"d�j�p���7��ѷ�|�#|� Ai�5Zk{�{SW�u�X�![sH�z���!c\8"�3�dfV�2�'"Z;��ݛwЬ�{����mr��˯hD71�H.FJd��R��!���3���'��fF��D{�17����59�1���^9¦�����wZv ��&�A�NA3)�����9O���%��1ӂ�eÌ�����̺���� ��H�W�����*�E/LHtJ�ي^�})��pY�,�?q�Y[�8�۽-�kk�w�w$5y�u�cw� 2�@��˘���=���˷&���bň��")ݎ&T�i4��A�*v��Q�7v�˫��7����g.��8��[�j1�D��5�}=i��8�e�{�Ҟ�*�[[X\r�:QT�Xi�����i�K���!�/{�)�g��,�1pA�p���wb��YW�=9g����Suj�OTG��Tԅ�&�927I�̧�QsS��_*��K��l�Y���a e8q�t.�o���2����@1�.ˀ/#qsւ�%b)2:SL�~~4Y�~6{�{;���x�B��츙˪��b�B1.�D*eÂ'��s���*QF�ݱ��D��Z
�;c$y�EW�|{#l��]{�Sp3�����;���&]��r�r��PÒ��2E�g�Zƥ��y�7�uy�����;,")Ñ�wi,{�{#��d�&��
�%ѿ���>��ϭ�N
��3>w�������0�Kz�bu��n�%=��M�o��A'�5y�BQñ[�mn��w�HwHq�F�����.K���GCm�[���G]�Gm��X���ؖm`Z𮥰,��h�Q���o@c]%�+0�%Y���m�M+mX�&
��h�Ers!�M�(���p�ɨ�Z�v9T��h�Dʆ.p���ivVQr� �U��Ԫ)6��s��Ma	��@�3B1Ƭ�7Y3?�W���|M�.�S����?nW&]����p�	�S�RmHL��f��W.���?ww�`���䥞�^��E�'�p�ޝ�uD�]W& ��+��mopŃ;���l�a��!�D�p$ D7�$V��Cb�:�l��SG�=������i��)1c2����u�W@���Hmd,�!�9-�UNS/�0�n/�D�o^���y7��̹�z�pl�AN:&e3ʆ!ϥ7_i�w�����jdHu���O���;��EN]WGdZĝ��q0�g�����,t��7n��v����4��rAq&꘏bd���3����+�_N�,x)��6Y��NŪ�]NMuu_�'����Gi���kR8� �Y��6�]k,J��p��bl��v����N�����o]tE�\�6O�5�k��K�b��� @/�E�U,�D"G63� .�^�}�*�^
{_��m|2wON�y��[c���Yr�^Cݴ�ʘF���^�(n�W,��;0v���?�u��VO���bŋ8��T�@S������w��.��< ͠�d�c �C���z��M��#)	4@�@K��Qk!��;�74/?��mv������jS�E���	�N��G�EV�=�΅�5���S��6w�����.��`��pN��Wҗ����j��"������y��)^r��,��]�B�݄�:ɑ[�=^����A�A�9.IrH"a����^��� �y���bj�|�|�߲��	.ܦ���UګT��t�Δ�9!��C�U����ϟ�{ae�}g���i--�7ag��'/�|����B�^�~ڞs�A�_j>{v�wpN6"�P���]d߽b)N
@�*f�f��z˿g7e'd AN5�
����V`����<�J7�x�A��ب fW�K��K��FlQ��4����Y����G=�z���هx��/��ur:�Cl��\�qy��[[qQL{j=|�;|�/������O��c�1û!X�.e��:�*�t"�� �H9I��E� L�xd&aƵl�ܻ���pŗ��!m�C�8^wb&Y��G�VV�9�{�j|���:u\Hʁէ	��$��(	�<�H+6�v����U��i�׶�g�u=e\�5�g=�a��,@��A1qI��*�-�i�p����o���з2�b׃�P����X�8�����i)�aŬ8)�0�E��z�� �3)�̧���׮����W[�8��<<��1z�a����F@��؋�pM�I�x>��??���y�=������*mr�y��s_{W5���t�b�i��{��N1��˹�ň*��Oրߏ��ZX�`P�x��&⧬������ !��c,l���L�RpA¼:�����^-����X���e{��y�ʛ��O1`A����m�ު�Ic�%b�Ѓ�s-t�9��j�~�<�;\�\�K�Օ���m}�p�X.��&2�����w1~�#2Α-�Y�c��!����X�h�o'R�s]8�"�m��=j�;�d&nkQ����Y�+���,Rj- J2��W�#g:_tD���0���FY��<$8�b$�1Gq���i�F8��	�&w3	�Mlf������LA1(�8,d�a��qu]x���T�&o5�y��>�i��}�&�
�5<	0��VC��g�4�	i�Z��4٥���NR�n�ǕչSq:	�3(;�p��&w��ȵgih>���L$�e�8 ��ES��A&y�.똧s�f"qTNg����e7���)2yˈ����TpR|o��4����#7n� )�2z���7�W��Y�r�� s׽OWU�D��r=N�!��
��wɌ�"�&3*;g�Ӣ v
>��UG7��O_T���<�4�#%Ù!(p#��g@F{*��/�t��0Ce�J�C��.��옝�`�~;���ͫ��O�[����4�ո�� �-�C�V�Z�ٸ�e;��{�ܭ�ܾ�]{����w�������_ln�eDjM�ڔ��QyF�}��4��m�ض��;��[�6�6��OY����p��sMܲ���|)ӎ�X�U�2�i+�u��w]\	�J�+�oR7"��&{�纤K��=$p�Xpa�*����������˷`�h*�d��v�5�Ӣ��ï<��&�j�@yƏ]��s�:1��6�34�"��/6oK�h�sr�gf�^�uM�L�7� �c��+5ut:T�W��	70���1�v0�L�u��ηَ:d�1Cӆ�����^�k���r�;�j�+5���W[[�fҔ����C5�v������l
Y����_kQ�W8έ�����z�@C�L����J���N���Y ْ��OI��c(����S������}}5b��V;��!!�p�B�qSLO3��ٯ_?h��S�������^��5t��J`Owo`�����Ikl�9=s�+�$$ ��ĸm������chc��nP5ۻ{-��n���\hu�̨�W�����2�i��s�'��H�����5���Ϊ�熲�^��V�ά�/Mmʷ@�I�Ew|KV{2�Vy�ECX&�\=ǫ$S��$���N�����꘼�Z�Wt��=e�S3��k֚�I6�)w|P6E*��M��]ڮ38�t)��ʆ�k3@�����k�n:X��>v��e^^����a�s���_+=�F�	����~�C�xw��)yO�;��O;�ʝ谞��x3��Q��c�ov�i����l�c���u<皷xN[�U ����(�b�,������6��X
���V�F���x������]u�����>>>=�ڕU��g̬�E�5P�����%`���yd��z� 訪�A���=�?u�����������)�"������J��
�NK�O
��iCL>LAED�L�d������]|||{~>>>=�SECDO��h
�h��* �/#�*�a���)e
��,ǏN?�n�믏��o����D�W�$PX��"�}�)��"j��,���X��U\��IK�a9�G!�)!�%E�m�"��QA��*��
h�i�()o\:��4RHDD	T��	�����*�hi������"��dX# ,GN2(Q��h��(,�AdJ�!
�|���E�P�%V�;iBz�BU#0Urk����
Wz�)�֚�*b�1&k4lQ��`m��i�Z�,��<C^R$J:df��5�De�$�Kj��[46f�Fk���6��-p�h�A%��iy��.�ƥ���ƹMD���\��f�-`Fh��Va"�ۨM�!�i�.��%�;ieW��	Fm+�]jR�/��]��2��@����h�`�[Rj�ܘ�!��[1��:^6�M��-`L�e3[���ͱL�K.�%%P L�ѳi�kk�Kn�2ٵp����6���֮�UL0��YbBc=���AU�7�u�(��f�����Ѻ���X�����n�AKv�2�tٮ�J�K0�HL\�(Y5a+H�� �ݯ_%ѽ��L����,Z�LG����Y��v���e�����[xьrͬ)�Z�L0�qZ��4��n�*����y�a��c��Vu��Å�ή�V!Ri�Y@��b�s�M�s���b�8�V�icH���f���2�2D�f��V�.�F�r���%�HZ:֮ڂb0�vghM5� n���@��Z�2��R[�X��.燬Ь��Jk2�ݝ4SK�k���!jd��ٰ*�v"��ĵ-�v��Fc�JSUFm�¸�q�qK�8�,lZ��6��CF�(�\��[�:�+]p�e��t���
\6�<X�-�\��U�k�27M-ݣ�s�%5���[,+6G1��x��,),`���6����A���4�Ư�#Rᖤ�N[LQ4�����KL�D�i��3,m5t���&��ƮD��ݒeG]��M.�����iKe�,&��՗eb�vu��k�U��	�(M(�8�c@���mB-���u&�A��"�6P�9��ʲ�.ѳ2�׫J͇94y�J3d&p�1i��,�7,�(�veyr�,%p��2�aX@ֽd�d�u]cpp�?��bbM��W�k�k�0MTƅ5+\k��������f5FWi�9If)�Y���3n��a�.�����3Ah:Evƈ�ڛB:jAe�܀��h�����a���-͹����HkK�ML)���#�� :0;a�Q���L-��m�[Y�]��9I��
� 7H�-�C)4��Ƌu䦤a��'w���"%"�4L��~N��kŲ�Ub�U�˗n&��V���u5Jf�2.�g~
~�"Il��L���&[���bwx,��)��_��d%�� �0��nDc�]��A�\T���w���D"=Ht�>e��y�{�Y����d"�p��Lj�n��ʘ�gk��2�521fE�sR��2Q�.Dy/-����wv��gݦ:��M^���x�fP�3ɤ�kd�p�T��3R���R:��\	�gijL�ss�G�x,��)��'"�}~t3=��c�j�F2:�y��!� �c ��p��eꓜ�dc�#���}��ޚ�l�8!��:�cK����AY�YS�{�Z�.�P	m����}~��\�%a�e��!���].���6�a��W@��źg�}���~���G���	{ȗ�	�];]zVMS����H:�"�ue�򁍓�Af�ID��=�B�Â6�E��:�F��A�}0k=�K��i*����OY�t8��4{���o�Xi�#���4^|�oQX�wG�
�Z���<��}�(��c�0�V:Mo��
�����������%sMRg���9p����V'�YpA � ��%����(���4�{9�|��>Lj��z��wC��N_6W�}�P��j,�U(�Cl�eR�y��G��;.�� �Rʝ]ڲ��:�q	n3(8M8��f�����)����1�W�yG"f8���z9��Y����=��wXq�Sq�Nц-2�&%O������{���~ߜV�6&s.�1I���2�nX7kb���n-Hat�\.�U�s\��G��;L�� ��c%�ٴ�{�	dzr���2սh���L@����p�e2�UI���3d��^f�Xm����u쬪Y�w��k&WI�3N�p�I#n�p�]�&��w!Dˁ�M�&}���0`��|��%��h�Ձ[��}0��=W8����S�bu�«��w���7K�^�4�6�|��9}����s;��1�crg>�~������s�L��1�@;���
@�-!�J^�\��{9� ̾�����n�Y9��\�!f��-ց�!����i2�S*�)��ÐE Y j�_����6ŗt��V�^t��[�눑���1�v��Dۇ4B2�FR�ng��H�t	br���3omk%�C.(�����jՕl��e���R�7SX$�Dv &|�H2�1q���N����q}�\�%�odl��0�^��?����#�?���r��-`ǜ�@#���RU�ؐ`�-�^i����t�AY��l�8�"Nˁ3�jm�ncl&B�I/r�[et �c2��ʋٸ�F�|�O
��iV�ՒrM^W��<��r�#�p�=J����ý�g�Ď��2�S!��K��V���0W:��f��ظ��i8# {8e��M���i������ɯ3�߆Jl�F,U�$��;|�*7����Xsd�3�Qgmw�V+��Z�+e�Q�{�|��ſ�1�c�g�{��Ky���BːM��!���69�gs�۽�ެ�*.�3�'�v#���<�M���Ri��>9g%��I#b��=�JF��*:ʶ��p���-م��M%!m�J�	��8��Z ħb &TL�qז��N�.����'���7�(*�CA���>� 
�	���v�L\b��Hn�cB�ƒ �wcu�������b�!��!,fE; j��S��ٗ���c�\3�[m�G���T�NZlx�q��Ț���"_��u˂������i!1l�pD�i<����C��2b�=N5\▖AZdrg3)�^ݿt�����O-���qF#o����� �#ؓ�����*]Â&z����	|d)2��z3t����n/�k�4Y8"��ϯ�2�p#�7��`/u���o���w!̋��(!iS]OVԫ9�pU��kY"��3z��o���zIa�w�+s��f���8A%������[�>�˯�Q�=��q�|$�,���Y�nh�Ґ�6�j�Qs�����^35�)9���_:#f��p\�*�2��#<nue����$�p��;[�±�iG31�Z�9���f3n6�,cV��l8{i3��.+c�찄�+-��V[FP��4t�2�w3vMՄp�R��0al�RYL�Ը%.\��J( ��-�6%�����پ��q2�i��cڪ�f�0�at�#�G��J�������ȝ�<�8 ��@�%�-0����u�����s9�P��xT�1�H�M��E�i- ��!Ú���U�O_�UO��1v;)�&);��޿��u�[�GxL�>�i"�����	����g����N0���2��H��
^��S"���������
b&� y�p�v-T�	-��+���n��q��K�pp�%N�+r�}��|^�s5����H��0W�D�[����L�S,�I{��Z�[�&@̯Y��U�tH���v���ww%yk&��9�,�G�Ù -����~�������O�>\i�R��M]�	fl�^���fY��m�K�8��W2�]m;��VG䨟���6cL�U^`��6�/�xP�=��ɧi�lb5-�33e
i3I�O���j��m��#>�=��\'�l�T�#F�ȕ�q_�	wx(��������l��x�G#E�t;dU�����������HyWB�o�����k�=\�u��� �#n}u���V~��l5[��)�t���@��j�9>��k�W2>�}L��
�R?Xs���f�J��zޑUV�U����4K�I�w��KKM��Vzv�d���N�Jff�;����ww����3���c:�fc��ٞ/��������܇�s^�J���,��(�é���K��r�du<ѨWL��W�U�>�ЫfQ�in璟�Ğ�w��u	�(L�ST�Z��9'Q�1���[��t�Ws��"W���������.USO�����I��������t��=2(!��]��5�g׸5B~�}-�#X�ڣ��(�G^Ә�W5J��+��j@(z�m3�n �bŋ���}qZ:j��T_����x�U6m`��=�ZK~�G��mka�0�L��͟_h9b�+C�t
b|�f���\��o�;9�v���0�6�M���ʪ�"ꌉcܚ4mv{t)��5osc׭�֮�B��Ըwz������T�[fp��]!�$�ٶ� ��q0\0�B/Ҋ-}¼���	��z��g�.�A��gW�e�<m�^�޷fYoT���M&��=2��LbhI����t��r=wLwgʙ̕kS�p�˹#]4�a~�s�����-��3�eՃ5�g��^��E:rP�{�1
D	�}�m;�@F�ei(��"�^U�E%��|j�h���E�<y�o&x�&&g�U��x&L�gz����V�>�h�t!���)��*�h�A'�~M~M�z�#g�sϸ/��FgW�KC$���������f�}3�loH6���=Vη�`�t{,b�HFS�wOj�ug����Jz�&"j)h�&%�)(��O���GS�j���d��)4��A`�J�D��ьX�b��X�-���SL�.<�>����S�2��^g���FP��=�lEJl�T�ɞ�T�އ�%�;�� Q����-4u���^�Ick�+�Rb����c��B�v���s���!�Be2�O��)�������/x7��g���O@	�1i�z�$��*3�'P�n#{6s�z{]FgE������lY�n�Ϗ�Or �+�]\���^ ���h��	�{����#F��˦]��,cWwRa,І??��G<�;��C�����{���Z�{�o^�Ϟ�/�6���F������7r�M:@��Tj��i�^������:��ίp�M�3&]��wCË�{+�ޏ���v+#��>6�j���ƧԜ�Y{����_����s�>Tk�^���6�-f+0��0�i ��Yk7�0��~�c�����L����0�m5^,��K���Ķb�S"	�ـ�ŪW�h2���ѵr
]2�iv)L�P԰�Fjf�#`UR�.A�p�Z\b�X���ǩ5�L��gd��1�6�K��`��^Ua�Q0��,�[s0#jJ4��93��su��å�
#2�0�[\WFŹΡJ9@�)า�.2�՞]�N�w���|?C���I�u�W6V�4�0�(Ě�ux��6��LJ�w�,��&�Be &K!�s�s���P��ᴱm\��v�����3�4��g�=�I���n�rފ�)��w,�����f��^��zS12.�,[��;�d��-�m[[@7���]�r��ѓ��D�g���2���fv�� W�m!2�]�|��l��|q}*u	�Z�g=s�������Ꞿ����)�'��@�d' �v��h��*t��u�)g�G3{�m�u��{�����2���h�|�w������.^�-���b�bji�͔k���Υ���l�*;�M ��|��2�PY���p�~|��v���B{�~�<���bҐ�@L��$��N�\�XƼGƭ����Z6�nS*�����ko����F����DZ�3�]�=j��hI�x�ȟ4������,X�b�
<7ɛ۵�^��X�=y�����C҄�E�c�Dm�<k��c��UV�T��t�ݽ�Z%�۱w�j�-�[�L��Jvv�Z��z��Q�fV7qrI��f�B��IF�-��;�+�����j�|6w�=o�'j�=�^��+�q����砟F��y;9�kD�^a�c;�D	t&i�lr�~��$����,�six;8���	�x��l�ņRc�"]������������3f_&���R����׽���FS�B��l��ɦP�ƻ�jښ�������C_Ew����"��}^�tI.��qU���k�=C�����^��Fbt��[�I>��*�%�e60�����(����n	�V�ې��p��&�놻W$�/Q�:A��I֙�����#Y�!樄Omfk��ff:�k�T�o(z���t9|dغ��Ѿ��y�h�W:���ClœA�aT�ۊ���o[㶐�Z�V'X�.m�L9�z;zr]1ZSx�����V�˩ԥ:4�Z�boP� �;�� ���:s�L0L���u|�쫢l�2�'�dWw��q�Ҧ����ɱ��b�%�ՙl���ɻ��:�	w��-f��J[�]c]��a�t&A�xk�q�!c�*h�7�l�`
��h|��A�C03�<��їWG]�3��sg6JC��ȭ�u��D��$q�fX�j&7zovh���I���J��6�n�7P����d���^-\5�K0���ފ;y.��
����fL���j��:C{Ϯ�7���oA�W�5�%.�d^+:�X0z����O�*S�]�ba�\3���<���3�`=Պd4/�z(�eh�,ղ��γ�Z�|�=���T�\��Y��(�`+��q��+A�{�TG4ɨ����M�v��O���f���f٫ш=Al-\�[�po�]�c��WG�g[�36e�X!B�tA.{C{�;٣�r�y�0<�%���И������Ǧ���i =$�gr$!��X�`�U��Oyn9���q�H��^tW{'�ی<{�W����o&���@s���;� �U1un�sɃ�p�l����Vq�ՇQf;d��ƚb�@��|�%O{Lu�i4��<��d(W���_���Z�~Z`�)%Һ���y�j
B1X,Xj��D)�hj�(���S�x��~=?|~:������||u(#U�cP��~�c4�Q�*����()��$��x����]u����������-"QII��ɪh(
i/�NJQ@�=<z~?�?u����Ƿ����5EL��UP4��IKMR�PR�!�)�ǎ8�~8�u�_ߏ���	Jy4��
i�R�iV���ҥ1!AT4-!�NM ��iZ
@"�B&�p��B������rj�������� P4%-�4�BPХ-�9ʥ)"F�F���)��))J����"��PIJ�
�IXTed
2V1 )j�V(����h+�:�X�bŉ�ɧ��˗�&��uJE�R(sM8>nm3ڹBetқ�ѷ��Teߘ=�sO���R��v|�;+3©0�S%�L�C��5S
ܾ��a�O+��J2���'�9�^�
�����;��ڞ�~�Iv5h�~�j�IF�h�4�nq+��\��7[2�6fN��P]��;�"��Z��T���+ӹs^��7��]�s=���{��\�1Kbf �Bg�]�o�b'�Gz7caKD!M���Jr���{���~{��M�w<�)�w.2�(%�|�(	��h�|y|�C��_�@�(_�2��4�/�8	��O����	�;�Q��f��������Z�U�U����VMWy�t�1;����r��~�-o^�Vz���-��f~@`��÷�M���T�ynd��ٵֳ �TW��p��k�"�T�T{?F11��~�;�/��u�Lީ�ۍ�qǶ�}0�o��}����.��[Й��:ު��{��Ξ�Ąc��^��l!2������B�GC���KJA�`t^<'���u5R�N7�^�p9�f�e�G��*��U3[@_/UUx[]�&"�&�WgWR�@��k��(un�WW��������j� "�z��|+]
e�6�h�eL�0]��&5o����Yw�tz42yQL�^>�ȻMq���%��g��4��+f��2j2����Boc��h�!��pj��UI�j����xL�QO��˪����0�c��[o<����ˇ����9l~���N�.u��Ok�)s˜��f��y7�̅�j���J@��q ����)y� Յ8�0pk��� yAAs���a�S��N�u�;�Kx��ŋ,X��5qa$$�<:�:h)�(�l�� ���f��lٺ%��i4��
PQ�6�T�e/	r�rKQ�ʥ�VXb⣀k�
���cj.��DM�ͫ,&]y�]��u��5��l�QiD��1[i�a
�3B��gWSQ�،"��m��
���Y��E�Q9V+4*6�[�:�f+�n[�p���~���?�o�Pv���)� �y�CM^+\QhmTl"������A)�y0�S)����UW��~�������7��ա+
b� ���1َ9F����c��گ;
�����j2�E{�-�g�����^_S��.�_��Bff<�R����g���Ɍ���3�hji�Ji	�j��}�=�'�ϲ��&�L&v�U^ts��$�=����_)�>��ʵ������U+k�Z���oѱ�{:��O��ѫW��e�GP��IBf��s�A�}�J>����X�؊�Δz�v3+��E�����!�Yc)���A�Db�-�0�S*e*�˧�e_���9|�_'M�^���ֲzEB�%4ʪ�}�'�Q�u޸J+2A ���oOU��^��۵��b�[��Ȇs�غ�l�
�}���['�.��qkc,H$���18�2�} ���,X�e���X���o/;����ۏ>H����\�����w�����]��[t*�Z���tA�O᠒�*��g���Q��¡{�ekUl	t�yN�z��� ��<�aT�ffS�^a�f��=46��;m6nԷ��;
�̕�K^8���@�F]^k��*'.����1��I�F�G�Mkl��{σb~|��G�#�	��*�z��gKG,b��7�B�ʹ����3v���?I��O���xj��w���؋U}Q̛'/^4^��m�W�qc��v�]���� ���$�%��Anz�߽�|z�9p�3�{&#y_a�m�vW��V�mw���~ܶ�h,M���W;�Z��[�L4T-�#����V�擇� ��[���na�Q��*�]�T�\k��p�,X�bŵ��}k7��>˨���C�4�3�2�eL�\z�w۴�^n5�<�[�����]�,tE����������g��RJc�$,@,L�j�d��v�ۘ�:��(k�\{f��n�8�fr�"K!m��T���U�z�V��]x������5sf��3&1��:k�T͘�+���w�{&�r�eK3��woI������TM݃/��3v�[u����	���n׽P�O�D>�n���5w�x`�U}Q��6�b6~������V��z,�)1�砓B�C��I ߣ�v�ՙ����$&�%�H�y��֙~�N?����5`�o�7o�~��~<�Qc��<�Ⱦs/Ű��?��R����)�k�t ��j	�ϻ��V��9��y��4�m���rZo�˞�F��*�7��>��dMPɡ5m�X�bŋ���<�S�υY$�����/M��1���8,F�ޣ/�8T&30���axx"}v�l'	��k��U�� �m���vr��5[42l릃�}~q=�zTL�c�T�crm�k;
��\:��M��U��p7�Bff!��o73�!Qb�q�@VY��W�t�W�Z=	�P��t,���ɦt��qt�U &T̓���	t8���:^�2���=�;d�yZ�U,k���eǦf��n�;J����4�՝�
�g.��3�h@�P�u����5���۳�j�)T�4�F��N_y�
g�I~�E���]O9��� }�)�2��[B7������96����԰no�����t[������%��|fu��n3G�]�tÂ� ��wG���8q���>^{s�w���U�K�}{�O)i�_z1��|L��!�qć���Ǘ����@aI[\�*m�� ˦U�ЪR�sm8�[,��,��$՟��7^<��&N��\I`^u��j�b��`�gPt�[�-�ÚWQ�c�G)��4���ն&E�����vQ�vw8�帰p������l�v0ju�&�ֽm!��t5Ì2��jͰ3q�v*�����C{�?�5!&�Xّ�[r�ɣ�׮�Ws�(��� �L����v�2��-��w\8��{/�8X����)�n���.�z�ET�Dl�lN�"ù�C[y��,�U��P�����U �V��y�Ⳮ�;ϭ�}l�͙w�T���G�^�N�q��B�E�꥛��UI#4�lik�����kK*�	�̬]<=�)��;�1�w��W!2���O4���ܬٖ<�69ǋ��PWSF_n�p��e��2�Qi�2�oxnఉ�a����<ﳭ�.c�JgS�]��0���#���k ]Cj�ZW�x��b�'p5��L&�S(<˴ߏ^.����gdw>V�7�[=��N>�
�L�����}�AY���̊�����^�#����(ͱ�[�Қ4�,g�m�o�X��uv����,ͭ7O�.�!�L#˹��Mo�2�Mvg�;re_�F1�c1��U�l��=\'v��V__�1�@"FK�M!��N�p4��Qr�c	�[��t�8�֩��Y$��u�`:������V�VfG�zK&2���MTy�ܓ���v�W���WY��]N�"�WO��7r��w��obƖ�⪪f�dn�y|2�"jxN嗨���s5� d��xU[�g!�g��H��O�G���O-V19��3*�� �#aA��/t�ue�bG������%�����i��s�����R&2�<V.�{��2b����@O�/K�j�i55�����FJ�M7G/U���uY%����t	o�N�deߵY�����ɔϷ�� N��@���x�Z�R}I���]X�o{�]3��n�=�x�TT�,}����կ{���^��OfT����.o�ŋ,Z1�u����U��<�y7�T���)�����by�t��0�B�4�3-[���=	��\g�ZWwN]�V�#�<�;[U@�&z�4	��u���.�v��Ω�3�R�M�e���6�T��ս�۵Zk���/i$3	w	�#�t���k�E�t���%1�掏5a�'�o��[f�qT�PMq:3z瞵�Ue��74�<o���E+�&SCL�ʖL��x�rc��op��M*ۻ�/�5sL��37�"�~H�>vM���ҀyL&n�>S��̱=���;�ҿU���|���i�M��oqYSh�k����A�	�*,��޾���Y}�w�Ň�l��|n���*;�u�读.ğ
J9�}�Gr�A�z}�9υ;��U�Vo�$[e^;k���բ3�Oq�����騳�b-��ň�l<�!z�i�a	�g�����v��B��C�p�9ެ�P��P]�H��e	��9cs��z󻿜�*�nRYi��11���q��4�L3E���')vH0�:�H�O��ZK���Ii�=4�_VOy�<�n>��k��n�?U�̦�o����;`wJ;Պ�ny��Գ���ה�"j��ݵ�%m��2/Ƽ���=
Ÿ5�o #UBa2�f[��1�듚!�x_�ɭ�n���x�	�r����MT���ZN[���L���tkEu�w�;�z���Q����r4m���B�m�H�Mg��Y�ڊ����Jh��y�g=�j�r�'D��:��2�fګC0#�H�'ӏ���z	��Z�*�wiI+���E���8�ڌ��xГ��V�f��]㛳r�ۙ�D#2�t��aU���J�殺�$⻖�[=&��6�)i}S�`dt{6V����D����Fسխ-�k�s:��#�zb5S,P���Cr�N�n��;�,�]�\ɤAU�M˺�s���Ax2i�r���2�ڱz{�ZyŮ��Z��V�Z�U�uh&�M�nӓN��
�{5U�"�-,�/�v�-&,��$���8l�4�P߃��2�Hb��]b�u٧�l橡]�]Ov���-�q�|�:��gn�y�T4b�E�2��o���V��M�Em�٩��v�nj��wl�6���O\9�)�ݶ�����]wx��u��SJƬ���HS鸫n���N�`ޛ����f�^s�S᪸��������k���}��?�ۜ�T�b}���-���=�Ϗu��k��Ý(wf<���t�a��8�J�h�ӡƕ��.Xx��U�#{z���}�>����T�̣�%�>'�u޳պ]�[|�o+u�]:��F����5Ŷb�m=�n��j�e:���k�V�ض�EK9�ڰ��6W*k����ZJ�S=g�*m֍�o�UI[����-oJ�a��K����l[�ޢ��L����)��{1ٝ�aY���$�^%Zݍuo���6��C>;�O��s�~�:f��9;FX�H���(|M��<5?vxw]4<�&=Wt7���Xu�O;�|� ���=>�%�[b���p��]4G-��Ĩ��2�3[G �J\J,!Ļ��&�`�h�m�&,p�,�ċ�5ލ�V�[�ģ����TY"X���P{�B4�-PPD����on:�u������^�ߎ�ÜV��SM5�9$AJSH{�AA@���AH��PR*�rd�O���]{{{{}����
JB����*��8T�R�M5E$I�<b��<zq��~>�u�������{{�))���(+dT4�E-R�Q��"�~Br8�ǧ���������������>M#]�P����P"����Л�E��2윖�"�������9r����J��PrI��Y�m
�AGt+`,6�X�|D+"ȰMҪ���X��;�H)6�q�PSL����A`�6�c'�*D@T@�%@
*�'-��1	hМqV@F��P��(��Mҡ<�>o'��E=X�;�eW+CY@����[c�������e�,P�P�pٶ�	u��pJX�l��i��.	3����e�-�i�䵋A�;�H0�Vd�iBW^��a2�,�	L�	���2W@�S[��W\�i-м�I��9�H� f�qXō��+y�lɣ�Д�!pⵀ��t؅�n��a4��0e����բ9LjQ�&0�T6��rHsM������c���ᆖ�"���u�`nlM�7.� ׎\<�5nyL5SMZB�n�8�K�ZZ�K�VRP䭖mi
�`���B6�MZ��iU�!��ڢ�BR���Q�	`�&��6b��nh0̰�SX���٭�`-8�`�m
QY��UʳG&rb#aB͜aĚ�! �,+	6K�H�+a���&����#4)2�CG,��1`Z�Ԧ�66Yv��Q���ѧ��ޕ+t&����5���૬f�l{j�2�FG��%��ڸ��M��f�H�N]��Cb�r�8�b�B��J�l�Em�[%�q���LK��3�ʴ6�f&�m��Xp�M=CD���:�f5�넻���+ѷKd��J�ь�n��ʍ��p-��mq-�
�(e�+�F�V�<��%�Bn��!M +]�630h��먼3�X�lUcict�XX�n�,���8a-ڳB���pG�6+a�	(%�����F�k�mtXt�� Ќ)��[M%����2��j,�Ѯ#5�ΑVj���l���%u�pˁ�k�d�֎�p��B���v��V�.�6�K�C2gSB�ƣ5�8�jZ̩�F�����S,�m��!,E[��l�p\�X�x�G#뜦]�i.Ġ[6x&�M(�!2d�Х	��f��L�ex��i��G�i^rk�B[F�LxfXa�v�X�(B��̸v�pP5��T������1#���y���7]�v8+	�����1a�ޭm�%T��%(�Xk��F�r5�Ms��]���Mk-)����h����0�$Zf���mA�	z�fK]�ZҦP�
�閕�i�J��S����T0s��bhKu�#\����c4�`36r&�M�J\Sl������T�[�Vl��-D�ʳث�3u��{|=�o���s��ߐ?��Ms���ÇZ�+��2���]M͍i��c�	�?{B�	�&T�h�/�=�Cў=B���x𖜶�������^������y�ê��'h�g~�'�	����ec�5�L�[-��aM��G���P[鶨�����55�Y�^p�z��s--S��=Փ')ΎG��w3��*�>
�+r{b��<{�T���:P�w���cE�R�68��/��~,�3C��;�~��k'�X|�OH��x��g��{�^�Wނ�H�ךq8AXq� ����k�`J�^	f�� $0QEC��x�������2�4�g<;�����T�ug�"�&f8��{�$��Mv��Be;D���>�+����h8TK6�[R/�8�"�Q*�t_>CkEodb��R��"+*Zˠ��}ܻ5&�J״P<��;u��o/9��s�r�����33!]���Z���EvOlP�g�p)�T��R��Ó�b
�|=T���|)�������\�����E>EO���>q<��b&f!��N��"V��[��P�`����o�G���9�H��{���И�{]�r����h�,@�3��Ga����3���Ε�:�Cё,������	�S�!�}�>�����H�O'Ϥ��!�	�0��3)J�F]ٖM2�V�QM�1Ḿڏ#���^|�y��i=��=�j���ޢ�"��Ur��6-���O�-��^��13�q,�Ǔ���;F��CrMnw�'�>�UgVkSuJm�w=�g����1�/�� �Ƀ��(L&���/�n֙I����Ȗ���O;k�~�[(�Y��w�7B�k3uʽ�H8���_׶���«��&}!�YF �ŋ !�s��^m>���-�*��U &PU�r%���n5��zBf���]��?dk5]��?>ӿp��������>�7�Ҽ���9���3W�9;>�EVt�7�0�Be	�=P�&�m��&hC��xu�~���CUi,�ev�8�^h�u���i<��;�k�(�h"<%��(���UL�ʞz6_C�u=i��[<{ ˑ�y�G��jٞB��'[Y]���Μɩ�]l��ףsc����Fl�53;@�MU���ywk�8M|�ޘ�M2��8`�s4�^˜����Vw��4���Tc2���R�x�=^�'/\y��0i��~���O��{�����z��*8z��)'3��7��CV�E{�^��+{l]��9Y;��J.WG_m	�׭��ꝕ���)_����m��Z��* �����U7 X�X�b���z�L�f\zfp�6N[�2�A��s|���d\�=�CO�3�i��������vԠ@�'��IN�����WXͨ�;xvԵ[,sV[��3Y�������Ar��de�(��]r���Ρ9�mҮ����ʜ��]D�n����f��ø�����4��Qпv|�������������]�CU�j�+�殗�$w[O��ܪ��aeu���."8�;�9��Eϼ2|��XT�;W 􃴲c*�e��q���sP5� ^�m0�,D�̨U�����b�;��=	��G�D��{���U��ֻ�.�ڐ&s:��L��oGn{=�3T��{�0��*T���5�t���y������Q�q9[�P�mGam���ͫ��D���*�G:|���}H��ob��9�;��:.ފ��<�H��8�&���$}n�ˣ��G4f��|Mz�ߞ��:^���Wn�]f�4�X3 ��
����x�^݌)�,V��c�Wh��].��:�84߻�R��і�ػ��U�va1���t����i���f�j�֐�e��#����k�	tKr �ģ-��4�Q5,�K*����cj�M�Th0�4rqc��i��f�Z��k��x�Ѱ�R����H���5�2�WfV�m�G�j丹���3b��{��y����/_1����~$�[q&V�]؂h�Utp�i(8+�� �f���h�`{�Ԁ�M2��n:�=��L\\��K������fY��}��UFv�7��ᕱ��}і*�F��b�Y=�=�SUYϜ<�[�L��y���cE�oT;�
��f�Q���q�J&�!LX�FtM���p,})�Z���j�%��[�s|W�j�emq����w7�g��neCH(��Ǥ:�xɲ�]�*eSPO<%fm�vsRM
���Nͪ�����O�jmۿ{�^ܷ��Ϟ�e'�~)�}�Lmf�[r��Ƥv��F+d�iL�[���2��5�f'@{'}��+��=%��>��1�ho��@�4��m�h�M2��)�M?�<��~{v����2��.��\A�q�`7��_u(;Y�*��f)6b�u�_�.�x>����w�����|ᛆT�zA^nb�1bŋ�v�8Z{3}/��M{�9� ��������s23�S�!U��A�>E�_G���}��vmMMg>sQ�Ag�B�2�-�����ϔy`���e>�b�)	�s�s�z1t��F9�i�%t��5>�T'��:���g�B�fˈw��L�]ꡣ����=`����
k޹�h-,��'�(L��3×��=[SAӸ%˂RwJ#��q�]F�)�����tcw�Ne��:�aU��-��d����|�~w��ho2�B��(�Q��j�y����1�ׂ}V�*Sf�ޓ*/�S򿡻������j���B-�g��p�^g �ٹ�ܽ~�F�_�߼��H|��\�kf���Cϫ���sC��7������ӧ~[fQ���{Q�xZ�f��^�D��X�ofGN�:MhB	ݙs��e{鱺fk<�ƥ��c�1��c�|������k������l��]-[B�|.�^b(���Y3U��Ѕ`���Ɨq��ԅxHdVV��Osp|����z#&'�|��noJ3.�28�k�N&�f�W	�C�^r4y�C��2��EvJ�K�ZQ2�q]qMͨ�L�xq����Cԅ��3pv�zV�5�\禫�B�ѵ~6,��ޔ�eL��j��\>���Θ����	2� {+�ݚz�{&�:3��k0�D!f ��+ۋ�y&�x�D�3/������Zbޏ�\�NtJ�=�҅J�BeL��1���j�ۨ^�&P����2�x)���F��&��v�｛�z���꼭g_[�\�n�Zs5��omǭ�ۡ��������ɺn������:�wg2���F}R0�bŋ 3��X��p5����[��苆�Φ�r;0�R�M�tg7�m��i�Ǌ��~ �ݡ#9t�E�w�].J3
��6� ���l�*�wH#��E��#|��w���Ū�&|wFzo�ޕ�{�V������ג�zZ��mo'j��UeH�ک��$�����]��W�UEz�#XL&�M3�w��z�8Y�;Ѡ�;�X�E�Ri��S��5O����Uy�n��8z,v��ffn�O�}B�׼��5 ���d�����]��Բ�sL�����)�O :�W��L����u��zl��u�{����ʢ���a��&����<���츗y�`�?Rl�g��Vɉ�ۈ�kC;s&Vf	~w�oԴ��� Y��x}�'�ff�Ƈuಪv�k���o���
�2��.����>�5X��#��N]�n����A�c��3_?x�r����||�M+eƊ��5�J\�v����-k�;k2@Y��duv�̶`�2�,�y�%�و�Z:Te�.Mջ�doY�їV4���gk�p�"��eŏ-j��	5\RW�hYI,n�ε!�Y�.T�9�[f�2�]Qc�C��%ChZ��*\l�� �4���:�؈��־��������yS���e�6�Am�v�f��ZX�Λ9�syŦv#u��9���~�s玟R�K/4�,A�\^�f��S��gFG�J��}Yޮ~䘁T���Jj�艇swq(Q����V�{'�i��p,fP*f�r�O~�O�]W�6Y݋EECzb��Ub)�~���_��P�)z歹��6�o�S���Ky�3\C�(�:�ŖM���]+��m�WES��gF���34	ŕ���1��������獫�Z꽵+����4�g�sU8㶮�T�u/����&����b�p�LI��A�) �J���)�Ak"C�$���=�t���&������`��^��¦v'-��W���@M�<�(n�Mu�{���g{����#��O��)շX�tc��նvv-;��+YZu����̼�J�u�PѸ�P}GP�l)k�0���C���[ �z��xx�b�^�e
���jw=��|����`"�d��d
&�������]w؛�1ރ�G��yO��}����ɵ�r�dL	��-X��-E>�����1wZz7������޳��F��8ۼ����k8�B�ML���x��v�KN�̺��f�UFM��bn�Vy�Uj��{ݏ�i�t��T�Vs��R�d��p;�딎Ь�(�e�Z�D��MV�6���f���Z���B�4�i�ٿ>_M�DeVM�?s\�������G�w�T[�ē�Yf*��������7s�@��۴}7���=���ք�d1����3v,�ji��f�'Z��U&P�sUа�.:c��ͫ��v[�m�{-��duv���sN^3��ΥK#�Z���:mp�N;}��Ʋ�I���]��]X$�7~�M�6ܕ}{��`F��R�%�\-;�Z�Η�&�b6�%�T �F�>�xkO�f]V�e.[�T�.���E�1�x��!�����0��s���fk2mi��x�]WŹ:�R�����n��;i�y�l9���oF�����`J��:��T1w}<�����#�6��	з;6�cd.�fs�{�1	]t��f�cu���ԍ�ͼ�õ��KW@�n�!�g8f��<��þ������"��&��vE� ���ʖ��k����H�0b��kw�Y�����tӚ!�u�kȔ����ݽ�D��w���n\�Z���7�)w���c2rU��d�Ej;r)����F�0(p4�������*&�v���[u���;`�A�#P�\� 4E��t\}gtY��H��7h����l�w�l"�Uө���R��V�C�Ql��I�.ԾӀ�a%��H;7��eAQl\/�tJZ�f�"�ޫ�i�7��Z_}r�[����d}1^g��'^�;nWvf�Ej+l˗��Md�����ԝۘ�F�_.=��򁛨���t�h#�8V���@�p������noe���ރ:e`ɶ�:�� &�����X�г;����D�@��ʴT_b�*���kţ
�ʱ��,Ha@��,aZԬ�_�
��A�{{x�������ooooo�������EDIM!�&OT�Hү$9|q����~?&������������=@P�
�%��v�pCHP4/.[=s��R�>��jrn}>���gggggg''��x��R2W�V�R,�!�YR��E"²��
�P����,����?M�g���������x{g�@>Be�11U���B�&�" ,���#lZ�	Z0QC�U��}�X��g[�H�E�eq���	���V'hT�
C�P�I��
AE��(���z����-��91ekRZi�Y�,����m�B�ͲTRbi��f����5*E P+8��ŋ,@,Y���lvk��UFM��g�c{Κ�g�za�	���z�߫��*z!9�k�jgno�]�s�5�~~��z��D���6�A�4����J���>}�B7V����V�G6
.*�8q��C�ҿ]ל�(�Q@u�2�Jxx�
�fl��\��ô,)�c`�,� �ic�F������>,]S�v�z��Y�&��_:��=7�ќ��V����s�&]�<a	SL��_=-ػN��u�Q��y�6nz#&�mo\�"��Z�TfZܡ�5̷�Y���y�pf�W;�PJEZF�r�:8{&���=W��P©4�ZLU漬��[�>�Ңe9���}����_ɈxN�jkG��`p�������J&��7`�**�l��v��=�ej�)�����`��p\Vb�]ӠT�W������b�]�d��I-w�e��ך}�!?,���<��=O��9��ɮg<���̉�:0��~2z�Y=$��r^��ӥ�!L�670��G�)53�Y�������X���;��(�&>�7M8W\n�Glҵ����i�]㘉I��i��T��x��_���j.[�y����Sy}���2�v�=�M���v�U�6�e	���KV�>�S���ۗ}��؜�ɥ��~�~��gݻ�O�aS�o>��]�P���;{�2d=�+�	��=xwf�A٥k9�h�$�;;bO�Ϝs����p�PމN%5h$��q��������o��ϑy5W���B�S)�Nq���+��Yo�lկm�����N�J�}�)ev���g��j�Y���QC����������oe��/����.F��P�WB�ޟ5�c�Ve4}�=��q�1&�;;�Fʻ�4#qL�� �]M��qLa���`/%k,�n6�&m�1L��X���.bm��@�͚�9�J֘�1cr�%k�een�hJ�֍�V1�9�:�M*Ges�l��4ҫrMQ��i�庣v�0 �iqe;0�
�U%�ĸ\:�s��E)�4a��\��������Ʃ���:+�ٮt���y�����)��~�
�X�
L�(Y���U�d��^����E�]bjS\�|mͿ�s����T��'ra[����9깥�R�R�����Qp����f��S��)hHϕ��H
�!T;��o�߇M+Y���O3.3|e�kg6�� �v��e	�d4!�dBD�3���{�r/&������-�����dכ�nW�ML�b}t�(��G=�k5�Z��_zs�sK�&-r��;>2�#փܷ����imcN�U�<Dm�({�$eɷ���>���j�hj���	�>��K�RD����Rf�4��a�8����4��	��`�ˈ(���J�疿�Ƿ���@zeڧ��]ʺ/�^���&�M�+���i��H� ר'�֚v�����|�����1�(S�Y/��@x׼�J�oɲ]�Q�Wb�u��7q�4�Xvk;>��T��65��u��Oz�&�1_�F1 �"v��k��r�}ܙv.�g�"�V����k*g�&\�0�#�#���T���2��\���op�͞��[6����M�ֺz���Aۚ��s�l�1e�F25o �5���4�4ϫ++�u��^����v��O�V��ɴ���+U�S�b�wn�Y8/!@ݼ�2�R�2/=�~��+���(l��Rd�>L�$�;��F$J�]��`�al�l���l\���c6S(.Is
;����S��hd�2�ed��Ü;��j�k��Z=���rd�0�MlXU%3�:܃�+�_h޹�z/�w�uǲ�y{���6/�:�}�^�"�tʭj)45L��ޗ  Zd��8�_���ڕd�{Vs͑�����7�3�U�#�X��g췋�m�;噰�W��K%�Ca}����ar��H�c��m�9�Ws����ff	��u��]���ji�-�4P�@L��^�I����O�Հ>M[S��[csx��6�Z�oRd�Ѹ�/��CX���cT�g�/5Wc��]���5=ˋ��6�n�z�g�Y7�7م��A�+��{]�be��e�i��L�R��`�l�.ZT�m�����{�\��A�L�oJ�f�vN_MUFQn.ٹ�ֵiqM���f5N�=
u����Blkw8�YT6�oq��ub����,���k�������𪈟gsI箛;��U�ޣ�Z3_(�MD���阜ɼ���{0��i�M���V|���il�T����/Ol�NUW��]�.���
�=�U��{�>d���_��>��zrԿ��ي�͖�1]���FgN�k��۠2��{,Pz�X��;����{N�q]c,z�cgш1�b�'��Nv�<��rP��ӳf�ѻ�B������ZY��M�1�L�����WY�ޤ	�q=�j�Di�Bdv4Y���Quuq)s�JKJ�dq�A wQi�;Ss]�j�;{��t���7��om7�����񄻻G���32�&wΰ��O��|H;���~~�wgzr��t{���@m*���w�%&�E�rj�&|�O���n8���WYJ-?�H��K�Hi���j��˘����u���+PH���=�E�M��o�Aǆ*�p��n^g�'2]4	j��LjSL�J��槽�	||�3nr����n�M�MU��}��|uq�.n�F�����:�髴h���ĳ�
n[��;���U�s�v�v��
Ƈi��3�h�:���3G�V��z� .}t�����A�0�>"��`4��Yn���Q��1��`oG�3)z>�ּ�gc2�%5u�6r��쒁��Q*�d�Vkc�#c�5H��A�K��͘%�ʒ�(7iSm������-�L��l�a���4�YaK����3u�H9Zg")w@�`˘@vYf���(�̶��S��CSai-�t�kM�CE��06ZP���V˄�[2�D�S����H�"�n��K�z^����{����,Ԕ:i�κ2��-a]K�qn�4�*�6CEnA�������U���vy�&��\s{���{-,�U�w�^���W�133�z�ΟCu՝�7Yǣ�y�y}�u��%�`K�c՘�^���e3���B�;���wg�v��˜���=�>�a撄��Sl�<�s͖�ж5P�+.).��We���K]�o(fX�WI�f�奨�P]�q��8�i�{�GT��p=^U�����]I�@���u���ҩPD�X蔁6�����y��8&U:���
�$n)�K����n�f aȆB<؈C���A�R�Qo��q��&���r˵H=d���a^N�4�&Pl���|>�������BM�#&ލ�TF�֞����QU�ǭ�	��=�y��W��l}op�+��_�j�V�}�ON�ŋ,Dö�����ԻyM���[���v���qT.�w�lx�K5r�P�BgI����x���p�����=^U����uCL�	���۽�/��0�=i�N31 J�Mw?n��jj55ۀ���2����\��;���2?��1ռ�w�v�|vz��B��n�I���5m)=��ý�km����a���CbۥQ�B���6�f³����K��A���8�{f�+�gP�-2����j����ʼ���Qf5�pL�b/e�o��S��j��{�S�ʇ���Rϑb�;���SW|�T�v�y�~��Gd;��gom�o44�����>�^.��~&/��hYk,k���)��z�}����ۡ��[2
9���9�����!�'n�u�U��֬{V1٤@ݰ���#��`�ͧ=��sg\�^T,��t�M2�S&��4m+%��S왫h�2��{ӵ������_o� ��u����z��T!� L{̄� <��Q��GaC�������\��(�?�u�a��CS]H�U����Fi�o'���!�/,s}�˶��#t`k�Tƪ\�֥bBh͗U���[�L��|P%���RL3�����Ug��9��*�Y��{�u��L�4��օBi���@j�m���=�������;�j���{����y��n*�J�'��`ԥ�Nbj��)�J��-���=[/���W\�
�,��dƢ�͡�����ޞ��[��e��T�u��1�j�^�"��@��F���:'e��)�\z)� k�ngᕀ�W�L
a�<E��a�s���^�^t0�S&d�n�9���H]�2��ƪ�T�݂��2�]w}Uz4K�U�_F��ۙ؊��>i>T��ݭ$����V]:����P���iks��2�kulJ�Q[Mf%�����s��;P�Bf�e+��>[�M]r���Y�\?��e���)l/lZ�	�T��_�Ӹ^v$T!��MO���j�}o�T�1�Ff�޽��cԅ2k�^\�ă��l�̬�-�4��z�f�h��������<\�	�L���J�y���dz$�a5�i��vU�j�j̚��M��SlP�F���u���	eP�aT��x�G�E56c�Nq�{�|f�eVTY{K)�=?���������!PW��E��[��
���_� ��@"f�]R,X�ɦ!�fbei��&�i�I���I�D�ʜd&�dRi��I��i�I��!	I��	���bi�Y��!�U��&�i�	�!�U&��I���Tei��h`bd	��I�$Ri�Xbi�I�i�I� F&��heBV��I�B&��I��aP!��	
da$$B$)�bdBA!��	� a��$  a bi	��I
eT&��	
eB&���P��E ` e  `P aB aB�haB e dBP eP `��� `���� eP n��(@�(L�{�8�
2��e�������+�`E`aE`e``E`aEz���U����������������뮀zVV@VV VTVVAVVB�^q����
��
��
�����
�C"+ +*+ +�]+�4�
��
�ʊ��
�Ȩ���!(2"��� ��@�BD `Bi	 �f�P뮑:f &��	
`i��I
aB� eRi�BQ&&a�NpHS
22L
CM2�!L�CL�*�L�CC(�CL�@�'�^���z�����Q�QTI���|���~�����������U�����?L>�/���(�`�����ϯ�����
��~����������"��E b����BO��������������~�o����@��������ϡ��?������_� ��0! �B@�"0�(B���@��� J���*� HHJ�����B2� �+(�(B2�	JH���JJ�2�*@J 2�!2�#ĨR�(C
�@H%(J��B�B�B�0!J �2�P�R��J(!@��B4�"!H�)J��%y��� +��� *Ĩ*�!@( ((�CJ��
H$��BB�2�
��$(H�$"L�B,(L�@��!��E���?Z���
 �P���������?o�=�~g���* *�?o�?g_��3�����i����������a�PW�~H2}�?�1�D�@@~����C�!�X~(��/? ��^�@}������_�=��y������?��?G�0E o������ *�A�P�?�>}����~�����`� ~'��@���x* *��������E P�a��'�z?����'��������x~���x�T�	<�}���
�ӁP����?p`n��?���~���AU!����*�/�����_O��0��>�b��L��kw���ǳ � ���fO� �#�         ��                �         o� �R�@ )AI
�@@ *��EH J� ��TH*�  (U@E("���T�JH
U�� ���)��U)EJ�D�����AR�
�Q
AR��T�J
�U**J�IBR�Q*�R�G� 6�E"�@H
$� >��5�tt{��b�&T�w��VƝ�EC�������{D�<�B��v��{�BS�W=�)k+�ݴ� R|=  � �s�� ��+{�O��	/�ω�t)��������:}4�[f�j��}�T(���]���/y�W�Ԯ��^��wJ��܍(�
P �$_  (�R@�DB��R��jV���+��IF���5]�z�M�*U�U^�z���n��]�:�´w�׍-�\�Uw�ml���Q^��ХIU)B�� ·ͤ$�Ͻ��RnUQ�V�M�w��keyv<�v�Z���{l��{�H��=�����6���{��-�;�mAm��B�
 �>   <�JPUA!(IJ�%9�M(�-PQɒ���ХuTV�]��*�mB��$VM	N�J�����-a�J   p|�G݀n(��(ws��� �'5Q����*��Y��rE@UI@=�  �R��
�J� H�C�}ʠ70�A�Б�AQ�D�pv�G b6 �f ��JXts��   U�   <�l �
���ʀ���	� nQAp gb@01�!����IR�  ��!JI$R��ERHE���@����q
. ��@��Y`	@#�EH� �� ���  E/�  �y�A� a�UT� �2 [�@q h7XҮuUP���r [�����@��$�P��T�24JT�@ z5T���(� �d�&%5Q��i���*E?�@�  �$�I�)H��� 3��������5�	$�0'���L册�w\~2��4!���HH�r���I	MI!!��$��$$I?ؐ�!$`$�����O�����{��z��}Z2�U%#YZ�ZtaZ4ٶ�5�ن�RyYB]�`�-���)<ږ%L�CE���˫�[����͕rIB*81Zتachɯ5bCc�[UjR��UM #{�m[�wH#��nݨ*f�,��i�>FYT-���t.�m�%���z�G�I�n;�Xm�I���B�[�U�E<u�&�V�oF֋i-�q^�<d�.�ɲ0��f��TOwt%�:�-Xj6��&m�N����F�IҳeX�g+k�[*\U*�¯p�e��f�lZ�{X��.^E�F�L��;���Z0ɧ	z:�w���)'-DhV7j�Kw����%l������(����ma�F�͂A�ì�v`���Jy�JS�wwy��Ê�I� 9%h�/$:�-P.��$*i<0j�p[kn��r�[Պ,È��Qnk��#L	���qV	0�0���S�f�X1Z3t����l�O������%��k�o�n��f�4b��w[h��Y*Z��(f�m���
w1� �)֕�ҝ�Y�LU
�rj
����:����u�ʶ��9��wdb�8���V�r��q-;UJZSM��G%��n�gp�,:�o%��zV��9����s4�PMV1G6ʓN���wb���C&�l+%2��Ԛ�(4�J͹�Ηk,�2Qk�s2͗�Z贵�-��Ԣ��:eG�h;c6�����ŏ��ePP��%���%�A�nN�.��(V^f����G�D���۷
z��HV��e`�;U[P�F��~�(Dje��aH�jL,eQ8i�ˋV�ia��%�{�
��4֊A\��0�*��d�$�3c�{gY�L-G��.�uE�;q���̣j�2��U���x��1;��m(��zZԷM&��:fZ�zh�ϯT;hZ�r}���6�n��s>I�ѹJ�D��T�ݛ�wj��͍EPR�I�e�۔I�A��"���ܢ�&�!L`u�H&u`4U�Ƕ�p�,M��qFj�-&�MM������ܚ+�{[�R�]L�;�"�ݭ�ih�̽Ԋߴl��"�r�J	��pT��%�N�ee��t(e�.���B�P;����EZc6�D���I�����J�������ٻ�6FZ$#AJ@ޢkU^�ef��ih�x��l�ÿ�"�3m����؄[�Sϙ�V���SY��ƌ#y����9(cq��Z�[�|������I�t��?�VLyYuP�\;��h��Q�u�P�]��@^���Qd�%��UMᷙy��a��E��mY����ִr�7]G��aVwuJ���7�8f�v�tQ�L�n-˙��H�$�����7ef%1mAn�T��VUn<���]�_ٳ����˫��]�&@��Gq�A�;T��U7�j��5A���P��;h�:�sj��)����x)Zv�-�n�Mj���1Ts3n��-ۺĕk�3k^],%�cŕCl<�e(ö�L�Y�v`zwK�^�����P�ܥ�U�w]�m�e.*h�f��U�_je<��]$د�CWɴ�ǔUip�B�W�wfX�#6�+wkh����^�T�6���#Z��aY�K\ZQ��)�~�v-hs+b2��n�&����J�=f�]j��"��v,�nR.n���f�G"����i��Ҥo@�oQ��I�q3��&�j�*�UX�.�㺭��t,	*x���NV���Ň�LGF]7M�Fݨ2�]Ę2�����g�fnU'�ef'Cj��6�!^Cd�A�*�5�/n�{�TOѬ�i�7[K�!�`�JtI�f�fV�ƫh�P��J���VӴ������⛱Ҭ9�kø��X�����P��41		d$VX˚�E�ʴN�p^�EU~l]^��sp�R@��찦#Z�ܤ�ʀ��7r�Ǖ����wU��8�,�k��P�-U�P�B��2����on#��y��0�c���zn�<�a��G�2���YD�V�ZmZ��
MN]�@(�vE��z*�.J�jVA-;�v;�چ�2��L�J;�&]��e���o2��̬��U�f��EFr�[��^(���V(\��(�M#2��Rc���d�M݉y� ���C�$ѷ�^��*�5���i�U��F�0mc�M����&�(���c3⫼��DJn�QrP���w+�x������F�����s2J�MEG7+U�f�2Һ)ͪ�n�!F�V��zݘ�����cV��Z�
<���7�t!ݫ�����&��%LͬUD㎡�H��v����ԲI���5�d海�ҽTfF�I��5���y��i���owW��PW�,���!�ܑ�ۅ��y�Br��ú�^Rcu��UtZ�u4P�kݺ�+,]Rx���6�[m���݄mS6փL��oMm<�"5�x�Ù���)Z����w3-ۅ�巋1�M^`7��,@୤&���/�n�l�����]Ӧj���C�f�f^m��\�u���ߴ6a�)�fdu� �KF!��e����V6
r�F��{K%Lf��J'-V�شd�D�a����F�ƛ�n���y`�.��2�fI��A3��n�:)��P��K4Pٹq��R�3bՖ�.�y��W��M�^ғS��Qֲ22���Օ�cJ�?�^eK��^��r����,%Ŵ��АʹZ�kj��c"�T���u�a���2a��12������33.�VV6�z+%������Q�R��nm�V�{�����#.�i���Sh����*���XΧ6����`���r��2R�bk�H5tk�e0�h���'Y+6mZ��j�cl���v�Ϧl��t뽠���W��trZ1v�Sn�T߭e�j����Xk~w��nE�3�6Xґ�U#KQ�Mw(\����˫92^����0^����m�f�w)���Y�B�Z����nu�!�&���Ԣx�n�v��x�e*�&,jk�;&[ǱP�S�y6�9(�Y&�,��Ù�չ6�՘�m�z�i}X4��&L@��vN޲��-7F�l̸��Ť�8N�d����:�£{�(���h�B�k��l�[��Ǳ�5��ڛ7t�Y&�̢��6���;e]�y^�uy]�,(a� �jI%ZĦM+�yuxeR��d�16~��l��14aka���R�b�i��J���rË.^�ֽɭ�`�u�h��D̔�iIi�	.���cڼw4*�c#�6*�b9�5I��pU,y�2܅ͺn��w�S1�FX�9��
�"	�-�n�V�˙�m���6TJ�bJ46�5V�̳����m�yT6�Uc�TF�D]�Zj"�����wU(+� ��u3H{ZŇ���*�/n&���u��Y��I��ò�4UUUP��2na�H��$��X���w� �@rޣ2�_;:��st�����������[���K.˺����m��(ԍ���c_�4�U�0�ndD�6��5W2��i��u�A����(ʩq�t�UZv�Hd�Ȱ��FPf�؟:�"%d��tv�C�ҡ�j�zn��3&�R��F���@m]+�ԑI�z1�ɘv�m.�度ֽ�&��^[m�^V��lYU�6b¥J�j[�(mLܦi ��u�^��\�E��g_ҙ�tkR�Mm=�xv��V!u#�f�ˬ���UH�N�(SXv��=�ٮE�ݶ�S?#l�54��c7`9U2�z۵s5�i�(�ۊ��fyc@�P��#Gպ6S�0\"�"j�"df\���V-Ɇ�D�ͮsF��u�ʪ�]���k($�,Ç�EͤU�5����ڬt�c6�oc-Lҁ�Q�I�9��;��&���0�FgvԵt�]�A�`w�] m����+��6�#V�RŤ�u,��v���v�*Si�T��:ʺ*���b�r�dW��,')�6%.ISov\�7-��2��:%�5�X&*�*i݃�q�)ƪY7V�,ešUC(�U���T)�j��]��Ӌ(8�Q����F���
�{�����6hE��y��̕or�\u6�=4ڪ����RbY�N����%VH�[aZ3ed�n�kS5s()mQ�*ӭm��ֶ���/U�]���1-���y��)�E���k�˸l�ML��p�;�����ZL�S�ke��d6u�a�&�$E�B��^�"�Q6=�e:O`��X7R��e*���B��ݛ�0�f������6��om�����c�Z��y��'���P5{Dl�H�������a�ˍ�
�t鰪\ã>�j�i�-�xtɹt�@�ƶ��
2���Uf�lR�'-uB޴��Xu�/��x
8�{��f�B�cVb�nf�w�\��4`��a@�d�:��n�B��`���ȂUᕵ6ؚAʙ���xJ���T�G%�{���$�K���h,yj���Ӻk ��M���ń%V�B[Yz���r��V����I��+*Qt`{Gi�P�wuy��F�cn����8����R����e�r�-b���Y.�C���d�,գ�vL(�w�dG�ة��)�&�,Z3B��}nmʡd�F��VK�\1���)cʫi��	8fa�kfn'���u(�^2�fn���&�S�V�ZӐ3�e`6�P(K������J�W��d,
�nf���l��Kx�z��eq�J�T�;Tc7�ܫ�l��2��6����",Vj�KC.�*��40�j��dV�2�����f�c�+T�ܶ�\�+q�-�Z��]A��a����vԺ�`B��M襹kkj©�d��ڇ��1�|�=|eUY��fݥ����1�ŗ��Y)�ZVA�G�Jej{+*��6�,U���u��ew�˵�l��4��B�J�6E�F�2�[�eR�w�����V�I�D�wXہ7�,�%�݄B�f����n�x��iԓ*����2�n��R,gLuUm��l^
�2f�O�n1��f���.]�˄n��d�x�IMm��TE��&ө[Y-�5u�re�:6�V+��І�K�9�}_Y*�#���^S2۫lJ�eU�V�;H�L��M�2��D�7.�J���F�<W�ڪ&h5������baҲ�2�J��mi���(�f3�-�Ne]`yN�edzڃd�.X��cQ�bt٬[b�nlܓF���M^d�.k(T�KY[Y-e�dlH&��2a(���B	��D��b�#���(#T�Ӎ�ʑWQ�"�Lܴ���q�_K��+ �y��D����̦��}��ͤ����\mlw�+����P^2�eeb֙��m*XU����Ԯ*s��T��v���U�Q׆�B����~�ב�Ŋ�[(�-��B�M|~Z�3*��M�nD0��6ғ1�Ň�Y81IH��P$�PJ�osu�����5{Wax/Sl�g*�V�OL�H��1f1��7�?�������z�7���h�+"P��^^ݺ�D�������(�!C)�lm���m<��C�z1��jͰf\Q�� onc�BՔQ�d�j�ѹ�Y$���ne�c�&�5V�т�+�\�rn�v���ct[�����bh�f���v���X��-廫�����WD`���$�h�l�aۢ`.f������^�)+Y�V��v�)^��t��Sne�̷��:p/����ݏm�V�6�<9��TU9����kK�'�uB�ǧ5���Q�H��iN3[�u�O%��c���uF;۵f�3vĺR��
�N������q�]�ML�T��y�y��KV�^܎��95�2�KU੸�+\�̖��6�>�*�u��wM�CGP"�T2��M�SvV����E��[)PG0���F^���u�Ǵ�(l�[0j 0�xs���n��EIB;w��*҅-Սd�f+,[�~T7p�3����w�����4Y��B�i�fK��gp�۹�ef�!�s��Y�;�^�U�m���^a[���ܽ�$͸i^��J��6�*n�'QA��r�u���lZ�ʒ[�IFm�'l�Wv�'J��2�����T 7U6Y�U^�[{T���(�wY�}--�Cp��V��ө��u�(̗�NXa��d��iy�f�L�ݕoY��"����"�KSf9�ܒkwWX����c���u.�D�,��|� ���@���GGoD�Ch����%��c3t�oC�)�uî�L���V�-����Բ��i�W֫U�R0B9Y`���B�[ĥe=�C~XVͱ��ER�y�o�FՋ�U��!�c!2��Z�@̦n����n��7��^<�UT�8r���Ϥ1Ŷf<�{��ș7�dY�ab��V���{>ʷ�'y2���%r�#B�jf(���̊�)�jAA��)W��N0�k[�4Y��/i�G�kj�)�yX��2j�
�dC!�vNd�,*��n�pfE
!��w�][R��5�;�uD��I�f��;U�f�x�薪���mV�����Q�aܧU!�j^��'PuYN��yj�������R���ͩ{0�F��Ph�G6*�tf�"m�.�yVt���2']�Y��	*����)T�<��Ně7f]kC4K*d��۶�n|��y�
���n]bH]�n��YT���\w�`�C�&UQ�p`Z�)��#V���CכQԒ��[�^MUpTS3i���l�,\:fTĝ�-�jmЇ^IM�-#m�O6ȫ���U�
��dm(SO�����,��j�kRHÕtܪ��YpenV��{z~��j*J��RM�Vm[w�XmU�lQ�V��Wb��|wR����x�ٙr����S��1S��a�Hd�VM�u6�B��U�1���
ڋ*Ҽ��j�J��sm哻x4"`(�h��yA�(��k0�M
C�[iأ��+*�]n��4�����n�˔�,��
3C(��M�wU4��t���\�%JCC.���w�5wS��܊CZ�`�y�X�!޷W�.�[�]ѭ�pl�� ��GL�
�#5;�k\�s4�{nD䧥B�*���C���YVϊ��n�gh�������BV�Z��h�mѫQ��6�[lm�5j6����mlm��mZ��[حh�E��j��Q[�X��k�F�V-��U[E[cj��Qj(�lmV6���E��F����[[j5X�U�ƶ�j�Z+V*ثm�U�j6�h�Z+m�U�k��j6�Q��-���Ŷ6�ڪ�QU�V�m�ڍjŬlV�*�QV�m�E[bձkFֱTU�[V5��U��kF�QZ�ըխ�U��X֪-Q������m������Z��Z*5h���j6Ѷ�m�D��'� $���B$������,�W���qf�f]	P��w��`���%� ;��N8���ӆܔ�V(�bpe�R^T���7]���[1�Hf��e��m9ƣ��(塘�n<��s"�(ؖ��5y]�s&4�.�5+u�����Kʸu�����T�D�c]^���d�c{Z����5�Sko86��i�
���Lf����6�0B���	�ҡ#�V^�oI��Wq�B�]J��%wUw��)�.V�f2�1f҆Le�!Z���X""f�{��r�L)�-��=`��o��y��WwZ]ίRɲ���؆B�d5#el!�s)N�b/Q$�ƜN�rh�Vqҫ��fC�6��.�������;@�r�$Ҧ{�]��'@��cr���&=7}K�u���Q��+��֝ԍ��S8ᶔ�;j�Z�_F���^Aګ��47%5����h!}M>�
�\D�_M��.��拤�=հ<ט"��[v��۝�{w���ĊYq!���1g��_N��!�i,T/�2�oma}\�F����wH��F�m�8����S�׽�Nb�Z����!w?�I����X�B���F�U�(��Y�Z���iVl������*�T9��v�ʎ��]�]׵rW+Y��e.��WW]��T��{�Z5�i��J�Vb���؍�̧#���j�m�`��V�ȢʬW���X��쌨Krr�m}�<Ѩhvs}7�[�BC:][n�ޚ���X��'ئ�W}�s�՜�_o+V�d�7i�MģJ-�-�UnMޖ������s���/r�g7�g�nn�K���#FIs�H֝7����j�a��弻]9=';78�ͱ{[S4�l.yR�b�tp*���};75�Ǆ-65����Լ��F�mȰ���#T��P�H�@�r%�����a�쬗SN�vc]2�v��^p�ǲ�a����5���'�/P�5�Q���땝�����ŕj&S�O���	�f�˝-Q�"c����Be�$���{iU+N��F��U�^��3��V��n���jg>�f%��Yuu�Ⱥ�K^���S��zn��݌�ܔ����ܛ�B/�%��ۼYw��y�3�rm�,�tT$qM7a����L�&�X.���c�K��V��0�)c9_c��!J{F]�w�p拗C�`ܩx�&-�d��w	`�P�d�-eʢV��p�};
c3d0���l���K&��Hi�͕>�ȈWS��Z+��JQ1{��M�ŸiN2��ׁ	�8�nP��72��[&:}4iڣM�Vۃ��Y�Rw�]J`�3��̳& kv�����[�=���/��d����E��]]����0���j�p;���e�j�]*ɢ+�m3Gz�f`��ݙ$�E%�o�<��(=��X��c�+�.���'pW-Y)5�3�����K��p��o3����Ob�GW�~��Ԛ�)���v�C"aVM|lnV1%���v��+}�:.��L�i6�<�V&�?��OWD鴳gV��U������,���~��mq��ؒ���ذ<ج���,�鮱���J�*���E�����|��N��lX)�j���d��'XN��*U��-ç.�S8�zqb��ۼ\�4�]�[KY����-��_`9�D�Z���jS;kq&�%1ۓ��]p��߷�y>Y�9�UL�hq�,���s�m����
Ui͉i�Y�jXLM�/O>�mr%<����/b�QLMIL��fRC�@�QKM����U3CIl�G�V�öe�u�!䐣V�mP�B�vU����-�ۊ�t[��m����WJvX�\�4}6e}r�%:A���ce���bs�V�]�ĒUL5R��k0�.��h�Ƒ�\&�qç-�Iw5����M�V�e�Ksi��&t-�/���w��̻F����L=FvM��A�J�p���f�Y��R��kQ]�N�`�\�v�B�se����4�t�e�����4�P[7rNWU��0��)�%¬⡯�o:��w�)nS�. �7�J�*��D9�`�k{kK���BU:�)��f�7K~:�+d�;ר�ř�Ylf��8pe��uV3��vV��Y�ySa��s�����c���������U�I�X�Ц΢uFٮ�mgeF���������(�؅`㥹.�'-��E��N�b��uL������y���H��N�[�c��D���t��T�qj�ʇ�YՉ_��3[��Ҥ�o6�X��evur��_-�N����R4��;Pݣv��Q�<y]r&���n���ն�`�p���+�s�t�on�\��P����yy��nu��e>���#�3��m��h��t��	(n\��r�m���(KdW
����g뒷v�1�ɣq��ysadfnVhYrK�v]�,XL���7�Z�WfT�p�z4Aŝ������;���BE����c��"�r�q�qf*kQ��
��{�8�i�g�'�̣"փ���C�v8އ��yW�><�Qnּ睈���7�N-�LG���Z��mKT�b2�V��Ј2t���%��C\��w{��,�f�Z����j�&���+Z[�ˏ���/�b{+wLCTг;h�w��
�E$����q�|����]"�S#�U������Wu[���m�86�]���ތ��4����o&�Vnn�Ǯ�f^����0�9���Kw�SI�Vu����5�:�Q�A�	&���:�CN�Qm���	���\�T�X�CŸ�E�e���3��mM������ͼ�N���kM�gp)7T*��́aW�iw5ll�K�
��wz���oF�j�u�;3���ܪ�*(*���×�o/�y����M�O�*�e�
�}��*���鋻�Pv��j霬�r���H.>�ÍΑM�J�6�Pi�yK$����Rmv�I
��P9h]�ڋ;��?lB�6�\�b���^
�b��UvӧL]��*+E��5-��
�s'F�fi��姤�[ɍ���ח������븵NEZ���+���67�����FJ�O;w{���dR]��KlSI��'�2oG�������jBe��.����A;��	}-����ފұf�e�z�^�;LMlmU�5�Q�ɫ��|�󲲗V�Tn���>�ڝ�v^-.ę��(�ם���.���U[ŋ"�Fw{>�ӯ`�Qg�r�KyddE�rM����u�����4XW�'M��{��a�K�wu��C���X�[!<�7�-��O�D��]���	]�4ٽǘ4��:�k�(�n-"���nn�]u��]�J���2�X��r�=�iU3@�[�M>�s��]�S���~�W0�Lޫ�Cn���G3n	�}�d��zP�y-���zYڕ{��X���B��tl�)R�+����T�M5"���E�r-l�1�#I0��7rNb��������	�`z��Rf)� ��(�X��Vo^r��s�e����0L�7���,�7x�n�Y۫�r�Y�V�֤�Ġq�5���&���Σy��]a��m^�e�K�u';*�Th,�'c̼췢��\MZ�~y�rm���́����m�;xPް��or� �{���鷦�.7TK�s! �k,��v�`�nL$�h,��'9��u���MV���b�QץQ;x��7Z�yg%IE��h��w����F�Q��+�H������z�|lSʄ�c<np����n�6E:��!
WL�q!�.L��_�8]��a��ٛ�4�u��t�H˰��p=�#�l�0J<e��%��w��<NL��f
�3�J�4A�gV�b9`����|ۭ}}٫��-=��v!9�*��*��;���]�4brQ����ゃe�(�h��^خ�*�U&o��y�D���3QwV�<�0[D��&��f�/m^2e�Gn��Xd�����Zt&��<a���Q����U��SyB�Tlė�+�v��h���N�F^K�|Bf�e�VX���{�fމ���z�i��jc�Rx�]�mV�e��n���Sڥt�L���x��N.�uRZ�\b�9��y7�����Sw/(n+�5ߐ�vJS����O�Z���t
0�̓Q��S�R�h6��=���ܫخ�Z}��|� 8����fR9��mcպ�2v˲49b8��k�˾�lފq����j=�/6��`����o�kI{� jVb}u�P����9���󠂏ep�m��yG�{��ya��|	uQ�|ŉSv�V��F<B�4��,�ʄ��ϧJ��R���B�x�	�9e�#���2��b�v5b>v�Mí�'P�ѕQ����c�x��q��:VRh[u$���3j�ݗHj�,��R�Be�b�t�6}s,h���j�����T/�Q�Rn�"��c*��h̋����42�s�h­��HYr�a�7v��&�ท�ͳs���e�a٪�L�6�+Ӄ�uV�z��&��!�V�a.�Jqr�{dm����+|z���9ٴ���)�B���:�����V�EQZ�(l�U���駜􍾼��Fe������қ��V~�Þ&�ed��n�/�e+�4s���ף�s�ϯ�L�Ec�o0^ҬߩV:�b����Ι\�Um��i��(j�h��_;S�Ct��Ê1s��k��ᬒ��Or�&����u�5�X�&;�]E;�V���%�v�&�q���/a%W�}B�.��kw��Ҝ*�#���
�הĻ�VZ`J�˅��Eƍ���:��e���G/Z�͙��9>X�W@ڏ�n��f9�1ŉ�Ԯ.(h&�)=gm����U�!ݔ��Rqӂ��'[�sH�լ�����}���u��=�VX�$�]ٛ��,v(�dV(��k�������+9�b�E
Ί�[�vk���!���G�&KX�ufkE��3iR�02�w%��J�bo7&�.���̰��;��St�`�X�P�X��r�6��z!��prwZ	��5A�7m��;K6��o�5s�vl����/��!����EO����cg.�i��.6�jʗB���q�S�ĝq�S�)ws4�֧JT��жm²ڽ�r��ܫ��a%Ƹw�ck;�A׍6��Ys�[봕�wux5���]u=��M�w�۷��-q��.㼖;��B����V��DV��(G�,�����`x{�u-&��np��E�.X��e}r[�]Jsȯf�|gk��W�%eJP�}�t��쪼Ĝ�\�_X��[�{E��[|gPxl�sr��F���{F6f-��e1�Z�n3c-��
����ד0�)Uq�v��,�g0t���d5�ދ{��?�d�\�Km��8��iZ5k�;�b�E7JҨ)n`�D5�1�qe��m�wU�jƂ�_.��ͭ�뚩�^в��b�!U��y��
4�Z����ޚ��Pr&�c&�v&X���Z&#���V�j"�b���X;sn�Ě{��h):v]<9�)�XL;Q�IE�uit�_��#s��qY1���g[��u)|Yn�wN�G6�;v��M��*�8&���(C�*ԣ0v��.J��+��5��ތ�&F�3E�>����!�OR���nZŔ9ŉm�N�/���z�7Yx�ժl����^T��Ov�n��\�L�o���:���
�
��D�;At�2��Ӎ��;**��[�;�0����ん�ʛ��=���R5W�g~�b�>��<u��,���Q{w˴s�WhA
l�������2�}�Nuƌ�'ec�5��(��f�����Ֆb��m1�C;*�Yٯ!�E�Dޞ�I��XQ�=Pr�:�x/�{\�P���(a�J#�ln$;m�ˮ�PD;a�x�t���r��aY��sHƖ�Ť�����,�d�����Gaˌ�n�wZ�ޑsr��g�T�K{�7nB��]C�`����gs�Gv�l钙�r�(^J��Np7�k��F�-*=��쫜�r��^Lt���� ��H-����a`b�����D8hf��2��9���s���Z�\�w�����2j��e<�OA�K:�\���-�����F����y�fsamMk����J����}EU|p�s5}.cn�N�� ���,mE��]��{�X]f�!��)�Je����	*��3�ؓA�@���QL�N��ځ��#$�v�Ԃ�^�R�4�R���ܥt!8wc���x�MN(��XT���E��ʐ�f95IӭR����ɮ��ј�桄Ny�{�f'Z���WMI��m\�m㪳�ϱT٪�A\_u�f��'j�Cg���.���M������xMȴ�.>{���7]B�9xJxɡz.�چ�f�չ~4�E�z�1ڇ�7�6��&s��L�L%�2m㜫��.�E����o�f��S��%8vd����ړ�5FB�N����l��7�'ru7qP"q�bL�۽�|���ɁIR7�:���-hlg$�~t�lͪ&tFgG��D���ج]I30ԫ�qvy,^�N�e�u���[���_�8V[w>���UU6����z�x�M�r�Ik�
���I��Qi=�V`�M	���K�V�]��i�$����Y�ʜJ�up^��朱U�թ��jɦ��SP��K�jfx��U�m��a;�&�)V����#��n���<DF�����0w;��-W��X9VhK���JjխW{�k-㺵�	,�c2�@��7���0�V�Z�JZ��b6壑�p������e���EK7���Xw�;�����l���f�jp�2����d.��z�N��`�B��4��0S��(1V�������t������3u�e���5�ߖT�W/*kwcU�`�t��kx��p�ݴ�<f�!��K���Ļ�W]B�7���F(im!d�Ú�&���"�IA��uz���h�W\EC�ކd��5e悰oF��{�uyws�p��;%V>��6S��sKe�Pe�[�6�"�;�w0����li��P�&]v�S��eb�1���ɓ�,ø�W:7n�\o����	J [��7INf�ݞ4R�hqGkme��5t�Rih���.Z�. 3�4ڋi�Y��:�c���e3b0uA���lF��It�͕V�eu�-IiV73���\��1a�CXJ]�;�"�U�mt%Ҹ�ز�^ѪQP΁��]��am��ҵҮ!W"�\m�h�KB��S-(�*(��ˈ:�\X\b�m��j�͗[5�ܤ%�Sb�6;mt(;�4jm�w\n��#KG��A{F�Ү�E����n��,`�tItM2��t��k."�wClD�&��%Rn��D�Ū�Q`)F��j&Rf�H�4�in�t�e.�ZX���
�ʙ�X;�3����T&n3em�Q,��v-lɩe�6��Q)hj)DUn��f��F��4���vn��kq���|=�dco؀9�]l3.uJ�l`����]�夼�n&q�il����Jح�lB#f5�<6ȼ��aJMm���e,6�`-��ĲW�S�Є�N
K6j�n��Y�NlK4%F��Ն��E����ᖼˠ&uֶ"��da+�M��Fe�[Rh�-�����5UMX��]5��/�`���R7@�d�����"b�8�kb1i-�rl�[����V�Y�urA�4*T�"ɬ6�ۜb.���]�l��L��T̶�B���t��&&��Q��,�5K�T�Yt�Z�݂ifeJlm���AQ�
�t81:b�,�d�T��D8��M�H�HUbkm����X�9�������(Y�MhJ.cn\�6fĪR;.��&�1mh� �0&�%�f+H��.�6T�bGkT�m��ĢU�5�6�*]{ma��%����-m�t�&�W$&-�uvR]�Ҙx� ��v�8��ȌcF�=L�fZɱ�:RY���vPZ��&�bM���
@��B�H�[��fm�m4�wh`uVدZ\�e��GR:�6�La������p�[g�fb]K���4!1���l:X�39ꙋWi�*��L�֭,�&stՉ�9b�(CR�.�i-�A�J6��)�k0���ZJ�Hk�*)-���Tp���ֆ�L���0iζK�Ƀ
Siq�ksq���.��Ģ$m��^�N����#�C���R��ҁj�&�����!]Թ�)-�S��9�b�P�0JvB�z�$*�\��b����4�T@��ے)�uZ��[5�mS^Ƭ1rlu�4����fF7M`7kr���k�2
�Hk7[��sj0,���˴̽���F�-섳C
�b2��z�:�hme�ۭ ��0�fݴ�,��ob-E�d����YBYlP�V�M[*ae�
�u�]�Y�5�5�,��5
������[u)-+���:U����-��f�.�P��1ƕ�)�6K�x��WYZjD�<J���K���/9�i�HՇ4��bWؐ�$��X�\YK�h�)6�4�J\�o&ZCmHfP.ۓL�B6�nc!��K��$FƮ�&,�ۗ9պ2�-�`�(�,�&�b���*�P��fי�SW�+�����5�c��)R���ص]�d�
�&�[v��Z�cm��4B���,.U�T���s��L\�a�����2�1n���8���(JA�Y��+.-�k���i5�YJ6���Gv��.�K��^ësHn�4�c��sf�Kt�fq�)��6g4�*�-��\5��c��-� ���J�b�C�:�t��f��Q]pZ�:�c���,p��RT�s�����R+.U�C01CL[����Yl�.�XFX�v��]u�j�@
f&��͵��A�mz��C,�]f*9�1ma-�(ؑ��3Al�f�M��E5�LlWBXiX��F�S�r�.�� ��í,�,�I2��kȌ�@�5&��n��Z2�@�5j�.H����Je3�S����%�.��Kfz��.����VX�&��a�e	K_I\��-���@�M`��ܣ����F1���6qC[<ǆ�<F���#��]qmMU{Mq(X���*�A��u��[�bL���TL�eh�3ֳMM�M���,&v[57*���e$�ԕ��Q���v� [+eq.,������DM����aX ��+��0�����F"hC,��h�	]���h��2�Ք4�b�4 ��k4aۭm5��]��h���n�c�!��`����i�;J8K�EˡsG���0HG7[-�\-��y�,^W��\K�E�i�r��kD��q�L���A�X���
++NK��#�i�e98�N(;bXحs�q�V.�,f,���Cf��FY��҇@l5�n���5��5- n��8<e</���6��c�D�Aխ!:�\fW13s ث�-ԡ.�^`+kR��"k�NE�0�l��ayq�c������mX̥���-�W�ld!M//����PL�9v�+̷0�RV�6[l��[ΊA�!д�j��E]D��R͖m�ҳAa�M\�ʰԅ��.��;fD�5�0Kl�U�֓1����M�J�Lޢqa�]e1G�o,�y�]u��G��A�F��HR�WJ�k�-�mxE��U�F�l�"[1WƺSl^�(�1q孳�;�P��e�ց��ɸ��璠h1����L4�D�5��Bi*�C9.���<���kk2T��Mmn�6lk2�*u�͠�j��%j�l�K.lM�]Q�3�^EFZ٦��Ҽd��(��ê��U{FZU�1ґ�Qf�*飬i��]Mtf4��$f"��˃Ֆz`ʬ[���5�Xю�n�f.x��4"�l�B�c@Қ�K
�L�U ���ct5�R����&�&����M�G7B�e�
�g1�4i���X�i�vk�V�*�.�	v���3�vq��6cD6
9�k��sS�f��W+,e���B�l32荘�ݭ T�@�jۤ��D�̂���P��
X,Ȳ��dK�SnƱZ�[�����5T��W[��p�V�b��X�R]|	��_ �i����T��s%��MqKD�X�uri�-ј��%�#�Ņk+�ZM�Y�F��P��b'e�ݹ�dM�=�[r`�$e��T�l�U�@�Yeq��mi��nf�4������W8�Օre��X�EF���������bm��h�Q`7l5��M�]����ҵc����"��h#�l4��4.�ⱃ��[�CD��Ƅ#�ʡ4ĥF�3�:m�%n�f���d�M��4`M
:eh��V�s@T��-��v��3-��d�ք��Ґ4�u�,ڦY�E�6#͙e٬�֖)V�`�0א�(ƶ�6ԗE��	i�Y���el�[p��b
Eڴku�n��gB�W�)%�K06l��+f(�$��C���T՘�ʓ-��E�8q�m�,i1j��Ō�cJc��XX[��:�hO�(z=�ۨm
IX�ڲm�.���Ԅƛ�ySa,s]�R14̲�I�S��#6q.P��+���t%In�M��KMH�[��8�n&�6!��kv�t)M(�]��gWjw�֩J+|h+��.�7n�� ��S�o16P�A�r�ueX\��n�nE[L�W)^,�j#���6���t�53PhW5ņT�ij۱V,�y͎�(��ŅE�ZZFƈZ����S)f���7�[M�[[p�eҪR�akn&�"�$�Rm���H��)e���n��.�:��u��V��Һ��V���aH/�D�h��3��iKjL���5�l-��֑� w��]n�b�j�\6"�kJ[xݡU�rEGL:YM�8���1m��n؆��Z�&��y�6����d,���D�)-�\R�o�m=GGUk5�E�ՈM��4a�5�GU.�mu�`���j�aa���P�lq�a�L$0�˳v"�gYse��ZT�!+�J)2D��l�\�WV��6����`Z��ʷZ�mn�H�T�����7�6ؗ��:��;h�vĭ2-�--vŨmK��d�X1%�]
���m
�����1�u�X�,1ˮm\�V�UD#��n��쮦-2�+
�`T9����#	`H��!��1-nSK�]h̫6�A-T7�S5õsh�5N%��+q�/B�=��q+����- Q�6���w[ ��q�m�	X F����u��޲����- ��Q��D�Z9.��6C0�K+
�c	]�Hp53A�����1J�m��0���e\���8e��C����W/a�tU��&�fV�K���(��L.�Wͼ�'��W)-�����)�
�pQ%���A�i�m�K�������L`���]1.�6:0�l�쩛�sƙûni�a�L�[��,�&���)�c]�^Z���6�u�+Z��U�E�ّYt˩ZCd�˭�T����V�f�41��Q��R!nJ,�Z���M��0ڔ6cZd�ˢ.m.�GcC��I��Q5�B��.`��ˠiW��Xj���f� M�)��]��3#vZ���X��(�J$���rF�/���&�N�4v�����������ci
��;bU�u��փ�1kR���6q��fEe�9��7�u�����]K��Ǚ�2gXM4�Q�V[�P�$�����;f��B՛�& �0��gB9�R�iw-�1vE+ct�U\�`tkFxy�K|<e��;Q�i���,k ��l�d[j�K`�^�����sK�c6�V���$؁���g�z=J���j)�ִ̻`D��5�U���j=��6jͨ���-��\�Z``�Q�[ɳ4�b�a��J	y���s�#���PH�m���D�X]�.��skYtm4fZ�E�7!�Q� �j��Ln��7u��f$�����fhRԎ�]k3�3-͏euYHF���+�Y��)v]Yf@�mV��sx�m-΋�Kx,�^p�J��aH>�Mf��cU��Q3�R��qWl�.�p�2�W�qb�9��]��U\��Y\���Gh˝\�Ҩ��I���:@ڂ?Z�4j�Q�R���(�60nn�Ʊ�lkMů*�$Eʸ!�HZ(Ѵ`��bMHŎrђN�ĉF��Mt��k��n����ܵȃ%wrE�[�����ԖJ#5&��gv�VKF��QA�^mȣY�ۘ{����sh�w\�d�ss���\�m�t�9�]�wu�\,guk��lRU�-�H�c{��Q�
R��t�Cמ�b���"�L�:�:6�,X�e��Mp�kadɉ���f ���,�&"���*K��WfW�q�,��T��fs�)�i�"ر�f�m�t���T��UT�0�v 	��=�^b�����hf1�4c�n�.&m��Z�5eu˄��\�	^v�6j41Ha�-	�j�9�L�s,��V)h�
bm��-v.�lf`l�f{0ւ`Li�͢�q]�-!V�Rm��L[Z��jV6��&����9�(� �GL1�����[m��Q�vb��P�%�a����Ar�u���\8I�ءu`;a��e�Qئb0ZJ��.*lJj�^����,�Vk5�V�j41�(�U�U�1ete��[�Wf�0[���Tlm	MP�A�\�dM7�mf��k�+Ѷ5�D��ChM2�KZۣ-�Q�,a��[G�-l�0un�ڵl�Գ��i��M�X�Œ������[6!������i�Y�JG2����f��Fܠ�r����iE�8!���[qՖ��f��ի����Wrl���a�EsHJ�-t5�,�.�K���e�]F��fbbk�I�PZc��ZzX��ݥ�b��Mk��b�,�C%kr�j�PZZ��˖Ksa�C9&0��q
��{[[]��b;�3&lb�]TZ9�1���e����샜����a��u4�72�@�Z	��J��`�lk+sG���*�5Y���bMe�A�2����C)���jѻ-t*%�Xqj�7j�VЖ�+�%�,i��u3��nan��J6�ׁK��<�t4�;F�9�e�3"�E�W4`��jJ�K)J]�Ve`�&�]��[-cɆ��nlv���<�f�I�Mm���If��2�
�G;e��ǳ�A:�p�l5e�9��m����&�� �Yh%��IZY�c���h�t�������Q���,�`�FSD�.�Yn���I��l��:����Ri�w�l0����2��J��R/Z�P����K`�"���W���!���yiPo��HB��R�������6X*T`5J�Z�FTIx���ͼZ$/����[,�A���H0�e��U�a��m�XUW�YX��Th���0@��)
%�!�����v0�T3e��(k��t8q��d,̺���Q��t:G�D;����6Y��c?�� ��*����6�c�w�������b'{e���*s��@�b#Ǎ�[�8�ؚ�ݑ�:$�x��N�]�o�6��S#���@��
Jz�^�=�� 2�:E��?%������5Qk���f��FSv\��%�2Az�� Q�IP���]�I-�U�3�4�$�s@����0��:x�ŻzƗ��� ~)�M";�����wP�R����Ғ�E((nD�ȴ,ذa⾿xzk�n��$w�$;�W�!?$�%"$gvY׊dpPu4��DZbe�]^�єn�)���se۷\�-����-�ep�~3ژ �A4��n�������͵����m{�,�zҹ���鷑�4h��#<g9͚�������6#D"��c�ߕJTb0�H+�r�M�2ޱ;7���VϽ��l�)����X3*�5���"�=���Z���6�Z[��x?u\�2p�����"!���8r����La��_	�+���d�A��,{���W9��h{c�n���>!����o( A���Ș"�ZcDN:�e>ޱ��)�\�h<w�~2F^�l��^m��쫹��~�#�,�*Z�/%¾�{X8�?~<D$����% ���3�{=�M��=Nx�ޓ���%����?9 �"��1hP"�����VD0��ۤ�I�n3MKH�
���.[�,i�l6f��U��3�  ��A�7_�V�"��\����$O�HwOL��3=yj{��ێ�DMԠ}�^�L�.&4�̽Y
uŻ��
��:�`����Q��$�_9�*�m{�:E~���*���,�����+�˰�"�!O7��Ҿ�d���(�Uxk��T�(i�t<X�����E���Z�r5i�^N��,���D��_�.�����-��ÕA�l�Z��^l��9`7�&#�$�g�;�'|~s �A!��F�v>��܆D�.f�QA��+�H ��sb����+�vi�RޠNd	#
��P���?��&A��A�d���D%�����:���~a��^�8��~s�U�����A��0d�&,��pSޑk�$��E���aW�]��S^b���Z46�h˒;2�����ߟ�����"U�c{�z]z�\�83�B��Q����d@i`��F݉���r9�ԩW7M�YA &ŽwS�]��S�7������6E�*</�)s0�t�D3G鼙P@�0ۻ"�U�wLq�ǡ���w�ʗ���t�sh@��0d���@�"z\}[_m��F_���ؾr �Xp�&zϫΓ�?x127|:����ڑ�죶�d���uж1*�C�N�]�����8[\������W9y�0����M���R��xFdF�SmN*�`��o=ʻ\$�����>�A�+�a�I%,���t<0��\8�(	�/9�K��b�!��@�w H�� d��~!�y�oʮ�Omi�,&��0Jc��L���6��QKV��,�J!�SO����Ƌ�wf����"w,�&!��}*��ǖ�Tu�S��m���\VH����A��%`?B��`�("!�5�^��n�{�٩��/��=l�}ޓ=�ؕΓ�>����"�y�����>Y�>�|�0� ��VA�M[�Wk6υ �2╞�܊p�C���v�T} � �@�h��fz�q��T���� 5"H��ݑ�\v�e9��u��x�1|V��F�ݟ=�K�R�ff� �PD+�H���c��rǀ�A}�����������( D4�D%c�T���f4���{sQ�U8��T)T%�;'V����s47n!�fd��Ȗ�W�g-'�P����r<.m��lAo��-�Ae&�a&[J�N�u��;���u�]bLava���RB�De![6��D�%v"ɱ
ĬŨ�-�0YahխF��na����`ZV�՗�[�MJ�ir�sH�֡��\�.kt�dV]B���,�5�E��pH�:�Yr���-����Z-h\�4{X�&�����pM��v���GRip%��K5x�`i���`��v�����>mc`�M̹����^ػ[�c��	�i-�-�x�YBG����@���2Ra������=~�O�i�A�h{N5z�˥C?u}@���2 !d$O�1�ٵ=/y@0�_s]>g�r�x�S��w�������Xf�p˾�*����{�"Ҁ�+��()1�����������t��	sٴ0�@�!fJ�Rrv�'�Q��B�N$��6/���7&��!���H�Vn�1�fN��^75w����c�Ds2�#�F�͌�n���T*2�u�\�枩K�{��^q(G��eM���k۴�x��{����l�++�]��Jvڮ)+r��+ikF��3α�����f!��<���y]a�=�G��x�:_|��]����~�ׯ�I��i�(��ʖ8����Yl���¹0k.�23�,��bp�V^�T_�v���#��8�Q���s*f��Ӣ-'-�18)��ndԨU�(]]-��Q	�X��p�������`������rD�ʹ�v�����6�󷨎e�&4ffh�����um$��=T���p �">�a�(C��#Z^^�2���T8���ܙH�~6��ޗ��x�:_@�k���c5�A�p0D4�N�����$�3%ub�{��iω��OϬ�_��\(oD<d��u}_�2�K�������h�6�B�\��;vi��[!b䥚�hqH�"�P��)kH�/�?���`H#L|~#wh\��]{��SJ�x��ey6W2�M�eY\|�����4;ʖ"��6	��#ٙ�Q���VR}������&ٺ�ۙQÎ �س������("!˷W��������a�nR����A�0������i����j�{�ơ�+��ڙL�
=�y�6�~3T^nDgtg˘r��{�y��^��]:�Z9j��v��,�K�_	�նw/��\(nr2PD��$L�" Eb?{ϧR!�Q-ڀ���I"��gO>ƻ%�J���lp �">#e��R+�X9����H��Q"�A|"W�d�/���[������7KY���a~sGK�dv�� ���$c�s2��<:�}�]��'�L�4ˬ-�� g
ˈ�ɖ��bgW��(�M� b.��z��@ ����I�G�аո�//�����?�:.�nP�쀾 �P{�Ȓ�CDd��^z4��]�ȳ�1m
�\�����c�IJz]-���W���a�)v��a�e�?"7�=�}�%}FH�"J��~�z�3<����E�~��}|0���LGD�CG�")a��-�U�~��#�Gk�G:$��.BĴ�K��������J��9���g7����	}t�GY���I�Z���8$n������r�z��cI����UV
|������$�6+�v��FE3�t����o@DC@�d��� D=�V�f�cϲ۠��ݺ�,�q��v�}�H�ێ�)�ϯ����3&Ǚa,tR��&�X�3;K�6%x�Vm��M��Zl�k�3\�6-ﲤ��=(/���"d"]t�H���)�{�&�IƣsT���>?$a�+����f�<�ۈyz{(E�.KL�����`��G�H. �.��ˡL_E��i�� �y|Ĉ D4�I�@�/���1Pۛ$uM�z�k���
��3��E$l0�
��P�C��dLdA^����_��V�φ	�����U[9��q:�o��̭�%D���Y��G�8"����ɣ�U�xN�Dvw�?�����0�����|\Sהj�57~q�I���3MV��Ä�A1�XP��&�m�BU-��m�&��6��d�����<zvՔ}�?���!��f��n�Ք7V�Dp*e�L�[&M�`ګ5ٕW��00���9��:`;]�u�Mm��ub�^vd���
JٲZ!�hP���R1�rWF[`�a�R.���,��ņ�Θ�1�4l��tu8��У��H��bh̬t�2c�kx��1��؆�pM[f�9L��K�L@X�ݚ��%׌�F2�BA!3]�-v+��>O���b��֦��G#\�IM܌j\݀�YiE�~�K��g,���ϗ�Yk�묿vD��>?�v�V=����V�\jx]���hG&)3�3R� ��a��_~0���#��d�fym����?3}i�A�+��z֫�k<�a�����@C3�̼wܞ?�W�a2G����!ʪ�/]���)� յy���}�	��]_Q�&��Bͯ^O��D����G����/�{9��oZ�q��v�}�H�&GeE�;�}��#���� ̔ �H�!�)���fZ���R�:La��^���"?I�W�.mv�'���Dn�QEl�p����m����[.�1X��u�Z��!�k�����sF�̫Dq*s�+�C���p׳����a+T�.O@�@f�`��Y�$L���P��������y�'�d1N{xOkqtGo͊��!^�m�-����:���\/e<o��Q���m�>v��*���<���<~8��Vk�s�l7�y��0�B�X`)��}�¾�p�#���0�~�d��d@����ft�c���m(U�La��^�|A�"I�fe�ʝ���_�ۮ'D���C�U�i�6"��z��v�{1���}���a^Q�;L�r�h�d��AȂC�f_���W,��_@=���A.緽�!�Z�[A(� ��B��@��;�!�.y]Ψ���Uhe:��0��\�j� ghM���&,FָI��A:o��s�#��d��(`~���o�=[y<����f,5�wϩ�ՠ�ݖ�B�3F��WG���w���.���Z� �t����P�i��i�r`u�� �A|A��"��i��D���Ƒw�ޑ3,1��f�Nk=��G�+�tx�}�T�ũ�I�г�oP��s;�.�k�Ө7����t���P��2�)B(#�ˁ�a�U�̩�p
��8�;�˕B��{#��t�Ӝ��uT�.����ຨ	݋:u�}����[��ֻ���K��N[x�D��8nN.�@茻��1�GF���8��禲d�H���U�{FZ�d��=��|��Sʸ�1ꠅ�<Sz�L[X���h�-iݪ��7�GY5K��{��n�m�(JI-�#s��Pm�͸�'mЫ�$	|��r��Z��bҙ���qb�6�M�0��K8��C�i�K�xr7��Xz�e��eRn������T��DU��6�2c�;�;(�>���GE���Z3���<!��f]�;�G]WJVS0���u������"�����	�]g�L|��ʳY�C��_7X�i�2�p�� �h;X��٫I[Y��挒��G�pϫ�!h�F�u�Y���p�M`ː$;R�E)h�fʲ�%�Z��ݭ�|k3ruU�2��Gm��bj{�s`�,U��r��U���u�u�wK�r;��~T��̪:oHY��\�r)�w#�lJю�Euۥ�U��e�8kt�7��m\��4�m��Z�N��ɘ��Ne��-eU'N�iu�媦�	I�LfDdW����XB4u����^��K9��E�3CcX��l�������c&�T��!lDRq�"󶪲�6�r�5�;T��恺Yu�	�~Y֮�U�k��{G�.��E��P��A�IQ�w1�W��\�m���ěAt�Eh���j.���gu.Q�[�d:F�! ,�R�z����t�"-�+�9�J��p�V���f��p�]�75�v�\�st��wk�7.����k�p�NW<ב=�N��N�5��닺7#s[�����7*�듸������7wwur ���6u�!�F�u�e=�(�u��F�˛��/w^�"N�szv�nDT�cct���p���^�{��������F�.�*�r��A���5���6��N�y�8Fr�9�<�S�撷+���}�;��o{�Cp���d ���$|,�2Sʨ
RAaF��C�����Qi5) �S)�TҒs��AH{���w�����p��Z���). Sw��L�d���D9�4�Xjo����߽�W/��?�}���Ar�?F�RTB�f�p�'є�P7�o�ך�?V���A`|�A{U¨��h*����h�M\��μ��\�Z>wj*Ĕ�XT9�j$0�����V����Op6�RuP��S��o���>�f�o�o���
B����R
AU@R
| Ss�3�JH(P�9F��o�{�k__'���~� ,s/8��Cclf�]�ecǉ�0�Vm4�],��r�������҄��0���4���H(��I���ʨURs�$������,��4W|�8G� A���}��w�>?zK~�������.H)?Qi2!I��O*�(�s�� �s�ZAH)�͞{Ͻ�߷�� ��H){�i ���y���߽[��>�?��C�ʠ�
J��.d�e$
��H,4�^U@��������٪�zAH?T7��|�R
�Qi��YC%?��(ZJH,+���Aa�9�-&����^U@P?g���kz���ך��>�f�o�H,=�X~��!EP��tQ
H-��). Ss�3��I
�s�i ��aI�P\aI&~ß���_�5�\4���H(=��$�H/j�]Q ���J~G�����������4W���-?�Rʨ
AH,����I�\��ϡ�^��-��*c���0�uL�A�hm١�g�vU٭�ե��c���gӒ��9Wոe������ي����!� �������!䂐P=�- �O�)�0)Ĥ�Ü��� �(*��(���R�$�Ü��LHOپ/ǳ �f����|�y+�p�;W���xhy$��\ �s�\Bc���H���_���ѬJ�t钳a�[5�âb�`��c�JM�(k�Yr4���z W����I�2S��I ���u����Qi4�$J���
@��O���׭=��f���$�X~�
B����9����7�����Q
H-v�ZAK@���3���Er�|��h���-�h�Xs��i�l����7[�n��W�<�XH/XtAH5*����`g{;�������	��� �$�D
H,�Jx��,II���$���Qi+���Mu��������S�
@�����v��䂐����tQ
H/�R�
a�r�m��
C��I�3��WZ�=w�ٚ���+l���/�G��?	'�0�7p�AH(w�i �44�^0,� ��.H)���
Ae�5�7�m9"��
Aa��;�|�X|;�-&�) �S)��,;�����_�k�����?�H,=����RU�QiE��麟�ہI1�{��i�%$)�H,40���I%�L9�\4��) �s�ZAH>��������yR՝�w��#�Oü��D|	ϖ�o?N�o��֞���i�E��
H,���0)II�o��>H,>R9E�Ѕ$H�(��T�<��^�S����Q�K�P�]��=Ű����u����A{6ߢ���d������B�N�N:ʸ��m�q���	�+u�����O{�Z^���\ �G%H�!	A8����8�&�
�z�u�+4��@m6Y�#�GVh�Z�W���Fjx����#������W+5�F��ER�˛)��G�̚�֤�͉+��5um��˜���v K)�1ƙ�f8��.�ó�)�ҹ���#�e&�uk���B��4�3�kp�6͊-C1�%�i��t���h=n�(�ݰ�>|>�ɢ`�KK�anį(F[�5���J)��c�.[*��@i���OVt��������U�QiP��Z;wH)q�g9p�>d���!�Q���(k[8��B�*�D�K���'b �?H)+��w�x�S}a�}p�'�RA@��,�A`hi ���eQ Ԩs��|�R
9E� RAe���Rj�׌��i�z��:�Xy� g(��B�%2�U@P,s���=B�|7-���>�/�@�>
B���(���D) ����R�)�9ˆ�Z����w~ܘ�P/�ZAaх$�P���
a�zᤂ�P>'9f�Q�����#�O�%?
#�N5��{M���{k39�����?@�r�O��Y@�O*�(X��
�{P� ��� s�yo�\�m�s�v��K��$��D|		^M�)�w�*�����vQ
H-M��R
X�L3;p�>d���!�Q���Y�}y�����ox~�}�$*��
H)(B�k9p�AH(��}g�h�};�}8�X�$�D�Þ��I�`SWϝy}*�t۟;��hÜ��I��
@�(���w��}��;�Y�Ă��S�
Ͽz�^����?����bAa��a�� �*�r�H:��Z�wH)b0�9p�>d����H,?kUʤ���տ�����c)���,](�El(+!�4�M�f�v�eۓW-��L�Ro�t���):�a�rᤂ�P>��f�
AH/*�}*�)�9ˆ����{����������?@�yE����i�~ο~;�W�����7�1���R7��>H)�����$Je<���ZRAa�rᤂ���r�H:��j<���������bun�V�텴21�ˣt.Nڽ*��G]��̻�X�|�S=P��ձ}#�͉�gn.����L��$�]� )?�0���4φJH(TC���I���ϯ�;��}�9���j��H.U��RR�[��L����S��I������;�)�� ������ �{�Zb$P2Sʨ
RAa�rᤂ����Qi4�$	TG� ��S�뛘��c1y�j�m �߽a��
B�T9E���]��) ��9p�6�I
�s�i ��aI�P\RAI��ç��ܯ����높
A@���i �44�^�@����_�J~G������ّ�����7� ������I��O*�(X���߿i���w
sw�q �e���$Je=���Y�g,>~H)
����
AH.�wH)b0�9p��z��j��7\����>�+�t�����
��S���P���!L5��4���H(�H,$�P.���k��$��d|	�����6���O�	�"hJ[��t*˦��͋����x�M�@��g�v`WN�C_�m�����YL��������zᤂ�P9�- ��H��> ���FC�G�g��mUO�$�?G䂐��z���8勤��R��� ��
a�?\4ϣnZ+���_KF����uy�H)�9ˆ�
A@�f�w����?�y ���UuD�U��p�>���]~�fϽ�t���" n��I�)�TII��5�
A@�(����~�9��<_�i��)�U@�) ���\4�R
v�H9D) �r��Rs�$���9�4�Xn���=~��:}噙U��<4��p8�&�$Ƥ�کfm6�Ǥ`u;o���fq�����4�!���L��1���Ђڭj�R�N����}�[���Me�z3����Ȃ�P)�7zFw�t1���Q̫�h���wk!,�@�D���omyp��E���X��<����Iݮj����Ϲz;�X��"9�z��'�4����(b!�P�����P�}�]�vlw|�<cu(����ȣ� �;'%�S3;<6��++�T�L�x�*���l\9)��Sf�lh�j3H��mb��n�X����"`�$A}���������ha�SV2�j*9�֧� q��	#�H�"��w1W����ֽ뛐�q �
";�祆�:�ܺ�����2��)�����S����G��؈�G��_1"�0�:�[���'3�-ޗ:z��Q���=��c�($��r���*;6vz�~����D�"D�����X���%��> ������7`�13�p��|Ry�F]d��V�;�ad�νCgVi��[-(����.���^�綍���Ԧ�k�x��}z8j�t���Bk�1����`�K�	�QE��}W_���h�=�T�c�3��ӇSb����C�Q�˙�x����7��U��]F�HV�����QGh�e���[4��$c��M�Z�9��>��`z �"?#��~�I�Ћ��n%�p�*���ײ(�A$��������^�`��{ˠY��f�ް��ih��gn~��"!}�VRM�����3�!��0�2W�����=�0���E��3W���ł�� 적@�/����"��n�I�}��1}}C����w����vؾS)�7� ��7�(�0'd�N�X=)|AH�D��A�� �H�;ù��q�`T�_��.o\~;�}d���?)i�7h"!�~3#��j�`�ݗq!��=s4ټ�;��p5��Z�F�Y�`(r�t��Y]׻oؼ�w[�N�uw��~,^�׿�κu�O����@$�s��hj�wQ�]nJ:�k����\EҪ�if�$з�8����ٳ.�M���^�p���	�����ě;f,θIr蹥���1cɊ�l�������z�[4��`��=XT�+�,z6i]D��sA��-���!&f�R�p����i��� ����B�يݡ�C���,��L˛� %")0a�ü����8Hf��v3��a��VV�mp˶�+�����X��4M�T�9_� �t�Rk�J��WN��û2;�[+'7"8��ѢNc��=P;�H���h�d���a�^_,�,n���)d�m�{o��S)�7���q
����V{��l_%'��4�(�_Q�/����'����w��#�G/���{��0��oYz�喘��`�H�)iޮ�B"� ^��}���Gk��a����l���@���G����i��p���LC@֠��@����6w��d���ksk���N<�[ln%Ȁ�ȿ���vn���߾�z6�f@v�Wj���Yk-��%��M�F��V��B�6�Dԗ�Ϗ��z'�=�:�~~8���r��N�z�d��KF �r��������2���4~� ̔� �0F���*gs��.����-�j�b��I��mM�k�3z�p���k��WJ�6B"�sU�)]�ي�N���.���ey�n8��p��l��|����?9���]߾�����~������
�$�"���!��;��wFA����H�e�3*�33G��Geu�]��W*'r��<�[ln%A#O���V!���0��*3(��/�Aȃ��vD����$�'�/w�����d�qe����_:s)�CD#�%ku�bGCul�3�r�����=l�eO��Aܯ���'�D95�|=��Y�m[���n�LB�Zi���$^�s.�l�HK`��ڸh�ҵT�m˹���>�9�-�ʙ��S�vWݬl�S����C�l�U@���bޣ;����U��fgƄs(>��R{LU��Ѿ?Br���'-;4�۞�Mzɽ�g���#u��x��Ђ�����L�U� >�@A�H�2R �!mߗ�\Kk���*��
UN[9��ݲ�A�ty��:�/u\j8��>ר�^feCI=Z�V6�jPo��s�i2��΍�^�� ��2&���^�;��7���t�G3/H�e�2P�{ޗ;�����������_Ηvc].Sc1�� �:��˳y�]������߈$i�D��FH���h��A�l����t�e��������Ylʨ��Ѷ��6缛�~�}��]qkaEL�ԬԎ�,���f��Z=S��ˋ����<)	���'�_��4��:�����gc,-}B�ue �/�רo�g�V"D�P����"in��?l��N�E7N�����)���}��~���݈�5@"�z�`�sh"��&9=5mR��w�ύZ��v�%�6���;W4)O�1_I`�Hw�+�8�<,���d����;ˣΟ�m�����
�Fb�f��?fY��Fc.:Y-�?	��n+w��	fT�㫼t%����=yU��e2�=㼬ɜ�s�:ۛQ�f� ��""�y�߀�A>ܚ#;�,fQB�e��[2��~�k�&��!���5�F�:���A!� ����W�D+��T�=���J��(��]�
mlQ�B줻f.�[5&NfgV)6�"������'�Q�/� ���V����^�^���P�/{jf��}@��������@�@��zdU:����}�h#L �ܺ+��;�����"��#�`�I��2�r�@��
�_1"�*�2F#���<�-��Vv���B�\q��AOhPv��!�$��4v�g���ʀ�Y�/��?g�Ů����%��<(c���%�ɭ��1�����A�%"	��ݡ_ػɔ�o�Ǿ�����o8���� ̠����d��d@�w�����U�{<�>�L�*����N8�}ѧ`��ߟ�Mv�fu+�OY/C5��UK0Zע��Yh֎�-�t�"��]�lSc�RR�dzk�W+�u_#�*|�f ���8������m���c��uY�bE�j����LxV���������h��lr��//B��Z�G����*�$FU��z�VnZ5��f�3�TS2ccMjw&2^,�r�����UڌgM���ȼW�1l*[�0��Z�A��G^i�8��L�h]�j�
�)9"�]+��&�NF ��F���ڵ��^��U%0�*O'$���_[�2�a�d�֯e:�w�E_ݢ�lC3���c�RX�}��:I��w�G�RG�<%Õ���-\H�vE���kw6���s,��˝':!�a�T{зHZ핼�e��e�s߰r��p�eѪ��{�2X��VD���1��A%�w[UGr���*��w;+%.s�P��p�2a�{1m���t��v]���{K1oQ��Z���]�+wj���#����I��E�;r.Q+/�[���8�7N�;:6&��2g.�9&ڂB�H� �`�k�_Z�u�f�M�y륷�>�G-��-���^���b�5qO-+�S������Z��2P)�Y}]U���2r�#m��e��q���{:�����X��8yv�Xkxᢊ9�;rO��o��֒�L����-
	5;:�]��&(e�d+�nrɼ���o�P����{�Qu,[%�b�Gz_wV�}�u���W�tU��7�F��UP_>�w���;�3�a�ݷ
��ݍ��)WYy6��YBڗe帟�9�qݻ��M���ݮEnuҊ����ӻ��L	st� �M	���m�F��wwK�*��p.r��.��r�u�wpNu]��8%�С�Ě)C:�ҹ���B�$ir�k���78�t�ӹ����.\��Rb������ .[��nPG.\�s��r�.WL̐͝�Et�X�c���DQ�r����s\���1�DG(��Ӆ�lh�L��� wu�;��1�$�`���������\�w\�� �wr��"Jhwr���k��DjH�3F����Fȓ��)%:�!��_�����[6U�䅕�c��]bK+��8u��(���i�=��n�AP�2�3j�\V�V��\�U��T���f�j�0]e�״�:�n����gKX��Ql̮v��u.�^l-�4QsM�6��SDK�E��lڛbXg0��ӄ̍���[��u��GQ��@t�K�be@�Mwd��]n�-΃(��+-��+���b5ZL�b]1�&��Ÿ�����C#
�fJ$c��^4[u��B-�"NHHE�� �j���&S��!͢�K��\�.�!-f��KN�K�5aa�6hs2WV2��IXT��y��lٲv�/��<��P).��Rh����mX�46&�=5��i,��/<.�+79�C#!��v1�k�I��u�� ��m�D����RMūs�Mj�8�����Q��2n&�6��Pe����ZͫT΀�����4���J��7%�d�M�O<i��@���E��5nr�)�Sk�Ik��r$,���iw&d��.�!���TiX�W�)md�Ek)M
�X�h�P�7<�r�gKB���I���ғ���N*=`�MnZƭ�����W<J����ntDɵ!a.{WFkP0H٪K��M)1SZiD��+��3�b��%�e�]���1WF�4�
�j4͊��&���Rk�6�Y�,��`ۻU�$3	J5�G\ڸ�U�a��O<Zx��"�ۨ�E�!F�Xg<�mlBF�q�� �]B1I`��Zܯ�r������D��۸t��k�7KA�j2��GfKڌ��Ý��S@�4��ԥu�j�Eq���2��S1�X�Kή��j�g%̧�3JBScK�B&��E��e�]�
Ҧ��c`�s44�W���O\������WMr�ݣ���ڣ��BζR����%�G0���c��LM�u(�	�Zi�ڜ�JX�5f��A+�R����4Y���	�0�e�.e�Ķ�%#vkHIe.V���D�ٗ5�b魐�d��V.��Kccc�iL��삠_��I$�a�١�)�2`jF[56
��#�����ֆT��^�++��Z���bVh�#6�)av1e7J̈́&��9U;\FQfÅ�����a�J�s���Eh�`��*R=l����gDD�l�
��]]�,�ЗP�j'��l�کK�P*.�+�]^:��֮X�AK��@�`bĥL^�@OY�|�|���ʤa� ��K���'�o�w��ϟ�i���V���CH�L9��va��a`�wV!K��f��e����a�?d�|�q�~��3yOD��2#��Hf�"��k��b9��hs*щ��ύ�QqP7��VQ�E�r��땭߽2�/Y/w��c�� ���:�����Χ5�5>��tj�W�+34hs*Zb�E�Z��P�a�J����q��������b#ġ�˙��U<۽z�t�P!�	?lG�n�
���dt�X����T�6�}+'=�$�j&fkB9�Z.%9�<�����y���Sk����%���;W4?���U���O/��]�me0�dWJ�fr�͇YL����Ps9���M-6&����d�L�h i�Fn���!��;�O_p7�a2r�'�,)��sS��E������"�*���P�}�/:ə��g���ܺD#��b`�k�*v)9�Zn�1pɷ�u�X,�����\�1Y�Wb��:u�V�QI�ǐp�e/���W<~gh���5�~�_���:S��q�����c�6+��&4���h�3�3.h̳U����[�"W�C�z�������;_1�� �+�_I`)|E��fOxQ�n�^]��7|�3��H���j�k��k»��6w��e�A|�z{� Gk� n���FH�"J�6�鹛��LG�:��c����Nj��?q�ޏ�+>aJ~��vE$��cPb��8R���[h"�WXM2b�5a�e�AchT�P+�C�>�k�2D�"D��aD�g��pRCOQa8�讲�M��k��@B���+�#��U��-v���I���T�.�5.`䍝���A|A ��,s=�A(�?m
���$A|~��1�9����m��h-3u=��u+��'(�3#�;�S
J�۱fV�;��1��zCO���m&�/3m����p+��˺���=�� >�ū[���W9�+j=�����`�H�D4�zo]���k^:�>"�=�� �A�s�iz��v�
K�� �ۚ#@�}�Ws�$��y�3�� �F����3��X9�r�UnU�uL��k�~��G��S^��!��\��+�$L%�%��=^�[ׯ��Bf��V	aک�L����e]خH��`go���3�;b�/z�%���㥖O�oO�����\ǯ{���\栭�p!:��z`'��k��!�$��+�)a�N���!�s52٨:�8m/g��8�w��@�-2�A�V��=���f
�J��r>�\DO4����eX�&�龄Ɣ���N��,6H�� ̠H�d���/�b��Sw����m2E��+�$c�{�����Ċ�q�A���\��Vm���QO���kF�'}�u�P���C�P�P+�O{\�Sx�{Z�Y���wՓ'wi�J���S����w�/�8��LT���!5y���*�O33>4.eq)�$��C,���6���vzS˳\��P��뚜�̪�fh�}�~�Ž�ǯR[�C���|�t�Xd�J]�����K��@q�؋�0s����|�O
B{���J@�D4/g�e�_x�G��Uhf�乹��L�`��ܬD�#�"�2D��?�����W��^��������S����XU�EU���f  �����g#\�x�|(��?���(� �$B	WդaA�^��~��	�<N���W�Z`�&��b�2F���AM�װ�e�p���a��� ��qec�y%�b.�������t�έΦ����r��P�3/B0̲���C��AL��6cv�~��.�� �<���~����v3�#ME�K7�h��B��X�r��q��17���3*�m�9�;��X��_h�v�̑�����
�s�+D:h�c= �S*����>�<����z-J�oHܢXm	�Y���bL�k�V�搉�\��@��޹��ͳ�m�W�t��%�ZM;,��ۆ�G@���`���WlYv�(��i�rK�:]clb��u�t��44s(^����������fʆ�%���Ƭ�+�6]�����
�k���P��haє�8ĥ.��e�FZM�6أu���M�Fk���߻R�%KnlY�.J ��i�A��8-ZG�]ۑU�:V1��˻�0>�d�	����׻"jUg���|NK�G/.��{�"P�la��U���J�i��H�s^��\ze�U�ψ$q���꛸�s��w��( A �d�yt݅i��"�H?8	{�P���U|~�ο+�3=�p�}��I��
���w��Ok���@����aTb�m��z�N�F�/����y��;�����}� �����3��N�CV��n�&w�4�U��1�L�ѧ6:�GX[�'#�C0�\=yX����:�Г�&e'O�E`�$_w���>�{�>{���f.*��HѮ풷Eɝ�`��0���V#.n�ޮI�V����ΰ��ϙ�<�O�~�ݡC8�}�[�����%V�"���On{�Wxi�{gޯ��DJ�g��2���P�;ۣv0��2���;Jn����K��̹j�K��G\/n6s��7V���U�`�����U��;p�D�.Y���gJW�?}��| xG�[�_~~�N�8M>S
�:���.� �ڂ?L�Kf{%&���H� �R q�2FJ_!=�빯}"/�veo_<���:�P���e ��(� �"����e��6�]��ir$����1��ġ��(�	fv���<6z��G��ϩ�~�Z18��a�d��E"�}�˧OQ��B@���:��)�\JW��@'n� ��#�?I����Ǹ.����i��4��ծf��*..�D�3<M��z�Vil�]�����,��Ai�F�A�)|A"�ފ]n>ݙ�����)�͞�J��1[�pEġ�=zD̲�bP�e�+�?k2�	��J���|F%B�z�ӭ��ܫ�	f8�A3��ح{���8�"��6� �����	���.�,X��,,��)p�y3��ut��وX�e/S�uey��!���a2D �����NvH,S�I�����ﾄ�c߽�S��;7�#�i��A�
��fJDY�
̳n7����J@���w�r�=�W�BN�L��{/4��-�L����N��҅d��dB~?lmn�,�]u��rd!�K�i�]�=Pn��x��@��2RE>:��>z��'�K}�J�®�*8���\�c�05mfрj.6m��X6i�d�_>{a�Y7�H�d��$A��#u�<�q�;7��=3�+�Q�r`�;PG�?I����4���t7Sn��Q?��j���L��p�w��("<E$R;gM�}񁬲�9R�9��	�E�c(�������]h�.�rqwwJt%v��?Wta�%|��$C{�1腋��j�x@:~��(O����[�I����l߳���L��~>�If�ަ\�u����Dh�܅u=(%�U��+E�OLr�m}�1'n�c����Y��(�A�%�ZN�)lX<�^�m�*��[����������HN���?QQ﹣NeX���"�_��㽟�a���^p隣��c\2���	�@#�Q�'���Q&}6�'H�㲊@��@�K�g9͡Z�X,���js
����B\k�SE,^��P����"g��3*�33F�fr�����uwOh�v�y�	s�58�V�g�s��C�����fe�9�ZcG����C������3PN���=�����~�.Z����?K5铽:v/����eg�G�|AH�2R ��?	��j^9�q�.�Ū3F]1�5�;�$�FH�"J�P?g�X��\�"�k�#҂�_����mg_������ێ��C0���P2%C�3Z8�ZcI��й�X"8�̲��WO���\�vC�W������~�-�� ��~�|D���1�K2�v����[q�!��.��y��VGds�t�H&"����5RS���F��w���Z�X�\�^K�����f1U[�RSfٕ57�`��6�}�'z���g�K]G=B	wP�m�j�R�����R(�B�IZ�`�
12s(�e�j�+,HH۵J´�mhMsT�5�(��g�]�;t�c��U.՛�-�έ���+��n�,�)�M�s.�Z�V[B�� m)�����"^�5۩���J*T��q�!t�/��z��
AM�8e3��٤��:���Qm�e�K�X�Ҍ�dԿ>~�m� ��\XA��k�A�(�4qe���������#AZ��������z���HA�o�G=]���5-������1�]�	��Q�#g����A2E����3yޚ�pg�B�>��͛����WtՔ��q�`~x����/_�xm=��о���C���3*w�qʔ��9��5{���W��u?<��l�.����̲�1�ff�elN�5�~u]t������N$4�.s���t�m)w�(I���2������pB�F�v��~�d��~�~�3�?%g#�5�؝��>�t($�u�g>6�ݻ)WݯDS�#;��̭�A1��/��3-��,�0��n+3�{X�R�L�uԦ����*�X��^]�����,�C�d���3�nȟ�ew�3�Euc8��/�@�N���I?�#�~�_$a��� �4�#8���{���(�T��E�Ğ��M��bP�tH�%!x)a[�i�OZ%׵��i��'a)�sd��U��mf�T|�)Ν�ο��D�2��}�� �|[������=�וw�(I���nPD�P2D����hVASyp�T1�v�e��Vfh�]���^�U��y�4��)S��A!� ��?����"H�	p�}=���dȠ�&D��?xU�>����Ef�=�|������:W��5���hd�0rW�=�{;9H��}���v���xT��&w�`�����'�H��쬇�y�^�_Uo��	q[�
�.u���e&���tT�L�XgX⛃�}���ɐ~��U���/�sx����)U��3���i�ؙbL�A�(���@��"H�&J��Cݮ����S��=�+՞�Wz=�眊��xW�Z`���.�g�.�Eo�"l0s�~#�|D�d���t�Q�7sj,b���z!�R���\im�L�mĨ(8�w��p�-��BA�em�w�.r��ȐZ�vv^�*�����:����r$�+�1#b�lU�,Rl�Xb��|k�c��}��7��V�_@�CF�c}&�K�V�Ӧt�l��XScM�rx����ee�<�c�J̩��^0��q
��N�V�ݓ;f��(yp�aD�9p;��a㆖u-x�ʙ9�l\�a41L̻Q���w�\�C�A���733�.C��fVt��1�Jյ�yti�s]+7����˪2���ӕ���K�`]6ԕ_8-�˧�H����{nQSuC#n3ui��������E�*]a{��`�ͱ�	���b0�r������p,ԅ�{�2b�\ݘ�]�V���V.�`�b�!�P���%�*L�&�r�����j���L�ѷ�>ƺ�u���*Gk�o78i�u6�m���Xh�i��x�ыU�����-l=�:�;�n�{�s5y�Dɿ L�����/����q���Wη�4�e��n��rh�!�[��M�K�{ Bhӌ������,��WM�9�?���V7e��qi�9+8����J�`�uQn�hL�0\�Jݧ�܎��c��D�-m��z�������5܁X�i�>s��˛�lD��l^N8�{lts=�Ⱥ]P&��򮝃j���W�!ՙjj�Yv��V;�}#�{�P�s��[j�T}�qr�d+�oWSC�J�ei���o�z��I�VrĨ;���0\�n�"D���]	�t`�=�q��2��i��h�zH�QII)�5��2�n�������1��U��C�W.�r��������wb�k�lS5
��"5j�\�K&�ݘ���VQX��	�HWwd��&�؉fa����c\���2I�$�wvb&e!�AI�2� 2H��BRHLa.q� 0��
D���� � h�E
h�3fI&�P+�#4ܸPh�")Be#˚�͆�I�W9�3f�˻:���͉)ۺ�JcH�h;�(���APQ ��Q��@$�߱v�u,��
�|2����3(��(� Ȃ�GK��k�k([ǯ�ZA���>���z���|i�v��V�$3@��o�e A"��"("	�W�H��G�GׯێM�B���m/e�5����r� b��!�x��{z�.��:����A�L6�z�Z��\m��1�bV�Ց��
�3e�͇8�}��O=U��` ��-���8���2���;�Q�Q�z<���"����Ⱦ�wv~� 弇1����#�x�V;�V���iڲ�c���`~ohPv0m�����O�K�k�=�����d����b�?Ql������-߆����F�~�.Z@�A ~�_I�V��[[F_��e��~�o`ΤA#L[��MC���r�ظ���܁ �2��8O&��3.
ׄ��1=]Kp8�¯ܯ�̍)4l�m��6�s˧�8��WQ����0u��L,&��6A�v�ՇQ{�BstaT_��}��-??sw53�[2��e�ٍ̲f���QKgە�c�A��)>��K�t��Y�� �F��@�i��	o����Gs6�H(�BZd�m2!�aiaFࣥج�sR��v�%�\�k�PN�7��0��,�'H�d��"_�{����ի������kr��o�F��=�#����`�_"!�D��{���XUW.�{)H��}4Թ��+-����P'r�A�("��6R����G�U�ɫ�"�������|{�-�r)ѹ%����v��y�����wF�� �$ڡ1�����/�[�]#��D�PB���w�>�^���ϧ�寷fA�lX?eW�f�+�D?T��d���ƋW0���F�Κ=�����b�nw�&e�?I�dCygiY�㕁�mL/2��M՘ʔ�o�n�d���:�8ҦSu�bnҜ���ϕ��wZӫS�b\�j�-���#b~� >�+`N�K�œF�v��%[�����S݇l�#-��Fm�U%�紵1Ҧ�P�Xg)m7cWq���G9-56U��6)�[+�Gm�L�	��m7l:),��&31���)z�#�ɀ�$q�#SrB,q��lG�\E���
;1��R�\57!0 K-��:4�Y�R:�u�F6��͙�KkMW����(��KA/���������P�Ѝ�����fj��I]
����5��\%,��Su*����̽#��\fQS3,Ѿ}��{��ɻrԔ�\q�8F�B<؁%�gv��~�X��M$Ю��b�j=�H@�٢�O���^>����iϧ��-?�;�/���Ů��{ޜ��}�q�I��3+b113��23�,�d�j�n���b�n.�A܀� �"��/��|#���vu�F�#u��0F��
�H�:�?{Ϸخܵ%+�w�3b��Z*$kW��~ �4�$B�����ad�����E߷��(
�-���n��U+�������#9�.3*J���4��f��=�3������Kli41�0-�`[Pخ�si�-��n5��7�4(6[��Pw�_h""���V|A��1k��l�u���b�n.��/bڤ����,��%~�@�"`��7��D�	)���������/���� �g�6lJ��.�[�<��⻣������H&5��[�8�e�۵������u{]�[��l޸�	���Ԋ���B=s�|TS���鸚j'���{�,Dq)�˚�5w{���3��;6�j�t�F���{����Q33F�2�MC��x���I����|0�֠<T��7w�P���Adeh��U���d{h ~�@�d���#��Ҥk'ϯ���3z���렱��9�>�C0AmРd��xu��wd�uV����ykؤ4W8薄MN��
T�\�@�vr9���mol�����	�d��%����{�V*��US��vc�Z��Z�� �|��?P�0̕���AS</���c���I�0/���a�f�U�qx0L�A�("�^�����e��ޯ�}�� ��:�H��Q%㞤�+/�r8w�A��q�3Ŋ�Pj�~AÜ��|My�F�~�o�"�ް�7*gX�W�$�Г1�M�З�1u�82�Ѥ}�z���ks��|y9/��N��Ʈ��q��f> �u��}�i�7v����!C�ځ M��?Pݑ �>
j�td�m�1����6��\-}U/U{�>���ʕ=�Y��U�SD�0̕c}�'��y�ڀ�D5���[���<���Й���fW�H"D�OY�`�!�Y)���1A�iN�:�0�HY�̺�`ܤ$
Q�.� ��I��4q-j��?�8����#�7v��ԯ���ԋ�v��&&�ȣ�/z6��QuP�_B �!�$�0A�� ��:p��wq?�?MAgxjw��b�8y�B=��w�r�t}_M��h�{���i͡@ؐA#N��(�_���5�k�^5�����<w+��"�~�~�t��>c۞�1��A�?I����֡'Iƫ��N;�@F �T�'�,t�ꚍ1�����y��2��иϰ$~Nœwˁ�X�6�U��uK�E7?V�u�-�K����ȩ������~z��8�ff�.e�33/�޿h��xre|�H9��M�����z�2Z�Ҿ��������n�{�ߞO=G'ٹ٣�: l�6�X�&�nݓl���K�%Z�[n�����#���$i�;ps���u5�X�P����mѰf҇���D̲�eJ���>���7��v|; ��"ݪOz�u�e]��q���ѭУ��L��t|�i=�ѡz�Aħ3/H���y�g����Y��x��Ng7�G����u~�_I`�H�qùW�I!H� ~O(Q�/Pn�#�74����	ܠ�D��L���{�8���c2�\̹�2�fn����p��;�#o���f�W��=]<�]Z�U�M'A#Ms��%a�!��¯|«m�7���"��J���7�nc���%ׁ��ə��M&9��r���]�q��v����3LFu�֮��y��|���ϟ/���߳�A*I��a���`(��G��$h�1��F�.�9�Hk���5�u�f�b��4I]5�LK��j��:I4���
h��s,UW4yp�*S.��&+�65��&@�d�f�-&��pG'[�r�[amv]-���a�s+Ke�"4#��"�H�[�Cm��h��tM�zث@�&�Iv3�Δ�TqX��)3�e��A	���0%��ܧ��j��W=�G6��]p���\h
�Θ3F$2f��D��6O'���$>�f>DA�ٯ�;�$t\
Y�*��U��

����g���,3���K���ξ2F�� ���s�>�6�7�:�LpƤ�s��,\
K���@�	DW�H�,����$H#��W�辒����H�����$J����-����ȑ8�;�ti̫3,���&�&��͚ �ȟ�\��Y�6���w��8۟�5����(�0��%G��el��#��4�S_>��M�2,�X'+[�f�K���t�$_9��Ѓץ�����!���c1��k��fRj��"�-;j�R0�F�����I�m����T�P��˛��ʨ�f��	z;��굲�2k\w�j�/�鈺�~���g6��h�#`�d�����:u�$v�5�w��Ŧu�B%B刻{����"Mֿ+7�U��J�7�/e�;�[wQQ1�1#1�X�;�D
v���E���>�#��M|A�{��B����j�z����A)~ַ�;��u��_4hyʴbq�32�G2�F"a�05��ݝso�v{���~G�����hc��l�S���d̲�1,^o*��u�����>���_$�7��/�ꮫ͕{�Z��B0���}��>��W�֓342��į��'U�[T���/��jg��u�5�����^���Ylʨ�fjw��~{��"fa��;�bR�CfW!�c��X�!J�r��T	e�E�,~y��C��a��РwbH$i�3����8M�t�2�����{@�]aT/�	dQ�ɂ�#�?n��	�GfDބ~G�}"�ožƧ��e^�ָ�$3 ��E��\�5�;+8lO��f�1稴Aġ̉�AD �Q��j�ٜ��Q�DWE7S�ֺ�yu�.=>J^�o5t�uR>ʵ�ݭgfzH�j�1ڸ�/tJ=����W�ҵҹ�6��X��Wt�*��\�g*gy\��M�~�~2�0A؋��fe�e\�������S�w�}̡@���A��08g13��t�5������=�}ݭC����'� ~�Q�&��S�{��b�9�h�ؿ{z�M�n�RE�-9����DӘ) A��oc�X�&�]
)&�l���%.ط�M`$гp-�a�
vS9�:;��.�N�41�h�G�C��53,��}Õ����z���}������2� �r$���|D��d�A"���Q����R�Y!|Z�C���1j' ;]�Y H(�wf�/Zxʐk�^:s�\g(�g�B&e�3*�fY��wv����iJ����\�bٖ�v�"�j#��eX�cBfe��}x'�Q}|<E�rE� ���n����'g��g��v��1�W�����V@�1Zh�������v=�m�}d�f���ay�:��w��u�Gs�]u�;P�l�u+��{[Ȃnײ�̹o!	y��掌�*&��F�ʗRff�eg�o���{�� 24��h��^�1F��7���;� �"�2D�D�ԩ�z|���_'��=�.�K�sQ1jF�dY@�+j����f��I�j����I��4;���==��[�v��y�F���!Wq�@���p����=�@�D4D��~3`	5YO4�<x~�����'��!���w<����~��L����^��ݮ5ܙ�s]�DS���ѡ̫F&7���=$T}+��:h:�'(u� ����(� ���v��.�0A�/���RFN��-��|��nu}�G!#/����Lh���K��Ϟz��D��V9��32�{����GP;<A�h���;�Lt/�}~���d����Hǀ�t#��Wf�+�ap�D��2#W�՚�5sdE�D��ݥ$.-��h9}n��V�媊����*]w5q���j��ɲgc�vC��Ξ�{B��+��G�|��h�{YY2�B�*|l�'�����ڸ��KQ�O�:;��C*頻Ee-��^�ڀ�k5�+)�赏J1	KU�B�NU�JU��h=9"�r� ,���%����V+��ܣfr���7T6j��&�Us!���������!tCd.]R��T�"��*���0ƹmq�ma�fԚ������v0�w�{)����h�	�%�AC1����8n�mΥf��V�6Fٵ1M]�p�*b����I��CFnd�9Y'H���w:�y*�7�P��Ś�huR�T����87��w��w�m��Hż �¯I'P��=�0�R^�;��T�PQ�ھ��B��me@����d��$���W#�w��(�:��UuT����*�v�yu�G�yr�ҥ˛:�Ҝ��W0�����mu�D{/bUh�F�,Ũ��[j�Ŗ۱l�l)ua���t���4D���E�MJ$�7u�:,j��B�[�SM�Mըw����L� �J�W}v+[�g����8���@v���a-�8j���Y�]Ik��\ƣ�.�&�
���������GmFBz��"j%=��*�R��q�%��o(�۱c�mN�fQ˥6�T������K��X��2
|�6�v�+�o
���ĺ`�Wvn�8��U0�ℯ~d�;�<�����c��O#��"G,=�����n�un`�ވ��O�)���}�hhH��wv��I@�w@�s:��2��DSFI"I$b2!"�U�2*	1�@I4�]ܚ)4(h��0I��a�"\�R�sr�d��JH��BIa`�H1J`�a�2�%]��v�т2��A��A%A���,��2)�0!�D�(wq�$�(5I�L�����ʉB#K#�MCS,`�LD�MAw]�h�JF�4wv1a.k�)Lib��̀�R�IM��J �#6J���6F�����M ��B��d�e9�$�d��wt�"H�D�DF��#E����c{��:�Щk�D�u��!�f���6�HM,ա
p��n-�R�-j�RR:�60���!A�`h��
�#L��Y���	�u�5��1�m�JK���I��
B:��{Ei�m��3.D�qKbcU4�)��:�+���v*%f�T�ܑwb���.�#��6�hѰ�!�Sk�	�\˭q^��Ɓ��W�:�5M�ۆ�A�B�8ىk�aG\V��-�Y��#�KL�nR����a�cBS�5p;f�m�Ѡ��*D1+(Z�u�!D��kSf16+bĳ.��j1k��]�L�L.�l��� 6�ef&����ފa(����K��l��f@�&o)e���X�f�6����y)�v�����#��=�E�1VћE�
��klТ�a�e����;�k	�Pd6��2�I]��������qw*X�fก�-n5 X�q�V�m��m�r7Y��S`1j�5sq�� �6��6�+��lE�XCB²�!f�n�m�ceXJ�Ɠ$5v,�����R�,�vʈ�I5���u��]م�<�Y�B���
XL��غeu6X2���Sn�"#���ZL�:�0��X��,����k��P�ĤS�\��Z�1����&�%+c3��X�uY]��
+
�5KY���f�BB��n�.jB�d���e�\�u��.�2q1��Yp��]��Ʈ�Le;"�9˝��-�@1=n�S���Kj�
�)C
H�&�A�M��f�b�^E1�����:eFhŤR0�3`]����#lt�cJ�`��T0;C�ژ���<룍�r�J݅¶�`ٰ�hi��t�I0��L�,���5ZK-�zkBhʒ�E�b�k�VSFL��г,Q�Z��i��)��E�1�������+
�FŰV�D�%5����A�ipJ�+S/i�	L:Kj�)���&*4��L�`�g�ћA�� XD-�m����0�C6[����(��!`�P�P+�Rڮ�GZ�*\�T���g�O#�����9����-�ZFZփ2)M4�d�m��lq�+�8	n���m���,��J,��d�J�� '8�2�����u*�.)���V&�����v�
'\�X5�.�7�t4YV��M�J��f�V�^>v��5�fr����h�
Q�"�� S!�5�#��4M���k�n8vD�KL��gbX�(�eب�k�(�'$t��jL�oϿ��!ò.��(��v5�"�7L fV�R�H5�Z\��]������'ғ��a甈װ��oy��~�r�>���	K�����,�� $��$B��9ܽ�a�Y .��skz"s���w�vv���� l���/&�M����{mz���E�L^R(���/3ٮ�&:ӯ�]����H�����G���{�Jþ*>�뙓�nN:}��
-wr�43mgN�n�� $�Q��lV/��),���˻΍(��_}ݲ_�[��%T���GUoxR\v�X�ʶ�4�1�\P��LGM3F0�h����eL*H
��nWݴ$�I;��g���˰m>�~����{��_����H����F\C���7��t���H����Mh���'J�e�#��^Y��$�X��}�,�t,nf��[e�j��	����/@�#�:�z�N99Ͻ��}6��넺�.���N�ꡝ@gD$��$�w��!��u�T�M��y�%�7�N��RPT�Z���ظ���z��$n����wN��<��}�s;��';�uR���������I患Wt2�ݩ�5˺g?S���G5���}6��!�x �篻���������*@4��K�Zf([6��p���L�D*
�!��_$���bꒀ���-��i����ٙ�[��y�݌�Ճo��m|$�" I_f�ͻ�%d̈wP�r�ӻ�O��w�nd⁻�)c=��}6|W!�_wT�	+�%�����m�<T<��wm�Lpx����U�ɱ���,UR9.21�G`�:۾��G�����]i;�+�
<�k��Vt�����Z�%����{Sd��U�BۃG�,�N8����%��b������D�<�|'-����=I;�����+�(	����-!�XP�w����rO>�gL����@l�IW�9m332����U^��4U\cmc0iv`���K��z���k���)�)�T��?}�_�I`IC7hקNF׼Z�fo_��.�����uYo7���wcv�wdZ��
�������;�ɹi�u�cș�[�p��۪��q��ʯbN�(	(I�y�x�?���O��y�s'u�ٜ��Ფ��#v>W��y��غ~c���;^0�zY0����G��\j����@N�誼����bv# ���+��	-��ܽA���݅T�mD�|4�D���}dm��o.&x��+:�V��Yq�
��Wr�6�$���ֆ�I_I����jwVs���c����D\����y39O{}��#v7n%��Wy	`C���1:a��U���J���i�,4F[�f���̯���?�WͯS߽+6��/��=�ޫ���o;��9��9b&UTq�3���#�}$@I@I@�C��Kr�03�}�]4���Ú�y!����}6����i_����I�c�{�N^p���e)<��{��V<�|3�t�$���$�iX79����99�wk���.7��a�Y��m�w8��G^h�k{|+�n�ך����W�H���m^U�:���j{�q��TɧS��+��wo����3�u�tR�Q'.�:�k��/.��^'�_�B�ή����n������*��W��z����l�
vU�uA��6e#U.��ar�}o�=z��c��h�Wl[!�
b�����k@t4�5�Wq	x@���7b�������,��.b�C�v�[]�`Ь:ٛIB������3(��33L3[h�RJT��V�u���fu��Ҋ�]�V-�%��h��l��r�B S����j�mJM�[�tL;��Z@mWdA�'j��8`6.�WhLK�n��R����ϓm��=��Х�,qa�٪��B�Z�[	�N�-*���2i���'��_I@M��<�Z��v�ۓ����g���{unR��]�%	"J�u��u������|mo<�	f:��O�cu�d]A};-���K������I@I�t�UW���{'b��M��@N�"�JU�*v�Ujw[t7v{�m��{��j�99����D1��ف{�n��z��%	*H��E|��MB�{�fsx2�u�^H�RT�q����Uiּ]]�K��M���r����)e��L�+��mB�%�e4��c��J~ݏ���Lc�ٛ�3��u;��e��������i�+Cܸ)Qz��/���4�)��ҏ{t��ؚ�۔"�)]�Ա��Ǚ����0hwF��[3�œ5��2�,�t�L,���[6�v@���y�g]�8��>�|���λ���5!Ӥ9�כ?%����vbz����	�Y}x�V��UM���RW�W�E��A��� +�J۰�m�j��n�n�q��\�f��!W���I_I�P�뺭l�]��om�s̙k^;�g���p>x�	+� �G�syve"ۢ�H�lW�SMJ8�v�� ����e�ېȘ3fWn�K�������T��7g�s���-;l�,Ƿ��-.�Ǉ��_u��$�JJ���ۦ��P;P1Yɸ�ȉ�ݍn�+���}���3�<N�^����耒��$����S�S�9{������,��ܔ�4,�����톤�53D'�y��+���մ1BSֲ���u��[����j�+0��׏-�1��v�����f5E�)���v���m[m�ǖ���L2Uo]B1�>u�s\}��n��wwow23j"��vm�!���)��;0�쒧u�m�z��	=��0�{�[Q߼״��#U��e2Jj�Zv����-kCt�R?$���q}�~�����}��9���vvb�c���n�6{g*ֈ����%	"JVq��B��mݽ�.X���(ŷ�F<�������p��
�u���dY��@I�E�~�r=�N��j�0k_�}^�4�H�u�n��H��޳{obxWO|J���]<�=��;-�1���pl`&њ�r:/&2{U�*:9;/vc�%k�[kk�V�}��r�R���R��Vֺ�L��c�ŊͯN�6P�/����%����~�GK2�'k�Ŝ�1Z2�=�73v�c���^�,UX��y3�WSh�A��N������ڵ��c�ԕ#԰F�a���J������,�]�����6h�Y7ܽ0ҽ�N����Tò��.��_IRW�D*��V���\���gt��l\s�λBۈ�}���<s�Ɋ��{��B�Bm��J�/��7�W�ȗY2�}�s�y�G��<�L��%��[ڪ/z����|=1�}��4SRok��J�b���6���ئt��2P��������w���T�Ve���1��{�<������\�����H��^���X��gg-Yv.�SaU���$;0�P��)���M�9�x��i�Mc��
��ĺU�%�d�%�s0�Sa�R,p�͕���BVTf�j�DRbʹ�J��������v.�
�RK�0Ƌ�;]H�s��c���,u؄�c�dqu�b�TsD�á���B\�¨�͖����-�*�ͣ����@��R�@��f�&�8Զ�p�mF�=A�76�T�m[3���]\8
����Sh��;r�%Z�	��̎ڛ��e��t4�)�]�I�m�`�'4.�Bb8�L��&X�@u�Z��|6WJ�/���۞��\��k�|�)�}q�U�������$�JJ>�%����e�9���N;P���}[Ff�l�y�\����b�ГE*�ZS��H��M�6ߥЭ���,�wg��FwUL�}�C��W�I,�R�y�U}�P��$����2{3V���v�}3�?��ה�- vt����Ov:�s>W}���o�e+͊wg��t=�$�xz��:�I��QM�R��*��L�����cgJm�]���Qc.��fͨWy���h�݀7w�%����n#q���cf�N�k��%?$���X�Hy��[|�9��{�����>ά��q舤�P��ѥS ���*�r��u0{��f��y�Nu}��c[��+޾_�5�o{�����r�k��@�Rܐ����T�����$����.	����[�7L�s�&�1l��+R8	)%)Gǆٺ��lB��U��ӽ��j�N�[ʶ1�����؇)�<��쟇t������g2��tPJ�U��\7w�)@�+��nd��)@	.�6;޿	0KH!�ۢi7D�[�BJ؄I��6�P+#�卋��ꁤ��Y�E&)�-�fp��廳�J>�B�[��&�3��DD@��t��V�o�pnBI+	)��������pjq�S���yV�78�}�w9IF<�ݭ������bR����۪����F�����2�%I���-eup���X��[�q�b�)��p��k�3 �[�J�37VC{�;�Q	/�]V����-��2������-���K�3k,>w�\�aU6��L_��D�b1�V���A��p��ݱ�½J�AaV�+])ύj��`�{8�1Q!���K�Vk 1����6�iQS]��E���tj�\�6y��X��!��է*�:�:�)
��*����F�+)T�'�H=o��F��m�ތ�u֞8��U r>ָ+l��:nG�w,���WR���t�G�W*%���GRyB��n�ou�����	i�PY�;��8�g3z����f���6sY-�Λ�m1bJ0��N����KǑ@�kY�L$��D��0�**`��@�ix/r��S���d�4�sX�nbޠ��/����<Fɸ��hV�;Q��Z;z抂nƑ������8����Ί�'������h�``�x��Qw�H���w+��wt�f*Íٹ[���v�!�b����`ЫY�ۑ1ݽ(UU�����<�f�H�r3n�Q�;jb)�k�6�Z���8I�+���:^i�Ϊ��3��J��:�I�{{���s]�l�h5�iɷZ*Lմ�S� ���UQ��{9d'y!��mG͎�����Ni�i�ΘK��.���Z�Ҿ��卾��x�+g7+.V`,87�*ާ'�����u����n���	�1$�˥��3�5��un��ުEn�i���Q����:(���	�û�&�,�Ha�CQ���s�!4lIRh�!���$��	`BF�#RE��[��Q��&�&��s�wu��b��*!� Q�vlHd(1b��$k�颒�%ˊ��F#I	���ʋ�2Y4D�21(N�n$��
2h���n�J�w �)M\��"�H1G.\�w)1�`\�m��	�F���((�:$��0dLY��!�p.tL��)7:B�d66La-AFn�p�cRTV`VH�D��"w#��4b ɨL&H$Z;�4�ɷwX̤�A�IQ��Gv��"LFb"1E�D`�"��_o�3y�n��*�����N��R���)�ܻ�w�djs�J�sϻ�F���S��}���s�EĈ۞���T����R˳��F-�Hto�9�ۥ3���[Y������IHI�EPꡄ�j��5C-fty��f%u
�ؕ�X�U*��R�ܙ�`�W�=�nj�}_n�wT�I�زK������Q�V냜���4g�cR8I$�%�U��^[���q�o��B���]��^�����΋��P�:��	��I_�+�b�*:�P�����u����؜o�;���(IK93�:�y���S���{�9�|��譖��k'�eyf��v����+��c�f�|�������/^�����}Q��LF��n8e���*�荝(�xF��^�L�	��)G)�b�t�\�t}��$��$�$L��_u4&�:#��̶��B���]��^��.I_�%�cz"�
��Pz����sj"��Xm����	�ɢ�Ʃ�F͢�D�X�Q���"%�ܑ��_�'�E���x^=���RĦ/�'!>����S���}�Ӓ��e��|�坺��+6�S�;:��'�~I��Q#���L	����� IJJ~	Q����LTv���YY�ˍ�x�]>^��$���+5t�b�kP���]%#���v�_M�.���}��۪{ǆ�M䓛sїu�yBJ~I%i!�����ݙػ+*���=N�}�g�+I`��v8DE�4Aũ�^㹙3.�g6wU-��ֱ����h�n	�W���6��J���`����jc�!b�]�^j5��ڪ4#Ůɭ�q�j��v�L�v5�E�]ZA
n Jj�-�h��V�P�I����ݳ���Rb�]�\M�2��u�4�!Ųf�u!���R4�g�5x�% ƣf%�[��`Sl�K���de��Sh)��º]u�+L�Ga��݅�R�&6%��bfZ$f��nr�ņ��Ԉ�6�XU.�GM��ӝE6�M%���n���w��.5��F���L��ln�,���`�Q�u�@H�J%U:.R��(}��wW۴h�����h���Z���r�uu	�C�6�ޟ�JR�Bb6�0���)Ʒ.����S��+[�������Z�12	��`]\����I%�܅��X5�<�/sر��*�˒���}�V�|I,���λ���w?w9�)�!�>�.0m��t�+���q�C��[˒I/�S�S:��j�]���N*=�䮧��F��}]w9IH	q���ukq�}-��{�E�:����ұ�=uB����i#6Yf �r�6B��QaTkR��' '�n��n��+�~YO�!]�ԲxaD2hyy�z��1�PR���J>�t��������]dB���A��<����i[]B+DWT����Z۷[�۔�
P'M��7�m��&̸�c\r���zlN ���q����)k��m䏟$��۽�g�'�J��h#���R��>��g��MQ�����w�	��s����J�9%��Mv�P���?���]W��l�{��d��6!(���y�M>Ͼz�X�|R�b
�.{��igv.����7\����^�}�����$�䔜��n���&���T�2Y-4H_3a-X���r�u#�Y�h-�iѢ�tѧ��'���v�IOZ��k8K�oaجM��f�g܌�x��R��%$����d�*6E�˜[����-��\Nof)-R���QvE���R�|I,*W������V��1s����Z������/���7*���M~s�y��H��,J�h���դծ��Z�k1�n�*��ZL8��1�u����IH�IX�*E��%�	)ϯ��p��ޗb���:9*xvwl�1�fH��J~JIQSG��՘V2�_3�:��7����R�|��|2y�=�a�M���+��� ������fCa1��k�`����{%��>��ĳ��	���>|:2�����ҁ5�_V��2W�e�{�>IJQ�JU㪫�r+kc�ڭ}Nks�������Ώ�zBH����|�O��?�%?$��$�(��)0lkQ���aNo��V%|�I��;�x5����@��&m���p]\=���0��8�.�������5+6N��VC>������;�%WCd�4���/�%�&�G�U8����W������R=k�mB�p�k��|�����u�Y(㛑�9d�����V&���v�������׬z���ϱ��b�fYc5��b쭹c�D��iS ��5�MXmIf�"�{�'�^�'�	)�$�⯁��t�Π��8��N�ߞ�䔤� ��������@�����Ǣຸ{��|�'��ItS�fj���"���sns�I+��7ڲL�	v��g1\��R���V&���v����PRj]Uȸ�����s�II��`��Q�y�8j������vǬ˧Y.:��>�����JBJ{\��	�t�)湮�\�k'���69�);��ۋ�����Oeڜ/bG.�L�]*�4��]�Q�C7P��&m�e$����cw7wA;����Y�6A�J�B��*�T�t[�c0	�٪6M��k��e�W[PB��]���$�`�6SSf�R2�ճ���rf�ݰv�Q*!n��\Z؋�.����խhYV�(�V��u����	B�k+��,�:�f�VPF���V�@�6]4�9��RҖ�m�.4�5�;@�X&0�e)�1Սi�
�0��m��6�#��2�YHK��[z�=�E6S�)�Y�1v������������J�F]Hp5�hKͥY�a�aѳJ�nR>72�U��gᏧ���k�E�Ӯy�.�co��Y�3�q���ɦ��%?$�^�}�*�k�/�W#WI�`� zOmgPaN�}�^�ؔ���^I�
��Sܳq�JBJ@K�s���Lp���M�V�u��d�RJR��1��\�(�+ݐ;�W����c\�z\���}�\��B��odp�������W%o�܍|"�A����
�{ᗳ�Z�%$�GT��ߟ/��V��8csnB����[� �ש-�z�`�`�3L:%S
��T�}K�f��g�}��v��1���6[���N��ht0�� ��n~I%a%?^�˝ڼ*�F��g���-VD�:�ΜZ���\��9:��o�S֞�]��-A��ķ��$-��ymE`b��Qx���ٙ2m* ��;�	��ʿt��}������o$����I�h' M)����RK���Cy*.��֪B{yHaV����T��|������V4�l��O w������#}=&ës�����~&fv�:%���n~JR����$fɸi(�m3wٱ��-0�bo�l��BJ@K3yJ=;Փ"DL�J3D�h�	Fb�є8������[cvbel�ں�5%O}�k�9BJ@IH5��E��3��C
�8ڕ�WuL^|3����% $�% Z�g��
j�#��-��H���n�M��6<���V���I�Zxگ���]}�ҵHJ Iva�yQ`��ם4x��-��Q��[zYWx��z~�"�9���6B�r�NT�L���moU�;P�u��加B��M�Σ8�:x�-��65�ױ�$�w�ܒςQ�J:���n��F��g��5�)Z�j��=��0�s�{"U�w�j���Z���R���|�IB�5���o+��Vt!����e�Vkq��?|�>IJ�d��X�x�t��䚠��U��,��u;M��%0�!��#K-ثĸ-4\gz�;�Ϛ|֕��nk���e��f�7�i*��4�8��ڑ������O�d�e\������)ޟ�9���Qu��JC
�;/g����_3G���fౝ�+�@�����Kcx����3©橆�yY���$В�I_�:�zv���ϫ�	,�|*�l���Y�I�lL�ܜ��)V�ʷ�S��|��7�Naz�\<����}c{sZA�/62����goT���s�v�y����}Yo�򕫪ޅ�م�ն�;R�.	)	)��Xndb����\�I�T!�g�)+���B�!(�%P0>�b�(��d�FɊ30Π��t�"�h���h�0h3PХ�t%P5@�Lr�N~IH	@��4��	yY��}$�;�O��B�p�u�%��IH	@%#�ɛ�7�ul�����op��/e����7�v�÷�$��$�G#����?�!(	)	'��#5��}�j;ND�JC
�8e���HJ�$�>�5՞B��w)��N���nv���wW�^�_�+��<�M�	BJ~IO�rҌQ���ܸt{�r��X�et8i�v��))���߷
�w ���eM�!�P-a6��LNֈ�JeK��W��#�TC�o���
���1�u|�MՄ7y�P�*S�6��j�-�]Kbv�6K�R)a�W1��c��$T�p�׌6ͷIC�Y*�4N+�O��z�1L86	a�]|e`�M�{�Yg7-+ev��l���ZD"�����r˝����G1j
�d�pa�Jaߦj�S�*����9T9Uك����{�ǖ�"Ӿ�Lyi�����"'�7a\n�TH��ϜTq���)ګ�U/Br�U�&�h�uܫ���|��o�`�B�� ��.���fة�8n&b!���ɧj��B1S�*�,�Wh'��fzǅ|v\��ƃ��xۓw:6$8�E��<E�p��-2��\��[�{-��\ܻVһO�,�2NH� ���R���QݼiHJN.�p���$˻"8���=d���8⒒��
j�F@�6L�Yο���Zػ�3X&�V��%��;���cK����r��c/9�ȶ�N��l!����!�
�ŕX��.�]�Զ�N$Qqb�YJ�C���Z	��B��J�y��L�Z�P�F�[t!��V���ub�O��,�Y[wy�%�x]f�W6����
�y1�/��/^��`�٬����rm�¬%��
ޏn�(3-B7���t���a{�09TͩE��J�A���t�Hm�C�=.��#D߬Ia�Gζ�^Qte�΂o3�*�7z}:��gf��IØ��}3��}�[w�b��R�1
e1�E��-�f60D��Dh�j(�,���IQ��f��&��%��(Ɖݹ�P[$�8�H*,AX,j��b�i�r�	�lRb+�4�Mb6e$X�jM��(�����,`�1�F�������Hh�AD�������`�Ƣ�$%U%$�$����!�ɒ��
(�Ѭ4�IfspĆ�-lb�ŌhdTF�I�dأC�Fѩ6�H�I�(��4T&4�ZLd���DX�5l�h �LRE�"�+B�ԕ�
b��%�
��mlT��A���[�O�^M|C�16F�8��e`YH̅�J�hд�c2��bk�Yv�`�b�È�5��1.Mpf$P���J%�&�ƪ]�D�q��
�+he���V� ݵ7c��[�m�@��Rl��0�����w;Y�5l6�L���٬���c4Z���Z�2�Rg7i��*�u�Wl2�.b������غ������r��kL��*]���%�@�B.4,9�7hLGp��h�r�k4�G
�,5�[�H2�b,-�4��bAkV*EPu��alh;D\�m��\LgK��cI��lKc@�]�C$Ī:�`Xk-�2Z+b:6z�}0�S&٬i���X��5����2қMv����WF�{nF
�ZK� ��Ι��%����bbj�A���.CH�h�],%Fյ�;fjk�a�P���va�5I��Ѷ�.e�0kl�pjA.βZJg��A�)ʺn�eGZ�<�[��(�Z��B\�6#��X�8��(F]���6t-�h�Ô�v	�T���z�h���.1���X�F�+�L�g��Ý���t�@�(�n,4�ZW#�l�����l�+A�mŬ��æ���A�]�.2;K1�mB:�&�bV��\ֲʑ��[�at!�A	GP�+U�XFG3�2����Ƣ�i����p�9���R�Ԧ�#���ժ�W&�5!�h�9��+K�,�]U��iM�[�4Z�D����Z�n�먣x��r��򅚶c`�tD�K1�4m����;	lE6�hB���ĉ���9�u�D(�df�0���f��fr��)��ł��0�k,�J철����7R�R!�\"�ie�v�%�i��j�h������S`�%X�v�6š���*,�UI�wmr"��eJ�oih�YC�k,�.
��#��4�зMe����c1�0֗\rQ�kc�GQ�1��ZE�eқX+�X䄴l�<�+-�#��� �٤��9�,j�� ^p�Z�63SB�(�E�F�]i�ژȀT�kG"j�tYE��Ά�[�f�S; �u02�j�]a����m���ե��Mn2�"�ڐ!����o��+�u+���LYX�%M(�,"A%�jY��i��t �]��� ���.�e�@�(��`!�\CT�YX2�+�������jjtF�D�)�XB�k	\9lZ��K�T�WFڙn=�� ~�bGk-� ��vol���`��٦�B!���h0F����O���{�{��%'�^�¾�=�d1���.�kMvv=�s��$�Y�PFE����r�6@J'xU�'�e��e���$�=1�!��2~ހ����� ����֫��U
��wyetj���ܥ% %	)�ˣQ{<.w>�$�����)M���JC{�^���1��&q�k������R�F����!9���gs
����lV^kq�-��VUs.-[e��'���@�[p\��Ye�	�5�X�2������
�i��h�_X���g��n�?p��%�Y]�ε�.�7.X̌<#@��O>J>IO�)U�;J�_+F�jY��Jd�����]f����a�0�uC�f�6��c\`M�Fmv����pd�B;6R�{�gV|���C��6Ե��<�}F��!������j����WP�m��e����RS�I�Og8�FM�Q=�r�����7u��Α��IH	)( ���5��Rږ�%#s_
��[K+��dk\\HdnOQTV���l��J~IHJJ���Uwy���ܷT�۳�ڨ1���e�I$�u(
t(z�SԮ��Vu+����0�C�m	@���̨�����M&��������ϯ�~�=�$���Sr{9����n���E���0��	)	@	)3�%��3>����Wc��jzm�k�q�>��鹊L����^��?v�JRM8�o��vNwU��Ǽ�R��N���+�o]��&��U�J`卪2m�^Pp3rm���Gm�Fb�Ys�=a'�J�l!�;��[U[[���Nm\x㇓ �ˁe핏U6�����JI%��֚���vO^e�����St{:������1�	�8"Of������)	BJ~IHJ��$�7��֖V����ָ}�wt����25�e����ETj$L���i�;���n�^����
8�J�-�8�u�g�sO�BJBJ~�z�3:�_j����wY=�"��u{����φg>��R����v����k仗@5[UM���o]I7������}��DqS"���Z��΀�O�%)@	(����W�4k�NmUk����s����J�΍���ә�f7�����O��oUd�Y��T��콕�q��6�LG���07p�b�̸٠������BEr�\�*�y�J;���6b�`��2�ͻA
qk�ќs���ɸ	и�t}��R����.����� ūͪ��y������ǳ�q�J@Ij黅6�3�&�ɣkSTh:�d6;Y�v�&5��m;mQ�](\ZbEU�Lj~m%i)�>fp�N�7��P�x.*�^����M�J>IJJb:��8���(;�}�o/��}/mz:��k�e���/ej��|��ꯕ�خ}k>NJRRlp&�}U���;nN��)������}���u����r;�%:�9�CýV����u�ܹ��9�5ֵH�+%?%	+� ��1���f���?d|L�~q��� IQ�ٵg��uV��ޖ�ӝϕ���Z�����]wbz��j���M:���u�0F��=�r�F�v�k.����/Q����YKH$Z�T(�E���ٌ��XpṚ���sM,j�6�J�s6�w2�p�0��vcv�!Mj��C`���<���)�-�Gim��&Y��[��h��q��kW���=���Jl��m�J�C-�5��A�6����e�heA]ꋚB�t���f���UM(8!���V`#��B�d��b嘖����K	�li��$6*Q�a���=��	Y�ݓ����ԍ��p��
*q6u�@cM*�(5LR`-�T�'7���o-ݟ�����r�"�'s[\r����^ 2�w�J~	@	)�Z�7��TI[��7s]����1�
xy]��ֻ��s�Iqл��]��#�|r���wH	@IO�%�9�37�Y��Q��ݕ�P��N�����BPR���3'�&iцk����9g�(5^�ӧ�<؍�mݮ1tt.�7�� % $�$�%��5�Q�ʉTK�A��D�����k��ﻺ~IO�|�l�S��`�v�M�E� h[̠���M���b"�j36�X�t�KD�2d�y��~]$�䔼��v��g��i����C����25��<A�t(��nhۡ@�[�$u{�P����G�[qZ�ؐsӦ�C��̔�;*�]y\Ni�b������>��!����xL�.�����yn�-�2n�����>����Ev�k���=M����w�� �� 6҈�W{D/���@⏤����n��I��-^��L�g,����e�ܚ���'��[s�7"A��'�"�����d� �{�
���W��;�o�=��J!g�G��0��~��.�3Ԉ �y2;���Kp��
�3����dJپ���d����{�ϼ+徟�wH���?��g�w�����o�:b���3D�[���Y�h7	�ee�n�X�����+�ʥ�n��}�~�䦁ߤQn$�[sHh���:�</�o&������"P�){� ﶅ'4-Ȓu@�ۚzieyϽf�]1�o=U�΅{</Uw��{հ�B�,���;�~��
���5#���@��8� ��Wŷ5�7"��{��&ss"̬y$�W�v�b�D��!��R_eYx����X��'��Q�z��9�Z��վ�o0t�v
j���t��Z)�v��NY�Uq�2�L�Y2���߅[鯈#�D�۪���WŸ�=>8u��33����8����4���{�����ɡ�H�>����=i�gڪ���mKk� �r$��W͹�r$qr����C�-����{հ�B�,�N�� ��
��A-����ߥ����?:�$�z�+l̤nd+�&���� 63��:�4��0��@Se�j��͠�ߐg�� � �m�^�~���!�Y����C�_��w�ys@�3�$��?6�in$Am����/{j�������̉�SZ7�U	��ʹ��_	�G7?%w��8}��{��`��zh��y_n��j��S�e�r�	N�U�ao,�V�|Ai����d6����e�{it	��@��_Cr(m8�ދ�@�_���M���䛯����6�]C꧵9e"�zp�.��D������on�n��-ު���Kb��w.�7��E����\����WŸ�~m��t(��=[�u����ɮGЋ�r��<��Nx%�<� �=ξm΂nFwz�zT7��j�6�U��!E�m�A���ܶ��fi5:]	Xl�l7Vٮl�|�/��~�4#�����W�6�P���'��}�[�+|�<� �5��>��r�G�O�[s@��}@��	��-c_��^8�;����D��q�~��5����5�<女�D�Co����z�ו}����蟈 '?Wͺq����mؠi��Q���{j�\yVȝ�\�x�@�>�E�?Sr$ۡB��1٫�Ue=���A��{�_W͹��Ͻ�}�[�+|�<A:�hO��q�b�H%{�D6���H-�[s�]}��)M! OH�k�7^�VEb�o/�]�+��MGt�6��mз*nFz'ޫ��Fĕ�K���UeP�t6�L�������z�J��9��K/���:mX��*V;��Ԡָ�ȕ���(N�H:u�IŶ�<���,b�iV�i�͍̈́��M��r9����&�F�U�!(�Y�"�f���ٺ�bP4	M!�"X�fr�,JZF�Tݥ��
�	�sr�d9Θ��CB0�dle�X��6ZZ-���m1K0�cr٘FTø��3���1^5�K�k]uآb�F@�  �n[u�hG��<-�+X���h\�PW����=���z�<~~{�Ϧ)Z�X���Y+hv���f�Z������V�*�KS]uT���� y��a	���<[� ����O�#�w/��ʶFW���(W	�7F��@���hWǓ��H!�T�?xn��&v;M�O0��?P\�Wo�ȟ{����jqydx�d�_4�P��;y�\O'��a���_st(�� ��\�dǽ�c��[-,��"q��K�x�O�;�O�6�WŷB�q�vn�c������ �?P��Iܭ��P��N�<�dep\�(|�O�C~��ЍU���N�Az@i�Kn~��I���S��#ڽ��.����,� AmMZu�q�ۗ�tƿ)���^��h����5�!��ֻ�2���sZ�,���Yh�g�ʗV�����{�1	���Qm��Ȥi�ם����Y�r����ޣ��!Y��&��H!�B�!�B�n'�Ķ�%�:���
�kݍ�9~ؠЌFlE�nQ̤g�-t�n��k��Y���Y�����tCUY��Ç7}ty��.��:�A���[��P�wSr�?P'����|۞�wQ��>����Iޯ���D�H!�U�mИ��5L������C��̧uI�N?,��ښ �ӡE��	m�|Cn��p�]E��]�4U�
�4AnD�6�iz�ӗ4����.^�~7��#�^�175�*�BZ�}_�:q'����_7�n}�һ=Ψr��w^sr�?W�P$}�@����B�
�b�}A����Eh����ԩKՖ"���,����c�neͱ0���0�#~G��{�>4/�H!�B�-���\ϼ�W]R�YO���.�}x���G>�@�� �ۚ!�B�-���W��Q��jT�b���� �9i��K���jn<&��oxP?�M{��3������H̡@ۉ ��� ��P-ĐAm�}>�=+s�D^R~�ٔ��5zᆫ`����VS����y�P|p�Ɇ�7��bd[��bnY��K�,1�so0��z]��٧ ʣ�G��m��TQ4Yq���˚��k�+��%�4t[A:�}����N�sk�ձ���[/[,�ws�����y��J��#:�pˑ'��E�xUD߫�T�GtGs�=��gQ��N��U�nV������[X��u$�y�b��gm;����.:7�EH������춦n��/������ݧ,��L%��Fm>��ʙׂ'Bm�`18#y�{V[��d�E�u��Y=�h��5y�o^���u�Tȉq�w�{��T��[2�\2ڧҘ:�e]��q��n�ۘK��+��DV6j��3/ih�9GY�6���<=��+J�$e��5�+���1p�Gj��ZBJK�n��2GX}ƃ*�j�F_f�_1�cS���_J��R�(A���!I|n����2�/�ue;.E�yw�"��8=�y���RK��7-[쥗�G w�ܔ�l����k���D���f[�2�;%ЁmVp�ݗ6�p�y����	�<0U}n&�j�f���b���,s[{z���3l4�h ��5�{��X|��MK���{YBԷZNac�Dv*ѓ�Pb���f2�#�z]V�^��˾V��h�WT��[ٗ ���4#]���uɒf����4�y��o����w]�d�����Vn˕��k�u��e�N�;%���W�jQ��j&n�,'��;�,EN#0\�leMbl�TT�nlZ"D�#cDFah@	3cEݹ�����F-I3HI�@j,P�32)(�VL��2PI��+h�ʒ�b2Z�0ʌ�4d�i��0�Y�5�I+! �e6b�Q4Q�X�6�EJi �aI�r��F �A�Cgw	��LTd�X��(���DZI� ��E��)4bC&0�m�X�(�"`���c2����"�3�2�l�.�E2i6ɐ�D�)
 �B���H�Ĉ�)5��v腏�?I��kuA7�]�s6r�9��}�E�?W����~�zϷ�����$�uWŷCپ1}瞅]U������?jɢ2���ǠY��;�=ｱ��������ۡ@���h�C�q�L{"i�mz��������@�s=4A��@m�͹�ʑŻ�^�7�ƚ��B��H0�;gfR[	�XóDfԌ�����=[E6�V��c�\ A<�� ���q �[r���P�y-_��ѻ�ȑ3��^o/r����_t� � 6�
�ۚ �/D���C !^W����B������:��Yo�c���Փ@�t+��{�SuSY��'�鯈�z�|� O��B�m�|AnD�(1�"�t�[�*�]m���-�Wמ� �H��m��t(�Hט�k��;�zk����q�~�5��t��_eu/-��w���� I��a����(�#M�9�л�&,�K�d�u�b�Zq�r�\�����Z.Y�mSu����q�UYge������,��o3|>��� ��o[sD7Hm���ɼ�^�d��1�~�G��N��~{ ��&� 6�����5�-=v"�mB�kO����4aT��m��1�H`�\\�Z!f4���G�X�M(�M��yb����� �w&!�+t��o���zkf.�w���\�pT_����#��+�܊��Knh�m�	��Ii� �D����-�L���ryym������A��>-��+D?v��%?.���܉!�_WŷA+=7[�B�Ƈ�5=�7��e�?5JY?PmТ�H �ۚ!�B��O��pׅB�H�A�
W��nD��ܤ��+��T���nw��禁�}����W��m
��Ƞ[� �����
-��{6��cg;�}��O��)~��s��nh��o?P'} O��(�� ��v���/�;u�E��MI��Aӛ ���:c��ͭ�s�t�m0u�K�^K���hw�ƶ��|���%af[�*�7P���Zv���դt؏^a������S�X-r�ת6ѵ�c0׫*ƖǍ�-s�U�f�[[�LM�d-d���&`��-���K�{Z�.����0�s���܆S;l�X̦3�s]YD[`�en*�ڍ� ���]`�6<i�z����m.�fS=�A�ڸ͎�����L ��5k��^��Ғ�QeH,oRi �l��ֺ��0o�!��.lzˤf���,��F�y�FͲ:�9؍�F�s�(���1�MI�.2�[6�V��O�������C���6����"���:^��=��/)�\x��S!՝�[�\K��/b�R �7?6�in�ɬ���3�O���4A��������7T��m��o=4�O�6��t٨��x���P>�	�zh�t+��}%�::����,]��&�'��[sF���}�� �G��P-���r$ۡCB��M�T}s;
��O��D���
���
��y�/a��'�/)�\x~*�����=��|o�$�}4Cn�p$Cn�ۛ����}��IA�Q�ＤO�����&g�r�;����
����|�D�u�|~m��m~vg�||����������Y��@ZK�!��hCe1����n��e��q�\�Gb����}_� �zh���W��|A�����yOM�{V�M��o?P��=����` Fw�P˦���H!�T	m�|EK��2}�E ����n]�L��?k��5��u���>��WoD�#6�)�\�m��U��>�|�<�&ĩ�y�[��TUF
�����*�)P]]\]���~������_v�y�/a��Լ��q�?jk�r(��eT�(fР|�k�=�B��A�n~����h�N'~WU}�KED�w�=@�y�A]"A���n��}71ණW�����:��$[sKt��zo�ڶ�n/�y�W��G��#^[�Q}劫�~/�_����m�[�?ۻڄ�u<Ƭ���t+�b��R��i�͹~��g�mТ�}#�۝�t�q �3����fܼ[�Ō"�2��
������㘕�[+���
��PX�9;�$ϧ����ȑKRt��b{��'q^�F�W:�4`�(�
r$�.��6���%�4ܫ��ײnp�}� ~�4�wG���}y�3w>��	�@����>�.�b�{��:�_��H#�(P �h�܉!�_
���.�%�����4���`'�J���ܢ,pW�� _e֑�Y\����'�O2�FiG�ٮ��͟<D��"̓�Z�QQ��/jr�&s�j_�Ǐ��hCn�n0Knh��P�${&|S+���7Z�@󟩹�';�g�����@�{�@�����X����
���-ĐAm�|m����n7Ԍl���8�t�5z3�'��ڲ&n��y��7�A~�@����<=�ǽxz�[���ub�@ʥ��fc�1I�LQ��f��7FV�'m ��ٽ������C��4n���n�o��R��mμ�~�"D��3nJ�� -���Im��0Ou�1��K#o�į �50A]"~�I9Y�1=>�N�W�ozh]"A�s(�y���9�۱�[鯈-�q$ۜ�ܪ{$N�1d�߯�lL�φ��M����+�ۚ��}C\ԟ�z ���Ul����#�ꯈmЯ��^p���̷�C��� ��M3ݣܽ�6M��������zN�#�Y�Iv���&��^��"�l��h�܊�]�P&������_v.�mI��"/0��nv��<ƤCf���<mD�:�hۯ���H!�"�mϩZG�z������b}j��w�(:�]��{�_WH�t+�܉�����{��̸``��EV���56].�!h���O'�kY1�LLEO�g��O��#zE�~ ���CF��ο-B&�<7��oF��~��`]��z�?�5�_ot�!���P%�4F	ۋ�*��h�c�W��|B�]�^jn߇��Sڅ�q��o&�!7_7
�S螛�u�sDj�>�!�B�-���Ț�}4z팬�TD�e�(^��?��ë�@�oz~��@m��ۡ_�HL����Rq*l���(�	m�!��{ݗ]~Z���x>~�~7��}r=N��sхl��;���@�9ȐCn�۟���޿P%��]w����{=ܶ�g���u���ǁ��� ������mϰef����Ìމ�f>󚶩��/�fgQ鲪u\�Z�%�Y�$���0��nH���p\����T�M�����9ZF�����4 ��U�Ule�Y�H��Q	���b�Q�K�6�n��B]��5cE!�%��p$��0]!5�����A��F浹,�Z3"��������p4��K�f,љ�����B[*�Dv,�qjV��V˵��ĩ�@l��Mz��b�L�3C��M���MF`�S-t����	L�5k���IwVWc\0���e��Y4��>����ʤs
ܓL�^y�F�j��Te�	�-��ºˠ��^6��t����H;�P�ۚ �"~�ԩ�/�O{�f\�t�����0ȅX,�N�$ou
�����> ���#b�s;�{}�U��_��$�sA�н�w���ǃ���'�A�u
-�/c�}��Da���j#�ڠ~��Cr'�s� ۡQ�.����e������L.N<A<� ���@�H%�4m�����} owW�� �܊�J��|*}�K�sç�+�ޟ�}�H����<���`�ݡ_��
-���A�q�~�^hh1Y5�˼�2���A���}�=�@�A��(��Mȯ(��ˉ�ﲾ��t^5jj���.�+S���u)�S9S�$C��k�[CA���o�@����mЮ�K}v����j!y8�!������3?p�m
�������n����+ӳ��W�'QZ͚��;_�lG��]{�0wި��[�?�����3��rھ��u��㏳rt��)<Sn��ȩ�QwL9�k�!�	�ԩ�{z�Ku]�޹�]"Hm�׼�y5�>����Ӵ(�>�>�#��Q�ۘ�Rw�plo�o�#z�AM�x>�
�~�${��ۚ �� �܎Kܮ<���ڞ��ޑ$>w_6�.�u�/����q���h~��u��lчj%�B���Kz(�-���9=�
��24O�����=��~�J�<:�G���]"@#������_��7k�6M*N�T�&�fj��x9�e�U�CQ��ښl��r��m��ƐA��.�E�����A5��ʮ� ���>�A}T�s����F�oV@��?_�I��_�	!)�AIM��:�-��������=�Q���*�͝����M@mР[�o��B�74Z����@�Cn~mΐ[�шρ�Լ^/=�v��z-�N�5�c�A<ĥh��eQ�Fk>�֕ᛷ����]������7}����U7&t�zDb(��6��e��K�EE1������޹��+�O�6�mȠ[��6�7�y�?,��} ��Z�;ڧ~A
�<w��M��DrQqQ�*
����d� �H�r(�����t���W�'r�G��j�'��Ά�rq��V��B�n$~-��>�����tD� ���C3l�Y�\���!]�\ڔnHu���\�۬���xB�w�H �>�E�?Sr&��f��O�QU,xwg�uV�
Dc�z�{�l�!��_�
��A-����ӷE�n�ǭT�����t�G_�_�jk���6|w�~�<�F�̍.���� ��H-ڠGǟMCr$۪�����v��7Z���c����y���S���m����[sD6�P�I>�U�� e�}�Ӥ�OպӅ�<=�P�X���
�x�!�t��r z7����I��3��UW�Iݩ�7٫8�{\[ͤ��覒�2v�i�M��U�bn���-!89�.�����D�ўZꯈ��Qn$�s@�n����r(�u1�5��ӯ^��y&l�>�
ߠH ��
-��AnGtU��g�����矷ݰo�%E�fa�ird�4�(��D3�[v�lѶ;�o�q���y柏�|�'ށ$6�W͹=>GW��x۝���y���Xk7 �׃�&3�'��=?{|��р�nh��
��	_��+��ڒe}���?w�OպӅ�8{�������}@��?R�Cm�2qX�|{����$�y�� ��
-Ă	mʍ�[�5�/�A����٪�-���9�$<�E|[sD܉���}C���s��}�~]�$��P��n�z|��3~�;q�q��y4G]�z�X��*z�=�_� �h�܊�~mТۗ��di���1ղ$j��kxxz�S�s�������H�u_�������r�I�����]����7(X�S_4R8�jV�"�ABT��}�y���j��*��ݮ�2��5֝d37ow����8{;�Û�o�����vgm�0rf˔��eM����΢s9��/`ėq�!��}]t�.�YU�������@�+\�D|��I�rۃgR}f�z�.����-]:�S[�}�_kwu��BNDv3����*[ُ��}�6��u��J�<�dn^�h�/>.F�X��8�8�c�e&T�Csn�)NT �Zs��$lf�
��\����j�d�	�����R��BF���n�6js
�e[��yTbiҁ��˄�lb�U��%�`����ܒ�2��-r�U9]T�f��\�F�`۰�n�5)���+w�LT3]y��/ܔuȋ�uJM�z��"�k�+%oG6��/ޝu����q�{�-o9�o�u�՘�K�Kn�l4�f�]Q�z� n�3�W�H�0�0k�,*�v��$M��s6�w��2�bb�����:�Pʟu����1�-�ȆBuS��{q�N6۔g��p[W��B�;V�n��B�r�����<H�l�Ӊ��g�[��N�6q��(mV�B�7�^-�ùǫP��ݻ����g3!y4�*Q#�#b�:m\5�e���Jm�qp����z��a��2\
��D��lRW1aaw����#i�gD���s�]P��V�/+5��̹�m���w����5[�W�{��޾�����w�kǍr���n �3�'jb;���ѫ�]ަ�T/n�A1�|���:���ʩ���	��ь]����G�H2�E�ABll�54 ͣDTS!(Ԙ�b�'��R��c3I(!#0�DTF4AR�э+I�6f�+�@TVE h�bH��d�hB���bD5	� 1!m Q5ʸ�$��X�u�H��QX��F
RѴ$��&�0I`đ��h�*�Q��Ec1��	�sn�T�
+2(J �F6IKFLlAF�ш
I�X�M)D����Phƈh�L��
M&�[~���=�� ���]uJ6Ppd1����&�#���&�"�pPWI�K�.&e�l��Y�r���� ����-yfi֒�T&{b�dt����Z��[�2j��v�L�,رx���Mp�7V�n�ssv��0�mنZC8�m�ka�(�0�!�9[(���3��c$Ɛ(���s�.�-���\����eV]��j�,��Sc=Z�!��Z*d�uJ�)��D��y�� H���qF!1�f���Qˈ�lK
�l,R������n�JM�v�"6�˰+l�����k��%�5��[+a����8m���H�n 5]]��1�B�D!�Ytʵ
�i���᣶��F�»�A�--��/,&�����GdU�D�n&����T�,Ú�.n�X:�e!+t��Z]�3$
���7h�ʱ�M.�th��fFR�UtѰ��1�����e��\��P�#)�M�YkcJisU5G��]mr5��n]b��Z�YK�o�`���Xe� (�qR�1X�6�(v	V!qi\�(���h��T6����Bk�D�A�h�ܑ�6��1�͔�jWs�H��(��]�:�d�ЋA�T+�a3a�X�l��w,��L2�bM;���sM��ǚ�1i�kupg3dHː��&D���,6��0h
���Z��u,ئ��4W]qRǞA����f��P���rF��`J՚��m԰��d���M�릶ƭ��ȩa��sUЖ�hCQ����J��0����A.YIjj[�WgT���ݵ�:�l;Z�/.e�M�Pba��7nҤ[����Km�Z�SA	Pэ�n�īJ.[0��+�q+2��YILT����q,�����S�fie��J��5(��A�=Yn�1�/�*��6������jh.���[�.,Q�.\��h��ie�0i�΁3I��.	aH1��3#n�kw[�ʉ�F. --��� ;c�ffٲ⮦�])�&�]��M-��Y`1��:�%�]3��:�6�5k��].8�f����Z�ΥLjSgX�t,i��a���	�����[)b������2R� [�Ɩւ��n�&��p�cX�F���^e&����)^�
�n�m0��^������9xaR��c�+2��<sXu�]5�(�R� ��&\�p;���2�fC����b튩�njгV���2�Ղ�P]7����<]�U�Ė���/^��P�ߨP-Đ~-�Ka���{UX=�""�>�P���^蕟n)�A{_wt���@��0Ow&�;�o�C]�~�MO���P�y^F���v�ʋ����Mͺ�-�zo=�/ ���#9P�~<�I�_6��nEN�M����ud���<t������x�t�6�-����z���;&j�d�A΅�I���l=��\��ǼP���G�t	#�퓊��k���p�� �;�$��(ۚ�O�6�J�����=�AK�Ǜ=퇔���7{���n�|[���ǭ(�^-���T�I>�c�Zmq�Fj"ڎ#5�	Wd�#e��$!#Z�CJ��������|����#���L~nD֭-�9������߇Wz�����uF���jR�k�<��!�B�-��[sD;��!r
�z"��R���Mo�����ؘF[���z�xC�N�q:���GՙV������=�.�滹f��ƺ�bh��M
j�'�܏~}鯒�{��ʭ��x�~��� �wP�۔$���N�)=�	�9��ȐCn~��t�C�h�T��47ݰ������� ��~�ۡ_�A��4Cn�J^-q��~�F�C���D��Z��y�ëm�����x���B(�%���ꯏ��_7?���t(�$�2����ǽ��M�C��]V��:����q���>}B�-���7#8�������$��=�h�\�=�nU�c;j�fl�^4,Jh<%]�[��5Vʊ�jxl܄�t�_.�$6�����<�iW[p��y��Wg�iϲ.�w��s���
��͹����n�W�Ӵ��^�ٜoxx����M&�m���U��u���@�x���I����J���g��B�͉ ��zk�r�~��G5~��eƿ]��W7z�<v��3i���q@��י���ܭ��)[U|nV�,�Z̽��Ue3��ZF����|2G}�����7�*��ǻ�B�����ܽ@�n�>�@����I������W��M=�O�+�t(Gg�x7��{r��|�x��X�욅�����:/�����>�6�P?�	mТ���ǁ����8=�/�ah��Q���u���@��5�.� ���M���P�{»�_q�wD������Մ��԰�̀c6���3MF�RlA��J��t��e����o�X�^D�KnR�7���w�<������:�؁�o�P-��AnD�u�nh�ëë�"�Я�~�}������7j��\�Q�A+�����n�Yv�!�����@�{�I��
�4-���>�"�}&�!��?i�y�L�b�wY�ݞ�A�S_��۟�6�Qn$�鿉�������QN>�[sIk���e�a�0j�?}@�p[G�LG@�3^���1q���FOE<8��yj�*I�mGtQ���[��%ש
?f���Oƶ�2�j��N]%�"��n�ܠp!�T	m�|?7"@!�0������P;���J��K7�G� �s�N��I�ۜУ�|�ϲ�������f�̥�G����5��1�a�$)�(�Z���Ȏ>K����,�������� �"i&��{}*+�	���羡����漷�͐B����WŷB�q$ZsD]�z߽y�^T6�x�D�>Ni&���yCk�s���6�	�B�ns�����[��������=ޚ ��I���n����v-��˨��M*��,l�5��S�����P-ĐAm�|Cn�ڽ��2�s "ݪ�ϧ��ej�<�w«�%5��;�o��u^�F��r^��j�xP!�_W��P��I�� ��|�n��{�]{nUM8�z���r�uHͯ�`�x.~6�O�wt��5���������'�1^=O��
w�ۈ��۳�d)!eP���o�˪%msQɞ�(VZ�/ª܈�!��y�c��������e*b�����ÿ2ph[K�5
L�ф�ګlf�Miu����"$��
hԬ�#�CK�p&�"5,�lU�i�lꮺ�K)��. �艆�e����[���{h��;E��nni� ���ƺ�XE4K51�c]m���nPYum��4��k�h$3.�/mf`��m�! �K�0Z�H�� ��X�`a�\�]eф�sc1$��&��O��Ov��i(�a��pQ��ن5Sr��65	����b�!0n1���|����'�H!�U�mЯ���|;��Uw*Xٿ5O����so�~��P��D��nh��@��	!������g��\+�}�4?���o�7��-�k!p�^�7�h�����@����/�
��EtH �}4A����~m�O���F{:�&�͡{(&�����}n�;�E��_�I�b�{}},Ft������"�v�gý�򻹔�E��� ��Oӯ�I鿻����D6���A%�"�m�X�܎�Ff���9z�y����p���ڼ(oT��$��WŷAk�*��<8�B�`*�D6J(&٪&�M� �l�� ʹ ۊS'�o-��.�]��]e������}��s<������4��~�=B��W���\�sovܺ�*� �wP��o�@���
�����7���G5Rw̛�%*�`��"��Զ�V=��Z�����)ڙy�mƓBb�
��辮��E�֦�/6���`o5em�v�<G��_�B�{}�ý��+���E�\x�Sʢ#S�E�;�Wi�O�tnjh��?{�a��|۝��r=x�ޞ]�T�k�l"���h��v�Wתk�r$��WŷB�q$O`��/�Þ�K��_�����.}�T�^��=B&�.~���?w��O����͏��-Ȑm�-��r$�޼�=�v߈��)���}�J�%0r�\x��O�u�q��nW�;�j5��%�TتJM���ڦ[֑�F�\���@�nt��b�s_��������By���nt������6<}���%�j��)G��㌃�\��r$�t�@6�����4�kjq{��A�D�A��-�W�܋�Q�D���	��9u
-�p�����j��
`��Rs�|܉!�B�!�B�v!�����!}����y�rB�33�����A�����+l�ȈKb���x1k
�R�!X�UO��:�U�'74m����*��j��y-]�&_5 �Sɢ
N�|q�ۚ6�F[]*�Og�}:Aȑ[��7�=�tV�%�@�Jh���]�K���1����S���in$Am�n�n8o�f<V@�� �T���>�p�{L��7���6�H#��`�r���3���Oi1_&�dctr�فk��Vh���!1aSP4�\ࢌմڵ@��[�gy0?o�Dws��w0�=�����w�sI�����v���������G�$�s@��@��I����Ys��1����
��k�G}<vq7%,��{�iO��I�W������(�'{��!�"�q$�nH���TYv#����x�t��<B&���	 �:nh�� ��
3��������;�|[t{��>��7��/��|A)��!�!��ɺ�ީT�ʻ�e�ZT���k�n�������w�f�c�)=� H#HW
��Ż�U�U�-�
�k$�:�&<<dI{�D6�-��r(ܩ7�>�sor%
�#�9�����grR�k��Қ �H�����n����1�s8����������ΰ�3#l&�i���6Xv�#b�A�F��.�a��
�b�6����|��}��+��} ��Y�}��u{L��17������O�k'!��}�� ��6����Ȓu@�[sD1}�vFȆ��b�p��e
����9�������w4�9|�xJy4!'_7���}1G��m�}� �u�ntnGf�Q���W9I���,�\�@�jhB����7"�q$*�t��.�ʝ#���^s �r�����:����o�?�� EQa��t�w&F���
��MȒle5SL����
��Ǽs}�t�ȿ5��ɠAIТ�}?������꽟B���ب�̉T:�C:�n	{���j�U\�rj�����0��L��
�L����HPw^M�,Cϯg�{o�4����P,'F��@�����k����H$��l-��.+`h0�]uxA,H�xY�l���P�7	�XV��0L�j͍M��d
�\eͰ�Lۘ�1�q���
1�8[m\�"�u���.��f!��a��h���dcPc����RR�䶵iu�u�%ĥ��v�X�ohY��ItrgB�К-.�͂,v����ѽT�B6���C��|��6�Wq�c �uI��jfX�ЈR
�bݭY����_����y��?u
����nG�s��d{�U6�J�>~3s���>������|G�	!�?PmРq ��m� A���4%����o� �zh���9���N�������W��H �:�m��#o���e"X�R'�+ʨW�4Cp$��|+��n�Q�o�]Ǽ����C{g]M&.瓏��og���Qn m�|Cn�l+���bs��D�P�|�5���OZ������U&�~��	������^c=���2�?.}B�q?Knh�ۡ_�j��>���A|al���'�O���ױ^���M�<��ۚ ��r��;EI��;��1Q(��4�`Qm��@�^ ���	ix���sw�^� �	*�JA���}8�kP����5{b���m^S�9�Z�Q}Im�͹�n �]�3�H����Ws�ɔ��kŷ���xs�e��b�e��GJk �8�yFo����7�r���u*\��)�=$�.��� �l�\�O�r��ez�)[rV߇s𯭩�zwȸ�΂��Mm
�H ��hCn��H?6�wp4`ڧ�\�ߣ۰3,�e�غ�\��m@�ϝ
-���r'�t� ��鹯�#�����_6�P��o�ޜ�ﲪ����>�/������ԉ�ѿq$u9����n m��[s9�7ۓ���|=r'��.����G���F_���}i�B�����_6�]����}O����x�g�M��ݜ��k�!p+M5�T.�����co�ٳ&X7nu�o��� y���A�~�E��ŷ7���竳�m�������{i�5>]������(���Ȓt(ۚB�.y��R�f�5���: o{}>�W�}�X٬��q�	�sD���-�3�6�:_*��)W@�n�����g�)V뫰V�！J\vGN���Y�bu�(N�n��Q淹P�w�$oȱտ6����`2������J�ҷ��ی��;���,�]�k�G�������8)�l��7(����O���_)��qɁ�*��t7:���k���[�3qM#�����*��ޗ0gk�������;r�YX�' ����'�������n�^k�X��V4��cת��uWz��%)S��uq㛩䙰bʛ�4�z:���z�u� W�j��Vn��+^��g�)��	-<�e�w�'/ ��ݷr�Rn�-�u9`��v�[D�"�PV�*��$�VgU<����n�*�=�T�dȥP�l��,����n����`�(f�n�s�ZU6,٣1��ض��Jv��F�:�s%��*W�t|���q��ծ�|]���e�����p)�x8")��륖�*|n��ۥ!W�*��wR��S�e#5��LE+���W��z�J�k1���'O��#� �+a7x���o2�V:�53�g\ܚ镒阱VR�V�U+��6����A���U}���q��o;��=��U׭�WR�X�r}q`Xf�gN��,'�5�ԵQ����3�ޣ���2��6ѡ2�:�.�N��[3c��u��):��[ٛ���f}Oɫ��x"L�=*��o���_�]��j�sC���5_gv�	�q{L��qP�1��k��L�&"��0�t3u�Y�!UB�Ü��X�l������mG���7��0��la��P�1�Ć�cE�Ai�sS1g:w쿨rj�e�H)"
��BP�I��j �#MĄ�ѐ�%F0E�-w[d��Ѭb̋B[ h�(��ъM��&ƒ�QQE!,��ӻ�W��&HM�dѹ\�M@bۻ�K2-�cr�&Q�F��b"�� E�KAF��y��=չ�#F/7J+�1��І�V#`�NsF��2܌[�0P[�˜�ccnE�c%F�1�Ń�꼬m�-�v��ЎiKj�/���}_Zs_~^�x+�t(�HUt����D������B�tI��5|�ހ��~�E�؛~���(gb�ҤV]���9��H�u�nh[� ����Ļsۏ���_�O<�N�Mcfn_s� A��~O�P��Kn]�z����l{ٴ���Dф�̠�٬�,��I��4�Yb�kaII� 7M?�+� ��{�3���A�A}=�����Rڨ����B��I���+�ښ �ȐB]B�mȯ�q$nk�D>�[]~�So��o�w�o���G=Wݱp�;�|q@�s�_����Ӳ,�ў�#�R(y���r$���_6�go��ݓo��J���)Nۚ��ܿs�ǗO��}B�q'�������M��U�$�7�
WO�܉�vs�O��=�	�1��ˤx�s@�g;��+��p���W��iJ�۳p�)]s�n&�F����%魰��W�rj�c�}��qt4��
*p��X���ѣ��<�}_w�"�n>��nh[t(��z�y\a�c���oҲ=W�l\0�߁nG�́$r�[sD��w��(���`��)�,[�J�A̅h���f%3�k,�){"�U�.�*A��r���.�$6���.}�l��~ڿEcfn_��А7k�C��:����/l�>�I��!�"�nD�7okq}j��GWM��]����^������ޠ~+�/H�f+r�xL��}�s����A�鯈x�WŸ�-���p}���,��ھ{)����� O.��s��	!�B��q���\ܮ��� �H����A�B�{��W��{~9��s��}��鯈�߷�b�]��H?y9�r(� Kn�ۘ��g��������c{�֦n�r�)��/H<��mȺ�W���?�7��0f���B`�D����8wJv�vZ�N�ʸ�㐎]1�����P�D�����U�O0:���G��lY�Sڟv��XoM�cüF�a��J�,�F��0�/hVSZ�M���2Min�mn��+�k8��n!30msj�ix�t34#�Xhf�]Y��u��5zk!w�Y�Lq16ذ���U�i��'`�
ݨUL�Yml �ˡ�M���&��]4H����\����1D��@736�Yp]Ƙe{A���H32�h��օHE爤\�l��]I�p\Oϟ>n��G����Kilٚ]�eU�3���ttj%�-�f�����B~�4)�|�}�������dϯ�`�
-�+�C���k[7~���}4AȐCn�ۚZ��Ǖ&#VU|~��3���_�j���0��wtx�{��_]_7}ܶ���_�+����~/�O��܊��� �܂"��t�9��>��F�^뙻���@�����$��
��ۡ_�H0�lw��{�`�~�z'�A-������۟U���Qo���}� 1x���8橠A� ��P%�4-ȐCo�|�uP��9�X���i5~����aÌ�8���y���|A����������f��GD7Mm�&�N�ƨ�J�v©�5�u&خ�T��ػ%�D'�R�� ���nh�܉w}�}�����s7~�#���M�����78����"H��W���
-Ă	m�;	�ywi�S���cr.`�~00Y*�ݝ�eZj��(�C��`�)䴋��3H�S:��D�t�c�1�s�vU���y�������������zm�z��쨷�_xP �Gs�@�籇y{x���|+�R'�+�E�O��r$ۡ_�����3oo޵��V0��{�< �9��΅�����m�qn7E�b��8���@�~��N�����c�/5�U�ww�W)�/}�ۗ4�=�?K��z~�/P��I��M��n:Y��̵�A�˽�6���IvT[�q��6 ��B�-���!����0�=��ҿ*�M�)���P"�%0��r�q���At��;�6�Af��r�Щ*R�/�߿?E�+zh|��W��
;=�+�Zͯ�8�wG��s$:��G�Ul��_{ч����6�P?�I2���1{�R��4�=4Ar7u�#��Z}�湊����r�����!���ʷ�	��7]�f�
�$J~�!�"�-��A�=>1Po��9zV?��Q��0٩������	���|&f^_�-�����!-�~t�gk����A~��7�#�y��3�9��M�	vTc�/�@�s`H �u�nw��$6�P�aA��T��g�lB���?�
ο{}�ۥ��aÌ�tx�������"~��1��$K~��r4�~ ��Qm�gYp�q�^�UTOr%�h���Z}�TM_�wx
�r��"Hm�|~��)[�j��eD9��{���b�M[\5�p�]��#CL@f��i����H�P����X�?�����$'���'ϑ �ng�ޚU^}z\�(�����69���q��~P8CJ�����Bn�ۚWHK��E�W���wP����o��t��1�8q��	�sD��
-�xV�%T��_s�@�����ۑE�4AnGq��#��1��Sh�תf����w��!z�ۯ��ۡE���QR��C��)@��~]A-��������ۅ�B����<́ �т6V�w_�+ZۗFk���]
wu�˕�҄79�m���r=�[7M��`�\���.��&݋1��0��Iʣs�'-�q���@s�#�u_&�n m�]"=U��";+zc��=΅;����r��0�p�=� ��4A�|�a��w˫�Q���OG����Sy�u����*+��T\X;X�,�iS����k����?c��0>�f�'���������{}^�^�l�U5�����ZS�k_�J�k���I�U�nE|[�۟�x��5ьQ]A)�������t�~�.no�>�À'�Тە������q��@Cro>��r9�������;m6�+��p�p���{�	|���#~-ğ�sD6�P�O�|+���t� .T(������Z<���^�̴��<9��>9�h��5t��ӊ��O�fu}_��WŸ��?��6�QnǙ/��]��|i�w���Z������l�s�}@��H/�|۝ ��nG]dq�x��\d�ꘘ�f�E
�ʹ[L%m-��
��g�rT�g7��m��ޯ�,�P�d�nŸ;1W�T�����y�2f!��Cb�]�St�l�M���c���m��1�գ�.���,�(fl�\��H��%�[q)�*�ML�.:�Y���H�7E��Wk8���,�v�t�N�RV��yo��y-���aֆ-64��[�z��rK���!e:�¯f�6���w]�el�%�h�Txk�XYV�1,h���њ͈*l���{g9ڃm�4�9�D������� ]�Vga�j��5fn�j�t���(�j!�E
Fꙃ���O���n~��6�!�C'���{�]t&8��|E@�>o�Q뜟���B�>�A-���?7�3M���Pg�V�F���s@�H�֏F�<'�薖]g���	�SD�Hm����k��������
\I㯧�܍-ğ�rx���Qθ�zv|���>�.nχ>�M�	���"�-���ȒuC\��=��_{��~ג'����?6�V�{�]呙w�.~]x�4GG�cz,wW��=��?����_ۯ��	��ۡ@��������t��ȑ��>���>��ifVx.�P ����!~@wv?������A���:D6�I�Y��M�AhY��e�5���K��u�k�X]6ҔF�~)t�A�������]���^u�d��J|t�L{���T ���|}ޟ�7 6����0�ž�ކ	�n�Oi�*�`�eV3,�!e�l�ݷ���yZe9��W���U{�b��]l�o���+��u�&�ȿT�����u
o=�]�yV�\~] ����]#~-��P\�G�
�Mk�(}��6�Wŷ4A��XZ�^	^��>.�Ixz������O��O�6�-�n>=>8�~��4�:�\��b�|�H ����WUy�����*�]�Wװ$���#��,�~6�-���n�y��EO�ۅ��\z�P�}����+��חG��9�9t��a�ʿw!hx�f�? Qm*(M��6T��WdG�����Jƅ(
]1h˫G1\¿'�o�ҝp'�A�|۟���ժm�<=~�t��~�~ag�|���T��L�qG��?�r(���ۚ"���[~1����$���WyN�R�_����%\w�{H<��i��j�މ��r$׫��S���܉!�_W�6�g^b]{�u����[�T��O'Q�^o^<����1uKnί�w:�YS���ޝg��G[��r������T*.:����kV�۬�1zlN�����֒Yj�7N�.��><�k��u�q��۟�z�S�ʕ'Z�q�^P�����O�b���xߥ�-����4���� ���Y����P�q���� ��Qn5�N�ݛ���ul���:w�~�mS��x'����G.��s�܌���y����>���F5�Z\A���nv6��hG�5	�����`+6քN_��������t��x+�܊����y\U���LC�.�
���z}�pw���s�}� �p�������-J��yF�E�~N%�գ���e�-��� �S�.� ���p�P����hP7�$ۚ �����-�1<|����35�w�m��5���}�@��~����:Cp$��
���m�ߺX �� o� ��mЯ��o��븥���؇^]��{zh����*#Ǉe�p���o�ᓤ3wQ��_��_	�vQɪ�sks��6a�N�;�m[��)��՗�ŰF��7+*�.�Tb�G������鯈mРKp$ۑE�>��D�2�b�{Tdz绯�n�o�}#��)�I?�$���M�����d�eo�!�#���&*h�"(Mb�-k�ֱI�Y�3Aa5?�ת���\].����?��<��@�ޯ�� �ۚ��/S�U�յZ��o�Cf�׽+�Eߠa�P���D܉����۝�n�����uf�_��O���hY���]�nf'�yt �π �΅�o(�\h�j� ��T+�	���:!����K>�{��)*~v,ܽ�����;�hBr'�t+�ۯ���u���&#�W���ߨW��$�[sC��/S�U��v��S��H�$D߻�!��1G��C�CN�����!����.:n\xD3��Dͭk��+s� ����SS��H(�A\��		O�$�����	'�I-�[n���m�-kj��񶶭m�ŵ�km�k[V����ڵ��vց	'��	O��$�$$I(��!$܄$I?ؐ�!$�rBJ���[[V�ߍ��km�[[V�߄! BI���	'����)��Q;S���9,����������1 o�����
���!�� EQT � 
T !EJ��U  PU(
�)@�� �HUU(UJ� T(T�P

UI(*�T(�QTU
��	
 �T����%	JR)
(�E)�B�E*�*(PR�U�R"�R��*BP@�PUUJ�T| �����"��) > ��A��y 47�{ މT���C�H�3�8�� ɹ�J=9� �A�=�@=��w�P	ﾚs������ްO-�*�� �w8�w�����
�4P�ީT�� tɧ� ͠.`�p ;��� ^
 

T�T����RI	
�UPC� 0��.Z%�Ήzw��H�BUs�Wv{��ʣ��%݀9{�TE{�Ur�
�6�(�B��� ���73�K��U�.l��-*�7g��IQ�z�����TY1�nK-
���TD{�  |�P�HP�I)PUT|@�h �ݎ�A݀��J�
2��V�@ ;"QX H� d
�Q@�� p<���UwIU �Ɉ��A�Gv [��F n� 2@d h�`�
P���  <�UD(�%$�*P
�����9 7Y�2 eY �AJ� 1 V@4#A�T
�r(U���r��@P��  w� �]��gQ]�v�� r�
�ݎ�ΤH�G v�,�2@*(�)� J�J*�����/�Yj 0
��7o��yR����v 7X:U� 9`�� ���r�T@�| � y �p� c� ���7X�;�@��:E\ ;�� ��ԁ�C; >�(      ���h�)" 4�@ i�&���%*U 	�0 L=�L%$Q�b`L�b0���R	*�i�1�@ $�IHSJ        !�D�2di�d�4M#�F�OD<#5�G���c����%�RBZB0kyэ��;5�ei��$B��#�e|D�!/Y��P(  ��B�"��?���H�%��,��3���O����-#�4*���Z֭kf�5~���	!K�$J�Ć��!BYb=_�r����������bB!+� sjQ�Ķ��@0���ȁJ�ƚ���D/�щ!&�ׇ��x�P��!�l�eKwz\��٨j����Q�7x/�3E��VZ�.+*06ڽ���딶��%ee�j%�a(���p�
��vm̩�p�rL�h
�wQʌ�ܦsn��m`P����ۺX͘�5gm�8Ve%!�4b� �b�M�\���!Dù�7F���Z�ln�WilN�&�2�f��h͇6S���RͥWm�K~N73"��C	wl# ��F��`Z���r�E�P��7{���*9N���`&����f�1U�
�r�ĳ44؅cOM0���e���!^Ä��k-�@aʵT�K�\�S�m������M�S`RP�)��i���٫�(K��d��S~�h3�;q�f00N<�6��P*d�6�G��:���]��m^�4���[,'�:�	`��iJ����.^M(���vj�ړA�v���ͻ�vr���C���3{���`�k^l{��U4�ф�Q�5�9WtRKF��PFdU���VU�Y9GkZ�t���V�D��%A��vv
S���d;�l�q�>�ɣ��3n��H��jY�rE�^ČٛsV�LP���IѸ�w�đ�<Ȩd �xv��t�U�E5�<j��@m�.��h����.a��ۻUj��\
I�
��)e�8�D�2��uІ�8��#�C��^�yx7@N�ҏ%�n�hnĺ%jf=W����ܬ����)�U�����.�)��82�i�y�]_�o�#wsq7&̃hzj�]�`2i�PvpE��1o��9PB.L��J��a�n�̣.�D�[�\4,"�2�uhV�$uIN}+*\��R�)j:����X�XG-b+"�f0"�Q!�V�"�
ä��6���D*��T���1�nl�س�n���i�y�-�3-�;h�Ͳ�N���Z��JY-�yV��NB�jL�b�KRJuE�(��d��%�4���m�8�-B�����<X�*��5��L�AJʱ�n��l@�z��Q�zw,��[�l�0,t.������Z���ax��3M�;�L�jD���͉.�	b���q5XT��v#ڰ���+�q���8KTb�C�O�s3,�(���N����ڲ�fV���-�oDm:��+L�ra�s��@߄��ᚱ�H�3v;d��-�v��X�J: �z��i�)��CL��l�5��Kk!T�)1Y�4�$[�TE�
�W������v���
��.�8~C�W�D:��v��ѿ�v�e�Z1�,�M����V���V��C�d��
�gI���0l�+m��&�EZ����#��t$���]�eD��\�a$�Wn����J�C�nrq�`y)Q�$<�f�T'4`�n���#�!�0hWg2���BLE��ЬN<U�R���ɨqS
�U2h�#1��TF&0J�.�(Sg+Q���˽T�.@�rʘ��C>VVFN�ӛa+<��ѺA�gkw�YP��!,�j���ؕ�XS#׵#� B�
0F�8��3R[��9�Kr��%<�`��I�bD��-d�Sl5S�T7-KY��qm��y)��,E��7f9+�-P�r�(#Sv]�yC���b^f�Ӡ]7���+C@,�	����+��N���T�#zm�d����+'n��T5�dMTn4b�S�d-ݫYp�X� d�
�m�dz.��@�	*��5��R7,*�MQ�� �Q�v�9���߲;Y�&ݰ7,�� �nԴ�IE9�8�&�!LL]b��V!�ӕ��.�\�8��XZ��N�Y�%XTA�-F@sH����rvf���{7~e+��V
�6����Y�[4H5g�+e�9�nӣJVQ�[���[�tܚ��i�8�S�w��묹k؋��J��U�{�F���l�֖*��KrY�A���ٳL8�hS��ї������5ԧ�Y��m;�[T�)�i`Y	�t���͖���{,ң�Х�Z�eӓ,�P'x�R5o%���.Z�8i;����Zڧi�-�f�$'�9x�i9�j$��r�mR��B�h�wַp v�n+4��Q��E
N��%��,�ˍ���a�30��c��(n�z�;hl��r��l�f��fc���^�(;�H`�b�]��jG��u����5�Dgl\�ZlK%�`։`�"�%Zm� �;f��a���=���L܃/f����";a��f�xl+�=QءXw6���QT, �[D)��I�l^m��2�9�
OIU�m�]9��[�"�� c�
%��}�*Z�F@�Y5!��La0=&+����i�gv��n�k���T�����䇉�d��L���B*��sXw�.�(̭�q1v�m�˗F�������f�`����E�񇔂'`%)[q!b���u�.�,e(�`��n�I���FUJ�)��*+��okv��	"�AhM\Ee�5�����
�9��W�9����wF\Zr�%\�0`�v�^$�ⵣ+Rb �ԕ�/N��*ͥ!w��ŲRL�[�"��f�Ն�Y�D�2���Y&ܗe1W*�C�COm�$�Df�0����[����rV�+9g-b��I2�NQw剩�T���Wa���f�[�Y�gqY��ш�re!��@�6��ݘt�Fm�;p�DdKF��2S��L�"���)I�tθ镌�4��,`�~�3����a�3]1ތ���R�;[f\�Ĕ( �E`EM4J �f�bTq(�XFI�c��*��R�l�jF+I���EF*�ܰ�Y�j�D)��+s1�x�Q��5��B����;\���G+Kԩ	xe�m1�j�-�3E`ʊ�.���h�.��U��yQZ�����R�{Zb��8U�h�n\q�L)Om�چ)�bZP�Bڭ��[���³7V�ʽ`��T��J}Q�IbbZ�bRbn��I��"�K��N7��9vj�P���jJJ�La؋�q���˲Čh��^�S/��A!��[D�p]�UZ`+��ڛ���Z��������q��v`�J��#�� �n]0Q�ns+-�̳�L#���Y�XQ�aX���;�c$�+A�5e�*�,�R���薄׷���jwb�p�C"�Lѐ���l7��-���P���wRte��o��$2.��f*�2Q"��l$Ҹ����$L]����p��f�^��q��f4�'3��I�L�l�Túyd�	8d(`�ץe��ݗeG[;h�:���u��5l3&2U�.�*C�X&�X��pJ˹4�p�@�Vv��چ�&�Amʙ���PJ�ͩ���q薀����pf�61��;/äH���U���[{Z�����Gh^��˧�}b/���aYh�L�!�u.̽�-a�����U����d�t�r�vm#f�M�jE S\��'�e�K���w�3n	ou�5�Ea��ڨ���S2�"�ȺFy�T�!�(h��@�[yvunʋ2H��2�7P�n�4�2��"��/3�>���/]ժ����A���=T���6��.�J� K2���vu�R���� �͡SD�.�d�zkbӹ�!�`�$�VݛVP+Ek�e�Mʼ�"��tJ��s��y�VY�jx6Q��G�tG7-K�kR�2��Xdwte͘��%e\�Sk4Ӑ�$3��nZ ��(jv��浘6&h�o!9��I�b�5�[�l^8c�%�r��@^�a�j�x��P>Tp�CAiD��Hjk�x��\nG�̠򖪕���m��3�wwpm�u�	`�4(�eXX*�Ӊ-����D�'z��q�Mdɥ�jf���u�X�[ l���,��ό�*�Ǘ���#V�Bl5O
���=�-��Q�T�ͼ�dGI�)e�id��N���"�M�E��d�2���޼ǹ �b�Z�wA��6N$BY6��T҄���Rcb�I-j�X��70�l�rmZt2���@�[@�/ED]�1#��`�
�c[x��SF��ʂ�B�Yf�5��j�3��nQ'����j�v�5[��W5-v��2a�(L 7~L��J���kqB�*J�Y�[����\R�rLۭ�6U�:��J�ɋ4I�t���3�{E���ݨ���R�q�V
#l7�v�ٖ�^�7�i�.�*� �p;͗� �h����r�ڗ��:x),�[J�v�K�P��č?�
N��i$m��ٕ�ܺs.Տ���ЄX�B�����Z��I�X+YGoL�j]��nnE��f����{��PCP����&�9351+E5q�+�9e�)�ٹ�)�]�y�#���m	���Tiy��ђ�X�k*�Be�ҺTG��x.���`�H�BF,u�
	Z{LLaZ2�N"j�e��蚎�(6(;��Y��(�+6Jך���dD�K���@���t�;'p0ܼBMH�FV�˩EY�ʹE(���v�("�+hb�0�������CQ0"�if0�Xoczjm"Λ�4ʑ��
�d�	����p�Fk%٭v��p+lܹ7�3�V�Cxp�-��s�i�q(,��m�I�R�2B��b0Q���Le��le������6�7+M?�ԙ�1�ˠ��+��i+U)l`p�Xsd�	J��V"!�f��83��9�Wz�����u�]�2��7p� ���Ⱋv2�p*��q$\Ⱥg>�M5I��E���v�J35�0F`����:0[���j�-��yv �R� J�������5m:�ke�� �v�2��S̒� ,�M�l#Ne&��];��.���Ȣw[���Z�$�k�m�Go1��*V����Fh�V����s)���3D}.�-cF�/231<���e�X)МH�5uHT���:���TT �fӫȑ.h�T�-�XE]Xk'�r�9��PZt�2��ֈy��m�(��t�~c3r�U�]"����(�5c0��� �2��LM�2U��J�]�	.�
��y�s�����o"�o�W�{���,��ކ�$Uj�j�T�Z��-DV\y��/)�Vh�NS"^*SB�V`q%�-Y�j�9%�L�j������ؼЖ�/2�]�ِ0�\�������K	�p\ė��i�{��.���\�Z��X�maV
���&�1B���;����]m0�Q��ő�2�oS��
�m�raȑq�YTISd���Pq/*R�P%�*JM6�mm�ĮłP{x���8�Щ�Y��lؑ{n���1��
j�Q�Y���T-�'�J�WP%Q�ZǙ���T�XE��(-«�N��F�,Sr�K(���҂Ŧ5w8(n�;6�̃f콊�������k�����ee��ov��Z��7
[�.�{�\�[Z	8"AE�e嚻;J[�&[Oh�j���t���̆��L9u6��a�Ȫp��4(�iŎ��`ZsT+/,Vй�f�U5Fڹ�Ѱ����^�΀�3)k��y�F�=L��	�Ȍ���;̀��Z�i�v��i� �^m����\�i����J�����E���N�����M���f�F�@Lšh�q0�j���k�� �AP��Na��QT��Rܡpn�3�a��1c�V�WtTPAQx�d��B�i�x�H���ޖ�X��F坛�ǻ��	�3h��ݕ�nk����
h�F�&�]jӺJ���&m��Z�jy���qGn1��fb74�Lښj�77*���R��#r[��3"�TI�r%kH��fT��Q��څ�"�����aP��lU�;CY�i����BL�i�6�
ܱ[2^Ѳǃ�x��ڸ*�dQ�k&��P�a�B��0]����	]���E]�b ��FR�l(+CD�{u���Uޝ��q� �jQ�v�8�%%��.�P�ܹ��UA����I�a[/p�܀K�VU+.��l�!�k�j�-`�X��40L�m@��*V�ZjC��ugnD~��3c-����Bݼ�;�@�n��z�@�1B�X/$K3x��VgN!J���uxU+��[l��)`4�2�L�34j:u3Q,5&,P���)$5N���lHF�F��1T��[��٪�l��֡KU	cD����.�e]�q��j*�LiG�{�J
�7ZqI�3 �g��-�i�j���[*�ҝ�� ���V6��t&�~��Vn��i3++VRД���f�/#un�^�$X��Yk+.���ĩ"�!g3k0S��ש�E����B�)f�X	{��?_a����pϚ�"����ފRd���J�m�,ZoN9�*�T����n!Y�1��ݡ��-��k�3�KAY��I�Qޕ�V�ȶ��+� Lǻ��`���r��n'0Í�qly��yD���V�J��q�*D��A�b�HE�.
W��JW�¬×�V
�+�mF+��d駭V����9.���H��CC��ݡY�TT��yun�{�����
ɒ�۫�d��.mfmE�AQ���J�����&���Cv����n`70���ڵ�s9$�.ݪ���/,T�pZ����ARn��6��g�H���>��|B�ߺw!���W���������D#ʦ	�����43��  �0BmM�lZ��Z���E��5Z���*��cUhڒ��ƶ�[mѫ�h��Em�h�Ս��b��[hڱ�h�lTZ�[Z�k�j��mb�ڨ�U[EmF�lj�U�Z�حTm�ckV-kcV��Qj�[kb�j�j�UE�m��Z�U�Z��ڭbբ֪5��գm�M�X��-QcV��Zڍ���EV�Z�5�Em����Xֱm�V�Z�Z�ն�Tkm�U�m�U�kj6����Z�[Ekj6ص�lI6�lI6������{��x�����=y1��@���fq7�����nD�����7!��*BH����5e�}W�O���+9��ѣCϡ�oo6Tb1�w����5���X��ӡ5�eظ���d��5��J��	UYo��A����=�]�(ZF��S���ft֮���Qڢ���vٍfЉ�d�x���� S�ͽ�ļ��m�0�iP�_[���e�Ɗ9���u]�@�����Pu����s(b;?>�E ov�ɹ���:Nf7R��r���.9�D�h���7"۬�,���T �
$9����ߦ�n@��QQQ�HRqձV�:��!Dj��/4�&va;Sk�!�.!!�Dd7xn��O/h���kVY�uoi����or����(;��������1�2���c,���zn�!e�\�(Uoa���cf�M�z��4���RD7�2`Y.k�]��(��"��u�S�a��"��2Tj�ĵ�Eq����}�:���ݗWn�mq�ww�/F�W���SU�:UCm�ճ�7��Μ�P�ۮ&`�˰"�PΧG�z�кhA�L�ZR��4�ʭ�0@�U�a�������yu��U��Su"E����2�쑈���SJcU��0��SFq�2���+i;�nJyƆ&�	�.�(U2k��Ļko"��(�mZ�32���)D[��5Wb�1`��.���]�zz�+:�����܂��mvN�򶻢�;w�υ�����r������k�AU�:m��N��os���Su���Wx�� F���u��t,;�[ƒY�n"d�u�qq�Z�`ea}�D8��V�qh��Ԯ9�fep��ݗN<*���(᳦�`�`�Az!A��ujݫ�b0&rlM��/-.�{��J��|c�i��a�~���sw)
�*�QZ5?��r,d'���m�*'N�5\kjެ����N�T�>��9Q� �]gA][E*�2�IS�G�<a�*�֢ե��z�]����>{JGxG+�cWb��U�gAN��tjaA6�D$���y�ғ�.r�T}ֳ���M�|�G���"iެ��u�a�<$`P��^ M,�y�4�ݧ�>	�?[/M',V�,�]�ݐ�*�[������Ųc���X�4]��G� :ї�-��梡
��7p 8�)��&˩�h�ê�\ҪL⊳�(ʥ� ��ͦ�MБp\�Z�0㡒�՚n���!� �M;�>e��h]K�����cὮT.����Q6���t�Rq$d�	��$+m�����K���;l��@�
H������2�B��EB+ei�3
Qc2m�e�h(SKZw1�ز�ub6b���,*F�XK`j�AF���m<�B�[q�*0L�gM����[p'&,8w��a0�ÉS�[2�g!� �ǿd���;ɽ���'d+6��R鎤(l[���>u�P��t�F��o��^��҄�45*!�pdwA�W�v���u�V�����UI��=�A�X쉘e(;�Ѩ�_bV/u-
��L���\���<U�P���(�N��VnK,�lN�ll�Q��"q<i����ż��u�)I!Ö�1:]�#�Wٙ�m����8�Kvf�F�;�}��Blԙ
�n��WN�P�T�q�j�
�]�����ܩxM�8Q�&P°���wYv��͋�KG�,m.�5���\�m^�t��m�"墭Mޱ��d�~��ݳ��� F�f}��^��GST��X3�s\9���Щ|�;I�Z���ް�淶�c�Y]�ϭ`w��QIk���'W;�Cgf�	�}8
;� �_��4t	���1Y��{�侍l2�7��[�%˕0p�y�M�z] F��a�)(��hP�b��mUG�I�j�ٛtyи�8,U��%!�Z��Xa�r2�s>��ۆ��m\�Ap���b摠w$td�@�4lG��>�ZЎ�xI �� �[XI}�y�[��^f����x4�b�l�i���
)�G�V�lr�y�5�%c}�ْe�)n�Qaδ6��r�Y�ɺ7)�
��ܬK@ <�w�SKq3ky{��< �(vs��"X��j�KXM�Z��e,�I�����K&Gw��*y��:	�����7�G�7�枢�N�w�H��HZ�eK*�
��Ԩ�n��F�H@�v���pm/�"�kY)�}4��\�#Q(�m����Z��&j�����t��x�d�}��6 F�y��L���5�gv�q��VdwA&�jبp@BE_ �#\���͖k;�t�$_N�KIY^x#� ��ٔZWUj����� �W��Ә�R.g3���5�;"�Zc�>�ݼ�Ҷ���X�F؁Fj�� �5,�s��A��e�TL�C&���h�qJ/[�&ԣ7J��gt�c_�عh�Eܤ���Vؓ�\��>y]���o1]����k7q6�'
���#���t��t�����Y�x��)H�L��]0�Sz�ћ��Ö��H�@��Y}����Ƴ	��jv���l�CѲv�+��h
��+H��I��3+ڮ60Q��>��ʚ���>�N���$�s[\ռଊ�O�w����V`
I��F���\�'�E��7�^f�u��Q�6��Kw>t�83F]G4,�b�4.s�~���NHŧ��R��to�Ta�Q�8�9���o�]}����%ˡ����lYg1��а܆�����RɨS�W�fZq�.Θ��.����K1�bɻ��0�'Agh՜�0 p;��=?W��	zw��>ϭ�uj�݂R��#�6����OM���"Dr+%jF*��f
H�X�'#V����@��G���x�QRemr��K�ۍ�RtD�k��m�hu;�B[fq7K|6�ϡ[���{�R����%T��Y��gi�����~���V��Nr�^��C[K'i��Z�Y6d�*�	�N��/�<qB��&�{6�>�\���Ɵ+�6�Z&�iu�ϻFP�G���+3@�o`�v���b�	QPba;N�,nkr��inu��ם�D��ұg
8���0�\:��r*rd�w�eLx���\0P��.��Ku���ctQ78�jm��(��d����a��T\=ǆ\)��`�m�j��"���!]rw:�}K:���5��f�]�;�8i��E+�����p�(j[1��d{(�kB��eNfQ���I����;�&�����Y$�[���O�mm��_u�N�,oF�����k�D��w5HTL��e䙆�Y�6�(hiظ�(��}�o���O�7}ϴ�T����'Mr+��]j���7�')��	&rh]$�b��:P�ά�j���^�|g#(�ZD7n��m�^����ˬ=}�(`:�������12�����ES݄M٫�9��um�y��Z��bb���B�c��3��v��FY52���a+�(B�j����le��`���U�kH5�v����5=<e]�/ P�0üe����Rs���̺�ruv��ghW�Zՙ��3q�'�3�ڻ��T4�*Y��0�kӎ�_Y+/s7!������9{{�a`nj���$�c:���,%Ti�z�C��ձ�-����:*�.4xb#�E�D.��SR-�J��a@��\)3V��-X��58в�%:��w#�B�ufQ�N`,G�0� Tu���&��2iګ�w�]��Νk��u�L[�ͷ���-(�Q;#��2Ҽ�b�Ckn`V$���%�Q��]�5"��ڤn�sې�1�[�?�2��5h��1v��E���]ts�6���5�4�0��]r�Pn��L��n�F��.g:(�g-Hh��&��|s�]abW@��� �F���a���Cm�'ڣ�&W0@;�����k�C6W]}�P����pM���|\Zn WP��u�J}�˧�/���K7�w�m�P���X%����a��E�SAm� �Z���Sh@Hb&�8�r$��2V��N�]���{&�":f�-k5(�H��!kLh��b�ND(��P:�\"
0堳'b��^���|�wKts,�:�N:�l��1b7qr��q])U�[s<=�f���݁�{}ҳZ���]9/�[��]�Cbmd���Q�|�cq���!�
Wm����Wkq&۰�5�U���&\�5Ձ^���c5�l�z���`�QG.��־�5�S:d��J�&�Z(�w-�����t�D�]����E�pl걌ɼ`��9~5�l9tb�*�Y'+*쀍�Q.3"��5�t�B��W���8	�jG���,��0�-�R�6��!�ࠥ �!��Igh���mkB5���j��6�r2�����Q������on���N��^;ѰTU�&沜Ň�����@ё9�`���� ��Y\+[�ҹ`T��L֑-�y��R}lw7����]������lM>
6������۠��
�yk|�v��Z�9�>��㵲�Ґ�y{�.�U�l��B�Z�Ңzg*���j��l��(���C; �Y[VBy�U���X��MƦ��*��e���mW4�A��[�M Gd.ػ�ֳ]�W��Ej�����j�Vޑ��,;whP���/�\.ĩ�N����aI.�ܢ�W�]\xl�,f��>�%�v�*R�[5�
��"�XX�X.%ʴ�)�''6�L�B4*��tnLަrh�
�ͫ�]t�%NlC��:Kb���
MTNm��\e� �)8I8g�҄�<7���z�*כ0�G��]��6t=��U�[K��8]b��KH�s �5*M�Y[�(K��-�a�m6���N�B�Cp�uyh0����U�h:�����d�#{����k�y0���4yG^h���9��f��^&������}��l����*-�r�o�0Fn���x
�8�鴡U�����jWKvƴ��6��@Vn��#�>N�#��Ӽ,f`�k�(Sئd��
���!a��פ��j
�yP( v��P�sF�`]o�[8��.�|���q�a��wK�1�����|���:�os!e,֎,a�{�Lk�$B�Z�<F����𡊳���7r	bؗx_AF���aW�hӒ޴�/|��r��Y��\�՗�]$+1!�a��c���Nd50	1�-}�w1p�x �m�0B�$"�9��K��\J�)J��ɡ��DT�[�����6��Q�ú�̭���f��3�Ӊ����U��o*P[]S�N�<2�W��Ρ���И�K��Q���Ks37�tt��d|u��n�f�.�{������.(7�d�#!A���&pmt�0Vn���E�-�m|.� YN�%VG;2��������=��V
�3n��&�^�� �3[���Mn��C�U :d�1��w��u���bvU�TN�jۦ��1qRR��2��1O���E��vV�\r}WtYt1Vν��%�
�Yʐ��ې���}�v.�CjU:VV7ٮK��_���"*f��tt�7��6{W��Al�Hb��a�+�)�lY�z�UڷH�3��fr��v�_egl4S[Nr��SUZ�S	��	�z�n��Br�v&�ys[��R9F�h�$���phT䣑���NF	�7�����)��*���c����֮ۂ��1��o5�;�{|kr#��]��J�=ڏ��ѭ�v����	uׅ��Z\u;�ω4i���&�5���]0�9A�]�{���,ޗ̦%� �rv��oXu������"����#T�M�ɵED�BL�L&R:�n!R�\���HzЅ�n�-��h��9b�e��޷\8LY�(&��Y6����g^p�!b�/��1�r6�����/M��n��x��L�����ICi7OSs@�C&H�/����3�*w��̈́��N5r٦����^�]R+���z1��Pd5z��e\#.l�	SJ	USu��S	�uu��ۄs)��nF)լ��`ݜ8r�K�T�ݘlĵ!	F�ND���X$&�n��FߪQڪ٭�"�l� ��,�U`�5*h�^�Q �mZp]�b����⥜I�v3d�YJ�OP�%=�8�!aV�30�w�n��/�wn�D(xǸ�:�A��V�e����P�x�WL�X�j��_��$2R�r<O�5f�\˫��۾�o��G��������O�@N5�le�ӄݸy�N3s8T��
�66��4��	_325� ݧ�j�8(���j1�Ѐ���"&�E��W��qISy�;v��l6*X�`]n��wܯ���Ϣ�;Ѵ�����h�7��
[V�X���C�K�ц�V�Ue���>W�$����YTa>�uf��IF7����Y1V۝o�F��}� ��hp8�]���t�����v:B
Auu\�LL8�hͬ5�	�j+�]{H�IrE��4��\�N�e�r.�զ��w�XgN�	��;Y�S�q!q�f�1� E.gk�kVj�w�;�Z��Iq��ϝ� �e��	,v2d+�j3�>��iw�	t;ꚪNY�`�S���EPp�:�C4N�"�j�2�������[�[��1�'P-�3(L���:�`��ɢz��luwS�vݓ֬	w�_c:zd�}x�����J���/$!�6�o� ���Ci48f��8JP4@������,r�ΨDy��i
��x_�y6���\��KlMkX:�WYl�4���ju5eP�W^lզň!��,�t��*�m��pgX���˓�8�ZV���:16�۫4F�P�%���-�3I�Eh�C���ҳ`
aKn�h���� /���34UiWb�F�i���l1�M5�a���6��Ej�95%�f`b�Ye;PM�����h]2\3l�N�F�uM6�1	l	,�m�Ͷ%�!(9;�P�R�d�j��l��H�t!�|����0��Ű�e�M�3��,+�U�����[fζk�GAc5.n̬��٣z�U����EYK��(.Ksy�e�K�km���7��*��t4d�S������D 0Κ�� K\��MA�!L�Kn��m����̬X��j�
�Wj�5���ٔ4�KZD�jLA-�]���-ؼJqf���0���H����m7WAu���˘�m,�f2��9�Z�pe��s�[3n�0�k.*�lьW*%]�`ռ̄q��*�2$��rkS],����Z�͐HB�ًpS]G,��F���Z�t��5�`�Q5b�v�����X�C�D"]sa*g�i�`��Ȓ�������R�1hZ��M\��aD�c��R5Φ�Cmn
17]SF�m�J��.��.�Xy]2�\����H9Ys��WLq�@Ŵ�LH�	�hX�6`K2�n.`�f���]�fuy[q��	��nI��q)ZMLܫ����f\`��E��M�@�in�l�B��V�6����\.�GeL�l,�R$�]5�e7#�l�{+*Q�ǳ��m�il��o&�-����m0�1Q%6�*�<j�W&c۩.y6%Z�]4Ц��n�Y����:m@�
Jg3A�b�i ��e�1����uЈQe�3p.R4���i-&�qF3���u�b�mB�KY�n���K�	�e�--bM(@�4�J��S@�Ѧ��c��-5J�K��)F�����aCe�=���amZ5�V�)s��hV��V$]l�;��E��A���\JJL�t�#0iW(���Z�
�-0�-�̹�L��ZNZ�X����ck�х-��-4h��	�{J��1�M�vJ25+�CF۝B&�e�)Y�e�V�+H�-���,� �Ƹ�#��k�kP���*K���ǩp�Љ1��e�G]k5jb��Nٷk(fXA�h3j���n����̯[4-.%p�j�6h�A���"���,�yO.��*�4�8�X%r���0���(%�M�e`f��46I�tZц��K��Y��ѷRfg� #�G�&�a����-I��q�јsF����X1�YWV�)1��r�\�P6#hvK�	s6�iz�,��Hn\b�A�5-�����iI�Mu�GGinͼ��-�	iYr��T�V�Uvj���X/[W���"��56ַa�0-�Y�pFPvƴpsh�i.[Z�`e�b�S���	b�m͖�P6D�6��+4�XMѕ�m��p�P+e�YZ�6ci�8k�A�/5�e#t��M�\R2��n��V�1j&kN9���*����r+�oVm]����a��-� �\FJf�aڧXF����\�.0b���.M��!�IM�V�����_�7�t%Flksc+a���4��w6jZ����54���K�(�U���Ds��u���rٰ�kXL��[�U��f�[-�̣�3F�Qbd�9va8Ԅ�b�mm��h�Q���U&��ļM2����؅h�Q�� ���],���n]�d���Z�L�H�%�4� W�]�F)�e�og:�[ͩ�+,��0�P�MM2g�.+���u��� �;D��	��α&+R$��Yez�k��HL;aЂ�t`%�6���]�J�fֲ��V�� 8IK�`�flK	��]�.�+l�yO�g�]�^�H�4��eªkŕ�ٛ�ZF�i�3[q@	���K��,��n�F�Hb\��]1M�L���Y�"������^ ��\����Xj�h5��wt ,6�Q"7l�Ч26�·d��%[��M��f�J��V���l��v�h��5`�[����k�.LF6�ȥ-5@`��%�����$�W��
�ᦫ4.�F�jWXC�%44̓e�ـ�%֥�N��q]YfK�[^�e0�v�٪g916�6��kC�Ս]"�C:p8�0-�J(*K���e�ZV3��e빉j���yVy�؉�cF*ĥ+A��,q�5��4dѤ�o�\�+�jډH.���ǫ��d�K-���f�Y����l�ٴ�em&٫g�u�R�E��6m��.[JG������m�6h�2��G(f�3lX�L�ѹ��iz�-5nL!�`s��,1�mLnv�U�X�]����-ts��@F]�+��2�GJ�����%tcv4m��D!`�f�LV�Ik��.���J�M�����К�5���hf��:�.-Y�����BԸ�@�ԉ�YV�مͬv�Üi�������,��Z�e���ԚR��#aI��]��sxe��5!	��Ps�ex��r�X#s�˷f.����F͛m&ڍ�*�J	e�cb����mB�Z��*��y��!�Z�&����4n��e�H��V"���:��m�����54ҋ,�ɔ���H-l`��[f�؆홍[@"k�������SiaD8
Jl"���&�c�֑����,T��a!�ԩ,V��F��&�-�1�.s-n�����ILMX̅Y���(�����qtѬ31V�6�6�H�\(%�l4�5��P�+��f�G4Z�4���6��Y�u�U�^D\I��1v� �D+���׉��M4VZ
9�� %�-�*�Da�+c|�i��f��Rbƴ���f�g��bY��	m
b!����M�fķM3Q��h;%�����D����挥S�n���j�h�mŚ��mM-�֭h��*䅅���Y�uê�����h���� �u�5�Tm�h4ق�u�+�p������	c5B�:+t`X���0��Y����P�u:�n��\aCf�]�
GuSI�t��Q���ft$E�3����#*�i&ֺ�1�j9�\�b�PSb]e�V�`�a�������I������u�l�n�4u�\l6ed���fk���Ѝ��u͗*��G��E�b!�G�l�&ZLKj&%��W�V�7&�Fř�M�^!������*j�mTWLƭ�i�[ �ױX��e'Vb�[3�K��ɅuliS��3v!�Yl�ъ±��6gj�t�b�V��՚:Xļ�5i�B�jC�K0JE���MD��Xں�hGR3���a%*^%�f��,�Y�Kk���-�]�XGMy2��4f�D.��2$f���]�fm��f!�#�Ђ����Ŵ���2�R8"[�evJ�kD^Z[j(]֛U������SS��MlàQ�F��]�-� �%4��8��cVض��%�r��ݥæu�gg3a�5N��b�.!lim�2���,5+e�6en�h��. ��w4
�f�F��l*Tp�8�l�j���].��Yx��3��4+B�8���t�D���&�*.��CJ=��F�oeÉ�-�&D�fT0t��H��� r۬J�Y�4�5�6km��+�ֶVf��@�f��	Fk[��ء���5�ԃh7VY�fٙu�-�F]3���Eα&���WR�,�!�0��Z�Cb�%��[S3hl�]���Rk�(��W�]kZ;[)��J��3]\{e&�LJ*R]�U��rŶ�n�(S���h1��-����,��B2�F��uGB��
�Xn�Uرk)��A�ʖfD�ֵօv��E��6gع����f�2hdc�7$����f�&���+6!SG�+v�Z�\;E`�F1�V'�攮R�B=Y�/@{[�m��]YU��.�M�1�	�v�����x>Ly��hym�+S�m�d�Hl��U����%6��u��4ɸ��Y�i�4G�g:�@j[2kP�Lr�Lז�0R��,h�`qe�#Mqto:�7TæF�+k6��b]�+m��Kxf��-%.JLݥ�WZĻ��F�:�ڻCqLو��ʮZ�en&����Uf�B8���pҐ�l��"1�l���R15���-B�7\6����тR�l3.UfC]-�.����Ɨ�S_��;��4�X��#T�h�@ݎy)lwjf;CfbQ 	l�S"�-.��q�T����mu �Z3w��K�LVR�<�w�6�٦yZ3�Y)�˘:����R\gF�90]B����)L!.
Z�ef(ͻ���ݶ�a��d!�2ؓJ��-Е9l_��y�1o9�J��i���L���D�5����e���k��dA6�G@��e��v.�C�o!�B�ŚJƱ�Fq+\le�t�M�۝X!Svb 5&*⸢AR�`��cm��m��4�E���W\�"d.����fuf9���f1�n���՚�Yk*Be,j�W@]�Έ����1�sj�fC�hh��̶����V�n�"��1U�t���L��Aͅη*���,Ius`���W[��b�UJ��pf
�2��ʪ��j��U�UUUUUUUUUUUUUUUUUUUUUUA-<�#[���6�A�8�f��Jء���aݡժg ��F�.nC=�uL���e�#Ԇ��U��6�m��fp�xr��a��`Sמy|�*��,�lŖd��؁���]FQ��q1]ڛZ��3�]X\�U�}��;���d �
�d�Ǖ���]��{������%FF�[��yb��1}��Li��Qo�1��3�޼�r��k��}�u�輾7�C����F����k�@Q�ל�Fn���m��f��%h �|W6�����ywu�y������y]�ni��F�EE��Q����y��=��ܗ.��颾{��c$|g\k��wIy\ĳ"ZR���h�6��D|H�o���K�%��0��)2��j��J����l^���U�JJZs�hf�*U�a^4���ٵ��2��U�.WK(\�����)�W��lR���*#���.H�.��[v%�n���]�����	[`�r�A�R�,��3�5�h፷�0upflZm�����0l�phܶ�ɠ$���#�1���2L�4����M#(�V��[i@fc���i�涂KLM��.$lĵD׃)LD��u-��#�Gv�,u�E$ڷ%-[i�� �[]�Z&NK�V+t�)f�=R�ln���]��+MӅvѪ�e�M5rˮL$q�M(�ݡj�@�LZSk�%8�lMV��b�M����beP��m���`�[G���rR%�cqAzĖ�1��콴ܻk-(��� ɳ3��;h;�q�Y�f���J˴t�Be�ٱ��֖�,G?�
�4��o[�0�h�V�.s�Z1l�-��F�-zeІW��4%���Mcmͪ�Ł�UM&�Ƙe�i�m�&e75�j �B��j��F,�D L��]��	��2����e�JЭ&��lŉJS6����%��.�m[��f��8X�X�b��i)3e].l2lcQ�$pE*�;�!���[+�	�c�c��\y<<��MP�YYh늦�0�蚖�תE�ˬ��{B���	�	ua�]*��f%�V��@h�+�lR0��#����[ck^ʃ3X���w[c��st1�5`p�R�v�����3�[l�B�Kw$��H���m�P����IF���$��Gg�n���F��ŭ3L�����-|�Q5��,(V%T��d6k���-�#+�� ���.��ƛks�	i��YAƦԁZ��F(�"�5���\�X�̦�ѥ5���ҮQQ�]U��UUUWM�2�^n��+ݶ�Ҫ�٠,���t�G4,�B�m-jKab7�b5�1���+
��(<���:�6؂�F�ZKB*K��X­���k-�ڥ[D喀�"��[P#)�X��V�HFڴ+[h�aYV�c���6��F�(X
+��)hp��U*�Yl�TF֖Ѱk�1Q,i�jo����!���p[�cG&��
���\emi
9��e�YG;>���^���}���_�!n ���UU�Y�1u��#D+f��,0f���A��<^��6����Kq��\X<ł:�gǵF,f���y�f)4�'����������W�φ�x�� �9��"An<�
'�ب��1������s�+ҥ���@���p,���7��DW��ւ �Bڑ�y�f�GF[�����>�̉{��NX� C����H>-� ��^6�
�&7O��H �Ԝ��u�λ1I��݋�4-� ��%i�;c[cuA��"��[��ҩk-���<�`;%\�j.wh��lF�Vd@�Y��H�n!�
�������d�J���.��������D=r��כ� �[jH�[���g�%]�ߧ�:֠|�pB�.ރ�.�]\�M�>j��6��u8;��*,��h�f��u�F9���Ɵ_,��
���<+��7Ј'q�9xfm�tfv�����H'6�ۻ"N����l��y�N�A:�zwP@��"}��ET��.��ΰ�ަ��y�f-71���/H�$����A� O�a)�C�qa��&'���~!�7�ٺ����W<w9��<�{�O�\Hb�M�ۡ\�>#{�(wq)�ww4�2��ww[7�)'���*U{7�x�v������lA{�$����n�sl�̻{%\t$f����5X�X˕�c�])�q���\�fh�!L�=8'�ڤ_ ��3�7vD�����������Cwb�tE������r$�������@;�>�Z�Q��ͯSkH!�
�]�����2W�g�����A�"7uqO;f6^)U��CޡK�ܪE��C������*-�W��Ӄ�;;:����;��c`�t5:�����z�;0�����6�"����f�\f�]O*�˙�;W��:�!=���D=���^�7P@��^�{5*^��) ��v���ݑ>�$�v�ܚ}�b�sA9ؤ"s�؋v��8s$3{��#wP����ۺ�����˴���@U�N�x��z&{�;ܽ/�@���������/�8�A��b'�O��&�W��륛�4ltq[tH�1��Ỉ� f͹i����>��$��$�Gۺ�-�Yu[����w���= ��[g�^�W� N�:�{v�7vgۺ��"�ή��i�Go/H���$��s�4�"�N8�s�I;dI݋�f8�ݰ���WZ����F�Ϸu{<7P�_��w`�m�ۻʕ�C�w) �������C� E���f�B��@����Ϸ�ϷuHN�e����w/]�= �p������X;!� ��X����Zjt��*����E����
9�kC����2�;�X�9u.��(9���ө���n�OW�w �����RC���f	�$�ޡS��o:ܪw�I���S�9�wan��QB�j1?M�BaJJD�ֵ�,�+a��1���'fB���qeW\B��T�]�Fs�Mt���wuz|���]���<�(�|	�Ga����V�Y�����Jf�t�0��Wq�1���3\�Q{�ۖ(�@����k2���fwo]�<'ې���wu	�0���u�/��A;��wPDn��c�� ��w�n��;눴ӏq�A{"N�/|wuI�"G
g"�"�:��D�ȟީ �a��]gg[�ʕ�S��v���s�s�T)P�#���㝳������H��$������IfyL�y����{
{{��l�u�@��dO�� ��/��k��C���î⭝������0+F�f�"D�Ҡ4�gV���s�$j7KI��,R�Ob��'#Ў_6���-t���9VH5d���(9�11z��x͑-�u��C�҈/&0�]�R�2�kT���15��K	�F\����RjhJ!\�f
Z�PIc��H�uɚG�9�7J���;&��kL����1�yh��uq�h���� j��f1���bm^J-�L�	�u�h����iuz�u�x�i@05��X�l�rܰ�G*���ܿ
o����1tK��ȄnԱe����p�^ufX��P2�ʕ2��C��R/PDn�Ϗ�vD�̆�:��w�b� #�0�D
�"�Ss�1���)>r%����˻���)��p�b�cӖԐ}��$ػ�-����ԯJ��Ov� ������1q��\��4�㏗�u�݄'wV�;�,�;�-�9�3y�<�������ݑ'wT�wP@�ݑ"k�ffc����|�U9�?_w&I���M�Oׁ�N8����n]�2D�$$����H�ِ|w` A��ȓ������Bdt����&�=*xH �j�}ڂ#wW�n�v����`�pA^��5ݬ�6�Z��#Y��0YZ�6�7CZYAx�ʩ�a�� ���H;��%�B�;{^'��}�(q� �}�WW�=ܤ@�@n�������(ē*b�Q�qPV��Zm�u(R�54�[l�ݕ�Q�tw���$Ʃ0R��GWCE�kcy���i5�yv��o:�]�~?v�(��jyC?Xx4h��/�I�ȟ�)��ʎ���|Gs^�`��H;����E���
�"*�;6��j�c�2��� �ڂ#wg��Ỳ$�ǰYħ#+�5:�}��O��D��B۽���V������;�r���i�˾�'Ŷ��x�ݟH'wT��@nn�o�o_9e���aVud�֞���q�ؤ��dO�� A;��{��uѫw,t��Ɉ�bB��sU6�AhP�%�]Ktv̷
�6B:�,m���h�L�C�� �^�N��P�䕚�":�1��+��������=��Kʹw\��wdHv�wW�/��n���F�p�A_)Vc��[�[��ݤ#g��v�"|wu�:�|���}>�A���� F�ϧۺ�nuڨ['��j����r1	ބ�D�A�Y�$��\� �r2����3��Z΋�vT���7z<����Ͳ�V8���{��k#��#���{��L��xѾ����{>�u��^��/�Q���3P8�ϻ�` ��y�z���G�g��wW��墇P�'1�2g�s�waA��$n�;�Gc&��8sXu�c����M����H ��@��dH;��wP���ae��@����9�nf��j��.QH�M�G]E�0	��h�F��3��>����A��>;�"f�k���8�=��_z����X�Ǝj觾D�n��]�*WpH�V�;H���..p2����G�ӽsst��3�;��{P@��5�I�ʷ�w�$�B>{�An��݄}��g�J��Q����=kvU��������;��;�ݿHrԩ9K��1o�*�ϬO���6����]e;�FÎ����Iٍ���U*dU4�Y�o74Ă	p�54���x��}��cv,kU����[N�<��ϥ���}0t��sA�-�.e|"X�#��@��=�0��@��ݑ>;���K{��b�"�@l���;�1Y�B��Pǻ���\�wtRe��0nq'翉����.��f�N��(�wGH3eݢA]-��b��+�4ٷ->_� }��a_>H�wax�㻪Uy�gxv-�W�(j�/:��7t�Ȟ�4�D�۫�7P�~�N�"�2r���W���j���ٗ���%�A/�Igl�;��p�PL����S�:�gݰ�;�"|wuzwP٣���4K��DD]�=�f���\T4�w*�rH˻�I�wE�$�ΧNd�U.���>�>�/N���]���{���C���OO[�a������M!�n�˻����5z�#wr��C�$���c�&���/r�37����㏷�H �{"N����z�0�_��5�D��!Z{u1��j��M_��R��:�1=���ݑn���v$�FlJ,�Vch]���)��w5H�Tq#���v6!��虒�P��2be.&�az�Z�6��-��c�u��0�j�(���Yb�:��0e�����ݙr�Mv�æ�Pe�C�Z�H�4���ajcYr�֛!Sh[��f�U���PtҖ��m�M��D&yJ�\+��98k���[&��3��f��VX�k��$ُk���ZU��@6.7-a�,�l	`]���˫���Cb=����ϊ �:��̃B�Ĥ�,6a�-��Mۭ�GV[����bT�zA�#{��u{�̻���׼�&��a�����j\+/�y�u���3㻲$����AAsn���H�{ f�*V���OR��B6xH'�AvD���o�P��p���";�	/yIn�7v��n�9�r;�]$n�������d�8�A;�4a��N�$cww4˻�D9Y�q��8�{�nF�p(���H9�������"'���j��=
xH ��BY�n�7���.��$O���wa	����"A݋֡$N_ �s�O�n9�7ݑ�5+ݔ#g��8�P���H;������|���x���sv�VfS�ҥt��![���� �����~~M,�=�t���/���7vD��-��V]�rv��8�z�M��Nbi*�v�w���^�ܐA݀�������*b��cǡ�����X6\ž�����Yؔhޖ&5�%��g2nz/55^ԯ��'i�Y���qE�WcWfS�)P�k1I�P�f
]��}&�\@�(p=���ڂn��=v�n]Nd�ᷙ"|{c��S�7u	;��|Eq��MMk���ێ�ԯvP����� {�X;���7P@�ݑ"����r`}ڂ!�H�n��͜w|�.��v��lq�{���t�j�*��n�7u	;�wgۺ�Zi_F��N $���ie���|��K�!wy)2��c|��n
�|S���g�X��SBnYs�ft�Q%�\�`křLό)S)��A��>�3�v�'wT���u���صCݔ#g��c��:�P���4}Wr$�j��@=ېA��$v��ɓU>�Œ1�N�C}"|}��$�YǗu����Q���}����|���J��:h���^��K����P��i2��#�Ɉ׎���g?���e:ʖ(��Z�d뻑��n�cgbJ���0�`�n�C���ܭf卪��)F��NY��o��J�ȧsX����������lcӝ6��Q.���lw�}L�`]l�7�ے����R�����:Z4�1�t��pY��r9�=u}���\ؚ'cao_ש̬jӊ���9z��ő����NF(�v��<�HYa=�8�tƇ1Cq��Ko9�B�@]nr�=��@�xz�7�M�a.����{��7p�
����U���F�)�8&*���ݢrq�˯�nEd�!o:3#���\]������3��uȷ\7A�*5P�y�&�;u�Q���� �z��.��XJ�3�>��x;���c
h��K79(�4Hg�7m_:�6+�i��1�37��F�t�4�K�"��R7Sk�w����NÑ5[H`�x �g����f͵JY�/N���z%#J��WM0�p�ܮH^d5��`ª�L�����|5��@T��쏸�q��4r�G�vc.`����i���*��9k�㾳=��'xb��s���y�3�+�J�o������W*�vΚ��0��Y�v���/<��5��N��]�8 ջk"���v Z��'uTmʙ��Ή�d�v�N_�%����z��9�{��^�E�6�f�6Ŕ�%�ٳ����Իx��U�.eƎS�]v�v��Oh`kA]-�ݸSم��I�ɫ�Ś����s���:U�}vq���5�����������6�d=����w�Оm%1:�!l�:�l��W
��1o:wm�x��^��*w[��g[RJP�o���S�{׮�Ȣ�"��u^��Y�������wN�8$�)`ף�S�'��(��{�Y�˗JO6�_�����r���w��ۗ+��;��v�������A̗5�DI�������O�c�э�.n�1���u���Ę� !,���b@�l�"5�
���#d�Xh�! ͥhAk|�˞l���'y�"k¡�]�|�%2����C��Lz�u��W���Fk�%�#��Rjo%==}{(��B6x~P���D96j����w$T�
) � ��wP�wr�A�A7wg�ńt��B��ӌe��u���E��OsR<�D��^>��{6k�'�_���]H�inH�G GK�]�PSV9�r��Z�lF�V{�OG�l�翬O�>f ���7a���i[�&�E\��W1s[�ur����>>��wc��^����;��H/�x��!J�^�����E����A<�"��v�5;ӅR�[��Fu�k���"7vD��싨��TӣX&��
�w4κ�{��&7�ni1��(��ı�wr��J�<���9�!��	#��%�)n�W&�bѼ&�<P"o���T�Cӯv�ƞ�xv��R�7f�HP��ks4�9�N]yr%���U�jfz���ɽ;=�tc������H&��/N�-�����c5��)x��)�č]��2�P�����P�Ԃ8�=�[{
m�-l�o` F8Ŷ�����"����G���d��aM�9�kq�#�q��@]�v٣3E�op���������#wg��7v}sg^�W���[�;�<;M��l�c��/u	;����F�'v ��odC��p�x�jH;�!h�KK�h��(7�=��/�^#wj�;*ʜ���ϟtȐv���IwdO����AؗN�]�W_r��[� �^�����BN�n�^#wg�+�HnC�I�r�I��"|F�ȓugwd�|��[�p ���mɤ5�#���5WE=���ɤ˻���w7{"N�v�6�ݙ���Ĵ�o�8��"&�}٪|A�@�ݑ>#wM\�Ko����E��ʱ[Ө;|���I-����f_JX�;T4��/�v�)��=(*1=U��L��$&�3�9.w���q�LϏ ������������U���RiF�b��Mr�i�YKW&��6�α���&�A�ۂީee���5�`3M��Qej��&y��͛;	��B̑�--2YKLP�6ר�uS��QxJSZô��E�p�
��a�p��l-�m�Lb�4�\ۛ4�s 2:�� -ɘ݀î�*�۴i�z���K��-#2u��!������"W�~+C�u�\ۚ�b��*�hhYX�k��k�Xi�nZ~_�BC�sw�����wT����k�y؝�HF�g���N馓P:CsP�m��n^�Mn�^��WX��7nmƭ��g4^�|n/nk`)�� ���){u�����i��~��O]�U�
Ү��У2�����9ǃm{ʹ�v�CW��f�b�86�ڨ�7z����Ǝ��ll�LN�WM����M����m�7�ݹ��3gJ�x�ޛ�壞cL���s��b���n�R��J���0�+.�9XI &b1h�W2��p뮴		]5�lGPjj�,��܏��>|��h��v�ϣ�����p��j�}1�,�%�`vF�i��mέ���~[��h�M]� u�"��\t�f��y�-�}��$D�f����!�w{;�9�w/�*�X�^��OE(����N��r�n|�$��⳿o�$�1�w���L��GW��փo$��V�sq��A��oA=�Wf���쎥��y�>k����xnjn<�A��QOw�D���h%��&�ҍGjY�иA�k%z���
v��h/GV}�wV���m��W[��#^�Q�{�Npê���w�Ǟ��@7�^���Z���N���SB�c�[Xf��E8�ZbS��b�5k�)0�L��x��}m�ڵ�֭{�;5d�9��uFy
��w��+u�6�mx��{���_G2���=ٓ}�Πb�d�
�@sm�Ӷ�.Q�J�3��p��6yݣ���5켙��Ef*��MZ6�B֯���^�}\pgi2:�o{��oXXt�})���G�u��X��sO��ާǀI!"���v{�>훹����|/J�KB���0Ww(J��� ��.�P.�[���b�8��[�q4!��Aз|�)4!���@R�wW<�浹��V����thC`_y(5��+���*}ň� �4!��.P��i�h.��B]�!�+���E���Vk��h��	9OQ�L�;�="���=@c��І��%
��>܂$hWw(J��������\��8%X ���F�
���5�1����5��0v�m{ ;L������'�:N�@�w �4!Ａw e�����޾��i�kا�p .��=�r67�Dp���N�BoY�"�.ﲄ��� $h����40.�D9����y��3Q`��́Mi�����e���>�s���V����thC`_y �{�Ю�
�+2��V&&7��v�Za��^�4ĕ���!���E� F�O����{z�J�*2�߻�8t���U�� _ܼ*�܂%4+��)4!���@S@]�H4#����7u��˩mkZ��#B��w����a���5{��r�C�Bh.����[K�9�S7�)?�JL�$��t�g;���KR�{�+�F�(�8Gv��[71�C0��3ݗ11;羭Q���7�\qc��7Q����BH@�Ne��rPR`�4_`Z��(��wr�I��A4+��'z�v;#8�c�E����n9��o9��Qz�|@F�:І0/���rP�
� ��6w(�-�y{駣Qpn"&��pU[)�a������hƽ�Lf,P�JEL��#uZ��#R�4�b���k��"�+��4
� &���n���í�z�P�d:Ќ�O8�(�b,���ІkR��w� P4!���Ȁ���B0.�ASB1xq�E]�a�y;B64-8  |< s���n����%���k�<��B�^��j�t�.�PsR��v714w��7������P��]�"SB����1�� 5�m��k�D8��6*�h��z�}@F����CB9t .��!�.�P��i4#�ή����\�j�c�+�
��=�4�S��PP0Ch��	0U�8���z�P�d:4!�/��*9��6л}�%C�eC@]�#��4!�wB� ����;���@k֯�fy����֯s��JѠ��)hC�]!�]ܠ��h��m���O��~>���=�b_��y�Y���������}G*di��(enb' Z�n66�o�\'S�-�ě0dR��� I����p�pJ��iV)�h\\����帔��b�A-t���ˢd�(t�cs��{+Fl�8�uc��cb���&�-�l�B͙a�&��Y�r+�jD�����W��ָ��	].�n)�Ɋ۩��e(�\�Z�Y���R�L�f5z��2�qeQ�U�cY��d� @�ⶭ+̷P�\,^���ڲ�� �6[}��~��.�f��Tcq�@���κDr��2k��͑��Xl���OP��x�u(T4!��KB��BT���Q������Ww�ӽU��#p�sX�|�ft�dZ���@w������I�]܅&�1���RЇ�q�hx�/HE&
��AI�[� ���G]��[+u�g�c2�1�JZ�r��]܁��پ_grbЎ���P�� R��nAPЇ{��-l.�P�A��-L���V�WN����/S�UHu�4��Ї|�B)���ALƋ� ��.�B��w��zW'\�#=�.��5�J �; e4!�.�P�Y��Ù��j�V����u�ېTЈ��N[��q�pB0�ܠ)�]ܠT�]�)Me��Cwr�Q��;T��T �Gp�.s/��d:4!����P���$hWw SB�����^����yۋ�j"_%��jbjbtB��%!���كC�n�c6��.�L��D�uqF]�*hC�yHE
� ��0awr��_5����l';�� l��̺����P���e�W�AC@��F���
��B����&�����35�c;��zܾb���u���ת�1\�лl��i����Vt��y�7��9Z-eù0Y�)�g���u��� o#K���|$��ʤ�nP���N���9�3�\�5�U��70���4#W�B)4+����:�U=�"��j�C �u!LIw�
Z˻�"�
��0Ch�����d���Y��Mw�7�g�
�d:І03�J4!��hWw RhCawr .�2��N�YZ�v��X�H*hF9��!,��ܠ+��kw='��/d�su��HthCM� �4#W�oX�5;B)���PS@��F���@��wr�I��A&�wr�+���[B4�ڔy���L����:���u4!�;ːT4!��HEB��wr��q��w��e|3j!��(�E�JPE�5�)femls���óa���K55k��I?w�'�:t���5}�!0Ww(J�.��XGڴ}��ine��V����»���9�wX��'z�.�{�v��l.�P�pІ���CB1ga�6�w����й�F�kw(_3�_f���h��f����І�vHЎr�����A:�N��>v���#)���	h�24!�9ۑWr��wr��@`�1Xdﾟ�.�
�f����~�ø�д�Z��ʱMj�@�՛C�˳�9�$nЏ����pu�t�p�÷=�T���c��]�	 H��9�q39�z�����70B0;ːTЇ��!
� �І�]ܠ)0����j��;���6��YM{�i���{((`��w cn��\�޾�z�z��3!ѡ`g��ٓ��kn:�7`�4.버���%I�.����*�����w Fu��E����RnЋL1���뼸�]�cN�q���jjP.�� 	9ˤ"���A@��` /�;�w��h�숌��0bB�M%̹�5�+eI��/h�P1�i�e��N��f���J �s(\M� -
��
�]ܠ(��s�r19���;���SքcU}��\��=�k[����*CB�]!4.� ��������SBAw �hF�o�����[�^��1�J`�� Nv����^;=1z�z��5!ք4��(TЇ�� ��X��c{�ΐ����4�Z���*�hWp�!������3��c�Xzٝ��W;��p3RbK]�!�] ��w 4��SB/��w��� І܂$hZ������9��\��s�s�;�\q���hC`w�����Uyh�0��B<��߬:��tǅ�:��\7yw�]��+W�[�9^�-�s4��6�r�~�#{�3U�:z͝�H� 7���a㝔0����4�]�)Me��L��ό���Mo��4�����z���t���1Z��B��(T4!���wrB�^ E(�u��B7�ۇܐhB0�A*LJK��[%��r�e�A��;*Qq�i5z���t��d�4!�or
��3}�!4+�F�40��@Q�s���<���������hG1۹���V�F���{�B(`���%I�� $h����w"�x���{��,����@��6�J��u;�c=�z����50���CB{�!4+�E����P'Y��9r4!��� �!��!0Ww((!��� U{nEG$r��Ǝ}�#�虷U�+R�9��.�!��%4+��%C��4��#3��:7��L=rf�b�AP4!����зp�c��.b���s#�nnuX��f�:1%�� ���w��1�w3��g���m� H�w(0.�P���A
��j^v��v��-�Cgr������X�qެE��LZ�.ASBPЮ�	hC]���j^�5��Ub4�������+��Ǻ���wD�MvpmY�X��:��-��$_r��7��j�|�KV�,vs�8,cw�/0�E�;B�N��9=���۝RQ qُ)���z�`��A�G�΄����	n��&����y�*w��5m���Ǵq�g/���X���>%b�Q����KLz����qw$B���U�8Ò�@���[b�ͧ�����bft�5�%٥���(T��nJ�Z�ko
����U�횑69�n��:��j��j�2��ؔ��㈔������<���M�{�υ�c:�YX�fh�0]���R|c�S-VE���(t\!�;�P�u��$��9Z]�����@K�Xe+*�q��M���}C{��6�����e�έ�w�nu�A���������yȡ�_�;8e��oZ6$��[�6�d��\�p�өT�yf��:l�`\�g��MUdH}���*�<�Me�H��3)آ��K���:q���̧+���:�oq[EQ�]P�%�_n0�6����Q�ਬ7����,sm�r f7r��:��if�S��d_��X䜊�8�Y�Ha�@��"(lU�
�c^B��N�L�Knk�ǯ�Jcs1�u�O`����*�K"vs��WCɔ^�Q�$h�TV�M��1LF�Kwzv�:�H����mB����"��X��sl3KL7�̲�DUX7�Χ`rR��j��fB���i7��Mk'������16aq�
]0����{���y��N��w-�u�w_�	c{��/~�h�&����]vэ%���Rq,,��,�2F�S��A�s�zr@Y���
'Nz�����������y;�8#��]�ι�������G\�؈�9.r�u�s��s��'w2��`�wk���@=ۯwe=q�8[�������������ܗ|�^�a�݁�)��]Jg�w�~;�9�Ύwwd��N�b.�����w�zz���0���Q�=��	�����}��}8��6&i	��Ŏv���:�wYa`h�1��"�ݮxճFvn��B�b�:��P����YEث�s�L�:l˦j��,��mb����9B�։ mk�qME���r���9�]�Q2��1\�iC)l-a1�i��-��ce�4�ST-��7
\Gi�Q܆#ux�2F��̶�٢�J�H1�m,A��8���K��K.5��*"��B ���{Q&���͛;�u5%	WY�sw-�G&.O�4�_+�,vY�h���cH�CTsF����̇n�6�j;mk�Q��,f惗�k	eti֮�ICmd2f�I�r]&e�`i4ҏ;f�c�u�1YW+��2Bk*�-i\:�����-��Է$זm#�2!�x.��#&--�큀�t�`Y�XC[%tRJ�1R� �ܴuf�	j�@õ�M������R:��hI\f�.�q�]����^��t�j�R�\��kx�W����Ƶ�����[Y��t%�ࡋ�m�7$Mp��AC�K�h�-�A��Vi,ːͭ�#���fb6�2��ZV�]�⑳:��L�4G6F:��QPa.|f�O<d#��읅J��T��3j�W��MH;c6:�a`Dr���c�ڔ�[n��G"�31���7j\�N-f�q�[�+s���c�2����v��.��Q[���!�\���Љ�e���)�x�Ps�q2��e��{iaA{K�s-Ŕ��LFgU� ,̄�Y(����[KE�M���LV�*�E؛�0�y
����B%��p]�B�S����AjL�]J]xg�ݣh�f�kŘ{+3�^.įĦ��؆ƛ�M�87X�:�5��`�T�Qʉ��"22�K,aY�جJ�U���LLka/46�=���bY��a��Vछ[���˰тٝH�+a{m��a��Z�)U�]�UUU�"�bo�y��$t��L#������i�y:t��x'��%z��y���jǈb*��gZ�WB��3B�)��/&���R6��2��mΖĄk8��p���[�]��b챩�LE(m64���� lZ��5�\�!�3q0B��.i�.t#H�]+�����݉��р��K0*<��=��]f���*��Λ]�������K�%���4K�1: ��0�ՕW,!AR��}�����4�V7I�9�-��; Ƹ����GE�Ф\`lMb
-W�$�v�����/@%^�HE0Ww")��� '$��'��#��S��@b�!քd���9^��6�d@gP�й�H�+��w��1�wr
��T�}���M�whE&��@4!��nP��"�`��s7������B�k�
F�s�(E����|�b+|����M� ��/Y���4���PЍ� ��24!�w(S��4Ur�Z|�g:�x�/=@F�:І��.P^�B� �І�]ܠ(`w!M�y���H4�:���t�S��PR`�4]��z�j�=��Lc[�:��nC�l뒅CB,���^��w�&�1��� .�2Е�� ���"��8��ޝ\����E0�s(
3��|郇;s��cu��Hu�h5�#B�.��`��PP�+� �d�ﯿ>z�|����̡�Śd!	e��<���.B�IW[4�;h������6���C��t�q$�*M{�$hWw RhCL.�P��F�ǜw]�T���LSB95��9[�� Іc���B�����cA��)Ý6r��]_����O���pC}�3��BDݣC���۴�����#;�.�`�RɁ%rMTO����N�^�b7o)�\?=� F�P�	��|J�h߈ ��z�w�}��Lc[�:��@u�0;��K]�D����3����96�g:��@g�4%ˀR���t�Rh[�"~x��x]|����.¿�G=Nr�'� ��>ϣ��k32c�p}�W҇��o��J��izs�9v1��]E������F�2�q�L��T�Ks�C/M蜏8'^����]c��������z!l�������+db��r�aK6e�\Ժ�`:�
&d ��E)���6�x��̗3}A�v���ē6sԻ�߱(������-��2 ��*Gj�K��^��ں�*�6��N���w�00�o��'`mj\���8���o���dobӂ0ǅ�O�R|�h�vn�{|�ֿ�v������_Pu�
��j i|���ꎿ*;���֊��srZg���{��c������������-~U ���􂺼3�'��倫[��T�I�m���;E&�窧�.a�'���{_*�T�+2bҪ��hUe�݋�ξ�U��;��M�S��<�*2����5DVC ���x�Pm���f.u,���0��i@ᩫ[��߾�C|$� Yv{������։� ;3�k{��{�}$ϤH>�<����4�w@�t��0n���YUutip�۱$�g˳^�uv1}�#I̩H>�:�}��S�½]�sӾ�]�o���ʐI$q�Q7�RB�w*�ٯ{��^��e�ʙ�O5�	�܅�eY���b�"pȏ'�V�/��=ɭv�lߢ6�ьB"��_O�>�0=�{3Ƨ����ˈ�ꨲ�\:���x���?�H���S����T�ARI'Ḛ���Vr����G��y �i��w
�eH��FR�I���q�(\�R�j\�q܉fl֘,E��牊���+�I����Y����5�k��N�0��~��n^E�H�vNR
�g��n�u���k}w��lH�;ӣ7N^<����^�̾Dv�n�H׳T=����}Ro���+�� m����i�3��h��"��H>�J��Ţ�C=��x8&b�XtT�g>�S�������˽�v*�^�RL�A �"K��y}�!��(U>��/��(=ײkD�O}^���I?��L���3�g��r���ї�4N��clgl�$V.�@�jz�����f�e1�N�e�ꛝ�w�)�fY�~����y�5�sck���ܓcYɄ��b٩	j��E�k����蔄A[�����s\튋�k2°t�a�8Σ��v�sɫBY��
�B(��F:���JT������y�|D���TKl[��2�l0�Tmq���Kn�V٪��a�,��u�TM.�����PțV��l��SE"�����T�f�.V�
WF�Y�~�~��v�XƎ�c[1*K-G)�ј`��4h��Қ�nr��=Ӕ��A�,XVC��Q	�X����|o�>0-쪐T��I�`6���]��!{ c���񨞽�ޙ��o���z�;�<�����
��[T��&}REcVyc�I��z/f�O���>�!�f,͹��� ��E�\�C+V�{2x����X)��g���5&g_�����̏{3�#0����6��c��>��m�|�*��=������d���&�m����F�[E�q(�m�B�GL6�H��Y6H$��W�I2AH�y�����k։�B���_������ø}��EU"�C����k����z�;: ��gĲ�Cs��\7[D����>[x^Q�)�!���޻�4��ׄ��Խg{�'X+��<�H�0wq���Y&���:*���.\{v=����.�q墾��*�
�1���߰kǳܺ���ŵ�?Uo�S}�$�ɞ��O8��*��{*�B|<��o��z�D�>��ƚH�lw*|>��ʐUH*��p�y�}<m�tO���(�C=U8}]��&}R��4�Cs�bŁB��aPMWC۰�SMsSB��+h��ev��&d}�ϠfG�f!��K��}�˧6�Pޝ������;�3c�231xfG���W�/�P;�{:N�ۖ���ڷwu3��kװ3v*��UK�j��G�1��a�ۢgC�An��f��TY&�p��G��n��	fn��*�0�ӭ�O�Ak/wV�\Q�eH]���/�fИN�/�� �['k{::.]լ��8w	&} �,���B���}��I��c/��B��|�YyN�w���,�y�P�_��W�$��A$�=�}*�h��}�O5�.o�d�UnU> �$'=ƹ&m�,�8Ne n��H4Z�K�c�L�-ֆ �m)h�5p�r�|?;�OϞ�z�{2=�*�b�sQ�st�x�)��VX����^@́��4������z��%������{�g<O<�vnh���誒H��xl��^���Ƿ���s\��Ut���I�c�T�>�xU{�V�U ��.�m��Ɔz�[:�8R�E���W�*��Y�$��h���kj�L��0h:�$���z6��:ީ;o_7�@3"�j�I�fd���T����YCZ����nu��gْ=��ّ���K���z3�cP���3����|��{����UH��Kt���l�v��\�A[c�X& l� ��aBM��6Y�fp�a7��+zH�A�'��n��y�P�����d��f�E�^�RL�} �:��`����*��`�#��Τ�wq!���]�I�Ӷ�g�g�u�5�T��RM���jf��(G��o��o�{�H$�� ��lJ�c�eH*�ɴ}6���Ç�Q面��RÖgs*AU �$�_��f������js��j�Hg��
��"����G�=���u;�f/f��6�1gk{����8�Y�;Gn�X��3%"YZƺk/*MN�E�-�X��^7�ݫ��F0̒� H��@h��	�m˙cK�q-���+Һ傘0�u�sbu��Ë�p�m�f���A��2��e�D(�K�Y����h�CEsm43�0��l�ok�c1A��ՙ�[A��Sh%��I����%���6͝P�aFkp�Ƒ�v�3c��ƛYn�\U�`�Ь��`��t����[����-.-��Gj˕�IA������Z~
*��Mn�&0��I[l����;�W6-#b��"�e)S	MG�k����Ŕ�˟��o��Ǫ쁻�����}$�{ِ��iKm��39�b��uU�OD��W��1��ôT�&G�d��,j�b���㝾f��Z���T�U�>�g�����if�s��}Y��=��+�Y1շݦN㺸�ݯb��0c����L�AR���;|���i���`w1[.����!o2}��f�'��|=�2�"��#�qEBʌ鮔S&�6��&^PAS�
T�bv�C2 ́D���;q!����M���8�L��H$��m(䷏N��L�@�s>�N�L:(e*J�� �3|��Z����
�ps"����u#l�ck�"�K��]u��t���՟���s�</;)}�J����E�uq���Y��q�����R��[z�yِ31�S�����.yo}Փ�}Ƕ������)��A$� &z�xݎ�]�� G(��,v:\���z�y	�</:F��/W�CRL�ARWe+Bթ�z�6�5k,.�m�#��\p�)��������hMB�	(Jb}ֆ�^�$9��3IIs��,a��Ki���Z����\�}�I2������]?m>q5�{�NT�c� ދ���ř f@}�s�z���b'�WK��-�U���fb�:��3q4:�@*�su{2dxfg{߂�ш?F������]��V�A�2���Ƣ%a�©X4qB���$�_G�%:&Z���[�O��u}�B�%F�7۹ʍY�"j�I���aݍ�Z7e�6� 2��J���tW)wM��*���(e����MÄv��D�.��k'�a�xh����Q���9n�����f�,ڜX��C�������-�d�6j��ًX����w�	IKwp�L�=�32wa������Qi���=E*�veoܶ�wv��9�O�M֩T,a=śC@V <�@�^̄i�f���pǓ!�����b���ō��uhF��f���n�dz��ыmg<*��w��D����`�6�"r�lN�Wu�RYA8ŏ�]�ҳ�/�tK�qܺl	ZN�>=]Eϸ�<ɻ��0:��x�Vt�w{,�q���.��۔v]j�zԶv���Z���W�c{��	��J�ć�v������R\�'�x�M��o"��uZ��}���M�q��%���;��BgSt_ej�Z^㋸�Q7�Y����	v��v�����q2���b�vY�{���n�'8�}��&�*��Ɋ�*bɒ��&T
�;X�Vo��
c�}�I���ި�6�S�]�q8
,H�L�b1n����ʵ�f
{n��-��ӭh�k�5ڎ��Y�|!���P{%nH�T�ġ���+xC�۴R4�RX���ئ���7"�hl����P�c5;����	�{
Dm�����
�#b����^�wnH9p����󮷻�&1;���s.Q�ݮ�{ޱA���;�r[���<:P3;�wqr��.s=ܴ����%��:.[���뻊)�T��u۴o=�~��̾v���k���p��Jg����]��>wG7wt3��|���u���u�G:�A�[�ιE��w\�wG)wq7���8)��9]"4�̔�"M����`��Q9vLR0!$�sr �k�
���cF$$�-��H��,���:�}���Tj��H��we��p|�&�6��	�B7���^5�|���c���
��R
�H�9�AI?wv��~h}:g�q#���^�[�6��Ｆ#��V{�x|��W���RP�a{�v'|Z}B`~���̝^=��g�x}�*I�!*��Zi�{<�UX�t  ��hY�;3b�2�ڱ�-+�1^��̚�v�#�]ڬ��w����R
�HVOgQ~�w���I�J���2�L��۫b��>�Q���I�*�r��+�}D�Gj{��6��ma��϶	+���v7^q?V�ϼ�8*���O}�P��|�lK�r23��꺅�v=��g�	M�~�8��U��&R^Y=P�N��St�~���y��zb�PqDy�k�i�CyL��Cj��;�ij�ǫ2����;4��;	���[�6^���A;���O�v
d^�ꪪ����߅I2��}R��z�TY�:U,�;?_�Oh������g���I�Z��O7�)=�O���\��..�h�9&!�VF��-�)ص��r���}��<'���� �uE��=�����,��Nn��V�ʐ} ��@��!�$*9�$�f���y�4o��m��d��H�4���mn�����>��u���u�Ҟ���=���xz�-����;�2=J�u�Ӑu��ew����Ƣgd����Y�NH>�d�+4lW��X�Vu��;Y�㝖�;ûos30��n��B�L���30��D!;��Y�/$VS�t�Ѣ�b�֩�k�-���d��8�I0�bFz�hX�݁���8w��,o|�8!щ�1T�Q$1̣�Ba�� \��m�rjGf5��jC�����Q��穨�.�W:b͇�(R����j@Km6�]Ņ�,.��$�D�͚%:����*%��	&�a,l�!���MB!�	s�S����&n�0��m���I��Ĳ��U�1�U�::m���(V�fiG�.V��f��{�߷�!o�WLh:���[�'\��������r$�`%�\� �G?�
��&|�,E���3ۛݭ�=���ŭ]��S�<>�$��g��<6mgO�t^Dr��UgV��r*�w�G���H6�"Վt�vm����}$���.̞��5<�pŻg��qA��K�>�H>�e(��]'�wU' f��d*��t�gKOu�Ҟ��;���ĉ9�����2�̌�^�@+����p!)�ԫ��p]��.�l�"��� �7�Z۩�ȡG�^`���[W@KL�����41��L�0,�h�R:\��w��yֆ8̀2�U8��9Z�gԜ��e{��g˕����zgx}$�} }_��x��Σ��g7���t����敃׶�
�a�Mlb��`ͫ�^F�~�U�7A�F�`F�.S��w��� x.��}_�Jl��}3��;�5��Q�Ͼ�*I84�7�+j���q��eH>�=Ն��"%����vTV�`ർSP�ö {L���_����Ta��WARLK�N����}pe���M���W����+�NL�A�H*In�#c�E��pv�N�n����V<���s�шv��{��t)�k�S[�aFZ�
f�0b2��ƥ�26XfJT��������d4�WI�u�_��%�a����_��A��&۰�t�ȂK��=w��N+_5#+Y�8ԛ����Vg�� �<d��fR�ªA$ʑ�������YCRﱮD��i�U�i%����B�i�M�k��b�7�2<r��G��ɋe�2�uJ�
ɸ�1w��DZ� +9�V�y�;zl8Q���`�I2A��ѦOQ��-&z�P����[5���o2f�p~\��ٺ�R{�O>� �����A����I^��z�Ke�[�,z��){��A����_�h�	$yVr�����R�K���ՉI�3ʷb5�Mi0�1\��'�,�I2����]��hӝ;v|�%���Y����l��L�T��M5��.��[&ø����ޫ��rs�b�k�@c3;���h���<����/fG�#٘5v�m�NwT���UZN��OjM��:�$R���v�˼ƴp�� ��� �Ke���ft��A��ʋ|뫝��IB������6u�v1D[��V	ٕ9{��\RE�l�Ě�5%���Uw�De�����U9��ه�ʹtg��ﾽ���H*I'�?v�w��m75C�$��
����*��I2B��y皪���,�_{I���if�*n3�YE�imK[R�fbQ��0C(�[(�gh�A$�G�v�	���ַ����E�*�[��I3� {З.��S�y��!{R����-�����g��!�-�cUW��U$ϤR�u��:���\�c�[\;c�c�x��0m`b�)�\�\1�txfb�.�7����z)�7�v���P2�~��ٴ����L��$�Ӏ���	���l�N�p�f6�[u��kr=�}$7ZY��٘�ԯ��>�1%���IZ4o�2Ŏ�7���+':�ns��a��6�KI^��IXr�t�r�g7�]:��N�ANbTIKD�e�ݒ�����Jh��� `�\�^3q�Ml�,�D.���X0�b��[6]�+�L�#�V�^,m%��0�+��Q�c�[�X�t4.S��:����k�Z֑�v�u�T��H�F��dp�k���;F2�ݱp�h��H�s�i35HZK5�hb���i�L�٫I��ݳ.V�L��}���������Qv�u��7)�bi���m,�ͭ�CÃ	���{w>�}'XN����<#�X���_��*��(̣���eH>�H�hI��6ۃ(�GկV^���9���,�({�p���$~M�9>J�n}�$I2�H���rS��cf���c9Ω���W����}$���@"֧>�ʭo7G�%x��>̓}qC.g��%��Ho�{��U>�ԓ>�I���m��d��r�] ��ەNΎ���p�u����e�#�Ϗ߾�=�B��Z�L���Gkl$M5�ldv����㮖a&X�8H�;�^B�����)��9�ګ��>�dwD���*��$��A=q鞬}�}|1չ�v���:ИM����nn*WiD�sA��2�n�e��[�)1qU�N�I|i�����o�&���+�3���X�����;^�fr�Շ���@�̎����I�M�@�K�m>�4Z�g��ՌmKRk��sř2=��(*0OJ�Qsb���&f�V�j�d݃}^�ʫ>�c��UG2A �&H�]�q����|P��m�=��\0���[��&T��H�=�Ν�b:�Dp��HƘ��Q\�KiٚP{W�\%�Yu�ֆ;8�6�K�Gzߝ��O���pf%w�uUN�й8�]�{G�=o;�+q� ��f,Ǻ9N���ڑ�ѿq�Y�3ճǌ/v�{�)�}&�t:ް�|�9/�
�eH*���/�)a�-���s�t��k�j�im���ѐTR#\�̉Y9R��8ڳb3��Մ�'G���f1�t`b��JE�]������2�4��;��'&X�������I3���m��^��B��H#y����ܿi���©�zs�;�!��������I3�UH$��Z=�{�q��\�{�ǻ��yO��33��T�KY��b�� �2���h��ۡY�a����+K3K@n�ۇB�Vz�ϫ���^L��Ք��̇�N��ds�#�N3[�Sg��
�I�[�p"C�Q�Y��boeB�g��.pv_��C���2�K�@T���h}��U �A$Ϥ��t��zZ}^��K7`�Uy{)�I2AV^̺S<
=�wr���'��o��2��}�>���F<����ٰU�n�)զ˚����6�6�@�b/7�5��W<�z����=0���d�2��i���bn�h%ţ0"s�xz�v|�̀31xfG�(}Fe���]�j�C��\�� ����{�+�d��4z\mr�1�7���Q�i�2�WC5�m�l�!0���%R�+-�����$�/&�U�T�*AH&�MOx�T��>��qۘA���������M�b�z�d3�������g��L�}�p��$>����.kR��h�NʩH*H�M���^�z�ޮg;#�K\��FZ�{��s$H>�g,��wK���u{�y��d
Uw+'�h��T��>���dilג<>��RHj�I�{z���S6�Z9��pR�p�!l��۰7c3�^S��d��7�rl�k
e����d��B�q>�x�[-�;�,ܠJ�U�Y���ӳV�҅�Vޅ�^b��;!�n�WMVV�vR��uй��K��U�.�T��Ⱥ�w)�+]ۻP����(5�d&���e�R��&�7���.�KB�n�6SݡwtN��ֹ�u'��{@�V���	9v�j���vK�ݰ�wk� *�59b��nJ��DkFeŲ(�t�]6�m���J�_Ϝ�+k���Ù�wȫ ��k�۴�<�d�L����h,P��	�c�ZS���:4ƅ���T n���R���8�X��4�ڃgs�~�Z�p��B:�v��2t�����i�s6����.��S��E��)��_x��l����{O:^�̍������(U��/M��V��M�&�u�Ƿ���vGO�c�R�-.W�º"�y4�
�Oh�;2u�PsW���Uz	�SJ*�S�P�˗�t{Z��9 d���U����n���̦Aǖ4�a&��v�#]8����>�P�m��5�k���'uJ�\��)�dR����os�KZ�=p����u�>��\�QfK;Yd�â���Ã�)���*Q)�&�A��N�W;Q��`N��g(�4^V�:�6mJ0�k�V�,+�4�7�^.�{ɷYoFS�4�taڸ��{"�e��]͕�^��`�q$�3F�a���{�\i�\[}QE���<��F���/�x��41�ۗ��6�FD̗���fRj=�ˤ��b.m�b������k����^TE���wVLE5�DTI�]�X�ʹW0W-�r�j�p�]�b��r�Q~���ZL\��k�F��6�F��F�L�]֎X��9Zf+~��������cIgunQ[>��� ��v24E'�Z�۰�ʋ��\����˛i�L�9���5��ܮF��cdBe�F�شnk���g�[��&�y�-�78`ƃ��W�vܓ��lcb�Mr�IcE��6����4\ۥQ�5�6�wwLk;��V4X*+rܫ�\��ܣE��\��������A���=Пg�|�~GR!q+���3MrK��\ׂ ��5i{$�mu��)2�7)�e�޴i��یL!54J��J�z�W��f���4'������99.yf��X�ݴZ:03*�öR��k��4��%ƚ���a�L�����݁�&�m]���x�:�ʺ9t5]�LkjTpK����%���P���5�ڪ�C)5�&�V��X�YB��]��ͨ*j��4�6�����Z��4�� �1.�g.кP���Ku�k��Iu� ù1k[`M�r�W7gM#	�Z�)���Řs��ƚ(�٩��ʣ�۱f�9 X��1[&D�7n��-�v�� �-^؆F b�B��X�e�B�,�n�l�.ut��Y�ʪ��whd$��l��A��C�jc:�ĭ�k�P���n���"�CKu�XkQ�̳B١����ĭ��A�c*ǋ��Ť���%�5���t+�v�ԅ�V��Lh�L�h0B�0v��jMM��c(�@���y<�[���X�Ԑ���H�].������J� .&���Ʊ-��@��6%,%��bT�Ѳ&؍�]C��U�ybk��k�8v��T5��46�f���`%Ҭƫ�ȳQ��c]5t�m�����2��E4�m��,6�k*Ckz�\���8�цT����i���3�C����e,`�����R�(b�y����n�R�8����(&p]Q�� !�ѢЖmC.]@Ynh1���,���YH��+�����9Ȥ���\�e�C;�]a��֬�Z����4
�hv��⻙���My�ֺ�]cr0��XfCS�k1i8��b�ڔ�q�V+���eJYwj�(�A5�h�t֊�-�	c� ������V˭�ln��4T���^�H�񄭚t��
 �2k�,�r��nF�U��r�ʹUUU[H��[���#��X��2j˕����x�"5�Lc �9q1����T�jL	1����d��n�$�V1�j���Un��Hq�/��Z���������4#�0s��dX�
�ѻ�(f�s�M�P��IK.t��H�֠4�����ƀ.%.��٣�KGuJu���Z.�2�͆�W0�b�<K�j��!ZqLkYx��pY�b$\YQ�v�r�(�2۪���~����Ģ�,([��5��%�"��r4lf�e��h�ͅ��m�=��K�9ǳ#���s׋yL�<1��a�ݩ�5$�bp�mȐ^�!����A-�"��|�9�]xƑ�f|w�W7���ዮi[��qǯ���n4L9����q�����@��CnD��"�R$��Grj�8Y��j#�F��]���y���כ�>��]�F�}uo.}U�T>�Ap�%��+���ST�Ǝم"+�%��7����m����rۑ ��y6���0�%�)�
H .��0��aU��;��A=|����כ�����x��a������ ���f�4�M�n% �x�%���sF��s�GR�
dO���IJJg�TF�BKp�Am�s-�]��~6�FH�n ����v�6�Ŵ��> ��^�U�/�K���
�����)�H�������vu��%������^�v�>�^��g��
5.���r��C�kf��m��=���>6�n��~ƾ�SS�a�م"*��y�N�j��ݐh�۵�@���AބA�w>!�*�ɫѳ��te�Z�gb�j��N8O_)!��q@�[k�ߐ�����b_8�* p �y"N� >m1��X�&�R���C�� ��C���;�FX��|FrŸ�-� ��"�B�mfMU�>��{&�S´v�)P8�{qȐp�n*���|��I�*.eR\�Y�-ƀ�s���5����lLUV�LL����d C���a����1ױҺj��N=]N�J�p �/wEAm�6����=ı7oq�sax���8�<v�D�1�.��	��/PD6�0�T�J�ޫH ]Ǒ�� ���Am��	E;�M#e6�}|�Kk�!���n�xj<�Nm v��ims�V�h��:�-R�[D�P���j��$����p�F��������ɼ����<IR"�� +�"Kq�Aۙ=��W��|�!�H��Wts�ג��nU�,���^�<�+2g�=p�}y�|Cp-�D�ϛ�����ع��kE�\>3�j]?R] ���P^!�"|[Cp\oXS�"6��JB� �l}�"A��JjEf���qu�PD�+���e+"a*L)��7z�������ћ�{&�i���\��'r�To�i,O�w�'Ǻ�6�!�"|�#��=�ַ\|i�tdϽ�N�U%Ob�#�ŕu#� ��RCp-��O��	52��S^@��"mϛ�B�Y�&�������ط��ղ�ʗ	�^ �� CnD���q^!�B-㭄�m&�sW���Ŷ�Fn9���:IR"�s` }j�wyv��$6,a�\ξ9�h�]W|mʚ��C���V�!sR�h��uo�).���%���(ܪ� +�������۟H%�@�A�Rx����W�w �X|1��Lu�䫨YA;|���E�@�[h�xx��8bn�h@��&DD [kB�mxmM���������l��G`��\�=[��F��>-�!���6����S�U�T�SQ�y�����UA�b�ޙ��7A-� 
�.YWgl���$�B ��T�Ό}9&�2'C�*D_y��͑ ��[S!l��'�Ǜ�^!����EP�:���7�*vr7:�U�,� ��RAmq�[jHm!�r��n^�Q�ӊ ��>}Am�p�]��]2^Ug�WH'v/�;�|Ѧ�@w����[�/�����.^N]�H��ӊcn3V�.��Β�E��6y�$������L�����l����CC������n�;��/l���I-�|���鄳]Μ]q�]�\u0�� �ҵA��'Oq��Cֆ; �YWV(`�m�6 ��2&�0�3a���0���WJ�Du��P��h��y�l&�cC��ǘ�͘&1e.K,q.%����7a2��rBjdh�`hL/$9F�#�Q(T��36���Ԩ��mԲ�U1�N��V5��D.!]j\��#�6l�s��Q`[+�%�U�G)�h���B��XP�l�V�+��k���߿��ufk+��VQ]e�6j�W�ņ�{5��g�w��{���7߿k���g̪�x/#3����=t�هw�8���6Ԑ�[�$w�`wW�#� w �u\�}�'��ˬ��� ��@�� Cl��a(AiB|������Kh [��-���!آ���EZ��ݧg�B֯[��6�^9��A�@fPA5&�B�7�Aւ#g���c�Qε�D�>�$2]]��#��r�{c���>9ڤ�א%��s��b�:�Ԟ�P&"��ݶ�R��w��Hp/a���m�����zf�=@�F�]��A8筅��ft��Ejˢr�5�30P�1
d����u� � �p�A-�02�!��-��bF(/��Y"�dI���/۟H ����t�c�����#S�j��ħgN(Y��.��kƣ罦�2�ƣ�rH`�ה��b�%>}Fn)�֪_V�eER}T �C�;�g�}�\ЬϪ>S�\�*�d{�o)�6�-�i����a�mj`�k�� Cm	�n<�m
�
��>H>���ytpw�ʑ��9�5~v���ψ��q�j6�镄_G���A-�09��!�˕�zLH�����@��ZY%\n�lg�8@��Cng��!���v��T�א�)���Nv_9��Y���R>mpmR�Tn�8���$.&L��D)AD�&9�h"���v���L@E%B�g!R��/�~{��,H��y�T�Jݮ�ʐ���L�0�
��A�ۋ �1�ϋh [�"�^����\@���G���̷�լ�[��Ĉ�lA��Ȑ[���Fػ��w>�A{Ch"5������S[�&�
�ק+n�3�屳['ZǤÞ6�����v'�����^�9�{\ج���z�+���`�ΰKo/���� ���|-99���*�d|ƻ�����A�m�7h\���k���{{�,�;�$�@���@R�P��77�!�����8�@���.�o;""X���ۨ [�|�S���ne�r+<��j�<9^��On9����jDg	̀� ��"Kp�n��}r�'���IsX�#+�t]oi��E��-�K�rҊ�J�]=ߟ#>�����LO~���PL�:�x������oS#����U���A��RCi���k6Tc���qn�BA�����T.���s2���x���CmlL���<�9���n��)��@��A�
�$����Ցf�kP�Fr��"|[�!�m
w�7�OGwP�����J����]f��9��W���REuR���ԕ9�P)ZgoNk*����}z�Mu�p$�+K a�a^�4U+������;_�,�<]�}�*��p��w,fk�
�>����>=м}�����"mȟ�Y,L|���,��%����Y�9����D� Cmz[B�u&b�W�^���,�)��!a5�Hu*�qZs,vt�L�j�e�D�$�fd��eG��Z��^n(�m�An��,�j��B,�ڤ��	 �ݟnŐ[A�BKp�VdvMwv�EޯO����;�-u��|�2a\q�r�h/�r���j^節?����r$��ޘ�֩U��-R\��s��Ȝ��L�Ƕ �A۟O�h [�]>�_zb꺳�E4}�͵!pqM��b��xR��q�DNL�&3p��ghI��p�m̂n ��6�Q}!��͋��|���s�]g��:��W}]�H!��D[hobA]�u���D�̊L��uZ��q��1s0-l�
�)�ɜ�D�(�C�M#KiaJ����s�(�S6.�8�6!����O:qѨ��]*-�3��BJ��	�X��^���Vg�����1-��7Q0�j�,
9�[�[5%X�Tc�P
j6��5&%�q�e�ˍ�d�X04�� :�b�֎�6šlٱ�j��q���.l6��..�X��V,+�],���b���6hm�(Sr�+]��ix5K)�F0-ٲ�����3*ܲ쵃3<�?O�u
��A��4qV2��GP4���fM2�Hk`��B,2�Y����f_������B���z�k_RmNfz�zB]���H�5�#�O /v��6��nړ��i9Ժ�r4|�(��7���".� ޹��fDl���9�E�L�6�>mCmy�ض#8gj��=ǭ�C��޳Y)\p>��$6�-���mH!���v�e�ʈ":r܉<�[Az�mt�d�o8{Uy�������DOm)�خ�`WU��Ƃ-�͵�m[��$���� ʥ!p�Xtk�]�R-rp�"@-ǓhM`��M�q�o0�dK���vKQ�i��:���]�DT�y5��5�2�N���|z�y����mUg��}O8^JW��m`���#�W�>�j�B��Ԑ��";�4(�Ac�H�L�5���7w�F+�fX������#�5�k�����r�N5�ԗm���*�w`�"�v	��2`��W<�l}���?mW�U�wy�ܫ��L�>���!�]2\Ҿ����h#. �����@������6/�z26�VpnQf�m�T-w� ��>-�6�m܍�Y�d���9�@��Ϗ�ASq��}O8^JW �r�G	Ⱦ�S�=Y [��!��	n �������'"�\�sXk(��p{����\��D=Ax�܉�m3�5yd�FE� JB ��Ȓ
�	+��y �덍o7\��.G�q��r��ޤ>y�s���Am����r�g�f��*�'\�^ӘT�c�p,�5�$�6�!�>�7��Wb�N�О���ɟ��q���|��h��� ���כ��b�UEUÏ��#.:�"mϛ�6� ~O�U���i*�ؔ���я���O�u�/�{L�E��������$�+h����v��k,
ѮA6��h�|��wZ�3o�WY
ڰ�3�C��\�a���B�^�kR���]d<ʺ�uŪ���fM[h7�pf�"l\�-{���n,�|9Ԉga�^��cv���w	Jq�H�ș�r��v�Pd=�P(6��#�Z��w|�u9�\�#*^<N�3$ӳ{ݤ��UqG<�1����uv}���e��2��*:av�̓�%�R,-v�9j�ZU�^�ƪ�4��hp���F�j�=��4N�wǤ�l�:�0m�<=#U��U�Մ,�m��6�+C[�-k[�(e!Ii�Z��5p��UKd^hͤ��nQf��f��AM���=�q�k�~
�T��S�<��g:��2x�גZ.a�V�n���y3"�&5�a�5����I�^�u��V��9:��z.]�Ȧ�ņ�<�:)]�`[��/&>�'bϯ_'�r�� \�������C��r}�f�P	AC��#Bs1�M&�ם�U�%�f����}�df-��}CZoq�z��V[���:r�v�s����`Ğ�cx[x������7��0-��B7Ru% ���g��pi���`�'gFP�Ơ���#J᳹.���;�.�S����F!����Ƣ7�uM�G�0�{L��"�����>G�՜�hky�~�����+k��}��.;�u�<�V=/ss(��pOU:��̡U�wF�p��@�JCP��Cj��y�Ė��Ţ(�$�j�\�1h�-d��ݚ�$�"�[�l�snh���EowT`�󕢣&�N��K�������sEF�LY�h�ۘ6�f�L��1_�-���d�kR����`�Œ5�ܷ$���~�\�5y���+��EDj�������G��������[E2m�>�ޮQ�~5�Z�W6J�6MX��Ed�E�E�V��E��I��r������LэE�V$֗u�X�幧v������-��ܝ�m�;F�C��66���6���_u:����?ܼ��J�= �� ��"s>-��n=�$��m��4�Q�݅�	m�հ�1�dv��Ī� A��b���0���ւ6�O��A��m���J����-N+��wLU<�R��Mw/O���p� �ک9�vihN0���݉��GCG�)k��ج[�63 �9ΡU�3k�z�S6.3�]@Df���y6���)�4J��[�G>G2����E�o��5E�����-� �ڐD��Dl��Wp=P��w)����<#�]�1B�8�"�s���S��v=A$�X:�ɴ����\:k����r���э%q� ����栋p�ڐCh:"A��Xv����$��/6���늙���Yy�K� ���R�"�EHkh����e��Qb�ms#Ly6����E��Q�4M<�3���X��]���n�۩�t�*@��u_
���>!��Am��Ǜ��(����#�U�JVi�%��kaLP�����Ƅ��hpn6���]��m�V�8�3��B��gL�mXf40Ax�Xn�i����*ey�A7Ѐ ��/ۙ��h+Rmn'�U��cI\p!�p��7J�^ڠ"�lymO�m An";��4�կ(�����@�AK��R��f���TO	��/PD6��s��Z��Ap� �R 6��@�㍧c���w��a����:�P��� ,͑%�^ ��^!���c����,UFx��k^��ޔ*���u/�4�G|v�O��x:4�UD!`�G�����-�^ �܉�Y2'���k�)/qoi�|�y�)���WV� �Aۑ>-�{�S�_
��&�	�w?+�k���@ ڛ��Cw�ҞH:��n�)��Ӓ�g鐸��B��\�r�hˀW�5��������a��Y��G)��m#MChFTM���l��<��XlE�P���M���Ym iH��L��l�6�`;�T��MR�Tp;Fۙp�*ls�Sf4��Ѧ���$`�G!��r�J��F`�S�a�jW��Sq��j�4
Rʽ�n7�m���!l"��c��]���؆�!�Z���@F��:박#X��e3�冺+�ߟ(^���[,#qx�Ҳ��թkYS��*���(U	�33�Q��j�H ����%�P�6K��0��P�zی������ ��� ����n���>�O;iƫw�;�'ǵT�e=ꬩu��q��{�r�9�!�v)vH��oX@������yy�p����k��Y};{5���	{��;��E�^"'��%g9ce�j��A�@�[j-�˃���ѪU\>7³�N��Ni�j����[���/[@6��T�zuK=.�p�gEҷ�q�N ��� � �n��wfV�v��"B�B
��*PS�A,rF]�X[�䃣bj�����a�*�׽ϖb߿�'Ÿ�p+kf��ڗgzv�k=It�ؠAz���D���-�[j|C.�w/c�|�9�%.���Vw֎���ι����Yˮ�o��k�d2Oe���aH1c��&r���h��Պ����z�����"8�Ss9���ɣ}\6eP���`/}z�H-�Xɞ"C���0D��*�D����� CnD���0w�Y�v�-���W�1�Rq� �k��A��n�mH!�p`6��f`X ���v=m��׳W�m:���mVz�� ��DV���ӗ%BpUu!���3���nڒ�A�&�����Ҧ@���3��rE^�F�V"�o`"�7A��B����RRʁ31aX�P��@LJKɐЍ�pL=��� ��kmv���at����!��-����_K��j�Tc��{!н��L��h#��mO����ni9Y=#o��E!�� ���V�_Y�5j7�ڜ�%ޟ=�AP^!��8��t2�N[�적��}٫�^n(Kmb*u��Yʅ��*m�.�j�鈯!]~wJ�qO���@>��S;Mɻ�����ݒq�����6��BA����X��E�z���鞢+�#�aX��� ��D��O�q��Q��G�D�����Ϧ|[AE�½���{3J�)8�	�jA{��L��qp$�G�=����/�r$�쭛Y��U�U���iʩ7�Z�עWH%�"���Cn}>!���mS^:n$�舟(02��TF״�m�Dʐ�ChF�,��,�ژe�m��M��w���w��	m���ޓ�䅹��J�k�;N���}�K�Ր ����y��6�|�zs�UЯV �GWH㼂�\�+��}�g�� ��$3�E��{U��,RGZ^퀈m� �����ו�OS�]*$oݫ����A�{A�ۑ>!�n#� ���yu� �k۱D�����9�ј�ص�װ �>7T�z���2ϯ�|wFܷ$j�ȸ!I���E���@S�!X뵝�KJ�Y�NvFf`sk�뜑���"7���ϛ�A�h"q��?x�P�AC���kcm]��s)�����"�/6�����-{�_-�nH�p�7g1L�3�B����L if*X�6p�"fLJ����T��$��C�UN_a�'���UzRA�:�V�LQiC�^n<����:���t�(�,� ��E�u�Y]F���Z���̀�"�ϛ��
ٽ#��R�dX ���3���v�qձF6L���O:�;V��jS�k���A�|[jHm/kWUڹvµ�轜���"�כ� ��[7���we=˹���A�̈́Fv��\LJW��`��-�ڒm[�'f0le�ީ����*["u8o�X-p@��@D^�$�>��ܯm?444��TKΧ`��&�V��T�d�ttf�Ƹ*Q�y�R9s9��M��
[nP{��i��K6Qib�ʐ�܁:d�yQ�`?"�nD��)ci�i���vѥ�B��4%�l��0�a�͑����E���퉦Qm�9��Z�-u]V\��h��fM�P��.wGfQѶ�53��[E�X�,H,t2�4�Č�b�m�\��;`ơ�ٕ.M��㰱�����Ħ�lkm��*�j ��a�˖޶R�m�� Ysy���H+k���u.q���䴗�K�h�%r.��q����Ԩ� �܉kc�XZ��k�t�}!��ty�
!�>�7 ҸW����,�T�w��wi%Y֘�@�	m��Ǜ�@���W�X���#k.��kAml�Ud��=8�r��$8���"evTfX��Q=��F�) ��@��͵rV�c̉��T�8�a�%`��@�� W�D��x���܉s�^�;�=h�s��
*n��s����j��q�jAǯ��.r��9p����Ch An M�[��t��uQĉh'�7�K=
���ϒ]��� A��b|[@��y3s�c���#ޘ�*�s1t���f���"��n��йV��,�A�fL��Tiv����Am�oޒs�s#w�x�g����~x狗A�dI{��D6В� E�1�@�xŜ�|f�^R�H�1��D+�{0�U�nLn�ܻ���O�C�0	���M��5��@��r�B���b᨞��r��J*��]~p�#��>����v�2�f�ڴ��sR#5[�J��m�۫�g�Ԃ;�/�"mȟ��A<f�J��gg��>&#�i�J�K� ��@�7P���E�@;�t��ElF��KAq�آ	m����9WK�چ��b�	ހ��;^A�ŵ6Z��3�@���>-��6�!����7zqnh/�*�\���ׯ���a��G�\׳`Yn ��78DZ��ͭ��q��@�nf%D*����o#���l{�X�Ե&�6Y�ن\��wy������"m6�w*k8�}[�+�$;/T�����^s�"�!�H���^-� ��6��T��\�o�p�V.��]�㶚�,R��/Z�q��do���6�#���	�m �_n�a�E��f�u��"��Ý^eQ�Z|P�QhV)d
��U��B',��T>N{�y˻D��� �aVvI�"�P�ou��f��ws�c1�m5���sR#5y���ڐm ���v�;�
�B�{c��^�ܩ��TWOn�^Iw��D<7�U[�L
{b|Ck��|[jHn-�Z����e5�����Ηi��b� Ot7�|�X�Q�8wMn٬�
��虉%M��I����cd�$v�sP�4{R�la
���ϓ{~���p���
F�]�rΣ��x���C��W��	�p��ʰA� ������x���(M�;���^ �A;;��8����R^Ip�Ml"PD6��+�u�S��� ��y�Rn-� ����k.���wW+bn���
,Z�=�^�[�&�@����#:����������|Ch*F�U�t���x���A��Wݸ�����aB�b��$�G2�"�5k����H6Aqu���չ"Ҍ�ѝ�����݁�[���毧���m���8�B ��������nD��9�N$���|��{�Vi ��݄��� ��@�����sє�������<>[�&���9��% \ꡍ
\��Rͬ��欶�c�r���!ןrC�����S}��N�uOm�Qb�!�{�N�[�v�a�ϻb�-�hYn �faT�X�5�4�r'�uH�*��]�1����q�k�j��ţ9x���2�〈-��� -��;��X9��S`��wv�I�<���כ�`�'q��ܙ��2u�V��*#� �� ���_g*S�C���Hص݁���:�|��X�B�8@���!�"A-ǐm ۱��qɺZ�{;R��K�;u�o�M\{�[S�3` [�A-�����ޚh��_E��R�h+��B���`_=���//w�n!��#�x��mF�����KW14ʒ�X�
�ѫFŲ�A�f�X,WiqG�ɗ�Z��(�vˮu���g]�hJ��͕a��B��i;ξ]����������L�W��&b�ڷ }��b���Z�y��+���C�!]d��xa��iQ���Ln�<�t)K�+1���q@ga��]ڮ�vKݍUϓ�]����V{Ȱ�ea�4
���&�K>#��v1nMݙٙe׀�yz�mZ6����4�9'��@V�Y�$�ʵ4E	Cf�Uh�H0��3xJ�#�قÊ�<�A���z�AW�*�J�gs�.��LK���s]����;���6��ز�(�"��}}���s�&�u(�FaQ���XE�qրފA�o�L�ǹ!RL�T���Ұ�G1�;&KQs�j����㪅��lѭ��b��.�����:ȯ��y8��2��
�]���sbm]ޟ`�AM�[�^̙xh��6� W��a�8�C"�bcU���%F�
�*��̤Y6�&"�$;5��nf��#T-���3$��[���u�g`��}h���P��E��Vu�x�ٷ}��#�Wu\���wZP}"��}D�#jr0����+n�0�"�:��ъv:=� $�-�����7k�W}�*��`�(�ǽ+4wd��	i�6�)]f�H�f�̾L�"_3'U�f���j5!1��p�a�y�f�����h�\�+���6s����l�lcyvZ7:Z��]�E���oS���&���^���n��lc_������/�v�ɪ�+r,lh�֓Z-�,j�U-�F��Ű����,UsZwF$#����\�'�sW��mWϾ��lRZ7�\�˕bM��G-��-�F��ت1�&���nkQ�;\�2_J�)H־��QU��1�6����j�y�m��[���h�k&�4������ݱ�n]1�Q�j�ܫ�����_��]����K��ٖck2M+�pQx��klVԚ`��F�Z.n��)����ay�L��p�`�5��G�0��\-%ڬ���-�L�+â�CQ�0*�� �k�]u�]��bW@Q)�y�
˓���
����i����\cY�6�ڬt�\B0M �+Hp�╠m2�	R޴`WCV�LT)�.��Ĥ%�#R	s�`�ҡ�PZ�H�P5+�&��KCi�X%.�%�Fэ�Ba���M0�87�0륵����e�	òCm��]]��#IE�X��#�����w��k
ۥ����q�LW^��B0��h�-&vL�:g�W�ѹz֤C�E���Q5XٴW��v*�kM+m��uֈG)�����X��D�ܵ��v�,���m��,Q����e J�4Ŗ,Ѱ�i�*Ֆ�����Jq��@�;eJ��3K�N�ٝn�)M���L�<���`�إ�9&G/-Q:�\���.�P��(S,�T[[�����,�� � Y�3X�WË��ն&�v�
�f��*?��[��̺�l%%�1	���eFi��]��)���L�%E��aq�a�V� ���Սz�d6�	KuY�a �T+Ik��i��L]�M���Ś��!s,����n�ָ��V�1�����X ���
Z]3P��D��j���lP&�K��쉈��U��V��m�-V%�%,���x%�5�Ŭ2[��8�a�
�Ke����4�".L�*d��������j�B��k����Ɛ���da̖�/7M�Y��,��ƚQ
X�pM�uΚ�]3-���2l	�Y4���)B�u5ͺm�m���Y��XF�+����Y�ޫ�ݴ�B&u�b�Y�☆�g�̷��bFj�JgVZ&���q�Y���m-�1�E�mxK
�������e6sL�ʪ������r�Z[�U�E�6��;CB���kV5��$��y��z�9n��B�c�U���YB���b�Fh��4�����3C�4J�l�9p\jj��Qҵ���6��7-5��Q��ԙ��!H�8hG;:1k��[s���*K�ʷ��ͬ�#Y.0�:ٳ�1 ���V��ٷg6�-vh�E(����YG$8&�륂��K�V٫��ճ���)3�;/k3<�<����~�i�Z$�G7;	g&0)��P��6U.	`T�vF�m.�ڹ��z��hq�� ��dO�p��"y<U]��{v�%�D� \�#cm �z����� 6Ղ*fҩ9=wp�xI��#���9OM&;����\'�^�'Ÿ��dr�m؟7��݉��hD����&�#�4�[ۓ7�]]�n|Fj�����6���#nb�#j�K�*�����qW^@!V��%�H&�<wE������7�g9����Q��^�כ��j�e�� �����[tkn��*,R�k�:�dO�p� ��Ӈ|뷯_(R�GT�j)�����R��2mu�!LƗ	�qW5�]?/ߌ>�!t������mRf�:9��eE��MTq
m�v��.�s��j�g/n�6ԀCin�6�z�s�:�����VF�.�e�~�+7/7�2ǆm<��y�9u�n�Q�����#�WJ�vXЊA��DW?ݼ�~͓15*�j�������oa>�S��*����2����� �Aی��9�׫ۈ#��׭H��KmN�)k:���W7F��wڨ��K���^��q��h"s"�llTOC�n<���Gw/O�B���{�t�Tޜ��G A5�H �3hBvř��3q�ouy�[��!�"An)d��Վn��!���w������K�[X�@������a�M�c~Ϸ����}fi���\��	�BR�\�ͨ����0�d�-!A�,�A�����1n�ԋ�ޙ�,�ݦJ���*�R��Yڄ�p�n!�"A�}���Ӆ�y�W\���
�$�.���Nd���MTp �Y�H9�"�P���p��V,!�@���ۑ �-�^�fY�k��>���jj"��l9P��3;G_b�*t�{��؝&�����u��rI���������e.҇Z�e&+U���2����~!?u��K�H'n��D6�|[A�(�j���(tR��{z<�m_c隣`���2TX�� Ol�{h8��21k!F�!�"|� !��Fε#��-�o �H��z������MTq�g) �A�Am����]SWQH�o��6��ŐV':]ڐ���E�[B�5�%l�S��j̍�^���=�"|[�n
��vOJ��6��t��p�\�`#v"�W�6��P �ڐC��kr*��7Ё��)���7�N�v�*,R�k��^�'Ÿ5άR��!8�=������y6�!�>����|�!��lF�m�K�67*��A��#6-� ��Ԑ���3�v�Ge�P#�В�"�A=��e��5��'�$8�D`��w!������%���#fACf�F������Ru��rٱ��&s��[�`�v�-ص.+oZ�;�t�bG/r_�ǣ�Cx�#�A�Am� ��E��?��z��5��p����b���\FK w���hIn�Z�U�GC��)�e׋.���P1��A�1�!u0�k؍e�B�Q2�)a9��\yk@6�	���S"$^�oK�7�)5q��U���n�8�L�X�=Ј �כ�e���7j�w��~:��o!+���޼&⳴��%�;p�!�n�3�(�[�d5�����p�Ŷ���"gz�nMr����ǣnP��>;�^�q���BqGS���b"�yF�Ch FoL���U2e���qszrSW�\���74��aE����^3Q�oyI��p6�H-��d*�]!�)s��^�9�r|�� ��D@6כ�M��{᝵�g,��3��ї&�u�\��hΘ� o��.e+HLy�{@=�1�q�;dޫ8^����3#�V�����~�s�ך�j��)���.���jTY��a։���tM�Ɣ��� 13�9���6�aZv&%bV�:[4&��j���E�-,���KMQ��� #5�n��͖�5�2�2X�ک�	�T��)��vY[6A�\��v�l����WV�=�`�XC��ql�u���ʹ��aA�b�����e���9͡�+Z+��ni>}���V�YmW]�q5��71��D�;v����.s�#A͹B��G��) �Z�	m��眧*�b3x�hE@Rf����J�` .�D��D6�m�`��մ^;��w�n�X�M�`�B�P��{W2���'}\Ԃւ�;Y��lJ�7P@���Dۑ%�@���T�޸�u��s��j�p+7NO�] ���pmψmy��:D칅�����p�A-�#2����Բ7�6����p;�F��B�����H=Ј>�@6�H>-�6�6ܥ���2�a���(!R���{��3{�W�\Ԃ�n��~{���>?'�0�	}L�#��f�`��̷l@����a�V��w�}�#,�|#e��������Ow'[oX8��ï$�E�ᗡ�SrpN� �h"-��my��	m��o����l�LL,�Ƭ�e@Ɖ̾�}D��>fv����Tf����d�����s�B�+�-�"#\��Ud��-Mye�[E����Dw�s+��g'c6�qv���w`"/uy�qǡ���W��sP�wcɴ#�O�m����e����U8��:��	���M\{�[^���� |�RCp3.�l#� ֜�:kg��d6�=Ѯ�ްa�=�~��A=p�T�x��^m��z|wPE�^ ��Ԃ��[���A��J���	{6�(�v��^��A�^݀�;�"|[�&и�2��u�@���jт�;[�i��1
f4�1�iM�@�&Tę�����$�D>��mȟ7�b.�7��Ux�W}���zӘ�����>-� �א%��f��dM�[�!��D����7m�9�w�K��p�-��m����q7pߛ��r�|m�$7x��m?{��[(�~��WDa�w�I�V\j�T�h��Q]t���ԷVT�^Z�C�}ҳ/1=޽w͑4�l�+E�ˆ�����.��]���p>;�nl��^ ��m܊��wí]���d�j�[��F=�	��h .B���ޗ�U�����A ���p����|��A���/M���ח���8܉��1A�Uf���Xsv^��;]��$�A=p�#��m�tY͹��s_���䚍��J�Ai�q�R8r�,�`�Kr渌�0`�33YQ���^��y���R�q՗[���s�2"�u���D�:���`���Hz�^!�2-�!{�G��o:�S�t�?��Q��]I7��|A��H��dd%.�@Õ>#� @:�"nD�[�n���`Zt�MuM��k���H �Dc�k�A��yj�Kw0T��;� �^ �ڐ���{-E�m������B��R�ʴ���)xI���Jw׵��k!��]����CV�dՌ�p�$��:�]�/�nFA�!�-��Q�q�����}����ǻ�Cnd[��Cp�V
�'�7�6����A�}w9�}�.�Ȗ�85�O�:�E�@�m�*�\%�����DDm�0�q)w%(��ScZ�k
K2QIk��6H�܍�l�ȸ�M��F�BKq���;�L��fg��6�[<�><)�]ovz[A�Am�11���==>�>�{��Ź4�.{��A��>��][�"Kq��*����<$p�AO$H>;����n�����b���̹��79۸v���Mdq潮�� A�m�7<�Q�����In����7
����o��Byw��H>=p�a�SתJ�D�ϧ�`"� |�R-���p��U��!G��ѡ��h>���^"ޯ7Am	���U1�A]�Qelt�D�Z]Q�,��63�h�/,M�m�֭�!�#q^M�IP�4ʇ�Jc����Ҩ%���0���Cַ���6v�h+	�0�,4��)B,Ի��Xͦ�L�j��8M���Qe8tm�X��6K�l��h���C06�lb�/]��tKh���6c,�Z<T���]��q�$v��0�0U�&(����J��YeF0�����nn��L���\��;%��K���qh<�5*b�#��Ynh6�;VU\��w2��~���r&��e�Z�B�Mr�X���4�5�ۊ�l�F��}M�} ��@��CngŴHQ���݇r���G��Nk�k����"�R� Kp#6�SeLM�N�ؠk#��)tD_U����]�g�] ����"s����9z�Z^@N �]� ��!�� A��>�rg��ml�K�Ǖ"9�"/� ��
�Ȓ�"mCn@�rg/N�w>�Ax�n}>n!GVNuo\k�r�Gx�k����*�;�~] v�~!��r$� �*^H��|E�UUq��Wn��<�C�l Az�6�|~|g���^�	�>���U��&˫)6��r�0fd�il�C�c+w۔=_�����h [��mE�uT�6�z�ȋ�.��ّ�j�
�>�!����>-�vս3^�u�V&(�P��������UE,�Z��%fNn?ScV,`E��`;5�:|en�6*�� �s����*�<a�����O�!HrS�?-΍od���k��@ւ�n3���b09#����k��,� /6�In �ܩ��"ΎC�{'���Q�nO�3Ʈ�a@z�!��!�n��%�Ul��"��yx�ԅ{�j�ܶ��3]|���!wt�U#3N���r��9��݀�mȐKq���q��է��dw��hB�XݭΌ�b����A �r��A�"�mNFg��5P_��XSh:&wk����l�GQ�^,v�b�7T�TЇ���W�����z-+��w��ʼ�(Ha�Cg�X�Q�~ �yo���n m�!�������� ��R"�:�5OY���thE���� ���-�.��m���E�L�^� ��m�[hO�W�B�O��)�9��+�W]IU�;N��P�v�5HD%v-@yn�Bh%�e%�3��M�>���"]�_���U����7���u|M����-cY�V���57tъ��6'e�ہ6�o�0;�l���Ԗ�W�P�'Y�g\�Ŭˮ'��ġ�0�p,�YԤĤ��F��Nun�ȵ�����Sإ��C��}ƹ[+�vːߚ4�Z�v�#*Ӊ�"�p�PJ(����Κ[(G���uu:�:];Z��Ю���*�(4�6�/��5�ɰ1��h�5��������5i���k{�MY�T˄��b��!�cEXF`_mp=��\�n��o{E���{{�V�R�%ʸ�(���e̕�T!|�ym��Q�L��|ze�vO��4�= 6�f��BfW,��(�U3gFf�;&�e�WP�������;�Tl��ܼ+)�画x#c��z�K������,f��"�+v��n���]�ŏ��W6���]ZGJ�ht�&�ww�i`��TzRJ���|v��y��n��������4o�G���=[DYa������������'(V��v�Ӛ���p��Z*4cz����F���H��DO��]��sQ���)��ӥq`Mz���g&��G��n̻˩�J���c��c��_e��ŋ�I�s QX]��hLj���lukdH
z�R�ڕ�صØ�N�
�]�*��T	��d�U�q�8�����sɹviݖ�q���t��Ge�}L�g3_S��_�ꀱ���߻^�n\.\���@�ؤ�#�b65Dc{��K,�r��oJ��הQi6�]s�D�$a4I"MH����,��v}7Ow���D���n��Q��B{�#{�);�bu�e�1wWDY(�٤|���K|�{�쌔I��DܷRa75̡��]$�]�w	��dD׻�n݀
�s�Lch�F-�K�%A�6;�7�{�r&[�h����Ch�˕�y��qh}��t�G6��Ѯ]�;�����k�đ��Ǒ����9�*�����+W�s^c���Tn���+sW-�߻k���O���ʍi7��-��F*�bך��ԕ�hѵ,h�5sE�U�^h��ʹZ1��#lo-�F��~wU}7+%EF؈ՍRm|Uʾ��s��nmW-r��Tkⷚ�6�k������߷����7�ї�S��?>4�H#\y��	m�!���B�Ca�늁����$���Bgb���;�N�U�x��A/�V�BS|Ƃ.�}���A���Ԃ��[���O�UN���z�V*z�uF�F���`/F� �]n��]�!2:2PeX e�@u�qM��"]�B�����V�*�B\�kZ��ϛO\i���PD6ץ�%r�l^�F^�N���8��w�l�X�A��m�����n!އ��Yв�w�_! ���&z"�{v�e����Ј!���QMRUVt�"��^ �z���"�"	m�����#6���j���:�[�Cyy����O�p�!��m��*�y�a�/�w*̸�#�G73��
(��gs9e�t�@��Iӕ��%+=�R���-���f�	Dw�B�C����Y;��M9��w��4�.Ɗ����ԎN�D�J��I0������x
�n��P�� ��jHn��ۑ �M�`�C��Vh�L�2��L�}`��y�
!�3�A�1fr��هF��a:`���l
P����6�z�L�fd��ʏa����A�/KmJ�δk)�q�5�21w�����,��������Cp�$���NQ�)Rt���ϷE:
��ǣ�y��Y�dp/�O� f��q�WN��L"�T�:��:�܉-����X����T���7=�{����fx���_B�m�����R��r�.�����8���s�)�|q{��F.^{ ;�M�j"�^nuT��/������An�D6�̡^ˉ��m���>����в�dp �ؽ9� [�%��<����2�=��o^�g� sQ�\�4eۋ5���rX�oJ]}�lT�2�NtyN+d+#N��ݚ�:��>�>�oqKB창n�T�n��H�q5D�k���dl,G	B ���t���G���j�B�C8liM�T�j�.t�7n���*���vM�X�݋h[+e3Q�j���6h��`u�!,�e�*�� �8��6��P��2h��,�[tT����&�f���H;Wp� �JB`M��"��6��*�X��_���K�ߺ�u���Jg^Ai�ZL9�M)q@M	FJG',��7U�fA����[��qdН�7S����Z�s��6D��}��^�]�5>n-���״peu]̎��������3y����1@��#5�77����@����2�8D���m���g��p�|���Z���X�8�{qO�#5��"	m�!����N��p(�3nD�p���A������.����Ј2�׺�5p0��}>#5y��	m� ��-���뎠�%�=2�]cw%Nv����1p@�����	-��#E[V�X�{K!DM	�d$"U�4ֶ�T�\�Ԯ	Bd[&�l�� 6*&R�������mϧ��P;���/������8�kx�~��t�頋�DmIǛ�@��ס��w�G�R�o�C�t�饋�O	��̐�F��4mw�5����h��s	<��;��m3kB�m��ג����ܹu�+6G�������A���bz��ɬ����/PD6��큑M�w� j�f�$7� |�Rč�o�U�t�k�)�*�����5Ȓ�"�h݉�u\��ɘ�ւf���
8��t�F�o���������$P�\�gn�h�uN�RCi[�� 6�H-ƕ�]�kW�+�?e��l1;�d�x��H%�yy�r'�ό�������w��nYh�[V�f�X�� ��&�5�z�͠��mXŻ�mV�o�9��w����A8ڛ��Kz]�9�ͥCy�Q��35i�:�ɴ!� H%�DlF��m��q�J�fŐ������+/8�
�o�L)���^��-�^��T�vqp�!�Ԃ9�	ހnD��[C��	*8��{rb�d��&)��p��:!0`R\|ҩ'۵Q7Q*�t_Ns��5m亿OpV�s+��v O��k{����X��+�{ʶB��g�?>�Az�6�||�Ÿ@������9G��5� _B �mZ�����x箖mM\��}N���y4��H<�{P^!�>	n�>mm�0L�I��&r~c�j{��*�o�L)�� �j��5[�A��M�3�p\_?���F�T������ڂ�mH"lݦ�Q�j孉#]�Ad���Sb�W��/FvȐ[�ktVQ� t�n���I�K���f��q��F�O��6�-Ǒm�"�粦���U.p��رq�k����j*�{��y�In
� 8��o:t��Ax�v��� �����|@m�]�W�]ӱ��k0�o^�SI�x�k�{6��yڟ�	0{{o,i��_@��ѫ�u�(� t�I��5$I�Fz�_B�.����i�`�!��l#o��҅t�ƈɂ����d` ��
�Tm�]��$iG�Te�_a�z�Ӎ���9C�Gc^��y�����q��ud�ˈO��ml�}5�{x��c�C	}E� �M����(�|,�?>}��n�fP�����!A�q�\PnɰZ�D)�eLL̠�?H&���s�A����!��z!U'��G!W���˕c�UǷb�|�^n�� D��J��߸������z�r��ND��.�>�=Am�v:�n�� )��z����-��ڈ1��#�������=���hb����/Zp�-��m̊U����H�3���A GoH�7
Zf��Z���URq���O����(��m�3P�';T�Ay�Cn|�kb�=�u�R��Ֆ�h��ʫ�J^�A�/s>>mM�$��b=�ӂ8����vLqD��UJz��^�\tPT�]H���'���o)�<�9�̠��c�|]�Ä�{��\ك
.��E��&�t�h7"2�m�W�T���04�i+�pQ#eŹ�h�R�&*BWA����f5��T0˩�W,{�m\�.��z��9ޘm���i!
F�1�LS::�Pu���zǉE��4̫*.�U����E��A���K�jb(W][JZ� �͵MK�X]�Xl%�G�0�!�����R�"�fSA�X�����߶K&!�#,�۳4�l����1x.ʰi�-��%��_��_�@�ϻ��4^-ǐ8ڛJ�{�����)�SC!urWȾٌ��k�_�A�7A�,���e�]	#��O�rJ�-���ʼ�j����H9�/��w���/�RGr@��CƄ��"�S�UGF��7Nb0��eU����@�7P��A�"�	�^T�q�j�#u����b�ytU�o�N�M]�����Z��ݬ�R����o! F��r$�y�Cod����q�x���g8�v��y��-� ��RA�^n(���T.�e��[��`�U ���h��5���3��%f!�\��WY���F�+d@�=1�[�!�'D�G3x�;�fM_�O	Jz�PD!���ڂot�>>m[�jȟ<�g��W4M� j-ik[o��7��!�TPs�j<��p����C�Z������2�fU�s����N.0�A��?�>9�"	��R..�>�o_Z������ք��d��/�� �9��}�M�v'Ŵ'j#9���Ό͌n%e��5+c���I5��#�ڟ�L�e��a�Sװ4/�	�"m:*29�h�u�d��ġ�/a(�G*����5�:�JC�H#�H� [�A���A�e��Aݵ��r3�^>�[t�b��/� A�D�����Sˏy������MpA.����H(!f�Ls�,nI+�:�%���1%B��͌���B�mϧ��U9��b�f+/��[Gz�YI_�r��!x�ā9��ۙ�9������|3PB��b����ɻ����"7`/�S��%��VǕG��j�p,� 6�R�X�7�S�%����.j=�����.۶i��:�|u���ѣ�h���*9�u����y�,��x�\q�I��V~��N*����˝�T#>����#5Ȑ[�!�nčm���/5u^�D����T洳'�8���r�lp ��b�}JL��jb]y�{�כ�e�|ۑ%���
=�S�6,jAy��������d��ġ����umȟ7�%w���~��ˬ�@���YYTs���r�%[���SWY��G�۳o������|���z�m�{�m��ӛ��JD\j��:r�@�A��"h Cm	�^"Ў�GD��s>=�VO8Wn�V_h9R�8A��$h"�_d��[��>��T�X���-��q`��л��Q²r���ܜ���C�݄Au ۹�p�[�+Ⱦ[����TA�Gv ��R..�����ۗ��0�c�½t�M��f�/�Ҟ{,n�9�@��z*XkK��qv�fB1c���.1�`x������7�w_]��U�S�ނx[��5�}}�>�Do �mτ�[��m �ȋ�?��{����-�;U����[}݊A�/�����Y��K�Gi&D�+�ً�(v��ɂ�;r]u!YH�H,[ٸ�R�y��P ���D�U=�q�V��eN_�O	Q�]�y(�Ta�#��|Ch/�6ת�gS����@�r����ټ���}[iH�� N�A�r$�jGn�*���]��6<�AkӍ
��KF�ݾ�S����<�7R�;�݊|A� p�>���6�l9E�� ���I݄n
t����[7ت�/�.��@�I�EH��60��^݁`����^��E�QW�$uJ__�����7�\��OE�᥂�{�3dI��7 ���X��\��C���D��w��ÉO'�2�Nc��﬚_m:r�}y���"@v�i|�A�أ�����t���[�VF{��a��36��H�[�A����*��N�qne����M��`�e�F0̾�M
e�u�Q���zqf�1�7Fʧ ��v��r�*i{Y�v�T^Jy)s٪��j��3%#V������w���>�^��C-)�(o(���Э���U���/�+*�L;�D�2�n��k�{�#k6eX׍B��;��b/\���#�]�A��^�f;�̨��JN�Z�|���$�J�ؚr���Ӷ�7s|rKݹ#^LvQd�y�4�Xy�5�m��U���tـ�Ԗ9f��&>7�eL�P�P�+A\�{o-�Ý�����NŞC+ޣ�+yimh����1S��p__YEa���2	�۟w|�C(�u}Y(\�]�A23�+L�d�ز_;��L8n��d��FtȻ-^�uCS�/_�!��-��ܸl��r�ը�,u&���"7]�:��ꁥ��X��`gX�:�{,e֤��nww�K�]�!Qa\��D�AJ��S�&��-��=m��{#}��u�nu��W�\�x��q��c���s�8�V��
�<2�Mq�;�(][�ؽ�W^�#���,4,�A���q��^5LR,�-b��SCڽ��X����6g`��6�(HꝖNIŤ��k���Rڻ�6��5�`���n����Nmwb��(=��c?>����~ͮTj�m�����5������b����h�+�slV�f�$��i�cZ5��{��_>uX�4F6��y���7�U�k^h#Q���hأ$5_J�h(�}���cF�Qj$��k��Wc|m��OκUߊ�(�-�Z���Fwn��m�Z��r��6�����}[�o(��Õ�%�={B^sL�.k���1��rۛ(���W��ԛ��-!�[��_��~�v�)��c	��vG$��S��b��iF�R�B��Cg@얖�1��C�],]�a0ڰ)�aJ%^8�L�\���5��mT,e��R���"_ �,R�͔k�^%����J鳬b���)��y�F:�=@�m-�,�rb���*��i�sc����ns��|I��i�H�]�-e�]lD.�Y`
1A�H� �k��u�Ln���u5��)3cUf�����[��E[Z�:����+���p�Ve�)�6�]�]��J`���ui���YU�@#EbSIYU��G����2���Dr��S �-�gY�;n� �62����u��v�PX�Hl�s��ii�*�ұ��x�Mq�]�jiLm�%],bP6���i�b��b)���Z��0�ʌK^��X� � 4F�ۑ�s4Qhhۓil�Xd�X�5a̎���9����Φ��P6�"+�1�j��,uV3MH��A�	e�R���׉�e���:��b]3p�X�p�qcEn���K3���b�I.hܖ6��ͼ`R��!���ek��b���Y]��m�F�[����SYcXX�S���+�m�T�6�F�Jd��F���u�6�v����X�v�V9�ك�B����dݨfdt��̀��ef��C��k���ktvW`bSl�b�[����])��p�^V����ڄea�^�!m�v!%�h�%+a��%h�V�����IpBU�Ýa-�,0$���sQو�cG\���)�Xr�=vX��ՉJ;�[���+z��P�:-v&K��D��t�+�*e

��\�֍���h�G�5و�kJmC-�kV�3:k�1m���k 6�l(JZ����2����9�`2]�j;M�l��v4��&�h��$i�2�0�f�QQs�+r�*����.4��#ZU����f��Վo;Pf����o�ߑ��/��7����cW��C�M�7ml��l�s)�J��f�ܭ�&�f։�t���{h�������ն;de�9�`unM-Bd�)SF��jl��loQf�ucrhD�����uHK5��m�����R<�ڍ�6�����S���[�&8a���pb�f��*Z��hb�R�c��4���4��x�87~~~��A��&bk�]�;GYu,E�u)-�8�aJhՙ��]���y�{�f'�ngŴ�����o�y�r�lp"���sc�ua�VAh {��ڒA[������x�r���A�r	V��΅?2����5u~��p�W[��y�#���X�A]�{�m��yx��Tg��J����]��jT���y�O�p�-�w!�8en#�&c_�<�Dv����������%�w�r�l{���$�����U�2��^>��A�-�@@mȑ��p�ʄ�fZҾ�̧��E��y%���<A�#v m�����lQ8rE�r�G�����u��`�驌X�swX�r������Ih-%�*eMڌ>��$>Ax�6ԋ��؞.�%���W��um����ϻ��-�w �� Ft�ݎ��Y�ݒ�͈_m�}�P��C���򂏷kj�hҲy�%�}G4� h�ӲǑ:7s֖��x��,;����~�G�#���܂w��m^˧��r�lp ��RAZŸ�bG\Q�RF4'\�mϛ�[h[%t%*-���^vR���Y~P�A�Z۟	���p�
��)���^́�9��A��^��kʵ[�V�)\��˔3)m!~v<�P��7M�yݳt�m\ڸ
�Z�po-��t���[ N����h [�j�M���i�v]�ͼA�xn� �3]R��n��8[)Īm��KH'm�<��nV~_S@~Y����-� ��U;��s]u�T���p�Ǳ�nn���+c�eVEk�@��|[A�"-�$.��.!s��S~{ ��"�&�^U��M�l�Ȋ� OtA�>n6��vi���b_!�{�`;�"7`/s���hJ#�D�����}no��ܚVcǻ=xnOw+�VnuѮlή�ƺv��{VF��Q�y��1�q	nX̸�ܜkR�r� ��?�=�q�Y��mr9R�>�ܧ�k��[�j�m qFP� W�"��c�!��.:�r���r�RC�{cǷ�d@Q5S�u9��-��������E����dd_W��w[s�{}��z�q��B����$��������S5���E*t2cC75-�yF�J��8��X��
��l�������}[�s��m����wc4��e�[�P�V� A�7w��>^�U�w@��� � E��sY{M�ձ@�B#\	ۊ]w�Y]}Su9~)t�� A��ndOl�>Q�D�o{&�G: ��r�mq�[k����&`^��vV��˧9�&E��x�36|�X ��m܌��ۨ{]�/c�>�A�ץ����j�����=�`�s�W.Ͻ2Nh�^-��'�2�dI��<����vU���λ�`<�Q�RR�#7���f�<#j>'y5�=>məw��>�|�G_�@!���n ��[���f;������@^l\_�����WU��H%�{\ �b||��6��
�^�꣆TȄ�FI�(eKned
�b��-fD�P6Rn�E��=�.���_z��^�S{��y�ݖ�sg&E�	<⩱�/3�21���C��op`f���n=]#$��G�H"�H���]��Y}9t��Q�)�A��$����;o4��E�VR�ڐ �@6�In��`��I4z��ie��WU���� �����ŸG�{��nz;���@�D[j}{��3�vu�W�.�Z�	E�Jꉅ��AF�u��=��D6�H%�D7 6��gz���H+ݭ=T�qf�ꅷ)�=|��f��-Ǒm�6�N/#�3�(�-u�8F���dR��m���SDQƠ嵳�� b��Yx�3D��2,��A�]{L�k��0�73� 쾫b\�9u�3x�S]A4V��A�a�T��sZ��aZ�hGX��k�5#�KA�%D��IQC#��b��^x"��2���J�!�Q[q�t�mBL��z��͔�%�4���
��#rZ�R�1&�Z$*��],p����e1\�`�k�Vܙ8�0�M9)n�e]n�Ѽ�7jD��!Q�5SKA�
��j����~z��hO�
4Y���ҭ��5�V��9��nTW,ҼĶ��,[ٸýO����@^ �{"|[�n�=f����W9Y~2�BG��4�kP\"��z��^gt��my��	x����Z�#5{��7�^�_e��wY�ԋ\��"3Z[���%8qeU���w2/c�6�!�3�C0X��9hGF]�:��śۈ��N;��ا�����D�RCi	��fV�U�x��
#q�=� ����ೲ��d�e�����TN�wmkɀ��ɟ=A� |�Rn-�옛����)��ηܓ�ʽN�b����������h>�a����/��k}`�:�a�\��P�"�L�P�SE�%�#���]Y��U���O��.�'�@6�|�*��>�Y���ە��̜���QxQ����jAv��8D�RF4%�y=2���nn����Wtۗ�
�	�d�W\�X�^԰�¾Sf�h}������<���3UD֝��.pX77=)�X�.�E��ފ���ߠ!T~��B��ޥ�����x�� �A۪�x�_vfߤ�}<�/�|>R-�7�	m���ٚ���i�{��=��vө����"An<������麷�kkdEla�H"9����M޺���}��w+#�'��WTL= �V�^M`�(��8�H6�〈>mȒ�Q���`�
�t�"��tF\�ߊ��Olyf��Cmz[B����\0��!"� L�J0�����%ԓi0[b�,K����e����./��>z��|��@���Uf��{BݬN�R#8 ���{7ͧN�k�qǓh"r$�z2�u�pa�`
�����W[�T�e���Ee�L{�v) �k���ɴ.ĵz���Z�K۰ ��O�n<��cg��o>��z���uB��kCT��d����]�:x��b����X԰�Z5�v��"�A��"fj%j�������$ok��5���r��O��l"h C�>��^-�9S�k2�m�@�A����n�лk���D8{���Zu�
��nF���m�7 6�!�92��O>0�r�󨧹k7�Yr� u���-� �����ccE����>�g�4��ᚆ@��Kk�����vf�kF\Y�:��)#��V�g�g��b|�����h*=}U��&^]yD��̆�_lw8�5�6�^gj��@��mI
��nE!��@�s5]�ݽ�I�d;�N�C� Ot�hIn�<�y�";�	=��6�m���<K5깣r��\�/H���X#̃�����u��� �Ԑ�	��}1==U��F�O�����
�y��uwaR���9�����'�Q�y�}���'%�W��	�e�F�Μ�#�M�5e]��9@Z�+K��g/���Tٵ�S���э�陟��{�����/��Ŷ�>mq����9ke\7aDX�ͽ��{W��Ԉp;Ǻ �qȒ� A�n�I
�����7Ҧ��!�s��aH�;9
V����+5�;6�caM��_��w?.�u��m��������+\�`��K#�1����Q�k<�G�>m�7h�
�
[%�ڪ����m
��p����4����A��,h�ȓR�p��r�� �uǐ9����-��Ŷ��Vo{eKݨo��2mmH���F�"An6���� ��0]�;�p�FdFn�7&z٪�X��e�����v)#�.���<���� ��{yI�@�q�[�b�w!�N�]�6)ź�WMwa�wu�2��D�^6�|Chg�=L��=6j$NG!K![����A9Ǫ�U�ƫ�d���st��_Q��e�)a�Syi�p��F]-{7��]"���AB�HY��[Xka�I��P���4���\*VX�K���i����cw���&眳���,��+mظaڥ�C0��=�a*�,�]eX2��#�b��t�R��l�(m���Z��M��(S3M�pislÈ%�C�yx�!���4�h�4�fm�@3YK�3�,�ƣ,/gH6�7$\YQ�̪�R.K����~��ii�D����84�i�� �ʣ��`�#���nZ|��	���p,�	m�O.{Fgf�ù��"?W^��={���	 ���>8�x���r	n=�`�ރsW�v88���zy�[��s��z��̭� ��R:�@�*��91���jAǷ���n��k�'�fP������3N�<�<{� AmCngŵ��!V��_l'�+!��yڑr�;l����mmH������A�H&��`5Ј>�Ax��ϛ�A�h"zL4���myof+�7S�F.elq�^��[�A���[w��f�������j�0[ZX@R��lh�ű)k �TW侽��ő��2=�d��pt9ݥ8�	h�K�D�@��z�fob0gP@�{>����ڒ;0���u=]�W�)����aJx�K0b��U���cu5zqn��.�ʷ�S5�4��IIbh!0M����Vm�����=uw��i�1�y׷0�Zڑ�{� A�D��5��&L�00ۙ�n6�||�eL]����,̬깊�m���*�V@����^-�[jHm!�fU���		�� �^m(]��<6z��*�ϔ���p"�t��5�����&4	����4n�Ԑ���h�C���Wd�[��iP��΍�}}s��Ԉ���П�|C<�=�*�W.��(�F k+SM��v]iR-pd�i��v�fgeʺ>��!���O�(�����+�힛����W3�Cɻ�9dS�Ε�}z�vŶ��[��ٖ��kX�fƃW���ww�����ji��fP���3P@���Q����1<i ��#�z�Ch [� [k<>��7{V}"���%��
j�Zܔ[���@0�P���������ED�T�6bᏥ�P	��(��*�2r����tѕړ�f�q�{H�ډ3
7�eN֨ݬ%B�Rt,X+�WN\[��YS�,��6�)6���֠�u�1+HU���r	�5w�3C��!�x�\�����p����A���������LtWY�-EM���s�]P'.���Y��REռ��u�v�i�(�P�4����ܫ�,uv3�gD�b�B('a�<wS+0��1��¶5�o;��__k�rE��);W�pX��B$6d�*I��(�sM�����#P��#Q�5�A���1!I��E^����*H�p7F�v��Y���X8�Q�y}��+
wP�HN�A�A��E�5�^�;v�	ً�Ԃb,��ݑԡᦲ�˒�쓲��,u����pd7���Ռ��i0lفY����w1u�۶s<6��ˢr�9�qlɮO�SՎ�X�u��BkJTjl�U���Ӧ6;cL�Un��Gܖ����ݟ��d����[��}@EbB����Y��[n*h\����Uo!�,�M�x�E�֎<����6��`�\��ms#.���lѬ���6��
YW� ���I��t��� #lP���b��;�2�v;%Ð���p�}h�)�wY�g�j�X��甕��.�R��n�����.�I�\C�[I,g�nAϭr�ף8j�e����5�r6�V��/
�J�/!
!��Q�[��^ksA�*w[��\�ݮm���5ƨ(�5�6����[r�E�|]ݺk��ysd������kEy���|n[�r����U�E�%_M���`��]ݯ5�o�弢��ռ�T�P\�,��d�Kѣo/�{65��r��*4D��n1E%�\���6���F�>;&�&�Ͼ�6(��o�W4n](��
 �4U��J��F�B`��ݙ�x�b�ڑ{��>n=a����]�����A E�^��+�ս6�[��e\�Lq�b�w�v���I����N�RCh An ���p*F���.����f�Xyw���ȵ4�}3= ��C5 ۱>!�8�!=/��7֋�%����R�9�X�#ms,U�����ae��$R�S=}�Ԑ|���yx�Ԋ��վ���h۩�6/p$�������p�A�h/۟	�:k��wj����3����/+��6�[��e\�L�k�Aւ-�XU�}
��)�X�]Ғ/�/��6В�"�h��Qڷ��L�3��=|�*�Ϧg���<�P@��ϛ��n=��s��f��'�Wy�@�[jEc�O��꺺h�̈�_@�nMF����XO2��5���W��{,�~�K��n��[{x�6xrq�j�i_4��� P{{�Qf�ޭ�p�4���q�,�8��Am ۱>n �h Cnm����G��/�n�;f����vU̬� ��R��"-��ܞd�7�j���`�d�H��RB* �Eu�`�uXgkll4�j�(M��!���Ϸ���n�nȐq��P����z�\];�L�_e�ʾ��A�4������q@����O,Tŧ�In �z����9��g���5�"7���7\��Q{�E]�눪�qGc�	Ƕ<����Oۢ�t��y�����=�����NA���Rh"�"	m�6�"nF�7�+��p8��BA{��!B��hk�_M�ӹ�� ���H��8��M���g�ݨ q�m�Kh"�$���U��/Gr��9��Y��rѭ��>;�\��n ��_(|3n�q���3g&��&b�%��cUG�5Y9�*v�(I����xbӠww�E��Ns9��S_n����%fe��:��~"f�&����KBʸ�, ��P������H�fS&�P]�n��\�f��LV��Ҏ G*��-���d���A�:�rk� ;`�E����qa��C�6�L�º��i����!��љ��Ye�L�ں�
�:(�K�ر�^f!]cqMh��K,�y9c����KL�(�ňGa]3��е������!�9�긷^�a��bV��M�II��:k�L�v��v�{'���F���m��3z6�\syq72�q�;��31�n&$�-��ͅ�-�$6��pvb�,��25B��s+�_MEӹ���t A��!�#:��֭z�=@�j�Cp-� ��M�m�.��z��w0ֽʺh�̈���w\�-ǐm ۹v�+z��c�nL0AH"j�p,Uq�q��y��M̧A;ؤ����[�� kaA��A�@�mȐ[�%���V�(�'cvitth�ۨ�w>S(q�-h"r'Ŵ�{ٺ���[W��F,�P!3f�<��P�,ƻ.A�v��u#O����)�9 t�d���y�Sm�}--�w6½�#yy���M�{ò�܉9��n m�7�q:���qR�z�b���Q��6+xcr�A��+�RrJ�-[9oh�T�!R\���K��W9Xٮ�������LA[�͞�̉�)�	�� �9��q��;��.U�6W���;��"An ��;�d�L�i�S�#a�ͺ��s�3�A���k�A [�FctM�/bV*�٨ wc�ڗ���iw7j�W��o N�F�_EB�;1G�g ��	n�!�!����[3»��	0�A�	W8�ֶy�a�T�{��)h"� A ��M?x"�d�0e��8A�8/0Քc4��k(��ך�v���̤��V1�7w�}�����dH-� �hP�t�p�ۨ�w>S(4�P;qA��b|@m�� |�RA#����2t
�#���x��]��-�{HF�@�w`!�7Z[�d2n�B�u1܉�8D��s���|�'c�8v��S~e=U���R?1*K{$�R�أ��C�̅��Wt�Yh�E�f�mp��N�/��Ȳ�q��m�rhJ��ݾ؝��8��RA�E�DڐCpLV����Ȑ^��
�M�=��g]Eӹ�̡��B=�����;�y��^>m�7�pQ鍢|wV{u�|ծ�y����۰�zА[�A�h]�o��������S�ƕ݁7V˂8(�e)�Ԏ�h�E��14�-�#��gm�|��K/�B �@6�O��F�,��vU�j��#C�����P�Mr�AkݱD�RCh��/-��7GGwv�\/sPB�M�]��geEӹ��������o�uɭ���@�Bל�������'�idc��:mns�a��@���;�n��� A�mCnD�����7<�2��b|[A+������}�eZ�� �݊Av��e�@[gJ.�zo=�*�͛�]vC�T�T�\[�
�#�w�r��y�H�Cl�����+���SO����W�3��yO�n��B|[�|H�U�c9�J�::��]:�L�H'�kAۑ>-�LON��E�!%�$������u\ڛ�)���a�&�--�YG;>������n�%��6��k���ֳ�P�K3�-bz��FE;�o���y�@�܉��a�� "��Bv�s���<��6{.J�i�x�v/O4n6k��=g���;R�mȒ�y��{�}�JhD��4�N3{..�Ϧg�{���Q��7�;T�B�U���y79<����9��m=:��y���ֳ�P�����]����u�q���!�"A�D6�m�5�ٸz�F�`1��zZ��[�H�V�{��� �pn��j��ׯ��Ra����3V�5on(��dɤE۸}:+1�LA���PȉZ2L0T�C^8,�̓�ɴ�����g�����Et��2�e�wk5iN�B�emmjF�p<CQ�cXL�K2��#�f��]��W�e�P��8��ۦ���Ql��A�j+0�4�ZKG)��Uت�h��2(�W$#a�l��	���eP�4z�l�%�%4[�V	�4q.�JhX��0�WG3!2$`Z.��A�*޲�����������2+M��ܶ�՛��=�]>��R��Д�-Pل�TS[����X����h"7U�Y�9z\A�vȒ� Am
"b�Oq͗y3��Hx��d��B��=��^#;���A�"��ڈ{9�#����v4�^jni��q�{n�ځ�w`"7Z[�}'UU�(`h
�$��h/ۑ> 6�LV���M�c;��ӵ۔���Ǹ�^��y����v�M�j
f���� �ݟvŐCh*B��OqΗj�W�g�{�x������؍��7�'��"�"-���h/�֤!�Ui��i��r���y{����ཻ�r$�y������Rк��peA&ɻ��D��^+6�]+�
�j�h���+�Xc�*��p.�>���ϣ,�Z�܉�m��͊��[ΑT�8��AZ+��WJ�; #��mI��n)��7����N8�������ڌ��>Ǧf�Ȩ�V�
��o��X���nĘ���U�XӪf 僶�a[��ü���1Kؽ��&k)� �h*4c�yt_K�y+�2���f��!��W�i�o5ɠ,��Ƞ}���Ap��iĮS9�}5p�D�+�;W�t;��� ��D�>n,���6�HX�����Q[#)��O�m\�͛����RU&�p ��^���M��9�a���T����p�-���O1�<�ygv ��v�7;�E��W��3<�{�x�p�|[@�9��*��"�3���&��m�
Z0Kb�ع@#3��[,�p;�H&s��s^n(Am�.�<�=9G8;����w�Ulw@X��{������y<��
"��Kh ��۩콾w%Rnc�{�IsA��Je�N�0guI�/n��������7�#��3Sm{�1(ī&�L����PY�N�ц��f��]f��--���2t�i�_��X�YkB�q��i�ڽB�N�/��p�Ğ�A�̀�Cng��E�D[�3wy�q��E) ��͏ [jFM6�_�G89��#x NlR*����4��sAx���A-��@�ب���U�^���{'���ͼ�tU&�;��^�sA���wk'wdU����"��v��:ۙ��� MFlչ���t�C(Z�݅�����������A�"An ������=�7��^J�̡݌dػ��� �Fk�	�mp��mI�w�.��j�	���2헗���7��o �9�ۮD��Bڈ""�6�Z�#û�@�Ax�����75t��\�dTSg'��u�k�*�sA=ؤ9�E��-�>!�<�K�̈����|�H-�!�47�oM�W��3= ���G��nq݊�+.z�)NeO��0DN�
�S�1.0�T1�8�r��n6˝�Ƨ�{l'J� �oD�=��佉���0q��|��QŶ� 6�8�3�0r�۸qٶy\��̈�@�����H-�7��:����=辡���E�e�FZѴKwR%ʸ���k�f��˘�*�y�����>|Aۙ�pT�9�S��3��Rnc�&Y���Aּ�+�mH!�����M��~�n���7�1^R����{�j��r�/!9s�7�\��A �$כ�[i��mӊ��+�u����.�ȍ��6#u� ��� CnD�'����]1��X�or���
�����u��f)70�!�TF3���@���!���p|3"9w;��B��7�X��3�T���Jڃz�FkZ��5�}���տ��_�뜢,�:i	K���D�B_��	X��K�P�昘�C�T&eN�¤�<��5GҒ�J��2�bH L$��Z�TmV����Q���H B����BIa�h@�� HMa��i�!���&i�����1@xMVT?(aD%�~��jZ�K�17��ĭ��M��ߡ�tG�$6�@�J�XXe$=��M(����z���BB|l �e_[�%�D@I�F��A�$$B_�?���S�������IhA�$$B_�ZB!	��`��!)=����������Y����������ܿ�>!���}�I����!����~��������14���Hm�hR X=����)��	��B���DGا)&��sRG�~��!�������$ Bkg�������K�+#I$���t|�
���m��@I��i��	|W�#��.��
��$ B�(Ym��żڃ�=g�^y����"%���B�`<��4z��#KԿ� ?�:a~�|O� ��O�>�{�_�?�B�K@qH�`~��5����|>�?�&J?k<�>��\	?/�����3�}���x�XB���=��C�'�K�����'�=Gڄ B��4�=�?h�0��<`[[�F�� @�#ݰP5�^BB��>�!��G����f�ľ�	��RY�@��I-��0� ^F@Y<�H�%���cm6��.*Gꄓ�l^I�!$�!(K%��z�`e,_K9O�30� 0>�z��L����Hb�(�V�0Rڐo���I���>��i�]{>�!��C�� ���� ��/��/������K�z����/@R �?`z�����c	�����=����%?z=I�=g�m���B�K�>+�����A ���������B!(K��g�jO���@�X|��萤���뀴d�4�a(g�񂆘�P��pj�L}��A����CK���޿��o����4+\CU�,�������W��{�<������h g�Xyz!y��}M0�׻1�ف���E�è�0M! B��M%�	���l}O�g��W�^�D$����	$!|��`�hih
 �=��CO!	-�A�O�P|�pe#��0bG�� ��	����b�H�
26 