BZh91AY&SY"���X߀`q���#� ����b"�                                        P)�  @   
    ( Q@@    
      U   
�      x�	R�$)ERU*� RT�UQ@�UU(QUA%E(�R�R���R*IUQU�   3Q����%% |�(n�((�*]�T��:�I��%\�;uUT95Q��n�Ф�"@�@���9�>��  � ���;f��D���j���Ч��T�%*��3���dR�սq�Rzҕ\� r� L�*��Ð�^�r t��� K�  ��P��*�R*�E Z�U� ��U��`�� �c� 8��*� lǪ� ����;���{ ��<%�l<�@���  � '�� �w�= �s�H� a������{ ^�=���J�0tu�^��  � ���`׀(
 �  /�>IP��TH�B�� m����:hDr \H� �t r w`�� kuQJ`:�@�=z�@ �  0<�G� b�

�f�2 r �rLtQL:u� �@�`0� ��|  }(�$*�UIJ 
D��z ;�9� :��A9�B��� b����:K�ҩ�G ��   �/�  �{� }� u�*�����w`� 0u@���u��� ���X@ _    �Ԓ�*�T	 �P%Rp�� � 4��� j�J�. ": d�ݝP�� 1ܠ��@�2 �� QBx   `����u�8%\ 6��v 2 �� 1������݁���� x       O )TML �0FɀO���T�4h h h D�2�Q�I�      4�*H�)H�`��#L�%?R���F�@ d�CL@ R��iJ&	�3$ڣ�̣MS�&��g��a�����<�?�G�|���s�a~_5�� �����PE�DO�E�����g�9UE3���GG�?���>���>��l��j�������UU���
+�0v?�B}B�����������C�@������r����?} '�EW�S��������U�m�@6ʪ�P�PCl�L 	�T� .� �(�v��`v��l!��6ța�&�Cl��]2�dM�&�Cl��m�6ț`M�&��v�;`���Sl)��m�6`X]���Gl��A�"�~2��a��vțeM�&�Sl���
m�� L#���t˶ 6ʻa>2&��"m�60&�Sl)�D�',�T�"m�6ʛaM���� �6�p��6�;e���Sl���v�&�l��T�*m�6�;`���l�ef� �v�;d��P� m�;`�m�8a���l	��m�6��`M��2�1�6�a���l!�D� ���
)2!�Q�� _��/� vª�@6�Q������$Tv���]� ��!v�탶Gl���A�(#� Dv���"��l ��`?��6ug����h���gvM����T����y�.32��7�f��ti�ьnN��� ݜ����͇���,���oP!��7	�uD81.�<�T��<:��K3l;�gP�+�q9z�{/�dP�� ��_����\�[���Ų��Ϋ���E�Yݫx@^��>�kU8���i���BG��Sk��qm okQm��As�[����(x�Y����\��7t$�j�m�\R��[2W;��g^��Ãsc��T-LD�ٝ�-�ۂ���Ab�
Ц�+��Ow����R�������gdѮ$o3Dgpm<��bqdR�<�Lx)N��s�	���B��������#���d�������m�)l���c;��M��=� ���<۸4Gu�ӣ6�2S�| ��)����`��P���s��]��̋�Όa0���k�Txy��!ݎ@N����p�e��3f���ۇw��ќ"X��}�FmEs�/���Q�,��{w�xrl]�\�Wcl�T9w5	y��"q]�����9 �Y��1�Q��2��0e	V�����>\�md��ׇfm8nͩ�n-��v���Z���ɲweQ���y2i)�}���Ww�<�z��m�?�v�s�ѹId��ۗ-c[9+�yb̓8���,q���u��zŻ��u�p�����ay�Z��^��4��1�� �+��g!ѕY��v��	��f<G�]�_��z�[ü�ŀע��1�-��4�CvM�
��j;9]�H���p����OD�4���`g'4���R!
��wd^	��q凹�'�//^Ԭ����~d��.�%�y[x��f��4�;\10I�;Myp:M�!��.�K����h��ԭ��=<��k����\;p��pV���$Ͱ���sI]�P�k+��NSxuYׅÇ# x�p��1v���o�u��ϋ�w���ұ����^�4�h���Y�]	����%S����ޤ>����k9Zv��6^�/f���,�\[�T��>�L��Sů����7N-W����m�)9l!�n1ǅ�
��i�J�h�e��F��+�v��.�[:�v+���㛫V�K�`�%����[eX8�l9�FޛD0\g�S$�ܴgV��صbݝ���q�`���C��̝�|�=���\ۄS�W�T�.�ݺ�"�n��z,�knu�p�$S����z�ܪk�ͻ5n&7�3/WI���n��@��o|����ɽ,ܼ�K��Yΰ���h�=�GF,�(,�r`f�^�*�P��58D�t���20�Db����'�@{sw�1p�l�(V�<�X�	�ktp���t���y�Aڮޏ3���,Q�h{����b�M0fN êf�7����0`��`!�&����h�����(쥡z�9w
�x�n��n�,ǸN�,��^��zu���G��9M�H����@��/��k;:õ$A�"w�n�z�Y�á�R3�=����5d��ߝ�;9�Y�pǫa�N�$���Sq��yz#�m����p��^l�r�V�{�+��\L�p��hѴ5{�^P�8���!�>\Mۊ��-\���sd��p[WK0!yH����<\�nB�2��;�R���
�XZ@��� ܶ$��1 ([�h�aҗcѻ�Л�3�5-��m�^i[�.*\ڻ:3p��s��)r�N�$��'	&�G�!�<�.=��f��f����$t�{�*Qe�����(xu�t�v�wa1������_p������as��910���:�٨�vNW��7o-�;i�5*P�!yd1\i���Tl�XoA��"�������9�.�'6�;��]Xr��V�N��vf����W: 4���u��3�I�&�q��������$Ŏt�� ���y�&Y��2�p!�a�wUϰ�N��?�Az�;�74��+R���/;�.nH#��=[��Nӥ�x)���:I���x>د1��a컋:��1!f�����j��4�Q�є t%�o6��b������9Mqs�p�8L�8GYxǐR�� ��z��6r��B��j�ug[2�ϹΗS�\�\g�#]`�;�Y�����cz�5�M����{�5��F���x�v���.�O���.�۫7F!zG��M{7��q=3;�!���_R�,���ˉ츜�Z�<�{wvp�� )9�i��͊11gD�r�6������R�JI5����M���z9vh��	}`��ϝ�PDv�jFJ3�]�*]Y�V������6q���zRچ�sG����9^���rS���72�c�ލO�Ī�B���P�BIko'r�PC��ޜwG.���M�c�U����Oc wl��^hd��UӴ*�.A�dɭ�[{�����y��e�|�=/��{�;�d�;{"��c|��'wd�9�+y;�ا)��@=P^��*9��@���v����h�'i�]5�2R�GT�/Gb�Ȏ��Fo]�Ç���rC���h�¡�T�4}�|�՗��o���b��p�˦r��DG4_e4��N՝l�4D�r M[ǲ��5pZ�����ML*sM��Q��N&�9���:^���I�;u�kpm9�j�[.��@\<�����A���a{�S(�w!�=��5�Xi�v�ʫ	��L:����2�pCd5���d��z˖ ;u�݄� q�y�����OpUk����7�����~]�8�0�Ϙח{I�`�uV����0-�v�{~'�ŉ+�R���VN3㼵;s�+^�Y0,�G�`�ڢޘ~/��ݶnެ층���Ƈ[�®v"�5=
.�����ǭ%�{N�7v
�;[��	��"��9a;$�j�=�%88� Y���k�]&3V�<���-��ds�����H:&8���)\�Y��jv�!ybSe`�Y��:�q6�D.���{��r�<��&nh��[�:�<�1e�ө���B�:�Wi��	5pt���n���l�!�QΧ;!����\��4��'���p�"��v�9�V��ͣ-�ޓ��-��>�l�`��Ј���d-ǅ����]J�H���9Iݮ@��ok�v�\su��0\]j�Ѝ�vq���7�s�Ή�g��m���ܳ�c�U٣F��[�r��)(-�����<s�s�S�v��p����p֖���*�M#"L���AMzI�0�!�sx^2�p�n���vw[�ұ��0`�)׺��h]�Fn�iC�ܶ1kr�ٮk���&E�4���c��\�Z��=M�g9iI���N�E۳v�Zj�]}��2F�]����T;VE~7Ǹ��������Cxd�I�:[����r���ߘ���CGyr�m-���`���d�SN藺vh�j�ܓ����J�?[���.u9�5f�͛����b"�׃<qC׫f#�_�4{���OW���qvv�.��Y����5n�pۭ*�f�0�=�&�U����r͈��{;�9٨rކ��v�u_A1�彎�Ң���,U�(t���YF�a���Y���{n&5��vٹ0�ު�K�׵D��U��	���2�[N'o9w;3����z]w�*HzW�ʥ�B>76��\�Z�nvЇ]�"��l]n���j\�L|W�e���ڰ�{�\K7���ac͇���2�N����P<s_
��a�ni�1�t%��(&򤧹oqZZ\ǹ���n��{�D�ŸmYN����n�yj�y�s��
�x�*��Cːea��{�ESe�7����84����=���}��Ո��ՁX�ŝ�uqQ8�D^o{��{��39q��V���x���]J]�.���J�E�t��������g[f�C�١���*8�pz��Ć;"+(�E�Ly���p��eu^\�zY�}�Ǟh�q�,�>o��)��oHJ��Iŝ�)k������1�K�^�0nي0��`�V�V9^�k�z��':���Y��v��_sMwk�����9^���v��3��-}�e8Wa��3�H��:D������X���9�	�Ǟ<�W7�7y�D �ѐg&��J�84�!gGa�rq��m���"��aٜ�0�{*#��dM[�ℨf�Yi�vŵ��s샸[N��ȼ��Ĺ��kh%yn��A<�n��9���S����sP^���n��75�SZ��r�Ю
�f�^���hKw�uR��'��&��� ,�
ǲ�7�(D��-�̀�cw���,�}os�D�m�@��c���Mp\!|m��n��eRܪ��8�+7J�o���Z4�=����5f�wuk�ݚ8ͩ<G��$@i�Y���eu�崻�F��f�q�gyF�}ן�=�fBS�k;�l��N��cҞ������K,隄�7��X�a&�'u�S�e�	�t�iف��< ��mY��\UQi�=�XΗ6��We�؟t�ӻu�S�l8���d�L��=��Mb�ՇQ�W��e��;�<�.�WV�p�1W �{n)�hݻBhǱ/��;�>����B�U��s��q%N3�݁�t�3jf і�٩�u<5��o�ܤ6l�����+�`���Q������[�1��c��*�x�G��;pSD���NZ֬�*A��=�k�7Ew�;s�Yۭ��f��$Yٱ�F����e�V�h�b���GM��n�Öi+;(�n�fuɂ��/�h66�C�����³��voRp��A�cx@�B?T��n��4��o`�;H@���Fq�I2�1�&Wt�$|`��d�؃r:N�%0�sm
�Wlx:կ�gA$ם�v� 6�w�T�o�q ��j�h��ӆ�<��v#;�QQ����B��'cJ��e�*�<omXf�-��!l[>(��P;@��	�.�Z-���� ���B�����@������魧,�t�f��v�Ei6��oj�d���mv���r �����KqC��rc۱��#x]��Z�ٝ�o��\��X�"��a����mS-ܺ)e'��#Ɏ��݉�&�ũ�'���^�f>t4�3G�;���s���#�o&;vb��Z����Yѻ5Z�mv!�Xol����f�[w�;��C��}ݕӗ�6^n'5��@b}eX�Bk�eڄ��ηl�g>5`��3����1�T�O�����"����l�^Y��.\��S��V=83_c�xX�n�;nYH(�3�n8^�]�,;��.�b��v�A� ��ui�I2;�=������ް�J*.��Gsg;�Ր<�ԷFo¾��0�5c���y�+��p�����3od�n��v(3^>��1��go&,��ȥ�q�݌\#p3��n��j��3��2t��P���8~����il���G]��՛ʹs��)�Г��^>x��4�f��r�F���4��������}��w��m�<)9�s��ћ��GdԮ
w�આ*c�{46�T�.3E]�c&;��3�����e;*��,�8�A��f$1m�������$M/�S�N)��8�|uP���LV���M�z�eȻ)�3B����0^�M�)2�\mړ�84h��U������okB�&-�s�ʭ/"�Q���P`��Gy#{ԅ狊a�2u�ޫYK��o
:��ٷ!�7C�;�Z�n�n��+�gP�׽��;��R��9-A��59{r��77;Ԟ=6�:�K�}����"P�r�FrI���I�J�f�:t�����sh]p��[u1T��h�Q�s���P3�����n�H
��q������v�}������7I|N�1�
h�1�&9'o�V��IT�`e�LV,I��BQl��H���WtA7z��Nᮌ8������M�j�JeC�8�����n���ߠ�W;����6ű���bˊ�f�;�Y���w[���t.9�䱎б)�$9���A؆����&�䅮�s�� Y��]N<T����IO,�׺v�& ��Ô���=���͌�o��j-a���%�v�'�<&�܂�>m�ܤN����twh�:um�*���N���:XU��z�/r֟��ۀn�b���6޺���Y�ƄytՏ�nQu����W��+�6c]�t��}�l(6�ݫ/���|�,״��Z肙n\]�X]�ڞ�o�=���܎j���g#����$#�wC�����/`[�ͻgv�Bv��q���ת����Ε�nvX�����]��t{�D��a�6����-˶�9��kQbxf��F�.�M���Z��7U	u��m�.\����=�NYۯ�ӂN�)�R {���a;q�p�(
�vt^ZO������kK���~�:�&�7J�L)���Mi$�);"�a���^�$�1�T��)RX��I�Hiʩ��ӻ����X��Zޅ��{Nwi)�+I���$�ZpL�����̆{��,Jd��Նi%Ib@�&�m.��8wd��F��	c*�������n�����t�N�;�v��+Rϗv�LJ�N	��V��	�,�N��S�zu`�K18���JP���:T�*�WvkK؏{�fm�����Ee^IwR�O��=�����C�P���w�����+{�,JV���J�?�����e�W��{����I�}�g���H��T\�!P(G$@hTJB�J�C �JUJ)EPB�!$�ZV�$Dr\�L��G$�Q)@�( r@2�T�
R�D����2A�Z\�E�F�D)D��R�F�F�
EB��B� ��J
�@��@h�
JU$B���)TL�
D(E)E�R��
P�2D�2@$(��@(hEC!%�)�ArQZE2PP�P)�R��JB�F�(U�UD)T( �T2r@�����L��>������M�^b�fF��;����9W����`�@�D�|�y����9��S���4F� �0�|�
�=07_8��f0�\���;��b "�����~����g�~��������*�����O�z}���x~<}�~|�ɬ?��eoz����k�^��h��5%�ؑ6	�}�x(��k�"�l,��3��zfһ��}�F�ٱnt�5�1�o�I�r��m�Zp9�Ѯ�W4I������.����np��H,H򺽏P���ǩ��=�{j٦�����C��cE���e׀A�]�b�3t�/��^��YA"w��w,�9ǒvA9�<���������{Wp��O��j�� >�|���o���&��>v^����E ��{��w��=i�/��3g�v{EΎ
�/G��#hT@�8困�˴���.�:#f{Q�/M�5�^��u�S���J�t�g���Z��s�i�t��}�&96B
�[8Yܝ�<�]��s��s�t��Y~���[ͱ�fJ);;���fu��١�=��<>��{��s��Rk���t���o{}�l�l�h��Խ�1�Y{1�T�b�Y�@�Ĳl��ћj�_3��F�x�6�)��m���7W08�ZaX`�<7���|���_]h�
{p�Vo}�wg�m*ůج+~5/?h��c$��)ۛ�K���T���{٫FN�lY-wn�5������w�;�XEbhg6j7��4�]��������V��}���*2C�H2��y/]���O��Y��P1a/�����%:;��������Һ�;��i�b���%�^����>}���+��@�U�N���E����ںg��'sX�GÛ�h��Q�S�e�>�oq�t�^U��c�̯dŸ�{�!vL�CfQ��^lr�p��y8���܃�d��C�4w��q�CξK}��{m&�p��`ޣ����M�����{�Ō�n���Q�7�9�;�;�3���E	��n=���{$�)�-3l�s����a}{�k���7���9�	k#��j��K�;;I���<ţ{l�/!�\>��nþv{ �~����NQ�����������6��ˬ��`�8+2�ΨM�^K=��Ҫ�z�t��$��u�{^-լcV�yfÞ�#�z�n���A�B�A��\E���l{�w�tsN�j}�!�z�֝�vg0`�-��n����̗Nʞ?����_5�-����O7"s<v����NM�����Q����_d��r|�{��,��?o���]�x����wwns�^v��p�ڨ=7�â_#R���J����]�M����{w�'���A�>�n�ק���v؃ńi�F:����<S�g.�M=�2�f�o�p�x�m�v-w=���}���<�bC3�Cv�;X�b%����7�>��_�����z闸@F�0�P�$����<��}ރ������!x�=r-oW�tݼ�{gC����k��S�f��c�-6X���������@s��/n���ý��}���m���N4���I��ixQ��'\�����W���ڷ�~3=�]����<��#ν���+pѮ���#|��{���r0�|tb�K9��Ȯl7{w���x���{'&��g��ټޡ�����4v��ٯԎ��s_Zɪ鏀y@da����{m��4�Yn7�@l՞�ۻ���E䇪���۞�|��:����ޔ9�=���|B95X���dx��Opn�5����`�O�*<�vy��hs�+�gc;��G~��ִ��z���ْ������y�]�e�;��0}�^,�B�1��ؼp���[��{�{�h���"=�K>���gZ$���E(y���Y�=����|>>�Yp�힋�M^P�9������&%��fa�Ԟ��=��.xwgM}�c[wpp}n�r�^v}�7�}��ON���+|G�Ѥ��g.J�\hw��6��60�V�C;�D�}���-�݇����y2�-�~V@�[�� P���~8�>.絃��޽�&{=��IZ'sG#��r>�^�U�3����9��m��G�7��۷u�ٮ������z�Z�q�K��x7����|����<X�}�7S}�գ�绬d�G�Q���3Gz��{����TQ���֖M�%��p�rp�C=,�{�QR����ޏz ����i�}�|w�6x�!LC����=���o��r��&��dt�oTȉsց�D7��q�<dI��[~�{��4�яig�Nv��мV�M�Z���h��,>�$,�K/��=/�{ٜ��[���=��!��;UӣC0�8�=����fQfq�'��L|�sVِH���c�f��s��Ʊ��;��Ei$/��<>u���dv.�+4g�˱x�u�1&kM~90��b�܅r#Jg��y4�.�&Y�w�"�xm�C@�H�|C�{ٸ,b}���e^~�'���[��(��#�a�7ޙ�gG��<I�l�)����;�����=�+;�vu�v!�'����f�9���v�>ݔ�r{ۑ�����
���L���X��K�W,�)C�.{lί�cCu���v��&��(�ݣ��>�P��Cq�����]�og<�q5����U���t7��.��˾�
ܩb3����W�ϼ0��L�<;od�÷s��^J�{�\����6-񳃎mD�zt�3���Nz��_���Z�fI��k�+t8S�Y��'b��}��$�z>'{</��p�����4��j~�,����5Ƹ�p�4��qZ����]�-B��x���b�F�ճ�u������Y������m[���p��3H�?p=}�'b��d5��|l�����k��8���?6N<�6m�F�%`��7���W��5�"	���^Ќ�K��ݞw��t�qR��n�,ɠ3r����w�w��{��%Ջ��Ìk��j�<�<<���$� Zs��d�瘯��S}�4w��g'<Vn{�~C��pk����fnx��u��;'{�/q�)���zu�Nq�;{px沷��Y� �A�\f��w��׻ɺ}��<8i�Ǟ���1�:=��Y�b=��ya+�ڧ�a�Q["������g'��y�܊�}�lR)���{��j�{���z��e���s���<�Q�k��q�F"�ދH�:�aÝan�~<�^j쁴�g!؎�l��`�7���ki�N���>��/E�P��n����q;��(k:'�薹�6���@wa�����Ƴ��C�{�b��q����3����#�k����w�E���#�.������8x��#�xFu�v�YҲ����lɩ.����y~Y�o\�=�g0�:�
q�7y�����������<������������=(���'L�{��u��ge�{q���A�����~�0�>�S��}d��5���g��g���_�4<�e�����C�/����N�9'x�XvMgǤkxH����}�秇o/ps</x��}Kb����31�H'R{�\y������Ҹa6�f����;�q/!��ͨ;�8��!�W/d������߻[Z$�js^՝���~��s����şs�����C����^f�__N���aN�^�􃌹G=����^�i=<xj�u+�1�7�$�y(&$�����5O��R�08��R!4�Ie���'�%�mCqN��؇���PU��}'�D\胷	�ؙs�av��n-�|I{=�.s�2ś�d���G����(a�@�vv��['�@~{�7(Ӟ���ovqۅ%��x�F����,��XWt��f�qv`��d�:Vzyo4�J�^]Y�Mi�����r���<1]XR�'�'�f8�&l��|Iy���k���݄��1��a�ݏ���{4f����Q�����\gq�;���7���J����;����v/zɭn�9�]4LHL�}��E�-��+�G/�?9��X�p�݌�߮�9�!�}�ܻ�
�7����Tp)�vU޾�+q9������튙�c��vm��m݋��gl>�O���5����� �������q�܋�=$}nnښ6���4��0�tgy�����c�盍�I�S����)8�׻Q�-�77X���{}�F�{���{z;��Z���p��+��V�%���8�f�Vs�{/�<���sd�|�|n����x�1R�Br��\�K9]^o=�rܺ�㏲B�=�tWrl��q�8��4����K#��㞷׏��#�7O���Pԗ���W��ل���b�۶pen�����x?gk��4(��M ��#�5%B/q�S/��p��`��U�<wW��&e�f�U.y��ۇ;̣ΐ��oӘ}�՝_K���<	�9{FAn��y��#�	A�pd��w��Z�F]mo���e��P�d��d>I�}	�8S߶}�h����1u�-��O��{��@��ƮǷ[�ǀ������r�	!��l�������S����R �K�R|Q����=��0����n��W���;ӯ������7!�;n��F�|6}���@���\�{�/^z*�|��B$�4+4v]�o���/-�8{�s�&��ڛnV<ym�0�x��"�喲�/k">W��M����C=���W,Iǣ� hp�)&��Md��na��.s�|=��{T�v�r��N�<f�lh���nwk�Ͱ�SF��,jTO=U�#���1.��8
��5�L��E�����{���8���c���m[������X�Wi��\���{�Y��y��Q0�/a�g��爄���dB�R�X-U*Ȓ��|W�Y�޹�H�v�@y�sh�:]��rgn�w��9��w7x���Y�{}�c� ew=�R'�W;}��K'vrc'�Gs�|.��C�i8�'������e@��3��\�4�?yn���.�}�"����k���{BYS���Pox�{�x���>�=)X9��ok��Ị[��pV�{�oU��p�g��{�{��|��G�����E�����zx�I��.�w,���z�N�c�".�\�v�k'_Z����^*�}++�xqt^��y�3�s���*t��o��t�j{������w^c�������郶��G��U���0�΄_+h~��?�=a�i�:<�����z�B�ƽ(�t������uL�-엶���j�#!�*򞮇I�<���w�>�rg�@ĵ�&5��3OYt�K�{{�sc�ރ�������D�!jC� ���Um�:�������u#�}Q�/r��t簠Up/��W^͈?U8vӠ��o%�.]v��vཫ�U]�<-�bf�s����xQ;O��`Cs��l��p;��;}��������]��L�����{9i���]��/u��[}Aݚ�7�ŝ*K�y���d~���0��g�K����Mt���^ks���5DK�f
I�^d�w�7�J�FB�����N��/��/��K�Qr�����g�VR���Q�/u��>BQ,�fbżp��z�;"U�K���%<�97�>�l���f{]�U�������/G�	�������B������:�0s>�;c��o���d����/]�7�ǅo�{���;oC�nd �yv�3V�t������h�t�#�S�^{�I=��}�B��)��pUm:�d���08��%h�������|R%wz�kG�+ܮ���3�)����R�]���֙7�ow~�C t$r�������	�V���v�-yV�;��z<��y?o��%�w޷���=�W���^yv�ƥ��>^������Wus=��{�m�=�(���M�>�"��!�v_8��|n�Y@��к�&R�����@�����������45��_y�Os���7Ԁx�;q��k���:[�­�a��N濩��<����@�7s�;x���﴾�Sg��!GbRz���w����T��}� !Og���6��7`�a�zrݼ���}�s��b�+�q5�ka�����}kAn��ܾWݣ�.��bb��mkD:Nt�W�{����G��ݛ�
8��qC��6�7�k
w��fw�5�x�羞 \{��T�zo���U>�|��&͑�'��v}75t��=���(˷/��v�Qv-s��x�a��������q'k�]�{���gj�=��c-���О�m��ڮ��|2z����=��8���퉯Qٻ`�=�|��^�����}��A���;L����ǬxY|l����z1�.0Iԯ>U�лz�e�Zͳn�'Gd�m8���~.��?VDԷ�ͣ�����a��-���o,�iƈ���(���A��8��عH��{pdos�z�/h^=��
وש���j���hɪ{6��ͮ��Y)���Sha�M��ɴ�T�t��6�`�]f.;4:�r{˻wts�8�A���P��d��f�Y�pp����xr��*�j�o��������e�Qђ�7�Hz��beo�k����:'��{|T���rh��ɏL��̨x�m;�=�H$4x��8����?{����-W�y+�9ǜ[�&C����=s�(\}ǧw�V_$x���z�o:����j�Fnm[��J:O{A� ��w�W���{3o�L-�P�J��^=㦍�L�Ѽݶ��u��Pyj*t罞8-^;��v�nᇮ�,�
rr��s��10xX����^�m�E���ʘ���͝�978�S��E�
��u)�`�yӰ�mF�/��E��NyOv��s���{���xHc�{x�<>^�4i�q���Z�&�h[�rV�"��q[�j��]p���������ݏ��{���	�{gdۈo���j��i(,\1O���{��6��-��<�[+�տn�a��k~�&���q��{m�����θ�q�9����x�
+����?��o����@ ����_���^���������������_����G�6�ƛ`�r �Q��ũ4���e-���l<2���Hn'�WS)��R�ShK=u�����n&�e�f3���5[r�]�m�i����ê��h��p�Iо��mv���룲f��f��uxܙ�!,fRV9FhQ�,�6:`�Ĳ�]�-��,*���Xԡ�֏ z�5p�h4eڑ�lv��Ds",Ł��.����p�
�I\�Wu�GIŒ��"�Žoeӈڧ�����^�f��)i��00QZ��M��pG'Ym�A�L�f��a�Z���r��h.#tv��tZ�xr�N1{Y�xl�
k/�6z[V-q�śoSˍ�X&�ݻ.�bI+J�Cu;��s2�14l`F�s�cmj�i\kbJq�Z�i���qp��9���4�)n�u�JeM4�b:���<CY���rY�S�Q9z�틓X�鎅�-�{� ��tX0�aX�Q����RJ���[[�]v6���_)F�tP�4���u���v�]le����IM/7K�q	GS(v̱`���4xT6]vS�m��'$�^nxΓR��.�t3Å�5&ᶽ
��=�:{Sq�o\31�1o@aL�`�/iq��e�KK�d%�\�������D�� uӎ�w���9,e�:�������'����Ň�s�������`�m��7$�:�І���Z���lQ�n�յ��tۭ��R��s鰻��j�n��8��qR�(JKq��Y��ȍ&3��@.٭��vJ�B��p+�H�2�r$�(
hL�w+��
��977��m��5 6�0����.��{��n87F5�d\��+�����d1��tt�:�����{�ӛK�&*�Yp��V޷X-����X�l��n�!mT��� ��6�sN�R�f�+P�q�ݹ��:��ͻH�Sl1at*�+�!�#��]fV��f �4�
N�]�4^ˎ8�Zӧ���h�u���{E�8�]m��q���b�)B͘7rVr^��{�x��nد`��in�d*3B�%�t�--��Ovx1mz���r����C_c[���p=�� �7�q�U�����l�}6�y��Ұ�m<2�`���#�;{17b.���BfV�ZMx�^�����:�2bpy�8�K	�Y8�q�=�u�����hF��M�00���{��ۢn8�zq�[a^#tn�r��+cd���0M��X�pr��!�Ǔ�A�:���+�h���L�kG=��΋����{C��8;F��ap]OWP��eM�G������I6��35h��%"�l1��%��[�#�! cl��nō��YkZ�H��P����ҊM�����^��p�Gdѯ%���nڄ|�n��;y�Ő�ܯk��_kLOf3F.�!�i�]���gh����Мف��x�.9w�ᓍ��{r:��':-����B�҆��sr����[���![����Z搎����S�̤D�#t�m#:�9�&���hw<�8�{:`��#͋��֞�y-Rr�nt�Wv���meCm@5�q,czRw�P����aFЎ�ݲ��]P�T����v[`ȸɰ� �BX���󶨔e���$x�����8���
�\'�W\mr�nMaLBgmX0�õ[n�u����[nj��Z�=='�=
����;=���kv�a��:�nf�y��]��jS,`�"3�PnnI�u�[�Rt�pEs�ɬ`�*�M-u�hZ�!sV��qtj�P�ҙ�Y���\��]��q{i�I��M�X����!�^-��d��ٵu��#Mn�d�8��d�ӈ���ԍل�l�.��:�<����)�g �ea�ڹ����"in�xwT�/�wY�V1��\\;s�38,��PL��Vv�q;1�p�A��*B��%�+�� �jק�D�qq����6U�,F�u�طJ����t��;k&�t�7�8׭Ҵ�s�&x���� �3��δu������$�񣳋�/q��]I\�X:s���vq��ŭ�wr
t<n�b.�c���*��#��ȩ[���{rn$�p�]�Wd��gq�gl��0˺
6�.�tf{6��A3�-�:9�e��N�ڴP�����s�:Z�$�n޻o�osڭId���$m�c6W�ݧvչ�Ûb�W�εˆ��;��ٮS���ϫ��K�0�u;�5��m�)�u̋�L(�E۳�+blFL��7�c�..]}z�:�j�x�ǲV[��*�K'n�; �B��!x��%�zwh��R�&A2�w%Nh�-N����S�Y�)�g�e�:�F1ۭS;�v7c�wS���V-��	��45��%�(ɋ@"�vOv1]��m�6W�ځбփ�oXK�Kt�K[�a����MZ�=�^��N�:���W=;;�Z�t��m�j�.�2���1�C�M1ӃjF�����vu0�[.�f�+'\p51��li�c�@���Gmm�e/Qv��m��kkV�$�U̔�h�P�p�����f7�\#^�SNk<g�G�{<�0L9oes����\ݠ�v�N��z�VM�C�v��L;ca�&���=6�2`�E�(n4�ؚ@e0�n�����ל��r�탷"�X�O�����u��\��0��8�{�0qS�f���M�ۂ�e��Qy���[/%4��a�KMYJ�κ�6�n��j5�9G`Ƕ�y:��\!�͹�ڌd΋����bz>�=���`6�cJ!fʨ�HVc�ӏH���ݻF��ܒֳLc�C��K�M�
�ά���"e�hs��e���a��-e&i`���8�<6��s��A�N��[����n�I{zBC�c�/�<�D����>h�>uϐK�����X��giT�|q-ǬA��l f��ś7 h�,Ҩ�&�v�n�C�M�("`�.��[���l4Eu�t[r.��5�<Bqu�/� 8ʘv�2��T&Ԁ�i�x�9��}����XՒ�E��\]����פ�d}:Sb�ȭ��0Ió�3�nA��s�kl��dS$݃�бe�.'�t�� ״є��56�F�:����2��k�K1ukn��ss��
K�qԋ����ik�Ǎlj��z���&e�k�l#���7�pc�3�n�ܮ���g��[��jZ�l�����`�f-8'uH��-m�v��&h6���Br�wniݸ�Un+��Gb{��p$n2jC�Q.n��>��T5ݝ���&f��`l�<^���L\���9�y�.%�Y�K���mX^����Ǜ���K�h;!D�9� ܳʷo@����]9cf�6��ns�7]���8�a�5��t������R0��9��VZ��L�oH��u�Q���wC����֋�9��V@1�ϣH�t^K�1M������0�6��0�����:=l��z����ܱ�cV��z��F���}c��A�&�1���Z�60��,���M�ի���C�J��ɬs�����g�-nڐ�T�C�д�i�tcbBCm��y�y�7�&C$���̼�ħ�׬ssOI��{\�ص��m�/9����;��������R�q\�:/ �oW��yۡ�*�\�b�@EI����:#h,�i:�	ûV���y�"���Ӡ۴�G�:D���n.��oM!C��-�hn$6���{i�b��jp����1�N�]؄��3f;8Ԫۦ���&H��V��CΫ���u�;��u��8S`�`�=)���y�>Ѩ녹N�)S6R��JKA���O]BW���Ɲ7)�k��F1mnnV�n���Q�a.ơtl#���p⩢\���1��tq�P��Q\+Q+��1,l �RR;i�חA괆�0�b^���<b�x�+�s�o<i���x$���vS6�qp��J�z�b���{Lَx.��T�� <&Iob�XB�B�Gr�L�@��a	��J��(W /�s�
���nƹ:�V`j٦2bSP�,C:����h��t�<��n`ӣ���۶�9�^`�!C&r;MJ�st�,k��ɪ�M��^�֮1Z
,I��d�F��+t� �Ԛ��v�7L*��y*9�*�����E%{�-�6M�m1
Ku�a�FV5s,Lݗl�`!2�3 4aV��t��F4Mn5� G�ݵq�km�s��- b����Zպǁ��Y�:�
���h���WgB3`�Z!@�̖ۗu͚��n�ou����(���1��vy몂��v\��Z[���ej���u![4@�m3�nձ%fѭH:�]�1
Ah�R�4#���������lH�=qi�HݳGd׷L�;g���&1�8���;�G�SE��M
�ۧ������3�R�ni-�G��ݎ���m�ms���w�-�ۊ�l�L��9Crfe6��4�S�ܽ]��g>k�kݴ]�N�n4���G`��G��� �l�T6U-�� �hб�Ƭw��ٓM@��Ib��ڷ�q�k��x��ց9��Rv���;�J�؞y����b�L�ŚZ��]]�ԲmK�-{9��uO��ŴNh���4��鋃lD%l��T�٬�n��ss8�c:��u@� �)���5��)���AE���lG5�^�yړP59���s2X���6��f.u�%7�� �]4wm((ôn�;��ے�[�7�ن�]�s{������A�CWT�\��+���t�-cOW=*%Rt`�9��[7-��AmtZv�J����XgU�͖�z�8%�cz2�D+���5��P��tD�̼��M�R�� K�ml5�{:'wWooU\���䚂Ё&K64���]��[�j�\d:����y7c�v��A��aG�3D�I6ĒEr'ٳ�p�rm���6Ĳ�ɚ�JC������rq��Ӥ"����rt'vYm���9s�$��E"2�BI+m��q�Ib۷8�k����(9�H$�i�mbK���"��h��#��(�D�"�����m�8���C2[V	Ěێ:r��{�I�On�e��I!I��e��������n�&�'e�A8�R ��[j�$䨃��vm�:2�yڄ���)幘�ζ������r@kug�wm����dD]�YZ��t�w������5��,rC��."*N�Kn�pQq�	N�ȤN�2��.η8��';k%�]�tt�j�#2'���k8`�ϲ�����l��m?D`�q]�����5*�Uc�Y	�sLB�X�`�����L��:���Ġ�-�R��a�#��^��t8�n�Ɓ݂}rt���t�FЪ����:�a���v�E����O!�xt"h'krR1C�M�<�l�d���l��ج��L���!��qivڶ:�\v|y�+�u1dՍXwf0B8���s���eM��m�IgNď	�Ѹ�y�j\�RP�p�8�%�im��ܚ�d�!f�p]m�`�	f�.H��V��{�%��{=ك���8Zc�������..��0[��B��V�\���SѸl{�vG�B�b��gh[�`mC��f���3����3��z�˫�'�b��t\E��96hP�=��u�u�]qJ��ke͂6�ŪL��B[5�kq�Ŷ�	�a]GM����&-�D�&���4�0(���@����%æ͌��7����6��2��/��"t�J�MR�j���B�|�vx�����i����Zn�F-�<Z�v&BXگ;rn�8^l�9���@P�zW]n;�ց��2�3�@s�JV�x8���ll��twR�� �����1f֘�
���;�8�0C�����{]�G�=�����e� ���ou��#I�y6���<W�^�\b�E�m����Gg�%�
tb�b�o>�v6я��p:点�kJ�æ��`y���=7g="�C
X�6�Ah;f�� �Y�.�M��M-%).[(�iI�aM�@��)�΍u�Q16��u��ѷ=w!n�sc��pz;�,y<p%r2���|a�Z�<�lŷ�P֓�i��`��\"�-�GBgl�5�wh���fa�"֕�}yӎ.yK�zɫsڄ�d�����t��tpb��&,á)*ь�\[a`�<[s.��$�N}�=�f����6��8��j�T���$��+a9��[e�Ym�1�l-"��-j�ݜ���l�{!Ȧpz�%��V,D--B�����KDj-��u*6�֣`X�HF�Z�r�Qlu ZVKő,e�(�^��gU��[kVՕ�DQ�J�ye@�mi��- h������H[G�eH��Kl� �H,FUp�z��B�
�(���i*��,%Fa�YC7�Î}��$P;8v�Sg�̘�I"g9�6r^�H�Ҝ|0	� ����fIūAp>�[܃���Z ���k8H�.�[��-��$�m���"Ĉk҈gE���,Z|���ͶǗ�t�*���ͳ�$�kv`G����`}~��z���
 �[i��W�7n/I)�O�m�ǉ'v�Ƚ�qTPB�A��{hf�N]�ˢ]���'�嶚��)#2����gfA ��O�@$ֻP�/���"c<����0-�1��b�+�=*�m����g���8�q�#�ӄǙ;x~+$����F��[M��H�Wj��guO�~+7"<�m>'�^̂��'D;8vp#���P�I�@ԡ֖��)F��
j��D����p�S�i�3x�lV]�Y��;E�W��٘����Wh��i��F��	�:a��2#^��Џ�/�	�y,�{PH4)����Gv���'n�t��.�Ln4G� ��v�I���9���S�dn���n�Z�Nd��$1t�_,~}A[�}���D����^��v�O�\mUe*ˆ�eX��[e��7�r]:�`�:�mg� �&�c��-3��@$�fD�N�]�9�W'{i����t~��un��ߑ;�D�hˆy�#
;�`7���3��u�:՜w������+��tK���� �kY�O� �Ƽ���z��=��޽��"2(�gd�	fgL�d��KFDel�ng�f{^"���N\k��M�6�dFV6��{23N�;8v|ml6I �FDA[5nF��x���Ӗ�D���l�#hnӵ6Bs�^^�� ;�,�n�OIf\�.�ާW��ӈx��� �==���s�+Fmf=� �r�b'2�:v΋�8���=��f�߸���  ��!���m>"]9ܪ��x1�']�]7��K�E��w-�Oy��nx�_��"����7� ���x7=�~�����>w�e��8�n��1���j�9���p�c(��oY:��V�s�����m!"��2t��󾼘�d�ge�}1��an6>�^����9M�YӸ%�p��@70�`���ý`�8sj� O�>ʛ��$�v_L�����+j�/�|�J&t� ��꘹��cw��!�:.��k(�$���	�?k�G鄜$"+O����/��[_��\z ���P�3q����;���	n�_�s�3D��B-���	�y8���-���z�������*�Xu
�]`J�99N�ou�2�y׌N�����h!bR��׃;�5��8��yȑ2H/b+�!�Ӫ	�#w�֙ګ4]��X3��]2�2<r�s�g�J0���ۀ�rr�L���l������77r|�Co��� ���bO��5����T&g���f?�V��#�̉wfb��(H$���5�w/��v6 �MқPH'w�xǐM/@���N��x��+�-
3��� �VIh*	�h��k"<Cj�p��)�mK�$��TF�=� �F�J,���ӧ�.u*��C!*�$�1�Fݽ��q���=4fIw�v�P<O�����
ԂI������?<nK�G#���}PH��{1�Hˍp%h��*A�b7s���F$��"�ӆ�"Z�Զ�i��=?.�����T��Py�]�y�h��zU~��.a����z��}?(��|'��-��Ν��P%1thPx:ݟ"{sN^�|��Q��,9y���FS�G���wb�뱇�EӞ�w5O�ܢTa�k��J��� y�e[�yڳ;������Z�%����F&�[3y�.m�,��@�7n;'nRq���HO�����vu��'r!�v�G]A���8�z��&l�=^�Jk�(��t�������Ps��CC�N86{V̗q�sg�M
���n`�ck�,ˠ��Gq�5�OcA��w�����F�,��þq��ف!�� ����Aˍx>���n�k\���PI#3S�EΌ�$0.���r<v*\nѧ���S3�lY�A ^6Z�|	9q� ͪ�֋��
�ŻJ÷�,�E����k&�D�����H0�0�����ʬ�@�~GZ�A>$���hNu���t�a ��X���
�v��H;q�'uT[ ��nq�C�=� �����Yٙ�b]·0?Nl��l�N�d���g� s�9�7s� �Tӫ�#^�ŴN��� ~Y�]XMT����Д�iE��a
=`8f��+�u�9�������r�jh�����i�Ǐz��ƭQ~[�o+br`ŪO�`�??͌�=;t�w�,JO�Ր�R��Pue�hoD3�NAr�-{ڱM�����d��oz+�T��Zj�d�`efS��l�^:/`�ۛs����s��=�c�{g]�Yំ^|��u/�m��� �����	�Hl���C���ퟙ1��I��UR�Q�I3[0 ��F�N��Y�t���b��'�K��߬7�f 5���PO�ݷ������A�ce�H9�L]�3��t����Q�Q�@3��`�8�79~�C�dA'mM����oF�h��Ȅ5ч�u9:�1@d,��MQ����D]*V�
��;:�M�<Sp�ih;:jq��[f�,�̟�Ļ��3j ��7`|Jݸ� �u'h�E��"DH�i����J�H�[��þ4��#j+v�	 Ɯ4|_6��)�9��ߙ��0�~�QGsQV�����w-��$�@h�ۖ���:��!Ӄ{��F��B�2�����}�`�D��G72�)��8��8�}ݰj��g����C�wk)f�\����t:}��� �4�H$�{0M���`]����4�r���SGė��Kyg-��$��F�ڭT�����״"�ϯt�:I����s5�� $�d��$J����$^��O�e��� ���5:��>�h�F3�,���Q\��q�+I;7n®��U�K���E��n��;Y�D�N`H��wvw�p�]��Qj	w�'�q�*fޛ�Q��̟V>�׳ �ȩE��3�Rt��A���&�52�����^b��q�\l@%�,wS5O�ج��d˖A&p�����x[� @;q��#m�p3���R\��ē��	#.5���I���S:.�&5dc��t>��Ppb�G��H�{�� �Ɲ@V��uY�*$�A�뽑w-G��0ٜ�{���qlV��&�Jso��K��~Zom��'s�!�g��S�����3jo�}��|AvrE�k91� �ڝ���w1�RM��(���H$��G�bB��m��_<#��S(�4�@b(��eه�5$m��j�2��nXي���ԧ�ٖ�S�EÆ,���I3q���:Ӫ<v�=^Υ��ݨ[;قA>7���ӳ����]�F�bs,&�ehf4Mn4�H�e�L�ESN�$��3qԻ���Qp�y٧Q�X�wV�Ra��^��d��Ě��L��Dȷ+�
֭BQ�$�;�d��^6lRy��[q�^1#<�E@�O��i� �Ƴsa�N6�:�܈^Q5:��;�HҴ%`~�7�G�����$w3��ŵ�	٩�'�δڂ7q�� (��Z����ģvf��U2�א���ͻͱ��m�3HKz]"��w\��%Ԍ?��2j���E�xg����?,|��o鱢fad���f̲�Ik�1�c�<�R�c��n�M]0B2�6n�9ؽ�̡�ზ"��θ�q��)���ŝ��n�����`�8Ԟ�"Bj-�:�,�n�Y��n�Z�.�X5��B4����X��@a�tqh:g]fl�!*;q���Qk�1W�]����-]�/nZ����:�]�M�s�b��F�k�;�\pMi�6��xD��p��\z�@;��̓���Ĵu�#�'�����������6��\�I�S��_�7"�N������M�V��ؿO��V(�ѲóPZ, �'�L9���>���u�#=�Q�I�$'q��&�=mk�DT�����n����32t�+�m��"w�>.���������{"	�n=��;��Iӧ��{��U���h��A��cA��5��cē�"<���i�om~`я�	<ń�N�8tY$��/� ����J���,������̍2	 ��{0H�r��@�P�d4�Ǉ���i=��;%����k�*���Q��{�S۔�&�Һ��Գ���Ce��Ȼ昫h����`	/e��#n�R�<A��&�@pėw������ !��b�Y%�mX�i�ދ��p��N]�VWxE�֟�|��_]~���K�{�����Ȯ��Y`��(&}��^���Q�ƣ����dG���q��mj4���h�Q�O���kˢ��2u3��	'�of@.�2�&�f�a�A�����v�b���ə�)�3'B��ݣ�K�5�U,�ᡮ�W��v� 	�f�D�I"�^�b���n˖������,Y�N$�:y�c'"yy^�\,[�D<��m�e@>���@$�9/�e�d	x9k��_.;}[�Ms]`x��ݕ�O�pnl:��u��p/m3qm�&,����߿� �i��ϑ���PH'�.2@'}[P�ŔmH��C׭8�A�q�>�NͶ�wf)�&tY�V4@D��zXT�ˍ������	o]�x$��}1�������ִ�DV����.�	!9N�TA��-��%X����ӡ��|v��۷oo����<�=�{����N�5��1����;,���^���|���L�7BWf{iǾr�	�;��e�5�VӀpF��w}����/gz��!h>^f;�olJD"�/T=t�u�z>g5���x}t�[�,�E�J+�l�^O{ݵ�b��	Kh�٭�$Ҫl^_���g5/D��3��Q�ON��ȓ��鳦�|r��Dg�vi!e��ΙfUϭ��4���d��-m*�NL/f,�w���X��'=᠅�q۳���m_ \���܍g6T���ld=߻�ؠ�Ox�����e��~�=F��KR���R�LU�$�����@�./MpU���/�E��	���E�cS��25��v`}읾�/���\$*��	v��i;�`j��r�3��=�шV��B�<**\��N�WK~~��}�l��O��`�Ǟ�*��VƯHwAoP:7.����ۅc��S����wӴL�me����-q7�y�wi��C�w������D폱/^���j�/8��{�}� $�UE��}�=b��}��4��:E�M���s�ɖ��	ℳyu�閟�mW�$�xSh�z���Fl�~��P�^��U�T��^�=}������w����ȏU��xz��J���d���OH�ǋF���J^�.qp/`Ŧ
�q��w�K�<}7�o)U�Ž�t#�Z�ɻ�����vg��^��.���0�v���f�ל�9������?[��v�����қ;���0�;_����^���!H�f�|�ˮ��5��p�=�Pu99�I��A'�\l0[U�Y$��ht���Y�qĜ�$����v�T%���f� �*);kSk9*2ͭ���e�A�mG9��%$E'S�G��taQ�'m�����&�Z�qQ�nĝ�v���kY�۬��� Y6�cC���tqvef������㎾<���������I.	m����>Z�N䜳���>1>|פ���JFռ���N$�Jv����('9}O�k�Ƞ�m=�д�K[t� RZ۲m�[o�Ļ�v���/;&�k�DB@;������s�ޱ���i��	��0[ͅ����x�I�um��	Y�,�bmd���){X���ݵ�y�՚�#��w�d����Hm����ei��{[;4�6��y�}q�gJP�,��þ�q�+!�uG@�"O�D.Ѳr�p̝H�<�#=.G�i��FdXz֮�x�(��>0��	rLa�;t<C�2�%�}������:��7�x�:�%)���Y��tF�3g��éUǫgO]K����'7�z��-�m{g�x"�2�.�O�c�Ȱ|�u�=�:�29��w�=����rR���{�4Ðk��s��y�/|�}�1,t�:�!5�MYQ����Q��έ��1l ��T��VZ�>_��۱.���8�u���Ϟ`jMK�.d�{�~t<Hj2C#!0߼��q	�$x�o�T)��>�`��Qk�H��J#�潁�"O�D �Ep)��;?::����Z�'A�����f�߼��q�}��/1�Y��亃!2LHrL}�=���I���Ͼ����H�$"��=���Dr~^��$��]�ݙ�`ɝx�<(��<�1�%ϼb�'��ϝe�L���JN�����r3]�2W��( �� #�װ<�K�d�>��^u�h� :���p����s�G����׽��y���c�w�ԾA��I��>yө�C���������)Bj�L�;�=�� {��Ϗ:Պ8q���iڍ�K���I�1�D��R����l�x���Ռ/@�[�2R���7�����w��Y_���0�FM<t����x|��	�s�~y�����;7�����98�9�	��z랧����J<�i"O�4�C�>�{bی7w��td9N�f|�=�P10|�|u/L��E�%<�B/����M�
��2������ �n�c;0�봮�@�VJYh�5�]�|��e�qL�Q,3�'Ā	�h�c��a�'���z��0�!��~�Τ5��u�w�[�����>��� ���|�MC�kz���1rs����q���G�=��&���������8�;���箇��c!0��֡5d&���w�u˩mb���D��Ne��,�ٝ0<�����T�Κ;o:MgO������d��(2\��޹t��e�1� :�y������m�v<C�2�%��}�Υ�Jd���Q�L��z٘���g�#¼Q�m� nμtw�z:�>�{��y��	�0�!������ԥ)N����އ�}�]��Y��9�h9r��|�:���^�{�����#m0�#�u�)��${ď@G�1������C��*�3E!�d&sߛ�P��%30߾k�4��+ ��=���)D�n�W{盅�強:� O��S}3��n(���u'������5�}'��\���.t��Ѵ��8s��G|GQ�"����O�CH���ȋ�H?�<;�Ў��,Y�7��3]�̠�m�V�ì��FS�r��θl��Ԙ�{77]��\���ok�4� ��<�����םO]��4��������lv�b/>N'X!�����knN�2��ݩf[g�!��x�b���r�b�ю<��:�ە�
Pm��a��lnփ453	�"A�rY���dhk\�`D���lKb�k�io��W5����*�鹇ͺ7�z���L���ueg.���B���.�	��G��9�Z�T�'�	2(����.��rR�>{�~�x��ᓓ��{����i侄�׽�],��B#;ZO�$IR�RgH�b��d��%���	.}���<ѵk.ǇMDE)[����=�Hud2R�V��1O����G��%�O,�16<j� �y7;L��.���4�T?	27��;��D.A�y��ӯ9��>�'�ݑ
v�1̳�ڇ=�3ĄՐ�Y)�a���b5�R��|׾��"A��x��E;�.����G�F�A#��O�`>�@��r;���K�0�$�rL|�=���CRd�.�{�]P����|�F_=:�ÀI h>G�"�x#�ڕ�t��e]y�Ξ�zy���Ξ�׺��:� �x"�iʙ:�&��<(��F�����DN��{�C�� �\�!߽���4Ð�׾�������� ~d�銬nS:#(p�J:�a�GG
=[v��'h=q�U�??�����+X���y��L�����MK�d�A�o�;��D�!��	���T&�	� k�s��gX��$$��x	����d��~t<JQ��:8�y9˓8�s�5	ǽu�T��� �����yl�-\�ח�4��ld^��3�7A��p,P�v!ܶ��w"4b�o��9�e���yr�ƅ��׏���=�����>�������]A�.I�9&{�=�C�-�L����κ��@G��;m;�.�Z��Yn���$x!�jV�����g2H�Q��i�I��L�S�=���h��!20��8�^��g��p����Jq���z Թ�&��κ��9&{��vv�.
vt�=Dz��Da����g]w�s�o��{�ܾ���@o��N��R��07���R��%03�zX7fs��	d�H>{�� �P >?�=IzB�|��	Jm��޺F�@s��t@d�x��r;���	ޓ�sn����v�z���|K����L�$��������t0d�",�K{��$�4�i��3h�>O��M���6��0GQ����e���/�)��u*�؞K?>���Z������m�N��=t<Jzf)�`��:�Bd�)Fw��\!����<��|����g��׀w;�|����z��`�	#��!իd0`]Ӣ:�C�:d���]�$ԹB{��u�0>����i�B#�^��j��ud�����k�������ţJ��=90<�g��D^��7'<\��<gBj>ֵ��Ju�c.G�~�R�%�JI�9����ܧ�ܜq�Q�+��S�"��mݐY�6&�B�9�>�,�f��;	��3���<�x�åH6~��~�_c1o��Q�*Ц"~z]��y��	�W'�����t��9!�dw}}k�:#�g)#�wDb���(�	�G�%��L1�p�!�h��B^�^Hx=l� ��BddFy���ԥ:��Ȯ{�c�5T���vG@�;��"<2:b	��|�'i���Ĺ)Ӧ��>�F�o��&��2\�$��;�D����4�uε�>|B#¢z ��%��d�9��}���)Y	�5�y����������.��]�	7�.�sFU�mͤ3m�ڔ�G6g��Bd��it��r�3��-"�4&E���;�� �p u��]S��<O�`K����p�R��� 0>o�����2C[k^�����=��G͛����>G�"o)���@
�56N�Y�fp��*�O-�c) a��yƄ�k����JA"P�ަ�$��k�iI$}��c���Sl��.Q�7�`]ӦH�a/!']9d$��b��tJ	�:���T;��	/$��m4 $�Z�X����.���ƅR鉑�뭣���(�y^�D�^f��6ZBI$ٓ��͎�Т6�Hv��B�[J�ݡ�C��Cpa���A9�mw/	��l��g����+Xy��^9�Qob�&�+�Fsђ��"%,d��#���� ����v��o3kԶ�S��L3�3����e�I �}�en_�ϲ I��$��qm2�%�ײ�I ��$L���C��c{I�O��ݹ���xL���71����ޫ�1���r4��5|ﯽ����N���Z����g�f�ȟI"o�۲&�@e�2�F8�����q�Q%
ƾ���.n�'D$�Γ;KJ~ݑ J%/;A6+�54U��wU�4�� ���O�@z�f�/��؇�lN��f��3�P
5l̇H$��́ JAg��d}1j��H)���xg�j��K����RK{#�U�u�����LPt���ukz�&���vV{S��MJ2%�̈���&�u0�"˪=%�ل��n�iIV�����wc]�g�N	H$N�ʐ�|v�|e�F:24$�[oKJK� �60̢�F�u4�1���&҅d1�ט�.�7e�dʭ�a�>
����I����{�'k���?n�� �~��iɻ�4�cA�4��\dK�"�gURd#v��x�{�N��@�$2vEd�������δc���O[Wetb�[�F3i��l��"��.��b�i���i���F�5�x�[���X���e�Ќq��iM�b7F`X�nhK4�U�2��ݛ���+	t�b��EP��Hzw��u�-���r
��Y�] ^�{l�zk�N;�u��\��GO	Ԑo#�zz3��nfϭ�^�Q��������u�t��nn��S6�*��l� �X%��m"Fj��-�t���~����$�&r8�l4\1�H��|3(�U�u4�G�9��Rf@�j�be$n���9��1Ĺ)Ӧ���W\���G�Z���$�b�cγ2K���D��G�r�Ns<�ZH�.�Έ)�9fu-)�cLHl�=,$��!1|���K˻c�($��)\ƶ$HGI�R��������3?*�U��O�I%���L��HcwSI$���c�s#&�^bIwdY�%/u~(0.�ɋ9L%�$�'�$�x��C�z��k�EZH�3)/$�����E$�����/z��_>oy��7��[6���b� ��\��;�M��oR�ũfV�@7��G�?gϵ�+��ó��|��$��I%���� =j�R>]ݳLSb�H+��2%��Y�ԤJM���Y'g	'	3��N*�������r�2���t��s���a:�x��s��q����zd
ܓ���źl�@����^�O�-ԞY�)�"�����>�}}?	I%�^�}�2Q�f�k�ZR$��T�M�tpJV6+-�t�)�v�.�%��j%$U��%�	 ��2K1:�sv}�6% �_)H�	u��j�U�nWa�3;�	���}1���vU�F���Ki�e�$����e��J��ȳ�>ه2Ϊ��\��0H.��R% �{�鋲LY;��UKel̺^Iy.�{0O���vf�]�&�=��n�L��2�[�f@G�=�QhQa���.��[˶;9.nb��:���Q�q�2�%��!$TE�Ŝ�9a�{0����&.�0�k�Q�R�R'q_D�^H��|1){��8���ڦ�h��7�ֺQ^IVג��q�-��p�\;;K�"L�@$|���Z;�y寸�A%|ْҒH��3�E$3�7`7���	�3bJU�lƁvp�p�9>[+�gΐIy*�|2%$� �g���������g�=\�K7�<�.k����=�v&�PX��6���Z��xТ�q���~ӧ6 >���$�o�]��k^W<�q����@����jߒA%�ݒHI$�}��4d��Μ3����ͥ��K�{B�R\�%��U1!�I%^ӏ�%$�U�Խ��ÊwSxI�S�d�2�WD3����s/!>li�>I%��R��ڎ�z��lA�i+L7�H-܌3 "�J����(`���suۙ��i.��郢�Ӑ��z@k�W umc���fi�������������ɬ#'r��E�ɐ��K�s O��I
ފ2I�]�"7��e薎���W�"���N�1w� I�_JG�BBCK�v�lK�%��!%����>�IP�������[b+�8[r�ظvv4*�ډ�>��'/��H$�>�ӔZ�
/-ۍA"W�vd��PIx*�3�)g=��Jw%:)3�3佒�P5�Q
!�- �J�6�R$U�f@I$���X���Zmz�гN$�<L9��p�����>��S����2���o�L�I���#-��$�D�e'���S��|����G�xx{�7�$sj�L�9��gN\��):.�T���P�'>Y�!���G=tK�S� ��&|����\�fQA%��얔���U3�-a��7 �d�(�tY�����k�֊�u�n#� >��t� F�s_;��˴�r�;�E���~Α>���,�z>�^H�+[�ZBG٭�>Ѯnau�Ȃd$��v(ϥ �׎�:,Y;��T_��1$r�so�	��f�R	$�۩D��!\ݒ��>��b�tݪ��'����mG:%����_^�'zg! �dK�y�@��LE�s�H�'F��(%\�!�%�g
�\�v.�z^ G��,k)��[m�!�y%��m�iI$��d��vؼ�ѺL�|~�2��{f�Jw%:)3�2�WTˤ�5ې&WT��nc�0@,�Q>I$��l�i	{� H��O����{�c���{=��g�������-��fu�t�D�4U��<p�q��<���:#W8'x�>��C�K�gzcd`�����o!V=�*޹o5��	�@z����V���{Y3���<9� ��N����������M�9���~~��{\\ja�|>~�hf�>�Y�{�=g�&Ul/��_�|Qo��,�Sܗ1�a�b���"d)ؘ����c��x��;���+�������Zu �d�k�w[Bk/�|�����//N�X��&y.�F��z^����=;z�?9o�=����G���{y�Ю��v�ٛ�:פ��3k�|�^�;*����1���X��G�e���{�v����[\�e��s�:ހ�V�q�Z��,�����N���B��c�O�(�◳��3۬wޞb�i�?y��d�u/:�l�u�E���_��?�kZ�b}��S��#�<_z\�����7swտ,���_\{4�zn�L�A1��p{։�6\����3g���w4�^��{����XW����n,��$哷_��߇��g+��|�Ê�v�>^����u?3P�pzx�l~E\
�5>�_��j��n���X���;B���f�/���۝���Ð�Z�Q2�s�G�zln͞\G{�>N՞wJ��.��:�M���u-B�b]U'w['�߭�>��^��û1�J��r4��V.�]צQ�Z��wy��@��6��]�C�<�Ż��\�L��{{�ϭ�3W7y��\zP�A��9S=�{@����� Ȑ� �e��S{u�L�؋vm%4q�n̦�R%��l[�d�m�LQ�l�n�թ��$N���xYȄGY�q�ym�^v���{aZ^Vrq�QCk=�8D����lC�����g%�V�݇�ya�i#�p�rw9�ݽ��܎m��#.�9"H�N�k�<+8�8��p�,��ݗv�I���y|dGg�ޑ|�:"|c��:*����BtVv�e|u�v��S[�;�o�����8�;��⣮{wY'Y�ptP�C��_=���K4�z�v�ʴ;��N��uV��o��{g^��ː���U������*&��)����^^uq���)a,��� uf���D\�usT��nݕy���[�aM@�j��)L�]�h��l!Es��D�z�R�^�	��5m�b;`��\�y[���حm�����:q���j�ݮ��k/A�� ���!�i�p`���W*V�\��n�LěF�g��
��ơY�m6b�n��1���ێ:ڝ"p�{]������a�.�.��P�Wf�a�\�ck7���#u�ۄB��gm���$#��p��Ҥq����pD@���+�)E�O3���7m�ѳ�6��a�!�6�bn�cV�,.�"�˻�x�=�f]qiX-�"B��8,���0�'W[��o��<[�����1��y
�>���H�Aem]��x.g%]�ó���[���@��p-��7%������ے\]�xB��u�Ԓl��F�q=���r���-�#44Zb,���NN�&d���JZ�&���f]�h�fi����h�3�1AHĔ\���;��r,w��kgU�������nl����6ի��σ-��{tu�mŶ�^��M��z�5�xwA��ɦ\��S�`W1a痰h0r�7��t�aJ��k�	U���hZZ��O!=��x_�]5/Lk���;�Y3@a{�ə�e-��.f��"v�Pb1��;�V���{�V��q�̴2��2���c�l&ь�j<��u���G\vn�SLKj��zTڝeMnɕ�^���^�5���=[G1�9Z��E'�}��c]h�FR��K)��n�g[�o1Ծ^��1rݙ�q5�q��=,rt���+��ϸg��
2i죂+p�60²��Mn7V$078��kx�g� v�pʝ����F�Ů۶���c� jp]y��,k���,����k�n�ۺ��u�<v��\Lm
	ɮ�l�����l�n0���3\�',�Q��V�B��g8��<��:X�bݍb�`.[��n0á��#����U�[),Zҁ��6_�N�W�#@����Д %�wC^���z��X��٫fuuq�A��lba:� W5rpD�[��.).��f!�T�Ƽ5�˥�P�[ѧW;+�:�݌�ݵ`M��F �P�����ΛY�T���xGv4�g\�rvأR>����F�x�����tI��ʃeն�0(1��X���9�WI��N�$��^Ԧ\��拧.����0��nX.q���-,��O[�=6s��BZL��.����`x���+�z�)�-Ic3a�#-	���;��.�w.�p��Q/���I'9e��o2-�H#��L�'P�MA��X�1A3��u�Ly����!���.�X�n��J^I�`��+�յ�4��^�n�iIy$��$L�����4��%�ej���s]�p�2w)���'�� �	v�@�%K�g`����խ3��;���%��2�
(���d���Z�S��ܦvp��;Fjֆ�`���PJ�tĺ^H����!$Au�R��
�4`$��OKH	*:V��p�YѡT��dO�/$Mcu #(�v�g��t��ͳ- $�5��'Ҋ�G����9���Z[���C+6�k���t�4ij��b�k5�[r��H*v�e���e%���g�ݷlS@����?},��I"k��A���u�J�I��9G���v�54䴤�|����|6r��b�Kt"
6����f�������Y�\�;0h�F�\��X
e%�%C�,��A����u�<�"9�?nWK��ŰܣP��݊��{�|G�J�* "��=�=�s33��"g� 	K��� J)%�Ĥi�vꉚ�ė�rWE��!ܸ%ظ�/�� �Iu�ʉ"e�1P}ݬ��Cʞ���H�^@�DH.��Pe�����'r�Ȫ��g��l�����$���	��%
��S $�W.�gg��y�	�N�$�簒Y2$JC,vF�r]8t��Y��CNϚIA,���n�~+����n��$�H*��R�Mj놐���Ŏv6��D�s����y�X�Dqs�U�i���PѬ��=�`�j�j]�3;�@p��dS�rΎ���dA��5�֢@H���!'��/O�HhsIڙ�R�$��~�2��u4�wE8L�ڼj���\˥乶
�6��76JA%��}�$ϒT��^RA&ޫ�� �eS#<%V̊wA�;�.ŝ�h%�R҂GȬ=�d$�J���F�>�q�S�Z�R��S��#�a�`bP0u �7~B�~�1ȷ��P��G�|��]�h��\������PV�V% ((iD8מzk���2���5�E%G��yIxۮ��ټ�\�e���C39@�3�U�$�K:��i@$�Z��^BD��;$7�3|E�p���q�)z.�1f��SL�<��{-�	
��1�]��V�$�s֩$��n^|�I-��(��g_�z���ێEˆE�:s�:�vx� ����g�/5��>�<�`x�������R�p靜�<ܕCNHiA$��뉄�^Im�H��6\gW0�1�yE�X
u�!$-vܼ���t�X�)û'&�P\�2 �Ob�#Y/��2e��o�y�2>Vݓ/!%���"QI[�/�z쟭k�emr�M��Y嚋wI8,��L����] �J���I$���E�훭�W����Z|��G���H�K�"��wgN3:��%:��j��Y�#���t�Wj:%��I��fnЪ	i_[G���Z==�)P���.����l=7b8�	x��+ջ��K��_�gՁwc�?xK7{Ð�<��q+�\>���vH��y1�8�|<댾�}��V�Z�I�<6l���?�H;7�˂]�������)�1?-�h۲14�r��%j��&B�ܑ>�I^Z���W64PŹ/�����=�t��k���R��������Mv�@=�y����M}~>�qm]�������(92!�[��$JA ��^�~�2�AUə��s+��)nd���J�rDԫ��.wd�6�uD�Q\�y������BA$�;r\&BHf`�߱L�ME󦥮CJ|�<�|��p�:�dS�vNM
���dH��IV7\����K^�1��~��ԗ�^]{�$J)$[���e٨�wt��̝�J�=R����L-6�J�.�H$����k���A+=���e��ހ���D��vE'A�س�	�UPJ1�������q>����8=U��~��2I��S(�$�w\������ΐ�ԃ�:�	R�&�����{7���&P�M�w��Ǝ����[��X񃂴�V�k�f�]�����{z[��8���n�/]pk�g����Ƹ�����"@R Д*�'_��0��9��.;F���Z��c=�]%��䛜�K$n�ݠ;z݄�m�U8�7M��O9Ů���WZ}�/f��kW�{\R�t�D�
��t�`��.w
���l�ǬՓ��8۲VۡK\#�X�����Yt@3xtΜn݀{mn+:^3�gJ�
 lSQDf��Uۂܜ��C�prH�i�u��=b��%�l��ڸ�qW]��@��@lk�L �rY�3獯�+�2b�oC�4!3��`0�n�c�i�>�7�f�rC��P_7 }(��suO�RI%K��Ϥ0f�3�9����A$���Y�M5��wS�vfy�Pz6f	rn�Քc���/������J	!V�Jd$�Az����"F9ך�S�r��׼xm��vr������2җCNO�IIaθs) ��\U�c���'BGu���)#�]�!$0F�X�Iû�&�����ê�u��$��_(��	*[�/!"R�̐�;�X����sE��<�j�He�3Qr��N2v!/r���	����"T��~
�DC81Qi)ǋS!"l�\<�J[}� ��ʨؖ�%�s���]���Dzb[�=:��4�V`��<�y!����.˶�?}����f��������JH�p�\9��	 :�$L��bg�*����5m��7����-W�/>�307��vo;��yO]�&R	 }w�[���s���0K�w'p���C��<e�KT<cKЃ顀�d��]��m�/�@g�C/�k�uf�H\����" �76̒�fٔY�%��zm��]'����� �ii�B��${��ڵA8��e������I ���D�(��L�$\�\N�Z�K�9��wS�vfz�
F́�K�r�R�I+�܋uΤ<�F�MެВ�HR�y	$��d	����7��',�N�i�t4��ϻ�k��8cW� B%�{ D�%�f`cŮ�����cG�Jb���������q̝���&�W��L���IV7Z����V˷��wIR_�RI �w$H�RH-��R%;н�x��ۛ��(�h·Bե`�W-�p�q�*X� ����<Z��;]���������Y�����L�	y"r� H>���Iu�b�	d�lu�=t�Ywj#%�$AffH�"�Rtܳg	�D�7J�	?��cr�7tgn$K� �ے&RI �߭A2���;c{-���� p�RAك�N	v2����"�%�[nCJ�K��G�T�B ۳S}e:Q*j�KɁ�u�^��s�j���>��`r�z�$G���ln�3�d���V3q���	����^Ό�sq�Z��U�=�>$�(�� �J�R���K��I,��%䗗[�j���]�9N]ٙ�(=8�+[�Y}�US>�q�I��e%��jI��뇭��+�)guw�R
��D�V�7��'d�'r�6z����2�J�D���[x#m�(s����2zDϒK<�km��Sy���C�L�t��q9!�?����&�����n�׋Z�G���l�C��Yi+:���~��>̲N����D�H$Mku�I($�ut���1���7w[52&Q@$��kW)l��&p]�fN�$,3=3	%2�ae4�����O� �Iv>Z�I$�[u���$���v�"c��l�y��N����3��U%8�rP	 �ձ>���;1���®�k��I%��jD��B��K�I1ԐN�˳]�����!��M���Z%����)$�0�n�rd$�_d�G�?i(����?�5ޤ�uQ{��]��Olri{Ή ��A뵝���b�N���{������p�罾��χU"Q<@� ?R�R��
* �(R�\_Ff�\��Ѭ��^oo'<�9A��3�9�FxBI �f�	��Ynpm9g��%���[�/T�	&U�/)%~f�n~�C�Èc`��S��.�Lzr�U�\3s��;�팒�r��;U��B��������tY�Gj�>�C�?��s��a�ؑ	$����d���d�*n�I��̴��J	���헐��ӈ`tȸww`hQ昁bR��y�c�gCi�Y�h��J$B��\��D���"e���nl99<����#na0�I�ŋ��ZcjdB1�̫; O�/y �Jzꭟ�i&��;䗒^��^BI$��$L�qM9gN��g�U�[�z�v����\k*$BA$J�rg�ϒ^H�7Z��m��j�<TbrFy��c����1%�˖��%$�]��->�ط����l}�IZ��yI��rD>I��je^_E�����3�A�g��FjK}�y�]q-���l�x8&((�T�"�fBa"C�2�M)^TD�{a��Q9TX��#�=�>����$M*"�R#H�(L"R�)J	B��y��:�ػ/##d諜)��X�9z���ni�=g5���l�g/[�85��K��dL�F,s���!E�L���RlD-5���Q,bݰ�.(]R(X��c�;h@�Q�vJ����m[�z��[�;-e�k���v�s��Yv��3;&�r&^�:�ܦ6���r.�q��e^'�Lg�xўn��m�q�0�9�������nB�6��:��kL),p@�&�H�]ղ�fn��	������m������o&gЉA.��(�������nY�>�,q��K���$@(,���K٬w�,�ػ'r���%�ճ�Tl�`G�����	�B�2D�I��~�5�b�绦=io/�I!a���;gv�*�=L�$ϒ�n�iI �R�S�����	%��"	&W[��VG'*��rX2!��HXc�f�dwiN��c ��K"�Iy��Տ֥y)	!K���eW\]cU�__���DdӺr����UD�7N��K9eĀ�	������1]�!Y]"g˼Ȁ�&��S(��Z�r�Ր�%�3��%�`ᙝy�p��7E=aK��W�u�n��T˱,����%�/翥	�9v2����"��Y���rI^IV�܀�,�6�y9k���DQI��S�Kɧ�<��Ô�3<z�GCl�)-x��9�,ݳV���;�UA�S���vz�fp앰�g�F�c�[�8o���W�-e3[�L��<�L�)ݰ+��U�҇����]I�����e�R	J(ZP(()��F�&(P�
��
A��)�J���������j�}���!�>��}%$�V�"�Z�c��Jn��tɃ�윗>�/�mf��4����x&|��Y27�˗���ř��#`�I$��|�ϻ�7���L�%�4��'����3�Ȯ!qS������	l4T����Y�q&RI%��!�3��{�,�C�cM�	��S(*9AT���`Ȇvq�^,$J	Vv@�S�t���k���I��e$�[}� ��wj<�ѱW�|���#�E[(Sj㫆48R6���v[�Ǎ��$�����O'��~����}��y(�ʐҒ ���I$J��2�17�ʪUn�[/���du�Ēd�x�Bv��N����D�D�����(����5#�R�q&@Iy$��$H�PH�[7.~�Ɇ��BR�������C�ϗy�̔�>n@�JA"o½��_����_����{=��o���x���.�fmcO���8��i�=]��Z˨�9|[�yPm����H9��x�%b�I�1b�YWW#31
��.����mP�<�G�'U�v�;|ǱH�����:�]���7}j7<��<tg�A�WRc�`��������o�QܙY���}���Vi�X^�t=��.�>���i|�ɾ��9m����Rv�w<t��% "4q�z1�/���`ָ�{��.Ӄ&òw=�(��t%�r�Ҥ�˹�u�7˧y��v�r@��
��sfU�����w��yf�{��p=�T����:��B]x�n��_�'���n ��'9y�Atah�!�Q:zOz���Oyh�Y	�����v�~���&w�g�w,��q�7^)sCC�W�9k��ڽ���8i^}�R��}�z�>3�,|�+�s^��=�jWO��%�o�����r�%��x�Q�e�#zq�Ӟ����DzL�=�A{#�#l�QӲ�]��i������|!n�	�����<Y����s��j�}�efx榝s�-ٿ(_jP��m�&>'6trm<��=���������*�`�(|	�g���)�U{�J�~�Q\E�E�U�;�磇\�w+d�&_<�R�]�6uq�=\��P�<���|�� ������k`S&�c����ܬt���K��Q���_h��;Ǜ]��A�݆,���<��
����C�z\Y�{uz	t��D���?_�";=HΩ����[sv���(2%���s�7���'Z
ljX�����'%������$�.:	�Ί:����Ґ��/+:��q��'DErtp�ӾmwE����=�u��Љ�q�r@68#��M�ӣ���ga:��;5 �8��"�ऎJ��$K���:�����^i�J �8N;�
��)�C��ˇPt�Aט�PG)QQt�[c��������AC�.�:(f9)�N);����N^��Tu]@ҩ@"4�R�1!*JH- �
	��O���S�^@/����R�I.�̑>���������乔KsF����Xe���y$��ؐ��K�ْ&R^H�7Z�/�����h ꧹R�q���gv
D�\�fR$�n��:�섳cuMP�'<�v0�2F��ԉWYٕ����r^P2�����f�PܓF�՛i��+q�`b˂g�H�Y�S�|�t�N��-�v��eL�9I$�y�̤^J���Y��[2	��N�䴤�w{�?	7s��.�PE$��z�{�$�r�����˺-�$�HWta�	/$��~��I6n��~��ym�� �.(��0t�:u��s��)$Nsmȏ<�I$��]���5���$|�K7��D�Z�je&���g�wt��Tr���2Wc53r�������2�I$2�-L��IW7d��#�]�`��y����|�M-.$��pNe4FηN��P��T�l&ځ!���tڴ#������R��/�[L1��]^)���y� �ZU)��J}�G�<9H/���ʾGq3�39)&.�束��Y�����n�'G%�݊3!$5͖�ҊIz��%�+�r�l6�-��_o���d�wV���h��Bm�9�BXMb��&��g�u936���>��֖��]�;;�\,��y�$̤�	m�ܴ��HW7d���W��A��1�	�$��~�2��*ӳ:,y��ƨ���|�%I�����O�,�I$�|�h	����]�ē�9���n�b��3&�eo:�Դ��:��o۾����՜�"C�RU���v���^`�$�K9��(���n�i	 E���f��N��g>���"��\�.�PI�̖�$�K�����<�Q�ԦRh�\;�t��g� �'���$Of���&T���D�����D�[��R%.��0@>���jn����$a˽uA��1�W�(ɛVj�͗��6��k�?F�׷x����"cۅژ��Z)�@��E�`�D����� >�4 � R"D�@���o|;��������;l<M<�"��Q��i����s��V�3M��)�&R�+<�A�N����OS���FN�O	��%Z,�ȼ�-��Vڮ���Dn��(���҄�u�e�hGdI�V��x�8����K��_CA�����Kc�Eup�%�ܷ��;6���pm4�\v���2����ŗ#�C;1u�Ξ+���2��
Ʊv�桬sN�m��F�����t�]��|~?3�frJL\1�_��ڦZW���qvD�D���F���"q�Tu9.ֶt��`�N���nKJKފ���	g.읝�+�n�踣2�Hc�\�mW3L�I$��̖�%H�dF�I^�"�т�:�{�ZvgL�o;��X�X�D�s�>H����=}�q�+����[nKJH$����^�.�]�`���Ϊ� ���d��Fp�i��/$s�밖	g(�c>I$�f���IV�Y�d":u�]�7q�%{�-!$GL�fr�&�K��L�K�$���P����7�,��3'�f�;���K˳#z�1I �z,̦�1�S(Ԩ(�⋗!;�g^s�X�s�������h���K���P�����ۅû�;�v{����d�'s_�I$����IGC94���ډv��k�I$fF��Ռ]��I�1�)GK�(%>��ry��%��DTvSEdHS
<���,����������{��zU�?�I��������S��|�rV3m�T���m#&݌�~x{�������H4#@�>k|w������^��e"R��,�"QI4B�}=3%��y~��$�;ad�ݓ��B�.w�S)�����JT���-Y�1�D���1H�W�IV�Y� ��6�ɝ:%���ec��>9T{Qd�ɯ%��j}(���cт`$�gC8a�I%��J@����]�1fvggUD�s�yJ	 V̉d�5I쫸Iv�Z�I�,���5xR)+=Hזז}�ɺu�
����U�+�c7Z�YCj�
�״��\ŵv綠��x�m�9����:L:�����O� �	f�܀Ҽ� �[�/!-���lv�ƛX��I��fd%�szq��tC&vN�EQsѰ���y���39�WzQ)%��fI����\�JA-�=�$�}(��Pv�6,b�22geHJz_LHI ���I#���Z�����G[�iy�&5�e�"��	�p���m���X$�ѸG�ի����ö��_�^C&��ı�� ����@�� x)
P��bP!5�~f��K� ٱf}(��fj]�K�I>�XY:wd���W�P\�R�v<�#Zλ��Y�̊3^I$��ے��	%�����[T����Lr8�[sfR{���3��[��&Wڙ��IX݊}*):��u�f&�$�цI�^�r^BH$��~�>��B�1ZNO�Rp���NɃ��\BQ%G/b���������y��	l	�� ci/�EܗffL���菳��^�ʔ��l��I"W[�)BYOj2[��-��&G���w>J>���P;���:L:�-�ڠ�J4�t�nkEf݉��؞�N�����$O3vDb�D���٥����`�^3
�g�2g,��頡��g̐M�G��JA$<�6C�T��f��5:3BH$��ϒ�� ;�ؠ�f�լ\&v!�giH@(�h�M�_�
�m!$z�Ȑ��H��RI2�k�G��[�۽9�-��!;�3,v.��9��(B�_�i�j�r��->��wy�����tm�F=u�8�Y�&���I
�.�*�۶<�8k��1��~}�?D*P�4#H��G^�a}�����L�靝�*>5^_;ԩQ$����	��k�����Hl�ԩ	 ��n� J($�mt����v�s���������V��ZO6�̆5����Qg�q��7`wI����Z��i�������|�)����û˞ڦY �J���BY��*��!#��z�e��c	�~�)'f`�1H����I�33�;:�����L��s�Px�6�T�Ą�$��n(��I]�"D�MR4f�S`�ݛ�Ix���;�N���)y�~�Fy��nہD��{V�2X$��]1���I���	�����"Rǜ����2g,��.�OO<�Y[Ɩ��8�	�:I(��R$�K�{���̕�c��#�ff	�H+��Pg�z玱tY��8c�����H2��,�ǂyY����j�$��*	��W}r �	 �+�"I v5$��!��|���ξ+a�Wm]O=�����r���X�m�,�����iF5��h���9i��ɚ�!��Rh�T������ �D�D9r�5�K]!ڡe����G+�hnC��� 賆�m�]��]��'\�u�S�z�hzKnń�e����KMlR0���,δ���-ٙ윺��m���q�v6�j�v�����e�n�B�M � ;��cY�i�(:����)�G��ɩ��%��/��NI�V�WO9�d�Q�5��r���^0�x��p�N�d��-ݶ)Jcvn�1���#�b��Mj�`wf�=�1���/��Y��;;�\�6}�7�R�H%��d���x3䪳�Ֆ�k�a=�J�(����2��Bn�rJ�	�|���	��^���d�� ���-ڲRI$���L��Uݑ&|�K_�+�!��'��"���F- �R(��������	A$�vcĄ�D�nV�S95ӳ��RI ���H� �]}e%*�����t�]�@������o�*�#Tj�[RA+�ؐe �I{2�$�����I.��\�|��t�a]LșI�,�����fz���yRA?��e�ۊY3���C)'̯$�vt���*��$�)%���ף��~G~;�s�qI�Z)0U��<�=X�;�p$��G@k��X��}~_���E��8c�����xD��̭x&|�	/��S)nw���s5��>s;{"	�C��$�H6�N"�Ι�݂�
��ޥA$���'��k��lx���[�/�
'&�n缫Y��w��C��QYOa�3z�3�JQ�V��4� �Uzr]�����ε��ٟ�`Z�
��_3�>RK�!�]d$�A}o�&����k3C��X�O��58b��+Μ�>捈&�A#X��RI$��5L�������pA9䗷�bL���=m|�R��!�L���ꨀg:a��ve�w�18x$�z�x&RIn5�	$���r�|�u͋�Q����y��$�1�Ǽ����we/*5��	���s �Ta�5yd�F�M	o��,w�S(���t����JD6�T��a��\�-�.� �ҹ�n��,)�D� ����G0Hj*��M̐pɜ�3�r�ƙFR�Z�H�Ix$��\��%9���HOf-��|�>I$���)R�c�ؗ_œ8c*B]3�"BN�ZOq����n��I��x��d$�=��&QIMw�^:n�i&�o	�Y��;��T*�nx�>��A#���) ���U�Z�5s��¸��}f�M&��_n1ɕye�z-��J{g�)D��$�`���l�X��^=�ol�j���"��$p |�|ە�E����R%��>�0[9�f��;�W�9��מy��E��xU\�I&��R$��	fc�I$���K�c*ٺ��SO��Rp�Q�&gvN���Wkтd%���>I�׉Ȕ�1D�Cݯ���	%��fe�z��5�5�Z�U�g03����e'L�ܦs�Eˢ�c<[�ۛl%�q�OOfX�8��*�~~�_���WL̓�.~@F>�)y$���R�GȤ/z�L�Lb�f�U/.��S�@䒽سC^�I��3���U��)�L�|7��6%�Зv����U�oBD�\)��W�	K5�����L��R���@%�g[��f!��v�-��X�,�4\g�Z}E$�Y�fQ%
) ��8�;:wwv
�P\�R��a�rڄ'�^�)I ��ˉ2�y��\�ؿ@O�])�\��m~�!�[�7SW�nT�j�T�R����y����ڗ{6no�lP��z��D,w8���e��2�兄;� ~*(� �_ffg_7��գ���gˋ�tJ�3!|�O2�	"k�S�A��3�1�&|2�$��$�/�$��H]oاҺ2��y�+wH;�p��31���7'�X���k�P�/�0�����/�ߥ��̡�fd��_%ׯD&R��x��H��߱L��T�.�|����`)̋2%Y��&R@B�G���3��^B1�T�Io�(����RJKwq��H��݊	&d���,�v1����f�,L���:d��4�a�dK� �kn(2A.�4�����k����>�@l$���*BK�%����u�����N��D�4h��芺笒=�(��n�dJ	!���g�$�U�֞3�ݥGR@K��d?xN&NΝ�ӕB�k�J�H$N[u�M�a2��.�%ݲҒHֶ�E ���=�4c�>���o��o���������������QQOq��15�U!���Kİuk�?]�`�"=�vv/aẪ��Ƿ�썞�)��sK��s�׶#	����Sۘu+!��ǟN���0�ڽ�U��x��ч=�+�	X<j/�l�W���������c{����{כ%}�g��w<�ɵ^tX��[1����{||��h��>��=�ǜ��z��y�{��v]*w�@<�	�-R��v��K�?]����{�W��6nk0�gm�ӘO�1���h�)������%l���"�/-l�=�,/&�/}��0�N{�;`�4��;�T����vnD�s;h�	�3_��f���>[0��;*�������;Y�*��/��QZ^�},��1Q����[4���w�O��=�'���gH*���Ǹ{ ���s��%'&��
�E8P�B!�śO�H�C"�i�#uV�Z�s�t���]�����{^�qu Z�+�(�;�kީp���Vܾ,��ӟ���N/'�����e)�e��X�.`��X����~��K:���=��u{��&�՛�O;Ȅy&�A��f��ɑɒ��Oq�^�:nὝ�6�i�웾�������qǓ��BL��Rw��/���W�_]z����b��1T˴o3�zk�9m�l�8�ۣ���_h�4S���3�b�J߅����\��=��'������y��L�-��ļ]���z�Y|ΝƐ�L��֜~�:Q����b[�vo��t�D*�ͧ:�.�ri�v7�ں�������O1�o��F\�YY/��������g��]w�gZ�e�]uq�<F�(
��]X�KL�$T�QMq�!d�N�J*H$���tt�%q��rG�wG)�a���K���Ӡ�(�((�Hq"Q:E��gV���wvV�!Y)tDPAY�I�gG���#�tp	���t$���;kA��	圝m�{g�t�9㒃��rF�ٕ�l�nQe�f���p"��o7I�rA�ebC��DD'L�Nf�v�$�δ�NBt�ڳ��裠��s����5M����\c�q�G9s���<��M��z��y��s�)m���t'ͣm�bz���s�]rv���ran�Z���๺�v��k�9.q����[W�\nz��Z�[)Dݶ�Km[�s�wL뎱�g/'��ťt:[�]u��J��.��9�p�b�:��=���R�IJ�GYHLS�Nم�zܴ�7f�����V.Y)��Ӌ�V;'#:P�����f�7�e�V�<�Eƭ����6�Zؐc���gʖ��liIf�3&Lَ���Kl��F���q����.�J��6�b��+C�Csśn^�x�x�t�oe��z�^�:=���a<��O<v
��|~1�$�m�Q�ٱ67�ڸ�q�(+t;����=�����'Q�s�������ڮ�8��J�ۍɛM��n1A6@/:ДP���ț["�\rm���;��[�v�GE�l;���>�nP��+1� ��z��%��[ft1�7!�0�3׌�8�
�qƭpn5���K b���4hFy�[����ssX�ˉ.��T�X2��Ĉ]�9��62�:2S[�����
���݇��9����e��X]QFؚ�fv�th����Ÿv
��P��&�K�= S�W\�5�wh�x�GF��7V�cax��V�-�5�
�������l���9���F�J��p9$�d๻�k̨d���7h����u�Gg���j�m^��4�j]�e���kq��x���hF^j����i!��>��]�X:���۴������P��M�qЌ�d��Ź�.-�T��/6�Iz�)J1-Ԉ@�A���B�s4�R�sHc�oh�Ѳ��G��{���9����s�,6��@�(�+(�Љ�XYI.Fe��f7kLR˷5��@z�eXk���灡0�*W\Tm����
J]k�����9���]Ht���&]�퓒](��p˖�Xb��j=E��%�{It�U���o-��Fmڭ��iW�8�.6^�;x"��@�����{��o����Z*W�"�R�6���u��lsM��0O*t�������T��a˧r(nwWH�&�`�F�����Z�b�l��/k�ĉ�nê�{sf� j�6��ā���p;�v�nl]s[ɠ������n*ˋ΀�.H�m�T����vE�K��S�K�V���&�\z��힓�-��3�G�l�fh�GM`��2�42l�G�8H�c����P��׌����b�k3�g����@�ŧc_�S߯?��	X݊e/$Msu���V��5W�滖��H,��S)�Im���338u�r��I�_b�`gvuխ���$�KٯئBK�%\�je�,`kv����P��;�����K���R%/$Nsm�J	/%,k���Ҝ���w��$��k�($��~�[p�c��pSL���-<�h���i��=jI�qA��	X�j'� �r솑o�s�]�RAn>j� ]���܄�1�)F�촒��b���o1N�/��%�ݪ%$^Y�֦Q%z��%��ֺ�� .ʔ	�-���V��]�e^9�s ��1����	�i�˰#x��q:vt��Z�c<���I���̽,$���-!%*EQ���z��ү",�$ʬ|�2�|~L��]�����X�d:IN�{�K��}������;*�\�f!��Cb����ʕ�BdA��*i�4���3n�c�	�t:p�z��<��T�<ovSV����y?)$�����$��o�Z|��Z`�;޶f���wn�B^w䶈N�����:����mO�I^	g,Ȑ�$L�+�욂R��{8N���|�"Q^IW7d��S
��.�3��r�Ϥa�
�2r�$��[_Hi^I$��vKHH����0�����S5r�T�T9�0t��3J5ḞD��[qL�כ-&���{�2�(e�d��� �b���~o�|�������3�+t ����؇)��rWl �LcA��ֺ�2o'�~�wi�9N��D��Z�I�[pǂI%���e,l�fY���|�2��Hu�䴄���;��.�]�عT*�;ԩ��K��"5�hI Wm�-#���߱H�I�����������Ps�o��["���NfV:��K�e�b�I"@>�1��S�a�A�4/A�bU�y�3YY�2�Py��f�e�u'Ȣ��������]�ci�����i�!
6'��Z�So{{j�սԯ׌�I76�2�
��ߩ�f�!;1fL���
�K1����.�bq&u�g�$���)�%*��K�[{���[���J��������.�0L��^B�~�>��I%�ےx�M�Q�X3�}���ՒҒIyU��(���~�"UC�&z7��=����z%�&�������:��lsnH5M J�v8�UI��{���C��h�ӧB���tϝ �K5��(�䐭~�2f�Z���W#�<����^Iy]��KV�����N�ጩK����%;�#S2��V�L��t�M[n(���Km�)7l���٣�y���ۏ�z�	�D!�(�J��n���RIu�!�]�Q5׍�H����"QI����z�2�>Gk,��W�<T��k�L�XA'ֻS)$�C����H%|��>U�y��M����$��/�"���l^)���۹Z���H�/�.�.�m��Z�σ��G��8�R�ڋ	g�~��#��~� +��͙?��=��JL����ř33�UTU��!�$��Yp���&�Oo�||�$�+����$��\"q��㥳�ƛ%;1g��o;l0��:��5���m�1���;jʆ^���l�b:��	�gwP��~�"R	$�[n|҂D�{�r�![�Ѭˤ��S���Iz�je �e+�Ɉp�:t�U��,�M9;F��J"�Zy\zY�%���d$�Y��
@I ���KW�r��_6�H�����N�ጩKe�TO�'s��d����^�ܞ!2cU����	%��jD��o2W��*R�F�N"��ٓ�*�fyUûz�T�x[�^:�"o�CJIy*�k�I'�����n�V�Yd����y��3Qg)��^d�N�4��2$��L���͆Ȏ/����zn�%osܢI����e8>^W�ŷK�4c�L5B�MdN�����^9�v<�O�9b�c7y�|�Yy|��<��괢:��n�n�ǳ���@'��;�<;E����.��#`0L|��]�R�BB��F�gX��a���hK�ps��XK
`��2���<�$��Fj���7��P�$KpjSPXcgX��YB� m,(܍гv�!�=�W�����'Wn��u��fˀ*�,�
B)2h�3��6���anV��p8�ar�̈́�8O.�\�m.T�ˑ�b�H�B5��D��@u��a��5�cM��f^Y�����6M*ݚ�Y�|>S���D!(�n\�'v4�^NH_���³�l҉6�W�o����%L�3�_O�J����PK;�Y$�I��S!%�\��|�
jB�~�"QA,�k�L¸GC�p�L��\�6r�)x$�seq�7z��fsv�JH��Ʋ$����Am��E�8i�����r�H7YJ��!�`���P��!�I%�ת})�I�'�ۈ}�o<�Hz�=T�RA$/Z�$��K�0���o:vw,eHKe��G<���䐶g�j�d�%ǼS) �m�����?�6Wi����ʞ�3�vN�ܧb�U
<��R	X�rdƛ5�v�!��҉��q�P(���n�>���u[P��q?G��k5�k"�j��k��ki,���X\�*B�<��ªF�������o�0�[�5����Ʀ@d�A*ƾR%$��]o֦D1�W9��d�d�F�J��I\�����$]�L�3�UT�cuH+�W���yT!+�=��(T���%�Y�FclR����M#���c�2��t���/��1����8jc�u��Bɦh8*�ڎڦP��v%�K��|�R@$w�H��W9[su^).�|R�����: �:e/*1��D��ܦ�I ��|О{gj�J�Y�8��C��H�W�z��I��j
�)e�LC��ӧ�����{.�>DXō���U�v��)/��S)/$��=�||޾"���WT��	���Zw��p_��N��	bT4m��A-�k����R�m�q���Hl�Z�I33,��R%Hns�ɞ�K:�Ԛe�1J:�W4[-�k��WN������8��gCۜsS�)��%�S���\9Z8�\TO��u�c�I���1S69��{��Oke���1���ˢ<X[�S>�w���٦�� �k[m��츒M�����j�%F�=�˱�jI��2g�L��PI콸�	-�쩼����Y������u}�gQrr���ٔ����4��7}�ŚtT��g`Ў��Y�<7��Nȯ����v�1��2��_�u�A<���G�_fH��プp���`��l���19�=�a>5+��O��	��ܪ��Λ��<X��*���Y���K�`��`��̎�ݙ�H=�7"J�d�l��@��-9⩯nd��M̦��:�7�q�=B��%�xj�.�bZ�&��Sn�cl�d���Ϯ�%WYL�,Q�p_��N��q�3��y�q$�N�M̗�(�����dB��	���T�2�L�p�H<ӓU�ٌs�ܑY�Q$���s��4�.g���y=��\ӹL�ˢ<�6�H�	���;�^��?A1�8�^$��s>$���ӑA��S��&ffp�-��Rs���q��fv��KC�ĂH;y92O��}m^>��;昆���hqV�ހ�Y���be�x��M�1��*�Bk�3��h՗�wK���u�_۳ �����//f�R��G���⅗/i����Oẽ.�,��%��(��V̂ۇ������;��Ή�$�wzp��,{h91���_Z&U�Y��e60"�k4Ƙ�IP۲ًZ��uhq CWr�݂,S�t-Z���L:}��$;vr$�5_[G���W��M�T�X$��Ӓ&����Ho:L�Q�4�U��'�����GT̼E�$v��ω'���*�ؽ���i��8��p$��`���<ӓ>�	ʎu�pLu�\_�Z�c%��hI������	l�i�&.���dctT��Z}X���7ӳH:o-��e������R�0�ޙ.����0A���Ӵɓ�0�ě�ۉ(�:˺u���O��nD��2�	��\����Ϲ<ӳoj�M�|ǫ<�P1�u�4D�bh>B���S�C��^/?m�o86�|FmH�f�4�g�Z��&+L]]<�]#L����%��(��*�׊]&�,��f�\zҵ,�-�\���+��.�1�R��`�ٻU˻a8���)+I�FM�!�Hbn.��ٝ�т���s�[k�0��Ԙlq�d�m��r���Wl�\q�#��(�Q�̬��0��M-�Z�C�Ù[���6�/��ۉ��s=��m��rV�j,����-Z6Y�fa6�<�yXhӶQ�{�!s�Jfxޣ�\z�^	m�{R�����H�wY��pr�\"Y�2�����;���$;�s'"h�!w�N������A'ܷm�WX�3tSN�g�ϻ"MW�l�������.tO��}m�˙� �R�g�9�ƣjv� �c�p3���;f|ʝ�$���q> �J)k6�����"<���A5��2.0h�	�����h��d���%ؽ}�Q�$���Z���g�6��;�ہ�k����'�Z�|I>5��9T���\�U� 	�k�)� ��^K����T�;�on��%� g�o;'��V+�.4���n8�36S:Z�ā�,k	����bY���b�d�ܻ��P�Ě�ˉO_e̘��
�M�z��Ҡ�D`��q3�b�.��%��(����r$/nJ~������ǯ�*P�[��ޞ�]Jը��s������f{�j�2u뗎��)z�1Hɞ���g���I��UF�$�M�m���s����rdxھi͙��P�M#V+���ӻCwFƀO��r�}�T��O�`W�#��I���I$�˙:�N`g��;�=Aq��|���ȃB@-��I ��˙����"JJ���s�؝�	��ɒ_�+I�	0N'Z� y�.}'ăG:�;�_grӏ�@�e�H$�w�s����h��D�����w|�i�&r�;�k�zz��n9xձ���ǳ]"�:ʗX�6�L�g�_�,d��wI��z�*�I^�T� �U��x��IV����d]�T�H�D�v,œ.�ݪ���>4��Ƨq)��O�� �H'���I$r���Ѧyz��o��D3��H'���ܺ �>q��s�wޱ�{o}��%�3�nߏ���o�����{=��_��f��)��h�={��f��W�b�;ſ]q�'{!J�u�j*4Q���0�:��/�̉��dԳ����|��<}3�<�Y��I�v��%�J�9��>�Ҟ�ܻ���w������yyz[��o�A��{i�w��WuKQK^���v��<l�a��C �_�=T�-wǝ�pɊ1wm����ϩ�e�=x�{)g�UPC�x9��
l�W�[燻��B#G�YJm���v�a?vy�tz8c��3U�'7�{�f��==&������o���o��Y[��PK��!o84�w�/&;������x�q{@�� ϐ�1���jԗk���X���>Y5E����E��#�"���j����ǃ��5�B �ؙ���1<��ɞ�v3�w�ûρ���.o�
njYn�>�f�*!b����My�ھ�-�b��������sg)�v�Y���|�Ǖ��D�u��LgU��py����Us���Wu��������D��sCRz�P/ w�%�6:�t��`w�NXHQ������ǌ{|�+�)�0[��D�(;�ܹ�%�͌#�{�y�y�E�O����)��� Y�gޟ(3t��'���!wef�cb4��1�/w�g3�=�Ъw�u;yR���ϳ�N�TG���e�;}{�&��$��9v鞔��\<~Bʺ�g�����94�fF%��,��K�2�{=�Y�bl{������X+E��{��ٺ\e���N�q.���ǽ�-�7Q���uG��r?�
�<=gwn:�����+�0`ƒ47�sD�%�l	�$#�N0I8D���b���I����p�8rXs�hn�$��Ԕw�YE9�Rw%��Bgbv۲���;m��QV[km����E�R��B�p�����Z��r8���s!S79NY�C-�9��e6�')9�Y�$�nr�֝h�G:&ۋ�:
p�����E(��&gII�M�-���f4;mmmm[�Dfmkk[n9lݹYnL�Nsm'�i�n�rڶZ��Tն�։GSnͳkZ�r�[n#;���m��&q�wZ�3���9�m7G'm�貲�쳍��H�H��+����۱�_x�M��s�9_��
ы�`Ί`]�D��ge��{��II$r̶�I"����14:Q;fd��t�pX]3�*d���H9�� �1X�le�'s�$	�$�f>\�k�Ƞ�z��DA�u����q���`΁-�M�2kΕa6-:�A+�M�z,�S�ՅӇvz+,���-��>\u�vD�H�e�$�]}s ��R/I�7�\d���� �=X�j	E���b�� Y�q��dYc��j���p��ڬ�$�|2�-G�$e�v@�D�l<a���?���H�ye�f,Ⱥt��@�.�A �ndH$��}��2��L������{��Ż�|�O���2K�|<��H�YHmݫ�l�����>6ˢ bI���	=}�{.Fɶ�����"��}�u�{VN��w6.��n�7��w}����_���r��4���e����R���9�4�f�B�)��)�w��8|NCn( �a��f�&	�Էtl`$�w.D���0�����A<��r��d�6�f��DS�z4���v1�u�㔃v������*G5+l�l�uX�9'g�lA�݋��+�pg%��8b���Sp�w/�$	n��|y8�n���[�N)�(�ۉ$0��b�0v.ZD�g��'�a�S!>e�2!;�I ��˙���ϤH4��]��r�����ɨ2.��q>�YY}r$�MzV̜/[uGC;ۗAw�	�d�EئEӧv�2s���ŵ:��=��(��tI>$7o�d|O�_[(Ǉl��6�6A>��ْ�_N�r����Q ��\��;�ڷ�lŔj�+y� ���	čW��@�Sݹ���q��Q���L�����zZ��,����&<D�f�p��*}8��a9��@8;;��/��K�����R�?W�q�2[�{<ɛ�ƨz���ާ1�;3'rZ�MmG�,F5�WF�
�����b�BX煍K�5f,N/>���p��9���v�������i�lv��b���qzy3�]n���fǓt��c�n�R�<��Rh���gJҫ�B���-o������T�+�aw���u5�ۛ�C���]�W`8y������Ѣ��Fz	{�:�;uF3� q���ru���Ɂ�Yf�u�Dn�)�GIoY]�.6Wr�{[��v{�o��2L���'ߟ�6mt��$�}�$�����<Hwve��+wn��$��y���03���ܱS ��r
��֔C]��ZV:�5t�Ă&��&@$�/s_[H'���N������w���V������ �<� �E��W�D�C�ο4Tnx�o/rd}z����u�,N]wI��ڛ�#X*o9�iB�O��̙I&���u�l�]�.��ρ%�wg��A��;b�:N��2d��9Vv\H5���zGb螮ޙ���j	$]w\ϋ�����O��V�d��[�veT����6C�Z�Ÿ��u��K +������w����E�!�)Ox�v\��jۆ$���&�mv�އSpʶ}�-ʻ�*|P$��P	����X0.3���vvd�z�'X��bZ=�b��-2��&KN;�k��B�LXϠ{v%����Hz:pX<:�"�=�L9e�C3N����%��5e]�(�t�~{�[�A���P	�}�̒f�ª��H_n�\�pm]���(:삙�N�c�|�uĂA ͹�.%ɥx���� �\�j	���'ͧF6������><�:�p��#�]�J�nv\�$�v��J�v!�5� �n� �z
�S�E��D�̎��Y}�A�1P�;ۦmn�$:�.d��D�dd�u׎!4���/wg�B�(���֮�-�B�Ǹ��O�/�m���[���?_�_|]8r]��fwg|V�c�A ��\O� ���Cn�s�E����˙ ����ܖ%3��|_3�du�Z������C>� �3s.D�O�]�Ǜ"�g&��cC�5��,��p���L�t�$����� �w;rF� �*r�x�`ic�v͗@�F�+b.�N�U�o/b{E�߼�H�k�z���᥽�}�S�w���Xu\�m�?+4��Z휿�O��Owm��O_�q:V``�vAL��;�[�;�zP��%\�D�|I�nv��$���X���;]ǝWut���Ŵ8A؇jR
����IV��j�g�h���2	o7.|$zۭ@v��w&\e���
L!.�k��nŨ�pL	m�܋�e�0InH�4\��*�����ftQ,�޶���I ��\O�'���%��dH�[ϙ3�A ��\����rYݑfwi�8�`0"�
W_,�ۇ��7��2H$u�Z�9�ƍۦ��*���lY�`S9JCom��ڶ�1�&Q��w���f1O[d���̂;���P	���K33��Wll)��RĀ_��dFse��$B�����	��5MLN%*��z?��f�O��x�k�x�7�~:�J�]1$&v�v�󫿇?�|7�����������<%��N�Z����w�ܖ��-ϗ06��	�A9wd��a��D���x��|*������$�{mG� ��}r�_Kr*lL�D���{v���=u�����-���5���(=�� �NS�D���J�p��|j"�I>5��c����~n���S-���h݌��oy��$G�5l�3'b�g�Y=R$�XU��6�6���h���{0	$��$��n��XP޵�t ���.q R	H����0����`<Q��z�z漲I��`A=W�2	%�d�0)��!��v�S��&�����t5�D�n�ng������1��z���Wm��$vB��d��g.��&_��d�?���Ȉט��{mkt���=��{s �|v��@�^k������>���HBz�<��:���x�� �u�+O9�7�x���4���a������<>����.��g� '&���hQ ժG�A��K�)��tb;\SԮ(CkU�z�ƍ]G-�=i�Lk��B{'\u�����Y�DШ��WH�t\A�N.���q�t��x��7jSr�%���-�p\q��;���P���f؋'*��	�"��&
e�R������d�l�Inw�/]Bm�s���g�G	�#�[Cf�1�猵�\�N�:��{8��i����?|��y��<Q�Ѹk��6�8P�Ӄ=�$�ݟ]n�V`ɷY����j�8NJ	˻ ��̶G�'2��H$����D��Ҫ�_ Aݗ2Hm�d�J�p��D��9�������4G�2�I$��@�e��������A ���4���#@*{_�� 0\�!y#v�}0�-ޮ��$�[�s>�_S�nܠS�%����d�iګ�]�Te�w��GvN��_��m��	\�c��뵒Pz����z�A D�����&vJd����vcT+��22g�"�4<�تȢ@'�w��k��f_=}��K��=z}J����M��6������Sc��X,q��:��%pʹKew�oP���o��b᜻;����wv��'k��x���M�ݷy�� �̸���8NR)˻ �A���> O��-d�6�v�����^G��Wz?̛���~��;���,�.wy!�7g��.�o����qm�!�Y	�gq��v�r�i\y�����c6#�$I�ǂO]�$wv�5t�:CS<��ƹ��(;8A�����:��9�P�n��sQ���Mf�č�z"-�L�3'b�g�/=2�5u:~��ؽ�My=�<�I^�Ǣ$�յ�s�ΔB�� ��@���@�)��33��9ZӞ�1�n�� ؝.�9-�`O�j�=�A3��D}�=�r6"���I�w+�Jb��ݓA�.����b����a�-l�Iv�|�����1I����e����D�=��%{�W6;��/~݁3Z�c��k��"����dc���$�������*��w=����j"<O���D�Xl6<tw\E���'I�ݒ�2[!gs�&�� �^���[�S��Z�Ѧ�x��ȿ�L8Fyn�#�f�ۖ�{��}㗯�ag�я�h���q�v���)�-�x���v�[�$/5����H�}X���3��dx��Jn6��˿�ag���I��!�(���f]��U�*;����f#���.�]�;$<���L�I�븙9UFj�9��`	3{&A��\���k��@�.�� ��s�kFE8a��9:�l���uM3NuԄ�alu[���O4G{���ܫ53�.'ϱ嗍R$��dzA=}q�v��-�Բ]���$;�2d�e���E�ҙ-�qʲ��i;�7���ȂI��ɟA���4
��`� �呾Y��EtY˳����f@'�������Fgg旊[�|�~$����$����1�Ӣ��$�ݒ���6f76��K��D�O��ۈ �;�D	�al�T�N�Qw�,�� �K�޾¯i[�R{�H��v�Z�L�Q�(�8+;Ѝ�mU��>5��*{�绕Td6K�Z���<��l�L���vp�;8A���$�>�FW5B��Yу6��b��*z�d�H�#�w�P�^]�&�l�ك�"
�%-�I	��6��%`]�.�����,K�)�	m&r�O�~�߸qgb�Y���`s�/޸A$�7R�)��K��f�+�I�����ݸY��&gJd��|pN������'Ăo2�<I>�� �f�˰��\�G`'��2�N��"��H[�pA&����Ap���v`'Ĝ̸�z{�����LJ�3�gyYѰ�o�Wv�c����v�"�>�ף荭���i\0t��-{,��	77����tS3$�3�Ra��� �_dO�nwtd6��]f�""<H.��|�tQG���5�������o���^�{=��_����
���F��i��ʩ�������$�'�6j�3rm���3�2�,'�w�)����t0���]D�ov=��ʽ`�}���V�K�	���{̺�ok������*Z�>4y9ꏖ�yV��5-��=��r�,���$�`s*�.�sذ}.]�w2�z�����{��(���C��i�҆w���!r;i�_v���ڽ��+�&9���;�^���2���� o���!�]��9坢t�&��j��ѧ�z�=��u�n�8���Z����Ā��Y�'8a�j~ƹd�%��41��=�Vɉw妷hC��յ5���:�N͓Sy~��*�\�d����&q*�X����Y=%�N���}{=�G�+���[7N��5���v��&	`>�����٥�C�*��l~�FqM�ߣȜ+������H�����K��q ��	*<�m�َ���Ӎ�f���A�0�~��q����kL�V&�޴f����3��#� ;;�^��sӬR���w=ܛ����MG��~y_���֮�$�s���m�{��w�ذ���Ai�9��A�����:�x��D=mVyt�aZo�rr$���0p��K�}��xo�ͤ���J�2/,�����7|!�g��t�8`�s�d'A��Ih�f5U̗�[��U[1n�3����Wᯥl�̋���)�݆{��9��hl8����}
��*3�{<��=��{��ש�N����o�]���]|�^��g?�{<A��}ׁ�3}�����(�m���n����-��D
j��v���_\-�&�f�?�?0�j~�ޅ����P��SM�k����6�Gee�6�2�[q%c��k�;,�l�������ݧ[k���Nrӱ��ִ�m���m�6k�Y�stDŝi�asm���#cY��ȗf`,�N�8����f.tT۴����93��6��J��Y�e�m�NL�Ą;�"��%6��m8RG��gnPvVnYɧY��F��M���I��f�7�7lB-m�v�`�a���:rFщ[k+t��m�[gZ�dݭ�3t���prH}�w�Ne��1���f��;0u�n�q�+m9�l��f̹Ŗ�5��f�ZB&�9,���ٙ�,��mk�q�ۭ��܎ ��ZM�6ț���",[�gbru����'}㧟��~͝v��Z�AoA�7I�n^��Z[�t�F�h�lf��pElI�hm�HR�l�JV7�Rh��;�^J�R|c�vv'���ۤŘ�X@�ꄰt!�B[1�7XmT4�t#j��	,�t�_駖_'���6Hus%sukW�9��׈���4&��L�Q���k�5���2X���1���Q^���щ:GX�N	y�f�S�ݽ� i�/,�])��\hHO;B{s�lW�����;nr�uQk�7㋲�Y3�sW2i���
.M1D��B���WS\4mŔ�vZ����Iq��Yvm^�&�6�e�Gj���]��nw��6�(qm����@�g��ª�\�{H�4u�1���b9%nĲ�^��1�@f�K�v3���qqnC�A����v�7;����ԇZ�դ����y0=u�u=e۱9�6��ta��!�"� [Zɴ�a���ėK�RK���u)<�T�kXhX2n��[���ҹ-�u�B�-�<h�mKv��t����ȣ�mXh�6z�������٫	�I�Iz�b�ʙ�8�3;�J��c���ϥs���A��3�g:��Q�=v�y&wZ0G)Q����3�*;�L�cQ	���)0r�v�nݥt�ku�f�Ж�XE��[+fM*p㵳����<��s�k��k g[�%h�x����h��;A)(86��kԩ�!ϱ��Q����G��[3�\�E�=�Ƿ(�d�3kia6.��fbɛ���¼nl><��Ց��jٟ[�]��8_K�9z�uye�!�kH1����k�u`�n���Y�u��I�Z���,���0�����;fp烊�賷<d^N����켌�.�oL]�3Fy�Z����)Zk�m��Lq�LF}��=�.��)|���ʩ3��x{1�.�w^��7v�p6ӂ}8�[\lv�]�n��y�w�働��v����ŗY����u��7\p��qV��փ]ۏ%]��۝˵��8cZ��L����15�)ٞx���\��v��X��A�=k��+ċU�۟LDXG�K��=[L�[��������F�
Cq
T�6���"�͚,`��1J+���+o#n\�
�;�&.��e�lZf��;�	��7=q�p��6W��*�^����+B�Q��;̞�٥�R�-���)�Q��z:����L�W?>��=m���n�ӷi�׆��5vi	s"�Kl��J����a�l����WS�Ϲ��vp������: ���DFu�L��ȇ��z���V���z0'�\n��;$��29��d	�`��g�M��H����}�$����7Q}λ~��<(0r��Ȧr�dkE�>5ۙ|H50�]�B�7[�	�woF  ��dό@�%����ĳ�Q �u��Fe�K����AnƘ�	���2	$����'�J���췃�A�]&E��L;��l�ِI>=�P#q�ڳ��.�Hvw���ݓ$��z���GJo���cK�Y��m%�I�^fB�ˣ�[1�N��AA�E�C 훩���}�������޾~zk>�A'r�"A$ϔ�o��M������n�u� 2��w�v��wE�����"|z_#�H�0+O>�1����.���G������z1Z�?�v�������(�&-�T���IC)R�)���<1�P2�1���~��K�| ��?vU H#����-�(�\�z��]6��	��2�3�vN���3�S$��Ψ�A�gZ]�l����^ђ]�2	���<~�vI�L�!2ry��(�MK�ܑf���G���� �D�=��gp6�fx�Q2O��AeΝ�	���U�H�֨U@��������'��3�I5y1 ��=��6[u��r{��V�Q.YؗN�0d{ux�t�z��чf����(ڡ�d0��y?g�q�!0wIçvձ{ fd?u*nz0@�|�y�O'W��^4�I�ɏF��&dY;3�P���%��]�8K�tWG��Ψ�zw����t�lNy�k|�K����.�S�C��;/p �o��H�zS����Kk��ÕA����͂Y,=� �v�Z��ݍx򓔴��==���h4(W���������;�5	�r�d�Lݳ�I�ʏG��=*��d�X;:��&�瞹����j��V�A��5�G��2i����G�r ��Ayݒt�9S �i��&�s"F�6m��C4C�v�O�#b'oZ�{��d�eF�;Q�5��S8d����M�yv)�a����d�;%��2]F��v�+�MV���˗'wgPL��۞@$�cT">%{��*����x��Y��@&�ڌ��N���'��.���KF\ݴ���}|� ��Kw��w_d�'ǯ�-ʬA�pt�u�� g��lŘ��ٝ���1��`|e�G��dKp���Ӷ�>$��z"<	�ɒf�tYӹg �xK�U����&���O������o2d�A��8δ�W'HFMy߆{$�V�J�����������&/g��'{���x1�����2�޶��Ut�Y��*6x"E�=�&�F��
[����/�ɀ������K���=�F>�����t,o*��ÿ����>���[�]WX�TL��Ff��J�!�����G�Z��Q�un3Lg�����4;d%����z��cL O_^D�	 ��<���r\=!F��O=vNtI-<�bvv/��u2Y����|"=��s2��H$s�'ă���e�Q�Zz���8�>��+S"��'%���g\�۳;��q�q��G1l���s��$	���}��*sIHD�5�������_���
犉�i����u��}���;F.�Oqq ���ۉ�2r�Y�!ތ�������j3�y��-��Y-[�2	�'s& z���}�M�0=:`��Y
c*�f����N>���nm8�a�"�7$�2n����7F��L�m�D�:{�
��<�c``}�R��iKQ�����e�6�n'S���s-�t��Vˑf��b� Sm�kt�ѶA[� n4����r���G���4�@��f`�q����'R�;��W\Q�v�ZM���MsoPv\v���aƶ���aZ ¡ol.��kS!55MCY��n�
Q��3�TWX#L,��#��»�yf���Ok�0���y��ݯX3e�<�R�5�m��!t���P�&�:�:q�t97��[qV�2��O�~�����D����92I&�� �z������j����Q��d��옂5�X�����])��lͶ��c\um��FI��x'č�z0E�b�y�TJy��8�bvv/��u2�S�$�j� ��rW�)f�(bТw $��'��� N�Z̓'r�vS#�7$��nͥ́�91O䁦Ƣ �7�����3��n��U~��dY�f��TH;2����D�Ec���D����A���x�w��d�e;\���Y�',��)�v�TӺ�ը���s�H�\J���	��w����N铗r�A�8�=��5�D�O�n�d��V��8��~�	>X�`�~��,�Ju�Z��`�@Gd�hw��V
��nP�yf.�o�
��� u0�~^�E�k��x޽��1�;��a=˦L�NÕ�=b���w��t���<GEw��粳��q̠�lQ���|H��`O�u�L��1��]��h~ʋ��s�l/;�@�Jg�s�a{�k"|O��s+X�S�=�Mݽ� �	��Hy�!c�r肝é�G�O9�ս�
ZyԦ��hh�`�M�ۗ$]֨���J5�������&��fI��w��?nL��[Qź_{j6�R���Y�Ǌ����$��='`,Bm�*)�6�w3](��H:�[�\��P�D���3CAlݸ�víL��w�7K��fv-¢�Ȓ��D��%?�z⁩�3���n��ny�5,n�-����'.���I�|���w])�n��9��Ыgq���>ݹ2	"��dr���fͮ|�7�A�R�\�vt	)�VGT�#/����x7����p��ɒ?���R?>��ۜT����烦���=��&�xS5�C�'����c��o<}�n����E�N���Mv�̂I5�Q����EyݒغL$FsJ饑�Co5��N�{}	��ާ��|H�糊��t�f��n�.$|����俋3�i�6 �f5ǒ˙��͊Y����d�OfT���dva�x�P��cn�o&p_�W0�F\��
S��մ��y�u9����@~������;�ᝒ���A9�P �A����wŹ�{����S� �	7*7�u!�3 �ٜ3L����`D��ػ��*3���j�	3���/ ̤�5��ɴܝ1t�9!�+Ƽg�<I���O��}Q�bfIN��w�I�� �I|�cāa�U�.]�;Jy��'����3�oI/1q���r{1�I�u�H�w�S�y��l����d*�U.����f?�Z�o��J<�ai7,�a��/*X\)��b��\M�sFE=;��˳L���y���wz*�-�e�N�� S�J$�i0	�����e5e�ҹ;�������f	�]t�w������3�����
��G^�BX�Ń<dS��gۗ��kꝒ�����)篧�>]��Z��p7=p �A�Ƹ�DFu�L�X"�n"�OM|�`!��2I��w�O��rdA�Ҥ�壝�	����龙�4��,�Tu��@��w�9�͐Af�vp�2va� @�پ�j�Ka�[M�Y�	�>�׳�Ol�L���X�Ӧ.�%�O��ڋJ�e���D;\"I-깽��o�z��Ei�d�.�41�Vo�-X� 
s7�zD��Η�<��a[���h};�|	�t�L�A>=} /fv�bľi���g0<��e�yI` ���M�y��r�E<%;��t+K��,�����Ƭ�:�0ޜ�,�c�E�`f�p��n57�.Ok���I)��n�n��i���#=���H<t�[cuq��K˟]�'B�JZ��nQ����܃�`f-���������͎��tR$4�n����n&F�fm`Mp�C��.�d���v6�1����j6-.k���p�z�'�61�i�t��r��LY��3��,���A�^��8�˩�,l ���P��]�#^S�KV=�q뱮�q��0j뢜�q���y�!��m���v,Jp�w=�1�As{��<_ۏ���]��]Ӭ�Սo$������Eu1C]�	�8L�Ew(V�nJ�!�ݾ���^eȟ_T@&S]�Wzz܊2���gA�;�Q͕���|n�G��h�W0��_T?A�A>�ܹ�@#o� 念H!��;��i�yl��si���~#2��I �F�Tz=�oF6�o����H��ɟ��V;9t�Ӡ�iz^�&�Z�(�R��@���>$ͨ�o[Q��cc��_�������m���\et�x{h�#Z�hj:5f��ǍKcm5F�I������}-�f[]��WR$�[�$��vE�-����p�6�g��� ����5�����C�ҙ�֘^휕��D,4𩪡�Լ=�z�����3�#��z�X����[ޝ�WN=n�vi�������^/��d���Z�,"+���3y=��u��6z���ى�S�~��K�C$m��,���>/�Q� ��j0I�=N{��e"�{hI�ڀ ;���>�תً;:O6�C"�aj9CUc�fA�����F�;��7w[��H7[p �r8���;8M2<� ��TH9�z��쐝�#ĂEu���}S"��whWv����,����.#�/M�u�m�/m�O8۟Q�Y8y�WY�i�9�2�����c\c���>���[��Zm[���3炲�q��d�v���z0 Xx�h�t�˄K<����TH'p8�=�����<lH'���`Iݾ��I�S���ޓgK�g��^�2t�`�:S �kL7��׹q$�-�;x}v���������������u��Ij{��4��,��5���mwo��-Ί��ʓ�}�pC��ם�/x�x-��y���J>���p�/o�r�:��	�xyu��_o7J�{G��<�)����$w���_��r��;T�۝��Y��h�w�G���7ͅR��q��.:��$ A�
k�69y��C»�4zx�w^P�x��{$P�ߨ���&� ��۫ѓ�xO4-�=�sc��5]¸�X�1�v �r�^��*_���1��9�d�{4��g��ޯq.=7���g�ݶ���T�˝�^�#if�_ݢ��lUvv����i0���U:�xnWk�0�}M־��1ycQ"}�/�������ǆ�n]z�^���<a����������ɽ��k����-~�7�q�ݽ�3�;z�]�=�G��gԎ��M�`zǻ�]]�����5�
�7�ԣ1?��z/�BDy�<z򻋖��[�۸�9B,6�抾{�Ƭ�3��H��K5wM������5!�K��3�%����7����Sfe��v�3��W�w9cTo��yo.=N�Ԟ&�o|�S>���\>Wx�C��=��w�Y�VUT�F:�a��2�X ����W��8��bKL�5�v�?,ӆS�����J5{�v�� Օ�q"t�M��7�� OoNd���Ls҆Y�=w$��2�m���D�n�z5-�twA<��bX7��t����Z)�}VX�X���3x��cm~k���p.ِ���I̻fj�BG!�h-������;p�mM�B,�d�L�r��;m���3�v9e'v�8��!���%f6��[2�'H�� �sN������ڭ�q���vւ�,��:�N%��;�n͵�)kZ%G!2�r s�u�h
9�[�mRRDHL�\�9�� �iH ����[n)�&���[��n!$9#�D��m�� � ��ٴ�en�&�iI���NH�I�%�:�ff!Ds���G�݌�)��;kE9 �,�Y���IM�S�u�$Fm�p✒P�m�;��(Q�6��e�H@iIq7l�E.m�+[ZY����b�Ӌ2�1��6��cE"Qq���
N�Ӷ�vj%"ͰH$E8��3L�BCf�j��kj,# ��"�p�g�5�>�V�o����}�>%硐X��-�w,�%���6��&�M�O�d4B��ܙ$��ծNQ�fd�����}	��� �LoZ���;wN̦}�׳$۵ D�,�T��gs�ߚ��H�}�*�A�;�n�j�y�Fzw��D�I��Sk3f�xeن/=;X��F��tu�"�5�/A��I����~�G�9�&�*�M��D�	 ��5ݮKL-��
n~"<H��"e�:t�ӯ8r� ����I�@�.��r�yC� ���b̙���8ʋ�I=u)$8�NK�p�g�]S+�+:��&�w��L7UF�#����$��������읜�,�Jd�.��]y*dD��*$��W��� �\�h
��Q��%4�A�w�R5�aM�16e2qe8L嚫,0�4�I�^�H��C631n�ܾG$�4�q�^U�?<|}.k�iвlPv����K�m� ;ݲ%砱�r�8vi�7��������t�����Q'�i�:��LZ��pu�wNY�(%X��m�c��mc�-�`�[u�B�WWG`�� ���<�ݝ�g.�0�t]�� �v��'�ηR���W#gn�C�`��ِH�Ω�>�O�!v �vp�g�9F �/R�q���n��Ē+��>$	��P	�veY���8�k�g��m�:t�ӯ8r�$�ǃ>Ae��b	/��y,y�0��"����q��]��	b�b��N"Y�O4tE�WS�NB9���z,&�|�H;p�	;����!��®�B�v �F�;'g��ҙ8kf<�Ě�́(�OjˠMmL@#e0�wo�d�2&�"���ZNڙkB�`�%�ڒ|5�r"�R�%G�-��:�n�����F��� q��FJeM6I`��v�F��յnD�_�2����\g���&Җ�9�l�q:�H�u�D�������z��a-4u��¶]l�`a0����qDi��	-.{v��;���4�u�!�h�(`F�gcsu��{u�7Z胡�v\u�j�v㧵�.NѺÈٓb�P���x�eډ��s';��uk�G\���mq�̯2�qT%���q�m�cB�&�c��0��c+f'7�����#����u���1
��ݥ�{fſ����>F���%����y�� �g2�A#��&A��o#o 4�q �yWS@$.�i��9`�]:�n�ْJ����09���a�`e]�Ao_d� �9���E�eMξ�v`�Bk%�t�A	;��>0r2�F��D��=\��X�ŗ���>$W��	$v�d��ͶX�ӗN���P�����xV(���P}�`!�=C�	�;[�	$�����|8:_-��<��%8p�g�֎��A Ψ��
t�]��	��s�L�A'�� �ӏ�N���e~�~���,�����t"�JٛSZ��`�������Ь?�O�Kp05mr8�߾��2gJ����79Wvd	�����Pg+�̿	�m$�;ۓ ���q܇,�g�dΨ�@^ʉp_ľҞ��>�W&?�y��'��=(�yý1�?�ۻ�Y��EѪ�_�z��P��B��5P)��a�H�m�I��ɐA���q�і�1�/]��U��4�ݜ�g.�D�m��ݨ	>6�/��Rъ��x���p$�1^u��Y.]��II��d��&���M�"�sb}h Oo\��;�N^�\'����a��Z��~P0���/6>�皻2���v�uvIi��٫�'�v�G�}���`��A�v58(�:�W<;=ycs�p@zӹ�R�l6�<!.��:,x��K%8p�g�v��'�Vu����P�9�66�r�s �u�k�K�vpY0v.�X9J:���hS����f�Q �ٷ�S�G��$jŬ�\ѸB*J<�C��g	3��=�I)��b��=��gj�=�".��gw}N�ݕO_��D�Th�-��k�}�{�W�<<�wrC�_��ݢ�~z���e����w�Y8������C�f���I�ہ3��`C`�cL�%����&w蒞^��W��`�� =�D|N�=��>'+{'����?qy�#���#�3;%�GV�7u,
O���D�z��^�ˎ[Fq����lcq�k����l����98ϼ�3�Y��� �C̍�����7g��Kĭct#uf�j�5v�^k't]�w#�A�a��ŷ@D���/�| �muy�G[�@&�Lx�<U�J`��}<��H/���k��ۜ�|q�%�r�`�r��dl�3��;<6D_7M�X�~�d��`�](.�a����A��]j/kb��u�s:��$NK��vL�<%+p�;x���$Φ�}3���`�,�f$�_d������YںX̶D$]�Mv&���B�C�=��E�5
�suڇ���1��{��=��:�ѩ4e�[*rx1��������_�i��Er�jת��-��J���y��_uD�H�{����-�5�2gw�]3��݋��'�r#r�z�i4����G�;ݒ'����b���c<D���aK3��/P{6���c2)�tHj���紻srWD=vM���I��>r��H'p_�^�| �n��$�w>�����B�W������}0>ݹ2gK-t\�w������g��E��[��Ut��H}y��$�\@$��T{c_�d�,��X9)��Y;�3^�2'3�< �A���H7L�q�Ee�L�O�˷�Dϫi�vpK0t])�u�j���T��,�H0��I��n �f9�����̣td�����:�j��)-9NAg	�dͨ�H� &{ء�s�(�E�?����<Lƿ O�V�uȌᤉ��wőw���@>ޞzD�6ue5�M��wGZ��sc�Vu!g�*dzn�pA{6Xl�t��J�b���#�Sl��m�,��Q�r�N68F��E�gqV}���̯]G��v�Q��1ۯ=��1���*eƶ�*���ͺў��.�Q��ꬄ�и�cY���
�4�����9oZ6�棼󉋉�ض��ٶ��B��`;<�Ӽ�;V�\�b��{G.ۧ�o�e%M�2-�������ÛeN&��Ѣ�6�Ѻ�';l���Z�+��3u�n��g�{g�v��v���ݲx��H���H g|���3;�v������d��ۈ>$�n7�
�U�k��~����I=�p ���˗wb�A;��>3|�D3�K��;���I����H��� �|׽�C��2k���-{,��r�
�h� ��J-� �A�U�^$_\G��c��i�/8L3"�WtFKvVz���72rz}��-�`�$�._�x�}�ݓ�-�B��ނK�\_���;8%��N����@�ۙ�'O	��`��od���� .)�� ����7r����&Aq��Ħv	K"ۑ�sXLD"�s�v��fc�f�N0:��m����a�v�h����cz� �cd"9[�3��]��>q�[�.= ��l"<�;�d��3L�9���$�>�w�zt9r�<eC�@�Ҁ�.��~���=/d���$���ā�����Ӱ���g���,s{�&9&�t>�K������w� uW�W!:�$ds�k���$ݭ���ݻ��7���آ�N�ό޴���� ���)�x�J&�&9��9���2���E��C/<y�OK�һw�8|�MF	�"|I�rՏ��z���v� �i��0p��l��o\CM=�T��d�潃"Xw���$�fdω��Q
��u+;:f�����1��LM�e��f��z�ݺz�*�	�^=r�r�.��Ͽ�ƹ��iMO�_����'�s"A$��ި��WYձ.]��߈�E�\G�H �L�DΘN�Vk����w�#:���@�pz��j� {��@=N6B�fQu�!�v5�:�3���{2	'ǳi���v!��xf�1�Ș���2wB�.�kD��R�+	�uN@k�R��O	�D*����.���z�3)��a�|n"T�ĥW(eF9�Kz�/�;��fI�Χ��k%˻�)��y�g���!��i�t�,�B�� �gTH$�Χ�I3��n���םy2��ю����s�!�B�y��|� ��n��'=Sp�h�`ʪ��O����D��)�A�#C������o������$�GhfƯ<l^����V�K�3�<[���j��9_=Ym���ވMh��[FL�$�kz��=/��U��TUML�I���#_g�wrC;�����n�N�Q���ˈ�Y*�bI �o2�	^HUuG>5q�o�(���t�O��O�9��Ð���i�c��A��Kd ���Q�,��)���:�v��SA��|�A&N�3L��[�v��>U�gx�1/ ���~0I=�� /`��{n��[���z��hm����y�gV�͈R�:d�v�Ncx/-�^'v���h�U�݋�:w1i(����%[U(��Խ�I|ˀ ��Oe3�p�^N�W��4� �nd���93풢��;��D�ۓ ���r�:uvC[3$��cd˅R8:�^�o.�z��q/&������yS`�� 9����xN��x��I ��lyFofL��D7����4����;�^�X�i�XHDa�'��rBK;M�)���(#^���	 .�����&|I��1W�;��n���1���;�!��NT�9P��j�r=&[�W`�,cb��]�A5R�`�{{2d�[��n����f�3���4�K2QW�5��>'��^�d�=�Vt�gY������L�<[�sPH��ɋ�v�l�ْA'�e�]?4��<���ݝ� �{��Ft����뷷���o.���W��)���t��B�,��Q$�JLe<1��^�9���_hmٗp8�r�	�Pp��۴���U�j�u����_h���𼽑i�	�$R�G�S[>9������`J��A��)]����oJ׻���c��yT��3������}�hX}v��Ƶ���vﮦ�>t���\�C�p��g��x��S�v���h��<��tzB��oP���81
ES;|y֑�|�i��橺�V:`��Oxg��ub%�ݬN����6U��c�YHՕ]�f����1�{��v�7���>��[7x�n��N_N�e>���a%�4s��CP��!���,-��}�/O43��'��Zc��z�~���q�GF|sx�g�9U����Pm�H�ơ|PfbW��}}��v�;�~c'�:�>�ټ�ʠi��(��<���hX'���F��nS��C���kj�Q�M�q�4f�����Fg+'��p0\Z�{6A�-Ol����ø�P>�|r`���ڻ�g{�;���=��]�}�N��Z �Л:��,#��<�t�߽�FG����w����$���c��X��B��~�ך����y9K�P�NV�:+]==�W���_�o�z��ܯ����龈��v%���W�^�a�g��NW{�)����+��=�8cȽ�9L���hZ_������6#��~��@�j��r��k66sٷXx���ÒlG������guZ���fΠ|	$�A���5�b[se81�X���i�ۆֲ�Í�5��ݍ%g�bBX��ݳ�q��6��rI�R�"�!ͨ��Y-���E��͍m�������m����fDm�b��e����RY�P�m$�����fq�[l��9�6�A��-L��R�ْ;2�V��ۚm�ݤˎ���D�D�v�VY%�lp���V3Y��-�[e��ٖI6ݷm�%����8@�[,�3m,���I�f�6�6�mm�R��3�V�D㶬�lX�qA�IN(:q���̊H�����L�&g#�
�(	��p[v��[%$r[gg&Z�!�Q#��:E����9"K��h��3C��f�)g[jٻm�XڲtH���țdm�t���mn�3���cv�ݴ�l�ڍ$�v\��#�im�k)����+_{��������v����F�.�2��i��N���h�m���C���v�s�� �u$q���mnhn4��BZ�(�P���$"��\�8tA�-�0�C���d]q����N5���m�d8��8q���B�n��̄��.��-֌��I�saV���n�pkX�v�w�XM�v&஍2�nӎ���!�^���(2s.�����'۲SƧ��	f�mX�BX݉��Ś���	�����YM4W/[��Ŏձ��Įu����3=l!���`�e�����3�$��.6ғ����Ḛ����A�a4#c�����fQ�Yc�.F<��qu{^�L�Un�X�eͦC�N��q��R�e�,�XH���А���A�4L�w:9�ܸxz�,�D���%cisRo4X���%;Tq���;���2-�,��P³q�p�)+�y�N����K�a�O�	�=���X��]v6N�g�)��L���^uܛ�{W\�b�z����
K�)/;]r�b�� ^�E0����K�A����Ό�,)q��nwn�m����P�֬5������t,�ۮ�,�y��烎uUQ����s��n6钮�8q�ܴ���ql&���R���I�j$
����K2U�q�;\t糭���k�ꮞf �U4��b�ۭ혋�W'��@g�wT����/�vRLoRc��딼{8\���m�;����Bڎ�ZK�����[ZF���{lf<��i�A\�WO�R���f;E��]r�1\rt8���d�����4\ӵķ�	�봆d�	�s�j7]f�� ��T��ێ�����z��U�]bJ�p<2x֚��^�\� z��0]���q�D�Og�R�nu4��ɒY��M��=F��,D� 9�ڈ�LW��GgqǭZw#)��f�%���%�!+2��v']u��iგ]�6Pf�hGMmE�c���(�	����>	�~G���.䍂a��ʗe�u�z�9�x�F�8����djώ����i�s<k�nM.�kO5�j@�&p��{��v�G�$S�7]k���3�@hm�"���m0����˚rQ�+v#�o8�D�l�(���6�;0������a���L,�2�teVky�]�"��v�qB�玢0s�R9��7G�bo3�+�eJ3&��O|.؃5�eD�#�q[��M.[{V:8X�;kk+�2�Q����>6c���~�md�NgfD�H�$=���.s�'Z �4�J	�������e�����=�ۈ�H�:�z��$�Ƿ�$�s�`*ޥ��,�ia#E�b(�p�]�`�<�2[��VtDJAšw��u�
�3#�|H=�0#z:�:fr�fpS��)-5^xڅ�:Te�*��$I>�1�%t�o	���o�	��ɐHf�,�܄Hvp�4�1�N g�#�Ë�}_�v$�nL��iusA3��y��)ۉ@��3�$�tCi�06A�[q�!�/b0�ю�œa�6�������]b%ٝ���:d�wv\G��oKl���c.����A �d�vMF;�9@�2p�d��K��|��Gs�K$�T����=O�y���xM�1����Է��,c��?i<{ij�����׌�}��!�O�o{oA��= �M�W�������p*1ʙ���lq �k�b<H$J��O��Q�K���S��H�Wx�搇vP���|� �9<�H�:��p��:k� ��丏�[<��H�;rJ\3b<׫���٦�`�W`�ވI��5ͳ�Q���ͺ.�G>�c��	�||���:�&t�fpS�� �U����ld3W���Õ�S�/��A"�M�I���L��֥��؝�_���n�ocDu�6aw(]����9��f�8)x7W��t�f7>�˝�D�w(3G�H�Jq��}�&\箕�Q��x<d@$ҩ�G��n���,��3�
�?_t� �c���ٓ;�N�мI>�clkH$�^d	 �=[�_n��0}rv5ݙ�y��i�'r 93��ϐ$�z�unmO��f��#,��PfU婶���i�;�On�x�t�Ɠ��jfsm]�6=ý��L�zu��0��%����(\%�bY�$�ɶ�	��ٓ$���vs(;�(�� �>t��jބ�c��|��x�f�rdI;�*R���� �y��NN�: q��FR�$� ���k-�D.�h�u�L��熪1O�oa[Uq|TG�Y�ٜ&31H�޹�y�S���p��`��@w���\0�9��;�����Y���Jr�|l�dy���I$�GDM�����]:�$��ٓ>%�̵������ ��J��T�z��//NA$׻Wd��q"A��Џ,~\Hk�A"��&.��2�vg��I퍈>$��S�3^�y�Z��A3��"A'�:l��wfr�A�p�9c�Ƌ"����TMD���� �<��
�765�|f���O��;�[�ݨ�F?T}�4@�����-�,cD�Q{�EJ���h�]��k��;�p� Ѡ`�N_!�`��L�N̒7�b��;���z2  �������m��[���5�BD��	�S�y@Q��b�$�.�FS#�n[�ͫ[tzӼ�)���u
q��n�Y��f�%���؆�͑3�4I�������[W(s������2���gĂN�cǹ�qL��wtS��qG@bOe�~xg�ڞ���ȒAWF�|O��y@$��J�^������2���7�;�	�A���>'ǱMǃ��:�.�����>�$��؀A�S�<	��� �9I��;L��ݓL�Slެ��� A$D�M�� ��ܖ���̒5tA���3�
S�y�<�!�'��"I35O{
W����^�� $��Py H��ɐ@owWfuC�/��ڨ�'�����0w���;Rې�ե�GNx�yB8��Ò�e�ɢC�e�E�ql��!g����_Q���hzX��T�~;���Od����dq�JW��ύs��Z0kf�=�rǚ���':]Ƕl^*�ֳkb�&� 1�F;5��g��,�s�"�����(����v�'�G�����3m�JB;MI�&�P��d�>��H�����e�p4uc����"�1ï!�� �gs�V��7n�0��N֬,�8殍%f�i�u�>i���X0�p������dUN�9�W�U+v�\m[g�;W�mF8�8f�J������o���K:0�1��x$�)�I$�ܙ=��drZ�٠�1��<U��"�,�,�f.�0y�n��$�R�wU�f�|$���PI=��3�@� �}�]e:��_o[�^� �����v2R�P	��"A>$#�
A74п*�yA ��ٓ$��2���;��݊y��7@���̍p�u��$����ڢI��ɛ��r)�&9����{N�L��ٝ�@ǭ�M��y��vh�܀S�(�`H�j��r�2dI�:=1���2���??~���&�YmYu�Jl�l�]�z�f��e��Ge�ZD���>_�~�\+M6�<�5�1��vdIO�ܞ���ɡ�z��:�WvL�_4-��X��9��&��-���ue���ʡyT��*���<3Kރ|dX��3�>��S��l�wiė0���v��Wc)Q���r�����+�x�*�&|H'��G@�(�IL�e��F��a/0�!i7}r�`��1v!�̀�bfI$��A�����О�Մ���ܙ�w#����fgvb�ك@��T��r��	�F�D ��lx$��T����v7vT�>w�������ӻ�*����$��8�46e�iZH�o] H���eƸ��sԦiF������˕�xL-:�F���%-��V`ָf�Ŗ;�����TS%2vgn�[�t�Aݍ� �6��q�vhG�DEe�b��Q �h���S����H�N�O�a��&�+܊�	𫎈��U<�I��`���96LGu���m��b� ��H;1�l��y�$+��cX'�nF�����wfD��zy�g�?��#ρ���L���,��?�G�����O����M͝U�8�w�IO5�$[۾h}1O���y� ���A:�y��NII��b<I��<�oa��K���>$
Y8��NwmƋ�6�/%�����IOqސ$��w�2gvb�كH�O��e�ă����h��'��qĂD��h"3�r��u�5�р��.$ȦA�̋�J�jbj!Mȸ14�͝ n��c1�۪���_��U��ا�1�� ��&�ω��ۙ1��W�17)��Q��� �5l�A-�j܅��������`$�?�7�533�)��I 9ukG�3ݷ@-y��%�����.c�Qպ7Չ<����H$Q;#�`s9�M�� :rq��Goê��m��b� ��I�����=�+C���%�V4	��mȿW��:�����ګx3H�S��6��8!����!�ڷ�Z��ys�8���o�~��yW�gvG�U�� ��^�f��Ļ����ً�'u���w�bڶ�O���$�v��ewD̟VG9�3���b�ĆM�	ח2-�c�ET�m�ͨ!�=w4�2�X��K��bzf�:���h:��J;s�\C/=��� ����1�ɝ�y���7:���{/�$�쎈��չ��vM��i�=M�n�nd~~��wt�̙�'�*z �x)--��.Ș;%i-�!ω-���t$\t���5fvB��v�[�9��'b�9�D�{vb����m';�����I#+z�H#s�=>��^5�t���y��r;+SGW0�����$�MnL��Y��뙵��-��w��H򭌑!�B�w�`� ��w˂	9�O!͂NCg5�� �TU�� oLʧ�<o�>�UCHvX�Jx�2xk��í�N��,H�����n{�Vq�n�^辽��hq�wzoX���w�9s۾�ʾ[Q<�lȒߊ	g��M��L("tf����[)JMn���������/6A/C8�WW>�2�N��ù+u��P�c,�+Z�,W��m��;�<����H�ѻt�]a���ݛ��Ȗ2��]��q��T�v:g��v�������F��y���u���2ͷm��]�F+��-���ƶ{&�����"D�Bm����e
��nɱ��0�4Ŧ�MX;E(���x+�]��usZCj�P#��t��	�K���F�n̖h��5�?>})��,��L�$�ޘ�I<�y���VDTʁә��l�~��Fyyn��{�œ;��v2���8]@�OKLmuǨ�y��|O*�h�[R��U�}/���I��Ȣ	��Ҏ����������ﱴ7Tn�@7�1�㦛��'͂w����ػ̎zݝ����&x^��n���ӭ�˚f!�Ygy�O���>�5��:vEIü�:g"<�ă}�p^)�f\
��.Ɇ�#�b �H�i�$���r7ޛ�uЌ�WK&�^�ܑŮ\I��	�7iy������n�g�NY�C���7%��$>��V�����ow.d�O6���xe�@q �ƛPH꜔]�tX<�爲H�צ��I�i�/�7�2�t�5!��H�>�}�s�Ρ��u��%�N��/��05n�GI3a��'r�r�:K��錈$���j�$�}=�s>$���y3x&����g�8Y3�o3�����z�#�|��lĒH�X�]9"����cO( �N�fL��~����02gd���u�&躣n	 �)���̑$�Βv��lD�!<'�MУ��fAS�JM��ػ�2��f|O��fL�6��Ȯ����w3ڂA#+�&|	$Θ��맳�d�.��3��GrhM��OO��3�Y�v&3��W�+��n�߿����:vEIÿp1j�<�w;2'Ē	����g 핕ԏ^�P��&�rd�����t�2�.bODcǌ�\�m�fR��ğ��̑>$�� ŗ���a~�u��ݹĜ1tX<
�g��I����dm{���_�����=��o����z�^�qn�&F�/�,�齸μ\O�]y!�j�7�@����L�c}4v1����������	�q�%�����w�lW7�-wWmR7w���9ZX�W���<�P�
���
�z�E��Nb�4����㑁�C�/<|7�o�A�����=O�v���yp������=�>��.��_w�`�#���Yn�ܴwz<� �捘���&�f]��8�ldI�{XMt�c�w�A���^F��@2c���׼y�;�x����z�/�>~?y&5p� /4]�v�S�����}�늞G����������F]���61<�����Ӷ)alI�:iÝ�� <FIU�Q������
�c�"��d	�1�i�ժ0�d�zvQ�C�\wٵ�CĞV���4�����ϡCVj]��./^ϴ|����}���[�BcO�`�(�2�:E���/$^���<ޗ0���9&B@�[��zVٱ���b���19q��Y��և�v!�e��1_.rʗ*�`�&�����x�&,�\�a�Y��j<x�}nB�л7=X]�}����n���L��n����O?{��ڱ'��Û|J��YBH��,I���,ɡqsr,>W�Q3sދ4���Z��s�$���_m�OFK�j��t+�w��Z�������|�fv���[�T�j=�x�a�`���GpR_M�����}W��DݙX�!ZtA�L�	|ƙ�V�"�DY�n�����U���k���$#	DdRf��J��Is�l:t!�$�M��H8�%;kP䝶�Y��ݚ�m�q�bt��̹:"����sg	�N�����=��;;2�t�rK����9�6�8mi�r;-ж�-��ֵaÕ��R3p�f�q#�����C��;Y��jf��!�lf"�Ӊ�㜂#�Rm����[d���)�9e�0n��f��m��:
�ͫM�� �J�:&[�փ�Ð�Ҏ�P\�V��!'L�*[MٷZ@Rs��$�&bw"(�9'%�l[h��.њJ�K��8N
(㋜��,��$ wGB3'H�s3��eڇM��ֶȐ�q�i��I8 QΛv	Y�G"�: �'[bPI)vv�ڙ�;m8�l6���rp��)�
&+�5�;�j��̑���oT����'w,�;�i)��m�gJ�m���ASӐ$�F�L$N��P*ct7,��s ��y6]8L̙�'�U����WP��|��@T%?_L�O�n�@$���PZFl�������r���W���Ja��n-"�-Yfۙ�e���ҍ0���Ų��|�q�_�6Ϯm���v_H�I��~���zP�j7ٯT֨c����;�<�߲_B5j:4�̘����	���6�FG\d_����1 �k[�?�Ȁh,�|pk�y�!��5��%��As��b�į%��C4�Fv�|	�v �O(�>�Ĝ1tX<���Ni�{����A'��4�H'�;$�}�"��&����f��	�+��o�ߊ�����ꋽ�/=-�4oT[��"(���Y���v͹�y�7nu��L1����R�o�����N�X1vw`�g�l�{72$�v�ȇ��\�Č��L�Gsu(�{s�$g�38���~y�݉�ER̩��M�]��Ľ�H�j��2��&��K�7-�������q��b:���ۿ' @#��e@bO���2�~hܺ]|m���UƁ ��t�
��V��v!�N������"�.�u��ڜ���v�z$=v�Jv�d�%wn�/�U*N�4�����5t�:vE1EüW��uF@`NnvD�� ���U�'nz�����H��ɐHmӍn�	d�\���2�[#p7����$�^dH$��Ţ�q��YR4�C�T�*;�8��.g%'�b,N_TE9�-��Z�Ԯ�o�6�`Ev�L����ZT�t�nQ*B��r�6(�A����ǆ��=����}��ܹ�^�K��+Zf�2��k8bBw�Գo��p~ҧ�C�>���	��~�
�d۠w-��'^zt\��Nݬb���:$yᒤp8J8
���W�9��ݺ���6���(:�S�p'Z��Ѹ�P9�Xm�4
�m��^Q6+m��͡,�0cVʗi�iaҶMh�K�@n�jY1h���X7��]�W�p���yk�K	li�%)A�Q�A��o�(��*���[btۻs��
]�Y�P��2KWI��6�����|Ts�u�e�rH�Ҡ�4� =t�)/�����Z�Z��ǩ��kvw(3�wp�#Sl�I��"@ �k���,�Yczu��d��̙�?dYt�3�0v/2r:�	;�����H9�f�&d�	������`�2������a���v!�N��?_L�H$��<X5���YO
%�g���	����MoTz4El�N�&(�w�-��ɱ�An���e��D�̚�� �6�?��γ�̩�M��]p��7b@%��5��%��As�� A#1W(�(ƥ5��/��f|O�>5�N ޝz�%-���4���:lb-��I��gp�^1��j��tz�ɣ���jSb�
LZ�tWD�?~{������ɟH9}O$5����V�f�72v��e>NT��C9� ��o�3��A�3���)GG��3��]ȃ��F��2{����Ay���
�X��̻9=Y쒶��s,'ݢ�[��9�}郬�����`~�"�n;h�5;��ə��ب�	$
ͨ>�j�$�acu�Z�����$3�u9g�IfgL���A �*�#ƞxRO�euL�{��n�@>&u��x未Eb1.��.�ؚ�yo�L��9������j��F��Kqw�=�<q��$m0�:6L�3$;Ń�A�Ȑko)�f�6ۋ���GD@$.ڹ@'���d���l!S��/�)���0������P{T�PX�]M�������4dC�9w�V��t�rN A����⮀ğ7{&|j�/9�UF�W�_t@�B8��ڨğ���rQ`�ɺ"�"o�����^�A�j���}�>��h�|��3^ۦ��;;�;:p�#�2�P	��ȐG��.yw�Pα���������x?�%�2d�x?��S�������,�_�֧��c<���fZ�@t���{8|Ep�X�ЂGm�L���r�YܖLΝ<���MN���&�Z���}I3��	'���LH��0���
	��QH:!��L�u�$�UM�i��X����@�n���y��&���+��!8�|�R��Κ((��b�pȺt�\)��0W�Xj�[H]nQ��*P�ǒ�������H8w����� �_d	�$��DP�{�%92��]�ʀ	$Owd�-�w�s)8�1 �FDXLh��Sp��Tt5��Z��$�o��������ל�����R3��L�̍g����	5�rS��l�UUI�oV�( �&��d|�T#_kvwH�vt��P�P�w�E�F�j�6'Ă/��	�u���w]�n%�:_Yer�#��œ�ؼV�i����^��)����7�^�tB��!����Z��:ُZ`���L�VTJ����Hx�,�8d��ӟH�ٱ ��X�{9�6[�� �I��q �:��<N�����L4T�.[�MV.�B�6�fW1cie1]*D���m�#�d�Gh��� �z�7ĹtC�%�:�w>vL�'�f�G�@$εr�[��-1���}�*^�d���� �d�3$;̃�1�ymr�Tf����	$N�D$J��H4�T}}794�?���Kp��`�.#�K���F��9!�2�r[E��sJBk�쨀A��� ��Q�?���N���"���]MΨ����@$�*�>'��%^�)���v8$k��g��f.]�%ݝ0xGM�C�Aμ�q\��t�R��W�rfH"�U��so�$�%k�ۥqpJ�T��ڪ��^1�Y��h�ea�O9����~���(�ID���f�G��q��V�2韽68=]�o�v��ǣh�Mħp/wo��w%��w`9c���Pf�blK���s�F���(,���ѵf���려�׉�[\�����I��Yڙ��3d3Բ��bЄ�K�C1���Da�cex�{' GG2Lݪ^�G����u��۰�ޖ�N+r�;c���;ps��{k��ӫY�t�N�/��BJ���1���cXQ�#��&#jͭ�jZ�CbSU�]^Ѝ%��k\� E��.d6&0Li���R���Gmg�z{����3;[��6�}��ǐH4z��A�ȓs{P`�B������ �3��Mp��!؂�L�m�ψ/Ճl��F�e�= ����  ��d�3U�PlO]*�}6v��&b��yk��`9'ǲ�"|A0�Jp�GJ��rO��n��;��Bѕ����#�����Z�L�U���>'ƮZcȓ㹙� �NwT�����'3[](����N�}��3$�����3Q���[�O�@$wfd�$ǎw\�*����܌�T��;�&r\�����ݻy������㳖X�\ciYF*it��>~|~.�$��vO�=6G�&�s"I$wT���`�����F<	&�s$HjCgr]3:t�5�n	�7�U����@�B;�����d�oo�2��G��}��׽��e%��۝&�&Oڏa����ո�j��;���r}�����3�Dx���n�zP���ܖ������:E]�w�1�Ɖ��Prȇb8v��{2$��$�F�C�;��9��O��2d�M�SǶ�T�N�2,\;̃�0l���-��A1�3�I�;{Q�'������iHQD��%�mk�b�ˈ������IÕ��cN�Xn:�r� ��_j�d�Mv*!όx�+��Lo�YŪ���\�EKBɓ�&6��Nr��#��v;K�����D����kL� 9M�����,�N���&d�o�	����VWZ��ӵo9�'ě;"�ݝpIwd�;�S���k!��ńx�a�ˉ�$����	S���I��ƋwW��tDn�u+���3;:t&|y��A'���ǜ�@�A���Z�F�����dð�m�g����_,�5Օ�����`��i����D��B���F�nTM�͵A�XP_5�:|I ��DA2�y���(;$���;D�}���jk/l�ksc��ӗ�|p�� ��옎��5��0��&7q�Vi���:dX�w�0o" w�F��"L<�'�}��n����)�a��dɽ� 6����lgE�K7�,C;�%�}�1�T�����-x�ZgL�2�<�������O;�u���s�?��o�du���6d5�+���րOV\�E��Y�L�L���fI-B�s��i����1��uN�G��9��2H:"��[vܺ���nA���;�K�$]�A�U��O^�@��_6�zmT�m� �%!�׈@'{3&|HjCgr]���<�;V�_H�!���&�#������>$�Vd�5��@v^���f�D�5h÷�f��΍�k�Fi�T������>�w.x�o;t�vMpB7������[S��w�V��	�;"��I:!�ñ����Fv����P�t��ݏ�{س �Gu�L��;�!��$�;��TƸ���cӛ��F�����M��.�ڎ �p�+<����A.Y�N�dԘ�vf�.��n�"�� H$�f�Dx�J�`�%�mD3����̙�s9��gF\G��/ �F@�3�޶wODP ��5$����Ux�����ki�OW.����ϛ&|MvܗEˠY�fN�klE��	��� ���O���r��U��0Aۙ"I9�Q��|��;�K�$]�NE7%mS&zb;;.'ĂA>�����~;�S<ڗEc�DgWL�5<d0vw%ٙ����ف��I��S�4���%{�1�A$���@�I��/�?/��/�f#�� ����T_�����2���W���G�
`ʋ0���
,��0"̨�(,ʋ0"�,�+2��(�,�2�������,�0
̠�
,��2�̨�",2�̠�,ʋ2���(,�0�����2���(,ʋ2L�����2�+2�+2�+2�00��,��,��,�̤��0�0�03 L��̬�LL��̤�̤���̬�C+2�03 L��,�:Ǯ��Q�@�D	� �	�@�T	�@�D	�P�@I��X� !0��22(�0�9 �u���(��
2�̨�*,��2�̠��*.0"�`�̈�*,�2�̠�*,��2�̠���,�+2"�(�(,ʋ2�̨�,���(,ʋ2�p��0�̈�
,�2�̠����̈�*,�2���
,�+2��(����2���*,��0���*,�0
����Pu�5~���(�"��� ̟��f����ߟ����wd�?��,�?�����?�7����������1����y�5����� ���������'� ���v��
+���?�?��0G�O�/�O�k�!���(������(�����3������o���� g�����a_s" �� ��J "� I
,  ��� K"H�@ �

)
$��
0� �0
���"/8~a��_ޟ�҈� �ϴv��>�������A��|��_�%PW��������>��vps؟�I��'��|c�6��s�gڪ����?O��s����
+��������~;?�w����(���~��Ǎ����?��&���4<��3����t��o��O���A�¨
+~������?4?g���UEPz������������y�=��hA'��`x| AEt�~�#���PW���t_�)?%���N���8���`���}��|��UExMEL�䘁���>�p��v���u��(+�L]r�

��?������1�?�1AY&SY��^`Y�`P��3'� b��D
+�T��$S[L�IkE"��AZjR��
��AJ �H%%k����CYBUUQJ���ʨ��!
V�� wE(��٩Iv���jEB���`RI-"$R)3jkA*l�*E-0�YcLRQ")T����$�(��TQ-�                                              �o���<�9�\�]���T, Ud1YQS6�P�m*�0 �CMt�K���m��(m��/�  ��m
�Yj�G� �UL��h.,YU�yE����=RUw� �lQE�k�ܡE��x�� qh�b�lP>�JP�PU` �         0UY�{� ���P.�EPq�hv���p>ؒ����lq�QN�po3JQE� ��Ъl/�sB�<Ϣ:�$���^  �<ڥ^�q�d�p 6�Zs�:�O�Q�J+�U���� &TV���TX�*zj���T��� +f�  x         ��f��p��)VF�]��UTy� �+-Gf�9�u��ݵyuv�f�;{ۖm��J�۬smU��3UyD�2eO�  {ԯ��ٖ�nv:m�� �]���}u:���N��m�X*��w/e���� vU�nZ�����.�{�ԯYGl��l�����U��]3�>  �        w���u��s��}�v��N۷q�ԥS�w�yWVӛv��B��W��;*���y�� �J�n�{��meu�VގZEV�1�  ����)W�//rZ޵� ޣ�W,盡K�w���^w=��W��m=� �{=R�մ�s��knf�oe����Զ�i�M5%Ma�           ��գsu��͚�n;��^]ƪ�n���H��瞖��n��ѷ-Ʊ��͝[�m�u \�� ��P؊�K,=�*��(�  z��{�*kܺ�}� �)T�ݭ�k�����;����hvҧ #-H��wB�W3�K�Ы���D�IR�	� "��Ĕ�F�  �~	��T�L��"{R��F F��P�eR�  &�0�jR�P ���������p���@������r��O���q��	!I�	�o�`IL����H@�@IO���$@�BC����?�ns�|�?���=��|�q���v�B�7xnnSֈf��4A��Z$�,[��� �ͩYj=&Y�FRf�d�-S¢�ۨ���V�x!V�X.r��@X�Xf�7f̓���i�!$)�NO�B�蚷Q��/�Pd��A��`ӫ%��-N1Y�_!�����ӄ�Ժ嶇�(3���m���ӆC��w=)´<�NMP^�k4
�S0�W�+�
φ�݇&r䀂R}��b��n��U= ,�m�Rk8ef�a��y3x��\�WP5 �l��e�a4T�a���յ4
�\ݼɋG�hϖZ�v��!;��wj��%ݺ�X������gǦbT��(!�fD%���؆�-�,S�ɑ-������%��'�n�'n]��Lo!��M���i��LU'D��O5#���fs�"��f	�1�ڵ�c�̝�����(�iԱ3��*�n�V�?LN5�/�D���tf�;
������膝tlZ̈́�|Y�`����Ƙ	�e>�j�\��w����n7h�u&��v������W7:/�y��S:>f���쫙v�Ċ���*��X`�..�М=�u�wfU�A���s\���i�ǌ+yi<gI���R�3+�x�,L�I��S8 8���v2�XL��6&U3f3���ƣ�G1nE���gH�a�ǳJ��m\P�����R咇�>t�l�Um��^t��v8�!�Hn�Y�t� &MR,=�t�b`U1B���B]'��/uK+��B���n�w�'��wN�0b�o���K�y�ȝ�^WOU����%�U�4� �����'.�Ǳق�᎘ZrZ��ѳA�DL`@�~�'�)�aB��`�̒L��)I��Ί�v҂����u��mx:�&6Sav+�@�a�Y@����l�dc�4��\�]���FQԌݫ/dd��dD�ݔPSs,&6H6����f;;XQ���*�J��\������"�z�֕�f�suԎB0M�Z�Š9M���*��0�ꅬ�����q#��8���1�p�:㒰`�D-���wV*7M�*��h�UC��w���GlU�7B́�"���AD�aZت�����1M۹�u,�{k�'S\w��Sz		G�MvT҅�"�8,*khn�J�eY��YE�oĥ���V��a�_]QoK�8�:�����Ż*��ob��̸��I	{���J�� �w�S�$�S[�\��~uq$��X���^�����ǂ����Y�3�{M�^�o�����&L�%s��4��Gk�Ëh�b銭����惉uhIv��϶��tu�Y��l�N�c��@<�%��tN�`rh2�\2�K:��M�[*;�,]$���F��B���65��Gx,WlaI�`.��q� tY"�,�	kfƁj��ј!�)��p�B��{p�΂t�N#*���0:2�}"��H�L�'�X�e��8v���TFk��<qG��,��는uK�<�z�RHoZ�.�lWumR2R�7kQ��
�����$�F�V�ٍ}��،�y�͊zs�Һ���X�,��xry�[Qw��J��y.�pqQt���M,�X��6���:U	W��*�0���:ɩ2�`�Ė3LF ��	���+N70fI1І�����6�H�,B�gSz@h���ǋ)�k���c�+vO�
��G�d�G��]45L
����8�z�w%�1�*��c�K]�[L��Fɇ�t��ٺ%O5֚L��ce��ýr���'�S.��w`���c��L�u��Eh��R�K]<!����v<�{��٩Q< ̲�+"k��+�t�B�)�be�&7�8��m���{�,���t��s��-�4mR�$�`n�WJ��f�K�&5��xۏjn}_��(���C6��#z�s�	���,Wj�wO�ڳV�r�*�0���q��m�*�׎�t*���n)�x��2=tㄠ�U��7&�,W�)1�#g&wkX��p������wrc(�ý��WEP֐jc���,�30fM6p�В.�6�*#u�ӥ�*@���1���ʎkK��_I�4CÔ���@+'�	/�yR��^o1M��m������K+ ��U�g���KK��DzN�;fq�����J���ZJ��p��z�`0��qL6$N�a�y�r�ױ6�)���gM:�m���<Tt%d��¬��a�s&�0"ܡ�-0��@���NH�� ͊�*t걹�V��Q��à���U��Ks6f�2�"�Xc���6̵1]���ѓ+��@��eX��ԩ�����m��ʆH����,Mں�u #wV�v�o��ls �04o��
���X�D��ѩ��$$�9��kxȭ'%�{R-��e��b�ˑƾ�2�־�dR���2ͥ��/h~��/��8}�7B���(�O��@�C�!*u:�9;P}�R�}0�H�e{��67_rȳc��ծZspJ���0P��H.��EEOU�L��X���:L6u`T�UW�5Թ�K��V�J�m�mPɗ��72is�绗@�A�0-Bp&��3@��[�DT]��ҡ� �3.�Dc��}l����Z0	t�hŵ��d�Z�l���mǗ��N����Ҽv1�I�&9;��Lcҥ�7R�E�B��Pw���C#Y����H��E���*;go"�%03f�T��<Ks"��I7qb�yIK�o6��j�ؤ�EbI��XNJ�c;a@r�eQ��ə]�����F����ldTL!���2T��"S�tstl�h�d�׆|T���.g.JPsI8�G�+,ƨ���[o�BxR1 D���M�(ԫҫ����=q��B�D�Ӷ�؃x�.�(�&G`�S�:a�x��[C��L�� �mmkլ��b�i���˔dI����ؐU7����sd��<mK��{[��	�,Z�`	m��ޘ����F!���z dj�:�H����fW�l;]�� a\:��$�wd\S����͏��Mօ���X˺Y;�f��i�x^�-<�HQ�2hN:&W���P:vj|"(�VJGV^j��R�	EC�@+�~�Uҽ,��Uo5 ��5�e��)�e@-���Wv`n��
]�Q�fm��e�������>;������ؔ
��=�����g)�����)�&����{t^*'B�������$I`ʥ�l����Sɢ� �كj��8ؕ���ڕ%�V�ɀ��+"��f��Sv�v�3��KC�c7%F6Cs"�NeВ�V�1��ի6��1S5oq\MpK��p�EBl��pz�;#�dwN��6�
n�L6,�u���s��m�5cڱ�X��&�,
��P�,n("���r�ͨ�|j��e�㊢����s��uj���c��&�^R���N���])����;�d]�3��ُ��bѩr��Z����B�U
�m�[[j��f�;��`����a�N�#��U�A;�.�𵸭�]��%��}qYTGc��j;��P�VD��;�;xK�j�+;���!�c�&�9�,w�7ppY0�{�+${S*n�����X�:X�0�m剹���0�Rdz���,�˻���2[��٭�iS50�k�BY��M��0ԩ���Ee�җ��	�U�֦eYp5��T��4�H-��9=j/h�..GA�5ݩ�����k{[�-%�Y貪��%HPP�5'�l��]e�f|�ǰf�v?v����v��\�i�&Pr��`ڧx�� �P���4h��"*L��͜�E��j��vi�d#T�0�t-4q-Ƴ�L��.����}������A���+U�����WWj��b�b&:H�_EbY,�3.�7[Y��Lr��y����WJ�_8���sӅ�%[n�k�T��jF��s~,?�bۨ��Y�!n�r���t" �K��
�Å)�����Ė��\��oN�[�S1i�����f��K�+ܱ��T#�77Q��
,����khqa��J˧7����%0pZ�F�H�^��4��re@�7{$���VK�ʐ�{v*cǑ��&�o(�%�+f��V^b�t�|�.l��fV��(S�.��]��cH��ŕ�d^ n�>��݃�!�����1��e�e�V*�Tt�e���w���j()�0�6�h����`Uq���nI���[��׵7��bط ӵV�W��QV)�^�����V�·6N;Ό�y0XĤ{��7x���&<Ѭ��~i0A�؈�[�y�Fy����fRH��HI��D�T�6�XE-,��j�35�t��C1�X��-H�o�U��N&k�~�{kU맥��K5{�=-����Kj��������^Rhy��X���AQ-��)]��J���[�+����c8�4�M��e7(�e�,�ڥ�je���(�JrU�l�H��߂�rE��s.١/h�iܡtscڦ[��5�,��!4�tB6��AtUl�c��Ʃ���T�`�$Z3n�7tv֐v@<E}  �H��dy�tH�i�
�3EE83Vk�I��@:�N:k*���N�Ų���N��B�w!u�*dm����ե,W�S��.�B=���ǓԼJ4��K��.�L���5�Utu\Ʌ1b����f��Z	�(j����mf��Dޒ�1�^�i�ى���C١��,�:�)���i�U�X����$0m��1��N0����K���(�S�tE6k>.-e���X�va�%-�e�d5{4+�N���3�&��Go�v(V��Y�KV�:j��fe���`<0]���%�b�m
t���2��yQ�o���S0<YT��*H��`3n�OTF�i�%��ͼ|�*ƅW{���Dk�}�y��B�)0~��{䜲vX�/U�~´e�fŉ��jn�-;Jzϳa��J�e�NR;q]&i���z*&�8��&�m)�w��ƒ�E�5�4w�k���F-�l�7n��P�{"�.�,Wg7.�$��յ4��AR1h]m��f�j�Kʗ`�+_ڨ��`�5����@�U,���^�����ǳ/BB��vr�iҭ8�j�ۆEA���F���rW�c�vB���p�o7��$2G�i����:�;�hx.%�#� n�4/�[�ZC� �)e�LՕ�	�����n��z&
G!�y�4��w�TN�����;�b��q^Yy5*��)��{0
�УMk�3	Ob �����8N�]'-��A�R��ih�,�Z�X��7k��3��I�Z9�h�����~�����`ۭ5vidpe����]���Ya�1��Nk$��bc+p��L�7�Y1�
��!ɗ��N�K#�e༹��E#�;R�I	�bIt�d0��ސ�2�GI	Y4KS�^9��%$&��v����P  �͕Vbp[�;�3Df���8X��WW�*jgHg\�1X�<��Cш�r4�Q.h,���R �;�J��PɈU�?Z�mm8�e�h��"5�y�Z;*\7T�g�Lejx�lB��i-��l&6�f-�kV�Ye��8��v�A	���1�2:w&,f���Ħ�`V����۔Gw��D@[�eyF�CfH�򯫹 �e���2�W��Lr·	�+сt���=#�R��*�t���|��F���ķKw@�ҩ0ȏ�9��N(z6�:�ۻ����U����n�Ydy��{f�����B�*����G�;���l}��8��3T+R�&-�MU��ٵ{Slx��Q;����[>��wQ(�r�J�븙��3/W�;�E��V�!�0m�(Vk�[X`�H����GMn�	���`6a�����@V^)��c���Z�è-ۛ��i��v#���8o6�mD���݊�Ζ�VI��.��S���v�i&ij���D˳4�4ځa��EgBU����5�M�7;��ٸ�Y���݂�:m����ӫCa]\4�sF�e��ʵMi9B�	���6�VQ�[�hAOY&]�I@�z*\�w�� ZZ�y�.ww ��j�A@�����ޫö�tی-�q�o`[j��#YTQ�9(l�7j�f��γ5�YF�/��5�&��Pmؔ�Zhr�kl����Q��l��)"�(BB=����Z���v�Q5U��{;V�������j��nl�J&�՗ �&��[�c�" 0�k6����(�T)_I�(M9���퇉qD�2x`��Q�y�2
���8��O���daM���v4�m]aZ��JmJ�3tۣZ�^��XjE왚a3 �ܶ喬�[�[�CLm"ɬ�����`I� �y�&c�v��S{d�����9� /ۻ�ݸ�f��Y�&n�?mO#�x���<6����;��oSI�mxz�M�\�8X˪����1
��u)t0Ф�[l���w���D�Y8�K�h�Ω����KŃ��U#���;,�&�5N�6��ʮ��S�b��ʌ(��6�I���Cc�JLx]3yC{���Fs�X�;�ׄ���E맔�p��WaCZ���:���*��p�Y��[�"pe���$�Z6i�Tc(�V��W��8a�v�����A��37���@����� �HdaHB(@� 
B �P� @R
B
BE	%`IP�B��
��VI$�H�,$�Y AH+%@!�IR� *H�E�H@�BHI 
��� ��P���	 Y	+�P�"�!	H��,�XBAd$��@�� E �I$��I$�H�!X�Q�J�IRB
P$$X��B$P�����$���������"��@�I! �a!+ E�P��AB@P��H
 �T����P!P$���
����d��$%d��HJ� ���R�d��� B!!��$ I9�����?�̾c?�y�7�p/yn���&R>Ō�y{Mՠs}�a[û��@�.yJ-����kyb�Q^�tD�76"B*�;��Dp�!X-j�Yi�C�0�~s8҆��j��޼�-���#��~۫�D���^��]�<|x<u"W��9�px۬�ܰ+*L�2�V(���C7bz����<����y���+)�w�tP�@k�,Ɔ�oIL��u��{+P�5�R C3�#�V�fj�ּ���A�ԅ����PBz���a=�A�$n"��՞�c�k͹���m�i���C���Y��$��p��7[��(�]�����/z���Z���zL�7o��}��V5���[W��00�ސ��c�dx#3�I^���X|�):�g,�0 �j��+��(Rǯ-�on�N�L�tFlwT�XKE|��|��N�={��B��7����Z)�E��H�ҧh^X�B|a�tgS���v�dl:���˔WZyj�*�}�/r��Bk'�5�!kߦ���ƈh-�uZ��T��M��V�:��K$�Z��2�z���=l�@e����![�e�Ĝ ���"��Ź�C�qśBoEd�c	�DGMN��o7��La���єw�}��t@9v�"����R:�n{�
;�Sǐeŋp�Lu�uX�B<�T�����մD_�����j7�;c�yY��GhK���u�LDJĂ�}��E|:֟�t@|qbZ�O���"�7�=-��Z�
�Z������Cf�q�'`�7���<�c���EM��*̽��5�-�=4q^M�Gb�m��6�e�e,��SN�
�1��S�Y�Ɓ�����s|�����';�˫̃;{g���y�ڜ8�r�u1_m�ݚ~}���!���M]s�5���~�ݯ`e��k׷C0B/��uf��/sn���U3f�%W�#~�O�[�N�1ooB�7�fV��v���k�����-���Y�@�z�z��ε�G����N�u���6 ZT��5�JJ���罃%m��=�;:�n^5�Lv�R�ڞ;�f�aIt�3�fʲ�I�(1�U�mU���g"ru�9�>v��wwD����'�{��'�Ն{���+_{�F�� k'$���h�q M5���PH2-U���<�y�QXc7^V��Zp���i�H��|�	���`��;FV?)��xl��p+��n�d.ˆk1y��E��D���-H5���;�%J�:�cܭ�����������٘9�ձ��ZԦ�WxQ���H-���UI_h����xշ�潽g��ݥi��DB
�61���~R�26����6�++F\2g|:�f��4�$�����N/@a��ط�Z.��&�q	����0�Պ�#جu� ��������å�]�
���~�d�(�LFb]���拺V���� �$ܻݺ�r#�f��
�Ž�
l�M�(CG���u�B��;�
�9�.ѻ��[z6M�}�d��k����}Yʣ�ݲ���pU�V����s�)SӔ!��@�������r�y��f�K���!�˨�x��Š9��K�$��o�7W2����^�},���o4"�`y�0c�1l��Lk�>G�Ө���A���H]|��[-Q�"��w'(q���"��]��z����=�T�ڃǛ�9�����[���%�=*��6綉|�z߯���sh�y�}4��݉Ye�Sɰ�#����:�����
�
ŻK�oer� �4�Ν_��=!ڬ�����;!s`��y=���J�m�Ⴈ�"�6���}�يD|ӳU�X�yT�����.���ҳ;A�VjX��J;���K!�N-eL��{�4��c�
�r�6�3���m�i�fWM�G!	��-��VK�e��eVT׆V�������<�6�z�ŀJ{����X���ǋy��վ�C_vM�X|�o�}�-#��wo<����2�Ucp��.+{p�\�!��ʼs�.Dlb7|qVq��⳺�ze�F��(b�Y���������^��jSF�ҢK<Nk�y%�@�<%��~c�G�\�O�I�΅����ik��G('�v��pp���#���"���J�]���uI}:�������m��,:$0��E]K�o�*��_�{i�(~:�`G⃹�w���{�����W5����E�z��lYϬ��e�eIH��� �@�m���H%b�����c���u:Ri�Ȧ��9L�Nz�F���xk��WǄܳ�}&j��^�x�Y'�a�@ӻD�ܯ%⛴p�d%!U;;�uȫ,=�� ��û%c.(2גv`�����Mq�W�Y���K���C9��MV�Q���gV���O�Q�w�6���0I˛��ܧ�)�t���9���>���G�x�/*fR���b1�S�/n�q��ħY�{Vv��c����|��"܊1'J�(����J�V����;���H������<|���E����ʫ���p��!~v�����;d�7
��yg���yn;V4�~|�O{�Eo�V�eZ�ۉ+s��obw.B!�z�Z��u@�� �k-W6���Ug3F $V@
��s���8�q�C�7�3��yhv��o����y���׸�,���{��]�ؔ�,k�nf�C���y$��_\ܼN�����;5c��D�f�+K;��K�\���Fq���8���g1j���z,�Su�a�֡Oݶ��A�ї}��Uv�����F}���mo�;ATD��b$��t����+6n�Je6a��<�@Ӵm/�5ZE<�u��)깝�.���^^�HJ�0>|����6Yٝ��3�h���O*��ëKu�ⴥ����l�pL��޾�&�����U��k�ѭ�A|�Q�1�GމŌx�}N�tA9L��g����(KF����	�NbJ�:�5��7�1�7v�CY����.�|�Sz.I��FJ.^`8���d�!��A�S0Xzj��y�C�ӕ9eM-X�R�����crld� \tx8��k���7��Z�*E��Q��U��W>}I�Ro�0��+x[-�]J%�x!��l��hȚ������ȇE��L��{����^�7���;Ӡ�b�q�R)z�K{�\��ɈV�Za�ͤ�h����%v+Fw)�C&X�/�ܩw˷�����J�"���\��CG��o��3�7��L\��˯.�t&o��_vr�1D�3�%�N�8X-镸��-Qd��Jҹ�V���[G�!2[��N�6]둏x���~�l�I��F�!��+���&���f'2����.��n��r:�HBev���X�^�/y����$����)��C}2����g�_I}���h���T{����y`R�Ǟ�~�SC��R��X%X���	�\�W�꼽��٭.��̮�{êP�L��qV ���3[8j�N��7hvn��L��ǉ�� ��+�-;����r�,-�nDdˮE��{WkK���7s����s���ο������j����~,������]�A���UPd���b����t�`��\>�˖�gq�;MY�R�Ѭ�.�n콱Ukd�R��]5'i�k��9���u��;Ķ��|��"���"IԳrIA�7��ɱXv;���`X�]���ՙF�B��h�4��\�G�K<��v�"J�#�Q��6M/�ֶ{�TP�.�}�Wa����������6��$#F�'4*̻��eĉr�5G�<׼�*
������#��
�f�ˬ��ZQ��,¢w��u������zp���|�cgNk(pӡh%�(��M��]Y�9��jæ���;��h�&Zt�Z�&�wX,�a	���5D<�<�S�J��S����w�j tp���w�9%X�隩 �oWv�SS��}���G�	 ��3�/{������@{��H�Pe�w�e�Mel�lt��NM�'�.��r+^`Z=$�K�*L.�Vx���7��3���&|+%ʗW��Y)��,-Wd
��&�6�d�t2t�5Ja��#wA����ݓشZ�j���zjsZ����{�ރIvi~��{V���ٯy��rw=���0/�^��L�Ƿ��E⹁��|����ۃ��k�;��@h�$����4.t�un�}��U7�I�K���gy�{۱4}v㌟Mɰ[�^dZf� �z�û�.�7��
��q���(uum:��ca=�5CHZ��&�Wx�8��u�ڨE�E�\V�׍�:����)מ�����_C�w��:#�2ʦ2ބM��ɍ�%�y��H�l%u��Sp�:��EcHh:�X!��7�NS~�_y�/r^
l`�j���7D�F�<X��Ѭ���� �9��Ow��JLVT�f���ʭ��E��=����A�8�C�����d�q��M�ާ$�~�?��7���Y&���e��!���ԗl����!Uk�<�/%��ͷ��ݩ�.;P�Rq�6_�+U�}B[���Z^��PN��%n)�O<�`)`a���G�z=ϣ}��WO���mq�|͝� �38��۽-ç��TIݹ'R��F�U��^̑�^�����5ʐ���Q��ڦ�8蔅�g��W{|��͡NM��$$�ZYL����]�����5�*������8�Ҿ�����![)��K6K$��J�k3ok����r�b A��z¸���-��K�SjS�����r��#�7�ΥX�����u��H�$�~�BV�;�[��B�غr�Z�+׌4:&ʵ(��"л���J�((��#�{LvT��|�5�ŕw��8�n�ͧ�5]o`�n������5�I���Ǻ������³�W�:ӹݾy�Z�R�W4��i��;t(���e�\Y&�k��7�v�ʣi��0�ㇶc��.��ծ�t2�{5ԨR2��L�.o����KE_�ZǸx�c�gg�_}�ZHeӺ��A�Ƿ����}_��>0Л��e$��0�Ԇ�tpL�B�)�N�U]P���b�eK�u:p��V�|��������#nb�}��[��Ok
w<}�qWq��Ղ1������=
��g�V�/�1���=\%G�z�w��WU��@n�x�f\�W��!������7�����Jy�����F�fw�2���� ��O�;s��\�)JZ�7���+FI���D:�6�ۻ��QZ\���qi��Π󯸹/S;��1k�ƞ�����%K塝ѸP�vյ�WV�t��[ڪR=(vK�Qi�(�ŮF�q��\��F]w
��dǰvZS��*-+:�)�t��1�(1Cܾ�"��:,͐n��U|�eV �1nm�»�(����P��ےZ��X�M��9�wYE	u�h�a6�Y����Q[�d{����n�/ �r���Yq%�Ӳ/!#Y;��/>Tc-U���eG�1���Y�^�К0x.z@�?w�$W3�+o��
�g��Gq�(r!��ul�ϥ�x�`��kĜ-��%�[-d2n?7'w�`��"�~�z��Lf���SM�,cq������d`�^;�2�1\�H���P�-�z�见�mӵ&܏rS�wu�Z�uRJ�Ru��֓�wTN)+P0{-M��i�oS�W�\hd�!��~܄����J0v�v�Ү�{%��׻�]�u,�#��9�J�ǫ�����O��&��ɉ��=�ޏAF-�\9���-s���kĻ�!w|�u��˂ �t��F�X���`��3��3:egk'�By�:̚Di��,W�n�M�f[9��U�S��t&7.la�n{W���}Idz�����hf+��s�\xKP�õ��n�4	E���fέ�)뫺�u빒���,��0L�*v�V�j�B���w{w-��n-�7o`� �IS-l�����,z:����<%D���6F!�wx�G@[c>B�X_Q{XӒ�NgXw�/.q�w��/ R��P��o0��,gq8ks9�76�[�5^��w5�-�x�U�kga4Y2��׊�N�}�sڱ��ݙ;z�y�J�3Zx̾w�o��Hf��s4,&f��+Zͭq�R��W��4��+��Z�li��gk�ۤ�b3�G5#n(�(F	���{%��T6��gy��j�`/}CFg� �V�<�������@�,U�P�uV�r�e��@|�yY�g3D�D�mq��ޚr�y �7�0�]r+%ޜ��
�E�x���,P�a�<{/a�QE�_F���͜�#���|�6դ>�:U��ߦ-��~�/�sT|NԬ߅
���N�&�����On�r�����[GJ ����`�oVV;�.��130�����"]���Xч��.�&-�Vsz�#e�=��#l��2*�]*�v��EgV|x����r�2K�������Xq�o��c]z�������`��;rwL%VrRok��MB�;�-���Jueҧϻ}��:Y%�O�{{$;�;s����t�d�aXݍod.����ɴ�"�\Ӈ��gx��O/i3��T���<2Nb"2��ʵ�>�l�
�._ �s����Wu-���V��ok��(��[���ё�^��9e�K�&��Q�+�g�٣��?��{wԅ��N����Hl��qm��n�ٲ�]�Nɻ�V6�/kC�"��`Z8~Uw`�
�I��D�=f�v)���e��ߎ�Q#Wi�3F�6��H�9��1	�wtU�U;�e�q�'�e�B �Y�]ے��9*2L�Ҙ:���{R����%���t�hǵ"�����׼�8��n�>y��$ I>$�gy��
ګ�������f�am���u�6��i۫oL�ы�{s��,pC�)Nz^�x�V��W�ۚ7 �.��c�y9}�͹2����	>I��;�m���M��Ѩ�����kl�Ŏg��E�Fۚ��c[n�$y�pk���۫�\<�X�D�y�v��G�<�=\vJMn��s�������q�]s��v���-ə)�l<Y��u�Ge\����1�g��[�h�"Q�;V�iZC��Nq�zʓ��ƻ,���4���7tnn�Y�M�.C�g��F�it��=;k<w1��GlXF�W/��5pj�u���z{���3�^y�ͼm���e�[ӗ�[.��mi0y���m��*#�/i��v��<a�g:�u�\��^d�H�M��m��h�M�.3A-F7�6������N7n$v�����;����t�l�e�Gcu=ls��ҥJmEpq�|d�8�u�͸�f�)����ͮ^Ե��	��ۉ��n��0m�c�8��[+��(�͗��{����no>Uvv�u\�n9�f�A2��[VBk�-��]/moQN-�7#��٨�:��N��m��\���9�/jp��� 5�v��:��b��+ϝҼ4�ձ���f۶z4kw;h{q�;����h����'��f�ɞ�δ �lv|����P�ۺ�ݶ�ݵ��\p[>}��mܼ�)k8ɽ�`�K;��On�)���������<�p�ю�xz��f���kB��i�ӯ9�TSp�,'���B�;����un��h��Gm�I�|�nx;q���Gq=G�u�r�^<�z���gs�M����V���6���{`�a*�hD�6��l@F��pq=qܖ�eP����\��Q� W��>��q���b烜s�Λ;c��c��l����p�n:�vf���v��m!�X:��2�s�+�3��۝��մ9S�K\7ۮݝ����G��\C�O�d:�s;i9�#������N��[��g!��xʬ��s�Hۧv�I;9˰�m�a�z�۩�PN��6:���N{jހl+u�x��6�^..��vd���5�\�Ov���m��p(����ϣ�����[�^���m��b�`����a�g�ΰl�i.�p� ���v�nuѥ-{����6Cst���,n�\\k�#�������s�'0a�8zt��&GY���݂��u�*]�npnj^x����-ۙ��h�5���o=w9�X��s�l��v,�3m��	������+��^������wm[^&[W{�n�s4�x��q�jNxx���lМqxݶxǇh��^cV爹����v����p�e�9�sn|'<�{\�d]l"���(!x��㝹`kn�u͹�)���z���;��GjCntn��hy�v�-�Wj�!���)�X�b�v�,]v����uٻ&L1Ѻ�"늂d�ٵ��������G'�����w[�՚:N��[�G<8�t�ո��ݮ���V�2`;v,��ۮp��k�B�-���kێ=��� �Y)��g�:�ۭ�W2 �;k8�o/gw7OI�w������n9:���!ֹ�Ƽ]��v�0�+��9��p������[x�n����ì�&7n��n�٬�V�;��d�E8rX.���F�;tU��f��ݮ����-�1���q=gm��tm��g�퉇����������GWsG �nx�"=�ͭ �>X�9sێ�@�1ph���F�k'4�s0�bLf=����͎+nܣ[s��ț��g�N֞P���cv��[%��m`��9��.�������s�6��pI̓ip�E7m۷IX܆8��%u�����9�zƭ����w5Z\�7U�����@>��l:���݅cFA)�,i����[!��Iݰ�����B�P�=K�֝�Xl6Ǒ�5��y�,�$/�`k']+��j5���І�k���tt��;�ܽƮG�:�����ީ:�ݮ�EPخ.0�2X���m&=�]/`�j.�u���c�n�G7 �v8��2��8�瑴�vo{q�w:�x�i�c��^� Blp+���8��N�R����㍧JL�n�F#��%.�.79�v�����9Y�nώ�r�حv�k��l�����l�H�8��;;Xn������qƯ/k���z	7s⻒��grh�o)�glk�v+cC�'<t+!�s8�SoK�]t��ɼ�+u���3y�����f:s�C�ɣP��ʂ��c��̏�箳�HN��뚌u�L=��rNt3����q���b�s�6:Q���(�n�U�+z���t;Ywn��G3�ok��e3���kk^.�w�m7v����gɘ�s����맳��xnծ�����Ä�ݺy�rV�RRN�YSZ�2��`�.������+��FtW��6y��ͷO�v��x� �y��.:�FmQCl3���;\n�/��H�C�\��s�3ǌ[��:����\�q�W]kb��S]����F���Z�ù�ƻxޭ�Ø{��Q�9��lœ>y���n:�r�6�ɸ�����K�n������k��mg�m^NS�]��Gk� ��tuч���=tݹ�vⱹݤ���ۉ��=rty�<WI؞^!#r�\r��N�n�6zN�a-�۞)M�v���/Fֽ5r�s;j:2���>yu��@<.��c=�7N�R�7K��ٻ�������ڮ{<�z�^����v��ۛ���=�d�h�,Cv���{qlN܂��^ݱ���`7<����x�����h
�!��ػm�].:�Z�����(�M
���\�:��͛:XMה�]��d%���pXun ��k;.���[n}�U��[q�7v8��npu�99�q�m�'�&V����g��>�����\g�����q���]��\A���p���{nպt�v�C�m��ٰp��q��a\��!�ն�c��wR���U��u�9� gq�]���N�Q��K��{s�v+���u��.px焙����[�v���zP�:�6��"��nttN{[U��u[�cD7+Z�����rv9���α����fk��.�{�B��j�;�N!ٍou�	v��V����C���s�3��Uz̹��`��yw)��g�cZ-s�<q�aK��n9P]���= /;��];t��N;qÔK���G%�:�<�۫���Kl���)�y74�<�i�l��J0[v��,��x���8��} B��q��i��v�6��ڳ�ʏ��i!�g1r�����VF��y23�8�sc���v�pSَ����`|��2�$4s�wl`6���s���V�v�u�v�A�m����O:y�ݘ�z�n{I�l�u�kq��q����ϯ۱B�1\��n�dM�ì�p*�3�"��K����}��r�=�����G��y��@3�r�8B��6�����z���f�gr���|/Q�FLv�g�7�v
\Q����!7&���(k��R:�k��v�����`G��˥�Eroƛk�+�e���KͶ.}��={E�u�q㵋Xݼ�b�û1���f���ݷ��&��6�&��8ص�œ��]ۃ���ώwg��,	h�:t��6ㇵ���̗(�{v�2v���;9��#���Ëe��`��Hn@��ZΨe�[��nL.;��=�����)����'u����h��\��8��P=�x��rV�s�z#9��ɗ{��Z��>9	�qq���'^��c\r[ku�ø�ݤ3��,ҽ�t��K��/V�l;�x\��M�Ny�M����{��!�R�4=��"�ɛ��7�^������b���;��I�)�.N�u��֙�1�2���Stv���0x�k�sg��qq�m�m�x���u��f�O��S�܏���P8��n�E�@��p��=�1��hv��޷E���S����^���<���v��|(GD�G@׺,s��'e�s���/NK&�[<h�Ccw�ɹt'<��ZyV�3�C�=I�3g�u��^�q�^l�Y���F��Sׂg`���c#C����7.�̛s^^դ�0^÷=�MAE��6��J9D��y��;`��0qV���� q�d��n}P���n���u�Z�P#j�k�#O^rf��X�������3��ln��bvݵ��!���n�����]e��uv�z5��փ���zU�D!��ޞWR� Jbxv���=��c���%�=Iڶ��<U�u��l���%��-�D�b��[�w����;uݬ[��`��=��������>�>��WY�v�c�"ơⁱ���f����n��h��ݮ�$��g>��[���p]\u��h���q�ᷭ����vM���\9��4�k�����<eyۜ��2��&��r\�x������7g��V�B�5��7��V��0�<��<�Z�v��7�46u��,�u�K��ۗH�v{�^�2���z��O��[�@	4�n��������rCR��������8�I������<�ƣ�������(��n�nҽvӣ��;&2�o��]��d6kXm�=���6���x⽊��|�qR�f��nDs��qvs�t��e��{2����ź�ج�۷Vy�p�,iy�ތs�{.q����:�Ÿ���lv.�e��p��=��Z5�v8�q�Q�m�r܇l����8t���n�tZGv=��;g�]ɫ�w�e����ΗTҊ�Ό*]L�w;���w�b�s�N1²;x1t��Vڛ�qx�,n����t;�n�ڹ���km��������q���;������2��;�ֱ�p�[5�I۲����;e�3 ��Q��Ş�z7j�;S[����ܾ5EF"	m���DU�""�m��Y[�-��Q(*�DcX#XQ����(ł�Ym����m���E�b�� ��-X�Q�0U��
+meƥU�ciV��)J�h�TAUb�E��Q�dQ�mU*�0X���HԱTX(1`���Rƥ����Eb��Ab�EDQPX(*�Ғ�1#"%@��J�DA�T`� ���H��������FE�,`��Db���#����������EB���X�AR�"��X���#*�����E��
-h([b���m�Db�X����AA���Uaim��mb*�*ԬX([QEb��U���
�Q`�U��Q-����1F(����b����TD@UU�)"+U�UbŊ�
E��I&s����nǤ����j�7�Lq;ն�nL݃��Rv��Cg��vNX7��ܹ�b�ی��:���7���8\g��cum��t��n��O���r�G.3����a�Fy�:E���'9�NE��"9���:���/�wh�έ��<��<���Iϱ�41�;qg`��͵)�Z~>�����vpp��k<v疹��n��Wr��q�p�\�i1��ܥ���tVq�:Ô�wk'r�K������=��L��c��"W`�x3�p�v�>��b��yn^U瀘����v���5�=�S^���ɭ��ey�m�bhI����q�<f��F���&�N�(2�b��m�uײ��Z�m�KϢ4{v��\�<�8_O;�c�ј�hݮ{/�[��݄[u�֋��\sg�p[�����tr�n�pc�['e�k6?�|�\C��[����ں�z�I��J�>�M�M���r�}�rs)��>{r&�7��ݰ���wlV�vI�۽�\hr�^M�7�u�>m�=�2%��デG=C�=��rT�=�$��R�uѷd8�29ْ����Z5v�7�:-����؂G�6L�v���6@�؋�y��;��XѶ�;	���.|Z�\�VA�W(��5��8M��d�>����%{�����p�nj�����:�;B���-]��ӏtz헨�,��{cr��۱�$ű���M�F���Ŭk��8�ý��o������L�;�������@����G>���zs�:�.�6��I�G�����t:z7VBܓu���n�:�`9v.���,�ӵ��'-�;g��Ok>4[�gY���9���p�ol�q�눶�Y�6�dr��ͺ��;��:�\���ݭ��`�n���ٷ-�㮼���kK���ĸ�a�Ѫ�Z�i�q���7\���;��u������z�j{;�%�ۗ�/&�ږmۗv��m�����n;^�����L�6���q��9D��{u���;������=�;�&w����۷g)��1�7=��ɑy^ˍ�p�<�r<�{q�{`2"��|�T󇓅۲���>0`ݷ<�� r�ۗ�'+���ݹ�yyqɀ;m�헓��n�;<8�c�q�=��<gl{{>��W�x���c���?����|caB\/���ʺ����w6���AM������5�!�{ow���N�j�E�'X>�!
@]|�wHW��6fC~c���mx�o���[��?��ƫ�YK��Ϫwi?��``��A�����Ҡ��F�����qU؋k�^��A>ݮ�$�^��	���$,��)�G�{o��$��&�$�ޫ$H]�ƾ#�^Uܮ�q&2�� ����ŭ���1�	�@ɻ�>�	�׶,�ڭp���n�ޫ��Ϩ @:��}s�F��u��{���@��n<�X}gI���{c;]w*�҇k9Xy���Co߿��-
&c��$�~�$J�=�� �9�K���� -�_(�T���W�"�~�&Jj%���&�s��\ �Y�Ѻ[����,��q��]	bT��)[S�ĥ���J�r���mP���-ɤ	���h���{kx�eޔIpN����� c� _�H
�~��D��y���=��F2}b2T��7�� �$�{V	5�g�n��Az\ݾ���ԁ��;���9���M0�Gw����3:����;�?�yH�O��yvH${z�ϭ��4���ARޚ��ͅ��)�G*��d����Ԟ;bS���'��{w� �����;5�;�6z���4�#P"�a?]v�,�ݔ9v��i��	;�i���;r܋ֶ����lj1Ċ�@ɮ��ǆ� �Kۿ�����>��A�d�P�v���ՙ/��&��a,
&c��$������{��� zb�J�}��@P����o����h5��B��/��7z���I</����)`��!�N�p���Y[U<�sw*�9�$	���f���煼�vLe�dÓO\������F� z)_��ج�b�� آT	#�����BcЈ#%H���bh$���O�2wU�I+�y瓦�.��Ev�ؾ��``��%���|�� ��N�}�m*�iU  ���d����d�̸x#��i"�5�L�ى�77-�q&ѧqWc���jN�X��'sO.`Ơd��p�>�����'w� T[�4{�����%*�y�vO˯��P(7f�l�H\����5#� (
~�y*  [�l�.�{{5Nu�ᴱ+e-
&c�0���n��|���`������+�u[�;���Hz�P7\��{�1� p��k��*��p�@����dHY�����^YP�z���[�x�-����G�2��$g±e�U��3�aZic3p��+�����({
	]���J�O.- �MNTE㢾9�{௳�`�K�$��0��N��]AD��� ��ۭ����=�R��<ڢ���W��+��W{�k�u:(4N�nn���D{�rGc�dμ���w�qd�E�ۜ-��l�7�feݒH+;�W���#z�,'Qv�5g�^����v_��$V��W��p1�)���ʐ�5�xW?zA'{^��=�������<򫷕�U7/!l̐F〦��i�� �꽱`���5u]6E����� ��j� ;ڢ�N�&��u��kҳ��,��v^�3@�
���  }��s�f������7�B	�;n����wz���nu���trc�� �4�?y{U� �V̗��V�{ᖘI]�BDj�>P9\���L��_��5�[⺎�0�.���
ѽ×(�vA���7�݌a�ц�Ww�:�o�Hn�@	�k��1uՋ�73�0l�:�]��D*l5ۡ��v�u�q��'7)�ֵ�;66y��G���յq��w\x��g��k�b��X䫮+CǞ��]qz��%ݎ�{e9����&�N�3��j�s�sq��^^�v,H���Ņힸ*��ъ�
�c8�=[��aKR�Y��3c
�m�nϝ�#��z�т�Ev�γ�.�9)�t^��T�޷���#��m~�}�lg�(Ld�	|se�$����A>��]�4�(�oVV��@s�͡�5��S���j͋�.��/D��FjI�5�~�`}@T�kK�>�����(��y{0_�x��R}�k3�$��~��U���S�d�C}�~}����Q�^8dq�S
M٧��0U�UoD ����|�������O?f��>so.�'�\�0�3G r�m�X��5@��?yg�߳�|�B�y�~@�r�}��^��F���l�qCQ݇[��*>��`S\\���ϵuc��#!\�����s�n�i/x׮����꿉$���h�
:߶^�@��۰H����E��+ q�%���w��"��붷+�;Y��H6БT�e��J:�E8�T�R��J�Z��w�sj��w
�ُ5
\5LZlG�v��U* W{�� T�sM
ۇ�w��r�U����^ЃL�i	v7��w� �~{H�CQ�w7맻�<O���,N?<+�r8*��7�f���j^�-xɴPX��@TT��h {�$TW�[M�l��eY+��2H�	��d݂�_���O>J�r[���
�撠 ��|���e�>Ǫ��y�������ɒ^:V�6c��^}�Թ��oѻ<5M�c��̢�A{ysekj4$R@���W	:��'��VX!�u`��u{��$�q��w��LP��"���Vz�����գ,��|  u��h
�PIзi��,{�I~��#%����Gf�'����A�k�M���ҩ���̅���[1��Ʊ,4n'���M��z��~g�U�%�w����i�i;Q�d��ړ������5���edN�� �~yK��VU�������)�%����#���G�s�EhO�$��^݄mv�{^�D	>�}H��ऐ�T$�}6r�� '�{P����\��D�,�@��IP>��UC�?G���`����m۝�~v%y+���Y{v���7�=�}���i�p6$(�C'�����-��d��u� N|�!�@|���Kk��	m_CZ�d�9�uՂE-Q������(���@U���\)9��| P#r��X'���,�����G��+{�����$@�wf��,Y$���`^5㰇��*��I|(}�������d��-l����v��=����� Oy�iUCnL�u�6z�����L��t4&�v�N��V A�Ӑ}[uv!FoW��B"��;�J��	�ڻ�֯���&S�]R��.��1X��:�a��u��� p��A��)�%ح��&�l�5�*��Hzp[�MR�y�R�ܙ�ػ4�˩߁�z��^����v�������8��f3^�0��wb��@Yj�^��c�J�'�.K�w?j��6�� �ug���쬮 ����u�%m�$B�
M�9se|H'3w]Nz�cw�)u�j�	���|P<��
B�t���~�|�T�Z�Q	�):��`$�͔	���=���Fv��0+�+���  ^�����P%	1����{o�
���u~.Q��uvU����(�Gvz︊[>ڦx��ת� g�G�,8�*W��v�����=E�Oa?w��b�7Ւ��u�ݛ����\:rq�}�ڏ:�u��+x�Zz�3�8/U��鞑�g%�0�.��j��Qü_B(T�YnwM��+�����~y1ԣ�\��s%�n�m���4n2
CM$l���I�l���(8����`�/gu<�э���n�k�C܉z.x��Ƕњ�J��� ��ūۖܓ͕i�xj��Ԉ�y�Fv{*��5�a�����룢"{��l�p;l%��q��V��]7XJe�:�8��!K�hܘ�����p��9���{����sl��լ�s�1[l�3u�,�RKn��&�=����yΈ�t����?��8�L)X�T]�/��{�� P��J��m�fo�TU޻ �	;��@�<!=Q���
�NR�������k��ik� �6mh�Q$ �|'�*����z{�s��5�$i�����}@���_ăS��Bfͱ���yY(�חvlꉅ��a�9�Uݗ.��40Z���.�� ��/��{�9܇���c�O�P�Vk^b8��2��˿��A�7�|ѩ�Ȏ���$e�ݓ�#;��E�{��.[�¡4U%�	��r&�j(�h.]u�s�M��O-��һn�"�a#R��A$���⌶Xp>��z�	9�]vA ���-�)7$r�͡@
��Ĩ
z)�-��b]��V]�I��Ca*m_}O�۴߃Fɿ��Z/��璊֏r��慔1=��/���Й����������ݬ��o��;ŕCջ�8�It[ʗ���-B������������AƩČBӆ�9y}v~$�;���AJ3�4{�v��E��.�$���:�� ���P2n�>w�_��32���'��r@ >�w���-��+a��eTO�{�vI�L-M��s�+  ���_�#O����~AC��N����e�u�==̠H�[S��r�眏�	��C;nI˜g=A���FMX#�Lf��V�$	BD�mmՂA�I$e�W�LP�gm�d��O���]���$$9L��u�:�9� r;�d+˔KƓ�?�n����>�Y�>��nݷ2����h�\"&Z-�.���e���ܠH$�g�U���:�3.p�6�{3%�Inф� x?�_Y���	���'��,=��*7dOY�ɣ<���$���xmΗ���-jʄ�^wH^޸P��O�W�u*s{��!�.��C�S�Ȓ�sɻ��܃g��&�˻Ӛ	�ptꊷ��n(�M���T�ʜ�2]LЉz��i��A�DP��Zb�炥��d�Y�L���~�0b3��|�)�sm���z\:���0�I���V8f����g\�|͛*��0�w�[�I/t�6��-� ��Kv�A���
ǡ��e%}��=uېx �6�םXQ�����Ū��FJ���N����(�t��@�$����a��JV�]�����:s,�=vŕ�`�� J��{O��9n�%~����@�e���x�sږ�wtù��~x�ܛ�h�02��_4�6=�̄Be�Ȯ��� ���l��ٳ2��0�YeWS�b�=��C{һ�}*��Ϩի�q �{�m������y�����bÑc��n��=�J>��P���綽=Ώ��U�����ֲ�L^<��zIjB�st�JVŽ�,�óC���Ι�1=�K/��U���O<j�F���=�<�X�D����wE�2e'�+6���
��9y��̹f�^�*X=c}�n��o�c��N�kp��,�Y��U�oYY#պ�#,�T����Dsy�ȬF���=t�d��S`��&�������EZ��_o��M8��<w=ǙsM��/x+�dR)Q�"�(��1���E��QF+#���A@PU(��DŐE��(����c,YF,���X,E*Ȣ���EAb*E�V+H�"#E�*��Q"�)TEPX*�AUb�EPQX�UPX�U�PF
UEb+�R(��)A��QT�U�UAdU��U��X,X"��R"***�X��(,�����ETTX�FDb�"�Ȣ1E��,A`�U`�+Q#1QX�*"(�*�XF"��,`)X�b�A`��DU��U�ȪE�$U"�EU�DX�"�"ň�X�F(�QX�X�H,`�D
���b�R���`���DE
*(��EQA`�PPPPUYA�E����g�X�>��֢�w�� �2�ZæI��Zp�ǯ/U�S�oíyj������ �~�E��K}~�Fg{l[�(�H�l�7`��A�
�k�k���ٛ��Y�l��4�P Po�m
y��g9�K�/C��*�v�pt���QΎ�:v;0l< P�9���.���iw{�a�,a�@�}Uy�d�9�� �jj�9eu[�%J�V�nQ���h9P�bP�Y��Y�o+����3���Up$�{�t(�H�����{h��WlWWo�	���O���[0:�묕�${�{Y��t�{M><�����(
�f� W��H�� �i�Ļ����Rͧ�S�^��j��h
�|ג N���5^�݄���RU웝Z@��U�J8���{��woJt����`�s��t{Y�V�̙Ϗ�l�=lb�6z�T���=���Oh#2�K�I��Zp�5�{Y�d���^��C��<�s��(�K�~9�S�{�%U��9�����{=B�����`��4���n��y{9��M{���&���\Vc�"	����iP��K�}�n��;�1���i�@{}}v	7ԓBaCn꫻.� ݺ�{Ao��O_�@�r@P;�I�g{|D�ۏ?��z�2�"ı�&e�~;�ޫ$~=WG"پ�����A o��� ��z�}��'�@�)���c����;֪��c�}�!@�N�H
�rՏчN��&�{�/�f�D�����ݕ���(
��Y��H���M@�Oy� #1o�}�%��2�z�*ޝL��|^��8L>��
c�є0���[�۳Ok�wó�'c�k+|����� yn�{7������3&�=4\�K:�9���hxãA�A�
��ɗNrht��c��r���ݺ���������d%|��O[�j�N��:{9��;eoB�S���\�F��O/+����1���n���;i�Okq�2��Ӣ��'3�F�nzy	F�qƁے��1�М8�<ݝ�c�l0��N�o\��zk*�Dpk��&���9�nm�g�u��굨D�-��λWk�ĩ;�7㭵e;�<]����p'���a���jq�� (I�z��>����۞Sh��h��z�	����h��AE�r�B�b�Bӡd8�n�(?w��$s�.� �&�̡��Ju:�����E��0��7
t*��w�$�w�j�`���n�yfy�x	<�������$�D-XUV�T�n��	^~�@|�s��@��L�VsE԰��候��;��'�DSi�䧼�~|�%��sx5���j��fn�
�;�4�u:cڋ�%�Ŝ��f�\��gizg�EW�6������	wc;��dS�N���Da#h6��fz��$�s˪�� ��8Ҡ��	����֒U@��YJ��!-j��m�@�����FӅ{�s�ݏ�S\bU0u(��+��ph�������T^T�i��̻s�c~��t��J�-�<�����\�tx���|���$���U�$����� ���Go��jл:�X�y�a�.�ʺ	��Տ��<��S_��ãø׫�mh�H;�L{���'�O�cbPa�Uw����bt�P��uW��O������$�:�wb>�I�]���G� .#IK�6�,Y�w����_V��`�ri�㺼��N�N�P��� '����e��M�� ��;��"?~�M;��lP{P�[\�2hܓu\�����;K�u���ٖ�����O��х����;�h��� S���íx��uܯ� �o��`��4�AM�{޺�'��y�����M��� �;o}v	;���$]P��Q���[k�C"��2�D�[qW����Œ@9�}V$���k�8H��{����dJ�\{��� h�bt���ì��Q;'���%�?�wS,�jF�*��|�G��|�WSr%YM������� �~���$��_]�|(�n#L5`�[c;��&1�ƫkn�$|O�ܼ�
�͆�>�a���*�Qn���a1�("F�NM�V~$�ڦ��:>�\�]+5>�%価C���P |#3i�������E��Mc�����nvi"��%��t-e�\��|�m'`)����M�o�@�F����I����$�Fy�*���&fnN�ʡ��7����������de6����,���(�� @D}���C��
���O~���o�]��6�YP*T�{���Ұ(��~��k05�A�H]o{�u{�{���u_W���~z3��"&"�n;��'}���m��VPd�=��d�&
IX?{�~���{�=��=aXV%�w}ɴ�������_y��@ yS.�e�(2 �G�����O�g:C�Y��+�$�T���5�B��Ӿo��&�
�@��W����L|����q~0�h��֗s
��e:�����{�~\�����!v��CFGw���c�iɓ��w�w�x*A�3u��`������������P�~���ɴ7��7��wqk�7����a���w�I��IP�9��{�l�#_\��P<J���]ɤ�`Q�
ח|�`jf�R��y�a�q�Wxn.����>w��ϳ߮2]�s��1h���,>��O�;�Hn0�mq�e�X�7��������[�,��n�Z�=ɤ�H,�����d�ɔ*J���w�{�i��Vϻ��RhN��{�i6�d���^��Y��N{?��e8�%,x�<G�_�����AHg����ɷ�~>^o=ɯ�B�B��<�u�M( V��0�62VVJ�������w{�}�}���&�0���!�0��`������?���00�Rz�a�{��6ͲXʁR�}߹���ߟ_{3����	X�
}ߝ�`k�B��;�y�a�c F�~�m�E7����{�{hx�޺�l�~��������������4Ʉ($����=�4�l*AIA߽�����~��څɚ�?R�<~�����z?]| �6��m'
Iږ ����8;`Q�h���&�RY��_t�M�B���>��Y�V���
������a��ͲTw�~������:o�w~��/՗@�A��`���f�N�9�&�el���Þ�gH�7�����`[��^�AƓ�����;*�c���MP绻����Xw�κ��Y��u�t	����H��C�鎋�(6 �W�'m�������`�;._��=հ�.��ɮcN��!+N�5�0�����[I�cѮw��
%:���F��Ӈ�rr�i����or�۶.��7a5��Yݲ�c���A�/H��E^��<�N-�����rQ�Ĵm�h�Mpt���y��Z�gmq���^�3�Ƭ��`��q��vbw�f�]a���ik��U�&
��!���w�
�&��4�_7�5��0�J�IP�9��{�c6�YP*T>�w�H,��ko/q��&��mq���`k��m�y�}�6�
��/��n�<��&�����M��+,d��w�{����ߗ~�>�I��y4Ʉ,IP�+
}�~�P��+T�]�M$�������83QX�˾���n���` !���2�D
�<@!�~���H)
Z3��&�H[HV��gNg��Z;���Ͼ��|*eM����m�+,d�T;���6�ĕ�9�)��A&LF���<��ow���1�e&P�(�a�k��d�e@�P(w<�tmbVk�y�9��ϊa湾g^�R���a�q�J���h8�I�!�� 
}�(Y@+(�YY+����hd��y�����3�I�=�+�{����lV0�*}�}ܛI�B�Q����Ϝ�`x��?^�_��e�I����?5���+����f�ʏV�7S���ͻ����?�5�<�鄂�Z�7�i�֤�w&�R �0+���f���Q�G3ˋs��s�4�"w�s�pd��%B�mo~��>�-�p�"Q�",�Y���Y�a%�1�������9���F�un�Ր�Ԩ��t=#��˙�RQ�7����@d���Շ�Y�EٌU�~���~��4�ZF�TF�z��H@��l1��̟�6�YP*T
s=��@�V�R���X���?�������ޯ���E|�`Llnxaǘ�u	��߾�&�`�Yc%ed����d�Ʉ(��D��Nzs�k�Ts�}�8�R
O�=�_w&�n!Y(ʐ^��k2i0�Nm���x�Q���G�+���׹��1��>{�u��R
����It�l`W���H,@��k���a�y����>��N3%B��u���Aa���K�h$Ɉ������G��P�B>�%�V�>�&ٶD������I��R
��;�H%`V�+_���f�H4�-��{�s��
���/|�|w-ĴH����
"�фT�(S�b�N��A�P��;+9���s�:������A��*���i�s>��AgFJ�2W���d�d�IP�+}�{�i ������AI�޷�rm&���+%e}��Y�Ȣ _P�#���bjX�d#����@x����鷒..� VV��|
BФ+c��{�j
j VQ5�y�a�ld�����e�s^�uϷ�Hr	+�Sxq�q���|�L6¸���e ��V�~�&�m��>"���*��c���yS��JP�㸭��w/鴶�e;��cbc-m/˙4��&>Rn� �G�eb�rr^����y˭gߏ��H ������
5 �=�Y��������s��n��MO�>1'�9 u�� ���g�G=��~�ܘ�9�f�*A]{�s(i%B�+
��P��
������I1L}��s��.>2j2�Xʾ�=̚M wON�����07n2ipJ�9�\�lv�����}ɭ��5ަ��!�l
�o�����@�=׿{�i�*AB�s��6��G��2~�fg�韯8�����PO�p��˹�Q�Tm�n��8v:\^ݵ<+�㞵8���]o�_�q[KO0��xñ�|�����MT�V�>�&�6�P(����6�����G����|� ������R��{�{�m�`V��Ա\)��x��~��#�H�,��μ��[{��ܞ>�wܟ�B��X���~���H,6¤�s��rm&�
�YY5������ons�g������ș@�=4��8�%����F4%a���r�(ԅ�s��Mn��)
�^7_�=����3�	�@�D
ü�}�4̓%H(X�>���hm%aL����b����p]Cl60�.~�C��_���7��<��2�hT�
��u��H(�_���F�6��F�UC��UE<_��Orw�f�ߪf��uc-P��~���GN�	x�,�Ɠ��V�1����d�+��\�����s��>gܙ��?��|%�������E+��?�bpHC�3p0�I�~��M�m��y�d�Ʉ9w���9�u�I�%a��߳0�
���}���M�VJ��Y]�ۯ��! /v�^��ŏ��"G"9�+��n{�,�]�v.�P�Pt.�= ]��H�&����Q��Q���q ~#𯵯�l�P;��5��*Ak��1����
���{��}��dNo��a��ͲT(�{���i���,�,$����~����@Y�4�
�<�{�����/��:a汮��f�+*A@������_}�w�NE�_(m�w�?3ݛ�|����������Ա4(�W�Y}��^��l@������{�k&�<Bĕ
���<���z+���g{�=�0�aXQ�@�>�ri �M����5�4� PP�<�1�TQ5,B �B?۝��㾜�:�7�<��R����&�R��
�}�u�5*Ae�=�3���|��������Vhd�X�����i�<��F0_<.ๆ�r0��k�i��(�ID+g�s&ٶM��6����k�g�aԨ{�{�H,�`V��1���<�R�w]�ߩ�>� }UO�9A����e�t_�]Ëj]�����{����.������MvZ�i+��T�j���,˼���:ym�ٌq81���;�㬬����,�Q=������4=�4U�Y}Z���BW�}�۳ި3�v��yGk9�7���Wb(��`�Z������H�U�2D���z*�����mp�^fg���?����~�x�QQI���D���M���=��̿��J�fpJ���sk��mQ�Hf��Suz%��8��G�
�]���ɸe=���R���h�4o⹬L�,_D��1��2�WB5���q3M�����;)��d�!�0���@+5�ԇ�u0:��z�{���UZ�U����3�Q_72��4}Q��,���t����������À/tnfKG��9���'e��]�N]h���X����c��/n{%a��8A���Q83��8yk�^�M�W#XH�g�������ɏ<�땃��C�H��6��	��.]��w	�}:��SXJ�ʈޥ��siK�oV�]����;����k�X�{��rN�����Nr��u�v�c�Vx�����Hgi5g{���;�+�L��z�Ŧ`n�;����-A�wU3NX��Y�=]���i�~��7�X�idv���p����Q�ރ��._nK�;l[��ni�u�c5�@W����NK�vgu�Pl9���`{q����͚O���-v2�J��1靲a��s/�������,F�9z �Y�r�F� X�ETbP1"���F*�`�"0F)"����b�(
"�ATDX��DDR,b�(�#b�D`�QV
 �*��b�*�
�,������,� ��`��ł�(��*$#"�H��,Q���"�Ŋ�U"��"(���)QDE�"��Ab�M�*�,�*(*�PF(��T
-����E�[ab����X������(��"�"�,H�U1D"Ԓ��+	R)" ��PDE QAV(�A�UR��*�`�dUEPX�*0F
Eb$G�S�H��F�d�	�@��#��u��=:�{��ԏ���>��)���i`��WZ+��=;qb�K��]�;v1��p�����9���m�pv��6����>�;�^R�]A���:qBj-�%�7���Gn������5�����'l+�Әء9����q��M�[c8���嫜�����Z����&8q��d^�v��<x�X�Q��\�/P� ��m�>0�uC�8s�u�,�C`��[����v��;fz�約A�*���q�ճ۟l������Gd�|�zݗ^.ra��&`8���yɓ�9���n�/l:�(6���g���3B�]ukV��FqF����� sl������Dn�>+����su��c�d��Z���6�ѱ��ا�M���T�wV8!��m�9J[mc��Ǌ�lv�Ig���n��rs�>/g`;ku�2�O=�G�p��;H�Ń���Ľ�A�۳y�P��h�"胎c�a=��[7;�9�'B�/9Iݥw;���:k�c����824l�+�nU6i�� �7d�bٴ�wB��������y�g��vC�B:xݞ�;�6p��l䗓�s��;S<Mˇ�'7W%�V�@�l�F�����\n#h�u���� �F�����p��]���xJ;�-��v6������
�5ƚ{p���۩��Ü��q���b�9�n�Rv��<�r��Wj�+k��plX���î;=؞v�p	�Gr�x��{=��w7n��;����<�WLn�������f=�SS�y{�\���(�X�.���ٽ%q��@1�z�W���GO�-��*�'wgz��Ҝg������Tc�H��v*`MT�,c�]ϲ%r���9ck�N㑶랞��Wc[OX,s�;�����s9Nh�Ʒ��W=�7n����t�4���z:�k�nM��zj4O<v���S8�]�M�u�(,]�-ӣ�����:�k���|���{ެ���|����t˸��:��H�R��N!��rg��&-5��o'�i61�?.�8���v��'Gj1�������dn+��v�7m�ݮ�.y�%ŵo9��%�-�60��:�����(��K����ق��5l�'<,p�hL�XwX�����G�
J�|�����r��O��x�1�:���s�t�(�C���>6�����7���n�%4gu��s�V�r[Ci��g!ntd	y`n.$^=��z^�q|ǎ'��?�O�$ַ�2m6 T�����cY�P�$��u�s0������i�~�8�Q1�wܛH,�Y,ey�1�ɤ�������0y��[�H,1���i!�~��'r�j��w�M$�
с^���`T��+*}��ٶJ��w�oG�|�}�g��9>C䕅�M!����H8��?�������%B���uϹ�c6�P*T ��W�����������a ~#�	���cY�R�B���a�c��yږ&����+��G��/hm;�~����f++%{�q�M2x�T��\桴��l*J��wܛI����gcz�6�Y1_��k2j!����Rb)�iƥ�@B?��ʆ�
Cv��w���A��}�����Y7x�������P*AM VX��_s0�6�YA��`�;���i���y�/4/ߴC`���L��0Dd�'R&f::�U'=C��=��C�\�������ߎ�u��p^�L:¾��o0*M%�9�}̛f�
J�Nw��F�6����g8�w��65�>ǹ���AH6Xg�����R��.��d3�f����{̛M���Vw�i��O|�^�"�m/�_s�s�vfڕ7M[��n�fȏ@2/ �>��J͂vU��0n5�A��Y�U�N̄��_��B�d�����?2x�T�ý���H,60�*s���M�M��ggy���sy���"���'D���Ӿ>;������F�7��u�d7�(ԅ���{�rkd�-)
���<������2w<��*h@�P+(���0�Af�*!�����IXS�c��<��h��V���
���̇�tw�Һ��>�,B�ǿkܛ���R�_{�}Ѵ�`Q���cy��<��w^wۋ�H>R�w��6�
���)�<n�V��bN��o&�
Af�+����i��c\��W�c�۫�2��%aa�g��H,6¤����6�hVJ2�Q�߼��&��Ʃ����������Ӭ��8�i�01���7M�S:x�[q���)��ѧ�;�������]�d�a�J�{���6�A�������i
�]��o0*h@���[�}[��>���f�*A@���4��%as�'Ǜ�Ï<1��.��W�k�i��(�I�d�ϻ���oa���d�f�,e@�P/9�}Ѵ�`V�+_y�o05� �B��{1������w����Ï��R��~����$��a4�Z�y�i�
��YY+����j2x��
$�7�ӿ��������1FT���ٺ׏߹�ݱU��+;w���ȫb���e��ZC�m��r\2�z�/[����}4���> ��9�0�¤���i&�
�YY++�sX�I���K��x1p��,�� ��+��P���k+2��D�{�M$����sY��ЁR�eO��9�m���y������Hld��{�d�2	�=�v�Z5�r����A���=�G�����Ƽ׻�}�iP3�{ܚH,�`Q���X����B���s0۶_u��}޺���iq� E�T����b���,��s��G`R�&�� ~#��R:�q�"����I�s\ɴ�͌��������� ���󙆘n0�=�wZ����7���Y��ɤ��+%R���I�� Dp_䠊}q�B�G����@۶�Ǚ7�w�1�z�u̚�R��
ӟ{���i�T���3�l�����3ן|�u����c9��@����?�anA!L;�x�=��#;}C$�T�B��~�2n3l�e@!��F��T��~�U?��X����ST�ie���9�m����~���o�`�`a4$�߲m=��|�]�~��2VVJ��y�C&��J����{�ja�aR
K��y�i=瞙�]�z���˛��L<����{ �FnoЏu�U�b������e�=loj�:�R�A�E9�4�A���Q7�)]���ʪ��~�~ed��y�=̚O,�ޗ���[L6���3���ݰ(5 �s�{̚ܤ/��{�}箼.�C.i�{��M*e��}�ff�+,d�T>�{̛CbJ�y�5�y�7��/�B��Vc��lH�,�A��N-kuv�������\GL[���p�k���߹9���|�/aXu�{��솘x�RPB��;�d�6�YP*T
�{�@<B? �oiyR3~�����k�-��m!Xw��3;i�~寧���.1[�M�7��y6�++%f�������q�d�1�s'ѓ�(��D������4�c
*J�w��M�؅d�>#�y����x{\��~�o���V*���3$"4�R�#�O���z����HR�9���5��� ��_q{��w��7�>*AeO~�9�m�++%B�9���6��V�O��j@�L;�x�<��=@{���C	<B��Vw﷘i�q��@����ѴĬ
Ԃ������&<��� ���ن��+K��߰�y��y��j3���M$q��﹍�����c��;<�/O��<IXg�y��laXX¤�{߻̛I�+%ed�+�s̚O=χ>�����e<�kѹ}FJ�|���X���dI/V�����cݟ���2�ȭO���{��h�{�2_i˓� |>� h���֞w�j�\��ݭŢ��W5��vsƔ����(u�ǩ�K�����/o	��'��]m�Wl���W����n�ĝ�,������^����ۜ�ZK�v6��Û�ܙو;lt�����*m�S�s�]����՝mN��zD �O.�ݵ�J���OH[������Ik��8�ۭ�'*4�l�#��xg��V^;'2��y[�
q�mIŴ]��8x��Ae���j�c�]vۤ.�R"�l�}�s� �Q�����Ea�g\�m��!K@�{�d��i
�l�9��H(����Y��N�[�a��͌�
���y�i�ϼ�s�Ǟx�%�຅a�¿o8�`T��1���y�����y����6�FT
�����F�7�(���ݬ��r/�_!Go?��Q��ߟ��0�? �{PZQ�bf#� ��3Y4�@��%e+Ϲ��CBJ��%a��W���^�=��7���+
0��{�M$����Q��9��K!��65"5#2� #����@G ����8���>$ ������!m!Z����7� ��
�'}�9�m��S���os~�I�m��B�w�#�O��u���Q�P��<�q�q��y�Rh�*�9�{�l�&�;��{|��iP.���F�
AH/w�k08yH4�-,7�y�a�o�#^&��C�9�i~�ߡ%��aYb!ӹ���s�Xs��1ۮ{a��\�l�p�s�&����c�b���7>\c�*u&q�~ɴ�ͲVVJ����`T4��D���{�u����􎲺��t���2>���o���B�Q����}�7�4'����ۇ1����4��+3�s!�l
5 �t�O:
knR�w%x���v��gF��v��!+k]�B�P�'6G[wER�v.���)e�;VsO��OHƛ�v�lֵ�@38�� ���{B����)
�[�{��M T���s��L�%e#%Cy�����>���1�y��C�%aNy�s�ǞTJ���*A{�̇�T*J�a���rlf�(�@�@�9�d={?	��h� �L
5�Z����`k�AH6�w��v0+L{�o/�����-���ؓ�{���}z��I�>�-���J�2W�}�d����*%a�}�s$aRT���rm'�sT�x��Y|ð��Q�������OW�X!�,F�֔0�g2��+����6� �,�w��&�)��߯y�ν�5�:�
��u�jM T��{�{�i����d�T>���M��%a��L����:�ϾǞYZ��W`䓋r��upsM�x��3Sh��9I{O�ЄO{�����LS������#3��4F$�T�B���s��L�R
�}��F�6%`\��;q���� ��1����AH4,>�9�a�l
�sܷ�b��b����cP*hw9�rm7++%c��s��q��w�u���d�'�Q%Bĕ���s�Ci��T���&�m
�`���]��sr��w>k��=��� +с^�`�|��� ��?k��`Q�
Z>�{�[)
+� ������A��V�_�K��(��t�su�ncF�-���j��w_{�ckt��m���w����)��C3�~�q΍�Q|�]c;�c>��	$ �_c�T� T��	�;�s�c%ed����&�ϼ�^>�xU���+����@G�]��'Y��y�߂"T*Aa���2m�d�*A@��w�H,ư+^{�o0>�7ݷ���)�a����v0+q�ܼ|�6⫏1庁��$���y6�+,d����cy4���sEt��ϸO�IXS��}�6�l*A@����H)�q������2 ���q�>�v�;��&�g��n������ۋ�z��c�ם,nym\�X�c3��}��`zb"����#���e㴂�P9߻�Ml�-)
�l�����L����0�y�+7湘m�d���
���y�hlIXY�և�q�aL;�x�<~�����Ă���_�h�5�q�w�����A@�*9�{�H,��Z��cy���A�����yM��a�k�fH+��ޑ ���ˎ��}?W��< #�+(�_���
���
���}��g>���w<���� °�*���ɤ�������=��4%@�\=5�0����<G����+h��s�^C�HR�3��!m!RO}���
AM�{��0�3��r��q��۽)914{U�Ǚ�cf��~�^�-��x%+<��t�i����m;Տ�鼽QӇWZd�@�;�W�������$�&��d�T9���M�����u�py)��:�a��7��4¤�T�
���o�63l�g��u��tr�}�@�%@�����Ĭ
Ԃ��7��R�K���a���wG��<?K��|Lֳ	QH\��r<��x�v�BM�����c;�"��?_������q�y{H��u�I��VJ���95*%B�J���|�4�p~� �<�&�?����?~�2 �w��,��B�K_}�y̚�S>p�<�q�1�0�FP4%a������������f�B��?eЇ� ��~{��9���
�@��}�o��ٱ����:cY�~rc�w�OP�J~��0_�RD�@��g���Fgz�aRQ
��Xs�o�6ͲQ��@�}�7_��n�����R�}�w���i��w��3��
���Rq��q��"/�>s���?k6�cx���f+(�^�^�&�%Bĕ
�����桶aXX¤�߻�d�O�1���~�����&A� ��=U��,^�Es�TX� {��{�o!�l
5!e�w�w�5�B�w�9��gǤ=y�y�sH)�
�'��|�6��J��P�}��&�؏��{���h5e���Ω\~���Kh*�n(͜ݗ���y��1�S�o|��Ⱦ����w3�����K�^c�x��n�i�$?y��}�>&�c-�+Ew�;�|�m������KVm4��y�D�	a��]n����=�b����[��{��m��-m��X�ۇk�ٳ�;"ϧVh�c�<r���w�<��O��Kۀy8��Fږ�]�1��O'1�6u��:��J�����=3t�hC�q��n:�	��a1��2Y��[��e��N�ݣA�E�qpn��n�v���vъ�+GnQ�z]h���� �$�v�:�r<���Fܼr�G$'��?��ђ�8���#�� 0��߹�haRX�IP�9���M��%e@�T
}�{�@ؕ��5�{^slc^sﳘ��JB�{��_���6ʍ ��+��>����1LUQ����7�aG�C��}��"��>�M�%B�*IX}��m�aF%�߻�d�Ad��ɭ�u~����q�/�W�Y���+AX��q�0�FP4%a�����I!��=�{̚�HT��W�{�wX�u���x��q�
p*Q��{�{�a��͌��w�ɤ6���������<0�_?�9]�+����w|(��T�
���s2le@�T��K#�O�x~ow*��ݗ�ԩٻ ��w��n�i{��ϱko�珗��\w�d�p@���YFJ���M�y��מg���mRV�}�a���c
�����2m&Ь���2��=�dЕ���|��y��?��v��ps�vh݁�:�՛k����[Y3�64�1a�$���\�2�k�tn���N�Ԭ3����l
ԅ���y�[
B��+�s���R����~֏����ֳ�ن����*���&�ؒ��y�~[��x�0�c�P�40��uP��">@���q�P�������ԗ9*K��c�\����^��f5��^]����,�T��g�f����P}��۬�n49`e�{��{=�ޤ�.��@�a�k�r~f�
��{��@�%`XԂ��9��iG��������>[�����_Vv-/���7�.�m7��y��H,�%e+�}�rhd�Q%B�+���{~�Ǿ]y�CL> ��ϻ߲m&Ь�����~�̚J���^>}[�7!�(�,�~�ܠ/{|y��W�`tjB����]ɭ�����
ٟ��H)��YD����a�{Ø͝�3�d���P��=�M��%a{^��M�B�]�<G��꺠7��D|~�TE|A����]dz�Ţ��Pn~i| =o^~M*7&���]u�}���CiBS��Y���.<q���z��k;��;O�A��/�SؑI�;��$�3}(�I#�/�KU[��|j��6on������V,��Ğah��t��d��w����ڡ��}X	 �@��P�A��/�d�h��)��U�پ �Yi��(B��U�(Oǽ�� ߷�̤Y���2�a~r{+�y��k^�����}<�y��]6��^������(t)	y�͌�0aG �ڷ���;ɯ���k�Rn-Swl{�w�k��.k�ُ�9��ż����U<-:�-m�[�#��Ij�	����ڢR=g����@��}�Ļ�zyx�s^��+s��y[�/��xaz�պ�J��Ey�,��;6��"ph�k��G_�V��wp!�j�qmy�Oy��w�����j �K�٠	���b���
��SbX@�N�ܼ�k���Q{mV�yO�E�(l��!X�S����AW�z�qI;�rZ��=n�|^,�'#���{��oeC~��Z:��\�3<n�Jo���zWV�^����,���!2����i��+����c�Qo{\]דENt"Rؽ�x�������Qv�BS�J�d�Ҟ���:�%z�V�4�pW`�tH�5� Ԁ;�of>�0V�&}�|ј��vR8/�YCN�%E���sH����p��(d�k�wl63��:Z�sڅe�<��r�F�j쮩�q�f![���|L��-&4T�W[*�)n��񁐆�!ρ�n+qE���=|k�<�QO����s�\�x��Kz��91�5��S6ݩd�Np^o�S��=�|�Z�\y��i�G{ǟ|��b�z�v�s����|����QK 4ӬG��7纡d��/d��i��@ls��{O�U\� �;o/�:���u��x~�;�7�w���s��oݩ�*�Q��(�Z��)PQb*�QkPX��"Ȥ�TD`(�(���1QE��m� �EDX�V1�EE-+$TTX��V���IX(�(�RE��-������EUUAdQ�H,��$+E,"�H��,��"��*�
��+��(�d�� �%�H,QAE�U�QAT�����"1V�X��Q���*,AE��Pe��d�b�UX#,-��b��Ec#E�Ȉ+V*ł�*(�, �b)Q1U�0�#���b*�Q`�V ��"�"5�Q���`�"ň�X�,+VPDOĄ g�k��QG�x�S����Jy��T��d�]��]ןq������g���m� W�M!C�z+ͻ��$����񭻕�"��|�H�a�d���sH�}ޚ���dJW�K���6�mo�U�&�P��>>�ǚ{���m��2mD���l�F^k�.Y3[���eۛi�RN/���h�I�L�ˮ��U�Р'�4� ����U� �R�[��~���=p��$ӄ���^�x��o%�{�4� +�މU E��C[�V^�W3�p�@�FT�3�e�dw{��$���z��@����^�~K�>��E��4D!�3v�nf�~�T	37ް,�{��|(|5ǝw�t���3,��.�R�g���V?/h���<}�$��n�o�[��6�ܪ��/���MY扻����K�V�J��R���օ�v-�{x�+���?�^�]�R�i��`�"���z�	���C>�츪�^˰I��uY?=���&
�*X�����&޳Ѽ]qVX���v6n����!�Lۢ^ˮ�$�#}��ȘQDXq�8��=v>��P��$	�4ޫ��X`�Gg{��=sZJ�nB"2��>�V��y�삹��2s� ��?*U@=����s��l��x]�S�a7�	�������$Û��A�6��|yn��~'�}�g�}���|+����
2���bc�Z~]Y"���'��+��$�|� Hޭ��t4�24>�뿉�e�XxPP��7_���]��P^�w�L
�'��:=�{y�6���~����,�7�{�2��^E��'v�{����-�Υ�3k��t���9��mc=�0���:/_�T�QkX���$qwh~����ꎙ���h�1��(��c�mN�s�7��ɋ���q�v�ױ��Mmx���"m\z�M��� ���Q�eݓ�s����V���aݴ��j�X���8�q�JF�L��,�*<�.k�r�g��X�L���n�Ŝ<�v�u�>;eK��O�p��uKѷ67��Jc�Pݳ{r�	��쯓Ք��u��<ѵ���n���r�e��N�0�<s�r(v����Nö|��Geq1"� �O�{4j�ی���E��yX��@U�g»��*|���io0ƽ��$a�y��_*(�3%P�i
�?*��)�>��@
z;�({y� ���g�LŞ�*,��@�!�v<vV9;}b�>�^�W���z���B�&��|GN�]�GTI�1G'��������ݜ7SI��ɴ ?6vz�Oۻ}m�Rs�<׳������/]t<+����
2���N����{���Y�+�7~�	e㯉=3�VI?v���>Ly{��J���	�U��ɚ��k��R잊����S�l�-s����'�f�a�EC�P�'�|Ҡw/%Bf���
�$�U�({վ� ���R�`�"���՗�u^����&Ǫ�D��}��A����~$O��U�	�����t﹢T}��i�=�;�����a�%XJ��f=|�'BH�}�ޘUO���S��{��8�c�k���p��vc�Z/��ˊ"Ì�2�n����A��3�w=�xu�'���Y�I?v�����4R����B���ٝ�{��T	+}�(n_j�P� �Һ&r��� 4]`JI>H �g]�M��P��x�vT^ �[]�}�|P��� ${����7!�Jʲ�K�@��b̜k��t�}Ϊ7���%6Ä[j��e~9�����
2���=C���uYE��1~Y�t1��}4��P�=�ͨ�zT�J� 8*��@�]�`z]�2My�p�����`���U�6s=P�y+���U*D��^��q���E{�=XI ���B	/�W�@k��d¥6b�7]]h�Z�,@qx�w�hr�Nͬty���%mx�t�w���z��[Z�u�}u��X�1�1����eg?�w�]�M��WЊ�KSQ�E��e�P��4��>͛�� /'6�"�ސw�޶��3c��$ݞ�bf�H�JCdF]��j`$���6 }9Q�̷�@��۰I ���H��z�񺸷;�m���P�c`ng[�����nG�u)��<��cBݱĔjZ�C;�'���|�,A�e��C���hP�6�'@s�X��C��=(]m�"a���w�+/�d��{�MA���M�亲A���*��m/�
���#o a�⊁���L�$#A@k����~$����!>�)ݼR��3	�/s�(���z����9�$W{ެ��f�U�m�:�hރ>�SΙ�=�����˸h灲���]�^-	�F������Oh�n'�G��!
��^�4��a�]U����2��}pJ��c0�F.�:�t����.ѧs��C)`�����|�|~�~�
"���\jAl�2�~^搠��jvF0aT*�,� ���`�s��vv�n��}5��UB��7��7�pȜg��e���dy�gQ����~'t_B�=�ȥ��!�4#.� G�ܠIͽ���s����x���ޝ�P �u������U*8�( ����{!�gy��c�m|E�����~�����+�o�t��[G�q8�nJU�:�,X �u���^
�C~��|��(
�Q�@|�^Hs*��0�T �k���^�	ᒼغ�7t��
�;�y/��>�i��^�p���Fu�]�	�g����E{�=C	"�}U˽��l�� �ﶅ����`�(R��%��<��)Q��]��ӓ;8����'�:TG������V؎��3k����>�Jc=�U��9J�C�=9���� �Ex�+4u��T�Wv�z6��9��x{!��۴V��������k:�Ohn{O8�7e���v�+lv�n��6o����rc�˻)+�v�f�o/&���A�������4���e����uv��j��]c`��5qs�b�G'<�ں� [����gn�n�i��.�uZ.i9ׅH��-��ݎ".�+s���6���"ӏ9��˫�[��K-�wg�.���0\J��K;��ghٲngoW�?�����.������Y �m�_Đ@7��@���z罷`�7:��;M�%m�#.�ڷ@�^���ѺivMmP�*��y!C��yZT�.S��'����X2�@�5���H?g��T��y�=�y�ey/P WO/%@ )��V�G0��_DіI�s��������;�u`�	��zP ��[�4��].���z�m�ׂ
?������.��}��d��k��>o������H;-�	����|8`>\I 1����1���iz����ܒ�j�&Q�b1��f��P�.9#Iwپ���������չv^�`��y�0�V�4� 
�=�6��$�@�l�#�ם�s}���>f���ߙ���h��f8�%����-[x=�bx�'/��]q�ȃ���,�*Ω�٭fJ������e{��_��~y�U���* ?�n�|��_ĉ�h%i("m�wdn����[�d�z�9��;�j�7\��H#=���7�rŞ�Iё7!�{�Ru*z_P��v�h�C��� '�yd�J|�y
o{���w�.E�Mvf���	B����]\���M��
!F�t�Aͮ�}y�}vM�G=r �a��"��������ltv�%�v}��ųت��s{v���d0�$�sBL�ޢR��{�&�J�P��څ�?p��Y���$f�z��;J���$5{ެH�9O�F��- P��!B{���A���*����S@�=w5!�8�IA�μ�Ff�U��%p?-�46�eJ���u�Ʈ�*�y�ѹ�^�Y� �ASÂ�#�W�x�c9�
�Q�j(�ʲy��,Kk���� �����A����d�F~��vH���V�f4�vͫy�H:�I&��� ����^J���q���1YC�~z�
�7Q��D�W����H#=���fe����� ���@B��/Ju�3}|�ݾ�CE�v�6�B;���m�J�cF��'�����I1�9Ȼ����_��*��f��3���?$�G���o=Uʦâ��w�_�yy*�w(�f͉@F���"=�2�������{�~$�ξ��H#��P�~<������������;R*���$5c��.� �7��_ %zn^_�yt 
��y/��7�D��I�"�&R0G@���U{S꾺~#D��> c�M�@P9Ǖ�W{�B��-����kH��g��ͭ�ː�?e�5`�0�S}SB�K��'7(�:�o�u�ɰ�ވ��53z,�ܕb�Jp�J�3A�M@���W��O�Y��w���
Á��bB���*9�n*]1o4u�W�eP�B��v��}�oK�zY��3̳�=Ȕ��r��n\��tu�"�rt�@z�H|�g\����~��ډ�¥.]�y�PQ=�7�(���y5Խ~̋�p�=�tR[���@P�窍���Ȋ1�d˰gUm��Z�Ԏ��[�$��JwV�Y �Z�,��E��Ri��L������� ��˲	��z|�
�w�֧�[��ۃ�=;r쟫q�c2IRCwݕ�h���Z4րH!W�}o�Մ�F�o_�U{��KY��J�9wƓ�Ȝh�2���H��Ԁ���g���*%��yd���	���~$v���7�۝a�r��Ck�1�Ӑu��`�M9���s�ze'Nؓ&�v�Q��#��Ͷ��~u��.�SW�5֔������V1�`s3�����	��o��j�γdYE�)��ObXV����η�VG��f�@o�I�_T|/U�fkP��ڐ�N���lP��s����m�*��c���V�8ů-��pQ%=b-g�w��;7qQOr=9���yX��9�'5L�\3O�fH
�{U�{	��z��2�ʘ}K.o���E�Y��2�����	h[��v������~z��Ӻ�HZ�U{4L"��=��uom�\�0�^�Xz��ư�x�c�r���r���:����zb�!�ü��4\踎umy���
}R�gN��_<���X�˂��LN�,��hgwԹ�yb�x��9�&�� �B��������c��k��jS`a\��bu�EG]S3�����VIG�C-�,��Ǳt9�K(�3��j�V�|n�QN�)�ڃyJ�j�yu�_|��N�z﫶�wL=��p��eՋ��W"�W��sn�:D�n��k(o2k��� f����-L��[g`s.�Qw�!v������e�^�|�5�O�Ń;M��εt;;���mul�1�n��ͭӒ5�YMn�3͌mۼü�d����d��x��>�j;D~�7<�t���}�x.ݯ�%j|�˻��ap��Eǰ�1�&4EsZ���1>!�7^gaߧ��9���=�w���7���kc{w�� 1"�RDEY�*��ŀ*�� �,UFH�,V*�eb ��+`�X ��UE��E`�UD�TYR�Ad�*��QE,P�
#@Q`�*(�`,X��RV�DE�I@UEP���E�őD`��(�T�T�����Qb�XE �X�",QV�1E����QdQA�Ad"�)AjJ�X,R"�TE ��TT(�QV("��PPR#��H��U"�EDR�
�T�*� ���DUFDb�,R���"�ETF,�E�"���۶��������:W�b���6մn��W"m����&ү:�8�z:7s��79�"]vsЯ@�v�7�۞f�NwbN��8�O���qs��m�v�D6��g��M�#c������矚�I����'���\I�(iջp�]�'+���::��n������eC��W/m�t觏mv�kv�4u���g<uvh�Z8��##ջ��}�m
y�w[||r�o���r���!��w��9yEz.c���Kv�8b�[Ŷ9�tƎ�4��l!�<g�p�Q��֑���θ�vH՝�ض���8��M�u������㎍��]g7C[�g�Fܾ:Ť���;���*��\rv��v���;�Z�у�9��<�ƽ��yԘϳ&��΋Fc�۷1�uX�\N�F4��;��t]vX�v�ˎ5�y�ݸ�Y���E����G�2�"��m�B\n�Cx�n�mv�{q�ヮ0v��v�5����ua�z�v�i�s�&h�`�r�z{6�n��Rc<������Bvy�`���7gFAL��Nm���q(��zScs�ck��V�{[�,F��&��-�:�m7/��ѷdG�aݞ�յ�z�!aW����]���]Qp�q�{I����9����t��m��j2�z��ь��Qnݒ�ϫ]�� �a+kv�c�@v�%�c�]�����v6�s�V��vJ�;]ӻWa+��g\n���u���m��˞ػB�Y�=npmf�Lm�25[�3��7m>���&J<띺���I6p[1��\m.�x�qF��k�!�\X/m��8{0�9i��[�3j�76������i��áyy��W�:3a�p�l��n�c|�.��gV��i���;۔ u�q�
F;r��ݓ�;��{f��������ݶ�[cf{5�&쁖z��x�]�����=�흨�uz5D	���k;.�n3
*6�Ʒh�2F�ˆ�y=[�) ۜ\���&����T^]��u��G���b��z:�[��s�.�w��w���_'t��}�����Y����N�kQ�r��t ���γ��u#r�W�v�nu�wWC�1�v�8����nus���x�t�%�qc!v:�{mlcm����u�6m[sRv���k�A�8n$�Ż!�ݍNJ:�ֆ�n6�P���я��N�|��Ɇ3�[�CpC�5i'��D�mڢzk�μ��%���#�t�W�8����9�uu�ٳ;v��;��#�Oj5ŗ=0�c@s�M�6���!���� �H�2_�nU��'o��$��moU�=2���?����s��A��JC��-AJ^��̧���V�Z*S>����?4������=���m�Q3�*�H�1�.̝YvI=��V~��ruw0�N�o�Y����$�h<
7��!gN;�
1�tG�:*��������y+s|J�ο]���
�-I$9�*�diP +�-���/�o�g�� ��� >�y!C��-�E��?t���ap��p�$��
&Z�I��lX��K�>m:�VN	{,\sf�;�����Fc� h�a�Pm�_ )���P(Pk�m �w�B�}��Hݮ�K�$бrD����rV}D�z�F;g��'A��ԯi�	;q̼�[k�$�|v�	.k����G�o{{��rh˾k�:߆ՎA��QT�R��B�w$Qq��념H>��'�~����!���{Ǔf]��oA#ʱ���$ �PP	�����O����A ��zf��Q̿�uv�G�����^�}G띍�p���ɗ`�վ�t��!@�Uz�W�$��nQt��'����L��~�z
M4!@h��*�3���̄����G��t,����������;��v���SF�D�6H��h��-�~-a����}��v���Qvlv�c�v��ﳷ��f��hs��ɞ� ������I�}�V��b�H�9��뿉$�{B�WxqH�2�4r���~i��浀 �K�A$�Ϸ.� Cօ
����f�����ݑ�wTA }�vI>=}�1�hg�����Ί��m�߷��u��[{�c��VV*�y)��Z���yRdܺ�{ªƗPK��WWp#��_oM�9^PF��$p��'��E�Vm�{d�8���,߀�)�$H
�/!Z}'����>�;�mQ�Lh���R XbX}&�A��곝��w�=���\�
�<�*�C�ܼ���c���p��e�R	��Q��-�u�vr3��v+����-ԉs
U�&�������)4��RP����}Dd�d	�۷�7ceU���aU̡@�Odܻ39�rG�CW���A��wy^�8
F�'ٵ� *���R���ڀ@����?u]F+�u��i�#BR0GF��� �m�X$�F�����M$w&��#ݷ�� бrBp�_vgW���:��K� �	<��� )��bݶ��s��wl��ԭ��
�ƃ]w�:�j�0�c@��Ƿ���m5�U1�kM�*���v��/�OɮQV_�����n�j9�m����w�?�V�V����2�)���${��łH�fP�ؽ�ϫ��r�䈄2Ԉ �O�AA3g6��o6��[��SdBm�H14��5���
���x̪�I���� �O�ՙ(��C�mGv����9  ���T "͚�$a@��UD��"�Gb�VP�H���J��G�� �Y}���-��8+��Or��"��R3v;����I#7=CG`{+��{^y�
��� �G�9[`ӎG
��Ҏ�^w��_�>�ޠ � �y� �|�&#�}⌭�T^����˰��(D\��$*����ڬ |'�5Hi�w��|�B̸)�l�i  ���VP����*���`��'����N��PZ�c���ր�MJ���6�f`�T�UI�wFO��mo)xC�z�W�9�Z����N�v.vq6yy8��l�v6�ܻ���N(:��&�p/^[�r�Xt���RĊ����;1Q��O>M��]As=on�3l�Y���x�����3�䠗��z��:�um���6㞏�-����mu�|�E��^��/�{e��Eɴ]CE�QMku��*��v���&ފ{Irgl���g\ιz��7���Tշ�6��ӫ�k�۶��e(���Omx���.5دW.�lv�3�w/���טpF�	��竁#�4�{X>��/sHh_{%g+ͺk)j�J� �p�<���b\!��%ْvR��6����  2��~���y�_
���x�V���)�F`4Z�z�}VH;����}���7����ם�kڰ�H�P)��꤫��P��;��H7{ޱg;}�-4�
k�Ag2��FmX��B�.4��ٱ������:ɯɵȫz���{�����	׽vW�:9�s���Jg!�[p���Czv�<tld��O�'���I��i��~8��"��<8��$*��.� E:$( >�]�i�ݍʉ{�(/�Q7}�vH�5N9L���n����}�ǎi^Y��G��v5��*���[���g��{0����CV;k:�r�Om˲.a���T������Лa�����z�&ׁ��uJ �O؉?��]�� f���%�z!T���n��۞H��@���Ļ��7n���j �;�y�٩\W��j�C�˺쟱{	E��D��6<:k��EC��h$���Ou�]�~#s�݌����Eq�?Y��F��e0����D� >��A�N�i����OF�{}�J�%���4}��h(mK2jjv�e�k��6oNc����t��޹��$C>�{G9nq��^����� 7_U� ��6Dt�8=��*��fb �����)�d5EQ3� ��2���t�OϮ����� ��[����iI 5Rں�U�;�]��N򳡧m��d ��jOu8���7}-� AWʢz��Z��Y�=S4�4�"MЫ�&N�G�Y�/��0�]$"���ӛ:ejr�����'�+�������1֦s;�a��cM���H��{ ���9f� R@�pܰ�u�3G^�N��� z��q�3��� }���r�'=�/�o}1/���,��DB`�`%��]�A.��5�7���ٰr�O���
��I��-%d Gvn{�� o���s�x�0j2�I6%ys֔�]�;q�*�`wc�9{g�[/V�7nlbE90������n(���Y.�I$N{��������
�WS1?s��r����D�	/�{�ݵ�~5$1�E�Tu�ۙ������z��W�_� �=I&��ѷD�d��-[)T仳�6Wgd�	'�h�d�$NE!���k�r {��y��˪����Tl�����>�m�$	��٘��>�-`'3�b�F����A�'3ĺ�� g\�Nb"�����o>���v{�^4�U����3��oH����#G}�����}گ+%M[���ox�L��{��-W����ʘe5ĎH��sx܁��UR�3P�Z������m�N\Tl㍜�M� ���� H�}M��{�Mқ;ӵ����A1�Fp���3�<�j狱�u�N�n7���a$I�{D�Q�0�5pI⼩�a�{�� y�1�t����
3��� ���h��i-4�/h-췤J�w��`�i�9�P�p�$@-{��� F�O[�";+���_��yl�������.����}��In��"I:�Zo��9��,$J��fb@ ��mH}=�`'�J�j*�2���3�nޭ��`J'���ɢ@?{�yI�O��c�<�f�h86�5%���	,B���܈��o�+Ϯ�7[N�o��Ы������b�Af���I4w*��U���A�n�^z�� 욅�&��n��<�����[3"���Q��i����~��#�6�6����]TЦ@�MI�Cn���{��U�eT5�5���.�Ӈpvq����a���ػqna��^x\�u�iL����;gv@f�۳��z'^�T������@���|ɫ�bZ6�Q�q�؋Q�w=���l��1cr���fK���M�&[�.�5''+����q���ZÉ�Y&]ۭ<��[�>��,Úݍ��'Iƻ1�:\;{=B��N�i�De\`�a9ut8��a��l��w����B}�
Hn�J����A"{���4H7���M��u?M�^km >�}h���2[(��L�$�^XD��3"F�q�Oe�0 ݕ� g��KD���qw���%��5��ёvާ�a�I��wt�%�j+H�˭�h �u7�@Ì�݈f�-Gr����z�J�W{ٽ�J&���I$��X 
�=��=~�tN����M��I!(!p�tL�,$�\���:[=!��f�ۈ��Û����޻��8w�]������� �~O�$rBb*�m��'Z��Rs���;�utQ�,���'8`�֢[��R�/=M�  �kn� w�Ͱ31�Ӷ��
�2�m��)�� �����q$K��5JQ49�ͦ ��(�?*��>8o/��#q��5���gS�O.���p���T�*f޷�7Ω\��
�X9��*��~*jHZ���Ok��V�z�KyW��z{.X��uQ$��C��C� �F/�Ĩ��V)�$!y�(�4f������~&+�k���%�.�� (c�XA@wo�h���ML�L�$U-�ޖ�9�/,#��I�g�� T��%D�;�r�k�����َ@Cm�@��=S�IQQ%�>�6� ݜ���{k������r�;�� #}Ӗ�k�h���s���
��i�0�q=�HS�����
6Ը��������U�qߟ������EEUE+��|� ;��l ����4�����"�a�_���w���\���mh�ٖo�6�]��9g"��r.����, �'�=�o�q� �/�W�:x��[Ʌ޹o�D�)�(�Q����Dn�� �J�����W����>���뭪��v6+��ŷI9T�>%u6*��{�����v���,I"x/�M闑��Cbz2��t�4^l8�A璱G�l������c��.w��ѷb��HCvi�)��r��_���NL��enF$�3P�XR�%�e��{:�+rs��c���'�`K����UǈL�J��Rf���h೽��j쉊j�N�6����}Is�/j�Rz@��r�D\��Wy���pg�>��q;�����&������3Nɫ���/�:���r`E��oc�[�t�]O:�����`k��7�s%�WS,�pD.�p�Z"�tc7;��s�E~��Aݡ�U��}�Q��Y��6�t*�.��v�4A�q�!T� 	�]��5��#b�[�/���R���{Y�U��R����}��qt�⺄�WV��9Wf:]����!ً����C�]K�j�FJ�{v���s�oK�=�~��s_�;�랎�~^X}7vg��R�A�KH���I��սz����p]����a�n}{���ޑ��)� ���woj�\qi��~cĆ�WU_W*�W�"t�j��S1}O9��o$�m%V/.zg���[HH�ܤq��ʕ^o��@�'Y�d���1A�k���̩���~g����VϢ*?��G�C{N�,��@�ؚ�rU=<�F�!�&39�	��Mpt�鸩E���^�M�;`�<����+y�Lgw!����Yj�Өa���7�8�G�љ&��cW8_^��U��%��RUQ�_b�*��b��dPETAE�X���X��b0Q�U�Q��ȱb6�X*�ŋTTH����*��PX�(*��0(�U��`�Q�b��l+"�"�Ƞ��dQ�*�2
�0PQADTX�R�T�1b**(�Ȉ
FЫ��QV��E-��2"IXT�
�-(��(�,���6�R")Z�QH�Z�XVVڢ,m�R*�*%�E(�("
��am��#���QRҢʕTPPYR�J��-()Ub�X�J���*�(�E���+*��%EJ�U��b�������֢��1)�V�l������D�U�*5%�X��d���(�5�J�b�F��VJ��C�H�Ln�#���y�� 7�8��f�6YC��a�Ҵ�.����vvzÞ̐>y�k� ���D?���jg�Ax`6I��Uo�v���*8�2"���ƒK�V�=���~�\�� ���� ޜo� �!�޶���.�ڭ;��)>p��}����X3�v2�۫�nu��˳c�nu��Ͽ���N��/��" �oUU�	&��Eh��/�o������� �nC��E������$0Y9�V}q%��{�=~���Z� ~�zWĀj�g�X
�r�<�����e�}� �N#f��SD�S���7!��޹Eb��U��cپ'~I.�~�h�o˲�D�e����n@�QZ�:��#}�N;9*m�7BD�t�����r� wo���l��sp���ܼ���[s�K'mNm<*KOn��]w��ztز�|Ы� �1����U�5|��`z���i|���!!���$��FՄ�.�	I{�7G��{ef�ce~�*$T>�� ���cٌ6c�p�2��R��r[ues����ُ.��dk�e�L�'��sPy��{�9k�5e�	y�=�,�m+�N� ��m���9���ų���6� ��7�����U5IP�;;ͦ��8��=[Uj7��z >]r+D��O��  �W�q���٢=���!M}2��Rl=�w/�go��@ q���=��~���Hz{$��ܻ��/�s6�R!"l�%���4����@���, ]=TH�nSznb��T¨Ў�=o����D��3T��CZ��L �ʶ�+����W���.���@ �|�C���})�<�r��%��mu�3�se�3��n̹@ ߖh�ß�Q�c������^��%�qŸI�Z���Q��+g��Kl5sU��ED!'&@��[I;e���ڄ㋍�ZyҔq��<e�d	�W�{/d�Q�ӱ�^H��\F��'���������K	��y�����A�b���-�ń���y6�v;��;6%F�c�����c��!����;v$·n�d�c
�`m�v���؋�.�\,mu���F��ryݧi�v��p=�kQ��h�4ݞ���U��ݸ�'�'Mu1��.�U㌹���7.�f��:��B�Z.��Eg����n\�

�D3�l�\�����| �=A�L,���ؾ���cK ��Ϳ�>aT������%�z�M�O�:�؉�s�6U��"��o��}M�� ���l��޿�>7��RQ5U$�MCh��6� �긆�Adcl�ǈg;��u�T�D�'�I�{�ɹ�i-�͉��%����� ��^?�A��m0��n[����ڮ��"r"'�����8�$T�*��*���� ����v��-�b����Dn�7�@ �|ټ����hJ�p�U��P�!��L�OT��sn��>4錶,B-�K)����a=�SUH�U:q^~m�DwvU���K�j���Y
��`ħS�D�I���/f0Ke���Vt���JO_\�K�j����.�W���!�D6o~�r�&�$b=a��@	�*�nY��ymK��u���U�D1$��vbc�Ǆ]�����& �;6�D0�)���]'s�����=�,�T�@TTD��޿S  =/[���]���.�����ͦ����*븎ﰥ p�#L7X]��ۭ�.�S�^<��
��[ ��o͓`%��T ���6,��V^lzwGz�Q6�$�\�� �]��j���|�zj�|y�>����N$��j "M:$��TI~�I�򆾴G=�yx_���Ϋ�X������a����a4����6�:���,Ɛ&Dɾ�ˑ�P�JQ3~ʾ_  8��� �wy��_U�Y�OF�u�M��!��[��(��J��(c�d쬴�Hvfw
�)W״��q ��Κ�;����� �zy�t�%�XIl��A��!�a&k�b�w�*�����ڊ�jd�4=8���gws����0�u퀠����깾�T��y��:/]oB���/a�.Y��0ߖ�����u^�2*�?]ωˎ �~n� ���hx� �@�IC	vu�������.�N� ������a��ur	��ih! �4t&��Os��e��3, �Wk{=wh��{:Q �r�V֘���۸��[���A����>�2�z���m��� Qa�H�4#	������:7��]M���І��pϡd���R��B[��?ρfۻa�o��@��u�a��uw�4��Z�_���CH�{ʹ���8��QQ1R8e{:���=5yj7*�JW��l�nkl ��M��Ź�3�k�[Y]�z�%L��L�%v����h����U��H��/���4Fz��#���m���M��ŇM��DL�!�`$.{�Y@�CB2v��""{v�4"��p�	 ��g�ge���Mn�Ũ�IV��&�К��X�&�vyk=x��:|s��ܓu�
[<�]\��L��%�َ�����U\'����*�%�Vd�(a.ξ��q$�V��\�]�z��>�}����g���� �F_7f�ͦ�ӱj���z/�y�h�m$:��i��=��-�g�\%A|ӌ�S? ��$%|�&>��f�SJ� ���G���L A�ݫ  x�Ο�u[S������wg�o[`�Ag�e��$�5��,H[�\;R��gwL/wc�.̞[��'���A� =�ݐ$�~`�۾���	x��!9TTLT�N^ɻ@|n�ML��I�^���Fz{Q&�v]�Fv���r��ժ��ֳ3��q~�>` ��W�D�:h��O%�߲�����8I&��H�+����s
�T������; A���{Ɨp��4Ve�i �63�n�����y%~7N�����XO�QnC&w��%~�}���j�Q'��[^͚+�%��~��I�n}`Giu�	ə]�w�s�<J�ނ�Ԁ���e�Y8���luFۈ���ɰ�q��*�O;�\�f�!�����Lv�v��ݠW�vl��+6�ͷ����mq�F�q�����oZ�D&�7&{��E��Z�tY�0f��-u��υ-�;<��,�<u��&��£6��x��WWv�;��|��|�q������:k���)�lU�뷶kĻC�^�9�S�n�q>Ѽ�ڒ�K�f�=ix�ۃ���;etdwcb�'jS¶~��M|d7
P�]~Y��w�K����K�>���ȅ�Gn�l @#c;���z	��iI@5-�y�3>��l��n��^��Z@$J��t�� =����\���x�W��nx��k�2�(ÆAvӷwtJ�'��d��\���r<�'I4|��/w��0&>��Nj
�*@������Ht�F�R��&�e�'BY��HI>��Syf'��$0�զ���2��5QDQUc.�ݙ���;�j�����WG *3��!��o��1 �.��v�W��z��w>q�@��[z�r�.r����m��Sõe6�gu�K�os8�p�8�Ҹ&�&�l1!��%ff_�D�����  .��qf���v���ݐ!{3���jկL���JL�w���G�T?����<����Qc}�gމ�H�����^�V��^>GD*��]r�k֛��:��Z͍�-)X��*��w��c6�a�i�u�w���;^մ|laX=���VF����4���//Uy(�S 9vj$�d�qz��f<����������@+�5i6�(ÆAw�\v��̯p^U����<���^��q�G�;�ӎ_ey����x�-�#�$޷�|Ek�D�e)G�l�l$NvX����U�@]���@|��ͦ��G�;��e?H��X�s�x,�Ҋ&	��%B��s�2]V�d��˻qmס"1\=��s�x�=������w�SUJ��9yۙ� ݛV���&�~� 唓h���|-�*��ff@�vm6^#ǐNQUJe
����v|I�'�//+�}��@}�v�5�D	��o�  �����ީ{����ܒ��ޘ�i�SP�g��+H$����BI�ג\�{(�5i���joH��w������{==uG�AT�_)��-���M��fN�i;
�^'w{_�^����
��n6j�f�> ���@G�/��H��Ų�p7E8��ޫ�:k.�<���C][�� �]�*��le��!�v�{�c���8�=�ʳv]����I�� �Q:vUL$�f�]�����^�yۻn" ���Ր|�۽��]]�����)�)��jBJ#����Q�:h�b9����� .T�Ye�y�.Ds���Iq�fz�C�"=z�v ��ݻٙ�V���D���c�Sa�z�}����$0A��Un���H���O\8�qs���5 �ї�M �w�0�#"G��w]n 0�<�*����T1�+6�!���<����i!�7�{<�ĒI��J��'������ZҜe�
.&�Z��.��B?k٘���^����n�����f`	 ��u8�ɲva�\��Vfe�[.�~�'J��M6b$�=-���֚����n��$��Re>/Os�*��UgJ��m��8�d��ۗ�:w��<F��U�H.�bl���QN+�ӯ=��H ���l�;�s��yqT� 7w{3 ;��m ��l`��K�ְ͕���s�p�sA�hD,l���X���ֹ��0�+���p8�pK�j�0ۻ�>���[���)e���U���C�n� Y����3�Q�"��h�%���H�V�R�`�}*��I5;�Ϳ� zOf�8�yseT{Y����6[����!RZ����z�/�}'�@UD������]3ӽ��TN��]��	 fl�o�D��!��V�;f_Հ���o'���π |��u�h �����ƻz���c�&�g����]�o�m@܅R�\�@�k��\$6߀�wfD`�6�_	 dg7P_ާ�r��2�9������Z�#�ϦA�y|\���3��Ф��5ʇҮ�:Q�=�K_75n;�Y9��NKg(]��#u
��K���n���3�Y�b�Ѿ��ɴ{�Q�-;& :�P�ܳ�lP���@.�ќ��3��������������r5��P+Wn'}}��Y]�U]Э�;��Vq���)b#4��P�$���J�nUF���U�y�����6��{���(���Cҵ=��m���$����~D��N:f�/�Wa��=���L,ۣ��Ƀ(�����9Ҍj�{f�� �z� %�6���2B��+Yoz��o��p�#H��s30���N�����eYΆ�;'J��	;���%n�)k�6p��g�%d"����
'5�2J���]�nԵӴ����u36�ۺٻa���現W�:$�=��w��
"��ï�+iX�yT���zn��b������&��E>�Ğ����f��m�^�� eh�I�9�\�??%�յ��/bO��=�:liy���M����f�%�o)�ڗDR��lDޭ�V��tA,��z����W�͐���*�$q��W��nP����s5=�h�w���qp�����6 �r;q��ݪǬ�'<�
+���ǹma���H4_P2솱�B�֭N%���N�-Z4��g�F��c%A��ΡVR�\��7y��`�mb�s�䘌Z��L�%h14�oJ�;��b���y)��*�[� 3�9'(��9�c�g9�ě���J��eEkjeaD�J"�(�T��b �e�UT"�YQ����b�R��IJءij[J1QQB֕�R�*��IR)Qb�+RTZ��Z2�[J�b�EJ�Uj��Զ�*DH�
��dXZX����Ye�V��am�
J��T6�ն��PR[d����R��VZ�"ԡQTU��E*QZֲU*�R�Y"Z������lkJ�U����E��U�h���Uj��%U�+YIb��+*��X(�XT��¥-
�E��!XVE��R�+H���b�Y-l�b¢�j�`,��@U�������Yj������+ Tm*J�
0X���AH)+*bȢ�Tm�
�hcǦ1�0OJt��v�O=�֓vy�#����GEc{V�M�;b6�uu.1�"��^sr�;�s�.�n	����.���x�=\t;�$p��U����{s�+ۭ8�oOkk��mֻ]���rBWn:����/�ey�<�=Y:�]���������7gX67���8qŮ��k�q��U����0WO]�x;A��p(f�n�y��g��;��7ƜY��`�ղ'5ڮ�uө{u]/����۴|�;�sGc8�n�\����ὐ��Ѻ�����\�ى��$�g�im�0]^��Og�q��I�f�tkb�)�'d:�s�gɐ�en]��50��A��'T��8Һ{$�W3<[֎r�t�9 ��1=r.Q=<�-��m�.x���g��i��<u[��J�o�����u׶:���9���nB����u`뭯V��S��s�Ķ{a�2�۞{Y�p�=Eu��4k���c�v��n��u���٫r�a��=��W����ݺ9���������]���,�p�>�>]��I7kv�t���v,b���u�8��!��g���b��kn��&5ݹ�B��n|����Q�^�-�g�wDj�lZ9���<!�a����kp%�=��Z��l�ph�o>v�9-��';�����7E���|F��۪��ڐg�ۣ�n�f��C��l������dH��磉����ě��iU�
���&��s�jLk�v5������l��uk��Fw5FW��a8ݽ�\��9\����y�������S�B�����K�4^N��mū���٢rr0\M�UX@�lf�n�s<{2��gY���<�m���t�N�[!ӷ���ۛ�ǥ��Y�v�L��BF�ny^���)Y���sj�p�:@:��]�ɳHDli;x�{3ɶ��r �vs�ӷ�=��s�k�������z��v�E��ۍ8kq�`��8޳��]�^q�$6�n��hc�K��>�n����Vš��X3���/;���8��݂�/m;��n8Ǳ
,��G`]�=fP�ճ ތ��&{�1��j���]��]�ŰW��OEc&ض������6ݫn�WN��Gg��vb8���n����A�M�<�U��\e�&楤,�q�l�>��^}�f��.����+ܻ%w��ָ���S��#��S�\�p�m�z0R��g���mt���v�x��������z�t]{a鬊�x(5 �3��ߋFF����q{�-�o��M�٨� 5L�%���ݻ�ؕۛ���f��5>�ƂfiM)(�l65���zrno��=XDD���`K�/��=��o��޴�����Շ��+ �lX9h�9b_����q
��u�)�����";U�����VEi�L��M*UPU1���5G{�ϊ�`�	��[�""�ku�v�vd_�o��[�`}�i�NUD�)�����?��=���}���{���m��~$0�դ��y'�E��r���������R4����75m҅�u[����b�
l �lm��������=14���ML��G�Λ����݁v�vf��A�˾��*��h" F�su�bH���S�&�����$��;�Y�����D&� �/�b �*ǝ(�!*fܼK̷t��;���v��t~�=�ÌA�&ڳ%��-��b3�긎�"3�� �owfb�w���ׇ>u�{a�5Q4P�������n�<� ����6FWVz�5 ��m� @%���{� "�����al2��j^l���u_tC��� �#�`|��wvf �{_f���Y�+# :���-$u�-DIJ�LL��1,y�m n�	��֧�� ��΢���� ��ͦ��C�h��W8��H�d�^�4d2�Ӯn�6�mM�9�j��&2"�z�DMH_w���H\�����4^�}t`A���`|��6�DO��Y�.��էE��d7���|ڍ=
f�M|M6���R�$�򯦾9;��t�D����l �>Ĩ�j�tn��ݸ��G����č�E�]�w�H$�K՛V� *�EO(:׳%^��ϓ��w<��Μ؏���TFh��,׉M4��$р��_7]6�c�6s��QoL/a��܇�q߄=o�ҹ-��}D�=��Ā=��Us��I�#RX��������~k��A���,�@ufۆ�͡Y�d<�G,/�?=�&�W��
�l3�j^l�o�K��]^��} y(��JF�tI�>��J����t8�Z2���}�źb�>"��L���KN����>lc���B�����b�X{\���Z�z	j#)�'�Y��D����J��| f�-/ETSk'}^���ɣ�۶��'	?���~�\K�	0�yNFsN�C'<C2.���V D��P;�XA�{���@�t}w;9|{Q�D�Ғ�52S�鿀����>7<�T��ވ��u;H��A{ʺٱ���##pG	8���$*,Y^J^{wI$��I�$�R�	 ��ݙ�\g���&:��IN|����zL�/dxB�z_L5�,GJ�'�3�Af�J��q!�y�Ǹ��^˟���B���DF(9���Q���F6���Ol6�f�D�B�UKa�cn��A���0uT�z7oDj��[� aͺ"#����"c�Z���*{���EA�8s(�&�wn{^:�y�WC[v�Hn�<s����\m\l�E`�e�"j�/=N!��[N�o��2"��z7[�*|�W��H�sˮ�D��X��IJ
U0M8�|������=Qν�f�U�	 ���� �����U�gRڳlVSޜN��6�@ӊ$Lͤ��?� |��<�  �=�`�R��� �m�������F�p8�	�Ի��]{��J��rI'��N� wwf` #�6�[����1��'⫻-W�)�8I�m"��3 <�j�<��^�w�k(ۯS��1�\�r� f�vf|���+>��>�'z����[v��ݵ�=�߹�vJ���9޷Ym��3���i��;�ߤ���k*m�n �\4�'$8��X&�'=�%u}�@�jl��۹7W�v���y�k�v��ctqή����ԑ��lV9�x��M�X:1�l�b����n���VRr�܆r�㛶�;�{Lt��,�e��iÞ�n(]I�u�H141/1�k�]�\ۢ��n�"m�*ݬm�]�7.���Ԁ�|c�vݖ,�{r���n�����x����&�B��3�T�������ghH0'b��vҼv�g��3����������ֺ��}��۟I!��	n+��.$�[��� ��8�co��z��ћ~TA���٘�J.bsD�f��/�W��	.�;}<jf�ݎ��govf����D4e�g_���G~;6�Rbrͫ��zςDyK��&�$�cڧz�zx�����#����i{c)����(��	[���p-�D�}o�	o�M��&�1���2�y�5tt�_��n�U� =���{䯙�<ӂF�n�X����| md��9�7���o�n��� �y:ڒ ����#��8�TW��TR��Ρp����{nx��F�BI�ʃǷ���(3�2GgsД�����==w�` ��ͫ` eg[��U*��U���t�m�����M_���7�� X��;6�}h����t�~=�ewS`���}eo�1�p,�:Wsd�3G��F�מ�D�V��ʽ��i�\ë��r9��()z?Y��Mo׌=ɻ��>��<�p�+:�>P���ۿ8���4Wb��N�)j��{$ &zbD�h���'��N�����y�m ��]�qF��'*"A�	�7��w�����=��|%�u[  :��᠈�ovf��;���wqO+ ���rzBI�A%TPƁ��6 �{���y޸7x+�]T@�{m���:�M� ��ݙ��<t�e5�C!L@D�"$��ye�;K�ɶ�`�����R��ۑm~�����,��fQ�K��$>H���ZA$���6�	}�=|]��{6Q �h�l�'���$��C	�Xmw�d�VR���}ux�6�n��ݙ�DЀq�Y;�M4��;�$�E�	�
�hD��m7:�r �����y�=��~�[o�}o����e�wrP ��Ҍ��C��
��P���E)���SvTX��^�b.��H��%Ud���O�MD�EB�+�+vT��{��|��.�~T��I�_��$$�b�,�u���> ��T
5�����	T�Dӆ�����AϽV�@����
d�Խs������G�����}�ժ��ͻ����hq�ě�i	�z�v��lu�R�o]k7�4������+IFB�Mj�Ǜu�{�` ��[�V=�EfQ��ڢ���$Ϫ!�52I-�̳�u+>I|߻�����%�H� �[�`#-��A h[�{6&y/-�f����yO1�ȣ�XN:�[^mI�b}��� �7�pٹ���6���{�3���<ڶ�����"GLH��Km^�}]��EY�U� s�i�'�My>� �t�H)��Y�I�j"'��YK�ʡ��.܇)�;�i�?2��$�~�aVK4ǆ�U�pV�zl�<<��bw�9�����ћ�ۺ4z�5�m�Z<��TT]�߶�C =�����,�ET�4W�o ��y��@��Ywq�o)&�>D⑦[ �km㊅�)�*�ą�䧱��#�5۔7)�>�O쿶��S(������q��:��>@ ���!�/˺(�)�l�I1?b_ �u��U$�1����t A���\��R���=K ��m� �yۢ ʛ�=�������״�`����S*�)���C 7O;������;,;��ge[� �ͦ�Gܲ����EF�q݅S{�s�&�7| ��m � Λ� ����,��2�M���	�t�O�CqD**�����^�@ww<f�X};+ݽ���l� ��V ���l�q��!�+�k��C�E�Y32���lTQd�fi�]�= 3�t�� |���G'���8�MGs/N[��KzSH(���Y�C�B^MZC�<�wq�u��b�{`(��L���v���6��vW�^Dy32WK�v���rb��j�F[�U
n\���nc[�cF+�]^|��vy�wU�m�η=�s�l-�[����֡-�1b��gv�g���tq�;�ɖ�`ñ�&�tn�� �=�ns\�ƶy-�g��q��G;k[�x� ��ԗa�M�/\q�y����Kx\��hָ��PS�7r@��g.�����խ�DpX�D,�}��\�ceH�U_�U~�v� ۟7"�7w�3'd��NN�M�ڭ��t�@�G��̆�X�3�PJ�2������ �H�b�����~��  @,�י÷{�ρ�ߙj��d�֬	2�
PEp������O�{{�}�@��k��~�u/�����#:��D4�����I]-.*7�(ą��*�C��¯�P���Ȑ����A��]�2��l���~>�q*���]J�)6XJni�߭�R�z���U1�Z�//) ��V1��������J&<����|ia�tQ"NH�d�s�Ϣ�����8�r[�±�2�:�����ߦ��P�bjo�)ο�� ���`|�&�~�85ӹy~��-�� �����HXRT�`aȑWFVt�p%�ق<y�׼nv���������ԛG�ٻ7ZM���f��N���<Zko� �r�jl�R��U��1⮺m��P�dFb��4��k׹>�� ��Ϳ� �c~ĉ l��4U��[����37�߼����7�L)�	�6v{���Iw�%XH�W=�?S�f瓘�@/wwf`DG��V�<ڂe�8@Æ�O^�[կ=�z$�D�&<K �77���3��՛��B��0x��켻�	*ۤx��f4�g��V�'v�X�b��ܐ<�B��s1 ��6� ����T�^�t��/a$!�$���&7����nI�59z��v�2Đ�d�@K@$L߷�a���	��n�g��ٝV��~܈�%�l}��5'��$$�O�*%|�E�a�DR�q݄����A/s:0j{~L=��$�k�O�D�h��˶�KS�k�#�����Q⒤�P�����=Gz��Iy�nA��Ռ�䩗��cwr
��t��#��ĺ2�d��a�=Oz�O�\�5z���q;��|����[�w(�+�7r�"�n�Wl���X���1.�)��j�#�釶��q���޽'&v��a���(�t�ލѮ������z<@��lJ�)3�*�>ͧ����SFs�"�C�z�(۴�\k�\t5�����@lҭ��|/u��N䘩��MQt��aS�n�4+`��&���C�:��3�*��q%̒�j��{ҭ��LUդn���ve���k8����_��{���v��=�:cB;��x��4�>�G7X�n;¬Z���i�Q�K��6�fwx�w^�{u��p�	շ�)��c�&����;N)�_cir����/���C�������1�хy�{��E3�"�uc9�ݵqw��_>�� u-�~7&䝋.9�Ƕ�w,ּ˛���Ʀ�æKf-��y�:6w��6���Y��0��n����)JC�iV@�*�l��=%����iܳ�~���;և@$�=ӟ1n�2�vL���ܩ���}j�w�{֝�7�栫���}�ŏ�
6�ϯc�{DB��}�	�m���kd�<G_mIu���|�n�Ҝ�ݑ4���U���/�p���,EX5�jiyn`�J��\r�i��\Y�Qq��4
,۸��/+9�&Dv���a�T��#g��0�ʝ�tɩ����O:�1�׎*|�{�W��N|1w�}���{�k|7���"��e
"��-�J�E)idH"��j�E m�-�-�*�Z�D��
�Z�B�V%maUFڍe%T�(�A`�*յ�B�mA�
�P�*kTUҵ��ڥU�إ[E���aD[klQe�TDb�e��21�QJ�j�k�U�������`���T�J6¥e4��Y(������l���PX�J�b"
��b��(X��ڔ�ږ�F,�Em(%h�ŔE�iT�j1jV�V�ԭkmBЭJ�����P���(����k���B��ʍ�6�mX�X���DF�TmZ���UJ���@��R�(�����%h�EE,Q����m�%��F"��AD�m���bT-�Ph�V+ee�k*��֔��Iz� D�5 ?Qx}�G[" �����k���W��-v0|'��d�~�TH ���Q ���m��vϳO]�A:ݗa+�2�	Q�n*L/o�@D{w��5�1p�('���Gy� @-��fb�#�$I���y6�uέ�q��\�n��'B6��jl;��mҘ���A�F�`���(�PFRX3�FMx�$�=��X ��$�}}Yu5fovr��I��b컉c���Jf��MSh{}��T/9�6GG?:=N���@}�>󘈎����S�q�<�t�����FÈ�������N� v�sŁ�۱��ݫ�w\^fF� G���� ������)*i�0�[�uaKΗ����DuAc�z�cN� ;��3 @y�ԑ${���#���l��GnۤFՓ�۸�����l2d��Э�dpz�;m嫞K��5[���.V>�Uǔx�vS*����ko��P�T�Q4�nvvg�D<긏(����8��p`�Κ wwfb�=�t�Ihm�}w`��a�i���;^�J �����j'k֍�Y�8�\=]v���Kl�!QƼ���]�/�';{��ɢ@1�j
��yG�u�T`�I}�D	w��3��,���)S��u~H�6x�P�ҫ$��7b@ ?N��ۢI&�5�J�$�gA��%#�o��о�(^X8��TWyF�?G��[@ W�Q�!{W�}�h�ٽ�d�$����$�G��a!�>l����Y���q�����`@��v� �^Ԡ�뙲��oҐ �ݶ�~��	��i���p{�����$���Zo���x$�MV�8�$�A��o���+9����&}oK��Z�3^�e��Ug]y����޹����=
�5qxyI��+�>�f׏:\�5lj�q,��-^j�v`^��N�iл���<����t��p�ln�+r�v�����m��8kq��]�u�0�nx�{�Mے�x��m����u��NOt�ur:�^Ln���1����m�����}����\�]]�q�U;v�u��u�|��Ar�xj�������{^q�n�݋d�b��gH�(����X�8���p>�֭۬�=��9n۶6�̡�q�'^�Gd�/[�:��;�����l��ӞE��n��Bd& lG5�]f_$����� Y��K���F�te�t�߻�'�$��{��[�4��j����a���gI�������H��fۆ� YYͲ ��ٜ����zy�^n ;8(RR* (�6���qEv>� �YXa��~s��bTL!e>���)��QJ
��D�6������}:�2Q� w�V�" ���� }��ٝw���I�W�o�m V�ل��!���F��}v�A.��}��Pw5�19Ry^�[���z���a$;w��'��̬W.�
�N��([]�[�]�u����z�c:��4�xǲ�쓸K2}��zE��U8,�d�$�Iz��ς [�ݙ�:���6�r[�nZ�$}�M���[O����8��M7Y��=���3���Xͅ�35�P��yHʎ�흡<n����t��;K�;/���D�)Ka���̒nw(��o�ƌ^y��������$�
6��i owfbת.1Y�eWmM���l3���(�V��z�� ���sİ A�zB���F��޸� [Oͦ@�	n�vdE߫�T))
�QH���ܧyOe�}�y�� �ݙ� ��?mF�'�ԟ�{��m$��wig���F�P��&�������  �����*�P^T�<�=�^w~A%������U��pշ��_YP�I��(7�2ҡݮ`�N�\�qg9��R��H�a����R��Ad{�ѨHnB�:$ez���D��u�Ȕ��u\0{�mսf$,��� �{{��I��$y�mc-�^��= R�(����EI� �;��` �+���$��Ʀ�	��E���i=
��L"j$�U.Y�ϳ0��:�!�E�ң���z�G/馦��|F�:�ԥE�g
�6�Xt�Ŭ{c/��i���/���Y�1*��Zی���+E�kq�`2;������3�{	�w7���M��ԦeLb"�⦤r�+�캶
�UW�~�7 v>� "E<~ѯ+�uw��8węɷ���YB���AE!�unS�h�����iU��S�<��p6FۢI&�fu6�����(��5�6�3�|�r��8��	YHA��0�7Ra�:��X���ۄ� H8�d2E�}�L�J��^�I <Lo٠"I&�{刕�7ܽ�!�n-QF�����^ΧK,�w�b,��O��݀u�וN�{1��Hf�?ac� ���� qκ$�%G�~%�
2�JK���V��F_7b��X��������D��q�̾m&�A��0������]��P/t��]�a,��V� �?^��`-��̎��7)�%yԿv�%��⬮r����%w�m����-k��������4�c׼�}Xm��_��)���y������z�J��m�|�3�j�!Ov�H%�ݯ0�n�gذ�쭈j�;p� '��Z$������VϸX;e��I@aZn{uFYأ8z�m�1�ٴ[Y�u�^�cg1����w�QP��"�RR��չM�����I&���6�7��@N�x��y|�L>�Pg}S*
�
S5N/z���@���X�L�����>�޻tH�=�m�I��7zĘ�I3��5�W��B����/vc�� ���b�[޼�=w��O/[L����s0
�E�z�PQSB�:h���X�I� ����� g��3 �:���r)�?TD?�f6رP�XL� m�;�o����$��t�	me�npXq߱�Y �k{���K��I�"u�S }����y�Ź����Jcy��u��.���c!�V/o�ng�_;f�$i|G-3�ѹ2�	�����.,�Pv�C�}����O-�kM��%�Ϙ(�d�l6�p�;sv�����r��Ҝ	o.��<t�t���RW�wFك�<Ojӻ���u�v���Y�ۤ����z�l����tB�u==	��WN�z.x7)�z����>x-���nG=��l�����llK��y����u�pV ��ٶ��*�k���z��M�mV雋�`8ݵj����E��axwVٹ��%��s]r����i�*���a���5���3�ƽf��x���v����r�d�ڪ�f!� wv� ����e�q>����oci�|�����~�*������չM��n#�����u�$��Ғ4I�����l ��'����Z=?:�d����4��bJD�[s��""=��� �d�>��3���w<��4���{s0 ���4x�O�������t{:�Y;]�v ���%������	���nfa�w�[$���;�%���aJ)4*E׊�m6�	����o�=0D牒Pv�sx� ;ӈ� �_6�u��n*a�NJG��B�(� h���uӮ܋V,��� m�:� ���=�����~�aH�*�g�e��0 �}V�@ !�����"���(��5۹�� >7Sh�ْQSR�EUH�u�v�Z ��1�n���(Z̱pzr0��Q��N[�T��+���Y�QT�AQ/\�}��u;�Wcen���O��j+EnfTׄ�����/��6.����p�@|'�ͦDF��g��������&�yL�p�jZM�8��@��ݴ�r��ٕL�{�{���c�o��'�������F\8�½����CG�Ѿ�� wz��_;i ��w{s<���&�ۛM�����u
�&��T��{sɱ ���[�7�W�2�o�တOo���{s3䏯&�8�^:�ش4G����8 v��+ʞx�9^LQ�z�%/X�,��s����)�̀�S*.��ͦ��" O׭6 [�ۙi)�|��{`�V9�A B�_[L>��h��"d��nߛL>�{�,��h���>�C��m ������ E�:g8z�7�=���i30FT���UH�Syͱ �����~%�1�P~2���G��y���Y=R��.5b���tw)kv�[�.W���z��O;,q�og�1YY�(3��4�S[E��)&Ap�\z �iM�D�I}�����HV^ۅL�@�P;gV�8=
"n�0��}�������l�Oğ���6 �;�S+��sL O���6=p�Ąd��'�W7��yN��b�.�i|��Sz�!�� �[�ۙ�Ds��)*�ܭ����b���8Ϫ(�4��2Q�b��p<��3�(.n�v.��ˌ��������xk8�����m�Dv�k� �'�a��l�=�g?g`��[dDf�ky��U��8�Nc�yo� i|�z_��{wZ�S|�z�5D���sn� ��w�h��a���It*�GA�V5`����P壟=��@|��'�� �S̛w��o8L�z$ק�ͲI#�ߵ"F��"��_6��Sc���Vd��o��-̮c@|�y|����j��>k�TM�������ce��-@����.�10�Ǘ��x�s��59[K�/����FpqݧS	4�]�<��P`��3���J��]��Hp���^���}��3�72vڒ >By|��;��48߃g��"(����!Ĝf����]��8����z������j>}c���M�V��{{��  �d��  P���@:F��߽�����ߵY>�dX3��,���!�����Kg_�wɉY^��ٕ� ���2 �����U��{��P��HI	1�S����� :�4���.2�MN���@ �̞mI 	�slؠ4�PQ@�r*v���¯>�H�)���Y$��HY�|H�����٢Xp�|����!����2�����G- �k۠*&wz&ʻfc��"�~����|'Y��� v�y���]~�+}����C+p�H���%V�|�E�&V�������G缝�|;#ם��_s�=e�7R�R엶-���>��>�9'm~q���d�������Q�].�p�%�%v���j*���[n��l���9KR�Wˣ�pyWK{#b��e΂��P�/n��[3|�o�9 �x�=������u��"����u�H{��dniw�f}~��b�	���В��w�=�q�qθ��zoSiP_r��%���j�w{~��۞���VCx���/s9���'��I�z�7*e�:�d�9���:"��f�ܥ�b�r��]�!����sA&�Gi�q�����Y�=C�-�n
ӊIK)����U��Q��c�6*�_�*K3헧nu륩[�Z��2I��7�f�>��^���Z lغ��!{|o,�4���'S���Lr�ۆ�fU��Ş��\��X�8���e)17ݛ����x0	�Q�kNYu\����(�:KsN�n'�ו�L<P�qa�����3V%`H�_6�v���mڻv�=i��2�*c5bub�IQm�e�Y�kh�!OfA���0��y���CʒP~��!���N|����Z̼.Ν�[��V����y���-!��*Z�,�<��8�.
�E�[��t�Li�O���κ�K#�e
�Wj��&�5 �/s%TD�k�X��Z����� �h;���������cKꙻ��NjW:�
 ���ѵj�B��P��b-�*(V�Œ�Q�E(��aET�,�-�� ��Q���4mhʋX��A�Em��QA�R�-m�ƥ�J�m�����[mYQ`��Q`�"$b�iQ�V+6��-AdE[eV[Z�J�Ҩ��*�T� �(�ƭ���*QV�eeE�#b%J�F"�hVJ��h�Q��ثm[J�J��QKJ
�D�iZ�J!b��(��KJ(*��ƥ�Ԫ,�ň�*��*�Ԫ�ڥQEUV�+b�QQ��`��*�Z�Q�%e+F�b(�� ��,Q�ڋ+R��TAUQDKj-J��Z"��R�Պj��*����֌���������J6�b�2�H�U�{�w=����j��z��.T�3[��N�s�����[����'�н�^W;o\��śs��6͊����R�৞z.+v�拞�XX�S��c��'X]���7��;zϖ�J�뮶ۜ�xMٮ�m��e�0ƶ��P�N��m��n^ֱ�6��,��q�2�q��Ӈ��iq��d^��9簐�s�C���S�;�/=�s�p��cv���{v�	[���g,[����v�ϵ��+m�X�[�Gk�@�88�v�ڻZ�bgb���,<k�������Vu�X܍���E��;7"���ɼ��V��9�g�^4���퓄�W;��m�M:���gm���sX';t`읩ze.ηj눵.wk{{=����˻B�7)�Z�OnJ)��Z��q�Z�»;B�Ӯ��m���8(V��W��㷭��qě\��;��;xn4�!�x�
���/k���t�Ց�G���V��M��'pn�ۢ�v��ז�l+��;�x"�E�=M���a�e�{6�F-fPâ�[�,gxI���u7<V�2q�&4)�Lp�kP�g�b�r�X�mn��/d��n�Z�rϢ�#���ۂ�%��\Z�:"��y�<�zcn$�/�i��nZݵȽ�wN�r�';�;���L�)MF��{0>Ɏ�n6-F{WQ��-��dx�rm	�t�lOad�˳rh��s�4��mۜ5�@���G;;Cg�y|;73y&S���Wm�y9Dǌ�8Ѻ�ܳ�g�u�;O�G���h�r��,3��9�ƱyE�[v��vz6y^���pT\	���]�,r�X�g��c���]��fi:�m���M0�ß)�*:g=���� ������/Gqu�������8�1�{q�g�	���wh�v�Iî��9��9��qZ�n�6xT�Ƈrs��(��p�ktݘ��r������Ûpq�i0�#=��="��;';X�tG	�#�a.s�[lysu/�湺�� ��v�Ŵ�=Wn9��5;�K�O\s R����kID��l�y�$�.W�c[���]����j�n-͍�o]�n���wH����̞w�Vo0n�5���3݇��]eK`���^5���-�Z8ݱ�nZ�jg��$�*�ٮC�.���lP�ƞ����jet��n��ѽ����p���^���Y�kլbs۪�[�j�w�����O&y�>�wa9h���s�q'w7\H�F���,��v��$�_͟ ���f�p�o=�߉�-�$:�o�e�:=2�QUF��"�|�d�4m��]�����Ss7��HtH,�-|I���F����3��t�d~�|�޴��g��YQ�d�_?6 v�y�	ݲŽ���x���B�uشI]����]P6�3p�*?�~�u�n�q�/{x� �)���4H��z6�7~G��p�o�?DE��m�RA����j)���73 vd��Q^=p�q^H�>v����f >��� �ɝ���ϟAN�Q�>0%IO�&&�$�i�m� {o]nLӭ�ru�];W=��O������������ϟ͈�ݽ� fW2�$�q7wj3�i��H�D�Oz7�|����"�������o�<�3y]S��:�]�oӷ2��>�|^��wJv�>�h�h�ySl;~�����dH��/K�T�QT�ˡH3,U�@=�KGJ����$��{����fO7��M���[�~�_9��^��n����,e�H��6�_$�Yx���%�s�{�vy�D�w{٘�<�}�5Q_L�AMKh��(�_tgC��D���O�M~$�3�Q"�?l���rN����i�]�mߒU�~�؉�7,)x���H�s:�p�p�����b"��gfDb~�o� @|'YͲu����˺�{Ω�`�K&0ː���:����7U��g%��3�LN^��iz�<d���}�����j+f+<�� ����� 'Y�mEl������o?{3 @#�]��>�����O��[��~���\���;��t;���L�@?r�ȢD		�s���b�E��T)s�{�@}��sA"���M*l�m�|�v��I$��i4-Ă�Im����s�֍ȫ�n�7��x�ױvO;ib��e��[�D�W7�!0v�y{P�����{9r>�1������pD�g�y �����䈃�'Yͦֻ�a��NqYڝw��痽���a��=� C�y� 3���KǗ�Xi�+��XW�;�/u�J�02�A5-�^��ؐ���Ņǻ/�iy{�״oW1���o6� ���x%]�����(�/��L�>0�\Nu�m���n�l�c^q�R;���3r�������~چ6$�&NR���$�3n�$�F�{ѷD����Ը���a�_��	!:����(�(������z��^�-Ը���nz�}!� }���������@�a[j�;zk5J�E7�3>�I�$�l]�����q�'�����{s�@ ��޶� ���{�%�ܹ*����avӻ�#W{r�db�9���� {���πՏ�'��s���|��a�R����&�u�6X!�Z�f=�k�hʟm�\,ܿ;�>z�e����\��^�j=E�V�r!en6�k6m
@&�����9��� _����iu��"3�f;` ��ۙ� ��>���"oO��^��ih��b)p�֊��2����`x�e�. Yg�R�J�E,�s�K����U57�5���{^` ��s"M�o/As��u�� �ݾ��Qu7�`��10�XR���H 鷹q�|�yl�6 >�{s3��#�'�� \���U.�>a�0zSP"JR���1�}�V�ד��D�/w��zfS�ϻQ$���<ۢI)t�붇��������T� �ܛ���N��( ޽��"#>�η���4�]w}KV�	�ٙ� ��΢�AQ��vU�$�El�k�)��ꋕ4��;������m !<�m3#H�¿cb��,���	6�M�Z���U9��f��u�P���R��g(bt�5	����u��{^^�靲��\1P�(�׽b�/U��b������e��ǟK,��NZ�⒆��z��˴�r].��IE����鹻J92Gn�kUk��ȍ�͏8�;lg�X���b�qqWd;��q�W���n����%v��V�h곯�ϕ��9c�:�O�[��m!��
�v�Me�jL�;/�*�q5�t��:��sj�E���im<�z�˳�ٻv/�X�M��ѳ$ۭ�i7��n�V�̹ #'/`6h�M��p[lM�*��'�n�^��mߟ�����F��xxci/�2&c�h *$��-UD��M�ܺѹF�o��tI$�c�@*� ���L��D�MK`��`^�k癢ڽ����A-��p� HO/�dVh��V�{�g��g�<��A�#%��������`	l(�/�)b�z_g��z��q�O/��@���'�j��Ϟ�yOV{��gĚ'�y� ��A=�@D���<�<7���$���i#��SxPs����� Sy�7�{�,"-^���s�� �����	���@��o�WH+"<�E(��3���ţ��Y�n{hMq�պ
F9�rM������\@T���\g���9�+���b 3�ݙ�#����S�0�z鰈�
�����/ǝ�!L���gk���H�٧^�*���݉��f�Ċ���m�����֑�s�2?!��,z�'Jy�%�tﲒd��m��<�F��e^^��kswW�A�������$�����lڰ�-�!`��)�(���L�O$ uD�9��8��w����A
�}m&@��o �NT�f7�FU��]gK���{�k��;6~ �Ɠg�.�{�1 ����S���� �Hi�_�i���	)J&������ DO{��A��7��ʍђQ&�I�j��D���~I�}�,����ll���q�ܛ�Xx���b��{�T��ۄ�ό��hw�q�ar����$\�}�Q!K��W�wt�A�~$��{PTK�{��'{sl�c ��7�g�]E �@R�M)o�:�6�&�1Oھ��͈"��f`�����;�Λ��s7��洚���A�pՅ��{��A"rgKh ��,�۷��%����z��. .�lurV9,�*�ֶJ�x ;u�ࣴ�N�u38
��ͥ6V{'u%�x��ϭ�K۠�����OL�vC�ͫ��1�Rqݤ2��R0q�|��� u{��A!:�it�/�\W�����Ū$����N1$�+����F�I��[^̗.bjy�S��<���^�dC�:�o�a*�׽�.<"j�jj8�":�.�:[��:���c�7��^����	�����
E5�5���{Ȕ�L}V> y|�{X:�K�OTY}�w�� �GW�[�Q�A+�5�}RP��+�D�����ou��W�_�R�4H�W���	�;2��w�'Ӽ�U�C�=j���
R*���rې@ O��l@Anob�7+v}]�_�� :�=mI�	��i3ב�dEI*^E14������;���<�@�U� %��i ogfn��h��+e�é�i�]����쉯p3����J�39s�#���ק+���~��;�s0��$��ut-��pN�5�s�\�[p��$�f����=�n�LFь��Զ�y�4؀H=��x�D�U�k�n�2ԘI��DQ 4��H��??x$ܞ@�ɰ��"�e$QA�{=��'s�A���� m��Ǵ3ۧ�l/F�����?�^n������K��� �m6 �;���{*K�﮴(K�ud��-T�{�J	)J���Yw��Ł�yͿve9
�v��H�I����?$�O��(�<[>����s���n���J,`����7�9����[��n��W�9� !fkw�wgf`gi[DIJ��"������h�<v3�����+�c���3�9�@$�����V�Ij6�.���a�[�� �J�P�;�31, ���rvzв��D��\֢@4矛�h�K����s���'��8��ލ��^�/0v+w�#eֹjC�xVV�y�O2�{˛��x�(��sՆ��!R��N��1o{�qVy���<j�)�	�u�o��FZ�'G%��^��M�y2k)�׶�ͻV3�r�^q�̍�m-�4�y�&����'÷h��V�������{M=��ιՎ �)m�hG��y�F.l��![V��u=r�>X��gt�F����M�{mam���;5>��iw$���6�g�:���s5�7^�|�-Q��,��W�:�N�]�C���wd��@�NY���m\E��n�0��2[Je�����.n�0���`�J���5�$+s�>�I"d��l�� �L�Q;2��y�p��_P�f�d��f`
N�Q1Jb��ҸUc�ƐK"��?�m|D�̶ ����A^��������q���^���+I����P0�R����c�@W����XFGY�c�Vקv�4��٘ ���rG��<L����R�
{�������ESx�  :�Zƀ@!>�>�j:�=8�6"!��癘�����
T1"��m�܀ ��Zomӿ��3Py�y�@ �N����_�L}^�A�9o�籿��<�:�
]��Xh���rl\]��/<����B�)�>'A0�f�ffff�E�AYua�a�y�yms�f| ���HV�7A**`)LA5��z�w�A�K�4�-������R��L�����,X�*A����w����}��ȳ���3�G5vl=x�3��Fb^m�֟r�D䣉�F���Հ kլ` '��� ��[K���g�~I|�+`���qT���/����'��`W�����]p�����ӭ�	��lF���E5�-ڪ��<}�m��W���R $<��>;��1��K��[���J��>6������M���M� ���ag6�#�Z�l{�{�^�l` �sw�����%<3���/�{�ڏp�I`�Bp�".z^�H&��ζ�v�);���\vs�;��zY�m�m���g�6�BB��fS���%$/:�&�A����A�髚7P�2\�Ϥ��	��p�^���P"T)&��k��� �4̴_������ߔ�	��h wgf`De��wnj�;z#���"q��u��h�� �7I��Y �d��t�$��~̘s���`�)�soR5Ԙ�Z��n����uo�{��9��
䂄�әlqɣ�ܬAڝ �y+EXs������h ����=h�����|嗮��&V&̧Y��t��&������]�w}pF�_HِTt��<���3ʰ^�2��YGvm˖6��/'���fB\)�p��>�L����:��c� ��މ�	�j��%.P]�4���յ�m��>sg8y�m�֣�wG�vPkqҨe� �-�����Z�y��Z��lK7@�p��AiIl�������/Z<��9y�qM��L���";nwI�:�<"�|+*-�J�&����y;����7�o���Q�+�2�����+��h�.0�-�#r�-����6��{FJ�s�J�=$�;T�g����"��硿��mH�d�:�{G �����lz	��l���B��1YAA3;4��B�n��#�2�K�d�����7�~r��)F����/z9��_Xցe����ǒW���	`ᏦӰ�f�m&��$��>�y����(��WvE���7W���6E��ʣV����y3ɑ�<�|->Ѱޘ�Qt�� 4(-Qo�*d���fJ��1���Zq�I�����\Ui4Hu����/�V[t�X�#�c��Ԭ�%���5&;�f�]uWT�Z8�I����w2e�����᳜�P,im��3w&���:d�h�JH3l8l>�&�4�^��{�L� �.�~����M:v&ƹ�K����¯Fk���J���������UJъm���h�-j#V#T*҈%eUV"��2�* �ڬX�h�U��l���F�E+X�����*�D�jF�ڈ�V)Qb�*1U�YKh�+m
�mE��((ŶUTV6�eQ�iQb��Ŷ�(T��RZ(!QhԣmEF��%J"�F"ֱD��Pm��mAE*�"-�Ʊ���V �[*DQAEk,X�AUTb[DH�cYZ �UPDQZ�AQ�)*6��e��UP�*("�QQPQ�**�*�**�Z���""�U-����QF(��-�APVЬDQ��1���V��"Tb��� �0UԌE���-�(Ѣ�eAEAh�b"�W�g>��H=��̀��f`	IØ�p�Rҹa;Ƿ���+u������
ߝ�� >[���ϐ ^�e��5���_!����3.���P6\q�E���0 �:�=nM��lۂ�E*"/��� K}���@ �N�!1_9۔����-� T��ɲ��&I��k���n5��/�3U7]Hn��Flm��_��w�D�eTT��
o�����a���0{���Q�DQ4jf��"L���tI���ZSPF�mC����6�h̿Y�)^����؀/v��0"�Ӭ�a�)��5T,]:��,�h�ZA��uI�o<�ϖ =^��$@�~�+[�o��#� ��ݙ� �_^�o��x�Ę1�D��C7��Ǳ1�X�~�}��` ��z���> O9��O=�A<tm:b`X�K	�4:$�ʚT4w&{re[��4nTu-�uu��P����A�g8���-�( �ػٮ�̭65�{)�����Ֆ�m�<�m�f$�a�CUB*��A~��) '�o�߶�����@}���Ȉ�6�<ڒByʹ���Z{VS������x�c�>����b;�.��W��yWƜ��Ae($,&�>�<��M@�q�|��9��?~�}��� �!z%�r��u�W����TO���� ���/��n�ǉ��̎�!tʬ	D.�;kN��;u� uzz�	��i���O������I{�SԌ�&�n��L��V@4M)�$�%j������޾��>6�<ܐ ����?+�ه2A��8޼l��#�9n�k��=o� '�wmFwg7�z�f�}9i���7>nAVt73T� ���+�c�� �{��y�<���\�}0��ש�!�g6�gwg�����/*�l3\e��Ӑ�k{�y�i ����r�rx;�D�\�٬[�=�g�7�_$���Gt�����i�ۭ�nw� Om�ڍ6���$[���^�Pɗ5�����UAͅ����m�8����y�9�c6�&-����M�&����3���`��G0w�96��W; ��&���Q�n�1O��5v� ���zCv�ֻM���n8��Sl��_G�[Z�E^�B�w�y�
�%�Ԯ8����+��ҕ���c��S0�\u���$-�kw!�n�x�f����b�9��e�5*v'r)�tF�2���V����ŭf�Nҩ�;Ǘa�H%\�n�M_{Ѱ,Ia���%F]�\~�h����ش�7Ɩ@�)�8�Ϸ1`�?J��W����n������ ��?w��jǳS{yw�\�qQܴ�J�� n�y�� fF��������8"-��� ����2#>�[s
����N&���vj�L�B0B<�?0�Hn�?� .���� H���^�z���Y�Dg�jŤ<!�f���!�.�]]~��� ��vڑ{b^��uo{���l��fb�~�mI����7����oϼc���U+q;�k6��n^.tm�N>��a@���J��#�~>���(�#H����W�[b���cϰ�>��k X5Ow�j�����"	'���d�i��c��D�Zw�n�D��y1���x<�k>ܸ�&�l�����7�ʷZ�ԄaXB��۾[���ՕC�˳m[��E�tH7x��o�h^߹6|��7� ����:I�ڬw7s&�y:
���/��k`i�	��f�m��"z��_��W�_/k��&s}g�o�����@|����J����*2T�`�9ؽn�eLl.������7� ���� R�E���Y���.e����'D�r�l�N�mH�v{c��A$���`]��
[;Y>_�ݙ��N���$�B�eݮ�W���;ٸ��)O�q��d�^y�>�ܮ^��m���񹭑�mq�w׿�4��Q2�AMR�����A���� >(u�v�=��/!][�e���� �+Z/:�4#N#H�=+j����U_����� m�vȆ���z-���,j?8�8;Oβ��@��P]?�/�̇�	u���X�)��qG<����-W۸���m<$j�%�����'��m�Ԋ��ۋ��qPc���yjl8�H9�]��SޞZ�Q��U�I&�z%���3M����p&$r�]�RzDc�۔zF �[��!�:�� ;�i6黮�84��#��Ud��n�*2T�`�9��b�v<�h�jf�#գ� ��k���t�$��{Ͱ
��ܩ�tpa�s����kI�U���t�lt�v�V/Xͳ�l%��8f��gR���jFۮn���H$�'^�����
���ؓ"s)#��mI�|'Y���9ȅ�D�jS�֣'�A��]��u�1���ʲ~ �P�|�!��{�3"��������"w,VEI4E) �������v�<�H"=�ׯj.y��J u���=��B�u ��bĂD����o�C0]o�'�׻�	 ��������2w
y��߭��}ouml��lY	�wti�W��3Kp�۹խ\�D��\��Ty�2��*�j8]��^ر;�u*�:#��U�w)�H$�I�$u:�.�?�=����J��4��>���H���IU*����~��=����i8]\I��+��%�T�v�zqU���c��&�~����f:9	��O2�Y#���������3���g�xG��$�Uw�� >�*�2�,��q���c�DឱC�>YƵg��Y ���ud��)�������,�]��Z	��Q(2Qf;�����Iy紁�ү.��cں��v�ՂA%�B�9,�B�I)��\��ޣ�U�~y� v�b�w83�&��	��۰K�Sc�& 2F��}��	��_/RO�Q���֒�*��_;���l�2Irrř��ۗ�#�Y@�����w�LJ�҆J!�5��KV��r�{Y�u|��q ��w��fRm�,�{b���/o�>*�ܞ�(w�#E��l�M#��~M<Nn�]V�Mv����9�k�:�O��aS����v5��9�:Nx���ݒ'�v�y<���!�,��6����w=g���Ot�]��ܣ����n����3�؅;s��+�����I��ۓ;���n(��\h�r��<y�{�q�;���ݫ��=c�����9k��':�k0�ج��6��vp+�;�-;y�!�6x�8�wR�k�θN5ֵٻ=���{�V�%HHM�D�d�6�d/`��r!I"lI#�'��vH'���h ~'��/�]2�7o�ʞ|�w]�~$����ll(��A�_Ɵe������bwX�{}Z���U�$�ue�&1ٗ�/L�&x~gS~N8�l5Cܝy�O��em�d��5�7�c}~��Ix�������c>w�YI�E������r�y�Kݵ{����kh���>{��>���z�#菆/g�k����*���eC"L4�p�9뾻 v�U���U9f��d�jG��&�o������v��@ʷd��č��䉨�)b�ϰ�����B�D�c;���j׃O4/]c[����?��@��ѡ��� �mm�����본������(�6����=�b�C+�n�HdG#}=�0�,��*mڭ�c!�a��9k��v�':®œݭU�W2-,����tz��ܗ\�b�:���=�-��%����G�)7�Kz{��Օ�}�]VIQ�YZ�J�������D�]�}��$ޮ��{��Vz��Guj���o��~��W�	G>�@�
��vT�ä��훷dO۝]v	�V��=ٓ��bhX'�������RE��j;��]J��h�ߞ�`�u[H?{}� 0U��G�Fԡ��r~�'�TSi`��ۂ������j�8݃�tс��.���.�:�g{�T��H�|on�����  ��6�Gf"�>Y��Iz������n�$����WNly%0Ah؋����1-����no�������-��@�Kýݙ����`�Lj,��f$���'�~+|��D}k�8u�U����:��L�ޮyܫ���к���w<��n���S�M~�m����EP��>���2���y�f�=᤺!�F���Iiz��� ����N�$Q%o���)��'0��eݚ��:㎽�׻VH'�~^��@�O�]Yn��mz���ʃ@ޓ�|<OYV��� �Gt$�em�~^���x��������P ��@o�%@�ޗtf�p��4�a�B'�	FO�P� Ʈ۴��%s�\��\
�Gb�h�s��{����u�rע�� �����l�B����ͻ�V�K��H
�n��m��6d��H������/�U�	�y��A�xhA�ʿ�ۧ\�*�yc�Q��{�魏"�& m��<{A�[ʕ���ӫ=�|����n���7���ZM0p6�Q�\���^�^�K*�9�"�>��?�z�o��uu맽R���$�>����둍Յ�[钑.o�E��&��X:�Nd��^=c������{ڙb�ɹ�o*�ʍݣ^nT\FJzjo�SK�.0a.5vkfzŐ��꿍*��_ߐ=Q�~ &���(>��W�C�{�Ut$�EѮ4�j�a����l��e�Һl��9x�4rԻx�n��cc@�R��~��|I̺�A?{���w����v��<}A	������f{D�5�w���t��x����rT ��$ ��#Z���y���C�r���4r��v@$�muY ��� ?c�8Pu�k���~̗�H.���* �@ɻx��7OE���_��W�,�����P w;nu��s2�����~5�m�̸��&d�[^�O�k�ߏ{���/�d�}ۻ��H (���B��@IO�@$�	'�@�$�	!I���$��	!I��$�	'�� '!!��IO�$ I?���$�@IN�$ I(B�`B���$ I?�B���$ I?�B���$ I?�$�	&��$��1AY&SY����h߀rY��=�ݐ?���a�? `  � �   P@  
  څ    
 ��h�� ���B�)U��@*��B� �H *�P( �P��@�}R�T)"�RR"��H*� U�HD�R�"  �B  
R�UT0 hD�*T�@>���U@4Jd�-�B`#�^�م� ���`��Q��`���*�F  ƹ ��mJ���@1�,��2��X#��w�J���U)x-k�h���7{uP+�� P| ��HET!@
�>+wG��s�:�HW�R_.�=ʇvx����n�9��*C�F���՞@u�P@H� 4�� {����  ���^:J��oX_` ݚ�3�{� ������ʢ��C!���O��<� y ^��� <��R�0 w�� �)T��z@���ԯ�f��Jvk�
OT3��f�d^`��u���mUDs����j.f�@��ʥ>�|z��>G;R���Ku;�^mUw�=}}W�
��֑.�E�UM����9i����h���
�$�>4$
��Q{
�}B;1J9eEV�U}��"��<E�Dv��c�æ�-Q͝��=� �-<����^J�X��� 9��U_,��)uϒM�J�w{5*�S��Z�����7<U^uPݺ�5]�B��O;U�$�W� |R�U(���I�EK6*��R$ݝӝ��n�g���=jU�+��u�+����^�
�7a�.���)��G���ﻩJ���R����q�Ү�����]� s�q���@
�Б��      j��LT�J �     E?&R�T�4�A�&� b'�T��U5F# 	�0�0�4�M��0�j�@a20A�	���i����MR�@       $�DT��1 j�MGꇩ�h�FjO��~����Y]7��섁��5]?��~��ۀ��������T?�d)��$!$��?�IdR@$�~� $���S��S����?��D���ʟ�4���TPI!�!$�
 z��$��a� �M2VX@��C�������Y�$A?��?��?��odBIa'�s����б!����ol�����~�z�
X$_��_������~�yտ�Kqh�vj�ں"�0���ItNy����&���&wn���KNv^�!*�',2k{�$�:�[��x|N�i�5͉�F�.[h��.���N���7�/z��<�S/�.!\�8��k��u�]�l�3`��4�5�x�5���7t^�j��d{L�i>�n�h���il�p�ͬ��2M]��FB�X
�֧?����G��2�s;#Z���$8���8���"�8��r �i��e������^�|�]�sU�d.ն��Q�E�Ꮣtgp����H	�DV��� AL@�O������D-$hb*���F��}0�MF�J:Oo$dBl�3��v�,�_+"�K�=��E�.n�E�{$�ٽ����rd3�40���VD;�FNnس���c��w�glؕ��wL#~{�!X�v�i;2��{�<���c�o��' �/ۏ�d��/j�3��^�6`wC`��;�}B��a�Nf�10uQWrXNn�Ӓ�n���;��M퀻��5����C��y�7��xF��Wk1�y�5��}�rn-[g`R<ǫf:��Wo��-�����=�n߶C��r�wR�О[-�˛����w�gR���1�+ygcs�ު��s�g�	>ӳ������a����w�h-�ϝ��V�Yq�(�r1Gt�o���r�_��+x�Fm!��f��`�`���Bm�֏����%�6��4���;�#��n�3���\����Y�Ǖr9�|݌va��k��t�NJ��rn���.�X�.���d��B�fü�vh#�IL���he��
Q�˪�Iy��
������P��j�G*t}��8���m�Α�H�v�l	���m�6e���vu�/*���>��دYm=�yL.�6�ת#wF���<r�DL�2�T=�øp�+�&�A��-\{��1�(<��He��;�f���}:-���æ]�!���a��Д7��@cZM�C���%U��HQP�u����w�E����
�Y�l��FOت<�e�s1x<��<���ޚ4,lu��Q<c�/-�@�,�sÚ�.�Z�T�ϩ�m�ۺ�má��07ƝE�]D�r�g;p�IN�'bM-/�	�>����p%n��Ω�^e���H��v�L��@��n�Y��vv���y��4u�z�]��n0�OC�odYі6-˻�r�1��Mq�7�|#Kt�W��X�{��:�f��5�:�N7�:4y���f�3�_P[}� ̙��-��]1�m}_h9Ɩr�gcV�܌���a�p���'"���oΦ�I��-�Mo���g����BX��92仯�T�oe
we��E�z���ӌ���������i�y��j��î��۹Z]h�Q��I�vK4mZ'lO/X�>Et�KY7�lVi�ܺ�N6kDesh��㽵�r�ۋA�+����m�����Bv�S-�ݶ��$�����Wl�dDn:��+Q:9"�#ۣ�o,6�39�7V(���[����pڣ=H��v���,�#��{�$�ḅ�8ٜW%��:�(�$�cY�x�t��
Ȕn����ͧ��B�߆Χ+�*1Q�sJ޺�іf�7� ��p*c���.y��{�m�MG��J���qhw�;6@:#��U^�6w&Ou��v\+l��[w���Q�8�K-�ns ���̵��N���٠��
��Ľ �����$Mj�M�$�Z�6�.[ك�uQ��ݍG�~��hk��w��C/B�z�Y�S���ws�p-f4oCt��jg^6�>/A�1�Y�ѷH]^39w=|{�H��#Ѷ�bۥ`�(��8�lA��npZ>��^X7�@:�����_��*�� �p��b8vQA�D�;o�oe�I�5�t��Dh|��>�>^���D���	�\�n,!�nk��O-���u�6���;�P�\���  {��GNK{X�t^ԟa(�)�"8{:bv��uüG��@�hq�	]z��S�x�o�D�;WG%��*�Wc�B<Qos�u�Y�᠞��I�&��U���]*%8�'�J�s<���Vsp|��SػCON��^�)�L�˔FL(?-�L!�W_-=���;�u��~ S�2L��wEN���V�^�C�4X�'��ʟ;t�sĤ<��7;65G�j�i[�OE�bX�c�6s`4n)���.�;	��n���q��.B+�IA�ؘa%�L�K��n�H�#����un3�޷ު�������_Lx�nt2a�{���d�x�,Tr���<q,J��q��v�I��I[vw����k	�;�ٝ�ܪ4͗�ۋd�+�K۷��BAuɐ�t3�����{����(ӤEn�xO�f�VNɭ��ڼ����ss�H(�E�H�9�Kt<Ҳ޸&��~���qa�dx哬,ogg\�)��x�o)W4��P7�W:s�I��K�Jܫ�F�@���|{��t1��z�kv�of�:��G`ܒ,v䗶e��L8�R��;~r���\���nYJkvt�˯;Ѭ��N���s�������j�5���q�"����].�Z[ӻ�
G*�[���`����o1��0k����IBȕb�{�-�6V�{RK�/���{V/?���+��H��v>ߡ�V�om�]|4g,R���U��$�&�m-̂^!�_k��-�sf�������TOhn8�h��gƹ��u.3�"���%f�aCYRÏF��8���n�eeכ�n��l׼����x�]�R��V�u�k!�ŏ���vk�a=ɓ�ؽ\ι��n�y1��V��N�wpWn=�D�kl#��"xi���Ok�ܐ�Q6�����w�Ҳ	L�#rɅ%�.��+�We�5"C�	�䵇v�	�-�T<�Ns���CR*U0���v�'!&H1���Ŋ;��G�f�04�.��X��%5����siԂ�XY.��`�r0�ׁ���ξ�dqR��Z��{�`-��0�uc�O@�γ8$V��vI%��Q<̺���5�(' 77����H��d��f�Y|�&h��2��/#t%б*��<�ԐG����K�����jg	�[����Z���u�đo'h��xrnx�Lށ���E7Sp��ӛ�0����S�Q �J巯Dv�W�a�gP��5&0�S��.:/����j�^�|��JV1}� Q��2��4e|����5`B*ُm�L��Y����8n��'�G�IX��ʲ;p�6PX� �.|�:[:voc�/��[����9x:-܃�~�j]�G�~���.ڶ��.��Z�fh�����-[���>�� IA�]ac�o-�������K�q@KWP��B{$�\��5&u��cd�<�t�6�<v��<	�O:1��Y02	 tzM�}01���Ö�}�Mg��'l!�qv��՜��A� �Ss�w^��!T�;@�ڳuc]Pg9Ў��1m؜]h����RG� ¥��P�8�z��qNvu���77�^�ݥy���C��k\�t�@�0�ו���'Mhd��v��MB��S95�v���wr�SW��&��Rlc��c��γ�����P�Xd�#��sD����K�0k�i0BKB6c�҂�{��n�7�u�q���{����0_r� ���j�q���ND� Uѻ;Nޝ��r#�nh�/,_oL�&xy=�x��W9���uz�5.B-ܥqs6�u�o��#8%�o3X 3Z�CUכ�\/�� �Ű�oC�~�ר��_b� *m�3^�؏B�|��.a׮g+φ���H�ipv��3z.�T{zN*sv=�^�_q��\)�&mYqcU��[L+���L}�e�-��fX��M��l�����!L��8��}�֍ɥ-=��{Q�@������|����0ZW�&�v������ʎh?z\lo��,�ﺬ,h*�Ix�1�W1�w"�4�=�^RK&4�Ďv>�j�nM3���huѼ�T�W/:my��]���k'��%��x������4gpZUeM���9(d���F�	GW~���7��.4�����oUdS���+F�⼻^'ڟX��1�8�ê��v�Ιǐ7h�u�ă�N�u['�;�<�*WŁ�\)��oV9\4l����}&�{�`�h0��"���w�F���bQNS�#R�ϵq�6m	�ڹi���Y�s�}��Y!ئp	�P7#}�Y }�T�v�j&V�g+�����Q�Ի�W����JloF!Y$����ټ���E2>Rk�'�vC��r�ps�}&w�Dx�����5Z��ƶ�a��,��0���(���ҵ̤�79 ҒuXh�6ocr�oAd��#�{)��[�[�
��r�����;Ði�V[c8u�n�IJ@7�i�3��:�t#�Ӳc��i�˅4j�j�q�NԵ��`��YPh�?��`}��Y!��8��K�c��B�'v웉h�)A�1�D�r�%`�ְ��ea�lҶ���se6�lU�O�)�C��2�:�$(�[F���h�9Nwn�L�n�,�t����7)��.\�n��F˭�3�.�����V��(n��a���p 1Lv���^��:E˸�2�m0S��[��,�Hb&ö�f*ō�ѥ� ;;˗$Mv7�]P�R�����y׏!��/t}��N�u���4��|��ԟ���)=ޯkYd�w��짮���~�����E~ƷNm8���]�8�II���~����ccf�9�%FX�}�nǄ:ш�pm�z]�X`�x�Y�Axm�<�����X�o&��$[���F��ΛZ%gb<&��w{N�^]��5�6��=7t�+قU7<.�,�Vr<�7I���W@�p��f�=�I�,����M��~H�ײ#r]�Ʌ�bN�A�L��N���7j]VR�N���L�vΧ��ٛ0�2�v��5�1='�
e]�1�NK�
uX��r���`��a#oc]��-{�i;��4�T�xpW9�İ.9nrېgs�uV{AUUOgt�^�-𨣽v��a�v��=œ�6"�k����rk�ڷ�������A���q��,4R�w�x>�k�p����g��?g�(���ݞd�pH̟���f~>Q;����z?Zk}������{ XI�� E�XB�*�d�H��@�$�RP 
H,!E VH�� YY		P� �)$�*�,$�X$*H �$
�@��*�` )$�B H��QI$�a$BIR@�� �(Q`� �E  �d��	"��� 	Y "��@�XI ( �� VH!* J��Y H��	
��XT� ,�
I!a ��,�Y  J� �B�,������C�)����韫�~�~H���A�z�5�BI$����I	��}��Z��!�$!$���3ӯ��y��k�i����C��xfȫ�Gk6�M�PSAG��)��T�j�e�^�E ˥��B݋!JN�<o[�ag�^��X�Ђ[=�2�D�e���!�����uh�wK�����v?o�׳��4�7CY����5��m�X�q���&=���,\{����Ux<��C2�|�Tw�P3�9/�P�ɞ]�;<l�ᝀ6��5Q�W��ݘU^��L0ͺ�#ݬ�A�8�W��M�Uv������[�e�y-���8���F^��z)zh��HQ��~9ܗ�E{�´�N���2D��O=�)g���Dx���;wu�Ǿ\���������_��f��7&�D3;��yvt��Ik�|8=�HXB�Cv��q�;�[��� ��u�~f3�}�~����b~���w�櫦G�6z`.C�]�gw��
��7�����.e�ۦ!n-�.5Z�E���l�;˯�����Oa��s��gW<��V\�o�x��=X�3�o�f��ڕ>��k%�+�g�s�6�k���{��Qy���ܾ^Q��`�z�S�@�]��XBBf��vW�aD/X��{6:0�F�޿_���5����ږrӜ�7r�����aᾫ���P�3��s�ᖭܧ
� �1�{��qn�|�#����8c��G5re!{�^z��з�qݷ��u^�v��%���;�|2�pe�����.��:Dݣ>���*�2��/ ���ڰH��|J����%xv��1�d����!>�g���W�U`nu���ϧ��'"�=�-��|���g��Gc��=W�u1�x�9uڵo��qo/?���_���W����SւQ�z�?{`ʏ�,7��ɻ��Ʈ���7�z�p��a3˷6�V	��0�g	���m�m�f�5N#'k�����8����m``� ވ��qk�����&�����{��N/`v��q��.�a�B���O4�.#�g��r�����Zz53��\�2�Df��Q>�o=�7i�/?iz�ߙ��!������A��ot������rk���#5Lz	�J9����G�\Z���3�G����++�L�.d��>0&w�� ���%OuQ�ߵ��tx{۳x�F;��=�`b
�!������q-o��3��,1���i�M�A��uk;//k�^�^�>"F��=dǒ�}̞������r݃<���X�png���K�^�+����i^��.i��m;�)ڼ7��
d�A������zv ��/Oi�L�^Z�us2v�u;�n�Դs�?��uU����kX�mf-���l��8-+��Ap�K�|��]f��?Ȏ��8 ����b��,6�����p۹�V�n�2�"]��cþI���n1�{����[�P��]����F/|{D,N�!zh۽���aT�z7�:�uyU1M�V��2ObhW�DnѺ_����\误;���u�&�hZ��;ޮ)���{[���i0ڥ�Hm�ޞ����+�W�N���3��h�h/*z�*ˉ0xk�ikι�n�x3�޹\�gyh�Otܘ������s�@ׁ"�ׯ�d�˧��x�H�n��{z\�E~nx��5��
�W�	�=���Vwt\N����OF�|TLi�3jʬ8�v���w3�Xs�ʭ�Qɖ�U��5�� h"�$�9�;zB^��O+�.;�"DY�*��i��o����V�dbͣ��j��.!�Z� s��?S�R>�������E!��V%�^��6��������3(Qt@�=���Vwg^Z��X,����9 �8�_vB'�����X2�`�r�����4���}�
��Ϸ�=�5��{�]��/}7�n��#Ŧ4�^�K�g%��_d���b�W-��IS��e�ғ02ҹ��r��ҍ1���\S��q *�Z}tŉ�O@wi���۫���<��Nl��I�7���"|��e�^ڔ���8��_wp�f��$
�/e����h?�=���\N���x��.j�t�d�Y�,/s������y�l��3������1P���I佖�M!d߹�~֘�:!���¶�E4�A���;����Q�a�*3�1b��O�୨g��r������Wӹr4�3���c�����/s����9a�(��8@d�bڜz"�9U�m��;7s�y��/3�)���Խ�F1�ߺ�ajM��
����h�lf�Df" ځ|,B9�O���M��� 9 �vx��2�N�7!���W�7I+��Jx�K�ϴ߲s^�q��7fTWp*[�L�n�K����7yǴ�� �����_G/*Z���^Yܙ�����n���=p�[����g}�_[��w�ڌ���[�wFsw��3�4E�I��};��xL�`�e͙�ڰigr|��P�/-"w��J�;0h����=�'-����L�]����3T���_D�k��fq���f��<���R�J|G�n#^�Ң��Ú�vz⧉S�r�j[B����/7�k��[*���;�:ukM�{�.���mL!��O��u.���i�yӭ�oqG���KPp�$}~��I��1Ve��+}���G���XGx[s�}����5���nt{�˜�<N�f����H����$���{!|p�OP��,�F�.�痻8��4N�#ݩ��w}��j=P+�_kVʏvH~LW�!��b�}}�9<��#R�ߕ��FEIo`(�%M~�-��I�LM��x�׆�ֆ�L�Jˀ3�T�gױ�l��|r5N/����}Y�L�
L��Udz�CT�g�{X��驠:�vh��^�r	�5n]ǆiL֝86Ρ�u�l�W#�o������j�E�#У�`I�C�7�3�4�c�k�[4�����<���(���|ͽr�F>����?n��M��ܢ-���w=[�t)/o-��ш�Ճ%��i������m�+ɘ��Ն�]�ƻ���?k>}�#�XN_b���7�6+sFm�V@��Z�����z�k�.\�����s���ܼ���i7#�q��=ϯ2�����D���B������x���K�sԮA}67��.���4�Ї��=�v�߅��o^����[	"m��k�|�m�=�9F���6�<�J��1��W����*�a���g����1R������s^�0�_�{�gʧ&Dq�"w����S��I˰w��G�d4v��wk�-6��!{��{�G ��k� �����	�&� ���,-�S�_]�7>���=M�dˇ�[9Z6x@��l�<�\V����E�F	���w6�*d#ǣ�1�ں�_xz&EZ�d�X�r�/�M?>�O.�s�R���E��R��	��^� �����F�X�l3Bͮ6|2���|V����l>o�KX���A4/ٳH��k����M�.xbŴ���W�0i$��`��	J�e�ա�����3�6�d:���4Y�~Sv�<��PD&�&lIw�� ���s���G�y��W�e�n�E����^����Z��j]Ax��ZI�[��*���_���3c�:��!�.���T�S��/�d�ܧhʬR��׹��$�7�@w��V��$d��b�_.�-ٜ�#�s�2{��ݑS�#�:���yo���x�Z5y^�Y�_-���J�6�UM��)c��;�x�'���M����]�1��k�j�*!\�0����(�FW~1�X���j��q����w{�&�-�F����D�����/0��"�;͛��(��ӳ�-⮇�fI���V���97S^��ǙcM�:�^I6�W���x�"q����k��O�G��^�QR���4���;ז�Ȅ�A���hq�j�e��/��ao�ᛢ}X����R�5xOm�ܩ�<��E�Q�Xğ/���+�tF��;w\�7Vg�W���At��D�
k7��/k+Wm�'3��߽�����b'/��y�؇������}�5���y4��ŧ/�>!z�W�.n�|��u�g�<��� >�";�q�3���;���Kٚ8�fŏe/\�h�E������"�N�w�����6V�F��~2P�k~&����x��yKap����<�j��i�3�1�j�t���/) �N �7|',/g2�b��rs�����q�N��������g���y�<��|��Z��c3fo�Β(�i�hS��������t9��q�:^��Ͳ�7tXE񅭽`���S�[��f9�<A�~3�T�O�gf�Ng���_L�i���^s�v��K�'��{)�WM�%�q�n/!d���i����{�K�ƍ�-�|���bK�Gn�æzW3F�<�vyh��F1�,]�x���p���Ozy�u,�Q��C�<ܽ���¾�μ�L��P�{��Կ0+}�Y�~�O��&�m{��|p�=��t7��&���z�n?!�fG��hҬn�KjdOמ�����|��������J�0|��Ƽ�9!���#���Oz^;�l3:�}/\�q��"D~2�O�8�˥���C�4����>+2����iʕ8�z�X�T�ޑ�nm^������M�<Q�Kx�����C�Q��j{j�(Ќ�;�
�nh@'��N�~$.ݐ%��A�w= �����CW�G����-lz��=:G��|���|O���!������̩��V�g�
4�����v^�R���� �]V�h;V�<��k!��L5��qh��/���b^ޭ�-�&�^�{J��9ߣ�:�h���=�1췔�j�O%|�.<~ۇ7۔W�/-ѡ�n��n2�e뙤<�~�W6$|z���8�I�	�9�s��g�=ڷ�}��/B/eO��`>��������'��$Ϸq�=�r;0MQxr)��55����������Cܣ��{���<R�o
��{.�C��;w�]ӝ>bx>�W�/Eޯ�"�n�3U(�#T�b���߯_��帱�V
������*[�#�&!��P}�ldlZ�uG��S;Nۿu���<�:��9I�X��>c7�ſy���%�ۮgQ=�z=��sO�r{�|���nEx}������4cZ/��OۧQ���@dǸ��a
ݼB��M�٦�bڼ���G��(3�S�Fti���V�I)���%��0�D�q|˒�sQ`~sԍb�d٘������qFV˷�0f4��v}�w%5?)��}���\aޙLU1���5���.\�#��w�OȁI �,"���M�@X`����ӆ���]�֝jܳ�:����k�9�uIKeI����`�*��.,7h�D��q���-���`�GG��fieB����)[,99����1�v����[r*�ZxX���1k�ئ�TɨI�ͯJ�Y�B6��^�Q�������S:�ĳB��l ]2��CB�B���h��l��m�f䲲a48OZ�Y�;=��b{���uƨ�9u�t�t6���%��:,k�wEv�5�(u�0���á0�M`����4ؕ,��k*�s��o<�Ƶ�h��n4�׋�b����H�)[a���Ė���Fl��X��� 1F��0�v��Q�)�j�q����j���56^4����&ff!�ny��R�ا���Ž�:1c�V�\����m��Tr�>���p�9�_X�v=���ۮ^,{)�'f�M��F�`��+�.7�R$І��TVz	X�y�u�윅"��7\�秒�ޓ<@�Ք�eH7L�y��K*i�����L�K%�2R;�up���P�[�m�@��Qۗ�8�#��Cus�� 8�#vT�������47a�[u��)��h�k���Ë��-UC��: �n;Y�n�������̧	�:���Wl�XRd!1my��5���ͼ*� ��m�h�����% ���fF�����]p� :�/5�4JV�i�b3Ŷ�צ;lt�[l��-�F�p@9Ɋ��F
�뮰#�5��>t�1�1i1�mI���a��m�Q�N4:v�:ʮ.0ڻ9�j�nݎ8�r��琶���+�� 276�f����R�5�4zA�N�u��5�5n�ŀ�kIB�����)̑٪M����n�Txn[� �]GXv!��]��6�J4���^�Ȝ�'	�bܼOl�1J4��og[��N�S۪����c�½qټKks]�=��6�a��#���#��®i��u�%�lKۗ�sY3�v|d���PU\+����99��22�6�F�Y]Uy�c�#�w,m�j7j6�<c�ִ�W[q8�n��q�n9��ԏ^��{���@v1��5$����	�&׃>�J����=!Q�)���&��Ҧ����Gh��R h���v"⍲<�m�&�Np 5����"F#f���+�۠�y�c;��ۢ�.b�,v��v�'���.�H��6nCri�띩�ˋ�b3���).K�q�`�,�eD�\�+z�y�p��c�zm��f�\K��lR���A�Dwk<��W��\��c��+���X�0(M�F��U�zR�і�»��X�m&�q76K	q����ëg�H����ώ����)-[s��<=���� ���p���G:*m��v3F�b�e�uj�#�$��jd�lY��%�;)�5(B/	���Js]���<�3F:����δ�c5ɺ���jN��+�ɞ�Ij��n�쾖�v`���r���\gI�r��gX.�q�@W�%ʹ�g��dVa�j�eS&`��L.�cv7`��F�����q���R���4�t@7Q�wi|<�Ѻ�Vjn���F���j�|pp]4@�7[�t7���c��λC]v��2v��W ��n���g��x��˚;{��ᓢl̈́�mezyz�b�rv���=�d�#�Bz�xΑMBh��7P\�X$6�Xrax�h�У{S�x���V��=#j�,�B [�SR[H�j���f\Eg�՛�/�v�^im\
�e;��2û']D��p�b��a�A��2\����^�������E�{���q`����kŰr�Ul��uu�8���v�CR��j�c	�V�7<O'n���q���W�'s;�湡э�F#�rlv�]e��D�	3����֎�b��[=.v:.��`On���(. {c�I�n9��`!�^ò!��s�f�V��vl�LT��f�5�A�0�����v8OW��l狧����N�]�w]��#`%ζ��3�Yݘ.��ཷl��g�ղ�׮�;D3'��&Rݩ,�İjB]-�6��6�iQ9�nt]A�Lqj��.w7ez�F�oQ��/D�Iݐ3]�`�*�9T�$�"j�T�#`��m�e!�v���� ƒ)v�J���V"�k�ؘ��λj(B�md����v謮Y�yy�ӈD�X����F��u�8�X����]�4A�p�I��$��R�n�L;)���ہ�.U�\���;H����:�Lv�����!�.��+-j��T��)M���7ḱ�{/=�׮�L$�i��
!��ގ�hY�0��yڳ]��J�-�ԅ��V�Xlq#Bmh�X�ˬj��4��)�q�C���]Κ��P�v7�];�	/�v�Nz�H��8n�x�`y��b��G5�	��`����u��6��<r<>q����2��1��.��XS9ƕ0�0AJF�8�o4f.�
5&f��k\�bЍ<ּV�)��B�۸�t@�T�nBLc�����W3(���.1YW`�hlֱ�1��]&�6��5-����-e���v^.��8kMXB�M�X.�GY]a��.�\�4%�q�x�n0Xu3�Cn�v^�W+,Q����bDz�#��Ɠ^�tB�ce����t�)�r���
��s��z�!�Kq¯f:��A����r{�l.ݚ8��$�Zu׈�jRⵇY痢�=�zkˌ8#�k��q�Վ�v�p�=v�iس�^$3��g��Mklrj�d���N+sFqҙ��y�1Ƶ���t��P�U�`�Zv���"�5�Oq���G�B�	�����������֞;C��^ڞ��݈��ڋR�X��Clܳ���zo���l�Q�e%sFUel��5-([	E�Ma���Z�̭
�C+�tvg�
D�:��)��$7-�x2AV]]p�#M�8����G7�5�4d�v�\l��#'��j�gA mI��,,������IH��S��J64�Jq�9-tb�f�u��X1s[��	Y���B�[fU5M�C��d��&u�!ˡ��*�4�cwP���v�$`/5��!�66�V�v1� ����`�hZ��\ZŔ�������$_^ ��Aqq+ۃ�q��ק�N�K9;f:n/��/W@\�׎�WOn��øv��[���7�uK�������s��4��`���WJN��w�n,X�WA����u�՗(���;>M�렮#��=��wX�2doNdk�֮�/<��C�N§oii��jv�ݟ)q*�ZB�ý==����F������p�[���Fٳp]Gm([�u��-���t�l��wE�O[�ƪ�����:n�ƙ��f�k�����8uE��7h[H���,10�Ҧm�讯/N��Ьv�V�kegW��Hv����nx����n-��t��\�@I��`�X�Fj%�.-\[\I];:2l�h�nԩ]��� �N���Rk2�L8e��v3��Z�`��q�B����\u�N�z�̹�M�Yy���w'B:s���׭l/m5�LWv	M13Zh��Տb���Ό`iv������ v�gA]v/h �iٕ�͖��75� ��%Ō]��9�v�Z]H͛K��it��\m�u�۶�<Q��V:����G9���1V^�����C.l�̲�ƮteqEc�Sk��0B��V�2�[��,Z�lC!BkB�1ڈ�ń�Z�D����I�&�\WG?^/ա�_�%��P!�):eH�9��
�X1�!R6����,)��l�W�V)&%VV�V(
 ��Zc*9IQBld��ԃ� �ۦV��$�� T$��X���2)XVP�LjkY��fY��RVERb�Nf��,��E+"�X�c1 c$���["���-*AJ�M$�[.�J�`�UFc6 c�,��-���j��0�Ѐ�b�XE%I��Y
���*�E��"(T��4�LI!Y�1�1`��RȰ��HU�)�PP �X�*�1�
(T
��" �E�RIQH�VP"�#&$�(�YUz	�gN���Cߙ���GCe���gK��չ���R�܊�[)6�k]�i��6J��
�3���	��w���x.]m[�`0�x�<6x #� ˠb��΁)B�ij��o2��x�{��jݸ���V��+to���J;�;h�-9�˻r%�Ħ;5&�h�eѦ0��6�0��-c�tWEQ��J�4�c#������u�$wc�;&�v蓍z�]��;%�;���:�q�X�-DT�4�6�*.���qp�Խ[ց��^wm�v�^������d"�Y�E��ۊ�W�ݻ4=���J��"�vkNސ-���ms��&A۷ѝ&N�܀;� �,{A���"]�m�A�muI�����u<<��{Z�hۇ�p72 v�9�������Q�,MS�bჂ�Mb��c�a�N�SC8f� F�lb
8�9�=��۸����!�]K�+��.�
���ţq�\^ST���!�Ps�����g���ۭ��2�R.�b/blUp:�Z��GF��n���8�[��V1]��:aMpKia`��ư��5��:�l��&il(:��Y\MA��1�lf��ֺ��WL����.@-ۇ鎵��7%�U�(��-�ͥb��,���(Ԋb��pv��n�V/��a4���j:�Ѭ���n�<ڵ�V��kl+����t��cv\�Ō�n�O���x�˥!�Ѵ{kH�p$u���p;ŕ�N8�N�Kմ)U�zӤ��y���N%q]���X�N�;L�e��2�F�Q� K)aJp�BX��A�+KaH-�%��%��%��/4cU#!x�1#md������%�Z�dTPR�e������"R�b��R� �%HP��R�k KF�bRZ�ز�X�QZJ��%��JDN�XBڲ�X�Q�b*�A�����g����]�D���������8�(�I%K��y6tM��y�_��	_�P��M}�U�uT���ۉݾŻyu@���$�=Q�$���;�s�z�H��i0��#D���$N���K�g���3~I|�K{�R($���d��E��19�b�l;]]��;�o�R�H%g.:I�oeLAiܵ�eg�D���{ll\�m��/'�I$��*��z{j�_J�X0����Y'	��l���7}�{��M�IH-1"l�n*������;,FF���}��S�|�˪��I.=q��}���$�9e���'���	9W]:�$#���$M�%���H%�s����sܒ{o����J�o kP�7T�=�s&bE��q���ﳊ���=�E���nu>-��~L� v2Đ7���&����apƫ�=<(sM����RcI%�Y��b�	 ���w����A$=��RI$��.��U���JH�����Í{�6$L岚$��ʢm$��*�����"�K)�*	.���s��aI�wi$O,�(z������B}�"��I+�˻E$ug*���s�˂w]pNМ)��Q"�h"�^5�u����赝@���\�m��9H��$���Q��+^r��"NRkM��~�OԨ�H,�˿�.^�x�24��-.UT��1#�]����0�Ժ"M����˻"P\�$�p��W���V%���"lI*����@%弡$���n_J�ǩ��}���3YO����q���ޢOT�^n'����|1���/IVa��`������'��O�)$眡�9CSi��ݬ�Up��Q��H��ڣi�����I}|�ޞ�G��@���k�ۤ���p�]��s�z�9�%/����ZH$|��R$�|�8Y���5(񔃡�۹՞��h��&^�g�E�:b�������ΩoQ͜�̺6IrͧH$M��i�}�CԻ*��ܡ�_VH�E�.�O4�UO�&vg���X�I%�ܥ$�H_;�I �)���]� ���24��,%ʪ�$�K9\F�I#�o����R���O{��H����PJ!K�rDؒU��w}��{R��_b��H�y�)$J�5�"i$�e�.uIXg �������{���<�q!�x�]����d��/#A��=/"2�|��C����o�ח�� =��'	���%nB����'�[ʩ�"s;*ū��]A@�3Λ��U��I�t�$G7���Q�K,���d�/�p�'јD�v�D���:[�Ӱ���F0䋆��%$�RDk�E����Y��4�Iov]�G�ҼL�uH���T����"s��[��X;'Q�1����<�	/���PH���.����7�9�>���E���q˗�eSK�]ەD�Jq���1�������M$�����}ⱸ�L˖=U6�8���$�ע4A%��vI6���9��Jӣ�$���*J!V׾R؎U����6���	^އ��M�G��T��$I�ܫ��I$�9Фf�L�"U��|���m!	��&`i-�h��N�.���=���/|DIfJ͞J�������X�u�Y�8,ưy����!��u��&����c�h����9�cTg=�2vˮ���n���:vY�����a������u�]�ܥ8�r�0tc�4^�h�g�u;=R3���0k��JPv���\M�uʹ�5�����凋i�k�M�6WD5�����{J8�GƋ��~��|M�q���UR$�Y��F�I#��RGMQLr~W�t�$I�vU����.H�V�})�_�{>���$�ۗw�I$�g:��*ڭ=������l2'>�˖�ݻ�H�ٮA*��o�L~I$o�*��K��}I}����h�%�Ḷ���[Vpnm@�5}�b�	 �.�	����LD���I}[wk�&���LʫK�U:_$���(Ex�z×��J���	 ��r�E���A.�y����u{C>lC�R{8�h�r��1��;g�:w�DM����~x�^��k�WI"|��:%|����+d.}��t�ӺۻE|�嚡�2CK������dD����Xx�yc��{�Xv���Vu_we/p����X݇�S���n�s�Z����=�]�]|�0��z�Wn�	 �ל��K䐵�L�_���f���X�*�Bl��&�&��:A"p��i"w1���2>˰%纪�I!k��<_��q	��N��~������"b��t�&�\tI �{.���W4��Q�F*�T�����i�\���ʯ�IݹWku�q>����RD�5eӠ�I|�{.�+[�T�gL���ˉ�ӟ"Ks��c�5�M�;�3�gױ�p����D�BI�ʜ"%$�om�[�k��HN�d��%PB����� fx� �caI^����:�ExoOy��%���h�$�~�2�P��h���T<\�f�r�A$��$��2�sz .7�er�yrR�ί�Rױ?��?Y���9>�i����<�F���"�`~��?a �c,��w��-xp�tx�-�M�M{�EUK�&�	n-��	 ��2��H$ug+@�c��|ML=�H��T\�L㉙�\��mش�Ir�SW[�`�J�k|�	&_�$ �s�����\o5g����@��ݸ�6Ť�Z28໮����+�̛������h�'��ʦ�IwnUm-Y�RAVnN$=�kb&�J��wiu�`P��2��\���D�L��Yw-IM �Iݹwiug*�Iէjj�'ey࡮8!2�RY͕X-��ާI$�2��{�x���ypI$�oeݢJ�r�Jl
��")�Yʪ��K]�-�p$�K7�V- �I�9U��+�t��zL���T��,vV��i�����ѣ$�Uᷲ��&|cG�1����fz�M���${וb��4���M��5�A�I%��SY�gR��
'}^�&I}���NO�a��>��_��n�4�͊�zIw�;��&�]F����sz�߿?{��A�#����ۣ$��A�I$��Ҡ���n�)*��P�r�Iu���#RQC��z@k�a�}b�K�mQ�I��r�i+�qM��ĳ-�����1BڕZ�UN�A,�r�H$Jk�W�B%n����Z��
E$�y�"iU/`q$h).�u]�Q:v�u>��jUI"P�wJ�K���^j����XIϼ�
G�}�"DR3V�UU�'�ޫ�I��׫bJ�ao	?}v2�G{�s�s����H�D��|`��~>�{~�G.�x9��i�S�=|gӝ�/Y����3LxK��Ü�֪t���Rd4��E��܏n�%�t��ݍK(�vM�.]k�zO:�[]��/e;=��BI��h�[2b�[s���ڧ@:���yN�C�z�y�$n�n[��c^�݄��ڢz�Oi�9����y[rC�������[vA�04](a�^�s, bbf��b�К;��R��ݰ\f��;,p�)�����{������]�W��W)��I��݄��:��Bi���o�d�7�d��3����G.Zs���Z��f��7ue�tJI�wH�N�]Q8��M�\�u�R$�.Gr�N,�h�]ەD�KՕ���u�J`I�k�D�K7��Z[��U�%E.�.UO�wb�xp���̛K��i /t������zx��D�=R��
R�.#�%��U��I|���Oj�)!v�E�$�^�˱h��,�R��9
NB�l���]�g0Z�<{D�{qj8�$L���>�")�9UW���ܪ6�+�r�Kg?�\���:�I$�[�˻K��b���a9	�	5�A�J��������KY��!���;jW=Ζo>zy���ϯ,nQ��˭Ut�)�|.W���v�w�_��I#}�wa$<��R))Z��R��{��R�
�[��H%�6���	K�)�)8U��$�G�2��D��9CՇ"���r:�3+�V���곛���3;j�Jך��&�\m�ʽ�<ۖ��Av�]�Y�ϘU�%E.��'�/�_%��TH�dFMS$3{n�%�Is�T)��$��V�א��[%�w�[3��6���Z�=���
kT�n�>|߿��wjo-ڻ�I$��uD����.�9w>
����_$qv�N@�ڢ$E#�x�� �P�
�무�K�g)A"l��M�A딻��گ_��t�a���m�߳v���c�W�����a����s���j��!+�t������9��[��O����Hus{�nN�%ٖ7`���9V.�{ZF��ܧ���������.��0�����]�}�Eѹ��7K�h��Gh�٣0����+*���t�.���f2�{�fӜ�!k�,(zg<1�=����g���D�h{��$��L��Odہ�F]BVs��צA�P}U;g���΋=`=yw��W��z詮��Jx�ñq�0Kֆ���w�v�#v����9w���5�P�q�-�i�eF�b{�֟��4𸷖����U�nG��$ub��EV�
�m��j=�,���B��*:�V:��������O@�>�T��η�Gk��V����xW���	����n����]�t��l;�p�~x��W�������%o]��{a<	|������;�[.{���j��<�NC�\�a2VEc\w�}_6�#Ңܐg��l�3��Lw=skY {���3�^ J�h9�f<ߓԴi*$ۖ��/r�����:�g�s�	��r���Z��:>��a̄��� ����>s�o{^v�K�������S��
�wi,����N˩���ߺ[��^o���7L�C�TE`�,�VB*� ,i*)Qb�ڑVH�E� �bJ��� �D�dĩ�
�$,X�E �X�,Q@AĐ�
>J*Ւ����R��*HV,����U�(,��U$TH�`���"0� ��Ր+ �b��(#"��PU��(�*�P�(��#�b�X+�)�E�ŋ"�D��A`��TbȢ��E�1H,�ed-�U�EE�,X�E�D`��
)"��&���߽����_����IZ�A!|Mq�C�T���Wg'|�s�m`I%�:%$�-���������4�S̓�[�ʩ.��`KI@j[U:��@8O���r7�-�l�׿�PH��n�|�'�����������B�4���	�'/Knf�Gm�Ne��vX��]����0��
�e�'H$O�B$�I�˲FG��\��&�I/]2L�0�4$�.�˻D��h�A�5�W��:v㤗�%��wh�����6�S�RK(S#�D�$F�iڪ�$�	{;*Ť�	I��Ջ��BH$�mӤ�I��ts���E�MbE�{lW�����Y6fd��D��*�V�K����~�
�m ʱ��>��_�ל]�ѫ�	왾K:귶����us�}��󥔲j7�4�N�e~�$��M��5�R9rӝP�K��e}(pn
�s��zX������h//��U-��m�/Mu�;�ts���#	��9������:�Z����"���shP$�B'o�������.�l��T�`Cn�����9Qi]Yw}pY&�����p�?R�]�}ُ3����M�7��6���"���y�g.&_�{e0=|�#r�21DH2E|�M�wD��ْ ���L;��^��L�ڥ"%�_&�F�	!?��w�`<Z>m५<����K�[�m~�ޫ�Q������ҝ�,3'�	H����4�����
�"4h�ä��P>���Ӆ������UB�:L���ȁ9@�ݭ,%�Vgb���،��	�3Ÿm6
�6i5�0CLl����v��&ѷ�u��kSkz�����.b�WY gd����z:�˻c����q�ڒ�E��!��eŪ�kg�v*z{j�!�vB뭓7�c=�g�D���V��7d���A�Z��\,Q��=7o���|�D��sx���A ����7z�?B=���>܀�w��vw���f#t�eQ��N�P�[�C�ޟg��n�;.�;���O+.Dk�nj�����n���ֽ��zM�������jc�"16H�#��ŀ����M+��u���#��5�9^��K���8� ��_O7��f�q����� �۪��{�	f��+2[��h �_S-��u>f�ɮ�kj9�z��S�V�/�_����>N�l4�(�m�n� wsU��Z��P�nܢn�b)$�-�����8�+��Z�Ɏ�^�{����GE��L\6�[�|�y/���}��V�/~;�^����o���̂I�uD����	��{�淒�'ڴ�c�
d8m�ٕ@�Gv�A'��w[�6-Y�TI'w�#j���(AR;�x���z=g���H3�S�wX���Y�K�����@�.�%�l���2��y��_�*/�G^k������z�Z/;�C��.�Ĉ%�c%(�L�`�FЕ�O:�av�[O�V������]����$"�y�B�$�:}#��ZRxht�_}�C| �L$\��9���<kے���.�a$ޑ����=K&�t���$� �r��Ko���:�	����8�z�9,𽪱eK��7U��`�-nWWIJ��������)�ft*�꺣�Դvu��/J�� �~bO��be=�$6�<���
N2��V�~ ��8Gw\򧜆ǓA�#ұ�*8AR;�5�����kv�_��	Q��]A'�\��F�]Q��o�G�HbA���Z��l� �۰�<q��!�H#~���D`��'�!$�ޔ�{��9j+Z��Q=M&�J�2}�
уS�ۋ���R�Uþ��⳧;�!
���@��uI �QRxn�z�߼�&1L���¾ �Hv[T�ڼQ|yXTv�@�wu� ��+����o���`�B>�$����w��ߐ���?���r�>~�=N�ayަ<i0J�P���.*Ì�s��Lֶo0��۾��@���s����fa-�����Ơ!�"l��<I�����R��F\0B�sn6!G/eV��O^�[��|Q���5l&�2:1�;ƃ���)n����y�k�n[��.O�'snP$Fo$:!��lH}��+���4�]KF�#BA��!!�y����}������w�SY�eqY�)oђ���n*��U@�s9�I��=[�r�A�����3�+)��MHH':tu�3:l���] �kL�}Q��t;���n�*���5�D�r9a.~�x�F��<ng��.� ���_C�沮WQ�RQV%���T��<sAc}����U3������/Bw^�`;�}g���lH������o���$�M�쵼oy�������A�"���
�U�+.:�u���:��ۺ��U��b"�q	,�uVXꥳG]�<��;IpA�c��</,��d��m��f���8�b��]�Zx'v٣�Hw����
�v�3�ga��%M0c;J��s���g��P�zv	ݼ�9�@s7!�Aٷe����T�]�"h{���~ia�����?��퐒���_S���]z����!�Vהr|[���<����d��#U���3"��Խ�q0�q�%�$�΁�I�����=��H�|� d���?�����UR�����'vO���9}�]x?m�z���f=^"��^0��$��l(�|���to�~���V�L�dwC�u�|u�����!�d���fF�(�CS@��Ɨ�څ`:XK�T������1�{�o��>�2I?wu�)�����S���Ft?�mOd�Ċ4�'�ʌ�޲���]��a�<3r�=��W\	�<g��^?g���>}�U�*wV����`���.�����}��g������0�W�����+���w��^k�}������m��-����ɌU��sz௫�<�a��fA��[�trY�X �2���n���~V	�8OHwZ0'�R;ݒ}��t�r��<�a,�''8H'7��	;��շt���*���Xm�>�2~�(�4���qn׶�8��a��f��	�\�9
;́�Y����9�ҖzCΜ�O�}uD�s�.RD�2�ڈ��B����uֳ�A�w]R;���M뾶2[�$�)A"��y�D�{�B	9�s�פ��`i�~�)����Ϻ�d���SϸE_O����n{��ӿ�z�]��8��C��(v���(����|>��r�߳���A���l�k�G��_rhQ�ɬک��:�>�A��s��ӎ���C�&.��	�2���h�$g�YC]�EU}T�E�Ja�}�{�{�����θ�q�������)Z�3@i �u��6��s�����R����s|�����6 �/���ћ�W�ޕTH$wO���_&K��IoB��r�\t�oc�@����+�'�+s=�Ն[�շ��ʖ�˗j#ؘ.3a1g�g�m,�4�.�p5���)1"�.�4˽�$��Ākm��� ��wW��t�;2�z��O�����1�\���ɡ�����b;/�C��	=g�6����EF��{B2�~���n�_�� >�|��g�����)"G��.���}4�{Y7����;a0[ݕFU�z���³�L��,�n8e��I�e�^�E�7֩��������2��M��I��W��0W�ԓ�k�B~��[h@��H���UW�<����]��� �u^�I��JB�^����<i݃Z?���pQ��&Vv:@��sY}�8���ޏ������9�Jrܺ�L��[h!� $��� �]��R�+e�sR�lv��h<�	1"�-��~$�l�{UZbbW:������
�ޑ����7�z	�)z�k�S5�R>�o_�l���u��Ĭ5�庥x��#�*�l�����oS�{Tws޾���i�����<���)��	����৲:�s}�ߘ�:P�J�Z��f?jtx�ؼ���ʳ�^��v4U�^�z(�ɤu���I3�O�yM:xz�W��S��������n�ڻto��|r�^���;�y�x�s�Lz7����<9�z�f���Ï[���gc�|�3:�0E�W���L�x�w�݈�x�������;��z���<��4>$�}5�NJ53��4E����t���Om^�������
g�Ad�9[>�W�sϺ���fU�(ﮏ ��^������vB�~�鈈=�QsL���5����k�����{/��徻�c�wKY��ea<NvX
w-�zH��hc���p������2�#�n���>� �;W���Rb�lP��9�DO!����b�=A�	^�#-�;��Bv���x�|!~�xxJ���[����m���2�4o5�6u=6���f��gɾ���[�վY�F�L;|�)����f��x̅�7�?c��Z6����|��Y���jx�E�� �"�b��AH��d�PRE",� �P �D"��1P�E��XE!�����@RE��P)��µ"�!P��d+PV�i+��)PA �
T���ʂ��T��*J�m�
�X�eAe@F������TVBVB��PF ���
�#lPm�Y
��YQJ���T���(�V���(V,eVVJ�%A���g]��p��ц��Z��Z���e�\X&�6:1�Bl�R��(��̈́��E�!5��i�K*��q����lC�.z{k���f�+X����V�j�#��@ǛWK�mϭ�9�5<��z U�m���W���r��1m��ٴ B��rmI�-��uYe16��n�u�y'��̎ʣ�r9�vwk�^"��4�&|�!ĸ�� u��u 1�s���EY�bZ��^66���F�Z����	fBRjjlVl� �0�ͣ ���U��vf�;I\cbF�wNc��=9��b�c� D���[ɨJ�Sf�lh���Z�C���2���L4�SF[B�<�Z���u����<��I2yw]���V�i�Cb���9v:�S�[G��q:u�OX�\�ܽu�T�Eduu�ۗ3�J����J)�]�X�YlQM�u�����[e���f���Xذ&"�·�KE%���$���qњR0<��j���K!��8��Q�9b�0v��ؑ�֣{Yܷu����qB<�9'SW�SF��dz�d������*�FSkD-m% I�&��Q��];�t��ǵg��(����f�N΅�݂�]�Hs<�'k4�����pz�u�1�1�[nu���\�E�}u��&��۲
n���dmF��Ǭ$ǃMs�.�u�9m�:-vO)��Yթ����fjV����c��"]kt�&�]�L���M)�pX$���1n^{CÂ��$��$e�i�6�����P�p�5���F+3lF��&�$�:I��!5�Y�B�ؐ���)g4]m��~wx������2K5B�ۄ*���22��]&�U�f��Vl@j���QM�Wt�8�{&�����<��r�Sn���{cI����j��N5p��]l\�v�g�<հ�p��t����K��jv�W��JKc"٦��<Lx��^�[��Z��v7i�E/ku���f+?>�'��؛9�����@�����'{��L���s�?�@H���+�<#`��fJ;�B��k�=���f��Q$�ܺ�	��'ڝ_�~ۯd�}���<��$�)_mU
 �w�1��[��V�8�U�]}G���.Mx��5.\���~w?\�"��������x�vrp��N`V�W���Sx�B9� ��|Oǭa����=��H �����<4
"��Zfǹl�q������3D�uB%ŻV�89�>5��^�κ�_�>�x�y�эG���	���?~�|a�sJ5�px����+~QH��:�8os3�{�ڽ���ZJ��m�y�8���wC���o�]X>Fxr�x���:=�`	fl�������P��~��������O�A?��$[�0��^l�u�վ���ˁ�����\a ����M�dg�@���s�nѷ"i��77k�Uy�����Eg����t`��Vfmm1w[I�jk�&�ˁϠ�����t϶<���i���L7��3��vG��K�ۅ��EHf3<5��7gN�&�5;V�I8M�o[(G#�
���7�I���d:�+E]�BF��	�k�u�F5��ܺ�Ë;��xߐ��K��N�;4{c̔��2F$q݂1��pP��t�6���/�}��v/|�u�GA���c.۶��-��ro�'rCq�����֗���Ms�~_?f�?��[�﷖#`��fJ=Ы���焂/z&�n��{�|��.b�~�	�<�a��U�$�$�k�����!����'��W7��u���@��
0ӖȔ��/�����஽-2����!�"v4{���޾V�@�;��g��
�KٗTM֊m.E#w`��Y5�̋�c��FvܠH$�O�ڮYc*lC�{!+����,��;�뙊���oG��e��o���2�cm7.n��n�37<�W�]\������;"�ժ����Mw��s1+Qq~Ή�Q�<yMKa��֭t�rl�����;�T��Bo�u�hR֥/'�������j�3���A�̃���	�5�1W���ظ	���>=��B8�lg�ey	\�$ԍ�ъ(��a�VGic�N�4x�9�pk����`:��袛���~�t��8��?`�3}9ߨW��{�����@�� �5!32ݙe���w�����:M�g.�`''
m,EE"we�����r>�NG"�� A�}���'��8l�Ò;�m�\��AӍ���uOw]3�++�餜�!}F߂�A$���qB~;�r����UԘ� }ѹ	��]R=�E^����VtfD�����I�{���{�%>}��oD��A��w��]�E�8m���;��i�ۘU�t������}��/�xJb0�)�an����#�3�E��v�a���x�γrX�Z�Ҙ�P�.�͂�qu�;��ѓu�c\nй�f��s�D�m��s�η��z�䃭�uj}�^[Y"}>��a�����h���=�i��k��`3K��+u�[\�#!c��^���mSt�]g2:�����N<�Z3�����4C����h�O����Tr���vucI��G^��z���6;�Kz�����_c> ;�,>��B��^����U�]������Ɂ���O�]OD"��^�ނ�����$�u_sE&�$�����X#�J���.�@Oo\	;�ge�=O�Q�N%tEa��cQ�]2��N���k�wdN��۔	$�s�s%�8F���l�M5�B.�㙶���Qi2��'i��H��WϿ�~���J���rB'snQ$ރ�m��Z��:���#��B���B�D8��=�A=�s|�<����<l�̸Ĺ�e7�Z�o�j��g�����,�q��̀���OOe"�/yâӛ���b�/����޷H�~��=e��r�j�A�)��c�]=UBޖ	�{���,��_ ��5Gi_L�R��HQ���tV�컷H@wkL>=}$u����[��O�;hP��I��!$n���#�$�^�VI<	���|{u���h�or�q��ƒ(Q0) z͕�����mctxд"�P<�ԗ)F5,�U�$]�i�>���Q���u{���T�#��o�#ppۑ���ę����
�k@;<�|_K�1��ʼ�Տ�ϰ��0�!�̃y�B~��� ��������/C�=�U��TЏ��������.[����w(��&	ݜ��=抲����jş��|�G�w����/��S�΃bS���w��\�؊y��X����h��X ���R��Q��<�v�s��� Զ�Ĉ;�D��u�X�݋%��sM=�� ]�uE�z��]��E��6��T��<��<&B�:�ٍب��h���F�
�ЂO� �޺��A����j�@A<��:ƒ�#IF��}2��}�\+���y�|I��Bw��	�}M��g=�e%����KS^$�u� ��"��Cwzk�G�ޖ��]Q[�m��Rԍ���}��z����w�T oq��Z�>���G���o�3����3g<۞]#�FzB�X�%��gc�:�g�9���$��}뙥��n�\5��N��3Z<Tf�i�dT�B���/�A}�Iot�G�/��ӥ�0��i���ѯ���R��q�\5c��8��t�5˷���������Egc����5�#�oM��x&�=(�Щ�h�$n��A�2w�16�i�'�}B�;��k3G�[
餋�RQ�1��A��`|Wz3ד��^����=�� ��iy�H�JI.�G��cΥiwm��Vy�������Cf��6��
���BKR7F�0Z_@�T��̗��J�$���Ǝ�.Y�ܧ������/N���Q�vQ��T�[uzʨ^�`â��^���Up�׌�r����F�.�S��V�/ʿ| �}7�w���b���BdhH���M���|/��	�8�)�"ku�� @���]-l4Xj6w��U�,�T�c�l�@�{�8,t����7c�X�WN�%d8���!m>�a�lI��������vT��԰"8׵�b"gF�@#-�s�P��]��-Umǎ��8�h8�sda��V|�W:�%ݧg&�_��4�MH��G��$2��O��I�l@ EwJےT��P��A��[�w�_6`rDh�}$����[�^��{�BI5�� ^�q���+���JR6��O���+�B	 �����ۗ�RmH�lI��c)'�"�Q�~�ɭ����z�A��	 ���OA�k0��D�\�dI�.�!l�BG��(���3o7�נ�UL@I�� $n��ef�[W��G����4�CD0�����D��5p�j�Y���C��8� {!$���Q͓A{=�=y'��p�tycb2D�Q�a�Yf�K��z��Փ���w��m���\���)7oa{���T�r�f��k[��4��t��w^��XI���p$��;�����ɯ����}��2��W���;Q_9��-�4Ў��@�Y��ە=T��=ݔ��&� ���t��5;�G��R�w2�>wv�M�1+P��S�j��OB��G��� ��"?~� �
ξ���	�V_���L6¤�T���H)��T�9��M�j��ǿ�x�5<ˆ�`!�6��\�8s�ֵ��s.�4�������f���Xk>ރn��
��6�^���R��4�h3���a�zL�/��P�6�P�*>��H,:ߺ�;��Lю���t§9�I��s���sz��bë�;�J2�T���6��jAHYi�9�l� �{��yν�u����P�c��SW�~��c����[V/�}J�2T��a�&ТJ+H��Ox��y_��iY��a�Q��L���9G���/���QK��盯�+���n�+q��!YDl��a�ϩ�����=�&�/�ӳtc�u��/�zd;n+wPܻgB���z�%���O}�^��y�'���{����{��M��)~�\��%ܥ:g��6�Nݢ*�G^��m�Yǻ�lc:�<��|����r�:�/�v�����\����ܘ��z;�-��q��"�iݾݶ�&��BoҤ�]�2{env!�vDJ'L��'j��e������wk�������]�A�$������ؚd,)&��{�v�G�h�ۣ��:���i��ܞy�� ���8�V��r�BWɇ崩�k�#xb�.�hvݍ��>��n�BE�Y�gw�;�~�*_�'�3�����g�1.�y�$q���o5L�qv����L|��u���{'#}q��7���!�Ȓ�~�^j;��
ژN���v�=�l�����v��q��[�^U���]�=�U�R�����^U�����(a�k;s~���*��́�1A����m�j���o��;�ے�]�{�w���S1S;��>~�۫v7���p9��n!��Q�Q��_���esc���a��O~�\�S�<8�
�Y�2�Q�m�
֊�Jʅb�"0X-l��ֵFB��b�%J��-���d
�QYU��JUUPR�R-��1�mm���*T�JZ��0�"�*�A���ذ�T"��j"��H,eB��VU[J�"�b�h,�@Qe��P%a�8�Z�EX��U�+RT�!R� ��J���`V(T���T�T�Z"�B��+R6�V��eiR��BHw���0��T�����ǚ:H,����?.~0�M�w^z=Mc�5�]����S�_��x�]j����|�� s:
$��Z��Ͼ�4�
� VQ:Ϲ�c3\�3�������C�*!��jϕ���sUǜ�"���Y�Ϗ�&k����
�Xuy��i��{��_s}�=�{��Ѵ���5!m9����
؇Y�j�`T�Ϸ�Yq��o߿��rZ��;��,���P�b>5��^�κ�__����m�ˮ��$�{�GI�2T����m&Щ+V����0�
��ﾼ�n�3~@ߜ�F�:Y(2�VT�9�؛@��_��ir浛:H,-�H)����s��9�sF��*Ak��{�i ��+(�g9�c6�P�*��]�s����uގ�}V�<��&�ю���5��ID+%X{{捌�A@�*���=���}gW�O��R
AN�����]��s��;�
��G\��5T�:�ӱ&s�h�3;���k߯=䂐S^���B�+
°�y߻�$��do�����c�����3�>��z��f�c��!l����n����~�'�n��]�Y9���ؑ�����J��G����$��O8ʐS��bm����z4�њ֯E`t���c���P�nAV��)m�ϱ�����,�? ��}�i6�R�e���C�J�H~�(�,��w�{��mĒ�����ٮ�祁�g�J:�P���������IM����R�Ci(�d��:��F�4�R
��l� �9�������t����`H)�!���C�����n}�۬��N������t�YY+<�����k���:K�0�I�,IXX°��&Щ('9�4t�Y:Y:�|��y��~��gɼ������-�K�5��������t�R�<�<Ѿ�
�0+X>����w��i��R�����1�d�X��}�<Ѷ0�)����J��i�L*s���}�޾��{�|�d��2�C
A@��=�gL��R
s�`�|���~�RD>��P�q�R�h��i�3N��Ϸ�i�ed��%O=�I�5ߝs�O�y����<a��a{�u�c�*A@��|ѶN�Y(��FT�9��M�k�=���w�֍s:�,�.u�&�{��4ч�t�v˾�0�݅����k�P�Ǽ�[��*�������G��q)#m�.��1�l��-<x�h��c���@9�<+s��Smw4���f�X{Ċ�m\����tw]������񡧍R�q�nl7<`�8�j�G��6���xK8.���0���Km`�K`�^K*m�6\�e�h�`2��ۋWb�1׮ �����V4>.Nsl�	u9�K�abX�e�mW������tu����?!�<��n���-���F��+Fk��9���@���~��}����A7�桌�%H(T��,�,�� =���YJD��<~3\�4�hVM�\=ק�f��>��Y�JʁD���4m��Ԃ�/�ߘ�!�$|	��{Jg8�`��>��!M�H����R��M�����T��s�6�hQ%aXV���Ah��(RO>�4�@���N�R
{�`@���_E�Ƹݏ����_� �o7�m~�K�H� �{��F��+Fk�>��i��Q:�sP�g}��z���d�"�!/z�՟+G��%���cR>����}��JVKX{{捌�&����}�;@�T�\�gL����<�0�iHV_��c�����>>�m����)�$H�\��z��q�X˷GW��ͧ�&�_��Đ�I�#��}��t� T��S�y��m
���+�s��$������}�k޳�ghu�h�'���2�VT���4������:\њ�^���=��n���p���w?��8}�g`�$�ʗ����뮰������O׏�����{�5z3ۖ���9�B_�ߟh�␭`T����4�bJ�YD럌��
AC��x�������a�
��{tV�j�n0�aS5���AH,:�m�d��*�x��Z��g���� �9���A�!Z�\�Cn�)��7m�i���t�������2O5�����YO!����$w�4CL �=��@~�;��LR
u�a7����V�k�������w���B��-�s�y�i������_O z�0*}�x�
l@���s��l�
��P��y��0�y�˽Em\�����X��
�"�7�����N|r]�
ٗ|��·Ztc�CI=�X�J�d�+��f�,e@�T>�<س�Q���Q��u�Q	�`
�)���!�l
��G_Wܺ2f�ti�Nk�h�:@����s�r����}ײ|�{��������ja��H)('9�4t����YY7�}y�~��w�G~�>�Et�`.V���}��i!K@���}�hĠ��W[�3\T*��s�j7.r��on����q��;˭�/����f�)�o��hO]�N^��Ye���g�[�陔�
� V�g��f�*IP9��y�i�{�y֪Z�W3p釣
��0&�_T�����}�G���G�
?2AH(���gL���->�0��_������w�{�T����Uϱ���l'�&��tt� T��S�}�ěC�sNs��{o������`°�5��
�c
�RQ9��� �t��YS߹��m|{���G<�[M�&�D�۴[19β��lĘq1��i����M��3G/��5��!m�~�F��+Fk��s �l@����ߝY��z�Y���bJ��=�GL:Vw֮g�Y��nH)�5��Ci*��u��9���Μ�^La�3�B�|ʐP)�{�Θ5 �-��s �AH*㧽�ι�W�K飧��4d�u��q'5�Z:N�++%e��=��lI��+��u�g;�a�aRX�IS�s�2t��FT����M��{���:2�n��T����h7�\�=�^�H)��֍�R ��S�{�i �s9�V\�w��}��W�t�YX5�w&f'z��~��Ѡ�+W���ձ3�jA�粦{�>h��%c�<��}m]��:�mߚ��I9'h~%B�o��4tè°����;�Kut�u�v¦���؆�T+%Xu���2s����8{�E �{�}������jB�y�`H;��jg9�c�O���������@�l�/K�)�4�Յ�vr�3i��>��w�<-�35�@�5捤p�����9��6��u�sp�T�}}�������c�q&����GL�2�Jʝ���� �z+�8�?���� �#��H|8h��5�� ��
�B�0*AO>���J VT�ߧ���$
#�@����R��F���4t�X|s���?k5p�]CL:aS�o �M�Ro|Ѷi��T�y~�y�4�:`x�jAO9�{�R�u�桎�,�K���2]:��9�oFӮe�)�4�R
s��Гi�aX_3�7a� �s��F�:�a�o��t��*ANs�H/\~:�F]�OEH,9s�$,- �w�<Ѵ���k}y���t���Ns����Y��g=�1�*AE^��՟+>P|��F�s����W7��zH۪s|/5ǟ���G��_�,yyX�k�'�P�~ߛ�'~�껪�.��`>��O^/���X����m*�l2��A*�k!��.r]5,ւ�؃�����)����B㣭:�&�y�jڹ�7L�KQ%��v�a8c3:�e����c"��qJ� )���/IV{�0�X�7h@�`�L��%�6U�Վ4u�:뛬�`fط]hw]�'a�ܮ�ۊ*S,w&�dUEy9���l��T3�m���}�Ł�W�����¦���6��Y(�ë��6�2Q� �}�y�l�����}�߉e�k�st�JB�C���C�
�]{6\�j�f�IГ5�tt�R9�o��ܚN���;V�aN��w
�`¤�
��9�4t��ed����P�셧{��F?�>���t\�gGi��5��q!m!m���ꐩ��Q�+�uߴy�w�=ObH,����P��%B���<Ѷ0�/��]��]\3W�i �9�����^��a��B��}�VM��
y�<��A`t5!m=���|��h��-h�>� l�>��B��Ϧh�t�;N�}�������� ���������_��>'I���k�¤�B��}�<��Ad镒������u�}޽�X�½9��V<��f�-�&�ҕ�U�6*X�f�x������4��Xk���6�B�B����F���9�`H)����w�~�^xʝ�^� ����|�F��7��;kn��Ρ��Tֹ�i&Я�W�?��Nt�?K7K��Kyx����x�qtŽ�Z��a���ɾ���c�sY�5��~C�o��R
�*<�6�������`H;��x/	QL�>����G�"���xR35�N�f��GI�e�� �9�m
����`��u����ޭ��V�*K�s�4m �t2�VT���lM�Y�yۇ���sW:;H,.g4�㛼���� �9h��h�Az��R��i��@���9�Ag�{�ގ�����$�Qs��t�Xw�tk>�.��i��
��XCj���ߵ��}��:�}ߕO}�J����}���R
B�O�� ٺA��js��l
��=��=:�nպ�ֵ�9e��n*{W	�+��{n�;7Q�'�R������]�$�9s_u����R
{��{m �}�j��5{{�bs��GL���ed��Ͼ�4������4k�OE`t��z�m�itk��k��`^s�6�R�`T��p&�*T
ʝs�����T;�.��}��<��z�X|s�-��[r�����Mk��H)�^sZ6��YP�@���A��;��=������M����ہ�V�+�V�~�f��C�=�j�r�<�>�T�T������H�7�$������� �� Ґ�:�~5�)7�rl��h�f�H��F���w�q�Y�����5�0ؓhT���}��Aa�%���4m�����w�w���q� ���bm]}ۃ�7U�\��Aas��x5!m �}�<Ѵ��xi��}��<����
�YS�~ޠ�q��~�6è°繛��Nu��:��vO1Y籭NZ�n�i���n��Z�6'��߳�{��ܸf�!�����!��B���h�+%eH(�s͝0:k����{H)y���)
��sZ��Sf��93FK�]�v�9δt� T��3w�m����]��}׸�ؒ��
y��
AI�
���9排'C+#�Ny�k=��4��Obm�~u�4k�N���9����R�
=���R�
�S�޻�h��1ߠi<�*aߜ֠�q��RT*}�4tá�a�g���k�D�|��g����K�=�2�f+R�|�OYXw�5�l����@�}�:`YG�D|C�� z����
�P��W����}�	�����i�[M����;��ā.x�69�͊�<�Fg���ߙޯ�߾��Ē���+P�}�� ����l������t$�:d���?���M���Y�ܔ���Jö��w�AH)�yލ�xʐR
s��m6��u�ϯz޷����-��;vw�l��0������kZ���]+4����e�nA��=�8��u�)�B��s��+X�
�}�4�bF��y�n߼���7η�,��P�%@���F�t0�=�:.�n\3Wp��T�:�؆�PB�u�{�??g�������`��FT
��~�͝0:k�!m>���H6�����\�P^��R�C��:3W]�3�Ѵ�@����d���4�ĕ�V��y�z^��o�,;T�
��<��2t��FVJ2�9�&�h��u���n�����sZw׽����a������]��}�h0+X)��M�T��';�����y��k�6$�T:���@°�o��;��Nf���Tֹ�i&Щ�;�Z7Y<�}�̺�{�<�m�P)�s͝0:k�!KN�� �Aܤ+D>��l
��K�8����U=~^����-ړG�BܶN;S�^��S�Ï�֕�Y�G�˽����^��o>��IǾ��_Hu��\�{ӻbi��gV���=+ݾ���#j42�Y&��i�y��c����y���`dg|$���"��R�Υ���i�g�K�4����Q{��Gw%��=���03٭qrr!У�ڰ�{�/��qX��$��w�k�������T��$yho�h݉!
�f^�k"��
�~���5F�k�%$��vm�r8U=�W~q{�3N�0�͓v�4N0��m��������j+�hf�7���UVo8���5�فP3޼u0@mkJ̞��A�	�F��`�Gε]��ӷE�AȢ�ʫ���7��g�h,�r�n���ݏz��:������٣~���� h+'^�U��^6E��*g��3gSg��E짳��/��֠�o-���w[� }�/#C�dLۦ�LH""�
w�x>��Qz�a��5��yr���Z�hW[�s���!��I�<,ђh���~�=6[�|��1R����Nt{��P�P�7�㝋A�\^ݹ"~QH6I���ѻ߻���{}�������YЀ�V6���&�A��G,1UƂ��d�-���b"��J�DT�V)V�*�e�s2bbX�����YYR,ī����EMP.6�l�+�V*��ܵ���eێ8��[hŨV�Uk�����\�E�V,�DQ�am�
lUEPX�Fi�p�EFc�Tc�N(�-ц2b���4��&�ƴ�ĵ��H�,Y����t{�����k�b�L�nuW)��Լ&b�XY�MF��T��c��y�3���f��֖�5��fl43�r��6qn�s�X���=���i�9|5�Th@4�UڂҺ�1�5.���WG������!n��*��;�Հk6W/���K�HK
�@f!�SB�Yq�q�����٥��#p��)��n�F���w���)KL(�ʦ�#�X%�E�E��R���+�\�Xn�c�kk\�:f�n:1x��T`wR�瑝t��N�ٚx-��A[prBq�����OB�u�a�W��*%�j�A� S�]\��pr������۷r�!2�pqՎ��8�\z��wEoYlq�kz��l�ۈ��0��B�,,�f�%�t�� �msd��\�)I�.0�X�cu�F#��l��R�&�������%̼N���g���g8��9��	hTF誸�m�2�#ڵ��;t��SX�_,�9'��c,q��wk��]����X�'Wa2cv�\���Zd�w+:�Ӛ6�ṓxP�\ :�F��l�f2]�6a˧��#qv.��)u�-Ѻ�3���˺:�jgJ�Y���f�4YpHĹm	Xnl\q��b�5})�O�}I���b�Qt5e!�	r��.8�Nbn5�	b<�]��&������c:N�us����F�[��9���ى��"�H�Ŵe�WUbw=�C�Ld�ͥ�g�{h�*&�ځ4���2ܷv�v�{l��$j̆�\l�X�c��j��6��\��I4ڍΖUvK���;�w���b�״jq��]�yz�2x���9!ݯ�p��h�z]�.�Z��JEp����֍��mgV����*N�Ɓus���qi��]�;;H��Z�r��7Lq�+Vlnr�,"U�u�T�ۣ�7��u�:��v�P�S=k[Pn}��8(����v�&p�vҀ�Ck��ԙM���\WM�o��������\���'�5��:N�
�2VQ�����6�T�w����:�z�}~������d� �VT�a6�@���򯙫��\���Q�~�'����1���_���s�� [�7�!RX9���
l@�����Af�*IP�^�r�h9��Gl<aXP���3.��4á�Ns����T�ïy�Y(ʁA�+/ov�~���xYG�����06���������o���_�� x��~��Ȼ�-�9�w���v��R
w�xm&б%H,)�|���¤�T}�4m�{�e��=�;����3|�m6��q����n�����sZ� �-�w�<Ѿ�!_L5��W�wǦJf��M�T�����d�X��D9�<��?~wO��L�Q�i�ɍ��-(�ݴ�P����&�1C��uum֗��y�-t��>a�¦����Ad�+��n2�Q��Ts�h�������<<���ӭw�l� �B�!�|ޠ�k��U�e���l fs�OD
��Y�}��ژ�ءu��U�<�����{賖]n�d0�g�>��V��<�Yc����?�޿w܎h�;i�h�ky_���S������+
{����
�RT�~?�b��_��}�.�V��ߨR�O�u�2 ㍄�v57�H$߶�2K�������{~�c�W����@��p�aL�N�u�UCo՞�Nj� �^ۡDf�z綥͡�A���V�9hq%>�U����另��V͍��� �t���6u{�xI�[$4�h�� �X۳��MZ%u�X�Hɍ���y��FT%!<W�B�m�@�h���-v�	�;-�Sf��YiS��?|T���3���$���No1��\��){|r���7Z�E�h�ifO���IW�q�-j�:B]oA����O���*�[)�(����e�[x�í^wƎ��?�ǻ������_Q���>2�2\ʉq7gL3h�q��V&GW�!3�i�_4�0��T�J�(un�4�9��V��lUϛ^�*��T��6S@��|���MYz��%�FJi�d?�m��;�pv�LpE��f��HAEv��8R�I7�$�A'3���i����>��z��ʠ�����FT%!4
�p�or����;��>3�SA��!뺽�_s�g��t��@2&��^����L�1����l����l�_�m�:�_��lUK�us`$nl��wuש����t�1�k���$�=C�ǫ��l$\�=N�y�V���(�l6�N��]���e��肔7�˺ ���o��Iɲ����n'w�����o�txC1[��󜎩�m���1P�W/�GC�~�6�jH� 8qq�E�`R��9��h|C0B��6�q�}��M0�|w�G��� �/{�����#�ݲ����!����s��D*��}�~�����=�MR"��]D���7�!�-5�R==/��MR�̏GE�������O@.��Lݑ=&J�]�ޖ�/��[��U�"�8��A	�E�4�n:�=U�$w�u�͛��p�:�����9�9�_��/E�vv7��ה�Rǲ緎<��[밽B��e���~��xg�x�-z4���R���-"�նc17UƃĚ//Tոx�����,VS9�A��#���[G �k�yy�ݬ	כ��n�iV��x�ǁ��o���5\jܝ�>u���!x��TnGZ.��՚]l�3	3�$�<��ͬ%�Q�x���m֧�-���H`��NxWPɹ�ݩT����y�s@�9�d�5q���H�pߝ���p�A�����H$�v�I'w�4��nzt� $��ڪ$p�]�aD��l��V���V_l�Y����ҙ�ޭ}�(�%�U����Iv5�U	7��͙�9�l��+ ܦ����?�W�&������ܷ�>$i�3�Fw�f�� �z��vcd��z�۽�_C��C&jȟ7�vK�ܗ�;/�������m���O��دG�x���6�a���F�f�MU��q�i��36�CG��ľ$ۏ�ٔv���A���ۗ2�2�@9�hn*ly�����!=@=R��m��2U�V����ׅ��'�ș�
�U/�ݴ��\Yu~/u��e՜�olY �?�m�T�I ���H���὾՘&�����tXEDLJ���4"���'��g*�}���kM_4��0���S�%��(6#�{B�$��I���BI�t��ƪ����Cx��8�4
ŦA�e�5���#�۽!X-�m *������1Ӆ��bf��/1��z52�W�\�k�Q���y��+E}��?q���'���� �	�����i�����=� ��Nk�'
7	zZ��ĝKM���]Kka�9�Bsz�0���^�W�!����I�w`�r2Gg\�A'6��o�W5���7���M<��D�R����?=��t9�zo�W�E�8�菌+��{FL���A���I���J1&�Q:=��_������ڐܷ@���ɾ�i{�f�#~%,� �Ĳ�L�>��/7������g�ˑ�ؓ U}u@I��4�Mt��G4�ai��i��k���;$qe��э�!�d����6$�08� ��H�e��.�l��ZMvA<0�v�d��ߜ1�+��Kٛ�׺�x�~�z��m_����za�_ �D�9@���*�$���A�Ņ���#�-�|���+���'.&�DL���;ʪ�_ &� @�ݖ/\q�r��s�

�ȵG5�oo]�������h�\t�c�z�-����fQH�Zmn+Q�ӡ=��C�|�}�>� �a6O��a��ߪ	�Z�}F�.��T��oy��>���NE���~B��#SL��ݑ�q(�RE� �"#0����I2T�G��������������]��]ڰ������&��NBÎ#G�=�Mh��{��^۶��oJa]<?��*����+�S�����{�we>�B	5�_� G
��Y���+������t��+�l�u�}�i�=����uܰ����ej�����6ؚ�V|l	ˉ�tN} �����X�߳�A�6�%�{��ʣ��E���\�]��hg�f��Z���+K�5����%t�5�O�qmiѧޗP����߲�eZ��y�������$�h���]�ӌ㣮��s��m'f�{������A�oJ�� ��b�Q�]VcB�Q���'������Mq3�>�ۮ���lt`J�gx�H��[��T.�3]�n+�1x�F��X��oh�P����DM�ƺ��um�D��uwk�K�76�W\�s�#;�g��vY��u���Pw]vu�v�\�7�{���b�p��S7��s{��UZ��{ޠI�)���6
�H������3��^#z$
��MǆH��P��517&Ԩﶈ��T*H�q�F���O�ޔ	#3V��ʮ������H'��T	�\\�p�v[���v�mS�����6�����J���:����fXþ�kfC`��+�~=��/����d%M>�ʠB��q��c�.�[�Q0&���v�4��`.����?�(��)�%�pXş.DG��H?������7��;�-��z��fM�=TH�e�X�I����Q�%ǲ�~�A�j[!�'=�阖ڿ*P����ri�R$����`�ެ�#6��Ry�t�{�%�c��f�:���_z^�L�W��F�K<�`���l�`>���#�W�rP ����3���k}�4q�t�5�|5��8�W�>�F��Q$ݾ&�N�\�u�$UN����oZlE�<�J$ݬ&j�F[�^������Um�zdz\'#�6�:L/f�\Wl�H�s���E�kN[����	��+�B�7���$]�0�8�VUWwm
����tC�-���aX�z��^ggy����:@�+��N��|Οn�0Yj��i0�ty�W�AK� ��U�-������.�౼�5��8�	�,՗<�����������o����f�ı8Bܺ�����x<y�W�0a��ۉ8�� ����O.��wNo�[�Ơl�X���/z�^]����}<�Ix��F'{��<�=�ks�_?)�XM����x��t��"=���3\�=��k[ ��e��Zw���>����/`F�u���
د�X)�O�==�ǝ�ݞ`:���D/�>�����R�3}W��/	��S��n�[�ċ�9�-�a =eB8Gh�;wgWw����B{�EU�W����݇5�ϫ`�sU<q�*��;j���7z�շ=�a���)Z�ׂ�Pn�[Y��S�bK�|%:��_��#8�� �Η$�3�Ra��O!����7��{��h�������S2�3y��\��&|u��zo50N9��'�X�������;L��k�Ō����z�̏ԫҎ��}���y��������[=��j��./Ot���&�4�V5Ό�q���	w�����ٻ݂le{�x�g���s�+c�䝾�� ��	�מ<�d���S����u�;œ�s���������e�=���k0Dczz���p�ݳp���;(j��9J7^�،\��> Bp�Kh���1լ-)m�
�*����q�2�B�z�e��x���e��z�ҊA([�U�#��3&)i�\eLfX�BJ���#xYk#-l��b
��)UG�\�[BD����y������De���B$ @�Y�Ʊ5E���֖�Q�i`�9y [JX^��ӪE	ļ�X[�UBFҖ�u���ȁ����n�cm�4��m�Z����U����X��eN�ll�-�[DS�KLe�]3\���R�
��
(�l�����y�
'��sS}o?$���o�l�>���Ӫ��t^�"	뮨F���ޚ<��Uj�c y�J��Ȕ��F�ֺ"?���J'�"�o�:�r�m�*T��|��U�گL��ĮyZ��F���cvr�<�.�.��n3��
R��V�ɶ#�A׽D��� =�ʤq��w�>3��R*tO`N��S�.�_Kݮz���UQ �S�0]ݕ@.��H�On^�Oe�^I ��ݕ�D~#�} �nƦNws� ���	��P���W��'G�U?���W^80k�G{=>�w;��UC7i�γӊ�� �O�{�;�h���Z]T��T7��aX�����M_OF��H]�e�������}�~��x��M��Ѻ��U�|sw��>�P�Y��nA��U	�z����[�i��CĶ��
D �m۰�4P��M���B�:���7��~|�;U��8��`n� �=�J[_�G��H'��U���>m�$u`�(�ɩ���es������=��}9�3i��N�'��S��x���>��9w^$���P$�n�D1µ���K��#\���͍P�]�7��(�bz孻^�T>=}�P���ƋI��z��es���eo1��>&�uR E��Ru����L\iP���>�:eY�MU6�����VO\�X�u�t���|j��w�c�\�d�Z⟾�����Xq�/X�z�ѥ;\t�]V�2:��۵h����7�63�u�67���Ŭ[��%��[�;Ɨ�� ����k��4Kn���t	V������[�Ec'V�^ݬ�.���uj�Y*�
��52m�0�vqa�񭨩��eSwZ:��]J�b�(��mV���9/X����I��XTōà�"$@����M��ѽ�ǵU�?��(G�����z�W�:v{Ֆ� ��>�]b���h��>$�a>ά��*�� nwR�����U��ș��V�C�#T�A#s6���>;�`�;ӹ�xu{�"�|� ��4�
/�0Sq�}�$�6&v`�\�I?'|�@ou�[�W��Wh޷+�sHi0��`8���v݂���{2� �� ��uF��=�%B���Mn���Z��y��F�����	��#t�v0�����ߟ�É�<���&w1	����Tc{s/Mt!�k��������!��n��uJ���|����o��]Mg��d�~�j8����N��}�u����p��]]Ҥԛ�y2����2&��O��^5a����|��y߾�|��`����:�ۈ�u]Z(�g nBCqw��g[U�#��;S���U{�`�.�U�v
��"����vN���r�x�9T����=�7��k��}hկ2b��#+2xE�m
��jy�i��4Џ���P�u*�:�v��36[��ߊe���6��!���tiE�g��l,;�ci�o��=�� ��~��8A9�pQ f��{VU���O{�T	�3x�m��tWuW�O�<��OkEV�0*�.�=����ڞ���;��z��M�T�7W�j����T<ϭ�^�k�]�{UB�ůg�VG�[vsg�D��8P�^�}��ݪ���;�N]�򣝛�r�����2��ro�8���y����>���5-�N2Cqg?9�z<�0Aί:���UW���v����H�Δ
�
��"�����(���<��%gDf�N������T����U�g�������a��m�$�X%�JLh���,��Fs�z�,m^�´(�)��;�A7��������O/6[k.�;j��{�����g胍՜q�N�kϙ���W0��nУW��*$�iޮ�M%%o��y��i���Ě�p��.×1[�Wwp�F�m
�j�}����IO�v{���Ǧ�f�����t���Z�FX�∭�ϥ���y�����#��=�s��a^ӆ�oY̡.'���h��J����=�2�hcIS� ��#wr�[���\�����_��2��+�֛F���;^���w�� ������V<��w��L���'��~�q�Q(���o
a��C���Z��������2'���TI5x�#{�їSW�g�OuW�o4�lTty���7��?P�3���M ��A>$�FB�w[�q��'�xyP��3k"g3�n� C�{1=�W���9��[�����[0L�2�h��ڌ�^�}W�l�τ|gn:v�wd���r�n��U�@H[�g�l�>�݅�T(77�R�|5
pl�B}] ������;�J��QП>��t��r�9}��`_��=�fj�������cDlf���u��ͺu_�}��}��\��L��6�q�WL�ֶ�K���0�o���<�x(м�׮[�d��^lr��z6�;˺kw`��B�m��0��ֹ)p��=���A4[��kl"��qW"U`mUH��f��n;,�'5h��k�k��:�gk���7+��v����3Γ4�8�78H;��	�pv%���Qu@�1����<�$7�y�ٞ�W���u������w��!U��0��#wh��t�N���Z�m �veR_{���Ż}���n��ͮznێ���>�w���Y^�~쟘f�R�.���.T1�q�ϊxǭ�<ww/tn�o;^� ���/��65�Aݞ�K�rW�-��n�8���@��lS�^��-t�@��9ٵ@�}pC5v㴭{��r�֘�M�8�lZ(9\g'i�^����~~����0�s9�7��3�ΐ���W�:�VNMvz�|v�=D!�kL�a���{��2�ѝ��+���mV/ץ��t�� �Vf�"+}U�k���1/�K�RNy�|��C���H����>�����@��[���$W3q�ת�R���[񑻲�uWז�$b��)Å<�� ;w�����-���c�hs.jy�LD}���A��J�o[M���kk������C��Fn��O�G���:�7K�z�! ���e�`�{���gV�꾐S�$��v3P�v.*�gÌ�`��-f�����>oώ^����>=豠G���D,s��Q���>�v`���c-O�w}ҨP9�Էv>}ѕWG¾�#����<�cӕ]��Q(�G0��Gt1�gc��|=�ZA��/=�=��v!���^���<�O��y�W�݇8���K�\	Hk�4����}��&U͵{��\�����y�������:��DwÙ������)N}`y���vwy_�,�}����G6��F�n:�P��w����/�`��> ��A�ٽ_SܯW�n���ĢL��1����)$[�X�1u��0�˺|���ns�"cG�ݎ�s���v�z�iK�?�wvU Z!/։m��cWOD�7�K���RdP'���
$﷨P ��c�n=�����E����Z�F��]�TI'۽@Q"-������yB߃3��G��J���Dk6?��}OѮ�g�����(�o���zΫ~ Ƈn��n{ŌXw'�H'�{������6�fς��d�05���Fdh�fX�9���|�&�g�B��Y	o�6��+��>�TD�{W)����HfWԍ���؎��+�ck2�� ����Z-�i�39������-)pE3ع�e�̎:O'�ٴ(�������K�gdl]W��$owUP���I�GV
k'ݝ<��V�ښA�6P$|��;�w���C�%m [E� sj��?�P"	 ��=��;|�/P|����_M	ͮ�`��?����ŬY���Ԩ [�C@�ʭ�Y��N�WP������!��j����@����1{1, ���T@��]��F};�:+�d^�S�ٹ"J��j/�R������^y�\N�t�q;��`���W����h
��a'�A��{|��_*	yO��9�<�'7o��nm�=�]�^��|�
��`�R�K�s��z/\dvщ��� �(��L��ܡ�n���ÛiI�G��ܕ���K���z��t�s]!��ǫ7A����!���Cv�m�ߖA=�/O^we��^��]JOK��|)�G?_{e�-߼�w���)m;���5+|6'ȡQ䄯y=�!�[^{
��p��Ȓe�ݓ��]�Ju8����٧�l�6��v�Ξ���m��Q�,�Z�֦�ܞ�
E��OM:��^����y骽�Ϗ���U���`�u�����M�xcŰD\�e�?g���^���:R���:���V�N=$���;-#=�ʎ�����Ei�|��x��6��wGm#����۠���˻m��>��ʺ�e�AI����u!.GDoyqAW��~��*g�t��u��7_:�B�ܓ-g��7��V��\����>+��猃U�[���.��n��	%�m*
]�c�w=o W{ľ�{y2xt�f,���G�.S�/�N�Q3
�0�DE��[B�J[�7-��Z�lAUE��Zʖ�/P��E��� ����!,8���� �\�[*�U�Q����mm�U��B�Kc{��m�L1n8*�����oB�KZpYV�-HJ[(,*ZRP�Bҭ�)Z#3ʨ�2�"�E���F�����孥S2�
��Բ��-R�m������ZfPŵ[m�ʪ��h0Q�m+�W�B��j��E�iXk(�ĶVڬ�h*��up�-j�Ŵ���m+nXbDdQ����AY�C0�
�*7a�hͷYp[q3p!v�P�뭬s���m<(e��Q/3��.�7	c�+�K?��5�����3-�n�WMU�j���RX��"	nո�wF󮳞	����'�3h�<���r�T�����9[/^z_)�]���&i麃m�mY�L�2�b�1!�L��Vu6�4�u�FPb)fB����wP#������,+s��j4�vPa�ή�hŝ{��j :^n�S3���M���0�����T��;�π�]Ƥ�uD9ո��1׍F����
��ю#2�IL��h0�շ!��V�p�<��u�+jڳ��
ލ�і�8����c�=]�V�ZJю�(qv��Xr�t�E�"��kp�Ԛp�!V����5 �uWma��u�����	�?[;}�^��dt]�k�J��[�3�� 4¶6���V4˝`7,����Z"2�V"%��A,]r�C��݃�V��ǌ�dǞ��[����c%����Gk�̀�Hn�����K�ւ�q��� ܲq�u]�D1L��-�^<�x�Vw[.�	fe�-�MaAƬ�b����t�`�cHb_B�%Ե�̧Em�0X�s0x��v�v^v�2Gkn6�i�x�y�����9|�H���.��A-�v�<��Œ�bR6$I�ޡm�H8N�;(�>}��W�.+U;�u�j�k��&�\7F(n՞��gMp��I/=u��tC��l�/Ls���%�NöF6;Mh����>ms�:�ָԃr�fP����t�_\W�9V��8hn9�u�(�<�� ��(v�]f�s���`cqŨ��9�8��dE
�tv9uÕ�ۺ���v�c��׆�������}Tj0%�����\v���6칓(,�+9�q���v1\-uqF�U�;]Ud"6@5��1�Ę4�Bu��]�s�m���"��I��U)b#!?�~_�/�B����t�M⦠ ��G��;8��ίR^����b�㮓*�$琮��u�J7f�wcT���_^'�c���_P�x��e0����h ��t|d����S&�r���SA�������&`��5��U�[�zɪ�z��ʯ�v�ݩ�=���?u>�h��)�r�t�`9��Gٶ��v8$����U I �wU7}��0��k�D($0$�.����"eu��[�s,��b_�`y�@��},A���|��_=d���ZA*w���}uD�g��ZQ�vvN�{���`�Zn�zz��!n�S^�A�پ�������2���I�4��W��ΰQ�q׍�|Nh���ѹ<����t�!g�ߪ�x�%�3g���'�7�>�U~$�ڠ@>�odt�6� A��T~�o:JU��d�-��6\�ڏ�m�������J��j���I����ǝ�G�t4Y;^ ��fJ ��U@�[������x[��J��킉��!�?�Χ�����l�p8�{o3�<TCI�Ro����ߺA�9��*��ww�|I5}>C����W����αL���bƩ�,�޻C�˝�����@������?9�Fwwi�.G��ۻ�ꯪ�X/������߻_�7�I�Rʱ��{շϟ�K}�x_v��������\]�N�]b�l_��ˇ}�nb7��F^m����>��x�5V����ܹ�{#�3����}YJ��l	�t���iw˟�DA��a��nmlL����|F�L��_ w��w\�K�no���בo�Y�t�N����&�<\j����Q8����q&�2qݪ��@���{����L>�}a��}R�W���c���}�[�TDm�עT�ʠ�Ԩ@��H{�u��s}�{��L��0%Ђd0Q]�@���u� 7�L>�dU�<o�0F�\���y{��2�n짼�]D_������Y�T��i={�ݛ��>.��?G�;����܏�7fS�][���-V:Т������K3l�ڢ8��r|r�yo�t9̡D���B��<�K۔�_]*@���R��r�g���Sz"b)I��(AD���U;fy����i�WA����>*G᩾'�A���?��T�'�v�v��ne� Z��v ���㺩���k�/.��q�*��/�
#�z|�hIf����bz\1A�kv�P$��D�L�����I�����ꣁ�	Y"�gǖ�]�3|�#)�T!f���=lOz{�f���ʪ$
g1���n�[��~/��y�/�����wJ��y�	��^���~Wߎo���F�ⶰ��>�4�3�ܲz����5����;�T�Y�L��^��D�ժ��0L!�l	R+����z��6qd�qʉYNt�� �+c�m�r�a�7n�X�=��];6`�6n��>M�F�1#4%Ұ����2Dn�[S��,)�Pn���B\�b��hX�s3�͡�;]6b�&y�ڷ��Vb.��	��Ͷyzΰ�N��;6]�8�^8�Πw%�c�e6�D���\���~��@��Gl��$ݛ_W����e�<��u�W�������s�o��[8"�y{_U� ��������y����F�v;_�JA�'��.��N��g_]�$�oAD�o��?qO�(!r�wU'o3���^D�m����	��� �u��Yy2"� :��P�J��d�㣲 ;vڒ��tւo�T� Jrp`����W�3_U����F݀i�1ݥ�ga�C�ۯT�@�a�O�-FۂL�Z�"�q3�#s�>E�֠@�ovU>s��J�_R�S�|+����Oц��8��(QW�����RtU��o���;�'�ݍ`�x�%V������˲\�S���ttR����~)�|�NFy����>��HgN�*u}W�5�����!��lN@��t	�*��}������v:�����%DCk��~ۨ�^��v���z��v��ps<�4�k�	S�E��b�.�[�_W�=�T{��}�w~1�"��P�;��
�>y��7��c��	ay��={@"KLV���ca�j�Ds$���:cZ�]�����F^'��^�I�vU ��r���K�����Q1����\�oƻޔ	s���(�8�䱄�/�I�#���2��w�e|OǾ4.�͝�}�IIs�N�L.��Vٸx���~�6ì�FS���w�Bwe7/7�f	囜����5O�=
Jy��I��U|H$��U/�z(�EI,%�$5���z���^�H��t�즭��%���]i�_���v�)���wj�;i��{W�	)��Q���W����w]Syx�	6���I�ĺ�s���Omq�&�_3�^����_������#��/n<� ��@|vE��y��{k�s����B���l�!���M������+��;�{� -��W���,�����=�h�<��	N&�%�0��O���=�;}3S��#�����T3NȚb!��s:�kL����� p�;�9�My�V{3_J��=��U�S=�')}鯥;�v*S�a<r1m�izF���a�B����+N]�Y߸�T)ٽ��p���	�@H��j���
�]N�@p�w�*�3!�a9�q�XVA�	�^y��t������;qu1�9F6T4�>_�JAOgQ#O[R }��7ו9V���Tx����($f.��W���ҩ[�z(�N��	���WĂO�}�&��XaP��F\8j�9��;q���gTo��}�$���3�ҁ3�3��
qGv^�ɏ&���LG�u���UA�މogXэ��W"O���ɔ(��mS�>��>����N�A�ޡ@���T�	�v�(��{cs�J�Ȝ��B�Oi��wTR�ڑ�R���N��̙_r�"�d��E/xf�m#DSb"�04�G`�Kq��!αeڄƖ�/6ɪ�c�ŷlWb��f�[��2��vq.�!�'�/=�ng�sqc�R�m�:�2� hC b�����j8[M�YV��$�y����\�[�B�[��)1�즺�ʹ�Wl�k�$�eA��K�F7 �&��ekg�t�uJ�kX���Z������Թd6��'�.��@#��"\�����mJ����{0`���<��|��R�t�����u�U ���EԮ�R�PSN@���\���TI ��RT GLZ�����5�b�/�*��������L��((/��=���=����: ����/Խ��B�uPT�I�MDK�wϩP���W�:=�ޅ���v{���\W �I������A
C�m9p>zO9�GV��W3[�]m'S�����I#�rmQ$��mQ�j�@]տn�I�D�o۲��}���@��rZ��c'~���_��,Y�����'7W?o5[�k�}�Ђ�_������.=)u�C��>����\�I�l����ἅu[��^x���x��S)�����FHΙ���j�«W�#{z�#�М>5k
	�˾}U�p��㾵{��l��>U�	'��E�zwكۃ�A��t:��" �E/c$�vzQ��^�'_�$=�U�?uV�H9��E}i�~�2�aBT@���6R]-�ih�[�5���}������'��t�6k#$�~��UԞ�������>'Wzӌ5>�GBy�|UOޞ�������ed&��Tǳ�*��Eپ�dRB��r(	����?/�t����֟d������C8󻷲�/)7����/C���kͳ�G�Ip1�`fP����k/��*6�d�y>�#��'�XI�s��K�d���Y|Kvy������.��c�n��f-hfv=Gn�'��e�^L�XٌLݦv��(�iW�׺=�4�X�s~�y���]�>n��ez��P`��k�K����W�6*k��/������]C6�%RQ�VY;����tC=��k�؟	ﻶ���tO<��䂞��r%j�����TE����&n2����=_tw}�I�+��#�Pfn�݂������5�Qc�¿.st^�qn�}����y��z0�b罺B�C/�(Yz<}������}�K��ݨ�wxըff�*t��o:Y��uՋ�]��ǳơe�7�!��Z�1��gz`�^��)
j9^�=W�(=��L;�1[�L7�S�t�ښ�{�c�7Nbw�=�m$�I�V�E��"��Z���<�s�r�&�k�97���%�h�=�=:��?OU/ ���N�"���զz�.���QM�,O���ח3�ߚ��Cŉ�7�)����g���xk���A_)�]�w���C궵�JU[10��zXTZY��k-H��-�B����Fܹ����R��fZ�!b�iUKF�H�hQR�T11��E�*�e
�(��֕i`�U���kU+�fdS[U��m��f\+l�s0��cV8�уj�JT+\�r��ִb2�S.4�6ʱ�DW-���J��km��i+��X���&�b1�-UƊ���1.5cV�C-�E��E����DAĹm��Rګ�J��a�\�(ҋ%e���Z��2[�X��`�
�F"��
1E�ԕ���H�a�T�L
�P�P�4�E������Qa�!�rƩ%N�o`Y [ֈ�QX
c�&ґeUT-�T�P_~����]�t,S�y��&_
�Ja���ҏ��^dB�B��U�'�{�UE��QӔ�Ā��	�HY.�g�T�����WT�R�ի�(�C�a���T��R���|D3�L[��<j��<\!����-���ı�-~�Ͽ��1�E��0������ ^���w#gs&U��8o���:��@�ˆC	Iƥ�����:ب�W�>:��|�񽷵�n���Z2&��H�?A���vТA��,�3�dm��#{-�$��R��=�(d�I*�ơ�V�"��(���ު�'sŨ�¶�ٝ�Y���'��9g�����3ϲ�
�y]w'v�w���N�Zg;��pŔ�˰Z|?u:A����J�r�=U@!����~�v�W�(O���L�����y�U��?�B	ȑ0�ӂz|�%����a�Z��:����]�Jm�oݏ��|o��Pw<4K�/t�N��$|��c�Tv�Q�C�mR"CS㋼���׻��a�o�#ټ�!�p�Lȑ�wN��&r9E�`��B�3�" �,����� B��j�'s�@ofA.&_ͷ4���P������ʪ ���9�t���vL�>���-£whن���谖���̆ﱩ]N�Rs�H%����3z_��fY�^<M3/�u��7r1[�k�yVV�;Z�Άw���awX�0t?��/�#�j�:ݶP�0�pY��%����1\yt�f�.��䣴eN{��,�qv�Uc�+.��Eᎄao�uƁ����16[�еΆr�͸��8�Á�nmW���v��dK�S:�i��L
],�jtn�u�[Y���p0t˳i�. ��X����h�9^V��r{7�[�9�@\��6��,�!NH�1��<w��L5�~T�tp�{���3[�Fe����lpȕ������ZŶ���O��DI�L���TI{
o/���{T.S왊�61����(B3:�N�[��T_f|H$U�0�޹E>�pHJ�*ι��U���y�f����@�m� 3}�u��z��h2�F����n}$��o2��A��]_Oz��R64�@������9�c���YQ����>�ә�m�#�s���[D����eqf31��a7�>C��
q)'���@9�r� ��ު*�a��UŚw���Di����A���cN]\ڧD��;�-�+祄rv��h�^��E}��s�H��*�&=0�M�P��{��{h+D��� W�ڠ3{�R��c��s�D�a���f.�mU
$﷪��m����w]*@���������>#c�٘ߟ�e'{�| ��s� �xM��rT�P&�]QOܖ� A��Y}:���<�q�j��^:.�:f�W�K|a��{����"Y,2���%��t�]\GJmbh�.ڌ�f�R6��H�����z� ����2�{���׵H��Y~&�S�I(bO���/ח.v� /7��w?��R�O���T����0���U��� $f
�#k��>�k*~���6Ty�vzM5-���,��s�6:�؊���e������E����|7�o%�k�T�Á��I�S�#%��2U���pXH�ʠOтa��]m�;��.o�s�Z��IND��_"=?�����mK��;���n=��c�@��R��>�0��kg�J9�:	�]�Ɩ���ńǌb�ųi�2��|���94�(�;Q����k� ��T"~/���U�����%#j}$�.��:��첧�H�pb;��R3.ί�||�+,h��$�RJ��5" �{��|A���{�5a�ȳ��	��s���/B�e��|y�W��H��7������Ϩ�wCUf	[�i�&��1�J_���U4{��㋤z�}�׶̛=��ߵF2Ws������1#�w�\H�|D	�7��J.�uP�/w�W���� �0o��H��A�~��P���$67A1 8Bn6��@���&��YVT��L�@�c�9�������s��J�A����ێ�$�۪$�9`���]���Q����WzeZ��O�.�@=��PH�
=�MM�3�Y���r?�nju�W���w�P���5�����"��� ���X���%�6�͘k�������_7@g�TH2�޿z�;A��vuAX#G|#��u�U���~������x	��H>7}_W��Z�3�FF���t���釨˞-?q���A�Zļ���*�r"�_g]��l��G�zVu6�n������`�O�$HI)�.�|\�5�۷NЧ7m��v�	���td�tSֺ��M0�X��t���lu�.0��ֹ)�:Ķ�`6vn.&��&��k!p�SOh��٬WC���m.�! �t	m4k7]�ל�1.�d+��+�. �5�.#\�A�i��R�)�v4:�qvgrPs;'8\��P�o�r1�=�G�46�c{�UP/���#��p�G�G�����k�"sw�����&�x#��+7��q�����{���p��+qq�ީ~���� �2�Ө
?�Y��]�z�=Q��$}��Q�2.�M@��8���DGSa��ڠA�\a ���f���{չ��[�U�4_	
q�%X+��ޔU�O\ubV�Uv�	��y�5�R�M6�����N��pt�I���ΫuWl�4��D>|�������"F�zQ���W�i\�q�j�! ]S�qj��jp1��>��C��~�gG��?����H���U�oɰ[����F�O4����W͉W4%�	ف�j��Ͳ��0J��_�����W���ӟ�n���(١�ƶ"I�g��w��':�Y���A#;�TJ���	�,-}����xo^�bu��
��@���R�Q�$ЄןOϞ<I�>q�O&U	Ggz��WWl`���eR>��W��jh��;T��^� ��L&�)J&��d�lr,�M�A��p�X��4K�m�2'� v�:����>P�o�]I0ň�X�P�DĮ�7��Z<�����ʡ�z
p���L�����#��d�ު���u%H%�}^��˪�W[�T%̳F������/v���w!�a��p?f�H���o!��1z�. �	���� �w;�Q���f���#
�B�s��O�T�I��k���r�u�IN��%[W��B��vO>�@#
��b�!�I�\�A>�tM��3�W�S�����i�g�J�n]<r>au�4���p��Z���ϟ$�s�|��Q$��l�E��w���鵝����u��_H�.a�vA�����im�-��#{ޥAq] s���+f�ʐ��a3��=�9K�46�X����A7��_t��U��^�f*�uU;u��qcwH�z�j�9KL$�����N��He��8c��
�;����xj���r��w����{j�cf���)�.�9b���n~��XXN$�1F�/``���J+�K4v���O��,��Goz�>=۹������!,�c-�!����v��ƔW��<���{E
%�x��t_���{���"%z�����V��pY:�(H|���8�\��B�?_L�ﲐ�C��T+�[Q���umX��f�RK�Qȡ?��H|gO���Y��G��0@�ݕ@�XyA3��+�V]�za��3w$�����7w�E{��1�)4:�V�f.���TA�z���Š�;a371����~v�b�,KVA_[��.ݯ��dǗ�����Μ1F��מ�*���}�����2x?v����7����
�����&�������9K���tlƌ��L��èP��'9>{�}�
x�4�����o��Zu�>���[��6n�f���{�;���.�&���s7���vW�Ǐƃ�|� �s�c�})�׆�?���2�!����ޡ]��6)T�w�VJ�y��^K�׳�׭�%�o���ؼ�F�{&#Gy���{��u�ԭ�� ��׌]�����̌�z�V�A�)��ߠw�rW��}Od�o��mM����ʸ������l?V=�8�^���})�"�'�3p�Y�%�m[�w/	)��h����X�6�]/78�y�������nz-�����86� �б�4�ڽ݊@ƖwR���s��U���7����n
��	�r������P�8�mW�Nn%�v[C6$p?K�x&�a6��s�`D��e	�����M�5��|G��b:-&L�eޝ�f����'���c�M������)>�� �ߪ(�'��{�X�Q�mZY�Y��N�f���z��+%���5u�ǰ�QN%G���!�����G�q��1E���(
�l�*i�e#JQVKi(�JҥF�R��$Z�bT%m�V�dX[eK�J��+%q��P�DX��kj-L��!X���8*�HT��Ku�E��
�*�al�%��R�f2�b�AVT*E��W-P�)�2�Q2�)�
��L��`e��X�J"�PĊ�QLq�ʂ%B�R���[q��(�U1�kX"
��DӍAd��X���%f�h�.5	��,�ĩXۈj�1��5�\�#XT*�2șIRE���(D��IP��h
��*"1LkQd�IS�U�T��P��6[%�������Z�MM� �g���(�4�:��x�u��2�-Y�u�f\�5K'\:z�+1���'lU*�	�z�(r3v��9eG���N+���=���:7s�έ�Tۘ:5�n�v\���xt�0۱5@ t�6A���Q�,p�ѳ��vڻ���s]e%ne��v�Ԯ�a:M�WK��S�nذ;q�v7]�.=�����&��MC�]bٍ4�Y�3sջ�ugoNm��u�X�M��ɸ�ug\v���o�k@n�y��9�k�v���f��67P�UE)Al�3Ձ���:1��m�����c8�pյ�m�|��v��m�yv�&{J���e1�:p�/Q��.��m��rzy�&c�X�lu'k����d�S��+w �M[gH�<��K��Y-&����ZM���EWb�5H%ɠ�Bk	Sm��Hv�SN��{m\^�{w]Δ�*s��\���k:X����X{!�z�Gv����1�[x)�R�Љ5� ĈMn*�:�P�������ns�xl�{\`��R��b�2FVc�]��k�CL�0��ek-�R��k���p0����4��
�,�ƹ�ֵRp�5c��8��t5e]J�q:��3⹷�y�
��+{t{]H�]뵭�Wvb�r�şc@v	u�c��ݼ�W$�ڹ�\b[�bC�۞�����Lӛ�L;q�*E���U�э�v��Ԝ���v�ǆ�����*�����sr�NM��\�),�=#�s<���lu�q�Dv��n��y8���}���X�unQ%��se��L���m+�Fz�-���tp۴\�\�p�K�ܝ�e����M*f�ǁM,�%�vNK���)�]�wV�����M�3,Ķh�SR��y��)�tٻ2�x�j�oJ��LU����Q��+�7c<�p�p��&�J#��ǻ�|��E?��H��Y��� }��TFhe9D�t�;��=��D��%��)�/gW�N�F�z3Zo�Oݝ�F{z
49J��X�o<��@^w�'�8�K�x�A�v�e�.Jڰ�}q;;@^oP~�>�@\jIv
/2r��m������A۽J�\vG>^�k���+S� "G.�ާ@i��rsw��UuUA��(f�C�V�`ͭɝ�`T��\#���q��t�m����g��T�WK��~�[�����������/���
5)��핡�8���4p����8�+=�"��o}�Ld/k5�F�fd���0ik���$�w���(����I-^U�6] ��.7�7^>�A~΂�6zЀU�j>�O��]
\5��"}΅�ӓ�A����W���P?=HE��p)�:o���h#r��^ '�ԨB�T'�/we.o�vd�A��U=����RK�Qx�=��Z��+�c�W�w�?�����ta$��ުjb�u��M`���2�av��Ʋ�i��d�{��$�m�/�N#�Q�����*���Q�و�s}T�ݚA��3�(a����F����N3.]� �顇���t���2!�[X�{������d���f~ƫ�Gx��B��{)��W+�y}�vǋYN�̫���t�+����u��R�՞�=c�k�V����Q��S�Ѯ�.���O��h��H�!�t
e��Aޤ5R�ݍP�ލ�;T ^��Asp)�4� �?�ګh��E+���A@�ݽ@U��ӵ��}�z��� es�L&-�	���wד�m��8lu�4������4@[jI�(�H;��_���QC�/m�Yk���F�DPM�������q��WfU #{�J�{b�?wK��Z���E���2U�UU	=�TH���^^r�~'�ު$���hI���da�<2���}ـ�w��/��P&�R���=�Y��	�5m�U+~[�����`�=�[W�����ޭީO�:���Y�S:�#y���3��p�؊Ga.�>9Q�u$*�<�%�?�گ��Ԃ��n���-�N�T;v�g��Q��(&ٔ�n�I��:a����}�����.\��U|;��@ ���R�����}�_Q�ު���8@�nIVQy�Z����{7�I�nЯ�7F鳝�\��{�5k϶���"�mɿ�B�%m/v^h�;z�!���ya&��2_t���+Tٝ�Nɂ��9�LovT�z�=�[ WU���v�%�D�s"������H^����å	�URO���vU#�Wvt���Yo�ϼǹ W��T5lK��H�#5gn��j�p�A3�x����&�rww��o���"p�>
$'��!��-	�wn��`V�8���35TiH�3��U�����n)��x�@[��8���:w6��ݑ��� �a�m��9�45����7$Gm��5v2�Z��7;�D����h�K�k�?I���8��=a�W5��):�)rV�Z�p���}_]��@��sX����~}������S���k�LpH;��G�����Xsz�^�W�l��l�r>q�J{j����g���*�����>4��yg1N�G�,��06ے]��8A=��@��ɾ�Zop�O?�'{�T	5�XyA6�{��SYy~���p	=��D�����mnd_o�ނ��o�P�%n�3����
�{:�L�b=i��nc� �ު������B2�Љ.���RX�t�ZA� ���Xv��k9��������LԜn�h>�����u����}�J�g�����X� ؊G`��}����>�IVT.���m��m���w�08=ծ3�^^��[e�[F}�NY���]�����eȸY���iJ^=� �c���M��9E�t{�V�nB��8�ʢA �f�E{e_y[�P�}�U��v�aٰ533-��&6c��{��]X��=�J�}}4>��!�̀��ڠF���PM���z(�dB������U #7z��_M�U(fZǽ�!y��R4Z�+V�v��U�ǰstr1�<^�TL�1�����!^�W�I&���Ou�W�>��ޕ�ͨ\pG��9�@�8O�dw�������ww���(`���̧��^�F/Ep!��R:�SޔO�تA
��G;B���νyY���)�gGԳ�9Mo��[�n2�ء�<�m�$;�n�N �e�Β.�^^|/�V�z+�`ý�U�tD������:o��a[��9���&���}+6��ܡv�U�w�4�i�.�k �v�Q�7�x��@�]ү�2h`{���K���л�L���\��_"�L�lCpq�}��n��4��I��9ꌰ�rq���	9����I?n�U|^O(�%�Ϫ�nM'��)�,�w�*�����qx�K�D/ʌ�ʤ ��-]�z{��j�l�-9rܜ��bh��t�^6�j�QWK��4oΌ$7��@��r��؊Gv[�ow�vy�8�� ���؏ă��� ;����V>�1�k���a��t1Ԛ�����֏'���z����>�E~�<������'�*��y延�{ב�-�[��?W��5��n2��8����vlGcv���o=�@�I�Ρ[[vƿ����Ք�d�]��qԉ&���)7�Ơ�d�7��rm�ӎ{�k����c���Q�L����Ϣ���}�ޡC!o�2�m�@�UUg�w�u�2��@���
���B�_e����)<-B�nd�]_�y�*�[��@���t��Y�{ު{����D�덆㑚9E̠����&C�wvQ���*/���>�^�Pu�U|t���%L��";��lS��kG���T�����F|}�p>]kH$�-�nnʿj����G�yޓ �O=���kW� j�]وm������a���|���1ˣ�.HT�6��l��Y_�wA���t�N8��c�`+�)5���E��	tr��׷7����Omc�k[������v7p4=,���ɍs�7Ts&�;7�q�d�ˎ*s�jo[0oLیOq��3�N825��].ug�>��y�34&!��K�Gc36�-ez�ΰ5�n�tZꭵ�����G$��˟�L��|	Gv��@�CG�����Wo��U��7�����w���i�.�k"'+����o���d���_:0���V~�ۃr����XM�t��V�P�����������ު@_M���[s$����T+�%�y�@�+�P�M>�e'{� '�*����Bq���L�����(3>��3�u�A�T~��ꣿ��=���{�AM���8V�v�m��[$;;[� qvM=y��bʾ}��!�oʢ����z��t)9�uW�u�c�Rb2��8��W����;�1����5�vv/*"=�2��o=��7���J�p�8T/f�K�R��mZ5VX���G��hL;{�_��\����r�Ͻ�-m2ӎX)g�#{}|I��}w՚:�on� �*3�3{ҁ�Jϛ���r����O�,ϡיT	;��rh��kZ�}5,i0�B���$�����=�*wk��I#�}@ogmOq�::gb)]}j����GU�Ǝ82iv�XU���ԉ�z����Krw��7� ���@��o5g�Ο�����H&�ު'C�Bl�����[ޤ�FWQ=�]��b� H��Q�ޥ_v�M］4�M;�N��7�+�;ٵ��/��p~��~����R�U�F�)�˃}X�dm����)[��#8�GYi#�R�K��;��$�v�V��m]�;����&�~�U������/i�$�Y��6L���|��������+�c
��i�����ux����1���7j tw���Y=�>�o�ޛڭ'·�3^nn}�y8n�����,V��qzBƫ"L���:�N���{�X1��/4O��ޱ$�+�;EF������z�v;K��T����h:�v�,��7.�#�c\�
o{݋��5�c�C�^�:���2�[zv��R�cp5�6�q��Ls�ɑ��]X���ۍ��i~������~B��W����۵l�������7���Rʱ�ovϞ�l�n?JV�b+5n�n��.ʊ�:�#	R��Y|=~{��s7��� �-�l�˛��^дr�Z�=��X�2��۲�j�S5�;�L�k��a�;Ϸ{�]0i	�_����e������vG�>鹱8O�����j��x>�����,�����,K��P(��J!��qҫ�����Ϋ=�'_)�A�V�)uSVh����a��׽\`�x�ދ��cFԣ�$�k�q�W�v��[��ME�<��Z5��X��2e�����A`�!YbԈ�,�-b��eE,d*)��b��be*J�F"!r�"���ۈ�*fP��H��2T!�C�n+�kJԮ& ���`(
bUV�q�eb��	\f8щhT�E"��bVcQI�Z��*QU�3V�Lf �Yb�Qb�t�PXMZ�]1Kg)�[$�6qZ��g�Xc��Y4��"�VH�H�b�J7T�-��S�,��J�jE@Y��Fb)+4�M0++,T�eB��U�
��C���$Rڈ!Z�)R�`���l��b\�������\a�j�UHT� �(��Bĭb�2�cRi	QI1����㿽�[T��}��Ͻ�X���R��Y�@�ݷ(�ު�B��qKR��U|WqfnA�'���Q��`�U�$�ݻU��ц3c�؇����)��$k!n��pQGyGsk��T�=N�>����2#|���@^�U|+�oU_jyj���˪D�{�j�g~�`(8����R x׺)u�T� �ު�(hZ�<({˳}�E�����AI�����D	�ӑ쾓�(��uP?�DA��i���7.H�yr�@���*,顡ݕd�$^�$��K4�#��{حO����\����i_�h��iQxm�`�#c���WV.�琱`��<;�q[� �U}��ͦZq�,>�����M=Y�y�}���F������GWԹG��x=�y�S2���3cA��h�'�F����;-d{7}��!���ې{�AǹTD�ޔ��G\ ��}Ό����E�A�ޖ�=>ȍ�W.�R�[�C [ݕA��I�K��P6$Qϳ��D��_D����?GN:� ����/���x>�,��FH���ه_����%��@�{r���yDN���+���Έ��Ɯe��R:o2��7�j�6,�5�>|D�摒۹��~#ː�N1�Tȏfm�e_T<���'��5�{��:��t�ntak���9�V+���0^c�ЩJk�궈@��j��(�[��o<w����'G1��-۫u�9��y객N��G �Z,ḙ���P�<r���2�Sk�qٽ�z楎1�cN�h��u�V[qn\�[dS��t��BL=���n_������h[XK�{V[Cغz�s�]�A	�vai�e1�BGn7+{v#��ݭ�]\U�������Ú]���{$���sy�_W<"z��@���	�%�R���u�3=��6<�ەB��H3���Q^�\C��ԋ�6��yҪ�׻҈�c)�x7����۾� �3���50؆G=3�ԏ��Y�!�⯶Q$�ݻTA�֕kSg�X꽞'��q�6R.C`��N��Um}}sj�!fw���}?�]1X��T��0n�$-A�E�k�Ǝ����p��n{0}���syԑ�������ƅN�2�s=�+�A'���P�E�$���A��E��=�1�]��z�����:�zne��R�����mѻW���a>]�նZ2O��˫�{��,
��>��HE�����z�j'�ۢ��Ȃے�M��Fr�� �k�cmjB��� ���+h�؂[s2���:����J��Ϫ�
�lh{�YX,�}H�ި�ZxXi�\px��3��3�Y��92k] /tؙ��k��]�R���h(#eH�K�_]B����_O�k��JH��l�x��6JC_�y��'R���t��ڏ^okω��T���C��Ti9�R:	�U|H;\c꒙�&^��?5m(A���@q�,����"S2��<^/9�&%�vI:Ԁ�w�Єfl\B����F����y.�H'�r����]�{J�2����u���ޘ�L�pcN����{�����>$�����~b����rQ��Y2�dNn���$�y$������;Y5�=�>'`5�!9l9w�*�	��oU������`��-}>��UNvu
��G6����%�J%���f�ݖ��-Kf��J;%#�l������Ɇ���9������TMOf�1yg/R�f�|	�z�%!�1>�UJ�����>����>woUl��X�E��5�%P���H�>ʢH�͂���{�ּ�a'V{r��A$��*��{��#E�$�Yy�Q$��۫��I!�yU�K��t��.�{�� ZA�o7����K�w��5lq��"�����	�=�kߺ�@��I	�on=���0?����'��٧��77D��5�O���O� �ۜ�$��T��R������#�7�ʌq�c�	�B�Q�7i�9�*���}����ӳJ�����r��ZI/����I$��wJ����:r��=���(-馩)���a�!q�g9H���y3��=2�v���	 ���+���TA!��Z�s�y�xt2�ě%!7it|e|�	f/J �/LdgU����"N��T��%|�H�c��R�褩���#ۣ׫n�����h$��ԉ����x�Œc9��H�xa�/��#E�$�)U|�	$��*�t�a��uO:� ��VJ5I$�W���An�]��^ap����}�?�����S���=��K�,�iyV���p�x�K�N��g�Ă�������?��K`�(e�Uu�*xN��E����{t8]�<e��t�݉�ڞ�@�:4��;f�'��.Z�ζ�XĚ���;�	�/:����Z\��6I�ܗ�MZ5���j�t���\ީ�a�S�7`��8��Pж�gs뫍�U26�n�ң�'���[#�5}��'>���c�6�n����Q��}��3���Q/\��|�9��I�{*�*���{+5#�~7H���ԉ������Ò�-�$����3���k��v�Y$${{*��6��t�aϫ�Q��lC#���H$NgeQ&��\/8t�9�$���S$��,�ˣ})Rؓd�$F�-S��D�țJ���4���&�>[˓;�}^�t�
I]t�$2�P�'�Ir�Nn�	$��i��.��]�,I
W��$��D�H�o*���x[�ϒ��kŻ$qaS��0����Bˋ4�Jm]v��!������i�㞜��U	 ���X��Iyo)A!��.����tɤ���]�� p(nTħ:2��#}���xxg�^��;���ve�r;�O���%e���>�:�C#�T=��c��[����ѩ4D�_%y�U$�>�ƾ�R]�;�z�+�����R�܍6�k6��Z_$�Kq�A#�x�6��$�=ݕv�I|�'�5KT���
����_z����=�O$N箮�($�d�TA$-u��AƈÛ�K�uݭ��`�$F�\�/�Iaˌ���:r�o	Y}�w�H$�ݜj�_$�uӠ�����J�d�=�T29(0�R��6�Q{k<뮵�sq��z��j*��"2}�~�p�JK���k&�߂����N����������ƩW�5�F�N9R�3*������wQQLʕuD�I{&���+�]t�$�L����k��8K�@�r����M%��P�$N���\J��2���؂�=�O[�{����ɿd��J���[`���򈹹G/0�o�e8���j��'���_R$�]t�%����l9,�J��ve�[�k-Bi-;q��$��w���c�7(8�䰍���PЛ�&���,��$�{�Z-q�Z��0�۷0�uR�$�O���$�we��$码�E��a 4��Hl8Çڍp5��6f�A��s�I�����I$×(D�%ov]���7M�K�
E$�uӤ��=FO�������IJ��_�{��$�Hr�Ӡ�H�vU�$�a�٪��������:*>Էt�Z�����]ە`ZI$���N=�i
��I.Yt�$�[��v���	p8nT��Ue�Ł��L�Fi"}�ʫI$Og5���V�URC,U�#�y�D:]�(WR:A�P
q�Ī���������]�㳤�xs�4Z���R���lI,�UU	}�R�3�a�P�IUt��Iwv]�+��ns�F�����y����B�lr@VPq��åg��㡱G&HV�-b-���,=T�$�^�ʻH$�=���
J����{)�D��ʱimRU���FH��E�9A!݂�l�I$�s.��D�s��};�����fz)oC���'�\����v�I�fӤH%��\u����4K��tI6<�
����E�.Z�e;�ˁjD�VՋD��Ǽ��A%���cwҺp�W��H/n]ص�����)�����$��_.�:��>\��uU�J�k�D�Keտ�y��?_�
�����������Z/�!	$?���Rz@�$��j��#gA��6
�x���=_��h�z&�5�	�]$������̚��lX��2v��	��;H_�!��`�?��W��Y/���q BHh�'�'�_��7��~{��� ~���8�D�ԛ6�B?`D3E�?�y�t��A�8a�R����ܝ���;09�6﹠��!I!�؇��?��g�~�=��	N�?|��$���2v@$$����L?�?g��_ȇ����O�t���?�������~��y������$i���@�$��?�!�W�8�?������?�d0�?|��А�`Ju�w���>��QM���Z�-��:�!������� ���?���W@�L��'��R!$�x~{,�$������c��D��$����C�I=J�6K0�����p07������˄����?�@�$����'B*�O�:��	�����7��G���n��?��I��A���~r�?I�m��6�Y��
���ݏ�:��?/�FRB�CĖF|d��C�:?�������:4�r~a��L'�,����������o�~�l'�C�����g�I��_����g�?��C���D?g�AC�������l<?�����
2�~A	!$�	��R!$��C�d�xA=g�Пűi�`��(~4I����(H~F�?�����@~�D$��?��!�c�~Q{$$���,�'`$��?`u&�����I�ejJ��	�P��uԳ� $Ė��v�h�`/�|���!I!��������ӄ����BI@�3�I?��!�O���?�$�C�O�?������2|��p������_��O��G���D0C�����&��!3����5���!���R!$��?��7���� "�yJ@?��������I!d��_����@�@=�8���?�!���ȇ�o�<�w fA?��SC	���O�@��x�?����A���>���?����̇d��5���ˢ!$�~��C��P���~��G򿿭�<�;
'������,?k
!�)����������d�����BI�B2O�200��d=BC���o�?I��������O�I?H$��u���:�=$�07�f@��͝H~PX�!��2�ˇ����;���ܑN$9ʻ 