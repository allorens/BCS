BZh91AY&SY�^���@_�@q����� ����bH��                @ J/�F�Lj�4������kFM��V����[
0F�b�Z�6����,��5cm��jm&���(� �*�B�*UII%�Cv
T��T��U�f�kZR�Z���SZUM�mZ���֥�h�ګ��Me��[iPiL�mfWUy����o��j�[p 'v+mZ�6� 'vmf�V� �Ga��p ;]�j���XmX����l�4$�����Z�&�ѵ��kca��,�� ��+ǡR�		
UABTy%$�  4\Ɓ�>}*�}q�jV�;����m�]AIR�S��j�G77ۻt����ږ�$ճY���=��v�9��4
����ZI]�V�2�|}I ��mF�����ں�R�v�޳�׶���Jxwu�Mn� Ӽ���hJ�S�o{��ZrFy�g���Ԫ�o}�ԔR��o���
t�-}گ���{ �\�z���hmD�h�-3ݝ��%  � ��_^�k4v{���
j���o|��i� G��Wo^�z}}��w�^�U(���^�K�^{�SĪnμӜ{��h�j�v�o�lo'u�Zy�����[fm�EZcOwu��II =��kZj�W��e좨ogn�v]����Ϊ�[y�C^�^:�
��l-s�U�
{G���EP=;�W��kG�����ޏT4w��n��y*�mioj�F�)���X�-`���I  ���^�B�^��q紥P��ox�OMt��|��:
UWǻ��-�v����o<��֜�Gq��+֥�r{���i��ny�OT=:z����4^���5.�ā�vmf%���R��7|��g��Ͼ�P{m�W��n��  ��ѽs���s���: ms�{ �=� r�� ��jm�,$�M[6��|��@�y�;�|
 l�� �p }�]��9���.��@�s������o`m��� �{� ;�h͚��L_mv��Hz�|����  {��
h>���
�\=� �����M3����z�o��� � ��Ox ��� P��TQAc�����F�}�JR �p=��`���q�w�n�{� ��x�@=�݈ z�{Ǡu� ��� n�m��P)λ� tUժօ��m��jŷO�)I@�x }>� }箼
 #�j�=w� ��v� <gM��\#���|o���`�=I@ � 	(h @  L%)R�` �� ���OC	IQTڞ� ��FF L5<�%R��@ �  ���ST�	�  4 &��$�)�@FM     "I�?T���`M2M1<�ji���_���N�S�?��ִ��/�{Օ���޼?Z�w}�雐���']u�̂�*�AA?����������4���!�#����(����_��|�I'�� *�cЉ�����?E�����I�X?�b���X��5��]c�:��&�u��`�X:����b�X���.�5�k���:�����&�u��bkX�05�kX���&�`kXF�u��bkX��&�u�3X:�� ��5��MbkX�q��M`���5��bkX�bk�Mb�X:��'k��4`����5��`�X����u��]b�X�5��Lu��':��.�5��Mb�X�0u�kX����u��`FkX���&�5��Mb�X����u��`�X:�X:��&�u�����5��MbkX���&�#��5��MbkX���&�5��Mc�M`kX���u�kX���k15��M`kX���&�5�G\X���.�5��M`�X�뉬0#5��M`�X��q��5���u��M`�X:��:��]`�X��5��M`�XF.�u�kX����u��#X���.�5��`��$`���`��5�c5�k� ��X&�X1��]b�X����]`�1�.�u�k ��CX��$`�X�u�k �.�u��]`Ì`�5�kX��&�u���u�kXc�\b�5���	�X1�!�1`�5��X�����/:��.�5��]bkX��05��b�X:���5��M`u���5�kX:��.�5���b�X����u��:�5��]`�X����c`�X����u��`�X����]`�\pu��0u��`�15��Mb�X���.�5��\L`���u��]bk�����&�u��M`kX:��&����'����u��M`�X����u��M`�X:��$f�`�X���&�5��bkX����u�kX����5����u���5��Mb� ��)�CX:��&�u��dc�bkX���&�u�� ��u���`kX:��&�u�� ��1��5���u��bkXc`���X�`�XF�5��Mb�X�����u��X�b�X:��$f�u��]bkX:��&�0u�kX���.�5��a�5��b�X���&�u������X����`��pbk�.�u��#1b�M`�X�uレ`���u�k�X�b�X�5�k �F&�u�k�	�]`�b��`�5��dbkX���.�5��X���M`��]`kX���&�u��bk`kX<`�X��5���b�5��]`�X<f�q��b� ��]b�X�5�05��N11������&�5���bkX����5�kY����5��M`����b�X���&�u��bkXcX:��X�Mb:�5���b�X:���8�X8���X��5��X����5��Mb� �&�u��cX�u�k�.�5��Mc�X:���u��]q��1��^1u��M`�X:���5�����5�kX���&�5��u��bkX���&�5��]`kX�`F&�5��`kX��:����X����5��MakX���&�u��Xk15��MbkX����5��MbkX:���]bk���u��]`�X�u���5��]`��.�5��#X��5�kX:��kXq���5��`��&�8�`�5�k�	�CX��CX��`��5�k�!�X�u��]`�����5��X��b�`��8��.�u�k�#�Ck�/�u�k ��b�X���0�.�x�5�kX�u�kXc�b�1u�kX:Ď���u��]b� ��u���`��.�`�Xk0`�X�b� �.�X1��M`���]`�15��`�5��]b��:��!��X�5�h��.�b�X���kX�u�k ��u� �&�0b��5���b��5����.�u��^3X0u�kX��5�k`�u�q�k�&05�k� ��]b���$`�M`�5��H�5�k� q��u���Q�`�Q�u��u���Q�*�@5��� 5�!�Au�F��X�]b#�Pu���� :�X�`)�X�X��@�:�SX��b��Q5��� :�SX��
�SX
񀩬b#�5��Q� ��SX�k �u�&�MbkX����u��bkF�5��P蓢ta�'D*���15��bkX��&�X���b�X�5��MbkX8냬15��MbkX����\\`��.�5��Mb�X�����:��X��bkX���&�u��X���.�u��]`� ��u��]`��b�5�kX�`���5�q�k �.�u�kX�����]b�X����]b��.���`�b� �	�X8�X:��X���.�`�׎�\`�X�M`��.��X1`:���u��q��`�bkX:���u��냬Mb�X���.�a:��!�`�X��5��`cf���ɑ�?����s��R�?c��h��PJK]اae�Vԡtsm����[����+i*ҲnЉS������(;:��b�+]
���scI�Ȧ��˂�L��z��r��WP:��PsF,���3M0v`��y����oZb�U�&��90U��2 j<�:kJq�s0�i݊��ޫ��&LV�T=q��� �-
117(��y,�j{w�Tt`BIn��c�Hʒ��R=��e�5U\'�qRΕ-�w���VM���t��Y*��Mf�ůXcD/�/�hS�m�F�j����t^����B�=M�d�xAh�)-�n�g�rn����x�\��ve
����d�F�R�Q�Ze��nKy�0�.�����Ҡ��&+,f�L�P1��Ԗ����kHP����f��PaU/6-���\e�s!tR�w��d�OM+�uu�i�g=�a^eE!�{�;Hd�rJ{a�^'7��ȭ�Kr*�F6	oP�U�K��1Vbr��tt��5
Pf�p��FE��+Enؤ�ݼ(����ט�M�{d�8�Ia����%iW%\�j"�n	Nn���1��x,��Svf
��*�ӣy ��E7eYH7�f��x��Y�(V��;����z,�Q�Y�5�b���pY"�G�	� q�#�nځb����5d,��pF��-���w�?������޲�hj�B�$�[��q��{T�ff,X՝z"6ٲ�k[�l�C�H����dby�0Y�V�� �'Q9�n3��ݢ�CAdYJ�<rb��8d��GXJ��֓	�J��F�L��o�m,~3k\Y��,kd����5Y7%�SB�7�ı4�ѺvXN�h�d�ȯ#�`�l��r�n�آ{P\���+�Wa�x�ֽ��!��U{u��o\�j�n�� �w!7���Xز���P�f�sF��m��dP̈́A;;P��n
ŕ��Z]�,;�"�dF�Lո�@�a9��V=wQ����x�^���KU�
�����){71��Q��jj�LICwY��l��[q�]�;�Dԡ�֫f*�
ǩh��r
iX�M��6�͔ǔv`.ڎT�N�V6Ȑh6�lU-F��-{���a�}+$e'l�&0Sv��wa��Q݄8)	54�s-Ix�Ճ3Y.Lӵ)J�E�l�d[��^�TA��k��Жa�M,���7��F��1e�V%JA6lj!"�YI��q[�e�8���h��oK�%I�j�`I�l��,�Pš�=�eB��K��ݼ¥��Q�U�M���6kd���l�H���(X�^^dvk{v#��܋
X$�' '7�oeȢ���ȹ����,^b�ݙ�ˆ�˲�-Ұ�Z��r�2��eі��(��-���Ӂ� n�mc�X�8�kw*]����
��#�V���F��ѱ�/a�(�E=�,I�%N���L8rX�n��ZLm^n�H4q&w&�3KEV�6m�l��*d�	�F�ݍ�v�`ㄩJ��&<��� �o��*�=EK1�jV(l`�Jm�u��R�v6;4f[��D�t�}�1�F-�F��m�.�U�L	�f��De��)��A�ʴK��a�Ze2��v(��c��nQ��RU�ʎ��-?#�,	I�铆۹u�m��XzU5����v���Jn���`tu�v�R����A����)�N���q&�*չ�.�Gkf�U����/V�Lҩ�?^j��%�GB�[IdmEL�N�0⽢+1�QUޕ�xh�ђܕ�.*���`)	v\��)H�j�/���̖���<8ˉ3o'�A&�&��/FKW��,��|��Jb��ǭJe��m�cc2����*�
@��s!w�r�ܙD֙ˆ	�`ʞ���a�ں�%+�:�̖�k	sYkRg��tE�Z sV�)Vk)k��U���oI��Ӧ9Uw#�ՋM��A�cXU=�I�ڳ(��Ƌw���l�(k����-�,;�f�Tk}�c$o�ۤ*'sCv��i�Ŭ%X��e9�e;U19��k�5�ءQ�EU�s%n&�fh��5a���p�Uy�/keĎE���d�2��̎-�S*˨OS�ZMա�r��j�b6�C�+�� U������2{�j�A%%u0h64�D�sq��w��P#��[��E�cA��Ǧ�UI]��X/e1���H��z)Y���r#���C�N�U��*f��U����4ؠMb唅�б\�*&�SCMJt��b��LDn�d�仃����f�'�@^e^2�)m��Cd^:mh�+��p�c�����ݸ.��E���k^��=!�%��b��
��l��[��5�w����#na�TTa��(K7�Un"@�qF�Ԃ������8�Xq-�a�;��
h8m�Ա��A[hfS��*k����-˭,bye
����J�`�Ԟ�M�enX�+TK	N�of��p��n�W��ˬdQÖ���p�=2�0L�)d���Ms�=�9�j�/����S$ې�lĕ`�Y�Va�N���9sI�F�Sn	q��ɕ�ۂ
E�z*̽-CF �f�z�2�AB����f�%�. �#�Nn��L2D�5f�y�0�U�ѻ���4k���N����YI�SGvf��#��!,[��V�Znf]����f�hC�zwoKvʔ@/�z֫�����f�@^62�� �6�^:�)�G|BI�d�� �B`���Z᳢­�.�nch�u�P����՘�x�)����X͈�%�ˡJ�hD¦�ɹ&�")��:
"�ȫUXǱ+cs ة)1��hئ�T���`� ٞ��y{e�ؔ��t�Z�o�ުV^����{��b��ප#gQ�;�� }����q�w�(�2�Y�6�dt�Խq�Y
lSqE{@�
msoZA�ېGb-Dj
6��K�P���X)��Ę�xt�e]F%�@�7^��əHV#�l�%f���Kг�+�FUj��ӭ���d�<���h��K�5��*�b��[R�0��^9/nKV���ySlTQbff��Θ�ڻ��֝D��XJ�PR̭� ��Kr'gM�a�ok/-$�H��73U���6��I7����m�zq�۵6ҽ�j�LGYDZe�x&��H�zF�7lvܵkf�'Yf�jm�#�豖��B�����4*�P�eܷ:Q�ٻ)cC$�D��zn��ZCUU^�1S��Դ�Y�]��w��q�*���Bj:�tJ��8�fTo.\��N����^�u�Xe= f��@�0pÁS��)��I\�MجV���k�6�$r2�um/��.�ERnL[��'f���Wa��C$H�j�W�,����n�T��M�5��9��{U�*�Ne�����^�a'L�*���H��L�aT����P�u?l�8#�UeV�m��Ki�U��l�z!F�u��*�3J%K�wl-:�vK5�ve�WBbڈ�q�t��MV1�n=��R�!yz�J�T�o��fJ��]�N|A6����=3�pFY#u�#%)oo'�ýY����r7Q���84�Q���4�#�Sd�lɴ�S�	�[І����Uac��^av�ju���/��+wjFETQ�F��PӦ�U�ch�yUIkU���6��0����Y8iRu��֜1YOI�7pT���q+��(ȶ���]���y5=��ѕ�-��X.����L ��Ȍk��[�m���^B�X ̼��T�lh�ѻNVP�̴0�2��.'S��]���je��AeKiY�O/0=F���A�!U��a���L�x�T�GU��K��Dr$�R��W;�P�Pa#-Ey ��+&*�	��fa�ӈ��$�ӣ٫r٦�j�H0Uڷ���Ks[�@��<;T����HۊɊJ�4�R\B��8r��)FV m��4�
�%e��f&�4l3N�[��+$��IX�3#pd^��j���46��Q��ZN4)��\��d����6cj��)5@�a��������Rd�l�u4빪�$�uX���Z.9f����a�<Cmmi3E*a�F)�2\�Gq��$5���i�P��Յ���hh�H�$��;�.�*�(Y1��<F��gOv��[EwJ)��f["ǯ�'N�hڛ$q��vvPk7�ƒ����]B�{)����/"~e)��vٖL�j�R�V02Ee���w���f�R�w1����y��݅��=�V�e�b���U��܍�Y,�GM͊��q�w���V�Y���[+�%��Vϰ�Lɋ}c`��f4�=�JX��T��v�X�k�a�Ę�ȍnޖ���[5���M*H�D
��u�7RL���8���-Y6�ˡ��BG.���Nɇ#"�����t�lReG��ݔu=Ȣ܎X
^Ǧ�oooL��KZ��!	8rK�Lma7i��Y�e��%[�^"ӎ��qÂK�s
w-��#���S����VTȩc�-
�!�u�S�n��*^��&
��-�8+�rkLSD��Ivf:�ې�8�̄Ř��j2�D
ݼۦ�p<���\I^EL�3@Z��	��q�d�$���6��i���ޣ�e�U8�՛:�Yn	RVR�be�nZ���̶�2lܽys"�!���������?G-
��X[w"�4�Bύ�`{fc݆�DY�n�$QY!�-V$2�v�d���J}Ї&.;�M�=���GJ�w�4&*]R�%��HDt�Ւr�׆�҄ILƢ���^��T5Ȯ���.2H�Dkf[�L�Ю���ـ��݄�SN��CƮbf�Wb,[(�F+��՛(�ͺت9��FU�Z6���%�E��E�p�Y4#L���X2C������ԋ����e���T�uY��x���̢��mlL,�.��RЫ����m�^6�ܸ��SYj[��0'�D�-��,�;��Ɨ)�%Z�P� �[�j�GU$�V���;�ܫWr�O�k"x���Z�]�
vڻ��ӕ��ֶ�N�j�$�rO��V���lZ����$�Ŷ��*�T�Z)bN��vv<�\��I{n�=kA|���q:V�r�OJZ�[�D�<�(��f���n]�os���5��E�j1=[K����;�"Ie��Z�.I�o��щ�me�K5,�_Ǳ|��p㤒T��D�S�icKV���GWڥ��·�ʹ�r��)�DЫw�DZx�J�J�`�[k"�F$҉E���Ģ�J-ռ�%���DIZ�J�Z1<SR�^(r�T�iF�%ir�n$��1F�3��b�M�۲�H�mKr�D�,jڍNN&$u&�V�isݙ�
K�x�,�mV�I�ƣW]�c;�ڽR#[Bg"�b�W)�uv'��*GSk�j��.�ڈ;f��v�xj=F'����-J�����k��j �Y��]hŉV(ӵm8�'��\�'��o��z�[j��Zj��;U,s�y�-ZM���V�⤝�H�Y��\�T�6�%|��ijT�)�j掫��f'i�Mf�%5U���s[�S�bI��z�*�i-]���S
�N.���ԉj��8ӋT�U�mMX�|u�eӍ0o�.X������SZ�)�m6���-H�+Jr�g+�@��-���N�I����U�Z	�U�J7t���i��KqLU57"@�)�Z�X�b�p[׺���I��F�4h�i&�.��[V
�_f�"Y�h�3��&��p��Z�[�R�r��VҥگDq\Rm��M�ĵ��mƘ:	�$�MW�Rhvvv�]���'�Y8�V�Ȃ�N�\�g_e�I����Qj�]�Mw�۶�V��#��cWX�Wj�v����iŴ���Ih%�C��O��Ԯ#kZ��е@��I4�i=U�Z��s����I%�F�VZV�.��Ig#��Rm0�������jAZ�t��j�.SS��3r�^&�_��|������m*�X��r�Ÿ�U�Z��k"ֵ��b���ŉ<��eQ���ֺ���U�|�[:ե0���A����ie��mjSSk�\�T��*Z��'][��z�q_Pj�]��]��w�V�Ē-�,�T�/��\�'�<gҍ0���Z��cfT�_.K1h���T鸩'K94�,�|�˹D�D�IjU�m>K���#k)o'�)*U�9*;}��i��@n+J�@q+�5.X�r���)�[M+Ř�W�cJ���4�O��\SVb�Wij�D��rm>Tb�[��[�mNm�\���%����iTJ,�T�$�����yJR֡1�Q��g*Š�I���X�ŷ�Db�N'�%MN[�jQ$��J�8�*��kZFb;�[�Z�V���W���u�āmrFB�J��9K��TմykXib���J�i;V�r�Xb�]���OV�@v,���O�ZT�6�āȎ+"�U�JbISF'�qH�Ǐb�T�űH�-�i+�.�V���)˩KYi�x�)j��R��ڭ��Me�r Ď�̎J��v�O���M(��x�%KZ,AO��QsG���\W���Z���]�mGZ�SRԢ��M�jj�W�$�I^.J�2�j�V�k^���-�u.R�rĳ�ibt���ڛj����&݃�_,��]����,WI✺#�bX���؞,J�^�E؞2�ڮP�� �[��g%rirZԤ�<�M�����'��>[��4�,Ir|����B����1f#k5�sC�F�խ:VZķj���h�`�]W�e�i��F*h�ItY��@�I"�I�q�-���"4��h�Q6�$iTJ,�[jE���҉b����kR%��bD��-0m��滾ĭe-�*�K��utZ�mRV�F-�� sRK�&�GJ�(�(���+���\$�`�M���VP�RܱC����	){e���6]��/��%��ț̙r������}��� �/�,>��+~��>z����3?6C��qy����qS��mb{1�R��"�XQ�]3�׷�C�k8�!Ns�9Y��7����Wi��/}��O�fk���㔂��/:L:����\H�+st�lc��d�=~1<\�{��l���<�U����,n�Zq����O4�M��tJKы�S�]�e�,�%3��sm����U�\�M��ilo�,̦�}fɈ�T���+�D
(f̍�9v�w��+�����OؽN\�j�� �Q9���xZp�K��I�.�f3۵��Pm�ݔpD�8� �E,� w]i�0A'	�jJ�=��y�;�nj%5�N8Wb2<r�Vծw�i�)�)�fu�N�:�8�M�ƥ�jP�޲$�2�mp�*�v�@�X�v��M��I��6ͮ�i=<Xy�Pܬfz�-	l�ǽ���#ْ����>od��v�R�c,�=�w��׮�o#�t[}��U��^���S���;ƹ<���i1G��*��ND�c�PF��d�ݳ�ea��⹒�d�*��*�TR�>T��ƞ�Eb�TV�^v^c;#w�vm��"��in�ʔ�_=��qљ���_L~w�Y;�r�E�ΤgDz8`����b{��)�k�v�X�FI6�!E�jI�N���O���W/J9�~�U���H�U��]<��ޭ����R��xѵ����x�ʝ|Vm�v�/�@���ͪ���<�����T��[}R�=�j�fgG��5o"r�6�vf⣙ӟ���a�r�����jf���ʷAs}���@i�昺�vY��i?nm���Wd����>�b�	zAT2��9�l�rȌ�2v#�":�n�{`�ek7�/�]&c�M]�}o��/*nѮ}�Ef�8���ԯp_��5��-s�B��W~�L0��Z��S�\�s���Y$�;#k�n�i��W#P�7ú�1��z3ﭲ�N1���m�um�+VM�ר�ҳ�[o-�x^�h9�#G/���]���S�IK�[�V]1c�Avc���]�c��E�-��CT⤠:�KWkN���n��:�`��}����Y���,�ʶ�g�u*U�q��ѝ`o,�&-�'31���΋D��e�&�_ѫ�;gi�1齊�ƷS;�Ǔ]�;��8+|�7�39�za��]�n݆<�X诰���b�P��κ�d�YJI(���5������蒧=�)ZV�v�7�n�:���C[��,����u.p��X��lJ��Cr��S7qwTjި6x�Ϸl�]3l7w|v�X�M���:?�N;`UŇyz��莝y#eЙʇz��W����QE�_�Vɢ�3WWD�w����&�A�U�ZWS�X7�wB`�[c�+������3�T}N�f���;�ŇYUϵ-A�ܼ�l��.��Q��Faw���R:��j�(b�]YU/r��gU7|�ΰ�k��L֯%k�����J�d�������)C�9.[���WcSV�N�|�\;Y�ޅ1h�7roV�!bڗ��`�r�tsvK�gTTe[�l<b�*�اpt�d���
�72P�J����ɛ|�dc�U�*�k;�zl�麗h��&U����|�a��v�v<����է��Ċ�8��\�a�>���Qxegn�PyiP�@�82�@ރ4��f����&��Z`��u:�Q��v���1��'YCD޵P]|YЫ4n�h�1]�9Gf$��y�a�>y	��:uE6i5I޾�c��W5F��7"�9u �]�I���Ǜ:�a��Ɂaȗ:�\^���pCGI�s�oqꨕm��x�K���3��V��h��W"�IK~�*��c����e�a��[st��WR����3�*\�J	{;�u>;�ݏ4:�N��b��;�ђ].�l�5/t5�ڊ�o+�������Ԛ}��9�BX6�RW��V�b����ζ-ܶ�b�b'3�F��v*�ſ��#~[�\&F)��qw�Y�R��rw�nc�+�Y3V�&]���t�Y$���E;�cā�T[���Α�U��鲕m����.���>|S�I�w2�ZV4�3g4(�{���}����N������a���S�d�yέ;��l��2��R�<��<�6�\sA\��pe�s�d�ok��d���d�Ht���N�kX�]Y�;H3��J�Y��;��6�����#��/I��ڕ[�d̐WA
�z����)�`讴��h����:T�H�W�F*�ɻO��P���9nଔp�ف�xI�$�2�J��[C�.�*L�Wk�fvN[y!�oi{��5�|մ�e��%�P�|��,��س��6���å�B����Y�/E<�:I��y+��G:�A�&���-=η�`ɼ��,�f�TԚ�[���#-��jĎ���rK��u0��{�쨻L��JZ{ѷzD�o&�+A����ZS ]�O�;�q��&GX����:����o)�-�2��������U���Ǜ�jR��m־$�,uU�Akw����"�~��O��ջ���hK��h����:��k�E#��9��w�eH�tS�38�9��S���N�nT�|�������]N�V��#:�}L7$����N:n�����J�`������n���4�r�<�ɫ�w��q�dguw#�m=� r����T���]���^�y�eg`�����lt�!if:��l��o��|$�D4���V��[21*����3�B/v�L��[�ҕR��YB�oR�qoCƵN��ٮ�0��z������m�fڥ�-غ|൉@�5O���w��5Y�Ϭ>���=w}ԁu��d�W3N����rf�c���$�����k"c/{b��Ʋ�`)ڒ��#w,�=-��4m�́�r����N_�tiL��7X���[�ۍ���䊲�!�59�o,�vi6���� OC��&�oLdfn<<w�8B�tܜ���\���rA�'8MZ;��	Lr�:3ko{YK��e�Q��mm�g�lQ���m���ͭs���Q�v[n����;���J�5���<����F�E3]�����lq���j�v�د%��;�n��Բ�޻����:�6K�`5������NoKm�r:o)���y#R�bܬ��I�#DG���s���e�kXZ�W'��;�0d�e�Γ���"-5m@p��z���R�˽���6��dvL�;�e�릱ut�jHE������z����&�Y(�-ч�C�8�����㳹�����Z�cLLS87�L��c�w�Mi�p�斋��)�p��͍`��b��Kf�f��wU6��XN\�O-�h!&vk�U�"����V�i���T�0���%y�xx]��1�"�0MR��Wˀ�*���ӥ4�!�bd����i\���lv�=$9�lU�t������z��q�㌄u�13r�5jv�:�cS����Vjw������������3E��t�3X4��S�@�#�4dL�ٮ�c�oY�8p�t-���9*�I�t&n��l�0'6]�;N�����*���� 4�C9��2�������t�.��`��qk���}�*2"�y+LF�|�Pc�#jr�������10��wl�d��-����rQd�V�t���݃/Cd�|xt�ݫ���in�ŷ�҂�)T:XM���6,q ���Y}}���Fl�A��T9�!���N�Y���MΡfvtº��&vȣ��Jqv���{���tR�j�D�'Q����sZ�GkF�NjsM�b7J���2�C^�o�W�P���I��l�_f��R��V&3�6s�N��7����w=Z$����On�W�Rs��L�16����Z�����iJ��"a��kyd#v���Ӭh;�)��/y����0���T.HPۀE�f���-�c p8W�w�>��GʥC{�k�@��tս��@�ĊX��]n����3r��b��E�Mn�4�� *󎻔N��`py�,T;8����Մ$�Z�l6�n)]"^uk�U�fES&�U�'f����$uk�P����1����X)N�\�}D���r,�K_�1��9ؖt][�hՃ��`�3g�.����N�<�;��u�gRjg,��sk����n�͉}�r�xDj�jQ���.	�پ��w��q�3��Hh8�6�\G]g�S�����%�j���F��,��ʜ�L�sB�m�ޮ���R���hj5��R9��Ƿ69�mj�	iGV�[��N��\��	/�Z�8<�}|��&2�5��N����P��s����;��0��yB>��^	%��K��Z�ʙ�wbxss^�{ï���i�M힗\���ڢz���L��g �e-͠�n��e=G��Z��F������ѭ9'
��#6k��l�[o�����F�Xm�˯q�=������Vx�kU�8�%"�m���&E���m^��k;��g2�$+Kݜ�ɹ���`�Pe�b]ټi�_�����8���.X�7"��amcxxn����4s)LN�W17Q��k&��t)}W�p�A⾦���a��}�\�m�&>u8gY�½9]w�x��2>�b�]�Z�tʂ]΅��I6��jK1�޹Ê7Me��Á��*�S:�02U�t�b�9�]�+Y��\ą��ћnX+����;.�8�$��I֋Wԅ�f��̜sl��e��u�%���Lpf*� R&Ƒ,]M��i�T����a#;L�:��#v*����s�s6qX��J��ڑ���At����;���]�O)n�ˇ���R:��:U�r��,J��A�8����ўЖ�6��m�K �|�:[�!��Tmo$�}��y!#o�t�;�n���-�n����6r�S�,��������Ùy��Ǝw���U�FH;8�<���{ұ�Mo�.�l8���\��^������\�4�X:/�R���,��/	���2��37{��L��$�I&�	$�v���ǜ�ХaZ־\���}[�N��t�t�I$�I$�I$�I$�q�2K��ֆ�}�;��#����j�w�9�"��Z�rg	$�I$�u���l;󈷘��P���-�:���C�f��&��y����<�3��S�$P%O^��H�x��OC���؀o�tuҬ��� #���Ǹ(I�O9�|ǫ�>O;���9$���0:�7�6{	{���μQ��t��yޓ���2=�� ��9;�d,�7�A:�S�qCo����L�s�pK�_ M�;����zޖ��`�=u�q`�!ȏ��W�z�&���p����t2>���Dy��A\�!�0G!m�yM<+J8� ���2����{O�D{ޛ�d���o8Xd��Q;�9.�g7����޺��s����Yz=��>�.ǜ�O=�A� g���Y�Cn��Ez�9 3̓��|�=�
ʊC� Sz����C��@���q ���K7=8��^B}1 �w��Y�e��C�0 �z"

w�?�����?������'�?�?����U��������G��������vtF�a���i��\��:amR&h�g_,9����
��.�6'�e^ELi��p��Z�].u��D�t�s�®ng�>���Ju�J���}~s�	�$Ɗ�w��u�Q�ir�ʕbO�J��ŇGs�qljѧL�V�P�9�t�pY�8�t���⭉��&0^c*������]���J`v0=��� ��	��hͶ[�s���.���-m��%��Φ]��].]�FLK���Q�/gr��(�9�9SNv�Ϯ.����:p��C]]O�z:�6�gF�a��=:���N,� b���Ṳ���^�W_f�`7�w3K�԰��|��Y�ܣ��q1q��O+Ҧ=��y���l���yԭ��d�~o�Q�[�6Pٝܦ�m`�+�j5��gN�P��
.�f�\��{�ז��z�cA��n�Bd��b��ۗז����l�����[��X�ףD
E�us�{��
j�:;o8[[½^Y"�:��x�|LV�S��>U;)�A�޽�k���L[�'��!�q������Y����n[�y]f��-T���{�|�<�=\kZֵ�mk^5�kZ־5�xֵ�k^�ּkZֵ�|k\kZֵ�k]kZ�Zֵ�|kZ�Zֵ�|kXֵ�kZ�ѭkZֵ�hֵ�kZִkZֵ�k]ֵ�k_�ֵ�zkZ�Zֵָ�k_5�kZֵ��kZֵ�|k\kZֵ�k]kZֵ�k]kZֵֺ�zkF5�kZ־�kZֵ�|k\kZֵֺ�zkXֵ�kZֱ�k�8�ƵƵ�kZֵ�Zֵ�kZѭkZֵ�hֵ�kZִkZֵ��z{�==�I�����'1��=c���@�;���g>(t�}Pξ�������]�^��b�Q�����A��Ey�,�k:�%����v�����I5���QW`W���3�v$��Suv����I��;��5%�8�ҹ=���� �ڪ�l�Ij4�"�vL���;{�/��B�˄J.���,�-��Cɻ��CVV�9���m��njk�h��L�H�n�\"���� ��`[���ͅ���W��s�q�+�u��]����&gN-��ه��2�3�&
�G�yZ��?,�}W5Á�0w1�N�i��\�˺���C�u���B�jei�[��V���9m>/��܂�QS�٤*��-�yں�[�W.�M�u>��{j��ro�i�lFes�}4�d�\@\T<��ԝa��V�"�:=�yG:"G�b=�f�n�vZ��̃&��)n��Y�!Ev�^�f+x�׍���41ƺKq 7;1�XI�kd�:���e���P����G�;�L� <�N���G�����Vxn"�
����f�ɲ���{U�3�ާk�SW���I�3z<u�M{|}kF��kZֵ�Zֵ�k_ZƵ�kZֵ�Zֵ�kZ��Zֵ�mk�Xֵ�k�Zֵֺ�u�kZ�ֵ�ֵ�{kZ׍kZֽ��q�kZ־5�q�kZ־5�kZֵ�}hֵ�k__�^5�kƵ�k^�ֵָ�k_5�kZֵ��kZֵ�|k\kZֵ�|k\kZֵ�k]kZ׍kZֽ�kZֵ�kF�kZֵ�kƵ�xֵ�k�F��8�Z֍kZֵ�kZ�ֵ�k�Z�ֵ�k�Z�ֵ�k�ZƵ�kZ�֏Y���}�:r7�ws�X+o6iJ6!.�pP���w���L�|:��2^9������>��Y�G�����f>T�w+�ߪ��k="X]>YW����3i��S:�pw(��λ�޷Y.��Sr���nkt���*�P�s}�]e�qV��Otia�nu�n�b�w��d��T�3�1u�Y��^N�M#z$�\�FN�"��ud��}�AOĢ��B�,��e����8��n$�K�mK�w]���՝�d{j�\&��9:�ljӴ�6wa�n�x�A�X,wVD-!#��f���t�Rr�_-aHY�O	���m���m���*2��g�<��_a�1+�m4w#�i�7�9S�P�xvۈ�w^Q}SZ��"�fqB���3\��øLv����uoN�sŉۡv��R�O��"=��/p�J4x�૛F����[m7O��S�By�q6�"�T���-S�F
��kx��$��
\��j�6����:�Y��Ӝ�5W��f=|��ˏ]3B�أ8��W�������|kXֵ�kZ�ֱ�kZֵ��cZֵ�k�Z�ֵ�k�ZƵ�kZ�֍kZֵ�kƽ��xֽ��xֵ�k�Zֵֺ�k�Zֵֺ�k�Zֵֺ�u�kZ�ֵ�ֵ�{hֵ�kZ�ֱ�kZ�Zֵ�k^5�k׶��5��kZ�ѭkZֵ�hֵ�kZִkZֵ�|k\kZֵ�k]kZ�Zֵ�|hֵ�kZ�ֱ�kZ�_ZƵ�Z�q�kZֵֵ�k�Zֵֵ�k�Zֵ�MkZ�Zֵ�MkZ�Zּ�{���w�����;w�)�N�[������9�"wY�Z��d�R�6��ˁ����QWO�Gn=�y;8��έ�]�5*bXX�{&�F���g�{�N���S���{h�z)�(�f��L��g"�N4���trR�l��Θ�c��n�"��.���>-X\a�ne�nTkV���ȵ�$�ڻڞۨ&^�0���Gs�Cm�.o#�����FfM�iv��;�O2�&S�"�n
�\��T�H'�"�gm7��Mu!ul!f����G	ڝf��v���UUz�����VVfh��j�n�eL΀�J�b��RDRj���n��ɶ�p����^�qV䳸��j)�Wu�b��"��g^�3�z�����7��,iԖ�Zʚ����=��Tk�9
�6���g�۾��f5]�K}R�j�b��R�Fzk�w�����ڶ����{!i?P�1�Ts�|�搙����s��U|�ϖ�+�_R6�ݧq�`��V�>g`�G�D�ʥh>ɵ��Ye�����I��V�s$
���PK�Y��|���X1E���ځW����f��UҐ�>�w���������z��u�kZ�ֵ�ֵ�{kZֵֺ�zkZֵֺ�zkZ׍kZֽ��kZֵ�}hֵ�kZִkZֵ�k�XִkZ־5�5�kZ־5�5�kZ׶��ֵ�zkZ�Zֵ�Zֵ�mֵ�k_�ֵ�k�Z׍kZֽ5�k�kZ�k^5�mk\{kZֵ�cZֵ�k�F��kZ�ƵƵ�k^�ֵֵ�5�kZ�ƍkZֵ�kƵ�k�Ǐ�Zֵ�k�Z׍kZֵ��k�kZֵ�}kֵ�k_�ֵ�k���w��ˇ�q�C�r�ҏ� 5���[5��{��)_-t�"�� Q��w�&�~z�����:�芦���p�owu^M�ݝ���{ć������S�6d̺ǣh�=;���4h�G�K�Vq�aiq�+���D1}�=گ:0_H�S�s��Z�OY����i�Ū�[ŝrST�Ճ]��)�9�

B��u��5-c-!T
\���������n�]��PB�p�78+�dҔ��9�"胼���΁t��������w�vV�e�}3����ѫgs��vb���Ȯ�3P��t��d��v*B��n��z$o�4p�'rK�m��ӏ���vmȤ����w"��<�����Z��Q|��31�g��x��yHS�>�4!,!����w*٩�y}�W��=�4��m@��P3H� �,���I��m'�hx|ꯞ2�hn�wk�UUK�{���7�f
ˡ53�]�L�,�&�I�gs{3_+a��-��{�`1z����Y�N���گVE���E�Z�n̴��tnlW��|����)T/��{�B	��<����C�cq������GM�ɡ�Y��ɰX��sXb��d�G�����+nqيN�{�� �!I�I$��pi�Tw��E���j�x�������yv77�Վ!h`���-[�N����V��nu�q:�A�W��PB�m3A`t�ϛm��3)��C}^��#hЎ������ֲ�����ȴ*%\�������S���9'=#���[j�u´e{��  ���V��E�H�b�T����
����ޙ*�:��:���N�ͻ�{�Ѡ�u�9��fǄ[����*��P8T�ś�շZFqWs!�&%�ɞ0�=��1.�x�",��!vL$ �媙�[hq�sV���z��e*�t�:\!�������P�mx�D'3�e�����ސS0�Q�m��&]��%�n��������xz�#kx:-�@��%��B���)��]��+s��(p7(�/r��Db��
�Ov�x{�np�xpۇf����bǸv�mqG��u��l�1����Y`_sK�̢����X[�� �V�@�;��3����z����׀�=�j���]�[uj��FYo��E"�d���)Aב��qD��k��a۲ �r=��RkO�umG����y�Q�O%s"�~�����"Q�YUl�/[ܖ�
����l���b���<�XWi�%*�����r���D�}/��l���������I�m��&�.�{c��{��g���!!ɖ�-oHC�i�v쥸B�k�����S�L�ݤ/�+��&nX���mNC� k@b�:f���vݨ�^���9�s�9d_^�λ�^͛b��m�\:�ft��V2�Na3Zu#���^C)>;5�ѩVCH��)�n���k�d��Ъ���޻b	B���Js19���T��:%���^k�y$���R**_V�J9��z�o,���Sj	C������7��y�Ќ5����v�6�U\���Jsi��N�|b�m��T��ژ���� Lh��*Ƅ����,�W���]�Oi|U�`O{(yw��kM�;���Jk�f;�*�T{Z��.�ݣƚ���J�:��	��yS8�|�J��2�6x��^�d��3/*�0���y���q�/W�=��1��ޭXn{�p�����'���p�ꊨ�!t�!X�{�V^tr,ᨭ1�4��]�o��Z��Y�:{p]ܡ:�3�Ԣę���]�L�;�F���"��^��0�͛hZ�c7��T��I.��X��r�Ǵ��`�N���V�N�cފg7�8�6�S��/�,����l�ɺ�}�KSo�߀��و�{�˦�L5�,h��V�Kܾ�4vW?!��w�eدxy��]���M*���[2`5.َ<��#c*!�qW� 4ө�������0Hz�b�Aa�(���o!����v��sd�BnUc���Xף�A��3m�6+��WnI��|Õ|�c\5�4�o������\v���/}�>�����fC����DfN����i,+��;/6:Ź�E6�_]
��6×t&�j}�U�2�fʈ�ِ-%�yeԸkKፊ�ױ�fT
7��[6�=�`��(�i��z��. Ȭ��&Qw�.��.��\^�(�<J���"���e�vz�����J���u�a���T)����9S#^��@����8r0�q�*�I^A�Y�fg(���S f���d�6S�4]�v�E@���C���8�RAo�����Q�Ɋ`W��LN�f�㽍a��,��T�T��E<�wj<��toj�j�7S:��UG�Ĵ�#
X���bh�b;lt��[�����]�i��t�X�f���e
u%�6J�2�B������)�h�m�<�Ӄ1m�Ϙ���X�����Y�|�U���Ve��T&��/#˜�8��.�����G�*{Ue�&��Kd�gd׋U��ʏ�"��Bbtx��|Ӊ�|��-�1{���)�\�vv^�T�@]*5԰��Ö�ǘ�hg;;��u��h5��N�=�qƸ����{�̈.�AQ��[��wk�01]�mn���Yqv5����%���V͍vC��r�K���v7��5M�h\&K9�l�T��0e�\e�\�����x�l��V�P�aU���Ӳj�E������b��Y�S͋�'hJ����G��aN�u[(��NL/�e�n@H��{<^
Say9;���k�A�z�Ayw+K,�� &�bټ�������r���29��΢EL\}P�&��{飗��x�!P�5˛��3Gu�-޾�;�ˉK��C��U���#�nnV��f3إ��B��6�J��7�ާ�!6�-&k��K���钸*3�EA�p����M'�`I���;�-]r��=�`�NC�m��e�me�N��5e�s�df#8�ˏA���ښ�B��{w��)�/���(+D�5]�#xùT6��Ju֌��6��p�I��㾽��^�M�SP,>�n۝����NZ�K8=�'d޶�<]"�V)�u2������q<���5���V3t�Zq��o��lJw�����9�h��7�:\X��69H��;��ųU�P�����9��=Hi6L�`�:vDܫ�ڵGM�B���=6�mhv7�m�����s��.���=sPש<�N��㏲ՙ���zK�L���}2$��L8�_f�*e�Y�5ʖ2����x[s�_d�U�V�[�]���PV�0Z�BV�6���)gh�2�}H�]��|(tuӲa�Uk�Nͯd�Ѩ��3Q�V��Z�!v�d��=�"3I�[����Q�1�w;�����N5L�\ ��<�\]W�|S�mm�3�!�~�ﾏ'\�޺���<=��_�?�  *�Y�����������b�`?����p�#����M�2l䓏9��.�+܃��kع�]��=��-�9�h�`F�ȨZ4XB�N�m��՜�g\n�7n�;��/g��\���TqR���Ls���y���x���^7=�����m;\�^8���
��U�7s�nyݻ���<���R��]����m�͹�i{5u;�X�f�a�ץyܥ����˵���p��:��q����7���ݪŽ�(Ů�$0ӵI�@�Q�)��r]׮�ܗ�39:�����[ȗ����ʛ�n��b�y6�|n�/=��;��Wmo��7�����|D�^�t�'[����S�����4�����ˋ]6JKyH�JIR6�@�`��T�F�rf%$&JM�#���$��9DE�^TDon)��;��׈^����;���M;%��`�����\\޽��5{�����^���;�0�I�SI��q�)@R�;`UP(�Pϛ,�F�O�d&
'��G�W�\�ix�8�9)��I*�іS@�Z��2��~��^�j�ոk��,���qk\����r�œx�����eԮL���J�;��ˎ��V�&��2�I�0�-:��[7)W�ž1h��{#p�d+���.v��Ә7���y	yg
��E�v�k�i�3�j�}:�(����B�-�!]�+�
aQ����ѫ��j��"����-4��X'!$�
��8���]v2��l^ʰ����39�4�Ҁ�DYϻ���z�ʇ��ɏW/QA)����S���oT\��nP|F1(t�X��es�po�e��r�����j3��x�G4�S���,�G�8⅞�hjj /��g�Ub��`�m�5�(X��ٰ��*jx�+���l0��t1�mc���RHWr��<���ws�MbCz ��6�FT���8��3�r�f��)�H�]y���l<��nK����H�%����˶��e_:;\m$$��۴�u,=	���(�85�I��p�X�>�-�ո��4�wr��ww]v������$�&I$ ��`��($.�f�e�WSf�vp6�˹�6�^Y�W�.랼T���s+��|�SvK�sX�ݜ�wv�K�v�ܯm�ocU�����u�\r��%^���h�[��y�s�1�u^�������a{�vw.�����.s�wU����������6^���o���xc֙�1�g�4��n��6��6�q�tP펝�Kz��x绥��wČW�*O&�0&�%H[R��[@�	�,/�	5Ң�T"��"��������;W��S��U�r[��7n�g���6Պ%����y���y�Ժ�c��V����7r+���ƩK]�qT�G�L4DJ�D6�j��&6JD�"$"��d�8!a�ԉ΢^:�m�6�Y��g��NmN9������eb�Do!��6)��Ls�n��j��3�m_-���)��[���۶UMJ��K*�	��!��j�*wZu��o�̞/�V��/P�Ǟ�m{�w�b�i�F���Ѡ�ā,����P&\�4bJ!�=��e��[y����i���E	���Hh��x���Cn2�㦺�lt�8�[֧+�=�(�kh���mN:����
r[�iLu���7&_�����p���d��Mꆌ&��2ڎ4J��
��yz��֎��c����д,���Yh��\!�P8�h�[�����om����{��:�����f��wnW�κs�ۅ�7d�G7��x����L���j��0mμ��v�vp4>n|��^�:���*�[����|d�-�ңM�d����H6�u�^{Z:���9Gv�/V�ڋ�^��og�l��X��O5���ڽm��2��sqγ����ۄo3��z���a��ؠLmlr٢�a'��08�
9H6Z("%��$��d�]�Z��Z�9Rۮ��!�.b�C$%!��c�P2"��nL~o^��1���ej8��EGU�o�|�������+��YR�[�9z�>ڂ�4��e[H&qǏ���}kZ5�kZֵ��kZֺ뮺׳�HI�d5��5���Z�A9����㊫mk<�W!QE�8��}k_Z5�kZֵ��kZֺ뮺׿#�w��f��d��́���u�X�iYfj����ˬ�L�8�$$!0��<x���ֵ��Zֵ�kZѭkZ뮺�_g�z�/��kE��z�/�ϝ���.��B�i�]e�E�������g]f�k�O���~}hֵ�kZִkZֺ뮺���ߎ��Io���%��+I/�۾�!ox�Q8DBM��v�"��ݻ[���d��-n��wY Y�Z��]�4͒28�*ޥN@�%K�� ����<y��-W���U��u�T�����Z�]J�;�
��ԀTc���)$ʻj*j5a��Sĩ$�(V�	�Ҫ�3Z��b��VB*��[)�٬�\.��5� U�N{�JY �R�m� [ku�%m�f�2@�B�� �Q����v V�J�<�GD��d��m�lH[���t���X�}2���/�}�yE���Q�C�����W����uKK�eS�^k�:��W\]6tԬ-`���ͺJ&օ둋�Ë(UF��ц�P��駮<��n�4d����F��4��f�?>�y�ɬU�P��QɌQEp��^o��������jo�~y���Ow��]�qA#
En6璀��������x�8U��^q���ݹ׹�{D�--;���v��ۮ�v��
=�ݷJn㆛�t��nTp�$	0��^�+M�����t�9VJju�0̬����c�-��a)}��*5�Jf_Wgs��U�׫��\�ol�u��Kr:���W���jgi���=mt�qc^;��wlv�]ŷcr8�Kn�3~m�$H��q�đB�ԔSPF�b�s�n���n6F�^�z�<������m�od�]h�:�ki�q��������Sl�^.;�ׯ5^:����s�j�+�MK�:����on1g\�)�1�طL�uv���wl�s�z�	�$bF1�==�Ӆ�z'��]��{�z&'��Uۏn*9�G L��r�֦�
P��D�����{�n�f�ܸ��I�1v�͢�K�/��
��Y⊕o"["h�\x��|���v�����i`��;�>�w!����EǯƜ&��M<ࠦ��[�csz��$� �٩z����gsߴaw�K|��SD�T�8V`9���\	��͑41�*�F�戕�J�r5˓ss� ���¶���ן_m�{~2.x�����=����w��*b�u��+��a��%K���_�+�h�������"c��ܮ_E�7�����;�qf��'v�u���u��ǣ�죃=L"a^fj:ZR#Uj�M�yQ�Ĥ#��L5�e�Y��AyKh�a�L
�O��^���%���hӃ3xm�Ѯ�r�[e%r�U��y��4iX\ϧd��++� ���ǩ��i(�ϳ���]b܉���tt~�G���6V��ͬ�@�`icEM6݈��'d�=� q jb��Y{���uNf]��u.�9�\B����+I]��$�����۱f��i����)Ī����uS������ª�z��'r�;�E�U��p�E��t*��m.��S�q��(�ؒ��i�ݞ`�0d7����ϫ�jI���X��� �H�jO�n����$5bWz�~ｸW����o�sR����0g�"hdlf�n�J$�<>w:�.z���8dϽ����W�i���v$��6��o<�>��khC��;�R�4��nѼ��b�h6S�{�Fp��|�����Og��� ���o�Ea�NqK-j���QL���	�'�M�5�q�XGC_'�L��܏"�͛�J�8k	��>4��f�+�g��a9�U	N+'�m;c�]d�F�ʜ)b.�-��T�*RJ������_�ԺV�t^��˛+&�Qӧ�{1�(�s�t���H������[n�zL�T޽d�c0v���Z�1t��:�:�F��2HHP�p�~?I���x'���K[� Q�ה���е2o�	��2�O>�Wݙ�C�}֯DiBW-q��=!͊g,�^�����nw��RY�$�G��q��x{�Ej22Ya �}��|BlEC֯3���ҵ�Pc�`�T=~�^xܤ�e"���*h��>-��ٖ|���:�٨���UV�|3��,�m���ER�p��[�ﹲ|A��L��v�#�=�
�q�xfp�����5��l��?���������,�B�d�0pር(F�x��gM�Z�\)󫝯o�/�nb��$yS��Ԭ(���Bl�t�����U���N|�Vw�q1U�/�Y<�yN�>�����wj�6ȇqR�7�Zcm�]�k�/%�E����Ubk�����IY�w�����0q�s�UK�ow��̩淹�F��@��֓�8zm|z�}��eA�}�R6�k�
^}s���8HV�����\��t��c�J�]w`��(MX�D�#	�^�9��0V̴;��K���>������E�.�,�%�f�$R���䯲�1�މ.��NͰ4'����u1~�U
Uߪ1#Ō =�s��:������e���u���������`�UE�`o ��vǝ:UZm� זh����dףT�1'�P�(}NU��'���#�J}���f���g����:��Q=4◷3d�EO�%M��.�q<S��dn�fƪ*�V5������1x I�^[���m��0�:�kg�X]�Zr����M�]ٲP�l��1{}��V ��X�5������9;�'���E:��Q^ϙ7n���+�]%�)CL����1L�ٴ�Ty���]T�{#���G��Ј^x(1���v��V!�z9��|��>y�w>WP�߅�����_F�sM�������M�F��ÕX�J�g��㧅H�8z�<�9� L�Y�B�E]�,�I`��A]8ʒ���l�I��`���2[4L;N�4��_Z����J�;�X�N9*h���ʹ,o5�{�+�4�ގ������Q�=:DB�]��T��6u��A�8j�{X��|����)���KS(��<yb����sM��;������r�r$Xޫ�sl�1v� �9�����o�#=pt��(�5��9�č�W��u�wV8�����n��F�m�g���s���<p;��|;���7���D�ޯ\�&>�ӬI��{�לgl����%Z��r���!_=	ϺzߊTN�@�m����O�C杖u�Ʈ���<����G��0�>�?3Y��+��o�첳M��PE^ǌ��ec;��y���0b�&g���0��ź��k"j�L����=��y��s�j��l���>�d�6)W[����,��� 6�k�3R]T��_g������ޔ#y�� #ZU1WOh�uN���5
)��"M=hz�gV�^�����(�*�j5��O��s4Ԅ��B�s��V���d��>�@�{a�ՙS�^��G��c���QΞ������F��U:��W�A�YA��#�,�x؋F�b�Z��'JY�u@j�_st6I�O�-�vF���g����m�R�d� �J��Aj^�Mƶ4�.кbͽ��/�OA��#Km��١�࿭
��f�Lܼ�x<�|,�dxa�S�8���;��z��.�솅aW��_Os��Lj��X�3k
��ö�oS��E� ������vħժ=G�ed�u}B��m ��^����N\�ѽ�C 5����WL�õ>�_� �$�X^ʦ.�ė����������,35y�����*�/�ٟe�}:g��7�|�]/j���01Eb�������|�fg����.��s��e��/u]m;�RI��n}�}�o�-�V�5��9�����л9o��r����e��wZ�����a�%^&=L{f<� �g����3��+G�^���fѬ���Ԑ5-4L��4>طʆ�#��^hc*FL�m-�E���|�`�Nzu9�ϻ���nu��x�o{3
�/qI$"2"�p�V�D�"@�?rt}T��ړ��*QJ���o���8k@>W�ǘ��P`$j���Yz��+Fa�z|:���]բ����|/j�֧���$+�a1z���{a}�o�tw�]9H���<�$x�4��O����>L�"�66C��k-m�wh���=�]��<�K�ݏ!��Xw�:��IJ�����+�}�v%V�
��T<<<@>  9Iw��x�T��U���p>Ũr����W`^/}_[�=�>����hh��c9#��4،�ԏ�*;��� 'ٕ�{�����N^���E�a��x[��ѾY2���7��#Jc�7��[$��.]:�}Sy���ɪ���[���&�Ҷ�ir;36z��'+W��qM*2�RI�Il�׈���]�C��U�[�@�W��8�wVE�p�G�abo�]����{r}L�B��I��_# 3c�rIF��B�V"�v� u����,����f��y��m���cF�����8����}��}$=y���K5�{��L]��&D_���Uq��k1��p�׏�Щ]&9�5�,�����M �l	�i�Nf��û��I�����F�����Ǒ�&��4�7��(�n}�C��1a�1 �����p�����/����28��@C�9d�	U��⺝��> ���}#��Ρ,N6щt9չN�����|@>>>>>!ْG��Ē�!C<�im>O�P^��FNA�k�^��Шur��Kmj�%L����R��-ܶ��� Z�OVo-蚴������Q�pTȩ�H��f�u����\"	����o�>�_ojU�;zq��Z�%����#,(��p$n ������V���+�o�K*���ϣy��V;M�}㦾_c-\<������'V�($�Vy��D��a�'{:�M紌!�a��R_���<�g%��^aT����C�	�>�T���D�)U˄nKk����.,��Y�qX�T)�}x�/��KoV��������>s���<w���o�D;F���3�$���L�8w;�vw/Ic�����?wzh	޶���D�����}����[��LuX�j�^Uv�șQ��m�l��邅�4���:�(޳�ّ��m`ȉ ��C5 �� �KA |l�3�2�a�7lǻ'KʝmȪ/��tF��5e�vup�8�����-Xc�x�V��xxxxx��|G�>Tzpv%�Wdnl����!��8���R�>��'gǱgM�K���M�F��s_W0ؗ�2Ĥ��7dڌ>2����X��O������t������<�|( {8�3����ǡu����oO-�*�v���w��o�{�	�o>����B�w2�g�&��fMex;{�	mm�w����|j�*�J�3!J�)��7���<m�͸�6�[�
�N����6�N��Ԍ�:[Q.S�l㨱{J�1|��n�CQ��Rl&$�^�8����5ָ�"nc��B���>�z�7�oI���a�@�>oPx9ꋖ(^�nz%յ,�BI�Nʵj:�v�Q�Tn<ikz#D�Ʊ�|�q"s򯾽���w�ƨcry>��VGx��nҎ�L���?� j-�UZ���pq$�]�7�M C8�����^�nd��ێ�>��{:�9y������N��O��C��1�(I�k:�z����7qsz�g��,}��G~�����ǁ�Wk�C�E�ԯ]�f�}�:p��T�:�ߘe;�h��2fZy_:ѕ�*�Cs�r&��a�����_ǂ6h�����`9WU����|@*�G������-W� p�����G*�E�T&�le�e��PN0ͩ��[|Y����;3��}���,Pk������]P�cm���#'�P$�y|R��2�$�0Q�N�c�zc<�3����E���Fl�9�`4����9�r~�N����4 ���h��h���KpC��kk���d�Y�#��� ϧ1�m*w�&c+'dKn��7"�Eϕ���m���,Tei�������
��J��Xyk7�����iG��l��������s6������P'@oM�סb������������5��q<��5�r��O�����DE�d��݅u����_}��=�x�]L?����i�
  ��I����l��|i��4�C��#�l�{�Pu�Rs-r�I��H���]u�&Ki�JGW0��1�[.���ނ�Kl>y���g]^NKN2���)���.ѫ����iy�c]�=:U���Kޮ�y.�:��mr~R��wEo
���^�䡺�z̶��*�Q�&��+Fp���jf���^0��%0x;ޒ�er�7��')��vE0gu�-����h��əW���CO-��:`�n�N�Njjˢ��.ˮ����q5.���������)�˳��]��QZ�*X��nb'z^���N�J����I��%����a�v�m1H$U�Դ3�TST�YVs��闖�I�7����Û���X�95ޥ����JV>@��#SO�	�';��up��A��oE�Q=�/_I�p���h(*jw�q5�TヴՑh�����7q���G�q��Թ+r���<}�WMU\�guܜ����C�e�=�"F�5i�=�woY0��y�~\��z�m��;�BC�荤UW!z���<(���v�>�ä������]���׫�C��#67-�%�H9�J��-�GG+��O:)Ďe,�%�pX�{~}��u�14#豖Dh+/�����T�l7Κ��E�������x:蚄]R&K��сi}�q=n�c��'[i[���C��.<�6�RPXt$1���1��zE�+422A��U0��,�c:�~�=�7��[��]�k7tb��x�n�t��O���%A�����{�AU觝�F�oi�m���f.'v6S�ּ�/r����rd�X��᧵��d@�g�ଆ�I苝����YL����w�\�-X6�wC�	p���7K)U�y�C<�BfHq饈ssP��m�tN]P��Ίd8�\T{5)12C��[�EK ��\y�,޳̤�8ͼc+$���[w���u��p"73�qܳ[�C=)�⬅s^.�c2{V�p��9�p��J�zז��γ�WwI@��M�:�,��j�y�418ql)2�Q�����M]��L��	x�<v^Vdq�Y��j�c�s�[�b�HG���dݭI*����ҵZ�F���]L��6�6+×G;dAT̶��H9Z��0���X�0���u��t��zo;9����-#WՐ���w39�EE0-Ǒ�%|p��Y���e�ܺjw�O�E����}H��s����y�M%�R�z�uekNtW�������������҃B0������	����q�j�p�R,�b�J\�ED�~k֏k��GV�ҫB��*Y�?F3O&���???5���kZֵ��ֶi��}��=��|��O*jQ�%�2�TU~[�2�m������-[T�u�fEE����L�3<��N1ǧZ��ֿ5������kZ�֍kZ��Ǎ~{�EVUTT}����m�|�sʈ����-b�v�lEFf333!ێ8���k_�_�������ֵ��Zּx��_�<a�d�L�mX�j��Јҏ�M簻ݳ�د�4,QYZ����q�=��>???>�?1���������ֵ�Ǐ��܄<�3g��5��8�M�b��D�"#��3��
"�*DAժ����QQ�-�_}O�:"�d�E�UTsK@�Y`��[�WN���hTQm�Eb���ł�;��b�Ɍ(���%��*�
F*�._��
�EV����D�UJ���7�Nj-i�c**�}�&iiQV(�[b�ب�R�/���t����ciUPc
��ytQtUc��jJ+P���qY�ҏ7�k��9P�aŗ9^���ڹɭ=�1�?K��]fp̎=�g]���ޓ>^88ノ0��0?�=^����2;��q���DTDCL:ȷ������W�m��`
� t�)f�oF<�����S��)�꛻�������o�|~1�K�cʝ����7��T�.�{%���<��ȇ��5�t� ��A��0M7p��g'�}a�y�#���O���~���R��3��6�ɎOy�ԏm�����Y R~Ol������t��Sp=T����E��s�栂ZaX�fr�{{�����n��m?�o�痆���=Ji�=k���:�p!�(;�^}�B������ċ"iDdDTVFG�{������|!��<~����I8�����7g��
����{g`#����8�ӊ�Kh̪�J��	C��3�	�����ǵ�ƫt_�G�o�7_0�}^�㱰�^
=�c�v%=d�'� A�-�(�l4�`-���N<eGk�r�r�Ȩ�Wu��,�/Sb��75��Q=���6.�YL�7/ssu56�5s��ly�C���9����s�p����u�<�g���>Y��]^nj-�
5�w�}�s
���V�3�f���m�o6����k&����1�ڵ>/�彣������R�ˬ���)�O�(ļ�i���j���^����{U�킷#^���NVz���'P����B�X��
��c5tz:�k�$�1`�}&�R�s&r�;��o.�M�B�>��Y�OZ��e�W����fq�1�81�'�}��o���#���w����?;��� c�l�#��9$g�{9������ټh����&v�������� �� ���ceyD��=��ςp�]���\�O���ƷI�}w7j�^��#���� 1߇���F~����v���]h{Z�g���_��5�R6����Q�Ox{ɰ?<�%�����}|�O�a�Sia#%$ְ�&[��Z�C�q�;N5.ܾ�B 3/���)����M�	�ܳ���'��1�h�a�MIG�"�%���M� ��ZX
��w�|���ǥ5��^>�  ����N����x�B.��ƋQ�ld>��6O =��7󆂢[߆�4x�_+����^�9��Ȱ�~��a ��f01�r_��Ym�Wڻ��M��1���5����Vt��Q�ם2<��+�G����똊za�-�D߀M�1S\uj��cxQ-���c��:{�۲�{�Aq�Muo�&�3�/�����)���Y����mN����!f|�8���b�X�H�Ǿ'�����^,�3��n��E����b��\S����,F�2�7��M^�Q���l��CP}�e��)	��}h0�1�Q�2,��m
��t��B=�aaX'[�kXN�v���Ź\9�OPi�3�qq������?W���8ノ88�}��>ݟ{�a��͕�**�%��.k:vmE���U)zэ]a���w�v%������/:��6[����"4���~�'W��ڱ�ޯ����;Ӎ�F�Cuz9i�^P����6'o�C�̌;���X����p���^������ߗ� ���)3��@O����!��p#t.�(�<�e�uo{� �<|���{�g�^wrN��C���zq�"��P��F��~�{���O���/���z���'{��yb��Vk�9�oH)@�zfܝ=<����'� }/=����Nĕ����x�!���T*�\�xE:����+_���椡2�z��'���7!����c�^���c�u�Y;]�`[Ã�s�zW��d+
���/=��T~� ��9�%�/P'=Dk��`=��~����w�r_�;?s�zw�g�ގ��� �{"axg���uQ臬w�W�W���vwJJ�x��K{����n���7^����0潸��q����_���&�80s����D��6}B��,?}�<Qn{�@p~��;ŭ��/��D�|����/\?�O����K3w��9l�v��s���ިB�`�(�=Q,�F�+�� >��,"���g_��R���3�pvԪ�K�/��-�{�	;�/H��k���a��^�'9q��"a���Ѵx�s���h��_s�钯1��;�����ڱ��[��fm:�t�smQ�ځ�4{�y�s�m��9I���>88ノ3���*�6�{Y�pO���5��b�AƇFK��@²�;�W����Az-�����ǻ���]�n��{�	>j�����z���@�V�˃��K[���C�ǖv�u�ƺ!8�z�[�� Y���)���/}�zCV�Gu2`��)Ǩc��:��
�2�;y��l�;�Pe���-�w� <-��r�f7<����)xQ���'�==^��C
��Mlx�+���mU���]��{��A�w�
�W^p�k����i�����~���0��?0N|�ɯ�{5<��J�S�И���z��&�罪y�}�tߎ��^�0SU��B�l//������o@ё�g���)t�^_j������xg��t8�"�<��`�Su�\�^���}� (��=�0�Lrf�k�x��{Ũ0;`\�&�t����,E�1@0�^T
s�ly3�gצ�q�!YW���ۓ��l  ;ߘw�����9���\M���z�֤��dR���KZp+��g�2��Xt��X~�q�c���fS��0����{�)���1����8\
��~��ށwr��,����r»*Z�Tj��N����Z�e�cj5l��q1Q��~��G�c�yLeM�z�Ϗb���Ŧ���)���������9��NC5h����9�[����|�r�O�=�q���b�ߞ�[�������b4��Ա/�/X󼁄!��|x�d|w�@������b�[�!���nb^�0r�Z�������ip)�g�a	���~�C�E�K��Oa�|�}ފmq��n'��6���ʽ�y��>���[�y���< �@���	Z�C�#������
`<IkN�3m��U��=����Yz�{��{�¼�l�Y>��n>`9XJ��O��d&�q�a]�
�kx#.�L��'ꚫ¬w�=W��bf&SFU��M�j�����~�}�>����w@	c��1�p�u}�W�{�����%𶱴�:u����JV���P��2�����8A�Y�jpae��+����t{;���>?[��%�l.,�������5�YlrR'CD7dsў����{5zӖ�p8b�W�Ew�k�4u"��=aǞ��y��鞋`��|#̟7z�!�fմq���<�\<D3�`z��xG�_~]�;#}�{�.~�^�@_��a� f������U˷W�� ��A���&����Ϲ�*� ��n�U����U���Nv/��;��n�qP�;�#\E���۷��e���K��)��Z�V<�(���;5��r���=��6:���E�]m8���7w�ں��;�L�qͰXPak�M	����T���_�������^^A��dBA�����߿|��������q��"&)�yٱ��K�����lk��(��C��|aΎMN�o.��op��фσ���|8R*<�@��a4 a��ޏvwR�8>ld��#:r��Yy�w�tU;���.�$����ɎxGq��d���q��zSX�=���O���d��.$��<,��3���~���<���L��6~㔉a��7��s{vъ�v2(����w����0��?��+�|�x���X�����aލgnb��S�.��B�W{�W�o.�l���נ\m�juf�z@�^��0�AȲy�^�?]�-���s��g���~�z����.�M�������zn|�?P�3}�vo#�����W����k.�ǧ�P6v27q�KZk���R�kx7"��D?70R�^&�����5{&�c���1� �d۹hBz�Ou$�������vOl������<>����[ӯ�1 �f�\�kMJ�z9rx� ��p��#^����:xbO༽���?��x"���^1�Q��g}�W�(���*_�h��,6zoa��f&!9��]'��(�s!f���o��+*t�p�3AtkS�n��V(u�=� �>�K�x^��;�6��T{�����܋�J��*R���_:�|�u%�.s�hm��=���}�M4���Lbi����{ďH$O�O¿���O��#5X�|�mmL��8�9Ta��;��}gQc�;>QA�N���V�#�3�Q�C�����7"�DK;C�Vc��%F��i�D�t�MWt�|��A��!��M��n�Av,�W2���%�œ��60�0�K�{�u�@��5���������J�w ���N��ճՄ~htq��XϽ\������h^v�O��Wz`ـ�x:𚔣��`=�vOf�2�xWW0i~q"�	�b����A<�z��k�xM�������J�oH�sl�0��z�EV������y)90�j�5꺵��Z+���
O�I�����h��)�+K� X���#U�\�ѱg�f��"�.8���
��K>p ,�?'��1��.>�i�����e�s<j��_�J6K���X�}>��4�Ek�E*�Q{����Y������5�ccB�/~ߵ5���3Emv"x&����7��_y��������k��Wa$���Z��ap�����ʻ���SL)��Z������_R6U�L;�꽚]/������-�_�˞��Ig�#����7�����y�-�ovgW�?XC�yt�'��mּ����xO��RU�%=��8��{�OǦ�e�����;N)k-m��	7���Hv닓�f(e�|B��YA١�+(p\#�����=�M	3Z�7�ud��mc�k��+:ݞ5/�1*d�2\A��|�{_� ���|�14�V%�j�1,�.DIE�O>���^�~�I��C�O?�y�����_�F�O�<&�� aq���wϭ�j�<���Ci��%�uW*�|�S�֬���B���|�g�g���.K�/�W��=Sª��r������(��҈!�m�]�ۡ��/;��k���`~���K-m	=��	 X����ޗ��[��pZ儳�{�t��O������DޚqL"�yw�r��~��Q�b�P�jWFAT���%i{���0������@%������K�g�6��I��+����	�q����f��R]� ��M^n�����yk��S<��|Xߟ���9�ゖ3W��G��;1pe�斥;��y���fĀ�<3�4�aOU)<4���P)�����h�CF�#�_���<����\��V�[	.����3�#��o`�5�Cw����W�F�x)���;-V%�;����*p)mς�lf?S+�K@C��B� ���cC��1�_���1�r�Z�6MZO.�
)�L���g[VE��S:�E>7��X?=��Ld*1'u�P"��i�q�3lWݸ�띰�BoBwԓ���|�X���r������ #ĀG��]u�^3���I����&�����F<�+�_,�VH��Sv�9aR�O=�)z����w�Þ�����L�:�ĳLCM1P�H�Ⱦď���w����z��I)0�&%���#�O���m.E��m��<�Ql�� ����$;�[1n�7&��l.���+�x�^og��L>5���+\������C�]AWG7���;�j�7}H���V�Կ����"O�H7C�$!��>��i.'���~^P1?uz
{צ��xj��x�����V�3ĝ�$�Ɂ��|�lǏ�;���y�����~zz�y��oxOH��[ɨ[�[���DSCΙ�^v��\�v�xdi1��"_��i@6�OY ֐�Y�Ծ R\s�'|��ia�m�t��07/�:PU��ٮ����H�wޠ[��
��������Bv�,�vl�����A��� �rmg���{1i����z�Y��C��s�=��	�@P#f�Vן�|���|��G���쨬;٩b�<�����C2{�����B�x��מKm�������>�8��EC�ځnv�[�'T��=;�؍�ؗpIVP9g��t�͇ �����d�(���<�n���u�_,{>ƨ䑛��K������Ű Cp^��ӂ.>��R�ٌ{M��o��y��`�_�1s�����;WQ���MbvHa*��U�R'6�K����g��\C�q�k��b/+K��ao�U�+�2�5՚��p�ۉ*{}�3�v��_N��ьs���$�w7�.�����O�?����pq��3�<r
p��= �
ܝ�V�xva�'�>����H�	�9�
���ב����!)iܭ.�ae�a�<�m����;�t��j�a_��+������&、����|��~�4bl,:�߾���=-���4Q��5�Ə���6��Cռ�wnO�DX��@,D��\g��v|�7fbɥySg�5p,-?P9�7��N�k�a���I�Re+��H�X�ɩ����y��0�\i���4L��a��D��(~a��������
�<�5���=�ݞ����d,�\ϡ��wF�+�����{�=�)�wK8O��]�������.[�1�\E}������s��NaS3A�,����ܞf0�p;�3s�s0���s��n`q�/t���:kj[#��iWI�����%���M��1��=����؛�2CC��g�NlOܐ���G��C�����c[\���z�}��o{R<�
���V�3����?/��H	��!���~�$}��Tk�g�F|���/Vwp-��L{�ղZ����Mdc{�_�~��{��:�Y�ü�ϳ�D8(���,�}w�/��u����j!r�S�%���-*8���؆	��2n6�\oi��� �T���ˠۉh%ƞ�pS�v1�]�a��w��6:T����Gw+:1s&����:�8�Zi��|��++I�|v�i�3p�b��L�^��t�!�����N�
��Ԡ�u���M�bҰgTh<�lֽ`رi�f�ы�ԏp��W`���]R��o*,���N��_ST�	]����Jg���M�MJ;����xeܶ�M�cq��
K���=�B�!eGV��'��봰���u�КF��27�JTvњ#���˘.�d�v�5Fu�v.�����2u�$9')C��5n�z��C1,�n�wَ�43[ץ{��3�e]�]:� � �͵�/��s�&�
���b� z��"r�bN��s�]�/1���޸8��c3h6�.�OZ�ip�ܺ�����*Z�xQ�v!���2���[q�;��[�:DZo��
7]|��=���1�iⴻ�uxj6^6���wu�o�f��q�TeܼF16CJ�S5��:Q�xcPI��
6z��i�{O�>X�t�M�L4�E!��+!��j�tJ@�d6T�(�Vj��Yt���Je�a-��:w�oYI��t�Y�dG�<��	L)��h��)P�m�]�w�|^A���+b��0�v�W�X~���>������9b���40��v�&P����Ŵ�j*�g7�f�$5��ẻUn^�2��5m.�(]�B��6�����*%�h��Aܲ򵙋&T�`]�to���.��No.��-O��x�fB^��ֺ�T�v�m��ر�d]PbYC����r�j�z�NZ�ٜ��Vp:�K�P�I�>������r3���A�i��}9�֕�+ͬ���j���t�-:l�2�宻̜�z�^��������#z��$�	$��ھ�6s������'3�/
�!�����n�q�d��{FK	�s�+��7z���jF�Z9��M���Y;Z��S�T�X�.JP�1�tގ�ٗ��V���Y����$V��J��^j��i�n
i<�Ϩ짘1���®Ț�k�qx{ک�{K���z�i�wt��`�5��n�j�Ii��d�J3����\CrOU}�.`����i�Τ��x�|��� �T�i�b�G�R]�S�:�CNw4ԝ�؊���\���s0Z�iݢ���AQ���>D�Q�E�kA[G��Z��D��QmD�@��֥QO�qǍ~|}~k�Z������������ֵ�<x����B�����&3$C��aR+�~l�6��e&c�c�<u�}~k�Z����������??5�<x���3#����-���R�Z�"�R���X�)鮥'��4��������k�kZ������????<t�O���{�U�������R�jQkEb***#�*�0\��p�KK����Y�4f��5������k�kZֿ?>�����<x����'y���#	$dc��%`�"��U��Z�(�2��X��ֹ���[h��ڔ@���h����E�R��&bz�A�Q�b=h1u�����֨[_T�#V�^��
*���8��UE�J�^���U#��/���-��ƥU�Kh�F/�(�9��^�QV%������U�({�<�_ITGUF�(���O�ڢ�Ty����b�:�sDkT�X[B����DԽK��T(�Q��("�jUK�~���sE��o�a�����������,:�|/�m~9o��n��^����V������S���4��Zޚ^znꕶ���m��k�N��T����u��-3�hf�k�/n������_0�-4�PⷠΩ����v)��沯��,��}�k;�WHO�4����i��ٗY�m^Ώw�:��&�u�'Wu��J��]׎z�]�M{��s�k��js��ᷞ�igqv�֛n�q�8��-D�νڦ8��|���˼-����6�C�U�+׸�n�]��Sm�u�j�=�����S�x稜�o9�(���x�sn�]׺�\W�������܍�]��[�ru�/^8�y���ǭ��k�9r�9Bѽۭ��i��׋Ȋ�6$8�׀�cǊ�<cǊ� N1�(rAB	"�"H��	���;���H�G���ܲLF��
�ܻ�`�4"�z�De<;+BD�s��Wfe��5�aG}e��u������[ ���G�;�%�%��W�؄�
IN#H|�o��6��6���e�d����LoU�x`x���������M��p
�?K|�6������d�Q��`�J�&�?�Y���;"X���d�6B鹼��߽��	^��x��~b�}��?|��	�ur��z�pV�SV����^��H`j��4c�k��ڣg�ߗ��?+�{�/����ʣ=_�����������nO��_��QM�=��_p�M-��}~xB;�>���b~-$�����ܟW&��iڠaWf�<�\0�юu�'0ޘA��ǂ��e����5��.����n�J�s�4q�z��!o ��w�Ȣ;��gg��@���\O�6���Ԡ㉹��V9������I��ɼ����SZ�&��*%���>3ւ�%�(%d��|`��AW;I�oTRIu���z�p�*��?���*�Y��6���LG����!���60�f-�8IР�S�������~9���'q�9��I�p!��&G�5���{�߾��0��`_}u�#���+�Wk�o���[��|��v�)rF�t4�V/���j�lؙ����}|.��3�T� 	��0�x��h�h�x����p���:�=Z���;�oi�(<�;{�R�sbξu�mZ�����$���W����1���8�<Dq�<D0� (�#$��`�<��[@k�2������J�9,�p.�N8�\j�lQ4�l�=%6B;�J���<�}>�I���p��;�>Ô�|��x0��{hz���5��PͼV����*�����-�xoU�k�M���]s��kiޘa��7#��{�5�tTO��{��å�a^ooy���'���\�牥�������<�	���4���Ml��@yk�y����'�ΘbVs�VI3�	���>|��%o�?�i��tļ���͡J���6�I��{q�1����k�	��4yf�����^�>y߶�r����@�	�z&:�i�"1�n"��bw޹o���ß�����~�����$��ǃ��so�Ǡ �����3\�������WY��{��,�oݚgp�LՓ�ʽ����C��(��@|-
�}�;�z#^���n��<�S�xp��n�,R���נ�@Pߘ�<;Y,r����{�c��̳�o��]o"����������^yU?y�+ ^ ��L�@~,gUz�`{m��g��=�Xa�~��k���Um������q��T�I�o=Hh̫���ni�}�&�+�G1�/�~�Tb*�{���
����I�$�||x���Н���(�,P�� ��ƞt3F�1u��ܔ�ޫ��f�}���r�Er��80@B��{�_���"! q�<x��<x*���� r	"�<�μ�����#��*<�5-�{�y{���Y�����Q���̣��Ҡ��^������LvGN�v�Y�x����aK�P���@w�801��������>V�����9�#��좱��:�	��|�ؼ7��b���	�>�a!-r"<��V�����k�&��8qo��mj�`��@��v��Cwэ *��n
y|��_�d�/x	*�/���r��-�X~��yC��?���㟏���m\<`=5�[ ���K_���6� ���D�ى���{7�.�c�w��}����Ψ,s�t·}�SlSԗP4,t�mGk($���7ryp,�fb��HO��<2}���S��R�f9=y(��X�i�����7��t�Y�8$���Ĵ^S�M~1���@f��s ��"����I�ٗ^e����p��^��5^�{�Byw��tc����n`2�oDn��l��x�V��<���ý[ &-��eΩ�̂���l[�W�!-L'��F�rhkή*�xm'�1����p��깘�O����
�4�;�_wf����]l��i�^G+V�wM
A�q��˨7�;B,�WS��'���kz�E\��36��Z�.=���˾o_`��?�"&<cǂ!���(c�<xr �"���+v�u�#��a)���)�A���8�n�z wT0���5��^�_�Ϝ砳�mpj��H��=���N�>�ܭ�~\}/d_�fe�0_���s�w���� ���>;��-ռ�T��]�.�Uj&%�"���}o ���f��'�~�^��%�����M�O">��Y�q�\d�W��U�ְ�����ΌL���=�<��~��fu������i����57�g8��G��������6�r�&��ĶK�oXmhi#������zY�ހ�=��Zy�Y�J�<x-����(�	��Xd砞���H�p,7��)p��jƴL���W_��{m�\D3�M�3�#���&�C��/DǓc^�Z%�>�� v�H�ҷ�y�C��ik��=���6��;��6��Xk*ׇ�Ɍ��'�>�O�bƹ���硞��
��#<�upL]�Y˿�w�)�&)����q�:������{b�؂�v��v��<�g���I�µ� :�cONȘpil`�ǯ�O��r�L.��CL�U�,+T�޸+�S���O/��g<����wsרʹ��eZØ~�1){�2A>|���E/dIY3=�����gGy~���֯��W��+yF�H)^�,�2�����ɋ3��oWq}��]�	'� ?�lzx��#���c�<x�� q�<x�""���� �:Ѳ����b�l�}���ng$K=�,���}ί��o17��G�Y��z�έ��e�!g�wY��PWE¬v��7��f�7\y�?�ԻFlb[�����d~�������#_���V���`z<�]�b��k���l���ѫY��&�qf��S[-�y�z�y�
[�"�&��0��L80��΃�?g3ڈ�j.�h�c�6���P���B��9���(�t�s���-Ň�<Y�T@�|t������v���L[l35uP�~oT�o6@�^�~Ny�ci��^������<��`3gu��~me+Z�Mi�%�qO�����*�@�@?��_I�O�Nb���4�1Y�y۞q�y��za� �!�ї�&�a��4���f�G+���'ާ����`|���Q���C#��=!`�T��S���1U���U�o�{u�/7�v0�ũ=�/�o�(�0�o����F?�,hC��)�%ێ^�*�q��&%��#�~�<��@��)'�/ 0[L���P�|��TWl�/PpяY]�t�=�����ڽ"ߍF4����6�Ք�P�	^�~~�{ଌ��w�����<�kf�	���6Ҝ���L	�A�1^e^���y��xl7�rg����W�����x2�i;�-���ߨU��J��w�h+Q���@�b���˪��Hcx*vOᡭ\o,��(
��R�����C��\p���}��'�o
2�h�n����3�E�g`��k����h?�=�x<�}�⫏�૏������� ��"��y�����߁�����_�5�������a>��pb�f��{u�1��]��^'洰���Qm�eà3f�@X�#ܠW��>676�A�8�5��{i�^�z�0ŭ�7ڰ�@z,n-5���`{���mf�"��/P��΃�{}��BO��D���M���崣��3=��7݇��mNl����!w���D��`9���|��;�B_'���C��s?.�a��&�=���I�nY�~�$�צ˳e�0���
3����[8�r��Y��KW�,�C&��&v8�Z�������U�ԏ�Q0��ߎ�����nop�N����0��� �y������)��r�mGs�Pb�L0�xc� ����z1Է��(w.�������e���"��UoG�X;[r��qe�gh��䡸4E�9޵�_�>z`)�դ�~8@��O/'��_���8���A`�Ύ�o8Q�d]���<�jznʀ�d���\0o��Jl�D�;���?W�����4�����4w�ԕ�ɲ�+mS�i�9Ya�T��.�V��S�Z��V�;Y��-z���+%�M�x�YK|E��^ԮS��}c6w649N��RB����贺�r�T��LN]�շ�3����^ <cǀ����
rq�<x��"���)ﷂ�u�p}ִ�-/>60��ׯ4�C���'|��@zc ���gަ| ��{��lc�͕|l =����n�f�+����cH�kG�����hc�1U�����T�ގi3q;uǏ������l��L����tX���7��������$k]<1�pE��ɣ9������b?z�v����|��[��A5��y���o��	��={eLz���_^����鯾H4�M���/��r���+�����r��Vׅ|�b7o�k��ijWz=�ugof{�zяv���������0��
�y��_���~$O��+�����nA뽖/^:�)k��h��'���� ; sr|�������P�jZ�|įP��ۘC��<OfTO�7up,3̘���}�Fu�k`��g]{ös@Y_#J�`�?�����������~�Gs�3��n7�g>g�^�p,�o��~m�L[Ŵ�z)����ض�� ��s��F�%骜���\��uǣ��%��ex}g�)O�*>N��.fۻ�|
2�.��2�9v�{x�=v��7ks[�v�:�TH��:��h�w��>�P���r�Q�yun�g]q����T�� ����p/��-նiv����]t���Ǌ�t+2o3������3r�Wa:Y��i?��u�ODx�< LxǏ\xǏG� �$ �-rL%ݜ�f������S!��"�� sG8�P�k��^�w֖�5��)����R�\�i(q�)NC����Af�y�Y���(�����Ì�$��ھm����ٙg�+���ri���0�������+̓�����#n<�|�������qϡJ��חٸJ��X�^/������v�g�?�j���Ac�R>���<��vz��<���;���7T_���5��sV,o\k�T��	߇տ�4D��JU��korT��&'���r�1{��\T �������Mzǁi�Ny��������=�C�vgp p���6/���/�a7�4����p�	�1qL�FO�' ��k8WDv���JwN�=ډ�B��ߔ;��e1�B�����7�*��?��s^���H�۷�o7JɀL;հ,He��7 ��z7 A�0W�~@�>@}��GN�Z����"$�]�6��x�iڏ���<�!�5xu�L[�� /�O@R�a!�z�t�k��	@����MQ-�u���f�t�Յ���珃[0��ʾ	-5�c�;��6�4�G�U}x��`���=��4wl;t�v���]w���pi4��]���;'b������/��{����-�z���8C����ׂ��⣏���ȇcǊ"*P��<���Ϸ��wΏ�������I��_t���ʽ�A��a�W�҄i=�R�R�.�,yk_��S%�a�~>pT	�p#ӑ����PF/�~�����f ���ߨeЩu9k{Wz�8��/^n&�35x'^�N9d [@dU���b�,`���om:ٔ�;��D���ۂr�v��W>ɏ��O0�~i�L�zߛ}���u.��nzK�����d�q�F��K���0c���_���x_yA��å�,�r�q����9mۜЙ���U���G��ܚs�H�C5zټ��E��g��ڌa-������x���H8~g*?�I��}�I=m��̚y��	�sǆ�3P���j��θ���:��"ow��󿢓��<�s���4
?����g���8�d�n`$��t�����|kga\��p~j�x6n�����c=����>�1�[)�����G�϶7�ф)�*^�6�Yⱷ�Y��{�$�����Ԇ��X@!Ƴs�{~�1�(>j��o�ݯ@nG�z�T�\� B#���9O=T��U#_��ោ ��÷����0?s�`�dK�F�5İ��v'�ȣ/C㹊�|b&���zMw咥7p��6��@�rQ8��o3|8��:��y�N��rW�4����
sCy�ϓb﫺��7C;Rq��c<K�㏙겏'�3ia�O�s�����?����
��"�� ����<x ��*H����ۧ��{������#2i	�7��^������Zی~?Z�6���m;�X�+��'7�z�1��wnb\3��	Ƣ�ڄH��KN��|����?��u~��f��I��o=�/��|>~�N�x����}(�`�p}ߡ Ak��r�3��h1�9�n;O=��s��;H���@��ǤV�����C��ߐ{ǂ�3m��0�x;v���*ߖQ���'�߂�θv���^�����}� Ɵ��'�>���*Ơe��l��X�7�U���
�������ナ�q��r��Y� ��� qS:ͽ��z��S5�3�M�Z�����N�耥�����🏟��\o�Sg��1\w7v:�ƙ��J�� :|�8�����Ф����'�\
g�5��c��?�������*\i�'�Hk{}���ս�g��&��Q���a�~�]�W�9�.;ݼ0����=�<1k{َ���{W�
��}�EF�'M�lז�s~m�O0$����_�/�^�B\�D@����㟋�)&��⫳]N�B�^
uKK0��!��Yi�"6ׯ�z��Ko���';�cw�R|]�[ԭ�V���orK7��hCBP���;��i��Б'��Y��[�)���Ю�Ӣ9�7 *��D����E���U�۝� �aէ]9��ﱛ��8���Aypə��>�ΌV�bNuv��x��\�7�z��GWu���VH��"�k_w�n�i��(�c|u
�̻\ʫ�2,V��/��Z����Y�c�C�⚳�;�s�nz�X��]�n-8js�$�kg��L�c�;�tפkY�C�,���q�o
��o�KmS�����%��U+>A�y9���3!F��w.T�KjAb�8���-�<�S*�.?�#�\�Y�����ݢ�3�뛔�]���u�1�ǁԺ���u�ggN)�YґZ2��#qv�2nԢ�`Z:
*�&�D�Ts��OA�M����YV�Yˍ��B̦�3x+ʠ�fXY|�G�Y9Ԡs��;�h��am�]d9�Y����,��.X�$:�;��՚���B�Ut��W ��RNS��
7S��a>!LΛ���)�!9rXvΘ����v��1�d��J:�˪ŵ�Tו;J�&S�����K�ar�MA���|�=n'.�g�n�fo���E��(�BA�t�q]��0�?�7��aY'��o[�S��A����V~�]8��b!}��]ځc�h`o��Z�j�5^�dK�>N����H�dKL���d�sf�x���zeC��3fL��Z��:���v6�莘�ػH=]Iy$��j��EKgem���;X�s)��<]Уz<�\��˃��S2fk����t�$�o#0esZ��p�h�ð>�5�J���x��]B��J�e�̐�����:cx�rkL�6�̫R��t�$M'{g��J���7��)�]��p�؁-<�탗h��gU~��Y<Ά�Ţc*�P��3h��j��s��ׂ�m����VF��(zgl7t���{ lj5���1)VX%�]a��̦�r�s!��a˨za�;}���ǻ�Ѿ�u�:�����d��Ut#-S��k4��"5*�9E�|T}�qjR�7���%����I
/�{��}Y�y�e�eY�24A�_rS��-Iڸ�=��ܡ��/o�ͤ�4�y�{ΫT��m)k�ׅe��үb��t��,�;��N��+�wwq�TeK�u!��s�b.츱��	|0���v����_p
x��b���,U%j��h�[+YR�6�����Iy2��7�S!��9�rL�<u������^�ֵָ�k_������<~{g���=�2����X�%�Ϸ3Y�W���jF�ry��6L:��|�x�����׶��5�kZ�Ƶ�����O<~z|<��'���b��F*� ��*���Z����X,��_��t�t������ֵ�ֵ�{kXֿ?=N�4�<�����Y�j�s^�B�U\2�(4J�ývUXD�c#��9�9�8񮽾>�5�k^5�kZ�ֱ�k�Ӯ�?O'�b梯�����+FV���mTjTF�+m��T<)^�iDX)�B?���bhZ+D����>qC+"�Tb���b�L�{�ĭ�T*�0�k���{"'ԩz�F�j� 1U���X-�Q�l��S�feT�(��`��l(�eDT+dEdV�{O�g��)<T�mZ�*
Z�UU-*
,F����J(�Ղ�(�Ŋ��
�QY)[<�e,Ucm[j���a�Jޝ���͆�7�r9�2���S���Ͼ�fΒ�q�,���t�NY�Ւ�Jo�xx{������c�<x(��<x��'cǈ��`jH�\�@�p���[���25C�I�e�0��A� ���>)�zu�t=Pú��fDΎE����Շ�,:r'��:οMH�p�oXXs3���9ϟ�����U㳬'���r�)�TuŬ<v�H^�S��1*�	�p����|� ��s���v	�����<�#��l�1�\��zjU�,#��XǞ���o���=�?���/؀�#'�f�?yw7[���dDw�����>g����9v��=�_�V��K��$/�ЄsxGoa��G��C�̋��9�o�x��k�5"b��;B u��Q��n�-����7�����=���1���P�&�;�2o��'�����KGy������$w���s�v��G�F�T#�F�z�uvX���ˆG�3�fI����~_|�yQ�0�y���g��v&��먗��Ao
������Co����t-ʯ���Q��v��>���>$�C�/��ܫ�cB�zg��y�tG���R�ˌ��S���s� �^90'�}�χfՑ�Z�%ڙ[�	^p`��a�750	wR���O�<���׍Dj�q�y\U�I��S�g�'@��!1������W��_X�����kk8����ԥwr��h�n���:��gt �Ĵ�;��n�u�����XU5��p�<�w���{�_����ǌx� �8�<Aq�� ��[��o�����$��O�:��������)������<-C�4_�>�H��G�6{�Ke��W9s3/��r=�h��4S��zFGsǪ��,y�:�t�;��Qyɘ�������P��o3{\�D��a�����^��#kW���O͍�ܶ���noW��y�t)�y�lEX�U����;��/�N<:�@�~KA~�c�@a����P�ڀ� ���s���fn]�sNi�ff�6�[�Ź�����s�13 �	�s�j��.'�c����{�&Vquw������:>+l�H3�Zo�C���_���Dw��[�Y���ؖ�s��Y^~��܆r�M0T��C  �>�:�[��������v@����3�<��A�8�72E��Q�*���a���C.�a# �@��~Oc�mxWeMx���cW�]��4��VA�f�#lå���\�~@/J��@+��@�U�_K�`�2���徭�hT�����?X���̢y��۹Ϗ�'Dg8lu�]��2�q��sy6�?���� &E�;b��܎�ɳ��l�~Wj��T�K��SSb�{h�*=�.��pu��tӖG¾��Y�NgvPBWNv��f�����d�kN6Y����q�3�'c��u�,��ɭwu�vS��\��S��&⭞���O"����ȣ�<q��c�x�Ǐx*r s�o�}���	M��̶,iIӝ�y��vZp��,s�I������z���������`����M�̷�M/6���+k�m�C���w����Њ?���~���E���� �D��D�?,�`5������
�C�>��F� ~$���K«`n���~V��;�x�!=�������O���.�q�H��s�s�w��տ�~�˯�<�YpږӁ8�>�1	�������؊ý�|�[�8f��-�א�)�0����O�L�`K�3�+���-UԞ�(�k4]�*i�"�:aG	P�S����[�=�\��}��N�1�M�Bz�����s3�'���'���$8E�!��?�e+4t��8���O��*�y��Zּr�ʈ��Zp��W��g�~�Ҟv5�����g�=�F��$dg�Sp���t�����y��f�ڰY�� Ѧ�����d������شc[��AG��c��%���~4��K��ߴ�ɿ$���j����l\�E�t���]�Ǟ�-�pQ��OIy��f�\S(���lw�no�7�0�_�� & �4'ìdsH[��a�đ� ��B�f�虜�5���_l�R�M�o���7�Y��{{z�E#�j<0㺒a��{ �������Oz��(�F��<A�>�:ޗ�o�'����E��/L�[�V�S�=[��dm��c8�6/���r����T?5�ǂ$x�ǀ�x��8�"��"'b�H������ظ����;�'��Q�`%>��W�-���@����)�gakDpv�f�]՚k��8�����w	:>��:~���P�Y)$}k�/5������Ԅ�����i��ke��̼D ��x�,�Pᾏ}��\�_�*@M}a�����`܏H�ju�a6v�n_��zq��~x�|�N��Ɯ�Xsa����Ӥ��Fk�(5�ʌ����立�ư�ܩ{^���M"�Xf�H���v��(>�g��=0	�3`�F#��2�**�^�|�,��� T={L;iظ��x��8�x�Qw�RL~	1�zp��)�����a�M�و�gx�}~���א=K�G��A�P��Q5���C�[���������{�5G��"%�>zeςn=��u�ᬙy��������ֶy`�E1]׍����|��p)�8��a�����lp���-uǊ�8�2ܷz���l�q��nb���A�+�5a~��0y�3j{�k��-x%r���~H*�=���M��~2Q�V�[���	`��u=��c�eI�-oh�ru-_%�f}n:g2�1g�k�N��V
I�f*�|$tfv�c�����m�H(_J�;���;��5�ǳ��tG��>��Q�8��x��<x����{�~���^���J-�TI?~/۠�z�~4�M>���z�%�ݽ��0B�8����^�=������8�V��,��w���'���98��0��S玣4�є#���Ն�Y������llb�K�#�� s�����3`O>w$}~
DZ}�Ǫq��w���L��Y������~����l|��x�G�~L�V�n�69q>���a���ru��I���?}��w�)&Q ��%��	ü�O&��4��tw�����<5���%	��g][�Y�Wv�k	�k��
xo*�w�[zˎaߵ@sG�gz���Pޟ{X\���Rt�6��eoM9ڨߜ&�[Azw�p���d*�9�yvK�A< ׌�u��Rv���7N�8�À2ㅘ���0_Ǧ-���ُ��B� �㾊!ד��f�T�0�]+s�Ҋ���w�Q��,�����s�Pj�AN�������1��;��Ƀ�(�������j�b�v�s��c4)���z|�ז��k?��X�d_u���1oPŰ�����"��wd�ց�Y�'Ete�0���37��nS�B�++(�sgF7n*}y-������R����si#��U���;��9�/V�R��X/y����T�9�)��f�WVu7�iY��}������}�w��� O��� y�8��8� �8�UN�����wˏc��,?k�B{`��ۑ,�����	���9�vk��Y=�Ȩ�̼�E^P�g��G��Ͱ��!�o���!9ͯ�Yj�Z
/� ��>Q}e�TU�oY�{f-�����=LN�֪z<���G���!����ς���/��GD�^��4���;*B����~@/i���K��P�����8(|���m�ʌ�����~����ǳB~-Np����Q+(#ތ�яx�CM8f`QM[�a9��S9usv�o`5�%�}^.�ޡ�M(@[�:og�O�X&�w�Q�9�jg�6DVmy����y�r'&�Ѹ#���+���C���m�h~ el&����n��ڜ�E3�wW0[��T��tݗWV�5�Q���\@������hl���nc��3�������=�.��ı�
;����FGW��>>G�B6�Qz���ҼE>d��k�b���;8����e���+yfc=�����=�el�>�y8�u������ pqm��0�{O�]wk�\���a�j,`{l����4��Q���/iK��D�;�xZ��}���%�r5R�.4rW�����
�K��b������D�qR��-�<��^bu��`8�u�&���3#�����rv����S���ǋ�H#�<q�x�ǈx�ǈ��
H�w�����6��M7��OgaY/ ���}��CdU�=�;���\�u��`E;�n�hoU��γmg
��1]h�ڍ�����\A���y2��K��&�.�z6�`�ѷ��Mݹ��fn�#���ޘ���U�MS��������������׶��NXU9s ��㊊V���B=���͐�n�QM�"������j�/ۯ";���~�W�����0�ṗ ���>2/��f�\z�����y���n�	[7Yej�(-������T��jE�n��ý��0�a�|������r��/��UM9�4��}�}�fs5�gsx�o��D��o�������sE0~�H���D<�����m��t�g{�Y��.���<��x���鶟m���c�qbK �L#xU_]l!�06OiD�v��{��,%���۸�&W~�{�� �L�R��P�׆.��3��.)�e	�7T��G6��v�e�{�����c���|��gH������N��Q���L�P��F6���Ƣ_���N�v�8�G8�"[��Nm�`����1�A�W��/qM���NP�]0Zc���^t�;�s�ձF��o�ޚю�������I<̄)�3��+!0>xG�*骭˸mm�x�T]��E���z23��|�]�;��8������Φ�%�\��ʃ��[��?���E�8�C�1ǎ<T�z<��xa��zs��]����彷��E�]����/Я�����=�"
�H��t��:a�ٺ�K��G✟}�t~��6l=�&ײ ��� ���"�@7wG�C��A`��3�"���4N��>fk�pRg���Θ�`O`n�����y�y�N��y������5�����_��������Y�zCp��>���4 ž~X5_,��|tv����^����u�`�ח�0L[����P�c�
`�9�W@	���&j9��m�0��u�'�t@L��[}NmZx�75=5Zt�v�rBx�>��<}�y�_/���B?d����@1���¹}/ϗ���ⳳ����\��\LĜK�
x�|��|����F/�TX~���}��8��C��}e�]�ŗ	�<gq=�����\@��^���A^�\ǯɜ?04~Ydz_̣{�����̳|�aq<<�%���2rgXן�1�=�Zᣌ�v"_�#��oj�Xw�Vp� �@d��*|3S���G����v� ����31�O8�4	Tw�[��5���V��Y�ި^���� �j�T�J,+0�S���掎��vZ�S�Ĕ:AE�Tǽ�\J�����9b�jD9b #����9.ܺ];��aF�X'���������=�|ۻ|ٙ��?�5ǂx�ǈ��� Ǐx��B3{�Ύ�H�������`03���C|����7��U��ϐ�xo_�/��>ǚx�ʛ���V�C��u�Љ��F?�/v&a\���8�/��QM~�*l�z�C�l����#
�>��]�1��NT���gĎ���o�c����(���s[V���7-�6�vvrW��9���6����鯹{�B?*��k�i�+^~i�d�l����8�Yhݼ%�.��@�g��T7y=4N��I�ސ�͵Qp�Ol��y�>�Q�����C�&��w�j'	�ϣ<�-�:���}(�9\�����v}L+?p�eC�}��o[N8C�K&!���S�o`�Ȯz�*���b{���mY���&���'���S�����t�@!����Ǝ0`u�l���$���B���G��9�g���R�Y�ꘟ��TA���Q�PU?]�C��K?|�������sU�0��z�cu�tC�^A������m�}���L2IC�#q~v�!��o�0�r��������O�k�A�h��5�����*E��m�r5��חGJ�-�ΣȂ�3����
pm@�� ৱ�L����s$$N�y�'�������,�u��+}��!y"��A�8��ڳ9�����
�q����糜��@���� Ǐx<q�ȸ��#""�{m��{��߯�a�f����C�Z���{ɠb�p�>:�7��7o%����y}V��g,�%|7|���m33m({��A��z
��c^�B�� �'�l��>������`�Am�YA���O|����K��ƛP2Z�'oP���M�k�P̀�D����f㯮�6�u��J����-������_\d�+'|�/�� ��=h�*&zK�+U��M���\�8��W��?�|���|Q���HT�Q$�и�|� ���=u�9�w;��<WK��c�|o��B?��'�U����~�~���'3�}�?��{��g3��[���u�+�x諒�ș�	%�SS*�W��|&Q�����Ы�{B�lR�;WVa���n�60|�PdT�O�p��w����m>��������B:_fs�-X���7'��^������g��)�`�� �ucʳ-Q� Il�%Vm=w��P�[��m}�g�F�&�|kAű.��XP�EWl�;{���=���|���~+���e-9},�hZ���%,gLwDm'4��;��=�-qm�[��XE`�gZ��A:[9��Β����ؚG*�iu@�o�$�n	B�6F����p��.�,DM�]�{b�uZY�[���A_�3&�����;n\ɉ�LH�f�v�?�n��-��w��%0���`��b�����{X�S��}��L��5Ư��!7�fG{���P����|�v��ӵ��u#���H��V��������ɼ�aR�]�%���膃؞�fo)�j��N*�:,$,΋wJ�E��LV�OD�1]qrv�}�愐�(ui��s�7u#[Z܅6Eu��d��S�����AL���}�Bm�N�V�/q��[Ó�
m����8JP��n�a�;�z�v^v=e�uo�w��tE�O�Ds�]H#���:W��xﷺj�8�F�ic��tk:1H���c�g5
��bs��X�sqb�P�Aڏm��y�Ko����UwG2�nuG;#.�'� ��\(��m���;-J%��˹o0�Ӽ��M�\�0�u���u	��D繙 Ysa��+���fFA/���ȷ&�|1����8�<3� �\_�t5�t��?'{Yw��u�䠇E.J��Kbq3DY�!��-�0�T"�H}�}����9vA�Ge3y��#��}�_E�8��!�*�[Ψ��ۨ�[+U�6�8�2Y,�W�K��Bj�|�H�ucZP��DEH�P��=��nݞz�Q������W%+��a�Bo%F���'d�XU��i�M1�s�K�
�q[��NrĬI[Jؘ�8Ma����G�;K{���5�!r�>S����U}��:���V�li�i�F�-c�6��tg���f)e��_2Xޤ�8y��C�|6�h{�A��J�k�G���4�q���堕nl��J�ŲY���(�h��fZ��#:�M|��#3y�;���N��w��,�i%�N �{d{�[����v���Q����v9GX�|ž���l�Y��ܥV�${�����Ng+ś�\:)�%�ҏ;շ-��N�8���%\O��e�[o�bf�+
U�`G���ef�w��o0��p=�g�T����h�.�Vr��$B���0�����Z�K:��`8Ư3�a�(��W8�I������A�s3p�-�';yϫy..�gtQI��w����x*7��3�*U��<=��OC�W��ѶҠ��'Ơ*��)X�JR�HdȒL+Ǐu���k�ZּkZֵ�cZ��Ӯ�����a5�*���+V�V�AA��U�����бb��*�3��Ǐ����??=5�kƵ�k^��5�u��]~u��0�3��_hUM�H\f��V
+(��X-k�D���>����ǧ���:ֵ�ֵ�{kZ�Z��Ӯ�:��0̆F2G!��J��?[�m��,�"�F�z��*}jamF�^�=�ק���ֵ�u�kZ�ֵƵ��]~u��xF2d	&a�!1�������
�*����F�j���lQ�l����ږш���d�Qu���`�*""�IY+-mTD�l*DJ�%J�b���V*�9X�f��x�����TUTX*�S%|-�1�~��j�0��ۓ#��
��$���*"��lF�=ۓ_,D���U�16�`���Q��(�cl�".>{x[��W��pۗ;'n����]/kήonqI��:�ܧW����۪��y��6{����ok�8㓕Z�qݎ�F�����iz�#�g^M۸4}�%}%ϳ0ǳe�At���]w�ơ̷Vb�o:rX������\�o�JO��i��"PA��)�&nk��獊�g�99:7�o&Js׭m��wg��c��b�*t���V�7j�[{�X�2ֽg[m��;�^��*�ww]LkD���-�+�y�51�;�u��wp�̬j��r'aRݞyر��˸n��v�N����;ۻ�#�����Үwv6ų���x��ݻm�����f^�{Z^Su�ƽzrp�p�?�����G�x�<q�x�Ǌ�""!�����^���n�������[Vx-�K;Y�4�X۝�Wf��s�r�whB�u�`��H	�<֋�-�U�_D����Ĭq�)�"D@��ܯ�q
����TC��v&�=�*<�6O�#��=��n�i�ͱ�R�7����JX5�7�Pg�������@��槞�!�=_N05�/�y�w�����r��/������_ �5p�6�4����* &��5u����\�j���<����פ��Z�Q�c�p0i>�)Ŵz���?�pq��8Ge�_
�ܽ��}/3�J��s���?����b�:�c�-z9���"��š��\��ь7k����B���;�;����Л�̉c1rK��ŷ_S�p�T癨#~�`�<i���R��؃���a�@�ns�z�34��2�ق:FK=���3���sOh�t��l߯��C���@��Ɇ����-Ņ�����;\�|<<�J��zjq��H�g��>��tp�$Bv�9��O�g}9�e*��ބ�ߐ�}/��������i��4\���%kz���s@�&Y���3��2�+�A�]iG���n�c�Y�5 ����f�`y�_��,�[��Jˊ�	^4/�0�C��t�U�wj���4";v���ɝCBK� !^#����گw��Vq�4�R��J�V@Ö��S�T�w%s�:�a�����f_o���{��g��
�#ǎ<R<x�Ǒ���8�@9�~�˳@o�7����Nțt��p�0�\oVZo�^Xza���g�묧}�1����c��;�^���:�1/4�ɜM��z/l�}�Y���៹f����$�m��¾���/!�m~�v�"�8����H~�S$0�}Nv����'�Ќ�ɨP�V�ӛJۅ<��=k�G���t�G�>Y���Ҟ�AG���5�k�5�k�Om
�7~�l흢^��a�������CC���f���L����t�*���>ϗ��h`���P���kh�ج9{�:	�<���c]�9{�W���]�a;�7Y�٘?c£�t$�Ϣ��K�wW0�a��7�~z�>W��l8,�x�+��pȫͼ�;�	wA�(2:�ў�	��鹏�z+�e<��l��g(��P\�減�1���8
�����
���(D���_�N;�@����n9�JU������|����S��.�/�;�Tv9c1 ��P�����X��w�z�����#�1���.�"�,m���K	S-U��-��˗����i��}�M��*�:��c`z�´�xa�zϳ�_[��O
n��Iݫ+�i��q�+S�iv�jҸoZ��g��3��1�ܻS�Uw���j�_ǻ޸����8�<x��d�����D�Z���ȉfx�{��n)�G��c�/4�g��G����ݞ�h_3�	nD����4�Vo�R���5��^�i���AX�}�"���DG����ȇc:n��I��fmຠ�M��}��޾'��?*<@���89��[��0��UD�(�����`s����X���_�W������{���.7�zc�%�g7e��ݽ�L�lwjeS�+�|0k�<��H�z�h���7�A�e���>�3�?7�/���|h�l�G���(�0��6�����I�MG���M~�Ič|az���Y��W�r9�7���1�C��:���^�I��`� ��>�h��{aP�����SG\�0٧��Y9�/�]@�5���c+P�~�ȩ����!�>�_�,4�|l�f�쐪*�GWf_1%�f"!�~���O3��}�O�n޿GW����H�GB���zkj�_	M��gX[�T;�oS�7��~�
�H�Ɔ�2!?2���}�k½�W����W�^���Uӓ�g!86�Wn�ӌ8�ja1���Ș �L��;����X����U�|�[��E���H�s6PN�0.���p�w\��4�Po��%�εx㣦��8nq
F�W�^�3�?⪿yy���=W��z���8���y��/����~��8vM��6���ZS<��nF���^�^s_v*"���M'*i�駇�N��E3�6X�<\�u���.����c���739�=�)�w�9٫	f��DS��O!�g�x�޽p�٩�C0�Ü�oc�H�	���~���s�ZKm=`s�����o��{� #�R6���;�.�c�V��T�i�V�-Ŧji�ΒQ��6S	��\��
=��z/nCc�n�t#�ǘQ�[oٴ+�!�ꧼ=f��Ǻ����F\��5x�z	L���2ݯ����`�ǽڴ����6qΝ]Z(�E�|��~�)�ˀT�8��1����C\J�hc�-��ޫ��I�u5��F�3מ��f�3�"7���ጛ�OZ&߫���B���h�����}��{-����f���
K�1�{�
��S�.(~�n�c<��"��Ko�����9队Ghc�޺r��u�P��>~��������%���n#�	��5Ms�U��ɫ���ܚ�89�ʙ8t��Щ�
]�qQ����?:����˶k�Фj�$�y��$z��G��s#Jf���)����jr��v����&� #tŷX�o[Ay�Ou_Lf�����:�� H���pX�8�ǂǏx�<s� ��G32ꥵ/ۗ7��C�ɢ�Eڳ�yea ����$ꗶ\���!*_B�l���T����lʅ�ʫ�}5r��9���l����G����Y�ξ�����k5B��ŏ�o�ޯgߠby�XԈ�fQ�"���>����H��4ǳ�΃f��K��
�?�DLV}^�	_�<��֩*�s�����g`��^�2�ϟ��3pD�O@��+�}�5���Z��=g�sҡ-R���(sq7�5��l���*}����U��TIidк �4�xr�Ǧ>#���Ҙ������N��Sߏ��F��j��b0��
����ύب�k�i�����Ɠ�;���|�F�	�\I?L"ܷ_-"�}B�z���t�=N�c�k�C��716y"E�cbʃdK?����;�0fO�"�xtz�"!�6��k��uѫwk=���xF�Ru�ڟI��&�{m	@ձ�׵�'�+`>�h�ף^M�vT���[oAaԠ�U7��x��g�&z�����o��C������&�#q��g�0BI$���O=��_���	�#�{}�5�k���y��^�l�3�w�2%�l&3}��#1�:��UP0Ԍ�Q��KnWš�/m�;�k{G�	�xF
Kv5S��k��&�U�`^��;(���__�NJ�~j�El�ĢkO��X����i�b4��|^��mg`���+o��E�2����S,%���l�|;���{:��O�uǁ<q�G�x���rH�<���߿u��a�8k.%M�O�P�-��b�Tt���|�<�/��^�����~�㘔{��d~z�`�7�<A���kܜ��������m�6��U����\�YwOSOS4��[�P�{��0�`&���$cK�
XF�:h��:n�V�K'7}�R,͜�<õ�<�ր��f-�����Z�h�) `���Y�I�^��7�ɭ��nG��,�Y�  ���Q_	J
^�9����οA\��D����Z,rmn�dK�e�Í�C`����F/9�zd�P:}{6��V�?�O.��,�����n�1ȓ�QS���T�A>��o�>�>��B �u���\0�y�*$�d>��:2����H�~�{>��
�CTz_Y��z�;����x��OT�����p#���͌��g2{���fù�ӥ�2�F�~]j�9��(�~v��~a�����DvnX�E@5кu=2mY'��>1i��a.�u�{���=�'ۑp�>�X4<�cGvHw�dyy	�� p�}�4��*��g3�<_�[�~����T5}���vM�E�Y�.TW��-^I\�l���U��`�|�G\�W1�fR����d�� ʲ��3�n*Pd둳B]�Z��^^�ڷ���o:�������<x���qǎ<cǎ<Dz��?~�q�ɲ�2����k�\g��'����|O�Kя2�]^ԛҌYv���:�[��1����9����02DG��҂�-�sH��7>c9��������a�X�&�{tc����x1�?�(9nn(;�жm�ʎ�d, ss��)�k���[�l�w���Izga�x�_�6;���uy��U�[����ia���ϩk�]Ϡu@�1N��M�80�d�\�Ǳ���~�c܃�s�m5v|w	�a��TT��=26!�0��ׇx�[9�x��|x���UT�5C��;��.{�B��F�l�8Fg�����^/����"�"�W5��ʎPn�Z3���{��mہ�O"������,���A��r�����K���yr|m	��P����/D R�~
��|���*Q������t��9�z��;�Y�?{����3~Յ^u��|�����	 �����%�o�|�.�ʞ,�*���g�b_i�{�H8�6���u��f\־m8��J���f�˧����f�7�k�)>,^b�;���^�F0��AER��ō�Ʈ����w9�g}�,Ч{jfީ,�o^s<sO�ż�}Fe���l�U���=�8����8���8�#ǎ<���I+�7���������lK����Q&(s��_|��P�_x���[�ffً�e�>CE��'��靐n���٦�:��>�ԥ� O�q	ߐEr��߶g^C��V�����(���|O���,��SW��<�\��dri7��nmy�+������8G0�2�
���ձs�W`���.�\�!�ާ��t� �[>��B�
{�]��0�m�h��q
g�i���'� rop�堿s��D:ilm,/�ǫ�o`�Fm���ܲ�l��.��uv��soޗ	�. �oH���<�D^�*|k��z�KwS�К�}<�g'��-q�ֳ0S������\���#|s��4�%�{���4�`�4=�4B�f�*��r�:�˽2�G+����0�w��^�|�+�Sw��U�z�~&�1oa6�tiyjq�u�����ﾯM"y�P���Ѵ	�<����=w�g���7���7H��xH
��?�����b4�2���p�k�l�h��OƬxO�~R����n��d�Q��,&���`�<����(�P�!�Y5�3�k�>ZV�R�̨N.�
� z�_��{��1�'�L'9�3$WS�>���L�}\9/�8hljQ�Εs.����YM��w}�������<x���8�#ǎ<�=�_�ѺK�u�;6�[���YN��ocG[�8 ������
�������k)9L���N
�n��ҹ��jnnUmq����I���j:�e���]%
q���|�m!���;1�B`�9��\rz���>b�(��!�Ym�����5h�L�f���t�4��p���?c��w�ǯ�0�v�����#��=(�.o(�;�nO|>�0��+��Fl��T��đ/�!�<��=�v����=<��N�[�q�><	~�1�#��i: F�S�>VP'�$,.�g-����LP�{�:�v��v��p�g0n�ϓL"[}�3��E��ܫ��&Uz���">~pO*5j��N6,��.#g-�i?�z5��<��]r�6�-3�^j��u �3���0�R�W3�7z��w53��Jj����{@��"�zl��I��x-�nݢj�s�����J�p�?.f
m��Kd����=w����`�X�IIo�^�z������nq�0��l����;�VW�R���$���O�/��l3
^�d���N��\�S���Y�QLk�W0�1l$��s�0���?C��< �!� u�;�u�-��=�sr<C����ImR�8D������k7�5 ����|����7�����5|�@adz�����஺`�Kg�}Zob�Wm�̋=����=�j�o�d�����R����X��}�������ۏ<x��<x���=G��W;�Wo���_�-�A/2��t���˝c��p̽E��dm7�,v4ꭝ嫅4z=�;��&��'-<�ڔ����ʼ�Z�c����ؚ� dc7���{����?�O-�p����K��Z}}�[�;�mM�ú�/@v���q�c>8m�y]K	�2�4pQ�^9�"�_������<�pI�/�͠0���8م�����ٚܵ�fxW\[`��L��5?5Ì��1L�:FO��P�w����j�.�xO�Yض�s�]+�x�o�G���Uy��/�\F{�{�� lm��oG~�;�`�y�UW�A��R���.���z�����YM/��/>'¿�M���}7�����Ҷ2�Y��cjzf4��w�I��lw2@����}�U��Z����=���v�j&.�.$ZM�YK��U�V6]�f"�J��1xk�;���d���fy�V���C�����m�<x1�@���L>��YQB����b�w��xw8e��*�n���.�1MDG]V<4�;�@��λ��$�������M������gKx��(Ξ0wq�Q�md���7�q�/S ��#�E��3�\e�36��I�#n���Wxc"�>$��c0�W[�3!��
z�{e��\�K��\��q�� �.��kYs0U�(Q�[d�eŹ}6(QZ��Ѳ�"U�)u��%l���u6Pze�}f����J��Lb��"2q�޲zS����Y�;V1����:�Av��)�Ӕx��^�vW̩��sٌ%�.�v�x5t5�=�M�5w;��ɞG�c#�v?�k�OKI�0��m�������R��f�x�I����$2-�Xħn�t�Z]N2��Q�w�v�n�׉2:	��RG7M=�2���k���lSN�pS����D4��v�2��O�(�2�S�ܮ�-���C)����k�U�|xn�7��2-��b�hu���]�S���X����=�Z���u]ϯ���XD�y�5��c뭛̴.�Zp����PTP�JJhc�TD)��%`9D��]Ո2.�WY}�n�L$b��T�)4�Z�f��w���Kg3ɟ,���K]�D�]���\�迩���1v�r�D�U�������'k^o<�'����r�B��/��V�)l_7��4I���t�ݸ�T��l� ��|�����Ͼ�8�Z\ҸQ�W��8�wM�k��e�
�w�\�޿]!����ZH�6�-����([��z�(jJ���_�6d|j��2��6K�ΝN�<Yv	���%�ns�\��iG����*qԃ��l���8���V�7oGIj.�ek��2=��N��]���K�T�By��v�"��X����o ��(�j�I7W����r���w���drU�g��eZ=XWa2X�{x�=ӌN:]��Q�>}g��N�V�Sղ�z���)E�)���QO���+x�w6�����m�s������L���^᫣S�eZ^��Hjq&�wFBZ
�vI��#��w+6	UV����jĥӾ�[)�t4[}��v+9}u�%����f;R�t�&A�CՔ�2Ag2�'>W�e�^�n���ܥ[
�eh}��x���+�i�Z��ˁԔ�]�j��A���7�6
�b�+���+-�V�K�raa�<��{��Ԧ(DLj��0�t'Ȁݷf��e�q��)�4��`A������� �_F���-���wnŧ���YR�.�=�E�����)��Ȩ�w.##�{�A>Uq�X;��sι������$d��a=�E]h�Q�یǛV?_'z~{zk�_�kZֵֺ�zkZ�Z��Ӯ�:���H�!�ɐU��Ъ"}�E�Q��ɟ1Ǐ��O�}k�kZ�Zֵ�Mk\k]u��_�>=�2d�C;��*"�DA+��1:�ɋ HHV8�׶����ֵ���k^�ָֺ��<|<E��Oz�+`�"
+'��f�2BI� �8���m}~xֵ�u�kZ�ֵƵ�_�v~�z�
�����b�Tg�>�*E2`��y,=,%�yhsF"�1U�����b�F+�*��ؠ�D�}�y�{j��mgR�@�b��AKh��W��{�|AaV��+�
�"�ϧ0��V%�,��ښ�F�*^�F�����~
x��r����3J�U��E���ʩ�sʅsZ�X�
�*��jgem�=�QX����֪�ł-iu'�������[�8v�S%�������{���]��안���O�X�t�Fe\=HH����f+��~����({=�G�xG�x�	���W�_�yo\ﹱ)*�~�/�kJ׬D���.��Et[K#�5P�!���\����u�JF��o+~�}m�9yF�4S�:	�b�s��+ՄdD�ߔl}-��~?�pv������0�p�^N��Ğ�T�ҵ��>3�KӼ�@�xS�Ls���܆�̳j�wN�n	���Bmj��'X�k��}\���6I�m�p���K����oX�:˿�~a=H�������?�y�\y�w�r�޹n@���ɂ/e���;����ONܬ�jv��@u��bC@�����)���S�@l�9��/Z��8��[q�N87�����������v%���M�Q�w>���Y}��7��vЀe}-$��2���"���!������"�x�ڼ��LnZi"�	ӧ�u�{��_0
A�m�CB�1���2�ɫ7��y�;�+j)��T�f� �,��/ҏW���7��e_��g-�0}��u�	����n#:�W���|q�Sn�h+�[�;����oz��{��##̪2[`��ۻ�����U����jӪbY�:m�1Vj"���/xfFc�w���u�~�e;�:�z?�Ƶǃ<q�G�y<q���<��_��������?uϗ�@������-���	�3���e%zCW�d�GOyګ�!��f����H]z�J��tA�>���d� ��t��>�x�Z�9�n��r��ב���
e�O�YT9�^���}���}�p��^=^��q4��۷��g+J��p�!=�6��
������?�kN�g�52*���7!��H���D�D�����g���ި��}׮�*_�����D��=z�<��`�\�JV�ni��g��wFUZU�ʣ,�;�vwG����+���D�;�ߴG���{���cT��ϛFڮ�sU�����{=�j�겉�I�*�>_eM��f��OU�N���7�"�{ w(�� 	�&�����s�o�g���؁lp<.7�w�5���/N���㳫���.����C����<_'mK=�չU0/�E���Ok���)�5�:4����f���ZU<ǝE�fbVY�(�FoY��|9dT�a�3a�͙�zs��Ғ��ه���T���{3y����?O/#���<�����������1?���ʎR%H�͕#���W2f��7��º�Y�t��5A��ܨ�VZY�Nhl^nI��#R�4�a7�۫w�����{k�a�7槑���?�B�l4cM��\�8�:XW����Q�R�z��L��á���6C
�������w� ���gr�V�I���ˍ&o�=�6���ؽ��-��B��w�.n��Z=�{�Tϻ��ݱk�=[�J�����5hf�ޙ�o�^���{�HL�~� י�
��l�1��	�������=jr�k����Hٮ��̿2->�Zo\.��O#9��p���)N�W�oTQ����֞�JUG�Y��'�g�=j��M���hly3PיZ��v�c&fnl������^��wB�)��+&����i��*�O���c)�{z�)�gg���!�DP�M�IN@�U0ݦ/��bm�:��3j�W���ރ;�MW��R.���9�.�����4�0u�'v�k��z��+� ��82���t3ζ�ݰge�ܘO�`�N���#@�C��	��w |��1�t�zgy��WH;}��Y1E�V��*i'foe-���\��\w�W���＼���� �8���������Y���}����ok��+N;������ϯ�v���΋�qZh;FJXj�bk��l�UO����������f��~�\eh3<�$)�Υ��Xr	���@v�m��{n��tM4<ܮ"}�(�H�:�* �Ɩ�3g�4�����$"}I�\\�z|]�: ���T����(_4��(�fÇ�V���N��ƙ���	v{hʖL�W�8@�]*1�
"��s0��"}�sݚ(�ZY���d�g>$f�l���kJ�`�B/wL�]Mۼ]]�}b�-T#Mz��#��OG�І�ܖ�+�{�ٹ�<�Ω��u���i�����t���=����Г�R���e�aZ����?��n0p��)ƎY�S����*�E�� �~n�~NmbFL/f��Dl{���Ij�0��d��sM���Ж��ƹe5'a�'9�@���8,�G��U�O75q|���.0��Ѫ�K±���o1�)񗄤Cȭ��]E��B_Va�W�]�Ż�"6��y��y�r�n��r���q��<p_���V�b�ߟ<�x������}��,oѻ�592-�B��}�*�V�˨��I�oǒ�����bW���.ͭ`�|�E�!0t.��-�����7s��	X*ۻ�<�T-��-��~�#����1e�q[vs��a��a���p���(F�j�+��$chޜIL^�󍇫U�w����܆J��q���/�.�e	�����ow3��R+}��=��C�{ѓUY�8�|�N#>M��"�^��40�fr,B����r�$<�n��u�k����DϏ9�=�^'2J{�oS��S��)������5n��¶��|�V�܋���������93P
� ޿��z�$_��ߍX���:����Y-�����6Xo�{�{���m�W?��Ґ�;3�4�tT.�Ž��?#^��wvn�~�v���D����Y���Ӌ��\*Q�-��ܳ.ƉZ9�UW���}���ۂ�n	u������6�=p�A���}g�w�C����Qޑ�f˒y�"Y}�d��w)����a���r����.��9-���C��r=j�6��/'qq��<q�o�����>���=���	��M���b�^����>K2�'�����m_=�C{���5�z��4=�,(�[�Giu.�v������0�+�5F54)�K]�rKf��<K���_�x�.�W�r�ff��,���ײ84�sy�Uә�4�XZ���S��z�������߯�;5d����C2zV�Õ����&-���;L��8�lQ�yv�l#���D
��7r9�+�r9�m{�Y����;�ȕ��Z���-
s��[W��y��{�C��i�E| �m�c���nb�����J�fF�Y���f��%��l���'t��y�um2�>U!�v�;H�������R4��SgC73na���q��9]؜v͏p��^��Nv�c��=1u�X���ۀ�rn�.*���ٲ*1��#v�����g�m��m��O��&�߻+!ֺ2QU*�F�F���
��E����a6e:u�uK���]>Ҟ|����/q�FU�o+�A�����չۏt�J\�:�f�@[����N�i�sm[���˄\��ng���6�OϏn�<x��F+�͟��$O�}��31���-�$��&f&�թ��e�W����Okno^s�W������.�^��N�O�1��,���4��+��Wn�')�S�".���Z@g��>6�f�ϭ7{��6i��ҏ�/{^���͐��S�o_���qRr�Si�s\X��Xb��Ձ�*��awp@�\��o�%��,.ɳ�=MǛ��;����ף�G�������q�S�F{��O�0�K���!4�9g~ý���.�ٔ.����p��ol��fc����h�u��e��ˤ]d�,�X�v��r�c�H���h���>�[A�\�u^0l�;��8<O���}��=9ط�|��/B/`�<E����rnj&���� |_�8o`��?^�1�����wt��:d��X������T�����33	�=yzy��͊7T���������7�og1�3t��#�T�F��t�m�t9@�a�^3��7͗��/L3��C�=(��k7cZ�������yK͵��l^(�G+�[Z�.��a}�jAw�ߤ.�;DL\[������]i+�<���fӒ�gP���4ܭ��ѧm��T�s�����t������@ ?y{�_�xy�����8����CV+��q�mX���yg�g��n�%��8��`�+�>�R�i�ۙ����j̮��W��c>/n���� �x`�"'5߽3���g�?P����_������j�r�:�[t�}�Wѽ7v�x��zv���W�=#)��E���v��R8���wv��@�^��P^�5ܕt�g�������sI�^؟.޷([س �
��]��D�x�gc.ִ�p&�N�Ր6��e܁SO��8 &��nYW�ud@֍g��e��{�����9:�-b6&"%�bw��l�U�Զ�6�eޚ��g�[�	��`���nFa���{�lnS0dʁ���#��Ư���GP����ˣx�����u��uܶV_�{��:FG$�d������@�G_ tEa�%��D�v��O��#G�{��=x�ZF��p#/'�0��$0xΗ��oqd˨Q�՗���V�էO3�^y����3�w�;V�Qc�sFG������|y�f	�'��.�)��^_V�*�ֱљbJG�����j�k�r�η]�f�����ǎ8��<�8�{�տ�BfwD�QrH)��3w��~�7/���fȦ��J��r�2�BEnY��l�w�[KH��l��X9ΟCG;�3��O�N�C3�O�G�b8��2���u�s׎}N		W���I��}��j�Y���m�鰙3���# �֟@���`>�"�\�*U��z�k�e�R+�
]���/�33W�9���� �ѐ��O^�:����D����8�ѩ���`Ʌ�xgYY!��zel!|���s���*�Q�@�(,nE�yh���F'9�A�rgj�ɭs��[/��k�l y����� = 0)@��8�������)f�۴1�������z�G�j����
����o�7�w3ؽ�𬼍/ܚ�h�.��bk�@z�*%���6&�
����7�����U1�m]
�'�^�����/+�v�ق��Z�i�)|(tN��M��i���	�TҊR������?��H"��n�]�:#Nq�8l����{�1\��0ݣ�r��.+U��3/���3�G$?�ǧ�pq��yľ_���{��vff�0I����ga3�z�ts2u\Dߢ����F�NP���Yېu�Kauw���,��y��������U>�}��9ռ�'G�i�;:[8� �H`��v���R���"]��F�znOq�<Fߧ���2�"�7�5�y6�����c���v����򜕛3O��y�&'o5i.6�(xKg��v�[�ˉ����M3��l�[���,�&=:v=՝�I[ϼ��!���<��a�8<����n�'K���t�(�#f_ZX4<0���`�`�}�U2�M�.U~���7L�=���'�[�ULTBni����l�B���o���{s7�O7��[>4H7��۲��)������zϟ��xo��t��ܯo`���O��Z�I���<:�9DVg�v���4.i�6kH�N�khF�M����5xȟy��Rכ��p��5�5ȃ3���w����U��N��[��@'t�E8A�)���U�ݚ��azf�����Ѝ���4�`�jb���5a���"@��!���u�&��.�W]��ם��]�:DRK�˪q��.`��QS'�.
�x���.���cRXEa
"�=��r���YS����W���.�b¤���)�Ґ�;0��#�1��q��s)^vC�Z8<r���]},d��JE���E[9TvCw�x)��X]ִ��ʱr����`��L-
$�ëy6�,{S��KI+�Ӵ��X.��V�EI�54-���I�Q.}��M,�n�d
`�^�|�s+&��4�3���p2�\��0�;��)���r���#F8�s)�kwBK��|�� �I�=&��Zp��{���+���y�ޢD�fi�,@� 
���,IPwc#X�,T��9�P�M������iKr�7�v���J���Лwzu����#��7�U�H>�7r]�Y��ZB��#�i]�7��&���;m`��}'J��I*�v��c*���ӻv�H��c�}��T�amgc��4h����E�S\��Y���ᢏ�i6Ym���;�D���B�/)��w���[�!`[�����ȎSx�C�o�̰�"��}�VZN��=>� 
B�w�r�!�Wp���62�3).�LS�0�J��ڲ,0�I�3�ż�x��m#W�Vs��V��k��5IoJ!�^v��]Ma�Q���sM�G-���!�Ub�)1A����,��lfZ�����@�¹���[�F�74BF�w���f*\*{j-b�b2�*mꅮ�&g k��yGU�q�Q���{�rKH+�o؁�i��V9w)+*`}�}b�	�U�"�7Kl�ۖ��f���g~��(�X�f�u>��zXv�L��e��5��!�����fa��M�Z�~�I���]��\���	V+�,�'�7ًMv�k�<~���І�7r=��u���]�1��ٷFLF�h�9�V������eM��9f>��-���L�Tٹ���_�C���;1fiǸ��#nX�9�آ�>��e�/����t��e���<�.���t��<%�y��S�?S�TG��d��{��>�nd��ε���L��Sj�+��.E�,6lv�̳қ�Vښ��h��#�x��'!��UvNN(���$���˻�F��y�����{i��]�c�l�;�����(v��T�!صv�Z�)nj/�";��F�Y8�1ʪ�Q�ޡ��$�H��<k�����^5�kZ�ֵ���kƺ�����}�L=J|)̄ATU���R���F �V1��m��0���������8��������ֵ�zkZ�Zֵ�]u��_�~��v�s,ٜ�E�h��,�9��C'5�I�I�<k�^����kZצ��u�k^5�]~u��{��0$��|OZ���*�Q"1@PR
(�+��Ei*/�G�Y�x�����׍kZֽ5�k�kZ����=�u9Op� H2��#u�F;mn�}�-PE�ؿ�_�3�����&�e�!)��&K)j��9�7�	�_?�QO������U�b�ŅB�b�DX��应��f��[~m0����¯�k�#^��k�2 �}\�^.�X,�$�k*<՜�J�T��F
yi������󠫓[Rܮ/��"�{Rwy�U�������,B,D_-��y%�ř*
F��*�_L+
�UrZ"QD��E8I�m2DZ;n�ws^/���ݶ�<�nv{u��p���7;Q{�sϝ�=wl�Y��F^-����S�5��m�L�R4J�Y ��:�^m�z��=�'	��D 9.�C���Ro�����r���������;�~_��4�Zk�e�����{n�7.M��u�U�l�ۻ��g��\tLw;ׇ�wR��N3z��ؽS�l��G��y��k�Ǘ�ר�;�\e��.��]�y��6�Rܵ���wR�۹5L����/c9�����&;G��C���{���U;<�s�nKq�n�h�7�������3��3���;88�B<���>~~^cn���_}���d��v�X���s}�S]��ws&��.��,�9���x�vˆwt�Kc*��GH�(���S��/*�N����o��;��z�8ф	�Įh�ZX3\��d�~�4��ޭD��z���0g^�3�;o�A�15'���"�T�5�޼��֎jXzw_zO����fb����x��8���rś�P��X{�`�}��HŇ��F�#= K�;��$�\Ky�Fr胚~<#��~������)KA��x{�af�;�mz#�^j���nϹ��s�`�3E�8����y�*��7c���5?�ת|��;T�q���gsp���@kW/g�w"��na9�%����b͒y��3g�Wq�h��Ln5���w3�|������4d]z�v�v�m[�ު�"dK�J*l�Kz4@�!�8iq�J!��;�(��5�3�)ӓ��he��U���{�JH/�<�N�tq�}���hu#3��@j�Y���%��/o�OsN7B1Nͬ��tp7;+�=o��&�3�\D{c�//N��V^�ZЇ�a�B;c�qZ�����,dK��E�Fnr�a^��}�������؈��}�-��z�V�S8�ߛ�:�[����?��ノ8��>�mwس��.5b��ϛ��@��KwP���ئ�-��ȝ�����sS�������?k�ff�"��A̕J�mB�\2�D� #�33kz����E���3��x@]��z炨z�+�U��05�lL��쮛�ν��E�u[ Oo�߬/U�`��O f3�d@�]�ܰbڒ���H�{���9�X��xd���(�0��|����w��؊8��ǟk��Lb��iw�=j����#���u&�)m�\�u(��j%���i^z˘������3�:w�g�1U5g�%O*�khNOY2Q�@��ݙ������54:�Q�3b�>66^�W��E����[	|�z����m�g�T�>ק�)�oO�ڦ�[$����D��i�'#�K�f܏by���â���_��{�=�W�Ҵ�t�6���n���O�g{��<�~��y9,�Tp>��1Ʈ�8��t\�c���z�^�4ù�f�)(��]������H^�>�e���v�5�������o9�~O|���Ƿ\q���xǜ��#{Ou�x�?j�W�s������ۦ��+������qa��C��l�k�:{S�����Tv��u�9 ���Ń�W��f��s]9׺�ٵ�!���O�홙.�]-�ܧݺN\�M���V��(�!��	�N��ڽ֝H=�̑(����Y��[��y��BĳF� 3�]��U����jm��R}�v���ڪ��mCD�af�}��a��5ٞ�����?��s�>���<{�,�eYq��o���V^ k}>������l�/��\|��N�+[Nlé����S�CXs�wsMH�kP��9���4��w�#�������:{b�T���L
�+)����������lx�{��)�M.qNoug\?7��I="כ"�f�S�F� l�Z(��Gk�a���{֯iZΆ/u�)湬�����$W�c�m-2�o_z�d�6,>�5�8�gv�X�x�����X�WAP��6o5��,��SoP/�,���s_�i�D
8[ �{|����8�H���=�ߝ_{�<����xM���}�0S���N^���B�c���?T��㸭-��~k��E����E�t:�
�USSC�W�I����8f��"K<U���@���x�^�s��P6|�fz��� ,y��Ni�����#d���vTU��t���df���p0AU1Z�{|l�U�r���<����c��Ht������R�>{�KSd�y�v����9к�D�*�^�'�����}�Wwٍ�B��z�WB�V�dqJ�*-H�͛?~"��W�
��������xq| q��<�*�[���n%�k�U�3_��|��C(�X́�f�u��o8��|�)s��c����>c��ېñ���ڌ{�r����#Nj�����X���3
H�^�9 W T�-�y�;e��C��5���^#��Z�9��k�&د���/.�e��2����>ε���� �G�ݔ���K9/f��+�%e�ǎz��H#�G��R���ԫ{8�����l�ܖ��h��CmvSs��U�h���B�n[�+l���zm0�������������//!��C�,T��E��r�n�*r��SR�����)��L����������T�qcJl�O��I�fL.�l�pQ�=Yn���%�[d�w��G�FoM�-4�Vl4z��+T��Rv#n�+���-��FK_X��O��	�ݹ�##ڼ���;K�&L9\r�[�i��|�w%@�언3�A;2!`1�f�n0���2:6���Ϡ�?Q��ط��)����޾ڮ�zvN�>;���+>���^�>{>y~���u'�K����\�x-��c�m9�]��i�m� �ѽkv\��5�Q��X������g����n�4�a�D׻�c'��BIU�wʫ����f��Th4��4�Df�ds�p�~Su��9���6�w�Au͗�'�d�{�-���aC) ��n�Y�Stw�G��w3��~ݽ(ף���2�$:�I9Z��TĿ	�������;�)�q7~��R��v�Tl�S[D4N� �A&R��Q+%�[nVh�m��d���q�	�m���6�o;�=G��)i����VD����,=
�G�sxN���a������[��S�gXs���o�����ٝ�g;�����y//c��8�c�<�}{߿g�y缒I����l��i�}��Ꮋ.b����`F�")��z��Zp��[�~�SyG�%
C"���g�,����#�5[�e�·��8aFrm6[ۨ�K�p�����}�:�<=m�������#� Q R�e�裆F��Kw@;����l΁<� Ĕ�7OV&�/���!�O�ƅ��ئ���^�Y�������MQ�=gX�w⥼�&}�#g�r��j�e�nb��˘�*No�5�Ēs1�\�E�����V��zl���}��u��>a�V��1O;��\��j`d��2L�ff����X��i,�0/f�S#&�*s7U���ʆ�`ޒO�{AȪ��~�vvbÍ{n�x��4��[�j'��2���=MN�L�?���C���-��&�2�v�Ӿ!�*���`�H,C+Iޤ07�w�M�yp݇'_JsQ5���N�K�I�kwn� �vwG��p�l���:\�7��ՃW]��	4$i�e��έ��u��s�޻�������<x��ǎ<�8�a��������tfL�2H�ټ�:Z���lJ/j���M���V>yq��稭�aQ��t�b���0c�����I��z[��sE�Gʞg�.��*3:�V�߭���:��a�N��M��֪�����=�R�8��h�<��z@�H�[w5-�e"�K0M������N>S�O^-��6e��%��\���65]{���u��]�
�M3�;�m��U˝��gU��Ch�%D�VDzx�8�eoI��I.c��9o�����͑|�:i+
6sNn�0�/��u��>0*��kh��TIfc���wsy+z�W���Q����}oQ[�nE��!�dԎ�4Q�#g����֤\[U�uu��V;��OQ VGGx.d*Bh��Bǝɬ�fe�mGU��iYU���f��gP�������_s]�%�2����y�oKH�e�+]u;��{)���]q���<	�#���i��\V�w��+'`�wQ�@G��>z���xA#��em|�}��V�w�==}J�fX�ޜޖTbjaK*�wK�^�Ov��;�?h5rP�������<x��8���z�~��{|����^[���fk�X�S��2�	3HC{=��S���2��ܬY�V>�R]��vJ�����d��۶�JC��J���w���N*t��p�D:}?\��mWvH�?s� ֚���'����j��� g�Zfh��5G!l���s�xh��@|푚�D6�����Vv	V�7�;��`騿>�����{���^��Ȕ�{6�:�ȣBpia{�N�o��y�H�O�R~�}\��˕�:�d�4u�Ŧm}�~���`�@��b��k�W���:þ���/��㡪�d�Պ^�荚����}�>ߍN!��{�ݨ��'nED��\\��OZ+yћ8N����7�V�F��B
�l�G�nT�6��I�J%��B�ޮ�3�C�O��zT��~���oT����y�=���qW:2�(-H�ĥHB:m؏5�`��+m���u���=gbK�CL�+ ü�5���Q��ۣ��Fn?tW����U���ŏ�'\�k�Y�>�Vv�[z����/���W�x���qǒs��;�����};��M�	�"�R{&�ch�z���<��Xd��s�R�:8ɷL�������x�n����(�p�%A
Uy fd�KHìYҍe�';��_���u�����	w���:�{���Ol��棹X�Ts���v��\C�ǟ����+��M�:�*��?v$�v֓�|Aoj�������߆8�����<��mvz��C346m��j@��T!6��~�n6t��4��QcL�{��m�&t�J�Q�ٙ��w��(�1����}���*������e��`=;;Ƶ*~�/<ܡ��,�W\jEgl�� �ы��^就��˿-��r���C�]�\u����z�Kǒ7R�-�W����{��c�M�:�կ��pd�]�v�m5ۦ��YF��"&�f%�)m��s��vM�
pYe�Gݑ�Ȉ�~�c4�2�f�q��Z+:}Ý���u!@VnO.����:�7�R��X# �����k24�ka�9}�"���xZ��kob9B�
�ܯpK�}�Õ9Œ|g����j�ݮ�<^i�Ǹ�ƻs��A5�N��y��u�ݡ	��6��r�;��7��9��\���G�yǏ� *{p�\N^<t}T��P���S��d�����Q���M��������2.����&Jݘ�9e�U��z���<)�z��Y.��*�*p���<�/�D9��׽U:��n�3���Y#r��n.<���4��QP�G-����O��3 7���z��M���z�
��uYE�S���ޗ���C'�ݹ0��(�7FqDA̻=��+6w�I�RK=^}���]¡S�ࡻ5(2�=7u���U�`�f�vf����j��o�O��kݪ9�@Fd�=¦�W�k7uaDw�#$?wJU�N7g�Rݐw����bV��7�O�ff����a��N�fn�`Wd�b��O��U�#��|]}�oA�&a��>gC5�����S���b��{�VT����1�����-�IF��L�Okq�U���Jʈ��4_)vJi-���	�����KYˋ�v�&#B-�ѓf;!��F��sz
4��%A�7ر��jA>}�n*V� �=�Ytܧ�ݤ̬��I�1h�cc��!��J:���q�sv�K��e�2�}�~�Cs-���-)���|Y0+]&k��gO�P��
������lmQvq
Y��W��ϣ�J���4{�Y9�a]��c]�����[r�U�ll&�&�����ћ���5������L�('���[�θ^�ܐ�Ql���Q[7;_vC�}���Q*a�I��p�¯y�+�S��O�V1S��^�ਦ�P��6b�y2���t8���T�:�*:�Dy��+��]��+	ǋ-�R�K&�ea��Qq,��2��Ӫ�S�˰R&0�k�G5s%Y�{W"T�$A�9\9vD|�"��i������N՛�}Ɍn�gC+�t��Ff�S6WKg�d̝L[�h"�`u9=��o`�0v���k�y�Ƿ�*Ǖ�ȎDS�o0faZ�U��|�#�lMXKX2��:�-x���H�&.R�FDJ[Zq�ѵ�1�4<�28�T8��w����@�3��Z���e��4��_Z�v5��O��'*<EW�a(���W�@�:�%��Q��Z���@���k�����ķ�v��²�v5��]�VГ���T]Wx-�}&�#<8-�Z�v�S����4�K%��u��1S�b����Uɇz�e�c�Ѥĭ9m\��b�ݬ�I�Eh9��wb[�]E�&Sif��d&�c��s��ψ)�:�g^��n��h0��kPX{���2�N�͝�U��RQ�'O7��P�k�<�R\ۨ��[�z��5a[U��{�W&GVw<��m�s�E����GVh��aؗe��y9<��5tİi1k�\^��;��d�N��l��X��-�j�c�u*�G5m�M�S�J��r��&�0nk�ٍ�r�O6V�qm�=z�:�ӷ�nt����=Z`�h�;(�����d����ʛ�!�yK��p�֕#n�2�p���uܧԈp�S��e��CQ�6�[y!n�I*��e�=�ro:�$���<CV� ��*�ݶ{��{dE9�l�Nso�]�5��F��Z ���38a1�Mq�����N�58ly*�tбL̼f^�6s����D m��ٵ��U+>0ȌQ��,��:�c�ߟ���Zֵ�MkZ�Zּk���������c_�b����DO�/�<~��3��d��#	 Cq�oo��k�kZֵ�kƵ�x�]u���g�c���*
*�+~Y3&E�Iv�U
�m,O��x믯�����5�kZ׶��ֵ��뮿?1�� O=�I�Ð�E�p��X�d�=�����H����׷����ֵ�k�Z׍kZ�]u�_�����L�Y�u�����I�pa�rTڕ ��)�/�
UV�T�
�Rf�}O�2yh[TS�QCZ)R�#*)X�j1A[B�9��E�M����w�9NTX��+X��E�z�3*�mZ�Y*��XTF1�������*�T�}s<K�V�r��%>�W��u�ȰE���PX|�/�߯o�z;�}���I�[�8�����>�d�ݬ��铙�;���86��O��k9�s3����qǑ������{�8�Β�xg�a���l�[�0E�.΀�N������� ��z��;g��۞9E�v�WG�����5�hC�x>�wևW;ٺ����/Kg�"�����s�^�H��h2!P.Y���T�i�M	l�^,��s�oX��-]�ڳ�I��9�aQ֜�ŷ�+#(�9���;i�OHw����āRo=^�|_V��fiѠd���;*��j�h�$��E��<�3���O������To�Ϫ��a
�{�sk�a��o�	��h�Ѽ��uG��-HUL^�W)�D�t�	�K1v_�
��N�U��#܈����t"���VN�z+Ζ�s9k�Qh}�y���2'ݾ����>�F���ff^�ɝ��w&��30k{���J.q��6��*�)��H���m��l��7��(�w8s��U�;<�ۚ�9V�2hT33�}�5l%��ϔ�4�s��sz^�#�$ff�%�}��#��g<5 �8�|:Q�<X���\X���*,_J.��B��{\�7c�˯,ns�X8�uޞ#��N��Z���pq����~�}����ï?���?C��!w���zs�����moO%ٷ����.�5j�y	�}^��C�������x�[��k��!�v��5Qͩt<�\̻��PطR�akh�-��2� mK��U1s=�Xr�oxΞ/��InH
��峎̀�_�Ü����ݫ����מ��;�����~���~�����7��%<��31Qr2�6��l�z�f�\�$��s��`��mw���Y�L�N�2��W˫���5����< " N��qS�����{�d5�Xݍ��g�i�<��w��$�i�ЄCU�/v͉��6`�01(�cU`jȞ/���wp/EI���C{��P��>y�T/}�N]O�}�wj2��$�V��@96�����~*�פ��w���܇I{����<�Q�n�U��qg1���0��PfN*�u�չy��}�*Wu���?k��ګ�w�����"O�lv_.���xR���m�E���QP��h�JG�E�����W�z�;�ͫ����\q�����A�~��Y���n}��s[�������ƳqV��٨f��J)�hu�Qo�K��(�w�b>�V�:�h����GU�I=ov����죃_N�V�7��\T��6��q��z�=Z�	8;?�DԆfM���(��>���z��Z�]GsN�~�=>�&���*�0�����;��+Q�Q/x"J�#�aê���[�lV�0m��tu*��+n✂/j���̨ξ�&���g���5@-z�J�"Df���I��k��p'����y�Uz�ə.��P�od{n�O�?�
t��΄�m�ޟL?qL���w���F�')y�rV��l�v}��[vS�T��w��2��yڋ��b��9�� ��GE���@�~?�Ue��M[��e����[;{5˧�n��t`	��#ǉ�D����d���y��9D�E���_����1fp�n��;���=��G�Ve�GWͳ*j�'<�u��pv����E)�w�)s�Y��MP�W9&gʔ�ȭi�#��O��#7���Sջx9����a�@gG��@8e�Q,9l+����{�HuZ�kt�7��Z��<��n&�v�u�u��{�����ע�\���+�8�r��z�`]���}pq�qq��u��߾���wwz}�n���窆`� @�w�8�JP+� �5��n(&B�5}���8ƪۂL>��3��>�H)�rށ���t𿚺�-�W������2c��2��O�0.Y��z���6�~�檾��8m,ȯk ��N��� ���Cǎo�j�p _1�sη��Un�u�gW�&&&{�˶���W�CØ{�}|���w���h�N���gk��18�c8�n#%�QH���~�˟~�xf��/�]H�T;J�1��{�n�-��3�����5r�l.q��E7�K���v�9ޕ-�yc6=_p�w>3O}o	����<P5�ݡ扜�ۦ���|]كuw����|�r�����wr-�ܮa�͸�"�����7N�!�t46_ڳ#�R��1�mQ��зُ���!�3.�G�b��kYZ(q;HI�a�C���GnΪ�}P+g�")䐬�G��Z��	]ѽλ�狸n�Q*�b��������Kr��u�֜�G�t��Z�6�63#���r�Z������~����������>~~^g^f�������o@�:��+qR2;6� =#�-�R�8�9�*�\��M���Y��cX��9�J�k�*���>��)nώ��T?o	L��T�ӆ��r<���^�1upge�N?�3�ɮ�ܢwK*�f��s3�I��Kp�v���f�ݧXu��j�9�px��S73v��כ�qL"�ym�[���$���F����8�X�o8��4���g��?��n'7�/�}>i���\d
�w�1��9���.�*FsO.���ws�*zo�����z��nԯ+�����������x�Ǵ��0l�j��A��=R�J�2r�8���L%���)�?m��HU:��<���:���gw��	4_^ӻ}���KƠ�`���T���--ܯf^�ek󰼱����]Äj��I���)����fjѩݺ�YJ��D�r��g�6t!�p��.�޽_AJ�Ĩ�A��+����'�B�Æ�Jq1��k*�O7@+���F�VE�3"}�z��[�s�w�|����8��/��z�����$E�zv�>���nǶq��0r�>S-�p��mb�:��������<���+n�T�0�BpU��r_&i��N�U���ݛ=�����~vB�VvB
�[w��t��Y�w�ʑs�2�Ky�V-��<_��;�a�
ȷ���P== %��0n�'6ռ�=���9��fi��8�e��7�z�k�[�^����3Ԣ�]T\��=թU��O�A `.ddG�������>?t�׭�뉕���j'�
<���Fx��f��8�A�p�<��܁�s<u>���w��?��6�_r�!9���I&k6�4�[�0>���Ͷ���;�#���w|�++	�{L�7�
���rU�f�w=�cdlT�sJ	�6�,��$;yz}���5�9�V�~������<�נ�:h����n�+�١��p�\���7��F�d��9ٽ>{�6��۰"��<f��3�����m�!@�I>$��$	>.e�`UA�EU"����WϾ��7�%jZf2��3:n���!�o���;˯�Զ���:��]�<��f~}zq�G�qǑ�������a?�M����չ�5���Lk,��uwov�ʗ7�����㍻��./C����6=��G���F>�XЭɍ֣�Zr��	��,e���@"�33�̫�\�|�	ݲ��
�a�'���Y�l@C/��v��~�ި����ϯμkrw��-��<v���4������S�d4�}����vza�z��.�M!V��e�n���u�=��F�ʗ'/��q� �'j�Lԙ�knE˪�㩄[����?��C$�w���}@+n�J��w�c��9�]N�٧Ͻ'3f��M��iH[qQ��5lfV�ˬ��JpF��5w����lzˌ��}�FH�"_�75Kh�3u=]��o!�s��a��5
�fn�f����r�6]F:q�7Z�NIzj���7�Z�'�Z�sz��ݝՇ��t��Ο
��B��"KMOrH�U���)#Ϩ��VpW�ch 6�P�u�4�C�/��ܘ��%�+O��R��f^�/%�}�ꇹ�(�%v���m_k׻�5�]�d{�� fU����{ޝ}��5WtԢYr��wu��@Kz�����&���f�<:��nu8����������?� ���6�f�%��67m���l�9��=����^l��{%u0�=��Vn��<?�*��V��A-�y�4���I�DO�MV*:K<5[���7�,ʡ�{��פ��ƳT�lUr&�X��
�6���B�7��Q�7�A��Ő(7_��Q�U��<+�W%���r����Y�M��9o�Ouӵ۾aA���s�u�Ou�3��e8���(�Fw�{������ۧ���#"BH�������Q���<�S���4���F]���;��35v�>AN�� ������!ϦV䳎��ro't��:wr�����R�[��ʹ����Q�t�(m�OWՏ���U,�ދ�oG�k�D�#�1���`��Y���by�0��v�~���q��RhF�z*@��Nh�#h�?���_-a��uﰼ������ke�/�'Ms��������Z�*M��v�kXͭi<��f�H{H"|���t�pJ�o
X�^.���՝�ȯ�}�ڷ��܄�]��%�G�j\ogp�}�o{ِ�5��q��<pq�s�;�W�٤��<y���3k| �<9��G�
y�ɘ���>�!�N1��w���g�=�ש�F�L���?��Oisz�y2�V�oYF���S�w���U��Pt}��>ǳ��i�fH��O���H�=~���g�R�"k���շ�TW 6֯S�"����v�--S{��'bCC�C4Da�p͌m=�S�<v;H���핻�	�pEl��a=�&䢷<ژ����tzh[鳳;=Җ��ԑ�4�{��	���\8)��S��nyo�����ؖ���Aw=�fIՀ�[����e�-�}@hZۋ��A�|�P
��1���%� �VnfG) ��'k``�9�� �;�ڶ.r�LMb;|�>�U�n�D�r�>��u�i���C{K ��4��{���T��v2m'�Q���[��-V�Mݍ�W�7�Y�C*8{��[��2��f�5�A4G��xO�9�X̡��I�vyf#�l>��Q�-�}9Oai,5ݲf�-�p����9	?!�8���8�%J��sk�(6�_�s�(T�6237�\lz��hA���O˪n/n�q�@�PY <�u�� _�=W��͏m���F�=�t�܈��NQ����M<�<��"}y�7��b��ku�1,��W���'���e{L�q-[�t���M	��U����x�c�l$�8]�;-��n��WZ�m����w{�oG���ǜ�v�=�΅�홇z�ì��V(��=�E��L4��W��U%�`O�k=
�G��O�@���=�7�wz��#fw��~��K1���y�s�w/�C��zk��H#�6���,�ا�l�w�<��G�׈�Į`Ϡ6h��Vu��#������*��:Զ�׸2��Ln�85������P���Ev�N�Ϗs��Qӎ���\�3�6���rp�[2��^���Ý���2�R��|�i@?��c�km@�f��LT�Q��T�x�Kc�)gw$�|otX��7v�E�8뽥:a�M1u�n1�}b��*����w]�A���I���օ{{c�6pڬ:��{:�,#�E��c��$�7��e�䳕�@�hd%�:��,Kk���0����Ѭ\ˣҡ�$�AS1�pjM�nVT-�3�{����;l����2������T;Ml<�������0ަ������tA�����F:�Z�:/5b�'T�q�cח���s
�Aח+T���/N����wA�݋gO:��9Mͩx �`��y���n5���ؚ������N���)A�1��"�/-�>�j����N�-�]%k�5�n�g�%m�N&î�ִ����Q���o��f;pκ�|��U��q���f+���R"���M�<�;f-V�Sft+{U�->Q��]���KM�{�R��h��g���<ob��]bn�w)�I+�o�g����+Zu�pF+ �w0���>�ֲ���{��.�t��ʱ���q��]���dt�F㳴!�`�2�ݨ��n��37[�܉L��+y7-�,_��]:1�=�Q�ّfk���Ę9���_P�����M�r��݄��Ym��.���C���E�k)��ZAM]\�}��]�@��u���1�q����51��V�Pϐ���:Q�*�6�5%���(��4]��[�H��9ס�|������Ԓ�05�٣�W������L��n���m[�4d�q2e_{�ⵃrK�S�o��ww�5���C����W.ܚv�m%��3x�q�����cr�i��D�¹���-#K��5��
d��>X�p�uaB�d�t�[d�mfx�l��L�p�ǜq1�uh=�a~1��@W��5���#7��^��+3�uH�S�e�1�9f�6���*C�	��(j�c:�;]&��fi��]fj�t��rk��:�L��]���M��쳄S�c�Z�w�(����MݛZ��vڅ���^������[Ʈ�k�g�5c����&grk��j�LZ7�1���JktK[jf�ޕ-�Ф�N�z-Z�[]�i�Wb��q�WTG;S�g5�a>:U��Rȴ��:�ٻ[���=�4h�N���/0ծ7y�Ϊ�g ��0��{JK��.��Yy�vd͝Z�=tλ=���~�&��4<�u]��p�W�>��;y|SA�F�)(ı��Ǽ��s��To�����w�n)�V�۾����A�哿�߉�|G�$B�����=�L���OIQm��I�;��1�:�����ֱ�kZֽ��xֵ�u�]u���{��;�3�io�d��(�����b�,b=H��e��~����s_^�___�ֵ�k^�ּkZֺ뮺����>{��8M�s��3	��Q
ز�+o\�bҍk��'���׷����5�kZ־5�5�k]u�]k��y�y�@�Z��a��V0P�k�yv�ifrg3!�q��Z��ֱ�kZֵ�q�kZ뮺�_�����L��)Ii{��m��Ũ���co�ة�Tb�J�R��KjH;��[
sa�*��^q�2-nث�kO;tzа�)u�;/��9�j]�J���E�-�V��.2�dD+_Nג��o7�T=<�h�Q�2�z蹵���g�^�Kl�-�R��݌�Ѣ|�u���h[g��婩E�<�_�f���D��۳�u����l�1�jS����[S9���v���Vʊ<�n���cm�ެo\ܻ�vn���N�ΛrSe\ncM9m�DDR9��8!�� �N�����U�ݢ��tG6F�S��v�-�h�ݮ��5�N��Mٗ���TZ��b�G������^��V�K��y��v����)��^)�r7��a[rsT뵸q�lwV���ʙ�v������;�ר��n�Wk�][zS���W;N���ln;l^/;����sr��6�km��{�	]�W\�ƁFIP��h$$(���څ/���KU���m����3���W�{����ku�7k�ս��σ�\@��qq�I$F}�i=W�mC�>܆�ۊ:�C-;��Z<����%��e>�x��r��Om��o�5l��;��`,�\mT�䇍�4	���3���SQ�O�l��l�;���h�Gq��y�
�{��u��nӏس���|�꾟)k��܆�2A�ouf����)	�u�]���S����w����ѱ(t]n�g}�A��:��&���o�[9O��7r�����,�b�ř�\�;g���zy��w�Ѽ�V�0Z�����M�-g�D���:��n�u8$[�-�	�s345]�*_�v�U<ǰ�s}�N�n5�:6�dn�A�
�
���'�\�6��U���$�{��t����K�q6�/����O��C?���c��{���}X ���V�:7n�g�1S:�g�H�k�1���d�Ef��������Z�]TJ},[.b�{uP�"�yƆf̮��U�Jb�q|R�V-�����<?d��9%��n��9y�m���/�u���MeǦٳ�9�SN�h�c����"Itz*�(o�1�0nt�B�r�Bv[�yM�f����vf���n�lK��>�&to�����,�3�������©��������x|�k:{����|�3�0?��%##��"��hb��g������ۙ�7+P���u��0���g�w1h1璘At��T�u�8�n������fo����ǗU7��K������.G�74��l���`��(�� c�����c�>k�ˮ
۰�i��=&wr���9��*��<rr;6��s���y��=4��.��x�����G�����t�ٳE������f��n��~�:���ҁo�zO??����P���#"�1�{8g��w�ϻ뿹������+4����aytaC��VNoY��k�W�8o���S����-v��<�#j��"}�]��䪽��y���x�/DY�:�J�1|��	���o`c��,9#���u`lL�П��[�!]���09o\����K���5�p�a����L�w4�Ƈr��_ҰfE�*��f�ت�o ���dvo��2�P�{dخ9;rVh��vNL����������u�p���u�ӭ@�0L��j�.0�X�#�r8�#��FD�?o^��U�Xi���.��Ձ}�́o�x����:��'��p�E�F�)��C�׮�ӧ@�����zo+�^����������ˌ[CO��'WHj�Ѽ�g1A&���D@�����>����p�ztI*٥�eI�|ȗ�{Z�Od��=]7�/c[�`y�4#�D�L�h2+'�L2�\�6f��3�y�/���u&�v\TK��� -�w@wQ��l�3���&]4.����(X	����6"�N��U4�'��$H���2�a�L�:C��8o7�1
S��e� �R�������M\O��8��s/Ֆk7��wGNy~�W�,ꓲ�$����Z��(i�Q
ǅZ=;�kg]�;��yP��@��g�y=�M����t�)�r��a���ݧ}s������������dY����6ym���m3�e�AN=����r�c&'�.��X`���0���KȲ9/x�ZoY�f�3��9�p]�}���o��Mjjb<�T�py'X��H�)�,��iN�ٞ��P�<c�c�q�G�;۶��՟4�&7v�M������2.T��q�g�yi�ܷ���ݐ��4�����q���ڟ���gy3����eޜә�N�Ow���}L�� ӕ9>�{Xg�@�0���aӄ�s�'f�`���I;-�ĳ�Ќ�&Bڇis�K�߱��E�~��l���ΚXz},������_옒��rm>���2�X�0��<us�-����g-�fy):FR��L�gl��`���wB*�g�=�e��բ�a�k �Y��_'�����ѵ�5ۻǼ��j���w�Q�z��=C0&PN�\������6�Œ��d�R�������eW�[�n/e��)�Q��s��}�
q
�,:����f��D�f�Mj�Uߖ��\�Ίǅ��Oѽ�;i��c�,�m�rMt��r�G�޳J�q�ң�����y�2�ԃ��߭qm�v.��Hgo��H$+�*��:�������}�T���m��TF��	k�د�tҕ����w�y|�wM��w�/���q��8��r3��«��;���q��35��ҵ�.�k/^��c.I��T�&��ҍ�ܘ�k>.K����B�Q4ݟ�@��T�Z��읽�|�lER��4�`eL��	�a._�}9!��+�7��VEh
����	o-��v}Sx9ƾ�\�YZ�Y׎�xt�{�<���*�c�g�\����ϕ���J�'
�/�nk���?H���J��Gb�8�{���NT�*b��o�9H6�HZt� `ng�~�|]�<���-�^e��H�S�g��m�o^��r[Z��@�S �1��Y����t��7��Lŭ2J������.�	nʾ�7�u6�>4z3i���-���wY�Gf_:�1ɟb���k%3����r��Q����V���OB|` ��6�y�����/n߰�������gc��RH�뾥����k½^F�x����?�.�ɽt&�\��In������~1#�C:���g>�VOt�N��7�"�]��[��5F1�t�����]؆�E�vX�6�=�(����yF����w˨��~m�Dh{>��ů:'u����C�a�N9�6�^�r��Pv7gQ��:wc��y�z�T��+�`�b�C��|}��~�CϿ��_�����JA� �Q�`d����Q���3E@�':��s#m �}9ޙQ}^!����]>������ɫ������	{��5M(@�],���bE��zF|ʿ��FYcwڸ7�[���Dvz����M�_�]E�G�Y920�x��7���yf�CÔ02UP�᛭��dv�X�\�͠�m7�á�^4q�lP�d-�.w��i�R9���0�p�kZ'j�Cd��[n<;3���K٫�Gw?��ύI�~*�W.�_���N���[����ڵ�V�.=��<� H/����荎��H]�fO�60+�m���FA�������OA��ghOi��ͦ�&��WP ������u����9'5c`�dsl��E(�={4{�,���s��~�>*X�v5�n����}K	��C)&*)fƲq�w\��Wv������nK��S�� �� g^��Ӧ��pY����f���S	=L�c�x�owy�5Բ�l�,؜�n���w��w��lX���� ��~yzg���n�����q�U������0��[�g;���~����;�7t��^��t��#̯ ���<ػ�������z��㞣<7:eN9ŅO���
���ç�>We�foe�e��oT�\NYH�T06|�v�)�i�dk�O���;Ƌ9��;�E�q)E���F@$�5��6��;,�	48�3�M�4΋ޚ�>�z�qK�O���!��hP��p'(��=�q���#��$lX�xՊ�MUMg�r�����[���Hk��Ƹ�;Z�-ۥ6�z�}#���&=P�K��R��j�+��h��ZV*f���"�檼D�R��;6��40W*�	���{��
�r˦����+���+R���fWjT!w7��ـ�&��Y�<�Z�>2�3)�x=N@��W�!�`YH���9�Eö��m�R�ض��`����
��ŏ^��W�f��m�F����j��������-k\�)S��kڡ.�-X�j�F���|;�I��������b�w痯���߯�s���o_��it��1����ړ^<�̶�T��[����1}��x�KWLG��EN9+<|J��0�Smj�(���g�˂�VDc�<Dg���w+����&���9ް��?f�-�F���<WSl�Tޣ��0Ӟ�@f��(4�C����S��p����<?��ܲqga�XҢvB��#�q�_�1�uu�+�Z\�GH�ݍ��҉�������4)d�f�z��c�چ4-��m�γeH����w�=�O6�u�o]�����
ff�8�[��;ؘ��v��V����y�w��������D��{�@U���ԔN5s��xC *������i���6�'̕��=��#�M{��5Z�36�#vXX*��e�mz��� <u���o�C���+şTM�w/�%Q;�V~��i�m�E�әݏ�zD�TO���Tٕvntvqt�n��R<��H�$ �e��f�U]`�utilv�㰗.g:7�#�nw��י���gFu�/�w&������f�w�9�y�FI2?:��G1�<}����5����\��a��Wv�Nnm�\-���q�f3C_"Mv��w��8\�=7$�r���Q�뱃1
ޏZ�q�l��^ӯ��a��,�:��o��]g��C�h��S��Ҽa֛5�g��x���Ad�{�gw)�'� ��C�!
�5��>K��|�<�^{uO���f���F���1�iV��L8�l�:IA�#gՙW�<�/N�[w54��nF!�;7U]8O�����"��E'�~��b����y�(��:D.xɴ��s�'I�Y@/U1��x㊹9�0b�*Ӂ}��[͂��Ct�,t�f�335�8@�spө�p��7�6��`����8�]�&��L�j�h�*;����@�K��8���K��hp�b3��9���jz��n�u7o��ή�/��~�;.�v3O��t��v�窊���w�Z}|^�Lw*2(�O��(�e= Bo3���-�R�����V_�er� �uÍ�u�G��CxH[')�%�\��(��'O
�ߘ�]����f�ʳ�&�#L'ْ9Ӗ3��U�u��ӛ$�ۙ���E��_n��-�7گ�������<�o|�{h�ݥ�O�}��x�z��}����5���[e'w��]���7����p曁� ���˭�9���Ӆ�c���*�}������ϊy�/y�C!�<���:�T��3�"u�75P(���_@��gz���P�6�=ȅl��3��f�Pf�k2�5e��g�{T�F�,o@$m�4.�!��:oRd/:�b�:n� �Ƅw�|��E��dCaq�y��}�^Z�n�y�nQ�Km�;��/MsLwpz3��{܆��яz!jKT�L2�~��8�s��E[�F8�0���|�n�b��@oSxu{J�XA˿u�K��{k�R(A���΋�d���ɹ"к��6xz����2�;OsLクs���m���t%�jznvf'-R���|-������U���4#�'�G��EZG:�{+�s]ym�o�*e�Kc8���ek�]eGL&��6�����֮�Md��C=N�����nH�v���W ��ŧ�����Э�AfO����F��źA���f
V�+�V�q �&I}��%�F�N�8$����{s=��X�v"�;��D:�ݩ�f>Ɨ'���fWz�p��	�w��
��oN<.:�N�m�M�f�/I�+��2���t�݌j��̽j��I&�U�Q/���K�����j���W-sl,�Fhn��`��S�]c�B`<lJ}D"�:�ںJpɤ7�<4���!�"�k*�����]Eï���9af^T�I0�۹�pJЈo=|;���A�0��=���O@�8�<�`��eN��I���i���5s*�co��\��s9�&��X���撑�$ʽ��oU(gBOB�]a�Ddr�\Med����v;
�*s�a��[DU�΋;K�qU�0ru�]=�m�fN͆�1��sO�x{j�7��ǏV�meA.�-�Km�+r��a��\xu�}A�?t�4�+m3g�.�(I�t��s*m*�^TWd:�L��M�M�pR!���J�ͷlWe#W�*Ԇ�]TEAp���A
O�Q�%������#��
#��n�T��Į��R���Pe k�v�9�Xެ9��o5)���F��S,G:���j"�gs?���g��g��ןk���l�66�;IT��q�I�J�y�ɡH9���Q���Շi=�}�#��͂��A�P֠���;6�uq����D�͹SkpLX-!��TV���^+����zo';Zy#H�t��.�QHÃ3�� g��칾���B53wk������b%.�/���Ь��N&�����鬎[n{���ո��%ǗEKzwe[���� �篒�<�Y�s`��{J�>�y�}���h�0��;�ۛ��i�8���$��7�Ц�La��ecV] ��MFmvH/P��6�'κ���ԦI��R��C�y�]E���"��˔pX�!�w0��4�t��"�Ii^q��A�c��#9Eܭ,�C��Ў��m!c���M�48ҁ�Npnz��F.Zvpi�1��lYp�y4&��s�X~�hZVm���P�D�s��i}�p���SNwwqm�w�N��ol�tO=��[�y��'�ڋĴqg�ʯ�6���"���XZ�ֶ2ΞO���kF��kZ�ƵƵ�k�������ȹ'��iÏ ��KZ�񡒰[R��VYg�־�4kZֵ�|k\kZֺ뮺���,�=�Q�s2}	��!��������C �GդQHΧ�N:���_���5�kZ־5�5�k]u�]k��{$a�9��s�%
��tԻJ����7�D樞[���smX>���'K4��|}~~~hֵ�kZ�ֱ�kZ�N�>�����lV���:�S?)Ԩ"�\�eAe�/��V�����Jؖ��{*M-�}~�,��vJ݌�oƆ�E��Zʔ&���τ.�eeJ�-���zlڨ,�TAI��>mu�eV�m���-�����_l���ߡL��Һ�*���O6�)Ʌu���=��c#m-�AE�Z��Iǚ+��V�6�U�mw�(��S%h��Pͩj[e�� |Jx��e~��}��O��E��߲����m����)�Lw9H̝��H-�����S����D�a~��F`�"Bu�������s&�9�y'9�����5�����>� �? U���U<E�e=�*�� ��O���� 6�JDF��|x��i���v��;�n�b�=[����v�H[ϲ��j�֧x�,�x�oͩ����2�s)�óJ3s�N���V{��d��O]}[�U�_������v.^rHý�=2�jt�F�ͦ�o\>@/�"m�h��[��N̞�,�<oP���	Q�vv�o��ň�z�{���m���B�͝�`���0���Z�h��y����V�����Iҕ�
08�g�+����L�z�f��M�@9������Lk��-�^22	s���7��zY�"�/w���Dt�=��=�.+��fmYqRԎq���e��ѪN[t��|���7v���2�^M�����M=���.���k�!ò9��ew�b���W)4�c-sQ�I���ݯ�RO��-vrn��뗹}��RP�.��9^�7��|Č�1���wܿ}ߟw���w�`!�Z�X�۪��`�fV�a��Sv����;gh�Gk6���ځo!ɢcH��V��wBj�4V�qp��1f(US<�g8B��� m_�'}��p>���k���g�,&��<�ӫQ��٢(�+ޡ���Y��²'���<]3v�c��׵y'y�+%]�i�[�X{�-*C�UO>��츍���ϼ�Q�g������Ǡ�g�3ʞ�`+*N��I%t��}3u��'�P�����I�?N矁���"^�wDI�@It�n��`ָy�\��$�;{��Y�:<l�-��܃�y��V
�+ ǀ�=+.���fa���#� �z�����޿^�c 1v_���Oq��:zC�b�[w���ΫJBS�՛�����q�ܼ��<"6�2�f
��`DlH"bY��bm_��̛�i���n��r�]��!(ę~�|4(��W��#�+�bŗ�dz�*�������А�83G=���0��ں��4�Y[�E�J�eg�`���ѝ��)߹�i<ɟ���1��o�e�k;Ek�%���5{�u�C��S������o�eb���=�3�)�+��'P�l�ӰhړE��y{&D8i8e�k#��ӳ��M����Cs$ЃM����0z�j���㕚\]��!o������������c�������%,q=[����@��fdE�oD�LB�{{��n��\
�8���K��;�j͕rt���P��g��[���(x�U�Sbޥ���W륝��i7:�d���[�j9���
�1q��-\�,�}F����;أ�)��r�"�OuI�SC*���؂��1�~�DM�ϫ�u�Ył���X:�ֿMi�:x����`L��q��4�;JE��Գ�lǟ���U������Ba�zdu��L8��U�@S[JIW#S�̊}l�"�Cl��'������y��~��3�ۊ��P�́V��qZ���k�#i��b�9�[²�F�(@4q�\���uVh��z���یɧDv��H�UNHr.��xEEOʧLSo�WP�N�e�e��!|/[�
!-,4'�5���+���5�^)��}GnN�o
��̈́_N����Nus}yC�E�C�k�沂�z��~#���y��oa��%,GJ��Tyw"����q��\S��9�8�U�>��s�Hj������).��y��zf�~��Jt���63��݄�_q�������q�kƽ��>��=�^��b���l��7�v�� ;:P�]?��3J�N������V댊1��Uyw$NW ����z&٣�2��-fٕN:=ȵ�_�GG��9�}�"��ݜoft�z�6�8����YVfg�U]�`����_�$Y�>~�j�x�OhPd��qT��YfO���������1�0mi��#���ǯ7<���AjȊv�7b�+4�7����!���i�M�R\3����uu]���{�4��;	?����Q�Ř43������O3d��k��7��=���߷�:������5�0�
�}^ �"��r+�X?�}��%ET�JOE���7��w��$W���|pf���ɡ=L*\yZ��$�}��y�<�]�.�廻�8p\���M�u"�H[������Ϭz��Y?`�[ݖ;��r�)���;��u���w��9���<c#�$󾽼�)���?�d@�]��?=̺�z#�3��U�X��\)�7ZT��mV��[>��(j���&�Y�9sw+���z����������y~�ä�����&���*߶�ۘ�u��dwO��������t_�U⧹�q�W��
=��6�m�@xl7܎�`�w��|�z�VϪ�)�����j���Z^�}`]Y�v���f�Wj[��>���a�q�� _<��K�kK]�56��Mу���\���zT�u��
���'����c��[�e�ۭ���e�Ia�͐މ�-��*�����秬�.WI�^�^aYn�O�Yy6�r�Re/�}����m����Ow��s����DK�U;��㷷���]�ot{ʲ6Y�ʽy�R!wy)3��Z�<�왝��qr�&_X��E;���rJ�]��|�j�#��x����Ǹ��:\x�iJ���ki��l�k���Hsi9]K�I���!;�o�+9k����K_���{���{zTa�H�絁�`��>���~��x���s��޽������xmv�̞�+���<b�y�ȾÄ�<���5�Vs��v����Lv�E?c���3�V��g��[�Η����ѷW~�#%��\�;�=\��F��!V^�y�L��w��5��ۗMd������Avy٪���G�s|�Od�u9���b�¹d����߬{�Gf2�dʽ�Ż���y��r<d�h�� �f�Mu�q�x�<C6a��E��;�351!+��hx\�n�����^�^� �p���
[�лƝ���Ս�"�3 R���"��O8���Þ�3Obi����lu�l��F��(�u�8����=Z���A�u��V��Dvl����+���w���7� e��r!���)�I�c�5��������9�&~���Xc+/�\�Iu��v����.��b)}m�ǗUG.�/�]�s��:� 4���,`�<���S:[�k��Ƌ�'(���P��E�k��Wax�q���Uș��=q�({e�?��޾�������Y�}�0ګT���,'��s��1M���5��8,ՙ��n�&�y"ݺo��`F�>���������Mx��\�%�����tW������/�G��T՛�6����s�zK�Z��ڶQ����epΟp�r��W���Z�c)���Đ;t��I��w���p����������Pm�B���cǀ�V 36������,��e��	�|�u����5`w�ܿ��sxW4a��誔��d
����=P鏵��{���J�r�L�����s:'�"_/&�+7�yz��^g�ӣ�_x�3��.�������-��Stc4ٮ�27D�	���#>}�"/̀�o�6���~p�-4��g��ƈ�Y�7�Zr埁|c�J�_)�k��N:�i�Y�����/WV.n�ˆf��{ ��+<�5*E�>\��j/�V��Ɯ#&�6U�o)�׷#(�Xz��K���N���������S�t�9o�(��r\n�;e�r05�y�lh�6���=긵�g^�,��F��2�hWb���9ո;a���,���H�o�Bo�E4���F[��5��L���qtν���}�T<<<<<*�ֳ����a�هhC�L��8�r#L�ґyj}t�̳:R��=sSv���~��>գ&�@T�q�p�Nj�U������}{{��ڎ�}I�%�a�M?H��8�b��S-���W��HiҐ@~���7/�~=��$����.A��r#���4W�x�v��gfSg9�/# ,�H�u���%Lz�+���+���+q�!�Y���^�񒁼�z=�ӦCT�]�XO���g�~��g�7/skg۔!���L�`�D?���j�F=V�ΰ^��H��}�gu��LbBb���W�7���~�x&�v�:�3ܸ%~���[�<�ȑ;RԪ��{n�d鳲�:��V����H�L�ݼ����>j��q����=���:�F��ndi�'{��o����3�r�O��q���IIr>˹����}��_+Bz`���z�d�[�U}LE��]_g}W�{�M��<&�_o&z�,l\��)�� �J��ʂ��(��p�����]�z�>�U��JT��ۚY#��}Q{-�l�ᝆ��gc|zrZ���ea������C������w�i���hF�'I�&��c�c��~���>�r�rOޏN&v��w���Q�����7����1�n0n2	��c`�.�X>9%��]tc=�H�7����U���Z1�Ȝ�^�06Mߥ�V�sꎉ=u9��*bi��+ ��w�s;||5��˲A�"�\߻��r�B��14���� �F�p�\�4
��~J/{9ʩa�Vfvح�Ƶ-۸�9-��t��$�q�u�h^?)�{�];9s+o��2�(��'���S:�E���|�l���ޭ��yrOeY�L%c���d?b5�A�����&��a8�U��촎ѤXwp��r�D�����GB=낲1�1�q�\���r���]{z|�6���;(�;�n��DRIC�]����##�G�5���m2��Sљ�Q1���W-��b*q� Q�t7�1��8c�"I�F ['�3�����b�,�vM��3wT0��G�q��.=�����Q.Wo��d4�j�r���]��bÙz�����O��0#c���=��_~��33J��U����;�~�2�QMS�x�fN�J���Osq��K��9O��1��Z4eg8�T�����1]�o<'l�`����;�9]"ܽk���|�}�Xǒ[�^�|�HY�ƺd��G�y����qhh�OLLW,����gP}�o|˷ę>�͒�W���_��Wc@�����t[-�J$��c��u��it�%���^�e#�A6���&/���++3畭�������U�#�����/��'�<����~�,3ƹ6�4n���n3U�(&j<.Y��/g��+�f�R��Y���gȵ�wwo�
,���hu�t���G�]�=��S"���D��U���l��a��jӐB��l�j��	��S�<}z����w������G��
��@PS�/����qEU?�AE��1�	!!C�xz�!H�@D1�a*����F	bHb,R0 �"� X�H�F1P�#H���1��P�H�!#B�E��$�H� ŋ2@����FHD� ! 1H�	��!Ȩ��D$`�D$`���2 �X�HA���A��dB ����FFA�$�	�@B��b��$dB ���"��$ 0d"@b	�$��*��F�$
�D$b��� ��@B
"� �c@B0��
d(@b!��(�� @b���X"�@b!��*�B (@`��$
�@b��� ��@B"
@b!�$@`���"�w�cκp��B H 0��B HA 1P����A 0��BH@ 0D�� ��T 0@��BH 0��HU����#D! �H 0@��B�� HD 0D��B 1��V 0P��A 1V HP !D 0P�� 0��B !HP 0��R 0��HT !H�H@z�P`T�1PR �AH E�1R �DHLb���0���@ E �0D �P@ E �0 �@@3 � �RQ A 2H1��0�0D�1P����	���d�� �P��� HHH`1P�0�0D���  �1T�1�D 0 0T�1�1P�	��$H�B)#	�$P�F���������`� `�A��	(0a"����*d�b�$�� ��B(�b��FA�������XȄȄA###cO����t���s��P�TD�H@�w��?����?����翎?������l������?�?��?W�����_����W� W���C�?�����*" �z�@U���c�P�@b�S��|?����O�b� ��/�����=8�s�w�bx���	��O����L$���UA�@X�EB"�$"! D�$P"	H�@"�XE�$@"	@�� )��E"��@"��Q�$b!�D��P"!���`	(E*"	`	�HAX�F* ��� 	�$�$ ��$ 	 !�$�	
�$(, �"(@��@�� �"$��,�(Ȃ ,����I UG"�B A � #�� �D��b!�D��b!�$b! 	� D�� "��$B
b!��Ab!"� 	 �`��$�� �$H�EH@X@B �V"�b!"u��B�?��~ޟ�D$U@@@Q�~������Fo��������S��\�`���o��������D���}�?�����mM?�����
��'����M=����� 
���C�>�����GAD{��(�������?ژ����x=������hg��������
����T?��wP]<?�?�����:������W�?���>�������?�Z{�'�����?ڀ *�px_�=C��1w��)�� �����?����@���<���^��#���)��4���ǫ�Ŀ/�D�u?�����} � �!�����_��C�����d�Md巢��af�A@��̟\��|��;j��A5��@�%*R�V�j��h���)����A	*��HR���J%H�SlDJT&�QV�*�TkF �Z�F�mkm�IZh�V�4��[b��1��U�#ZœM4�l���*��[Zm���&lKYh�(��(�UYh�-�&��,�j�;�6U-���l��6m�JX�*[i�4a�Ҧ�m+m�Y�[f&V�Z��RX��K-A��Sc[SfZ+T�1�E���m��)����m��Fll[\   \O��6�M�m4P���%ҶƫV�uV8l�6�s+�(Uh�mZ�+U�7u������.��@J����&B�.�UR�kd�Zfʹ�-�EjMeh�Y<   ,���v7clm�a��y��B��B���u�ti�Ҧ�C)T-�l��u�m��ki�li�R��Z��v�i6�j���Q�5��VՌ��wm9N���U����ږڍ6ii��V�   g��Qa^ۥEm�2T��m���h�%��ͭ������Z��M��UUEK��-8���QUmv8�IEh]ӻ6��٤�͵Z)�h��  �J=wk�]�U]����Z�EV��Ӯ�Un뛦؉m�������Tt�f��Xi�i��j�M����UEJӶ6�5V�R�f�L�ٶ�5�   ���U�UU���Z�	[��5`\� �r�b�:E���R�EZ�۵!Y���:u���������m�T�U�V��Qmjh�����mm+�  u�j� �u�  �q�  s�� P�,h�[�8 4��� 	��  7n  1� 4&.��tjl͍�������  gx�-�75�� 7� .;\  ���V:�u@gN� �f� ���t 4s�Y�֦U�M���4�  �x+��]�r� ��-� �Vp �isn 
7j�@ ��  wr� �wum�� ,�  h;�ULS[kmDҵ�6жZ�  �x  =��  �,�  sv�  ��@5@3� � �]�  �ժ�@ ��K� �Z�kk�Dȵ@��  �� �  n6� 
���(�v� �`�A��  8s  'u\ @w� :���&4�J@  OdbJJT �����h4  O��SSM  "���b�U=!�d��)IUI� 5'�$�V�Fȣ����=�f�Ҳ9�EÇ���^ႚ2�Oo:����>Ͼ޽����{lcm��� m���m�����6����66��� � m�����_C��HU��tm��� B�lR;t�dR�U�a�2\�^\? D̙��R������R� ����d���`ők��k�����D�v�dǧMj��Lp:R�95���[�.�kn�˃D�[�Z��Be�th,�Hc�q�
��̇2�seӫ��Ĥ�>�J �P/� !��P��<���x�\�w`�%[!9t�a}��=َ�lf�tK�W�v�G)B�t�TF6���VL�<�V����Jۡ$��,;�van��B�C�K�R���ݫ���5^QT%ff�ՑLF��q�3oN��9
�d�%��-��M4��d��w���j:/u1:�8�;K6����ECi}�N�л���(ڒ\F�_{'tU�e�n�uc\%���އ���Z^�f�̣):�hhq�]��!���0Y�����nR���L�]b���hDő��:����7l�e�r�ZYx��.��r��"�ff[u���K��H[`.L
T����E��Ԃ��V�W�H�ђ�b��{��7���J����kD=˳���J�d{�5[[ut�w�J	��ab]n�.�����2B�S���2�E��,�3T�29Yb㡢�(D��ٗ��(�i���=����V��A��V	R�;�hh�eE�wl4��F���:@��vވ@Q�A�����G7�f5�l�{#R��Y-�8B+R�&��X÷
$k�h���z塡�^�t��ݸjeh
�2m��������ku��l�	��Ij^[R(�ϭ1mn�,5x0����&�ͫ���#k(�94���	�be$�H�����@i����D�D:.Dk@���2JY��V�J:�GR:2�îi�B��(we��5���R�p�㧤R�vRv����Ў:͠�;�:j^�hx,��X���U�ܡ��QMiKGMFj�	6��ͻ`mD����E���M�m6���{2D��jW�櫧���Z*���Գ�&j�[��
��6�/jÚ2�l�m��,�@��r��s*\ ��31L2Yi��R0*�]	�9Z�ZA����QjY��hV�{oL��L"g��6=�䭣�j�Z��/&1mӪ���@᥈7��h�z���F	��ZS�i}*Ë-䡀O��o*a�3DL�!�� `Pi��nP1D�EK�ّm��(���Jݢ(��ch�H�֭-�UQ���%)��:�n��Lqk�h����A�
cg�+�c�y�qٷ	_KR��%_n�Q�&-��I&�-��,r�+%h`w"(iz#�j�]؈�`�x˻��Yf��ܡV��X*m"a@�i@(�"��8��m�,ǺRJ↰#r����-d� j*���y&��iM�gA��7J�2/�%;�{�5,TX�4���(���Ԃ3��nc��v�vjm���5+�m٘��R֧VK��;��mݜ-��q
�ḳ���'>-�x��ejy�Lx�bT�!�Da��kU��
8Pr�j��SrͫQ=Gn�ZU�F�J��9��8�8�Z�qmЂd��I�n��:z2��,5�Ҏ�i�e����Xz���^h�q�u�14���|�%d��Y @�P�	������;�y�P�2.ĺN*G]n�Ȁ�V�f[�幆SmDF�����MlyW��aT��C����=;���t�Hd�[��s/e��I�q�H�mY�L��P`g%��Cr�; �bIY���Yj�;��t�f�.1hӅ��̒I����5g����ʔ���JR�Ң�@����tŐV�,l�*� �:_#�)��g��z��x!�6�>�eѻ��<!LB���{D��Jw�o�o����c{&�;}3U&�Bh��4�Y�(����P[7�m;[XM�AL��㒈��C�2��%"� ַ㲝]�j����H[dB#��(J�KbL��,���=��]jrP�^��y/3��F��Z���[�H:(BU�%"����O�[�xoj�<YE�WM�f�DL��-��ɦ�(��Spk��CA�.+�m+��ڶ2�7���t` ��R0��:T�6l�P�yCc�f�'r�T9�r�X��m��7R�leQ�n'����ʸ#��ո*=��1-�Kh`�p�^��1����l���a�z�K7R�Q9I�ux��,/Y��6v�MT�湴Ӑ}��B�T2F�;[�1V*�t�0n*ـ���E����*��k�C30�X`�U��<T����yi�SuJ$���:�ɌY��6��c2���oD��C,�xDckV�������Y�8��pb��/U��3n�D(#r���*fdċa�t��u�)˧��M	����B#n��Ӭ��AT�8�2�2�`�+�ʲI��-��ЫƖ�EX��Gp��a*�Ǵa�:�z;��!��[��yvw孅E�Э\ڑ!q�6܎]���|Ш��r�eBZ�ᣦ~�	9zsFb���vJ�9��IA���W� ��A*�k��2���5��e巳��ܩ�o[�[A��Db��m����)��ۼz�v�����U�)B3/iB�s��4ssv�Fc��Ӌ���j��k��9L<J�8�Q�w1�2��Y6��lz�/w�Q���(�G�/I�<B�mPZ�F�j8��P�.�nU_�,:7G��� �l�*��oi��b�*b�(��CF2ʺ�rehKDN��.��d���%4L��"ܽ�����^���i�un�V�J�C�{!�y+:�R�L�f�H.�4��q�������K-�v�ǗM5z��Ԧ�(��S�F i�����hʼq�s.���2�kj��c/d!�T�-F^4.�J	[Kv}gf=�tTRff�0�K6�a%�:�H��*5����o s�7A���e�.ˊ�c^i��	��F*KUޖ��ڙ�2,[
���76����1wl;�L�2�C���t�� ��k
�cg-"0��
ٌ��òZ���/0�j�����o|h�!��b@d�.�`$���zFL!d��f����ft��0�w1v$���B򤤩y���㻅�81�z��X1ro�4e,
L����$�t�5	�j@�X�Ut��9t�2��$��f'6�dֳfZ���h�y�1��H��F�a\�2F2��ʽ%�SF�0dB�إ�طO@ר����Uz�������.��X�WykY'$�Ytk2�9�	jfmLt�	r���L���Be;��%[h�`i���Om��e�*��QA�&���� ��ؒ��n�0�Yf�z�b[�d��]f�q\!���ڻ�X���j�4m�1O��c�(B�r�3�2��[d]<.]<	<U�d��X7e�(���K�q�����u�lY�-�jQ��x��� i�p�v6�:zEkWVM��X�vakV� ��%�)��vdX�j:ǯb������	�(�y��2�H�VI0���]^�U0�C���j�r��u09+m�
�+j�;�]Z�DRx��J����+���Ŭ�Q]1s.�&�ph(��g�b,��Q7Ub��7�2�ݑ!ᴵѬ�����JGx��gK�E�t�E��-�D� ^b82��f�<�
XE�[+o3q͗�V�8j�[-���,��	��9*�HU��i�2 7o��N����{B�4��)��4В��
��z"�Dն��JǏ-ܭ��l�E�-BT����ZQ��llw�		��G\1���Qμ*��1JpL�L��4|b
�ҩ1j
�oe
dw'���W�*h��S--*�v/q���*]�kn�:6���5�N2o.�
�d���r����ի���2f�'.��.�,ݩ�1��T�_�k͟[ui`��\H7tVM�CBt���`f�����&�`�_�/5D/3 �ڔ���D=�[nPd�u�R��m���LѦ����#����Fzq#ݺ��Oe�udg"$�X���I�U�ֲ"ed7����ht'���`������̉9��	��dob�M�`�?�D`��.������Ս8m�a�-��S;S�Z5�2���a�I���R	E��QUy3��Qo]:��[��F�;�G���X�r
�o���{�&ɏ7b��x��i�쁆���`��K� �C\Yy��TplOJIh�c�#���"��2��Nd�b�r����x�I��ٙz=@Y�4,�u�8�f�<��$'^ݛΛL����w�R;v��Y)Gl7:�d2d���Uۧ&XLT"�������ѲW���B�V�B嵐���>��o
�
��Ì��EP�$�(�f¹�KЂ֕��:~����w��o��9��C�:���[��5��*�Zԕ���WBEY��D����x��.%[��.�G&���9YX1���b�R�;v(U�eƞmը�Dn�<�ZF��6�ٓ��S2��N��5��Y�Z��7�E2��Wmq��E�p��x�X�Ĳ�i�hӅ��BNS��'4p��Q��'��ȶ�Zq�n����V�5���Kں4a(���v�7�b�MZF:�`�X`�z)Z���S�D1b|Hp��#�n��%��"=�#e� �v"t�Q�!�L�`@�mT��`���aHZ͇
�P�ܙ3M��V�Ԭ�V�OB�E��R)2��E��]�ӱ-4�ǭ[�+�FAY����˰U�ɿZ'�R���%G��Ʈn�2�	ܖ��X9p˳K^褪DIȝ�p�N�}-��a�	�6%�����7�nD�Ү�[9�r�L�ZfE2D.;�k,P��724�̓+!�ԅ(T��J!Q��*7V��lvˉ�����V��Ř�Y�/w�R����j�W$�������.m=7��wz�������"�M+��M�wv���d��/RiU��f���E°6NV�WBK��$e���1�_ш�m'3�0p�|�GC4�0�͔eina�I�K\��E��}��N�	�36�Kv/��\��0�`Vo
s19�F2�0���C��J��e˶ѐ[M�,�n֦�!t��'	ANZ�b M��P��W5ٍ:tu���K�%n�+�b��vn�٫vjGZ1���j�h䨪�lIJ�l����8��GvV�0
W��[�v+d�Àf�8�
�p2@�W&��E�c�Ѵ5�InՊǻB�h[��A�����ki٧L����N\�nR���/6ZQ|6�3+O�!�U.��Fk�:ZS���3��k'�@8)�V�
՛�/	��Q�M����v���":m���F�cB��:��
�ڑ:k,�j6�e�j���.f�v�h���-n�Vr\���C[�{���YnݨuX��4#%n��R�����Re��%��m�Z`k	H*�-�KE�-fG(��fe�A��w����5%��0���<{F�b�8��u0n�д�]�������9ɴά{itP����:����5%�R�U������\`
`⧆�{!�V�l��܇]�N��VTIf<�н�wI V``9b��=���FD�
`��&[�Z�L���X�P��7-�Y���i����v�n�Ԁ�c#nּ3�R��.��2�i)&�X`g0)��&)��ǐ�A-�"Fa�D˕1�4�21j'r^cn�U2///Cw�̵A��XA�ͦ��Vw&�
�݋M��ءJ�eV�Ԧ�]dN7��y��[ŵ�4ؔi�@ Sd��@�R��=M�	��� �˘-��t��+\T��Ӷ�կ�j���-ٵ�;�&�-{bV;ւ	`	�b�,��`P�1���/C\�1 �h�қOV7��}@iV�9y�P��� �yZ�:�b�� Szh���Q��̋,}u�\��#e,5�<�)��!]��R�t��s��5��!y���H]�T��ȑ�x.8��If*++d%hl�����ǐ6u�I�@�g�c��<�� Z�̺������F*�4t��-=��R��Z��AU�'5�bY�JXƈ�euh8o4a�>�n���F7���_3��6�{r-�M�1̶.����Yt^���E@E��b�7�&"�=͏[�ˢ�`�P�4����DQ�J�ä��'�sf#�AN�6�����ò����!�Ͱ�'�Vފ�pё�R��A�2����;b�6����D�V��֡V�#����Ze�`��ro���f�@�<;SePwo�AP�f��+F���Ln}���fӬL���;s� l8�	��FO��sM�٩���$պ��t4�X�l']Gm�N�r��z��u���G ��X'؞����M����u���35�˳�fP��Y�Î��@���f�-��lJAG�=�`��&�n��LT�[�(�4>��# �!X��j4^���CY9�!��#Xo ]��Vhfv�	t�cq������b	�4� X�"<�W.�U�Y�U[iJ��l�ȴ!�R�a`�!ņ(U��j�z�ٻ�k�٭�Ɠ"�t�7i��P-�����<� ��k64�Y��Y�05�����kuf)[�� /�d��׷"$���jP 釦�L��24R���z,��h@�*�%�ػׂSa�D��aY�#6�;���b/5�N/q���-	0���[�oe�u�Z7c�T�UL�Qb:ʀYW�/�]0��7�LF���(���p��+6�8&�o/��.���r�N��n �(u��h�O�u�v�k'n�[e�Z��A&$�y����g�:82*7ƲS-�	aZ*�Ejđ�N,ˋt�JSҥ�y�)�����{�Ly}�X��
���{�@.��콶����H}[@�r�/��${�N�C�k��9N7P�X��UU���w|���d�R�;Ww��W�V�Ѻ�z�"v6�qt�Z�ΆIލ�+/Oy��)���Z!���܈H7u��������mh=ܘ{�|�\�Ƀ©޻�{������W�����ܛ�1n�t�X�{��̋���Uv�tB�v��S�}DJǔli��p�/�3T���lq�|��Ơ+Y/3���$])��p�nLdT��<Aw���ga|�}[x�{�%2�5˰�R���e��e�Zgo��̦Uv���mΓ�Ӗ9�4=Q��e�2ܪ���o9Ci<�ReBt��`{V�J䠻 Ѳ�#��b�CD�]�n8��u��Z��!�t��@gmL���w`=�s��W�g�+pdӽ�fc?v	��]�ʍ������՜���,!\u�)2������v9X�]oG}DI4����u�K�C���^
M�R��C.澏�#�v��	�93���F��.��v%0Hq2���NN���|!է˷=v>��>�}i�x�yp�����H�E�q��l�!=�N�fT:,�����3�}*�|�8�=�����{���J�صY���{n��aՈc7�::��#,���fQ&�O':�MAd%
�����Ij����%���f����K��g���Vj >��¤�����/�sd�ҝ��K/\\�Q,�v$p�*kG��+�-�#��<-ܫE�S����T6{���Cl��jr�*HTwX��K�17��ns��ξ�Mv�Н)�Z�2�G�`��0�5�����#xY�p���յټB��V��yG��ϋ��-3���6G���?Tp7�-��<;�Y���o��ƍoOr&��n�)��쮏��]�v�U��g,�i�I�Wq�0-���Ay�~�u�Mw%i7^t�R�I˜ޒ�e"&/��Ɩpv�$��<��7����Ak�*��ΗݬM��,�p�{+1wE81¿>�aiǾaKD�^�Ҙ�7��f�"z͙5��2:��VW�7�-��lhA͛uya0OQ֝>.�_v�',k�>��.RɆ�t%>e���$|jp�!�ŤΫ�w5�Aܦg��E�;�2!O�sݫ�t��p��a/�w������®��R�k�M׏o�ky�f]j���L��89)��q"�vyv�\J�Ս�s/���m+�׽�v����ܿhF��,�z2X*��<n�Ejv�;/Px7���h�o�<-�G.�qeK�u{&�»�M�R���j�A~�/��-=٨ꌇ�N�a^M{=�K�t$��wh���a���Q��4.l݇.���=�{N�l059_��r��l�%����hut�_}�[��?��0�Y��
��r��6<��{J /,���u,4�t�=lQ���z�쭻5�_�E)�n�)�">[yq	�����ڦ"8 4ɶ�Tf.G������c��oB(=����DT[��!��[)�Z��-\hr8"���-�9�%�v�JlC���-��O:ѫ�������mn�g�]ۦ֋�6�ɛ�L�۬�9�$]fJ���2�)op�ͫ� A�z�3�αK`�[�ad'Z��Vn3��Y4Mk�]ꥅ�bv��J�֦|���qoCZ/yQ\8�R��XP"n��j��5p���CՉ9Wq�U�j��|}����i�~��g&��\��ctv�"N��0����|��E�v���,l�c`������]��B� ��p<�����,b�<WLZ��4mrtvL{��"�H�`&�I�����r�)��|���;9��R�U���p�z�\s޸�6T7��|��ڻpVm��9ۥ���Je���&�("��K-q����m��Y�V��٪]Ε�)�A'Vs�4n$�}Ϻ��KR�?s��e��H�
��4.�ŋJp9��,Xb�ח�4�z7y˖��ϴ�AkR�J�eM!>��X�ڥ(Vo�M��b%KC��B������Wm��I�c9;M�<��g�_B�u�4��:���G���~��Fe�u�)�$u�=5�=on�>;KY�'f������]�&zm���rn^�� ����)�!fBȺ|��Hv�˕�#	'�ӽ�u�Y��Ԭ�ţ﬌��z5�͖�&������ ��+����C�q�R:'ct�-^,X�.�1��*�2��$�����u}��Vu���嘫�*.BZ]��:�ue-[j�Ҡ��F	��a��7\���n$peHk�58��3�&�����[8'���F�����%���a����K6�^4��`=B��Z�qJW�9��S���1Z��탅I�ۤa���pPfq��kWNvŋ��k����]ڊm��~.�d�ؚ׌CX%c�0��j+��[���L�;wI�|q���_;	}�a�܆D�U��yЮߦQ�epZ �j��*N܆��b�]�r\��je�EA�[�����iɍ�z2����fmΈT��f��`�W��ay���I��LW���?:�,�x�1g�:N5���d�w�9�Å4!`�P4���ڧbܽ�C���^�])�'p��a�Ȕ�/E�_>���=��/���Gf<�~B��C}���e߯�=Y���)u��G����ǣP�SJa�5srpI��,�s3����fvyv4,m��@�25\�I8HĶ\#n��4yMÏޕ��Ҡ/.[�͇Qʍu=�/[(ϰrw.�ޮ��]� ����ʦ��0�o�Na΅��u��S��[)،ت�f�3ԧ�[
���޲�Rn���U0�8Od����<Nϊ���.�⑫s^jX��5NoA�wv��6|��!.{�j#ͭ촻:5"Ǵ��WX��x3K��7���;.7{���k����$���e�7���t�ۮ�5o�s��E�:�rMgywo]x��64_��6��1��N桝v�y�;��s��(m)6�V@���n�*gV�Ϫ�נ]w�2�{��3�@H�ݱL���㖇���4�U�M�0���	��t�y{�/_*R�a����=|�V}k�ڜ,�k�0���u�腋�;_3��k�`�N2Q�v�$r]]q�;;#]1y��2�!��^S�ܧ����w�]�F�w9t���m	��Wi��e��(mEg	h��K�g���u��|�m�I�7^�wx'���.�{������"rtC�}��Y%����;3�is~V�z	Ⱥ���C��-K���~���Su�Y7�����k�&5��=�����(��UҹQ!�l�լ,\
�\��~V%r.���(�⟆k�G���cL{P��e~.����\o�ϝK
���Q��Ҫ'{/o18KAr��=:���C����Uw��78�ćwr����3��5	�א��@9mN�֊{d�<t��C�
-�-��lb����r�^��A��,IK���钏3;�C{q�E��n<����ީ�=�^�۳^��`�����xPR�w�o��㛅j�[�3[���'	��a5��`����*+%�����#����ݼ���LĀ��Qc���Ë=~�w=�� Y;
�
اw�yg���
�t490�@�|sJ���F��҄|U�0���~j�ݱw��9�H���ͨi�<6�۲qGՊH8�K�=���yϯ\����JOg\�*���H"��c�}Y�h乆%]�7�� ��F>�4�&�2�b����n�ac�r��K��9`hp��cӨ�f��P՜�1�dy9a���m;s��J˓�e��qR�a���0z�͞���h��yD�ny�C��}�q�qu��rS�ŋ5]�6�9f�Eʞ�����hn�ٖ�c���yqr�������~ӈ��4�~�h��޾�e�ZU��]�]��{�,���#���m+��E���Lo-�dk�\���!S���${�Nߎ����^���o!9�Soj4�;�&%����v%�гv6ۏF����%�{��V�p�^3>�$pƵ갉�+4�B���G<}ё5�su�]e��*�>��/�k����w��a����`�*��4�׍YZ�oivUl-�����&o\���JN����A`yl��N�]�բ&z��- H�lJ.{�^](��J�Wڂ�{*N#���v�ZwF,�ɕ�\���
����Aܾ�.�(�a�T�=5��QO[�в�ï.�=���v����K#�#Ι^:!����h�gW7�V�N���8����[
en�)9�嫩��3yX@Ӷ-
v ��mIE�Zx�e�����Lق]y.����	s�p7=�i�«I6�;�[w,�+/iA��6�~wtvᘽ�Ӎ��s}��\Ɵ+�Ѣ�r�Q�!*���Z;����V�:�o���'S����������lOW6qΞww��q*v�Tj���kZ�w����]����v�N�6`�ݧ�f�,f��VY�� ��1���p�� X"�GX۹vy���A�v�B(�W�,A����XP��h�r�0�Y��oo~��b��ew\o
��8�iӃl��@+sd���C���,e�� �+s�Ue:=�,��˔Qu���VlF���H������Z��ُ�f=��V�"�iݎ
�t�ӈ��^^r�&���p�j���!673HƉ�[Sz���W
q�O�ӫb�(O�����_�"�
8�[��HK���g�Ugn��]^���y�k$Z�>>�p���J���/ ���|C+�'p�˲ws/)Q�<���Q�9�v��g&"��Yf����hb��B]�ܥ/19��<mS����Z��֓����L�i���v���������⢂���Z+3���zw,7ť�'_r/[]�ik;�C��v^�ּܗ�U����WY8�˰�JlU5q�֙��}��}�-��0�eQZ���^tV�F����#���3��-٢��/[������|���%GG���)�P&M�e�F(�u��$t$��A�����BXZ�|�l<� �L8B��HM�~h���&^�i�6�;�c���V]�� 0��w�z{-}��8�����iP���Ӡ&u�2�����[p꾺�{����mW칢[V�
N(����ٷ`���Q��G��� �J᪹t��#{B�퀳]Xt��#��4�A�V��*�d!�������W�D�����ř|ϻM.0PŮ#]u�҄�ü�s��giH:t
۩��]25��X^�ý ���(������J:�I�N8�	K(
����]Jx��p�*��ž�w9Z�
�3Qz��c���+VY��4l��R�M�1l�5�m��@%/5g���|���8�$e���b��!"�6m��E�%V^\x��.F�g�^�ܨ�ޢ��k��A"���^�.�F��Pi�rgkR�;��t�O;*m�|���Vs���uX($E�?2�p��|�Nկ��`���nw��Y`��.�J2��ݞ>u�b-L�`�p��ʂ���n�V2	W@��;�����ٗoT�!�u�v1��-�F�'I���.n�͖\����ة��_#���ȗ�(�,�y%����l�x�pQ�M�Q<�)�Jaν�v^��ң+32t�bZ���Ӯ���u���ሢmňZ�ϛ�����.����]oUS���Jd�>Ҹ�
���d��#
m2���Q��{-w����+2�~@�^º��e���%��)��9�m�h�/�Ǜ�	�����Ky�RAˌe�'���H�6c&��A��<��cy1���v����}���P�1��Y#*8-=s)� ��i�m��u������8&��"���)Z�˨�T��jI�y^��*�j���8�5�gJ��c,��jkf�N��uvH����[����U�.Ĩ�ݑM��9WК�s�w�B��`=�0y�=d;��z����r��5��3�*.�R�qٿvo�����X�%����F���Zn�K��\͡ݽ�hM�L\�9|:�G�����T��7U[�ݜ��=�^�u*<���┎;Gl�;8Yu���mtS>�.2NȞ�L��"�9�Q2إ�pө�O �6�7��R}���\����3_Wؽ\�M���[���O�)�d�s���1���!�\�.��Nx�֝���l����ul�(��<�y�y@�g��k�r�UAӭg+�&mU����|1��3��4�v*�&���ܦ�8�SĠ��hH4���wf���f��s��)��*5u�i�����Ǭ<�'��j"5<m���;��z�����*��G��>8{��շ�f����"�/ms{��T���ﺴ�wlF�3�N�Yc�k���S`��]�i0W�"�������\�ti�}� ��PGe�#���Z�>Ϡ|e��|k�����ȹ���}5lvwso-u	�)�n�TCD�����E���#o�pJ38HE{�6��m�s[t�����y�r&��l��V�w{\$yxʣ�W`��%�����}$��4t�.��Z��{ט_W�P#�g���Po��H��#G��tW!�;N�>�]�:��E�n��k ��Ag��i�1al�+�������U18 Y:�|�󚔹0���#��s�9�d����7�>���{g�w��gGtԨ[��U�yۊ�I�NJ�U���U��Ykz�@[���Rp�s�]iJ��q�q���ε�I�	潺Ɇl�Q�p����Q ������xo�f�^}e��Uv��㚹��U������d[Myozy���R1Zn�]�֫�}g��+U��Yn�/Xn/+e?���}{������m�6���m����<���~DW�������WiCD�U�r�ꧡ��7vj��5�j�:�����,�c޸���;����z_CG�Wh�$0S�v�f���x3��j���e;XcgE�n�����/i���+��r�~"d8O>v.���p^Y���dr3Q�ö祰��&�A�ǜ�5q���ٸ$���|���ӨSe>r���Ad��寐�7�ڪ�m�g�YM}tw��n<�K6c��ZD>ɼC��\�1Kj��%�͹�sFj'��~��?oO�ݼ�^�m}�(�9$Z#�v�/XX��2�1'aZ�C 4P#iR@muS/�X��\.�����ܪ$W���*���"����z������4K�b�@����i��������*���Ys���o�\�պ��u4�^*��t�ɵ�^�Ǧ+Ů�3��b�J����K��0�6����� L���Qң�jh3�"�B;,�n-��pZ�+�CHM�	�i[[[�v�s���3�l��]�\�G�nY��K�nP
-�a�I�X[���!���l�!ӹض\Px9�dZ�M�޾��5�A}Z�tBNR1:����ng8������t�a�yIj�C��p��n�_)�\�Z�x��(����x�O:�VH�h�R�:��5
�v�	��t^}z�j&g<�6��V�l��{I�)����f��F�*4)8�}��Eb8+�y!������:CMiû��&A�Nh��r�u������(s�Y�Ȼ�C��f��LX}�p[�i[��Ց��l�ц\i��㒁v���)$��'p
�)�͌΁\ c��'�Ѳ�;�\{0���~�W�${H�<9�4��B�@�G���V���;E�$,�t�MT�a�Uʡ���P[X#���n����f���ʏ_j��ֶ��Ri��,�Jaى�p�k^���������|�V��mx��E���_"���r�)קb��b&7�ٓ��4w�z��C�m�hM�����c���� ���i�kcJ���W��t���J��5�lt��y�i"zյ`�PW9�?M���Qם�t=��QW�f�ᮒ
���^|{M��[YȀ.�=����Z�����oU���$�dD\9W����`����k{)9�Ej��;񌻠R�&��ߋ	Z�]�T�̭�6ՉMmi�H�v�����^>Pllסq�l'�jG���l��Dh�V��־2�ق3��(3w��Ok��l�7��B^�����ܘ�dѽ��ܹ;���(����=��/Ǖ}Y��]VθA<�N
�+7:҃L!̢�f�#Hư��}�J��[8\wA{�p�4��
z�C�����D.t:�}6�J�	�A�-���3ou�t�Ji�;��.;V�s�2�v�Nv���	*k!��`�卵ff�!�K�ε�ou �#�"�wb��8Wn��;5Uϭ�^�7��"g�N�US�'gB8��iu`�nv廮31)Η8��ㇳ,d��wÃt����-<]K�a[HU������=��-�Z�V�!xԦ=�ob��b�����.e
޺}��]����U��(Ց�0E����9���l�w�,��#D]���8�)b ����Mm�K\\/����)'x��;M�[� ,��<�z���z���W*�)v��ʏ*$��b��yp��%tOy}x@`��2�`=�d���w����:YNx�V�����R�{2>2-�KyJ/�i��"��[�缴�y��-�>LL���x2S����~�
e�ʕ�HΞ�9�>�@Qh֣�F�w���tB�_Q	_N�S�w(�HH��M��7ؚo�Z�sg��́��k	n����[�sΏ	Uv�b$c��z����-]#daz��>�r�k�> ɯ��kƺ���K�eޯ[Ȟy�dֻ=v\�#t�PgOX��kX�sx�g^�aVY"/�nA�)Y�x�Ҙ��,,�l�� �-`�m8c� �Gh��\�q^�/�萨��jrO{x��x,W%�f@�h[��x��qDC�f�D��0e�3�"�w��aIp\�0�͛�}ء�?h��8^���J+�C�h)�q�5�TNa�HU�V���f��_!)*���y|��wmԴY�&`�� s�f��W�Y"Y@�ob�"&�^�{	��*��W���)U���-cTvKk��s��L�ɻ2�W]f,Z`z`�[���5��nRj�Vz�8��=��o�Ώ�B�_5������ع�K˙4{-���������!/2��.�{O.��\��e��˳j��Y8�g*�E`j�f5�g;웃띚si
�|79��-oc��'��;���՝x~��Y4�x���p}��� ux�3��{4Р/�B\:�^���nq���n(��C0JMT6K��[�w�nӶ��G4�`�t��r�+TsUP1p�&�ܔz�:V���&^&�
�d���K�5����eXT(����Y�K�Kr�Pjj�[8�E6�ns
�c5�����ν�����f<*�X����`���m�Л���GRw��JՓ�YJ��V�D�2u8/u\�|��(�1HTK �rWB����n��3�N>�r��8�����L����#r�u`
�;il�W%�[�6���s�,��ho�f�/r5���{(:���(	R�-^��H����)C�R�Z.þ���yfa�b�����1���ŭt=�]�R�/t�n[oQ�"n�N��;z���V:9Uֳ����Z7E��/K��[g\ �4��&��������p4��/�2謁Ў�6��:&Yɑ̇l!�Z˂�9�i��Y�ٳ�X�d s.�NT�ÙL��35R�/g(�-�!X<�c�`�����?��������K���p}��pݧ�bɵ��Rc׼]�eH/{����H��j����,՞Шq_p�9x,>���1��5h� [��E�k��A(������e>�PKu-��N__��A��v�PS�}�|H�0ǅ�Ǽ_���2�Z �`P04
�����M��kxvvmM0J��j�Rv�o����K�˩�)�d�VkS8�A��;�bJ�c8A�go%�g]Cy�b�nowh'�_71����·�����+z(훭�Q�}��c�㵥��3�ҭ�!7q�.���)3�j�J��W:��I�B"��p���-q�wV�ؕ�;Z� Ruq��d�:p�I�I�g�#{�R��}�-<�
+����F��2	;)h�����a���q>�Fb�9��WM㚷7�X�R��v��n��N1mc���$���Q��{��s�YG�Q4h;x�0�HFbq����kv�h��!�ǆ�])Z%Bjt���B��Z�*�6�p��ԙ)�=~�wQ��pC$3�o���;֬�W��SƎЇ�1�~)>�41ƥױ�򉻐
���k(`��ɰ���K�7	^'�k�3�n�e�h�u6�JI@�;N�]�5k�����j9�z; �w������j��k��%���9bhr�V�09�vYn�L[���kNXV�wC�u��:y5��@ҧ^�*}(��%�.�4,���GmL�W�;&�ۼө��1\~,�"�*n:�$�Z���1|�t�]H�kW�dY�`_gf���u�k={"Tq�̟rM�.
�-�k�`x�zD�Ze�*�Dbێ�L�޳]m�t��^i�2�a��r!W4we�pԶLެ�gH;�U�-�L�V�O�]A�B�X��d�qY���ټ��W��Η{�YY�8���6^����jE�s�z+���t�p�HK�t�h(v�=��m��͐}Kqg/�o.}�N��@�o�Mښ��C��i��yܕѣ0>��ҵ��z�c�5��뷜�u}�ӐX�S,�ֺ'3Q��"�	}ͻO_Q�At�+�􅒥�"堘�+���F7�ߺ���f@����1˩�gc����d��	w3�� qT$#.h��J�4y�}�؁���̼��X��	�-ۥ>��K�6��s�ǖ�q)�N��ӫ ��R1Oyޚ�%����#ӍރV���c<�wg���T�X���VN�v��Y+��7�"��|�0rżSuB4�x{�PH�tºf������>Izzjk!�z� �S�ک ���δv�:�C�K7"]�ϧl���o2E�E>j�r�osaV`��X���ҾӲި	v;Dըl�)�*��w�l5i��ܰ��;h�/a��� xJ��h<ʵj��=;;6��G4��4k{���m@o6,|�;�(pB�U��N��+��P�xꡛ�P=�G_=ߙ��4�Y1�g�ܢh����U٦�\��u�.�k�T�̤1 ��ÓB���9G��!�+)Qz�K������*�B��ʝ�������s/SZ�O��|E�vi�p��KB��d8��F�j#��'m)gc��K�wN��a����mCn�j��~m��2Ё�������x���ghZ��-�����٪�烣VE.o�J�[�_��6����$w�tf��"Ou�2tun��� m�E²�qwZt:Q�|�A��5ȃ*,��f�,�Ιx-dz�Z*������'R�7vd��i����<�)�t�)���Y���=
�L,����0K�=>��g
�o�v�я(��)����7�w�����80�ɶ��/�P�;�wwʃ�DR�M����1���r�M0���J�й-5��
��J�k��������W"�e7���
�cUu�+�����D��\4f�m�ǝ�#B�n|��]=	�w�k�)�uI:n�<=�@a�}O��+�P��U��
|vbx��U�Դ�r;�:�ŁMC&�Q�Cq;ud.WQ����%�b��� ߈ߕ��^�ޔҾ*���su�h�����wD�%ZKOGr�I�#d",<�y�`�(�#)�к=��F;�����n�F1���r[h��b%����U�3!���}�^��-��X�q��㕟pg@��;n��6`���r}�^;K)����2@|���'4YEJ]5Ug��w���XYS�5��b,��!o9 �	R�+j�S����N9��NMH.9J�-�-ĕ�}�z�c�������˶`�gvҌ/P�p`����Iz��1�������w`�{=nRf<����Ր�0U�-9�:��H\Z��):Qo&f�����ˏS	� �X����)A;h܈�,t8L1n<ƊjLWwq���WX�'n�Jm�k����Tw���4P�yU���9Q�gEĝ��d�=q��`|c���% q���"�)!N�	�tzY33 ��2���=���k����s��p�x�;fv�n��,�I.�I�5��%����b�L��GݛQ�0��㨭��T�4y��tv[��"�T��fK��Ǌ4�Ib%ޗp�ogjb=:�T�SP�t�{k(7��m^2��F���ܥ�W:�,��>��K.�Tx?�!A�+V���Ws����V�^dp����N)�wȀ�ai�<��Ĳ>�&
���`���"�u�U��V�و��x��tVR���*��N�I�"�W�.��^�I��y�^eM�vڔ��M-���o���M(��/(�;��隅� i�&yQ�Z�l�h�OU�z:��f�ո8s��sj�<+.��+���-�R��	��'V�:k�\���*Y;V�5�]˥�e�ѫ�s:eH��:��D2tc��P����{��{����̷��s\wyr���� %�ȕ����rB�](+�Wb*�mᗃ_���x�C��g�m�:��uݬP�X�F�pU҆��0�������G.�xi�i g.]�uK�s�*�4���U��wm�z`�)
�-e���Y�<��l�����{5+p��v�७m6��ul����;��w}L��,��L�nձW�9p\�X'S���t;�лB8��=�������W�wK�n���-s6�+�!����\�P@�w]'�-v�c̝�B^}(.��Ԟ7���|�������C�,гu��; yR)Pڂ��G�oC�jV���2Q��9(��N�ݝ���Xr���X,���.�5��_����!�o�b,'��1��}!�N�"i��7wOi��W����w*�ˡ��D�xj,�Â���x�T�8^�L�o{���%<dVmDhnqB�0:�T̰��(�rr��Pi){s+N٢2s��~'��G��Q�ǥ�=rS[�!f��\��pO�mu�Q�D���.���p�x�r�U��/w*4$z)��"a���\����=�~�+�*���ܜlw3�T��-b�Op�p\q�� og^`�2.%1V�3թn�a��L���'5�W%r�@�*Yd=�Z45i�fR��ܶm>��R�yY�	aɭ�r�[d���6,�[)_b�Ԛ�5��R2�\����.�#����"*�%�8�����c�L�G`CB�����|r��##�%���:����5��ita׭8ކ-�W[��.$��Ą{��2-�j��ji9��Iȝu�O�����E[8!b�p���4���bR��tmK�u�� �\M5���6J���v��n�iq��t�x ����}Q�5��Rq��4��G�<_q�Y|w@k#}�T�gMcz����rރ��uwUpK�܆�<�'�	J��u���XcV�9K�J�
���̅�[�۳N�0����\k�[�Ѣ�;�s�œ#ߴQ��KX�[E+yЃ5�����g��Ie�[h��4J�u�e��c�i�u;Wf�C�X���˲q\u���vX.��#X�	����7�e]���wR4�#*���>�U��7m�`�![O��O�}�}��W���g�u;.s��6{��C��2q�2K����44����w]�&���h���Gl�6��T�%Ǔ��rI�e4�v�~��W��{���>�N�(3\>�kpЅ\̅[����r��v�bB��d�u�7���v����{($��N��\'Y�z�%J�7M`�k3��ȈN�DBc���;Z���z�e�(��MN���C�|�D4X��Bw/�{���yE2��3�����Z�|=��0�c8G��n�;*4���i�sj��\�ʷ�O7y�*��݋(,bv��m/�؄0���Ozo	��v�����t�ɚ�Q��r��ޏW���퐴5�#�c�vz"�!,�&I���z��g��K�j�)d��)�7!�f� gm�ݶ�֓/'lK�+X���n�&�փxN\8�3i�yO9K�jn���R��IQ�ca{��>�#��'�I��dݞ/z��P�.)�������w�
�F���a��]n��ge����K����'KdY9�n�V�����q�vE����s�~N����A��lq��aqu+$��wǹaJ��t�MQ�m�X��t�R�K��Љ��e���+�A�x_W�`jd���X8%�9����Y�� �R�v��u��P���xz�4��A��L����=��?'���Y2����t��]���Tz�a$�4~ U���ML�j��	$HQ+���U�$T(��ʼZE����u���A"i��"���auMTE�b)(&H&KU@�«4�S�HҺl�� ��E|���ebef���$�*ԧt"���<l�#D����j`Va�d�E
ȡ$x����R�MN��F!�&d�s��r�uZ�p�0��E�*Q�	�TD�ㆁ̶Pj���Us�rY<×��j��.^�TJ�s��(
��N�Axʼ�)*����\�օ�$hXdT�'��T�$*�/WE��N�B��*оA
&冕�B�s�E\*�HB"�t"��8����ED$���_��
�B�h`�Uʋ�QQVr��
�x�>";����AfU,�C��Vu��(��ȋΔ�QQDr-	 P����9�t�J���Σ�(���Cw�oi���E�G�J�S��򸬴�k#$݋]-�Z:�9��S ��`U���q�Y�>)����o� �X�w���n}h����Ύt�{��nJ��x,�}�Nꩠ<q��专uC'��⯒R2We��;��a
�b����:�g�I/�ݿ!Tc�5�\ƹ���y�/��~^�ώ�ȯ��]��Տa�]��Bề�N�zwۀ�\\��1a���R��o?���^�J�m������>�"�G��Ӎ�T��3O�!Q@$*o<�_W��=���	��n������P�Ƃ���܋�FN��|�X!Ri�)�x��U9৞ޔ*�y�����z�{(5(��y^����a��{%W��îK�'�\��K| �W��Y�t�m.��Nu(�}�'�����$;��)�H�t@o�'��|E=?u
���/P���`A�>O\j��^<�b�n͌gК�3iX����b�t�v�f6~&�G�%!�c4�Ҋ��Lf4֔gj����	��a�Ş(O��׆O{�xJ�V=`�t��G}��
��|��*4����.��^<�=X�aۀs���yﮯ��-���Dn{HQ5�[xcյ8OۀNԷ��9������ѣϱ�2���!��2F�C��!�l���:T����Nw��H�9dQ���r%��8U��b �:�dh�_!�R��.��Z��-F�p��kՄ�1�>��ޯLl)���P|�ƽu�Ln�B�ȟw�h��/�������Z F+�)��O�X���gª3&��s
�I�?-��ogi=�P����2vg����T�(c���`3j��d��W�x%j�5u�Yh (����h#B�x��Z�OǗ�����P��HiH�- >��XU��xx�rn$�:mE�^�����X9�X�G�j��7���5Z��g�K�w�@LnU�xۀ55f,��0������u������o��{��yXG
�|��3�x�&��9X�����VV�1�ڊfl��X~�V/Z���ͣN���N���sb�{���t4G��K���6���|��s�O��-0?�+�R��[�ۂ���T�� �9W�}좃�,�J�33NH�����z׽���H�d$V:Y��mT�r>�yP���O�r�A��yc$�r|yb??>IR�S�P�W�`��H���	O��J�J�+ڻ����=1Q�b�����Ꮃ�'U΅A�i���6xw��)�,�2���y$||�e��H�zP����	�R�0V9��SD���{|��S���QVE�Gs�a�b4fY��o]R�Q�}:�&���u�N�w+M�9H�ja��i0�T�mu�S�̖#X��w`AϻWi�ib�دi��;�7c�m���1����g�u_��E�;�JN���8��� ?R�"�[:#E��}��W�f��W'�
��o��b��Lf�;�S�k�<y]�w[kԦU������>�mK��Qxu�!�9"�ڇ����Bɛ�Ď��F;��J<��S
��Ϊws��r�x�oj����E��()Mh3u[��+wHm��1p����v�	�`��[�8eS��Ǯ�s#�mq�j���{���Yo��w5{�\���>����?�cѵ�cKExJmxr�W���W>ʽ,���u��f�j	�3��^��*� �Ǳ�b/�wX=]ڮ����r��}�OH��P6#D�7>�[�2��:`���w]|���7��8�>��m���%{��̓�vlǶ^&,F��K̚nl	mߊ����H��U�LGs��c�x9��,�͑�M�A��"���f�,�4�-���L74 ��R佣�6�ļ^�IibT���.8�'k�)�]�{t�4o��3�c��Y惔��G86NI��#�EY����d����K6%�4S��Lz��t9�!����$�hVlP-�du�XWhK�K
nԻ9+�<�F�#%~��Y����,:��@�}�r(���m�|9�e�йF�Z�?�?�A���%�| ��_X�[�H��m�f�`̡�p�U�FGp�ٕL�?�p���W��M^�e�|/m��ه�pm�5��Q��(Cz*~��^IK��p��0�vn��(k9�Z���w^�`l���E�̐!�������1����U"�_�qX�J+���/�e�^�^'I��x���*���\�� i�U�7�[u�pl>f�}�+��"&��=ӫ�:}&��n�:�p��`n���(�����4'Է���c���,h��`�q�צʙ �j���f@Z\�'�;��T��2��g.��:F�3��Wr߇��ӊ<v������5�+�������=6G�z�5w]��pU㙷��`�wQ���\^4�v|3�=�˥�/T�ù�:�=��v�~�.�pPtK3��N֩�,g�ʀ��r%���0�&=�wV��>+w+7|���4�K�>��YP��7��\¸|�:����À�	��/��J���ctPѹW�Gnh��8���e<(n���4�
K�gsV��"���7��ݯO<`��R�!(����8���|$����W+3��+>��lf-�`u�������};n�vvȍ�T�'��}�ZOX.wL�m��m�w��B.���ȏ���0Y��COO���c�/[��{�KF�>O�U����[��5�0ԣ�~�{ʰS���K%?Hz���#+=�a�G��j���EǛƂ<i�~_�{�%�5<�X�������/������-xY�z���{�՞S-}9�;��N�=�ٮW��<��1͓��*3owFi�d3�������� ��]���G��g�S'�ā�^�G\*�x]m��W\XwgOyiU�3b�Ş׽��\]*�}L�U�u�N���bI��-]�7��ب*xּc,y�P��`��]��09��
��l\�1e�x�'���|A��Rb���K��V���1t��}���Ӻ]c���j�g��|߂ۥ��:��X�{m�|>}��bI^��*m��ؕ��?x��{���|8 5R5���W%c�[�y�u�OǮ��z�A&�B�88�mg^W5�Oy�{�r��Dӆ?/Y���O����)tǙ����=5�4�zbuK�����8�	֛�N�h�e*LR�%���>~�5�t���m�j�r�۹�(_QU�|߽��/�*�g�̌6��7�*�*��WL9�:�ꅤ�2�뙃�3yN�Y°,̃��ѽo�����>�1���:�"�`l��I��1���qxׄ'�+��a�.���
� <�g]�٧����{:׻��f73䛷碌ᇉH��������~�07�|�_�����
�!>��|���*��ͷ�,�Ҍm�ϓP�ʮw0{ܭ�E��ӛ�d�*��4��zfN��W���o��������UѲ�ra�-҄�_�xd��W��������L4�
�t{Z:�����5����^��w��~�t�S
��0��,��?Uƹ�!��jN��x����^�߁]�����O�:� !���Kx���=�}OWʇxؓu�>�vzR��������Vm�~�g��Ǿ��ڏ)C�=�_U�hh�ϭ�\/c�+Wd�Ӷ��>�"Knk��gfԴ��{�O��JU��ܨq����kA�G�;c�R�X��C������O��u�,��s�}qx<��V�I��W9�*+�P����!څ����xV��J|[��>�s��j���F����e�p׀�,D��Hr}&K1PL!{�F'}<^�W��y�K�R�uh�]So�$��.�5�_�wL��ф��^�f$�ѣS�:lr\�I\��=�(���]ˏ��+
R-���o��t ^�K�7~�rGW�6l-���,�䴾Z|� =t�pW�Gob��e�i���>a�My�v��?���K�yz�z�ع^�l�\�wu������'k���I��"6��Y�����x[���+<�U�l�^�����`�h�tZ�9#������qv�/<$e��u+�b�Ef�W֬$t1qr�D�s�Q��cMV
Y����I�%ۦ�j�A��?y�~��އ�i+�CS�1|�EV����J� ~���f�ցx׍����ʷ6y�=��wr��	����ߗ�����(kčzv��ŏf��J��:V�>��V�K4=�p�j2�,C�\���MW{Uן"\���p��*��xfu���<�#`�����C�Uy��\6��Y�(-�ut~�c�r5�!a�[$�^�}���k��o�
b�O���|��Jk���V��-0���{P���?N 3��j��yl�'�ˬ�}���=v�3���ҷT��޺��0�
���؏��lBn��x�z	�]s����yT��V�']A�,�@��q�¼%SkGJz�����n�Ԧ���ؽ�t�g(�E��52��eo]���P��q/�B��[�(X�gQ�@k(��ix��{���Zڹ;m��9W���J���f�e�V��k�ٕ&�Y���g*o(E8�t�A��(�-L�e�gE��c�)�}v����onf��Y�bǨ��#�_������ex�O�� pp��U�B�����8~5�׬�r+re=�e竓�)ۼn�Yp]�C�{�l7$ZjD�T"tO�a��- )P�?oA�e��_� �L�/=����T�L���g�霕`��J�L����%/;�B|���j$v����^߫9W���7�@3��!<tS���-�rщ�yE�4�-�ُD�sL�j\JEя8*�>�3t�mIp���HC���t�Yb�I���m��>)>����6N��s0�����r}���:�뜉��m��C���^N�&x<�b���ԘŨ�������ez�� �u�LS�������r�}��KvW���1��V�g�r=���G��v�<y�wX)�!y�
Ѷ���~�mw]}U��P���¹z|���Rݥ�gr�Z�Lj�=ͽ�8L����Ws�½��Z|3�g��k�a�0Oy`8r����X��Hy��qYoB�������i�>���*�,�BRޙ��ǅ������O-� M���G��T[^Aaq�����߀2���^���t��[Id�s[�>�XV�����aѮ�og��ku�+��[��Z�g��.�:.)__6�ofq� ��4�:�[`�yO�'*3 }�q,M>�b��8��\��;&0@z��8 ��b#z�s�eK���qZ߼p�,�G��M�]��Wj�����G�ߜ{��MzL�9��'��;�+��d|o֨
��/����zc�s�������z�s��ɺ��h<��r.]׻�h��Ǿ�b�u�I�^G����X3�KeM)�D�P�X������n$�X�hf~[�S����{,cQ��*ҏ�~k�V��B�Y��M��Z�����~͝�sD�0+f�¥�=Ћ�g�SM���f�yTX�ޡpt�n]�>(����m��W{�T���C�}t�;y~�d�;�U��O�_�,��'=䏊�b�t�.R���J�
�Y@y��ѽ@��F��9�𨵹M��M����e��/��M�7:f����W�P�ʕf�����d�ta�*�p��dpt/����ۓq��pX%�c�N�Mч�L��;�����G�gԵ2{Mה|'�}��V�r����p��ez��1������X�D��0,�V p�
���$����N[�獅��	À&�S�[i��ϳ9�����P�q�P*�{���������+�<����x�g�s8�I�~�2��"~=����x�z��;[G����N�Yf1{��$�o��N�mս�*�ws	���z�Ԧ�˧��v]1���%@��V3ws�v`�4��h6݌���/,�t����#+����͋�Y�,���B~U��~���L�y���[n+<7�y.��u�V� U��y��1^B�_�9W��->_�Tw��i����޿���[߬I�Mй��\���G�s�\<���+��������������r�:�,O1�+�#�mm�Ts��U�#D]�TF��(y��>A�l���5om^��^Z�jY��좟�f���ws_�Y��{��9��G����� +~���~�8��¥�=G�����!�9�*R��k��7U"��.˯'��)麡]C���tx睋�����#{��iwr�=�;��gS��3W�z��7KA'kf|4�)\b��U���v�#mw�۹t/.!����պP�f��a�MY�eX<e{�d`z{!��"o<n�{���<��[ Di�S���eu�i{�d���AA�ϫ���QL�y�{��m�ͭ�{f^�zUy? �� �]�|��4��W�w��+u�>���tS3����3��C�	��[��ܹw�]0�qau���-U��Us��2���BC�K�bbnv֩�<�I�]]��F��Ũ����5e�*V2�(���t�jm��')�k��,��m�W�]~�/v #�$*��0�{�W�b�5�[Ϲ��Z��:�D �T_t��8�'sc3��t�v�ޖk��&�5����������[�HM�2�i�x���1�k�(��,k!
�#��c �w{{�;����kq���c�x��i�8\[���F�W6��'�vt�ܺ�S�i�3�c�3>�e�����d���岑�&ݑ�9ӆ]����4����]�����kB��������:ө3\M�0�AO{E���*}�53�n�Z��T��b!�V�$����gubœ6��]ԭ̏hhQ6���&�TG�e�`U�ž�{���V��.���(x휻��Uݢ=�ĹmwH�[U�� �>���rw��l���~�n5V�nv��<��pj2���j��&�R�o	ځ�:��l�j2�-��7w;kq �V�O��Bk�	�l/��R�L%��nP�f- �R�ܤ��6ޢ���G
�oe.�On#�F�Wm��v�v�]ю�� ���2P8�_������ٴbтZ;W�ypv4�OE9p�+���3/�V�u��Vܳ\0?��:@�q=�P?%{k�(�np� =�B�f�^.S��N���tW\ۭ��Q�u�LX��!w\?P�����X;V�����ڞ���N���i��@�1����Ȭ�1����;T;�1nwa�_�&t�K��+��\�Tt�D��XQ�ͅV�/A[/z�KޥZ����q]��T�:+l7��FP㺢�%�G�O�wS���{�YxЭ��j ����M���F��o`!�u)|�pE�#�
�*^������[Cs2�|�z�{�x-e�H��󣙼2�K�v���(�YBVJ����M�Y���h)Y�0F�`s��V�X�z�]���7V�86rV,B�o.$,۬S�����up�{Ǯ�L5�h�&�N���.�s�����6�˛��1*��Ap���z/ o�Y�:;��m�fi�Xz�F�������+�H��t=��إ����mebR�2��쩶΀^��	�At4��]ƏV[ų�u�i�M�tᨶ����tw���{+k�4y�sn�_675`��������v:�&v.q`W��[\�wW��\#�~���vℇѡ�%���6�<�r�Ph��e���pu>��r����..mժ��B���5l6>5ǏN��n��s.s�nFz�]!�'�T�u���95�+6C][E=�Bz]k�e<��Fw9� @��Me�[�p��+����Ж{,�&qH�� �e����l�jS��x�h#�mg�۸n{)���B&�u�W��I��L�3��4���-�����NXP�g�r�1��޻??��\�DD�B��+�꒴��_opH��Es�F�\.s��E�A��2����ЊQʢ.A�W���G)$�8z#�))�����TÊ!t�1US\�8P�e���$|���9�+��%J��L�9*R��ZY�3�TTW2H���U��B�<���!U�Q�EN����dOr=�j�aBa�<����6U��R.Eh��Ԓ�2N��G �"x�W.��TEvEQìʩCB�V�bPS9f�Qʄ�Z��9�]J��AWE1L��$�9�E����B%��Qs�R�W��Ǻ�ϝn2TUEFd�*�+�Q_^���AF���W(��Q0�ⵕs�ZYZ`�*�
�(�(,���	��E,���"�6bdi-F�F@
�I%A� �[��¸;˾��L�⇛�:v�P�W!�K���0r/�Bx�MX��75ܹ��0��x���];ތ(˂�,��[U��s�_�?��q�;��WcӿS�
�߶9$��&�����l�C��߁���$���}t|�m�I]�x���MކM��;~~ޜ~8�.��W���P��6r幀=<�q\�o�����?���v�NT�w���B]�;�����x����`��O����;����I���d�~A����yX=��]=���I�G�x��� x�rԕ��M����ϋ��ϗ�=�ߞo����@�ђ��,Dh�����x��k��7��w�������)�P�w������bq�?��zOI�������i]�{�w�����p#�T�
�PW����~����dsuB"~_�g�P}N�캥uJ������ߐ��w���bO
������	�����|��Nw�������N$��o�oH�!;��;+��&����zC�W���*�/������Cꔧ��,�'O��^��@P��>����A����߈^������yǯｿS�aw�=ǎ<w�Ʌ��~y��S��z=���l�C������UAD}�
�����!UDQi��ۂ�[����U�紺#DB B|DEa����G�����N}HO�oǝ��'��'?��S�g��M�	�v������|q}�S�aw翽�����+�_�S UW�E|����V��v3�s}v�ڮ�#�?D`C��A��P��������=;���&~G��I]���}���ra����2�!���P|I߮�[��x��'}v�|�p">b ���_}¬��G��-T�:5Q�e��^M�S_��E}b�U����1�|@n��}��Ǌ�_����o��O����>����c���!������I�܇�s軏���aWr~!ɿP�~�A�#}C������|I��O���w|?�z�~\t%כ�A���""��*>��$��w��S_��}���ǎ���8O}�;��w��߿{'��bWo�c�~;�M���}���C��{;���?�w��?SӏN�Np|�~?Og���n�h75~;��9~�*�V
�?}����Hy�}��9'oｼw��n@��=����>�H���97�/��w���c������~;x�^ϟ����v��������ߨO����ժ��������h�f�h,r>�╃�,�:���L�FQИ���J7�)]����)GK[�P����̠9a��+�7�`�˝=Q`�WYo�ٶN��o�=�XK)��Z����-�@�O���򮂾��*m�}���H�Ӊ[ӧf���e��	�X����dYz����������Ӿ��>�z}����=�um>�w�?m���{�~��=&���:q��� x��o�㽧���Ϝ���H{w��;/�hs��Ͻ�������B}���v���Y�T3ُ}7��w�|�;c�Ǵ�+r����ޟ�ב��M��M���Ϟm�޽�=��7;۷����{����|�F���lS��0��f���^׺��c�raO���?�!!�~�����|O�睽 |I��׾����ې?�O�Q�o��Ѽ�C�>����#ӏN���w���zv������Ꮰ��ٻJJ��}��U�0t�c���D4��M��O�p��N>!���}������]��A��8�|NM���Ei��z�0��]'��������o�x������ɾ!;��z�zj���US�^Op�m�K����������N>��v�I=�}y��?w�|z@��o�ߟ�1�nBS�ｏI�#�������۟�����;U��I��݁p{d<�����F��~>��~�*��~��ØaK��{��麰����}�����'�O��߉�Đ�y������v�:��	2�C��~|��Sӿ���߷�oH���϶<��r|�'��������q�I�����!�|@V����K��pY���|?c���럮>'�x�|�5`���ۼC��������zｽ;ۏi�Ϟw����|BO�������������@���?>�����n@�DH��!�AM����W35Mu��������}ߨr��|C��ݏN'�8�}��0����?|N��N�z�����ލ����F'��w�]�ra}o�8���~8�}NC�>���E��4��@���E^k�>q[	��93��پb#E��B�t���}�~��ǟ{zOI�	���;�I�BM���x zq�ܓ�$�]�w���
ğ�o7��=&��G����z�1:�8���q��$D����½�s/S��5�����w�[O����L.�~��z���A���ӏ�X�o���~'�I�S����zI�I��?�x���C�x���~�㿿c�ĝ��z�>��ގu>����u��󘥺��
o�Ǳ�8ݼ�KkH6b�ƺg�e����~��c��8:�N��<9�w���r���G���7ص\��W�N#)MdW�h>Ƀ���'{��;˝έ�����L�\s�2�|u@5���� ��-��U�2�=پ�۹!�PX`Z��J�/$�!��>�uIn���vP� �3-d��g��t=.x��_�cG���3�
��߃ۯ41׽s��Q+=��yc��Ҙj+)�}c3�����<����kB���h=d���3��~�^���v`�{�Î߇[�w?Q-����3�	o�)T��8��c���K6��|�߭���r۞f��ӳ���Ru���,i���]�����S�ħ��<G���� ,6�ұnj۰�;�,���3~�-	{��N��M����_N/���tҽ2� +�U�<6U� ��LvyV����'Oo�5��^��W�e���P;m/�\I�U��J���ʚck�xֻ1tq̟MI/c(���Z���!.ԉ�Xʨۘ!٨ײ�{�>��E�D�|tK������8���v��׬�텷~�w7��������<���]��W��k~�f�y@U���5�س�en�b�jNA�<n��6j�V)1��#6�Ѡ��+0�ֳ�Qb~~s
�^�k��˛�J�u<;ٍҨ��GQz))�[��)�zu����������ټ��r��7�%���.��.c:��"v���,>����'d�Z�9|0<�H.;rX���-��ܠ�s/�q�N�R�Jn�m�lM�6�����V;@P�#ߪ�ǯ�{e�yͳ��_R���=���j���bb���e�=t5�皣�(7<g��>��m�<7�p_���I�B�aS��yԶG
��]~���>����Dx�{�7ӆ���X8��V�?���ϖ�Oi�(�rC)b��G\+��{o�����%��7ϯ}����M<��^��� g���{�x��|=�$��T;a]��ȸNL�i�Oo�;3�3���*/OU�Ѩ��r�dz����QD��{L����7����7ȯ���عT�1�K��n}��y
��<D�v��Gֆ?s�V��g8��g�*Ӟ�[�k���Cn�������>��[H��*�J��x}�י�x���MP.�'%�}����4z�uڂW��u\����A����x����Ujޔ>�aL}uHk�����	Q2^��o����6��Y��~���eVY��ў T9�X\���D���tU\W�=§�N_�o�����r��	��C+�;~Yo��X�x�y(?.�ױ�H@{�[�`v�ݓ�oK��r��tv�A�T�	����yJR�����^��X�8�Cv���W]��܅�e&���Mw!�PM�čC{}�;x
�2��3oD�i.�V�-K��ɰr	�sP	�{�	/�k��5�}T�GP�oE=��i�
��9�f��z�Wt�����a����
���1N��N�lχ]o�3��mkJ����K��zj{�&اH��2�:��W˸�(_�xg�Θ֗��Y^N�ˊ�5�K����m쭄괴Z/)��U)�[�)����E0���t�w#�ޟ�ա�NFFvǧ��3xV���xϯԀ�O���`� �t�D��b��zk����Lf9�gs�.�������#G�P��I�?L6�x�������ڀ�j���ܺ��V0{A1o�b!.�tJ�;����X�3�nP��t�F�|�@MG�e�o>(���O7�F�����V`��l*�V��]j������"}�V�I��6��O�B�L�%�󝹹W9�����*nt��4}�>�^���ʼ�D+���>�595�.�@X�34gXʻw[�]��o�_k��#U����||�C�ɔbb�|��.-zU�e�u�v�ӭo�-<:~s�'�4F�Q)��5�l?�+�T�Zř���VV��yQ�?8ܝ�[r�^��D\�V�°e'k�a�p��݈^���B�S��s�u���E�=Z���w���_m��n��WK0ͻ��PĥgQMNԓ	�`[ZX��+%`}$&�]h�ٛ��x�F���//xW����w�����Z��¶�_B�����ﾎ��bL�;��좇�z�m��$:��.�x�yVHe��	�[xk��u�b�;����w�{ �{����(1<������^�d�׎P�a��Qү� �e>�%J�+���uww�l�i0���<�72���"�<�ECk�ػ�͛#�Α�D�<3��_rnoW=���U�U�������,�%-|+¹	y]�b���::Z:i�"�WG9Ow��v��7�[��X�T�� 4:�5���Pt[(,՚N�b-�j�������`}��mf�fh���9�zy;+�1V%%�O��R��Z���N׻��hT��ǫ"c/D޽9�U����ޟ�a��׼��ӓ��V��4�ä��r�78k��W�.��rڝ��6{������>f,o�}��P�}'MG�ћ-eu^2�E�g� u׮Z��ox�"�.�n�����8q��9v�3�{l��>�V|�� �#��j{Ҡ�𷛺��{]ҟ��<5��O�a�½fW��x�z�Ɋ6x"x:�Q�qu{���yC+<e��`s������Vüpx��{k!�X쮿���ɹ]MVu�\�M��g&vn��7��#��8߉�~A*qXe�l\78=�,���"py��
�qX7�׸���q���?��1�����qHI�s̩2��F=T'~�������<��l�~PM<P�׊���?[�äō��5��P��*눀4��[:�`�w���u��Y�~�D��^,���	�?��R���~F'u�}(�`�ǅ���m�A{�ݿ\�����ĉ\��e.l��D�03��#��\���/�m��ږ7YX�aҋ�W{8�Q4R�8 ���%�A��yT�2=�D�4T8��g�y?����<�K�ݗ��.�s��`����:��qS���O���hk�j���%c�U&זv6�����	�^�<��}�ք=U���~��3<��]��=��C{�>���)ױ&EYp�z�y�ثڳ�����՝�|�A�U�f�@y�{Pz߆��g����s��Hm����q�4k
&�W�;+,4���=!���J3bS���>�<�g��zg�����ӹ���O�7e�����y��y���V^5b�'�N����)�b��<vZ��:PNx���z�Ζ�w������A�-�6<�����6y}8�'���J�� WeZC�^./�{ܳ��j�Tݥ@ԙ��^T�k�2 ]����Ȭ"����':Auf��)<�w����l:Y��0RJsʿE�oBꉞ2)�x��hp�M�ו�ad���^V;qu��E���4�g#G�����)�e��Ŧ��ңz/�<y�+�Yպ�s�c���\���_}UI�ʫݷ�<E�O�m���_;:�xo�s�3P��������oLz�J�3v�ynOz"׼�\����rV�.�j�|{��PC�ȍ{,g���ueQ;Pt`'T���m�E칞�;ً��~��}���P8{�*E����<����DW��b��4��a^D�[[.֑9�j�}�j��<P�n:��
����)��5(��ắyV��Ζk8-bǼ(jG	�:�ٺ�({R6\y�6b(�5��@to���>カ���bĬ]��5(�u���ޛzppm�������R��ё�^D�!(�
��_�V���I�X�in
�QzN��|�'\iV~�$��
#\����h��$��jC�*�l��Zw�`����V_��*�z������xtx������ t}L�^�^%�����I&0���X�3o���yO+�����o�R�Evy$]����| �{�+<Ő��T2��3���15������Ȕ0w�?vT���y�Py�y����U�՜F�.������^�ݼu{l��c�B1��>L`��)��%�+J�-�+&��xT��aG}��覛{w�#�*��X�[�!3iS�Շ�/{pպQ��!��,�0I�V1r����0���eKܣ�-s�W�{FH�5�%�L���W�W�Ug�xb���<^ӵ��3��ۡs+��~!��<P	�J��k�k�W�I�~��J���]����{���=�7�4,0��A��ϼ����A�N'eq�#*�<�xxF��5�(mku���x��z�QZ\k_y½�\~Kr	U}l��s�w�4�Y@����f[��/�qB���- /��'�25)��\������M�<(^�_x�o��k�ZJ�/w��t��J��\6Vy���U�]w?񿓩�3ѳu��sh�:Z	;���C>�$��%��ݭ&4ʢ$h�R<7�
8r|��V�B�f����b���,,������a�ٽ�N-�<�`�y��뼦u�XO3D
��};��?/wl���+"y���;˻���~������y�L1�}H���� ���eSKx���=�S��7���ˏ@�%��i�M�n����ܛ;_;u
�I�?O��x��!CzW֘j�گCG`΍o����Q���fڞ�;on���k ����3<Km!�OЫ�'� �$i�n�W��Pt���v���~����Wλ���������!�I9�pGM�f����>2 ޮ&���٩;�yx��T�:/[�y�2�nj�G.��]����@��uXȫ3)�s5*��ژ��;��>����Nݗ/]����u��َ�4��N���U}�4�>]�{���}a];�Vk�W����\^<*w��r��~j�(Wi@Y�M1�u�����g���4�ܲHw�|埍DE��������.���`?/����a`ąi�y���F}��ύDe�X>g��r�v�U��r�OՋ�Nip<ݬ�۝x�N�O��˿N����͐�4B������P�e�6����&8^y��{�?s�}lz$拻�z*P<��Cډ�OG���"C��.�x�y}��W֬$z�n�jw������|2<G�υ^�ղ�%y������݌�߁��U����Ҭg��^.�f��>������sI~U�2劌J�y��vaّ{��Ո���Z^�zH�j�E���[z�����ʦj��ǨX�$/�<���_
������N���z�u�o7����I�G�p�禍�mxfz��a��@hu����W΂���=�mt~�o�k{�����yY���"�ܝq��xR�>�ә��;+�1V	z��o?��5;��U%�TG	�V<��V� �Ȕ���՜�f�n��\h��Eٕʦ�5aժ57���躍��ɢ����%�ŃpR�Y���K&�}����S��b(]-���V;d��'���e�f�k��8���Ϣ�0�̺�����u�\ˌؗl�7��_z�:emX�qA���|(�N>T���f�0��BT�%���JKNb���P�X��H����ʊ�e=M�pʴ��YLsrU��`փՆ�p��am����,Tҗ��1m�oz�𸯴��R�Y�3�|�R��zqVli��ltS��]�N�ټ0|W�u��AǬ����wޕV��'&�<G�G;�F\���뢛�<���.�'/�ml��^�õ܂&�$k>�3�sg����jƓ�׽B�!y��F���Zq��ޜKU�8pv���gJçZ��޿�w�c�z��v��	��qӱ.�CXa�s]Z�Uw.B�h��}ⷆ���bJ���GoF�5�u͕�J�e���㲌X�.r�1��X�����y��U�ܽ�]q[j���t����9�flx�������j[a�su��&�v3u�8�ָLX��1Y���)h�r�g,���t�J
L�Rk�k,+� }����kl��0��`ϗk6Įƾmu�q�����D��f�)��u������lW+��1�7��oa���Z�B�Wd�fX��}* t�KOU�i:V��C�vؼ�l [W��ӊrПq���@�L9��m��&����%3��U��Oo��=�ǟ/��fUɓ�2��02{���8ik
��b�Nq&�%R���o&��a���\em��Ltv���)�\��j�.]�8|'(@�r�[���F��NǦ�/�,5t�}]Ȩ��j��`�����s5�}���_db.����7Z�+>|�>��UЙ�}d�l����g��H%�跲�L�YU� aV���i~B!�`Y���ݓ}�B��d�p g���,(��8ͥ�q,�[[ڨ�e�2+�8Eڻ	hL*�y[e�k6T�N�2�����6d鸞��ea� �m�K�`�o)��hqmJ+G���)]�{7�P�r��n{�F+Έ�^n�9tŗ�ƙr�� 0b�U�
f������Z	��]�+U�V����\������,����!)�ј�"~+i�y=��Wy�X���_�A"
A�W81w�<���h��ҽ%w�����5s�FVZ��ˎ�[��Ѭ���R��rޭU����;�$�i@{��o��v�ɪ��˹M��+4s�s %Ht��f`�\;(ϏF�&�&��D���=�Jǔ�����\�f�du�'�?2��wY4��|�S���P���n.��v�7�o��uD��I˩ˢ�[K`����{ɻ=���K8����w�9;1[g�2�nC��p�ݬ�i�+�^��޾>����HѸu*��;����S�!��y�� ��KWh]��B�S����)!L���C�K�r��EQej=$+�'Z�\�ª���h�ED�*��.�(�T<a]̋�\ꙄW(��5�&PjV�Y$�L���*��d\*��E���iét�"��"5*��j�ӗL9΢BnaS�j˪Q˙%y�/Q�$R*ՅSTADʨ�v�BȪ��W"V�g*�"�*�(�\*�"�d��2ʢ�"�T�E�*%Q��^���*�*(�&W"I�"&T�UG��I!�&vr9DEA�r
�"��h�h)�(�D��QUEp��>D��V��T\9Q$,�Ԩ�Ru�"�T\��*(���ED��a �QQGđ{󧄞���.DUd�UL���+�TUAS9QOV�9"�MC1��P��(����ʯ7A
��	R(�Ȋ�!�TJ�.D�t�PG#�%�TDUE�Y!�(���%��(�ǫiT�/V�#�U�r��P��ʵ��j�иm����
ლFAt����*�߷�ޡn�|�i�;٨��S2��s�8���숩��?ﾯ�蝹���^�u�<bI?����H�o@�;�����/6���%Q�W#��L�oX�7g��o�;'+���hl���-l(�z&���!�2��ncw�r��V㉛Ʌ��ׯ/ۃ��M�:�`���w�!ƍ��tW���o��ysRܬ���~��]���0��?Cr��1Й���p*{�R�uǌ42Ȭ���1�<����|��wNX�m*[�Fr�^[�{%�u3%��Ld<5��ε�|��v5�s1�f�&��r3'Nꪋ��>�։�-LA�����ʝw��׏��k���|.���ɻy��Qn=u��CW�	�=�F����l]W�o��K���̧^I��Vh2�7A.���^���ƚ���l<�W���1����=8L�H5��[�zԞ���v�ws�TǖV�S������������-�r������d��ݠ����rD��Q����f�|�(����}�=6m�r���C��y:��n�*4bh�������R����uɐ��9�y�';��.��N.��r�g�nΝ�Ed���{�G\8!���b��i���3:���r��E��Bw�}�}_}J+�$�<��z��C������Oَݲ�y+�i��%���g�7o�y��ֽK͆�xޟ��BT{�2�P�v_�V	�˱���n�4����4U[�ݬw�s6�6�z~ei�=^��P�.���,�A���������-�u���#l��,�u�lꭘeo�ñ��ѻ���>�~&��M�qw���^����F�\�s�ӭg�Q��ɪ���&)�b���a���1��J��$�{���߷�]ֽwMV��C����\��G�^<�n�����}���Me'mfNʣ0�{�_t���g9n�h���V��p�|�:���{���=�R�:5{<*s{��ʾ�]�WСV��ۙ��^�۪ͬ��gŲ6�����C��	�]v:���z�(b �
 [x�;��{����q����g������D*�@F�V�Ϊ�"c>����� Ғ��֌ro.q_c����,�%:�oʺ�L	�}4\�]:���A�V_]l���o/�؁nߩr�lB#'k��>T�A��t4f�˳{�Ն�X��W�s��/����M���g+P��u�pr�7��+�AR�Mv��MG������ml�#����-����lmi�EG��L�}ܨfr{����#�si��#nΙ�޽�s[�OZ��Wz����ᾅ���_=�fHy�;�2@色���$pY}m��G.�hiq�S�Ѫ�WQ����������M�=ޙ��0l���{>�,<����G;����+{<y�ŏ���3��6N������[�h�퉟x7�)<<�e.����N��.�(�"yc��'3���^z��Kv�Ɇ׈�7f_˼5�_P�ï��=�����͡��u��7N���:���t�U��}E�і�A޸��yw�^�qj=�mۉ����:��k��+��uR����/j�
#��^��!��VnQ��l�u��׮��y��y;�ssBP�+KЧ^���p�v�g{�Ű�d�����'2b<�V��/�޻��(�fs˅�����+?xu��WP�A,�%���V��7u��j���W�6�Q��l[��yݘ1%�Yzgz�Q�g2k�@{���X�2����;G��齧-�#�
��{�,�$�#A V��&�ӵw[��[�WchJ�r�I���������㎜��v�^�Z�}�ǩ��Dr'�d�3��ѝ�J���V��t1q{��=4��>�n[�46k~͟��A�/�n�9���@��w�����{m��K{Uly���Js�a����1J1@ۅ���P&&r��M���b�p����{�o�a�nS�f5#���k�2���uC%�i]�U�ཱི�������6}
5�Ru3~˂�7t䍺�t�3_�3��.�6��S�1[�_oS��|����7D�Zd�T➙R�]��~#%\�۩�����yӟ��_M�2�Jn�3OV/v�-��U��Q���]Е��o�h���^{O���#V����5Y�]���r*�=�fb)�7Q������+����r].�d��]a�Y~݈7�zYe��,�OS��	��=�~� �����ً��Cޛ����U��)ֆ%�����("� �c�C.�����Ƴ�iSB�~F%�K3�	D9Ve �$�Q��nץ�^C�y277���ڻ��[�+x�Ւù8b*'x��+��� T�뱏kQH��������C���(��od�-D�i�t���U}�}�E��w{��v~�:�e|�
�~�V	�����_zlϗ�{�!v`?{6�zB�nh��g��.�V�����-�����;/���Y�Y�E�I���	��'�R��(�0�t�}2�V��Ft�9.xSڂr~�e�������Q��������΁�������M��HI���6ϡ�ܺ��M�]�=Y������׵�^�Qhkz歋��w��/7Eb�k��Z���t,׹8q�y�{_����>R��{X����w�R�� n���n�����2¿{}�L�i�[�}�ח������!9ݦh9�߳|�;uX]�3�n�Ǜ�B22���Y��f��-�˸�:��]����r��f�E⸽��Xݍ���)��1F1��m�Cݯ�c��3G�w	��cx�x����n���^�pv���8�ʆc|kmL�U�7��t�oH�誟W���4@�#��wWEY|I�x\�v�;<���`��ng�ʳe'�j:g��r���L��T7���X���I�Zo���kt$W5�Vˊ��yϿ��^�����	�dZ�J����>�(:v�=Po�Cn��#liRMI���%�̟�_}��W��-Y����mA�n��B���-!咮F�_k��o�����z��sO7|?��TM�w\[��0�T=�}��* �n�߼3s�rw��qV�o����>mrc�Y���N�w��h��l�s쓖��{�~Μ5g��D��K><�g��(�e1�kq{[i������u�6��o=�(�d��������>�-n����վ|��&3�����x8������^�~���׻��sa�_q�5\$8t�=��U.����_J�վ�"��-�.�"��{�T�ܭsݏ�h}�j�{^)ex!��z/TkkK��j��H*���Bzj̭�ڃ��U=;������g�����#f�+��Ke���yy�������)׮�Ǖ����/!ց��c�BE<�<V��j�~>��&�5s	^j�s[�v��f���Z�,�����r}9��E��v�a�n!�qe��"�^��O�ݪ�z�ī<�Tе`�xΓ��r���,?l�Vuu�+^Jۀj�/��f՗��̚a/�@{q�3�BH�*��zeWi�[vdYN��x�H���
Ps ]}.���gG��'D;���#�o�r��ײ�
�-����~�G1�9��{�����y@�%G�_-�ξ���/rs������t�(�_?�x+��sݟ�}}��c/c�#�̓�9\�s�ƶnal��s[������d=���m�{+��5闫:���?w$�/V�~��	����t�Ƥva쇾��O�o0������-Qm9��{sw��3lmi�����,{����7*�u�����u��t����lz��Y��K�ƢF�X7�k�t7Э���f��3-=�,z��uX�N�zyg�@\�UQ�G*�yG��}7���?C�궶��罠��yWG9e:�g��mɿ �&����tW���s%x��M���M��q��н�x�����M�,9���iZ�+��~7�c����j큾���t*���n��s�^{�n�{����24%G�r���OU���7���@Q��Rg%�[B���m?��/2��U���\���!BL��'��h�JW$X*T�obHc����c��@�ge�X:Mޗ}!`�9�F9h����,��V�'J^B������ƏD�a�ެ�7]a�5q����UW�}��E�r`���_�jʁ���~m���=�����u�bzCZKy~��"q�-��NXݭU[x�nMEy��^pbݸ���Z����k����F׆9 �Sr�ӭ,� y=Ƕ7E��]1I�l��w^�.u�^b���/[�Nhq����t�����u�Fk�/oFwo��������2g ����$�J��Ǖ[��k���-�NǢ����'���̭���2�����y=���������O�庋46b�������+��"sW������#=[=��7B�z�U�=��jӝ2����1x6�m�5����M�^����Yt���ws�m	��n~NY��H���[1���z�Vm��y�E���F��^T��av7E1�To��%�W��R����K��C+]��,�|8�OY����.�7{Ɠ��	Y���=W���gd��6�Z8�û]z(��I������|k��錹�v2�-Ԟ���Ҽ�7үc��Wi�3u?d1GT�C̹��6@��wd=3�M�v�!�;;Z�Z��{7T�hɶtp�:䤥����ş�[�I����]��x:
V��k5� ���+�������[�غs�=�_�Ք~��r�7�~ ������ڗ��Q�-ˌ��x�8l��s���qy�n�5S������vߦ�~߃K>���i�ݎDn�x���`f\�wX7!��������kW0�T��<K�<�ۥ�yLLI�t��f׏��.�Ϛf�~Ϡ��=O�K��my��y-�r-��n��o'�vt�r����<>�Ŏ���V���e	����>qzl�^I�zג��O�Vu=Nu�c�DK�;faR��yq��n�&n�hvy:O��d����P=�sfsL�)�j���}�x�fU��T����^+�ȕ���������{�rg�:E^Lk~Y_:�6cUl���F�alf�xH�։oQ|�����d��{�=�z���:�,��o@ٍ[
,����,���5?j�g�)ݼ��1v�w-�v�;�ۭ^n�������k~���~ �A��a8�v��
y7+z3�\����ij�e�N����.�����Y���^�B�C��U���q�soc ����{V�j���[JW��Sԧ���k&.��kp6�Slȸ�{\�ˬ�9X�m5}�2�,s���;�,�bZ�4�S=��W��U}�Ћx�;��聯��4�nO�^{7����O���3A�V�n�U
q�r�vW�N<�T@˄+Y���t��Yw07�պ�Sc�1�^^����)m�]��6���ݕ��sT7��tz���u��U�m-�έ3C^%��㚿��q%�#K>��nW�� ���K^}ổ�"呻~�MT8�yx��"��xiqn�O�CtƔ׎ �@/*��yd>�tǗy=@�vޝ^/�N~�Fo7���|5z~x*�fb�yPJ�-���nEl���>~���,�s����Vk����U���YT�[��g׷<�N�"�>����N�1,��O���ë�����ʇ�^;�g��*�������3Z�/ 7<�u��RyG��|��ϕA����u�^/?͌}�ed�����{���[��a��zk��*������+ll|%kf�u�O���cr�mPR�Y�!��|D��]�ms���<��fI�^�^�a�hAl�ī�5i��)�m�!{�N���P�)b3�iɜf۱�i�d�f�m9�|ƻ�.w:4q�#���eb�*��`vb�i=7��.��8����O�[�-,r��c޵s�@T�9��5c5qΦ_ci܌C��-���o�T��1��5�z=�UDP٭>՘.�;f�4d�Y�KY�ﯽݧg	�tQ�m4g��t�wԅ_y�9�;RY�:��d�½Z&���F�S-
���K��f��{m�N���w�n�_���
�^��|>M� fm<���F��Z!�](ZU�7oJ�.��+$pN&qMc:��7�,�[K�׽�,��嗢�㳗�]N���n��2���m87M��m�o0�B��pa �k��ʂ���F�[��X� a��V���:� ���O��15�}�����r����N� �aAB��5u��֙�%u{��w�Y댸�⣊RvҮ��e��V_�ekrvܥ7*������Kܞ
���=�}A~ 9H:?N3Ds���z���c�Yr��u�_,j�{�,�R9��tu����"���Z2n����"m�=�C��:!^Yˢ��ga��¬�����L{v�#�ަ�a�RS��m�7��3��L�Rb��ІK�iTc3M�Ξ�u0S✰�0���K�p�̢mrenV$\@�y�c����i�1��lS����{��M�OA�{&���r�+,.�:s:�;��+��K�{�~vO'+Ԫw]�P?�����d͜��F�VeY�����-+^q.��B�|�V*Uy2s-�к�9<��=|n�7���� ���흛2��=L=�m>�mݐE3��J��8�lE���Wp{��<9M���z�W�
�_T=��ٞqe^�r-�c�3��S;�	�ێ��[괹*�MDl\Ioa�jP��E�%�F�7�B����f��C�bm�ȝ�f��؛����6���`�
M>�M��ݡZ�^F����� �=��Y-�%�{xF�M_&��ԗ������V����2�B��J��[:d���+Jvdܴ��%&�y��*���u�#�h�8n/@�� �m�ƺ-�W&�8����_v.h���8�.!�<��0���_$��Dp*a�5���rr�h�Ἰt�J��*�.�5ң������[�-�7���3LP��9�����l:^�ݲxb��0����!7μ3� ���%�C�����yU�y��ē.nnq��(X;8g:F�]�"����|ɾk��,�\�ё)��v� ɺ��cM�o�f����-��%�ݦ���C�۽Vs]}_<2 ��ɾݕw�����(�q�jܸ�1�]�c��kD����b�/*��.�J�R�pG/�.n-m0�j+���ךċ��x^�G6��e�C��|���a���Dg,����9�Ur�h�K�$�siȨ#2�����r�'9s��fU���xeR�$\��2�Q�J��p�E|�r���4J���dQE�ӽ��Ts�$��B**#�#0����"(�YUs!*��P�QL�" ����
�9W*�0���*���F�*��"�
��DG�t��E�	m"�"
��.|t*���n�ܪ.UI"���r��Tr�
�E�\��AUU\"�"ng
N�3�B�LQL*(��H���r#$�r.��fvAsVfQS4C��
1H���]�TG"5
ft���\�PWxʠ������L:�
+��.r���e�sʇ��o\��Gs
e�*�u	�DL�ȣ�Њ�e�(�**"" ���"�@6޻v��{Ӷᬬ<@]�[�fH�;��R��k�n�m>�=�� ��6Z�˾]�g��n��m��6�?}�}��~UxN�;Ǵ3���;~u鸽�<�D����x���x�|Q�G��N���)N͏cW�Ec���y�̬y�S�_��|�,�ZΪ�eo��jQ��^7d��Ũ�jS��O|v��:e/V�pU]�Xx�5z�۞-΁�.��B��Y7�~��+"Em8�-�_I͟9Q[�g}�޽~ߚ�cE�U_�񙘯S�sU�~�n��.�U�8?������oy�֪��/�n;�}m��\5N�㺭:��6�.����/O���;�W���ߞ"�H�����sk{�{��+����٦[A�V��b�bp�m�{yQ��Tf���v�z��2�?y}���{�u����G���u���{M�%�S���룇Ü�jD���}{�j��I�}�|ï���b`�3'�>�]���D�������1໖mo%��Q[�X�ާ��F��(A8{��{���iU���6t�S�ٗd��
c������"�I����VE�@䥊�7Y+�1Pen��^�\R��3ίiEؾ���g<�8=�����wɌ���W;K�`vBz�(�*�Y���R�. S��w�z�r3޾��+��U��}�ѳ�p��3�)d�hm�ī��߼uҿ��^S��Q7�����[�Ff�k�|vs\��U�ب_7D�ݠ�%{*D����_��s��p���tZ���e뫩�^ۭz)B/2t�C�s}�yD?=�2�߂���̨�,s����gsw|3�2��v��i��wV�T��ݪ�?W�+j߳�7�g�=A>o�q�k�RP��-�����g�����E��9�{^)L�U����'��2�����֭�p�|�=�V����ͭR�~ש��~�{ffߵ#q��;�KS�2�x*�ɈN7'��=[����Eμ1�v\u;������^��{����Bo�ޱϔ�u�f�����w]_���sb���f���ﲷEI^x�n��;6��<��ԫu�z�#��M�;����B�ٸ���^�[M�o��fo�Ѹ��N�n���߳r�A�(���K8�)m�/V�]�qw���9/��|����˭�$*HFIs4ާ4�Ξl���3�VF�ԁ�8���󉺉��Ed�³�:�z�̾Л!�[Q��nmv����ґ�[c�5���Nn��-釫bb+�+��3�r�ܲ�JV���&��J�@��K��;���}�W�W���۝X�r�:&o�5��f=�5iΙ���oٳ�7��Ѡ}XYz׽�2/.j}������f�'�ٲ�:I��-��A��+�^��K�u�ft�ë��j�4���;���x*ػ�e^^O��l�k�ۜ���d2hWȬ���z�u���gxr�ץ��/��0M\N���UG���Q�&f�S��Q%����99^�*>W;�n�/'x�71܊.7r�mź���
��M=��~�������_���W�N�;��m=�K��\����[�5��^�sEL����x7�d�ۯbUI��^��l�ꢝ��]��_���Ϥ�?m/	�z��ݠn��15M�l~�\����m��?*^�����)��ؓ�Ͳ�y�<���Sko:�~:;.J�wf��^V�4)@��0�zV�����*-�����q���꧵�;�..�4k�ޛѬ[J*[�׼����SjJ�Q,�z;��O2�OM��� 7r�y@emb(��XC��z��ޡR�ʄغt�Ne������.�F�Ѯu�!���n!�:!��ԋ;+ud�b��>G?}�}U_R���Ӄ}3Fk�_�f}^|�߻U���K+��ϊ0utuH�b�u{��ɍ�y�t�����=z5n��y:ߖ9�7#Ul�)�����m�Ǭ+�� ��-/[�:�rlۻ�Y�����'�Y�yhl��l�ر}��>���P�U�/�����d[Xdߺo�Vެk�.�
�2��~��-���R]k'yb�$=�J���ʫMa����O�����\W�������;z!.z����w�w��j������:��1*���y^����-\�p�eI���̖���۔c�*m�r��^ls'�/3}�/[���pGmz�~��$�fN�d���b
�[jg\G��no�n�^~]9]ź<�;���~�*�������C�	X���QѰ�k<���v-���|�)���~�ޱ�ާ��W����Şc��f���$��į�q;x���0�﷖ّ�lQ����ʄ_T����ۣ�3��7�[�A�(�������Y��mƑ����9)X�0Զ���jQ��/S���؅a��S!P]��Y��p��IE'U��v�_�l����}�}�}�Gbv�{|��.OԺ�:������V�����z�:�+yꏫ����
N�l�7ĵ���~ߌHy^���?#��ۏԺ!�y� kN=��Io��%�{/ke�&z�?�~ғ�>V�R��ϳ�9]Oy=�H�݊��Y�?Q9��<^��}��k�E�u?�Eg�7/�kMÊ��܀��CC���u��=�y��d�;�����Ẽ(�kz�����8�.�ի��?)A��	ӧóɪ����Fo����v$��LK�5,:�x���F��.�؋����t���;�^�nQt襄Q�5(�OM��i޽3`[��p��9inm}sg�kwM����^�#5&�H�|��Kڧv���m̭����S��[��I�̝�b��)Yez�&�y�U����2\Я?����-՚b��يY�
��C{~��{%�7�FV��H$ǻR�./row�d~��n�ܑ$��e�oa��y�to^���c�~�����s:nt$m�W4r-�g_n� ��o5Y��H�.�}
X-�HK���`ͭP�W�/�d���(f7�ݎ�b]�s3�ꪯ���{y�1�e^�C�7)Ι��s�=����նiN�J�Z���f�M���}��)�����lz����}���׌e8�w�5�sQim���/|f������Q��m}��:�O�F�bN�.��ޡ�Ռ�o� �߷�iW;ԆL�Ak�qo%��?��X�ާ��J����=I�����N��o٫Í�jb��_�`sKh���\�9��*���v�{�\њ뇓N�,^�]�yIB��+{ꔻa�vߦ��T�a�����t��]�a24��U߼��y�&v7.4֦}z��ϒ��@=�2���h�yG��AR��a~sY�;x��^�B}Py\�^���my���qU{���5�3�X��εwe��vi�8ܖ�����v�0�����n|��v�^H����]~:�>7Z�=�A{u���ӎ�h�V^�K�S��J�:v�q�&���t�g�[���_;�/��*�6�"[��:�lYT��{����_c�ơ6Q�s]����ޛUm��U]��L^�fٶ[��o=����]V�%`w\u�E�(�dr���;JU�l�}��K��Z�/FaE�,�ծ� �d���1�Y��ߪ�����Nzu��	��'�Rϼ-"�alnO������fcu�s�^RN���*�{�|�����xۣ��@ٍU�����N7^�W�Q�R��{�'ss��ݰh��v�^��k������i0�m�(�=���!�)ٓ�3/N�<�F�w/�}1庋46b���khߝ�v��V�u
�Ƚf%�{�N;�3�+<��UF`��>-i�6���߳H�!l׍5v��V������hE��S�?w1S���0�c�g�9e��ޞ��Puғ�k9=<��U��C���0�����w1�����5�`�ϴ��d^zU{v�r�!�m30ua�8�ʆg&��.�6��i;��Dyk]t������Y�rq�C�0�[��?F�QX驃��6�.���9S�jT�� �n�6�o����Q/�g5ź�^
���J��A�J�J9v/7E�(�i��ٶ�V�C��ݶ�M{i��)h�d���:n�ׄu�ևen.,��O���˩@�.���roT��L�����u�Wr�g19M@�v���˷����
����ҳZ���k;miRwMwl�/�ef���}_}_S��M�Ow5����_Zz�<���W���ֵs�=3<J��F�]d*����hwE'	o3yoԺ���=���s�>YRz��x�M�מ�ZVZ��G���.3�{R��xx�-z�8t�޽K�o�K}LO/m{��K`j^��z�zAKb�<��tK��V���ןt�=^��ն[��K��d�f]�;r���2ٚ�^���M�W��u}�x�Fe��zW�����#y�;?v�yf��}�h췞�y1��e:�6cUl��~���<�_�ANFg���9�~����}~�觺w�]�'�j!�c�#o���ձ�����,�Xz ����|G���u�r�}��[�����q^�C</z���K��o-�����<�/���|�k��ӊ�{��t���˂�.���{j�P�Ἳ��㏬й�f�ԣ���۟�[���_/ �oه���to\�%*0��3����|U�E}�=�lVg����B;g��zq�E���t��b��&4IF�u�em�:�Z�"����ɠ.�6�@5.�C�L5��R��N!{`��^�	�g<��]����ڃ�>�W�n�N�	ݻ��f%v�UU�U)�~��ynk<;[6u3�l����|6�3����\���i�����z��{���;�֟0��,�,�8��D3��~��Au�>T=�|�wtf�:��ѫ|��3lmDiqn�����Z�8�˰���9`����-Ⱥ��m����˪s��W���uź�j��	�3��|���y����ț=�
���1x�.F��~�_W�oz��w���)s��^|0���<�����v_s�i�b�O�����n/D��otK������kj����W-��������3�ۺ)<>V��P��>�'� �m]�l���o���^��/My��[�$~7����j+t��j��Len{���G]�����^=��w�9_mxm�^���գ���4�����|wc�\狥3��y���g囚5:�;����e}��k�G��
��.e�R����]_jj���-�:�9�ztzSV~\��so�|}e u���{�߮v�o��^|�O��{_Pj����@n>Gu��en0�I;oS���>y�m�|h]�
����x'#N�Q��zឹ�ps}F��ѷ��n���kFm��������;�^�x�z��X��8�s�{�G��87�]���T��.sГͨ�����w�]��=�T'eaV�y5����Vh9���5��Y}t�E��̝�f�~�
�mG�#(Iܬݱ��p����N�nć;�웍�k�W��.s��f�a'm��}�;t?QNLw����ܧ:e��[����mĭ~�,�b�"��ƨ���+xz�<����zb��lz���$�f~Ԏ�A��J�Q�V���q��'l��u�L�f;Z|í>�r�ѩ�V�HL�Ʌ5�q��G��3�@~�f��+��w��5Ű�1�5�f�D�����G�ֺ��ʞ�U	��h�C����~G;�o��%�TϘ�G���{�G�36�C��qP�I�{A��Tv�����m\�OB)�HQ��e�)t�iǨ�[�����25{c���L��������%D>�R����Abᚎ�K���׷u���J!#�j��,)��[M典v���e����R��u~�7th�L�}���-A�a�S�nL�܅�O��j��l�ԡu8a#��jk3 cn�ҧN��/k|m�p�Y �w�y�	w%&�kw�J�.��`�]�.����̍[c	C��[Cr��!R�Xz�����;NT�#~|��ʔnf�\��u�O��ռ�MN�F/�����V��1���dq;n�eM��r]�fw�ΡJJR�\��K����}���w�D�)�����:�+벉�V۲��4V:;2��l�}8�G���|���-��ɗK]����k���]�B��͌%�h��iX{�Y��7^�qՐ������!b���$Z�jX���뮆0]�=i���E������-F�e��WQ����^঍��2�����*�^�:�ŝ����Ϸ��=�6	��@�����q�HX���!�2���Ӯ�j�=5�]�$��%�� ��3{��6O�+y2�_Y�C�X"�y��y�u��ϱ=on�Lhl˹x�y��˃���́7���_�R�v)�\\vjurw���\�_��:����h��.��<�!o+��$[4{Ǣ���굸�*l�7��d�N�.��]1C�썥|u��5뻎V�����:	Zi�\�S�u�LR��m�V�v�-�wZ�KP�i����V ��b��(���^N�^��2�Oۻ������!7ms�x/rы�jѐt�I��o�u���ǋ����bW�ݣt ����3k�ڎ��5<Qn�����j�4�:��w��pr�b#��q��mgb4��Q3�qz�a��Kb�q=��_PifH�rf:{�v�����ً#�̛�B:�4���t��0�O�P9�f�
|��%uq��P���}Z}���w�QE.��WlMj�����7���Xy��+�hFo�M��U۹_��*���=�ځګáJa�1`���t�vp�B��ޘ�{��a�-� �N��z���'[�P]ޯ�#��NC9f� $��>N�_q����;� 4�˽*���S��ݍ��i�B��_uZ-$�tJ�����{�#���]�:���BOE���⮁�u?���3�{؅�#�[��[)�u8v'sGx��\[�wo�|��F!�9\q�ݦ���1�qc;C��=��P՝�'K�6�
MX#eF�鋅]1�Uɧi�KH�|����b�3�5{5qv\�/5�bA����*
����|�K����2v8��Gp�Z��p`�%7CT��l|9[��5�od��P|�]]�V����9umVt�uK����NH7��v��,].�s�e"���z]	��v�t���~z��39J�*%�)�	+(�#�l�
�������(�QUPr+��*T��yFQE�Ե���TUr��Ȁ�吚�i���DTE�2
�(�
���TTPt���TA��9r�Z"�DW)�AA%ʋ�"���Qp���8C�r+�t�ATvQ�AL�ȳ�J�AAr���
���9.T]P�Us�*��r(�ʸ�AW"" �U�G��\�VʎFHP�	*�<�DDE`�r��3
"�9˺�DDDW"�8^aDQA��\�B`f��DEUQ� �Q�3(�J�
����2G2+�2��*.E��Ȼu��E(��b�EUW�r�DE��*�S+���!�¨���숫�p��<�����ݹUUPQE���+��DN�˚ _�r�bB�
�0�z�Ǔn�X��5.LS@5|��t�ZE�p����zl�{`y�˱�����:z�P���_W���#6o{�l�CY�cL��7������tC�x�V�L-I�s�F�$�F-����X�Z�+x��~ߟ���=y�%�^��k���V6�0�|,�~���J�C��Ŏ�7�"���{7Λ�y��Ly���d�ĄG��:�M�]:-g��K*�|	|zL{cG������ͭR�{/d]�	>��:���sL{[�7ڮ{x���|��K������5;�L��wǳL|�zo�OENK���y�������;`v�6��������`���n?v�����2wPױ��hl��=;�z��^t&��ޥ�=��ȸ��v�s�3xuTy���p;~�W�[�46k~�gb��~~��cś�]�+���z���q���Y�����7��S�-��)����6�K/=GWOq?E�F��qѫ��S��qt�ws�m	m��$,��^f��Rz_,߯������!�
�Ok�FIZ霡8�2a���Y��Mx����]�����L��	��]�6%�U���׾Mr�Zl�^�Md���JV�c�-�.�Бu��{j��L�fZ ����5�;��*�f�fI����Y��D��3롎���$�Cr�x�F᣼�_�3U�^n��z�EPi;Q�X��[>��24�0����A�眝����`�X�.���pk����!�c��K�q���A�A*��LA�i�&2�7���Wu��'�|�}�����s\y��S�T({D�� m�u�(5u���el�S��27���鶽1V�Mjg���r�T�<�&�z6�����W�0G �GfO"lv^��),>V��x�/��<�OS�י�^z���{w�5�幣tί9�k^^@%�x�?pl�	|{ֳ��7ϳ�V	����]X�<�<�������~�ݱ{u�yZ[�{^|Tz�R�����hu��.Yݯ�v��v�U��{~�&��2��	�]��mx����+�&!lnzrS���ߓn�{�fͻ���f<ѩ���؍o�*h1w����W����S�`N9���͌�Bj���U�`���=i��֚"#�^Ftr���.\��ۘ4CL������>�#p�1�<���ݵ�yn�
:�r��ý���N��l��~j���øg^�Mvl����k}�uur��.���U�}������y��3��ܟ��En��=w��y^�V9�{�
��k�A�/���v�za��/-!���;k�S��ms�.O��J���B���{OێT�r��>}���X}y��B�y�d�3���]-{"�yr7�^����)f�'�U�϶�f����+MJ��O�\盞���͔4�������w�����o���	�2u��=���!�TA��?�&O�O��,�m����cw�@o�Wc<1Ɵ1-��.����8��3��U�e=��M�y��7{�6�9w^ўef;Q�ź�>��<r~L�މ���B�5�����*����n��+}�;��EM�uǜi�x% �
�eǮ�-�q�lZώ��_��K(���\�9��VV�����[	WG�q�9G��Y�J���v_��/J1,<�.�s��-�[L�¬w��}0��W��E�R��mx���ב�V�t�Δ��ļ�/9�g�|���>��~N��}�xJie��m��	���.�])��U�ZL�����:�Hs�*r�[~4����y9	(��[	Ȳ��gL�����fO�}_}[48���K�Y��p�����w�v�3��n�/z�?O��c*�fA��S���='�m��C�����ރ��MyK�o��I׍�\�+v�֯D�^=Z8zQ���.9-z������19{kݾqU{�g�!;6�:�I��֍S7r���^^�{�N>�<^^�K��S��3�oóɪ����1k���x���=��x��oʶYO�N������wL���P^<��~9��R��2��e��z�f��C�f5l(�7�����I��I͟��En�Z��ns
u��6w�gS�oE"��ۨj�ؑ�[�l���މ�{}?#��"g6��;�i�fg��YO77�\{׎���󟟰�u�uf����6id(p�V3��t���&�7v�N=�;n���~�������Nt�͠�~{�Q������HĴ���߼R�U�����Oޟ���~�o�~m�O��3������[M��}:�E�����U����Nz�a��w�X�FX2�A?;x��IZ��ṛ��9Iy��4h7��}��"�@x���{o!ӛ��r\��f-�U�e%�@ea�jf�� I���7Θ���d]L:@f�׹}�Iy;�����N��磌����t�43z<a���[f~�^~�+1�ڍ>a�i�I0̛&�;�ZUϢ����C���/����^�6���z��Ao�Sy��	�뇲�d�
Jy��ܤ���Cbal�1�����t�j��W�����M�bT��s6�Qq�η�>z�1n*�(����'�s=�[�{��Q�>�>�n�����	�N?��됵6���|���|MzJ�ߘz������׵�����GU�]��_��ړ��O��y���s�PJ�v�-d6n�r䜍�}�3�t�>��^����c�LA��n��ٹ�hj���^Od�/Ҽ�5���.���� ��L�]P�.����\���c=r!w��$�v����~tn��1��2�ԍa���`�D��Kۙ�v)��^<�h���Qμ�j��ߎ�:�6uV͕��k%'��MO-�=�~zR&c�����K���z����Ѳ�Ԡx�ݵ�u��;�ͥPEM��ڻH�\��o}��gA�!��.3ˌ#z�{�ˈ�2R��A�O����kcH�*��s�4.�cѴ�y�j��N�Gs��ہ�Vw��ۊ��t��nUf3?o�w_7�٬yhl�zӱ��}�.^�����3�S�'ު�+n�wN/=���������uhl���gxmlN⦖>A#�t"|�z�<"sڙzsѮ�>�s�o���s��ڍQ��ЫV:�*i�-i���_{�MC������<�qvQ�r�����<������M���W�tB�fa�vcvGmx�F��׽�,u߱��M����Swo��(=b�kgоn����f ��,�g�=9ޤu�c�D�31U�loܮϾZA�9�kK�t7ѮV:jN �W06�tKs�����ƪ�u���+�~�ٌ�TM�g5Ǟ@�R�T'�J�{A�Gbp��w��MC��=�i\�S�(�c�Z�Zr�Y�g�EJ�����WW��vgIt�����>V�w�/��UI�~گ3㽠��=���=/��o�Š� �����&�5�32OP�b �&��q���u�j�9�;}X�E��.�i�-t1>�۴!�o�^����dP_E��=o���o6�޴�c���"V堜Ԏ����=�m{C����"�}U_V���MN>X�[#�������1:Q[���{:��F�]F��-Ǧ��I���v�{�o=��[�yZ[^7���e+W�U.��=ʉ� ϱ�m/�Ș:���&���ϴIگ����U|Q����~{�x�#�˸�%ꅵ)}�~t���>�ߖ9�7L�`�m��Uv��t�ʮ��u�O��͘�̘�[�g|��z�Z�;4|���!G�2��f�'���t?-��3y���m�'6c�*��]�o>[�׌z�cO���g[���s�����Z�VoD���a�Q3�+%}�י��(^u���gn�pM��=���+�9�o8�k������8���_W�;�;������ⵞ���=�y����Br��7�~{1F1@�"��蝱2�{B7ق�n�c�뱯������L6�$�f`�f~8��C1�)�i*�Z�}G���P��.v̲ļ��ۥ�#�R�����HWUmo.t�4}in��Jn.
<L��؝wpw�U��+���X�k�)e���q�yg���V'ZX{���!��NT:�<d��sDn�����Q[�çX)��|n�����}�D|�W�4,��"��S-׃�����֗�Ty�buKN�%DEZ����o}9g���_0h.���T�[9h��`����ؖxO��C���婼�v��;#2�	V���|Ӿ�V�<�^#N�B�y̩��	�gAj�N��p��㊙����{PMۥ���.�s��`�[y&���o��9΅V�ǵô�T?��Ϋ�����Q�항��.��P�Sյ�ýe�W�����,�W�'����_zk�^K}�N��E�uj���sM�9'�z�_�귊P�;~}LN^�g��^���M��_9�.���h]"U'�;��~�
!���Q�����t�9��`^���K�k�5�����s�d3�-�ϼwX;DNZ�͘�y>�5��u�~5s-��u�X���V涽�yE�δ�[/k���};pN^4_w�Wb#��Ԯ�r{�l��Ӷd��apʶ�7���:�ns���v�_X\p[�$#F�B(�z+�cg}n��_d^�ԡf�"�W3�b�l���h;��Rɝa��pxE1Oz^�<������y,���[?�����jw�{�9~9���wP�k�46kp���oD{h��2�ze7��Q.}�'}:·��&��ҷ5��py��N�n�,�s�f�F���_J�^�w�;-&�p���Uӹ�ݕ�r5ߪ7]�����Nt�͠���1���R�xly�hE�\1O�5��Q���1gm�D3~�@r͓.0)Mh;���Szy�u�����P�󨯏�x<ﶸ/_�-���Ղ�����v>ۙ^���9�:��x�uC�E�c}/�1��R1c4�x�3���^��\�裶���~T}/(����	��v�斞�8�o%�ÝgM}�V�o{�X^��EDۍ3��s�����T/�Q+�T��"XpKDo�%#�g���9�Q��=ng�����%w�?uܕ�}���c�e�z��Y��Y�������/x�� �y'���������g��}��"~���ʸG��uff,��k�+��aֻ4�L��Q:�#�-�Hk;6���O/3����5�E�I=�ӎ�]Y~���u�볥���a�f���㘊c>ػ��_'֌+*4�gR.�c�K�¶t}�ܔ/�l;���' �ﾈ��n��]��n�Ц2׾T�[q��;s��$����Ӽ��K�z��1������N<g��3�����,��xg��z�1uB����G�W�|-���%�E�y�=Urk�w���f���)eW���utt���c#�]��Е7���R�/�o]As�=�'�߇m{zﳎ�ڈ�-���\��-^�&^���ٛ[��+�=����g|˺o]�X�$n��9ձ�b�Ǫ�@���)4��T� ��G���fN�/wF��_��k��H�U���{4fj����j���W��쯶�y8_i��μ�m�L���P5��3����d�x��
��G;����B����J26�V�03nb��]����/:��gB����r��b�w��f5#��C��_ �ِ�LW��fH5��n����e��/�U�z�|}	�dig�Cr���
�>�����IO\"g�w3Kx�=��tV��6��I��91b�m��qJG�mh����)N�f��}��;jo�o��է�ނ��T,K�x����_�J>
�s��z;4z�6.�sB�("}x55�3�sQ撚��`�h� �/L�mZ��/�<8�=�=��|�c���,˱V���Ѱ���qFi���`~X8_T|�ޮW�"+��}vK��Ǎa���/�#|��N�fX�F;1.["�^��Ș7����G�L�x�ٴ�.0�MJ�:2V9@e��Uº��<Z�}�����Nz�Y�`�.�[����er��v�ũox�$�S���J��**�a��'�՘N�	ل��K�T��2�K�6�vՁ�vIW�^�n��(I��lR'jZ;F3,s�ٹ�.���������kF���C�V�x�@��+u�I:p�����LP��*uY�v�)Ǔ��y�2`AP�*WrJo5 9� {)JS��h*�1�0z���&�q{oE�j[�r��[(Q�yJ�75��=�L���z���V���bN��)��������s�;Z�9�4�u�ʽ���F���咃<���_nN���/Uu�5r248,�sx��B���}��9�v��ZP陸�a�r����u�����|�[�#:q���8��Q=Vw�cf��+�]{���=6osli΢�,Wz�Â�}��U�o]�|��x�䜡�̓ZTMǊ�����ݬX_c(�]�c�L�vC5I��	��������do�N�7lkL�eZ�������&�\�DVS2r�PnR�cE�ЎZ�D
|ˁ]���x�F��U�(S��亖SW2+\������l���-e�
ؑ���Pa��4��� ��8rz�2ż��:+�;.ȷɗ�=5�X ���t�v��k�� �;'���)p�%���rvs���Y7��m����C���h�<m��<��o��1�M���4�5fp�edn�+����>Q:���ś�|���lk#�zJ�c�ٳش<�S����׶��c9�V(���{�*Ju����Er������v�S���^vT����5p�TWP|c���`�kz���i��Nѷn`��7�͕���Rt�'�osb�;�I/�Ƶ=�� ;�ײ�z��ӭS	T����[1,��bû oNt࢜�`z@=��)^��9۬�lmv
[HP,M(�ZY��7k�vo��Sr���4f��wL����{�/$kts�vM�gLatl���^��ڮ�vJ���]j����k"z����W�<�Z���C�=��Y�wR$K�,�8ڼ�L���w]��3^T�ބ�Ao �7�r��G����s��n�����nnJ�����^��Y��26&�7����f���d���^]:IWgv���N��6�%�J\[��%)�¹�Tێ��	=�w�~�*?��K�\9Ȣ�Թ�*G9L(��3�T���"����9���(�'	�iAW
�DADE*^Xz��QS�ʠ�=[�iDEd�*�Q\��y�h��	,��g&Q	%r��T�p�ΕフEQ�We�S�J�eE@\��Uv�|�!��"x��$�������UAQ4���"�Be�<IU:���>D�\��P��5"��d��S(y�%t�!#�;���G*�+ ��WIUI���]����U^��)��\��*�¢�OX�BpH堄Prs/�8D�TjA+B�q�I�AEUU\��Y��Ku�Р�h�t�D�y��U��λ �XU$W>R�愄E("��D$�0�*�9���!Q����)(�*ey��� ��9�lg\gg<�V���`
�h�4[�ҵ\���kW[o3�"F���B<n�jæ�Z���EI�H�<�f�RZ����y2(���Զ�~��*������-q0�1�Rq��`�'A���A�8d~ރg��D��7��Foa��3\[�3炡�q�
����ܾ=9g�]ouQ��_"�vWͯM[�3����Ս7>�t��E��gg���o}�@v؝m�n���.����q�"�k���E�R���kj������y-�� ��g>:V��՞]am{{�=��{|�Ú��x��Lqy+���6l�c�XU+�l&GjS5R}�mwO���9)��<@����������Bu</-�xh�~����;��غ⥙�鸞�����U�ލ���6����!�_T ��:�T�k�&�wm�Y�)�]N�w�$�^�A&D>���r�ѷ-�.����tJ^f���޴F�Ⱦ���P�y�ۉ�c��t���a·���x�Cr�V���M�=���N�r�p&1c��IN�'���Ihw�Eǹ6m�#�O�g�@������z�j�UjY{p�nK��r��W�����Xp���=�)\��w��_���y��!�o�=z�1�R�O�6b�Y{���)j�k7MdsZ0�u�"it��޺T�K���X�,�T4�����M�^-aR��r��O�ﾥ ��ϸO<������U����z���QҘ1��~9�����U-j�3�"���\�J�����yY�c�ϙ��F˨�t����/��x5p����v�d��
�׋:�z��g�f��6�6��}7Y�+��=gͮ�j:��b�(�gy��x�?�;W��/=�yx��U�췳��
�}��N���>���5�wTd��
�S��ْ�X.aU�I��|��0t�BW�i�::���O��P����_�\s���3�g�ϋfg
�̺��5�78�t�:Q/BS8ą�O�ף���&/��R��c�T7\�{��-K�۝�S�΍c��SJ�5@��$�gzM٩.�I�.�����K�B�eF�i�����=<�ۮ@9QΤ]}�#ƪ#�m'���~G'zvlZ.����<�2X���z��^���[f+��8ϡ��	�w�e}���G�r��D~�#f?����7��cv���Z~�ݽ����ŀ(�eG=�n�gҸ�omx`�����vN#�|���NW�L߬�������5n�5��[R�˖�ڳ���\;V���d�X=��;��i]c�C���r�ݳ� ���SwlR���O�V�m(7��eg}i��p�th�D�����,���P�t�e��:5G�iO�-��}���W�֏k2?O)f����s�(�9�D�c�e�/Ds^���k�k��~Z]VnB��U���'c;o7L�&�L]��=Q573���;j�1n@X�qU���}f�Y��\�76]��?\�۽��n�?w��Y���3Q�]E�kM�p5�'���6#�6W��,�]�\���g�E:G�OgF����^G��,[I�a�Q~�������FÙ���SKmn^�f��m��i��F�J�|�;=�)�=�+��^{$\������c$�*\<��>����j�43S��}�r�z�����W_|���w��O�8@k��Mo�A�w�馧��^��޲�
���9Q�C��ܜ��|��]}P���:�]�O^���-sYa�Uw��p��DY�8Iܐ$�n����Z�x����Y5�8¨P6�L�&�}�=�o�^�B�̫Uʉ�l��l�+��U �|j#�9���wy`,FC������g�E��͚x,���\	j�(��%��rT6�l��]}����|8�8L���A��1���ʒ\]N)���6}O6�ezf��E�<�[%�,��3�;篨���P���	MU3wm_�(<#g�!�i�i���H������C��H1b>�z�9�AC픯I�;��w)��»z���֓�sBs90���u����u�� l�g��5��I׸��~�;��(��{��|����z|:I�G��P��e���bz����<�nL3>�
r��rG�51��s(��tKF���W��E�gH�c�ґ�~�;}��_iY�@�w��]�f��{ُݬ�Xr��ؘ���+]E}��*�U�c�g9�ׇ�;nR<bw�:ǎ;�9�丅�K�czn}����v��s�Ɩ���g/Fr��W��^~���N܇�9�������׭+�T<��D��f�I|N�\��d��q���X�)bN�++��^=Չ��{4~��{د�����\�83��7f�=.�+J�a�p1ې6: ��>�W���{��drs�x�����������#���rt�K��fX�J^�-�oY<'�V�.��;�v{�̘�;�
��_D.�c��z{��Z{����QT�bN�L��$u<>Yw�z=oG}2��{�(=����?y�P�������vq^��a��{�$�Zێ%g��!��3�ef��(3���Y��-�H�V��^�z�}s�Y�}]Q϶����T�ĬT�dw���X�8��&N���a��٬�,y��i���}W@�aY�U�W��Uq���i$n����hz�_A�/U��|.k����-�*u�ų�82��B���87SjM��^��X���)䢇_;�*�
�{���{���V�c^�4{P���L8{d��vj%-���vlz�^�|gт�9�u�ύ\(�}�=��r��*�<�� ;��p�]B׿(�.,��=�л�T��{��z����f�,�5�`��2�zk�i$X��Ry�Z@l=P���@=ڻ��4��7�'oˬ����6��}szj#RxK>i_��l	���)9�F�[2C�}�hlqЄ�E�<�ц�W�wז�f�m���3x�{i#�}E�CK�g{��.'��(�;ޞ�KfH퍜���b�����̽A���v|)4�gK���Ḓ�G$��/�|=)���*�����ڛ]��f�vR�H���Go�R0w�M٩.�f&<2楊�Sf��t�UG���czP���MR.j�2]�?�c�_wM����V��Qމ��5]�f��9,Tj]fnc�=n��W�Vy�^Į��f̱;�+�;�>|��Vo�:q��S�(>'����_L����=p��͡��Fl�_'�|{��y����vpw]ʳd���|�����w�u���_�׆�_�޺;�q䶔�m`��#�R��־�ܧ��"y�fon�Y�ֻ;ox�av�bP��P��]),��B�ks3��] �q�[G��<���3{\^v�OU;+/;;�5z�4���!m�Sp�Ar��s���]No舺����_�oZ��@Qܨ3�9�D-t��:���5��G���{�Sb��������Ez��fBҬ��v��!�E��y�T*���y5C�m��1P���K���y��I
��w�7��=������9��]}r���R/�7,*�s����;I�|]��8p,�^��ڽ��}'Dw&Iu�Á�ǮJvQ<5���;�"�ɳ{�.�TZ��P7�=8x�wM9Fl�wl����1��4�Sb0�5��t�3&��7ltb}���&�ҎW�o<:G���zG���.��i�hC�ؑ�������Ga���>�ݗ��%򳻺����hoTOVa�.笶z��t¾���in9��}� nQ꙱B%�������ƺ�й�4�z�7ӃDj�ϚW��t�����_&���=��{޷ۇ�+׎W��}f@`v�=�ᚥl�E���]����	z��3���(�.Db��S9ל�A�5]&�)'t��z1�1
��u�0������qJ3X�L��L�Aw��3�،^M�wI�\��������@��/����<�"=eg�}�@Z�y�N��vkḁrg���:��A*����ծ���ۤ�8����UR�t"۩X�狗V�����z��}�0s�sx�U�4v�f����]�"#r+��4v��x;���p�@��ܑfA�Y	)ރ�vPvzNE�f~���q��˽��o���nC��C{ r5�� �C�u�#ƪ;f�Bc���~�G'zvl]D�d٬�>�5=�l�G���;��ҍ�Q]�u��gD�/�9��ʑ����G�r��~�������M*��ӗ�7}j����fB��}�k@�Ɏ��A�ެ���<sn;k�_]ׇ��q��7�Ҭ�$���Uxn�ps��y��N��)�_��_�ʫ��C����"�w��ׇf��74��ȉ�l��<�^n��=~VK�G)��PԺ�����)�;r.x����[��.�cTL�w���3$�����|�����yLW��u#}ޖIf���5�)u�+�jK���E��j܁wM������ӭF��v�/�X�zl�/�΍��6��w��K�2���㨿J^�3Ӭ�t�7H�\���$�׼U�ܞ�w�2h{N�C�\sϝGg������Y��A{�)`O�rX3��ڝ��k�6OVX]�7���GD���h6�bG���nz�����WO���{�>��ߨ���7���
�"��u�A� �fStMݏM�'Q����fn��v0��X�]�;\��Z�.�P�c�FQV�<�����.��WvWo`N�5ǻe�?��~���\/V�Im���/hU�q��a�pĶ��s��9q�u �<T'�}���]�����wH|�
��u����s+q`��p[k�������P�$����.�Ԛ��w}>�,�G�׌��<@x�<*���;}���9�.��d��8>��"d2l����{���z$�M�'����g��(J�xT�x{�]�#�^��oHU<��#.U�[�����L�`��̀������rQKfK��*��Wڮ���e���=>6�nm]�n_�w�tW�$z/�(־�3��q�&�����4����"�e@k,������mJ��]y_��{�D�նg뚘u�e�����6�ʎu"�3�x�=����?I��Ѵ�p�m��2�5���VY�Q-[9�p���TF.��g ���U�g�}Q8k�wu�#Ty��Tlb��v��δ�}�����Na��Mϰ�O+�.X�k�̓[����g)�Y��I��Ǻ���Y~�ž�t����)���w����ܨ��L�A�;�, �ݓµ,dGo��V�@��9R.�'޿w`��T{羗�n9φ�����}�p�4z]BV�����ac�V�uqRs˪g���\U�:X ��.!��'R��=YE�Nޭ�!Rڣ-�坴���Zy�V��b��m��a����;!��Ȫ���;
!O���\��g�P�������r��u"��cl!�XZ�V�z���ͮՐ��<W��ҡS�=�Wԙ��5{�6��=F���BrƳ��𼸇���vuZ:=޹,�s6.�̱~���7������Θ��W�Ʒ����6r�f�>([}/��uK����]e3����o�ל�h�*��{ټOg��iX镚ע���/ͺ�Q�,�so�ޘ�a��D����q�{���x��2O��S�O�Vi��K��todT��juP��r���x��
ɺ�9��OzK�u��W�ѽ}%�q7��S��h
�i�D�xfO�x3�{�{��)ۢ������7y��=��t�ḭ�;�O*�� 5�"4�y0&���t<5�VP,TLN(H:����}������Ş^;��ʞ��̢�s�<׭ 6�^K�#B3�k�.�_!ww�:��F�P�.��/	ga�|K�G�&;��P��y[2C�G���1��0���{6G`@�W�]]�om$cُ���it�j=�Qc{��i;�7�94����|��K�%H�P^O�+s�k�L\�O�
�ɔ&+�J�\w�zSÝ{�^���H�E��.��� Js�%˰��`�l�D�2��v)ܔ��v�p�z� *�e����:ѡAn��έK��Q,ZK�(���]a�}�!�b���2�q=�Pe^�!ɕr_'l�n��VD�}�';�}7o��NԤDwzH� ���dݚ���bc�.jX�+����Fn㧼ۡ�/�z�WP�����17�6���
��2c�nn�IvM����1s���Vv���1}w yV�6�w�z9쁜}�3�w��^���sh�7�d�g	��͚���5y�l@۝]ʼ��鋨eg)oM��t�����8;��Y��K����:d�^�݆Oz]��K��W{��M�B�TY���3�t�0)k�Ĺ\=x��4Wc�Z}��{m�0���k��bwrӡ�eM�jp�Ө3�P��u /<�S���D&�wk3zc0mf����X+0�vE��������.��Ǚ�S�c�J^�Q-��7ܤlG��;�g�(B���)��>{U�k=�MΎ�I�Qɒ]D4������e{����,���ٗ��$8�M��7α�/�Σ�o�p��O����]G��5�����Î�д�ԕ��ݫ�9��%�B�����̩h_M�	����7Q������_���W�C��[`s�C>�L~U���+ҀvK��$�
���]p���\��YC�o�9W�`����E�#A�,�iQ��]�7��lW���j�-f᫺�B����j`�tQ��n�15)on�[�U�t
d"�w:�����<l��p�=�׼IJ��>3Hs~�k��3�qaok׸cL-S���6��*������Tۜ&#$a��3Eـ���s�s)�p��(����c�v$Ē��C�,�V�ht&i��%u�Zzm�,='a��%o��5ϳ�� '�l�z��-��V���6�kòh�w���{��(s&E���K���:ʜ��D4*��Oj:v��ǻEbs{���F�<5a�0���]��K�r�G�[�X�Aδ�^�i�O�ٗx���3#�ǭJM�v�GӢ!ç<YW*3Bө�'v���Ռ̶�]v�-����jQ�_ K��'��$By��!�<BE<W��g�T�CV��ـ4j�b�D�]�]#�������ˡ}�B_3w�B��A5[��Ȕ9reoR�h��:I���5�uք::p�vc�bɻ�oӭ�f&5]�3����Ĩ/3����UȎ�x�;�v�8cDΝ�Y��u�*�g*�e9��9���C+b�B������)Z�t������$�8�>E@KB�0�����Z�3N�Ae�=pOgFgA��ߖ:F�=��Fg^S�C/~oM�a��V3x���[G�F,,���톤�]q�ja�"l�uC�	��z%�Dȝ�	��o��Ml�犳�Ė.�}��Yg-��jtp$f�9� ��i�>F��1p����zp��Op�z�D.�e�.�3s:�;rآ�2)��q1 :��8���Kv��l\a��Jssŋԩ�+�n���s#���wn�.G2�L�O��)<vXL}9�h5�����c[<��qDm����}:Ss-+xˡ�l�� Xz
6�vu�"���)���Q!} �~�� ����;S���K��^����Ї�)ե�����'��ݙ���2�ٜ���ˇw�ud,��qf郥V��]����<�Aګ� 	��b�e� |���Rӯ����N�q��J����kU�\��tY2=�6�<Q�euF��iR���^�[Z���K�V�|r
]dǖH�	I���훍n�r��
vs��V�/R#����bMժ�|n|{!�=eio�_���4OOkst�8Q�fr��3dW�V�����S�Sz�L%x�1J�x��=��\�4��7ݶ������C�;�q��\���Gm�-���.� �,�K(���=�g]&[�ʮ����ra�t��e��`�t��y�Y֢�7�����/1�%�;�wu��I���]]y����z�!V�A�V��l�G��t���=֨�������РT@�4 �C�W�8�tH��O-�fD]P5(����Y��Y«��"�PC���	'"#�2�.L�NfDV��"wq�.*�/X�rYVl��;���B#�>;����bӲ9E�9g\*��WnNI��)�Au�t���	�9kYATA��s8\���焢�Re˪�
iQ�HwY�AA�s2w���rH�"e@U)R̙p.|���PyїaAg�&(�4��,ˇ��dL�*��""�ts�.n�C�%d�4Ȉ�i�yi�s�ĕ18S<�$��"��cQ
t� O"V��ih�iW�G=��$���wpyA՟%�**�1�]�QEAt�'%wn���^~z�?�Yeխ��P��(�����{=�8��5G��t��Z�s�Rn�)C�!Eo3�y��$q�N�m<���Ͼ��/�V{vޯ�kP���⯼h>���1E���Ck���ꅕ=U�
Nd�Q��fCE�=�O8�7��:zP��
��j=rC���
��E�D4�������dŪ�޲�U�u�a�^�v�����H{�2������6�e���$7yY:�\p�R��þT�O3����� �����5[&�j�^�R�p=0�c߂�K+�e?�={�����v�A�u]G�ɽ��{���v�{Ô����@�s�J�MP=�В��1{��=&�˲'ݞF�;�'��'�s�f���軙��h�����҇�:G�v�"��?I������ǝ�Y���1�}�[�-i2z0�R���u���tN2�.��ʑ7���W���L�;sB�W���4��o�/9����薬���0�*����F�Vq�ݪx��ݵ��ޚcѕ屔�u�X,��z�w����C�~�0T�M���\�\�<�3��[.�s4:�T�e8�Jq�o����w7�7��ߥ�w���x�)uSs:jZ�����@z1���1����)�z��)��m?���/Xy;;9�}+a�sFƕ��U1蠏*�L�.^qc��ώV��CxU;%Y���4��,���e1��^��Tƥs�N�V����Y��Ƅ*�0�ٛ���M�PO�r�!l*y��[�9��>���벻-��զ���4��yLW��u#}�zY%����5�]E�kM�Ip5����m1I��l�{}�v�){BU�w�C��[�Vt�|Oj|u�NV���6����`��L��XJ�[���FDs�~�Q)ݼ�n����[��M�*�\sϝGg������W�f��� ����}�H��bv{��y����_Z�������'j(L_s��oQ��{0��g�>��<}2;o'�D��z�[�۲��~�Lp�<{����s�G3��8(���簚���Xq)��J>��T*U9�����]�N�!�x�� ���<��r"�'����y��U�{�]�n-�sf�E�Ϻp
]��*s2��j��}i#�+E@w���m'f�;�GDoט�Z�w��ޑ�G�zt�368�3`>��m9�%�d�^�J��j�p����/��u~���핼�6:��0�e�żJ5���6j2G�z|:MBړ�}���7ke�G���{ۘo�hv�����\�èΙF&���-��o#�H��1d���JG}�e�Ĭp}aN�r�^z@3�����,)��ќ�V�5Z7����;vʒ�U�_��d��V��r�>օ'θS�|W�`*e��-���-Oܲ礶���:��l+�t�#���MSs������Ԩi���خ!����3����Qx]Y/8�YeН���(����'�^{��<���o����V.���t��G�j���>��/ܻ:�������=q�/_���g��B�sw�n}��%��1����̓_n�g)��$��ǜ'l����5�]C��}ܼ2�����G9�K2���*&�}3f��'j.XG�'����<�Ѻ]��o:�s�:!9�||���w����O��j�l_%�=.�TM�٩.iu<�Tf,rj����L���� (�Y�W�g���sS���}LmvuZ:=޹,�͋��2��Cw�J6*;�{u�nls�Q��/Y�v����
����к���jsOq���y��f$��\�G�f�Czʞ6=+��D�{��Eڋ���u
�w<�g���vz9M�>�/fD��W�iي��Ú�8����$��,	�
�lzRvQ:7���N��=7�=��/��80eU�3����㺮a3ϫ*;#ƙ1�Q�;mPm;5)hx}T�:���#���eM]�k.�v������H�j:ܡu=T¨�<�� 5�"4�y0&���t<>�vF�R��u"~I_��'r�ܩ>�+U7���X����O(�(V?�޽��d�Eˬ��Sm:c�7��U_����<��EyoK��|�n�>��V�NiÐ���=㢅P�GC3Q�/q��owٽ����Ӷ��e�u��,w�m �v*���^����;w�߿�c�Y�,��9�wR�OnfQb�Ԟk֐!�ª�����&��̅޼�v�e5
;]���.��j]���i_�/wO��I��5�ْ��X���"���"m)��|��p!�
�]���O��׈�;s(�c�,�4�w�����H��xv����y���X��Y�'�Nd��d�4J>�b,���]�y���'kh9�G%M�:c���1cm.(��o6�߫��{X�����$e�I�%H���P~=v��qsR�q^7�r4��c#i���[8s/i��%v��k��_s���ILs^j��Y�鹻5%�6j,�9����AS�"�&]M��'f�w|1��'f�H�ݓ<'}�^]�V=�͢�ߣ�N���pMO�l�v�(�}��i�^o�z��=a�
#ٓZVq�oM��wL�ͼ���uܫ6�H��l_�"qw��Ȭ���at���D�����ѝ8�
���'S���W����ZNS�<��k}����ݽ�2���+��T񐬭7<�;V�vպ�G�uB����?~�@~��F����X�oR��eL���ǧ=���X�v���i��x���C��hF<*�vG�.�ڝ�����ޭ�o縉O{#�@�� ��|��] �[�&Jw�V[z�	����b�SARKk�����Bi##c���N����׎�g޿\�ﭹ1���Y�w�$���<�r���K�S kȹCF�)�兞�f(��ͩ�w�Eua��L6}�s����Y���.��p&1c��IN�D��Y�t9�{{ˮi��͔��^o�h��f����=���<3�GO����]y�Z��Sp�5ӳ���"��h��;۩ǵ����U,Q.h^�l�'ǻ��S�L���N��zd[�����z/6�{�@�j@9������f�.����O_L+��(W�̖{�c���TNtQ�¯nn��́�7
��
�l���ō��E�|Ҿ&��� U��C��E�fk�n�꽞�t��|�d��3 h�=������V�U����J�8K{5��w�s�j�_K;���c��Q`LGw���3�mj�{O�Jg���+O�ע=0��Rc�D��좽��fE��ff��~G���UF�p{��u���rV��{W�R3�/x�IvzL�l��Ә=�
'��J����4�C�Kǣ��F��� ��C��#ƻW�B㟤�~'ta� �Z�Hq��o�l�{;}���F�X��T���������W�N�c6�)���&����n�&����.ز߉~��7~<�(���V.�8��;'��s�1*ς:����{���D^��pG��-ʡ>���{|B��w+��n��c<�{��a�'l�����69sS���Vt+e�<��;��A��m�r$��,��5��Y��ߛF����N�Q�����
�yY7Q��b�;�;�7ǰ�7��^&�zd��G�ӓ�1�,̜���������G2�LLC3�d/f�Z�v���p9��-�|�3y��<яwy)p�y�6k��źhg�����;}�)��Q�]D�KNS��J��γ�v�Z;�]uun�y�u��m���4���g7�Xq}�R7��d�j�3Q�]E�J���.����[(�Q5ʼ��gn��ْ��m���.�|]�NV�漋�Z	;�h/f<�}�O��Z�7Լ���kc���3�x}S?�/�П��em.7���vqT�o�W�f�<�H/��YZ�qSu��d��=�tx��5 �Z��Ku�Q���'j(_s���Q��{P���W�ֻ��{�q���Y���^S�O��&��U�:�x��Vڰ+�n{	kE�}A�Ǘ��n�W�-=.��Tw)?��!C���X����*�{e�3�o�p�.Gg�#;�\�S�#=�dl
ɬf�<�W]Z��ّ4�}����^3!���]]����~Mq�?b�s�]cm'0b�	\+����r�#��U3���E݀�kLF6S��#����B���`�ݳV�'�t�8����t<�����W�/0�ّjxVf�7G���9��ɯ�t����T�e5\���#H�H.�p��Vj�s���κ��[����茹�sZ�[Á|���xN}�AԋՑ�P��ޭ�A�me+�6���6{+UQ��}���ṃ1����@_l@s`Oݲh��C���M�=}*='�]Ϋ�x��hu�9����ؚ�]fnja�t�11X�y��ßW�n[��-��cG�Fy�Bݎ_m,�G��Go�V3�m�-_�b�ss4�]u��*��W���ٞ뫹)HK�.�{�����u��딌��I��t����;�)�`9>���:ǯ�rs`��;�{�hf/WN�"zj��R��ïz�W��J�<�.�v�r��xjK�w��n|6:@y�Q)�<��:1+dTBs������w���}ursѮp�莙�5��%iYk6�WC��Q�)�a��o��p=g�N���r�"��ϡ�O���sU�w�K:����C�D���EZ�w"��Q���J^��v��,�[�
<��B��|}��;YW��y�-a��hꚝa��V�K�&�&eMz��[�˷PG��X���HN�ޯ:-����}x�'�2kD-w� 
�1��w݀�ҹ�
�/�t7��V�[p�J�i:݈]��IV	5aX�⤬��f��2�lm��f�L�渉��m�����������6���e=k�Pݯ��(O�m�*w<�g�;�Gg
Ω�^��<�g#�^���rc<)=ܙ'��`N���D���JZ7�SCY��B~�r��d��7k��tZ�m?YG[7�k���}:��a��k�4 k�S��*�f�%-���K����7�M�O�ʻ�y�@U���h�3���]2¾�ʼ�Z�JfɁ/�C�3_�=�}T=�6swWPvy���Ә@v{K<�wu!��\SI"��<Ւ�VČf����Ƙ�LN��{�t%�*;Uz����5�vϡ�|K�q�c�}�
Ng�,��N:;C%�m/q���p!Э�ٯy>3x�s�2�Lf>��'�_CQ�bie���u��S��μy<4���o�2�~l��%1�|}�ĥ��˯&.�P�nL�5�G$�2+�[��=�*�+l���uDٮc�[�$f9�H��JcG�Z��}��޿�q�m?F9�+t��x�G{�wetG�hr���FW1ꊮٴ�3@�\n�;f���IvM�s���a'�M_P���u���^������#��eR̈���7kd���N��;.���޴�.�BQ�r����ֺoX���`,2�m�AI��+|���S�}�]�5p��z)��w]=��\Ɛ�G��w)��E1ǞWYz>Թ#��a/�,Tƾ��V�lr�]/�G��W���� gĸNu�}�V=��6��~铦a�����~ӓ�Ys��g�b���[�OD�Y6ll�<��ұ����ᛊE�]�a�wfRËsoh���� �G��[~�9�K�����W�ةhv���s��K]>>�N��徯Ք͸�TiMq�#Q��gs��>'u���
�!x�=�gjԎڷP�t�Z�57x���x\�;��۵\�f�U�a�zgOQ�N�jc��]>���@��F��)��z�H�B����t�
W[���x'����c��MΎ�Ig��K֦8�=qS����[��^螣x��v���C{�ɡ>ռo�<��a����O����W�~h�lt�sޱ�g�ҿy����eEٙ:7�vhL^'�p�=F�W[�.���|�#����x���R��WD��<o��T���XN05���;Y�(�����a=}0�"'���Q��VN�݌����8��p�{_Y`s�����=
P?�z^2<��Ѣ}���>i_�DJ���߮lz�v�*t	��t�mƍ�AڹgG\�Q����"#�W��X�g� �\9C��]Nt~�k�Ӛ�Y[gUZǭN��.aV[�R>z�!�qRq�\k
X�v��c��n��	b^�|���1�%��e��Y��0k�΋W�`t'�U��:�Bْ;}d�!���.}x��������P�_�m�:��+�M�7ѥ03�j,	��w��9��5T��}	L��P6_UǦ�;��ث���U�l�����ڔf�g�U�u�a�@jE�gG��rE��bJFp��Ku���)W��sg�Lɱ~=sSY�6k��#Q} ��"�7�6���x�s�sm�9Lק/x,��P�D�dٱ�r�F�b��tN3�y3�w���_�M��.������'ъv�k��[��@��98;�D����yY7e�q�b�;�5�Y��v��]N�2�U�h�1����������?v�ׇ��!��W�w��a��?�9�]��D�v:�Yz���B�N�@t�
�M�|���.����9���~�>��Y/=�b��NbW�Ӓ����:(ItrS�lM��������:�{
������hu����b��27c�,��D9^f�������6w}`��	WG-�y���p�>�{ /rl������v���+Eg9�_���%��e���ܗ��Za�s62�b�/a.�+x~]]�k�yi�^k�v˙�) �ݕ�5�ێ��hk�����y\�ˇ^�����Żsv��� �rW����mY�-$:�8��#��Xf�Mn3��Mcnj_LK���_��*��؊�/��s�v`�u_v]|w�j��>�Tz_iP�1T�l�]��v{J+9 ���ҳ+��j���=Be�C�7b��"�ˁ�K��S���i�'FJ���5t�|3���oJC.�@��B5}X��v�,����]� ��8%��wr͌�Y�Cݨ�Jh��C�{{�E��[�tH�q)�γ;���7����˖W+��S%2�@cVx�������l٦e9L����fc�ZU�� MZ]�Vz �c�T�Ee��jY��n�W��>��4x���k�w^I�"�O��Xڷm��m��Q�(+A�.?-W��7��!��D�r��q�}�gbe�b%��ج�srV�th��y-DZ�k���q@���4.�wej�w�l�.IWQ�R����VF�mx�R{�����U*��A+�| �n���c/v���.I��օ��:Pڃ��V�Y��F��n%��6yy�i�
:;eV�< x%EfuA'����zd�y��iX�fڮ��)ɠ�A���=G%񾭀�u�t�Hv����c�,b�,��i`��S6h��Ե�ًr�=|Z�3��qN�X$Y�o���譚�9��c���8��xRڝ�E�@T�v[N�n:��9Jd˹���J����:8��t۩��r������)�y6�u*k-�:g�2��}ޙ���s��WK�[龥�����a����%�o:�e!��"ѓ�5�Υ�NX�� �Wy��G���I��=(!m(��x�h����1f�� �zǓ�����E�
�տ9 �\RMe�39:Ҿ��s9ba���_TKt�.�&�[۬ �;��u�p��څ�8�*�_'��dx�1��*���������@7�cJlm�u�zL`���\�@�>�ņ�ug_.��L�z�N+�j���W��{'S������( ��z��BZO���������MM�2������"<[iL���Z�J=t&ɤ�z�Ȑ�UʵJ�ޓC�z��vp����	K>�>��y'�.��?)�&u��Q��*���jU��K�.Vq������H�y�j�A��K�I��!T&Y��w.w�݄O�h}|�z�2�|rҽ�m���`��0�>�o,��h4S��_C�rغ�-S7���2'\[|���G;�6�X��DF>j�xa�����h�~6�n?n\��`E?��)y�?�F;ױZ�#��&�w�w�[y�)��}1:���]��Ŝ��'�Z���קE{��곒����T�ݷ�a��Ǭ|��#&tO#����EQr��THr��E��ޝ�YQ�!=H�[�4��B�v94�p�$�.\
�8��r�N(��rp�E�*e��%:E���|x����D�wX\��42JtĂ'3��0L�u�EQ���������Gs���TDM8���zܢ;�vA�"���pu�r��Ꜫ.*�Bi	^t�E��.��"r=�wA^q�I�!&S���]9�F�.���u+��Q=vD(�Ů��wnd��w�Lt\2#�w^y�2X�R�"�9��	ur��ܯI���^9�n��u���j�)�Վ��:����.�Aw<gω�rԗ��#�:ʨ�N$�-'q��g���p��Eq��s:���?���-	[��z��!�9�ݔ�Z�_$7%�(򳛬�*�������f�;�=���/�J���F�*g�h�A)8����J��2gx*�xy�9{��A�;r���1��V�хx}��3�ۑ�ٙu!]�{+x��S�O���"wyH���v���s��=F�W^�+��<��q�X+�=8w����_k1���p׺��t	�`�o@�9^T9�Ι/~���+��yYG��Rm����y�T,)˘Wܤ��B:��@����`3k�T���`g��;r�������m�����c�l�=q�`�j;�p
]��*�3)�fI�v-!�~=����xV�X�ٝ��|b�Y�J��B��u��Ѷ;���n��_��{�f��}��j�rQKfK���i{��Z�V;DI�����T�t/�r]����Ǭ��P��s�Q���t5�.#�M1���m݋%�>���V����~}�i~,�����͏N�؛/��ja�Ft�15�'�����Y����ƻ�Y�y7�ޥ1<'��yޞ@�~���ޒ7@63���j��ȋ���F.�����S:m��MO?T{a{�g׳�f�x��0��u�x{��G��B��~{��[�zc��rc������!���1�PH� ��cvU��fx�c�k�Y�N�&p�mVb�K��áv�ʾ����%r�,�;�����X����y����A��&��oEM�)m;	B�A�p�(�њ����i
�){w\1�d�3�)l˓D����Ss{:��0�Xڒ.A�������6�+@�͹ˣ��o6�Wx�s��8���/���G���,�*kr�7c�~�'A�^ڼ:��^,=]�]zlW�,�*��������φ�z}'3�s���GLݚ���V�q�H��ˣ�T�7��I�����ً�g,�)l����O�}Lm}��h��z䳵��O`�$g�j��78��P���͋���QS�=V�sG��(7��=+C�*�z
�����D���l�n���_�H;�Pw�K6=�:=�dQCv�/�(Ly�P��.Y�}���U �\�>�O��ǕZ�_r�����<{�$�+@xV3c�);5)h��Mf��T���D���n|3������E�rx�u΅f�WTw���Q�u�a��� _�ӳQ)hxi�P�u,��Uq��+״�*���'\����]nP����aWt���@�ǥ2^L���	{��G�q¯{6ީ�2��^�a�Y�>%��>��l��C*zk���̢�}Τ�\���Ul���y��<F��B^�P��W�(sw=��R�%�4��~����t����2T�`�I����eM�_��*�߆��KdF�L�������]�]kٽK;*}%��Ta�f��B��	u���E�	�O���k�[_{Op��=(шip�zEYR���+���k�a�#�xFEg`;�ƚ���-n���݂�nя���&�Tn,H]nF^�_J<��x)p |�x�����C�I�}'N��-�1��	q�vM�н��sު���nD :������=�JcD��vy~�7�>�����f��~��nWȢ!��9�*�J]��`gzTM�����ԑ���H���`�,��_D�g�ђŉ���ᗯt���`{=[���t]���h2�#�hr���|�LK�;f�S�x���k�Ǎ��B�/MnK�V�C������d��o�\/R�5��q�K����^Q�uc��6��~��:^�~�q��&����^N�F�����5%�6jˀ��0��@9˸�wL�͸���8(ǯ����~�Qmz=��ͻ+3�vL���v΄���r��VyPg���`R�O�r�z�����F��Em_]�w�r4w׻t��yY/}�l]DqR̊�S�����C�>�P��ΨS������H���][K��v�Vi�}�S����.���3\���&��@��F�b79/\�R��^��m�c��X[k��s��3�>��w&Iu�N�A��J˦W���ד�*'o�&$���2��M���ٴ뤾wduHol�c�Y�PP�t]׮;����k�E�:;�w�+��z�r^J"��1�0Y��t7�ڷ�.���n��#5H_\!ux ���hU"4�~�:d�n���s�ܮ�p,t�aN:l���(ApE����'�(�������,_[����<��a����t���F�]}� j��0�U�����\/iUe/gh>�A�/ǢJü}�R��vhM�|w��l�[�=�OM2�W��o03�r{���޼{*83� nL	�|�B�u����b�.��]��_T,��*�`�D��y�P짳}�P6k���+�p*�ڏ\��z����i����X�Wu8�,�}��]�E�ȝH���@�'�P�^O�ԭ��D1�;���W�+�fŐ�s��+��ޝ'��+���3Q`O���A�����I�>�)��?+O���>�}��1���[OtZ=~��x���g�U����jE�tz�sU�Zj��^IH��Ց{U�&���g��9��3�u���]c��7�xg׾`~F}~��8�P��t��ٴP���j�-�/_��]djx��.�蝟��]d٨���\�ì+��{:'��&xN�;�H����ɿI��vg��O�6�����)Wd�v~g'#~8��eC��hw~��x^e~�<��IE$5��E�����y�^{f.�o�Jʒ;W;���5Sr�Y-~�g��Y�m�Ӓ�Q^�g�)jK�'�1dݘ�r�m�@�`]R��Z���Ev,�ɣ^k��V��p+1e}аn{l�_v��Cyv^�[ؘ�{�0��8�p���3ۿ�	����r��oU�ߦBws�to�w2���S��J��_�������&����@:��t>^��9���w����d���7�]D��73������*��WwfL��6��E^��� �����՜U};=�����9oe1W�u#}ޖIf���5��]���-�{w�H�{��7�OI��Q�|����eT7<B���NV���6����`��]�z�ӗ�t���:#�����J^j*&\�E���П4�B��\sϝGg�����#8�����e�oU�j�A���� ��,	Ò��ݨ���yz�kf$z��n����*�7M��d���;m�oB}��1�)r<�������@tmw��;-A��>ףNO�O����yY�w���[d�_T,5=N�Wr�ƼЁ����� x�*���㣷���]ψ�g<ͮ ���:*5t�|V&��� ��{�
�s2��樞f�p����J��y��~��=��et��j#�u��o�ޜ��{�f��ޮ�s>�Pu"�8��ӵ�3H�^�?z�jb�H�Eepp�����'>Zs*HM�F1ǟ�)��{s+�^ZF)c�/�k��m��Nܧ�˄jsX3�K�N�nFf^�$���h%'�V��[��W2���h�y?`�=�a]Wn�ܓE!�)��s���V��]�W?\죔K��Ы�ٛ����3����@_l@s`Oݲh�W������_3-��v��ж��z����p[��ʬ^���^���b���r5���;y^���{�[���{�~��Ά�x�1��H�7�#��J����_����F.iHcы��K�)�G#��ɺ[���<%.��L����'?zhv�$z��������j%�����d�
Wo����u�'����α�Zs`�ю{9{��#��Gb����{���w�r�>2��D��f˭��q�#%z�]��WV�}����'�jY�L{�wz{�9���O��dط�Lݗ��N�]މ�g7*sMz+/�Y�	4���ri�=f܀��q�X�|槅���cj;:�}�7s`���Rc�|��q��3b�8��}){TW��=VϾ�0<���}/��T�� \57�ׯ}��9�]�پr{�;+O��H-�A�)�i`ٕ�ר��}1"�ۨZ�d�>F.�d�Lﶞ��R������7�;"�Grd�e0/�+��'f�-Ҥk3r:���%s���ʾ�M���u���[��D5�-b�4����2�l����vj��4)���Ukn�ל��ft�ΛC m�C{�Ȩ����j��Y7�G9.涸W�om����������P׺�g&�����N3�m��^�ѕ����}v��ˇ�x�G\�Vi�uGz0�K5�u�)�cm_N�}�v�L��y�����zz*��sbN9�6�#�\u�B�z��ܑ�h�TzP��.�3�VL�����>���@��>�a��=9��%��>k������ʉ�*���,bxv,��巸=�V���[]�$L@{0���
���^����s�t��Yd��ގ3`5�B���o�gv���WΊRh�.�#��#prЄ�s�k�O��"��2�LFc�,��7�|����
����wUw�^���u^�� w���.l��tJcD>�b,��5�&.�P��Ǩ�B:&}�%����\�=��D>\w�:��Q�=0&9��3��Gh�,��R]�̨a�����+�|&�t4�jxS�6k�gHeTy�X����c�_vͤ�9��q̘�]�^�J;�û�k=�����=d��Yl�E�O
�K��ѻ�q�Gd�	�vW�TGuՏs^Ex���C����Y*��~\p�+������M���=ء��� JΞ����}���<8��g�W�g]5���b�*gJ�IڑWF�:��i��\�m�w�S.�\T�AJ�{�U��do@9Q���Q�^w<Uq��^� ��߬w��_d��]���a��=�P���k�o�5r�"WrV�1;X��d���y�/�pu�e,9q2G��Ю%zM���YX
<���ӌ�����]QPƙ���E�����x������n�4Wc�Z]�c�غ�⥙
��q-v��#��-��AI�6����^v��8]�7��r�ݷVi��}�S��w��51�j9OU�}){MK@k�q�ǻ$}��k�����Όɡ���dC��{nz��}�s��R,�w&IuL8�E�e	�<�߫-r˿oh�==�J^��a�^�ql��h�������1���@ז������^���>���E��}Pk�k,ԕ���*��S�Bb/�m�6z����K._�6⼣����*C6�ۃ�ݠ����2LsA��_�����'k0�|]�Y�k�Ϣ�ٌ��T������k�,Y3�Nd��H�P=��{�8������w��v%�}&�w7��G�q�ڕ�i�Td
]�U��D�D=�2�ڐ��xf�[=�:��U��vO �[���q/�Htf��_�\s��ރP櫤�-ROi��Lோ�@�����}����RX�x<#<�e+���
��2�^��)"z�Ϛx\�?��l&�86$��W^���E����^@dN��q����QΚ'u��Εr�e����5J�hZ�����p�/�W�8յ�k*
x��C���Q
�}��^>5��'&��7��;��w�����>�e#��x_Cu�a�e_���?s�rT��{U�Q�c�aL+%L��7��t7��C��?��.��^����>���3�^��b{�N�~�CUj9���>=�mW��ٞh��{}'��Ń�v|.�WY6j��1sS��gD�>�y3�wƺ�[��?gK���co�>�y$k;$��,��ld�n���eC_���J��zT�M�0}~K}//�.�=Գ�}�Ⴏ����ݓ��qPk"��"�|��D���D\�:����M�g�w6�`���ځ_'=|�ׇf���6��w�����y�.�Dr�Q5s:O��Ef��3~�z�e���o��`�d�R��f�Yˍ�*/��F��,��|�y���4ojt�����j9�7�����N@|l��[�<�e\Cs��=���ӕ�9�"�������71Ӷ���=`��3�?��ޕ��4��F�����ҳ���6P�v�q��c���Ӝ�]5��Y�����׻Y�¼��ݲA�)�qrX5 ۵��/E�'j(L_s��j�˳��f��Ѯ��h#?%�%3o����-�vp�@wϢ��.�{�9gp�ՋV㿰b׵:�P:��,�U���:�U���a�E����*��J`'��'�˭9��n�b5���`Q����N�5��m��9�5�SgVq���q�y�T'�9��fvo�&�y�+��1ތ>�����)� < z��T���C�À�jd1�"_Nٕ�{���8�K����t³���w)<j#���@� =��xR[+� [FQ�rl�׺���C�7��_d���8�ǉ���{�
���j���y�$i���¡���惘)�bYo�� Y����>�c��y�ޜ��8�fl�<��t���딽*�O��y[�K��^&Fp�S	_j�>�fb�(ss(�ى�(�k�;�6_�nV�ٵ�-{T�f�9g#��ä�.�:wȩA��c�K�6_��sS9$bq��f|ȹ{�n�C�Pyviڞ�}�R.�7�x�/})�~�;|J����6*%������h1��W@�2S��:�nES��9*�r�+<��p�s���$�]"p��M~���ʧ����Q���>7,��y��vNM��]6F��r�g)�z;�W��~�s^�����kr�}�:U"�0�U���N��'�NU΀�y<+R�A�Ǹ�w����9�ھ��9��8N��X�YU��tꠢ�4�e��E�5�rn�'o�,�(>t��ηe�^=�
2�3d{��.�e��+�"���T\J�7��5�r���]�VxD�9��L�� �����wϨ1:�8&*G���W�3U�����ci�cS�����Í�l�nx�զ�˩[N��i��
-���X!�)4Ĵ���w6{9a���9$r-[1�/Ml!��o�Z[Ps9yU����y�zN�ק���4�����q֌D�Mc����廷\�9sK0Ѯ��|+4Q.Y��ؾU�o�	#�h��#���#](��2�Ӆ�}1��Q�Q���j�O��/��͚��M�+��rz��N��J_)��k(�rR�v�ç�m��\(V�<�,1>�����[�x�h�����4a���Z��� �:2t+��̋���Wt��]��3�9M;8���[�Z�քx��gyW�j6�k^���\1�I�����YňWnlη�02bq�	�PՎ�m���M�CU��mu��#��q�'��c�UU���6we�:ɍjYY�W����m��˃�)i�����Q9����2b`NX�6 �yR���5,3c��m����p,�~�2�wY�;�Su�"ժ�]����=�*X\��7�����0S�9ܫ�KMYh>�[�z���s!
�$�	e�o��$I�n؝��:�ܹM�Go	���y\�C��ٯ���?d����*G9�h��ћQV(����ow����-��8$z��0nk�W�u@xk�Ə?I�U�nو�àr�,鼝�W�Lja�ǹhf%�S�T�S F����ꕗ��̱I6�3,^޴�����*��_Q݈�j��luȋŻ�m�=�B�+�	*D���y�6�b̊�g�o�BKH�ܩ(��#PinU�sv1����V�{8�%v�yu���o;��KF�|_Ilr\���W}�c\+���B�,�l��ʴ{�D�v�C��`/l�������>j'=��m���v�!�A�	�`t�\�՚�t\i�����շ�1!|�[�٭��í���n����
�]o܌:�&���<C{Y啌��^v����q�̡,�w�h@T�ʶm`�E�]�X��Y�}[�w �\�=�I�a�=q[�5��.
�D��E��ۼY�x�	N'��S�<l��G/gQ|�@�/.�����j��aQ��sT6ޣ<\;:2B/���H=�7�8
�� ���s�(A�l;b�}�Y�>wL�
�.���@v\gv�4㭏��+x�a�r�@����%ڷ�ĎB+����c�R�w1S��sJ��ͧ��3j"�VLГjw
�c-��7�4�)qiw7E��YjK�®b�_2Խk�	����3��mh
r��gU���Sigc���r����˜���u�����=��Kn��^]��g;dx�pi
DQ�� �ϷwRK�&:�����'s�)��"+����vy�C"���Ad�ȏt�9E4�p�y��J����<)�9ʨ��u��,9�<�N*��)8�.8�u�n&z�1u$:d�s�N:��!�{���Ke����=��¨���=�Q���A�H-/���]L)�[�c=4r'9�^���r�����{�y��q���*(T.9��wr�tv�4]O�ӗi�����m�/��u�*���3�t*�iP^nܛ����[��DE�B�.�S�Aze��L����Ao<�Ό�s�g�)��%��<��f� ���9���!9P�2�TZ�.(�ŕj������e�2�*����4BԂ��ŚU���U3Gp�$0�)��yB#_^Ut���Q����}WǦN��vݡb2qfw$��Y�i��%۝Hfr~�%��	ӰU���]Y�]	��5��ݧ����x���M�٨��;ME�����������R�z��1�������N���9����y;��6.����Kڢ�ZUE������.�|wEFbs
��/�$*�{��j�P��O�Y�}�rAu�S���*Y��^�	ֲ��}QC�ǜL���L��%��c���kU��Q��M��a��k���=P԰'
�l{�I٨��oFm�G`��6nUp]۹=Aa�B^����{'�W\�Vk������,�G�5�G)�cmm�Ġ����[���{�~��=��J^�d��'f��q�a�nH�=m!잪aw$yS kw��=��>�7��C����<�J�X�5�a�Y� �g������\��YhW"���=9�S�/"ڞ�X��%�贀ـ�aL%��Y��(sw=��Ի	g�+�Z�^�O�[��&ܜ��Uv����:!tΣP�d��G��9h@�[�W���׈�1�2�d�i��K��Vn�4͞�5';��.{���[�̥͑���S'�������G��g�z?A�إ��j�ֻ�����L���P}\뭾�������L��~�u�����)N��	�)..J/>,�O��{"�<���Xl��k��G���8�F��g�w �I�E�UC|0��	��2d����vz�K��S��k	�B�j=Z�Um�7|:G�]̡Y�4���gC�^7��y��3��Gh��n���%��rbӘ�Y�[�=:j�'�R�z3�ٯ��!�Q�49b�C�#*9�TUvͤ���+P>�Y�C���zn���讗7ed��w��b�R�5��q�d�	�Gexew]X��Z�:U��4��V{���抳]�̜3�'��f�|f|\�u����Kzo���g�n�f��_�A񽢽7�m;�t��f����Xr�d�L�Б�6.%�ڪ,�y�A�X�	�2�N���r3����h�-�b������i��^�9M��*Y�SjtԴڋR;\jY]Q�e</��wꄫm���;��T*��z�fGvkU�a�zgN��$���<�G)갉�9x*�Lu,�z������MV{;���~��,e[��X�y�ۉ�c��MΎ��}%���/b�p:7�㧸�_u�o��y��to}%u���>>��;�"�ܛ7�y-����S�+Ĺ�|#u\V��U�?f�7w�ep�yC9��Z�5%i|}T�:�vhL^'�p�C�l�G[�/~�r:GEO{ǯ+y�=b�'A5}��b��$���{����yp��/M��\0�m���X�� L�Q��˛I���^N�nfD���1S��{a3����у���E��>@0Ku�Qi��B�� �;C�AX+v=�#�s\�ɱ2���̖��vQp$���O�xwꀠp׺���pL�P�׊�hwTN�a�����fX�5��;�7Ý幮�'�}������g�9��2�@/
�p*�gj=rCk�/q�~�0�w���H����x�W����Q�)w��W�T����$=���;���u�G�2:~��WН]��>�ے���Bw\�-��_11�w��j�t���I�$���c��K�U6'��I�о@��}]��:������R��9�UD7\�@jE�gG�5\�Ody���v9��z�[�ˤk�%"߾97f�힓a���L:��5�r#^} }(yCxc���E�3R��ʯ1���c��t�(s�Yy�98;ӳb�S�l՗�nja�Da]f=�
�t��ȝ����V�OxM��R2���|??$�dG�N�㓃�*�ਞVMզ�ݕ��Tb��BF5u��z�{�Ns��>�;T�͸��u��jѻϹLK3�dT�M����]Q���s�3������|���_-��^�����s^W��:}��y�Sg�^t�x1r��: �HC�ύ��d�D��5���(��1�9»L�	2���Gvp���M7�i���r�v��N��;���s��K�w�ؔ�j��sô�\�������;z���ל�|���/���k2&R�kb�Y�{��R�@�{�-Gagv>���O�@^�`� 61�▧���w����LW��u#}ޖIg�2�����^�s���a�Su蒽���f���n@_y�ʨ����]���W:'@�M�u�6�������G���I��s��/j����}�����B|�e
v�q�P�ͿQI��c�srkz5�)���W��_y�]r���n�TJ[��F�����_l�C��'eas�Y�c<��w#e����C�1���<j<����@��^��W �8Eߥlg���x\�U�S���Vzo'@|�y��K�Vz'��*��'��9�@`��@ް��/Yٽ��Y�����ʁC/���}�F�9��qX,����*{�
�̦��'�s�1/0�k��J�,���#��y(O�˴��ƽaC���wy`/Y�z��O���C���'q��5�2��9��{����aO�_j�4���P�ne���s_H���,�	P�^_\��� ��&������'ewR2��xNŧfnja���(�7BƇ�ԅo�cճ���׵mÈt����B�9��T��N��8�O�6���k��CQl��-2i��X���K5c�\:X��LK,��sC��L�m`ZrE5��C{~}H\�����ؔ���wn-ǔ�����N��4�9�]M�Tr�wtR�(�jpW�Τ^r@��})��#���gz
�6*Z�9�\.��q��(�l{O���ov�!#���*=�CJ��qY�TN~�п�nR3�g�Y���
��(3��⥙��׋Sߗt��g�&�	���Q���������R9j�v/���{���w�A�$TOz��N�W�j�:�Q�q+R��^��, ��<+R�E|�X�>����v�φ����ʨ�+���Q�n���lWE�ݚ���
��l��\�Qe���܀��Y�W�e�d�\=w�=|�h敾������7��ڴX�z䳾s6.�̱h��	��lY�L�~^�Pf̳x	�`����~��=�z!:�7o�暈|�̳���y;�W��j�	M���uP��3׈a��א��5�I*���ѣ���-�˕�s���)�1ތ>��w&Iꆥ�8V3c�JNȮ���0cʽ����ǵ�c7�hf�̋�p�O���
�D>����9�u�a���>��3���7�>^�߸��Y��,��K���ٱ'��nH�5nP��,+���{k"f=)�踹������f��-�LNF�#�PQ����7dݤG/�@<�b�<�ܡL$1鹓6�s�*n��}�ح�-���GjT��'����A�O�ad��*q?m[���'��W�+{i�;����6�α�F�_(�Ņ.tY�*=�������xC2w&�-�z��Q=9��v{O��ju��~�4�7�%_�f_l��+�s2�����z- 6�D����^�����'��Ni�_� �'����l�e��^��}�
�Ng��[2C�
F��mo�Q|v/�e���ێ�SW�����cq�z];��ľ�D	��OI�[2Gh��T+s�u��&���
R�=�:���k���L�&��4�\w���5��c��#1��Gh6=�ɏVg#ϊ�fg��9���n�%���K�x�{:C*��hr��|�eG1ꊮٴ���vJ��n�y�] �����&����zɳQe񵉋�K��n�{�9��^�u=}pf�[Y6;(�.�w�ev辛EY�}�'K8�M��f����p=�هZV2-�$�e���&��hn�����٪�gs���8=�ve,9�X;gBG��L�ŶXy0S���>����'�����09<���]S���W���wKO����ܦ��,�VV��h3�磪V{ ���V��.�+�B ������F����8A:�},���ƻs1�lV��
[�(?�^d�㟢��h�������bw��8y'��E��gAE�AY�K�ogo7���[��ĥ)��3ר�a��`��]�V��f�U��p,�x�oArwg�f~�=��Ks����fG<�7�9�]N�w�$�jc��]>
|�Օ<��u�f���=���Q(1��E����s=�z��}�MΎ�If��$�9��vo���e_���9�+�`ty_T_�$��R��g���_^�ql�KG���g�{���o_���f㸺��9�WS�3U��]� cUҘ1��i٨���>�ZD�И�O�ᷨ����/Lϡs3q��s{u^�5j��+���4�H�&���*�u��;Y�e\>�j���s���ۿw���O	���YS�\P��K<���|d��Bay�P3��H߮���+Jo��f�f�d>̛+S�,�W����Q�WL&��;fH{�� h����ڤ�6�MǨfu�~�v�o�L�/q��/$���J�8K�2��&<�w��i�WI���'�����ӰW�).�ۙ�W`�V�7^����&.7�1X�T�p{��u������3�O���yK��8d��%#;�&�����.���L:�Ι�Q� r5} �����g]�ԛm�k�ͫ)d�c!�坹��4�ƶ�X�n]���ĬA8��Έ����V�����Tl`������q���\�]{��.a�SM�����sT�c��L�~<P�w�lwZc��th)(˝�&�%��癹�+�����Yi�3\s9��W?��7{��B[��/�B98;���غ�Nɳa��7+�U��J-i���:>�'�<�?]s�*:��l����T���~������R+�X��d�ʰ�%�~,�Ϯ��/�Kjz�ud�/gn���i�A��Vq�v���4,oe�x{��̿�����3�dW��6OU���^ ��n�ݽ����6t��p��02˾^�;5\s^|�S�a�Y/=�b쪪���ӛ:���v\�&f�G{�?��ޘ���? 9չG��qKS��R;�������n�fHSԡ8.�L��8z�y����E�J���=Y�xo���+up�yv���s��M
�P��*��*�f��w�ͣ����Iue�?a�Q~�Kڢ�g�Y���_M	��6Pe���0�w������~�z)r�}�C�G)�=�+��^{$�0/�9,ݨ�Kw�����xE�>��Jhp�u�VV7����E�mv��g��a{>}U�;#�#��<�@��x@��Rsp9�@�7��YF�3}�-n��3��n��^N �`�Cs�Mu�Bº\¿���5h@�Q� hQӗ�ߨsQ;�B���܉W�s;wj�1����Z8���6x�i#7ɾP,F�%w�X����<�>�E؎N�����;����s��Y܋�Z1p9�A^�-ԭR�ivun�=U�m_�G�#�嵏w(��$�Z���3�b���n�:g�,׶!jqK����}�pnWސ-��X4�|w�8�M}�ӀT.�z9�Mc�{����^�ʫ�z��[=�bC���%y0g�|v9�.��倽flp=�fl�d��w�:½.3���u�g�*${V4�mم?%}���~7|9��Zs�Q�A��g�(Һj�sgOj��/zM�?wI�'\�����F �����8.��<��jׄX+��Z'TW,'.����#�	��ˠ,��R.�:G����:Dv�|/���b��㛓T����c�uX+m������ɚ�����!�^j���C��Q��=�m���[�f:W�O���U�py�L�G���ok9���n��&"�'�js`���r�r��W��xeGuߣގsx�edp����8Mu�����yQ5�5{�ڹ��ݓ¾Ա�_-�/����Oaۈ�>���9�;����������F�G��b�T4ꅑmٔ�P�Y��<��J\�x��2�#�c����C���0�:|����:r�fx]}�e��J^�����3ǧ��Cc�g�V��] k??e����A�2顚��ZJ�`<���]�{����ъ�{���kku6Q�t=�h
޾��k)�ƴwh�ʿ�m��
�1�7��?j�8s|���=ך�u��!r\�2Z���q�-R�Jm]��,�gg,�V岢�:;�(���w�T��p��Ǽe���ePx
g�X6ev�S�X�{��t󳹛�w7r{˹��ިU�,�s���ܦ��{��Qܙ'��`LaX̀���R�U����v�<��J^=4+L�_9zq�<m�΅f��uGz0�K5�hrkܾ�C���Z�7q�:<�(
6��D����R��vlk���G��[�.���Y}�p�x�C.��Ϟ��<�9UU�8����Aе��J�x{L���|�<�_���yx����_��]5��B�k���׿���qU�2�7R5�H��م)y��VG�(wk��W��ͅ1w�l�V���t��=�['�f�����P�Ng�:�r>�468�Bչ�5E�q�r��Eo��{���[�"z�2�M�,�z��1q0�E'{��N�GnA*F �P^�쎉�^���-V�o�g���Qc����1[�(MgH䩵�g{��&�Gh������3��Gn�^��
�S�7�l��W���C�4{�dݚ���O�1�9M���t�U}sC�/C�#+�b�M��6O�{�����)+8�3)7�}�+��m]7h[�f4����RV���b��8�.��u5 )���q��R�K�#��ѯD��|��ߦ.>��"���8�Jμ��y]AF�g:�=�wW�HZk:��f�_<ɜ�;y�	.�BR�GU�O�Kһi��&��*kg ��}12o���d�%����t�h.t8%V��_GUf㪾�/O����>�&.�0u�a}�S��|�F�.Wk3o����mEw��lÂ��c,w7�ӏl��v8<���Z�3�ټd�CE�[b�=@�<���{R=ټ��o�$*y%5��<�js���\�2��\I�O4*�M�ظ��E����L=T��ە��_i̔P�D����p�C���9H���<����^�,�T��'0��L�1����O[{F,�q<WzJzS壳].K��a?xT�v��O|K�����1ӻ����8E&@��?{m<ou4數q@=w�s����,��5�Ń��{g�k�Bր��e'���9�m{��=��|i�Zc���ˊ�n]�����[N�O;Bu��,���J��씌�,}[ؼ��Rt�-�/ׁ�a�_
4^��V���r+Z�,���!��:��36�H�'Gh�,]\	���m�*q�U���gxլN���\�I���;;����!��f�g^��Q{ĳydU6#ux�j�Ag�\�髩F�ko�.aA�	!��5XG��ߗ'������Cel���,EL�5Uvr�������L���n�Xz��g�ޡ���K��-;4;�㩚�T��u�C��w��Zb��2A�+P��K�Q����kC��\�c�fC2�I�P��}G�n�f+�7S��W]�6���J��cL˦���ѲIt��V��$1w�ږ�������L�ʡ�,�zg=e��C��<�+����d��!Pw2�]��ǀ��w�Yp,�Ɓ�ɚ���6PG�69����ټ挬u�P���8�z*����vT+}s�f��a�xI�k7�?)"�4���w��i�Q��;��tI���Ӷse�z3���^�=��m����ls�d��t�Ӊ�����{�5��1��A�A�'$ck��t�.=�'_��f�z��
�a��W��������>�.�����ԙ.����T���a�n�9�e���WR�)w>˴�������ê5R�s�o0
J�����]��F�j�1Ĥ�n[_E��3����(e��u+���g9�Y�X�wnblQ߂h��6�e]� �9u��1�*�ܓ.�1r��D�.i�������:��NW�=�ۍo)�z7;a�*1��I5���lj5���t���u�8/�?J
�w��A����U�%��M5����EҌZ�}��w ���*�E��k��4L�{#�_ k8Z�l�=H�%�M��J*H��{�K��E4�Y�+��#�I��s�(����i�ԧSd����e�\LJD�\Uʑ��\]��Y�:����؞dN�;���:�yЏ%\�䦑E\I�n�p�wq�U�"����GPn:�t�14�C��*5Ȍʮ���'���<+�@��kU�X��HLP4(I��"�;Ρ�'H�aF�T	�u��R��Lҡ ��G"���H���sC>y���/Li"�2%d�#5#�h��k"�Tf����[���aB2��wc���tEj�MT$�����'�T��U
a�;�aavh�<��L�A"+�p�J����Ei�ֹ��p��ej�Fd(T�:iP
�54Ӊ�0�������Up��ڴ� � � ����Y��|�{B�>$Pl�nۆ.�	3�k\q�$�=i�T��j�U:5*CaVR�v�~+�R9�����t3�������$�R�X0�r̨�}77f���f���k���kw���ɞ�xJ���e�۩/v�qo����[�?W�<Ea����^Z�9N��)��٨��/vL:ұ�-S��IJ{f��U�ʛ�Wc��U���3o������n�}ݙK_L���ZįI��������w$/��{����Z�4y�'e1���ᢻ���~VK�G)�uT�"���2����;�{�ռ,�}�fU�@��q;/Z�j�v�7�?L��ɒ]51�s*5�gq��^��U׍���){
����Q}4&<ܰ��3�q=Ls>���G`�Y��q�Ө���K����M��p;�Y��+��xk2N��f���f�&�Yq}��62*�}�W>�.��*a׳v�9�ﰯ���@ʣ�0&0�5��t�9KC�����|w�_a�;�1x�a�.k���ou!u.i�������#� l��~��x�<hw'�W�w�j�܍�����s%��o.�j:��eOUqB��,���΢<d��i�
f'''_Y6�͐�i�%P�Tz�7:�]Gr�Łj�gg����!�_�rկ�[�$+n3(��)O����2C�`��A�V����ܝ�k�yq����!e_^�ғ^y��;�p�{T��>�t�6�	Co��$��vFeN�i��S�flz����=l�}�GLE���Z�(�������w��4WI��̐��q�4]�;}Sb(@���=�����B�\���WǪ/$���J������3�����Ajg�퇔6�ev��q�u���ɖz��P^J�>7^����zX�)���*����ހԋ�b��(�A�M)�9�Ǔ�'U4��\��䔌�|rn�IvzM���*gLٯ��@�O�O�]��G���3�Z�gUW m�C��<i��(\s��/�����ȿ�_���o/��,\ڿo�ˬ�κ�1��bs��&xN���R2�?~�����$k#�H'X;%]��ɻp������ܻj�*��+w�8�u���Pk�ެ���<sn;k�}�w^��s.9LK3�d{;��Y>�W���^�om��r�.t��D�c��]���ׇf��6��ߧO��Y/<z�� �-���w�ˢ��Z������S����m�k8��������9q�L<zh���2�Q�������7��K$���7��_��i�.�V��r�l����ȓ�C���o��ؼq�K��ƹ�2OZ=�xvqn����zs~5Wd��g(eLP��.k�AY����sB\KĮ7�M�f���G��X�}���ذژ&;^�w9B�͵�jc�ʺ���d����,��<��܋q��Gĺ+�����y�\\v[�c,� ]۽�p��ο�O�m���It�X�u�/j����g�V�W�@L�{ʤ�bћ4Wl�K~Ƕ9x��Cܔ�w9��*���
�,�y�]G)`O�rX5�n�"wy%�=ρ{���&�u�m�OPY�M�P�����6�=Q׵
��W���8@k��)�&x@n�Ѕp;wt�����Y�g���W�9^T5��N
/����j:��a���P�;��5h@�|��t�SUãٷ�p� QxW�eDz@�f/�pTF�9��qX,����*{�
��9��F����
|�ŵ]��fIzz�fl�+��T�Ƣ=aC���wy`-�����]0���<)l��۞ʮ�9�WNg�*)l��^�m@�R�����fo��1�2���T��y��k7�7Er�(�n�:9x�DO����j!mI����^r�߱�k>c��S�e��mL�@�����]�]̣�	���t��^t�&;})��#���gz
�6'#�7֝tZ�=�ݔ��tb�s3C����:CK��o���zhtvܤg��Ip�7=�����z���zc<�q�;rؽ��:��ez3�m���V�YJ��m���!np#~:�>ce�<~|9֏���f_���|\�4�QL�@E�\���LnN�wuP���Ò����,�}�:qk�{�T�%[�rڇ���Y�b��#�g��V�Ug��Ճu<8M�K�̓Q�=�����*��*���ڥ���r����=�iv�+�b�>3�*&��Lٯ���r��\.5,dL{�}���;�?j;}���*r}�շ6�>{ur_��	��雳Q��*�nf�iȲ�l�n@_Fr�!�㑆(GQZzW��]oh���z!mK�Θu�V���"δ�<��蔽�*ZU��f;E������V^_m��[�mk=�X�jsMC��e�D~�2����?վ#ޢ_���U��Ug�:u�jA�lĎ���Bv�r���Q��M��If��L���R�\s�y*�=����x��/ǢR���45���U	��r����<r��
�>���FIeg����i�+n�W�jc�KOhg�n%-��Q;65�}�ܑ|k���'��I�����:_���?p_�?6uJ���R�G�P�kߊ�����Ұ�,ÐK��\8@���:妲�V���٬��$_K��̢�9G�ش��z�y/<P��{�W�(j�mv�gP�ܫk���C�*�pr�m�rj8(�Uǰ��7W����O�U���Pi��<7e��|��v
s��^k���R���d�8�^�0��)󞺓�y���$�F]Y쬠����e1K���ֈ�c�W��6:�{��d������w��ړ�x��|K�q�{��P-.F�̐��f���	V�l�'o�IK��\'^��w&���s(����E�|�������FHԺN��#����Nk�~�.0�N�����X>Ş5E�t_O�
ܙBb���\w��l�ݣ�c��#�]K�}յ=B�v"r�r�~K��ĩ�dݚ��{=�K&楌�o�gHeW���ϔ��b���~��c��2��m���{��S�5�V���ʎV���>9e񘋜�+R�5� g(MvO�z��ƨ�g�:��{�o\о��G9�U��rT5��j'�8k�/��V\v(dp�D�6֦z��6�s��^g�L�;��ھ����ٔ���2G�v΅R�&�KC��}�/<�ޢ|^\�����50{rs�
�oS�\����ᢾ�wKO�~VK�r�\T�#;���c%=��\��{���{�B��Z���� Q�P���l&�wm�Y�)�]N�w�$�� @����
GOb�x]��R�=��ǥ/3_K@oU�6�H����	��{OSϣ��Gfs�-����[yx���z
w�ˬSz/�פP8/tZli��.���g�t��G~�K��=B$��=�k׭Dn�s ҭ�P[W��Iy:Y�Wɽyu���f�1�d����b�@+�w��[��#69"+^���Tsl�k�+3�Y�B��޾�6���c����� v�L8q�z�f�.ϩ-�H�rl߾y-�y^��q�v2Tj���5�C莟V�h����Ȱ0[�;Ӳ���̝��
>p�͜w�ڿL�V=��g��r6]u�B�)e��x�G�!����ڨP��Rڠ{ڵ�������+�H�ǻ�K��u���	�M����Yl����}��W)9��s�:�d����PN�_�b�B���{>�ap>ӕ@5��lX��%�i__wuF@�]�T�OI�[2C��|\b�>���S\���`�y(J��3T�OU���}(Ln��/̮9���]Pn�6ı�����v��36�t�ɩ'��)��*��u�0���_zX��R��X�M�g����>���=9�۞�{�3v*`tGt��Q��{W�%#;�&�ԗg�՗e��:������1+'�����H6���ktT�%�@�u"�3�x�v͢����x�"�uDn͋����5_�f�A�Z ��~xFWV=��{�e��c��}ng��}ߪFW��||=�ܤ}_�A;?�N�D���Ov��A��SB���3۳(H�$�����9j�������#�I&�d���T�0���R�FV;c�wz������7~Ī�d��g&�i��s�Rrei�m�q�m�Shn
_��-����J۳�C�n�u���{qr�+Q0K�#��X����vZ�n�Wi3ذ�ʎ�����Vq�j�9��^;=�}�8�e�>=�۳Qީ��O���=��倫���}s�y�{��u�˾\��[׆��N�N��vo�	:��3kc��g����ʻ5�)ꉩ��)�;r�1n@X�qU;/K�9�g*=Vv�,V׺�w����z�o����'�C��k������5%��j����*<��GL�����j��Y;��h���y=�˸���Y�m��K�Ne��ǮR����zu�QZ_>��c��wm���;<�(Tm��9�Σ�ܧ����Ϟ�߹K&�n�e���8� ��;�u�ݬ�f���C6��P���u�^���:��]>���>�����)�=�/GO��<;��4���Ů«�4�DyP�j'U�/�ǽ�=��;ꅆ���P�#�I�>�Uu��*7����[��.� p�;����*�a�}�پŃ#S���'���cwݣ���I�:��og�s��j����-!�v�=��_a�XP�.瑘���]�y�+�Y���[�����g�k��G�B���k��.��6iV�)H_J���Z枷W0���#������]Y�vwm�>��+�sAC�@ �K$%Iר��M�c`�x��\:ٵB�����6�w&�RQO{�H,��b��Z̚9��ٮ�`��������9�t��[2^�G%Cj v�)J�U��x�3�C�u���w��]�7:�n\��=W2Q����<�~�a�����b���֊ce-�O�ۊ�!#�*�{ޅ��;[�9#ޚ��ne��薍k]e}Τ]}�'�	��JFc����|J���..~�ίO�h_c;���z͎�un�F&.b�hp�]u��*�5\Vy�D᯹�ׇo�Ed�u�N���bdQ~s3!no���/Y����V��-bb�S��7g�����Z�͞�ښ~>u~���^jʾ�辛ĳ.9L��*&��6k�/�ڹ`��c �c�x�z�D�ۙ؞��[4]Q��>Q}uc=�l��雲99����ė��Yp6���t��������n�v����'�p����:��\�w�f��G�/җ�E}-��Ǽ��u<�����g��P+2�|�K��]R�m�9��.�,�������aR͇y������:36}~<��ٺ=}���^x��"/�(y�0�!��垎�Q��Szc�R,�rd�{K
} ]Tͩ'E@�	��tU��D�&�~����ө�ǆ
�TD:��K�ߡ�t���:w"d}�%�NI����S��\:���*L9�voXm@��s�����6�Ru��7ob+Q��f����Ǔzs@K��b^���Z�gU�@9�	��SgL?��� ���Nx�tk�#4��T&���x�;�
�k������bo�&���v3��5�@��L8�h
6��N��*�Q;6&9�7m����p�У�Sv��-��۪�!�.�¯��O*�@kȍ7�y0'�����}�VONa�u�������ߤy�go�,��^�$ZjY]fQb��u'�������'�(د:=}o�l��̥TF{�����ٓzj#RxK>���/���>�|��#P�d���3Cj rЁ�������W�Rs��sf�h��]�b=h�1�2�Lf>�Ϛ];��\Ot� N����-�#�*2��[=�aƭ���r�öCz<������[�(LEc��Wͮ;�F1�~�YV�&�N���h�3#��M9��D<�T��M�A��̖,Z�Ǿ�Sf��t�U}sC�.���+��~�9Z�M]�N߫�3�X�Ew/$���V��Qޛ��R]�f��6�1q�u���3K�KC��Y뭽�L
�x������漊�a֮lJ�L�I|M��.}���\��g��鮿xb��Rv=MO��)��M�&i.��ެ꽹:� O��RϪI{+e��}���Pi�v�=W y��9uj"��͢88���R��籺stQ�Zɺ���O�.�%ԥ�	�n܈�H��Y5e�4<�O]*ܑ�i5VJ�Ӷ�辋*�	��Gt��١�}7guܫ7�2G�v΄�����h��<�롹H{���oZ�Ӡ(�nT�`g�]>>��x^[���]��it|K���ض�g���v���-2a{mפW�Y=���jp��v�H{_[�Dy�T%��Z��ݶ�f�}ޙ�{w��3ϊX%t�o�/^��$�DZ��5�r���ҙ[��4mE�П7,*w<�zN��q�j�s�Iܜb�������8j;�$�ja��X�/�IL<5�����/f�ǹ6ow����+�X��g��WJ3g��e��O���a^%ל�֕GT�':�Bӳ_IL�X7=�P:z5���v<��;�W���ۨ�ꎹ#��i���<r<�.[u��T,�ʗ�/�^�R���E���������v��-]��;��[=d��a_}=T�f���G����U�%���K�����f�ap9�<@u���ϗ3�����ꌁP��P�*�zk���<�Xj��I��ײ��� h���BW��mߞ�ּ������צ�R������m�����6��66�����lcmlm����1��6�뱶�6����co��6����co�lm�����6����v6�������[lcm��m����lm������co���co���co��6������`6���cm�m��b��L����hYt� � ���fO� Ēw�z�$ U	((  P  �J$��� AI
�(�E � P� B�@���J��UEU$T
{aB@�J��@(
U$D��RR�H��D�EUP
 R��H��
V��% ���"EJR�P$��)*T P	H�IB�IW�UP�'�J�"P��T���	)J�:Њ�5J���H�TH   ������ڃE��gv���'l��S��屭K��Wk��r�tV���Y\r΍il4�:t[k��
�ݸ�UT���!RD�*J�W�   ��QC��V]�4��&�QEQEq��(���.ox�PQG��(QEQEuۆ�  ܦ�(�Ѣ���=;�QEQEZ�+�w��RE֐u�A�	"�  7z��tv���v�ws��t�p;���n�ݬ��;��m��.S���[�֮8�m����n�m�nSƳ�u�Ѻٲ���-��i���5ػw!����%B����)�  &����gZ�w%�ۙ.���k,�9�9�V��]+N�8�S�uͷ*Y���`ݹ�N�d����Jh٧&��hi������ʌ�m�v����6�P���(ER�Q(��  �xG��i�grs��khZŸ�w"��V��]k�9;�tv.Kw]��r�N�l5����V���X廮��+v�p��h�ӻ���rt��h�7�5*���hJA((��  nyz���㶛7+Uq���8K�-ݧ]wv����Z��Fݵd�5mt��u۫���K�J���Vr�]�v�j���Ϋm���V�5�vWwn�ӷ(�(B�fEH��� ����Gv�-9.�WY�h�S+v6˻r�wGkl+�Xӻm:��m�eN�]n��Wu�8;X�[wr��L�j�v�T���m�Un�l�;VVۻ�@�%H��TIM��  ���mv�n�۵&���:�mKn���gw-�K::ͷi��k�읻m�P9�r�tݻfu�M6mI�];�k:�7:�.m;�u��#�e����:�(�@T�	(�-�  �-Y��z���ݮ]����[uW*��mf�]$�r�'Y��m��n�	���\�t�w]���Y����i�M�wm�����Us��C�\���UU����o    ��ݺ�ghM����Mk��,e�Y�q�a�I��ttsfΗ��Wl��w]��t�Z�p�
����"zR���d �{FR�� Щ�3
�  ���*��A�!���UT�P  &�M&ʪz�`�FOh;;�D� q��8%��B����N�'�w￿c������!$ I9��BH@�h�		�BH@�����$��$�	"I��������nj��{]2�Z��cFX�t�6�֎���Z����t���iĳ�h��)�ki��K@P�2��a�[��!EZ��tss@lfӢ�eKx���B�f`4�e����4���u���.��^�GkKd��X�ʲNa��N
Ln�ц��c`���yw��Ji�"-ڨ䰓��Y71�aj�^�oma�!�+H�J��H] ���'|KTtm�`c�Ծ厬�Z����e�����4�l2� [;��Tu��oi����8 n��ح�
c��,�t�j�1���wcmSd�ޭ���N�ߩl�g6��l�!�/�G5X�YY�B8�lCJ�*]+�U��!Y�e��f6T��I��L}{��X�8��ln[��^�
 e�.[���ű�̂,�e�9������ڙz����Zl�{�4�����t�Vӵtҥ�Q&d��BAB�j§Xͧ0�N�����9X{%�K-�N+�\
�x0�[�6cұEk-9�>5�vpi��G-`�4NDUֆ[��ƽ�\.ڦ��ӳg6P��g7*R]�]u,V]�V�-�؞*��YY����Zn��p��� ���\��ˬ
ő���=��/J!U�8%ӳG1��tv3��w�*׋**Q�.�m�+���0wF���ZVV��._�(
TmSS 0�ًI��:�ۥ���M�gq�m�O.ӌ*h������;��&��G5V�kԐ���ܱ�As���1I�8n�J��Mp꽻ok`�ҥ)��n���6ح�v~YLV�aإ�5{�@kS�1�Xe:��u��s�*a�vt2 ��������ݽi�U�u�PF� ����n�˧݋Zl�6�]��Z�V���N�� XU��4`7��n�ݱ7fa�{���6���t�Ҍ=m�ho�����c�v�e�������׷,��њ�<�t�Y>ݭ��e*?��z"��Zax(�,J��e�X�r�r�a��l2fm�oA*�^ۙ#Ѥ5x�+M+u���h<ɻK\����j�xU3����^�<�ku�,u���:"��~(Z�D��Z�"��f!n�^�0&��ⶎ+��5+�j��Ssu͛B�ɕ2�@U�hjl"���bYܙ����sT�j�ͼ����,�n��[W�">�s6�dw6n:�Kn;%�>��p���]���&G�Mu�Z��n�K)i_dbT�q�wv��QE�n�0��t���e��sEdk2�[�u�����[zY��DՆ W�J�j<�ym�-�X��ܕ��T��H;Ib�X�^�)e^a���Yv��z��Y6�IN���;��,�����w"[>/4���sX�5��K+f	Z��I�-GW5�]]�K;z@�/*�Um��%@�V�Nս�#��'{y`Q�4�˥�{X����]ָ7�6���@ה����CUK�+����P�m0+1�sv����U�I5��ʱBB�.�1�M9��Hu'w/�1{Ckoic;b�LNSAUdwrQwz���.�ͥL�f�˵�[��R`+��p�6݌71
.ޤ�Ud����U���j�kD@*�6E�wQ�N�(ְ�n�E�gF9:�/v��;K��z�����H�I4�ި"�OD�r˹4*S�_�mV�赺+1=�ʘN^���M�l1ge����F�=vw\��V��d�t�|G"��懧B[������ʖsE���9EZVn���FH��n�M�30m�7�:"�L��Fˍ^A��	�̀�G*\˱Aqb8�����Ȃ����P��Sh^H�3Elq��n�<�A���M�"��7>�����&��Cuaoc$�X�$W��ֵ�A�5y0��%�B��l^R����F^�a,5�hmih�asL�"^f2T:�����gJ3^ࣗܭQ�4��D��޽m�6m� ����� F�T?jy���Wp�׍������=s(�H��ցEX*s V�H�m��J��iZ��3�b�g^Qa&���-�=� ���,�� c��u��:����+��X��H̏Wfݔ�	�Z��ؒ	�n��ED�je�rt��x��l�p���u#��w��)X&bnnI�s6YM�Vs�CA$rtel�v^��Pu@$��`4�v�ww{�b�&U��:�cј�0M����.'Z��ӈ�x>�u(���L�����=�����9lY:O�p�� �F̳�b��k���L5�pe;�H�r�[�r�;KVij�Z���
�uMө�˖V2�Vm��[VAe�#�!.m�C�)���(3fT�X�\W�[�d!�c�w�C(��n\g0����N�[ZSy�� ����*�^��ݰɀ��ิ3*��w���˵�e��yu�� 5��VU�������G*�v�`����2wҮ�p�֪���)�lz��b5w2C�٫�B(e��Yn�ل�Z,0�1�1hĵSA�U-3,&�A���'�2�bݢYzqK^}Xr��]�H�U��J_j}G��J�ap��Z̅�1�tY/2��5%3*�ou)M��
%"R�`YJ�(�yA2�!�b�23Pr��\�Q^���-�;2�emvQ�]�r-����>���=���c4u���"j�0�n����������ai���f-Xuh=���}��	���e^�X�
�`ΰi(]��Jk��[i��-U�vPei��&Y&�]��� lA++�J���<���&�J�,
�o|�{`2̈́���h��x-ػJ�����ݲ��JR(�2G�j��%K���m�U��Sm�7X�zfbҷ`M�:�Q)�B���MWCp�zH�S⨗wz��1�ba���V�X�j�.�uvS"0���N-�<�m���777첐�if֒OGeic�ʽ�J�vHb�$+�0���u���8{ww{Mմ�k�X��R�CÛC�hr��5�yW+-4Z���D�ʫȞ�.�*�.���I�U蹳dҨ�aF�cM�2[�̷�³[����1,�ӎ� ��Ǔ�4D�)�e�Cmu��m!i}�lg+��n����c�r`��f:SI֍m�yV;@T�=��[���g&\�/T���</"�	
�+�c`]'�feU��v2�<.CW���mn[;	϶�]�q�B{�e�d�Xo�nْ��b���[Xt��y]��!\�_$�Z����	��{�{h���u����v�)MU�J�_>F^��h���[`�� ���Ǐxc�D>�9.�Ѿ�wh�(j���1.�)��t�Vmh$^��B�ɚ%�fP���{��	��Zh;�N�Hfk��C��(�U��ֺX��憲�T%��yX$��V��ݫ;��,�F���;"�J�Eޒ��P�r�s�s0J�f�cF�:H5��7wN�U���Jr��V�F�$��V/0S�k߈V��2�%	M�%�hD����V�2!�,��b۔66rc�E+�Pѱ�V0��#���]��W2��kE�!Y*n2j̰H��e8%����ɰc�N!hej%�&>պ�j!Cq;�[PTӕ����q�wG.d��#"�Fۓ�"��2�:$�N!�s�4m�1��U���hr�m��7��Q�I����Su}r�ñA���(^�X
�XAۉ�z�'�ҕ��f�Ŧ�x�@uW�Ǣ=$Lٚ�����1�q��6�]����}��ӻ[:��|��V��
���ek�ÏH�Cd�������3Vi�1�M#+Jf����́���&78i���F���E��P+r�w�z���ھ� �0liB��rP�ω���8���cP�t�	�Y�Y�}��p&o6��(]�:�n�t�!2�׵rL�h��Ws.i-�GךPۛW�1�9��v����4o+r�ڶ�R���Kh�Tu�jG0��^����e,�N�,��}���,L�,�wj*�����$XfFN�ږ]'IA<���L3Xʹ/a6�[����o/w�8��*�\�K���эlĮ�:�n�<H��+�[1����@6�j�6���[���C]�iV$�sɢ�G[7RQ��Y;�F"P����փ7;�閇r�n��kPz��M�dL�"���u�n�e�ub�����3��ka۬5Wz�a����=���:�e-�zL;j���� n�-)�1��t��K0��,`�j�7(��v�y�-0~�[V��H��gb-԰]�u�'��������mv���Ȯ kn�	���1�CwL�b,v>���[�dL#n��[������ư)��{ylZ��K:f<-��th�th�soqMa�VQ�;�2�ɥ���n�3u�&���*�n"m
wq,�bI^�+�ՙ+b��XS6��5y� �G�`ڻ[�C��4�fSȷ2�^0�j��	�Z�%6��Hh*lP��V��{@�����:�
�	���Vh�_Dƺ̫���.�47�U�McE���]t������`*��mK���;ٵ��^ݣ�,�m��NS+!6�*V��]�{Jp]\8u�'V ��.�l$�e��]
���d�hVms""���ΚTM-��`��K6V)�G�[�B���׽�3�]�\:O:/��5��vq'X��Z�G��u�)�(�T�ݵV2�AQ��@��3i��˟��&qY�(jh�2X�XoDim�b:mcת��Cv�6��OF��
��;�pś��ڣ�a ����Z�o�N0w���u �<f�/u�8)V�M�ϑ�9�T�wmAv��C.�`;�bժe��ݢ��r���D��*��v����i�*�M�	�Χ��6� �)�W��������]\���!���W����U�ʷ��[.�#jîgWah*:�:��id�A��.=ѵ1#��ɢ<�ڐ+��Z�]��V��Z)�\��U���CX�X��+E�������z0��N�ݼe�d�e��T�*;���n��`�J�!�ވɶI���;u�v�7Jn7,�����U�j7�F(�͠ ߋ��rJ��@��2��V�c�9�k��C
��E�o�@Imh"3tS���q��2��ʺ2���۰�Y!���h,Z���jGI"�$���a��2�����Ԯ�8���p\�Z8z��q����qXN���2�����FS5&V�7L�fl��ܒӺ
�C6���ի
��Y��YJ�N�ʯ^�	����5�J�%iW�����:I��m����sPpPWѼ7sҭF2�3Bٷ��k�qVQ�׺+�V�1�w����jV��]���JD%�[��i�\r�Kٍ�\��ն�GB��k$��Eõ�9[�E�^Zy/��?]`�qlBV�a�w����	ת���ӛ3&�i:�S]�j��ksY@^V��1�R�Vb��e;d4Y7v2�Hi�z���rh���oXz��PW��@�u�m���.��c��&�z�ܲњ_e�9ɱ�s4��-F�H�Wx؈�\L7+���#.��3V���T��U��B+5b
ө�͹w�t������V.����-�7Yj�7��@�P;��Ů!���ؚ�G���sZ�w��ީ�*�@qP��I���eՋ�QV��(R��7�� �ɢBH�T��e �Z�"�����jQM�Wx���b�n�/v��U����6�F⭍:�ԥ����՝v����V,�O	w�w�TÕ����������l	�� K
��R��V�9J����۷vՍ��^���f�aL�O�Z�Y�e],'�F�Մr��r�hc����
�8m��p�ݘ�D�[R����k�:�c%��-�6���� MPe]�����6��i�<Oy:�Y���� 2��5�Rel�0�`��։�eˬdd�T���^P��K,��$yNC��Jx&�v&�ۛp
�;2Xʰ�/@4h��ыk+x)�)��W���2�Ҋ��ѻ���&��U�j��C2��J�M��׆�]��̹T��*}/S�<�Qe+1�$�����Z�ZM$ۢHô��6������W����FN
�b+�jŶ�qR#h:IO� 	��}Y��RlU�ɚZAܠ��D��t.�iH�`�v�ӊ�Tɧ�Kn	j�6����nQ9d�i�r�^+p�sv�Ů�f0����#�ѷ�ڟ׫f��.�
��&��`*oD`��+��2�	f�˹�7@��c�YFi�ҭ����Ll�d�$Ub�ϱǯ��ñI)1R\(h�(\�v����������ۢP�WZwS��)�@@���i� V���(E�7��5MX�Qe�ZF���;Z��:�R�Q����nb�mT*�Nʘ)�8 N�PX��*�*�
��f*T��6iȘ�O%�tT/(���ʄr^	�h{�&HC{���A`L��dj�u�][����eZۘ]�[�Cp��q�*���b`Yr�A[�/+h̭���2�-Q�쭗&����b��P���bf��3�D�n,B�K"�/��Jn3W� ��ү�ٓiGz�
��Y2f�ͻ���ks`��F��� �iV[�tJ��X,e��!�՗n��[mTI�#�w(�Qj��8���3W����������0R��^�������'\/�5�Q�O�-'�lx�����YG6^����l�VcNfRm+B�M���ٓ+-�OP�� 4�xXkYݸ^�$�M8��P�oT�ֹ��X�0�m�Zض-�Q�޷��3E�(Dѭ������������k=����ҹ�V�
[Ǌ�d���9]�mAp-3�Bƻ|w�'��dӔ7]�[ڝ�[�3wALM�!z
�Mn�՛Sm�ȹ�����3&��d�3�\D�}��{���he�r�c+:�w��`����$�ܓ�fP%���Y����`Rv�x�L{Kx�7�D8iۣ�|�4/oUvA���������͎Y�t�8:�=O
t�z;X�ˊs��{!}�Q�6>�oX܏��!��v�b��:�u%�:-`��l�ha���3�VC���Gτ9�At���άo���{1���X]ӐB����o*�{��G`ȯ��\���b�4�fv^�6XF_v,)��R���d�Zoiڷ����tU��a���1գ��뤰#C���jQ�#��7E$�*�pݽ�/(ӍH�!͌*Hq�o�� �AR^�t��%�/���F��Ē0��Yx	�0KR�[�WO8C��U���&��Tn*���1��v�sR���8����'N�$��jTAI��(]�u0�Q��f�eH��2��s+v<�8�����Lͣ��N�\�P����4ַ!ޢ�ѦM-��sSKܧ���N��=
��t�ݮzV�<i��vz����]�-�gd�MX���U�XW}%wP�����.�o�\��cKJ���Z;�sh�-�Ts����H;+��kP�t���xt����CXw-�	�{l8��!*�L�b�bJz7K��>��D���2,QՏ� ��R�R����J���mTLo��\ˬ�Wn�;�¸��]�4�b,�=ʭ���F�G2�p�Q�7��w#� WfK���j��z��}m�`L�_�n�ۘ]n|R7���,kn��|�uI[�gJ��]��Ko�]�7�mw|hC �����36N�w^]iqu�[iN����謺ONc��]Gb�F��`��=*��W22�3��(f�KD��#�.<6=�q/���G]��n�Ŝ�J܍7Wo�J�ՠ�wYc���a�f�G�t� �ݦ��i�5�E�Ӊ����U�4aE'񕤼8xI��$�ҋǉ�j�VL���|Aݬ���w*q�{_]�P��{�yQaP���,����鵓U�4��m!�ܶ�!�P��gv-St�n�uN7]>���MbsMBv�c�v6�e٨X:�nݶ5�h?\Z�')�6�6���m�t�(.�;��X�Q��7qi���ͮ�)�C^��/����Tb�*�y�gr��^dw���-���*qY\�L�{�+�W^�W�k���%�ˈ��P���]O1�{�H�:s�Z���G��°���s�kW��g�A�V��� 6'�+�Ռ���l���U��3t��rD��6m:zr����ޢ�l������VI�G�f�m}�n�6�t���E�-j5g��Oo0��9[�d�N����Ǩ�2�
B�Z]][Nr��l5�1�u��3�=%4�D�6�Y0a���o�!jp�rH�-Ixv�.$^򴬭@e��j�R�]+�*h�e4�7[N�4.�"A�� ���J�˗�V=�w-�r�5>]gu�E
��e"��;2]&�+D1�P}w]��{a)u'*�cslU��\�(Y�1Pܾiך��`�sZ��5A5�V�x8��ht���ŲS�X._=b��қ��M*Q"�� 6�jӸ��,w��WQ�r�V�e�7e�odH;�H�F��}�z�Ĕ�ZΒh=1>{��E��� ��p��������-vj�j�xbt��R��Y�ۀ=9���q�s�O*�w{��]��ﶹ�Z��'i�������[�4���.��Jfo �;���d&Q��;;�D��Bn_1S�MꙒ�eA�޾5jUg:P��ۍ\;rS�!Mz1!:vaΡ��}�]�"�Yv��ײiL���Z�l���F6�*8���0�A���k�[�W�v��<s	 ���
��Y�)���Ж���mf��N�kO�gR��&)�v����Y0sD�\�R��f��R�\��{3I����2��L^�:�˻��n ���c]�V,�4<�DZb7ND�\�Vd[Pڊ��$�.���9S�*���4������c-�Ǫ���c��8W:���oo_;X��)�4]�1T�+{���Nnb���nݘ�FV֛.��]M��g`'�KHȱ�t��F�}����%[\����l��mEG\��sV�˸yJf,��.{a�`�}[��������
b����N�
����;8��a闖8�y��� Ӽҋx��+���`�sS<��[���%on���W������7��jF��kw��z#�A��ۗ�;i��zy�ː*�%Ip�YR��KwpTX�b��n�]�8"�J��W.���'vA�p�φ�{�Սڜ*o�"��uk�j�
�أ
���A2��n�Ac�Ϻ�<EV�$�V��NW�����`Q�G�7_|���@�Yr^��P���]hQDuMH�R}�lW�M�m$,���o*�+�5x������X-,Y$���2���jf��\���wZYԲ��X��tc�z��6�]7.κ�	A��kW+8l4:�	�C��ư�5�Ԏ�S�@j72����,받|GwVA�Lc;`���(���v�
��6��+3���J�߯�#�	�P�բ�f� t�,ne˝���3:��B���Y�fR]GU="������;H�-]�kswRT�X�<�q�u����Z�m�{�Vq\Ӏ1aV�έM��k᪮���U�z�e�7�)�*�Sj����S^\&k���[�4i�M3�k�2�x�e��E�Y��i\�4%�b����8�)I�Ժ[��)�i��DN-|�7/f����W	
}����q󩛷F��~��r�M����:�mbbR��K���
�]d��SC	5\;�=krYU�ҧ�L�깘�OP{�`�qHr*�O2�T*�ޙM�96��K�/��Өf��w��f�+S���v)���+f�\�Yu+{��d ��5I}g-�󺚍wm!t��Yy��<�>{-N��e#��]*��C��WZ%>f�W���ݓ`4��\� ŀ%u��q�Q��w+��IB�jSX�ʜ��IN�.���Ww�i��ɜ��9]�԰��=�ǅp��4����ag ��`6;3��=�<�|ھ�*�2�B��V�D�*:(P��J<��8�H��ilJR���l�)f��q�l�"Y�j�3����0F�5���:v�Im,1.f����}AǕ{޿�7)�־�5q5 ��.��1B��Ʀɮ��hX)��MP��MR�B�����K_m��m�@�3/2����c7�D+1&�����`��\[3$a���)���yg�%l2V]�Z�J��8�u[��T�Ǐ_T�x��<stȝ8�;�p�ei�+y%K��ɓ�A!��EW���"�{�o��uc[��b�]���k�a9����(��p֨p����w];A1W�yP1R���#w�S6�.��H:�NF�k7��G�xI�HPWv�׈05ժ�'#�F?�ohye�5��c�rc��0��,u�횻'E$Xk��u=����+ �&.dp��*��9�����h	�n9��2CМƍ�ی��+D��75�8��c+YR��V��P��c�g\��K�b�����:.|�GOt�mE���4u`�:��[��ȘJ<b��J4	M��}��T�f��[YZ�ΐw��P�����r+f���`���o+uJɘUʟKk��l�:��w�]���HP|�[Xz{E���F��4o)��u�w��ˆ�^� �w6�-�x'��O>����e��I��Mp{e�\��y��ک7԰w+����lQ�wh>�%X��yq�v����L�+���@�`�J�'��m��2赚"#Z��em��zʹ8�+7b"�Aw�u2����Z�C���ItƼՃ
�b�:��������6G��y�!�ǎ����7$�F���V)!h��%��n�c��4vb�Z'gv�C��v�=[��*@�v]k�����������2�1-ޕDtpF)o/��G'=�ȉ�]���"-��4wNTz����#Se,	*#M��{���5ԗ�ҁ�&u��;�f�I�բl��1G�h�+i�۹@�5�ﴹ��U��Z��y���8�c
Am��b�M&��+��tv�,gq�ڴ.�4(Fu�)7���/����iVtP�mp�ܒ@�ś��v�P ��'�r�j��� 9��w\+�B�Z��k �,(̷m��=�`�W8],tҮ0�ܒ�v�;�0��D����*R����v�GF�L�ɵ6�rM
��7��uk6LH$�۳^d�ξ�V�+:�%or5c0�G;D۷Y�<�^���Q�(�����-3|L�M8�[Tyl�U��/�mA�>���9����d�R������G�ܲ���kZ���6�{'[Wg�����E�(��'r�Hb�y1"�M�|����ha��K����R�$}�@)�.S�c����fBonF7�#�|P��&T�)f��ed�]�f�f-S᣻���74U���$��͓�n�;/�kp:���f��0ۼOV���ur�ieD\��^�{��C�fM� �K�B�<:�����6�j�nް�k����\�􈱎�hToq�̰��3&E��Z����P��u��C\�����8��$���^�+7�\�����o:������,F\Ű�m\]"R�ޮ�hPF�۠�����/���GG��$�i9�M��<�AN4w+�q������ɱ0�vf��\�ڈ�x)WO��}��X1�W�%�7o��	��VZ���I������8�uI��q��*�2��)�]-d��AGr�Ϩ^��a����	={�N��I;�^)�fb�)A�$#�rc\�!�*�ݸ�b���'C��'{��ךh!���Muf9��B�rɯ*k5�k�']�ڴU%d>9w�I��"�P<���9t��żv�o�Ԅ>��������WO�X{B��zS$�ͬ��oQ�ͮT4lͩ �[�5�sW0c�n>�Տ�IL��[r���G�D���U�(Z֦}��0X+U*�����T��1a�{A�O0��g�S��1�c+�W�u4���b�R�ܼO|jy+ �X2��P�Z��,�n��s���̸Z��/�UEj�̣��MK�k�6���>�Fك��:EV9�#��R56���h���[��ki�v���g[T�pn��$�d�r�_���=��%y6JK���¨��ו9��]�#��E<g	%>��:��꺬i=��i<�Sul�:P�p��r��=��n5��Wbg��[��^s+E0T�Vgj�����-N�=�8�G���̙�G�	څ��k���qB�(f�x�Y7�n6B��:)���NX�*�CJ7Ȼ[˱Ƕ������#��N!Tr�6��G�����f�ҭ��QN�c��� �wq�)�O$���9�+��e�Fµ%,S�LێQ3X�w��*��g>�M��V6m7j�빓I��]�����X;�zb��*��u�\�}+T�V��Yn7���7w�Z�efe�&�L� Y�h�l��v��%�V飽&ޢ#�-�[\�/K�OuvAb��5�_JOe����%��{�ʚ$E�r�J�m���P+r�	W�R@�о'd�ova"7����GظL�W����$��x+�Ս�a��,I҃�E�tAQ��̙/&�{P���;a3o��|�
P��ehi-��#�(�8�+^�w�{WeŔ_^V"�up�﯊��s��7|y��^s7���V��-a��)5׷}�W�3����3WɧY:MY��h�	�%e[��
��k{~�+���݄p��vd�=u|�����ʓ���q�˧�-�6Ukyӥ���wlv"[���@]�㋩���v��B�m8f�B\��_]K���y�-uCǢ�,` �ᢎ��L��
�[yY�Qs����Dʌ7T=�k��v�����љi�:�N��N	E�gZ�$i�-I�um�<���Yf�4�����Uܣ ��˖�p�ݱ
t4)l
�������
�saNJ�4�G3yV���E� V�7���sn�nS�p�F�V'QK�|�7�EK�u��#�OX{5XYcP���w�ܥX`����`���G��rf�W�L#�c�m�r�bN��*�rd��H����u��k�ԣ�|�ގ�r'gy�젳Q:1�Y��J����-��F�Jf�M7}�f�iH��W�Wv�����C#��N�ѵ@cY���6�q��al�����K.�nVj\{kR�8�B<�j^��u����m
�q{Ը�(GJ=%��U��]V�!�V%\����fC�V>���R�7�Ewi��v�E��|Μ�Z[�}7Pl�BT�,`+�}�5ӄL�N!<˴;m�z�F�2˹���@70&sv��[�e�v���Qt)6̹3���{-�d���[��gn⎀�rd�Bx |ˍ�+�:���Ua�[fs9ٜIʙ8K[�@J-M��&Ρ���U����H��{]G���2�_ho��^��v9{wP�Dv���e���}Ηȕ�Ჺ�H��N,q�"Ǡ��	h��w����5ȹ̼f�4TW��6��# �͊WM�gp���˼�-��:�z\����-����W����f���j�%M�ܫ��b*I�v����u:��ι)�K�(��ݽ0hM٤ԥ>�tg�lZ���4~ҥ�㲱Pa�ձ��AqR9��CJ\�e꒮1v�Q��,+�ZB�e�w��L��&޹{��wI���! ����$���~����7�5y���d���+l�m͖��ø��!Ij�j��DoR�L� Y����%.�y݂C`]��N��/a���iqT�6�SB;ߋU����=e�{LV���%��� �kvX�|�!s�T�]i�V�s����A��;�M��y����:�`�����1���æ�AL�Ǻ�%_e��Q�ӂ+ �Ǹ nrTf�DʝĶ��̲�F��9,�������-Se�OnP�<+hX�_k��d�(��o.
�$+T�h��r�A[�)��|�i�wwx-��ۊ��$,&��)�K2�h�y�ګ��q�l����;���[��v�I���X���Y�&��2G�9�94l}1��L�z�}N�4�6u�3���q�^�x�s��)S�C��ΞA^���(�}� ��V��g=2�%� `w�$e
�(�{o��#YF�X��]=׿wv�m�v�Ō��w��\iU��"(�m��+��%on[��Ԓз���܏is�R��3.�f_i��U��٪2���\�L1֮�o
�{����*S�L�/��@cb�Σ»5e��Ĥ�T��IM]+(Y�9��(�q̷���H�����.���iӢiAw��a�(�����uon仍MɎ�"��Ю�쮶Grs���м@ma�}c��gt
e��.ޭ��yְ .")p]��|k/O\��S+�ne�$��p{�o���!u�M�/��z��}�EM��`:2^੥�
C���kx��]�5]�p���.��@�=ID�aeN�M�]k-��M��}��u���U��:���9ͦ6Qx�)��<
��T���׏*]��؉#r��ݰ���є�ڴ;.s^s�udy�˦2���"��C��zF�W-�k1���Z���X��CkQŔʰj�Ɨr������Xnf�v�]��s�:kkD��AV���+�o���9����rLv�>������]M+�ɰL��K{��mt�f;ǭ	7�.�S�$�]ӎ�j�B��ANo7����W
�Jl�u��5��[:6ᔏ<ܻ՚$�o
i�����.+��7n�"T���*5��n��o۫滇^�&)�ҫ]X�kr�).��5���XQgR��u*�Nڋu��G����%�jck�ĭ�(aˤb���]�N
7��j�7]�����6�CYts��ΛXeő�*:87�fs5�C(��@m^S�Et�x�����\1\���&>oR���ɘ�3��Ո�7��js�M����4��j@㻝�]ښD�
��=�ކ��
�諗(�m��aϟڨh�lR�yn靰v�ȫ���:y,-�cQ�h�]�&v��]5N��3׽�D��ki޸U�a�ġ�M��]�5cX���J�;]M�
�f��vfvs��n�ޝ��I f���Y>H՝�h��F�&�1�2�lBxvZm]Txb3XKXܰf1�Ym���0�`�<��;�|�����!�j���;��'�-��������֒�en�\�z��3�雃�]\��&P��pì`��32Ż�.b<l*�}@�d(���5�5#���tw��F�eܭ[�*�⻷t��&�1�ұ�+���T��ڂ�F��JWnf�3:��mN"i�S,Y�:��j`���l�[��T�gN�U��2ڱ|��[�M�|���ڒ��
LS�z��e����!����b`E�άo �e�2�c��y����[׎1����c
�Y�l
��܇��s�b#�
&87C�<��L�:�؍�����!��ѱ��Mɽ-_�2�0 ;�S�˫���Cc�0U�[�ɾu{���u���(tO]rP.�q��5�ȝ1|�U�,��I�@�h�c.0aΑ����Yƪ�)��Ąh��o4�=��	m��s@�b�YD�' ���7R���o5��=��aEc�B-�'kJ�7�sq�y
�i��u2n�Е�4���|��^��i-��&�*��A�{�%֬g�����\��q�v���g�,��h��r��:�vĖ�W����)̸v�Ce$��T5�=�Q������.�f��s�����V:��C���q�l��j$[Y�LÌ�@t��b�n�S���P������u��݊18j�u�U��p��L��U�$�-lO/d�9�@��h5�Z�R���m��a#-ea'(Ki���a�6�<ߎ��Fo ���Z��n�M�_Y1
xL��J/v'ݖ1!Ő���q�G�'���z�[�2��e��󩋤1�a٬/�@��,�G\�5[��h��]��?��(�#�n^�&�W�

���ֻ��o�T�������+��,ˮ��:#�
n��dJ��lS$��[�U*!���Z��ђ�rm[F�M_v:��*�֜�IIS83V���v��a�/��K3��*�.<�l�c{k�*�r��.������j�,�ܬ�7:m�`
8���B����<_v�]�1i�*�\.�Js���ޘc�CG��Se���%:��P�}ҡ���D�P�h�V<ɍ���0�(]a�����y|��ne�����-�ph�m�ۈ�7A]�%H�fpt�ڷX��l��12 ]X��yu��Iv)�D�f�I)�{Q��9��v�Wl���/@b�;Mlm���nՋ�4�����N��wFN#s�d۔�:{�G�Wp������e��c�[�����iUٿ�#ך;L���[՗M��r��ޱL������64Q`�v�dj�p
����U�#�b_>X��t�omh�'n��1�κ��n����ղ��y�v.f`��&���60�_Ž�&۽���rD�C6SA��۳�x�9�̕}�,�.�Ss��7p��N	�[mq��*�9K�#6���h�uȯ 0�{ڧ�Yy�ˠ�iY�T+^���)��t� in�B�>�y� ��^۷j��as%upN�.@��E��J���
]QP"1�FC&rt�M�)�D���&V}�V�I���>�����x���qr�k퐀�6Ø`Yo�WG
��q=N�.�n[�vSZ�|*۵oB����R�H�����1V[f�9��u��b���U��r��W/Wƺ�NՑ'��뒮ܡ��;�.��w�Fo��M���v����'��Gg5ܬB�I�r��v�	�Ճ5iҞv�F���G����
�ع7�c0�y\Yܬ�WTHr=u�g P7���g	x�YFq�-ㄞ�\\}��V
����c����Œ�g>�zB���M��a�71�F:������`��j����\�+}�6y@B�Q���P;�[�\���:&m��\���֛�b�53-�ȆX�A�V������n3�O���:}��۪m:��V� ,�Q�w�,��5���x�eZ���N5+Zp���U��Y��x�f\����HK�x��C:�J��v+8*hI�$,��;��[�c��i�+�Z�x��j�k��3+E�,��r�)�0��W����U0�}�ʛ6�b6f��li׶8 Ӣ5�=����ù�O��ղm��=P�5x��?w:�9�(� +�m�D�^��R�¢�c���γB�-��ǹ��9[����ʒG�43��1m���o7�sy��A4m��Ӄh��en� r�(���VX��(u����� ��86�r��Xq�<�;A��!]��Lܽw!v]����=�[|������J.�\�p��`M��ˤ>#��,2��L�u�Ka_ى!�[6�9w��Gw�52��c�]���ۙD�ΒNgaEǨ�Lt�X���V�Ι�,]н���{Gs|�V�t����&J�(�ҁ'�R[j��	�;)A�01e���I=s�����6Z�i�2���6�]��)E*r(��Zs	ْ]s9X�M�-��ir�ǰ�}����@��:gV�ୠ�9�f����Ҕ}���TkF���
���V��L���sr�U�^�<���o��,��;��f�B�f$o���ٻ/Oer��.�U��%�'kq�(�,3t�wiVX�eݪ;	��O^o	�E*�SB]�p�!,��4VB�F���,U*b5�v+2`<�gui7:�;:�&VM)�ی�ַ���=OsZN�[��v��4�F��:�L�2��H�T�v�(�n;,-�"I�`{�n� ށb��&#�iك������?^�x�l�|x�89o�U��a��l�Z���Y�۬s7�l�MwF�S!��A�{{�n�}��5ɍ߱�@5���P���6��T�]L�N�[����B�����LݷG@���I�I$\įWw`�
j�0��k�'+m�ʇ��K�[����.�h��'p�U�	Ʋ������-D1Ź)ҫ����依)]���IL����Ȓ��i#fi��m�+qR�ʶ��ebܔ��IQ+� ]�b�Q<nE7 ,
�k7[��^cJގA����C˨�4�cU���O9��xsM��c�c9�5�Kv�T]����5۰�Cz��k�ɛd�-�Y��Y��njX���n�"��V�O-ӵ{x���Douy��ZC��|B��^e�fB.�Eչ&����3�c�Wu�mk���]��dAik��tY�tV�^��]vb���;u����XsGK���LG�31��kv.'W7c���j�E�������2i�7�XvqF)�2^]a��IpN���"���� J�����b�=���ȕ���樻FWH�wdZ�1b���7y��*I��ե��C@h�j����[#n���ŧN�Xtq8�fsZ���.��(� �N[��5��P�!xs%����/��tg
���q��x�ł\�jL
���R�j34��l]�5,�W���b㘋hȏv�/$�:��*�u�>�
*�a�4^7���te�<TϺ}�/��[��%�����YtT�KCx_cTv�З�4\љ���<�&�7n�@TЎ,-P�+P��S����iKh섩)v��!�b������q��a�d�Zfn䡔���)^��`�L']�!��bWv���ѯY*P�JB�����I�� ��S��/�gz���,�Aͱ�ZB��6ڻ9���l+��bgP�"-���s\�Y\����t�8#�/�T�R�Cل�{!��7)���i������e�*�G5r�o��W[�/�k�`
�=��U�{S�*�%gB�g	W}Q mR���9fLʼ��#{D��km�5��*�5���U��q����)1�++�^l5۽$`���#sk����f���W.T뷂�9`�"�wL�z}qfC́V����Y�%W�^���G�ˠ0��l�]�c':��R��4����^nH8��{�7(�yۦ_l��"�-K�;.�{Lu�����Dy۪�TYFK��u'�r��at�:��ŻZ��bj����Y	�\�/)��;����i�̕|؜�9�ׯM8MA�gx;��j=��^��k�E�&����컊�����/QW��p��:ws�,�Hƪ��+-�E����J/v�!�/��+���#�i�V�]�5��L[���xj�;�d��c��3�t[>꽖r�JA�����T	�c��k�72��܉�*}��j�k����Щ����}���ʚr�I�]��9ι�F����wB�riխ�GKyK#D{ԓJ.���ہ��EA�V+�S4�`5Ұ�NΕk�h����6K��+���<
�'��u�VX9�`�*-�1��z�(J�ҮK��w��BѼ]����]��i�/2<d[)]�EXHu��S�xf&E��N)YJw�^�,v*�q�����>6T�P�6�tC��k��lX��E]���3;� �T�4$�.�b�a�&����bI�+of��t5 �b�$zY����r���B[Yb���Ǔ�΋.��/)��\$� V�,=��9a��-!z�[��{��e�N��|Ĺ��W_���	��}��s&2�X��2���<�+r�t�����[]���*�QblU��n/���z�Z�h2�V�Р�x<�^��
�p�2b��a��-
�lB��.9ޤ�YE��9le�9LU�5_tF�m�Oq���(�K;��Y��P��j�8-M�Cm�����ie�Z��u����,h��i�b�<vWrWa@7J���yP���Q�lV�,U�3z�x_����3+ϴ�u���U���6J�%]6La��祽�<�ϸet�<�y�(2���{n�0��{b�F��j���S��Q|��=���4��Z9+���qn��x�0���S 5��%��bٮ��:�&!V����J_K���ئ����+�U�s�&�u� �֔��aYή�R�+�%�72����8��΅'stD&3)N�-�V�c�좀eѣB,PZ�q�{�M�{�-k@/�{&<[+tV���OgQ;��\��ݴP��r�q	�V��P���! ��P*�8"�v	�0idO��Аt�ܾz�Ԡ�
�Q�V6.������w;Z��	�8A[ۨ�� l
���b�&�l��g`��.c�f�W����2�Y2M����7>Պ�S�9/+�5xs�E���ʚC{U@��M����V"�1PB��X�ud<������#<��0ltY�����[0�ܤ�1���1[�V��3������g4-�OQ��J�}�d�]\�
T�,r<�w�;&�;�s���Y#r��r������,�����<ҍd3 �U�v�X�_��c=��yƞ�:t���f����ѵvP��z=�G�=�W�����5���ۢ�D)���N�r���y�O�F�!o]k��W���tR�%�vP�;iD@��;#��	ີ�0�����2�v�ѝ�B&�]Ԑi��� ������O�C#�mgnSb�	<L�Km0j���9�ԣ�����4���6��1���M����� �=gQy��#�6�K�s�i�oG(.1Q���$�ӝ.�t������s�c�L��Y��{�+�:
sH��3M�i���y�]N��{ko_NW��Nx&����g+iK��90a�"L��v�o���GF�-���Uy�6U�w�o<�fu'q�S�ײ�B�f�r����;ĝ��?t�*jKv���y��eD�W�t�]Ff�SV�t�r��gۑ��[}ɧsk�Rȁ�=Yf��H�噕����Pa����R]p��&�u����N�fKe�����lk��b�s���+M����\�;���|�w��>FS��y{jq�ю��9.�y�5��H�]�R�z�{������Sv�̋*�7��f�^�3�PK���cָ�fv2�0����z�o)��(��w�]��l��aa2���N]�N�)��T�D�;r���\k��	�+��L�Ƴ�9���fʹR����w3�*�w H%�WA��=s��d�Վndr*��$��� Q%��@�6��J4��X��Z�8屨ڭ�"-�T5s ��-�l�h�V6�Xե]&eX�R�(!V��*[kR�JRV���EmYF%�EV���dJZ��e�!��J�c��12��A)J��[m����UV����kl����f�Cᘕ)im�֨2��*�1EKF���
��0�V�"�kmm�����-��E1���f%UƢ��m�kXڭ
��,D�m��(�"�Z�Ub3T�:��j[Dij�eV"E-h�ETcMT���3*U�U-�ղ�QDkj��FQ*[h��� �M8`�jZ5UTDb*���F֭�DA��m�,Q�QE(�JA�Z-R�[*e�j���eՕ2�F+i(�J���b�J�"�+k3����J�lQ�kH�YR��j-)UQ�e��"���kA���(��Q�E������[j[UE��)h-�PD�Զ�%V�U�lZ"�����- �Z�(����UQDV$KJ�UF1-�DR҈)[-hX�UA<������wMW-t��5��nXC#��g.�r�گ8�k�-\���}A��ͼ�},�l�K��|n�E[3���f8�m��"X����A앜�?q��vy
��(7�a��I2U�u[+�=�tvf��^Y��.�@2s�t���1��&+xh��n��;\�f��]}5����+��_��2x)�N���$��X���-N���ސ=�r�F|=y�o��8ocv ���OnZ��A�vWX�N�fwR��,S��ـ�
�tq�J}��S�x��fL����wA�ln�7�v�=wYк0����a�)KT���c�wI�s�B�v�t7����_.	[��ON�#&����a��EOb��3Z�D��~EeZ�[�V����u���B�1��=�ϩ��O��:��[0P�9�>N�=��)��,���8�^r�s�q���<�GwL7���rܪ�0OVc�܍J���z���9�h��kQgʣ�+������_
b�k�6&�n�T�a��!�S�����Yf�X[�X��ޘ��(Vyޒí�X��btpV��/SyQo�KJ��G0w�TV5}�5krR����J\#u\��]jv��,F3{L������ʏ'+$��*�܏/��r�b���vw;{+;w��s�x�}�=9q̹��:�Ф�bkSy!~<�9j���AyM����I%s���r��-���eZ�S��w�R�c��
���`��3h�mc*�n.Y�ﻜ��"bf����j�c�{�'�R�%���p���iV�����9^j��T	>�=�OBHX��&��r��P]������O)���knR6i���U����S�&�]�ѩe�*j�M���ʮP+�V�>�yQ|z���>:}(׷���Sww'p1�m�3��U1��1K��4�,�ʂ«��i�����Փ*.��zI�����c{q*�ۛ���4�,��W��u�6��|�E���������i�B�a�_�{r��!�G�o��Rʃx���v�a�IsQ�wz��[�8,�{�^l�P;78��4z��$����X��;��|�*Js"�Z�_u�|��m��P�q��h{E�P�V����gV�i�J�2..nlȁ��ɬҫU�)�f8�]C{j�:� 0E�8���S;@l�H�x�Vsj|��K�L�znv��d���;�֨�J��Qj�_�e��q��Kq|��0��zv�����(�0���{�{��Cq���)x//�ze���[�n8m��f����g���__�ćf��ی�nlR5yj5�*����$�ӚvY7@����y�
��%�;���i��髏,�WNl��]*���f��-�.�pmjh�ɫ�=O�!��U�n�saluڒ�������o�^���Ok�I�TG-WҞc皽�Ҭ��Sjp�||����5��:���z�jq^E5�HiJ�꾕��L�|6=~_��m0�pʑ9w{b};�)k��Z}F�|2
kbW����4�S�~�̫4�=k�
Z���r�����E�EC����^�Z�okn���+i/]��;iPy�c"-!ѱZ�*�+�r�SC��:�ނ��2i`ӵCE^�Q��.���i��#�۷*�$Ȩ�3�mК�����9$+ǵ���ZF��^�Q��*�^�'�'D��q�Q}Q]ϸ��{�z�r�B/����4���4��;Z�@����q��x��]r�H��Pv��l��6n�H�������=�4��.��b�<.�v�Yl*�_�L�O����.�=oӇ�u�z�T�aK%����*w�<��{�����-�t�����Qߟ�߮Z���BKB�X�ս��d���8!��
��~���Ӂo�ɚ���z����q��'�'yu��m:Oca�f�qa�6�ܧ�x�eߊs5��sqic�]�>�~��aڹ��4��R��lK|n����;aG>�k׍Y̵^��]�"�j-'��=��3��3�Iס�����I�gս�VJά�2��ǹz8�䆔wM���1��s�k�c�0d��.��O�9�q�nm�k/_I�p��\g*�F�7��}��[fy=�03Φ����癯<ِ��b5�K��Ģ�6/�Σ�+�OO5��~VrU�wB���eܻ��lɮ�Ç�1v�ݚa]:������n����r�w�r�c��2W��|�n�;�1����H+yl�;�K3]���e�cv�4��O�@9;��*�ξ���iaz���*�X�s�8\.�w;Zbع���������E�M�_D�+Z´͛s����<1���Y6�sj)Wjs�rY���l�)��J�êZh�_�p�k%Q��rf#orvov�w1�*�:��=�$��_��o1�\Ϻ؝�n�S���Cӝ�*:n\.N��-�'\g_��	�Q~�kL���U�W͛�c0�u�:��
�s�QF%��[KS�Ox�7��|��x��E�x���x���]�:�����a��Q�o=�Q�J�c�},��_��u�/��.�ƣV �[2�vW��|2��1��v%o9�	��p6K�h�Q#W�,��H;.�����V�_��\�VOk��S���۰֖<�մ���A\8�1�����7-�5���WiK���4�$~�Q���b�lOs�� xl�T��������f=y���Af��f����V��l�ɲ����2�Q��h�.�ZMu3+)��7����%M��@��/K6meMXln�z��7��e���~�(j�����g�'$����_-sӢΞ3��L�J�۬כ�j�;��|��G�	!�p���;H���J7���Vt	��1m��}�^l�o����U�د��<�c��蟡�/mF���ą��{��sWբnj����^[t��ڤ�Ds����f�8ӍFr��F���o�W����&Y�'g�K����!�T��5���Jw��:t=���](9y�tȡ�ȗ�����eΟ=���'��1>�L\Hf�j�2e^������7�q��-�Ҭ�Sjp������uZ��2rs�q�uQfw�s���P���ע�+�[�c7�u�=,5m1�M��x�7�P�F����*�d�닸�I���^kNotq˵���D6f������v��ˤ�4�3(_T�;����9B�]�z�z)��jf$gDi&1�%����!�H���%��*"�*�yp1(��c�nJu��>��T�-���9y�o������s����x�C�D�
���R�Ѝn���Z2���O����`>���:ohڎ�t��/�ټ9����2��%rsc������}x��FPe����Ԋ�<��慫&�ׯ4����䰸��f�I�2������&f-1�J�}�YPXU�+�1���UX�g��A��%�R���x�U�m���qZ5:7��i��:ǡ�t ��V��k����8�)�̯T�йW��m�Ļ���z:8ܷ�f"�]�������/х����˗0R���X�/�rK���xw�*[K�K'v��I̥T:�֚�J�e�of�T	�-�"�kC��ޡ�w�N�a�SR8��g")���/-A��^�q1�1��Ή�њ=�����miJ�������_��"9��O���c���ح�#
�C�G�{�����S�U����3蠫8o5h����;3����"m�7�kp��*p��&��O�{�Y��5luߔ���(Ö�N��[�6���Y�Ζ`�l��M����{'M�s1��
�*���4_�1h�Š�m��J�5��/��N�A�k$�6a-�$*Qe)�����!a�����gO˪��(A:�.�2'���!,meL��*���q��)����Ⱥ�Y�נQ*�qo-<�htK�yԳi+5z��\����@��q�8>3&�lȳ�UvڝWJ�чi���J����[�<��j.��5{L]q��;�2�T����i<��q|m���7W���o탗�a�y������D��.�J
8%�8��uľ7s'��Z.�7$���F�X��o�2u�+�DW�!��X!�����Bu��yG �ߨ-�{�]�5��joL����Z�J}}�B�=3��{>A�\/�l�ofpC�E�^C�=����8�v��Z���on]�\6@��8	|oF��2&C��{��b�p�9�ѳ6��m�c{iݰ윺���{������\*�~.Mv�+x�PVL�bs^�*- ��o�zgu!B�S�[�r�˪�� �q��mf�E<��W2�s%@��n����xM�[�g[�9l�2x���=���c����Q�R5�_�e�9���D���4�^�����8:mgZ��1��܉Q�δ� yX�����*��9O�8�^��=����8v��js�2c]\��x�yv�8L5h[4;�VӮ�vV�f�y�l����+��l%��nj:]����+G5�l�gL:W:o��^�7;]�W�yp�����f�=W�'*ڌ�r3�����
�uṾ���#g������)��1���5}�N�#������V>�`I��e�r��;qg��uʍƦ���}���y��N�c��۵�� 	���ۢ�{�
�B��~���\�hL�6��2�z��}@�u['�����㳫c�yU-4bkS���O���(���ec�9[�>�{�zqz�֧V�M����Y�k�Ҹh����汧�g)`�*;j�{')��:�LF�ζ˵6�A���r+��z����]�[��
ħw�?mgy� I��vK#$����|����jcNn��Vc;���n�&�٪�ju/f�yWmy�[�r�б�tc�9����9�ʋA���Θ�v�u�Q�J����1��c4�qz�߭V]�}���j�֋w��Ӻe�hZ���]3~��4�kk/�]ݍ6 ���_�����FVǴ�q�N��%<���	Xp��hF�Y�C/�
9b&�\Jmԅ��0j��IH��x�����8���f������z_R㣳 �U�]�r�Aa_�b�f%��
U���	0
�x�'%K_[�ۅp��R�;��Kb���Y3X��OU��qu��-�r�}�Et4��\41����tq�K}����w��c+v�+�$�{T��f�\r�=�E򇁠s͛��X1�����e��o���|�{D�S����}��w����!"��T=;W�'^����!<�2/��Y.Z��\kז��Qј�\�H,/1�����ıt���i�[0��r�}�Cy��ʼ�/���C�y􇾘�h+td2z9��������*sk�Lˢ�ҝ^O�E��(0��J�;��V�]ۍ��|��v�7�c�Ԟ
���1g�`���֙3�
���GmR����p�ot�*�ڜnoy�-.��W���hD/3�Ss{��lW��Q�P��5�`��#v��;�p�j��q��w�l���,��|�eL�]o{x��b��t0��:-`ꎓ6X�s H���ݷ+�P�)�X�	y�2���������ح��(M3�c9v�*�n^��<�PF����Mu\0'EY�I�s����T�����01ו�\'���r��V�c
��V28]���d¶�e�T����	��ѝS}���bXA�ɛr�4q�h��Vk���f��x�&7�|�h��t5κ�ڼ@�S�֕b��1��G%O��:��.����|��4�S`�'8m^Q��Y��8�C�@R
��[$ ��n�����wtL�
�.�.��TZ����*��k��܇��YaeZr���i�/y�{�7re�Z.�?��|�[�,�]@���P(��!j��2	V^�=TLN!����Z�R-�fI��L�'<���H�#��f���{��y��؉ږ�𔲋�.��9ɠ��Z��VT#�gt8��T�t9�w_!��S�q�i@)���|�J����`��,Q�*65J7}3��mV^�{��g@f;�+y��y�iԳ�gl���9D5�i��Ѯ �Et`N��K0��9�ötFu�X-�˶K��T�W$R����L�Nt�ky"�뒜���KYtp�=O2lF8�S�d��>�����Z�n^�\���&���C�q��w.5���Җ��r�x��]l��m:<�5��@xh�[.���3��mR�ĲwӦi�bvm>���R��t:uu����bs��CL-��qNT��d�}���Ë"�7�f_'m+L[�N�f��uC�e�S:_8K�����]pWP��++Z8����N[�k�Y�}���΃J�dً��V*8�>��hd���i��_M5�IVA�+�&0�ݤ�g�P�mu'l�7�"ݾM�]L��@�����7p7�7�{+1��Y;C��#���t�n�rLM��%`�320�>�]�}dK��j�����h]t��*��ܔj+yJ�v�u�R#�3�P=�G�8w5�]��L���oVO\�Uϫ�-S�$�!�R��zE��2���뇃R*����6@��x:"%5'f� 쥦�VamB+�fK�V��C+�}�{� \5d��zķb�������,�6�ƞKw��f>yv�=t�
/ev�2��p�"νQ�2�ۦ-:���op��@���@�Yukr�HDL����FZ�Y�1X{7pW%H�v�jnݲ&cŪA�w�{�x{QPn$���,s�,�+,���0�엻1�N�F���tέY/�%e��4W56p�������YB� ��!��.%vNlk�H��������l`�386�+�6y�T����F�fu`�uLy�XwB+����d(�{�ے��YP(/#�x�!��WA"�=r����ԋ��t�w����}���Vb�ڕڂZZ�()XV��V�ZTQDZ�#R���lJ�-�QR*֍Dl��(�j�X����V"(ZЪ!�TDUEW��TQh�*Uڨ��B���U-��A`�m�)R�H�*�%,�"!id���j*E��������LqX��)muj(�"�J¥t�b+��,[J�*V%e�"�6��b��D���D"���m�TX���]-U*U����+�*�fB�����Qb��(e�l�U��*((���[je���J%�R
(*�eT�[b�Z���IX�J�P���+U-�#�R�(�[*8�dGV�E�5��Ub��Z��ԉmV,+lZ��YF�J4��TA-�b"*EX�U[J�Jʈ�Eƪe�,�Z�b���Z��"�J��� �¢ʖ�J2��T�Db���R�l�H�	KPTE#[.a�2�PP[j��m
�j"����(�(�9j"��G�[h*��5h喴`�ID�W�(�M�獽b1s�X.X(�$im��+�e�6�p�+C��܅V���r�[U��!�$/2��R-FXV+)��&��<���7yf ��1˘���1�i��θ�eڛR��Z.�^���R�3ٶ���<�+�X
CCϦ{���)�sqˎ�οc")�#2.��E�]1�hP㧖��y^��q/��]��w����F��릲�=��^,y��3C3h�zp��=�A����e�;����7�J�sTQӓ�4��U�ES�zɔc�����8	\o)aadE���'�d��7��Ux+��M^��Q8�$���7�.�R�8_��e�7G�nu��}�ɐq 	Ͻw�^C�8���߃fh�&�U05�e�ýjN�g/+^!i�E�;�@�_u��X�d���j.;��~Hey�l�Aw5u�F���[x�YP�*a[�p����GaOf��Ɩ��=�xu��[3��On8���.�j�H)��;
:�R5y}e�9�]ik�o�}���)c:���;1V��x��$d>�3yu�R�ؔ����͉�͔Ȭ{�<��ѯۭR���xp�,���n�i�8܌';X��읱b�i^c5��C��]��A
L�╝[,�4*1�&M��̾AuN�(!f����ܧ%��d+x�;�܇,�<C�{���^��[Q���ͤj/-E�j2���bLhԠ��v�J�a�r����،��d4����r��n������͓Rt��Ѹ�ޘz�k��Ь�zt���))LNfѵ�4��0э�Jn�VCo�lvs�Z�:S��|����|���6�$f].�N�ћ%w+	�ꧪ�ː��;*�z��o�7Z�}����h��nf��Z��q�fzkzR��]~�¼SY�t^�r|��u�Fd�XV$���B��_�x������EL������LcSX�$-��cTq#M��ͪT�m�|��+�1�i�rֈ�_k��u�����C�ru�KY�,�~����'��y
ޙ�E����a�XUJ<km�r{�<3�ۥ�4�K�����2s�pp�6Ա�Y8/��B${�E�G�#6��4`]�P���Ҧ�R��&̳����>�^?�/0���d�Y�˭=n��J��`�AW83�\�*_	�KK��Q��K�N찱���J`����>�Nv�`�ksR�^޾(;
�ν�Ѻ�c��}�]t�v\�ZS_G�{�{�\�=�'���{i'�4yC�+�^ӌP�u?P:����1	���!P�N ���`N!����y��Ię�~9��O�.�����wu�/	YXN�ĕ������$���5d8��6��RN!��=a^�5�ć�c1{@�!����<d�
C�s!P�'�Y��&�i���|��������==�,��7/7�.쓛~�O��y��u�='��`z�!��'x�hm4����C�c1�������l�������k�[.��_Ey�#���'�?2~J�g{�+Y4w��x�i����I}�N��I�����'���Y06�yOS�N$�v��<I� 
j~�-���v[��S�{�",z8B)%N��N$����,�'Y=J��y�~d���߷��&�<���I��M'yH������d+�>g�ީ$6�����Wz�n<���u���b4D{{�"4A��A|7I6�k��i�m����8��|sܞ��'��OO��|��O'y�|�~`l;��'�$�O9�H���7���]ٯ&��:ce_Ө��#ЄC��!�C������Ad���:��/���a��q4�6�?s'Y;��w�8��Oϩ9;��䟟������.���"��͜��>3.j~�X��">��O�x�����VAI5��Y8����q��S���|ì>N&$�a�ӌ�݄�)�'z�d��fW�:���u��I�_*���y_{�=`�=��ޡ=`x}��LB~C}��(|�|͇5�d�C�lՆ�RL5�!ĝe`y��q��S��2u���Ǉ��=�m>�8M��gëV���X����s�z�d���`~C����H~g�������Cğ3}�i�qɳVM2O�É>e`zn��=������®�ϰ-˱;��b�����ݸ��u]��*y�:�����ޗ��d��^��� �w`�t3��wݛP��������j�_w;n�y���%K�'�����oml�Z�{S�үsb�Ir��p:�u����Q+�����z�raɷ#��B�� b�8�a:��ө>x�{ڰ?0��'��RC�;��A:�y��GP�N ���0��'ɳ.$�a�<ՈB,{�A�N���Yƾ���F�x����hm���v���>@��S��	�O&��R~~Bi6N� |�l�?w�=C�x{��J���i�+'X~"UU�W�}½��4!�����nMc��~���m��w�?&�O��Xq���
d�'������h����N2y5�?0�u	������$�w��O����Ԙ���v��7����~�������'Rw�`�q��o	�OY���d�M��=��,�Rx�a�,06��Ρ:��)���&�9H�#�l��l�����ݽ�9�*�� 	'�~��I�RN���J��VK�N���o���'=M�ְ�a�(|���=��Xz��@�C�??�4�b">��sL���U���Ws�ܯ�B(D1'�,����|���y���aˬ�����%d���a:��'��f�'=Mn���'y7C�+��ѻ�C�"�P�_�gqVFf����Y�D`!�=���O�X;��q��w��I�Og{�2N�y�IR�����,�n��gp�d�'����	���y1h�y�C��%�>v��	8�p}�ǩ�!߯̇�b��Ad�0��8�����,:��T;�B��'{�a4�߷�Wl����"��v��@]Uu�����e�wP	��O�E~���8��t9M��'y���<By����*��Ad�0��>d�T'yg�:��T;�B��''o_�M x}�u��������}~�?}�L��>�R|�ә�����7�C����4��'���~C�N �=����4~��RM�A��8�ĨN{f�u��iﾟDp��{��Nk��\����%[�z�Nu�+�X��хL�J[pLԱHQ���i�����	��=׶��[�S���S�yҤ26�q	`yF愍�Mctu� ��v��m�Ӡ(t��l��z�)`I�����_R�w�L�꾘����Sd>Vd������tv��WV�������f)T�,��� �olN8�i;�"�o�㹓l��~Lf$8��{�=g��Ad�ݓ�:���hO�q}gSL�l�a�N�Bg�n��C0~��J��=�=�ɏ}f@���'��z��߷�|�	��9�H���0<9�6�z��boT6��3_�:��O7d��u�<���'~����];�+��ߢ�X�y�G�UG̜}a;�q�����w�'=I����M�:��f!?!�ԋ�L[<I?!S�<Ad�5���J���o������}��W�{^��ěeN�P�$�O���I�_�q'_XM���I��'{d���י	�C��4f!=Cg{�)�<d�7;�4�8��ϵ���x��se�n�;����G�c�9���1���~I�N{C~�2q�����I�}�8���	���=2~��m���z��C�g�38�ù��zs;c�����������C���r��z���&2O��Y>J��t8��'}��!�N0����$�'��aԟ��M��@���M���YP���|����w�����3�G�S�zD@�5W�DH���-��I�?RN$�4X|�a8�2�Y>v�xZd����l���Xk���$�'����8Ρ4�����{�_u���׻|��m��=F�{��xRN!�}�D�(O9g�VO�Y?wXq'�Q$�M���5$�5<�������`|���!��y��z���P��/P�f�}�ǣ�DE9�"��M9�!�q;�ށd�!�;�I�P�r�aY>J�r�ğ�7�1��&ӆ�:ԓ��������5�6&=�:���;?Pބ�>���@�D�yz�i����a�8Ͳu��!�?2y��@��I�s�I�RMw��
��VO�I�O�=򛚰�d���o������7���}��|��N��c�:c�]�����u:��\z�T픷����M=�/n�ES:��٩롽�<,�w�r�t�ٗ#�cx��'
z�"�츁{Y�E��"�s��L�Wd�Iq}P�52�{��]�ɰü#R�����k�J�����u�~G�u߻�{���+�$��rÉ+�C[��Xbq�������~��ĜAHxs�
�Y? ���a�O�w�ON��3z���|/�E��h�����מ}��>�������'̟yN��>@��ݞ>����݇�z�2OoR�bc�8�W��i'R>�!P�'�<��H�h�\}�_��{���:A'�5w�럿~�O�޳�/d��&ޗ�"���<���M���P�`m5�=a8��v��<d<7x�u?!�<���IS!�xu��R}�Xu��V��������P���{�m]_G�Dz�����M2xw��J��u�y�)6�`=��>I��j��!��=M0�$���i��?Op��:�G�u�������&'蹷')��ءn��({�"G�/�=a���V��'������I�O~�D��I��,�M��������7�C���G���$�
�vOP�'�6�����N�e ����7�=��C����hx}�d�+!�=Ì�d��I���̟�<;���'���tO�I4�sܑC�q��s&�����5Htz<���U���zyh�C4�7��ë������z�̜J�hO�qO��i$�{�:���	����I��'�w�u��'��	6���ޡ�'�s��!X�C�f���Y���|yƚ\1^vz�q6�3�$��2|���|Ì�J�'�'�:���s��q�֜d���ϐ:���N�d�Ԟ�!���1�FS�"TOt��'v
SS��1��;��"�Y�'ɸwXi$���x��|��:����O�q��Y�!�N!�;��8���ağ��L�菄{G��V����ˏ���s�߷��3�z���y��!ˬ�q����C��'r��q���5Cl�I��Xq����N�q��l�8����$�F�^v���t�o�5�g��n���b��#՜ֆZ���tyӫn���D��)B򻄕��f�1UJ�5�tZ��'���}Lp⃗%p�-W.�]��-*�^���Σ���Qps�B8?klJu�&���Bë��Go$g�撓����?�W�}���~�.��7����|�$�~�>C����l��|���C�s'P�8���`q2z��,�䞦���4�|��|��P��:��>������7��|>|������=CЇ#�b=�ƽ����	㳽�!�m�a����8���$�(OI������N��d����8�����8�q~~����9�w�+���w;~�Cl�~Hv��m����������k�?!��	�d�2P��d�w���C���Ԙ���9��Ld�+'�Z�8��OS���f��~ϵ���]k�)�M�~N��~�I��!ĕ���:��M���a�ƝBu�����8ͤ�=����<���RO�xw��++	����{�vo����{�_��_fsi+'�\����&����2z�7a�CG�:���=N0=C�?~�u!��b���B���Ag�9�8��G�������sy����~>̼8�=I��z%ea59��J������$����q����RN!�n���Sw�P�bhd:��?}��8���o�}u�Y���u�s^������/aP�'�Y�,�a�N����$�M��ԗvIݿd�'��<3�N�q'���VC�S^P��	ěa�M!=��C�c1�������p�����=���g�)%N�w�>AHs�m'=J���a
��Mw��x�i���Iwd�_��>�>��,�m�6j�1��3#��#ݜC���8�M'������~g�>A~I6��=O�RJ���N$�+!��d�N�~Jü�z��'�߷��&�<���I��M'�y�Rz�`y;�
����<�9sν��u׻��{�������3�<Hm�9M��O�y7@�$��t�h|�\�SL�l���8�����=��N�~$�w ������h�GG�n<���E㖖�Gs���oQ7��ZM����Gĳ��6�;�%�5���[u�-!��8��c��j�z�@]�����Q�����W:�ݑ²9����wV�dHB��1l�kBB8�@3���d���]i��M��h+Ң�Vk�ޥ��V��l�A��$u̞ue������=��9�����a���f�C��٪C������2u�ɺ�u��_l'�8�A�8�d�g�Y�N�a>;�2u���O{��䟝_;��{�g�_���2������8����C��!��ɴ���M��h)&k�Y8����q��S��a��q4�q��c��g������o����?f�r��?G̜I��'y����??�^d&��sz�����"���O���L��~M�Xm$��$�+��|���J�2}�c��z2��1�̬�K���Jέ���I��a�O���=�(I���}�I��:�����C�Y&!6����C�x��l;��$��x��>;K������Q�lW�`����o{��9
�<|gO��P:������v�I�����������M��Hz���|��d?Ng�:�2q���!�8=�#=SB=�=<�>YC��g��9E[�w���2O�̟n�yhu���v��i qS��	�L�:���I��r�q6����Ch|��̒��8G�T|"${�D����W�~��.s%��q��t0�OXz��8�I:���N�d=-2|�o�����z�a8��k�~a��I����|ͤ�{�d�A�^iw������/3/$�'w��T�2��sXq��Q��&�����8��X~d��!�[8�ԛ0�X`m��Bu�Lp�1Dz�j�e�B���c��=�o�?!�K�I�>��&%I5<�8�����哉>d���Մ�����XN0���+�!��8����Xo&">���S����p9ߖ��ŝ��&�;�ru1? �gy�:�̞�5��<g������:��}큳<�u��Oώ�XN z��XN04�W믅����o�^���T�_��N�Y��[�s�t2�]��:pĎ�8�u�B�.�	�:`���ƽ�D)�9�N�mb���{k�k���V������2��jRڷ��GzF�U��s%cP���SOO�7�or������j��v�T���X&Z:g��_���DGZԏ�s>���d4�&0�O�$8�/0�,s!P�'�,��p�I�&��z<d�a��ޤ�RN���,�n��gp�d�'���'Ns��ow�_>����׆�~}�}�W��!���C�����1�����$���a�N��<���Rzʇ�y�*OY5;����'�纒��N��"��v�����|������-U?D��B<G}s�GDm5<����<7C���O7�$�
���Y%L<��8�	��d�N��ʆ��T��w���$�s{�s7��1Z�<5����N�~�PC����^�=x��Xx���Ci�z�!>I���<d��i'�u~��RM�_�Ì�J���=I�Oߩ?~w��U��3�cO�����ޱ�},��ziÿ��?8�i<;̑I����s&�P���Hq!����N �y�'�u��/��'�8����i�m�\�nG9���n���u}��g>������8��'ߩ=���O�?;��$����a>q��~9�H���0<�d�!����P�$�_�:��M�zÉ:="6k��n����ҡfG|�q�<�zǎ��M0�a�9�u���&��2u���OC��:��'�p��'�;��:�B~C��&��x�~B��6����W�]�o�d-F�>T>���`�;���:�����O�u����'y~�ĝ}a7�L�Ԟ�2l�rN�?0��oP�Hxs<�q����ȧP��p�'�1����oR���t�{�Dz�������q��X��d��ކ=�=#�O�_#����g\6^f���������YكD�|Ð�WN�.s�J�%I�7��\��زk�*��>�Ih4����{0��CYl[��p�t"N�Ԭ׼e��i��`�ԮGg���L�g"vZW�l��]7d���U��ݺ�Չ���VԬ���m���P���%r�^N�70;��"v�a5��3��U�ג>Q��%g�ծ����着=�>�p����8��h(��KLL,��W��]������
�j�S�q�E⼚*�R�O��U��EZ��X!��W��@|t@���cܷ�Ui�~�ˮ��Gԛ&%��L�W�1��vQ��XR��1�L��ˬ8,>Q9\�)G8Z���o4\dS{r��͑���{���X9�p=^�s;x��� ����zb��6�+b��&�&j�r�K�I��˔���f�>�_���vM��^җ�0��l�����I��!^Wh��]s�r�ʪ�� �q׾t8�n��9�q��ƨ[��D�4ef�;ס-�&O�1�oi����q�Hׯ/�4�}�':��m�����WQ���y�Aov���ZvkZ�ۇ#7M#yJ+���4-7�dw#��\ ��u���㛸�\7�Ρ�g,�:�{�3�U�:σCKG$31��*yvk1��p���3�H��f�F�z���*� �W4<�������^*;Sv�s�)�T�.-̧VN*��;e�l�b���ݡ(���r��F�ն���݂���R��u��-�w���/��o{"��-����3�.\u�{o�Q��к����vl����I�0[���>�S�p��*�q���4�^���b��0�/�5�ծ��Ŷ�Ԑ�,���z��z#�5t{Z�i&�\��� �ق���@q�O���۩�\��LRKWSð9�A�̭ch�Զ]Ц�=*֊���°w�������1��+��j�e)oknP*���U-4xp0��k.�(�������S,v�F����wD�o6�0:ģ�4����k4�d��@�;2�Nt�T��uʖ<mmGV�<7h�.����t3_B��{�����y�.�qU&ͭМȩ �b��d��ou��2�q�/�N�adw��!���,n���ek7�6䁻�i�n������1��Jݸ�^]i��s�T�NZ�]ݏ(*cn�`���M�����_}�45��3e\�j��quʞ��X��_�:%�7�4��fxd~�${<3�˦�n���t�6���qZD�F��P���Dn��5�G\x)�-&��Ź�BJc��}]���K��0���,<�V�\������`O;zsh�Z���M�w%rI^�f������s3����7p�Pqj���j�
����U��:d�`�(Zi].�:��wR�'�+k*&��İ��qu-]��VQCtc���l��S�$�c�*��ϯ1���VlJ�gd��Rc%�T%���I�u�ai�c��:��1��p�+9�0Ym����d���_4��U�,�x��.��.��㔻b��`|��U��.��k�&
����%�� �F�D�܎X"R��
U����jCs��=���/�����4G�]���5�%p�L〽�m��h�
9���f��k�߫��]0����*��Q!�-nJU��stS�f��F��I����;�Z[���$3��χ0��^-�az�6�����8�ʽ��J#�C�v뻜�*V��'���J2E:�Z�&�\�PF=7�/P�㓚t*kÇ3�3�2�[g��v��m����.�S�l��$��7�\���T�ݗ�*�3>�pID���/�k��8�l�hȖ��;�g�]N��]�W�6c��a�P}��2��X�#d�9��
;e���;r��?�	��������37�$�n�'�+�&ڗ�1қ;�ٹ�*\��*D�7��a�Nۮq��d�Y��y�M��pc�:����o
x��gd�V��C*�),�˨N4�b(�Y����t�79���ZY2�Ŝ�=j�9j��̄�|0�.�&��,�&�C����(QE�kQ`�m�Ee��E*T�Q[K�����"��E��*�+*,X�P��Ir��P?32��h
�1s$��ZJ**�TA�1�B�:l��Q��:lPb)��QMYQQq���E�¢���l���������R:h���[j�6�"�c���31\���!mX5��Z"2����U��*��iX����1Z�cQM5����FQ��1��DE[J�"�V�1Ki����ƪ�E��,Tb�i��"����%Aj[cD�5)�1aZ����Q�*��1b�ҌTDUQ�,DR,�X��Z�0X�FERZX�T�b��0�����1dU��Э(��X�FҪ�X�������RZQQ�آ��J��*,*TjjőV� Mo`�b�4��s��_���w_��"&�	�1����N[�saȫ����w)u�<c�[�n����'NyFĝ��"�{��Dz��u����U�i��1��zr�t��V}2_���\��4H��F��<e�������jme�UK���H���R%ﶙ=�G�4��dkV�V�!�ׁ�us&wl;7�W�<Q���x=��_ѧSs��*���0�)�ʣBԴ�"E�r�5�֫Y��ɍ[��:c�U��-Q��䠮���
�n��]t��rgm�]L�:�vL�/;6������^s]�,�k�lˇ�D�<S,�jY�`���Q�Ym�ӫTU=I��~{k5A:���C�{���+���r�2�6&K���0�^��]�/�	�v��OD7�������2������c-�q��E�/��X��h356�Ks�'��x낄����ی,6�fׅ&sD�5����P�
]:�^vs��);ҳ��Q&�W p���o��:LP��#�5��wײ^o+am�L����%RwE:����P�U:�b>���7����H������F�S����mkUei���1�{q
��Mv3���+,��;�\��_ˆ�+(]m�"�3��mtmY�=��q��Q�]��������H�6m�
&a6?�:y?W�7-fo�ɶ�*�F�n�A���P�C�Y|d��W��x��U�k[Dwv��m��.��� ���$���K��LV����6(0��|:�et�ާZ=oh�}g�8�>�=w7��B�,�N���̾QQ5܊�`,�6KFF�}��uグz�!gj:�k0eq�V>�_a�[�^`�%M�@sV�_l^�D�]ؼ 
��w�����1��eRa�]{ʎ6�5�k�P�S���;d3Z-H1��9�b7-!0V�=ө�RB<�5v K������
8�b��F�v�Y�!@>ͦ�m �!;��:X���������;gG��������i�=c���Ç�o��(��?gU�]L��e�R�&���4v��]��8g>켪�!�V�{|����s#A�x��a�9���:���t�P�|K��Cé�-g+cq�w�o�XP��ӵ���q^�>l��]�aͻ����b�Q�}uDu��R���uN{����)�rS����*X�&5�p�\V-�`¢�K��̡yG$�u\�R�Gy�ǭ*��tb�b�T�n�ӏ���S��Ϣ��ڪ�7n]���팝��'�8M�=�\�	��7:��Bw����㕤j���3�� ��Eh�Lb���8Պ�4N�	��2�fXɧ��l�wx����ʷyv�7�fi������p�f�-I������W�3ݱ�D�[�`��zqz���f� ����=��oSp3ՙ��ʺ��c7�Q�]%¬3Y�J:9��Sg�����&��Ui��m���~8*�z�� E�5�k��v
�4�������/bXaDA{,����M����{�x<�%�)=�x�5��c�X�i���⡎���E�r��7Gs
	���i)��w`0�������#�G[Z��H���]�Ә/+�{A�U���l���ҋD��3�P���Pr$Y���o{�su�\O7�p����B���/���APα�ҌX����ę�Y�/�+'N�	ۃ�ek�e�;C F_X�5-S����ȴU��UU�
~���F�)G�x�L�W���`�R�St�:X��zw���ꑂ�Ʊ��L(�����}��!.�S��Y�����=�N�q�<a��zLY�n��@f�V�p|�xܡb��S�	Ѣ�}�N�D�.�r�N"���ԩ���؍��Ӻ�M�1��2��D�u(`�W�R�X/TE::=��B[|.�9 1�jQ�������$������3�]��I-0��%.DE@�v�N����
ޗ���&Fm��Y(��3���^nO�� j��6��9���m�# �Ig�k��b�B�\3�t�d�Lq���*�U�Kt��DG�\�V������+�	.���j\Ղ&X�f��*�!Cx����]e�6�jy9a�z�4���Y�?7HpgCexb��1Φ-�*k"�N��������觺M�����ܤ��E%�+��@w�ס!�U0��u_��]^��Tެ�(kc&�^
|'�0w�&��=bF�&���藡�Tmy�.��%��PV^(#�z S�.��Mꉁu6t]�Y��ׇ*�M:x�5�H"Cz��� �G��3�S�bg���c�R�x���K�'1�J��ٵ�E��N�I���,+�@a�b�d�
�z����0��b{n��u�o�dU���!Oi�^�n�XpT�p]x� '<�m�+�f�ͼ5�|.{eʭ���:��Ʈ/z�
�3�n�t�r�����]%`�H�^��=[�m��^�!HVl��e�~�������xr�y���(��ؒ��.�J���V��g1۪ᥩ/����F���e��f�j)ꀭT�� ��O��V�_A�7�����\� <+}�V!��@�ܿ"��a�YG�L�S�䦰k���v����@}���g��w+�_R.-���!"^�4L�@�M�ZGx7I�u�$@U�}���q�eU��c+(��TOp���{ޏG�vַi�Y�{"�K,����&�L;
�o���T�e����Z�U��4��w������2�H��Ӧ,kF�p���t�ʶ#.��5({/��O��H��n��8׵�j %�������8�h���r���փ��cyx�7�w��e<�C�<���jy�<���8�ZDP�W�˱�i_�#��;S9��:.�ʸ��c`o�s���Q����\9�X��j�DpZa&�qw�:���,K��OE�z��蕸Z��x��X>(�)�k�f\�Jj����n@8����"�m���Nm�uځ6w	��x[��O�;V伡����bB����s�⮮��x��b��.a��ͩ�����0$qE�.��rib8��YΘ�eRvk���\7(q0V��4۶�v�6�vz��пo˳6�^J?2�э���%k�s]�,�k��p�h��L���r��C��,ԬJ�t �k�+5}/�8�d��`���rW��
ֽ�-bd�h�#յ��;ivV*�OWF{��S!Wί���|������3��b�Y�7�{�1bt�p�*v^(VKںӘ�}�$u����:ح{x��y�����7е��K0���k�_7��[6�J�>7���V��C)�"��)FO˗r�+�{���7˵�f��n��������(vmHA��,�u�*�E��2[ȸO���8ؒ�����qD������0[4G	��=��3lyלU�רc��f����Y���S�C�����Xff,�-L�U�CMT9�ejL�@�1�R��slՖB��츕�ݗ!��縇K#�W����2%..1kg"���7l!xv�>ͩ�<�b�:�\�����ŮQ��]��&)l�\��tE��P3�u�t��&��|6޿fW��ޟek��y�����u�J������C��6'g�g�,#����ͨ��|i���6޹�<�P/�8�>��4�dl���(*��%��"��M�'gzμ��{pe��g��V������ sS�F�-�u{j�߲��G�eaq"4���(����{;� �����Bc&��1"�Uwk��u��x��������nB���v0�;���L�u��;ި���������eƈ�٬�hq��/�&*�t���p{�݋Ei;�cӭgg�-L��ۑ7M��SsC���nq�kv�@ьa�=DL�fܣ��i���e7��<�p�Y��_x�D�'�,Ѹ���y#��:���@B�"�IX8�}�j�KS�i�D��lҭ��i\��]N���.�nx�e��G���k�N�զ�P�;�V�{^[��dh)�7]�tk�4�
��t��|M�S������al�z�b��\0��u�ԧ��\W�Ke�s�g-��Cy�҅T�� i���h�H�a�3+<��?R[�<^�ڿM�Y��{q�=��X{�7��6<�!.�R��]�s�̑�&�$�m��bZU�hC޵���5�ߜ~��k§4�Y�Y�&���b��C�-Rh���>�.�B���;S�Uq%���*��5t[�0]�jf>U��g�v�n�m�{S��m��p>&��^���R��j������0^��T��E��#�;2��^ofа�6�1��b)�"�T𙩚r���s��m\GM������eq��9�6H��e�b�yM��0����!Q��p��WLv�ȹCg��˘�n�Jߗ�`}����:i�㡵U{+�z��Q`�%��K��>O-%<Q#�3���N����8�"z�%���jX�e?	����(gϝz�B<l�Bp�[l]����`��LV]��vY�ı�њ�C�.�Lu������j(v�5�e�����E���~!Z�d>��#���wv�(g�Y/A�j���R��C���0(��L�)�Vu �Uq��ϙ��֞(l��1�����.�2�K���{�R�g>����G�;+�=˧53='��y.���z*5��7l���M�`�뻥�;�bBk�=�����(�O��n�R�vO���ρ`��a�t���3�ߵؕ����wVřks�7{�ޥ���7T�N����`���1e���3k}V����@�9P�z,I�yb��5��ϙ�*Z�M.b�#qѻ8���)1e�T]V����9�����o%�?_�T����Rb��yU!�N��9A�܇��iVN�3C�XRB���S���]MźLk�$�F�w��8$$�r�مp9�՟��֡�w�����Z�%^��g?`P�-��GbeW�~� �F�c��ae����ޡ�Tޭ���T��J��s��̖j2(�XAª�L���w��^f��	uY�e�(#�z ޯaf��|ܑ�s#��m@`=:�"s�fbC`�O� �c�����d�(q���W���-Q�$y�r�)�-z���`(�,���q^�
��4BC��Y]���õ�ۨ�p!� �^��9c3����犃Cۭ��Q���X�}k��H­5�8l�e��Se&a�4X�{��R`�������/v�t�RW��st�n�-��{����vedš
�n���Z9C�9F�bA������z+����\�Vf�~��C�߻hCb���t�E��`�}�^H�r�%���HK`�G�7�K�ݞ�n�!���ߩ��0���R�w��7�:��p�O���`�:7S8�2�]h�8�m�~*��'����;^:�䭩^��7p#`ISU:���m{�,m�^�NK2�?�夙�PS��P��m�V0f�j)���� r�mU�ee��o�r�jt���H��u��^���~aA��7��v�G+��٪��0�@��O^��W���D�8̘j�C�ۋ֍0�*���^n|*�~�y�����SAₛ��}�v2��cVX>5��%��n9�Z4?r����h;�cy_�H��RȱV�ݬ�՗ν��ZC2����c4��;��hy���{��N��det �}n�V6V��}������LˍU(v�\G�֘I�\_5C���P�qv��d�=�ի
˒�GSM��T��^,�>h���ڮX��b��O����-�F:i=�bn6�R���΃��]hp
iq�ϔg�+|���.+��O��>W|�uwZ�}��ՠ<�F:�,�1vf�Փ+_G5�mM�,�)oH+ �+/�ojE�:#�6�!+Q �Ն�ө��R�g�C�4u^>+���d#�K��G��K;yR�N�L������s��z3�����ө�M��/�/��ΪC�K���y���n���aA�h����g:c�EY�b���*uR�!�[&��q�W�"+L2���GCs:^�{�ud��㭆,������\�gK'Z�̸A�4x�x��M�Z��c��e�Կ�V��&��<�F�b���a��f�'"5�j�����P�kd����5Oe��p�4=R��-�&6eXI�ͬ��2�{އ�\��Vj!ָ	0Xyv|���B��i��y���5�$Z��cBTPf�^��5��bf��`ͺu��U�ר}��	�p��Z(b�Y�2�4����m?86�x��,PßdX��x��(ي�w�^a�1wq�1W�:�uD2]�C~���(�_��,�^��EC�U��b�Xe�����E;��A��Ұ_���#��;`J���� �{բ�B���8µ_I*�z�jS��!�J�GzfkTMg2�k:�#�:lN�zϢ�0���� Z����׾�b����y�Z�b���GU�X�t���s�w/��3-��0���eX�:���u�x���;��Kдe�je�T�u6�OC�	ņE�����&�����<ݵ����+)\�t��%Q����@���#�3zu��l2���nΈ�u�(��w�+�X%�ųS�������3a�u��K��g+Ǵ7��J%�8�se��tqjޚFB�Mjf���]3g*�71"��ӠG��;x��,SJ5;,�z�iJV��ÅX;t�8"2���6�CX�9Wc���5��^ݙG/q�򸑁�,��SfG�������
{D�@1�W�_R2�@n�<�&����Z�,E�J��ݥE1�S�gR�����C�v���'b�.�Q:T�Am4�i�V�#ĺ���|u�Z��;�G]��dm#�Y�Kc�<��P6
Ŧ$c�o�cz��.���v�o�V���r�(ʊ�2��[�ȵ���_8ܥ]iΖD�E��=n��Wƕ�בP˰����8Q��k�xN��л�[��J�������J�+J'Z��[�zy��5SOw)C��V���rSbPw�lpz�bn��7Ы�[}g+4,��s]��s�]P2�f+ڽL^�F�)�T-��,�XG���ז��M-0�A�s��P�S�Ot�NͲ��[�қj��W�D.�I%B����V|��-����e�l����Q�F�dѻ���ň8�"ݺv�ܤ�;R�ej��qmÒ�z3j�	Wi�	�lN���IgY��s&�]2sjeoZ�t7I�؃-�eGqݼߺk洶�$�]�i������ݥr�ʊ��UH�F��/nk���X4�1K�o�z�����Vm�p��^��g&���9A�&ɽ�Kt�����j�R��T��r���*9�V�*慓���ɕ��m���N��&�ePf��&a��߆:���ꌙ�j��;�3��T"-W��g��G@0��)o4�(& �˔s�rm㛙�3��;�b�BX�彖U���7�=����K�u۹����(��h���;t,Y�t�E6�]!��07M9�J�\܀[���b:�55wi��W@��y��z������;���\M2Z�Ǎk܍@վ�N!mn�ݩ+��tF*SD�ܜ�<��j�iGyڈP�t(�y���P��]�w���D��]Mt���uhXO`�6��ά%��HI:67��F�:1@9�fu�^]�Qst�Hi8^���2^=f����xg-��-����79�������:ě'9�)��u�����rKK{�˸X���5.X9A��H+mmt�Y���r��/�5���u-R�r�1X�x+�����u'}���$��o���.�2)`w+v���멻Y���._9�9��t%��oM���$I7��������{ X��RUe`�#(��J��"����[E�#jE
��AJ�[T���%���mb�(+PQ���TQE�Ժ�X�R5��j+b*�qYU
�*��
DF5�`2Т"��h�lQTDQ-l��V�eB�����R�A1�dTb�"��m+UF(,UEjQb�
	hR��X�e�Ģ"�"6ж���QZ�.�2�b�ڶU�E-
",PRڰU-��aMR�1�J�lDr�R��D��E#�ڢ�J���H���EZ�b�F$�AUX�UQm�"�Ҭ`������QX�F(�ت����EU���Qe�Z�YQb��lVcX� �˖�ER*V�
�j
#�MaTE��F*�����+PE1�� ɗ˥D�p'MLpo&B����)�bQ���c�ܵ|7Q���C�Ɯp��K�a.�&w���i~z"""=\�����UJB=T4�����T�"�

��K[����vq�z� =����R�NV6�9t�T/U���Y�r���z�K��hp�ło�.����(�����|�U��7q^}��jn�ڀ��>�����a"#ѻC/Ǭ� �f�r��i��dJ�U�� ��]�O�$�)�O�F��yg��ƎzkA[C�Y~�>�0"�҃���Cz%)!�v�A��経�m�K�Ա��GsWh�p�d�`��ȼ;�9������ң���#�� �v�x�GG��T�,�asi�N�0��?y�ƹ�g-��47"9�HE������޻��캢"Q��tO�JSp^���N�� ��ż,b�wX{��+�{�o��Q#���q\$8��ۧ�J��:1w�}W��q����c���D��3�C�M4�a���[��f�:S*�lvTSf��5\ �������uʹ�F������<]b�<>�|��!�a([f�)J5�(T;�҆�f.
W���7r���� ��;�����9٣>�Էxzz�6c0�EM���|��[.����wH,p�WXD�Z�O�����|8j@��Sxc��%Vq홻�۬�rX�}Ʊ7F�s�"��\��Ӄ	�飅�+�m:w3�h̢�W"4�ܔJ�=�G�/�b�Sj�Nإ�
C����n8.�R��@��SS���z�!�x�%<t7�o�,������q�Xb\|w��loE~0g�(a����FnE���&���5���	��,�Y+5Ⱦs�5�(�>�s�q�uUW���GU0q�Qh��Z:l�}�yi(M]g���*��u��^*d�0�O�Cl�0ϲ�]A�]UW�uT8�9 z ����w�RN�}�gdv`硅�9,�@nI�b�p�T o)�6#7n�C��l`W� (�������B^:(Q2k��Χf��8şCzgK(^�� �`���٬g��k�+>�Zf�;�����d����"pϜo�Ʋ���s�x���p�^�ۘj��M!�5J���0Y�|v�9��T*�S2ĩk�]1�#]��&V�ރk}�;�����F5�¸'�}��\�#���E�_tT9ݳ�sg!�v�l{;���|�3C�dݚ��m�ͦ������*PqՖğ,�(_T$��\[+غ+��;��l������"�6�wL��C�w3Y֣ޘHԤ�*�B�ǉZU��Sî�d�'�������S�eI���]��4>�u�\�PE�FVd���5N���Vl��'4���Q��}��Lk�M^JJ��\�,Boy�. ƏQw7�;�N'szX�8w��U_}��J���sS>�U�T�ġ�ձ���\jdb�FHA(/L#2�Fb��y���<9�<b~(�[�c��f�\�=C��H{Pm�י��yB]g���S,{h�#����S����f��`<������٘��P���mj<��:Y:�=�_n=��l�}Ű�m��
�z�i���t딕�`�@_�9��&٥S	���g]������Ǥ뚼�C��*���B����r,8*`�a���nZ��g
UF
����%uR�R�G��ñ��j�oVT��*��΃��Rw��54I���[�m���B��e�(H�����2|/9�k�U?�"��|���kހ��(���oZn��HV��Ή�ӵw�����d����)C�]�pU�����dZ��u~�X��'K5���Er&|�$ȑ�I��2˜�y࢖Iv)ڦ؂j9&�m�@�d�W{���]�D++�\�v$@0�ٓ\��CӦ,�i���1.�Y�LA1�o�9ǧ.b��HQ�`-ύƴ�q��A8U��˽�W��cCB�Wjܓ
�]��[F���l�l,]��WF��"�]��v4L��wmud���r�aa�rB���æ�#9�2�*V�҈����̏���v�Rc2�*��T�?}�}��*���՝��sr��Tc��x���Ï�`��:鹶��F7�(@�7Kr��W��Soֻ�i"�>9���w�C�l�ϖ4�x���M�k�����cn�1^��<0U%Pl�1z��p�������u�os��zr�t��Q eٱ�Z���yEqa�g��Qw/n]+t�ѓ2@���C�]��y��"���q"W])�]�v5�켮�ʆ����G1*���<��s�]\-�08iT�Pa��6m�@�j�v���7�-¨���t��u�3i�ҡ�ЇC�5��dtH����v�h�k���B�̴���ReC7>�fv�.!���+���d�^2�$��T�.e�v�F�Z�R�z�{Za�K����1fʇ���C=|"ۮ����Rc^\�l�JȯJ}ˠ>ȯ2�3䎗��U��Lkʹ�I�A�s���u�*�z�GS�اb/	��zr��u1Q�����Ȅ�'��|�xc�@E�ZN��٨�}��44H㋍��^ʻ̹yjl�.w�w]ձlj��͠qbŕ睩o�׮�1��e�a
�h��[c�9G��]���}]��֐�#��^��b��W7E�E�s�e��y]Y��*uˮ-
�YY5
�6���V�����`���~�DG��{����NTQT`}n���qq��31~��Z�1V�s=i�`u�V��{��Fq��	����<�ua��c�'�.*�]D�@�Pa��r�5<s�lh�ö�������wAsS`����H�;i��zz���P��SQ�v�ؕ�f��:GاL-���v�(p����yM Z=�p�]n:�%� ���Xk:�#�:g�:��Z�t�ۋ+%�y��:V���U�f��4�h��o]ĵ�ȹ �a��:����]��὘|�M�wkZ]וViq�w)�1޻�hp�6'����ס�۬R>W͎D"d�̞S�.=Z���T�>��Z"ܑ�h���=d(ٴ܃��9c�����f�í�Y;`�����}&x�m��U.����sˇbߘ5�`Ek�����K+kQ1ȣ.�r��!P�n�w�N�N��j��o�[������d^�I����굪-<Vڊ��j}�q��g_�w���S����+٦",k�g-��46*��]�^z]�u>�ft�+�U�L��kn�f�b�r�02�@H�9=��π�E�!X9V�2g�)��6��v���ܬ��_v��S��"=��؊���:P��|t�mo(�o>�Z�����I����зY�k��V�]l��8��ߣ��z=�v��>:dg�T��}uD;��W���M�M�x��P���?V+���n��ޓK��v��!Eh�����I>�6%�U�i��ز�T|�n����D�hªVŷ.��[ۚ�u�ʄ�?'��L��n�ʀ|���QLm�W,�W"�Wԙ��͢�௜�{��gvm!F�{�p[�yY�6�P���R�kxP�tʙcOV��G4�C*�9�Ei��՝~��5��Jl���j�2���[;��s�eV�sZ��
A���3^i�0>���:|��E&w��0E=u=�aj�#�E�Vmp��!k��7�;�����9��-�,�C���K*���߇]��T��0���a��'g]Q��eڞ�2tu\4�%�e<Ck��E�;~��<[��E�T��Ak�惓2ōF-Z3lm�6����k;mMK���ɜ�GP�aX�1����7�h/���,��}0��vu�K���H�u�TR�s��.L���`�D��T�nc.x\�B��E`�Jo),YP⭂RU�=�+9��Y��&:��-��z�]<���ź�5s�PNy��0�w3��%͓�P�H��*�9Yf�xBz�Aʍ!��Cr�Wj'��oޠ�K�1J��ufV���,�ż�[��w0.�	�8(�諭���.�]M9҂�y;�h�/v�vr��F,t>ޓa��`I�ͣV��ӕ][�ۉuK���/_<| �j�+���k�E��;�k�Ø�I�����מ��z��0(�G�z*b�%�R��T���x��/�Ѹ/W��r��k6ǳ���o�"��R�u��D����^�H1�Г�E�0�\[+E��;<�j��T:מE�Y����L/{q<�4o.�0Wr�d,wV�Q��jdb�Fw%q�x��}��3��cݞ6��IT>q]�X9���l:��`�uSk��3��ܠiҙ�(Awę��U��>L�Y��S�փ��p9m(�t���ɡO�
�ܔ�qR���3�Crj���w^��t%d��������ʹZ�X�u�J� B�Y�]r bY&���|n�n7�+�s�z*4�Y:�3��*������+�w"Â�����������%�t�\2ubQ��	�o�b7B�e��e�:��=����Y�]�|����%�o�y�B7�7݆�ԡ����t��.��T4��5�� ��dyg�7n���-��3銮P����(���ደ�u�$���B	7,<ܥ:=ڵҰZ
��ڼ�ސS�GI��)�2t���j�dVhb�s#�|2ܴ�Hc0(��{��z.�vs���U1�>�񹙰���I����9���N�"��u��x\	��^Y{�=�~^�`E��о���/�w_�Z$�	G��GÆ������2X�U�4��#.�g
z��r��x�%�M�q&�t�X�/�`/-a�`����
�o��P%��YC��ř����{�COb���F�� ���d�r"����h� *�e�/6w'[%���
�o��tO�{���ƌ��Y���ێ�^v��Kt؝\h�{��7C)9o%Gx�<�qy���X�r����b����]o���9%���;������S7�#R����)T�i��Us,�g�V^���W�u�l\]��sӔ�܎I��Y]Z�ғ#��-���kǈ��.��:�mU/��"'�H��A�.9ZVK��B�ݍ>�{^����kj3Z�ʢ����	QRtc�u��up�"� p*\��.b�^��L�b���>��:�,��{�85��՝*�'f�!p�C���W�4��v.�r�j�u������]�m������s�5O����f7���d��N'7��j�#'�Ղ�\���u��to#��=�jokn	�sIz�ut�*�;q+��ٱ�e��I"o����J`*�k����ΐ�=+�8�嫅u�~G��G��:Ыq���/设��t��ۆ�m����+��,�k�2��,�@w>>�Ŵ���/�~�vو!�-u!�K�^'�b������a�W�n�,����S�9{�'��p(��f��(���P���M7�*|(;�W�I�ͬ�̰���]2��D5��vȍxs�6��F_�Ȱ�;=@��E��Wb�C�=@�@]jX.6��P���Gl���Ӽ��&.|�I��r�B-K;�L�H_�h�'��S~����C�y�|'`��Z� ��{~��ǃ�	���9��ͧ�lX��X+��e�:V��OM�6{�N{F��Ez�,	1���`�l��c�sD�0�:>Bx��[��Y�2!�7�o���� ��o��3�wՑ|��/l��l�h��~}��B������S3���n])���@�>sR;6�.P�:�3����"�

���K��E���u;��7��J��~}��1��f˨����,����ؗ�C�]b�y!W~��x{�b���a7w�dQ�Fj��=�&^�e��t/�,�gk��9�����]���ˮ�3X�e1w�4�bס��ȭ����݁�|�M�y�Ժ�uf�+':P��8V�uGԵ���+t՜��!��G��ش��@oF4�t��vmmq�"#���z��vC���~�p���»f+�X�mʮu�S�RP^U�(^j��Y��Z��	ј)� �g�ꏠr��=5�����y��~�`�g�\8k�o��WJ�V`���tl2U�K�����k`?s���lƥ(tuK|$w5v��v	����<rc�'@��܎�[]a᫋/�T�]���%xW�˒���5�a�:�*�������c\��c��ƤTO�D���I�;�Պ$^����r�F����I�X�,-��ۇ��y���h�����ocӥ�GP/��X.��1��5�U���i�]=L�]���<����0uN:q�o�ic�1����
��]�rJ�0|K���z���K��;!)�hQ}�xS�N{ѫ�:4w�f\�0^\�yY�Xv&�@����^�Q�AC��iBGz��)�3xxǚ��?>�xA�b���ڗ`p�,�J�Fx��㷗� ��E�O����E�}��^����v��P��7L�EV`ࡇ�
��0�j���Y�=^�f�s4���Nu��i̢uT�CK-�bAÊ���Ww9M��1���n�5�+�Ɲ+�CBTke��dw���!�N�MJc�Ͷ���b���^`G
Sv�tv��\�|\�W[ĸ�ξ�\�#x+�vΙ�J��;���Z���V(���-�ύ�죡FȻT9���%�t�r�9�n��v�
��dv��%@�dtm�C~4�$���M7r�*��HZ�2���T�F�!N��P		L\}+��-֝�l�~�@T[B`9so�A�r�K�)��8M��ң'ғ��W�|���XSi�ׇ��cJ5+�IHR���w���0>z�3F�1v�N�Պ�"��-���y����p�v`N�N5)�S�M6�ƩP��u%J��)v���S�a�&pg[�����c�L�W�9�vN�4r��N5�r�,i�/g-th�������Y�����i���$ڱ��4ٺ8��Px(V��|�=Ŵ�]8"á$2���Hl�i��8UY��*��`��r�.�sn�1<�̙;�P����e.T#���Aŕ��9f_$��T ���L�-
��/F��ޕ֪Ql�M;H�P:6tq1��7:�4$�,⫗�S��#���1��f亼j�x�+���d��Pj�E>���r+x�o����"ǈ-t�|����4dgn�r�o8!�|*�rf��,�SVv�j�ʙL��lt��x2rF��饆�f�d�	�F�R�ld�Z�ғ5+i�<���}����6Е�M��)tGg*��h��g�wݴ��:O-:�}�M��m{�0��8^�G)!.�:���P�00�g�NT��ڙJ�(�7R�
�o�:
�
J�41V8��yn��[�#��/�ѝV�O��Q�v�Gk;�
yh�E�HXq�;1��S��$dw/!�1��׮�!�rI�ͩV+V��E��E!c%�T�L��Y�|8���p��qP�]�M3H8�h�6ؓmV�m�n�\.W\�ۂ��U�P�yHV�:�������;\k*�Z(��Wn,o��������v�^����RX0�+�olY&�=J�ŷ��ꗲ��3�ܭeT��EBޭ���O6��M�S�����2fLwv�cz�S�m���{;����Z�y���m,Ր�5��;��:�Ҁ��l�"�����h��j� �
oQ���4����ؙ$�6��GQ�lYr�W��[$��-.ٯ�a�]�ۧ�C�\@��RO]��䠕K��9�R���}�: �U0�-���6[�9�huW���U{�͇�d�'�C4ة�slW�Ý; �ĥto�U�;���UK�nixwr3�<����(>��PZ�Y}�['9�@ޛ{
�g#^r�[�2������_��=��
0�wg��z��p��sbl�,���mv8����;zZ�w2��e�=�t�ov3���!��V�;��|OY*�X����#YJ�Qc���E��T+cTbX*�E���b*�U�X�TD*DTb,���q��UDւ(*+O,�[Q2�12ш�3V����[b�iq�-�DE!��SI4�#�,F*E���"���b�Q����h�*��R�(DDDb�EF"T�")���EE"Զ���aA�RTiA�f��TE"����(��*���2T�
���bSV�QQ�4�%B��,F�0EDF
�V�Ġ��"�* "�U@b�(#H*��@b
*���AQc �.2�Ks&�1DV1TY���e��A�H�UUb"��1UPEAE���lm��WV��F
(V
"�>�������1�v���fQ0���k܄R�DF��G��k�c�!����}WL[t���}���<���G,b{���_ʪ���6�]���4D+�ȫ��˞xt��Wd��Uce}���8�(�xIh鼺v�q�;Y��veRu�|�ZJx�$x�2.Ź��;���2PᲺ��`��]�s��t�Wz5�L|���yy(�-W�6�,��du�&�����1��A�Z'�[wԡ�-J�ϝfb��%�h�ͭ�T��C��}�,X�3K>����5��z�ٗ�n
�+�u�7}�V�Ǆ��X,�7�ِ�*3'[�Ző`�ޓ|ݍ� ٬��x�^�;��E���z[r���1y\]�KX|z(�����קug���������ݵt\�^"v;�[t0(�\�	ϾyJ��R���Ǘ�
���ci���9A��xX�����M�T���j	�sR�4��}AM��-	>y`T_T$����Xz.��<�jk��]��t����{�_5�nT0h�5PB�D����ձ�y`#-L���8ṿ�r�&T�r����	��iTc�{Ճ���U�u��ê�\�g4]KL�T��;�=T���W��jc�����"V��+�;y5V@>�����e�KۚG8'�j�s`��621�h�3A�L9S�����]�,�hǍHw6�W��N�ͧd�+j�Yq5�������������[��CN��Aj�Իo�{��W���̱��a��u��# 8���x�^d������mj<�a{;&ս��#�&1�ޒV�d�K�;3m�W�6�6�.�r��X
�E�eu�{L�x��./jCK����A�u�^R����6mn���x-܋
�-������*���=��k>H��#���m�F��+��~\���3iD=��n�惵Yj���N������8��Zbؿ��I���'S��S�JtX�έx�E⭧F:Xޔ����,qõ�b���W�$`0GSW�O{�ayi(K	�m#��]�pR�/�|c���͆{_�WK׊�jҧP�D�	;�t�I�4���@�~],�9�.���e��vT�n�އ�nM>`�yx�z���`�CrO��K�;DM��f<9b2��XV��;���k��K޳Ц>+�t�Leʌ�.w�+q[�+v���Z4:�.Su�o`�C6-���Μne��WQ��κ�#���Z�,{}��-!�(y��C�4ҿ�;��ꂯl��+����,�+ʒ�q��@�@+�;��:���-d����eN��o8#m�p�C(��$UL+&;���RߕQi���*ᇠ��^���)C�h��X�bX��3�0�V��:�k���� �HC;0r�]¦�d�������j�Z'�R���G�X%%���)�~�7��ʸ����/��YMx'��Z< xxG]���)?a���]9\���"�C����c�����#Ew��u�ڬX��鹝�|�n�G',f�ŐKm��SHC�{p˚oj25�|�,1���!QRt`}ֹҠ�@��x�w7�ƄO���^M+;�w�ҝ*�[2�t4�u=�X��Yҡ�Ѕ�j��L��#�s"��c:�
�Vλ�"�]��f"����feC�|��{킹���KT�yl5&�yTY�̓`��}�WA�wZ�Fr�,�!���R��|�,�L�c����pFTf5����9��2��X���@���G�^�}A2�3[�O�`��Dꩽ~�̵K���:��U�4UXv���\"�
�sȈO'��ʗ�:�@Ft� �mOg�׈�smV�6-F�k�Q�ӁQB9K:OZHo����Jg=Up�`u���S�~2�{��I=w�U��L=�p�i�;�P���j6*��Չ��Օ�w��L^Y�����x�%k�`�{1["�F��m.�+&��"�eJ�Ë��5�,q�>o�<Ս��ֺ�{�u'�b_.�)*��1��c��؈�<M�3tY5�V���LZ��0��A�8�Zz<n{�UR��3ܻT�_{��Ed&_'B��CG���ۋO�py:̠��E���^6a�t|��"��ki����u�!��jvPY�Ad�c���:��C����u�0������e�/Q�6�z��˕�UT�X~�8#!�3� :�j�}���ܺp0`������ndC��y\}�l3��_�$%�W�l���cO��1�^��[�kj���V�RFV��t�EM1x��d⹡�v��/u����)!���Qb���O�5]7;�bP�֦�/<sC��Gӽ�MW#�e�.�t�����3�;nWy��n1ٮyp��W��o��l:D��m+ۂK\�`"F��چ/�e�R�>R�	�]�-��d��x��T޵Yz�mᚡz��l�eS��ub��4�.i��a��\>u-����-�k�54�B|���1��1R�:�.�@����&v�B��S���e��!�j��|:aҥ�4*���Vk�91H`��q�7��
�4b�a�Ȫ�4���F*����Us��@��՜:Y�Yaɛ�<�D�B˨�2:�]��Րiq�}+�����k�@��Q�~WgV��WΝm�\~f�(�9۔�}���Y̕�+�|��ʜ$�F>�y����9�XR6p&f���� �r�,�����=;����ɋ�}��i�9�7��_Q)f�t����ȿ��J�c��k\O�����$���\=��C�N��U�x���s�_U��{!����-�sM@��0^��+ ��U�o����E��Y�t�+�Dx��\�3xG�`��M7��ۢ�������Xj(���*�����0_y����5�70��2kO�]��!L����ӧ����t���!�Kt���z�,���=\]o{ Y�u�Ղ[@��ZJ5e5Ս����k��I�
z��y:#�	A�����f^>!���/�1�e��Xbx�Ϛ�m멵�wʯ|�$��Aej��vj��Ow�('��Ƈ#���'���n�d�9,��rO����P����>��"wqH�u�v��Ix�9�+�L�1�^E�GKU�;;��$�-VCڌ�ǅ&}�1k�U�W�6��պ�IeXPr�|�3�� �ۍ��n�q�X�,}�&,�cz����j����[-�o��]�N���2(/+���k��W1�#p?^�Ӟ��n�/<�\�����=r�TB����>�:U�:ɕ|��3��.���9ٸ�[X��*�[�o�Y��Y�Yk M	D��n��GV�I��\*��'g%_P�Na�,WT��^FS���x7��k�<�ΣΕ5���f�
S��6_���H�	3R榤���v���Vz�*/�`��Qw��5Ω��j\Ց3m�>��"��0-��8�R�Z�����p�����P�-	>y`W���.�HI�����κ�OK>�Iŭ&����{qN��ֲ(t���lWn�	~.R�w���]��H��A�!vt��������(����H����]ؗ�H4�<��
T��]KL�O�F���`&�XJ���,�#W{/K4�?�V�NvOyP��RS���t�WSy��'T�Fs��.Y��t�f{m�U��֢��[�S���,��u�X��.2�]Ԝ
�u�t�=� �����\��3��T8o�������H�p�:��S5z}��S!�L.d���7v�eI��1_����O�0{ye/*κ�.H����uN|�s�ܤ<ׄ�bj��p�OZHtH�Z*���T�XVp��[C@�[N��uê�l�}g	I�qi�/���g�Q#A�L[S���IC�������V^;�Ǎ[5��ӷ�]He���V�x�W͏���1�c�j�Rt =�5��=5:�l�����e<�u<x\��a �����JV>�ݶ6�C��ukr<��ɾܧ��������	�{o�k�8_KwX*)�� ��w33o���R��w{ޡ30����E=\
�T�@�t���b�^B0�xK4�n .�;չ.�ħ�����B+��l�3ۍ�
�fKW")��Z4����w*g�ݹg^�<���Ī��[�IC���7�"�q[�0�m���ѡ2�EOPݱ��E�kB��%�M
7�a��]T�{n�;�-!�C�^˱�X�I,#�6dl�`��Tf�q��D�b����:/�r�%LC�^X���k�9V�U��.2x"��F9k�33M�s�
�œY�����9���|;à�#�h>[�O�e�5�Y���7;���&-�!�s�j�5i>����]N�Tw��|�|ct�#��)�7��mN�F�M�VF2��˦�1�
����K�̝Q+�:���.:Y���㚢��ds�9�Y�b�%@�;� �6��̝3ܷ�V��!SMӶ�]'}3~�L=�a���>N���k��=��j��� U�M�YW��~1R�0�.F�U>!�,.�:�K�^�'�b�t���[��};�X�4���9�͗�@�7�U��z3숡�`���u�f����dgI���d��d l��[ �W"TLځ�}��]7�Pt��6�ܫAp�A��^�'4 �����L�Z�.��iƬ�ò�N�u2�u0m+юu���r�%��G���n���A��?Dk˘SG�0�^"��hlʴ���ϩ3&��/:R����N'����{�6�MRxP�𝞠ly�E��S9��C�=@���p]/"�[����_��W�g�����-�����*jX��g�@��z*ݡ�"퍌����]v4���mc�jZg����O�sn���
�eEPi�
��?��i��u8�%
^�}�J�)���`��z�]f�)}~Xu�"�u�A�R�"��dk�+x\�b��ح�6竷K�Dt�a�YF�0��nX�{l�u���35�*&��p
�lԻlb�tz�m��rJd�d!�m����X%��,툀�Ռ��u�f2�M8�Z�T�2sn��դ�J�?0�;��rP9Y˒�5i�$Pퟟ=�4�*��P5[�kK�|~U�ԇv�����!�;�t��-ªo跥�<ߌ��{;�v�V��f��;��6���w�x��(M9{�Z����/_'�A�M����.�xt�5Mw�1�d�w��f�1ٮyp�TC.�����m�X�����8՚�����2�#�:��7	�Ѭ���4�f�)^�]�3���u)�=CQ/��7�5;�x���+k^{�1��,= =48^�6J3))J�$��dװf�޾��ljvk7[�oIEmtÀu���Z��}/;[�K�=���=�q���?�V*P3��Óh;T�X=N�m\��2���=�4�i��JJsK]�*Y��`���4�
.�����0�3 �\>��Y�Wٱ�<�g���5nK5X,ˈӖ����L_JR�����tO�6�zm¨-	���Ǜ��[���QmN����X�='��]8�_$�9���*�y�OT�}m>W�8(7���Y�,K��a�E�\��9�F�k��\c&`_��2�N��T�6�G�Pox1�+H'�H��=rDp~�H��U0�sf�Z�E�啞���m��m��.�]*�UG�����^Z�w�`��κg��[�b]x鉤��L1aj�,ڴ��8ld�Q�L���=��1&�Y��8:ǳq�g����p�;[�E�>6�5���(a�\3)t���~�6���2p����p�]��5m� �x�Y��3ʵ$���c��+˺�ޭ�^��L��M���ׄZ:l�]B_�%"E�"�N;�6�	��+u��]UBN)p7Vտ?�7mպ3v�A.�)+t2V��޻X��LcWp�UO�-�b� �������W��3�l.'�&9b��Yc�i��qS|E���rf�7%oɁ�2lF���_g�[FgL��Y�=�����xY���w�$6X1U<v�N�^��f3�i�v�� ��[;����ǂ�r�"-y-����=�!�/)����aX�5��a� �Z�`gIpf���CJ�N�s�m "�ѷ�q�z���d1�o���
͔��M�a�(�w�����`����{d(ȍ�
��X/�� �ݸݜ�uËX�,>Λ��x.�� <�=���,tT����}B���Ș���F�ғ�77�vR�b�eSC�'M�̕U5��b�OڇE�lf�甩|�T���������T��sUa[��Z6gn�WL�חI�|=��87��������,
��I���]�����}N�S��c��˴wK�z�>2_j�6
gZ�"�N���6���� �g���켲]��H��q��ܒ �hl_s��1w/��qi��ޡﱊ�Ճ���U�ZA����M�E3���r��zo���[.���թy�G�)�c�zY�9�3���N������2کOZ��k԰�}'$]���o�P4�d�(q�m�ꈼ�B��b׭�)��8���ϋ�k�t�N�е��as�.����݇tiVQ�܄Q���`>��裸6�oh9�X2Qn��\�o�R͕��:en���˝�ݍ(��f·��ymE��g*���vCz��Y��X8P��-7ҕ�~�)V|�f8�5�+��+�*ut�qPu�;b��5���lh�|�^���Q췝!r��Rٴ��9u�$v�|�T:��\�X$����X�(��Mb�ˁ�_wPt�9c��%a(�Ԧ��*����d�gV�s68�;�ow*�k�F8����r�å�
y%w/���<��������r)���N qq�eDY�Sq6���P��t�g�s��U�єT�#f\�CiSg*Vտ�c`��:v�7V�4;$e�ۄO����ѵ�k��;��a��(�/��^����p*��(ޛ��0�X[۶��/�7ƞD�̓$���pjb痉ֆ�+���ka�+�Dmۡ��\�ޕ�=�۴��zL�ָ\�Z��ڳ��*s<[�H(��X�&=Xf��8�\ʚL_@kq���a�$��}ԫ���|) ��5O�>�ᷣi��4*^�%K���0�2F{U:զڢ�<����N�o��X��lV��݀��S�O�$�]n�|��#}s@H��V5z˜�3Xv�}���KS8;���us
����ϓtt��MF� �b�˅��D���-s<y�t�k�)}�-�K�΃yʼ�l&�N��%����劲��?ne�AۣM�ե���!lh�.��o(����U��h������ۙԗd�1L2}��(�f�#z�B�QaGqj�1��edf�9y˚���.;Ɲ����K%��И��n�̔&q����,�R��Q�tT��m�,�(�U�J�j�G��z�fQ���S�Ug-%Z���\�n5\ܽv�<R�4������Ҟ�=]n�s���X�c��Ř�(X�e�!�N��z7���f�]�Sse��͘(LN��d�6��8���^YY�����w]A|1j9�dw0�NR	����"��˺2�-����13ܖb�[���7�=ֻ��r�\d��p5�T�:|I�Ĳ�&3y��b����C�YcWABl`?��5<�y�=�IW��կ*f�p�:���y�iis�wP&f�.o�#Ϲ�a��V�pd9���A���<�۾QNԡYgKi�����^^�y�oqkn@<7��M&���u�a��.z��d�[l���.S��k{��jw�����`�VΞj�(�^�Gs�j���eh�r�D��z�R��0���μ�u>SrT�{6�ٷA�!�Z#��M�4�ywl�dh��X����䮴�+��	ͭ�κ����T��Y0�JSro|h��Cġaا�kT����>��5Q�4V��M�{����ۺ#�Y��o�>��@�q�i���ZPt0�o�e�I�;�������j�w%gjU�< ��G����X����(�UQU�[J����r∢�IV[V��� �EM5b�4��j�AEDA`�c#2�PR"��T���1��*����aDX�E�\fcUY�YU�dX"�*�r���
"�mX��`�
(9J�E���(�1UH�cUU��2�q�J�R�b�Z�h*)�2�q"#��2(�����$�DX�b�AKl�h+m*V8��"�5H���3TX���%eEX�,R�T�����5
��M3I��
�i�SKj�Qb�je��k]YD�(�Uf����-�DY�**e�h	�1��U�q�1%T�e�Q���Y+�l��lкp�KИ�C#5EW�69]�,?vK6l�a�N�t� WmXu-SU+N�p��������9�b���!����ވ�O{�#��^���}�wt�<b�p�ϳ��&�h2��
��~R��ϕC������0�xݔ<�;q����y��2yu�&.�ʓ�TQ����o,��Y���}��ۍN����<�<�3�u�FE���b��b�>�Ic�H�Z~|)��c;^:����;*.�ǦV�6���'gLM{�5�9%�0�ۧ�b)�a�˙�K	�m(x��23O)k�Z��;5d�\tWY�|q���Wک�����R$rę~?R�0�ʤ�)�z��~:��UCxw|0Y5\�2Cf�6�w$�u�3R��>���(��n�*�!D���&cP�9�����+��3r��g����Lxe��Ɔ㸓ܨuGf���Ḳ1�����h�:��7�tn:9���H�u`�{n�;�Hb��(��~ݥg�՞�������`}=�.@��l��`v}2��.�^ů��銋UnAU����t��Y�ʄ�n!H[n�0��/���q����b��4-��&e�5�u��V�ڣ8u����{>sw���v)n�=�ۑ.7��@��&�=�׺"�x��Ř��ʪ�S����X�m�VԁX�m�H�a��΢��k�P�7�%���=��
d[,�m]�7�ٗ��%O��EA��1bҡ�e�P�/��wɺf�9����t�ɍ�"�ܶ�t�{Q�Sާ �7J)u��<�U���)��T��o{՝/���B�]�0ߝ4��uYP�����=�aL�}*�W�!碮ɸ�o�HOv��f[�8�Cէv��h�P�͸a��ۇ�P��o:t<0�ך�Y¬3X{�l*eH�(!�!�-u!�*_b�I�����p�|�zE7ύ�x�HE�w���k�ֶz�3ҫ�i^�#/�hlʿ��ٴ�5��v��ݡP��f���7��Si�[�yV2-�q��\#��)܅2jݡ�QLe�����(�ã!p�JH9G�fÁ�b�R�i�W�~�s�����3�!~�m��l��DE�fv������V��K�I�m*���'��1!Pe`:{��.���m[���1�
��R�!�JYz�.�Q����(<���&eLGDv����C�����/M˪����`:�}酽T�K>���^ �����׼��_�ᗙ��Z�ڦq���{ʶK�K\�Qy�	)::�3owF�02i���4tg��bȔ4	��^���Vo]�:�=s�#w1�����]��\84��>C*nɝ�S�󛙯L�V. �t�n��D��,���4D�H�s��]�h��Ū�a�� ���ə-�`��@�8�l\��Y���uZF=���:��o�_����wb��?rN/E�qz���]�yU��J5X�k9m&}yVZ��w��ќ��T��0J���TG�n[e�=ܜ]ɗ�!��T�>[�/�H�����O-,��^W*cN�pf�rm Ӫ>����&������݁���ǽʴ�d_`������;�kC����o�V�P3:�rv�w
����`0ڹ��L�{�:q��(1�c�9M��T�a��� ZO]4�26�(Q֢W��5�نÝp�)���u���ܠ#��S�����^��CT�9ltY�����ʠ��m�+��
����!wzT���	�ۄ�CQ��\�N �o����[�d�\��Z�t`��J��b\��n݀�l�);��fۃ�gF:�or���|'���Vr!�հ/��OybJ�0|K���C�Xe_�uSo�ь����E˦gr*�w�0��o\�yr��g�a��@�l�$:��z��qʹ[S��W�m:��%p���D8q�)�~��25n�s/:\���|O�8�F7M�b��KǗ:�5��@��=�n0��cv6�mj�SAvMԒ�mE�P��V�c���f��sxӁ�`��ǹі�^j�G�1
}\����g�s�����, �O�VVKdplA�ݓ�u�&�:|)�. -TE�V�4�����}�\��#r��@��Ze*]�=�bj���7����ӧ�%E��l�!\�����+$�m���4?R۰ ����p�]����ki�6��r��\c�ڪ�k�i٫.h7/s�Λ܍Cv�G�4�zvw#E�n�!<���D�|���go��ﲷeM�z�̙3�^����e�T�APn��1y-��'��伧�N��vk��"�L�=ٯ/l�k�u�{ؘ�Y�h.�0
�p_�^�v���5��y��پ�L	�w
�'z�rpU��<-��`uW5ؕ��y�]��ِ|�n7g<�p��,�۰8`<��x\�|QGi�<��A��EA�+"b�ꖰ��Q+�6L�0M��i��R�z���s7�=�1���Mc���X7��x�S�R��������
�M�Ӷ�\�OJ���JvT0A�ͱ��VN�3C���$YhK4_W��H��b��2�}A���[{�K�jg��:��S;�j,i ����07Oֽ���w�r3SUwj��������xZ����Ff���[���8�H7� �Y���F^0�JE��ү�A�բ����Mo#��&��)����V�\ۣ�W#?��¸���Y�T:�0��t8�Wn��K�x#Oò�0%C{��y�A�u������L��0���8/L#!oTb�{Ց�l�c�bU	�8��͕�D���j���X5��\�}N���:B0� �^�|-�x0>�l�w�6f";R�}L:��T߳��2]i�Us[��	���:Y!�z6��E���X4딝�-I�ްyV������"����D�hB��
��4��j13���p�mR����n�ly�rV{��b�Ʈr�,*xS0�D��.�/�db7�2�L��S�0{y�J���2#����o�bت�����Bb��S֒<��W/����g�����$�&s�`,���kiR�҆��Yq0T��S��^ZJ&)�FjŶh���Yy��r�B)��d����QO�P4��( u"#������!Z;(���~�_�zeP��:ʃ7��Pe��5���T�B��z�<��kݢ�k�Jϴ��7F����O}{��݇e����`]�J���:�ح�W��ֻ�9�W*��ËE;���VYܭ�|UgOA���@tV�q��Y��M�N�j޾��&�8��F�옰2z��
�:����$C;�G�/�d{0WE��p��T3�ˠl�w�ICLnPȄχ��K�6��t��@�㽌5�%!���h�p��P������o+��Dor�|1޿UgEJr����g&M9�ڣ#�St��f�1�R�o�v����g����ze@3�\sص���+�U��ח��������L[$�˒U���=9`:\]��|y߯�+�:̨��W��1���o���W[)`3�+�'9H�.!��l?T��֩�S�C�"�r����un��j���#����@�鹴�ن�^�{8�9@�'�f��ѝFf����`3���ܞ�ll��b��W����w�Q���v��|������n}�P�s*p=~�9e��Cܟ"P��)�v��f\>*$��gPC�_˩��ؼ�t����Ln�b���ż�h��ڻ�|"�w�d�k��'����wJA��e�@�2��v�̬��ƽnSy��H�̨��^�-.�{އ��tʳ��G>o"��j�
w!L��v��K��u�N�4u�ʰmJ��Jf��̧(wR����:��f>���8��ɕ|�.lÖ룷�79{I�N����]]��w2���hm�n��e� a�s�='p�Zy@l�/��Ǚ�#��ts6��1�d�'����7/�V�m��0O�C��m˒���M��Z�6x��E�n�bX��T8.T"Աc�����t6ұZn��c o�}�s�����7��xo¯
ȱY��?��'�����]��oh�:�_�ﻃ�W"xA��s�k���~�z�3I��V8<��{Ƀ`6jj7��g�u8�=�9���~��F!f�qh��٪3�K>��g/g�]Y@���[��>B�'�Ў����ph�-�-�a� �"�;�P�Yr�\f���LFA���Z�����U4oUI�9E@͜`���o�E٧�q�>ʥ�n�gN箐��cye�}�p�U�	�j�X
���+�:��r�n��;��)0��_m�M�b�EwB�8�Q��Ӭ�37�9�u��
�]��ڲ�߳jD|�2ܻ9҄�:k��[^Y.E�j�쫂y�Y	��*jÍt��Y~�5Mk� �u �iԤ�R�	�\/8偺�Q�ݺ�-��e�̍�91��uժWAW�}�D��M?�نÝp��s<�}�Vp�yJ"�񫺾tXktSr��ض���X�����3��8����OC��ͤ��"�1���aÓ�J��ͽ�����VK�+]śLl��L�7����w��M3z���[�u*����^T֨�����ȓ�����㦢��ý������яmƾi\�Wd��+��͖5�z�`��f�竼�.	6�i
��X��_3y��V���Q�n��i�Rc\Wb6
�ޓ=W.�Uk>��v�Q|�z��<�&���]ګ`����P����w9՘G;�6
��d��2(��Щ�|9�W�ɫO9�#\:�5HA*��̠�Ʉ+���qn�eg��Q�yСJ���/H[�ز?d=(,wXy��E�(r�J=պ����2�j���	�XwT���k�|yWfη���C��C��@���xI���ӧ�����}q/|�h��𱴌��殦�w��Ԯ�׹S%Xc�ԉ& ��Ѹ��R��բ�;g����\�UQ*�Fk��fU��H�,7�U��K�$�t��z�|�ZJD�8��܋�6��0��Ԡ�������IB`�j��r�'[�ר?�!��z#�޶��0�>� m��/��N�u�	�M_���j����L_���I#��+t�X��/�M��dۡg��f/A*��V喢�[�N�BT��o{x���;�m��juA���W��{��������a\��rQ�Ҟ6�W�>u����i�INn���M�����:L�fm:�Z��7�7�YJ��W�d�vެ�Uy���M�m"�ܑ���@����ss���
;kC�v�l�0�ln�����ffzg��+����R�wj�a��|$�f��Z�˵�����J^8E{O[�$5�0f��gXm����U��p������t^&��\�R�ʥg!��B���ei�v>�{��gҥ�X"f�=��'o�����$��W��ˆ>}RV����Ȼ��i�V��sW�z���;��`�w�0�������ÂA/���W;���LJ�=�����Բ^a7�i�/L���|%�P�1����!��/������%"�6�]/.zq�#\;����B�-2�iz&G����zY�9�0`=���v��n��k����~���:�z�J�����k�a���f��j{�x�>��F��z�t�������r����,���a�&�<*��`��u���z���t
�
��>�z�ZTu��ͨ�)R3nէ82�E��$�減m�X��
��:��\ux��M߆���)�::�i2Sv��������C��uN���Y�
s�mwg����Y����X�6�}�	s[�D_K��r�0<����n�P��tfMn���1H��'hu"儇a�����a:`^Ϻ���sf�mgLf�_)��UUG/:���d�<jz`��.ظ�Uˌ�p�LS4�,��%��#�uI��|���i�z������<\�ݸ �^�Ly�/�;���N���~n�ɦI��\̰}*)d���bZ��f�Vh,4�X8u�o�+/����V��]�@M�H�ɗ�)�A,k�z���7�Rg�1��L;�nz��!g+�=��m(*7 )��f�o��3L�;+n:z��!���3�4�ut�f�[�t�0A�Q�ʌsq� �����iHחW5  �=���p/mh��<�x�~�3T�Dorʦ|1�{w�Ť1�	��ib�3��'C�fǭN��F�.���>Se��0;� �hl�rk6i�0�IT�It�ͻ|����wQ���M����uc=�zrå�^^�qW]��7.��u��swrG&����?Vs�R���i�O�ԉjb7��#4��dkV�V���G1�\��V�����MR��χ/���V�����%�C}���,�{|{e/o'�շ틵xZ��u��0]�W(B�q��B��\��rD���'.��:�yM����O �4N�g��gs^��������umƔ�̛�X�|ib����
�F򊝂�rWM*�v�l3z��&�)��5�t�q��᎝^NZ�{+�#�R��r�Q��q������E��U���g5�}F�g6���G�^����]/P�r�e�5T�����g��\6��yَ
�|$�駖�+F�4i�B��6�_]l&|0
4�n�R�'#��zbw8��}"�r��r�p�p\t�{lre��OW9�Y�G+p��ǣ!���GPd��Vo�K�Mc�ʗ�d�/s'n�ٵ&ܕjə�w02�]<k�X��hl3���#�1\�tؠT��#ٌ��R��s�5�0�:� ^EQ|@�/ZT��gR��t�������ךR�G��0�|�-�%�uƸ^�}�����=���G9�n7XA`�C~T��9���&�C��r15��ݮ���V����rٳy��O�9ylee䒯� ;��=Z�e�%WPR�*냶�m2���GE�5�Уtw{]̧�]�Xv��]��Z���L�
]_Kh�.u�+�E�;!d^�#:'4剦�-�]) 7�A��E��בe̓$�nnN��^���F,;WL2:�PE7s�T'�
�\��i<����ł�#��c��Ϋ����+�]�ʥ$a���r��{Ma�'Vc�
�����0���ګI��nG��S�vt@�Q$��Σ��W���*@f�d*�k��n��woK܍T#����Mw2� �m)��J����Yy��C5J�����E�@�8���%�F�թ��e,�&��[I �kw\g`w;B�CEm��=W�����̺��Y�۴��pn�^��U���i�z�ӽ�BJ��b��rq<f�$萛:�0:�]�KP��3��8`�x>�k5Ri"�u����)�u�Ǝvjo�(Y��2c=p���gG3�Y4:�������@���攤���
U��-���F#�t\���&�s�Zv�
ܺ6�f*�Y�é-D�{��2KPm5�5������I��ͬ�x"���o&�b��e�O�9�S�7����;�"�]��s
`,ƠۤU�9��%�t_S���C����[uq{J ��4N��4�\j�O�]^cn�@Z���3�	>��
���Z�+R��3�
�x��~]i�}%�z�aWz��AM(��rj]=�2ֽ�W�ۢ�ה"/�K�ė�6`T7x����{SCo�q��7��S�U�9b@�]�xY��w�sؼ�6@���r٩˅?� W],�V~Σ��:�9E����F-z	gt	[��84Kt�^νz���]�[�����v���ۆ,��I��{HS�I�ey�8�S�)��P�Ջ�.��{�����"�}�8��%`�1�[n0(��X�R��E�ɉY�P1+-�V)-�.P����̩�a(���Z��"T�\fam&8�Z
(�U*ҭUTR���D���������T�*�1��(6�m�E&0�1%�[[AQ�"�ņ%q
�R�PX�r�TSl*�+�-�c.�Q`�j�QV�ȰP����"�����Z�(��ʵ(��YX[@���c�1b"���H�E�ҤQV"X(��T�EjEU�)Uk] ��RڄQ
�D̦"T��Q�&f`V�X�*X�*�UZȢ�+he�*�	YT�B"e"��1s
�+*���J�-��KA��al���j�h�  �}��;��S�h��qsW�I�t�u;R�sɉ�����*9�ޖ� 3+U_D�܃��8��n�rZJ����SgR�{���L��+�3���������m�����Ssm�,��U��ѧΰ�;�6��x�sPl�v�N��.�M�PA5�\|��O��ȴp׺����*:f�8\�����>n�,���{fZd�h�F��"��~+�U׻ �.���]Nd���*Xw�X6�U��Q�[1P���pS�
d���z;#�W�>�ǻ�r��W��(�t��`fm"Ϸ~2ķC_��e
��<��ᫎxX��y��peۺ�<1-,�h�_���2�b��+֞զ }�8E�Pm�n"�;��Y=�W	T�g����6�+Q��]ç/j�'���W��o_�T��dR�$EJo�3�I��hd8N�k��T�0:�eS��m�~'K2wM�^��"(0��٣/��&���u���2%���|�'�-�`Ü��@��V=kK�{����B��07Lc���o��"k븖�Y%��N��C��f!�E�F��Y�cIڳ��8���
�*<��vk/��9Wת��vd5qZ�l��q�vp�ۛ���d�h�o��.v���2���{�l��"�U�t㮳2 r��Wehե<Vq��}�T��IIS�B��O�c�v7�s�p��ڻ!}�ιm�y|�`ϼ��Y:)��X]�*����m�=�ݞ�Z��wՇD�e�#~���+^�z�G�L�HC�!�F.����!�9�܃�����t�5Mw;�@�\{�J���d�7��V��e�NF����|��rk�;C��[-������̰KP��X���s�������?����83�P��~9�K����ZO]_Ν�B�����.r����w������Rˋ<�vud� ������c\��`��f�繿��0f��s���ҕ���h�۱���=@�v�������y��q�2���B����jr*��N�C6�OdJ,�{j1���Uf.%�y^At^i�m[�V2�#G\W��0-�re�'E/=K�)�os==�0�po�-����%¬?�]gs���5խO"�-�,��[UUm5��<��d9�"{��%��]�P�vǩ����>�^:bi�,1��"ڜč��Xwk��6���⸐8����焟U���U$�,(��vuΌ�бq�X�WR:�N82��bM)�����xh;�d]!��%��pK�N�,�t4��l� 2�B��l���Z6��R�wE}����W1���4-��jo0�67yj��]j����a�iǮ0�r��ֺn�jq�\^JJ���mLޱ�2��rE���Ǘi�J����=�����ǝ�r����7���X��5t�i�c�k��<&?S=灖������:`躪p�yXWjJ���u#�n�>K'���Xt=��u1���Ȗy]���M8��*k���U���@o�T���U;7�6!�/GP��Mv�է�a.�J�w�]F�Qyh sv�1��MƫN� Fy�oD�5S����'c*��� �<1{sG��E�,Tܧ�
Åok��M�3�3�FGkfCܨ̘���A�~�{��yr��[���,��bϛ��P.c6��Wחl�1y\]��kJZ[������Ov˦��]���Y�ܸ��c���X7�Viq�A����|5f�h��m��~t�]���[Ղ&��xX��d�l������%���h�ͻl�°o#Y�P� `E��.�=A�u1c	��"�N�����q�y1�x����u���Jy��t��q��ߍ72/B����/L"�{�<1��՟t5ʳ	�,
���j��L��u9m'Y��x.X-l�,Ig���ɦl	9�t+�J:�V��A;��Y`�2T��J�7��+���IVL��Q��lV���U�MB���.r8y�}- ��]���+������Z5E�Δ� ������>����OP��oϣOÑ�`�^Jf�!c)r�!�i��8����ם�Uk�'Teo�u�>H]mW��rR�T�k��3�w��fV�W�6Ъ\�� d��ͣh�V@��|�2%��Ȱ,�� \9��LT,�<*���}.�Σ�;(Lېw#p�i�U�lP~j����f�֭���O!�u�d�/�q;�n
�lT��K/˧uj;c�om')4��n��]e*�7p�Aڃ��bjR�Be�K�=<����.�s�N�O'4k��; Vx�����Jڕ�P�3w��4T�������P޻ȁ'J��o-[T.3iAYUe����!�VV�p����"#;}��p�^;�zZ��I��fZ� �?.�3���6	�B��a�{5q��H����xf��\:r�x�#���w")��5�L<
�ut�ȫb2��(�˕�Q�{L�J���%���fb�����jd�ܴ:q�h�p��PZv�^���]T�c,�,u_
��5s�#]�B����;Ql� Lr�Ⱦ4M@��֗�-�ӱ�W���M���OF;��Јҝ6�oZ�6�!�y�]��X��H.����Ce+3N2�䬠c���u�:�w���.Rt��+����VF��+�WyiX1`�z��L+	��Ϳ�\�H���R�t}���������]���6Y�0;� ��n��Z�U�R�{�\�=2�k�V$*Ｔ0}ʮ0�S/�4';������W���#Գ1R�E�<��A��5�MC��½MeO��@�Ƚ�n�@+��~�Nm��s�f��JA�^��Bx���6�`��^�W��g����Ƙ{�]�<ly�K�.p�t4�u=��v�;�b��gNLjܦ�1�=VMx:��2�(+��$*i�m���Ș{���Vc�L���쓶9A��
滥�1�.h�L��(T��	���B�<olMX���g�q[s�.!�0w��g��Yn�,������hL�M$az�A27}�8H�/������tt1���o��kx�m�<�n����.�u`�r�x}Ʒ�h���2���C�E!�`S�$ha���J��v�5b�����fų�gTv�o�JP����
�8M�8����7�՚WՑb>�B�5e�ƭ�rԕ
�P��#Fҝ{f�R�X7vd$A82�{�N�8�p[=��{Q�����]_N��jv�/!�N-��[�!x�l�Rk����w�9£��Ro�):���{5P9����u4��#I�p�����M:�mj�X���#��ݵٵ;��x�8�����?�Akg=F��9vƋ��fԈ*pUfZZ�0�K���������f�J�S��Q��Ȭф�6����W�J��V֏[:��m-�G}�U��O��fN/�ϒ[�s��qo��3�wg"�0z�rv�@vjB/յ82Q�Oݭ�[lc�z��$���s�ZEl^�@v/��l��ƚ�eRa��3-@�ݫ�\Y�uByOT�/�l�c��ł?$*�ێ@jny���k����ud��X����k�A.Z0��-D��
H��}v�Y�!@1�M��A�wg=���<&��՗'�t��'uokw��1���Ӛ�f���7'݋~`U��`��:���l�u-B$?:����/T�=\�DVc�~���b:��\��xaߜȼ; ZO]Xt�2=^(�Q+�=3^{���G�N��oe��b��[9�+��͖5�C9l9�t3�1|}A#�HW.��Þ�}�czm�o��"����eC����\t��x�CxX*�4dB�a��z7���Ӂ�f�0M��l5�hRtf��%�;w���ӘA�jM�@0Tj�c��q����u^-pV�6D�P�{(	F��6��͠��7{���S�R���uaU|q�}��N��<��][[)t�j���ɷ���Ю�J �KNS�tɽ�޹̹{�����j�N�e`2��úw7�� ����}7�^$U�c���^�괽����]l�
��GU�x�u�Z�3��A���e<�~}1���o���C��;'��bZ"�5P�SA�y��1�&�0�������^��6�R�K1*��*ɣH[�v�>�Hd
O�<�����i��\GK��-��Gxߕ+�fv��ܱ���:���3��~�HTf�\9b;$��������M~��v��貹�N��b��=����}���8�(�x	-������@A����Gs;:"�6Q��:_���t���@�O��Z�u�R���!�n�UH���H�뱺�nQC�oٹ���X�@��ԫE��3q1���0
�� �?\Ҳ:Z�Y�����ߠ�v�J)��6Ζ.�P�,�X0]#�5��u~�aF{kC��``��l����C��l��`D��&yN�p�,���n���l�r����R�|+<e<\"����=���j�B��t���8+���]]��.��o����.=��]��'�oF�pY�A�U�����f7�m9��	�>����g(����H����ʍL��WuJlv6��+��J� �y*	�Wc�.�u�&���6�8��fQ���8f�ʁ7�G��Ļ�"qW8!t��x��܄oF��7��ǦCt���Eu�o%��R|�P~^Xe�ʅ���ի$kS\�r�W�*�Iv϶���cq<,{L+'o������N���� o�v��y�����Y��%2M�-2�]�^���^�<|4lj�ډ��F���Nz�����g�sB��=�89ZmZ�$d5�PV^�G�!oT���#�TjW�;�D1��ݙ��ONL1R:`ꡉp7�=�i�v5��k���
���hC�i���S��9�3;7��Õq����[��)��T��)�S_���.���b]!ّ�ǌR�`��g����6�|�w�s"X
,�ஹ 1,؉���~<*��{3,�9'M�IO=�I˰�����8p����[k�r,8Lτ^H���]r^��F`����(��e>�d�=��;�!)��[Ք�3����P���wd���`�[$��$q9{��{x��'�
B�`>���;~���㭩\a�f�$��/��=�L��(�u��5�v�n�S^p�|��ctu��7�YpP!�6����(����9~W��jG��/�<�N�Q�eo��y�nYy�y����oøt��٭K&|%�Q�\�&s��oo�b���ȕ��#:��l�|���M��b��zB���t�c�ԦF���V^+,�nE����U8@}�@�����D���_8��^�}ޫ2�!0�O�0^o��`uv�W�,�·T�F*ߺ�
�<Rvd���Թ�ú���<����֍0���F] �r��˃���B���L�K˹��l�����:Z<%�q;7��:ѡ׹pBm�A���ޯ*���υ�s6a��36=+^����^�y�dZD�=ʡ�cM����>Se��0;5� �Ypu���ھ=����%�}
�P*|�"�����_*���}9Bs�,�Ѽ�8��c�qf�:w�u�#DY�l�fK����L������;HErۄG*shf�s�c��S�t��55���0U咄8T\��s���up����u���1eC8:Y�=�I)c;�c��c�rib8��YΘ�dׄ.�%u�!SM����������O���ϧ-�����&F^_�����9I���S����'���>�T��h�g��X+��-zv�\R�e��˻���R�9�)��JS��p�jdҨ\��J�8�cV�û3v�mA*곎��?f�u��T5:���fX��������2�&h�}Y+�[�U��s4�9�[{�D���R�*cN����bG�c"���.R�X�l�kS�{{��w�|�X�űB��p�Ou��$�/����-bd�h�#�l؅�*4�����V8�)����jLO�`�՟#�M�𿟗{Oʸ�f*y���+)9�.[W�Gr��M�	�Rz��T��4ƴ�A��i3��e�n��T8.T"KLs�}ŭ������C���<����&s7�u��`�CUdX��x^��1���v|k-ۧNMSy��Q��c�اvD>�2��)d���SƩ���ڑN
��wH���ѕ��oz�;�;�a��	�Y#|���tE��a��;(Ӧ�lE�d�b�1���jQgN��i�^vo�7_$���9�ό8����}��>�8##��ٴr&LL͕��5y�<Y�r�����u�a�c���w��"��M����|5�֫�çM5�r�E���*�}^�M1�j�3������ȋ;���+u���G{;��y���.I�/��f�~����V��$`�7he��!@>ͦ��e�.�t�1�����O�)/7�xI�i<t�Xx�rᜠ6q�6zj�nN��1)ME�э��@b6�Z�R:{ R�΀Q;�'¶���7����M�՗���W���T3-]ؽZ-�u5���rP�F�X�I��nL�3�nn�w�"!��^�_:f)=�jՍ�:���2;��)�u�p��1��Ut��yFns25��-}�[9���j�`�;��]�^M<8��ӛ։R�[��Ÿr �Z�J}OY�����Pk�εHsfJ�s���gag3��8�����ދf��!Qږ��5R�7�G^Ʃ�Y�x�%<X���C��r��ⲫ�X�d�+�r,1^��7չ��>�Իo:�8UvX����M&��]��Y��"���Fi�����l�7�*s�X��6)W+���|PFʚU�V����4���y�%	�*�X],��:�c+���ږV#�zɽ#��&������Sɂ�"m�����&��{�\�ةS�*XR	�-娤|���t/d�����7ɿ^0�������i��������fޜ�\G��^kC
D��$M))�؜tA�U���b��E����x�8Cɻt�,dH-�>���R������;â�ٯ�%�XSPY��`����E=��-Rbk��Vx��N��o7��SE�0�7C�VК�)S�A�p�E*
"��m�M�0y�띉n[Q�Z:�����j���,tv	|�:�]������i�Z1���^�q�T�n���/�2;��5�|�-]�C4���;%d�W���Tد��c���4O_Nѫ~�un�2\�>�5:]ڹ9�������d�o6��yP鍾,iV�c�>�w/�Q�j�_]�ˤ��`�vޜ2^�ƃJ�M��P�Y�h�b�Me\q+*�lh�n���-�+�c.�puh��Iǝ�Y�ͅ��o!���I���R�����+KI�[��'\�QR�:�I�Wn���u^Յ��F���N�Uw�Y�a���>�ه�=5�}b��&q�5K�W���U��kdT<Tb8;[Ru{�g-�2R�ߊɒݝ�}�4���R��r�r�۲�v*ok���kЪ�̆:��n�Q�����nު�H���,L�W��]Xyc0l���u���'�����v7�`�U��i�i�Hfn�fot}�',�1�t���+��	=]H�k4FʽCx� �m�/[�y����ٹk46�	b�m�P�W��7��4����+Jm�\����ON���MY��Қ�Վ�J��jv��2�2ٚa�iG�uyyO-�Dm߂}OK}�kn}�b���G�v�r}�\���]�u��4�"��\k�UZC�P��Ԥ6�nko����Q+��A��[�+7���,m�E���z�ZfT�l�%��HTd=�f��{�j����̽=�%dJ���A!�NL��r=�1�)��~<ןy���4�q�D2�Z���cD�����j�U�eq�%TX��\�-[T4�)X,++JX,�˘[J��QkX*���&[E��-V�q�b�ɧZ�)Q��
�4��KR��QKlfR��* �DZ��D�[sTb�P�YE�h��Km�����J�`�[kK��+U"��ke�
�FTl�(�F�Qk* ֢����ʖ�UIklq���@X4�����բ�F��#E(�X�֕-�Jڂ�*4���Q�c�M�[h�b�P*�b�ՙn6�)3)Vڮ5���lh����mK-
"V�㌥��QE�q-�-f4ŵ�كl������u�К���F*U`֘�-̠�--cK*���[T�3jF4��-���9p��1�5�T������rس(���*�f�Lp+A�j"
,m��KEEִE.SEP�j�����o���6|5��Gw�J�Km���$���q�O;�	�[ձb�B�p�Pc�lL�^F$�%��\s�ol��9b��+#�&�p!�K?yd���K7��ˆ�*��ɨ0"b�ڀ}�H9�A�(,��cX4��y�+gV�AJ�!�j��o�[�Ɍ�91�:]_�+� ъ��֢Xp��e+һqFm�\�R�p�i�����⽜[,k�g-��5mUOo��_^`�x%��KĝH֣��^�:��x���YW����M�M�yK�����[��TY��R������C�?O99n#�^�*�NӪi*�4�]�_A㨹{y1��j��{���H�v�v�G{7w4��
jT�c]rLJ� ��N�KH��u�Z�3��A�������sltG��V�w�oڟ����`���^�5�U���8^�����[�\mg
;8�b�^=*��͡bUbݫ`ʻ�Ǆ�*}�m58��u4���x:����Q1��IqS˒�0�f�0$ς0.���Sd81��d��Tf�\9b��#�G[��;9���!��q��{C#��X�Cj����l�`��X$�pTiA豢}@U��*_���S{^�Y�d��n5��8�rHeI��Ռ�)�l�/N]d��j��*�d=�s���,�^1nm����
����v��S!��Է�c��R�o]��0�*Q��4�󻅎S���5��ۯ&��-C��&	p,=g��uw���C�l���(-t 9��F,K�v7�y��GKYi�V½��'1{���]��(������|���*��<~_ٺ�_���0
�pN�-�A�Ȯ��q���j�%W5.c1e�3�`�0sU�+
L���\o�M�5a�(�z}�W^Z53˚�y���,��)ѫ����zLY�v7��I�ͣV��*�9��թ��/]ݚb{4t�1�3rT��8�S�P�����m��yӺ���_����S�W�*˽R�(�>���=��5��_sZ9ݳ�og<�;s�Ҭ��hvC�
H�ima_E�N-�cWv���OW <x�W]����ŻC��(t�#p��l�k�HW��u��JjQ������i�vS�v�	�*�o��L#2�A�(��Qw}YxAEx�^a���W�v<J�L�u�H{ȯ汘.��%��`��b~��s/7U�#���,����u��^d��9`0y&�o�(=���L����L�f&����]�ۈD���up������n�[��ܼ��0��^[�ҭ�,�P�Kv����憲,�#Й�hk!�aXg���^т3ͨq�!���r��:��S����	5�LuY8l���e`Ƀ��V3��td��N�b�V�T�ݼ�Tt���A^u�_��)̣�
�a��s ��A6�ҩ��_���z��o��Q;�P-�q����B��+�n�XpT�l�輑9�ې[��KIL����A~l�Ǹ��C�`zlm��kj�C7�D=�n�惵Jv)���%֨��p�y/�5�2�VH����;�K�:,`��U��jW�C��:$�FrTգ�s��t����d�1*���^ZI�<^���n
V^.�a�u�E����� Q���#n���c�jt��S �S���^�����߆�ڨ�"+��f�-"E�����ܧ��.�j���~s�lɆ�DT=:b�kF�yPΣ���lF_���<�5z����n��`�X�\ �5`�|k��%�p��:ѡ׹pA�ʹ�1����܏`�8|㞝1l�#k܉�? eٔP\8��o�@��6Y���Ĥ�tnxu^b}���Y�ܱ��P�Uk$�ظ���k�5?����//l��Q״�5{D��a��/|w����9��N�O>~
Z�j���zF�/_!�`�XL�d ��:�w}�΢�+t(0�^g; �Ë��sxoG�p
9ll�O����o��\M�����5(�Fo�����4b�W6m�ğ+��}8v�c�89�*^�9x�4�	���Ҳ�U�X|/�DO�:�-L����NmJZ3Z���K�O�t��[��n�s�
���"��s�A�W���u�����p�6�(�i�k��/��,�*?3�`��Y�J���B�י��J����gl�>�nzmC�d땑�\�(�\0��m����+���d�[=P�2�p�ى�㦡�W/���EZ�����"��$���^N�a�`���mԾ#�~�|S��W�^��j��ˇ��9mf"t�S��f���̫	3ٵ��kx�b-�<��ue�)񎦯���;۰�k>Hڡ�Ό�M�q���>����԰�,���&s|e���u.כ�V݃$9܇��v޵��U*��Z&��t��ixf�-&f���YR�0v��'�U��sN��A�w�zE�PkQ�PY������8���9vƋ��mH�خ6�+�cEk�Y���N�l%���"�K2���/l�\�sb���GP�N�[�A�w��d��I`a��\���m)�wfօW�[���M��j ��U�le 'Y��86�8򯅳K	���ITd>^F�,p���Gٝ�j�pɽ�{��v۵5����WO;�R��*�>[�!@Զ�ګ�g/&�Y���|� x.�4��#�f�c�
�ǏV�)���L�h�+d�Fe�C6�C�'qED׳�p)���h��~}��0�`��Bγ�og����B��y�9�'����#`AV��su�rY�t_�g����k;4�q˧U*�~�UVC�q�k�/S~�Z"�`���tZ��9�N���=�ӽr��,qu����!�V��$`�>�C. ����nA�m ��݌�z���w�{�r��m`�Ez{�����]�Y��vj��Ü|��5t>�������z�F<�ϰn@���K7 ��P0��`-�{=�����s#Be����qGPU������xc��cw�s���A�E��fu��f�^�-�5�z�`�:,��t���"����Pb��0_�.�|�'�j7��]TeY��M��p���>�+��:�q�xX4��w��W9��$��cH���+�����b\�e�ز�A�6�[���]-ԼT���#1E�K7naD#Q>���&`_�ҙT./?�T�6�G�Ip���w�ξ9����<�����ww( wwӒf��U�T1[ʈN3N>7��oP�;m1F�:��Ldڽmn��=n����K�O��u������f�����)�QZ�����no���g&��Ԫ�nK�H�`�u��Ѭچ�+;`���9���63���:��Jm���>jwa���*��uս�g�t,E�k���-ꬬ��9�z���������9F�U�3y F?K���0��
�ج;q�w�`p�,�J�FxMN;yT�M.�tF�]	Sxwv'+
Q̛���1��/y͐�"Xc�� 0aQ��~g»����­�-6�5�:�s��B������(mUl_h��Ql�F����V]L��BĺN�QY�Z�|��,?R�v��ˇѕ����UV�k��ΌX�ib�xc���h��ǫg�˪��#�ɕ
@�-د5Ϟ?/��v/"�_��@!ӊ:㇞ڣ����	l�d�.�ٺ�P֚��m�U��b�g�g~�Ae퐣#kCA�tU�"���v��vN+�C��2=ۍ��n�q��dX�gO��7��f�U�I����1KIz)3^��<�.���JfX��#�����lF�7�vq���&,��T}�����N��%�[.�S�i^�ܞĪ|#��,�/_t\���.jș��!�c�aY8��3C��W�ʤ������j<'��_D�ۚ��b���Z�Ȃ�d�]?^�9r��l���Ce)+����5����*^���j|�t8t&������WFŃHc�Q���({�J�M�e�Kl��\4�`�]
�mP��t���:�����)�B�J�c�2��x ���=���S�^Šl�ȡӱ���'	��=�zYe��M�82��;<�����;^���T�uX`���u/�D�T�N��);�����%�泇&-fS�8��]�è�Be����W�~�c0]/(K�(+0�1�*�%��痼�{;c�NF��=�6Q;��l�D\P�$��&]mJ��d�:-�eC�7�5F2�G6�kW����@�:�-�)̖ AU_�0�d�PLjYE]i�>�+ʽ�(5�= �oQjwPΏhB�Ms��p](;��K�\LC+;�H�;�'o�ͤ���r�f��嵺��Օ(gx�y��A�剫§��K�u��ff�}�g=M����rÁI�P��	uI����:,`�V�uE⭧F:X�0,�Dd
��I�ҋ&ҵa����.z��q&z˙�.��0���p�7+/�|7"�S��'����yL��p������&+@��F\7�a�5&a���Y%ؤ3r��Õ�G����|�-�9����ۃ��ߘ��A^�
�X�!���=bλ�C�ve]y�>�p*�
��y�*l�ѕ't�]�k�oa��)r��mQ`�+|ֹ�W*Q�u˸�c�ه�˸q���0��4���}Z�<s^C�k�`"����>�;�۳7��L�j�{$`l8=�ߣDP}�}�zw����)D�ܫ�e*p�����{�q���>�e�=�2+��T�v!n[.����B��b��nb�3~k0)]�J��9=������qI`�'D8ɋS���0�qJ������ξ_N
�|٪�n�]�f[���J*B��6Y��	Y{ʳ�u�Q��Ob��^t� :\]���H��]�!��?j�#x�l�]��ӳβyy�[j���R"wH���#��b3zO6���C�]of4������p��ʴ��s�}7��϶�up�)�����;Y���Z��G��2�z[�oh[U8\*Zxf���Y�t�<�3]Ep�U�A]y!SMӶ��Y�q����m�a��w_2d��\ �_k����}��؀�=��pX qJ��5Ui�鋧�{��տkA�=DJ-�K�<�(o6���|E�I|^,k[=H<ێ�̿?o{T�s"��h�:^�#>ƃ��ٕa&{6��L���zs�Վ��Q�u�]f7�o��G�H',���� -�˽�3x-l��Y�{t��H&s��7���ꅭW�s"/�g!�DeLw\'�����S�0��Ƀ��W�o�e>������L��fI
+-�KXBoH�k/�\����ɭ�<s��	������f�(ĴiV{��Aߣ"t��h�v � ��[3�gk}(f��ޛ�te�㧣-aNus����鈹�����L��b���[�4����V̡f`d�b��d����/��3e��\�r�.�L`H�QT�F�@#V	��Օ�w��ã=�6����z�;�O����DG��U����_Ǽ�6٧�5r6���@�2:�eS���â�f�7v�t��䯡Pg=|=�t�)���TMg2� C;挍��M��8#���ܱ�=6���P	<Z:�~���������?VPϵ���ȹ,���X�����GvbuJ���ִ���. �����/��X#�B��9�lkw�:�M���k|�}�O�/v�(��wՆnVҳ�=�XrF�v�Y�!@>��nA��A��^�z�	s�+~��}��Mw;�D̗"��U,�0c�\���>a�Q���[:��J����"��tuIlȥ&7�N��ս�f��L�F�˛��J�������3�syS�1��^ۆױ�NR��u`Uρa�0����e��u��!�oR�V�/-%2�q޸ro�ܽ��=��[j�>��2;�7%�\�M^�Y��pf�7-�d�n]uI7��X �b�ʦg5����Nܫ�\�����-�*	�W�E�2ن���'-�͂��>l��r�`â��f��sM��ͽ�ˤ��F14�$`�i
����:'��bmX�ۅ�y��\t�����yd}6�Nw�T�L^�Q�ʆrH�g�lK���ӣ{P�"y�R�~�VacK�9�ӌ��;�ׇ*q
��]�rJ�0Z��P���v�����Zԙ�m������i�v's;�i
2䝂�[�yXXC�@�)�Z����ʗ���	�_-�#+�Sã����CVu����z%!b��Z���Y�S��i��o)��i�y����qR��:Z[���zr0�:0mD�iH\o9��w`0���|+����9�4��z�)h��g���ۮ�.��I:���X����E��Ih��_p;L{Nz�t��������M� Sø����]b���.I=�:��x�!<.םv�lZa�e�K;-MKk	�Bɜ�`u�n���U����7]�ȴ[WԶ�w��H�pR.]1�+^^�������V�]X�zI+;�u�,�� Z�ۻ�%֑a3�U�����}���)���S��JuT�q�@MU�|z�2�.bL�B�v�����]+;9bx�7V��NUF��ُ]��#E�C�0�`�*�5q��-�p�Õ��km����~N.篣�u�ݍ��ܶ�C$��z�@�lc3UtĦ�=�p Xt��YfAOf+�5$4e=�ȷMʺ����gkY�е͝Y��&u)y��Q|t�o���/TjP��-e'@,�+��t,�'�]1�.ҵ]���i���o���{��0�YЂ��$���Q�i�+.��8�j�p�p
Ų��3[�hR��n�״��+�l�C��ܮ�)�%��j�=���cv��Ψd��/��z�u����>M�a=��/��k�;)9y|��m����Vq��]���]��ś���0� n���wy��j�bВ��l�̓z%Ģ�5%��Q/�Cu.�Ϲ�س.Ym2E������J��ʠ'�BY��E4���[�ܾ(���g^Hޑ��l����n���2sh���x���%��n�����ni�(L�%f%yB
式%���tE�6d·iL"��&[�j�����ڭ�c��/NJ���6���G�O'c��#���%ˇ8;"*���0��q_m0@pQU6��a�hJ�r�Nܰ��AJ[�;h$ox�u�S�S��t!�X�->�fu�.ʁ��ը��Ѥz�C2ޡN��"�M��؃�1�&L�,���x��M�	٧�D]�`m���gi|���j�Ԯ��r��F��v�����З�;VL��g9����a�pM*9@���谤��oK�N�S&�&��a{�u�� ��LO�Z�
�u�qyJ��2э�ʃ,Fs�t���sq]b؎}Y3h����҂�ŭP)��u�b.�(�z-���lh̦q�7��6��	r�X!� ���έ���԰հ�q��gt��W���;�����r��|j�F�薍� Xt.�N^:�T��C~���z���lgZ�'c�>nV�ﱿh�ٕ��o�J%{�L��7`��Sf�����:l���Ȭy�8�^X��+w�q�y��KX�]|�W(=�Z��B�Is�|��L}s抳x~��!�{��A��ٲ�]�f���9ʔ5�9:Dfl�業�#��(��)NvR�)=��#}w�S,�����bG]Yՠ�v�J:5�M)5:5(�=B�]|�����v#�r	�<�f��Z�e��2u#Ճ���y�1j{MFa&�a豰���O
�T�f̭��J�o#��r����Gx�"�&Qԟw����9آDG����*��1k���C��J�7�G���\��ʀ�y�����>O���k��n��x���
 �HH�I"AH��P�*V��h��9q��h���1#���X��*��	����R�l�QE�EDR��U�f&5)eƊ""�W-��Tim�-�e-T�%�Arܴ����[��R�ڌ�F֗YsIp+��̡T�i�1WN� �*(���mXTB�*Q+�iE\��*��ҔR6�e�m�U��b�X���UP�2�AR��[QL���33I���)Kmk�S*�q�i+R�ITS)�+*�R�ʂ����Z0T1�[*Ѫ-j�B�ih��+\�1s*�Y�9­"R�VZT�DF*�l�+B�hV1V�"���im���Q��iQV�j�t��ճ�)Z���Qh(��UJұi�+�.e�V��UA��k��#F˘`�[YT��7�ZY�Ѻn*#+WM�*.4T�UU(��U1�����eSZ�`��P��D
"��O�G��H6/�U��r�h296d��nc0EيS�нY�:kyKZ8�����{@	ӷl���p�5��q%�V����c�J��;@���t�R�s��/�M��g��sU�+	^Le����P����jVbf�.J����N��~G�n��X�ǽ<gg+�Yޯ��m{�~�{�$m�W�y��׍����R��ؚ��[��d���y�Rb���O^����H��mC.���z�*OUJ��5�S\���t�z��n<,{J�p=wb�6f�aްaE�/"��	�M_T$����^�D��rw5l
ծ�vW�RWw��ٸ�V77�!j�ԑ��;!:�cz��FZ�L#$p�^�\j�ր���U'w\�k��	�A]�Y�P�*�:Pi0y&����{.��>�4�d�F��������E��7b�.�6�,�.������>(?�)�S_���5����2���ՠ.D8J�= �.6�����#��s�n�NdD�Y]R b�*1Q)��7ݰ��v_���w�g��+��U�f�e�8���o_�@�4�}�o���e�"�N���V��]&�a�2֛Vz����{%mf@1K�۫&�$���D��A�k�J�],P\z��{fo-u8��X���m����w~�b5}�D��yG��O�0����x{��\�ۤ��cO:��)wr�wR��P�;�����u�:�A��ԽC8UC��?(0\�5Zb��Y}���!�b$k0z�[$���%�
v�sc\s����pc;�,M�8�I�MVRԥr_^�r"�|���LWĘ� Ld�(�;H�p�7*���c0�:]�iʊ�:@/˖���Ů\�r��5ě�9bL��y]�+�(3q��T�=V�Y��=�>O8�����@x�Uci��}���kٖ�DkӦ,kF�y�gPr8��2Z�w����#���<�`�~XJ�C-1�y���|}��Z�����M�����g/}�W�lz�*d���4�T�UH}�A��Ic�QѕN��8rK��q��E���(4�wp��t��)T�a�C��2�&|%e�*Ϯ��uq��O����V3\��4�9��X� �ғ#T�/���g�,pt=�^u�ڪ^/�DO��R%��::����8Y�W�A���'V�\'�4��kT���n�#��**N�s��u7)�����9~��%x�+�S�ނ��W�:��X>p �>��L�x_����N&�]���O��׵��Jv�o-3m�����Eفe���@Es�W��ƤT*ُ�Z�L+46�r�B���Λ�:���jP�]�Ϣ�O���PX����H���]���ӽ�3�zS���ǈ�,�����U�3_��Oz�9���1~TT�2:���T!0ӳΜ?H�x?x�[��]�eo��4��ۆv�<�k`\־�N�����]��k(�����.4���}e���]HuԾ�K�<�(`���S������Y�V�G;4�[�sg�T���D��ſ
	�__�וq2�fԄ-���\�Y0� �9�Y�s˔���o"�}��\�BK�U�gPP�@�]�Kfm"Ϸ����nRܳ����QnCf�dZ�E�b�x9��������峾�.����Y������o}��r��	;;��5F�'�!�3~Q�P]Ehع��Ղ�Q���t�����l�H���94m��Uq`I���5��55��%xل�m	���C6�!f��]��<��@���Hh����V-�VE�KF1APΞ��5�^�3�wd��3�S(F{A���{r�*Dq.�e��ͬ�C,�0�en�c#gD?P�u����^s3��ʵ�*+�#{%�s�=Xiv��N����>&���Yq�\�9ٺ�
�N��nneF��Κ�����.��u�c=[C��sN]�Y�����viV�wl��|��ٯMMW̻M����0��+�iwQ�dF'{�X��*�QI$��4C�f����ٲ�#6Y8�:�v%����b��i[��ǲ��WE+��sqدT�@��Ά��ۋQc�m-���V����a@1�MȢL(X�3[�V�wrQ��!iUӸ[0^�}հ�wb{���=4��<�p�-��[WZ���{J�8�bZ�e`<���lƥ(t�c��-b[��dhL��рmV��@nMŽ��]<!XB��X����l�aθt�q�����<�[����G]�Z����
/P����OD��|��}�Q��^���u����U�Z��]�O�GP/{!�f��%��RK�m�ĺJ��3{P�"y�P��������z[��Gg_D�
�����u�&`\7Ne@R��clҹg�\ ���\gd����3=-��O����u����s�|���X ����^�5�(T;�҆��]�fy��.5��R���_8�`��
A�b���ڗ`p���#��f��y]�`o"�O{S�4���,�Z1rp� �Pn���Ӽq7�d35��f�@�w+zۢ�['�B���`9Ш6*��X��z[ԙ�ۖaEn��K�0toY��U�M��m'X��6d�R�����3p�E�%�Z9	0�rN�l�}2���M^�M�ʩٸ�Z4�`�0.���6C����\S$
�7#�b���W1Y���sp��&��i���^�^<�g�jK|~��ܡ!>;]�24lѴ�ٖ��R���*��0	Yt��Q#���=�s�j�������|�$�|����u}teu<0_J}:A��f\'S�~o	�Bɜ� i��b�p�*7����ev;�\NZ#�� �г�{��wd�%�Hr��[-W;;��$�-V.���Y�,.��٬g�b݆�d�n%;�ѝ} .��	��2��d��!��*3'a���!�Y>ޓa��A�Y�g*B�qaN��l�����Yc�T����1eqw�ꖰ��%s�7#�ލ�o+C��qx�I��q$����ͩ�ֆ�c�/|�R|�Pug!�?s[��R�.&a��&z�%VO`�Hi���:�,�sS�BYƇg�XRD^�V��M|/�o�.-��tVz��;|Õ��˖�N�\���v����rZ�4if�Uv�pd7�Y�ulvy�;^��YL7X`��Je���k^iV����E�N@�4���-�v-C�̯	�K ���g�EM���]��1m���*�u�4��7!��*M�����E�ur�s⾬���Q|���mXضҳB��Ėq5Y\����׸��Ї8f��=���{pd��Bd7� �(k�fuA���U6�R�v��2����ݽ�L�G;�dR��Ve�;(+�8��`���Ᲊ���ϯ���Z�N8��Və����/�A���x<Ͷ=^��@��Řn�Nd��,����E��S�R/�{��`S�~�1_��/�sW�\}�3b���+b��u�e85��N���{���$�K��6�V����Yӫt���#l;b�B2���hxF�P�zϛ]z�u��n�?Kd��H�J��S��Ti\�ಗ˱��T��B�=w}ʦ���]$7�O��ڸ�C�Ě���� �'�:r��E}�x��8a]Ojh����R�~;s�#�`m�A�KH�5��#�&_����!0�O��g6����T\H��y���Ӹ����g��<YX�(�gI�|�5(�2�Q����z�ut-�������.���~��^"��d�\�1��Á��X�\<�8f�4g�<����j��L�\�����%$�գ�(N�4��C�����7#5��S)h�T#�lgj�̆e�j�58�=��;��� �EW&�Ŏ։��G3x*0�Ϸ9VM�M�,�5�w�����u!]g��Fgv�l��E����5="�;����T;�ř���IT=�,i�`<�wU��p�m���V�2�=o�R��GIs���隷���攌�8E��
xxG]��:�[}[�:����|�K14=����ayc�jyf�˧|�M�oXjκ���q"'׻<'��6�dI*Ѩ�m[�ZcuY>�r*N�=�;ѧSR������1x��gv����S�^�-�n��y:�c3jE�Vf�TT�:������u i�����j
zSJ���%���e�W�
u��k��]��-�cXʒ��C��~x�ʗZ�Fr�,��8y!�R��|�,�S4/6٧+�����G:p��t�rǭSC���U�� ax�
	�|�ϐ�갓=�YI�o{�g����<�Wr\XJ��󊥟z�T�vZ����>�6�/uj���с�A���u��w��É�X9�{���l)�ι�[-UҊ
uF:u�]2�5}��ɮ�3���
.on�z�±����h�n�x^M���*������V�>W���U��[�z�:�i�\��{^���ٰ�x/� ��1�ޫ�&�R�&U��ND�cuX�f���G3q��Z�.c�!���t��sE>�%�9��`�ސ�yAT��\/_�=��"�5�(���r./Ϙ���Q���	�~���FrԤ>����|�^yJ�,	:��r2��LF:G�E��D�}tw5z��%��k�4�]L=��q:b��c���*��
���>hC��~G	�V�7��g��6�S<�R}f5�a�2��Q=�^���^-�U��fJTSθJI�t_H��.�"�s�D�gNL�7�M��oq�>ʤǅ�eUfu����p��{�����.�a�h,I5d��8��!0^�=ӭ�R`#�r���J+D\9#�nuV�����P9M�a�~�]5\�L�$�9҄#��sv��q���g����[�~�[��G-�����kմ'F7�t����n�>1^_qԮP1��06��L���s#A��ɮEoҙg(B��:A݈ b�ܕx~���χ�4�P��W��հ/���c@6�ս�oPW8*����{hnH�.���m��SS�t+�f���oګ���U�1[p��y�cNŦ4�Ҋ�1C�8���:0��G;�"�%�WD����0r!����d^%F�
ݺ�Ys���G�{��T�W>NIk"�[�n	(�#nq����;��5��V֙Z�`�:���.�u7��Y�mğ.��`\\-��f�Ó��F�o������J���Ĵ��\=�[B���CM���x�Eeu4s{:�-�ݴ�1�r�;}�2{�TI����
�X�u��G���頰ߴL�D��g Xz��6/���._<�|���P�ޥ�%�k���wR��J�CO1\��k��$5ԶLJ�3H�a��Z��6�}H�8Ϫ�\���L��B\� ���}�\����{=n��X#O����,1���n�,ܽ���[��R��R��yPo:�X�Lϱ��L`�����<�Zg{��<�k�9�@ȕկ��mі����=�I܉�AdŁtk��G�����cp66m��ã��p���j�ɾ���ƦW�,'[��0�ccϤ�VzZ�w��X���>��s�枯b� �^�o����6�R�k#�a�7����4�o��L����k��q-n��fX��ul��pZ�D^ҳ9��P
m;�B��z����yd�	աL��ŵյl�Z$�M�\Ϋ�ŋ�;'6A���|v�����Wz�@����e�Ղ���{���ޙ}�T�pe��������f�Ҧۋ�]:
yB�ؿ��ǱU��l<s���=���M�m��q�юz�T�T�_���1B'Z��L^r�UX�����G%󛻋�̤0������o��[<oL�o��u]tV�ξ��?���鰽�3&����k]�yU������0��)I�n+mUvM��1ǚg�mN�rK�{��t�̴��[�C8��7m
SкR�,�Q{khq+�w�c2<c�.L��Uz���n9j���l(ޔ�jM���
�Sƺ��`��ڄ���q:8��ӆ��nb2�M58J��ҍs=I�8��'ӫD3��^��o<�nV���9w�P�z��{<�{.YwHf�'��a/v	k�u=�׺^*��n`+��ƭ{=ܻNUbR������p���f)e�2��~���0�+ �e�I�j��:_K�@K�4
�e�T�r�I��Wa�Ж#x�̷�]��,Jf�Է����A�nN�.�b��3��t`��5�w��	.]x ���q�Ժ>��4�0{/����՜(ù�L�՗{:��g6��0�nhI�Ү빠t������)�f�OM�,Mm�o�H�ؤM)zw��Didfn��mH��ne�A��͚fV 7A�ب���J�<j�*�@�Q��t���#��nTɻ���":e�����9w�W=����ٵ�����[A���J�f��
�E���6\kM'יX�pA�%ۚ���
M�����e����TU��w�Mp7jf�&^Ρ6�����𕴒�]e!�˱u�p��V��|u�ؼ��I�s4���W��X�
�n�1���d�:��ku���=��\�Xq��ᷛu��L���Ю�SW�c6�D;}�m���h*2*�X�5��tn�ʱ�9j��P�U� �l�|��ݵs��i�FqQ��ʇ�wm��9�o`������2X��0'*Wr�}�M�^Z[��{x��U�㱋�r�V��Zf<��3C��YG6�ӭ�u�����ۭ�l�ܡ]C&$�K�M�|�B�[��	��K9�B�@;�Å#�t���ڻPKGu*�=D��E�քM-_vݞ�y^;�mU��K�8T�VWQ�1���,�Ӊs��>��Ύ`y"���|�<�HI�Y�va�o$��qWB�&��c���Tm}�e�����B}�����UK�^w=���,��-nBŦ�WW�Ŷ����h�q,���+�c-ǜ�x�,�|l�iM�N�F�sr"#��'"�w-T�Z�79�j+j����D��L���7w0�+���oݽ[Y[�U� ���.�$u��E+E\]W���wzn�x�T��f��57lh�%���"�7!a�U�g(�<o���ԓ��b��c+y���/+Um��/r�V� �r�Z�����(2U�g�p�7L��K�<%��]�pJ',L��$�3h,�DQ��=��m��6�f�uu!�P��[a��D$��j	��5$8f&I�*�t�eK����^p%P��M�+���x�+(fd�.Hy#:�);�f�6���ʬF�����>X����M�����0���E�uv�ۢۼN�N9��.�M��Ǚ�Y�7�)LG���d;	��2	�1e�[�-�|7s��Wb��@@{��vZ��U�;{�y�Y��8��ȻpC��م���b�fgM��c�**lZ�r�H)J'��dŔRΧ��#z��V�!G��]�F�պ���܎ɜ����&�Fn����}G����&��V'�d�Y��ܻ6���'(qҥfA��0ݡ�����<��;]5�x�o��49�h�Y�Va���؊ǂF*6������+��q��ڤ;��o���~IU+-�j���h��}�\��A��*-J+p̊,f1�-mJ��1�EKjV*´F�#X��[Z��"��m�iKU�����*T�j�1��Q�*�
"�*�Q���J�l*T�]a�ff1���*�#+Ej�e��
f���5h����h*�QQ*U��r�%L��P\u��"j��J�TTLkQ�+l�QF"��.5E
մ�̨�Q���)L��r��1���Yt�F�i[]k4�%�]SNLff\��p�b�Xʙi�5hU��Ֆ�
�4f1��̢"*��V�m�nV�Z(��iu�R�`V���W%�0b-�LDTs-ʦfCUDm+Z���h&Z+�c`�b�,Ze1+D���q1E���j"�*�
6�ڬj--)Q�+���r�J��d��$b8����pƍ(��l��c%[(-��NeIQkF�#DKkZ�eZQ��1TD[h�UQe���E�����TZ�X��	j[E*�c*,b(�(����
ĺr9aA*�ZڢTU[J6�[LL�Zj⸱UJ[Q�X�"#Z4*8�De�ī�&=={*]�7�)�õo-��g^񷕆��_+�WO�V�h��K*���h�w����ol��.�-&�}�b�	-�Wh�@����-�٥�o^���s�8��+��̩��iW��ۂ��3,�It� �����g��+r:_8w�T�<�
�5�yp3�����Ƿ%�Sfed=*�l��ե1�"90��5s_iF�c�/S	��7��N�I��7I�Hv`��8�g��+x^n��x���w|���������5z�;�Y��TSБ�Wm=ۆ�i���V�8kذSU���$�k�)���}�:�œV�6��{���\s8������n]�zT���to�gS��/o�uq���P�Н�7�{<��*�r�8|�s먔��;IΌǕ�O{֎G�3��HY�^��W_��gX�;-
SX�����f������N��i�حt
q�����1���A���+Xh�=�Bq��vuB�d��y�x�A�q��;3[��*��/k���b/-bKtr�]���y3t:z�e�h��P��>��W�K��jvd)�}g@�)�I�IN͚�6�����}z���Y�N�G`�VT���VoF�s��="탂�\m�;\o��ܮ�rt"�ٓG�ھ�%AXT��W�;zȼՏ9[�㔑i�Qv"�5��Q�y|�e�/��N&��ܾ�v�B�ۛ����ڀ)'Ro����o�TZ�-v�k�l+�<��J���%�ǭ��@N���e,�W|���r�-�U�ێ��g��>�����`l��z�m�i��-���mZ4'1�H�<r$�|�^gڑMMgu��>��_�t=1*��b�3�!�z��z����)�w�W#p��`&�7)e]�Y.�S�� �sqq� 6ឮH�y[דͺX�ĵ���������Q�M#^�}~9�d��P14���9,�
�Ǎ��s�L�|��>o��#&���c߼-+�5�f���f_o��9��g=�/k��(i�\���5}�N�]wR��)�Y˳��W�:>�j��&����Xw� �z$;��A��_z�^����T�=<N�|m�bI���懵U���2;���^5{t(���e �n��0���R�p�]�B� ����Ε�k Fh���/uQT2.���d(�eܽ:*	��,֙1�GXˇ�`P���%+/W��(���l�n��=�E�k�O�`�I��/]��v�X�mo��,��5�K��F�A�[�ײ�6��D��9�I�O�[u:u�<�K�����ߜ�Z15�����{:����P󲪨`f�D�I�/��[��e?m[B��i_T���5�ؕ�7o\c��ݞn�vQ����Z�N=Q�p�hP��l�hr�uľ���/�'�.�VwEZԋO7Իy�ٲN}�:�ORBŎ]�k�{]GZ�0�F��ܑ�̨j��,o{5]-N���گb+�k���gsSZ�(�8w{M1H���7g
m�ʵ�~�2�ku�Z�J�Ү6���&{$��fk]�2�]x� U�-w���V�G�0�bVk�ͽ{�?-�Vnt�5�D�_����:��yT�*��p�x����lf+>=u9l���E�U�IJ6��9�o��ֆ����~Ϋ�?f��)�uiU�:WV��J8�m�[��˧�f�4���*�u�h��b�]H/7y`_!�n�M�&������(iܮY�VQ]��t���-��cj�N�cs��[�&6�pi-��
��<�����!���r�i�F�.ʿ�q�fb�������8��6�7��#��8��`H�l��4Adtq�C�F�-�o����`e&�o-�`΁Yϼ�zC��CX2ڃ�q�a�ܚ��T�ig�{�NI���_�Ԣ��Y���aay�����ڸ[�4-�#���;�=1��G8����ypX�F3��n�}׵˽���/� (`]q!ف��߼������Qw�s߇:�re���|�(_+��R��M�Ken�g-�2�F����q����C9��Mu(�j_e;S��[8�\\cY�{�YW���q9������_CG[�z(?g��7:.���������13}�:K������D�1k��k7f�s�^!V��X��'��^��7��l���!`�TC�}�U���к}����Ř��yuӱ��n�=�x��t7���y��K�Ilz;��ZC���������B	3�e�A�WS��3|e�s���>��������o$(b���d53Z�/���eԌ���u�uq�,��.2_j��{�mi�Nȥ�	q}U���k8�E�W��޾n����)ӬoFj!MH�{G �l�ʾ
�����Σq����SY�D���tW\�O�.�m���u��UR�x?�����G�3'�n��A��Q�G���ǝ�U���)Ϳ��Q���_�RÝLѥ6��9���r�.�3N�a]{�3	-��v�D
}o��m�R����˳X�ė����]��F�IQY3E�;����2��l�V/���)�H 6'Y+���%�|�q\�-��P3���X��S�<���ؑWGV��.�Ԏ.���Yȫ�Q}e�9���&/S�zF��Fg!���I��*4�V�ך��Fn�^^]Y]�+�V}������..��b͝씻{MN�XK�{��f�Κ�,�Nl�S��~�o��<��DVmZ���0��c*Z~�*�C"�F�k�9����^w�f����}ڃ�s.�1A&����÷knoP<���Q��M�DQ=�����\��k��7!�ඛK6q6p�y�$`�wP��K�G���y�f\.�6���D��t�S]j���qɭ/S��s9��l��[v��aX�%���
��uܻOng>Y�tpg=�%[)����c/t³\�N㯱�i�^��d�5��5y]]�=��\�\t���֧V�.㝘��9���uSr��{�*���p\2�g���r|��e�V�E4��j�p��j&�oz�u�mT��[2o�����Q�����iz��X��r����q�]��jz-�ZfT_*�f�㷵[�EAǋO%7�e�򨕜��'������3֣Ez%�����{�-��cы�l������=�\��7��v6���h_3�F3���P�{
$�g�6p.+~޵��glR��sno����7#z
��k_#�4�[k.mM�Wv[�3tYa�)w��o[��C��k��2���4AY2�X�1wP�`���9LtB!����3I藔$���e��D/�k�R�W,�eә��ZA��%�)f�������*6��U�\ر��|�nU�@�^ �Ni��Y>C2�9�+i�bN���^��|��,��%\�ɥZ��T1��c�:�zs�e]�E��s;��sq���'T9�9[����Xi�����X1��ѵGY9�W�)n�=xL�3�V�7hjnw�,w`��y�a�G���ڱ�U�3a9�4��E���U�먃 ?B'�~��}*��[��Y�w[ӳW	FG��操��'Z��,]�E);��ٳ�ٍM�<Os<��7�p����S�j�B��о���	��x/�[p��[����6�;y�+3+��.{T�*Y�x�|��{���p��6o�DSm�/IO%�+p���y���s���uv?:�q�}8a�W�ed�w�p��a�n�zg��*ZJ3����ز9�'���3�OFh����|�R����6f@"8����u�aԨ�qI��q��:�OBHX��ϐ�t�tk�5kڐ�U���8m_����^Þ(EJ�M��S�$�6��V�4@�����Vw���m�	�� a���5�o�t:,EIz��0ʙ�@��\�E ���Z����^k��jN�a�Tf���բCݚ]��N�3�A���Lf��(���s�l7���f��Z���L6�zY��iLŪ�Z{V�s���k��PiX��6t�Q�n�j4i6L�:���e$m%�����u����E���/bY��yۉ�<n���;�7λN^����B�\�X��f�Tο6�������ۓ]�����t4��[X�S�)2�tq���L�WeX̄�ڏ�;���u�#:�f檎�����@���px/��6n�1���p�#:�����7�#[�u�ٻ-��j��眱�0�ʇ�j��^�&�ץ��ٹ����2{!�ժ�U(�]F85��,/5�ۇ�h,�W���9,ţ��R�U�6k9ejޯdc�4ʻ͗�fr�o����7�9�gg�¶��3yS�z�uX�qLJ9T��7K�[��j���U��CT���)9z���!q���r�Si��C%P��
�42��z����^HkT�M���Yٺo�ɻ�b/�	��Ȩ���vAg(:��n��t��,��h�8����p;���OT�����-e#d��j�ÕZ_4�q��U����Yw�{�nkw�V"O���6I[�i�k���d��L���5ma�q[j��эA�w�GA��o1�Bq��J������Q�������=��w�U�\d�/���{A��Q9{��w�<�)Vr�'�a���5�u�+Lw*�G�~�Kێ���Eyl��݁�ɌN�5Z�um�s]y$��W�ُ���緬S��ݒ�LO�O}�k˞u��}�wJ�ݝ�*��U�ES���b?r����uO���}p��9C�[zi��2���s��������6�]�7`>c��i�Y�,���V�vnQ�nH	�ހL��2�{6�]Wp�R<Н���ýaI�f�8��w�w����~W�pq�99�� δ1���^�.�R�_���*��*�Ɯ�^zy���l��0 �Y[P�+ �ǒ�!�Vz@el��#��Q�+p>�M=N�a�ʶ�������e���F�a��(l=�Q�~�E����f���}�TLl��:c6�@z�=�I3��m�ŖB\�*բ-}��N�=4�Y������]�p�x�*1@����=uS�.	$����N��*�e�Y
��sWiF�:���øwy�$ K���9����9f8|z�L���i�YV��=+h��[�=v��I�d�3G�poa�p��/���!d*cJ����{�qj8�['h���0;:�$����w��ې�g;-��,��K���:��jɜ����u��O�pX�����ꌞe>y�{���_"�\����8*]�i��hD�}T�nV�$;�S�Z�.;�P�[x����2]�1y�gx�K �x��[�V���������y�WҖ��n�cx��f�'$<���I�m\Lxro������Xs8��kQ&B�ݵ�N��ʩ�ݥz�f��EF���/k���=������	!I�2��$��	!IHIO�BH@�xB���$�	'�!$ I?�	!I�d$�	'�@�$�܄��$�	!IHIM�B����$�����$��$�	'��$ I?���$��$�	'�$�	'��PVI��Ezʓ��6` ������������UT���`0HU	��HP)R+Y�6�*���b�d��%*$U�R����5*H��cM�D m�dQ%a�M����W��mv:�&K!�m��k4�SeF
%�Zm�5����ej������)�͊��V�SlmV&ɥe����hҋ0�w�{�Q��[ ��4��kVIli,�b�Dڍm�*�afe�ō6a3fcY�e����l�[,�"�l�el�b�J-�mV��Il-M�mmv�N�-f���   -v�:��l�Ү(�C�u��������uXЭ�gA� 6V�j�M*i֥m���,�)6���r������YPP��e�T�kMkcKL34�]۞   ޗ������m�TL����C�V]f�
��e$���P�5��\��mkI٢N��[���5o(w���hP�B�
7<���Zͅ6e�����g   ����
(P�C�כ��СB�
�W�(Q��B�(�l��B�(P �ǽ�B�
(PQC����
�C�h;UZ�5��#W�
��)�Rvu֚mrn�mB�K��6�mV�f�5��F�4�   �Ų�*���-��MR3�v�����n;�+��R��T������Km�5D�Cl#�pR�n�:-mU�ӅMil�:�E��w��Z�ha���<   ��Kj$�i�[R����@˙3T֕AKU۝(�0��k�۶둶�V����UY֫���6����v�A����E��twuSJͰ�l��m��km�m���  �ԭ���8��5ch+���� ��bʶ�jU��뺠P�j:�ֆ�:]� 4msk�@PZ��QB�'\ �����6�֩�Rm�6�F�  &z�)�nQ@gm�
 *�AUt���T�ʘ�+UK�� (�YB�T�N*� ����2��ִ[h5���m�Ֆ�B�  ;�U�v[p
gn�C�v� ]�ӁJ���݊ Ul���(6:��,����5��ݻ���w3�l��6L�6��ֺ�  ��T����PWkm]�@��n]TP�]rp �]8PP)k	P��ҺAUC�q�(�v�[u�h5]�ww,�&fCM��Xjj��  �B�N��ݘ(�juk:R �5j����S;74i�
�V�BR����M6�i��W �R³j�`�V���Mj�;�Lh2��j4 2��R��   �O�B��1��)� ��@  T�M'�J�4  i"&ʥ)� ��a���W/�,�����
[���r��y�PV���JNW;N��yKP�f��Z�����B�{��D$�	&�! ����$�	'��IO�BH@�$��HH,*R�M����)0�3��x��%"4�
���9Yn�5.�DŃ	�#q_��c�,�^��ւ���! ���e��o�jYa%�#�i-�I)���Q�B���-���,�z���FL�����5&ts��5��T��E:,D���Z�F0#��M�c%Ռ�X�9�*�]4UZ9�6�Sh<+2�#�.,Cr�/^�;v�6V�CY�$�%�Y�|�]�X0����+��h"��W�k���B7�� �BAa�v������kMm`�sj���I��`r�]4���{[Heek�jVhO!M4kA���Qv�A�{��~�jxH�8�׃�B�!�S�BE��rؼg(�L3 <�0R���6�v�߶�*���
tF�.)�=�w��;��C�B�e+��V��R��6���c-�;U�띷@V�aʘ��A ��9��b�E��Fu�p�ȒT��A]e#֝U���.]c��@�`�S+d�f�Y=�J�>�r�z�5�b�v�i��K��f�Xf��'��P"�՗Xt�U�j��#53AXN�f�V^
!]`aLm0I
�:����N�Emm���MSͽ�g%��Q���U^�QG�(�빟H�ƫ]Gh�@����h��R��,�M���F��sU�r�h��R�16�_�@��-huyO!rQ�kN,"�S�/jP�*j��x�*(6�ŘP�B�E:��Wz��
y��գVi8íK]n���N#���r	����T1Kb<֤���Y��j�	h�H��© m<��+U[cX#N��<�L 	�^�#�_�^�j�Y�t�f�ޱ����$"F\A�V��,�%���M�Ho�j�J(c.��&��L%c�jŧ!b�ɚE-�nˉmGB��&�X�r1QA�H�"�ƺ�G�eF*8��ǵ��W�b��暛�݉N�
́3-*�I���,Z9Ǵc��rf�,�
�Ж��ҸU�Yc���V��=Jx�BLF���ݘa�ZS�r*���Rت�֎��JT�,Zj*�x���y-,(�X]	xF�V-���V�+N��9�	`p
�Y�;*:DY9�����	�~������xŊ$g���wT��S�p�4<�`@sX�uz���
�y��Uw4س�mG2	J��DLw����b�r�^aڍ��}�k�$.���:9�vp,TA����)^3Q�H�n�e<��jL��x%0t 6�˽#n�4Y�JأV�0�
�O����ʙ������mb`�6�c����b\�n�[�$�V���H;J:�p<PA=�ю�@��(�яZ�I�K�mYN�
d=i�蚒��4�V�[՛Y5kʘ�FjҔ��e�ݑ������ r�7,�+k&bT�h����@��M�hC���kf�2�n�95��Ot��twخ�XCp�f[X�i4(ӶN���*����P��m�
[Cul4#�d�pQ$��tP5X�I2�-Yv��1sT���}�f�nTwq�ӳn+�RJOf�ǋ��CfP�XLh"F��h�ƣ�/l�l!�#4�kM����I|_�G.�kE.�fƦn����V-A��z�&r��/v���P�,�Q��΂���#�D�X6����V�۠m]h�5n0�C�xT(S&�5�ZN\��AFe�Zh�T
.�Å6L%6�f�'[ǥIM�@�M���T�3%bkըK�:,5�u�Q�b�8�\�:b���Cj�
����ɺNe�okcm �@���6���^T�I��؍��X<�vp	�i��ZU��0Ѝ,�򅍡�])
w�a�1�W�(αm���Y軺�vn�槐Ñ<>pDF�ha:w.r̺%e=�V����˩��-�w+z�Z2�`�Hu���(Sw[�����n��wE�C,j�ԛ�#O�D3�df������b�N'6d����h*ԍ�Si[��<5f��)$j��W�W��u6�)\e�u,����7�"�'Tګ�G]a̔.��u�J��0<
bcr���w�A�ӏ �q>8%���Xc���|U)����E��,�k�[o)5�Z�+i"���j�Fjf��j���w�o���k�cE��Q��k]k����3{z,HU��gN��ÀfIMB�{�
d��`Y/w3pj;�
�`�}2P���e��)�%�mϋ��?���H�7!�4����lC+��qcr��r��Se����7jQ�[�-=E���x4NF^m!e%Z�x�̴��˥X�Ȯ��6��Td�0֨UDt-�xU�����p�zp�v��k�0�x�yyB yJ��w,]���j��#tw/u-��F�wH�+�[�[MĶ�WY������� ,�"�^Mˡz�|(C�LʁL�Sۧ��}R��-��-,�%�(�ڭV�Yx���U�d��
�R "��c�YB��	�S,�%:�j��DmH�򆫩VB�p�[H*չ���@���t����/(}(3D�m��{�l+�J��V��c��͆�xl�P-S!��຺P#t���1K�c���*�]I�)�v�B^�Tq(4�I1N�X����Y��7��doeܡPnVT�]?���Z1Xq�Ձ��v�ۖ�C��aV�Oqi�[�e���8��8�TF�5f�[J9�ג4��dM�>AO���N����(9�ު؉m��4�ێ�7JP�cw/4M1���B�b�Y�j�=&YI���Ք�q(!�P�T�\�V-�;pf���I���g%�\�*��p�]�h��ᒃ��Ur�0XFl%�2joc'P��a3���}y�̘9��\BI���1/,Y�A<��G�����mNCV�kZ�m̨)K�aV�l)�/w,�wPҬ��]S�R�E=cZ��́��2��V&�yQl�h(�0^,,4'�d��SV��x��/4��ǡ�Ôv���8����N5 $���X��Tʬ���Ȟ��A�ZAтhئ=�X`F&�G7JѦ1M#����T:7Tj!�Y���N�Y�b����׵��K�ĞZ�lD�[%�7R BP؆����QX���d��U�����&�e�ˢ�^����,�q�&|�ő�ȍ<��Af��;�KuJƑI^�v+�7{A�P$���RA;V�p:[����,�.�4�KWp�)��1Tx�� :��+2����`�aGe=�bӓjM�����PM�i!R�h�{���X�*�f�ZS9��^V:U�-"�K
Çn���(ܬa�	%x�V�͹tײ��n�R7xj��ѳ�h���0 ]$c�Ԁgn�2;ˊ�5'�$����=�~څ�w�nA���0�{������Ù���MaV�YF�s2=��(�*v-�	�;)n���>v)-�ܸZ�dVGJ֓w6X�,�ݣ��J�6M9�X�6�� ������]FY�n�Q���-�ӂ̩cbt�5[y���5r�n��V��e�S�!���Q9x�әW������0Q��y"o���mʻ�cմ��-l��{�5�����!il)�r�;b�Wki�,�PB٭qQ�.���X�;�:Y'S1b"�ka��@ML+��Sv�&ּ`E�"/9b�٭�h�x ql%�Y2`�W�L͂Bb��h2�0��P[[�����Yh)��ZG$�&�!���9E�ں�$M���n��f�m;��-�7qk�H��v�GhS��z	�+LSX[�y���D�Y�cr���%��X�s3hL�N�R�ۤ�T��a���Y��T�W�J���{���Ͱ�;d�f��oH7���%�7N�<��Pj�/s&kՄ�������!u�B�*i��+(���c�Y��V���ږwB��W�\B7�I�.��n3�i%�Uڨ��@Ԧ�`O>`�9���\�;P�ÊP3"�&�[��fQ���4Z3VV4�:n��[K)֩19��9Y�l�M���t�0���y[.Ʊv�=�OɫY��H�َ�n�ha��ї��0��ir�
e�)�i�{��J�%Xn�Ve<=v�ǵ��:N�T��N��IR��xf��6,ȶ�M�*	�Me�t����[�HZy,QJ\pbH�ӢF�e#�MY�a�A�[Zw���Y�rj
��C�;>%��M��9��wFma�i����Pב8i�v��%�{�K �r��C2�;ak�����m��д��ɨ*�5ˡ,�b�k�Ŏ�6$'�0W��B�[y��{��T�h��r��"��E���8/c�1��yxUiYX�+1�.8f㼼x�H�˺��4m�őh$��R�9�69aZ�r܇u���4�v� ���+����Ue�/ndB���s�-�5��:��V���n��3#m�2"A=�X�P+Vswa��c�z���ܸIJfK�����Ռ$╌&��� sI�`��]�g�kw����p(8A;e
�{wJZ�q�R@��X¦��%�"��IX�a�pI��V\7�y�I�b�t���ïH%X��Z��{{��sU�dIS�t��twgJZh�W��XL�L$�Kby$���[�@��$Y �G�R��ɇ&#Q��ؼ�[sv�4��HN)�l\�[Ca#�@�GT�ْQ�Fːpm�ٳp1����ҝ�p8��W�t�5�#�#ړSB���I2f*w�t���ۥ�����q�͂n�/�}�7U̱�)�In��7/XE�i�3*��T5)��n��K[�e���/4Ս�"�I�U��q�&�$Kc;t�Xh�Q^�l
��,S*�Lf�ة��� Ut�\�+pe��'YO1�lvk�Vk1%h��\ȎMYh)6Sa�25xF]dT^:��8|�˛B��v�{@V^�TK
�pTv�!��/��*^��ٸ �J�@&CqM�Á;�j�K��p�W٢���^Kvj���#R!G�����W�*P�Cx�U�n!���F�Tn��7,��ݷ��Z���X#/T+M���

����Â@����I��e���dzhķ�Iѥ����r�HVj�b�Z�F�؎D�d�퍻׃32�V�-��p�V��������Nҙ!����QW2��,,U�(A5��r��2CEU�!����9�b�*іc�J����G�k�5oFR
ɭ�f��Xa��m��̵Y	d+[W${-�sq	c7ي�V7UTj�˚n�ZwH�� ��B�����i����n��\Ǹ���w�5��J<� q�'�����LF�,�9xw��q��A�$���b�:����*4زi��U��IE�-a�v�v�``�V�*��ٙN��aR�O�����MͶ����b�ki����'L���R����A�S��6�`)"�AW����m=SD�L��.�n0r����?u��DvZ'�꽉 A"f�7T���Y���ǡ4kZ���AT���o	�ܻ�s��Z�L,ӋB�8����Se����B̺�]�n�T��J���]]ZEfԛFX�1`j�|�˃�;��hєY���R��SpmT����t�1Y�+m&	�b,G��)Qͦ��Ճ�l)G) ���79�9{YO�T5f[�J�R���b4/[�F���)l�F|λ1P�t?��Y��&6^�5���Y�*�]�M�p�r���X���uv(6��[Wh*�f�K�u=��
ҐN���aKu,�J�^Kݻ�$�(ь
���\�9� "&��Aym�9Y80/rlaVl��.�:�D-Ugn�i���꧊�jX����i�]�+@/Pe;jU��46)����fVֱЩ7)�+X��x���Y��h��e�&��a�YsI���e!��tI����>{f������'��ܤ~M�',�a��]���:�L#>8�����cf`����,3�%�ϗ�j&@TO��&�
mTi'fg��a���p$��(���$���ʕ���T�F����9PP5�pSR��B�Z[�3n�lf�G2��OVd���:�њ�1�[ḓwq�$���'Z�(��ut�l'2�K[��$s/��ۋu�!��Z�Z����	�SGآvE٘K)<b�Vlj�;N����$XVQ��u�j��m8���*г�/�lW�Eعi�	V��J��X�"EB���\n��AxtT�:y�zJ��vv\+4#�~��C
��T�փ>ȎV�=u�Ϸ�/b߄8��ḅ����[7lbא�a���vn��0q�cnQ(;�a퍕�ZC*�2�l�1&� V��Ab�`:ĝ�A�2�֊�P�,��i�!�������%[�t��ˢ6|�qa�R��-b[,�(��{L���Mw* �[�"+$DL
¡$8�+UfCZ Ұ�HWH�P�)���[�e�x##�Pjdc�c�hr8���j��
�
����t1�`c#݅�D�[Y�YI&L�v�C�=�i�wH����4n�*��-X
�āNb��yW�,�Ye�Ym�� K+i˸2�-��
j�M�{��,IPy�h-%�,���,{X�1j':6�2�.,��[6���ųV�M�H:�(K�6蛍��ݥ���:lL���$�a�5�2�Q�cb
u��u��a̅��A3��j�$if=��pP�4���/��Bh.�U�	9��2�,wރL#�.��;�#�������O��e��
�1qN�F6�۷3G]_=�*������v����fd26�����D�.����<SC�7ow��Ovl�F�9��(^]N�x�R 8����+�-|�!'�0�wd�=^�M�>ms��*l��t�Z�q,���$qS�����l5�V��=� Ee�ɉ��wMaμ��op��ظ�l_<�pdU!��CfR�9ż�5���:���v�!.�N��|BwF!�'[�-ai��Q�=p��6�ܑ��G��H� �˝�ɼ0��|f�o�ƣ�T���<�̤r�ƟZ��M���x�-c8���檽y��\�񨻕a�GJ�.:�ԏm�kg�˻Z:�$�1R���Qe��9:\\����R�	p�����[�m�'e������:��J���a���r�d��{S��<�ȧ�xT�{�����b=[3��1{<�4Ъ��Z�9[�p�Ic�_T�㽇rn�f�-�q�I�Ub��GN��-fܾ��,uB��k+H3��hT3N%6,��Z�����p�V��ʖ��6�>�l;�=ѻ��y�6��ʈp\��2@M^�p*9�!�����m�#�� ����o. ���L؊Տ��gj��@�ه����^��sb�]�K� ����Qד,t�=v�<8����>���h5�d_!L�n]��NP%f��w	�q-��K���M$��8�˽M��=Jߎrɀ�7"���$�YY��g2wv��U��|���.���k�;�&"�{�:3�m~�_A�Z�ُG��u���r"��97��zݷ�g�ΫS�����fnQ��>*r���
�D�<�M���	u�7bP�w���ɦb|D��x�dTY�.}ܽ�ʷ�0p���_�O\�1��ѮН�%�^5�*W}��̄�LW�&�����CB�sv��Ilۃ���)n:=/:�Γ��ָٱ�q�c��s�;%��\#��.�� ��%6ͰHec�v����MB�Lؕ�z�)[�i��f���,n�0�`z)L;�k���T��@m��������v�V��8�[�����Ok��KݞR��������F8ŗ�yt��O{Q��>��!X\�ƥ�5������I;"q�YN7}s)[������T]�*���EbҮp�ƜV�L �^3c���6*��g,D��&V��Lf�o�\����)ǥ���Vږl��y�}@�X�tIL�LC�؆�m��5�Wg����\���W��+O��<� ���������r�7Н{�p���0k]G�<_���n�����N��kX��Y�Ƣfs����i3^p�[APݭݻ�$�9��$��Ҧ����W�4>r�̽F�`[��ٻ'K2��ܮ�<��JU�p2I�fh�Sۣ5Z�J�L���ı�H	����ӭ��ܮ�wH�o�Vms��,$��ոH�������٪c�L��K��iS}%�s���sv� ��� ����]Ew"7���N d�&��ޱ�+٢`�}�����q2,��>�6��ʧp=Ú���II��A��"�e��f�DК���m�X���$�7N�Բ�Mh��7=���'�!��x�wb��;1���h�e-���ت=��c����F�M����v���r^c�<����������(N[�ܷ0�y���&�x3[ı����>�!�X������;�������D�����vΥ��
`�S�X�Yr��x�6�$�c�͆3!q����|:��(�KW@��i����BCO"[��kGoP��*�r*Q̎K�B%7b��xL~S++��ƞ���M�Uxَ�>���E�}���w�pW����Huyup 0t��TK$��o���yƃ/;3��ާ�K���#���K98�u��x������Ä���Z�+�dq��]	ݗ�Y��3�vx��]ͨ��mה�_�������ސ�e��3dq�mn_
�\j
>*\���d� ���h��!��3���Z.c�:�7����mm���N�x���ݢ�w�V��`9M�`ckE�R�R+���5�̘��o��-��u��١�Nc���S)�җ�.QsxvC��V�τ߉���K�D�ˬ/i��B�[�Iq��e�,ռ�OP���짖^�j/(��
f�Pm},�������6)=�zEc̢��JuX%�X��j"��-�:��ׁR�@���������54�٦3�沆<��Sq�:b�:����k��t���JZ��7k#�Z3s��Y�j8��z9й��a�Z�����~j�r�=2�+j�0/�ǢkeM�Z2����Χ�H���r�hd��3�[������.q��z�zo����(��xe1�P4�aލ��9�"����>,Q�=ZE��ekِ�x�! ����9=����	8%�����k�M�x���;O h-�F}�=�g�<��q��yɜ�Y�MP)S���A�˱�"��`�٬��Ɖ�ˆ�_^�.e�qԨ�b�3��ͺ9�~,�����{��e��<=�x�:6��EN���Υ]�4g'�b'W��Td+�q��W'����mH�U�f����jh|�6�X��E]��B���z<�`��oe	��&S\�؞���ݼ�9�tW��v,wR�tJ&��j�,g�v��+��*F��.��{1�eX��&��ݹ��6%w�w�v�$���W�-_��{�88���rh��u�����O0�+rWp�y/-�'1��SF9<�ĥ\�]����a�����ɸ��v��쁺Avn�28�;Y���a�h�X�TbOsm��1�)2�3�]-m�����Q[S�.��X�����+W�y.栮)���6i�i�wv���Z�L�f9ϲ鎾�90WLz�R�n�K�NÜ��zt���:���d�N=�õ3V��޾�M�C8���t�,��w5�2.(�7�U
���O�r�u��4÷��.X��� T�����	k�ؾ6w�{taa]�)n?�?
���r�?�-{�ڨ�J�ʽy��}v�J�/2�Y�Q��u)���4Y�t��9����d����=�p?��4uu� ��Ed���9�%�
6��-1��,���᫴� ��x:�+����@�*����{�[U=Q�n�P�Y��q�p���2�M;��ػ�::�i�{�g:�ae8,PS*�>,o\0��ޝy�2���O.b���%g)�J4�W���wZ�:���çK9Ƿ�^��M{n��ky��2]�2ua��ê��_w+ۇ��Pv���R�C+2������ƞW.�M�!\uvS�Fu9jۨ�G<�������e;�Q����]as���0]��`�G^<G����V�]k,�p.ԥL��u� �b#� ��7�%i� w|�ʭ�3ũ��7==0wZ�)gx�u��Twb�����b<uw<��J�j����W*_K�:�Qe����ۓr�\���_vv�p]6�����wS6���p>�s)���PP����-SS��8W9�4�E�]E1��Pr�(01��}ԫE[d�S��}����F��$Ċ���`�&=.½<�'1�����♵��7dL|9}��Ó��5j�f�2�L: ���d1\]�������`�\5�*.�Og�7�n������稃��m'�]P��n��z����ޗ�$7�+3To����)�4��Ń�o�|�p�>7;:yY���|g��]s��M��\�E	X�Yٕ
Ct�~����
��-���e�nTK|~�?>�fq]�v�v}3)��y,�b(�"������V</{'�$꾥�%��ǀ֜g��[�|0ϑ�7;�Cn�q����������j��P��`Ei�-��9F����c=��!��=ڭ6�C�0.��Qq�%�;�F𻓲�͍��e	�f�`u�Q�ee	7�h��=j��3Ҍ�t�nѵ39G|7��Z�~ۜ�?!�]0<�OA�y�P'�q�+F���םP��������}1ծ�F���J�A��S���1��(�mΛ㐷����vL���$�K����E�`��&�-Ƿ{i���@���g���k0�@�J��yW
�ty�R�h���%���e��1!��z1y\�t��R����AU�,Ε�j��b�3�+*���q.]AG-n��9Jѭm� ����M)�v[��~OG "�-��c��n�\�CV�lC!墰K]�����&�	R-a�gN�rK"ސ�խ�S����z0�A�,��Y=`h��}�S:~�x!�;��I>|5U��A~�B�P|��;.yw��Ɏ�O��]��1w�p�z���A�xy�0����1���ݙ�J�t̠�@Y��������^��aeN�4���9��f���RƒmV'�+���I���.�(�m��-���Ź�.�^��W�������d��3.6z��V��[�[�o��ܱq��͓��[LoJt���c��jT�N�½����et���(�RΞ�It�����˚�Ι���Z������2�Y\��zJ���@��VA�յ���rH�|e�a�&=��f׶�z��Aݼ����VGۈsB�A��Y<]��uf;��v���;sM�cDj��.��#ʝc�Gfu�:���n<0EM�N�®I%b�eW.hVⰳl[wh�إ�)N|.�]��gD�
��;Z$̖߰���Khu��ݪ���]�W��졧�`z�B�cbs�/����2\,��՛���V�<��]]���9J�]��p#9F���]ԏGb��\�M�{��zy���x�q�p]'�����0� ��+@A�8�`)����a�ٽ�z�kn��4��a���)0j�C¦ސ͐�ZD4+����y�����ݖ�]�Z��:9W}��:�z�MN�I4#���]���x��-�w"��'�ӂ"kX��7]�c{y�S׵�d:.�f���m��5$��/2�x���J۬iuCԗn]�fD�C���_4�}7����P�U�=�-$�.q���Ы�ǘ��������0�e�ui�͊+	 �^V�ת��
Z-��X����=�A컁r�ʻ�u�چ�Y�f	�`u�*�^��3�6S�J��hQY���Ϩ\:��j�T�"�j�Y�1v(S�[��_^��J���B�71$���W��ϗk��)0�h.F�P�!�t����>�p̡/mk�����/>���O;q3e<vwyۏ;�Ȭ��XZdI=��F�m���`@&�L���a� ����v�:N ��iw��䲻��=�^4{�c#B����u�M�B�h�q�8��c�W��MCU�A�oH.�]W!���y����=�pअHy�H�:IJ��f�o�N��¡���]a�f��7�:T�p9�-�|T#8���ux���C�[��>U���$�&���{�y�'��2��S2�E�v���Q���\�O/��=����.�ܭx !��Y#/O$��g��H���hv�t��r�R^RF��<��K/�{=��Ѷ��f7��z�3���q��wM�	�����v�<�]wh����50�!Y�N���d9{���2�ۅ$;I�fәbk5�WRC	o/��ur�ٖPx���8������	H�9�T�J������{��:���Y��,�Z6 Am�.������g��7@��tF-�����wn��Գ����퇨A���f�o;3W��r9�&t5jĺ���&��moQ��~���s�ޔυ�SB5���_����҃���%�ַ�HX�{N!�g��]Sv���h����5���,n�'���;������o�9b�E�N=�6��d:#�8�*�����ma��/���81�Cڟ�H���.sE	���{�2֗�����-r%W�`�[��NT�^�"Ѿ�5�E����2��p�E�9�Ǡ���g�_���V�]��lr����ح"r<%k�d��i�g/k������;fo���[�M D@$o��'v�X3�n'�S]�����SC+���	�1�T�˔{c��Z�9�U�ev�N�G����
-,�E��w�ܬ�]or�&Md�J��w�MR��t�M����wwq��E�Ul	�h+�lR��tn�~ػU���T��]�W{ي�F�	ǧ�n�\� �;[F�ɄB��D�������Z���&�F�]�U�1t�2l\�ι�ZG9Ѩ�;c��b�b] ���+fn�oI��Fj6�,����#8T�!�fnl��<o��YᗜG��x���]���.Jv�q�;����8�x����Wz��+e��LL��V�Oy�����Q���jqwٜ����X�q�f+B�Vt|-��eem*�a]5�w=ƛܴ�V ��4�m��R��ޥ@S��=\;�E7&m����\�FB�w����X+s�6y�7�N�Q�C�9vfʒ���b�Vڬ�p(��y�XF�|)��N�S�tM����h=�=�1�I�d��pp�j�#�U��6ZLv�=P�O��PU��}���i�"B�5�)����:o���8c}��ToAu��hC��mqӮj������0�u(W2r�+��z�A��eޙ+�����*���tFwɥ@�u�3�S��{�a\c��V��e�{���ɖY���T�uiMNb�'n�R���'-jBN����{��		�	!I���k5���寸�p���[��up�}89MEbȆ���..T��8��,�� ����OB��jt`���y{r��2\��+�'�6�If��X=��N/���l׸y��λ�%d���T��/ov5�����|)��_z3즿M��O43mI2ڻ
��fgӒX�3S��S�ɘp�R!<�v$H���u��G��$i���q=3E�lVTw��߸��G)�nW��J�P^�^n'�˧�Q��ެ�Ҳv_F6o��WΖK�\cv����o��a<�� [�S���aԩAS�ʖ��mĶ��F�K���f����!%8S��£�u��7��ԫ����7gy@�<~�7s6K!!@�vh{Yڻ���ʟwr�i[0�8<g��<��m���`Gxf$n����܇�@#�Y1	��t���D���.�vsi�xp�����$Pu�*�����ʈb���x��(��U�4�r'��˅	vY�]�sq��;���Ku�4���ZQ,/A�W�%�g�Nw��0��.ϓ}�i�/n�Z"�M8�y{�u�
҅�飵��M^T��,�f>����ޕ&�C-ؾ-�i�{��9>WO�m,#����]�
%5��/
�;��W¬�R�{�+��dy��C�j��D����V��:���_v�GcO9m��3ԉ��sCf�$�j���Ir��=��up�H�]t��1�n]����y �P�V��Q�֋1�6v ��Z�gh����S��(7C�H�]g�:o5�B�,�S|%ŷ�w��3���mbZ�Vq�M ���i��s7���*u�75k�z#����\E<�Y[�9+��P}����$�ۺ�Ƀ�8p�YCatSc���>PK+��񢡮�Yj�fҾJ�tT9��T����XMFj�³H�h������XF�%= �����,��L_u��C��X��Wǰ%i��}��^��7q��u7N�R���i�ZX�p��`{��/�\�7���Bg���:1W�t���М�гG���vfws�q܀����<�VF�^�<y{F�����gP҂��1�6�.�% �q�=�b�U���K����^9p7[/Z�U�����''	��ˍ�	��^g�b�9���X�	Ƹc��G��T��%%��v0���㻜��ܾ�)�@;��e�w�������v��K<���^,�aX�i�<�7�K)�sٹ��y��r�*��Ǚ��i�3����qM"�b�;ќ�lA��5�o�hՔ��)8kjwm�f���{'�!E���׉��;Y�����1�n�Sr2�7l52�=��:;]�j���4�L��O��Zk�M��(��%�)U�y���G�w_}dh��lMv��Q;�Z�a���MYq/�'~�D��r �r�1�ɛ�ޘ�v%�;䅗>ܜ��l��L�r����s��r���5�����=���{L:�z�ɬ":D�"��h�tɮ��0.M� gB���Q�ٰ�gț��\���w�)�Vr��j��(xe�5���C�J��F�˩<�����9�YI
�ӽ�A�.���r��yp3*���&c<[j��m�V_nr���.�Pl���������.ڍ��1���zE����]����ꛟh��n^ �9�/Wty�p��gB��Ue��&e���#_�q�9�]�M�����r�6�?�*K�l����r���C�Ȟd.��kh4��}�ꔴ��q��^�s󲅋���gb�|DR����_G�6�糅&�'�k��ݲhmt�Yr�7�\�)�5+@�j���Le��Dl켦j��Fw��n!��w^���;��ۮ����r�L.�hz���1ݻ�ܜK	-�ʊ���}��G���x'Of��L�k�b�T� �1K�atpe��~W��IMeL�4.�����r�lh�K�iLԁ��݁�m�=�_��:u��N�V`���^�(�x0���>'��Il�o��-��B�N��v�.>�M�yD�Mw�s`c��u(��&�t�Erɑ��t���Çʧ���t��z�2��?e���'A��}�c+O�(�1[�g�]D]=|��`��8��P��.�<�ZD�llg
���!6i�Z�v�<`� X��^���Z����\E��;�#Sg
5t�����[�+'S�:��X\*^fׇ!X��35U��Z�\��H�f�ñ'���W
����y�l[�z��p+�DG,�A���}�v;\n�DW<��-����/;m"���#a�p6z�璧�o�ൢ~��{ ,���&o
q�;1��9wA�F%̥���kY��3m'˽�����m-���Ա}��d9sr�j]�]{���t9�v����ڳ|y��ò�s��8���p�}�)!T��f�l �l�oA]���Tjk�"�Sk�f�E�5f+��i�ʷ�u(��ǌ:��� �Qu1"e���Hg7��ʻ��l='���᫐������x�Պ���@/��W���Z�r�<��o҄
<������Y�$!Pg�ۦjAtiǪZ��χem˹0=\��S��en.6�
\��r�kvg=��"0��ףq��z�C�m��e�0�f��V@v�.\R黝��E�����m�nB1�cUiv��C֋ Wq�zs�����A��IW	c��l�T�1�v�K2� 1�L��Bn�hR�'�4�v7sf��X ��Tj�3;8{m�8�fYe9�lH��X:���N�vñ�\�\�|7��I�3w�[�Vm<f,��Ի@�U#J"��a9{Y9���q'�a�9�E�qtF�����d�0n��{��Ε�q�r�,o�t^ȊTvìͱ\����d���0ef;�h)���x�gvy�h�sOS���~<��o/d��I�܋��Bvvt��V�v�/��A��.���u�+��K�rs�[O���������Ie]�9w�����"oQø���9�\^#3p����o6g�$`V/J79�Xk*kޜ�#���V��v�	}ʧ��f8
�[4ln6,;���ݳL�:�B;l�ХR�V��-\W�.�1%���nl�n<u��kR����ݺS+�I�^�#4P�f֘*}����h$�Vqӡ��L.	�����Y�IXm򖔿�#:��w:���w�ۉk���pm0��eG�ƻ�*�u�
\(�Y�p�QyX-��޽�:$9LQ��Kp�Yì�8bՑ���ڻ���<ٓ�Q�޵Nb��s�ohĜ��غ����1���ݜ�F�m;�d'D�]�m�u������[�������AS+`.ܗw�Wq��[[�9��=�|Z��9�Da^s~>kEq�g�I�.�ݬ*�V�_�_a���H��Q{t��O�.A�X�f�נG���T�v��*�xQWV{Y2�;���8J��z��:���;�4��$c���/�����Z^�I7��CN�گH�0U�M3
=}�Y�겶���5�^��+���,`���z�R!T�J*�-T�ۗ�%�wf���I��%.n�%��5ji�Β6fG�(A/����wV��z�����J�Ci®�����7�4�x0{���><:>�I���\��O��ZA�H=��Lb������W'����ċN<�oN����T�c�9��_����X�K]k�W��cwR²���<t� ﴼ�N�PsR WR�X���N7�1K�2`��:�DUд��zhd����zQ�Xd���F6�$=VIF9�o�#�Bx��`�[�&c�C��L��Gjލέ<N��l۫AVݫ����4�5)ݕD�䭖�n@�N;=a���eͬV`��@�9#�f�H]�+�*�\���$��UXwv����WLr�Cl�$�"���Є�W���Zn��[��oe/�J��.w"�S���l��R��]֍:�Zݾ8r��5��"4خ��ըx�Uu��ֲ��_�{�%��Ś�0��e�pr4�u�ޮnо�O��IXޡB�Ҩ*I_i(�:uF6�ܹ��ɺ�݇1Pj���]CfU+��"��C]`M�{ԡt0j{\h�w�}���ó�5tQ(c�m�ب��o+Օd�(���n�X�cK�pG���dN���zwt?}wD���"�U ]6h��Jy���dB�jtrM��U�t�e��Y;�V.1x�T�h�^i�j-�w�t�EwC�Y����j�.o��`��3[�;��{7��`�`����C�lH�v,T���gWY�Y���w����޻�3r1���� *>3�w�k���YJ>[X���������:=]Wd�hݯ�=�N���S�	(4�dY��Pw���U�x�iX��Z��������Y:<ߋ�[�����e�M�_�d;�s ���G�r�U*��8�%'c�ư�yW�����c⯬���Ќ�t=f�^+;&�>���Jǟ���OEB��&�{�#�}�˰��3���Zڝ]�(a�Y�H�u��5� �f�`����qp6�1G�=�����,Zs�([�<�A��fT�u� �)�zf�5\�b+��ёku�V��4SK/e������&S���y�2?M�!����y5�(�d�wA��o�����8�}s�)����10S�6{U%w#�}�MpV��*���a�n>�P�.���T,�l^��Yv�q��ܤ�t�w���3�����-h��/2=�G7�!?`3ܰ���0,��=},�)vL}���Q�"]/�C���z�/$���.@>����)����=�/���U�g����'�Thl��ͣ���[�ц��
� �%�/�G�������h��\=��8��<v��Wo:4�v��������F�Ȉ�R<"��)���	�F_,�ȃtVf�5R�
w,9	aZw�*;Y�0��̘��t�F,�'e�j-j���Ѩ��X9vb�q�+xU�.��1ZVo}���Ұ�����nd����x1�S�����޸m�H��y��U����2Dn���Io�,��*h0�ۓy��ή�Z���sJ�
m��9*����o>F�M�c�0��R3��'���Vu��Ź�;��P�p�6M��1e��T�<�E#����%�؅ѣ��+/w�%M�u0̑��*@����Ǜ�1�m
S�r�"��N��^d��!
�M�:m۴��j���݊�z0�e�	��Y+p����>�:�mc6oF#�+;�H� e^�F���Ŋ�J��l�/����\����N���透5����[r�㗼��.���i�����x��:u�M[� �s��dر� ^�\5�*X�-�d��C�,��kga��X��J��x�^�y�/��5&�j�a����C.Կ�^B�k;�լ�
(�`$k)���F���9����fϏ[r�s�i�it�ǝ$#&hʻ��n�C�L^]��<��vP�75&�q�E���U��Z��TU��v.�A[���z��`�cTT�0�7�*��4cD0
��s��f���S�<1G�j����P�����r���v_<0Y8��
.��mg�Hi�O"�p��U��_��/t�$.��Gw)Tz�����<\n-�T��p����f�{fP�1�����e������lDZ̄��U%3gfa,s֋��-\��)�l����WR���.6�У��_���g���ȯ��Xq!M9��F��7��}C�s�T���y0�dC���Z��k����������k�۩3GjR�+�����v�aB�9�����ݙ�8�����xr�MPo]������)�U����.n����9M��$2uoG]Og�w�o;;�JND��Y�vʶ��N=(%"A���U�؃o��h�#+¢�%�!\^�Y����I�>q�Z�tx�˺��?	*wӷEA�D�1Q/�lLj+m�mØ�Z�2�/��V�fJ	���w)�j�{P�$�V�`Liy�8�< �A@m����Yٰ:�{e�*{|ھij��cY��2m�&��b��p�[��p��e��"�i.Nj��/��3��ʥR��Ȳj8_J��][��Y4
�-��/&����U�"�l+�c�0(�:����z���P���h'��gֵ�h�(��S
�����Z�i�Y�����a$�r�V�I�}��j��h�v�签�+,���a��gaЂ:�QO��ueR�����Y����qa�)����kv�W�Nq�������k�9����MS���Yu��#��}��3=���ꁥv�,.���'e��K�zŗW��-e>SXV�hn�d�a�!��9w����o���Tţ�i(rk���mop������Emr�ZX����
�Z6����e��,��ɩu/��N�6V	�L.0:�*�{o����H�3��оK�g�����B	�q�x�޳֭-ͩb7� MK{EM.[t�cs�6�[���cz�a�5�)�uq���z�ŷ}����OD^�=�`E�H�-$u`�sF<��ěp>�NQ���s\��v��6�P�,�ؕnX���k;�^���Ml�k��8i�=���iD��p��&V�Ʈ�v�ҍ��Ք�6�v���y�f�,�(�7&f"'!(��2�4�1��.
� �tf�l*��lo���쎯5uk��2g�\�3�vƬ3������s4�tQ�Y�;#n�;��uK���[����&g[�>O�BH@�2^m�Jq������v��x�;`Q�U֣޷n��2�0e~�>���y�<vo��[�O0�����.�ڀ/$�L|5پ]���I���Gwp�A͒^��xމ{;�Ztp�B�֝L��v����(%|�TV`O4K*^����9����/]����C<�ȅ�L���1��q��V)W
ưF��n�@9����P��V�<��8�o'B��#�`gc�9�X>��nA9����	Ԗ<���%�]�k�����)�qS�[7\��=�3����ml#QU��y���Ci���q�Sy5�����Hp�'��Y���{�fbp�3{lޔ�@�i\[}|���"<�(�P��j���ɩs4�Q��lz+��fuD�Ӑ��C;��֐2�[{Y%keqg5BB�]]�̥�V��o�Ѓ���$�2�rm3�o��r=,�]�j�����Gժ���XB���粰=x�](�'9�lWHs�cvo9�CsU�z�6���K�����c��+S��f�(]����W)@P'	\\���-�[d�^v���yk��sg�rb��ݨ]�LSP�y{k�8�Pr�᝶B�^��gj�W�p�mI{�\�g+�{�/'���E�u�	���nj������u�v���7
L���.պo��v�3FJ��(��X̮�|��ֲ��f-��Ϸ�ٷ��d�mQ)J��B���R�Q��%J�(�1[e����YV#Jږ��Z���ETQ-(���ʕb�F��PeJ$Z�Q-�Tl�B��b�TD�*(�l�b��[j��EX�0YmjUE��QZUDZ��T�eUV(�Q�*1jDVT�UlU-�*�Dkb֊0e��ʬH��UEQDV��,��
0[j"�ւʈ�1R�UA`�b����R�QDb"(�	[UE���������++UQ�ֱUR�E���UX�R�����,-�j�b+jX��֡F
ň�DE�Ķ��m�ԫ0m���TZض�"�TQPDD�(�5���m�*UTU��V��eKm,E*��XUAb1QQZ�j���)Z�S,�r�kLʑ(�#n`�Q�(�TF9j,EX�J#iUb�-,�W-��ź?y￼Dy��1�yY8�� �3
����C�ډ��/zu<�BP�|H�5FN���س׉u63Z���y�3%�O5���8�ɠ��9�%p�A�M���>�Y�Ǉީ������eә��%���9�����證��+�Ц!�7�d+��p������g��E�U")E]U.��/w0�vB2�@�:u%�
P}�Tt��茛�dX鮳�o��'uL3gB��J�.̡i`���z5���P��<@�J$'����2,���b���5���L���s;
�8 ��C���?�:=��(�]�9Sh8�OTB����=2w@�U�F�q-�}�n6^�"����������Kw�;�#�Bsbj+"(�5n$@3��[&�j��~�{�Z.����ݤs�
�����Q|Y%�������Q~�Qs�M]�Rb.�]%�y��D��i�ү%����*���~���=�����*e�4�*�r��E0�@�ȱ�V�u$G�4+jp3[�
v�����sh!�7�tgT�Ǻ�G#�2��;�2����
Ͱ~��=`֍����K0�Z7C�6���nn>ֱ���e^M�｝K��c^ޑ�񾢓��E5���c��']��k��jN����u���=x�,{0'w9����e�	}�(��+�{����+��-�ϻJ��Y��q��mʎ����<�Cq��m��y���ʳ���K�^��T`�d�fӈw�w�����d�w��!�r:�F.����Ej������}���-��Y��2��9�
!hD5 ��ca�Y�_������ec�z���lHW��{���,z����?`O���!,��-"T{B�s�p*��=u50�v�F�/����IA��Ȩ86���+l��82�Z/�����3m=9h|_��XS¡�����k�:��[���!d�Q#�[[	H@S=#*ȃl�hP�W����m��-\X�����Y�G2-�)�G؏b�uN6�(|�[�%T�2w¤\Ex-�1�29���+�M#��#��ka���ڎL�(fj4ZF�V:�D� ��с��xlÛ7Vτ:����\�/[�t)`������#�}cY9Sb�)R���"�q�<��[7
�=�*��B>�ձv=\�h�p;gvC�CL�\��cvtE���D��P���7���ɮ���11U����P�V$�p��>�eŎ�U�̽5���}N�]h��H')id������;��^�"���?\;yd�ʇ�;�i�5�BŜ�:�WWXs��DN�h�m�r3���0��tY��OO9�n�OcG�C�����V�}��om��7ZqoN|(���z�t�Ս��3�%�YW0��U|��N��B;v�"���DEJ����]iaP��ʝ��ʵ�zV���^AB�M�)� ���o�S�����8@j�0T�����1[6�<g P�EC���Z��Vm^j�K�E=�Q�p��B�Q�Z�"�l���MT�1\�<�&{� mM�<�l�AU}��zë{��`SOl���b+$(`���+T)�A41D4}�Ɵ>1�PI��]���ݘ3���.MH�b��Z��PΎ#0���0�BaD3����qw�:��C�q4�$x�����unf�RK#kv.|�h�RF�{&��$[v_��}����������-w�&�g���,��M��q���5���x�v'x)����7���V=�a���k�3�xE�N~��#E��^N��};R��ok�O���DɱO�ƈ����C�GK��Nb���qݙ=�WP�����;p�2V��&c�+k����#�/��aEٕ���3�E���*巺w��;��T��Tclb.d7*�t�Լ���[B�1 'ϵE:�����xܿ��2��e�V�Sa;���pK�����G�jXX��{V�s���g9�r��m3���W�8��}��tcy�>�x�/�M�=Sk��A�O$� �z��GY�>���D��Z}�D3�/lhZ�`�tJJ�� ��z8]
Y��W����˭�s���CUd��'WR܊�]�R������c��t��٫���t��0
�u�ePՃ���X�>�5�w��v�zKY-��=��y ���>�*���S~��(譠,�7B�������ߏ��{E�������r.l��->>�H�}.�RU1���Z8�#&�ʃ�����=�1�>��&:q�;���D�VO=��j�Hw� ӫ:
^�R�>E�Z���ʔ��k�զ����s�vB���Ǧ<b*���$;���yӃ���qbh��.�H0�޺���f9��y+��W����Q�S��5$#x�&cf�sb)W��;�*��f)��]���0��4��ꛌ�f+�z�(!��P�����M��tl�?^�$��S�)S>� ���X��U�u��]�'���Q}4_�����v��i���I����f���aA�ܪ���d�����������l�^B7e��lduf�iw��ٻ:���OsX�g2�W����!���V���dPZ������^�I}�{S���K|�lKv�^���Ŭw=�/q�X6+q]���D^S�\VY+�ᷱ3ǣ1}/(��-�擡Z�86��sxi�\�)}�\����s7��>Z���"��L��kx�����]�U�
f�6���}��N�?�m���O���(مYm����`�ݝB7�":seTX
�<����+�H�#O#>>��ֹb$����j���=f��(7�>�0���E�	�pC�=�UP؞l��b�:7S��1���{�[�Vh9@��n<}2���:(jz
���Y�L��ȷ6qȤ:�c��5j���Wp���ã�ޢ���U'��G���V��2���=�J�\�_R�[{�\����r�sKV��{�y�,C�ODlJ���aA�=�bFƹuZ���F�)nJǹ��r���w ڥD�:�����g�.d�@���IM��!���Qt���Z�.GAV(l9V\v�oj��1�R�F��q:��.x�ķ��>��\�H��>"���D	�c2�[�,����q���:ʘ�h8�	U��;T#DQ�JN�r9k�6�m�Z^��n��[�����~���(?pV^̞��ڎ��B��1X�r�W}�+��^O�V{̄ևP-�#Y��=[�b-ɗ<j><��9����p��b
j���P��1��jԊ�zs)�6����L|.D��	���d��笚�s��q��;	��5��Z�<q���su�_r����4=HՋ ��r�j_��Ҝ��i��
��C�Uo0TA'�ۊv��\D��T7s7#�Å@kҞ�u��,O%��I���eA���t\Ty�	^-ʺE�mc]��)��f ��N���P�n��#�z��v������.2.�x̷9=��9�Cb&�{��]���#��a���8O���;'|�ô4R�K0�g5f�U&C�՝͈W��:n� ��16�C�+���и�{#&k�ñ-���^�"U��B"U�F ��7�zvc�f���p��tz��|���5�w*jF�*�cc��]���;r�Y9��]�����j�A�Y��α`���W���AK;�Z�v��)�8��j�楠�X���2��9����V⠅�*��{�1u�Ih�ipp��]Zzr��ť9˱��K�7��wT4��o��.��H쐔H��V��B
��]R�`:�zөV�P�&�\H��{�����d�}N�Nf8��U�uLb58֊]��s����\��#P��~��{��34���y�ߔ{Qؿp9I��X�}�0c����=B�"�V�=�ŎŊ�{�ӛH����~�h��1��y'DU>�Z��@q[������}$��{���]BK�����z�s*�c���H���;�� .���ܛ��α2�H���j�vNʣ�Р�s����;G`Bс���y��&s3���j��S�V�(����,��Tq��W�87>�����Brb�*Q1�U&����=*������<�=Vj�a!��׎qh�p�wd:��8+����`��E� �s.��t�j��
�����V=*�T4��A���G_)�2��
�b,�35�1"�ī9�n��F1�+�� Ex��P�E'f����}�h��o�v����
R�N��{�`�Vu1�T7��T������R@h2$��z)��rsC�w�W��s���fHc�����b��ֳXd���Q�>|*`�+�����v��MT^��u���հ�X��l�r`L!���r�B���A|>��c-�q�&y��W�'ˤBx�-MC���Z�vez�] a�P�C#����f�t"�E^��[qZ���I�^�މ��Q�x�k>գs�6/�7=�\'��U�]^.��08hH��e�đ���U�^b�9 o.�#�8����f����Y[6��D&Ccv�=����/��O��Ɯ�o�	,�Z�*����'w1�UӫP��#g:Xk�b��\介Qo'7�ɜ3���ۻ�FPŮ�uM�tU��p�^�ތ:�4���c��qO��:���l·��+�5w��|�!�z�e`~��B�J:,�.���O]���X�Yͬ0�XV�E�D���ʒ��ok�K�µ�:{d�SC)��B�aX�4��'���Ue>t�)^�GM��U�Sv�`d���1ѕ�~�D��S��z�EKJ[�0ÔoX���<�1���Tt�;H�5�2��L�> h9]�ev������5�w}]��� K�TU�e���N���ׂ�\s�2:(j������[�Q*�}�Wxz�A��3��e�$�*4*�X����Ѯ	UX8M�{���wO�f��^ս�΅�v�����ީ~I��>�{\`�"6Q�V�9J {*7��.��t݆c9ܷx??N�ѳ�|~��T���C����ྐྵԆ�T!�T3���V}�:e�u�pt��(��1e��T�r�F iՊ�R�B�P[�����)���ѕ.����lV
c('�'`�ߣ�	��"�x�
��� ��ˋ�+a�ڱ�[����h���)�廊/O3�ԏVWNE+�ԯzv�[ 8����{��F��yڑ�%�/*v��R�C�:P8;I��
�H�!p�9�SQjN���>W�;
���Vpm��Իuxn��%�,ϺwSgrG|��"��%��h�;�z�bx߳C�0���MBަ"��f6l9���)��ʉ.Q�ҸӡL-T��X�ӻ.��4f;1��d�#IrŁ�dpt1y}����0���(�Wl��ه.e�)��zU��P{(�7�����*6/v;=�cՒa9u9F'��	�Y���odhL�͏P���ʡ'\aaW��#�c/	�Ex�z/!�
�f

m��(��́p�v$ǫ7:`ܮ�zS0X�w����U�b1�
K�߽���+�Vע�a}���uc+��7��
�(Ъ�����ꕞ|TLX27#>:��9�&V�4�[{�v�`��x����s㊡K�k"ݧa���b�
�lOXn�MwG#9<�K�9E�'v��m_�i����fK5F�=6OOX��G�����_ e��Ӱ4��g�s���⊊�:O��|3Ζ��F�.��T����>x:��9����Ⱥ8f���{d�B;9�w_�X�>J�����ؘ�v��SB��h���+��p���a�T��鹚�J�ǔ���6��,}�)m�����-\�}Ck�y��Q��� �� ,� �������(�Y.�2�Iߘ�@�eNH�#w������=�ɐK��)�\6�`� ۾�۬�LyLBݻG���4-]s����f��6�H�79�P��a^�w ڥ ��#���_Qk���uW}����(��ٜ�[((|k�906)u�T��str�w�\�J$��T�+}��1��Üo����y��z��\
r|3)ż��OCr�ĲpE���ņ���4�{���E�����3@c�&L�haS|�L^]Y�d#�Jׁ���#��3�k�7(�ٞ��N��ȵ^��H� ��}mAw���T�Ҝ��r�b�!����ݙ�)�]N�^i���<�d��b'W ����ȷ�'�.�ȼvTE�[T�)f�I�K/���\Ds��u�m:o��RDp�U4Ԗk`Z�P�ȻU��)�����n^{�
}x_3=Z��%71~L���� <7�Po���#��l
�vA�/DR���,�bӷ ����P�3iD;��v�261�����:�9}&������ ,��ϯ>�U��4E�ܨU`��]�'�!D%A�
m���vv+��Z�V)kY���欻t���؜�s#�Z��e���;Q;;��qਲ਼EX��D��Ը��*c��RLI��N��p�7�=հ\lpŕfT���2<#�ś�0+�<�.H-Un��dI�-+����t��.���Y�}��e٠��2�9|y�1�$�;�U�X�Ͷ�e]-2�>ݏkvd�᫻��I[Ћ�Mv^��!�gin�Ȧ��m�A�mY2��{�B���<[N�lv�rfto�@�̒�m�qt���7�tz��ǂ\�M�ռ�ü�����n0����j]|)�1��j�rSes��'q���yI`�i�j�܄֜U���t�K(+tᨲ���}sL㼀���&q�9�z��d��Ւ�Q���K.oc�c�U�ˑqb�����y�/���wq�*ֶN�a̔nAL�`8nI���}*^r/2��L)��&#dWѝ��7��t*��kX���`U���ס�j�Wo�+$�U�q�۹FD���.��qh%@P��b_2��;���l�������G��Y�W�s*3���r�U��_ci	kp<VG���vxP]ws;y[e>k&t�wT)_T�V�>.����4Im�ݠ�b�3AK�!ݎ>��<�ɉb��?d��:s���=F�)
*��&s�f��4^Q���	1�+�@�%����'6҄w<1�b遜�-���˥��	p�E	�M�t�����M��2�o�ݚV8���E��o3h���W����҅ Aw24coO"���-%k���]�`} �ZL��|���ʖ�P�.5բ��s��ؼԷ�b�R��b��})��ܭ�q'Wo���3L��4�M���i��:A�+J��9�p��2E5%:��8!ʶ�X���͸�n��y��<����b�v���+��y�t���2�A'u��c���f�����.�b˭��p1�r/3`�&�ӝF7ܳ.�(on��8��%|
�̝���mk�l�fܷ�nmo*��`�F�GY���{�2�Bh��e�;hn_���﫼ϣ1<ٗ��}�S�׮И�"}�'w=`�+��&Jy�o����r9F�a�Gu��s4��LPw�ݺE��m*�M�� �U�>Ouw�Ƿt՜�8��U��h��z%t�9[<� ��:�
1vPO� �4���Sש<}t�Ȟ_;pVI����|8-�7Q���Y���9�M������龁^U��{%��;�ɏ�lm��C6e\��V�s���	�dR�̨�(Y��C��uH�-V�F"P�p����4�Τ�����⺲0�=�yVp�c���ވ�{�	K�tnlB�߰��E |u��	�w����(�5S>�sl��F^d��;�MIS���c�SF-a�ñyú� !\�q�T�/v�S�@2���Gz�E�2k��3߼��UTU��*�[��1�*���U�b*�ص�Bۖ�1U��1*�*,Q[B�m%0��2�Z������b1X��q�cE`�µ�q�" ���2т�(�H�qZ���QTQ����Qh�Kj�iX�5�m��[J*)��
�墰W*�Tna���������+�jUTZŤ�W-aF�cQAUV+���mcmR��J#m�E�Qj�f5�*V��X��QcXQ��������r�b�EZ�F�)hVR�QX�q���(Ĉ֍�T��Ze�YR�"�DQ�ʕ��mb�(�*�cTQ�b˙�[��j�e�J±��kF*���EX�9���V"�h��QWbT�UL�����cr��̖2�ƥQV	lZ1`�!Q���m*
e��+�J�`��DX�*QTq�QP\�{�W>�ߵ���y~�:�F�}�@Bט���ɗ�5;��~���9�|[�!�Z�����:�1G&�&1f	��K�k���"_�-X����)���U,�(j�����gX�s�z:�*����*���̅\O�@f^�c���x�R�S�=~	�EA>#�R�=~�����Z\?p�+N9tM�#7\��ģ���	�о91S���m���4:d��=��� )����Ym���]I	�t�1��R'hp�֫��뮎��c���R��ԋ��+�`PM����Q#`�݇L��%�%	F,[�b�9�c&�C��Cj���G&z�C��6��U��8���h�G)�t���'�=Y��@�	�6lS�L:�l�:�������}��X�NQ��XTa@R�u8�.�{�΋/-�Q
Hj���N,9�#��i��ݐ�d�7}����v��ur�z�n��m!ݴ2$�q1H�P�w \�( ���m\����z���2������խx����8�
�j8"��;SuOʀ
�P�Rvk���{��eqx�t	w׻6�t���B�Ij�)���UȀ����T�
�d]�`�z"vK�3���9{6�=yQ�q��T[~�j/ W�W�6�u���˛�Т����zn�i�^�]M��R!l�7<�B�l�K�G�u�q^l*�hj�ǫ�vs;��/�N޲\|�Yd��M>[��8뒞�{ .�xL��	�;�0F�}�|��/ا�tKC�4=4��9
��@{���*���5R�
�'��s�uBiO�6n�ݗ9\V�6+���\8*�����V�5p�y�Ɗj�]:!v���g����H�'f��m�g-5��o�v�z8�0���0�(A�
!�W�qe<���f�� ���s����l��R����zh� �
����4��!�ޯ`X﫲@��۵�GӜ����fW�G��)4�ث~wYx+5޽,ϼ�1n7���VVS�`v���hJV!�I*;��;R�,��犮��N:�7[˸�R��I���d;K����\.sT���y���ҶN�K�BG{Uy�ݸX�[/&c�+j�R�!�>��B��!��CR�~�c����ܠt�׫f�9�05Q��Ndpn�s~T�����Y��ҷ���j��}��AOI�t�8*\X _�}g���%N�C���ɝ��ʜ�J.Du(X��Lu��#�w"�K�ZQC$ MpHj��_���t�Fk0�esn���d����5u���z!R}zw;rp7ֲT�z�q��@�D���n��F�e�����vZ�Ut��,�F�$��g�_PSТ�=vt�L�5H\��`���0��p8mv�6�ᨩ�z��s]O���ѓ���]i��_}U;ɩ��y4����+p��ދ�D=�.(�`��M(��T�qˋ8"y�wԅ=y����ӹ�F�_��d`�j�M�����Ш��%B��Q�~����#$�{ļ��;d��!�v:�	M�w�t`g1��4�S���4��n<�M �!:�6�^v-�ٳt)���R��L6G���X� 31�PΜ*-6Th�uh�����֋�l_�42��1<��4t���މ�@�w�P���
�6���~έ�������p�CZweo�dnb#"ٯW��W�K�/��u�/�ܾ��v(�?g"�@o�s�aNWt�.�� ��R�_����uvTl^�v��#��LN�A+/�Lp�kka�	S�"�j3�P��qt79|�\��t��*~����^x�et�|��j͞B-��T���M�گc�#�4f������W����\�3�j��qݩi���g��{���ר��?D9��bEPy;G�V>*$��#ϣ.���q	L!�Oo�	��d�@�7�R�����eVnˢo��K�-c��Mnva��S�r�G�н֌>�f��rM��X�sC��+1j��X.�����jA%׭��m��v��h��1�:��k��ݓxآ���A�9�[�詐���U{���p�gM5�>��F�Z�lu|@�P���E�NÂ�F)Ъ����R�j�,�/�=�[�y�*�\�m�������S>�>�z%azv}���q�ʞB-����;�Ot���ͺ�#�]�I�W�0����\!\�vL� P=]~(�#%�]~�7�n������<���}����u�]
����G�6+�;D�FĨ�s������Sm�̈�z5�H�$dk�~[G-�d3#mR�"
t�^���Tt�WDd�j�F�P��Ӗ��-��E��xk!��r6
�Ca�+���{T,�=*TH��һ]�6��uٜͨxyi�J���..�ׄ���=��<����<D :IP1m��$�n�aɔ��1���d���¦��s�Ϋ+pvB>��x���>��K[�TOs�w[�{<!�wEdE�n$A�<5l��5ߗ�SgJr�zx@�gB��W�O�5'ė�xF����7�C��@
�@M7^�u����]��`c�����M�I)����^�'a庻VC�g���L�ˊ�؜���tqU�5�5���溅�K��m���v���_v��%!R����Sָ�"{�d#]��eB���u6G���1�2YɗPQ�s##@g�)��OC8gn�-���e��Ϫ��Z��S4w��_���#�!��`ߒ,t�q@ԑ#�^h�,��� ���z������SO7�������Pv�9�� -��xo&�ߚ92y�P��������Gw�c�;��1R��Ӑ}f��FK� �҈v�C��:���ګ	N���������ޱ�(���1��0�v�د@k.��P���Cč��D5 �X�l,�'6���N���C.urv����`r�EyY�������{u�2��Ƕ0���SY�nj��~ߐL��~�\i��L���}�h����B�\��Ga�GTKE�˪Qq����ŝ<��֮P��G<{��&�܎����������vHV��L�?W=��
�KEД�X��I����I)im��(tu�my����:ħ3}��*��mH��t
��b�B��W��]�o�Y����R��גg��<y�Y�5�Sjǽs�Ug;'a�w5ZF�V:�7�0 ��xʜ\��v��i��:�q�t�
�%��������y�����n�a�5X�43�R��A�+��|Z%hP��3��#*#�%
#���`�;F{���z�,�0)��s��
�c��.�{B�-�]�>�����֩���G:*ȝ���A��:�v�snG+��?^D �!����a�16�]MlJ�<�.ykHik0�E��Q+��nH���ܥ��Ѵ����2�`BV�2��T\���)����U~�v��J�B�*^���@��¢���?	�u����3�f���z��2zw��3�,4��Tӑ�B5�Rvk��¡��Ƀ�����{���[�Kd����)�q9Ȁ��S6U1���Ȼ�0z�LV͹�Z;���wx�K;�5@~��P}� d�';sP��D5��V�D�K�3�L���8��bdE�����״�>){N
�e�W*%91~��"�Hp��9
��S����V^ӡ��\���Ꞁ���{��ڌt�x�:�=�^��@Ì�(�}����c��0���Kxїw�䗶}ƦO��_��~~�M�^٘ll���̔��4�������ۣ֞��r��P��U���\>�K�Gbw��ey�b���t��ޮc�:GU�u=�ͩ��vUDf��V�R�sf<=Wx�ZV?yBt~"��tnٟ/k�(N+�`6^`�g���*�)fP�wT��xh��̨�
=y������W&c���z$�qs]7D��vN�=B�pB��y�����]v��ΐ<f�=cip���N��:ޭ�R�.��7d:�eLJ=�*�f�KI}J�'`���� ���^�&K���
���5�{1�ݴ���U�.��^zf:2��r�@x�B��=q;|�ۗ���\wGZ���k��7���s
[�ٵ �x����Qnq�;R����I�h��Jn�Dٍ#�R8\�(#E����fJ�Y�GE{Ud����Q8Sѯ��]}ɪS�۹�T�����N�!E�����HQ[Us]���|'b��g�3֘�ݼ�,T����\�T�;�w�7��>��������e
�-p��a��x,�1�;
]��<��X��Jr4�?\�9x}������Ѝ)�!8>�hTl�s�������j���$���v���=�H�F]���2܇���4�
�Y��{�:��&ow�j�G.o�����3E!Yʗ�*~.��>0|G����ٯ����5��^k���/�
Ƿ��w=Z�K�k42�6�ƽ�f�+��|�nlh�� cx��L���AuRx�kݣ�f]�>��K6���#��	�;��Ʋ4�1Xؿc��9Aȧ,/��_��=�u�3�f���RѿCӆ���F�M�bw�a=��lH�0I�֓�u�u�x֛�����Ŭv�(z�e��VI����a<g�ó@�%aR��,�Qpf�R�a��R��{���s���m���z|1�fz�*�gd�9����ռ�QL�[{1�6U{໌lѶ�d�
p"*)譩!��]���v~C�57՘�d�\��:6r�^�(�&49�հ��ف�W5�s$k�#mW��{������N��wt��*��hB�K��a�k�m�k��oH�|����:�
f�5V��N����J��c{��-N9�&âq��ô\?dר�1c)D9ޖ *Uм������=R�R����d:��ɹgU��7�����c��s��m�8VS�����/��nӰ��Xz1M����T�<�ԥg:�Q:�+Q'�P��e~�q�&z,p:(豲zz��W�sW, �.8֮A&���ū�"�oʸ�R���)�
\:�zj;&R�(��?v�4�$Kb'�����rѩ3����ۢ�ؘ!*W4�WD��+͉�u�K�sz�Y�C����y���#��P���Jz�lk�`]lo-���E�P$Br�[���"��i=Q���p�٧L�O:��*�h��*��X�.;[7�C!�G��(�b^���E�@�̣�o���RP���5";�Y/A�Ub��^�~Ȗ�m:��(z_T;�Х�=鼽����S[B�1�u���Y��Gι��kW�l"dŠlRX*=�Jm��;�|��Ҝ�`�TVu���;���^Q�[�r��oE��Ht�w��{��w�Q���̱�?Lb�蔈�n/���3� R�w.�>������'c{�1�&�C�}��W���#��X�Q��]�&g�*o:Nc���b�>��	���b�S#� ��N���әB ޒ!��Ȋ-[�06d��Y�j����rY�֨ӧ'Ƕ��.�I^-10?eS[������\D�j�d�!�5�q�h�cj�[��'=�3�&'-f����V��G�LC��N���6���G�4+js����zFԙLZ'm�wz�(�c/���\�{h�|6鹋L����!Ἒ�a��$s��յ�v�-ٛ��znЂ��K�i�H�/�6"=B���x�J�,zw��/�j�'us��j��n�
wE��4�+�A_�o1�T���6+�5�|:��|��y]wݵ��~�Z)
D�6�)���|5b7gb���R�;س��x=�O|���c8�Si+��� ��
���λH?P��,�c&��P��ٔVm��*��?z�G�G�x\��u
�AM����b�����X��9�m!��i
��<�mE��Xi>���9��i��_h�~5t��Rw/�`c8�P���|�~�n��"Ǫ����VH2q5�@��ȳ��$���Rb�j������k�m�N��C�ێ������A�9�N��svV�[�;gw	L�s�R֪�_v��fG|D��s�]�1���SޫD��I�x��K��j,Z�u�[E^m#=�o����.os}T���!�O>�I6��u<2��+��S�P�� ��û���O�Qd��dS�O\`�C�f�A�����{���>�sy�8�*��ѦNX(
����K�f�~�h����{��d�-���rM��
�g�`:�d�l�O?] (�Y>q��|�O��9��HV&��M�2z�ՁܸβW�Me��`
|�F���$O���Η���̧�U'�ގ���*C}�{�����c<5a��<jVo�'P������b,�
遬��J�;�&�P��������>e��&�XB���`q���&�� ����ef���n�ڧw7����G���UT�� h���,��A�����~La�9�Af�n^a�>B�����m�Y�~N����ɟ���6�|7Cim'Ss��l����V-�|�m)_3�{�� T�����l.����i�T1���]����%M��

/�N&�Ri%Cyd���B��e�O��R
x~�OΒu*,7���'�/R~͕�M����@:r�k����߅@���6��׺�>��!�g{a��=T�'ǽ�H�zʘ�3�T�B�c-��,�a�;�X�{l�<2����2d߹��I�*y퓮�O	�6�廊��Ņ�%%��<6{�����1����7���a? Q5�`uY���̇wa�P<;�;��YY�3]�1jW�9�§�:�$�C5a�E�C�]$-��z`�j���v]3��N,����  <��ӷ��o��i��<ϲ���
³L���v����4�}̛UH)�,��6�CӼ��
���&3}�I��<O5܊m���s_��u(Z��G>gp��`(�Q��*4��Y+w�0��5i6_�+7�& .�n0�
��?Xz��m����M0�*f�~��-`Vi&���

/�
��@ĚCYa������>�a��8�P�|VE/�Ɲ�DyT�	�'N����>�C�ֵ>I�?%E��Sl�8���g���7��w��ݫ&%g%g�*,�eN���P�O��N�:����L*��~-n��0f)S��hL�W^
�ۋ)��za�� ����{۳KU��r�N�9����7��ٺ{�k7JB`��bng�J��r���	�V�ѐK0{�w�;K��Ƃʮ�QM���)�(��/�B����@A�_g��a��!�N�Vl�W��6���.���p��cY݆���t�Bܷў��yk���٧����i��9<ՠ��E�F��^VL�oNF��fҔ�QW�=�&*��9Wo,���7�J��T3D���4��38�v���B�Ú�r�pқ�d��G]�`kk(���W@��RjN�3@��FVG�u�fp�{�:����)�;��ڰ��h'r��ğY�%�糋̹��leڕ���{�0����_2���>����[��*ɣ8�n$�7�RWY���Y��r���.�tӝ�z:�J���w΢�}or��f�\c�R��N7��	W:�k��t�r��V瞑���el�3J^\ծn�&�XPAu�qV�C��	a=�$�c��{)��&=�3鹇aȜ�L�����Δ��j�������3�EU��J��S�����a��՗���V�ñTi%�����^`NH����q��ީ4��]�!���o����mD�2����,�b(4�˴�cqN�%�^����yے����g��\%�z!�a�������ͥ���м�nZ@#��zq�p2	�[��˳��>n�Vh�0��^L��<:�6xp��91z��V�9%��U �C7�����}�t��+��-g��͎9M�_*	�lL]�5��`*��d��P��4ĝ�D���%^!r^���C$߽NΆQ�ao�· d{�o@}P��5�c.;O�K�Yp!`L}�U�x>)b^ͻi�4��Y}������R���������֟;�sg�b��t
X��%������7�#ST�x� PnK\��򅭠Gv6�u&Z!���_9\kqR���Y��NԊ�kü��ݧ��u�觽�4�;� �X�/�H���;]7��_���wļ��g��Kp@@���ƥ+��b��Ǜ�`��T�s�;�(m;�=N�=�a�ꗾ��zڦ�	}���vO�;emm��=��H��(b�7��3��U,,&.C���0^�/v>��t�(G�2}VJ�:�*6����e�}������},�K���˿�­=O_&�K1IWo�]s������hCp�8�������W
��[FoB�d�U[ܸ7l�q_9�$��L�=�X"���<��}�xZ@��p�C��{���,��î��A�t�X*!w���u+�q�)|��>9����<7��E�vFT)�������|p�g�&�Ȑ�<�w9��㬫Ix	)7�$u��2�r��ӻU�s &�	���/�O�*ƛc1vW�H�LuY�;w{\���v1y����U��mf�K�TF?������6(+(�dX,F
�lm
���ZTb"��Llb��EPQĪ�3*(��DE�
�����������nZ,QQE�UQDF�S)X��ۅ�b
�a��`���D*V	YQ*��##�D���12¢���UUX�X�,����b��)Q��X��AH���TX̰��r��b���TLs(ő�D����.2�ffb�����QfR�QƊ�Z�e�b#�+*�1�%B��cEn&
�9i�,Q��%�����+���aZ�b�eE�SAE�VV��`�5�AX��"��"��drъ,")����*
����-jX��Y�3,�e�UTq�T�*�DUAEDX(�m++%Y\qTTQD��"V��DJҶ�����*�ŋ�EeK-��3䵭C-���)��b[Kr⠨2�UY��c*"bT��\eEX1UUWYl+Z���6���UX�X�9�g�}�E#]�P�K�$�$.�j�����w��]�r�h�VG�/Y�	mt�Ɍ�L���g�$a�뉽�p��^���M�dk��gr��� �He�O������V��Wi�'�;����9�B����|�o̞�ua�vϙ+�&��B�S���	�eH>��'ua�B��hn�k-��론S��ru�S����3����X5��l��?!�~�a,?0�Y�g}��C�Cnw����������)4��!�S�4ϙ<�2O��4��
Ͳny���8�S���V xD�NRΤo.q�.ߥQ�J�@p�q��3�B��Y���2�Y����O��E'�ϰ4�0��CI�zsx)�%b��)�H{h{��P�<�dĞwxiaS��<��O�	��	r>p��ԥ�l:ھ��uv�x¡��0�n�g�y�i���&��)������
�˞��'�~����L�N8�IQ�CI�&8����*A��g7���l�Tx���]\%���[W�nn���R��MY1OS���bN!Y7�2��La��뤜A��֟�2b�u��w���
���w�i�O�v���r0���Oڳ��d�gzb�c���-����k2��FH�Rt��'�eH?]�o }凪�f2}��eg�wh
,��Vq�'P������E8�i!�C�<��6�1�a���J��T��,uE3��y�g����� \yG�����fB��³���K��Ag<������8������z��R��}M$>���<��|�C�y�&&�q��������?}o���U�rsp���Q�P<}oN}��g��bw�E��T��r٤�B��?N�E��
�r�Oڵ�Y��4����'�E8�Ri_��?2��6ú��e<~s>N$���]M��6�O�lx��E$�/M�8��Ϲ���T�����x��XbO'����%f��{t���YS���
M$��dYm��1�g�ɴ��m!�޵8�P r�8P��5+o�H�^���8� �g�C�N9��SL>a_�<Nk�4C�%z���C�(��;��=VT�9��H{�T+�dn�Ʋ��p�mE&��E�V~a���>������x'B��!������qٰM���)���W��u�,��������V�()U��Ӧ=֖��)����5S�V��מּp*�����2�Z�U.G��p-7OZqB7x�x'���g������F�����u(��[��{����������@�m����s'XT����	��|Ɍ�Z���+����	P��&�x}@��Vm6�C�� ��<��I��U �����,ӌ��2Mv�!
�'?�-�x��E����������Cv����4�~LC�+�k�>CIVO��E�N����Ru
��Ɉ�QaXT�l�>��J�a�����
Ì<�`u&T�x	�[��9|�g�%ӿ^^G��\C�{��z�Rx��Y?2��a��<C�f�+<I�9=�E �2jo�m��
�uwl�M��l1�@Ĭ��X�(�u!濁�'#��n��e������}��7l�Ɍ9[
�h6��~���d�
k��F2~q:�Yr��i?2z�l4�x¾�}=�yH,��_{dި���&	8���7��_��tw{>���Y�R<2�â#��l5�����4����܇�ҳ�M!��w�<H>�b��TYXT��4w�
M?�L�ú�C�J�����O�V~d��sD+XVs9m靓'�C%���X�g�y����|�`m%U@�*i�PY�~�@��B�g���3��Cv����Vm���i
�w����0�b~�*x����k"śLa����{�O�V{���Z����V��ou��ź�#���`��=�I�+ua�Q@�=g��4�Rw-`]��|ɤ^'5d�m�����<�~e����0�X}��Cy|/���Lqs4�AO�>D�㟃�(g����wo��D}U�s�La��1<��{�ҳ����iE�A���q�'�{�N2�:ɉ��Ϙi'Pm��o!���J��5�
u������8���M9�<�4�;F}��W�z��Co7�xǆǄ�G�e*o)���?}����QH.��>@ؓ�eC�H�H{�|�1!�����+:� (���q+8���~�Ci��;f�gXT�߹�}߿^��J*&>�ݍ��,��=0�8��=���i?$�?3ý�x��Vc�G\��W����u�s�y�6�$��7�1>@��73�Rԅw�8�H}hz��L>LC�(I���½����"rgjV���퀼��%]���W������tJ��B��Cu	���d�5��1��x��_k��Q�ѡ�����һ)dSvE�@����ܻ^aH]K ����o��&�Z	����N��]c�ˤ(oZ��O�xx  X�sz�����a����b�yO�!�,�:�y;��ۤ�
�r��3&�
�]��^P1'P����Xk�(�<�j�{��oT�8�PR.��@0 &={�}<��"�}�>�]H���S&�~���0�I�y����I�>̇P�>M���|��q
��ٝ�m1��C��ͤ>�J���U&�w�,�|�J����M�|�l���{s�s�w�DJ��͍Q����G�)�2m��9�̞��=I�';�$�'���=J�|͇�d�!���䒫}��CG=ʩ'̟ss4��4?,�-���>+2j^�]�����Ht?kZ��R������A݇�솑gXT��z��J�:ɞ�aC�J���"���f�s�;�+���L�'��_��:�Sl�P>�G��r&�]���u��( ���=Ԯ�lyt�|���ڠc+���&�
m��ri��1!��9%b�'bz��Ru
���Xm ��4g�T�h��_��t��`�T���gr�ӹ�ã���Ǿ}��6���Xy�`,�%ACS9�����
��2!��'�^��LaX{����`st��$���N�R
z2z���i2�4�ý����<��}�]��ݏ��7���� t��>j��n���1<E%a��ʆ�=e�i���u�I�6��d�βVl�d�OY<q8��t4��*z��n�HVa_ǟd�'<�m���������|��s��|t��'����ĨI�M~�H6��S_���Ci[�]���1����+1����ECă�7;�E�aXl32�=I_�=7M�=I_=�߾����Y��{�d \1{-��������N�YϮ3�J�d����P*q>�λH;�|s�6��&0;�r�Y�LO��%H)�h��Z)��>���\u����ޏ*_����y����o��}�V,����!�I���y�Rm �ߚ�i;�$�����m��
��i��Z�Nw$�?2T�>���M2o���x��d�.��� ǆG�T��w�)dh[5�U�$OЛغY����,����"2fQ;r��T�
���f����,Y�x�}��[.T�4EW����쓵}Dt1tﶕF�>�o�ڼ��9-��氂��ˇ��EW+Y^Ǜ4�����	,������nl�>LJ=�!�����������9��w�*�Ag�?��pZ��TR?kZ?2~q��
��}�i1���5H{h<�g%@S~�I�T�)+7ퟐ�'m�g7Cl<aRu?s�kt���̕�����˝����U����o�x��
=ꊀ`}����1��Ȼ���>C��f���kT��_�1��yEIS�
$��<̚H?��Ê�Hyi�N:egP��Q`q�Y�{{�}��Ǽֿ{g�u�-[�����>E_����³�s$�t?$���{߰<@QB��)��@ğ���{����a
��w�a�x���a4�g*i%wj�S�
����v�~���~�����������y�s^�x�ͦ2m��Af�q:��A�*)7�{�u����1����k�%b�O��;���&������&�Y̢��(����m���'Ʈ�|¡�N����}>�<����g�N;�֢�wO�G�=�>� D(�*q���I�;�O����HVaܦ��甂�'��_~J�'���O�=q��f�A�����{���>��E4�*J�����s���T}�+j6��->�;�q�dz`t�鏌��2z�lߟd�a�'���!��ğ��S��8��x���!S估�HV'��&ߙ=Nj��wY�u���5�S�f ��`�Ϲ���}>���˭y�s���Y�A哿�����B�;����k+?!��V�ƥf����u��{L�Ì1q�|݁�P�%z���&�P�5?so� bO���egY<�a
����0�;ʾg����,�G�G�{Ǎ�4<c�G�)�7��������T~q ����Y�cڰ��a��4��TR��m�Y�~N����ɟ��=��.@�2=�������1��-��y�Lf�d��i���P1߰��l.����l8¡�79ܻ��Y�J�=�_�
�M�I*�&���5�B����|�2�S��T��$�TX{���Ͼ;�}�S�\��韾��>�a�i�n0_��餃�i��!�,6�����m4�U%I�{��d��1/)Ru
Ɍ��(�i�T>�0PuH{l�<�
�xɁ�si�
�HT{�����;����TC�V�o�'	�����]E�%�[��N�7ݝ���bG�W��%Q��;u+��[�Ԋ�;�
dQ�����yS�	k���x�iP��޾͸+�s8t�'SXO�Ī�O�)Ub�m��^8�ǷݹF����l������<�>֓�:�s�'?R�¾�i>Փ���ed�Y7��ل��D�P�I��d;�U
���a�����!�M�@ijWP�`�����6f�5s��P"<�����	
{3g���eg{���B��W��1EM��ӷ�$���g<�d>�aXVi���@���1��s&�R
q��1:�͸�����
���&3}�I�������=�#\���V�wڏe�ވ1�Q@�s
�a������|�V,���������
��Ɉ�n0�
��'�P�����}I��C���;�X�I����PD��0%1���٦#z��r�����������z�~CYa�ϰY��+�����|�r��f���O�I�*,�Փ�O\a���!R�5M0�l1!��4��T��=��Y:ʝ�-*�{`	�y���ι��o���矵�,�&0�
��È:�2٧�9���V?w
�1���~����HT�����ߙ=N���݆3�J����H)��Ⲥ,�퓻�8�`zR�턧�ߍVM��wk���z����S������w�ٶq�����?w0���b,��hi!�C{;��S�L@QN�E&:t��{���g̞�'�vi���d�Ͼ�q�L~����^Vj�	��R��y��8��Sl�����|���~�+�u3���)�?}����TRs��a�1'����R�J��<�Om!���p�i�~�����0"<.<&��ёr{IKg4|Z���������OP�=awN�ـi�XT6y����Y�<�f�PQx�׺��I�>�y�����
�˞��'�~��s3�8�M%G���!���f���x�H?R[�{���ߞ�m�ܫ��)o� (�Ο
����܀2ǿ*J��&"��*q7<�&�|�d��rj��La�~�I�H}i���&�S����u�:�Rq��ɴ�'澑ᢪ+�G��Ǽ`q�m�������[�{~�����d�ϙ+�y펨������|���g7�>���B�>�Ʋ��;����f���1:�P�����Xq�"��x�I�>�����*�=`��`O���Ʋ�;�5��W��G���xoIb�yq�Bak��D#|o�(��;��B<oiwC���N{�� 5�iJ��v��u��p7�.6ވ��|��%��s������[t?%t�=7��yѴ8�n����gj
�����0��H�����{���~���~I_��1?��:����Y̅���+1ӟ�_��8��������8��E>Ag�0٫�!_Y�>�i� �&�|�C�~7d��3��������l澌���S�xFϽ0>�٦q1�$>��~�q��Y1��"�L*gl>�d�N�XbP+0��9����`Vq<;���PQ}d��)�
�H?fI����g;�>�/������G>�z�R'a�g�q'R�oH)�����`i� �~���ua�=�j���Ұ��͠(�VT���
M$��dYm��1�g�ɴ��fG������u�]�ݿa[��=�@���$����Xz�T���r�����W�O����|�^�滐��)>C���'�ʁ�S;Hy�T+�� sv5���p�mE%����G5GT����~���e�/�۩uJ�黴�l=a��3'�!�Cf{����&2xZ���+��꒡Y�Mgp�~aY��Z�w��u���&�UT�������,ӌ���}8��O~����e��l��B@+41_���a�x���?!Q}5`bV��o�CiVM�k"ͧcs��'P��,���E�0����$�V��ɾ�@�8�ߵo�_�\�C�߃_7��>�yT�x	�oD�� PQq�}��u��<svO̽�+��`m��)=C�g�vLg�?8�g��H��Mo�m��
�uv�6�a��b��i+8��}�t��У^��Oط�D "@���T|3g���m"+|N���cV1��J�c�W_�a�B��+9��k/�ClV�ˌÁ����FMj�I�DTW��ڒ��y�v6��/l����J��к.=�;:�z�L ���[ҧfE\�5 ���F߂�����0�#�5۳d&�j�%����a[����R�[�z��k�������X���^�O�v�H��{
���`S6�w��Y/��yhc@t��={�O�`�d^K�2E3�$���ɚy8᪬��~ �]��7w9u4s]m[:Qanu�˶���r��p�����ﾢ�Q�>h5u�zc��z,a�#lm71���.>.��h�V��A���Y'��l-�mh>�7A���ɨ{�^�]!�����(��*��v�u��k:��=/��Z�S�r.$��.F�F.|@k]]	B��@p\�<~�#��<�x�){����=p��[R����2W�B��v�K�T(���A#F=�=���]���n�2��in�냼�A���^(�Z�a�-ͺ�K��n�K�Br�2ԗ��Or�غ�15�~����;��mlm��S�PJW�\{���3I�=.�^��p��F��LdIk���o��	��E�trʁ��Z����b±��6�@�	˩�y�LmҔg��Ŭ�݌6��_�R��T̀C)Τ����{����>5�Ǜ����ĩ�"�R?fBo�{k=:�?WR�.��#�E�����^$u�o& R�3)ż}O��B�P�����η�̐:<y��7|�)���U@p~����o*O��YX���k
=��D��1�Vq0��GHM4�{w7P��h�yL+ABif��EJ̣�㡢�$���ql:��%�V�:�M�N�t}�^_'R�j\d����4<l�ݽ����^�{o&��ŌmE��	A2�1Z��Quh�}\3E�����ފMfqQS��`�W#��|�VDQj�H�ꝇ�T2�T���\TA[}Ӯ�m<�o5jbo�@�[r�@b��9���Qr�����Ʈ&A-���v`r��U����+�pkϾ���~�2=`��2rx��*���H��a��jLp�P<}ts,g�](�?A)-���1Vѵv�����pmB�鹋3�]Aޏ Vm��u���պ����yߡ+Y>�W3�4R�%�i��6ˡ��.!�J!�n;�V묝6�O�� �w*�WZ�sާce{��|t�5T�q#r\!C��9
����s��ܽ22 ��-�z�X�l�Ek���C�W�Q��|�Et�C�
�%�[md������!h��5�@�뾏�S�qUt	�;�!�G�D��f���׵,��M'&��t�{���93�c��Q��:��+.��#�B�4:d��1T[��
yZ	��{zKg�����v��a�F	g��{��#Utu�Nf8�g�V �mH�=���B��f,��F��D���K�*�2 �-��4�^5��&j|ù�b-[���_I2��"���]�+&�v�+�B`�I��97��0u��ud�����	�}��)���:vf�E�G&����k��<W'���>|=��k\�;�:�;8V�]U�?z�\EŹ��RUNC|>��L���"l�ǝܼ�s2�iC՝�.%��� �с����*Ed*�l�:�UwC��ٚ[��1A�����E��[�X�ʛ���J*$�!��Vt�g,�wC�x��8[=oa��9XM(U��+���B�R뛾���1�ȐeC���@� 5��pQ��]��y��#�oo�1�2�i��ߌ�:F��O0B�L��i�����DEJ�K�8u�r�rW��ss�E�UDds���.M�;�c�"��sUȀ��L\�U1��p����V�6�=;9�Lr�4�P�+��D�8�
�f�8�#2j�Mh���~|�n���n�zX�s���ʭ�	���{��)n�t��O�T6Krb�T!�0VߣX�q�~���V�c���[��[�6��n^���-�Ɛ��MA��u�z8�0���3o&�Y:���װ��81���8]L�K�rEs�q%�>|&�p#ǲo��G�޳��P^z��	w�S��۶{���Ҕ�ۄoT�m
�]��#��_sl�� 9��X
�
���6�u��G<�E�#[�n���(r������G�����mڢ��&�qv��Jd{�s'�a���&�r���
5c�=;H�>�'x{��ԚB�]<F��F���Y^.�W4�o�
��0�����MK��/}[����A�|�nϼ[ѻ~��m��*o�+W+X��^�*͜�IM@���76ѱ�mcU�Ҥ���4��(5���Z��W�y-QUz���uW��n�,����R�u�c�+iڞVs�(U��R�>X��^�z�D��Au��U
[���w�h�S�dQ^�����ޚ�K�ez�o���*gj^	��[a[& |�p�>=f��]��w��,�^^G���yAC�&v/ؙʛ�1.ԗ]��hi�V���2ݩ��׫;���T�C�Jr�\T��ʜz���1#qB�g�`K��"6T�6��"v��|ۆǹ�mU����u�X��tu�˞�E<�st,Fڧ�B/��fC΅�=�	;�c;�o&X)DC;�،��Pb2S�=�H�1˱��HM��LUKBfwP5�x;���~�-oUK �ؑ(R�����Ld�t+.�R@�.
�"�1ǂ1���>�̞������7i���ī��h�����2� �)h�/�9���ޞ��F�.ם��˝{5�$ǟ
y�����������9Mj� �&��5[��j�T�H�zފ�eh�v��mB������}ч3ݪ��@W�I&�¨�9@X ���&�>hb��ھ�j��VN�9s�\�iQ����L�oj>�F)fe��f���p<B:i�K2<c���@���M�x�h�"��w8�� "���P��-����xY�y �vEC�a�Ps��(M��ج��>w�F��t�JWS�Z��������TB��w�g�#��e�[�Gۉs�S��G���=9�;Lw������c��b2/&���oVU�56����\��$"H����oK!�<O�&�ev/*nǑ���n���s6�Z�K���p� ��8w:��M�V6�Hs{�(��6�^ɬR˧��5��o^r��&脚׳�|���m�	)��U��,.��������kg�;FVn�9����i���+������z�v�����ul��������߹���S(�$�Jx񮗊������ݛ�
%ں��ZGN"#�}���Ʋ�#�'p��X�5f�س�P��Qz�7��*� .��}�ܛ���tV�6ZH�3�8�U��bu[���o���7׻���k��8�ə�dۜ��'1%8���b�|1����]W`�H{��s�m��d�խ�E�oq�
��V�f�u���	ҋ�������N�7kj�;�"��N�-]��� �ɷ�!�5�=�YV��3w5�Gr9��<����v�170˥��c�pp�"S��T�5e�N�s`���8
A|T�x�GN�k��$�r<;���¬��z���u��S;حy0fخ �����ʉ�Lve��q�fe��԰�EЂ"��r{�����Ś<Ϯ�^Wm��"t	���x�;h�{��Ip���}q�;3x�\¾�T�����~!ٻ�$dӮ4���G���4k�O$&+W�jI�[B�� �"U�p�ŋ='���#0GR.S����M鶴�-�G�"�=�Ƿԑ�Vo.���w��nQl����39�H{͍�rP\Yf^��WV�"��]��Ϳ.$Q�˜\�[����5/k��N]��O����#EX����ug���Q���f�K��a��:^��Z^�:�'�@��,R�!G�|Z�Ћ \�B�$�B��!��p�}u�F�������=��F9	�]SRd^*0LD>Äќ���7�8//z/mI��3��9��6�}���25����0�Fn�h��Ӗ�A4��/�%�b�Hx�޷Wȑ������E���ͻ�m
������Xv8�z0<}�o"�%���7�bZ;�T1���Y�j�F1t@�`-޼�{��~�؈1�h���-Ub��"(Uuh�*Dk+R���4b�F�Q�)�Z�U*��b����*"%�"�,�����,X���DilH�*��Ĉ"�TQJDm�"
��Š�b�E�r�DTAƬ֊��UT�R�d��A��Q�	mQ���֋Z�J9eb9lKej\��#q�UF��唩j�!��h�ks,0kk�X�����DkZ�J�,���h�*ۍ1��TUX*ѱUQDQ\�UĮeZ�Z֍kAZ�c�6��2�1-��d��Tb��EX�H��������h�KXTF�-EL�kc��T�`��qUX�J*#+UR,KKJ����b�E�ciDTV" �nY3-6Rҵj��aTE��UD,m�jT�V����J�ZRҋZ�������2TV ���*UPF�-�+Z�Ŵ�j�V�-��ԥ-#m�+Z4,��PJ�m���1�AEEa���ڂ�T��B�U��|�wN�^l歯�>����غd�t��*�i]���N�{�X=V�X4�;��k�Dn������٨̜����x+n�U-y��6�h��b;b@�Ùqr�l8飷�t͓��4��QKrb2�/w .7x�=�-�b �``�vb�J�y�2�@�){iK|� ^���6�%Ɲ����ԅd�t�c��	Y��ղ4C%��0�N�C|cf�D\ˁ1�EmIf�Ų\à�GY�|��/�v�Mn�!8ԙ������or�b��L��u��^z@�%sT���\���2�K*2�����3�x7��{�e�sj�pÏ�����h���\/����~��ӳ����Q#��(±�^���J!�7�t8p�A��g��1���O��]�m��Y��D����#>!��=�=�
��!����>w9�5�}��a�s��<?5c���F)Ъ���eD��ЄP젭Y����E��p:s��ҾW���R;#�#b�S�׋>�jdst���X��(�)q`2+�+;&E���wN�m�q���@g��(�}������JW�~�q��&�f��ؘAt
�]Ѓ�bf�������C��秦���\Y���8r�j��f���ؼ����{6Yp�;><���d-�t�7�^x{J��12�X��5{҆������\˸��]$��
�{5���w	���A�؋<{��U�2�aW�{����<�:\�3�؅��z#lM(��a���{*�lk�~���9lXV6���@��1{yK��M���Ḱ]g
��|WDY�yԭ5�#�X�z�`��t�f��x9�w�~�}��ik��v�o�V��BpC8��*b�k��C�s~1��-��+U������t>�x"������n�J�y�"SU��<���x�y���E^ӏd㹇n�[=������V*��n��`�S��؂�Ȋ 5n$A���e��W����=�a(z����~ͷ`��\����ky�����d߄(-�m9�����_� ��x$�qz����6a���[�9<zb{���i:m��jzu˗ �Ȍ������Ӣ<������S֪
N?�^�ˬLu�y�Zg`�V���H��Ν�o���|Pw���k��4R���4��!�� Y� d8B76�CάK:�iFn��M�U��F?%Ddl.��5�Đ�;=�D���a����P��GèX�Y�n*��-��G��d�$ks�i��q��lU�5�^�ܶ*�c��ݣ,������u��!t�5^�[�t�Ǝ}�{cM�q�v�ᕎR�+c�\����gwh��U=W��Z�X�Aِj��Db�*�N�u�
������F7�V��ۛ���	��]J��P�*~����8���7gb���sA���Q����dWL�b����I4{ҹ����~�PT9R��I�j/ǧ�
��O6z&8<���*2��z;�;��g�3.��,�����4��Ӱ:)N�J��2�`XGd�`)�35�� �N�䬖t���H�-ߠ��)�Z.����uS�C�ԫL_{Nq�&w�.�i�/�hHIoy��NTuH~��`PD��
�*#f��^<[���(�Md7����/	�����c��ù3nr�A��*s.'�`@Z06B�\2eH��] �:�D���T��qm-ͬRjeWB~�uϯY9Sb�(����d��ٗ�޳�ĸ����[P{�xa/�>�N��R2��swэ��1�ȐeC���RAk�2=bk����r��x:m�UdK����O���)�2�M`��`�b8"�L�EM9Wp�5�㱦�����x�I�">);5뤀���l��r���̭��n���@,���>�|�����1��*����pϷ�{��y'��u{zK�Ѳ�ɼ� �G'�#�
X���l��X�Wp`;lL`�뙘sy��Uȕ����m(s���tz;g�$W�֤v�iZ��,�%�����&����ѡf�0�{�D̥�iTtJ�� ��^�8�yy�T�W��E��S,3��6*NHW��[VP���Lt�@{ggj�
A��w����/��/�o:��Bh��$+�u=��C�!�V�~�bPC�4��[㶮��.{�r�]��3*������D���V�3_�>g�c�z8��}�<Z�yo����$�d�۬DQ�z���&�s�H�^�q$$c'�p��Ì�H�}Y���<�c�.[�P,]0��� ���r+�{�]W�\���q�������g`t�����籪b���u�=�MU\���^�@�+ü{Jk:{�i�!���*	�����l�g�T����� 6��n�}s]��J6�W�Mۅ�-^Ҭ'~��'4T��̾��{��%yP���{�B=x"�"��P*�Ks�ٵ ��5'�.�n�cy�D��ȹ�ܨ.\�ʔ�GD�[a[& B��&aAl�}�뻋ԕ+G;GE�<��^�I�k�ɝ���T�tK�).%ȈQ�����9+d��F��4T��Q�g�dn�Tl0	����"��'_��'�v��zX��e�7�x�u�W��՜.s�/�GskKଊG��n���u�CN^��]�vL�{��eh���+M�{�y ==��;JHu~s��i����of�w���� �U^�/�u�.u-~���f	�_�=f���'ܩ�W�wyS�Q�>���)��_kT��kN���:".S�x@>kc�Gl�������U�=^v��0A��ePi)exW�-[���q�� zXL�0�J�9U���x�X\��2���j�������99/l&�f����t੿��
��_N����:ȣ�T��\7���n��㾣���4�DF;҄+!\�5�2��x<X��o��m��V��]��ع�����8e����P��s�	B�����#��|V<��������*�Bņm{���)���%8czϫ$1IRŎ�0��N�[�S��d�POe,Fk���S>yޝ��y��+kvZ��	n��Ϳ�,��ʶRɎ2MAP��ܬ��Ћ~�vNVذ)��o�3XA�;�e���%��HF��sw�Q7ڎF˥cw<�<�"g���4g���fέ�����8f��0�'���J!�������hzLV<opb�n �䮱��7���-��F�<�·y+e"�WG��ηC(��vj�g���#:w���%���R}��R��{��z�*%j���E�a�9�+�56�N�I&�+��V)�-ד{�BZ��#����7�{��> }��ݼ\�4�n]�l�뜏�H�J}J$��Pg�:�0E��nk`ڨs��u�oL��9��;�v�Jع�1n�v:�ъwʨlO6TO<B����7��5]�����
�9m1t�ڇ6K���;EL�M�nm��Y�'�M�R�О�7t�vTf3k����*��V@�P}��v>2~���!)����F>�0[�sO��1�a�0z��k������^R�5�%�tC����=�r65˱u��rذ�mr%d���}Ъ�I1�,Ψ#rUK`S�u!��y-�~T��h����`}>��~�Sq����{��-�g�w�B���ǥJ�����`t��*b�����d
\A�#XL�1�S��.�LFf�9�>���R�ĲpCN��8�q�S���!��O_"*�q���&5jI��ݻX��p�2"e������x�sbh+:�O@���tR����z�²�(��>^�Q�]s�{c�0���)��]Zhx���=�,� ��4���>i�fez^���5i�G�9۸��o�=�i,H�@�:�`�N���C�ڢT���V5��Ny�-vs|(���4>2f�h�'��{s��T��7:݆�N�e��3�KX�>���$\��g��:x����zxВ��6������ܨ�PQC��xxf��u�g��Q�Q(`���]I�ľ���X����}�!ge;�E��J�(q��G;xr뼃X����+�x���O��AbN_]D�㗉���Ƚ�%w�
��÷�R�F-f^x?9|�T
�8P~�vK�V��4R�ݐb�N0��f��FK�!,�v�~n���湮P]����F1�y
�TE���V�z��R�r��D��Zv�� +��uy�Rq��mL�ل ���;!�2HS����dV���
��cb���2���60l
ǳ�wy+��7�u�uCY^�ͤ��?Be�+��Ut	�n�&�}�,V-�d�@��ҕ�%-
�m��q���q�o*�s�r�N܎���IXN���vHS��	��wC�kg������U��"��-BR�`9�u��~�Ӄ8��\��9��m]c��,�ϻ;sk\�3eHjG@��("�<!XD����z��ɵ!E�Y�U9�$�R�{�$����S��*e߄�;��J�*�S�3��P6B�O��@�
�=�&��Żu|�)Co��K�*q]�s���'M_\�5ge�������ڽjs�}&�F��*u�^��r��Laą6�1��H�:�g��Ek;�vm�瑋A�j��O�Gx���˘��1}OQo��g�U�k0�k����%B��N_������YޛS���*��g܎���d�HNj(h(�����6�� ��/����:���5�lm�b6��^��cvC�CL��X#��ȑ
LFREK����-��j�p���h�,	��N�A����x��l�3=`d� �X�i����c^J�sվ촚������(m����'�Tl�Z@X�q�Y\^Z�=5 ��<@J��W=�H�<�m������32���%#﷼�J^����rsB���9�nQ�&�˧�O]7vۮ��mD��^�uV�&���!��S�R�8*і\<*�o�,.����֚:w	�{�Y|����:]WB�Nj��LQEpf4��:juu�������x�g>�Q.�WGz�� a�ibQ�8+����"�E��I�f2|C�F��D��D/G����P�X��g"�T~:8�(��=:�`�����Q�����TG��������AВ��S�Z�-��e���Oy��W+X�[5�@�+�p�Vﳉ�����r�xP���g�!�3BW����N�D��lu(l��Oc����ǃq�a�8`�c�5�"��t��\�ۊ�Lgz�Q�dUoh�k	�,�j�S����R�RLx{�/M�:����4F�ugq�с.'�����w�  k�o/��]�5�T�J��s�t��������9��g!��]B�j�;P��쨗��G������Y	�K�Y���ڿr�C�}�}��z�E�VDl���-ʬ�9)��=ed�k1a�2��
��T�nT<革y:%lq	�D ���&aA�G]^������7L��N���:��Ѫrgc}������aIq%Ё
(ZbJ�#����q�>���/e;�x�Z��v*9&z,�ݓʜc]�T����`6}\o:{�]mYҥ������`X����'D����ʃ��]����Ys����~�W.c7��hJŅ%�G�$f���@����:��=�в�:�k�5V4.�3�l���(z$y���9���s�9�
����M)q!RCrzpVU",���(iq�<��s�;b�Y�}1�u7�����?����2�=K���_������F���L���5]w�rx�e
�O��6=�j H5��A��0�%
^�DR�#��QX��\�V���{!�!������}��cn��π��=�U+�Ε�4�mŰbvw��iO����]�^ӝ�j�����f,w{��杩{Ղ������������`�|��q?vTz ]��hpA��*b
��4#���Pv�ï���}_}�[��Oo����ؿgY���W�K�;�aG�u��4o�X�4�DTuɶz�`q�4�m�<T���u�v4�£b��vxu�EByNCIS���95~��̲Ε�qߡ-S�f���߆g�+b�<O�+ųѕ(Fh�nb7��D�PΙ΁EB<��j�wz����^�q��<��q�# �#�� �V2k�]!~�QqwlWX��.�yf��0�e�M`��v:d+���h�J�D�CX����宮��y°dӕ�������r�
͓
|�*6]�"ݧa�u����ݨ��
,E�
՛�q��u���r�%�<��^��u,J�-�#�Sъ���l�s`:�IEz46aK�m��ƥ,S6�l���R���!RZ*���?��������!)���{�����t�i֩��1�Z��&�;��&2���Kht���W�����{CX3��uۜ�WU���tM;���'(ws��N�J]K���Ll��#&��q�5���@�E,�������Id6t�5�.�Z%s��h�ʙf��6K�2�Dʋ�2�i���a�`��v���
C���Ӫ�Ad���Js0u���k�+�V��]dN9e�MK��-�j�BO#8$��"���&���K'�����H��.���Fr75o��u���1C2IEV���WeJ�aF��슄s:,`��2ƪ��aU2�=<�7K��z���i�����Ab�:,�y�RjK�e<BД_%e<�}�fk�3U���\}J�P�u�I���5���n��4UrGiՊ��s���ŕg.��Iu;!W�diNȲ�u�����b��[B�uE���7��ɞ�ƽ�C�&�����JC0�j�{�dͱֶ�v���+S���p�w�f�MǍu�w�ٷc�s�H6E;�=��7wN�c��->�OS��)�ѳR-�5I����x!G_<
��l>V��ǜ���;�0\�X��]n��Xݖ���S����(p������*�E�E�TX��vby�*����f��pT�
#����=nQ�t�)c��m
Aʮ���4q1�s��hC�p�Q���_;T��u��d��=����p�[� �V�3��\{��O�v�o�݃�N�J9w�eM���{f4m2\Iie�~����GU�Ϯꝁ�Y��nݩ�a�]_	U�.Q���a�s;m���ӷ��ބ7�c�D�!�|����'F��e�B�,�-� ᳎Sޘ���E4�z�����2�c
��e[���y�}}�N�Y���b�ɸ3�k�u�F͋���j�}%����y��a�Q&p�������Y�$�f�y	'�
={/VQQ���z�ȃ����n � ���J\�у�ӈj��9��BH�پ�os��Fd��i:����$gzQ����5��vb�.-FL��=fK��]S]��,��z��NJC;�-8��H辎�6
S���EYu����؆"�KR\z1�4X��|�<_Z�FWe#0Śe��b����]U�5�t�:'+���Kc��9�����D�P�\�͙��aρ��.>���ٽ:s�ڪ��l7*{P^u�<.g�N�[`�Uܹ�.W��-��$����]9k웗��`ۏ#�����d�OP�Cü���Ѕ�h��tG\�G*��*��es�p�q�βWw�ꫳ�n�{d��rz�k$�(�*(Hx��@�?-b�j���{��i�j����V�T�?s~���y��_����Y�2\6�����]��R{Ժ�^�}���v������uңY\OI%���K��k�����A/v�G{D9��x�<G�Ũͅ�Ҳ�Zsr�x����qY�Ӓ�� n�T�Y��V�f��V�k(��N�+��l���*�
M��=����ݶ����We��:=H�)��KSl��s#�u�Wc0����vXw��g����>��ȡ��|5J��C&��S�����Ä#`UQ�[J�J��kX�mJ�ch�h�T����U�5��X�-
4B�TEUb�V��(��*�w2��((�Т,��mT���(�Yh[[PQ�J�5���EV��UDVP�ؕU"����Z�m-����eF4�T���QF�ƥ.d�UDĭKJ4J�mkE��Dh��EF���5�P��hUXֈ��E%�*UF1E�V�+X�FU�Ukib���Z[k*"DAQ�m.P�\B��ib� ��ke�X�*���h�UV���+--bQZ��+*ւ���V,--e�ն�3¸�e��т��F.Z[YPmb����U(��A�B�����.\Vb��J�J�m�U�qr�DV�\��D�mq�6������f�j,*Uk*(���F
�e���V��J6(��&Q��J��+�E�����J���TR�X(��l�iV��j6(UQ����R�e�PkVڱq�Qil���[Zy�>s��O1�y8��L<��H�]�:a�5j�ܼ��-"+/rN��ʬk�@���v�Ӛ$����)Q����g�  ���z�����W����P��<iR�w��_!ZxmR"��lyg��RJ��.��ᯃG�T�<��yg�Bz��CN��4z�*��oa��x1����z;���V����Ν��)���}\X�!9�D�EcV�DR6!��i\,�v�������{�*L>�mǯlQ�ƃ��L�]Zhxʬ�S�*�y�0p�D���2���Ԟ���Ӧ&Bah#`����y�X_I�b_���V'�)��= v����U�uq�ќ�nN�N��5ERD!��mN3[�xP�ȡv�����s�F�6鹊\�=#r���(�]�n���Xo&��h���C��t
�vA�8d77,�.3�ww$`g�vf��͛届(C�elCD�=	�����z��ާcg���0��5�\}���o8�/�㸤�W��tk�# �ڇ;�-��*�cc��]���+�Y����b���S��/�]֙���b�ϝ��R뫱��!����7ǉ�G7ޚ]��ǚ�䀘��}S7@���
iEmwf����n�¶���,1XxV��ML6�ʶ����D� n){]�^]�����3-�9ٰ��F�dѼ]�I���`�L�N}Ոt�����)P��i]N92Z2r�l+5���)�߼�t|����]���kYЃn�n�^�YT���Gd�N��T��+<w�L����{�ڞVs�JG0:ht����9���-B|�X�FT�U��/��ꮎ�S���o!%��ܻ�����L�ʑ�G@[BlV�I�6o� ���°�W_�;v�b�{΋3�$��p���1��O�j93�*�E�F�puN$�v V��Z<6oԨ���;����v���l�ܞ��.vV	�dr:��5��!9�����Jpb�¾Nd��+$��L;{��ә*��E��p�ݐ�CL�\��`nΈ�uJ�u���Rզ�LO�b�ZK<��RL�Ǿ����v� �_?	�u������	�44e��!Z�����#��;C8�);5�J#"���ɥ'2��鈖��D��]��G��c��/8��g��٘�R��.X���B�<P����x.5��t�v���=��vp��1ڍj!v�X d{�H߶��K|A9��m#,��xU�{����K`���������mr���;�/!����R�S.�v�/������S����'mn|tg���a�.��^�L�U�X�żT��o���v�nlp-ƹ��N���a��í䓟h;��uvK���;B��*��-�]3qH�W\�ٿ� �,�ef�#&?�������P�5�&(�}�Ɛ��MC���X�j�ܾP��O��jn_Y׳����7CD�HF���8���l�{"��q'ə��Uk%���P<���[<zV��XP�`U�\}��T~;��E,f��W���6l�m�b��l���c�m����Q&�S�TŹM�c�YX'����U�ӱ0���N�@v��Hj����W-:jj���$9
A�g�Ɓt�X�P��r;��V�X:k-DpJ�On�ܦ�����.wНR�q�u�D����}=W�`�Mc/3/���7*\�JX4l��<���
J�d=tclb.d7J-˗YRЉAlu�l��
����w8r#�]�r���(���t�`h2\��GEj��ؿbg*l7@Ļ��K�hg���r���GE�BcI�P�a����r�\X&����]+=%�*��
���؂�1�ݙ���tYx~�
^�u�����]���֫�C"�_��QV��[�G@�H�<��Iz����Y&!*�]�$�]{�˕#�Wv�ɛ��A�g��z��[���Z�8��8���;+�]N�5�7��\�&�?����f{���;Z�I�p��pP-��G���G{y��FGu!�{E�	�5��d��I���V�B��v�3B�9sB? y�N+�hTl��hYP�a�^����|+�>���wq'�V�G/]ź���Q�i�WG�p��4�+<�mEO�^*Z�uV3���n�oEs푪0ˏL6x�U�X�~�� ��2��Ra��Wc����I��vx��~�N���ݏ��4��Da/��MB��X���1�u��K�H����7��@��%�7}oQ�:o6u��Ә�lb5�є�%��fN�C|cf��5c%;��.���^^�aoz�(��X�����<���TlX�ݎΣ��a<�!�J�����Ӣ�����Yp-(L4��n�u�׌�#�c/	�An�7!{M�Aޠ�R0t�u�Wz;��5��-�P��{�#�4f�3�O��FAG�5�P�&�E�ى�>��{�z���ye��e�V�qEB��#[G�Vy�Q&eCX�y�~~Z��J�x����9Y�Q�[]5f�Y�ʣ��:���@�NÇ9]������eD��T(���A{¦���RZk1��+E��T�0є+��l#}���
�Πgs�dv��mrk�o	�� �؏01ep�o3Mf��.�G���[�\�W+f�o�˂N�u�<����r���̈́(7�9$T.�ov#F������tbS�����T��}���|YIwY�6�F��v+�N�Q^<�خ���$1Z�a�-����X�+�1��ڜ��U���aً<-Q��(m���T�hu�|�u�<v��!)����q���N�&�c���{��G�6�k�I�>]�M���=�<%�5�=(���vX #�rb��N�Jx^�a� ���AԠH��R@{�b ���ɒ�:�����a\��n<�Vu��1pj����y!>�����X2`Y�>��R)�v59�I�VR�}R^���X1���qlצ:�Y8!�YS!ǐ�Q
^��j�u}�IMdu�-��{h�"��x��h(#&*[�;�\X�	͈-EdE�Ĉގ;��t��/o˙P!���W[P[�zk󬘽< WR�C�Vo����ő�Y�0�*��i^{���h����u��������/�(�|��-�a��WLB��.��:���[����8Jz��m�R8G��YS����P�ȯ]��t��P�׮S������~���)H#+��T���>�c���O\;�.��{�́�z��s�_��P5����/����֋�Ȭh��h4n�\������s�RCJ��o&����+t����C�MP���tJa�:�5��i��)7����9E�ϫ�#�{w�(�9��0]z+��`�^��{�k��4R��,�LO��X����q�I�������k_7��t�۫+:!0��sB�#_Pٚ>xv$�����F.����C ��+5��X�g6���Mŭ�k`W�4>��q�>�r}�B!ԅ8���ݝ�����W�������9z�*�g)~�'��(~c�gPαc�;��~�S�!N���D=OS�)��I�'z皃���0�����]��8�ʉh�V�>�i��kC�}��O�+#�=�ޒ�r_{�0~�^"\"��z-H@>U]"�VDg��69�ޘ�� ��cn^/rSBV}Y;2��b���ԅ�j����Pe#P��ǆ@�F/ϑ��[�9�i\�^���m`�r�o�'�2��s����Iv Uh��
�<6vg�k�Λ�X{̗ѯebգ�k`lWN��.vUY}��k������⊉!81~�F
��鍯 SyD��L�i������'�5o�J���Oa�F�k|�<ݝc��@*u���E��%�IJ�wmy #��
�}�Á�=��[�}X���SKwI̤%^֩.Rn��
�����\�沸G7�S9Wzcn-u��j	A����B�����7U�m��8���k*[��r	 R�u�DD�U�c���u)FEw�r�ɾز``���)�;ϕX�F�o�	~^8O[�zF��b�*+;��ZѶ�QC98�;��~]�b*l�R�k����b.s�(�6S�W��M�ۅ��n�\�鉘O�r�Eb���:����D]"�}�RR�=�
��B
��������L��d��+-)3<�u��.X�_TC������D�}�H[0��pU�2��i��ȚosS�
��Lq=�b�T1�1�W	H�5	�&(���������:v�Oo,���/��b:;����֦��:8�0�A�}���D<�+󂸻�9�S'^�e�J�j,�f�ߒ���0��ގ�n<"¾���k���H-A�F�
E��@���I�#�vܾÛxzk_(
���lU�ߙ�cWEϬ��@u���X�A��#����,���{��yVl�T��{]2|�(ʖ�婋��#V9´:�����
ۺ�\n�[��vVvQBC�^e'n�Y>�F�X���_޺k��Ю�P�Z��i ��N��&w�\z#����J�\rƑ�	��5�_�gJm[}z95�1��ox�|k���)��7_��]W4k=�#��N������[���s��=�et�=[����f5�����䊷��f���6n�+1�g�x��>��Ϳw��[��϶�I�ǲ��1��Ê�(�8革y:&��XN�ʀ�,�&�>W��u����U�#�S��S���R�;ʰw����-3�7���~R\Mt�`����P��B�ޮIEn���ц#�q a��j��_����>����yxWg���zE�B�S�ޱŬ�ފQ�B�� �e
���WF�}5h����r2ȷ��(�=vqY�[	�/��T3������:��=�в��ãkޛ�JH�ޝ:�D#�lSJ�ry���O��Hw� ӫ:U8�E T?i��nZ�¶�j����H׏?{,��!l��\����b���pj(	�e�� v\���;�;l�o6�X��j�],nW����VU':4MB@{��N�1�x�(R�m")zRՄ�`�[V��]�?"xp_�7ÞGCU��X��kչAȧ,wTN��Tdѐ�o_�����a�((^��_���j�c.�FGan�gQ�W�I�߹k�^e+�{�M7��������ů9[m��s�^�P^n���l�������g
� ��:6�nfuM� �"3�̉��&+���qvY�=����r�ã@0��W������8)ԋɜ�QUK������с��OYrdJ���Uy$U�򎣳�~��n��#,��c�B�a�O�<-�O�|��k���*~��-����@����N��3#<���<UG�a����3F�����W��d�q�3`�VMzpU����W���1z�gP�j�!I��EB��!������DŃ#pr1s�q �4�:JwU�d'x�e�1�J/f:}�B���}���r�-OT6'�7j%�
*�n���e�X�rj���[�V�9@٣`L��|'�tW��^�����Db�2:�"�ۮ9��6�&�]���w��\��\C�Tr�z�d?�(�WG�U���:�d%=G�f!^>�p����8�w7���N�)=ˠW�6+�5U��J0A;
�{*�lk���!�A���k�sSmާ,Wz�׎Q�J�!:u/`J��!Q��茛�d]��
 Ic�o%='
��Qu��z-K#��6{Ԯ�v6oj��1�J�H)�����Q~1s#m��7����z��h��>.2�͌��JNe(��}Q�����w�"#U���D'�ǳ�Xϸ������*��B�`����d��#�gA�b���R�a>D�[�6׸7��~�h��u6��w�yt�o����op�E�~������=��#���f�G�3w>���|r�[����N�lg���t��_h:OH<ӑ�^o4�
��q�F�Prb����>�,G����{��N�+r�\�.����b��"���*�r�j�.g�gJs�� W�P�5��
�DU�OLJ��0�a�ss�w�4��* Vl��R��P�=m�bNP]_���؟��i���k��l�/o�\Urųo���\P�n$UN���h�,�����q�Wh��uM���9���f���!�t�ŀ��.��?�nYA��'7�*Ѵ4U�Y���#l��`�7ӎ�����g:\�oqUשf�siD;
�!�tFF��6f�V�����ы���50��9v�w
���7��T"憐'���8������*�ccvv+����26+2�i�h-\l�;����T�C��gPαa���h��?����
tng�S��vɐ�ӇW�vޗ-aξP'_+q0V}Ǝ��i���KE��K�����ӓ�]LB��6�8}o�j�0�	�]�R;$%:g@l#�aH@*��_�VDl�hP�S�0�o��R۫����}�����+Mv�1l�bj����ƻ�7��I�/'2ގ��WXw#Ά�>��oK̴�[Kr_<*��Y�հ�x���<;�αz�j\���� ���Wu�6a$:,>~�.=�ܬ��N�<5}k"7G7S�]����E�z�m�����˫�3ơ�v�o!�)t9��+�)CA\���z˝!�F�Qns���7� �+Sf�.@�;���pmM����qr�{\�B�{j��O\uW��<1գ�,Y7FG��f�B1y�w�;�)L��P��kfb��pR|��`1��^�2v�p��xQ�N��}!��^���ީ�Z):�3�g�'i��ԩ��n����t��Ŷ8R�����]3�xVP�,��蔘}���Z��y�ޢxvU���"U��^Fm���j'
�/wu���9�nd>}���!#��E�Sչ��+]���w<�)+6BG;	q|*����>�q��Q���Ew�[L�:sjo��	�T(���Wv#����|VʓR��{^r�;&�h ���m>�Zsqpe#H�{$�ԫ���}� \Œ:�N(Wf ����i#4�x 8�#�-4U�{�%�au�I�ôdw�QL͈;͇/{����r����~��SI���+/�e��ef+[��d�ԜN�f�v�����fXލG-�o׮�f���S�^�Q�U�=�F|�ʓ!n)8V�J�\�ru4/n��F.*\�S�]a���a t;�2�������i�X�s�y�n��=�Ճ�Q�~�<�w@�zT-���B�����4���Ն���os;�X�I��w��1�|`�3�j�^�B����m�7��ER2��v-ѡpŞG�yz/�Ж)�\^�AK�"��DV�^ّ�ٻ�:�m�]A���GT�q�_�X�N�'�b8�ɷc4K�� \��U�;�v�s�ݳ���k/9Ү���Cv�I!H,V��Ø]�gS�z�e]�Xʤ��~�]�شnF58�V���Xn�VG�KU����f�sCsV�A͟I����)|mWJ��s�z��_�8F�fX�od��ʟ	{�Gvh3�xxj&;�4�>�,kΘ��y�S����N�F\G"(T"v�zp�2����h�;��L�6啛zyX �^���e����@��;���G\���7���Pqۼ�{��p[XH�jN�HZ��Vty��4�,]�!����%���SĆ��c�Frḃ&�\;���6����2����acSP��ڷ�y���:#�Ȧ#�'�k�{f�W#���K�6Nn�l�=:�t��V��>B󈹦,�f��3�!�"{�Yv�+Q����X����LӛD���5�w�֖l��ҹM��lp��C�G��sv:π�� ʠ�jU�R���PD���A-�ե��������%k���X(��5��m�֖�֢����[c`Ш��Jʴ��J(�UD��УADEQ��Q*�h��UE+m-F�[d[mh��"�k�[T1�h�m��cm���T�+Z����J+-
ڵ���"�)RĶQeKmU�Q��1j4�[Q�J�Q(6ҊV��Q"��4��JTh�6�#Eh1�+mh�J�-1��U�-*�ڵ��ыjUQZ�T�hT��1Ɩ�,Kj�j�IPZ����!Z�A�R�mem�T*�X(
��kRŋEX��h���(�J��ʫ[J�-+U[Kl�,�X�EQJ+(�mkV��(�� �ڥ�Ub(��KlZ��h��V�-T-�)J�kcK�acJZZ�E�i--��Z���Ţ�`���5�+j��J,U-(�R�[E��mX�Dm��UJ�����(�J��]2��Z;c�Lq��MNc��UDP�8��Z:������ i��p�e��B��0$�ަ�S��E;�U�Q�|���d�}N'3��U���ԋH��[�+��u"�"����ϔ,w۽�Zś�IKs}#��	���#��Y3�*�E�F�9��; *�`l��n����D�N���;{ǳ��;����9s�
�	�g܎�����	�E
*&;[۾̃[�����{|q�X�AT�H2�։���V' ���u#jg�;	�:"�L�׈�Vʍ��8��ީ�e��h`��r�}������K����ua̺�X+�<"sP���Շ�f�k�r8"�I�Oʀ�g��E'f�����S������V/qRqU���u��JwYՑ9�(mT�
�9�.X���1Y6���Wh�u�<D:^u8��bhNb͘U!�������b����(��5j_	��hs~������M�S�=��d�`�>�6*�F�ňB+$8c���B�������V�3�����v������d��~#×kz8�aAq� ��χ+�?K��N�'��J���d���ښ��58��d��+P�L�O����=Ls�c�����l��챭}�)��.��tflu�\Xcy'ٝjv�\�K{F��&��Mʧ+;4��ϦkL�:Z����Kk3�_>��y[1�h.ԬٝMp�y�d����\��r#ެ�M^z�̺ksޕ�ԁy�������FGl�m	��!&�K%^j:��7W�]�t`�F�^͆h�~'�±�[�و[ '\����qk�Fy�mr�{e���<�Ι�^�����Ol�jb�Pv�+E߽Yj�jz�sRI�襛5
m�բ��U�.�%l�1ѕ�c�(�����^�¸B��Ǟ����7�2N��S�i�}����)�lڐF�1��̎n�_�{|��K��p�uػ��*�RG��2zd�3WP���ł��b��/�:��Fq�pe���>��0}G/6[�q�%t$E���Opy�P>��P�6�����$(�}v_���8.{�Ń#vO�o���R�����@�]�`m&��f�u�{�B#ed�D�Q��{*	�.�WGZ�L������3p��s;yۗ��W�a�0A�O&�X)�)��Z8�#&�ʃNSs/�A��nv��%���D]Jc��̷!�:03��ʧ�
����	��������~P�k��C�"���'2�$y�@� �O `r�<W���g2�g5���w�H��;RA� �����E��'���G�����KMs�4�,X�q���poٺf�vY��vͩ����_[Ss>��M���G%^�d ��<mhJiP�O�7z�|���U�َ��� K5��@kЀ��TV��)T������ܢ��Ox�#��rw,���R��h�
8Ksz&�߷�P����9��*� ܨ�S��ѫ��CN�0�G	Ec�>Ƭc�������Z��a9c;�m:����W��n��C%�r�Xҟ��YuKE ���#~j�O[{s
��[�����a>�un���pV���n�u�>dm�T��,��vPu�U	y�n�W/�<�`�鿐O��_����i�c�5�o*�|�)T�=��Q����B�6s���dl�r�|(\c��p�d�)�v]:�]\⃇B����h����Hަ QQ~UA��ch�J���D�M���r1s�O!e��n�Te��jf��ӷc1�x���>��s�S
_k"݄�8s��jx*��=~n�L��\p�"�B/o57�zŏYj�lp|��)�
���h�������Uox��y����ּ	B��or�3mgO;;��ä�+܌)qa�\!X��ɉ� X������z.��\�%5�q��o�}���#�G��CL�k+���#v�VK<�m&*蒱�L��I��3�ݐ���kqg�(.㪁D��8W����gT$��d�%��*S�D�{�΋qq�elm`W��I_:N������@�����j�<�[I0��^9��&����?Ʋ�wo����U�R��¸]�k�)��̅V��Z{|�+6�H�78g�1�b½��A�J�N]N��)A�����,ϔ�LWuj蟩bݗ���ղ������إޡ��R�q�ٽ�σ5ˁ�]���������7 �^�����똎}���aYw[�K=c�Y�W���qr��gjb���؍:>r�&����B\�7����m�ߌ�7�ǎ����&*[�;�#�Bsb$��7�G<��x�^�\QVz�}JyV4��\>E�_���Δ�/CX gP�5���:lQ�[o+Yy�(^�,φ����i�u:� ��T߲(]��x�;4�2b�F]j{1�3��G�LB�����E���RDp�%^�x��X*u����b�2VW�i�\��Y�Q�~�1��70�d���d���s�{��;CE*�1@tȭ=�4��/�������X��u`�B�iD;��w�茍���3D<;|�9����c���SU,��B�a�{��6:�ͺ.��e��RŢ&��춝Z�Z�{1��WxH����2��Tgu�Ni�v&u�dݾnws�}y�3���y�ؒ��ym-J������/z�ćN�br�)���(dor�;�,5�'���|�_��:�we���CJ��Zv�����*��B����B(��*�ccvv+��x����&y����Z%���i��~��7�Y�*�lP(2:� ��m��e����7܉o��ܞJT�\�gvz�S�<���)�+]��Uюo*��(�Ut��{cL���"�֫)�Πa\������{܎�	D��lul$E!L�X��YE����%I:ʮ�ܗGdp��{\�u��%9���*�:�R-H����`��a�6w�=�>҂�u��[�\��˿4²�C���mW�j93�%C�� ZF�VT�H�B�i'��L��gzHOICf�N�z{���9s�
��z#�}cY9Sp���T�G=|�SyV�R�u�������Y�������𒇖���A�y^ܧ�����6��,6��n�os6��������J����*�v� �_������ <�����q댪�RV�։�Y`�s��5m3��ʀ����뤀���~T�>.��~��i����L������̝B�������+�P�2���b�0)�{�����������mlB��A�VZ�M٭�7v���
c7���Tc;��x�}v9�F+L�Yb���� Ŏ]���N�)�[i��Kb�Ab3�i������n)��)���¦.o�T�
�9�.�L�DLVM��g S��[R��m�7���Z�G��e�=R��]��#�����V�S�
r n+�n���K��#84���ۅ`8���a�*�!�w��K����>i�,��{90/�����w��!�٨���U��Gfa�@��e
!�_���͘}F��R��t�v�݊��Q�Gq��>U9�x�M��	��aE�0�)'�;)� ��Vf�]OM"�ّD�+�@����y��~w[��JY��1n|�!��V�`h��q_{�3T6��J����X;Q~��Y���%5��L��(Q�l3��D`�
'�Ŋ�k�vMռm��ٺV�N�K�B=��^drV������temX�J$��>�� "9�Ǫ&]^t�i.���=�*ȃ|}G��9�jA�F6����ܨ.{Ιږ tO�hS���������Mn�Ő����C�I.,���;̕:���&v/ؙʚ�I���KZ�.�Sd'b�D��Qv��sz�:㕋j���ۮȢ�jS�$��Db����37:�F��WɅ��gP<�8�k]�_Y��Pw��.]L�_Tj�˴�@q�/��r�	:\���9�w������ouY�t9��4l��5�����P��1
�d��B�$G���)�s�.�����F>#ͤ]}̕�Fr7�Dh{�B#e'D&� �Th�8��9�/9>��������R:�N�^�;��ie���0A�O&�_�D����:��=�в�������F{q�A�����\��;��?���}+V�e�aрub�|U8�(R����z'g!�B�������[Q������bR����[��-$;���hs.*ޝy9��Ro�r�e��4v�N�͓�^��
���:"a��X���1�/ ;."a�CS��Z�zy���/"��
�;jv\X�ӻ+|k#Nb��x����E{$�b��aᚍ�O�۾����N^�U4ZV2e��������hl[�NƟf�-�Z����d��S�k��3G#eʙ�z��J��sQ��2F��6�x��G�^}QE����U����Z�SQ��6y�j���@3�Mñ˞t-�ҙ�Jޥ�?m:��Z�d׏x�YUx�͞�dX���m���:�ՕK@c���K8W/����Zζ��k���:�O+�S4h����=<��c��;�7n:���(��y�E�(&;�E�N�M.��g�dJ`���꽅t� � �9��{�"LF�Q��־�<=/a�d�J������ٿ�ە�C��L@(��L�s���OT!A]����i)��O7�(/R�\�D\� X}�'��M�ֹOl�b�d5���Rڃ��_���C�ߑ9B���:���)A�N��ʄl,�jY׺�U7ܷw��+'�OE�d:
��b�{�}�|�����&~�<��I�u/yB#\�6̻S�K`&���a���{Ph<֭���ϣ}��W3�Ճ�C�Gbw$ZFAM���js��oxc�K�ܼ�-�[\fnV5Y���o�͜�i�RP)8�uk���� i�{�C��q�T��˳�^�m؇Vw"�"�wt�ל�>����l:4Ŕ2|�����i�[��*j2�GD)V���A^���ݱbky��(k"&��
��m��Q�Y�(`��c<��L*�n]��;�mL��|&�Z�c�a�E��m��>^ڼ<V���hX��[}w�5����N�5�OM�g��g�w�����jH�C�C��2G��9�5�*�������H���5�g��n>e* 1V�}�g�� �.W��ĕ�F?f���q��-�dD�[�W�v��l������[���=�,�:�4>�ui1�D���hl׵��J�����13�8�i״�}-ﾕ۶6���0yc+��y��l5q�#p9SoV�w�X�%�^l4��onБt�cCsPd#l�ʞnx>��>y�}R팷��L����w0T�%�S����t3PE�c�k�9>�_%���
�����E�z��M!l�6��D�����V�Z/�=w��-rʾ�Ï�<�b����9�\B�ح���[7=^�jw�츖�������*8�q6��|�J�=������VWE������3=�=��azuI��H}����8w/��W��U��(u���+�q�V�1Mv��1��w�<H�n��j��1;�J�s��h���35�I�)C�b��P7�f��V&�엾����#�4x�����`0����l�P|��g>����qNW�xl��[�*)"wѮsq���Pl�z��A-�jtXK��5m��|o��b��E���LV���Ny�6�ͱX�u<ˉd��z�7]�O��J����G�^�;�Y���W.7����¤��CKY��:���kڌ�]X�����u�%V-�9�/��Nn��U��ܳ��8����BPU�5�� ߎ)�q��i�ۍN�<"E�wb�]��If"'9�ʍ��Н��	4�
�5��+(d��1�1�p���xVw71x�em>�Ήl�27�DBb�Qbhsd�P�}Yn��.��[w���b��:]���C���&�cQf�����z;u�w���8�%�^z'��'�4�e!����Eu: <ѳGb�72�D�/;�.7��q
���A���@]�7HaЬ(3�B�<2�f��	�;�7�8������\���5�C6�d&�(��t�A�=�#duqԍ婗�����j&�м���4�ޠ�{`C&s���}j@��b�^�ʵLG��+|�k�kv��G]?�l�;B�l2ٷÓ�^�s~���N�Oq�����.�۔j��2��҄ҡ���|���6��6qBІ�F˅���X����eu*u��1��	n�Z�b_x�k{�˫��9qc�F�x��ӗY�t�_�E��޼��[�T��j�|�X�>nSw��}���ˡh^�gi��z�n\c2u>M"�Vo�XXll��#m���Κ̥۬aZE��:�uuL��v�:�i��-�ngX�!��j�"�5��P�iv��z��`<�K&��o~�g�>��JA�x<�F�N��nA7��JC-���{5�����ֆ/n��7�������[y����{D`v�i'�mn�
õ��]k��<+bO-����n�gj��Y�CН\|	��\r�R���m��ȏ*��"k*���u�\V:֛;�j	�����s�'q
�a����WJ!V��6������d�EY;(Y���d��q�i[Z+��\H��#�v��nmo#��n�W���W³
����=��Ъ����D�I؀��!�5zr
���Bl]��Jn�>��W�8����]6����ᾰ�	��Yّ�L�N�"5Y��3���
}�o+X������dEzB ��e�AK�<Z����m��[�	�v��������vlE�y:�͉p4�ڲ��,��p�	�l�0}q�����!-��-�٪���5�m!��#v�{4F�� ���\�R�_k}�$b�n���n���++_�}R�+�;jP�{%*wI���p�Il���m�����-��S����Db[�Zxb�d;={��p
����
�B8�:��Ե�v�X�[R�
�GU�o��@ޕf��bd�;4剂��Wzͥeq����+�7���t)Jɜna�Vm\��l��k.��9�0�e(�Q�˫�����ã �ͬP��c��	c��ZݑK���/�ަ]���iDaRɋ�<��E��.�р�Jغ1�76���+�7Nޙ$��]��r�o,	�/[CQ�I♎��b�<���wRQ���G�[�k;-���U���K++^f� d�h]X`�S<���V3 ꖏ����*+ �ʻ�������x/���%�e�%Oxn,y����)%�pu�}��x�����Xn_!�{�s�ٜ|mJєz��N� ýZӄPO�(J,v�tj���ly܉@'����%���� ��D�C�N�3pJ�Y���sRe�E�kNHW�<s��z���O��}��&Y��4���fs�s����}��}�S��I㑮��#��ՌRe*��cӏK$��#*Xq�.̢.$Q(W�%Ш6���s��ǔʌ�һ�Z�u������G( խ^C��p�\'Np�Wh�o���{���=mbV�kF(�-��ZʅcZ�RUdPZ�JQ���*(�ID��4m���V�P-j��ƫmF,�V�UQE(Ƶ`�[l*X��j�RڌTKJ��l���1��Ir��r����.%p��JZX)
��AUb)F����ȥ�iJīAVh�b4TDZ�Z�����A�J�T+*X�Ҫ)U�"�V6��l��U+Y6�F�
V���5���J�m�cZJ���aVҰ�ղ�DJV5U�X��
�V�k�RUJ0Rբ��n4�D�QTH�L#`��YD�j,m�҂�b����,X�j[�*2QR�ZYFѭ�b��KcR�J�KX��*%��#[l�T[hТ�+j��hѦ�
��S�9=�ܶ�Ny��-jY8ڲ5����xe_9���r55�Q���ѧ�#�ڙa�T����`r/�C���>����_����OB���y��t�{�^vC��\p��V��#���y��<�Aԋ���l&�r�����Pv]s|GN���.�/4X���eأ�^,&�i\u��ͫv���Эif��ծ���ކ3#��U��b�{�]�T�p}��Yht����7�5w:s�۹�/�2�)qA�V��|�*Ɏ�l�Vw[Zx�Sf�%�٧kd���{Lg$�Q�6��[qA�kڴ�D�L=Q�:*����7�,n�IX�y�X:�[����y �Jp�ֽ���.TA��"�Oi�XV����H�
��Ͱ��O�)8(%}�9�z��J�צ���u� ����H�`���3��L�E��ޞ��e^<�w���<����K'�Sb�Y���>�m;V{��uJ�sՒ���O/6�v�2A�*B�;��m�.kn�N'���^ɝ}H�Zҫ���ݐ����܎��<4ӂ/(jV.a[�W#T���)����+�9TʕwÓ��U�q/��E��9o�N��$�f��s�����f�X��=��.��M��zu���ʽ���x��ӕv��l��C0�4��IT�-.�QH�[qlwS������k��z6h:ݷ���<��y����8�ޝ�x"_;����ޅ����ɢ��{\^�*o	�VU�ɭ<7)��|!����`*ч5��a#l�Z��95�<خB���9=74r����F*�`%x�a�Ƿ�
�:y��A��"IF;��Ҟ�jˆ��\v�H�ŸtV1�m#��=��p���	�e�ۋ��4��ә�gK�]�T��:ҝ~IMaqT;�N'�Q}E�+���n#E�����׋�5w�xa0��_��J�=��nG�W`>�b�u}�|�ݗ�t�hG�U�!�����|���b����}r[fZ��`*lpeW2�t:�n�Cb*�N]�N�[���+���n��,�щܑiɹ{e�jG�����{,������ˉ��K;�}���rO�ͨ@� e%*$.l����7ӵoB|�g�������=��h��Ey��
�Y��v(#��;۰i�|c�1{4����-y������N��Q�!����oB��oVm�x X�54pr���8�^hn�d4�{}V�
Aw����8�n�tZfD�d�*��K����t��y��F�!�>�������O6�)O|1��`%'{�zd�ƽ���;]^	��^S^8�Ѵ�	o�T�lꪺ���3t�q����5�
��YjM筹;J���&7)Čͼ�ݬ�'�y��ŵN4"������_��O/p��QA�ױ��Ո�x��W3�`�r;)�LcQ2���Cf���U�+Nڞ�o�ӻի�ݙŏi
��#�5��^m��W�#hf��)fn���}��O�ج�<����
�A�ӳ�:�/73/Y;x��~=�&n�~�\�7(�o�C�C5����eE��쩘Y��ܻ�GV+a���z(b��W��ផ��҃��G &�'H�7����إ�ӧY��.��}�lt�(@#��/����e@M�u�o
w�a�4��s�1��
�`��T�8�ob]��Ǯ7�Z+���'{&:��1��6�����e��z7�oF�RẈ6p�4co@M+�7s�2��u�@B��ML�O7�����ǋ����P��v'Uc'��M��;�����3��;��*ur����V,n:�p
z+ͅ�C�*�=}\�w/qN��aO9�������jq�{Zp�_yOE �5s�0��9P��j���Sv�E�3�؞�@�f��d�k��dq��H�����[B�om����������M�ߌ��픆v�U� ���!{g/qE��4�Ҟ��m����ޗݦA�)8�{Q��\��p����������`�Y�����i.qs��i�I��AW���P�8��g�m��k�ǈf�)-��0�S#��y�#x$���BP�"p�2z�[R%�uw^��@^�����Qe���Bz����Bb�j,O7Y(k=[���<�4\�{J'؄՞�ۤ8>�%sڋ55j���Fwz�uaۆ� ��jX
=��%ڭ�&��'$rrL������ţ����Y�*t��,�+�ǩ�釺�{��P[fu�Ι3k�����u��-�Q��Ib������:��ٻ�,�`ꔸ(����#�k�oV��s�RJ�N�M`��o@�˵yt�d��[�]N�=������z�(kvw/GM1��Dm>4�v�
ݯ]�7HaƆWW��ĝ�
���\�p��7ɪ�^Q�yqA8� >iWu���-���yv�y�{Z� '�}[�eW����iu��ބA�u��R�s�"q(����sz�f�壳���U�H�N<ܞ��.}�]v�K���ד^��]��4��'���ʠP|q�Qgɶ���^5���׸��YH�Tpw��#���GW`�"�}E��]��F'�-�f��9e���+=�zu�gb����ʕ϶R�D�6(~�z@_m�����V�@܋�I۝�����i�u��F�k�����O���q≷�bC���d�0S�X��96�H�6ữ#�>u�8L�n^A���u&R��u��B�oR�,~�i�0"ת
�F��IWK��l�,|�u���JjŃHj�:�=�1p��8\�}��:�q�j��pgu�v���!�Cvd��l��� �C����'� 9���;4q��&��5���9z�R|927t�:�J����E����Rp�{m�A�c�GrN��[�Gw�ѿ��;���+�K��U�<ۿC���_˼>�l�O��p�C����T�ǂ�Iޚ#�F	l�#y�}	؎�ԉ4��sݜ�u�^B�fI��N&���ׁҨ���B�2rqJneQٵyԭ�朡/��b�"_�f'w�˵����)	{K`n
�̓*�{<�/Ehy��eSz2k����{+��=k1Iֹ])o۷;��+[����0��,eu:/M5qZ��WJ�ڙiR���/L7�_rN��=�fӺ�cb��Am�Z��94�_}S���/K�e@���r'�(!�I~��7;E��b���T��Ǜ����7~9�qL��g)���SW�9A\pGZ�s�
� ��!6��[EDct�b5�G�j�M��P�����Z�>���4�p�&���>rV"55�L��(s��nE�y���|x�װ�c�
�S`_!;5xYy�\vL�8��v�r����w���6��.l'7�K�,�$���Au����Vg�3�"��Y�_u���&vN�&����P�J��xOX�_QAq+���Z�Q�:�_VY�E[�&�|�J�����ʆ�>�x�����[j�j�����D��G��;��ݿ}oL��2�th[68=U�:SJ5l�6�sv����-�ۙ�]��`�׹dq�6��Cn)��mU%�+�n3wi��Y��?mp�'I��p�v�U�D�}a��E�d_j��Z��Ί\ޫ�͘�:���dn2D=x2V��]��By�Ƕ���R2x��kS�r�7��\���^C��R��_p�41)q��(�	;�Q'��Z�ŕ�q5��p0J�N��([s@�Us�E�U�l���a]4%����y�a1mA�hESCY����x�%HU�m�F���t��Q�h�n�ೲ���QSO�U46xT�j�pdS��c.�^@���Jm���v8�)#̽�i;̽��s��pPR�K�KbXԚԽ��a	�xnȕ�Ө�f<[�i�V-@b	�י���Mϸ��_$്1M��S<�k��[fh�u��)^�+���g�8.n���&�ZV�-���{մ��Br�]N�ͽ�`5q�K��v�����7n#����7YE+2��Af��6�K����<ɋ��vf�/Ө��C=��VR>��лA��PU�0�!���<|¥�oq���������V�`��8n����(>��:��;vE�n9�Yv����F�ǧ,����9�\�u��'(}��^,�䡿6�-Ǟ��Ϫp���Y�ڷK��d�S�M��C�+r�$�7Q�����0¯c4*��i�j���Z���%�gD�9u�VrqY�p�����Q��V��v��VG����Q115��Y�c����܅�`:��E� J�ڳ��`68����V1�_����)�Ot9'��Ȕ�8kڣ`�*�z�cx��ߤF��	�s�Sf�-bC�@���3@宮�ç��-���C{\�X�m�v�k�H�Ր��7#�*_B��껩���
��d���]%�$�c��~����n�L�3}~��+3A���ҹ�eMX�Z���u�����n:��n�t+�j�s��C�pi�)8(&���P��8��D�n����V6�N��[�'���ک�����&��R��Yj���Q�dVU4t�M�Qy��ԁ������=�ՙNx"&,���5�l���u�#�O�NkE��^j)i[��G���x3�R���ma��6�oK�C���wQ��51��*��˖�r��-��Y�����y;�Ȧ�s��Gq��뽧å��z+v���.��h]VL#�{�Qm����#�^�p�M�סy�B�w���C7�B1b��J�)�2`��'�5;Z�e�`�����سW�Y��V/nz��ޥ�qu;K!��Ƿt�ʣ�8�aW�YV�#�8�s��J���au��7WH�t�1�&Χ]�%�W�X�;a� ����M�`:X��X���#�	�^glɫl�|Z=�u�ֽ�ѻ�-�\���?�՛t�E�3R�6�0b�oO�{�'}�@��>�j��|�ɘ�x�}�r���QT+yG���oD:���|�f���>��H�x�?��vj��o�+�V�Ҽ��g�=q�T)����)(�����.���E=@���+��t�q�֡D���Fgع��k�w����L�}��ߐ���XCdCT��o�z�]���F�o��թ�~�N9�z����CB.�a�d��H���!ٲEN��9Z���u^���Xֺ��H�mƇ��j�u�\.y�7��]�i�Z������ụX:�U���N�m%�p�_��ծ�f^jvM���it,�Ոƈ���L�ک�݁��	�W�r�ΐ�.zNZ��.����l:�qH���4p���%��q�WT~���4��	CJJ���r��%���4��"kme^P��Ҩ�)��P[����o�ZO���E�����0�&�������x.�e��b��3�f�������ǘ�����٢��q�l��x+t ��ں�˷d��~T�yk5�9P��~�B��;�iNA@h&��;k�G���.��8��n���:���ܷ����9;��;�B=�Wn��VZ5�)Q���jb���&�1N��/2;S� ��qݎ�w�Jѡ���Ro��u�)y]��b�8p���ǂq:#�|�EV��n�Vn�
U/��q�'����^I�,>��Fڳ��1�Œ
�#e�N[���CN�P�hN��#%=���q$
]b�2�����"�Õ{�^`�Շ�Z���%n��@��ի	v$��_K3���jvu��ꖸ�����^Y#����Θ��s�܌U��!���͏(��9���h�D:G�f�l>�͕a�[�#V����¢��:�\�c,��_G�ƌ���:��҇�oQB�
����"ō-r���M抻۲��I�l*wk��宕u9��s����E��tA�o#s�vDI����Ӡ	�t�[7�w����y4�W]6r������.e�����@ޥrl����=� 5n\!;�,�)�Wu�쮔,i
A���On�Դ���C���]��0���{�fk�1�.����`d�kP.Q)IY}y�S۶�I�iYpI[\\�%��q]ڒ�V��lK�u��)K� ˺WG7�7x��#�D���2�X�4B���z���B���51ОDua:�l<���ܗX����Z⊚N�+^�ww�ֶ�=��c�\��TqC廾T����rg����$h
\�]�&&������j҂�M2|h�ޖds=)�[�rۜ

iu�r5�}�ʑN���Sݛ���2.߭�-�y��I�l=g;Cӈ���z$/�č��ͯ�t���P5��'h���g�쇞��D�鏚:��7��U�&���
2j��⫻�֨��8�%�5�2�Շī�.jz�Ó��?.��N���p"�R�z���^�)�6��/G7L�`������JI���zܢ�
�6E.ô(�4P�4�b]�Q[�p����Oww
��u�	�v�Ex>>����w(���R��<3j9ҥ
�a^f`�s��u +���=�u���w2�9Wg:�mpF��^�+�]�d;�����ag�e����g(u��gq^��Ȏ.���$6��i��YV�Z�׏����i$�nC�<J�Ӵ�����1k�zS��-I<#
�D'lp�轫͑G\����ޜY�ڵ��V�\x�F�(1F ��QV�����>���X'�J԰��Y4:�trK�4.��ܾ�t�y��ՎJN�E^�X�b�ʷ�]���NG��
�	��3M���8鲌u5�ڙJº�E��Z�_�wK�S������`4n���v��_3�"Y�oz}�{�Ò ��p�]ݫX��K&U��g0�ܸ�Ú'd���>`"��E��*����kjT"µ��V�*�h��֤b�Kc-hZQ�YF�%ejJ�(-J�m�,m��*Q�h�҂�"��J�����F(�(���[_�����jZ
��(���*�JեX#-iQh6��YiYF(��aX�YX�Kh��*�V�VF
�+b�XҭU(�l*��X�TUTZ�m�D�����U�J�-�V��B�Q��jYm�J�
5YV�l���ڣl��ʣ(�6ֶ�lE������)J�h�dD��8U��V�kX,m+j�B�ԨVҒ��eE�i`���Q�*"De�j�,�
�*�[l��j�[
�6�ƤjX�Z�bҪ֖�K
+J#�p-�����ii���[m�**�mQ���T�-l�+U-���
� ����WG����)��u�ȧ�-/����M��L
�;X�誡���,<u�vOU���ߖ���HF
\m� z��:��Kc��^퍦2�y�XϗS�����j���\uO{3<-:�5�p�a�ǫ{tI Lf67٨"��9k�Ưf�l`�o��57uY�E[yZ��p�3��e2��-8����T��x#�o_3��i��v?N���h�U:��U�{;E�L�Ydu��03|S{��K�\h'n��'{�x�A�S�p��(.���D�.��m�)fv�~�(�(��ջs�)GF��e���U�!�s������m�K�%��q��=ݞ'�:�����̻
z(-����âsAuZ����{tq�/c5�Pn
#ψ^�nr��w��0{޴�Ӷ{=i$��N��W]��\GW����,��v���7W;tx�`l�s�cJY��0+�R�V��D�-p~zh��%����q�lW�+ ��� X"��!��T�{�ݏ+:���<݈�p�.�{x��]p?��K �/�Mی�ۥd���o�a�E�e�ጛ�+o:u�ϑ�%����{��#g����Y��wv�+�q(�i>��X���ӗ&�ޡ4&7\+����$<dw$�;=�v�I��p(J
���\��h��F�]%\4ާ{�I,�"s�eT�}	�-X��N!�=Yk=Y �3��9�Oz��z��؛Ż++n��.���{y��A�U憳[l�{��}wJ�ՎY�x��v�t��� x9�s^I�j&q�����^EQ��q}ǅ�e�l�%^�&rP�e��k@]N��n�N��V���������}S=��'o.P�hp����"7:��2����i^��Hlz*p]�lVUx��Zq��)�<��5�/np�*�v,���_��R�te֜6+j
8����F��m��H''���󗢨�r�$#S��~����G�mE��C����&����t��ɞKw�&�R
]ЍE��j�,v�O.�����ٛ]�t��	�IT
qL�~==�ɧf�tͦ�x���I6$2�+T n_[ق�]c�fsz�{�g��w�(�}!s���#Z|�����GcTY��CD��B|���t>�j�ч�u4ҽ�4Zσ�.�Zh���2[,�
��no+|-z�K���[�:�
�Y���(rW�/�յ�N4�֭��k�(@� ����K3�>����C˅^�82��V<5��Kn���dB�e��x�P�=q�q��]ݻ����̫
\S�
�hj{e+�7M��}����=�cO�)���i`g$�ڎM���(�'׭{Q�S��z�ξ��7Q՘1�
�X��$V:��}m�֞H4�>h*kێ��ͻ���ެ��֖�Xq��)�S=�S�!;y��M'���Tpݺ�x�VҜ#�X�i��i�!
��D`��E�y�}	�E��R1k.�㌪���d,_��M�=X����z���YTr�;(pw��$'#0���v9�w���9���A��F�7�wE�G)
����uV�\���^�
t��ݕ_/�l����臣f�f[����˗cC����D���,�ܑ���B#i�Ә�A
w�k�TV�䨪,���J.�(^�H:)�r
]��A�5�TW�A��� �q�ͱ)�y��ާ{A�αi7��fD�=��u��A�V�Cl�;7�tcv������N�}��^�{�x��3�M��^����M��3�E�����Ѕ|�OkU�3^氊7@ob��ײ|�b��^�8վ�9F��,�u=͹o7N��~��3�u� g^�iR[�8�[[<�ގ�J:+Ƨ�l�{;�F07F�H��w)�_dj,�� 9�NF�g.�Z�v睜���X\�jJ���^/�����#8�wJvA������̸L.w��7���E������{���g)by9��S셈��Pp����H��Kl�P3� u��]p�%Y6zN�f���]J�m�ϡ�KvRl�պ�;��8�y6�H�ۊn�>�>S�ڹ}�ӭ�)��by̆��2cuf'���u*�Xl��H#ԔS�A�D��o�����V<�]h�L CL��X���mߡՇGJ�#!�U��P� �.��3��l�K]�8�'z����н�8V՚p�!|�e8(w%ԩZӀ�y��j1}��x�ՙi��dp��! P̵�z��*�&���=�����`���ޏ���j�>U~�@ѵ�C���\��]͗����R������䩵��ч`����:G�%���7]kM�B:^�ێ���Ӓ1��`��^��ׂ&��z�*ۚ:f����B�ތUB�b�>By�b"p<
wxPi�j�hESCX�/���aw[��9uä{s54&�fʪc��alpy�N�Ll��P�O����}cn���b�G����~k�IX��6�V�,k�ּ94@j↸�NM,웼Z�k������ʣ��ž���{�y};ɟB�A��mdZ���=V�76���Z oA�v��nv�B�x� �*�n���eL���ˏ��qY�J���@�u�.{��؂u��Bd���F�%�ԋ\��ǋ���N%��z��Xd��6�z�PS=��]	��Gdu��g؋#����R���5#Gոj���[Ϋ��]�{�h�b����"��Ɋ�"޹m?P��n�e�ۣ��شGc0��w;���r���O�|l��%*ЩbU��	egI����4<���[�:�|���^2�`��G6�}H_G����H9�oz𰷪i	ۖ�4}��|�}��p��u�q���KQѡl�"�t[����
T�#�ù�dOX�͟Yz�� -��8�w&�2��Y�S�n�8!�w>�����Ϝ프��F�Ym�;�S��V����'����u3�{��/�L�+�Rp�Z��$��&Ջh�1�܇Y2�c26�Fufj���:���`��H"��^�Cm�rqMow�)쇲ɩ�+wCLKKh+al�ڎa�|D&�
�5�D�Z�Õy�tZ��quI��oN,詼�Lf�#D��=	�>j,Mx4*��,�ۺp47�.-qĎ����6��g�і�m�pr;�ŵ;۔5�B;�P[o�������^x�����.�#%��ob+��I6���Fu�qK�4\���{].��zT����5�(���0��1k.ܞmL�}�����ԥ��M�: ��13�y�$����v�4�V�y�_�air췣��R�]��6�__m�c%�3�I�D>���~�����w�u�]f"��1�py(n�ސ�*E2��;8`s���uw�a�nvk;��uz���ivl�ܫ�s���7ɯ���^���*�u�E��[m�J��W�J���N��P�Y��C�<����z(+M���Zpح�=��B��������t�J����PH*b�:,~�����za�=y�zi�m�{!`��c\F��m'K�9�ˢ�D#Ȉ|�����e�{CG�����=<9����[X�io�	f�2qT��y��F�KL������
�U��X�΍vuSo���5�M�5#3\M�K�{
��7u�'yW�.(=����C�|'���BΧ�Fϳ�R�˳[9��\���(N�-{Ti��N��:M�w��i��fn�l��yfe1X�������ӹ��9y�n8d�f�Yfv���;�F������)��l��h�vO�p+޽�*��	�yae�D������ ��#2�Hxd.ȍRq���SJ�n�����Z�6�<�	]��^��w';:F�3�\�Qb�J�8�Dݒq-Ë�:aՌ�ָ3���Ĕ���7�6+��2;�T���얥�wT���b}��.��f��T2N�����H��[ p��Bw{Ry��?OzlO}�~(���D��%?�5�tR�,��oF���b3�N_�G�yy�����E�}�*�ȉ��&��w^-�9Hc�V���8�>yx�/Fg>�T|ލ�!���!��s�^�ݫ��#8�����n�<z�IŻ(���,3��w�NM4c<�Ţ����*�L�뚢qt'�n��d]p��n��AN����B�W'{S��j�k���ե�vl�>���u=^3����3��f��-N<�����^e��ܚ*��=�e5|U=�*!X�ЬsFJ�h:|)Iw��=����{�s7ܳ3��Y;a%�.*�"��=b��(&FWm�h�ެ��Ek�Ư&����j��9�G�b���C����ʰ{�T��v�K{)�Ǯ#�Y����t�׺L����7��>C�c,?�67-Ժ>h:�<v1��<��t_��	�A�N��WT�n=�"��D芅Ni�WP�%]s���8AYA����t���l���C;N�m�1,�+	�\1�D�ǯ�t������Ҋ4�N�ٗaH��44-�,�숫vx�{E���oN]����`�[��8�y6�H�6����`)sǍ��u������[W�1�̤����u{�O$\:��Q7�{ͽW[�07��x$l�Cl�H�GmT�n���!9D��X���4�f��n�W8������V���`��V=צ��wo��f���~�AF��E��nh	CY5��U�nh2����̼�OWuMv�+D Ƈ#y�	1mA��@45���tn��a�S&_=7�Q�u�)��Oe:)1�|ъ�U����I揯6T\��S^՟ �;�gk�Sy���M�"�2��^/7�獶m������?j�ݷ���Q���=�[�LC��
�Ydp���N��y�W�G�%:�ǖ��dW��w�}��Z�B�d܈\�h��'�!aY[����򁛑p͙s�jݢF>�n��&~9�J�\�_��s��s�b�2���⊧x�OH� u�5��Y�}}yv⼺鯀�Q@r�>���7��G�;^-
����9T��Pc��u�A�Z�/�yf�Kc�y�AX�-���=���of�e���]�Z�\��Y(wN�ܑ
q����z�p����7:���g��aU4�ʛ�:^.]���ӌj�S��z1.!��Þ�V��l*
F��v�n������������;b��^�}�k��]�G}m���Sѐﯮ�̚��<yv*�u��Vn��F�:,�]����l�W㍕�C�GN����'�s�c���C�Y���s��^�θa��V�{�4hz�1ԡ�g��<�ܲ���X�fD��V���}������v�t��>�;n8����Fk9��F����i�I��(*�t.N)Q�u�{*!�:����v��Ua�{j�<�	���i��JϢk-O��+���
�n;�.H���Q�zФ3�#����rL��<T��P��
�l	��Cc�r�Ԅ ��;˲�\_��L�3F��4�v�V�{���rL$���hf�qn=�A��,˃���1��Tq^݁�
�o������Ctw	�7Բ�i3�=r�\��x8���=�W֮G]h:�yB:\�+t�8Kwvk���[�."=�F���$k�_E۴�-�Y�=�8V�Mz�W�����yާf�Zi��=�)S\��օ,�S�D�:\�uzl�-.�Fv�
��!H�'^�>�Wqs�h�=�����!����()�x�tv3_���Ъ����x�8�oo]6���^[��ݨ�Wq���J���"7�
�Eo!E��APڈR�%�b�L�[uhI���s����v��V�����6`�F�E��}�c�e�|�Q˥J���߷b���?%n��M?@��\/���iT����i�3f��� t�i�h����m��NB5K�F�!�F��/��č)i݀6Ȕ�v�`�k*���Fn����e��z�T}3(D�]�(��\���F�V�=M�������*� ٖ�t�����eVs�X�9�����S�A�5���Y$�岻˝}�jTI�9a��ZلK�^qu�Rmy���2��ٹV8�i��ȍ���!��N-]Ќ����xnl샨ge����ѝ�+�xP�d�ײ**�ϔ�|�7K���c�x�����i��J={��qه�J:��W#�Ɇ־�ӯܗ<ћ��Ap�.��B��=ن��iۥ��}�h�^mя6���]L<�N��'66�v�ٴ�T]���;5�y	�"-�G|�1xS��.3�yא�z��:��Wq���� ��[�/�c�qc��d�ZT1-�e�ѹf�|$]�̉;���+�A�h��DO�"�rm��yVE�6�9R�t�ԵɋE�b+6�N��՚�Z�(���7����7��o����3���sn�\�*���9G~S���<��L��}��τ��L�K�q�yKs*> n�5SB�ѱz�!ӝޒ���y$�^EAW6�ӻ�g^����c6VD�2��%��]����(#�:�t>����&Գ��\3��`�E֕#�z=MU��tG>j�]^��ͥ6:𶢰oJ�4Z���}z�k��q��_m+"f7�� o���1��l�*�=#���{�ݐ#�9�����ۑ����V����<Lop��b���6mج:�a gt9��ː«ucs�9ťmȺ'v0�8�✢,����nM�Ԃ���\���7Qr�go�$�Xoj2�/�H�*���r�-�[0�ஞ=2{ݪ!`��� ���������A[K;���U�=�2Ď��v����1��m�Vf��;]��z��UPD���Ĵ�l�VE
�#(�e�U�E��[Z�T��-H��YF�"���E���R��
"��.U*��R�[U�Ҷ��TJ��[Z-�5+��K)b�D�kB�bZU�kj�TQ��̵�Dm(�E&%LHQ�m�ՙLE�+E+Jт5�VҶ+*Km@�*%J�R��F5�
%S0��EQ҈��8�L�Q�k��R�h�j(TVҋ��.TE�
�ƶ*Җ���b[Rԣjh�kh�meJ�Q��5A
��T��Q�TF�eB�"(�ѭ\j)��j� ֖"�j�Ķж���(R��*�-D��Y-���k"��Q�e�V�eJ0Y-�%T��V��
X�� ����b!��Ԩ-q�\�h��A� �+�7z�2��:�����g���z�д����p������,J%�o3^vN۶�u]��
a��N���9vu�]X�1��6tg�;GZ!�;�#	�j���u�J��D|��y�����RҶ�c��U�ze�����1��6#GgI�S^�̕o<%^��S��6�}�m����.�����t��ګ�Z{\2�b9f��٤�`�6����t��P�7Ha^��[���Q��s6>槬#���h���n>��/�������͊���
ӯ7ڳ��zNǯ�Ρ�jl2���n�g��"
��i��{;��}��ס\��S��@�\�E�b�~�C^����\�����/d]%-.d���hc\F��m�u�ƫ�P�ha��ΐ?'��֋r�E��C�!W`���<9����V�'ׂVs�ݎ�� ý�C��wF������ka68-�}*���gU6�V�A�Fɝ=�㭰{���	�Q!��Sz���K�׸Q���\�ą�3��\_Z���~YQ���{��qJG٢�!j�j�u1���fkq��[�r��jo����$ɯht��܇��ޯ>ܑ�
��$�� [�GS*�Wm]�uPp-;BsSV���/���q�����59�|���U��w`�׹��c�@�,�.�Z�u��g$�j�PiBpZ��;j���39����R䰭�N34�5�����7�8-;�+��9����1���-���62���4pe,^��O4D'`���^'p��5�'p�L]vZ�QyE}C݁o%��[#���a	�3y�c�f5l�L6�M��o=�5��L����\Q��AeQ�l적s;��Vq���KŢ�kAj|�\�6�N�96I��oFiG\bG�f�/�V��ΖӢѳE����<����H�}�� �п[1��׍�������p�f�^<���n�+k�x<���˔PV�ў���̝��|�e�L�أ���Γ������]������Q��\���.��b�U��[QQW���U�D\�"��	d(F�{�[��1P�07w���`�h�����
ƶ��׊V�S\��U�׍����}�:;���T������m�ۡ�!x��j��8jB�zy���9��bQ�R{dqK�ѧA���seU��tg(�4�8:�h��
q��Ĵ�1äu*�Z���J�9֔����:����W)�_gxz���,٤�}��D���0�Ǔ�Ҋ��r!W`3�(���t;=���Z��3X�#9Gջ��#�b�C�t8%=y*�����OsR���8����%i���q�؝��l˵!d�44,gw�A�;|�x������]=\w[��\��;���Cn!�޷T[�cw��4vO{��j�O�y�+��3#wJ����}~l�O*9}g*� �Yޭy�k��JC�yt*���$��D6������>�Du��ʨ���n�7M�p�#u\�)8�AW�;��?<Ou׏?�f=(��؟^����"s�ɜ�&F5&���b'
�W��&%5(:(E�8��ENE���S6�!æa>5���\ǭ���� N��H�O)�[qJ/8u-�+�TQ����}���0�[�3�[�jŅt��ݙ���2�Z���	�[{;�p�G�Љ�]+�R��%Q���y�����=8��ՅsyӧS%��0�Qbh�U����>̀xOrp��x.�y����"����U��}�Oe:)1�CF+\EY��%���\|A(�o���Y�Nw��������MXhnw^�r^���̶����cnj4fٜ���,�B�o���iԡb����}O1;�K���+4D��A�VϽ� ~�[�㎋B�j���ȿj
�)�Иor����t��o#x<�V�*����c+��=\��d��n_Y�~�YN�$��x�Ol�q���:��Xd����*�zh�g��X3�o��%H>[�qg���;{%(����8vvӨFÛ��I���>.�o��UpV����<X�����Gc㡷��qf�ﰝƭ�;���cP�]:,�OX�u+���6|����nxv�g黝���ME��A�ʞ;pJE�����9�|�^�6qo�M��hf���PUg+���5N�R�J܈3�σ���{����F�2�N܇-�#>�y�	�������q�=cr����a��೹{l�>����4���\m-�z��98�=��ֽ���MW�s��۰wJÍ��$��Go{i��s��� ZfA�%	�+ظH3����v!EDUln"xsNb��?�]�v�y����i��NJ
���B�]��؍�#c����KIa�,�24mP����	�������C\�7�D���OUmŵ�]�=�������')պ\=�]ps��0���u�ۮ�h��:����ӣ���[o^W�۠]*�ov���9�T�a̬��[��;������B*�Ch9�Ş�˵yt�B,��s$���$���������uטS�@�<���N�n��Qo�C��UL�[��ksw|�����w[<����٢	��=h*�~����P#�t����t��c4:�k��rǚ��כ���b�1p�)
f�Hج�ӽ9�r9J��;�����:S�*�C�+�b�`���.�C^�2i��}*\����\oX����y�@�;O�i�y�i��[���O�RbG�6��4,t���a�R�u^wDZ|Ƿ�:5wBU�כ�X�,���+�vb��)�w�������j��˫��� �L\�r���9�� U�/7�-)��à���i=���x�����Y	��Kyv��K	fu�g>��vs�S�rQC�����OX���(&�i\u��{g�ְbFd��SH�z���]/%��ձȺU��4l�Sd#Jd�ӄD�F�j�x����VF��ܖٗ`)qO`*��C�@�]YTioD�QQEt���_b�I��J��u���1��H�m��Z��m륶�J�����g��[|.�o{W����uc}i�I@řj�if�xo�w)ν�,��v(\�D�&pe#��휞m؇V&�MU`ʜ�]��c���%�d
��Q�r/�')Xr��G	�ۆ�۬s/n�K^gi�㕃��bhsfױ5���ym��VKv5��ٝ����}�ّ���\Ȩek���@ +�Z�A\m��,�4saS�RB��..F��u9Z��j1�^iF�k��׫�UL�-��7��%MV�s{-X����(��y➸���ܴ���"<�zm���f�fE�_����swD��D�c��M1���4�EPhk�oj�v�^sҧ��M;�؛+6UVΆ0�t:[N�|6h��+\EPz6kηm�P��������}ݳ!�^��>M�V�������|��/4W�����~e�^���N|{����q�}f�eQ���Ha���~سz�Č��V�Жg���4���<��\pج�EΖ�Zf��E!�ja���}���ub�}*�{�Aؽ#�8]q�k}s�
��Wo{+��qYk�e%��U��Q{|���[j(;�T"��5pS�zgi���/Z}��x<V��>�Y�5�/��J�)��M��*��w^�.U������1���= ����58㏮Kl˵=�T����_,=N�\t��3��s��p�V��/U������� ZFD�1��r����fZ��@o7�jژ[BR�:���d�/xé݃$Ih-Wn-yύ��/8x?nv���Q�ITLj�M�ֻdu���[�1��;A�2�زĮv���ļJ5}�:�N�Lx|4]�u�w'�vt�d���P|���Y[Ѹ#���Zy~����g�
���$�|#�a���U�t%[������Z�G�����}�-��.�޿��m�M��R����ƅ6�����D�8��1��%8(*�GqȼT�8�)�64�aQ��J)���I��Q�,�����NJ�Me�x�$��g*	p��{��Z����f�G٧��B�����	�-E��4"����8:��w��/iD��0{B�x3��)Oe: $���PgTV���s��18ֻޜm�w���S�ϖ���}�^�-��X�]N�R�J��_nX�b�����]�vf�C{%��J���qP��΢�ƆjǪX7ƒ�v�uZ���Գqu����6/_
���7YH��h�26vMt�㪶��e(B�^G��y������^���q�uԣ��v�J^�T�l�O5�u�Y�=tiWe�K���a�0�Z���q6Zi��"��H:✡�M�i�S�~�-?d[�*��w�����g!ٗRn�fqC�!�6���F��.��D�/gsc�9'�h]�S:��[;6��rBs}+����T��+��QH�8�`S�=i�Ӱ������3=W�	n���aW�!`�o�W�Ĩ���'w���l��%�+�n�U��q���������uvDY}_7�������_��c�S��@���@��v�s�-���6v(v�M�|p�%X�l�Z� ���.O�^zoh9�`�E}�<�F�c�>�FS� #��A�2Q";Q^���۷9q:��u�9�]	�:��ꮤ'5�*$�81H
f+S[�e�m<�Ky��}�	|��e{�8�;��d��X#�:�q1H	�Sw��Iգ9����=X�\T{���u:�̑�6	�W�L��3�7�""/���s��N�YL^��ÍI�V7=Y�.��pw��J�`�Y��:9���*.e����ЪUFb��!����x�:��h��B�8�6*NH_���{��C�~�����볚��c�8;��K���%�h�A��o��WD��n�V�R�t���N�`�N��Ȯ�1w4��C�b��)QR��z}�s�g8;��M���b���Fu�ػ������J�z�{��Ѯ�?���y]��^���ɡ�bN��^i��c� ��5%�G���-ӂ���]C­�o�,J��P��_�ҕ�
�M�S�Ű241�r�
SP^h"b��>��cK�5�=���G�%s;���˺K�^f6I�{�u�r�X�< �����S7���]���Il�O�|(ԟ#ǲmR��DBR6/;��ŭ�N���>h9_''a7�/(Z�`}W�]���R�g"v����P�y8\�f��ײ��1��EBܚ��{����U�LٯD�o�ῷ�t����rԞmRJ6�NL���8� �-L]*�V�U9�b�����e7nз�H�x��wuWܷ/:y�r�/+M�?pߥ?A��]��0������S
[�6�U���K�'��%E�92t���3�/�tM-����R8\�TX"��!vف���j��_KO���`3'%���Ud���g*m�%�R\I�W�1
� a�D�T�{����jšF8������P����>�N�wySx���m�DP{��Vs _�Iq��}�+C�.�h9�^Y�
�>��C��v�����
�j����yw���x!��P��AN�ޓ;Quj���|�с��U3�(5��y,a��A���Lqx���Mi��:܏r�s���,&�g6�ֳ��c�t��z6�vWZy�h�Å	���$��m���؝��f-x���[����
�C:�H2��O<��+�"��!��r�V��ʵ�"��gr.u*�sÆ�%�=Y�w8���ׯ��S�h�G�<*�ܰoSٚx��X�V�Rʣ^�v����y�9|�ņ�_��j��!N�k2{�/M�bl��u1�k��#�j���
�a�ud���`V��΀&m:�\l�!a��q�9kXn̛nڥru.H���*��3�;f�R-9��o@�^QZ��Q�s1��gf�+0K�N�)!^L\/1M�J�=�>x z��F���f>��Q([ܖ�j)�������sO�3�d�~����c�N�Q�|��N�U83�3U�u��S�R���6���N
y�J����.�TԎ+����B/*���c��w�_?*1e�kr��c�b���1�Q|�˳�����)+�h���ݔ��L#�n�b��CpnlŨ�Sd�K��c.��)n�\��kpP?Y}Y�� ��۴�e�Q�CM��Mx����yЉ�wM��Ñٚq���.��9��ƥ��W������޽=ٍn^�Y��WN� /��w�GU}�=�"�c�^lY�M	�.��^W]h���,:���S�#�*&3����N_,�T0�P�Z� �0mHo�B�ůQy+_g*K�z�"kv�����R1�R}E��u�z��b��VV�{3�n�X����M�f�9\�83�Gu��D^,�i��|uܢ�]���1��K7.��NΈ�����7�˺\y[.�W7'ud��{Y�9rS�كXˍL$��Lu�U�	������/��Oj�۸�x����t*��[�ʏ��s�g�x_#{�f���N^���`��F��V������>`����R9@6��/h���)�`�u��!N�7g/����S�Qp훓.�E��I�⫆f�c�8���{�9�!_��t���V ۰�`����C�*0
wC*A��H�nN:�P��m�Sͽ[���e%׊�8������n��	���ߖ��Y��xS��uң<���*�:�$Y-^0%<K���o2����z����2�ݕ�dV��R�ֽ�{O�P�,�J��B��W6mDkc����N=�!�r��q�E�����-9F(��^����;��|�p66� �f�t���	�S즊��^1�[��>��:b��C��v͐��Z��7�R�.t
��{���a��S�a�O�hyn���{�)h;���ތ�t9��<�9�F�>�6�ԕ�Tڣ}��_.x"�I����eO=��@����>�mk%AXUh���UeJ������jT(�։E��Q���)+%-+V�-���ib�e�V�J��X��UکR��Q��FV�Eh��U"��Q�6��KZ�`����E�ֈ�5Z��iT�KV���[kKIZ���իIE���[kZ��V��,TJԭJ��X��,m���(��TQTb�,U��T���m�ڌmJYZVV�Q#Y`��h�UPEE������m�ZQX(���QF�V�R
����b�ն�Q���V*6�D�TT-����$eaPb��Qm��-��-�kU�j�£j�KE[e��Q��j���*�Z0��V1�[Z�TX��Q��)Q�keX)h%-��U�UE�J]��Z����ߗ�t�$����v�e.c�WM�3(�Q)z��갪��R�yށb/}�:��U�,�u`ʙW����o�{�%�)|uh������~>ӣ_.�C S��[d`�R�hDL�9z��u�u�v�lY0��,?��C��Bʇ��')���E#�!�w��f[��ؚ1��Pwg[C9(�;�� neX�`�8�@�)��_N�ʘɠu�F�$`�M���b��N@��=�ݝ��x�"1�!_��B�TUV��H��	E<��	gF:����U	�2<{U�*�ss�s���AN�@	���T���sb��"���0�J+a�0^Ot}���M�,lu_-a�Y���dR�0w28:����)�U�KA{)b5���*qT�fno��qn^���`�Na���l�٨�d�A�򭆔��<l�cݴs+f�#�$Rg���Vذ���3@iñ�����H�X�HF��o.ÛUÀ6�ଢ଼��S����`�{;���=4e��S4!^�2��p�d�+���HGX�QHަ C�9�%��3;�����r�#fG\�?$�T�Ԡ�L����^Z��}��}
��!���΋^k[�=�^�Ej��)��A�xkv��ȅ%7�H�V�3��w�r�'HrnfS��s�qVy��5x��u��>�x�(L�+�g�#5i-��ɤ�or�����S�һ�&w��A�b4����M�7J��4����uҚw�tA�p�ܳ��fm�W�k��+�ԩ��:��^�E��
³q莂4���!m�խ=Z���02�8��+���v�G7@�s�q\��E�)ql��	����H0�f�AZ���913�;J���u��s�PJW�\{���3HND�wJ��}�3N����2
�yJ�l�o@�Ex]P����U�Fƹw뭍#�Ņ~A܌�u{اM�(��W�-fm@�gR�+`S�TF���Z�JyԟU�յc�7`}~����QS4H�%����T��e�Y��7�B�\�J$����t�c&��x�:�|2b)�#7��]���K�J���87������=�x��W��J��9�F�x_"*�C�Զ'�֔�[�X�φPq�-�dT�1P�؂�Ȋ!�q"�"da��f�j�a'_y.ȣ�]s�{`�ƃ��L�]K�T<Uf��{�Y�C�@��ic��Q��4#����s�!�+o�fm�*鿬)1ؾk�����>� v��w?V��]���RgOd����Al�'���~ܬ���Z�2p�cXī�1S3���t��V��8�Ĝ�I�����(ʩ��b�֌n�9��;h�^N���zԓYdeD��U%��.�����C����>�c�T�-����O5K=8t��BՎ#A��Z�k{\�k�i�{K�5��b�}����vj���71i���+H�:�l����璠^�5�(=�	��
���)}�fbU#l׼`��P�gèRznbR���W�PT�l��cw��*##b���������N���1����6+�T*�{��F��{{x���#�A����C!ԅ8���7gb���W����l���7�Jݷ��s�g�8N:��d\1���#��C
^��]���s�p*��=i�EAx�,,Lqp+�o֣����^ͱ�n4L��;�J.<��e���JtbJ�t�@p6�t��]*���i��T�eX����� *��t�"��G�P�{>���5WGC�f93r�'�ִ���ƺ\��ܭ�S��������xB�J�ٺ�q��ɵ!E���o1>�SڦD1N<ܒ��V���L���sPm#t�<�Ll �Z06B���%P!O@�|o��m�f.,���M�� �����~'!�G\����7	Ɋ�D瓃��$�j��[ֱ�Y�&���D20PУ:kg'��a�Q�:���&�17Xm@�F��;ĔWV����$�~Y�Ut[��+/�Q�EzXovw�NC׭�l�L^�W�{���ΟO��˘�[;�
T�1W��0�6��k�p�+���{uv��M���缻�8�s\���ٳ�z�S����<o+Ɔ�>�n�1�:"���D�*LERFTU����^<����?�;ʣ�w�(����V�C�ޑ�#���Bg4�"*i��S���8�����j������6�e��C�~T�>.}k������7g
��ϥ]1lė�{ݖ[H���e�G���R/S���B
�9�^�]Y�nl�0���M����u<^-�����R��QF��Ɓ�13�9@FYp�q�x��'��z2�\�;{<��
�H�au\=T)�C�&+CO�<��iA�����gF�f_�LS���q.�WGz�� a�,AaD3������l�^� 6c'�9Z7��u��e�'�S7��9t��-+
/��)9)�AyC����ɭA�t]Y��A%��p�{��S���>�j���ǧ�V���1Ur��镳^�@�+Ë7a��-F�osW�|�r�봦�oJ�jB��'Ol�jb�Ls�C�f.�Zg/�;c֯#�d�������謻x��rϫDゑ 3(�8M��0[�uU�_K��r:�<�<��EWd��0K=Sï]�͇z�����W�$��fK�=���`�7�y�=:n�R���ų������OoIx��<ttD�,O"�M�8�S��_{��:���eh�J$��U{�Q����ȃl���Rܸ2�q�)1��v=r�<�G$�xPًI�W��O���}d�}]�e+�����*TX�8.`���.�--��+d0��@�d�׈���&v/9Sa�%ߔ�]��hi�T�5���ԏ��C�8!�^�)����ܳ�)�s�.,#vyK��]�T�����z"��N���A�t��n9�;��8��t�P�mh��=����ߏ��9_��2<�u�F|��ޤ���z��W��T=��d�p*�Ha�]St,��	Tm{�|>�����V�����f�n���s�9z ��ੰU8�i�lj�v�\�:ȣt
��\<	���������B�Y�}1�����xC���@��\]�@�8����t͜g㳢�s���3��n���!K����P� ��x�&ce�A3υL
m����a��=i{ѽ�ڪxli��Z�����ƽW!�\�}�aA��^>o�lѰՌ�NEFbO!k�&����һ�n���*5Ԧ�����%�=��:�S����6�<B��foj�Nf���	r&�r#z�ѕtޢ�Mwْ��q�9�=�vŕ�%|���cʸ`}ڒ�@lڜ�[rsy���
$M&/��Kt��|;���X�Q�O���s�mK1W�;a!�vP��h���X������ão.
�䥼J<�z+�%�y��Ю57ᙾ;EP'����4�m�i��;�!q��:vJ�P̅zyg�|ֽ�3F�o2�!^��FAr8�����&�E�ה���ř���ޕIp�<���v/�TN��ꕁ�Q1`��U|�J+l�V��8�lvR�w��9:]fɅ>ۘ�Oڈ�a;�tZ�U��ډ/P��e��IT��5�	�嗐C���CǇ�:mJ��;eL�j�Rî9��O��م.9w�J����"�vM�W����JP~(e��KER����-66TS�'��]�i���>�0Ct�i�����6�U�j�n�j]�#�W/��.�ӛ�2Q\.��{CX3��,�{�\I��k� ��M�%�����u8 �*u%���Rk���)�RU��V=�p�����g`Dթ�;{��;	���P��=*THN(4#�T�34/k�írĮn��+�y��k8��[w���<�����Q9_,FOW��s���-eLY!]��]u�	x���wD�kn��!�pX\q��sV]�4����/�vgnb8`=��@��_t۷yJ�3��55���$G�=�M�T�8�P����5NJ�Ļ���=qo=g�Bz�%��,4��Ś=
b8OtɃ����W�
�>�֓�κ�9+v%
y�c�F��#&*S�;���x�NlA����ո��l8��2ɱ���W~*L;��[׷�0��6b"�1J�c&�@��z�5�0�^0u�t��Mh#`��d[��Ryؕ~��½�>��-��N���E�Y��rݝ˝5�K�#�^h�u; ���E]��uM���0�i���W�9�D���>d�פ���Zp����{�k;CE.K0���H�� �Y� ^��{�E1��__'�f��b��+b�]�;	���6f�V��R�:��D���a�Hخ8{Yk���e����ք+��:5ʍ�sj��"�B�v61�;���
��c��N���z9�4� ���d�b���G@AK͠R]��S�qN*��=`'}	�+���r�tm=�:��e�K���=��T�-�-.}�r�ӐH�*N$�,e��ْ��\�e�=1�{)����x�kw����\z�A�n=����:e�f�Z"pH-ݜ3�a�垛G��Ft��x�Iy�Xþ�6Rȩ�u�dX�_$I�}t>��*&Ҭ���4�Ss�:�L��+r����ּ��N-���(�Oa'�ҋ�Ш�I��pUvf��A�(t;^���Utq�&+��fe�Y���̜ܻ���N��U_Fԋ
G@��("�+D����H���sc&ԅw2�I=�z���˄.ˆ�[�)�3\�w5�7J�:� ,с��ᓵh���o"/�.�O6��F�V�(9=)�\����#�}z�ʛ�'&(TI�pb�6�i�Ú_s��\a[�ގ�7i�؎�r/�6����2Eswў���t2$*LE��78����W=���g]���2�@������./��U`l�3'�l
��Bgh�3��%)S�=O���R��a� ����׭ ,*������U��U��"��sPx!xee�2��]�/8��:�����0T���= ��lۜ�Wh�
��0���Y�sc�&�9�b1���j1�q���E�iߺ����D8n{�pxj�	�]0ĵ��BIY��Ɇ"��P���9�!�&)��k���|c����o��o�͒�J�P�y�y���MȬ٤��q;�GN-`�*V*.x ��i�;��*bf�*���9M�^�xX�;�
��ttK���s)�����Ն�pS]�y�|.�E�[�����k��x_��&����%h�x�S 6�B<v���
;Z a�P�C>�~p���� ���Kf2}58ꬑ3Y�;��kE]K��l�k�θDj����Y����T�������^b�W^h�^�:�O�u�Q�L>F���t�+��0:Sڮ�Z�L?C�}��#��i���z�z�Ŕ�_����=���9
�e�b�b5:�hu9��+F�3�_��� k�oy)��1�w;v,�}�rֽ�r�C�}�*��#ׂ,WVDg�ʧs1:S[�vV<Z;[�H�Rz[��]��\�!�Qnq�;R�f:&���
�1 %#���,���rq]��,Z�P}�\��G�Y��^GEj�'��}�Ho�_�
+����]R?L�uK�ʖZUPV�Zlp��=�����k0�
��=%�*���h'4�E7��9r�u���n8"8Dl��D
r� �Th�8�����U�\�2)���6x�Q�h�8ڍm���f�!��YT#�d��:��~���YU�nlG�)1ː�k#;��r�fvV��ᩜ�o����d���{0xrƕ�%��!ʮ�ٜ�1>�ɸ.".\o�_$`�s+��&)C��/R�u�0�KK�Z�3�u��Sx�PU���z����gqxՋ��wb�5Y/����/aX�+��x>�%XE�V�λƇ6ӭ��m�h+�}��L��5 `3��ʧ��o����1�GYn�S�P��C)����#�Wk�����D��bćs�$	�e�)u<�y/�U3x{�¸4i��0)ƻ`�^i��tD�$�LEE����@��T��Χe�K,����,/��	
x���lR^4�#�k���\�~�3
m:�o�lѿ5c'{nM�Ⱥ:񋡓:����P=�],G�����f��1Ѓ���}ҍ�Bue�y���Ӿ�Yp-(z�T%��0��^35�p�e�>��[=2P�;M�B�fpJ�^�J�઱-�Q݈�kH�M3�O��p�mM�`�
�k�]!�BD(��W�]��n�Q� �̭:�(S!��5յ<�DعG#>s�,F@�xvu݇�aY��;՘~�Q��3��Y�'a���b�U���v�K�T(���Ah�ߵ��4��͓���Ùq�2������G���	�C����F!߳�$�	'���$���$��BH@�RB���$�܄��$��B���$��!$ I?�BH@��	!I��IN�$����$�!$ I?�	!I� IO�H@�rB����B����$��IO�����)����Ё�Y��8(���1#��ޒ�P�@�� �R�( �BA@}d$� D��(AT UHPP(B�PP ��"��Q"�!KL��J���*��*�T�U �JD�ѥJ���HT�J�I%T"���U J�4"EU(zeA!AT �HI�QT�H	("!E�)QTP�TR�RRU"J*B��$BUH *�*I"�^ƨ�P   yC-�����m�ݝ�n)��v��V�k�:�nb�uVtw��u��v]��`�uN�n�һ���n�F����v9��s]v��[�T��TUT�H�E�  gz�uثmܵwu��u7jj�g4�Uvwm�훊��Mv���:�nƭ�ݶn��9R��w�4�m1��]��YvXj����k���jR�DJ�B�H.�  ���;��`-��v��ݧiu�;U6�K�9l��ŝ�AwmXX�k��.�̹Gt�n����b�((�F���(��
(����QEQE���QEQ@8r�*"��(J���%�  6{� � ����:4QE ���QE��{&f�v�q�B��B�F�Kj��.��:鶶6����(6�X��h��U*��%UR�N�  n�孵�������hܔ˵���T.��e���MЊ��
Ejf�0:��vu4�tn��;���l��u�TJP�  l�=���[�ilrֻ��$J������w5����6ӝ#�b�����C��Z��[��1��u�W�Ԫ*T��QU�P�x  6���ۣF�ۭ�q�in�;��������v8n�vs��+7w]��\�iګ[��08:�wm��;��G.��й��m�m�7v����Rmm�qĩH�"�I��I
�  ju=�ݝmwb�Z�)ݫk�w*KFv����Z��vwg]�w-�۝m�:�svE]�:�̮m�h;i�&��5���V9\��í]����v�Р�IEI*RREU<  ��R�kwuN��0��ꢻ[��5�eJ�j��6ݶ�;�4���.�C-�t�nA��]�n���8���ڵҹ���f��m��-��n�����T*�������   �WM�Wcws��]v�m�Sm��n��w;ml�ٛa��]���v!�lݚΝnj�U�T���n�n�v��s���[�u�Ww!��ݫmv7�6��)P  "�����  T�����  "��	JT   5O�0j�D ��I&�*�=I�FbY*���qZ�JP�	"��f�H(���M��{�=�^��_�	!I�����!$ I<$�BC��IO��$�؄��$I! ��������������<��l���33�v+���<��kA��[Z.3�.����Ȳ�n"��B��t��+���	i丒�;�X(f�5���1]!L�7�ׅ�R�pT����4)�
9�P�sdU*J膩-f�����?)*Ȗ�)��2���yc_0�$6-��X�����NRd���Ȇ[�Ӷ����2�	�wR�շ�8�� f�Р��2��u��6�M5j�a�B�[�X��U�U��]���	��I�z%�QM�P����$h�t
���s�;����K�0&\��me�U-���B�`iOsA�z� 鳑���oWO��Ջ n���At�]���sfi�p-��/�z��@��U�,
E�1��|�����L��hR�]<-L��s0f+n�'�7ӣ����3q���(�R�T����ɚ����V�x����qҥ�I��^1�z�Z�%�A�91�	,GP�(Z)i4��D��6��
f�f��R�|�ѻ������n��+ųa�� ̋3sJv�1U�����J0��8ҵHX%��Ҕܧ���4PU���`S ����[{�g�s�����U���qZ6�U�3��
�K���B�Xi]�<V!*��,������e]H���r�*ɍ�*��YҌ4�M��A��ם��2m�u���tn��4�]�x[(!�E�KL$)��J٭)�q}�֚����Uy+U5���nº4�6�M�	0(XO����r'x�Vۣ��2˔�^0o1�I��h��Mg@�A�R;�R߲��+h��̣�5S�5J
)��^h�nd�%,,k�ݚu��5���:�7zP�=b����p�6f�̫Y�����+3Lh�#Q�0���k���(���r�i���;����ܖ�LV�y""�̳lX�N;�6~�-�̼��l*��lf�/a� �[�!�q��cj�`xբq��+V{"��c�]���ᴲ��λ��(�p��!��B�
�t�uݼ6�$�(�Ib�p閯r�X�fCg6-`/�Um�-U�:"��T�4�Ouau���ʘ�b�ȵ\i�P�4�u)��5v�L;�r�<8l��h�y���i:#8�#3Q��tE��x���jao̻ir ���Y�^��Y��J⬳/~�����Ci5�M#��1�AT�9�ȑeb�h�+hh.Q�j���aĦ���H�v ��1Pm	Y��jة�ԽsNdWW7�cP���.��t�'�O�=�F�N�>䆼d[௶��c�A8���9V����-u6�V���i:e�j���W����թ$�^�Pޅ�3VX��L��p��^nW�	KT�)*ڬDU��������V֦�آS����X�i��k^�Y�@�*���*�(��*«W"8,21�M�e�틠3Uܘ�=�wJ��Ł��ڟ&M���^d���H{����t2Q��,�1ٽʛL���	z��&��0�x�x-���n�`eΫ���yK�un�0�V2�^�N�Y�Ū�#�x�5D"�YI��V�KA���eg!��|��+am�l��wZ
j��F����[V�m�fX��N�	#�ɓi^?���lw�����Ķ����(�B�!j��ѧ
�Ǜ	�H�ӋSK��|{.�b�Y�xK
j��i�b�����iRd�y������5>�h �0�۬��^*�X�5�'4 ���4B��)س�%�l��DA�g4
R�.�Bʩ���e�p��H�����2�m/��an�Q�=��wFpP��Y�O͇Mq�[�����x��h��XrZ��*U�	X�b J��sr����Y)�e%�dҔ�MMr�ȅCM�ʦ�w(� ��/�3"��b�l:Ү��z�c�R��Q��x�	��;����k2�a�͔������%�i�N�݈�j/Y�0��.�*�+,��B�ё�%c��à/T��j� 1�)<�JZ�T�n���d9��ll-�n;{qb-K�Rg
�L���T�tmhf��D\��"�,H��3)8�wo,�����n�mu��]�C+�j뻲�)k��Čt:al$T�[О*��:{*��(K��Au�E�Ю�eK9P�0H�w�e�����2�=x�;+r��\R�l�0	�i�/&	���'��up�7JȳW�a-�a���4��㬺����3Z-��v�Q}z.�5��!�qK�z�h��D\�9���t]]��c�}�`�x��&��Z��i�r��gp�1�EJf�7^�� 'Gz�@���iC]��=�-ƨ��+wE�2��ڙ4�Ǵ�Ⴆ�B�!�u��.��c �:�&��y��,�T�|r�$��'�uth�(m�`M�/v��F�o�;�� ��F��oy�Xf�uگ��i%ۍ�ۻ�=w��Jh!�-��V<�������ss	��)��7��+/�7XB�V�k��V\7�u��.�*2�4ʣ�Y�Lr刃��uh0�hPӖ����]J�1Y(Z�i�8��&֮��2��H4ik�a	i(Z�,�C è
��I�ٽ̲:��U���<�F�1�j�(h]�k�j��i(���9�VV{v�F۰&�U�U��w����n�MW�M�G��n���Ŷܲ��ZY���\�а��^�^������Ϣ�&�M�X�ou�Z���4 �w[��nV:46����8�����?VmeE5���h%��`�v��(n�5J�]��+2����f1���S-�f�+�[N�I-��p�Z��WlP(�:���.���gV�ٮm�c)�e�׊��P?f�gRWYxZ����m 1�F�Gfc�l�#+T�����v�)�1q�h�[��^��[5&�45v,!��/�� 
��.�w���Xݠmm+]�0� )�o'J�z�6����i4�f�>�O�e1�x3[�M:��L��lHE�ԙ�P��x*�`�� 
԰*;w�oĢ=]a��@���W���0�Zְ\ cC;��cm
� ����,���ǴG<;{O��
d�z���d, ��kp�a��vU�Du�7Y�]]c��#lU�3�J��Ww�6��WQ+��tm���mC�f�`�:�-�PX��(��ȾV�+�a�v2̧u�C�+6�����XK"��O��(aZ�4�K�"�U&��]��!݁�ǯ!�JUK%]��6�KܫEn���lSr-�#�{�� joȵy�`vw%$��+ �pʎ��(P���4�q^L2���o)ݪ9�MF,�H�n���vù���Y�t��b�h<VYj������\t��p�Jd�ُ$
�YZ�p��	�Z���H���WWB��˼�V�2 ^Mܴ�[��a��TW���7XlVܠ��m��LڱoH�܋&�!��OHLL�XF^|��*PMw2���2�V|�JkV�i�{�ã~��v@/+�.�C�U���s�󤍗�8�FY�ڐCJ+�w�@�M\]��o��:�n�e�{��!�yݷ�ا ���4b�>���n�m:a0��El'P�	���f�+T�0#Z�X!3XY.���Bd�l l�gRjѴ]��3��Y\��]�0���4
;\���o]Yx|6��dcF�^D7+`Sݖ%��%�T���*8-ݬ���_��F
k��Z��\;���VQ�ۤX']�h�:*����gBWA��|-��/���������x�M "�]e��Ӣi�������Y������gr��mB"�.b(�)$k�c�yyf�kut��n��g7iH�Le�e�P8j M�p
���n��2�^Ů���2A�;Q���H���E�8 7�j�T��;9�6�T�rEr�z�aG+ J��)���6Xw�mnV�@N0�й�ށ�s%K/�w� �д�C`��YHh��ޗ`�B�m�rΏ�J�� ��x�aZ��Y������n]�fU��k�*��Ү�e�- :8i��6�a�;C�����w�� �
�&F6��j�(mލeKf��@�w6L��) ��I]�Vsu,q�4���Ee��o35ne$dI)g4��U�*m|�M�Y$Q֩6\��j��Ɣ݄��2���1D}J�c�-��Fƫ��*�݆�N�����|��,׏v���P�SB��jW��+��W;g�"��o��9r/��s��&��f���`�JE.�H]ؼ�ZFl4�ơ'/l��
�f�S�NݮR�6��À<xh�Yv[u��睍^^�1I��d��lv7cn���ŃB��0���X�B�,��i"�%��=gI�q�6���z�����Q�q=݆iߘ�e��'2�c����^�B���5>�E��`�m�z���%�
t�Z-ܵ�L�ݳ3�`��Wk�uohF'��|	G.�2��8f�����幋4��Y���M��z�
�{J��Q�g/2��orܽ|��<�u�t��
��'Y���2�tl�nYp��j��&�hQ5	
78�a����KE�
9[���#B:v. v���vV"������g���&e'ofH��oe�.�� ��F))]\�@�߮=��Ju�Y�T̳�B6<��i6N��kTT���%�y���hŘ�.efbX�]�x����^8͵��y>D2�Kf�H�r�*Yv�ȵ3,�"�q�wq�Xt)��,��2�/u�������4�Y���쳗��f�F���s���.�l�H������9�lSv�Z�ζ0�"�e�5�c[W�%�4�]:yt�M�E2��������۸@�;
�����h"5�NV� �ϖr��G�v+{H㥘e��/�j�8�%�7�2��gE�&��Ԣa�K��-9�7m�{T隽�Q��h���CJߕЅL�+YVoriR�nb�>sm��ٟA
KVX�74����!���x���BK�� W�Z6l]�u��t�Sn�XYӨv�ж��i=�ؒ�k/��gA��z(�N���앒���fBV��L���x�)[��ǣr���9��сc�)�$%yt,^QV��ҕbH�HK�3@-#bhXY�M!6�V�u�%Y����{x7G0&�xce�E�Yً�ai�� ���ȕ�tVS�l��w��I4n�*�T�i���Lڔ&-����K�nP�����E'�V �}�NdU���Mؒ�3c�������c[�ho$�z1kD��̼T$��-U�bA��e�V"��vU�U�7�Nk9�=*��kJ�fV�)�iU�@KK@]�[�&�H����R��ƃ��:�ʛX��ʴ L�k(����v^�s7�t^!��V((;A�J^����ufe]ܫv�mP�q����)�`g�ݼ�ӗ��oLZ.���CN��Z��8#�YҥJ��*�ٷ`�j��E�R��7h"�,|ɶNݽ�/U��l���u3�Y>�*�X�OY�TY4���n�� ZݲV��]�Ա'D�6��,_7xjD��f�C��o�mR�����O]�Jҥ���Gcx!'Gm�u76��eی��^i�rӧ�񭺟$H���$�ی�cl"t�\��W��jc�ǵ�n�-�U䱀8!-2/+(�� ��]�g�9���@<ëyS��vh9C,H.��u�VHPBά�r�Y���G���gQy�jV-��)���N\���{D��3 ��-��3�v.ᕢ�V<��g0�)GӫO]ɸ)+�to��c-��j�ִ�����LTc�GB͵)��6k���՜�q���B�4���U��:Kh���Ytwv��4�Q�ƭKkMʉ�I���7-٧���Gv��18��R,2�+�Uy<����l؋e��!�
X]m�[f��,d��th+]�'JI�^<P]ҡ[P�=�+(1�Y�o�K����uS��^e�Z����	�wN�ww�2I��&2�M�P�h�N��}�-\2�oӃ@�i�ڵ�e��L�{�Z#�WO6�fd�n	�6�N�(^��3�e`)7
v�~!�cz��XG��kN*�%���R�-]� �w�2��)j�\�˱�f��u�7H�YEՉ&�s4�0c�[i�N̛k�Uk����e�g�q�YN���M�B�(��9
e���%iq�8̨~&<�헻�u�G-X7u�U�>�P
��ƕ��I��uh�7/t��x	�VGW�h����a���aX�͌�@�Rwٗ���E�������������;�(����T�&+f�u�	w�0�J��=�����O������s�  2���۪�q!�w0?��,�L�X`�!;nѤ]�&ѕ�:��ۡ�N�OS�ò������t���
m ����QPS�xf�ƌӐW�J�<�*C(2w0U��d�6!�kմ-R�
�`�xh�@�T������.���ً-�ɓN�QDsv ������hM�4�Zi�\��Y�6!t&+lcՐ������h�Hi�qHu��!A������nM�5����b+ �q��C@�;�bkH�z{U5����i���D49����;v@ɹm(�Z�c%�m�tT�v�.�B�EPUcS�r�)٭���B�ݻ[���N4�h�\���I4���X:�m��X����b�C�Ѽ�޲��e�<�_=NWb\�΄wm���8p��:���ň�gD��|�	�y��\������0�XZ���iZ5��rlg]�M�yN�ĕ�j
�D�yf�H �a�y������e+Qf*8ᱺ���� ̳EB�8�/3@�9��![P�#@O�w(� �fS�eSGr�p�F��3�IGt��'����+t�e7,���}�k��Ε�;b{�1�)a�\�Gs(�#�^����ފ���7� tS�۹���Ʃ���q���-�!JTz��9�Xx�V�z�9�Ca���6��;�W@b$QW��q��xd�ե���Q9����T1�8=̩��p9U�3.����%���yZU��%�j�J���mJǠ�8-����@lV�lEV1��蒥�3.���U�Kw�͐d��hZ��rn֚� �ఠ彬U˪h'u�!-gf;�Yʂ�d���u�G�*v��zJV���Q��>{i�\��,�1_V�����FKǗ�����q���R�y��4|���`�#�1)CR���R��'�v�:�:�\��K7tQ��C���7���W-ޱ5E�|�D��iE�Ǘ��啜I��2{p.+���6Z���p�Ϟ���SޤqFj0���k@xG:ޒ_`�1��-"��}�ʃtt����W5gg���Ҿr�ʲ���8�N*�l�*�aՂ�%�Z�^�{3��+�����R�}�R���h
PW�w�;����}��=(ހ���]����q�ElO���̳]��l�xA2Mۧ�l�ؐ��q�I,�t��R`�:�	���R����)pl�%}��VU��n�>��K+�:�n)
�1�H�|�u���Vu�/;f���U�/����@���b������fZ����(��+�56�M�4۶[9;����7�ݖ�­�P`�%��t��� cY��{�Sy�Iħ>�Gl��Kc�nP5�v#��8c7�0��vp�T�g�I�qԠ5Zj����4Cyk���xƚi�:*	i��ׁp��h����b0[�����MCh�u��"j����Ǥs�c34 [���8�R�!�[WO3D��vi�j���f�gZ-���
�Þ�B�yg;p��}���me=��l�v	�ս��%�h�;���gb���:��!QD�7N�S�?�[�$z�M�M]cA;q�*�pl�J7ِ[��Pm�F���qG��	�)[\��H����:���_���Qˑ�e�ؓ�f+I�z�]g%�^r�W&�c�Y㚂�m	�����δ����(l��)��_f��"u�Z��(��xEVr��۹0�Wm&7b̏��მ)�J�ʇIB5�W�z�Bģ�n�v迢Z�_Sj6�:\���Enp��x����0@[��W;�zC�f���f26�:zV��h���a��C���0�c��t��5�f��1O�d�}.�s��0k����>cFW��ufʰƍ�}řa�IN�fJ�WJ�oj�<�/�=�Lc���m���b�y����=2�;��+}s�(����m�KӺ�x�"ȣ�\�����)�:���ӹg�Q����[���;wGt��M��yҲ��Vۙ��m:8B���Փv���Q/�f�7@��3f��;��K��=��FT�&���WIT�S����Ɗ9����������9���Y_Mn�t�X�C��$̡w��OQp2e.��Bjp�����C���Ïj�--@��3b5+n�&���5���6���)�A����kz톶��dC]V+m��i��R����d���C������ف��E�鼕��n��TA�0�P�CR�v��x��V��ql��[9j���E՞�2�䜣�[H����a}�O���+m�|���t\9W���Y�ʳf�k3x*K8��n�=�R.y���&A�X'R�h��WF1��0�����)�޼���ت�Z[÷��4���A�դ�뾰!BQ���(�4gc�d�X�l�Ƶ.�Wy����m:������+kG&�;%*w�F��-���u{5_�b�ظ��+�ͷ�+�Á胶<:p�4��]yX�S��Ώѵ�y	�n���\�����
���1ΕaP@գ��z�ݏpK�GQ���j<�FKŐ)c�V�5�Ӳ��-7�sw��g��;siɚ��<�����n�%>ѓ^*Lmd����`��ʇy|N���6���b1�j��LRȸ��zȦk��f] �3�� ̻]hV�tP@������̖Or�nɛ\��$PF�@03� 8�.����`�\J�El�l�RM��K[�Ҕ9k�Z]k�;��;�u\��&.�X��O�l���`�h[�1m��x
��&_s�.R�ך«MdAIe[[>�l��ʃӭ�PnKS3����s���CJ��C�.�sC7��Բz2I��U�7��Q�b�s���դ�K�"▤�]���O�m�c�J_r�����,e���$����V��^gk`�����q��� ��.%X��B��7��f����LQշ�<���o1hw�s}�]����6������8�ɶ�Ϲ�ڀc��uf,؂D�[	�ם�.ef�q�y7@dKKNo�#w�C�����K��.��\�m
1ލ�~��\Oe��c��Qd㹫��p��1,؛qEb��J�\e�[Cd
��B.��9�}mfU�8 ��z���x�U�Hd:��2J�Ù(ǆj]j��T�B�έ "�����1���-���o������u�V�C7noҵ����y((6�����G�\��A����:$�$[hx����L�����1j��j=�2z��Z�wz0��Yg�[��B�_*v��ىڶ9p��:T�� 
��e{s�ѽ��eJ�@�� �����8W�p�4�87'��{�)r:��ș�@�F��*��EKx��6��ɹU�wF�ʕ�h��ojwV��.<F��f�s�]�V%JzA\3j�^��+V����s�DS�(����B�W]k'j3��&jT����m�
6ò��ګ�����/V�i�y��el�ʴ�ۤ�si�5����v�*��N����ko\�:�Q��'�?�� 5�_1QC1ma|u�y���z���-���`[��4��ηy�7�AL;|��;&M�j^u�a7�nl
drs8�ꗸ����
!�����u6�{�5��Xk�����w/�Q�\
Rg���se\��Xw�0�	�
�fA�5��f�[����ɛWP�h��!(`$��n�=Oxs�<�Sל6S��c��I�JF�*�n<r2��;t)���z���*�����K� 2�.���nr�7y�.��m	7k�\hWwa�eZX�ƛ��z	���G7w�ڗƷ Y�e�!��,�f�9�Ww"��B8�����hN��I$&�ݶ��؞N�K� L��������G���7��"
�s��B��6w�v K����:�̬c�^��!�Q\�W��ܔ�iBj}���ǓObk�w��4��Ψkt���W'`��+kA�Rə�]��P!��M��:��y��������2�q|�Z�yF�v��:<�Z����P�
�xćS{ze��W��}��Y]�
Z�fBK:�ߵd�a����\
�f��=�Yե�]Y��K���U���>s_9�U<
b�k�*@��м�h+����k���4���u��g)�X���D
@Z=ܕgv݉��ئ��4��oI�r4[�
���u:\�I����.�.ó�
�5�jISYK�MA૱��bh̐�-���'1m�)�[��S�w�p���;�%��q�E���s�
ӥ��y*���ފhn��3�n��W�\+�"SP�6/h���{�r�d�f�%�mǮ�$�!Yn�u:�@�#��-iaRSs�Ԫ�T��Zj�8�H��Y�3*�l铛[b��j���L|���K��Z��ۖ�)��kR���t(v����u��c�6��1>i�3Fڽ��
qN�6�����}`��u|�YSsn�Q�Uܝ��1e��TwO5� �����8فJ�H�M�9y���:|{Tr�S��ɴk.��N��N�u����obh�u��r�뒉����zul}֔T���GP|hS���B�J�h�+�\��޷�J�ب����za��n���μ�}Q���[E,���5KQ"��
T�4�8o��\�k�w�|�=0\8gn"�}��퍠x0��s�΅���_mB�bOC��Sd���-����SEEݣ��A��1^�_%��>.��L0j|9�:v]�Yq55ݑ��b��G��|����ӵ�rZ�Q��8՚93�Ԣ�W0��t4��u����g,"�S�e+6_.�m4֙N3n��ͻ�����Zc��,��޼��칥,{$
6E��n;���(������O	1q��S��gS�]�2�m+�0��F��h7sk&�*R�~[�`]�EpJ�E��Q$+�of4s��d|ﱔ]Ar��X�T�z�׌9�O^��Op}�U��QZ!z�}onɣ�.�pG�p���ąI��P˶��L����[�n��}�uˆ�4��]����hv�&~�����~eF�8��f�h�X��0l\�1)W<;j������W�u�u�*,�rV+ͻ��v�,q���&\�Vj���e�.뱥��ý���#\Us�|�r�!Ov�`��y����Et������ē���Yon�m�;��A�ִ�`��Dv���o4�x$ �g����B+oB�,���V��"l7Ema���;x&�#t4[�,��d�H����|
R9��j*�*��B�)v�R)^V8w'}l6�|,u*0�pOo>k�4s��뇭�Ѯ�#�N��cx�j����IU�0�_5WqTu�`~i��Ռq|P-l��q��v�ޗ	CJ�<�ҥ��7�ݼ���,��+^�kXp���[���k^�i�:���ėo:8'��hɔ;���*nWWXج�\z�&���m�`��c���ڹ"�u�n��=�Y�Q�[��l���_ x�(��MDxN\�u�r��m��|��������Ho!F�J��뮢e��������F�`��ݞ�Uy5WR�UL$�9��Z2�w"7Q��ܮ�Vݩ2�s�R��8{�v򚓡�u�L�ǜ�VWQ*_��Vˬ��)]��t%�!������"s���R�*�/"5���^Yh]
õ�s<U1�k�!�k��=�ɶ��N��:q�1��5)sV�N�%����Bhw�'��Ie��.�No����zim����Ffs�v��t�8�5(	�����ŋ�0��˳W3���M,n/���Ψ� ��Wٔ�ށQ�fs��/F�v�]%�5���F�V:(�>v�hy��c� E]���-���@h;&vdv����(N�w��]�p�����LK��%�W]�� ���\���mp8 ���a���`�H���ʣ]W؂;�d\;���89��ĺ���r�A��7��E��zhLvL��� ����XF�<�G�f�If��p�� �b���Y��U�^bS�N��7�^��fn�p��'��ͱ�ϡ�]6�"
[�6gIV���V9�<�r�s���c:���M��']���n��9.�2f��
�/3e�CV�dokSx(��9�,xr!�_)9
��+{Q��!ا�b�8rye9�$j-R���^s���:�.�G��eͥ.�][� #9�}�
�&h�2E��p�
%#�:�-�%.52�@��w�6��<�c�:�jNf`Cs��4���uǵ�+8o17�tS�P��먿�#��H�n.��Ɉ;(R��T�ڇG:�B�a,�%�c+5f%sD��Y�u�1\��h�q���R��<}�T���m>@�}+.�p�v�⭠O4�|B��n�OD�JF�O�hzx�4Mu��Ӭ��ʂ�m�w.ro�������A��Q���zfi\ΰub�օ�n[��i�R�ʂcY�U�]�����re�d>�['�0�fa���WM���D��Wh�W�<E�)Ý����l�v�F�*;ʅ�,���3\
D��� v��X��6��e0�<���Y�짻�],�����3�y]����}n�6��ݗ�j�˳[�yPC@P,�L�^=]�Z~2L�ʍ�lv��Y%B���ѷZ���P�	����FKV��A%`Hݞ�u	�rs2�m>\n�,�:��V��JT�*-E�F�Lr�w���tN��G�-S�P�>�)��^�X�ո2�wR�i��v��!�ڃZ6�H\����ܧk�g���+�O��ڱ:�H��v�����v��F,���@�e{��GP�t�t�o�1��_uѱ�͒���PNWJ�[�F�#}�dn�5&{�5����˴���i��C⫴���St�Mmw�+��1Ӂn��eAP�l����"-��7����
��t��sXu˧e��
����[G�͈���Ln+��g��v�+�s[��Jla�CF��bi�{zVV�˅Ԥ��볲�C}F�82n��=�|�'eq5)M�}֨}���ޑ�+��4M�N�G�
����S����-d��F	Xw(WNz+�DuA쫖fj
�mcm��o��
9����"�R+緎��ܛ-���+sj��c�Y}ٰA6r��J���{�30D;ZU��0hGS���� ��Xio^�JP�uo�N�f��1�Ћ�:�mB ˛M�wiNΘ�,�B��Kחyje+�K #�o��$�\v\ub�W��:��Y��5��zyj�}�. ��!�6��o.u�J���}jd�(��˥�c�Y"^��-U�MNr�-m����r��#$�|���/ou�l���M�_Uv�Vɻ�N���Ơ)	y�U�Q	�f�w�-F8�&7�[Ϡy+b�������)&4����I$�I$�ʱ7�qN��M�>��}�������I! ����IM�Ԝ���$j�~=RX�Ywd�P�ށ�9N�&�-d8��ŝ�����t�n �.�-" �m�u��˖n�z�֝8+p��.�06e�&����dGwD�b�zj�yZ;S]#hr�r�)]2%�ժ9��������O�u3�g5I���Ti����,���c�"�K�/��!��1<�m#z�y	��L��[,_dy�^똌rqxp������
��t^�_V��v���3�jc_݉M������x��]0��Vf��SZHh�^�)Kh���8L��ObwO� ۡ�4�WV��q���u�^f$�^��D�^	]GG 룳�6�6wku|I�r��U�̂���:�a��C���l�+�I���Ҿx.-�m�RV�A���a6t��֨�'+2�jy�̴�Y�bt��huu���g\�q�%*���ͬ�;��I�	������lZs+0i�:�i&���HWU�[��ųQү\�)�[y!����h9���cu����KB"�g���'�E��	��\��ibNP�ȹ.M��,t8zN���	Gl�9K�+��xV�m7��U��e��ֶj5h��.X%�熰TCmbӋ"Ϯ�(RF r�mf(�=K���qd��3�˖Q��c��RL(r���O����&[�.�L��]y4�wF�We@���:Q�Vh	��%z���dT��,��z��n�xћ��"kcv�@�%%�m��@>���Wɓ�i�#V�8��ӭ�����ޙ��I<���C�������\���"�S��u^�8V��ruۧ�ӆ���1@hB#4hxznU⸺�XX��*�s�n�	�-����`��������t���<!b�4�ewC�J�|��К]aeZI̥�Q��;c2�M&w^L�u���u6o,�8��&����F<��F�̮�5Y�����Z����nQVל"�h�ó�J�(�^�,$If]f ��qŰ�y]�A��q��Ѿ&���G���˛N@V
}��>��p��& sm��D�ђ��dE�	�9mU�Ac6�Y �	��x�����P�F)����K��ֲ�j�m��G�=qi㵸-n���z���º���*��S63� Ҿ��M��P��X2��6@�bJ�Z���g�ap�Iݩho��HR�\@n�ǚ�kNW4�.�)��(Tc��7:���!�ܻʕ4N��2w�l��ղ�x���\��/\쭲�Ho��U� U�|�n,�Z�+͠c����4�
���N�󫂮6�\u�+F �-	'U�Z���Ϻ.��{��F��+�wG2��g�����m�#4�GT���S5�:{4_J�Z�rM�5���2i�V����n���j�Ѓ�V�di�W������9�f���ȘiV�{�Ɩ�G�@�R^�Un�����1BN:��mF�R���\!a��Sgiv:Wr@��%wPЯ1&�a_E��r��9]����Bw9c�+
*&��*,���g�6]]����K�&�]JQ&*��{2�B���Th�Uzȗ/���p�&���IPRm�;�ɚ�Y��' q�]�-oLTr����.�I˗�R(�Ȍ}n�\��ߚ�7��jgs�����͎V0����N�L �nw=�&wi��lZ5��V����Ej-B�yu��U/����;Um#���Σ|PFSM-t�ӹP��w7�����
ת��`�D�=F���T9N�ֻܴ�ZZ�z��)`NpK6�"��]Ω�Mg�����,����܁��o�t��n��pn�m�*��\Kpp��gV`����5`�Lf� �\�����j��]\reuS�\�ۜ��K��P��������]t/�%a�M��t��ÀQ7Hء�x�\ ��IY����inǶh��b� t-ލy]34��y\�(ti�Ô�����ı��#���^*t^r��癕;Kg�e�+x�S�nQ�-�T!K���&�v���E��9/vR,��d�4
�m�މ��sc&e��6���(A�0C�I��v_`[2�m�9�K�86�;��33�EY]�Z�T38�͗
�
�wEm�Ҷ8��I8^-����?-\���f��1�;r�=ˮ"�I�qL捼��k�}/-��B8C�;3Sy	,��M�`̩}e<xu����Z�{������`o8�a��KlY�m�Ô�S`}bD�z�+N��gi�oTmX��pum%�,�W�+]se�E�Յ�(3M�w�^Չ���R��Vv�-D�Ұ��nf�ڢ�+��	��u�z5gq����zZ� ��"Z�r�GF��c��o��<��NQʛZ���T��ĻEW��%d�����Y�\�\��+�
a[�����: ��*����V��l+�j�9��|�)�f���]�m,;�l���f��a:{a�*�t��KpH�O�q�i���#�gj�*�T�E=� �M0ͺ�}�cU��ئl��X:��#���*�P{V:c{[uCuǸҬw�m]���9�b�t_!�fVς�;�9\��
���:�5&_Br녃5��e�}��.�_]�ky�wDEV梊hۨ�V>��m(f
KEM���ݲ�f�V��E�	�Cu�d�/t+V��JB�wlE�8��U�d��/�s�
��ɘ��գ2���5E��%�r�������\�> ��e�KIĢ�7�/.�$���K��*�ڊiz�ٳ�}(f�ջ������@u_j)��]L�s��k+k97Q�Bb���sT�X����7�i��e<zӺλja�Y�#먲�P�^Ѣ�}R��W9������T��`�K���MC��]B6r"��9��U�t	�Ön.ڹ���q)9�)�>�H�&�BF����|�"f���\w�]���fd�1Kݏ�L��/��,C�q��p�w_.'yVq��<B�T��o���]]�|�N�7Yb�x������g�����y�._�2���Z>t����+ �C���7���%����sn" T*P��Zn�~�	�H�uX��i�j�zJV�U,�<����7[�ٕ��7ٻ�a/�+kFQdF�wz^ D��1lmS�st��-�[��R�a;�ay�k��Rt���1�.Qή΋f�/OT#U�9�d����qf�˕������q��w�jL�2TF�<�볱
HZ"��fO�ʔ�]�I��U�Q �T�b�s6,c/�5ʶ&70�z�����wʥh�КsN��%픎$5�{�EN1m��Tei ���ӻ�����4z��F\��C/�
�0�>� �vS����얤�.�0�F��Tk�� ��GXy�D^�Ֆ:�q՗�:��ߝ�؝F4=���j�8��%���9sgnN�vet�I��1�2�����v���=Σe}�t�,n	�;jܦjP���2#Y�s���WƓX�Wΐ�r��]Coi��I�,ݻ�e9Q4֑f�X2*�:=դ/%�U�b�v�ƭ�y�wZ�֞�RZ���+���E)�fe��A����P�i�i���fB�r��w�0e5Wה�b�͇!t���'`�'5�[u��ꉞB��j��M�J�%[4,lA��ӕ�Gׂ��![�^pu�|B�V1vgD�j�s��u3˳x ��_�X����J.$��פ�(��к��Ft�.�%˖�Ý3@����S,-հ�9�_}�cKE�)չ{�Wf�$ՁR�����R��C9�kRT�Ԉ������h.X��ǴR�����/��vT�F��Evډ��;��dO*�����:��żyV:��ʺ�(�?V�N�ʻp\��E��I�P��C�Ι�����H�A�@���dtt��=2��6�U�ʰi�S��յ�s7�<�\l�☁���9�u�^p��Ct�		��_!�U�T~��giީB��1Z���-Z��T�%<��`[dݜo�)�v١G���q+���z=�;qiA�xrv��q���f4����@�R����c~��v� [���6�sR�X�JN��@�7�Y6bʺ7ҙ���~���y�˘.�e]�W|��Jm�;�hw�+֨k��(�k]�wnVN3���v�N1�5=`Ht����p^��d�CP�Is�տ	Y�dZi�7n��1�(<�`��:�;m�	��A�nI�խE%}����V���Ȳm�d�J��=ʉw�cX�@J�ݝ�I*�+���#�g/.�W��/��9+J9�`��*�[P�q��X2a�ȝ��d��m�(vF�4�o ��v1��6���Ƅ����g	y�{)-;ޱ��h�5/nq�D(�Q�5 (���ʝ�����-TM�8#I��P�hP'n+H_e��LʊT�{�dPT�vq{��U���ZU/nd6�$�-`�cM�4�@�͝T��aŲMm�F����l��
�׷ �
J����)1Z��!��{�����Nݪ�K],�F�S/�eAϝ�c+Yl�8oiǎ��$�|o!E�Z�:P._[�����i�5�#�l��-e@k.a�%�U[�u�P%�����n�>��0��1	/q��槖�I�ޥ;z�U�*��ghi�ܾ|��U ���,�IikM�-Ko���痛�!�J��
��mW,��`=A�٘٬��4a��E�ܴ}Q�����ꌅ��+VuʗӮ��u�v�ܷ2gt�R���uuغ-F�Q��v�^n�Mf���6K��[�cU�}ضu�6��t�*�&��K"^f�_})�-k�R���v8Z<IB�>Ȕ�-^���"e��+}�F��Wɡ���nލ��������w+�-��gt�Q��������F�b�3���:Q.����.��o��r�duDŬ[3�q���<y.�R�N�G%�/�e����$}�uw�D�n�U������ ���2�]t_R�������K9�0q:k������@Uk1vFq���N�Y`R��A�=[��
T6��,
��,V1���㵠��f�aD�7� ��X�lpbܥ-ji�!��[QR�3zqf���r:��:�2pq�r��)�a�H�����yC�J
%ـd4T��5M����b���^�sc�V���>��$ӵ)\ޤ _l�s���������P��:ԷE#g�Qp˫���;ծ�Ard��	N3X�����т������5}���tmݲ4���n�S<P���C�ó7t��2�:Vw��I����@*wJ�7�p]<���ŷhV�l�49b殞-}��u:�]er\�r�O�Y����{C*;�l�
v�1�3���:2��`�������ʃ2`�T��f<B��d4�X�z�n����AU���*J!:�q��gf7z����a��d^��ElY����Ӧ-�j��X��'qMMf�S[<m���ZW\�SR��y,�> �z�Z��G�DWS�����Nm%*�;�M"�9�c��ޤa��N��;~	�O��s�SGs�'�Zp�����u���b�L���6,"1+dP�!��e5i�.�d�8��-yk��8Q<�N��Z�n'�l��:��3f@Ȭ��$�V��X�R=����V��Ń��e	ڬ�a�d:z�2�^Xu`��]S��q��YM1�)q�
��$��y�N�6�[�0���eG�l�^�J�%̉,Y�F�8,-Du=	��7�H�V�!]��j�*��1����-ۙ;H��w�ST���F��BW9��on	-��Rٖ��Ӎ�`�5�b�P�m���ٙ�Oq�%wk��* {�>\�p�e)�id�2V��eS���s/i��6��Ҭ���}W�gR�{��i��%mh6���ث��oa��4Һ.5pZ��f�]oD���5Z�Z��M3���j"�c���C�ǼȮ�xZ���6���=��O��2�6a�s!��������j� <���ςQ���U>��w��
��<abp�{;+Y��fk�j.2I�!�e���\���6��}$*�'�Ź�!�X��i�Ҟ�V �j��"�a�dc��+Ejl����A��V+,5�r�8s]���T%bW�6�<��.�k�K����ڔ�B���B*.�i��o����U���RğѥG$Nۤ�y9���|�%�$�9ų]���^V��XJY(�{Yfa�a+�d��7���X�C%:����e\U�K3\B>=�ۋy��v��5,6ͱ�� �u��W��I���2^�m��gB��t=F��@Ȍ��.΋��-w�f�#U�"^�Q�A0_Rdc\xVTC̎�e���/�KE�#�s�GWJPX'�gb�0\�������Y3�t�6���I �Z�z��+g�ۭ�v���Hr�Gm�؜�s���������f���,�K�+*V�U���"��=�)9����'���
YtV�ws{�;-�HGOl���-��4���r��Ƨa�"v�g��
�qjxf�ꙏb�l�Q��Vin8��XާS-�f�0�����}�F&����o+�c�d[S�2:Y��:����p5�3h]Q7C)�m��d��Eݰ��E���e���W[�:�Tlg}�TP�,oX��WK8�Z��	�B�ΦuZ�n�]a=���e@z��D*h�̥qmJY&�L����@mN�=��{H�%畽9�]���V�P��ɇWqq[a�����iv�Q�ٹ\�s�|���K��Mֳ�`e�Ǻ+3�͒W)t]%�e�K�LRM�N�����:�'Ԩ]�[n��
������Qн]&���}�Xe�4)����f��պ��8#]�IK�yu6�Z���n�e��������{n0qᲈ�ջ\W����쯫��z#��ǝ��="��;c��*��P�'dj�ebr�k��oǸ*�s`f:޵�Բ6��c�L�թ����Z�QRl�[���p�2���n���1��tB�C���[��V�J�@oxN�4%na∩���Z��.�]ًB4V�^�8k��+X�7fQv�Xް��ivh���5uօу,ܢ��RX.m�����I�����÷a �0����9X尰3��[*� ��9�v��56R�)t_.ӊZ"����~.�|��w,,�M��zOB��o9��p;�j��@���������)��^����fc�}&Q޴�;�V(S�x,�N�_ni4����$(]+2����&ʺ9u%]gJ�j��h�z��\\���?�jj{­egvg#�ucf{O�͛_9[�ҵh,+稩�h<�[��:[��U�L�9�l�ԘU�]���2�������]�u�]�EZAt������y4�C2Ɣ���]��N���jJVVM�;wv4qMw�ns�]L��;q�vIٍ�%։��tzmte	�R[ܯ/�hָrWA��@�df:K�V���i�LcTl�s�wQ<Y��N���ݩ�bҸ�jU����3�b�mu�KT�PI`�;���ii���(�2nNpmN���!=������ru���E_p�؝�g]���站��Z����st��-��m��j(��[PQX��J�ikiF�*+]�2Vت"��Ab���%I���Z�%�U�[eDeJR�!V��������U(��-lm+-(1-��(�Ԭ��clX*��J%KkkF�iQEj�DU,PT�V��[UV҉l*��Ƶ�V-d�jV[`�TJ�26�̊�6�T-Z2�kkT�s*��F�q1UAE����pEX�Z�V�K���".1lE[B��b�ш�(U��(֩J�JԊ�TKj�6ʖ��QTQbD�q�,����ZV�`���0�JWWWR(�9T��5���B��X�UU�1��
�����m���[[*���V��[T����ʶ�`"5���+2�bѢ�ME\���ƣj5R���rʩ�j��PQV�X�Qb5�-����+%TEm(ZR�[E�AE�����J5cQV6��e�҈�d��ָ����Uj��"ƭ�Z#Lq��R�P-��"F[(�m�T[j��wWB��3�TK�����7�B���\!�����ly�sV"e����&�̗�×�oJ�κ��3Kc�d�κ�i�J�M��L;���fS����q���s���������+�ʮ��ј
#w���+[(�-��+�\N�j�
��*���T�E�,���޳/♆�6G�ج�9���]y݂W�ݸY�p���B�[��[���<T��Q�|�����* �e��O�Mô��-���1J}�,�,�����y;�jx�)�2m�q�����l�;Q�&�0����]�F���5b'q���<����aD����pJ����Cn1;sSx�c#�8��"���S��+J� e�:j'��"R�Q::j�o��^�0.Y�3�6�����}u�ލ�/&����>{�!�\����n����ȑ�<��Ҷ�����{�MNv������EVn�יm�ab\�˚��g��7L�ca�d@�9���<�9�o;.���ĳ6`�rR]{��s1��5߂/�RҊ�\v����rYI�sr&�i�d�]���=������^&�c�8���[-{���<�$
��k� ��u�&�d�Pr���r�����b���9W{z��R|Щ�^\#c��y�o�>���F��o34�@Kx�5{�hOub~9(ii.��Qr��Ǽ!fp�Mv�WG��m����H;z>����t�s����B�S��#�U�Zh����gL':���Л�1U��ER�]�U��P��\h��!r��sƮ������Z_<>l�FyB��Y����5!�*��W2c�]���eM�U=��5���be`շ���Vy7|�Y>y\��7��Y��:릩:�$,��<�o��T��ǰ)O�bw+�޲r�K�p7��4�X�\K����.^uf
�L�7ѪR��Q��>4߼�j�Kɽ��Y�s�1J13����W�ʌ;SeY��Z���:B�KG�r](W ��{k�洗rN3c���π{Ά����wr��-�\js�YQkIJ�^��r�{{=Xۡj��<�t�6r �q��u2�Ɣ)C�@s��R�{�?���U�ҸvDܤd�wn�7iƽ����Ӌ �~�Q3܌e1VÂj�BT�:�&�$+�ެ��i��v����¥�m��Z �2�؜^%�� ����gPTwa�T=�����b��o��,���'�����J��5u7�:J�k@oZ$��Li"M�7�ǝ�Ǒ5��L�d����Bg;=z��V=�GC��;��H���-�:|�J�,�;]�)U�����=��1��Y�ה�?(��v�Fً;L��d����(_TO�x�L��`]�Ƿ)�\5I}f�)l;&QIٮ?�K��AS����l��mF!���`S�֣F�צ�g��@j���� {*���TR�&M��`��#$��K���7z��v\�{|��]����(g�*Zi)Kٵ.S��F:�4��D���n��4V_�_�x���d+R��*��['Q�:�O1�wD�1Q�ɇ~n�� �>�v
Lv�8�a��Zh���q�C{(4	���k�],u�~'�aH�g/�U3�h��_#�һ}g�U۲8ɔ-�e1/�F�4�zA�=�d�c����E���kn�-5���[r�
շ�2��3!6fq�@�&5��3��v�ô�O!F��-/h�D�n{L7n����]��������y�����&ltB�������kDXwA�孳=�K�X���K%�C�xujs��q\U��}s�p�13������&��_��_&̲��F0�1b���0��/ �V=K9TԻ<�x@���k�:z�T!�heqcsQw��ۅ���:˱��Ҕ�d�t�݋�de&&zcX�P��}���]���E��v��ǳsVg�wp[��<)zX��Е�x�������[%v�k�|�ӌ��l�V\���D�I�p��q�ۊ�[��do�)]�W 
�ԣRU�D]B�C����_t���k�wx"ކc�����6�Ť�i^!7�m���ҸF`�L�lG�.%+�&\�u3��N`odV���1Їe�יH��O(ܶ3ΙSl&4������
���d~N����;P�&��Lud eQ�=��U�e�\�^W�>*^0������V�9 2�S1������*u�=/ݾ��.f�[2֬j���4��߶�u��ާ0}oL���ŭbQT�ɒ�<N�+�W~=h�uM��6&��V�џKU�Gܲ��G�m'zxV�rת=!x>ʨ�K�Uc2�b�i�d�ǣ���J. a�"Dw	��T���Z"��A.rgUk	Hs�;�5 ���k�0��ˤ�,UO�KD`1U��Ut�%ڳ"v^�ύ���|2^��Hݫ���ΪZ�<��9c�GY#C�����c�Mi�ܯ���h��{Vn�\�D«adN�v��=곝n:Ƨ�H���$�rp�L�G�ϝGQ3LvMQ��m\vUs����S4��b����aG���k3�U��"����{#v�(l���3l����|��;���SھV.���]s�c(Ɉ;_)Q�f:Ëoe%�&��S�ځ$����]�8����e����5[�Gq_c�W�"p�oAf����Nټ�M�f��C�Za����B7wT��<�#3�uo�U��-�y�
�}rs2��SM_K��q��S�Te��b7\R�a�<*��݄e��т>�0�$����5'g!�~���}~�@�va������w�س�23q�G��b���z�����;����Е��I�fj�r���Y���uX�yKK+=Ŀ��P�7�r_Tx�wD'2׶oI�5/x���a9�}ۙC$cu�dzU�Q�����3s�D�b�%�b�e���o��u�345T�Mª2�[f�z1�j{`�������%ʗ��n�V)����~�Q��ݎ�H�i�>18똤����|��|/�.jB��K�H�s��k�]�Zj~m�HP����F���`K��qxU��u~g���.�������P�7����!kI�op���Je�v�����M/��6���9��Yx���Vz�R�u����I}d+�R��95�ܼ�k@쯣���^ĉ�r�K�Y�^����u9~��4%�$V��^B/Z�+6j_�26n��`�����6�&總`\��a��5�'�U�ȩǼ�p�~�7PyRv��GzJ�hnt�н�JiK�]���9L�e�w�E��\*�ʂ��n�+E[���h��MD�VJ�}2x�m+����s�'I��wM�SDM��['\҂E�vR|B���oWrW�V��ʑT�wxy3�d����͜�,On��&așn� e	���)�}XE�zf�g��D��]&g�8��EX �M�PU�]~^������V��4k���/����R��ڃ���=",ɸzvW��o
p��f��x]ʹM�a�C��d_j\���p�ES�5=��~�Y�6��}��W�ߥj�P{�@����E��,4����N=z��{���.�90Dm4�g�����g�ۖ���q��k�l���D��L��MQ���_)4W5ي�e�u���GER�2�H9;2�E�L"��	�����g�):E�'���ނ}�ڞ�Ƈ�g0/��d����[Y�.P�����ن@����T��fa"�z۵�p7�=�9�3ωr�Tw��)D&w�}�#r���Hգ���]5���]��ԟu�A�-X"b
���EZ�,��s���N1Ox�:B�h��Q�2�%�m�XFd��=��O^���@V�\��(:5��I����"ǯ*�����V�F\���g��z�|��n� )�X'	N7۰Y���S��N��kt\���>j܁��j�vTΕ�4vq�L�%�Q���5�@����϶Ά���oQW��*�� �{bcucy�j����ٛ��"��7��3��mMa(oS���ni���+]u����z�#��/���Z{E��n�l�N1�n�[�51V9	��SV!�E��[��h�QF�<y�:�.\�ʅ6U* �3
&�r��b���e�f�I��Pdڤ�ruG{WB2���Z��mq
T��n��0q%LJ1�Q& �t�(n>�l�{��E�[��)�^%�/�ԑ�g�1y[/E�j�o�t�.ax���$v�Li,ɴŝn\�H�ەc���h�����:��?r���F�JU���쪊�J���&J7�u�{�K��&	�%�ntA �����_Z';�%��KC	3��mJ�~��T�����	�-n��^�݂;� 3��R�+>��>>�@g<�D�ŉh0��>��#Ǐ�}p6�:������G/�T*�}�&zf�;B&rV\a`)1�F���L
���D֫��j�3���[�����9�GB��y��@}�@�ceP>ӂ,^�ʜ:�O��ѡ8�[�'7�r\�(��Pld���J}�����7�֓���.s)a�0w�W����Ax ]���(�O{l78�T�������[vS:#�Tʩӆr�W�_[��c�u6g`�-Zڒ΄��q�"��sk��o/u^����|1�E<���l�+&:�ӽ:8i�o���5�ɨM<�p��4�;��eo�mpΛ`+����Nܵػ�Xp��qס#,�¢]�F���3/�\��{Y���[F<:��0�ɴo.l2N���],��M��=!�y�+S�B�.+����U��]�sc����$''Yy][�٭3-Z6���x�~������ W�6�c[�b���#�4fЛ,Yܐvy�;�^$wV.R�����nG��Iv7��@{�x�]����K����S{̩�mKI��Γ��O�;`��j/Ґ��a��܂���.%+�g�g���_ ��h�ӏ�	]%���2��Li-�4
NL\�*��.�!� �H4�'�����%2��Aя����\ey�b��0������V�9 2�S1����Ku�L�nL6gX�nww#j�қ��<�{�IX��G�g��L��v��ES&N�Ô��Q��J���s�Β<������	|�:3����KzP��}q�	L��
U�{mp���Z]�r�l�e�n��h�m�O���!�`��\K��5alHs���6@v8F)D�V�آ��#�o�Nhn��)�y������3�=����d�l��n�,fR�s�i{�>��\�E����bf#�c�	0k)�}s����뗚	�n�W	��2�]9*�!s��C��#�[��ǲ�3w���'Ƨ���gyD}�.�F{�`��t~���z�ZO{{��K�V�s](�D	ra�a��(ǚ�P]�ı�=���-�(���Zۻ�5d�Z��v,]�!<D�3��Nfj;X.\�'9�:1�L��5FvF5�V��ѼG��kg>*ɨf�7k#Vٍ����}�s���d��h(l��T���F��3�ETe�N�z5.�zv���A������g�Fj
���>k���]/鲝�o6������^g0�t���F
:>�_���yh�0��\=�Xޏ	�U��ˁ���%Puy��-�Y�#e�-�mG���ԙS�^�`��m�S8:�����˥�8qO8<�d��'�̾��}��l���;�9~�/�#P�W�Զ�\���g�xk^�1�- ���0�L�x$�f�t�:��^���.%��W(Z��s1׌��]�q��lLI��9����j��.��q���M��bݹ�Z9/�-UMndf���.]*�*���j2=�o��΂@,����Դ*v7vDV�r��!O�R���:x�N|Vu�nGD	'm���h}x���u ��Q�շ�A��F��y�YgCT��f�gJ���}�7�6s�oT�K��4*.�������׼�p�?;l�)���#��P����:�$u=��+���@Be�L5:��왺&�x�	C���l��2�_w$F��Ҹ������6y��b�u'7$��m��J�l� ��~Ã��	��������e��k�U��b����3+�&]�{�
�]�P�Mg����`����՟):��Z�Fm�ϟG%����m�A�RE⽑��U�q�Ǻ����UCeR$w���L����}[��~xמ�V��qzz�H�\J~s�=�Ya.����8�p�+`y��H��<X�C�;dlθ�x�7R��f�K(֜3�i������Mw0a����d��|��U�+�Q�{$+6�y��6`(���K�s�)Ŝr��G�ڵ�7Ɓ7������\ ��8섛�ܺ���u�c�C�j���q��t
b�Ն�Z�>���+��Uo��7�
7p꤭���/��{�UĨI`��][=��rT��A�ٗ.s��gL&i��c��%%<sޖ%8���x�&bx�u�Z�̙Qp�Zī�1O{U�w'vV�P�,�NW�xP�5G3���ڬ�s��6zc�i�cxG+�.uy�Bv<��:�7 L�%�!��(m[�^��i��tOB;��tyv���2K{�6h1��ڥ��R���\�D�.�R�
C�����
<^ ��h��ï�R�;�u�N��J�i���M�V�Ȓ�nG(VK�]Q�=�,�t�
++lɦ��j�U����˥���5+��m�oy]rL������ʆ�b�Z�,�[[�e�
�O$��:�e��(��O^V.��{��Pt���-a��^Eto�-r$�ѧð�no&����Y�xf^:�d��ܼI�c�}���cf[N�]e�k+B;~�y���ݍBlX	j;U�5w�ݻt�G���c����ZkI.��w�[�5w��[ܭ��#��X)�Y�,H;����l���˒v�+]�j�	yvz�G_b3I�I�`�ڶﴕ�n�Q�$��ԅ����`̾��]���Cn�]6��z��Mt)��ug�b���$j�8d�elW��7#�Gd�}�"�f+]�b\����ݼ�CYr��5�(���5Cs������쑺|��xη��7�Z�\��,�7�c��=zH�"*��+rA���M�\�V��},XB��¹s�q�o+:���	�7;Yf< R.g*+��K+i:��I��7�eڲ�y��o&�ٮ�1pÁ�N��4��i���ݯU
��|1:��M0���\8iKoz�x�rGn�Y�&tֻ�;4:�έ��$@92��[���Yl�u��%��X�J���n�+L��;�X�a4U�ݣW/���Wx4ߜiPJ�6���Iա�LB�����¶v��Z��]'0���c��yB�A4����_'�v�v�t�f&���\�f�YF�+�8�J^=n�a�X�T�n�K9L�6�U��Yף$�a���X���g�$����H��,��Xg���d���е�Q�M�v�)���U����r�\W�3o1�@J2�b���
:���t�*��+�tf��N��z_*���	�J�� w���7�Nx�ɛ�t7���^f�;\�ՊV뙒�s��d��y�suX�������t����7�����-
����D�{[�˂9�c�z���]�m�O�1��vcѱ�	�9��Tn������Y8AY+:ܽ��C��A�,�������m��9����^�S(3��<�}�&�c�E�g�$zk�
�V36���(��N[-��̫�h��T�� ����2�r����U	����1��$�cl��o:�xa[�����(P�=ң�b�T/z�)���Nj�Ĝ.��%#�M����1��H2ʧ�e���
�奝�勉ֱ��Eh���YZ��-*��(�m�kQT

���(��mX�-(����*�Դ���J�V+l�TADE"���-�F�U�*X2�[Uh�""5*E��V��b���X�Rֵ�Z�dKJ6��(ȥ������*��X
�°�*�,X
����QX6�����Im"�aZ��J��X0X�bʥ���EX������A��Q��F*��(��Uj�LX��V1Z��-eUTmQ���ȫU(�QR�m�(�R�kV"+b��)P��E
�(�"*5%Q��VB�ŉl��*k"��,X���2E���,Qb�#��,E��E�@QE ,���F���X(Ċ1+`�E�Tb���F���QT+R�Q�5�IEUUB(�ER"`(��Q`Uc�kR(��e�[H�
(�H���B��`������������s��I9w8qb�3ke�p���fl��R����[��l�ξR5Ҙ�1����R�eq��¶%ֲ�y��8���bC�T�\�j|+��̖���g��F��Up ���/�5)+���B��r��Y��}q.�L+��.8ҝc�c�%��Y	��f��T2�-4�hWF�݃IwUE��lġ��rV�Ρ��9�=o���:��g<V�!!�8��Q�wm���j�^<�h�T�r������vyR���k���k|xwY��uu��ߎ��~ؤwR��& e�숖K9��d�����z�"���(k��f�i�H�J�Hr�)�쪿��P��9��\Q�;�yn��.�1T��jT�c�2Ao�5��1�:3�Y������ÿ=)��]�����d��D3
&wQ��=�h�"�&6O"r��ʆ�^���Ŷ�\U�s~�$WkZ���g�i�*ĥ}3Ȓ;�SKM�s+ܵC롇Ϭ��ۼ�]Sd�f8-Q�ua��F�J^����=�Q_�Y%E�,�d6�ow��(L��y-茯F���Y�"���yW�� ���0�Ɲ�)K�մ"��B�ˡ]TD���q�����;�㙏6-y�����m+����h�g'�No	{:-3,���[9x���Jb15mH9Ӕ�rA�%�\:-mNz��]VS��+�@����P�5��ɲ���De�+/���X�!L��鷻ڮmN "�xE�k�X�U�U�s�3�;%�
�p�s/�Mח�~]�[�/.yJ'�X�~�zh�R(w+����Yt��k���FqA�.9`�����Qk�Z��ҙ�F��|�����<�>tT���������M��]����$������Ղ��hs*�3"�s����:��u�v�YK׫�]�,�9��[�����X��&�e�x{�W K���u���^ {|��u�v
.�m#���������߭�0u�Z�DL� ���;y��5>�(��*��?uʲ:+��ɧ���>-����B�A���SW��u���~���%�cԳ��̋�o���G!T���+)C�7g��c�~s͗uWN���5��+�tz�3�g�,[��چE*b��+{�6�
�t�.��'M��؅%�ۍ\���Ydyk�\T���g����Ɂ|�@�k4���ZT��S���<�'JL0��{�˚*rb�v�F�~N���K�h�^;gp�]ֶ��yv�e������1]L����B�����j�>��ٓSm�9̔'m�Z�<���s&����y$�e��e�YE5Ћ�Et'�;+0kK��\5�K�'ɵG��g�-6�!a>�v�W.&'j���w�I�u�e�r].'�n����h8���tجhw���0������V�9 2�S5V}�GV�`���ܻ4fEIc&�TY���ɞ	8U��z���z`��.��1�u��j��]���7�v�ɰ���[�����@��YT���C-�B��u�L	�1Z��$,�GO�J�r�{�*�c@�B߉�D�I�p�/�8��9& j:�7�T�����+%g�R8Wq
�!i��o4��щ�#��U��*�w^מ��O����X�fw����hD	r�T9@��Zaw+�%A~�NR[�[�Ң�3D���`�t���3�`"����#�Q�\ U���<0������l/��Ln�Ҝ:�$|]j����;q��~ڋ7Z��ra��46TK��$v�D�Z�h4���^&�n����.���1��
~;F����xg�FP���d�/<0��V|r*LOe�Uk��㓽*,�-��-�mu�-�ن�ޕ,Ɠ���UFI��S���b��O�uuY2�����sxjN^˹�2[br÷�2�#��u��*�F���ȫ-���{oGP5 �x�V$fЫ�G���U�u��.�"%�:0�-9���*IŲ��%����M�N��U�vr��[�g98ps��:������%�J��Hk%�\S�9�����8�N�����#&�1[�gEQ�|Ydq���U��I^}��X�5CP�=<�lP�;G#�>��^꽎�9ٗ�ltz�n�����--�����GE�����K܆�igj��q�}�ǱP�ᇒf�$�f��Ҹ��	@KVz���#$����+��r�)�.꫊���03�D�#�U�rؿ3g��3�p�/��e�H�r��IՇ9�g�&�������|(�S}Z��[�:��q�cD�2��v�V,�jn�v�ۡ C[]@L����s8-�=f4����ê��{�#j��+���fT�mΦ똥E}4ߖ���c`:�$inzbixðA�����@�V�^q���g
Ou_I%�i���sR�CH�NDK���^�1<m\M�qz2�֠��j�M+��|�5����U߇���W��l��h>�P��H�9ϕ�w��m'g�4�r�V�WF���3}�yeڌ��q5	��ӛ�2q��3,� }&�S=��W+�)
��ߓ��j���~ė�-����	heJΡ��v���y���.n%I�;I��S�f�P�G[&t��GnN�n�e-�-�}-/���2%���=s(jc�Œ�"�L�4�9�;�.J�]�f�d)�$��Wb����T�}�U�3�zu��qN���9X�dh��w("�)ib��7b��\I�]b���6{�ȴF}�6��C�Wib,��Y�.��G��e[�@���.��͵��7[�����O�7�� ��ОV9�8���(}cՆ�V�Ϯ[�T<7�X�SE���
K���ϞfK*�n��
�������+��g�7�
*p.�~旻<:"�Q��i~��s;e�)]Y}/����u3�����O�镅�v�߄Xu󤅜����|֪洹�{ԫ�}��!�U���a_
z/�iΰ���(|b����I�!�ߦ�,�����x:3�#�B,͘��g�5�CM���Eg�q��qȬr��eY��v,>«<EK���w�����=;��VY�h���|K���vF��{�tf`�9��=%]D�mn!sx�Ld�@?J��,�6sœ�Q-����E�Bd�ZEM�<q��{u��x1��T�,��y��XaM0���M�w+��G�&����r�δL^��j3���M�ٔ�֚85�eS���]�s��t:Wp�K�V��R�G�҃��l����ݸ���P̅��)���# �Gnj��(n&z�ʹ2�˫�Sy�d\̘�ӛeh�әm��ܬm�0h��a�D,�(E�B����}�P\W�bx�_p�?%\�^V���Jay�m��j^%��{B��gPCq��&78.����u�aU�lm���wb����������Wө�t�Rʴ�[D��SM�H+��t:	ݹj�����'�]�9Ն�Z�kT�]��x�UEqY2}����Kʫ<�c:�s�d̤�H�A��՜p]:3�X;~���`�V�JR��m	ػ^�1[������b]�>U�/d�k�d+]Jǂ�R��s��ș�%�3�AY�ʕ{Y�Z#���o����GP��G-�~F�	,���*�^4Ж����q."�]ii��6�t�]:��v��L
=Jf��������<�R�(��Ll�|¾�z�*�٤�As��ś�H�D�`�Dc�d�1��]"�dR�s%�@�&#Y�(�94�d
���蓅JI���Y����_S`������%$e�2�#�ׂ|� _{|�Q��v
?v�MK<�ng��:�Qܪ�J�K�����YX��y�թ�!@��*�'��*�o-�f��[����q����v��̌��¡��:��Ujv�$o&�ݙ����q۴Q��������'tx=�:?��'d!��kb,�Z��}�cD��kWK���ޔ��CSsf[E�nT����vs*�T6�����������zrP�?}ܫuY��W=ҧ���o����	b��<5��5.��!�Bȩ�za�Ӆ�2�Ɯ���.�U���k��oM(�d�uN =��V���u�횶#���=�Ey���
��7/�)�
L[O�;b=Ƽ������kfi���~�g��٩S�I��jL�h̜t��r�g��L��0��z������/���1r�̉��ᝯ�\4�$�_�a d1�����M���4'�K�aC!�����Ð��/�e_����׽[�S�����Li�B�_y��wJ���P����>������=��r���}��ۥ�yO�K'y#ČS��\Q�,�N嘊]q�~��!�*f��.�g��tS|��[0>���F7�i�{B%���2�Q7�Y��Sǲ����6s�C�;����Y�׌L��`ur����t���E�@�R���7�J�fn�����	�vB��N�ٝ�;v�c���VH�
^�"�>l�r��f��Mv������<ų�^n<��Z�m��I*a�7����S���JsU�C[bǹ/y�u2!��_��s_�� ��:�+,e�WsY�;|/I�����7�z�Fm�W	q��1��J{��O,�b�ԍ��˭�ij"�9��Ra:�t4GA'IeC���\N�5�:�y�G��:�q���4AF��g�a�m��JĞ܋�Љ�d:�?������霤��b�7s��c]Grz5q�u\���ֽ�ѳ�t�#B�tÉ�B���kD�)�4�'Vv)ܱ�ꣅ3+��3�t=8k��o�����r�@���b���.�����f!�u]`�������z��*������[xa�͋4/��3DW�q)9����
�G�dd�wn�Uo��g����p�EVz��l����iS)'��=;�a[c�,����]Ζ�9���o���^3T���۶7>�ԟ��+P�h��YxG����a!�ܾI���@��<0.o���{sp��3�IVh\�Zw>����V>K�������������ʮ=4�t���|7@�r18����-��l��pg��4_�f_&�S�{��;B�TԈ�Pg��O��}I�ܠ�5T�J�RU��ۧ]J]�ܸ&hz�6��RŶ��͡�p�J� bS.f竘��!Y�/��hk��C�έLl�=ҸXU��R��Z����Ҙ7��0u/_8kGG)JK�� ��:է0��YR���o7�L�J�0H�mf%�3�BOո%�眓	>�f�ۙB�W��8b:r��~�}��i�ͅM�5w4팺�}ԭm�+,\eavT[O{����}U$�Q�犓韍CJm"����C��{�b^�D;��o�!��vդ�b��c�<"�I���긇���ຌ�z�Ŭ�)iݶ��'x;����^�-����1�x�2(M�>�L�·�ކ!�Ǻ����UCeR$w�y#�l[�0�e�vT�r���a��ǭ�"js�aa�Ŗ���c��)��d*�2Ȗ�gt���oryΉ��h3<b&����u�FD�N�D�?���KK%������qnV����o���i�'խ��ekm��t��V��Dj��K�uq'�D���{�S�s��Չ��B�q� �R�	�+G�H{h>���aҵ�|��v�.>DaZ{��u����H��郣$&5�)�K���tl�&�9
*u�g(��Gy*_o�il�P6�f-�2m]��z�oqP�d��zx��&�V
��6z�_���R�n�o�tΝۭ��>e%t�������ب4�X�|K�����y�tV&w���T᳼Y�T������Ʀ����QL��$�+�ܼ(�ʲ̿(sY�h@x��QŮ%�:���
��6i���6�5)vY�:�����xE&V�r�2;1�nsB���5齻��0 �!5��qX�E^��V�o�Cn��^:���/N%f��_��� }�� y�ݜǺqw��7��U����CM��t;O'��}��ȯ�v��*�����`q���.�t�mcGuF����Hy�Ӗ~����J�H�\M�ޠ|�c�%RSÀ(����|�%��J��L91�s9�t�+Lgd�X��,�b��o�jb�r.�Gk��G��OVs�Hgt���Ώ���X��S�)EӠ!uB��ܮ7��a5r�bNl�S�d)s�F�7ŪV�*n\nT1j�
��>�C����+��.4t�����:��]A]:���Ǹe�	������'+���=����f�Z}ʄ��)���{wǘ�/*�fI1�T�2i�w�Wt�%�D�k�j���ua��F�`����d��h�+5OJ�;;m5���J��Q7��?x�F��"�~
�T�s�J��h�}	��N}�;J���O>]���|!�db�"\��� ӄ3��u���W)@[';��-ͅ_��Ճ9>n�g�J4��u�Hdö��Yd*A�S�%i2�;,1c��f��O AK.F�[�����`+x��6i����jV[����x�X���eԙq��G;�u�В�⢐��(���C���8��c��������TtN!B�Z�S�*�m�RDu��N��hX4ku*�����6Q7�t���\O��@��Y�m�}vi���: ���hAi
	/�z�;̞;Ô��:��#��@�끡M�W+Z�R��� �Z+�[=�nN��m`�Y|KP]��Pt��X�W8�{�è�ݪ&���̻GGW8{6� �wsB�rw:+K]Xa���c��Q�R<�F��*�|/:`�T��ۏiU�1�ڸ���]�6������K:�Whi�E%�E��-��F(H�����W2��b|*��	om��c��j�hF�
އ�c!:N���0�M�j�ՉE�1}���Y�T�ٝjl��ᇎ�J��O���%P	��Y��R�Qt�^�ݺ�J�2�YW�޲#���|/�c)n�D�;��F��2��'9��;޳֨Нe�pa�~#AWو4&`�5'͍}h���7G�k�Fy���]F볿1�a}w���Ѐ������C;�"vQ�r��ĕWr_ vK��c��6��"Jv��S��c��e>�����u�i:�'Q]�Q�����9\��O��dx�Rj�������sܢohk��4���\t
�Q�k@ǣ�J���� ��z��Q�SX�e���d�OLJ�����f|���m#�apД��na�7	H�ȟ�UR����� uop�����"����̹�Y>�/��NY��ܕ�M�.'�}Jw�VVي$ZMm�CҶd�u��g+���F`�I<���[t:�r�9�6�Vc��=9��R�P+��U�A���.��U�[��f= �,T��7U��ʋX|�f�z�)_N�n��y8ǽ\���I�{،��P@�.�v]��|��5ls�"][]H����R�&B��5Zre���r"2�{�M��Z�M������\�;�Jz�m���v��TwO����O^ɂL�M즫BIS+Z����l�����h�Rf�4�HY�{�X�5��ETܠ�u���o>乞VY���qm���!I�
C~�wto�'Q�Do�K��i�;l��LUXV��/g�u�p��N�LJ�w�
�Je�J�8�-�m��[HU��@��� t,�z��9;_$A	�v��wb���ju�DRs)Ӻ��a]�󚺔��6v��yܦY��
��^�{0����3N��/�r��V�԰����Nf��r|�̰@��RVe���b	�m+|r�q���;餲)���o�/��+��/"�-�����:���N!S�-&���]j�p��?��6a�n�
�ޢ�G֋ͩxN'h������2gr�(qI����U�X�fm��}|$��'�A��	 jVE��QAAb*(��Ղ!mж�XYmE��,�Ŗ�R�,TUDEm�EF*���Y(��
���E�b���"(��+`����Q�VV(�`����DQDV(��UH�!Q

*�Ī�EA��Y+E��0�*�X�TTX�Y��QD"���`��*#T,TETF���jT�BQKh�E`�����(�DV)�R,)Pb��e
,DT�
�B�EUTEU�)dX��*
6�
�E*T"��"��b"�F���Pm��TlTP)T*�U���(T@T��lY����(�hڬPTQA����+R*2)����Te�*U��b�J�PEU-(�[J�X�ER*�J�U�l�e.%H�QQ1~� �>���ݗ�<�f�#0`�ҡ�n�����Y\� �EC�t��w6TB��)���u�$��U	KѮQv.*�����z=��7�ǝ�e.7��� 7\I��'��a�7�����Qr����]1���p�B�#F�F8�x��S�"ՈGQ4��tQs2+˝̗�ĝg ��g&��[��0�x����a�J�Q�f&r�����ԑ��1@y��򄙱�`�v�t%�]O���W��SRm�����<Z֡��8C�ëS�B���R��{q�/�����1^ˉ�3
�ʱ�ւ��V���4��zc��c���\�u�5��N��=������><h͛(Q۝�zs�ڴ����oM(�d�n =ؼ�+�{}.���˰V�ZW`�2�8G1�4D"n_e6!I�i�Gl{�y!cb=q�Q�'��U��h���&�Ɠ;'3'9�c��V�����6�cHY˚�91{*�6y̺8c�$;�VUAg(抚#���'Fw��X<�Ok�6�2!����a̋���4�����I^�n�t9W�p/Z��Jo����B�c�<7��1�.y�zqQ��]�ͭ[ryu�9 ������U>�8��\rX^<�{�V�V�2�j��އnB�r�t��\��	��T��)Glp�LY��f��.M�ہ�T���zj���Yj�T�b�f!"ph��-�:(�������5�%�[b�t�t�&�6�Ͻ���ވ�x���^��f��r�}0�d���F)��8��TQ�,�u~܏�_Ps�D�Jodq.����\�����=�Z�L��Lh-2{
Q>3Є=�Ǎ�>�zq��Zu���e#f-�H�kGJ�,��C9�4��ut�%	����/D�{�y�m�`-�ʷމ�W�ӗf灶��l*
Z�D	r|�0��U�f��M%]�Ur�7�,ۤ��,�w2f�qAuY�Vn�a,!����#�S��%�E�aER'���� V�j���a 5�ĝ��^Y�PI���Ҷ��b���b�Â��G�b�c^@P���j�ٷ�櫅����=�{�q<,J�cC��Ld��Z0�<smxc�ni�]g�r=�h�x.NѺì�H�>UȃhS�Љ��)�g%�� e/���9F3��_��r7iK�'�˺�Eɥ�>K��u��\66Zu8�J�X�2nS�1W��:����Ǎ��_���I^���I�d���x�FߚH��㉉l����UT�m�U͞�Bgn�؅�{��nًH\>D�3��d:T/�	uY�Ш,R�\��/c#m��prj�Ձ7E<F�;�I	��5�yI{�qW���R��F�|#y���/w
��!���t�:ь�ʄ�buή,)_�d����t`���`���CrD@����挕�>�z=�z"ʷ��4���x|̡���C+���<gڗ	\�ww�~Ɲ���g�"�6�'l54;j���>��o���J~t�ʡN�p8��Ę�y�A�a3g�������Wc�A��lV�w�o���j��[���k���t��Z"hn��S�t��Vp�a�;*�s������;ދ���T)z���Pҙs7���6p��Gng�ff�Kw�����w�m�y�ow{3�N�
�䎅��eE�8��o˂�"RA�pg��~�����74I^зr��v��\�;3�[�"Em��}*Qƴ�B���Kh����q/��ɚ&�W���r"��f����y��a�]�ي�,/�M�Eޓ�"nfaT&D�u'�6
+'*
\o����Ga����k��MNt,,3��&�����>�.��Uh8ONR���ʄ�V&��d��{6�3�&��7���5��+�~�u�<@C��`��+���֫�Z�y٥�M�sG{�5.nD��0�حgf�n��k=.ƽ�g9��)P�9� ��<���b��}u &2��=�g';���B��>V�=QN	��@�lT5�7�S��8t���rLOv��>s�U��΅���aPX�X)mp�s�NG[���I���8J��S&i�v.=�΄���rk�VR�{&�GmTO*ES_�����RK��u�ѡD�$�ֈ�U��F�K�g���FH��=�§i�����U>rߺ7xD�)�����}%=�`�M��:��M����Q^�����#n�ռ����;�h$�A~�z�Ƶ���2rF�ˣ'gK�/c��ױ�d˞���>v��KQ����NƘS~���򉷵8R�����+<���y�tS]/�d�a��Ɛ�m�=��#p{��Z9�ׅ.�PC���ڠ�c ^�[�A�^�XBzJA�=֕�]/UCѳK+]�h��D�)7�C��H�\M�ޠH�3Z��jb�����d�j��5r�"�
M�\��aP���R,�q�7S-ޚ���A�9Ӗ7t���J�&\wqsV!�G���,��M���
r�@\aD�@�W�.�0r2T���Y��m*��������rv�����P�r��ఞ�F�
��u����B[�#��:�e��hz�؁�Fp��Z�;�hBr���+��g���T&�N�*���zW�^���&�L{lmD���WDV꠴��U��<��V�[�������Ѷ�c�lb�k7-@:Gja�����0=I���o�a�r<��V�X}4�^�>��M��]\��)^��d���ǋ����o���G�!��{f�չ��諭��{2����&�)~��
��t1g�_�D�k�j�S����@j��ue�Hz�-@Կt�}����Vh��N�ɒ�7�~��F�y
�]h��}�����j:\8v��U"iR\�s!tv��eeQ:�h�ǜT"�FJ��tR�3aY�1ќ}*��(^��K�-���qpmm�*_���T�{Q��:��w<̮i��Q�4a����[�=�����J�K�-#b�,@+�Y�5s�>P�����+�h���_>tT�5=	�4������_=_R9�(��u��S�5[
�mY�'\� =�`\�#�2z�wzb�V�x��3�����N�Z�ɾ;@;�)����-{�q�O�����"������8}�[�.|���*Gt=&���\�o��������[�Һ��⸹E7�'oM��6�=���hS�N�ns�P�[�X��=�r�=ҧ���?+'�/ �V<~��ҝ��'بf�+z���i^� ��Gf3hM�,й۷�>=�Hɬ]� �{�����d���-���f7�wy�#x�ҭQm2S��'wU���wuY&�[V�O���
:�mq��P�����*����b�_tL�X��gu��/�]�q��cY8���aD�w=�0ӥ��2�:���$s���N���w�J��L1�-c;e��c��W�U_UU��.���.޹���ؙ1�5�T�X��}�؅'�:m�q�y���_=�2�Y�#^��]i8oOji.��:*LN�UJ��L̜t���)\*7<�z2��Li=m�"��)U�hח��oӛ��Z�,�8�l$2� q3s~�M���4'�Kr����Ϟi�y<9>�{f���`$���Cp�G�U*�S|������P�$xo5�n��Ƕ��..\5�fDw6������ë��z|��^� ��Y���%E�픮c��:���l�3�9�r�BC���K�{*�4y�Bc@�V�Ox&�}��.b�����Yrp�cê�㫢��T��Զ%�&P!�������'W���Yt{�O{MO.fN͛�>�����6���E��:���q�<-����hyl�u�G9�$�O!��Rz�I?s?jE']0<�k!�
�y���������C/�w��b��~����w���	�e��z�f�OY�:��l�	�g�~d�1!��u%gP�l2,����d�I�w�>�h��3g��q�����FeE}�6�Z����'�X7���1�S�~.a$6�_�q>d6�P�g�&�y���z���u�d�g��M3��La���Y;{�{���G���{k??�i~����x����S1_&d�s�6��QŹ���3�2���iZ��T\��}pm��p�ޥjAcf������nj�q]����
9���%���_H#�����bqc̡*\�y3M>o�t5bJ��1��\"�1c���{ގK3Q�)�ً�O��}��=_��y���
����<Hc;g�\�Hm���=���g�N�i��a8��4{f��I�m:ɏ���~��|��w�9���>{��8|Ȳq��@�3S�s�"���wD����rOXT�����!��|Ƕ���a{��Y?!�'�Rq��J�S��	�Ce�7;|����科��x�Ͻ�10'�r~Bw�u�I�Ĝ@�d�N~��u��LO�w$��L`h��m	��>O/2�%w��i�@�n��?n�����fw�}[���~vLa�+6��̋���l��x}Ld�i'�\@�'��~9ܓHa�~���O�'}�P�m��Nw	�>f�M�'̆3��ޯ柑�mο{�1?g�;���k��'����O�����E�~���&�ԛ�$��8É�Ne&�a�w������ߵ8����GnoQ�}�]��X��/���ό��btt�OX~N��CL�$�9Cl�x�٫O����!�����r��gm��0�q��k	�C��3g���UP�G"�`���v���#�>�f��l���=a��00�J�/̓�G���~O��2~N$?MP�Iǈz��0�>��ߩ�N0�������������瘟�J���߾;�I	�u�������°���i<9܁���W����xy�d���wL����5f x��P��!�0�c��K����?�$QF�N����]FN2��클:β~����9��D��a;�+̕�$��䕑I����N$SAw������Ԝ�H�o����Wv��Y��n�d�EO����`x��L�z�x��m�C�������g�NO��&0��I�|����Xz�^�y�rJȲq�����\+�Hx�����g��}��+jVG�;�Ԣj���nc/Y-=�@��^i��c�N_��J��2�l������C�9{ȋ:�W1����=�)ø�i�Ur�SH�v׬�ut`��R-����̰uH�'|'G)UT��3U#u��=���8ޞ|߿���9�,}��'̇�UHxÉ�~�x��:��|����M��z��=g�Ra�&���S�I�<3�Ԟ=d��Ǧ}�s���]��.�_g:'�z�)8�:_p%@�(}�	��Xu=d>��8�0�?R(OY�S�:�z�P�̕���C�:�[�Ͼ�G��{�~_	����j�;�����v�;>��"ɽX}�&�1��������Ծa�����C�OY��x���ȲgY�N����ѓ�	��C���H�5��mI�/�幮sW=��E'gw���>I���I����k$����<�XM c��̐�Ci�{���&�xe�����z�϶}�>�t��s�2`�?���<:h�1|�׾{�o�����&ى���d�$�݁�"�����To�&~�E�}ܓԝt����Cu>O�2CI����hOY<���~d�1׻�^cw�{翽���}����O�?0�1�2OY�Ӭ�}By�:�d�c0:Ȥ�����"��������rOXT�ݡ�u8��?!=O����R���Y����N}����Ψ~d6�ܤ�+?>n�m�P�1�a:��錝}BxnΤY=��P1�����"���u���;���}b��۟jdJ���{���g\�>������1�'B�|�|�j��<f�5I��+=|=�8ȡ����$�}Ld��	�d���N T>���G�c�V���n�d]��o��}��~�6��w��=f����0�	��~g�����g���'��$�+�=�dP��q�	Rkt�&�#޴*b!�{g�ucT��?'�:�Ǩ�\���1�s�S'��{&=��rh{�d�Cl�'��0�a���|�3z桶O$?��"�����C��?S�"��]�[>��~מ���t�/8%��2�oj�L<"�M��̞ڌ���ޭ����n�|�|!�7�zzF��ž�)��z�Iw����&��SI�����k,=j㌱�3�Ԭ3�:�l�vE:�����ec�����c���vхʇ~�����܎�rO�K�T������m>I�9���Xz���u!�'���S�|�m���Q���x�i�{��u��?�CL��$?��$ϼ��W�++�Qh^c{
�t����T�E�~g7I�?S�8�a1���8�d�9��!�~���'̇�����6��q����a��5y�0�dS�����هiv:�K���.\��2}�;$:�L}����=���XO<�gq�	���l�d�s�!8γ�s�I�8�~��V�V|��{�q�S�	sw���k`��]���V.9�{�dQ���l%C��d�C���O�!�$>a�s�O=gY�q	�>=�6��'��;�����ړ�r}�~��}�;�M8g��.\w	�9�������%H�|����I�"�/0:��(yw��N{d?j�C�M����Xjg0�����m�C����>�O�'�̵1˟�_u��4�R[�n��}�c�a4�XN�ﺑdǨ��R,��_��|�/�n�(=��O�M��C�M���d=C��i�'��0�Nޑsr�_�v�=�ߠO�b2c�}�:[!��4}�5>a:��;��u$����Lx����<`bN����`E�Ծd�|�i��5���P��T�Ϝ�}1�����>�Bۄ������(M3n��N3�C��Vm�!�d�|�U�u�ý֤��	_�5�~d���1'&���!�y/�O�G��(���Ր��m�G�Eό��G�7�������ΡXO��i�&����u�Y+�=>�8�d���F$�d�kD�ԑO�I����7�`x��:�'F��ͻ��;��ܻ+~[G�z2}��xvO��~���=d<י	��y��g�I���Τ�1���8ȲuĚ>�:�d�}�y$P9���$S9�~���{��c2�g����i꫑羥m#� _ob��uV�BK�r�J'�9���UYN�GRI$/��7��f�v��S��99���g!�J�:#'	�&�5��G�(x��Qu<��sC߉Ál��jG֞��fI�R�"���&ԅ����v5�lqM��M������?$1�S��s z�m��Y�Ԟe����u�Og�	���1�a8��vbN��O7gR,��=�>��c��$r���3�}&��.�������	���d���05=��3�</r�M�����O���Y8��%g���	�a��i�$shz��s�ﾝ�4��|Wn}ځ�V~=哧�@�Lu>�������z���͟w$��f�o�|�b�����6�c�]����m����̖T��DG�Ǧ}l��K��Z	w'~v���bx�m�O��>z�yˈd��O�;������~�?0<��P�m��C��>g�i����	����!�}>�����\�O�qY
EX�cᗔ~��79���Ь�&;gOhOR,3�7�$Rh�8ɾ�O'�8É�Ne&�a�s�����4fЛC�w$�71c�}��{�>���k]��[�~ZVfr3��vky$��$?j�ċ'_�紆�C_��,�I��N0�u��'�C�8��k	�C�q�rC�'���}>���|�<����s1����ZK_g��a���ԓ����z�=Oƹ��'�ڳH2s��)@����'�O��'L|�`u�|�޷�z���#��R�;	���_u��������?!;7�V�Vq'�{�:�+��q"�t=N$�'Ʒ��N>��f x��l?y@�!��x�2=s�\F��}aϽ>Pd��<��ǰ��﹯w��g�`|��N��!����ޤ�0��7�a�JΤ�JȲq�ܤ�$X�C��E�.�d�C�1�M��y@�!�=>�ft�k���7��������^���Cl��Cl��~���:��<���N2La��oRxϘO���"���$�N<|���>MK��d�]�m�S�A����^{p�o�*�5� �M�-����1_^�݈���̥���f��.���L��XFӃ�m�[T`UwqN��7�Y���*��s�:JL[��̡��Q�s~��� e�b]1�&ޞ)�d
����!"���*ϰ7x����f�����Gb
�$Y�fB�g؉�]��S��V.��ջ�j��WS�ui�i�;�@.�w.�ޗ��$��6$�T�ͽ�tր���gT��ð�x��,���vI��	�"�5)��9�q� ʺX:�)�6`%��K;��I��x� Wu�ؐL'�#�!`�uG��ծ]�u3p�낭<�����3ehyh�0��u�1�vMUHn���c�d|K����볋�hR<�����:����S7���,c��Ƿ�C͹�X���aQ֮2�D�0�7�a��֟\��ޫW�RV�*����7��G�n����F��9�Zo���є�N��WN[�*J��z�jE��N����re�*F���u+�a�]J���F0�i9�*v�*-�Z��ܗx
�z����s��:��.g�*u�r���A���:�h�&(A/��@.6 ����R������5���+C��j�;̱Y8mD̊Jx\AnX��&��_fgn.zӵ�F]I�l���b��A�Sz�$�p�W;�1h��|�Ҙvy�gq�ݶ'6ɕ��,�K�_����;�T��$���.Z�*c�aR�gK��+�Hv���9FPc�x��T��Bԃ��RZV,�/V�xr�敒�e	v���p�}�����dx���"7��R��F��	txBEX���>�8���Y���6\�@Z��	���Fw��:��B��ٔN3AP}�, �fk�6��'��y����]պ��GB����q��s��4�CI��|r�ɕ��p:�p����;4Nxڣ��*��bI��,E��u��#4��f������k�b����EN���1dڑ�����0��kk��.��r��w�.j����Z��[ ��6-�`�L�K�ᗸ-.�{�@%�aP��e@�^Ț�ǐt2k6Ij�5��=�[�]����+�vW����%���r��]��.�v�Ňf�@ڢF�=]
��m%�s-��r�*A��u���Q��.��GVdk2�ï��0Lt�kV�N�Xc�;���t�	ǵ4�-]���1��/1�"QIܚAł�71E1!�6?x�N�}���ߵ�]ۖG՛R�+��bUkA�Ӡ�]��]]�p�u87p-��5MH��o��S��Ms���l���d�΀�ضoA�2((k{V��U8� <hn�iiƱ@���\�9���9����B�T���I�jp�tw�+&�;ZD�k��;��w+t���pEF����I��X&L�M�x�J�����y�	�+��6i��L���8�0�~�((T�+*R�U�H�
�TX
�����$Qb �b[TUV*��5*�Qb�V$F(*�E`����*� ��T�UDE�	i*
�b�����T
*�b����#��PX����k
�)������� �B(��
�dX�������ʋ*���J�B�Q-cmJ�U"0U�*D�QD��!���"��XB�P�UX�B�Tb��E�"����EX�TZőb։"�"1F�IX��EX���j�()QJ��`�,(�b �ڕ�B����1TR���U%eAQ)X�
~V��W%*��b+�QC2�*"�� �-�*�",X��+PR�*��Q��hEL��,���cE"�LIQq
�,X�,ַ����ﶣ��"����:8-�C\i\��w9�0n�Nm��fQ��R:�5�6�Q:���y�9S�wm�����U_}_ ��jp޹��$|�3G���@
#��'��YX�m�g��g�z[!��>�|�c��z�>�d�&? s��x����?�B(#���W^��y��}�����W]>�4��7��M��E!�:Ϙy�Ȳ��^��N������Vmd8ì��<�d�I��I�:�l�~ԊN�`k�ם�?yt~{�7���Ͼ�5�z����;�d�������|�i���6é�!�0'��C�E��7���4�Hk��u%gP�[��&}��'Rw�޹���<��{���w������$^��$��z�<���0�|����{/ru>d6��(m��'��$=g�Ǵ�6�:�7M�i��h�8Ȥ�c~�{߳�ns�������W=!ċ'}�5�%`h���3�$_>�I�
��������~g�CI�ڡ�C�'�a�8�̝f���ϣf#g�>3�>���7_�����K������M�����dY:��1������H�k�wD�����z¦0>��g��^�Y�����~C�Oڤ�̕��}���&k�/��������������0���c�$����z��q�I��M�d���!?$<;��M�����䞰����1����y�=a+�{��������|���������3����z�٫&�~IY�x{d:Ȱ��;d�Cߩ���$���Y=��;�i�>Oӻ�?$<�}�P�m��Nw	�>f�k���#�s����O����Yf!�v��q�c��p=d�@�j��E'�y�	ċ?S��J�Svu&�I>jq:��G�c���:r�G�c�r5�f��&ͼ�~�y�����߹6�0鯲M�l�'S��q�m���^�4ϒLs�6ɧ����E���y=�4�����,�a��I��L~`q���&��Y�>��~�������\�o;=��J�],�ϟYU�P��ڵ�n,�w�
R��U�w�5t��E����蚨|�R(�����ۼ�+��B�QX��[����e�51&7�q��ae=�gh<O�CO�w�c����Ͼ�G��Զw��ƴ����9�O�yW�#�}'{�Y�O�g��8�*j^g̓�'��!�����k�d��H~5C�E'!��!�0��O�a<@��iq���ُ��k�K��t�O�ԇ��>��6ϐ�y�H|�x�����I�;�8�Vj��Bq�O.�x�=O�]��'}�?MY�2s�9f޲�/����i�X���T�Eϣ���6�x���q���C���C��'����!�:���}�z�0�������$�JȤ�q���$S��Co��uQ�(u�璡���M�I�����<��5f x�i�?O,B�~a4��m�C���紆��z���wS��y3�Ԟ3�'�°���@��k��L��\������;Yǡj�qP>N�r�d�</rI��C�<a��?P<Hu�|�>Bz��i�8�Y:����C�=d��<���c3������{KQ4�a�R�z6�>�7'm���_d������%dRm�</�	P>f��݄�3���m��5E��'�<'�E	�8��:�z�Դ:��%�l�_���ϣ�n�z���M��#�O=��߾������9�I��$�w?h�'5`y�a4����;hE�l�a����3YXq=d?����:���E���'G�c�O�}�q��Z5귇彯��_o~�8�l����l2)3�sEd�I�{�I���2��N������@�N#l�$6�����	�L���C���>qU}���}FO¡��~��osE�����|4�̓����M3�P��Y+�5���E���c	P59��L����rORu���d�!�:�'�s$4��=�6���}�n�9ú���Z޹����sz�x���O���Bu��=Lg����q��O�g,�La�XdRW�w	ӻ�����rOXT�ݡ�u8���g����o�K߷�}��;�N�^�Z_ݰQ����"��z�Cn�mXޣ��R���S��wDnr\?M�	����	���R���ѸNiّU�(,�7�2N��S]i�l�ͤjP�2K�ŝ��Y��}],]�m��C��� >����ڽ�|�O���z�~d�8�L��>��0���4�N0�VN���gR,��d��u�:s�|$P5;����&3�=���H�~�k�ȿ�Uw����&*}�uBd1g����O�P�'�m��:��J�ϾМdP���m�q!�1���'��@�O{d�� q����g>:�8�XKj��-�Y��G�c��%���l&3�y�z͡���!1����^`|ϙ&y5�C�O�Ʃ:��%~C�l�0�g��&�N�o�����-�t�7��s��O1i?	��1�1��O���?�������~��6���'�z�2q>���l=g��L��g���m�ǉڰ�"����C�!�zf �m��#���ްw]�+��51�L�������L~`u��9�M0:��t��������P�����1��י�I�����L�	�~s!�O��Y�yԪ�&�ndi��v�@��ϼ�z;=�1�5�ϻI���q��&>O���q�Ú��!�g�gtO�;����ԮP�D���f�_��{G�ھ��=޵�>��7��O��;��cF�f���n�^�>������'�;�.(w�z��q������*��5N6��Ƴ����H����a#]��2wV����.��Η1X�W"��ͳ��*�18�t�w	�^L6DO�����)S�J�ꨋˏ���j���ӳpp����9�zwS� ;7���St���C���6#��ܕ3�WX�	�sYջ ��n��/.J��rػs�xb+<��̝�]X"U�j�A:̦s�Gx��7©�+�orq.��-Es�U�����vT|�R�$��DDD{���+�t�^�F�[��]{��aջ��d7s��_V@�Y�p�*���{�ջ���Y�+VN�Ju�FYn��«tz�%�ݧ�[u�P%$�z�̚�����/:]{2�'#9@����l��ZGO!2��;;Ԗe�����X4O@^PǷ��L�Pg��XjW�-�^ѵ�xf#�	k�>P�%{�2E.���Fi�q�F+z]�e}����9;.{5)of%;�f�4�g��7�/^H�v��0��+�>��+Wn�h.�0�7�#)��[���sي����2jU�ۋ�9~�Qէ&1֘J�:w�k�ۃ���5t�{	���ϭ����}���@<�t��c�����IwUY�F5p/�TF�g�I
y��F"�{�Ov���q=F{
m\ڵF��NR��[c�����EQ�q��2���C�F���h"�Q���J��)k�����[f��ћ��+�Y��L�\p� ���9����UC���u-7�W�Z]7uХ�_Kj]wC;�jX�� 8o�f�l4�[�:�z8�pty��}�����D�J鑀��F����z#p�V9iv����w�Ԯ�q��]:�uE+#�"��i b-��L���<$�Z�/)��[T� �/�i��"0�3��x��{n�３�f�U�Ȱ�~Js�w�۷��OO\-���a.�:�N�����n�R�T]��Z��KW]�{!�v;VM�����Ʉ�E�uK}��,�����FO�N7Օ�����:��3ʴ(��w\}	��w3^�y�`���Zeԓ:��Y��[�ыs����ҝ$e�-��9T:�(աg4n�.������T⾣�ߣ!E�
��.J��c�ˮ�8���K���2��G����H�>�o�Ƽ4qe痵,��^|V�U����[\��7Q��X��e1���)灃,�z^
�)Ou�$�1(�{M�X���� �����|Ń�$W��e�Ì6��d�����]@�Hu�Ӷo'��\B��V�º46�s=�P��6��[Y(v��a�v�ε�Δ.�bZb�2�e
��x�5c��u�|�7ot��6^��n;�ZP�CCp�^0�۶��:vc����'9!������j��K����������שֹ��_�/k+Q�k�e��i��+�؄ �Lm]��oRS֣��l��Y*���Q���'O��;wv:ka����ګ�%�ha�Oup���÷a�Qkf�^�����T^��b���bD�TJv��ל��E-�P�\1������l�k���4�viKb��	8��؞Qn�|SON�hMJ�W��ҫW�	����[l�����Vȧ��`Ŵ�*�P�s��ҚQ�{u^�:y<�/�=�l�o���FU�&-%���OT͔"�馎��#���`��',�t4�4eԹ�Yq@�'�.&3S��Xm4�==p���N�C/b�+.r�iY�ʞs�f:���2�/�N���b;}��r�>/��f����$�*�3Q�T�u�Z�\R�l��TI[F ={~�+�1[�fl�-8vmq��D��;z0�A�ۊ���խp��&�>�tXW�r����-�W*�ۓ㹓�C9Ij���wE44��ݗ���n�{�gk�F!�Mr�:�6/�%\S�^jvo-ܚ6�tz�Y��agn"��]9�y�,n-����V�w��=�z#�[�~¾#T�Ϋ��{���	[��/�A�k;���J](���aU��Q�>��������#�yz<ڜ
�2ux@������R��N�ś�[�vo�`gB���"�dV=�����V���8Dl��w���H���b�����w�;�p������/�W(kΩ��+a�WW��ą�\vfΧQ�V˼���Pb����ik(�O7sݓ�0��o�z�@=��o��<����-�<��:�YB�En�`m�[��r ��>YX�E�y���;+����Y�k�����X�djWl�F�O�}H<w��[�f�-г)tK�ˉu��-(T>���:�A�SjR�y٨�mC����9$U���i�tSBjV�C��v�Uj׹t�$����Q�r��?ZHsQ�19/��8��x_<=�?R���#��+lKԕ�,�٣=�����z�i�+c��'>��p����\E-�ofZ3>Ηv�-=J�:⳺Q�����Y�nt�n��,��==4�s���v�7k��7�F�qy#�h�Q[�x�B��EQ�cU�G��{Ȟ�|��h���s;n)ՠ)-#�֙>��7��ɦ;Z��Y�UY}�h�|��ʚ}�%*QQ;�LE���v��\�u��Z��h�F�B�>�V�kp�3Uk����CɄ��y����Yu-��\d<���$��-Ρh��n�i��Ñw	�^L6f砭����.�����lҢ�gr�)�O�����j��[�f|��@r���<��gX>��yq>�<�YS�,P�nl�ej[�Q�G�ד�ҝj2ϛ�sp��ꠔ�@��[�Q�R|]I;y���_���봨_B��nE=5�B��F�m����pU���~e�ȭ>�]��QV}uh�:��s��S�}� k;�\�f(~�b����Q�>���b\vw��2r+	�g���w�É�'�W�Z9yr�{���P�e\�Z%^(��gL����O���Þ�Ke����@�UۡT�实��&�~�M��e�N���#-����g��E��+�;�R�/My�����p�I:��&��gvb�J�(hd�G����Wb�1�۰giYy�8-Ҕ��'R`i�K�4�Cs�fo
ʒa��}Q�D@�{��ή��*��x�+�ݞOt\sͣ���6��7�}�7���
�%�5T%L�j��]*m	��̓"Y�5>��nm;1?;1��V�WFP"�F�{�%p���&ѷ<���p�����\��w'��G��WeҫWc��S�Q��9�aQ��F�>��/��֕귚ޗ�[Q+�w�d=�{���:�<�~ݮ��k��9�aa۶7{s)��jnz������lK����Em,���	�CH�c6�����{�is����~OOZ��k&�J+ӯ���Ʋ�L����tj�ۖ*�9C^��wqڰ�-47�ޖ�,��
cI"u[e������	��z�G����3j��*�>f��\�.и	Vd�ED�{ŻSpo�����D�Iƈ����B׷P_\b�y�/'LD�In(	�tS+"�nk�Q�*�.w�=�Q+a��-e{�Y��TA������`���a�6mw����͒��O8�YR\*�ˑ^"�4Y!ʛ]s	�;|*׎=���H7mM��˺��K��vND�Ֆj�lݧ����G������uM�忣��яuPi�v�m�N��8��+��9h�gz��gZ��.�̎R��>b5P�<�ю��$V���n�4qe�5������C�%���*Rt�F��ǆ�)����)�~
��u�z�QꩢV��ͽu-��*��D�����6*Y(�)-�������k�}/�ouTY��8c5�ב��R�g�=�|�FB[/�<�\�C_n��K(����ߩ\�P"ޣ�Q���f��v@ΗU�G�-d�5y�R~oz�k�,��԰�}j:�ν[�>��cD���|��D4G�sݽH�Kv��[�끊ZU��1N����8�o �hc�hƽ�K�!zB|������zw<ZQ+�_����[�0���y��7w��V��6�Y��|M������r����Bj'��;�xGJ�nw��ܕ�*Z�m��>70���6�خ���*�K_0r���ӓ��Y�jU�P�/-�e�Z}����J�]�7zh�oEm@2�`f���[�(���ҥ��5���Ś�����Y�v��Jk���xe�{��u|뵈��W9%	�p��t��W�.�7�V���ae�[G)�ʕ�����;Xp^v=�*���Ù�:o�ӝ�*�gW]�p.�a�G�b���J���5�\���)qw}{ST0�\&��QIu��On��K��
������*�F�=\�YT3�oy���/�	�y�rz�*f='IL�V�M{9.ä��������Ӫ�9�Vi���]�/�]$7wP�l3s:����j��V帝s
+0�A����Q����ۮJL�jT4�Z����2��\2�:��K�Tr�,z4�����]D�`-���Z�2f���:8�"����^���D`l�H�6���kM��U������&U���}N�� �'�4[W&��k�؍'�OTi}����KX�7D��6";U�Q�!���kOo,�cG8�U�:�����\1>
v��^%]����b���P�ū���������7���Oj-[49q$@ܺ�"�s���e���x0�5�t:;p*�Z�$۷�rv�`�ޟwn�Vy��pT9��UsOA�&��3Ua�t.����J�m��^�(B�����ƶ��片�;u��#i�|�O:��rz3�'j�1옭R����r
���XǑ�8�R�E]����^\�i����V�:�Tޜ�2-]f�l�ۺY|�D��3n�E��S����	�Уݶ����`���:�Z���.����E�w�S�6���-�߶�7��n)R� fL1��:�f���3��@�j`t�ڲ(��u4�6��u
�Ԃv5�i��@e��v��qV�)��建]�Kr�L�_\��T��Ga���c?Nfܔ�4��$c�vA�"�uﺑ�M��_F6�h����J�Lݚe�i>Ipg�*3��Y��G���)����NkO�gEQ����rqt�oD�n�TWد�v�����LQ���Q��,��k���q*�s�c\���nPq���W�ƃ��7�<�0�Uh�]���c�Z�}Z'l4��'Y�α���r�c��U��p"��MD(�Vp��Q1��C` �9�B��N�=wn�)��	5����Md�۽;��50�d���Vj�5�7�s�d�*>�Ǫoq�6��^�Y�*o�w�\�T�"R�}w�O�Ӝ����-�I����/je�_]=��b�������[T��͚ߌá n�W�53#�4$Tn��^���j��y�a�d.��a�����z�\�~��˰��Z���ؐ/�4*���� Y3�G��?�{��z	�C�՘�u&�:P �!�?���(�UAE���
Ԫ���edR*��kF�#mE�D`��+&Z�AbŊ#�\h�YU�
��E��F�*(T���jER���Qk�ڂ�E��UE�*ac-*����°E�*,GV�*	-$��AVacE�F*H���±aY�*�QLh�PT`��X���iAb�%�`Ub��+*�Lu�L(�[R�*�aYB��W�J��*�m�%f0��`�����Ԕe`�j�Y�5�U*,+��LL(�ʅ�P��J�J�RԮ%AfE����d��nUX�+U�X��+�QEH�bJ���X\�6�Ć	b�����h��y�emM�wl���Pq!����D���d��b����br�v����g��E
;@d���fQ<��P�?W�W�q��u��!VO�(ڗ���ie�jf-�ʋo�	���u��������_�u��sn�CU��˗@5�({Ok�y�/5a������F��̹5�v8�z��rϾn�ͮ�ys��*�����X�(]�Fq��6k��U�˳�WPS�t"OGY�c�S& �|+�幃zNUK�u�V<n��2�Y���9���un��â��Nc���{±`%<X�{X��6gl�q8�n�yO�ͭ��B��*�9�z�����5�.��,�Tc4�G-�x���o2���25�`Cs�vEc�e��~SZ��bY����9���H����ox���a�\"���%[�	���e���m#w�3Z�Fltu�@Fl�u�Q���\b(1bk�'{�w;��I����Qw�J	�U�%�e�����~�}S;�j�{�z���D�QN�v�o�e���^�y����;�)*k9��ͷ����E�7��;��Um��U����}Ӳ�2p����HF,���:DzCػ���.O�z�9*:���$��n��NZ�<�l�o��{�M>ל��;2�}��b:���y���;�]��<;t�x⍹�Y��+�
k�o|�Eэ�U6��QK�ʛBl�T�̷ُ��tc��岯��;Z'�Yk�)�8Z��B���F�`�I
w��1m>�О���ݾ���
7��dk��&F'�Ŝ�T�=�V���H����p��*���t���SV��%	~��{^�E*�~�)\�i�i!z�{���21˔WcVs��5I������d����ZP�`<�	ꀸ���J�n)܉�{ݘ=gZ*�8��p-�W糲�Ʉ��Ez[�%9el[]���b;�a����L�~�篑�6;~�tQ�<�����n.z��`�3%��	Ys�+u�����̉�#<�v�K��y���d7=�L]Fq����)E��I;+�r�
�˨)��U��5��ħZ���9�W�j�i��}��- ����_[��ˤ7x}r5�[�Jr�����B0	s�]^���s��nνe�MQ��
��W"�ѝ�����Y�9��F�%\��dȎLIt�z�t���q��0N�!&u4��)�cV���Y���!j''5v �a����W�UL;�������IK���~�a߳L'����)ȮQ�è*�)��]�"uXUϖj
ofс�W_�V�o���1EY�խ~��W�Q����q��Q�o�Ly��\��r��3��6R��߂���R�(���� �u�:�Ǐmp�|኎����9��d��\������.��w>�̲�x ��ny��8���d�~A
�n�r{���ш��Y���b˰��*)���>��4��/��5��ӷ����}��仫Ƙ�}9=O�c�8�Q����@�=<*n(|���1�%q
�ۄ�rϻ%e����K�������}~�z�gA��9��+>��<�ݥ��!���wK�!s��i�H�&��K���S�̭]oԙG�"��>Q�a 㞞s޷���;�˅�κx��潲>�j:vă] ���B������e��S�Q'� �Zת�m���i��6�d2}<��->�Ӧ7�w���9�B&'w���Y���}�Ρ1���~��j֟���1wӢ�v��-���t�R�K;���aN���QJ�dg>��١oJ�F{��V*yb��#��[���ebۿ��c,���E����V�K+&5압k·Nu�hz���9�;tMf2]�gS��j��M�O\'��n��sj��<Y�+�a�]�^�({+bس��������wQ��0,��\�5�s'�87����P1��q�:���^�A|b�Fc��t�y�1�ُ���N,�|��O>U�ዅ\ KX<f�T��Y�{���5�,K���c,\:�2���a���H��q�Jh*���p5ᣋp��݀wI�X�����y��r�nr,vEc�,���SAYfF��|�&&j����Ǐ��:��
z��*b�8�>b�ג+��ĭ��`�'+D)=׋n�8\����oާs����c��qobB��0��a\��� �I`��{!���^MF�:��跫�V�px���<W��6+2p!A�V#wWG��r�\���t��\�ʫf�==X�1W�e=t&i�N�GQ?\4xXP�9���&����˴h��ES�T����u#VH�t��rJ��s�W;�����a}%�Gk핊H ������R��Z3.�e.�����}�G��-D��^-����Gf��������n(���Qkg^ �f����9wa�9ûmB2O{���"T�Z܆8lRү�c��7Ɠ�͹�{�W'�WH���`��HS}/W�ON�BkҺ��]<�Ui�XN��6'H��+'�l�c�W̛Im#�y\J|^�N�К��j2=�wDZ��S���R��h��p}��\�+��������§@���:7=a�����ٱOw?x�f�H��cq��)�v��jyq����d,�{o�v�u�z�yӓ�d�G�Q��FD��7�����ǆhX�m�[5B3�(:���n}�~�����F��R������I�����LA���<`�h��2k�Bx�fܧ8b{�x�~��!p誠��^�/��Ŋ�qˀ�W;����Э���b�y:e@�s�a��8�,�H��~$
�t��d�+�؇k���t,!�g�eb�uႜN������W��T�����:oxJ�:Zu^�b.�ZH㜢��'$k�}As��~�i��q�ݽs���Xa�a��Ջy
|q�edT:����}"��ic�.�/x9�m�T
��b6�p���W�z<����r����<�gk1�*7�O`��hvEc�l����}!�pʻ�`7����+O�����j���ʴ}�j�*���Iv�n��T0��Yu�ެ�~��P��W#4ĸ�RoS�����\b��U���o.�3���E�o�]��UKK���Pr���/�gV?�j�k]\՛2�Ud��Wg�\��v��c�ɩW��ԥ��(�!K��Տc��]�p���V��2���תof_ϳQ��@�Kd�K��|�w$����1�������4m�۔Л��̘�kZmT۵F���,�uj�$p:�_(�I�iU��}yn�m���K��#o�k��S{ژ��9FάاX��E+�:��&�@ާf��1���ͫ���ʧ�>�/k��چ��%,ե`���hG�'�h���_|/TC�(��^{j��V� >}tp��z�b�ue�-ھ���[�q���Y-8�.¦�^�xR\ݙ����Esh����{f4�w�3��v�"�3��Lp�&����.Za�uI�)kV�J�hy��+K�ӨK�����*�H���U��?F����[��K�	]tTK}wV_�
�ǂ�17���/N�Ʊ��nXe�|�����e�y�<�n.{=%laW�r���~�k_\�k�p龬�k~�3(Ö��6�s�V�!���!��s[D�ӭ℗�8���cˊ���+�1��sǗ$.���G'�Z�|�����Y���:ر��Vi��>����3�1�7h����/�}�v�2`l��<�{/�Ei�o��5᢬�.�t:�V8����trt��[\���u�ëW�����o3�߾W�3ҍAF�9��H����E��ZY��HC�NT3��Q�j�YL\������.�V-jk���;RWf�=��i#��J�R�1˕˓n�r{��mk�.Yvt�Eٮ^�:�W`q[�];������e��_�撵oW��U��+�v<� Xb���.Ȳ���b?R��6�u7�^񲆪�T�ٟA]�t��d��lu��I�ʝͤ;�9�7���*�ԕ�O�ʜ�9@���G�ݥ7�vw�Y�k����7N��]rذƆ5f2�1�\���W&���臭�g��f�;/�u�����0�����Y�	$)㖯#]�1��ۧ+I;��ⷚ��Y��vZ�u�+h�q�u��i1o"h�q�y!��p.��g�I8a��Ұ�&�%u��K/�����`>��xJ�r���
}�Ŷ�M�B-��4��t��s����X��%6y�n*��xҫyҵ�Gc''�bJ�gJ�pt�m�fu�ݢ>fT4Umz��E>/b�uJN2���V��}X6,�+��S��}�δ�y�>�KyІ���s7n�z�(כ�V�=Y[a�)�zuc�u������ݲ�:�b�Ե�	*�`���+���n*�q������[g,7��G)�����X��\:=T�`�}F�1G�Q�*&�#q�ꖐ]��������n�A玏U�#a�΁�-&�fw4��xW;���ob��amD��O >U��l��)��9y1�JA��8S���6���ŷ��O�H�*1�\�W{gv�&��d��q���e��C�pC|Z�OWl��z�8�=�L\N����E��#�_f��Kt��&��G�l��|�����u�U���D��6���A���E�Ec�e��R�E<�T�yUB�Z�f��Fk���O^�QF5��91�-�,M���K*��:�Y˯ ��j;�����.2�#7��ײ����PA[1�h��WS�ݬkO]m�DTP{��1 �ἥ㫫=�t��].��*P����5�GyȊ+��p�wޣ�������o�a�(Ⱦ��b��3-oM�g
O��۵ܫ$ ��*/oɻ1o��Rݥq��ˮ��tc��"�Y즻�;��;E8��oX��|M=;��5�]j�.�OrΒ�Jb���Jw���B���1�}�ׯ�>��������gvB\Б��Hʼ�x�>Z�='3����4��ֺ�J�f�}oyߘ�Rr���:����r��|��ʚq�1��%;�L�,�;�=P��^j���B�N�F&����,�6[����r��;z��-��+ �����f�Ö��S������;I^��Ģ⵸���p�`.�p�QYX�ѩ��Mq�����\8Ft�L��H�1]L�I��G�b�[H-��UB�]J	��N�RL�G o���)d�V��V��3�NK>y0���o��wV_�
�e��R��U֍Fv�-�y��v��,�AG��L��.Na���y{h�������zv�,	O���|�Ek��;s�"yoSr�}&?*���Q_Ta{��Gi�L�g1�4Q~uY����W��x�X��49�~�[Qnz�fslj�mZպD�8�}Dg�q��5,��?WSP^T^����u���f�K8���ج���V1���c�f�`+5��Rq-�+��ˍ�[�+�4y5يF�Y"�Xj'7b\3s/T���<M�-ܯ|�^R�Ǐ��ܪ�}���_t�U��\ķ�/<`�ۧs�R��0�j�"	�*zҵ�p<��O�J�f-=�p��|�X�a67����O���9>�0�vM=S6T�eT޻��1��~`�[HX���/p��>��S,mK7n ��w#r��%Q�K�k�$�:���w�ty
�[�V7S�m�Ų�%XO��I�����UL�MM�)\�Ⱥ줪1A B��2�VX�O�+m�_f����Х[k���)gdt"%Zξ�>5,�i&D��������K)��١��q���Z�(�Y�`IE�fq���ke��d�:��/u�rX�R���4�N���}ն�Boda��ą�U݁�Y�BzP+���栥i�]�����Mn8uQ�C�e�[&���X������VT,k}�3�n�M�]��c�g��T�~M1��t���^�z���0�V�E(]���͚ƧfBnC���kqaE�m�r�l��B�\0Т��─��$�C����ᇜ���V �Wp���S�x�M��M�Į�]sB���`��&reM"�X¥��wnᚸ�h���D�eV�	�Gt:�n�s�W��o��x�|�\G-aG��q�*�2�8b���:�e���fWm�!�]�n�B[)��_uW���q��({�a�We�Y�.��9��6��qA/�S��2�n%�҉V�����V*���`�Y��gU],Hd�{L�yv�S�s��v�o�LEt�X����/ZQbO 7:�Y��k�>��J*���rZ�T����T�gv���m�#Ut����T��lp�6�_Ċ>��Wv����v��m�X�1gd[�cmΰB*�5�M�L�U����\����*�q�m�����y7k�x�h}J�� R��'WA�j�q:{����^^���e��U��=�,Nt͈��Vr�v�%mI{��l��@�rN/n�L`x+L���wה��H�7Y�&
k;�FuY�ӱ��8m�O9��a�TY�C&슷���&-�X��Ԉ��6S���`[A�sM��;��¤A,�lg	��������Iz4���M֨u�glb���*0�^-��� Z#6�@'�7�xF�����Z��Y�
p��I�`��F�7W)��4��}�1u����Ω\Ol5��	�Yܻ�r%LTMĺa���jI�a�>&n��p�d2H��Uwh6�dUAha�O�]<��v���/�T�L33)^v�7Yt���g9�Q��P�M����oF:�j���j��*�E
R�9�*	�XhN|��@��p����ᷨ�<p��4h�C�t��g.������=��ӹ�]�ob�t�d�
ƚ�lw�P(�w�7ۦ`�H��Ȭ�l�����Ö(n�3r��|t�Շg*�CQ7%��n�z��9�!	��k ����O-O	�*͋��.9e��R�\���ѷwkf]���ބ�w�Q�v�`6�wƕJ�o��նE�wZ�RUt>��!ǚfw��*MAy�K�:ui�58���<��^>�mm�~�K챴9i��֖�F�$�wQ�X��R&�7ڦ%M)FK3XH6��[�䵩+U���
�.0�%`,*�I1rڔq
��N�b�(�dD"1�aR�J+"�T��-�)"�@L��̮R.%J� ���#%@�m����VH��IP�%m�"�� V���J�TQE��n�ҵElH�1mD(��Q�[11�-*�
+,XŭdX�!�LH��+TE�,"�f�MU����Ar�b5
�)�5%eeI\j��*�Vd�q�b,YXV&R�V�,ƫV��R(9`-`��ı�f �[
��Bb���ul5e+m*
,��!Uĕ�ȥA�PP�Qb���䨦[&e1��`E0UD�
���r�!�p�VbbcYFPiK�*&5�#�@�T(�P�KD�G�\+Wt��b��j�:WQ�1���) NI.�fH�5�^0uJ�A���c$�qݵg4�]
�um¿�
����WU�?�[��(���P/�W�k�Gʋ�|����_T/;}ij-M��%���ܪY�3�VmI��r�H��S�m��Xm:1/�]���u�z��5�/bk�r�5m�:�uE+�:Ӭ�I
�z]�WD�	DL�{9�%�~�oj%J*"wT�꽠y�=��/3Y�.�n��^�y�RG�S�K^\f�6��oge��	�訖�۪�1�뱻-,ݫU��nD�un�>�N���裠���҂�,�<)Я#���㈇���d�\:���ek[�fQ�ϭC�j�=�l���_TK�f��F�3%^��TN�N�TI��E&b��^N���6��zT����$r��f{�rq[꽣�A��x���#8���UFe
�ND䚘�3�B��x�iX��#��q��T2�c�8�����m�k�T���g��{����4)8��-�������+#U��T��֞D޽�i'=7w�Q����;[y[�tAZ輭ĮT]Ϳ{ʄ;^����`���w��P��nN�4�D3]�]-�Y5#�L	�OxN��iV8H�<=��l�;T�eq�ʄ��߼_wm[V�jǊ�r�}��ȼ4�S�Jmy�����u[3F��P�n�]|m�QdZ��O�q=��eگ�YL����7�E�f�s]�Upa�y����m<v�
��y�}�6��ob�[��m�˓���֋�����+��#���c�Bv���(���Wu�����ԛ}�b5���]p1KO
�ۊ/�r���$�J�o1Ku�ώh���n�ٽ%N�z�}@�e���>uɍܷ��S:$=��d�I�w,�֐�>hW-��O
E�5���E,�E:�qTR�S�ƉH.����rR+;A~��Ŵ��m�;c��NO�ؖU(��Y��Ԇ�=q����Z�@�.��]@|LcK.3S6�i==kg%��	.#d��4�,Y��W�o2��ˠV�.��1:��v����u���TV	�j��G�O��:e,���	'�r� 㹱C:Iy9L��wT�n�Dc���-C��uC.����p�xP�]�R�e3r,��bǐ�r�]u �T�Q;��FU�ƘɖGoN�@�Z��F�[[ӣf\���[,�3Wl��^���(����N��ȻK��4�V>�vs3�m�8Y��`�۳�V�.�X�U�pL��uI\��L����
��eV���T<Br�9mv�����2ϡ��~B�� sI�}�T#�^cF�:g�x�+/��wB��c�2�v�ϛ��y�T\���&�851�fh�~���'.���ƞp����E�Ȭxl���J?|�t�P,��gs�Gk���H�Pͷ�݊]��ƸA/ܜW�1b����X�j�7N���+�����to.�����Z�px}�1�o�W>����f��	�&H���� Cf�x���Yߌ�]�7�Pyq̫�6;���G�(x����=��������O5>ϥ�K�|b1A]���1%oJ�e�s>A�j�ۄݛ|�s�KVN�Dz����#G�8��e�ǜ�B���,g�kO(�e��;X�-�n+Q�c~��t����`�s��W��;/���m�U��a�@6V�Q)vR��;���c��v��rڙ)��+6)�5J�K|�Ui���+V��v�O+�$�3gG�f��%�+�\_�Ǻ���f�Y|�c�$U�8>)��i�0��4�7�p��Q�G�w`��,tc��Q|��������h>0�nvT��T��@F��U5D�."sv�j˥O.(������[K/5;{ͣd����ntb7\�+ԋ����a#��W�uI��Yt
u]�q9��ծ��)�ǝ������C��	�K/&x
cY�G���=�����9s'���Q��������,�(�>	�p��E9����VԽxNRЧiT<F���>��B�}r�=F�K��/L��	EU��F6�c������y�	�p*�(U҅��.��g0��;���fފ�ꜞ��α�gtR����n�}Vi���԰b�������#�Nl�O{.���5Vm�!uȭ1.7�+vma��Z��j��	���])vJ�����&CL��۹��t���=ov�BIH4�U�xx��1A^Cͷ�Y�df_�;M��oE�lS�l�[y3�����u��[4�(���bJ�V��&N�Z.t[qL̗��ަʕ�"�ʎvW#;D͵-\��T��F�OcD(���h��Es���Fi�K��U'��<u���(�/3���a�UOQg�
�SO0\F��^Ǡq��}.2���|w���]ES��r����o(J�Gѣ��,w��g}i�h��,�lr��^�R.[���䑼����ֶk^��oc�������2�i:n�tMf�����۵W��'iOK���(|���X>䑅E��AQR64��!(,�L��3ڵ'\�Խ��K���(�G�Q�i b9������k{殭��t��h��alM!�hա�[�)\֝Twd\�cW&;J��ǜ�qp�l�ɹ�\�ryb���4Ǘ,���*((��2����>�˹������Xb��|�oge��	�����Dh��YӍ�ܨY.��Yta��w|�Q�`s.����oѮ��r�n[������d�wGc�A��Hh�|�PY�(}�Π6�D�T�X�%u�����y��!�Uk����JE��{��[��O�
�j�d׉_7�}j�s��Z�t������2u�m�a;++��m6FZ�UG�w��↻L�Y����e�AZb,_1r��:��2���P
:��-�q� ������Љ`+�m��y`�9[=��f|O�/[s�	Pqvs��N�]��.�S�#�b�
���	\��m���i��>��N ��������|��T���*g��x	�X�'��)�
x$���Z}��9��9��ʓMv/�]��i���[�;"��En�Sh����[���';.�ٓq��=���>�C��cA�Rr���a��pH+�Ə9ݺè$���Wё��S���ej<���B��َOt �3.�s�m���T��,᧻�Y�}�����w<q@���]*ާo�	nTf�wy��Os�x��7�����r�]p>���(���E�׮���l��׶y��XL���^ߓh��{�Ov�ĥ�q.�.)U�����D�N�2�w��W/D4���e���J�C�;xfںͷj��D����M5J�V��!e��;b{b�S0��\��3i�d/�u�V�)�z18sP�6�t��s��Ct�CjL��ܬ)���r�SīC���TUIs���)~��'���+�G���sK����i�Y�5+�\�,��V����#2�4��m�˶�c#*/�>��>��O��;:��rx�lK0�Gu��p�%�J��Mvh̢,u��;���,��N��B{}p�ق{2��ڷ�m݊������F9N�/b�s��ZK�٩�ڰ�hV�Yr#3.Մt㴯R7�5��&7Q��o����]�,�d�ƞm���@�8Ƴg+W3��1=G�H�B�$律��+h��n*���U�{�<e�.⽝�)��X�e��~B�� %�c�K�1 �{��+��Gޕ���Bw�����t���OH�xl��5�:�xzϴѮ�MfwoW��E~���[���}�C[�nr5�����2�]���v��J�M��u��p��௫�{��늳8D�@k{����@+�=�SL�v�^h֭��,+b���ݥ��.��H^��<;I�.���E��Xwt�9��-�y���X�%A/�|�}%����nRm�Vy����^M��o�l�bx&�%�7*�7"ro.Z^89��w����%�Ub^���t�A�͌���ڸUz����t�-[����^��֛Ζ���s�����|�J{�d�����<�%�
�u�z�`�������U3à���F��۝B�\��n\*�8�G2\�|b��2��f��R��Q�m�ן
�	��5 oR��z����%�p�^�u�H9�	�+��5��;��yu���8Fr�p%c�ž)$�uQ�2\��F2��_+�>��W�r5r�9���sFx�TD�f�(��I�-ڣY��b��y���@wLhR�|jw.h׻��z�)C�6zN����8���s�s�!��'�|�J;�+-�;�I1�q����T��2��&��$%w����3x솻
�s��Y�S\��bqx��$`3
$��W�'��U�7��k�'T���J���{ٝ4R�3_O"&'�B�)_L�$�uھ���:��2�Z�6-��K���n����]�8��09��#��k�h:}*�r�J��Bɒ��#��b����i����Ay�u �u��^ �rk�fZ�d�Urc6ah��-����O=��C'@�[��1m�'-�or�`Y�P�)e�wG�ݞ���m��5ƆX��u�1�5�c5��Q�W���)S��{�9:�x���J=���GU;=�\���q]:1�@z����qk>��wog^�Ʈ�������3�ƻ,�.�ٵ(K��_���<QG�����=�Med��z's�N�\C0�R�yT]h��w9�����>�m�� �`����N��S��7|��V���@��JF�e���kҧ�h�:��\�B�Ū ukqtus��co���掣W�j�Ȑ`�D��V�W��:�2�����-�瓄Q��gY]}u�O87В�ID�MaR�a*�|�/r�)`��r�Ę��{��|�>���zf���[�<&������*�4����4�L�rE�t��,��=~��OFW�T0<�{M��O���L����!@�_r|�\���Y��Ʋke���������޵��{�Z��;� >Y.ȥ}IL�+[�����e�5s���3f1�:����-�$��1�'Q����xEJ}�	�hl��*��@�Y㣴�}��z!�쭭{ض��VQ+�-�1r���dv�D�J���.�p�8�I�[U.LE�38��m��-a1�t��k��bC�Ob�oۧA���ᛎ#GK"��̸aȭuB�>���v �����N�{�����2��G�שnu&R�{��0һ�rb2v@����n�ArM�vc��ؙ�H���6���f�@3�� ɬ��h�7eE���}��'�}�x1����Q��æzn�4�]9�ЁS�P��.�!SD$:�!6�r��Q�Y�{����=�P�^l'�Kr����`��\	<�y�b���_��44ָ�Y�����{�{]����N�b���|G�t���j�_�Zԏ��]��f[���c]R�fz�2W:�s�q�-|�f
t{�>�ioJs���f��v�b{���UQ�U����s�u�&���De
� Y�|**,vJ������$�GX[!�&J��ղ�v��=c��c+2E9H�y�V�&vx�tx�5��F�YT>�eF�tlxg������yy�q���s����S�A3��K�X�uq��Ξ�%�]�S�QwG"���˄��I�[U�B$K�ks���H��}�[��r��hm���b�s�k���4)����ɒg^]Q����5�@c^@V�x���#�Ce�W��e1��Eix�y��iY����V)��K[�����A�� X�4��H���"���x9�:]7�1)�:���v�JS��g5�<M}�B����`pS��X�����.n`�da+Ӈ��溲�9tc�x��Ѷ
8v�wGf��aG�)���ѧS!!´�g9՝��Z@o+��b������OCǌ�t��k�!ݗ�
�rE�c�M\{��R]���'m���Y6�pK�L=xj�j�Ѐ��$~S�(&��^v��j�����=#��ۤ��H�e��!=��M����If��(���c�Q_+;�=殦IR�zR1[	`6E>��w
[݋�Z*uv�3����	l`��)B1o��]�����r�LJ ���\�R��a�sF��e�+�M��;��,6�@���v��:��L�.�f\��ò`�g��1�@���{}��D�e%DðN�!���X���\=)y��f��@M���q�f�l�(��ISޙ�u.�o��oN�Ԙ�t��:��ù���B����V���X��Y*������9d�5]f��z�k���-�@|�c��wL��"͙�35"v���V�]R��I�Ռe�o.�n=)�cG���0�K^���Q�#�p!�jY��h��ٜ��c]Bv�ؔ�kV^$AV��m�b����f�],�yR��J�wf�m�-Pw��o.�d��Y{��g[��-��Yf��.ٷ��7/i�6�.�]t˰�I�ы0ե����C�E��Gn����J޼7h�y|�1�V�sq�xh���|�j����Q��r=�}K��=l��W�LAƳJ�$�іGI�ye�;��-�����ɥ�r����Γ�'ÆGܺ�����򔛳��<27�κ�X���2�L{�<�fj���_�.ij�Ųl���/.ds+�Թ� ���lz��i�w�s��;���[E��Iئn��F�s���<��q���"S�k6�k��u�[��d̗.�v�Ej�=��<�>�v-Nc�]gM]��z� ��c5tZž��ˠ���<��/c�4fS�e�Jp����]��t��D�}�AL̒���	�)x���]q�S�[�vз ���j���wi��t�]\�;*�I��a�Q���r����w0��#�]�f>y\��f���{�Z��7�-X�m�Gr�M�.]R6�Ga�ɝm�]:*��-K��1�+�-�N��Z{\9�G��4��������TQ���F�+4�@���+V(m���Y���s�[�$�hAqk�u
�VX�d��^v(�)r��1����P�m:�f(í�w�+y���D+K %0����o*_F�L��ó�Ѽ9�W�:�4Ew���f"�Ȋ�=|�p�HCN�r�񜹅�h��,�pS˕w�"�v]�`ӗ\v5VZ�<�Q��yu�>��yo	�|3\�e�2�#l�Pv5WW���s� ^��{Y&�,�>��S�d�*�����`��s�'t570���]�� �5RTA�B��as2֤�J[X�Z����#j��+
7,��vb�VA����F�k�6�R,���b�U�Q�(b(TG.Q�*WME�6)�X�Y�\)U�J�J�73ڨ�!��EL�kT��Y1�
�X�*����c�r�X�,EĢEh�L�)m#�3,r�-*���[�bYWJ�b�U+U� ��T�1s1El�sT�ڠjܵb����U��*U����4�dQL�-�ʵ�Km���X�)n[�T��F[)���2�km�k*��k�l�6�)e�f	qˆj�CV���W
fB�	�YW
Q�ʵ,��m���(�Tq*R�Sg����<��5Q.��["������ƫ[�..pr�������]���WK5
sxԺg�n�٩V
�g{ﾨ0�;�2u�����9�;F3��Ί��q���W%V�}~R����_��g�p��������⢛Y�V���Զ�x=.�2��o�t�(k[�\��.�em���Ι���GZy��\rg&��٦�e7�������;��!�v���̓{ܮ�rk�	�lݮ�w��U9Sj�˝�M�i���{�C C�oD�ʧ)��9NIS���[��E��v�9�h����#z��/���Gzm4_�Ae�H1+�J�*r��o�=;����r.c%����c��_[��s��o��P�S��$�� �iP{�GU܅kS�E#iL���6p�����-&:�)�3�#����&6u=1�Yw�(F�syAl���,ww	��＝z�ՠ��iA��2��R�u7}Z���o�g\�R�k�͙^���jya��m�_FQ��Cj�n{�M�@2����g'�M^��,g8�(��˲H�/���t�UCH��<�����]�=AǾԀK�V{#a�㻅���w�n�Z�_]QŖ��	mN��B���a@�\Ӹ�]$��3w�`52@����:]nZ�}QX�|�˭Yl�e�\�+Qɻ�J�yV�D�N�1)gN�4�K�|O;�ԼR�{q��J��`�1q���{��,�;�e�T�o'՝1%J)H��*!��}yS�j��N1���"�y'5�l��|�K�F�O�Jq�G-�n���fv.�ܶ*'����a�ɓ�K"���'9��1�z��w2^9��;>8�������^�~�<z2�׀,z���>\�D��R`F�u̩Y'�sF�
32���S?X:1YV�)�S�~�IM�Y;7Φ`T*���p�u���M�<�E&�1TL�p����Tc�E��,��_(�TGRWltV�JR�g��ȉR���ڞ[��}6��\�����<�%�VVz�`#̙/���!�9{ǫz�{�z�����9�n.�ê�18�x�ݠ�\�T��Y,.B'��*eb)�Sr^��b�Ղ���ȴ�P�f�t�f�j�!áׁ�A��Ou�{i���<��!K3�� +_֫��+�ʖ�]\ԗ}NzST�
���υ�4�q���6����>����Ǜ$���
��ZT���Ta��*�,��qy�PFF�N�d��nV�u���ar�W���ʬ���W��6�TV�%"�1^S�;kߞ-�S�$�q�j�%�Ѩ�{Kc]K�B�v��{b��nJ�Ȟ�!j�!�ݬ>��Tz�
ч���(zV�,�Rl�Y�d1�J����?��"k|��a��Yo�؊��F���b�2m�C���ܭX�V�}[�)S��7]��!��X��F<�;����X��o�Mt��"P���Kqe���#�8�B5��{+e�L����o�����&f��C|bsӵ�h��4�ಊ��:�M��w��N}��y�Y�X�֙Kk�h:}*�}ʉ+�B��@��F�^��J�x������[���Lu�Y���VՐ3�zV?���:�y���>�tq�b�i�[�zf�
�-/�����D�I�A���0,;U�U�s��ș�ǉm����WU5V*Յ�����y�󜚌P���GMƏJ�C>��"5�,1c�U���cU0+I�D�fh��tkW:ƈ�/��TEz���y皕�@���6P8,5k�kY�PP��=��y���=�jvM坊�g9{_ 
��׵Q�畒���[�Kχ��d�I��P��_SG#t7���f3��fI��ه`N���Àsp�p���=d*��)��%�yX����|��6;zd�|�=��+B`��Y�-�0[�m
�z�omJ^��g��4F��T����g�oʤeS�P�ߨ��Y���*�Uk�*��C�*ٺݢ`���H��^����Ǐ�Q��/�Q����r��jh�iG%�s2t����ʇ��������bi]hh.+���s�h�Y���e{zd�����q���S\�x���0�S�d���/�V��ʧڗg�"\ܾ�>y&��Π�6drX��Kx��dA&�e���{Pu�ڣA��6�Tq�w��/�$��	FxbL�.v��8��u+�.a����#��&*"V���q�UC���K���fAZ�fq_|���Hn���;�Tc��*g���!�,��悚S�ѨF�tq�āc[J/RoK�l��Ս��ok�ry^L'ԥ�a���Y#�� }�{k*[U��9���7��o�r�M)�������*L^�b}x�S����czw��t�����U�b�Ev��V��x:�uY�`4��})`#ܳ���>�ioJ|�s���Ue\[�}[]��������(7Z|i��	��{Ncb�[q^�Q��I���}!�/h��rQLc�J���1��U	�w�\a0h6�L&��r�J�p`y3��΍���ӌ]7e)�]{y�T
+��[O�� ���G��+8)|�܎��iv��wt��{�����u��m�Q�^� H�_�w�{Rˊ�`��q��-����Bvg:\�E��3gM�)>��8ɥ�e+�+y�ˉ�H�k���vH҉X^�w.`�����Jy��0���c�{]>�,��Wr�u��kq_\��-�ct*{�3w��089��b��*F	1ϝ����MQ���o�;��7Bx�;�l�8�:���j���vrH�V��]
��d�ݓ�ѯ�6Qey���5R�PIg#�/G������f�Y�	��k~[�g�!��p��!1���7z�'otO<�Z�I3����k��m_���yhX��@nU�u���>�����P��sʅ[57t^��%�1dl�O-�m<E��ւ�Uo�L7�3�&�u����1���w�6�A��+!>[�>2�Bj���j�����7[��dzlҏL�&%�ƘQ6I�Cje2R�oJ�&_us�r��Q�;��������(d �g.Y=7J��OR�y�m^fƚ-v�ĝ�}��N*r7��B���+��M���y�5 �㒤/i������.h���*�D�X�P<���_;�����M�/=�*4?b0�>��`+�&W�_��!o 4uT�È�[ǔܿ	���;>����ܬo��e��l=s_gR��[������;��4��kI��ߑ��W-�x��τ̒��mrWO+��L]����q�)_����4�L�!)t{&�Zg7	���[�<3��� n�V����L���eYD���n�w��Yx���VR�}��G݂�*��W�A�͛���"{��~��9���J�<˵ӡ�|#�S��|b-)�̹���|���ޭ����s�M}х��u~W���w�j*��F|�����ՠb���V+�'j�4����et��ҩ;ç���S=��]pn)�}P�Vd����1Zܕݛ�į)�a��,���J�6/ wˉl�ca�d@�k:͜�N;�1>�Rw�]�o0?%y��9�[X@2*"�&*';�0���'��d�L	�?a���%N��l�Qg[�`
i��`*��ߘx2�1^�^U5�:αk<��/ǻ#�Qd~���hv�����a�ծ�머[�N42{�hld��^Δ+a}ʅL�u�x��#���d�	�Ȯ���7�rV��`�}J�?�s&:�]��෎2����V�v�e�������_w��1�(xW��0+�|���B\�5aVz�`#̙���Y� ���y�vb;�X1���uw]���+E�ZP��EN���Cpi��m�\5�&��7��Ιo�����&Z=�3���Wa�%�&$���w0��Wg�.Bhv��D�V��)�n��b���tn�Z�vv��/�D�D��3�Pxnpf:T�MB��پ��yQ�#Et��S�g�%��>1r^q��o;�1}�h�������tfN��Gm��UF?��p8���F��_
A͠f3�.z1�-9i���w@c�ԗ7sn����P��v�H��u�@��y���λΌ�p���[����f�Źǳ{��@9zj��y�bR���ұ�Po�]N����	��Y�6,��[;*�Ƕ�P��!������P������Lw��w��[s޻L�Or�F0�D�v;�A����0�vڜ���~>H��3�Ҍ���̨|6�ξ�6FiW���e�u�kH�Y��\�r�!�tV{ïȒ6��`�m�Ӱ>&坷��]���GnE�@��Y��k�0�/�]Kյ��Tk�W/t,�._y��,>�s�T���Y�"��b�TA9�%�*��OEc6��u���.�Ԧ�i�O��96����<)
0�9�3���3�c�o��>�m��]�W��@f3v�����+T+�OU��}]U�4�"�e�]�u���#N�a!�[�ˁ[���xn^�����{=`0d���&�1�ަ�fT��2*���l�[���8q��rk0�}s�����L�f�wG0ow��E��˯��hߝ�3Ȥ{(C ����׬�*��&7h��7)aq0���'���ޮ�\?m)�Ub��Xˉ��u��#P/uHmgԭp�I��k��ڦ;_du���wVN5'�L�0���^��d����G�ɦ�V�\�F6y��zU/q�K�w>4&6^��#�$e�b���7��	/�:z�Y�D�˪��F��^�������9�6����¾�E����
@�o_\�He�`�Ú|JDc3�v���ւ�C�A.v&~VN�\��`���Y�vyX���C�/B�q��ͦ��g��p�d�O=�M�u�έ�����3m�9oy�dPα�O����{�_��d����r�s
M��#�К��ji��Ҳ�'|m�C��<=���s5d�)[�����Y�l�2ҥ0u9J�Q�B�S=.y!Jht�O�s�c���H�Z�+���x�;'�n��ح6�!W���}JZ��}"�w#\	<ן 'V#~P�]�W���꾥��DZ�6y��yv2*a�2<�iv���E(�����#����%�I_4�[�0�Pr��9�pt�fh}�v���S�f����Z�+T�o�����xd���XsV^)���h���.Y\�kc���*�T��~�ge܃���om黤?P�}j�4�y0���&/q�/
u;��i��Q�G����,���M��$,���"|1}�?.8���+���WŌ���GK�����oϞ�k�9G8Q���
���olTBd�z\��+n"�����I������sP�[W=}<�C����"�\됮u�L�N��|jM�����f�6x���.5�s���d[ݕ��#�m�)G�%Ɇɇ6�����Fi*Ȁ�u}gӫ{1i��ߍ�7S��?�<��1��y��(��Cr/C_D�`��gΏ��: ��CBH���Q;�/�f�U�K?b����|�8:�k��s&�d�iCe���ř���;�T�u�����7���;����9�Mɏh��5�T�<�H�M�EK���C�{��~����o����k��`�`˷�α�'%V_���'%��q���U?o,��o0�o3�՞ւp�Eo�L7L��uV�����m�"�ӋQ��s��qp��*V��Uه�-*}}�k=Ly;��4�1�4Rr'�OC��dr�1O@��@f��U�J���m�� yx6��L�z�Ú��)ѝn�T�������S�S��CW�����aK��sO
4چ>�NC����	�f�Y�swlo!�����ALwCDCX�u_��sr�Yy�����p�`�d���Z�;�7�I<:_I���|z����z(25�����޲��K��+����2i���bO� �9H\#g��=6�/��\Ԃ��ˋ%����ߧ&��P�q��\%"������fe$�+C���1Q�Rٝ��Fgqlc����n��P%.�Ŝl[(u�O��n�pЄ�wJˬ[�He��Ơ;(�]/z��n���xa;�EC��{�b���O���X�5W*l�.B�M��B�������W�ʏ��"ʾ�4�-=Ql��:G�΅n(5Qc�2	��!�t�=�:�\n}��%�OB�rgc��ԄɇJ�H�t�R:���]�<(�kV)��ɷ��\��꺛$������Ŗ v_���1<B����1V�E�j��M��c�n.:���ʗ�w;�����&�[��܎��MR��D���7b��%D��U�^�����vެ�g�:�RU��
������*�˴R֖�ܛ[��8�����\o��;!�g%^9J�,+���{��:���Q���E��9rR�j���Y��Wg<@=�a����5r�#�#�X-���m���k�;u9u���-�S��g�ĕ�r�+��I\Э�Cn@滣�ʰ�o�8iõ}���&�j�vfq���J���+��4X���X�	ּ$A`�;�[X��Н5YR� �,��V�Wv�d����#K�mVlw҂Un�b�n�Ki�mabX!X$2�@�2�u�3��ؓ#t�eAY��;�uӝf�����-0k@���7i��]{��J82�SR����k,YWw�J�'!�/
7V&�ԙ�.��ƗE;��C#:$��G�bT6�G��f�TW@�����d;�\Ŕ��q�75�<�S�g(�Y�E]s�/$	���s�3Y�]�v<��N'kf�=P��зSg3�n�)���w:懫�8�����:��{VL4��6�.����;����8`��ގ��wk�jJ�Ȳ�Fn�;'V���gJ �ж,���g#,hTv����X�Uj�f-U4�@>ؚٕ
��w3�v&}o@.�K�΋��)���$;�3�k���>�/x�]H����5Wz���N�w�.�<�zS�\�[YҲ��+.ȡ�ޢ,�2�z��,r�V�s%��Wdu[��ÈpӸ�7�h�:Z�\�c�sOK�P����u�WK�/.�+����k���P�����Y��_n�.U�1m��2`��b�a�5�f?��h�>�ڍM�P�c�C��:;�N;�Eu`d�����o�����ߛqRN�n����q�����=�C���ӝ��ZXUUW
�W�l��"��c�\�*k��m�e1@�u���+��+��\��n�}FP�\�sNw5�z�&�¨4/99�t劼�Ǩ��;sr�}sFhJ�YO��xh�(ۧ�m�J�w!*J�>ZP���u�l�*e$0�]:�^�l�����ar������d޹XFl�D��B�Wc���U9��ZI�s����8�-�� R��w7F�S������`̴�o�WK�����]� ��(�ӗMa���$[�/Ǉ�`��*�e˔�`<Ő�S@d)���cwvv��U��'Vڃd��p���Jwk�{v�$�i��YA�j�J�Z{Vn����x�[P�0uEt����3�NB�P�Ԍ��v��iPT�q��;\�xpFBvmr�
)�#�Y��g5��i��s��	X��pV�pם�z��3�ѥT�N����S�Av�6��Q��][� ^�����g����O+#׎V��?���ݲ�e�F�fڤ�G�N칵�ht�`��Z�}��Wiԑ��ӷe�L�&B�6�$�t���/lA��/���oTi���Y�|���\�W�6�]],�ZS�ۦ�rO���y��aJ��p�1!���B���d˖�Z�Z+U�ʭZQJ""�-�bܥq�Tb¸[0\���A�j�}�amm4�㙎Z��mU
���d��ln8�j¢�S�p���`�Ǝe��n2�s,�*7Y1�Q-�\-�1��3�D�0�19LQ���1˂LqC"c.�EQbR�����2�m2��*�ʙmej�K����m��T��\AE�[���TDP�p��
���J�1��-
����.\�(��0�\�L�R�FTiq����n*b�1�UŶH�*�[��	��Jʕ�jZ�%T
1��8��"���QJ��--Q*�U1�\̅�c��5QKZ��KKm�fdl
���]YX9kP�[s1�2�1�1XۍJ������Q*,
H����*�l�3 �k\�\�u�1��;��7�5):�4�m�j�O�M��sR�Q��Q��uL��澴�Zff��)r5{z�}�M���u^���ȴFm$���T�b��7ս�~^�~�={T�x��U���p"$���j�6��䧈��cz������������P�d��sxK^�7�oOQ��5��;
k̪�u�HPc����v�t}�؛���3�p��`��U�k�5ٍ������z^�<Φu\#S�P���{&{�'�Z�>&�*�[��S��I��e�w޽�"sԾ����h.w���	�9�i^��1���5C&�0t�Z�����ؖ���c=)���Z�Y�A<��ZW(tr�(���6,y5Ys������qrZ�=�z��'�G�!�n +]��҃��]�T��r߹�=�V�
�}�,�^븭��z����6B
������pYw�n =��4)T;���|�����7d��eNG&�37[��ӿU�r��t�<�(��F3��8�P2�Y�Rb����s���O��sb��&?���:z*�r����.6x��1����
�������|��R��"�����iC����ݡ���B[07Ԃ������GUq�V��1+���U�w���̴�����YI]tH50j޵*;ͦ�V�X���.��zj��AV�=�(pi�ME���+boo]H�_ay
 >B�LO�����P{��i8qXs��OchvG�����?!^��W���Ț�-�^%+�D�Ԇ����ȎRV�h���[��w{猎�o�ua��F�J^������UEqY%D�5�Vwޕ��{ɰ��� ����XX>�{h���3�KC�/�wt�V�ጎ���[ͪoꥢ0�KO��G�*��5��)�Vzʠ���eL�:u��c@�9��̽�J�
}���dÇ�Lu꣨@�#�ȴh�o%S��Ĥk�_��r����g�zI��9�E�6^hj�m����}Ԧkˌ	r����u��F�i���K`�Ş�ذz� ����s����eD��.��d��ȉ�zS��Q3P^F��3�MV
���+�{ӓA�����7[C#r���ie��% ���1@y�B4�*s3P����g$P�n4b2 ���2_�nC��`~��K�����y�iep��Z�b�.+��'��>�o�M^w�F�޷�5�NJ_�U��jAJ�V�<M��zV/ �V_�
e0!�X@�x�� �Al�]{W����M�`G�P�2X���'*���:�ʉɯD U�iT�/+���6�=�H�nq�t:u�z�$��Z�P�A���s�%��斩�����y���wIy856=���ies���Ǡ���w5x�;k9���Ԝ.�.?�NxѾ26]��ú��u�c��)����@{�? �w�ߜ�3��˷�ؗZB/CUO��M��f��T�5�m��_)�C'\��*��ަ%WJ����FT��s�1�2}���=NR�F��*eK����z�{�l��!rc�h�a���j��>I
�:�@�c}����:lU�W�	�)k�#�d55��r }��I��o{�`�[{��ۥ��Li�
-��u��R����W���ELagæ]��2��&OY]/�/�4w, ~���� �b��>��2��O�����f�rw�T�(�R��Zm%���yn��;���b�Љn�0�FD>'�t��R�}Pg�\�\�c*�Y�S�oM���x��t��ʉ�3�t<�WGMH1��B���A�3|<�F�p2��d�^o�����6n�׾��Ւ6�iK1%Ɇɇ7�Ve��i�ܬ�A�_�S��3�s֫:�)]^h��s/���
��#h�^�>apGkˑ"�繟:=D�1�
)�*}[s�7F�����L3����o�D";�]�)2Km]f�2
r[�;��Fo9r@}|(�X \Os���%��z0l����Esgw�YnZX�������1��kyf]�nS�q�`ΰ����#R����L��q�so��l���\�T0�D�ZQ�R,�m���u3�c�+���0��h
%�10�{P�7Y��n"w�9L�^&�}8s��Tp� ̯36�O�+��²:�7�p�{�e�V1�)P(*w�s��jCW�h��_���e�*h�'~�k����@ꬑ��*Y�z\�B����$Ao
��Z�G�_(ՓeA�{1ҟo��{|�><l��K��c�ZY��;<-`��yb�ܭm����Ra��z��|2!����n�����2=*�|���Z��.�<�eaI9�vX��~���M�=��75��Ö���Ε�\w���Z�\<��K��i1ȶ��l9�\ӈ:`�1/��P�U��1V��b�>w���M��0�:7����V�\�y�8 |3]���S��p(���;�V�_}�ërG@Oo���Tl�}uxk)�:��͡`pH*�2�c�1��EK�~5^J�MOJ�����R�6�#��T��R}3�R�KYN��/-���0�Ø=��#Ur��A&c yy��ql��-hV�i��.�g����,vwSO%m��c%��u c���3�J��6f0�u�~Ql��DV�m�3�՞�:�nn�S��J��oݵ(Axܡ��x�NQ\�G2�3met:��B�Ѥh)��-�d�-i�U�oTo�qY��YB�T,�g��/Kh��<��ߧ���9����eQ�fE	����S9'�i�{��s�E_]HSއJ�H�t�&G_[d�]W_����>�
Ѱ�б%��w�a�W沍��2&6x�s~�N1���#L锬 ��ͼ�[{�ݟ����^�y�U�9X�g�D˨�0&���_�]��mS{��b��c��#�����tbI��W����<�&s��y���E�)��w.���(��u����+���/���ʌk;��f��F�����E�S�*�]�Ë�5w2�z�n<�y�w�!b�VoP&}6+����I�\j��r%�\���P)aj�v�{y�x�.oj�E��'%}<�Ɏ�D�N�X]����E��zR��2Z�U��ܑ���b΁ޯ8�}�HX68ӝc!�.VmA�W���gx�dюyJ����wK8����y��rS\(iY��h��<�=�3�\��|�&�(��2x�+�L)��\mf=Z��;V���F&���qu��9��V�4G��54_$;�{t����*�O�J�'�����{��sZ���qu�ނU�z��-m���fՃ�6y7��k5�h��YX�(g9���>�Gg2��B�'������)A/�֭5~���l)��>�
���TޔvyRϵwr9��62�N;\q�'*Wu)RWR��~�J�1+LgdK%�����0�L�zjc+�����p��Q��Q�.!6?�ýr�8�9�ƚ��^��~��r��g���۳�=K�T����w�2�nTܸܨ3hr�Z������r����.�g�<c�Π�d��WC�ý:�y:�����PU8|�z�9V��ت�u3_5{�L/�􉙅k��3��<�f�Z�r:f.���Ǔ�"k����XN�G�}�R��ۊ�cSN-384I9��Ms���պ���=�1�8-Ѯ�_Z';�(`2�Á)H�u2f<�Uǲ,���b��Q�!���:2&K,��N�V���*�-��=�2ؽ�h�p"��}��uv��$t�BFL;���1�E�4Ț�=3o��5���7D�Eyѽ�N/Y��ŷ���T7B�*s+����e��3�գP/u�鍡�6�Ue��?^ڰ�]�=kb|ܺ䡏�Q���˞���N��c�8��[���h�)��#n�Ծ�`^�Ѧ����t�;���;��8�]N�[����ٕ���{}Ä�����kAw]�n=�Cx Z�Q�bNR�zg>�׺���c��⾝)���\H��j��ՈGQ45	�[�\̊���L>�$Ƴ�Q�g&���(�����H�$�I�nz�=�ُ��pX0�	x��B4�s3���!SG���L�PT��V�MfSm`�g!���������y����؅�>PdՕ�)PM��{�fl�P��_���-��|jk!Wp�u�t"���%�cԳ��szm�$�*f�m߲��3)��^��|}.��wZ��ȖO��]v����K��ϲ0�5"�s�v�]����Bgf5�h,^��=��6Ƹ��.� ���G�oo�XzX4�����xD�=&vLbfd�089I
3��T�	�!e�����&�p�QǢ�>���۔�����SD/�z� q|nq��X����/<�:�y����:,��달{�㯹7X	(� �Õp��z�"������U�H���p�
���2���e��b���x�QVoP����%��8�_u�(��P�Fx>�h-�B��o�����Ϸj����8YYV��o%�
w"���gU%���Y��{��]#-)��VҬ�":ˬ���n2�ٞ���ݦ�t��	�^o
�y�����݈:��;����$�|��1h�-Yϴ'�S�7�E���"�SXJ�
=�8B:��{ķ	|\ي����t[�<kS�(~G�Bj'�3Є=��ف7J.��	�b\����g.oô��s�;�57N�~UpiN��y:` E�fD�[�Z+�tu�<���?w�x�3�Y�G���_y�a�'�<'(ǚ�kL.�t|��gL���onM�M�g�x[���+�QŃ¥ѯ)G�tJxė����V���sh�����k�ݩIs��
����f�a�=��t�^�f�@�Q.���#�	O��T�kӽO���޷ȝ4Q�4;n�Ld��Z0JY��v���j��\R�wZ޵���r���x��W"rqN@��S����ׁ��[����u:3FAU�7iKʭ�'���T��<Bm�h�9��9��L�F�wegR��h �h�G:�n-�:�+=y͇��nnL���㪹��;�J�M��s�(f���y�KzB��4��z�^"�IwUX:���C}��cع(a���×$�4'Oi�~~��O���uȍ|������<y'���]�7֪�X���	^���,�[ocK��d�\���S=�8䬬ʁ�Р�Y����Vs�}�u���]�k#�,}����bt�s�]�';��ɘ�@;0�ߖ�=�r2���1�<�R�J�n�:s
jQ��雓S�ӄ����=Q=����bqW1H9H8fϟK��
f������Zpb���5gޛ8 kܠ�<&���p�&�s����B�}�ánH���b�.vʶDОL�"��-��4=S�0�C����|p G�Ϛ_wJm4 ���߲�ї����}"S����k�:�0�E�E�~Qv$tLp�^č����C]�xh*��X��WJ���Q�o��5��P��(�Zs�`�- {�߁��'P0]���m��8�Wo>�b��~���ϙ�9&>�3�ϻ��m����*�#�4L��~�º۱����I1���WV�g���I����=�1d�IXC�Ӿ���"��Xe��!~�������>����o;[�}�u�*�tB�jZQR\�E��.�G����w��&i>�7c���C�����2�y��ؠKد�,n��c�Z~V-%��[ն�HB��H˝ֈ��@�/W��
d-Q�o�OS�bb��;=�XZ��pJ��t��p{(�s@���Yq��0N9m� i��;�W�)2{����Hһ@�z�f&1F��u�\��f�z�c�;&Np����YZ�00B��3�Ya�hکz򳖮��e�%�7�2�=s���MQ)��1uͰ��o
ڎa��4yKs�w�����a�����	[ҁ6&�t��5�J��>>�V73�0i�7�c���m���L^����Cc'=+�����{&�VR��З&oj���s�6���Qr�ƘR%�/"���*g�P��o�9����ǋ��N]m闚p���$��q��P˖���Cv<i�O�
&����Hk
L��'��ӥ���쮢[�����d�ea�-��tP�,��/ȑ�-�,
ޠH�=�d��Y��me�s�VP2��.T�[E�l�S�@Bڋ�K9��Q-�	��,��P����+hP�}�\ՈiQ�5��w
n'VTtߋ�@��aD��W�.�1 w\��sy�Q-�ҩZ��NɌUM�HU�V���Jay�m�Ʀ�p2TĢ��V\NѾ`�k�3��}�2� 9�+FV�;M���el��������of�݇�e�0��\��ɽ 
L��۲��خ�v���ά4��(֩K�Ք����=z�<`v%���ٜŔ�$�#�3���m��;���i���T�N��kd�@V��2;�T+;c��7aPd�b�ٝv2�-�&��v츲�]iXo7R0euv�ƷLLn��"`��gy�^P���.�]�Ռ@���Ŋ�^��;��*\��J��DLшÄV�2�Pj����#O��e<]�N�����ޮ��5E׷Nq�r�֧ .�!�%�yJ4m��i����A�;��ǃ����#
�z�*�Ve�E��ߍ���xzf�D0�z����iKɮl�V�+���ꂎ�-�U�\�V�7)��W3�9��!rF��%У�\�y�^N�ac=��5b����a�	�M�"[�el84ǀ����U��N�� �D�{��f�N�
�Z�����[V����b�Մ��c���v]�.����c)lSr�<��`��/i�_ �Ҽ��vR���]��NG\f^���_V_0�:�es��*e�k�}o#{/�NBb�7W{M��D8�@�������]r�E�2۶n�Q��x�Е\�=���Y���pҥ�b�l<]�x�ŭ��@�`;�*\���l�͉|�����u*��������W�Wn�[��;�١I��p˜�������;Li�8�]�7�鳣#ww�k6�]�	������ӃV<б-����JX��1��]np9������FT�#�cZ�#��+�cغI{���p�ۼ���C�7�/�حjU����}�C*v�G�Wc��c��/ٟZ���ͫ�4gt^�S�uجJͧ!�cF��o���.D��Ȣ���9>���[��b�J�B�2;(
�sA���fG����2;X���i��E�WLVM������&9q�c�iW$5�{�Y�:Zz���x(�s�q[*���{W���]�p����.�i=���פjd�c;�E�Fژ�h8���@�0񕅻|M�.��T;��(�v~���8�3`Cx�N�j�2���/:�7@���x�v&aS�q��_>JH\���U|�d��1-���Wn�@T;VyV���f�XC�mɼ���U�ڧzr��O��eݍ����RԼp��\�x��v^�E��f4�@LK��<#��(��*�˃j^�������{v�
����o
��\'���/s�\i���5i���M�9�r��v�wu��$c�ۨ���lG��E�2�_-�i�LZ�lXv���p��S^� ��r��T/y;3-�.?�U0���L�H���ECvu�Q��]�#C׫lr���2��M,m�.���]��zJ+(@Sj�5\N��T�"�u kk��J��B����!h!��RZ�ٙr�8X{i�M�0��`9�jM5/cW�����b�V�,�gJ��JՑ$pie`�5ݽ�QG��� �ul�u!� ���ۻ/��=��9���xUo5�1Ԏ��n������H�Lmh��־���g����̬��M�Vq��UYU�(���*QK[RȢ�,�-hԪ��,5����Ƙ6�Q��`�PZ+d���-n��Q
�ec0e�`5�
��"�q�V�b,X`��ӎ%J�ŬQ�b��s.*1aX���FAh�VTm�.Z�Զ��P�m��-��j6�2�Xb��Q�m-�q�m�1m���S�rܲ�mQ�����uL2Զ6�JԺ��"Ԩ�ڢ�j嶭kU���
Z�YY�m+�F�����ʃF�j��q�ZE�ʔV�[CL�]&`�+m��b�Y1
��-�K�TKd��̥�1P�*Ŷ����,���e���P��Umj��B�0�mnR�pUՔM[��U�6V�����˕ib�R."#hU-��cK3*.*�TF-*����bVbZ�ڪ�Q��))mnfckG�TQ(�M����m�Y�_[sF�]��&�"�H����M�]]p�3s�\��Ntu�]�=}��ٓ��I��Gpb��-pr'TҺd�')�Jb�J��ɒ�x�Ϗb>1�Xl]���Nw��C<
���>��eR�wV��dj�����,�G��u�i�YFJ,�ߍ8C>��T<r�-�������WⳜm�mi�4T�q!LV�&�tu�
��:<��MA��*�^5�hKW��hX]Yw��e�e�z�k�t:�MY�ħU��.�Dx:��r&��f����j*z����e��˷�s���aO�
�Rj�5�䑱�ɏý	)��'�XT�GI9^��7ͅ6�ut�
j��l���Y�5�q���5 ���C�T
4揕9����s���v>~0��o:�w0: �ô-m�8m,�p�o<:���J��}�~
O/[�;���L�nis�Ҭ�=bf���5�|˱�u7���~VOL^U��� ��ԻG3*�$ͮҪ�Ժ���e
;�۷�>=�H�ɾb7�7��j�S&pP��C�n���s��ˌ�����꤂�B&���}7��@==��.юx\Uᔣ+Ԋ����X�9ь�t�gk+�� �H��V�.����������ҽ�>-W��o��Y-N����#�6�6��Z��Q��S�y��+�[�n�k6!į�v<��Dt�6\���$J���e(�[�.I.��:�j�ͧS6:��p���:R��Ɛ�"�sB��oB��>@b�G�����p]C �a!�)���c��`�C�⥹U�M�rc�1����*Aڌ�:EL��c�+����>����X���f�E��0��Rە��u��띗���Uj�Jҋ�L�&�8�G�j�>�QA�e`�Vs;����7�-�;��j�T�ּs��eTB�`�Ɓ��W�{��5s#^=�L^��=d`��{m�:�.N��T����s����}N�p������7�:` E�f\Ԡ���$��zucF�����fg%+A��$l/B K����U�eO��rz���ɋ�r_���0m_c�Ɏ�O"��9��y��%0�$�D�H��'G����\���[�8?x���-�� w���{1��9j��dN��l��ADÉ�ي�r;YNf�j3GS]w�Q�vy�4(��^fm�S��0="�w�V�1����4a�=5bG�y��ԯ\�][���R�����bu�z�K�h���1�	P�~�qp��������w�ĕI�@��٬�쾼Bw>�c�+����E1����paF�' �nt�U�d���v�	SXCG7-.�Œ=�A�H�kk�$���w:��l�	^}�謡+=����㮇����a�+� ���U�wk�F��a�οj�'\�<���&�j*�,y7�銾gEQ���Å�+��ɆI��d��O}�{"@kӳ8(aB��4�K�����kWR~�o1x;	GH@�Zٛ����NǸB7i�yP3q��:6=��75��×$�4Ε�v�*쥹��K���f߻�n�|}�:0\ބ�R���;`�r1&1b�S�ųg�rt�/��+rs/���v��ܗ���}��nh=�ǯ�P���\"hw/�۩��%��T��v�j&x{�}��k����zT�b���	Ҡ�\��OW1��T��U�	����;N���`�vv�n�|gv��dpZg��<4��p�/�hD�~ta��0'Gqz2+:6�0n���z��׺{r�A�S,Xt��	��Pݬ�z/�B� �yi�������m[���y�p��H����-�у�[��:��ã���3�^Ϧ�"�I�A�+����9�76��b��9ǜUĐ�QEOk	� �
9ܠKq���{���J/��<�^f��֌��Ŕ�^M�ѷ\�u�WMk��P��¹>[�f�Z�Kn.����O9�h��KV˕Ș�s9�Z����kV��:�ST�`#��5v����[��v�V���ݐ;��]	�)�[�Z�����=�1e������;��ܓ�:�F�O3j��{�h}Xfx� y��,t'��yتݫ�+���,��bBy�z���R�Xy��eD�|l<��3���ekmC���"�=�#P��z^��qg:�� �/�7Z�����������{��O4;1�M!��S:�6��|��3f��v��͹���nk��5���Cc$&9�V��Lث���bo�rT�+�p�\+�*��eto.�꨸��P�`�i��㪞��:��l��W���i�ɭ�3��S���V�4��T�YD��u0#���ٸ��Q9oL+��i�-���\��F
W~��h]����5w!M���rH���Jj���xP����ð�y=��S�"�y7��T�+d絽S�%O>N�oBѳ�i�D�zw=.��o�����˺dK��9�z"2�=���/�k�*����tf^�59����:T�Zc;%���G�'�&[ˉ��$e��gACS����U����.b8�ݾ`,	t��yM�O���3��`c)�=+˾���������@�!�̀q2���L��#��p��'is�͊�_F�J��`:T)>����}�˫�jcP�z�ݔݹn'H�gD���Zܺ��y�js���N���xw��R� �[\]@l�0�g��q#{�K�X�d�k�EF��������S�qR�gJ0��G�\nqx�<Aa愇��o�3���T4��TfzbeytZ*�I���膆`�X;WSr�:�3!G�s���	�Sw��e�W�$u!���ŝo|���B����C��V�B�iA��k.����申�{m�Xq��b+$��,�d�^'��lǑa`���&��P��;�+��Y�6���]K�z����!���2Yd�p�B�Ԙ>�<iչ�7�7R��.�q�]���g�^ɈW�Jl�m�� r9l��h�o"j���̢<����)sr��S���H�1ܷ�:LnѠu���3K�	r�����u�+��{�����{��.d���;�7V6�a��X�QF��
����]g <��������h�)ִy/k���Lv�)#w�?w�j���P�m�;�j��������Pk���צ������c�w`Y5��pѽ�,�:�t�F0�a�aN�͓L��L�Hb�ϐ�s��_{��ٜ�vL�
�;�yYR�l��� m����3Z�:_q��n>���LTl'BP�m.���Iv�S]�2���mv>�5�v$67[�W�яpiM�5{�$��ws3�d*N��ׅ����xv�0<��<ᴲ��`[����!٢�����0�R�����0u�3���}W<J�*�^{Z
��[���4�?+'�b�ȟ��Y+�����}{��]�x���1\�����6X�_\��Ӏդdꌽ�d����h]�vF-z5
MB�v�Lֿiٚ���&O�F�z� �7/�9�*�}����%p���'x0��Ć���t[bj��^i�֎���D˓��1���>�r�£s�b�T�La���wV7g4�Ӆ�J�Қ�*P��W*�'|n��q�W�&61�b�+����t�̩ݵQ�'�n���X��V���W�a���TɉڎQ���F��+�t��IX��,�7����7d���9�9�^��5�w1}�bQL(�9�Ŀ�9����j�>�:3k��t��7­WR�3�o{9P�l�v9�^����*�:`�Ɓ��G�&�|�=XJY��G��Qw������ކς�싁���\Y�~�P�Cϕ�:jK�'~����~���f����1QWnJ�׵�G�.�ҩQY:��l���wy�:\�z������^��b�L��k)�Lu�R��\B��T4D�3+z���5�٥�nt�e�ի;.�t��5�kS�,#�� ���fb�2�,�N��1�8��v���C�h}�frQ��zY#niK0\�l�sj��5Y�C�r����z��Jں�����<���Oi,�$�
ʺ5ʤm� GD�\I�Ƚ	����[�����Y�B�^�q�L��Tga�cz��*�N/Y�{;E�a�G^�yM�U��S��z���Ičh�Sr&3�y��S��0=8h<�\[Jў�%*���b�$�[�ZW���:8(�@؛)�g%��K�z��*��0�KvZ�n�j�!�ޣ��\�R����)\P���V+�v�f��I�{Z?�P�I�a��������uU��qv����R�������*�c�'f_ήTF5ݑ��;�����.���oϠ�l1�]���GU�Y�����;ţ�����.IV}�M�K�NH�/�TF\ǅ����py�	r���Cp��z��|��EN[s�<v�wn���l�ZH^�SRw���*W��Y�L�o�#��{���[(Q���S��Yn�x�X����1�2Q;��*T��W^:=����vf�^R�VgBy�ۛj1��#e�w��,���tѭE �a3��`5�2k;��xuN���e`z�F�Y����)��aw�Ǯr=�8j	�[.�| V�[�PbO)G46�}صu�kv��*i��<T�":^ @��u �)�3s��l�/��y+�[EE��'��ݣ̬[u7&rj]�W��ɺ��xi���Gc@�D��װ	wi�g��Na�S���*�5W:#,x?���q��������3�t,�-�{���Gݹ��գ���:�Y�@��Z��ͫ����Y�X��ׄO��y�xFѱL��W�K�MF�>��i����y�og����Ț����=�Y%)+��E��orK�4)���,��}���_��c�3(�A#�w�i�`{T���WT�_y^=��0�Yl��~<b/ntq��<��C��c��ȸ�MK��5:e���^�}��Z� � vQO35W������㩑RR��+������\�y�4=�
c�CՆ��t���vv�L�x��$[�.v��7��N�4HX9�V��M��]��o܅;�h�㎅o��y\�.\\��&&ΘHi��㪞���S:�	��+�O�L�/�ѭ�喱
�b���NA�[�������>�O�.�V��\	�%�gV�[��U�/��Ԯب{%7s���� ��*Y��9�pĨ�=K/� �GD4A��f���A�0�9�gd95TE��g2�1��Q�VؕǦIՓD��Rw���%Β_���0�jRWO�T����XӖ�>%���ȭ����//KڢSz�l��wE5Y��G4j�\�T���4歍��W�q
Kڠ�޷�����,dúC
{r׫��l�T �صh��X.�V���a�@V�\3[Y��[+&s��t��b;�E�iU�5r�s
T[E�l�:S&"V��ȖK8Y9�NS�E���&�n�5b�ˬ��]���!;��y�ް9Jh�cf�]* ��0�r�)'}Զ���t������6��_ѡ��i�˸�k8�zzSn�榴�S���ܨ=��ɱ�����]��G��eC�7R.�M��h_FV��x���Np��F�+�}Y˼�٥�[C�$�c�a"H�Xŝ��v�V`�^�Q��P��8�����g̪؜��.(w�B !t�A�dA˅���v��}3���{�����g+t}`�R��-��R���!Gc�*��*׉�"�PVz��۷}ک+5���8K��Dv�W�h�d�[�Ź�-��Ƈ��8 x?gV���9��4�m������w���[8>�n#�!���w���|n�v)FN MYxё����+�i�Q�,ō�/\��{Ҵ&�(�F���;w/6��hb8�T��yv���A��?b���ƣ&�GX���["�4�g�:U(<v5�/!H79R9�(�2&��3����N�ک�H9��\�|F]_|��ۈ7�u�yܹ�>�����t�ʠwN��eRj��P�:�6�r&<�BJc�Q9t��"�����9�.P��Ji6��y&�f+}W�K��B�Rׅ��:�2׆(4�;�q���r'�����i�R����L�������kDXt@��p���������F Xw�b�{�v̮չ�@\WO��\�#��L��Ʋke�ǸU�vo�1`._*�j�B.�%-33,�li�K9��dva�6��b�F˺�+����?_�X����J�S�j�{vwv�uu�z�;��z����d�I���|��)V����ЎDGY޻��S���'NMZ|m���~N��q)mT���eF:s �9J�Q��1S*]dm��dN@�r��eohD[���}���hU���0�a d!����qȝ}o���um�U[X�"����|oT=�sf� �u�Zj	:J�+T���wk��kՔ3�t,4U���r�������텄Ml�`�>�U�k2��<2�Ub\E�R�dgk�I|��c�[G�N���'>%K|;�+�&"wک�V����ؖ���8�a��<�u��g�6�\��
��lF��ꙛ����	m2��`c�4�n"�<�9HH�d�C3��m��G6�-p��v������N����y�o^�;#�M5��a��H)����w^���;55�����*2ӥT��h�b�u��/uihn��5.��޶Cy��%i����⮌wDa�����h]]`3��{�"�/�tt���[(μ��6���S�n
��j��S�K�\T9�����s�Gn��k�wF���Ngq��(�|��:<��w��o���_Wy�͜���@S���ܣ�v�;M���SRߴ蛵o�B�؅vՃpW0�GJf�{�͜���D�@�ofoa�C/V��r�@B��ږ5���w�%�u�`	�7H��t�ξSD�RZ���α�O�n�BZ�C(a}W�o ��qre<�%�֖����м�nV���)G��LޣYj�sWS���%dQ�HfVe��k~�>�R�g�Nk|��T5�� ܝ
j�/{�J�m���
��ri,a{ ���"e{�K��b��N��d*����(��<9��j��9����w�10]�Aq֘ P�9zN��C/��˽��tEk]��
�Y8!;(�ά������6)�*^��@�=��X�v��*���1}���u�6��r;�[7�b���5�S��T�=��i=vl��v�$΂�`z�͖��I�å[ݤ'h��0�����n��.�270�5�I�q���p��moW�:�ُ��m��81�)x��d��f�:[��%3�]�I�wr�킌�lJN$__v]�We�lg���ܻ/o���j��YF-�<�ZJ�S��I� �=3+	u�[io�LαX���4����pt�`c�w��;�Ϋ{b!��>0Gt�n�Y.��wGQ|�rT�(�v�����H��7A��tx�x�ހ�'z��s{��FJue��V���u�y�ƺ^<�gK���Z�ݦYr��9M�Ù�
ƫ���Sqc�a�.xO.*�Y�tf����¤=�sGwFa��;�p^�y��t�]�b#.�*������Ln�N�����XT��w��ti��ӧ���t��V��)Q�X��]��Mn�Q�'�vY	��X+�e�h��#m��ދ-8q����GM�S�YӍoŠ�t��pK��5�䈧ol��5O���� i��&ޫǲ�wx}��zfJ!�w(�^-���Y���"�Q�_X���e<�kWX+�� ̥�CE�r-�����K�x�GS���nVӷ�d���5W���u�j1��G��ֿ}��b���P���uQ��\h)�`�n�
�E�U��,-jխ�1(ۃ��""�Z�U�+[h�U*�SN(��ikF�Z�(���J��hU,J�n4r�e��(֪6���m����Q����6�ulm)����F�VFJ(�R�-e�DmQ%B�V1�жʖ�Q-iQ�A�����#YF*�(�F�YQ媍J��I�b�2U�Q"�����d]j��ӧCij�MTQD�e�-
)�X��5�й�EC�m��F+q��kj�F-�kE��Ī)R��8ܲ�h�b��ڢ��Yq�ekXV����KbQZZ-��e���8�unE��Z*
[h��l�T�h�V�5+R��(1J�1�T+YZ��K��\h�ʈ��*4m(�Dm�+F�V�iQ�iAEJ�+YkJڔ��"Q*R�������(��"֬AV�YQFT]�*��w�7��t����O��wJ�&k*.%n���2�&�����L��;V��U:fKu��evV!����mӃy7��9Ȼ�%��{Tм+���
J.|M�c�PX_[/lyC��VI�֖D|��n��̚�JsЎQ�#�T��:eV��v��ES&J�!�!��D���� =�z�bz>�76�;]����AI(]�rת=!y�UD,t��Lh(+�=��NoS2x��<v\��ayH���.�^ZB*o��$�GX[!�'v����b.!U��.���܉�Y�_o$��J�<�a�:?{\`X�Tl{��`�RϠ"�-�em�ﷶz^=��{�����kL,�g���ҙ9�YN,0���U6� GD��/�5�����jh��wyvb��R0Il�W
��;}5Fv�q��{QD;�&��h	goX�j���s٩;pV���*��%���]�k����ѡ�1���h�T��L�e�JދW�ԡ��ѼJ�96�qq;].l�i���Xe/��Y;N�t��5�70̒l�8<�u��������UQ�c]N:R%V�y+�v�eo��g������M�Y�+=�����S�V��3�l���=$�~����]/s)Ie��39>B��)Lͥ��I���U�`���:�4�����]�y����ɔDӻ�s@�A�C"Jms�v��H{��WQ�1�^Ҵ�����zb�D�t��s�TNZ�e���TK����T�e>P�����j���k�#��6��-[������=���$;<#��OVyP3hg�����b����R�#���SyS���vaɥW�薭,�{.;��=����,L�ɸu[5J��)���r1'؏1S4�P�9�i7�x^]#�:��g��zm4_ܩP���Y�
f|�s��{���j�Î����}d�O4��`���QXt��*^1Q�����P�9��d�*^���f�z��v�H�c�jp��rf�F3�N0F�,i�����1p��JV����6�c9q���ы�9��o�#,huK��(g��oo�B���OB���$�vW[z��NA�:'O���i\LwS��`\��a��5�$��Z��׊���U�Qy�`����]��;�| W>�@��6��|k���{1�59�8e�GR���ln��<uy��vwa�F�1h?J9]6���u��f��ҼX����&�(֜3�~B��ƥa^�=]PT�1.e(�P�f|�K[y8cr�ej���;�V�z��	�޻c��:��1�.�$ΘzZ���'}������Ԇ:�w����I���\��S��*��T��靨����-�O=�*��d�bo�P�&9k"�ڥ�Kz���=�T=�t1�p��d\q&�#,y{Kg��=�]��)F�d��G��^@}&������~ʰ3�Mv�`.f�D�d�5/�EO�����ʎ�]'"u��OU�c�-o����q����Cc$.P�CzX&lU��g�7��F^�n���^��:�*��*zl8��>�D1�M�<��rO3�c�Q=פ�s����tgf�N��DT[/�3=�)��&uPo��a�����?���_ڟb�7��,��Ȫ[���;�g"(��1r^q��^6���7^��kUl䦼(iuVz���PP�����q���Ny��H7��ư�˝z�ˌuF�AZt�����O���a�����\)�ٕ��9�*e�>��!먣Ԓ��5r�+�Rm��6r)Ҡ�1���cf'���%5�R;�M%Uh�&{��S<��E�T��J��䃸Sq:���˥@a��I��U��kتx���2t��N���q�]c ��o"�J�b*r�$*򳔥��-�qd�c֨������U��;(޽�jUe��iX��BN!�Km�u�F	�pAjt���Ŏ�v��3xe�k,܍V�����r�3d#Y�N;���u�݊�wv�L���fqJ��d��]�7�쇣qT���NY�vn�յ26�֬�6͛��UmQ��F��n�P���"��{�4!9]�=k��{�\�)���ʿa�gv_�����^�@L/�&yGRHoLON֭�����т冎�e�)ǧ$vov9�=~��ǰ�.l�JRޓ��J��Yd�e��=h�<��*�n���4���kn��o�.�����WZh���jP�����qh��zY`kxR��;���b%�twW�-1�4B"�N~ʙ�t�<Ɓ��F�&��:�VY���@��<��Ļ޹�W�w:4tœkƀhm�&rV\a`)1�F�����Nf����'���
P=��2����6��/w9Ơ�:.h,3�Wj±B3��:����M�U2��dTՄ�57������;����(��ɦ�V�\�F6%�j���.�uБ�*yJ���A�sz�g3/��C���ׂ|� �����v^�~mm|cô`yko�K(p�o��}}��m�,+h&5�X!�1�Z���x�%o�b9�H)�9�)���R����L��ޓ�S#J8��N��m�$;�{륕b㫝��d�vy��{��-��c�]���]ݹH`����
U���K��)$�U����2٧�*��:hyq�qLQd�`{(��SoӺ�ߌ�/]����	��/V��YzI}���zhc�� ��o��^���߯����]o�>��k�;�^{H��*R���1מ�=�����n���Ucs5��LL���꤂ȄM��NaJ���ܓ&��9o���WN5��B|o�WHU�ނ.%+�&\�L̜t�\����ҧb����j�H��w�����Y�,T�-|h�����\6B����tج:)�$wqn�YU�׹��x���J��V �FH�ׁ'�s��\$��֪4��\0nT����O_�D�s[[�G�Vi<��Lat�{ֱ(�L,�<M��j4?��,+�mMr��ܸ�ݹ�tSU)���k�ٿ@��3<�� ZK��y�SJW�y�~��z�p�s�)P�@z��<)Qcr*b��7�a��=��L�5;N����5��T��V4����9�=����~�bxJ��������fg%��K#viK!%ȭ�r�ソ�$�Խ��ՃB��P]��(:P�t��b����S�\�m+�O�{�44�w^@��w+�"u��7bĸ��ɪ����Yj�J�s2#��O8^�"�����Z�ym#'�r�]�6�on��7��dB��٨Q|�^O�e��(D��R�V��'J�ޑt\�ƞ�k[�+G�o���.�@�w��g\��wf1���X"����֦��۠�*��Ҷ�-�*L��dJAw��Rlu�[�;Ơ��}�����{#v��F�6f�O�(1ھ�4�1��*=�=t��\eγ�Fs��:���|�X��zCBy|�GF����]�����rv��vmV(=���zf�����
7����3ٵ��y-���C2�3�g.f'�gW/^�����uX�.���{�~�|ڪ�.W�ߓ�/��W*Q�Y�(�QRpv�d��իa8u�Z�H���E�V�fP��u�_k!���I˘��DN�Lg�[y�mR����q�;S�Y������Y=5e(_�Kc~#|�VN�%+ӡ�sh���z+��AQ�-�[.E�,����W��C��ϛ��;�oe$��zm)��[����\�V�F[�:��q�cO��ե��斞���:�,#�f����>I
�$?�v�R�=&L[J�XǽZg��"��7�v4r;���'9��j�L��<ЊVz��^�Xi����L]�QfA�������[95�VɈ��2��Zm[�)vMG��r�[��*�K�LX���>����q�b����;ڵ�8Cm㲲ᦍ�$n:�>R��^��N��4n�Z9η��S�v�z��}��m����45���3���Y�(�P�A����s��9^���&���ܕ��P��q�bxJh����Tf���-tt,}�f!��'�[����W��f,�ȕ1$L�~L����R;�v�� �k��MNuaa��cF���S������c[��
��Q�ES��N1���"�j������zH�P�*ӆ{3��:��vH�~O��坟l�E��--T����(��7G��I�BǗ����ǒVd�|r]����÷�{
�k������*��>���Q��Vhw+G�H{vM�NK�f�S<�u�u�󈝍&++p<�,�~��cvpld���Sޖ	�خ��k^h��b/��9�T��W�71
*mcQ�UaЮdǎ��㏆��9[�^�������G����^��v�:m���߆G��trc)+���V���*vku!z(��Z�v��*q�D�Y���y�tVy3��4j����O��g#^4�=C��Wr>��U��a��/k��=ʖ�KB��a�&�2=�*q�`?S��t���»3��5�℮Y7l�������OϏ�����f�״�H��هx-u���cY��N�	$�8�p0�w�oN��Z����ݻ�J�W�T���T]X�dݭyZ�\���y�B���s�Y��#�d�+N����ΉtP�,��{&A�eR��tj�o���Y#'����19�]EpIW#W/G0�[E�l�W�`W�x����*ݿ]m0���1�Q�0y�w��@w�4)T;�	ܸ-5�2`V����T���9N���w�(T��頻'� �x�D�|�6��c����	S������HU�V���J`�Et��ل<��k�J�����S�fL�}=�h�"�&2.�I���ƈhajά������*�IC�R��)T��)_L�$��4��6�����'�΢:�����\��[f�yZ�8��;L
="�]K�WVPtʨ�謒���&J�ߑ��""Ȭ�d歙k�.v���i�����d���C%)f�xMq���v<⨼Q��x�6(i�{pﹺkop�������T�MX��Д-����D�ŉn�c;��P��"�dJ��%z�����U;J��P��!�n���C:�x���.���O�^v�#��� ��]�s��C3�32�bqr���k��0����ҪE8���S�w��oC=���1K5�޺bԩ&��T���k���Cw[zj��B�V`x%�K��8�ܢ���+M�}z�;����p�~$��YS޾㽱RsrvI�κ��qrp���nf�s31|��'T<�&H�PIC���k�a{�Ll�}���ɪ�es��h���V��WyW��{}�Cw�DR�����B���y����&��xbS�Q�)m��:������M�;$w�/��Q�PPֵ��8Ibl���잲���/ͭ�cô`h�w=d��a���\�a����"[�¶���\U��}s�p�f&o�F�:���\J=®�]Aɾ�w�co�u#�����/�V?�,�ZO_���6X�B�nޑذ��l��o�P��֚]�mZ�̃�"x�"���C��W�.f�)12b8F��$B&��z�/�Ny��F?��.kQGSճv���3�e�nG�.%+�e�����(�^��	7u��_z��Nآkn�pЫ����[.h@�ɋ��\�#�w��q��q_y�:��-������圻mp]�A��KȆ�7^��u�I��s��\$8Z�����㥶��÷��(�Z�qî�X�Gf�B ���{ڷ��J*�]߼˺C�]}\D#W+�ZI9	��i�EQ|ˆ���r����n����a�����e"��ő�U2���I�v������ٺ��V��4�㵭k�ES���hn^�������0�}���]p�mwH��2]�Cp��fˇf�6c�����w�}�m4���rׅG�/>ʨ�����"[�5�ڲ��c��g�gg%�|�Z'�)��,� �sp�೽�-�8|�ښ��E��{f6���!�{9Ϛ9�:�?BUt9g�������|��g���<l�X����/��S�o�cB����'�>�@OK�"aM�ՙMMi�ܬ�A����Y�QŃ¥]�]��I��*��y�<��A���sqT�y�:=D�1�5Fv���c�����**�-l�������L'�D�>��U${�%k��2�+k}���J��c��~T�Wp���K>����yXEj�d�b,Q����C�u����e���Ul]m�l��o��q�F߾���@���VP�C<3��lYȍG�|:�5�Ot�����)ZZ�Y���HY�Ow�MI�s�V�|C�6��L�e>mUs������|;�0��\"�2����O���s��F�R�b��t2��˯o�W��_������u=�7��	!I��$�	'�BB��D$�	%!$ I?�	!I��IO�!$ I?�	!I�$�	'��IO���$�܄��$�	!IHIO�	!I��IO�BH@�bB����$�����$��IOHIO�1AY&SYעyt}�_�rYc��=�]�?���b>�"�JT��J!$R�IIRAP�"��$�U)E*���R�T�@��*��
��IRn�UTE*�ƤJ��QR *�)%BB%JUID$H��-`��P�D"QA%(
$�dB�U(!$��%(%U)*�*� J@��E)R�QJR��H�*P�BJWF��t�*�E|  .:�(T�b���mVkT4ؖʨ���� k5[A�LɀU�@ �6�PI@J���B�  �H蕭���b��%6�Y*���$�5UB	@l�0�@F
��EQ*�&�$T��  q�)�L�R���Kk`�
�L1EMm��4դ�V�EV5�I�[U�@CQ�VڨI�*Q2�RAp ;�
�V���MPf�UZ7(
�p�@P�� ���Р(P��w QCC@(P��0tP : 
˸P��@4.9�P��YIS���JJ��%)T%R�J�8  �R�@̶�3HD35MeJ�l[R�kT��Q��VZ�JQTm�m�UU��T1[	D���kB�Pb��V�KZ�
�*8  �%]5T��6�M�*Im�J�ZT�����UU-��*�M�XcZk�&�j���`թP%L�R)	*V�A�#V�  ��Aj`4�[Ef�Pֶl�m�VX��J�J�b���-��R�U	l�4�UT�ɪUH*���a�1��*�l UQ$R�  �RKJ�j�mJ6��P,��Z�֩Cl� �SbX��5M�V
�2Ѳc5�Q�������ɒ��j�̥QP�BQJB�W  i�J�V�j���d��V����D��D�jP*Y��5��X�UB��� 6*����M(����*-���  .� �SAE3 Pm�(mfk64mF��-�� �ն
U�l SSCy�(  &�R�*A�@�  ��$�)��1  � 昙2h�`��` ���S�A)UOP       DH�&��M5<���54ڍ24d�4�	4�	�)B	�6�!�NGW8��v˞Y�9bԌ�V�e�ئ-6g)/zW�����b
b�-�AS*�����UPz��Aj"* 'TAF�|T+�?3�&B���D0�PF	��# ��P����
L �
7����g�Z�X���׻ F�ȚZY��K�q0w��;n�,�A�C2f5���-�ZIM�l`�FS��� �n
�Y
���w�fd�J�`��]�mL[m�݇Z�TfE[�y3[�˺N�TL�i���+�gL�����ԝ�W��ۭ��V�K�a����J0;zH���l�۳�ꕮ%��B��j�.��m8Bt"���
�?���&�-)]�.V�P+�@�ՇwOM�N�fm�޵���ֹlh�KtƏ�튶�j��ѹ��0m��<��S�b��Tcx�%�c���r�CM������&)�Y��l���f�H�3X��0-�+eaY1�td�֭f�+��6�E��P���5��l�,�Q��b`�#v䩛7P��-eCpZ����ͥKV`͖�@/�-n|�&JhQ9I��5�z�2�tx(��^i(2�yu��ɶ�E�׵l7��蝨�Z���-��u��o(J�(�։�7-�d�Xĭ�knZ��l�)[�b�N숗Z�\l|�`u����,t�ހ��<qf@��f�zTKY��ԛH����Hdw-.�'�Ky�TTm\��8ă6�:#-�RSm�K5�^[�h��X�lUz�4�*A��Z�5)��Px]�2�K���M*�j3�+B�i�[	�����f� �71B���sfGa5&���s1K���v��GN�J��t[R,�����WU��G>8�j�(2ĤZXv@�ӻt�"����~ۏ^d;SU;yH01�]���!e\Zg���cS6!.9��X�a���;�O��U�$]˽{����SJ���V%H���L06���e���3.�������4C�'j��� f.���Y=��#��h_D�¬/cjd� G�Vk�
�1�bs/�77cѲ���M�����u�U��%=�����yl��e,�30�Bӽ�����#�)��L�R��tօb�cs7f�!�r��wT�p�6��8�Jq����Ԟ��Z���-n�)���M�f�E;��v��=ݩwN�F������˼qK��bpIa+�L��v��4��B���ܰmB���t8b�hS[5mѱr�%7&b�u��3Z��fbŉP�P�[�z����@C-`)1���x�a�C�l���q���
�ۺ�LYCpPSa����C���7x�N�u%���)�pX��1��0����a��^�i�5+h&^�������11�]�"j�=[C �B�M�y���v���s�,ج��i&[&��m<F�t��[���@��ǹ-*M<���[y���qh%�1[b�Y:�Z���NPݢ�ځ���A�&��+�-k�QYp�Ҏ�4fIX��1l���Q	�1��J��(|�V"�7QEW���/bZV+`�o�d�^�Q���V���/Y�����oqC��͚HҺ{�o/Y ��L���ُF��.�'�)�:BI�IQ� ���5z"N9���GJ�)����L�(T9�^$�x�c��3E��5Au6��2KB1�⧥��4feB�l�[/&غofZ7��`e�n�2���~��/�`�)�7S*B&Me݇�v+,�-���o���S�ষ���Jr+�u�clbJ�L�Z^���oB�/7i�T�y-Z�bH�q��6�������r������ǹm5�Âh�%�&b�*:��-M�ʺyD�
�DU�{$m�T��{�����/i^SC�U�:�r,Dm��(�B�7x/b&Ũpڛv�*���©'*��T5c�e�+��V�KlS2��Kte �W�Nd5��)e��dqe��Et/3+k�X�P���Z�BjU��AL�q=�YGH�v��-��(mk���ҙ�D��6���銷Q�ҍY����2�"��0��6���X#u��A�6�5�m��[p��h!5�v�N�VK�p!F��Q4ÀV�q��^պ����ދ�I�+b��fͅ9yZ2X���͙�,���MҺ�t�op��x$�?d���YC)&)o�N �ڭ��月��[�CsK+v;IJ��V�h���YZ5S�Zҳs�ī�YzU�l��h��^���Em1��*ؙ5��+����{���Bس�⤁b�7�f��ܬh�.���՘�V�DV�5�72Q�bSn��e]n'J��%��jd�~Sp+���BaF�K7�y	j��=̤�<uy�A��Vq��wPn���eX�Z��3l��
R��I��U9�q���o���Z>��7p�[5)Y�+c6�\�)ݗӰ�F���t%74�J�������(i�הu ��t�L��kFCD�b)!��Ӻ��-B�V��w�-ܳ� ����w��t����V7�3r1�c���4�X�]X������ek��� ��Vn�tE�i�Yy�iՌb��
�mT�0�hhA?��z	2��[�.��zX��yyu��V�v[1нʃU�vn�	�T$��hc�M�V�h���%ڏ����lJv2��v� ��j1�q�-k�E��H��[��F�˃ ʌ����2M�Յ� n�iۨ��0�w#aowF����Д�U/f�B�'����kwV�yV�Xp7���Ga#�#9�S\t*[�s�*��n3������+M-d�n�\A�m��s�Ee�2Ռ�l�Em�D���c�5�VP&¥%!�A��Dљ�#w6bqK(l��r�f&�	�R��:F�Q|)`�m�)IKwMaZ�eXV��x[���k+* kbZ���ꬎ�6�e�9����Ӳ�M���E5:R�E�Y�l��e��VL������
�V�����u�M�t�Ge������]XE��1�;K�+me��Bb���e�2�j�9d
�[t�`l����h�s;E,	$aVP�Q���n7v�m�,��ƙ��-�(X&���[8E[�e��2��ҽ�G�����X�.��Y��˄G6���;�woN���Q���,�#��J�#/D��I�����^鼗�Vf�K6-lm��`�S+M���Ȥl�N�b��)��Y���1c��͈��җ��,�̸M�)H^���$�K�hJֆZWt��gm@�OpR�Ul�=��ݣ�h,Z�U��(z-�z�ʗ+Qfˣ�`6[w.=U$e!`ʆ��bkF���.�!e7d�:�֋m�9��s-5*m"�F��"Λˌ�QL����jՒ��!X�I­ (Ci]^�-b&]��b�L���	'���٥6 H��pitN�nCY�[Ê荆�Z)��D�:)lՃ�q]�t�6���^�:-kv��M��x�yr�ьId%�ˡ/r`�n͗kJƾcj����Ġ�
@*^m�s(�,�2��%��@U�WX��v�3M�t,1`�0�!Sm���ʌi�BI�V�[A����lHVH邏fj-`)���i!�1(�@N1la{g)٧���57 �����je��aTi�L�(h��S����b�gn�5�{LX�����Ĭ=z�d�m}�m�{yz�{��&se�z�m��t�=?0)�����斴Gel��#��lVshZ�ƶV��M+��!	�b�Ҝl:X�\Vi��u�P�cR]���z��ṡTS��ӡ&i�s$v�JXH����ۗ�^��HN���Y��t�HV(,�o)m�a�g+m��Tj"��PP��yHl09��L�n����3RǪ�|�8F],�^֍#>��ˎ�*y`޲-n_��*ї)&*f&���7�PxEj2U��X]��-.��Qҷ.���k]$����Z.�Դ�I��7lRn�η0�ܬ��\v�1�)�"X�Wb�EwG7�Y��U����O$?L�I$5��2�]�n�Uf6إ@�l=��K���V�����˗�ZH���E"�݊8��Vu�n��j�(��	(�����/�� ���yi�Iۭ��XjH�BXj�T�Cm�@NYSu�@(���b�j�YR��4s��������V8��kq����J���Ʋ�H�TQ���ڻ�+h0P�m��Un��8��Ц'L��ͨ"'p-�J誨V��agh�P3j�t�W�r�L▙,BN����,:�+a�6�%���싡 �O-dh�ݬUh�0���Ā�î�G)bf;V2�26#c$Wd�(�����o%-֝J�3(�b��)4�z�B��k��,z$�X�n]�Q��f�5�L������Vd�f�����X-��Y�-��$��ՃX(���7?[8�G0%Y�l
P.��%�0�ɸ)`�:�	�h+Y(��}Fҷ��lYZ�\�{i*8��ԧ�<�t�w�1�J��Y�͚�hK�/����K㶷P9�aLcrU��8���4��b�����i!���nU�h�d � #wFLK�`�;!���c0�rDF�FM��	-ۛ�!�&�a�� �OA�qĳA��*��1Ndy�t쌲M�Ȳ�r�$��a qŤѼD�EC�&��6x`+�8Dn���ن��x+�f�]0�m��n�)LdD�WV�M'm���567e;WXdh�x�P�l9��:�F؋�V7K�h�u��&ԣ�p<�am1�(��w2dQ�T2��W_*�hX� ���� �h�����ы.۴n-��-N���[V1��N�;��,���{�����X>YXg׮���(�}M�&=cH�MVO��K9N��n�p2u	�X��.,��2���p�mH�Bkjԫ�Ά�'�"k���^T�z6ҫܑ\��cC���F��xԵ��ᗥޫR5�r�2Hȶ��y�DJ��;K3v���L1
.�VS��P��7AYq�b5f�ؤ֥MU��Hi��C�+KA�.���E\���e���`�q*�[�Eeл�hs*b�cE��0Ɋ�-[���i�F푂]����`��\���+Btŉͦ�S�L*f�¦|���J����
 Ė�H�FTP=��7pn��j������V��0�K�l%�����Bk�P+`^Ʊ�8��X@�Ҁ�W"�ojY���X�IE��=��N:tĕ�3Be��ϡ:��	���VV�oZ�Xp8�\��mլqb͌��.jn���q�Cz�զʑ#�ڛ)^V#V�T�M]m��ۇ[aQ�tB:�$��T�#��c����Y�4���RP<KZJʗC��mL��9@黂�h�������1ѡ�" �e�pB����@�{���`iң����m@2M���w���r�`|��M"T`�
�YZc� Q�����*(馨��P��E3^��]�%�S�&B�A,�mU��0��dZ���/5��(R�@�[�n�ۧw�)CaM���I��B��-'�ƚbP�w���O$į�%ѳ�iZ�b�<��i!��CvQw�=�[n�eIAJr+n54շ�s!x��6�嚶�6�푣C��[8��]����C�
zر���F�Ʋn�=�u�{l;�JF¤���͈([�h��i-iT6��cܬt/Dt�B���$�õ��<D5B�Tr�R�R�������9,j���`�� 3��i9аm�G2Ŷ�4T��)�Hڄ@0aYz^'�GtuY���VSܦ]�+ �d-��Ww�m�ʊ��)R�8�`��Y�P�k��ͫ�,sRDP l
7,�Y�u\����
�%�u;���ͬVd�0iA�������ee[]�h�e�k0�LpDeÐ���PHӼg�-]�G^�+�L��BݰmZ9����:�Z�fEy�J,ԗ-dO����7���J�r�V��e�Sw�n6���4bKMl7��`��Qw��Z�z��*�i�LU����x3pn6[�S7^)�^n=8ڷwVl�����+2�X!1���2����6J���-�0�1Z3-V�	��nj�C����X_uZ�Š+�cr+��Тȑ�=�ӥ��36m ��]�e0�4�挭�`��LX���B.�fQ�N[��/>iI���i��_F�
Vu��b=�#TV�;ے�*@5:�nܱ���GW��k���j�M���۶��.�
�U�!����ݚ[�&]�)�b�z��w�FLM㵎*6�t��jV��[x������/�G\<�Y6G\P��|Vd�p`�G�\TH���~���43�m�%�_%���'�N���uub�0͵����V��C:P3�
�2�reo ���n�{����8�۽F�u����K�e��I�\�o���j���N.+ �0�h.݀������ɮ���vӧ|�]���	3��4�ղc���������9+�1n�hܾ�	��0��w;A�,��.�m-���^ג�|�;���Z�J:�Y6���E�7���V�\�d�GW[�D�-�bH�8�A�wmѓ�8eJj��;��:�Rլ�M���������DP=��\�:�D����D��)�x�F��W���9��C�<��{�vm���j���������l�1�N�0���q��8��R���6�\�״~:����`�����Ug]��K�z��t�yB��N�Z�i����}ۆ� �OzJ�VJTtz���Yy;�Y�����S�Xg�9o����f�U���:TJe�\�:!M�Ѽ��ҹG��36��ʍ�=y���P�25ԫzu�s`z���nt�KS�b���Y�.���Us��#޺(5x-��u�9$�~Ae3t!�7 gݎ����� �D��{�����-�7�ݴ_�W(�8*��N��8rR�نZx��^1Ǧ�Z��Vs�!��A�0%ו͜�6�9�-ݥ���.�KB����9�z{�����E�{��b�3r {�Qc:ӽ�%��$�馮�h1���ҷ��(<�*qw���^s/�PI�ҘA��܊Gv��ǔ��F_e؊,{����t@����W���=���:![�h;ʅ���h�ޣ*���;�E]r�k5�+��u�Ǜ!nN���u�כ����f��m�
��x�)ͅK��lB��}��8�m�Җ�]��.��$8�&S�g�&�#�͙��si�,U�m��n���&�W�';X�����y�;���H��&C��nP��=F.�ׯ�ǇN��ma��3 �@fm�2ƺ.=uԹ]�-�efri��11c앯V.��r��6�����/e�µs;׎�/�빨� :�\�=�{o�+���^�^|�#�r���j���5�нJw��v�y�)v���\	(�g�i��Jo{�S�<��o{j�vi}|M�4���3W7��(l�C�q����*p>3�n�?Y��E�ǫL��۝å5����)h���c]Ү$�q��X��z�]12�Y��"ܙ.]mbF����-_f!�H�cN�v�ս���Zq�)KZ��L����x�s��k5M���t)�k�Yr�b;v�+<��H�����eG�9��l�h]�iwk�.�T�9��b���;�b���� ����	:���e�-N�rr}����4g6�:4�CO����'p%p�PP�I�*>�KIvY�sb���Ø{�u�ۻ��dU �XQ7s�y#�-y]*1J���3+�Z=��m%���o���ʴ�J<�IÐ��uΧ˓X�!hU�b��CiZfW����2�;V=�>�	��V!yW�;����R����(_h�jin�ڙt��+N�6�P�����&!G�����k���͖Q�B�+i��st�ˣ�9�،����!��j��E�vPV�}��#גL��0�ݶ����|����-έ���8j�N��b1,*�;0P��8����b�&(tNa�L�@N���.���v/c�|z��[��Eڝu}ao�m�]�٤[�yG��®�j�l�t���<�4�ӚV�c:�3��^ su��=}%{��gu�}]��3���p]Ң&Rma��F�4�P������@Ńia�Nf�����Y�p��+��:�_̍��ݑf�!�����}k�J��D�eAN��;���s����,�S!�z��
�/�,lP�Vf��rjk]'9K��dj�*ĉk�}+����Qx�l�|�K�tnj�T�;;C���h'ck�ˍ�������6+M�O.���޼���Bl�j�}$�:G�n�*f�h�6U��$��ro]�K��.�W[n̳:��a-[����PwvGnVW_).}�k�<�9�86f�>h��˃��]��W[�/sD6���9VZΩD�49>�,����ʌ&���4e����eeS��.��X}ѱ��2��a�R��J���w\�d�������3o���7�"l��e�]-�If"��A�Io,��6�ir�}`�������X�4eep���R[�o�]�ĸn�on��`ª:9��� ��aШ.������cKM�viCdn���K�g���9��O1'uOǝK�G�^�O@̬Zw�� ���],�����LtW�cz��p��T+��Kld'���
΍�ӻUନ@:ȧ�|�ӈ�m���U���n��q2qO���'������J��Mi��W99���Ú���>�ݩ,>�{]κ�Cc��N��mZp�K�ｏ�h�^eQ�mo��gr�������	�u\�W��,g.�E��zz��NAVhV�kՑ�t�}�զ�pC�*a.�2�67�띂�A ���l{�F7�2�k�jl�^}��s��y�N*��e��B�hJ�J!��k[É��EFE*�,�g��V9���qR�+��a0]mJKDq��M74i���,�N=mc��g*��٩��
+���}"No]���LQŭEnd]B�l����r�_��w��G��4n�32��u��5��3]=�7�f�M�D4#�r�N���y�P��Zs6�x7���<�hk�:��u��\6��%u��A�':A�m!��!�鶓Y�����{�]ݒ3��Z�qhVe8��:��K��i�C��d�Cr�WV����رZ�,��d���:�{S�ҙ��j���c��P]^J�L}Z��2ڼ4����E�����da>�ڲ�s\Ô��"��gn�����W}x��,��0�G��(�3����!�6�\���}�W|�3��zC��:]�<��M��N�Y�6�5e����B1�G_�%�i�=ݘ-5Gs>�R	b� ���x�nNzy�t���D�{�7�Ѭ-���/�[�6�iv�L�5t��nTsz��I�P�C-�$�.���XGÑ�a	Y�է��)��օ��$�1y]=�qd�CK\Ԟ�Nb6I�˾X�f� V)h�T;`�u-����8���`w�Wt��(k���̚��*`鲓&��WJ�Ǩ���R��P�\w(����#k^NeR����L�I8��x�V<.ʮ�\���K�3���I��r�5��+��4��ұ�in�!u�4D�a�c�y�z�}�T���A��K�g¥],������\��}�5���]�N�������GVKnB��-_>�e�`�1�e���t����vR�}5\#"l�\��3�K�WuXaP�c.e��]c��r���|��I��r堡������6�׹���Z�0r���$�Z!rK�w��9{Op�����ְ��F��G ч�4�`�M�w���/�PUtr[��Rb���lba�;C��:�����>9@i�[�Fq�{2���h;bQ�K���]*7퐙X{N]Q�+k�u��n,��X�Q�Z������ջ=�ޭ�*K�.�q��عN��کj�7���}5���1�e6����X�>���C{���{�Z�Od�+�@s��Kk�*>���6�y5o$(:w�k���PNm�K`2��qZ�I�+�}��g9�{:'`�ڮ���I��p�`�Ҷ+�r�c��Ot�u��p�<7UM��	�h��(w,��G�����m&�D���<P�ە��κ�Dt��2��h�	��q�)���V���wV��t��n*9�Fq\����+�5�Q��6}��޴��jwլ������_�&��2a�y�g}�5(u�v<���eos= ��3S��#�CD�+�������X�lBu&��z�;��%o�H�P�[������
�H��oB\/����W�t/#���p���ă��"8n�v[�&Z�Z]x��"����t�*3x��o-h���������FU+s�� *����j)L��*�q���o��h����� 6�ҝΚ��D�h��ղ뒭(V��1k�c�5����f=E����_>�lv�wf,�;Ӡ�;Ҷ[��G���꺾��O��탘r�֨'k����3*�*����P()`�5f�ja��ۧP]�NQ`0c ���̮}o]>�Rɨ24�oG��v��>|���Ul$�:|y��C��@R�(bi�]��t+6#�b�v�[[^����G���E|�s�)�x�b�Xo�7�ڸ:b�6�X��h�
����=�KNv!Y5a��ݞ��b]׷���q	��i4�}ۯ�o].dҲ��]��=�+����Լ<jS������p�kwkM�۾u+���w[�K���(B�c���:e�*�J������t�(X�0�B�M�{�EBi�	l�\�)��˳�����1��7����y�:����1�\�ntu{�"�c�D�F���0o,�R�cVp�xw]v�����oN�]������-i欷i� r�1S0���J�]�3}�Xl񇥔BU��!���T��ʓ(��d��na�����x֤�ڋ�c�^'-��bh/<�t�H.�Z�ٱ-��f;���r7�{�@����_�%�w
�K���.��!�b[�Z���+t��֛ac��Q$@u���iEmjB�E���(c�����gb܀�'wu����M9�#��_]E��'{\D�7WB��-���oZ|�jT3�Y@u�싮��c/zգV0�zlq�&یV�c.S=X�� ����-��D�}F�5J�qB��V��Ǭ);�cfw&xZ=y|�X;Ws�/�V���w�����ڮ��g05�c��[��+7��-��i[WϞ]���B�3T�@�ՙ)w\�_nAI�)�j
'�%L�i���vGw9��h�(+�S�&��&���O���A��{�X�����3�[���Uնl,r�$��	�_db�����P�g@z�m>�}w'ܑ���K�q�9�kk��2���p�0٠˖5�����W�u):�1V�]JY-n.孮�@<��?\���t�Qb��r����+��Б�%�Vd�X.*]��l�-s{�Vj���}���fv�zl!]'f�J���%�i5��y\⒴Ν�h���n���̇51[D�g(��1m)!PՈ���uLC^�le�����V[v���3�^dW\�^���q�.#�-��!�AlZ�Ĝ��Ƴ��V���+l�Hv〽a��+��̣D7fd{���so�r�=Lr!�$���0��7�xӜO7+J��@��F2�u���ks[��qݔ�� �/b��n�� ��+�q&/b�1Z�*8��f\��2=t��nە֜�8�;L��o�[{N�円�Ճ7�*�T�������{sn5�W\�b��b�Ř�=K�Lq�O�+k�9\QUxAr��W�}��S��Z�����ۮu�hGf8�����薬���K�Җ�un"���uN��S/U익��&�w�"��[��RP��ɢ�s�c�sK�r�`��oZ&t4r�Z���0�6Z�]�c�c��((z�s:N���8�7ӟm�u�U͊�^�ή��St�i����d�
i��;7f&d��K�7�9���(��ݲ��5*�;@�j����Wٽ:KҞ��j�����]�8vas4���}XV�:�\+�c����>�\�.�h��%�w-�����ާs��]���e&P��;8K��}�L���v�[���=�c� �G�l�/�e``i���B����Y.������W���u}�v�7��ܭL���s��'�u�f��ԏ=[ڲ.̶��R�*g�˯���<8��wQh,��z�u�f�~ �Mg,�#�h�*��T[����b� ��X�I*�u�(X@Ė��ҝ�5��v7����3��U�[�̦�O7�ARʽ�L�ܗ���|gN���b�܇Q[ҷ,�+��)Фi��v&}ȯzV��6/�.�J�K����e�2���Aڌձ��EuYS-gf�{`��E��Y����Nr!r����Ǥ�T��v��e5�f}����6cV���ڢ�
1�A�i��Qז(�G3��(�
?���XӅqM�����i\S�2̜�(Ju:p�ֻ7s�þ��L֍�yr.�u��u.��]u�h�}y5u��zj.�����Xᣥ�[:۲F�;���ӈ��-����</Z�OlsZ��!\�S̈��d58�!���"�WI�Y�����ڴ>{6��w�C����g�f�6r����s�+R������* ��Z,�>��o@�-�bZ|�z� ��j��u�L�6ޛyuc�b��M���K;��N�C�ܱ��_���7��we�Y���u�Vif�\�(]	�U���;c�X�u{S�l��MڎiP�m�Y��A\�*9EQ�Mh���G�kN�}fsf�P|(��
�1��2S��T��k�[�9{%X��k��W�����,U�+�K����6y��\�t��o���h1i��x:�ck����
�]vK�S�q᧣h�eҙ�"��$�W|8��~<6��!���p�g]j���ze�V���
��!#�z;yA�3M`�j;��絪��v�0�3����Y��-k�����B�P|��ԏ
RMWF��q����#���x��y�w3�r�4��ꈭ}#)}s�#�r��aeCip��r��(i44���Y5�ڮ�Vdu�A�x̱|kgE��>-]�7úq�ѐ�&�BB����o0�q	�B�����繂bٶF�^�pV*�h.�[�����w������pW%:������x�l�E��% m|;sQ�$nk�f\G�ɴ��P��4�W	Ȇ>�W]M�e�����DtU�����e����A�G�������)R,��0�+��ҙ&�^,ɰb�V��D�5N՚��;�{����s\U �6zi�;xV	��Ǯj 9� �񧫶�w�����bz�sʹ �,�.��@"��Y�@*Cu���e�437���{WR�CDՖ�ls�u�����ۓ:���������ֹ�V �*��ox#��ES뚻�ޭ�e�Da�]t:��S�(�ح�1vcW�/Q�mC��ko�N���_eu�M�T�t(f���fW+p���w��[<�M,*�Ɛ�/�L�a��<��I�c't.88�Τ~�ޭ���mR^�U5��xp=��+��Ot2��8��^�a�@��b�"DMn<ja���8k8ӝNgMI���I���tg�ͭ��K'hk��ʕ���B���p�3��W�t[W7IZxe�� ���>�l����%6��K�(>4���M��-�6�+/�n�[ ���}��s�T�t��f�-���:��k-c��f�Y�9�2it�����ŷ��gô(U��ȍ9e��u�wsW�+�O;5�!
��k��]�����S��(��]3^f1.�!|��Ql��Wy�V��d(��� �Bʆ�th_pŖ&i�V��ho.V��B��[�����`�r-����)�\�D���8Y�[��3����0��Zd�%	��-�Rgm�dE�Zg0;� �v7x-N�	T��o툅mԼ4�Ώ�	_lmYA�ٹQ��--Lu�O-��qF4�F��>�(Ӕ�)���������V�K箸�'ivi����hS��u�qݘ���w�(K�u�������p,N�����m�{]-�����h�����m���1�e�.�0�sX鉀�G���z�� ��*Crv��}��	�4���S��r�M�:������,l��&͖�K����)ې]>3@�MS�����/��0��m����$L�WRJS��Ch7u��4av����.@o5�3jb�����n�A*�Y��+)g>{�M��<m�XpZ�Dx"�n�s-s�+D0�h��=�̮4uGZ���*r���+錙@����.�^婐�G��D�ں�1��uv�%O+2�0�`�L��.C�%c� ooo�����
�#����G�R�]9=�x�XǓ�C�w%Y���&�;��/��m�1^,.��5�Ty�M�佭��9�-��B�|��q�R�Z6�ϴ\5\��f����M֎�8�qv%��-��*_
	��]CV
p5K���p�]D+��)�dq��V��p�(���`��wl�dj��v���˱�j�,:4	v݉�k�o�����otQ�/hb/o_r�����;;R������w�D�=G�<��7��]g:R����W���ɺ���9&�M�S�$	<{�(�
nê��w+��7V��2���SkW�!����p��8�մ������H0�y�*q��S�J=&�\��ĥx{e����r�ӷ����{4֨��u��c��zLܦ�^�MU��,D��f=�)Y��� A�¦��j�e<�.W|)��޸��EᎻ�L졝L��_L}eW<x룥��C>Ш9�2�.���ht����-������A���yJ��d���(�X�5/i�X�d�eӫ�.��K<)ٶ=w�D%1QUд:ͽC]'�N�Hf�a7���íf�J� ���#��BQ;�^�zp��5\�e�4�8�����9�4^d5����zY�HB̩v��mo;�t��c�bκ$޾��_=��B�X]lF�{T�Ҳ�	kT1�b�L\�h�wh�ה�
���)�{ęDVc����P[�Z���e���Bm`��CP�TN�r��@FQzkr�^vr�x*-�k�b���K�֣b��:�jA�Z��2�K��p@P�� �^ǘ�u]���kyhEO����T�{�wF��	F�w$���W�q�3\ܛ����9I���c��E�,�5ĳ~��$�ػ�E-��_-qd�<�|�5r�l-&$i`{R�j�Kz�R��;@��n
���)��WL[F�
	r	.V�J��d̥]@����:+)���T�>��&�oD��M�!m�݂ق�M�fe֪YXh��'�����h�����uY[K]fhR�'8,{nZ��B˰�p��7�wzBa�$u�p���ha�Ʋ�G��\�WX�Zv����8�Gx���K�U�	�"S���3/n�p�۹�TWKD�߲0�r��s#	�;]�.��ּV�@�I�j�9Z��@�`{{�뾽�h�I�5F�<�}z��Vr����s�f�]�.���]d�}Fv�LԆ���e�8-mG۪>(��9LV`�����^ݤ/��.[r�Q�go_i�)�v��/�mq�$i�)����ۅ�WP�C;"��pi�k�!�^�Yo/�{9�w5�ƦTKtL޼��/3`޽k�}�Y���W
���dG]����������WS��n�MT�{���7*�R70�艺�B�Yr� ������N��Q�2���0g=U��;��Z�]_f�A�Ci �̣}w:^����չ�j������/
];����X)����h�wv�)p���Sq�(f�j�pҧʲ��2m�Wtٔc��N��Ѵ���DT��#���vu��Ն��j;��*����e�]�"��n�JN�zʥ]�s� ��*��o��2�/�t5j
P���K�m��@<�T�6Ͷr���ե�h)��nU˩����'UЛOtӬ�!@M�)�uj��Z�c8��V��8R�V�Ċ+
3�i�L\q��l��2�iu�Ѿi�Z���V�рEC��>��8Z�w�oXD�����WMZ�d�ڹ�tꡌΝ��6;��t]��ز�a.��$e�3��y6�*����ڍ��X���=+��X��˙�[Fތ�9�Dq�)%u���¸m=�V�ݤ�ˌ�΁{K$7�Yv�I��L	˲hׯq_
r�mmҸ,�ˈ�݋yZ��*U����*F��״�Gbި�4o�̂�+�^>�u��]Y�f{�/!A��;N�HjٌPt�C�/j,"f_hʆ��fTL=��3�ë�1�Zu'q���u��.Wq{���ڎ;�k���Y�Zu�j:I�Ἓ�mB�n뗨1oV�k���8���]�G(��B��%��n�5iVI�gHt�ĝ�C�d���:������r�+t�r���V�c�L͓d���z+��6νͷLWZ�s�-L�c�Ҹo��[i��5݀8�5N�M���w-[|���{ g�͚,S]�^W
O�He��;�����t�Q[VrQ�F���u/{��1�/��o��Z�o���F�����<xy��h�|z�k�fh(�gA�t��M
-��ݹ�@��<q%iyV�)�;��n��Q���ǥƠ�j!���[��g�H����]k]`�foEگDgïU�w�j�9���͹�:F�Y������X"�(oNl�q��-�N�{�)oQhi�cܡ�N$v�.�Ɯ&
Uc��)�u˥,*[�9�o�H�y@�ӫ!��cצ��J�b��v�32Nn��֎Y��c�4�x�3p��+�n�oBóy�u�~��Y�oVkã�߹�J(9�GB��B]�/o�/�c�|VC��'q�@�$̤��4_�*�rh��'z�B�0��hR���;��y���dGn��i
���Y�{A��ċlLr�ޭg\`����e(�<��f�1+���Q��te'�$AhV�g|*$z���*�;M�R�����&�sd'�J^�]�[2���93���\۹4`T�����L�@�}�\v�.O���S�G�����VWכ�.���W&U���Mt�۸횅W1S^a��{
])��O�#ZhOxxm'C�V����}AZ�1�����Q��n���s�k��C�y�7�h�zt��R���s�e(���)h*��:)�؀{��W�Gc�e���3+*|~�l�x�;�)�\ �Vm�/Nvr�Ɏ������N�$�no�F+����ʓ>��E�Pfd��	�G�l��Y	Q0��;M��X��ji,Lc�/e�w^�@������w�u�R�.�i�p�6�V4{����S,L��E��iǙC	���s{��mS�ѭ3�4�rF^Ӓ<���vk�l{dF�́욇=H�����g:�ݵY���z��j��)cOY���x�$$ ���Y��t�b�IW֖M��ܵ�oB��]��N�ƘVͰ4�{�:
Ŗ"�[�;��mZ�Z�1m��p�]�Z(�1�����4&� �M�J֕t%��}���5�yjU*�v��`0޶�9�����oD�X���ޮ�xsՕ����n�����i�d5��E֢O�v�P���e�V������Y�$�L�S���sd6�2�i�f�qm
�:����m=u!�w/l��uВ�J'�����u��O]�dl�����6�Ѯ���2N�>j�H֨:��ΓJ�H��f]�@��n�=���Q�'d���l�ĥ�Yo3S��w5V�X)n�8u0���b��YǙ,������BU�RP}��;����A��gU�:���v6l�{�@�4�L:6a�yY"qӧ�*�K�e��r��+u�F��\CO�S5����8��*2�F\�ŝܧ0݋���9����9��6"�zc(�ע���{S��[�d�q6\Ή�Ab-Ŋ�;BV�/������}ԺV*cU�mTC�M�g:����KFWr;�tt�J]���)qD�u�d]�Ry/rg�!�Q�Z7��]Vp���R���fF�h���rWPc�i��IP�y���rяNc�U9EE��4٬����uMt�>
Z�К(@�2]��<s�,���h4C�4H�P�����f��bV*)�<rq�ڭ�ˣҸX*����X���8��	���v�7�T��f�8T�Kp<b8�Ӭ�ݛ!���󳦕o��OjXVo���|=N��4��ҷ/�Zsi0��p�>]�CT����T�m��3a��ͭ;k��a�[�ZÆ�@ ��%�Κ��4bf���>�@���Y/Q]}�eaWe�Ƣ(�dE�mj�hg
�t���Rv�5.��A��Ĩ@�"�9��=�āЍ%�h(�=]��O`Jx��+o�<w��i��*+B*돲c؞�������Z�䂋m�-`���]��3bg�����w6�i��SyS�uo�X�7�]_)Ԗ9>�-]#�Ԓ�����75�%}���k���:*(
01��u�/29i*O�R����Ƹ�Yͬ��3u+T)3#�2A���ws)���o���ٙ&-R��7�45����^��٠����VY�oZI��c�w��<ŕ��u	��'/��}�e�i�p�U��7�*_N)�Ύ�Bm��T�X�Ǣ�7;s�"��<+�@<�}E!�wo��vm���*�+'b�ݗW���O�&�꼊�r�䌤�A��Ʌ]LKU����M��j"OI��.V��,��R���d�YP���:��CSy�����#Gv�+Z���Gc�b�*9�Nk�:��[�`ۡ���$��R�;_n�Wk�u���&�m��Y��r���b2��'�ĺ���f�|:�˟�Z��s�CGr�$���͎�^m��W;w�x9�k�����Bmr����86+�}�ؓ?:\uA�V���L �$�}]�̦q'Bfw��X����N�s�CF&��B�)����ٸ3���}���xR�wiU {�.�j�f:ژ�]�p��:��Y�V��q�
;BV��V���SGk ���ɺ�3�����Ҡ�_�����<4.v챕�:F/��hچ6��r�6�����9`u�,\� 83,v�{��t�8�4g�Qt<������?�[�,�d����ER~jEEER*���U������/�Fr�����Z�"c]j��*�b�F#l�#(uj�-��<��Q8���VLj�	�+aV�E�;J���P�����1��q��AlA�Z��`�m,Q+[-�-��F"�h�c8���f�"�b\�ę�.5����Tg.aD*Q�Q�h�`Z�AF*[�qU3(bV�+F�P�UQ����Q����YU�l`�V�Ң���j2#[����3�m��1D֕��V�����#E(5���\b��U1�,SV�YR���q��9�o�a��uz�T�v|�V�H;\G��+)t��gB�}�<�u��*q�iY��P�5��h$�Ar�����J�g�D�v��*�Z�Ѫ����G���W�MTQ�Z���&x]O?-*��mz��_:�/jgo>���7[F�ͬ�{A�8��*-`T̗92/�7雖\���o#���yyx������w���g^Ϋ���k\65P�i���vk��	샎�]y�g\4�;����㊞��ۑ�u�B2��<�*�qs�ѫ��;�װ�mM �Wv߻����$�KdN�ٮ�T����ŭ1�W=�Z��mZ�-��*/b��L�R|�Ċ:\���e��\�M�ax����.�u�4���\�&Ǝr����U�+�N�W^�ϻ4��崯kp�CSK�|���\�5T��Y��uC.��qW��n�s������Vr�h��%���U�������Ȝ�VCmuh�K�^f�)S(�U�w+�К�e�԰_J���주9�=��X5�
%�!��ʄ#:�un����P��]Oh�|�!���{wg�^�b�q]�M�$�+8|W�k�ʃԜ�'s��A�ޫ��e:�՗6�u�i�p�"���.��.�t8N�:�ܸ��@uVr�����Js���\��f��8��6��lƔxKu�!�uI�Q;JLZ�+��&Ri!wt	N	�Cj�ݪ�l�Q���P":��U��j�=���q::q�D���W��C6��v�X�*��f`�X�t'��Z2� �{�Z��+L�Y�g�Nþ{�R����	��O+����\\2]���|ޘx�T%������M>K{�J��M�%S]���)��T�'��寅��ބ/��z�A������ԌN�w{�چ��F�+{��g��7-�C��e���QM��yܨ���ۀ�j4z���R�(kܠ�2�+��-��&��k�;WE�Q���^@��Ҥ�2���9������=/����v9���D���(�L;�����r�#Z�TӼ�R�9���69R�R��Tc����}��:�J`ȓrZTnjGow�r ��k��� �W�.�"�_,]ާ�7�j/�=�p��EbM�hs��}h\�`����[CҲ�#�틦V�Ƭ�OM�Ո�a���eA�vڨ��[V.��sǞd��N�v�;���#ړT)O����U�O��4��G6�"0@ڻ<D\�6�I�������T,�=Y�oK��Ɵ$�Rs����'�gO9/j��wMD�1i�
��e��-/J�	�f�M�����"{�oY6�y�j7;�rϱ3�WL��̕+;x���33�~jϨ;Vh.�D�:&���^:�Zǁ����8f .�R�fyT0���םCc�6?�����򑺜�Op��Ĺ�JE�":b!WA�=�ǻ��uLu�6:�XD��k��Id�~|.�������z���2+} �ˇ�!q���ٞb3�ǳ�XJ�w42&cQ*��M�mU��q\���lKG:��O{gV�^��4_4�#w>F��,�\{�Ųfz�p�d6�S�P
s6��u^�����z�o�L��^NQ���jr�.c}��5�^�kS)�+[�`��R��X*ˊ����`�}����I���E�+)�#aͬ��my �y������|��xKZ���I�e�Ng(���][h�$�ޥ��Ov�2�5]�8�}Zo��u<�<�}ْ�L�m�ֶ�6ی��*m։����я�*�����v��qk�{���I7hZf�h�l��G�%ջ�7�,��*뭼N�皖�Z�ڬ��~ЕNJbE�m�q�E\Ї*�{��cf+5Qƞh�I�W�>\s���-[�s7;�$�P��a늵���9����:�9�N7ؓ@�ingwBp�Ʉ7\!���qF���{��z�׫E�Ɇ-&�e�*%�Y�Ǣ���s�vt.��NR���:Q�Xɹ
C�U�*���A]����s��[v�}�o�*���I�ud��8����6&��}wZ {N���{b���0�"�ڝ×���u�V��E���/�p���_h�A0�t\4禠��8V:�B�3ְ:���`����ϵ�y^.���H��'T-���WL�XF^,��a��US����c��0M�T�8J1ЂbqJ�ώ?�����ҒfoTxI�[s�1@���t%Ҽ���t��v�m��Eun�n*�T�^�����,����XޡT��=�� ��Ϗ�hw�o_�/}�`+w9x���R�>�N�]G��Ԙ����ۅ�¢��1f��\�Cp#�r��/�|�k\�̸lGf�O����R�Y�f��q[Ϥ�6L{�t�s��g�-�����ϔ4�1�W+Cn��AB�� �HA&�i�F�tr��Ã��,�M�\}i��>������8�P'�V���[9ÞkƼa4�+��$�7,on�y,�2��v=�5w�����^�]�췹����F���$-�`�1\�Vs���wռV
��ok��4�����=�yki�pX��uh2px��C����pg�_A[K�m�|�jy�]�����c����)b\�w9�ީ�a>�(�ߥs��i����'��=pU�u�Z)3�4k���%g��+�4�W^�L�lɢq����&�t�j�d�[b�GZsK��ֺ���Pm,�ZR�kV�=>WON{�G���s}��^*��׃ғ��������*��ݤ·�8�f�,[Ց�Q��.�sѪ65!��瀓�$uj�b��a8��=W(Ŭ �gJ<%��:�h`����6��Z�˃��]��5~�v�֘`n�@�Y2�l�-2nJ����=Z����.m�y��:��6Ǵ���72�p�/+R�+6w!���S�\��16|�����;}�k f��x]��4$�C}�G�����Z5a츨j����Y��|W�x3�(�6����aX�XX�ciɊ]f��9�Q���6�̾՜�h��ƕh5��	���V��K������I]�B�7]����=/��}['q8�Nۂ���;��a�0�褲q9y���0x�WW�u���hCӇ�G4�QNktQ�&�vW�[\����\9���t9��\�gf���n��:�N�%��u.�	�q���k̓�zW�Y�^�3j�Pb��E����[Y���m������a2T���aB���FF��~�]O7��D�Ā�y3y������!s������bQ�\�1w^�ۉ���J��I#o��u�L�V)�¹�3s���%It�p��]\:�䐔:�޳5��/4j|b-9>��6�ӓ掅c��yj�$���G�^eN��ζb;:��4*�I碓��5�T�[r�+}!W��د14�_F��{^�������'�HSG{�k�������X�����½*��P�i���m�}FSg�v�A]G���E��yX\�n���wV.���vW,��:22R�b4ou�\U���[L3;�-�/��T�P���]Wva*)s���j�ۃ�@[��i�S��r�'��	o`[��UT7m�PU���u|��==�_q6�'=��M��P!&EٽІTm�p�W���j��Bv���ZG�[�1��Ky��5��]!�E�!�$�*�چ'���P���u!;3�G�(�Q��@�B�<��E5��'�����f�ln�=K���h]�{��ю��.�w��fYaM^L��hNB��kC3e��Sx֮�!�gy���<�J˸�.q���	�
F�V�ʞ�@d?{5]�:л��hH�J��|��mfO���S��x'^�g\��F�e}�[��n�V�&�<�RK�X���F'����n�Al�P�z{`C�VR�U
��SX�g<��vǃ��VH�C�n���Bϑ���*��c}���ugw��lFt�yk���]>��%H]��=f]2�lEO3�R�� &V<=�����>�}iRٽ���P)���P����s��N��"�Mw�;xM�w[�x_j�}ޭ\�v�zݰ�B[s�*
C;י�!�]O8�݃;j%�L�$q��5&��^�b1���i	�2È�j�9-^Y[V�v��s�o`�T�$�gj(-�k��^��u{'Ԝ�����7�V�\���lP�i�9�3{U�2`9�j>[?3���#6���/��=:K�)[��~78m`zB�Յ�Yֻ�%A.��<���P|�6�]Pҿ�����l�Zv�dwr�3}� _��������_'�p𚃻z�gA��L{8$Fz�0֥�Z�Q~��Ҏ��{vk�:yg<x�.�d�U�GG<���w���^ߟ�V���="��8(��}ܒD�t��'��o/�I{S ���y{h��)O�L�o��פF�E�u�a�sw�ֵ�С�B�nu����^z��f��S��]��7��y����Z�^2q�����Rn��΋�l"�n�����G�e`�8��蓗y|;��we[�v,M�� X�������,���Y5�;����N5�~�����{4`Oaн��cƶ�Z�3}9n�m>O����,�n��t<��q���{�;�<k�rs�=N(r�����넙Gz����n:�P��1�b�:��ꄍlЦ�՝U	���i��>����Z�[��@P_q��Ƙ���,�Ǫ����^�X��c�-3"�<��z�F�"�8�|����1�l.u���u�����8�}-k�=���3q:�Q9(��W��J��	��N��Vj+4���mD��L>�I�Zs�K�ѭu1���aF���r���OB].Vi�m�vq��׃ғ�Nci�2�
W�����W���Mlسήs7ƫ;k��s�:��Cr�x�����>��;D��G 3�2H��4�qޞ��O$k(<]}rf�x�Q��H��MM���c���ݷyyv۾���!�μ��q��X����Y((���+�ۃ�'��o0�9���Q�-�����L�N���]f,x����$��[��Jz���=ܪzR��8���Ԣ�Wa���zve�y�r�7Wnr�N�{�G�}Np��gb��ۉ�D�6m�|̧���}�;�ܛ�������l�1e=�*�Jȶj6����q�<53�d��;���=��]��8>�С`F����'��w��4���W{|4�[�;�Q���ԭ�XٝY2�����W�Y���;�j6�[��}{��D.�k+{�L̾������D��y��"���ZXK;���2�ַ{g=�g��
�oiھĪ�ku+,\�n�,G���B��A�3E���̣L^u��w7�V��ֹ\؁R�/C�n�w\5�rHlj����v�L׺��n�+g��z����I�^��w���`t��H1��e�u�����;�2�=�(��eJ����3!
5��4(+��K���$�Z���(� b�4M)�ܣu��D/I���2�f�g ��@q���w�V�īk��5��s�#�տ���Qk�6b�n�m�@�����̓�cr(�0v���CK��qT���l�e��/���������UfV�smu���x9�<�7{[�� �Ϟ�W�(I��A]�N
���w�����8ض�`�h�iڏ&�,��~��`W|�ts4ֻ��y;}�:c����]8J�gvs{�����u�p=���7�ϳd3f���B�Ϧ�]�.���
H��'��N�L������jn��o�7v���qrіsfw1Qȭ����v�9�j.x��)��"�u��'�7w�\ipgl&]�T�l�ڱ�]q�-�����b�W|�����2���Pm޻34YNp�B�c;t���\�b��y[�{t�R�R�}X:ذ�}�)n���[ۡ,ﻔ�Ǝ�lC]q9���	ɴ
�����B�c�"�;A�.�TL�����V`�kS�Q(�׭�]]�SqZS8��Uۂ%Zn�|qǉ�Sbq�� ���g��n�ε\���\4�ۥ��A/;
���|) �*ת|]��`��AC�oS<u��.vH�U�m��ʨ��Usm^=�'GF���_�]�������I���|9�]��u=��ƅ�aIr�Fu_w&�ā D�Q�v�dHd��y�.�ݭ.��CU'���v z�bN'_E�C\�.��]�����M���[�2�-UX���k#�#��"���E1����{�������wC����ODQ�Y����X��UTAV֕��Xȫ�0��������墉����I��X#��ҔQ[Kib(bkt��#Y�QE���F�Z(��)Q`�(�+�*��Z��5�e)T�k[J�Fh�fbQR�n����\b�e\���q�V�[kҨ��ZEL��+"e�X��r�J9u��VҊ��"�r�Z�Q*DTX+%�Sn�e	R)m���5ƶ���WLTPQ����)���1UR���j���c�D�Z,��(����+7(��0Z�-h��
��o��=�g��3��dRA��R}x�-����Я+8�����&rƦw_(��{����{Kd�p�l�J\�-K9�h՟�&g����r�� ��4��ڇ�C�e�Zmꁌ��Wf�Q9��.%R�I�Cj��ȴ���_}P�X�	�E	�|��)��e|�g5�ꟇR���C:��eT_��F�AV!�jr��s����N>�))�k'5�Ҝ*뮞�Dv|-k��T�Jx���wi�i\��������s��L�h��D�B�[�����`�O?m0qzeG8�������i�}Ոv��ge�������me ��S3�3N�%��˪|3lK��0ɝ��ĥA#P���J�.����}A��9�F'�BN	�U�dk��oz�e��j��|n{�UD0�T�%1��b:V멼�ۆÅ�ڡ+���x�ެ-�v��V�K�PA�G�5s��V%������W�����¾kqnkۋ�X׉<�=ب�d^���4�~��1�XyG�ӦW�y:����w���[+�>F+JG<��4��i������L�8^=\/��v�ۓ�go���A����Z��l/ ��3��v�{�7y�/�O7|�]bfڰ�aFoM�y��{v��9��q��7��ŝV��2�/�Y�nW)1]�����K�}�v�]K��g.*�*y^�Vu���^	���y<��@�5��q)���{�]z�n�nu����s��Y�(�.��J����vn=t)YB��稅�Rgo�΋�g1�Wt,\�NӮ|�_.�vvm?^�hfuL����"�gV�k*���5��u�5uk��/��G@P�U�Þu�����<��T,^!�3����{e(�Yn�����P}��r.������3ݫ���/���p����c=[җ��jgv�s���#<�
����	���9@���m�2���:�ݟ!�;M�.=�M���NW��+Z�.��@���j�%�7��{=��xF�Ƙ�0�sp%KO}�ׇ �-^et�o�G����ɓv�]�F�վ�Q�8�k�;�콚V_!!�ȯl)��+S��s�ݧX.�Lξ�q��%wV}�p�B�	2=��,�F,ol��:{��U�J�xGnoqez�ywev8�{����O+��л(�x�'�tG�ݶ�g?Q�-P����Z�-n�P;r�Tǜ��n��o9͓���=<�s���P�;���A^�J��"O_!��!r�B��{;�\b�Z�G<ڄ����m[t¥��b��V�IĊå��r�N��j��L�f�8�'�)&�b���Ou2+]�p�j���J2R���*�TN�T	즽���@�~���X�������n9�����<WS���
����O6�j��yW
�1�y��4|S�k��9W�I��Nzh��R�[���:�Et;������,������8�S�\�z�:�lmb+���L�F��C@Tc�vf*Y/�d;�'6.��ʈ�4�g���u��d����QOK����"T�}�Br~�h��`��t�=c'>ͱr�m��{��Rs����'Wt8��G�w@���\H���x�wY�Ӻ�{�G]���������{j�T���N)U�'�'�V6I���sw@*�mZ�̪��8��{J3��fv��]�k�͑��%�v{o��_]�u�<��Q���{TҺWn�1Yƈ�����5�)p+:KW7�M�G�[/_�T��U�5���i��guwf�4;\�܌\Ǐ!���(�vh��ã�OV]La�
����Mt�2Zz�rx��mג|:��:��Z�zY��[ܠ��3q��m�{�����L�N;��(k�C{#����uC��E���e��}%E�.�H���YԞ��\bӽ�}��(a��q���o� ��8���IW��2�Ǫ���<U�{�ډʡJ�J��8�w�Š�e(���1�i��'��V.ό��h���}��|VfWZ�>�ї/H3x�}�X��c�SM�rG>�_-f�ژ��v&��J��N�s�]�{��'���!ݚmQ�Z�}wV��=/&q�t}��v���Ҳ����f�Z�}�r&��V�9P*�cf�I��q-����-�W^�]��$�[��R�/��mv�W����){Z��,^YDVmqk��>7� V��e�<�*�6>����zc�81���ڰLWp��.ZsT�%mX\���ws�:�f6
1�KS�GF���33\&�m��"�����y��+ϲ*��o 8�1�t�jˡ�F�Z��З7g�����]�),᦮۫L�������ם�k�����Q(���Z����~^�?jZ|}}�^j�6rv� 
�]�����BJq���bl�&��{a���oe��Wn�1V،��r����=�N#���C}�7y��7���H��췽Q,���U��{�K_ோ<�S`�+�q�B��Ĕ��(��j��Q3ɦ�w��35X=zp���i* �[Y:ڸu��*��%�����n�[-]�%1F�g:ĥe��+rus4��
l�xE���*�� 4�����N�5�_>�D�Wf^���/�u� u2�(gViڌK+ϗTBMLܒ��r��5I�Op�S�P�Te@�[Ƃ/_Vs�3��P���뜝�7��c���x^5
��ZJ0}����uW���/�SO����K]ZX�^6��=Q�;���P����s���-A�O�]���~���HY��3mX��
�;�s۹�7˵p*v�ԾQW4*T�����f�9΢��Zs�IL733�Fԙ�U\ӅT&��N����*����8�M
�q�:8���E���bn~�ن;���pstѩ���g`���g��6�T�y�[�y49�к.s�C�2�;x��t����^��m@Mi�}�k+��	yP�GC8�G�.�D�2m�Nyi}���×����1��̬^ʶ��*=g�2�V@���Ԡ��5��M�X�Z��7�)��Wn�����.���ܐ܌ƓW��N�j�U��g�&$Z��`�t����M	�f쌗�ʽUv,�Iq�����v�� y��B���@F╪'�b��g^�K����^wz�5�q�z�Vm(�҃w ��Ƣ�''��:}�K�u�9?�^Y�������qL�qV<1�8�Q
���0ɽ��;�O�Z�����C~*	o�{��1�n��%��3X���;�R�zo��l�66��p�I����M����!���w�|���X�Zڨ��z�.f�ˇ�oyS�{'���9�����
q/o+�SyN�*�o+دW=�)�1�
�4F���6�7Sʟ��;kڗ���x�9obwݶM��h�����g�"Rc,���7����\kQ�y�Kyߣ^[UOu�zC�y�� ��1�`ި�	>���Q���3Y���0�hz<���*��E����:�Sf�7J��У;�.����Z:+	U#�Ҡ�{Ƈ^k���
�h�Q�,�a��i�c���ե��>����d��A�Ǩh�|3���X�8���]n�A�)�W܊�	D�q1ǤL� �Jo.F���b��\����<+�U��E^aWV�u\�kޣ���A6v�ml}��<��Zrb��<WS���
����k+f�����J��<M��s����������n�T�P8w�{JyYe8�f�,
���#`�r��3�:��lm��bm�Q�P���L�ڰ����f����cj�p�Д�Z�fr���j���y�����N��yt6��I�b�������,A�ך�������A3�y�էhs��g�?�R��Ջ��Q}��z6�Y��r�W�1�ֽ��?xY{��2�Z=�X���}tcC��S�|_Nc���>���*�赁9��F��]Q�lWv��Y�����	F��ے�k|��c�n�'î�Uy[�Ffڳ��	Z{q+(�>�(h3o+���{{-
�Q뾰n�tj8:0/���t�M��d,a�dR������}�yl����s.���H�D� ��K�)>�S�n�����u��od:{z�f�`ʜ8%}Ӭ�I����7/ԑ��7��r�z��}G{�!�VS���4�'�6"���F��㛵g]y�Z�bӽ��US�NV���dR����CU-*��1�Uv|����ڭ}�-!��7���֭_���vR�Y�YU}����S�� �_9=���Ւ��:�7�*13�u&(uĶ�%g��+�N��h��i�4���i��|�f�d@OEBq֜�{Z�9-���������ɱE8���[���l�uW��A鄜Nc�t=�s!�mLf��5*�P�2���<js#:�Vc`��rZ�s�T'X�f���(����G[��ʠ�^<�\�b-�1|cJ>�-�,�T�P8F���P^�q�ܓ�v��We��T6��>�=�1u&���?f�ޮ�+���
i��xC�n���֮wE@�C�q�k(�Y�v*}�[�췶o�`����W����i:4�jO�\�s� �ДN�����ܜڰ�k�]wZJ|-�%�|�
ɇ�JPέ����xf���Nr�o>�����7�'9	�������׬��T:���ʮh�1����B�S�d��jt:��%qecZy����;��q�V�tV���q����E%��\�&�=]&�-�ӑ�������ϗL�q���d�=����V������%r�[�V�7��hQ0�q�gob�C����"�VZ'��
F�\!^��������eh�?N�4�ޕ�47��'�����Ū�\2څNT-��ģ����	1}U|��*IqO�����~�x[v��\�LwlK�PE[�ս��r�jW:k��W���Py��L�ڱM���d��&��8��������ܝ�Ւ�j13��s�4W��i��~?���=��Z�]��nܙ�OF�1�Ѱ���gh�5��Wa����n^�;[%6��1�T������Z�;��crڍM�Ӕ�/�/�<�;�B"��'e�R�-���ƶ�_�+�9:��a�IJD�f����Uè�B8V���oD�:]w��bp
,�w�,��i�[�X�I����ޝ/�2>���UeE5�o%]vy�[ǌ+0%�-ir���n�p)P�Y��5>#���O���tٳ7`ѡ�
m.�g|��F�w3a����z�6�����Y��\��{f��76!�ũjod# Ԝ�����l�+2�fMn�
ﶮ�]\E��.gqg�۾r�8y<��<���j�lꫝ*��8��V�0V��7���t��4|��;�:��D
[�o/a�ȥ|ި����4�T*�����{9��Љ��L��"�&��ֆ]Y 1!R
oB����8N:m[Xĸ�∥�bȶ���bl`�����wv;��E^6\u�^�͙�S�+v��)P��sr�Iҕ��bͦa��P�운]�3<�N꿯�v���cX�}G7�Pmf��inZ����!��.K���ڠ�pjl�tQV1*pB�p��2�v�{�9AEY�\�w
�a�C�
�6����N�J�X:i��U���X�5�y��M�V3�\��[$w֭�PPx�Xn�1��v�K�+N+֥��;=p_v����%}�`������+A8���	ۄ$�f��X&��y�,#�b��Qgm�/���$��S�2�ݵs44��V5���p�(u\���r��]����+�Yjp�Wnb��ʮ���d3�7������5F^�"�УY�u���3X��p<��-��q�3b'�W RѹnĦ+K��C�	צ1t�[];���*�CQ7���Ŝ��"(��c�z�: �B3ݢ-xↈ6�p4u���3�rOunU��^����=Z�Sj��]ǘ�E�)�L�����M�+�a�B�.��c����%�>{[�LV�����P[�����ۈ�0L��;j�����没�Kx�S-t+H{�&7���9r��EcyJ�#�so�_A}f��{�N��廙�$us`��y����u��۵U���>�<�{%i��״1��5�g�8g�gow�6kq��x�]4F�t�p��W_r�ס�+z+�������9������!��42�E��+�G�9����GZ�:�쉈L�u�^�}>��>A���gj4ܾ�;�~�ZW��/m�7ˍ�u��ӧۼ�*s#7���;���� �;�$o_5{�����?�~�߿�՛r.ڠ�e�4Lq��R���*�Z�,��c-(��2��U�YZ[]�mq��մ�APj���4)mSm���2��5\�X)m)�r�[Rk`,iGn3��0ܸ�l�ZԣQ.2�h�ۉ�S\�+MfG�n᪍�cR�C.QQTĬ]f�w1��V]���X1W-���iX�h�6�m�Q+
V��Ҍm��R�"'��*T+j	m[F�i*+�ƪJ"�Ҋ�5��n�f\ws1��km73-P��6�2�J��"�J��TX��k
�#����c�Ķ�"*�ԙ��"���A��k*j�J�Գ�\rER,X"�����J�J��Df�(�MaDQV#���EĕX��e��1ULuC)`�V��M6��DQT73�b��U���ĩ�!�R�GTq����j���9�W1�~����	���@4��K�6�1wVn��ɕ�^�{��R��3��R���ʡ���a.ңqr������&&�����"rv��4��C���V*���N��]=���\�k���k�U鈤��n;����"����G��]�u���\S�p���vr���<�S�9��� �W�sQ�ݻ��e�#l&��������C��,�)W��=S�d���Av�U eZ�#!B�7}ӇqB�a�
�q}�x��P#�7�Q;]�\`ڥ3CP��7�����6���������;O�6��;�0��6����v��v=\e�q`\�̷��}O��3h��}1�끏ѫ#�rHF��Y�W<�ۆ/P�2���;K}����y�*�bۭ�'�w���)���F ��ܵ7�vڝI]�7O�^�;�̴>��y�ev8����*{��C�մ#���n��,�Y�Xo0f�z�+�A�m49���N'�"u�+,�;!���e>�Ī^ʂ�VlqYp�J�XL���%�A&d�w���w��*��hB�{JӢ ��w:���)�2r�������1�fb�:,(D�ԗ�=��Rq���P�P�U��F+�\�q֮<��3��,�_&��J�f�Ѿ`��Q}����Q�O:�6�M��;!Pt�4v�[]
�.&�Ľ���rf.����w9�����^�K�Og��0���o��TFE>������L�>���ۻ���F���K��[q��-���R(W��Q9(��(Ӹ�{��0Q��Xj�k�y��:�_NBq�'&��Pt_x?h)g��6��>w��pn\ �ӁAC�\^�΃�������[�*U�N�R˩�<���d=Tnp��Q���[\� ��P}�v��^�<������U ���7��ڥ\%��Ju���2,�ov[��8�r%]B=u롵h國NLb�����԰���[,�ƫ�Ŷ�ḵ�'�Wtr�8So{U;�V|�;�p���2�]tJhz���{�Ib��`�h^ݥmA%1��).�v�AGrj���o�,�\����h=��T��Ε�(�J�R��
�*��)G�iL�%��ހ0q�z��T�α#���e�T�C�*��맕V��׻��{NL��p���\2]�;ִ+R���C{\xM���]p����y\���[�����e�w5���=�_.}��1��C���c�Ԟѻ蝙��;����F֪|�[}�I=�4��=QK�y���H��� ����*�=���8�y򆻽��FX3�{s�5;��5y�ꡅ
�e ��M�-\bӽ��Q�E5ڷ5C��\��SL_G%�iW��1(�Ǫ���-͘�:U�eK�=�	uEU8�}X��j����'O��nD�w�vS�V�a��R\j��OxtF&mԖ�rک�E^b��ʺ�����w/�Ù�ٽy=	���������y��ʶ��D�����U1 3TЌ�tj�5�S���ŐY	��t�ua]�ʣ�A�n��2��@G�]'�D	^�W������4�iagv'\	��!b�G9L���s5�[�����wz��M:{�sRw\�����I�"U�Ϡ�a��^�{aY���8�|�Ԝ���HT�;z�4�����teh{�tU��X�5Y���k���s��խ���s9Q�f\I�>�Cr�r�@R�[5?u� ������۾�v�Jm�~�n��)�S���Q]�N�WF��Z`8�]6�&n��U" M�p�ڦ�TN�'�^=��}B�B�9��n��kn���Т��F���Sx�Nk���.VyK�_?,�fd����yk�(<�ƹC���ǡ��ww<���J9@�����g�����tʨ�˺��]D���5ٖ�t�Njv��s�Mv(����O���x���[���7�ve�ùta�~��f�y�C������T�ꔐbN�R��� �s9r�Iy_T�^�Y����t�ڙ�o��t*��]\�Ŝ\�%Һ�ي��Y0uB��6�{��ud�'=\r��J@f���x�������#��m�0n�ȗ�3{����Y��[��m7����2ul��꾯��b�m�S�2V�i�cY����8Wj�*����Rbs�KޭEr�[u�3Q�x}��^�x�^ݵ5=����|�s����^��U�}kғ��镩��P�]{>��6]�i=���f���ά��*�vv'٨_4h�'�u���U|k�2�p�n��0RJ�*ޝȴ�W{[r���=<���/o5y=D8�����<WT1���騃Sw���+et]���%����'�:�r��S�9�/�l�u���탶�D�ħc�#�\E&\xJt�C��+fv��:��̗�[�X��X������W�Q�@>�0�^�P:@n)N��lKT 8=N��g�JFA�E��e��wV�Q�Y��a�C<��ȼ'S��p�UӉ��&0BU�vp���1��].���by���vi�¬��T	�ئ5Uy�Fb���jp��}x���iC�W®�]��}(X���Ŋ��.���e�S��fu���&&v��EGn��{ވ�6���n&�O}{�	�t@���d��[�y�R2LZ�n�+.j�ea�qK���������G�����:��`��&V�g��&��G�r��9�r�����&h{iL�Z�2���f�N7�m촷�OVyo<��ב��B�ڮ���&Zw�[����J9T���p��:�kS�K���1��p<�z�zsؘT1�c��eFX�ʁ��u_iO{��by�Y�u�qK��޼\�$j��5B]�l̘}�����<b(쪎/xš̨9#y�ٗ�ef�UKGTërW��K�Z!�[�w� �+����R�3B�ч�ò��{���#�jkB@�|�c�L�R�fy���uY�ȭ��L\�����{}�^>��o��I�a�Ld�G"�xT ��):<O\xM�Y���'��Mmu��>S�ו�A�4e�<�5�+_r�8�E4U�mWd�9C��%��>z�D.M��O]k��s5����ҟ8�]�����[o{꽕�\|���\E֣i�v��B������v&�Z��r&/�h)@�f����D����4�a�虃7��MF�.�	�(�	33�ßt��bIڼ���ؼ���__WK�84�`f�B�1�Lha�p��"���ɞ�p��6_gx%K��Ic���g��W�N���|�8��	@��y�w@	�ɨ@�����>/�v��_O�1�C�]�����������4���_m =����>6�|4P����>uPY9�f*j-�q�9T��R)���m�l�hW��W5��z�
����2�P#�V�A���\9-.Y'�v�"�0o��r/T��?�!Q��
�������Z눵�BU�99�zkd�S@u4����@y���_��c���>6��lrC�u��@�˝���Nfc��sk�3�L0�cǛ�>K\��Ĳ\��nXo�yg*[�Etm���ݚ�� �~�M����Ho.`t]��m��Z�Ц��=��
�.����/��WC��P���z��.j��=.�
��\���� ��`^:eZ�W���w�ΝP] ������DF�b��M,}؆$���>��~�T�
�s�{)��Wj}x-}v[;W����|�V���z=���71�d��r9>��2؇~@�+،�nU��]S1AUL�Y�u�I���bs�Δ�w{��b*k�!9)�8ګ�kǕ�t��p¤��� g�M©�ꝺ�i�ܟ%���D§)�r����0�ɷt&��fb�˕��+�����W���hVB"������ˮ��u����I������̕��l�b�r�!�1b�z��l�0e�L]H�2����D>f��̹���g2�jP���}B�\�x�<+�lWkP.�`�����I�X|O���x8�c�ïE~\��I�8�=�3	���CC�븸,��s�sI�g$�*~��f�*³;���z �)����!�ዉ�YԎ�>�ۉa�,��� ��f���m{Ñ(��W?>��
��k��{U����v�B���tY���� �u=[.���)��X8 ��*઴�!Ww2)��E�*ꝩ�یX�ц��vl���3F_�,��5u���*q&����oı���pz�[/l��+N��$���u\�|�sh�2�?R��_o��m{�#8喸�$Φ��77T��5Yմ;���)r���G�#;�6Ӛ7C���8�2��٬�@��jY�
�xM;�Fspd[�pV�*�X�u(lPזȭU�W��5���+>�`׉M��*vyY������c�,k�+M�z�3H̩��	]�z������莼��wO-
����������1�8�٧�V!K>��ȋk���:�"��Uق�, ��*���s������~��pw������φ2���l3挡aL��uE�5p�u�5[[�V0*��b2R�eC�Qoj+��3E�s����9��D�86¨s�X걦�O&2��K��/��ó��͸D=�d�����nD��o7uI>�� ��ȟl�H��"�9��wON�.�o_��f,�4&�M;)G��J�]���C�ʀV�{�$
8�5<*�<&B�^g݃�;�<�5��s�4X"��z��1���N�@g5Zye��8-�f�3O
��{^�����R��X��Ƌ�]����Kt���VP߷ۺQ���.�pg�On�����pV��M�i�?7���V7�+h'=����*@Y��2k�%tX����щ|o֩�qf]�ʭ�[��W-_����E���n���$\�&jS��	��L�D�VF��\C���WWS�ݕ�S����)J$[&�L�u���Ф<�|}ƽ���Ϊ�`Dd���p
��rA��^+;�:�rC�z��w��/U�I��/7."|�xD���Ц�n)iu�>i��N���bJ���+���՚�ߘ뷙�?|��w�U������I���޷SD�Pk2�������i2(Fw>���9>����h�9:��K�hf���Y��x8�;PxV����PxA���AҵLp�+�5�����!(uv�Z���ݜqg�`�*^g�`�^\,1~©�5Q�S�X��|����ïhSc�5we�:�u�Ԧ=M*Ε�
S�x?��G��<<<ق���F�
�Ҿ�1*���'�9<���!4�����$+�O���P���z��t����F����d��z���p��,z��0����&�X;K�F?{'�Of�=f���q�_zP����H
,X�uz�w^�;�k������h]�����ჷ���-SQ�TQe�Z:�'�Q�F�"]�;�4���);&$�d�A����Xhe����*�0�Q_b�+s&���A%QS�Seްj	��5J�rl5��(�9��t0���(�\:��naR�Wh����6�Qc}Oqp��s��Ϡ�Uyupv{ǩY&�]��x�[�J�E�;x��@��v�D˽��s����P����DXT"z�|k(Yy�WV���Jf����n�Ym���C�S�Wf�i�b��!�:ed��_��դ�AE��Cά9��:=$�'c��oWci*�gf藋���U:�3`.��0ȹ��3�I)�B�\ښ1a�w��i�F�j�$�ɁmL�A�_ס��bu��vH��w�@�l6\�ʏV���(ʡ׈̽�
K-mKPG0r
�]>�:�kx���N���q�i����+w*�T�:J��郷y��ۛa'�������\[ve�
�z�o��P�{�p�hm����mp�p�ʳ�S��)4��y�9��lũJ*�CHW���;W<��k��V]����{��e<&����F�:������!�������Ӈiv}90p�F*��u��lݿ�n
 A՚�r�ܼ;Ѱ6ʺaoq�Pw�e9Kh؉����]¼��1pB�q�ʕ�&5#�!Kf�(���ɬ��an��rj�4��pE� �o������l�b�#�LQ��Y���hl}*u�W���okK�Vx����R'6zVȮ2�|�mmE�d;5p�`墙����� �n��n%sT����W���1���9�A�fsH����.�Wu��Ӿ%�ڔm�[\6�]Hr�=J���IPwc�ɧ*�N��.}Ce�4�^֡�Z}27�M���Y;m����4.�g{5���}�wv��I1���fQWv:�w,ion�쓜�e]�&���U��6��H`^�_=��Z�n�\�1�O\CV5M�ŧ,Qթ\�˷�{��smpy�4ڽ�8*��Y:�+�;�!V��K��{B�ipYoyM�S���4tb�W=lPki�R�vV�4n˃Q,cᏄ[���]cF�U�v����Vt��iTq�����:k @Ě�Ŗ;�l��Vﻃ�z;��Kmbڛ�]>��%/V�6���q��u��սO�9W�a"�Q�����/Yj��x�i܁A������X�1�j��u8j�T��±vrj��>¯�.�s�we��r�ǏzqW�G݁.�*�-앜�ٮ�-�9�ŋϚwE+^�����S6�0FZ5J*e��&�¹���*��X:��%b���-+6�1 ���I���ECl�Cɒ,U��+R���-u�M�U
�*TG
.e�
ZعeeT�1��
L�ac1�\q��TU�iKVDjEĢLeaR�J��P0�naPm�\I���e�,*T����J�fPY�ͷlm�
Ԭf�*��jB���
�1\�Ҙ ��XT�Q(əVbAQ$TqvШj �Aq�YU5+��ĨkA`�����E��f�ā�&�
°5�"°1amV;kAk�b�,�%chV*ְlP
���Ԙg\��_��.�V�~�xisT��o*����N%�w�l�3�=���َ�٧5�K����r@�.5b
3�/�{ޏz"��$��&Et��>�n��U��2��� �_`����S�(쪎/xƾ�w|2�R�t�L��E��>���᳌�<)��B}s4�ٯ;.o��;������Lfפ'B�����X��9J���e�cd�¼��/)�k9�T�1��i��e6ġ^�9.��*jrz�A�A�����t&x�=��T9ش��&�,�=e�dز�⅌9;/�9)�f*]��Qf
N�js�E�
�Q��9�z�G�,�{�M^��u�MY�c�>W*{`�:e�>rbD�5:��GU�]�7}BQ��h�����N*�LNf�GH5�>zO����}���N�Ywܢ�������d���1�玘�SqXr��"�V�2�rPZ�����jr�3'�AL�fQ�U"���鉽5�H�����-�yS
��b�>��j��UT�[�S3<G�o�.W���j�{���G����Dߠ���Yr������wwa�[���O*
��[�Ƭ�*� ô���V�Uo��]��5��)@Ǵy;��ʷ�٧Bg��e�]��-j�m����wc���L��s.I;� �p���G(��!R2^�Fa)���}��=�]iqngg1W���q�ى
��X
���Vvy�2�1�ݮoP���1�ww�us\D��g�"���{x�}hj� �d1�ٵs��d��}�Zy(*O��"q���C+����-pTg��KC��Z޵>���/H�{`lMK��;m�j?���|�z�!���ҩ.���35�۞�)��P����ݹ�0�E�9J��&N�|\p��SԄN#�us�v�(r@eY��֘%*��z�S�*j��)�����;/������1�Ӥ �ӆy5s1�z�#��*oq~>U=��;m���J�����j�r����aK���T��\�r�vNd�ؼ�xA���񍚘7�]�5J
]v׈��_�.`M&fz�`N�Q�RJiO�bh����N}ӳ:o+(,���Х�>���u�>f�(w]������7�i�Y�Xf\�`L�;(*s�/F�+����}�NWA��=й���~��)b�������/\���h��s��#n��2����6���y��ٕ|y��@���s�JGu��r_�����}ӧ��W���U
��ZMM��'O
�{�Z�R<�f�K�:�a�S:E%poe�[����G�=E>��坚�<�"���L3:�f*3;���$�u*�xX��NV�P�n������e���+��R�*b���RC_�N���W5��Kpt�I�^f�Mդ�7R�CI�(e�ӳ �r������g +��#s���������G��3���� �U�Mv��T5��(xQ�< U��k��ow2*��z��n���_���)�2�"8�.&+��a��g�X��5�xϸޑ�������M�Κ���"c�^g������q�����v�>d��tċ'����<���
���vjz��Ă�,���W�%������9٩��=�AH�����?�����������Rν�hx����):u��PSɟsC����3.'�q�$�
�:�1��*��5��PY�����߯z��~�~/�N�eH�v�qW��'����z�}��=IY���=�H()����S�
~{ϲJ��8�{�H/������0<jAz�3s}�>����y�g.��tu/y��:f$�PĂ��|{u��%`~k��?!���;g��0����YĞ�Xx�3r��RT����`T�l1
�Y��߳"��VY������|�61m�}�l��=
c�,���Nr��I�(b�I���t�AOY?8�>!Ă�'���0Ĝ:��%A�ï.�|���*s�Ӵ�$�
�e̝3��̰��������
r�����0m_��2�bw廇^���N�S�M�:<9��aR�Y�8$v�eJ\��*��jUS��lP8)&��rNmfDm��u�5u�޳���X՘Tw������]t杍�ِⲰ�3����K��ވ��N��~����7���;I���q��0���*B��@Ĩ��~CS���@��b���O���y�1 ��yC��� ��u��'�1@�*C�C��Th��5>��D��	s�2��v��NߏP�Rs�5���~g�fT���
��T����:����d��ȡĕ���OP���|�����Jϓ�<r�P<�bv��|�H��]����y�N��'�S1�3��^��w�=N���p�
�����쁩�Y�[J�H,�o2kRV�9���+>d������Nyg�a�=B��,$����~�����:��b�MC��P�e��4�OX;C~�����=IX
�p�Ooy�I�'f����I�"�����ɚJ��XMg�G�C�1�b.g�,Y>ed�>q*jLI�
�0���d�|�݆��~q�!�Ă��_��>@�T
�{��8����܆��J��ѹ����R��og?u;|�r��z��O��F
�_P��Y�禾��ިbC�C�p���X5��+'��~a�&3����bAa��n��+֧&~�R-`VE>0'�1c�zr}�O�r'd|���׽���soӉ8�g/��|!�?$���i:{�Rvr�'L;OΠv�=@�1���v$�o|��:`|Ԋ
�Y*w��AJ��bi�CR
�ߞ���g�u�����~eb���|y��1
�Y9�nɌ�?0����ğ!X~7̆�hP��5�v���HT>gl�O,���VVi�09�!P<J�{�k�PR:;/���}3�DL�!H���C�>� ���}���>!���PP��'>ܒ���*�|�q�YY8oY5;N�bO�vu�'̬�%NSԚ����u<�Ԃ���7�������ל=<N�*T���'��8Ͼ�b���׷�O{�_Rx�jAz����I�P���������Lk;��P����s�Mu��}>�>���/�:���U���_�b��C*�W��ʘ�S�Ŀ>�Lu:�rZ�4v�H����I0@�/+*�N�ݝ�f�yX��#���SZ9��S�1�%����M���)����}�A���҉놜����#).0gm���UW� ����?~���8����՚�������|eH���3P�������$�
�Xp���!P�%x^��'�m ��_�R)�<OΤ�������g��H)x���~��9�Ͼ����8�0;jRb
%dӭɩ<a�u��MB�釬�/�+���?!Y�Y����+�^Oy���$�
����*�݅B���Y>�{_���߽�Ͼ��s���3���;@��s'�gT�IÔ1{�'[��PX|ׇ���Ă��^Xz�ψc'��
(q�=�`~j�S��>�����F�g�C�4��G���s1�1�?���%eg/0?$ĕ��g7��'R,9���N T�8e�!S�O�<:�1�+�8}C�Ǥ���?P�Ԟ?�Xwq=@�Rx�󿸍ش�ى)��m�cЀ��/���Ɂ�Y;�ۇoS�����݁Z������q ��g�
�IP+����*G��I����+�ی�OP������!P�yᷬ߹w޳ϻ>�ޞ�3��=m �ى����x���'�_{������}��ϐ���N�n�(z�N�"�H)�O~����
��fI��_T�=�51>�D��u7mD�ks��ҟ�Y?2��>����bO���C���+8}~I�x�������P�����:V�����P���}��>I�Rtg�+������=�s�1虇�z�����J�rTX�Mu�o�>�L@QC���,��|��pi+'̬�hvʟ��1�6���|��a�i�|������̕"�����bJ�?s�y�@�S�nl����MN�U�s��;I_��͓�^�
S�LzI�i������'n%jAHm�H��cְ��AMB�{�fE��O���sp�!���|ÈT��>��}<����G�]��d}dLD�zg'�b>�1�����J�n�� t��+>��|�*��(k;I��`rwq"������OP*��Y��M��c�1�Xu=�H((|��w�{��W�K�1-1�����}S��)�Th��V��q�(��Kή�{�7n���.d��[[�2'��l��#��0��BՐyN�|9���np�H���H����&��P4/|�F�����X�7�t=>	1����ĕ
��߲k&2�zIy=�֤��g&�ċ'��:��a��$�<��;aS�
��Rb0�O;�j
E��Y��S�N���/������;}����gt�N T*N��Xk��^��Ę��Hp��Ҳc�?=��׼�5E�o�
����0��+'���;f�i�LgGvz��|��c���Ž�{uv^�������TǄǄ��.n|�ި)�f'�*w�&��T���^$1���}dǧR
?�R-IǴ�<�p���Rv��sb�RE��1}�Lc�[��{���n}'S�+��l�jv�Y��8��*A��Xj%g��
E�ʝ~���2��?S__1&�^�����B����q���ͤ�\���
�
��h��<�����sW���}@V�T�?3]H()�t���O��|�AAC����ʐS��?3�*��,1��V/�p?SX5'�+��|�E��Vs�0����1&�_�D?���ԣ�t�
}}aO���j��v��˼���Cs��3��S��Y������P�'짝�5Ԃ��T=u'���O�S�'�0����!�
,�=y�����_�������+�o�?0=k��'���������VT��I��w!�d����6N!�J������t�PXtr�'����8��<B���X~jAC�*4z�O��f��}�{��S!����c�R/�<}MN�*z�}��=�~zb�Y9�ܝr���c����u8�g=�Y�jz���C�;B�bV¡RWÔAH�'�S���|&!�.����QK>��W���w��]}@Ğ3�=d�Rެ�&�ԝ�m�Ԙ��N�o��8�S��st��H)ߴk=C����H(({��ӌ�� �0��Ăb����$�Y�+��j�8�}*��fN2�{O��k���8SY�R,���?P������V��Xx§�s���*����w��AH�S�æ|�V��E�	��z�{d���������M��>��I�%��^��0P���󊯆��A�9v��� CV[�.'�L#c���>���o.ݛ�@�b���SͶa���n��j�;X	���2��꼭ޮ�t��#��'Iqn��n�6�FK����O��I%��߼���]��ϠV��L�0֤��é���?8����q �(���k�Y��ɨ?RT����d�?&���I���WC��铈bJ�'���z��d�)�������#�owr���)�����3'HT��~l�=$?vs	�L�����e���$��:�a=@�S��x�AaXu�<O����������O�}$L)&�����+r��>?c��z�b&�CV
���X5"�s͕"��*7���{x��={�Y���`p�����'o�{@��t��|� ��?3~f��u���_��X}|�|���������=Mg�����P]�����%e@��
�0�bJ�wdd�ff��Z����3ƤY=N��Xt¦w@ǝ�z���O���I�z���<���y�y�s�}�7�����֡�1��:�� �k=C=���H(~f�2{�� �����Ƕc:6ɉ�'�sw���
[����`z�d�T�+;�o}~��E�?������H}c�|E1LW��z�d�9��q���J���Y]g̕�J�YS��f��T���q=d�
w�)5�O�N��l1"�I��昐S�
~���o=�e;˿w���������=�H,��'6�I����|��ALM��Y=e`V���>ağ!P��I�=aP����Aa�n?�R,�ʟ���5ǤC�h���K哿���瞿��3zۙ�|���zg9�����Rz޼�PR)���'OI=ggV��q����t�ɾ6�H,�z�����yC�=f$���jAd�����.c�}dLC���̬��eg��ǔNߏ�~f5"�����§~�;�3�1
ö8}��!�*޲�z`Tk*3�b�<�0��YY��:�݆X~�jS��9R�Ǿ��w�v׋��?G�N2~q�S��H)8{��8�9����J��%z>�'l�'l��v{δ�$�+'&��Y�J��:]I���|�S��bE��T��b`��+�?w�'�������R,Ջʱ��aK�ڎ��9|[��4J�0P{��+a��{u����5���rY��Su���o��̀A�)��'LjҜ�I����p8j�i��d�ir�P���`Mq�s�:�G._��{����׿��n��S��8�D:I_Y;x�?��1"���O��AN�u=��?8� ��܁v���Ώw	���AN���d핁���O��$�
�}'���&#/ky��s�;��z�y4����ڂώ���*E����>I_^�1<>��g�����Cԕ�!��a��t�����:a�cĂ�7�%I�5���CR�=C����0<W�E�zͯ7m�g������AU%eg��&'�;f$�u��Y>N~���%`~k�wa�g�H�������;�a�5'�V�r����%O2�a��X��܆�Y�1R_9��<~}��ן~��������L@���3���Ag2�I�X�<B����?>���Ă��~q��Ԃ��*(t��~��Π|���ˬ�2�vʟ}�$�O��e��|��V˃�_}�ȂG������d��}RLgn3�#�0�'�����P+�_P��'�:򘇩+���{�b
E����'I=C�Pߩ<q�=�$;�<O�ǻÿs��e��}�o�߀����P�Y���ʓ�l�S�5�$�ϦfT���
�gXT����9���/l�Oz3"�W�)=B��%�P5RV|�=����AAC�_K��]������Ο�SXjqԃ�x��>f8����_Y�;��'Lj�^�(T��������Y�[J�H,��2kRV���I��5"�%�����*u����1��.'����s��
��QT����O�w������n$P���e�'���'�ӟR ��ϒ]�+Y�l���Ƥ���{gI>d���:�$�������;ޮg�ny������}�QB���>9a��A�ΦX�~ed�<q*jLI�:���k8�P���I���|�[f��Y=e��O�8����r|��&}G��G������{��z�Nw�������AAH�O9擷�� �ϝY7�Lq�M�PćV�'�����X5�lSP������8�ϘbO��jAa���5%`z�៰ُL���ϣ�ZgyV��/�h�̐�8�mJk|}n���ReyֿkS�{޺��/Ԩ�,���}3k��+��A��B`3^蝽�xveN��Z|�9�Y����%\:xV��}H:g⮙���Z=2�,�	Xg6.U�(�7ed���Z&N�[�F����z=�6�~��׬��Vt�$�����'z�g������8��+3;�q�AAN�C��Πu;�'�&3w��7�`|�0>jER�T�����s�1+&�d��ӵ��^lp,��v��>9�:eb���s�p]I�V~jN}��c+�*u��� �'�Vo�N�P��;aۏL�x�C�x�T񒧨��m����v�p�q�� �g���=&�Aa�P�<3R
jO����|Cf(
(t�����+����{�p�d�VN�MNӤ�����'̬�%NuORjJ��g����5�j�(�O�7�i��!T|�X�jx�R�_i5O̟�gs�&!�J�a̧�n$4��5�'�������2�����	RZ'���k��58�d����n}�߻������:�|s>���흰��Ԃ��ryf��+����)�T�<C�b���L����
�Xz}M���v��t�'�m �οf�Sx����}F"�6b L{�ύ�ұn� ��_~�ٝ�ߪAH/�u��'LڇgT���䬛:ܚ�S���Rb �}Xz�b�����<u'�+>k:=�=ea���<�@�O�����\����KZ��s�ĪϹ��ށ0Vq���PR(v��^�v��Vr�O�gT�IÔ1~��njAAa�^X~~g
z�Xz��}=1}�3��eO�v&��Ϸv{7�RA_�h����i-�󣩀�5����tc��|��jӏ�ꛦ�'�G,�Y;��ۧ=�T	WP�s�D�Q��
uz�=v����]�Jo7ۙ��q�a�-�U*�k7�Uhrbڻ�ŲT�&�0�����cfD�ާ�X[�i�V
TrpI��<xy������z�cvW&��G��w�u�r�U���8���7g`����%��Тa�|�z�~u{�{U�=��X�+Cހ]W�tR�ܥΒ8�����2�m�v�N�}U��UH�y&e웟�)t#49�V)��P����*|�!7��F�r�Lsr7�;�N
t!;��>9��^�\�NOP�X/�����|���u��BU^Q�b��Q���^�	��q7����o�z���R}�ʚ�f*\��1����y³t����OWh��X�A'�%rxy��J�5=��Ч`�ha�
�K�8/T����]d}���C-�ꯑ�4��R���r\�#��>f�+�tK�n�(g*6���˙C<��@"���	�3��:����*���j�~��.5�\�BP����ʙ0���h)��2�U �Ha�LMi@	ۖ|LZ�eN��!�<�n����LT���V>�@��}�֘9�������C����q���F,�o�&(�T�s�;pf�UD,Gb'/��B����¹�C��XW�mfL��ͺM�N	����%Z'4@#�6��D�s�᱄��:��A��De5��so+��LR�?�F{t���)���4	��FU��ujE<�w�Tڠ%Apv����������
Ǭ��r=/t�2���i������s3:��j��`�e���[��u͔�ƨz3����W�F�T�������]\��N���M����ڈP6h5U�v5�]E`&�
����̹�[�e��ҭ̤��رg��v��ٲ�ZȮ��w�L��I��I@eN�][-��1ۺ!�}��
c��R�+ݚ�8Ѱy&q�ze<v�;���~��lɦvr�-������]�b��i�T�?��l��ۤ5^V;����u�����|ﺭiPcK!ӄط�(����1�&�(ɕ��S]�#�.���Qi�Q5���n�Z�h�ʑS7eL#�.YĤ�"u-MMåmn����pc���!},�H@릮����D����Ӭyܦծc"��ɎpT1�u2��F��q�S4S*��P�G��l��dԣ3em/ =l�1��ٵ(�j��R
�vӾt:b���i��&|˼��zZ�	Z��ԝ��ٹ���zn���(L4z��fb�Ǻ�OyP5��s�����8&�R�Ц᷸t��[�B�c����Q_I��Sr�״4m�s9:1+4����R��|�Q�)��#�s�so��z���+\�\��n��$m����sUdi}�htZ�s�*��׋�9gWRwR���k�v%���u��X�X�T��J{�=�Q�Pi�&�Ex.�,�݆{���y�.�T��{`RSw��y�]Y�$f�O��b��q��4��b7����Z�]Ft���}{O	-Ǔem�*0ܣt��68.�Ƞ3*ڥ��.Y��)�%dT��b��}8�h읝�N;.:�����U&,�2��R%�#���c�5;.(�1��\7���Ku�1�huu�Q�]��a��2&u,���a�
��j&dU�=��W�sR,򹨳���Eq�GJ���0��{{�R�\�L���p	�"�ո�7�L*�dvv��2�֫�!����:g)W���`p��/�3�ܧ�oR��=���S�c��=����T��
�3Ti�:�e������8�c��7QE��C=�ǓDU�9�@,-�z�m *Lʹ�2�y��1:���⤝+6���l�2��o�>���3;fS�P�_8h����ʻ�N0$�[v
|�c�R���F�ù�cS���:V:X����"ӹ\�ou8�����One����K�;M�D��\����}[%�PR�O8�uq=jY�|�1����*�)W\�޿���*ΐ;d@X,\q�1
�bc
�a�(������*fXMJ�����m��++V.$�hjT�dLb�k"�cU�B�P1YYj�ԣ��]q�*c��V&Z���G,��X��MqX�SYD��lͺ�bLdP1+�"���5��kY�"�Ɍ��QLH���Sm܋
�IPSX]��5�c�c��Z�Qq�qXbk!�1�,+3(�+d�2�Ԇ��r�jH�\��I�p�ZT�We��S2c��f	Z�&!�2T�[h6�f��AACFP�f��c& 6���Ʀ&3X�l�+&R�l��0�Qb�Ad5�������UE.P�и���Z)����*��¦����d�f�;TRVZ�%b%eE&%m\�W2�ħ9eq�3�G�����ίP�sUY[9b��mU�2�F,�1!}K��:!B��vL�pؔO�ހ1Z��W�G��;x�/O{��\�q�;�jg�\B9Je�:����D�t�:+n��+s����ܮwpj����m.�u��]"6q�T�����f� *x�¶wr�n^�<�SqST;?s�m�\��LBh@E{���j�AuL�Jp�3��}�6�ނ�=����E�/
��|�L;/�mUϜ��:Ba�l�e��S!��ؔ�C.�:���} z. ��̍��xzK�;<n)r}n�M]�����]˹1$��3�<��5�v�dQ��g�[�*���gX���a)�2�T�bJ���	�b�	4�̝t��l�Z��Ec0��ը�W�xP�&V��*���Gf��<�8y�fTJ��<vXT����܌����;�5���k�)MT0��2x;��:�f9=c~�вz�.1x�v�dc+�j�b���k+e׸Թ�#%�R-=���(�uϛ�$h�7k���p�'7��@�S���X��� ��4�Lr������P7��Xtb�h��v"���o^�t���-��z�Ǘy���p���r���9}�M�Р�"\l�q}�tBl���.��1ʿ=��=��gpa���M���iM2�U� Z����q���!ns86&<�$tҹg�6�T`�v����*�������5�����V�?�W5-�Z�>�F�;���0���S�dS�["���,>Z�t��*S>�N�C��,�����t�{<��w � �ڝ6��0N[�]gص[]���5*�D�sq�6{��w����y�]�Ǽ_J���8��N͡���/��� ��o�%�$��e����z�����n.ƾ*U��,�VnD5hTo1�*0�4T�����Gy<��X3�\J��xhʽ^��x^�y��E^�+�bu���rL��z��#z�4�]��6
��ګu�\�:u����½+�����[v��_o'��4��&&��s�1�ǔ��!�z�Ñ��k6�]�C���;5=e�=|�M��Ѳ�1��4�W��EhUF��X����\4f�<b`�y�AYh\���s�.�>�������Î��8����x��v^�F�T���<fS�A[�+I��n��ھmW|��.�z�_U�^C��r�i�V$�Î+Y�J�yd��cO|�mͭ�ɹ���ޮQ]ܾ���D�4�Lf�H>��rf.1�R��;�L̪���� Q�!���ؽF�M�͌��.Sri���9Z��spD4!�>wO
s���9z�ݣ7�B��x���dC�`ŌB��6cL�SQ�Դ��)0���%Z���Q������{��ж��`d���U6,�}b�*�R���!e*P�T���w[�P�#����~"Z�JJ���̿)g�U��~���3�R�B��bZ��S�Q:E4د�4erDh���xE��]�%`��+���7n�Y�z���*/�]�bf�>�|�$�h�b"�T3'�+��A���v��`��4j7y�w�Z��o���d����Ұ{"��XE����	j߾��٠��w|ub���/�QL�l�F�R���ʛ��
�SUՕ또탰�-͞�pJ6`��&>F�'��ɫ������y��sp��4��fk	����v9�t3��ݛS:�^��t�$ΨO&�9u1
+�&�%x�7}��dȪnѕ��C �{�c��'�Mu��wh���[�]eX�Ϯ�e-G��n��2�f��)p�ȭ֬[/�9����;mb��.d�Č������舏Wgr|��G,+����5��3Mľ��Ρj/h��[��ݵy����|�%]��F�`��>G.��4�6�Ύ��X;K�F:��|�����(=^�bz�CuQ�v_�t�~�rZNܡf���q��铀u}��^�]ߔ2�{��y;����.U"��)��V�0bڻ�l�%NG
p@���΋�Ƭga�Mޯk��lR��ƉgG�^N׃�gxG�V;�ɥJ��s-��1���f�=ʸxr;s�G�^��0@�U�|�9r�'�T\��Aϻ8''�������N:넥y�}�Վ��EI��eMF�.�@�cʲ1wy��OE�^s�>hi."W'�ף��N��kB�;ź͎���yX����r�vF�)�a���bu�� &*s�)���\"V�Ȭx_EX^�/���1�"�R�⪼� )�bX(����'l�澏���b�8w�]�o���J�hݺ��8�/m��x[5��!�R��#F�j�T+�=u��j�����}��#.��iO��¬'1<�
pӺ
��q�����dݥGWr� Z�՛��r4�<�\�f>'�V:�w�_E���w���z�셪S�5���l��xK��p��ʌ�|mT*a�D���ԛ2�3�0o���ͻ��g�I��s��+�Ky���C���ݜȭ�Nz�gxV�sG<e#1x��-��F٪��gӗ݄�w��¹���Rb�w�ͦ����
\^�2.�1��	�(&~����NZ_)�8���R�Э�B�*��Z�NΏY��KpJ��Dl�U��KE�� ��!cQ̩aq��gPn����]/nNX|=z*�|]{9]"6q�1R�3(-��"�g��ͮ.��p���1r�8�
�)�6��9{LC� "�H�i��?qm�e�o;�����W�6��ӵeL)�7�zT캌.q�W>�1lyVV�ݞ���Rq"�!N��Lƀg�\@����@7��~�f�gg���.t��Nzn�Bƹ¹0	�=FaʞŢ8:���\��XO��\<�<������`�}�5((�TJ��Y�����>�`��|b'�ч6���Z��@}�����'z��
|��G��;�p!:U���/����k��Y���lq�6� �&��2(*#�8�+��/�G�ށwV��2{r`Oרt}Ą� 3ˇ�+�iKv�]Ecο)���o�q,ܶ/0�����<�\'f�#y�,��N�jT�&L;/��Lp�a�])��z��zzcK'dl'�ٷ��W��1��P���GF�3ȉ����U��U�}_U}��G��:< �
������<��� 9��&YD�F�g�Af���-Y*��i���|S�tB��v��h�xxQ��^^��_r�@z͙�<\k�o���C��"R�%T����q�"��X��ܹ��L��HHh���X�y���;.�H��������ܵ��KpTg�iàY���Sެ~��s�چ�����D9��!P�T<5����Ю�݌�r �&9g²nq�w�00��Mj.i�3t��;<�ߐ�{�����YP�#��.��i��oX�;j�T��lʻ.�ɲvkj�wO~Y/�5�}u��55T}ˁ���k8�t8�j��K����[F��G*:.��Ԛ���	��WZ�l�Xr�:8����u��u�Wk,��+�p�_[���"���{�+���ݹ�q R��E鲖�՚���c0����:�j'9�pY������w&�T��5�a�ً�"�d�߅DY0�s�Y��V"�;)ڈ\��$�9�1�㏹2	��8�3�)S(������xk�zU[��=�����u5xW�JQ�i�ի������=s��0���h�����
��.�'�a᾵u�隙���l�7Jl��^�K�3Ex�-�\�c7"i��B�c��\���b�p�<�.1�L�C�Ég�����W*�#1~,ƁHC���MZ132y���3j��xy�󺕛ːԖ�TP�90��M�NV�.���spD4"�3�S��Nje%m�`�u)|Cڰ���5���4!U9xW�ƸL!�<����Ľ����\�4�	��ұ���y���eE��E��j`ʓĆ��y�\�WR���N�d��+�f�FHy��)-|	�'�̿)�L g�N�֋�7��خ��gg�4�D�x���Dhu\�$^��h�D]���G��.b�[�k%] �ҍ�m������w�8̹���%��:ʌ��KC�=թa��*=�8�Bw��Y�	Vó.��|����.-���w�Wq��Vֆ�Z���6�)KN�ȵ�z��r2�O�SV ����W���(�I}�x�_n�E�:f~����@��+w�'�wC�x�L> 諮X�0�:m�H�o��]�o���T�8�^i��d����ŵ�4E˛�q��*_oj�Vw,q�LT�ߨ�C��L�{�`�+�]�2�&���[nQ�'����=�f��
�`\��y1������pȕf�ƅ*����b�����%q����n�UyŨ"sqK�J��`aY�}�g5V(iaӑ/�{|����́�E3�����wڝӗ5KÄ�Q�9u�0t�����:��J�sӱ��Gj5�U=Z����v3x�q��$��y��A�HXj��ٙ#��bF�nk���0ְ�®5��6Y��^���Z���s�Tcg*s��8 BQ������IMd�33"b�Ã�8T��C�x��_{��|��Y�x:��DV�a�m5 �����%��n}-�TO�����U���5��x\��v!�,��r� n����R53�n>�J{S�s���UͣÕ1��q�w)<2]�snu��[6j�e�����W�����h�����ĵY�����3xWf�_7�S�fwi�a�����Tt]�J9ߕ�UjY��C3p���5����=7M�3�g���&�Uu���1����@[ ����w�
@�:k78}�Ԓ��>J��~��u�g�?Y�xxW��<s-m��Sy�Q婡�^7��v�)�����`?���<44����g����pО�Yb�<���;��A���8�@S^�(O�N ��d�j����r�K���o���.�gb���i���\�
g#j���l���q�E*��B�]P�Bbݡ��~U�ݖ�ݾ��0��6�BgC�H\��c�[���������h3j:�u�Ľ��[�CpK������yl��j�yeN_v)ʽ`*�º�<��]{��nK3��� �Ꜫê�ר��c#�PL���?�SG�o��	]�z��]&�.ꢯx<�ьxGf��L��腵3�-�6<݈��*S84yN��w�pM>���I�82i��F0��ϕ���U��TQ2��Tî\����94"P`��w���xȄ�A��}�D�ẗ́������A���;]W^�g�7���g�ğr�v5����h����<@P�Pyا\O��u���D����7���`:JwX�i7�Eٛ�N�RB��"\f�����z"��]��̛�Ҿ�/B�S�m�r� ���@�+���N�Tf�P�G��)�� ��ʙ�u�Y�\�ѐ�W�,�uk��j�|�V]S}��[ȂF��8�#D�+�w����q�A��P�+e��4���\�a�n�J�=R������*|<<:��åۮ֧���
�Z�$X�����4�t�+9#�t��5���@L	�&gYS�90���VPY�9;QT�����&d���rʞ�?T:��aP�!�!�bN�aKdp�؆S ��j�7������@��N[*��΀f/C���wN����DO`��-��-�ܤ�Z��˼ߥ3/j¨p�T��LW������8q·�U��<Mw�ܧ�h���Ovw�����'�,5���>���Wָ ���J��.@V� ���}��7�ή<ӾG��6ewR#_�#�>�T�䕷[b3~�0=�L˿D~�5(_(W%�^(�~��������8�m��;�[����3+{�2"��q;���s7�m�v�%pb��4[@��[q+�Gi��d�6��ߠΠ�XHg������[�q��h}Q���Fe���0�ל�g�1v�W]{�Ry�{w�7C3��ۖ����tz��ٜPG/��$�Yj����3��/��oxY�ݚZJa�0Å�>�W�^Dyn��Iw
9\��
v�:�(,,U����;y&���m�k�?2��=\�Xd�39��A�X�3���e�{-vSc���{B���SK0���`
	wjF�b=80�;MԹ(��	�� ��XMi�]�B���j��.�C�g`�8F��5���h�>g��g}�
�~l�7��V+bu����ꛂ���Y��KҀ����X�i�SS���ܹ�n�TU/����U��p�8f�9�0Y
�7u��'pl��t��%]�����G��EW���)�����	:��}S@����Dd\:Ii�r����vaU�]�W������\n��5,#�+�u��֚�����:��yZ����^2�9�+-����r������iRÙ�m�ʏ�������(Ck�X�x;�Ec��0��`�wo����R��0�Z.����t�o��M6�}��{7�Yz�%�.�$��ț�[xAK��:�x�>�U
�r]��Ǵ�ky��v�d�4戓�Wq7���f���t=2�Y=�)+�����d#��n�RcU�3X8�j�b��; �9��lL}Q��;&�c�7~T�Ș�I�t+���ԗUѪ۴������6e����5�9̗\�]}K2m[i9w۴7)�7�t.�T��z�Tݾ�0b���:�r����/�]&x���.��i[�SὋ���T�P�T�Ӂa��ia��%r���L�wxkk)���'�g���-�9��q��ő��g��΀�
Nb�p��ҭ�t�ay+�:oa�ْ���Y�s�vu��u ����v���Pgf覆Ej�u��Cgoc�PQ�%l����,�%U�;�l�Q�M~�.������K����%+ݸ��J�ԻN�%��&MTո{P�[� �u�
k�����ۊv0���dj\�3�gx�Q)_�9]͚}\�:>ה���:uc�+.sSs�zX
W���y��rc��<�:��kv���;��篕��\o9�R��ʼ�ٜ7���r��+��ȗl�[�o"9��{���k�T��e��֙�-*����o�y�����Zɻk*��E�Z�$��e�(�YX(V1*�q��P�E��!Z �e�Qe�Ԙ"����l�X�-B��
�`�q.6E�*�%��	X�ka��U��Y��\��aX�3n*kĪ۸b��X�JѕL��`�+��Fb��Z��\¨�)hc���I�J��UAB��IU�UeJ+R�`TY+&!F,Ė�ʥjk*Mu̲�Q�Q�l�`b��bҍT�jC`V,Q�+*T��U1��e��VTSm&kkZXP���32�bl�e�V��k�f�s e��[q��ZɌ�Vb��J"�ڤXcq��XF��,�m7
�!�U�V��i�m��� *��J�S��P�b�6�)�]�T]b�f2�Q�Z[��3a�VE�`�V(��e�A���DUʊ�9iY�mIm�Y��X�L�wi�`hhꏫ�}���8Fv�Eco�g�q�+Cz@vc�(g>�9l�z�vV��Ț�`��+�ՅBԿQ���z��6stM�������CYBsq��H���3����y�F$�qוzԧS�b���t��p�����%�[B�x�es�Ku!خ���'{��Q�5�]bBY�5��D<�=댿#��A�-�1SR&Z�|T�Kg��R�ǩ%�ງB�%��vcv0�X.*aK�yqb�aI���~�f�P�̤�d.��32b��!�0禽�\�b.s�ҝ�ʞ#x���;pL�S��f��ơ,G1
GK��<�xoKu�\�:V��=�ec6ᓄe�ܲf�f�����ؿ���uB�Ӱy}��iOL���������#/�j/[5��Yډ=�4�lg��^��!׼ߑ�h���Y��V"�ۇ�{&��㏒���ی=-�W���`1�z�<hD��0� &c2�I�o0൭)M�\Ш3΍�LT칽���9iB�Ȇ�Pgj�1V��ʮ�Q�OׄU=�x)N58:y�>�������@WI��]��!�i۽pv�����5�0���㏸429��۬�K�l�SƷ���2[��.�~�\�Z�P�]5w�W82��ԋ�k�B0�Z�����;E}ܾ�z=�o�BwbOA�������F��"�S�)�B��j]�"Pw�N<{�"�va�cn[��&\^�.(�#����ˮfɦ>߭��t)�Ha�T��ܨ�ow��#�=3� �]��j|4D���d��ٗ�c�79�9�wE�K�^'eF��s�2<�J���OMB$OM�{nl�7�q o��n_6���.Ҝ��N��N�zs~�p��Jwt8|*�$lĬ"M[����;�&F^�4��9fz,:��Y��_^ Mk���c_ǰx�´��khh���GfWH�d���E��#}���:�j��>i_�]�bB<>ك�ҥf*�Tʜ���7�ٍ=�v4T6���F�91���U)�
l
qSܺ�=�׿y�X��@�L|�`E^�eK���I;�&tWH�pdE�H�sT7�DY>SO�B0D�����R�vA�`��=.v:��6��#n���t�'q}tu0`�<���7E+��9�z���`.�{��d�6k��m'+�)�F�~w��ƃ�14�E��=�U�K��Om��)5���ױ�1u��������l]�4���k��䆕���zc�Xo&hmlf+�*)-_{��z.�r�M)ښ�"�߫����苍%$��#�U�h3)	hƁ�2�V@��έ��s�W�a���X!�w��x�B��Ƈ0bڻ�l�%O
NPji"JRf�aO`{|mJ��T݀2P��`�,��5xxTV5����X��</8���`�kք�2�ˎ�ظ'��eUe�����αW��5����r���Y3j�Y��+@�,t��"g:��\1�e+�S��6���(�aU]yp���<7��U�+���r�1�O�_��ߘ�>�$��'.�㾮��G��`f���ͮw�|��0? �~���+P�`_)�0mRX네��<=k؅͑�L����k�F ��z������$5�P0��@!�Ha���6!R�/)��"��Xr��?;W��v�p
���E�i���|p��jn�˓��Am��M�vH�ˀ��BgD���S��X�)Uo ���P�x��Z<��;[~���*֫���������3ڱ�n�q�T��іjj�y��޵���h/KȻ�q���mwWm�VF��Au,¸L�G\����:ޔ��v��"{J�|L���Xs�8�:�v� ���q�~����,�䛢	͠g�ݡ<�Ӿ�>�㮐�F٧�_����
������l�ߧF5���;����9���<�ٌ��0L9A3�7��M+>����)v�c1��M����������㷎	]�tF��`l3�������~>�7�N�JK��V��TKGJ>������7)u
��ʊ#%�eG.`vBd}��o�E�}~�{����B\R>uf6U"�)�=;h�Ӟc؂b�}r�&a����B�xrv���ڀ�䀃»�ю��|�L�p��9���o:a¬[Z-;|�i2*�������8a&�f6 =���.26���,C�����k5�w9��4\*��OFC�>�T����Z#�^[�֧�߀�^߅B�o�ct�N����Lf�H��1pY�5���PL	�&f�ҟ��
�t��g��+�w�Y�=��B��YdzʇP�#�u�3e�$�T8x�Ձ���O������Wj크W��ɾ��yS�P��:A%��5p�t$�+�%�PGG1RQ�Ώ΅�+)�
���熅���5��5;+�jZ�ׇ�:�&-����g&��+e3�idĺu.�pnG��)l�S}	r�=����Y܋�ٰ.c��>�;/��؎51����D�vLtj31�	�
;o��1];պ٫?��ނv�J\�Y�t �
yXI���J/�^�2�<��꨻��W.�j' $VH<�#�O%���'ə�8xQ���n�߸)�e؎��7��qK�Â:�^tz~�.J�����j�=ڎ�FP��l칀�ۗ^tR�׊����e��^U�Á����["��Y-h5-�H{��w�_�?oxiq��3�߰��dF�S�Zꊇ����m
�<����"�Pu�T�ߑ��[�/����M�8d��.������J��/fʹ\��~u�K8�'�D¼�ڹ7]U�L1�Y6Iv�Xr��
vpV;\:�����
��R�S�]�b����z�5˂F���láPɄ�ܶ`�� &sL&�Ƽ0o׫¯����fڼ͠f��W���U,`u�tB�4e�!L����k�!�,0�t[ڇ�P�j�K�����<����4u�{�U�8Q�|�W�˸aw�!�ZP�]�8gJY�)���eYB������<�frk����)�j̡�n�y"�6���uN�w�>��6�[��;Uޟ�/��휮������N,qΪ6}?/
��.=�G�@�F�h��A�)�|&e��)�{r��%�d�w��SJO��w��5�b�����nD�uL��Lt�'�����D�瑁�{����Q��rvrz�4��[��#9��,ƀ�lc�5h���0Ь�}�^�l�g�w��z��JGHZ,`������\-Ɨ.��.D�B43�S�g#��q��i緼�D��j���[t�F��І�9��މ!N�e�%=k�j�gvײ�/=�*0^�!��Z6�+�u��XMA諆U�]*���o���(��

�R�����a�1�˚��&`�����|����w��/�}g�n�]8D��ň"��ꕹ��)��K!4)�5���D�黂�ܚ�xo���zz�;��XW�B�����u�}�����>O�91Tj爇�ͬ�w�k�+7Z0K��XWGB	�>�X��: �Z�q�W�Y�XV�:z���ej�N�r�o]fA�A!1����n�l}��u)alV���.6��R�h^�[�E�l�NG(���e��Ʈ��Z}��e�
��v�Ιj�xҌ���v�1�Xo 0�{�i���R�K�z/SֹK9@��뚔�џ��sqD��F�5x}�t�X�J�g�`֮y^�N��R�u�������2�ʍ�.�%Y���*�y�v�o��Z�@��<8vj���s#a�0�ZWۦy������o�������ݣWK��f{ ��x������K���W(��y����8��3ɁF8A�{�ۥ���*����.�J�}~�x�`R�E���NP�yF�2��T)�wuMs����3[4&e��똯Fq�y����=�Do3zŵUa���#���L��ZIĊðe٥V�{`��5�Q��}g�Y������	�@��檻a�3��֒�sP�z���u�]��U�ݳ]uR߰�xQdg_��S�]+�,��O�/���^��o@���}�@u������<#��>��6���s8Fv�3���z�=��><����N؁<�b5'S*,9�I/��8_��G����{^�+l�T9���Ʃvk��w��vؗŤm�ܮC�,�}����+�Kr)�I��Y��J�Z���5�(X����t^����qXz�}-�����������g��6���(��G�^ݴ.E�d�ET�K�{nwGBp���?E�0���(��|�ĉ��FgDE�DPS�D�B� ���Z�%[63tu���3���v�ʣ�˴e�Ɉ�́�#����ǀݷ�!Wt�N	�R4EJ��V�~�\��L綩�ζ.��]ͅ���b~�N��C	�j�0P���6/���C�٤'���R���}���b򫣮�A���Oo����J���*��g5]>��l�"p�S	�Gʴ���ˤҀ��v6�6S5qfd�B5��4ٌ�����[�'V1[;�$���"���a�V���m�S]1St(4�!hrFC0c���g�����er��mzLϖ=�=ڥ�:&����Y;.zD��Zo�ygAKG���������;�x���z�ׯ/�����^Ly�/��uhl-�)���=ǳ�bf%jㄜ��:�bH�F�6���a*��3y�,g�v��/
�u��Mp�<r=%��#��C��\��㴋�	e4w;���n��[6;�}�L]i+W%+�U��s-S����f�����9.�Ѩ"G;�3���Ugi�|��ګP�f����ҷ�"�81ªj��<=#8��(�]�G�$�ϒՙ�]���!�Ӥ �Ӈ�Yj�b��7��kp��|=Η��Zl�S{�ʃQR���f�9rm��7ӳ1s�ß��^d#����	�fc���3���B�v�Π�4,��j3=^	�&�@M{�9�{�9��.z�nq���Nu�]NS��q�����G�E��ό$�f�%Kd�+���9��q<�V<��+j��6a�R0g���y ���SCΑ<��*��L�b-Cy�f����nEIo������+�����/�VS��N���A��^���iZ70�u���mX^��Fh'b�~ɵIa��uӎ�`��EU�3'�N��E���;4�"�j]l��."�j��D{5s���~���}��^:�B,����&�vJ;���R�A�8�DX�^�P�Ows"�{��yqP��G�Μڹ�M�N����Z�[�&�C�3�_���S3�S	��I�B~�XN�HV��V�*��ȧs�L���\�`j�)ʊ��[3r�0ֹrG/YpW/�Œ�^I�X���nlT�.[�+�E��"��܅fhF<����4��O�fs�nKͧ�U���,gwd�0�;�蹯b�M��*���4r�tvO �d��~z<1wϗ�_$vX#�/��c֮����YC����#z�-|=��C`��=i�D�C�6�P��Ka�c8��h������R� �p��Ywyc�j&�ͤB�uW�����µ%���&
���sL&����Ã�^n�Y�x��;����o&l��q��h��8��[fX�^5�q=���C^��v�`�e����{��Θ+��F��������&���s�,"�2��g�ap��ӈ�a��b��5(Tzn���8�ۄC�-Ʊ���nD�K!t@	
%ML쓂�]���ۡ�V���8��S	��ˀ�N�-E�_��3��)-^��ӕ f˨:h~���ae<��sd5���*�d�Hl�j�xh�
�5��GP�����'��׷׹��J+������hu�+��"ى��9��Sf#L�S^�zËO�Cd񂻳�K��d'���]S-28	���5��T}�5\�0+�3��ۯ�Ɛ���4��?=�28�
]���W1��t��me.�D�7L����1յ�::���CA3���Pm(��gǩ���ɶ��]n��[��]�(�`�m���E'z;�
�{�i�򬻚���;7Lz�u^ԩo=���d�{b��:�1����RLdmQӶ3���z���J�����3X�Sa7��Ӕ����5�������X)Py���q|�%�z[��q�n�������K�#[Ե�z��b]�D��`��w!՜B�D�̨%L��(s�2�{�r��#u۶^��879���o��I��R*�ϰh7�sƖ伛�>֫zd��Mם�+X��.�=�J� k�r����+����LUn�p=�k�!���S钹��(�`.�uv��K �Y���1�#�.승
OUv���@&���¸�UM�(�oFr��o;�\$|ig%�_�Jf3�x�+ˢ��ߖv�
{$�W�G��2��,+�)y�;+�w�mJ��{v���;��[�L�+�����B'���nU]A�ڷ(kyX�ڸ�YG{��cX�U�K��"�͢�b���7Y*G�;�k�e�(M˦�q�t��,��#�{��5��}7�(�3��.
ު�evF+R[7�)��r s����v�~�oK����M��V=㱐7{���1۫]x1��wIܡL�|�#ќ��u�dѳi��-.Ae��r� ���;& %z�#r��VH��خ������zIhDM.z(��<�d@#����n���YsH�ct��f��X�Cb,6�c�AyF�tX^���r�Wb����}B���:�:�r�0s��.�T�}ו˯�}� BP�֩�i:���M���'^�4�{[ef\��A'#�\Otz��RZʺ޻u�e��:�X\j�+5��z.�GՎm����(
I��JU�Q�Z]b�(��8�}9����@|z�(������s��S�9�:�JWK�tf�Kz��<FP<�DbÆ9��SHb���\��)hH�}�**b�S���)�| Z�Z��R�%������z�r�em�bC�,�v�w�:h+yF�۔8c�;{�L	��q%`r���+������!���\��3vG�����|�v˳]��1�ֱA��rQ]���)��Hp�8��|�v-1��i8��8vF^��u ���ΕC����^����Щ3R�Ҷ�Ha�T�����".7E��d��}^@�k8���`@��aw����B�Al���ԴOR[�^.�zv5k{����p޾���RӃo�^PPp�U���؆��VX6�U��.l�e�miM-(���q�əTZ��6�j
T%J�KJ��c&�X�cw01�J
T�,YZ(��%V��Xl�4�B�X(\h�C+3
��Mq�k�,Sj,1U��1�@ċ٪ʆ�&1b�TR�XVc�eef8�`�b�VT"�P�ʚ �kL����m�&#J�ESTk\��-��,m!r���	S�r�4�E�[aG2���E*UK�a�qp���Z�`�1����
ȡ�&1E����Q1�0�+++
�w,���!u)�E2��[eJ�a�0r��J��f`�¦0�Z�`�RT-��pKJATr���J�j,̥d1�.f,
*�+������ւiT��n,ĕ]h�AHѪ���6�3H�0�TDEm+�7�7���޾����f�{�//mu��L��:(����._:淵����w��K�7��k?%B�a�N�1Ev��������W���Q!��f�'��@U�`Dd�r|4JKd�me��l�g0U�]u�nv9#�0 t��wjj��C��(p��H��#D��<(ʯn�.�:s�<o]�D��ߩ
�Q�L�ڧ/��3��)3�cE�3�0ðswi�x���ɸfc��F�XY\�bp}�}���u��G'�-A� :�����n�[�C6ɇ�ݡ��2�g�{6iҿ|�;Q�}��
�xf{\gv.�.W)�ei��vy����T񣼼L}����.��	��-���?{�/�>{��������,)sKz�m�H�;3�����q#�ύQ���֦7\WO=e}��5�9�����T��B�Ҧ���#[3*��<GT�_�.e���CoϷҵ�����c2�F�1WE��C}~��x�/D\h��Ny��4��v��j��O8�VD�c,��d�̑��1^�\��
x��
��F.4F�7���w	WN��9Q�!��t�,^�:�sz��^غs�NC6�������z��vn�P�d�1���+|���.K�y�*��-h3E��JQ<�4r����g�;3&�дQ��/��Be�Y!�A|�:mv�fs����yN�wsΦ�/�{�ټ�7 �w	���&:j0��I��׀T#�P�s��xFhSQXq�L�<���G���U�z+˜^_�M*�3�,�,l�W��!g�)�L^�*]G�s��.�{��XW["A�r�2�`s�L��%N�B\߫7M��9�l�|�E�*��8eM�Xqp�MC�=�.��c���>ht���)+���!VeR���&�Vtb��GP�S�\F��>�&	{����uN���b(��2��e�����Tgs��=�^Յ.	ʼl�+؎�ty��yW���BX�O�N�Ū2&��z��z�����'x�tT�RX<�Pp�;W�.I��2}�N}]eL���܎|��o_6�uT�d��ѧ�bkN�$Oe�:�!�%�a�@_�?
U��'x�\��R�fs2�gw�55:��iꡢ��9��Mr�Hh�]�4�r��<�<�6Q��O5pU<+&2�̿1HC���Pٌ�����[�'VC��2M��]rL���a��+���+#l�<��+0�u.UeD�ͭ��.ƽ��*�j^K���csۦ*���ya:�����̅�'1��K�����ONt�m��f��+@��+��f��,��}J	��&��)-u��n�
�Gu���K�z��Ăqfj��2w����#��NaW��>��<��.�p�����/��6'7<�<�<��*S<88��k�[ا��z�Wu�g���#g�k�[�*�j��P��.,�k������톴{*��C\6��^�s똘7u�+{7s]*X�Q�Ȥ"�eVY+9�E���k�$��5�ʞ�.a�G#����s4-�9y�sy3s���t�sw��B���8zU��f�(n;O���Jk��7'��}�mD��q\aKcg�R��Yf[.��N˕Q8D�Y�BWA6�/+o"ë�r�m�C�f���t���`1�z3=PLR(	��t��6a�w3I�;Y�㉏z�Y��Q�m��%�L_`��f�  ��Y������,	�����(~��HY�Ͼ���>�haټgg^x9Q�j`Ɔ�"x;�\��{}p�'/�Vhs���|������	���g�*��+	:�|?:����^Z�8�]wԾ�9��G�gu^;�r�(����Lh�&�]���u)�P�(�&��@�pSZ��`���0��1��3[����/��ި2�Lu�lXf��y+����ՖR׷]�o5�q�b�œ�o��U���������w�+直�]���^� �H��5a$:���}�>Kp'���w�(x`�����f��6��Şy׼��ۼ��X��fc�.��}���;4_"=V�ɮ_�g3VƷ�r�X�v�Y�z���$B.fN�BtD���)*�P��L�
��u���z�3_�Z�^��*��K��
fGr��1���U�1��*��Ӵ�I�`�����M��X���+GmbB:��H���!�^��abz���i_l��9�>��<<�I-���9��Z)��Sig_ k�:���ʱ��7WwV-�sۥ*�R.���`��o�}�K�?$���iq*��u���9�:5�V�Žn���h�ǐ�NȝaN�8��\6e��1
e ���WS5b�z��p����K&��Uoj��s�\��o-�MB�PPǜ�140V�hN��X�s�+�,t���=�+6�]�+�-�k;8�H�n���fw�����'t��W��j�Fmg_}qBUb����@ŕz��/�E_=9�̻͌{4ML�'T}���,�C)faJz��xT�5-5��)d�J�U���6聁s&�c��a���P�ԇ�/�����M��]Mt�zc&�cc�F]���3gΑ��Kʰ�\x{�z�cs����>���H�p�Q W�[�;>j
uC�D�Ep��Xw�:�͑�V��t;�ĺ�zo��}.h!���j�x�u����t�'�\�؅6}�h)�u��֐x�G=��y��a:'G_��:����6�:#�Uyd�]�a4��+Ϻ�ՓSx��$�����-�V�s�'���)vFIU����8[Yy�nc*�U��˥� rˌ0 ��{M�o�4��9*�+���H��"6nSG����S��<��d>�ᵢ�~��0,��.n0C��
d��}.��5>r�T����wT�ۼA:F��{<z�M!т��#�+�Y�l��}��b�'�H�#�ͭe�R�you�#H�5*�o��5��9kB�V���W�/����k~y��̫�9�<�C·y9=��O4W��|W�сȰ.cvb�J�N
J�E
���a%�e��|鹸�T'tnf`��d{`Y9��g�_Pj��}sUE:�5i���+*k�mD��Ͻ���(]3�
�\��h1�����P�4C	��q��D2��+����j���$*���Y7�Sc�Ѽu�w%��{��׉'3}=��j�e�R硅.V��o�ӓ:
@�!n�d�X�߶�L��P���OT��Q���a5P�U=��3�)sJ�J�(�3a��V"P�[sn��,:��]�9�٠���f�o��֌��<=��U��SG`�Iۜ�r�Jn��Q����JZ�5�Q�u�- �T����k��;�_����oC������i��v�Q�Ȥ�\h8�s�Lʚ�0��؀�:\��9���Ц�1x�8pKwe-yS׶��U��2iR�=4'$y+���/)� �/l.��xN����&���C��N��Ne
���ԙ<J��:�����~��c�e�<�����Ԩ@)�1��2��A�����Yu�����%�RW'S��:ۦ�7S[`U��,�ӳ��0v�j�k��T��V���u���Ώ�CF^����w���1VRV��rGCH8<�6�ʣ�˴e��<^}�z|=݄��J���ں�R�*�3�j��!�X��3�AާW�v&GQ�0�;$*�Jա�{���o�/Jch�u��Zͫ�Wlt�S�;:�Ek�^Z���o.r�Z�r���	���p�Q��}��ժ[��:M��l����Tİx:X�
�fq�Kq�
����\ �� z���iy�ݦ�)�Q2ZU�L\��ޚ�H���u�P,d<�B� /ұ�U���q"��s�6����7qv�_�ϲi���eh2��a���rD����2'&{G����ȸ
�{��j�kw@6H���Th�!_���f2j��-nНYV���4=D�Oh���O��3�5~��'��)�:4�cơ�=����ɵ�����v���Lu�D��oR1�lo�l�'�y�R�����`��І�[إ1�T�}�ّ쮉�����Ē7����TîZ��G!a�
��\�m@���Qi{L�җ����B��^�z�l�*�+3�涏���)�l�.�*z���!8f{'Y��3���P�r���m���c˴A\D��VZ����0���d�����w�����aEk�7�f6j;<l'�me������$p��̄q�p�S�נ�o4c�hvm�s2��I�]C.z��"s�QwU=�͊��Z*@�]�o���vn����b�t�;\��g`�R�����������oE�\��%��}��f�L��%�!n�xq=����D�݄�������
��^����b�;0%13�0&�@Ns�h�����lA�]+�нG��_#�ca�:�1�  �!���I�� �Ff՚��}��D�&Y�ظ�JxlW��X3�TWV�b�x<�'��dݾgd�ޣN�).ojf+����E�d��3����������MU-��ک����K"�2�u)w7��v�دT b�Hy�\I���9���%����^Y��!��
U���<���Urh���x#+�
<tQs��3��hЕ�\E@ͻ��1Lt�X��O(��!�T<3�<(a��a��kO$�LT5�'7!����*c6��[����S!��b��a����|/>< 5!�b��^O�Cڍ��\V༃�o�fxr��B�C�9kC먖	f�sĄv�I��\>�姦#ׅ+{	A���F��2kPCLlU�	�xeC�]���������)x�d{#�xV�}�NuN)�m�i�7c d�����2�����u
4�3[9z��lA{���E�vd���N�Wu�4��`f��L��`Y��>��7��@����[�;�X�30Mm@<���}
���z"�j�˻�+>0�[�~o���>����R`�K O��.%W�o��xo�^oT�A�;.�s���eNp3�)�G��^�5�\]����0�u8a���*�.keF�oL.�cxTb.c�4��m�9����<:�<JW����b��/$N*֍�+�0V��WF��*Z9�c&ة��2e:|�R{������+�X{ʬS�R���ׅKQ{��#��f4*ZTDKlO,���׻^�Q�#�Wq� ]�.R�°;eh����Y�
έ��u�u�|�u+�詇C&Uy;R&ӓ3���MC;P�����,�����Sp�;�Mf��7K*�l�R�D�였����� ��iwq�n[FհS��U��9B:�q����!G��x�r�����)Uv 6�S�pO]���GD�ά9��o��ֈr��}�UC��Y$�(QM
&6%L)�j�'���t񮺜1]��w�S+(�O_(�b�u���ɐz��H�~��_�&��{X%l��������SW*�<ŖM��ٍ��f�1b�S/"�Tg����dkN�P��*M�F:�&�g+�t2�r8{%._G�;�[i�]��2�7��-Wg��3�5�J� �����|@ߪ���![��������Y� �)�G�^1\;qxd2�>�����v���L����R����h1�����u�&��ٳPxq�؃�j���ln#����k4�w9Eާ(��{&��j�U2�lƾ:р��3!�Nm�NE�.o������x���u5�b����]s�R�)s�C��Y6��B�@�4��&�j+��+4��^�}���b�e��0�K���]��2��E^�����5���|�]{��6�?]��y�Gh	!���Pd������I�|�1�G_��^���}t=b��)֩1%̂F��L��	T+�'�d�G�1Z���ݢ�.��#X�gNI��J�[UT��L:�w�`�%N{��SQMs���<�h����F����j�Y	�G*݇�[���>��j���a��6O�B���YWO�
b����\�����O��waki�*�u�����U��l���[�3^N6�k��X�_TW8l����W[���C��켖��k��5�vRG���t�A���&j�#v��#�؋Ѭլ��At�\�:���n.�ƾ�]t ��q�M7nSl��r�u�������<���t��A@8�w[�ptw�g@�V)]�7���e�l�2���Ӥ�@�z�&ݥP���H���;oy%���z����b+Uck��}o�]"ū��n�_���<�nYn��)u����N�V����)��u�X���� ���l��K+�w5�>=|�̻q��{��u1)�F��%��K��M��{κ]/%ݶ:D�ѳ�`�v,m�h	�n�ṋ��nᣫ��>��;�����k���
\��l&�u>�nX'�	Ѧ�+uj���ۯ�6��6�yV�Y���dL�ٶ�bY�z�����y�x�;"��E�KoxY���.K]{�van��+����7��ѫ<��%'�ugk��1���j�[v�z��]c�1�Ng^�1f*?F��v�-�9�͕qn��F��'2""&�Mӝ%��+�K�=g�:?hV��٘�;����itNN8���Lٔ�ƞ��)���3YrW��aY�q�r�B��D��M�}�1��[��9 �=�Z��¯��o�Tn�n�P.n�㓎L�jL�� �����[�F%�*$����Mͮm!Y/m3OUe��gPM������E�/s�ԥ���v޸��RA�� #E�y5��[rl�ֹ�P��m�ү�$ohT���a��w�j�]{�|�ذ����x��ש,�k*��T(����y\�S*�����s)�ע��;�>�+K���8�����5�)�,1��B���ʧ�m.ۭ���_[m�b�XL��4�� N�6wi���͘t��u�F��>n�wB��k%op�qt��w�sber4r	�Sr��#��z�vƕ�M�C4�.k�uŷָ�T�%.QWpx���ӽ�UNLɼ�X�����6����{xNB�g��7��e�e��;�a-C�aOk8�9%�V3�L���X�0�x�0GfҊ� Bo�_\�[7Rhp�
�ᤦ����ή��Va���ã)��7iR��պ.�����q�,L�Gm�U�B�ֶ[�Sed�"l�ysK�F���u��72�@{�d��[3hP}S�U�S�7eYi5Z�q.�CC��_m-�7�}xM��p����f+}֪�j�����=���%
�r��%tC��]{+����\�Z(�i�%�_4�=���p��R��"�Z�U�6"�L���J�T��%&&��k,b%�ED+*,�a��jE��S2����e.��hQĬ�ċ&R��(9LB��b����DLE��EJ�PV�X�UJ�`���QUĬU�)r�6��1ݦң���6�6��E5�1��7%�E]lEMev�m�UV+&Z��`�Ŋ1�����Ң*"��AEE,Qb�dY
��Va�Wm�U�T����*Ȧ4b�i��2вe*�b,����� �XĖ��DX�m�TEU����U0�f�Q�DP`�*"++TVe�)DX�D֊�\�V
("��*��UQYQb�F�ň���""�)*�ʨ��*"��DX�T�F"$ƫ�AUe�����N���,�r��g��e�(�}9�7�{� ̨�+y��C�5���Z�C�e\���s��l�ts��M~�f�� s��9�+��fdƺS�u	s~���~ ��j,�'���uhv���E�v���L9�*!yVwy���}�����:���c���j�ޗ���<��v}�lF�0v	�Q��.�2�����C*ƕ`K+^_����#Z<����>�,�*+��#��>z<� �%�&��������'\����`�LwlZ��2%���LTQOW��'��_c~{�Io����\~��L �4�����6�4�0�$k�G��3c!�*Z� �W�A�xX`�-���:Z���/�:B�V)"07�f�"}e�2&ȎE�[�+F���)���V"g������B#��M�<gHK��V�����ڀf9kfM�m?,���b�4�;>0�xTi>8�Mz8o�!�{��<��	}w���3�*J6�(d�ٛ���l�^�K�)�੥cF3-wb�?v���Z�=�o�N�]�x�hZ���e��Ek:����<t!n�Y'z�ڰ���ʓ2ST�w���V�z��0�����^�gl7:�j `"���#BbgS��U���rs��7�(N7].�pOu� -P4�p�Q�~.ErT�·���yh����b��*U�׳u�w�gЏ�W�!
��H���m\ӭr<���EƏa�EL.�^CU=�>�@3��ty��sƺ������M4���*�8�u��*q�ӝ�m��1��4�Z:R�@(42C�3ڥ8E,�6��fқ�f6T���U��T�\BW���m2F���憔U�
�)�{����0��$r����p���/7���+2?9b=�ğ�l�t}�p|��3��Ec����t���]C�1�"�-e��V��J�0�ouq�/��@���^K��P�8)�,*/��x
���SC�:M�N�ًۣ��[�y&���U)T�T6fzj?D��RY%z��W���AX0έ��'x�v�7y�NNT	"�ْ�� '� J��Ga�G�^D)*��*��wD1�nܨ�(�ɀ�YS��P���
�/쏴_V���ǡ�]9�b4��;�xat河�.L{�^:�z��� �;�ūCNb�Â���=��4i9�۶Yz��E,�c�]�[�5WԸ\rby�P���GB�o�95�77ܙ;���ɇ ��Z933	E.FvE�vd��R��\����]�� �?�Te���JP�@�.��"�Ġx)|��0Й�Y}�ګ����~�~��j3d!ޫ{+�FxS>���� ֚���_���YV�����5m��_QG)�$HVjPd�؃X���	V~�i�#(`��ܙGE7����>�<u��?z�Y����G�ӣka�p�V��xtS~=P$NMh�����ת�6�>f��nA�,��Q���><�a�{	wF�0�pm�6���M�����g�-�}o��M7���ׁ�aM�8��6&c|�t�
=���8�����C����\˱.��=��+�cxV"�:���IӞ�
�A�E�#-޸��e��0L��`r��i����-�k;5����X16��B��j@4��Y�X<.�ʬU�PZ0z����e!�EBf4���4��}�)h5+��r�s�V����r��)E�
�
��c;jpO�S$���ب�1��;�e��êGi�oFd�^�p�#�&`��XT&V�_w�������]�;o��GAƹ�t��鏝�qf�p��Eө(��s˾9V]A��`��q,^���n�9v�]\�`��;��h��F�)V�x�x05Z<qW��#\�g
�ʏ���w1�3���2�MBe�y�%d��L�4�p���X5G�ٮӞ��W��k+�i�(�t8��q�ӳS`F�w�7E!�i�*v 2q\4��&1�E�����%���n{(Z� Ņ.�d�%
#�i��W%YC�p���s�s�Q{��ۊ�%K�cf��sǎ`T7N��0p)��ʧ.��1
s�D��֟9m��>���<9GԴP�Uf+�n�����}|=�L�U	��@sH=�}�Ν����y�@F5�0E˙��]fF3Y�/،j�}c����q};��ϔ��
]�VO0�d���bС��mѕٷB�&[�����jFQ-�����H �5�h�r�׃�jR��9�ͬ�I�!d��JG��W�T6'���݉&K�� �N��~����|�i���3�s����S���	��K��U��:�LԊn�V�G�

�>�w�@D����s[���xB��N�s�:��+:�v��t�(^R6ؓF�p�;�V4���8>6��M��t��Ţ�V���n�G��f���b}D�2��ز+�VC;����rp8��t������Ge��액E�/9��MC.s�{�0��'���̴,5P�	�!t�hs�pc�M�_��s��%;����7%rɚ�Aō�1�]�r-��{��SXL$��fQ���s~���:qLRF���sc6� :-��Ɵ;g�-Fw�������yY0��t�9V/+-N��=�ġ]0i�����Ϯu���6�̡Q�ϩ	��t����._:�8�I�QY6(�?P�6^	�t3a�5��5�<�Af6�'s5�}�{�I��fS�\�U�z��E�h�Mz�\Vq<?_��RP�K]�\קݰpjӧ����n�$:�A�|4��zܳ��|v�b)��1���q 9l^]���@����^Q?xe�_ NC��M���PSVm�A�=��S)��;��*��s��>vɆfQ}U'���:}89'��:󠭑,�Y[c��U++��X���Jo��\�����EP��Sa��j�v���l����h�kn� ���t/�c%�і}H���[��]��x1�K$��%�{x�����;�$�|�eFP��W}(�gAn]⫫�&R]�c�:��7��b����g�0���H����13��6��fd�\�	.ԙ�3�9�*c4�h�˭>��S&4R���6|b:�--�:�7nAҒ����w�Q���	������$G���y�b�-��N�>󚮞Bd3�sv�ԉ�Dz�Z�Ϲ[����K�)���V6c��wb����SUOk��mƻՙ廗<u��{��L>K�O�l�*��@sW�����[g�`Dӳʧ�l�U��Ţ��C�c��U��mT�7�TLנ.�J&f��
��=�!Ens��$���v\�X�Ҧ��s����v�3îY�W�ѻ�8���]^���m���I�z�5m)�S1�P�N�0�͵tg!�vf/ӳ�;�&�R��Ǫ#�/�ZZ-�0�7 {�){�^U��Ygf� �&�E�%XƗ:���&��_�)ϲv}t\q����d��U�#�_g�y�Z�Y���vgK�]�'"�mSfE�.��!�lE�Q����쫏]��ϫh1�&��ޮY���{�t�f����:�0^�^�s��pf:-��k'2q�#w[�VP���ֶc�ѵ��ʙR�P/ fu�9Ӱa��!����1��ā#�>'����M.jS�"S��$�>��%�����Y>T�eG#3͙���� 2�W���M�l�#�ܠ�w(���H.K���B�iř��
c<�3�L�N� �]$vT}�:!HU�n]۳�*���ࢃ7�0QV��}o���H� +���۪���ObJ�c���ѣ^6���ՕU�1���F]C��(8P8�)a|C���"JJ��[ӽE^]q�h�ra;e�3�Y.W=�?�ィ<)|���7æg���/D¬u�`�/M-�M��P]�B���1�l���*�3GN�T�7>K	��=�O21"WU`K<]�Y�>�ei�W��j%z�U�z���hY�TC�2]Y��q��M��9@��3vz�����B�ʷ�!�����J��JIAC�R��&����-�N:���Ʉ��)SQ�������t��)�qY�����B:g�ǩS�ve�q3�|+"��q]�A�G��7!V��1PS�W��rפ\����#U��0f��g�%�f(�a^��8����W�1�}�ݫͨ�2Q��9�zouvh�ն��K��O��]Q��Ec��ÃW:u�#�S�]��X�����,�h�'�
э�^�\�^��)'nr$XD!��\In��
��Np�z&e��^���h�0�ix"��hLk6X�6���qL��Q�+�2=G��^�ͅ���X�#=7:����Rx��s9���tJ��!��Y�8EM��� ��!ȱ�]B�<���ݾӦ���F�-�3Lh!�P�5��q��x�w��5ZW�:w�rp�Wf')=�S�; �,ӹ9����=C���Q����J�������y�&6�:#�Uf�'�7��������	� �F�.�iN�L������)�+���+�g�G���r���c��*R�s�T��:(�Z:���7�44�J��|�-�+W���B�K�h�/�ٕ,��>�#����T�9��
d�S��ЙXU���Br���x~��\��܆̯�G�h�}�����.v��1���}�`懕��&���^�5�t�Vᶲ��p��",�;���&�|*���&�xdX7��ط�S+W	[��e�ۧ/u�{:�l�Tr��U��)��;p[雈gK�GX���r�U��e�B�XM�#BX��J0έ���h�I�M5w~��� ו����\M{�0Տ?��A�T�Qg��Ag��_vk��(۲&�>��J����a������E�
d��_�b���CD(�/ۃ�d��P���08k<��_:��ڸxO�U[x�o�:D,��<*;��@�9|��uW�!4Ǩ6E�]Z_x<�Z����7j���|֊.�\UnD�����g#��������2P�V3�5����V�¬)x!b�D#��@mrnU���"���3�q	�����2|;>�ZǮRۭ�!��j�x��%sꋻ�>�
a�U	ȶOJD���a'�32������ϲ�
�[������C�������=����EQ�ؖZ�|a^VL,Gn�cP]�n�����9A���t��0f�X9ӵ��q����@�y��M͊J�7�Gy�"Ǟf)��:�k�y^^�����܄���� ��uHWf���c��ov�|;�B)n2�-��W�uڤ���[T�O,��Ѷ�KC��������[�*F���"������x}��}D�k*�-��ǭ9te���N뱤��}Y��n�LeI�K��ռ�ޥ�",�>�d�SZr�g!�W��;>�7B�;­,Qh@�}� YM�9���i�_|`=��Ո΍,3��ȬU|��}��кo*�5=R���2S�a����$K�	�es\*�X85�����3����]�>[���FK���ϗ =M�?�J�l'[��*�~Wܑ%x:󡓶:z�2DY����f��kb��Cb�V?
U��b�C�Mr��YA���5�=b���M�'�};÷"R�y��Y�g�ʀ��z��_��禡��i{W�7�X�k�)F���rqhx�a� Xs
s�i>�:r889��{n�^�7w�R��0�'�OV	��/��@���gP�r��z���Z+�@W-ش�gs�ŧI�������̫��j,9U[~�k-ӏ��My��c�@�~��/�mJr�̀z�Y���f�s�P�!K��,��ǰ�s
���p�J�-�к�(���t��G��^mFһ��-�l���
?1ղX/��Zl�l�}��3d�JV��A�k:�c�k������>/v+bDu�u�ա�+h�@�t:m����s���~�q�kM��w)�,`��"�ڝ�Wf�4;]Mg"�I��4ު�Y}a�k���K5�:y�H��;-g{�7Ɯ���]l��ٜ"�a��pn��Ӟԭ*���o
��D�� <ŝל� I�-�y�5�C;)gAO���Xj�I���U|:��)�+`5���v��+�.�z�TXI��$��oVLWR8+<�_NG6mt��7Ҡ[N]���ٔ.TFAx�Rpa�v��.t���9M�	�o�wۄu�NH�q��x�/8v�E6��Y*e�f�
��.-�BN�&�C&s��n 5��
�]f4~v,ROY"��ǈ}��)����o�ӀS��� e;��.��8WT�K�=�����wV��u����/_u�J�h�����ʨ���R�yId����yJ��X�a8.���%��Ax�3
���H�X%�vz���ѮҸվ4�_FL��v�;��TaG;qj��6w�Y�7�!�R�96�W��9u]��f����]�l�!D���pV~�����Ѽxc���Xu��֡�0��EV+mU:�<�%������%�V�ˬsM�^�؃�6���77�m��U�r��0�r��.�+�}�Č�b)0��Y����]�2���,Z}gK�-�:�lDf����;�'S��+5c���	��j�j�4̼vt������ַ�kb�r$M���������r0�U�Ԝ�m_h���5����uu��ي�u����4�bcd?�Ѻ{��} #1�M����)�ݢ�	�X�uʝ*��X���������ۨ���z���ZWasz�E-�d�,61�>5,�ya�C����=�*Z���+e<O+#p(�W���s�j�,&�q�f`��9�-KS�;If�Y�n�������c�#���Dk�|��K��������ˍW�;�I���,�y��E륯o��0��:an.�0�s�y�ջL.g(@�wY��+�*vV@�r�L�Y]j,Ѕ-b� eC�I�˽rd*e���SU����`k�Q�4�<�Z̈́s�TE�y�b�'S]����ѻ����x ΰ�ԙP_i�s-]�i-��������/�W�N�2�{<	Ӌ(_k|ӊ*jm�7��@ C��Q�L�(Gݶ��*�I`�g���P�|����&'ZT�hPF�oZ���Oo;��{9��qv��/&ԫTz:��Ek�ξ�gwE*�2�A�֡�*��K�4M��� �|�(�1�**v�,1���b�EQTQb�PQ�1DDPUX*2�"�f�()"�

�,u��TQ�R�!R���Q�u��6���P�Er�Ub����*���f�b*&Z ���X��TPQV(�3-��m�̷T�V#AT���DbEV*�V(�TEQ�,UX�����(��Gh�Dc5R��S,�R�Q
ªjɩUTRm�U"��b�aTD��b*�Q"�9.b,�"���-���2��VTb�)m*cEPEDUV��`��TATw1�ڎ�#�&Z�F*���,��Y[��(*cPv��"*"���]U�AU����A*�����"������ƶ�A�����/��h�U�
�w}�7-d�4Չ݁��m��e@3%�7�m)Ev^�WH
�mE�˘��S[vo�k7_굃�E�嚯</ؽ9�����>��g�\�Ҟ�h7n::�S���;�+����]�:�J��)�f6i�w�
\�WFr�f`�鞧a����%|"�F�S�B=�YP��vוA��.;0&�s�D̳coj��ۇSp�5�)�F��q�u�=x^��~���=U�ѵ���i��q�ڶ��d��%�be4}�ā�Wi�,x`�8)�,\��=tR����jm���*y�Ĺ��Sv}n(+�\���f=;���v�E}Qx|/�`���I�{�.�y�+�9K�5.��P����D�TN� ���Ga�G�@h�.�@+"���4��f��ѽ\��>�
p��8JQ���O�s�Ղ��:��t<�/.tK�z��p��7���m���F]C��J/
ʦ7��W�Tb����r������^���8�4\�؃W�
��S3A�as�:fGR��T� ��p+u�]r��-]��9�,Gk��Թ�~�̍v�wv�'�&qT��1�Ci�`6swi�­�%��H�>�A��ΈX�.*�[�o�n�����%��-���".ɷ�lD'+�DRY�M��3������"�;]PV��9�3;�%N{RŐ��K���- �Xs��r6I��{�qwuZ��{��"���^c�M�b{��=�V����|=�.�Y��y5Ӈ&X�������-��o&�o��hTGs��VO��k�����Ad6(���*�O�ׇ��Ppw��G�3Ǆ�}�x�\��5τ^ή>�Y�@D����c
�Vc�'�#½����9	'np)��2�`�o"	�ЯҌA��2G�����g�յ
�8��h�-9�gJ��Nu��%F���5b�CWH��Mwl.�ʬS�Hc���V>���3�#s#+����F�;�
�嫍y�N(W[�� ]�:C��<)�
���mRY�Y��U)4��F�S�D9�9��J܉��̢#g�ڇd�����˛�:8�N�g&���
{��XyJɈ������T�;�{�m�棦��n��x+>T�VW
���۳EE�����w<�ws���R30@��D�}�_5��d�(-�J�}��+]���gP�z����C�Ҫ�Fǯ^����c��
�
찺��P�9�)���b\;�ܒR�=#�W�n�<�8��qJvj`�d0��:)�+ӵ`u�oWL����$���p�l���S3��0p{UJ}2�f'��p�V�����q,�/�.a�P��#f��sg�`YwE͊�8���_(��ϯ���!�>�oUn���z���Vb�{,���Ά;�Q�6��t5ҕO��6fQ�b9*����P�.fu�b�!]6��	˝��g��o;��lHz��r`����A���MW7��6oӯ���Fɹ��DƂ��J�֚�Y	G�Sd�u
T5�h�r��
|T��1{4ܤ�ա�ʁ�kp��v�$���=�T�p��,��/�5̩����%҇���s��[�4䙛=Iz+�M���0:�����w���|�އ�:	V���:�o�J�ed�x
�tݹ�r�MDb3)��B�'�d�G�1Q��]��פ2�IU��^#���x�^�t�lkq�;YCZ*+��w�c.�2fl�Aή��>h���,�� �#^���<7��VoZ��ƆAr�����kue^%�Ժzc�����ǚv,
3J��y�9JsgV�8�s��hڋ�-����b�9����,`�%H�G6��{` r5�/gsٖU����(v�ܼ��
j)�b����O��^�0�+3�,�'d{�\.˛��Z2��.�;w�q�D��<��X)3� �N�S�B�9�FffM�����Z��9^�<=f�?U�dp�;�S���ˉx,V+a�=���0��{����.z�5u��)���e��ϔ�#f᜻s�靖Yg��c�L�aV�(��0���7��v��"��U��n0g.F�Fxht�?�Zp�TV��X�u��S��7��s�u���9Q^�HrٞUYĉ|�9#¦%���b�)Ҋx��j�yr �=��m�Z:9�"�I��.9���j�R
V�㊦��$�p��7��+n�V_u�j�l�劚�\XS�����U3^�1D.���J������u׍ɽ���۾iF�ň�|�f��i��@v��``\k����mF��z��S�&f
��feF�]�d�Kx�sV��-�<X)�4�F�o�<��\`�@�j<ʔW���5�S�I1��1�Vf��-��|*�'8�_a��]����G���_KW�Ι/�uu)�̫��������}ʔ5Y7hN�B�w�D��@

�pm<ϗ	r�E���B>��'9N��]{S�f9�/�]�K}�3K��敍�p!���Aus�S���G9]�����*^�um�G���Q�:����v��SW��!�*�7X����Jo��
�9X1�\��0�Dpx�J�~TL�]^�v�jy�Z�z���z��5�׆��Ϗ��h���8�6��n�}�\��D��y*8'HK/j�K_��<7ꙏ� 2�g���P��6��#ga�vaK�j���d�p�r:��L�%�F��91�`J�y�%q6��@�eB��|��s���	7kʄ��T�z%O?@�M%��U�~;5Gq���{ \=z�����õ~�U��+��7]7 �▪{�����@:{M�(<%Â�,\��=�+�P�7��~{��|�& �|�<��TJu3����� 3v�+��&=h�J����E��P!-�B�/�}�~��/hh���&q�d�Bd;F:]ԒH�{x��X�c�Bnk��a�cc�u����n�Mp��U;���k�S� ��:[��W-hJ8��J��f`��j�(�z;�Τ��fK�z�B��3�V�s���|�s�!�D�T�@	�]$vT}ӝ|V�s[�B��X۰ �&���*�������t�P�&aLB�⠅$$��&���{�d�VF�(��>�T-*�j�.���JV/
X_�P�t�*0N?_n����G��"�y3��es؁�LR� Ϻ�x`�Zs�t�gn�r�z����w/�5ǵ�����&E`���\� �b�y���l��M{Ô������E���qe0&6S���y�Eב���}���y����L`���ZwKj�pH�V�iF��銎�OK�0��[��Ɍ�}�8
���
��VC쫪:���[@mL2M�T��&1\*�*j51Q�M�=/���#���������Nq�������0�d�Y�U�n]�"��~���]��ڥ��u鋝������oR�&E*ɉ��s��,(b#"{D���Z���[P���U�Y�p�\�E:ͦ+�`�^M������ԍ����{Y:Ɋ��3�
IT��5�X&�ڇ��.�S�J��3:�.��%�i *+o\� '�GJ��QU��]�)v��4��g@��)U�Aohf�oP�J��[=|�f��{�g���9@	
%M&bL	ݨ�=;/3�J^oE�Q蔩��tէ�f�H>~#��lƁ^AKZ����1Q̴,	�F����A�^�j��p I=�˷G��0P0.��*Y� �v�+r&ӓ3��hu厼��� P;�����B"5ި�X1��l������E��bN�j��gI7mU��s~��6��9%T׻q�p1a�.����L�`0Ўh$8yM�����J=T�_�?��8]5����!�D�P���'��oM�~���������C�U����Ԉ��ևu^y<%-R�\Y�	Vi�
e ��l]P���ʋ읱hL�O�=Ƌ��a�+�S�:*��m�g�٭��2��8w����z��<.�
�p�R�3�^}�6Q�Q{2�"�/<�{���v���^�`�N�g��/1�D#K	
��J��N�OZ@�aU�B={*���\9Oogl�">8k��V<_��*�?]��9���֮������8�Avr���r��#���)L]�d�w���Кk+(��Fk�)�4��uc��ه^g[��Fe܆�K���r\�7Ug����6�;�Q�Z�!�ym�vm�Y>>�(��n9Ahc�l*�-S�v�V�ά���WP�g0�³m_KH���սz�K�����Gu���uT �T�^�n՝M�يog�b���7U]k�}�YM�!hTb��"ZR�2%1�S�yL�%���IRK�x�=�{��e�jض��U8�}4��s'��\�*�S�
��s��U�+B{��u&(u�j1V�wTn�8�C<��9w�uԾ����f��)�N5zӞ�["�-˭�ǚؚ#��u6z��uxq;�U��Ω|��q�p�ॵܷ�S°�C���iC)3���Ŏ�Y��B��:fyڗ�����N�m'\Hn�@ڨ���e\�X��.yJ|v���R~���FwnoofXĻIO�1�mWe ��Zk�Y�P/�e6mai�[}�G�]��3)����%µ���};g4%� +m�
��WZ�|��2����6C׍��iƺ�6��;[�_8ErDeݠ�Q\����q�N�1�'j����:� m_��fގ�\�x��s���j� �9oC�B\j���gL�8I���;��<�]`,c�r�;]�iPv�C���ʍOh�f��f=�y�~ף,�Rz�#Nü�L�緝4�V��-$�%3���gK��Cg�����`��,�Q��Ӂ�~�G�6���o8��޼���dj�-l�xR��(gvΌ�3�� �15����^�3��^�;�E�
r�����g�HZW��7iob�ԙ�WQ�qϺ��TF'����O�jT�}�����o�ӫ�6����F>��������U��$�\!s�k+[j��;J$^���h>�,�{W;���+5Qy�5�z��u�e�=��3iʵ�I�guK�9<E iR��1���˧�Ϩ\l�0�W�8�z޽�O���okkr\��8���D�h�O.��S�Ǣ�v%*�*Д{Q��
��nj�F`��ϱ��*��a[�V��5=!2�����{���$�8,/ �nQ�8���o_GX���Ts���h
�q֭d��d�����Sڬ6��_��TD�{*�)��=��� Mv�C4�N+]P\��܈I�N`���7��5�Stw\l8̛�m����ZjU7����s��S�Ӟ�������j5\>�?���[`ns��������+�[MN��2V��q;����{	:3<�@--iQs݆�B���KisyW��-D�����	��]@�U�-=��ciFP�y�����Mf�J�;CK���2�Wc
�k}�վT���
���s�w!w *n��X-�Nm���2���eaP�s9cAT��R{9���}ec�W�7��Ͱ����3�?EA�ރ���٩C:�/,-�+iHې*Go������5���F��(IV���e�+���VWwk�Q%d��,澮�mV�i��f�.�#��hз�������m�yDJ���Mv��!��)��ca�)�X$=ygVyu�mŸ%
t�z��c��������m�r˙4˰���v;��-9,���:]�u�^A�J���n(�)R�y��,�0-��ݩ��h|��Ub�n�ʶ�s�	g�Ư��]��-J��/���[9;.<��zU^��1ʺ�>n����5{[����G%:;o"o��,1F�V�qhN-�U/�!�Ӿ�^Џ0����e��_Le�33�1H�g_��P�=_*D�9b����g�$tD�9��vzv�K"���˔-��\���1?��r�Gk�5;%��{��V�ވnL��c���g ��Bq5����V��l�b ��P���^������硼�0Q��z�oX-V���>ޏU/.�������Py�J�{d�b�/C��;���qWwPٶ���ʑ�HX.����V?�\:/U��w��i���z뉎��R��q�.\��Õڛ���JP�Q3�r��HT�yɐ7��m���tgK����g1���}b��J�P�����n���$qea�x��v��\�ɢ��� ���L�k+���<6��SOk��rd��]�������h�z��Hc1*��7
V{Y�#�2�U�gD֬2۳J���J�p� 3���J)x97���L)TI���z99s#��U޺ɸƐz��������᧜-+p)¥��d��N��1t�}%;��pX�v���-iAF�r�K�sja]�lwe]#,�>|!�W�˸'��(�lζ^&1a���đsAU>�X`b�d7�!K4c
]n⤵n�����9�ϛ���Ѵ�`���k�yDK�_��u����u�gdC�X�;�e�uΕ��;�,n'ZƩŽY*Tؕ����/�;]�����a��)ێ+��ߵ�������J������b5�tv�gM�S����o5-�
��Sxnp�8b2�-6@^W�����/,o!���"�Q]9:�ܽ�,�t�)M�y��n⹌�Ȝ�jb�j���^4WM�� F��<,+(+�65�](J�W��F��(�
Ƶ�Ƅ볡��3yk�:���He�J�J�]6��.�4p�!��C�q2Ƕ[B�����%X���j�3��*� ڎ�%^#*��j�>�՜JU�#�Њ�zl˃��~�"�M֊��6,EDTA[ZV�A�#���"(�U1��*R`�c�EOhV�WZ��[FҨ�w.Ң1TE�TA�,DEu�T��(�y������b �b1X�U��Ek*"�l啂cxы������Ȫ�Y�,N5�2�8���Q-�1"6������UQQ`�����-TPEKe,b
,V8��1Y�������ڨ��<J��DX�X�L����u
�EQUQ�1��La�P��X*���+6�Ac1A��AX��\�PTQ��u��
�lE��l��TG��DU��DU��$v�+h���y�/�s=;�r�ԝ����۽<�hvMJ�����-f�ݕ($6���6�hː�t2���Ӻ�p������ƶ�~���Z��<�I��x�N��97KZ���M��٧�5��:�o������s<u��+�ն�/[fI���p�GOm����}���|�h�F�E%k���9\�q�)�F�J��틞;5��^.�F [f�D�eO'����U��^j���J2V'�c�7j'��]����ZI�R�����v7�*j���dsj�%�y�Q�w6�4���o.,.n�@�w�ꠜ��JNM'0x� {5,���Cڱ�na�S��6M�5���9˴�'0$���`�on���&���U ek;����Xjðu�k��p=B��f����q�OȮ�i\��i�|y�{�Ow��./�ki���R�v9�=�.e��zM�CZ�bAMV]�w,����ܤwn3��Zi�w�r�LfFy�����E��Z��'ՋA��Į�F1]�u�1�����.��ӻ��kʸ��E�����36ʅ���[�Q�ٷ��u8�Tj��v?,�8�Jwm�N�l+�\UaҸ�<x��!�:�ڂᄤ.麅�7��� =>���`�|�j1�J(����b��=���j���ו�6Q�Qg:�5iX%%�U��T3��*�h�����G_7����ڼL�����3SDk�v��М��*��1���j���U���Սq�Nj��5���B�y�s;H�u�Uݜ����j�����Kv��n���\�ǃ?W�Sw�W_Cb�&�����FcL�
��O����"�1����A6�����-)](��!{��ځ�d�A7*���b�*罋_c�ڵpŰ�]�o�k���
�ݐ�T�W��k
7'�7M�Qx�����R}:6�(����"����k�$g���Q�N�l����쩏΢m{S��-3梬�[F�t;�;����;O�`cv���]`c4b� ыs�u�~�q2��^l����J����v0�j�4��|���^�J�Rՠ`R�aȯ�p+[2wU����f�2�?f�߯�w�u�z�z*����ɭ���4�T#7I�5��l��y�\U�N����l�u\ڄ�ҭ�	V�	�fPi9�������Ws�1c�@i��K������WI�)o�	�R�WL鰲�e\���	�QN����J���M�xJj!�uN(�(-��uaª��ӍÙ��]���;{m���#u�t!�\A�S��u)��eTu�Q�]`=���5t$&/T���̪�X�XңJ�[܇�N�t��m�*j&��8���hM�cE�Ȫ��L�宔�O:t��j���칼ei�qK���P�N+c3n�FD[���^�wYI�\�A�/ou"�+]c۵���-|*��B��73�u%��.��x�����rZ�=�B�������&^aGgMf��@����P$O^x�G9	W�w3'�'�݀�(�	7h���-�gc�,���W-��s
�R��g��3�tB��ɶ��*FQL:r��Yw�l������|qܜ�T�W��TcYP�u$�f�y�C��uR	P]����ib�Q��T8����v��瘝�z�Ů���T֜��|U���A��"
�xg�f�]��Sý�Q|�޼-�{;��<��/���D6n�/\���J��oϧ���L��k<��'�b](gGs眬��Iջ�A\����*K��]����KpBu�5o�j�Hm �q�撘���`�Wg���zS�Pb�
�i<�9��T�:za⪀�Ɣ��N`�q]Ln;9�r�v2����<�A�~����6
:�S�CF"S�Ӟ���{��\P$���x�~��~ڰ��nk7;�w(�g��-�b��3�
Xř3ԗ^�˶���3;�����p�ȫ�X��ao�Ft-ܽg�N&0Oz,�o�V���q6$�C���X�A�\������zF��9
��ALȕq�+0�aUr�]*ǣ�:j�_P�vj6w�m��-݀�-\���]d%�w��N��m�N�U��3:��}ن4�p����]%�^fz� =t2�z�Zx7Thc.]3s�2��4͝�1n3�-)����xw�,*�2ޯ��<�H�DF�t�@[���R��-�Nmǁ| _��V�K^��z��t|K�u�}E<Cp�o��w����6�A�	1��k�is=�����<�T9��	�Z��I�w���N��z-�w��b+�^m�5�]A�41�k����s�R&�R�4��r��A2qk��o�2��_�mk����.��p��t��m�[��A������m����KF{`����n�1s��xD��+���%��y��z�ڦ�Q�*��F�27GU��w����C���1Y��3	�I��ri*9�Q9+��t��.�ٗ[�\ss��/�,�o"( W.=T��jIɚwC���m���̢]{@��i-ޕ��w�\��]��X0�]R�R��m�ʱ�⍱ۜ�����E7�u��Ԟ�sR,�ą�G<*�`��,wo�ك7���\��!���n63���q�9Ȥ�(�d�|��t��ۿo��!��C�̻]��o6�VCW���΃����:7iYK���
fʚ�_PM���nr�����[�]E�l������� �j�s�vgM��k+��a�Q�p��b팖z����Tm�L��4���lr����O�ݼ�v�B�`s��΄�R�)@�Z����%5�n�]�]SU<A|�?/&��� ;����U��Q�Ei]=K#���I�W7��,;1#�@��B�����t�Eb��Y��Jo�mT3+�h��&1������՘�$�ڀ��POaн����ϷӼ�+�ͫ3=����Յ���O:�8�����UNM{���ܥ]�`��۱�F�F]V��;���=�==5ov����n�I`epV�q�����=:)��f����2�'x�~�K�V�(pG|蛙�� �I�i��r=<͂�S��[�b�>�`�>@3dv�}]�٘�q{8�Q��:�hodr�6ێ��*��(���9{�@N�k��^���Q���ŧ{o���B�%Q-*��&�3��.�q��t*�V�D[�x���c~�gͫNi�Ӳ�B| �+��k�V�N�2�V��V��]�o;ƞ��L۩UwT�A���rH�����U�+�4�%u�ϻ4��)袄Ҏ.���JУ�_I�^�S.��k3��
���6+j�ne}�C�ٱN͡����i9�;\�Y�~��Ō��ݬ��"��i*q0-�rU1�z5F�Cp���jVU�����׫�kNӋMʀӊ� �Y��B�!3�Lb�ڤWe'{���,g�Qcr�b����^��@�-�(Ђ�v���f�ԙ_G�-x��ϼ�H��}[���:�`��h=��kK���΋�g2��Q��sF�wLΚC1˵/b�V�=B5�Y�)1W:up�K.�%�ܾ���W+Ew;��[i��p_v=죑7�-���&΁bTv��fޫi�YE����Թ���5�s5�s�,�]�3��G�ךTm(1�V����I�s�SD�V�i��o����Nþ{�e/=*W��ތZd�-�Vl��8���Z|���vx��L�k�#<�f����������煙h��ϼOܻ<���!�}������&x���� ��WT\�u��(�Y�Y���.I�q�ƭ�{U%�VfM���[��١S�%R���畉�5{Ū�\3�Q0��D�;<��1�poiq7���ĳ5�\i�q=3�Ɵ�y�쾌=�(gw��X�O�ɇ�/����G�W;�\b�U��֔ ܮf�d���8y��M�a����72y+�7�o�����\�!U�%C6�Ag���B}�����6�m]�����G�B:-t�5�Z Z��:�*�ea�ᰥ�o��x+Tm��42�^��ɗ�I���P�M+�hj�BH�J�(V�j���+3-b�{FV*'B��WY:�6H��T�L�ݴ.hԛbs������F�J��cl�k��@M
4�L�'1�vC�Y�� ���͙kq���ٱd���=O`�a��P�_�s�=|�ۥij���՟�O�mu�R�YY;w/1|c`��[�ǐ�A��L>�kSY�N@S&�z�"�gV@V�*��- �<�(��Ւ#m�U�Z|�R�%�nK�վFz���H]O(�NN�kL�T�P���۪p��	)����������qbꗗ��wU��n:�e;�0�qiV����ov��xT�9X�Ov۝ý�`q�T�+-M��5,����������+Nw5hN��n��8F';��f���Z��Ě	��n��4���\�_V`v�]v�p=��Pux�U��V����=����ݤ�^�
���uf!%
��Oe�z�0�$;Z$����s݋e��`�]整�~�Ys\�V]X�vۗW�՝-�1R8Oi�ю|��i���8�Z�T�"��,�z�Op����Ý����
�V =:S��9W�n?n������*\eP�Y������twqMKh��v����q��4��-q��j;b�x��7qӱ�+�U�n��%�4a<�Ky�k�m]7l-��'%��=r�˾�T�A�{O��7��3�4RMTc�1H�Qͪ���I��R� �;s8����������)T��rs���\^_v�m	����N���F��;�+!�����s����ġ
���mاe3YS��%u@J��u
��Z��ڰ�fZ�b��ՍJ.vmU�����B+� �We�ʶm`�#/; �8%Sv��9U!��S�%pǡ>�R�TOZXκV��Y
��<�n�+sI�1�.�9d�R1�QZ&2���+�=������f�&&"����M(��(�̞? G��l��		�O��z�Q�l�0��ܦr=���+b��&"P�M��f QEA� �`t����i�Vz�>���K���m�G±)�R9�vǶ-��m`�3�{]zߤ��kp�8�5��vɽ���"� b�a�Qg+dW,�Tx��|�ӯ���H]x��
? ��@Q��ԌBJ��k�cНW��V��4`��R�����,����I��(���2��ሁΣK���D���L���,`|ɽ!_ʴfyR����Pi�Z���@�^��*�bѪ��v��z=�@y@�в��T'��^K�%���IT�P|�j>�*���xx7蛞\v?Z4OD:%�p��Lʹ�Я�:}�?���&�i��
���É�s�M����;:�,R}���.@������sx���.h}�'�x�ݢ��r��r7�*������1��k��g#�H;�0A�� �F;�*���?j0p�{!:D��(5���C���`�M��̾���ۛ�C�����0;# AF[H�ȅxM��\��Z��xE�,����!b��R�Ą�������@��;�9��:�T�����R6��W��{�Ov���38�8:s�묱��CM�%㯛ݮ<��C�ܔ����{�R�*��]�Db<E:}i�Pzց^�.P���cf���5��@i�:d6�\���<ʔ (������^÷^;���=>���i��q�Wqv5Px�͵q�߼b�O]K� �0l�܇�RA��]�~��Qd>������UG�aU<���]��z���DUG��:�ap���x�ݵ��+��R^s[&����U�R��.�w$S�	Y�p