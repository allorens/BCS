BZh91AY&SY7�X�٢߀@qc���"� ����bD��      �]j}��U��c
��
U P"�L��[�`�
((j4(QIP����[M�KT�h�-a@Ule'tw1e����S�Kh�)�T����Y,����`����Zƶl�%Eil�2E�mLV�1i,TZ1*ٵm�56�fժ�m�| �꽚՚����ݍXZ�Y7 ۍ�lUk)UJڔ��5��`l5km6Y�JF�ک���a	J��[6ִ��l(j�5,-[e;G6�&�U%�(� @ [�a�@�� �*�÷A֔��]�ö�Q�ڪ���j�Iִ��0 �T]�P�l�t�Uf��ws�Z��R9��E64�kf�6�o   �P =�vw\���V� P*�u�gC��-\q� (���4-�]�B�˛��P(�����;� �Qpq_n�W��fC4�"RM�   [���^� ��� -��w]: �Y� ���� ����� R��t����J��Z9��t�F�8�t)A@wK���v�8�%*�QY+   k|U;{��^� �׻�{�R� '�8��QܖP:wN�]�(����A���3Ň@�����IѺ ��4m5�[m��B(CV�  �o�E�Ά�S@���t�BwNT�mv;�
Ҁ�� i�)u��l
s����K��� �� YA�]���6�6��Tc	�� ���*7.`��F�*
�R����jt�4 �ڥQk4�wpB��+*T(
m�q�H���gСA�8	��c��h�! U�|  �"�M $[Ҹ����0�d��۳�4tH�7 ��0 s�‡��:k Q1�th�up r�mb-�� ��HZ�Jo  <u�/E���-�ۀh)w2�]8�P�;����vk�@lV  6�� 3��J �Sm1T�R��F�  ݝ��{�  ���P�G���v�. N��A\gp�Bq�P s�m��Lj� �n�kV�Y��3l",�Mm�   �x 11� i�  .�� �up4�����s��@m�p n�]@ '&4(�        j`�J�&&L i�&�S�R��  �  � "l��P �F� 1  U?��J�d     ���Ѣ�L�SO�&�    !)@�*��L���d��OP��3S��O�����I�G�iö�C�띹c�{�\��^��������Ǿ�(*���  
���
��( ��_�?q�g UQ_�@���1��������*����U~<QUE~�t%O�U_?���_��~�'�a3�L��329�̎`s+��f&2���&`s!�L�fI�2L��&d3	�L�f2�͙fS0���&a3	��f�2��&a3	��fS0�`s��fC2�̦a3	�2	�L˘L�fC0��̦`�s�L�f2���&a3!�s�fC0��̦a3)�Ø&09��`���L���`3	��fC2��`�3!��fC0��&`3	����̆d3	�s!��f0��2�0�̹�̹�0��&`3 `À9�2 ���� s ��Y�2��UL�#�3(�a̨9�0"L�eA�
��G2�fTLȃ�@s�a̈��G2�f&�)�s �a�*��0�f@©�T̊L
��2�Qʃ�s"e��fL��3
�d̀9�S0 ��#�s($�9�0 �W0��E��PseRaG0��D\ʃ�Qs(.eQ�*9�0
L��@��s .e� ��G0�fPs
.e̈`̀��G0�D3"$f\ȣ�s*.`� ��0 fPfD\��f2��G2��P�2&a̨��s!��f0��`3fY��`3.`3��f0�C0�,�e3!�˘�f2����L�f2���&e3!�p�fC0���a3!��f0fa3�L��S09�̤ٔ̎e3)�L�fS2���r	��f2��d3!�fs��fC0��e3	�3,��S2�����_���~�WT���hu���S)N���M�w+�TFfܽUl�i��ޤ�[��	w�}�[M��L.�/�'1�̉C�MG)�iZ&e=r3���rғ���qѡ�cA�G )��^`��Q�!EV]*�z�Yo�޿j�F�B/Q�u�V����ɼ���ۦ��T�1#{v�.�ڽ	�MGw*�桦l��β�״-7y�p|U��\m.{�Y̶r��C&S��-8�e��Y�T�(�GE�TV���B�i*�Q8��
��b��6:������o[O�5�e�XR��t�U�d����G2�͹�r�n�k��<�VͱeiH��̭�6�F�f���z�&�ܧ����B����MW y-��{m�׷{{6�\��GU�8"bel��*����=�82f+tm�¦���M�+v��P�"�:���Y+U�hM�d�̽إ�J�3--��}�p�OAnD�k!P�D�!��M��v�ASv�ؔl�x��H(;�qޚOi:4���;�kP:���K��6���7��:6f,3cU5�Wjƀ�mm\:ފ�r�x/7t8a�צc��Y������	���Jt%��j\��=owE�Z6ki�c���'aծ�XkPK0���vi��ڳ�_ ��	5Z�q���FH�j�&"70f�С��&�36�iv���e%�YqԢ��-m��#6�����$Z��k{�S��3�Cf�7U4���N��kz��VEh?:���H�Xq*�P�{�e��[R9�1[�&��EL��o-��n�b�2�K�����F�n��7W�%xfݨ]˒�k9~�ؽ��@����gMڂ�w�DѤ�i�M�sN<K`(�ڥ/5�f�7R)���7!#n�i̥�/Il��b��ۡ�,�X���f���r�9��id�l�knn]M1�s&[�ՠ~n�cEI�6�v���Y���Y��7�)�:��VtU�Z#5�z�Jn-34�-= <��2�l��e(U�"q�wh�7���O�4[��E�OHX#�S�zor�06pET�b��	�C���0��)�Jh�"�X�0K��m��\�6�,�Ku�V!uoB���9]����7tμ0��V2�9x2mm���B��HViIh�i�����r�w
:����ia�]��[k7=�h���j��ͭ�/^��v5��Z�4��jgm�D1�a���
�Դ颡��a�xf�7	��z)����'/!��j�T�yZ*2��hӀ�n�Hn=����"���^#Q��Ϻ�Cv��v4.�7X���%��VSXuVK�-�7o7L5 Xa#H@�2��Y�L�s4e�7/=.lW���ݚEXN|A:n�����Y����e��$ �� 9w��P޹(\P�ջ5�cS͂�e;XW��iּ���U���ԙ�AL�8��1W�`�Utv��h�lyR��^lP�&��c�7��xs/me��
Wv��k,(1k�V��QuK6Nˢ`��VBڷvDE=m&<�`zƬGX��wG1]"\����\x�$j��.�X�6��2#�/��;%����ܦ[�����H͹��a:��V^08��q��x����9�%�Dӻ��i��Eho�
��kq������Ԭ�	�V��	bQF�Z4��Ql&��Ae{�t�~
�C�h`�
�\����R�Y���7��5���(N�Sk3fY�qa������,�!e���V�-��浵!�@�&����sM��aR
Ӭ՞Ӳf�bx
��2e�L�h&hP����V�Ar�o"^'z�� �i�h«&�����	&�g&^���L��A����[0Q�6��R�
J
�fd��vhV��yKV밆d�5�&�F���Xzr^8�蠪GSb[�+4"2�f�8�LCn�X�7m�A�!�4$/"�A���1�Xu٦"lfJ{ej4S�.�U�Ɓ�{Z��(�q��f��a=9yh�fKV��q����!�7Fk��7m����N�Vd� zEb���^V�e����SD���n���WTk�.�cM�x�WX�=�;e}��R�ZK5��j��2
�0��Y7�ǻb��j$��-�«Ӧ��2ً��2�õ�$��Bcmi �Fc�R����6���E݅��.���):w��D�B$?ҭj�֪Ѧ�XGH�z�/%��l�wh�s]���y��ƋËh`��sv�wn��
r"ҿi�����ij63q6X��iY�e��N�>��w� Ԏi6X.,��¶nV^�+@8UZX��2��v@Qd�aF���S��z�Ѫ��Ք�b�q9{��G���̢f-1��5�|�T�R�=��={��M�a�)8�(���vlӡzeY�k��*�If�#���4��z��=yGu���y5��IytvH���JxLZ�,Y��8a1ae��ŽX�1�uu�9��ܶ�;�E�+a��$��;��2���mm��lj�M`mCw&;�� �M�R��H��g���NKdu#˕l����62�
�n��G��Y�-���6L�%����c[���a�,YL&��xK9 �V�ۀ9�3)F-���N�Pˠj�(�10�X\��`�%J(#ܛV�a�dP���g"�y��튽��8� �kqa+�,�F�j��ݣu�����4[�a'I�x�oS\�V�5I�ޅo���a�D�6�*�ú��*bB�����wI%����5��"��O�3^[�YZq��bw
���Z�
����i`|��W��\���0bHl�f+�0k)P^m�f�Z���*���ۉ�����Z�����&l��̺�ff
�شf-i�`�h����p�6V��BP�.\��[5��K�[�h����bٸ�AJ'�H72��j�YXKJ�/Y�&��:F��K%��:&�ŖR�,v�&�!��V��h�L�2�M�Rhwy�aѪ�R�0���H���p�#vՍ*ƚWv���^�ww�a���on�M���)z:[k,t�ݷ*ܲ�'5�׾�f�M��k1��7gd�zLێ9hV2�C+��=rTSb
�<�A���tdU�e�Bb6v�۽�4(K�&����*���M�>fĆM#RP��g�m�T���J��4�[T�+����譇M`�w3Aؔ��''m6mKwS7r���V䙔�*&�6���]I`����o;���\��MVlӑ]��Zd��`�Y9n�Y����V7t	��E�M�`� ��ۨ��v� d���AI�X&�^�$:����\�C�ժ5nZ݆��c]^�;�c:�����"T���֕e����Վ�m�7�zM� :n΀�ت�ssJ�mSժ�VY �ͳ�^�����j�Ȱ�[����M��Ô�Y��kv��ǉC�-MG�A,�ř4���R�}���l��l�T��&m�7e^�2ð�U!���)e�7ǵzF⎚����Ҷ��Z&�әy��"��]�uw���d-bmb)�`���3
��G�@�Sڛ�k������j�Kݠ�^��=��2�<L;�k:�x�O;I��� .�M�<�}���ĴZ|��j�Y�U<��҆$�QA�J1C �ynfM�b��p`�m2�E�d��q���q�J���z&$XB��V�+U6hm\x�J#E���V�D��I�:��7��4�����{h�a~�6�x���ֵQ��ۭ��wV⫏r6�"����0hc+&CA1Zx%�J�Mj��7H�J�]d/3�6QGufJ�$EYcr�$��ߛ#uK�.���7v��t��
��6vej*Ң�nH�U��ֲأI����Э9��;�a1�mI�e2��r��l �ɔU*xZ��h�!��$Jñn�	�C����I�1�-5	�;��8s�u�'��!6�^�J�}+l�K4+2�H���yiǱX��j-X��ҖQy[Z��i"��X�kd�9�,��Ɂ�i�5�(�V��[X�f,n��Sr�̒�)O*��a�}�GfMY�K�2]�N�:��n�*���A[6��6���5�Q2Cf����:����o����XN�fXx۫�$U�B�k�ҭ�.���0[�����ŴV�����}en�J*iz���"�6hm![�7,ĉ�sF�ZԬВ���ɴ�4�P���ú��(�cZ��Ҹp�"�B�Q�V��m�YL����05��[.V��VЁ�!���E��i�oc��4��qܻ� 'K����dBL�z��ʪ��z�����(��cL����Y~����ؽ�q��,�b��M� t�c	�����vŶ�za9��X1m�St�V�r_������wEI�{mL(Y�2��ֳL�wrnFֺ�(���e���q7�ީX�eU˖���F����SiUBg����uFu�w(Mѕ��x	)7*;�M8%�r~�H�l��p�O�/4���N4���e��"ܖu^�҄5�U�4�Y��:i���ȁ�t�K
kG�<.3m�r��!+L.-pU�F���,ʗa���[�*%����ԗ-�P�"̬�Pm椨i7�1��m�M
�]Z�OE�䤰r�7�1@�����q�@���
d}Ʃ��Z���&Ⱥzs��鱶�FtK��r�؎V���Q�֍3�F�$�p�5!y��5Fa�&cy�G�6іFȪ������c��t烈��tɀnd�w�(@��`/��ڽ�T�� -�\��R�E�01y��3m�B��^y*S3�c+l�*e�Aiց7U�X*�`0��e��V�U���a��]b�z|I���t����e<1ŖE��K��Y;�0��ƛ-�[X��[q��;44�e�s,��R��z��6mrݽI`db��2��Z1����S�!�1В�[�.<�����e�*���
!m��-���*�[QmL���x 5tL�olԈ�:�?<�[Oo�5�<�sr��Ԗ� �97Q��r�$�3r�Y�@��FC���Ј�v�)��l5�$����յc>���tRind����0�e�#��`jL� ��j���J��&�YJ���$m�aKA4�Q5k��IS��u��ֆ0�_pa��"����~)��-�&�� -���M͹{���b4C��Jv2��D��Ssj:o@o���M�Yz+J���e�J�S2G��jK��N�ŪŤ"X���쥖}�eҁ��c�b�ə2�Y2�O(�����°�X��ې�s Â�j�R���9+ ��` ��4f��'i��վf3��?*Gd���1h���J�� �_5|�`�hU�tF���yuTR��N���:���nTU�½'#5�N��[��NؤGV=�KM��Ϊ��wP�I��x�!�	w%̢wpڂ�A����c[�Zz�H��Q�������n���F��VI�7I�c^X�J9��ּ�El�F��]&��x�k�2JB��4����mOE�;feh+R�6 Vj�Pݩ���F��t��� [�sV��Y���,� U{BQ�x���Y;�l��YCVͻ �\�g�ܫm�����t�AM�ݠni&)T#�rdZ��ne��d��M
� 4�]�G$C�%�F�|����R4Rg����.nS�0�Wjd��&�b����% [�k׻�YP�qn!��GG��`a���&��v-G��n�E��m���T�WZ��6͂������)����D��r�,�on��`Uꎤ�7��:YQ�F�'T��-�D�B
	��b�VS�#hj5~��em̹YAK�5���l�`��¤��ǃ-��)䣢N�5��1SXV�N�r�Qmr��nU�"ՑpJ����ٵoh�Z��x��dR�D�ܳ�-_���6�o�(n��z\n˫���x��J��m��^��l��Ne�l四�1�
K��cZ�jC�Ҙ=�+p�2�/Fcj��٣t��J]�4�s(� ����pmdJ���Q�E�|�����7i갨mI0L Vdٷ��j�H��z�A{Z�iD�3j�u5���V<rf\�z�G�������Ԑ�N���rSЖ4q�Z�\��M�Q���fV�zġ��j�spm��R��f�xI֩��H�rҺo�ѯ�(���xݼh'�.U��Z�#oD�0�)�����i7û�v��%cs@��[Cmh�aRw��̫�l��T�C����o.,�1�{��uoyn-�*G�j��V6]Ȃ���9yx����ص� � �u�&����t�r��Z��nb!�Օ^��:-ЉeQx.h(���VM�Enci��ej�:vI[����c�S9a[�r��%=@ȰB�����HZn��X7L�QD`�L��À�XRW��:b�M�r�Ր(�����yg&��=��n����H�X%ơ@˒�H$�_Y�[��Xsr���<\(�Y�9�����S#B-��D�km�1�H`b,+��aa,��⪍&�q̚�t(��7Ux�\,��,0�E�m]3=uIn��ڸ�%T)YA[+��d��$�5n�j���xk
�� ��]8C#�-�6�$�i���eq��黮�0\���HHE�rEgL}�,�!��Xl�˾�aI�8Y\��1�VE�W�\����@&�:nhwg��b���[�G_3ŝEl1%qgK���$�yE��Ml��-�����X�8�]�5��SF�bm�1�l�p@ �@�I�$��Vd�uRCRF*J�@p�K7�v�ɹT[Ƕ��a��IZ�sE<���54f ְ8_D`` �E���a�D ���TqJe�Z�b΋F�"k�\��]u	B�5v#/��1pp0Dpd㷴0�1r%Y�&Z��r�ZA"�ʻ``0!�Ț�Y���g��|��G�?݄���7���ߥ�>��a�?G������U��R
7�z5rU �W�3r�.���[�C�������m��j	��DԲ��[n�뼵{b��q�D�sm��%��:غ��1Ǚ|>�!�n9����76����vЄ��E��ޫWZ(B��-���ܲ��"�Ӫ2v�2�C��v�_2�WAb�>J86ő���t�b�;�7�����F�'Sgkٹt�{!��JGS��3��n>�Wb�ۻ����x�C:�kw�]�T-#������j李l��K.�o���S���IEM!r�κ�`���a��%�.�t�<J݌�]'�TB�8��c�QL���ZG
[S��e�k4hv��`ۈ�_����5���.
Ὤ���if�*��uk�t����	9�#zo���ϝ�g��#��)�koG��f�2�۩�y%ڣ��..�rn>UxU��g�t����вp�w/�!��Q]}Mتӆ��ai�EǮ�P�4m|i��\a<\�v�Z9�����V�J;�&��L�hYG�!x��֓{�1m����t����`�t��<լ����On����; c�Yܡ�M@���;�i!��8��͗c{�z^-�A��)�}�^�F�l���8V���o�����9�<�n��	��FT��7��>��M�)�!�H�h��;��ZY⸘9��Pt��v��ui�Z�e�{�s:�V���W�����e��uzdR�ʻ5-�8,yIf������'.�W��Yȭ�P�U��UHT|��l��c�3��KJ����Y*���3�u��Gq�k�݂��Q��ǚ������������,�3��f����RK��8֖��c��N,��u�тm�3"v;Z�&_3�ju	7S��1y0�ҴI7��^�#�BI���Йt�+�rb\����e�#�Kk8i�7LJ�7�Zw�����Bܭ�[>�u1��/^�J������T�7��k�!�Z�O�:��|!]f���]�vdq������'ϋ��fe˕:��)���F�;�Ԋ �y�/ce�l�u0��T�|q�P��ܾ�tn�9�� �2;��D�-Q"��fت���6q؎ف�'$��f�t� 8_[�qf��j;�s���z��f��Ɏ����$-�{�v�ۄ���"�3��G@h�',�����ř��DSM�y}�b���P1����A�VK,���!�&�R�Ǧū暭N�mX�4qe˪�bF1Rc""�Pu�0C��ٹ�ln���-GD�>��oyf�=�p�*��im��+E�٭�ӳ���㛝�y��Ѡ�m11�Ʃ�f��;mM��|�¹�z�����F6;7`���_P����}9*�bm������ɻ���g8hE]cEkɌ�q��%f�y���p�$���WP�d}J��)L�\deuq�M�[A�v����ҍ]�U�17a�q3k1I�鶶���s�x�	z��}�S
�B$]��z0���ǈhR�R�g9���s���*���_d�.�l��Bݼv�Ŧ�6x���]��� J���-��q�oN6��yC2�V�IR�ܙ> ���,ǘ�N�8*�$���yLN�� Km��TB662�U\1�@�)n_$4&K��cNd���8�����q&c�Թ�o+Z�Y[CM6�y����B���9�B�n���1m=��u.�[��:P�.�ˠX��oe
���wѤM����;����hnMѦ���DE���-ݳ�ѫ�KK1\��;�.t3���l�Gw}��^���o�����[٢3�fnr�^��a�Ᏹ&a�<���痪8����n-O�]��I�z�b���zi�e��W*h�3Ô��׵{��$�sy�Ց��\%�A�j��FcӸ����Y[}n[4�=n��w�c��2�'Ve�t-V"m��L���[�~���S�V�RA��%�3�N���Dn�ү ʽ�8�,^=-�h�N�U2�Ćܕ)�ٴ���mM�Ɍ0:�깣�O��Uފ��X���"��q�5�mW�S詍J��9��\Q���nm>���Շ�,Δ2��s�5�1�ځX��uC�^hX\e�V.m��܇��)�2���IN��!�#[n%�q^X���zsީ�q��:!�e����Q�Ju��R�K��kZe�HU�dR�����an�]%���6�g�����4����^]��eA4�*w֝_r;�q��!�D\+o_^�Z��r��l�ȇ�i���O��$&�y;U��l1n��Y��+R(.V�m�C\޸�d�T��})<�5X�͉M�fC�m
ϊ�`�]-(պ.����4v�D߆���V��U���{���mZQ�n�ש]a45-B�������M�L�X�1�YC�������*�BawXS$GGzx�^�Zk;�?4u9���=�Lκ�vt�"��%�Y�x����PV�"	���b0m���M�Q/���h�WB[���7�mټ���-I�;-ݽ����zV�bb�OI�8�m�ͭ���Q�\�&�*03$�&	�}�Nf�.�xp��lD/����J�>�g3��)Jx�N��|�h�X�J�[�8lJ�M��Rq���t�^�z���u$RM�����uoNVcF4�|mmD�]����Cb��rn,<r�s����%�_�k.�6����;���H���-��;��E,����cP�Z����U˩�d!V^��+)s�1ݾ���k)��� &�Ⱥ�[��2���
,m�<�8s��q̎�^\Sޥ�M�1��mr��6�Sʮ�.�wY4��=�΢����3��wy:�I�f�����fL��Sb�U3!�r��;�s����-d2S�l'\�Y]/v9[��H�	��3�n����iRn�`I�
t���9�ק��.N\!�Ӧ��F��UQ�U>�y4cWl�s���
Ȍ�ʔթ�B�	o`K����t�%�	!Vj��۴Œ�_	}ʹ�vr�N���=P�օ9w��S�\GH�tP�]
�
y���F��Vh`�\�'�5��n�vǗ��3l3Nr�ӳD�0�|p�]S%tf�r,�V�W�4r������'�[��I�e$M�YZ)2�������0>�Qƛ}gpӏoq(�3���[/t^��.�.6e��J���ؚ��-�UYkw�m���<���B��ɋA��e�Ŧ�^�w�S�A��Z��=z����j�8�ݽ�=��k���v`�!���e���û\.QַX�cE5��R��P�o��1�/$❭����Dq=�[{������6eN�\�x�og;/n�3����fc�	k�r�Ѿ�Զ�(�cG��� N.[�1K�ʨ�{+��K��q�
(x)���m%4L��罌Kx�gP�٣՟|��p4n(���wbU��fa�-K�tZ�M�/w<�$;���}~̄�+&��/��{���t	j�c=Wɉ����2�j�W�R���xã|��:��K��8��V�����&���jP���|�C�9V�wf-��xn�R���q.���m�t�"42�����r���gv�C�n���K�2��4���q���9ޖ8�m،�zt��z0v�Zcn7.n�f'��"�ܧ3u�dm^��Y�5����7�M��v���m�[p��5� �"ˠ��t�[�k���(�#��Ӛ'���+nX���	��q:��$��fHGR.�:����O	Rf�ɴ����Y��«	��h$-����`8#�+m9y�`�yt�-����]�'f�Ct+2�/�{wx��Քow�{��w�J�W-ȱfB�'KKM�u���{�e�R�������BC��3�)hE��["���,ιI�<׫�Z<6*����$�җ`�kvfsV�9D1Ѱcɝ[:����l�	����s�0�]��u_*�d�K&�F�l�clh\�9Nnl�[��s3Q��L�I��	D�"�L�S�@�S?v��K����a�3bu���s�c7+S�8����nk�ˬ�*�Q�'\����_�8��)��lb��3"ǁL��f]��y2k��5m�t�Pw��%�J��e�(Yف]�q�d�D�Ay��yԌڅ�z��*f���Xz���̬���x\C"���%�VkV!vr�E���m����Z�\�cޗE��3h�Ŕ/�e%5usMh]y��4G�ׄ�ˢ�j�ݒ[���Q��:�}�ޕT���Z�G�0��"��p�`�H��\� �H��j��Z�00RgZ��Y��ye�G_v�8���j[�R�]>�G������K�U�N��*�|x�"��e�,,)�y��pU��Ÿ��#Ow�Y�g����ń��W*=�l�x+b{*dv�В���D6#hq�;E��.KE:ಳ�ވ��:�|�7�����ƺ|�^�VQ�WyK'��ք�9C�C�Ko�������4�����vL|�^�c�s�7U�����*A�N餁.7�b�Gֺ�v\W�h��Qep�:�2��:��A����ǋ	���I�ui����s7s�%eɏ;��6T�lzyC,nLs��y��_(]�wEO�SXV��B�M�Y�{�"�=������c�����Z�\4�mJ�FX�Z���N���ԡyz{c��{�.����Tu��g{O"�x�љ�t����":�b���zNL7k��l"�[u���������u�5����~���o�<M��R�����v����I2����ڛ
�zo�]�!��&�ؑ�奘v�?Y����(p{(�6����tg驊���k�.(9���TG}o3��&��(QڧtLu5r9�3���	jrv�P*��*�Ժ�X���0�-�j�Uר�tlu{��
��D�FRa�Hx�С��J��Z*	������L6�����t��@mt�܅΅.oc������&ج|��XE�BOv�L,&�m������kNз��s�R��r�d���X��H�}2��967OJ��6�_.7��w�qyQ��!���w~�Y�}�7�n���uE�����66�2]�z�a*ќ�a���ųo�S����@v4��qk���۽x�*�-7Uk�e�
✮����yen�C�F1tT�a��s��|�Iƕ����'Cϖd�b!�ͻ"�5v�ê�Wq�(&�,����-�S{kD.;�[�".��g\K�v������LJ����@��(����We���y�HvG��H�����^W=��6��2�"E�uz�]����:t���vgv��e�t\hr78���:��ul��P�l8��ʬ�3u�S}9�m,�m��a�^��5%�$�Wu���Ȅ׻���[���Q[��S����u�f�V�;:�Qf�riF�0�n%�f��i�`�{������<cC$�bW)W�G�,I����ʩ�MRiթmN�۷KAUՌ�6X�:�(�	к�N���������|j,$P}�M.�;�����v=��w!rPc��37U�#[���t��[ˑ&�l���ir����vD��&�ۊ⽃����[Ҡ��,*��/�y��.�z��,�wDz�m��U��R%��˭K�T��Ž�E��a	� �`�եj=�%�*�dv��S������[.���0�d�캧B��ؗ$����Yy��]�ntKIbK����4u��L�d�|c�6e���AN�;�N����l��a�{/.ft[6����i6%)em���_v��X����k]d̽��3��D�tA(�N�۔ �ĸF�}�q
�!���z}�cΩ0{���{��ƞ� ���ZE�P=Y��py�C���+]ll��V(v��*�v����տ���J9q���m=��*TΗ,�黫#����NY\Y�j�Ft�Y�yU�ٝ����ihF��/4�;;{sL�(�^䳙��X,0/ ���N�Tjc����ٽw��k�)E�O2LWb�$�H̼g]]g-�.��v��b���:���2�u�p�C�&w:�6�U�\��x��>9�]��c�c����a�#�Hd�ӱ$���Ž����%,�r����a�8j��v�&UЃi��v�C���H����|}���Rǯo��{i�㝯M	ՔT�}I��:Xl�7\-�S;�]�z�ۨ�S�2�c\�$W�7T��dٸ�E�<81�)ӱp��]��t�u����9	�
�����6��+5E�d̩�ck+���#�k(���Sk�ڻ}���y���jJ�����{��+p�y��a�z�5v��{���A�Y���Sq���%���7������4��0�1#6��ҥ�k�0c����h���p�W+7��\�8��	�f�b@�8Ԏ81�ڢ�K�Oi}'�uA�N*vlAi��t�d�*�b�QB�:�)�W���؛W��ޙu��Δ��'�8��e9������I���7�-+�Z}8��*]'�w�9)�;
x=�|��8O8q�|F�Ϟz�'��7�׋�^c������['/��"P=��|����: ���/�4�=�@kǜ�����P����7�O0> /^|s�=����֗W�/˛�ߝ㇞C�����܆�>z���|��T������7 �R�����p:I����D����?O
����}�߳���)���?��p~@(�/�����<}�<	^�^/73��;�\�O"��޻E[*�%�Y�D��T���%����l�6x��`˝)�$t��*���r�qQ�)����M��[�n�AT�r��I.���D�9xuP�GiuM*BNJߕM\�,��~�k��Ŝ9��H�;/O�#����UԼ�sj%�uViL�~S���3�>��V,A�|e�;�d�'O-�y`y7V�BS� Z�����"���*��.�a=-`7��D�Y�1�^�'�-A=��7&���٦�p��3U�m�]�@��3��3S����y��n���݅a��`��J�zY&d3e4e�w�q��,��B6��%h���ə{�;���fZ}ED�D� S�ՈVvGN�=�U_�+S2ַ:��N�������
�e#���j�f-�H�;�5i�Yq��RF1�ͶP�y1��t^#�Y-�m��v1b̘��T�2�h�lw.ڕ�Z��]�yh�@�ݦWp���%,w0_q�:���V�+2�h{Z\ʒ���ҙ�E�x`yΪ�LN�gI���S��뛇-hU+d����]K�3�3�l�Y���,j�'O&�]�;2��w_t�q��q-[�nհ���b98��ϖ�8҉�V�N���Y�k۵�����f���JS��V�[G�f��Jx���^~�w�����x����w���z���z��ׯ_�G�^�z��ׯ^�^�z��ׯ��\��ׯ^�z�}�z�_/^�z���}��o������ׯ^=z��ׯ_O^�x��ׯ^�}=z��ׯ^�|=z����׬��ׯ^�z�z=z��ׯ^�z�z�z��ׯ^�z=z��ׯ^�~=g�^�z����׮z����>��):��1K�t��x�n����UAn�8��7T2��*�{�t�]�%@G�J.�o�mms�YBՇ����f�z�ob��G�� &��E�~��yC#�o�*Œ��gn7
x�;WD���7�;��:�x���+�ȓ��=��]�u�.X��CJ!%.�ξJ��Ǽ�w3z��
�GhM;�9N�=miaܮ���XIÒ��D�_f���u����N�x:�����@�t'�[`M�Gq.�ºA�Vd�j��0޷vٹ�f�ˬy&8����z^����\���C�{�v2�{V����)�*��[�%۵9h�J��LM�S~�xY]y��ʋ�rT����/g@����]���̈́s.��i�岦p���T�
���J��m��s��tN��o�h:$�=ئ؋}�A�%��͗/uU.���o(ݷU]æiۆ`���Ǐ[���zyY��b"�[��jG���}�^6�՜�z�!�z�������ͦQ�K{�Ӕx�K�ZN�C`����SkJ��Ѥ�sg�.SM�y���ulv��D���H���ev�8Jm�;8�����J!Vl���lI+���.��T�yݍ�,=� ��Y��̭�����p���m�E�,4a�b�a�"{NK����h%7�T�v�u�7y����<����9��|����cׯ_/^�z�}�z�^�z����ׯ�z����ׯ^��z��ׯ^�z�z�랽z��ׯ��^��ׯ^�~?o�}��o��^�~=z��^�z������ׯ^�z��ףׯ^�z�����z��ׯ_/^�z�z��ׯ��^�z�z��ׯ_/^�z�z��ׯ��^�z�z�랽z��ׯ��Y��ǿ�=w篝�%����f;��W,Z"c�]�y ���O*�n�̇+�j���5��ugD����&�4�_�Y��a���-Zp�u².��{����
}���'+&C�Mhy�{wn�Z���0�^n�t<)^��Fڱ��FM�EGB�e�}C*�-�k��͘�������Z�X)�G���F�����z��0�o���a%� 2�k�O��:L�䜩k�ƶ�:I;��u�v�6��U�� j�Vhr92 n��V�y'h�����aa�}���e�6�n��!���a�<�4�ܩ�8����u+s��h�`�6��u�°�=rj|�ت�R���'mu1S��%���ٹ�cb���&]嬭$��1�5sћ�^�Ж����s�Y$�ʫ����s܁hѮ��Lh`S�r�I��'}:����3�ֲa�l��]�+k�맙&�'+S��7i^ *h1�Zmh{z�`F�!��$�T�IӔ�AB^�k2n��b6V-�*yz�ؓ���`����دV�%�N�F�1�ӟr�Z	�*}��,n�h�Lb�����j�5ƞ��4��K�¹FH�-�ڠ-�\]��בVA^��rl��N
����hd7|V�vޚO\����I,��ko��WU�-�g0*�oB^΢��ܛ�Z�(��=��ў]yIྫྷW�g	ʧs[��Iً3;q�.|�I{Od�H��T!ܧ�En^Mڕ�-���,Y���9IV���',n�W�{0��8E}0'vA�X�0^"6�Y؎̹���^jڲ/�)	cJ6D�F���4^�Z�X�%��\���`�s�[�P��[/79	M�2��m)\������I�E.$M�ڍ�����a��!���lo���3�B�s4�t�'�6v[]ʆ�zaU�~Rx�ˮB�����A�t܀����y��'�V[GjfXGm!YHf�;B��O\�TU�h��.�Mw$�C�곸NYC��k�W��EW�U���/0^q��ە0v��}s�^�JVu��P<ۑi��E׊��rl�#s�V�Pė�*�[�z�.�m ��7���'Pb�r��)xE��R�l33}Ӯ�]�,���׻��ez��SZp��l�K &�]d�ھ�$���B�2�[P�'+!(��z�l�{x�_Y�K��e��:�F�ek�wf�Zxؠ�*A�]0���[�z����f�rw�(�f��狵��N�ڻD���Ew��v��ڜө7���K�s�����"�한
�#m��s������S���e���z�R%:6�+*v�k9�<�H�!Ot�\I�B��L�Z(jY�cA&:-���|$��)]�m	]4�J�m��;��3��(�I��沇]C�]��D�������pFN�f(/9��ʄ����%Ԯ���<rpU�8:ҋ�gJ}_�k��ؕ���	
3���Y�f�7�~��d�ǇV��JB���l����9��/=��f;���� ��Z��v\����J*���������J�sԮ�<��.���Τ{0M.����np�S9�n��5t���mW�-ґ[�V^[���x�cH4H�ֳ���!���*/Q{fm�n57[�^������u�������1e��1[�O��sqv�`���Z�b�� ��`o�}�fw��KV̎���P�XU�;ZՂ����P��NBNZ8�hY�y]�8�ܬ��N�멋J�n�z���4�-�*޷�|L��+N��M9�H�H��qV��%]��o�3���d����V���N��U�-��'�r#�h.ں��f[�������ˎiޣt%Y�
��s;/��xj����y�d964E]�vh�(�[��͹d1sZ�F�w�Ǳu*Ƃ �.�'m��v�ǹp8G}��̤z��r>�o�ۂ��nn�j��a�Ǯ�t�x���5y��/a����vJ&h蚆<�=��IY �n��_,�f�%�JȮ������
���Cǈ*v2[B�?�C%Ž��r��c#����P�+�ۼה�+J_3��t�a[#F,��0e>����p�F�uK��j"����s=|Y��o�b�{H�={ʪNqYa�7�f ��M΂��ʬ=lq�+w�z�.aoHo�kN���u�����%rw0�{𫙕�s��u�\��xH,����5��ǂ�l��7���s�iҳR�ҹt\��eF4��)J/�l#�^�Nh�޴�	z�ab�)�N;WWWU�j��TSt�b�}Oo��o$��&
����īR�2<҉8o�n��3��$��KP�kpd*E��Ԟ���`��h^���o@og'�a��shŵe�[�	�.��o:�*R'�[2V�c�v1pY��Vqf�ZD2��\���hv�|���.TR�ӈ+�A����ث�3���{zC����㒶Ʃ���z)7^�����!"0L�{pV��w>=F��迚5�J��+j�6^k�f�&w�7rܺ���m�@�-��h�DwfZҮ�mޡX3�ϗV���d�=�Y�u~�uЙy4�.��{'�)�6�m�o�۵���OI�z����`�`� �ګ�Ȓ�P����׋�[b����;f�μ�9�
�d�2M��C��l��t*�r8��F�$b�t���wR��[;+�j���-�fVb2ݣ)��M9��G+�o�;�Vez3�)ӗ��z��oW\�ї(��<�3J�~�4Wc��c���Vn64���}���Ҁ�};y�akx�(I�1IB��ՂF�T �rݘ�nnӬ�{-j|��w�Q�qB7@҇{nN� 9��o�Ou�C%�V�M�d�0 x�UT�oE3�� ���7����H�[:|�����4f�U�U]���3���=�yQ^*�6U�)�'b;���*��j�LU)�Ta�*]=�״�ӕ{�Ai,�3eh�U�>E"�j{_%�/�"ӗ(�v�S���%_k}{����HA$�GGN��14y]��ʋx�=�\�t#O?Z4�k��Ζi��؟YC�y�EK�}ݶ��쬌�4�8����V��-�	[�K�7��w��w�K�����V�C��,
�zH��U7u�B�kz%���uP3���`����`P��
i��y�Q�o�O�x�}S�oL*��wv{���bڳ-��Wg̑J�7yu�R�}P��e�=jTI�E��6�)��ʖ��;G%�{�GRT�Ӎ����i�N�-��6ھ'2�,s�&�:˳�P�p��z�b����H�ޝ��uu<�saz��ďN\d���:����[�ܳ��dcX38lv.��uJ����)Tu��[8�(���u���;�ݩw�*k��:��"�]�A�S�ktr��i�r�9�VȘg'a9@;.��VK���|=*�.h�'-p���-�56]�d�T�
*�	o�rN|*��ئ��'�TKs)eYY�va��2Ă̻f�m
��mp�N1�^օZ�kkm�˕u#�f�t�Ζ�S{�WI@P�<x���V^��V�������ŧawK��n���o.�[��`���\�Ƀ	_m
z�y�1~j���|�==���9�=pru�Lhq�!e>�#˸����"r�kcz[ެ��6��Q��9����3G��d�h�4�ϻ
]�b�w�Jp=�oShPUֆ����pn�sV-�A��Ķp�|H���c�n��X���������RGJ���ё�|p�|1��\�J�^��66p5�E��E�1ZCa�9t���\��۾���!�^�Y8<\�Hl���nf�SQ«մt�y�C ʪ�r��*�:�a� ���۱�����?CG/���ޤ���}��Pwʹ�E�].\B#���;k��p��*�^7S�cğ�+���r��l��S����1�5�dr�s��:�U�v.�UjZ=2���>\D34�$�[4��تx��&j.��Z����;����1�r�[F7us�{ � �#^��l�8lK�M��I�3(��
�o`�;tm�$44R�a7uء��!	�Ƶ_]�[����x��n�P�ת�r�����^!���f�'lr�kvv�t��)��ٟVe[t[�"_k�/r�� �g�����f��!	#8������E�K���ls�F���A�LN�r��^��6��;�fξ���Kn� Ne�8e�ئަ�l�Ժ��e����v \���JY\Zl�l�9[���,ê���m=�r'Dvk)���������{L�vh�|�:s4Է̲rm�Ū��eݙT:�]J��"Cg��4ia���Ba+*���z;k6S�\�4���-'���ԝwU�m�;��b�SN����S���?k[��΄��a9Ⳕ�B��}�t��o J�%�8@7r��ₔ��g��b�͸�gh��/*Rx_L��Q�z�A��7�=��1��%���Ӊ j��c46,7���λ]֠0]�q@!�޹[
R�a��v�� �:mbkM݂�1�ݱ�uf�Q�����*�ً��tb!�\ђ�"�|��g4�-�G�t���Y�����X1Z��	U"u��EOa���B��R�;ܮ�V^FEJv霸�Tn�+�Z����(iU�K4oA�r�ȹj�^͕I5�۴�_��z��퍙ۜЅ��E�e�4�WG5\��3+��ݒf;a@��xa�U��	�6E�Gɋ<�<Ǌv�}m�۰�=n48];¶5	�,_O*m���0��1o���85����dv��&n�e2�̱e�b����ejT���J�/xڣ5�M[#ޢ3�����b�ۼT&�Q9}8��NZ��\��Q1�,u��&s�txJ��+i�!8#�t�+��P�M�M��иF�f��}"���*.�ۺڼ�(�%�z���tQ�+-x����
$jb�U�a#z��tQ��o[G8�tV�s]�;�T���	��I�ٰU WK0�����w�]/7��z����V.`��,���F:f��s�:N��k)�J�9�T{u{�-����FX���kp����p��K㭰g*�e��c��O]����qr����Y����4�\W�t���R��Ў�:
����{�D�,U�3�J��%�qij�Ɉ��]>��)M��%�X{*k�R��y�[|	�z�*��[�3b��e�U.]k��W|�+��������폤��C.���o9�KE�#M��u.�������q��@����vr,m�+{��wq<��X��2$A��0�s?6��ʍ�B7׹���mͫ̆�-�q��� ��=��I�
�9J�4���[f ܙF��8�43+�`��⥷]��l�k�;S��zNaG���J^��/�^���S��Gf�s������y����׿����G横��t��������Z�������o��O��S�"D�q&S4R0��2(�R&�f"E�(�p&�%����)W�)#H�����R&��������83������x*-�� U�)��~�P4<DP)���Z�
:��L��h?�FL4(�E}]��7/�wL�]��8?�	���"NT3�F]u��d�	���h����ۤ%u.oXN��,��b4cYXV�;�hp���* �_Zg�Dv�Wg�mvcp"�qМr���]�����&a��j�;�)�m�+��,��z�o`��S_L��5\z��J�ft�cG1�	�$��췜��
��qw*�J�x�lLq�Wz��f�r5ڞ�5ǵ�g�=��(��뺐�p%'s���`�!�%��*�f�36trT���}���+���8�gYƏJ�ʁ�Z%`���H�:�(7��\C���L.��]�+A�3:ROye+��q�;ϲ��9�g���]��������:�.V��O������Jٹ (�ÝU-��Z\��м=0����|��V��Ю�x�d��|�x���!�K�L�ОWn�z�;In��b��3#tQM�R®�Q<�vm>�Cn��{]/M��z���.�Itb��4+��㮒�� %*�x�K4��cC,�<VU5�s��%vs\�Yw�Nt�����Aw����+�ի�)*X�
̏h���>����˻�q���x�h��q�i����i�_�eߔ�C��9�|�c�Yq�V.��G�Hnѵ��gK�n�Y�s�#-�H7=�	��[q6T�ԭ�:�4L2k��Ph� 0�?���	Z�%�������ؠT�t��H�@�G��"�*@ƐR~!D`xT�P��Q��dA@L%�QX�"H�p�q��7
M��P��A@Rm2�q7$-��&h/�6�P b8YG�"E$Ro�4
NF ̐��� �i8�K�j��ƕ�]-��(�ց������.D����Q�Ć)mH!9!~�)�,Qi%!�D(�#-?�#!08K1fJ���Ggњ��Z.m<�����ͲUld���m��F6vqm1&x�|��������}��o^���{��5�v�N�V�ƶ�mf����j6�m�*����lV`�����^�z�}��o��������]�5����1��(�6�E�54r:^9��ƱZm�ڪ�V-	���1��\δ�Z�S�Z���q�VKF��0cZ��1�cg��G4�,F����l���Q�i��TDU�mZ��p�N�"�֬mFب1�X�h�&�� �Q�jѢ-cUE��;F6�4UTM[�9͒ѱ�*6���XųQj�,lF6�cK�U�bڭjڢż\�X�mPkmg��ccZ����i�!�	��$�M�h���L�֍�׀�xG��s�1��ss[mfx�5�n[q9��sp�y�QSUdѱ$�+�=��x,^<��c��并��<�^����˅`,T�[�1[:֩����ږMx�j1�xp.q�s�p�A5msOG8�9�6c��r�r͹�D��F��s����F�A�o�Vg\�96�b4ch� �s��F���ڣ�-�tDm3����έ�Ѷѧ�(�u��S�X�\SƊ׍���؝kbH��9�s[�#\Φ��.[kFk�,s�S����G���p��D!�ơ�DM2W���Ϛ�6�ٜ��K�3��{����G&�.�W��K%`��dz�3���^$�:����wkU�����iHBEDL�KD!'�6�a�����1FQ��b��L�0�~?��3�������n�� J�$و�m�ڳ��7�#�w}���u�퍼3�(����w�Աs&��|�x���N�ߖ[��Z==>��{�g��r������6%�]��VƲ��N�p-�?:�!6�V��+xQ��#���hq$�o4���N ��<����/��f�\��=b�<�'�=6	7����ח�L8�s4�F�2'�+�襏+t�F�g�y������\����Tg��7��s3ɹ=�y����<� �	�p��y~m�go.]�3����2zuK�<P�ߢ��}�z'���o�]��t�^q�J�����|�=~�c!1���O);S��ۼ�	����Ѓ�E�0��佾^�"�8������疽��d���zM��ss���ܭ�sPo=�J��A.��Qxg�1P��$��C�ǝ6h/ރ��?_y�<w��#�6��uyb��Ht�����:�v�{*Ⱦ�K.�������[��|U�r�����'����z:>=�w�V���V3�a&{�k���fV�]�
���/gvk��+�ɲ,�ו4GC���2e<��Mȍ��μ�Qh�E{��yƞ{�=�%Z����+���z=�]Y/F��D�;��0�����σ��D2c�Q��P�`�Ý�J�T���~��4=�^�f��>� z�AI���G
���#ƨm_�
~ӄ�u��瘇���~�__l���]������w"�]z���^U�n�C�����;[�A��8.�_ǻ=���}���$�|GH7]<{o(�f�v'���^c���w�>�T4�z����42��/�Ps����{���Z�Ӛ�6G[!�B�˫�T��[_��X���s�z���}�k�J^e�޶�w�����G�{X����;F��TT~����5�������k-�ls����a,�Ɵq�~���߶��"my�MØ�/���c�s��4q�H������y�� kɛ 7C��mf�5�á����5_[T�v�j���D��n&0��]��!R|��`�v�3+9SNi��
����Hp[�܊���H�H�=��wem�n����(Q�4C�X����:�o�h�B���c6ܖ�:4��ߞv�7C�&�\����y�̩��8��4 �)�LX��è	c|�����v��X����ْ�O���pz��{�R��/
V`v	�)��������͉O=�W��5����^
��@���,[�v����-��o�e>]���UoN��<Ʈ������/�mk����BU���j��e�����c�b���o�=��R9+��ǷŁ}�E/�>? ��P�C�Ay4��mmu������47�~�d�\�lr�F6d�E�A�=~��~��iv0���{o��r��|��-��Ϥ�!=�/Ӝ\�\a��z��8�Mk1��cLx���{�7�ȍ�w�����{�ថэ�{<����O.K�<1�$V��.]?_�#(5U�S���8H��5��E3��\K�S�D�%X9l��^�Qu��W�\�(��Q��Ͼ�S��e���	ȴ��w���\xNm�3u���[B��yJW.A]����R�%U�����G[:��{�ͮ�?uV^VҷR>���M�hCj��ц�[��n�`�Z�V.�� ����j�.�_�:�Ot|�4)�ɮ���=o��g�V���P��J�7�t8�h�y��Vܪn	K3JN�E�g���g�zzOm^����^B�0�lP��UpE�fk�v�`�,V���O3����mx{'��wϴ����33�1ꗝ�F��:)��2��vI7�x�ד#��>@9-�'Q��Q�Nfe�;������c���`|5߳��ֻ����=W��Ձe�g�O�^Q=��q�ǟS�
@����ߞs&���9rE�m���N�oʞ��)���둿D�Lf�"���ڂ����p���ް�J*]�k����xL����*n��j�n�{@���v('�4�e��Q@�l�����x�ϡ~[=&��v�h�a�w�x{y>���u��ث�����(K��"wj�?zh�<�~��r�j��Pt��T�6����9}�̧sC�x1����f�6zZ�p���t�Ug�fl�vK7]>P�%$Ԇ��a#'vY� 
�7�,�VY�so��V��'^ŕ�7%M���<�݆[��W2��:�#c9Ňf�͉ũ#��մd�BZ���i&�{�nb�;C�=��)5kT��e@C��X�Ӵ0�ˤ:�Ek�~����S��Pɻ���d��꯾��~T���M0u<gÔ�|����{�^]k�^�bR>��2�{{��ӷ��X��|�bC�Cҗ�K�+�{�|hI�̧����ߤ'"�U�9;ѱ�5b��M�{�z�K8}�}��ã��h{�}k*��.~�_zG�N�P����v��2n���kNmED��,������}f��������{E���c��VLl�~(�����3�Z#�3<Zʿwj���-���=��l�\�$V�ӳ�A<�{�s���f�&��K���O��c��(ۿ��ݸ������
�E��V��c6	1��j(���<���݊�?}�&���n�`H�8[���|6�/65�-�oڭIۙrO6�Û��	�=Z@��������0PF�����|��LB��'˵�[��4&�}�+���1D�t�Z��KLr�̆c���Ӆ��CTwF��4���Ze�i�|{��Eo2�XU��YۚMcޤ�*�b�P��;��ʮ릏�ꚬ�8_W�l�{�Go�]��)9t�>�k�E��Q���M���:�����7���&�=�e����i����$�cݟ]�e�L�u@w�wz+�wd��K�xAl��~C<�y�t< �t=�OE�{>�7�d������{�m���I=��>j� dy���0"���� �q�oh�~�߫�8���=�ԝ*��A.ؚ�����EK�� 1(�=�6��,E�]��	ĝ���$���6�w�Z����`��m�}.���k���Ѩ�!��6W+3;�����o[���=0l�,I�6����ϰC�������1�aߊbg�7��M���Wׁ�y��������� Ni:7>�:�K�9y�CO����ǿ��;���xL맏c05ƺ��$kY��m�d팘㹥���h���Ͻ��+<����͡ɸ*�����N۱�G����=Br3�J�~ټ����3���
���N�)�R���o)��.��AN^�;;-�F��u�~4����n����7U���֠��a�G��p]eMi�-����(i�*�l��Ȧ��.�q�R����m�iui��>�.ݮuR4���%��f�`ޢ<=�8^��A�C��Ս1u�j
�t�):2s�{�����wY����>�(m��e[H̲�\��uE�/#��mQ���m��8z�KA'�<p����l�ƺs:�q��ӷ�0�gq�tN�9-6 ��u���m���_���9��qc�WR��og����E{�^���^�6`\5O���걳����?w����z�;F��ٹ������}S���Y�vO�O |���DG��ɫ��=��n�K|�T�Oy�O	t]P'�t<�k�-����P�Pqv��R泷�����n.���~���V�����B�!t��=�3+tu�������<���J�k��Ƿǂ�x)��Aу�ۮ�S�w]6�swz�w���ޒ�3 �>�-�����Es5��`��o�+n��
�sX�N�1�=ՁQ��C��{'�������2�ݭ��{�֯g[�N}H]5���;5x6s⎌�0dYt�Ņp���ԭp=�m\��^]o��Z�x��	�����b;��%�M���C�]��HV��.on)ǲ;c�]�ԣ����g�g��]0r�`s�y��9RĐ؈l�����/�~~��~פ*��ۣ��^�����M���m�=�x��iJ�[�+q����Idm�f�
��ҽU����n����G%~^�1��h�����Ҝ���hg���`�}'�ڨ����}�����_wե�_�fl9W�0��%���#���z*����1Οޯ�tzN��H�;T9����j������9@��d��d�٭�s��%ȶVX[Αs�gVV�e�
�~�� f��E����$׹��q4k�x�y���E����}x�[�h��䱃�Ü�zph�2��vI7�v��`F7�yy_��g��~jx�;�"�f�k�`�*Ƽ��ExaA7����qۉ���\]�X��.�ݿxy�a��������w�䬷��������_[Ճ�.�|�6����v�2�#��m[�t����논�h����x�3c�Rv�{s1��u:�y{ �%��T�7�Y4��v���uw�wj�C#$�랉��H�3;yu[���K�,V���7��B�M�Y�M�&���Oo�J��m�pI����O�9�0A�14h�M�=�{��m� ���;>rǎGMn��7�ᒜjx_-�����OL�7/ؗ .w@7��@��P̀��0\כ��SY�����]j{�r����n�����S�uj���<�g�����/�Uv��c�z��7����T߬<�o�Xо(��딼�.e��X芫>��5��Q
Z�X����+���\���dnW����r0��k�}y�c��N�]�.����/|�s�sn]���a�7�� ���~�9��&�	������L��p�~"���7���C*����㙐*���5��d�"Op��~ا3���ٮ�y�����>�B�_xY���[s>;�o�<����ڏ
�~1g���t�w�N-�%�؆K'�<��Ֆ�s�8�M�6_�h맼�!�x<k�y]K�N�\ �Iׯ�[O0M�f�z�Nzw7�/�S*#��u:�xA�_��,՚C�W��4h�ų9��&d�-o;�܋�!�z��!۫a�Ʈ��gdfv[�1Ҽ���_e�%���]Ku�5��W�"�>�-��G�0S��f�?8�}�I�)���^� �k�=��`���U[eP������
�n�F�oo�#3��"Ɵ{Ì�Az���/���x�<�^|)Ә��<�㞞�X���>H� ������s�֑�s�[��Z:�d�z~ӳ�l����;��B��`�Z���7��{�S#w�ڹ���������="����#�Z3Ćs��I�����W��w=���:Nݓ����r�����Y�Q�"K�&��͖3�Z��D�Пy=}���A��H���3�7
��������<��|����_�z%9{^;�uR8���ٺx,s���;��;��*sĢ��Ӿ�si���E�6��#���9ەU�13�)�C&h1����;
w�`��
Cu��"��I�7\v�7Γ�L�ي�~�l��in N�\��՗���_*ꊙo6��������
f��P�h�5
c���a�ŷ�xY�����Vd�{ 涔��2�,0��[�؂�S٥�wAZ�1s�̥&�hu}�vD��t�=�����4.���)�7WQ=N�[lvt*N�}a���;9A�9mFG}/�o>_|7�јwO�vQ"n.B��b��|�=���,:88ᐢ�.�����C�X�;���ہar�W6E�{#���u�RCQ!:�Ì���ckN�7u�ǆR�*H��K�W�bfl�f��Q�X���s��wy��b�3Ftʅ�Q(K�P��ԑܺ$�)fP�sq���f@�.d�d_ua���+�=�p.ʹ����wtD7ͨ�ZC�×���#s��N&�v=���7\�=
��9u�bW[����#h������#\t囬,pR�ړ���s��MeK3#�c]%�����2>�k��Ӗ*\ �x8w&�3���I���IG�V^Hxc�u3�R�M��=��oٟu�2�J�L��╋ctE�OԸ�hF�v\��\KgIP�:��mm�Ci o�*��Xل�@�+z�����C�E�� ��.�W����DJ3��R9��Վ�콁&�����q�I�Rv+{7��!��'�s/Eٿe5��y`��/����*�
�L�֯vpqC.v�(bޡӲʶ��ztXEL���!ҭ"����@��<���b�j�|'��\4���\��4�0.�o�����T˽#6�i�4�S}r�VQ�����J�"�鋯9�f��ۺ� {q��ƫiGZk]h)d��ܔ�Щl�\L�?����w�v���8��4�03۹�n��N���,Z�m��:�Xu��J�7.������W=
vr\c�Q3G�WL
�)�j9������)�)ּ|�ӾG�C���
/0i��q�V呮� ɔ����1^��M)��V������9�yw��Lq��8^CuL���n�hI9M�6�t+3,�$?lV՞�l�4�o+YZR̠L��^Ү��U]��fl)��WtΧ��8���Нab�M�E*���E��\OJ=I���I� ��Zc	1�t6U�v��HgU�k���!=��+#�|E�x�̺����,-]�Q	d{s���V�\{k|�tQ(��;�\ݭh*�q��3.�Lyj�.�}Y��7�j#;C'�;͠foR.���]A{�p�v�jD���s���f���|H�1��hc��+wV3 �T2�-��"L6��[�xr+����ג(�)je=�M�M���b�v�����T�ǵ��l��<�Rpk�(�#�.���r_\6�̦�5���z^�ɪ���2޹G1��!ZF�w���� -�mSΙ5��j}��$�x~D����8����j�A��ny�8by�F���D��T@UA��8D�7������}�}��o�����~?_����lX�9�jy�DQ�%�Tj�
�N*�m�sb��9�O\り��Ï
����χ����~�������}�_����L}�qb(�(�H�(��"��1��i�Ϟ<#FH(�b��f�yf� 4j*��9��LܳAx���ES3��Æ�9W-DAA�4E�M[�Ry�EITG�h�TF�5>�������Zb�c�[Q���ɚ"���$�(����b&�QQ�H�`���bi��� �(�55DRLQM$�$DkTUTI����UDQh��#�DUE3��"�4C�QU�tQͪ�
=��S��{�S1O�̔j65QkE1�������"*"����J�h(���d�(��D0l��6�ATDDTEM	QPI,3E5U%bŭ@TSM�&*����7����^�x��^�z�㲖�/��;.ﳎf�F+L��݌�Q�݋\�t����]��+"qt�5�����t�(�s�o��}��b��[�$zvcq᩽������X�{��h�<���p��2n̟;� �uV�y�)9��׹��H���M�Y{nO^�^����oW�6nf��Xuy,��#&���m;8��M=\�n\�]����7�j��w��C�҂��5�3�"KO�t&@��oS��s��cH\�3�0�h,�`Y�Dݱ�W�]��=�!�d޽cո��)�08{wâ�o����Tc�j+Ӽa�6ɼ�'�-gc�U�Cٝ���[!����u��zi����;��e������.�!Cic0ut�b�h�e$xщd. �q\�Y�)W��XTi5؈�|j�hOT��v� ���.͛��D2Pa<w�!�n`P�^Pɔ�殈��>)͍R)�5�&�(�]o�0�?>5��"O�_�����+�-[:L�O=��C(�,�^���}},�
o����uI��Rr��E'�'��^���P⬌;1��6[�<�ã��4c�f��	���ٽ�`)=�R�q�t���JO!' ��ަ�˪��6I�����,���GS	��S�
���r9����o@��9V��E���?ew���)x��y��䛐^̫X�/`���\�6�g@��&gi,5+Nf<������N��0���ުm�A����V���9�7��q�1n�Ϻ��Lp��y>T�H]����MXHT�Fwj���f�W�/���kin:7��y�^k{�٘�G��c\:r \�?ybC��F���idA�ÿ�m�z�ȝu����ܖ�h]eh��C��U�W�]�sNh�`�m�\�V����Öi�V�׿_����A̎�3c�PW�-[�L:�Ʋǿr���OW<��� ��� �<W}�
��q�ko:^�H�C��}e�Qt�1}���%8%��o
�"3�o��1�[��o�����-�`�D?F6+��M!�gg^ ��LLt޹q��l�׾�"I3Eٽ@q�bĹ����O\�"�߾����_~�-=_�r&>2���=	:o\��S�U�P����7��9��
����;�bKz���i�خ��Xoˋ��l����O��* }岮}]c6����'9�qU쌷�����k��l������Fu��=�l� [ ��sӼX02FIݳ	a%'�ġ�c[à�w\#F��<j �6���t�p�7�,qtkY��=ǟ2"��Ʈ3�7��ɍ�R�Ok��kr���)xL:�Lk�d�.��A�=��o&KT�M⪓jT[w8�c4�TF��E+���A�y�wfLsv��z�coaq7/S����M�qSt�[�Ѹk�BRc��]�=��[����PR�*��d�:}C|��p$��oV�%6!�r'��9��Y֚cI7�����w�7�N���9�q��s���<��om�ьfy���DU,~��.���^���y��_����`vތ��p�jv��n��-�C�$��)�6
T�kV�)ţ4����[�%_vO�=Z��<0Cn=�hT����Pp�C �V�7�Θi�I�g	�lef�9�?��^�s��j���oP/�E��-� O��B5����`�|�ʸ˵kҫ�n��k�I�G��	yC�qu�ק���#N���3�`-� �g�!�i��yO�Z�n�{�v*dZ����b=F�T�q@wQaU�+�Z�B/<T�X�;Qq)��G�!���������%g��K�����y�KQu�yO�%��s�V��E�Z��3j�"y]�4+A=@�>�^���WS������e��C�l�cs  (,��R!�oUxZcrG���{�PK�m2�G0�4'[-�j��Ә����=��P��`�y��0Y�br��.̲oh�6�rR	�#5��i�+asȈ�4j�w{��=��}kdr��^� �L�y�O�y�Ƈ�����댟�_P͈�vOP�v=��j9n���#��ӯvC7cׇ��B���g܅x樓�y��g�~jS��**-���[R�.�lJ�"�w3���O3��&@� �<��Zס��ڊ,�$�'}�K�y�=�]gn㞨�]'�Pv�Xl���&����r9Eۦz�AF���VE�-�E�a����u��:���C�t��5v�Jgv���r�fɡ��	���������6u��Fz!��.+h��$:Nm��L���6�ƶ3�`0%��غ�^����j9!꩎�Bj-=��N4�VlY-C�  �%����� �c��>F��v+�������]�?��C��)�_���xUcan�&�w+���4��*D�Q�Czm�U�K�uTr�qʝC�O�X@�!��_�G����,?}�mT<@���%6�#!2+
N�ܛ�'*Y���j��h�[`�Su��wN�z1����v�
 ��'_!�C/��5�`7�
�&N�ݺ���d��z��W��0-JR~�(�h��p`ʅK�5�~�C�Ⱦ�b(�	ѽgSgZv�����ɔ����OȺ�C1��6��;��w��KN��̜?��#�H�83-fc^��!����bD��N��]0��=L���e��ۋ�1�:�a*;���|mQC�Ϧ/��wT��!�ً/G-�09��_*�c'qT*�zY���,qAo;k �w��yĭ+��cٽ�G�\>��=�5�0�Y�>�d��T�����[�)�E޽j;���r���A��^3_�E�T5Vt4���N�a��.b�r�Vr�ǥ�ū�b�����A�����KeɎ�zt�3.�ýP�丹�<eg;�?���g���FN	@es���u.6$2ƊWE;&��(�d�{W[=I[��q^�F�$�1;b;}:���������QM.���q��=8x�Dk!�:=k�z`	lU��,��&��ҵ��:�gw#�1�A}�ù�(�C�^y�������'ps�]C��xr
���a�]3�6�ج�M�g��]�%�e�};���oP�tx�6&��}J=�=�9���,Ƽb�;p�\Ń�����"����ͱ���<�/r2��X�k�=����Cy�^�O��=%��Z<;+�W��b�:� �g��9l�6N�u������cӸg���B'$��%�u��A�FmcxCH�_��8�'Ě�A���k������6Ի��6gSY�C��γD�MZ&�!�z�x�Zޑ��4�Z���d��ς��p�{#U�Wm�.um<Cm�Y��&�!:l�����O=z�1�˒�m��Sy���O�
Qr9�n��=����v��u�b�����
I����a}�v�NS8�.j/�<����~��[���)��^��!��pD�vtpld�M'�]:�s�9��XǬx/V�� �d�,.@����s;e�sZ�<b �dl�#�qC�K"�R�)��Y�i�=����{gO4�[�	9H��{��oUV�Jn\E���-�l�h@w+=խ]ε� |�m`.�E�ͺJ#�o@�F�u;=�f�*��s�5'}��Z}�} [c��Qr��enR�����j
喘�]�Ӹ b�j|֝�g�N��ҬFHڃ���:m���~�>�?�����N,N��5k�W�	����Ϡ?D�Iz5LT��H�TQ��ϵ�h|��]�p9��ˮ��ț�Dx�y�#`af50�t�K0W�w��4�ሤ�g<�R�b�f�s6ƵNV���M�v7?q2���ϩ�`��9m��������K�7K�F-?-�=�Q��OTu�1�C��1������G��p����
�� ������@�?j��(�w��S
��C��G�({��WHíw�r��Ŀ�q"Ƽ(����u�����3�:�t���C4�w�<e�1Q{V�`r��M�~�d�͊S�5�}�}j�Tٟa�^��0g��x�+���Ӎ;��({��D_z8��K�����w�ƲǾ]>��5�>���|:�;v�;&��(SSY�h��,�D[&�!�f�K�>^���I86��0$8���+��_��cgkb%��I����a��c��L��L������_�ڷ&2U�A��ȝ�3Eڀ�.ū�w_�6z��_N�`u�P���p�����6�;�A�4��I��zm���'�����F#?}�1/M�Ii�z�ݬl�%v�i@�J��wW���0�^�R&Q�e��cY���d/�|o�d�����&��E����
D.8+(��P�m�34!�5c�wgaKw��������]���;z��u#�SnC`�l=��d���t{mw�^H��u����xxz�������6��Ŕ!���橙S�nv�{%�8{͝��ʹKOհRX<�������5s��Pts:�.��4��^ˌ������!�1���6ʲ���zw�`��!';]g-�A�WQዮ"lgoW�h��
&�oXQX�B	��a��qt�Z�F:����͸f�L��[� P��m���.18�hLO!�)��d�6ak��4B�яD�Gm8V�kY5I�5{ˮq�j��sJ��WQ�=����5O��?3�~oR�"�a'i��p�����@�Js`�Bһ����j�KE�MU�k��#ǟ�š6D�v_WL?�xg���#^�+a<}�� wR��u�ct_S�GLp҇��k^,y�D�n:l�y�-��@���>�!?C�9�_@�SI��j�5��n,Cݦ��J/69M�.���_��Iy^�߬�K��
�>���/}��\�����e����<@m�*s�R���
�����^l�,hy�`����|yp���퉝��S4,���,W�2ǯKκ�R(��I�A*����c'�Bayf-49Zjrپ���_`���x�Wg����V\��8��m6i�9�� KI���b�����d�86G�7��wr���Љ���>;���cI��
jɶ���-P��I��,�YP����r�f廎���d��.�>��57�������}M>����{0l���y��@�Lj`ke�I�q���V�����*9���z{�+nq�\�����pG��F2�ԃ���v�&9����fY7�[�Z�rT�e�x��ø����}K��n�Fo6�/n�3�����+zA`p�B����쌟�_VlGX������^9���פ{��0Cv'^��nǮ30�C���^u��0&F���)�R�K���g/�	��C�o^�<�i�@����	A(2=ؖ�ƚ�xc[����Fb�VD��O�c0o���z3gy]ա+9�Z��'�����p��^i��t�����r~��䧛j��Vi�����{�cK�w5�sQ�]yU-�K���xaT��Q���Ɲ�m�ֻkG~u#��K��b��1L�>�}�`��q��1����殂%6�FBd�h����o���qotճ2
�wL�X��4l�~v~9��%�t���Y�hi�S�}/��R�-3K����x<����mM�<�iR`�)�������z%=�|w�-�����!=��Z�&8�`���{��7���hҷ��t��Wە�bu��&NI��7x^�Z� �_����] �����:�m�W?J���rn[d4���<]�s�ɡlx�D�I|�<����1�:ɛY[%ά[,&�;w�%t�	Q�yٳ#��x��p ?���{Ьm'�Z����71!�(w'�{�'XĲ.�s�1�QF���q�w0����� �6G�.�}�2���S6�1Hyژ\����}|��3ص�k�K��9\�L�S�Q��-N��wv��u8��嵚�K-��������0t��<h9�a��*�*�u�I���,kT�~f�*rhHٛ~Z�^!�`��Ԡ:��`嵦�5���ꧤ��o9d=	mº��a��}��WGբǫ��ߐ�)G�}!	�x�<U0�c?�H����ں��	��M�L�	|\r,*�e����jR�1���y�
Q�>7Rʹ:-���p��}�:�1�v�Ҍ�p4/��<A���#:�����:�,#>�tT�Kr7,�=vEŻ��V�U؋����Su5�?v�C��O��]����g��I��_�_�_�no_��Fh�b�2�;�r;�v���o&�<���*#J�`�,�����Ǣý㣽!׉׬!�a �94$�P��o[z�NoGK5��J$�zz�P���=/�g��a<�ԆAgkd�$���ޑ�yfY���KJ*�E�y,����s�����ܽ�9�tȤ�ŭ܇�`�������gG����v���5����g�k���hu��;H9+o�ݴT���a�8�$��G�d��iފ��1�x�i��#orZ/���h���,e_])hGY���.���2����}��|~�~?���c��R�{B%�?�&��mᵡ��bK �6FFS���s�crR͆���ǥ��1�}��Z�o>��}6Ú�'h=�6���}p���[G�:.����U�n	�\u�o��Qʴ!�6�g�z"�4�Y�i:��a���Ui�P��?�2G�eY��jM��DK����C�Èuy���U���'�s���+U�"�����Gk���=On����7�Z86N�0�ZP�
q�K�l>���B}'���S��D�65H�T
4���m�/;�u��.�u��eaƸ��{��1�`�;P�R�6��c]�V�w�ҋ�>oC�E&�Y({����%C�]���B�� ��\�C�H�O�|;Q�;z����-�0�Bn��ٴZ�?T�x��ly�ć���󖼄_Qh�]4���`�CD���xr4�ܫ��J<���M��f��:�8nv�v���Dȥj��ܫ���$Xׅ��Bs�;'�N3E���\�3/�_��r�܊ePUW���t��،y>�>����=C^�ٷ]�P!��x���<���dW�������Y�y�%��c���i�p���Y�Rk_{8<R�N�a��
�9��7{6��ޗ��� ��fk!oz^-ٽ(m�$䤍Ԩ�ugIޱ(�����%[����-�4/]7|H�J���AD�_]��Ysk$ =��<���aJY|6��V`��'K᪕�n���X�T�U�2s=�{`�!�S��m:N�v�:���
��$�<�:��h�\m`�Yy�q9�w�G���8��Q�.�9ս�R�>ҾJ�0t�c0u��OJ��vK�Mld��?2�ŠTt��<ĕ�Uv(/�
��'��F8�ۣR���/f2_#����4��j��V�|��0�6k6����*ݠ������T�q���:�!WO/��ׂ��u��Wn(g�]����*n��V�Z������	h���	Ȱ^1i-&fe�7m��@6p�R��;Q��KZ�Z��-p�t&���ƪ���e�Lg �s�<�mDgb���F<���]r�E*ۅqD�.oe`-�`wg��f����A0�&�9�N��심��zq�P�2VN�O_L�K2�CYl��q�I�fuq=%���١dš�V�9�����1���>��V���j�i�25U�M������nXT�]H]ѻ-�.&'h��6��"<�.��U�Y�h75�zj����/U��P�(7��mc%�P6�2W�6�c:.C��cTZ%"u��UP���/0
c���^�J���0\;f�"9B�!�v�����?�`]����r�8,�a���~�̆���Ok(���zum�s8تRn�;h�5�4�t��M	L��:�m��G��H�v�k͋����E�P��V�/�m�*�
9}���i�}�3��Fg7q-Y�P%SN����xu���*��nIlե���)n�����/����J�*��uZR����7[p`'�-�Mc�V��VO�M:�9u�{���IX��M��i��k9� c\���u��%�|C���y"�`�ѫ>�����医�U5�`�^9Ŭ�-i�<�Օ�v�`��T�6(�SRyRc8f�)�7'9+)��Ooj;8u���s�sV�Թ�9P������n��c�$���u��w,Klx��Ͷs\��T,`����a��I�6�Us\u	�r�R��=J���
�6��&}���v�N�'Z�J�s:w^�%1�&�j%T���s��kf�GF=�mฒ	ɚLV�r-"vJŵ8�	�%���ϯ5B(,=(��.B�{�	X��e����C��h|����ƶ��
=�)P޷˶�|zL(�æ��U+����K(��ow#�y��\��V��]��.g'YDD�R�VX]�d̅�CqorΕ�A����6^�C��©���R��{;�V�
F;_�Ą���W�/5��t,�&�Q�}�!��sa�m�h�H�����G�"&6QAAEL�PL_l�QD����3A$�,kE��|�_o�����~?����z=f횦-ccA6�4T3MU�ֶt�Sb4h(kX�&h��^�z���~?������~�Y��DQS�ӵ�TL�RQ��i5��KLN�� �h�4UD��EscA�����E%�f�vDPR�EET�A�(�DQs:
)
Ji����y:)��H"�V���mL�MUT4U�3UUR�LE1,LEk1T4E)TTU4{�6
����U5G,�4Q5SPQ5DUU4AQEV�*�"(���5���J)��QM5V�
J*��)�I���%�gl��LQr5A��:�����������(*b��cDQPLL�m������Zb���)���!����$�"*)�i��(bh���DG'SL4վ��kx�x���#?8YM"�RY��)Sh��wIή��=����aw��v'�Ϝ4s;�lR6�h�a]5�Wˎ&��v%B�]�kso.�T���~9A��(��%	d��1�h��ɠ��\aR $h�U��B$CR8x9�ܣ��@�Es�� x����\�R��������ߋ8d��� �@���_y���{�,��Ë>2o[i���\�����C�@5��(�r�.��=v�2��� ���6�K�|�2#o����L��
�ń��_���\�\�G9x�r�GGM�l�ǰ�#��΃�;`.[DL,s1������D��˪�57�䜼=�����ѐ�wD_�*���`�0>2Ƌ|g�����F^1��^�2g�@��uK��~������n��B���K�&�D�0�ԟ��6�hl�w�}!�|aa�-�xC���[�������V�kI�H88�77 �I@gY�e{i�V@�t�νq�@�O�����8�u�gs���ٯ,��Xʊƥ�B~l.�un!�kY��=���9|�vX��[k5��l�b�h0.}�$��������uϽ�yӽ�"�I��T)_��,)��;���6�ЮY��"�ꌇUq~Ǌ��0�]z`��|�L�&�SsW�!2N]�9�j����M=�����!�[�.�l�Ǧ��t�z= �4ä;��l�pmΈf���*��32_sz�i zJ�)�(n�Uux�F��[>���w" [v��g'�L��
c����=�ҿ]^�2!|��m�w��4�Ҧ4j�V�dк�[_��B���v��1]��b\�p9R.���V�0u�1Y��_x{�?���� �3���"���-�k�,U��"��\h���� a�����0�'� �s��v�cع�����(n*v�f�'�Fm�����@i�3��h{er���������~��f��To>43��Xl���zRv�2�OY��j��	Ic^Gi�>M ��c������=��o�Q�65 �7��z[�����z��,���f�WZ�A{���꽅����UT����NN��`Щ�~�e��,�1Ɂ��zhZc�w�Z�T�ͺ���4ܯY������nj��	MZ��z�hlsL?��9�fY����q�ce*.9<t���9̆N���W����k�J����e轆s>2%��D&#m��'Ff��v�d��t3�t�P���	7���ێx���8:3��yw@������Z�	
E\l����A��e9��6�/�k�A!�(2& �;?P�}CX'fba\�����~�{�a~�x\�;��O�f�g���@^:A��#���PDךE�S�� a]�!bf�j0��Sl�[�N��ZM���$�Ñ_����A��r�!Ŝf���;����z�d�;CyW5�f�+�B��d����1�:�*�98p�p5>�=wI�̺���{N�,F)6�v�o���/�0o(ls��	�Ss�!{�}����x?���  ��qv�8�V{3�r/tV�(X]�;�^8�ι�km\�.|1�A�
���ެ�bu�/�?y�jI�״?v{f2���M�#D�i����Kfa��t)�x.�fմ�y�ڶɧW�kQ�'^�Wc�+���v3�ܱs�㖽���H�w�8\_�5l��O
;y� Q�<�����p|b�e��q��5)J��d�8��𞅾;�amI��n'g�9	υ��p���#P�]m�7���S���dO�o��ƚ&�خqO^��OZ�۳���_�B;{�9<�jf���6�9|$J�����]0C��"�啮�mJ:��V�{��L-���m�ڃc�;�G�(f� �T�M�|hQ�4��S���-?5��,ml`yf4cSF��^�g�3\��ծ�q.�z찏2mg���v�bK��,n�/��TYX��W�*��LZ�Q�s9 룐9��8x���+�`��o�M��d�2A��s�O�Z3n�e-���XU��tPK�<��50͜:-��@`���~/b��p\��F&/n����T��%ng#������y� ���Dw��з �ݫɾPI�Oj��/�feS�l��=��ޘ��J�>��K�������{+jU������f+�ڸ()N�[��t�W�/aۭ�3�U&����(����9�P��ߞ������|L�_�&�?)LHeO���q��6��f5�������X9�=
c]^��|9�Tz�u�{�n}Y���3�����Iz��;(1^:X���g;��Q�v3V���_S�@Ȉ��
)�, ��H�3e����J�����!�wA!�qhI&���n_2`�#T����T!��"���D��BKHC ��{d��K�{�`u˽�X��6~��_gJ��ٳ�G��?^C~u�Zfj�;����4�FS���s�c�iĦ�\��{���{7 zHb�)�m��ٴ��޸��ȧ}-��*Ĥ��2��w%���Oo���N�ʘ?!�鲄�'⢃&>X���UӬ(�^=z���o��P1I~y�w�K+���78:�P��2p��vA�]~{����)��J%�
�&���|j���ⓄȪ}��m������pP�O;6P�,��H"}}'�=q�I�|Q�ug�S.�J���7�ĒW<L(��d��t2{��I�b@��*Y��82��`�����i'�b)9S��O���b�l���=��|+j�o�GY�z�%��{ߵ?�����-���P�mxf��'<h*ک-�I�2���|`|$�8�T�����T���f�R�E訛���L9���,���-Y��:���� a�U.�9�ϐ�+�q�L�Ԃ'xq����������{������,v�H�x!tt�6t?f�K�2LY7XQԹ�4�0u�{�;\�5 ��l�����[W��M��kc�K�(vmZΰ�O5��fVj-���^�O �������L/��=!���1���G4�3}�ٙ�$ۧ�6�y�gN5vA�-H�0������v���(���;��K*�^���u
��5Flo1i{(	�)�	`Gu[]��)���oDQ���"de{b�ٶF���6���
Eݽ^�y���`l�B���ͱ���C��a�}eo�����k�cC �������b`����}=�����r3ƈ�'M@C�iz�d�}�#w:�pm��l�X�"�&9]]��ub99e��0kb�^/�ܱj�������������6=1ጕf�}y��Bns8�[�gm���_2r�5e#Z����y��=�ߕR���ҿ���xt�p���sR�>� �n.�􆬷���C�c�.�(M2K����L�w�#[�y����N���F00s��_ݓ㋛.�,Ǹ���')��{0�-�����srY$5��=fͲ��l������ήE(��PF��_�����E,˖Y�_6�$�&J��Q�Q�����e+�_i�a@�yL�:;�/Jm	���m�H�+@�Z�Υ/����՘�{xy(���T�C��a��Yhp�'3�s]���Ⰹ/'�N��6!�fr��\���=���W�������  �L^�M�X�7���y��0�r^TV5�B~ka���(�3�1���p�zS��W,�����>m{�'���\���cO���i��F��tB�����*S_N�+��W1�ü5����N5uE���3߰P�ޅFC�v��f�>��M�~���;؃��i��;*��ڏ>�"�*��[�S8쿫��<1����x����5o����^ci^2�~��0�Rg�O	��y��W�6_���H�!#}B~�������|]9È�_��7+�N��RSգ6Ⱥ�^2��7N�s�s?>x8{g��h
\F.fٱy�N�	t?<��QE��c��ś�I�W��\���W(��JKGjJxw�k�aNn�噧��>�����l� ��/:�<hY�2q��%Qak�����
kA֏�����>�.��ݞ��5��@Z	�A�?�}c!��sO�B���&6Ⱦ4�Ù9~��_�s��c����Ћ]�n�է���Om	��r��rp_���|`a�9�fY[%�2Uy�K[���[3$�7�U�7!��+��a{4��&�=�
�[}S;���M"1Ť�.zEsN�v���UŘ=��(E3���ʾ����諈��=��NҬ�Ô#1*���e�/4�ms�����,�0���f�����I4_�|> �������ǽ�{�#��X�u{�ֆ|m��ڱ�̙�z��C���4<��0Ҡ8��
��6���e�V��������v(a�L+�Iz&��8��M��,����$�|<�Zl�+z���g�snxW�7��b����(��w6���C�k��	A(4�fN��ouL�c����u��޽!�h�>�8��Kؚ�Ƕ��ּrC�h�9��d�("k̩ ����r�w[q�;�sZ!�+�J�<k�]�	���#�����cWXʩlj���~�2GD��OV�=�k�f�Y�(^!���=oM���uM�k-�_��``��4(>ׇ�����Z+۩x�L�֧ծ�޽൹�Xז*�£�.�zs^���i흠 b�S�/�&C%�g��U����֧�x�[fy�B�[��ʔ�5)P�ȿ[�F�≼u)i���yL��w�q�C�HL1�ȀD��^��2���x�E��ģ)� ��)���Z�ɠɳx��f�D��嬼��1�D&�2�/��W�]�ݑE�?��L��<S*���ʉa����`�Ыհ����N�]]���[�ħU�y�Bt����%h�v�\�kkQdߛjSw*��i}�g#�Z��7}l��Y��!����c>�Z*J�\/��8��j���nɷ����>�v#ۃ����J7���1��j�n[��WkQ]�|�
���� |�?��=��մ�X��Rކ��;��;�B��C��7H�4(�N��v#t�Ǥ�ϸ�z���ˣݲwc�����zj^5�"O����������B5�������NP��PË�P�c4v��f��z�:�(R����z�{p�{XA���s���\�9�F�|�=H�j[P&�7k�Aƶ*3�б�˹U/�|���'s����Wa?��6�K�T��͸�ي���vf�t=Gdc~�T��:��Ց����ǪY�C��Gӳ��/�K@�u����?�w�s}�|Ã��/嚰D~[��^�/�ǤǢ�ŠuW�O���-���Z�-���۱�����Ce<;�����^���ް�#ٵ����h?qÛZ��Y���M�;�T�c�۽����{���T9�L�:hj2O��~;�K�{���JϓY���.��.�Tu�m��qn�ah_e����m=sͻ0j�1a�ܑ�|�*������W�,�6(	��O3F%�ҹ���,-���Jɶ�v���'яV�S�`qm���s��a�� @�����E��b�������dn��.��Oy񾑧e�шʏ�9��F�R��=�6����[h����c����ڛJm��^&�-�Z�j����m�ú�t�Y:�{y���&.ʵ/ph6ZnM�nV���3vj�$��+�|>�_�������  {�Sݲ�0�E\�vu�]SE�w14�L){��TX����D���M����ǀ�����;��z�)���oKVI�QMC4<0�7���h*��tB	�#Ƚ���_�o�ɓfzbӂ�2�x��v��ܯWn��2��i1n,�s�Z��`��|(#:N���>��	ei
����2����'{w�6~��4��]\�/�y�+�;��e}�e���@��4���߻����U��-�4����+��+�a�a�G���|�>��G�9�hLpm�^�5�={N~��f�Y�~��S�ܯ�<4�Z~Y��`	~I��4�|@~j�v�6��=�C��3ʸr��6ʽ�'cl������D�CJ�k;�ҁ�С���/�$;G�H����;Z�[#<96L�D5v�, "]��hL��U="��;���wIO�`b I��Q�񪑔6-�;l{�T������ft���Hl=^=���ȇb�=.��zdR�9�è�e�|�}]bMsX�k�
���Fn���]v20`�r1k��^��>H�4#h�I��23L w1��3�}P�凙�`!�k�J��[�2��R� }e��v��]n���>}��O�T&�.���wQ�5޾�I�5�K�]��z�*ͨ�a���H��/Jխ��y[3�#�um:��C�|�s�_&ױ��3�[E������8�������#n�f���B_��(�\-|k��A�eoรC��5�/`�c%^͠��"l���݆h�;�7��hJ�lֻRR�ZI�$�/^�o`C���E�5��GБa�r>������s���`�|�/�uϯ/�N{�O;PJm�j{ћ8k圥��b%x<�~�>�yy�����ǠW�0A�%�����R�fִ����t�+��3��3f�P�Ο5��aL��_��_���G��h_�C��k1�rd��g�A	��a�ז@�S�]k;���2�r���U!���)���z���Hv@���\e	��i�Y5�\��2״b��z�'�yݰ�{�/۝����a,��ƣQp�1�$AoG�~��?�F�O��⑐]䳾8$	GJs���Qm�^؉���J��UE8���6-��ȶ�э��C�L9�
Δwo���v���������L4�����o@LU�y��&�������qń�i#0�ަ�����f��\u� �,���^o�Kʝ�&
zЌ�"�xҴ���vk�������nfVt�cG���z�u��rf�b9p-.��nd�[փ���]̶3KjB�(v�k�Y�"S��]���NK��W���zg`�dn�4i��5��+���R�q;��k��w-�u���J���[���"��EB�H�D�Q[ͮ�����!����Cf�g.݀՛C�Q'�v�U���jm���k9H��:ҭ �d�b��u���`��}b�Җr����:|�γN{A�٤��n �	k���+:��Qx1�gI3S��5>��Q�Fk�_4���l�.�Z��R5�C�4y��A���|U�t��&U*���H��IE[)޸s�Cl�6D
�V	��	�b�$�w�n��B�M�ēLrӥ=�����~ξ$��ȫ�R�h#�\}Gz�N��_S�ƖtovKM.��S��%b97Ǔ6���t�Ӗ;C�l+���R7fȃ9�~���&!��V�*��f�Q�
�'��c"v��g1��/{/l96`��(T�>8���wj _V�����3d�Dq���#����+RIC��*	��L��K��W!�o9�mk�ؔ��։�,�Z����e��7;q��u|�=r0{/&^��qj�d,^�~F�$�g�e�{��1Yt3�)�K����o�����;�5B��H�0C��%>�<�Agp�WSA%�[�e�U-�2�%�i�@w��N�T�T4��#��׫�o�D�j�����Y�\W�&�l��RS�����d}��4{RGtc�[v����]�]ۏd ]C���O,w�l��V���0�o����<�N�D��]�̜;��EV2t
�ʌ�ϦTP)lֹ�G��5�܈��N�-k��Qs_Q�����@�y*�z�z�3M�sl�"�u�3p��9\L�{s�L�`hy{��*�{�����h�*qї���3N}��W��_�}�@�m8FA��-+9����Lw<�wQ�ÁR@#ʯD�f�f�>�(���8D����M�=G�^��Jf���H�喉�Äx��O7 f7բV�(��\����3@�3e�GJ	������t���%�Qkr򪲩�"�nF���k��YX�ɵ��$,����欆�U1fJ5X¤�$_
zĊ����.v�c��h��.���Ve+f��������rW*�0$k�@�w��O��Kz'Rpd�	�����ե}:0�*<)�:>�SU]�3ܺ�$Ր��:�\y��a�+�U';\�	j����P�v�qĻ9;&dZm������R.e���\�n�Ju��8$�HZ�]�{/L�i�(j�9�G�/���ޓ�ץ�������ý4Y��ݧ�&RD��8,ଊ�m7RشC���yق胔]qJ��hW���x�K'�`�9�LF�,A�4�EE4TQSQQE%-0�<�����z�����~?���������v3�-DӶj�"�"�(�*���r�|˪)���>��o�������~?�����Ң����b(��h�*��������T�TA�ڢ�LESM--��b����!�gZ)��KU,EPLSQ�ب*�m:Z+N�
�5�j����4�-�LLTQƊ9�QU0t6�(���Jk�����"j &��[FR�I���X�N=cIsj���I���v�Q�*d��*Y����IS[Q�u�PTP�I5@���s9��4QE4U114&�UM4��E͘�"��y�**��T�m�F"�;LME�e�����F�c4UQT�RTU�\�Q`���k�5qv���5EUS4�$UAE5ED^#�T�HH$A?�?�m����b<�*��z�V���{��P�J0��f�Fm�*u�Tt8jpΈe^⡽�+���������<�����_O���r�����)��-z�x�<��z�_�xУ~�I�P9+�Z�j����>GjW]��=S��=Z��YZ��Cx��`��[�D�^��]T�f���`�����d�B�����oE�{wVƩx�ځ�o~F�3�?�Íl���c"�s'u�w�Ȏ��C�٩[���{k�>�`��ksPw��@!�+�_>^��	�kJ:���5)�Z#ѐ{�syce��AXe�X�>�&ew�4 �1~U�`�OA|<�cD&b�.)G2r��L���L3�e�s�SbK�0���b!��c���1���˼�:�al ck��B�{�9�� &��yi;?}y��w����	^J(���pE�un��s����J83;�+��R���e��c2R{��^=���֛�$<��#�+�M2٨�j��]r�ժ��̷oOk�y�E��u��9�vQ������Y�|'�:kr@��w�}�a�;5�>���wMvD��o�:v��������g,���0�*��`�,��@]Ѝ>�u_bgk�;�vg��7��mWa���Fվ��y�۝Y���Gf�5����W���	��i>$�r�[�M��٬v	t^��6�G*Ч�j��_��8��>0o��SLk��Z�(e�.7Op�sNP��6�F�/o6'�m�t���>| D��N�"��υ�ӟ�������<�a	���'RrE���z���
{gd�&^޹:���ʋ|Y���"�|C+�<�:������R�&��*q�x����z��~����7��cFJ���8BYz�|�範$��WL�N���	d]g<S��;W�/Ѫ*f��|��뻇?��k�Ɓ��n���K��7�D���~�Sz(�a|�Qu���$U��J����Ƿu;e/Bk�����fƑ!7P�	�}|hQ�������]/K��m�(���9���΄ƵJw栜K�{X[���:`|����'O�;�1��;�'u[w÷��CuR��Z��3t�wy��^G� �	zp�� ��:ڡ3� �����p�d;?�/�Ó��6�9Z���U�	�X��^�I?.�ﱫ�u�]Uʯ}c��"#�-2|�g�S��ù�e��G?k��D�ئ�&��`����(�|�gӏC�sO�T�1a���75F�<�Br�u���v�2:�:��υ���d�^hn��m9�2�Iz$@��(?�����ڡ3.��7X6n~=)�Gv+2�m�PX�1�������\�+-�嚭�}�v���Y�)%z�G����t�)1�n�pu�Uы4�r=M��[��%f����o&��=U��e�(֝��o+G6�\��"�|�p�ڮ7�={��Ǯ�����.s���竾�� ��E��۵�:�rr"�#,+4
9NK����8t���\I��г�A��ߥ�+���?Nmci�H~y����'���77���m�p����]Y� �-->C ���$�|��S�͡��B�UF��6��On���Vl���>y����*�-3�Sg���Lde9�;�{����:���7ҼK��:� �LۆbVM�,Q���i���U�*"���[U�z.�tۻ�;��ڹ���3�]Σ���gXj�N��o��ɩb�O�o�Fcз�x.�{�^��U�]��{���Ϸ�%��@(<���y�������'�bY�R�d�Jj�8�s��WzN��7vo��\�Ξ@��dD��:C�N���96�4�p�M��=y�%:O�"S���ˋ�{���뺱�q}��Z���kk�<���ty� ����%L�m����0Ta;�{�<ۋ�^�<J��G����g��R����5�/O����G�`0b%6����q����e%WrE�d>���R�]�.�㐛��Z~X�y�z���:�M0�����k_�B9��c<���97ى��fQY�ΙU#Nu'rՇ�	��U�ʤ*��\<�a��t���}���������ǧkg���@k�t�ѽ�k��j@n�P�Q��Z�eM���R�*�ȹ�f�[��˖��m��Jgz�����z�<<�x�#��mI��|�c��᧞���cyʵ���E��c���|w �v��g`���;�U"�w���Hq`�n�ڟ�P"u�OH���j�J�(�R��yU��U#2U�ZEܳ]��H�l�
ٵz��pla$9/"��z��[�KC�,8��+}�}��*��ZZp�]�m]߃��._��!�倚��E��^/�+ �:�|}K9�ީ��s,��QS5��d��/�p�t@7@%�E�Z��a ��L���E�?b�C*���X�a����Aˡ��Bh��#�h�����{C�*��Z~�6����%H�e �8p���ágLiN�\��2�Y��]#k�O;P	M�@"f}o�i�m��^��=@jm[+��3pa�"9�=����5s�͋l �$PY72W6�gY뷫P�l@�l�����3�r�vr�I0<<�L�H�(E�p{ה�ܼ>Z݆O^YX�ݬ�w���;�S�wv*g]o�^ʋ����f^!�]%�W�&'��.�d��\��A����>��ȳ~?�D�I3��
�u�/��ڸh�<0u7j=���]���J�����YU�4����x�0�5e[x��є6�v!��Z�wE���G�����n�\窌kG[t�~yQwU��o+So_��l���K'��������� ��� x3{�Sz�S�����/�7��s�T�SP]s�]��uO���[��������yUq2������}|f�E�������I�+T-XUE8�ئ�d�J��H1�0�X:�%���6���#���1CnY�4ީv�oQ������(�Ɓ�GM��|���/OB�7oܛT��h��K/Fz4'���	�Cv��&
z�#6Ⱥ,㛀Z^F�����b�t��B�����p˚y�p�`vd�M>�!����T�F��aTJ�Z�\��iIc��S�:��������ʫ�Ѧ�X?Cd��;(�T��7�>��V�BՇR�Ţ����s����٢3rb����yCn��O�� �P ����Oǟ��cNI�/Mϛ˛뮮˻�:�
��ʲfcn�n-y�Ok�M�%�?0к��sPw���y��F�4��s���@��6�6�ؽa�P�NN�־�>�t�:.���KsP=�z,��&;��ȫ�a�V�da`+`��bur3j~��v��vRa\bK�0����fN��5�-���c�4w��5ǖ���e6=k�燋��q̊��&g�:�ە��=��>�B;����v�[�����ۻ���'tȾ�uk����8��F�Wr9���n�9���k�Y}�/�eB�oW�y-��y�E�����:^�E�v�� {�� ������ΐ��l*�?|���?��$_,!EG޼���\�~�Hz	/H�8z���x�p馁[��.�m���2B�*�mẼ�;�P��e��}��߄�^=��ƴ��D8��s�����z�T�f5����4!gk�����S_`�E`^"���5���
īU����U�����|�,o4��Z�jK�CK�0CY�(�Ty����	��M˛�O��p�k�!r�/f�>�������PǗ��[��!)�	�
N���c�ٯC�ᩭ����O9E���e��*���F�Ҙ����x��Q��!	L�1)͂�0MAJU�w7��n'�㎴���i[n��OK�w���ή`�{��h]p|�0O|��קze'Y��,��犿9��&l~�,b]�H��3���:�p��a9ml��͓X.xb�_G�C��.��Ȣ���"�ZeݫbF��<̒�a�nj-�r]��-N�٩�����	���M�/�
8e;�����������'��������a�`����S�0��a��C��ǌ����~_uտfҬ������Af�kQ��u���&a[\twd����ɮ�5��W�o��ֵ�;ȿ)��YK�����ߡa�?�#�:��KxK�r(Y����εg��w��]g+:��Z������#��9 ̮X/��={ן~;����8~����9@�r��zw��+s�	t�����d�k�r/�6��8j@��-�4��v���*;��ҡ��5l�l����/�B}�xFc��M��=>>��`�ܩ�eл���ze�Mk��ͰeA/t�J9��f����6�.y]��,����R�����!�?3�6��fx�1ȥI������3�Ǡ8�4��K1��Ɍ5Oh��CwMeb��ڽQ��_~�O������<���g���{(�[���H�����粎;���vz]����X�bƃ�,�D��XF���}y�ڿ����9gP�Hs��yO+��sI�8n�Ք_4	5%�[�F�Mup��~0�1x�Y��̵<�l��9t�u�	�������q��(�è%���zK�y���z�m�ֆ{�8>?��G2�°=���?��LǴ����Lz1��f���`�Գf��PcK&�(��ٴ�=[®�N�p$⭞T�8�،�Ae��b�Ӧg#�j+ӼD����ɩb��(�]<�����R�2$$#j���ޭ�P�]�� ���0D�����l�+%W5tB	�b@d\��%�sk���K���f��Qo���|�x�Q+����c+�v�gD_��WA~}����C	`؜����v�w��M�A�����#��j��W	���w�c��3]�M����[we��R5�;��ܔ"�4�˺�>9.�94�!���WP7������������[g����W7}茷��-l��[�	!D�f�	��|$>��~���=<[*�S;P�{��c*[{��|��-�.���#�|N*kps�ǐ�O�;Q�?K�H��kti�^��k�2�h�ÅWJ�>I��pv)P�\Ú�1e����4[#�C��Sx`MsuqO�����7<�^�v8�_��}+��y�{K��(�7]4�O@~m�x�/[1R���M�mɡȲ��
���zuM7X�5�ga�I�n�A(�zO��Ļ��n�hn�v�v�J|�s3zz�3�\>`�ً�ɑ:��n�#����}c�ɷSߢ�_v��!��>Qϭv���,]������"~��<F|yA����ʢ:�}zhZc�qx�X�� �覅l�6��_~��mx�[A~�=cYA��H��T?0^��'���������"l��͈����q�ؖ$ ��5�^7��X��q���#���Ag�V��9Xi��V��du���ǐ;A��T&�3Eڀ�.Ť�0�A�^���{dD�#�����@�=��j˞'�2,��\}�̠���y�>�^1��0�`��	$3�����.���-�9�@�ym�y�����`����CCt�dQ�iNeo/���S��+F�g/��
me�q��@�=y9��bW���G,M8���G� ������?8���2�������M�LasM��������	�wI�d��G��ړ�E<qۈ�@��ӗ��9�j��j�d	���$��� cQ{W>���ZҶ(����!���z��r�<f׳w3���ۏ�}hQX�T�����$saq7 ���l�HN[q�O�ķ��zg4vwW�S��?é(�Q�.pV��b���c?�?����!�>F��4�k#���U�6�����Q������p�m�^��.oؕ
Je0�[Qm�ꋇUq��"zBa'nj�y���0G���>�k��L�!�%����$�b%9��ZS%8��l�	�a��*�N��A�kP�w_.��ާ��}X^��5*�f!�T;`�i2��LU�y\�2	��/N�o7!���Mf3��M�.�CD��s@L9�C,Ɲ�vT��~Fm���I�ԻF�)��Es��U7&/����N:wL��m8:�!�n�	y/�<hQ�a�B��W(��&x��\��ԩW��1]�/ѽ��6O��VQψ*�X:n0ހ���%�㌊:��� |�c���Q��;#�aY��{31j�4О�`�SN�Nh�M��ݦ%�j��:1���:���yVDG7�b����\6�!��Ȓ���n�,ߪ���n�LV��1�O��U�lsqP����C+����NG��g��趫(S��*8>S$+*�6J�u�X�|��|~���������X�&72�yk
��?R�gfb�������A_���-<cTcNfss�Yf#Y�Jb��GE!e>Oc�~�V��ނ^��*9������z��|�F�3�a�e�ʘj�]����_�1�k�kP�P6.�ǰ�3NW�Է5�,���d��ֹP��j�,�'�:�� ���3�e���,8�s�	�nǡ��KP:#��<��u7�fj��B���o��2�a�ExK�zaQQl��گC���y�� ��<����������&m��O��6�
�e��3%'�ME��X͍i�Hyj��v�2�ځ�+	bZ��n�Z-ק�G
��M�S��t�ê�x��zä�b�h��F5vLhXU�̚��8P����%�!��=��LyW�ˡD�=�,�G�뎚�tS�Á�)�Zi�Y8��3�Us�g�.�#z��[��Є��FBeK
OaQ�g�5���6)YG��Kaj��a���?���O9�L"E�y��<��%2�1)���L(JEld�:�!�����:6���� �.f�U����L8!��t:�{�����DV���p�9�ij':�C�[�yf��2��&�2rGyb�OJۺh�}���+9I&JZN�p�u������	Da��A=��`��yX ��F�űYF����R�t2¶2h��/_M�U��b`��6e�zջ��ԡ�nMޭ,^]��vʚ�_ ���#������N��]F��W���t��U�|����Dz�q#��ԖX�/N4���j7A�
S��e�H�����!{׋�6��Q��J�:��uº��K/{�vZR�En�vPm>�1�޳��P�RC���?m�r��:�졁#��R�i,��T�g']�JvX�Y��E��y��\n�r�!
Ï��j�͍U�U��HNR���+��H]�h\i;.e�o.���L�z�,5j)숊�������
�)ܿ�9J�K�DG̛�*�
=o�/��^Գ��ܔ�;��p!����u�f��4�/.�"?WO��fFq�ԛ�D��-���(S6�wCGIy�G�e7�]�_��MF$��K��w��Ǥț\��]`k�Q�q�*_-<-ؽ���c!/w-LV���S������s���W��c e���I���ǔ����p���go�����2���ꈄ�.�g�[VQCdj�.IPN��w]X�b#K�1,cV]�e�I�:�i��R�̹bS�%��<���[�#�/���'�so)��sqŵ(�&��M�Xb=|$����]C�nm�I
I"�t���L�C�s�/N�6ͱ�߷zd��T���,���	yM\5`�:n+-LeYM�A�Pu�U� ��9t.�`�:�BV	tڬ��wKx��۔�Z�"V�o3{��:fr���:����r�eq�-���e�vT`nf����i�9m�D�st�{(
Z)�	���^9mSս��R���aWO^�:z�a��5&k��*�i�Wkz�,�c�F�����Q����� ���n�f���ΧBZCj�D�wmڜI:��ZJγ�������^�;e�:+|��`�Wu�N�)+��L�8��E,ˎ��LE�rj�n��s��3/Zx���w��E�%_j����+fn,��^�ïQ���OȺYNPvDW���K�5�u��Q'����v���pgC�u�yx{p^7��X���)�:0+��C�|�o����^�a��b�3%8��&F�6���BGX��Sb	p�n�WT�c�ޒ�,��bB�]���&�6m�CE��C�m���I���ug��[�Avq��@�u6�7�;G%�v�휖�\'gne��%��5���U{�:	8�e���Sj��ի���!�Z���w������V�[�+q�~�2�n�A6��+pu;���Y],R�(���3���|�v�������sa� "1��#�W�6�hg`�G��"�*�d��(�
�"hj�l�TE�����}�~?���~?�����j�<�DDDvtMk#5):�D4��TE14S� �`�1-^v���Pm�������������~�������~�Ҷ�I!�:��b���14�����b*��i�K�)��. ���,�֪�`� ���!������0��Ժoi�*�b�H��"b<ƒ�F(��ulUDG�ny��$"��1����9���Z"�1kMULl��6�M���QQ4EQ!�QRPi��N��"ib��<^#�D4��SM4h�T�R�qPy�Kɢ� �F#K�v�h��HR�R:hW6Y���O�x�-gB�6"��(b_⢔��j�&��(�4�+B��4Q%��%��Ԙ�h�K����_8�<r�<nx|��IHK&~�G�4�P�b�F��h)b�W[�&e�J����-^�x�L+g`�k-6�qk5Ӊ�iP}��F�eI{��4�ci��l}�gYJ4FOБ$!��P�,E_�k�!�ĕ$��r"�Q�H��&ns�-�'����}?��3�
��G���"�Yܙ]��rՎ�&j�n�c������H|��B{����5��):���E�{@��c�7aV8��*��f�l����in�
Wq���j����N���"�%�n�|$J�}E�GdQt�A�EH>�?�T�^??@�G)��MM��)x��	Qc��'|Ǫ1�����+��+mQ�����ٸK��&]�O�eAc^�)ߚ��w��C�0�5��z8F�j=�y�E���o6����9�t�zKj�P��2�j;��ҡ��sh/N; 8�!æ,���i���P5y ���ѦM�<��`���,~J	{��J9���Y��E�~̓7IZ�����M�7 ��2�����%۝4����Vt� ���'̣�����q�sT��v3-]�U�n��wLֲ,3����/���'�������������"��'S�N��C[��
o��5v�W�P>
��t ���	E��4}?s�?��4>��؛�6:[����ζ%��k�k���f��7C�I� �PŴS��"���%�Z�OA���|d���	a����̋!�����7���aO�I��3Tm����w������n�)0L�Gc;.Q:T��~�'��o�	�B���ɬ���c��G&��$#S%�y�љ�F`�Q��U��l�mXpv�9��Uݳ�;�}���x?���{�&J�<j���x�dc}���f��,;�YA`Ç�y/�\��`�
�h|=��d9+��"]�g�g?@ì�lu9�����{ˊ�l�7M�-E���I�яV���YO�wv���t�2{��h��^b�Ҕ�0K%���D��P�&VbK�+�мU�˙�������G��Y���8��"P02}b%�Ȉ��۞�FʚnwA8A�E���Dȉ�:-���r�W��k��{kVW�{�Ơ�ߎ|�Ȝ��	z�<���$��fB�_��{u�N�j�\_�׶"K��S*(�kk���8��������c��OT~�{�ʡ�-X칰��{^�lOK���c�X�RO�"��
�+����z,��}��`�ퟄ�c�+K���e����VY��g��߰�v8�_yE������r��>ᇾ��ٍwwD���p:ý�L�����^7�[��ʵ���E怵-�����PKד�9To��򾗯������>gad!��y�d�hM�
��+�t�k��k��I���o&�䭓�-/V݃�v��7��'eX�TV*;G8� N��w}�R�I4+��Re�p��J�u�����=k�a���.����@=F�FR>�	��{t2�l(<]3"Ψ�n��fvhɗ֣y���X5��h��+U1L�}"6�Q�gۺ��w��x?��<<��av�m[Bf�fd3�|퐨d[�1�a�8A��y����K��^�Mo�s%����:�wЮ��Imok,*}]bWs0lf��a� Їc>�`ϡ�<	�(~mO�K��]��7��4��ń�xs�W�+y°��0�x1�]�\|xR���a �&S���E�
Pȷ�R���o&H���L�}B`+5٘4����T$���w��]�I0a���_9���.�V�K�U �Ks��6I���7}d"`�V&-���͟G�/�MwI�jJm�j0��|kN{���k��M��/��+�N�9�PB1�!�-�{���u�ִ����!�J���uA�{%k۽��Q����}{K�V:�)��%c�e����@�b�)˃�ȥ�����Ҽ����}�c;�b�=\�i��B���;Z�@�[�W����\g�
��a�!��g�4�k�34[���j�������.�#�n��b��ĨR�]�L-����^�-�q��(BoEA�k��.�1��LԸ�,�fB�soD Y'��Nl�ZS%8���a#�-�W�p�������Ju����fү�'�̫A3Fn�I����ɼԡLk�R�Z�q�#:��.>�JC�q�=�����/ۛ�'��@�enL�ܜ�@��t��5ڦ�cf�5��/9���g˃����n�*@�Tljy�`�'�Qښ���1���������{�b�q�ȣC
o�>��D>3[-�t#��zL�<�q^�E�4�cq�e�wf�{������{WC�n{ܙ��fv�?C�9�\C",�v��RSգ6Ⱥ,�!{�i�{9��'w�l~��_%�r�e��C�Q�ܪ)�����I������eʓ��6�Wl�v����ö|}��3���&����X��n�qz��uBxв�i֔e��ԝ-�6��9f�L*�O1�[�f^����h&5
�Zz���������^f Ic���7��b��L_Э�pcҹ�Q�/m	���.�:�9�;���0~�hs�j�C�1�9SO�tC0����:�0�ro��kVqT��t]�/}ƥ���/^/a��ݞ	�'��.7,�f�Y�4�fXHy�oc�fZ�e�ei�i��
����D3u�a��2�Ds���)�&�	������S>:�(����~������N�ޱ�H�-_C�$����?\A�����Q��)� ��ra�����tM�1�ll�Jeć��W�,�b�����!`�r�Y:��Al�y�[B�Q��~#�Kd3=�fS��\���mpģ�H��j�)
�e��23;��VQ��Ɲ���t�0�K8�`��n!ۄٶ�Mp��]��U��O����}�.����C_��Mh��w��8�����&�'�RzI��t*^����W78MA���p�My��)�WL\:��L�����ʹsR�j�g�Y�	#{o��C��[k�;0
�e
%I���l$\�1��gA�ka7{��j��6�S5gs������L��0�r��D��FBcAb�I�*;B�ǧ5��e�K첐�-�O���5���2[O����	�P�}^!��soB�_�ħ�U0MJR�k�'�ɟ�ܨl�3��-�x5���#�#u��lP�!��zȃ�qk��wd�^%��ﶻv&�Vj�v�n��%�j��)k�B����CV��8���rg�<��;B�g�VwܹO�f��.�������Ω�:�tY�vE�\���ׄ������>����������}���\*��m�! �n�w@⮗��i��rčR����8�xb�ѴG�<��s����ቷȕ�zg#�H�p�1S�FA`�@�r�߉Te�Z��3*Gs�Y�KӇ��!�ڑz��a�gŗ��iOpV�a��p���b��Ml����,t_��Ҏcsڍ��ڜ-���_�I��4<}����>��ux���M�([u�.	��2���^���ͤCŘ�X�m��פ��A����޽�V�N}���f��l�"Ԭ��$�V��oe���љ�1T}��҈�Dл�]ˊ��*Wח�t�P#�v�7;">�}��y���H�),[9^R�7뀂�a?����CZ�4 ��n�eqʓ����z1�[w�UuL���w{���Q�z���~���@�<�c���55g����y9z���e1�&�[�6�ublo�v!�y��Í�LW�LZ��;��xA��ň�6^��(��x������"1kws�nW0��[�D9�pF��P�}��lEC�dK< ���2B8� �)���Q�f7��v:���qHƼ��i��L:�YA
FL?��YߎÜ����Q������a^֒����Ư GL����&���B�1�%,٣��dS�vHs�ٴ�Um�n�#�O�s�j�؜�S�v��b%������%�.==^5X�+ڊ���l�r�5yb�NM�\fl��kkma�4Q��͟Qǘ�~�V�*��1��2`p���3��<��P�U�C�N!&kun�=H܈���QW96�a3LT�M]���X)ZF|9�NP�����Nٻ�R���l�Sg��:��A�$�G;�D�7�|)���4�����_"��s��b�}	ܕ���T�iC�/ܷ,nW�j��cL�Qiz3��	�uY��i�ǚc���OIT8a鹋��˲�j���R����׍���2ܕ���y}�}E���d��M����� S�h�+d�nS8��޻����_�������]�F�<�~`�1��Y�fB��i'�I���y�ث�J�;��W�`�����m�m~��_!�C���9������J}T�I�M��9E��.w���.�a:'ۀ���SE]��|��}L#Y��>`�Z}G ���k��M7g)Ʈe�ԍcA(�|���γ��9�i�-v��q�lK�@��5��Ѕܠh��� ���:
=NM��,ߋ�{���*�7y=��(Ֆ�^��W�s��d�T���ͳ��p�W��XAλ�[��%�_$M鱋��j����0�1�7QaK��v=��}]rk�|_h?��C�k��P���Bb����9�,�Oڴ1ݣd6������Ȃ��'��"eq���nu��BTn�����]2��wU���dR�U5u�։�̍gP}|8��դ͗l0�[I�$e���oF[;B�����8֍b�4	�x~NpL[e9�������M�H�ɜ`=��[u��<�Zϧ<Ϩ�*.�j'�.Bq��7,~j��&�}F��ZҶ
:�[��"{����p`�5Ӡ���Y27�$�7�mV�sVc�]ҳ�+�=����������f=�yF��7,��롽U��n\{֋�+��K�P��9N���zZ�:�Ӣ�Aw�Mt����.�y�튆:���Jjo� u��ǆ�n+��{9�T��\��p�9XэOOq{~^o7�i��g��V��8�;:�Y�`1��-�<�zw�`��!'�C�=0�DϮ�8*����=t�Kn��s۶�k�uj#_��AzYX�F���S�g�T\9��̂qub$���G禎p�g�?�0fh��+:�,��.����C,}�'X��D*�u; g�m}V���L�4���}�7���ss�x�)�]�̉�қ���"��Jse*
��Jqo�L0{r-��:�����bo��v�� �\;�v�6�ޑ oJ���LU�y^��C��k�nҮ��'[У{��;#HC�kH�)�LȾ�,o��u���E��]X������/�i���;5?g����ʒS?Ό��#���%��|i��o�&����:v��u؞fj<��7;�`%�.5y�X�kT_������&_��dQ�l:$]�;�� ��'q��%E�z�O1��_V�<�郕 �?s�������p��q��ޣ����%[0t��S��Xs&�W��a(%�Ts	]Bt� �����^������ad�!�v�B�[*���l9�}w[&�X�9^<6� �Ew��ȫ`m�͘[��%2���}�r��p�);��:^v�+^n-�OS�b��:��)�V9��c0܈�r�;�)���
�B�.�S��L��߽�}_|w6��#4T��V|��pJ�fH3�JF�B���_~&ŨP4aD���VW�C9*�.�ǰ�	��R��z�����Zh��5�vj��P�T�g�`<!0��o�0̓��;d��Qa����f�s��b�nùm��Nv���S���<�0�,��~xE�����m"��0�M��0�be�]�ӳ>�����8{͜���N�_�}����'�^���|�*�FT�O�n{L�>-go6��I�Sq�Z��<��HA>m��t�P���Ǭ㻳Qa@ ��Q~n�Fbr۔�4e�Q޸h=���	�醶��H\���,��8��"�h���5�L�Ϯ��\B���Hs�q��6�{d!�#�N�266�XN��Q�� B�B��T�z//�{Xڭx&v1�;\�#�M�W/�|gh#��yį>P�D����9�t!)����R�&�O[�2��x-��F߂�k9��ÃO��W�����XI�_H�5�ޙIщ,�H�k��Nv'+�Kov�ݎ�tSu$i0����!>�� �5ȈL�{}Q��ar��m�}����C�2�p���\�V�dK�D�y�%]�N/J��l̆��sF�2p�nS��ysvqU5漛o�� k#��b;a�4��^��#m�=יM�DQ&�e�:Њ��n�gF�A��q�g(���yȝ�hyv��ݡ�~^���q�]��n,�E�긤�3�^�e^��f;�y�78��(`@~�T��a��1�S��S�nC��I��)^N�@8������T45Jw��X����Sѭܻnr�9�]����B���S��sg/,�|�2�-F��*�s�Y�|^�=�g�k"n�ob΅ר>����8~���Ķ*��L��i��+]'%�ҁ3�n֤��������tͶ���CC�J�ݛ]6{&��k:m��9P�/�$���9/!��-�îOn�^���d~ wFM�Q�5�W���/���~7U�������f�qGu/�Yw9��bώ���� XU�y��Сレ4_�M�~a�踑�˫�����ztԳl��1��f�}���;Y揨j�a���ı�=�S>:)~�n�쟜.���P���l�':�H�;�j�v��u��E���ϴ^_S4׷���K(!A0�wl☷y��8��n-I�eVl��t8F4�������=5>�z�1�rT�Y���`[J;A���`�쁁l���U�斫�����*�7wo�N�qV.�VV�	�]��n�S���]`�&�ũ��<1X���p���N%�t6�ܜy�9�CK���̥iY;Γ���l�R�0uH�BS����Nf$V�n�wa��J��2�uV2G6��Y��!�b���|'l�*��.�A�Yߊ��Sf�EH�=���ɜ�c{:K�.��M���˵o}�y3o�Z��ܴp���ov�T���v�ڊ�}:�#sh�d=:�{\Y*L�f�Ĳ��O]^=_X�u�/��cnf`J�s�Ⲱj�r��(�/4E��j���7D���N(�Ր�,9����7�8{d�ߋ�k+o���Ao�+*1X���C���CX�����8�0�r���Z��>y�^Cw)��f�mr�C���]���n�-�����no��|!=d�S�̗OoR��t��C11����^�u5^��G�`��:��i�D�wT%�˱���w|U�P.����_7z$�ջ#5�֙�c�g;+M�b�ۦ6�d�w��(؄E�(K]���H��n��u���U_g3x[Q�۵:�r���B{sdj��Etj�,7��#L�jf�qK�v�4�Y��U�<5�Գ����Gj��G�o�W`����n�ޥ�k������,���5B�"�;vid��篯w,�P�ͮ7�x,U=����E�G[	n���:��x�-:Te�����%?���~�ʝ5)�e��y���߻~�)9�V���i���=��;+NJ�\'tZ�c+�Ιi,�xt��茥vh�x1�mjX 8�Cc�̨��XE�ѕ�V�ds���՚�ul�#�0 ����yTj��3v�����Xs�v&��:�1���D.���x���K�hV2���r�n�Qɴଛ.��e�E��M#� ���gn�*�N�C����}���#��t[V;	���D͗Ui��{l�5�������*�Y���޴W�)ٛ�?�f�nOZ�S�n�>���Aw[�όO;�R��=����z&��ۖdZ�1^)N�!�U�a����e֥A�M:X��Y
j�w��\` ��VaL����
<�,ʹ�����K�0՝R�mٚ�!� -n��I��{���&
��u�b�nón7� ��e٬����輲�0��s�����p���-����S���GH�򠟋��S��y�u������2v�{�fl�@V��em��H(�tv�f=ڠ� f���5�/�Nڞ��
�/6�<:g<��5���OiZ+���Ճ�r�����9\V��X��r�*� ������e��{�yTf��E;�Ӹ�.�&�zpZԑCuV&v�Xt�%���NJ�R��u�}9���i]^��*�wa�l�&d�dr�B�^5����-����@SII��AP5U����
��=N���Hg������~��ǯ�����~�_�} (֢i���J����$�����ׯ^�������~?���Y�����T�?I9%JQQ!T�v4y�H�ITQDG��lU!CUMW���SUI3MRz���9t%�E	EQTT�RP�Q4SAAEE5#TDL�Ĕy�4��Sd�"<Bkԅ�E�%�8��)b
y��4PD��Jj����2hJ��(�!��CT�JRґEA@M$4�EDoX9Sk^6)*�)���Z|}���}���v������:�Z2|⇥+c��Ѹ-O����/3a��=zvnZ��,�W
���.ٗ���~�������b�w�w������猯�[E�%�.=2�����%6��MDP�[uo�-�ጶ���s5^:��a^�ǫz����vgA@�"X\���.�o2��\ݍ�͝�.f���f�[�n���Dk����~IM2R�<�~{��VWʍ������9b?��mKw���KØ�X֓_O8@��'���I��Nl�S"���|����� y�5<�<\�K��ڞy�,���ž�l��̄=�S�FY�N�q�&Rr�(sȥEW0��M��;���؁�;����?Unw,�CDy�~n����7�$�_)v�nY'����h�ع�nNhX�Ij���,�s����60Z�9��-�k>��w��w���g*G%sͨ	�=��.��6�T�������ۚ���c�H�vQ�c�[_�H&��N�M��4�'�C���`�Z�S'C��G\!�Nq����SlEóH�`��?������&tگ�m\ω�hb0�Mo�x`�1�P�Xu��ܺ}U�x������DǎO+���HO^�Z�y,��ӗ��-��2:o��弭��+X�1�R卢�0�s�C�X�Eᴜj�!�9i�,̏��-]g��;k������̗7��ۑC���Nbbu�={qҮ��p�a!�[���:���B�E�a3��X�����޿ �<ky�7�4َ�ؿI�l��7})86ˀ�aH���1\��_��P/a�G<3�K����j�w�Z3��p��|��Y�mל�4	x.���R�O_����ZWFۡ���p����=�յ �#�/>��D���/���zg� �v���Fl���D绤� ������Rc�"�k�h����{kס�6�5�
<&Bl#�ql���zn�q�9���gc�~d�M>{��\�twV��^����I��y4ʇ@�t��zw�\U�I��Q	���rg�H�L�����>}��e�_���	�,�,h�Z�F:�H���:��P.E���d
��"�c��T�2�k�.��q��&?;�ε�&�[*��R�U�)�T[`ꋇ��z�NK�ʘ.�����9PR�C���}�l���-�^��=��Nl�AW��O�vd�
�Hʎ�e�;L�;ݯ�Rӽ�����7 ���e"�Y�4�{�~jޥI�'��U�Ȣ��a��h�^b��{|�w�q縮vk��5��8�!�~�0���B�Ԍ�=�B���2]*�L+1\����}ʥ���r�pP�o��%?Z��lg1s��1�:�K���4�]���F%Em3s[G��hQ��C�d��+�a��^
��M��]w�_*��h��>k{/:v�L���������|�=�S���Y����{���)�d��j�������F���f����a�2�)Ό*�*�~�O�re���V��wa�^JO-f�)���g�/'�q���m�]�m�q
�c�b�x�ge����{�B�O�+���.�*�
�y��*����3��T�z�~�Xw;��Q_9T�����6]Ln�{�-1�n4ҵ�(%�?0c�&��ß�뵂����M���{��s �C��pQ� @~ןC������s٩H'̺k�0'(q�n7Ϋ���ʉ�/ޝ��u��_k��^�����	��
Yk�2~�KƎAz����$���8S2v��·CJ�=��i}} �����1eyNQ'��hY�Ol.*-���N��U�3p\_*��7���!y#t=��I�i[H׊�D�c�l􆐄^��	<n������% p���p��q���lr�v5���X����<�Y!
�&��q����NK��
x_��kϧ��3=�j�>�A�byצ�J�/j[q���:W�eG��E����E��͇^@En,W�p�~u\ޯJ��r3��o췕8�붭*(�[Sox+��h�KWj�c�*	d֨e���̷Ov�������2\L+M�U2�!����4�M]�d�Yr���	��V�u����љ/d�>�~���S9n��vi�l�l�;Nut�R���;��10�v�s%���b���*��5��+�:��Me�~��9�k�z���{gh@űan���|C�p�����%5�K�-�"��e�FS&X*ԋ��1�;�_x�?zw�]�K�Ɗ埩ZL@��tC�	�����D�����Y��f�̨�Y��?c<7s�QLJ2�6<�{����8x�}�-z���W=��爭k��뎆� Vܗy��0�0��g�+P��N[C�mxw��3
|0T�C4�uzC�Vv�x�w��@�tB��N�A�=/A���
�Ic~����V�2��/|�"o�&�gd��:���[r`��΃�;?:��a��9e�Uzk�U祐9��w�ڴJ��x��M�r�C������<���X����d��L;��V�����}Z^�:b"L�X����yn��P���!�9��<yF����r�g:?k�u�z�2y��]��7����ǣ��^=Rǌ�	��~�(ӞT"?,���(��ae*�f��͒�[lr��v�����W׋V`���N4���sVr���-^�t���-]����毈@�\�˻=(I�8l�n��Vn���W;��{���Ѣ��sB���1��q�m�|%�ݢа[�z�d�#�B�7����~�7��;�!���e��� ��\��0r�/�5l�?�s
��*Yg�R��W8�����[��.X�͠�9Ռ!���8�$��-����MՎ��Zz�J�g��roh���FG4Ö����g��6�y},ӃzKJ�!�ɇ/"��Y����H��{����/>�3�(Sg���'�n�^�%Oӕz�1��S5Y���M�-���4�X���	&�W����~�Y��=F`�4����E��q�)�`M�@��Bl���l)x�S�ٱWuhjd/�u�q�P�<�V���D���\aQA��y��
����`�dSަNg�=ʚ�c���:w)@Ȁ�|���~Q���^��ȩ���A@L�٬ب4;����_b����[�A/esן��Of"S�H�U�&��r$vEê�G�;^��*�ݻ/��ơ�e�a�1�+e�)���GuI˺b�C�E**��5�.�m(��q���gS��m��۫��m>d8!��	���ٽ�)�_)v�[�I�r�O���ox^��U15��MG}Ǩ��Ph�_��wUn�<�����)��LS���ֽ���,n>�6ek�m��78]������BnSS�gI�ht��'��a�5K��+�ٯ7.*�]J��\�ڄ�N�qe⎓�	{�������/7��Wv�l�;��A@��	������>zw��`$?j��(��*8��I]l�S�X�˽Ӣ���M�5����*X�cɤX�e�|1��:�vM�ȝu[�����t��r��ev��N�y�B�{��Ҩ��wChv�:H0|���o+�Q���OŋۦV.VU^�w���𖾬b��V��w�����_�����(/�m�� ���O,5�,�2��{��� �c;c�]��oM��)��]4��}�+����b�8B��X�&m�n��R�b0Gpr�7���>��,P^�_�ι/��&�:�e2�_N�礼?}_�\��ҕ�1�J��k�ذ��>O��_���	���=5�7�>�y�ơ=�y�R��1M��cZs�ўz�d9���x�74<G�<����Z�`h�3��[�'�U�9��j�^T�h~���q���%�CW�2o&�W@�t���V��,����x�9>6!�L�?{A�"�]PڊƤa'�a�ۄ�@(ֳю�shlg�
<,�3t�6��p����en���L���\`~�������/2��n�s}g�)����V��v���MAέpV(J-m���;���?|�(��z�`�0(U�\ʸЮ��*t�M=�-H�6���[M�;�.��KY�D�ixL�2�Ɇ�gͯ� ��F|�N4�P5w~W'�_/nn]��qt�,D�3� o\(x�i͜b�����!�:�F*��R���
j� u�7K�=�WK/"�+�)�c��Wڹ;: ��cd\9N�/dp������x/ȥAPS%8��Sf�)CĜ�}�ܷ��s,�4�z=!��� �!��K17�D�J��xo2b���cL�t\J�骢칻w5��սM�خz���c�{m�?P�s��	eWƝ�30	�Q7Q��o��Qy���Q.i巜�x	�iGf��?>�����_q��)��������zۢ�<�P9+�Z���\��%Q�qC^]�{�]�xu0t۶��g���l���cy���������']������fT�{mi���<��Pè��w�z���U��>�����H0gy,�Ll�/UL`ۖ�7�贠�ƹPXJ��\pv=t+���Gk��We`�`fi�,G��`��|O0���VW0MY�Q�5�GƯ_�::my�G%&3q;���խm���*�^����-�
YK�'�G%��(�d�
6�'�h�l����ݙg}�}	FeT(*�v&����gu�ݚ4�҂����]䕠��f������B�$�KL8�fuG��fs5��5��-e��-֦���Nj��z詡��+2i�u���=r���[��i#%�+a����o0��f��F7�n_��f�z&d5�9��������<���S�dS�g����e/�N��)ki��T�4o@���CN�{I�`V+C��D�^0O��9�w�=��K����%!����c{�O~�݋��Vs��y����<��HB�&��q��t��_}9��5�P.��&�m�{�� C�8{���&�N��5�r���aTe@�:��b�M��_:B�q��ܨ�(�3�-�X�L�� ����J��U_�_����u��s*X�Ry����ǍE+���߷�+���x��R�4h��hQlXC]��H�.���9��Jn7u��
sjN��1[Gs�^N_�,5�IT-�*�Z���S�Hql��~���A��R]s�2�ή^Ws+]`OȾ��<Q��u��5�B|��f�t�k���tL�wkd����g8r��b_���p�w�b���R���L�>�Cϭx�@�a*>�V��U�V����8P����DsmLc-z��u�S��S���O�`�,uBw���Z��3z���HEF~�r%�vKbv��P��Wa��z�y�X�uܭ7X�����u�ڃ*OGi��Ǐ�B뒻��W0C�v(P+�+��i�u�m����N��aaoiZ�y�s)q�:�����[�7lwAteN�ge�1����s�j�����{�"���d�f��G�̛�p�i��ꀪ�����W*��Z�cU�a�������i8w/��A}���s���.�����WTp�;B�P��;��x��̂��lН߻�;²���մ��a�HNP�d-�a���$N���?4U�Y�����I"�#:1�����B��w>X�S�ס�|g�uBx�Q��	C�����P5�<�=f�(��u����K[`���{v(_JO��=-=��oEz{DSsP����	�3z��Ò��`wV�<`,�D��$�5���A��l=���w��{ަg�-�jQ��kIu z�q/z�ҭ�vp�@��]5��"��o'=�^���f�ޒÒ�hFL8��P�{nk[j�[����S�/�z�	��N5�->���I}΍i9*f�fn���b�)/uvk_q�k���+a����C:m*��t�A�Z��~^��������^}@�����ag�2��uռ�܆�!�J�%�$g�PތǶ�x/��f �\����ޝ{|�f������}�����sQeX�ş������M�����UO\+��_wX÷~Wb�I!��1ە_4� �aX�ְǼ�R}Ư'QWL}�D��MڇLUS��cIvAR���N+E�k	�㵳��Ck�k\OpI`��������1|��g��7:�� �R1,���YJ�'�{l�ΞE=�Ǥ�p�y��J�Ovk��f�0��$"�W=��'P�8ˉ���ʊ4���Cne��l\:�s���u4r&�.>�n5����0�2��`p��q#��$�b�V�������_�
�&�Tn������o�|�Ã�������O=_)v�r�<z�������TgkX�o�W�ܡ�;5d��4;f�Ot���
5����xe�^�4ݜ�L��"�v,��D��Y1���j<����z>�_�X�cɤ^;(���6ܠk�ƽ2']o���{����f;�GB���k�R���O�Q�5R2�Ż�F;!�����k)���<����y�Q�k��M�-uŐh�41�Yc��.�UA�4�ܲ���h�
�)���7Ze���G��:點��_*Y�S�~e�L)���b�NY^�"�pu��(v��P�^ g�va��![���Vm��� ��v��	�nc�0�*È��LLm1a#*�mẴS���)�W�8�[�8$A͠ԭ�g�(m�EM�g:�	xm��s6����w��i��Ȣ��Ч���"��O�aOU�ޘϐG�b�'���3�=R�E��z�*μ��m�%�-f�<���g���s{���ex˃<C�
�Į+	�y6���k8��Haӵ�ϡ�V���0���7S� �\�2�2�YIdUL��Y[|�Z�;��Q��Ӝ<l7~d��;q�n�z�n�w�6���ml�ӫ�,��%L���ʬh����ƻr�{���9Q(��O�'�U�au�^��T���Hm�:V̩S��`��5K5��m.&�fn<�R4��8�8��p������zl��n���K_\4 �����g	��8I\�S��i��V"�%-/�iY�ظ�1Z�4�Ʉ,�ڽ��{uV,U����zo<��S�w%�ν�Dv��m��R�g��]���e�9i݅��S��+z&�r�Nr��2�C�@��Ʀh䷌����<��ch��=[�B���ݬ.tޘ2n`ãa�Q��e�c{��
Ơ��Y�4I�z2�h�ٙ,��	�uv\�����ޠ�M49j�\���#c���]37��ʯ9X�/��-L�i}������'�,�(,�JZ}���I�4E׎�.sNڜ y������_8��s��y��:�֍���iC)������T��N��ʱo6m�9fEڝ��_]�f�3��NҤ�а�q,�J��r�RFS���=_-��n�n���Q��0�e�Y�prf�3\͇i(/V���a��OA�ժ(��f��Q!܉�t�-��lQN�3T����WY|!ʆ�d�i=���X�Ӑ)�1Q'a��9�R�P��1����k��s/4�yf�p�Ty�s�:Y�4:
=��V@fީ�����݃Z�y�';T\qm5���Q�Cwf&,LT�,>J[2ܤ'V����fë�:���j�%q�v�V;�;���w�m��,`o'3J]5�q��۔אc)]�-�P��N�:�*�҆f]�tb�ה�=_M��rѹ/$���r���z1�Uza�5�m�s�]S���Cn�!ۋ�������#�:(E�9�E}�嬘 w�&�]K���j�����e;�s��8ܧc�qB��Ww}��K�؛8ۼ��� 7b|�<]�7��f���.u|���Nn^���2�R�}����z�4�ܜ���[��<=�UlKR�,Kh�d�s)����w�k���P�W�A����]4N
\�����ru��j]��h��)ّ������b�I�OX�딃��aH�z�M��v�I�Y��6pLags��o�^|Q;OgEZ����O_�.4_*�F��T>��U�=�z��ˤ¬-���V���sӿR�٭��� �☦jyX�ٳq{�WR�3EPx��h���"��F�x�|�_O�����~?����~?_���,��TR�cF�EAAG ���E4�L��>�z���~?������~�O�/�m�9�("J�F�9����H�(���J>�bZ�JH��
b�*k�� ̥D�$�IMU��(fb
�ր���C�=@�#�cz��A][Q44-U4�Dyؤ�����d��Z��DT�Q^a�PPU��E�AQR�CI��H�����u[JgM���C���L�U1-l*���<��(=��%D�{j�l��LD"L!A�M8�!"aIT�xs ݡ�9-�t����/N8�{�v�r����0���ˢ�X����ޛ-��8��/I��G� I��5���,FK�B��$��n)��m��fD�Q�D���rd!����?���+�}����������n�^�=�#x�jg�D��A�4{�4�&z�=5�63gח�$��k2�vվe�Q5�xd�f�Ƨ�0AY%���U�?�s��b�%l!��["�5s����
��h[�+����G �椲Hj�*�hg����,���I1c�X?|���l��ox����r�_�/D܎�QX˝'���('Z�.��ru��.b�θfOT�MA�Ĳ��8�#	�vgd7��8B9�B��欘<��2B0�׭*�*��\�)���V��;q*gj��Q�ݕ��ν�5����	;M�/�ԛ��!2OaDO9��m�D�)��U�-�v���&�v=4vt�z$=���2��f��{�Х2�QM!�Mچ�����Ʉ5n��x�l8�|��\h6��&�231�>}�懇,�C���|~������<7;)���K�G*?�yc�P瀛h���;0m{p�Ѓ��"�.y0�;m�����o.b�u
Xe0�9+�Z�\��9bW����kA��l��#�s>:-/�697����.Ѩ/..�X{�p�}sk�g_�(�F����Jw<�O�h����������}_4���j�r�܂ud.^�E<�{�C��|%��t��۶��Fg�M��Í&��ϷY?�76��q�}��}_W�L3��	c��̵��^y��w�qd�,)lkt�U�[kg=8y쮍����ƶfb�փ����,���S^��̜qD��{	A/mbTs
(�BM=6�`x\�iT�u͉�p��c!���}�c&S��h�)��y��sY\�6rR	�k�@��J����P�B���P�_�Ɓ^��0���,��#'�l�Yy�EfdC��:�owyc7bu�(f�z��P��h�c>��l���ހ@������{a]ZML�@]�sn���]���n˰W�m� �z�!�1l*:5:L��#�|<����l}����_��=0��n�Q��Uo��"��@%�Dϛ}q����8��#���;}�}��B����ܮV%?�z�uC�5{9H\�0��,��RuÖ��ƒ^�ki�Q;Cx|6b����@��aAg`��k�%�U,7��ټ�&X��3Ц1EQ���r[_�3u�C�v�sվz���{gh�L!��"|��C_|��p����~q��;d:؈����W��Z�늲�.W���S�m�z�)
�yGwwC'u�bYz�+{�%A�����C
���rWM�Lջ2���B����tڲM��I�5C��V�B��xo�r�������}�z���y���罦��/������O��`X�����{��t��{w���2!�$�F��A���r{��g� B�5�bu�bi�|��EL~�8T��]���*�3w/��_K�$51���K*ar�K�e"�H3})�@�.�r�E��L�P��N[C�m{�y6�t�k*�U,�Z��a�BKq-��"M��p��o*0�=7���~nCT�.%�G�}�Y�I�;�:�fc��*�|�~al!������g�Y�(Y*L��X�wƨc���a���YZ9�wu�^94���������/�uG}ShQ�wJ"�$��~]87j����tv{��PD3e�[�6
����(������Q�~���p��kx���F��gPTx��`#?����|g��3��@5�P��'�x0s4p��&rx&�:���L��lǙv�߆zv^Ͼ]`���>��o:�htx�Xh�I{�s�|Y��Z�M��)o���B� ��f��W�hOAx�B�'A!�@2I�i�[��s-���f��v�VѶ�Fb�9�YAe�J��h�L�����U�{��'\�����QA�F�۩ٹt4ũFC����3;���J�S��V.��;0#!��Q�q��[r�e�MQw�J}5��
'�g.��B�e�����u��g5�ྠ+� |�{\����A�z���4@��.9���z��z63k�y}L�[�Xu%��ML&�S�~W�h�����>��ե�f�BQ��Z����{�Nc�T�y�װ4�J�����Iޅ��[+�����v�C=lSd	;A�fͧ�{g]]�Xq��'��%���ʙ����|,�������?=�wOG/UX��#(2jY^�2�z����9��������cF!`^�%	���ӑ�N��^d�@d�殈!8E�~)�V�P�
6��w�,�bo8�uM�4��?�:_�Y�ٱ	�a�/D�&�O=y�$��)͂�S �2���r!�c�:�b��N�~�Wϑ�ۊ!� @��$(� ܳO��1��fqzL��M]$�b�TA�ת�Q������7T0,�r,�>G�^�P!�9�k�c�f�D��|��{ ���A�崎�Ml�7<�b�]����#���}��;�]?���韚��#xe�Bw����Qq0a=L]&X��rO7�۷���I�V`&0��w=y>;���,c�����ܑ���6<}�|c�{k��r�Υ�lZ����ͥt٨5 ΢=NK"B�r4�ul�KZe=�o(k�2\��z�6$M��i+=�ǭ�G^x���(��n��*;s�بہqNԘ:�i�)V�ʧVzN�<�C�.f��tf��r���K��W�>�ѤFj^��_�_-j�V�7t,���z���ܔk��=�k��/*��T���wf���<��X:�[��|���[]�Q���t!�]cԾ�H���2Xqg�V��=4#��}�����^nu[rE�̂o��p�2�ScH��%�]��ޚ^Δ��.�`�{�vh�ZH��:��5����z��l��;���-�vю�S�8L��mא3��%�GPZn;�k�'COn�.����7��~��T9Y^�`�|G�6D�OP�֜�Ǣ�W)w#.��\��b�g�إ�B&a�ƴ���y7���	�"�C�[��uF�h���7�G�fN4��$8�p�!���@!��F�O�f�P0-�<����XP*'a�c��C��Ӆ��y�D܂���\V��A�&�:�z��\ކ��euDOv\u���Ӊ�q�c��,��Q��,�"��&M g�Gol,���-��]���d���ʌ+t����+V��g\6�F芪hͦ�ړy���Ht�4�������v�ʹw��Ƴ*�6���ڻ'���`�3sb--dk+:+�F�_���L��Uͪ�9���+�%��Tg7Y�Ӗ86�$5"��]x3U��=�BJ]JJ�1Ǽ��"R�;|�������ޏ�1�/�#4>�N�W�+'r���-�H\�P+G��W�o(͵�PK�3�7{��w�&J�-����e�F@t�}m��(�3������7i��\W�A�J�J�z�b-�v{�@63
� V�cYA�"n�\�F���'�����Tqtu,����RW�Ψg�l�3M���MJ�;l�]�<4��d��ASS�	�0��r�mw�[��m��N&z���[w('']��8�f<5�x�pwd^�)14��'�W���Pr6�kc�p���6���m��ohL�������7ܴg$UĿH��
"���h�޽�^��{^J:|�4l1"G�����)i�a�l���v�a�qa��<0t7U^�)2	|{ў|�i�;j����g�5Nf�H�c#�qY��yo�B�"I/�T]������G5�	�L�ϳt�X���l��Z��]�Bۓ��������X�<�z��.� 0]N��L����a\�ED�³p��RF+����� �:�1��ŞP�u`�[�)�R�f���3N��+�7���;T������������[�B�\3a�K�ܬ�>�^#��y*# =ɤ^R���%�M���՘�!��p�C����Q1��ȹZ��("�P,�Y�D{jj�o	��G�^}����yDA�G�Y�ҷ����+���tzo'�^�c�U�n��}����^m��
�s5l�@׮B��H��D�޶:�m]����]0/v[u�Ɵ�O����RPT��h�e4�:�"��'��sQ/�7{����eXV�����#F��*�k���n{�n��3�eW\�qq�C�-�:t��4{#I�4{�	y��u��쟍	��[��y��b{P��z��#V��-SA��zN�(�����n�ŉ�4�Fc�l�%L$�
�����Q��^�YU�J1p�c:��l������t��Z^<�g���a#z!�������O���h��|�Cx~��v,�g1еQ+A��)���v�D���Q�S a
�Z���X�[uo��ܽ�]������0BB!�91g�<=j߮o��*�����c\��\�&k*�*D{,�Q5����\����6����hu79��}WW��h&���}@|=$��쥾mΟ{��;@�jh	N:`\�'�>`�qXo���R���LG��O��{<퍓7'�랹Kڇ��z��L&
v�%2�;�bp?���H�*��w��u�,��{��^��H`rܟA�M�m�ף+���4س���cზ���'�%����4"$i�9$����v3E�j��(�]o�K�Ht�)�@�g�A�3��o����tDNj\�������9�x�mi͜���s�6�7
a�z�D�{�lD����Ɋ��4.V>>�v=[�;A���F�7�z��r���	x�j �� �r�|�E"�Z�z��=�æ;�Ʉ���.#���K�$�s>��~����sĭ;��]|�B�>bE���� Uɔh�*��95~�n�:E,3�7��ow������*c����/����y��r��*��jh���@o�Eݺ]B]��H�6)�{[-��Z�z%涯'����^�doGsNh�h�ǝ*��2"��^�;f�+�;Y���.elع����1ȗ�m�P�hl�����.��F�6i��R��R9;�C\O\ܜNY?UW޺����Eˎ��]���=�3oUY-���`3��[��'�s�P��	ъCns���q��{8������ssz�ÉW��#1�m�[w�]��:+�Wsh}��Yk�<q���y���19���)E*|;��0���l��el�>�)��a�k��[tF��2:�E#�t�ǂ�-�f�vk;�ִ�g_�h��C;C0��~�J�s�U�T�[�(���a���W��y�u���]'E%�L8EH���T���Q}Yɰ�:�`������U
�uCY܎P���}G+<�ϛ|�;��#^Ei���y��e�A���!�n֗w�ٻ�I�4h2���=h�~�}~Ҙ-}m���B/��'��x��T���G���/x�:(�Sv@�ྀ𔇚F^�ȟS����gh6�rxk�V�O��Is��9e���΋�!D�F�E�h�x�E�ǲPݲ)��gr�����nWͅV�
�u����[o���)���Xq�N��W�EĘC��y~�?�ө�������i,�I���̸#�{;��zUR�LD�gCwxE���ۦZ�ݑ�r�����\�G�?��_W�|ǫZ�0����B&�_\�"+��䬉�]�r�ڭ���M�LE�WN���V�Db66|G�z�O�@ɋ�ܖ�� ɵ&�GZA�Z"���D��q�b��f93�m�~<���b ���+q�G�x�4L�nfy��&D�ln��ov�]��=N�궿pU (7>��[�=Z�m���d���~�/f����U���-���:#��8�=ҟn[����$��x����PS�Ƹ}��s�v��gL�^�]"��L������Ns-2.	8��yyx��ʲc���p�4q�Ro�o\�@.��ƽ� �Qn�f�Hh�dw��UJ��g��6� ����
�=B�*�])R%wp;Γ��vTM�*.r.kgg.��k��p®v�D ���f�]P˕Z�1BV�򱰱�T�E��$�ѧrp�r��0��]޹|SziS�rj��'�]r���O=S3��1�]�uՒ���(SP2�F��+��c�KN�3�r�j��]�&�U�oV�D�b̶�\j䕻`�|wj���1��tUK�N?�����h���`�ujn}k���e3!ӹ9�V`}���sV�ĦjQP�� ��9��Ю�;ӗ������7�
�C��+��f���ݼ�t�	���|�	7s�L��I�m'c�Bs���K��z^��q�Bs�B(���Wz�t͜]�N���h�Y�Vզf'bwW�nC.62��XQ�L���	�������}uE�GuPΗ;e<��@���VQѣ�07٠[���]�l���^d��hC�5��\�v������oP5�;��G�$�`+䯙����P廨ý��Z�a���|�g>���0�+�[�¡=��l���l�6�3��u�eք��8�ȉ\�X���G��.(q�Hd�LT���g�x2��]����1�z���	Ax���\�(v��N��w'�M�y(c�[��A�Ynn�F��2�V�|%S���J��BgR:#������(3ē���ͣy��~T�����	�����+㧱@'XTgSU��U�ko,iÏz*��o�����&��l�ш��W���̉:�K�w_`�U8�Vܽ81v���p�#Xm���]0��`��u��\4��ˠ/%��޼����څ�MC���՛%IN�ud����z��S[�3��l���v�X��5�򠤼uJ����.û�%�*��0�����Ư�,l����}��Z��U�L��cszVXÏ1v�P�RjG{��(vQkqh�yfqq�3,!�{�B�_y��	�:(v�ޘ���;�30�gv��X�}�2ž�u38�{ orCQĤT2����n]�u٥�
q�l���� ᕓ��h�e�i]�=���s�ά�ZT }jY���{7�C��A�S��N²,�{�w9�Y�bs��7@5���a��Yټv=E��i��.�N,��{z�ӶP��0�ڨ����)��u�ݾP햞T1��>!/��S�����I�uvi�ʮ�IWF��ˏ�t�T$K7.�kH��o�=�#�ImTR�n��*�(����|�3^��$���5v\C�<�v�
0hw8��I3�m9.J�s*�`�i�s}Wa�A�d�<�z��<:�Ls���ԫr�w?��u�UNE���˘�^mh��AdAx�1��+�t�R�@�r� <�<�8{km�
�opmu��Ѯ֥wpuh3e�r���m��-��㙑�
µl�V�^"Yw�jA]���Ν�փ�N����- �C��=�q_v�uh�_g%W<�K�E�ٽ(���\aix��4�sL���]R�,��wAT%m�D&C���V��t�r��l.���W�n������L���U�F�'�#��hih
B��&��C������z�z�~?��������~�٪)��Z���(i����<* �(�������ׯ�����~�������gګI�i��ր���銝
(h�K�U����Ųhh����vն
1�LZu[j�zt���F%�����E:4���i����nf�l�kI��A�N\��cN >�N}�/8<*5��B6�I�|�rLS��:K�Ѧ�����Q)H6��ؤ�+�<������\�'���i��hxܹiѤ����Ѧ-&�6â���f�x|g�hq�1�����]�si*�	�Е���F�76&�\���z��G�^��|��ڠ�s�����|�	V/�s�<u��9Ǿ�U�z���Ԧ���˚��o�^�Fʤ1v����}_P z�vp<�ts_0����l�g��G�G3��o8q���]����s�IK�{�tj��A~���f��1{Ϲڬ�6ǈa���F�_ �29=*}�7�j�����1!�6�=ZJ�2gķ��}�#�ON�s#��������2N^^+g�D��.�/�EY�������y�`IsbXg�}?�Ȭ�//r�{Ӭ:��Q#�Hȍ�^_ooz����Y�h�=��Z̧�����^믬�Eۑw��|��*J�ɨ���^FJ�S{�
���qc���S��*UM�<�tJ��G�N��]
�X��:B�J�b-օ����n����ߺ��i�D�[)��O��ȩ�5>�� r�˞!�Gl �Qы^����_N�K�2`����vj��ǼSҒ���\�i�M3���mjpKp�=��݊9�S�=ÄV�>ޔ���k�+�k�5Ө��C����0_�����\��t�R��
���кn�mMaU3��[v��������p\�?mua�n�`��Di���)Ù8���b?K�6��huV˫����sE�p�X��HiaF�*nQ۠ ^{/��^y��{�n�ƙ�H^�Ol����� ���17�yp���Wt�W���r[ʑW��*E�ѣ��i�kWu?�;��jN�bH�[ ^������Ҽ��t�lM���q�ߓu�Uy=l��*�'��N�l���5��a����7�<M�F���GuL��5ٯ$��6���1���!�q�8;��A�0���<�"��5âx�eJ)-k H������)>���Go�b����ֲ�ם4A�|��.&҇�v��ܷ|9�]S�ǣǤG4���h-޽�}��p/��H���{����"���p۝����=�af��+�׵���9P@�xVh��T/�o�q"G7%�-w�U;����s�{mϺ�-o<���!�
�~I<�k������Pk�1�q�g6N�V��p�	/���lS��g���T��>b�����}���<鼓E4C %�m��_i�O`�T��	�4)<��K(��\4�X�h��twPs���Y}M ��m1p���7y7;��(�67���^�Olu!�M���v�h�=��	{G��["&��9:�s��Ow��ߏ��}_ 4�������W�{{��K�����K�cܤ���4�{�\��y�Q�����!��U�N%*nI7��7�W1��ů���Ad���ג.i��y�_kwUYeq}x���"���F��ڦ�l�k�U#(�)JP`��W]%��ce5w�v��7�����T>u211%z8E���#C�WK)�	h���y�㽼�����mw�7�������BC�Q:-N�<zL���s6jg�dV����e��k{�q���]@����۠�Ð�Dp��m�u�LU&�v�l�ټ�7ns���4�Z}��_;.S���\��MF�l��R�t5|�U�u�of�{&�Ǝ��"���IwJ�x�e���������ɟ���w �MQ��������Nݐ��Z�1AVǍVN�{����x������pF�F}u�Vy��P/�+ܻ�~�4�&MAP�F^{7o[Q�5w֖M�k"ɶ�`y�[FJ�U�*�p#*��+����-Q9���ϳrS[u,Xoy
�[����QG�ں���R}�[���\�%��Aj_90��7���Z(*���:�&TX����L�z���{O����0;3��~��_��>��n�s|:`�@^�?�\݈�����z�.�;)�fl��)d-��^Q�i룚�3�����^t�7�4`e\������9�'��39�Ρ^�뎵Hՠq/ �#�L`c����ђ�Q�pD�u�_i�P//�@�<#s���{��ϴ5��%�Ov�N�M����hD����Ǹ���#$$�Ex�
�1[���n�����xWО��^^��ߞ�q\���#9-��	���w�L���4��)���N��HD��~mS�i� �,Bf�-�]<�,�Q�v����yr� ��x�W�i���x�l���NM3�A�Pn}	�o
չyM�u78%\sft����wV�z[�$���w�˭�u�{"�$-�R�]Ê��8����y���<y����*��W^�{]������>��~���5�l����U7p�m�����zW����]ޭ�ݮ�����D/�ީ[�Fko$�ti����@a�s�њ5=�y�D�y���ng9Kq����]ZҊ�����ݛ�eA����G�+���;t�ԕ
hT��gH�9O����� ϼ����&�T���j�VSu�X��K�N��-��O�ae��"��L�wv�������mˡ�0z��I�*Ϯ���T�]�w�G
Ʋ�^w?P
]���C�F_�xP��-�*c��=u]ˤ+]��E�\D�ɹj�}��/t6���^6��,m�~�v	t��S�aziPrn��A����P�5=�|� ;����ԮWG�H�M�7���b7��8T�\ИX�En&׎�9�r3�Pe�k����M Xc�.�r����v���]>�ɡYY'�;��mqXJ�'�Ď�b;��s���5��UDe�fP�wۢ�t�r8f�x�T"�*�m��}��%���I�<������|=�F�m�ը�P������'ٹ�7cׄ���u�'V�tg����ϲ��������;.�o����Q1�+.�����Ϋy��0�xd/�̬,�ɽ���ɐ:�7���b+MM0��O�%��-1Uj63*�w	��3��a���_w���|G�N�e�O����'_^+r��0J��K�l�x{#-1kv��p^�X��^.�òU�u��j��0�/��y����7�U���3�{�mW%�s#e�!OA���[��oTa�Q����;����ѹ�$B�+<��OU�M,�7���>�mF��$����,������bE���!N���`�J����*��u���Kۡ�ԴA���|�6�;�mzO�͐�W�
]���b��<U>�y��b��ȕ��\i���y����[^��w�Y�ݎK��(yJi�M��[��7/x6J���"�����dܼ�HHp�����ރ�M�<����so]�fI��n�;u��Fs��m�K�
3�7J3:�+�0�,��p��?�
rp���)�(sb�[�n-�����H����vA��XWc:�o0[�;8<l]!X�m�'_�9�8�U�V�D�Е����w|GHͶ���5�[3��@�!�O�T$nG����>+ң7�A��)��ΰyׯ�]�y#�p����6եY����7W�2�ɀ:Sf���y/k�����.�¥U��\!�F����DYef�@��Br��7�$ƻ��CG��*��n�h�&�g���6r��:�y|��R(��{5ͳYVҼ�j,��R��������9�$t�ك�f��I����L�-��w~2�g�w�1���O������xzZ��O��㗐]W�9Su�� �A�����`&��J�/o�{����/��ǋ=߅g��O��؍����˛�?�� �WP~ITUɯz�޻b��|SGwD���/5u~�+���]-ys~�g���j�rbl�5��r�t�J%�*�B\�6I�h���ͥ�L����]�SWK��V&pb�6 k��3�6Uz�2W�y\t��U�ח����^����f���Q��B�{M���H�%(\��y�s"�u��."4�୳���ʠ-�p�������|����8h��2צ��{�s5CV�P}��S�/��_�)���s���2~�~�WƔ�}?��7��#�����g����m�6�.׈[QÏ���wq�����C۔�Xۢ�6�̘A[���Sd,�춄ٛ��kv,v8�5�A�#gwc̫>�)ª���6��ĵNS6�e'���a�x�V�D���"�Gf<�.g���a�&a 3]�F�!:	Pp׽.�'ڪ:�!��A䋬���B<��oA���x��o 2�G��SAJ�@�@9��咧��Ah���GXf�鑚f36���uF�H�b	�=&���[E#�{��k������{�:e�f�vE�qj�|���Ha�s�Da}S���T;��Kw����/9ŧ.D�3�䡽]���F�y�sH� �q��6���Ҡ�ǨՔ9wP��~�[W2ګE�Z�͐ꐤm�|������eh2�.�ə���lm���ky�d�ޤ�8���g���;���'꺄rJ���i�w,쫭��ȹ�;�)�80`��f�����%�	;,NC ^F��F���w�V�h�h�����5j</#׳[�'�I:�Mɱ�oӢ�)l���R��z';�����щ>g*������;T��#�%d�*�ss7;^K��p�fNv6��N�c�f�(z�ꉳ�W��m_g�ԓ�� B��z�P�{i����9V�J�}6!2Mam���ŧp;����t����3#��?5nV�� [���ҧ����m���}§̘y�t6UwdG��MH�;k9	of�Y/8��'k�X�LcV`��il���Rq�Q]S0�W�~���eޓ���t�s�6[/F\TK��g�=b	󹥸}�C%w1
��kVZIsqٻ'�{;]<��y�OsL����������M;88;��D��s]=˰��.RE���ґ�oݙ�-$,��+�sWW7LP����9�4V͎&�:EX� �3�'EK��a���!B�����%�F~���4/�"(N�_����h�\��/%�xR1/'���"�C�F19}��o�2�����]!�u�\g�_%TqtM*F�]�F���l7d�\���c�@��A�8`rV�z ��ȳ�~����j�.��kW\C��{�W�ÎL_n�T¤���`��`�f�vt�;锘L�˹n̥�-9ۺ��Ug��t�%t�6z��o��9��l��b�E����h7��\|jүg$B������hѰ�=����'�ܾ�13wߕbO�[�:�&\�¬�Q��:��*��˯dɗ���~aE���0�i�����r�.fmž��ձ���OHѪ�wp��U�VեYw�3O��M�����;����
гM��B�\�ũ�������':���y��h�4\a`QA���U��g#\dω�/��OH�nz��Q}���65��U��|'���~Y��R����<%�C�e�C�w�g�G-Ҟ|l�vp���a/��� ��>B��⋎���&��^��w�mh}k��Ln�c�3gm�^��#��6�u �]��D�H˺�,��A�ns�\wr3]�f�Ҽx�*��]�y+.i��W��Tz�0�8a�Slq��նv�_��7q#K��Z�S�:��u�z����V�����D6mU����X�l�s����M���-N�G�%SdՍ�B�ӭ���w:g7{���.�\2`��V���)+�xGv��)��2��-�1E�*�w��S��m@~Kjx(�*�׻<��U��6�_f�b"�i�[z�擏����@6�S����ճ{�j�l���&~����G�FQ�N���nm�8٘��g�n�����g$"c��Ә�r�Y̗����2��{�D��XV�n��^Ӫ`���������9�p��u�cPE�G���D�htq��Y�n.�Í���:\,ޔeL���p�[_�����q_Gq�{���l<���µvu�{z�/�]XLo^L��ԣ�S�fB�j���a�A�k��"�����i�}����+d.󍽛M�h�/b��i�/�=R��7C���^ؐ�Q��+F]�"�gi�]3�#)*S��3�Ej����������+�ϫ���/(7�l�Ztr^�}�(h��l�V�2V�z��\YgJ�v���v��{V�P�N�ɢ�+�'J�M�"����ueǊ����{�pt�}#*�F ��e����:�l����z6앉���[��9�˧"��}�rm�'�Ǝ��ہV.�q�����m4sȶiʗnVe>�+�����&�D�c�*��Cۨ1(훱h���ڝ8xz�6�Lb�8�	[��{^Vm�]��1fMA��;��젨�,f��M���2�MD,'2�
��ݝ��u���[nc��7p�͘iɃF;�@�.���t������ET�rXN����v�c�ro!dg&%廫���fI�-�$�L�/z����Ө8`e�uY�p"�qlv��p���z'��>i�Em�F*��6|�<��n�l<y��7��T�����+^5�M?����^j7E*���ߪ`�;�'Ϸ�8a������xY�a����N��㭨IAT1�Տ�{��u�(��i��H2�Kƛ�r�̩M���6-�G��f@�W-k=�ݳ+�Y&[�����`q�&hy�bר_Nt ��v�.$��UR�b�7�7i>|��y��s�K�.���R�m!rɇz�ӗᓟ��s�l�svEz��+`��4���{�5���9a��]M�\�M�۲Y}��52FƘ_t�΋{��ЍRb� ��5r�̈́�b�k"�;-ޮ�"^my��gX�$̮�nh�8�C.��3]�����H%��w)���Ԇn��ʔۓ-���'s%�E�c	�HJ'`��gz����U=��b�r���Dج
��Υ��Un�b`���S;pPk��cfe��"H�QP[�]m��Q�(d��V�IX3���L��N5(g:�yry��etE��ͬ��e�������9�.��r�5�&�I�o^ov*o�ܶ���枺� C=mj��R�k�����VE�2}��J���E��IæT���Ҭ�s L(-��%�b��7����s��:5y���r�X��|�ْ�>s�u�qm�'=tէ�lR�kq�]��#b\�4:�p��Ԭ��l _t�$lK�����*3O���6
h���A���<�ן��ʃ��[ZӠ�Q;Q�5T��^We�bNs'Z�F��&�~>�/��_o�����O���?����Q1�`�ƍG�s��3v��SR��A͢hv�1�'�	g����}=}��o�����z�~�~�E�ö>�.Ti5Wq�"y-4���X�Q45c:R�b���lD�m-%'$��4�htj��S�l8�+@i�5���jZ�6����Nو��*"CN�SF��E�΢�-��4W(����
h��KMcDX�mI�b��7�4�Kȡ�ӭ%�Q����i�h�J-1��Z*�l[`<!�W
4j�Z(-&����)�֨u�m�kc6���e5IN*m͚|��#kPg84Ph�)j�[8ڏ�sh��u����Q����#E���+�5��N���jTkLkTC�m;h�Z]��Fا�]���5r�Q�p��m8K���0d����N�j�3̺Th(�>=�*�?=�D�Uy��
&�,5\���D]�3uPfj�0є��&nҵE������H�($b1�
0�Q��4\�4H�8ag��6�x�[��n[x<r>?Y����õ.��bd�K�[|���G�I�3kgG����:�t������w�S�����Ș��;�2y��n�E��U��)g<���k����o@a�����f!�z}}P��
�"��o�J�q[޴�������I�w��S1�ݷ7�^��㢎�2�uH���4h?-��X4����vO��b�3Z^.cr�v�m�VV8l���8A}� @W��H�^�^��`�4�u����f�[C�ȉ5ݛ���FM}v#��B0*��"�s�3�L��BR�rW�K6�Z���~����� �W7&�\&�J�/p���k]�?lXl{�k�M�������{�W�N��qc��E�5�{{�=�n��N��k��P�r�(O����5⎴��St�6Y饰_:轫��X�f@{�1k�\�H<B�E!\w���;ݬ̮2�L�z����<�Q)O>ڏ�����˛[��k}�W��uu�BY|�Δ�ѻ���4�Mw��0��d	�C����R.f������y�:�m��!T%��Ě]XNճd��G`�Қ]��a͝��i�y�v�h�/7�xk�i��we����u�{�\7˵Mí}t
��k�)Q��+;u<me�m���>뫝V�"��)	�H�T�z8G��KjE��ӓ�z����7�z���p�p=�g5V�I*m�t�F������j6dQ���z�8]�0��UR[ݶ�41�����=f[-�m�A�!kF�F6��,��3w�����uGH�-�9R�a=��l�H������QJ�U���l�ޡ�_AS�}���oZؐ(�b��]�Y�^odn�x�\3s9uv0�l$BP�!��y1R#���IR��2����aڮ8Eҽ֝����Yl��#6އ	���n��_Vd�Q��X�Qy�u��kв<��{�FO��l�o� �<��Ѐ�����٘2�؈��y�{��e�eP*���^��A� �>���o����=��o^�S����j�f�=;��d�k���鲫u�\�(:�m_^��	�^yY�fO�?�޸O{�ڶ��˕��hw�,�\�Z�$Kbd����i5ú4]I2q3�q˘��v	�)���y�_n�'h��1�g_tηvyy��v�ic����8I���qH펟w28�ϧ�E��g;�{a��'ڝz��^/��*��Nn�	DIDA�x喹��s5���g˘;�6�vh�*�&� �}�"j�2�GW��Jȟ�x@�z�Q=[lz_�%��,~�*Y�'�� �S�Bj�V�\��n������C\K�~��U6#I�����~��T6����'�g�+�b ��Z5���<˫&�)ۚ����w={�4���&��Tz�^%����	�s)q�55}Y��|Z���9]�]$���+<�5U�S�n�ݙ,hY��z�U<�W�ɢ�B1\�
��Q�9�*�<�+���j�57�t[Q�s��������.��;����S�:=]�h_��%R�\lk�&�[z�f�3Ҫl-�������!s��\g���*���iWރe/�ꫲ[�Z�9R<���	Ѕ����2�h�,,�v=�g����6��}L�ڋLI���7�r��3���x���a5�(�Έxd��]/zu-��D���^��GZ�L���Nj�U[3����h�.�A#���w��k���y��{��swn�-��g�cd73�`?.4"O���Y�X��OU�v�л���\�n�$��(J��9��p;>�a����#�?���T(���\�:�k��m���ߟ{�{�B���~q��� �4���������7�˛�e�!���F�����.����%/,����^�{/3	s�B>>�e��yE�}�mp�G�x���G\���1���2�s	���)�W�8B�:��H�6U��v�D�#���w6�u6�����m�̋L��y0����^�M��>�Ą40�fW�v8|�K�u%vtmn-C�I?VL�q`֛�]߫��$~D�
%�"�hg��u�;Q��"���H2����c^Jɶ�v���q	L�=�gV����g�iB�7�&#9�REb�AOd�m\)_�^��֝r/����)���у^�Z�/'�ú��綠��M�z�kJ�H�<d��}�fe\9t��e]����PE�p����E��d�Cb���1�oEf1��IDSZ�V�4�hû��m�\��yڳ��eb6osVNsڒN�7]�����o Kn��{���l��權��ܼ���/V.&�`g!jL�!݉�=<�)T.�Ĥޯ)0 V�W�]M4D�ӕ'�Y����kH̄���^*��4����b�1ㄽ�k�9gwp5�����{��ϖ�#Y��tV��Q\z��n�%4��D�RF�t�Rm��ӻ�xq�g�۲;k��l�An'ѫoz*~�:��Y�4Uګ��ss��yh�(�5&��m�W@`���g���"i��m��{�w]l��onsբ��eQ(ĊY� ��k��0n2�C.c�Z�����f��LI���/��v{�q[E5/�NL^H	�n��%5��Q�_���A=~89��viN2�;E'~[<��J������}���
/r�:�7LY�!%��Dpߏ�����am�1��X_$^����U�lC��S�2�����v��[R�V�r����t�
�x����6��o�^~��TY�|����)8�{��E���q�G�^�l0�#n�[[s��^���=ҖE�=�6z��:��4��k�<ߤ)ww���h�=�v�e�"�ÔY��F�gb�K���Id��*{�n
��Bn�ֶ�z)sA5�>��}@G5�d����^n��I�x�<{�Q��~����
��*���H�ջ�8����r�Ӓ}��k�+A�*���f����+U�����Ս�y�ɔ*{�[ƢT�܀��\���5⎴�ҹd��z�tӆ閫�̘����+��`L�d׌᝹�]d-�PR�:x�-�����x]֝�{�ɧɠ�uEW0xB��,���-AGK�s����/ۗ���pw*�j�2*�Lf�7��}�
���Ɗ�9n��W��q:� �����TQU^s�-��x
ؠ|�*�]ܞn�]�Wnx�t���,0�<
�J�:�Z��㫨�-���~!�� �ɥ�Y{�0��TF�����Ө�\�rM�k��J�s����%^*��[\���/���]�幓GOٓ���$��˱��-�JUq��뉍���i�Ϝ��o�_/_s�-g���y�կ�yӵ�qjKşb'!�UI��H�h���2��ƿfؗ���k׺B�~�	�gv�Z�4�ޗנ���sx���
)��t(GG�
\/�E5k�j%�u�=�U�%<��;o����ȍ�g|��y��K�q~s�5����}C�:���Mu��]Wwy*��1�\r�7{��7�6��j���[��4��#{|�(�m����<zND9v��ʡxܬ�[��g�od��A�}���?b5f	�~.C�[�
;H�7{��ɟ�d1�Q�A�t3��6�]1'*�gf�L_{���6Va�uVkm�84�O�����E�S��ͳ�_[YT�s	���8��~���a��RR/:�����"3ǹ�Yi�:�n
��4Kg*�ȇ���M'{�hD��^dya#�v GJVD��̪�O�h�s,w�lmNN+~��{��a({���$[�/�A�}��ve�L�*)X;<j�Nk�nT�'A�TK���&�pA��V^���j����K�{i���tSߴ6W��g�@�*�ד��U�j��˺�z��:�����ܦס��I�:�y�	ݎ��:��ƈ�)G��R���4�ӆ�<;5��|�gEP�dXə��=y�E;:��}\���5�ol�\S.ԓ�8����f��G4ndn��0Iŝ�����76��}��s���~�����Y[^MO]c����a��E"Ώ��j��-�u���R�E�e����=�Ӓ��mhJ0��o
ތ�H�:EG��3��d��//v���3�\\��t~������x��eT����*��\lk�f�+6=���V��;ݻ�Ǯ{�A��W���t0G<,���S�F�W��l�VA�1�wnϯOI�u*����k�a�i�T�8�����T�T�8m����/	U�]�+�K��a����f�7�WAZ����!�&�^�;	}����Y��u�d��>��H��m�w�p���5R8n�>V�kޚx�;�]��Q7�P�(�.�*���&���7M6�5�WY|�]oQ5i��c�1���:�	E[\
�Mq� ��#�-f�4ō;���wm��5^8z>�o����0����wE�7{� �>�^���v�U�o>��/;q�0::��U�Y驓�7#�!Yى���w��@�<݋��l�߸<��8虧8�ݏ�a��Jo`L�P��	QB'Q�b)��Ϸn�-��;i�9�ɶK痒�D��޿_���W���۳��ͪN� $5WG?z��=�Hj���� �0B�y�)�>�����8�ų�ς�[>�5Α������$�&�^T~������"(�q�_�"���`v�bt�Btwm��*ˏ)e�B+�%vK��)4�}�:י�;�Ca�=�s�O�[�n�<c���ʽ���QH�0t앵r*i��~(U�'[�͎��^� �����״#ǰ����dj���pR�2U3K3
�sT��+6��w��=4��
��O��N������m.�m���}��4���s}�^O�>�N������J��z�(ųEC�մ8�ܱY���{7{�h�~�kw{k�O°H^಄j� �
�����_
X����N}��\eI_j�='y����z_�>�͇���v.�vh]�_�Vxά��Ѵ_A;�mt�Ƙ8�`�Pv�nf�����EX��j=�άr�g�b��.׭�KKw&-�۱v���6�Lݧoݙ}�i<�<��Y(��k��E�ْ�#� ��/[�.���yh�����i����(�Xȇ�خ�Xx;P� �ӻ5N����}_P��q
k�p��0��7�ߦ2F�m���Kh��76)9���B�&��m@�Fm�j:ȭ9�:��W�å�dxL����4���>+�*t����X��N�p{=�+u���e�H&C�Bi/�\B��޸1�8��|�e����ޭ�Kpm�}����A�vC��#
�E�"0�M[����`�5ۍ�(���,`�<{�Q��O�2��C}|��sK]	t�fV���E)4��������j�Pا3�̓8��G=[�/Z�7�dc�3����U��S׷���i2�u�ٴ�م]jGwn����ӏ�rٸ��q�\���T�5��\B�E![�{�����+(*_X�=�����Y�����v��n
�?]� p�ڭ�� �����7�_�l�>.���r���}�-��N3�Ǔ��B*oG�֡2�sO�C*�/�>���J����]O�s���{�����3��`��ؙd��P���b߂V��9�Z��P��u�νqE����D�Anb�)vnN����C�{�V�5r��)�kC�H������s�@9t�c׉�<"��}�I&nT��\�N��ST�칃z�-5G��'1ZI5|��*n�J#2�M��o�h[�j5
���^�ɼbć�V���9��g{3��۔ҭ�x�n�/8(��,&�v���^�!�+Nΐ�q�&�K�tu
Z��ӱr�J6e3��0��eq�C�����m3��PEh�<̃&o);��l����oj��M5[��nҕ�Y6�@�F^��؃���e�*gYhJ��-໛��+�9��h��L��vh0�7]p�D�ٷ��V%�u�X2-\V��50����.���a��yVK���[<���`��2]ظ��"�س�ڦ�b°sE�Y�D�S��ӥI�;d��]���:����<�����c�1o��hΥ�Ü��l���h�Pp�xm+T�w-�ՙz�Bm�Ye5u�pBr�-���͗T�Fetc�-�uHI�W+65kO��p��zj��!s*�a�86Sf�X]aۭ���H��k\x�y��]��Y���H+,����]U,:�DQ��k���+�AJ�!�8Rb%]0���`�Y��oBI��{7{&�KȜ!s9E���\�e;UH�1�]�ǔʣ�om�km�Q�EM�,���\6>�^���y�"���]Ѱo3z���js�B&A���EP%ʼ3�1s']Uy#��V'�ι�Uhf`����@n����[J���]P��+F�f�݃�ޖ�/f���9�k9z�u����������+�3� ȼ�vbE<������
CC^�J�$:bm�9���̇3��î�"���F�a���p����{ນ��+V�T���>�fvwH�A�)���
���|�vM�����,�\��M�@�}�lJ��o��{_[�1;%#���ɡ�9�n<v�Gtq�Db,n� uڷQ^M�j�y��]Y��Tao��DV�g��޿C�M.<8ӊ�ڹ@�w��ԩ�c%��a۪��U5��q��C��mF[wnZ���N��f%Yǧ^Q\S�3*�S�9W4�{�Ȳ�'�q@D��cS�h��+��
�k:7j��[�o!;i8V��ѽ�Rg�m�E�{���wu.1�wmeu5��
��z6��Pl�0�q�=��UP���������.�����F-a������ڬ�x�GC���'r�R���\�hk�p���H����+���ؓ�8�T�H0Kʖ)_��˱�]�e3�Ys4rE�2p�P��!��*ƶc���E��J��f`�����ʻO�Ԭ�I����a����V�z��I�$*�|9��bv�F�ε�4m��|�sTF�4RTA���/�������}��O��~�_�?H1?d�̓%5Z�*v�]�L@�U��g�U[�s���~�_o�����}�߯�����I��Y��E�iJرG�9���t-U�(�4�ېrJ��Ѷ)u��c�Pf"ִ긜ܨ�1}�c�4Fձb�(��s��[Kb���ů�%,m�t����؆�0΃A���ژ�5��9lc��[C��8�[:�3M�E-Q^<s��m��"#�o5�<DC͊��F��<�q��cP`�T��Q�QU�Er��v2m���s���4m��x�8lnn[��UO���x����p�b��5\��0�h�\MmA˔sm��k�lUF������$��[����m��׫xɩ�&����h6QH�
_�& ��-7�.��y��m�Kor��&���+��;j��;S��Ӳ�����Y�b�@{��NGa�s��y���x/7���7��cM����@��*���}��u~� �:^�E��tefAI���8��N�x�R�uƆ��:��p�s�Q�gA�x���m���'��󠸭�5��e�T����W�7��� :�*ّ�k�5�2���6&�@}���oOW��Ϻ�Ċ)%6!w5�!hM��kNd�,�<vq8�d�K��n�@#6�qw�~�5��2N�aK��۰��3�*�u� �(U�6�g�ʹ7�ي3u�R7�R_!�]�=�_F�a��T���Ļ�� �d�����`;�hG��;��ខ��{:�25���ex�_%��;+�wc��~�;���q��փݓZ�ߗIx�';6Y���,�K�]�����i~�᧏>zX�(��������d��f8FP�SO6�^�c�v��=ϟvؖ2,��^m���w5�et4+�g;sВw{���m�e���v"��
��y�i�`b���mM��%Xc���1�Rc�Q�gT[y�8����a��r�܇����<������5yt�d�v�OS��X�vj�����sF�mj�A����O�z�~����7��a�4������{�^&��/2:��
��츊�
a�`����f��a�8�â����OKX3A(z�ꉳՑٔ�Ƕ���>��G7�G�Ei!�vq�g�mm��y�Q.�� �����2�襊�߈ �ew�V��㷃�9d-���#�m��fyUf�tKКg@�Ū�7E��Ҫ��g�}��y%�������6�x�ۤ�x�"V�j��Jw.}��Й����L�gH�+�9�"-�+�+z�a#|��A\i�[0I��`k;*3��w��Ԏ�p�+�ح2�_��*��W��3Mzxݝm�n��V��ϻg��;K�
��s��1թOetr��,8����g�[ݮG]f�'��~]�^��u�70a���ޱVwA��ҋ�8,�n��Dq��]V�ʭw�[��{�C	l3c�4�9�b�dm�mF�f�6�u3�z��j���z=�7�>�խ�	�hro����k�q����Y��l*Dwr�Q� uv.���Q�j)|�z@�Vf�ֶ	{�k�7UR�C(�%n�M
*P����٫�@���{rg>%1����wj�:�����_����������aߎ%�N|��rD�Zl�3�Wc�q�YV��M�t�V_���c)t�#�c錌S/���׸�&x�L�a�`856x�rF�tާ����&Yb���m�9�Օ���9y�0����*��V"k����������Z"�f���=��z���yd*0�`��f�U����f������)=�F���n����b�p:]y`�ח�g����C=%1�tk"Fd�:shkYѭnјy�����M7��ܚFe.yz�g�~�	9��j�6޳��>�pѸbc&��)m�� +�>+��%e�U :Y�"��|�Kw;A��hY�v�c_�qȌ���%^�SؗU�ܸ�v��=}�M�	wH��K&�������,�u{�H��N(s��ׅ}����/uk�M�V�.�FLw��,�"��0R�q��jbh\,�W1���EF�L�o��2)0�	��\�b��@��Y��їΒ���^���T�t�]�:���*����1�r����v�.:9��+�y��D�X"�\���+��qٰ�[l�W>�W{�%�A�>sd��y�ީ���g�����o���I�'ڞ�k�S���:+jx(�pP�%U����K�}����Ry#(�9�Z������NAۂŐ6���<��w5ٹ��'���SQ�����<�Y�[W���m�Hq\��2Xa���+lwN>��0�p�Da]Y�*�F&�s����I��Y�+1y�M�����>��`S޸�N�Ҥ?u��^[e-�K���}J�f[{2n}�Z�]�F}�ӣ�s��b3�qYԩ�o6*n�{���N�Aɣ�p�Ux�Ⱦ����9� �m�
������u_4�x��xM�owz�Z�FVk��h���Y���ȴ+.&[k�v�c��ӱ�+6z�+��(�Gr#�q=��Q�6)���pa�=o^A��8��^�oI�-�&����6g�č�q��U���Ow���u%hO�/t���%�i;��؆��{������cݟOT�R��P��xTC͡���k
�����<2���F�l��@�X9z���?Rl�z�ڷ9x�U�iyJ�ڔ�7u�K:W�_WSK��t)����㺵kW�C��������y�������c~zy5_�1�hC[]�"T����r�[�%g���*/Nݶ'r��� t�u��1�U�8����!j*Y,ޘ5�b�4�[ͧ34
������y74�@��*��v ���w�!s��=���q��yߺ��$;g��R�)3'*�ڧ�
��<I��"��2/�Y��a7���]���� G��}ݬ��*�EKd�]:�.m��+�wY+3D����`�=:��P�wIJ�������=GCd�#��8�c�;�$�5���#�:�lMk�����9�(r��6�kǼ2�S�k��]�u��RG�9��jc땬��C��.���=B�ֶ́(�c���g#�av��73�oW���(������E�u��A����/ލYU���Y�%��x��-Wp��ڙ�����O�L��i����� ���}���׋P�&�W��ԅ�����#qv�G�~r�v��o���ڗx/�vi'}�f�>x��|���O�tv��*��p�
�����!\��t���v���JS���Ԙ�5����
�����vd�C���魡�3R�d$�_V��H��������H���?�4���g.��;�3d6��6�37�ϵB�C`ډZ���8�����U�H�K�����z8�s�>��3��ڥ�V�L_Z9z���o�00�4S�~���Ao7O���:Gp� q烢�B!�e���v7;�j�CQ���1�M�R�t�ޠ�����~6��U}��&N����hl[�CXQQk�r&��� ,$tՊ�x���j���]-�Ek������3��OK?��P�z�l�4$��a��(B<c�=�D^�Y �Ptu�O{�9�m���Y8 Һ��X�p��K��n��Wz�h�9)�fM<��v�}�OMcn�YmQ�9Ź�8Є�A��o�B=Z���9�%`�"R���M{�S�ά؆�^�ؚ�ɝ��w��բfŌV�Z���Q����Kⷮi�ؗ���L�N�����c�s�]#F�]У�,����r�gD����S']�٭~��:hr�@,���)�b���Z�ܮ�	�Ʈ��Ώx�Ș�Z�Z���Qޞ�ʸ#쎵-(�e�ad6�oe�ѽ��c��2��z�~�j�>ky}��x��Y4���<EE�ׯ��~�w, �G�.�#b�ʾ���%]��d�xۯ�%��E帛\��1{���&
�� ]k����=������m��}��79u��@�#@��K��v6]h_��pֲ8��P���yO�8�;�o�υ7q�V��P�g���>�`�i��3q�����MC�%T��F���oT�Α{ԩɹ=�+��R�] 􍞦��5����}����OE�`p&}���8W��~���9�:�|ȶ�gXQ�nO�Y�c5�]�nD0@��02/�%B��+<_�Mn3T�P��G�s�FJ�� �=�t�4��U�Y����.�K�x����>k+�[���Gz�Hh$���k���3�Ba�-׼B�fc��Y�z�j�fb����vB6A�M���tS��8��Ϭ�w&:�C!b/��v��_D�u�3�D���q�Z1نЪ�E�����3c�cIM��ʠ��!��:8֗!�v�щ�6��F	[)��2=�Vy�5%���Q�
˓,�b�����c�G�붲)3��3
�5]�TM���S�z�~_������͞��3Yp٠��(҅{YfAG@���sN|����Z��+�&���#E8���)�܄�_8�+�4��b�AOcTN6(��f�o��a1�f�M[!�@�7�\����ºR�u`v���v���N�ܽ�kg6�&�[�Y�W �0�
�DV�z2�>{qVs\�{?q7�F����ߠ}���u:����8!�؏9��Vӝ.nz��i��+ �*�<�O�n��Pww��S���]��_�^���eLi`�7�P����hYMF���:��>�t�f��s��5O[:���74�gp\��t5��Fwu�A$�1>���	ݐmu�s���L+��z�+c���g,ǘr�z@��1��ݮ�ܖ�L��^(���ۭ��ϧwOL����s�+�����d@ˁYԨ?#�B&�`���46ã	�r���wR�q_�}�M��Vxn�>˦�u���T�z�^�ww�W�r�G�zn�Ϊ�Q�vR��5�o��wNU4�&�[�#9DK݆��c:b�q(���i���,:7�Zb	zթ-C��1�u�om{��7�Z7���9�z�N�K���L�J!�G����#�$0�_�8�ϸ!��9��7�L��mϷ�gݢ��5k����'z��x`V�65p���=9��{�̽�SC�<X�=��Q��O��eU$��09�{�d��~��& tyW��U^��E�ԕ��|��|��;\�Y�;{��e�P�b/�&�OO^�.HMr �F#a]n�`�J��-�ݷ,v�$]6�4�W�=z�d)�n1qZZe�"P�n��v��W��H�����G�$Z�\*��XU#�D�]��w�S<����zz��b������L���j�S��p��f�+�wO`��o�sl�ڊ��@�FCw#@s�J6UүU;��U:��9Cr)���Z;���D��>|���	N�?t��q�y<uw���sB]^>�޾�?4�i�${g��g���Y΂�;�\��OĈ�����^�R8E��;�k����	������=ن�_Jl_]����"�*&��:c��&�1�w�RG.a�n��m�N�_r�k=]f�zc'O9��M�X��mG��}�����n�@ێBۂ��t��&kSEi*+Õ.I�B����0�މ��۽�6I;��ǮT�w�an�l��腯���%]?i��	����Mͧ���kn�=�"U��ǂ�3���C6�댈�O�x޺Nϭ=�/�.T��^��[}zs	�Q��3j�Q���`�|l7�8(���wR�cwq���|M]~r����soCSk]^�o�؊�}��3r�����MQ|@�e���Zr}|WPc���vO��I�/���F��kJ���l闧p��#a�Xl��E,���$��6������]��U�3����Q=��ƞ���Y�g!D����Ѡ/[�y}Ǆπ�=Z&��og`"z�1e��t5��{�hD��u^������fg�ڈӼ#wr�>�ѳ��0lӞ�;���������O���_���AUEw�
" ������DD���1�e@H<ϓ���f�8�C*�(ʰʰʰȄ2�2�@��2�0�(C*� �0�+ @ʰ�0���C�2 C"2�+�C�2�2��C ��2! C*�(Ȅ0��CȄ2�2! C
��E�A�A�A��a��� �(���� ���0�0�0�0�0���0�0�0��00�20,0�202,2,0��������2�锹�|�@�� ���#� !� !� !� !� !� !� !� !� !� 9��@a e@`@e@a@a@d d@d@�ȀL��"4� L
4� � �� � ʠL
��0#
�0�32�12��!�e�eBi�HdRD�&	�e��<!�Hei�I��HdB@�!�a���e\0� CȄ0 C �2��w��=z���� DU&@) ���~����~�������O�O��}��_�>�����e���w��9������?/_����ETW��������Q@W��QX��/��� $�2��?�?������ETW�<�������Ā߈z�������O� ������b�0�DYE F� ��T�E� @�" �( A
   JJ  �JJ��H��� ) C( @� �+"(J���B2�+"� BȄ�(I�	 �$ I !, P�, HB�2� P�B��8~��������'��" ���P 
~C�7����|
�G�����TW����~�?�����<{�z_!� ���������o��O��9� UQ_�?D?�?����
���j���������TP߈~��A"��������i��|/�=������S�g�| ��TV�����_�
�+���=~�_�����~��>t?h��$�������*��������UQ_���?w�<�������N�S�0�������~8��������*�����g�� ����y�{_������_؊(
����׀Q@W_���������8q�?�1AY&SY��n�J�Y�pP��3'� b=Y��U%P�@(�tФ%$�ЪA!�5�@R$DUP�%DMeT$EQ���B
�J��RPH&؊�`����c-�[6�3+m����m��1�٬�2��k`SUSJ�5-i���f�ؤdjͱ�j�Ya���c6�M�Ƴf����mJ5��jִ�)����̬��i���f�b�ƶU+f�M�E�c2UE[����3i�,ؚ�����mj�m���*�i�����ƫY�ٖl�V��[P�o��(STl��x   ��ҥ}�ݩ�uށ�`SoE9צ�Ζ�g�.�osuvی:��(���v�,ʝh
kk׽T�J�������S�nX׷��5F����Ӈ[x�F�]x�Jm�"��4ͥ�+-5��  �C�hhd!�������P�B��|xz(}
 �I�z�q{i���y��UA��75���3�o�\�n/n�O;u+B�]iۜ�=g��N�5�]Ԟ�c%�ҫT�j͚-�Nƾ  ��*��[{�W�ݽd]�݋{n�m��V��v��t5�[�m���ۮ�+W�\�T�݅��Os��{k�3/;���ѻi��cj^��Ӡ[uݝ=�4�Z�cZ�Ҥ+��co� ��}�䬭�{y�M{�M�ne�tu�[R�]��r޷)[f���9��1�s�ɭʰW] �Ov@tQ�֨�*�{�mj��UE{l٪���k&�km�b| n��5�]���]�hg�w^��ڽ�d��� ��ӌ�f�w\��^��Rm�n�@5�]q�^�]s:{��Z�u�T=R�wR�LM����H�F����W�;�]WZ���������E:�I ^�x�[K���=W�����j;�nITw[�e�����ݪ�/T�ŉfb�Zh��4�� �{�Ҵj�����Vx�w@��n��ujǭsy�=���� �@v�MӀ�\�<� :7{�(t4�{*���2)��e��m�  �  }v�[Ӡ �7�[��y׭��r��=An�� 4 [�p �K�3� �j;{μ��z���ΞkZ���cY��[b���4��  ��  �N� : 1�8 �g��� �� ��,)� W=^��x� �;�� ^���� �;����km�hKca�Mb|   ��}�+ y&��@s�n  z7��p׶ :��4 �^�x �zwz  x� {�� :�ɼ   "���ʥJ�� E=�	)*�� hh"m1�T�O@��S�A)JQ�  jm�)P   ��H��UD  3S�����|��G�~�M`T���E-nZ<#��r�4���nӝ�)���UW���y�K�<���Z���V�����v�ֶ��ګZ���Z�ٵ�m�����<�>�k�u��(� wVn]"��JK�h��@ّh�"����]]���Kj
.Sx�7w�(5�w��B�f�&�@nٌw<a��F�e��(6��7(�ݣ�vBtiH���b��Δ&�K~	V���ov*2��8wsB����ߴ��T-j��:���
5X��5�+A�4
xX�4�A�l�h�7u�A(�z���QT��Î����~�z�]�L�n�u�ki#���-Ʊ�(�Gq�w�JOT.�����zj��7�k?]9��E�KHu,�5� /RQ\)����ŗ�n7n��n�Z�#�U�a4][D�U/)��3(	.*�5K�*6bU��X��n�6��^�c+1�v֖>w!��6�kL���e�4Z���KV.�L�PO�	��(񕊙D�6�P�n	V�X��Q�老%:��7z�*R���0�=���AMY<��U.X��yYRٚ��!gĮ��R׬�`0p-�x�hۊ��7>���h��srټ�
�ei�x��MGm<.���:�&�L�I��7�7֙=��j��T�C EF����ܵ�t&쳆���^<�Ih��MI�5B�Ģ�-�V�	8��U.hB���r���Ģ��`2-!���HX���MJ��t��lƆbۧ���r1��T�W���MQ��V��E�[V�-�i݅Z$�F���)-�PKy����J��.�T,�¤u�+�H��nCZK��Յd��M���4P��M�b�#c@iv��M��c �6���2��c-%d;�R��^���Up �o�
��ʷy٥��ni�����٢�SY�ˏtʑK��Գb����ГB��t��	��2������Ec�6�KV��Bݴ@�{�l̰P+����]�7k��YJ��KYzMy�d �$&Mk���ȤCwn�B�I�X�PD e�$nŧ]l;m��ɩf� ��d�%��T�l�T����)T��^�ҊX$�Ն�fQJ��ͤ
x"�!��$,�cp\%PxB�w\LIEa�yW+�#kt����`���X�܍'zn��	0���^Ւ�(�����ڻ��@��1TL��{v��e����-pR!*@�.����k����/��e�ψP�emAS@M��܊�[�˨�4P	2�.K�6"��t�����=j�+��%=�����Lm��J�Df���MR����%x�9�7�I���PX��D��ͺX8�ZK�GAٻ��n����Ϧ��u��H�fϠ���4)L��i�:e,����u�AT]�����ю�%�i�k3�Lm���9��a�Q:)�mY�L�%^��ӫIH�Rl3Q���&�si�K �tcwM0�[��mػY1a��3�� [����af`h@�*��g�fP��^Ь���b�)��hQSEI��y���^�e�m �����[,���6nxVV�K RƋE�j��n�:D��"�|��3�ŻG"455u1Ĕ�����ͩ����-] �U�{�`L��v]]Y��j�BQ�͕C#y�/nƂ�[��;��iŻ^�:\��ƥ�WJ��a���^�$ۨ�ʷ)1��u���yxSnb��I! ��Nh��xZf��ז��.����u�m�D���UD�♦��g%D*���洖!wU�S59�<ƒ�]!n�`�I��c7C�b�VZ��k�����v�iM�$���̢4ܙ� t�������&�P�$�r��!{�H�ѷ���+[��J��&���ש@A�GF�*��� ���@��@f���"+�c%.;C����Ewm�^�NP�(bh��v���]���Z�Z���HP�uo ,����w�-��������(�%�ٴE��V�Y����ZZ����f!�Q�@�e]��6��#�J�T�C+p�WI�f�*��NJ��i-������
֫-K��ĬǸ�����u�n�k�baJ��K��n�UxP)�4k0ޣ*
���MVT�m+L�b�T�I��֤���ˇ���07"!��f�cH�]��v,�,z4���:x�[Lk�mն/��
��w3!�c��EV��x��:ZV\n�%���M�P:�&�62]��R��!�)��{6�m�(c����mS��k��C4/4Q�l,�G塝wZ�d�bŶ`��fՃ 5�P�H$�O)�mZNŵ@[�Xn)��HC7���5�}�E�]$��_�uK���-@E0Q�V��<�M0�D D�
[��N(�y��F����u��j���Z���'a%V9Dj׆���,S�QzXL�E:9�-�B£�'B�ܭҮD�j�
݄hd�6���M�/��v.�j�fCp�.�B҃4�e�i ���^z����|��j:�@`�+v�ق��9&D�@�@�a�"g[�ˀ	Hf�2-m+�7�Ҭ���+^ۭ"ӭ���a\h�;b�W�`�Sn��gU�l\�>�iR��c1Ya��[�ߍJc���Uv΋��^�b�z��T/ͽ��I�o�P�Id��mɲӚB�;סX�v8Ѧi��y�B����ᕊk���qغ�o�.���0��@�J5��m���HUY"�CɵcR��;,6��E�7E��ұ����[YL�őMvځ⵻]-.��|��W�� VfJ.m304��ܽ��vM����̬���)�"�A�s&-�aJ��hK�:�n=��k�q�-�6j��b�6�N\c,�{��b�h��������[�sbo�>ͱ�J�왮[�u�V���6�Cd����n;6�R�mق���Q�8º9�|aB�*v�'36��j��`�i�)�=[��
׬���)��L�o,�V��X�e΂GD2�Tk��:�X\ܽ�XV7�i�P$���ͫI2�ܫ�$0EM��/
#���$n;�ѱ`ŕ-�&��m��8��i���j�ȝ�C3^Lf��-���ۖD���K(�B�ޣ�A���ɹ6d"�9
��cx�w��/o�����l�݂c�� �6W%R)X%q��e/�8&c�3�Ben���;՛v�;#����t�Rz����I�����ڽ@�w"�+7]�r3PӅ=��`���qR4�����L]@���=D�f�&P� YV�;F�7�+���)��h��;A�L<��ƶl�n6��>K�%n�D͛ġ��ӱ��ʷ��2,wz�
M?�㡫.�i\tFm�5s[�y����;��7#�V:6�S�*�u�L��0A����r)���ii���d�l`	l��5-j.
l�m)	�&^���!)��F.=�YC�R����*ka�ۄL�\.��@��F�D�˨V�(VV���W p�\2�*C���6�܌-���a�x��M�LA7]��1�F^GzL{�ձqRJ�l��z����)����<8^,U���q�f�ͪ4��FJm�"�ơG�����V1���T�ŏY�I�Q<a�a����Ӕ�n��3f6~`�@���+*G$*�ީ�\��|��(��V�6�ĕ�t�=��ù�2�bYt�˵�AR�E��]�t�(F�@�V���**�+h �r��4�ᖉ�wlTR"�D�V��C������V�0!�P��NO�3nVIS9��"�E��Ό׆ӎ��ǭXb�n^�enR��Ʊ�[����3D����X�c\�4�a#��;Rm`���E�����D�k�A��g]�n�L��@q�.�֚ܓ�òhu��րl���+�+�zJi�dF�sh�i0p0J�@r�$��PZ��a�Gל�:J�cX�!��ˎ�ɠ���YP*owL$�]�-���Z't�����n����R4DQe�&Q�Oq�qZ�Yl�V����M��U) V�G0�x������7�+�X�Jh��䂑�ؑi4쇖�Fd��E�u&�Fh��+���^!�SԀͩ j�T�Sl�	���
Z�j�$mF
�:2ܛ�)R�p-H�����R�H~v�!f+�kX ��:;����V�hT����`1��(	#�;��U�v����7�ՒV�s�S�nҢ�Z��)Oe̙�q�����)
$I�B¬��l
��&AN�7%�(:�_`�be�z�CU���ͬ�v��E:�*����PބNc�M�Y�<�4��8]c��ݠR6i2��mZ�i=�R!*�ݍv��C'sJfƻ�ѪP�	�ni�
�쥀r� ���������)�6�@����WjR�+#�2�Ď�1�`�2��tq�^9�v'�U`F���9M�F����gn�
�����V�5
���q;8�,�t� 0&P����u�V��"R�Ht�I�CH�k�2\��֥�cʴ�"�,RUf�^I[M����H����0����l���j�,������p+k%���@��V�TN����Y�
�Y��՛�R�RMa�F���KS�_f�&ۻ��ԧ5vX�×�-"n���EꄷaRܱ6[J�^d��Խۚ�A��V橍�-H#Cv4n9p�#&b�+�q;�h�n2����t���8�9	q�w����JSD���m1J`{r����ؽ72�cĤ�Y�佈�t�+�Tc�5P!���(�* U��XM�%��)O!:+EcѡI������n�cPj�0��7�(!����{5f��`Ӑٴ\e3�Y
�Kr��dB���m1r]t^@�t&�hkס�c�*�cB�i'
yJ�%�	V^���pIO(a0��15oW"��*�l�#)Ċ$��I�:����\&�4���Q�����`�N���VI7T:�ln�OT�V:�Ye� �JʻqT�����������K	Ԍ6FW�k�^k�h��ܻ�������,Q�����]�eL�r�a��YT*�@oBO*���
ޘ>D���Q1W�[qP���
)c�5����=�����j
�c[e̥��j��V�y��M7Y%�B^�nc�
��{�(m��@(
A����(�t�����t-�=Lb��&��k,��@U�9G���t�Ue͑i��ɑ�&+K9DS)E��7���y/M�[z������#>�]ArdVm� �	�
���3&�6�"�I��Nu�A�B*;���Y����p-t��B}�ތ/iԵZl�{�E1X��!X��O5]�������J,�(ԻO%"u�ɰ:�t�n+-,��.����·St�JU�Zl:��*����U�̽�iS����	�?��ԨyA��i���^��jx����rz�MV���M
3 9�L�����viw*��@�Q�DQTE][�6����C"��e�1chM7�	�Ov��T���f�v�,Wbh��Lךt�Z2�Ĭ�
�U��ː��JS�%�V��G) 2*���i� t�/RǻtN�~U������WI�:UЩEv��������dh4i���[F��J�p#B��Z�ߓț ~�XD=iia��7>HV�lLf�4!�;w0Tb��ɻ����xºU��"M[�avV0�	<8$�ٕ-6�V�Dh7��Nj��}���׈I��޳�ʙ�v�Dݳ1 �t(D�2u�5�Z��u^�n�Წ=Z���i��A��a�O���WZf�4��h��<-f�/- v�U-?^�H�kY
V�Er��m9���Rlx�7,6���#�,�����\�R-i�%�ZE(v�W���4c�5��V���i�YE��Z�ݓV���9!Z�f�.m�������sE��0��a������k����`t�[� no׵-�jʂج�O%��l}-���[,H��PP!�W�!��"T�5���kU1�"�XoV�2�1*�>�weT��	�a�Ͷ�)����mjt5�yP�.�2��,l�N�JԾ̡F��j�6%�� �yBU�J�ף2�09��lj��jV�Vq=fcM���o�:��aZ ����|	ъ,ú��֨R���\��\�m�y�)�*�<D-T��㢵ѭ�We��!�.�����`�%��(���Ҋ�QxeKoN��B�c�J$5�k�c0n�Cn�t�DV�Jыu�S,^�ŗL�WkX�'p��M(Muyr�AQbh���ۿa��<)��k�Eh���˝��2�َހ��[Eէ�*"��[LlƔ$�Gh3+e�r���:�Z�KJ�:��3r�*4��]�Ğ���jH���E���ʃ�^�.:*��#V3vê�
n�E�vjm��c����B�ߛ8�Ou�.[�5+B9W�Jx�I
�nZˬ�q\����	Hխ�S1囀Ӱ�7���M˫[� �{W���6j�1|���^[̭W��sVm$���`�	�b���81�e4�l�8Y�\���ۂb�,�hU�w��ʏj�9�$���e+���M�D��R�;��ub�l���u{T�2ɹ4�U��Jҷ�Ml��Ua�Q5�e���E�Zs$�b��)`� %X�*AE:��-��Ɣu��*w�n�K�O{�o�S*�%m�%6��G[l*�y�3y��� ��hiV�hJ��I�f�<6��3�[���T--.��5��WC�;�𲉈����Rh��Xʐا��d4AGiA��3dr*��-�=`�zջ S�&\G6�� 6�FiS(Z�U���SK���vF��'ĸ��r�Pf^9JX�݌��$��Qm�{����;$"�j"�Y�����M���0A�
��o{N9]�~��0#J{]ֺ��:�m��Ux"�P�!}K(C򮽬G��B�ck:��s����7�	�xДj]�oy�����g�hj��������@^o���60w��9n�eژ0�f[��o����F��<˔o:&�^��[�;B̊b���wE��UՐ��N�ˡ�d7�<9�B���Y8�&�=��ut4����������R�]�U���2Z�5��.۽�Ӱ5z��ʹ�i�뼩�K��܈��c.���G��i��O���}�����}\JzT�a~6J+��o�Nu�#�ĳ���W��HY���e[�2:��Tη�so6�Wun��[с�D�#�kt�#l���{��㽥��B.�>a�,�S�n����C2��e�0��e�{'&	PհJ=3���g_fS��qj���;S���޷��`�x�:�at�w���O:��جO��X�j.ܣ�ka�K1�e%��t�p�X�;+;X�Cv�31�B�WC�|z�R=�R#� /�D�y�7�d[g@+\#���ȧ�;ι�u)��ՁoYd�i������v��[d�n��J�Ep3d�T �9LW�_1/���2W��WR���:��`���N5jP�yO]D�Y��*�9^�w7�/��IN��&d��G�wW�����xD�b{�I���U����S��_E6wx��vB�)R�U����^���rY��Ɯ0�����P�zJ/hݶ,����Lwf��(�ȭ�$�+yD�]��{x��0ݪ�#U�ɬ�3oo#9�5��$��@Z���f�������!��w9�Nd�/���Op�<���K �O����Ui��Q�;Vm��ԝ�F�wA6���x�uE���G
���;�Za���i��qN2�\A9a)�m�9SlcJV��yhfDw4R�έ$�˧
�&�Y��G�h�����WÃW4�����WZ�E__�އen^�����I<؜`}:��z��y�Q���m8ka�]������ah�}�驪�ʙ0�J�6u����!�X�%,���̅|u����)X7w�)ݩi��h�w�z^��p��ҽ�P7�Z�%nN��ݥ7�+���hf����z�^�)��/��6$�Ϟp0�To��S6*�0.,Bk�S��d�-'5��$��j��v��řz؆]r��/B�[ݗ��O%l�윯�Wdڲ���r��=Ë��%h�䬬v�<g]�Ե42˧���`��/wk���ma�(��]�C�w\�WdS%���A9Rnͫ�i�/+JsEԡaS�t���k��*'B�wDgs5�Ψ�G�-��$��o\X"B�:u%Y�oZ���m��6�:�D��9�p>8o�����񝓶Y ���pMBqeZe�m�'�B��o�4#�`����c-_�&�WM;*޺������{�j�	6�F�7�r���̓; H��6���M|t�����N\�9ױn�b��![|�cr�u�{Ԇ_f���(:��֫o6�4��.?�t/��\8��ne�^��*��PWV�k^+B]�pg��V��IAŏ^Nx�r�ϱ\�}�$�p�[ �	3a��M��`3�p|��ST4/�;7��X+U�Њ�iG�VО@�I�C0fj��0��`'��XE{k�&!�ڃ�5��͕ww*VK��c�`�|.�'���+U���I�ўr����=}AE"W��5�Xg	ȼ�>S�ɠ��9���z�upS!�n�ӆ���l-�M^vE���jJ�&F��%��X�U��A��(G�U\��^��7�v�t��6�K1yX�^"��6R�p���E�qk���T<q>G�υ�Pz��ҥ��}5�8�04�yX���y��u����*�ٲ���r�^>�.�j�b��x�΃�svK�S�n�s#��g��iS]�-cp_9[U�RCx�Q�Ъ!F��j�.t��!d�3�hNeЬڃ�oC���-��g����n[L���z�9���6�Y�B�P�]��qc��C�2��T�Z���e�+���z���	��s`d�[\�&+M43���x?Dh!j9��
s�{6zy�.�G�I��ridlG�����u 8#�Z��.��m�]��u��m%2�X���Y`���+v����X�;��.�[���ۈ����t[�����`��̧�;��B,.0�P�n�Ö�mk�M�b|��^�4b���:��n�<=�!�m_W]j�n@��̔fu7+�ս�E4�y�3V�;aoJ��B��-��q�����S�W�@3�U�`!�q�B���VU���+���Q��ώ���B^]��=74� �H�4B\1�&��Y�u`U�W9ͦ���[A<��@�H�*¹Q�oj]�F���#�s&nd�=&u=�}B�l��P�'3Aa�`��!7��O *ﺞg
r�%�o�3YS���^d�O�U��L�z3��t5��<j$����c����D��%;�Csy�t:�=p�dWq�Fd�b'��w*��{2Tj��h>�7�V3�����39��ї���"��������5�>G�<oێ�?w{��I+��މ��ɽ�*��5.Wj���ʊ��y;_	#�׫%v~C��e��U�hI�^�z�>s��^��*�"�}ܣ[Rq�v��}t��{4�њ�DCG�Wd5Ҷ�$����	VU��QL�{�b�׶�e��td=��*���q������s���i�
�]!
2�ƣX��T+c�����듍<���*uyS7���泊�^�nѨ��k~&	*cy��Q�Y��6ry�KN���f��������1>�A��u��b-�<�x�os4�¶���U�2�:Uۺ�5���"��x��
����*�����u��n��L���N�.�t��n�z�����Hٚ�WSPPL��VF<�����k:c�]�U,dse�O��C����Qk��	.�l9�ӧb�ds	W��CՔLowQ[�i�"�侘pi�l"j`��R�$v4�t�"U�$�Р���;n�6 m	����͗1X��O6썡�Uݻi!Ʊ��_v�����ٔ�X���g7��0�I���6�<����]�C�(���[��s��I�\��B#=Ȍ8}���f=En0��H�TN,�Ew[����֊�4�BܐTr���x>�H4�W��{�z��B�-��q-rp{�#�eӥ����6:LJ*�\�MeH,˩y�2N�j_��w^|�f�f�
�w��V,�8-��-�����ۛe7�����vo��@���i_U�5�|�^�r��N	f�e��'�k]�k3� �7���8���<�wi���t�<��tVi�H0
V��xl��k��]u����3.�D��
y9�$���&r��:pA��˗z8q�H�{��h˫3%��.�V3����B��ю�O�2+B��Ipy��Vkw�.4�R��*�v���uŕ/oP�������PJ�1h���v�q��eYD]����$��:l�D/q�ė%�;�ŉ�r��A옦���Z�)S���Ԏ3�9�:�'_:��ޮw�f˷�bw�P8e��f�H��K_X��8�n�>��w\�7Ir|��F"���!��w[ �w�	��t�ܺ�c4���}�B�c����}�	�b��E��o�X�fptI�A�& �uJ~ӆm���V��{b�H�;Mr�9"�o�ȳR�'_��%+ǜ@��&�=,uL����w÷w^G��>�3����X�X�{ћp���kgH���|� �v�0�=�e"��SF¢9*g�(5\>���v]�h�3QN�\[wn�I�Ul���Ϯ5�Ҵ���Пd}H��Q��!2��<[Lj�j�$��J�ma��tG+��fǉ�_.`c���(�X�r39�6�k ����Hz���i��q��G+<��L���wI�l�X<�1���^2���`���(�\$zbΕv�j�X�ӎo�K���5(��xy�%�͒@B
�.S�2�l��@;Z��e]R�ܡ�]d��mVrƫ�`��)���ȹJD3O8��\A�≖�S�f��י١[�X�D�bWY��C4��1"ƁN;��ή�	
>��X��΁�Y�#oa��:����.�:gr�v���;��
�d�(��'\6�k9����J����r�u,��y��Y�#����++lN|Rٕ3I��c��^̹�9��&8eB�V����R]�X�O7���P�_\ZB���ƳQH�ۜ��P�����{�2(�&
��b1�� ���+ʘ��B�ek�U� ա٨<��+j�*V��Hju;b �"�\/���.��E�l������݀eu��qt�C=���Q��h�tw)��z�3��r3����Gj�w��b@3n0�f-�W825\��� SЫ0�x����ȥ��+$Em����ns���m]�f�-�s�/��e��H>ZM~�^b��[��Jޮ���d��Y�K���q�7ί/V�u˜boF�b�gf��H.��٬��3k)d��G�e�[�����&��=���\/x�E��;��n��Y�����+iu�K&�am����ZJ���������٭�*���k8�J�NHlv���\��V�Zd�RɌ⒒�sn�1��)ݚ��Ӳ�Q�.�a�QDdYY±k�[��n�'6-2ڀC΃RK�[y:�Dc!�DZ�ή��y��z̂�q��X�u^����Z�oS�<�q.�t|�˺��M�h˻Fi���2�k��p�{�҉4l&�$J�#@��N�����[����с֪痡<g��2�4�HԼ6�K����J�}�*;�z�fՊ0�\�O��pL�v�#0zrv;�+.����qM)	ʎ�o4&mDm�cw�1$�L�3�ŏ�ӣv��̳��BCN1���Z�E���S
�
y�K���Qr����3��t�ƊnⱨG Z���d�yrQ�_Il��U�SF��$�Zk �Ĭ�@Q��c�׺@�b8-���3��0��_w)R�XRd�f�c�������r�qy6��T����SGܥc��b�c(�Ƭi{�^�d=@���G�������˰l��
�W�T:�ֻ��C(���ڣBA�\��u`��V��O�:���`b|m=��f�ztCij�̿V��o=���k�҈���H��w�.>f�y��.�����②���zԲ�%�x��{[':��a�3C���0*x$�K/�'\�˒J�n����qJ�{�o0xU�Ű��u��I	McϹ��2ތV)3�m�:��{��S\�w[uq��#��o:����Dj[ ��Z�o%hv͕7N�U`YQ���Cx�+sy
W0aqp�6�ͦn����R��ju����k�8@5
�U���ͥ4
Բ�S��y6�F������p�ԁ��`�Lno]=�� ���;-��$�]̫����ׄ���'��Z�M����[\-��7n�i,̎�:j�h}x�c��Z��K�X�I�vVC�$�p�9޷w�B�g
������n�ܳ���i6Z�һVq�&[!5�{���y����Wp����n@Բ�%�_ݕ�4&u�}�מ�Ifm��0�Gv���-j�-Tm�J�8��ϭ��b�/RFΎ�hלV�n�9vv��+��=�5�I�TԼ���{�`�4!)!���
���Es��AY�܍vمkQnZN�)�R�H�f����N�`ǹ��]��%�����9�Y�vk��oq|�Z9M�g:e�孠��{s�/�(a��lR�B:'z�P��LC��F�:�Eu�89���.W%��(�������9�"��z����h`��m��R�v�����L����G:�,���Q�Z%����I��Ar����	nv+�m����(����[�W�0H�1�ry�UdN83��Y�p���r�r^� Y�D�;�9�W�Pz'`%E.^��(����*t����=�#.�y�^��Ƕ��>��Q<�Z�q�:d�S;/S	�0U���杶�
9�����b)֬H�r��T�������{Xvd�,�=u	����Z�g(�o5�4��&�rgB��i�]щ��d�J�.۶.�©RX�ռvYɉ���{y�Op�����'d�(=5�
���hÜYJ�-�-B���.��z.҈'.;�z�:S1�Fé�V�6o�<�ٛHQӺ� �B^�[]uv(n�M=r��+ֳ��!����!C��k���������o����޻�N������R+�D�_5z�͠!�P<�t�Jr	�;����(���$\�ڃ��<����+�i	ϱiɑ$IER�����4�[t��L�x;y�
([���S]��z��$q	
������Vt�n�f��bYppF���b��ooQ�*fNBJݺ}eȖPs_�N�olL 4k�ת�n5\	W)@�ٻ�δ�{�Q�HM)#O�L<&u]&�Ɨ:�k[��'Ώ#bC�s�U*D��:@yK��]�2t��v���sM������P��ߊ�p�C��I�m�� �݂��sozW(�ʸ�oV��BS0�*D��t{�2Oa�����fx�R�v�U�]t�lSѠ� �f�4KG���]Ԁ� ����M�B+�V��]�ţL�x�Ԟ�opq�m��r��1}���/6V���C����~�2%��T��3��[�]�5��pd��!n�/��Jgv� {{l	�1��lQ��&���j�� ���
_.|+4b.��e"�ȹ:�W'��akki�q�1�wi��+*��?/zն���ej�����s�\y��n�~�ϗp�N��s�I��Z���vt�(��)�T��ut���%��R�|�&̈�IJw[/ ��FqW�'U�u��Ӵ�65�.�����Ba!��{K2����P�)���ǃp��	��^Y�n-��-4�WG]��Jw6�K��VpR���h8�m`�\H���CY�W%���e;�.����T�s��"]����Ѣ�M<��pя^`���w�Ո
d�x��2�1�&[U�rmh�TV�/s�K��ZL��4�`^SJ�KgG"�e�#��t��[+��x�r�ۆ�ٳt'/�t�A�&Е���Tm�W�0�u��g����Q"I��m
����8U�u�V�1��m��e��0���{�=�t�W58ʜ"��c3:�ݴ���}ܪc�ͨ3)V��j�>@�b�fu:ul���엷Wg>����.J&�6�	�:	���^�U�N����vq��Q}�(Z̑=����A�N���)c5j� �^�Ai+�-"��{#�!�D�^n۠�O[9(T�R�u�0!�2���u�k����ժ{�y�Ga^���VVemՆs�&`ց]}�3wš�j���.�g)�c�R�#�6��^V��e�՛���۽)jjzM*:МBݚkQp��j��5ǒ;�y2֔���Y�+v�)����7υ�!bX㻆� w6�ԍ�E���i���2l{b��	�%.�^�,�;{QJ9g�r�YOn����Q�nَX� 	�n��Cy��x�秕��()�[]��T]��m�����1�b��8�9�j{f���U���mS��D���6����G��\������yvPn���9u�|����F���V�H'�*���އ����hF�e��x���%za�y%�]2Go��Ug/��>�li���f���C
����y]�5���%���'t֌�ڇ8k�'��k��M�E��e��b�3O�ңfnc�����.�Sk�A׮r�/K����C|N�ս��L���o@:�P�0�L�j��
�M4�L�������%��kE�&{�0FMl#A\X�5�,���G��GU�i��|:a̢�$N4��Y�6�i&��R���{�!@�2�,�s.�vn�8Ou8 �A"�2�^]��x����1[�����6�4�f�1�g`Ӂ�5� �cj�-�(�{��;��|3��R��`lX�����8���`�գ�4�u핡�#"l�`\z��q�{�b!���pr�î��^P-�X��]L݅�M�"��6��+��7u���:�ןsDj\��s���ib7#!PZ�����n����8�=MZ���[I��T��\r�^�6��MJ���z$�����Ec�{3C{L�񝠩3�o�*J�k��1r�:�s�,ٷO��b_�0ᣢ�cX�u�mkR�X�=f��j�t�(�������N��6�'�]GP��Blu�np�T�̈�Y�["��/P���RA�w(��ni#�C�
xy�l���Æ2�YʾIY������ܦn�x���
䅞���:�1��[�h�٣��s)t�5n�\+&l�ҔA�l�CI-�5Zz��R�X��ȕ����iX�K%k�N��l,����������D��I_J��[ˊ��Re(��	ĚYـf-Ԭ�3O�
�b��*&��C��u epJ.pΕ���$�w���zi^�ap��
9u�]��;�*s)<�l��T����Y�7*���ݧ�y��hd�(:k�Ut*�lX�GL���i]�:�<.�~E��x�L��["xm�S"�R�Z8�ٝfQ��ƍuϊ ����e[fKD��6�r�F�������{������:j��e�����o	��3���p�ʱ�d�Ɓ��+�*�q���6�r��90S\'h�:�q엲2�Ee\��)��F�f������F7]�,%Or�����ŜJʼ����5�nYa�U�kJ�gw�*�O-�����-N�`gL��E�m[�hue��Ֆ+[n����G6�dV�!�F��<w-.��'V�m�"T��LU�`]���g@;�a	�nS��s��м|��R���9K˥j0k6�
�`*��o6�-V�`F�=G>f^xL K�3��� ��.ے�=!{'Q`bhK�݅�[J#��sMo�]�2ժ0Q�� |ͨQ���n^���4�qm�g	0r�8^�!����X���W�]sfR1�̂�`\+����K�jo[�G��iR;�|��2��u�S�Jˠ��;/��3��ͩ�@��nN���I$
��i�ԡ�9(����
�g��ȴ��F*�摇D���ؙ���������PA"U���ʇ+m��Y�Z(�w�4�l;S+p\[g����_]crL�:qq1T�I읋����+��l�,
�^�.>���q
w�;o!�^�+�,v�zƌ�v�bhQ�!u�م�\�4��.1Iu�Q8��*���=��Q�t[�-Ko�����%�{gQ�W�ti��3u�H�i\#̎�Ջ�>us���"̷��2r����2�!���)�-� =yuf���ׁv.sb��_+B��2���C{Y�8K�b���7Sn]e�)�i![OEX\�Ҩ;#8������>INʑ�[�k�4����N꺾�lO��T����Yov>��N��3�����8k6��_j�`;[&��5u�C�^����7x�-�uuh����)3o8�ُ��,���0�mݮ"�~ɔ��@m�/��Š������z����`��A��}�\��}�c�n�4�7�V�`GZ0D�u�n���y['وhR�$>�'��2쉈P{mk��1
];��7$�w]�a��h�I%�y��K���H��Sz���V��1���Eϣh����x�ӻ�EQ;�����)I�;(N�le�.Iۨ����]��Ҡ�{Y�	{���fIi�<�ݼk����u��e�|Iٶ��BIX� �ޙW֗bo����� ;͍o.��u����R�ts�M�؝dn�A�	}4�KQ��^���I`+�)�G����+�̶��ɜ��Z����e���#
F�.�<��n��Gh��m#���e��G�Y �,�Ru���z�e!�Մ�_`�-�w���u�*cb.Ն�����S�r�9\F�p��f/�l�1	��c�,	�L����d�Z°�Y�����ʜ[��r��ܬbf����Ve�)H>�M��].2��KL,pzL޴/����T��G&�cUAR�[�&��;�Ro^b�g1r���֣�(Aآ/wt�O���wY���=�D�]�vy��]\2���"�k{ו�U�p���z0��jP���Gz��Wi���U�r�/^��POlK0�6hl�)�6J�)]���C.���B'�(����Aϵ�/��jI����� 1�ڧ}P�֨e��̐�:ɫ{\�c�+st�Y����q�ҡ$�ޠ�nV3���%+��yl�yz�cBN_e�\�:R�)�Ѯ8�7�t��Z켏w-�|�ةZ��X��*�Ҿ�(�!nl;+ù�C�pi ��)�|��E$���,���O�D&��hV�)�vV<ZQ-��������_R*��V����I�;�kӿ��^6k
����^���B�|�iΗH�Q���Gm�N�]�ҝz(��,�Ӡ�Ղ�;���k]n<m,3��7=��d��:�ӥ�W��v5xU� ��n���۝��۬���j�VR������EYf58	���2<�v�(#˙�T�[�p�Z,0>�wԍ���+�I;2�m�YKK���:J��l1X���h���C����ٕT�yƱ]E���S�x�2r�ذZ]�	��]�&�� D���2�WDvѫ6AťT�����W�t��Z�/K�]|������z6�V:�m!��H𾒘�a�(�0�U�q}(���{R�[ϔ$�Ԕ�
��ިl��!�n[����p䠬mhJG�N��c7J�@o�#B:6�%kB� �"�p�;���8�z2�9��T-Sy'V�����(Ԛ���pԘ��,�ܭz�ۙ�0�:7۴�ߦF �pjՔ7+�\�����l-�K v�``	�����~�b�T"�Z.���d���Cr��e0J��ÿK���y�t]���s1&�<�T�9B0o܎6���_F�f^e��P���T�c&�����C�e�Wf>�P��3t�Z��_	t��R���*G��kA���먜�z��7�Xk!�I�u�Z���/���;3tr%$�4�:�W�`��LT���X;f֮�F���2��䞭�r��D�#�#����l"�Q�R�j[�B�_�Ҟ�Q��t�oQ��:ܭ�q@�^-�
���P�Vs9��� �k .�����He��\�%Y�zU0���@�ŭ۷����'w�n�i��ֆ�F�a���y���R���6*�YY\1m,�Ù��]��gp���p3�Mʷ:#�&��xWL�t�W�������'R��x≤QDT��A]T����fe�{��/��P�f��!*mҘ�ۈ]Hgu	278��gp=�,��*�ٍ�ū<�]v����H�Eghд�� =�bNWŌ�)�n�t����[���(����V+�,hI�c+zuLn����n*8ڏU�QTȠ�c���<��2�w ���\�lFK*����8f�VXݔ��7̮$�2����+�Z}L�PEY/yN9��70[��UvM�F!E;���̣�+m����`iސ�}ʙTQ��iuj�T��4�ˡ{ʜ���.�;�m>ǈSZ��y{ �hހRe�he�NV�epչ�I�j�� ��`�>j���7�U�U�K�*\������f�nՐV���<n$B����gTN�VV���S����9��w�`�z���VÊHҖf� oz�s�.�+:E��#� 	� '{XR㽋��
Nw�X`B��'�ب3TX�i�;��e"�fL��OǤ��I�J�/&�t����22�f�^h�EEݸV.�R�%��w��V2�+qbEN�ZԏUʻ��Є\�ܢ�͍i����-:΁_#��צ4X�fcz*�AW�A�S��Ur���,S��o7��������]1�==t"W]I��M#+��Փe���vɮ�O,_La�gOTrS�;�IU��ᕎ���7�Yu��<ˋ�V��"-V]t�-�۫`f��qD	�-����0�zI2�<���,-�6�����/q#�M�h ��=f�����9恤�q3�q�r�ֆ�a�)R�/L5�(h0ޖ������YZE�SP+j�x�7i'Hc�*����M��:����.�,�B�Q�������D��Nӭ�jnT�s�9�O�PpS��% ήm:Gr�r�����C|�IZ�]�Mz6�4z�,:�0�v׽���zE�;��\�b�著(]��K)���$n�
��H2�&�-]�G,2Ѻ��5�ꆥ����[ST�kY�l�\�`���w�Iq`�b�J�rz+�U�͖��F�n����N1:/�K�����
�N)�ʞ�H[�4e�+����6�m+���V�Lו�ή�\�8O����=�^����Ebj�k����wV@��s�s���9:�j�#Y{W�Cn�K�6t�&gR��Gn�����p$��D7X`�VmL��[������RUgM�ںH�h:�Z��۵+��9e��{(4����E���}a�(�2vWL+������u�����l �<���=�»��Le�Y�N�--�_SZf���L�,T���~Y}V�P�4
&��G|b�d���3���1)����'1u
�z8�����fv1�h=�b�]u;0M��z:�����sW�}�������\�G�d�i*;��p�2���U�*]�P>p�u�e��:�gU���9�v��^���:��s��pˬ.٠7!�[��gv���K	{h�t�
��5Ƹ���PQ�2��<#V��Ū�Pk�o	��R�5��	�Im;�o(�W�d5ha�}F�-�X�t�,�Fz:,L��ט��
fk��S�7zpg��u�(e��K�ff歘�Y5v�dTyB3�_��ꏲ��=Ǧ���c'B	 ��T.�+��i��n��Տ%go6>����JsO;<��I@ц��4=%$�j�C�ر�λ��Fq���U��}���:��ɰ�ۀض<��(,�Y6�Z��q��	�ܳ�Y��"�' ���j&vS���-@�p��d���X��jeO��+;���u��j�ls�t�2�VÅ�v���]v%E^ج�o]��c���M��
ѩ�8�b�=M���b*�νu�}Ef����y<�`t4�˺���b�)b�F#j�q�f��]��#�=���yYū7˱t�N��  ��>�M��ޢ7c��	$g%7x��Y�.]��]8�,Gؘ�T,�N��o+(7;���=����~!�w�����.��������@�k1kh]�O$�9͛��ʷ��J�ݺ�y)hz��a�L�n������p��T�q4I
�`ښM>	]�jVcld����)$�=F��c�ϰ�
�&%��v�m��;�7�<�ӬU�'l�j�:�fx������l�����롣r�fo]��	�.m7����T�s&��v��`��*hvF�κN3�����d<%�F���D�\ŗ-���k_4��d��J������o�qwX�����A�[NY[���R���Uf�W�I(�c��ܔ��fV-�e;�{� ����ի���7+�DE{����޸Ӳ�`�A��#v��K5lIk����V�)v�*Ś�v�kr�}̚��q��XRp��OsJ��䮬��	���:�ϯ_f�^�V�������a�xg�g縶Ձ�\������̴�s_g;����-)lc�;�d�k�����N�@T�krA�o��ԡǍN�Hp��kk@T���d*��u}yL�K��dq7���@�p�-��� ب��4q�fmM��,�k�f�7-���5��-�N����h�[����s;����vr�"��^V��)��N��ֆ.�
���5�F�_*��FSUw[J�- >Cue��;㶓�^}���6��E
u�8y��]Iӎf#J��cWh[@�Q^w������a�|�(����aR`Wi_�,�p������r�L�t� ��А]��l�ɴH���46��6kζ�*c�H�����4�����t����.s4$�G|a셪|�ܶ��t���[pt0s�*,��������IRV�;R�r}��ާ��;c�'2lo���C*P��wr�ѐ��'�K;Y���g �hݺs-�;�2��w%�:�Y� ���E6%w��S�xP��%��u}D�-{t5��;�G�`���1k�һ�N��12'P�6���X����m�[���^��=�:uw��_8�FŁM�Je)dɱ%���h��c�Rd�A0�0h� ��RђD�d�DcRb"��DT`�dj(�Ib���2!��2���P�h�H���Ԗ�0͍F34Db� �1Q�KJj"��Q�6$61A`рQ4lF(�D b$��X�5(Ƃ�fQ�XDDY*�&��c% ƂR0b����0 c�X�IF,A���QfL��3L(���Ō�l��b��PmIL��	��c+ c$I&�`�4b�A��`Ѵj#���# �4Ed��&K�{���_?�}�����Ӈk_Sˌa�qμ��[�8LΦ����K��{��!��j��a���3�^-��%֗�sW�l�|�j�]�*�ށ��b����-����i5]t���>�ք �S|Ϲ�d%��ܮ�<]�KwW��#냀���ƅ������ם�>�5a�})Ψ$�e�F�;C6��G]Y�S��E@�	�G�S>5�Z��e_q��[��N��rws"f3��P�F�iz�_��HxE�b�;;����*A�zQ#(��Z��XC�~����T��ɯ�3��%';eDV>��L� ��q��\w%Yƻ.��8�u��+�E�%�g������
��7����c�[}4>\��C�L���a~Ok��uF:Qy�����|���t��E}'y���e���A�����:��/RՀWH��eK��n��T�找������^�ΒtГ��2��$�ƽ�!$vr��G:zf(.����C@��`'q���*�C=ޭ`�1�'	�0-��T���j���Wd�<�/K�opj�7���<��_|�h[�
,����0.����|O �j�W��3��]v簼
Y�"&b(�zsK��P(t�MvI�yhLn&�R������(�Z����A�C(�b���>|sG��1�u���C��ٝ$:_T�r�����Y�t1�ʖw��z{�X����Zq��9H˩*�Z���ɱmK�NNf�g_oNBɓR�g�(�;�צ���ȶ��G}�cJ�q�e.���'�}�@��{u�q��Y�ֺ�W|�f�D'u�	��3����GF	m_�3z\n븜n���i�+1�V�5��nf��hb�)����ă�z�Q/�h%k�Dlrj�'.�"�8�D��g���0T,��ާ�����!R�,������;&'Ҷ����_u��yr�Y*��x����;�nvI��[����z �>�P��.�NK����؍��Z:L�9�r���|���?Q�^J/2��J��Y)�F�u�:��"�9��*<���>�0�ݼ�7��sCV�gf�-��i�����N��s�M��N�YGx�3�����!u�#V:VS��r��X�i�`�ӑU���~����7-�}��Q�[���/"��D`Fl�c��K�����0�b�=4 ��r�;mDE^�-g ���MGq��5v�]��n$z�Nw'��}\�N`5Џr�~QU�Ox�����E��x������e'َ�,�ɉ��$p*e�bf�͠lM3-�;�&�n�2��˽�P���WRdX���Յ[o`�GY=�V"⻸�Kf��]�۵8����b�1$a�����t�J�@�F2�´
\n�r���Ž��E�G;�;�w=��8+/�;33�ߨf���:�z���vh��j�Ck�5��k��N��^_�+s�7Z������>��4�J	`����n��[�V[|/�7C͟mFu87�"Xl7<�yZ��p�9�D5Y$�<mg�����ju�<תV��a��luT�s�d����ۏkT\8�8�j���SX��1\0$-ŉ]�T���*���xI���"�*aiک�]]x(wT��ҸR��z�3ٝl��^�W�+��	��(ף�T�!��R�&�<���*�E-}b��ݎ���z̋h������#�v��}U�T��ǂ|���LD"'�Jv�+K�`.4�W�6��9�;�+T3����9��������z`��I�D�z��P� ���[X9�j�
�^>�xR�Rܾw;��Cބ����ro���,��K�k"()�$>��Mo����+kxb���q�b�\o��!10:2��;��:0���"�Iٓa�]�B���I�(�Z�UMyM�Z+����v�H|r+����\Ǒ}�����Z�a�p6�*פ��C�V�q�OV�ޞ��Ӿ�v�3��#�����)TGkWjsQ����lb�.��7Oy�U��^�b�&+���96�Q3Cܰsz�TK� ����8�Tu�\���{���4{�A�Z��X�
7���7�;����3�ˈ%�=a���X�w�<F� ����l}R�0�t�����b�՗�p,-uՄ���TDEZ���c*�\L��7"��HT�ω��0w�9��|�����X�<�I�}s�!v(]'���҆������D�U�F��9i�+0Ei`��Ӑ�&t詞��}��0s��_Yո�n}�C���e��*1��6��|�`�4R�=�s:���}�lx�̔�\��yM��y�b��qx���n���;rA;�Sf���°��u��}.v�g�k}4���;��8#Kª2��=�Aw���+�*B.9O#�W[~��Q��mÝ�iO*�F{/�q�@U����+_���遳�]+�H+��bW��-z�ʀXl�B��CUO�K��څ�۾V[����rY�#ĕ@ρ�
G�ꄲ�R�����܇9ձ�{�䩛�$S�!�b�1��ߘ�O]r f�� �r�_
�9�Lv�W��Mv0]\re&/*R���M�r��ѓ���a�$9�P�V�]�B�5��h����뺂�&q} wW��X�%��,�7�Q�A��nNh���ȩp�eƔj�b�(F�W&����B�B=#���>�{ّoFڣ�ző�!�us��͝��:<Ц&vS!�i���x�b�S�FQ ����@z���*\�i{H�+9��򇗣�Z�;��j5�]���}��E��	����٘��J5�R`t�5����mNKӽ۽��ym�#�^��\�{h��(��,�#*�ׄ�*��ܺ�`�Te^�zf�C�)v_IN&B��J�l99Eq]�����ql���Q+����또2���*��Ub*!�r�$2�ڃ0��yB�un���&�,(;�[���.swe�:�v܋��oV�뎐�q�<qD����&6Q<#�N�p�z�n����;�d/m,ʰ�g+;:xoSgZ�́o��Ӌ�D:7ᆡ@�On�����@p:7���>[7N2D�Ë��p^v�K�YD�z�3~���R|��e5T'P���Apl��(�]~{jK"��$Ǧ��O{�������E^���y�+��q��nE]�p�M-��*��q�/|ŧ݆��*��:q;3������ ��W�b�y��T�R�م[��n�
.���}��Y��%tC�%U�(WR|o2:�F3X�z���|[�~{�f��5:3e��X�X\ELZ���@�&�t�sܒk���ok:�t�6�^�䙷�Ts���Y�����U����Q4�jfd�<���;nH�U�:-ʚs0�S��nC������A;W�q<kmTBC�a��F7&(-�ny_{��ky�)��/Wu(�z8e����J�	8]#�.����7Xk�.�:J䔂��c��W�e��o�S�س,c���S��Yz:��i}�'	� ���O���D��';��<�s(V�e�=[���e�cO�m����sl�AF�1	�3eL��������Ks�����w�>���yۯK.:.5�v��s�Ҭg�kθW@��"~����=7~������FL���J}9���宺:j��7��目�o�x��\�A�랙��<7wzV����f}�.�����b��y|h$��FF�rj�c�H���q�ѭL�ňK퉌%�����u�DD��F�vLH���ߨ�;Vu���(n�+[%�����~:pXr�7�@7���9/�;ŝ_*=�ú����b��Yώn���ɇ\�l7����Y^m�(��4Ss�C����,�;1�f��xE@B��C��	��onqT���1�3c��7u�ĉ�o>m߸L�fK�k8ryʧ5eWK��o� В*|t�	ڑطFԬ�]ح!b-��h���N�/:�wZ�9��yЍ��P��f��ag����I�.�X$$]Իj6�)��M�+�]�O<�9�uq��V.��ۿ!˯,,�����}>rh<�"v�N�͎>C?AWs��u��V�K�ez��{���BÑ^�u�����ɨq�S�O��<�=�U� ��G����%�S�3se��ݿ��!eHzj
9/ݶ�"�]����o�>r�y��c5�����Vz��k�A�W�t7��?�R��2�x����{Y�;:���-�:��(`�B���>�Қ���5��~Μ�(Qd�e�L�5�;C�S�F�\��vԺ:zf�ݹ}jv�_h�`�(�)�_;�8����mXAޫG���@h���5�n�<��E�����rj�[5�i�/�п>r��a��2�ۿm���*:Gkd��L\Σ^��m���׻�b�:K�D�S�Y"�q:q�å���v�Vg�����8�����᝶$�7J�\�J�}��GʻL�dt�>�ס�\׆E����sy%�>p�Ì��o��J�6�����rQ��ޟD��h�'�%}�K�鵳=�Rֿ>MC��̕���u��V�N���c��h����6�Sș۶IGZs/�A�	veju�J��ԯ@�kY��nl5�� d�*��������f�of�C-���e�Ǌ��6�6�n�۫�*���Y⩪��f�'AZ5�9u��p�%��p����Ɣe�:ta7� ��&���Q��$D]��a��Ԉ��Iе��*�a>o=��)p���.�Ź����^�A���E�7'���G�@J㢶�c�W�Ƹ�ԯ+���6;�>��c���cr:��2Z���i��4��ܸ���X�������"�a�]���s��|jH�$��7��v��y�0U�����M��f��+ع�xr�]�ӥ��Ī\�eϭW{�}�}ܮ�X�B���)@7�G����̫�6筚�o6�~^'��n���r�3��,��C�Ք-uR����[1?zU��ޠ������Lrżi���6���a�u����X�.�qw��E���Dՠ�a�]�uwCf`r���S���u�"��lÀ���χ]z�L�7����v�\�n�}�3�3�!�
@�ؕ��T�2�ب�z�W���b�5a��7+�\J�gb9H�N����_�Ԕg/��C������*+����34'z��i�:\53Ъf�J�Tu�%nc@��\�2����m�����<�l%��u�œ�12:"�>��[�|P���˫�e����KC�)Dt�9}{|��Z#VP�9���P�gY_��usR�$g^���c��i��N�����u�e,ӓ-�)����9�ݔEl�q���O)P�ވ4z+�
�
��G�΅u���rp���X"b�7��5�3�6Hi[ZeC@V/���*����r�gºt�ug��w�Ы��x&���8������l����=5:;`\�5t��G����{;.Ĳ%l�UTA��y�ё=+7��e�%��:�Zq���n�ޠ��@��UHV��\�j픝����1��t,/�+K���d8�7]�k��!~i�|H"���í =@F�Qj���ƭn��VT�.4����Jv��Z0ȸ���N홋�(��gp�}=,nG$�U�X`k��&Nj�]0��;����hp��WYG#*�׆�8��S����yZ����[��Kʓ���=d�rP�����P�.Vaņz��R�sZd��ɼt��{gm�=5l�L�U���q�� G�����k6�5�[RyZò�+g�̭�]�fU ����5~.Ϣ@�d�>ZcB�u�onW��ll�(u�G�����?���g,%��]ɟ\Ns������]��;�Q"̃������
�j�*��K�<V5���k�) u;U���>c��l[�&77�]ntf�.;ٴeJM@�����gC��׌i��n�i��W �]۲ٯ/ZR����W��7O����\�!Ѱ0�(a=����g 8n\u�O�dHw�2ׄfOf�x\�u�T�S��<poKf�u�����LV��5v'���Ј�6v"��̸n	m��P���r�mA��F#����7>�zՇ	�+ʜGp%Wؕ�>�8%�z��m�#����!��Wim�{O�Ӊٔ_0< ��-�������\*�G�g��z�'�:�;q���2�f}T\s�B�}S���=��B�	�E	�_e����"ǒ�2VZ����������E�8n���S���t8Ү���c:�I:hI�hʯPC�CHB
6�n=����w�_/"=<+^�7��u��&E�T�sҲ��$b;��� C�
�DX��ȵϺ��q.+)��)=����sV��RY|pi�-��.
�E{�|� h���@��{�T-,�v�TC��j�X��L�s����ȿ5��;�sTc>��(
�OH���x�36x;}x��wBp�����P4���	�ӝ@�-u�ђڿ8�.1��$W����@���X�ǡ�9ȳP�4�����m>9�·�[q�\����9�=�����Ss"�l�����i�c�sr]����j�����I�,�i����g�յ�NR<�-p��m�[�ԅ
V�\1nb����b��ݺd_��y(�Q�ז�k0a|
ySt�w����Z���r�:̅&-�z�v�я5������y�G;)�"�DZ�[��"%��0�0�Q�O�Z`�e�/l�!R�u�[���n-�ź*j�?D+#��7�d�FZ�j�>˺����O0�6H��֔���]�V��f��6�n�3�o�j�܊
V�I�㕑������\f�B��e�f�1]��(�Ը�r�;��&t�J�L#o��%�6 h(3����t;*�r��aY�/����w��wS��q5�|�%v6u��O<�:TJ��a�C?@�E��媷/�ΘAk+7i_
�/C�H�U��2Pyx+AU"���K/�2��[�|���T�؅t�V�e��[�
9&T�����FTB�Ë��x�`�X�>(E�j�<W��O��𸢖�}��H0�"�5U��j��Qt�h9�SΊ�v3z��`��'kp��� �d�/��4+��]k����"Ñ<��d����F5�gA3V��*�cye�+p�`��y6n��-�f���]���<�t̓&��R@5� B벖Բ�q��;�̡���cu�I�m�Fål�d��A+>��,/Rͨ��t&�<Hs�60��9���{��R7�#�_:�[��5H:R���0M� �gu�\֎I���RQ�T��$<{c�u �<9ŧ�:���lΒ�T��VA�tu�i��\쩧t��z�ɑټ���WL��%�w��H8��I��g�=�9�<�Z�>�7d�3�`+:�X1�	;泷��xd&�.���*�]m��^ILH��WL��uv�rN=�?vBn��¶�g���%�{)#$��X�k�BӊS5����+T�_Lֻ�ч:e'hJd
tg[���KMGI�Ȍ�6��ݗڪL��@�ӄ�!k�N1� �������(j�L�û�k�X�M��,GM̎^���f��1ER�B��Wf��R�k2�$�X���Ȭ�:����H�S�)bU�5+����I��u�ع�rMs\��;w@U�aXT�;;��[�i��ٰ_A��K��pΣ��v�t��M��M�V�,d�X2_)Og�Ƈ@���*اi��t��Y�|�Y�4Q��rk�-����6k���E�����_b��ĵ=̛c�j.Ð�Dg8�)4���7Z�=�l�6Mͥ]�j.��P�o:�;Q�/]��1R��5Z��|��#�,����[[���L�ysE*] ������[,]^�\���زp�[�=�T�8�C%�zĽ�d���:��I��eL�P�	,����]�_��]�uw��]��cAF��b�"J�#Bh��b"(�H,Y����1i��6��L�X�J�dL�h�X�����!&�fd��RRh��TEcFƤ�`&IEEIDjA�L�hH�"�Q��F��͑��Q��F(ƣ&�1D�ZJe��dj(�#F0&�hK%�&��$�1a$ŦlF�dДQ�X�,�[�@cIF�2XM�12(�"�BXLLK)4X�H����`f	�ə�ɣQ�	ci��L��Y,$�V6,�5&��D�4��&�u��������z��rTb�-'��e�V�[{��L��ղP�&�kwf�K�G�!����2)-����޻g�SXj|��篾��������_˯�޹ֽ?+���o��H�/��nＮ�͍����[��6�t�t������+�|��t/����|���W����m�Ͼ�7qW��	�^�8���~{?O�1�������ھ���t-�s�[�|W[t��}���^���9����������i�-��}\�y�+�ˮ_ͻ떸���W�^��.����x����W����#� ������e#"mZU��r�x{��\Wŧ�W�߽wc��M�~���}mι�-���z[��mϼ��y�U��.7w��O^r��z��v���mM��[��t�-�/�v5�x���d/v$}�nn�։��ߗM�]�J��K����vߕ��o~y����kA�~~���J�W�ϝw�-�].��t�y���/Mq�/�ϗ?uoKzW�����ͺ]-�w}�kO9�o����DB`}5�[��}}�M�z;����߿{���q�mżv�|��ۡ����ݿ7��ߕ�|�7_�m��o�My��[���o�����m{}WKG�u��v����mל��n����W��ok���{�>���`I��uص0{��K#3�c \D�d�
 ��Q�9v7��U��]\�6��6��z��~W��n�B��?��kx�?6�u�뻯|���۞����m��|Z7���۾r�Θ����U��[��_߮���ӏ�������>{�]z�߿^]7����\/k�]����W�9n���]/�s���o�|��O�|WKO9{�\�X���t�W:�]7�����sz[�q�۟o߽zj-�DyMW�18c�#�MfM	ޫN�V�g���/6.�e�#�>��C����������o�;��^��|nץڻ[��o��+��_����֍�7O]r��+��n��t��qo������+����.w�W��q�/=�=�
�]�ƌ�=�ݐ�k>q�\L `�O�v�yͿ.����}b��<m�w������*��/w�:��zo��׺�Ϫ��6�z�˥�7N���|��5v�-��z���/KF���r��5��j����� �������-H"<#�"C�{�]�͍���uםۧ��.�z���}�ͺ��}o��ν���<���W�qi����y�{��m��ϫ��n���=r����n�B��6�o���k|����)x=��E��%�֝��Q�/�;�xm'�}�hf�p�p
u��P�7Ky[�������ن��#2�i�4��'��_Z۝75�n��Y}-ly���w�� ���3Is��U�� �P�%	�f]	E�t�3H�p�WSfz�N��S���8�x�Ǉ�n���˵��_�w�[�Lo�?�۵��}O�w^���뚽�wѸ�k���O{��v�/�t�_?{���kE7���q���>���Ik}���0#��{�^i���=��c�1���q�c{Ux�W\�m�������n�V��}�Wmn���u����u��o�{ldxD ���	����6����O)���b���~Q�(`xD���+��nr�+���]sv���\i�__[t�J���/�v���^����KN��������[qW�Ͼz뽿7�b>�S���g��D|7s}���*���2}�����ӥ���_���-q�[㧭�Ϋ�~^֍���+����ޮr�������s�����]��-��ۥҽ��t�sn��>\��h�[s�滏�DxG�,��窼�=R���1����mƼ���}m����?uz[�q��K�?wk���>/_��^�<�7m�y��m��گU��M���-�;��E��~�眯M�۝r��r�o�]b>�퍢�b���qƱ��wn2-������u�zZ+�o�]6��}n�r���~m�?uW��{mι^~��ok+�����z��\[���]��t��Z�����n�Kx���\�h>#��K����+��9�z��8GMv��wΖ��.��n|�����}W��^����KF�W��>�����]5{�~뵾��~W?r���ߕ���}�uֽ*����9�^�6�n��^u^�	}�$}\=���i��G�:����/��+�9�/M�z��uw6��n�q��5�\�;7M��u�kx�Ζ�����z떸ߖ�u��}5�]-�<����];WJ�~�ջTE/�w�u����g�*�~m�{��}B�}.�t�_Uq����|�j�h������[ںZz��ﭽ��|׋����M�{��Z-��m�ﮯKE�W�y����~�k��ny����6��v��>��nj��֩�t��Q�x�=10>��OkE����}���ݶ�\�W�[��t�K��\���Ѿ��{��W���z���n�����z�ֻ�ŏ��_?��{U�q��s����t��q�{��_�|��n��m�ɍ����J�!�xn �Of{��Y�d�Y�%�%4���(�]�2���5�%�ч��G�c�R.ѪF��.��fצk\2��׶;l.j ��XݰGF����EnAy+�F&KH��^X�(�-��m�d�F֟:Z\,ڗj��)�����j-�������oνr�u���zm��n���~�tѻm�}��{^��|W�t�W��s�{�7���./�.֍�����7��]6�׮�c��D}� �v����n)���C�>��������������ƾw�}���n��}�j�����������^��s�{��|^�����/k��M��ׯ�]��\�|n�]u���on���]|�2S`���^��z�}��4}>�>��z��Ƽ]5��t�u��]����?ux�KO�����v���t�K���V��߹�_y{�~�W������^��o��W�r{��C|m�Wު��]6���d�z �9�W[���D}" �>��1��j-��w��ͽ.�r��u}m�����_.���m�ns�����]��U��:[��WM�nu�����x�k��|�w����o������|W��i���?|���w�u��z�z�x�ǆ@��C ����]s]�������]w��ۥ�W��u��j7��]o�q����ܮ���_�������hѸۏ^u�/��_�������kx�.�����~�����Ω��ϔg�Ý�ϼ��p@��S�}]-��}W��ݷ��Mpk���ϛ�b��[�ﮮ�[zU��{�\�k����M{��J�_���6�y���k{W�q����/M��;�:y�y����~�{���ߵ����q�7���W���~�����E�7���Z��_yk����k۶�oM�y��}k��]<o]s��؋���/��i�5��˦�x�O��}���ѻ�ͺ��~u�����z���Ϗﾮ�yo��h/ۯ�����[�[��W}r�ۡ����~�������Ξ�~�����+������z�~��t�ۥל���ns�>����*�m�r����lZ9�����u�_|����{�W�Mm���D	�l{�}ז<{�8�W��wo��z^���z�����W���v7��������w�W>�_�~�oj�\o�����׾ot����m�nu�>����D�#�O�k���LY��ׯ?�������n6��_�9~}zhѸ����o����p{��U��������v�����U�w����~W���㮷�7m��WK����k�ן��]��=�:���2>�z`P��e9]�q�_���ls�Y(gZT�j�]W�b���X�1�*.���Hwji��7oq��\�NnT;��RO�Bb���wͦ����Nw�	{$�GH%1���^V�z��zBG,4=�p��M�o
���"J�gݵ�w�.&�gVpݺ)'���&:=�|>>��]-���/���W{����~m�vޛq��6�w6��o���[��6�����}��~���y�\_/���o��.���]h��t�On����Ý}�=��ik���z��#� �鈡"=-;��y��o���^�sv�Z7�����-�]-7}u6��[�t޵�u�/����_��J�\_�{�}�m�n-�\{��}�oK���}�}����_�fAח�k8*	��22=�(�������6���9ţzm�r�_��h+����o:�t���s���k����^������hޮ���ץ���t�mpo�q�����W����,z���^��������=y{���׿��ޕ{\o�>��~��6�o|��q�<�~���k~W:�Ϝ�]���_��_��4h�Wy�[��t��z��CQo��z�r��~�k��)���=8"���Fy\S�����s�G<_��0^T�f����@*7�����hW3xa�&��*�w���|�����o/��Ǫѭ{�9��T>>��<"���k+Z��'c4�"��o��լَ����Y"`(�9
NI�D�d�l���k��V�8��J�7��7r����ӱB�������'1�W�v�*�!^��B���	B� �m_A��;�y�Z�\��cOU6���v�#�,�� ��i��=Dx�3�yA�t8<smTBXuT8�o��Zg��v:���C�ܹ0�N�<�\s;
1���.Ɔ3��9H�+�Α�i�����G���S4���2�]�u|K.*g_�[��2��:|����~��)�I��(�ht�%��#�Ɍ�n���irwO�&X�u������w�Z/`�x�5v!u|̏0�>!�a�qS�rtl�ӻZ����'mK'O�^���]�nA����Ô�# 8V��L��8�V_B�8H���'k�*#Q���b��E����R�����"�kÚ�����O�m}aE���~��^i@}9����k3ܮ, (�P+��u�\��?J(`��b�㚤1Ɩz�S�c[B��tT��%��>�`&"���"7��b�b�O>���T
Z룣��~qZ\`��^"�тT��V�6a��^�J��1(�"��.����z�Dl<�ƂK�Ddw��%(	<�ͅĩNg���.L���>qp���lE�n���<|��vLO����L��ttT^����q�fX̆���C�%6Ҡɠۮ��C�S��ꜗ΁�ί�-�R��^zwWe:�%q�/�WI���MQ�Y+ĳ+���Ǜ>�P��Uq�V�O�Y�
����..6�*VP����aa[WC�����}>rk�%����l�R�̪���fR��3��DF�!�D����W*�E��P��p�ڧ�3S��娨y��S�x;"�6aWN���c�����qG�`4�yt�XVUթѶ����!"17�M�aGlR�'v*� e��E�,�v�z�;�0���̫-�զE��������=p�Z/��Y닜�*�4_T����u��XX����i8�g�UWԎ�U�'�~�?	���Y��@��3�e��q���X<l����u�ފ]p���9�s��UT���wT���w�>컩����ݳ!a��x��$�N��R�N�o��/;�����߾�!k'm{� �غoͪ�涺/:rH�(�z2��V]��|@ ���r5~�+�;'F϶��P��%�)�_k��a�@ݿq���LX� 
��qT�S�������#|�����*�<�4�}�_>�U�nS+���*/�])�zq�]Z�TooP9�颎;D ��x:K_E�n�ҜY"�k��5�J2B8r.;c�9�NgWoh�m��wB�f����q!$�p{�� �����K�����,`�*��l�:z��3[�[�,��Q�p�n݇�.K4xoI��BR�@OJ�~�_)��N�x��K���+��?K��>;�Ҏ&�9A�G�#�֐B�W��0+1N��΍�C���LI���[�^���E�p(��m7{n��M2J��T�Ӆ'��O`���[;d��;Q���~�*�6}y�/ �E�N�<x��Vb;C)��<��9�p��B��%���U��tc��� H��S��HH��gZ��.��;3'tx�.�wa
+
z��p��l��6 gS�Xq�$�n�h*$�_P=��W�_|{�z�^��۰g�"�ؿ�X�2��mI��4 ��J�>�o�˖�ݪ��{�d�a���{G�&��5�t�W�z;��Z{��hƤ�I;2[ c�3ٺ�m�޺Y���k��a���Ip������]C ��Ր�8�(I�T�1�v^��P���S2�S��yU/�͠]Z�8�Z��Af����g]z*���*�}�mauԼ�yvlv�����<_�!�k;ʘl�
����;�Q�u���P�<(�BL1b�Kwg��$P�9�}콴!Y9�HB�j��`tTDx����N��;���gS{v�E�[U��S)��iGcV*��Y;�[j���xߠ]��[��%��ʌ\�`o�`���ko���6!~cگ㋀�X]R�՜x�WI�=v�d8Bw�U�����ܢ�5��.,AңL�*a�&��W��J�V�%�Zj�,���{�Y�]t>�"��]�(ز"6O�(�|'�-�>�
��N�W���^+�o����{DL�Luib�x�l'u/���s��`�7h��I��X�����M����j�\grJ��Ք��x��5��\+�ooqnwk�hLf������	.!Ȭ������e��Ħ��r�jwcaaڧ[&N�D�w�Xwr�_x =�����0�n^\|�Hq�1�C�N��ګ��(�u$�|��
`�z����2�����'��Q�O5%��1�B�x��m�w�`A�V�]ۙ�:��{!��1Smr�����K�p+��\q[V*�2�ۙ;N'0+]Ozs��.r@��	��a�>+7r5��bf#dF�zs=G��ޮ��N�# ��G<\��	��;9Tˊ�i^z��f�d�J�G�ֈ�c��jb>U�r���r��=�/�Z���W�.�S��:d�Į�6JcЫ�}ҨMq�'A#����l93�N�W��B�$	��t�X�������*D�"�� Eܪ"t�9@�����魌����I��.�:���x:��c�q���7�."Rr�4��$ŏ3�^'h}�lڃ���5��Hx��u\��T��v���=�q�#"��s��o��3*�+'{$=��+��Z����3���������ǭ�<szS7�n�eHxE�b�����=)`�"g�!��x�n����H�w[�S��~n�zz�~�ܷz�0��f�:ҍ�q2KK¹�֧zz�᎚�s�O7s5�ʾȩe���-��y�[ޯ-@�pV�wmm����@�|�Y�Q������U@��eV���ތxsB:G6�R��Ӷ����sؒ��Ph�yH�#��FNC��}������W�`q��+�S��ys �Kл����ah���a��5+.��+�vʮ
�{O�vB��}B� �o��'�Ǽ���L����N�8ƍ�[�S:�:u�ҞOFm��d�t���Ɏ�������)t���A%x3;Cݲ�Nˋ������b��7=��xWO7��G�v�C$XI�F��\����g6���MQ�P��H,i �]��,9�ӑ�<�A2�N7�2�U�u� ?ư.o ��}��/[}���U~����C����{��k�����RʍT�*�^r�]l�TE��*�uX>*:$�B��]�뮪L�^�r�!�t��sU����Hc.Me��CU�Ώc���
�T�48��b����O>��2�W�����m_��VN��cJ�4��gQȶ�wx����(�>���z B��D�:�E;�5�u����=SvQs:M���Ǯ йr��*�����\�`�ғ4|iV���8�=���|"&���j�ݨ2-&x[���V�ap���2ZV�%d�ݣPN��
|4�K]�Gi�X���&�%a|e��uk/m����H��kF�G1��,;�%�!�wi2����6��˷��	ܽMU͘�!�lO�*�Yj��K������{� Y�+FS��I��W��xTe�T"j!%Z
�@T�/�@����U@w���M\����+ڬ/�9�]^gv�*�[;F��/�������S&���Dsf/zE�i�jB���O�#cu�Ǒ��$qR��p(B��U=���Ŷ���������N��O��y,D��9y�
�s�Uo2�,��YVex��U�V9ѯY����j^.���{����;V	a�w�����VEz���Qi���Kqp���aY���{��{��Oz����
�����l4e�~�O��jj;�{��?�F���n򊮲������el�b��ޗ��D�#�"���1<�6Nyϱt�j���ќnH�d�_zea5�g��R�7��:�Z;��G�j�f�����!D2�Д�/�לrs�7g�W��[.���C���t�kt�,��f�M��yګ6y�i�b�X�J
"V{��e`v����VM�݊ҥ#9h���Tq�MVI(�AB8W�z�/�wN��"bw���(��8I�;��T��+:�a�u�d�����#�Ԧ]L�-Uo7ѣ��	uŃ/Vr���bm��Nl�W��9���J���l\fQARz�����qMW��N�Pqa�(�K�؇���2���ŸtǛ�_�3��Z*`S"D�!���[ClX�����wO�!��:���pn�M��Җ*Մ�Vj�x��[�-ۛ5*;$a�X*2�
IJ���ȸ���'Z�xe�V�y�u�g���1����Hvn��Y�9�^d
�üv�FumDOm(���2�sww|�j.�E]�J�#�<��`�3	zM4���|��	-R��ժ�JP���NChn@m�9+9x�[�Sb�eJ������J��XQ�9Z�\�a�U�+a,:��o%L�i�N��(��7S��7���-���x�Q����I�յ<��z�tUx�3F �	�ѫ)��`�ѯ(Z
�E�{��2��ɧ]]���ng@`Q����F-q���� ��8�sS�|&:�7l M�v��.9��Z�a���c2�����Gd��&ਂ'Τ����Flؒ�R5����#���j&2��.n�.�R}n�J��qzt�veeɊ[��sy��\��v#�zLF�W=�嗘��������D��V�y:�NW�'���a@�pR���J�JU�)⽩����D�ҧp]1���-�+�\�ٝc6T��<���xq���C�9�{.u��F�\������0�Xc�vZQ�W%K�żn�Aɡ��5Se��K��F�ɣ�����q�����+�����^��sU%�����-`8x�yE��V}�E�˕�*q����_s�S��S7��ɡ�,-d�4)g#0���Fg7��K뛽$CC���Be�����[��8b׏�ܗ���|V@{�P��lh�vAMVeB]�tZ���I#F��t�K��Q� `��ǳ@��p� :��bt⩇;�3�"��E-:)䊻�*�0Z���>}|_f��}F�t,�;���Τ�L�!W�Պ ��/v�d2������	���גq����=v���<�f]ɠt�Z�MY]H�r�C<�9�m�P']*�yd�����8�{[rt�!��=�'�W@���m^�hy�<K:9����/oL�oAb%�V|�M
�5ѡT���-wZn�մ�F�WW�z�V]�}h�"�����D��qےV��.�<��	踊���ƨ�#gi��V���b��K�}|+NWJ�luᖩGy�n駶��u�l8SNu_@�l��Ӥ��]]`���ǫ�!��GJ��&��~3'n���V{�h0(`&�|������9���jX�ŉ�����s���Z�f�V�i��nK���M4	��7J�f�,w��]�e�4,Z�h�E�a �#��;����
�1��i6��e켚�[d�慅D��{��la0�Dh�Y���QR`�Kd����#X�Ff(Ѩ#T)��4m���Q�E��������F�%�l�$�*)6�QELŢ�"��B�D�*�Ehō�X�U��H���EL�bMA�d-���5*��e��cQ5cF���b*�1�љ���l&�F�,m��J�E���F�AX�[E%��j�*,h+%��ecX��L1j�cm�QFţ1�o���������~]}{��^�l�Ի�1�%dޜ���2���ĨV�oLvge���C�6
[���U4�&��sɖZ���ޯW�^[R���=F�5��Mc>�D�8I�W �t�ϕv�mR�t��ý�V�,jHNJ���Cm&Fszˎ���t�,ף�zL�"AJ��'�X�
�*.�#��az��k�U�N�E�7O��t����DFS���)^�_
��*p��m���ۚ�"nLƼ�W�rt���rg��{�v��)>H��~+oz®���v�Q��" 4\Jӑ��S6#z�	u�-��2m�5�L5]�+N��>�z��\�a��p�!p��J�BE7�7x�)!�2awr�'��pFM�X{g�*q<�F��g��48�z�'�@AvA]"�����hw]�FV��-�c�ǺY��܄^��T1	����	u�UJ�͠]Z�8Ū݁f�W��a�*�Vp�����0��)��<&���HE�*թ�
rn9LPu�4)�Vx��x��uۂ���PL�o��x3���L"�T�6����>��xMʜ�{��;a�ntXy ��?��J쾠�ГW�젺u�[(���+1>��6:�AʙJ:,a�X��wz�t;�. U$M.�q�ۗ�1��fX����~�
����v�x�zK6��Xkh>�{Y�����ޡ�,��D�-YQ�M��a;����R�ej����oi0��;�Î
*��S�W�U���l=�}��M��9=
�YU��L�J8��Շ�*��Y"c��j��Nq�w8z[kr=O��h�~��������'����-���;��7�AַOP�HW+3a&s�fAzڎ;�*�w���7A�V��$�=#��ɠ�k�D=�s����������5��]�kG�xk�m�2�����in�A��\d2����Z�����@���c��/D=�'~zl*��B�EF�R �����V�ʐP����Kg+�[�i��]�f��Ϩ��h�F+�����2{�}�'� jGf�i�M���~i��7��W2�^U&����J�T�!�y#6Ҳ<�k�M��Ǫ��tT�kv1g����}�3�/È\ioWGd�m�El�a�n�7a^ķ����S�r�x�^��>O$x��h����A�L[�^+J��z=�˭!��d^��,aH�Qd��x)��*���*N�G=��"�'aɡ�+���P�xfތ�!֌ّث�m��m�y�Y[��D�'��Qw��n��|MFQ����=�G����D���Ne��2��N*�t���{n��e�g�y^^ԃ��xo�w��֍�0��^�mIC+t��LX)pܥ��BJ�&�"����� ��q|�f�j�c�=G��J���Q _w�V�'.�C���t�]�ƕ���r��H�[��=��ԷA��nÁAs�C���M����zMG� �X��流.����Sw����ٹ}J�ٗn��]1����@s<�V�y���K�5������A{���(�*5���q�]O��zS63�߯�HxE����]��̋&z�����n�#,�E��^E2C���RrO��<Y9`v҈�jÄR�#ČK}�Ֆ>1�tvFX}ٶ���N+��*Č���<�'d.@xe ��K"73�y̺kd<��Pa�R瞌�L��ۦ�{]�3Ǭ�R��'`*���:y;<�{w���
O|5�¥YL��-�n{C�p�:�������a�8�m}�xe7L�}�M�e��x>kg�E�@b4�]��Ξ��l/��r��w�e�,������Y�.yɣ΍��3T����I�J���^��^>��Ƹ�TMj��RYر��2����|�s��1q��v��廮�K���pގ�RS��
��_
Cs��媲�'Y�vk:9:U��D4L��em�Nv��̓��ʋ�8���p�8�^��G8W:�w�'�l��}J�+���WT
��^�>P�����}��V��.?L�a1߁�:k���~%#gA�Wt�u�\��V��@9qёa�v�e�zf�����)f(�m�ǲ��J88��b��$�f�L����V��T���ݜ}S�H�T������?3h��N���n��ti�(�{�]B'I<�ߨ���gdLM��B�8s�����]���MR��D���'Su��ؚ��#�����M��WH����<_-��;V;��(.QClr�ɦ�t�C~ h�L��U�r_{|Fל,���|��if��u�WR��7�+��'��MP0��M��jp�]FSG?*��ou�:"I-HӓT��UOa�zqm����Ziu兜����ɋ�ݫ���ӳׅ�L�m^?}�A���"#�.B�FB���W��i"�l�w�`��F�_RpI� �}=��������(���mr*͚�n ~b ٪3� A�!]Hzj
9"zF���
ylҸ�Q���u���lr��F55�W�ߵ�d�3�6FW!~�����Щ��=2��W>���;Y�1pKY����%3h�̨7F>S���Ԅ7:_���w��||krZ��+m��S��Q�g[���W�7���ex��p5�lny���ᢶWf�@X�ʻ�tY�B�;�/VQ��DXl�9E*�e��� x*�n��"��fW�DH�}f,O:�ϭl��U�,s�返ǂ�G����&d��{��ҕ��t��������� 4o�e�VK,��2����:�N�̵��v��23jk�g������h��h�J����������UE���J���a�L�~t�!�<Vp��c���^��E�@,��A�W �
��K^��?>W֩�}���5�w��Lo�kA��(�n_9^MX}�k��*��'�ʈ����쮀�v�Ƶ���=eED����Z���R�"�[M��1���A��۰�DGŏ�4����'yf��������m���c��q0#k�+�_X���t[���9N�'�� �)��j:d��Ѥ�7T5]�*)Y���	j�5i �}W��/2LƖ�W�rt��3�8^�A�w����wg:�كU�o�I�n����GDW�{���y��gvҒ�Cg.����zz��Q*bfvgK[~r0=Z��tTp��o��a�!��C��(�Zlw:0�5$=��p{��ez�`�ʘe��ʂۻ�s�#��ǭtV��Zu��6a��v9Y��]���rL`>.%����5�����Kǒ��+4u��CӅ��:Q$����S�\�VI��p���L�{Ǐj�C��E�k�PDu��kz�r�>�� �ɵ��tV<��#B���I���#'�^��(t�6���jֈ��o)hi��֮tgZ������@LÙ��Mʩg�@�^'U�>0�ו�̧�9�6�u��X��;��E����*vy�<��,S���[#B��x�`�&^\gP��B��Q;I����uo5# dX�͌��q�a�<��h�'��g�5,�e&�7�3߫���`5�7Z�0QĻ4vr�Ui���J8��Ն��2�`EF��W�<�n�
�
��i��՗޲�vc''��(y�K�u�^fĢ��jxﰺ����=�̍�]�\�S/�v�4<}����O@ݿ%z��� � 8�eE�:T`����B(i�kk���Ctܱ��xJǛ�
gn�څN��L�u���#+����Yg��Ek�)��P��n!�5�Ў��;���K��&�/����H!ůc���מ򫮄(�u$�|8rz����֪�ԣ�ڱbD\��)�]�f�ϫ�*xq�,��c�������I����Fy����׭�}��t��ͶT/q��u��9�ޅV��ſK9A�;F0,۴�=���'{}^/<�A�~p{.��L��u^xnm�㫸f*�{�ޥk�-�hЊ����'�qpY��v��^���f%L��[6���fo*���(,t�/�z���ӹ�*���#2~���@�@�v�U��
ڱV&\ws!�i����nȾR�P�}�l^�y��[���E{�i�bJ} �z�!q[�ѽ�N�# �{-,Xw]�g&yw�v�@~�tnU>��I�ȑY�	��%>U�r����}�xlj�[%�jr����r2n6J�,1����T�\eI��L�v"{�;MQ\D��t�*\��Jʜ�Q���c%f[=GԒ�K�r�9���|Q;B��`���+�m-w����/:1��G�T��E�+uz��r�7( �"��Z:hz�*ϢzY=}�i8(0i���o�sp��l=AӲ��xn���®�ۿQ���@�On�v�L��,�o)ɖ��Ғ�U�
�Z6|-}�/�v�F��s�׸��LV��Sb�aSy�.s�xɫd�/�OVOVu�6
6�<�(cBʜ��<Y9`v҈�jÍ�˴S�M�kcxn�j�/a*����b�{��ma�q�.�U�
��
d.@x8���U��;��\T��*E�]��[�.�0D�p�t����zz�]�*��GrU����6�"�9	�h�An�v�Τ�Uy%�����l�����3@	��+F^YBT�r��wǶ<y���e��3�㙸�8V��)M����nW�{�xy��̊�����E�;ܽ�S<��R���ǢVm��T>'�U����ͧ^x�zU�)]e%:L�B���S/n�Usv�[&+�g��w. WC��+/�eLm$�հ����9Z*v^�Ӗ��`�תH|h!,��v�ONF�p���L��t�ƕuЮb�
���i>�,ED��s� +���;��JIG�;"8�����[�5%��4�>�ިC2�������k7*8/��½ �j:'�x	�������ٞEӟKˎ���̩���Y�뷈r��{��1�_�\{+��(I(��b7�Q@yU]��N�Uޕ¼����"�f��i\+�#��U���q���o�xأL���D]�'I�<��z"d뚵B֪���u��'���]b#o.���~Bƒ�*�.����b`������+�zrj2r�"å�:���_�P\��߹Pd�m�Aaˀ0lq��x�d����W�B+<.Uwte�Z�L��0�����������;�+�O+�TR�L�)���wc&2�D���%ܣuR���^��|c�~���wu�mٓ\�Ŏ���J0�2���-�����52��[*g�|鹱XN⇼�ӥN*L�2�#.*K
�������n�ev�@L�{��]|a�����wV��M`��m>��G�c�&����z!NA�� ���[Io55U�o�/�\��*����g�_��:kl���O	�ai]WAh�����u�^Oi�C������{$�r�N߇+�68�3�����"��X�^������p��"���"NU�՗��[`ھ��WOm�G�>yf�D�?1 l�3��	
��0�C-ӳR穄����9�Y�,o��]�^�-g �*|�`jj;��^ʩ���K'v����� -[�>Ҕ�{v������@��'��!�E��1��t%U{>]0�ݲ��<�Y�Lx+6�ř�Ü���u��%E9��@�
��#~�6���&�S̾ח�
��ٹ����u��;̴�m���rv�$�=X:}M/j�[9�i�/�оj���8;�2���V+�Xs�?�hx}\tQ��x�8�U�\�k�2G����T���F�+ch��{��1�A���ǘB����v�V`*���X�0���<��H����:c��R��}��S�T�:�J�+�]���s֮��h��1����b�g@���eu_��V�<������C��t���_\5fj����L�c�c��{J`����u�3k^GX�S���	LQ�/y�f��r�;tk�C[y�K��3"������g<�8����u��]��%�I�n��K�S��$�(�Vt�Rե���j*î��1�Tg�=����d����[��OqY�����W-��7O�M���faD�Gf�~�p�`�!�:qt�v�{꺤�z���&�Kz+���E�p(��m7{�S�Ί��R�"��V���I�Ol� ��;���n>����[���v�p[��f��]n�+��K���S�DW��&+��0H�ՑR�8�:��v��~Ό9aS�59�؍	��Ɍ�8>��Mٓa9Z�4�2O{�'�2}� �"����bT�5>��Ֆ{p�O';�M�wa+21�]���+�9�R(s��8��v��7���q̉�2-���^�����&����z�l^�ᩗc�F�9Z�ySdhS�<M��s�~ݖl��-r��Y�A]e4l��2/�S63/mY9�HB��]A�_����M�?�TS5����B�`�� ���P�VUi�S<�G��Ն��2�qQ��b]�;&lN���1�1�3g�ӭ�(T��:�F͓�]��|��/����D%����"�m�KQȽ�qx����:2�T���-W�OS�Ns��<Q�|Q�f`���JmS��qp���v��\ʙ,��`\��T����΍�������;BcS��1	�>.�km�l�N>���
���U�;�h��[P�W�d�q�%���R$#2�uJ���x�ϐ��pd2�&e��+�a��|�u	}m��t�B���d��e���Z)�*Dk�l���m���+-�8au�i揑s��{����\59S똶���ح��G5i_j����<rM��P�j��w)bi6�����}��Іj��z�h��� @_@���� 0v����f��B���k�_Q;��W|U����ݩOR�/K#{oXU��A���5P�0!����w(b2�i�yq�\+�ww��k�u��p�n5Y.��٘�N਎�Z���v�Y�Ty2��0�P�˲��2�	X��ձ��.j9����Q����������ɲr�����f�U��/n���Қ:���F��D����q;�6�]Mvk�b��G�Ӂ�y���eظ!}�2�R�٥����՝|��5���nȁÍ�u<�RY:P$`G����kb�gD7��d%�%�����ibY;:��<���t2�Y�ʋ�( �@�Z�`�mR�jeN�%S>�:��ݣ�t��b��0UN��j�!O�*ĵ	��[��Y��L#���s ��<��lkj[��iJ�y�JsK��+B���{EȘ��231�e>�ٕ�f��9�E�1�`v��F]h43&�l��q�S��{7&J��b��̫ǭ<��@�fϻ-��r�����-U7��}�h�_DL�;����h����]Ei��݃{�֒����S�Wy���2����m���/��n�Wl�g�3E��[�d��@e���4�{OgL��m+Ţ�8���C�g^Sˆ�I�!���_3ݤQ�.�	��sq�m��B>t�̳qn�O9Aо*l hv]貉���0�/aٝ���*�9��0 ]��o^�I��"�`K^ql�&�����J'��K��K��(�--��_7��KWP7�U0Mp�
�9%{����0����N!ݺt�Q��J�9t{���ZF���L���=�;�WJ���G^��F��Y�ʓ2���P>wF��Y|*�@��O%G0����0�ի��6���\w�6I��r��Y*L[�!!C���g-���>\�,BH��Z5r·-Tl2 s�=/q���ץ[���Zp�!tN�2
�]AQ��4���K53���nEBӺ�~�D��ژ�i�� [�do1-���wo�gP�!:]�qZ{�\Tƀ��:����u�u[8aZ�V�t���[�s/�"[��r[���i� �Mf�[�͝E!�f��c���ժ�H*ds�Y���Փ/�����p#�����m�2h#T.��:%���a�m���Q��@�
�� +��+�QX���MF(**�+�ɬQ)*1��QF�ZH�5����h�#E���Tl$m��6(�TIE�fh،cEIDlX�Q�h1cd�شY5�d���4b��Dhѵ��6���1��Q��H��66(6łɨJɠ��lF6(�IZ4��FD+l��Dh6(��"Z5��6*4Rm�#h)5��Dlj��i1ccX�46��-���E�X�+뻿����=O48��>Ƣ�Y���e胞�E����9ǲ7���K�Bmv
�E�tvtM���9�y�)s��/燀 �j����iQ�*��L�)ڠ���>�Ԏ�gY߬crK���U�82�L��s�~�щp}\P����m�vHE�G|��-�1K���"��fA�������jQԶ�U"��}j����c }e�u�:��ʮ��(ׂ<IZ�V�u*9%P���Q�����W�R�ыÔD�x�R��x�Oy�,��1�B�x��m���ˆ&��/mj��an�u��@�Ȩ���q���\q[V*�ˎ��;/ +^�Y�֎5~��^������"��f�L�"c`�:H
�u|(GDh������Uw��O*UU� Ez�r�U�M#�AY���?I℮H�|���";�LGʼ.}�xw����^ZOc�z���\�z�tz�ڣ�Z<�u�@��{G�Թs���G%PJ��-�O�py�j� ȨZ��0Up�w{$M�P���q~g���T�a��
0."@N��D�U�Y��-��c����\�myoV��D8ɡya����55%."W���0��"£��;K�{�<*gJ�k�^�3b�oK���t��<w�0�`[�ӗbMV�N�F�D<��e��5u�k#�wY:l�!dv=�.dɳ��/��Rt��K�XЉ�VTᘄ�-mb̻� SV"�n�V��c ���lЪ������z�unx���.1��`�[���+�G|9Hء{7_&K�ۿh6�u�9�,��y�bkn�=v��ZW(ׅh�����UԸ�;�2�u��"�EY]���d۞{ꇹ:N���%-��|j��պ5��Z���?XZ|M���i^['e�=Qg�\�߻w�Q����m�M�R��<(	,���{O��l*�ԧֲ}}�6x����N⾃'�y���+<)׷M���7�g�N�?P���d֫��
�d��_X���e��Q	`�P�X��1^[<���~����˥�>���&�OS� ��wP���%�p��,��I�iAF��]��Ξ��<�A2t������7�@t{;Ofe�� ��р���^������PӣB}��{I��o_�j��u����=r�����5��=6��>�t4LA<i�l���uRg�^�S�����{�.�y��v.*��m�4��q�.�҃G���k�( k���'}��z^=����0�R��(���i�џa���scM�MT(�ֶ9;^-����'�1�tg����
q�,�;�� Lj���4���u�ۆlI��kN:�Bq�|��/�t�)(��'A��Z�D�f�7p^ZG;y&���0��E`�n�B��לW�����Q7hs�m��P>�ttd�����q���o�݃���>���z B����C�X��MK�ΈvgqSMv�.��y|h5}� `���_|�W&����U�`�ȵ;��@��GDnR�٦�z���tf���⼹E�!�ͺ�,9q��D\E���7rKv8�n�2tyMK��#�]_*=�ß5�;F��q��߯ɪɢV��I�~�&Ny=,5�R^���pݴje L�B�
�y�5�~j�'�������\:�k"��͛�\�Xŕd1�|�׽k�N��f�YVf�U��|X�k�+ݝ�
�[^�7`�5�[���'�����2��(J^��.uE��㔲��sL@43�ʰ��s��m�q:k�ܚ[Fz�-@�b
*X��"�]���o�>r3�MGq�>��e�L]��f�ޑy�1�OIK���n��Bc�{�d\�H�)�ݳiuh�^�H��[�z�P�s��8+- ��3�h��v)�#}rF4����Jy�O��Uzг=����J!��]�^V;Eq��l`͗yue��Q�8{�&��W���5�1i�qV(��� u�7RC�%\n��79P}��)j�">����=˵/K��j嚢ےA��M���/z�ի��i�5t^��mö�V����ꪬ�<��~Ѹ�S{�X?U�pJ���@h��	`�2�E�֪$��ݱ��!C�n�c�b��rz8D��Ӕ��n��T_�:(�t�q�Ep
���עd�ϔO�޺�ӛW2�o�^Oͬ����k�*��|�9˪�F"�h_q�N��wU\����<`�ťfd����ٳ�C��;�v���:<0_��a
&2<3AR�E�����bΠ�Gl�?���{����*�-��7O�ew�&_�oɎv۞�C���s=5�F��D"=#�����+K̓q����9:H���y7n]��u[��ݙ��;0�����:V�j��s= ��qy�S6#z�K����#�Y�H�y7��]�R�**۩~� ���_/���[�����ʼc�l�{�V�V����4h���ŰW�($��-�1��Al�1��>ڃ�+k:m,(�*�<f힌y�����uZ��ML2������4_n���&1+��c>>��g(xuz��/T*�0�r��W|���}FIy��=$�=��ߗ�J�u�E1����Z>�.��w�q�԰[�Tռ$ݮ�"G�p��Q]EM�O�FEH���o�FE�m���Fr�m���o�P��dG3q������U}��s�Y;��m,_N�z������[�5/l-a��s�U�ǭ�@�ی�e8���}{=�&#_P��m�wõ:��w�.|�gz�C�x�F���޷�7_Bc�
��W�s�5����.\N�4��z��s(f�0��;�J^�{�=�oȐ�z�߇���J�:���J�[K@۝.�fn'�d<����CT�_�v��y����\�q�|k��nǴ�&��P�5�r�"��]q��x-��4�
��d=7��x#�͔�N�������Ib�bM��r�Z�b5����a�y4��qP�4eRW��Wef��3w���c���J}`u�t-�)<��5�1��o��*��Z�uf+��W��Lo{5��������]j�M�u�o����Yq4+�3�'bzS��o0U�zr�S��ހ�B[	��7�rL��F��<���y�خ�#QUvɣ��3+P�T\т�;6$�>w[���ֵl��݆�˱�"�LK+r8\N䩩�����f�r+-�R�d�[��G�]f�)v�\�^['-A��hK����թ�up�qǀ-�� �%N��n�^��K�C܊	������6�>���mT>o �u���t;�FwtfZ�p���֊С_�
�(��נ�j�ӱ�Y��I��)6�W*�2�/2kw� �C��Q���p��~ؐ���it.;2�.젃�@��k���T�y�)�����o�Tj�דc]7�*6�ȕ��M��g�c+�vd��q�[ѕ�%fd�{��hz��X��V����G�m�ۺ�6޹麝m�W�Y�\t�-�Fb6������'��0*��藾�"����k{F.a����ٺ��̄�ј�nr�y�H�ҺN�Z��^��cѯc��^�t�~���#�3Uݩ��m"B�d�k�N�ND�b��Z0�ZZ��N������(������_nߓޡ�gj�wN�m��� 1.�u���O)�ꌮ��2W_�p���Is��}�<�Nj'���mY�v\���
R����6��WkZ[��OMq]��Qf�����`������%�^�&���_E�1f׫��v�tԯ~��:�t�^� ;��Ǻbˉ]�h�0�6\�*yd��R�J�ۤh��{݂��� z0N�];4��7�dFI}":_V�R�J�kyoa���>��ogx���v�+�w^���U�]�؍�P C�RR�;1���5�i�q���O<�mb2�rYȬ���{Ag-�m�\,����u�K�wG�{�׶f���b�O�9P��aά�%�v�gU�R�u�(t�ٳ�Gv�\35z5]*+�{��_O�uPZ���qZ�=�`[b����;~�h�T�H���u�;f��]��^�Мo,qJ�ލ�ɥl��~��(&�W�Ӓn�xL�Tvݖ�x�VЎ�<V��+rkw��6�s-���65��f�wۖ�;i��c����$:Gk�SP��D��C�mw<v���2���q�V��Q,&���7Z�ĎQ����OfT��Y�m��8޵�;r��n32�t�ZÚ;I�P�f���U��V�ny y�z���w������zڹ]4ZFv�t���8NɝTݫ5�w<�7��>�i�^9K�*׌x��BVu�[ �s��ݾ��Q����Xi�u`�(2qh�<9��9x�L�	��Rw�J�^Z�\ȩ`��m�튳�/���#pq8��t�}���`�8�yw1_xb�W�nڗ������-ߡ ꖖ�'>���E_��V"m��v3�{b�Y��>�����+>����w�gV]�X�r��b�v��\aK.�7�M�P�N8b�ax����]a�ܻff���
��یVZF���,=T㲋����i����%���I��y�^�j�S��,T3���F��"�_l�V���!�^5c/&��B��~j�m>�:Ol��[g�<�4=���j�7�k_��a��|�Ω����O>}e��=���Sm߄T)b:A@�U]� ��%+�����bP�z���T�k�S�k]�g���h��?z<2��� ��#�w��Ƴی�1��'�q˖����f�n'�m�k��6[���7�����3
F�t���]h⺖�m{�J���ۂ�WW�w�z�>u�Ҥ2����>n�K���Vg���M��8�w������"�m�7�l�
��l�"hun&%�2Y��Yp�7˩���������F����7Bek� R�o9���-�����[k����������v�H�&tGt��\�U��<2�˙i1��g!vX�M)��)0�lX>���a4�m�0���=�[�.xwqS�2�i�v<p�P��-|q����b=�M{m(���~��y[5�V�$;1�P��)s��c]�#c������W����-���vFw�x������{]�n�u6�e�#������X���k����Ւ/v9�]BVeO-}��h^ն��Xr�\�y/T�/<=�.m�%η]�&�N2}�3����YC�:��w��rx�#�xjfh|����I�}�����o吝-��!��Ҋ�#���}J���崯)�v�JW�ŋ��Y־Mn�oP˳��3!U�ޠ%�P�A���w���ִ̙�э��)���]�a=T3��S����θ}�|�/����h��J�u���J�#���oOS�{`����2' �*߯�	Ǽ��b��8��vg�x�X�mIi�mm��yn��*��|�o kdy�іW'�T�:y��"�D�^7���IuX<,���K�[�9�����G���Y��9�'�\�ek��䛠��4��H	�zh�<~����덥��UҸs�RV��\]-T�F����o94��7�6uP��p���%�<���dI�W�E�T��RymC[~��hH����<:|n�v�e��U��N��T9�����F�=�j^��o��H�٤ީ�V�^�u0�PΝ����R�S�ޟx�;?_��1}F��t�-V�m{����Er�+��<+���T�q;�0	���s�%�~H)L�\�P]�;)f�o6�/��j7�ؕ(��Ѓ�x�J�<l��ܫⰳ��S��[g㉾t(�9k4N�lk�lJ�8v`�z�͸�����r��c�~�r�F��O��{�;	�6�<�����NŽ�N�y�U[�6�+1,i]�!ڡ/3%k��o=<j�{^�fŪ��Ol�^�����jrݧ���V^Y3s�Bs��O��|�oɇSM�[<�����=�u9q��������!Z�0�bLf�[��@s�������JntZsj�r�a�L
����K����9����(�uq�����_fC���t.#�Gbs�+ũ�t�Ձs�G6���'NB�C�ހ�;�-ڔ���	�uhkYՆ�3-�T��O,���TPݓ{W|��&GoG&D����U�f`�W����s����ׄ���luV��o��U����Ц��Ȧ����ƢV��XjýD�8�(\�:�1gs;��L�N���g����O6jz���w�Jܐ\�4��"Z�U�$��*g^�؄��2ظ����{L�ZPr�˝�i����53�S)����#�H�����7^\{����2e�G[���1�c���r��Z�����C�f�KD�c0��\��'K�>��g��]^�i�f����u%q�MԷ��v������(��#M�z�)�`H,���V�����!M\���x�	T���Բ�[@:���#����D� ��Xn%[6i�;�oF�=m�"��n�XT���U�gpH�Z������""�+��L̂ս�]ӭ�����gGk&Z��]���]p�6�S�9ɹ2U�BI�`NvU "U�ҋ|�nա>7}�n��ͩYxx�ou㏜�1�j�ئ�x��8�KH��w���$��w�(N�쵡���f�Nx�˾���]W�oV�QUb�賧L���R�!T(�4m��q
C�Cz�J�A)�[�&�<� B��BHa��mVs�E�iU�M���dGA��ׁ�n�^m���` ����]'.����"�8�����H�u�O���"Hũ�z�[�+>���H�0�N�r�Y�NԉS�v��ѓ_#J#]���H��7+�HI�����.Y@�t��{�돓K���&i�B�i�u9���|��_������ٚ'-WJ>�՗ů�.�#���|�iT6�н�GѴ������p�%�!�K��8l-�x鎂:�t�+N�w���*�ӄ�'e��p�x����Z�Jw�M�;�j�#"�d}9qW˫ �p��\ѫ%}W{�➭���f'5��o�׆`ٕ��!�6����m]s�(4���4t��۷G�(��A��w[X:Hʏ��`���\��6�wGڅ^��G\�Z˩���t;���sC������n��&�q۩l�{�l��;闃�]����W�,^��.yWQN$����Ř����F��2T���-(Wd(X%��ɉ�u�D���ty^Y�H���yY��c�82�SJq��;4!\e�]ˁQ���� ��ʑ �
@6�#�Q���\�|O'k�s*-�gI���̡���1�B�.�v]SHz��<ŕ�P���M�������&qj0Vw`Zz��f6�#4|�si�X�A�Ǣo/A$��F���- ZTh�!a���l�-ƈ�Q���6�PV2�-6M���4`Ѕ�I���DlQa6(��5���6��1�����k��5`�5�V"��ll[���[c|q�cE�pk�ɵ�5j6�Xێ(�Ÿf,Tm�E�\hՍ�ѓF�Wq�X�I�����c8�Qh��c`�渣m#�o���}�ק��tLҜ�=Ҙ��Q��Q���G6e�y��Cp�6c5g{@s�ʖ��[w8,s�iX>Ntq^W`�[X��,Q�����ɍkQ׷�U�x0���Wo:�u/����q��{�����WO��wN��>�JD�׺G8�T��nϝ�A��Ǒ	�z��n��7�O���O:��_��ٚw/
1ۼ��
���.v��j�Z���K����:억DI
��j���KUlF�)�$�����k��5�yݬ��^��u"�^qvN'�g3��;o�;������>6�<x�=�Ϋy�ƕz��1��Bul<��^7b.І�tL4�4EX��&f�Ķ�GKg�k�)况���gU�m�Z"�O��2��m�+[��6�5J{}�I~�}�~����u���m���b����h�t0�@����Vz�����k�����u-��M$��(���p�e��~x�#��I���e�E̯5���U���1_���ՅaO8q}@k%����k���fh�lյ�e�dY9'�̷��y&*nD�fg(�醷q�m����ˋ�'g>�/��xB��y�/$�xWT$��2��1��#�6n/�f���b�̋q�ۛ��g]�k֬P��o��m7=�٣+�Q�IhWRf#�����V�)�L#bv�OS;P\��v9)��,C����2�F��S2��>	G�/�q4cZ��vc�h��!�m���u>ީ��z��ݎlN���v:��w�,a�ha<�]�q�"������Nd�F�wf��-�{K�>��cU餾]+.;'U�F:޷��*�X�1I1Tö�r�x˖��N��
��k�Ɲ������Ӝ�B|����/d{c�q���V��6�Crjlq��u��9�q��w]5u��SQ���$�4P͝`7���>��z s]/%k��>�}Z�����+#�T�Ԧ��[5N��>s����P�v���<�A�a�m �e�⺽�ʩ-�F���8��n;P솲�O�O(�mv�ꭈ��˓�s2�F�7�X��C�F�V���OOn9c�����)?L�:�i�\M�_J���3��[&Yӱ��r�EQ�����%�W����7XK'1,���.mܕ��1�·����m���+r��lY�:qV�0�;L�?*�\j�ra6�&e����+)�l]��Q���Xʭ�ԧB����x�'9{���W�2��o�}#��U����4�zޠ��NcV:�
��)�O��Z�h�%Iw�n�т}�]��ׄ�K��j��c��c[��}W˖���o��>�O;m�A���{S��K^�כ\.O����"����{7�K�͓���؋�A��W��W�<f\�0�t���Kc2/#Lw���-��wl��[��>�W��u��C�.fĪR:�ڃ�mX+\�GoN5�rt�&�.WX����-�_Gw ��.���xd�ŋ�: o��N���ݝ�=A��gyf�R�o��$�hZa��lm53��LgFAi�e�b�5ir�޹�mv?8�=���.oo�XsO)Ξ���f}������]�~�a��T&���R�Z�Ś�������g��zb���潩��ťdƺ�����$b�v��ON?B������
�q�S#�2�\����y��@�7���y���|�/yb�R��s=\�=�q� �D�׷p��z�����\.�m�as�N@nh����42��F����S�m�wE����BT3��5�c���$%�~�����^�%t3E��r�)o�]�L�q�־o3_f�˳�5FeA�X�+6K�6��Ã,2�I۷���9����$wjP�-+s���휗��2}F��O��U���x��+i﫸��j��Z�Zi�<�]g��p��%�o[�":���6�KT���a��okɧ��X$�O'�o����g�T
;���i�6讔sRx�5��fa��E[�w�i^Nnõv*�k+ܭ���!{z|P G#w(=�v���ב�v�F�*���=��mZ{���x�W�Ҡ�{{dzب{T!���m\�8"�щ.�T��wX)�ⵧ��[��f�0���bt��u��<�%�7�s�X��,q��Cy5~e�;�<P�R��Gs��WF�s���G�[������LO��:��E�s6Li�DeHv�������Ek�lɑ����.�\F�{���b�V�MЉ�~f���|v .�:��}*�,�1:�S��Cz/��sY��T&6�5�!1��+"��{U��NU��Ѹ�w9~~�5+rh{w�.Q�Yԓ��l#^�ݵ��F�%t��/]��b�-�C�+r9���[]���ׅ�̬���N�ǒ�~�z�r���{�����U�[U|{k<����T�.y��K6-�1�<!�I�:T��sA�;A<�tkxj�O�/彃�,��9�����T�6���}�z��5&#�)�u8�3^Tk]��v:
C9��qiYŅU��b%te��	��)�),[iVm�[�n[�K�?0�ѣ�w2���:����}q�v.�����y���3S��'����"9�݌�f�=����恿:^X���F�X[�	s{��i�l\FTN�ve�]��Kk%�j��Э��<��
�^�W��PƮr^擳����^G��s9��'�WԮ�� �a�I��Yl^OT#s�/���2�yM�S���8��8�C���dX�`h{bʾ�}��<���*E�mK��cZ�p��}@��̴b�[IZҪ�Id�viT���&Z���<ές�V���KB�&�b�v	�ew\��l�p��c��s��N�v�J��̾�F���R��۝������ի��l<��-������Y����/��K��3����;��6�"�t)O,%�vk�-���!0�����z���v�Obxd���_C{V�����yk���op'�-��]A�z:3	�J2��Ewxg}�P4�h��q\��7�J�:݈x�x4�5��o��nu�u�z��D�/*�<�Е�^��Kz6�K��Vw7e��FT}�&�:�c|=����\�/���@�6���Jy5ڶ.�5@�֫���Ǫ/)��Q�I��M�v7:����l�g�ߍ��T��$�BjA{��2��g)�Z�uZ�N�,a�y6�O*���늯y��w�]���O=K�o��)�mmc\�}�/O��<�?W����v� ��<皬���M����B`Cً�Bm酑}��h�q���5[��Х��%&�KNXi�G��u�|�˒WWs���Nu������M
ײ�����RW�;�e�A����o�)ӭ���]+��n�Z,��^N7,���nWQ�En[�y<�0�-���:|��BU�}HMA��1;�o!�Gq���wm����]�3�ꮻ7^N3(��O�Mעy��g	�|9�v�7.�Џݎ�Ƚ� ~�#�q3�}S��ո�ٟ,��6��uH�*�����Z����k!d�\?>��Γ�
�v�O�;^������OT�x�t㪜���J"��ǵfz�+�G��Og�^�k]���:�iRlL��u�k�.��9��N]��R���5k!c	���6��1˲������;y��#��>->��E�
��)޴��0����^	�v�[܅m^�/gH�#������Ե��o��>�K%w97�7Ӽ�x�̼mleyU9��)��}�#���⺼���$D��f�6J;���^�ͦ�C܄��sNh"9j��}���.R��/���:��o!�oؔm%Λ}�<p�P�Jz�ڃ��fZ*{kF�#�l_����j�D�G6C6��U�1ȑ/%K9Z�1Z�,���^c�;�+0�%����a`�n�N�"bws.�<]�YnjEOI�(� ��|sTt�d+�h/\y�3K��L�-k�!WOA�F`���X�6�]�V�#4���Z�)�',���]�}'@I8���#a:1c�l�H�[]�w�-�\�k*���s�&�2|7U���xZa�	����v�>:�����oG�
#��hOeb®�	կ��ym^��\ޭa�g'�I�U��z�uͼEe\�6��r�u�q�g�j��>S9�+���z��vճ�8�;��+��4�φ��]F�f�v��~��0=�6}�:ǪE�������qΨ�ػ���n3ε���ݿ>ٴ�gZ[�9W�������Q��IX�V��'B��_>�=�B���v����k}rMy�=&M^��O=C���|�u��U��V#e���-����η�>=7]��5��z^n �{�ͨ����:��e�-T�F����i�;kG���	GoЫq!�[�֔��������~x�呷G���k;��T"f��C�q{iYZ�IJ��ۮq^��كOR	��x�3&�]���rn���<�/�e�v-��΄Jt�m��>�㥽�b�U������;�����!u�*�1���N�P.�VySn���x�N�ff�U�r]�orm�NKN��*n++PX�r�m�P�{z���wmy�'k��;q�f{%���vK��K�X�x��J�
{��K`s�sI�;��8��.���ƝT��m$�{�>ثn2��4�)�yv�'�VC�N].�h�������sj�7�8�Kz7�I_C�x��M�L�o]!�B�]~�������;<��^��K�mr�[}z�;�n��]�k
]���v�w���w���sY�<�k�m{���[Y��1%�W!��UpV�*%�Cz��7��`��E���	�Ë]^,Nތ�B�0���fe��V�a����yT5ٽq����%۞Hb�A*>�Y�QQ��㗾];Nջ�R��&5��}G�ܪ�[�3(�ڭ'i�E+�����|��m����~��^�=��g��}�:|� �%w���F5�V��fv�m���_�7D�fMNJAklwp�o(�\�a��Pֳ���|��9\1�ٲM�;��!5t�(̓	ي�8+�qN�Qx���M�P����¥۩S@��>ı���l��g),�*���wC�ȱC���#��2���v��}�/]M�W�S����.�<���X��]�G7�<U�!}ۢ�e���������&��.��g��H45��qIsz���:9ʜ�W
�~]'�����E{�lF�1�I}Ci��])Tu����S�WE9=��Bym��'��U�.ª�#d�D>T$�p�}ۜb��bT��q�o�]S��p}e�a�y.X:��:{ �ё�g���Sn^�Q�o�bP�#o]�����l�������kG���}�ۈd慕�UF�߻}9<�ݬ�"3\P����WW���-�(�����[q��)^���Η��T����o��_	��P;ޞ��ѕ˺Ѽ^ݴ3�v��2�fjVz<W�����:v{jyl�Og�q�Wf��	M�kp����xfY`4�;����lO�(�u#��G\��hK���N��;s`RY��o�%��w�KP�<�woz9�3, *�Z7�����em��m�G|<�t�g�)g��M���nO#~��$�)�AOP�}�S*�*�1��6�WF��krG&<SH9�>��I�۫f(�t�|T�6�D�3���t�q�E�ʲ(�p�
]����� M:\H[\[�C�t�=��α� AƟV�X�1]M�;+0ueH�Õb�.&���X<4|�@�:��کt��-ʔ���7`7���jZ�3.T�۷;O2.Q�Q�cn�
�:����E66���x���ǚ����k�]z������$�zjIe�o,���>oy��nO_+5
�.��Y6�	���I���Hh�X9���YDr�u�G''7]f�(�R�g9�&*Q�\�o\xꖧb�%Н;/+kR}#�}�U�����k2�5
u�������=$�زh�G+

�����S�Ưx<���<����V�v�i,��sӐLSTqm9>��v��4�,��돻�
�$�'�u֛wV6��<�X�
 �/���"%1�#�*)�d��^)��Z���;�7�S7�xsef})yoqι�)ხ�F%pQv;�SRd8MC(H�4�M���X�P���9K+RՓMrxf�ٙ׉�EVճX�X�R��n����I�dN桜��2�T�ڢ���+8vJ���&U�4`YI6�+�V�����Oj�;%Jj&;ώử�Ls=Hh�\�j��}B��,ٗ�D�4�]����v�0���M@:q�\Hei] $��������M�r6%�{bb��2�V�R�.���6����
�h���ѥH	0���
�u��c�ŵ��+�U�_)	s�KZs�Ce��b��:x��M�dM������B�����ttu�#tR�!���v]t�#?1*�Lκ+$l"�;�Z�0 �G;�}%8�Y�rG��A&��"vR���RQ�Vͥuɸ���.�Mt�kfG�I<�Sk8�x�P�OC3��ڼ{ ��h���MWtvv�Ge�b����W{��[�N��¢ʽd��d�U��r�gS�kl�v/:����L@���7J�opn=&Eݧz����m�P��kOS����K�ʎ�쩎��/�ź����z�q�̙�=��r���$��Y�YN�E�_%�gJ[�&�W��Q�1ey:����K�y ]�E��c�nm
���.�=��[u;{���!9k��[X���d�7��և���y�Q��h�8�}!/�3�$B�޼ynm�Ӣ�vᶕ:�jW&2Twڠ٫9����{���OE\���9�D}��V�r$'3�c�$� �Ek��m�t��+�����ցP��qn;ݹ-��[Bq��V��W!�ɬ��/-[H����v@r׻���k#�*�j�5�3 �cC�$��YWp[iԣ4��뾹�:���w���5�h�E�b1�6�%��\\E�(�L��k��j
6�6��ƭ�$h�1�,T�lh�X�ێ-b�h̬V�܄b�V+cDci*-A�ƭ��k����q\j�m��U�6�\js�ps���l��b�E�椴Wq��,m�EpF�qlj8ƣj�*+��ێ6(�ŭ�m�*KU�Qq�9ʪ���$�M�;9]z���w�*�1�`�6����6���'s�e,¡�x@����<�x��V]b��r�_��6sx勫��;�7<��*�-�]ܠ�lk��:��(܋[B�(�ٗ"k'�_u������u-�ם��j�:+s��#h5���g��r�7F��:�"]nľ��y���+2�R���緳M"�9��r�ef5��׺��F��yd�ߖ�E�	��b����M��9��9/\rz�g��r�1�!欈�kK������$�֖�9~]���O\6������tD,n_d;��,`�U��c�5�~�sV������V��*�:�.�ӄ�j7�,�UNq�����+�sp�=�[�|�����Cw ��@9«�H�h���X�����l����!,m=s��7�v;���y��Ⰼ�p��;ꊳ^�)v�W�����ya�=M<����.�3բE�j�j�Q����-Dwnm�U��5��˂�w�, �S�r��~U�V�~�u��w�q5��X�7{uf=m�xA���{�0�U�/g��N9W�)ܵ<��!���w�CvK{��D�\�����ht�x�*f_,�M8�N�u��6Yu,vZ��7��M��J'p(gnB�.I�	�m�<e�(��uk��WoS����N�؊�+��W�p���)}0��Kg*��d��q�R���Xέ��ί_!�U]5GO��l�.�9m���=��Ǌ�]7��U�0Zj���A�ƎHz�UJx�l��	ճ�_����ERs�/Z�N'�-�{ѩsH_C�'
����A�=�J����{|�rΨ̹s�&�;S�.P����I��|������w�݁���m�a�Ž	�/hG\�{s.y�м[]�jg�i�i65���cOi��]U[�/ܨ���Vc�Fmg%���*�9�za���W���S+9��o����)���Ѭㅾ��U6���jmf`���BS�z1���
��&5�}Gi��NѺ�8̠_�1g��%d��3�ų7L&�����x������u�������vVδ����^	����$���u^��aP�Hfa�:3j��zr�J\P�9�՜�߃C��&��:�C��J&�gdtHx��uHLE���S�k�w4���ͅv���q��鮏<ssI�6^$\F��v�W�ڹ�����e��o&��ר����5����7qڍ��S���"P\1�尼{R�T�ٚެ�:�u�ɰ�V��le5�q�8[k������I�����j�yX�n)o7���ι�W.V�<����5�Gwe�,=U�>)��r_PH�J��=��Y-�s5Qկ�.�bf;w�O+���aM�<�#a
�ʤ��î��*U)FU*�M���hJ��0�cn�P��)�bsm�T)^ޒ���Gs�Rv��s�^Q�zR�W8�oL�ޙ~k��u<g*]%qP�w����T�k�Xoj���V�UÎ�w�u���i[7�S܎��*]3^Fׯ������Q��o!�|��=����;����W�_C�x��o���8��M��&��n�-�r��Q�AZ䭹��k�f�\�6�^NF�k;�u��2�چ���}T-8v'eD� �Q�rpL�ͨ�����.h�*���MܐX�����
�w��4p�Xb��,��ݝ�X�.Z�Z���r��J��Y��ˬ�5��2��9�up�+�uMͳ)N��޵2kK�TH]��ʺ��4/q�.I��Xa^<΋���ĩ��J�HM��v�ӷ�U���h�#r����Wgr1�v���M6ư�c���eU�{~>���>ӰH[��)�X�:�c����9����k�w��z*���_)�׍Y�2v�|)Υ~�n�{V�����>���*�ٺ����F�j��n��.�2孴�d���~��c�f�O��U��ڛ�4���IYD+�������1�=U��v�:s��u���غ(|�9�����O��p���c6���@gY��_��{�X�aP��n3��2w�R�����wv���l5�����
؍�y�Ff�C�uʴT�rO]ž�s�Z����	��S�*��aT+b6����
z6��]ӱ6^�[���S,NT*J��&����{M��V6*Ȏ��5�Kkj�Rכ�kPq�#1�����lҔ��ֵ���o�)�on�fى9���Ī�yX����o��R>u������Y�I��ǘ �gk`^N�%������Q��]j�V����a��f�]o��1���]�K���lm��\���2}�s�C"cz�n��HHmZ�%���b;k-�@��$�b��3v#1�������2��y�OM�t���=�:��w���w�ݚ��b»敾�X�c�Zi���!-����q]Kz6���|XV��91]�/4F�aH��r+��Niʈ\V��`��jV�_��M"M�W�����!��l���b8v��E�#����c�<O^���H��P��,Ò�.p��)s��lkQC5َQ�"���I�c2���)��*�Y��8�Wյ��j�u5i�i�#Z��vaM�fN������ު��m.EM��y�^ջJ^����9L?]��k�1R��R�ǒ+}P�{����o֗ma����;S��N�T��7U��$U��'Z��B�t�^4����ٽqw��	�ͼ��j�S�,��U�K���W���N0:��]��z���s��\��,��;�T�<��Y/;A�[Au�7�^cܷ�''��Å]3M�����dPZ�r<lqy��@���_���.�S�K�f�G����A���,.i
J�2���7�x ��6tmP���M��4j��BgA'.�7/*ᐗ�;�ϛ�-�DVs}��������|��Q�.؎C�18��7'֫�S���v��u~����2ٮk{㩴��ӓy[L$4��-(��	e���<�U�.�cmWK����y�DS��d�8�I}[T�*R�7l=���<��{��{���^[�.��=��-�� �}G���RR�t]Kf�����j�e���{�g]�Ce,�5ˢ߹Sw
W��
�Gv��v�R�?\��̪Z =Q����֜Oo��e�M�^IjT'��
�=�B�ر��4`��1��؜IBbV>����)�a�ְC܊�n2��sH�]^�4��&�6ۓ���.^<�)P[Ѵ�̾�`C�
�fĪC*��(�՚��ȝ�x���[��Ԯɡڝ.P�'�i$����c��P�\���*y��V9�;F�Ϭs��̹�^�[]���j�ާ(���/Hd�u���1���Y�R(Wu�v}�26��ub��G��*΀�T-�Ɋ�\�!�m��*j:�9����9�Fl$B֗w1��]�
�2�\�_:���ޘpc�qȾ٘��Q�p{%q}�!Ί�����.sZ�=Ě����ko�Wx����~�fS�.u�Vc�F"�s�T�2�cn}����"�u��,Ʃ��
[�s���Ow��V}6��>[��v�`��!>�M!1;���åx��+K��&5���y��A�7\�2�/�ř���l+����H+�KT��J���j+;
g��^��~�kf�ߑ!l�H� a���v׻�z�>���צ�(D�}b1	�tW�jQ~T�\��O:�y��#s
�y�9fѵZ3��%N�WGta]��n�x���o{/lD�Lw_V�%R��{l�E`'T��RV���ή������Ť�x�����R�/}��C�綦�	��lF�(C�RR}RV�nn�kb�:�t�B���:K��s�a�QD�C[x�ڷ�mͶ&�w���*���ya��h�\�*����絪�>��ƭ�CX�x���Ba`�oa�"7�S��4�u���/X{J�d]{[�eA���4]�R����:P�e�-a��=�*'Y(��V[r�K1��J�8�N�m.e�ZƬ~�i�"�Ψ!�j?Y�TR�7�iy�wbR���0���r+ú6��C0ل�	�jG�v��r���>��h����������	��zی.Y�2�#ne��`����kcX~[1�A�BV���*�ލ�ɥ`2��(R�:�3�Qȗ�mm�ڮ��[8�Z��T���T�ŕ�h}��m7=ӭN~z��)�X��2����޿B� )Q#�l�)��+rhO<��j����fcd%��Ŏ/2�J�,N%61�i{]��r�����v�%^o��+w�%�s����3��ǋ|�[K�Մ�����5����V�5�4Rla���<�^w:c�x��7��}��m�{4�//���Ϩ�=�UF����9�F:N5�7C�˪�����{�����W��fyY�}>����)�&uT��px�>�O�����KG���ʒ�u�!#�(�|�m��"T� ����D����"}����sT!�o�-pA�,���W·b���7"�7צ|ܖM�b��eov�t���ޮ�s	=w����R�:9:�1��&�:s`ʉf��co&;I�a�8	u窷�&p�rb�k\x��B�]F2T��8����U�4�q�ȠU�i�^V��)��
���G\�)mJ}(���_��59{�{�{cf�˶�A�=uL�RV��PH��ў"���bp�Y�oW_�S�y�i���_P]�UlF�A1��2I(čW��h�m*Ջ��Nu	���9ͽ�>���0��m=������*k�P����;���#�Dn@i���t�lҔ��Z�f��T}-%�3Ӹ�\=�����w�ܒ}Y}��e�	lP�}w��������w� ��S�t��޿�G���F��;~��@w`�خ�Om}٣!nW�Y�e+j�k�8�Gv2���M�=�M��5���=�C����eއ�����ǸBv���m-H�{�������5�*Q#������Ϣ�0l��f��r�bV���h�p���$��>�6']���7]n\�Ɓǭ9�	i:����r[̹�[W���U���z��lFך��ɇ��t�����j���W#*�e��9]`<�;�Z'�=���m7KQV]m�q�v�.P�l��)�k��*��<�u��Or7&�y��u
�(�eӜ��ܷ�9X��'m��c���e/�%��Q��i���L$/ws^�{p4� ��Z���ȓ'"-��U�Y�Ե����ڷ`%/l-a�5E�>�W��!��p��k*�]��1�L_1���o�IY}��ו�R5�����0kuhTt�Z�.��y��\H;���}����ד���=";y͕J��8�x�n���XO7�]����դ-��KG�6�o�Rm�չ8�6uZ�So�:\bB1����>��=��U�]� ���$�~���ڭ�Ӧ��0���{@�J+ݐ�6��\�v�̤`�R�:�Jbu5�u�Y�_Hyפ�l˔�Oj��o,=�����B㑜|���m��|�#��D>U�)wT��T�h)O=E�9Rw=�Q]kIs7)�hZ��n��
W��
�$�%��K�<��W�'i�re�W�Wd����o��-��uJhaw���CKc=���9ZWOs�N��g|��������D�2޻p�ϔ�k�D���R7GoL_vն2*�n�G0wM��o�R�/$Q��S/;�,^v��:�:��o��78B77�Z�ݾ���)\u؈��W[�-�-Q	�U��쏕�!�p���	�F�5�|{�F;��cB)ׯ8�Q��씰�F���5`�t���]f��,=����M��tK;�OJ�=ܼ4�껹�*��9���Hѧϥd�]=�P��{o��!s�{q�6^L|�7i�;k2*���}��k�!��CMoMgwl�pZy�f�0��8A���쒹w�ʹV�ט��%��7��M�ܾFp��C�.f��tn�j�p�+�μ�X�wxb��η��ikI1X6�/�b�·f��סVt��faIK4Ԓzt3��]�sݚE�."��@I�/ �:�*�C�ufI+��Ww��i��"�썭P��}�^e�f���ξ5AQ۹M�3C:P�,5�Q�y�_�w�q~QaU~cn�P�IWDL��V��pp�/vt�gD��͹(��
)C�=�,4��j]byxK�9��Nѕp�3�8n9[1��|�.��M�mZ�u�G��Γ���f]$�X]CP�n�]�J�:i:-:\��^*�t,�-���ܽ8�&7�:�c#t�ب����u|�YNU�V�o�<\�:�Rqtc��wdZ����O,����I���X��˃]62f�p��ۜ:��2M֨�Txr�u���ݨ�T~�O_;�Ǥňw/����d��c�����1��5���A<鋮oZ�r*�vWt�]0+X���PE��1r)�%wӔq�1��uu��m�1s����ع�jů�����/mb���S	׻��2:�-N�l|��M���kmw1Gk8U��!�D$TDڊ��lL��.�t〆�f�g94��H���η�wI��mI9ް�p��4z�k�l��bUh�Z�z��)hu����3�h�x%�����W���L�B��;����/��Y��X���=��Z�8�6x�!j�-�g��j��R�j�o��(�� D/�}2��c&�$���\��*��Uj.���D�,�0l�;��:�m?_,����H�2l��C���0��v��pؔ���z8.��v�"1[�[E�s�mn&�c�������E"Tû�&�q*Z�9BE���j��vgբbrE�2�R��N+2����Y�͕B�vb���m���M���s:(�r灣t��"��W{1�6*G>�wU�W� �wK��M4:7���U��	ed�K�[�w��R����b�o)�����ԫ���ۤn�X����"�Tfw;���ł��oN�	��G!��V%o���w	�A2��&�y���z�]i���y�HC���5����w!+*��ܰ�0�2���n��0+�N,�K�+�+���u�� y�b��k!T	{�-���]���u�ۜ���w����������qc��j��n-0n5q��6B��q�q�k����-�h�,[��-��4F�.ƣ�4b��q9�\Aq�9�q�qƮ5�6��M����Wn5G�k\V�Wn6��J�\b�Kn+�5��qks�ۍ�q9�n."�\h4��79�"��K����I�1�˚�Er�4�Ú5�9��\\=r��|��Ӌ������}��g�zQȺ�ἱ6���s&+��A�ގUt�:*����y��o��}zf��{�����*Ë��uW��u��V�k!�E�-�y�'\G/��`�+�o�欦=3���K�wC/nh	�󡥛�\ղ���
�6'ʑg�M�X��kYʞ]�S�����AZ�vM��r��Iԓ��z��6����`R)�ï��sE���mC��[�~�y5x���x�R�U+��튒
y�t°�a|�޸S#]����{h��%���9ˤZ���xu�k�
���:�fe��m��9����7[�c���'���3Ҵ!�1�����mj�g.b��ʅ�s���&1�}Gk����n��3(��"3{2���1w�R��j�ٰw��b��y��Z�9���Qn�so�2ռ/�E�{�7<ũ~.��3���"X}q�_.��(�*J�Z�iAYc��4�w����&����.�A�B\�m ���W�-���r�Cб�E�BeZF�WV������nfuVu����U,!H��&�5�-��se��o�Aɴ#ٔxS�3�]_�v5.�~��Ú�)���U7fy.������R�l����Nёl4�\����N%mЯ-�x)�Y&kiWu��,��p�����K��\��
���v�[�y�T$����T�ZaLőM��e��˦P�^4�ä���+��>[�⁇ʄ���T�V�3K�����+M���47������=�o��m���+��P�k�*�g.WooEg'��t0"���ܾ�om��vc:�x�W��V"�l��-��/��k���@���O���寺�k�x���h������3��'PM��sų
F�p؎{:%k����f�i8Zع=�3��'
��J�bV������⡞�z6��5+rhn��6g-��;��.\�����Xi�v!���XE�xd�*�e��MN�J������/,JJ7a,��Ʊ�mQ��8�	(���VD��}��S�驼CB�f��Ur�wV����W���U��N�����]A>��~ �?\Nd����x�����B{cI��:��wT�:���k,��DQ����߻
мg����J�m�v�5��[�b��|�/ۮ��D(��QK=@�'�'�3�Qi��&kd+�����O:��M�22fޖ�$5�:X��-8�Y]�����Y.�Q^=���U��Y�mVO;ejt/j�E�bcZ�>���[����)��ǀ���L�w��ݺ|��:��F_�P�V>v�^E�-]0.�ƣ/4\O>��	��{�4k�]®�P���%8��b;��p������Z��N�ײ��[�>�&�����;��vW����s�(4���3�KZ��)�Qx3�:	s{��j�uۭZ��;B�#g�T�9��V�A�j.P�cږ��2�ւ��R�����	��'�⯨v����2�Y��R�yb�RfF���5nK�:���ͽ���X����
����4�E<ǵ�W�؎����iu��jV�)�kZ��s%mP��(��/���5Ҽ�Ɲs��R���-��}c�,{,��6��dd���1�<�¡�Y|�"�E�<XF���D Ov
�دGoUni9�o.mJ�6t�0e�hM�����	s���(e����+�㝁�\CDf<�o*��.z�F����N����0S����^f1t�evX	��G)�ui��`jN���j��)��C�����1������,���feJ9(��gu��[]Yk�\s	��V��=ȯ&�3.TB�Һ��K\o��O�s|2��W����=��	s4};p�P^T�@�����|��������ċ�����h	o'���8i���I����P�vB��&��ygO]���٣�7��D{�.q=��[K�Հ���L2���<���$�v������Y����=��Sj��l�~��=��>5ݞr��lvܷ�����^��6�m��uz-	�ڴ�j��nV�G�R��e��B�4Ű�b�լ�d_'�cTv�檣Z��|U�<T&�1�i�Ü�^(��A��+&�-�!7�;�S��X��]�{N��}��]T����ȓ3�"�u��s�"P]b1��j\�9OyWn�k�DA�8�,��6�1p��#�)פ��6�J�=QiGd%|�}a�<��[3�Z;5�t6ؔ��V���[S��^�*=����=���٫�1P�en��Эێ��T�*�<u� X2�J�8�k�q���8�Tu�5��ے��6�2��W<�/]��n����Im3d ��C�˗�F��xD%�c{\��9��lZ�87��gg"291���ڧ*ժW�Xa�\*��\�O,�-w�Gu�ꊧϻ/����C����Bި�ݻRV}��+X���X���:i�S�B���P�����2�tؘK��⁄�P��{ �9x#X�ف���{=��S�QO�1z�m�PuJiR;���3�G6��n�Nsbӵ��;�8�[ݼ��3��yp��~�L�FLځC�=��0��2v��{�NoMOb����f����u���w�x�_�أ�:f+���ꚽC\�u�(��9C�W�Z�+�hv�K�4�J\�v8Nj�$r�����R]�h_$n'��"b7��; ��;�+'�;G�ʿe��q�����g�(����37ݯ��uE�J�sm�K�4+]ԃQ���ô��'î)�a��Z_l+�[��~�]q��w��ޟB�@:6�����o�_�}q���Q��F
�����ݙ~��'NF�����ƅ1ڄ�d*]Ak��u��i,���6�����ْ���~F.3Ig�+�f��d���z�k"��Ὣ�}��<�����Ko�$ ���u-ܗ)��htGd�,��9t��"��T� })ȹ;�1�vfwϽ�U3��,�l�{o�F_�rq8�8}w��^ibћ<����`�� �1Yj�v.A��hJ�Z���஧�pY�L��m0*����*�~`��{НX����11��`z�.�	��#21,4��'0��ŋ�Ma�J�}ᔀ��W����V��+�G����۩�Dz֧��r����J���vQ=�f�;0�N��Ґ��rݐ��۹�~s��0��q�^�7�A�U��*�B�eH�:IӒy�3�
A|v��(�\��HT��=���Ӫbj\c�v�´�_�c�O���1�����H�$�}2�����C�eb�xz�Կ�����u3����V*�r���,�>d#�Ϯ��5�_���֯��*%_K�]��^րp2p�q�/��3�n�Uķ|0y�v��k���㸜��wh¬������!��Γ>��Ε k2H<�H�'�O�;�����ڴ=}���7]��z�*�!��NN���m�w��/�v�&ٓǀ�� N�ζ����x�%p��F�MR��r\��T��^mؾd#Q�V�[�(T}�okzQN�-7�\/2�k��W%�:�]����7�?��{;I��	Ɠ�fu��=�����i8�ʚэ�k�[X'.�Yv��C
̫�A���'S��v�="=�S#{�ךݹc/�{��{��6ݓЏ���:�-۸��2�z������D��tn�ӕn�s=!�j��O��U]��7]�=ࣜ6�I�m��0�^L�}�J'@%3裪�^ׁ�3�l����s�����x�NQx����G.���[&�&��t<ؽ?�G9W�'����Ȣ65Eg]��f���!I�	��B�m-7���;�1�)Ѹ�����w�oK�0���j�[�i/m���y�)��]q+����:�wٴ����~5/.;��VC�=�Bkܵ�\�dN�{��XG{�>6�'2��1΢�W^��J�������|���'�9�� GcL����X~�ٶ�4�KY��jw
��ϵ�+K
'�4Z�7��(\�]ϧ���;ӗȇ�Z��wQ��ͪ�ކ��\gO��O��ڎ��U�X�G�1;�g��b�����J�K'~Jy���p�^w��k<�ӣb�I;S<��-�1o1��Q�}|�y�ϲb��	Sk]X^��p�/
e3�!ڸ{q�{��4���i��%ߩ�ʐX�˭�{iG���,8䍇F�M���G�O*���DD9�k1vm]�i�����ޕ0w  ��vB�,�	���i�$��'j��vv]k*v9-� F.e�
am:�t�*V����m��6��sUZ-�����`80�T��u�G���X��N���Hg�v����ۯkN��[���I̐���c�0�I�P��z��'�{�\�����K�k�(Z��Y-��DG�O�����ww�s���i����n���f�7��0�L�I�'��xuB��Ell]�{۞�V����<s�hn}I�nta=n�ˊwhM�����t�rAJt@+K����"إSw�q��<��8^.1�Q���G�9�il���v!7xĺ�f�S$�Q�+���"�ޭ��)��C٭�g:��xpg�L�7��q	u�-�Ĳ�.q���x�{\s�17����u��E��q���]n=�s`���qN{\Gm-7�s���]Ʉ��'��_���{!zA�`�U^�/6�R�2O'���	~1R�/��T�߳i��~$�w�N��U�]U��Dyz�egVR����c] y��/{� �l�z�zam���t�0�\�/�����*[����=8�DݪI�����Ue�����N�b�}����q�c�Fb�m;��i{	�΅��p��n��+2 3�ZOkV-�qԒ&�XeY%%"�zv�պ�g �|�vØ��|�W�A��GӦ�U�ԅ+���`�kV ��t�=��N+Q�����bإ)����6��)R;�1bY6x�w�t��/�޴���&���{�{����.��1����֪��O	�*cZ����u�F�/O��K��2�j�	��3���F�.7�-Wvs�'��#Ǡ^��O�5̲]#��j��uf��~��q�N��錻t�^�hu��d'fÓ�p	�g�J�b�
S̰]O#��}q��y=���[M�̪�Y�����wo�,z��,_�2��ڠ��١�������Ct��{�Ś�
g��h[}���!XSza�ʔo�:I�3	�3ԅ��q���)z��B�����t5����`�,Pk�xq�tC��;A��B�WJ8��z���H?*��e+���#z�|;�����'�QNm�>���;�t�y���0�%TB���I@O�*`Ճ�5Y��7sz��s�����V5B��[��Ц|�i��a��vF\C��jÙ��yT��!m;�2~]�E��Igr���`c,_��[�ü��F=sm��;��n�亦dn�&Ψ�CWE�c:[�!lt��<�h])�s��XW�޲5.�_C��Y����`Mµ��5e���7_6�偢�+��p��9�1j��,�����f\ݫ��a�������׀��X~3/=hm���j�Q�W/�ɲ-��Z�E��-��Z���}԰:��>+]6�d8 �enP]����>����)��4�;�D������]��e�(G�R�5�e��&a;�1R���5��H;\��/���C��y1�6*���v���W�!�W��;����7��x
��rGJ'k�d-7�~��[Y��Q�r�=�H[o�1T^x�G��_��sUto�'@9�큥���dGK'j �pr|:�f�m�}�O|a����Q�:�����,,�N�O�k��(Vo��_�i`��>�:=�v��+�]s���x*�Ck�u��.6�i:}�)�muC�SOz98�ec븝�{N�>F|_������=����#���fw��>O�%�c�z|ճ�|_S'=�H
�}�cʫ��8�'V7zp����x3w߿~g^W�Y��?z�K����3�_'�p�A�@>��@Wb�\Oj����iX����;���kK�����}J5\���)Y��׌�t��m�(ِ��x=pj$����r׷l)��D8�ө��?R:�gD�_�vT���$�<�A��R��96�x`_��y��-�	�y�w���=���F;��}�Lo�z�/�UD)�Iڙ��}T���Oۿ�r�9�8���4��u�P�Ǉ�Zi_�P�:4���s�ǚ�Zy$D��s��
��|�Mr�*d.���6i:�҇q;CM����!�YK0L�,2�
���t�$dPЗ�Z:�j�[���y�C38���R��LM�ww��,GX�:�Wn�k�,b�����Bc�U:M��q�f��	ض^�B6�(k����'q�SJZ��C*� rձ���a��W�;v�n�� `�J�R;a��Y=Xd��&Ԥ�i�9�+�W��T��%�-�`=�1�Z�[�j"�����/2D&*��SFS�6�z:�Z�[�(My��p�)���n��J��\�κssq��p�ԝ�v,�Z��ƀ�����+���0��N�Q������[bN�ë��(�On�N
޽�r`�PW\�e+��5$�g	�U�E��ѫꅐ��6h	�x��z���H��X���7�1��
ܩ��;���)xu���l���j��m4�ֶ��F��y��;]�6O�8 dY{��]��S����u��|�Q�n�0�W�,d�u�YV�=Y �WnQ�b���'��Bq)�.����W�����W�j�J�u��m��M���hF�}k5�2x{BW���!��*��]�7]��_���AVW#PT��z�����B�Н�O�f͍��n6�gn�GSǇ#�}f���ܓPf�B��8�vd��tN������n^�W$��vCWN���W:��[/�L�W�J��U��9:�բ��(A�2\��|�����F��1�����7o�]FuG[ð�G�e�vH�V�]du�/e*?IHś�}W�b�����ָ��T�AT��ed}Hپ��Qm
7�Z��r�l�I�+6~.� w�4T���2��Y�}A�)�V��`���[4�C��C���;_ˢgc�b����Y��	%�A�� KM L��7z^���*L�9�T��Q;��N���xj�r��{��i�m)�et�+��1vJ�]N5�t+Du��#��o-�u:m�[N�w*��KlI7V�Ɯ�a�6�����������@;�M�B/��@w�`����;1���܃REaG������E�vUeq82�}��X3��LB�ޫ���2���t�~Ǥ}�#X��B>9����wղ��K�jRe�iY�*��C�m<�LF���$���+��X-S$VM��"����-M<����J�%h�eCu��)�h���Sz̤�6�N��q�(�MVU�9nV�8u�ebޫ(ц
f�����u�}��^a��m��x��m��ۢU���U"D,�
�q�*Q����v(���bvgN�B�[Kz�O+�*@�J���	�e� �/�r���C�/��A��s���z(l��n��j�9P��Ƅ�ڙL�jTX���X�vj5���wF �:W*J�nJ��阭κ��^�����u��Ϟ��_ac`}��s�D�	�9�k�\m�iLq�W.r�7�)4l2��(��X����lRQ�IA��i˘����cL�X�M#Q��pb,�l[r�䊄��c�9�\�4l%$��b�c�'9rT�2F@����� ��0��(��K�6��0S61rn@��DQ�H�nc3���B6���Dɤ�H��h�qĮNf�����'.BH�IA��L*H�M&�sqrh�AO����[Ae̾���Wn�:RDŽ��5��R�c�Ĝ��\�Ղ�l�� �Èc��x�/V�a4MwV�\���3�}#�{��������l��S,�+Ub�+z}����1�gn<��o��y��D�^�thR��Kc+3����	�l�5 �:-��g���
���|�;\u����Nm茆{�n'0�;t��u{���b�Q�@ޣ 9-�.	���X�F�ڴ=}����F53�˩��2�q^��%�[ptʥQ9�F������13ζ����x�%k{�h��jHu�dS����������%�9����u�:u��\�\!#gd��[N��Ei��{s���M�ˮў�1��x���K��m��L��x
UH�D��}v|7g�ʞ�>��c��V�uo:%i���o���MUI^<ɢ�M��U^��ɮ�G�"�л�w�����#/{���z|6J�ᕝ������W����1�¾�l����&4W���;�׳��;���ɟ�v<a��K��ʴ��m ��m߃�����zFь�'�Be��m]�T�'�W���O��Ne�f9�	�0����U��m +����6o�Oz�J��Z�B����&
ƶ��]n�� �C����0���st- �ҸA�ջ�(v>���!#bl�w[�r��R�[t�B�4��;j�`�<�헗#m������+w�dӁw'�f��bY��r�awC���E`
�vh�YW&����	�uע�w�s��cK�R����マҋySjY;�C����;�eV��L��wT?	;"q赻�����D9�\ܗS{-����5����vE�����Z뎝���~���=�^���Tr�@�,�
��M�S̽�~�l�]Q��g����$�$�:=�<��^H�V�ۮ��GA6<�_L^ڡ.n���\�zQe�L�u;WB����f�_U[��}��9�m������H8�`�,\T�p��<r#���st�|!��A���FH����]�5��q��.�����P��z��`�E|\����]D�V����N�];�Dm�w?;���9Q����t0�Ǖp8n!�w�䲀���f	)V�d�=��\Q�r�#L*$*ɱ�潅dV����q�Zq�u�I��tF\S�BQ%O �2���c�r�B���=xu=U�R�.��'�MF�p��F�'iC����A{X����ճ7
d�*:�q���f�l��,���z����q=��Rqdi�����[��|K(��K�#^D����?���8^O��/�T����8�;@����4�ټ�6�i�ଷ#H���3�@u4����Fm]#�@y��y�ʆ�-��$��z�Oy}s�S(��90��V���ǁ�̼��H�Z� n�"*u�2a�l�!�6�f;[u:�&��H�bx�ӏ��L��ҥ����:�*T�4%��������D;O��Ť��6ܸ��6\��)���l�W�ۏC�^2M2���[b_�TJ��T�ߣ6�ۅ�~y'wBw,>���V�������:Xɗ�R�;q��,\k�H5,���[	�1��<s�Z_g��ƃ������x����z��=��t��B|r9eX۹�~��r���Fd�دS�<���w���ӝ��g�.�/�S��iS�����9S���]D��_�R�W�,��a�s<�������k�����e�Wv]���eV'�<t��j��L�(�E���j��������3�c#xI�7FA�r.|���xYF�L�z�Ύ����N��P��n�e��wI��+��˞��pſ��}�����FYS���'�̱�gJK㴤#��C�yR_݁R뷷�{k7
"������,��+�vy�b"��T�~x����T��*e#}w_E<\�M���V?�D��O��ۿ�>��Jg=��{'h=>U��.J5�'��ྨW�H�q�|0�x7.i�t�}��)���-g�p]�xxU���<�%�ҝW�����r5�oXeZ��r�  ������¿��v��+����B:�Tc�5���Ð�79S�^�'s�%���8�Yq:�z�:^���՝��mt��b�I���<r+ị��g�N���C��q��T�v���1�M����0��UB���D�e\�t/X�v�n�ܰ �vU���+}qW��)�3�r�������Z3jdIgbe5]��E��]��ݰ�$8�����2��-��ވT�#��m�p��&�wgZ��8ncia��gݚ{�댄I��jH]p6���Ϧ��Ju���e����Ki��/����=���~�t���	�߫	C��(*t&�3�����D�^�����Wd���H;�r�~�v����0��]�l8[�rCN�+��_��_'�k�����T��29�T�D��w�.w�>�9�uƨ�.1��<���y:ͧl/�����:Y=@�-#�Ep�}�½&Ӫ��JX:���d��x�+�~��rwz}�-t�o.���{��ޖ�a�� )��.�i~tk��!��]='O�6S7��Q����k)�TN?��7�1����O2(�������h���<:�N'�pd�d�iQx��ǡUs���;������OS�2��փOuM�jK�>�z�d�����%p�z<Ȁ�$J*��\�B�r>{�VVMۙǺ�G�u���`��v��39 mN�ʠ�Q�N<�⸕����ze�)�+x�s�|BS���{М������:�
h�SN*�����A>��+��ߋ�L��9��+�����7� ��)ث��ﳞL��9}���|�#'��*�Q��S��О���T鸲��3ƌ�B�3�#mP	wFO���ק�23ۑ�;<-H�v�"�l�s��H4�1�+���vT���$鯤�4g��)x%m[��/;ck�\�������v��^���|�K/=�����S��� �.�砓�Gq[b�f��=��^��϶�{ �_�2I�(lw����Z�k��>��YZ}�C;~}p��k̾c�ۊ��ӗ
�7{�О���p� 3Y��niO}}t�t�9u��v*�8���1-6��7��8m���tg{��q8��w����]���AKd��'�O��P�Z�ڤ3]/'5����ͣ�Q��p�gW����i�:eӡ?3%�����t����mK��K������_2�ֶ=l�4�9uĸg��&� t�'˙�$F�
�tkX�Ƨ��ە깻��zZ�R�޷�r���/���[NK���p/�L��W��T��JgF���}�B^E��YD-��7��WF���j�ǌ����BsDp�އ ��ܙ��1L��#�����u3�z�h�h�S�y�_�����q�R`�V܌��1�^�ʡ�դ��U�_4;f�َ��.�7q,x#�h�y�l	�M�ӊ����e�ٹ�ܹ��?U-��W�Jg(�l�7����WrVɣɺ_����d�מ�N����H��w�����T����\>Oa��Ŷ��6������wzak�tS�P'^za���en��UZԁڵ�S�.8��a���L>�X�KÂ�i;��A߶���D5O}�{kJ��;_`�/^��YG����SBu��.!{�>7�N`1��amz��4��}�hWKX���	���x(���g=�C�U+�}	S�)���z5�p���R=},�˃0�k���]j�c9�gb�`���?gS=#��x�c� *;Y<뛓��O��\9���rr�'G��+�f=nm@��*t�I�ξ���Xn6��H�.�.�7	O2��)�Tfl5�B�:rN��V�@�F�C���{���|-��A�+�26�	Sk]XQ�X/�Y^-9L��ڸ{��S��o�0� 4��c�.�3ƴ�w �b|P���[t�O��X�Z���t�F����Q���^鞽�yӬY���Цه�=%�t��e �(�K��w��]µ��u�>ܫ�yFk�/t�~��uU���,W����f�7��X�1���+c���V����.ɇ�Т�pȗ��/��no��>��A��s5#��0���#��b\IN"lH(���2��4x 	z�XR��poh��_����lntMN���f[��ki3��x�G�p8[�P��e{0R�&��{��0rc�GEz�tx���eƵ�r�{�����놓~n�����p�J��� ]5�	��kjnu@j��ʾ���_��/�&[£y:H�s>��Ȃ��M�n�٫�2J@��ekq$m*{5���d��D�T�IZ|=��S6��F����7/�g��2_��~��rv�]�]^����R�!�����]6=�Y�,��gݴ��s��}w&N���U>T(�I���q��_n�p18F�Њ�$�G�z�$>�������V�����8�j�!��:u\�y��R�B/!K��%A̦X5�`�q�� �l�z�+���b���lv�A����W��V��"��PU����h{䪞��C4�U�[)����z�{
'��>	��9�
Bέ���2
���L�v�s�.�R'�;e�~�VǢUS�}ʘ֧"�����{E�����\d����)��j���ȿ��x;�Ua�['���p+�����gYD�\�{�ڸ��Yƾ����P/{�
ęzA�Me�d��N�]���g�T}𾓼�r j�o��p����I=��(&k�:w�`y�n+5ӛ�#�=���:v!�wS�{.J��3�]�h���w��&a�0��(�k4Tۼ� �BD6��\�{ ��Z��2,u�Շ�?&���l��P���*]�A�(�*`���`����g���O�h�<Vwp<�p�qv�{L8�ʝ7e�peT:P������W���1�+/���wU��������4Kэ:L��w\�M{�_˽R�A���B�{������EK��n��I�!�{�dꨚt#X�W�h-�'�C���MΎB�P��xP��,S�U^홺]��Y����%V��R���Ijw���Ϥ�kwl?@6JD�#=3�骾�K��^ր��62ﲬ>>���;�[���S>g��G��tG�:�g%�W���W��W�b����t�pG�G9�t�{�2��-���T�#��m�s��@Ϣo%��o��c�5(Z�[����o��~�`��L}�d�	<��zT�6	oQ�Ki����,i;B��=��1�H�e�q+!��\��e���L�����(K����ޚ��A�W�<9��j�O��w�6�y�a��rR�h9`kB��N�A��D��|_�
��U�V��r��PLa��dc�L]�z�����P7�f����X�p�!q#Z��l��
�ǶY�:Eٖ���4�ܮ��_w,��/�Q�)�u�R�֩�XŜ:$U�t��wMK<�Ř{�뻻`7ub���iQ�x�!��T*uŕ�ѕ}��c����W����q�p��s�cͪ�>N@s�Bv������k��<Y=��-%�_��_�K����!O��/謗���+
�߮;ܝޟB�@:7�ˤ+|����q~��K����zg��lggb�QpvX�8�X�}�OIӚS+�m���J�xc�G'���Q9H������y�۵�߷��6PG���,~���]O�࿍u~'=�H��r���
�g��	A�sj��.����������W���S��?�`�yQ?"�ݧ���K���`~�.8��/x/Ny�C��^`�L�S����p��T�,�����f��W���o�w�/#\���X�T�@��[<��A�w���ҽ|zdn�Βt��y��Y�ζ���_��>�v������mj��ᮞ�����}>�v��*��Ĭ���j��$-���f���I�3�$fT;���Gz�QT��b�oO�Iei�F9�T,�	�͈�9{=�y�?��x� o��:@-)���ϡۮn����:ZN���Oէȳ����]#\lo^�^27��q&�u����6�`�h��I�M�s����fV}�f�<:ژ��ĳ��_vtY�w-�$���4�7:I�[���K�r)���	��ҥt��ܰx�s#˱�q�col&��7�wVNA�	N}7��w���ҿԮم�%����Kd�A<�}��(r�\4]uU�+�����;��{��9�7!:�&���7��M�%������:LL�tV��l�c��G�A��,cwE�Q�lc���5�4\rj���]q/��M�n�v�&�L��������C��I��Y��8�W�ꌅ��̨�-r˩�mN��t���^L�}6�tM��ޯF�ٌ�y�m.��Y��TD�X*�3�{Jñ�.�M]ɿ�JdѸM���UC�`Dfƈ�9q�)��n�n�ۚ�.Ɯ�������iذk��/=�O����?����)�������~3y�Ӳ���,ޞ��؁��2�+����r�'}�����w�������|��Vtӎ푊y��=p��XWs6}��s�9��W��4���2��]U�7s+������1��.�Cʩ����X�>ו��/�#�,��3Ƌꅋ�.h��S�2��g*�f�q=(�v>�.y�7'�c�mN���g��,�_DH��طs@h>ɘfdX�wR�L�5b$�uvl�w����>�u�[�,�e;ڛ6�$"j[��&�k6�Pl������j̤uKG7�ks���٬��X37Bdy�Kq9�f-�oX�\�(u*{���-��r��᝵1�t��}�',����l���ɭ=S�O\��Q���H�q������2�Nь��`�5����>�C��)� *�˜�}y�^a�q����D��;W�5��i��c9����q�S�ji�����,��)���NLY���
���0��@%u!��K9���Y�O%-�tl��v�UzK�^��Jܼ��X=v��b����������@���X�\lne�k%�6׋6dф4���ߴ7�ʚ����Q\zu��ݼT�Lٺb/��#ovbK�-h���)!ޠ���D�X�6�( PXBE��囹�2�����I+[)�{XE���l���Dq3��/0gd��瘖�ޮ]<غa����C6e�4L����윲rS6�#L��T&E
�2ι�m8��4_[�s l�Z&	����չ�q�|����Eg:�E$��tº��KG��kP�;j�C�FoU���V8�k@�����U���qL��qt1t�g�@��������j+Ѡ���[�V�?\��"�z��|,����e�V�j�3{�P��5|J��XƠ<�s���ֶ,J�ٚ��]�z���)��0r���mͮ=�Ki�6-�r4�$Ш$i�+3��r���妻2pȭ�P��q�ݼ7�f�Mt�-�Rܞ��}N�>�M��g���i@�:���t��Ӕx.�wr=�A�dC�0��m��2�=����wqc��tZm}�mK0䏼ѱ���,�Q-8���X�����k%ĳ6��+����b���
X�#h�9����z+o}���l�AveZ���k�tvs9+	����5���[�����;�>yİ�=�Ʋ�r��^�ř�G����:p��E�#�3W�+�Qgl�ɝp�:BR5�����Y�yҨ��v�r���j��k{n��R�5�^�Y�_S�r�W�PRi�{m��8V����/�q$�k�|�-:Z�ݙΥf�i�[�j��n@ ;Y�,Jc�>��Ga]Ek��*�<&�W��K+) ��2-�CҋadX/s�o���N�����v��G��V�T�.���,�e�EFƾ�Vb��:�G~˧Գˏ��v���*�#i7g��1C�է�i��k:��ӑ�B�to�嫢�%oYb9�vf�f]�6P�t��Z��W�(�^�b,#�r�c��)�l��F��k�;�I��Y�v��UCZ�y�lw���y ���^��5����ѱ����(V�s���{}�݊g�ᮙ�̛�݇+��[W"�{z��CmfÂS�.��v�w�z��Ϟ��Mq\W�+��䈡�q���9��B,S"�4E�
�6g9�!Hs�PYH�82r�(aD�X!D[�Č���&�����̓h�DDS$1\�đs�Db͘�b���&�9aB4��r�!�2#7ēI@�Ps&%.8I��ɒHqƆ.8�2���f�4ē+�Fs���r�E.r�1�PI$�s�I��q�9s���������23�3��B`"\�$�i@$JF`�� E� ��P�3DQa ��b$ɽu��}�{��׭\s�7� ��x��Sf��3�ɥ]R�a|2%�nS[{�$��P��l<;�-ʚ�ͭ�+��d����n��յL���v\x]2m)�^�����36�!����5��%<{�U��ܟ�I�X^�L�w2�b�mP�+\�]5����Yx}	�g�ŽnM�B��������/2��X�gb/d��� >(mOW���r�Z��]��]�G8ܛ�дq��~��	Ci�gm5p�)�a�IF��OQ��=Ċ.R�멉r�m�\����rv:����A��x<��G�5�����p8[�P��rY��7��0�L�I����s������g����t�LmF�p���\����>��q:��y�#.)ݡ6�J�� ]=��U�^s����yo__v�
ٰ`yn8�.+xLf�v�dޖ����7^]U�P��##:xz�lg�CWev�'B�{%��
s½+N�i���-�Q��]nKe�,���d�r%�������|�� ��$R�S�	�y�¢T�4.)�a�����>��9~����S�f=��fU�*��3%����L\ivd����zam���+��z"�S�wY��zn~���
�䚦���VO��5bZ2դ�D����A�]��M�������n��d�;U��W�/"�ER�-k��kQ�����p�wP	�T��l�
�ǳ�a
,/u���h[sŪ�kƳ,,e��̸������){�Mw�82,�J�лk�L�m����<���~N����u�𡑭nXٟ����A�]+kc\Nr'�x�q����U�sث��[�����C4�4d�Oj�]̋�FJ'+�|*㘘c����U���C�{xe�����n�V���W�հT��;ʘ֧��ۇ�����O� �3!�S����3�\��8�~5g��Ua�'�<n�@�Ʈ��5̲r!��=�W��3�/b�^�Z�^~�®g���ˉ�=BgGIrpdA�A��J�+`�%\��^gM�n���5���7}	^#S��kL��>+����Ji~�>��^4��jn���w�>1[]���c�r߁����t��C����1�.�J7t���L�A��.�{��{=O���x^�ѻ��G�����]��_��l��S�7:9@�(�:I�0�f�W<�;�t�������q��޻�fխ���J�CRZ��:i����˄��~��VtJ��E�K~����>�j� nK��'����S=�4�o�*��>�S>g�������܌�R�EEL���t��C*I��0��vvK�{�[u���=�.�67��;D�A]�ш�b;�n;U`.S8}}GfI���ԗ��[�����-�oR��8��qr����ɔ�"]�<�i�Xȹ#�A�bT1��*%Ym�����S��m����k��ҼH<r�ÿ�H!*�`&x^�\moW�*v��9Ͷ�Z��m������1��*�R�FB$���$.�DL�}4.)N���2¸[�F����=��Eϣ���y�hn[�Ͼ.q���zB�Q5�T����s�;�+iѸ�+�iO�j��SN1`��׃�Րŷ�r/�2_�9`kB���O� �GJ'k�d-7�~���IzyЪ73�}r�p��ue��*�����[��]�t�N�_�)��wR}���V�9��d�5�Y��k�Ά�g��{[^t�:����Q�]����?mۣp��
�B{��3�����/����^����}<:�d�W�c.:�i:}���m����*i�G'��yz��f��q�ɱ���j�!�V�q~�a��ߌ��G�'/�?T@����N�]_��v������`{���}����M��XQz7��-�j=����^q���ÜQ9�az�K��zk��@>��8AC�\k�p��=Ʈ�\���|�*\��;	�p���T�����3�
� ����yߓ��r���#3M`��*��Of���ľ���S*�S4��'����X�&��j6'��X>9מ�N=�u�]����a��g'����7��"����c�j2#܏k!M�#X�T��9��&6u�>�u��z]��Z�VJd��
�٣��}ճ!���nq|�H5��7�J���,˒�@U�8��]�S;3�3��f�2���:T��U�x�{%����}>��c}��_���~�f��3ٱ9�z����N8S���3�L������w���j�U��oK�YXV9���n����;:�q���9�ip(s��2��<��߯��>�n�U�w��殫�f�ɾ���{c�헾/�NF��;��uH��%� oT�)l�d�������~�S�E+v?a[�-;C��m���u�M�y���]:��d�\D�t���u�hﱍ�}&�-��6���T�N'���W�-���5h{�.����&�7X�w�s=��H��]
�a�����J�V����!��ר�Q�r�j+xLb�]nM��p�1��W��UHyӔLU��˭�x����A��zn
�
�[X*��L�핦��\?&����L�7	�^��={|�.�iMUy]9qҽ2j!�#�P}(m��;��Â����Zo����N�\�]x~k�a~n�9E���c`F=�"xGl�ˑY�q �,�z�'�Z��X��E��井����$8���F���u�N��˲��X_wt]��#��xq��ܶ뻜�h%4ND*o={$�s��֫�-y��\��ڞ�ے�L{�E(}P�N��'+�7_���d�����X�T�8/��ZN�6�y��tj{�1��El��!�~�R�F'#��by�z*4�S�ƖN�!}@D��VW�z���X�{+�距�<}J������u��S�)z�M���pʹ�~����u���u��+����ٰ9�ˉ�����D��S W݋���u���wQ��ͪ�ވko���>���:�iy��#3;��(S����A�����W��p>���+�.�7�S̽�������u�.�\h��A�Z�����:^�'k�@�Ф��j���Z���t���Yx^����U�ю;��yV���j��
�qC�e�������'��{��~�8�?'��[�ct����?Fy�XqLg��gnWB�f@��i$�A���H��.����ή���D�Gfǵ�Ӎ���ԝ��[M�t0�ǝp8[�P�eB"�|f���sރ*�Nr���n��.	�+ށ�����q-��yϩ�܄놓��ڟo�}x}�=����z{	q<����˟��/8_�=��#]�z���vݴ����ve[�j�z�Y��]q*ф�2�î��*hڄ��`X̥3��
�;�?)�h6�Q 6�o8�l�m�w&�q�KW12�Y����U�F���R�#E��1�g$2�b�2u�b��ξ�����!R���i~����������&��T���n�P�xf~��-��fһT�8s$�_mI]6vH�N�U��+N��L�-�Q�u9=��Yھ�<�]Tc�IY�;nF�ϖߥ������x��/�T)W;^�Y�qN{\v��}Έf`#9�s���j}C}Ѩlf?I��Q�ۗ^h`����*=��X���-m��b��潨����NSO��׃����'wB���s7�r�;5�/_�A���酰sr�hU��S�w�KAwR�X�M�e�q]�L`Q�[����-t��A�N�	�X��ީ��Nu�����m����N�r=��}�W�q�R�>���o���_��,b�s�������B�nu�9�U~tpY�.�Ӆ8'l�����V9��`�T
�����S\�%��;�	�O5/�j�Ny�=��c�⵷{��0ߦps'��(z�Ύ��tp_ƕ�0�;����
{OWU��^S]���c���t��;��'zȱ�jx�~%(./ �<\X3�6ڠ��ɑ�f�ʌ!���n��V����;��5��2�=D��u	2���j�Q�o�������wm[�p"���+i�ͼ�S� "�s
]�-`�����tح���IS�h�sM��U�K�쩒��b3\۲�A��CO@�`]������^���;m.�Lg�:L���׸��Gl�'j�f��!$Kz���p��M<�uE��h�����^�����|��m;A��W��F��O,����S�Q>����X�3�Td������K6�m�\�o����9a��G�wl>��b �+�o(�����R ޚ�O��H��h.=
�\U�w�|�|�i�NF���v�W�{���{ܤc�W�o�2�4�L�� %Z����}�Z6*P��M����$t.��3s�w�c2������o�N��ӻfE(��RB�DϦ������,)@�}��AΩ��͋uk�����a|���|\�%{������T��c��
VӢ�����E�̛�Uln�[94�0���O��\BJ�/�,~�� �ԃ��D�} �Zr���E8�C8���}=[.�;��}E3�~ˇ���ښ��y:ͧl/�Mk��U͐a?U��>�ׇ���vJp����)s�9���9�+M�o���aѸyt�n�ܣ�x���^��l�7k���h׼���
m����hl��p^oWW|�	pG*�r��/P{ %N�N�oj�o~�XS�
*Ju�c��5�%}��1N��խ\]����Ƅq�K��-EƅN�֕�fR�����t��"ܴ\�՝�r��u{�;}�_�X�W�|���}(u�����Ǻ�a8{��L߶���%M<1�qGŨ��ʑ<���b��w�9UD�~�a��>F|x3��L��0�RnO�A�����o��N���,���G=�05U���u�����}y�.>�z��Ne����K�צ��� �p �V�B�Ǜ<|X�:���sϟ�8�+�N�n�B{\/��T������R78�����&�u����z��/�/|1�"�l�s�ԃ^w|�J��eHؖ=���D�P��o5k�M�'0��r��|n+e�(��w
5����e��}>v��ި�3U��S@c�{3��8��GN�N��C�qS)K�]J7
�X���ޗĲ��=��V���CWfyo$x��u� �����My�Q��(	�t�5 ������>�n�S+ ����ٱ�wSݡ�df?�V��z�;�ˊwh%�p 5
[$Ϧ��L,��}&c)WG�C���x����5h3{LgCu�M������n�n��v	�i}U���h���h�̓M~]��i�>47����o��񷧰�=C�c�lIyv�rc�(r- ��E��\a]��։�~�L9/�y�`�0����C�pt3�Bw�x��M,�K����1,)(�̡`�3
M���C ���u
H�˵�ݝ=5ݙ����/�G�����qɫA�<KP�D�&� t�'˙�nU۔[���7LfM��ǰ�
�T\QCәQ��rB�o�]nKnx��_�*��W�������R���g��|l��WҶ�U�Jg(�l�=���uS+
d�^��"�H2�+t{y���:����L�0�N|}(m�s����[l^l�+j�:=Ì{e���W�aw���\g*�QNM��v���z_���id�DL.��e`R^	�8N$�lN��!:~>�ߺ���1�c��C�%O}�N��Y������X��T��3�x'�a[����V��Z�귖s�,Ү=�hx���T��%O���������W2/�'޺�19w)_x���[/�G�z��z��jZ'�) ;Q<뛓��O�Uü���D�u==��v3�7����\��ġ`�@S��cnP�4�
��d�JS:�a#������Ⱦ�����k�d㋷��J���MD�'���%�Қ_�V�!*uk��t���A�QG��똡�:~(�_2Ƚ�p�u��nkB[؃���;㉫E;�V;{�fe�X�� 2�^��4�x
���4.l�)�$�An��c���@J���Z���5ʵ�%��㒻9(`v�� �Н>���p�컊F�U��4�+��f��i�g��\=��W���2��{$����<�e=��򳷏$�-����Ƴ�z�mЧݶ��.��Dc�Φ�t^f�zJ5�'��2���H�i�Ex��7v={x���e�W���Q)S�5Rw����G�5���s���N�1rY�D���ޮ,���>�ʽ���<�
+�����/�P��-}qW-��3r��'\4��7Deû�*����i����򷽦��e� Y4zH��Z�+K���B�-�Q���}g�[8^��X��o���~�ǽy���x�Uh�$��'�M��"e:�W+N�S<��F�%������wK@
q�~��{
�^�<Ys�O{�k�R�D���S�	�y�����ȧ=�����p����hsqۦ��1~d[k�����vd�r�k�B40WO�d������?a%���8;�rX�:#�W��2-X����Xo���.��A'UC���s7�r�;5衮�A�K'c�;W�$ɏEQa����ٝ�Ia�q��on^���Ƌ�߭��^�k��[ʰ�g��X빑y��o�x�P��s�9�1�h�2��y]EJu%��ɮ�5yE],Gb��Z�m�Ey�7��b+8e_(��������2�c.}:�^��ݓ�blL���b��ħ@^��B�����@T,ej�x�[���rU�T�{&����3�N2��ڻ�1��9-�JPͺ�ި�d�7y�Au�a�ia���%5�&Bj�^�����	�5��u�Ҭ�����i;QK�o&��\�m��4w$��A�X��7�LA��U����-I�s�����v��m�Y����&-{�u9y;T�-2i_�]z(�e���T���3']����U��Kf��p���Y��������'���ܱ��Y޺�������>���U&���m$�;��/!�\�<�Y��_b>�W}�]a�c�{��Y�w������(��z�µ���(��p�x�u�A��̳+4��0WS�L	�-��J�^�r�lC�@��GM�Vhؚ{��WO�㢨*�\����(�X.���Y{)L[���̀ԡ�7�J����2X��ɦL��o�$���jb�2ә��Ls�>�X#�ÈҠ��n] Ū�$�d�3�<��X�(&`��cl!��gc�q���̮Z�ϵCt�R��eۼ���/8*;��v��������BF�1��3%"�YU��ls.�Ԧ���';6�ubˌ�61���x��o��PDqT;atD�&�9�VB�oVtr��U���g��w�0��HC/�4�L�]��rlbm���/F:,�����(��r�t���R[s�%�\����1eȂ���m�Yl���ԡ��MR�:]�&9��	��J֢��ᓻJR񾺴��R��:�P�v[G�%�K�A��SYΨ��|P�v
���kY{�Ǧ�)�5�5��#�,���ތ��!Ow��4j�v+�F�����]"�4�6B\�(�S�/Meԭ���.j�i����.v7
L��a�\���(b�d��!��Յ����	�9I]��X��b����3rw�s�5�C�n�j���=RXu��e*]�T�"�TxsV�W_`�(>hU�mQ2L�r<n3�>;6�8��3�fa[��(��/y�0����27}�;b��8��#"��d�H�a,�tD��r��ܚ�J�L����s�SG ù����i���KHf�i���!��j�
�Qr��u�f��17��]&����o��w��-��r������L<�L؁�v��D��δ�C�Sj[�˜��X�M#U��3�)+=ٳf����	e�M�N��zY�2�Sٛ�ꣽ�� !�a�l襇22�2�-�-���mm��<�b0�b�b��-H�K:+s#�x�Y.�{�u�[� )59���c�{�{Y|��f���f�feGp�p�b�$�!2m��F�	وDa�*��|*�BR�H����$�&�$L)�`R�L`���BD��B"R�D!H��9\4���"�䘍�"�#"(�i�E3"�$al�.(�h�)QA�F�$��"�$H,�$	1C2MQ�#Q�2	�Ƃ$B�)%%����2��KF2�1$��Z�XH�ȰI��21Jfb,!��cI��(����A%��Q�!��a"�0��)H��Ěb�&���E	D%D�Lb#*b�`�"�L� �E�f��0�E)�Dɱ$�+$b�C,`�����P@P��3ض^�˫Z�f��_b������7/SY�G+�!��06��+l�+V�KB����`�3��TU{2�ձ��������̨W^���K�p�#�S>��c�U<'ܩ�js�wPw�ݑ��2�U�#|y%�_��Ł�~�ÿ�~�~:�`5�<��0��\?D��e��sW]�£<����)I���N6�w|�Fƛɜ��8rR^�Z:5����1���^�r����(�ul�4mn��ý9���E��y�_\n�^F;;*t�E�Ou�eT:P��|F_��`���Mz�q��[��Yc����Aw�+`���Nyn��)�q��2�$���L�)l7�M�� �S��w_o��i^���~�yz�(��Þ�l���Ӵ���<����/�pF}%�����ޥo�;���'���F_�`Yv'�a��~����RZ��c���>�2�}�X��3)=�����И>'iHzj$�&U��;o����EtKw�}��=�11��eX�M��Ȏ�����9���SL�|�AF��Ā�U����x{�eq[��n<�ad+��3���g���s��9��)���v̋�2Q����ѲA�htE)�r{�M�ܫ�u@�O����!�BlU0���Z����x�PVJ�So[hȯ%g^���º]�Ύ#�{Q���mO����'c����s����xk2�A6�q�Ό�]:�[K�3����9��c�D�����65��R5}'V��@49�m�ou5��O!|4q���u?K_��E[2��+��+�G�WʕD��eI��L�8;f:���x�m�E����U�[Ψ���ɫ����*!����E�$���>F��R~�(�M#�]y\��=>������igި�n���r��p��s�cͪ�7��7	�K�4=3���U(����>ˮ��2���� �}���C�N�M��|~G�zXμ�����宀t_�����������q�7��zmЮm�_�_Ѳ��<X��Nq^�3�V���S*=���(�ߡ�[�u���yU�ձ8�?�]���^Ӱϑ�\Y�?��,�ճ���NnT�W{�.8����8��9� �w�2��g����neN��w`�~���{ k���z��':�
���s�9 v����u���|���t�^�\7O���q��7�Yd�tnP�-�!Y9bs�h���pQf}P�"���T^�mPaxcvE��nw���;�iW\M���a{.⟭�᤻m����	8jK�Pg�ї��e@(��w�5����7�kߦ?��s��c�W���34�՗0LS������Ȳ�!e��Ě��n��,I߻5!D���*P��"����B��/Mo�	Ы]���[�8v�c8�ϲ����@��-���_1����r�N��XpU�Nc���N���,t�^>l�M[�נ7q��w��Ƈ�K��P,��tv�PT+����.6꧍��X�j�������{����wH=>f�Yp��v�<��o�י~���P���jiO
�Ρ��,Uf��>�gTV��m���k��Y;����N�^%��|d0
[$B���Uط��v�fx�u����΅p����ա�϶�܆봛�wM�;w�(��_�}O��f���y�:��z�s��0�%�z��e�	�����qɫA�<KA�M���ݻ��=z��N"-����o^����H�G������*�v㙸\�F�.�&�\�L�z���u���=۩�Wn�q�\9�3��llJ��W�T�r�iXw��ɫ�99�$d�J�(���;v��_�M��ઇ���~�<a���P�|���V-�/6V�����Y��x}��Q���������&��������,���]c+�����_�p��-G��ؾ���D��\���c��=�{��}f��Ǚvl�[�8����6����?�3��a���:���b���b9��[��+�OXkod{%OQ�ܔ��9��gsF�r}YJ��z�V�jF�y�6�-h�nؖ�M�"z�
��OG����z��bLR
�!�`I+9.L��y��I��U#uڗS�[���g�����\s��5] U�VǾUN�r��V5V;���p���H�����N����;���k�$���ΨW^��f�2{�2�ܺ�<�Z���b��j�t�6�LϤ��:����nOA�b;���O�~��+]t���3풠4F�x9d���e�L,���#������w0�㮡��{�5����I<�����z|��ʵ����u�t|�����5�/��
�;��[TQx|ܦ{����|U{���e�A܃(	�_.*z�{G�x�M4U��Kx�^;�K��U���VƏk�Hg��tۄ���^f�zJ4��z�2��+��SM����G۹��I�����먖�^��;��ki�ٮ���a�w���������HW�ϲ�� n {%�%3����־������n_O��<W�a�G�s��zo/)��u:�z)��J�� �_iV�p
����.+xLf�v���g�[8�:h�t.��7rNL��J̗��ko S4�d)�P��+�����\*J���2���b1����)͝m��a���v���)�WAZ&TynS� T��&L�bv�T�K~���l>�7~�g�r�%�0�˅�V/G��}�m՜hɨq�L���wY+&^ ���M
�%�����X}p���0�E�N�zv�l����Ai,���/�v2T|8JK����{?2Y�8�hM��m+�T�ٙ�w�¢%N�B�)�a�p�g_V�����}5p�-�y��TC���L\BIٓ7.#���:~�$�d����'�#�`%~�K�+ڛ�_�]����͖1mU�
wt.<�3m� �W3]ԃQ��ۤ�1��1��;<������>F:�f��V�ٽlh����S�ռ��|�Մ�w��2i윖�o�\�p��� �w9�
��S�$�'ǰ�T{o��J�xO�S��fg�Jo���Տ����򃰟P~�.�W,X��;V}�s�]z�M�L�'��J�Q����+��u\�U�mz�iqq�՝%��g�	���Ds�ギgs��/�=��EK���*�5^$�[yB�q�Gc�XuWvBށ���:�T�P��7}	�#ޙ�A��
�t�s(�m�l����R��:�����l�K�v�C�=�	�g�����0��Q����K�jd{��K�wE�8(�3��q2�������!{��|�Kg1��U����s�X�v.-��6�x�0��/fE���`G2f�f�`���!�IS
1�_�q�V��;@R�me< ��xݍ���tG+�A��(U�{+3/��&䘖C�F2+u�k�3Et��53Ho-�Y�ĤU�:�0�6]1-6��լ���*�Y�MX�"��{�@��[8xa'Y���}P�(�G�޻�f�Zۊ)S�֤�;�tӓ�'�4b2k����ѝ�{��q��~ĺ� 騒���@�{��갸�}QE��-
� q����:̧�ǟQ�	��ֱ܌�4�����=Q2�	V�`�x{�eq>���j��K�f�x^�[��Ҷ�{�9����p�M���v̋S%�B�DL�}4<~��$W�zJ�w��9°{�F�]l!�r��>�.q��G�WʕD�q�'n�s�Ժ�x���<���#x���}fd����&�;ik����'�r.!%L��偯��x
��p.ڬ�hz�d�����~3��|Jp��u�z'����3�~˅����o����'@9�N�Zb�oO���9՞Nj�������i�'�����9�w�[/���)|lg^XI�U�E�ɫe�����~��������hV�9o�_�\l�x�A���2p+�S�+Iù��ނ�9�ڏL�TN0�yg8���rq8�(}w���y���3���O�e��'��}GW���*������K�>n(�Xi���WuL�8X��}�Z��,�X��+d�[K�Ցs7���/�v��Tg)ܒc	m��d^\�Yy�r.�/�#&�	 /g(���&s.u:�
ރ%�������I�5VE׫�
�1��w�띚�3��fO�&�n7�6x�:&�:@T^.�0�W�!��:ӫ��j�cs*tߑd�ِ���6�� ��kg�ia�����*@]�v+�E�>~`���2��:�|���;�:ft1ӥ�h�=���=e�ꎿ��W�t^��A���g��w(>uZ��;�8f_�������c��,�w:I�Bg�z�\Q��h����w�]<>��Yy��Q=�"���z+x�no�u�����R����H�$�L�$>�WS)L\m�O��N�)��S蚭llw�1z��x�>D#�Ϯ�6��liAz��8�7 ������$��߭�·��Y}j�U���k]�9�a뇎�r��0�.J5�Axʸ�Ku�sFk�ի�C�{T��q�9k�;�ա�>�cr��n<���qN���2Q�ꑹǹ���<���bk��ΗG�G��������|��=]q/��D�&� C���ߞ}I����^���f�Y��̩��!#gd��VӣQZr�7n9��Lf��ro��p.�*�b:5�6FV��z�M�� �ša��������κۏU�k\յ��Rf"�̔�^Sw�T	
<�,��u��&�V5�a��ͼ=�#�H��� �����uű��o�c�L�u��]���ZR�CI�3d��q�/Q[|�R�`'�#^�6�]6�t\����𨕵���3�{J���P�v�b_a^��Sݱ�lf?Iq�[&��n��ઇ���]0�MJaσ��Â�m�doa��4���s�>o���]��M'w�=��96�\	ۄ�,�ѥ�ύ�d�L.����Pe�|ϧ�+9�>��YǦ{k5&��O�6�w�����5O}��r��	ۅ����w�Sド��ꙍw��3��ޙ�׮=��7�:��R�%���`
��cЪ��>��>r����}�+�Y�V��Ϯ�^P/G��ӑMN�A������W������@�@
�.�9��wQ���q�L��z��<���*=��_�_�ؼ�����Y<2�exѝ��u\o�P#K��0�dϧ������oݳy�\�c�����2���u�Z�8��5u��󠖏Ji~�R�g�^G�����zimL�b�̔�{O
r<��@�ݔYX|ܦ{����^�h�F�d��P⇥]׎V��ʨ���O'��e�m)���V+�0w����t�M\=Fm�|.J(i'��}=f�3��0+"<"�����;G�Y�\��y�,]
�4;0�ԉ4N�\�U1��i�C�Vh��������L�`��j��'o�}q�h�Tf�z���ʺa�h�/�}���U �(m�[RU���M.��M;Bج��1$�����u���Z�ni���uj��˥�z�%ڵ�/�I�C[M�t0���\n��C�J�� g�'Fs_[:\" gQ����>'��xuB�k_\U�-��z���높��:Aǚ�\�ۙכ��{�����L��� � �J��V��}j�[£n9;H����W��^�y��5ݟqq�`7��ꭚD��I+g��)�
���h)�Vz�)yd�s=��r�tzÎp۷%���W��2_�� �"G��N����v:�+�S����ߦ=<\K��������s�����Έv�]ɋ�$�ɶ����j=��d����v�zam��~����+.��k�wU5&����)xj����w]�!���t�e�sa�;멃��%�VSȯ���f}�>�S����9��������F�����m�����Sҵ�f�<��j=���[�zQ���{��a��R<�'�,s#ޘJ�O������v�g�]L2�K��U�f�d`��r���v/�-��;ks�/�����t�N�/��a߫*��2�% �����n��Z���.���dս\g�ܑ���wF�{�X���&�c��ה	���K��ӻ�W�io�Y�xS=$y�{�8n��F���nKk�8���o�iqU��k��D)��)v��k(��Y,��<��vk���2d32@�â�����V���br��Շ�Б;�g����}���
����ˉ�=P&tuԺ8��_�1Kћ��y��x���K=(�*�TwV���+��z���u�c�;*t�d�o�P�,�<��t^mն׍�S>�{n�+�6h5��"ևLg�:L����S^��R�~�D�~�՗����h�ĵ�&��x�9LI/�F�����b��x=D�sю�{i�N+Ԣep�(�y�[�/��c��<j8�'��8_T+�(nҨ�uZۊ����h��2�q�����y�r�}�6��vyt���
'��3e�@L�D�v���aq�+}qE��U�~瞭=R��B��(�Ұ����eӫFmL��@{&@r��L��#{�c}
}�dw�c����T�#s�m.w	M�m;�dZ�(�uI��Qh鉷�Vi�x��hJ>G�-�#m.���Y�8�P�.B�Q5�P���<�%���c �G��k����z��ݓW�P�z�Cc�Q�~��9緝xz����-�������ֶ����[[F�ڶ���Uk[nV�Z���k[o�ګZ��Z���V�Z��j�km���k[o�mU�m��j�km�j���+U�m�����mU�m���Z���6�ֶ��V���Uk[o�V�Z�|�V�����
�2�Ⱥa�����������>�������� U
�
	  %P � :��!T�"�J��P�)]�
�.e� QJ���I(�T$� �s�*��몥���KYkc6Zͭ3�5m���Esb�� ��cƫp r  	  v8���n�1(ɪ��A�-�EQ4l��%!��`�i"�T�Z$n8��Y�����]ۤ�HMV�X�*ZʔkI��W �WMr���ʶe�)w8�ZJ��٣V�w+�����I���U(C0d82;]ۉm�!ws�G]ve2]�NB�b�3 �C�P\�J��m�,T�i��Ŷ��١d�mSi�b�-��Be�+��J���E�*I2�il2d����ld�Y�T�u�FlRJ
���eM���"T+mJ���Rd����j�i���M�i���+@V      "����RT��4�� 4@E? �)I*4��@ �9�&L�0�&&��!�0#�JT�hL	��`Li��&�&	��0`��$�@)D�M	�	�����2i���?������c�����޹�ֲ��B �l?��Q��@ '��%@!  ~	 	a���XB � ����o�����3�T����C�0���	�  �(@�C� �B��0D �2B �C������r?���'�����  ��I�/Wa����ڇ��s�i�?:����((�$_�Ǿ��Oݓ%�����hv-��N��ԽT��T���ݵ�%e�J�n<X4n�1ۄ���>�.݄nf<�e��Tvs\;ZC��M.=�,9KyK�gk�/Kh���%%���J�1Dd�V��dR��mіͥ��sv�] PG~��ނ�C�AkN b�m�
�{��aF�����f!K%�Ia�L�p	�+#6ڭ��Dn�Jѽ�ח7u,<�i��׏�'1yF�nb��n��å����lӒ��`$���.��ku]��M�sw�n�.�Q�1ŲPط;�һ�v�����ٔ�2 t�WGo.�Űr�Ғ��Z*0�ͽGm��2�[�ݕ��AfE���JR��ZU$�9�Z��t��l�;2��h�����6�_�J]J/$�V����Y�E�e�&�4�j����2��B;�r0v��m�I+]��`
El�ٙJ�#y�S�MQ������8a=ZZ�&�������3W�S�Y�s	ȫ2�tm�S��٣*ﴓXE!�J�sѕme�.��,��!��U���ӣ1�4���
��E�!�&m^�t�7p���JD�6�B��2��.3�(&�Po6��1��DaۚND�9]k/ ��D�|�c�m�+�C^b�qՀ�fT7�Y��)�5u�j]�v���:������t�Ҳ��VP�f�.�X�Z5��"ś�ww����{S�	[bm̤��-K ��N��Э�M;�F��n��ؽjQ��U��W��B\w{�JF7���*��>g*�ooek�#J�[����iIرZ�F�]�4m4�m ���7w��	j"6^��F�w�a�z�',N�
2Nn�a�7F�QU�9�-���2*(7v�����0ڷƲ��1�^g0���}K�|oOv���Xmi�ƫ��0�6��1FeCcm��*qhKKX)<ّm��(-j��T�&�A͘غF�-^U�؎	Kj���eHu���x�V�a�GWy�֫��mn[��bK[K
L�YE�m`#��a�pXEh'l����|�ǅy��X���-��ɩ���sv1���@���)#2��^�v��e;�ʹ^a��I �#�*b�2}�B��@U����x@.�ɢa.fE����_�A��w��ʆ��d�%�^Q�ZV��e5���dc6�\F�Vq˕��ڨJ�r%#�'e��yZ���v�cq�N"�Pm"��%��b��­�D����p�*�q���mA�%V�*�n��:ݾ�,�f-�wv��V�Lؽ��<��Ҕ^�X���)�76����p뗆֫��	�sq��MPY�Z8w2!W*Փ�"�.Ռ[�6�L�{�nj�-f�E�[X�$A+-e �M�2D�Toe�� aݻ�Ә��Yb�������kkd�xm�^Fo`S$�[ӷ7�Q*����%�1��{w(����y�����e�N�U#��Ki,���3����4��
̰�����*�'eZ;+N����$%<xA6�n��dY��S/FX�ӹ(�xV�g!�G&c{�+a����m��	��)����Ԡ�*IKn����q�x�t��iX�V,BK�yD�,L���W�&]l�`<��jyz��Ȧ�y�(����ť��2�CW���0�2�a3v�Kƭa���Yѫm_Īum��r��ju�����j�ͼ�J�s2�ڗ�����K���
9O7�$�Y�t:��ַ��N�g]��_w/�P45���W����d�p�j*ֆ]�n���`��V�{R�;V,m۰�P�]�����*��N��)�y�Z�cd�:�2% ��,�RS{v�i��-�@�۵tZ���մ��Z�O,}������LmX�uOi ���^XI'c)`���mc��+������kU���ֶ��oqi�?�^F唬�Z�a�9�7p�I��/1�R���
åSR�Y0�f���e��;(F��{�b�1�p��lEeH6���[�%��j�p�[EQ6]��ȩB��cu"�ͬ[F$�q,���M�Ku��/,�
f��(��L�d�X�I5�Tׇqe��M}�����8�I�4��C]L�B't��P�i������AyW�J��R��`F�^^Z����6�f�����T��ֻ�.1`R�O��4m��Ua�c̭��F��®P��R�R����ЫX�k��q�Ҷ�:$V-^ޝ�u,`[��f�^��-���|��XW,��лRVV�8l�,��t]�Cyۊ��>��v�6,`�ʺ�s0,ٻ˻O�I�|͈�o*%&�rj��!��o59c�*��!�kO�{r�LG���L ��-.�=V(O�)����kr��D.YWz��a�ѸVM:e�%юg�*Vc�VK��v��e�L/X:��V�y��ѺM�o]-{����;���f��!|Hq���*�������F���?>���n��Q7U����}�5�Y��3����                                                                   ?T  `                                                                                                            z���HÈ[Q*�l��V㕈�������r];`i�h�b��{ՙ�0".S���.��^vC/�|�e�y��i3�� �.�2��A���V�J�mmڵ2]Z���1v�f�Q�|&�n\.��Wy�̠ުG�/z�K�]��<�j/cL='$ ��]���Uo;0���Cq�j�LR���H���%#�ւb���D�Ҏ���bPܾ[ф1�&,N�Z{�K(7�X�;�
�p���5��bX����������S�浘���}y�4n��4R"�Ks�V��<�:�+b�H��Kuj�S�3Iꗊ���GA2��
�tq���KZ��͡����xhwV���PJ�q�vG,σյ/��ꃸ��k��+E��}Sw��f��쬻�鐹�&���4���ޜG���@��Q;t������)����5�b��L�{x��T�U�Fgo\嵜�uq/�m�.0s0��VT��f��%��w 7W"���y��y����7�����;����(v�ܳwv[;�����i�ũp�]\8!.���L��᧪^�֐ -��e�q��Q��b�'�Ir��PJ��G�rTKxNg�6�� �yjK�&i�zs�ʹv��i�+�<����)o^W��7j��Ս�'eD��|������QH��"��p�����7+yf��j��ē}�y�}E�V�5�0�ff^��½sR�l�����\��y6r�����x�-Y��v{��&�\�NΘ����1�:`�k��Ρ����WfV�X��/
ڽ;nr��ev^%4R��ԃy�W]U��7�gn��_>�к�*�g M�s��[�y����t�}@��=]����u�7�x�YC0�k��"����кN�V�7eCGR7!)�1��}I|7v����2p�u ��.*μ˸lk��YF�TTC��ol���Vޜ�?k��8S�f�ol�MFC׈[+ ~�V�zQ=j\H���FL����;w3knp�����
3�f�Z�
����6V�J���͢i�]��Qk̝����qML�q�9���r�ĵ+i��?��u��)P��<(D0s��E-+'U˳�3�W9`��y˥嗤9Ѵ�#������I�\����@���k�5���`�Q0ξ7s��6]���9Cj����r���L�(�sY�k
�jF�]�y�W��Cws#'_-%�u�;]��v�H�Y��jv�':EE�����,��H�,���sT��X��]K��l�q��N����85C�(�S��1����GJ�����ti���s�תؔy���h)ȭOV�ُ{]g�7���B\�gT�&�ݗ�;�=�Y��P�c�c���h�S���.�XN�^m�)�m�O���2ѐ��d`ô:��N��d��8O_d�姖����z���UՓ�};+��S7��\�y
�[6���˼鲌�Ǜwt���Wy](榦h�4[���)�rV�o:��1A�ʴYq4��&�@��X��7�%��/��RVٗzf%n���=y-�{ώR��B�˭�a�i���ۆ� �v�1��w3�����{ͮ�%�Z��х�c ��mt���0Y�nr靵4|+��+�� �t��@�Ӧ��_hʻ�P�Cbd�M&����S��e�6Ձ)u��LgoH���(�N���e��)�]�3q[s�,"�-�8�S�C��ݕ�sKgi>�k*}t�y�]��mvB�Kt� �C�<U����(�1�3�l�ڒ�[B�΢�� P;Y8���l��ǂ΁����t5�P��e��F��Wc��SFgc���l��R ��^q]��O�ѽ����w������g#�:��H�{Ni)��<r�Q;�gU���@������ԱsyKj��i����ǲ�aVlK)�.�g,��,�q�s�Q��Z�)Rc%���7Z%���*���)2=q��}��ź$c�s��c S������N��p�g���͜����ΰn�8fD�+��do-����\&��LT�*�8-6�qX�V��(��
�����㉴�t��m˼H���o!46�}[���0�so�gtډ�OPpG��7�It�Em�I�'pn6Cb
o	Z(%�:kjʏ��Y���i���N����q�-�ӌNL�{4i����s����v�����A��������XO^��M(��Эm��'���6jwn?��j\�]�}ٍ����$�]Z/��K�U���뷖�U��3���<mfY4�nՐl�{$;���pE��G� 8 �C°�xU�ASP�d	I��3����wS(BU�.�Jun��1�n�Ss�)95#L����;��ٻ�J���  ;����{����߷�?fgٿ�}/��k��Օ�� /�9�d�! �]v�!?��)���@ '�?�Ο8�F
�c9�~���4֝�]]���滒X��OU2�����e��c\m\�����Ƶ��k��V��hb���g.�����$��,��p[$�t:�A�iSb>����4��|���n��hIy���wug2X0 ���ݺ"!ٗCu��1�4\�+74����"��C�PuJ8�̚�0���`�b�]��eF J����j��� ���=F�J��[�k��.�,|��DY�ˬ��<
�b���x���v��C�[�ʛK�K��W1�R�n,��c���T�����Lt�3!:ɋ�G�%l������{W+����t�)d��2�j��@c��MZU��6) U�u��5jm��)eh}�a�m�˾�hY�/��X���B����m,�sT�2�#"�CRu�=F�]gv�U��
��Cmq,�y��D��wuҢ��f�h붉U3�v��!�.�3*7����n�2ͱ,���'W1��^��E��x�Vn�����O��2�l1�����z0�9�ӧ�U���7��7+m+��Yǭ���z-��:����pY���d�|t�R���i��n�q�������j�I�y���?f��=��D�%}e�t]�gVY�W����ٷ�3�Ч&�ו����y]ЩZ�̎���`dF^�4�e�,0tৗl��*^�5Xƪk��V/�N�"��<x�� ����&��"]!�HQx��.+�(�gRz
�r�4ڵl�-�7��j�7����d2a6U0�a�����{�����R�nZ�8Zʗ��nP���� �3}Y2V7(���ܖ��8j��ǋ�ӎ	Km��ݷѣj�$�����]9@ov��H^uJi\��ׄM2ku�	7�p�Nw �r�v(%#R��f�ۺvv�b���}���&`5�ÎU���tjm鬤�-�u�2�Wa�C�� �¡���6�͢r��\�u���P.2�Yv����*FX�Ɩ����8�+��o�Q;yDT��Hx�G
�j�r`$�2�Y��vx)ͫ&/^g#��n�u��j�6Z*�]e���y2�W
vr�Z/�eթ�������.s�L�V`ɛ�4CV �5|�ڷ(�y��w��Y;��W���DR��!�X��W̌�Ա��.�P5i�ux^W_ϫ	�����e;��#�Qj�JoW\�,e�.�Naδ�Γ/0�)o<�o��
:��$T�<��c��ZY,$�0�c��������.���.�}ڎ�P����Ҫ��X���"�����*U�l�r��5�ʂ\���GR��.Ԫ:�����2j�yD}�,�tӬ�d;Yū�~f��- �d�`��1�3�߯�}u�=$���ا.�����z�P���Y�%N��R�u���9�N��N�v�g��k�ɭ����V�;@T�보z k���Hnp{K#V�7'kl�ڜ��]�Y�3�YD��$�� ��.��kY6W)��1�d9���H�m�	���Xx���weB�I/�_G���JR�f���]�hS�tO2ɾZJ�t�(�5�n�ث<og`u1��C0TЎ:�a�vI.��y;�N4�B:퇴��+0f^u��grFs(�XPij���v7d\�8oE��/b���4.��G'[ku�:B�7�xPUf�=�[����Tk�(�k��M
��,-x�vaԻ����&�]Ƣ�Iu��h��z4�b���h�BY�]ݏ3,����"��ɆM2��2+�.��ꏷMq�em��=?�|�gL�ݍ[!d�*�N�^��i�Ӕ����.����[)��}��U�Z
]����-�Xn��Z�4h�H���k{s���o/,G�����g�xvsp�Q�mT��C}z�����3�7���zNKuȗ�\�gQ�Vj>3O>����	:r��g�L�#�4�`��e[�Ƒ1 o+�X���B�F]_n��*��)�q"Ȃ��p���җ�9ِ�D��`�h�J��VNv:;C�LO��z"�Ӛ,VV��vT,���4���y;����C���,ZWے���f�%C�ayZ@�&̕6�X�/��bL�6�d��Ue���K�˷����0	eG}cgq�G֏P��#��=6��Ut{FݧL�$|o%⮶�׊3(S��x�͹��K0��5�����(Y��Ւ��d�j]��0���3��p�$7��.[����l�`��&�KPLJ��Ve�Ŕ�;�gh�A�;ۈ�f�3X���9�W���9��&��՜t�6��֍S�Ԡ��*��P���e#��wj� ����6n<�A��WWW���Fk>�+�X���Ջ"W��䫺��[Vb��q��C)�%<b�Ꮀ����wr�ڌ޵f�K�զ��jIVp��c�n�Tb��V/	Ӻ+�O�@ �,"�|��0z���C�����Lz&KϷ��0               �+ҽ^=����-����7w�[,n���4�m��՚W)� �����uSr�w
�k�`a+�һ+y|[$�4���� c
:���*�u���0�ʙ�A�.M\q/�r|��ǋYx��\�֗u�S��L4cmq��D��!����ό�H�\n���՘�N�Oyt�sв�'�l���@�ۆJ������;V�J��n��H7I��ռa�>�K�Mz��v�qCV.�՘�rlq�r5� >���� EEʫ.�M�IlXZ[h5T)tUQwwm
�U�#M(����ZB�-R�hkE��]
�h���JF�E)�TJ`�B]�EE[���Z6�uV�UB�M�D��,��Y��7T,j�m"��Im4��)�"��,UZV�-��.���"Pū�^�-�5Ae�D�YU"�L�E��Q��u$�Ee2���RR���,j�Q�7Al-Y��4ȰY��W�3���ύ���՝جբJvn�[q�w�D�䤲O�C�|�����>�]������_����?z��+ZݩI�d"4�kkooa���}�Զ�#����[��T��W��T�5��Z�l�D@}����R��V��l����UFe��{��������:�ee&j��>]�;t$��X���(My�� �a�oX%��`���C}j���nW#E�[��~�����Y�~�ȫ C3���¶t:����-ʻ��.tj<1���ܕ�5�,֕�԰���!:3�vi=���'��P�u����7�E�+Y_'7ѓd��m���~���4F�������=q����yj�p�_K���ڷs{a�c�pQ:�R�fv�u�<,~���d\��0�F���:�V�r�,]�	m��}<����8U3Av`}�qn-�;z�:jҫ�}�w����e�vU�ȝ���c�ۜ��\ܗ�k�;2;]�aN00e�J�h�˹[#��>����z����ѷnoS-�{{�i���C�/}ؓ�����~��t\F늚S�u�+}=�����ߨL�\yA��+
�w��|��3��U�w���k�h���Pa���r��Wv����M�]���Doxi�b��O�F�+���}��J�q9��''m*y�7��+�5`���t���@�÷n�Ͻs�fknvs��k�:pi�mE�ۻA8$u��5�y�=�Vּ]D��ݯ�ܫi���U��e4`�]䢵�q4wof���ҷ�h�[�J4W���4�x�~w�ޠ\ќ���W?�9��[���sA���g�ѱ�T��'�Ϩ���1W�i�6�ޢ]��[�~��t��K��1���xu�͹ӽ�ׇ���˛�]yE6�v.ɳ*��r`��ˬQ�����F;J�WM�zophus�4ocT�%�	l]�;8�SX�C-�:O���}93�춃N����n�/��c�t����}����Ø��7][��G/��u5EwVM����T �5��z~�Z�/'��L���QIlY�Χ]3=f���!���{���
�Y��q�}����׭8�p�,�W��A�u�����C�I���^�0��2U�4}f������f[�4ԡ7�y#��x;����O��ϫsI���T���:Rz���������;�8v�ܤ��m�T���oz���2�_+XW��������kT�{�z�ݾ��1l�'^aJ�烰'@���M����k�c��
f����8���eZ�H	1ds�j�[��5mK��y�F/Y�+�t�爺�3�L��蝭^ˇP�7�s�)�W)tר��=�x̿��:T��j�+��{��ǃR�5i�[��0L��\7���'��W+�[3�zx���
�t�`��DA���7վq?������j�	��5��Ѫ��r��3�0&=�y�1�o+ݻ�u	ܦ.�ۚļ�L�V3�{��r$AXA[�^�c�(�^�=<��l�)��Y��Dв���k&Tx5D�/Ne�\S�+.&WǺ���d��G��5�^2�sƘuK�.��^ͫ���[���ú��ނ.�gU�!��,47�{��f�y�_����̙\��GE���5��:�;sbߓ�\�Lׇ��	A�\��j���.c���1��ڡ�J�F�[.Ǘ������uG�lY�q����������s��g6U�׽<�H�^�����ǽ�p8���=�ՠ���ڽش�}��XȲ{r���Xi��a����T�����5��ȖP� ����qgvQ;�jN�}#CɪBw�m��W�gnJ'�u��)F�Lf�`�{3K����E�vj%����ٓK�`�T{��q���.�d_>�A2$V瓾�ծ-^��y�3��u���؏��~��|=��Q��u�����^�a���U�焨�@�����53�TR��$H����n��WA�eGabs���`��CX��b�&s���#R=�ڨ����(�˓�ת9�)*E�&
өve{�-M@�dHw�/]�(���,���徒��{���V�L����T3JG<��zr�i5u��۞@����l2�&�@�C�^���3'vcy�*)�����n&|v'��j�s�lҲ���Й�A{��OЗS׸K3��j�$Q���u��f��t�}�@�G|%j���W����01�־}o��ϛ�y�n�~.�����-��x=6m	r�tRgm7!�ٙj�n�ΞЋfǣ��Y�d�H�t(^�y/s�.��R5�.>��:�a�tMiu�\W�]γ3i�b?���� ���J��%u�Z�,��]ی��sx����_9����	�ׄ�}�v���+�]vg��n����u�,���W6oK.��os�T�KI��e��I�J�v��%V�Ư����n
7�H'9�G-��	�Z�VF\ś�ƾ����o�qG�o��               L�^�}�W9ܶW�Ȏ��k1٥:
�Eq�7�����ĔQ/P�9�B4[AQ5����NmS���٘Vvq��b�wP��e��+��J�skl�w���SX��}��y���Bƚ�U�>�kq#h��O5���1s���7J�]r���r��4�ۙZ�]��twi�Vob�:dh_ƚց�����Q���\њ�ގ� 4�h��X7��S���G�a�9b��q��cd�X�NDܜ��珒���B�PF,�(U��utAeUR��?e�"�iD�����L��KA��жS(d�P�*��J�!M�U��Q��h�e"�R�2R��	h,T����Ť�P�JAhJJAB�)�����PPR��!WR�5TS(VS"��S)�$*�5AT�S%5UH�P-6�`�F*��K@+�Q�
���$U�UL
��aL
�
JEQ����E%�l-�0�T)�2�:'�|����W�~���&����顾uj��qON�C�����M|�.ᓽ֧�K�<F����_�V|~�#��:�W��`���3_�WG0�ߥ����a�q�էs8�����EE<c[vl.V���Q��q��W������پ�5�Q���~%z��q��o|�ީ�quX�U�>��/%?�]��妿��s0�K<jQ{�/�ȑ�w,��s7V�zѡc��>���ۓ�����ט�̐:�P.�G[p�������9�߫�@2��:P�@�_Ǥop���~_K�q~_��S�gUj�C���|��2���g�5������\�O*���-]���/}~O�������X���k��]O��MH�ˠHK�Q������\��~>����5���+{oӘ��i��o�a���_UW�_���Ӡ�"���ߠ�CYc�Q{��bQ�p����\w�7����n��>$M�����@��}i��G�c�sa�+�U_W������_�O����:���,k�w���j���*����T���N����h�u��M"�8��B�M�RZη�{6r$����5�(}�*S�b"����bq[c5�kp��c�Fm�ͼ��������y��f`Խ}Pֈ���^3�וֳ#a�/}u����Y%6k��'1�T;������������.�q*����Y�u���j�{q9:�d;����t�)�� �w��ña��[Cw�W�*�2�}6s���O	l~�my����$��߶d$����'RC(N�B�C��ߨ�ڧ�!y�g�{?5�I;�	�<Ʉ�{P�	<��	ԁ��|��{G���~o�i�a){U��@<ɖ�d��e�i!�!�d�n����ܐ��|�u (^�He8�u����%�):�N2Cl�@2����?=��c�y����C,:�99P0�Bc4@�n����|`u����!��ϝw׻�!��)$>&ٴ��CHKI-�y�M0';P:�m �'�w����J���~+l
VNc���5';ھ�S��D�ܥpk8�ĻͶ�n��k{򐅰��>$0���/�&P�)hq[0�Cs��o�׳�-��a �I:��I��)Jd�!��&7A:�^h&�u��k�{�>sćn����,�I>0� M�e �C)Ē|N m�ZH�Fu�o�9Н`)�Q�4�4�:��!|�!�L�L2ACL�	>$&P�wwX����$6��M��6��*|d2B�RCI!�T&X�c���~�!��C�Wh���2yRd�Ha�T��L��^*H���=�����za���I�He'���8�>Pq�l�Ԑ��T0����p�ӌ�d�yD:��M��l�q/�4�0�@Ϩ���a9�b��o�߾zHZM��	��'�	0�Y2�q�HCi�� ��!��4�^����e$0�a8���@���RC�$�(	�@0�q�i!�~�>o��͹q>ƩpuE/�lg+g3��*���G��~���{��`����$ř�<H�=��V�<o����{�=��I�
��|d�$�)}T�g�� �J�I
I�GZ��㚑d����-�/�̆�8�=�B�S�C��I/�Ԗ�Bk�HR���&Y
���l�!��@�������C�03�gW��θ�5@|I���&Re��C8�L!�!ڗ����t�!h[�'���:�d�XJI'RĆKaIl��3���>k�!�@�>f��=P:�q�l�d`O2	����>c?3�s���8�e	���^��/4y�/դ���I
I)!3��X�~�t!�q$)������<��!�����!�L�d��ŭw��l`N��y$)�āԚa�'���Y�BM���Jd��^~o=��h'R�-$��� |Ja�������Hm�l>$��3��*�&?;D�?*A�ą;�O�k��>��W�f>Dን.Zчh�w732d�^U����p�$�a
޻�{��0�|d�!���I��Ra��0(a%v��ꃉ��:�W|o}�}ޞ����@��\�����mB�_{�ϼ����+��۠ex�>���K���sY��A�v|=�ӗw���}}���E���#flQ�:���-���߱�2yb�<����9�Ƕ��}罛1�2�B&֯7-��է�ڢ]컾̲�RIXp[YZ}�k��s\ꙙ*t^���ArR��g�C�Ӆ!O������g��X�كO����򺯪���GoI����.F�3�s[Z��/.Kյ5� �Ԛ��%�*�w�>;;�վ���L�9�j]?^b�{�ļ����i��ynTd�u������k��	������Mm�v1.Rj><^��y��ئ�CB�b������Ro{�~~��c���x����5��p��[`����D��Z��eĹ����@su��HL5:U�sk����?���W�__}_�W�ϟH.+O�\����X9�����vQ�ȯЪeq��nߔW�Y���5�f����k�ɏ6�q�T��<�7��UT�����⶞�Y�[Q.�.��|W5�J�x��	��{/�A)hVoW�.κe�!h���j�B���.�!H��<�=v��5���G���v8u2�q��s)��9O���I�I�>?�Ob��"xJ9�ZzL#6}ݾֹ�w5�f��v��B��E�� ��(�)E�Ȣ�U����V��w���:�����4�X<����:ws+VP�]���W���s��杚��5@	[�~��z��Q���+uu>Ƥ��5��[{��'֏1[F���V*�o�����Ǹ�t��.�+�鮇��p��}�G{b8����wn�����^ĺ�J�	��xޣ�G����_��i����oj@䟁����n�����*LVv&�/Wo2�[C᚟\��E����)�=cu��>�`�����j�\v]�A��=�̰)�T�,^ҵ�H�o��=ή�"��lEP��녈o���%!�7O��r�R�y����s����+�Ggh���^��[ ��]:ti3C���XT}��f��3x]�O3�/{,h1͉���\d����R:R��Q��GE����g;��1���q���hZN�a��yL,�J�G�i����              fh�/���;�eW�:a?Z��6�P�\��wW�+��;P��[����H�3w����*�eu���@��^ʸ6�W�nhx��/y�
��"�;�U3`� +���ܪ݌Y����Yܹ���wl��ڔ:��}/Ri�_5��I|���^�&�%:M��Y@��9G�m5<S�?��^�e�[�M;R��uX�l4���c��ܣtl�u��"��u�7|���R<9yNC+yF�MI7��\�O}?q>C�<���i�j�!�-	i#"�IJ�	I)�) �%"�,<�.�*��U$Y �P
B�	:���D�����Q`�P���D�X��L%0�e0T��SI���LQU��R�"�U�H��b��U}_W�����?�nzr�к��	34�5�ײik��[���UW�}���L��b�&���+������0!Bu�Q��|1���ْ��o�p�w��7����QѼ0�)��|���OоFo��*G^l����p��V��r�wZ�U�m阡{�9�j6p�׺�^�؛ɹ�/uq�+1�w�߶b�[ķ���|�^'$ڵ��+j7�}p]��~��&�E�^k>���ygL����s���M��.��{8���-i��������UP>�'��u櫶�N.��*�����R�u�L��x
��C�v��c�;�v�Nl.�����Í�7ީ"���=�� +�X�:ѵ��y͡��p���x��]��s��>]f���xa1����ĖaO��r�2b�(��b�|h:�"����||��D��]E楤��xk������@�Oɷ����J��݈vM��k��G7������!���������h��^V���#�����4�&�"��ZpV��9�#��~5ٳ�T0-5�D����yױ��t*ݖ_��|y-���J���[{��/�޳�{�.�7AK�O{}}zQ�u:���'k[<���W��t2�]՛��Ow�����ʌ����^�\�iw���znS���/����r	���$���R�m3���Ӛr����꯾W�ϼzn����lXitە<%d�����Z�3��T�Nf�v� ����s�£�G��^/2gzktp"�qlg�}��w�����W�I����3���.S�W^<���ҹ���j�5��d,䙋�s��ȓ�{�)pv�s���������w��\����+�31]F��m+��#��i����}�����jԄn�䰫���}��Y�}��ψ!_���t�ͅ�鷣�[�]�빨�k[FN�˧&O�a�ύ���ν��o#]�G���{�٥���we:بxi�y1Kb���;g�ly�w�EpQ���k���K���үO\��K�ٿy���3��kw^���X���װ���y;D� ����ܨQ��T����E�mv9:؂���� "�Dä�m�z�1N��{��ʲ-jt�t�Z�4���W�_U�^�o㞰(���F�~�렻�8���ꄀ�A八��I�7����7���{���Y�٪*�T�LF�}�X��~W�Z��r�U��9�4�i�I5�^4��}O�iڏN�>T;���=1V�֦g��a�41l��4�zjnq�NN~'�.�B��x(�>%�*pU�U	��FCS˻���p���;�Hg\c���ɘ����j��	����ꯨB}����o?`5���U��-�٫�O8�N[.�Ϻ�A5�zϹ���ߗ�m�5߽���FMy,ozwK�gaѨ�JĂU���^�������Ԯq���4f�9�w����G8��@�Yn[�Ɲ��ƂV�˞��K��O�V+R����'mUC3b�l��_VU����:��c�,R��;=G�R4r�i�k�T��{֛Z�掩Oz7vI�I��W�W�ܣ_�­g�8�l|.�'y$��Mh��<~����5����>.�'�*�~�������T�ZNu�ȳ���W'k��	�_e�!=@��w^`/_�����Ks��okɬ�S��]�f�2���y����묬F�����wnz%�����*׷�4�\���4�y3�=�2�X�t8�rL�E4R����
=� �����ҵ��b�{J�ZR�[tVN�������/t;��~�+���)O�׳^P!v�����N���o�Nی��a>m<�~�Λ���8�ܫxy��aڙ�~���˼㫘�Ee�>!md�}���mȟ�t�������1χ�m�oUT%1#�o�2���9V�z\��zVv�O5o�yn�_�P�B;7����c7�3��+ω	˰���q@`�v���$�S�<��ُ[��{�q��bU�q��}_}Uof�'������䴪B�~!xfye{0�e��;�NR5�bDOZ9��r���c{�q�ܢ[?La��)p�@���Dv���϶u��΀�(Vy��xv��粍?N�=	���y�Ԏ����]�-�W	��s�XC�kϬ�t�Yv�ެq�-�����ﲴ���̫֘�0u$���J��)2����GQ�=.�\uՍ�>B+b��T�7s\���(u�B���y����s��$�g틌����nЫ[p4�V�X-��|��(.1F�yB���W��%c�,��V��=ї�E`eS
)�[��y)�a`Uj�t�2uh=v����&��)Zn������&��~�/U��}W�x��ؐ!����>�oo/�Ƿ�p,��#�V'f��&�b�t�[����Q�y����4Ӽ�W���#���               "jOz��⌫ab�K�
SU�ވ+[�q�5{`�S�o�՞T(ؖ&��X�.������{f#�Z���;�ϰ���W��}�m�w�Hp���E�Ur��z�Y��fr�O^V�YȮn�n�rIq�tG9�7��ĝN��y��+�2�F>B��)tx�������p���Wΐ�cF�`K�u1�w�91-]�V�C�EGPSo_o��%��ٳ�PF�Ц���f�gEI*Af�@��Ӏ�8 5�����113��f��ł�PX,��cT
���UB�RR��+�b�M0� }RP�b���H(,PR,Qd�% 
#@YXS
AP�$D (4Ф�
�Ȉ
Z�QA@XU��ϟ+u��ڼ���}����x��mq{ْ�8���}_UPŝ��+��m����'ʳ����4��\yըh:y���ʾ�ȼ�e5����c�z��*�j��.E�{�[���S�-ro��D�4�cl����\	�
�a�z�+{�~��puϼj6���v���!�_J,xb��ǹE�O��{%�����7��	�	�J�E���f�Τ�Z���:,�c+uΝuy���/�d~���3�s����LT���je����nR�����9Qb����kWO�0��f��}�.Qxf��X�69�A����P������S}�����c�t�m�e{�K��e�x7J1_���h����L]�������U묧k���Sg|�#F�=���QC�ǒ�b�7�{^���d��bR�]������������pB%d�8�8��iIP�+nK�ꯨm������Q��ۏ6<̫�Q�e^oM>�^�H���o���칿+�ӫ&}{��]G,L�]}J�;��Qx֟&��]�W�sS#QVp��O{>�'�s)��6�w�N_te�����!�fO*�J�V���,��6��[�({v��8�/��;�z�Q�ħ�����t]����D�R���Wv�J��o�����%6��1I�U��R�^�����۲����h����n�G}�+�>��5��=Z�<g���������1*���Zl���En��ʵ�(òoزv)�c;���YZ�a~���[�G۬���y�2��cJo7Ms��o��ӭC)�m$���w���ؒp��pC��0TA&�t]��Ͱ/a�s�hS&)�!ry��\Td�˅�͏���å����ًF�N��ҳ%k��w�g�׽����N38��2�)_�ڝy�߹~��(t��iߨ�8&�*g�t�^1z�1�p�;�pM��&Ղ�zj���ȴ�M���p�h��ʭ�wr�W,��H����ה�L�s�#[Ap� �	�x�`t�P�2h�V{+�![�F�m]5
G��*67>�������b�����b�"�)�����WQ3�l�*��>j�H��wS]�>v�)���S9��;�94�*��sM0��xQt��*�ᆅ��M��ã�mےNJ�%�m� ])��0�gWnĮ�lH���<�fVk�����fˋ���}���8�����5	��*��Ӻ���W\��t�����O������L�X̪�ٕK2�ϴyal�|�[f��i���O�}��sfd�i��Y��|�M%���u�6�T{g5[��3��'�=i6�2n�r&�kQ���w�>��{:���P�T0|���D
�z�[ܫYb���tQ�#5���t���M:������7�r���&��=On�~�)����^Ϯ����L'�YAJ��+>+�Rإ\{3@�}=�"�Xe���K�U��^��m��w����6>AtW�b@����;"�G�u:���1���9���9t2��}_��߷�7��5�_�ƨ圸i,N�N`�_=��b�=�-�h���{GDj�}q]��JWw����������j�핺/��:���e�1�_>m66���Z+�Uo�[uw7(\�W��C%�YI���;����^���Y���-���6)�\.��Ej����J6~�5�]mʳ	i�c�=��wy�w���Y��g��@x@�I,p���ʱ�5�n�t�u�exVYB���	���s!�{| ��Ѣ)<i2�xS�Uv��1{8���%��a۵��7yvlE�!��=ܑ=쬹]*��M��[���s1x�����!��>Q���Te�T�n��ӟ�fr����w�<��y�=�M8fNU��*���/5X�����oS�m��
r�N�9����z���3�j��(���S5�r��fG\�C���[��VY�Q�:N<N��{<�s��m0�5��^��Vqb������Lh��J���v�+�n�x(-=z���r� ��3��+���0��+�+��%��⍡��n��bc׬K�����p���=H�E��ia�|k�h�h��T��X_��I�tu��8ګ�p�虬�}H�^���GT|�^���;5nm���覆���+W��!c��m�o�,۴���o��;�d�9��z|�h��&|)ap�$��N�U6��K)���+n�x{�m���y}}�;�0�(�q��n�ܦ�My�yja"�?i�O�V�g�f�HTք;�%^z�{:�2���WF�L�����㣅*�A�{*���E��IRмױ�{�Ϋ�癦�&޹5��CF{��8�]�Ng���{��)��S3n��W��W[l9ީѺb�`:�ОJ�^ݧ��f���>�͵�0�L,c�VJ��9|��zhmk��֢z"�qr�{�R󮝢u���&�;����	���4��<���B)��AV>������*8H�5L4xW��]4P���ޘW�&�<����[Q���]��X��ڧ���YV\6P���-̥�@@��չ��y�K����#�}{�:�f��~�SF{vezz�m'��Y�۬aל���%����3I��@}4�
�!�Y� ����[���cᆗ���B����	��H;��hW1��mJ;�m�z���Ǐ�8�ny�szK�`JM�ݛf�W��;f���U�7sK�U�x6j�ïe�87��//.�7H^�<_s�}0f���+(?��;����s|��-�=��ؾte���Y�;b��J�_^X/�vwqM�X�e�L�R�� ���tbgU�v1�s��f�K��*�Cu�7z�A���֣j���S��q��|~2�VHCA�{�'fEOO_e�o5�ѐ�n�gq�����"�p�{�$�=�*í�C[�[Z�����������m�-�6��Ps�vnȳܭH��F�W��X�2�`�����k�̀   wwww        Q5$/l-���w�v'On�Ϝ�JG�ء�ʐ݂7�n��*�K����<���
�����+�����3�s\E�¯x�y�M�b}X�E�9����^�a�X�=�^��u��A�$�>�|{ώ��db��+��YZp�l�^�8��f�l�|�����YO�kJW�V��{���eL*�)ٺy M�����z������1;�����"兄��;ȒT�D��y7��NP��nK�8�s��;��ϰd�#H��b0�HS
i��PPP ��[
��dAdX���0R5P�

R:� P�S!�) U�%$�,j�*�"��%*F(���R��U�?C�wNy4�g���b��7�N��8���.<ֻ�� ��=>���_�7�^'�_9e�f�ލB�����8��^��|+p�?po;�C�j
YTtQM�+0mi�=�����l�O�^m;\����C>��}�k����z~�@V~�i��-<>��w���
�j
�y��w��:��B�v~L�D�C�~�.B~��(Uo&�zxp��f��4U����w�2�ӡ�i�f ms��7�z�uG�y�Ӂ�˿Q���}��#�#������C\8P�b�R���a+9�2�ԫsf+��?�N�R�k��t&�W�5�����\0��mm���%%���}_/[�������.���o3�_��{�\1����F0}疁x1Q������O�h�v��ޟU�1�(�s�̘��v���y�w0����]��N�9��֝�Ė��g�4Y�H��!�� �����\Sˋ��I��/�r���]�,�j�;��:��|�w�qk{5�o���s�6��t�����x3��]^p��:�\�ԦktX��9�v����q骴Q�;�.��\GY�]c���Y�G���Iiƹvq��,�s�aںx��:�9�+a���a��J[V�\��rv�K@R��
.��2�=�IÝ��s���$�7�kAv�~G/��z����M�7Loj����4AF���P�oɍ�Ԭ��v�:L'3]�C���w��K��ˬTZ}�)<WW{80��4i
Љ�����x�זz���T4k��>ۦ-����k>�=�:m�2���:�m�S�	�Q�U�ݷ�k��xvUz�:�S����ꥺF���^o��\�Q�|>����t.��u:^Z��P�M����K�2Q��۶�9�N�����\z������r�&+b���V:;��nv��zm�d>ڙ,�����U�+'ti���.�,�'vǹ��;� ��l��.s
q��#�c~��5�i�w���m&ǎ�j�}K@{"8�.*���X���47��� ���톓0 �Т>�5��ѣ59�3�/yǽZ�,�m�h)��g���;uri����'渨�Ș1z<��쪖.�xb���^?o��镢eeR���2��_޳T�����7�=(<W��pg��b�����r�{�����1¬o����iCWj�W[��U,��Ç�U�V��1��p�ru���wޝ��i.��^�u����P ��u�{��Y�n¯vN�୮��F��ov��/iTr�I�n���]�U�����?W�	~�O*�շ�SZ5����q2���-���9�կ���_���[Q�V��*��@�����ˮ�9���xW|���0�}��3���G���(�ר�jl�q���o@��yx��k�fS��y�(�ѵ�r�|���>x�t�h�q�C��5�w+$�V87�s��������Tm6�2%9l�q#�
�.f���=u��[�q��U/����w����U�m��T��{u2��.
�xg��rW3b���g��f�l5���7/��z�¯��痛��ô�dx��[z�{;u�z���
�Y��ՓnS[��\�$����u��_p�'�ٔ�L۪O�����g\?��ӷ~�ǯΙ���y�l{��q��1�V.������j�M<(
�٥�� �?C�&�3Fg��`�4x�>�P���Q/u����y�(z����"�^Z����T�U�tݺ]�E5�x`���B��*�A��]׼��)P��S=l]e
��.�6�0�ܱ)����F���t��W󂳍g;��m8�E�zP���xxk�,���2����z�5Sv��NY�3~�Y�5Y�kz�~�x@sd"@Qێ��c^o��zsǯzp�
�Kx��]��B�&$���?��:��W�� ;ۭ0�x/��`�-(p�[/�K�FѮ7���Ơ@r�>�F�(��K�$?+���~4�l4�\�@�]��A�+�a^���*^��w�9@&}�]�?	�&	��鉗;�{�ʘ���:�ڏ{%�	�לM�M0�+hQ�u9U��Lֵ�{>\ד)��=F;Ee��qYn&��1�{���<���u����=7��-;M��48��nsTy����N�8/�"�zi�5�q�A�&���5�cE+(^�����'מ��V��\�uJ~����l�V�����ڈ�f��jJӣ�I�[��0~��4�Ƌ=ƿE>C	�W�DSF���������	L���¸@�Tdg�7��r�:�Oְ�!I�3�SnN[�q���s�ͫ�j�3oS��"�G�B��6��X���4�|��*#A�c�+U/� �qv�e��Up�1�a��43քZ�s������垿[�u��줴#�V}�);�=����k��r��X��:������jx�7�<�;�]xP�{eT��yX��w�>�+�t=5����5[�B��L��zZ��ܖ̳z���^i[D��^Un@>�,5����йP��;�1rg�ۄr��\{Ϋ�UUp)�(������B��ߌ�1���5��M�3��Ո<�>Ks�qF�r��tg�[���)�H1��,��4B��F3�i�Gm��t�_צ�<4G�\e��j�ųp}�|En���M���'�N��Z#�=|4V�k�V|)
B����Un�"���^���v��x�m۷i��]g��&�&s]�������枦�[�u�V��oY�W���>���#LFk}wD���{�,��xxx441h����\>|����}�&j���|�k���ǮM���ċ]�tǰ���їxn�\k�?N�ʳ�xm�'�~��>DIo<�L��>�U.��F��X(���t��Q�l�J�ENk�Ò'���w����S������f��9�|3�O+F��]H���{�tU�W�ǳn��V:�`�/C�%=F߽�S��4����p�U�v��V��b�e�Ѻ6��,L��e: R��������׃��}�Uai�@V�3J� ;���{�}�4�]|0��]ǅ�>�*�x�7Z�J������ET��m�����g�_U��u{�!���(ǃ}[�^������u�C��ox�`˃�H��*G�vWiP������X͸е��^�� ffT���H޵���}Ĳ����Du�e�\�A�<tA�bq˿C�+��9՟[y{7�2���&��M	ۃ����մ�*4�����&�v�u�CA��b��z̩�oSv7{�<�˧�έ�x��BU����>�|V���}-����"�u�Ǧ�����o��մ��݈Y���� 9�d^=�ϑټ��c5�VV�76��a��C�v�
�w"��b+���>�H>�#}�};͍�               "�&(�Z�cӷ;��ˣ�O%���v��F� H
�FQ3]��e,V4�K�����\S���s�}i���f��X���6T�I+2��uڬ6��\� C�4���SceEeлJ�Y��%q�f�.
�>Q��;Pl��l���X�Wi���=݉ �t�Y ��r�;{��q[4�]J���KibX�4��˧��ܜ�7��$ڛ�K��.�ʾ�
�r2���c,�(宴�'��$N)�~hk�D��QQ�PUb�"������,Y
�
���QQU_QQ�R���PV,F(UP*+#UCDAj�(S�S)#iR��QEY���E����EU1e�CItS�Mݒ�Z���y۹���
+{Cr<��Z���|�{o�f��o]z��W���U�1�<������ѷ�Z�L��`Wu�4�M^����<��`"3^�<j
A�h��G�H���E^j�!����y��gT�.�n��}�����o�N��Y����;mf�[mδޯ��9��6�N��6�h[�t�.��<��q^�n�C��X9G���r�Y���{�����G��CA�MϘ"�{ty�x���wzs���)�Sc$�UD���0��m�u�vU���bg��lXc��uG�����k�3��4�OooC���o��7�JAj��o�̮�Z���8�Os;��:�qG	��RK}�%�C@�Y|+���*�!�a�@6��S��}�U�g]g��
���홢�,.�ѽL'����oe+ˢ�S:�˗�Q�L��F���U��g�4xx|�����P��h�B7�{��[3G;Z��<�W	��st���V�}�Q���LUܾ���Z�m��R�rv��0^�F��b����"��Y�
>K.�YZ<0���me�L}�/�TY��A�V���k��zsd4�j+*q���>��q�Y���6���7�wYr�Y�㖷�.r��yb����׽Ӹt����߶���nG���-�m�z��6�S̖Ι����U���r�¦��?Q���|���"�"�Ƶ��[�銱b{к��녢�pB�E%9O���~xu�9�����nͼ&.9�=VQ1?"��t����*jc]l����ʯ_n;��w]V��.h\�?���=���`��3V�ɴ�_+�٦?WC�Fik�7�zڮ��`�i�맱8��ۢ����WY�{�yoV
���
���`�����F�T.�i�I����*��;�n���g��~�������Uō]���X�#]�z�*��� ]�0���^��2���k�Ij�F�oVu��}�&�;?��<̿.V+����X���b���Z^��5F���Y�����8���Ǐ�X�5�c�����9����=�1;Sg��}V�*��y��ösT�e��T�k:��u�(�÷�u0��K�, �X��6�K5�xn�yy�8"N
�Z<�ECEP>竧Z�R��զ�����H����Q0��Y�em��:&:蜚�Á������6~{�R���]pC�W (]-�P�nP��(L���b���M�I�@��h�Uo�٨r����;�5]t�i0�|�;\�6c��)�yH+�S��w�΄#�5�����ws � �᝕�r#�ǁ$�tޏ���;p�t��=:K#��o������:(CDf��w�z2@��������wN���˰#c�q%�)fR�(P�g�t��m��j�#���yv������O,P��(`�Y�B?{W�Up�y��y���6���6v���Jv�Nz����ox�v���땢�ʉ�RyӦ����OG*���lxS��j
A�c��?d�دO�� *W/J�1��m5Sv�SNW��3�k�ɗ����+�T\���N�"c���n���}1a�4m�Cz����@"���Y�t{�^��-����Bk���-M��n��ABTN[w��t���2�6�r��y����l��_wztӓc�m3��Y����k�汗)��'Zg[�[�9SZ�����7�{~M���ݦ����'/��|K�f���E.��e�A�U�7�����Ջ���KJ
ٕ�7r��]+�>6�}J�����]Ĳ��xT�3�u�}�ޝ��7�&��Ep�5���\(`Af�������wH[4Be>@
�
q�����=��S�y��;�*�>@��4rk��=</e�!�[��ehѶ*�Կ_�����^���u�w�<�z̫Y]5K%��K�7����3�����r�fe���;�nk���ι�k��u���+]�|�]�n�>� ~�v�x:;��@�������®�`��������o�մ���>a!C޶+�U�̭׾�F�C�U��Z3�t����3C�o}�ԧ7Ѭ=O4r�l��n]%2�Fs��(�n��y�k]e�r�7�Y��ܠ�N�kئ�2"��E��l�vS�WSr�0�u���������o͊���"��(c(U���6�0�ι1�����pg��پsW��5���YM��X1<��K���	>ŕw��{,�\����W��*�{��d(�؛�U���9H��s(M
���Ó�y�5����y���|x���N�m:��L=��\*]dϝ�x���^��<���0{�e�+ο��륹,̥��㢘����w���h�x�CG�|��kHT��q�$@��/M1F�=f�4��]oU�oo[v͉�g��)=���l�q�sz�s��xͫ�u;���5�
�����5d��8�j
A�cC��MO=��Ou�Z�'�ƴS�t�d
B���T��x�Ƙ<)YCw��	CY���(�6'� �x�v8_0����mb�.���ܫ�Һ|�5���G"p+�'\�O��:�M}�t`"ŏx��@v~�I3���_!ZK!��5[��X�Ƒ�r���ޏ����O�VC��wbzs9�����>���4h�}�X�|l�@lp�{;�\r���y�:�&^��
��ϰx�q\���9�8�VoN5F�"�H�i�׮��i�#��m��j��::R�^޵:�x}�VX��FP��h��O�Z���Tb�B�*ǅ+�¢j�z��o��;�Y�)ߦ|��_��:.���S�c�9ْ�-�pP��Wv�hЍ^i���&`�z�x]G/)Z#�N�����wx�I�JG�qLѣ�4w��}�؂�0T�B�@�ߊ�է�wr��>P�����:�c�D
�C�����h��p�9W[���]x��G85�z��or���-�Q�6�(�:�u��}��ǳ��5��y�{�r�3.Y�V���cՇi��oX�=��.��O��E�lr�n�S?v�YJ����*ـP�J�
�)T%�*u���x]I�J��ok��vX��q�,\���[��}��S���q��e5�2��u4�v��}}�s�ϯH���
��0{MO9;��a�J� �f���ܽ����l�r��7�
R�'B[0�ԛ��F��y�t/���aK��R�����[��:�2��������{�kH��^shڗ���l�SCG9�P�S��S)g[�܋�`�v�2�V�/��\��3��Gn�T{9�q�n�-�B�ڄ��LC��
�hX�lT��e�V�t˫��в���FS��u���L��gX�Cy�;DT+��m!�܀��o/$�so�t��]����^�U��1����z>�6���з��=����ʃ�,�K�                ����w#n}7�gh��T狎�N�2kn(�,��ܻT�`��T��n�Z��� ��9e怺�e�\�c"��F���0����2Λ��0�Z�����w�C�O����!���E��F܇C+���w��e
�7��<�QX�=<����w�M+���}�jy�c�q�3V���}�>��\����HWf뵊�&�&�DZhb�5L��d|DFj*A*u�J8KN9"M���{�Je%%C�R��L��WCu����u��RT�����Q�H�H,�cE,QQ��--M �ե"QE*�E����#EJe"�[K���V (Q�rD��W:�N���gt�+����������u�H"~�+����8p��Q�>��"���\?����<>@
��P�+��$�S�Ó����5��q6�Ue<��.yx�uCH��j�4�b��G�H�����]�!]U�̬z*9Dg��]P�X�g;�t��.q�t����T��< �J؈�;s��Ѣ�،��e��_M&[}�w�5ntQ�OXgu��y�P���Wo����xU���~���|���b��fs��sz�}�z�3�����c����.��j�/��2�-L.�1ݺK=KtI��ӛF���y'f^=w�fB�s�S�
��ci;��+�'�n�}]�^�[�D�����ɲ;F�u�d�|<�����9��s$21��?�+�P~���2ǵO��!u0�u����=J�dT��t��բ���%��y#�����d.�L��^�z{���q�!�MN�{���{;�N�9�U������o,lo�U�Q���{ވ�eG�I ��������_U�;�*�����җ��'Y'8���%��bʃgs"WY��M����]*�W|z��I��<��*y=����>��_�)�w�{"�B�ѥ��4�>p�4q�N^/vћ����w�JɝLoS/����NKԽ��VV��̥�.�I�[��ɘysk��EG>��-�ռ8{:�၏E�5��=�X�t*�B� |��Zkn�wq����\�l���%w]����Q�k��K�������Q�p�]\�Xĺ$:�J\��ۍ�ؔF�����������Xg�=ੂ�ׄ�N��Y1[3lk/�׹�¿�"jom�~1�X��m��}�g�����3_M��Zޘ�2a����T��[�U�uyW�y�:頁�,c�<94Gn{]:�Y��xQ�}��Z��^��i=z�6��;<��(wg�s�N�1�}Yw��b�^\���p(wsj�wØk�X���nCr�Q�Q�H2V�5�xg�7y��k���Y��kF�I��ǠQ�=���4o'{-P����5'ݩ��v�����֏zܝ9w��퉡�a�C�Gv��uQ����<�j�.^*;%�˄�w����.\��Y�*j�;5�]Г���#&;t���t�X��ے�B=@.�"�ۭ���3a�x��*�{\�z$�gun��=Fz_j�L��8&�ʡU��RR��[+/��<[�i�\��A)-��7EC8�S�7#�n�wH�(�:r�j����.4��	�k®�l}JRkp*�e=V���7��ka���[O/�H߻�A�{�1�T�����D���z�_d>�3˫<���W�Ź]�����m��v	�k=�T�V�����Z��A:�˧J��{c�1*U�e���z��5'��u	J��%��8�}���!l�3W*h%�^��Ň����ݰM�_U����X�]�m#���d��[H��.�K����3<��u���U�*j�������䴥W�
u��������mߦ��Fy�f	d�Z��;��*�=����@�_�������^��65o��)ZӁ�����;t��{p��mr��xM��Ky���;/96��v��w��d�8ܼ��dzr�&�u]e	�[t;9۲�]3V)�/"]P��;<�m�֦Ig�dQ�Ϻxl���
�F�_��pzz�̗�$Uպl�d-���wў�ʌ7�S
5��\���Lw����0��o:6jS�{`lm �ï-s|��v�ͺ�!5�!^[��8�:>/��4ҧ��C�q����̲����X�WZ�J�W����|��݋���{�r�s�P���|
Xpv �4N�����`⫛����4{鹉�n��T;>�Ϣ֒�����g�����u�j���+=�J>�|��Y��k��fe�~jj��SCs]�"�3����c�Y��� �w�J��#��V��Z��Y-b��/�5�B�'�q9鱤6+x���Q8{TW���;�j����ԮtcH|w���5��`�o�z��g��cy�fm��b]|��y<e�M���UP�^{��Z5ܦguȘ6�yZ]G&t�O��Z�ҷtVN��o�ߚ^*������x��N��D����T�J70o��W�G=�ޝղ���I��M�f�8��e�}޹�޹C7ݓ��uC.�������v��[�۾���g��*�O�*�k*o{�oogA��:�Bl��]�~��E�;�T��}5m����^W���T|��~.�|�Y��?�k:��b�
�'!%����onv$��.;y�6��k��ʔ��ˈ��#�Zi<9o]�`��H۸B��g�Q��S�ǅ���xՔ9�by���[\�Һ�I�w%\�L�2�>�"����>f�f����#@����{u���N�<jĎ�:F]D�g�+$W�s�}z�S����v^��\Y�XI�H�wgJe����vp��r6��kS�&�ݏ;����]u���o���y��A6��*�!#rZ�⪴u�.�~�Z                EEE��"m����Bi�]zv�Y�B\pmp;Y�ԉr�\/���n��er�T�U�=����u�TZ(��5�Օ��ݘ�*�hw%��[س��k��C�A�6�n�Ӿ4֑���╍?"�켆Ni�d{us{��Qv�s�M��m�MpEQN��w��wI��5_m���Lg7O"�OGgy��E����r�0��o7�����Ť7��m^"(ɔ6>Ň]��{�w_S|n% /\�D�NI����� |IJ�m��E������IUPF��1�u��t�5T
J���CU�UB*�)���ŊE�)�Ī�j���� ����H�QB�Zb���H���0ϫ������O.�\T�49��;�x�Z�va������-%92��-�A��+���P��=I�i�T�o�q��I#�r�`QNb��o.z]z����$�ݷ5���(�F�"�k��Y�(�K�%��Z鋊�ZU?/P]t�{܋��o�l��j�^?���r����ݵ�/E�&�dT3}�r�\Oh�֌�_q\`$�Z�O�^v��#�J�g�1�ݣ���ʹx�#'�nq�x�ʶ��Y���iyկ�0�R�A�;�m���?��4F� �k���U��ؚ�`�x{^�i5w��s���k��%l��}��x����DI�6�Xz�5���Ǌ�-%UWa0&�=�o�<���>��,I�l9P'��yX�gF^�����I7��x�n� ���)���e�����z+��:M	�F6ߟ��ǭ��[x��W4v�}~��f�$l�N����f�on�"��\ș�k��Tϸo���^�xm��ŖOY2�m�S���x��"h�V��훦�i��P�N��H��:��#��\�3�SI��x�Y�Xd'�y�]v�PNO���뫋����y�k���.����Q/v2��&����uj�og2r�Ͷ�JgGz�^9�����f�k;-���x�]��0�]��pC�x�n��A��۷]}�S�s�5��Gb�/3��,V����(W:
q�^�ʦn�^�MR��G�����a�w�Y~��õ�⤬���{�H��da�:˿䤟�u{�v+c�r#Ap?�y�G���=�sJ�r&ך{��0{�}�=��to
s!g���>�žǽ�y�^�?U:+_\��>i{�bygW9Ee�r�X8�~��e�YVq��	�]ֺ�v��@��ewV�rKջ[M��f��u)!ý<���^��z?vT��Kp�WI��3[���Kog���[+K��>��|�o���%��G���sy���m���g��]�O�i>���Wh�f|R��stl�觸oe\s���ힶq��t��Gz����]���Q1���6�a��"��ax&���%�u��L߄���џ ��+O�^�h���vt=d��W�ُ��}��K't]9f����e^�����*���6p���,k��j������d}ݑq٪/c#�yێ�k]To{c3P��)O1-�ǰ�']J������}���&�o����B�����%Y��<h�U9k�DR�7qa�g��Lv<ɪ7.�Y����^� \9����cM}��e��;���;;d��)�=�+����f�K7·��wk�����l�q
��M��{�5tkZG��Y� �gv��6���6��S���ձg��ǳ�t^��W��t�c����|��%�p�܌Kf隯��O]�?B��#qf�J�Tͤ���0E��4ZT���:c����&�#v���#�k�@������;w�י�Q���5�y%@���δ�uq��me��?b�u����$ղǨ׳f\e�V]�C+Ͻ��Mz�u{�h���8�����؟v�n�v(.�pe$8�S��bv6�42����.��&�z�8}+�er;�p�N����Lqt�)�7ޑ��D�t�׍��\���'��z'��{���_;�s����C�ϗ�"�ִ�\��κ����/�S�'���5������q��B&̭������b~����]���gKh׏/%r�w�J�dV��]���_ ��}*ֹW���7�g�'f�y�P��.]3k��j�o���DOS��Y�T��T�K��;�sNf�ܳ��ܿb�7�������XI�{�^�ԫ�=t<�W�.��kƻ7�r�����2����r�)i�v�����T�}�V͞���T�kB�ʽ1vp�7p]>�o\>�̶��ٱvE��t�V��E��V��:����t�}��6���B�3�t!����v����K%+�qz�*˓ �^�ӗ�qTX�R�ke䨙�����ݎrM�MCt5!�]����r�l==�>^�	z��=ݗ�yZH-vS��0"��'�v/V4��h,M�s4�:y�÷��ή��u-�����;��x���ۛ\��3{�6_�����,�i��Ưv_�w:�]��iV��E9d�n�[^���>u�6{1��$[��*��湗�y���dk�'|�>�E�j�B�g����{b��ލ�<Nur�#�;%|��*E{M���5�K:k�sB�� �Ÿ��"�E�:���Vn��������+�]y۾�����MF���,V+wNۋ�{՜��X̻�&���n�)]��u�).�wU��AU�k/hP?Zn��)s��/KwudU��8�2+)�˥���kIe��ڙK�&����,B	.U�}�h0���jH�����t�II�p�G]LdwҠ]ub��@
S��,`��V`�M��<�)�`�j�;�J��+em��Q�č�                *f��o���ҕ��}D��AH��7����@�bi��X��|�R"�+��\��^�ԩ�r��Ur)mq]Szq�@�b�N�g6G1o���r���t�t���z�V/M�%v�e��>s�̪m�fmkx�7��0���I{@𡕚�h�QV����sCpry���؍�Wu�.S���O(ه���;���hu[���f�nmaÐ����K��Q��?�����>��-�rH�I�"��	F��D�G�%UUJ������*ƪ�4���+4�0���\��.P5T�Z*����i�E��Um��Q)��Tj�UR�T�Q����QKE�(F�Z�*���]�M��U�-Uʪn����W���hZ)1tYL��M!Wwum�*�(�[-T(hQ�;�{��o�^N���5+}ۤ��MY�IM��O_w]\��k�?y����»0�Fsk:d�[R�_��0�ճ�g}��<U�}�!�J�{Ji��Z���.ש���U���U���l^7#W�'��.��z��}ֻ�-#U�=��{u��3��À編'a۪+�J�k/�o������횫�l�j��Ǝ���ʉ�3�EP�k3ý�tǭ��ǆ�C��ˋ6r*=�ool�t -�[�������g���t�B�9Id��w]6�{���M��k+�5=ܚ�eV't�Cد����{=�՞Ҕ5SGs����ެ��H�6G�x5��+��N��~ݝgqol�	�[�.)��yH�E���;�n�|���е���Y�z�}��<q��'�.p����>�8�/}�ozLa/)����=�!��@�c�|��6��L'����=Ӕ�թ�:�7/U7�ܔ�[m�29�9d�K�����9�.�'ұ�[�߸�����(ey�d����^���.��2~殼���ב,pb�(�`�T�".Ii����N��W]醏aږ��=�f��TAV�U�|_s��J�wxM��k�UiG��I*�W"7����=<��w�s�W�K��Iv�}��ͦ�l��;��s��}�;�ϳhk���`V�>��v��ꔫj0Eyn�"d��&�v�#+[��\��,���V`>dyV����.�s�v�����uCj��~mus�ejZ7���c~��V�Sq��m^^Py*uc�"/�w��Ċ�k-X�N��|ڿM(�~��ԩz}���7����vwz.�x[��-�7=��\�a�ސ�b�1�ټB�e"t�kc�'6�m�k����x�I�I��.H�V������ܜ��wl8�S{�p�0%��4�ծsJjP���7+�5݂("iPU7#������|U6��Y��kww���o fy�EcQE<}[^��^�W{�]���L�^C�v�)����g7y<��h�E_��k�U��7�sNV�X��׾����ܸ�kr�)���Tv{���}�������x�����+/����D?i�WM^��ھK���n`8K�y���妟b��S���pE�Lu�w"�aw�;h�~���|�@��^�1���N�>*��3Ov�.�+�W�W���@.��ʝ��X=~i�6�7�C+S�>��O��8�SJ�J�n���b�~{����t󧎿^y{u�*�S��2�N�p�����-|�W����[But�QΗ�FU����M&�ކsk+��&灖��^�I:���;�8$hn��N�]�tN�)����s�L�R�lj<��E�j��v�_�z��Hueo9�^��C�W�l�Qݯ� +����W�w���$UM>ʻ{�k��l�no���G�_�6�wל�������
�
�wT�|�#���ۉM=�Bhx��QyG�ė��q��/�߸W2�Q^���~͔�Y^�v-q�����}D�K�s�/�q,����ʞ����/�1Y��_E�B�3�>��݌>S�rGkZ�T�j����sz8O�{�dY����'9Ь��r��7���|�wEL�O�<��/�I�{��T����S��t�=�+j���l���<XQy��کGgǛ�����A���t��8g�`�d�f|
W|�˖�iE�/eI�E��%�q���%©�/<�ӛV��x�k�Hu����:������>w�=c�;C���] �Ӵu܊��2�Ci>81�բ9;�N����g����2G��LJ��I��R�F��b��?ì?�����{�C�B�����ng=��~�a"m�u�@��hol���3�k�\�g]���#]��Y�^����؂�j ��W%�~����#⩻*���}˗�n�os�_�����E=gϬ��^#C�X3�}���R��n��]-7��߽�P�I��;�ך+�5�:����mS�0T�M�ݳոR�� �zu�+�m��:�V<[6q�W��|H->�f��5O �~��ĺ��n��A�e�۷ի����6����yğ�2u�n���Ә����9�\�c����o��Q3/�t�n���*���;�x����۾q�c�Po���V'/�A�q5�E�,�=��J�ng:�#�I�<�S;�詮��}_�о��Ç',w��˭+��A���L�%���p,u�fҼ����-PP,r�F���;u�VMw'Q��^r��t궣��BR�E���Vm�7ݤ�0��)��u��n㇐;$gaD��Pq��%���K�"�e�޾+i
h�"u���r����m�����Ǥ���PS���ffZRt����}k�;�6G���Ɩc6m���k�c�u0xbT(ԫj����62�S/T������I4�a�+F͵\�m�W�:��~\��+������{�               3^��Ǣӗ��ސJE��w�4�F�r��n�[��k��]ʐTEu(ٝ����p�6v�yt� �t�c��IQ�xf���v�����&�XU�hvzNn���J��c�t��#��ӹ�GlL�'<{oO:���|A�m�H,i*�9�'���
�7U�͍��-�����0oi�#���kb��/���x�s��4fW5BT*�(eeh�Z�\�E�K��z���D�ҭ�rN�D܍~���� �ChU�UX�1�i��l��,��-���j�B��
�T�j�KD���bԵ�)����m5WVU�j�)n�m,��\ݍ�K��ʻR���m�t]���P�-�)�R��-J�MEA���(Z)J[V����4T�Ji(��d�jP*�B��P]U5�n���#T�U41i(���H�Ut�iI)��֨h�iwRZZKJ���n������Yb����+w�&h��'K���E̊u����6�V^����4��O���r�Q�x	cC�U�T�{]s��*�=ّ���h��G�.(W�^�x��/0)`��u���~;�!*��L糌fQ{����H�������Y;��ޕ��eo�E��������|Oz�΂Ni�Hy��i3g�f��s�����&��x��PS	���xxG��sYw�mbKK�x#�a�&�A�9)*�m�b��]�K͎(�A�vК��'l�>�Ŭ}L�Ox��Ϟ%����ֱ�~��-��I-�[k�K��(I"qU���u��O��[
�ʰV���[����Vyz)�|�R�m�2&(��y�����؞���Mdac&{����o�E���޶�L�^yL��׀w�pk4Fʖ�;il��^2evv��J���Χ�)�#�sL��1{�9��ߍ�{��D�F��{~�|�Ν�s9�hH|o�ռ��'#���=��|�䎏+i�kS��TY����=s��vv- kۦtL�y��m0v}�AQ�<X�7㝷�q��z߽-{���e;L����=�JF�^�s�޹$�3�}��~t_N��'��ݻ��^mz������B5M~$�[�<Ru�9iYa��%fJ�:I��G��ᵯG�fM�[�p굶�9+�=0W�Q]'���Xsw�9f�����S������@�q���::H����9���&�f����>���zm� �I�WsmB9Q���wu���N.��v��⧊o����v��j���ՙ�?z�V��~����6�/s]��y���=Ϊp1O-M?|�h]��>��U���oL�g�	�FM�t��F��f��a�+\� �+�Y���Y(�$>J�X֌��W/�Eĭ��l1t�WI��>�Mx���7��I�:�T[Ug����:o=��WW��u\kJ�b���8��5җm��b{��]�9-禨�)غ�c�;9b�ܩCv�|�7�u�x�c���z��G�g�UԲq��E8��)y
Y�{b}�;tKQ�kJ��q�z�w�t��$�2aٔ�����|��Z���YR��x��X��|�6w-^J�B�Ej,΢s(��d���宜��a��ŋ~�ƴ�V��=7�9**��i鑀Uw����E���=���m	+Ը��K�VqQ���4�������}�K�~4�׺r�}�㩻�e�m��`���E/+\�Ť��Wy��-�y�Y ���D�),ݢ�^f��0�Ʌ����[�F����۴�l����t��Mq�&n����/ap�:>�79�ޭ��9|/2.�y�c����o��0��#���m�g�3�O�*���T����6{OVȍ�1Y�g��MS�q�w�~C@�#=�[�7[���ܫ�C��p����fv�(��f�m���/�ߛ�XR߆�}�7[���S�o|$�w�ҧ�z��{\�~pTz����I���B�{�eڋ�,��a��v�GH����e�wX��Yép��V�Xx�7v�e������v<d�t��o�v9��p[n@7mM�.��+����젖w�*$���dp6�P^�����YJ��sꋪ��ŕ����w�������X㞼�~�pEMm�T2�W.�_�z*y�]��X�#�p��A}��I�	���q������)O���w̲��|�]�M�0Q/_g�o�GZ}/W�6����|o*�O"�y�Ir��C�Ӭ�dcz)�e�p{*�
�ʎM�Y�2H�k����\|��뛷x�yq���&���|�~9����֨��O�wX��{}
eP��)	׻�|��gǳ��=��c䗭��x�>n�,���	�D*����W��ֶu*�H�3�݃Ӯ*ڣƽ�:/;����w�6�N�YA��<��]�+�7�]�vy����|�:�P輟*���//yc�k���u5:+�U�u�T�w]hp�����ƀU�i�I�Y�ѽ�+�_=��Ң�5��Ge%{J�d�-wM5e)���}]WTz�u��I��?;te���P����7�䫫�h��r���F����]�x�qSZO\�r|Mc{�%]��> )�JE�w}`�m؅��E���G�% 9��.W��h*�@��B�P�	]��#.*~��Ν��V(����Ԟ���U����3�y��?��
��Ҫ(���A�@ 	m��`@ 	��
'B  O������
0f�^��bC��C�0f	���B �(BHH����
@���w��/;.g12T*�XT����}(�?���FcR��H�aRW��O��  �E��Bu������~������B�K��&C���ϼ"���l?���E�/�Y����ߋ[�l(���Cy��o�@ '��=����/���;_�$� � @ '�&� '� }��¤��������C�P}���O��'�!�2Q�_K�.��y�̇�P��F���B  N��:�[�?X��d,6�d,�?Q�I�!�a(����d���Q��B��B���"�q���? @v�?��a�ZԢ���%  ����S�&{ufR��ƄO�!  &a��䓠�T�ܒ���F�aa����قi�_�����~Ѐ �&�hEY(����	���}}��?�!�U��~ʝ&C��a�O��~�O������?���������Ώ��#( ��J��.��C�h�d?�C��p>���F�����h�zHPl!�������f���.I�ɐ���g �����$������g����~A  '��2 �����D�!�g�$���p,D� (~��xB�UHc� �%��  ���'�����'��Z!�:a(>�$���PH}L�2>��4�Z �A'��c�(��8O�]� J�&J�$�	!�xjL�����}���I@  vB{A$֥O�%��!ٰ3�%���0�4H =,?������C��  G �3��H��?/��ğ��П�����x����O������A�I�1D��(���~����~��͇��!/�C�Hc�~�9���  ���Ϸ?��_�/�!TQ ���Hr� *O����������C��??��}�>��Y�!��~�Cz��2�����"��A�Q?���~�����C�����O���.'O�g��]  ���$>��?\7���l>�������
����	�|X~(C�Q��U�p�@(?�2H~ϐ�F �#$�r����q�!�?�~��}����l �r~�'��&����TMsr03������ԇ�!����Q!��>�'϶n�.�p�!+�*