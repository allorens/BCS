BZh91AY&SY~e���_�@q���"� ����b?~�      ��"��d5�% ВTU*�la%4�@�����+@��`[P�T $ѶSD�I�� $�ck��ʭ�u%,Tؕ)lUh	�6حj�k%2fm�����iA�m�f�J	��i�Z�R��U�T�fX�il+l%Zm���7�͓u\�UIY*�݌�k*D�8v�6�i��*�m!j��UKi�[l�V٭l�Rd�ɶB֚�[jRm&i�յiET�L�f��Hi[�g`��UA5�, �   ��z�*����� �tӕZ+]-��u��wi: �����Ӭ�h�եr��U·]���(.�bZ�ё�ٖ�0ږ�dx  7�
@su�����fp  ��@ A�1�(� �+�P �I�@  �#�t���@U(`t U���[Z��Sh�	m5�x  ����  �y{�� ����R �	��{��Tʽ�����G@ v.=�����x= ��Sۃ� i;�n������
��6�Fj�l32� ��CA��W^� ��={ޔ(:�������vN�(N틨*� 9�w@Q�j�N����P��wf��Ր�V[dhf#�  4�@i2���� ��ۙ�4h[�p�����8�l���5��i@
��q�@:Y����a�:kr����VlF��ٚhl�< �� )���6ƇCv۪�t: h�ӃG]f���Ez 0�@5���PU U�� Nu0t%�dn��@kwH��VY�YS(�Ym�C[�۬=݀��s���u� S�5�`� F��v��  &���ӄ���
h � PX谣�+6j�K-��[i< kǧ@uXP Y tnˀ�P��q�Tݜ  n�����[p�awg  7]��ہ5��V�����Zm^ #ހ wv�P 9�  ;]n
����h�V ��� 	��T v����r6�U :3E;6�J�تh�T���<   ��<��T���j�Q�Ӏ��
 V�7 ��٠;��t �\ 6�p�W�        ��R�M  �b` j��b��* 4  �  D�2�T�    hd ��R�@=@    Sh�mQ�����@�&�hh�`BT�jI&!14�mSFM2by3P�^ַE�a2�'ĖT��H����h�ҋ�w�w�~�=��^�9�{��QU���� *���" *�����0��+���O������x;T�����媪�>�UQ_�	S�J������?_���~l�e3)�L�fG2�9��&a3!��f2��9���&`3	��f\��f0�fC2���&d3	�L�fC6d&C0���&d3!��fC0��.a3!�L�f0����Y�̦`s	�L�fC0��̳e3!�L�fC0���&e3.ba3	��fS2��̦d33.a3	�L�f0e3d��fC2��d3�˘�!�L�f0���&d3	�ɘ&C2��̦a3fd3!��f3�f2��`3��fC1�I�2�fL�)�U3(�eT̠9�00��As �Ps�a�*��0��Q�D3 �eT̂9�0�fL�)�3 a ̣2(��)�E3*&a̠9�G0�fQL�!�FdT̈9�2�A�#�s�`A̤�3 �dD�"��0
fL�)�3"9�I�G0��W2�\� f2���2��P\��s�a�"��G0��&@\���U3"eT� 9�2�fQL� e�(9�0 �Q���Ps(aa��� � ��2 �P��s��s(e̈`3(���2*fL�)�A3*&aT̊��0�`̓!��f2��d3!�f̆d3��fC2�C0���&c0!�L�fC2��&e3.fa3)�L�f0���&e3�a3!�L�fC0��̦d39�a3!��f0���&a3��fC0���a3!���&C0�̹�̆d3�L�fs�fS0��&a3	�L�f�1?���t�}y���X�u�W��3�#���Ɣ�`�J(���r�^��4Mcã(���"V/�OL��R�!fF�=���1���K��tp&�qfn�&޲�Z��5�t)cs+v;F�G\+ f[�u��2�:�ݨ�bpVnf��r,��B��KR	�Le�e��]�����{�$<�0"��F]5iXrV�]#Ni�+%���G4�T�)�݇�ٔFwAf7�5o,)@�{3e<y.��Hʹ��D��T�Ne�ݑ9 Sc�U�n4���놙�FSz�-�І�4�D�E��'��BNL��і7Z`��9Hf�JON��F���v���f�)�YNf"��?DwwM�Q�		�fbݻ�#&�X������1T��F��u���E܇tS�&�����ҫ	�4�.�͙TY�̏&�����.�&���E.KŽ+bn�odF���F�V�M˼Us(��м6V`:�(5hh�9�4^I��5Z׌Y'(��MKt����u�$Z�6]]���m����eE{�Z@�ң+t�L��	�N#���a�-6�U��R�]]�T��֢�ȏ���:�;��b�\�c������sm���"�4*%vi���od)��;�*m�5IR����el��xiX��5�.lVfa�n�s7^VV:9��t��PPf�Sb
l��a�1�ʷ�&��]Һ�Xf��qdò�u�� �ǏK�δF!��&u�˚���CJR��R�^��]堩��$f>5�F�x�kݷک�.��ڦ�dYU���n�DSX��m=x�Q�����O���
����3F)�ܭ�t�ZU���N�"�!5��$�!Z���̻u�2/u�zmZ�R�E�,k@�-���5��j���"�BpL��oa0�4�36��Ҩ��(̛������ω���n���������tdw�r'{[)wb��?9������F�a�lũ��юG�=���^��	���A��V1l�n^����N$��r&*��YPT�"�)��K�KӋr�7w�c�2Y�4ؽW���FqB�����A���	���x^����L]e0��ZǪ^��ku7�0P�U��jݽ�e�n
͸u���;l�Ϫ�	���)]%z��X�o(���H��U���x3H��f�Q^�`�Z��l��{/H���O��R�v�w4�l`lj�2�����b�����M0(%r���к;d�n�3[����ݭ'���*d��=��!Ȍ~�fR��=u�;�I�
���%�Vj�G���`��%����x�Xچ�ɩ{�Ø��d�hAe�[�����v�i����n\K,��t�v3r捵L��0R̆jZ�W�3	6�l���赵6�ny�ֳnKvf�8n��֋�Å���`=t��x^P��#�ئ���G��M[���2 ���aBa�F�����͠�J�#q�r��&%x:�\�]�&5eeI\o@���ߌ7Of�4�I8B�c�hI��M��5l1X]fCk��p2.��Fp��/���W:�iR��e�.q��F!2���Ri�����I�	T9����IDTM�� sc��R�[-�V�[k5�"F�n��kMbэhfL[���)Պ�[OlVa˽�$v�!k���Ḙ{�����Č�h�K&t{�3��Τ��ld%��Ħ4��^�ѥ�bl[���V���p�tX���# yN���)�Ǜh��2�7a��y��XN��Q��"����YH[X��9[�Dw�EZ�-����3kN�-Sqe�x
�j�' �=�����s�R7z6m�I�xD��.��#�4�M�YZ����9��q���ޔrV�m�,A���kD�h���.M�F�#jC����7���f[h[��p�7ڻ�j�b-�`:
����0*��h�+�2S7${�V�jA
��sDYt��ah����1�{`"�Kp]P�Zt�e�������Cy�`�M�P�5k�2+n��R�w�(LrA��5�$�H�9,hH�)E6�&��Gwq�e�u0����{q��-��q(��J��̡������7�Kr2k��V,:�nMu�9Pމ�!�藗�W���PI8��#��/�{R]������.3���ŇF�/��Ѳ��I��˗���XX{�^�p�.�f!wKRa��"J"�c+K�X�G���j�0�qm��D�7̌M���7I��
hF�b�@ؼ�11�c���:�e^�Ѭ҃��+u�cژ���cЭ0ї���Y[{�����M�v�J���PAQYˮ��5�ذ���n����N3�v^�X�L6ȴk`�{&DU�8��w�f�.��ذl�P�
��.f�j[���Jʙ�V����oH�1�f���#?!ch�6��"�Ja��$�XW��7�+w6��6�1{/vn��������R��;xo�J:���tp���e�0f�l��ud�����r��4�^�YXP��a�籓�[��{0��qh2@aE-�V�GwWky�����Z�2��e�m��4TZ�	�{7cͿj�X2�5LZ���k�="F�_���t@rD3!W�iΒn��wW{����e0�d:�'a�V�k���n p8��ͩn���B�N�Y�"�#�r�o%0�o��f���Y� �K*,����dt���P/إm;�zm���Iv���L��3�/(�/��	ڙ�Zz�/�u�z�庋@	���I~����vfa�^f�,3ڵ�U^`�)�F����+&�$Z��)�kPNh��d*�`�Q(P���D��r�����e���j3��;,@-�a�ڪ�j�5-䫹������L����7yKb#Z�6ێ7�hSoZ@�.�-�"�lmEt"�.
"�l,7��]4&2��b��r�h�(�L`�lm�똞���̰��DE����UVhwa���:���y	Ctv�^�l�@���`°��^iY2�qKZ/኱�B0�P����Ql!G�k�t%��A�T�Z-,om=z�7�ںhM�V�Ӫ�hh��f�B��a���̧�u�9$Rȼ��*�4�T��u��3*��f�ݘ�?#�n��bi�Or#������/
 ��ô򌕂f�0��"���`�v�8ni/p�-XL:�U?^�^��Мb�	�œy������ /7{��\�&\fE[aL�lM�2���{`�wux�p�K0�$��F�����d�l�
�[�KG�=�:�sN0t7�]ƶ�����ؚ�����"�И2RrK�Sf�f^�� �im��qL�L�2e�c�C�퉌�˼fQ��*��R�F�,=��ˑk$@�����g`h˱�e<�{�ܦ+$�n�W�D��Y[B�h֍q+��KvlST  �s&P��/%N,ڼ��®�L$��QS�Y�>6�^<�X�e�����+�MR!h���{N�ǌ�Sю`9(���p\x�1;�8�&H�{���ٺ�wk�t�3$��v�1X4��.����i����
�y\�i�!7r�'��@̻�Y�����)�V��y���L�l�xa�F���Dfn�p$r�X��r��rf�v.=��@ X�K�̰waK*�*#F���AU4�&�Z�x�Ԝ�.�GN�2���*�b��	�.fU�	t��r�0�d�Mb&S���:�&��]3YW�˒֘��:���ۘ�R��닧Ma��I�)�bT���ނaܪA�F�p�Z�ئne�i�32��[r0�Zov��4c1��K	T�:���E��o���Ti�V+���"vC����ɠ#x85귰`�K̭Ӗ�n���a�����uX^ڂ�N�{�W[�.:B,M6�s�b�=�S��Fm Rc�WUV�+��K�&ucx.��Yr��2����j�$�1y�F��#�ۙ�YTt�p��lV�f�0��x�M��jA7�3r���VXZHq�BE%Y&�ˡW7&�z�-:u��F�GX���8쉄]�T*ʼ�owle%D�q����f���;Ʈ���V�E��1��b�(*��i����N�[�Q�5� =Wt1^���5�B<�[�t#Jl�C4��H��c�U�x��B��Uڧ@&*�ɒir� p�Eh��&��s)V�1���֒�
�k�YJjB]-n:�z�a:�X�Oj`t�V2����If�7SPp������,��XV��!�Ī���Sk K�S�2�cp�*-�=�6�\��f�kN��nf�h$7����L̬oF�3�A�^-���Q�����
�!-���ՎFM��Ʉ���-�6l#Q���
�oF��R�܂a;��%QMYw�b�&��5&�8�d��d`����r�Nj8:�������!�׸��.��	۴wEh��+ QX�i���۲����l�h�X��s1�'$������'��f��l��KxE�t�D�:��Vsi�8�ܶ3m�k�kcZ�����x���l�)Pۋ,3)��e_���/)�v԰f��U{��L�����Sl-F˫��^k���e�XT����ٸ@�N���a��*Ǆ�m3h#~���8��2T�X��c[/2R�H�0��$4�cI�ŏ	O�y2��=l2��y;�;F��iM�26c��~b�0��&��l߶�o8���
n���2�.mY�*��)�IL��u�svłk�Eu���Tn�nf���՝[Ɗ��c���ݪ�3�����E�۸���,�x���ꐳ�KȚ�j�^��,#|غ�����M�%�;7Uɘ��4��L(Pm�Ӓ�nB���2�y@+mS��F��ha�W�]6�,�f���*U�N���i5t��F���Jey��c�+E܎�ՠ������c�/wl-�Pn��U���W���`�Գ_:q3��ƭ�>��*��oեY��(J
J�']�[���殃���@�P^Lu:I�E:���͸�f�h���O+r�G{��ne�%t���T�htmL�	���Z�I��	ʑ\t6X �Ro���-j'U:TX�nȆ�#U���[W(d�*nڣ��u
t�Nf�(kh��Ir�f	X��ni��͚qګc��F]
cʵeջ���[MAt�Y���f�Y��&��I�����ě��h�ouOb$n7lՋcX��Ypv%��&�����oMU�ӗ�H�0��GaJ%�j=ʵR&�� p�w�[�^P�ɭ5LbhY�N͵3��N�EZ]k�pHNG�ۺ%R����W���`��p�C2d$V:�6�}.�FD9j2uh�a�}0+�6�f$�[�j�d��r=�0�����ؕ[n'@;�M�%�fj.�X�iXY�#������hQ��[�䣴���4ۚ-0X���-nT�񊹴^�=z\� `�6�Y��̅,�$�MA�2�,RM�[Izj�Ń9c�t�Q=��|�
��3���̎��Z�ӡ��j�1lQ�#�v �̥e7*U���L���m=�%p�d��BX6(�IU�c*[����Rxq�Ռ[2�e�z�F�,wz7|)�'n�V�U��Y+u\�A�ʗ�����V�M��b����dl�ɱE̶�32jPŰ���Ӯ���i�����ӊ�Em�/Z(�՜Ej8��aCe�
J���6Ŝ�z6m�+V�{\��6a�,M�IB�ܻD2��1�r�%a.�-t��X�z�[������ucsl�OXk&��1K4%�hjӂ՜4��*�a�Mԓ�B���U�+-ॐ����/]L�Z4Z�hݙ�0�����r�;�%<��uvW�v�cW*�N�lm$6���N��'�4�Tə���]�z6��³�ѽۚ��nܺ�b$���rX��{�t�@�dԩj�oU����\2�"�@Z8�n��w��-bn�-��@5�<$���^�[�t5�[�Z-2ZƔx!w�y7�&�p�3E�-�fc/oo���U����F̠�]�1����
�rb 1�&֊j^R��i4�:U�u�h��.���%gP�aX�t�XӦL��]Ŷ�&���饊�d&�b:�/w/,j�/07�sj�r��n<���l�՗���t�	�a�7S��9�#8�D&V	��;їV��.QU�F:)�vVa�Ea��A���`���;��aʂY��j�AA���Y�0��a�w�lZUL�؞�{OpŖ�$2Me��JA ��ؖ}R,�;�Еj��[L1n�Lǚ�ҶT{�Z�O7n��0V��(��+j��ZgV5�j��=��5���v�,�g �]4���)�<�ń�WôTt�����2��^�y�(��0^�nt`��r�o#���WK]������m%%�9k����bk��������v�{���mmLG�L�{��f�Xn���J��Ŗr���3�6f^(Ji�Q�F%h����"]�]��u���G�>��"Y=f˶������������I��7�F���`�ڵJ</n��FtԊR���Uw�wTT(�;.A���4�,���vw��8w� ������)�԰x������KG���%��kNsC�d�DpR�YH��I��U�\i���!�r":�Y˩*D�9
E7F��dh��K$�:ʇc�7�ˢ_�=��6�s"�%�e,-�qKbz�-�Z9^q�`�SX���|d���/R~u�܏#�}p50P-�������
�8�C\pUi�� �5Z�:�d9u�%�JLR�YŸ��L��N�B\[s�U݉�v�����%�M-���YV�Z�u�y�H�7��g:�A�z�q�H��/-������z�ŀXv���q�"��(A*	.�3o�s���|��KdOev��ԭRE�8�с����%$ÇwuBt�+	g,�W��͏���[��@~��B��K0j�#�~�������'Ff���e�N̻;ù��H��%�ha�x�FmmӧWg��[I��ɹ�%�6�X)S2e���e�#�t�;#�_6|���}9��I�H��G�#�ڲ���)�:�\����H�@#�d�Q�ڎ��Ѯwv�^|��{7o�����r��=�+M�l�U���6z L,�7�v��\©����)4�*��*;�m
2�:�[GR���;ДreB4(P�sP���S�V�Y�O\q���wb���W����1���6�u�P�NM�)tb��	ie"�A�At�����c�;JX�-�V�j��������[�о�w����m_��2s*^L�4��lnb1���4ȣ3E	��z!��Sᶴ3��X�Ta��I$�f�W�-��#����Ɍ��#�پĹjB[�ȡ��)���x�K���]�GCjX���.֜�H�}��N�-|�x�y��O��̕T2|�����T[�fv�K�a#Ac(&�)�Lt�����r)���V�6fI����0O-���,v�S�,���i��N�uu�y�B�q�����uT���Κ+����9'p��lwy.�	����-bo;V�Ma�v�WdN7o��x�	Y��fNos�����h���̕p!�zW<�����޹f�8���ӥ�겘��$��M�i�^q1�X��b	�!w\L(�m�A�띎���"��jbj��֯S�<pu�;���q�ω[�dYu��<CDń�5�t�b�#�YX�D�f���3�����yOz�s��\���L���ުѶ2��E%�칒�]g���N���{u/u;��LN���XK����6k{i^�*Y�	�lX�9KN��Ğ����k88����v$2�mֺq�N�9i�9�ٽ)��@1CfurŶ�/]k��,���ݛ�2[����]��@��iS�j�dѣ���phY-�	-$(���\�nC۹0�g9�֩�m�hg]"3kv��v@�n4�����Y4��C]-��uǼ���ofr9Ih"T�1�e���PJ���^�C���Wϱ��|����B��Ӑ�ˁ��Hxҹ\�ּ�`�{��2��j�t2�;@�g.�����]���4.C�����	�A���޻��h�'+�<�n�)^��)��vM�ƳV�mG��H����C�P�� #��b�9�u�ys��h��a��+�-���v�M�!�'\n��!��.�Z�8�f֝��a���w�r>{ծa:��+���^m V��������=�Q�u<ܨ=th3x��{��M'Ҋy+���^�]=�����%���.뙮^����I�}��Q�.��^�.�f���{f�]W}��'h�	�z������ۻ��@�9�
�6��ܵܩ����1�4�0�c��'z�^�����/֍�O{Cʺ�ql*Κ�E���c/Wfjv�;��4�[�폊w1���Q�v�7�c[[W5uDo)�SN�J�cՖ�nCӳ�Efy��z`�{U��u��\h��T7U�ժ�(���U�o��h����Xk/	�f	p'v���9��Yc"��	Y�o8�pK���{Em�ɋ{Dͮ�yқ.!�lr��x��9��A��0:���
�[HI;wtES�g�tY:fc'摮G���DN�d��ë�Fh,R�s�Vj�� hNK]�Z�Un��B�v�Ԓ�]�7g���RBlV;��5#<5�	"g�η��6�g-�T�dj��qRQM���"o �f;��=V��d6�9]p�ͺ��6̴m��*��==��6lOQ�ՠc���d��¹V^���5K\�C���/���Ԕ��_����}b�����O���;�
W0t�p����+2�&�t��"Z�Ŗ-p ����(��#�2bP��sZַr�-}DW��WQ���Or�
�kr-�<��⚖(�uUѪȮ�D�Q���͛��=4bW�;;��z*�ꅃ� �Hǒ���_odG�;�3fɇ�t��u5:.�[�-���)�4�x*w�+��)�widԅj=ӥuI��:P�w�Fm��0�?��/�o����F�ZW��Vx�ר5U��$+�ޭ�R�;�Zwl�A���RbP�-𻻹5��b�'jj�u.Uj�ʻa]�E�̈�����a�uA]`냪�cyG,͎�7QIV&n���>}z8>ڇ�UX�+�����s�V2q�귵�;f�����4���oH�Q_T��r��`�	Ms���m��7�1�!�}�~X����T�F�*��8\�.���Cj*����d���fZ�ڱ��F�U��P��
�Dn�y��]	�3w�R`���ugdRmPt̬���*�.�]f,"a�.ٻl�Mu�7�e�j��u4�	zx��/��i���Xy[20��t�a,h�yλ�����˽��LٽF���E�r$3�4B�8��nD��ᯎu]����̅D���F7H@��m��E]�niE���d�ix�k-��(-�Nb���W����kV�t.<JGT��h�Y� �F�vB��m���5U��.S�9*܎�]n)�#��������BZ�p�Ã��4�h��3jf����(XȊt����+�z��`��"��i`b���z�X���>����\��TIu�w����[�3Fn#��Ry!x9У{�N��9+F��o��ZI3#������y��35��*1Йʳ�cRD`����sU�>x��k&&o�ئ��[��}99�n,�𪂦�@�ole =&�{ݎ.�	i%n$K�P����lW+�����W�$Y��Ƅ�.�yE<��r��W�,A���:��v���Sdnt�l�M)SM�SMq,�޼�b������u��F��A��aЊ�޸����]J�L�Wmd{I�{�MY.Ѝ�xR��ngX��ou�CIX��*5�!���2^���nˬ1�˵0��ԣ�G�	p���1�P�F�%J�,�FY���N|�v�0�-�V��R����qm�Gw�j�j�w�ҭ��ݍ�S��%��o.����JM�Od�VzL����{�w��ëά�GEs+�{�jsٳ���#x`��f\�ٝ�fh�4�3Zm�鹈v��,�+���X�s5��2�u$Y�;/U�����*Y ��:׹�wl�]���vlp��܏Z�[d5]�'u�/#�{{�:��{�01Gz�Z�@�ŭFm�ޒ�H[Khn�H�hVm��S�[����U&���<5aW���r��{;�n�Zx�y��O���nr㊲�2���K�.��)�h�J�~�N�a�GLU�+��n#��WR�{��bm����.�L&���
`%m3z%>����F�s]ĺ2v*��%Z��A��@ںUw{���I����u4h�3����ïU�-D�1�$����\oRD� GSVH�P�����Sh��k3���M$���hC��sv�Z�!�0���x�7����܈t��aAlq̈���2v�Ў����t��]gt��Gg�:ƽ�������^��!٬�g)F�x�Y��Ua��݈�c�sڼY�1`Uӱ�~x"�ck#S��9oi.�����kR�Y��nv��I�^Q��j��2m�(w	��`�kD5A�̤�9r2u����O�v|���4*��X땹��4�"�,m��.�AQ�-#׸F�@��[�ɫJ��UR�Tfͫ\bSe
;�2��[���6�@��͈������  �Ƞ��CK7t�Qm�!ɚ�����*{�_ZO�D���BU��Y�Bخ����\U�l��W��_d��b=-����Z�g`�-��*�-�[eT��L��$ڭR16��^a�Ղn*�/{LyM��ֲf��B���*��<�W5ˌK�/�Ba��v��30i�P����'0�a�.�5�C�c�,���8�����X���(Pu���;��;�#�����JA��DD�jï[&��/�,�q =��e���_N��ĒZ��i�7���VP�d��M��1(�6�l�u�s���u�]��70
��9�w�6�)�I]z�Fn���d=u)�x�<�$uZi��4�ݽ�s	�MІ�Ы`��2S���ҧ+�Ip�Ω��'�Чb��*�*ܛͽ���k+wP�q�E˩g�x�GEV�]��U!�j���;x<�GUe;C5aɹ7d��P� �w��hH5ҹ�;OWX8b�o5�D!��x����RҀ�˹`�A��:p��ĥ�Xv>ƶ��wڊ�Wڛ^�/h��'=d���fL�N͍�Lؕ���S�S�X�eo*��
�NuG���~��z��v���sٚN�n�*f�N����K�h�1FM���x���aE}v�����Iƶ��t�nbU���\��Wݑ�nm���U��ټ�o�me�Y��vZ��SYX13Ou����1Z�^�*�D��_3���O�nmߥ�@i����ArYՆ�C.W���5���Ȫ�{7[����nj+Ka*�խ���ڙُ=��Z�5 "��b`�e�nѝWl�K`T�:����1c��하�������-�A�A(����s���ͱ]�9b.�i��H�.��Uguk�n��M�8��8���ڬ}�`ѝ+���\���lh�8��c�!�@O�M!��u�{R�a����M,��o��T��]�<�]J<[܌a����Xw��]8^�
�87�ԋ]�q(rf����ku�J�fM��F۹�٫��c�]��ȱ;����T+�p+���4o���ؐ�d��S4�]`���'�H(���}�x�M�:�1פGA��q���K�a��S"&���,��֔���2����F��=t��]b�g��d.���z��n�{&��f��l�L3M܊��Rs��45t<�Ӕ�����*�e�ml�2�����\��[��	�N��*�
������Vuv��Ĩ�5\��p�p����cyt���7��c��Ҿ޾s$� W.�T�Z���\2ЛU�(���zx��k��r�ʹ|����juUĈ���.�]���s����l��KȬ��T+&�s-QMp]�t�kn�nf!H��w[��U��׷N��fl�;Ô���e�s,b�a;��}YG1��NT헹b��8�u�w]	)��s�C���F�n�����+�+��ܫU�+�n�p/�Y̾qe�]�r_[yO�d�ц�sE���,R���
"Gqe�,%G�V����&�+����Y�a^ޥXj0{�����v1hT�Ǣ7���^�0�g�sJ��j)�vW��W>+3���-�B�jn:�ur>7�x.[�<��M�}\����zn�� :B�a�Z��}�7Ԫ=��5�m��,W-�)�X{lt
X���F��ܕWQ�x�Q��zg5�R̼{���H5�Ϸ8�`�S��mЧ���u���S������S�;{O�wu�4�r&w{h��R�S\��v��̷PR�΅v�;y�����me�2��G3Ew[��7��0�F�N�}�(��Zm�h"�acjoU.��V(�s:8�@��ŞXeK]�ZNK�^.�h�ϕ�#�5=����CN=�f�v��O/��7e؝`��j�xv�������w5/��6D��F�`��Ш���O��rb�K�n>�Vt��G�Ks����7JU������u�P�4x�[RHH�;��ɪU���"�����&���ڨi�
�4�]���&y��b��C���N���`�;�"۪����&f�nR"�<�֥W��:}�q�'�����f�Erc���twf�d�e�yT ;(=������%���WJ��;tJ�2U�&
�Ruhe�8�ww2�F��j��.EÛ�=g,b4h�I'�[�`��'69Ѽ��9a3YM�1�z��C����pw�*�'�$lu�}�q��:�_a�in�|�3sL}�����Շ��شmb��r��qiʋH�w��b]j��w:�Ջ�q��-�M�Y�Y֖��<���^K����9D%�U���iL�=(;
�ƥ�O�f�v���4 F����)����8�o��Wěvr�e5P�u��[���S�M��Q�a1�R��Qm�q��u:��DU���q2�U�5�2%l��oz���.�"���F@ڤeMx/3{a��� L������;��'%#�1U`�s�uDb����y�+�)���rS������ZB�����v��5
@���,[5�Z:�'�E�=;�"�w�h���Xv��Sm-�D""I�Y}�3d�����kQ�u���	+^��x��H��^[:�Gطz,�����-;��{�&9��"	�XRY�t�����Y�k.�52f�uh��D�U+�a�R�����; )��p}Yn�P����N
5�˖9r˱mpr���ۗ�72�-���kf_�w�<N��N��jLur�rv��Nlf�;�қ$/]���r*�*FՁ�?#�0�@�az��C�@SL�����ϑ��N���O2��,�h$���'�Qy����B	�� �P@-��u� �?F���X���5��1 #T@", *O�!���cP�-�?A	&�bT~{g�^��kV��*��f�^�j�ax}S���8ӡYd����0�i"���6^m��{���B����=�ǭ�qq�6KL�G�"`�cH}կ� mqFb�
�Y��l�� u���iߟ���~�ADA����U>���}}��O����DA�����������w�����؏�����yO��m]."Js���y�`W7�{3"�d��7����|�b�r��§wM�m�7�_^�q�483t�v���Y"��9�`�|�-�:o<�c|���!J]u��F�*�W �Ԯ�f"R��fW^�u�#h�L�L[�{dۋ+u�V�ˮ7	u���s��Ps���Eh)���6%����9�v�.m�<��̾M�繈�b�f���{T�A�B>�,��:*��
g��&궜�Y�F(KKt�Ƴy�P��7�����*�y���e�$���T����wӫ	��gRA n�J� X�M=���:�u"P���r���U�^Ȼetgq���4��L�wT��=B����N�!�D����ڦ���hm��wkő�5�7�5�먧����ʛҁ�jZX�nj:wD�YgPOdް/��;(>��D4Ȃҩv�=��v�U���;\�O4��u�'�8������X{�M�=Z4+K^�o^sR;D�j�����Z3F��zI]��j�a��g�i�H&��븁 ��]����9n�����!�h:Gn��y�ڳ�5���ia�g
cN�lr��s�:s��q)�VY˫�L-J�R��%&v%R� X�ֻ/�pJ�S���'c�K�5\<dEk�؊����*M"ݫM�>�ojmMD����x�=��1�/]�_o���}<x��Ƿ��x��<x����Ǐ�<x����Ǐ><x����Ǐ>^<x�<x����ǎx��Ǐ��o�۟o��Ǐ>�<x��Ǐ<<x��Ǐ<x<x��ǏO<zx��Ǐ��<x�x��<x��Ǐ��9�Ǐ<x�x�<x��Ǐ�<x��Ǐ<�w����{�pn��,fۃ5՛3�_c;c%D��O�tx�Un��Ǧ���']����S�!��;|�ͨ��Ԗe�%GH%�nDRRm�wi39�:7`̡=e��}o�kT�<�"�-��_j�gI�gS�!1�Y�B��UM�]���Ӛ�@f��杋�s|LT)����:���ƥmV�jÊ��\0����\o&�N����9AĻ.�v�xM�Cd��/�\�U̠�=�[z�';�{��oJL[ۓY�tI�V�7�i�4�X\I=�Kr�WQc&�+ٚ�u��/�����6��u˃ gKP�z^� ����`h[���cDS��>����9W6^UI�>��q�=��ܠntd��������8ݝγQ1��pUt��B�37'I�ׁ�8*\�
aR�8)�׋,��zR��ˣG�ʸ�PךS�Gf�
�J�jk`�eY�r�r���ۗ�-c�pxI�'Tx<���N��֛DX�w
5}�G	C`���t����%@Hб�Oz��Z"a{�e��4�+�o-g�����)t�nU��*���P��W�P�8G���5R����|��bc�Ȋ�l�Ԗ�i�ɃA�Ջ��8G1�\Fm��f�8,�*ʪՇt�쀠����<�hW�+�r����aNzlEa��3���Ä�qr�
g��5^k�'��~|������x�{x��<x����ǌ��Ǐ<x��x��Ǐ<x����Ǐ<x�x��<x��Ǐ���x��<x���������������ǧ�<x����Ǐ��<x�x��Ǐ��9�Ǐ<x�x<x��Ǐ<{x�<x��Ǐ����Ǐ<}<x���Ǐ<|�x����Ǐ><x����ǟw��.�s���Wd�>{ځ"ԏ��r\.s�d�oqҖ�j��\D��{�kD�V��s�蓧�"�j�!u�:ὗ��⩉KHV��&NY�Zw�m��9P����15W,�ÕMv�ٲ�]v��N��3iEu�&��y���0*j��NKZ9]$t��/�u�p �Q�Q�v�_m�U�{�3y���]�F�ra;�v�F*�=ab<�H����m@3Yu�6�Ӱ���y��:�'�����q�a���.]9e�O9��U�7/�X��-| y�&����ˈ�btC�4G�-�[Á��E!Lˮ]C��N�����M�l@=�t�?�h����hyyǶ$k�M(�m�X�뚖��i���s�9�-V�5�HeR��Q��M�0�|*�d��+{���Zu�ȥ��yHe1Zv��P2�c�Ї��;ؘ<�
�q�h=�s
",48��b�Ɖ�T��WE�Q��Q��F7,7I�W��(<9(���I0N�gv��SO1r�������s��X.�0�N�6,��z��.���n+�7s����U־J���]Ӄ9�<�c�'��ZޘlV��������V�ք�W�u�}0n�g�Վ��2҆�j}�[ց�� �G0����v��m�Ɉ:�V��|)8��M�S��oZ�e ƓC�f)LL�����m�q3�8��;�Z�`��]��(G���<=W�T�z�-���XF�ۉq��˨c�xv%���Zn�6;8U��KAręQ���{5�L�9�U)q�Ő#x�[F��{7�Ϫ�Q%S�Pp���f��5���^����ʦ��t��JܸR8�4_&�� �c}�r4Z� �7O���
4��[�o�2\L}un{�����R�'!Q�(�V�P�X���q)J,S8��3��ԣ���S:���\��x�����G��6��dα�,��I��»;���ǻ�dv1��Z�&W9;&�6�/��-�]����t�4N��L��O�v�"�Z�[꽽�m��tx���e��0�g���	ܟUV*��[,Y&l��M|�X*�����2�$�ܸJ�Д�h��\���ľ��b�p�"���?Yg��D�qsz��gu+I��>����pt����s�=y}Dn�qRL�M�Cn�V�w�����0�α�	���IGѺYP`*�琜�TOQۖ/���oe]־�]b�Q!,/jT%I�R^M�x]o0�+���&���WH���w:8ͬČQT�ri��Y�+1K�Ac�,�]���8�Ѽٲ�w,*��W�ڕsv�9��*B�3�xNȾ�t�1��E�5��f�¹����]���m��(��e���aش�����:��/3���X­Õm�<S&����M����u{u��s��s�"{�8)��-��M�A�״o5U���S�0��NM�:��|�����R���XN�n���3KK��VE3�x��:,o1k�Rn�H���'RX�S;��u���DM�.��5z~���s��:�6r<I�y-��kL���WO�.mbi�ɭU�v�r��q@^��c���y��w��5eDs���r�J}:D�t+U�%�l�W�.9HV1],��zZ��pS��^�%+
̰�C��V�eY�����3�w�&��g%�p�G��귲%I�F�˨b�
�;�l��ݹr:�Po��ȝ�G���ɸ��+��Z6P�~��t�n��(�I�y<�^cg�^u`��Y�A���^K�jr�	XB����P�V�o{Z���V�E�}N�-�Ο��mx��ؚM�}�e��ף��vt\�C�����T���Vv���6pr/MY��#���a�v��qs�s:�n%���:(��b���+r^�qn?�ڤ������fj�[[�+\ �-t����:�������6UA��M�m3�ө!��6�Qܰ;6	;�y<�pȺ�R�=�� �xjdV���/�9�I���
1A:w<'j8(�al�]Ƃ@�F�c�cÈ>0�U�T��Y���ET�F��F�Xi�P��Z�S:
� ��j� ����XI9�9���[�\Jˍ�����u$���\o�.�U¥w2�x_`CWP�{`����伡���܎�u�kJ`J��
�5�T3K�9��FEE���v�y��Ct�:�]�#�Q�{T�HVt����ffo^���*��fԏmK�5�yGb��,̪�C[�8�W�XP�t��Ν[�{����EeΤQ���M�]���$l�a��ЖmY�k�`j��F�O{���)�
�v(���.�*"���;�B���(nˏ��t��:֫��1w	�p��s��M*����<������p๕�����΋Ƀ��Yv�9ГQ5;&w���-��[xD֝Ǥj��HP���Kvъ�]ݭ�Y/
붐x��e-[���F5k
���K9i�A�p��N`ƨ��wT.ʾ'�Z;�1�4ۼ�)C��j�Dg*�csZe:/���%ow^�ԩ�S�:vF�f�,�n7�J��%�S�D�'����
ͷ���7�%o�����H��7���YB��t19�g;�9f\/{Bu9ٰ\��8��6u��"��{�6�μ9�u�un� �DS
<�M�0���%l��qaA=wgl��`�TGr�;�q��ՕX2a��T�q��|���q�,�	�Ȅa��ٍ�}��D��bp�&v�:�R;�R^<�g��U����	���-��Š�)X'bgc#F�\H�1��
���E�b|e�*��Tp��J��ak9��^Mum��1c�����c%AIIZ3gjP]���A�Ż�m��9�|��ot���y!-F��I:�.����M�'�+�.�|/�qs{Ւd09RJmrŒ�y*
�Kk�*��`�B���{5x���;���N���{��j@�ފn�Q�Δ��ǫ[a�*y���fr�#
���'�G�y҅�H1�y�q������(�]/%7+��z5'T����ɻ�����v�����|��ls�K-����Q�[��HX�įT�vw)M���RP�w;h'���cF�M���d�2�
���6��Kk�i;�xgy�⛤�̛��z��i��J�q��s�R�9���;ֱJ���X�$˃]	㾶�5��\o�3�=�&�F�щ�|w���3!�!X��I��㉺�f(�gK��:�a�
�6K��Q]Vq�L�7z����*���K1ɰ����Ԯ��;V��4� @�w3���s��nu�s<E=J���\j�L��S,bդ��]�Y�2�rH���Z��L^os�z�]���w�*N2���O7���+���h��Ք�Y���m<+�����q3������s�[h*n���׼�t��A���+{�v�p���+'3��a��:`�S��5�]���LݕQY޽�:2�joov��YW|fp̙d�e�m�scw�8a}m=���W�-M䤔ē��[6h�}|p>}����&��]EL=W��#��' �˝{W#�T+�&,gFG���=�1S��{�w�5B�7���zZ�j�鬏�c�8��-2�Z��rc�7�,ތ�Z�)f �Kke�q�(r�)��@��Uu��r��T�9����7E$ɱW�M̢ؾtr7�;2�b�6%X6�prK���W��q��c�0�j�v�d��Æ��*�ٴ�����9R�X��W>��ԅ�Rt]7��r��b;��_
!����z�ȩ
��J��*����[��{�f]�[�����u���rq0�)�F0�R΅���*S��fX�k�h�}��Z�G$Ń���r�G�[ w���zl:7�Y�{���h��ow�k��bsnEYsUG�T�/��.�u�c�l�PV-t�);pi�YheEAiC���w�C����Rfp�8P���w׼��C�ۮ�yN6��wU�j�,�d�Gx�͸)����W:�D�P�3��9&C�%\\����.�5�en)K��6�V]�cu�Ɏ��m�clf5a_Kh)N�r��>ֹ ���p ��-rޕn�����LG��P������a�Arյ�\�Z��V2�������g0�SLy�vy�*er�'�x��My�V�j����+Eo�/XǏ5�ֶ�7/k�0P�&`\���4�A�[����-5ϵ^���rs3)�ٔf�6q�p��9ڂ���G�+��vzF��w�摽�z�S�Z��^�b�)����VJ1��{+u�I�w�U)���������;6y;HN���|yǅ s{U��b��H������{�osNSKq�FSkHY���W����ٍ$�;-�ɩD���N���J;�.�<��K6<=�TÚ��pӭ�&��q�Y�(�r�7r�����Eg�
I��\>�Ne��Ի�naw�Th$󨻹�/n�l��|�^�f"z��y|��z��M�L�~� eVG8��x���g'}��Ґ�A%d�l�������{��`��شw�_Mו5T9�=u���f�wm��
ˑ�#R���/*��=�a�C)��eQ�p����[�չR#��{Z�[���7\6e�����MJ[���8������E:��\B���tŧj�5H�©�Y(Ls��/u$��fᗛv�滫{;����)��g^&8�Q����������i������g���Wni�ݺ.�q�6���ڣ�B��So�e1g3-d�ͳ:ɳ��U͠��sၙ�&L�_(��P���U+F�3yv_7K�r�x��w�gW ����^P�K���kcwVE[7"��qv�����OOw��{�uL�4�NM���<.e�n¨hv�o:���_�/4f� �ۈ8��kfij>�ۏi�����69�0��e���>7-eq+����u�V���L�`����]w� P�_E6���K�dsN�5S��!���C3���1s�=�:����NpN�d��3�V��^3}��e�]���Y{bu��o��T��4�c{隦f����sJ�u�DN����r����V�3�]��oTȚ]C[�)*���fn�vM˓4Ή��w$�yN��A�{IV���S��9��ݷ\&r;1��V��{IK]aF�l�եd��L�Q.��u㱇�ڵ:�Nb�Z��V�Ԛ�5�fGʮub,w8�/v5[�m�Cs�[�iV���B.��݁Չ)gp��M��؂҃T��՗{��V���+h�y2���0+G�����x�=\#�W���-/973�_�n�ۢ�j�`�t芦ũ�Y*bRe�7�yҜ�4ު��[����t{13X�˨l�40������3*ҧ�Sː_i�ӛ��(�4����Nt�լ�t��aV�B�-731���_�W���������/��W�)��>�W��_�����@�u)�鯨Aj����&H�pE	�JW�S
j"( oⓎ5?��l��k�K(R�E� (:6�Q�D���%@�ȳA�̅��B�2�m�I9"0Q�_���V��vl��t���pi����pn�ŝbe]��ok]�L��oe���=A��b�f-K%k]զ�����]�l�Z�9�Y�`9MR�u٠��*��d$������kTzC�0����i�͗v�.�mZ{ױ_^�,�]�pX�x���ۚǖ�Q/U�~ݠ��B���;N<9�l���9���˦x���h��=�wrڪV¾x��mS|������
�{��i�M��=�g>)Y�J����a�ɏr^�5�bλF��%jA�K{x��סH�Θf����V��y6����RΜ��Ղ�Ewm����.U#��+��VR��^�szQ�XVt�k���eVӃ�3��PT���w��K[\�m�Kj.���%:��v;�4�VJ�c�t��g^ӎA!�����n��C�շب\��&.�CO.��!\�n���%����ֲ�6j��~�˃��ې) uhё�un�q�ܷ�3Gb���{֩����ڭ�-�;����.Ы���-nv`�qQ�muQ���"������e�.pt�շf,��z�뙗�1����X�Z�p�ݮk��7��� �rhZ��u��Ԩ/Öe����!�r�C�ӷ���Ր�P)��sF��U\`���9�y�z���Dj06P����2ʈ$��H��"ZnD��#!D�4t���������9

D��-��)E> �!p�����/`B�)Ӫ���
Q�1��8WѸK��n!�r�AM+��_�����b7	�aa�R�*,(�R܂$�E��`'rB��I����'�����@�'	��Ɉ�$(FʉC���u��u��UE%SA5QED�RIDTD����DQUD�������}��o������x�&���&�������"妪nX$�j"`��)��&����x�����}��o��ǃ��@DEDDLQ4�K5EAU��0D�;:���먂�*`��)*����UTm���+�h*j(
�b�����i�d��"����d������*")�ᩪ)�(�b�����1DP�QLURQQPQATE%Q3/�ETUU,�QDET�%PQ$TIUEqMm@LDI}x��UTk�i�u�F؜cZמ����-j���#WUET�h���KlF�Π������ֱ��h�Hj֠�ز�֚4d��jlڬ*�N*'[lF�Hխ��ڴD�F&��%�b*M#�X�F&���c�[���ڱ�z�D�!kuuѫ0��i��f����^::�+�m���:5��"�6��m�m�"���|;��f�Y�u-�I�Q[��;!�;>ͱ�n\��xwe\T�����Kn�<��ses��o�Y�f�i�qb�i�Ր�-i8?FA���h�K)@�P��|���[{�{�ʙ�+fIZ�Vִ5����L�����
�v[_9'�6��e���햮��)x�%}頿�E���T�����{���~kv4���J��_�3{�V���ú��fܷ�.x^�}�V�E;��	2�i����n�^7���$^�E���5x� [��������w�oI�|�I�5���65�d�����2������/Ax~A������ռ^BV��
vJ�c�/��Y]����sl>�Ƀɗ�<�-����c��y��S\����<I9��W�#���������+���W�
��DZ~3��W��Rs�~[�O8po���y��;(�x(����8���gck�l��@}A��I3��S}�;$~[=&���`M���-��ۗjN�p>�	T~~$*>P^����{�/ޞ�~�O׶D���N[j���D�Ğ>�����ǖ}��^{�������qmd�m�\�+��-�pML>����X�/S����u�/'<�㗹�ty��vDHrv����u��V�mCv}�Xl�E�]0��V&~����[g��s[:^*Վ�>c�KƝ��z<����
����P���w�<�����}xmt{�:\��ø%�]����h6�χA����\���|c����O۳����R���>����3B8��l��9��/��H�kL:�s�»��9�;�7c�Ay���{�ឝ(Y�]�W�����+=;H��hI�et���I]�n&6k.<�2��7}<{@��^xc�7n
�������J橁��_��Ɉ7��<A����4\�����x��X}RW��]ٹ�`ޢǺ�ڐo�j~g�~��g��]���
�6G8	�{���<j�.�m1�M[8;#�y����7�z��b
kU���I��#�2�+��'�^�+���ׂ�O�:"m�}��ݾ�	֝��o��:Ǣyh��	���C�����m��Ժ����������.K�g��f��	a���:����Q�ے��Ѭ��2м��6�bY�9���L�{�P���>�/�da54�1��{P�<3���ƚ�UU->���=���Ÿt�ݥ\���YW.G;9�R��'��g�Y�0>,��x�V��C'dئt_u�P�����>��<�����}�T�3����O8[xvl|���C�����+��@���o֞=�����(pO7Dy���������C|���Vhy*#�?��<�}v���6i�wD�φՊgd�F��.���{��b?L�Ŵ�����!z`��T�l����*�V�[tK�T��D�
i�Q�ێ;=4T��1(�9�����ӣ�֕���N2��{Ẏ�/ޛ���_H���1�'}������LdeH��ᤵ�)��0��m��T����ܸ$H́��3�7ׇ�N���ˡ���J�p%z��M���G#���8�����=���n,����xc��:����K8�b�Tz������Y$eq���z�2���+K�oӰ{ᱪϻ�;�(#��|m�����vS�?Gv+�h��Ƥz~�n�LQ^}�ni�J%�yEyo�ʒ+i*�Zq���*��rb��D97+:��2�w�dO���\^�9\/i���O8=�C�x!���ud�ܥ\'������Ow����X[��u�qn��KVΝhE�D�#��;�|����E)ܝ�>�f�� ���LL�\��<���L���@h�ı&��Ά��]����E����G��֙$��zNM_�M9�V���*qڢ��j��َ��?:���X� �5��rI��3��ѣ<j�*6��E����9fw��^�h}f1f^ ��x'�����ү�yɔ�����S�r�^���w~�_xA����zϻ�r��t�=������31xgm�?Y��!��Eo~_N�0/�W��o>�����=���|�Is�H�����:�zv�`�������L����o
����	y�k�l;�{l�g�cq���=Gt�	9ss�9���	����̛�&���\���|��g���Ⱦ�p39�G�A�7o�ǖ�=���kܢ�z�u���|��Cv��Y�>�'����� r�G�����P�va�C��]q��O�]�z�J0�f��q<�W�d�xz�zS����yom����%���3����k�ެ
-i��8����{.�7Aѓ����r�W,��R���uFm��O���jWta����3Z�/��orSt� ԯ��9��V�ݗq�[�^�D�o�Y��}�Ȭ�C����+�+>Ȅ���O1N
�j���K3}h������+� ��N�_@�ݕ���=;�eۿ�Z�v����9�<�,H�C=���^���H��vd�UI�4f*j_��5�{���D׾�h^k����������O�<�h1qB{bg��'�ws����z����`��_d�OW�֟f��*a�FB*��/������3j_A��C֖ǎY�|��m�sI<o�����������2��e�v�>[E���>�����rs�ǺIy���q�q��Kw=�w���/7���'�; x(A��N�����t�=k\�1����es8���m\M���y��2vک��/"G�G���;�./za�ڷ���G}�r<����xobO��*{���e�eS�/��T�=%>�Pb��-x����ncҰgw������[4�l�iod۶GO[�H]V�8-��p{� ]�N+K+�34ek�flm֌��=�h+�԰H��bJ���Ԕ��k:�hVKy��9d`bD��]W��ӑ�˘�-�n�E�d�1uZݐ�h���|�\Ps?l�=W����ɓ�{�t��� �p�@0_=�ۏ���Z]��qp��`��~�<rܙ�ν�=���g�Ͻ�]��y睞�jK�
ؤ��!��&�<+��ɓ�jo��D��G��{�u�1�}�!|�Y��3��^ݩ>����9����������W������&.ɗ�)o�Z�"��EF1�G����mt�s���T��a���ͻ�'���E����9w�C&����>��G�0�TI܋5F�MT���W�ǲ�P������� ���8^ϰ�߄��E-���2��3�ʺ����+{w���_����;�g���a��)�\uCP�#�{�ꉍ�ˏ$e�����A��=��!'�|��x��k�O����hwC�l�fɡ�3x�x��h�������)n�^�[�MclJҢ�fL�,����	��N�P����p��c=�Y��>�]��hg\$u��'n�}���c���2j㏫(ns��9J0�$p��cܰmfi��v�a�*�vI�a�'���&RͿ:�3)�&fF�o7����g7��ݿp��d�E|�a_��4g��=�z��r7�����c�ªO��n�Xĵ��v���k��g��񷱴 �j��sޔ}轓���+^
�>ϝ6��D^T�)�Jש��x/b[�<������ɝ��ȫ�B�ە#��Ej��yMC�*xX�����Ьjy'ʽU�ȝ4x�c�w�w�U��f���]tw1�f�n�`09r5��͝�7:a���P��LE^Uq�e�9�Ի�o�.�CA��WQ'�{�s.׋�Ž�֗N��3A���uj⸜��?M��e���_@�@�������Z�!ܗ����}�%�d�c�+��#�15b<��uzwc�g�zǽ�މ�}��Z�o=��ޚ<fg��-�2)��Uw�ף��m*g���7��Uwy>�J�e:W��YB�.�4������C�&ś|vУ�d�U9g^	qD������̃�pKU�{$l�����c��铓�c� ���(#��r�@h�]���:P՜(V]��>d4�um,y$�]-�r���nm�s:����^�E�7�Ϲ�cG"{�@��>:+���\�A�ܷ��7m�">^��&�U�U㊺���s�dT4X�Md�����t'��z��0���
�����y`F9+����MChźw6Ox��a��X�������הg�}n��(N�8{�{���3�L}Y[����Gk'-�a�g0��^�u����D��٥g�+�m�:Ep��G��i^B	�7iƱ�������I��Mx�L����K��D��fM�۽v}�*�(�}��돴V/ս��I�x=C��c��)��Ҳ,Y�n���6<�=IX���3���bpO�H�ׁ�$��<u��[���߶�I�w2ԟLr��
� �\~cï��>�k�
�Q��1���]#N���S��#����g�;+>�
t����K�d��,s�o���Y3�z\S.F�Һk'���y�*q���j,�Uz�7Jb�ky�RL��\��'[PVmK�fMY���2�E�0L����$��و'ûgf��L鋌7�ܮ�3��v76�)H����݅Yt��xj�}}׋n:a�Π�)����fl����Y�F�|�^IN�2ڭ���J�y�n֭A�O|�w�=�O=�{�?"�ͰE�#�׷�O��L{��y�|�9�N�x�/ݻ'��~��<�; ���hO�|+���ߍk�>��^���˝S}�Nb?s��v�����|s�\]j�ͷbe)�R7#�����`��X�^��sޚ<^v��-`[�x<تW(��w�J��N��mx
�y�+çɌEe�|ǽׇ>�%��m�s�ٖ���^�u���?l=x��ۤ��~��}�r�Ʃ��
9^��n��.���߆�y�"A�x�u���5����ݓ�=�	f��a���Ng&�7g��ʲD`��p�&�;�)�rhl[��kf������Z*�#�İi歍����T�'j��{.!=g����p=�X��R�}N��NCc�4G@w0rɠ2ce�����g����);۶E�EL���3��7)X��ݹׁe�Y3(�"K����8�oD��o\�C�_{M�;=LQ�~�&_>�q�^vz��z^��3��stKl�o��tЗ}H��G����f�/W�[�z�Ξ��A�!]�=QN=���}�l���a����JLJ(E�� V��;�\�G95�6n����M��Kogm[������e�M[@��$\�pzƱ��2e����^k��X�ښ�7 ��Ƀޞ�Z�V��$lA��3�VT��A�������7x��3ƴ��l������^|B5�xx"���U����8]�e��n�U�i�Ww�E�;ǧ�7���T�H�x�Y���YN�nv�����%�w=�[�:N�s���~s4o�Ͻ͇l'j���]�����{e�s�5� ���ͨ��^��4��ݦ�q�Ҫ�����>摙^���^"my��:�sH^�B��{���z-��Kќ.��<).���;�y�����N/�|Ģ���X<��S/J�]x�z�������(���9w��T�u�L/�H��4�K5SY2�U�Jvɇ�y8hZ��-L�V�ݱ��0=/�ƪ����=�KT�h�����3��5�.]ȕ��3��a��A���h�X{�:�nT���Ί�r9����T��V�ߐN�;�����4]�-�0����ɽ�o>��Eכ1s/��d��3F�Ǘ˼�̏(d����ا��Rk&a��U
��p{}���	vb���Xѵ�h�]�� j����]Y���+8U�pnE�{m�[�Y2��N�!������ȓO5�]���ׂl�=�6V�b\�Arh� �z�
+.�o/�I���XWV����Q�29v���ŗ%��j��l�Q���n��ێ�->�g7y��Yyp0�
�I�SB��J�z���Ka^w<�c�� V�N����l���wy)uث��왠Ѷ�����z:ڐ9��_�e;P.���6�S�I�#����/ANB��+�]jRj��ѡ���ԛ͑�����%f������;����	+�(��c��G{����e99�U�q	���4�}�SU�v�̎�ڔi�o+E��T]e:��Xhک�n��`7�(f��U��Ejŝ�$��h7�n�줐ڰ�_�J��\�$�ʣ�RX�7��
�4t͛|��匩�\�&�5g�����M���iB�哲��qN�\t7�p�\�	�)سvլޛ�� r��/s)ꗃu�[�Z��^�����Z/�ب1�r�8��y�*�ju�����t=�_T�}ꮾ�8Q�$J���9[�4S��!����wae��;\���}�/����DkR��Gx��X�Bu.�l�Օ�f�	=.Ll����9BQzxv�ܗ�-\���J��
�1��f����T�-5���B�V�u5�$VA:{����9˵bV����VLY%K���)�n`\�{&�8nK�̣���I(�I]�F ���fK̢n�Z���\�TA3�̋p	��{��ǩ���{��А$t7�1���ޑUBm}���Ce'D�;��Y����A��Q���E��ʚc�!�Dx2�Q2�������M��R;��J�����ǳ.]U�$�]k�n#�C ��%���d9�i{R��j��-:�R�9�'I�$Φ�z\Ǽj��Pg;ȸ-�vb�*fIK"�_�\���L�6�|��:�0X�6��z_d�2����%iGo����:�S��b�1.��������YCM��Y�<][K�S:�ccA�_Y'&*$X������x:v�\�$$�T+th�	��4�\�L����e
R�[�5���VՑ�����;�*�9�pIూ�E#u�����u[\c6���f]J!�7�`���%�n! ݕĂ7:v1	���ݹ�qg	u�܎ !��/��j���
�yե���A��\�^&�C/��(�H �]��U��lF��F����A��Zk�cU��Ϸ���������}��o����Ȉ��Z�W��E٘��J��'Q���E:tm�+N��������~=�������ߏ����Z��֍`��h��݊���M��3Ղb������� ����r�1Q1CA^z�%��1�PS@U��>@d�
hh+��`�� �i
M`�v�P�TQ#G�����(��EG�P��d�lbh������	����z�UIIMUU����DBUQQELIU0�M1,QE�i}mKAA�cEQP44�U54@TACQPU5EE�UUSJx��J�����מ�x��p�Q��n�V�-��U�E}���&fr	��͇��ɗat�9��nb]���";o���Y7$�|����>ӕ����FqP׸����psA����37���<'�����h}�Mv&�%�U��3���aT	�ݒ�����C��j�ǵ�z�4��iV0�`[�j�!A��`E^N'��с�� <���j��fA�}��3�Z��<�Bi���10=���΍i�L�ge4�q�`$�b���f�StL�4_�����1���޽{���%��8�,:/1>��u�U[x%cj+ӼD���-��/!�/9�~Z7��3�����k�֏5|���Ui��l�Y�~c �� l{��i�	Q����O<�EWY�i��YC\W�w��7���4��Mn�om��[:zkw�H01<fͱMP�����H�#��c�Ą;!s�DIt�g�
N�@��]%��m�5c\:��ONwE}-�o�б�$Y[�ޮ���5��u[!���0Ct�K0S��0�}�F�p��)y�sxsQ��E�n�{V6�m�Q����C���ϧ����>�"���^�jOxT�M�LC�zOȆR	w�4�14�!�o��q�BԁL$�XE�>O�`C�G8���N��u�9V�~0��ف��S��s��a�:�[�*����FDo��N':슈-��,ޢ�#Iqf桲*���T05�V��u�=ݚ� �2��)��^g^��k�f�=��bl3�6��L���yv�"�,�S3:�����F^��Ef�xJ��ޏ��hv6y�_7���\�3.H����sד㿇A�<��>?��H�.�[�˽BH�uS�)�*���K�%�n[����`��w��<ɏX53��f;����.��3�%�'~{�~Tg.B7����f�7y>��G0�ƲǴz~�����=��H���/B���A2�{��c�l.#��C��.��}z��7:RpH	��
$@�q�KsP/�ܵ��s�'����g��s;;y��Bt���j�	Vuל8hM3Eډ�`I1���Z�Zi:淈OT��ᛦ~c
�/֥���@I��^�� ���7�^�)��#�u�mN3d]��q"&LH�GY#�y�3Pd,���`��-���������H?���V�����"	�wV�F~�%����ߓ|'yo9��O�fF�-I\�j�z͐/^��t��oN��7�����>[���9�H��N�����.�C�� �QX�W(!?5� �c�bWN0Lu�5ew�%���  ����̎�L\�7ѷ�P��qK�]��`��z!Z��N�-�+�ʩ7��[<�5�M���=_��mߕ�/�*h\��7ܞX4����/��An��
&�j[t���K��Yo�h�[��
�=R�"�[�Y��r �"B=lW]B��ɹ��3�A�Y{���VuG:=N����n`]�fu��׉�r��g .�mhu3�qO ������Ƞ�J��ϗ�-�8� �Z���
#��ϞV&�d�]	�N�s�v"��b�ߘ��D�7�R�j�QN|�'�v�C��&��/H�K�x/UŴ*���	1���0v!����;�i�0��L�qx	�4�y�8��J=먓8�Y�.G��tvP.�����H]�  ���pO�0�}YP�4��t�o=Ĳ�Xa���'r�K��!����;fط�,�~�e��n��s�s?>�a҃�����K���'m�&�	ۛ��S�W!�%�z�u���W<��W�\��`�,i�`���������w�1�co;�S��4�mod��a��Լ� О��ĜqvJ���k�e7�UZ�|���|�2�5웷��C���Ŝ,[������i�� ���NK�J�a �	���Mf�x�9,���T?Z$n��h�n��` c�D����&��j�rT�'�{F���;�rr��*���z�kC�y�S[,�ʼ�~��'�n�	a1��!���@u��d�Vl�l�e�!��0DD���!v�r<�e=۳f?tD2��a�z�ų�sK��p&tFa�>0���G�6-ٓ�V�et��w^[���_��ʁ�,���u���l؜]A�7N�&�:)���͖�p=�G��e�gwu0���/�w�Q��n�4�1Q\**X�$���ؑ�8ݺ뾐�H���m)uZ�l���K�m
aov7}�h���R�,twu��y��9Qǭߍ1#�����f8[�	@�za��Dl�tM�1�63�0%��`�X+�Uө
�C�����Z{k����3Km��I\�)^iަM�����DR�q���V���\��{���=3N���.�%>z�1��ʩkj���`�� ʂˡF�Ty���l3V�w;�����=r���3ǉf[Z�L&�^�^}�˯j���?)��O�d��'Z[���@ˋ`�Ҿn���d=�*F���z��ᦞ��8(��'_+�		���ا��L���-�����7'x��N,�LPR��ɶ�5k�<'��x)�:O�l�'��v�.��̼͛|\��G�����m�ok�Y'Y�ƒ4�P}�/�P{���=��3d��������5rzZ�u�sXc>� �w�ì1I�U(��x���9�Ϋ��� ��Q,M��H�'�/�q���#�-ٹ�	��e"�У�S���S��֢��YPXחI�������-��#)%'w�f?��#�9`9���옔ꧤ��j�r����ը�s/�M�ϯ��U�J�%3�񻳍��m����V曎��� ��U2��S��|��CR��,�3C�&=~Ē����=��c�5c2tٷ-S�yqU�+�����9���RV��5Ò��	E�h\��P�-?LXi�/w�W�����o\�\��C�5��D�1��=�9���Ǡ8u����تv�\���pkXt� -z�|S1z«����gd���}�����z`��'O���d.�<9��|~�_�h��Y�
?���4�<R�,�|�܇��bړlm>X�#銇y�{j��Q��`�8y����p#�#�/:"�L��7��Ook�l��f�*�C�_7�'��zK�"� �yO�ϴ@,��Xh�q.���3{(��v�P��l>^��#�L��p�"vR{��t����ӛ8�F�"�H��>'�	�[�]��S%82 !�e5I��л�v`��ŕ�a�á#��MC�ʄ�^=�s���͛�Y��)]ȹ�X�>�
+F�S�A��<��{*���@_����>�����/\�>��^�%@3m��̳תGjn�4'��g������7�5v�^͛/X�o�U�-�p8ƌ��PU�+Q^W����ש��i�e�{x���������i=����^��-逷}(#5�M0ʈ�wk&���¾��{`�s���Cg�5Bq��p8��\�I��m�s�l�����$M��,�Ph{�f�İ�k��i��-����`G95��!�OA���z=ݒ���V3���������f��������myb>��}��W]R�[��%6s���3��������}���W���S٘ܢ���y$�^7���Ч�-d=-6����_X��$vJ箈��$�D�Z�K(�`-�6�
�p�U���c1˭�]z���:<1�Dx�3m��H����A���4�ሤ�sG����s:�j�9m�c]�{PtoCqn�0vf�&���=̍�0���[����X;/g��(v���u�-?-�
�� ^��U����\_��� �Q{�]�������G!g�����G�g~�6g ��V��\CER�=�e�z�G0]�ܿHv���Jhϼ����Bs�2~15�im��xR�2{*��CĸQ�o�t̢�،y4�Ъdf�;�n�yÐ����x�i*����Vٗa^^�(zm���B]���hZ��K�1������	5�>/���!۵�7)k�^�mvٹ[|G�6��̚a�f�K�|�R#w�ԓ�	��C��/:��nY_�׊�c)�®ۥ�C����� `��ЇAi0��?�2]�A���r�6
�N�R�Y��+ϼe��{]9آ+�Z<�h����yW�%��36�[�<:N��\��>�y}Bq+�|t�/β�ڋ?]prRR;�o,�ax�����l7���y��������Ʃi4�bǔ)��B�-c4�uR�MCD3��Q����օ�'\[E�Eo-n���;�0�Ņ��Wh)W|f��J���FY/��젥3Y�$zk�'��G��{�����Q���1TS������� ��w3N0Z��H�B�k��Ӻ��6u�5fE�����KO���I1��I�<!�vy\��
�_�צ�ʙ�|��3P���+��*��`�ṭ,��R�g�ٶU��Y�P���ނq{��SҶ�#U����	�y�Y";z�ֈ{`�N�����B~ka���(�3鎷Ƭ��sn��H��Q�X���љ���P��F��DzT>@� uC&��\�:!��bыN�-��*��ۜh+4"b���'�B-�x��r��5�$Ao@
���JN�t�X�/�75{�$�b%9��XJJ��9d�N\F�({�θ����M�8މ1��,C��@��n>��ޕ)�z��oa�/�W��F���=�ĵjǑ\�O�8]�)�ی!�By�s��w��e�_6��|�ݴ�/�zͿ�:�9�iɍ݊@��"賎e��0�vk���͓�=h@\�!�b^�/����c�|Q�6vN�!�X>c�mP�~ΤB��W(�ߊ��=h��	O��|y����7���6̵���{Kr���K�:�<hY/�V����] s)�J������Ww�����{�x����+�a�W��{j;��Q�]����u��y�����LޭY�x��<���{���2y)u
�n��k4C�1��T�Id6u�So��<�q�j�uUMf��%�77���.�R0q���!��|$�K]k����?�����}��\.Y�T����f�h�T:ni��XИ�7���0m���_�k�+�%���*9�b|(��.m�����ù����0vC�Z��9�0̲oh�֡��i�k�]N{hI�O���t�Cǝ�y�-@�NZ�9�dK����!0g}����2N�ٲ�R5���n\�Ě}�t!���nD�)ٻG�` ��g��Y^ZZ_��y�����a��òc<m;97h{�� 7i�E�Yyލ�"ʀ�#��XE��:&����l�=�5�0�5�f9�����nvQj/��lkM�q-^��9�+��z�po�C#m�W�b����kSN�`�h��ʸ���d{ZY�=�CC��b�h��U��2�Zڼ�H\�]J�D�Q��?��SƯ��8O�����g(e����?����բ`�ܰ�%�*�nV6�[���M�=��A2��Ge�O0�ij6��c��������	��.�t�U��3)YE��b�|�I|�&B�|Cu����y���*��H��M��'���J`�BR)�*�u��(z� w�m�h��hL9�y<X~�YJ�;8��n���j2���3��=H��%sQIMkyo]�� y��n��5Ä���z�.�]�ǶR�����!�+���V͸w�we��Xֳ<frs��صED��ya[�Vt���P1|f�"h-ӧ�n;|���}����fq۽�c���������� ���=l�)��{�|���Ҕ�N��,���b��Ã�_8����~���@�ۥ�g�ʔ���<�x|�ʈ������D��Hy�E��R���s̱[��u9jw���&��i��wU�b��li��p����y���&���^�����Ich���in���V�uS�u�7R�e�y@`嵤B��1)�OIib�-j]�wWQ��Q��k����{Jێ����X8�~���T�cq�<����A~?i��Bm�V ��0�*UF�Ϊ
w��q���9�򸮿>>����t�N���a@"8��v�M*a��]�:+)�D桷]�1�*9Qcl���z-�1�팟yP(���	C��Lh���p���Z0���=m�����#�!����Y�����ϰ�b�:�;xw}ø�����Dv!�l���'f�e=�/x�oN4vl�xCp�C�"���[�b��β�KnP��ܛ���f�험��g��->C ���'�OE��g�i�nf��E�WRQP�Pq�4��]7?uĮ�;��2��b@ͺ�v��%�H~��'$��氹�;�eeH������^<�����I��Z�˺H��2�����F��'3�����2_Ԧ u�vG \�-	Qе�1����%�۵0X h��C�����c�Q��Һ����}{����dC��8P�r�Ӷ��Q+D<K�8z��|h���^Y��	i!Bi������y��=,�%L�b���'oUf�S�S��{��jW��5�����I���P�H�x�K0�ma�s���j1�U�4�x{��
��wZӝ�]�i1���`�6��j�V'�+2_��Ui�P�R�~��	���S��<�"���u��ad:}!
*��tA	�Q,���Y(�kw�{l�uފ��;Ʃ�eP r�Tm_!���I٦��a��d})�|"S�P%�i5��۞k��ցK�-�囮��#�ix�+���j
�m�1���_KW�*2a����$�b)9Y����ՊF��=.�.�8P�qq����?�C��1�lLpm�{<�_��S}�-���1%��t�B�u����=����d?��݁��s��7�d�d~�~z`kÐ�3�U	�(����zu��Y�����(Ɨ��ct=q����C��$X���t��r�˽v��]du�mB��T	mQʭ�����FM��)򨁗�wf���x4{���v�J��UB�2S<տf���P`W"�P��	��z���n"��f����1 �9Ȇ���k��À���&Ua���=i]�H�4�7)�rƱo���v�=���3%��ۉ8�/
����7q�C��N�u�2 �;��mt���
ً�L�k�>��i�*�ئu�f�Ӎ:���kѬ���JZ6J��Y�Ϻ�Bhq3'IsnGD:ܚnݗR�R���[�LG��.>�(]���E2DR�L�Ă��5S{�ۑ=�.$��s��Q5��g}vm�9��F�U����0��i�BMed�9q�.Kw��9���v]�vԒ]��أg�ۡl�2���&m��(��o�i���\���쮽r��űtު.��PӸ��ˉʹ#+B˱
Q����3@D̆�`37�	wU��蔺�V]�#w�b�p�:�h�zd�`�h.�9H#VUlCk���oU-sL蹦tv��%���WPCϺ ��5;�dyp�Gf�$�'��hwp�b�����������%;���`�َp�h��Z=�X��o_]e���KSX�q���,;[mKQ�������n>���5���$����:��[�d\�$�+Gn��Pc��c;��n˕d��|��\��MVx\�Z$�
lB	��	|�q*��Yx���e]�2sV��{r�؎	B�͗�����\����m�Y�Cij�$�"7.���j��=��.Z�[Օ�6�S	l0Җ�ۃ���Y���;��a�:,zwN�k3	w�m����A���'_LU��IQ���z�M��%���2��[�)V�w�I�:!���vQN���͌��*�\�����rү5��JqPt)UC�.��6k�k���n@FCfwd��ÿ+��h���F�B�([E�n3̌�7Y��u�ڮ�;_e䦅S��vծ���e��m�c2c���n�r�^3��`��J�b���%��{-T�v�ڌ�ͬKv��v���H��/m�ud�t]��1��ڭ�r`�Q���{I��Ek�CS���uc <2D�-3F���9m��e<�n����F.�4���.<6n�l�З���S�;'d`��턂��1v��c�V�4�7zf5���gL��ӹ�W1�H��\)���Ws��Қ���2���R�a�z���i�3��OU:jK��U�Xɖ�Q�Mj��-H���j�YHԔr;�[o�-{n]{�Qp�r�����K��������H>w��7�2���E)�[؟iMNw��;'9�>�E��u<�c7Va!D<o�uJ���v��pb���bj��e�;k�ҍ�	��Z��ޱܯ%�j��?4�뛥<��LW-q��K�L�nu��&U����H��v���w]e�sI���ϗ�;�M��
"�*��i������(��"����B����i��x�~=����������?�r�(������X����4S��ꈙ�(f������|���������������g�*=�QRU4{�D�<�E4V��"J��b"���)�*���*)��MR�RU[�����)���������&ez�TPS;& �h��jd�((**�đ%CUW��:��II���\ڒ**��(((h/;QRRtiӭUx�4�4�]I���EDM:�Qs�����1tlR�P�ABQSD�L:�x؊
��P�QKQA������EՏ�V���� ����&��THTE��Ժ�"J&.��W[I�4��i)i(�J������"�*B�+��E�- � ���o-4�)�̅ �!Q$@�j�)?��R�K��=,�c�^+9̾X7-*_A��I��ʻ$=��3�%���%Ӽ֟L��-\���`��$�[ �
@�c(cQ��YP�J��
`�����ǂ:<A��Ꮆ|k�E~�������UU�{��韀{�g�1�ٌ%~��v��ٵ�<3s���P�nd��c��Np�\�%�u����:�@%��ًlM�����r6�Ö��.��E��)8%9�aB�;���Q����=��_&��ux�c�l��;���G3�{��"�R��Ld�d>���Bk��v��@�S��9tE��]��YWGC���������{A�4{E�3ä�=1���s��⯊#(Ry��5'KPg��Ṑ��:�
-�dz!��ִ�9��l�w�Ϲ0�a:¼��;�,�=];w�U
kg����ۛ��V�kNr��A�fnj	\��Q�g�ٶU�-�<�zw�\g ֵOC�Kq7�w�)��!1����1Xʊơ+�I��]r���kY��=�eEÐ��[����c�n�A�I&=(
�NҺv\�c�{�A�����T)_���
n�2Ǎ^��YF�	�׽�&V2ʌ�ʸ�x�ހaH���N�/e��?Bnm��9w��ۦ�ܲ/��1٨]U�ž�0�zh\:q� �5�z�e�WK6Ʀ]k��ϧ�����ճ��~�!7AZ�ש�W��|uU(9Wi#�jo���S�%N�ܵ1f;��ՍԻ�d	50wf��uҴ:�ɮ�@LݮQR�n��پk���!��R��e	�e�'�C����t��We����"?g�(�s�O������o�ߏ������� �\�$��.��8^����xa���b�'�pE>�<Ԍ���.�{;�+3���^'6��ܶ���,㛂��6�vk�����\=� �k�I|l`��&�_vs�o-��^K��hQ�0�aTJ疡j��*KGi�?&�v5�����d
�2}������ͭh�X���u�xв^���*�
�y��*�^����Z����ץ����8u.7y��<��	��9�s��d㎰ǥk�*	{n�f{�":�fauڟ�Mtv�aW"/��� @�38Cc�D���f^�a�@g%@�uf<A�0�Ls�L��<v�,�]��4��<�KsQ膲�3�2%��D&�^��s�a�ӡPՏ��ڋ���7f�p�N�h�0C�Ir]����C�-��l��^]�."�FGp_���ȿvwE�窈Q���DG��~R���z@A��i��˞)�{`3wm�7f2\�W{�4��B�s�'vi=���{k�x�{�D<�_A���B����������SA'H��U���%��r������9����×[�m��7l[��*Tϒ��UV������/3��u����I����Y+���h���u�LC#�ŕ[�aC��X�Tz��w.t�����������Fj�YR�V��h,��7�<�?��|� |>��������y���P�!�����xG0�ܜ=TIx�S�5vL�Sg�)�2�2�2+2���O+���Mo_c��b�Y��۲Ȃ㦽�p��`h>_���R������hQ��˼5��9�7�����A5W�۔.��(��)QE�s�����
��l�|b�W�[2�i�Y;woe��F��1)͎2�&��*`D�
�{^��=|w�!Ŵ��,��a�HMn�h��{4j�� f�f��N�����: B,�ʗI`���{��������ch�G*��Y��	Lн�=K���@���]�_EL/�J.�s�1[��&y�p[0��&�.�ѐ��9وg�!;�m\3kH�[�L�7ƅi;��*���������s�}�����n��E.�t�=�}TCH��-�?���tϟ��9���O0-�܊�*�;i�bz��<�+v4\ި��U�:��zp����:����ֿP���ZYq*�Z��5�f�谲��gr,���t���r(�k�tͶ<!t�` ��~��:��(�����,/�����Y���;�ʹ����Gp��	U���J��	V�h�
ב����D%DAt��ݗC�l!��4z�D@kwQ}�w�u��fiC�����G;UX��N�]�����xN� 6n�3@�U�ǒ-r��Xil�p��p������� ��p��A�j;�BZ�����y X�����eK?x������>�Q�s��y���QVUڭ���,��{g�K�;�*�P��Sܻ'm�yA�$�%��Ǥ�/�;lq��ވ�-]b:��S�i�X��ݎ�5ZY�vd��C3��CC�'(���:[��f�0�~�$9!�OT4��u�tV5аq55�HX$�z��ʢ*k��"K�Yڙ'�z��c�XSj�zg�L���_��/�}O���G�F�vA��w��^�u�r���id��FFS���>��gL5n01U'r+&�'V�Bf՚ޞ��d�����6����@�{[@���ǧ�w﷔�Q�
���g���\�Q�0t������9J���M'�t�
�au�|\8J����&���޼���y��2��q�wl�+%W7;��o(�E���_�Mw����t���e�n�.�Ƿ�ބ���tp4���wʘ,�	O�$�׺"S����:�[�&�����Kh�������e縸uC���i����`�龖`� Ì�uI��Rr���Q�}�����q</�Ȇ�ƛ6��]�f-�	������E���G�cq�@���f���E�\�¶h�wV� ��!�eh�h�C�.A_^�#�C��;�1��:�$Z3�s%�*��]�謫]O�*�afam���9S��^jԅNǄ�!GW���?N9�����__<w���>=�������bbS��� v��j�Ȳ�����[A���86��;�}¥��a�߭�W8h��Z���Z�н��匤�����f�p��"�kO����k��nGZ�ó�A�2�g���u�m�ֻe7�M���Q����,!�ڇF3�y�!�X�`�k�`�]k2�_2t�3)��)�	2)�Gu[]��+���jR���_O�*�C��ٶ}���v�te�ͮj���W�+(����wfN��6��T-1�û�cYc����3�p�0o78����¹�6�%{Ӻ��8N�.�����Ŧ[ץ�>M�Yԓ�`'3L(���q*�:���n~�o	ڿ1���CÃ�k�6�`PZDL,rޱ.1���A��ga�9u�Rfjg-�n�B�YN�2Y��$��9KO��J���c�Ϝ�/�#���+����%�-��l���j��^e	�oI�j�S��R&a��Z��E<�.�3Y��S�#Xb�h�XճKiNݶaC]:���έlNPq��2�sXJ�D�s�oN2�6��-.�(;Va�Es��I��	�<g��3�Ź�S��%,al\��N�_{:��*W�~�5��Ԩ�E{������ݑ���|�����S��D�b��ɜp�Kx썹�V��P26*��(tRm�S��u~�G�Z[�C�5�ʵݼH3gHwW� |>���� �� �9�e��ũ�~Kϡ��W�nB�ʯKcP]_�sf�A=����w��<?S�Uϑؔ�������&���C�3��.lD�Bby�B��MQ�B�#�Pe������D�j-�J��QE��[�Cmڋd9��?E��]/�����;_�u6��N���:!2Nf8WL>��������h�w�S��VVz�q����3"��oH/�b �@�!���Y�g�j�5���^El����n�U�լ��~�E��q�n:p�6S�?������OגL�^�1rՖ���j���W����
yF/�뜫x�K�ӑ:������툕�g�k�����5s�+9�>0d,���A����h��<��/sM&��o��b�E��),i�a)��vm�k)�OV�,Η��Wi��6�LY�&N�����uBxг`Ĝqv	�&,(Z��S*u��-����c+�YZ��Yz��?0`��:? Ť\����09�E�jÙ8�1�Z�.Վ������ƣ�����z?�פA��֛�.� A���O����Q���@�����e-�[挟�E��t_��%ǧ�������{o&e�WK����]�엵hVOh+��e`�w��vyI�#�:Y .��f�y�����ܡmk�������jDd��0�
rp�e�BJ�#2ږ���U۫]B�����}����Q�p"+z��Z��WϮ��=����ۗJ��D��Ft�{��+����=I�`�x�	�<F��PC;
[,�Geif���%z׵mc
ė �f�}�3t=1��_�����i
���k=_:ΐ��Cκ`��Ƿ6����y����� �醐tE��MD�)Ğg�N����9�3,g|"|�
�(��E��X͍i�Hyj��9�+��My��sύ��c��Yy4�e#c�Y1h�L��S��)~�h�+f��}���F��B�:�2�uL���υC�%�{9���w};�{z@��e�C�lS:���`�È琶1��mT�4���X�4�	̞�5���S���a�)�Wm�Ӻ��V����ց�iN$�{.�$)�M���ng5�t����
Β�)���%:*�)J��E[�e�'�p1��G^_��A.o�묳7�:?���!t/D$v*�锝xd�!��#)�y�/��a;:�G�p��}��f�e��}�z����Oy�_�ջȾ�.�X�R�����4���x��hAˌɫ�)���R����KU���零����S�ԕ�&h��;���(Ȩ
;�K@�� p�L�-��{]�t�X�JK�Ү�����cU;�J��!�e�E˨�x��O�ݺǗt�B��P�Vu�d�Sz�j/�7�s�7��}��U��A�|<]���٪e噃k��L�vlk�!7T�y�ugo6�ߠ[�=I�>��T�\��=E�\��eܭ���rń;�;�XG�̛Z���u��$��H,'X�'h]%��43�j�gy�;��fl�ʤ�r����AWc?������˨�5�������1�M��M-��6�x#�Z�9/R�Yu,�C��?OH`�à<���ێ��j�T�ƹ���������ϫ�m��Ĳ����>�z���,ƽ�p3���t���lȊ�n�h�w}�u�c7�B";�'�|�d�"�C�H��_��zK׉;x��<tE1cw���̜��O�p��TK�,( ��<(��%�)�j��������t��#���lqI��K��[v��B���b*VD���	���!�Z}��՗�)O��θ^�sް?%���1���Y>��l.��`\dÇ�/&���-35B��`�??�|��k�2���<E	�VZ+i���b6'�N2�^�3m��$_��[8����|آ�1��{�2U{(����}��%�϶SԀ�y&��#��E	�]Ѻ8֓Y���Q�V-1U�����J�f���H0�[�����ff�%��
�6��v�F�,��Ϩ%+���|�����⍝�Z��^��UU�gw���׾����nx��u��}���ȣ��Uz�ާ��NY�w����v�_l����Z���,3�/>�j��+Q^��%6�徤5����UӬ(�ǫz���o��n���˞2���ͩ�-,2� wW��\��q��Y�R�er�&�#q�_#!8O-PR���i���?�Y���k~)m��䅏"�C	��W������)�m���ZԊ�5j_v3����t������U�/��m���U=,�H�$wQ��&�����Q`���j�Gp�Yoz�dWW��0�b��|�>���A�{ �M�3<#c�K�Υ�:.՛��<�f�v^��m����������u ��	���*�M�>Om��s�'Y?2���w���vܙ���3M�3�k]��^jԍcS�?y>;�wv��vc�ŷ	Gu��vT���n7,���C�u���)�������'�FM�إ>�S#5�ݛr�30Q��_ ��7� 2C�:א!غ/BO���:�R�9�ë�cYc����MsY+Ge�@�;jt�X���
��A���r1k�ؔX�i|�/M��u$�1,2�A�c��֏�E�Jp�ua[�p�\͵������bvŹyx`٫x��-{�p� �)�K��F��x
xYHE��&ttq)+�Nl�
����T�9��ڻ�5�/�U�[��;�y���V����\�v&M��c��P���'�e�(����r�)��>}}w��>��>d+���R߀�騽�q������0(-"&9��^H|x��}����ͳw0�9�HJ���;Ŵ����y��I��P�yA�7}`,D�N{Sf�[؝�����֢��{>��4&�oR.�jq�gD�6�}kO^畑*��B��'7v)��I��?v�P�y�'��x��J�fִ�n�SPC"���o�_#�K�㘿�t�Ȓ>��U�q�ߚ*��	�~����?+�_}=�V2�!>�0��E�)����e�r}Cی���w�m�TK�T�C�8fH6"K��y.����M^���]��r�N�tշ���mk_�{3��M�;Zܘz*k�,���^?X�~~��?ߑ�^�Ԋ_O#��}��_�~5������KV:<�R�H���[�S�h]�� ϧ��A���A�c�M��ˌ<�W��7�y0��I�����(�%Ɓ�������w BF4H��W[��Ɔ��]����Ì����/�;_M�OR�d]g���-/#k�m�~'�Q��-�ߥ4���C<+v�Wf_:\�	<�3�!:᪜�=�V�ni�tܝŜ5KEQ��
�>�����0/qӣM7����mM��\���d3kWi �؞p�]�T�����Ė���׏v�yԄi�Ga�ƶ]�m-��Xa.�E�u]j���)�llR�[��f�&��+��AQ��#�{�2�w��1_��-0�:�(�g�u,ClR�a�WHn>��5�綉��%*Un��1��}ՖN�X�	����͍���(Ĥ�F�A�\��c��y�
�N��l�xݬf�V�;��3xed�䡱��w���<�^�v8a��/�G^��3i+.,�S�w�6vb���&>����=�V���2���]��W��2-D��j��Լ�ŭ81ΐ�m]���^�Z!Fx�D��LӃ�����n]K�ύqvL���G�w[g�;v��������n\���)�"���D8�ֵ�4��I���E���']C͹��tMTv1������Iv뼹٦�zs�[\,s�}b�d"uA�z���mHzu�uZ'4���/��,`g�[��J��,�oHn-�V]n���\È@�� U��N]�*lӓ���唶;�z�/�W�M��.+ V��M&�����9��%�"��Bi<��z|t��l�p�W�M�\kw�a���}���3uDlnSZ/rh��J�=��h��A�Vbg�;��/&CL0Zp!�]@&�z�m哸s���6���2Ną��c�W׎I���U�$���pJi�r����>�ӷ3�/�P4ޓ|d���u�Wz�X9o����GRzݻ�tŸ�e�wi�X4e��&vq�v�V�*m�6)��(pwP����v�;Oa�X�|��En-8X�/��KB^��Rs��}�B-ef��Ӎ̠��ϹFAا�%x�r����t�v��[�3M59T��^8G����-8�l��5���9��Q��3�I9���E82+S���^(�-��B��57,�6�3��[,2�������}��sJ���r܋�ӯ����1�tL7�,9¤3� �A�f��N�}��}�����V;u[�+�W�����l�[�E�8�����,B���9������n� �4��̭=�sz�Ք�SL��mt�_Y���Jc���ĩm
����JG$֎�p1��o& +)O�?�u2CǮ?��jK��z$���'p��}���ܮMLӇ�,`�d�J��n�vɢ��m�=S�t�ҙ���p�v�/b�,Z�3Y�pkҐ6�ͬ�!�*Rn݋�z������:�n�I�)ҕowAdd9M;5��R����v��{��N6U
w���S3i��jooi�$=B ���{VR��v��*Z��sxЙ8�O2��.ɭb䯐�W�%S(Ơ�j�w9CJ����\�<�������U$HUAUB�4�.�CƘ����7R�����{~=��=��������>CT�TR����b�X�)bJC��Գ���|�x�����������~?�--	BUSAO��4{)EM- P�4�)JĴå0l�T�4�%RDR���C�xʺN��DD�u!�hb��&���(
 КZ
F*A���^�t�D!0kJ��)�!i��@��褦�<lXt�ht�K��AEAE-UAM����]�@D#I��E�H�V���P]j�5�LK�+��yw����y�9q��X$�u��>���m�z�_C�%�;t�0w-��p�����Y���5w�Ql��׮�r�}?g s�Q{�������|���=0d[�`pu�:K����^��i0�%s�U��^o�IcA�a�\eS���I�-��m�P��r���ʼ��S�M��_�]
H�^�y�����Z��S:�`�V��nMEdf�tw`��:5�h'�P�Z{㧍������r�BՇ2q�ӭo��L�M������
�s�G�
_����z1ֈx!+�#����B�sBy��oer�b�6v�휣���d/��StM��f��0��z��^�9�"]�p0C�wv۶����\��T�֝���Yo�L3�l�nvO{�����2{U��hv}@sQ}hwE:�~`� �R��t�t%Z(Os�J}`���w�i�@��/47��PiG�A��j��sO�:���\/1L�5!p�FǄ��\g�2R{��^=���֑yH�k�AzF�!�%H����`�;��yVd"�}_�Z���혾��P?�U�I��.�ت�j�ʩkj���{*��T�5��vS�o+j�(Vߒ��*ޖE���tR�������E����<�4
�4�d�SÉzB;�͘t9��u�/U9���6��t,�3G��L�k����p��'���vq��Ý��pifns�r]@����aNۉ*����kr���E�׸��󠎲R�n@�J���#{2��Իv�v+|���Qµ����x������~�u��_o��C9�*^�|��y���̳�ko��D�ky�8����'�rEh];�C��v�;;UɄ'ʠ����؋tYot��,������]Jd�u��LPR��FM��m�'�|wW�結�yf�c��j�w�vx�!�> �B`h�_2��}~�5*��/�:�s�1������s���98�ބ#b%��:����H0͒"��r��Y��.���酎U(���ƕ�l�B��|j���g��PPi��;�ׇzh࡛Dp��vz�Уc'qUeWC�O6��%���k�o�m7u��{k� 7.�na��8�s�m�{�ɵ�8F�C�u�������*s-]]\�Ӭ��{�+Q���s7�T;�`9��8~�*��a�Tz�Z�+s'0���kVLe�l�j��7zmB9V��L�r��U�~|}q������Wa<C{'�.��+,�9Z�x����C�:i�f6���6��&6�:�9G�ߋ�v���1a�v/2C6�g^���5�[}ڃw���^a��d����}{(�{����D�o�7Z�B�;ᬓ��*���Y}���;�G_�K[l�����j�*mz׽�NG�ν�O\�\���]��5�E��&�ڐܭ@3������^f�W�+��SP���c��v�K��F�7��z�l��4�0\nK`c�cl�]��:6+��o2�p8��磇���w���E� |?g9�TP f�z�ͫOQ��t�2���f,\��Ic�?�`h��ix�f�!琨�8^��+��f�0��tC�6gD����C^�]�	Wu_����b�n��}�ǃ���6~Y�Uj����Č�Ad�v٬����oJf�/'XJ�!@#&<�ͧ�9��u�,G4�	�ddcz���� �r�ګ�g�[��q��dcN��V��PcK&�x���m���)?��K�,�f�U�(�|��#��S΄\zx���j+ӼD��P�&!b�OaWN�<�o��"�例�nUE��,�w���b��Fqj�K�
!v�#!O6�L��P/ܢY'����i5�,Y���Tq���*��Kqw�����a���\�/�+�@� �y�7��'2O=tD�I��Jt���K58Mlk(�Ese�GGa���]I��j�<͏p�ǟ�gJ�a�2��f
{$Ì��y�E��T��O����t:"���7H�Csj�&,�x>G�e��@�G��Jm�	����3��*h���̛��{�7@n��y�Z����rHe ����uf�O�@~��`e��k�s���#�찴m4�S��z3�Ef���΅���m$.f����X[����>8�Q��,F�Q�r1�S	�z 4M���)���ٴ�	�e;�U͇�G;y���f����}',}ڮR"�n����F3{7���ou�g� �������������,N�Ƹvv����1��Z�`��V�kr���[��zj��kx�U�i�WLv�3�д)�v;� ��Σ�KvGu[^���b2m��)���@�5X֥�U�6���{`wf�P���>����C��/R�zhZ�2Xuy�k,{��o�&@dyM�ĝf�ڍ�L�����h�V>F��t`>��(a
�R�oE�����#ڿE�d���h_�����`�� wP	EsPO�ܱj����4G3�
y�]k����I��]U=�ù+{r+i�r]U�Bi)��^�.�3�|~dA������C`�~�,��2)��Y��aδ�f�.-YP�j2^ۥ���\�[�K�x��A�"f�Z��<����N�"m�����k��-f@�'�����5՛8�j(Z��*�AFu��w�j0�{2ic�/��9��_��~n�A����TE|���dR� ]'�<��҂{����/m��w��y��?s�g[o�YQp�7�@X�.2������M�2=?B�%�\�G����[L�W�'��z�j�6l�^	������YC+�3WE�����`ʻ9�՘�v��J��G�vms�Ïp���X��p�#��N�BV�y�����\��}.�l.hi_l��k�9�>�p�۹V���v�ں+1tB-�+$�5�ӏF0��ݝ{����������f�X@��f��M�Г�Z���WT\:�q����A�},!'mΖb:�a�����=!�V4��G;�Z�\Am/`�Js`�BՀ��qv:z��z�-�WN7�A�i�p�(jvb��zB��ƌ6��+��F�i��L�
0�Bb�SȢ��.���Q9
���O��e��qȖT�r��]�3��}S ���!�_v�_T��hͲ.��xsHZ^F������]�Z��ܲݜZn�3�je�wb���L"���t(��I�P9+�Z�\��eIcr2Otյ���T�ju��֫z~dB��Z��ó�����UԪxгf$㋰	TX0��j�?D�%��A��B����`�Ot���n5�!���>�3��8ֽ�o
k�)�0��WQ3��"�6�r%�cdn:	A/mr��H;Bu�vz0_�:�8oG�0h�2	�8n�P7-��+lG��]�v���[���`G%@�~�ǰ�3N��R��@���g&;��`:��vԵtL[[�I�oOOPT�<F�V&�uC6]�;$����܍��/w�f}�ϫ����g�܈`���Ρ.����&���q�u�ӲZ2b�V'y�N��2e_~~{�Hl[w3$/�>�����<+,�O?W:۵���� �7k/���3�L*��	b�ݳ&��})��<�5+�:�3��z
W"v7k�蒆�]������� ��ǀ��Zf\if�w��`L�!'�)���&�i�^=���;�$=ʀ�O�醘��<��a��ַ���<K����{"m᰸f�
��\A��c*x��zn�lk^9!�z������ߠm\phy�e�/�+�B�vϙ[�^<�5� �E<�;��#���b�o�PFv�n����Y�>��?O߶�m`���B��C�B��G�={zm��\�uϩ����[��s�ٲo^�m2���]�a�t�1e�Jm�2Y�%��H�N��M<5��;@�Df��V�P�xڙ�z��!P�7���_�j�y�Є˃���oJ`��R�}���j�O��;���j���~U���vG��S.s���/�'݆����/�:�x�5�#�
lf��.%���p��75����?ˎ�x�����T^��%_Iw����E���?I�wg��N��nrx�-ڋI̘b�u9j^^� 3 ��Z��M��`�4(��&dP~U=V�0z�;UR��U��Y~k �_�y�4?!����!�̅�鏃�����iE3{����α*^���x�F%m�ܾvy`vCP����p@���r���L��mRM�3oM��ov<�P��j��=1lF�PڛG3��mt�V_��b�zb�ѬG�0�\�l�WH�Dfn����Dr�bz;!ܥJT�tF��WK7;��O�|~��~ }������r���~�:��O_�SE
�����H�==���s7J�s׹l�ߕ�j�Lg�� ���:���^����tb�eM
!ʘ�F�&�y핈&��x�+^ʂ^��sH7Rͼ�T��ΐ���m���q&n��r�{�������vm��Λcb9Rcl���џN=g�za�ޚ��Xԥ���ZF��ߩ�P������MY�q�gא#��Q~,���H��.w_���E��Ή��o(rD�'海��u����8��X`��^~��ᇑ����O�������x��nR����~Z�64A�_E���x�P��P�
z�3����$��[іz���:1���7B��T�5���i�j�K�U�B�2a�Ͻ{6����F��ň斔&��9X��M�D�ħ����]O�1��{e��Eճvj�VE0,U��C�ٴ��V�t�z�_s�\\W�K�Zl�zb͊S@m�B.==F�#`��*P�m�R� ���4�®�a^����lǾ���g�B�~�t�9׋��/h�a{�F��K�A�����N4r�d^�Ji�!��a^��x[��O��s��Tie�u1���U�2��P�k�u6.���6��߼-�GtA�?�=��l7#=�|N<��3:���8�9E�*^��v����D�8�6A/�6��I��n6&���yy�qiq�⼕��W��D��� ?���9-��o:�ߢ;�Y\�+I�����D��?_<3�O=��O�7������6лx�>!�E7QF�[\m�5>Eî\�a)�;���Y��f
zb�g�>pڅ[�/�Ӌ٩��2��ct�8��sz�k>�l�#����q=�Eq�h�K�:��V�r��y��R�6a7C�F-? ��ryA�Xt���2/�;���Xy�q���=�%s!�':bZ���=�ֵ��E慩������:|K�{.�Ѭ�����x^)#/ڿm������z�d�k�"y�zL�SuGu[]�zR~k�d��ҐXƬ���'9�s�ެ��"��zwmr]�"��^����_�Իs���V�K��5�w�g�L��-����^o}g/};��L[A}:�G��AZ����>kNyP��Y{���Je��/aK۵�������L8���;θח^>4QZx`��f&9�C�#j����<[���Z�1�^�>Ê��.�aۘ�$�/^�x5�%�!�"���$.�E�:��XX��%�o���R�3y��]Aw��d��O7ެi���^�������8�Μ��;Px�A����B{rr4;��67θY��'3�Ռ˚q�9o5DZ����M��s��l:C��Q���!�����>�����8 {��'+�b����"cS��ŶS��ǧ�/7�lU��O;QS��PD�4��Zz�o�����Rxi�=Z�s�fא�u�dh���[�&�|m�ޟV�'�!y75�Pj(γ�Tj�v��ln������b��4c���xec��D>��y�L\�o*+�B	��a��_V�g�J�껱v͇C	�)�Yנ����~Ƣ?������_�+��;W�ˣY3ۭt�ų+��6�"�n���آ���ХbU��8�WT\:�q��"�JT�l<�m�-�ۻ<���z��*�F�f!���Y'.�dQJ��b6m��E�*8ސz5�4'�a���y������!�7V�^r7T�H�I�����E�.4��^5KM�>����q����L��y����(t�L9����2�]0S��6�<a�9�v���|Cc���Ie�]>�jn�,��U�9��~	aX��+/����?�z�_���:L*���'yj�QyF����^����sy�Gt�[R[L��&�v5��/H~=��]P�4,ى8���ܧ��w�9s�.�G�Da+��{u�#Whc�R�j3%�wZ&+����`�%Nx�*��TRQ��NC��?U�e���p�g�q������7�αv�eаa]W���uCq�a����D�Lf,�{o%��c�[�>���y��q�Zy�����L?��lR�a<��� R|ACO>!i�>c��[*��9��Z~���/�F��oR^� ����c���L�*9��,6�kX�.��p���7yi��:s�Y�(^i�3�-��0�Lٮa�Y�P6���p��3N����,�x��r`C�>����f����n����!��ó������XW��/^&�^���I��dP��XL��dD��
uo.�4!���yO�**-�͗a�����	@�2�����vc�yՉ����u�`�l<�&�Ys�n6�e��d����E��A�po�/��c�U�S���PǓ��k����n�nF�My��]7C�:�tS<XG�:N&.�̾4�DP�3خB��~���E���#���aTe
6
���{ӌ'&*�E3��pLu3Y����g���Y���؅C�9�٘nm�"Sm�R*��B�ߥv��>����V�����3��11H7��թ�C\J}�0	}^A�v)�Є�@�'@w�R�&�)P��d�: 0�'~�/�𵷖�RI�G�Ϲp�]"�W�{�b���;;T��	.]�ޱ�I��� ���
�Wd�^G���km�r�h�Q��ݟ_�s��}@��j��5��*<��3:�a���Yz�ڱ5�
I�wz^�[���}&�i��W[C������m�-��2:V�G�j�?L���un��q�iԹ,ڱdm���7�x�q��[uDb̀ޡ�uJ����:�@�쓫(�D!|i*�{L�x�s
K�6�x���A�1�O{m�=�79쬆�Z�uδ]�/PL_��T�+����ta�՘�2���5�Wk�nn�yͤc�抭o1��4WV�����
v�'I����b	��^�#z�k�1jM���a���2�l!�e�-[\�U�T��4�&T�s��D��g�d���r�����V+5�Mʕ���b�Gݜd3� ��8��Q��Ξ�g[Wk�Ю���WsKq����_ԣ�5��\�����ȵ�08��'GЬ3pg���J����w�s]���j��w��[�KE��o��-S,w�tw�x�C!sQ�S&G�7YDw:*Up�/,C���m��x�惓�sȧwu]qӁ)��Hj��]��Z)���z*
շ!)�)X�n@��L��h���C1��z�{Z�t���~��)�N90�٤�:�41���0�<%�#6��\��Nv*�;�
�|���P��qw��:Q%#Na�X�G:���,T3�F�o���V���g5���}O�3q��u��6s��Kw��&Aq�.�wtb!�)�h�멳���9���c:b�MG��tQ�b��2V��{�PJ���SR��7��itW��9�K�k�e�8�s>��k�,_ za�&�U^�m���K��y�AX��w�u��n���୊Ł�Y�U��n�fT�$��HFo���Z�{gly{�l��6�sï�dA§s��;,t��(M�nG�V�͊�1�zM�8j��qڙ����*�ea<�X�nL�3&)w1��ҍ��ۦ �G��SH�N;z�`g=��͝���Q���G;����原I4�u�ip�䃈�;(�C��v�Ķ��/d���p�TNU��c�QG[������e�wT�#�7�Q��ZMр��Mb٥�X�u�Hs���A9N�neۍ��7�-��Jb���,�/������c�"�=�Sf��΅p��ߐ;Εذùͫ��`��9�z��AH��\�WRzO>����z3��os�Ԋ����v��F[��K,M{ ��ergU��KxL����͘�ε+:&��
d ?�d;�X*��������I��!z���p���G~�ќ��g���H��0��v&���y���܇&)��S�'��[�:���ľ����`��M�L1*��@�qߪ�@���k��^��)hkݥh��])����j�O��<}�_/��Ƿ���{{{{{~?�|d�K�� �
i)M:4&��B�R�F��������Ǐ=�������ߏ���<�Z�i(
i(=�5wwHQO[X�������44R�F�����
t������

����4���B�ZJ�M:�HSO�č44�KZi��)O��Ph4F�i+Jh)� b��:i(63�P�=B��l	Z&�J�BBR�H�4�T!@R�V�14V��Д�R:uR�����

F�B�SBS[z��5Bu	l�V�hѤ��.�0�%B�IM#Դi��~�u����B�`�c�BIM���ڒ��qiC-f��7�M8��V��B1g��=�
�[�^��εZ�:�P��M��j����Fq��+e�A;�"C3�PE��j0ˎ@$@2�A@�ǥ��0yv��/;������hd�[�;(ToD<H�/ʝ��.�$8�����L�?����^��2����,���c:��?*�-�q�Pj�붱�l.`��^�A]Ǫ�ե�<����?r��@/��T/����Qt���}�b�V���3?R=��W�g��Ʒz���u9jw�}-�c�N�?Ǫ1��ޡ^���+�vf����6�(���uq�_mt=z�Z~k*���Rq.��}�0�t ��kH�5��.�F�MlEda����9S����e�J�=Z��3`R�����@z���X#�.��g��}�u�_�����%�Н���ɛa����`�%�^�G4�u,�}�t[���ޑ+9Ә�C�2"�{�;L�Ͷ�ˣ�&6GS�1��1��9��D`�0����b�M��f�z��� `<�y��>輙�Ce�E��Ǥ��c��Cg�R�g�A�f���A\�� ���4A�$���<�/���t��?�$J־h��O;�5�^��t�����CH/��o��"���J.�?Zp5g��Ff�ӪpG�g矬˽i���-�SV���{a#�H�x�_[B�����lb�^�o��i�\,Mg95���3����א/u����"'�\Wy{y{ė6�w`�����W�V��7L(�.��6�I:��%�� ���1��eGٯ���C�:���y���3_e�\��Uφ��=�ul��f�����낲�	B�ײ�W)i���S���������~�Y����s�"g�2���Ҟ��,ذ�VEw�u�!�͛O^ǫxZ�U�AEgz���?^!.�K 49/".=*���c�j+�|D��ʐijX����~ْ��}�ߓ9��{
��EIų��V�o��|w� `d�`�as	+�A����D �W(�E�M9�<����687^�����[�]�Uh�����1���y�#�G�| �ܵ�v# �,{-�h�]�t�뭈��T�C1�&��s�O�p�G��	K6צ82�e�ǔ?�"�����=�C}������!;=ʒ��`�}�A�S�*��LYz�|�>Ϛ-� �y�Pm��죲-�#�����Lpn�_O5�*]��&�t^��,���H���?k��DP��i��`�6�xt�X_�흈���;�Mל�Z��^jԍcEGs�|w�Z��P��VL��W�N��K_/�wh��|�H`�ٓ��4ț�����Q�V�^�$���o1��v5F���| B��g*푏Y[��yգ�okS�Ը&��W�|��]���3�=Y����3֍�uz�x	����B����}���^F}���s����5e��*�w`����;#��v@�f�D�ϴ��iԓ2Lf����o8��n���!Jw�q~^��?U�H��}�����Q��������7�z�A�r�Nhf�f&�K�����}�~/�~�^����E��ЭF������K�|��!�iwVv�mM,�B
����s4���@�|^�?^5�a.ߕ5
�qF�����W���m^���s������f�}y�v@���\eش��0�N����y���!�#��i-BXx�	�]:�n�pμ!��L$�bb�)��6}���׷��8�5y0�V�5�>Q��ν�6i6s��^)\�w�"��!�-�{���u���Cf*�-�?5��p6�&˜싘����['��(��/��<�z�uea:,(#$�>c�
7 ��TV5.��[��j��qiEGD�ڶg�ѧ�X�B���A#Z�_��̨�s^�΂�rÞO�NF���O㙋W��|�����Djf:#�t�6��p%:+M
V%Qo
j[���皇X���3���"��]6��>�cѥ��Yv]r̅�&���,���D�%\�&w���͊L�	x콮�~�v�xI$G�L:�~6�\��dAb}%ͱȵݻ�.������؀�=3�[�^�d�vxWU�\��Y�v�A[�@�?�&~�e��nBw�y��f�I��ͮ�!NJ�)�;�G�ԝ����X���Bc��F][�ܩ�A<���i�nVg}>�����"�z[����C�n���K?ݦa�5��`�&*��"��\h:p���!n/{1���]X�<0[p  ���B~�L9�����[�|ꂞ{Ǧ�X��~�ⰳ�;I^��zۮa�r���n�����؆]؆��7K�~�zxУ����ھyn�՚��<�n�]���������-�v����q�����/ǒ�y2�~�;�/����I���'13�ډpWoQak�}Ψ�U�O�����AiO@B��<�RP����g��NTV`�Z�D1C/+�ߥc���Z�9/M	���m����L`; ?Ut�����'����@�5�,�8��u>��e�3i0桜Ui�kf��q���qŁ������9��L�z�q��޾�A��:<�L;�'�	�d�Vl�nvI���0��8��vL����̙VU�t�w=c��hr+��1�~bpY�"���t�����!�O��,oA�-���p���#]׬�z�jx�K���-��)Ꮈf�\G"ˉ3%'���{kM��`����&1ϫ���4�LyW�v��ՙ.�q\�{([�F�듖��xsi��SS�e�DEbٺC��VkpH��������)������U�vPQ:�˼l�jex�)�-m�!��K���{˄7]�r۱�ܮs���k��s�T.N�Q{�����ߖǄ�7�Wb=ҧs4�wv��m���8���@�[됇yQ�4���M]1p��L������/�g��e��q���֘}�;�����y{n�����Q�gaT�(Vߊ������a���:%�4Bn�]�����"��A�2��u��R���Bl>�U	e^X�R{���g�u����G��v@r}f�Z���2[ϙ0
��;�7!	�y�Ju~*K��鄨Z ����U@x�u�w�?�W�Ÿ��!cX�|����և��W�6d�8ıbޗ$�P�ɯn21�`�b-)wRaO�|��a=k�D��>�L<1��*��������^4�+nҕ��a�)����ܕ�f�f�?���zu�	ɥE�����p�����ywO��F����Co������qV��?Qi���,h.��5��y�?y�|ɵ���I¯X^��<b��,�P����6��r��F�Gs��
T;���4���,f���`�@z�/#c�L�q��0��%�7�lU;E��1l4��J׾PKܽ�O��ug-�-$����7c��8��~��9Z�VZ�ކ��o�ۃ�՝N_pk9��]���u���0]���ܶ����e�-�+��u�k�r�l�Ω�E6�5*r𘁼�l�dJ��B����ek�Bl�l��}�q��ocf�l�Y��W����N�"P͵��H`�k���1"]��L;6�Ȭ�V#�&7�Q��hϧ�c�x�
����qک��K6�E�v3���|<�\��O����<�}y9>���@D���cf1=�Tp�l[1ך����n���^��DS��!��D��A���\LJ�/b^��A׮#��АF��z��yΦY�9B���4��VBB�CH�C{ձu���- !�O�[���ָd���݋��Խ'�Ε��Ὢ���d�`�J�R2a��Ϧ��|)<7A�X�B�ߜ�.~�:*%u<��kR4��9�����V��y���\��f���`[l����ӽ��s.�Y.���x��w�[E�)���֪��[/>�"f�!�%�i>���6BM�Շ��հCv/�i�[�{����,.F̂C��잮j�q����s�n��ox�[���|�ƭ�/Oƒ�V@���煵)ZN1�~sȜ�0�)�/��6�=�0�,f)7`�eڍ�%��a���)ʒ4���ny�ϑp�<�i��jf�ֲZeȓ��77��p�T�x�]���%��ڔ����5&��L��D^�l���wD=���5�&���J��4'��|��	wZ���(�9C��!�j���ʠ-��NM����lG;{y���Ԝ�v��+�l[\����en�\�?~��j�=��4�L;�P��`��vN�1����r�@�X��sP&,�>G�g���x���_��h�=7f��� �T�gײZ�߰�v�ft=b����A/ZT��f�7U.f!�"%f-|ەڮ�G�-y�[����r��<2ס;�M������/�U��,YS૎��6cb�s%y[��~���i�N$uiDP�5����n��צD���n���޷��I���n�oE�M �u2�������U#+]�N����.#�=�m_�*Y"�еad��q�8���Qhs����aԼ�:ݯxz}[~���j�sa�#Ƅ;�`����`����zsX$�BȦ���~Z�����^Τ�Nf�Q"+��~�mE�[�����#��ϡ�����ܜfg�t��H�l�Ljus kٴ^}����&hϡ댻�ca���.y���ے�jl��Ts�A��0vZ&��)́1w��s�s輾�5�'���d�g��2Y��*�y�S|�m���'?Q|�}�Z}C�RO�&��е�,x��I��֟b���a�.�c+S��
��,E�I�N���EҖ�����/�
�y D�)�+Fs<��G^W�� ��ńJ��v����(MtP�-Q�EV�������XRҪE'[�*�7>ZW��t��Vj��4j�i��n���e�7���GNw�m�����W���~�=(宫��o������6Ʋ���{w�`���|��za^���ʊ��;K7&�W�r��㺈��Cv8��%�Fp�ϭa��mz���'���,9�2�s��v�ЪPw�zݎm����2ş��PC,{�2oPXdR�J�aM@�^�Dn������;��o�|#ib��ݱ=6E!1��o�!6d�5�L��xNx�AP
d�q^�v�ȶ����ʽ;�vWds�oW=o ,=�s�'��2�V�7���'�ҩ2�^d�sȢ�q�ցM�ҕ;�v�݅2������!"1���L$Ϝ�U�v��~O,������W��U�c�|b	�����@-�M�����Y/~w���,y�s�'��_t�a<�Zv�
Ǘ�3.��Zq�*��ڍ<�eGk�T5��O~B��LkL�~c~?��c��U/%�.�
zc��򸱰��뻵@vI����ͧ\ʥO0�m��.X0k>6�`�±[Y	��0���p顋�0�hZ��N8�zV����'�X-T���,W�ę<_��e�H�K��)�j�y�哚����7�+�k��mޥlW��U�I=��~����c"��p�rɸ;��8��)����;�X�Փf$�|�C�|��%.�bV��]��r$�2'Cy�	T5}*v�$�&.�"����{�rd���xx{��"U��6���s�x�y��B�-��<�C�m�O0-�9*�O�X��	�;��/ȍ`��se�Ó���u�ɽ�v��]�ꀔ:��Ͽ�ɽ���<��q~�l�+U4ė�_�÷k�y��B"e�lO*���}���M����C�����(�z��/l��y��EU��|�I��s7�b+r����]�e�1�}����ϵ:L�`�1�j�#)���O��L���[ym�4F�LӬ�����}�*��=>c댧M��c^Y�?0����U�n�q�v4�s2j5o5�kv��B���R��Byκ�Y��뇠3f�M�T9��g�d'��h`��m=b�R�^����%��ϏF��کa>��)7�+2$����Fc�k�U�m�<��^^�n��tf+�,���:-����p��z�Cv(������bS�*Kx&����������?,���J	;�7�ɘ��\�R���!m �!�O>��vG�z��Ru�Df>�^Ԋ�sp��.j�CSu$i0mU�`Wq�U� Ǚ7�G�U�߀'�|P�$"��}{�U�c=��{����?���gbuU���厭B����_,�I��]��;�*����e>+L��\����l
��R����W���-	|y�:�͝-��˹tĬ���rE���'u�tc7`Ђ��n��ܴ��)kzYۭ]�EK��w�G_>�\�M�^^o0��9��|QѬK���>0^�t��s�1����c��Pw�w�X�3�r�o.ʗ��ӷ�Ϲ��b��
6;iC���=C�Z~k*�a��$!��;��A�m�MgO�ɯeYi���"SP���^����g,�w�Q��j5�P*�s�� sH/N7x1��6+C{�v���A״G0R�G�8u��&%��ȖO�4û��r���S9���&�C�|��9���b�6��������q{�m^�i�;6[Ȭ鶅byX����kXC��I�Ȩ�
�v�O:ѭ'�Y��T
=���_����kNyTG��{8�	r0�UU7��{�g!�b�ܟ��`cr��}w�%�z�F�\K��+��q"%M����0������q����?�ӊ��4���|DX4 za��o�ؽ�7�yG�j�CT�w��>�Z�|�V�Y'�K�{"���^�yf���;���]+�ɇ/b���m៌��T'�JU�{�پ�?�&3G��/��?��ocwy*f�,7P	M�-@v����S�ߧi�9��iҳC�;�]Z\��$MY�-�o�6[[�sY`� �����O=Ϝd'Sviܽ�&���Y�R����gaX�v���qZt.I�,�l�^kڰ�Υe-�|���9Vխ�c%�ھ1mn��
��ªe�n�T�-�xro�+{��V�7K�7�/���q�.#�ڬ;2\��o;���Ȗ��ɠ�V*e�h�s�ZR���C%qx.�mR���Kxp4��pU8u�A�ɗ���#zkN���6��P?�n�p;���I7�.�����g^��yol��9#�q�z�WK	�sZ�ta�K�O��ً$12�[�rGxn:�l�3d�s$�A��Hk3��棕vw���ٓ�G��u�b���ec�\�HX"���oB[Y�V�����v��B;N��&�|�6'<��z���&E{�G�⹊V�����@ML�o��������UՑ��	����Z��s�z����3�F�UR��$����n*(��V+^q������f���e;��s�{�#x�]�i�w'n�2�h�� Fء|�om(��/[�,{hsi�&�ib�xf魇x�)�췵�q,�����r�h�a��M���q�y�\`�c5[�M5q�(�-��T�S��ӂx�i�7��n�nJ����+�פ��i,J7�UT���h��%�9���"CH��VU��o6dE�����n���ïg`�I_��+Hz�)w�;{ [����W{�c���,�*AhW�{��f��v�5����d��l\#�hcu�$�P�hW'eT��\��{&,u��K�T�=.iPnS��w;8)J���������[z�4r=X��KG0�vC���A)OO4U�>�+�1���sWQ-Mp�F��(��xE\Vi�nʃN;����fg���$��SUV�w4e�s���(�\q.�0٨/�Iz���N���or�����S���9JE줌�X��:�CZ�P7˅����RV���q�5C���R^k��ӭG\��K*��y�����-��ѵ2�/oJO�s�GD�lԕ&;���I�S+,�"�Y�,x3z���f���&+y�>C�cʬbF8ܒ�S^ں�GA.=�Z��Z=5������PI�B�@�[QE8vȸr3Wƪ�b��U�s�����/6��6a�f.n���:�ޅ�\YS��;x#B�ܽ�Sn�Q.��+L,�iU8�ռ�S�tK;!WS*��1���VMB7dj��=�E�ϑ�-�z
��׷X��9�Y��5��V�v)2��[ePm���ӝ]�Au�+	KzjԂrn���C,�P�k�y��R[}Q��N��8��D��)�����n�d��(��>�T��2>Q�k��Jr��n@�����n���z���Ұ�V�Ǻ��3:sq&�k�;�3�}|=����i
V��H$�M DR�)?>/ǏǷ���ooooo���}���a֔�t����4�u/wR��SK�������x�����������~?�r]&�P��H{����)O����t�	O �:�:��4����ZZ
F����
GE%���B�Pou�J@:����a�*!�bF����+A�l������ILM-%&�OD��A�*���
��$AAB��-,M�]ZhO��ź�@4��B��/P.�z��-x�� �>g�?}���.t6ml�w_e��d�7���M�j��q�
���-�v����o�R;��%X�w��Z[�U�v��������\ͅlf�4_�c�?HR)��j3ГЌ�L��a�򢼸�M��Pd�w%l<�֎'E�@B�/��%ׅ��a]�x��O	�vd��X�ffoU�z�! ��=#�d��0�sU�XR�L��X4\q������LK(Ъ
7�=���O�Ȋ�gN�P�c�swS�Mo6�k�u�U�]��tb%9�QT-����k�"{"��tzql�8Z�a>�\�V<��n'��I�z���e���q;�^G؝��&�:�*��5x�)�������i�Ƣ�Y�4��<s?_n*�X,G�8Am��gײ$��m�wF)?"H-!iy�/�j�ȣ�f�/كiS�e�[�_����xe�S�4�~�T*��\�V�&0�Y��C��N.�y�4�}߮,6����Z��x@D>���ݓqɑ7�=Z=]=V�Q��:�h=���{�sX8bi�jx�ڹ�}�2�ϥ�N��3�ܷ��~�Q��tâ����;FN^۾�{���L/������F1���W�D7gC������J~�D%_|�˟��U])��)n�ka�"���l2�W�����
D�:M}���^��/ޕ���	*�����m��x�(1�⸴.�ږ/2qk�᱌�v�&�)����n3��N��\q��{A�n��
���82�7����,�#�V�h�^�3s��fm�&�	q�'�����L�տx�$\7D��o����Or�5$ԟT�� SX�r�#;,~��6�����@���eۚx���tE�c���HP�Q�4r�;��2��["]1�^�q��������������~��U�� �ޟ���6�M:Ξ��4��[��6�d3`N!��Ƚ�\��Uɦ�j	1�F>*���80pc�'};�[/,�g��ɦT:���9{�n��~��T�b�)˃;%o>ju�?��gs��g���.e���g{҂{r������1��E�T9�����X�/��\*��ܒ�����E�7���d_z��PɅ�^~�k߹BeK>t�J�υ0���������	T#�>fC�b���۳V�-oc��;H�������	�{"S����8�����˲j���ͅ��P�P���zCǭ�'(8�rO����N�Hޅ)���.,O%��pWU��!?ed��~��1���gI�7C��@A�����#�dC#|i�o�JzΓ*jy��̆g�ڟ&ٸ��*X��ώ]yKX*�j$�p\|�{�j&nX�q�v!�1��٨Ⴐ�ʤ�	d3w���]ö���=�f �[�����3R�)�Eֻ\ʾI���`�uԷc��3�l��bIl+������W���*��2�+��1��M��,?n�6N#�Rg�Dz�f�?���g>�A�lL���\�M�G-^@m��8�nv�<��E��WmW<��*~�*�ަD�}��P/��_��?�o�_!������d_v6��(M������*�
�d���Z�B{mi�=8x������]�ΑK.��l�_X�i��q0����Ƚ4-Xs'P��{w��`��p�����u��T��Uq�%�ۈ0��f@�����|!ٕ�O0M��P6�����Esz�UL[D6c����o,K�fa�W/��P�t-�3����@�xD&��bc]�|�v�ʓ
ė�	��&i6e��g�Ag'i���L�����^y����S�
Ql��Ӱ��cb*�.��1Y�� /di^J>��� �i��S�v8f�	A�ȸI�5��$��k�ݼW����s��=nYwC���.�4;_9/�\��>:-���� �
v�ͬ���9f�3"o5��%�(��UU^Ե��B�vd��I�Y�l$\�C��]�r*��ڕ�kf���Z1� �]�ljp��J���k�o(��PI��A���B���V교ge��[�l�T�זV�;G,F�cR�Ziӆ��[�n�	:� ��;t��p�<�nr\�Ӯn%�*��r�r���m�%Ev1h�֤f�oV}���� �a��%3�W�Y��Ѡ�i��k�%�U,8�D&��!2�*�Į�PY�;��~u3WYHGjk݅9qmV��ףZd��\K\�zu�5��KzKPs�SW�1)�*�k�*�áz����6�qT?P~���Rye�U��3	�-�"2`$�/�&;�h�4l�Ó��Jj�Xѓݻ���y��%���)�$i0�ؾqOw0����0͋�0\�E�{��V�5��8���OCݛ����㼥]0�ʥX9��[�:�D}[�#�u]Z?���Ϳjg���t�i�W�e��ֵ�Uvv�f�ˬÉ�S���-?5��,it�~j�N%��}���Azt��YM���m����?�x��?������$��	��E���Q��Q��2@R	r�mma��KK�D]�.K_iK��p�kޗ=k�LKb�NЦO�4�r�����O�iE3ɞ�7�c�?i�,ʀ��W���]� h��g��r�}Y���Y���1�2úZ��!ѽx9������l_����3��ݓ��4t�BQz�-��>uR�yS�e����f�귱����u��s����[�-�[r.��p�Q閛U
���q/kc�B��`鼢�d=�*H�NJ�ָ뫙+�R_(�����5��l��Q��P:#̽�:c�������:9�9�^��a�����@((_�ՋR����O���Q������ nP�u�hP�ΰ�ji?�.!�_���__�~����3ot�z��Z�K�*��A�Fua����w�z{��X��K��[���%���F�3�%�����A�h�֘r�=Kս,��{�r��hwIa��U�B�5�2��ZzyB*b�$�h�/�33�)�L?�!a[�������W��4�rT�B� �^Jm�kGrq��v��m�>���T�_~�x��cΣ�`�}=�%�EǦTͰ&�TW�ˈ��WϮ�3���P�d���ѧyXkj׌t����ϴd^<S�3 |�_`�a��G���됞�y6���[CĲ�����V����Q,���YB����}k��t��{w��`dO��vj�G��ף$L�*�ܷ�ά`v�|�=��,���Js`�ƁF�[X����ty�.&���NWw�Ъ͍��S/AR���V�0���q�ԩ'����t�2Usn9](�ve���ѷo��}Y�ΆŴ����"]	���!>{��]��$��Z~X�G3{�� ^-�g�����^�~"�Wj'�&��aV��Õ ��\�&�0N܏v��u�y&	R�0U;%���c|f�l�X�Ms����Z�.�ޱ�.9��$B{7!���.}-�c���ͮ�o��%O�U���]�E�brʯ�'���?�|����6OCҵ{���M3�4��XE0!8�C���1,O���5��5\�ʢS��m��ʛ��W���ׅ��ʀ�� ��GU�E�c6�@��;&�}2'�A�-�2��%�	�X2!���bq�*�x��]<�l+��cb�٣���}a>�1t\�ڜL1�j* ���;��Cw�/��L:���{�UA�֯���ۮ��hp�i�`�B���@�c!�Sץ�>7���t���O�L;7�W5�nZ��`��%E����,!���v� n��c��V
(w���Iy9f�1�q��rv�ϓwn����^{S�c �?����K��i���ċ��k6}y}�~�i�8�y���]�B���| ?�{�>:k�r�����7��O�Y��"�5s�y8�XU:��1T*ͬJ;��p�#C�%r�`6�ɦT@�t��N���$�v��.��;�9J��=oWn�ڊ�6
�O�ga�nc@��g�n$\�C��΂�}�Iv��).�Q���p��k��,����b�,�ɇse^��^��SsNVs�ک0C¢�Z�	�;v�Z5�zW�郡U��#��_jUR>����w/DOtE(^�L�y��3�a	�(<�Y��Lǒ��`��Yv���E�jL]ה*����??.�w�J��nK�Em�d��K��4���q�VL.z�D�_��G�
P��K�g��v�xvs�-��R��~�ϖ~e/`�ހc�]0S����}	���Й'�)�FB*d��rՌ.b���B�#������N7�C�A�AA�C�e>��n��0oJ��x	�ۈ����B74�[�1�A�^�P��7�aޭ�c�@��>�.����_Lb�ވ����k�<�'s���'w�^΀)�u��iyA��ȐuZ
��~~��r��݊�L��w���-*P���C���BԮxj��/eAcK�C	O�;!���m�t�����x�S��K���Լ�5=��q��⨰�]<�oԫX&����N5��ͤn(Q��Q����ƿ6�a���Le7���̜qD��{*	{hO�4�:�Z���m=#�I�7b�32�~��`��g@�g�3�|�fY5�{�X�Y�`瓙�t�F-f֎�ДL�-Wx�o�hաX�o<�+��Lh���3��s�<��vɽTXC�ɣ�/�;/�^�c-��D�e���
�.O���1|3ax��Y��c�����b{h�bzw7Deȶ���+5+���0 �9��7L�1������\��҆�q�1R�=������`��L�A[�܋8�l�=b����G����'���Gfi��yۯ@��}���sW��`~a��g����g�ŉ��F���jb��h;M٩� %<.}��*��1�g{�%�
����Z�663�	��\.�q��l�JHWv���^��Omyѭx�q��s���W!
Dך}q�髦.}�,�Y�Tf����/sv^̅��h�A�B&��T	ڽ�kװ�H\��A�,��8��6m�O>m�jqf��]�7[P���x��c�4�;�%�B��Kfa�o)���!2X�Jw�+m�!o4��X�e�6��x���C��S�;hOma�	k�	W�i�S�O�Jj�I˴��?k>m*�R�w,�ŝ)�j��vd�=v�t��p-�����"*`$�/�ئN��N=�)e��ʲw���E<K$�5L�H�a^~�.)����a��!0Z��ҧ�u�v3b�okN�r��e;�ފ.�_*�]`�cKz��r����TX��Z뇗���AB��_�n�8`���	�&U�D�=����*z�E��T4�L?2a.����D>fN4+%��_��-���N"��x,	З�i2Fe:��}��h�Uܯ�k�\�dq���l0X��}uj�=��kG��S��I|����N����}�X�(�r��{ݡm�����1�.ֽ2�nUk�U1u}�+����k�MU��|L#�9ni�#Y�Ӻaa�y�5gG�8�*L='��@�ϑ-O/���]�^2����CYz��>�t��õ�G��k�LKb������gr��qCC�*���x��dB��QOT�ꐜ�D-�<5�y"u~7􌜵W�6ʁ`�-R�����wZͫ;�����	�333
ײ���jY����#`3?�tg�t_!��^2�%�*�%e��Xͽ/fE޳�QnWt��>׳�c���bR�m��gI���a�Ʀ����'V�g�����A���K�|dhf�}Μa�烑Šza�`����&�w��\;�&e���A�����V���Y��y83k�//��k�K����,j{�.����J�u�ur��V][ͼ1>yh�闥�[�{�NlMO����cO�%L�,�ϯ"2l�1U�=]V;���U�S+=�6(���:��N�aŴ��1q�)�`NKϐ�
���k&�(;��ܚ�Ep�Y�7!�<�,�.WF0�z/����yݰ ���0D������M��@�S��{��q������-ݩߓ��:w]�¼�,y%�Uwl�����o��d')nngN���&Q�i�\�"ǎr����M���qj͉��͟d�pne{P�缭�����n�a�縈��-�����N�vM���j4Dn-������/��L��9���܄�G(�E�4�įP��n�d�++�R����Z��5�Ki��zn�\�=�*m٥Lh`d^�H����'.�QR)�FSSvN�e
틇N��2B��Ww����u==gu(�`�c\c!2��3T9��,���F�*'����(�*��5�.�n�mw8D��i�
e��y�t[@��yȄ�Bc�l��D��|��زO����_l�L�
}o����Ras���l����6�	,W��0�a(�v#�_�ᖽzw��n��B���X��Vph�]��<�� �K�)�*�� ǓH�vQ�#�/ܧ�~8bk��	���;nf]��O�|ޞ��Sj=X�`-��U����=��F�t��63���x ��yb�N(@�e]632����^�!dд^��5�����u�����d;���`̒֜�^��ݾ|2�ɤC�\�%�>^��:RpStK��8�sW���hF�K<��p���t�Jmz�#��a���Y�z;�s`Ld�6�b5�Oa�@���C�G��\�]�~���U�l+鯜���ؼ�|�F��I���S-^�Pd�)����퍛�e�Ë�ǖ�����n:��H���O�P=���f�ۋ ˹��d����+�2�7b9]�,�`����j�㷠�itx%c|�i:�놧�_u��`u��d�bӶ��܈��?��d�c}�pj�EF}�B�c���\��%XX嵐�髮�:!y�J��-��}�*ܼA�|I]�Yn���݇��&�KL��}Xm��%\��7/qf�읢���S�΁n�8ȃPV/&�����q��;:bZ�:�r�.�u$�ȝ�8�Ҭ��:���6ӷ�V�U��ֆ��2$i�1c�N�7��%:ݰ��1�J�[�;�j��������Wo��M�ڭQuc�c;+K���.᫚��	��T����a���U�C���`�)EZ�L��n[��ݦM���ҟn�wwA�S�-�L,�2��ذk�T�\L$��8�E�R��.֓7gfՃ�'a�X^�U5��Y
�-���W]H���k0��X��Ml��bgnԻ|�,W-|��G���2�Q�L!��m��.�ƨ��a�$peP8ۭ��9A�>���C��m�U�9IQb�T�W wnk�)�;]��r�ڰ�̗�]����aGV�����ŋ�%ͺ^`��ta<�k��Wo9������Pr��o��zk�z�������-���!oF(s��k+(}��h�~� '�R�G���]7h�ڤ�����#w+���<<�"��a���j3��WIRZ�n�7:��"��yaѡ�9Εw�a��Sl��6���,n�ֺ(:o�`�y���S�%�v��s�ջX�T4⧗9�7ئa�,V���X ��d�;Rl�nfb׳`�o(ݪ���0�k����t7J#���r,�&�#����k�j���P}�|���HgoB�QnG���.����r�{u$���l�}s�7}1��������)qN��PV�,�s�9j-
�ځK3�5��1�F��;��i�>�S6ձ��t))"��1�!wu��Nh%&�brA�N�j��iUp�yk�vu�':f-�n����{fi%k�" T��*vPJI)ۻZ��zޅ錜�(I$B�Jﶻ
�8�¡�g!vOgZ��pѺ��Ê�2��f꧘XO�6���͊a�m�L�� �{����@���gəD��P6����٥��n��MGy�QK32�ƺP���p��������if�*)R�m
E�u�%��W5u�)wm��Ql�Ia�{�8�Ǜ_-�if�c
�4���y��ӋM��6��移;� `u++1px�Y�=��z�z�i�(Z�w֍-9)һ���c6��٨��S�/�M�7_z�w0�1y)ة����=�t�hmVnE]���cn.��90<��Sb�i%F�d��̘EW�@�S���F���Ƽ@����|>^�=�����g���������NJ�@�#�h)>N�$��O����Ǐoooo����������ZA���К�((Кb�M{�4>$�4h4ht��
PҴ�P;d�l�MP�R����90G��T�y�'R�M	B�4m�"A�P4����z�x��ń3�
C�:�+�� iB��CAC�4� P�]�]mѯ]��Ux"�|AUE	��+5�^m�Ge�F3\1�]�dhfj\E_E[����kLg���y��4�6�,�!�9L��S{Z�"�3��.��%F�(�@2� �J1Da���m�$�g� AlSq"�4�?x��6"T.�U�u�B��Q��� {)�e��j��M�$�|a�{H5<k��U�=5�7�#����v*��|�$_?�W:(���5�沩����/]��9���2�Uw_�AK�(?|g������p��}����:�� �+��Cs%P�h(�i�L��[:y�x��3��љʪ-RO�� �j}{`�7�**��k��-`n�	�d	cEuk= c����*��f׶���UKpp����guM��G�	�q C�;,�d��<��2��钳"J��SQܝ��KC�;��%k�Pbk�<ހ`Ⱥi����$�M���~1�ߊ4��u)5�YŊ��Φ;˽[���m��o@����] �D9�V�7���*�)S@���~ˡ��Ⱥ~,��?�����'�
��_={��3 BF4�'�sυ�	e�	���(;��=�٥��b!���Ω%�TS�9����|��ä�f�j�?#�`�����2;��,�ޮ������gRaVas�p�r��PX��Q��<���{{p�WK�����`���A���S�Lǈ[�}�Nz=-����]ҡ齖�/��}���~�wk�o:���ڲ�m0�\���}4�FS�Z��r���-gg6d�.����:���T��J7v��y���.���θ��t.3��������<��y��-��YkЗ�ꀞ4	�(�|U�a^��̦��Z�B=N� ���G�{��3�bj� ��0t� pa7W�1�2)1>�����{�PK�X��:���I�q�,738�[�5��
ڝ�`�%>`���i�����Y<�6�%@��y����/:�Viʘ����<��[���������0�ć��A�q{c'�+Dү����!'b�p��)2�D�bK�J�Y��jD�Lk���l��s˼&�Sϡ��_s�f)���vu�{�X��� ^o�kjB��\�v���f}��g�%��E��5�y�����x�{�٘9�p�t$�'���ٱ�"�
-|矊�R&��.6�5t�Ý���р��^l��e���`�a��qqw4^�Uz�{R��)�����@�*N����0�ٽn�m�|�ף�a𹋇�yg���m~�;���1���R�F��o���s���=I�HZ�u���V���S�ܳ���G��~5b�� �+��7b�nSO���E�Zo�s��w�?zG*pc.�^�.'�v1>罭Y
[���NkI1�L�l�{l��.��J���ئ傅�i4{��-�%f���׳۝hn+�X{J6v���tފo�����]oN�=����H賚�ӗS�����w��FA;�7�܉��*KΒ�Z������Ϗ>��x��垄C�����.��Q�3��u���n�@�w��Jd�X^%�{���e0������OZ�� �5�s0Z�ݔ�]]�����u/���@9})��[�e��8�\�Lk�z�P1�噃k�N%)�u��,�s�t�"�9ق����	�E�P��S���a����_�PX����_���5�V��;?[
	;�<6��9L#����t[!ຍ�a�خEJ�/V�YD3wnWWK ʩ3��#�oI����� �U���:9��2����j��,�wU�KoT�mZ}k3aF�dv���ٌ��t��b���I��Zx(Q��X�C�y�mt�^w�z�Hw&CfT���}g{T�^�48'���F}8�8�4��$�T
�k��c���/͎�������1>��>˴�*̇l��/��eH|~r����SA5��&~�w_
�Bި�
�XX�CN���LelKc�u�kCOt"��- �$�4��o�>V5��C��\��o�����~`��=i��?nۥ���[z0T�c�in�T���9��K2>���ꛛYQX{�=�_:
����y�0�.M��/�?v珫�+՞�L-Ֆ�8�'h�y�CW6<֩����7�#�r���P�|>=<тx'�쳺n��4!pZa�$��z��y����f��Xut�I�;)�e��٥�=�w���+���KP�(S���}����-9����ׯcWG�vg�<�x;�VP���c���X�"�c!����n��l�@��a�{�"�/�)�a���Z�)	�=���z�P��ܼ�Y�u�����Y^�����馞�3���vZ��{-����r6)�?n�P�u�@d��tA	�'�E���+�
���\�ΞE=���톺�4[���#�r�֦�/D�!7�y���	�{"S�*E1(�jn��+����1Rζ��������H�� �f�C�c[�`ܞ��J�|�1	���"��mm���e�����L%�|���F�k�G�D&�~���^�|��}}�;�;F�p35'�p7W:�Yoz�l�c��n�Ԉ�Av�?�Lxr���{�3Ln�+�0�VH�q��{7���5�x��^�Q���`/�b��G��>`�a�q�r�B^����k{��uz�����g���#���K���V�Sǵ��ft��5�u�`]x��Z���A����d&���\h�ܙ��%I����&��$p�mM|d��˻uTr�v���B���6�7ۮuI"Ɇ�rù��%�lQ����«J��)�T��T���	
& "���)����[]��)8�k��ʧ��b��v�/�D<���K?
����k��G+�
u��α����}�Q�j�Ia�Ʋ׾]>��֐_(?�mv�f�̇��b��KPG�����Bli�ȼG���鑝��I�M��D8k�ײ��m����Z>Jn���V��r�����$ܙO���E����Z��̕f�}y�v	�.��lv4\���5����*�ݖ��(ke�8�DY~j+�6���A����*j��^��~�|�!�c<��e���%n�!q�쇒��HG�-�kZ}�o��f|�l���f�%�CS�v
��Ձ�z��n���ƛ��U����Pj(�f�����ŕ�Aʒbǘ\׵?0�q?�����WѺ�)�B��
���d��\V�aA�&�]�>=P*%����]n��LK�3Z�c8�`5 �0��M{%t󐲽�g�̚��peq�-{�ji暈� ¹��z��jѥ"�xG�=��Qz.c]T����NV[7q�8��S��C��X�4���/r�[�+w��s�X�sK�g7�ˇ8���m!�5�!/�E9�op�M"�>5�aDյ�l�yTZ����ή}`�V��� �r��U�/8�(�3Tg=yB�d�d��q:�!]2�W�;��� �v�Y�;v���q�S�ng�#�/c�!�!��(v8�j�5nL�x�n��$��ua�D�h:\d6V�]�Nc�F@t�}k몤3e����Gs�q^�����F��U+65џyo>����a.+9�TK.�SK�9��g��{����c���;����B�[�ʛ�S��/=���|���f��5�)gT���6$�P��;��8ɠvU��E��+vU�i���ó.���ͧ`a0p�t0K��g�M*rnA�Y\{�M�ն=:ə1wz�*��U�[��0Й���8�M�-�_���p�äS��Y)����n��܌%�;U������F x��e�$1���ܫ��̖ݎŬv�;9���Ș;�-�<c�GX��s�ԁq�tC�dC1�k�4��>J^G���yo��;�"@�����"�ݞ� *	��~%�jz7Y^�̇5Δl�f����א�70��*!2����G��b�������t�U���R��=�����,銣hkF�<2�t[�u�b��4*��a�dS��rkq����w�dpeS�j�=�j��\��i�ۈa��&�<��~�`=���:7#_�N򍫥c7o����U�>D���Cd_z�vVM�?:#D:�C8�r���S1�dT�Eu�AHWf�U��g
�.�����s��J}sNge��*�4�+q*Ɋ�+et ���9D��f�8[{�]�/��B9 �܊�s5l���Y�$G�aq�tٞ�2���Ƿ���6Q���:JZ��L����	��>L�TDC�ό<gP��:ѕ�(�Hޒ�gG�OI<Ux��v�� /?e�?��K�E-�X$>#���A��di44��~,b��3sR;�k3���a������kA���}[[^��,��u��^k���(�1��~�U�9�'��a���bJl�(yY��.S�ݽ�*�F./7��u�m�+���\�Ӧ�i�,p��0ހ�oH��g>���7�����0�5�N�oKjn❔�.�[}�����d���ۻ�Y���ty�ҬA�>H��ڶ�K����|���.���c.����R}�B*v�A.9�h��cmk�At�ݦ�|ewh�{�z��l��{��^7w��������z>�y���=�ƛ�';������jat8��O��b9�G��S�D3��W�7��AWy]N9l�8���Ǥ@!�9�G5q�fVٴ��xpn;��Iw���a����Y�zz�� i��|��3E_�z�(��{>߳���c����%
��*���c�D�,`�;�a�.hؽi�/X⒨�����]A�$��9��u�$v��ϲ9��h����?�dd-��cǗ+�-c}�	�,�EY�����/*㚤��h�<���D�~�����F�Q֑�JA��}]M�m��V�3Z������o�j�q��=R���[^�J߳��H�\K���ov�
�ܱ[K!^Y��
P�A�8.�/���@�*��Aeޫut�,A9G���uC��|v"�?>���ގ˟�F���*h���_�3�O���DK��ݨ6��n�Ufch�w�Q<������Ѽ��o|�sO�� �@�O=������Ϗ-�H�W4�)�7�y_t�ے�]���<��,gpY�r�<Q�g\"鴬*2g\�͔n}!y���jk8�_vs��hgC�|��y��
����e�4�ܼ��;��/�S����*�ٞ�災)+�\f��<Ƕ�q�t���Eu�@#f[1��5{#�l��s;��A/6=����mm;�7Zw'���ٺW��,���X'��CtC��DBމ\�F��S��ۚo�M��It���W�iU]_�7߻���U�o�MA��檝��b'��J���]�����9�M(
�}���g�*�Lf��;�{����b�'ܤ8I?]֚T:9u:��t��rE{T��.f�fs�xnۆ�>a�#w]��x,�Ӓ/���R#�c�$�(�f�Fb���bM]f�!��t6�i����}KM��Y������/��f�VT=��d�6�v��nA�[/kI%Ή7��� c����Uj��q, �\k-�z��T�ۡ�x����-��Nphk !F&/Yk�������rw�foy%{7��9٫��X����9���� �>8�����b��%�'-�:�u�N�� �ts�o�}w���F���g^�C$VoxE�ip�MG`�Ή9��,<�d��w,�V�2�椻�u������3��g�>����4�O�S�Q4��r��|GJT���@��:��C3r�ڥ�o7�s$#���4��Q6�!�=��� AJ�&��i �L�׮��&��I�᥸�u�}ɜ�a�~�ѡ�����dӋ�'LPך�{����{��2��7�B��wLK�L�����$ 
�+VȠJIl�!���36�Y���}zzLq��YZ�2v�	���w~n��0!��c���T��//۽�zy�J��ϒ�!��Cg�������^/���+����k�okOsGm�7����%Z�q�������ɔ������?p��Z��ظ~�Py�J+��_8J�
/"�zؕ�s]%͏�b�W9�x(\ed�i��c����t��z
��d�괮V��[����ͪ��s.�eo�"*�	�6��������H2b@=�d{t�S�Ֆˋ����go�J�[�u�7zvt�(M]x��J�'��չ:�nF�Ü���w]J�E���n�C�
$�DY�e�Pw�6'gL��:��A��]�܂���,:=�|ۇg`O0��a{� �� �6���
���}f��n��1��/
hf�u�p^�����^�^�1Zo9�t��|�0u�j�Ǝ'�sJ��g6�}�ޔ�k˖���c�oku3��eTh�H�=C%�V��ۚy���3�*�Su����գӯn(�u���C�r�x�V��r��p���9�ڭ���N3IsZu��*��[m��Z��3 4��׍w���d|�rz+,�|6	h�z�\�Յjѩ�y6j/(6B{A�(�4zi�p��:M���EZl��(�c��Ǽó�E(/"\S�I7+wl�Ma�K�/�./�й���������Y�%ו0e4��{��v	��P�5�ͺ��n�Ci�{��kN`�.1u�v��v��n��ÜgE�{;��y9�j�U����yL�m��D����7�[���166��Ț�"V�CVN�{wԧUs:+Q5��9y�-�@%�oV
��y�jt��N��'�SZ:lӶ$���*�N���X6�K���o+�ɞn�m��w�a)�um諦V �*� �vԞ9�w�U�I��q�*��˨�P���;��C%`�ꙷK���8)c�n}$9�n�
f��`{��6��^]K}!���e��f�c�k6�F����|���t1�p��<��#v\�Ԧ�u�mB�Ls�{�N�������.������í�;�nM��f
�7�,)3�;[:��������,3����kt���Mo^��W;�2К�9�dpV�0p��ie�LVR��\ӕ�eǤ�A�[��q_:xl9��$c��-:ܜ;VmY�Z� �
)�xr��{��`P�W�w�*���͓��L�jU�Z�q��ӎ)2m*)ܻ6q�κ'iA���Gݹw��t]���q�|�.������\��bu��Xr��S�<vm���$�{��f�躇R믭�ɉC
�U&��v������<ʬƭ�L��`ʾ��q�&Z��ܶC�&��le��+�ځ;�YQ��i�KtF��hv�������4�QxҸ���m�M���/I
���A.=����.n'�4ޘ��̸Z�m@r
4l����/"=Pmv����5>�ޭގD��È�g�>B��T园�Z���n�����c���f�	�QYn,�uUG���5\��&	W:p�-��0�ZAUJ8�G]w8�.y�(�ܛkJ�j�7��Ϋr�J=�e�D�,!�իx���Kr�q����C:����ZI�=Zּ�*F�;Z8�s�J�^�uƮ�̑ R��n���eaD�b^�e��2v�%Wq����5sX��;�׏^���|�s�� u u)�#��MRS� �	��|�^?�ooooo��ߏ��|��N��^�GR4��AA��,�~>_/<{{{{{~=�����y!�܏P1RJ�A� ��s uԇ���[K��=@�t4��Xj���Ѭ@Rtd�u��Q�^�u��4�#BP'RkN$u��.���:���������M!AZqkHǎ�JU���SAHP�+Z|�SHu 4�h
k�1�
4����)���j�҅�'R=u�m�^5�5x�J���E!���:>�l��l������}{���o�ݣk�sJ:�9�V��s�xi��LVnnES�:KǷ��ۓ��\6��vǾ��xY�y���9�z���dl�7o�s_��a���P&��D8Q�Aw�Jv��k1��R�>M������ɠ�op=�h�O/�7�e���lK���kC�m�ZL*�����:��ng����2�\��/ڟ{�=�*�g�6�������g���3��^c43�3|�y�����tKv`��"4%�ٹ��n��"&��DH=ɫ�-��jx��)�ewE�Ʈ^W6��l,��L\I���ǛZ��)��k�u�/"��vs���ۍ>��"�N�:�y��ض�¹��+��יxs�h"�f�[�b�B�;w5 S��[:�d܇$)3S�R���n[��I͈2o[u�!fqB��W�$�O��w��eL����1p�u��:�S8�d�#�z/�ӽB���~KxUC���MA��\���+/Y,ϒ���׭t5cq�Q�}���TY�4پљ��M�]ǹp��
��M2��:�����"���D%���'Y{}����'���}r�������@�;��eVce�Ut�%���o7���$����5���vВs�������¹8�V����s�M������<�M���͈�7@j |B��dޓB�h���i��ͨ�R)�~�\ו�'�0J~#2~ˎ���,��6�R#;��5�v绒�w���<j�Nz�9�0Ef�ϸ絤���;���`����W��{n����-��w��IqX�y"fh	Y��T�������qb�Ls3�UR��{���I�j�F���]^c�)��Ǐ@�t���&�4���#V�f�������8Ǟ�f��O���z��Uu��ލ�v���H�MЫk`�we^4�m�p����Ψ�O�#%���3��<X��]*b���x��w[H퇙�ا�*�b�tߣ�O9�}WDE2��l�/=s��}=ԯ.�.%�o-\S��%��Dy�j�^%�߯�P�k�X�{O#��3�}�|Zl:�תwd�m������r�z�9���	.��.y�������E��v��rs+N) �N�M��քWVU�L�]�a2�A7���%�'8�9�.
��^��V�L��N�?}������j�~��|��~+��H�e>�+V�ur�U��\_
<7|M#Ei�ͥ ]2����6�F\t4C�I[��{�Fo!s+�[\�S�q�8�g�z���3^��'�o��m��MM�6��BقD�R.� W(\�R�B�r�6+1�X��~�f���[);��g�5"�C,p�_.�H���8���kI�s;q�^�Nf�.��3}�t�>�l��?85g�9��Ik�8p���_V�;���!�v{�uw�i�^; �àv3�Uk�'���;"�9�k��vo1n�K��>�9�w7z�[���]sST&q��셼[n���z4��̎��&�3EwJ�u�
�������B�M�|���<Xwp����^��GUu���+�n��iA����z'��U�u�)Q��x��h�Ak�F2��Ү�/��V�"j��I9gkS�n�_^ڱ�tmM^�p����tu���q՝=U�3�E�����ƍ2�D���[ӯ'<��	���j����V՜�K�ą�Ъ�}6�RKkY �)Q%fJ�u�M^v����J�Ɏ^��3���̡cέ_a���h��͊QWR�;y��|�o7����bߍ��y��Pc	y��b7b.�iɾK�����n�Y�cŏ[{���S<���O�c����Q�ϡ��C*��rJ����xn](����m6bb����7$ύ�Sĺ\)a�P6��`��<%q�=^+����Aɻ܎��¤n�y�
�׎]j����b�z��?���G8�vB�H�H4:�/z-F'5�{x/x���:R�(W`�ͳ�^����J��wJ�/�����=T�6z�LT�KW�AH2I]�Όo����x�.���sXD��|�rg+��<��k%t������:јpi^���N�)Ntw���l}�	�lc��&�Dj[�+V��ljn�v��#FF��׫3M"����Rk�U۱"�$��
��E*C�������|4�P!	��\G�s���z��\pSق�L������O��h��V5�k�/<�,�qF�\섧�/��I��+���K(�r�T$ު�`�&(��l5�v/�`���q����{�;�dDβ�DG2��onԕ/��\4[���4���9PVö�a���q^���|�{y��3]�<�_����xD>}9�˴�!6�A�Mޮ��T�:��[ϲ�Ha��>0����R���덄r]���v|�P���#@��y��]o����?'�����G)�4]?��En��D%"8�:�ywֻ��cYK�땆�#�n��6���S��`�n@5�%�����`�w�W}.��.����#������B�dl�7F���g���8T�������z���G{Q�=��׍e�O<f���4U��Bh��<�VeԳ=��dM��Q4�XD�g����Pɟql�mq�D��s�;�|;�>޼��������c��ўA�6iW��Ҝ��̶���>�H�͇EhΩ��\�ۚ�m�0�}�6���l�Y�A���{T�R#�����$"��Dw��N�Ƌ��%�W!�_��X���BMw!�nqj+vj!G������g!�W�>;��ܽ�J�wn��5!]�Y��*.v^�=����Ef�ԻQ�pw�7����dk���r>=��~���t6�Y��+nqܖ�m��y�䎔6MȫAeS4�*��S�#�MeR���]�.	D�l+��%�<]y�|@o7�4�.�>��!VZ��GX	ͭ{oK����P�\?GJ�H��j���=2�X��t����d��b�B�c�uSNj�V�dٻ��3��lh>�jY�_��ٝ�=�����{�'.eλ���k�B6�M[[�3v�[�]��a���	���!�f�pto��zPJ��X���S��c�0��(C_p��w�!�Ty�-�z[���}��oI]|�c�L^ӝ�wZ��o����˾�v�A�X7W?��t1�p��&5l������ף{�a�.�ltd�N`n�=~�K9\_������,��ʘ���b��D�[5tҕ���;Ƙ��E��Q��8�ύ��i���!��o@�n�����2z;8u�m��"�e�ҡ�V�FJ�������g����#�؛��7<�uE�n��P�.ͥH�q��J���n�t �; �!��h�%�3�~�vb৪t:/������'�کЫ�o"(�e��	��1٢�u�J��btr�&VyB��U� ��9:��!�,jF.���W�Q��V����˞�]q����w����ظ��9�SL��tu�x��;I)��P�����s��刼6{=v�=��B^���g�d��,���j|��=@�L��nN��`jں#��g?qxj?��#G��U{%�b�ۯ7����}���캧�ٺ�d�`���gu�R��s#!�hB����>��~�uV�OR6�^���sf�D����E*CB%�VR��s#%�s�AW���
�%F�=���M��vv��HP�C�4�G@ͥ"�l�C�g���������ݦ;�w~{��Bi�ڙ3eP����2�$��㸨�����O5��+s22�N��T�=�gW~��b�8�~����������i�������Bu5��Q�n�S�� s�U0��z�"��>�]\�y�\F=^Fs��k==;�<e�iv[�7 �c�����F�8�l��-;�FoC'N�ue���= ��Y��x���_��BHW1cxy�-M�_]v�mk�
�T���nȳ�i��Tq���,k>a�w9�%g`"J����+pnPM����M��v��XQ�]��v���sEl�Һ�9Y�w��v�A��)�9ϱgn]�*���T��1�u:{:����X�c��Ѫ����ݺ8�A�n���4z�2�����|��������Ag��=6e4*"s]�.��X�	�#vM�=kcA���+�B�x����6�4Զ�!�
�N_)��Xm�C�F��TK�OrRs:��*�oGB�/R3��v'Z�����;!�0��j�d0d�Gd
ݥC��z�9wT�L�[ݴ�v�)��Ur�07;#|�C�#@@Y�}��e�|ԛ{9Ū�c�0gf�w紷l���z�v���1�e��w��m
C:�B	Jl6?9�}^��Y@�tF�W�GC��8_�.%�du1�i�Ї���dK�k:/p������\�~�.��X��������J���+�º ��7��:F��ɮ��"j��E�GP��ԕ�%�H��Rvaŷy�K�n#-;�g�s��ꧪfɬ��\���|mIձ00��B!��eu�j��̑[\��[oTؠ�2�j�YMX��3���!:�q�N���!���,�+��E�s;̇]f��k�w��SH�!oW_v���Y/8������LҢ�;���o����������Wk�Ό�-NSD3:3�E� �<N��r��_��eED�N&~	텈0�вѬ��9�X�	�B������l�F�ޚ5�;B�����4��A���
�Va��eM�]���Y��T
K8�Mwlv���d�S��sOv��cBn1հL�9��2�eoc68��I.h:��l��T�Ff�`E���T&��E�]��By���+T��-���T�65ѕ��'g��M�c����ݹ8p�
x#���z@�3��O+�}J����)���GD�2�u��=f����iw;�7 >���ASL��u@o.Qї��bo�N��хz�0D�J������l0�
��ze9�<�[����E8�F�?��F��׉�r�
�P����p,����*2G<>��j�]�����b��p�M�k:2w�I�iPdu����SF��w�w8?A!��F���TV\ri������:�`�1����}6����|�	�:�(ݕ���tm�#�z�K]��ЉGo��Tle��p�w��oe	̇��6�M�Z��@��+�B�ݚ���{�@yG�.Q�2�~�OSy��&t1��z��|���l�Ո�o����z��L~��y�w�=�t�H6���f65������QW�-@f��f{+�S��yl�k���ّ�eleވg�bs��T4=����E���O��`M����6y��2��޸���E;��S=�觏l3���=ܘ���ǁ̨D��MQ;��f�Dx��RWcMϱ�Ĺ��΅PF�����)� ����Q��~���x���Eb�O�G$���ә�������4531�̣�;�nڛ�;g�T�w;���]>n� ��J�<����s��r�L̩3Vf�/z9��Ƃ>�1�'�
��D��XoJJǋ�X���)y.�>�B�@���ZA�͈�檈/z�[r]�A�W�^�g��r�P�e�5�lPO�z�gM=���U��u�b�*PAۂ�յ��M�p5�u�ʛ0䟿����;���(ӣ����Vt@����j�u�z^oRV�z��hR�	����Z�3�j�hm�V���;�]�ұ0Xg��9��s0���]b :�[NHk��[}���:z�N��]a����� 8m*��EÙչ�2ԩ�ֶ���1"6�I4��a��`�s]4��\d�D̍a�uG�6�b�t��^m;ڼ�jH��KV�<�y��NY;P$+,����w	�(m����
��j+Ǉ�V�.ck�#��H��K#���^�%ӌa9:�X29��]fh]�-'/Sn+��!z�W1���(�����[���<�i���]"����)�T�u�W�h�J����|�Z����b��'��8��;/N�]� �C����<nQ��RE��xT�YWU��Z��I�W�X�*������r�¾��d�ݥE� �Z-��eKՕ��Lח��d����ZI	��y�9�=N��_r�x`�<!ᚭ��>�p��-M��b�MNVaR��z������%ú�M�֪� u�7;9��ؐx�+���x��=wa��&#=W��syP��:蓭���Be%�W|5�A��� �_W	*��o�ì�E��)�:�UK�a}ϕs�`�f��_+1h���K/�����9'��Y�A�0ḻ��L�c��6�aܽ9�{�E�ed�,y�N��y�t�k��u��|1���=��'�z͹ۂ�/�V��ko�n{�w0�L��"�\��ه�0���\����y���*�k�NOP=�:]Bл:�^ i-гj`xG�6�dmc7��i�ζ��1���J�Zv8��7��n)�;L�;�����D�o���]X1�v��ڮ1գ�:vl+�pwN��t��JX��=!'@�|7���mL��	��O��8����;De���*�(�w����.uy��&\��\y:�5��v�N�zuH����+ٵs��U���\ t�˝�c�(���qv���ޱ k��U��m#��\zp"s.�����kL�^t�S��s���8��vUyA�ڼ�6M��]>̹�ʜ^K64���,t/Ǉ#o`�Nߣ�ĕ��lc�uoˎ:Z�2�6_z�Q�t8u�dy�2�npt���K��.gD�<�5�s�C�7�y�/qp��)�밽o,̗&n9���b�J����� �>]��;(`���ւ�f�J�s��W:�vQ��l@�+ed�N�bs��3__ܼ������yKR�g�e�Od}���=[&�JuD�e����d�)��L�,m���[T��X!�*���A��;�piZ�K��{�ή��S���$�4�k��A�����^Ts�aڌ)33SƬ/Z<����X}w;�*$��87�u�f�޽��9�q$� �e(��������y�{�������d�	t=F�H3�������}��o���>ߧ�����S��:�h���N�u4n�駛��)���`��?O�������}��o�����>!A�4�PU4:Ӥ5�;�Y)�OQԼ�.�4��QѰ�/V�ati�=Hh���#e��5CRtC��.��U4�^ :��7��Ju��K6�kKQZ�+u�CC@SMQ�� SB�f�j�q��Ā�|uuI��$���*�n��J
�4�j�����U��F�(�&Ѥ(
+����j��"�b�����j�*��J��4Q��'�
  UcD.o#��"D�1 ��8�&�����L���,;�z���v&�:�9~Q�����B��-�wLf���;Nr�֒gZ��/�K��qumon�M�H0f|�"����L5 	�Q�B5!M�P!|ᐘ"�.4����?���|���MUil�������
&B��(���(l��~V�>�t�YYB��^�cLV�5)��]]�)$bic{���]��s��aƱ�س�A|G�nN�3"�A����۲��-�
&��?��r����$�FD�#���E�w_=�V4���Yc�>��-�w�{ڲ��q���Ͷ��MS�ή���Dd�L�8A&�W퐖�'�8�ڋ��X7g[�j,�0fKd�QȚ�׃�������;�#a�Y�\�S��}}S�@�ǎX���v�wm�������K^_�d3��B��U�rD�i��\[�*�3;Oٽ��W�	�-�F!#Iz�Z����l�<�EL�n��7W�t������%�}��rL����>ͥ"���棜�"���wf/�)����LZ�(���y�����z�%�H9p���+5H9����ٓ��H�$�؄}Vo}³�F"W���ێ�I͋�:���9�3��{O�v8�f�ƛ�j4ͭ9\�E{.�qWWó6�Y͈F�A*�:Ϧ[b�����'Y�D}y�!׳D�	W+�e��hgJj������xm�.�C����jW0�B�V�u�)R��T�D�MK����N�=������s�V�V�:sR!>� t�0|���4���ۛ�eѹo�U�/��!�����F�9T�u˫� � ��ӃW-vX��:�v�x�A��>��οs�xּ�uu�3@��!e����T�m�o[�[C=�m�H�-\�yF�mr��`,���=���3u�W5�3�JqOe���
|��������K ��F
��.�� f���l1� �B�M���z����!�1cɄ���b}<��N{�����z[�(I]wL��$��e^�ڲru�S�7����3p+
���=A����o eT�&���7f��>���(T��۾��2`Ǜ�
�V��"��b�ר�nC��oguQ��TH~�/�v�Hcc��h�|	�:�Sڑ��ͫ�ikKO�w����̻�[��|�Y���ڑ���֡�I�TU;�4��+���`�Y�� ��k�`J̻�#��E%�����]9Yw[�:$���e�q�)�̊�^�
e�tHK��H�1/k�
슛nf���]��^o0�81,r���3zFR�<5HK��FGSyv@��;Y�4g�f��~�B��x�i��f�����ADA�x�ڡ��;�i��G�/t6"p6. `*�����̏Z$u_ҕ W��m�O�V�0�E�.)=��Y�'��g�.�e��hdŮK7���30�ɼ8ob�M�^�9���9f!���z��]H��x�� � �ߖZ:2WN�N���w[B��Y�'����2hA�F����/ M��0���&j����[{}D�����o�|]��%@�����S�n�vdH�1I��v܅�iV�k�HO�Ul1����2I.y��.2�[^��N^�[���b���l>b�2�L��lv5K�ق:+��k��t�^�+��+5��3M1hƈؗ�XM>kn͈��]�ϙ� ���]"s��J����J��ޛy�ikp���vc��ݶhk꽅.�1�Ѧޕx�c�!�Z�;Gen0Ц��NB��b�]�Cw+�q�$7��j7_O���PRB2��� U��2���f�,8�����dD�u�E�����>3+t����-��V7¤��s	�yz�;�~���{wo8I%�Gsz�{3H�g���\0Y�z�&�&NuմJ��͋�N;�_v�zUi�%n��,m��3`0��]1س�q��M�3��Kgp1�������sg��q�r�� u��AUBQG׹���~��J*��iq�;��%�'���;#���4�1â��k��kkލ�kOu��~���
�� U��z�A#�}� v	��3#�[�Qp�Y�:F�zU��P�O
���#{�ѻm;�H�H(tBT����x�n�7��_�KE���vȴ���zY"�P6w��Ą	����l��^]��n}�꩹�����)W�p�x�g�� �=ܘ�匃J�rѣGQy�����"k����W^=�*��3�΅PF�����b��Wf;ؕ���&#��,<�!b�P�H;w"��]k=�ߑ�nӧY뭛t�n��P��@��P��^��G�T͕�M�M�w�s��-WѨ��Z�Ԓфr�uM�Hj4g^Ԛ�)[��j�*g1twmm�5���p|s��*DX3�]�B1#V�	�s�7�ط�w�7��Y`������%�ɡ�7��﹬s�<��.*��t,RZаbˇ ��]\y'K 
�.��.�[X����;-�Hˏ;u�HɄ����7�%e�*�=�����sE��N�n��F��[!��5��2+c�5�����+��	Y�
��3n�vP9�u�vo�۲;o��lx0����
����9��y�ef;_�M���� C���uYD�\_�#1㭱��ل�?�4�SyX�xUR�����EE� �b����
�}�i���ڢ|��k�OR����S8���7;J_v��}�uyi5)�b�͌)Fԭg�V�f0�ږ4w��������T�ˊΥA�������(r�A����*�z�ht�z����v�.�a|��z���ѯ���*��{;6��{�#H��#�R��۞w�!�,��ť~�Nl�~���F����9d��7o���z�w}�;5c�_Pܘ�9�ݶ���R�ýr:=���e�|�\���������f��4+w^�=��]Ԧ!�S����5���Wpg�D=������>�ظ���94s�uވ��y�U&��LNo��$��;�9�,f������	/z�.�>���v�����^�uhH�%��j�-������� A�����'d9Mz%J�܅���!��<������L��LLK�x�h�.o!��'�A-vP3d��d��)�䂕q��㺨>c����x㾮��x��|�A����A�v�g��\�����^���:��:;�K1���`ޣ`�	�H�T��p�|�3mbQ��$��M4lt�ݞޛ>���*OUW�j �Z\�H_��m]9\�'v�
��O�	=��W� �JN9�^x�]�=�Y�6�B�nK���з�/U�kGуb�:}���Z��erM�g>vB����8�tN4ш�ewO���0�#��D-�����9��������
�����	�u@���/���m�ɶl��Ɩ�<�z"�/m۴#���k���*��Y��~Z:�Y�K�OwGr�;�:���l`^0�]	/�gΰ��38Eő�V0W`�i��Q��k%S���.LpN:��9I���E���ؼ������hЉI���W��?������{�o�|�A�a�K��.��L�{�����Kt�m���w;�k����%���09*O[�����W��$r:�is��x�d跤�!U�3c#�{,�Ҫ�l��3XXw�H�0��6u���Ee��G\�M��a=E�R#���d�A�;h汁TD�#�`��	{l�:r'E�V��7��_Y����ᧉ|EM�3��m�c\�ɜi�zj;(��	G���0�� ��7�2��� ��-�v��������B"�"dE(v�z&��/�|:�|GJT�S�2�n��̼��Y��܌�,�F[���z���<�&)r[���q;,����s��i�Sj1$u�M�Q.�nL�@�=>�$����>��g�~����bf��)�fW��&�uU̑�OL�@�(7j+n.�CZȬkq���&^���`M�P�[';�8[������O}�s�#(�ꠡl�z��/���&PWD��q��L���'-J4�1 J��y�*�X���/�o��g$����5�V�=���ב�r���)��(����;����\�u[�'߼<=��v�l�[\�"6���E"Η
)�T`�W��O�-��fž��<��v��*���!9~�F�f�G�"u���M�[������3U}���ę+���m�����L�Z@�|[@���T�:��	���šx~ܾ��J���ߣ�����Y4~��ϼ��R�16�_%����k�ܱ6�w_\ѽ='yԅ��l��,����^�R�����)��-8�+t��wv�q��]��(�*bou½��.6������č�L����+8u�n�w��W7+�Ք8�R�+���a������wL##C��~�/�c���q���|�g$h'麟.��ov铀�c�ne��y9:�-c��v�,k?�<4 %V�b�D������4�[�a/x��ҷ��d�y�Q�k��iu'  ��W��EAi�V�u���˺����px�Nx��L� u�px�\�;ڊ@pU�V�Ņw�m���;]�G1H��\�CN|i�	Y�7y�8y*]Η
)).�=�i���l�9�8D�R#��������q;��u��GOow*�nU�����C
���MU�Oi��V�,�k�j�{w�<���ۢ�^O��[s��0c(a�>��'���Ӣ�{o��L{��ው{7�A�ΐ8�{�^JΊx����V%��sH4C��CF]Y�wVwt�����i�	Wf@+�]��)M������5�[{7�p��h�ّk�W�K�� �ƧɈ�r@)6dנ�Hn�"�MI~���'��{���s���U?1�Tܺ"1v�XQ����h�ʀ��])��܌���Y��M0 +%�J�{|gzRW��EC�D�͗��t�gc����ҩ��|�N�k8/M����!H����&X5G;���A��'N�u$3���^v�m��m�� EA���ӗ��s=��o��E��آ���X��?}����M�>���O����f/[U؛4�s��A���j@w�|�wخg�tH�����kO��`��j8Bb3Q�Û�{�*��s[��a,V��y�Q*���:ѳn�}~���s��'��k�c�Z��G
:����I��ʰ�dh��P�Y����؃�U��{��fL���S�R���*�0��0��':�
��u�@��O�ؕ6��s����5z�a��Z�/�W��W��K���3b����g|[*C�{o��.D��~3/��������r���ps�����y��Xb7�u�+���G�z�*:_���52u����r��*h_�����!&��qX_&��U36����FV�9�wV!�7$����:�l;���gVn-*5;�F�����o��ݚ�f�L�%>$���(�ا��3�A��&u��\���m�����]غ��;}5'e�I�u��%��>�`���ḽu6!<���ZȖ��D��S��܅�	�Cd�F�G[6Tz�6jUso^�d�fb�6�^�3�"�(��2fɯ=ˉ��Sͩ*�{=��4vk���V��Y��%s���/��ّY�S��	\ؓ��ڤ\-���K��#�3��Cs���z���Iʫ�n�������B�W�����;&F�tR���-[�U�5Uep���]�9H%/H��
��)�n�3c��t�N���-��鼻�.Cu\�\s��*��;l�M�ȝ^�\��r�kZ+q(Y}��)ҧ�j�x���1�_8^�L�iH���'!��N���D`���݊"�N�@�@R�v�/
I�OWfl���vWJ�ǅ�%KXPA�\��]<�ϳ��3�>��@��Ӻ����&kk;���Vحb	,���3�=����卥�{}�1{�^�\/i��Dw{0\�4�0�u��{t�md8�N�0g.l���[�scn�]�񯛵TZ$���H�,Y%.ۮH\)��£�\{�v;����QP���83�v3Zp����ٸGv�гR�])�V,�삊b���p�tv��+cZ��ǲ�M�&�&�owq:.-�9�V6�OU���]�pީ�+���B�g��[���9��(����s�<&�ڪ��
�Mv���L�!��mM̓xf��e���v�&��r�Y	��¥Hdm�U8["�*ef��L�:F{��&�>��X���\7���M@�۔��W�^m�t������;�7��x�f���d؉Y�a���"��1(d��K��or�-�Kp�`="�)%��Bp�[]Y2
Ɉ9xf��3�0f.��_� ]#�]Vv�̢d�6��uY�p���jfMȩ��.y��ʃ/:ĺnqz��Y�q���Ѿ�$p�P�Uy�%3�r�@�a=��U��U`D��wK7Z��2�u�i~����}π��5p�:��;�?jE�a7������6	�ꮽ��jd��̔���5+���t_U�����S��2���N�I/r��y���iP�ߓv�ŘwEf�?i�*/�bK:�S�l�3gb���_-<�\�V&2K�l3 ���t���:2�*E9�Z�`����V�^;'3Pc�Lha^v�k�����c���V����y�`��X�J�$���ҳ��5tfg,��J�4,�+����WInW��&P�ür��"��L�R�t�����5{kұ����bL���1��Y�0��������r�]��kF��n���E�*s��R�W]�r�x����f��ե�`�6/l@�6��؋�[u����\��^6�f��J��X^����<ݝw�٬��Hn���TĮ���g0�{FI���Y��Ɩ�C�+cś\��@��8	Ӑ^E�]NY{�ܜT!�5�Bu�y�(�)]aCK�.�WtW0�is+�x�~*he��K�r��m�y��g�̣p���z�ُ!I�/�����VY�%�u4���+b�Ő�t��Q����Δ���w���Y�6��ٮ	f�PJ�MY;q�Ӡ�N��(e"�7�a�{�����f�Г��2;r�κB��b���������&a���t��'��Q����+Z�cSMICs:*&�<����|>�>�o�����}�O����D��u��]Ͱuj"��:��΂���5��'m�4A%'O�����}��o�����~?���rU	HD4�#�|�"'�f�Bb��(�u� ��g���? �TACy�Rt�4LTy�DE�4��f"������*����!��
��B-��*�&!�*"h����b
���b*
+F�jf�h���(��A��"65-�j/8�b�LT4EK�jO86��f��l��EGV��ƏQ����������^0b�J�;5$M��j����*z�&"���[�EUU]mT�TG���((����<N�(�`b�����
���������(��1�j�)��������Uz/]|�ѹ�0��c5\X��S�hR�a�Lq�u1�w���U��s�4�?پj��Oq���q+ǣ�����5�/�8b: 7W�����z����U�ڎ�u�`�HW��.�y[�&��q�(qA)��}�)o:�Z����=�Cc�>݉1I�t�YՕT�*��P�%L�l)�m����L z�+	�<�_$vJr	m��Y�����޻���l?S�����r�k�XR:�ؕ�b�|�����[�W���ó!��|�6���猈�Sk�OOD�䦘O[�K�p}4���3�hg�����'��v���
/�u��t\q�ל/.�FCbǷ����ǺlA� d��m���t����E�vgS9���Xٖz�_�Y�/I�/���<c��hϺ��m�~U+�SU@���k�yt�1��ME��}fOGOp�>�^�2:�ͭ�m���ַ�A>��W�h���\����dz�/j֍�ײ���;/qҍJ.Y��Z��"��v�׻�jP��l)D�g{4�|�u��S�����3��D�oa��T�f�<<z�l=�^R�^�;�;����v��)#���_��#c�s���bx0�9����4jkX��;:��t�N_�|�o^��$���/����5���h�M�g�r��#�(��Q��7p��T�fh5� �]�*�S��g����%�y�3g�&*���LM��Y�y0\wzqy{w���&�(��Ok?�V�?0�R|���	 �Ugپ����ˣ�	�YC� ɳ&�U@�gD�ul�����ك+,�J���o@f����I+a*7�.L�)P�ꝺ߄�g��y0�\�?C-���P�R��)��F���ow�(-�-h�丫Zpo�� c�r�O8�Gw|+�����F@r�}l
�*��e���U�����ѓ��v�?\�3��ɔ�~H?����z�%�ڄ�<��9���UK�z]�7;����~\�����A�a~ܕ����Ğ�m9~�N�v5��޷9w8�"/�z�n��ܢ�nʽ��6ϐhf���v?�;�*�e[�9�tL�%�3$��.��Vl�K\������nN�y۹�-�[/F!|��U�S����dG���9��Ћḙ�G3$�����8�2��9}W]ʲ�B�[ݽ
���Ċ];�B�x���TT{2v��L����|�xTbt�-��|!�칾^�ԩɹ=�(q^�nA?w�����=�uN��Z��R�?���������Q7��6#�5��7��7�"��8�ٚvg߆���7�S�E���� _?�%��l�/Q�&L�#�3���k�[�9fk�]��C�~ɔ�t1>�e�Q��F�Y����՚ɬ�������޹���\$Q�tI�P5��o��1B�RWW]*��E���uF��z�������ol�M>=ɦ򔎊}v�݈%�t#p�7t�#��o�����1��ۃ�i�c��̂�o)M�9�l�T>�ۅ�����ʘ�1}"����hv����(�J��*���Ϻ��;��9ƿH�:��$R��~�mK�&�:"<��]��)����"0k��z]8_9��m�!��v�`M2�H{��Ʉ���d!=�O����<��3L~;JE��,J!ǘw�}W��2c WM��^�+v'��ׁ�Z�k���
�|d���%;���!́N-v�K�&�i��f�$'���g�l�c���C��{M�B�Q�W�(�^7�t&%��Z��w�}_Wݽ ��{������3�<U��k�R5����[S�EpN�X��L��>vWF����z��������J���1m��� �,̋ɴ5\F�^E�s�+s�
�U<�V�����>���&��+��38�4�V�y�{/]'g�����f3WP�*�J14��������f��l���{�CdN���ެ�>���Pp��Da�z6T��uw%�1ҘK[�F����v�骱�pER�4|�
��8���gR����Wכ�i�&���ݨE����:CnsPm�!�?Z�p+᝔�̴�vZ��(�L~�Mޯ_���9o>�oOPgY�������Y�`�;b�m]��q���]0��_����Ykǻz��=�� hsϩ�7e�oY�ks�۝!��֥QW=B���_�I�D�z}{�Ekdz���?Z�Hz8*��]:�=�fb�að��^~�����4����һew�/��Ƚ�Q<6_;Ԡ�Y�l9[1�8m'�q��̮5����<
a�=}Ii�������UuL��}���_��W��>p�f�r������5�w�q-�=B��s�+��߭�qzު�M�׀�g���y�T���PW�023*����&6B���m���Y�26o��܋�~�x"�1wU�K�)4#�`���Vu�d�-�'���m�ݮv?'~�o>k�)T!���F�\!L-��
cU�n|�UL�z�+�Ncd�Ȍ݈��|nl~&���{��Y�EUځ�N��_��Kޘg�{f��']�K0|���oJ���ЍPמ�uO�3jQhys�o<�;�=�5��t�!�[Ek�z�Tr�R�PY� d��T����c�NF�ݛ�����;0�-��oO��hz��֟��R1kn��4i6&��DwTbǁ�ٸ�|7�0F�r��z��;n��MK*��
��83��F�k՝�O)�rv�>y��ހ�+`�2���_Nݫ�ZN�΁��+������C*Y�O�]9�ι�##Θ볔�ȗT���*��(�PN�˜U��m�ndS�6��w�]�&_�g�L�k}���_iC%�1��C�&�WB��F �+����dNb�\�񌫼�9|㣷��G��y�z����gzϤ���W�j���T ��6GPn��w�T�c�v*$;e�ޯC15�0_%Ŷ�Gl�v�Hcc���@�#��k����`Ϟr8@c[^��f��Q>=�4��^�<n��XSX��Sܥ���v�0�Dy0�Rjѿf� fYy������W�ѵ�����f��w;�Yy�N�CX52�37�ͻ�nG�;OR݈p�}m�ë��z]��X�������WP[U�0��`��$�Q�2�z���˯�ߺ��/o$�A����B�S%�GZAꊉs����	����v�Rfם^�z��ة"�����rux����>�=�1����x�mv�ɐ��Izb��Ŏ� ��ZN���@�(���4�*b5���-C?�%�N�g���|3^�pC'�B�mv��(�$���6����L���)2+#���]^�Ff��NE�zo�%�9�f��wKi����Xwku;�������}����8�����{O���2d�T�$�-ǘ}o��:5�8Ã5��ړ6LY]ɤؗ�n�snaY��j��;v��'Q+~��}_�)��[3˲LW.�au6di��LGӍn���A�����?v#���*�|Zt�7T�6jF\S�vذ�9�u�t���;=!�;K�
����Ӷ{$��b6i��;u�,������y�H׊�;εCO�v6@a���kIY��s!�-{b8���n}M�yP�ܢ���u��L�3A<x�)���Kwc����i��4��M�=���+���Y�Et�M�B��نq�=�ǆqӹL���[�PẜM�*�rF�~������Vo�n��q�6�U��n_��V]Pn���1��� %V�`V"h'&�2{;fU]eL;�Fȁ�$Ϋs#���,�£QV����N�g��ض�?����|��S??|�ߢ�	�â��6)�s���,�%e�W@jk�Tq������^�ؼHD�FH�������>�I�=dۧݍ47`�ڶ?fnZ���:�X�'��,���P4�+a��"�6vV�}��b�}Fi��Xkm���;�o*dM��u4Ɩ�j�0�=�8�vR2o;�6Sĝ�VL<���w����}��Qq�є��7Uu�:7tT6����<���ӧe��2�G����s��%���<��&�ˀw��uK-H]��/)H4��������3��W���%�Y�t�P�Sl&q������0��U ����<�4�\�r���xލ$�Hnۋ������d��!v"�t��
�B��h���h7�Y�X�v�B7:���F���H�vL�#ks���"�3��Ý��F���n�^�?qg��L�����m85��$'�����ҫc	�����V��L����}h�/=6���v�C�jA�-�G%8�]N!����q������=e6�+^F�:�����Qy`u��X�f�p�֟ze�Ǎ���
�a��vz�̔������%�)g��vM�Fv�H�y��y|�`c���(�S��R���ܖ�Lć旷Ƹk~�H�a�<��O��I����p�=>oz(����������ւef�Nq���/-,��B�����|�k�H(���2�Cp��2��cnN��v ]-u�wǧ��)6-Е�p=E�������]���Aky��xw��k[UW�\�v��W	řB���YWŵ9�GDʔ��L��x�n�f�̋[�m/w��rN��Ɍ�؆✠�@=#�6�sh�!�f��x��˵Tqq�[�y�S��������]²w�{D������T���f�o*�e�G�����ȼl��Q1���H;}��|��]UZ�΅���d�:5��W���:%TUʫ��]wzkx�QX��K�e.�����~}�y��MPȎ��ڨ��s��܁�! WJ@�J'���csW;�Xr{���VM�n�PUv��s*l���\B�ȃoJ�U�����9���(��2I�U�ד趧2(2
�P����v�����z+ w�֍�n��4�1W�)F�)J�R�^�e��u>�g�Sp� �Μ{�暣��[k@�v�ZuS�hs��*O�6�F��w�g�us�R�)eF�OA��܇�}�n�%=��7�%|�y����=�l���ۥ��`Ǌ��;x�u5���\������U/�V7b�tUצ,�v-��pc���g�Z�^������G�6�c�R��kgd��`����Y��;�5���n���t�K�Κ�+0�fp�j`�PM���z&q��(~�g�rw��qu��K�B��C:k���4W���\�n]�����y����K�Ҥ�'�B���>�[1�=|�GZأm���Ɍ�t7So7�QP��J�r�;mhfߘ.�\]�X�5�Հ�Nt*ѻ��yv�q��G@��*���a��3`��F�iLV76�� ��?4�FҺ�Y\���Rv<rFO��m�o�m�y/����hH���M��.|�j�f��rR[��v�Dws
c��h��z��CCDZf��Fz/��cY�s��mB)W�Ӿ���v��{>riJ#je�������w���Q�l��!<��� xJ^i��ck�>�p^��p3Fٰ�L�Gt<;�ڽ����s��|B�]��&�w���G��������M=��14��UcP&�I��S�4����P�A0�S������~K?���+��""��?�������� �>O[�d&VV@�!�a�a�dB �@ `B�!�a� !�d@��a�eXdBV�U�!�aP!�eV@�!�e`��a� !�a �!�a��P!�a@���A��A��qa�a�a�a�a�a�a�a�a�`a`ddXdd`XdadFFF���A�A���A�A�ב����� Ȁ�Ȁ`@`@d@a@e e@`@9���(��( �]� 2�0�2 20��* C  C" C �l&�@Pi�S�TS���T �E �eD	�T@� Fi�aVfeV`���A�p��3��,2	�M2	4�$22L(LL�u�@�C
�0�D0�0���C`r�2��Cʰ0��C*� ��z���Pc����D&PRd���|�/��������_�������������������o	�������~�ވ������������"(
��QX��/�?�>��@�)�������?zވ���'�O�����zH��ܞ��?�?�N��O��}�+�eTQER�P�T��IWJ�� L�0�� B� R  , ,�,(H�$	(B�# B(B���)��K2��HJ,�@B����A�
:?@��������?��R� �@(P��7�O���/��
��� �����(�����?O�����Oa�؟��x�G��{c�����"*���C�'���~����*�������?��"�����^�UE}��������>�;��C?)�G��|@x�"�+~�?���ETW���v��������?�������	?��������?�?��"*�����c���
Oֿ�D��`X;O������I�a'���"�+�=U2{�i�'H�<���A�;_���_Ԣ(
�#����DP���<�y��!����(+$�k)�� 
�0
 ��d��F�|��kki3��1J��J�mj�`Qi��UfY�@d�,k`�ZY����ڰ5��Mj��2��U�m�k[�����[b�5�ͥ�lƯu���[kZ#L��i�6Ս�+b؋,��jc	�YUM,3j�fְ�eۺ�hI�(ږ�LIL[R�n���h�k6��k6��r�m�%�m�E��ղ��ɰ�3��ѕ�EjiMm��1Q[ɣX�di6i5���JhT�նږ
mm���6��m�,���ijٛ-�ݍd56լg�  ;��y��9K�]�*��L��[�P֕�r��_{=�=�2����zi:���۪��w;��	��z3�������δ:jL֖à)۩6�#T�ɖ�l͋X�gq��  �B��
Ƕ>��=CB�
(�����(P�
47}��B�ǽ��|����'Z�-�;�u��Y��F۵�nU��*u7E 4���[S.���Z�p���kl���[dUV�kW��x5��j�ic�vv��0��:���;�Ju���gp0u�hiY������T�=���R=���Yԫn�S�a�����U�Wn��Mm��FQ�[X�ZY��[m5��| }����mn�݇w��{�4�Ght�Z7:��� ݆e���5nU��.�n�PSg.�	;J�@�Zj
��"u��Y�3am5T��5��۽6)�#U�����C�r������v��3;�N���q�V
j�wu�v��\� m�q�n;�2N�6��ؕ�����(�Y�x#ޚ=u�vi�B�uX9�h7N�Z�(0�p�EGn���N��Z�n͸w����� ���l w3F��$���CFm�ٵ3o���kFZ�[��]�tN�
κv���Uwm]���x� �������)��iׯ=PQ���(�)^{ӏ*F��y��$�kk!������ �>�����^��t2��*��/B�!<xnJ�*T��;���QX;�yW�������Qk�[�HN��ԛ�IJ*��<R�l{�mԛk6��M��e�UD�  X��R�����ut%���z��W�zܽ���Ha�ӹC*U��{�
P�u���R�J�x��m����s�Į�l7�ޞ��O`e*��k(�lm�����zs��_  �ϧ��J���;�@Ξ���	*����޵��=w�*����A$U��U.�)'=y�HT��y�w�!���w�w�A�����R�D�@ Oh�JR�  )��	J��#@S�����   j�Șj�P�����U  �5??��?� �����uD���B��,�A��2>����r;���������DO�� "+�(*��� +��U_�PE��"+ ��)��?{��u�ғ�ߕnX��)�w�<p�E��*1V��q��o(�i#�ӟ-P�Z���e�.7[0e�vܫ'�D���$��kr84J���VYRب���3�K+Z���5{��(��[��0e\����3�tZY��۰(�d[i�bP�䤆���n�V@i�*��3d2+�f�d��U{_�xU�F��������BM�H�ٽ��E;z��M�`̣F8m`�0�I�MK��
O*�,V���gA�^�С�N���ֽ�����Ȓ�������N]D��A�I�u��*N�.�t�T«X���Z�ԧYH25"Mf1�m����lS���3X����˫N��<&���&�mՑR���P�RՑ�p��7f+��̓�Yp7��1h�n�"5�4����1Q���h� ;QJ��wFiж�H")��nM�
��h��J{mN-u�4�7Tj�����L�1e��(nf�f`�R�5>z��r�iB�F��UK%��V>�t¦�Rw�Ul��h]��7\y!Q�n�U��Y��&1ySC�$����a�a�ٙ��0j�4m\O�R�O>v����lJQ%�Fj��I����bC�d�.�D�v��XX*,������ͱ6Tp��MZj�w��v��[��*ڂ��n�@C+H{�`yA���64_�kmd�C�q�[W@��ּ�E�[[WK������{�^�'-|�k@��1y��:��/e���`�.*��"���|iG�)aY
5��ӲRԶ�[�3zݽ��M�t�3SX%�L\�nʕ�j��X֬f�#��h�溄_��J�(���e�01yA��U$NcMq֚��*�V��\D9m���!��wB��i,���`'"���7F�c�)<jEa�H"��tjc��Bkj�U�xUBN�"q[& ��繂�u4�u͸����|�Q� �unA@4lt��Xm]!>b��۰�ޅ�����I5�&^6�+�l�KXu���h�=2�x�ܛwt��z@�%[����&�U!��n�G43���1�z�@�hCa�����*��}������J�=[i�2mU��:5tM�g-
LU�ԏe�YU-�¥^�)�Em1�/���a���i7w�U+��Dd�0��
���%�!��#�o"%��2$�rZhY
��K���N�B�52�<,�гX6�h*�&�1��B��Ym��ofN���m-����t圫���X+U�ޛM�SI�j�W5-�-6��li:�+�v���B4)5y+:ɲ�)����8.���I�6�kt`�E�U�z��Qҥ�f�8�m�,f�v�KL��W��㻆���
�q��;#�ӥ��5�e���2誀���`�J�l;�.�m,�7v���%-�Q��!�($�tl�*2SYkX�LД�[���rX��h�>n�B��w�Y]VlX;3Z���rM�B�yrJBE�Uj��x"W0@q)	���	LC� 2���wZ+%*u��Bk��kr�Aql�A2���t�q����x��%�lӰ�t'��7mY�)|"���^iߡ��"�7&Q��ZT���M�[k5�ՀV',e)W��N۴̲�6Ŭ�)8T���ܭ�6�	��݆JS�k%�C~Ʉ��L(� ��2R'N<��7��M7i�Q$�e,)�T3+�q�I��vEM��dVd;�� Өn�Y9��dJ�1`[u�n��[�r�!Ҳ��a��2�f�["v��sJ�g�`"DF^mjR����'��Hg4��y���j���ذ��v�L&H��B��A�8f��µA��a��40krȷ]���՜�+�t*�,�$R���%�GYx�8Vj��R��*CY(3u#�O3"F�[��9��A�I��Q�W�E�~bP�v���ހY��4��E�O�2ʊ[�-���ou�ʷR�9������a��6ㄣ2�ۭ�L�!�y������ۊl	T��{U ��aZ��R�k$��j��ӥk[[saJ���]�ƕ���(�rD���m�1T�֬��Qr���e�Bd��L�Z�vь���nRŊ�����Q�r���x��tS[X $j��Nl/*��h�m7���޵h$�QV��kDAC��m�]��nù+3~�e�_t��O���hX*dk�-�X���Έ��4�q8v7��	u�ܤ)ň��un(ذ�d���5�FÍ���ݢM]䈷x&áţV�f�eXH+�2U�"�x��Z
��zf`x6��W��M7%n���2�+��!�W��u�y(�m!r�B�3>a�;Y�a���
	��(��%E���ܔ2�6�j�P���Y�ݦ�P�T��^��C'Y��a���o��1*��Hva؎j�r#�m��W�T!ۙ��)�sH��˧6�;QFK�T^Ҙ���!�XTa��)R*�R(������ɨ՛*��Z�ց�0Vkݰ�:������^nmf]�Q0�fVV�*�+S̅`��5�U[�ʳg�1Mc]�]V
��.h�D8�͡�t�(�TMYctѩ9m�����Qf��٭�57�[�{�*��-a��Op���p<�Rf�� !�N`zX:N,�qcV���j��o.&�{�nȔU�u��h���5ux�u� Ε>�0޵J� ��Z��`PA�T^�\��E*��QQa�j֗F�{@�f��B�G[b��e7B�M]=B��"%�� A�eT���P��pVK�Q�Qͩ�֝Zѕ�j�G���uX�
*��+V]l�2b�)0��B��uÌ���(jEt���u�:ۺ5*҄�]i�Q�4�a	n��6���:�K�n�kD�Z�Xhm�M��Npؚ�Fn4��1�bv]�p���Cj�Xʈֶ��a�7j�7�e�-4�@�YBkU#�g0��dz��.�yd���g 2��^��� �����_��4���%���k���l��8�����حB4T��nZV�����@�/q���dX���Lk��kc��#!���Ӕ�5���q�h�s5n]�t��[�C�C�����[r�e����*�T��Ȃ^մ��e�jZz�m�%�Ôi���4�'��x�5���K f�,�2P�	n�A�9�[R����]������i���:"x��7Gp+�Lޚ���Lj6��D6Խ+P� �[�į6��.ن�bm��h݌r��s��hۦ@�����񁅡*e�#ܣI��6Z�(���1�ŉQ� Ҭ��ʹ�QJ��xY���uh����;kEK`�y�S�[�|?+�ځ]�r��COۄ��<�̗�e��"($ �����J<S6U�ꨩ$b�K��M����r�5peIM��W�^葜ǋ1��[@�{��bۆ��LBi rӛe#���0��ˢ�f�q�ޛ+"������Z�Q�b�lAN���8��˕.��B�$割� �Y��P�7&��7��X�`Y�܉T5�srj#`�!o(vEc��^L3�ҩdg1�e������P��7K��LШE���6ٷV��B�s+d��#[ˈ�{ZQ&�4�Co/)��NF"J+�6S��hM�ɷ>ܹu7rΝ��5����:��I�:-
N����]�#2�dȠ*�y��6
��E��oV�Ǻ����4�f`�w�ZT��K�"�j��C�eF4����E{	��s2�z��"���9�h`gYze|
!�	�8[̚4�"���P[:���SF}�eӆnR�+;K��c:�T��.��{(�7 ��Dc-\1�3i���j<M*f�a���� Ɔđv��`�v/H�jU�ԧ���0�Y2H%��;Ն�X��m��p�hƌзX��U�� �݈.��$�C�[6�&����N�CT�n�M�EC�h��r��j��n�M09��n
��ٲ���������32cN�R���}hi�RX�	u���Ӓ�Ĕ����`k)k����J,7u�aRj@�֫ځV�36D{am��f܊;��4��3.�	��i��i伋&�$`��!ѧ̫�)Uے-�
�[)ɚ4�qse�T�gp:EPe
.�cF�����'딋R�����4��/,�Һ}BSt������o�
͒����K�7&�6I��Xؕ��r��wD�2�M���x�`�lK��,�V�zF�d[B�^嚄���fd�7(��^���uַ��i���	��Ei#m�	n�t�Ւ2���Gq1s࿎�Y{P�l-7WdG��&5تڲnnH���8�i"[���w��n�l\͉�`�t�U8����i%٫v�$���i�&l�P��Pݷ(��l;4�]�$�32��C%�Թ6I�u�1<��i�:՚����V�����a�`�P&��� �r��Wf��t�j�F�'���7�� Э�/h����uXAʵ��SO�i�M �m�kZ\�7J��8r�\�:�?,p�
Ԫ�1��L�;[g(�Gj�EL ˱1��ĸ��Oȕ���鲒����+��tm����x��q#Ku�.�����ы);E��o*&�..m��g+p뽁m�%�r�QCg/^���(L!݊T�׀V6��ʥ����SwtV *ͳK2%d�ݡ����D���	M�V(�͢H�P˪9r����p����	��
�)!�ץ��˸/���/e#yT�[�1r�6cr;�t!�kl�mL��#++	`\��*T������N�70j�1��@m�Ԇ�F�悢��ܧ(� *�@U�3X�ڻ�H���QF	̹BrI �$	]4�/EԲ�i�
V	�Ypjj1\���5cS)��{).�X��hE*�G������'u(Yf��+5W���L=Rdʈ0&)��$h��x(��m�A<�=���R�4V�Tr�ŋ�{i�z�V0�3U�7 ���{�oѸX
W��=uw�VVE �@�3XAY��#a��w[M����"�f�5��HK���Fh�g ���k,Ef�� "jn��A�������*vs`g�7VT@��� K\7Sd����m]�e-�-���X-c����-T�T��U&�y�am`]���MQ��T��;pjۇ^d��dT�5*%f�8H�Jm�t�b������!)@�<Bm^V�Fn��Qh:�ֳ�tt�Z5�\X�h8"7���k^�4�Rbe��K�k[�D�+Z;�,��̦�Y۬J�d1�n7`�U-[V�`��oD��,��5�IW����S�Ȓ�߰h�#RJ���Y�D[Ķ���f�S���FC[�֐�x���E鬗L]�"#��8ls�Ud��0P4��0U끚���r��sj�)�X�W��T�!N�B"d��_\��x����h=��J�0�iEo]E�1!���ćKSt,ڱ 1�2�keR��kE�+��r(���SA�R;C(���x�� f��S�`�&Fa1`O֐�K(ZoZ��.X
�)ە4^ҕ�v�En++]�3
#�Yl�b�i$��,je���������Ō3@��ju*j�{�)��`+����5��쥘)�Yj����֙	� �Q�nfXZ����Zd�*8v�M��+5�[��bf��j�U��u�2�4�v�T�0V�DK�"'���jh��g*ٳM�ڙ�wY�j�Mib�����%�㄄�] �&�x(n�6�35J���"�V�"G[ ��Ԕ�y��Yn�f�ٷ��O �K���l�Ԭ?7%$�Y���3�ن�ɇh��T��t���rf��J��P�Z� ��-l�e�)R�Z_^��(n�ۥ���P;�-�p鎊���Ij5�(�xh2r�ۙ% ��	.	PEK�m������aM�����u���v�c�ȳ�:a�ݤܹ�K��ѥJ�L��`r=.k��X&�^,[��*�䎁{\%^���7p�i}���Ra�R�zM^݆,$�&VC�Lt^�N�D��i�j}�u�0cĚX��2� ;�DX���k@7$^��P嵭�J�l	.ݕ��-[�@� "Fv�nVǪ��5iN,`GA�����rm������Q�M�I�KF���z��W��l�@Q{�k�'e*2��Am�YZm��C,�ܤ�܍\1��<uv�R����V���B}(YOka�z�=PU�ɸ�d�� ��MHr��{�oB�5�c:�ĞV�F�!�V�x�ܩ�>SlMv*ʅe8�����3]�%=�vhJ/vR����m�q}�L�YA�J4���N�(ꩭ&�T�/��Ֆԭ�m��yp8���5o[��Ա����/Y�D#�90��Ik�kufĻ	���,w�n;���5{��*��I�O�t\:&�2���!��Q��d�WM�(�5e�l`;��;��S�rYTV�jUŇd���n|7E�6�e�!m�0���^�J(E�	�^p)�Ir64���h����n��,D��z��
�H���(��`]#LZT0�؍��һ��8�\��9PVb�ŢK#e�vօ@13 ��xbp����l�"��(m�z�]Kwl�EL
�1�M˷��Q�&ԸI՗��E�P`��t�v�/���Z��n�e�Xȉb�w`�g&�t�2�,[R��2Z��r������:	,��*��
2ںf )����MnSoJ۹e�n�N����Q����q���tԩ?�_�aRW�kvKS��P=�yP	�a�L�@v͆�7
�� C���ya�1GC���i��=�J�k���:�b���󱮇�hT�U���*1�ҝ�u���j+��*��Mj`�j��Kn��J���Z���O\X����|Ʊ�$L�����a��� �o�X�����}��֖�+��yz��^���4���	�y�SS���I�+N:{)����6�c"��M��C��mQ=EuI�i�\��^ڽ�0d�@��8j�K����cpԓM�x	,��j,vp�@��U�a]K�E�K�Q��T��d�w�˕}�u�E���'�]�c5��vK��lC"	%*8p�+�\��c�5D�sdҭ0A�!��t՛�c��rgW����j����.u�g��t�]M)�4��%��C�;�]E���\�t!��0�veCu�J������9���f���3Z!U���J�[��j�96��I�T�.8��RL���v�%!�i�
�MP+�+�n�\D�4����O�&�Z�����t��v��u�:8�],T�v��%K���3H��F1����\�S�fmU�����Y�)�����U(V��mC��͑�W��s����!;#�4��S|�&�f	�Q�i�;w��ͬ;J�e�[�,Hf#���`���<�۔��u�^�MDr��L�J����P̊[
B�'Z�YQ�1����d�Mۛ�8�L��4����J|�4�I�c�밓���a�S�دr���Xù�J�\�8�R�*��z��O�=\�,/��f))�[��ūE�6�����8�Oz�3�m�B0R�^<����srt'8��j��9�1�kz���`[�V�#�vr����u.}��"� �� ]$fzj��K�u�Ŭ�����@�証�TA�C<��� YTH�7��)�Hp+����S�N�I#��R���:me�ϲ��`���ؤ�v	��d��ڏ0WVh���A��Q���KT����Q#E~�U�����
{gx�aN��4��:RY1�r����l�]�2:K	�����};j�t0��S�iK;�9�͕̀}�e^�ףiݼ�g0ws%G��fԳ�����qK�gv'*lӑ��F�-C-�!�w.��Q� ��G+��M��ۖ7�ھ���VS�F��Z�;�),Uty^���b��-���Fi�ʜn��C��ޫ�.�����Y����`έ���v�9Ú�P�=rg'RaJN��`K�-�|�u0=t�;޻]�0��/ 
��Z�5s{ulH>5.����r�=2����f�p'	p�+�⛶�6v�;�s���Լ]6-�Fd���+Y�x��xDm9l�F%�s��3K&�o.]� v��Z��X�VҷM|S��ե���7¦�c�@�����o�$�.u��R�%���g��J�!�hP���g�lP��'B�;��3@x9Q΀Nw����N����h�+cX{pf�:�ki��̹]0[:�z�Λ/��]d�¢����`t�ݛ/A��H̖��*ƨ�
�Cr�^� Z��ݥ0KkFf�f��L二�Jn�I�uj�r�x��p�,ҺN8:,-Yhl�O�xU3��t�\�-�K2�VS�%���DYY���|p����b��wbd>�b�H�3���nʝ�6���U�^�ي���(]�]Y-d�c-!���;#%�Ź�qȈ�Ch�T4��³ �iֿ¼������z!�E�on��J�K��)՗��Bi��8�b��3*;��uةp�����uщ+w����Nd
��r��;��9WFk����m^�S���^�jj�Z��]Y�n���bk�T�}.�wk��u�ứ�1Va����K5�`���\�i�\�H�˧F�*K5)���MՇ �u(�K�&�yXG��ռOJw�a�]���)S���ZZ`�ӧvs���-�0n�Dc���b۳G���d
KM�M�����PM��T3r.��9v�9��-�mc��
a�ʶ}�	9eY��۳�ީ/�9gv$5�`��6�|��x�J�������m�e.�[�}�UL�1�Y(�T�����Y��öf!����[1��1�$��B����jʱ�GR���1c�;���9n���`���WVPj��}�Y�"�{OT��@6�u¢�m�,|��Y�$��)�>ꕜ�-\]���짡��\�y;�肺���m�s����4Wu;����**�cNp{�!vIK��:�m�v�x�q=��U����P#;�YQ�L�yK�*�h8�j���� j&�b �X�F�距.Q;��8f�6�VZ�S�O�Y|�]���Uj�͍�M���\p,>9}h�5�GV�}�vm={}h���i�֑m�B)V������9����H�Fv�6����oj��Z�����2�h� �l�i9|�k�G=g�a_(�ʗ��S~�6`ޢ+��5|s��uƺ�*�:2�m�Fh��wz�#޺@U��v^�4@zvK��ϋ�.����zk�EA���R�R��[�]���������c�0E���w�㮜�a�C��t"��"�D�ڃ�躷����3gS��UԺ(yw&� ��e��U]�L�T��z�[��EoR8dw����o:yu�d�m�zF����L��m%y�V������c���Q�S�VV�$E�S���oJr��:)��{uV͌Q��f�7,w6�ٷx��q�����2v��))xj������C_pB�S�.��8Ԣ�6�v�|2�s���Xm^��w��#I�
����G6�Օ�:�	�Uw��R��A<2}	ǳ�AO�d|	�w�J{ˮ�wƵ� n���Bʃ.���vby�lf.un�ӯ)�����H��Bfu���4�ul5�������C��ߊ�[�;<�ǒ�1�O��Z�}��KVn�6�

a�$}d�YR�y�Xĭ��N�NZw)���!ec-pu�u��.���c���yA��y�R�,;�v�Ã�Ic�(�Z�u����q���B�^�{�f�9;�(��D^G5�D�[��Nuuy@�膩��;�s,��.��k#䠓���v��Խ67+�w�.����#n&`rX��Ǎ2֓Y�mX\�j�y�'G=�V�`�B�]��D`"7ϴ���mR�v�A���3nj�����EPp坙�����-H� Ffݵ�I��j���a�Y���ns���\y���XФִ43���Ά*��[�Xk�9\D0��7�%�>%�Z�]�k��>�\���[���@d��z�5�Ǔ��r����mI(^�oH�'u/U�r�Q��Yߗ]H1mlژrsv�W3�8u6��M��B��-�Kx嫂S�jS#lp���"o���*�ηMX���X;|�
��[�Q��M�x,un��K/r'c�ˠVR�[yK.��k�����QY���8�gۮ�gJI;�a���#͜��s���[Prk���s~��"'���b�ǭJ��9��A��$qe�۴8�u&m�N���Z2�!�Ii���6y���7A��/)�� ��=���a��:��nL_l=�V�Z�pю�WjETy�y�@�����;*%P^�\�Es��
îD��ݣx`�K#�I�����_CA�iv���g�hQݩ��+���A�Ձ�jd��h�G����h����$����V�Jݪj�����P�sy�&<�g%��H#�k�,��[��&�b�I��9a��D�5
C&L]�7�Ćt����j�I|��W�V�2F�F]q����!�\�92�]Z�y�FP� 2�Vfd7E�#��:xwu:�Q�v#L1�۽�u�J�,�[O�c}yG8�v3mr�JMr��Ɔ�T1N���5[�������osHxIC��B@v����1���y��A�xP=�n��<�ɵ�#�'t��[1��LiR�gS�xX�.����ý܅<R�m��u�W	ŋ8�o� ���b+�f�f���������B��:]�q��}��wu�L�4��/[h�d�[��c��.Ƴah-������ N�)��k1�z�n��y\��{�j�S��C{5�Opu�ޝ�z�2�F�^կ��4�ɧ����@}�u�6�e��c�u�}�`'��q�bA�鱸3�'^U�X��aW ��Η#\%��u��s���Ze�8o�^��#���y�yr�Z�#��7�Dr}Z�A)�0ِt���CUٓ�Zr��J�`p/��|����*�W���5s%�dڤ�8���F������M�yк��+Ĩ�gFNC�]��,���}S3gEt�.;u���Z�Ć�����N��*f��o[��_Ka�z��#>G$^����;��
�s���ݞMp�}Sr�h�mq�H����7?���Pu��iC��+�!v���@c��n��5�]���}��l�rL��7��C�P���ݧt�*y�-�(���}o�Z��&E��[��q]J�tu��4��`�U�Nni�ֆ�\ē0���{D47�$?���]�(nܻ�
sca���3G@K��v^�J���(�-����{psܒs���ڬ�S樬�W+1M��:;��b���Tv�_9�Ɋ��|r�<����OvBv�w��εg�N�ƹJTs%��^VwV�)�	ܻ�h3�Zm�OohX8\��MV
��<y�g����,֠��C;�j���(ct�J �s���;�zh����}t�~J��׍�������>�`U���-�r��I�	�Յ��Ù1Ӡ��+�t}O�%h�Q8JK��+]�{���'WB
<Gfwgmg!)�I��%����WY����r+������v8�X��b�P�R��%wI�7M�"D��(ڵ���v������e�OT@��b��f�ΰ��j�����]�2f�G�����n۷�-����B�Q�[8k;WF��lب450��M��bv�k�������X�+>]�ޫk���YF��H5D����ek+u���H�փ�9�:rf��g|��D6��ʝĺv��x��Pp�|W9�Q	��*�Yu���o(�H@ʌ_��}�bzҿ1�Rr�=Kr�v�`ڎ�>)ua0*2�I�
js�YG���;C���0>ɇ�$�]�l�k����`|Ӽ�c���T�fe�{��[��4�܂�.%��WO� -��oWV�N�OX����w{�N��%͹}.�rZ��n	���Rܸ��яU7ʶg=�]��Xkn=���{~ڣ��%G9	��%��n �].g�xR��r눅4�\�nQ��LH��cZ�$֒DRqN�0��;t�5����*rA���.��`Ezh�/7{w����s �yb�N�f�k\�q�D��7hm-t1fi��m�Cv*_3���v�h_6�/���!"�p��o���R�����CMY��F.m�8�Ɋ���-K}�B͑�<�f���-��i�)fWaw�ŷ�pX��w%f���[(�����6c��Z����@��̠,4�v��Ƒ�EMKl�*W֎m�k���������U���"���i9J>�9������MŬJtղ͚ή�u�	ղ�]��6�n���ڰ�tv����v'����j�6�r��Y��"B����(�5r�v��-��LL��4(�~)j�� ֍�]h�GW��V�΃��{X�+��'�=e>��I�'�i�ŷ�������'<ǿb"b�xHIi�8.ٕ2l�In޻�wpe��ǝZ7����YǑÙ���R#���������7�D�2	�b}��W<zG[�A�Cj�2j������*[�tޘ3bԩ�2�y���,6���qo�V��6�D��y9@A4ޅuʻ"�1�\�9���3`���t³E@�w�>�Z:�U�{�yYS$W7�+��,�-jU���pt�fI�7}p��s�K��
�h��Kze�D!����\���yt&?�g5p���[ռ�ܖ�x�f�}�1.����B�ky��ژ+{	&�z^�׼�%j��'b��6��U������h3VHj�qNun�6�n��5�IN!�j���S�l_�=F�Uޓc<N���(KQn�dӟ�7X��x�F'm��Ք�ږ�̡�3wrEu[cq,w;1RX\�hS��)w�.�v-O6�a=&�����=�Y�+���4:k�OtF_v�����FV/n��c�݊���BH�о��.�WY�쵣Q|�W;�q�sTH���Uv]��ogY�6�L�����duojI\F���",ם�@Ht��0�7�(.��FC��v��vx
�S�-��}|��;@;���D��&�vޡ9�ml���__��4�mLE�p"�@�<Z]�x������f�un�5w����&ݕ {�eWs�4�]eÐ���
.����YW3fO���Uv�[݉rC'��!l���Ί���� s��ҝJE���^����	���L�ma�V�eɝ���7BEǙ��f˃�w��m�00���/'%�(��NR������bC �n,yXU���W0�u��2T��9}���N$l�B�Bǈ�=�j��x�X�]U�a���O5mo[���VW
���T�ΘP��<{�Q��0[D���Gў��6��u�2��P��[�:�L[�F���kh�9�U�2�u��,�%W<���u���Yd��TN� ��*�|] e�'}� ��oM�K���]��\��a�9��4���Dp�E�h��k|9��
�S���gc}+��Ӗ���W!
 �
tB��|�.
m�sti
�u3ϳ�P)��w�|*���@߽f��Z����u�5��D`�2�vd�vn��C��|�#bR:�n�7E��sWS�6��l�� �\�iuuP��� ��I���op�
�[8W[��ҹ�{t�1�*ud"V�������[��ѡ���O�p�X�[�,e
 ]�ӛ�Xg�:�ڏ������W>��b���:�Y����S`�d"�f����G�=�y���ܥP-�����O��	��ZU�*���!��jo�б��tC*�85=�0��v:ոwQ�:�.�ǋ�-�-����@��Sř�9.\���fz�Rb���P��*V����g��7���3a}�2
��Fҽ�
�>9S3sqSК��1�Wi.=�pR
�߰gi�z��׏X�G{�\�:un��W�,iO���(,sp�(u �R��v�̥���x��׈٦/*nop��+�ք'�I����Β��P5 �S/�Oz���[P���S�2�x&���-]fa:Ѱ���;F���3��$����j�w[�V�2���Ԯԧr�Oe��Q���3�t&UL���!2�)��L�������/UbQ��I@���⻨�\ĭ: w
4��Zq(_��5�>�o<���Xsht�K��m�S'4Z�Jܔ�'���u,*��0�}�<���cnE�˜��������<guv�WH�i��N_q�M�6�$�cl�ƚ�"��`��L�շS&�uIQڦ�r�h�N���&/��&����Y\��	%,i��6�/�ku�W�oc�}F61�fT�\�a����M�kg,Ցj!y��kg5;L9Φ�θ��B�(t�vk-�޼�f���W6�_vw�jQ^����6FޥP����]%���/&�L��@
:��s��v�ԬpB��1#�7��c%b� (�n%���bm�d�Va��v��(��V����y)@��I�5N�f���nku�n�eh���ٛnI,���_�T��ur�%C�13�l�f���#�v���Xb��]}��u��.ዩ�o~}���bq��q��^�Zt�<j��7nڔ~��)�Hu��wAQ(��Æ�@��y�qq�P���EB�J�:R�Oi-���]��,�-�Q��V�}�Y��и�x#�ϸ,��f=Y��0(�u9��P�l�o#�m���unC��Z�x&��!;��%t�|%WZ�Kq�]83w����]���V`�t#b�+{AV���ӻ�8��skP0WK��vjv$tEӒEm�љ(ajD����j�-U��ID��Q��w�w������vݾ�,nv�΁7�R��7�Q��m}� �:��L�a4���܅�Z���C&��e�sumd��f�t��s$���7��؅�H�����F��lm'.����>�P�?)����(��ty�EwXh�Of�� ,�{f�����U����Mb��L�p�e޷�c���w3��v)!-3�Lv����ʯ9h|�$h�v��W:��|�����%E`��|�`���U�Uf�*j5}�$�{�Ge�ܮ�am1��z��Ti�\�	hL�m�B�J`�C��Wn���ʸs5VZ������J�uo^�����t\�]�f�\�nA�[�9��fA�A�M��oX��8Xo�GvZ��5D�i3&��t�^n.ҫ�h>�q�M����o�f�W�:��]'�Ӛhg&vV��+R���~B}g���R
�T�|�MP�Zڭϭ��2�p�/���С��)٧�YYwY���-@xA�!"i�.볱�Tĕ���o��.��6��ǐ�A�+�6:�j{YEj*�<��%`d��*��n���jS���i�A��[R���p��g��)nNc���s�h�ͧ�)Z�N��#��*r�g��%��Qg�t�����g%��VV�+�.��x�8�
��BvL�l���ۚ��\�(�B�8]r���qj��j���W�Y��6����%k���E����3���:�1׸J�V՞�͌E���ƍ�.n��Ӡ��	��)q�xT�-�1[��ᴹ����kx]�2�}a�;u��C��-�d�&V:���U�	�rn��q|�q�jB�� �6ʙQի!�.�rS��.����b����ϥ-y�;L�vڼ4�'�(������L�]2_^^�.f�S\��-,�r��i5lVO����s dN��{3ԻMI�ֱ[t��6:�U�ث�Vmg(�k n��m\˦������� �&�YWH����*�WX/9M� ����S5M�fY>U���! ��,U4E�{7�3LZ;�>��*��َ�rHm:��GB/q�� z��W0WJ��R��av:�`��X��q�
@��6H]��h��YD/��nd�W׍�徼Ŗ!��)%��1�˻������!�r����U�T�Kew=�׬3���G�f��r�;I�ɭ�xL��-�7эE���x��[�j�ò��):]�a}�Yٕy�3>s{i�(!D����à�j��n�pVv;��1t���֪bWdc��W}N㠀Tݽ�f���ځ�Kh��e���#4�Q�KE�����e��3Ț��j��.����S��fȏ_&;V[��*e�e⮇m���j>k�y֎9�kr�h�5`'�X��;���M+���=�k|B�0P�����*��]uK���t4jr�\t_S�#fв��]E��e�`篩q�z/X�g��e�P�?�=���xfh�E���'g����{{�5�b���	�ܩ
��/~؈Ui��0�2��Z
|܀7.��9�)�;�4bZ<�qU�o��2�̺�wݫ�u�=��/v��KZ��Y���7��۫��G�M=A>�6��8E�m�Ū�R[������y�83��VSY�`j��@��T"��ۛCeޕ����> U�9�uԝM(���A�ӵ�����A�辻�a�W�b�1��s�$�8�!z�L�+IDn���o��tI��[w{y$�ꆰ:����)J��^�#G�}�4o�Qg�i�����u����ι�a�h�� ʏe%�)�an=ٔ�[�`uë��\<����l��vѣw��4�Ңl2�V��&��n*ur"%;#6��i�e�V{��ѮV㈧��N;7�fs�Q�P���d=��dc�#��� m�eo
r^8A��aZ�����郑�h�>�c<��'��Mù�/f�n�5�Vw#��t���][�zd|��Q��Q���Dq�cj[�ƅ�
gh�1L�ע�L����څ��V���AS�iv�|-��hc��*fƍ�oN�h�Q�������K��أ|o�n����}�Jź4�6�M�m�-��V�t�!](��.g,�e��}G�L�T�⹽b�g�(�z,M��+k[-�����#��xWS��'���N�e��(�gL7y)�
NWX�tm�/���]:.��`��xcN�m��x�ܺe��"N�5��|�XPf�.ĢEʴ�ʗG%������}vz��ߜi�Δw[�-��.������|~��<���-}�Ma$W0"6UœRy-k�[gm�ݛj��f�Q��Sh��8y�WM_ک�ˤ#3��iiY�n�1��/soip	�������f�b��Nθy��;s6�c�x�>Ɂ����C��˾�3b���<��uihYv��p�7�*�gP(ᒮ8 ���Y��:��-u�w���Qj��#��� :>Tf�7u��f5:	��e��9/ 9�`W*Tx����,�ql֖#�nP�}���v��{�@V�\�]؂�d�H9�x&�"W���;�Ċ�t�1js��f.oCʽ�ݫ�l�U���X�֜sr��l��,��I�\�;��͌G�V*}B������2F����<t`|,�t�;	Wb�X最�ٰup��.�J��W9�� �°,�"<�ʆb�1��~�IV�t�`�T�|�&�>��.�EԭT�L��:�p�iA��b@��ǲn:mnfLś���[}X�u������Ӻ�hEo5 (,�T�p0���@��y��4�P��he�i���zU}9fs����Qp@4q�fL7��.�OF��t�0�a	��Re�kLY�es6n$�o��]3�*�N��/�m�>�y
��u��2ۙ��t91W8��_+��&ܓz�l�f��(-����L<��<�x�.ȍEu�%����oCboT �:��n�SU^��O�ݠnm�q�s�][�GlJ���⯖�޸*v�Ka�3UBi9��}�
f7��N��(��^��-�tczd�W(�I���D�΢��I���	�����
ëHų+���nX@`J���pQ�i���E���m@�Ü�A� g`�5��ܲ�
��E����M���R91^�r�p���j�/r���$(��u�뺦_m�f��HpՖ�@�1N�FU�m��t.�r�r��s14�Qޭ]�+]�]�Po��춞l��6�V
euӱ5�YW�Vb��	E��V̣B����{pj̏,9���bM�;N�1"/x�R���n()*E�l�" ��9;V��eݠn�%�˙.��!Kk�%����bHY����@Օ| �۷�I仼���W�9��}/�,_(Ҡ �9��lV��Y�n5�Wa'wZ3X��Z�(��5�̮J��P�yB^����纂Q(FT��ݧ	C�9����K�h�r�-6R��[m�/q܄qn��MQ,V���y��ό��A��)]n#�E1Ԇ:��luE�$��Z��ɏ��������5���kEQϳ{8`r /H��H�VK�H�E>ڭ��8� ʔ��-�oF���d�����jm����11���뛲�I+.�������1B�Oh�8�v�R�Ɛ���Q�*X6`���Ê���[ ٕ���o���K/#�)22���t)�N�� 2��¬a�Q`m�����a���y�z�h��V�*r7&�\����ن��d�Ggi<�}�]�S.,#�c��s#�=�@|��[L���n��)�W�ᢩ��R�Bg�m�q3��t]�5�7�.Y'�ZL�Mq+���爛�.ܽ&��໣}R�k��r|6͍k��.k�z��.]��!N������c���ތ���g�=>�
���D-v���4j�Em�r���ĥ��fJGu��O��n�@�n'h�9#�������u��5�vsν����d�w9� Q��اӖ5mvw+�i��)��@�Y�U��Nr�3 sO,�3!��R���g�:���e�7ov;8���8�G�t��F��{9b0�^��Dʰ��Cijo'V5J�D�b��؇��|r�)��h�K��n�ӭ+�4�Pz\��Nd�{}6F�%k䨥[�m��t�*�Q4/���yO�$�`�B��P'(��(�T�0q�Qe`� <��s��Fuj]m��
BF��{C#���Qٴ}��i�ʖ��ى.͉q�ӟi�6��xs]J�R-�N��Iη�%��>%�ف��殶�a� ����7.���-�6V-(ut�
��G�����a�a�9���V�7h:"Uޭ�����1��Q���ֲ��(5���X�j����'w�1���*oJ�����q�C����ˣ��m������,&�>c�Dc]-F��A�V�	B��S��D��WϚuyl>��(�fv�v�K�, ��=X�hLc����4)IU�4���M%�t�+��q�D���*M�|��ռ�����C3>%�d�W>]����|�,�ە�׍D1N1s�t�.'yPlݕ�����J+yMN��tu*e����޼�4��bj}ƺrŤ���{K�m)��	���
���&��bvQ���L �],Z⹌���io�W%��kƂ�}�=z��S�Tw�!�M�f��4�!]��p�g�-!���"�]����)���0zr���]�4ΔH�]�&���.�-�]�z3)�2V�ӛ����WYh4�f����Mj4�9�i�l��w0:�;���p��or�W;/����R���`i]�L���6�P����%r�۷�J��W(��t���<�;��2N�.���`�3-.4�`�F�r��l��9���R�Y�Fݎh���Y��[VWv��و���kr9����ҙ���&��蜾���]�GMX�B�4~���ۄ9��w�G������g �8V)8҉�����j���N^SU���BGVp�õ�Wj�M�N3��ivt�d��3>�j:�V_&鸲� � b�]�v+J:s�S����s�\�q���z��O���P359t�E�N�/m����8& �N�˩�2���J�:�G�#�Z��|�R֭�7W3������*,s��;�#M?��b��)ie�%����Z��k�:W4B3��I�w�
�G� ����+���+��1$~:�t�	�ʘ�WS�A�jY�&`إ��i�y���	��=���o;W\1R����3��&`G�`���ϊ�79v�\7E�G-1��-�6&3����wgw6l4�PW�U�K�ou��Y-A���d�fw_'M��Hs�1�9˥�S��'5Ia�6�ur����kR Vv#�B�M��ي�@�w��֞�].���¯y�OE
�%�2�[WWՔt��x%��lw'Z9�v�T�:��Z!B���H��IC����.���.�~0����%�E�.����`�D�ZƘ���n��̍�(���z�.�;�o�h�n��V	�wzuki���n,���">��������ۗ��Tm?nN�Qۤ�&�t[P}8�R��S����ɥe��N>pv}��<�V����I�|-D��^V�|3r>�xF7���v#ޛ� 9Մ��9֬������BѭH�m*�t���~̴\�wc���r��v�X�/eJ�}R�tmQM^�*drh˕/J��3��v"��������sLT\ I���:��4+�aX��WT6q]�bl���֡)��g����鴹�T�������$<�`B�e+N�ga错��)z'<w�B�R�\x*���X�l���ʼW{���J�҈�71}�Zd$!]����U�d]�R��:��T{[(R��_r�/�;�
`�'�V�6N���]�=�V;]VC�gh����Hd�w&���	�}of.�>}��l�!�Z�������}4(,���j�����u�.�	t]�|��Ӎ��F4���	�n%fp��0>�~�-�C^��xۣf	TFb�0�B5�fJؐ��9c�I�|�K�hV�՝�ʾ!�P�6��L[3K��v4�0.��=�L}�D�#�(���YU�s��զ
ִ����є�&2�gN�����Wq�;+2�^��}�M�c6��]w���|�uHU�Uͨ�
\��
��˚�Ǵ��tCc�b���N>G���T��F��.n�܅h�X��C4;Y։�J��� �o-o�m���VMRDf`��5UUURRDSUK�UT��T�fUDR�U3!DCPUBSEUY4��MU,�PQDDf`LLTQIS��U0U1fbSHPd`T�BSDE%PQR�S@D����4��#IETTRP�L�#BSH�E$TQIAQRQI@Q4�CA��14�%�1
QE41L�L���KIT4�D�14T�L�RA�R�JP��еM%,I��4�0QBSMT�P�#IEUU�THR��AM%4PPЕ@QLMQU-�UDACDH�ITT�P�%-RS15PQE14PQE145M%4%-S��TEQAUC~_ñ��R;��so�.��+Mb�ؕ ^�*X�c�4nd��m۳����q�7�ԉ���)�ϥ�R��e�z%|o^y��꿕C	@�f�*UG��2����Z*�w��ݶ��� 8{�T��p�a��*��<o��v��W�F��વx��~�6bc��B��>��ƠU�Ӛn���/=BV+���r�ԇ�� ��Ib3~on���9pa��1厌?vҷ�-�&��<�Ţ�u������-�;z�*����pL����yu0�`�a�j_�k����2����<a�:J�����<�{�e��0��+����#�MގW����T�B $˘��?!P��ᬹn�R�W]�׵sXlҠ��1|��<�φ:��Ȋu��o'��w�a��*4B��k�'��p�,�`�B�'D:���TY��c�*�7=���bn� =;[S�����_sق��_ν1���'N�8����kк�]@�S']v	��=����)<��q�'&ަ+Dp�ڸ�aʟ�����&�q�I��\�z:믚\~u�Q��5��������^�7{9J��B_s��"Yz_�D!���.s��� hD��A{��ߟ��|��Z��|گb4�v�L�ͩb�bݠ)J���)��� ���vJq�ծ􎟑���)c��6��)� �=>4�����%���ф��1BDv_+��+��p�"!\Y��w�N�.Wm�(�扴�b�V�������7:$=��ϽP�U���m{=p`�K]�w��*�%���uP�+%�� o[�CM��P�/r걼��	�����Gb)k�1�W��y�����'��c�w��Q��=�o<߫<�}�"��&�˼�6�h�@����rj��.�1p��\ێ�����Zk�^#��kҧ0�q"1|~�4vH��mz���j���!1��*�K.����D˺}�9Q������ ��,U��.+䪀��ʨ���S;F�Wڕ3�_>De8��"��׿8�U-ɓЛ�9�����$�1<>�c�����b	=�2N�m��6nŷ0��F�˅�;�c5�̚y*�y�;P�J�4Z��-H��K=�!5ݭ)������Uδ���a��_���Fjt��������}yS�W.;�G�bD:���o"q���P9���M:J_m�^��/�e�ҧ�a�!0����Gb���W�����M;�|x�2��C���5PZK�Nς� -�Y��dƛ�vr;�Ԣp�wa4�-���Ω�#�ق��b�w5]@$�Lj�]û�)�����n�u=9��ƞ����V՛�����_Y�Е�!Lt�b,�s����1'B-��*І�Tb'8�[A|�5�m�3Ӂ`L����[Oe�ޟ<\��i�H.�?	0��u��e��1��G��2��ڎ�2�Q�|Q�p�7c^�R�֏{����pAA����_�jc��θ\����$�<�%��U��z�n�a;
ǯ�W�SJKyD�Q�&c������S�Ӕ��n���!q��OQ_�p	G��n��f7��|"È��B���r�LP���c�|!����К�|�?t���)^����g�wV�I�* �a"��|o��.���B�T����h�}�u�P;ʧԽ�����米=���NFœ���5I�p'�i7�+1��B��p��p�9O��R��	������i�[Z-��1J$��� F&@iV����"���z�~�}��l�b��7�����i�q�:!���`7۽��`��S$�Q���&�?�ԏi��xܾ]r��i��6��	P�[�َ�/ *��H�W0t�c�|:��zO�g�
�v����L!�nuSTӳ�!���1I'fKf#B5���58	|��ׂ���vO^�6��C,�����J���ȼ��}yx����
�<�4MˬF�w;g5P��yS�#D���/x_�b^�8��,�}���u)��\�!�GRiVw&��]����n���<�՝|�L;�ӣ6�u����t�k��[�g1m�
L�^���s�~������mу�^�pu���8��f�9`I����er��v.K�)·�[@��^&1��,-���s�
���4`�,o:�"��̎������+�<�r�����V/�nШ<K���#1W&���6�
��.�u���c�tf��ŕA����\��%�m!��n��]H������a��T���X��e����OB�o�rJ�}K��,�5̲v�c=&���7��;��9q2�T	���Q��V�7 !���۪�Ώ|^1�YTux����U"�<W]r*O���Q���w
����F�ƴ9���\<P�X�����!�5��R�鈴�3���b��7�_.ח��!~�=$�����x���ng��Q��+V��,�kw�!�c.�b�մ3jkK�g���N/>p{8�IF��J���|�R=[U�)l�P�Sú�4���NM
yb�N��l����QM�ީ'w��H�7�Q�UJ�Hu���}�A����޾n��3�ZEr�%=W��D��-�ʏ�:+P/�wȚi��x�2$h{����SN՚�g��p���Ӗ��@��)�֮Z/�P��y�1�hksa��9�=\�Q\�ر˵r���U��־����@�+��ɝ���(]�̲�ڙ�;Kd�އ��e��F��"'��<H��Z��H^�;{�ism9�hW^b������]6~����0E|ۨ��wv���F�U$G@}]ˢ�<���C:�[��8���BY�/x�
�S�����	�VYω�D�f���*���U�X��3�w���sx7���Uҏ��U#��t�CSQ�H;���b�g��I*d�X�����NV�ߓ��z+ ��]R�<N�#�!�htƃ�^��mu��O#�U�v�FآZQ`]L͙��|����,3>�ˣ�?Qx���H��c��7���=��we;*O{y�j0���t>�¼�9�@R_�(�p�݋��ٜ�0�hE��~�N�#�r��|��=�˳j����)�εZ���.98�el=�(��;`ɡgI�����@T2%=�;z����z�S�����J(��E�Yd:�q�qϒ������Z�c{vc�ܥ0/�E��t���fa���_U�a��"����E�4�Ꭹ���}�y��wEu��7G�: �hK|��1]+Ŗ6�J��q[�|�O���{ݬ�Yz�WXf��弩Ҽ٭mbz����{��}�֯{���+ j�θ�7yڌ��a���|WEpT�nRj�n�p��w�J����-���X��e^�',�v����b~'D �㕪�K uPb,crEC����rx�o���í�w�G>oD����cCn֒t�Fx�������uj����xdG��d��[��ҕ���ˇ�	�r���e�Y �5�A'I�7��뮚\~f*1�3�^%\bn)�]�^�k�}�v@�!���p�f�p,R�	%r�29�9T.��В\�g����������8`�K]�v9�Ү2X��!
(�t��p��K[u!V�R�Q� �f@ـcx�PK}9��P��k�1�W��'����� |�k��w~*Ƈfh�=�_z��⫈�#�-&��ʣp�K�\��T�*x����0�F�Z�CWOwN �X�&�0Y����GQ	v�3l�:��/�Ӄ�2TK~"�cgsatQ��!�K�邲� ��s|���*�;�(����7����5�گ���S����)[���K�Oo�MTH�R�2nt<�ű�Ւr��13���y^����^����y�r�|T�guQ����N�i2gT��lu`�V6�dX7fP�9�fw�W���5��Kv��։��,M5��h).a���ժ�{ŭo\ܱ��;��d���b0YvBqD{9�����O-�橗����ɷ�6����.���F�� g�\���wu�y�N������F3\�ɨy*�{V�~C�*��Ә�������S����lѯ�
��ZL_ٲ��١a��O�25:Ž��ի�c#K�ڽ�sde=LKۙ�/�'v�3�adEL= !��v� U�bіp������ׂ{��p��;��wբ�p���N�o�\Nc���n����MT���*��gu���vեQ���43;�ᛕ4�}���W]�pU�c��-F�3�`ˤ����}��Õ^�Oj�q���������l`���S̾߭��+/�f�U�~��8<D�D����r�S�3�~�U���l����mW��z�4毣���(�EY�NS+"���!|P�[$tyo��庼�'-�<�O ��L�B��J�Y1Bj!k�>�|!��`3���|�?'ڮ�}���r��/�<Iڈ2��_* �����T��U,`���1����s�ĉ0�RrOq������"���[�X2K4>��3
 Jt��y���}¡k늸t�8d��T�^u�"L�w�V�]��T�����l�JE�5rw{�˛n����^���X���K�B9rYӤ��Q�٢+���{�!Qr}��1���f�x�]�U�;�
�2��N�xc��u�<���rew>T���8��sL�N�;���M�U��4�S%MG1" 4�A��� B�]�m��jV��r��4q���|^����U���S$��J� Й�V��ޑ���=�����ڥ'��N4�3cxԺ��nc�18�x@8�$u�0��*�(��+��6�
]܉�Y��zc���핦��u!�,�DH��Q�܀���ȡg��`�GC�f�T�oi��Lt�����T`��/Y���u��ZN�&C���%Wo
739�;S����M�S�]H5����U���?]/)��½�u�`Cp�:�]�Q�Fk��n"�]���rX)����n+�SZ�Ce�B�q7B�g��B�����/�S �:u:�V�Z����������12^�iS�ƮB�߲+�#���I�Z�j�VP����<�Xy��c��� �|=�YQzy���L��w�5u�:�6"��
�x@u�Ņs8��O�'��!�\��f[8.��1���:ꆺ�R-���S��Sf��0�1Vz"���M[&�Ray �("�`����K����¦�̻i�y�>+��D�lq	����JY�1������Z��3���q��b1*n��v��97�F�]��a���h�8����L�D:_T�3s����H�����Y�����X���$�ͦ����ٵ����+����Em:��!�]�|�:b.!9L�}Oe�[����mL��>=Ӥ�b��,P�����uM)�,xWs��t�kw�>��a��z��اx�[x��q��Zn]��2J5�%Q���Q���t|_���<�')�c���%�T�_1K{K�RY��{D=/zdbu_' �<� 6"8�r�T*C�5y��[y75��X�����V��_�Y�7
f�8ܑO��SH�$�Az�d�o,8.%�W
�WwIb���{��>=���d*vٌ��h�b�l6�1�'�l�ك�u��^x��^x��ħ���"��9�hJ0��Ga#������Z��|Lb%\3_FG�����s�9�Kեj2�U=t�ML��'#��w��ų�~IK%�p�ɼ�V4���_oU�ɠH���U�x�t
�ϱ���^�^]p�R{-������|�z��P�q��/
 1Q	�K@Ȱ��4�u��0�R�0�Ǡs=����	����y���T����'�w�O�>����#� �P�4ݚ��ȧZv1�E��\�[��Ռ��R����df��[,͇Y重j��+Z8u���-��u-��r�2���U(���<`;�YGz'��ĕˉ�G�v�^]��-��������K���'	��9� ����m��ƏD��
���P���~�������u5l��O�|Oޖ��Z��0��'X�OW���i�&7�;�(��$]��I�#/s�k:8k
x;����	������z�C��"mJhn�V�*I�������\w��+�p����V����j�v���t �=���K}�>e��"_W����@@�@ͧ�=w���oi�{jx��Q)_�~�?�A�5m�,T�ܑ%|���2C��5"]�������LB�U���Y.���$�h�W?��סi��x�C���_+�%K�݅騶���a��ۄ�_Ε1�]pJ &�Iܙ@L�
r
+ltq�8��ݖ��=���T�f��Bj!�o�|Ԗ_��_<�,��^��J�[�4�Ŋ�Ʊ�z��6D۟��[<���QX��K]�w��+^��BfOA5�E�`)����vQ� fx�"���D�Ȉ��K]p����͖7!:�$}�}��SE�����	<-^�j`��2���,�TR���o�8�]I�ۂ>�"��;V��v��.��uF>u}(�m[����v�k�о�k4���*ޗ��K��+[��jZ�"���"����(�q
���,1�"Y�'r����\(�GW�����jSv�"��,��
X�<W��Y�6w@�޳��<J���&��	5���J�B�:�B�:��,��6�Vb����*c3t!�^5��I����#6��p��#M���ѕ�E;�"Է�c�b_����z�tB�Hlj���]H�� �c�����3X��ո�gQ�U�/ �}t��Q���Lu�Y�N�qR��RQ�l�;C�*�-=��=�;��a��t��L�#S[GD�W<Ҳ_j�.v�{ӪXD]�Z�M�G�ˠ�ӬE��5�,�}�%�� XA�����\5\:���$#5�42)��H^��,��V���=V�j�u@�:��IZh��f.�˾2���>�F��s9��$��}�(N��rԨ��Y+9��m6^p�p ս񝜣�+���U��
�;J)ӝ+5�E��RC*�}�_:��o���3���#�����;y_0I���`}D�xna81�������%����{ �y�@�-F�*��IX��jDnE�T�3�%@�#�O{_$]qY��.��Z�ᕉ���q\���N�u0o00��1�;�.���R��[I>G�{W0��mj�b^���Ί���cW})H�V���v�
B`�e�{�Z(sO+�{�3�؄]2Eҽ�t���%��j�=vͰpC6:�����oT���}�~���0٫���H��,��V�<|��ƹ@۠�oR���d·;�~�Fg����X�|_���X��s�W��o�\��xµG6��[�U�mt�wHb��vo�%X���>�bEH����6�;6�-�|��r���ٹw�8S˙ �!OI�%X\�+^C��0�vo:����z�c�i6�۽����AM��K�{`�_(l'$W���#;I[u���2ƙ�6]*|�8(�Yr�p��h\������&X��r���(G�g;*qۀ`v��dr�:4��9�[�h�,�ʡ�y��jm�F<޹�O����Y��g_Vv5�D�Z訅JגҼ������iV��� d�KZ/_H����T��m�89)c�fn�0j�WN]�N��]4���c�o��r�;�e��J���*����� xdB���:���챸�Ry?�v5@��dm�⭺3���y�[O5P���E*O=s7v��g<yYJ�Z+9BYh(Ҿ9�L���'���)��G7+��-�u�m���mN����li�WJؚ�z�n�\dy��^�[��O��6偕�s&�V����iF#���V�+�X�R����W:�ѺwV�u �V2����AX�g.h��f�8`C�:����P| �4DD��U54%��D�%4QQ#MQLE�%	IIT$EQTL5A4T1BP14��T�IERQMP�ERRP�R�Ҕ��ą*P�-DKBPD QT�HRҔ44P��E(P�0�	E%UQCMR�-1SCI@Ĵ��4�PP��RR�KT�@PPR�4	MK0�)���S@DД%%T%D!IL�R4��)AJSBQC4U5EUQCHQAAU$TRR�%IB4�IT�--11D���4��BST� R�QERP%HPuw�5���{ߙ�e2��{Ge���v�ja;"kk���9R]Ha��2;��]�B��/��O��JW��指�����H�u�����S�<������<�"�#�5���Zr~����w��5	[7�����������%�`����u	}����� <���~�}�>c���U��2�0��Z��7��=�A�亍T<s�9�2亍}�6&�������r;��qӬKX<�4��U!C����K�`�;w��$�9Q�{z���ɨ�"�ؔ��� >���և��V�����pf�}���~�d�_`q�ζ5�Ժ��s\���sX���u ��s�˳>�pdd����d�gQ�?[�%%厥�~�F��a웩
�J= Tp>4@��t���^�y4�f�Z�Z��� ��@ T��	��gS������U'g9�èwHu����<�Q�r���iyI�d{r�`���w>{���.�P�v{����K�n2�.�>�$�{9����W�s���]��=�ӓ��:�~b��T���l}�.����oKO!�ԝy�{Gp��'�ﹳ�;��P��5�����5??iw�-9;���sA���ހ��<4�����$}p�USk���>�3z��^k޾�FK��8fA�K�>��0�O�r��ч%�jK��p>�w��5Px��n�˒��:ٮ�L�K��{^^Gp��y�6�f֦����>XD��+�|��o=��O��x&\>ø�'Q�F��:�cRj<�����%S����?A�K�?u��G���kA�d��5��;��=��9.uߜ�
A����'L}}"1I��]�1�r�^�%�߼O��=^ے��ѹ�\���5���uR��Ǩ�:�p�x=��ny�Py��ѸJ~����5�'�:��z���A����7� ���ԁAAAk2x=�v��T����f{|W�G�T� `�H����j\�4%�r_#~�ͿK���w�4����\���{������C�ը}�?gf�����9�#p�p�)��)���
�>��f��^��䵰���N5�j">� D0= (k��O�r}�s_lr亍K���w>�\��|���*�K�a���B]��|9������^ƣ�wj|�<;���K��FK��\�vts�y�wk�n��
��A �a
�l:�G^���-��وP4��*����!G�V8/x'c�u��ւ����p��ewK{�ĉٔd�9��\x�g$l�/B�)���y2����{�90L�����{�v)�}r�ix�'()lcۨb�1�I/gwa�}§�&O�8������7	]������;�4�}�p�>���n~�5�x}�S���������Cs�rMG���h��P{=��9~��5!��k����������E�#���v�ұ{q,;�%��|k�Zf=�A���y#ۿ�m���=���7#�߿��� u��L���翰J�����}� �#���fV��]�{�^S���(��pd>�ט:�Q��:u��9&I�֏oe�:�#�Xr�K�jN��]��%�佟w�����gg�kk���.O>�������ݻ&��3[�u3�
��mC�q>ދ�&N��j��h;�Gp���5&�A�|3�����w��%�-95�_C�亍A����]}������%>˝}�:`��ACH���z���Ȉ�c�|���T}/-O�xs�:��2�]F��p��GI��:�����}�����7����3�S[3�(9}���\�f`j~�$�r���������N.)�q��gj��;�����l|��2�(:~�����K��������_�́�u?��a���%� ���i:��wa�ܺ��	�^�Ի�C����)�r���>��޽�d���V�űڼ�@Q���$�c�������ZCs�N���=�dj� �����w�;�5�}�!���y�W"�p�I����:��P���A�;�/���w��:V{w�S�8;E�u������9 3����� 5�%���\�f'�g���S׾iw��{<����d��o��N�P����>��ܚ����4;������c�K�Z<�������n�n��F���{dz�&>�@P����u�%~�P����\��B];��e���=���r_֧��ؙ�e�_�{��%�e�������d�sK����6}{�~�޾p��_������p=���`��q��n���b{�S�sX�w<�I��N��ѸJ}�d���y�(�r]���ׯt��!�G�~}��#'���J����� 1����ܒ�	�T�X���Y��r�r�h�+�)�4{�v��������#��O��2�/��}Ͻ�#}�}�^���gb�v�km^�(ᆆ��n���������U\���q;�U�a���t��Sj�=|sx3O���w;s��nۨ���'�߳$({���%���sz)�\���廿��ܔ�.A׸w�RnL�:���~�F��%gx&O�ru��<��)��:���<��Խ�;��4Dh�=�k{����:g{�����;�:����5�����}'�����^K�u����9W1~�~y�Ǹ:���Gg1?Gs�_a�l�S�ܝy����_Ӫ�֐�?Ov���	�>>���z#ѧvg�W�=�oגw>F�8��[���5&���~ךu-��6{p�1��ާې�亍n�)�S�h>��J���=擯�>�������O���ڀ�Q��
>������W�xk+����}q{��y%�T�����K�k�	�z�G��������^hw?K���۞u���g��p����sX~����I��k�>ơ)�<���P. �@�A�g%'MK$��Ȯه��}�-I��[���G��bn��ܝf�>K�~�.Ӭ7.��!O^u��:���_`��4����?W��RRS����i29I�2�����t@\	�Ȗ��)zv�n{u���'�>�kz��#P�u�����y���U&A��l�4%� ��h��@}=�a�7�˩-����+�_��GP�B^���_���.M���v����yu���>7�#�/s���9���us���u!C��կ�:�~��?^���ܚ��R�����5�W��k7	T�Q��9��K�N����~��W����{=�����t<�4A^:���gFcy�*���ׯ�A��h7�r]T�'g<���#��j�{.��~�O���;�
vX��Q���NK����n<������a������I�}���4��*���+S� }z�����{�}	��rMG��������o�MG�{�>���9{'�5�hMk!�#�?sk��'��s�]������5:�5�!_�Ġ�d��Q�Pk��R�e��}^^�����"f��IINC�f��=�I��W��P�=�A��4;�����9#P��ZA��y?A���u'�2N��� ����Xu\�P@ �V8%GF;�OH#<���uoK���*<�c�W[�x�J���ـ�p-���},m8�H�׼��V�V̧|U�x�Xmԭ�7�6�L��o>����؏z��ݼ_���a��z�^�uԖt��GXe�ݻ"�=�lT�G.��{7^��~�����.���=A�5W�����u@oxk����r����/''��`�A�b�}�v�HP�>��g�&G����w&���?kZJGà(�(詿+z��TE\4]E���u��*����:� ��>�����:����q�J}��0߸?��%t�Z<�9��5=u����]T�z=�A�ё�{~���:�!�v�^�z������vT�2Y�8�9�= Tt.�_�y�ӹ�\�_o��kY	Or�a��9u4%Pl�P��O�tf:�	��~�]�G!�BS����G�y��u���C��7=���%�@�"k��!�X�궻f1���@ y�mz���=��͆NK�̀����<�#%��3��5;�#���/֤�� ߸�F�R{A�����@������a3ȧr�]�d���R��}�����Ɗ�̨�K�|s�N�rle#m��^���a��&厊Gl���i�ךɭI$n��;X2�����ߠ�S�X�N����i3,��u3��G���l��}�q��pvENQ�<Y7����ֲs*�9L�;�U���o������5�ʹ�q�Kơ��3�W��x?���������"�y�A[���ꘕ�I;פ��;�`���8� ?�H�_�f'�m�,�T�K��F/"�k��9�I����s�����U�ڻ*F�Βt�������{Hʕ���+�)cyv!�Φ*�r��y�7N�򔤭��+^��j5l��C���Y�l5���է;ȍ�n������@�k�k4#{���}jd�Hf�u��}��}8�k}�>k=kq�k7�wGx<�L�={
8_oP�v�7�=1�v���f-Ҧ;>���g����`]�ڛ�J��.��;�9Ng�U_��Z~kTap��u���9��_��O:�.q���(�L�;�F�:W����dީZ& �X�@����2��n��r���H�9U�K$%Y�.���]j��dyt�Vpp� j�2��ai"��}9�������6X�����N�L\�*�f��[����|hq_B(tt�K�<�7�5��p���t�a�mou�M>T!nu���A�˦LXc&��Z�wP`�>H��
�td.9DH@��o�	�E9v����4*���M6�y� p�(�UH�3�;�CT&�t�;��k/��]qΘ)�J�mt�)<��U"�Jdɿ�t�U62�$���ů���Œ�-��M�8W�pc���C�����]��9�>Iݣ�~d�<�v۽�.n���7N�8u�SE�-+�:Z0�s�L`b�p��(7h�b��O�3�N�	 ���4�d7W�H�}'�S�E��v�+����W"T�z9. ���`�|*�]�Q�h��E��ٚ�Sq[������qu��i���o�&5݊�j�l��!8z�[�T}�Ʃ�1Q�v�JLq�J�����S��4H~=w�S���4�u	������%/ݽ���{���c����dϨ��!�v��j	C��@�uU��ꪱ��T�j�7zyZ�,l}<�+ܘ�s}��Xݠޯ���n����MAt�����q f��7z��OG b{d\�l�,F>��MW�s��䘐��j&V��ڀq���/��������W�����+�JG�z���¸/�f�5q�ih�I53�AA�U��{B���^�xpk�3�]L�1ԤI������U���2�)��B����p9�lS���V�A�:H:��bb'��Emӕ8�b��t����00�u�3���ұ��W�Q��k����t��p$$�e9n����/�k����2?MpD.�n���a�w#�U��I۸y$�oa�P$�ZM�<�̄k��Ef�F�{u+m����T��~��\-NS㺝!Ľ0E�M|�J�� F>��U��f�÷�6�#u⡺�L��Ds5���|���9��&�M� �b��"x?�G��o��G#:��yM,���X�G���n�)�^�E�ՍP�5���2���)s7�b�;��J2�V��=��[5c2ڨ�Q�mF���.hGR$Jw����qF��Y��9�h���⻫i]����f�I��D�CsX(r�oMJn�#��-����DG��o8�u��(ì芒���g���c5.�%�P\�%�U�R�D��]uƢ�9�u]9��]�6iAE�����
�T�(1�b�핧y̆��
��vd�b1��"�0:�.A�������l5=�I���OT���f+�]Q��T�40!��!p����L�ָ4C%߻ޯ\�1/V��}ʩo��]b�:�*���?5�T<+�*��(���M?7һ�d�:�����*�:͹�
vo��(W]Ԉ���r��f��B���h�7s���m��x�>c��Ċ�7�}ld	����T�4Z�JmW��u�Q�f�̟L(>����}�38��?7��]��j��>�y*k�d��z�W�_:�6"������'g��DP���ݑ�&�㠗���8.��1貨��:�UHs�����l�y�v���&V��N��p��@�#���P�B�*e���TQ�CHk��Z�#���iF:����l����]�<�p]�c8�.ʔ]3@b���+��;Kt�G»>�|خ�Yl��݋~6�8���uʗ�{%�
�`�9$V�b�Rl����v�":��/��F�-�-��M˃���`sf�I^\⨠�.�,tC9u��II��Y ��͝Ʈ*��e�\Of��9�B�wE�f ����,��վ������.��߾������s_��3I-���{D=������W\@�(�#Ĕ�A�Te#݋4�uf�q�ᜋu�{��<�~����_�3�ޛ��R6�;�����Hzk�(Z�Tv'h��g���+�����(wOn��"۲2��uh�EӖb��cS�8��E��R���F�sԐ��Bq����������pl�r��Pۨ���"`ٮ��r�L��G�(s��H�u�R��uHΉ��0�p,.�<>�]L ��e�H�엞O5�šr�z�$��w�qW/*W
�v�U=FY��ty:Y����]:��q�����W7/�uC���m���J'�r�� E��DpD��/**WV�\�ȿ���\���JE�z�[��+�, �e���3C,�?	��OW�c�cB�|h����m�E����`���㔦���+�JcEneG_'w�5:ɱ�P�o*��{3��#�����\a�ڶA�Ӥ����>��}hþ�@��L�u���S0���q\��j�'�b��4u��Wˇ	]pf�)wUŽvHa�[�qm��n�_
��p^���a~'���2�����ٮQK8�s�#�2n�g��dx*,�0����,���'���= �{}����1����k� x���3��iA�}���mٗ��ƚ�2���k���G�D�B����H?�|Mc5�ʆ,����P����iQ�d1�:�q
g��
Yc���t���k��tRp��1�s:w�`�a�:"�k�R�.�|���/`�,-�I\�)�&�"S���.!����<n�%+���'�0x�m�&�f��.c[�B�*�Sh�U�sRE-�n{m���pc�V_�.ʑ�x�n	�;~��c k��L����잋��� �Q��t���<�{p���t���Y|&1���F�':�썝٩8��R���e��6��<(MBJ�����某�y�\As����q@*A����@�( hA�_����S<���NX��-v��F�:�ƨ��B�������o.�ٳ(F�rY�� oQ��0��D��̈�(E-uÆ:j�45�ózQ���sW6�B�)���wB�q:n�~_:�C��E���i)����.#�BOcp] �n�=s&��䣺 A�j��r��c%78���MA��A�qH����9�ե]N���DvgT�̞[.�.Z��	�����P�q���Lz�������Y��U) �%�m]���%eo�<B��:9׳�Y���c�T�������*㶉!eC��Ǫ�n��R��*��D��[n�N���c2��"��u�w��#�^7L�ܖ�:�W����&3yT2ju����8\@B��UH����� ��</N��*:�mk�`�Vkx��:*N��;��������QjS&M������h�L� �Ok�
;�ۅ葏\y{�
�z�l?])�~b��u�ㅉ;�cY�����s^�G�ؘ%V����3�B��i�6���ATf�\�I�͔�4߹���U-�e7����=s�S[ژ]�(Í���A�Y��+q��C>쪰��;��4�a�]�6ƪ�mw\�d��?!��Ƃ���S�1����9�����q�����Q�?�+X��{Ԍ\�ǌ�O��	x�Q94 �u�sΡ�r����^�u���i��}g�莩.����3���7�����p�|��ڷ`�*�=e�V��)�_o�����3Z��TG qF}�1ߕ+�;���ͲI�|K�A-��]_���5�~�|�`q�)�L��n�ݺ��MPɉ=��ܽ\���� �� �|e�0
�=<2��ʜ��&�k�>�|!��M����ꖠ�u�:���k�t[kU�O���X7�|��س/Og)�[iͦ�ǻ�����	}(;@M��U�T*�RwB���d�ilOe咶}-_�6l�U�z��}r Fc��|���:�j}�m�����O�o�i�Dه�L���!�[�U��GBX���X&���>}�a�K��[�Q�ۙg��J�W[�Nأ�3oz�s@�j)11f�tDT�Χ���c99vwD�I���\���Y��l6�\�4u���s�f˝��M��Rg1�v��{x+V����,��CY0���B�5��Rc8.\J|u��c����%b�;�����V��A1��01��$��'f�h]�����C��p��J�]�xt����U��,�qPg�(I���֪k!�ÐU��D�H�[�1��V5iR��4��:���ՒuS,��8����uʜZ��&%x�&���n�͊�:��Mⷓ���H�JYId��k �)�������3
�ͰA��}�Ol�]]�e�ñ���.s���o�^�O�"�b�H����B��R��v��'4]��:Z4�*�i�Y�;�G	n˸{~�0#��]�+�X i�H��q�ŀVwv**��@��4&�/�H��,֜}2�aB��9^��P^<����T锹��k\Y��{�Gt#\�X��Ȗ ,�-�-�� �[ײ�#�kz��JUgY�i�����s-�.pGs�ն,���Em+.�=����z<�\�RȐ �E��op��-��+o�+e��ǞQ�~�:4K��\�ԗX��T#������� �D�9�>hub�U��-b�\�!tт�Dh�z0�܎�7�����-�oM��f�Ϊ�Q�ï��ˀ+۽UI���-�]$u��V��om�e����:�3ed���en�{u��O����T4��P����ɺǋH�k�r�U�'<$=�
���Û�wv���2iB^������_S�gH�����­�t��@�ȹ&0`"��3��q�kK5}F���BQ���cw���Y�T��ҭ7r�T�_L��l��65���a�׫���� 6�*�}��V4�}�Z���3GF&n���y�4�.��CD��c��s��\�M�����ӫy]�'��V1siL$��t�0
.N�M̻�	�x�M�$�(�1���;y�fPޭ);� ���O,qWR<3��1�-V�S�g^�Z����a���кЕz�V8���uP�v'P��eS�N�f�f��4�a)��!��e:�W�d�	�[DQ����2�����Ak�&9XZ��ǁ#-�/-��l������CPQ�3��SA���а�v�[la`��J8�Wz��&M]ܾ�A��g����v�p� Nцu٩�s��wIג����l�[�S����Z��OE �}T�UHU	JQH�QBL�CA0�KB��4�SH�� PRSMHU(PD+�(�	CB�R@��HPCHR�BP�IB�T�KH�!M
QBR� ��PR�IBP�@U- P4%)IBP4 P�� P@RPHB�"4)J%*D�P��ҍ(R�R4��UPQB4��@��]�w_W�����jB5��k����ơ�^AQ+[������N�d�J�4V��s�C�'AY)-b�L�H����o\��=o�U_U}_V�f0ў��n���;��sX��(B��z��(	�{��0��W]Aw
�p���9ækj[�ҍ-��M�ϟI���84����$�C��
��i s*�f*9fC+_N�U�5����늹nㅩ�|w[�8�{0F�!	ȅ2T� #���s�p�9v�ZV�
��V�{��><��}P���9��ϋ��nw�_Ϊ�g _��8mƟ���*����,���$X������)��oP�[�p��`3l�
l�U�ɣV���D�${-Q��[�B<yW�xL54��d4tL�p�vdҔZ��t���B�����T߸m�Ȇ�pj�|����.ۨ��m�8e����[`U��P���秲�1ȇ3I�MG9��Iu����J;���T<+�\ڰ�>5�{\J�qKjơ��Xx%2�tbt�s��s+��D`D�a3gv����d�v]H2n�W<{�ZU��{�ٸݵld��X���j�'o����~j�z�5��e�A�6Z�x�)ո���Os�t����N�3��w)�p�_/lݫ����T����S�
&�*�]pgD�1�1��a�3��S���4�h�-a���� �LW5;�!��*��f��!�]
�aeJ�@wc*Ⴇ�R��ZFOi�osy;q*�4�wm���������K&o��ˌ~�����[������VE�kÆO��K��q�Oa�0k��F��ڑv'(�V�F��L =e^g�`�%H{=vP
��D�N���t�Y��;��S�4����lŧ	^�,;��P��҅�S,EFҠ��4���6�M8�4n^��5����r��g��L*��iqb��ڣ�x������|.υtj�4Z�Rٗ�{Ԣ�1ݴ#�w�	�2��m;�鸕u�E���<IUc��IȮy�i���W�n�zvv�{��%����J]��C1���Z^���N���H�3��f_J�	�,�^Z���� Ɉ���}��㐭���2�q�3v���#�-��x���߄��L��|��^�a+մFi	���0V�5п�ep�N�1�l�r��̬��j��-ˏO�n�Fޖ=>/�"�����3�0�ׅ�B�:�l��8���v�HJM�N��,��OZ5�r�J�\��J���t��"鞆����ʪ���ۖ
9���8c�(���.����U�9R����趯���]s��ej�(I�e��;Wq�0 j��U�k�!��W�i�tCC�d	�)��wM����������!���GZ���ӳw	��o�w>m[�ɵ�fC��r(�.�foJr�.QK����������MGn���G䔲\2��舰%:����+;�yQR��m�
T0�Wk!��^�V�ͦ�`��.��{l6���`',/���t�z�姪�g�$�!��~�c�cĆ!\�=T�Vf�c�s�����il$�N�+����f[�쏸�ۣv�\�ZϽ�a޵7: ħ3�(x��W����Es+Z���3X�3A]��j�^��Ga��`��	�+��"���g�O���)Qz�C�WyՉÂ���9���ҟϪ��*�a}���р.��!0!��ꝧ��`x_� <)�X�w���J�ov<���Aժ��6VC��t�yPlġc���W� �]��0�޻��b����.�v�V�*��_��)l�s�n��n���J���vT���t���O2�mV�]B���!�x�һ/�bѡ#KU�,�s���a�ڄ�uz��6.�GPd�ri�;K��G �uo��x�%�U��K��Z��`�4ҷ��΋�0��*!f�p��r���@�ʽ�v����T�qLT*BL��jr����ո�l�y�1���@�>���4�J��8@�u՜#�w@E�XF5��w���j�(����"�5�dUk��+P�t�h�]��f|��1�l��JgP{����Z�`��FG��	�W�UU�������=|��B����K~<���u�&r��j��X�q6���e3ד]�&�U�F{�}��uº��(����@yP5�H�M�B*��݌��V&QoK5�b�*qj���R��u�M�w��7��
`;e��S�3l֏e-J�g�GT8*m][��7!s�� �QɫC!ˤL\0"j!7Z���W5�}�hx/���A�����]���l��jmMQtW��\�F�d�ͺ�^?  ���U��.��K졐�@����{��d-/���)V
���v��t�)<��U*ԦL�����6U'n�mu��.�w�D�1G$Y���3���~V*�7U�㮝�o�J�_y����c���mzz��']ͻ�<�� ވ0�`[�}\�	�S:9e��s���T������r.�}O���|�7������N`?t�d5��{ .5�`m�Y��;�]���ƧP��2���s����^�Օu"肋�faa�-W�J��F�>Q�O��y¥Jݦ�ۗ�oyF�9ء̾�73p^�p{��wk3w�]1�~�<Y/��-�C�n���6�8Kcgݙ�!E޶E%9C*�}�q�$����wk��:r��S���Q�iֵ&��o�m��m��Yb쑻'q���a���������x�Q�vv��3+	�1��ȸ�u��X�}7	���x^��E��&�0��O"�w���4���C�uL��sѸ;.�Xd�y��-��+s�3m��8J��:Trl�޾����`�%����T���j��_mN\W*z�r�Nhkb�k:g*�wi�ÿ!��u�
<[�A�W ����=���:*�������� ��2���^Vte9��fXL����p�"�3��(B��c��
.��t*5G������uh�z����I�a��i��N�sN�Ë%�F���P&
U��S�륂F�rz1+���f��蟐-}qW��St����!��Cق6��
�<���8�_'꾖��#�o��]S(
Ⰱ�-�_$�"�s:!�M�����D��N.ӻW�������������E4{a]��p1��[�َ�.q��{�˱��^��H7<��������!��:]�u�#��*�A�<&sWi��懯�(55�yʶ������n�b�p�Ul���n#o���2 :H-T�݄U� y`���n�fÖ�t�y��oP)�W	��aIs�JZDY��`�Θ�cl�Y�0�+�ΐrk��'�7:T.Y}��iĪ�wur�L�t���R�U�>��胓�E�%��2X�@^V�$Z�L��rDy}b:H��u�r�6�3���i4��S�I2���]H�W�ݪ�&C�����,���r�U���?�Q�X��;i�4�<󎈫C�CF	���ULE���fn�;7	�P���XQ9P���l�P��G�����$n�c�U��L��}�ټ�V�D�X��������~�� ����v��J�t��l�;6�����Z�X?��8[Nc뇑*k�d�Q�g�5u�URbF�g޹�ě�kO�U��PԜ9s(e	_B|���c�g�Wץ�/�[ǁ�8�일�P[�����E85�7g<�SN�Я
��\-���ixS���{�=�I}%�!�yܢ��z?��+GJӔ�e:��|f3�R�F��4j���(��[JB��6�c�:g3�&s�FDS�wb;>��|1j�m;��W\}$�_B<ITg�k�d�(�U6uj�ߧ��4��*a���q�j��T��!��h���{�#o���p(�܀o�3�5t��=��ggR�q�-g����ƫ(�$���w����'.[+�Xh����$u����Dؼ�wo[u�p[m>��5ۮ�v�^�%7�|�پ���؟`���u�����[��
�k{H�tC��Sp~}��}��+�ʏe�Q�4}<@���V�V���q��1�r�#�"۲0���k����[f��/k�*V��(�<�H*����*�\j�p�T� ��G7���1����U��L�Y!��'-]�4-L�k�REF5�蘿�*���J��ﷱ���͓�s��n� �6[��h���ԫ�:PGt%S�e�ϑ��[=.w���zM�=�oT+�9N����dx_�3�~IK%�X�S���ڀd,!�ŵ�/H����S��T�j��}\�4�1�'2��os�a�5E}��L�!��V#��~�^'G�BĊ�}��Ř�x�g�cð���?V��{���{Q�8#�9;�:��䱔P����T�,�=]��xk�M8�Y��~�^���r\?U����Ѩw�*s;��g��y
u;ճà�5����s�6x�Ug{oM0Y��i�5����Գ��P������u׆dWoy�����ب��q�ޝ��^��US�ۊ�9k
�UpT+�x][W�]`x+p��5<I��e�9ȝ�x�?
�̕7�bC�a祤.�����Q�0Q���&P�e��nUHc�,�u[��6f��:Kջ$-|�v⼺��D��㽱7i�!�vĵ�m_I���uty�nJ�3p����N��*��N�\��A���}��ﾯ�F��}����V=<�φGΩ��O��-�iǹ�#�w��w����-�5���uY�x���R^�P��C[rGaԧ\[�![���u����q��F�؛��c�xߔpXS�����@(�B�w s���a��f�g�}qg3/�����o)2ѥD����M{�	1��W���iq��Ta���4��Ƥ��某�{}6/L�&v�56-��WQ�8��`<o���I@H��`4���L�_K,p�n�EӘ��ȇ3}^��;ð�3Ջ��~n�WX�x��@��<����@�\�婟H�P�L�m��8�Nz �J��,n|�wo]��T�� #�B(tai4�󌚐��~�����}8N�Y;/����T�y5hc�H���MD&�@��[ȫ0Y��?.:�ue�Izr��x�A�}π�d:���W�u���&3��%��p�4r1`J�@��b��+���n�WX��S?0E�*~����r�Gt�7	=���Q"�.�(����la�ٚ�ԙ�V}�@a�x�$e�|�����q��Yx>m����ٛW]'N�(��A�B=.5� �AX摓2Eų�
����C��C[�*�&�5�{�JH�#�V�g\;�0�v�gq_QP�-��P�P��9��s��������r�筍�EVI_r�1:����f��?�]�#�RO7f�����}����I]���z�Ϋ�{� �c�Wr�B�1a#
�U��iA��'s!�vI�K�Xv����]��jt������l�+q��uY"���y���w�����SFJ/.�;���8�l_^��/�e�)z�����&�E_�,���q\w��hSW���~s���9g����̤OA� ؎��E�S�l��c��MW�s��䘼�MK���lvO<�yT�V�a8,��̪�qN�����+�Xd�Д�/�-��+�<#6�H[�P� ��ϹB��$�^�&& ��L��iz*���Ӯ������ܨq�*��u\��>�7�06�U�q��s��౐�0Q��� 뢸�pt�p-kҧ�d�	�C�@@�R�떾�iZ^�(X@#���k�Mc?\@�LB:I���q 3�N��1뱻n��ݭ�Y��Z�.!T��᭦�c�8z��1��N���%�F���#�3�F�jt��ۊ�*�!�Ɗ�P{Mߡ��������>�[�e/z��:+s�u.���|�%�B���{Ճ���Ws�0T��]\�{���SB�\HqQUoy�m���t��kMk��.�pr�5����"��ɂ	'U�?W�}�UVu����=^���}�9���Z��Ӹ�p�)��n��m��̄'�R5�݉��͓�hv<͞�k¨K��Кz�Ȋ�{`_jN�9gD6p���w�A\:-���w��״�G�V��^ԉ��2+&�?�!i�y�S67�����ܛ��8W���B^�Dz����t�9��p\����Q��)T�Џ�^e	���<��e��gd|�嚶Z�uӠ7�ӝ̣��*���WN�{
%���1|��ǈ��(ڬ��|����[�l4+�kT�k�w�ӻ�p!��r�Fx�eV���/�b�(Mw�܁�$�r�lΝ����kU1��fm�Ps���U2#�XdK/������=�����C��u�ђcX��L�fڶ0��LCG������8b��OY��]�ćX�p��S�j��T\d���O�e�2Qó1���䩮e��c�D�hn�w��=�Ę�x��wL0{�"��NG��%�iy�_1膞�������%��ï�{��f���f�1��w(vbc�M҂�Df�T�ֱ��e>�3�`NR���؏8��1��jm�.��%d�{B⺎��j�
�]Gl�IrJ��*�׭����(x�I[����֥���+�C�����v8��3�4S�b).yh	��d0Q�<����̡(EKh>N�á������Tq��B��/,6H��:�j�d��<{�v)�
��v�^j+��H�D��M�6�%��t��\ݖ���%�}tZg�ʲ'E��i���X&�����x�fKZ�-@�_*9����/�����B�����]��Cvym�d����Kb���A��`[�2k.n�GK[���mh�)6�y�|��.��.
vH龊e�K"�`}��h뵚`nk��������U�C^�;��	�ͳ#�/��C��N��/M��́�lro-��Ţ�Iۙ���t��PQ�f��>t�q����r�h���d�״2�Z�2�����eGr.�[�TIU�h����ԘBN��;b���3��
����IہZK��J+��V<�lG�T�f�w��I��e�(C��)S��sfب�ވ[��>��.i��5湕+����am^t�V�*ܷ ��������@ޥԄm�rn��c�/Q��y]ѩݝ;�����`�x�	W,��뜳��!��$���s)�Õ;"Y]Y W����+nb7��Y����U����"$R�]u>M�Dt�v�K��Gm*���@�oK�a9ۥQ�Q���K_sn͠8��hh/Ri�otX�]ۻen\��ꓷ�Vfu]"��w��1�:|/�����eca���-Z�#T���U1=��VȘ�v�;BԾ=E�"��H�|�=�g\.�
란�j]��i@a�K�3GK#���.��̓6X���ѦMJy�4���q^*����o`�/P=,h��,�Q�D�o������RQ=S:�<ZjJ�;̎�D.T�5v7+���1֕���G��Ha,8�\l�^la��k��*1m��6�����.`o�ژx�K�e<�b��#��Xzh=�ӯ�����,�!�ɿm���|��:y�4P��JC��:�.y�YU,�9�����X�*ټ���-X[�@!Љ|��*N&��v	Hٕ��r��.P[�G�U-����$k.������E`�akI�pA���C���@-�F�}��r�䶇y��[pM�!�Q\ν�6na��XW]
)�iD�����흲a�7�u=��[�1�����i��^'�5���wq_Y�r�qJn������a����y����u�����h�}¹��F���	�)΂�T'�DƁ�H�����6Q��񹲥h�*f�r�5z���i�X�c���wWɩ`�+���qgm�*9;������Ъؖ:����G~y�gFw�ދ}~�@�@(����h*����*��)Z
F���
JF���h(�)���
 �J�Jh�JZ
P�*��D�B���F��F���R`ZZZ
�
hJ �h�(�
J�JV$��)ii���)F����X��� �()F�
A��  D��  7�`ؽ7�M�K��.�5�ꅭ��S�
���|��36�<!��v�f�0z֗��:g��X��.�r����UU�}�����{,�vxr6k�_
,+m׮�tW`�<>���=G�)ɓ�^+�3�C1�9��R�鈶�3�N�5�c!���Y�+G��uEG�S~��s!������x�OnQb��q���(���aC�!��'=7*���Q�G��Y�=\�^{X�[F	^RW�Oh���컉F�-��R��9ƽ���T����mO���[L�ڼL���܀;��>P�T*C�|�t9��vW���ez��{��Vzj�H�yy��i�p�E{�Di���w/��=�\5�k�\;>T�O*\�$�S�9=�qbv�wxIܦ�*����<�o�îH�|��B��\k���ʴO.�&�p��v��Z�2�e����'h3�[;!HV�t$3�x��GX,XJ_3����n9��l��E�A�.VC�=G䔲Z�X�9����v�B�`��iUzs�'5�Yp{'p�0�Mf\!�s�cUtp0��4�Fh`v~^��SQ�.T�P�i�Q\v�R;��(��+�6�C��Ke�&n�d`sC�ڔ�eL�h�N�w�h���C���}�VC��-��t�OQ���롤���b����g-�aV8��#���s;��C�8y���:C�u;H�D�`����Z�G�r�&��H�Ae:�3��|RS7������jt���
�E���AYYX��8���ww6���<�hT����Rs�����O��L�vڿ�L���pp�lo��Ѵ���	қ�=S��K�]f�Ƭ/���Ժ5��E#�#��ǹ|K���<�%W�;9d�҄:gj!�8��V�l�y�x�.��\½���[����� KQ�+2�
K��A��'�V�<�φC�l�w_n���^��'�W�}`�ڽ�)jJ��X�f�f.���D����Qn�K uPb/��g��طLBs<Ү�P�*F���4�On�*#�t�L�+�9?�Ƙp
4�]r𯆈a彸L��KT��mݹ��9/�����ܫ�dǫ�A'_�x��뮚\~z�`��4���jK/�n�v>U�+��A�r�\�z��;��2��A�
<ҟ��S<���Ʌ��f�͡rt���\��0=�V��FQ,}���b�� �ߌ��ZH���ӄ��������Q$�Mu�}�FiL�ަHRR���zk��[M��c��'핁	����V �X� )��FX�H�ta�W$�=�Ou�'[62������}�(�:Ru�e��+0H�k -&Bz�N�H�-G���
;�C���荒�r���ß�7\8c���6X܄븗��p�@����0
�-'�������{��r��^��.�pX��\��ɫC!ˤLXc&�7Zëyf13K	{1�ہ���ms����*H�J����w_�Wː���Pɨm��� h�i�l�i�:/�yi�}�X�bx��H�?\����3�o�W���֚�"�JdɊYget���y��B�Mž�7<:�c�L��Uq��U��c��?E��0�ꫨ\v���7������a����xT	��(�/L�0L��B����l�`Vn/��(X�	+3��hk��6�T�#5:Ž���_8uZ�pi2a_u	w� ����)��En���d����� T^��/�e�ҧ�c!���s^��WR.㥓��6�c�ƵJ�;��*�P���U�3�2�=�&~�]d_S�l����m{�s��h����x�	�rJ�lz�z��xe̼5v�]*�z�CG�ˀ�5	O2�m��,��&�P�z�XTH��ekl�6��Gm�xWK��3pBۢn�1��oٳsiL8-�s����e��t/lг���Ź�%�B��R���E���G�D[����C�R�	��Ǯ�j}l��}�%1����Z����s�U�}�SpŽx�=�]pxZ0\$��	`����>A��_GC9�.s���\qT�I�!{���O2�����Ƒ�OQY\�|+�J8-�.Z&�A��_OuS��y����.5;C�������&�b��~��A$�D@P�$��M���Fi��/d�ϯ-�����@ţLs������ʴ.+W d�f�.fz��*����<������(�Ǟ#_p����*�;��)����C������BN:�L�b�8N7��-�3/���@��A�V��\zu}P���|�tCg ��
P�\���٪�wY���������D�$���'� @x����e3cx�K�ɑRe᪬�,��w�#*q���\��D���)V����AU���s�1��Ip~�m[��%æF>�*L$�-��M�����
�����.� ��GcS�в���q��N�Ըx��m$�_֜3I�;��F�#��z�7U9u[s�jSt:�W0�p���ǆ�TUI`
�ƻ�N��<�>J�i�<W�+#Ӻ���W��Iq�$ΚWM㭧E��Щ�V�"���\�$���s���w���3�aE-����#�/�ufcT8��L��>�e�8ݤvӝ�+����3����U�zw2�{��s�{X�/;�Ny.q<�vop���'�V됈k�����|3M�+�v�_^�4K���4Ԝ�Wl�v�@���\��w��m�v=[�x�&�(Oxv���)�x�׏+��K����S�E�^�NSV����`�Cf������c:��\�e�&_o���9fmb2_��6j�˔#v��W5��dK��ǚ��x��aJ��bahn��m>��|�+��o���|;Э�%���A�)7<�M�&���˸V�_�[ǡ�OC�M=�*�]�R�s>!ܕ�դ	�2���J}}t]D*[4Ry|᭷�k�6GO��=#ZU�j�-b�}���_oa%W#���{}3k��:Ϣ�Œ͎��a��ݠ�ƴ2�U)��
{��0�KE�0t�rE��F��nJl�H�l��3�t���c՛�wG>Xwen��*�����>ʜr�un__+� �E}��a�Q��3(._Z�mK0:���ϥ]cӪ�V����{��	vؕ9��2��qp]!p�9��e�8��)��y�I�gM�YkV�����Ͼ�&��
5k�9ڽq7��)�r�S��B���.��OJט�n{�!9'T���t��X�R_r�|� ����W8�|�cC
�b�J' )���>�U'��sy�A�'�jL8n1�7�w��J��a��v)7�������;����筵3�i�5	�ց�2Vv0�Y�|U������Z�Y�8��}ܶ�r��9��ᕢ�RQ�YT�����r�u�L@��3�7��I�����܁�f��.�����<�jS��4=�Ox�v�Z[��e��������.�p���Z�E��y�����49s3�2�E��&�k�@��"�Q���Mwpw���$�.��&��Q�6��v�wݝ�e��ș�4`E��#w4VJ���:�\����������-��>��s�z
��"����0���w��fS�"G��걫��1Y���?�g'i��SӍM%;�dn+r){f���r]	a[:�ijk��Q�e֎	����_Y�S6��c]x��S*�c���Y��f����Wj�luJ�]6��¯�&�c�A)��{�/�W2�!g�w���_���*�_I}[J
����o-�o��T�gc�0�-`ɥ�y9��r�7�����R���mIꎮ������
�@���j���ѵoT-��g-�����aLB�x(��CK�:�9�9w��fn�*m��.:Z��vDk��leC�J�X]�����,,�-WFg;��YÛ�S���ZP�r�3�.�@.�n�M?'W!b-Q�˺u��=���)~�N��Ҹ�_p!Q	���4�eJ�=��ӕг��_̾��Z��nN�5�1r�i���n5�XtC�����9�������@뒷&�Sɨ�[Q���j������j�*IB�hܣz��Eι[��~>܉n.~�M����.ǖ�ۆeb]O%Rqګ���<Pv�ʨ׆��c��k�ᘪ%�z{�!�:
s~ֱ�b�E�@�˟9SA.n�\f����[t����x�{�s��p�3`��ar�3r�
���]�g'-.���V"�,k�y�����;��Gr�x[Νm�6vj.S����Y+��C�����0�Υ�)�A���qkkZ<�fEz1�|��ީ�0��4���s�Y����K�Z���ۉy��/����B�x.!'=ʽ���4n��5�K��{F�uh���^��q܌J�nr��:��c�p��|�ϥ������'�:&�ޞ��N�s�Z��C�*��Yܕ��
1��sz��i��:=D��Ò�*�.p��jr��Dֻ��	����ޡ��!�]�V��K�ham�o���w8����姶VuB�*�����|�$�)������n��F^7�{1ɯDu�������Yx��Bi�n���⢭��g�b;�Y�I����Wb���*�R٨R�_�k\�^�<㔝7b�옝��G��]Ex���Υ�V��eKھ�2�r��߸/G�5r��2nY�M�0��Q��j�ɗ�����@ih�]�q]_B�I4��n\��yS�,r$��Zl!�/,5��l��F*}o�<7���S�L9���Io-�4���Xe{<��|J��?}�:�\��d��4J��Ƀ����_Tf'�)��M
r�7�e�c3)mv((�|��{ ���$Ɵ�`[��*����e�w9��n�sY�sH�1�T��R�2���}�nVq,���TT\�rR1���l+��
�6Q� ��%k��1>�/���!��}��S�<��qi�Τ�4ۍw�O���������
�c��Ω�\�Vz�e��Wd�<��Ɠ��N�M��g]ld�K��Y�̶�]��\�ek��Ve}<��}���kE�bp�C�s���V���7Y$:��ۣz����b6���ڝ���S�Vjw��u��+Y%m��ҏ��K#�勥��.���,���=��TOݏ�NL��ਓ����[}æִ�u�<��u<3ǭP;��W����M�[n�ؗj�f{��ȸ�և|�.�\�x�,�����C�a�;~Φw[gj
�^����j_ѵ���l�lR���M�{⳩v�76mh���w�/����׶��U��wq�'�gNT��ZSɤ�^���UAV ���kj����S�{V���=�fm2ӏ�eL8���y��������:T�KR�N>i�=�� ��ָ�y��ѓ-��\���޵�0�"T�Tm�S�ϾW����C��|��-V�_-T�[�����z��O�⯓������<���H������
&ީ=�㮋��#�;���Lrz�bwWB�"�d�ؕ�,)_oO�A��n�9�>�r�ܬ�ۺ����K��Nof4�uZc+�T�XS�ou-�r4������6����R�Z�Kj��v����uNi��]�~3ڷ�<�]�PSР~��v��ڴ����� �' �FB�g�;@�gNpM��ճ)�d��KS�ײ[���U���$�w��h�J�w�h�d��y��i�Zr�p]s���)��݋{���eŦ�}	��N�.�Z*7����I���܄*��/��>�^���J��g<���8�F��Y�M3�I'����Hz����*~@���,�Y3j����Z6�3S_A�T6e�rW9d�
�;��,s��T�J��D��V��c�����k�3���t ���J��K�[�:�9y�d��eF�\��U��e�uur��v8�������J`Mx��L�e[��)�����A\C��l/�\b��ܗ<������@k�`�������x�L�V#�go,�]�6�]͇i��7��F��\�i-n*r�e�ᢨAݘ�K1�S�%�����Ж�5r�媻����`�w�#��X��뷧�uEb5���G��A�YB�&n����T2��"���K##�<����xz�a�1��m�� �q�,Z�@u!�Su��:6��z�+�0�Z��t9\4Ff�H��Q�C�F���u����J��fрFܯ���BdP-1�4S��6A�5�O%kC�+;D�Y�.*B�닆1 uճ9=��LL��k�'�О�şr�xh`�ξ���t�i��ZtE�Z����TT��p��4`�.����0�Uy�ͽ�g=;���E�PI]��D��j��yQ!��٠� ����;>L���,=xT�IS,����κt*�@�',�����Ǹ(�=3}���\��4n��f�C$����<�2v��A.��.s���A��߭��شfZ�2� w �;���̮9N�Ӝp����:�SK8px�lVSٴ;D�q����i��ۜ@�Fέɹ0p�a�T�l�|0��4B���u}h	)˲��WT/M�,lT���&�^��d/rW,nF�ެ��p��nu��L�;@��]=n_�yo7_���y�Y��ѮV� ����w��{`�t�8U�O�[�`\�p-<�v,ܱ��:�G۸���g���b��,[X)P>�J�쭢��2-&VK8�XR��eu�dZX�gj��ɓE#Be2��AM�n�@w*.�}m_
�@=A��&�E�BkXޜ���dYՎ����D�F��h˛�(�Z�5�m36��K�h��Z�N}K���ޛ-gF�j8M���m��|;6�ͼ�6,��e�l���,���Ԗj�{���;�Ɲ��'m�f��9I�)Yy������k�u> Y�UJ��|.�-����Ck��B�L�c��tq6��D�ǽ�Ӫ��l���bu�ڠ�Iǭ�$��8b�wY\��;W/���"dM��ku��}��!��n�A�Wu��+.J��G�MZ�-�L��鋛��AXS��.֗L�����H�Lvm:�rl�ɦ홼��_ZX�u��屩V�h�2ڧu���K�c�e�ޤ�A\F�a֤��-I[������|b�@ZYx:%B�:�^?�T�<�]MP�F���S��h²�JX2�uz�:j�c��=�ǖ4V����1�����n��è��X�(�3o�;_H���,��i4��\���I�eٖ6����q+����e��yi��kW^a�]~�?�!Jh)Q�JF�
TJF�F���
P)�JZD�ZR�( iA))�V�h�ZQB�
�
b ��w�{�e��<�u{{���Y5��Fg;W`��]�O��jo5�uNx�R�P���7�'��n"A܎GĀ�ΐ�;̊���������y�-��ٲ��IƵ������%U�.�9��φ�:<������ouD����Y=Շ�z�3յܹ�ڙ|���2u���ͦBR�����h�k_��{7�b�-Z���(��|y�c.�O�m���á]�.�VBUZ��ض2�J��;Q��+��|1��7�)��v��  ��,*�W)G���;�Y���j���d�^WA��t�kot��V��{>��\��:ﻎ��^r����A��Ry �z�a7{wJ��'`��K|5���Ev8��[���|��.۱aJ��*�.]P�Rg]�f�w{�{%��KZ������N��}���u��16Bp���+�v/]��_R�������<��r�Oڣ#�B�vfD�z2�b���z�j��+��[�y4�ğ���ߏR�njf�v����qS$�\���ͼ=γ�b�.C��l20m�c�9�]ec�4=kP�罰ź)��,�蔵���Jd�1]���p/V�����W.�m�ը�%V�y ��RC.�NI�p�,�����ӣW2�u����wz�mM��b�U2�u!x.n�S��k��ŏ�n���NjV�F�:[�i.f����P}S�C�C\�e�赽��>F�U1=L�~���Vw�l|���S]��!��u!):p���/�M�M��af�"�ص��N��M�ui�1��)Dجu�RAk��X�T�ÚMAچ���c�Rڈ��۹��ao��5ꩿh�<�ku��[��/q8jIʆ��:��}�2�+:B}n�$��igv8	uM��+v��|���i>k���ޥ�����������HfQۆ��Suy��������Z���F��[�?a�b{�j'�Mb����܇e|U�;�.p�}�uDLN�hp��#�N3d�e���s���kL��m(�ݦ�OeX}�=7�\�~�%;ɩ]v�I�w��I��l.��i��Ky_���p�EhDȽWU���<�^���K�=��~C�(K�S��Id�W@�S��w2U�M�K�k5��JgV��7�*Hi��nH�e�݊�}^��FLJ����/%s}��q���ܜ����-j�R�Y,�Y�#u�ؒ�)u���ո.hΓ���xIiܽ�<`�1�軘�\OV�q��kyoCyq��ɧ���:c���ұ�� Q�ǏP��T��\WPU�l�)O.ko��<��k���:el���x�����f���
�b�s��I>����J�G��7ܱ��Y�F�B9T�M
��,swq]K{jiA��.n61��=NZ�����.�a�N��9�D)���4\�b{_�S��J�AŖ3f���.�МF&���a�
F)S�u#� �sG��^Dx�j�Ot*l�un�y|�9�2�Ꚅ��n5�7	����i�P��]�;Z�x��&���Tn�W	:��ᚄ�o3��q]y�nt�]M��r�F8j�����'^����������i�9ܙPq�6dC )��mI������>�n��Z]����L�&�{���%鵐��S.�	3��e:�^�	o�X2˥�)A(왢�rs�R�W�t�Ҕ˼�/_iliۃ�Wr�"�w�u6禷���+�Ghy|�t�mM�Vd|�+h���;��(	���[����+�9m:���I]ée�j%R[̱�j5N��߭vm�rv���J��Γ�<�j#us~ʿ˷-����Τ}N�<�M%OD<��s�;-��}������k4$��ڡ� =�9
Vc}��x���\ŭF&�J�R>�=�Ӳ$��,,������	m��������&������.��8J4��lR���M[�}AWԻh��9��8m:U�$-A�;�	f�;�+�YK��_�Cyp��&�r�o8e��ꖭ@���ϒ��5�z��;��.�#1�<��m��;WsD(�x������y�����zJ�:���s�O���;(V[Վ�ѫ��U9��-bz��臌�J��﷧���eiN�U�лI�뷏�K���uÖ��9����9P��"�B��h4�po}覑�ñÞ����"v����|��Sw���.���.m�X9z�%�K$�5�4,�3�)�@��o~6� ;*������؇M�;o�����es�Y�}&(�u�WOq7�"��=�GN_k�^i���*3$�ܡ+��K�:�z�(p�߻&��[�Z׷��ƃt�٬Y�wJYė5�*��smA(k<j6�5=Us���k7�n{j�u�~���n9d������H��$�X����G��v-��x�U5�$�/6�Ч�VGF��v���N:!y�ض�{j����q�]�{�ͭ�$��.g����D��^��߽.�л���*�zj����l�C_WfU��ɪ�l��,��ݽ�ض��Νɝ��2�p�teڧ��[ou��ģ�\��$�ڣ�v�\%k7�c?>SV�:�yz�mym�ʹ�
+Ѫ��q'Q79_D���b�䆞|��K���v��t����|dN0�6-�q��p鏃��E���j�kU�lT%��DSM[����'qb���3;��i*�N�P��Eh9X*I{��{yʨ����±&�o
��ɮ|Z{�VG]c�@��{{���i@ǡsV1`l��q��
�*z����b��Yܠ��i"t�����ػ��/��]�o��*W�m�z���Z�1�k;C	ː��w��nUݨ�g3�fm
Fw�Q�V��W&{0�;����!{t�7��t��Ը��3%)̽�T�r��.;�ۅ��p�~O��M�	F�AP`w����J��J�d���?C�߻<�{;˹{�����O�����f�c䓦f�޻�P;n���r�LP[���-|��mc�=�O��|#{b�oV^7�՜��Y �ϒ�S�+]�Է��ri[:ݳ�\����A셇Qgu��Ǔ�թ� ƟmD��������ڄ����r!edɀ�ʓ�W��WZ�{�TdB�
�>:����,����on�S���q]���vV���@��k�'�tD��o*��ڿ�2k��^@ݯF7OO3�ky^l�8z��ub�I��{������1��}{�Ι�������vNw0�<߳[�ڷs���èy'+沺l��4�WwNd[5�*o{9��=A�6�~�3�M�|J��|�5\',��,�����z��Lu�3��z�0��^�/Z]��d�B�̀f�x��d��6|]ӂfS��V�X�s�GIsݑN�\��oQ���1��p\��Yt!�@W�==�\�/]=y`��R➱��nX�Mj��-t�ci�	�oq
�-����ݩ��p�p����<����}��C.���I�B�"Wr�|�'�V������r�Hڞ�U�.�����c:�(���Z�I��l�Qo�=�s��k��iD�7�	�����ޔ���̴#�­������HĿ��оb�Yp�}n�T���p���\sn&m�.η=\m�EvS�M�D�2�Z��kyp�7��8{I�����$٘�d( �㳔g(�8=t�i��uP�l�)O.!��އ�8�IC�c���͟g7�s��E=T,ﳃ��WßW݋�k�r���م�����d]�egr9isi��T�������+��k���q�!Z�Vd�=���*3t�=��FM`{��x̹�D.!u;1���vh���l�δR�gv���� <aXw�Ҏ�Ά��/V\z�a�ǵ<��3]6$H�Ċv�̊mĄ�ګ���tL6���fdv�f��J1qV� �cN�=��Iŕ�>���N�7���w&0���Y�6�(8UK�	�ϟ@*[B-��%ۍ*�]���Q����d����!��-55p�F��ђs�]6v��F���2�!���I1Pۍw�JvG!���.�]fM���]k\@U%�î�s2w^+�I��Zp�n3y�\;�Ln��[�M�:A����V|���ȃ�͵�/k9'9i�.r.]BPʄNL��U�N]�ꝭ��6�|"��fsW�um��}������}c�]j@�}&x�g�ڣ��}Gk�ͨt��y�Fb����i�tXdV��2��=�AR����'[��*�W!�E\�|�Mv�o0u
p����7��=y�6���=/D}�{{�dK�Yd.���gu dU�g�baZ�87��>I��?�mt%ce��ب[��SM\:��U������ˇVE���ۊ�6`� 򯤾��PU|�R����O���&)n�3C�hˤy��zw�AV��	h�Wϑ	>�����*��5'���*��VÇu���Qٽ;Qħfh��i�V'��q��ZE�m�-�<�#�>�r�1�=�5�H1Z��QR;���s��٪���'DV�k�����;ut��k���4v��x��@�Zl˩S)�@f��J.�!R�	��r��ggS���-f��:���ꮗ�yNdy{Ƭ�]��z��*�&��>�g`��շ�W'&Tf��/���j�q���T��
c�ޘ���0B�G;b�j��ڼ+��9�4�Z�y�J�׸�h���|��ЈS��u
�EL�o]a��OPf�&���Ū[�j94�|��+��EC�td�W4�T�����ޱH� ��/�M}+rj7y�C69s5��q�ʚ����*���28�i���ے�&��y5ڶ���mL�)��ZGH�IZ��j���.ǜ�8xa����/�����S1���;�w�,�u�;ë��X�R��OuW_؜3P�A��r5�v��eU���:�%K�����$�5Y����-ɧ�K�Z�ZϟQ��UD*�u�fQ��Tn�j�u�k��ޭG�ܼꈒ�e�ڢ���vZ��m�gM��ˬ�-�AܩH��p��Mͫh�w{��sc%w^_�{�uzϣ�N�$��e⢇$��=�εQb:��9���̝�VLǥ����vlE��N%V�0��<�9v�Bo8�Ԍ�%�h{ǎ2�,#~YEn���
�ܝ,5�>j�Ss�S�c�!G�63�X��]�q�1���A�5�]�ܰ��ןr�K���P���
�ca.o*uda���	�8���֙��~Q��=�4}5u��>t��o�1���%:n�s\����&����}��
��4/�v���-`t�t+~��ٝ���@��ky=�����-�M=����XR��**Z�d,���J�Ry�Z
�wtR���S���k�5�s�7��v,1�e|�M\U���q�pv�븎+�k��������y��/�����J&I��S�_]�q�t���0R�_����o�M+f��N]CL�؛��&�g�n�	-��M��B��]P4��I[w�y�-��tT���9U�ؗ�m�Hsw\J�&#����+\�����v[��ܾ����nJ彣���8Q���R+Ω]�d�ؘ�?<�q��Y㘣N սye+�q��+iI�K͍e��d��cGo_>T�)G�ݨ�H�HͶ����\��2�e�V^���
���r�F��s3�{uӨ�L�������8�|ƻ�W���3i�O���O�
����b�&[ 	:P���*���!�a\�Y,�)�s5xS�_JU����u'����r�s��T��^>-
c2m��M�T/z�q�6`�A�u[B�H�uj�Te��/�kl_?I�̀�q��`ٵ0U��� ��:#�x!ASKU�s4V6��{���S�۽�M��Z�����bmq�e���:j�q��R���G�g�$��uE�^�C�$��WSx*{tJ<���y��i-k��&)0��s�'�v���A%�ܣ*h���1����y;`I�&�"*��@���y�!Ntu��x�ǆ�]�:u�&\�%����p5"���&�2���K�#"�/�V�{���j���4N�nP�Vq仁�iYȫE��۵(�ӄx��\=��!��:�	cU�$������9� ���̾4�9�-U�S#�e4�P��L�@GX3�ӫ���t:j�sy�8Z�M�YÛ�����`
W��7R-C��9�u�H�i�hTi-��TD8��2��\Xʀ��C6Nc^�5���g0��l��GCeJ_<�u*5��m��}өLsMe��t�QV%_B�͛�:�S3��As : T�Puܺ�\�S���|*��v�f�%ӝ��k�x��}��O�ٱ'�p�H��p&�Ï]��Ӟ]ہծ����.3���	d��Li�`乼jj�]H�A8��U����t�un�9a�{N��j��u��u�98 ����v�sD��]0�nV�P]��e	��ݲ4��xf��'ׇG�hgT5�.��s;)#�%2�]2��۰�D�A#��x2Ę0��>�{V\:ӽ�s�ޫ=��ʉ�� Y�aHw��hut�P�Y��)B�ͶY�Ӑo�T���:1U�J�N�|N|�uɨg3WŌU�n:�:�l��k����\�jp%m�P37����rn���u6u��f��qb�D�V�D/�ĭ�C�L\���[b������ƃѿ2c~W;b����E�R���Ft�:NP`ѽ9J� .�����˔��A�q�������� �B[��0��⻍'�nL���X(:ݜ���k �����}W��Ea-h���wcN��;����`0Q��lr�`e��=b����H����FZ&�qe�S`k*b��
^��e!���<0��ݧv� ݳ�$_<� �l[��U�8p���@@�h�Tn���������-����fi[�swQ�t���h��y��E1t�@����ʝ���_2�,^�;�n�X�|E^�.�() �����T:�
�)A2@(��rJ���
@
�����JE�����JX��i��Jr��;ߚ�;]#N��k�:��[1��Q�f�ڳ��1�GgP*K�Ca���oMK���o���G�izy����J�N"�
��g��t�T�В`�n5��e-�!}8j�_k�6�{%�Z׽�@���
Sժ��Kku�.�W	:����ɸ;��#^?kS�)F���kL�Cޓ9z���~�9!9�ʧ<��>5=�f18f�yG����
)C�D*��ۓn9��z�f*����	X3�5���jO��Y$]R7���hhs����S}:��w�p�u��֚�Ao���}���n+�(��g����V�Mf��vq��G�����TW���9�g��j2��u�f{��hW.l\KO�lL��mR�=��ɿ9V	<�f�V�3�-{O����d>���-!]�,��O��=�*��aU�m���'N�!��f�f��rZ��k��V�\o-�o/=M<�7�R���堘{�2GJ��X�Z2��"��R٨R�\4=�꽃���P�3�;r�i��J��U�K{@���գP��]�oc�F�+ys�ʫO�zd�e6^�"ؑ�zQ��t���CP�\_i���.�L�����R���On�EWTK�z1oS*�;�E-�١��ra�B�J#y��u>n=<7�
ǧ��r�YG.��XS��I�	wd��T�v��������r��4����"NY~�c9Pꔠw��CKE���Q;_p63%P5K8�����ڶsZ��l^��(��F�Ϧ�R���on*�Чi;��OO5�3a.j�|�x�_�gg����\Ej֕����OVo=X�gIN�5��C}S_$�v�hTbvF�ܸ������E����n���ɬŽ�6�jӆi7��Ft��.:�S�l��I��[�"wF�om�g%�X��)9�������h}�>���&k1�����7���-��9ٻ�A�n��'�{}�����k��k�����Zr�\l��I�5���z���}�P���S-�nD�Sx'r��l�9y�"���c�eJld:���fƼ��!l�J�P�6x<�h���D���gs���j�����ð����E����W���/���,˳D�u�J��[i�7�y�;c��A��K�v�9DgvnH�T���9�@��GR�|D��AG�f�:�)�aj�<zq���n�y��������n���Y]��&n��_u�#Fؗ�b��\jC�%��ݴ��ͷ�v�4(��;�'�-��Ibж�=��.-X��B�os�i�<��AMl�9��ij�ܹ��N��y���!�m(*�j�c[ˇ���VL�߮�<��=q�������\|�XS��6J��|��);��)J�'�S[՛W�t�.�����Mb�-P]�87��е�,����9W}�w�l6��gY�G���9�_ʟM9}������ί�3��+�aO}�&�Nø/S��,V�w������p�k��>�_<g˜F�әIƷ� �B�,��z��}W�e�Ojˎ)-�ɥ2�;������.xe����T�Ԋ��س�U4/\�Jܝ�kxf���|�� ���.��-odn��%K�l��@�rs��Qڶ���օC<�D�m���T]��s}M�Mg�f)C���EG~�@���K�V\��ߡ�&��gJA����iK��8Ļ٩��S�r�zf+���n8>�挕�5Y���"���Q�v��R2ݪ��]X��`W��ަ��p���7a�zbu��Sir��/�M�I��#7���7�Z��dKk?o/=[sx��:�=Y6{g����w���ᚇ����W���F��Y��*�Yڋ�Xi�J�Y�ѷ~(��я5��r��%/��5���v�1���
�&^�nU��Jy�z\�R:�{��V�ꚽ�=��g��?t���=� �II�A�W��~�5��r�Jc�b�Ć�|��X�l .�t�w�ʼ"�p3ܽ�����gY����
�ި�Ol�j1�(ج�v��9ɞ��&u�r�3q8��sכ�*�ó�j�=�nM{�;#�Q2�{O���x��%�Om[	�P�7��}r��+:�v:��N��@��Ž���'d'��k�{o�Y�t&��M��Z7,utŦ�OB��BBO��%+%D)O.!�k�#\gT<��6:n[��z�o�oe##m�JO+o�[B��[7V��<����V��w�5M�u���(�7/4��m��<F�jNP�j�qa��y��mR��5��Aw<�m�ӡc��E �lO�r��~���>"31��\�k�oV��3�s� ��\9ys��#d��)Cc�?�τ�y١Ϯ�8���k�/��,}��'�%�3i�[5=c\Z�����8�R5C����%-��+��͈�ҳXiO.���f�3\,�����Ob�͹��
c����w��ۙu�y	��������5N���M�m�p����
P��Gh{p�~��\[��[ᡀ5��o"�������è������q����']1�l���voU�u-�����{�
�˜嵺�V+�IԬp�55��\;g]\Ǥ���������{mb���W��_f��٧̼x�3P�	�,Q7�Փ�l����M�M �s�G�D���C���}��{���F�u�~;�7�OT㋽O�"��i_�-�q�N���Ao���ʻy�1�{g��|�:g[���5�q�:�ʳ��fQW?�����=������Z9˕{n���d��5y�i�*����:��T�MX�9�C_*������PvL�_����N%TY��{H;	����m:�ێ��L�J�=.�>j^���e�ͨ6��+Z�|���ld�%��w���j��e*N`������p�:�.8��a(���K�->�Uٶ�*�D�MD�to�z��5�NC�>�M���	\����+�%��6�[�{e\u�z`^׶H���ީ��RWW�;L��j����ކ�<���cQ.fx�3qU�@ݽ��-��6~Z���ʤ���*[4�<��[��p��fc
�w��o;����3�征aLB�zJ�&.]�+����kn*"#.��������{3����|q�7~ͳB�M�:_N���f��q�	v����J��k�	�{��"��W�E�ŋ�lp�}��5CS�����w5�2�.j��öq0������=���$�1�£u<��p���_d�ݩ�A��-$ÿ�q�
�S
CX8����	XxԻ�#(cmr^�\D�ɬŽ�|ک�NKO;�wOh��|���N:��)��1�t;;�(��-Jz�B3�ԭ��6*}�����E�����1jR�p�(?j���f���xH;f7v���Q���]	0h��E�F���:�L�'6��,��ڳR�@L�2��q�g�V�5�}�G�4ܱ������c�Fmg��\�T���R���e�v�{���q�����5=��vo_�e�JK�a�ټ�δʌ�
�+FS"�'<��qʹZ�yrq�d>���f�:F�9�ʂ�03�Sޗ��h�tsz9.�YX��'�����lgΟ��ke�E��֔��X]�B�z�ʫ�a&l�D	�}cM��G�!*]v��yB����W�y����}ϸۊCPuq 믥�TN�J�l�l=��/N�l�B��`�Sw9�����V�aڭd��R_Tm()j��5��� 9L��5�0�=Z���z�ԟ\�XS���|�JN㮊�CoŚ2˚�k�'.��I�ރݝ��9m�^7p,)����PGp5�m�t7,�pҢh�؂��{}3���/F�����گn��}��)�l���a�Yށa]���1�v�ķ#�"��N��f	�LE=~rR�ɪ��uuOA���Ǧ}��0
���j7�Wn$�2�^���z4�>(���|��󲱮���wr&$��<y@vT��y�/bu#T�#G�;V���@A'��9d�	��*�]�}P��2�P�k�O�T<g*S���*8O<�;��%T��}�#����Jח����O��/��hF"s5�S�,Åy�Rt���^���=@�CA���[s���>\��r�jlJ"^w5r.�[ju�� 7Ъ2�1�͎�ճ|�*��Q�83o�oP���b����.�}���&}	��p��F�U8ET/��_�)���u�!��yg�Ӛ��7�e�w ^϶��NW��Ì�˨=������~��zn:��q�c&��H�c������ۈ�ori�R�ֱָ��ǕJ�ܗ���h�F�ѫ���,���ͭ�+\v���|�!L�����Y�\T��j������ܒI:�e�{��|�÷��R��	Զw������	��50�D�s�H�Խ�N2(��\+��*�9���ޯq�����B�Dr�^��ZEL���PYO"���=�ݚ���y*�1��3h"�\I�h1S��vƚ�2��ā�"R�N���h)�h����nC,�����:��SY�Y�n9q.�P�M��%�R�"S�B�Z�S��6��uj�d��3���$gHxb��N^�w���6�U��g@���U}%���P��v��ݔ�^�F�ƫ�jb�x����R�z]��a��^
�R6��]����n$ڨ���zg>�m���5���Bi��U���v��m��Kn��@����}q]Aҥ�Q
S���k�5�uC�9��@���o�U�Q[عOl�P��%��%�9�o�W-}=��XX�p(�?�_*���H�Z��i�T�|�S�.������-wq\������WN�8)s�t�˜3�ym�B!Lt��	O��V�'wt:I��6U*u�y��z�ڄ��m�w�xð�&�1Ԏ�烮y'��\,W��}V�>�W���=�F�8�I�龩�I0Sq����$\G!�5oLQ�@����[��|p{�8����WMē�������Tc��'�]=�G*˭zU���9�������d�/�/o�kV���A*�8Ѫ��X�i<4g#b=�߯i2١��ˊ���&ޥ[�&��7\)��v{�B�ngFh�y����s؛Ok���-Ρ�Xr��9]�;�v>�PAV��ݺ���AR/�L��ddz�xt�{_�R�*yk��{W�n�������tL�`Em�G�'�d��2��
����ۇ�~��h���kg�ΝbO�3�9�ޥW[�r暓��<�4kX�ߊ�M�T	�:�=w3��;�e^��S��jg�/_&�z9�d����̨*��w��:ɖ�&��+-C9]X�M����	sb�Z}p��m<U��j���{��d�ut)Ȥ4]S�� �-��BW6z��*>�	e��9�_a��Ŭ��on�oZ/{�:�:Kp9\���e_��+��������S=�yD��tr���<�'����?-�
�"�ԭ�S���BUE�EV �3cj�p[_,��},)���Q_���{)u���
N��Y3�/0�-���J��ې��x��SH�?w��KF}�AA��O�Fw��Tn�V��(��yi��5�km#l��%6XT�����Y����f�n�[���m2C{�rE@�7^�
k�V9k;WT��lq�	5���}���I�wt�B��)F�t�쾚z������*��k:�W��Ms�
�o���=n�m�Ոk�M{gN���.i�q�]+VA��%�F둾\��9���f���i�	��wu�P��k�w�f�G4q��s�8�&�R�	͕�ty����R�/�|��0�.����u��I�WO�#�4�R��Pg �j�����9We2�W��we����B�8غ�2F���J:�(Vb�)�U3�ڈ ���,�g�|3�݆y�FY�ە���1n��
��t1>#o3V��n�b-�*�9�nQKn��IRx��ʚ9��$���n�,��YX�t�՚�*5D�-��Q�9�ݝ��Ӵ��34�OE=(jȭ�8ްF.��G��M�*r�}�o65P�o�f��H4�c�?��}���e��������q��T�=���<�x�ee�鮝�����Pq)�[\�a��0������,�v�kr����Tjm�f�(TLD�T;gC{t �6��ve�ki��$ٵ�W]����=���R�v�Eğ*VvAGz#���oJuL�۾�t�vs�>v�R$j�ekO�f�+E�q��t��@}�5�ts�
�����V�=�j-�\�S�¬Oi�w�s�[���L+�#�m^�D*��f��<X�G�V���'�O�'j��{o�����a�@��v�t8�}M��T.@�wLYR5��d�|�LP&�T�k�
��S����4�Ӳ�
��ͬ�B>�|{Q���7V�ݩ�N������-��݂9��a�����A����YJ�v�v�.}�(e��a����3��Qt��z���,WRg(�ۺʚ;_T���c����:���WaS�_.�%������:w��Z��:ջiz�S��͒4��ȹ�� ��R�ݨ��yUr�Z��0�'-ԋ�>d$��;��F��G�]�����k��>(۶U�v�;alMl�4�Q���:bBKh�>��>�Y܇qT�Kt
ü�����\����y�(5LV���̀�N�L�衤pf�eZ*���N��],��Jd�Q�
J�y�B��P����78��Î�(�w�7����,��EL���u<�kX@& ۬!V5-�1��5Ge��p������SF���f�9Nͥj]�WżT��paIg(/�X��@�ƍP�� ��*i5�]���S�����`��D5u��[��nhB�Æ��ff�)�.�������0V�0c�6 t�A�ƪ9��ۥ�����i������'OU=���S���#,E�QW���S\�rf�6s[u�� u737�R>B7��^	u�;����{�6o��V>������B�(T��)�)_dS*EiiiJJ �
B��D��S C$F� �)(�(R�)�h$2(
h"J��
(J�D�$H������
�(F���
H��)j���>����4`o�y�˘Y|�L���+v+a��N$�n���g89`2UjHN�<���m��L*l�|�'��Tt�rj���7gb��_�ow"�L流�
���uNi��.;�e<հŶ�[��_��s��0wo87�4�|��+�T���-kQ�|(�z/�ny�w����	���G��]1:��B�C}SI&��ys�*,ݽ����W0ӽ��n�!����l+�+s.y��,�筵2�:�Ȣ���Q3T�(f:C�9�p��~"���tc���߱s�_I̶�����U��^2w��V�'��s���s�z�E=�b����Nb{f,�yڅ��3۩ﳧ�랿�'���5����׻���c0?��׮Yc��v��3W�^Z��e�N�O==Ħu����ם�G73 �&��F��q��.v�շb��w�D���b����7�]s�\�����c��ʓ��ܩ�,=T�uAW0��dꄬl�c=���W��zSXˉ�-
*�:�V�Ĳ��CC]8��T�|�egÅKU��g��(�#��e ƈ�%l���Vw<lgC,��J�$=���U����$�'������O[X�c�X�ьC��|`t3�E1ܩ�-n�g�j�K���ac�+��X׍Z:���惡/�:���v��<����z��v��l�n���M;x�x�u3Ie�J��S���|r��d��Ӆ�{hS����}�?L�Z�o��zi���w��|�z��9m�^7/���4Eq{��7J
l+�kKC�x�;��/����K��:��9P꒱aC�]�Nt��59����m��/xC}\�����J�׹�}��3������MV%y8���zԽ!/��h0yl�Jח�*�o�M&"����gfK�.�z��.�T�"�P)P�J�5��ɨn{k�[��}4�]\��.�z�Cg!�7�+�R��?����&��M�Tzf���㑵}:�(U����U5�֓7���ׄr���n+r��t�J9��%쩧�ʯu�F��i:�NP�Aچ�^�c�B�32̋'݃��4��v�ޡ��p=�@.ןf7�q��w{εuL43Ҟ��{���i���u�y[b<� �� ���V��L��Ώ;y�(tDr����.�Gʢ����o۵8�r��u���_n���l�}�iR�KF�7&؋5�3��^�I�Y�y�t�{Z��]��y���W���p��ݲO#�<�{����[�p�O��}ip>n��Q�j�aa���U���(T `Ѯw=jkw�nm'�7��*��܆ep�d��D��]��������K���^����z�Q߫�z�t���6�A�o�-�ƭ���z��[�Z3q��\%�B�7��x��q�����SM\:�֭vv�G>�T��{�5V�d�{�^���=r���/�ʌl7������Я{l����v�.�;�X���㲼&sG����uQƫ��޾Z�i4�ʶ�����Z�9KH��|��z����lWPu
��)��5�vk��۞�k��f�v�(�]MX����T	h�ϯ��ח���j��k)y[�V�;��_vc�9n�X�(�G|�C
Z(-w|z-��j��������f�T�r��W��x.Z��<�壃�vRܙ�D���B��L
⽥x���ͳ���&%\V���*�c���yC!�������R�+Nq<���]�:�m�%N��:���uu���eP#�G֩sv��ʐ��.��E�4��]�5���o[�gpSoa�s�"ѣh����f4�]�ѽ��\s�ܗ���:��6��j!����;��B����;�qV:���`��jX��Κ�Y5�k��P�T�I�P��wdN�#�������_.:�OJ�(�����`�f\�{W��څՊ�u4�ÚM��v�ԕ�D��#1}A4�e8��D�wϬ��Jmg�ܜ�����xyKi�Q��=�_�cY(n����SsB�qn�e����]P�����|A7;�4�x�S�o��d�V��z.9>k��������i_i�.�8�� �Ct)����L�a�O݋��)�ldD�}p�p�/�S�J�q�>#6q-\���e����@��c�������q��\��.P�ڭ��V^?�xx/M��;8����믤����%|6z-!��,�m9�T����f�
iѫ��:�}�t�ȃ#���tA�U���Bu�F��n�,�L�a�w�;E��l�l�d3���k����S��H����ɹV��m�5�/�]���v��)_݅�����*���R�*�9����K���"���-
��{rN��������yT�ꝦU��R���������_O+�3X�*�',J��>}�o��
V��T�TIK�"���KW(�iX+Oy�q�[���/���=����{O8�'M�
a}�%A��.(<�*N�yp�==�X�[9˜*}5_u���>lg<f�ʕ�!O����2��s��SXV#��T�+�ܮ��{�Դ��sZ��7�m���S�������_n(��H��'9�Z�`sKx^�歗��x���Z��]�OjΪ��Ǵ>��A��V�|<��Y�f�ޯ�r��)&+�4�*H��1Wz�Z���#q0����_)d�!����պr"��ڽۇ���_�u��v��©5sa�a�rX���5\��a}E���4���D�q���_���7�l�>Ee�kAU}AMx�6^�wa{�t73go��4hu.'9�Ll:J���O����9����C���Jo�P���5w�~� �GƦ:N�q��ك�D}����7���'b`�|���q�j�H|�,�C�Ǵ([Øa�MDWd�b�����f��ouJ���`��ޭ���3���3�	5=�ڒ�έ��o,
�K�a�q:�q�hAG���m.Ẹ�Q�/I��x�4=���J�do0���ڠ��~��A��hifջ�����/M��>y̵}�:��9G@�>'1ODO�Pp�g��u8���sQ��uzF��r��bhW�r�z����7tP�L/"��Mi�N��φ����.W;`��鲒��x\�=Ќ�״�o�c)d��[S��R�3���H��΀n:dx5}�##�5�9��q�&�=�^{{e��1瞻C�t�|�Ԏ���O�f�ޒ���������3�~���t���3�|_b,����9����(J9�I�`L*�S��y�#M͸����?'����[���,���sQ5����=E����9_;��.o��,v9x>�SWv)��c^o�_v��C^�0{NEu-�Nv&�r�b�����5v��A]U\GX��62��k��+�6�QxE���:��@��}\89j��zw�ö!�����k��tp�s���%�e�VК(h�&
���/���n�,#�����~�u���߱-�3Fnɸؐ�$���O������U�r��U4�{��q^�{Uv�D��6m�Ӊ��-Q�A��Y��G̒������Z;��}X+vssk���s�{�a���V��9I���Κ�����yAG�nW&`����SX���s���g�����xM�>�%����(?:�im���Hϥ�z��E���^;SI�@YX�d���Qs�s�e��Κ5�nv����XC�`������/&�]�_3��뺝s�k�^I��<�a���wmT��ڛ%��c��fc�1;�(�*t����S���T婳�=y��^y���n�OEh̗����w��V���%�N�B�n��avW�e����]R_z��r�g�����p6�;�������ǯ�ۼ�ydc�P^��yU��*|�ף'	8|$x�Э$�4,m\͔4���:�N�q��7�h;�.� ���3��O�j�rնF>���W|��({�jc4����C�s.���,��W�Zn�X끒��x���׾Oo3��Y�t�h�C��};�ӱ������'b��> ���������AG�ڜ���hD���.��"�Y5�嬼�N�3�vG�>}~�>ÑU����?a�ާr]�':�;�J�!���s~��v51������e�l�9�������Я�hX(�v�GS��oήV��p����v���=�wI���WE8i$�ro$�\:�wRZ�e����g"NY#:��Em�N6r@�\�Y�p7q�0��~��{�����Չ^�O�Z��9+�7O1��N^D�XeAb��N��ή����
�Ep
��k���v����žn�dy�9�s�s�=�Dx�*�{�!N�Y�~��גF��6g�v~8�$Ԩ�u���
���g�W�[����^�P���^�f��q��M�����$��" a����Vf���c��z�o���V#f���r���ū�g/���a4�ʋ�u]�<�"#�h-AwNA�]Y��~h�N*]'�U���;K��Fo9�<��͆�n6�"T��$OD���MF4�y�K��9�,^����J�7ﴭ�_vlH��M����ղ_����$*.zf֩��p�'5F���vˎ�J���s3'�ٝ��pn�0���H��Ί<�oc�XU��W�I[��1�qm;��a�9 G��	���=��W����_�]�c!�]м~�霋퍤5�C�^۬j��B�;�qQ���&Nȏ!�B�B\ݚ���͗���N}P0���O��M�7�����S<���e���B:����0w���]yD��2�ɳ*��'nhey4�Yy�K���5����'Oa��%��+���[�a<s���c�Y�����lY�K���<��<��!���I��\~V�g�O�k�}A}��������̞;û�� �3.k��-�H�`��B�`[�����v��3>�y:�^�a�HYB��"�R�>����t�f���Cu�׶gQ���˶uޟ|j^��,���{A��ҧYd��3���o�ϰ��~Jⵣf��摽yE!,m��#���:	��S�:�a`r�k�ܵ���8�����W�s��s8�|��.��5�1��2�xA�ЉznyS�t�V1�Z��������t_�����{�.uտFs=>dW�nS4(�'$9�l�P��J�N`��ި���ɕ�r��
i4/r����n:�|�@{�=�c�re �e�$�a���j��q�[T5��z�w�hރ3�8����љlN.���'�[�<��J=ު�~	u@���&u�w3�zG�I����<�/��͚�g�OhM9u�x�3�w�ѳ�ܨ� �k��%���:���;�~}g��Wj��4���eׁ�Z.=�=5�f�����q���|l��KnB� ꩙����|��Η�΄�:��
��/�h_��v�j+#n!5~����f��VDdH�4���0O���5}��9�q*��Qj(�Dgi7mX��QWas�����`HSԞ���*]�})���� ��7�&��0�je�txUɄ�L��-�P*�&mSügN%��X_ƶP��������mT�K�N[>]��flX����
�v���}Y!N���$oX��"Wd�4$�ڝ���6L8|��A�./8T�s�l���9�|M�k�3}�C�\�JY=P��ϲ��_V�Ϩ��ݸ|}#��mn����w��ħ��(`ntԟsQs���ϊ��~�F�NP8��u��*�t:�D�����α��oWa�e]�s6v��CF�Ը��u1�_��N���8ީ��>��F�R�~%���uE����^�xM�Yl��V�~�R��'Y�{TW��W��5�x��g�i��t���ի\���Dς��΅'$��J�N�`^�\x'T��}u�+��v�~���VŠ�G�빼���_�#����4�wE����B|��=1`�`Tbv���v��Kb��+ד;;{]�uw��͗�t�q�Oi�[S����R�0���>�U#q\��Uʃ�Q��b�췽$����c�G�Ǟ}�<}�п�ڑ�<I�Q%x��E�5�RS�1��]����խRX����Ηg��,����x:u�%���]|�'�e���{G��Ք7D�l�*c�$́ɚ�dQ�Kyov���(�/3c`�Mc��k��2�yD H��y/���3��󝑀�-�1Vv�0g@H4c��!�n�"��	"ʚ��ڮ�ofZ2۾�'=�*��X�[��*�j���c�- V��n�N����I�,
Y�e�-9|�؝�.�+a��ގGD�Ϻ*l��s��K��L�ǵ�tY����d9�H{e��1ެ��u��8��ך~/u��Mhлi�l�M �e�����	�.��";&��Qo5�q�\Y��J���'H(���k��R��#wyK]�)��F;Zq������58(������2w+F�,��t[�H��T�̩t+��Z�q�"L�ݼ�uآ'�����&t��:p��o<pn�*��ɜUe�ҳ���c�*s��/��Q"�7�:(:��Npt*pͦ�"�_5o�5������w5t�� �����uٷ�6ݣLQ�\�4v��:u��ǕN���8BQy�-[-��bC\ g	��V�֞U����o��ru�U�>V(���p�ݺ$��K]K8h�;�l�Np�up�8�EgV��`�G��s5�G���v,�6R�s�dFI�)\+%_��|�R)-�z�7C��L��6�[jf��rwf���iRn���;������8�J�`���z&f�}��"�᧱���a�<q��-:ѨB�D�酤@bwWs\3��J"FĨL4���G}Z�JA��Y��v_�k�f��@��N��Y��U��U���^Q��#T�����δ��t�#ռ��c8�����>��.L<ߞK�-7�5��Յ���4F��xd�������aB���_>�Sy��(����3q�y1�w��*��(k��Z�X����k�ʡhn�\B"Ӻ]c��_bH*��}7y	�	�IT~�[ŕ�ߟ�����������v���}��7��I[W�u%Ū#=]�v;bT�m�4m�Ε˧��b���������7}�+}B���}� �k�R����:��
|{��K��q�]�*ck+��J�ޔ;�r�t�H�^Z���C+f�o 8��N���0=\Nl����qY�<��̲y�f��!!u{��{�dvX��W,�o$�vSm�V<���/���9��(��,pF���"4��zy�6o�p��޽�ã�O�����h#)d:�Kh�d���Q��i<���@u_f�~��uZ���<���D�2�认\2�
���r��W�e�{N�Ҡ�3.��Q�s����-�I�`+]0`�	g+���]�/�ʼ5�ȘK'nMڂ�뒊��*�J��-��7�ح P��"���6�t�\��*�
4�%�y��N�I��&*�&����F�kS�.�b�2ޜv �!/�K�4�ƛ}��c����u�[N�G~w��{,4��}�~��M*R�4#@�TE
��-D�M-4�HP@R��!TRPUS�ICMU%)@1-%@5CM5@UB4�	SJP��f!$KDJ�5T�SJR4�U- �4�T�K�R%4�+HU!T�IE�PDSE44�Q5A-,�S4��}xg��ܽ��Os5Vl;m�r�+!�`���[BpU���jO�0q�]�^Y<V�3�W��u	F1&e���)�Y�V�w;��~��q��J�C���s�]����[�x㽑ץͲ��A∷����P��G�}��G�� ���jL��O��:s�4���ǻ��i��E����
�}�M�7�9���+).u��1���Y��9��o����|����޴�W���^~��3j�x�Q~����^�KJB�}T�MqG���	-s�jOa��5�ϖ�{<���t�<���/U�����i�'�\q-��~t�[�2#��K����㴫���'����*��x�c�/7�Fwl�t6�`����_X:�
,�e��ǧ�i��S�ꛜ����c�'5�%�]�����u���5�\�F�����8�ǰ�$ljueK��]+�1�n]>�a�q+N��]~�/N�ʄ���1�_1-v�B���5x6.����&��˷�U����A���t%;7<��͖<��ۼ�ydc�P^�����C��]묝uV��u\TW�^��B�&�(ovG*N�.^��ܮ��oiĂ�~��3��Օ�gk�����sI���/�ބ��f��0�tRb?���6�]����A�ܯ�5��X�w��^ ��8B=�G�j�(�<9\j�WK.���Ꝓ�u�1���/X�8I�%���K	�C���-��:��ziS�Q��qO��ꝳ��\�����Ԇ�̋�,��a��>U�+&l��2v���=�Ҵ�O_�UWw��v�C�yF(-��ѷR-��>����|����_�᎒�7�[u��ڟ��iu43�v*�R\�O�&#��,����^]:�9��}~��h�Ub$�`�0�zq���̙/�q���Khd�˻�w��\���6���¼�<���D��/8��U�˿k2ϢԐUA���X��U!q�u(ڵV*�5�q����f�O{ctyܥJ}1������AU���%�g�*��D���[S�Z���v�t�z�S6��h�4R�8^9��p�=�?�W{m�>s������~�Y�8�����&����h�Yo�a���Uc�eFm�,d��G�+��/��a4�ʋs3�7�$yN���RF�rd<��
o�����Wx��Q��!�X�ؑ�������o��M���u��s>fh��#jZ5��r���-@gV�/z�Ez%6n/�
�5�fČ����Y�ū�>�� ��4��t�N,�m��_��t���L|mu-b9�LOQ�E��]�s�VE9���wnS�1
>����e�Y^إE�^3�*�b�n>�βrA�u2�5w}.$���w�~��Jv-�E[�&`���͜�������w_D�6�Dm��deЋN��e�ʟf�|�2�yP��+�q��kl���87\�t��I�䣼��+�(�8�ϭ��W\���rŇ�ՔQ3ǉ��Wл�H]�Wo���=C��C�����γ���Qxe�j�=��[�I���w�*(c�Pp�v�y�n�ܗ7f���/lfӌ��}	z;^�<�^-����N���3�o��W|�GN&�L`����Z�n`�9��������+F'ȼ�f�7�-�TM�G��vڿ�U/	�ޗ�[ꐲ��~��4�{�N���]�f��yu���;׊�kؗ.g|ew��\"v��f3Į/�1��r���o�7�:.��PuӐ���շ~8i�q������\���mtF��pp��\:�g}����yS��+����c�!�\hQd���+�L��ty���@�_��z�6�4���s�N�3�2�3���C���^W\au���[R���OW�a�ѕL]L�g�|%�<yb�i����^��Y��,��w��7�I����]�};�"��#�v~(p��BJ�:k�n�J~A�p�����r���6�nKا9&^{����̖%�k��C���[�e��D�2l��Y�*ѕ!���R{�0e��&��a�J�l�u��๹�������ҵ�y�uM|Û�M��o����λ-j�]�q�ek휸��đ�����S�
;q�m�����͟[�N܉cg���|����鑏��@�^� r�������<��tX���f���|i����y�{BZs�w��w���v�G��S\g����ż�6L�/���ݛ$���遝H��e�o� �z�1���|l��M6�+^[�d��'��ح���:���A	����w!�w���	��c=>V|{��7q���� ��F��������!N���}	u<D�d�5'���.�ٲaǳ��p��:ȱ���W���r��i�c����Ԡ����*;� �+�:��L�ub��F�s^��:5���s�q��MI�s����8�/Ê��c�Pt�v��>#M���&f�`9S�"�;�jS�3�0����U��w:�>���CF�����t;�}�9t�T���і��j�_仩����VW��+�q<r7���emȧ�0o1:�Xj�����,���c����;w��޺3��98N�p94����d߅��E[�4t�?86N3�ݻr�;����LX���R�3~ٽoaN�2�.]&�Gq�Yo3��+��ɣ&~ǯ�DR�p��S���1@��ku�, �-bu��*x�\�2��e��=�s�ѭ��������A5(	�n�ic���g˪��3~(dὈ+x;^�</4��,��n�����*���_��/OE��0���6���m�vBM�I��d���5xox�=���<�&�.�v�8^ܬ5Gĥfa�3���H�W:�xd��ҵ'�.Y�MVM��b��F���[W��Ly�޻C�t���x�ą�UC#�[�������-]��Q�;x��T;�F9v}�x�.��=^u��OU �8K��<	<��n�z�k*�}qj�T�3��]C��e�XŗR�÷V+��i��{�#�)����sl���wP�^�f�Hܚ�H�{A��p@�$zP5 ����O���B�z�hh������HһHS�u��$�b��+U��wЮ�X2O��-2� �H�%yNb2¸��[r��9��F<{�v�U/J����K�59�%c��.��W���" 5_B�BZ�$Г�]�L��Φ�&.1?�2�g�h�f:c��e�%���8���7A��S�$�ڂ����a|�%ɫ�ˡ��~U�N�>Tr��&|�i�h�m��~�."1�GO�9.��y+�){�c����\�n�`9���.�\��jiQa��vo��S5�C�>8oc�z11�+7��y�;w�ZEG��p;���q�-�&�Qkq	-��D�X��Hbj;�����Ey;)@�6wq��Cn&��a0�z2p�Л��Yu(rG�R�e����b�1t��V���J�B��r�������y���_����~f�e��fL,��iR}�g�m�X㉜^��v%m��o)�{2{���U�_0�/�D+��8l�P&hT�Q���O���3��E��v�W�S�q��	����@e�zo'����M�u]�U3Oy!�X�����C�?f�W��@��C+�o׍����.t[Lu��4Lݫ^�)�o&s���^F%��,oKֺ���8��6�ңթ�w@��2�S�<��J����ܬ8j���S[�r��[�/�ζ���oW�>��������s&N���xGwaݛN*��k˷U,՞���gN&!��8����,�����:��+��{<��rO��0ѝ�NvVK$��F�ЖCD��`e9�ʾ�sQތr�ӹ,�-�g:_Pz%�N���@�r�%�>��}���5�b0rAL	���T�B��Nq�o�~2#��^vdv��B��5!罝�WN4�Ά�5L���x�ㄝ��!;�ĀZmNE��>�o8P�ڽ󻌩^��Z�{���6�wJ�AL��gud��Z�p��;ǂb
C0MC����k��ʢ~b��Y��%�l��]/7�yő��eY��S篻vʬ�b�ޝ�`�w|��{'.�Y��G5��#a�N��,�ɻ�Yu�1�I򋢫��
5p�R�ù;+mr�K}�ܺ��߱�Y��aY�Ν(�l0#6J! {�	��v�w��H��+�rY�~�ӌv����&�����+��/��a5�*.�uU�<I�cLDv�-<��g%��2��mO���,^�} �^c5F�!C+��]����-�k&��n�"���3\�=�u-r4����`��͟O��#	wK��)Ḽ����3�e������ղX�Q�Ǉ�:�ʭ���t�b��C6�g�)�fb���47'������0ws��-��Ǝ�Y�,z��y��f?��X��h�gO�#�vP��EK[z3��^�y�LsUX���6n=Lz�;�/6�[������lk��E}��A�L��C��+�55~7:���R�����]Ǳ�Jǘ���m�N��r7��*������ɨ��J�U�&����هO���6�&��zt�O��9���˝�:f^﷥ƾVT��n��]K���86oQ��C�C���n���,W��f�Z���k�N�����9�9��ϟ��,^�F��cL���9Ԗ2�=f�;��]��w$[@�O��݌*O�ޖ0Q��M�����Uft.�hU���.�X*�w٪H�C��SD��8h�q�,q�u�Z�U�5��N!�Ř��ʮ]��N�����.�w8n�n�J�](.�\�-�Ҁ�dVծ�4�/�z~/1_��`a���x<��GE�t<�i`(�^����>���g���@�g�������Ws�7{����J\e��g�3�o�A���q��*��N-��[�Q3X�B�s���/�=��F-��f��Dd��3WG���jr����$;���W�`ɗ[�wc�qϪ�ݐ�7��G��~�=Ļ�%��g�*��8|���x��g�_�v=�����a�Z����	���e�/��$��N�T_9�`����[�W���i��ʮ�����+����m�CҞ �9u�x�3�u�l�*=�:��7��I����~�9]�@[�O��jd!z���FZ/���}Ig6�!�>��'ГV�Ě�˩k�_�;�g����"t�������Q�v8���dm�V����������T;n8��P�/��4���8�����
F���Hk�<D��%ɡ'���.�Ku�洙�� ����3����;�Y/�i�c�hx��e�_/(z?���[�SS�`��D��IJY5~ruυ�(�`uA�ټ��ҵc�N���V�wGa쫴�l����o�h=O���)6�gO�˽=��KNV���p=���ME(lf�{��5����q�ݍ�w��OJ(���{�Jy�"{b�N�� ���Or5Ҟ�&������?����;n��o��׹�C\��Yz8��PǷ �)�*�G�1�Z��);y��>y�&���kp�7����WC|;�V�<����+K�^[��$�e�%�N9[�5�8|z|������ۅt��7��ｕ��J�dxo1:�[ڠ����ω���C;	9oR��.?�F��q����?��:�NQ�f�~'s�����o�����E����K�X�����8_����1v�ͫ�*�Ҭ��ɻ�P�H�X�3�K�=���{v�]n߲�������)uX����R��K�����N�}{r�Т�ݢ�x�Y#�\ΟT���Q�ˌ<k��������TX5��P��Z�z�r:1�ޭ��*2�a'���gg��C��w�gr��W��!3��T;�1˳��]��z��^>����	w��e�w�M���X�PIO�!}��-���}R���]6*����r#�O���%�_{U���@`mEE�~����X���X8}�8 r�_��h7(+�~*=~�+��CC}�h�۴�nY`�{��"����$�tqP�zX�mu���M�u$�jz�h�oU��[�m�����kTv���ut`߄�.�`z|F�y��Ʀ'�^_>-S�jĵ*ICe���{%��L8V�����BN�{��C�<;N�D
�"��|1b�#�f�ʿW��w�����$���`��[�"���8�a'޴J3�ɓ.��s�a��2�/e��j��ck,��f��t&���F��"�9%Ga~��2&�U!�rEW�uUc��;�ߌdP�}]�:K�5qĶע0?:
G$�ڂ������^�>�jH����x-0�����Gj�]p��i���M_��y��/�C��*����:g�� �P�;��T �V���R����ӂ�δT��ln.�Cu���UI��˙(��ss��Ȼ	*���p�g\p�>����s'LY���c�����i�u�����WC����_1-|��AE,دEO����p%{��l�G�p���Xڸ���P���r�t>u^��K��)e
��Ág�����Lk]a��,��������^4,�7tP��b}/.X�HV�x���xo��;��3� =���ϝW�A�������_w��ڹ����wE�����т��X"��;#n�������N�]���1K\�h�C��};��lU�r�&N���Mʙu㙇7nϫ���1�׍�Rw���mK�R����EM��%�N��X쭤G���&�le�']�r�����fe�b�)�p��k{�	�F$����c7=cc�w�=}Z2�;����}���y��p!`��a���6*NP�6�n�ϝ '6ڑ.#+�^�;�6�ms�4y�0P��FG�WL:=��C�,n";0u.�K,�E�H�9i�5`�5�����[�-��F9�|*1�ƅӅv\H���G;^f�w��M�P5��q۲�>9�o�h`��7ušQ(�)a�,SLD<{�Rbpz�g:tBN�S9�\�VZ'Y��)�Jg�np���LL��b����3��̈:��
�ёs��1y��.,�z��#so8��� v�Ro���|C��^�p�y���,Vp�hLJ�y�r��J���s'�=Ĝ�]3����������#l�Z�):N�k@%(n'u�� ��]�ORA0rf�7@��ڃmH*�6,�eS0&y���m{����BF��I[�$������l_H,n����ֆ1�_3��Q���,h;Z��BJG���@���@��Z2uFr[�2�+I��M锒�RuC�P�BYz{��C\]ʓX�ۮ1���^]v-sP>���]��q�|��U��{��N�)]�q���q
�+6�R�<�N)Pj�ډ�qQ��K;�^�|��6�PZ�D�q�9ծ=++��
ɀ�wnů�V-�*tt�3�镳�PY����n��jf�G1�˼�[���]���\�٥#y�͏7�u*eXH:��'^�V��Y�;��d���'�t�w1��q����QWz�%�0�v���0�u)b�.�Xq�t��sR�4�03ǫ�[���W	��^���1^*/�4)�1%�+��5�]W�t�Ёwgn�R{1�+�pv��].Ʉ�"��ڸiA`�9�Un��s�X��éء�,�ww;�S����/��@-��u�+S:Ү;H:k�Μ/^(�&.�����$�F�'84��@f��L��M�r��������s �t����ޖڬ�*�oM��-��� r�t�3�	����I�Rܤy�v�=s�M�:y�4����R̥/���u؇jj=%�ڬ�UǑ+Z^�h�r�fp���WRޮ��q���w�(ű�_[C��c�W���������^!�-�h`�:�ɲ�5f�����wu�l8��C�q-�������Q]�ǃ�ؼ��Ϛn��,c-���n�]G��N3�A�F
�ɬV曌9NZ�m�,y]=M<����s�h1 �o����N㝽;uk�b�+������0D��މ�����uw]V�#3�SRΙt�=�;��"�9M�5n���ɻW��+M��n�[�Ƶ���=�t㗘����B��^�!�v�Ǧ��9��3�WR��@�Nh�������򤠈i���� "����	(
h����*����h���J���b*��B��i*�	"!�H��bJ" ���(j����i���"�b�)"�b&�"*(�������"
� �)�f"*a����$�����f��$��&"���"j" �&*��������b)�f*&�3*(��b���H"�jj��L$����H��j**��H����i����b��(*b���
j*H�������`��
�����j)"��*�*�)�������**�h�d�d("��P*��d7hK�����y�VI�;�����5���s-PZ�(��LN�Or����\���pI��p��t˙A��g/���ɵ�����ŢLGT[�M �k/,S�������ϼ�t4s�K��:�d���}�RpO�&�N:D%�����
]0�Wc��Ӄ����6����Z�P΍��;����S��Ze��A�X �$�C~��9ǎ�S�W���=���qв誾�q�Q�k�g(7�x�2�If��$�X
D���mNDZ���;61�$�����C�L(��
�W�����ƣ�5��+<��z#ȳ�3`���\H�~QT�[��x���d����d�9{�r�zr�9��iەN��-�#���Z�����'�w<��~��`Ԯ�������א����旰�m���M�Ȋs>fg�����[�|�NO���3��#Τ��*H+҅I|pe��xvlH���h�i�,��l�/���7��4_�T�Ik�=kI
�,T
Cxj��˖31_K[fhnOa��\�m�̐]���jE�E��:��;Z�/�p��GH���D�i�r@�!�_B~1R�ތ��^�y�Lr���U��-�l��c=bkl�ݬ*�������BX�{�/n,���������ʹ��ջSwr�*"�(���|pBI�=�/*���9�uv����]�̭�`a�K�M9ʇ5��[v�������S��:]��k^k�͕{y��np���.��̌�{:L.�b]�x)��_﫧��#��T9����늊�r����ُ!�oƷ���8�O~�oۧ
��o�~��k��tdP��WN5�����)��C��{f�B��q��ڀp?o#���ڷӳosO��?����2��gۉ�Yu���3/	�N1�{(+b��#��4�k��fJh��&ݿA�$���b��X'Y:h�p�m���u�M�-[;Ϥ^n��t�y-z��^c�/�5�(���X��3�]O���yO��u�y��.�1�'
��B�+������M6�U��N���[S��ωJ̱�2�|��u��4<��b�q���f�y��,;�lt����:���ʴ��\f0���C���z(J[���|��ٯv��Ŀ'��Bo�,�X����X�f�I���:�x|�ӱ�8I�(p�Q�0�Oe,mB��H��Y����lS���z��4:�(M��g�>E��|�L<4쨺�?A�=B�\�j�[h��/�~ퟫ? �Ԏ��f�`�-��ߕ�_�֑d�ҽ�:U�}r5��bW?	�[�]�PÝݜlÂhᴦ��+�����y͈W��*�����;�`�2�r����g3*����yHH�s
��M?~�+�n�Ǚ:O&m�`gn���3��[[]�@�qt��Bi��Z�b���E>�k�;n��sR@u4S�[1�r��(�
?������`�1�O� ���0�=;��FR=�*Wp�{�90�3Nn��X}���UL�q'���a��#$�)�t�w!�o�����$��Ĝ���u�yZn����dxD����J�p5؅� �'&Ğ�Sq"��؛�8�律^������Wj(wt�_����hz"y���W� ��4�}���f��S�Ż�z�˓�n}r6��t�S'}�b�ΜF︩�P�t�������;��=.�s�>^�y�mGa`^�Z�����/M���k�WC}�s��|�CE�WD��/a�̡�׷H��J�kW3���k㒂�:Eexm������~7֮=�:������[}ϽF=v�OP����:�����as���i�W�����	8�"-\u	���J�����`^�\xUD��g<7���(۾ò����q��9���:�"��M�,�ۃ0��.�kH� yml�~�S�>�5BU��3=��Z�-�~po�R��K���ݭ���Xk�E����<5z��^�P&tm���-��Hd�Ҍ8�ׇ���Hs�w��P�?�xdk�\/R�[�:���*�[ [^�s}��Mo0�+����=M���!�W��d�/}������sĳ:��+��@q���f��R�s1ĲA�����}�t��'�F'���.��Iq)u��J��tgr@}�U�7޲=�{Ӯ�Ly�޻C�g���k&Gt\�'�~>^���?<�Ц��3e~^p~��k��)񬥢����xF9v^�� �59�u�^Z�&�p;^�,�*.+*�Ȼ�%���ވ�`G�Ò[���Y�u�Q9�.νE���7��S �M�՞��]ޡ�[>��Uk/ ��UX��������z�HW�Ԇ	�y'<44�`}�z���i�c��V�g���d�j9T�}$Y+�q,��4��U��Tr|�ʽ�����_�_9�&��AY��	��3�vȅ�VW�߶h�	�s�i5�Z�g�\J~��Y>�8�ơ��|�������D��=:4ۛ����<�KD�>��]PD�S�������n��ao�$�[75�CY�����zO��p�5�̰g��PW�W
�.�i]g����<fsM��萷&�hJ�nN��87]�m�̚㬔X��#�w��b�8��kI�~�k�sƬ���uO���j��77�N+1u��t;ù�i��qHh�Q�?M�I�ua׹e@��F��}�;ޠjWu���h�GT�\���嵊\�7�B�u����`y�v�/{�s<��o@.�l�����3�]�N����w�g'�,���irTAx%��_|��5��6�۝��FP�r�4J��{\�m�NJ�ο<���B����avW�,��C������N����'</'��l�wI�Lʑ13U���Y�N��}�Mdd>��{�V'�7�����Z�����a�(�i�Q�^��z�v��2V],��,�����+S��z�n��/cάr9��B��ʑ���د�߬��������%ܟgy�brgJ]���"v����u�o��E�^��N����m�qgF���6�\��m�e�{�����V@DX����x��||&#��,���^]:�xK����e_Y2.�Z�{_f�k��>Ga�X�9?%����Rz����cS-���K.��`�D��^�Oѽ��m"��/\5�V�l�2�q ��e� �.�Rw^�9X�&}��Y׫N��ǲ9ty�s�}A�r�C߀�,�<IUX �H-�K2&<<.�5EI]1����[�v�&�<�����8c������ϹӠ�͎0#6AA��L�P��s���}�9�>'8�1Oc��^�cÕ�ӗ�v0�ܨ�3LS$��/uEe����Y�V�m�b�Jn���W�He���FK�p�^��x�Zy�*�[� �]~�6�D��=Z4ST�#��Ee-��v<�wk���n����2J��Q�`۸"�0����l���_�ڝ�.κ��عʳq+��=k�:�/e���)���^d�/��~�<�K#��������a����4���5ՠ���������`���6z��k�:��#��Lx&�bQ�>�dg�6$ewm4h6���w^NW:u�h'U�ýx�	�#���Y1;K�*!��g�+�31_K[fwY��&}2Rx �U��	7�&����\����E��[��$btQ3����ǐ�	��]�W���Iw�[�J��/f�N�>�oU\8��U1�j\�D+z�qQX�T����;�0�.=yp�d�����ԛe�l��R�������Uӏs/��s�w58��&�j����&󦹏�	��{�T��4�����[�w��o�S�'N.��}��ǇL��|7�ƾW�ꐲ�߲#S�����H��u:�{r\��ˠٺ	g���	�͘�d��|�D�������,�����k��#�c��˪X����ש�s�_���X��p�K�_�-�~��ѿX���F��9VV
��]����;�g���8���X�\wc��1z����gĥpe��x�qS>G��e�C��ˇUb��bz[M:�v9	�+Z���)~��cJ���fs5�ych�2�Ui->�}J	k�����-W��>P����_q����l�W��Zܻ�S&�O{^�P%Fu�U�B���&k1�V�t^�k��r��0]�wV����ݙW'i^��'�Cs�z�"�W�����W��;<zoH��nW�����C���x^����V�b�ݾ]������]p�g�=����ǞBl߃�0��C��ޝ���,�Ĕ&��0fj%�V{��9��������<zz�N����"�g�I��ޥ�Ω�ΠO�c�o�u*������;���&�x��j�����:��>���['��$]��=���E�{.�v�z�/�7��٫S ��(#���=!��l�b2Ѹ|����q�$٭��[R��c���zYk,�΂���S3�26Q���`ƽS�3�S�U�/d���7�afSˎ���f9�:��e�x���3#�'��)W#����1vK�/�����)Rγ��<��ɯg��[N���w!�,���Ƈ�$~�O���S4�헏z/��5,��z%�-9E3��#��?K�>o����9�j�:q_AQX�*kK�c�\)��y䛺�˥�6�͝�};�c���#�K�y׷#��a�sѠ�������j�Cx˞��9�e�k��T�� S!��Վ�(^-�x��57\�o*+��
�{�6�JyA�픵�0ւ���G_V�"�����`��Fn#\oz)�gsgie���gr�o�L��jYǋr�5gi���$��b�Qܧs%�6k��6��U�0�R+F涖�������(jO������Y^q
��<sz_���{A��ҥ�7�#�+�j�d��/X�����̅�}g�5�x��K6��N?LZ�wS�t\U��ϗS��E�Nwo�\�o�پJ���ٜ~plS���5�����`�����y���֬�~R�u���L�vi�4)j>��=��Rׯ����&�.� �N�^ܬ4(�R�0��:�\U��ti��s��ފ�V��X�Gv�LÎ��n�W�����C��<D��-��C��>��Q�����;�s�d�kL�r}%v�I�\k�Ϊ��.��Y~�P���K�UqaӃ�(�1������9��䆲	9S>�yS-φ,��]9�\�{K�YZs�>�����u�$zQ��o��<��{�z�vA�o���Y��@�.���-�o�y�Nv$UE�H��s�������Χ�񨳵�A]|꫈�@�,�( r� z~��. ��9����z�i�̾�h���/z�C#��ldzo)�X�;����e̹qG���\Lg�͗G�z�K���Q�|mu�s%h�n �c�̝�od���nڳ���\�ð�f�F�Y�r�z˵�.��MLy\W'�J��iKn�<���8�vr��|�b�j[�u;��g�!���3�3s�:��$��$���gLyWО�m���E7�&�n�N:��Q��J���+��(����z�ǚ|�����=�Nt��j㉯�sq�#�im?9b �R/�`ן�cѾ�ͯ:��g����ɩ.<�C{�FW��Mm��x=^ w��� ��&@8dxZ��Mz����l����t��S�T����=��ݳ,׹s%�жϽ��X�<4U.QK6��ƨeÕ�%eN��:ǥ_��;5�����M��,ן�o	v��2j<)m�γ���	h�v�B����40�+ƾ����;E��E���\O:�Ϙ���GWFlt��ݏbs�)�c�^����[Q���º긨��,u�hew����zBV��Y*=b�F[r�:|k���|������1�z�n��/|��#��.6�e��L�'W����y���=I���.>-Tz�*��L����[�;�^��I�u"ޯ};�Ӱ�e�钾�!Ʊ�Ù��9�@A��/����p�V����U1�&�)L칄�n_f�8�i�b�*y������c����8�z����"Lip�D��[/�/+�Luo���W��q�vm�&?^`�=�����[3h��vlZs7���2����1��Ol����㱃zӭR�6V��wP�2,6����	��S��jmӫ\�,�%��_v�۪��.t���Jdr�V�ٺ\k6Fb݆����� �(ؗ�q���
��H��8V����y��W�ǖZ���}$�WD/��=%l�Pʩsʟ��dۥ���M]���΅{����C������\C��au�1�Yߙ�J�2��R$(�V���V{���%��JgzC��6g�T���쉎\����ӌ=�gi��+49Ӡ�͎0#6 o�)�S1OMпm��}�:�`��&�'��zw��	���8�=7�s��&��QtꫢJ���RW��}%&0�Gr�b�s�ja~��#��fČ��]��/al�y7Q1�0F�y�ګ�Y_�O��:��W�'�I?��A�"e��*K�7����P�행�:��;���5�Fϟ��,������2EB�s�	�퀫}.{ƅץi�]O��@	}��Ee�����ǣ3�[��"���F�i���2<'�Pd���}	��koG_o���[��K��f�Q���7j�x�U1C��T4�k�����PdZd���2�^){�����yڟ��V����[���q�C�WN<5̼>���2�;���^�sɡ}��ͯ����g����{���][��m��|of�g~�7�P���w7���"��gP��7PJ�Fo�=�gmN������L���LDs^�4�R��n�1��t)ě��]�:RNm�=��M�¯_^�*k��>8��m��΃�N e�W���p��G7XSEX�8���W
rmB����Ö\��jT�����$4b�s�g8�2�|ۭ�״�]���㻀�9��,��)4��*�H$�B)�*�A�]�R�WAγ��%��-y�R;�&�2��x�mSZ�Ы���5���;�M�:��B�{j���6ˈj5�5��ER�͕�7�f	i����r��E��Y��K�C{�7*.N�gBS��o�\h`�OZ�5qi�E�q�[ڝ)�G98�մà�����_��(Uٮ�F�m�����t,G\�//�6��W+^����wD��u]�J��v�]uus��
�s�[x��%���ל���C���X�
�''���t]�)s4N�W��,��P�7t�
�t!u��\y�i�z��8�;f�.!�pU�q�B�9Y�zSnIV(�G���"J5:�:�J#�v2/ �c�V�bl�Z��Ĵ�\�ݱ`�𳖧fcC��`᪰I�>��m�"ܻ$��_/��M��6iX��4�
�ս�r��գ`R�F�K�*�+��g\[�6㋁�L�v�GNWP,����b����2�K��9u��wg]>��#�s8��t%�k�uU�66��MĨ���-��ږ�H(��N��d��6FS��}�%f�S������S�]oEA��}�h�J]�x�P����a������r�nn�VМb��`�ra�Vκ�P�m�[ǨKYn���Դ�š�C�������u'�R�	�c�D�ѳ�RK�Րj�q��	f������������\ �}0>�Dُ��9r�fV����/��T��JU�xt�9�[���H����he�j�`M����:���>0N�/r�9��֡����[y�BJn��{�J��%W �7tą_�n����Xo�J�o�8M ��3}g�k5�zX���>V�d j�ݑEc��� 2%�K��&��-�f��X���e&��xY�f���S嘎�ó�\�F�7u�14�w�w��t�.�#�=Ҡ�O:�˗�7 ��\��0��"Wjs'�Q	f�V˃s���cQ�}R�ۓ��UU�h|�cQJ�Q�����N�AJv�`AΚ���w|,��Jn+�X���'kkj	"��q������pF��]������d5g7��l�u!����ڻU����b�%v3%q���C��^0�t)�*�ƪ��}��l`�X����M�9^���B.m������A���&G���r}Au��QG��$eZ]�%�!ْ��y�\�d��N���:��l�n�6�0ֈ��X��k��	� �U@D��E5%Q4DMPU��QD�D0EAAQ-%T�EATDD4�SUUQDDD�A5U%DURSSPĴ�FI�PQTT�PD4UEU4�QRP�12E$AECIQT�1D�TTSD�L�D�TIK5CNa�SEPTLQ4DPAED�U%HQC@DU1TQQDDLDU0Q���4�Me�LEPUA1M4D�Q4�PMP��D4RQRM��ATEAPTT!AAD�LQ�ACEC4�D5U@SKLQ4�eM@Q�D5EJQTąDRQATQTD��ID��^�������Y��wt����[4\J�;���\�Q�]����L�|%vB���4�B�]�uҘ���{]���V$��-�Q�ڷ$���>4n�:�K����cqs42�iǺf^��c���!d1]�R�:�#�3ȃO9����+���僧o�/�WB}3��N���6��g��Y;c�vd�='�n{٬O����PޟWy��������T���	h�V�G@�#�x��J��Mg!^Ʒ�ٚ�E�j,wI���\wd?^��jxݟ��X�x�Tϑ�Fޮ�Bj�궳}h�Q�4�������x_�9�w�K�����Fvܮ5G	9 ����B�RF<����b׈��X�L�7W\�Oýި��\y�&����L<�9�qȉyH<�Id���Z��%"�}�=�-�N���_���ggfAgWe	������ȾY�a�{*/�s�{�Q��[uJ�z{�A@�s�@��O��E}t�c���ﺞК˭��J��=�9�{{&�;^^y#��Y^�w#]M3Z�Af�AQ z�7\��P̄e�o� ���!q�w7�2z7�J��̏l�Yd�n��uT���2�!��D�����9�g7}����͉�Ϻ���Z�igS����Xc�LC�e	��-';nX碥,ݬGe��b;uS�}kĵ]c�I
b�Tv"'pRg0�;�������Qք�|���Z=��vVN�kzR��+z�J����Vɖ��|-kÏ�)r���॰l�{�Vp�ʺ޾C�7du���2=>TY�ū�{�����Axi\�T$5��A��R�~-���lv,�RX����-�M;#��UH��x�d@���C7|��"F�'&{���7r�<�1�Y~�)�ݕϧ>���;���C}5&��9�j�:q_AQY�n��7}\�)��}�j�,bd���<1f��	�56��{��P�\���L���w�=T�d�Y����d���Y]�c�=QZz�����?'_�q��\]��'�3C�[A�O:��6Gm�1��6������ِ�G��x\OF��j��~��q��I������ۇ|���n�Uׂ^�f�þ@{�~�1�/d3��Cuc�#��1m�N�9�fT	�,%䙞q^��{��+}z|k(,����^��ׯ��R��	s��[����VtQd��u���P����>�:k}��VHu.e��و������[ta����9�}��o��VǺ�ݒ+Kr+,��-�����Q|d���$����\k���xF9v|"˿�9��"�_�E���a{�^^m�-���a"`D�E���5�+��ޱ��*����dUyd�4��'j�*�ne�z�Rڨxh=�|�͇��7H�eGɼ7�Z\\�p^=�q}���-¡8�cF���r�������5P�ys�m�|���3U{+g���U�� �.��OTJ�du})w!C쩕���٨�����ݞ�����-�3j�^��8kŎ�x��P�zs����UX�(�������B}"����.\���Ȗ6]t\{{v���;A۠��U3If��Td@o���|/ک��\fn�؋���q�=p�ւ�;q�c��N�f�S�5�3�5Ps�*���[
g7��<�.�&=�J����2P��ȯ��WG�s��CWM��E�Azs=xg�4Ҫ����:��T<4Fb�>Oa���(k5��#(om4[k`���F>ۑv�o�ܬ3��_�uX9�3��ϼl��R��T��ut�7�^ۏd{��Zk9C<��L��`���%�����f=X��gP�~>]@C^�C�[f⾛��)��i�z�Z�/9�,��˝�1�����p���uthavW�C'r<�m 6�;��i�Ɨ�-��E	��"��{ۉ�4���P˪�8�����ݎcZ��0��ދ�*p�F�N홄�� Z����R���J+���y���s�`�w��:�� �ϰ�\�HC�ߺ������+{'AO�WKt�7ê�冓cu�x�Z�L�FXOq��gLW�[k�SL�G�\C!}[�L�1'���v�b��fj���oZ�2��Uu-Z��d��"\�9����eƎ�up}�/Z��b����v.i(����_3�B]������e~C~��GT�f�J\�������:�6�|�"� �EO����a-��km�Y���������u�K�g�FԹ�9%��#O�(�K%#̽�F��4�]`�O�g%�Uߡ��O�7��b�T��I�P�@���|�/�B\�>��#�K1��W�{��s������<�p��A�#̭2����x��X��T�����x�׻i���Y��z���=V*�s�C��g�3����.��=�$�L�%TA���FK����u����=�Z�>�u�w�������+�NQ����~�Y�ϒ���0��*�y��+0Dz֓�y�����4c�~�,C�y��C�����ixn�e�ؕ��^w���%�G���"7T�C��|}��4n!Q���>'4�}���'"���>�;z�ǒ�p>�mހ�m��H��(��8� ��ģ�}��s5ٱ#$h����d;���3ч����e�ʓ��� �;�35���2�ʽRÑm���T�ut:L1������e��{�KJ�,�A}`���U�[��Qݮ�`�4.��+�q��¶��2�ڼ|�0̒� ���RE�;u.�ʮ���:B�w[��\�Ksb��/ܛ'�3�K�>��S���sӦf����>+NbU�J��F�b�^�S�/^�$�G��U�߬��b-�]O��'$G�쯄'���,4˓��Z}L�j�`��NV���q��Up��Ϊb���4�sN!ek𘑏Ҡ�d��L��Ü�*�����u�����4'Wa{cv�dW�ʺq�'g��qL;���\�L��F��{���{F6z�J��{� �1��GP�za�|v�3�u���t̼'y8Ǫ���Ȫؽ\�uf��guVy�ݾ��6�������o���A��w�eW�R�J8v\
[�q�J.�y�>���l�S��^��t�'����E���@Y�%qCZ6n�Xʁ3�]O��N�����O%�X{�I�P��U�g�b<���8�A�î�+"���~�f�jڞ7gĥfXʈ+E+��#��ŏ:y��N�M��s�q��0��-Ӄ�d9q~�<��K���=7�Wm��_Q�N;����V��.�eC�F��$�3�]t������w�{y	�~$����=Kc���Oyf�49�zI5k�'ӵ��]�U����)T�y6V��2��G|����P&�f���WgV���:�0J\�<��bh����싷�Ae�D��2�0�"�«xNWjl�]%sk:�%6v���7x�»��B�3GT�r�@8��*��riN=������8D=C�I]�|+j�f��(M��e�/��$������7�����ӓ��+�%�9 r�����@����U��|���=^������M$���XG5���4ݗ��6w�ʏg������,҂8����n��@�;}ٙ���T���h��y.����k,�m�WN�����#�F�1�Q�a#�T�*۝0��;�W/i[�xVáٴc+{i�G�Oh��W�����WHR4�G*�\:NC��o�~G'ם��J�Tn���Z�c�Ӳ<-�]ȸm׉�O��c7}�p���yf0-8ڗ��=�Z_�AQVh��H2nϤ�75���a�~��,s����t�0�X��Ǟ�'�r�yb��v܃NQ*q�;8׫t�l�>GR���:��c~���ո����3Z���6O�]1]��=Q_iv��bptǋ���:��\] ���x���߽�t��쥷�ݞӵ^�T�����u��V�~��L��ϗ���?�������~�%���! ����ȍ^����P��:VJ���6���ϯ&�P��OEH`^��G�=h�Gh ��zkG.=��9�J=(�aѽ�q�}X�o:%�r%�^��dc}m�X}D=]�E���'z�>y�rQ7�hRh��}(�o�(g��S{���o��U�G�C�^�g�n�wg;�b��M�"�ݸ3&1���[��ݖ�v�Tޚfp�ר(�`v'h:�ӃΥ�ޗ;��������a���{���Ϋ�;Z���	����F]B�%��8�#��2fw�ۣ-me�N��Ͻv��ίf������eyw.���ʎ��a'�u�l��$����\hvuP��.Ϟ"˼��m�����w ��e��7-�J}
�L,��Z 'μ�$��^��ȟyV�mq�ɇc�!Wɵ4�Y�~��1�l�z�/��x㽑�y�b����f�+�j@�>nP���;;����~5b�J#�o6{f��:��M9u�q��u�o�;C��7A�Wޏ#�~�b3g��y3��MT/���\���=�9ޜ�F|����/���d���;��v�+4�	�(������_�GW���8��K�BJ���m�4t'�lg�ԉ�N�M�ޭ �-�"�w'׉�����ċ�k�8O�c
��L���'���ٔ5����FV��F�s�[���s&6����~S8tU�^̶���.�<�+kibs�����waܥ�ۿ�������S�N/��cv�+k5w���i�ZY;L؝zv�}o���:jg�{�+YZ�M���^-N̸���,�pS������q��V͡;��tZ���;�`��ҚidW�.f4�x.ɸ���ܝ��w�1�\�x\��\�>���ǒ_���(�j"��V'i�8��FT5�늕�E־��Y�p��3�*�%��}��U�~��#��KE��
�<=�l��<�0�l�~�o�w�T/fK-�ݙ��܍C�s���ys50k���cZ�x�׺�*(mzW�:N�$#.}���햩�ᤳ�}[0�����4�A�]l_^�_�|�zD7^^��uc����Ð�����$�-+P����x��cl����Zn�_�^s���&1k�m(y�u���Y�����߰{�)ѪvOQd��/|VH��L鬥���v��漼�\tq�̳��ׇ��s=��� �3��yj0]�I�.�PJ_�/ܪ���K����g���j�ݎOz��s��m^�~�Ⲽ�<��E��Y�$�,	Ȱ�yơ^��+r}
�Z�-=Na�ڜMm519���G��s�~���9�u���a� d�j�J�@ư��^f`����?dɏxG{b�%�i��i� e�q�!(2���u�1ՙ����Pܣ�uP@����Y-ZǏp���qr���P|F�y�}�,���{�o�]@�b�)jͫ�A�5F(�:�y�jGj:(;}�v9WR����\����J��b�����~�<�@e�OZ�����-���ϼ����d���aY��Ӡ�7�n��z�)�w�r�E�0"���a1�W26�����d|�k����Hq9�zQ�� r�~X�E`��Tv{g%����b�'Ҁ��@?y��n|}��4n!Q��~���^ҧ0
�"�W��1zy����/&���uq�|���蝔{U|qAs��G��=`a\�n�TumP�0X8��;�{\1�s��|�zK>�d���G����k
CX�Q��?���$�,�q{��oR���Oc�����{f�P����H��tQ����q���D�i�rc�v#LI���=����z��ǥ�^����5{���	]�c>m�LW���T9��]�Ҡ골M���v��Sx�+��8��&،C�_B�#�K����/4nӌ�d�\f����_9�U|�GN&�h���VO����{{���R1�'7�py�;����#f��:s���o��W���O���'ߢ�7�!='Ww�z�~�;Y?5/��g}�����ʮ"J�(��e�ﾙmx��Gߏ0���J*[r�.�m�r�ֺ��F�	�bF&Q� �-fӭi;y������8�����q�Y{���I���)�3\<T\�X9�Z��zt؎8��*}����㘈�(�k����jR�*V�V��ꗳ'�]���X<�Y��9��j�9^��Mp~;�y[;Ϥ^c�a�5�+Z6n�]�	dl�I�(Se�DMa&g�_����VHE��BṴs�t�YM\wd?_3����ݢ�=}�f�B�rL�e�vu�^Hؒo����y:hy��_��������;�s��9{H��\fU-t�)�x���A�X�і�/�i�Uˊ��J�NuuL�����7��L<�=ʭ�ҰKx�z�d�������y2�zAA�E쎡%te	ΠY��<�}���'�{Ҁ�T6d��c٘���w�\|תF���~�d�@���
�R=}���~Wʱ����u��M�k��έ����^����F����(��٫s �J�dCs��~(Y��o��Fh�4�z�����&���ޤ}���G�����Yd�n����S3�3��5p:��[����&v��;3�:��O�\О<� P^����M_����<}���̏���B�+�$|��!u��e�zєҝ��3��"��v�A��k�C�\��.�!%,�����b���"�����Р����"+� �����U DW��_�@�� ���PE�@�_�\PE{_���5 DW�"��@�_���PE��d�MdC�5�	�3~�Ad����v@������`>��(U@*�P @�^� �( �j�C42��	UU���-����D��=��*�h���
�R�*�$��ʢ��{qU{8 ;�͑��T�E�����Ыf����:
S���tٴY�Jۀ6  �  6g��@كkjJ�-j�UY� �T͠�ch�m���)#c4�R�5i�J��������0����w� -�s;�s!�lk�]YEP�*S���Z
�30Wk����vmgC�Z%EUu��SM�:wC��T��F�� m�f�:h�nh�lK�e�[%i@��m$�EIP�� ۠rk�� ژ*���6�`j�i-�R����%"�v�h�M���l�@Lj%��� ;6�
֨�hM�ֲALEEi�	���Kb���KY���iY�����(�   "�J�P40�20� �&hE? �)J*� a@ *H� "a6�Bm$��16�M43A�O�D�U�       昙2h�`��` ���M$!�J�&�FOP� i� Mu��˫���͞yu�>�X�x��В �.|/s�:_�%�e	 !���#/ҟZ�$0�Yp�������_���#\?�6��R�����I$��(k#]�H�Q��$�*�ʂ3�r�ϕ��"��}�;{�:�I$�1�&�-/��_�t-(��El�d��ޠ�r��7�B�	�k����������htS��1-�W��֛k2!Q�ၦ4ml��7�oN�6��c�F�a'Y[�V+i�j-	Pݻt`ݼ�g6��٫��̽���je�CvTAV9��[�h6�M�zI�d�.#5e��V��E-�DbwW!�20�Z\˨���8�XUt��x����{��3B�`m� 5t�v�yH鎚V݇�*�l9�$CyDG��n�jŊY[E;[C�Yi5�\4�X�(h��m�B�h^뛇b�)�F䠆�&<����qU���KDZ�ImMF���F���4�Բ�<ثy�^$q�م=���ʹ���s]��u�[�Q�v�uGV�X�&d��I �!��Z-;�XM
�4���>�B��uA�2�Ѱ��]k2�q+0Ȓ�]�HYx�aؼX�-�������"ƕ7��Y���kux�+�����6���$Uu�z5e"��틧�Ik#j�%(� fY+6XԨ7Z��j���t��&b�0�L[.ڻJۅ�-���YVe�Z)ӛd$n���݋�{�iIy��,̫�)Ӛ,nA����c��<��/+#&��7h�TU4M�Żwd@ࡤ*wX� �y����r!B�K�����r�r�2>��(%)O.�˷�(�<�R	1�d���2��q7�Z��v�Ec;mڨYW���+d���'�{����xn���L�'��4mm92��͊�v�S:��aY�d����5��5���4i��Jn"ʴ��W����z�Gp�r�Yu@-Ů�N�&�l0p.��Q"�+^�_[z�r�h�J��Ʋ�ԡ��)x��bSC;f<�4��X[�C$CZ�P�q�i���� X�C+*-G
�]���l�f�oE���mޘ����W'������5}��+\�g��bBJ�2*���)���B.cE��Wa�/]u��ֆU�=��5K�T���m� *O6�5�6yf)���vj&���\��]*�[(�f��f�)E_�� a�f��2�t웸�8o*Sƃ��#N����W!�&6�K+�Lb�-#P3u�LT�F�XEŢMpAB`��ԩ/!�m�x6`��k��*�$~ҒtK�Ȱ���M5�+]�om�k&�jDH�+r���}-� �F����g�hefCZ�t*��b���kn������-�R�rM��iPx��el�8#�1�M�Q�j��@�e諫��ش5��i�,�K���Z�n��֍�6˼�t� ��ʤ��`�Rӂ�/n�����ik�3jL�֞�j	v��1V]��0�S�+5-�¯$],zhn��wG�-iRNB�X��M���%٥2��q�1�%l�H]h!��r�jY�j�֩3-^J�"�>ۺ"li(XS��� Sn����^)ip��*ZN�,vp�]%�X��v�nY���]��L,����܊�*��1fXjXn!BT�oC���@0LQ�U�����A^��
�ɽ�!bS�˅�e���6��tK��7e�*a��r����嗴R�Z�:˄��fśMR�拤%dЎ^Q)���ɒ�6.�,o[�ܝm�`ӣ�\�<wv�E�LE��9qTu���Z�d�r�^��;�F���Sq˺2��Z��=lhܲ��z����قf�����5��V�ӈE)��M\��+wh�E���v�'˖rdst��"�r��X��-6n@�V�wf�ЙzQYٺ���Ǽ��/2[�G�ĵ��p��u�o*ҫ�3鹌����;��ʔֱ�T�[ܻGP6�-��xsp���{.Y��Oe�j)�^�e�1�ti
���Y�'�m^��[��c�kl��(��PG5�@^��%hj���yu����$֜�Y�ۊ�c�[��m�F�ǘ�����8I<\�����^��
�"��Y��1m kQo0�ib�]f;r�������!��v�+��o�u����j�o�鬟H�̩��bұ������r�R������#�M
�;ڼN����@�B3H/7"��Z��k^P�tǢYv.��Y,�gU���Y��#�Գ�Z�cV���5�kwTw@l䖳q�tͫb�9$a��s%��P�E��BV�]��Y���_f��BK8��n�ٸ�V1�1�T~w���;iɷz�aY���ۣ�5�4�	��U�;�/]�Z��8�=�R��:`��ٔ�E�aJQ�r8%GG&j��͂�@� ��$Ë/E@��i�iQ"�;+,�%Ϲ�������$�Y�Uԓ-=[��/,�XB�5Y�0zf=/�X�sʛkU���/�pSﰞL��ĳ�^�ز�4W2���O��g�,b����f ��¹��e��[?I��G�&]a)�E�o%�]�,lZ�h#넊�J��T��Wu)U��eL)[������ᦲ�� �U����f�I�yD$e@ٟ]mIOv��4�ͳ�⺒Ѐ�yi�%�ٶ�V�����ݥ`Иkd0�n�W��3�U��N�S[�c4�ʺ�c%8���o�\��'t@�xF= ��Xz�K��r���7Y6�n�"nU��M�V�W�$ӹMƫD�%�`я]�˽w��%#J�����z��M�řFe�����G�]�cgF`y�)cjJI虉�Ә�M�Jm�-|x�� ݑ��Z�Lp������yc8Aa���Knͥn���K$LX+`deɔ����k|���x�w���?�g�����_?��rS�$fO�!�G��f:�yl?�<�6g����}R�]JV[��E�'�g7��ݕA̗sx��⎾Č���&�]��#���VP��:ٲ��<����Jg>T���$��\��˸�i ��o��Ļn�/)��g1P�81��v�)|�Q妖*O�<y}q_Y����)L�4�Ô2^�wҶ�2�hu\���8tg�'�9#�,t\�\צ�4٦��7+Cq����Uu%	YH�[�:�8��#q9�]�"^�7�Vđg8�W^��w�p��[L�.���%v�L
��󯒻N�:g��\N�0*¥���o�'(P)�����RL@9��I�i�G-�Cs@!^�pՁ�����ҷ�6�Ԥ2�.v���K'�;�*T�}_�?�.�Xyh���C/��ouve�yl*��)[��b<W܆F������*�5� ~I �ή���Ya���-J�"��kOl��Y��N�u-;�3؈���[;sN^k����1��Y%�j0�/ld9���H�%����Zp����gl���6�֤)�֗J'p�6]�w:�s�|�c���T&�_9���©�X��f�nﶧ*lX{���zFڮVA��!{�4���Xhk��i��e�z֞��͔c5�c$ԙ��I��a(��L(m�v3#�.ꐺԨ�M��{e-Ճ�2�1%�,#J�;�8p(rxq��ډ<��.�G8��+���4mm7*ICN%I]ZT~��
����=3Wp�:@��vq�=�ʬ�7�ck��%�}%����t;�-��׮�+��Xi]�ѦcN`���[\��/y����[.�	��OrYb�K���ŀ�i�`�b��m���k
l�H��{����}���%����� �1<Ņb�CI]�t�K ��s�un1�X�nr���4�΋�Y{h���͜EYEd�K5��C�r���/�+[�Kk{IO��r�;\uK�#gbE\��$iQ�Aʽv��l��h�qpS���0U>w'm�#�t	�s
�zZ�69+�w]�9�;�c0��c�p�{\k�=:�h�8��Ddͺ]Y����ѱٝ��A�a���Vw#ց��ж���w�*Iq�4\_
�v��:���{g0n u�t��^'��-y���l)&��w����˪
�.��W'J[Ϋ$l�r_G�J=9���Ct�KrS�XԃU��v(�\��pU�t��?�1�k�d�R�~�5�Y.=y�s6U�Vz*�Qw6�lj�%�ē%�N���k�F%���^���\2�[�#�)��7/A��kmNc��u���n��'�Ù�0\�u����eCX����J�Q�>Y�x�[l�-F����lT��i���� ¯>��ZObm�Q,�iX�K��b��m���V�[�
��D�,��F�ɹƢq����B�l�Z��Ro-]��ܠu�9�O-����b�jt0�l��x7�r2�GWw`e�y4�M�o~�m��J�����Y���c��\���Y�x2 ʜs��|�ݍ�K�ZD����)#�$�� y����ӥ9n\��,���T��yysE�U.n�����h�K�3�Z�Q7��Ԝ�Ut��oU=�N�Z6��QF.����L���r����Ml�\�H�̹�f<����:�����VI9]�e4h7.�}f�ln�\��>r�����2� ��z���-�|w���'l���z[k�!E��X�x�������o=�q<q'kN�ja�ˊ>�탕��l34���x�J�{���0��/� ��i$d.ܻ���e��3i�7]���_]��fRw�`̬.\�� '�ѝP^�;��Z�Z�t2�o����gc�k7)vq3��}�qU�0W�%s9����|4gi'�C7s��`f\��$7YW�����WÞ�t����_ ���p:��H��b�	Uə���eY�N���́��noP_gӸ���:Sc@��
v�Ҋd���q�,맏4�u�T��"��� ���}D*D)���gc����1���r�ە�����7+l	�cpn,���u�(���ު��*ؕ,�>W����ƁI��z��Ձ[�¬L��O�a�������ɝ�vY�:��S�����I�Ю�U� �oB�M�5����/e�7R2��Q�_J�E���p��KA9������m�}��]��âl��ƒq>�K��n��A*�P�"pG6_R�\ɝ6J�ܧ�rT�Y��$[$���$�I$�I$�I$�P�+%t� ���$��I��[��|K�o��M�~��r{�8�.�wy�(c��͙���JLN�s��.r��x��6�G�S�uڂk�9�	 *H��Ȝ���x�~g���	&�X4ɶz��]�M��R��r���c���3bG��(7��wS~����Z�.����o�ὃ���k@�p�;�y8+�P���mEPͼ��e֦*pٔ�|���ٶ9v��*�5�"��(.�c�b�@R� ΂Ky��:m�
Ө�/��#�w��a��>��9g b��۝A���K�J֮@�ř!�&�{5]�p8����I��̻��<&P�R�8��.���gmc��:/�Z��iSeW���c�U4r�����r����p����Yc�.S%�pf��s^Ϟ)Ro+��y]�Dh�45T�Y�0��ۿܭf3ϱ"��\��`�]v�@��q����X�;�ou3!v���i�ݧ�/�(z���f������^��|�!��|޽Z�yxqwl��+~���ӅK�� %��/��bI!ߞ���֍��)j�(�@ ���3��O��g�ܯ����o0�kY��Y����_+K�Pn�X�U�ga�xҨ1n����� ���ɽ�]��'�#n���9�Ċp�����y�f<źXg�_S�^�߇3}�"[�.7	�qWGu�*]s��j�A�
�����b���3Cg@���~��t�o4
<�2�Л�z�w��+����|mq�{&]u;]L��q:�s����V��g<�]}��i�\���.wP��;���#�����
Vg<�a��.%Vʖ�Y�ͳrp����b�k+������sB�ך�>��
�r���R��I�'	4�����wY�uN؏j<O+��=x��F�h-�|��*��ǍM쮁���Nm�`P[��䨾�3u�Nܢ(�imާL�oj5�݂�a�q�ed�y�W'b"�e�W�CW`}�s�yr�����EY4[(j<��bdJ�V�y��c�ws��v�Do��R�ZY٢-���._SC��K9��KVX���C��J���<�K�7)ٰS@������!���tk�Z��C5��e�o���? �Jv����B
n��k�u�"�dk�G3���${M�N�\�u4���r�:�cA�y;y ���܋T&��'���j��O_�+0���Q��OXfU�k��9��@PwW�e��d#���8�y�v�q	�@�Y)���ˡfj��
Ř
ǜy�K�(^�r���9�\q��;r�_-p#Ilհ'&t�p�rm�eD�Zt�J&��#ap(�T:{G�WESY�#�p��]jj8���'���ween[��e��Ű�ˮs�Jy8����0;K��w���]����5v՞HK4��'$��J�;�up�Ws{C��l��wfCJ����\�Ŝ��wD�����K���V.Ά�iȈ�r�af�22����Ӓ��B���_%�ܮ47�mBY+_s��>�ȭ�#�E���ZH';k�YW\-tz]!j��Ct��d��Js|���L�*nYUm3�̄P��['^nWv�G_fd�U�����@s/\����;$�x�V��k���듧֭I`�6�qR���Ď�z��
����X&�,�[o���|���l��PY��^�64]��Cw3�S��2��R|�n�قҧ�n��<46�c��(�����ν	8R����kwn����2b���q���B���k����=��7Y,��9���f��)q7�(V��&j�$��V��xyJ�uZ�)���];�9��.N�FeeM�͘�*}\y����B�֓������-�+b�+�7GWV��B���Es�dG(��]`�n��f]��@Ȁd�S��PrGs�֚��=x��㽵qZt���R}���ۭ��̹�v3������c����']:Ǚ�WD�93��9����.Se��a��%C���ݳ��������G#-�l�X���Ptf8qF-%dVM�(U���M����"��Jb;"���qk��2!�	�Q���M��K@�
�cT����(E�Z
�
k�pW��`�33]s��c
o���E5fб6��Wc��uI��W�E�G�☷�2���4s��`����ኢgps���/n�Vr=B���+MZ��ۃ[���{VQ�m�)E0h�O+\�+�T픝UruuY��t�.�;�o}���������#fN����QtѝOS쨍�v�u7����sׇ/sWX3��Q�RD�/8����M�ڀ��&��k�\AS�K������WbfG�N�9H]`�)�[�6��/)C��a|c\�f�����BS䱑�����f���D� �')}�s��j��]��̣Ǯ��vЫ�.�u��7E0��c�M�Wl����L:jlf�&U���Wn.k�vZ�-԰�y(K��r�h��u��Ik!ݴm���T�XUe�穾[L�C��X9�Ҋ7�f�ǹǲ᜻F���c�w7
9`mFBu�P
.��f�_MU��(q)l^1��f�`��oK�/�F��0YJs��J�g�w`��3C%[��^`� ��˥��d}v�]�ѣDP��L�L��5�u֒q�z�
�,��]\e�n�q�.E�G)�
�]��w3y	����=����� ��坂���6�D,(u��lc��)�
��1�W}�Qy/A�k���3�ή��=MWZؐ�`���6=���"B1���U�� "�"��n�w��s�<�R5 ���W!�7u*�/6�;�9���&|`�1J*ށgC���b��8�ޖ2��ɩR�q�
��r>5�T�˘�ȧI��gU�9S����y�<��OE(,��[������pf�$柼�!V�)֝ʕP	F�3��J�xro,Զ��n:��VUgW��wK9L�	�1Rvq��[˸&���V�J�ʉ� ���̇fW^.b��vP�8�/��1v�t�����s-Y�k*S���Ve=�锘k%����C%�I�z��j�i����Uiܫ���@��]\�����@��zq5D�.e�=,�i �:��˺J�{Z�[����h�[3\Va{Nڲd�4��b�E(h���2K`�)\8��� �יw�mǓ/��y�B��w}�4��q���Q�6���I?37p�D7X�������ʭւ�+2ڬ@vB�_et�dÄX���4f,����7.���f��^���o_i�u���qk��4���:�]�f������Ekܛ�$�H��Q*���6RK*�������h�d?��<�g�������fvsnr�ż�/��4�VM��ʋ��`�̮�A��vc�ڵI��"Wo��\�g
���Fb�,�v��-���Ȃ�=��6&%9u�02#��j}�uz� �[+�R`��5]8�a��y�|�N��Pr������xT�)��ohr�dy�
�O��8�id�6������4,��Fiw&��K�ڍ\ю���G�7�u;j�)�M��	������ܞZ�h����}�.o$�v�3Pc�8q�4&��*qu�i�eIŻ�� $ȡ� Q�R�Z=K�m�f`��T�aQ�f%Y�,��\��k,E��qm�,V�[�0�4�2�X(�mĦ��lH"��DF^j��lK[[�#���RҔaG����%UkXbUV4Jk0�5p,�
T��-l�+�VYcJZDEɓ-Kf-�*�L˴���y�qF��V�6����4�d̪*4��YHe�Ց���aLd��*�)��� �ŀ�����6�0�dR�"�m���!�����_���w�*_�Oo�&͋�Ws�󏓁%F����)����������ڒ�%{@���K<�k��t���h6�!$)n�{�۾�[��lmz[J'�|��+{OJ��!���#K7�qN���ov��0�h���5ځ��!�tQ�ۚrש��L�_Έ�������Uon:�rN4YH_U��
_��U���m� �����,�Ǻy��<��w�c]nh	0��@y:Z�E:H��� ��-	�UĆdw}�ؒ�*Zv�ؕȕ��5�&cg�^Au=Db�4�V���o����X��^ȝ�K��.�cT��T��^���׈�C�h�7j�_w�<�5bU���#l���xd�t�/9{<T+����8��h_1YVF1u�@٥�\�Ś�c��eGn��j���w�S@Q�i��^$�u��z���@g�;~T�]��u�F.�W���N����X��㘽:�z[�x��Eg }v�>�rO&�McltNż�";�l�y�6��^�6F��ra������y�^K��fҗ���1��"���S�OޗfA��"������v��LdO�dj��$}l�h;��.�ԗ�Mj�g^Wd�2�X$Jذ���~�x����ݥxTW��:�_��*��f����@���ǈgZ��JK��7s�7>WY!ue;�w����C����Y���]�c��p۵,��eZ����&�O�;[1lW�ֱԪ�zH��h�ުԱݢ�����V76AW /��(�[*s�E���&5+k��|	g�9�M�Z5{*�t����2��I�]w��E6�k"��S^�Q�f&�q�xj4lo����z���AwZ�4(��*�KnuP�%g>�oG0���5�M����[�4ٝQ^�]����ς�J�I�*ҥ��V�PR��la��(�(�fN�D|z,fEu��Q����F��k/��=F�aG:.e�?Z��;�b��G���,%@lLR7�+\su�=u��m�wp� E|�o�w����ğ�3��8�гb�n�Q����v�,��H�^��6g�\H%Q�%s
�h�VY��f��y�`�JT��+;_��{�;���喥�f�h�V2�N�3/h�nv._T�0)�]�y�%*W�y��U�;����oS�|��JRBsv������+t��5eZ� ڷǊ3��p�%��%,�k�n���1����b5��=��2_
�(��>rJ���]���oȧr��D�G�xP��������x��s���0vC}]��`�:ĭ�7�l�<��:��+J�O��Ξ�&�zA�70��q��.�1\ ](�-J��g>V帲s7e�S��1��1��/���rr�B��q�R�4�<k�h>B����=^@E���#r����2�������L*Ǐ��먦<�F�J맽Ok1�u�6"v9�� ��xq��'�ڛ�i9�\��{��惢^R�X�x�h�D��0B���.��]�[RC��j.��fx���������)�~��Vsvi���{;*�[���ث�]�����SV	�Oe�e���]����t-�7xD�Au��K������rl�z�'����x3 ��ǩz��e��$�צ�t^y���XS�F�lļp�ʕ��n��	��^3GI��}�˴Nut:(��z�خ}^�12� #�#���w����ײ�YEKq���y��잧-S��,�$��sZ�۔���]����{���>�mf#��8D���a��VW[��\ƅ�a�O��֯���,6��l�|�hV���G�7(lnH�&nH�0�5mX��6��n�y��P��A���U��2y�B�ش�z�j c��פຶ��jeY|k���`�#�3Ҡ0b�5Fx����h^��f���+u8a/v���OT��z�X�a� �]����Ɗ��,z���wL��q��p�F���q�d�㰐of���`8r��5�bLҺQ�f`�2{k���=��s���$*ݰ��7�-ޗq�9F���Hļ�ԕGx����t�[��MY�&$���TS�qPS9�Z�k�<>���i��k����tiv�@����cs5[7��*¬��^�lm��p����DAj���x,��b`�_�ԡA����y�B���/�+듎^C!y.�Q<�]�6��>�ɥ����TJ���sϸ��ᙬw�~�y���u�g8���o݄�u11����n���mp�pt�UŞ��u.��U�d���Y=MV�Y����V8�;!�\fR�{��W:�@����٤�������4�A'��+�`�LQvl�X뫳��Ê6���8mwi9(5\N��t�-Ѡ��b��M�vXK�u�X��� J_azv�{`�ڔ8I>-=oLܩ���-��H����n�o;��T�l�k����F]��nN��v��P#YCs*-7�r�"���m��Ҳ�Y�E<Afn��J�ޜ����E.9ηKRË�!yݓ�l��J�S5��5���>���g����c����t/.o)R`�b��wgbˤ,'�������� nn匾�STc#��Ǟg�r
�)8a�OU�tR�q����kSȃ��:N��+V��oSk��U7�N7
��4Q�H��4�Y��Cf|���������C��!��[��%*F�\i*�Vx7��+kVF'	��R���0�a���-v^Vk���L<�8��t�w|�fjNv���"Z	��6�|�<S~X�h��r�\�I��*<��� ���3\o\}�X�K/����Ɂ�������>�@+�Y1��(u�Wi3T��+&�15J�U]\\ma�DƎf�a�ZT���$Q��]��1T���m�d�q&bAuh(��Y�M�AEPwaD
��)1Ta�J�J+:r1Q�4�N!��T�U�r��H��U$�6�S-TD*B,�UCLuEFЗT��R�
�T+ *��g՞�����"b�zB��X���:j�̤QnR��^������j���2���U�^�ԲȤw�k.�J�O��x~Iu���˯����_�6�W��
��O�c~jP��%�#k���s��rq�!���Q�u��*ᗐ�u����Q���
h{��=�<���:��wE_�F��qgB�3��VH)�ā�U<��3�tN9uqv��>�0��N+��w�����]�v�{��ɨeg]kP:f5�@��G%rp���^��vI���/�WgC���+��bs�.�i=8{ެ�خ_@[{�J�����M=l��{�ɓw*yf�nD��+����`�l�7� ��z(܂[����9��XCx���r�5�_���R�7�u�����D�t8ZP���Wt$���%�='ŭ�	�U�y�>8��[���������x'{�������ݕy��Xm�����V��Y��M�M�R�r�=�J��}Q�%�7����u���
�Z��� ����k���Ǹb7�+d�ٌ����t�>�э�AX�uZl��"}C�;�NC#��CZ�I�k�����rP�i�,�vsi+����������mu�N�O�;^\B����c2��w�t�5�E�{*��~z��������;�#���d*ҾPȜ�(9�8��s'e�~|k{�����-j�9r߳��Bݡ�~��o{��ƽ��[1f}��F�����n��s~���<� �'5�y�����>d�Y4�P��m��l�Đ��!������3G�~��o��8�x��2~Im��@�H|�8�=�����o�����@�$���!�
��� �q����l�04�m�Y ��c {������y��C��Cl��x�z��ԇXL��R|�OY!�&��C���.��I�a�@�XOP�HCĞ�yO�C�0=@>IP9�$>��������t$�u<g�L�����C����:���� �����V <m��UӼ��L>�(���I3��0=�Vo�e,�3݂��=c u��-YN�l������?_�����CL&!+
�?2i���t��!f�O�s5y����{��I��$�%@*I�i`L�?2d�	�CHM��������پ��ć~��!���'�&��C&2m��O�a�}�x�0���x����x�;� |Ì�8�P���!�&��4�m����huo}�.���~���X7Bx�f��}g�@�Y!s�$8���C*�;|�繜�w�����~M���� o�!�'�kt��Ւ@�I��La���{��u��龜FO0ē�I6����$.P��3�Y<d5�$/n�A`z�{�����w�~��M'̜d��R2�$�B�~�35a�@��C0�׽�{������ԛgXJ�|ɱ�:��$�a�B',2�������;��CĐ�|�z���RN�d=C�z�8�i$���!��������<��k��<�(aǊpÊ�7%��N��]�1sg=��롳��Ԗp\�/��Q� �o�=�߿��7���$<d&$�?����I�Y�C�����$8��Hz$�u�^w>��?��8�������a� ��3�$6Τ=Ho�RL��|�P���K����!��N2J2ABq���!}�1����0���P�X���ϻ�����I�Y'FBx�+$?!���M��ē�����ގ���7�~����aԓ��NO�!yd�a*I:��	��ā�!�C��������!�l��7i�l�`|�g��8ɡ	+$�d&����|�=��^��~���P;����8¤n�0�v����1�`o��~ֻ����A��q h�d?0i z���!wO����$<d�$����k��\�='�%g�%`O���$1���O~Bxn�>C;gP��ެ�9sۏ3�y�$��P�H	8�|�����a�@��!�Y<e/�_}B;���~x��S�N_b�0^mN
��v0p����.�� #��=W*�w*dT��Y(���������|�2O�b�8�M�4�I&��>�b������3�����ёu��ɢ{���3z�9����X~����u�\-ACj��}�(Oj'(щԯtF��׷E�A~�7^���We�w\�N���mz��������iRϺ�i,�Th���\�({%粭�	��d����L� ��꘩s�L�&x�5���c��iY{�d�(�2�Zg�����]�{�>��B��j�Ѳ�爢|�t/h�����꫙o�P�������>n����W~B���j��K<k�v��T���t�,~�C��[��'_����J��_�p���]��8�x4����wݝ�9�C+Q��%�Ȯ߳�(r�b�m&��y�OVT�
�G�<�	�	{YKL��ԥ;tkt$�^���g^��531�9���y8�E�m}ថM}�ά>�G���9:-p�v[SWe�%wIJs���Ҿ������?����0Ew��Ѹ��&����Y���H�����8�p��Tǭ��+H����bJ>����̋xRO�ۼ�w2��gf#l�P��-�����4D��Ox�^�=.����kd2�����t����\�2�$~�>�vطl4y�A�9"s�\Q�m����x0z�j�~<As�D>�Ì�8K���:��]A,Y��ŃLش�v�3���Z1�yJ��22�暎O�W�W�C��'��wu���
)��6����2q�[$�D.�Q���=���O/��<8VP��D��l�)�=�ay5�n�Н[>W���Cٳ��&yfۡ�,�r�XP}=��vVm��ۛ���_P����2�#i|����7n�t�ꚣh�ڋji5dg����H��!��SrJ�N��%t��~+Eز3$ ҇�J�9�j��s6�o��^��EYnT}h�#�W �ѩ�bF\�9�Ӝ�z��#re�����]���3��*E��gA�k2���K�KW[��7`Xgf�m�tyk��uc7�vgi=�A���Z%�V�H,��jg{ո��cMuf,�Pib�Z+Gͮ���s��i�g�k 9��_t�I��#Б�Pp������g8پcA���L݃�oYk��m�ۍluj�%˔���~��XkRt�Vh�v�Y���ݢ�ׁܷ͡��
SR�r��V�ٖ��c��t�h����e��֫��z���u��dٿ��&e= u�)�e7]w�I����XOA�S �H��� �(��˔M�*��ff �����s�z��#m0��%���b+������ׯ�ӽ�]�:굮�|m���64�M��8qˈ#
ُtݽ�V���Lleλ20,����U$�hJ<f�9�%�]Ոn320ik�אַ���N���T���$1�R�׏C�Y��u�	" �bm�m��ȷ奲�I6��N�ᜓ�B�D�ʓ/0Ȣ]��H2ٽ��雕���|W��Z������F�Ѭ8�*"R���Lq�j�M2c�@�+0Ę��(6�b�L˘(��Xj�հ��,��J�b�٤#h6ʊ���]f���QIU ��@�jɫd�""�
�� i
1Ab�b�	*%�Xc�@�X*ɉPX(#YX�V(�U�B�mbATTDUdbT�)�(�T >���8)���nvR��R���ɜ�q�m��6�M�E}_}U��~�z]�����ᮋE����s��}�R�{���%Vκ\͜�j��oq�M���`�wL�-�p�L^�pv�.�w�d-
�k�5�A��6��+b器"���b.��1-ޮC��O5]���{��w:�B~Z���AR%Hd�M���fici����j��C��^Q�~DY�F�:潬�iÛͻ}��S��nèl�D\��Cje��g���d��9"s���������Xj4�gn�����z�"�Q���{^ȀyԳQ��.�C�<eq��w�5J�J�\J�Yfs��.����ں4��48;����]{��`����<�$�����3�S�B�w��~d�~ڱ��8z�n7�1췘�>�~4%z;~u��Mӕn���t7
f��<�R3in��+L9lQ��c�Y3�T�䨳�3k�/��Tn�VqT��oM6�������y:Y�3�3Ư����C�g<h�6!���Z��e�w��r�����3וy{ A��3�.;M,�^���/&�����j]�c<���XZּ0Q�wF���h��<��{����V�Gʕt�R���J];2M��i ���wҼ+�� �{>+U������<�e�u��.��]�r������F�>��>�A���+l�l*$��+��G��L��e�NA҄�ަ��着����
�x9bт�w�=��omr>ث`���xm�m쁷�%m�'�\W�̌�N�{��+=�5���p�x(N�v��p�^��k�$��I�9��d��O;�$Ms��-t�:��P�G��2�����\�OP�c�P{�j��A&6[H��O��o�	��}�{=���0��3Z̺�=�� V��ɻ��q�=N�;e[��-�j���2�lu{��[���Q�����������������~ʨ�\&�a���Qx����{)��ۼ��ۺ+a]%��Ӳ����sg��5�π�ʷ��*���viɏX�Qf����u�{�eY5j:ޫ�cL�^�zh\��[�[�0A�¢�q�Uk�j����{}I�L�}י�����o�BW6�7a�"�fA�s��5�f���F��7gj��	�ʂ�STY��%��\��q��y�Vȴ��"�ڮ�r�7��o2�I���������u�^�v͑�. H��%{O��x��
�X���Ĵ�ǻn�Ֆ�L��bt.
˭���R��9	#h1=���]�l. ��AdQ�n��pR�N��Y��*�9]WW����ms�@:$k���Bʗ�p����4/k�/ ZT�v1���Ͻ��g���/	{|��8!��\��q3��]�w ��af���N�mT̔�)y��:7(cnH��U�U}Y4t����}�W�vd����j_�&`��?q��VJ��p�Y׼WA��p؍kn�����ڀ������.�{d�c�Ǽ�G�knO8]�'��7���k$����P��4;�^����i��́��c[N� Gz�h�=��,��8��f��/�״>��4T4���U[�ND����2��7}�2�S*�ZS�E���m�O7�N�x��o��}_}�mz?�3ͪ�&���"�C>��gf5���V?f7��I��W	`vJQ����+9�Q��
�F3���O0�/&����|s��ZL�S��W��_F3h��o��!����S�u���n2�Ӧ.zu�iv��LK�p��jn=|��Ў��o{rCO��։0�O?Q7�Wq5��M�/
݅Sh'Ҏb�u&$@��땛-t��9+[D^nknStM�r~��������BƾS�G��/�E��6���2��~�zy�8w'����ĸ��2�i�n�u��M���
y�<�:�+�}�kfD8�t��+��S&�)���F	�����x��z��9L7�|�H=a�5���67���V��Ӷ�gn��j.zj��(ᓺT��!?e3��g��^�O+��
�Ai�3N5�,K�N�s��`�D71�L�ප�մXMU�I�������m��@U^������q�y`s<�H�M��W�9�fs����ٳ�n1������D�!{|}D~��RM���#A��\ǒ��ek�~^T>8|h��U�^A�.ؽ�s�Q�1�����3�٬ӯ���Iq��V0�<*gm�K�q��t�5������}��;1�(�k?=Y�v7t�Nr|��5�ޮ���s�l�N�1�ȴ���܆�T��><M�:l�Θ8���n�Q	X� �i��#@��ܣa��h�ή��<l��'B��Ow�!L�cN-�Xi,�C������+գ{h�
���h��+i��)cm��wr��4͜�x_�';A�Wݫwicȋ��&z�6[�����N�i]�#`=[�+�,ɋ��e�g�]����3�j*nV���㚸���C��s�m�I�� ge�����,sdp]*�N%�e��5{�f�9���Y]����x�3��ރ%iv���nq�1Ue�/�HeC���p���u��"���mmƴڱ�Y�M��!�YK�ѕ���bq]��븅Zb���Orb��"�[	c�w�Շ�]�S��26��r�4����yy��V/���"og=��V'�m�W�H^r����9x��ᴳtc�t_+"[Dś�Z��jlĖG�=cC�ُp�z�q,Q(�D�.���~��I&�j\���!�m�b�ۻ{�G�۝%�3T�rT���,z��Lg����E

AB"�VV(
)V���F����ʂ�d11�UR��aY*ERbQJ�ȰQdFA`���i(�XT�PQ`
,�� Y�0� ����&�1X"�
(DdRU�?��>��+z)�4B�ga�����1']��A7���US��?���_��ߕq�����@��5�Ք�W/���~!�����j��\rZ<o�$��_9���}�%	�ͫ~=J��^��˞��T'�p��K���=�2v��.�{�����KЇ��B��}��럻I���elyh�2b۹K^��+���ߦ�|_������kȜ��iЫbFLUV��Z�,�U����[�IYL���8��0`�E+��ɛ�.��&K�SL����掍~J��I�9߱yE"=.�P�]F���m0���W�hznj�ߍ.�{7���R��*���'�Z�|ŕ꽷�>�l�L u?	�&*��8�/�OH_C�f��Μ�xU�`Z|�s�Z���Ǐ��yT˧�Z���c���0d���_�f�J�W���x5�k=�oc�fug����+�jf���I����W���Ng�.����7zme���v�Hܟ���������cF�~�آ�\�;��Sp�P���۱`����g�[�zZ���\��>������������E!YV@ݠ�+}�ŧ��U�����������3���4�˸�]	��G98S)��چT�4kHW��z��*aUH6��<���=�엒ۮVo�S���O.�B�+��yʹ����K<���u�)��qEC��yە�l���z�E�W�U}7@����/��W\w7W�B�����}�nC��\�'���Nh���M�R�B��)hh5V�c�S��l.��ͬZ=Vu
��2�g���m<��u-�63�i��&����i��S���ۓ5����[�}ǌ��5�`TI3�c�ܗ�r?`�8}"�U�@^����`�W���<�S�`m��e�}s����`�w\'!��1mf�� 9��R9?U}UW��yN��W��������P�귍�g��P+Bƛ?:p����Æ#6�/%�Z(,?p��* +�uP�3�v��#i�8P�+����1�>ϸ���w�X��i�-O�Y{��:��=s|�.�������R�6���|�;�xr�&\_�����h۟Y�O�����4{�멺yӹ�s��%�1U�x��DUA��Q��OԴ�|| �ܿ�������V>"���楼3�
�d:)8.WW^5h��j< ^�7%e]���y��_��de�-��.�k�嫅�cOw z9�>�,��^3�Dy�^&�m�����3��1��x3i]}z�Oyg�S���ϼy��i+�)�wbɪ�h�i5����q�����k����`�<k,��,SŞeN�]�>te�λ��W
�X5���!��W�V��B�xT"�QB��B��Q͸�&�k}қ5�j�uu ���}��|��g熷Ʊb3^&���4�p�W�1]��� � "���
�+�h֚B�`��x�hw^?X��)â��*���v��R��]}߽�zO�Y�OrTNRk�֯[�n�~~���D����kNh�
�U���aM��x���c%Röw�Ü!�t(ԙ҄�ֶ�}�}���b?~��`]~?p���+���஛�}�ٍ�6�a����V2�]_�%�(DxY�kz��
�#i�רk˴�i��Y���~�/I
`��x����]J^����4��򫃏�Oo����+D��� �~6iߞP�CQ�U�k`�@}�0Sf�\5��\��������5�����U�������3��{�QV�{��w����0A��95o��璬z]5p�W
�L�4ń
?<��|�=� ���*�ٮ*
P��u�N��#�<p����ɺ�A���I�:�>C�Ǔ���J�b:��o�P�"�2�m5�����=�2��ߎ�~�ZO�E.����k*;������W��\4}�ت����\���b0xT�u�������rƷ��}u[�4�Z"�̔g<��xs]{�5�㦸��﮽e������<����A��������G
�z(�p�s�6�A��/W]�	u<:�༬���Q���Xg/��%.���厼�y����9�oϾ>���5�*m��t����5.w3�Xy��;ö�:(�CEY)e� }LW}����*�Mf���JZK>y�gE4��N��7� ё��\pI��Y�lo�Ax��ͤBo��WvA��&�� �R���+]#PAH`n��E��o�3��)�/�Si��㛥>������.Bw���Ç�z���������!ʒꇥ���4k�R��\ �"�:*����t�����$T)u��1`k��R9���QW=�kG�h�
���d4��e�{��`��uLW�/�4��Ҳm>ȼ>��G���]h�;�c�}}��?EӄG��r�`�q���d�,�D��ꁎ�[�uߝ'_<7�~��;�)�L��I�j�Zͫw��Z���FʼUbyC�����f�vo7�p-�L�-)$n~������B��~�r��o��6*�}~3/������i���#TbZh�t�Ov0p��_�^�a�:~k�������}Oe�p�4�r���8)
�de__�/_��$�}Ѭ._u52�ۣ�p��\�"��}�w��G{t�ju��r�1塯���1���PǴE8���,4ݖ�0{Ʋ�P�~�=�����ҏ]l2�S4hRk���	�u�1�z�˸eM5ve
��f�a�g�a�-��P��}�ݻܧ�S�xv��ی�����n��g�^O�]�*Ȥ��s�9f�t�Z	^��)0Z%��bX�~����rL�S��ֆ&r$E���4����M�4m!ZT�?nVe��'Ф/�rE��������*�[2V5/�\�o��]�j=�`
!�vQR�kQ���
�Mcә.9Kw�9�� �L�Su�|MgVܦ$�ǈ��,�����Hp�w�g��j��3�{�N�
"n�D�����u�-S;�<H<9��� � }F���bt�ER$���v�_�.��C����`�����v�Z?����O���J���8��	�o��ͱ.+�v���ݷ�Ν�bR9��Nw)f��O�ꮄk6kxU�v���*ʮZ�W��6Y�B6��S{���t��X��[O��G3)K1�w���(F���{-�&�.�q0=Qm���ׁ��o�����U��>I=p�i7�b�K_\��Eu���-���Q��u2c�k[�	8wR2�B��B�J)Q9$��k��(�nIy�o�˛9=p����t��*,��09c�@卯�C�W�,�LJ�

�ŋ"'-�TPU (E&5�Ff��� [E��HVQ"����&8�m�B�FE�Q�U(����W�XXb,F�QHVE�.�1��O�&n�tʆ&&*+j�V�_������ѯ 7�L�u*)���������o���i�\G�y�1}N���'������@;���oһA؞
���(+���|+�$�h��oz)������=v��ǩ�5�v�{������`>�� �x@�F`��h���F���s��B����`[���=w���hS*�S��eTV�eu������}	�|�_���'�*��>�r�� ��������
���M�����>ӳe����.ߧeՊ�P�+B������N�cyM~>!u}~N;E?�=��O٘x�a���\��U��F�7
a�j���쭱�dՂc�N��o^�󒾀p	a.hz��Z��9����	97������w�b�R�l��`x�o-�M5��mu����v��������<p�0�v]R���\�0��tD��W׽zѢ*��|��@�'G��ʳGǇ +$� !R�M�>�Vx�PR>ax��� ��A_��r�L}�#܈��`��2�A�3s9�� �k�	B)��i���>�·4�`?yr�oMACƀ�iK�@����N(��4}�,U�HV�әpb5�\�Vו�Ⱥ��n?9���s)��i��x���.�{��u��I^�	�v�v1f�LL��k���P�/
^
���N��M�\���]Ke�v%sb�C5��������d��q��������_��;z�<����k����P��stR������~U�N�L�ɽ�+!��©r�(�8��d��}���Wz�A�MdZ4�hD�B��y�Dz�u�`xXA8"4��
��n��w/(8`�~@
�
4R��+ ����7@VW 4T��6O�8y���rn�o�)l����>F@VtW
"�c����R]c�7V>�]/�� �}�����x�� [�>�
c�ElA��V���y�'L]ׯ3�c��Ӱ_3R�W��݅*���M'}�K��9�Ǚuw����ܝf�i��y �����T���3�lj_뜧�k����uQ�Q+~?SMy�<���?o���\ @�ġ�u���>hP8i���7��o��a�5{�������^4�*Wb���l�/����W�R���Pe
�5!�`���U�:2͊ʕ��΅-��#4�"��1t�AF���B��!���>}�O�Z�u�-9�И��fac�s�ҙ߼��o/�kt��1�+�1��xҨj��Y�����}���|�����_�t��<��[���S����;��F`u�۱�w滳��'�4Z�Җjz,�ں�K�TG��8�\_	�ݺ2R|��bI�)Crr����<+?S�
�,b5���_S��w����-��2x����s���>��˧�LW�U1�w�wQ{�}�׆��a�)�ׯY���S�������ֱ~��n��n����a�<;}z������ξ=ߝ���\���_S���q|�nY�e5�j
c��c�(x�=~k��oƆ��3:Iu�
��H�+t`���3:3�Iu|t]lU��l�b�w]
B�T��w�{�I�@+<�܈
e�����'� �j���$�O^c56腜h��ˋ�G�2����PP�y�ߩ3i���Du<a
%����)�}�)�x�B����sڷ �K��5�Q�Q��|}~�=�4�lSN�?�o�9�a�0�/�=�~m�O?���8}�v��3M:����2_�ؤ�>}�@M<(%Ӻ��G�m<�4(��e|4��h��`��)�Z+<�g�5��&'��=�F�@Cw���lH�>�k��"�]g����he� b
��Pю��{�Vk��M�c QT�.f�Ō+���DX��T=WV*���
�,5z��s��6�7��;�/��u���,��zΩ�֛\��
����1��+Eg[W���^���:��Zm^=����;m����#f��_l�*�v#�T��gr���nL����۔�k�������1���ۣ�f�
�~F����_dݘE!D^^�2��=pVK�{���ځ�7�u���WK�HWx׬���7�����6'��}´[&�>y�5�}t� V��;Y�=���������c�E3�|v�#���K��V#�¼��i������[���W�L񬆫B�?:,hS������r�Ը�b�8�hSM0B��hDѣ;۰���i�R��@DO]`AWCZ���]][��L!�G���	K��T,o6P�R��W�`.Uʄ���Kr����^��/p�5�n�pD��;O��lۜ�˧��X���S{A���I�֫�Aee�a�~O�+<7-��#���01�^��Ӣ��<0W^�!G{�kY����8�i����2��R�Yf��x��]�\�d�s� &mׇ�Ka�b�&��Z+O�O<�M<.�h�BKc�+iQb�� p�17B�|����L1��@h��tA\'{B:�x ��>�g���?4h;Y�I���^�[�Q+����]n�|�~����{6n뇨W�i��DRV��;���f��R�|4T�"��W�e
�D~�^�f��y��N��aop��=����r���Rk�;F^B���]��+v㏜���w�������Є��p{�	������\��O����Y�#M ����ƯEi�k:)�#���T�(!Z(���Քi�'g7K��)E|(
���uK��wT|[/�뇷���+l�C���M��+�񤆿G���l!Z�u�.1_�1PV���	=n��zi�481��H ��6<�����f�P��M�Y����pO}���߻�x�Xk�q7�,*�x���ﳼF��u�^}��G��R�
�I3O�Z�@yoƴ-�G���k��:�c����6�Z$[��e���*�%�D�8M��6Bi:�4����Q�v��i
�Ѕ?��4Q�4V
#F
fo���Ly�����
�5�,T.��:�C6�E�J�O4b�#��`z��)��wSrr�x>�<*ɫ�[Ǵ��u����`��c|M�������q*mϯ\�^Zhߘy��J������=CEhc��ų႕��szO���!�ο�i���4z�Մ 6^֧��{��x0S��@}�|n���An�ܮ���v/-����G�̢~����0{�������K��F��ב��}z8}YU�\��4����;ׁ Ug���[�S�Ff�t1����k�a�a]�j��[bq�yO�6�h�9�8UA��f����vA�����v�R�G��Bю�)2�S*�E$2���'WT�����x���Õ}���̙��j��.�*����8Q��=5p�k�8�)Z(����9�yPr�o�}�����a��V�C$��°w)Ҵf'�7�a��S�n3JĶ� Rw�*mr� |-�{���g;J�T0���H�YVΠ;Gfuᾳ��!�R�鄣�iϳjI2���!�^o0Uҥ}��ᙠa��O���:_et#�w�Nb�2��!�qa�7ᖓ3u����
9�im�l��Xء�#���ͯ����c��un6�p���؍ݜVMs�-񤰕��4�z2P�su�����m��:����D�J]j[���d��p�-1��x.>9(���@���rM������,C白�Y��(�H�����E���۞d�q%v�7�\[TVl�=&g6G_)ytI緅����%n�8�S����iF�(��Ï���nIk{C�!�LQdR�K<4�A�r*|�f��+%r��c�?�MO��(x���t�i*m�� ��	�ɉm�\�2��["�*�s3bۦ
C`�L@�PX���˃��PSbM�SV�t��\�F�m�J@��@\nk%Er��Ԋc��f��e��#1%��C2�R�«�4�l�Ea���`�f����e��c��!a|�X��w�돱�6�H�֩�f��Ǉ�B�b����0���g�x8]�c��;��b�X�z�����&����?^�zW�`� ��>(u�� W����,��/F Mx}����B1Xb�ݍ�~��<g��*�ᷯ��/�{O�i�<�B�gz9��0Q�Hb���V�XVD \���X0}��:��*�u�Q�u,�M���A�����A�̬��٬��ƆܒX3u�4|G
���[s{y�iU�n���`�����+��n�w~�K{����{{��/.Nx���@��W,Ye^�]�Trr�s4���'qέ�7u�r���76w~��֞zX��^���.��"��b�'h)O�Fق��4��2��z�4d�LX���-��{=�^xT)$�A�PA��c����&v,�����Dh�>���(CP(X�J���G�nw~l�y���)��3�v�!�*�����o������@0��ظi�Lo�
C���O������"�M=5�h��W�n��BN[���C�C¼ |Pp�*Q�������z�,[4�z��
TuƔ��ozsѡ
�F��h\i�:����aK�h��kǯ7f��}10�i2�쒦>�Jwr�mj�3�]�184���m��)�1�k�Ȥ�����{=�X?q�ZxxDW�ֳ�kt����]+N/[�TwV�2�**��u�F����˔��Ĥ��]���|��/�g��.����<j)���bޛ��ށ*�cs$_�ꏌe
�D!V8sO�������~��#���2���F�=���i�E ���.?h�m�L� yL�)����B�]S4aC�B,���e
b��e�M���v���3v|���S��ӗ��-�7_y����/�Ǐ���r�:���u��V:�Н�G�]c�1Z몂��3���b����n�]X���Xg�<+.n�By�ѐ�"���B�zV_>KnW]�R>�����?�j^�p��(�(~1�d�B�+�'��=����w�k�y����n;�k���:��8�K�|+»�T�ç))m��S�#PW3��1(z�
��2(Y%
�Z<��fɤ)Ch���Ol���]gF
~��x�^�|�b�
V��=�$Q4b�g������
l��\��on�A�X<*��Ч׉���H�Pp�s�&���6��_��ۯ/P�.�3Mw��{Y��B�u�>�dXb���δ�+O�w[C����)H�����c�]b�ͥE��ia;Mv-�SN��+i�S��Ʉ�)��ﾹ����^�_~���g������So����}�7����s&j���bw��R��q�^}y���{���Ki�����_to=}��^k��c.��>>�����}"�DP��i�����/ňMߣ6zr�l�:>��Z�6P�����mL���qy~�W����m]���bgo:�~�o�w��M�8<jCAHp��t~���=8�zP�B���E��)Xt�M��w�`�B�tkO��ϩ��=g�����߹׬�u>o�c�o0[������)��w��^���Nf�NSb8��8C�������a9ʞV��:��v�h= o��������M� u��S���b/�l��3��q�g���tҔ{��W�ôDk�5 ���M1����Z�AFQ@��*�_���)�l��Ml�A
M7�}}x�5�]���k�y��e�i���{�6��6v��5c��`���gٓ�J�±�(`�C\7��h��#�P!^APt� x@F��!�����N��t���`B�(3W�c�J�G��^{Ӊ�n�������<inں�)��Y���"��5�+v�V
��
��q�TJrg��t�9z�<(���$�����r-��*I�;�7��rժ9�����~� ���|W�_�U<������x��6@�.i(���P�����k��,_�_�"5PD9���YZ>l��2��4Q���1V����=��Mk�ޢG
��*��]A��@h�'0��x|��u��_��__5xԭL��׹�S��y3J�����u���Ð���V�"�5���-KM��m��Z:m��4��J���G!�����Pcs=��B�q\)BE᪂#�(���}xVx/��@|�y�Qb������P堯5ܪ�~�Zo��U�h�,c5���&q�,�`�*��+�Vn����;�:��Y���_eq5�b��pp�Ӣ�(�r~����y�+�~�j�E_�υ~�=f�T>b�9^[��a������PÀ�����H�]�yV�,�Uaz�5�`��4��Aqс���y���������u�>S�=�5t}J�'�Xܗ�m:�KƼ/�t5v
x|�
�1E]�ۃ���� Et*�M����9n����3O�����}�=Nn�EA�7+u��R��p�j
�٣CCH���w[�,�r�*s�M�Ǝ�bق��4�,:(�/��Xz|*�-��`��+�P�`���ϯ=�-F�I�}ޤ>��י���f���n�����жS���s�6��I��ԟy��~ ~�7�OƩ<���\q�?d��G��(���}1��V�Y&��׉���ǟ�z�k��u˧�)�֏�Z1,}�@����Z�pԎ����> �+Cy�;��u�/�~�:E���qp[\�TDw��`����<U��u�����: �y�G)yx�Y�G���]a�]�Au���ia���R!�*'N�I��B�����%׶���fZ1��G�0xUy��,����� �����T�i?]!��4E1��[Ve]*7Sv�f�{�)�-8w�=����*�ƨeq2�0�q8�̀�Z���շ5ffQ+zHzP��|���}C���z8~�k<��,T����G��DM�'$�� ��~m]P�ŢŊ�@��^+�&D_(a���� ;wZ aЁ��(���k�g�"��L>��8�(��>x�����߿s�9�1��x��8�&{x>
wqa+��5_�
c��C�0W�h;wX�����W�¯ŀ,U��(8T4K5���=���w��q�]#f����'�a�����������L���A]Z|�d4EhC�wj\'3ˤ�(�Oc�5h�`����#XUL�_NnXڽ��w�TΈ`�����pl�Ľ8o��H:r%�Q�.���8��3*�R���p�3����
����8��Ѵ��5׏�]S�����]�;�q���[|񾘟'H���(�W�W�t�.[�m�h��Y/a��oLRh�s�J��!8�Lc4�nl�b�<E��Q'8��}�YJ3X�;�CU�?mN�7��.hO�ͳ���[T���3^>�q#�ٶ�`N�ϊ��9�v�^����o)�2�7�cV�]����v���*&ɠ����z3*U�3a�|8�,���}]|Ʊ��cǕϕ��[����ˡL��r���(��oǎf���ʔ��E{���;���A�����(J腪�/4ɛEd���u�쵸�ƋmT�׮p�N��oZ����t��fi.��(G�G�JWGIAE��5�V��T�4�Q�5�V�f-
�Z$��Ÿk�E���q)>ADȴя���"�M����}gڒQ	���o�����fjO�'�=�j.�m[I�]�7x6�$�i��~OQa��-�m6�2�t�e4?�o�B�,��)0{3 ��oj]�r���O����B3�T�y}N�R�9&[*Jե�YU���b
WT1%`c]��5�9�,���µ[�̳��l����ֵ��m3228ʗ+����72.9�L�Zb��i��nc��&����eˊ�̸�ݔ������[i*,�m+����ŘԶ�n(�c&m��]h�-�&��չ�ɧM0��kEJ�����\[j�k��z��aX���ܩ,���C��?az}|��͙F�����}���vK��`�k>k�"��� "?
�;��wx�����ۣAM?"H�E�_���l֫�ar�릏�NQ�Y4� 
�u����@��<4*�ǅ=v�!Hx\�LO� \��T �it�����>�fY�^L�bu/� $k�~T<+�	�؏F����z�;?f��~A8v��=������������烷z)ޖ�a�.��Oy���}������y�;Eu��L���u��pn�>�H��Fj3�x�V˨-�>b�*}*�Uu�GR^���B�^�껉>֍�\�ô>K�&�\%��o^Ȏ���^�i�諭y�O�&�ل�k(������n䏐O��8eh��|��8Or�~��V���{5kuw�ʷ?��oDMg�����j��Y5�yEߵ�g���,"_�[�|�-2 xt�4us����{����.����b:�>Z��QW�E!��C7(yh�)�s��gl�D��9N�n8��>B�� q��m2�{݊�.n�q�1�X��&��J�-�:��b's�q[73S.]KS��^�Sl��UWאt�'�v?CC��:��e]S���d�0��զ�t��X�?zc1�.��5Ԝ����X�>���YK�$!	<��븏
�X�@���SD,�wk�֯q�Z:�Hb����s�i߳���8�6���L��D��,�T�}�Z����vm��������� ��>iqW!�վ@؀����7�ݫ�����Z�(�a ֓ۺ����Б�K����nVQ��R�t7o��?�I��g�Z�>�DH���{���h��,�{����L�b�V��d�q>��]����0W� ��xX�0����Ф��C}^�yP����[H�'�(+�&��vI����rt�}�	�ɛ�/���uul�����o��Z��w��v�3ãY�����*�
����L������eZ�{�P�1���#�W�.C�|fYOW�܁J&�9?U}�8B��/�N�u�ٗ寊/g=���9��^��l:�x�}� :�t��A��"Θ�����2-��e�ؼ��V�x �	s�
��a��+�cNB������~�Bd?zX0׵�Y���p�(����H��R�y�XK�uu�C�i$��~o�J�Z���a�~8�q�K�nV=y�=�po���3�;�];>SŰ(Z�`5a_So�Z��f:���W�+����5�����I��#XO~�
l�?�5���q���p�h�:�r��m��Ь|�;4�=]Q>>�g;X��jt�e�OP�B<'^��wf+�9R|[��޿��0V+�Ӟ	���҅:^�����;&�^$��n�y�6��&w=-�2���� �oЎo�Zk�.�]��xot��Uv]���ӣ�Y@�V$Pו� ��B�+&S��:}�I�ݗ1�\�|��]�ؠy����I?�}�W����a~�wߴ�f�f���'f��f$�K�[�*Ofo�ߒ"Nʽ���}/܇sB6�����7B��U�`��"�4.%ƻ���˞�5wJ|/Eһ4��*�2���ku�X�� �hQ� ��hNt���Xse��QQW7A�����3�����zJrǟ������%/��U�}ɗ�'z���춉缨g>��E��1�z�^��8M��i2�u�I6����̃�Bg�?~2�4�<<��nI��=�xr�կ]{m-���z���,������aPb�|�^=r�C����U�@[+sr��SC'}�ԉ�d�|�{�{��5��鑧r�s���#��P[��EG�5oÇ�[��5��c�(�f�$�@J@G�mN&K뤵���ieb�e��pߡ�ZkA�I�3�h���@t�0�8b�{(��k���8a|e�����Q���~���f������G���ض�?*��8"����=6
 ��N�0w��η�kZ\�Xұ%͢��{Ex�������[��A�o�_�)~_x`�7B�=hs�/��;g��/�|�zج2�ty�V�l�/����Ȯv��v0{w�){y���M�)�]�<'��O`aj�����X��	�w���a.�]KC�7Ο-�p�h��7�#]�op�MW���M������C�ٽ7�f��m��fgd�5� z*]�Ŕ��.|!7��S;U���>�2ϳ��柩��ud&jx��ә��oA�,�@��8�uw�4l�}ó� .q���E�Qέw�`-����r����=� 0]������ُ�-6ߗ���\
D���e풽�ï�߈�qw���:���7�^�*��۴�]NX짝��R�w���آT<��P�ɀ)g�Ӧ�_6�Y�[GT��/\�v�D��F*��Չ�ʔ��텨�՛���=w��O���h
,�]�.묜/�g0�|m|w��U�p>�.��S[|D ��w+D:�3dy�eN7&N���T�i;̺m�XI�$ٰB����V�ݱXk8G��"�f�����=��F=�X�'�Wf�$A��n5��LVv�W 7:�M��D�����u��v.�Fs�β~��5F(Ĭس7gn+�X;6
Ԩ��2���3�4w�0��#�]��l��]��v��.S���]Ļ�t���'`f�uꫪ1�'D�$|)wmf��W�G�\f��m�@�G��:�}�/:��g��>+zBdC�ԧ"�ed�/����n �jgZ5���qح����[vqX���O�������M�U�u��WM���͠�W
-�Vwe�1�;N��Z�Wt�
z�7������m���c�A�&q�QIZ�EX�57}Ҳt����s��дS�����ﻝ0.F�~�ř�0�˙)u�f6˔�LulSY�a�&�j���"�S1³"-j(�Y�ȿf���]8飡��5�`�V��e�6��kHEг*�D�JD�7HP��K�J�L�5�v��6b�1�2�:�r浚�b��Ŭ����Ŏ�Cnb�+��+��ĨZ�0��]�m�J*�m��Vf�4��"��x���h|��LWew(U#�c�ɲ�����Wޛ:��W������Bj�h5�'��߈���Y�F����J�xe���Rvk�������~rC{�c��e�[w��8�~���.�0��k=���.��ar3�L��zf&=HX��b���n`�$��e��3��Vz�p��������U��B�x����*M��
�{����r��v�C[��*�7k��13�� ������9�yP9vuۉ4����z*����r��@��4���I;��^*��n��<��c�wѵ�NO���y�)dv_s��6�,a#��l�5.R��~�n�+�C�a�7����[�{��"���J�٪	�U��������V2�A�� �U�56k�W�9����_��������p������g,��ɼ����ٛ1Yh���`�.����w�Kf��!�t�k�i�淸p/a�f���
��m�L^��O�;X��h���=�x����b�x�w.���e'�iVT!�U��"mI�@7kag����)	�D��]��s����k��;~؅��h�+�V��]��
�N�4�4��Z��=�m/w���	%tVL-����u]��?���o.���WGs���y��K��o�z��[E�Wř������uǫ�qYwQ���癩��)���l<G��X���'Y����R�JO�@fߺ�f��ͮ������՜z��â���sf�%��4{�{�Ag�r=�<�� �$m��?ɓ�*����3`;L��t~��`�>ûdg�b�����v�H��3�>j��˿Hb��������R���T���	�R�2e*�������5Њ�gzR���_6���nd��6a��+8muz�}���]Ϲfb^�mJ�1��3Vu�{��m��ӂv�
|���Z�b�����Q5^���OGj�;5�Xj���홨f���*n�m�������� ��C��kAXZާ6��8O+C�ŀ��%����s �k�P��i�cx];�0�m�z��=8�Y�*^�l�����[�=��j�lzv�mg�&e;�~ǽD���*�z� ��s9okF����a@/f*���vAbOq�y�x�ɒ�P]�{���jE��n)������>�n��_���=��Ѝ��؏�%��K����� 9�XX��׵�1]���waCH�-�7Sy���H�4}H�ݥd;NC��ݓ|=��(�W���.��nr����Ý��}��yt�F�r��.����}`3La���qv��;tʞէ�3�>˷���^�l�C�-oh��1-��z5fur.�ia�zD:�2m)�ȉk:U�G� ���nF��&��4�}]X�o#�ǧ7�0K�Y�}b���=�;|�I������f�ҕ[y9B�޹Wڷzz�}׾v�t����1�M,�Uܟ�DȟVU�p�~>�����-|���kŊ��)n� �52M�]���ע[,��:	r����-���|��mԡ/9ҧe�;���Z��>�v�u����M���ܭ|nf��S���X�=Њ�OWlJ��!���umL]�XB�I�(I�>�U����U� 7��1nm�L�w��c�[Dz�Wxf��s�__GKk�|�g��0JG�MhD������+=�(�Yp���q܇{F>)�K�a��D����Co�p?e�J���/�{��=���ɾK;�¯Ց5�=��E�I��Y�qE�^1`������<��[M��č�0P�-��n#z�8�q�d�d:��QY����y8�r��MG#�1��3}�xк�~���Yf�9�y$.�h���t�#��y@�=�[��_\��7�=�~�r�@k{:�U��e-ezt�4k6��Һ(�y�L4j�㗻!ޒ�iT{pxȒU�1Z2�g��t����ds�n}wg�hU�Y�c�J�x�=��u�^ƍ�{J�T���޹l���������T�X�^�	vŜ?�3r�\�G����do%�1�����1楶�K�/dmssݜ5�icxO`�}��Sb�7�@�]U��!a�o@�e/+�ξ�^�׻Ѫ�~]����Kk�f�(4SG�&��r��x�A�uf��Wb��-IgR�4����{gP|i�h��5�['L�Nf8^I@���%�ғ�KX��+��W&�z�{a���_�������}o��4�D���ɮ��c6��@N�,ˬEl'{`�x�5;���BqY2��DYf��puь�H�<N��a&�����Uj��߻�K4�`ɽ��ьG98��z�Xs ��U7��xM�
Wך%юd�=Ə�ͻ���=gt��	�A9(�ׯc	[ķ��	3����<�!�Oi/p�3�7K�1�vq������[�l睂��ϝ�O�oy�J+δ�.���E��1���ПR��û�ؑp�P�Gu������w3�iU��Á� N���J_u	��[[��^=��� �Z*[��t���^��쳛)L�����7��cj�
�,�F4ST���b�3{D�4��/i3!���T%]d�����]*-������2�ҥ)fd;e���%�Zy���kv�a�V�_�m7�(x��2�|xN�`�`}G�<*}\(^���*f1����	WVﱙ7R��Н��
�1�.���f����7��,1+8���?HΡ�P���F��\������4�@�m�-��iǭ�$w�^�i:Y�GlT�՛�q�4ppC��
�8���G�r�bf�*�P(ȰX�*Um�P2�
���-�KQY~�:"�dPY��Q\��6���k2�,n��h�!X�J4��j��]�̺LX��Y[�)��#[Y\LF&�k*��D�K�[���m��T�-p[q�*V�3-޳&��{ϼ3]�]u��_��E�9����������i;������p��;��z��u�g�Ε-��5��%� !lө޾D��z}k<��E����{�{b�B��=Y\b����=e�!u�-Q�W�Z���È�Y�e�A���Ӟ�;����,ݘ�%�>K�dC3�˽�n)�u/��։�ךw�[�TDR'��c/&q`y��T9�\F����*�����e���t�i�;�P�wLqY�vn��F�o4npF�r�Gp�_�ȧ��z9%7��~�}�V@�z�/ЯO��� ힺ�	�]g0��p��n��t)�עh�'Q�_�����U�Q ��ӈՊ6�^�Eϴ����/|�й;.��k骗���e5s��A%��.����7B�R�ˮ�4h�hU�V��~ٔgt����l���_��:��?�.�$hP�@3n���૬�gJ��nڰ,���MR�ZvsC�Z��=����	9���w��0��;�6�\�/��N�Y̎�Ó�+C��~��/hWZgn��=�S��R���F{5{�J��\�
c��L�#�;``V���w���i���V��;��H&�d=~m�)�*�C�{��h�8eW��7�5��rp��Z�f�W�JG�6�i�W���/'����^ڼM,{7��;#�TZ7�׈��+�,v�w�+z�f���,�*;���\خP�i����R<jP�^ו�n>V������T��׹vy���*���C��y��\}������\�q�n��mrO��w[�㊮U��ԫ��N��5ݍ�R���	-����)z�B�ݙy/6M�z���6��������4˅gT܃�`-���sK�W[��.�W�x�`��|d�=\��ZKW����+ڳ=ے��
Q>7�;�k��f�OL�,�����>���k�\|˫�����'\�͑��fn��-b��bv���$��R"���4�U�->�(�K����yV��Ƚ����Q�/�f+*�=��Ԉ4�	|=���d��$BZ8{��.D?x��f��ƞ�{ia�*�Tq*z�"]�0_|0X�_�W9�8+���[�%��2v]M^���L<[�9��S4�x/���*�~�X��.�m`{�V�&���)�n�i�t�P�ܑ8%�H��}��3�_�rY�{�*�-0��&k�W���V�W4Q>���r�;�xU���DdV��kU�3�����H�z��{W�bd"6z��'�}޸��g���j�{q��˵���v��#kE��%���+�j�hQ�|�MC�O��z��7B;e�sެ�Gz`�e�ɯ8��X�_C���$Uw��]�ޤ��V�$[��#,�r�_9G5G�	y��|�#8�s~Tpٚg�����#3�пIJ��KÑz �P��2�X���oG��{�X��Y�;��wi�m�|p�x{PK�������8A���B{�z�"�xd�[��ƫ۽X��5����y��j��n�yKƅ�\�=��:X�īѯV�'62���q)��9��HcF<d�gXGfi�xpɢ�d��"�w��f^�nStM�r\;��X�\�⌦{��!c�u�DM�*WXv���k���	�>m����ѭ�3[�N�"S��u���>��y�z-j8�u_�l�n�������\u�b��ai����F��eƲ�C�*T�J��cF	����JhF�y����v�-:3�?}�x�V#;�9~��,VEu��J�V
{�^��V����mX-p��9.�4%\��p���+8��z��et��@��G%K�9���|n���.D������?/�Wꃵt�^�շ�\�3=]���Oo
��nђD��#؟��V��� \���3X�B�
 �h�5j�.���g�%�iz�s3�i��y�����9&i֑{^��1n�/C����E@�@���8�׽�%p�h%���PZ��pR�w�n�ۙ�+heu*�a�O����2��dr���`D�K����9��`ĝwcM�b|�U�,i+9���B�'����h7[��-�� xۼ��Lx-��mԝ4e�{��υ@�)�¸�t�־F������ɍ�쿡���ǐ0�����H1�6��)�;J^\�0�~��*ߏ;�h�����3��i��P��e��vp��<F��ls˯I�~��Y?~���@�*�})��v%���͕��d1Z0>�M�xH�]��ՊLD��kv�ϕmG���׶�0Sz�MD�<�Ǹ+.gg[ k9d��J8�W3x�ҝ[Ct։q���N�̠���t�f�YdJ8rİ[yV�G�J��ۧ����:t-���.��X��k��x�����.��]uj8H&Kb�γ;ZX�E�h<�"��}���,a��c9r�gl�]iĨ9�M���R&2k78˾�_B���re*�T��r��`�W0�
:�{za]o'>�MT����;yC#��H%�z�Bn��
wL�����g�9t����9]Ycj��ސ���\�;Ӌ)�P�h�Y7�]���5�	��.�&�5I��5)��"烛�s�ٔ���ظ��H;;��A�ͬ<�U�d��D+ѢS=kk op^-�h�s��n�$����70��r���Q���6Ԩi�������P��k�l�j˹��v>�*�i��4��vMq��t�e7���s��:;u�� η"M��m6�M��2Xm��\R-�cE�M;;�csci���ҷ{E��\#r�uC��n�4S�>������p�WVE9y��[J�њ�l�r��F�r�3Ƣ�T����r�[�M��Z)��RҬQm�Dt����Ue-�K�TJ�aQ7L���LF]Ҫ�R�֬eun-��Vi̵�L��1�Kc+h*�:1D��e�Lh�-U�����ք�����f9�!���TwMe�5���QJъ����Ֆ��kQ-� ���8p�ih�rr�\V+�.E�5(ln8�nH�P��Ǽ)P�˯{��L�]�P.��JT�^#G;v�.�5��P���n�;����������W^\���9}|p��<ۮܫ��pl�\~#�RM��w�:�L�YZ��3L]e�nb0r���k}�{B��h���Ns�37��{@{Lg��~�p�.|p�#w깁a��j��ǐ�	-\�
�m��&,� �xm�!��<�[\sFf�=���旎�&�"�]s����5a:�A��t��"�)z���=�������MT�1�xQj�i�^v��^�^�H��Z�;�о�
�b�Y8{��sCH�U�Q_�l�k*{�/8�'��.�g�����������C����c*iv�|]2�Թ��2�#w�s��Ԧu�T��Jٓ��4r6p쨠ŋ�^�*��O~�NF����rgYd���2aз�T��-�]��c�`Xm�)3W̤Qn���1�Tf���Ѭ'޺����'�?v�І��>�����a�8ViCxO�/2�I��<Pg,VSY� ���9G��mk�Wޛ��|̆y2,-j��j�+�k�%Jxd�p�	�CM��]��y�'1O&��7ˠ�O�%j�l��c����#�u�+:�ص
t�9�E�=o���`΢�kV��W�{+� x�K��X0�VƸ�f����3'H��)�7O1�\�����o{�{g�j���R�m������F\EB���j��W GM\4B����Nօk����:^�^����p���w ����8xi�lo�����pf���I�a`��rn��윟ؙ�^R��x]9�АP<,_��[}��W��ZH��ȯ{h���b��h�=x�|E,����lu��T�dUֹ�o3j-�b)��͔o����+�܍G��=o=D.�2�*6U.�(�($�F-��	�Q���U�6�����Lfz��P=�Ľѓ(F�uˠ��o%���)��p�f��|J&�2����ǡ���y;�]
وУY�)\�y��u<˻�|z^u�锠z���*����b�5��c}�����S��=�g}�2��?U��V&�[if��ؕ嗫�wv,v��bgF��L|��F��jM�A�q�%Kܜx\x��
�[$^��Y{��zGx��C�ys�w�\��c��3���s��lʽέ.�]��O	���u����/�G������Kӻh{���]AE������>�6]�N���q��ygk�a��(B]�\4���Z7�E�p��N7[���גi��X�^
��dQ��l�j�Y
��F{��wj����3Fx���ZU�%�'.�0G�^gM�t�m�N�(��y�庰fÒk5f�HG��5P�|�}���9x��	˄��"�lG���=��a�d��B���)�啌�����}y" {�,P1H6S�1΄rSI��;yd�����
��{&���-�a�'�q�u���(��!��n��\z{}=)uw����̹RƏ����/8x�lK�B�b�\�Kve�&��FiaJeoIR�99Cz3!�ԹoG���\�7fzj#t�lL?z��3;r�y86����"���|N/Ԉu@b�U��4����w������+���n��N�SKk ��.���7�	�g��Ud]mz�I��0���B�[><���I�W`v㏽�E��m'n�g<ųݰOjuvy�]�0���=���JZGW�Y������/jVg�E��!\.SB�:1�4�0tv3�ne)���M�%N�0�Hsu&x���Y(Ze���rRق��'m_=�g^o���.�X{�{Y�V��Z�<�٪��b�mn��������Vu��LI���7��/�c�'�}0�8@{3)y����Rl^3^zm� �]�t}��E{`���9~��@�]���1sqz�L�\/C��Voe����q�	�
�%VZK��y4� j ��%S}����:�;���
�,ۭ7|]s��f�DX�f��PO��T�73g9�
e_�����L/j���M^y݁�]yoY��Ţ�N }�
�p0�5@ڣZ��]r��][B�3�J�]�\�>���*s�0���V��Z���C��}�y{�_������*��z⻯H.�7 }o%q����u��]�D�H}*�������><�;�|vg�j����i���?�*m+QE�U�,-��I$1��?愒I$z�(�k�$�H�eh�ʊT��2.X���_KneFU���OfI��lSe5���H�TI
�đ �HHF����	���a`��8���C�ތe�f�+�V@�7%�X{�^�$�H�RUo�(��qՍ��m=��E�F�a�YJ^g&:rQy�D3EM�?�=��P�?��)9>�Um$ӌXU�6�cI��� O�=�����$�o���hH ��Ri ��:b*��]�?����'�'�=��g���u�i�`�7��gg�$�I#Q����Qڤ�(mċ�B�]$a���%#IrY��]�0�֏j�/I���-n��Q��Ntt'}J4�ޮ��|�g/y]�O�D�I$SS��%&5��b��^Y�L��I']$D �?�tL�O�ҩ��(l?�<�Z��s|�h�Y�~���7<"I$�7ɜ��*����3�I�N����#kҥN�Mi����7�����ma�9��g��x޴��6o�J���zZJ��#�F�n�~h��+�dY�S��.�!i4#�ڷ�_6}]�d��q��ӆ��7��$�3��������$�H�:�%����J(���&����S�,6z�H���#-�$QK�x�I$���S�E5���D�J�#��-obXݒM^E51$o`<��}�@31�zQURl�WE�Q�jM�H�Rai0�
H��3�/-m�V�Tg{U�,(zJ�fd�^I�r��
K�Z��4�&�r��#���I$�6K�wS��ڑ�#��I$�l�y�~�$�r���R|�f���͜���M��>�qE��)72�W��Wi<�N�£��K���F_[�Te���I$���8�Ƹ�����Y����"I$�-'�}�j��1��m=�?�bpF��K�����i�ԣH*^)��fJ���vX�oPǧ��u�Q�����=/���w��j�h��,o˸ߜI$�E���Ҍ�.�ӧ�*��vg�F�=S���Ĝ6�GUE�nY�^v婄e��0�ݶ:(��	����R��\zy#]:��x�8�~go N�:���)3L��q��d��%fY&�PƗ�^���R�Q�O����"m�4��]��BA�A�,