BZh91AY&SYĻ���R߀`q���#� ����bFO�                  ���f��ڠ,cl�f�RM��M�����(D(�U[j6+Ri�DTU6eU[�EM�       
 ��wcZk@ �+iw�l�Z��[kI�A �4SkE��*�����H�Me���F��.��W�{�솖+\ wY�ҴV� U"�S�� .q�[J�� �馪A)h�u��k&���L�ֵ�0B&& Z�e�͡2���@ ʳ��     �I&� ͵�@���Ez����&��:4�q�:{lʧq]� �wF{���P��5J�:㺣�[�[�O4zӫ:�mmR�,�K��rЦ��$�@����� �^�{ב
�
��=۫�P���i�ݪth {���R��m^����t4����
���R�KB����+�U���z�W�hT���V��ejS`̭���I$ <@{��4(kT�����j^��y�|u {c>��hd�gg���]��R��w[ǎ�O@t{�>��O��U�><��(�����hԀS73�Kִo5���1���5�f�䔒 <�|��,�4���<w`R�뷖�*��ӡz��;@��d���T+ڼ���
�s����m��{��h�U^��[�kV�^���z��T�RPi�,�((�>R�����j�>��s}�%C��>�UD��ی�ஂ��^��g^� n�� u^ڃ{���P�����x� �ǥ�'�Z4��{�@U֥�y�[j��m��-��3��RH>�1@:�|�� q����q� �� ����4 �=Y��Q��7����k�L�&[ T[fm}�$�������OG��x =�{�C�J-��X (]=� �� =�w  ��׼�f��@��.�DMSiU�ض�}�c�  }�}� =�=n�4J�4{� )燸�A���@����Ow������ꚶ�Ū�-�)������) ��`�| �m� P;������^�{  ^����0 Ҁ8���| 4��� UԶm �fR�1���JF�3��>�8!� ���l�X� 6�p 	�� s�[�뫀 7\� �p �    � ���@� �JR�<��L�L d`'�¤���F���4ɦF����������� ��
IR� �    ��HMR    d MI��IHOCS)�I�'��#=M?_������������˪�?Bhx^�>Ž5�ߎ�{�>|������@@Uߐ��W���*~�EW�?�_�h$<?��'��?������3�S�����I=�4@U�O���O!ȟ (��߷��GO��SX:��&�5�0�&�8���5��`kX���F�u��bkX���&�u��0�&0u��`�X:��&��1��]`kX:���u��bk8��15��]b� ���`kX:��.�5��Mc�u��^15��Mb�X:�`kX<bkX:��&�c5��]b� ��5��`�f�u���5��`�X���15��bkX��&�5��MbkY�X:��&�5��c�N:�c`k#X����5��M`�`F��&�5��MbkX���.�x�b�X����5��M`�$`kX:���5��`kY�u��N15��bkX���'�\b�X:���5��]bcX����5���&�u���u��Mb�X�`��]bkX��щ�bkX:��.�u��c ��b�5��5��`���f�#X�q��]bkX:���8:������u��]bk�X8���5��]`kX:��F.�u��]b�X:���u��u���X���&�u��bkX���&�X1��`kX���&�u��`�X:���u��`c5��15��`kX���k���&�b�X���\���bkX����5��x������u�X:��8��&0u��`�X���X�`kX:���u�X���X����5��f�5���5��MbkX���\��&�5��`kX�`F&�5��M`�X���\H���5��`kX��`F�u��X�u��M`k���5��`kX���F�u��M`�X���&��u��MbkX���.�u��X����5��f�#X:���5��bq���&�5��`�X��c�k<bkX���&�u���$bkX:���u��M`�3X:���5��`�X�:��&�5��`�X��&�pu��bkX��&�u��1��`kX:��&��X��&�u��bkkX�bkX����15��`��&�u��c��)�SX�u��Xk15��]`�X���c�\bkX����u��a��5��`���u��x��X:��&�5��3X���&�u��MbkX:�XF�5��M`kX��:��5��bk ��bkX����&�5��M`kX����5��Mbc�&�8��&�5��M`kX�����5��MbkX����u����8��.�5��bkX����5��`�X���X<`��X����b�X���'����5��q���x���5��`�a�`�b�X:����X8���u��MbkXq��1��`�X����5��H뉬M`kX:��&�5��M`kX�X��&�5��M`kXǌ�&05��bkX���t`kX���5��M`0b�X����5��bk�&�5���u��bkX���k0u���bkX���&��F&�u��`�X:��\X���5��bkX����MbkX:���5��M`c`��Mb�X���1��5��`�X���&�0Mb�X��u��]b�5�����u��]`�Y���.�u��]`�X:��F.�u��b�X:��&��M`�X����u��\\b�X���&�u��a����u��Mb��&�u��1��`�]`�X��5�kX�����5��MbkX���&�u��MdbkX:��.�u��X��0��u��MbkX:��&���X�`�X���.��u��`���u��]c���u��`�X:��cX���X���.�5��Ma��q��`�X:����X8�5��b�X��3:�5��kX:����X&�]b���"�]b��u���Qш��E� ��X��]b�Tu�.�5��x�X���
�� :�GX� `��Tu��b�X �`��5��Q� ��XkM`�� �U5����(:�SX�kM`��5���A�:�X,b��D�*��X"kM`��5���D�*��X"kb�Q5�k�X �Mb	�E5���A�
��X(�`��\����5��bkX����5��M`c5��15��MbkX:���5��Mx�k:�5��b�X����0u��M`�X��&�u��`kY���&�u��Mb�X���8�X���X:��.�5��`��1��X�u��X:��k0u��]bkX:��&�u��1��bq��b�X:���5��c`�X:���u��bkX��`��u��b� ��u���`�5�k�!�Mb� �.�5�kX��k �'�5�kX��u�15��^0u��X:���CkX�u��`�X:��&�0u��]bkX���&�5����u��&�5��MbkX��5��달CX�u��]`q��q��f���#�]�H�����^y~��	���#K,|tf�`mV(�1���!5[둂 7G��4n�(5�a�B�����D��֣�G5<����kh�7w�M��ˬ���`��ƨ��w��wY��wX�m�kf"�ӽ�nb���H����r�*X�T�ef�'�iÏ�hXO�'��q&�]^�&',�{V*��CSde\5��d���c�#3m6S�ں�3L+4���`�h�V�ӰV֪��!���Xf�6�ј�pK���g���\��ƣ���<m�9��]�ڷ�����/:��|5$N`�K%ťu�٦r��(�����I��5���yQ�4�;3A��;�ص=eQ8X��^��S6R�Z��e�h��hQX��V�Cd�dLk��;������;B$n�I1]=v��(7(�V���4�^éĶ����]��Aݭ#5��)�ˇ�r��,�̙˥���1��;�c[-4<�2������J���@ؔ�	������qLæi�k�7n�u�͋���|I��a�lR!vdA6�M�������(́7$��6QH�R�)⛼���G`�����J����V���!YX��k6;/iv=ѹ�>LB�v���ZK-0G.̠.�ǭ���#��ܭ����[f��Ij��\r@l�4n&V�i6�w34�&�-6u2ܫ�ӧ��Q���.	��eӲV�V5;ӇB�a:�)���suRZ(��Vi�8_��M"�\�;�)��j���r�mdRX��������ğj�KT��8��4�WWV����D�r;���Vaq	�N�Q�,ʢ	س*�����M:n�i
*�P��m�0�U���mݽz�P۵LjĮ�Y"��QIXK�bٵ�I��Q�ĵ-s%�n��Iȅfh�2� ��U奈��Ջ	��z�Ro���{��Z㇋J�S����w����Inݦ�T^=.�k��(��م�%M���3w�4��6)o.�:�JNf�D�$Xo`��U75ͼ�Z��4dǚԻņ�19I����
�9��2c�juj9���p��J�P�΅�ˣH5ϛV�$f���T�]�V�ʃR�XԘ3!�Z�����ə�(��q���F��Q\HśW$���ُfIHD�PG&�í�'y�-݃��^��01d��B�8���Eb����Ó^�ҰoJv�GF�\+��.SHU�wv�Z����hP�Y��ܧW��ޠ�צ�+I&�<JI�N��
J=�]�vKcf�a,=s%���;�&�bYG��,{�b��e��WR��Lћ2EvTHV�:�U�b�͖�[>��/I��+��T�*��1*pm�6��6�n��Kř2�[�y!U�j��ی3�*��W5��5�j���.�j՘J��G�Vli�YT���+�sN�˸r�'ͼ�;RY��u�<u��%�ZF�5#���K,ɚ��N���Olͅmd�6�-`��{�V3e�՛Iڋv�l�jw���w3}�M��O��Q�e��)�-�:n$��W����	�%v�/�M=h^�Yj����7D� �6���sc;9Riwu6��wl�W�v���#�hZ�4NX��$�A�Mͥj��u����f1�Vj�M![�ز�v���u5�T�׉�X^��ﲍ�v��EY.�]"j�t,��Z�3F�kW�\J�Ե,�-����w*m�p�HT�s��t��=���*`�r]Kr�a�Q�����Ѫ�4��P�yL
��5P���b)<G+JZlԖ5�4��2�7d^��鳛����X�D��o�d�LR� ����yuo2��4/B�ݬ�Fqe�q^��đ�)�bz���LVe콹x6`� zl����c6o��Eu�k��1
�٩YA��&oR��R�2V�dahW��LX�i��O��1=��'0��j:��߉��
���E�䡘��ki��ô����)���*n��vd����I=�����S��TY�5e��ѯ&[�NR�I�W ���dj�a[���R������),��`ز��/d��n�&j&��]U��eq֛K.�J��ۗYI[��Y�$��.Bo���N�\E�t�		Y��dŖf6�fV`�,���"����>�'/WviG�= MX,��u��E;��b-��n'�am�!�t�9�6�E���TX⩂V�VT��ͅPj�,�$�3E:�:W���m�Tqn����O/^U�,)�f�uJWn�,CwTUj2��(�߯f��1e���ػg]֪c3!e,��zN��U`0�e�Xt�:m]Fm*��&�M��lֳ�j��ǌ�m�{���ܯClS���z�W+���%�9yI�M-���l�6]`�$ĥV+���"��g�$���w��%�i�〦�)n�݊���6��R��X��M7F�Y���yr���ț��-3+qYX�f�G+.Z�[.�m�4e��n�,eI6��^*u��i�U��͸�K��*�{e:�st���6��r���-wxݽF���j�e\�QX��ċ0��ZFR�Zj�n��acH������r�YCf	r�;Q��H�1���]!��9,�TR��RV� �m�u{ugۨ�uR�5�]h�V�v�B����{�mɣ��q�JͶy�W��]�(��c�IrQB[���n�b�){"���Ӟ����؋�s�[vq>.�-]f���ok�s���e�)��l:'Y�Fv�u��Z�3��MΑi�+�w�
k�R�`�mJ�{dY�fX�z\1]n#h�uM%U)�f�]
�ش�G��RFH�W�A8��j
bϷh���&��)�*e��-�/p7yH�I��u�oZ���Re�`�־��a���nR�TI�f޹�hU�t�-ѧ�c�J��dt�� 5v�:��qyCt�G*��@I4�0���k1[H�b�E��v�jRJ��j櫺�؍�w�d¨谅{See��!Eʥle�ޭh0]��Lf�5,,�b�6V!����TZ
\�$y�� ̫��9�*��`���W��ӏ:�%�����/9!F�����Y[��3;�2&(�)RL7U��-7{n�[ceX�M{W��������)�Y{��H�(��)��)۬qӱ����+]�D�
F�YBe�	�b�ЍV�^\cnbqX�PQ�C�F�T���%��ś}ͅV[kS���C��k�ͧ�a&��L�w
&M�Lj��-cH)21��m�Ƶj|tQ�o�U���N��Vm����QG����Ő�ј��ɉHm&#:��D��&�،�͗G)cRh���4Q��a�̳db�s9:��w���m�V���ת��$=2Ŝֆ4c�ORۋJ��݄a��C*ۅ֛�ij��w�=�zJ�����g�7L�Y�h�[-,���5�F�H��Ink���JS2��m\��//]�/q2Eʺ�w�B�!j9��ܵ7�1*�ݩ�[��̹)����FB���d�o�֮֝�|6�x]զʘ��d���.�L�v�h�T�ә2�ՠ���YY�P'�]ԖU6��p�&i���R�oN���V�l�T��"A�&�w'.�1�G$4D*zf`�&��њnѺ�δ�'`�L���u%�5K��Y%H7Pګ2(��Լ�#�y��?\Wu��r��f�c�{��g������H'�:Tj�W
�/v�A��a�<U�т� �k\�[\�Z�NUV��0�%��S���j����g*�n(!3#!-w���d��i�V⒱{�R0S�X�3x�&ƍ+Y�晅�-܇���m*Z��x��ljg�vk\b�i`��+�AC�S�H���"�PV�B�䭗x%���2��IT�k�X.*Q�r�r�p����$j��QЪ�6�["�́4��w{28��.��*^D�4&�ҷ���Bl\X���,�[��v;ɛzbY�d�V��;�`V�<aץ]��1�i;�kRG���n�nbo,�jڦaV���G������2,��%n#���Kj\����uVA��v'R�����I��-YyFz�7��X�"�$�\t���T�rpE��.V\��
A��,��]KT�N$�d�sr�/ʛ���Ͳ�5]a=�UX ����ȃ��˒�ԽZ�bJC���]k�Y�!���iF��R�z���VL��뽲2CT�hA�+3e�9���z��(��n�ۙ�&I*ﵮ6�3_j%j��EQ��Yb��jX��UfK��$ ØV@�,y��_�\��J)h6k)�/L9b솒شmc��$l�#nĥH�#tL������Zûr����&�20�Y�L�t���8�l��7���N��Ʀm�D�X�"ȭ��s$0��i�:E�.s�b����	#qz��A�t�F�ɸ�vAb�Sm�/4]�R�y�Q�X\��覓�AH�R�mG�V�EB.��ǥJ�Rj��m�[��f#�֦�I5�b����m�-���w���R<Mc�2�R7��!��x���6]��m*r�k2���d�m�ٶr�r7�Mܕ,��Ks��W�ʀ�2�k��X����f^�KDUmJ)�۵,JJS+f,�ʙr3�i�r�nX3<�-�h�()�č�Sl]�k0׵f��Ve��6�e�qQ�ecEa�Ȥ
�ތ��K*�\�z�w��3�,�V�9��&%�u��˻�W�V�3CU�Nq͇��4��]JpC"���W�g���d�i��%{4=̕��v�#��R�9f8�)��Q�%�ő�5��؇3\E��ӭ��R-��E�d��T��X�~�f���r��#��ed�ŭ����^'Y{4�z�^���i�z\��J�hR�%�yl�2k�mTJi\�����-T��7qط�4צ8�
�ҘP��1Ռ�Df;��Y�䥻�RWao�yЭZ���cl�u��*�Bv��U����A�2�2:�f��M�yKtIAш�fʷ���5r{�K�,�"�u(փ���C�y����x���V��2��R���$���:*��iE����2�26:�R�V���e�jjMD�-;U�6)IlJ�%��Wa����Ui�֩<�n�bԺ��i�R�ijT�U��KU%���H�ym��/9��cQ'�ud�R�n���KR)��J$�Ēz�)j�$�#�VڋUjT��I4l\�ԥT�RŜ�'ǘ�%����LYiܥ
F�ԵZJ��ܪsF�Ir4�T�q9۵"1k��%��f]V��	G\���Rv�0xt �����]�,I"D��_5i\X�	���֌�u)r�M)�uN[�j���jQf��b[KA�M����GĒ���J�T���u0hW��Lı$�ډm��$�����V�%�"6��"��
[5��Ji6Σ��ȥ�ĭbYj��Uҥ�f����KmNKQju�tm]�jU�����ľ=#�M8&IJ�X�/�%f�r�����-�I`;�R<�)�R�K���St��W�t�V��z�+qjN��6'Y`֮�v���V��X�*K)RX3�$�P/�*5��ZU��]�)�%�j6�;�mMI���6���U�+�>��sJ��Q
�E����jU��2�9.L�,�
�j�I;WL��X;I�ޥ�Z-,J�$�ؕ'Ƀ���L�T�������X(V���9P�E�%K�X��_���>�ҵ@���m(����oVڠj���IZNҵqe�I�i+[%T�Ղm&�)客�U��4�Z���I���S��-�{թ.Yib:�Uj�b���کkb���Dw$M+
b]ˁ�),^�V�S�m+XAũf#F�r��j��^5-h&��֟.�A���K%K�ԜOWܕ�I��^t��u����Uj�P���V'��E�)JD�K�����KW*Rf'ʬD�.�`���kb�H�HҮUc6meLN*\r���䦭՚�%��,��E���dޢ	�|��UFҤ�ĭ��R�Q�K)f��EV�7J�t�6��-���Q"5�LR�iR�{b�t�*�rN��"��+�9p�r�q&'x�.�v�`���%��V�K�P�ppui��V%J�o.��֦�MU4=���f�bz]D;�(���/�Z�SW�L{��H���\���J�;��]�+���ȗ+�Z�dT	��|z�0�I��`.%�IU,���U+���q%��X�����Eʁ`�#J���W�Uź�yDu`,(��J���RĶ$�;_!X�kV�j�Ě���U��.�j��],�o$�,�i/&Zr��+�U��V���t��
�u�f��:[��U#i�Rf�9[YX�U$�%���S�X�����*��jj\����v�Zz���r�S��i:Yj�]�1R6�ԵU��z�%%ne�J�Ǜ��B�Z�ڤT
�lYnM~�d�X�����u�iM�Uj�X5ib�L���Yi�e���A1.E���_.h�mQ��"��%�Z�"u��X�iZu�w��&��j�x��MI.O���)_'���<Ib赪K�_^ͬ�R��$�I��I^%K)x�ܹ/�ʎ��.��W{a���H�'R����]��u�Z��qv�[nlX�<�}nr�lM�J�,[J%�t����%h��:��D�W��H�ʎ|>��6�Z�F�\%�)J���ku�-�Ҕ���A����.X��]J��R|O<�a��uS�m���6e�|U�bn���-dJ��I*']bm(�("x�ԭm,�4�`=j�O��p5�D�$�M^mkK�bU���M,�-J�K��)���D�RjjZ���qJW�bV�%b�,Y��h;�r<,�弣HJ�1<�r�^�j�h'�u6���_+�Z��Y�1_&��t�-�RX�*�5e�/1@k��5$�*Ki+Z��i-J��9MejùBq����$r��_���%�Yj��+�NV��H���Mu$���AZ�)j�,T	�A�妑�T�J��Z��.�m��EַR�bT�[v ���y�`��Lpo�I;WĹV��;J��R|�%�ȳ�㵹%�q�^�$~�m|W����w���}�,��_~w�����I$�I$�I$�I1TRqŒ��9YV�y;'s�)q�S�tw��������5,=f>u��}��')���8��r���۵s��(P��i��L�pm��Z�LF.v��e��@a�bީ��*��H��(��S�L�������r�b��A%M}��ޫ�s�؈��U�^�&�J�+�Q/T��o-P����JX�-��3*���IC����_s+��k8B-;^�W��椬ř���n��噖�0�9Y
���ʀ�s����8^����Y��xz��a�� \��kzgK�U깩��郰�	8��:Im_;X��f�E�L�iD+8�)��;���&G������\��xJ�~H���IEEP���3t����WPX�����f��,�'3����v� ���.�i�z�)��v���oG� �`����^j`��ܸ�]���V=ã!D����r�ek�%ca�3 ����ZbY��7�%r)̢��%���3��o=J2r��銶�$�B'6^;�8&��"�B���r�͈�j#������:7Iќkr��9W��0g	e�д1g5X�^��W�rZ�Jދ�f6d!�^m�O���t�ν5Qʍ����v�>�h�]�*��J����%��>���xMG)���L9H��ѥi�
��]D���ţT��2Z�SU�v��w-w	���I^K
�q	%�:�\y���A���/m@��I�s�r�`%//E�Yy�Om��Jݫ�Tr�[�Sb����'cģ�K�6�v/��(�	��)2�7/	�O>ڝ�
�|xKG���ܴ�Jn��l>j<��q�<��3zp����Tʍ����-ҡ�+�#��[_-:�Ya�J��i�1B̠R���lvre�G]�Yo
)E�u�+�-���ʕt� ���u��w�m�"���6�}��A5�Jm��6�hݻ=�S9�J�*Ef��[�����9xjU�/1�X�+v�W�����<�[{"�����Vؕ�d���y�׭��E�80|�K�����+���6�*�������;���.e��ݼ���7���2��TB\�OV��J�U��kW>�>Kr��s�GD��X�c_|�՝Bt'����So�R�V�[���S�j���V�N�uB;��^?gYD&MP�6�yWn.�Z�f������6b��6ʋ�9����)"�*�3�Ԧ�G�͘6�����Fa�d�'[=��.�W{2�kj��%����|��.�G��O��O*FJ5���)K�b�BE.���͞��w��=]bi��Ykq��x�˼�:i6��I����8�U�[���r��o�v���mr��+|i�"luh,!����(`���/��t�A��W�6�F�m�=�����ޤ�U���R�Z�iw �v��s`�qt�od�Gv'>�s�N&M���M�WW�/KT���٘�4�J�p��NQ��PCO9.�'5�c��V	�����`C���K��#se@�-��u�}�Fk�N�/< ^�S�|b��nV`��Ҙv57Vᵽԫ�YX�*&�2̔�Y�S�_NU��#H���r'tz�\�w�tV�-�N�+ku�p�fvJt�m����u-���|5����&γ��%I�߷s^ɛG�re�q=VT[/zE���XY�Y��t3�����!-�%7=����Q̦�'{"�J`O�-�yY��p�\�D��`���)��ay9ݪg����Y�-M���vz��z��1�.�Z�xX���t4�'c׹�fK�㽔׬��mɺ�p(������6�!�ɨ��Ѭ��[�L�Hd=*+�B�]a�x�ve�q��-i"�hWo.�0��%���f��X}WG�T�Q��7.�;�sb9H�EZ��j�Vt7o"�ݮ�"�(�N��u,!�$�r�>$��k%�-��}R�G7��h��܆ul����KgI����g7K�J!������\g#:�l/�h�e��W�fвF�!ʵ�f]�4�Ta��!��
���\�M���o�w��7pb7wҝE\�w�<d<0'�d&t���5�X�
]�A^���Y���(�'RǱ�m�.��fJf�X}!v��r2�T�x�zV[\�������vT�x��A٬���9��.їl���i'Z�ZU��0]�װ�՚�ԫ<h��֮#D�3c��ςf�B�v�y�Տr�81Fo�gVa��7���j�^d�G"֥��*��Qs��;�/� '�M�ҩ��Y� V�y�N��CwӲ��՝o�.��e�Ք&f�!^u����O�Y5�1e�v�'mC�lʑ��r������SN#x������Ew�z�^7ܳpi�4M`�m�N3
�0�_U��UP�q�}�X��k�d(e �z�8+9l�ض7��7�©�+OR��JT����f���cN����=��O;,�b=���u5u���A�+�3��硡���J�U���AD��N��Ã�T��6���U��a������ׇ�6�EO�o���ڮ1WwtY�r��`��a�o�J�i[�uP�����r�u���Ӌ
8����v.��:-�֦釅��o�wCF�$MĨnjXT+��f�c�g�º�h����6�r����V�+D	}1B����?5����"������uf�ɵ�r�ۘs���Pb�8��9��Y��΢��*)E�ǥgZ�7\Z,>o�b39�|b��u؍�H��!4�nh%��*ɷ�����gn.�Z^G��R7.�t�ǐ#���D�ڂ]�S��<�l|l�k �/gSL&n�N��y�����!��+�3���-�eqZ�,��	���35
�o�{�sd[	����$�q����p��ۡ�!�����;ri���;bn��3��P�w��T��΃�v��/h�p��.�]p�w!ɣj;��ۥ�7n�h!WHMX�^�9��,'Nf��w��p�Emvm-�n��Ϋ@&|�T.�U��e�%�Of`m�\�*�6�����U��ڻ���ܤ�W[��\��P/�Rø��pe��w��ˇ ɹ.wu��Nu��ꎗb�+$FN�5��|�5ʮ�#O��5o3�ܱ7،G�բ�U�\'��
A֧�(��7��=FQ1a��6�iv �ʾ���n�uhd:|�wSt��3j�3(�Kt���T�nr�lv��2c�����|�w�����/����4�cd��]��%��̳�`/Zi���)t�g�0S���F�-�Ӣ�/�����Sl��7��w�.5�� J��d�W�}��2�w�Rӳ�$tQV+J۪Vzr\�:�4T�����a�l��:+'��1�!e���%
�]�ۥ�{ֶ]J���6�\���(���
��S����R�In�ST{7�^k�h��5��ŵ���W\Zt��O��2�=���@�<��ɥ�LrE;��v�c��N���	+��m�饓v
<1sg��i�L�=7�k�2�Fr7`.,�'�o=���S�+k��QS��D���]/3�('5]����g�K�����R͡�p�e%�W���71P��҆��YUF��a�5]���$A�ʚ�}_v��.�뚤�=�6ا����ڛ��=wzԧ�A�-S(�u�E�Hf�2�ɖ�x�]��%F�n��� �N��l�D�&�X{�lS����0�1q��DmM=@&ˤko���|�e\ɢ�Yx�d�PS���l���%a����(��E���	ӪmcZ���)����خ-x���j",o�G�y"�3q�¯�>e�7�o'HrKo�н"L���	�����2ᵚ.�"�\��h��Nc)\��F`��y,��ܱq��hͮ�Y����^�ִG��;��Ei;��j^��ծ�+��	w�"n0H�Mn�]]��l�ɵ6@�<�R��tF{�앆�gj�n���Z)Mܭwu\JAck<R�۶�A�
�7&R�{�VqMJ�,�˶-��:��|�(�������tz�g7!8'�nr��yMm�{�N���̥l��X{�wb�:n'#Rc�.����q�-��ڈ��+�:�[x�#�V����';dw\54�8W��\��9S��.]�9V��'m����Ղi�'׷��h��!g1��3��R��'��L��z^�52�j{B�_R�M�R�}�f�G8ƺl�B��Z� ��W6k rxp�����b�������Ήz�����㠩��W�M�(��L�s'ɇ(u�T�\�j�H�2��|fn�d�:]�'�Fk+k��s�+�rIAB�^���S�xV�ZC\�^L�O���lVy	�f�c}7.�OO�)O�ƻ����.�f+q�uf���1v�;��ZZ���e�Jw��tK���Fe�+�T,�zp�<��0ֹ"�"^��J[͈ͫ��K�F�ځ�Ss�'G(��w_gU��vS�t�3H�E�eٽ�WA2zX@�i��%ŝWO��Z2WcՖ���Xxhat-"���;�;���yyI[m��(�'K��H�Uq�b�X��[�!V/ �~��z��X�6Y(��+��u�@���)���2�/pGu1X���gf9�xm�x�1:�;�U.K[P�A̋���e6)��(�0�Ns�NͭҢ����勲.a��9_So-WJ���\�i�'�i�Pï;�`#1B��KdB��E,<�ŃHΦ��"Pj�7ہ�,㷼k�׹`ov��fS�R���w-�㾺���e�6���=���Yg.�F-�ɨg��K=�9��vL�5]\˱�op�B
q�Ry���{����V�8����Q啊n�w|�
kI<|�^{�c�gpI�Q��t�}n��n���<nn�[���5�Bo1��N�}�e�n(�0]�`Sf�]�*t�0���}�e�b��.\��#�}{�Q���Y�D� [��)P����A��xL��'(^�rI&�Gܜ�I$�I$�I$�I$�I$�I$�I$�I$�I$�H�l�$�h!8�`��k����.I%��n �S ��\ɑO<��N�=:�<�� ��z^f��-����xC>o\�2Π�H;᷾|�"lC<�L�~�`{�g�@��r�[s���>�iJ�5�Y����B�~�H~~��>C�Îe��{nm�"\��U�����|é�b�������g'����X�Q�y��IP����)���[�Ǔ#"��;�>s��b��<�Oy���/ɗȯpL��9�'�����	��|�D`=�{��'�C���P��o3���s��δ�����B����x@&�}���c���I9؀g��s��yx�[�KO��\�`Q�<<ێ[�,�]����|�<���+�+�}�d��ND8��>,���e{�qn�ߒ9��G�� 9�Ȳ��CS��<&ZY@\�r������D�'^�L;XG�P@��XS��H6���  �׏������j��U��OqȯQ�^�/ȃ��D����_��E�/�O����O�?q�G�)��(���_��#��?����~�����>w�����~y�^W���c����":�y"9��R���tS��v�,��e�裾'Y�]�*��%a����kR�܃yq�ם3/�Wt{zշ$�E���A�N� ��jKvӨ�,�c9���<k(�S�Ӥ���阮�[�=)F����,�Ƶ��eC�q���6��Lz�U.�}:%����j���e:���l��\C"��n�H	ݳ*iXҾh�O�y��D���gl��H�����Y�>�HTD�Y�����n�Orm�Z�Ő[�V�L;(�.�nͣ��UlkPsY�xU\�,���d�v�� �c��f����m��;�Ȥ�Һ�uzГ��gy��=�z��(�Lq*���;p�J�GR��M>��|.ur�kh����tἺ�Ebn���60,�[������j���e�t��WaKS�7�������yBc�2A�S�^��x�&��Ʈ���%�Le�mI�}Ԩ{�w&�a���к�Q�-�p��x��Fܚ�/�^�Q�՗Kj��T������);�����㮿__�}kƵ�k^�ֵֵ�xֵ�h�kZֵֺ�zkZ׍kZֿ5�kZֵ�kZֵ�kZ�5�kZ־4kZֵ�k�Xֵ�k_�k^5�k]kZֽ5�kƵ�k_�kֵ�kZ�5�k^�׷�kƵ�kZ�kZ�kZֿּkZֵֺ�zkZֵֺ�zkZ׍kZֿֵָ�k^�5�kZֽ��5�kZֵ�kZֵ�Ƶ��Zֽ=:�k�Z�ֵ�k�Zֵ�~5�xֵ�kZ�ֵָ�kZ�ֵָ�kZ�ֵָ�kZ�־<�
k�Iق�SW(��k�4b}�ý�T�4���zE��eW);$ըѩ�kL�ռ��6�c�ˏx
���*W1�k��<�΄U^�����3�b��X���^�v��m�*���]����S*�F<TM�#�`e�]�0O9�;�,�Vf�E!�ٮ�x�Lw2
��V��l��ɘ��b�+��U��Ɉ�ÉGP��cͤ�-v;wPF���Ne�@(�+r)�ou7R�*�usU.2#s'n>v#[Ld�yh��H��D��h #��v���\`���	V��>�懽���#�X���׬Qª҃��VsK-`�ud��Bޑ�D�v+��nT�5L��;�:�1�4G+r��PTYrb�<ii���d�p��hՔp�9cA����@j��|J���Uo��m����<@P��]^4]�jWiN卅�5�j�U-��tȐe]
ѷ\KȆ_�G�m��N��.�fC��]W��vRٴx��U����qӢ���7�ASq�e�e�$���ҎL�&��N��s�'�������ƾ5�kZֵ�mk�kZֵ�mk�kZֵ�ֵ�Zֵ�MkZ�Z��Ʊ�k�F��kZֵ�k^5�kZ�kZ�Zֵ�{hֵ�kZ�Ʊ�kZֿּkZֵ�k]kZ׍kZֿ5�kZֵ�kZֵ�kZ5�kZ5�|kֵ�k�kƵ�kZ׶�Ƶ�k^�ֵֵ�k�kZצ��kZֵ��ֵ�kZ֍kZֵ�|kֵ������ֽ5�kZ��Z׍kZֵ�kF��kZֵ�Zֵ�kZѭkZֵ�hֵ������~��ibk��hX�AJpqk�L��CD��V�����Zv�
ܳ��@�*�{]!t�x5g�b����.�Yc�ծ�@�t��~�ܔ�7�iP�@�(�n�޽�=��p�����Tu[8��ڬ��$[�܅e�F1��gf�������g[�َ@��=^s��_r����F.�������]V�W 2��4���H"��yV&���C1��Xf��i�p=3�����'���VG��.榪��Y��s,󻒒�j
R�UV=I�W�q�]I;�IY�q���6l��hNY���,�2�q}\k��4�;��ڵ���aٵ:����c��� �Uu���ݞ����Kf�m�p�w�(Y]�r8E�5� ����Z�!j���¬-/�FmKa�x����}
�ԪgVgd���@�c��z����-Zuu�v��;E�PI�i!-9���ΈR-���U��dSX�Wq��a�}F%ڲ�$Z��N;V�g�M�qE�+���`�%�'\�g�9n^�潱����־5�cZֵ�k�F��kZֵ�Zֵ�kZѭkZֵ�q�k^5�kZ�kZ׍kZֿֵ�zkZ�_�k^5ֵ�k�Z�ֵ�k�ZƵ�kZֵ�kZֵ�mk�kZֽ5�k�k\kZֵ�mֵ�kZֵ�kZֵ��ֵ�kZ֍kZֵ�kF��k�k^���ֵ�MkZ�ZּkZֵ�ֵƵ�kZ�ֵƵ�kZ�ѭkZ뮺��Z�Zֵ�kZѭkZֵ�kXֵ�kZ�ֱ�kZֵ�k�kZֵ�k�kZֵ��~�V{��7L2Y�e�p�s�|�7+L�bڑ���3㢦�u�$ٔ�ZAwe�<s�Jw����.�j�RwNf�ǩ�5���4R���n�]O'w�_
Z�U�J�a�p�r@��n�󧇪[ƹZJfX՜�Z�.p�t�Z�6�i��ǘ[���n�����ǈv�D�:�`l=����������+���j\����J�o��n��qWRf�-�����z�*#����˯}ί]�W)����znc�J ��� kq�Z�xL���[	Wk�\ؼr1�Y�u)�i)�,�r�n`��W�I�SEk��ܭT�����XW���3�p<I�Ki�o��ն���A�HJ۩{����x"����XqB�"������{+<RܫI�-�G��/mqѰ�4��á�]ep��m�b��� �]�q0-��P�h�̮�W�)��VC��7.�X���,J����9��@<�J�y�]7v˰����O,n�ي�n�ǩiˬç������w�L4��;R�� \��N����F��u����#clSEe-��Ư�\!�X�4����C2X��P�k���^��o�zkZ׍kZֿ�5�kZ־5�q�kZֽ��kZֵ�|hֵ�k_�k^5�kZ��Z׍kZֵ�|kֵ�k�kƵ�k�kZצ��xֵ�k^�5�kZֵ�ֵ�k^��ֵ���k^�ֵ�Zֵ�Ƶ�k�kZצ��5�kZ׶��5�kZ׶��kZֵ��ֵ�k^��ֵ�zkZ�kZֵ�Ƶ�ֵ���k^�ֵָ���]kZ5�kZֵ�k\kZֵ�mkZ�Zֵ�MkZ�Zֵ�MkZֽ5�k�kZ�Zֵ�O����u�yʼ�k�ab��z�Wm�r��D���f���G(��F��k�R��e���oU��u	��T�um�^z��r̜f��}���Kr̠֐�{޺y�(|�x��PFm�9}}8D�=���(s5�Av`���.�~�<�`�"ϡ�r�m[��a:!��k7{���z�j�qu!���[n����Nι-*��].�j��ǯ���R�t����-�C�W[���Eel��*B(�����v�l͸�i��n�*p��z��w<�T��,���MU�U,�'����ez���/Omx^f0�ݐyQM�H�	�x�7�i,�ۼֲ��͢�[�Z1=�$#M�ѩ������1�Sh�]*���!=�� b*H�v��{�e�����=r���T�K3���L�z�kDU�Ŝ	U�폱x{�ص���j�VI2P���uf�bu����ԕ�����/	Q�gEF����9��{�E��-�����e{6�2�d�6f�uT
�UI�9�&��03��Pژ�dm�e�$���������
	y��.n6���p�C4�P����R62ȭ��+q���M��1/7o���<!��{OB�����dw@��S�,LneD�=�)U��vsg���T
@���7:˿&�ry;;B��@�>'Ăie���U���m�ZM�ӫ�Jș�:.e��w[�������W�� z�A��q/��/[�&�X�V<'�C1 �"���Cޭ�b̣*H	'Z�7P��c����e:��d��V�R��u�vȻ��t�ѵS�9��!��t��r�z���]�_=R�Q�v.f��t۠"��s]�<��g�>4+<*�>�R���zm�u��H#��T�����7��6_�C�J�n>�Ӆ�90�T^�6r��:���^�U+Pj�h�sZF�)�U�6����P��(ۘp�ڧua����ᯊ0�����DE��P +�d�< G��vϺ�����u���l]z�l���0f!�+��4
���9��������n�P�/\���z�E��*weN��\"�Q�v�L��A�xƫz�Ԣ}o�^�/C������'v����9��n[�2���J�@���`�#!�]c%9x=�O6�mѼ�����+�s��Gt{�}�9p�lj�캣���ݑPDP�����G7�c1��{X�4�x�uiA�X*��Qԝ��sWD8�Z�S����6fY'���hT6-b����f:��)W^���D_\��C��Y���3`�z�\Q̴u(0���(�:�Y/��ګ�9\л�U���e����}b���;�X�%f�Z��saw�-�,!�겡*:�½&i��N����ҩ].P�y#�v�|f��f���Mx{��3�whJQl�5�U�(B3�NӲ�jͅ9Ә��V֬sK=Jnk:�lEsm]��lD.N������7��{7���[��n9�tOjs���A��=uQo�9���a���qlt��"�fhܙ{[~���s���:�@��ݤ-3��F;^�7ya�^	}:��[Yܯ�r�)ꊈ�N�@-u���u5�K�j��m�Ϛ*6T�N��]f��4�d1#�nʕ��>�;�+����v�������[�b=�'&�{��Q+����ŏh�؃�!]�Qd��l�Cw��.BX���p���қ�y�,���$T^flU�Gz+�^��u��D]nsP���K�YS)雖@W����ٞ��W�e`�'5�t�Ў��s�����"�x��	�ރ�՜4n <U�T��q�::ǝ�PZ�|�㼤�V�v-�5���FG�+�����=� $�!
LQ�}z\C-c�o�(Q�*t���ǹ�#�|=�酈#ت��K�FƷk��鋧y��4abM:3*A5���P�K���-	X]��9$Z�6���zJ�w�3
C�C%��ң:��&�q�iutFx�����)�����1+�*ld�4톩��½�(�S��&=���Z�]h1#����M�F���p�.�/lsY�Y�d���snUJ��Z���485��NJ�λ�a�m��8�}E$3��:�\\�&ܯq����<12k��&��v��Xœx����Y����L��H�0���թ��[}9X����5�,ך����|.��������F���K΃(K38 3��įc"$y�f���uvӹ��TU���.�+�6)�6����.��G�`2�;�
=2���]Ηq*c�Ǭ���gIx��i��g��Z��#Z�,�Xu��I��m�U�&v�(/;�Zj�PKBu�?x#��S�ʋ�Tv�-7��)�P���YN`������)�{)�
�x0��3�K�u��8� ��V�)v`^c𴚃w��\ܲ�Y\8X�é�qݤ��te#ԥڻ'mX8�\�}B#g��7m�,��1F-a=�u��R2I8��3g5�˱+�ۻ�%7��l��5C0�D4�5,%�\�y��%גY��R�7����z�Bº�i�	�<7�|�b%�x�n�5�"���W�v��6�;�P�(�z�����'�̳�ܒ�n�C��@u֤�.�s��Pnv���W�_���@rwj�`��[k}W��(�����C&8�AYEu�{t��Ět��1��xxl�3�
���n��\����u[;���wk]�&�$_]�B�L}-[���%��d���z�B�s�W��
�k%7:�;��j�*v�ܡ�y��i樷���@����;HKi����λҗ��ѫ��M�N�ӱ��Hoʜ*݋:��;V�)�X���<7fS��K*��1`�S]p���᧭����y��AZ��`�fc�&���3�e^��TI�	[%���}�{D=�%j�Y+H�ڗ3���P����
�Ր��+�l.���ȮC������ሚZ֪u�U�P�Ô�t��zf�E�(�L�oV���uʙf"��[�Y��LB�*�8[��Ly�f�y�nd�+�r\G���zq�\��W@��cTL`ǵ�iЋm-�x�b���.�{�������4109էy}��C|�����Жo�f�s.��\zr��R������*ӳS�.��Y�W2��X;��%N[�Db�SM�0m`�r���\�L�����-+<�z$YX��ۣ����#���ׇ�"Ybd�<�g�nUܺ�oh��C�UY�$9:w7�ޓ-j�r�ۭ�����9`�S#G�r��IY��=ט�L�pkΣ�+�%d�Z��5�6�����f�=�'L��j�*R�Umv�3m덗��*a��6A<�J���a��{+Ego����˕����5�tu��o�GpZ���q���5�N���C���.A̬p���e8��-�2�Vm�ZBA�T��8v�ę����,:�}���#z��:WA(�-��Ec0.0@K뭚���z�t��������Aw�?�� 
���������~�����_މ�?�>�'?_�g��b�e2$�KD�a9!���%�Pn!m�H���JNE	i��p�ԉ�#&!�HT���h���ꌧQ4�mҍ���HĎy4�E��B�UP��m���G pH�!E &C�d��NF��D�2$�6�m��dF�H�1E�e�A(�pG��FTT��"���J���z�m�$�č�R*]		:l�Tג�$�T���)*L���*�n*H���&�2&�eR3C��U"�>!$h�$L�$��nBH���,5�I-��E�$h��I(��8�&L���B�Θb$$�0[�/ �l4�!��(j9�+�#L�� �H�!ȓ!��`����%Jr��|Q(�jD��e	
����e}<�2hQQ��6pO&�i�P!-%��0$�*��2&�
Q��~(2�1�1�7Q6ЈH���)��� �R,�hƔ&d���.�p�A�a����x�P����Ð��J��H�)��#~�4/vv�)ч���;{2�]�o}�%����Ћ��4�]*��+(�x�vb��'�]�ۊ�ʔ�]�d��K�&v��պ�wVg9r���ԇ3kk-���F�kn�޹�-j`�r��_;ƆZȶӬ�4w�$��wr��WR��/n
Yچ�بmq�|�%%�\���U�TQp�̤����m@���2�OQ;�q��:�l�,��\���
Is�!��2Ϋ8�v�\��ش���]~9�nZ��SV,����˳]�6r]A�Pl�ψ�\)J-;g�u���s):�9H�60�^r�	����t�[��.�:>&7\�`L���z�7Q)}�]�h<��'r���cZ�1�˝J�WWj���X��Ѧ��=��Õ|���jd�2�J]���Z�{����G��k�A��˧\Q��U�P�Ba>Y�����̗q�[/��j��+�p5� );�L۝agS�XZ���r�D���Ű��:v�#|���
<�����oV=�9���4����m�����ED�,�d&B\ƈA���* �%��1��p@J��j�A@��
2C rH�2F��G�L�"	&#�i��n�D2�hI2���/2"1B��aD�?8�ƈd��.�p&�	F�P���*4Ӑ�`����0?\eED�
m4��0�م��6�D�⢌��%Fg�H,D�0�qrG�5<QR>LC	d���nZ�T��I�-Qd���8�	FZD8�CIA,B�`��Q�XR�-SV3�O3"A�$�<�m��a/4�/4�GQ��D�X�
z �p4H�(DiG@�*BLAFch8�H#��R�&皜\P��H �m��B9p�LD�Q `r#!�qBL�Q��&�IHRfDS�C�M�	(�Ԏ����J	��08 ��1\��r6� �Im�)F���Q��R9�RI���H	�	"Ϡ����H~A��A�,T��Tp9�HR"YD��@��m�`��4�QKIE (�R%�l9Gʌ"�����
1�"*B�P�Sa�"&�e�#rQ��$A	�'i��"1"!��(8([a3�B�����ɉ�"ny�&"#J8��K��#3��! m�,
z �p4J>�G��S�ȐqF�""m��%恑�#��Ti*��(�
m��$N1��m0�TY%E��N(�Q�����P�QP�a,�6���BD_�j�m�J�ό���@�"�Q&I���A |�Q��-�Ym�aN�f�m4�L�ɍ�2(���Q�S,F�Nm0�Q��2�F(Z>�(��q�A$�C~i6m�|H�&T*'��$a@�n@�~0��%�	���)
2��N"�EA�d�ߢe��A��H��BdD&�*$J%6�EhFn� ��L0Ȅ��^.6BO�d�\!$c� BE(BJ7愐�[�)$�,�h��&1
i�,y*" ��Ay�^��m/BH$�T�4@	�J>�ڥ���wg�^<W7׋�7���������ƍkZֵ�kF��k�����~��؋�q%�Sμr�x�9[ǟ��lW�������3�ddd3��]z|{|k�F��kZֵ�Zֵ�]u־>}-�WJ��}���ח��1c}���n���~�Ͻ^�L�@̙�x����ֽ��kZֵ�|hֵ�u�]u��o��H'��2�$N�?A��V��o�x�	+�O7������b��^��9<�Hp��c��OO����׶��kZֵ��ֵ��뮵���I�����W���$Z�P\�Zvu�3ζ�h� �k��sqB}y�E�s���U�u���"�^-���c���9�Ŷ��wwX��wV�<�]r�-ĵ����ߝ�N�5�滎�^�1���t4Vץ��:^��2W<y���B]wwr�<sj�7W'rڻ���.���ۗs�v���iy�V�:����ήw���G�5��E ����!�>h�l{���M���aH�^��FEd�fs���87#�	��!a��r�C�8:���`Q� 3կ}\8��מ;�r"�%<��� �}�@�%�X/B0�fsp��I�09"G�y#�7$��J��#HF���kĐ}hSG-�Omr�/��K"Y�߂ޑ=o<�5������J뎯<�IOm˙�|^BS�Ǘ���x�u��x�]뺗�qw�L�w�r�^C�<����	&�$o����L�j6����D�E�b%��cȖpI!�I��(B�D�)4	I��MB@0��l@����	$��A��"�^%0�HYr!@T1ׁ���L�Rβ�.z�LQ�����M_@f���V�Еk7RwrW�ܵr�s<u!&Izcm�&`�2c��*4AM�!�e4�I"	rI�KMA�(�j"�~f ��GH�4&H��&�m��L��(�M�T.8�"DC)�$MڊZ���M��Q��a
�(I,4�$BqO�QjFO���QA��$�N�6SH�C��Pt��
��p!!�!LDD��a�擘s��1��="wy7��͙sWjI�)�&�y���%X�3fԘUSQ--
���S ͷ�cͩ���9r�R�(U�}�'�>�gx�j>3��~������]j���ǐ���G�%z��jϯ���]�}� �{6����TY���p�/���SΏ5F���}#Eۉ����uib������Jst�3�^l��������或����ڍ�՗I�/[Jf�;�e4��>���d����G��C��=8��񃲠�Z��r���iL�6o�^�[$ٶ`�mH)b.�� �J��z���(�E��^�;"��ג�;���}Y��O-;�^�|��N�Q���q�gZ�"�)	_�V�e�eF��}�i�J�s~�N����}��l�^;�{�If�I�6�<j��AĞ����M�-����/�>�`���	�짗WH����!Y��߭�n?5b��EUҢu��e0�p;�V�u-cE�si��F�|0b*�bj���I��tѰ�QZ��}Ix��ܾ�+��Z�!����Q�y���&]G����r�u�t��ڌ�wl����S�¨xxxxxW����)�_Wgg�M?���܅f�~C�P/D+�;�?�;��3��N��Qz�:3�S^���X,"�7=,��oQ�M���Ƭ)�6��{wy��D���ٓ�03Fظ�Ժ��3�U5ܥ����}����:Qo��U>N�C>��q�%���Y��s=�b'#)�If��0��3�����U�y��ݕ>�N����Vʥ�R�#��_�R��+Sa�H�����}Rgض�0c�t*�f��A;�iA�Qp��3�|�{Q
�=�����������������xO|��{>L���i��s�}����?9EϾi�V��������ن�a�������{>�-ﹹ>��%M��.�}�ä�8�34��Vu@�߷k,�D
��2ﲒ9��|�6����Ӭ�?;�Q������(/���ZvVtWu��J�r�g+��i�n.��w��ڔ��m��{EV�y�wH{�#t&Id���z�(Ѯ�},�����;"m�'X��b'���^�}�+�G��}}%݂��������Y;w;�=X��@���4ac�?Hvv��z6���m��C*2ԣ����a� k�G���'Օ�D��I/%�`2Y�wi�(��I�ve������/�|�����}���ֳ
Ņ�j�9yZ��>�+m<�wgv|4�fyd{S0o!Q�ˊ9�S@���o2���t"�W��ϯ|�'lgS�A�gx�����g�&a6��X�5�p�C0y��X-�ϙ)'`ǣ�p�z��Q7>��f����A��W�=s�dE��~�m*��wC*���XXq�_Q��-1Cd��S�����G1x@��r�b(��S����P��y�H�7�Z�x7_w /B�o뉴;jܝ�wv�D��8��:� 5�9���IK�;�\:cdQ��}�����~�o��U}�,R���C焅&��PZ������M�M�,[���f��p��4d��n\�$���;���&k
V�Ǧ�mX��*�l��͔��Oz��7���J���0s�;���[|�g3�@>9o/5��ADP���LCcȲ�oQ6��u^��P�u��|�ۉ6���>�C!B��-O�#mno��i$�>>���kEzR��{OA�r��*��˕�i���v���p]�Q�;�U�C���0b��e��J�����Ek�:�n�$c}�˿Zjǌ�@����R�ǚ���>En5g�P����H��b�����*k�ly�ŋyX2|ǡ\�>��F~5��q��i��Q7S.�����zICI2٩� ���᾿[,��R�ݙ����oo/Qb������M��yν{��߈��2���j�3���܊}������Wط��xp�s��p4��t�%�-WVu8DS��̵�5��'�c/���.c7U�W��o�6H���E���Q���/�{}��\��Y�u�|n�#z��L��U������
ц��V\���(���C�I)�|�[Rw.T	�uf���tT���$�.L�p��jWr�M���@~~#����7�'G�ׯ-�в%\�Ĝ��L���r�Q巻��l�|x4u�ٌ$�hE{H��{'W˖\��؋���.%{K�h�PM���X@�����]
���z��φ�Yr.]��ň�V���|TP�^���+���U=R5��a-7a&����:��4����p[a�|�����ݭ���S��T��!�Ѽ'j�v�1S�E�L���
0h8���q���c,+B����jU�*�Z�u_/Os���9&���N��e^%}�HT> ��rv���ax�� 4*��,e��L����(�V���*�=Qҟ\0h5J:�E1�W8OZ��L-+0�ʄkYLI��8ދk��m	��R
 \�y@H��_�X�;����앺tIp�U �N�KCl�V�m�d ���.�����p���.�J���4�Cyx��$�ol�dz�4����9�^�E�xӐ.35�kyv��Y��7iEJN��5�z�KJ�A��XʵK �-E�R�g��s+�<�T���5�a!�q����7�b�t��P���D��=& ���r?'ȴ˷�u�m�$��F7q�S�+����xxxU5Qݓ��l�RW�l�@���vA��*q�hPt9��Gb�&�N��!� 4;,R ײ@�3:�dP���Q��x�	�ϲ)��^Zpb֛�%�d����;<N�1+P�=�Pꃊ^�ٖ��^�)[���{�-9t���e!w0��@@̥���v����h�.ZE�{��C/��9�v���N{����^RA�r�<�{z���ZR��a����<��Tʢ�|�Jw_3`l�����g�ԓ���hY7�g.���=^H�L��Fx-���u�Op�3D角7;�zQ�=(|����g|�x�UҢ)�m5���*�U5Y�I-P�m�B�5V`2!����4�� DݛN��c���ӻ�/w���}0;7�(��m��=7�/Dq
���wԹ*�����^Z'�aX��6K�e�o���+*����3KZ�-�צZvn5%�Hv����*���@�I3�x��[�J�\,��h3wۥ���3x��Բ"tƢ]{����S���+�+��5.rHx�1�H�_�y�7��yo��['9"��yO�ۓ�؎/��6
)W���LX�rVֻ�w�{,)Tf��|�w���t�di�HAG�xz�=��񋒦~�:�^�p�U?���yݫc�w��9�	��{w��uO�	%T�{r��a��"�rA�x��Y�0�>���j���Ko���t�;4�������9��s�8[��q"��}�G��~��/���d�1�m����e���eZ���R��H�8��aF�'��}��E�}�c��z��O�O=������yX���~>^_��ۊ�N��0M_m�6�3���N����i��|�E{�jp	��;vBm�	�Xl��,�.�O�%�1o��V=G�M�}������ �^Z��l���"�׃[�3q*2������\����c�P�����M����u�%>tg_w1J�e�RW��֞��Ӿ!ޫUQ��e+;�nTH���ut�icnn��x)kP�[|	ن��T6�������F��2m�7C��||||@> ������(}_Wo���c���Kg׫*$��m���L��ӻ&�Pe)e���牍y�^�Xhg����!+*����2�y�w�r�����u�'��G>|ކ�3闍M��L;�ö��,���7���׷5�_��(A�>�R7��L��i�w�5yU���3'w*�Q5��#�ن�&��-�����l�{H�b%-#���u�E��|���H8f�.��RX�yX��j.�"�<!�kT=���D<�3�58N�:��Wo�p4�=m�xV�i)�C]1u�|Z�p��)ރKyj[Y��Y�V:�7u&N	��B,-z�q�U�n�R�j��N�SW7����� 6_�y�ց�o2��.�eQ��\�q+�O��lɟC�B�&�輸V���9n�k��������j9sX�n�2��5B�iϵ��@��ԕ�>��1��:|�l6��R���y�iM%�c3fEO[*ƚ\�b�����')��5�Z�e <�����e�~����-�u{F�fų/.�PTK�
I��v��f�Y�;s��G ���tzRK�nQ�M�z��x���;�J;�^KOF��7(P(��U�
���݃;���C3ز�	6��}Dۭ��-j5�X�*��k�9k�k؀��B���x1��@�/3���4�ox\���)e��3�+J������=Sy�0��Iu�x7����7�81�Y¨�P+<�Z��(���ۻn���$�w{x�ό��XS8^���pUЧ��u��Xf�)��t\[�I˨iw��/}��=�6S���������b�Ỳ�-& d�@�1�|�=�h!~}B���]�!ਝzU{�Q/V���BV7�&w���w���W��=�;頯���(| -�y�sqI��H.�%٢&S�{t��}T]��n������gn�Vm�ՙ�p�x?_�4��o��
����Pǔ3Ǣ޵�p�FD>,Y�v���������IKFhF�[�6�t�Ψ�h�fċ������:�99\v�2��1�ʩ�n�oGv�L��eH��q�$�\��x-�<�CHG�5��%ӗ�o�Ϝ����x�c��fc���i��p�����#��>�wƯ��WW�E��70��c�D�?\3��Y��wg�Χ�1^���_�5��K��7�����3/&_�*���݄��}(�͕)%>m�ڧX}^�p�3��0�Ңv͒I�f"tޖ�D��r.>��n����X7�6}�73=�� �	ͿH����*��[��A�3,��4Z����T-��B�Ր@ȥ��99�IJ[�¨yU�RH��>Hg���B��Y^�>���Wת��P5m���l�&R����jU���u��}g��W�Մ�C���i8	�-x����zX̖}!�d���g�R�n�� �b�&=�����`��+���ή��=��%{�,}��?x{�����}��L�ʹ�S{��� �d�fu�]�u�֞�= ؁kv��j+<�;�y�������tX��6��g5\���+P<p�JD�̮�.�l?lD��7+RkXGT����uM<��@�V6e^�ڈ�Tm������i8�\�bμ��A�����2��������X��<�l����}fP6�9(M�z����k��Ucyn)F����$"�8{V��J�u�0��Z��\�a��+w��6�<o4�ﱪ�cN�|�Q䱐�z��Lx�F-��9d�\��+��v�z)���U����_[��Cݏ%|Q�`�d1	�i�*�K9�w](f���;��b�9�u�k7�����3�Q��bٕ��;���f��T�A\�>*�3�-Pr������q]m�}���4���BR#(�!�'%*��׹���h�&<�-�4��o���ڵ�1�����QAR�@�o%�>Ȋ�U�1���sP���@^���Q\�s�H���j��p�ޝC4.I��0��ɒ��!l����6���lR���f�:���7�]�WR��5@��/8\Am��i�y�U�^�[���%r���B�^d�\�Gn���Y�-�E�p�ʑ1�k���[ ��c�O�WM0�b4�oMR�5p&�ۡ(,iT��:��}��<�� t<�6����~���ua;'�af�*�f�N"�\P�}4�����I[0t#f��nؼ�N�D��-�k�ܑnh�M^E9j?]21M(B?Qۆ��ȫ.rf츒�����c�;��i��Ӈ:*16W��oAGq�M��%�S�sq�y��i:���7��s�A[Iˌ�1�_7D⛕����}tuK{Ŭ�Kl��]j髍��O���:�nX���8뻾����)7��"s�W14��W�:�	�'+/�rY֕�YK��S�9�9X�Н�L�״ym�9s�#��GpǇ]`��1O�h+U�<�a�Oz.�����V)�%�3�ۘ9@i�l\��u�4�Bvl�I]5$�-�]~��H���\��qǈ�,u������t�}�5��;ϣ�ͮť#��@��o!U�TI����X�XM�'z��V:�bξ9�-O���+l�ɋNYK�wx�l��#��r��,��*���u�c��ѽ�ٷjW�1"Y�t^�f�(� �kt꬈(��N�@e���K�,�RI�I%��ӼmD֙����̒�����J[�M�=���y �zp�^�^"}똄��p�4f�9����\����s@Ǯ������������������kZ־4kZ׏<k�㏞IBO2BL����G����#Qwr"M����q��H�H��zkZ���������ֵ�|hֵ�<x��ǰ�$�c�e&��$w
��yҭL��q+�e�i�~��~9�:��o������}}}}}}}k�F��x��ƾ�=���d	Na�BDG㯽�I�\�/6�sFo�оZ��5��&3s!�u׷������}}x���������5�kǏ5���ߑ$H�%%(��"�rgwR���44��h���뷬���s�Ͼ�$������x�h����Fƅ�_�$�]������T�����W��,����䑋)�M�G.�wu��<�E���0o*��{W�1#x�]��� �#ݹ�wL�twx������W�<��R$�.�� ��3��_�� ����	�����} �籞be�7��]��
�O�]�Z�&ڂG�b�d�Z�.���#:��>^��vy�pq��q�#q��vc+N#A <%C�ly��� Ud�O�*y\��[~��΄�X����-�={ЙqS5-��o��x-��*?)���T>�߱_�˚�ϼ��0G���h�p��/���g�=�� ;�G4�@x�=�%�x2�����u��	��
zhj|1�6��x&������әu���xx����8�Y_N����d��}�{kּ��^��q"g�@�+5[#9��{� *�[�E8���~��9W�~�|>�g)N'�f���,-נ1{��0����<�k�`�����+�+7;�  K�m��7�q�� s��L����Ơ{ѕ疨p-�zp<W�y�?�΃�wi�����J���x{ũ��8���y����4������oW����rF��z�ǶkY��F�/������y�)�P:[��%��S�W��(�_|�Հ�'»:Sx�({�Ζ��w\j3�����&�M��z���!�h��ֿw��_�y�WA`-�͞х�4�9Z�>�+%~�\���1�x�������������Ț�k�<3�4�g�ϹH�!���m_N���\	��C��8���#0��ւ����)N�v�5���;HtB�5٘pW��xQ�b��n]RWNd��)E���œ%��fyj�K5�mr�3��=ӎ��:lR������Y�]�I3Ŀ�}~C����1�#qĽu������T:���y���:>�G�4�x���ᬌ�f��6W����|�
����x=I>�w�>oxx&�4��r\[Zu��.-�dK���?�a�c�N/�L��`�����}�}��o�a0�%2��l�������g�����d�����`0g���`�m���o,�|����~t���cs/}3�t�@UχH���M����鐕�E���Jz1KS��O��������0��+<����ghA��"%z���1��ОV����]
�����~��k�n�қ�Zu{���o�-�� �I���z`q�*L���W�����S� �дVie�%�.�-����o =?_�M[���2_�dq��}�~�$��vE�+�/�3�_���ݙ=}�]�FE�;�=�y�����}a	T��`	q�dS,�ǅ��z�b�lxF��B��{o�w���)�7n��|����p7��� .4��F8	���f�@����a������2*j�X%�(w(���s1g.���`a�
�˼��0+�E��r���^� CG����]
i��TSN����=�֡n��N��`��Ky@����}��^����Vu	D�����ٷ�#��+!
z���E��-x��zFr��}�Vx��%��� �w>���s;5�j��2S[�3�<YX����c��n�g�5�#q��q����g;�OF��?}��8�޵U�*+q�3I�}z6�n)�[dl�N��2M�1+�=�"݌��աWVD5����W�t�fZ<&*����GX�Ά�χ����+� �Ha\>���ƻ�N��ˁ��Ba�~*,�x׆9�@8�����,�FJ��}��L2-�(�_~�@,��A�CW|��j,:|L��ǫ��7Jq^�i�����k�*[�{���'�֣�G?yN,���$p�4=����0�d���p~~c�O7��+��2l��u
�U����c�Z1����f�9��d/A��Ϯ��p?��0��Vs4>Y��y��\=�{C�4 &���^n�<7���j8	9c�������(^9�
	`�(�6)�1� ��Ź�������O��7=p[�¨oN��N�*K}n���m��/O^�1�4�)����
��������9�-����zC����!��f?���5*cɨ!Yo�/���AL�'>��`C>�!7�ߦ�9��~�l;1�)�5��K\��\W�G�Q��֋�>����� ���M�f�7�Ē'߹�=�N��~��oE8a�0:��ކf\�n5�ҘM�]��k���M�f���i��Q��#}C���#KH�F0���_�D"�>C�,!O�0����]>�z�&�Yn��VӦF�1U�[�2o\�V���UE�!�����c�{�7,V����k����]a�yMwC_t��M9��b��\��F�$v5�2�,���gp�ŪɁO������c�8F8�c�8ro�>w��}� �;��N-83�&��y�3n ��	^��_��!��3��L�WvQ����7�]?K� ��\��Ӯp��ߧރ����� |`�v�O(Y�M�SJ�zo.��{�7U5N���ق�|�p���z�#2��lO��!������7�!�Ꞻ�_�����k~��+��=M�l�t/[���xey�'�v�v��ݕr<�D	x��MX�S�{{�y(�ތ�D��Gdw�c1��z���O���a#��@|�>�F��o�<��V]�~�*OR�;��<�o={�gY�>�/���������}���&�{���V@��K�S��Y ᛼�=��{5;�g��� Ų�� �yn���_7���a*���G9ap:<.DBogN+*���Ƭ���]����c<ƅΆf��&�~a���b���ا6���K�o;�@��<�$]�\AW�J�����{��G���j����4���� ��=s��� l��=��Cs���l�Nj�m�n��z!����xE����u�cx�������sv�'���m���ٙ�SG���&�@�/��O\GiC��J��v�y���dlN�U��:»�����3��u�@ڱC�����玾�
��mr��6�e5�VN�c#���qNY��[V9�0�Rײ<��/g��ノ88�*���������GN���,ٞ�w�M��a������z$Lz@,u��~�ꌒ�u���)� �����[[�{�{���S�?�uT���-�0 �������D~@~1טԫ�?p��vYV��F�.�xN7�:O����z��������j�F��&��P� x;E�
ox
�֟\B{ЫlQ�;;����?�w�<�E_��V���E�T<�X����x��N��o�[�-�%�����R���nU�?�_+�~�^+-���,��3y�� ̋�oF<�ȹ��"���Te�>^����#� �Ѐi�?1i�i�dzDxF���9��@f&S6ܹ��Y����D��a�n}�Ɩ�p�b9��i(o|��l�^�i�����+M��%�G�����TOq^��V?������P�r�t�C}ѩ�y�\r>�����s�O���wu�ܕ��I��������3���<���{���-?�r ��~{�Y���m%Z��a���kFЛڽYڭ@�{�_|�޸Lm����u���s_8�ް��x�>]�f��ф���7�̈́�=}���I��oWj��b�(U[�}��d�t�cy���\��ëC�[���N��5��	�����N;Gy���V�� e��V:
Ix�{�K}Ҹ�5���)积v�����8ノ8��0>u��ow�P6jqp�8S��Sk&� ��uK�����L�������^���w���C߸ ˺����D"��:�r�2��-�l	�����XÕ���}n^�[��${����D��Xw����vN<�}�Bh�y��~�5.���إ~>}~v�9c�����wc^�.�r��ý�{S�cp���a���g��z<��
�
���������'�}�	����k0��뽾�C��q��,5���f?7q^���ӄFCY����~�u�؝��K�^�e�����x�O5W�zy �`����.-�����57��d�Ng8�eUh��<<<��ɗ�zw����O��kئ�Ϡ7��ѭ����z�3���ǯj���i�V��(�.��z���S[H���!�{��`}�;�}���&�c�C��=�[՛q0	�5c?f�V�����y�V��;X`�3y1gn�c<�[��b`&���]�T�j��p(�ږ�n���[���IǢ��[��=�^��x��q��@`'��&}�Xj�?c��0R��Y�m����¾�JO{l^j�|.�k�5�O��R'j�g��!��n���(����>}d���qkI�W-�	Y��ʜ�͓-��꠪oL�A�uv���ɘ��Ee>�j]��K��~����1��#pq�q�ں�xwZ�!�e����d�a����ۨ�r��ƍ=�[���n�u��r����+u�9��t�Ų"&v����_x{�D�*�@��~c�f�'�� 5��	�1'��}��	Vߐ;��WS�)p��{��ğY�3[ru��#oѬ$o\��RP�Ͳ�`[ �g���a@���k��AE�R�l����L8ey�>0v��h�?56 �hkz��n�@��r������	�n~_/�;�xx0a]�	q0}G����`=������܆�OV�Ҷ�\�ҍ͵<zû��什�6���-���	Y]�͟W�̉���y|(��ƶ��W���붼n��,���ux�/^l��o'�m
c=�=!��1�ð�/�רP�OO1�< ^U*���<��Y�dM�^�R'�y�(E^�H(<<3����T�A�3�q�E��s55_+噧�<5�p��
/,uͶ�g�y�V���8�}�˼�� z�9�ml�N�e�j�K/{�a`�SwvzE��ټ"�5�C3��\��}���O�D|?M�����K�%vZ{��R�;����(���fX�N���'����nT�k�g�ZKӻ�>��۩��֪�3Q���4fo��:�~<+OɳV}-j�I>���X]br���mSUy{e_�^'ݫ�sUd,m��`*��!�~��V4���vkK��y���j4��)��3{.>̕W*�v��]՛r������||������,q��Gz�o�����9��g��1����k�e�7nG��l	����צ�P<�y �Jk�J�oR<�-zm�7��{���A��;�ݺ�T�	�[��d��')KQ�σ8�=Gt����X�n�⮮�<5�������G�y�2��H�
���#Z�v�3����m�}�Ѻ�f3��pd�"��8�� ����[�"��W?�8|'�S�P000^��ь'�Os��f��▞ɝ���5����3ۅ��ͥٯ�O9�]�~��� �5𭯜�ԓ�o�pA��@pӪ~�`ދ���g�BW:Du����&sBV/qY�5�%\D���_U�ڸ%;B,k�kl�qY�f�/e��||,#�#�/��$+��b�7�����P�>�á�x��5�ȼTG��}���Ǧ�����;W�B�ו�_?&C g��[㟻��*rltS�vQ�u�Z�#�y-�Ng�C�f=�x�KU�;@��	�|�LR9�#ɦ��&y�6�;LŮ�̒{�����{��KxsP�Evſ��,��RĠ#��߻��T��@r	����0�v�UwD�6#8��'�U]i�]�(�y��Y�]rtRӱjV0r��"�0*�锑�󔎂�Pha0�A��/Aq"6}L}��6s%M��r	��a�ԉ۠e��5����.�Sn�L҆���I���|����q�c8�c�<�1�=�y�7����<s{Wˀ�+}J��麌J�7�B/�v���~�^�`���U�����=���NM�N��f�����!�ky�������/�����]T�
eIuSkt����d	՗`�s����p��ϭ����A¿X��P��@�����-;x�+�\�kwq���ݽ&��V�'��0��p���^�G�_�0f��Ge@��6�)o
a��B��r��7vy�r�Һj�I@y�h�V�$M�T�
��y�|-/�S�� "]h*���6�x�~t�oW���T�gP��錝a��ǳ�.�;qj�8��_5�~��30/
a�������1�\@c�>���(�����7�u=�k�*p.�#D�{okl+��l=� #v�3y<S8���"�v��\��Lf�)�_g {)־cg�zZD`�K���{Q��S�Pa������s���D0g�w��3�kOYmǃY4ދ�@	�7A�mg�iO!���˳�rO��O�
��o���������T-W�Ɗ�^����2"��=y����3�(]ܬ�I��+L9�����mOQ�kFм������J�9��A�kc�`?h�;��1����e��8D*NômE���ӯ Pq���U�MK���_,m'쫭�2ϝu���v퓝�L���8�x�C�1���q�x�8ǎqXAd@ѰEFƊ"H�z�S��q�f�<�N�z69�-���a|@e����
����|B/��7вB�Z�W�x��<�ν>� a|"����_�߳�|�4Q����|m& �@�z��yq�oO���܉�.i�ĸ*��6z�\OdW�?��FǔV�|(}��h �DQ?�G� P������*����v#�{M8���3]�Bo�<7=#��`q�Ϗ]˴=�d��[��z/l��w����x�6Vv��Y��� ��U1� S��`&Ƽ}[�K�_���/���_6���n�Gk{&6��Dܘ���=3�ކ����J�!؆�ݕ�o��n.Z=O�1�
��Ow�W�7�;q�����!����^�����z���c�|�+��oߗ��W9`)�sm^������F��o�&V���n�X�=�F��<���l- S?��[\���p��[rZs�˿I�l�@y;�'�����@��A'���˙x|RS�>~C�!i���~3�ೂؚ�^o <�)pLx��`&�{�H�03����|w�c���t��� �� A��xxx r͓n�~_~�6ɡ�mځ_��N�'q#���]mJ�d��N�%�qD]p����$7�}1�ہ��S�̅���Y�b��H���9��B$��c	֊�u[�]�Y5�����^����G���5&���@�=Q[8p��u}p�^Y����z��e)uq����c��mWed[�刏uF�:��Y��td�7L�̰��x�l.�(/�и����*i������4�5gO�U	Ze8�j���L��B �C�u�7�O7p��j�"]��J�1H�w<�[2[ܝZ���[]5�ƞ{tNWpX�&��<�%Ű�%��Rh<a❗�e��ЌN
eU�:��m��b��*�YS8\�	�ꡞ��RR���nr�su�;!|�4*�T�zQ�=6�j�sf�p�����Ⱦ��T�W��-|��%�"�{��q��(�O���I�#���#���_rm�u�ۊ��KV���e�sU���Z���x�׉&q��QAtt��UU\T�f�jP�o:F�N��Zx�`�ruP��F+��!�7h�1������))��_r��p�e*��«J�����t3��μ����x�\<��(����B�xP�9�������.;�1�r(0�����Y^ܣ��DU��K�@�H��f�����5�s�S�U������FK~M��8�5�nGK���JC��7e�R���*�@h��G����D8&�$�]/�ںB�}��q2�Q_,��7p�ڎ��^<w�e�*u1�v�N���Gu̫Hޓ�X��m����y�sweax�@ۧ%�2+y�f�h�j���j�BSBd����͋�SC�{o�)
��BlU��6]�y�}:kڒ��.�atv�a컈ݔ�ֵY��Q�d��Ē�ga���%�ѝ�0Ջ�9�M���SZ�%�Z�5���aI�������r*��{h���4q��C�:0V��7��V���$:�Y���d+[���"�G���}&Q0hn����C��i��,(Q���l�Ϧ�C�]*X.ϞU����K,��`�)��n,��t�X�s҆wrrJ��D�n�2��&d�Df�m�h���������b�\z��ޕE�è�3@�B��ә7����,`�]
Xǩ
� ��Së�vRsP�W�r���r��fY�)ѦDYe�-����xWY����pJC�c�W8�	7N�u�yn��p�'��q�J͂)�4��JD�}��&o)$�ܒfV�sq�*ٌ���ul�*�/N�����^܏nO;ח��a�7�ӻt0#�����CM�}�w���ƿָ־������>����x���o�����d�q � �F1��˲��7o7�������k�kZ�������>��������߻�������+� ��(�g�v~���,%��!#$$ Bzx�zk��_�k\kZֵ�o���}}}u�Ǐ���� I�\у����k��\�D,��)!	<Ǯ G���?���ֵƵ�kZ�ֱ������Ǐ�O�~I�`+睼�
Wwb�2�JID�sEZE󺧾�LH���	����'��>�D��{�y�X�%)�!�SӲ\�O�c�W-)��f?{\RC$���p��1��f$���&�]�h���恒�D dh���L�Nl�����z�L�	'���u�[���߯e������qȉ1�D�GB�	7�S
)(�'���i�I�$�	����j��A)��$Xi4[%ĢP�QA#b��DK~E�m�ٌ�ICpniq;�+)�����7�� ��X��RʛX�1��L8&̶�J_n@��tO���F� KE�	0���6�B��)O�N�R&��!H�Am�c!6�@��B*4�A����"& A�^18@p�'Ŵ$M�)0[aB�
2Za	y�B"�'2	��K�4�M�-4�4����IH��N4Z.�,��p��,�A���Y��f"���S����E�ʅ�[� �A��!��3����y8�<@1�<C�1��9 	$@ �x ���O�M��J�s��F�푶�G;�5$9�DQm�ɽ��@��ঽcyvjqIc波cx�{���{˯3o������_Zd=��	�
�z|0���u���o����>�u�,�m,��Gaͤ{��3ML�� �-"��!۞��)�6�dKxN����^���Z;;Ǒ�=[����{�o ���&s�d��"�N�u�ֵ���H\+}�q>ǂ�Kkb��5��s7���X�3��e�3G�����ݻ�zt?��LL.z��_:�dz+��eC���5y������������Mv�ӎޑ�9�I�0M�9�}�6E��r��M@����3w��������y�K}����@A���
mx��\S;^��7�����z�d�grƙ��p8C�z`�ᝂ���������|���������_^��
����c>ؤ과����7\�������4�6Z�Bփ8؟������_�h�����F{�Q�=2�!�U;;ć�n�b��煰��P���诿1����3�r��樗�hGow��b�8���/�N�5݀ufm�!���^����,:�.i3�!����_�HnP����nf�7�!31)�W�ڜ��Nz~O.��]�
r@	6�P!��o����QW�l�u�|���t�Q)�q`Ym��1�牎�:j'�Uk�[87[]�]t0�4�A&�� �����yd�1��NDI�1��1��^@D�d@	0���0�L(�z�G�9���X<dW=�ŗ�=z-�a8��(�a��b��y����u]ț%��ˌcF(-��7}�^F��2΁�#8\
�mvj`87��^QڶO#pn]m���G�0�E�$(���_��g�g�u�k���Γ�j��x��O���v`�deW-~e�]n#��zXo����zC0��.�T�n������>ln�	V�HQl�sC۬�G���(���<��3��L>�v�k&}���y\�ѐ+��[ɾm��Λ[��KH����W>�3��I(jEL [>�g���U����@�0��G;�4��=P@`�����m#�q�FLu����3�F�c��������`p��|���f�;s����L ̹�9���{8�L�{�ɭ��~d�A�	ߕ����B
-/�/�q{���8�����a�zֳ3=hB=�X���*S<�W�}C�@W|��;�@O�a�O��W��$�?�_�c��<�O^��y�	�v�w�~��� 	�����^>F{ �+�#|`͟@��,x	�(�u�uN���=���o���<f�|��ty��B8;8>��:J�x�!t:sU�h�[CN��҂RӺ�J�|���z�K�̓�X�;���@UBIK"0�=��d�9R�t�jϓ�E��X�*Ks&b�&s}w��R�����r��>�'�����}x(c�<x ��<x� � �7f�y��6�Z[XڋV���0J�{���t��>T���,���'<�r'�z�J�.Eל/>o��h`6&�'���z��\tpN���`Y�r��T ,�1f�����4s߭�_�G��@�����7���p�~ݾC4.�{��c9v��̔_� ?$�ϩO����Ѽ�ݻ��]�nq����Sr�Ѻ�<�g]}]�5��P/l��Ow�l��S�i��[3Xqۘ�U6���	ؙ�-�E���끭����xxA�yL�m�;���t0S��AfH�F=�5�1�4U�_epp\W���W�����/����؛��>�藖\�s�[����ڍ،�]9��N�òkmǙ�h����Oʽ ):޿Vs�,qb��t��yvvF��Xp��_؄/�����	o����>��z�=^Q��2���"��j[�k\�}�'�^�Y*�M��l]f�������m~�D���G����6�����ß�/��-�܁����pb�<<�up8�q�D�O�ӽ��l�����f���p�7���(�b�}�ω4�s4�^*F�UrI���݀{���V�*g��O��}b�[uݚ��i�N̷�P}I=ƶr���|O�m��eϯ-�ɝ��	�%lRv��Q
۾NlD�S6�����]��Z��"7�l��cѷ�:37lA�q�o9x�<F@�D8�<�D8�<�TH�VA7�ߝ�����>���縯ҽg���5��`�!��@���K��O	ʁ������q��w�}��p!�]C����v��]��|���l��&�M`[ d;��i�Ҷ�@z��ۗ��1�a���f�@�����������4�����$�_�F��S�~���7���i<��0�7PMr_�M?��!pYۙ0������c���k�l1��uq�q;W����� �����h�ˎ�g�B��+@ 3�~[���i���$��8��Y#���D�εڸ,P�n�|�7�1.;odNZ���x��q�#���������]��BʽZw�l30gf���>q���߼N?���0H�0O4�s��ß��Tbл����N�n%�zCS�D�W{d�F�n����.�iW�(�{l񝀩V�5��owU���4Æ�=.½\��?��#ڞ!m�>>x��>����V����_o��]�\�[eD����3�v�%�ʁ�TyM����[��.�p����C��8��@���I��,MRbn�C���cu�j�w;|��yu�"Y��~���)M�oj�%h�k�ځ��z�Q{��	A��6׼ς k�aħAC��w{/�}-��̻��z�[��Y5�u�4#���Y�Df]��oa��2XȲ�4���?��y����q� <cǀ�<cǂ�����k�Պ�+J�U��o���w���R�x��Ai(Y�eb��'�y��ĕv���ؖM*��f�(�|�=���fk}�Kv�Q*�m(�HU*�c���e��^�X����گ����������k½�|���u�2�:=��~ut Z�sv�qu�(�&���o�xs�#i�_���,Â|`9�a��0���F����d�N�ˊ�	�����ss�������^�]�=���"�����>�xm�@���4�<�.��|��`Kx���g#�	܎�O�l�Z��'�0�yw������̥��/�����}$8|9N���2�2+�y�a c�r���������__�~k�$���l�!"E 0��c�����y�~����Qח�z��a�a
��z �48tپX"�(���x}k��^;��;ԅjS�5���L���]r��x��)���W�`� �A���f��Mݭ�������\��8k��F��֮�4M���N'��<@>=�r^>�T��k�����"�c�!S	�=��f:�'N���X�ol��<�I��	�9@zp
{��p M�kˎ�b���O�$s��!�� �����(�5���d�]W����$����@��m	���t���k�wvz�0�����;&�o=y�}���f�.i�}����T١��nq4
m��QҶ�TO'�+h��?�B/�/�܆����>�j���k�D��0��=�����(����j�rɭc56�<���K�'N'�Z�1B�#x�3z�l�{W9�L
?���?�x�  q�<xr �q�
�*�q�<�� Ȉȋ"� �H�Ȉ>s�u�}������y��zo
�8�/�M#C:�67w�l[�/��.."DGE�A�E臨|O���Sz(?y3��\l�9k�O�� l�x� 1?d�v�b\Pʺ��(\it���)7�y�v$���R���"q�����|���1Bn|%������\.�z=F�w{��`&��݈�/���i�V�Ǧ�V���f���+ ?�� ���TXt�u�����h��]gp5��,uƲ; O����J�����X[l�͇��!�U�y���C�����	th�`�Ws�A<�k��j��0�Fp���48�M�{���<�%�Pr����Jp�����}����)�t_�u��3�o�����j �>�
"�֮�o	�M�k'}W�ٛY��z�t���1��0�}��Mz�Ј���w�c���ش�`o�Vs�9�J���H����ϩݺ���I�yާ�@�Sy�X��|g`n���]A��.(�rr$!�u�NWi([&���K���]�`�1�� ~X9݀f�K	��徦
��C��`���9;2�͂��/��0�y.v���[�
�w��2�)~�{�͓�W���q���$�7e.m�I��2�h���7(���҅vR���ϗ|�.�|��`!��><y8ǏD8�<@y8Ǐ 7�����j����֦js���p%�3\���,����21���������'��%����Rۇ�?�	0s�s3��類�_��E:^���L����˹xg�C9�>_ފ��Pp�F���ytm�'��[�����E5g8Y��!��y<C�@e��}.���	�/�k�� <_+��\�e�4&�otل���`����P�t�Ԍ���@Ϛ3���{�e�����G���)����X^ ����¿{�����~m2Tdo���+�?�߈v���p� *sRÛ�J�Un�<��޾�-�͋a�<=���q֥Ӣ��x��P�@o�?����3y��Yh��ܒ�K��3��kF�z ��r�o����X��3?�H�L����Hx�i���6�pM�n�9`0��r��`��>r%G���Q_���@^��B�F�+�B�<CD�x[��m���z�r���-���ȶ�\��ы.�0	�=O�� ?���'�n�wwW0��n���k�L4<�%�ѫ�i��z�q>���y�@��U��S�~ob������:6|�}��S���̥���ٟ_mW,1���:��T�/GZڳ���r��[0Z��D7� ձ� h����[�*���b�jE|�l& �̽�{�+랏�u�|�i;P,���$ӊm\z$���coD��3?��z������  � ��<x ��* !���������$"��s���w߷�;\��?'>f�����n���װH��@4s����Ʌ�I��ϭ�c/��u7j;M�G�����Ӟ��m~~�H6���W���a����ߪ`����@��,�F3���.���s�����~H�1������z�	z��!<�q>hoO�������ۑ �,�����<s
�<�k.��8��f�Z�zo["���"U��Umzm�{_��_\���Sa9;לNi@z�f/��6߅(��
FHh�Zuc[���vi�Li��n��<��B���=�z o�#�y,[�5K�|���I��� �&���F��-{��o��u\I�=>�wo3�9���+�0���j�`ӷ~�`/��wPϵ�o	�e��>͈��c�^���&�G��N�A��u�)� p)�=�$KA [�ٓs;D��=��τT�:���'w����ÆlxP���n5{v7)+}=@~���[����1K&Ln�`z�qKwRm�<l��x��i��F��zo�$�M��p(Ǣ��� ��, |U����t�'�r��A��n�S(|�q���}!�K�x��ݹ�^w�Jǘ��(�������C����;6.�Ö]cnKHnWS1�:1�[*j��1��Ĳ�j������h�C�^��D��x���*<cǂ�*Ȁq�<xȠ2� 
H��%<~g}{Χ&�|��Q'�O�{����(�NQ�w�ř�B����	��T���ynE�MU{J�-�meEm������3���t �-�`H�0+�'[�n���|��RQ?�� ����H����Wy�<y���)�!)a!��{ ^J
��B��	���������'�ϲ1��E�{n��P�2����v� O����|�&�Z9��Ɯ}N�E��;�h7����N�R��2�g�½��./�sϨ1��������4"�Უ�z ������5�;�	$��v"LT�(��A>¸|�%�ӈ����򠗬�1�5����������v��2��qwǰ�o����U�-�/G#wςi�瑨�~q��w�EU����4�2�1i*Ip��w��Y�z�nJ Lj�Ez�<n?7��nmJ �p)�3����ƶ�X���P�A���d����{1����oc(x��)�� /� V �Ί��m@�yw�m�/�Q\����RD�ӈxfx�������ޏK��\������+���kx��ʵ{��0�l��/O/����k��{������<���	��������b��)�6L��߸���7�+���p]��U�T�_�����pτ�^��h�v����a�U�u��N�6ͱ�b8���֓)�g������Ӓ�J�|�d�fWM��7�ț˻3����'[�JsJ�)
�zB�l��Sz���؊�8Ƿ�� ����"��cǊ��+����
"� "	�H��o�z��߾��H��{V�(�z}�ƽ�~C_�Aaا�E������?1^�~��qj�k�Id�^��E�����34�̻c�8��k�M��]�q��s�럯1�hQ����ύ*!��)��^��x���{�F ?r��������v��ԛ�o33�5kjhf�\r������"�jP	ח���: �]��b�C��+ໟ��׮�܅@���䌑��\�^��zb8 �@"}�,����?�s�����W��u���AV��ǜ�dvS�:�*+`3 �8oU)�ÁO����{ 4^���}u?E�|��<�b5ݙ噚w�1��cZ�ÂY8�}� � �a��P�����6�g�,�z8���n�挭U�x�0���p2��B�8�k[ש��{���
oH�a�� s�?��|e��K�̷�}�u�������߶< ��ϽIW�>x�/(�;�0��z1��3;1����X{b1���@\*F������S漰�l6��V��j1e��6�	����7��m�P�yc0,)�͸��9��t#ˤ�̒>�U�C�`	Ho��d��֥�r�h�j]	9֎#���鳒Y��x1�ŬF��EܺWNj��V�pTK�m_8�.�n�㽩Y9��δj^�@ղ�۷Iј�;1��w3�gs���Vm�]���&�I)-cҍu��}7:��%v3(�s�|7$T��{�v�irPdl��D��.��K��,!|���՝K1�c*Y�xY}hS�������pu�U��>ۆ����d*-b:-{'sw�+luP���WE n�;�C"+.��R�w���aC�>��SK��4л]�	o�j���ڑ����n��D��dU�D0��l{��e�QO�\W�0t��v�v��u5V1ǒsX���
���rU��E�4����X�Z��]l'ۥ����B'��"*��k����.�D�n�+�����鬳Λ�յش�C��<V�"�Ln���pfM�<x�r�!t�ǋ�ԛn�K�ۯ-݋�k��)mΎ�Mab�{�d��Fi=����X�o�(���֚D�
�h�ѸR$�����YCy7Q�-�R��n�)-Ua�>�xߕ4ڪ����	X�3OG~�	�;�Jͳ�X�w1�(�+�A�+��������|[I����"	h�&Ę�Rb1��@�y�� @:E n�I@����3���k뙝',������kYm�%�����h�R�
��SZ������ϱK(����/ �T�$��'N��W%)�-d�HC�v�q�L�R�̸��\fr�5-����w�V���!���J뇫mm�<�v�*wG�#�Zw���J��ג��+���}	�r�a��.��]k莱���Ȱ���j�#Snp���ys�5q���1|9P�ޱ+dt	�ܧ��wz��_���8C+qm�$�0�{3���,Ө�C��R�f�v���"()ovp�u��u*�+��m
���*��Uq����|e"�T�$@���eҧ�Oh����lJ2��<���9D��v$�r�:�Z�F�w	zx�Ǎ����i�ۂ������������U�p�Q��'*�.=��MN�b����� ��앜k]Va�7����a8��c�J�d���h�Q��Jjթ�m�͸k��x7Z1U�>�j�ڒ���t>wD�Z�]ʖ��IN�^�K�Y�Z�^�Ni�2�Y���C��ͣ�fHY4��~��DH8|�J$���w^��^��@�#	0G	�20���5���ֵ�k^5�kZ�kXֵ���]���}�Ϸ$$��f�y�v�������?���vHw�B0�q����zkZ׍kZֿָ־�=:����������~.I0��\�$�$d��$��ƽ=5�}k�ZּkZֵ�ֵƵ����_^���}��O����u<���/��$%�q�t��f%C�]�ǧ�����ֵ�xֵ�k�k�k��N�����HFB@�"
�$�a}t ���&E	&�������Q+����ݾy�LR6$��C�t	CQ�4��b�I˖cj��ƻG7l�^������TL� /��1&�)0X�AK��/%�'�t���Q�#1�DS�f9���Db�1����)b��t��@uE@���d��+���:\J�y�37��JI^³��˾E��o>����8o:�{�L���ۼO�@�k�Aǌx�1�<Uq��' H ��(��~w�~}�Ϸ���I	I��4� ����/���5�}���s�8��~�R�Ƶu;xU֑����n�r�Q~�$��ޖ^��f�O}<>?ẍ́8��G����!U��un7f��S�h��K/k�8zȆ�{� H��zy
��1���;^��A�]qv/�4撕�w_�<�{�}0�ׁ��/�2���W�yos<3����m�W�eN;��&�g�{�m��>$H?B>?�-��������נ��Ě�/||�J��9��a�sx)�ta�tss���vl�b��P⿞��f"{�w~xg �1���z����St�ܿK�>�	��N������<<N/���i�~��"�2Ƕ�������tX�W}9�PVP���H���7^[:y���y���9���8^����%��-,��g��AlԄ�l`	��۹�(�y���*
��{���+�`b�jj�Xt���hp.�c�x9�R)��/6��E��hY���ݤ�7��b�>�>oF7��#��>D�_ێ~i��~04`s��2�ؚ�u�n"��5m=���u���2��y!�j���bm�t-.G|l�VkN�O(q��;s��N��Μ��:�c�pvh������6��\U�Csa6�R��a�R-�\�X(���m���Ƴ��M���*&��7�?�H��@$E��Ƹ�E#ǎ<P8(ECx���8�Ey  ��dT$��y��=���o�b��?�\h����įvP�����xi��>�0SmC�Ke��-��uG{��'z�n6� ��cu�A�,|ɣ����'���Y���~��_���V���o��D~I�HM1̌��?4ԏ���֊����n=a=67��j}=�]�\�^`��8˪���.��l*6z1��p���[yۛ����v�Q�矛<|�r�|��CN3�2s�;����O�����ѱl���@��@Lq���&99{��OEm�b�$��@g���۞��f�^���X��y��r��w6�[�ZI|��jWvªZ�t�v��"�G��Ry��t�P�ܫ��~�~"���c�O��6�|B�����V�B�SV:�λ�D�io����%�{_�|��_)���^�|$.`���>��=O.���P��"�>[G��|�,r��[��^������ȵޛn��UxhlO���N�ڪ<7|����hX�".��\��s��f��ge�s�}.��"�z���6�O���EzE�a����>����gGԬo\t�\��|�u[9�:���R�TK5���H�V�J:�a��B	T���Mk��U�74?�og��lZ�ܳ�^�QqVR�����i�EIwר�:6r���ǝ� ����/W*� �x��(c�x�Ǐx��	"!"� �� O��7��*�)	���l���Z�L�OhZ8�Q�̜���a<ܝn��N��iL�]�!ꝚZ�:i�k6����G�ɬ��=���yz�	+jam��~(4���C��c�$�ü����� �gɭ<56��$6]�@��ǒ�i�k:����68k{�C4��|կl��+�� O�H��y3��(��U��+�g[��v
Y����mw������u��~ބ��zg->����U��gBB�~vx�<���j`�s8���{�ݏ,�@��|�ɘ��Ú�P*�)���:�"���a��F�lӜ��y���:L<�h��1 D���E����Ϝ$	��'�<[�Ow|�� ��)ʯ/��f�y�Ǟ���9����ٌ�@��#�[�v\cF>� [���U
��)�ݪ~=*֣����G��SǪ#��������h�P��D�a�����V;���2�s&�'�|�Db�nF�},0����w��G�x��������; _���2^����^X��`��>%��z��>�g�~��w�i���Vz��b������魎����o"�_�y�"�pO�|ǟs�A�*X�M;i��;=��,}�����~dӮ��`1���-瑻�S��y|�K>���,E^���w�����%,�[��kv���έ�]	Spk�E�J#.��۵�7T���31�r�FȆ�y[� 3c�f���� ��M��7'�RcN��6��}Z��Kt������l���}�n΃eJ�=����BP�3������/q^Dx��<x��Ex��G�@"����ߗ���}���;�m��D/7�"f�c����s�^{���P_^r-0��5C����)fN7,�q�N�<7���G�p0i�� �B�P=5�Zo#��@��os+��P1�t^;\�p�tsc�I�gH��-�YC0DM]̻0n}
f���4y���~~NK��������a�nU���}Ù���{:���{������<��@��?����Κblk�߄牌�{X���Oc.7�ukItɥ*�f +�E�PX? ¯I����������G9_ja�/��5��uً�����[=��Ĥ��-q��[��f��������r6��m:�ђ���0G���K���z\^�!C�4��� 0�7��	ں�;�u�����g�?{���<���[��js�>B��5�cMFU�g���}7���3�?q�\>z�8�L=z1�z%54ގt�!�4	��̸�U4���Zx�����㉹���5{`3:*(G'��D��ύ�l���t<p6\)L.E����"�K�?,Gw�MgX9�mn�io��y��wFo4P�,1�gh���=Y�V����lM��P^$����EZaY�fD�wf�/V�y'G������9 1ǎ<D#ǎ<@��8��I O�� {�k�;z�o���H*�T��Z(���b�Y����zG�jI�z�!��{^xM ރ.b�)=pD߱�P�uv�xKp�,#�X�vR1�r
�F�2�Q�E�u6މm���ҵ,�8�g��K:[�9mL)<��l܌	��w%B�ŗ���kxa>��\%_0�j�<�z��o�6�@���Cy�LF�����E77��09�w�m#8]r,(o\����'"a���/�Rvin���ر.�a
�k�����1d�Oe��XD�[w�d�X�pp�ވ|��i��As� �~"��3���=q ��k�V�k�5����ŗ��s�������~Vt�ySV"�1?0��	�� q��'�kx����zߛ� ���}�X�qP��t�2��E��^�Ϯ�  Ť��y�|ůf�M�\�x��4C���l[��1�ߧ��� �u���/X��1�s�[J��2���Y�QXpw�}�`5��<�r(�a���D�T�|_pA�B�!�������ܗ�A�M�[��M�t)�7��J���܍sa"$��s�J_{����Y"��}>�<q��7�zϻB���k�����9�]ǽ�
�a���j�l���9�ҋ�XNt��<������Fs��ز*~�5Ǌ���
Ǐx�G�x��"������|��~�}���p������C���.<��ע����
p%�@8��ހ�F�f�J��vc֛f3n�����/`S�]ld<_��#��Lz*�ۼ�ܞۙﶶ�==�����<_M��9e�f]�#��͜�y<�q�`�TVdp?��U?|�. �5;���Ùˎ-G{ܞ��
�f�n�xְ��n�LS=聍��3�v����ƺԜm��{6��Ň:7�Cy�C���'�f�y�+��1��`=[�H��h�e����V��>����5t@잟k@���"}N����	�g�Wl]�k�?;��
�5���Գ4��Ȗ�D�������~�\̶>9k�ї���t���AQm�;���Ŝ�w��'38����վqF���@P,�&���0h��Q��<��W�Z*����j9wkN�E��m]5p��}�h:=ȋ�d�`&��@*#��>Pj�וeu�D�k�zNk�;r��m)��֯'�@�ah@���w�?����Ru§���@\,�L+����9��LY�*���Nfێ���k��y��9[������gD*�̪�'K� �C�_/u$��0J�}��	����R;ĉ�]qw/B���.�m��euq�J�ޓ^[���Y�Cd���}q�����
Ǐx�Ȳ�<q��BH ��� �Iƶ��ΓW�d\m��F��4٫jM��{��ܵ��j��6�e�2޽�UR��̲�m34��Yӛwc��Dod;oL��INw�|C?�;���ߙuݾ��g��ϧ����]��-��^=�/m~�)]7ΕGՙ��B-n�۝3�jg������|����Hb�~5YL@�|pWe�e�����pK��?�Ɍ�4���PV{�g����h7���pn��=T	�u��]Ŭ�0����"�������������n���f|��Z��P(7}�O���8��{����8�������LШ�4/���-?�R��.Y�t�_J(Ѭ�z�]?^�>�,ŲY�X��>�E1�'�kM��?��R���~x��T�۳��'�y����3�|�V��9��O�o�,��l.,߾�����>�JV�7Ic� �v�E2ź3�`7���,Y0��m=����{�����V�T�BZfa� O{��=��Lzdt[��q��q�>�R1���:/:�7Q�觌~�;3�)��	��0���쑹�R���ɯ{e����P9��"��u�xe�4��R9՛���ܺѾU�H�c7HF?;����W�������W�ӷ4l���n��v�J�n�S�ä<�HȳOYĚ.�X��QMӻ*v���O��)��� #ǎ<V<x�Yx��N@�RD޻���y}���M�xo�cu���������.9�;y��o�ƈ~p9�k^��ՁW3jW&nGP����o�������h*Ҷ��=�~�q�7G�ȸr.��":��f�J�鲳Vi����i����:j�6�@ �Eu�kfkL�IF'��������!�l�1Ι��s�7^El�r��|�Ϩ(��^F�3M^j.`E��!'�33��p���9"�@Ƒ��.�ϔ�ێ�Up��%�^e��3��%��gSetF��J���cr}c1 ��P��,��k�\Mdb񇰮|��Wʛ9���M��יJ�F"%���G�q!��~A~8Ez���E�]�m�-H����a�/�	�&y�f���Gz;fm�(�u����k�0g�^g����5��y=�_�˸>M|��_}G�n�N��w�E���\��yŢg[z9�j�X!��1��qE�?A�|����#Z�/CM���f ���QR$c�?-�O���v���g�L�|�~�8D���������-�z��]m���Oʞ|��˭еa@�Fg;:��|���fs���ߢЗ�:�/��J��_A���ӌ����K��M)��(����!vilwY�����ߗ�_��/}ݚ��O�8�<x�Ñq�@$Lq��T�$ď}��}k'�~|�1������_��9����Q狵ܳ1�3~e��c	��o�Ϗd�|QIf�>$�����������^lE��qq�����	�I�.nYb*&$�Ꝝ[�f}}lxdgh/&D����<�ݪ!�eJ,~_�?)�A��W�����םS�$pkw�WM?�{���2k����P�@�ߍ0<HT�|B�<��8@^;]�8�eP˜�9�����hx")��r�T)�ܹ�D�߻��+-W�ydQ��d�� ��~S*��ClJ�V���x��� ߞ]�[K�����]��;�W5�EVW�����Aa��g髕�����N;�4z_�M8}]<���-Ҍ�=s�rT(<{fɉ�����g�+__4Ǧ�x��>m���L��g/�>����yn����%�B��籇dmu�������D�<SD	���_��7�b!�qpV\���q�_�����(����E^�8z�8�a<��b���j~��"/Ϛ��������W폾`~L���Gd6V��]0e���7'[C9tƏ4R//冭�����7`�yMWËދ+k[��u��xlmcx*��/�,k�I�j�U�' �ͣ*�tƋ͎���X�4c��%��tJ��Q��y1�&����������<<x��yq���q�=�;}�N,�{|��|��HOm�1^z��`̭�����s�r�o�c�_��OQ�չ���d��8�qoAO^/�P��yw��e^��W@���x��8�bs�l��<ev�<Ff3�~�~�Օ	���#(5BOZ��e ��?�y�w����r�/ ��ʺ�y���KZ��KW��h�w�����P��'�'𱀸�r�ghwn�T��p�}�{����/�*�&E�g�ϲ��ן�	���GJ���>%3p��?;�"���\�AbA�� �{��|��[�P�<�.6M�me��VF�Y�,�w[O�q;�1Kus}������Ζ0n;k*��"���w_,��&
J�vJ�1��^%�,��? b=�:W�,�3~�
��gU���ئt[W�t&{6�O�$�a��ff�L���Ϯ{����n4�`�9�֠_=bYW�#�X՟F��e><9�,e�nZt0�^��"������ߔ�g}��~�������	�sz�E����{����ˋ4��_;a'+���ӧF��VR)s>�)v�Ef����2#���d�%v�+�<��$\��9,��OU�n^�ʢ�_H��l*C�p�g9�����_t���E�:���$FA ���	G��g��:�a�-���M�̖�NX���	W���w&�F*Щp�����Sܺ�ic�؈𫝲룫t��ȃVO�N��L���w��ooQ�v��ɺ�U�y�T'�\ȵ��,%�*nʙ}���lBۛ��E�ɸe�sy����&��I���`�(��U�VS�u���2��E���o��Ie����p���=z�-Y��4m��<et�B��h��P�r��:Em�]+K�˙������(PA�'���fsv\<n�i	d��4.�έ.W�ŶK�\��G�*�!J�⋰�(�U�<�Q��B<��ش�q�xM-����X��IwcTf�겭����=��ƟS��|�V��m�A�<�P%�ևQ7�.zj��r��4t+�=�5;5J�O��J�9|df�ʗ"��m���@c�?��b{���'��H�V���b�~jP!4
S")�U�[P�~E���}$	�ܲ��P�/cߡ�JlJ�dvv�
Р�lOv�n�W	�}-�g���2���_$�����P�s~��D������=���z�+�Q�Gj�/�bn��Ӵ��Ք��E{���%]��N	M7�0��t.��,�`��{���^�sдHq[έ&\R��s2���HGfR�%c�"�gG�Ͱ�:�{ۉ��`J��Z��h<����v���T�fv�zQ�A�;.Q�Vƨ��e赕}܍1�:'8%�+"W[�uy��#�[�sc9b,I�x�>«l.������:��J�!��wi�;-���Ul����v
S��5��-��ڽY��Dz�ޜ�Vgi�y�ik(�z*���R s�hGx��	1�������u+�N�v�<�Mw[��u��k���Vl�<*3W�"/D�����֩�fhYz;R�����%���=}�r���(�tya}�yg
C^��0����B�6m���;zds3��YU֖�w.��Z U����J�/ R9�#�m�ٲ��MN�Y���l�]ٓy����f��ݮ�KF�Q�B�̒ �(+��7��2����tlLҡ�9��o�e�}^�_={���x� )��(1Бhs��w���^���Zֵ�Zֵ�Ƶ�5��^�u��ǿII�&D�ⲗ���{�Dli��������kZ�Zֵ�MkZ񮾽=:�����fd�d'�6�1)�%��F�F8�����ֵֺ�u�kZ�ֵ����ӯ��>yBI$�����A�I�:�ę�ہ6���#Ǎk��_]kZֵֺ�zkZ׍u�ק_^>>����dDm5�!��|���ݽ.j~g��uf4&a���)�,�~:�(�Hjؠ,&CA	��DT�:�BF�����QГ��]���%�,���&�K3s���tGu����|�Ġ9����32!�"&%���ܽ9�;����
aQd�4ޝ+��+�ϟ{Ӽ�S��1��	�����J�qD�0���ec��"�h�b4�h�, �F�-&Q(EL�b���ų,��R�3$�!.�(B�ܵ�3�<��d ���[����\��vꢭͣj�ֱӬ=��՜�Kq�v��JABA�"H�	r �&!��n�BHQ�	�2S��!�LQ�ЌE���A�D�*�(0���Qs���I�"n*7<�fI��6�)�QPH�$4�r"�f"6�2b �.D@�MQ$�
6�"�i7���e�r D�p���RG$�@�&"�Dp�Q(�ԍ�&?H�0�2&�)�	�"��|�\~8�x��9�x�Ǒ��8�yYD	��t��O���}{j�7��jG�bb����;y���䃚�P�^X�nn�fH��Ҏ���mF��E-��Y�yxR��3���2/����I�'��Wb1�CE�U���?Κ��bs�-�Q:��sR�jܤR:{����Ǿ�+���H��^�8>��|N�Ő�Q�^����+9�*��;1ع\�;3�[�)��ޠk�:f`��ז��'�]�nkc���]SQ�u���Ľ��Ƨ%�'�����c���/;�2 ���;D7竁o�;.��`�I:����$��g���ㅌ��CeV���#���~��:{�B�݉�G9`]������"�'�9%����ף�ϳ�"YL\����|���b����qX�8�6�`j˻���������W�~�����<�F]/^�2E��|�=�G��n�7R]<�\����X�5s���)����!v���'43�=N{����ϔ���{�C�2��l-�qԪ	 ��k���{ȁ���~�����~���p/��O9�zY����}x�O�c��A��_�S*I��_�k�f��/�d� ��_��j)���C!o��ɻ|�-�Aw�$K@3�d&���Lu�r�Ig8i[����87݈�ˁ�AY�~M�URI{���?���ϧsR�̥���\��=�CQ<Q�o^�fKݷ:�i��С{�]�˵������&�����߼��Ǐ��ݼ��y�y��;v�v�bF�x]��.��^�`���FDNG0���>�8��o�e�f U��ٕ��ݮ����E�^s�;���`�NR�f�4�L9��
}{6��3��,`���)oՈAd�#q)�- 8`?]��ߪ�M!mx\���Hj�*-�w|쉮�Or��(�[�n��O�6=��b`�����l~��A��:�8w�����GcG	�
�0Ə{xh��A@�xN.��?�hȋgUm�6w����RG���-|��	������ l�<lX���T��>��7�|&�NX���<���2�f}��`9�tX����Et��)ل���Q>c��o��t�Y;�v���d�C7ܑ}�;�g3ۛ;�tš}���o�C�Z�i��d�7}ϲ�G1��O���i�̘6��ϲ{�M�7U�ê'���p��m~�<c��|.9�Ñv9�ps%Q��˙��+g�ǂ{?7������S��xa�8��9hO��^d����m�3�a�����Y���0���"GMT�l�?\���w����:�Dޥha?�cLP���-�\>U���z��]]R"![���T6!�� �-!҄�k;���n#����*�E�]�/u�b���lˎT�/�u���t�Y�Һ"��>Bs�|q�<q�<q��1�<��`���)W.,�^w���=�?b ��,�>!����������<l8��}9Q��T)�(�<���1�&��z{i��ZEiɎ��~�K0Cן��Q+��T��VQ�W���X�^8�ﻦ�?r���U�M�>.�C�E4���ŷڨ�J�w�q0��n=��R2��݆d�	�O��@1>�ϔ�H���� V�˷f��#Nsbr6�D�~�<lz[��{�f�~W���a�^�t�~��g�p;�}�^{h�~��B�P������6�{"�|�B�@Qt@C�����,���)wT�M]i�J�6
���~
�� �S�5�(�#��7Ѻ����/�h�����~jg�5ǐ�8�y6����>(��o�G�s�^�=h����;�?/}������ֆ����giͯӤ0-�NDj����l�k�G۾\pG}�?U�����t�x���d��$O�>��s��z�P�O���T��G:u��:����o��@�Gsי�"�cK?��ob�{�v-��4&벍����z{�����F�T5��o/���S�;���1|�tCr���Oބ ez��b�fF�Aewj%�pe����Ŏ����Z�#R���'����n��W9��ȵ�oi�P�ۯ��߼�~�Cx��<��8��I9�����ϧX��7�:��r�/�/^�h�8���xq�:p���WOrR,:�Obsq2����0��0L;�3z �v�ˈ�G�ca��u��=yn�6`sh~���z�3Wb�b����u) �wg���3�Ϧd#�);�5D�>�/������nu�]�\�[ѕ�ط��Y�/�V��EX���S4m��$7�C��%�S�I��E�Y\v:�3�3I�f��EAaT���N��'�֒��c�d�/��a�?1�ª;�}�{*��TW��@�R�vZ�Gs�z&�{lQ�0���Y������9����5f��}�]+,ȠI��$�~�~h�vjSi�K\r�Ep��A4����y��|�1Y���~���Y��� �k��k�t??���}��֟��{[M1�7wg������Sחt>�6�<�/�J���[$W��I.�h\3��٧����Q��n�6�b�����WI����.������>v���Ə{�??J�:��fGbu��RI���"�7}��%a�񚥶����̞�6����� ��X�ޫ=B��Sdy�Ѳ!�Ů�'t�x;{ 9�^��;q-)p,7ۼ⹶{��$~�z������xG�r1� L���>{}�w��Gӽ��%�h?�VYs������X$Ȝ�.=�ZV+���tyb��������mn���/j����҉��������gT½�=[姎{��ZYUa���<>p�꥽��m,�卭�w������j_�[��V��:�j$��V~��4����5�y|�_�����ù�yO�Cv��{�Ϸ���p���S�+*�/ #u���Qh~�O1uUF�d!�B}n��Zݷ�_�����{���lS��X&�]2Ԁ�i�-�^��7��p����~R^d�]���~C��}��/I�*��*�����~Z��Ͱ�0��w1�C]�qr"9�͡�����ɸp͈j�hyxJ��n��||aݾ�n��~'�rպ��/^e�y���]���8�4?6�k#��W]�TxJ�R��ڃ*�%��Z҈mu���Ʉ5��}�����ٽP�}vn.{��r�����(a��6f;�Zވ��:n�����O�0K(�l&<	���ՃHgj��E����rÀ�������وM���y�GW����F�c�{
�*�R����SB��^���e��3���"���R͚ƾ�xi��i���i�X���#c4c�i�!^�yv|p���|�E���LA$>ߩ_۟s\����{�f�֧Q�;sǭl$B��K�Ԟ�6�Cl��\�9!o��O�?zq�x�ǜ�<q��c�f��4����l���~��q�H��쟙�e����s�H��ίc���|�
��⋽���ӝ�.j�	g������G�G�^�nObs���7�7
56.�st*��nI��vx^����.�Ty���^d�X��XEC�ia����3��x�M��S�g�.o��s�I<��M��g>�p�,ĳ�o^���ί�э8/H�Cq�KՈY$�sj�u�����>Ƽr�~mO���d����7��;	[���\�Ķ�h	=CGq	ɫ��~���a[�_\,�B���A�A{�LV�y�2��8����Y�X�8�.7w��Җ:�p�V��JG���|����cB�|��?I�����T����/E����E60Y��\��Čw����g�� �է�Ȕ4~b�!�>�\Cu�K���0`!���\r��j�ou���c[c��"J��mF=��,���sO8���ցFf��yٜ�KpǏ!�c��O����s[\nH��@/�`?y�C�h��u .7�j�%�8�3�N��ӝV��Б5Y�,J�k��+!���h20��a0�!����s���>@dx2�!�G�ǘ���������p�gz*o��۬7'oR�:i�����b����1:0����??zq�1�G�r1�r�s]l����,P#�� A	i� k���?0��G������I1��[׻�7�z/�q猋`�4!E���*"�7o��s��	& A��	=��>6x�ŷ�_���s>wH�Lf}N���4V(�2O(�˃E��������sJ=�Lo*D�Gc�Z��:��ʟ[�؉.��f����?�DYnr�~��d!i/����������C�d����c��S�l��Q�K�Ț�/ۯ|Ϡe<ON��n��g����d�_d�c��3�&�ڲ�2�k��d�ۻLsi�p�!��� �{�ճ��5/�e��#�鍃w�<��K;�!5��6{�Vnl��Ϊƈ���N/�w{ʁ����F<����L��JT�
X����2G���E�����~���^?�I��`�y@���N���n�ɤ���	-,Y��3C�4�b�Se;�w�T�8?��-�}/��=�P�
B*�Hg��8����?J�6���ooo���}�#��t�{�v��@����h
�	���JA�H�ST��
���y0����r�[���*di|�{)�%!��Ыga%�cŸd2���]�y�pˊ��=�2�B=�����A��������O��	Q���Qp�)3���K�gJ	�-�h�/]�ٙrT��έ��%.�sλ�ϗ,�u'׷�?����q��<�x�kG��I��!�Z���ϵo�3�k�R�·�B�w����^��:����b���"�|��X�-�� �{���rܠ�"����(D G�
a����t3��q�^l��mek�7Ska��X����o�B�>O�����&��<����I&a���{^�~:a����ٙ�8_Dv����D�����-��f��	�yyX|�)�qdC��0�Q����1 �*�.�sz�"��[[��d�mQ���h|a��ͫ�2�#6�O�g�(��L�¡5yU�xՆ�WO��ռ���?�K4�C�E{e1=�O��%��}hn�'7�D��Jq^�3;�b*��
g�R��|EV��w��a�8?�r�}�8�*�����v��pW9yݘ��<���*�^�(,kWSˎha��0��,Dcxt�n�O��:��??r�7vҹ�:���/� �at�����p���ǹ��v b�妇+I���i�B��_��2�����#V6t�-�.�g8����l��W� ���߇R�&����kP�'�����$���
��]i5̎��Y�YI���h�OJ�\Nⵑjv����~A{ �|�����L��_�7���i��U�J��B��u���(���R�u�B�����U��u&Y[�����q��8�ǎ9�p���=�����
���]It6�*RS"$� �.5ɸgb�"�9*ڭκ�ά��;E�D�8F��'z����T�X�ћ�gmή�۪RI�?��ˁ���O맄qʿ�p�@?5Z�����m�P<�8m�јKfUi�a�Oto��a�
ie�� ��@,����/�Xᆼ4nw�اR��V��˼�+�1��j�d�L��an;��P��]�9텈{nU�aM,���m���ӓ�x�k��۟w�r���a����#=�x��L�����$7�o���/ܸJ�6�������:�N����'ͷ
I�	���@���@L?��֓��v��
w��Z7�~a���(����7E]�K��T^4Pz?OLZ�w�����]�0�oN�v)��A�&��(d��n��>>g}M~��ý70z���SĬC���e�iv�3��2 ����0l���������rfn��ĵ�W�q�{k)�s��34:h�P]%�`,h��.�s�up|�i�h X-�2�կܬ��5��oXO�=b��s^��U�M�|�I���g�0;U?W�}���q���V����\�!�<� ��݆ԝ���k��P�����Ú�c��ȉ-#��a�DSa�ȱZ���.[�-�gqNX���u`B>G��,��'�D+Sa��7-g@.�G��v<!�3P�6N����e&���������ά����'G�����G�r1�q��'ϓ�-�{��<����I�m�я�:J`37P)֘@30fp��8(�"[AMf�)�|�L�s9��p�L�c��+O�'-M���J�Y?55|D�S+XZ3��~�Tz <7���;�}/��󄐼���@*Xa�,���&;1g��cB�ƧSվ�u�@ɇ���lߘRzwZu�4v�"r���n�7Kt&|�ǟ�����4���Dnz��Ftskf?'*��nȝu�:�y"o}����a�>����nx�jR�M�>x�ϞCg>�(,F�3�w=�m�C7�E�vW�z��_�2��$O�#��-��Y�_�SL��'5�9�x���Z�7�����2��zv{���1RL~
�x�O��`��~�Z�o��~\�S�T���F��%8}G�`O�������v�_����-�BYyčP�m�"i�����x�������%�9�$1X�/�Fˁ�Jk�+��������G@������r�,��F3{C��S�	�^Y��^���g���\���H=�U�ke��m�q����P��.������-���Mk�pYX:�r"���1X:���u�ي{EFkp���R裐����zȹ��JF�[X�cG2��.+ǍgU�]ѶZTz���䃧ٴ�]G�\K�MYyx5�|�;W�,.��pS�$b]�̴VӝS�hkQa���4R��N�N�|;�jC���J��dt��b��ξa�9�w����p�:�Ǚ��BA��r1{�����s�ڜÓ���� ȅ�	C��v֥33N��L
����[��HQxG&��o���M�F��9��a�i���͖�PA;�+��r
�	9�mNkWs�V������P?f�pP����{�3��)��u}N�g��x����kf�a���x[��on�ZS�����rɗ����Z����T��`۪���rªTk�j��G��]�V53�Etz��$����1Z�PΘb��\s8l�.��a�f�d�HۧAh����m�g�s�\����BfΗ�b�ؖ�+�=u����;��)b�S���-��7{���V��&2����A1!���/���}8ۢ =�I:���J�)��X&��n�5�h�����=��SV�v++��'Wܨ}hc}�H��6�B�t�n�}�U;҇�!�W�Wb���B�v]A��qS���M�w>�l׍%1��������W�Bb�]Ps�ݽ�W&R�{AP�]�3M#r�oKYV ؗ����E�s���ݿ�k{Y+#Z�-�7��A%u�ޠ^�<��f]풍W��f]'��"�E�E�)-G��E���ٷ��j���d4sx�"'�)1}�y)N[X��ځG�Z����eU$�:�6:Rl=��:�u֯�wH���h���ػ�[�NK����r
�3fm���-b�����BwEo@�u��5IC�f���p��6��R�:�X�ז2��guX<��ެ�dG��`ۺ�j��O\q�0.�	HU����*!`nq��:�C�:>�mw�͵/+���Kv):�c�8��t��֊�s&�ώR2�-x��^u�[�W�m��t�w��diD^v��uf����%Pj���H�j:���dB�.B�ĘhS9�kq��܎����K�禾�N�V�U��-�^Vmh���kF���lzU��'�j��+i|�X���&Y�Q�>�z�6á�M�UV��{����)���MN%+�n�yn\�i�ok�õ�A�;�#:l��,�9+7�E&�$eI"��t��f���њOu�����%w~����<_�&4bd��)@Df_<P�ˡAvbٌcǷ�ƾ�>�kZֵֺ�zkZ׍u�ק_^>>>d O�r���$�R#��@$n�"B0��zu�Ƕ�>�kZֵֺ�zkZ׍u�ק_^>>'�󫒁b#�W&F����$d$IB1�ֵ�xֵ�k�Zֵֺ�u�]}�����}�Qr�}딒Qcƹ���f�v�(���������Zֵ�MkZ�Zֵ�]u����ǿ$BBI@��W�]�7�B52�&d��?���󫆒+�v���3L���A2����9�t���A�MC^ŸQX�4*&`ѽ7|�R^w��E�����c��r�&(�QAH{����ؖ��K��Q�c^7"� ��z�z�A� �+r#��k���/v���{�f�j���1(�ad��F ͍�sf&�l����������F8��<x�ǒBE��{��/�|����N���/��|��_���~���/�%Kν����z痿_�AU��Ĵ��ɛ�kx��,��3�8^�ζz�+9�f~
ȹf��!�/=p:-�e���k��+��'7�	)�cAܝebJ�Pj>ņ�YE��'�|����~�1����I�h=w}}����C�Z♙���%���]��-}�:��!331��������qP�lN�B�);����jb$3�y�b���S�����r܆��JS{����|��gت��r�4��'T���2=ϔ��Ӎ�0*�H��w�!z��f���E��l'�Q�FS�t������k�pڂ��'o�Ϟ����L��p	&��J�"s�w_��akp0ln��u�ج3�"��`Sݭs�����wD��2�yx?�"I{����y'�{<�sc�1�2�^���ݶwDz��Ͳ�����~���ݙ3�	���|ͬȟq֞��75�j��ãL���)k������y�U�y���*S������F�=\��v������Q׀���9wt�~M]�h�Y�kS��t��ͧ��M؋�(!@L�o%���l9WY:�u�Q�`��{}�C����������y����7I�]<�ڽ𐜶�b��X ��%yF����~��t�PUyIPS��6L(������D�lF��!�E���d[5�V�}�tg�P2�ppn��cy�Y2N�S5O/QN��D���p�8�j�抮Oz�.��H`���}���33!�Uy)|H~��GS@/���,��}��h���F+hzZc���]��U5�Пa�XVR�ho��[y�P�^|���U,���a7��s��Hf�g� J��^J�|��
�s���8S��#PEFs����P��� T!���{�"��n(ԯ֎d�4�XS����@K���;޾/�@���ޱ�����v.���{8�2J�{23���_{;�/T>���tV�˳�؉�߫�[�P��Y<��
:R�u�e�X�����c�݁���bfˇ�Ε���&Bp0���u"t�{��୧0*ݕ��6��ov�is ��7�[��M�louvt�2��K���A-�Q�<�[2_>����!wzO]KTQ;3j�.,������}#k+gZ����xw�ܤ�wǷ�q�x���=~�:�r�f���o/̈ҡǲ.��R%[ב'$�}o5�P��vc���RT+�
]�]봉��]H�>Y���b�4�4� u~_���+�g�d4���ˉ(�}OvP�P�u6$o�Q%��%��^����;�}��ט5�������q��y������9�B��c�>�֙��xx?t�du��S������K>q覘���Y't��W��gVA�>��z���eQ�~SS�'��T��m�ږ���M��H):M�L̈�"�^=R0ꩽ���匴n��T�8���F�U����W�r:��8q���̺�T�22��cl�{�zs�Y(��^�M��Ћ{��S��8��Rx���X�V��[�,����#<��׭�S�0�SP�����@�Ǣ}|�vr����]٠x�w��ǀ�:3��3Y6U�E�:z��z_�s�.>������(ob��L*����3d�ݨ7��Y���К��i����$���Zq2N�Z�.�d��Y*�ֳJӣ��Y�+V��~ Яz����T�3�os��Z���(�:�ns�eNS�ka�L^�zk��+�8y�>_>rX�V1����F8����խ�]�>3�kaad?�IO���b�>�	\C�N��ךug�I�Ļo(�yέ�k�T��N���%��0�j��~1���/3����r+�;�M���ףb ;�{�L��d�s��s S�=�"F?r>�m�=�&���tF*e0׶��<��o�@>죎2��%k����)��¦�o��8��V6xω{X���������4"}�,���p�e=(#f5=��N��R�gf,�����6NrY���f}���7mC��WrM�å�]Dfw����W�Kj�� ���;�G��BW�����)ԍ��9�ǚY-m�����_��w�@L����ħ���rƮs<�كyI#e��L��[@�?�t��� h���/���y2��w��Yp%�����Vv���4�l���}�t��,@�||�����f8������-�V�6.�����q�r�uu|6j멷_b,��7_v�i�w�m#A��"P�%��73�7��E�<��z!�H��B�r� �j-9}X�y#����I]� Q9�B�9�����ノ88�y��������]�ÿ��|�b<�|7*'ͤ�9�#��l{ׯ-1��6�gs����tع��N�tġ�p(�� ���Ɲ��ك�ܜ��ah!U�z����eU�=4���~�"4��W��C��x���V�M@S�p����O��]FצE_���mҔT�:�
��{Y�أy\L�;��5������*]�X�9@��N�g)��v�O<^�C�Z)mo-&B��x��r�-�E����Dt���M�P|#}\��b&5�������8 �.v�2�[����
�m�q��<׷ҵ%���.��[7���<㧻����x�?i!5���������L�/f�L%�C�,�����69%��ʮ��fz���o?�!���	�9;�������A�$H���d�>�6m����������^�@ީ�Zv1u%{�޲Qܹ��t%�2��C+
�Y�fdC�g�}D����»��јP��仨��CWbLq7���؊Y��P5j��;ղ<��3ק��q��88���z��|�-�=�k!|0h��ah�����=2�zټ�����VB;���=��=��g"�-;8�k��m��|^���f:��PYE�U�[h��u�`y-��" fv���,����K}{1,���W�N��Z�/L��q�ŚK9AL�ް;Xct��>z�{���*k��?M�s���kN}a[ֻ�q��=S����`�ig�ҕ�!?�O\.fq�f�����{�`C�ێu�,[� �ϡ��;;�M��N4.[w5=��#q���;�{F�����B\f�hx�/5ʭ��Z����\��ݍgf�Z$�Z	 �v߷,�>!J<��Ly�s^btQ���_Z7g��/�=�L���	G�Պ�>��g�H�i�z�KԚw�|W[12�N-*�կU������2g�sqNl��������)y�l���le�鵦�D�ޮkfؚxb�u�������&m�ܦ`��2�>�_<_<;�Ϻ�<�D�j����C���:����F��Ii��+������T�*c��	�)��B���_������<���������¯6}r�����׼��	Ke��m\��l��[�k�{�g^fV�źie�OB���Q�z��-��d��1�1<�{�-orP�E��.g��~��k�K���s�L���vb�ԕ�ݷ�z*9	�;zĵ1�H�1��K�#d�n8���oZ�e�����vl�I�."{8�Y�Tʊ�w���o8�����B��,�`���Y Y޽���.�]>�=�l�X���ϼ=Y��_�_�����>A��hN=���k��~�ܫ��e�N�X����67����[g�m7�?X�d����p:��^�E���y��&S�ܖ���>���;�vC
ޫ����9�<-�N%���݊= N;3~�m�8	n��"��H���em��.v�`�B�ײt>��>��}`�YWNT��y�[�Wf��#������ȿgH:�kU��r c�~Ѻ�o�ÈM���pH	��o{B�O<�,5�����d���筱%؟�s��迋G-X�&���T\���vt�7=I�W���;�]�+Y����S�2Vf'3c���h�5L�V$G=jE��@<�M��"K��&٬Zd	�iwC������{=��@oG�����y���Q]��z0o���J� ��+��P&:��*�5{�h8���GwU�36y�o<<H��xq{�]Y�a��Q�Ȧ;��Ӻr�#��"nz��ϑhPEy1�)�P7i�l4�<��i�;yq��/l{���{���@����^������//��>�}*g�� 1#
~�4��T�n"'�Z�U=>2�fj�f��d]�D������,������Rx�~�*�覶����om��1���{���l�Ͳ��q���o7�Bۭ�W4� ^��ݓ�G�gpQ�92����8I�u�}�ԠM �;'��G�k7}�u��=�1��]�᫦�q97bu�+�i�-��v�ٟ5�Dk�f��Ʌ\�L�;��n��Jϻ'�zQ�Q=������%��{���"ռE'�1�3�E�Н��pwJx����Y�DY��\��[�"��:��� ����� Vl�1�����k���˽U&jƃ�r�Dޝh.�5��k�կ��^J�:W7S���X���V�����W����������?���[RJ�w~�$pz������<nUuzdwI�M��n�	̈��9*RH���-b���z�_���uDt=�x�v��c��ʑ&��F`����e�{�%�a� ����ۙ
x3�>p�tt��#��b�`J��NYU�3'����H}�,�~�U	T��}���\4��I��z�u������H�CT�)�H���7�\��ƽJQ	��L���s^�ة��Z;��3?i��h���]�32)�ia��%j�d��ן��kε��-{�O���Y٩z�b5tõA���5�x��^���^V:g�;}w�B	��xxSq���oaV��$�5M�F*&��<4�7������G���Sꇩ��u�ٝ�͢ڢ.zU�z�潈����v���$G�!C�L#&1��[s��YMaI�*WYj�G/r�N����e�"!�St�yk�Y٬"��0��U1�U;����l��]Fu��<M����͹l�۩��*޽�W]ܼ��퇊����+�K�-����z�����Ǜ������y��z+cQ�����������G��+e�M܀U�M3�@g�U�j�6v�sLa>�ʹ�7x�j��J�y{�~���� ~�  �	�76�~ۚ����C��!|�n����Z���M����P;�^"��f[a_q�<e��]I^ά����̱M��j(蛩�/;�����u��;U	���!f�)�vf��k6�'ϗ�l>J��#\3��!o��ᬫ�U�ϷY9"����7���`[<�۸���v}����4���a��C�0�I�,�K���Y&.��D�MC{��P23znʡf����~=x�B������_}���,g�0S�3?y�[��i���Y;[�� ��x�o �;�zFv)p_Nuwe���jQ�
o-G��]���ɖ�Z��r�?��&�c�|�����|�W��كI�`�:���,5\!�6�G���uf�9�;kT�VaĻ0��g��1�1l��>*��N��7:��Jf�AO&�4G\�¶K]N���"�cI���A�HOLθA ���T72��fAF�ܥ\�^q�F��I2iݡ�g�e0��\���iqOp��s��¹r�f�z�o.Wu�Ͳ҂�RБ�w��KU=�B�ʽ�D���Ocx%��.>�h�(u>�F��q�|�mM,��`��a�V�[g.7Kb�tK�M%��3/��K2婴�~Q��gA���]��hk9�T�}��eK$u�C�+7*ٖ���@��H���3u���y���lp�j�u���Ϗ_N�Pv�^�z.��ʘ��ǹkM�'Z���w2r�W��6�r��V�u�sL'���vM]�Ńa�mfR���3rM��oC�yZ���sҫ�l;$���
oʞj*1��r]nGl�A�^�������;s�m����V�Z#9g�cn�sɽ��Z�"6���g���t���f������˗|,���h[��x���z7�5T�n�N��(��d"��67Q�s���6i�5���.���0�"(ZWsL�7/@F��Oh�1�A�ҥa�yy�Ո�:�f�5EnN�ȴ.	S�7d��8�l��!���hi�*է�����^�;���x���w��tٔä�Y6ճy�֧�@])�l$���9V���@�S͒s��6��ދm�!"mH_��A2KȤ6���D����]�8m��vD�Z��廰�t2��"a�&Wh�e�b�����<ׂ���2�^eg;��DV�;���ݙd=�n�Z�OE�g &��R�݌�R3{L�2���E��ma�sXjh���*jh�a(7Y��oZO���O4EN.{������W֯�"	kqf�S�q�b��y���T6@9�ɼӖ����kL��il�M<�Ҥ}ޣ��]��B�f��[B�G:�66��i:Ѻ���U>{�1v�5K+m�d��wń�Ck3k��r���v�Zw���q�8��ЋW�B�w+ �|��d��@�۾,�O`��J�8�=������]mv6v�)�}�a	�D��9�(�A1w��犪���Fjې:�/����)]����v�����eu�5��Pβ�.�z��--�JyR����$���ʜ���{�N�r�ö!�DKt�b�h;nm�"�5TYG�tP�@���лX� ��Ti�f���	.�� q��|�D��b2N�.H�rD��mK׺��Ĩi�ͽ�� ��>�	&�@��W���o���nT�������ּkZֵ�k]kZֺ뮿�O�>>p�D�FH�a�'&z�l&��?{��c7��~�����Z�Zֵ�MkZ�Zֵ�]u����o��ܲlE�\J	+�u3@DEHSv�����}}q�kZֿּkZֺ뮻���o���4Aj(�I-�ݧ��h�b���zVrBH�Z�k��\kZֵ�Ƶ�ֵ��뮾������$`BE��'�]�w��g�2���o%?�m $G���t��ҍ}�M%��S��(��d��M�Rmx��]zեu4D��ܾ�w|oo.�th#_;�J,x����&�^��ĉ븱G�l��5}W�x��D�2Z���I'�>�>n2B�H�0�m4�cq�	m�1�ۈ%l)���m��"�S�?D2�F%(�\�؈���&*��!10�$��3�E�d(A�4^NB��$Ê����wʖ�W�a���B^q��ֶ�$����h��2%��b�
���ĝ#1�����2�iA!��@j"0�a�(�	%<�J`B��|R)��)H�`�&H$��^�F�2�jPm�PRD`M�"F�m�R
FC�	H��Bۍ�!����d��$2�����#�f'�"�F%!��)#H�Qb0��CM�0A�:p:�"6\�"#ND�J2c�d#湛4����1ǎ.8�����׾�c�����5�zPx�	�k_��{�f����@���o!��z��O�����fĝ#Բ�2�t��	ME٪�N-�7�ٙnH*����>�g���>��Jg�W,�`b�ӝ�=��&�:�F�GuP;쥗�7z|��}��/<E32(Z��SS3-W=5�+.���&�Fn�<�(��F�|v�l!˹�ԍԖR�7F��2���OTe{|"wL��ӵ/paj7������3�����\�4ˇ���^A�w.�Z����^�vS���3�<n���sy��lұ�-)�'Ђmv,������\DU��>�Ԥ@o_P�;�M��K��Gd�G3�O֗��%�b|/9]�8�"g�ǥ5��3qy��T�����1��Mv�y_���k	6�ʄ^�ڸ���"��&"S��g��xT����;��H��6�6e�������7���V��ٕYWԉ[r��R�鵪A��w3��t����|d`[sj��oJ�go��-�����rŧ��-�e2��^N��vt����贔���̹�M�PH����M�dl'=a�-�^�E�vˇOP5lQ�8���VE�N�^]��c�+2op��,�����HC����#ǎ<�8�<x�����֕�l�_��gL'�J';�W�|��{ �sA������)inn�^3��`�{���㽦9���s���F_�I�r�G�������ٻG*̽e�<M��2�G�ȿ{�#�=�^�k�]p�=$R/�_ �!�kF`�Y]��B������8'�Y�q���yr��c5�řP$m�v�n^�_���Iq������� ���h���Uj"s;w�MǬ.~�|�l[�Hs���gצ��3�e&y_����۔�p�sw15=m��}��@΢&��
ù/��I(��<\�'z� ���g��y��e�ݿ�����O����2�s�����{�.~����?
��S��%�ß�4z�+��ވ�cӪv� A.���m�j���G8��T���o���|*~'�Ɗ?����5lXO����ER�.e�bo-P�Ԡ�ɶ�͜k��ܧ����Z(���$���K�+�lƤ��d7ź�U���/��e>?q��W��I�0v��^�<��p��~<{pq�G�xG�y������Y��`N9�����:��ٽ�Q-p���uK������]{�ʷf'B��YՇ��$��x�3޸y��S�e���u[س5C�`���w:�qE���Ӥ���ݧ�l���49�ni�Ҝ�w�M�>��~�F¯w���W+�������(󘾦禥�����(���w����U~���e��ō�B�~���M[�)7�9{�����6�N����(�������x�gf<�|`,k��'�ͱ�����0"�ks{{I���Se�o+�Xj;��6q��1���Xc����2JpVm�D{w4����Cg���-�-~8��wg7�S���wh�b�kFl���~���n�z >��{{��*Ѧ`Y�-�6���%5���c�����J�[Rb����Rq�y�� �Ӳ��h�hA�/$.hår�2�w-e�Y�36����O���9���*�%�z�Lz�޿�j,,�8�&$q�5������:�`�Q������B���Vhc�s��A�����o_<�_�?�x���q`c���bT�K�����g�W�����G� �<����{�s鼉��9����iYl��vwR$��9��3�B���؁7�JzɧÞ�9�������ih�yj�A�L���������wQp}~��9G��+�iQ�� �� ;xxv��#���p30/`�OI��F|v�³�PkCy�%g��g����(�V��:M�j/x"���?�������i�o7�����
l;ߣ.8�y$��K�p3���e�^%Q�n��Gi�f�0<�߿?��gXEZL$AH��>�^��\S�E�n=�����M��b�����4�b�{�R:Ot�c:����g?��y���A\��b����O��M����oq&b�,���$�SI�j��˷�tK���?v��������2{W%�>�̙�3�����p�o�s��_�2oE],	&�%;��s�"���X��P�R��ؾ�׷-�W��f��*�[/��i�#Ȍ *�݄UR�v���sa��$�W{-)�P�d��`�S_�hI"�j��%�b�O�����e���Yzbw������~�8����������gJ�snV�U�MY'���Z5�G1��[ʹ�rŴN�Q�(��6U��Q�(�V���e]�v*-���v�.��Ǒ���������,�H��������l�o5D���J�e�{��z���U����[��h8��"�
Re�.=��ex�R��ސ���@��FèSYwy�T�yXq������,�R�ݲ�9�37uw'��j͙Y�d��oj�t(�/[6�ƈjʘ��n�]O-���xl�7���r��U�.�f��=壡&ҵ��D�Ü7��"O2���ƅN[F3(L�zM:L2n��H��;'�ۘ�B���&�E�0����V��[����93�҅�6�K۴���_Ձ���E�;3�>Λ�� z}Yb�+�h���urء����ˎ��ӑMwy]0v�:�ك�͵{�67�v@w�
I��>Y�D�L��b�҅��e�{e�"�s7x��uM<J�{"}#j�n|���\���5�I�'�k)��㏈��m�ȷ���͙ }��n{c+^}�+�X#a������m��e��c	�^dQ���o��m��M�P<<�p;֮<�ƹ�Փ�E��P�w���i�=F;����<���'�d��z|pq�pq�3�b���9�~uf���v�@7p$_r���%�1qV+^�l�⺚~x�'Um� �ũL8���A�[�0�-�|W��w�VnK�Dso3�K�Ma���/' ��S�<4����J�d��a�aR1Z�SOx$���ٷv ���;�,G��1x�;�o�G/@��;=�����h�n3צQO�S�{�ш0/}��S�iF�{;��R�W�]|��;������o��Y.�<q��|�����X�0k�s�y�71�+�i�����jDE���� )7޼����O�`��q���V���:��%����@
J�#O�y�B,|�9c��;-����6L����#W�07��D��ZIj�S�G'�aװGBSs�mTs�0Ю�aOjqm�6�����qP/���kU*��WK]��NK�!�s5�sGw��ft�:MXo�e�[��s�+-7Pa;r��G�Z�Q��B$[��'��`s����I�e`":뼌��Lps�>�ԧ	�{�9��}k\q��qǇߟ=�=���>�4�ĴDN}B��׉��=��{�g�{z��)��^�[��]9'�~
ӳ��n	��C���C����X��N2���_JcC�Bw:n�ngƽO�o�k�����ɴG�_0 ����Û:��S0�;�v.��sH[w55��V8Uo���].��mP�*��p�f���b&��f@~67�,����@�S+���c�f�u������r�譓�sK���X���/{�=) A���~�l�R�&$����[9=���b��Y����D��}�v��h���7��{��s*�d-���zw��G���{:�[ш��5-��ރ&i��!�M����V��A�p�v�ۙ)��׭i�nnyj�T��L�굻>@_G���(������9��~Um
�ZU�w+l��r��[x�?�<E1F��Ք4^'��0�&fֱE�r���c&���-"���0UX+��{EW�}D��0��zY\{�������>rY�oo;U�c�I���7i�����X�v�*��pq�q�#ǎ<��_��{���>g���Ss;���592�ط|��=��͙�x�o�W��\�2�pԗ{Y�nǲ=��l����]C�t_v����MAw���=�y2�}��KE��	n�L��dk��tegM�b2&]s�� �G��{[�x����f-�Ć��l���[�XT���4�����2*�c{$p`ѱ"�(�Q��R��<N`�4#~^m�n[��k �}{�V ��G��B���9�7+��:E��0�y�f^f%�2�FdwX%{��/hjn0�C�U����}���(�wQ���GV<z���1|/�M��	�����wޅ^#�VΖUW��\��kNf�������Ϋ�`,�vB
oL��]N�}#�nn^�xxC���F��������M�qQ��:�=��B�~�>Nw$.Yh�0����4��jN�ASF�zp��{����<�<�$�#|Ԑ@��G�=��h�|<�6ܱ�ei��$�^��/{�������ܾ�E��l�� �1�3�{�ѷ�_��8��<pq���w���g������m���r��⚜�N��ѡ@�7fƽ�əe��9.��w'���sB�fvo�Jף�g���w�Bgzl���T�:$����\�Ml��#�wʎt��������+n��}9���3���m�d�꺚��Ӏ����g=g>I���� O���1�С�{��n*c��^�k�ջ��g+�{�-K_v����y���v���E�?Eq"���nn�j��g��{#ɧ�@��g8����ҏ[��H�/��+S�ߒ������z�~�X㯆Tv�7�z��9\��ݓ>�l	5L���=��`�h�p|o��Z"{:Î����}����,���m�o�`�v�tP���H���#�n;ǞE�y��ݕ�c�<a�԰�A���w�$o"�V��,���{ޞy��r)������^+ҏ"��ΐ�3�+48Ӱ4���`/RB�L�q�p[J��̫E�����4Δ�l���Q\�]��|����QViN�����J2�d��<0������q�}ixMke5�srf���R��X>	��D��v�]5+U����3�*3�z���&}x���<pq�������"��O�'隬]��B��z�z�1�6&y���,v�n�-^ԅ�`:�{2��W_���L�Zk3O���W-c��M�{G~�׿u�5)��bU��~(C�K���kB"���vݜ~��d�$�Kz�)z8U�𭀢�ϓq&� i��Wga��z�"�m�;~����T/�lz��j�G{ ?+��sc{C����^v�Z�j��sT���I"ƌ���6�7p���M�NmOZ)�`�I]7Wl�a#�>���^��dv����j�+.ɺ��L;��[?��v�(i��v������'�I�q-P[����֞3��^�kO�y�7}Sc:�jҔ�q�"�2���y#w��ϸ�o�=�
���z�'*�#�p�6�P�u��x��*%�wK�0n]�EC�k���a�w��Vu�B�{���]*2:��B!�>���}E��ж�{j�u�Y؅�����\�Z̥�(K��5���f`��Y�nL����Yv����qk�o�I��s���
4��-n�O ���y��MY�_Py�_Q��t�<�3�;q�v�L�H/c�67*se��U.��y��w�=�|m��ڸ	�Enʽ�Ȗν��Ns�p_A�j�V閵�Ә�:[i0�Xc!4�/�mE��Rf�Is�veen�{P��t�8�Tר��32l�~��FX��z����_v�!\�q]sηw��{jU�"1���4��|H�C:�,`����,��VHFæJ�U����y��ڃ�����Bz�*���uʢ{���l�'*Vj<�mZ�;������v�=�j*Hv�b�:�\�w�e�eq[nI4�Z�-���M.7�*�v�R�}|�����]�-�c,N��,�����r����Iʎ��R�\��t�L�l�6�i�c�T�W3�T�"��%�"p��WH���$�y�����A��a���|�<Q�M]`��dW��b ~���0�b�U�8�,5�ܳD�����p���]0�|j'ԉa تR?@H��rB,����%�Π����΅o�$V�=_&��fJSc$:x��PL�n��#b�3_���ڡ�l�/��j�g�f�]���rv�fd�W��_wEs�P�w{�R���q,�=r��n�L�2���@���:p�t:q�G��강���T��	eR�'3o��f�Wm��$�ɀiѭV�ٍ���p�m�$YY�8Κ;��Z_8� u��z�)׺T�7�Zqf�d�'��e���%1��p��Lt�8t�P�{��ڻu\�����-�9�����w��P�J�@�[���y�Eexlgl�S�q�r��)=*�5�4G�����%���`�Y��5*�2��5��W���8��+iQԻ�����qJ�$�Й�X�:9y�Ƨ���w[ͳ+�J�{�Hk� �Y�fB�ĭ���C�Ыw
tvNr��w�>��|Ǝ�I�<᫥ݠ����>���Q��s)��f�T`��ǎC96:�S�d4�1Ա��w���v�%d��%�S��sVm�"[�����K�E�i˲�.�1�w/�wȞA����ѯ���nD��sFC�!_�^���Ƶ�kZ�kZ�kZ뮺��� HEɡ,�[ů��Z7��G�_�_Xֵ�k_�k^5�k]u�]}}c��{��fI$�$	��b�u�k���ֵ�k^��ֵ��뮵�|||�d;��!"#`l�S��CϘ�H$��צ��5�kZֵ�mk�kZ�]u�Z�o����W�޷��u�J��z`���6�t���ۚ������� Vk����\��o�i(�ڽ+b�<u�W<m�ƍ��ƻε�Ѡ�v�������~u�\�����W����F������}^4b���^�
�6�7��_7R�ٕ��3�
�y�x`@�4�`t�Z��²��Db{]m�����^�]z�~�C���^^^e�U��V}���׊J4\n3�k�%�f��`�����|?Do5y��<Ř1H��i��� +�j����t��@��]g=C����y-C���gهO3�x�q�3(^�Ѿ����'��ރUp���S���VeN��1�{�4d'� s�-�ך��{�v��O���#jq:5cޣ��U�)i�y���h���`����O�jMz�ҋԧ��2���ϯ���%�z���פ�=/b��h_���P�j��}"�������u��&v��C�^��>���M�tlz]zXK��>�u%O��I������$�k�߻[�S^��V�����૮/��%�jߚc�K�Û��mhg�g�f`�z;xW,�&�Ap�V��ߞ�G�=�e���c������iEz�mo�es�/O��t����� 䜧��7�3��dC�O����?gAXc�On���c]��?"�`��쵹_9
��/�P�`&йZ��H���c����].�W�J��"�����*�w����p��I2�wb]��y����^[�<8C��קpq� �y�<�W.ޟ�Sz�Cx��s����{��ߴ���K��6�p��1:v�$b�7O��-���ڦ������v�e����%_.���5�ɚ�z-�	��]��$0k��}�_@ܤ���=����o{Ē����)g��<u�gƘ���V��o_|0����Hų3ag=�� 3 ��s�)R�[�[��ǻ���/d�=Co�E#��0�jqF�^��l�������s�8l+��X�	����0i��"��+%�����7n��7�-�v���J9H���焀���7�]�=NZ;��9e�e�k�v��jD��P^��4_�ḳa��m\�<��!�\������G�-&��lzčCs���`a� ��U��͘��������^c�Y6[K�7�x%�N���;���V�rvfA�D���V��-Fɤ-��:��S��U�7@)���q�V��zS�G�cJ
��D�{Np�}\�8#���R�+w�i������q�#q��|���u�u����BwP`5����p�K����*i�T�!Hk��$cV;1�)̾���z��$,�T�!�����������������('��)�Bo�i�x�uvq&� |��!���R�հ��z3�C��昚��%z���w����qe�� �3uR5�K;�:]�]�}�R��Zܩ�Nb�yP�i��y�Ky.��h\��T�X��!��'�m�W��R+$��H�꼻u�ߨ!-|���&޿b��Wvҭ
�ny7f�a�y���R��`�����3x�+������x�M�T]�ٜ9���-�͠�|�������6CS��4�;��#��oR0�H5��^EM��.�%�8�o���ߟ��h���s����z����;��ٖ8]gV�P��9��xu�����c�c���.���e-Tyz*��ٕ��N�WH�������n>K��;7�j��!@M̹�r�ӛ�6��f���w��ԅN��-����� &�E!(�_�ߪ��]��J�㯼
�壱l��`�����,Z�Er*S�T�AR��fj�pK��� ������=�8��������*�*;�Ś��}~�>`�=�<b�t�p'E�����!Gs��YX?�&�,�{���J=��`l,���ZF��mv+z2�C�~ys335�Ur����������%+!�60c�<.1en`Ȫ��=vsu��y�@g��>�B3o�3�3���>���=�;��C����"��᳚�����U>ǎ��	�_U����� �,sSxs[=���G77%�{| 5����!��q���Du�1R����8龕[+&��]�؛���\����&Fc�z6�OP*��R��Dٸ5T!�������N�7�If(��^��h��:(t��Mvҩ5nt��s6�"`37d��������k3�M��H��ߎ�&��?��}#���~V����N$�0l���u���u���[t���1�2[tN�c�M����n�鿋�3%��h�xGݛ�h�\�	�ܫ[G︻�e�a�z�g��@����%�<��&dwi�T��o{�o��/�7	�~?_�8��<���Y׹�gߨޫIĊ-����3O�+ ~�� 6�w�{�l��c{3^2]�h���w�E-^���Dߺ��^}]��J��
*���+�
�MU�F�Tc��Q�m\��d_)F�Ƶ_(fn��z���}]�*=�ϖ�ٰ�����3��7M��~ݭ����Rݢ�|N/3մ���S_�����3s�^�K�s.6k��g�����w,jP
�<X3�`5��\ES2RWf�L��94�NTy��\���z�r�����K��ϸ�6��C)7<�L'��.����O[�t�.���oi�y��n�������$�L63>~(`KEv��K������,��#��qf�F�NFZ��z�Պm>���6���U�*�~��߬�o?Y�}�^#"X�5)�)��5��w4,��n��X�OJ���qp�5q��?Ď���`���Y�;����߷�����L�+S����
��{���|�߰��G��mm��a�p��20���ʅȩ�����~>�ǎ8��<�=���ϗ�>ޡ	ѝ�Cኈ����X`�Fw��ޜ����ʵ��^���n_f��q^���� ��[wQ.�S�|��\ɾ=��emm#��=4���fv��^���.,��1a57�U{Z�e��4-5�j��q�����>��*�=;U�7��RzzBIu��C�L�y�O5�y���R��C�>���� �No��y�E&2�CLt=kL�xs�v�3������ ��b����oԇS!��ށںk�Z�m�N���:h�-��%��s;��n��m(�XK������*��&�7�I���i��+[�Lnb�JRݳKx���g�Ǣ=�Xk��.�Y�2�ٓ=�i"ru	��z�.��Ш�S�5�<�{}ZƃYS��i�b"�H�e�)-�'�y��S9dn�ܖ�>���eN;J:�grZҙ�94�E^����~��Xp��u����}��^Y��T�}Wd}��h�$.������ץ�d����`����2�k����6ږ�.�^�҈��\�;4��`L�H�CV�l��uvk�w*홷2�?���g����^^^���z�����\���w�{y~dN��q��/�������V�SOQz0�˗svN�s��Xݶu˶{˾�X-�CaP��<�a�������5�d��y���+�Hk����27s�Y��ś�\��D���`!��f�.��fqR��ܰ;a�[ml���'Q��Q�VJ�y�y���K��IP��zҢ�+D��tp�2{��d���o���O������U:}����4�m���vMZ��w�!Ө��6`��_��۶���hgEx�(�ҟe�3��f��iۄ阭̽=�`�N�zu{'�Eh{�۴��}L�e]!�q%:��?w�:��x�0lYq���,�OUb��f�(��!]o������LsF[�����9lejf<�B��9b��ĉ��֖��m�7C�����r�t؁N�úC����U|#�I|1,�;��z�KQim�)���6c��~�c�>��y�~]������ݶ �o/F���i�Q�ܳ�'�t����s�և�n���޼h�<�'���h 2�}G���gi��K*��1��H�Us��Q�;�wWv)�J[َ>��2��@U������=��]y�� �?�lnfoZ�^�J���6�$7#�����O�a��p��g�j"�v���Qc�냛����YT{�$�M{g�W�.�N6ln�k��B��?�=w��|�0N6v�Ϣ=��3���'/�*�#o��NpqNZ�{-jil����5�>���F\��j��������8�������FF��І��<�vU+ݒ��λn����No��E?������؝AxvHfq�d�t�︫i!ǀ�Wna,ⴳ����}F'/ݱ���&���cd��g'���7Su?I]V��UdE�Ȯz�z;H������o`F��2S�i���~���RMR���K�WC�׊oE
��o�/
�"�incg5��7�O���
������u@����>���'{ze9`�z����{�*�z5v���m��riwj���|�T�<��,�(]d����ǘ�7z�N��enp��U��K����8:z����gkܢ9F��=p�\�ubR�><{1;i�WG����ݥ�{�|ɻ'צ��A��p���� ��߾����D$)� �WU�[	�ʮgB�����|��X/;f��1ƿ��]�l�5dd�n���^���	�����>�p}���J8��$v��^�g#
�E���$93�����������u��s��y�^:����%��KK*������}�7�o����w���1Ý��zo6�8�ا��g��9�|��P�y�VGFכJ���n>�E��.szI*MO����ؽ�vn�6d��rK�������N9�b�F.�'�N�8(l����;�ںc����G��Y��.�o��0�w�G���n%mc��[s0 ��}~��S��r��:32�D+���/j�D4���DT]�X�[*�*z���$ml{7��<��3�U�묣�����*ţ3�y�F�jVdW���Ŀ��[gs�c��f��ٽ�S�ѳ����>s C�桃�>*j��</��˄g��X�Z�Of�*)ت:���[�8�a�Z�b+7B�975�C5�";:�W�RJ�a��v�C�ƕ�nr^��؄6#�#�7(_������=ǎ8�8����I :�����}��<��l����Vx�,* $-����u#��UK:�x{���"Ќ<*�|�������<g���Y�����[����&b1�e��]��n
,|��jʜ ��B�=sA���N�+I;x�վֱ�O��c��p��j�`� �UΎ���1�,��cvU�қ�f���a�}�96�2��XLrj��b�n0�U�'�}��&h��T�YĊ�u"�͞�7����7�И;� ���Z:�(3�L�	":矩^X�{A�i��%ʟW��ٺe�\��b"N]����Ds����r���MlxD��d�G��[��K_��Y������U�Q��gvw�>V��U� l���8���ݞ�&zy�Mbu��2�
�����B�l�l�`(mO��8��R�ڧ�ؽb>HgȕL��a�2���&���Y�r�,3Pլ��ǣnv�W{A�/��F�e����Ȭ�Suө<�������vT�Aǽ�0lK��7"�ŵ��5U3Ͼ�%�@���c�����l��+ �/3ڥ8��a���3�nT��Щf9VQksR�eu�X�I򮞊����B"0V�qi��B��(��z��oH���2��{|ZrI+��!�hL6�I]|2�M�c��[j��ii���r��]ݔ�g�iLw���[���N��F�l?[9��,����`�q$Dɽ����ٽ
��8��A������K7ېl���ڐ�R�c8�j�����bi�Pՠ	T���B��r��&���u�TbG18����T��gJ��9O���*躞/�����846-?a
��׊n<Ưb&�&�W"&R�3�m�^�����f�k=���1rZ�CV\�e*�V.љ�M�9:���߯���M^���އ��
�e�����{8dZ�\��v�mc�#e��_u�e�o���+�<����
�'<
uf��\;jT�-�Dlނ�kU�S�K-ә��ԫk� �*��y9���:u��q���4M�)-����1#ڃZ��}Jq�ʻ,3m=��*������hB�ʪ��[[`�m���d�)�1�J���o�V��B��$�FG%Y��Bd���6�4<"AatԟW�Р4�������^�2����f�x�7��Kp�s��Ζd[�l�fڹ�lHt�D�+��d��X��j��hH�=b� �L�]��>���u(��mZ�)�E�v����y����36�����ՑV�;*�uQ�<�S$4�&�G�����ؙ��	!�I�G��n�2�'��aK��6�gWR0�`M���#�5��\�`3V�E�5�[Siqܙ6���'V]�x�9�wN����!�غ��L��0�Zn�q��[slN�+�m��amN��%�+/)��C7)c:D*PY�n���Q��O�+���xV<ͬ�"Ch被
���˗b`e_q���KV�CA�ײ�.�j��k%�ޖ�/e�	� �]�FC�,���F�$�}�VAK�W(�wHQ&�a��r��0P�ǲ!�y�=)�s�Z����f��^��V�����c'4p����lHμ��UJX�ܪ��*�����Iq����x�[f�õ�0N��3f��/H�z��r*G��K��V	ѯ��iRI�CD��z���"AU;z9gjڮ��Ij�m�.TX�b��NX�=>�5���Zֵ�k�Z�Zֵ�]uֿ���y	$�D�ȳ�f�FA�&`a�@'�N8ֽ5��ֵ�k^��ֵ��뮵�||Bǻ�#�#fA�ȒI"��	 �=:־��Zֵ�k�Z�Zֵ�]u־��~��ů?{t��1�m$F�! G�kZ��ѭkZֵ��cZֵ�]u־����gY�XE$��ƞw4c���9nhۛ5�W��_i��{���r�Mx��r?<���ɋ'�����w��yݷ��C�[��A��jC�m����Ǎ��)���#k��r�c�\�úܭ�9��zy��ޛs�� �2����0��jF��@�P�&B��J��TB���1��.D�qB\���(��B�NZ%�h�0�"$��1����I�\IH)��B ��ȧH�F�l֌ ÅΒ�r�Y1�.�GM"����Ԫ�=E֚ow��#�竂]s�_\H���"�A)
UA�J��`�M/�M�O�(�M��j(ۄ�r��(J�5�i� ע�$�Ĕ)0O�j#bR�(M��F�)MEI��B7�jH�G�a�(��1
I(Pg�d)2�$FHq���pBCpH�L6-"���I��-��i��p��GЗ�D�iI�fg9��!�ÓM�3�/�׷$_���>~~^g����#����+��?g��mf=Kt#���0���"DUқ��[y�xx�$�t|kzƵv��Vn�toA[���6(����Wv����5�&Z��-���6�u3���;��1����ub��A-��'�����N/?a�""���d[��gw-Y��m1�kz����}ʑ���̯rU�j�ed��'�:�24��y��Eu�1�����\�آ7r4Һ8�5ScT�7�\C�5�AsG���1C��ߍ��s�z�!�Z��f�1ێ�W_؋3�����L[���T��P�C�Y��E��Y�ѥ�#��oa4o�գ#�Az	�nPff5-�C�Q�+�9��ۣ��(�6pW�����4�Q���F���r��������3�b6A���ҔT�ɩ��x���b�:��3�G��%Q3�{K�F��戜�8r�5/wc���y�����*�>�_@ ���y��ѯ/��~��3p?\݂/^���<�LE�g�����������&nw-C_nE��u^Ś��I��'K�{V�j�w�,�c?�r�\�2�/�Z޷5C| \�8�,��:��Y�In���9���������~wל�3��X���1�N�]p��w���o!��B~�g�w���-�^�!`�_ %��ƴqǝxfb�(�$�eV�<Kp��s��K��-y#����B�Z�7N���:�]��,�&s׮�w%�:n6�}@ˁ=p;�����sh%�MF�n�-n��!�T��#G<��{-�+���9/���a���x+E�a���}z:�g>H;<cͧ����;3��M�Y�a	h�{z����V����-�;š;?����>�e������	>����8'������~
��Eb��6��i#�!�}]քwa�ґ��&Yט+�B��9�/��lZ2�|f*ӭ�����H�����B��;��<���3��1ܔ�˒�N�[���+d�E�������1i'b�ܯ��n���K�^�t��MU�E�S�>^9��������Z�zmW׌r�����v��b7[[Fmf,į�s:�5YU�һ�ѷ�>���ra�%MRo[l����L�u��G��mI���Q= �=7�q�S1h5��¼<=��^o7�a[�w�wX{:�,�2�"U�ޑO'ȁ�3�83�^b�����-0�Gn*��f#e�S�ܫ�;�jc�@7���K�`���A�ow9j��'�Bos��꺫��,`�ލ��AҏGXJ�^�.���%�&�z_�z�w�0�j�6#�z��a�#�ܸ�ͷ�����F=��Y%&��~�Η�H������)󹎾ɵ�n�M8+=7q˷'Q"�#/����>��z�]z/�ltS,;�!�fꢺ�2�6/�1{�|x�����-�n��-�=ܩ�3�������vf��!8�a�"gϫ�έ;^�ZIQh�U9�]���rWT��Kh���7<ָ�zFG/i�\x�~Ⱦ�n�ksI��Me�t�#YO ���/�U�_M�Dn	��K��gk���s���i0v���8�*��\�9�+G'��֮�X��kГV9�'��>��$�߽�(����+�?&�㼁�ٻ�4t��)�6P��\�rq�"�#������T���|��:����&�O��G1�&s���v�q�W���z7(6��x7�q���"�]V�;9ӕXN�Xi��έ��9_�h,7���w��fP��/OdWR���z۾׀��yܖff�yBu���4����l�)t�u>�wn3y}��P8����=U��峢�[nf{���J�B�z�9���T{)���v]}�՗IT�3M3�o��6�~�ky�_*g�2��y�Ի�Y
lff�������vI�i�V^uNu�DÛ\Dȇh>��y{`N�+��l�-yZ��L�X	�=qK#���"
��1�n.��i^M=���ӻo�0`�P�3K9dٷ=kyl�&�������02}c:@7{Fo,ܱk6!OC��g.E��fê�՝���(�Z�Nh�W���~�9�u�g�t�0s�
�[�0<5��s꾝�g�PYo-K��°my���4�V(H �C��J|�;����O �3�
�|r�}��m�D�S�����&JK/s$�޾s�����\3=u�1���}7ߜ��x�����Tf��꠵틗�w	)ȳx�w��u����8޷��W:	�ڮ�����`�ll��˯A����Ϧ�F��1�Q��d��)�E��o-�&�/�y��/����x����+21��D�ì�Y�zݷ�㫊ZQ�>��8<���m>��&X]�C�=��w<{��)�L�r���&����Y6e��\�ϻa�٧�P|Tq�ٹ��8�a�����v6��:��j��:�]H�D��P��l�4r����,O��ף�f$Ѕ�>Ksh,�fi�����w��t�y�l�.r�No(,�������݆{�~�l�*pfm� e%C]sźs"�;�4Ql����>�zDnQ�h�ucBR��w1��fm��L��-�Om������)	>��~v�� ��x�uݬ�Y�� ���i�����.���v���{�13��DQ�]�b���g��E����<�*�ݶ��q,��3m[���N�9��g3�_Xz^)�U�ӵ��%
[q}Y׿:�"�ڽ�Dz] 7#sF�/��r�!������X�[{S�)J�qJ�쎙�li*�����չ�'?��#��x��0��[��-��!@$O����f'`\���l>���;����I�=��k���p Wnq��7�O�,k���q7��'3�|��@��y\q�g�����kbT��/iO�2;ѳq���YZ������q=kd
���X|�I\�󊩼����V�- NR����Fʑ�:����/ ���+���B�m�XR27b���;~ۭ�s S!����"8��D���˕���4'?��:o�e����D�mzf̌���wu��}�ܧ�&q�v�2���47{xl�<z �ނw@�"6z�� ��y�r¿_L0�����Ż������ݤ�#�O�??{5Q�6�6�]I�Y��)�����:��ȏ�k=2){�ի��ݐ1sk錈����L����xv���M\K*�>�������|H��U� ����w���u\U��G�x"8���Bm�ZS�Ϲ_I�Yy�ox��S�l��$c����6�Wd��>�oD�\�ٸwrod;����7��7��<�`f���_q1�`��'���ި$��[Xb�}�"�;�f��*���T*ݛU����=��|�[������r��u�j+!��6%u��-�W��Z�v��zg�q��r������}���	�?���p��4�7�ר��Kՠ���+���-���KIc;�=V`r�뗻�7�����,��)"��r���y������Ru�Ƿ}W�OM3�b��UQ�=�S��0�'��j�b̛7�G{h�hӵ�۴�R7�ё�Qj���n�������9�&����� zPe�p��8�'Ak�)W��oK�G��C�z���?�MS�٘z�~S��N�|u\d���w��Cc�z��f���\K��j�=��VO��15#��3�:��n����JA���y�j�4�5+���G��d��Rտ�/��3���s���F�W�N1����+Q؍�ECG��mN���X�o�2���e>͎���]7�$��du�����`Ps��f��ie�U��/��W�vS�t����G�����߷�ߴ�u��ǬUP�-��o����U���3���H5lw:_i��է;мJ�kg�VH��A�R�Cg_&�lnɯ���ODN�'�����xy��޿�:�c�!���i�������	�f���[�K=�f��>�����q*�\���~����$���� G���|\����q����e3S��J�芨���r�
fo3Du�������ޯsoezV�����M�ҳ6X3���M�̱��8Nzͽ��x�/=����t�d�%Q�O9#k`b�sw���R�u3WGW`���)�d�����G��{�H��B��Č����t[i���犳�������r;-���'��"ż���P$���n�!�2�-&hR���d���+u�T0e������fų�Œ�׺��a���W>RĮf�}V@�r��|MV�P���ZF��(��B[�6��6�k��]����]1��׵~-䷃�)���A�S�d���,�2.��X�ㄾ�qu�%J�s�HR�ˤ;S }w�V�N_1�1����xg~N��#�/��bxP��mӀK�3�E(�'����h}�[}wK��>�6֚pv��5���5���(J[O��"�D�����T��>��߅w��:[�^jM���\.̮Ϋ[�яw����Z�ŷ/n���U�J�}�m��bj�j����3���Cz:���dU��;ޗ��=��Ϊbr��dI�(鍻�� ��#��z�U�]��Ӡ$"y��Q�Y��3�
��g����j�Z�Ӝ�ED\���+�͛�<b搪eM�����XD	=�V޶��u^j�8d��_/w��W�Dn)�Ț>�*�e�?Z�)�W�Lbݻ(�_wn����n�lϙ6���;}��=z�~��(�n��L_vQ7b�s��o�M�3�n'�q>�3����\��wf��:c�}���Xf����If�[do�����v��ܥ�Ob#,̎�6Jɢ������}u���JE�]����G��d$�%f�lk=Qs���WL%`���}�Rw0P�:L��hv�t�.+2�7�*�-,�M�R����7�y�����a�9�;��{��v1�q�G@{&s�73�*���mm�Ue�MS�;�7�C3���1����Q`5r��6��)�d��zl�XQ��_�����<z5�y�-\o�:�R��2��-���4���н>�*c�I"C�������!���J�aq��������4�p���W�� �Q2b嗳���o�2��.E�7W0�I��5�Z.�^��O<Z]�P��}rqV�9�E�󭆆޷SxODøh�Iv��a~�D�Lz�8Β�I��R�[#�1�6�����+SbS^x�``Y�z�eO��x�㞛B�7�x.�f�D_��ӀuS���';�n�k,î�c���Uz�F��bu���Vw��n\�H	��{��{��?x'�Wt'����Xw�M.�a'೿i�)B��`:�{�n��^�i.CYͽ�mf����x6ҝb�fJ���K/��N��X]+��z�	x2�[���a�wI��ސޚ���'��a��{U��OVnj�뢈��:��I��iwe��{zU�mtW8spJ��6($��=b\ ��3�3�WKr�Q6u!�%e1x��!���ȅ�s�s�U�I{���˺�4����HnR����x-�!�쉘7�����d-֜�z���Mpzv�=I�(]�q6�y����N4ѓ9M���v�9@�-�5!2��K�ͭVÕ�h�׹���M�^�H��u�ө%��)��4�m����Y#fX��Ê�ꗜ�(�l bXE]fVu<ރy8����Џ(��Չ�AE��`+��#װE%�Gz�4,LgK��O7;��W:�cTK��ަ��)�/^=�����c�u���. ��CxE�e��Twc\U��ȩ!\�^)v��d��Y��ja���:ݽ�F��Z;�}{���c�K�Rς���-V<Y_Go��n���e[�R�
V�0N�;�=�.�p��X0ʪ���;�n�O	�D��	�bJSS���V)�D����f*
��c�����ФAԉ�J$�@�H[N*' ƀ�*��g
9n��@s,C�"0#uP�ԭ)�1v��I �hw�Aߑ��ʌl�0*�X�z�s=t�,5�ւd�'>]�w�wݏG'�y�B�T���Ήi���.q+K�Hw��}ӌ{w�-�1�g7)��{�֋�� .�#V�J�rY�T緩\��rk\m7���;��ڻ-�&�G��-���U�#k1����=��+{9#�N*�hG+%jT�r���)2��x�nq�IW-U$=��Co����ud��\;g���沍tm�	Ɨ2�����]Ls��%'��v4��^ooba�=|�6V���	�xܻA�Djݚ.����݋�'/MZ1�K�W�;K�j��H�����p��]+�@1��Q]�e���3V���YOi�(����1�*a��z�rԡdma��=\끳/�2��&��[Y���H��f\���7�82��p��+��x�/���T�9�k�Ӥj�U�Q�&�=.�/l"���ǚ)��zR}�!��}n���Y��؈�ƹ}�M	��T�x؅ם��۹ �l��oqekv�閜ζ�#��j���k^��RI�H����6:��"���ӻ�u��1=G֑"�C�d��5xo�z�9t��t%���]/k�H2$�8��oƾ5�Zֵ�k_Ƶ�k���~�a�$�L��L��,M���q�4��$fc ��������ֵ�kZ��5�k]u�]k������U����u����srK�6~n�<��\�9�������������5�kZֵ�kZֺ뮺�׾�p� dHB=G2o���u�u\��,W6��28��ƾ?��ѭkZֵ�hֵ�u�]u��}ܱ����+���kκ������F��wK�˝�:�wt�ӕ{뷫��+�F��3��'�Qbm�	$@ ��x>�c ������\8�'P�t��W�S΢�|j�պW��<��żh��˞{�w����1h��+Ɗ/ַy�齽"�w�;^-p�9�ۏ��c�˜�w]�D(��DbD��Q�L6�(�QD�|Zd6��I>"R'Ȅ)u��tЋr�<�5ы�؃Y�{��q\���)���פ����3�ʊ��)X�vu'0'��`�b��;�߽��Y���������+�����n6��M���wv���B|��^d�"r[>�D򱋛�Clt�zQ���|���v����F����PS��\�y�w�'ӞM���g>J�U:ȴ�K�5ɾ�D�"x`��:&9�s�t�N���[�4{��������W����Y���F	��~��Yf���W�������E��f��R��Q�̬�j,3ѻ(�:�a�7�8+�^�k���uy]�Q	k-�lXH,�}�wgfF��.���|+��pE�s��v��솺+6^j����qV��y�g"�Pd(�g��r�Wl�]F���(��3Ʀ{T��l[���%Bܷ��$���d^l���0��(�P�q�s�����������Igc4���ٽZ/��r�N_��D݇Bi�gt���X�ɑ�R�ay���[P,��O*=�Pj������n�4z忡_W�+L�7k[ݮ�&n&ju3:�<��$�-i䜲,ʚ��<�����/;Q͞��y��7���J�R6�Y�v�5�!Υ�33"0�y���S��`�H�6�uב�\�'k�yffͯh��A���B0�K�M�;����-f�P��b�q�4�Cq��H&���b[�+�<W����*@���ecG^
����v�p��p����U����ό���g����&��)����6��ӊ�~�R�)�(��d�{_�뎨���&vUz��,�q��C����9Pd����hj�[��[Oo���ql}�m$I�7�׾��l~ጆ[v6�7�En�\t�p��3����Vj�Gl�p��<���=�-�U�1����U�^u9��Nm�ǈ��M���E]�M� ��W�!y��z�����a����~��«�g���=�Qh�� Bս>��O)n���ђγa�SOfnqӚUb}q�n�*�N̚�f:�3��KZ�K�BI�3!�T�-J�P�I�q��1n"3l�1��{�.`ux񐐑'P�����ν.[��^��ԩu)\l/,=	����{��&�a9�=�t���2p��w�<|<<<<*���n�v��"L]"�ڰ��
�n��JA�fS�i�۵d�S�^{;��U�%8%tn�n�\�ዮ��0� 2�\��b�sϷ2S�`,���Ty�=Y&7S�Ue�^"��c�`8ډ����G��c+�} �X���2ea��eV����d�x��l���"�S�#9'3|��;2�!�E]ڮ�:�(M�����2�y���J�G���Tߝ^Ŀ_�9�z4������K�ͼ�y�j����>���nNcY�Q�Q�U5Ra�e�\�F7��1_$Q4�I33l��"F��nR�N�=�`!�b^gk	���7F��jS.1vw��i����x}��X@������㐮换l0�3�I�#���Z�}Y�M�[T1�I��Xt�s���'M�u}�v�r�~�zv�3S��̛��U�+Vvg����:�CV��fQ�Ҏ��g^�e`M4\��پ������v15Yf~�z�����O��i�9-xs�g���Ē|�ԳF�U:��mY��XO��M<���	7�����k�_�I-f�ېs�)��J�C��©	�]��2!�c��;d���/d����}��C¾��έ��g${R]Nl3����^z�y�`�v��`����T6���+��pߓ$z�W3;3��4�w�#�!��cG���9�4˵v��<P��� 8x�_]yL
�R6{:��y׍3�9�49�lƱDQcV�Ux0�\�b0!-�����i����EXTٞ�h%{*�C?�.��Z��G^RՂ��1P:zSg�m�t=�wm�g9������4�uj7u3=޾`Þ�#�H��.g�ݵr�|�������;�{�WWl՞oJ���ǈF��o��E���b�iwʹ����&���d�y��v�g��aa��������p��˗6�1��<���K��贷_��HtXhZޝ ��f, �w�`�M�F[N��"�wp�����k:��-���y��*ا/k���O��\�����6� m�ݧB.�魊�nm����.u<v#������1;�S��Gn������\%����3������u�/�>�����*�N�|�"�iGe9Y I������ª���>{+�s��kz&�%H��7��Ui���2�ќ�4޲Wk�2�Z�������V��nve�m{}q�Ri��֌���>��TmkWlT�I;Z����m��9�g:�� !�����U��'�3k3#�#�c��UIګ�^��V��8�T��q9/u���D��L�F�U-4�*�� -yF-���U$w��>��z�c�o+�Z_��j�U��cy�x�.�Y�ӧ�6�]A#ӆ̆�{��&e��L���;����������ּǉ̨[��1{�5_9;����ҋ��zB���N	n�q���A�캳��>�Tu�p�w~��d��s�Z&C�W�WJn����7���&f`�9�͘�h������s�����Ny^l6z��4/��N鈧;|��0�ϰ�r�3w(u��Ɗ��9q}��Z����>hɉ��'2iW�*���e����,����v����t\=h�&5�RR:��[�w�������K��v$Q�/l�l���p���y��j��+_����v#���׊���׋�k������4�n��QXL���@9~�Ke�H�D�
�>��U�g{2}Mw�W�v��4z�	�p�ڤ5��&��.�O�s����"�ԶQ8՜h)�3�d�x=!�U��f�{�;����n�k.ƝU���&`��N�K0Q(Zj�~����fk�gI$�,��Y�w5��x�Z������1d�����!�"a�4�O*�s��fΜ+d�3�sv��u`�܃^�9���ԣ�i���B)�p�����5"^��l5UȜ�J=�����"��%f���Q��Q�xms��b�z������۝�pq3���,�H<��)k��5ݑCGx7����İ�9�����d��;=)�6@�(L{��È�-���\&2��7�(9y�A嵒���z�Y~N����;��d�zB��	e�W��/W�H�,��GÈĚ����rí�.nL�]�V�}�uY�Y�.砧b��fcHl�mGÜ�ݯ߼|||||||@8����L�ϷpS8t�-L�We�p����&�	��Z����P˸�h�fU����s3X�2ut�2r�.���F��S��uO��u݄u�����P|~'����_�����D�LƦ]�v@vfn�F����DLp���8�T�\��j�N���l`�x�廧9��C�6@m�G�x�GM�s<���.���r񪏋N�4U��uBQU�֯n����R�#��h�R5�i���w��cW�}�Ñ�(���X�72Us�U�&��6��E��YERI�/��\p�:�t���7�M���v�:Xh�˘��ɫ$���;��B�ng�W�m�_~���!��؝r�*榸�v��oZw�5r�7ƴC��A�o�E�C7^h1�y�3K���Y��i�+�#r��[��ȱr�w7�b��,®nn�p	�����P��&��a��I�����I�_��Ԟ�+�?�1K;�� �Ub!��:�iD:ǫYM܊��Ң�,9��������6�d�������n��f|�C�ƭ1�
KnLKfs!�ڶU�eS�傖���7�X��R	��%u�<���ju���C��Ê�%bDWy�%�v�2�WFhq�ޓ�G��P`5����Y5�ƳQym@�s�S��S� Lj�Մ��Zܜ��Y'u"I�xfs�#��݁Lu�ϟ������Czrو�w2�[zO����TODǥ7r7}}�Uy>xFf0or��'P�4 [��o+����-�a%��� ��Y3�
�>�`����-�Y����ij�Dߛڷ6�aQ�Ӧ[g��u{M{["�C�3��[e����.%��?l"eo����}~K��ӫy��l�]e����D9��صG^��W�F�ai;��u��;ewt��U��Xf5S�S�7sZo{��(�p�y{�#w���ɜ�uy�#��&�e��(�ۺZ�+�rd*�<�u�>Às���������Y+D]E�n���4 ���].b�#���o"��q�k\�ŝ�|}�*�fc�t?|$���$zIv�'ǭ�0�B'���W����>s_I|;nA:'kTԵ������4或�mHN�a��4��Z�ݚ���y��o0���q���hV�6���xx��4���
������Gs���[�pd�mi������/��Y��o0�$ǆ\3��V����6�gCB�����TrW�Xn�7���BA ���om\4vN�c�=�KHUG�h`�����������qd8�e���&�b������w]��c����z�}~��԰���#�^yv�Ѭ3��<owR(�h	�2i�6Z�H���O^�6�W��zr�F`��Z|do����K��Fob�wvw�x��0V[�nj�=~�jј�?\) �h���^��Y�Ƿ��z̝�����8���S��ѕ�f]��JҦ1�4�wz�Y�*��R{���O��9�>�>�Q�Essqj����ΐ�wJz��~���ܷ<����Ѝ����ߚ4E�������R-��ۛr��e������-��&7\Wj�8�XĶ�����B6����QG��'}��y�W:��k'et당���Wwl%������{XbMg)Rم3�p�y��` o4<֘�*ڣ�p��6���zEH;��C%m�P������d�r�q�t뙸����_�P����rvk�����S໭����M�8%��C;?S�FqsB����o���~��ɺ�躑��6�����z������U�W�}�E�b�	{�#F���շ1����Ugf.3��5e|�;`\dW�F��%��B"�$�A�Gi�U��R!�zr�ʯvo������ex�)$��	��GŘK?Y���o��D8���6��c���@m�6Euv|�$I5��.��&{3xՊBf����7�F��������N��c�4�ہ�j�V�ޠq¢��4��3�@)C�'��L)���a�Xwvz�����@ۍ���:�hǰ���O��O�DU=�w���~��1�  *��"����{��(�AW�`��	�xp������;�֧��ܱ���5-�X���ŕ�Y�mT�f֘�f�MFkZcVҳjҬX�V��mS-��,�S32�1�mi�2֘���jL��͵f1�եXœ-�2d���I�kLe1�m+5���3Z�c�Y�c-Y�2�f2d�VV�k,�����,��,f�LX�VcRՙ�K&mY�3m�������*Ҭd�L��M�f՚�+i���j����e�2X��X�V�1�ZX�j�eS��+6Ԭզm�3kJ͵1�[MJ̶�f֕�jX�U�X�եejVj�SS-R�mJ�jVkYY�J͵+-�Z��VV��6����f�+6��֥eZV[R˺ݵ�jm�Y�Jʴ��J�ZVmiY��em+5iYkJԫJ��VU�f֕��YkJ�H 0����+�iY��f�++iYV��iYm�f�+-iY�JԫJʴ��ҳV��ZVU�eZVV�f���iV��Y��f�+-iYZ��ZVm���++iY�Jʴ�MjVjҲ�+-�Y��eZVU�f�+6����j[R�ڕ�ZVU�e�+5���Jʴ��J��V�ZVZҳV��m++R��+5iY��f�++iZ��Y�J��VU�f֕�iYm�f�+-���R�6�Vjҳ[Jʴ���f�+5���J�ڀ��Q�0Sq�uZ��-j���U�eU]��IZ���U*�mT�*�J���U�j�VP�s� x�� b���J�֪U�V�Vj�J��T�5j�Y��*ͭUݪݭZU�iVU�YkJ���eZU�ZU�ԫ6� ���!�T Q 6���Z�f֕fڕeZU��Vm�j,�]ڭڴ�%�iV[R�֥b�kJ�Z�e�-L�V�e�V�e�y�[�ԫ+R�YZ�em*��U�jX�6��*��եYm��*ͭ,YU����K�K5�2��Եef��kWX���FV�,�e���{_����>O���QQ	PDH�#����/�����A�O?O�����Y�?����.��p���L��������?������P ������������ ���DW�_�?�� t4�Q�����?� @U�w��A��?��� ������'����<�3�� �!��~�"��0��P�HH#ͭ-eZUJ�ԫM�+i[M�6m�kJ��V��mM��iM�+YmJ��֩Z�U��KT�V�U�$F �A��F����Q��F(� )&����SkM�Zk*�U���kKVj�*��V��U�ʴ��5��6kSfڕ�jiV����Z�j*�jU�ڙV��V�j[5���jmmMKV�V�DDE@_��@p�j�ړV�j*�Ul[QV���V�֋Z��JV��hڤ�L�M�ԥZ-�f�+5�MjjkSf�6��U���5M�6���U��R�j�Mmz��!	��?��p���h�����"H �H �H
"O���}���?�����>�W�����  *�N��=��������H~�7���G�ڝ�?Z�����֝�AW� ���h~�����I٧Q ^�@��P@U�@1?o���z�=���~t�~�]0��4 
�������~�?�������z�������y�`W�?xo�?h`�����C���DV�_�@P�i��;C�H�������?����:������ ���|�1�og�L@���?_p8��x�\K���(�/�``~=h
 ��_�7����b�?�1AY&SY���|R)ـpP��3'� bA���j��!RTP�)D���*�����
B
�"�R�RE(�(�H���*��T�(�DUJ$��P�A
�UU	IU*�Q'`e&�
J���T*���H�
�ET��($AQ
TD��HU*)$(�H�UR)h�����%R�TD���)*�B����U	BH�A"(���*!TJ@!R���II��)*T�B��Z���$S� �u��c���;7;�YT�mXh[.��VM��+j�-;��t��iMkj�[�Į�]��\��I�%*m�w8��(6ԑ�v�U	Ҫ���@�QA"�$�  
]��t�{d���KXc��ؽ����wc�k�:�o){i�5U��Gv����mV�h�M�k��hY��6�]�Zѻ�������9��WM�v�N�ۍeN�sGD��@�UR��
WY�  �T�\�շTҪ�h�L�m���;�t�Z�K�]�mgiY��j��l��.jwh�#u��a.�[GN�FP֝�]J	
IM�FH���P��  ��Р^�����mS�;�%wf���a�����Z��YQݡ�M���M.�R���٠`�;�;���U֚H)*D�'L�B�Ex   ��κJ��6��V,u�#`i�̣їl�v:wZ.Gv���������ww(cn�l�Sj�kfU�B�!T��� �J��   ��J��0� )���� �i�  ؘ@h0 � ��� R�  ��@uu�\ ��UPJ�*��D���   ���  VL  �  �mp� )e  # ��� :4;BƁ@��� 3)	P�U��!DH��  5�z :Z � AM��C1Y@ �w�����  UX X-@�vu8 �P�*��@ER��  ˀ ��u  ���  n !�  �L
 @�@ 1� ���)�)��� Dʒ�I�"�EBSx  8�   � 
�t�t�@S+(  m�8 Z  �G@@:l  Ύ x)�4�ʥR4#MhE=�	))S@  0�0&2i��JR��`  "y�*��@  ��)5U2 h�1??���~��'�?�����H�I j�uN��$ѐ�+6+8��vVq���}��W���wןo���ֶ�V�ګm���Z����Z������[kj����7�����U��d7�r���cͥ� 6½jM�(�f#X'�#hC ��Y��ѽ4 �/��5���΁��,7S(��j�kI����́�F�`݆]5�
���^iV��3 m�甁En^/�Ɗ������(լś2����C+"a+�7��	'd\��)0��x�c�@_�d�W�h̫�V�"5�:4����wB��X��Z�&�Am'�p�h�K�FPv/�, ���z^ݳ�	 ��o������J���N��d�v
J���5K�ͭ�.˻ov�1+���;Ui�2!0`DX��"��e�����VQE��z��Eֶj`ڧLL�E{����a��@J�zȨA�$�*鉈�����Rm��u��q��B��B�=Y�A�0f�úa-�;������ �B,�?KF,א����{v��N껅���Rq^*Lc�6��R;�^�[�5-�R�&V�6���.%�	a��c�����H�=���m�&L�X�i�4غFHTsi��[[ys1m6�<�E��1N2�f�(�A�j0�ɶ佔.��2��X�k[ʠ5�/Ӽݍ���#���.^V�[��Y��b|��;/r�l�V����\xZ�DI4h��P����E
�v�.�DKASf܃G�הp.�2nH� �,֋5r:cU՝85�V$Ь��!d9/[�M����/RQ�?d,��/Q`M��],�0� �	&	[�qJ@l��L�� -%\��$� �(�*dbk6Q�k�3v;:��tE޲���v�zaG���#�R�f��u�$�<�-�U�
JC���fZ�l,�4�{���&�Mhu�0�e�jU�t5�Ea$9���]�h�l, K��1e8����+"㰚Ѳ�7E^�qG�KJ;Y�k],�N��y0���X�v�)^k�6�˘�;u3cDXˑ�Ge
�vަ���n���/�/�5��gDK��l�2Ʀ`ք;���K-T��Ǆ���Kj�ҁݬ���pѡ�Wè6�Ǣj�C(.�5F"�S�TNSt$�f]Z1Ƃ�[���hA��7 ���U����3hk�ʈ�M��d��&˧��Ksje&E�vh�����P
M'j,��RS��I�-M���7����'�Vk[{��{3*(��Z�����E&?���6%�	�f��+��E�I�E�8AMZ7�k��u+��+��9r��lX�X�lhM�(������F1`dB��4nŬ�����y�� P��|�Z�[50il6e��1#*V
��B]�تM�F4��ү��E�mR��2A�
BMu���ċB;�@V�^�re��E	+��.`�2K}X�ߙ����x 	�ܬP��kH��ˋ,�Y�nJ�n�nǢc��3
��m ���V���ı�8��n�j�!�wN�M��t�3QT&�
�̀�V�L���+sZv��F8�e��)����Y���<�H`�M+I /P�3D�4K���-+�s+n���k�i�;˅�d��$�IKii��n�-[�
%�7nK��ϴ�R�Yo�`^^ �Z2�Jm����"�t��Y�aAwMf�:b��pKee8��W�:h
��
�P�b�Vv��*�������b�Ĉ�u�-zcÆU�KT�%<�q^Շ1��Y��Yhޤ�h�\YZY�cVp`0I�JѴ�/����u*h̡z*&i�r����5EZ��Z��d��4���{���JUn��jYd�n�F�S2��ƯhSGu� �v7DfՉ��^Z����f�)n�kb��
'.�˷�=v�OML�Gk�f�1ASn2B��Z�4�a�p���-f��k���)��B�������H�à:Tȱ�͌����o�`⑀�ЭV�kG£:��no*M�	QGXU�L�j�B��I(��C.�6wp��X�w�#�ީ�V��ujnJ����m�.�X�4�nQs"�
uy��0]*S]�UwG�ˈ�j�D�d�j�\b�:��X���ݩ�ԺK��H�p
V����&6�-�V�0(!�WV��ޛ�Xݭf�lR���k�ղX���sNV(�,�Pz۷ZQ�s\�֝�n7,�����(+Y��Rl�3���,m��ׅ[Ηb������@�U�K٨���ʺK[K%�gnw/TX�^ӛx@�V�j
�b�Ŧ;B^S��Ch��8��n�m��Gj��*� ��Vf��L�HUfS�״��r�-��Ym팊�&��5�H��;*��zph+��k����CB�+Vm���䨃2�2�HƵm�pV��a�5	V&���v�	dI��7J*�m����He&j݃Y{f�*�+p�4���c8�D��B�6��PGI!STk+v��P�pC���t���a3����l,�+K�,�(e��BA��t�7������@�,f�2�Qm"��L�-���t�l�kz��A\Ç��B�+f�P�h��m��Q�e����u�
�1j��W1�S(�KK�� ���d����ٺ�
2R��MX4�
��{E���ssv^�r���;b���ʚ�t��e�q�m�i�����F2�	ު+Q��V[�E���p$�x�Cb;yW�,��b[Jλہ]�j;�Y4�:r陳E�q͗�[��W,|�e<��;Kr+Ӵ
̢f&B�m��+Z��5�H$�1`����O�/sl],��ӬSA�����r�
�:V]�n����`*����3�u�::�ڵR�he�!X�!��2�͑����k�[e��*Aw�[�U��8�Ñ��ywlE�]ɔ֕�X	�s$�6�fEy��<���mK*؏4��v1��)���SV.���+{J��%�#��rc�a{e u#3W/RWw-��dP�6��٧�1���f���d�	�:��f�^ ��[�i0һ�����K`Meen&ꘆ�R+�	�ݕj0+�sfҀFh�wf��In;kr�w��r�-X��6��̢6���щu �zV5.��X��sM=���V���D9��*c/,P�i݃	{��ܭY�pi�b�x�ײL�� ���P�7bݡt7!�1�Vdw�L!�a�I����U:� Xs4�G)K5�g�*@@K,�:�Zxh5>y�������Q�h7��2ּ�f�R����2�駭;f�7�Tq�7��E�,�@���(5���܏ Ue����KJЦ�+b�g���1;(fhr�m�D�nY1���
�~� Z�2Roj�Y��7m6ա0Ggp�)�n����&�45qc[��sh�Su�)CI��T͘���ڻ��4ӌPL^V]'z�L�T�`�TL����W��Mc�i^Yvj=�[n�`�h��7of$ͬ��.���ZƂ����z�J[(���5�Y۔�B���t�5�L����tVV�okT&X.#Lahܳ���Q� ��PC���Z&{��ᘶ˘�� 2�İ�?����o$����՛0c��iD�s=̇6Q�Zb��\`jz&��]�*+�dU��G@�Jj��;����&���m���s*�.��ܪ��kY �nH��z�-d��%��e�B�Wك^���y�/FhJ�U�fbYB�IRLy�h�Z�D�f����Al���e%�?���F*�fĥ�t5
�C�P�$�ֻ��knʚ�E޷��r�԰nh2��T��˼�F��%:�f�z�!p���B�]YL��L�IS ͕��L��S���5�je�E�^���!�6�E��/CD��jT���az.|�YF�7��@ �x���Or�A�oۖ�o$ݡ1�~�Sp�A-uynBbX�sP���31m�rLlC-ʏr��{�Nwl�6�a��Y�r���p�*�"���fZ�V6]nu�h�J�j�cY%��[�[c[w����7 C�tqM��AL�d�S3S�^B�1h�RjA���K-bQ-�D4r�e앚Y��fր�j:nPW���E�m�6p��O#��n]����L]L]�Õ���S�X�L�!�<+n1C6��`�pF�	�N^ϬҨm9$aDZ6J�Ԕʼ�:u+
�-�z0E���WZ�d��u����cZWsU�#B�Ű�iTs���Ѻ;�X�����RT��G2��pAb�o 81̭Xց�Y�h8ܦ�[A^3SK�Ef��U��UA+�,�:.˃m�N���^3��>�K���ێܨla=/fz7[8+i5Kh�&���FV+E�d����PѲX�f�gf��năH��S�T��)���0E!WY-�
��Ame�1C��qcܖ��vM�M@�X�[���K�om0�Ԧb;�@Ȓ4�M/U:-��d��Y%
̬YJȢ���%{HŚܡ��&�Yf�1�9�ŗ�pQj<2���ѽ��8BY�Ֆ��e)�J4ˌ�d��Vi+�iI�te-�B�L�l�̺V��
z�śMB�O0]�şn-A���EhY�lIri�:ohT i��z�\b��{r�CM��7{6:K2,JUo��l �ITͭh��&�5^V�@��n��n�����r,�2I�X.�^k��ݴ�o4P)�-hP��4]��(	����5�#��-:JQ�	M�v��YH�����t1��r�{y1EJ7n�{��
�v��n�vDj�`����D��榝� rK1�+%Ʊ�"�=�B��1�)�ѩc�jf,�{csiJ�h�Bٖ������5pPm����n��4-��)�-J(@4`)!WXe"�N&q?�ù�x�+$�Wv[��cG"ϕ�V�a�����wMn�a�[��2S%��c#4ʽ��f�+�l�oYb�v���QfT�^lY�33*�7S�x^���$�ya7�[�ߣ�Q5��(b��]:���ed�gf4��4H���$�Mc�"���f�H�TrRME���e�BŲ�7.��2+z ���t���/$�F5���Z�cSح(-�	t�z��1�&��2��6��#C�CwB�j�2V�l]�H�ͥ!�h�`��ܭ�����Z�uos]L��[a-��"��8�I��ҍ�Z[�{![�������#���☓�X����ҥ���DJ;Q��PI�+�t\����;�M�4�P%��FǊ�#���Ūgh1�.�e����m��f�&�Gu)����fQ�/i5m�Z@ܽyM�h�R}u�P3��/��c0��v�(�6���j�xsQ,��l8���An(�k!�V� [e�l�0\�ͬJ��A�U��wТ�(/Nkц
��Mh�V����lȖ�*���i㴛@��f�
L���ٰ���4�&
��-m�&k�{I���`�@�XkLPO���	�KjLzI��Ŧdu1Rp����d� x��,Ҿ��E���p�Q����85ۓéh��fKÚ���S����r((�SQ�I(�
�+ׅ��]�sR�{9OKI,�[�I[Yf�IV�H�.n��gh̨���Ar���E֢JV9c�*%B�&����s�0v�9���E��mVM��L+HP�@V�@VT�Su��5W�ص���a�m슎���P)wJ�/D��*f61�ԃD����[vu ��2]:�p��̎��4���2� E�C�T�D�@�T�*l��m���bۃ ���PY�&��.��:˕(f	��p��)�33d�����1���ֺ()��riLCu���|�VըpS�(�6�ְ+6����yI��R�i�/v\�QR��*���`��r�Eح6�.+m�M(�Nva�T܀�ĥ���)Ģ4ՋD�aj�������^֪"�`&"�J�laӦ�ɴ���-��]cYj�n���u�PO�(/�B=�fƬ�49z­N��H���3&;q(�T�3B`U�Q��;��#���2���X�{*��$ۤ�֜�M��҂���|�`Ԭ�����B�Mۨm,�t�m�EF�����w$����7n��g/pB
J�u�� �P�sj�kf���Q�[�(�S�	!Zm�(��m!�bYxdyvN���,*�f	O%2\��0�e���ލ���&�����
İ��������h�//Z��Ѣ��WO �gB����%)�w6�Ӷ���ֻm�,�U>��j]�eDlO�JV�EN�ؔPkG6����/즀Y�ѫ���L�n�a)h��m<�-��F�K���m��j'YY+S��Ko�K
�Z�X/T�3��h�2��b�ܡbRR�4ж��>;�'���V�V�:6�t 1�q��
M�maUp��*]�	:�R���I�r��J�0�!1�w�Tt��ϰC�%��e��X�![V�6��XV5�K-��WM��,�(ab��	F�����v�J��3�xj=9�Y��aC�/X�bn�Su�y&k���7-&M�/%MˈԉZq��$�m�D@l�YY�A�b�eL��,��<�4	�Un%"�Y���WX�b�Q�"K˃G�)ei�f��P��5�p�D+�&m�P�3uZ�A�V�AZ�/��@+n�=�������6�*T��e�u��K^��j6,	�Q+#4��wnїf�맬8չ$w��zUfC����+r�{mP�QC6�0�j�c�`�t�6�,j޸J����(�wYzV�%&6JG(+�gHQ��̀Y:��@`��NjeS�K�X[�l���yImY��4��oR�jڛj�d��]<ݙ0��
q���v���c'w7pI��u�m����VAԕ�ѩ��S�����|���V����S�8���z�����'�ĥ:N�&m�d fjw3�wR�=�+��`扆�w]Yl��"Sij\6��Ƹy_�3M����Z ���H+�K̍4��ϯ�n�*�o\y�'Rv͇S�y��.��@��#
�cwg�v�q%����kb����/��9�����;8���<v���a�k&ћc/M';����}s�y�㚞f��HU� �4��>��r�T�n�q��:�+6汵��͠	��I��u٥Y�Eu��+nK�k��XA�$,#(Χ�N�O�,�"�%�M��ܖ���3���x�xx��ԫ�ioYv���ˁvĄ�|�ޅa�jԭ8��t�.ۮr�tT��������z*�VV�y��̦^ݬwxb"��ɍ	�����C]��T��v�'��͠M,\C�諾̌�G�HNS!U/7�t�-�h�})�\�y�曻��c�)�*;H�j����7�c����l���;��4\W�a���:?�ں7
�:���\w�u�D�e�,k"�L�p����ڛ3y=�Vwt���(�$w�]��;�52�Ph$�@�W
k�D�C�%�o8�S�e��^k��-�+{�zyX�Ϻ@�_`��.�J� ��Ws����[	�H����Morxv!ڂ�qju���v^v�?;�F�W�v�2����Z�|�_w{����-�M�wՋ��z{[���\k�2��T���A���Q��Z�˙z'>��+i+��9��:���k�t#nK��*4ي�����tsV��*ڧcS.�i�v����r��b�.v��xH���r��u�7Z�-W����ˠ�M�{`
�C]� �}6��H�4�s������D���P�د#��Ϩ��xncR�M��;mf��ΣJ��uv�[Ru\"1����N�PZ�"@WMW�e<\3����?ޣ٘��I;l`>�W��-���G���&*]G@�����To���(��\�p��l��EiL����U�,ҋ*�i�W<D�&&�T�W;�݊R�@a����,.�4�j�����2��J������/q�{M� ΓV�7�9Gg�ԭ�0���Kk�Z�zi�H`�?>��Od��-��uX����-�S)���C�>�4�d�$t�olj�����%fwuf,U�w7��af�:������m9.��dK���+��;�}1��w}�RN���� �{5��l�ۼ��v����Z��PB�;�u� �6:��N�q��h���}o��:d��uM}��p�8���-�*����_grү��D�Z����ދ�9u�E��r���)\�:��&.���K�W�v���h=�b��p��4�Y����ϔx�b�B���3�k�j��.��Xś̲��J��Q�h�P��y��pY}Op-S+J���$7�)���6�dYEI*��6X���0;���>��kdVZQ�Q�gy%��j6�#��E��{*��v��V�7Z� ]7MҺ��n���Fu�H�v�[���e�h�C�Gn����\���ց�{��XZ�b�k ��Uf��9_G�wma�y�OH�Eh+��S��V�Mek}C8��cY�dɼ775�w�4D��i�m��V�e�rN����Ug	n�Ϲ���`nM�wE�Ȭ��v,<`Z��D�ܾ@J��W0+���ѧ3:������Y��w����MIȥ3T:X:��u`V8FwN4gu�[ݧ��MG����;�f�M�\���^!��\[]"���J�WK������S�**�ݙ��u�:t	N�q�\8�@�����i�4��b"��$�U�^�譼�u�a�qMN�*+߯i�;�Y�db�6�-�\�h�]��Ir�M�*]��Bë��n�N�v)�%�v����:rEOf�]��Y9�8��`�'����i�
����Y8�R��w@�/�F�?-w�-�ٜ5w0]�Y ���ue�xn�������뛽��M��v�ܑ��4t��Tbb��^Aw��CF�I{O��:�~P�޾��7��Z�1�޹���j͚�Β%I��o G�J�j�:kUt\��\���lр��9��s�K�.�d��}�����fu���44�π����O��U�-�*���{��Z�c^����fnD[�g�����P�u6�q�
1�w���;^=+k:5X���nF�.T)<�f������[���Y�ZB��]�X�zZ�{��n�� �ѻ+�����n�[��7p�P�]|�]�K���G�6M�qZG�:��VG֨r�gI����$�۔��Nz{{.i�k����Ok6�|7`�b!�ⴵ��
���<�/,�s��Ov�޹R+�9���{4�"yq0�սϐ��k딷n L�o�䳃�zܪY���Y��oLc��x�^��Ex���_l�ٛn^��3�Ov���˸F���ˌ�@�=�;}����]e�}6Hh���c8�`�ǿm��@����G���TƸ6�P���S����V�.��Y)��_:f�|��֪i��b��\5��,Z��ޫ�G��b�B�0�k78�Qr��.9\A���`�ֲ���l:lQ����(��9�c�{�jjS�F�=X�,X+�O��P[�fb����NV..�D�-���97���ͻ�]t0���]Y�F��j��!p�ݐ�|h ������!n��^�]��T�a��^Wi�mT	�hj�Fij;�0�ݝd56b���L��C�Ge.�G�������Zz��ٜS��B�f,�1�����z;�ЛT����#h(�����H�@�*;Ճ�c��<|࣭^vΡy�f�F���� ;t� �vC�Z�
b�l��"UG��Ժ:�/��:E���ǃ��ܩ���V�+�S��K<޾=��i7C���"Ǵ y{�.�0h|2|0w
�"�ql�Sk�).+wr��6��k#ں&
s;
�x�§M�"���%���'cR��0�|��\�r�%���%sxѽ�2�����;��X��y}�]�_e5q�ڗQR�;wr�N��,�fL�s[�q,T�=qޫ�7|g@�.<	=�Js>x��dJ�������s�*)�٨:F��EcWd��o.��:]b��`�x�
S�Fc��\�e��ဋ�)�(����]L�1'v�csa6�u���l��{Y�M�
�k
�B�]]y�.���ʛ[����[f���]�ܔ(������K�Q8R7�q�KNkN�n�5i9ͤk��ݷ�M޷/�qqYN�KīJ�l���ޭ,�+����4t�u��f'��6�]��R��ǭq�`'��Z���[F�[:��0Mx���qks8�����Q�ۿv��@�Uy�6�ZV��fJy�B�ȬfŽ��K-L���G6fն�Qa �[ә��{���Q����L��[i�&�ZJn��[]]��Q5��������␵��D��+��X��ͻ�����83F)���K
n=��]'�TM�ىːzU��oJ�ŮE=��'*��kk��1[{�6U�����c�bIn�cw���#�j��Y���u�m�+�>��Oz�gwR-ݮ#�8�v(�w��Uۓ���F�$/E[��j8{�=��4R��-F&DNY[�9��-�s����z�����k.V�\��ĞdV˺o�Q�I��NӮL;LZ�=�M��}k\��%n�mVh�������X����� �]X,E@�:����qc&���ff�_;n��M\]���-v��e����\Pc�3���"��wMc}Q�l���R����TW��&ҭ���)�c�muбA�%�j�xI�l����&�e9�h�@:rN����ʅH0��v՗@�b&'����0�h��A�
Y.�1-0g��e]�r��5 ��d��.�s�l�Eu�O�N3�-d6��>�iZ뵠�u�Im�c��f�]K��Ҵ���C�B��W\��|GbN��v�:k�8�e���W]�Ȯ���-�*+r�]��P�sU�.����
��ܡa��ˋ����;ug7�]���ۦF�JE{�Y�@����l�]	Ԃ�u�Y�-,L���4�(V��r���L�_ݔ�AQ��\8���2��%r�G���q��������U���Ia_��0�3��SΡMR1����th3�]���r�����
.*�W\��=`4r�iq��|S�F����f�'J�:��e�1�5��N�]B)��;���)��O[*����S������#,�p,TԦ7�7�iӝ��<5αl��G)��e�U��V��-;p�o�Tܳ���dI���y����Xw1�)u٥�>�@U����Ⱦ�����I�xB���頮6�{��|��֍�M5{wyJ^1"�` ��&0��W�Wom��Cg,Z�ۧ}P�[]�L5[�	�Bi'�V�곓鮼T5	��vl���C��H���b�9�Mm�j�ѥw��	��E+�9��T�X)�ʳ#��b�:�i��]R�d*kŝs�`�z��"�S�.R,I��K�@���t
9L,y�5 S����7Y]�yQERn%�V�rA��@{4���wy��g��9sǪ&�hp=����W�k�wV��)=���
��P�jd����b��ŵul�s#��mR?a�`�m���[���`*�Q����ƈ �K|VX�;���;����fAP�)qn�W�٧f����Z�Q]����S�b�}�(K���Gn�\��Z��_B�k1���8��D6�N:{�������le�0M����U;�C/1��q=�lG�6Ϊ#H�U�� W�W4��
���t�)̶��N�E/�	�+��$�{�;�h�m�.�6�ѽoM����)��.���$�k�F�df[ܔw,R16�XӼ $(\;������چq�*��)��5�i|��Di�E��1�N�a5|�e��s� �VG��ӜB��}Ǒ�)U��Á�j�ݚ�%r	�R
��j�w
��n*���p�*h��D�}��eb*��>�o�7��RZ�^8EO�|9ed��@�/tͷӀ].���u�����-ʮ8��5���U��9#+jl��dv�uΘ/W̌���9�!��Z�W#��Ү�X�;2�G�\Ajl��V�b$�=�S�T3�v��BT^�[� ur�L��m��#��}BI�`�2��&�5���Ln%]P{��q���9��̄=������[N�?�ZsP�W	:�����t�����(�Goo��d³f�
Ve"V�x�iY#a����jc�u�G�Q�@�:���ɢ��"B�A���f#5a��*Ù�l�+4�x����;;Er--��#v,@cb��P��1��܁jvm���Y��(1�i�w�3Z!뷺&�:oV���*�Ǉ3rY��\U@i�z�Pp>䁾�g�U��pBl�ׂ��/���G[���n4U��Nej�3���;��ǣ�F��78��Pʁd�Gυ�aԠ�l�A�������8�P.(V[B��u�Ց1j]_ZZ���+w����%�{j�o?�S޾豗>�67���84n�Fq◺�p,��m_�MV���{��-̾�­'�q�諓gJ/�-1��o�ܩ��-�lr�0ժi{ˎj(�i���������8��=Rh�u*��]�L�wΣ���]>�c���@�FM����76S��R��t�\�6��S�l��-(v��_W3������!ӎ�Ӣt�{�����evs�v��L�:Ӧv0�87X�φNZo1h+��1�Ӗ+��[Ý�3#܂�%P��wCL�G����y�����mLq�m��P�ss�=�)�[���,�5�V�ކf(���;���V~ÕoZ:k�%�n�����9�bH�9ܺ�sgK�ε�'F��4:��}�xxf�96Ҷ�S��P�;IK�WvWl����1��7���J]I��r�{�k�EV���ڍY���OAfag��շ��K9�d�O0�l��b�����F��8n�Q6iWj��hGv�ܙf���哦i�*~��K�;�$6f�k�E'	��euc֏�ap���,5ȹ��&��]|�&��L��n_��{VS�b(lkg��g�{K�R�h�*I��⻌�����`t�2��:oJ��z�����ȩ�t�ta�Z�g7��2r
�\���-wJw��N���)����O^-Wy=�ca ��e�euty�w�$o��	�.�]�8�x����]e��A]��,rv0
�x�WhF$��;���T��˩}]����y�F�[ȡ��݄+���6���86�	!iA�8�X��6�Jݧ�s2��kPs��;-�<7M(gr_'HK*At��w]�޼�n�!�ypںQ��������>�ǹ�°�"N9����\s�����"��Q�!Uσ�
��yQ���\P���o�b�::�c���j��,M���+c�m�b�+;�#:�^me>Z�̉S���Ζª}%�k����C�8xڢ���n�6�l��Uh�����6��Yk�e���عϓW������Z(���ά�݌C�k�`�".�7�N�-�W�g9�zJ"$�
5Է �9����9%�gc��*�4�x�ӕ���r9f�����w'm����M;px;n���ń81����&u^�+�q��}ҵ�p�M�'��k�@��&�-�J����>��ű�R��2���3�U2a�'WC����\1V�͑A�Oe�.�Hb���(Z��<��费r��hy���Wv��oPx�y_M�1U�%4j�pg��e�<�U�t��*�	��V�j�#�K��^i\�>˫����b�s�M����Cio��m^�����`�JJ�A�C��j�%35\�|s9VD�8F���1Wl�Fv�e+\��L�����{��!Ӹws�����ٲ�o��i���:��gN�������U_}��꯾��������M�3�[�>�:ӡ�('��yv^�S��f�tk����v�H\����w]v=&��f�t��XN"��ml��������pMd�wg���9��S^]5���ka<]w��*w�O�9,�Ǭe�D������}V.�['�!\��YVK��$��L6�R���uݶ�Ǝ�͍�1�͞������
(�Ī!m��i�%��!��9;E˸X��olSm�E�+ךg|[�d��
�e�=ºѝ �&a�?KѠ|��D�ƛ��b�V�7k���]6��y�4Ơ��*Tu�&õ�C%mԃ���V������`��e�v��5���O���Y�u��yTpq���s>ڋ{Wnd�v�]Y�Y<��ԭT��ӵ�\8��]�\ھ\�`��[���#[�ӵ�0����Q�7}�D����삶��0�N�j�U�L&��b�����Sr=Iz�n�m-��a�l@͎��s%)�J��c��c�x�E�D��t�r|R32p��,�/cޱ������eaz!��w�29<�Ҵ�|e�Ջ#<���L�� '��Æ��=������˝�����"���j�����vN�e���ZHK�fc�r�+�C��,�{��;ik�Ƙ�ǯ����ilQκ]�Z�ݷ]���l��p*�r	t�KR�2�`�F�P�m��˒�v�\�F�]��=y�ϋ��h�'l���\z0�՟D��k�9X�%�t�9�Z2�[������6l�	g��'�v��b��y�q�1s*�C�,�{ƶֶ�\�f�Zͳ;*�q �,;�9�rG��P8x�a�wW�l��S�;@� �h�wpY�S:ͥ���;|��Ξ��S�]]�l����H�_$�+����]�GU�ݤ��D�-��ac�5��#p�7�[���-�-h-^:�Χ��� ��u��e���;�4�P�E�n��Q�a�<���yV��p�%eٳ��3��V�(4E L�Е�x,Y�[bl���kj��9]��>���#J�Uh<�O�P �:�":�19���]мÊq�����Y� �X�,_X|�]gR��9��{���	�����FT��捥EG4��G�W�����J��u��-���v��D��b5)�`eڜ��ݰ�C�(�X��,$�s�ʓV٬�ͩ"�S��YF*Ÿ��m^�K:Gu.��7�I�mhU�^s��˻8s���A�=DgC��'�6�+�]\���\�΃tv���@���
,���N��wՕ��=�VI¹�u�_sQ�, �f��b	�����YW�-S]�}G�,����ὯVwb�H��ﱴ�on.�ҹE,[�"˲�F�I��(Z�í�5ѡ�v�gp��#Tx����9/�uY��'7Z�J7#^Wz�T�H%��W�,�6�19w�2-���n����KJ��¤+T�f��뀔���z���rFIq*����^�0b��%��l��iu���hnꢮcxI��t�gHs�2���6�д�J+��ԩ^�T�.���y�bI�*��b�ɉm��oyl9��fm�!��_s�e^XL<�\��޲I6ՓV�u�\4�ѳ��*ьF��W�*����7���қAҢr�����e�Ӎ ����CdV������p�\/��)�.n*(����ڻg]���)�wS���i�-�����_Y��;,���j�� 7(%��;��Y�Ky%V�ܣo�B���X��]�8��]��W)�)Z4������ ����q�(#���!�ld�l��am�6�|�+%+ZZB���(h��}Z�۳0�[H��_ʢɆQ;*D\7@H%C�]0�a{B��(;r���� ����lVk5Z�qw%O�e����Ŭc.����9u%�]����՜ͲuT����NK8�r��4FZ%�B�bW�ظΫ�qv�2Wj�z��ɻ��f6�1Y�G*�h#Mq{|z�S亵܇���>Cpe���@o(�]��qt����|���W[�C�j�U�T/&k8���Ӝ�4;�oX�Ά�B�77��-P�jW�^��)�}������E[�b=����A�g�G�:�]�W-��E�=WW�WD��M�U�M����Ƿ�DW>��<���aT�ӈ��2���Z�t4+D�蚁�^���k8����ٹ��I^�z&��	#Žy����m�#Y�7���z���pWV�{��%m�G�:�[$&�]�Ҍyf�3��r�ܗgP��7����|6.�P[ǲ^��{t�-a�uj)K�T��װm�
����W���u����9y7Q���QY��'��JP�J��vzK�]w�	�-��0�K��I˫Fa�].(	��m!��k$5����s�=]T���^��ۏ���SKl֫TZ�x^���j�y�R^�(;�-�V.H�2e���#p�9:���د1��n"�Nt�%���p��uw��j��\�sr��T @Y�[!:�OCC��-��0�WVu�5���Q({��&��&2�%�t�:�|9�K���!���zjQ׻5�z��f�j�s�\��l�����ԥs�����4p��\�\Vf��c�eY�(MX��\o�r�a���/�(gQ9�S���2��9ԴnT[�4�*ι\ݰ��
se�z)�2��Sy⮫Ν�I�edj�|�J�m i����5��S[B�ƍ�:�q�6��w72.�H|"p�x�f�+�Bq�X	T����e��&����7�OQ�2���/�
��a�&�����SE\���ᬉ�fV�M��YK�K�Q���έ*�uwJֲ�ga�G\i�#q�M�:sv��w`e���% ���tk7;�ۮ6w�Lm�c^]�H���&I��k����S@O��n�Ȳl��nPmh�)p������.i�c�'.ޠS���*��i�j�?aHV�.�J���桉�vY�Ʒ�З�bv*�8ɺ�2oXK&顇�:�YH��W6ݫީfKt*�4��\S�3���Px2�v�+J���(ls �LDq��t��t�����]�:��[(���R�����{k����UkK(B���7��	!Nd��(��(qF��*���K�7��L�V�|e
.�/e�:l.��;���B������81\(A���S�5�s���Sz��5���ހ�4�b��o4�yt��Pq�M͕&1K �b���.�f��Bx�ݐ��=u�
<.��6X�lJY6��I�E��(�苦�M"W�]DV���W�@�ً1=��.E�N�6���W˶frC�#\x�}�)j�t�n��dn��r��Y{|�T��[�}�#�u�ͱ�6N���u�;�[F�L�Q�u)��@�Cp+WS�[o���	ݫSRYQa�9X20+�:[�aF5�n��J����&�mI����ǂB8%�T,�k�@s���V���k��D�O9��y,�V[3�j����ri..��S͂�u�)S�/wp�� =����lբ\�.7���V��8�\[�3C#s�m�'���L��v�:
&�oAyY��=����-�y&@�zv�⮣�mU�kt���u"ݣG'�6�J�*<J��:�Hr�,�^�s@5e�f4s/8.�zoV]�l`���wX�\t�Wv�+g:�o^�
�yc�����&ˣ+qG��\�9��p&Ef��:��5�4"�󹍴�Sn����ts�*Um^��^ �x�]Ԟ�+npj���;[�fN�݁��I�������;�+#nQ�H+&�+�^�Ψ�a� 505�P��X���E�ܥ����D7Gn���f�J�3)]]�f��X;Wl���ʘ� �~4�B�^�0���eΥ���2��P ��H�CC1l���_b�vT�܂qѦ�k ���h��[�Mq1��FR�Ʒ���L���":�1t�]�8�j��	�:3+2�#���ʘ ����\��&�^=uv~%��.M-�7�#D�%d�v�%Ά^�l'�Ca.:�|%�l�Qd`퐷Q���֙���m��Z�7t�.B�l��ZV��7wĤ���:�㍢k�nӼ�͊����yS84�g�}����:��Q�OM �խ�2�f�m%�e�K�x�D���[���w|��>�wN=dU�"��jg���Vm�Zĥ�Å$��ڳ+^S-8���}�X]٩�z�mi��ȕ�+�wdc�E�o�eЫ����V�.E��n�+�X�RԷ+��� M
�K.�1t�i��J'�� �X �����Xp�O-8���[&�<7@�q������u��TG���у�R�)o2�q0:��gN`���N���U��rv����fA�Y5<<T�"�m-�0��"8�2n�P��)��d� �ڎ*��1�s�jʫ[��3�鬌VČK�8O
	j��s��rử�%-l�Ћ\id���-'3��)m�M�1蘡����*�"�w���W݊�3A��t5��a�Kr'l͊}ˠ � �B�*� �����]��M-h�l�(�'��Ix�T�k��N�7m��Cd�6�b�-l��H(�_P�uצѫ��_4����<�pZ�7һ�LS�%8�5d=��u�w�*d����W4C���j]��Bޡz��/��$/��-�gf�<�D���ZCX�r���l4�R�[�M'#e��T�Ű��.��⏋�z6�M����d�æ��3��<\�Ŏۙ�i8mB�s	�;�a�Sz-�Aҽ�'f�A�E�D֕<�".�J��-8�y	wz�)��^,�{538T���ܬ�O>љ�D�0F����ʕt�ӫ�}xj��r�Nu�f�{�*�Nj�^�m^�Np���h��2jZd��5�C�]X]}4"��G]N�fo8��fo:Ѹ2FzBV�F��{f[�]�R_k��������*]J�({{r���o��w��Ʌ��xuH�G/w&�+	�n��](��>�[��`�!
���
:�eT�֩:�<D�5ya8-�n uC�a�f]��I��k����^��{D T��2̂[u��H��g#��L��Y��0�j��F=٪�	��ܑ�ot�A�U���8�w2��֓.g7�mh��a8�
�u�v(ۧy%")KGY`���-���4�������0�k��ٜ ��,�� ����T��;�d��1\���6�e
�u��rW{�4ݡ� H���5"7�k�,Rr��t�]���x1���]��mm:ݴ��U�F�Hmk�7�N2����6��gom�|����ed�{3�e�A��X9�`������9�E>h�1c[Gs��;�{����\�ε��J�a���;�ʖa��h��l�Z�e��o_Y��o`+b�m_+c���j��B����6!2�m��a�Aƅ��R�.��{�Ed�éR��J�NA�C�:M��B�%�p�Ndi����m4��{��	�r�yZ���x��}XV)v3&w����
9sq�M�5v�Ձ�T�Nt+9�\U��<���삯�]�|��{��@��Ze�@��}!y�;_)�1<�%�Ƒ�Z�wA�&�T��7:�1�Å��8��`r��s7�(�.[�����b ���x���Y������ޫ�=SK�4����c-��t��XLڻ�P�*.�t��+�uL�G5��ѽ�Q��J4���(K�h�[w}ė-�w�e��y���ڙ�q���ػ6���LT�`Y�O��N#[�7�#�u ӕ']e����Ú��H�rm �͚���r\)��p�!tu��oe����Ciޭ��q�qb|�t�����֨�._8�f�k�8���wm#dvV�"5�n޻mZQ��}ɀ��3�s܊�ľfm�XA{�m���r��:*�N�f ���]7��i΀N���ގ�@�X��o�u��vՠ�w͵�@+��zy	F�q� �{�.ɇ��d��i���-r��t�ս�W=�o/�W���aV〲��S�9ii��W�ܮ���-+VV5h�CT�`�A�LS���]F��1��vVޒZ�wJ�^q��e^��ʓJ,�&���i����Ч�E�q��BR~ٺ��}��w)܅r��ų���ȹ47��`m� �v���wMJOJZN�Ϥksq����;5�OpI:���/3E�E���d-X%`��c1��z��+Z��sVd��y��X�®j�����z���@iiA��Yn���`�"� 	��Q�d���b��3vՋj�P�jd�(��>�A��|�V)ȭ�N��8���n�Y3+UԔN5,��6��Ko�!L���`8v$�ɝ[R=��wq-<]gh5#�w:p��*V�[z�}l����ĳ��kM�3!�ں&�zuЭ��Ÿ��K�p�G;-�QE�ɝ3��0��T��لT.������c�Y�I�f�����Z��;	��4-q�asfɜwx'}��9г����w؁Lt�3V����+M>�M���!i�KUlQ�s:U��κ���C��f7���|8��WuF��f��v��cŻ�;pt���+c������N���>�	�T���l�>E�+��Z��S��a�o�s��f�j�β�qu��h��r��F��ː'������g�f��6L{�9MQR��e#h	�������z�D�Tׂ�С`УS�5�G��5;�!�5d��;�f���ϲ�c{��z�*�U��^�M��\�	�K��߭W�a��`l�L\�1��<����;0�$㚙��}o�.���k/N��d4�*t�����-�K|)VA�wtP�<(��}w;�U��K�Y�����%�z��`D��coLaEfJ��G��G���,k��&R��`^q��܋��A��Q�&v:n,Ι�0Vb��dꦱ=��ww.�J�N�Eu\��gY�T��z=�����g��s#�)��nQ�`�`�a��L��A�"��Xu�B7A��u����IJ��u����y�nϻ�r��S�4�Merf��{qHa Z�mf�Ӹ���b�E�Xp������Q�d*���n=���':vج�f����F�]�m��J�ь���wG�.:���#Z�1ձ;�3azp����\z�� (-�K�֣�:�v���L�Kv:����Q�kx�"�׼w�1r��6�%���Qa���"�}BeL�ٻYb���u}�vote��'\�4O��<Z��[Z�L����y��͘�>}ܲ�b��MU���iFT� �v�S��R�L,,�0���V���\�R��n�E��"@���a|��);��̎���fL���$�-�+*>���9���9���Aگc�%�݋]�!&a����5���bI��G�t#C+z�,AZȜ�L�.�-oC�V���32�M�y��V����l}y��9�	�፦
S&5Jq׵wǅ�aiۗ�}�X��mnmЃ3���e䇹7�$��������l�70��h8D��T��6OwbVV�VWaԅ�+�k���ܳ3�:�F��=g%��b�a�ZU�s�����h�zRR����=y�������M�Q5��s�9�α��4A]��ڏ��ε�1�W*�\���9vr�Ryݢ,lȇ�WB1�sc�3���\wUҮ�+�L�cEp�����ם��W-���͋y��s�k���\��5s��͍Α�],WK�7,Pc]�o%��m7v�M�Qd�wcE�rѮl�w�]x��)nWN]ݭ�9p�˚���ۖ��;^6�W�ú1����Ȏ�����m�u�ܰ�s�scstǋn[�\�幻����r.F�nQQ���{��������ƶ���.��-�|&M,���ȑB�]u��2TWQ`�����XR��4����A���-L�؏,嫷����v1�nt� ����G��P��,��j*�m��W�_*Y
ΎW{��6�+Er�2z�<�_�tz�Uc>�h*�u�_�W�ڢI���ٌ�Xj²�-��0���=�
���A�tI��f1*��b3��>��B��?n�J?n+�sV���x�a�q�G�����[f�ΧN���-���}�V ��g�븼���,���yбK��y�x1a󈞞'/&�.�ac���Y�j��{��Rl�}�T�+��&�5eE�����^��=Vk�	4�ւY�h������q�!p�|�kѪ�;[Dm������jZsJ/�����k�)L�G�����) #8���=��H���뱉V^<W�3��^���bY�}�*��e�Ndo��ߓ����]
�_/�z�=�R�癬zo�h��k�uR�X�@8W[���ݽ��z.��su��'9U�i�G�x�W�Z5R��v���vwq���2�����"�#m�j�͇lO}2NW�˲���̉�Y{��b�b������t�bT�S��ƣ�4v�ӭp�ڂ�I�z�H���go��n��_Rvߴ��p��^�fޮ��W&�o�m21N��,*to���dދO�¦�互���k�(즕�8�e�Ӣ��6���|�[�;�j���#��[0g�k<3��+��x�μ+҆[A�m[j^�s� y۞��h�� ��^��4�c�c�U�
�T���w�^�g�d�-1�/k�$�ʴ���8_�Ȁ�́�-�0���am�W���{Z8��a30��\�L��ʅm�+�3�]�������b��]ʀ��GK8�J-¨xW�T���Z�mF����Nf�Wx��f�:�\�88��&!;�-L㩂��`*�L�1F��x���fR;��Uh]jƥ��
�6`��9H�|���|k@����w���N����9X�yK�g颭G��v'�6���+
�:��6�:���)69���CH�lA]��o�Ѳb⃸�殾,�=F���驥�ʫ��E�Q�;m�V���x/Wv�wvq�95��l���E���ZVa���¡������*\�jL��*~ͺH�J~��Ӝ���iq�[j�#2�����G����(����.�p �?[�*�*�
�[Z�_�ߠ�Tt�Zn�:��yʗ�^��_�켫2vn[��jV��lw��VՎ�����J��T����n�G��hE��.�:�>Դ��E����&J�hO�o:�.ղ��q�	Y׵�JJ&p�M'Hl��W.E��`Bk6�6��U��/Д�1z��J���+|�W����ޔ���U�!�~I{�7q�~i��0.��}���3�y~��Os�p\�kMO%a޳_`je3�r�kn;3_�����$�1��"}ܫ��J�b;
Ɠ�"EK�z�k-t'qԀ�VM�Ē�#A5:Q�S����:������B�l���p�s���nB\�I�ʻOTk<��Y�O�\�r�8.�UzfP瞺�F��jP���Y��)�Ua�M��ܲ����E,�pԳp0Drfa@Ӓ���$��&K
vaiA��P-�wo����Դ����U���/�ʀ�y��V��� pc�G��t"�;V��]{��ow���~Oږ�G�u�IX\�h�N�m܎�ub&�Ē�CR�ɐ<���	��{���/�psܳMC�E���+ڦ��̧u��Z92y f�L�=�j7�
6�ؚ��@vѳ�޴3�C�DH�r/$���rb���쳐�b5�1q�� *9��EZ�QL����>�^�#�_1���_j�o��-j���v=�K����wZ:��U��dwڸmZ����F���q�(N�u0:!�������ٹ��
�I�bǟMc�س2+J�ԧ��yG(Օ�yM�[�1;�1�o
�@ЮS�c&f΄_L�Y;LC�<�DWxC���:tO�B��k�����̌�H��g�6�*:lN-�9T�'�b��.Cu$%�L��㳘n)��V�@�&x?�Ɋs9�s�k���׶��pt�k���?����9YK}ج@~�Hk���l�������QQ����v��ŀe��P���1=���i�;��]x
�Ȇ'E}�}7�z����N���٭F�׭����N�(��#< ����n���sCz �xb����͑o���j ��,��튯�33��=g���~������gQ��<���h1����	����ᠮmD���x�����E��iO��&)�C�ٯnƫ�'����\�%M���Q�c 2���'olz��ˡ�V�
�Lq�__
��|��c�k�����W��.����v�o��� �+�[�;g~�R�S!`����Ğ��Ճ8ԶT䗆id���m�k�}+Q��y�n}Y��]�Z}Lqy^|6rJ�S��jJAB"�#,A�*P>�\�Y$�Y�R����pr�v�Nw7���)x��\�%��%N�EM��
���ni���7�l75>�V�]G�p뮄5��z���3G:�bI�y�d�V����뗺�7� e�!��\�>��&D��ْ�;�S�;���)�t��iW��.Wk:Ua�;.�!��"����C�:����ͪ��N�$e,s�w�X��iR��U
���9�y��E`�U0~^F+/�wsRu\�3�/
��1��6��s�k��A�^4#�![�3gi���MCn����)��/YݾT�M;�nADZ�#�h �A���Q�^QW�3��,��+���c�ƽ�Q�\Ԓ>�u�~�~>Q�3婓�Q�z!�h5j�-�Fc�+�jLv�|�Yc[�D�Z���M�w
~fcj�0&9�95����0�fm�V� ~�<=���Ȧ2e�^�;/k�\�t���X��ɑKd%��f0�Dϯ�T�Wˬ�4H�nU���m̵)x\���sA��Ü]c�����+���MbF*p�1鹸ńP(}3���yZ)+�kR>Qd��A����J�'/&��-L��Gs�gY�yC���~�(R�6	,U�2���l޳��o�g)�btB�Z,�c��!��&-ֈ�ʠtJ��n�=��m�Nd��8��`��R���S��2U���ؾVr��Ë��,n�m!��L�A>��[���o�/dӝ��k�Y���Ss|�i�(j���KGeִ�&��l��%	������Ȧ����LK�L����]�4�ײ�J�*t���m)�<׼zA��q�}�Hgٿ+�fu���"}*@{���� N��j{@�ln=zc8�s]�i�+�&m�����}��ȍ���!8�'��M,WPྋ=oݵ��ߥ�-{<�~�	v�Q��j�L�K�c�Ҳ�Zj��\;�	*�����U.�CEZ��tHz-k�\���Ch���M
����"1�c�jǧ�Յ�}�7�p8����6��p��5�S�VD�[1$�3�}ʢ'��mg��$=���)�Nx����NMc��m968�6i�Ph|ny��F$Hh�t�Bg�I��1;�����{�ќv�����kd��q�Pp����(��`:6���tvJ� ^΍�U������0g:h�܊M��$Q/ݮ�k�W�D�)��#	�WT���\f¬NX+`�@ʹ[�<����L,/�v��ֆ�c �NO9��"�v����k�ҝ�!�����]���^�\��4A���r��L�z���l9��>�V���O�f�z�1e��2� �\�y�a�U�T*\���6[�l��{cc��|d�8x�p����r�s�����N1@m\���m�1���)����.����R��� :�7/���j؁��M�/s�]#�'����f��,k�c�p����]�v������}�>��]g[�N�Ѓ{_ ;���ߣ�3���	��0%T����Ga�N��v*�b Ȏ�lJ6�8҆W������9�tz��m�S�9Ō/���7�).>��ׯM+����Qc�"���5�j�ˡ���t��0�z:]`�r5�qv���4NLF&_(9^K�G���>��EOl��������_j��a� t�>��ٹ/�b�<+���! 4X�.9�>5�,f߮`���3͛.���5ia�f��O.Ϗ����1bZ���.����|+	�S�A�B�
��Ո�ƫh��_a���� OI���[ڒQ������en����ub�P�dO)�yt~�xf��w��-1�����`mN�^��c��G,o�☫(�G�o)�Duc�����&��NzZ�|��G�7g3L����
��1A��$�@T@��tI1C"&e�U$r8"G[T�_��g �W�@s��M����Cz]Kd{<���;jQ�"930�fΫ iXw�2�1t���SP�a���0�7��W��<�O��^��=��m�-���R%���3>�I3[��(�ۗ��6�y���w�ou���.��t��������������Vi��ֻ�¡�]Ⱦ�eg �=Y�0��@��E��t[+8�*λ�]t/��Wgb���FQ]�F"����Al�yK� C��{"�(��;�q7١���5�\���8��f��!ᴝh6�܎u4"s�bIB��M��>LA�b^t=�!��l�u�"��&oK��0����)��Z��M�6�iO2���D��o���#w�-!�[������T㢮��R����I��r�F��F�"��d��d�D]�ț:���Xf�>\�ҁ�0?�����|=e��/�?�:�m3��O�x ��d��mV%r/��Z'����'3)td{��Ɗ�ٔ�
�v�XE
�4 eή7�$�h&�[�;�f��YC@;5	��q��s�f���"M�uok`�t�_xfg)�o+�7:o��{��0xvgj�6�����cS���g ��N�=^��!+|g;onV�;��3�$=�Tcʋ�3�/ּ%?n��'�7P����;��贐��Ԭ�k+�x׽��<{�UH�M�U#�zP��s���O+�s��c{9��ai�u1��rWVƞ�۹�ᆟ,�́0Z�-��k,���-�T�8�[�U�'>�\~\�a�^���$��+Ν�h�\��챜��7w�
w#�ۼ&�^Eג�o*Zո�B���j��_)C,X���aE����Nħs��C%�솞^s�7���t,`��*	�➖#��TJ��a`w{U��:ϪzW)�Sa�{����FI>��j���H����:
Ev�/�^O��i^��
�Hxl��%>9����CNt��Z��=��yq.�F��e�eWB��Li�c/̩�6�7�ĸS��L�V�ݒ���;-�5a�\�3~�P�pڦ;%������Lp%K���i�=P0,&z�̐��J��x����G��
zh8�0�i��D7�R/[�e��"�j$qW�#�S�B_o�3wK��k:>�	�ؠ� �U�	�^F+'����5�񔻺�/\�_��U�]� ��
���`4w}!u��l���p���>���lu]1�����s;�Me�2p�%tCz$;�� �Zg< �$�4c>�s���;��ʯ�R����9=�EXy���(�̪Z�=���>���Z��G\)U�.��v㤚;/_jڥ�ڒ�Ѡ��R���!��0/�C�x�>�����[9�Bg(����mҐ��t&��˼XwD�ưK��K駲v���z}�A]g��G]/t�_]_4k��|]Z�@}Ov��6xB�;���HB���Cg^8(�v�v��ko�ٔe��&ݾ�M+����l�����[#��8_C3��4,��^�#$��Ml��J�qH�aNgX�B�ո�3<��;\| �u�l\��g�
l�h��'`�$�Q�
qf�X;tS�h�9�i٩��L<1z�y���ߝ!��|�����.��+�vťca��s�|�`�9�iU�g�wO��*p��d��z�S8=]ε����ek��8OI�Y����������ݸ��*��5�PP�6�x���CuT�U�Ԓ�c6�Z��7���}Wr�9�گ.��Nc3�!̡ͅe���c�*�@x�3b�_���y�	�!�r��YsA��n�6��2�<G|h����}���+�v��/)�\�o{]�XO����0�JXL�K��;%m�M�Q�EJ�U�\*c���|,����<���!ĝ	����43�dX�a�mT0����M��{�h~���k�ݾ�Vn��߹��`�����*�4�xʦ~�kE0����u),������b͜9:'4�,��^������z$��0(� ���y�!�^��HL��8X�G�LNN�=v@2+I�M촩��Z=�W,�I�i�7V�Ҝ�Ӫ�.;�1�j�U�s&��#��-�k{�F�"�WR:*݂�pf�*�
gJ��pc�#Y�wZ�=�}�Źl1�Mc.ѫf��+��m9M�+�������P؎�.��76�J`�7�w$ˬ��gfW�cck(��G�d�����%�V�rA-�x&�8+t��T�^06�k!�4A�I�z�VU�1��g��d-*��Ot�c�2�ͼ���,7mO��7�����W����vq��Lk���7�VC/�r��W�uݐ$���u�����쑫E�� ��++��s}�J4uv�;q뭡;�����@#���]��ʍY�`4Uǀ+��k���V�b.�-��(Llvv%m���_v��*bB��ݕЪ����IS�E�1�8&�g 	g<��-dF�x�C{jQc�n�ゆm
:�+������%��R[He�a!�{�$Eリ�C�lU����m
�B�\X���.�i+�t�P��or^��y:�%>�n�q�2�� �L�#۽�=E�V���tTE_��ٱu���~z�w3 �8T]̙�����qfT}�4���	͡x���cA���5i��a�A�{I���`pγڹU��a�{��h+Є�a>�]WB��C����K�r�:qlYZ.�m�仏N�+8�g��:+[m{i�|&R37�_^+�X�0��Ӝ�h[��Z4��1*��r��֮��n�I��L���\�Z`Ŝ[�W'(����GhK�9yXV�حl��/�j�Hwc�_7pC$�}CA�N^j�I�ٰX�gw39]�Ch:)P4+CyR�L�P���l���=�w7���.��k2>����E_�Dp��v�%ٮ��댋w(�,��3y��[�5�Wwf	y��e�"E9������Ԝ�\�t۳J󊸪�߯dS*r�2�;������VN^�j�.s��I�0���՛�:��]�y�+ʕ��q0;S�j�S�A��Z.�
���n�b���ײj�Y��K�8z]A�β�v�۔���r\�:��߻��h�c����b�T�u'�u8�d�tȆ�if.�]�kG���.7J,g*�0+��Cqc��y9LM�]^�G��m�XF�g$΄��L��=��l�Ŝ��;�Mk1A��{�Z�I�w/`{�"l���.΋ 9n�I�ڬYohX[T̢���Ƭ̅�\�����$;X�>0X�/�Z8�0P_	�zc�St�$�y�9j]Xom�>�G�jZܖka�8 x]^�Z4��v�di��X���.�S=N��/0��k ��g;� �T�D+wi�K^p�%�Gi������`�o �н}��Z�u��;��p��Ӷ�r�p�� �VT��{�a�Э��;��|��:�u�H̷��g!X��T�ʖVdB6�t���pL���3�u�0Vثaʐg^�����"J�"�"��(�EU��#��T�	��q��.�\�W�67�t�nsIr+��]�<qW�D�.h�\w\7	�N��Dn��wEF�N�[�s��N��W1�ː��w`�.Ne��ܗ��.b�E�v���v]Ӣ�������뻡�Β��q�9^/���.��vw\��F;�WN��.�/⼺��r��\Ԛ�\�j�i5��ؤ�7n\��Dh\���̝�bH�p�]�*+��H�ps�!�Nws�:uv�^93\�<x�q��9@�s�E�]�d;�.��n��#cr��뻺$�Nq�\�g;���r�󫘯;uΖ1Ww$�t���;ws����a�q4d���Ӻ�J)J�tu�˻�J�w�y#x�뫳��)�D�,�E&�$5;��c#6>��$�J.�2m�y�\�3�ٶؤ������ܪ�Vo`,[��ɜ��ޝW��ޮ�:e:x��ǆ�ft�W�Ǒ�<���cwfk�������>C��K������h/ϝ�^/��oϯ�+�v��~���ν*�Ϳ[���;oJ�r�o:�W�|m�y�ux������_}���.^�_<���r���_>�`?g��ru��LU�}b���^K�+�s��w�Ϟ�{k�]������}>/��{]�k����W޾yzs���ԅ��}T����Dk�~�*��"���`�b�H��L���A y��!VvT�?2m�M�^��U.��"�௮��z����|iL\����c�UW1�~s�}|�ʋ}��7�ίo:�5�}�{�{^�������w��n~��}o����� �E���!#�(�C�ɜ���n~Fy��"�� ��Կ���+��U�+��o���k���׭~��^��\�cv�󘊘��O�S�#_|�.~�?@��o��yoj�+���^a�ڹno_�<�����{j�}^�|����5�y4�>��������{�
��G�>����-5�����o׵����}~�ޚ��Ǎ~|���-�_�����^���h���͈���xߗ���z�����������{�#!}6<x��" �"יڱ��;;��-���v���U!T@��T��Moߝ~5��<ޚ��4o��yu����}������^�m�/}o�׋+�>�VER�}D}^Q�����4U����;���O��_w��T�U�_-5
7�k�����>�kv~��}bC�4�(U�r�oߞW���/Mx��������\7�^�y��_��i�Kŏ�}5����s}��;}�����W���۽�Y3�D�|� L_�k����q��y� ڠ���5^�c����Ӓf"���ۆ�~u����կCQ����o���֘k��ʪq���>b�EV���
���
��{���_���o{�_J��ڹow��?�������s\�'�����D��|�w�gv �~�&"���ƣ�~v�[��?�ܯ��5y���צ����_���*��M��W���7����\6�����~3Sd����1�����xU����������)����r�=�x����]�\����L�\�LEKc�c��w�^*�so�����ߟ;os�����W�n_]��{W�|W}���>v����4_���?�������m�{���_���o�྾z�oK}��j�[ߟ>��|��Xq-��o�4���T.]��Bf�V"=��sj0�N��u_��9Jc�Ҁ�*��7Q�Ve%C1bO�e_K�r�5Ê�9Ǉy^�Zz�T�F�т���t�3�Tj�J�1��o����r�rR�"�4�·tȻT�������3���-{��
���E�/?�oO��h���޻�������x���~����W��v�^y�~|�x����m�����k�y���zU�r������ƿU�W����W,zW�^%���=SY���� ������?tǨ}��ſ��<ޕ_J�ͽ?�/�Ÿ!Zb"G��u�z&-O�B#�=h��z�=�,�����T�k���!of��޼��쟣�1�LÁ��S5r���<��x�o����^oj��5�{��׫����_���{��ޟM\׏�-߽������^���k�y�~w��L�s��~1�_B��#�q��@�t1G��������_!�W�+�V�CM}D}\*�>�|����Z7����+�{k�/��+�_����=y�i�����ח����^.W7�x��}���7���-���G�b*c�^o�EN0Ȭ���{s�n������}D}ZO�E`��	�����ү>�/>W��V�-����}1HG�'�S,DW��sb#cA���wm��Ϯ�F��+�ο�:��;��>���9���"�(�\�z7��+��V���"!�#�#G�D|�{P��U�z��ޟ�~+�������ן���U~�>��W�W���*��#�u���/�rޗ��x�ǟ�k�{���k��J�?{}��𙟡jkz&�:�j�{�r=��h}���=��z4G��뾮�^~��/����ή^-�_��<������W����K~+��W/�:�>����>|��_J�W5��|�����x����Ϊ
�>�#���mg{���`�/s�^��K��3SS
beW�s�����߾^��x۞�u�����s�P����߂��UM����*��A�~��h����_��^7��y��QF�c�9�X�@��n��]zh9��y��A��G�V ����(��~�1�C�ɯ����������W��y�zW-�������W��5���^7����������Ϧ�_:��[�\���/^��7@څ?E1��&`�}��MqkƁ��ۘ����zo��ݷ?�/�y�h�����a����MT����X��C�!��O��AUIs|_�wy�^�*�\�/:�[��x�׾ן�\��^���^�.o���"M}s��0�����vX����Ap��vj�w�+�8_y�	`_f��'Cr���v���u;�����q�k��Q��ڜ�X�|���(���vG[�V�F�ѓM��;�X*_Z����3 �Vq��	Ħ��LZW!C{��w��NP�%X�1㫙���t먘�)��xI��j�ԧ
�{q�*||<٨nhF����fg���Z����yK[��Y�%��j�=G��޸4z�ǂP#l���
���-��Cz��S��2�k����Qi��Mr�5���-��}r ����y�x��5��q����sC{�X�68'NH}j� >���޽�F�?�J3b<\u^��'G�\�0.'��9͆7�9�5�N+"w��-�qZ3kkzs:D��h�n���f��:dAD3����W LGg�ҹMΝ�it> ���E�K���I�>��3�*>��]�Z5i^	&��
�&C~�@m�>�]�����暌�	>糇,���nVV�;���'��ףF� �����ݘ/�����ߏ���r��M2�H���mS�����IHƂym}��S=~f�xsq����{�6'�8S9w(+��V+���8�H��E�7V��:$EE���^t�z;��p��{���T��ʁ@�G�#�ѱr�����[�Td�^F+-]�5�����H5���R+T/��w���IY��Ds��ܶ��ѐ��1G�/�R�z���0q�.ms��"������#c }��Ք5wq�v��*��V�ț��X���u汷�X�M�;8�q��(L���E������T�����38\b��d��1O��q�F �U�?<�}���m ��h[o�{N���}�oG_���qW�SE��Hmi��'�r���:���g�.�R����f`0#��wUc�W��gB/(��y�|��Q���2{M�G�sA�Q��vc��҄{tAN�sV�OT����״������p ���P���V��U˞Ø r�㵟~�v��Qˏ�m�զ�+j��sh����;� +s��F��'�]y�Ȯ܋�ke.�V��E�{��=���lt���ϥ1�/WP�4��B1S��F=7 ���Җ�xgE�9��ҏ��
#]V�x6�f�R����v�㪽?�qb���w~r���!������s�N`����Oj$n�9�"a�2&���R��(�w�s'�!a�Ύ�"l�{�ݫz���Ϲ̞ܧ����S�^��_�*WF²������
�����ț�盋i<��C�I�vsb�L[�e�S�#�4D������zkC�yW�j7Ď���2�Z�E����':Gd�
�/�xbў
��J �3UZ�t�*��]y-���a,����r��$�WKb�v�R����z�O-�rێ��t�N�av>H^�������k�rYæQi���&K��ygZ']P}ݖ��[���[ٓ��Q*�4��;�
��#t��A_�]8�5䩄�K��4��U���k��$��sv;fE��6>�f�)����ɹ��F�rxr7��T{X�b����a�����qx6tO�ܯuw��93xy;�}"�{NR�2�b�f9��xD��4���RY�
�ټ(z�4 ��y,�M��5�s*Y���@�ni�@ƀ$ܤo�3����������,�k�q٩�]|l�j�8\
�>L�gmH����k�mW�t��n
�w�����Y+3�uV(��9u��C1�	m̌�v�*�dHB���6rO�d+����ě�ǘ-Z��3èɎ�Q�����x�P�I��W6��JE
\Y>�P���S�-��ZоQ.eoN�����$Ln�d��������g��'�ߴ?z�@�l���Rȸ�A��x�:�|=ɇu���������ѧ5}�]w/P�_���Xyp^9y�UX�<�"�BU$wo����5{��1֖f�Z��f�)�)��VR��������F_8��Ή�E�������oi��B�mb����~��;�T��튕�]��t�3�b�^�啋�KYW�{�deW%�+[�U+q��@*�v�0�솻��ݫ�-���>ާW�]:\;4�7s`J楌%m��<���uǜf���֤c�ڀ�WzS�+�X����Qc�"��x��^������o��ƫ�������^�QYN/v�^��׀-����Y�M����%S�ck�f��ρ
��
����i=)Fe9���ŀ.�p53x�C���sc�^��Bs�pfC�8k�y\U�LA��
ѕ1Z����p8����uq=HCQc5�M�^�z%��=��^(�{�-�]�u�"lw����.U����Y�u|�*<3�Oy�]�m�xf���������ġ��B%�2#69�3B0S�Q�i�X�"�U�>s��ʹ2P}����ӯGdm��Y����Br�=�p�ռp"i������ho��9���b�v�{���O.�Ԟ9~s���+�Cq�0X��y:�t"|qvO
�p�qk��K2��;zCy�X�E��WI�{0FS�(f����>�g�иK�d�I��x^l��7&�a����SӺn �!ᴝh7]��wV"jĒ�CQ!�Ė�e�;472���D�#��j^ҧ�������x4yo�Kͧx�5ڲ��f^�H�^��+X�]���z]۬�i��!Ύ\-;�w��#�e_[9Wt
;�4�+�o)􆹌z�^휎�v�D�2����V��onA�k+��Q�t�rE2�_==:a�C����dʘ�7��?F��6�cB�d�n���hK"ޑ���`��97�����I#�#@u@s�$Z:"Bg/$��\��I��s�f#_eb�;u��#.[]��Eԯw;�#�.g6El�i�4<=e�5��_��7C^����Zp�O����̐+��}�+ߟ�m^�#�%T��F��;9�B�}����e�&�:���ݛ��
(zbb�Ok( �9-��.}�ٙmN���uÕ9��^� xU-�b1��o �*��J���n=�GYuS<���o�m�����_��]i2!�<_;�r�-]��ɗ�$��w%�}����*����s_5�s,F�k�e��c���g��{7���g.ĝ�|�8�6E�:�N�n���,�ޔ����F�y^�����ʖ6��N.�ic�f�|z@���N��~`��͋`�4:+f�C=��`uF��&#��9�)��
5nU���w��e�%��%M���5X��qȩ�Ds���꼟K�J�� WBG���*���K��{d��Ps�,ײ�n�;��F�I4��*�Q53.+w�}ư�v��J�-o���׹�])ZZ��t(m�iPG{���6�y���r�C�wc�ܚ�w�ż�\�Dm��Gwۣ���ONu�9a�.�,���=����÷�*����X�gŲ��ˏ��q�ԏ�E���8'¼ez�z}��J���L��U�*B1����qOn�g7�6}�N�S-JFoت zoͪc����9%\)����R����i��_(���x�����GYl�;�u"����p�7ڈ�:��B�{�x��j��� ��]���.�z*#�h��t5�~b��8.W_�otE�Gpy*����dWCw+V���s۞��^������d�V�**��݃��������<������K�> �=��ͫ�(�GZ�!�O��s���H@K4hQ��򸲯�Ž~���R��e�'�3����# NX�)�tnzh��!����^�َ[�Mi����=����X}i���������}qX>�h*�:�'O�ڲ�Lf1��Z�4G|�$'�l��������a뙓�z�B゙����\F#8$��lJ�9�G�\#��qȽ����}7��F�,G�B�~�g�����\{������Ndu�;l#U�����ޱ'4�v�=p�Vv;�U4�}n�@n����}��n��+�l�M���V�n;
2�[����7�VV�υ��b����*wP�d��n|ݽ�c.e�O%!��9�)���.�C��2�sg��I<�4W,>�N>��z�Fmz�(�VA���E�0F�c�Mf��dܫ\<���+8��Z�Z5�ʲ����f�qx3��8��cD�`�Z�.����n��\|���8�pC���vY��ҳ�v��Z�W�&�`�g�s�+������H���T���8j���dNàu.�0$+�z�4���j���	�Nw����ƥQ�Ǭ�{��S�q�����]���x�ԕ���I��~��4=�Ҡ�ײ���@N)�%L&K��7�V���u�r�%S)���0���-����pL���T�B*"J���4:=�R2,c0�ߛW\9����Z�#���^lu��Bl���NeQ�i�U�Qpj�P�#���l��.�;@CI���խ�b�E������}=��V��;D����0 F�,ܤd�F$H|1���"�^�8If����k�he����w��7*��3��"+�M¼zmޅ��r��m�?|�n��&57�K�Ո�v�*ulƌ&��R6���EY�!
�� h��<B��ci�dfþ�*�4����3O:�j�=��Ke˴ա��ZԌ�)��U�t�W��Eq�3c�����!�=�q��tn��vk��[9%9z,N%*0����c��;���Ų���Y����<�ζ�l&�f�˜�Z��~���9cRZ��ޯQ�O�1�o�P����8_���^5`w��w\��UB�J�4X��ʻ�-����Q$�S�v0�kxO��H�)��)t<�k@g�I_ID�G�����VȪ.���.$MNU��	���21x����M%.�ދ�y*�w��ro�-��'��a�(����)��5�l?�+�Xx]����<�n��.���.�o��ms��� �	Lh;~N��s�pJ�c(�2Em׊�5�j��,���e�������)��uږ����9X9)�z5�<n1϶���̎u�gu}��6�7���[\0�z8�k��\z�q0���\.:fx1�ߛ�|c5͎�yz!3rl^�:��3X]1_-�^�a����yv{�TN�"
,$lk�D\OR�),^o��Y�xΎ]^Pn�N�-y��9:oB�W�%b��-�s�����xn_:
�N!S[ռ6�ʘ�
հ ;EgU`��{M�3�r�KL��h����x�*ĪJk][�7s��S��}Y^䛻�L{�N��n<� %�8o�E}�뮬I+�y�����k���\�| U���(2�Q�^fwuB������"����R��soi|N�6uL�g��ega���ZQ���<�a�&��z��C�.�� O�_>��Ԏ[�v��s��9MP�:���#<h�.��w��gp�f���O�ap���IK[��T[��z>S���n$���;�\L�Ӭx��=aGB-��:�6r������.af%�=�tS ^��m��hoq@EI���W���eE슍@����Kr���t^XxM���������x��Z�%�e :�ŀk��c��\,K�%���e�4�7-��p��j.�w�vuɽ�t4�����Vp��3 ��2���f����\M��'��v�ݾ-gn-`��Qu���mϮ<׵�TU31����S��V���e�Z���X�mucQ�3e��H6*Y�M:Pn�̓*�����8���Ҷr�7I�J���F�M*C��[;��g.���{����/�f#��1g���Ws꽩�Rov��A�m�ܕ�!�+Tқ�S7m)ݦ���Q�n�k���F�T� Qlj�u�tb<��p�`:�[݉�(��< b�4К!d+�1�S��]�/���I�U��Kq��V��κRYS{Uskc��b�C�#C�zꖎ#�j�R�u��h�*p8�-]۶�mH�=�/��fg9.��[Wd�`����j^8�Ӌx������P�����T�q���T����ުKw�v���_���}�qIm5d�Wlժ��쫘:(��q1�����1w	蚮�#���Ae�5�`�@���ic�|�m���CE
@<V�.*�YI�V������g3x��\X03�a���1р�/�������0�-3���9�N����^�7�Ҷ�[�[:�����ب�@P#0CN�P:v���׊N��]���
�"�R�aG�KV��P���<����Oqaڙ���1�}c���1��\Q��0�AK5!eٙ���X01|W�@��4��]h��N��jE���kkLa�}{h*�u�WsM�ĎfԶƫX�潇�릕�$��#d�i�u����\��M{QK!�]ڒ#C	}Y���V,X�<{RB�#RL|�F��[j�\�1E��S���T��W[��WhK+y�E�Xǔ�F���}t�9c(�M/�ھW�8/�ܔ�7f5���j��9��	�;�G���4�T�0������*R����Q�������>�9�w5uyy�u^���=�u���A��T�Cb��I5����[�p����v�G���Ӛ<���Ă�'�o4[`ۗW
32����t�W���l�J��Z��΃ �0��wx��Ӗ�-i�K�:[�O�c��'2w ��W]<�f�t�fB�Y�'[OG�ͤ2V�0gdU�2�Y��l�ۥ*r�m<4��D���M5�ږ����;GR�8r���}}}������������k�eùԒ�y�]�,�;��;�`�2nk�wld�˼�-�np�uu��鹬t��ƝۤI����uy���˕�;�Psn�;��IXV.k�Ȉ��+���w�.b��cr��t�+��sn�n���&rݡʻ��u�t���/�:o$�^#\�Aw]�����d�c$�w���NtӺ�wA�/:��ww;��d�wTg;�������F�&wu9ؒ ��;�BF��LJ�"�%�u�r��jKr����wno<�O:9s����.��ʹۻ�1&�s�A˙-�n���ܺwu˺��lY�D�r#���˸�wne�s��wv�5�Ûw7S0h�����<��(WWQ�%5��e&�O�֭���{-w"�0���]G���8U��`W�nS!DӮ��l-��ĥs/+SV,ͥ��vջz��UW�
Ԥ��{�1��U�w[�|7
�M���Մ*�/���( {۞�V2�M���B����h�~Ś���n��Kr�r�}�P�W��b��i�%��rY���r�>�j�Z���۽��<�};NTƷ|����y��W��*����Oj.�=�
ݨI�x�םS�IA!G8�[��x����
��oM���)�ǻ\^�~G���B�C��zʻ�9zto{A�P6��>��1��kf�9�
ac3�Bڶ���~���a��r��[�J[��[Ӄ�<�C�(�v;���>֗ZY����t
�칻��ڗ�����<�c�#9Q�2'���A��3���eJ�<��Ʋ�ݧ��IE:��>^7�1{����B���*�Q�b1zEB��b�,��:W�D��%gԟ��o������l~u�;W��	���P�����!�U)�jl�".Kn\'�m7��V�;>o��+��Wme�Mյ�+�@�z6�w�0I�o��yd��n,8ح��Ob���i�}R�{$z�1�
T�n��_1���]{r�N�<q�n.�W���_�}_}�Ջ��%��=�s��Ę��^���W�=z����|�tv�F%$ס<�b�^�q<~��6�,�ɃAU��K�w�?>��}�;�V�&/_��h)��G;KN����VVk��fTק'�%C�q��G/n�.X\�+���|��(=U�HK���r�og��!T)�L�˓}R���`G��W�팒9����T}�7��s���W�7%��hP�D�N�ʡ����įM�w���F�EV'R�<�_w�E��i����ªq
Mj����a�Ĩ�=:�yRW+�Ur����mv�p�^y�����\�&�iR���%G�'^���"���M݄��wyۇ��ƃI���F��_���%�Z�V#�-������y�� �:b��^v����]ݼ����
M�T9�5HU��Go�>2mi����s9u�{��Jf$�4��n�h�k
F f�����sv�7M�-ǔv[�����9P=F�P��F�f,�[\�d}��Of(o�:�u�L�6�Qwv�|��fe�-�{���*݇k�O�-bޜ�
j̾��R�"��z=��Ƭ7Ku�bol��hW���Nد)�5��[5��麂1܊�{z5�h�To}�k�Ȱe7ޱ��k�r5�E�;s^=A��(C�$l$)���q1�jEj�EW������9+ꔝ������Op{�2�xܗj:�!����C8�[�~�{|4:"cz[�;Y�q�{�ݮf��^_<{ :�s=�:]b�_yZ�i� \Œ4A���h�}�Or%��d{S�MO7��e��n[Y޹�����f]6an�v7�O�u==�E,w���g��W��N�%�v��S2���1!���u��и�p�t��ծ*.AK����K�Bx�%�����<���S����Ǥ�TOC��K�Pm&ji�t�d�{�4i��®RV,�U�I]3��B^\��|��uc�I�����ܙ7�و����x�pi��{ ��B�ـ�M�y���I�3/+.��3wg9���&m]�Hl�im�����ѷb�����Ѡ7�s7��]��ڢ+�t-��ү2�GI��+1�2iΩ�Ӹ��w�{����9q�mou��c���ﾪ�����r
y�����yp�c���gz�w��q���Q����Q�5O#}|��M=�9^�M��Z�G*�r�Cؘ�I�T�]�G�3^q-�ɻ�����~r�m��L��亵�Vc�dlL�O���ddݪg)or�Yo�Z�'�x-iD3�*gkͿ'�{��J6%,��)Gyw;�x֤9{4�K�ׁLf=��$-�~g"a;sP�\ɾ��t��މ��<�����z��ېe�i�=�N�*,�B.5ߡ������л�MS��jVG�i�c��z'�j�<��ESί&lJ�;J�ݑ߳7A)��U���D���-X}dλ�;�V<�Փ�K!g���	�(�$2.½Y�ގ��>�i�ڎq�Z��V1��'3*V�gO�J�u��q)�]�a}p�:���xC��}�;<�+�s87������ѡ
ӱ1�j�3���?<��k�;v�v�=���K��2f�]~O��,2�k��m�wG��;�����qEo\�0&�s�N���Rޥ��t���Gk�
To�U�%Y�8��C(T{@����+7��m�I�rKx�=�W>xo�0������g�o�-^��q�9�3ֵ�QG�;���k��W�Ø��<��B]���]����.&�
���։ת*<y'eS�n��f��.NM�em��Y�*r��n�2��rz�B��}Q��d���8��-�a��N��tc�5���P���h�P��3//��S��׵�g��p�O�y5�z����K�%����cp���
��n�Ȓ���j�+&�	ș�����y��%�|ҩ��\-j��X��nKr��*4jZ#�c:������p�����2��T�ې�c���C�J���ֽ�+d��H���=��+"`[F9mKj'�k�c˄���x��:�"�ط܁�&��f�ډ'/���f:`-2mi����K��A�}�}wП{t�˳m�Nv>�)�5⧍x��Go��3�.��K��ƺ�>� �� .���)� A�C�JEx���F�{r�m&�w�o�8�����7(�4���h>m�����Z��7B]aۙ�`�T3N1�Hq�y[�/5z�]^��.�k������|`�x�]�t���,��h��Ƕ�лK����#���iu��5�$z5ߙȘN�|����{eP+�;���M���)�N ��U�S������D$�]�Z�J��بvߡ�1��i)�'+��W~N�j=�ш�E�,��}�j��x���b���]�m�f���<,���t5�2ܷ��c��VȌjriV�����R~u��V�x!\��'���=�����򤌑#Z�����ax/1A�z�8���޹{�b�Ҙہ�	�ZU�޷ڽ����<���C�����[���;4���݊��}��d�v��{�����<�ygؖ�᝛X�mb��㛚+9���b�q%��i0���=��
���r���z�)��VEw*�EgJ��]w\{��xlY^����y&���|����w�
��
��=���A$}=���`3s$�Z'm/T��F�"���z��p�]\$��6p��!�Y�*XT���ͻKʗF���b�|X���MlM9)wc%]�U�3���{X/ISi�|�;i�M�T�WS��ωz���/�&�9�-*�"���A[��w�jk聵h^����ϧ؛�U�o��9O%�ӹܹ�3TWF.���6�Z���������r�)�Do�ѳ�>�w��pN��Q�qp��q�:�Os��`��-vOD�Ƴ��Y�S��qoݕ*��C{G�ks�g���Y3��)[9����㦌���0�%Jd��^j�v���=����b�jH�o;]�9����J�jl�
m�T9�G���W\G�mD�/�
��2��mc�r�F��q��{��~Gw�Jv�)�4zB�f���s67d�,���[�kB���v�}�9��3��<�g��s���x�$�l�R]�i��X�����t0ZpL������Y94�\��j�jp6���	�\܉��׃j�BYm{�F�Wq��/l�o��̿,���Lyo���a���w�&\Pr���
v����lM�o�{Y�֮�R�՘�ɝ�MOB����~~�j����W�2s���M�T�:Ӕ�9�:��A*������|���7�z���u�n+�h�4+=�_[[X��m��yCsg�3a�A-B�mu�f�VV��0�׺�xkK&X�Xv�X��6�=�E�	��c��2�m�O[�;�����+.��hl��C+��2ɇ��G����E�:��u\8��jފ<��v��#��:�԰�'9����ޏtC�r�<�}<��u�G�.��\W�.W�*�n6����R���JuRofcy�
q���Ĥ��U��6�T.�d��Pb�f�iߋ��
�k���8�',��6^�z+䧪�����XW\Fk�e�=��=�5zL΍��L�7)4���P?;�}C��~�h{{�/��Ռ>G-�x��)5�H�0Y!���j/�����<��7cp����ʉb`ZU'��Ȱ.m��N/_<\��\��_p�֘ʇT����׹UEZ�eZ5u���چ���疛��3x�g�,̈�عO�q$0�U�W�\�v����t��u\'w�3��g�<2m#�b�,ǻ��W�
ᜉ�v�ּ�(�h◚g���B�qzǸ�]uI�hS��3��W��j��<갭ێ#G�
%��*>��2����O	���u/)b������*̈(	T�:�U ��r	�5&
�7�;Wu�P�N�\��F)Ջb���L
��n瞞�jPǔ�
�q���{֪� E[pBFk��$���ك�����%7�"�a��,w[����K?�}U�}�ߜj�>�������F�����L�J����h�ڜ���׻d�͙<,�q��[�K�I��o-̝�--�w�Tk���v�a��3��Kk���_#�,�劺靾{�<����R�W�ֶ1|P�J���<N/H��#P�}9���(�ӭ�T�C����պn�z��X��-���i{<!^/{�<�%j�bx�S����W.D�Z�(������u�]B�����hO/���'�6��q3�5���6�_,5�s��r���D�ᮅ��t욌Y�`or�W�;�dU�Xz�.�[r����V���맅u�9̦eMD��zT.�����QkY���x����F�u�����g��a{ԛ��|G?�N�>��ֺ����c��Ř[���^��pmƵ��}��W�8�+SD*�*$n��*��Qs��6a�=/p������Oo�n�G�w弟3C��L�α[�˨T��m���M�ܠٻ��!�\dL52=�`��1w?u+��`�Я[=���R���x3u����Wg�5��lT:�TR�w�GS��-cvh(���@W�*A���G2�6�[�!Gr6&P}�t���|�\o�5���y_�W�UW��ߢ3�;����k�����M�O����mypT꒰��^�w����ی�X����S�L@�F9n�7Q=�^\$�Uyx>��}�"-�5\v.��=فow�TY��L�Za�ؼ
}�v���}7}s��[zo+zuG.���b�ښ�R��l3>����I�^��^�3nr���PQ[�9�.5�#�0��P�ܳ�{`++�ٝ�x�̲=�0��>X�=����
ww��L�j`�$�]�9Q�2�x�6�m�1��m]lk
έ����}��_t׳���9Qz����i��qs���(nj�������C��V���x�w��=ʽG�`^1x�:�Ԇ�ߝg��hy_�owR�Gө=z���;\�eq�w9�^��*1A��������;��ys�\vq�(�)��j^��T�Q�%9�E�#�&�dJc�1A��G�I˗5�]<l�~��IT٬S�t[�t���}-+�B�fM���Z���)�;�ҳW���zm��r�un�5�}���]�c��=y�rڨ�Wq�s1ֽ/�	un}819̻�Q=Ǵ>��S]���n���=��W^s�VU6�C�^-j��O�m��e��3�,�݈�c�S�lֽ��.ҭ.>@ҧY�.�զP�Y�=V3T���j԰L�G�:6�1�6����r���Q�H&����وa��L5���TV��/B�m��1�sn��bӳ��C�>Čn^�}f���jݭ")]�&���t���g
G��}��F��=�.��K^�y�̦�����Vs�bdj�����Q���r��Ü�+�6���:w
�7uL43�jH�"�xn������K�Q���G.�i�{u*��yj���\�� 4��A{4�/WӤQsw��qq��.�$6�)�(��+��Zf�*�Y�Ɔ+_v��s��%��u�B<�E����V]�uaH޾7�#�Q�F�-�����F	�8C$�J=0�H�jWe[��r�q6�K���ޑ�xZU�Ҵ��kb�6T��-w0� ��;0�����u��ݾ���сF�<�Ĩ�&�y������9�r�'Ώ�[��s�!ͬ�$/ 2wj�Zbj�����m1	\�Ӧ:�$�H�<W��SJ�ր���Z맔��B�l��L���ܐW9��[�ܔ��,�o)el9�.��N�Lu7�&�P*�$�٥r����J
�N�3�}����8��
������u	]�n����qÅY���L�gF�>�`�Y��2���@X��)�p�n�-.�u���iFL4�\��|&L�`�ݲ�2�ъJ�ikzN�.�2V��$���/������UE����亵��+k/�u��V6i%k�w�>��a��k;��ڻ��a<���9���u_Ww:k涹��O+�t�
��Y���>�Ε�U�Y�*�m[��۽��̓U����p$�J�6�5�VA�a���+�P�q��8{�o���=u|�ܓ'H��ۮ�c��;�92􊔄���9��N*�X^������9)�������uІ���̻[��mE*��H'AT:Z�G�	�ǿ�|��@�WEa���c7شN���L;iH��:�z���o����N[�.۰�\���
����n���d]@�<:�ꃖa�w��B�"-�#=Fv/�ͧX��F�]��{Wè�­��)�˂�!γy�kn���JR������.-��ӷJ�f���ӫ��)g�>n��Ţ��X�yӮ�%b\�
��k�
4�ntn����g�6t�k3t٫
���v�Қ`�V_�\P���,C��w��S��t�PY��SS�����a��^�Qb}����**�&����O�/��x�y����ӕ�/��(]u�K� 7NW(,L�O4��^qÝ�: TDP�wsE�\��ha�S��&�9�4W.R@{뷝tr�xY�$��e㻻b4G����w�2�0$�/;��<���v��),x9)s��΋�E�n��ݻ���Rh�<�/:�"Dd�(���!Dם۞<��t#���tHi�DG�sW;x����diΤ��M)I���^v�<n��u�Ɋ5��!s��wvyֹ�ܺs�36W;ws
5�4/�Ly�3u�ї;����ήk�] ��T��l��
(+�"1�h�n��E%@K�7* �������R)1��"���	;�x�O;��@��\����O;�H��2Tn�bHc!�&�$��':���"_��߷�}~}}�~}sj�^�lgS�a�������C��n��I�K�>b�������nG)�e�h���ݚՠ��8J�;���}U_};|��Ⱦ+�k���f���U<f��<�V��2��'g�C�2���JB[��V���u*'�j"y�O5�Kճ��#�ܧ:�]eT[�G���{0�<�ml�띄�0��i#I4���c��x���}��K��ή�h��Ë����V\�D�[yW��Ť�yb/oͧ�^'u��J��U����u��i�d:�5���;�W#�q����ٖ"�%9/b����e��N9��ǆ�{T{�����?�xT��wݹ�L�	���sv*�Wf끒�OE<gjR�����5Qf:B�ZӁ��g�b����Ws��#�[�/[�gp6�6ۚ�2SR�1�8����l_2���򕓕e��W��f3>�z�B�'lT)�#�\��w����O�\`s���y�i1�	Ť�/_*�S}�S�OǇ��1E��U<x��*v�����`�&0�˾���%j�pҋq���Y�/�w��n��o!#�k����zF�~�M@��9�Yڲ:�˙]$ؒ�����o�O>��S���=�ɋF�a�{�����=� �[9\�O�Z����[����{WS����M�����ꪪ��ka��������V1�>�Y���]5ɭP��N�mhU!���<�(]�����-����>����+ұ��kɌ�Z�zq	��ŞLl[�{��'c
���w���D�;���7��Ğ�r���}=�>qD����0��%{S���g�+��w�&y�mU{,�p�6��Y2617��e]or�֒3C7��q�Z'/x���r���k���{u��moIq��۩{���R�.r���F(�P}�\Q��)w�ڶ�v���w�7����D3g�w{�o�Dk�mgWi�ԴǺ_r#�r���-	T����S&��Ꜿ|.�nO7h�,�)mUfzq�j������OW��v�b^����ݸ���;�©4C����a�?VB����gD���My���_^�6��[�\��9M�q�V�����@{-)ͳ��7�%��v��L3�m���8^��#'�����aXt��{�2������)���Q��t�S/Z�-ݕܩ��L����
�Ȣ)-�}C��N9ܒ.=bj;ո��[M��t)��sO:��{2�R�hrU�rڊ�n�{ݏ:��Ω�N�f�='2n�j�U����������o��r_�W����׻6��O�Ȟ�ʂ7�o���q����R�M[�Egr\���kÞ>���;{�3�RC"Up�V�`�������l�r��11�H|E�5�9E_b^{�����PM��Y�nwb�fO(4�g�e�u�1>��-4S�����L+�s��ڪ�-۾��
��$.(��V�H}p����rY����G
>3=�m�#�v8{�ELTrq�����ȞvTi3��w2�V{ [>u
ao�S�-�r{y��?D���x�t o�p�a�Tx��zB�#T��B�X`�uT"�:�O����te{5�d���=��^2�����w�q�A̵�Z�L�.��Y��}���UY�N�V�f��E���:^V�,�b���p�>Fy�԰�l���\9(ꚛ����Z'^���=�
!�����]L�ڞ7МΛ.�N�$��������Q\,dśQЦ�%#�@��";6g,�`ݧ�˿b��6*��-���a(�f,�N�Wu�ӭ��ˮ���mG�:�ۚ�."�y]���N��憒�Z$7B��u1�6t�y�������А�w���O���m.�8���xg&�k]]��{]_U�"m +���D��T����Ps�������I�����U
mT3/.M�J�QI�1�S��f��ۼN�L��\��U��v��H�,i�KM|� n�!tB�ua�K/V��@���!-^��Z$ߔ�=ܹ޸TDE�L�|��`y���ܿq�}'�������(c�{\�ޞ����sˆ:��^o�إv���9�g�M�}������$_3C�Է>�̯�/�=4�
��=y���:�3�7���zJ��A���Uc�-2mi��oǻ�8Id�WH�7����x�p�p�M�3Ns�K4zB��1�kfST�3�
jFH7��Wau,ԅ�q��u�
�q����SnjH}p�-4HiwQ,y5��j���ƴTk|Zϔ=����ޱ���]�9Z�"a�f�Uٶ���̽�
��Yt�ʾ8�V��۠����<|=Zv�x3q�m琍��(Q��q\�B���H��K���˴�Se%��泘"3� �장����R��챿v�����oH�w�.p@O��=�"��;kh��;���#��v���������񙩱�D�tױd�M-f�T2�i�چ�5���Cu��uJk4'��.���m�U�!�d��,�w�Ի�vxJ�z��R;b���sݝ��om]���w>�1��Ok<�j�ϥ�"����̂�֧��d�c�S���{��.�	���"�8I���\k�=L<�Ր���oɘ�2t?c�)c�j��{��{�륅m��~+��kI����ٯ�R��?g���$2&ߓ��puk5����y�j^��x�_oa�5'����6������ZΞ��}Q=��_Tb�i#^I�~/�{�[�,Or��sq,��Ҝ���T���μ"�"e�ʱդ��E����ah��t`Me���v��·�X[�!3УN���檹W��c]�R�
�%�x�r�}��U���amT��ƭ���Nڋi�T&���g���W���DάXB�3X�c=�Tu��iO7��Ӌڇ٧Ey箮J�"�7݀���B��H�V'\��;�O����WF-�Mb���C�ή�$���i�_>�j�5��Wk��In����}B�י͋g�������̥�����D���33;�ﾏ���m�iK;I[5�r���傭���Jd���GB����=�ٸ&�wbW�k���|�KX��/���l9�4�J�j�Wc��-R�ܻu�{5�Cx\�W�Lf3>�z�aߑȔ��s��a�X^W[����j��a�^�`�쫵��.�n7S��{��=@5_ro�o�M:�շ9:<�˰��|��rś���_W��v\ކ$�T�h���~7�{��bڝJ����W��~����D�����~YK7�|2Bn]��3�u�C���E�WIPm���x�i���3bo���Os�����)�c<�ݼ=�λ�,O~���i�<"���x�g���/_�~�3\ԇ,{��+Ӹ2�;Z�8ꊃ�t�zx�^+��a���7rj�8T1N���9H��ʓ�2%GuF8�Q~׮*.W���6������{4Ҝ-l�ٽ�f_Denk��⡣_�GSR��5��z����MT���zĜ�߶{�kY���~��DQ3^U�${p���E��z�Ni�|)�/!q���NA7���x��H�DS����.�I��M�uյ�t}����ﾮ+}2է�泦T����̬�D���%�(ȴ���}&Lc�{
� �{�ڽz1p��9��U�@*�Z
��7����Z$��q:LU�Dk�{�ɨרH;4�r匼�~��Rh�ХD��˒���,"�;��-�Wm���.Y��e�K�!p{P�T7M��*��Q�*$=�)xn;
n��ٷ�7�36Fj�b��<�w��b�O�'�����պ��r�
ƹ��z�5����i��ݟR�?h�]�C=&C
%R�g����76oWQ$��*�������7�x�cڎ/B�G]�'��ɿv.���wql�[֨�Vс�=�?D���>�Zs���H��D��r����k�W�7�Z=ظ�N.'�������r��sg,{��ٝ�:�ܒ9�c3�����i'�ʍq�΁�j���;��'q���zt7���� �.x7�s�Kٚ��;۾䳍`�a6jJ�y�S���%��&�**�������eCdJ N���hb��ކ�h�֐e��j5����{N'�;���/�n�Ck#.��1_5#�]au�P���}�cS�Z��U��_R�����&�a;�D�q��-��\6�o���|�*�^-X=���:�SQH>u��^vw���l�����-���?^�W�S���rΤòu\J s�.�_:4AZ�B�wf��*%���[�\u@�m��{Y���۶ʓ8�=�i�{��	"�SQs���{Z'^�����*R�R����^]��E�6'����],+��T3*jrz�Bꌗ�}�
�n�O�z@+����x������������!TB�T̼�I��9Ϝ��Q���'{��k�OxtYG�?*��p=��}�W��ªD*R�	�V8@��PQ#��y���q߰I�vқ����-�����6�꺚٭r�嫵�����E���]K�9��/��;ޔ��5>΅�y�8AR��ީ�0��d�=ܳ�'��~=��+��3�nsߎ��Y���w]�n1��.Sv�+��k�дp����YG�UmK�(��9��t-�+.��3J<�:b�uuy�[�Σ[5EǪ�Uڰ�cr�b�5���&MшP�vf��.֠�͊
�w]��}]��H���^v�Nd��Z:�fbM�2���T���fҟ�_}UUIi�]�ݳ3o�7����ĕ�y��1дߍ�5����%ꁝm,��w\�>��X�V?3���6�+����R��lC1��6�r�z�Ы���2���1_s���)y�b;��p��w�r&�)M��=!��q�S^�����Y��	�i��)q�ǆb�0jq�ќ��q�>j�Ԭ�!��պYQ�z%���g�@gq�!���Y�U뜫�׭8M�;��i���a�c��M�-�f9XJ���sٕ+W���Z�^��Ԅ7:�2��O3oVp^�"�ߝg"οH<�v��W^�����(��>6���v`�>�ڒ����W���<��5x�j���~��I����p��ܴ�Wm��=�k�H��r�+o�[���}^ƶz���9�̩�����(��j�/�vףt⃫Y<�qT�q�U�og���$�>k�$����'�\�:���7�ck1�b�MqTeLW�y��z��ֹ*��.���������Q�[z,�2\㑚b�"�L����gEƠ#i�V��>]��뚬��离��t8�4ç�-=7R�i�V���2�
�g�����Q��DG�=z|�-Z��4R�ěEG-���I��w�/�{�R���,�Yxا8�m�:��Ѫ�`3j�=8։ڽ����ˇ�Z��H���yr-r�=.3��ᶇmW(B�r�cN�P1a�g�����OtWe�/:�Y�M!���W����u�ʮz&�_3����:%Wnxu�i�\��o�e�w,�iNOQ�A��u�j����z�1G:��P?v���z��f-�hZ�gpT6�)͹�S%ST�8�tȍz�M��Uoh�1|d�F�cW�nc=�B�#�;G!:`AyY�no�MK=#�]P����Lc
}�&}��5�k�l��Ҧ�h\�Or}�|�j:�}�=Bm�]���摬�,�\��~�$s2H��d�y�{a���-���'�4��'�ߡ���D��9y�~^��5���,g�%:�~jr�=*;�C-%i*��>�/[�J
��*n
�h*vDN�8\0��
]�,_h��a#�7D]�Z���䔘 �N�8�ͧb��h78��t�L��lHJ/%NN��Vm�"p�O��74l4ъ�]���1�XE��'�WS\�&���h�8�%�p'�J�v
���v�e�m�3��%1����%XT+z�]�H�׋;~U�W6���<󭶞m�i��ǽ�ֿe\�)^�y��?#t�_x�ICՀ�U���]�6v"6�bP:[���tŲMU���Հ��>�h!y��o;t+2=�/��Z�Ke]��ƅM$��6�.^��!�1i�b��E�ؙRQ�(8�b#/.�Ä�7jD6�IKc�jlH�syWuMg>���;��h���qbH �r)^	��|A�ir@���6���P��~�ݤ#7ݓDK�Z�4`g�=��b·n�̖�B���Zkr���u�w^��w�vx��ݻ*��dX���������ޗL�ma�Z���`RU��<�z�G�9G���j��58�a]!��׶�u��S]ڭ9Y��6p&�k���;�Vc��e1�8Gp���m��%A�ej�Z�-��J��_1)�m�oz���'|�!0%�]�[Əf_%+�yq�/���S:�	-�J�:�kA�Y�&\��\�-�:`%�؂������*N�̔m�j��c��N���w�8t<�gm��XyA�g1O~�N���-^A���A��ZcI����ؗbŚ�`'��>�DnT�N���	͖O(Z�x+9ޭ]���T��*�M���ԛlS/�]m%Ft��k�N�jʚN|��n5���-}6�F��s/f�@����B1r����No_
W�����ԣ��Bcr��A���G�+k{��iV��7�U9F�w��r!X�C�ü�`y��Xu�*��R�p�Q�ʖm���DE��n�]:����C��eO��v��{6��ۭ6�^��V����M��\1�!㳤�����&.���)s�+����sg1ֆ6K6�"�a
�Ő�o�BS�\]�:�6A��K�9)��22D.�7�V�3e����0k� �WE�-��"�A��7s���zh��I���3v�&M��Q��}���sެt��yV����t=:��r��m!�؇`d��f޵a3V��1�i6�P ���[ǎ�@>�{v�[����q��	_KYQ�|ok]n��951�s# }�N�NLT�Nl���v͋�[�fÐVP�1c@�I��P��Z*v�tI��@�t%�qZd�Ě��j�x�CY3L�Ä�jS����>���5jQ�DU�}���݀Z�ŵw*8�K3,�{�p4(;IQ�ٙ��#N5�S���ʯ�(-�Y��Ѵ�";J�'�����^�ۆ�+���F+�&�Rt(�Q�w�]Lj�WO�m�6�8���{��4��
Q&�C�H��7�ِ�;�1�v�û��I%t�,Yw]�"9��<��H4PL�7+�fd! �	�6ba��tQ� �l�x�RM��Dc0�Jh��kκ�u�LM�M��"d��L01<vxݤ��lBL��BM�.�dVL���!A.�
S4���Kx�� �YCIx�ݹ&A���)9��rEΌ�BDP��D�%	�SI�7% )D�QAs��n$�"��%w\Re!1����d	y�7.�Q�(�Dd�� 1��(���&D�	�I���M$�Id&Ie$$�a]۳	H�0d�B  ���9�Ζv�o׬���y�����1*sv��'<��o��T�hg�������Ȁ���O2؝/��d�Ș^�����Z�\�W�����=���(e�U�5_��dBˑ�o�6�������bOݷ=��K��̓���'���xE�O��D�<�6��@���n���/;�}}�=Q��凸n.�|���ڡ9x�{��)�5x�k���><�U�f;OiZ���H�MD�-�����Q~~���M�j���u��7k�= �p��o���J��G�*Td��Pm&USHKV��1����q����^�BoeKD.Sj��V]����1�M]�]�����}@���Mv"�����/9��*�D:�*&�G�jP>��wv5��OIЎ�۱��ėnB���q���,˜��H�m�+-��{!��IOn*���޹+t_�xL�|���}R��'�@$�Q�Vt��+qs
C؟L��u���⵬�gpTCl��fmэU�tD7�V�+A�<d]O4Z��VX68�qn�Y0�Zn�_F��GB����*��]3y֏<���x�.b��,�@�U�j�>ka��͡l����JĐ���e*U��[���u6�JX7��Lt���=�lު[$�C�r���G�������� d����\ʾ�>�����1���Ё7-�,���ף���s����}G��S� t�+Ev��{�У�c�&wk��k\���X����W��h�LBqq>�nh���@Mm�ʾѴ�P�[I ���̹�t�]�(�w(�q¼cz5��m�@c��>4��[n[�9?NWz��3Y���QGx�x������dj��"���ه�ԅ��2�_b���V���ʕ�1=��Q��s�}�Y��z�F��%��y�z��bĆm�k��e�0�����b�O�������#W��������Uٻ��"y�oR����>���Y���Xqnuzo˨Q�q�FZ�Z�Y׾�$�^��x)!�{|���ڥ�yoY���W'򵮗Wo{ZPS������=�}G����~��UC���y並�U��C2�TtuQ���HuT��=缟T��ǞHp�6b,*Lwj�҆P=WJ�c˱�C짭=�l"p�
粂��]k8;9P��&��8�lX�qM�e�x��+�!\��%;��J&��ñ�)�(��.�ʻ�l�yѢ2S�8Qק{&�-��u�{�}.��{F��磌V�3}��煿�'a:�/�1դ��i�D�����nI��P�w�KZ�ucRz՗%����Q�Sm,�ZW�j�+�t�F�br�M����po�����ڵ�\�fN�j}�K^��M�nUg�k�k�q{Gﵻ�C�|�������C��	�5��j.�������A�K%7�w��`~���:�4�Jk�tY��L�Zj]�g�K�zb��,k��hP�����hV�1P��f��Y��_���Ưu�:N��7ۛ�YY9Y.�O�X�{��W�Eƻ�r��#H{�5�kJ',�|�:�;�þ�pe��|���j��&kS�q���� ��Lm>s�U�Y	,�d�*���;�n�%c��
��+L��u��P�Y�Fy��w�$��o��5�����<�wm���7��D�!y��M*�/ �gIn�Bӱ;y�Q;��K�Z��+�f/-�諨ù�uV%9�}�c��`\o	ɓe�	�,��rxͼ޻�΂�I���D��1�۬t�]唎�:ލj�՜��|�] �;�cG�[��bWk�Ϋ���܄��-���Us�z4At._~����VjN��8����?c߫ߏ���o�n~��Os�֮��֗�x��w���'{�|���r��5�V;˸Ovwr��#�5s���L�����w$���Fhc��ŭ��`��m[��G;��/s�w��}�G���wzyy�V�ikZ2T�K�^��>�q��Q�Yȉ���Q^�D.�?G����h��=��8v�#��"����\�ꈕ��_V(6�)4�|�e��J-÷�f�gN_.Nv˸v�H�ъ�$�T��qG�c���ދ���ᯪ#���{��	m��]���;k����v�ծ[X$�ݜt�����}���p6���n.��n[����﷝T[J�vR�M��@���_v��/G�=]�Y��/��;>��U��ʄ�^k�������S�%^]p5�%Ȭ�i�{W
�f���w6�*�O�=>��Sb��K� �Ϡ�B�E�["<�wqn�i��K~����=�=y][W�"a=+~\�8�_��,>�@[�:������:�޷��T2�r�Vpqs��s9�dV�*}�7�<���ՁWB�|z|:Q��ڲ�2��[���ﳢ��x�����S;��Zc���ٌ�w=
��0и�\ZV6tԬ�Ֆ_,�vtښ�R!=�񓏲�-d�
}�&b7S�����q(^�m�v�hV.)!p�\LqH�2���?D�{���}ި�(o�+�P�oJ/��y�p���6{�o~���F���7�v��D�9y��\�4�o�:����f$���ԳN�sT�f�g�f����� +��W�����]�bl̓��~��-)�T��j��{'���xCK��x�jy�oV�,t{�{������@��/f�np��o]q��;n��j��U��"�]�J{qİ{�U�nۇ9�999R��(��(:��A��bW{R���w6�SR�K�%�z��c;��)̯C2��o�%B��"�j�	o#juD�׷�nip���.�೹7���!T)�Q�V\I���|������B���-c���1��X�j������M�T �vS���� 	�j�Ź25�4uQ�"~6�gh�~�pL~v�ޑ�%Nq�2�l�-c���n�(�ve=I�U�^c��ue�nB�k�48X5ˬ6��aǖ6e�{�1vt����}�� ��.��7ME�F�2��Ol��p7
M�����X�y�C����p����.��ꞩ�cK���r��q�V��Ul�f�s�4�kC窧a�
ȑmT�[2��d�'��-�b�D�Gq\nR�Κ��UvW�m#}�WA#��/��ڕ�_!�Q������֍�����m߻�i��7���|J�T�����};_Oh��kM@o�/�ǵ l,��ٽ��FY�v뚵��c�9��9	ӔK�=!s�����48��aSޅe�Wc9^�B�~Γ� �q���N.'���=!��3����}"�q�1�/���[���5�({j<Z�^��~5\1?Q�Q�2Շ���m���&��q��f���ƣ/�R����~���3���~��x�^�/��U�s����-?bHyY=���[������xOp��0�x/P�Z�{\��kz�<sE&:\Z�Z�39��>�i�ޜ�m+*�ڹS�Y����c�0�������׸��J�x�Zs��4x�J�v�gnn;�%w	(��+t�Y]f�����Sw�8U��t�sd���ri�68wIۜ���_�̞h��G���p���p�t��&���(>�z�#���A0�@�:���zf�{�g5 ������x�k��F��s������ԛ:Ǜ�M�9�&b�`;��u}��C�ɯx��Y%o!�ױ-��F�r��ͬns{�#�8�K��ֳ^�\����V�o'��!#Jr�P��MY��Fy�ʓ��O�߫%N�BM^ܣ��{}����/9��)���I!�&�Eԭ�uR�O%�뼉*�|�rQ�S�˅���Xl���a��릵��d��azcx���g��Cy\�k�5>����+;Q���-�bk�剬�m����{�^�Q1�ċ�j-�l���{T���Q+Y�q�訇��:�(���Uc��0mi}�ѹ��r塗��e�����3�k�^������
�@�BtOnB�WnoN/0ߢ�{Q�m0۠d��c��MyK��J�8�����T�A%E�:�)ѣp�u���o�����g}�xg(�&�֓���nC]&h��#*��8P54��N(I4��38�)��l^�f��.�����L��Q�q׺Ԡ`y�^����+/y��p�T"y�;"�)X�sАq����v�B�s�-ig"^��Nkiv��%@<� n�񶲮-f:Y�f+S�q���s٩�Wn�t}�VM�＠��|x���!�~1s
�;�&2ik7�z���lf��V�b�S�s��9�j�[̯D��ٕUa��ܴ��z�]��o�[��yRq��N�޼�o'\�˫��K�/�����|/�]��n�u���\����'�6��'��6��z�˗�l�k:��ݫ��K�~�Ѹ�"-hת4���<ގw���],+D$�1��> jq]⧶�z��ͬY��ut���ƭf�˕�O5�@<QymJ�i#��ypUX�T�#��@��Z�*9V���ZH�M3�m��s��}���v�|;i�x��l�v�U
TO��ˈ�|O���gyߜ��k�^�<'�A�ߔ��s��F&z�����ƬVN{Tl�V���c�:�r�^<hp����{�VT���vy�`���z�`V����Y\�"l/.�Vǐ�6�]7]��zoh�
��B���)Z�XG�3�����/�����]���P�~��{m4�;O��U�B�C��P���Os�0�x鍙�Sf��˖]���LBֻru�y���,��oQ�^��P{J���,?_nVN첔>�����<���w,���OQ�A�o��N��z��s�+"E�j-�Y�4-m��ᷱP������n��X��ܓ�x�ۉ'�P�~�0i�_Z�iW�xI�s����_Nţw⻙d���$~������f*/��ٵW�-zG����,�4a���Y�//M幓z��5�9�qq1�����ɝ�s/ҞMF,j���;��:E-[��w�g��I���9���ȟk�g�X|-yԉ
�}�牕+����Y;�,Tt�^�Q�b���gگ�q�$,26����vH�T�����c��R�e{���Q�`��z�5�=q�����J��,-����y2	B6�t���A]YY6�!���R����3�����vQ�4�|m�G��]�kZ�]9/��Q���v�JH�)�]��N�i�}��y�n��A2I��[�`EM�[vx�%�:�<ֱ��c�X����/��(<��T����U.��z{̳���s�ɳ�-���Pb޾�O%��9��S]�3�XҖl�zA��^�������9�`���¡�⎜Pc^���z�,]^����EԢ�摑xM��	�j�v�w�9�̬�I��P������@b����+����LZV_�$Ô�����oe]4B�Sj�eeě��C��}������+����u|�N�/��^�Ci헜�nI�yJ�J�7�72y�̥"L����w�?n�ڬ���gB���q�征�W��q�cf��d�糼������_G�;��:��*�ȟ������kyU?���};��SH���Ӵ�L����s��uv目+ZЃ2�6�Õr)ŵ���ݬ�S�
d���5;|񵦃}x:vz��"ڙ���C����^�n��a[9	ӜS.h��Oh|F.����=d]
�힊g�~M:X��������h�G�ڒڳy��DDj��ކ��i�J��ɷ���ޭ;O�^�i��qc�Or��F�����NW4*ꎚ���/.���VOIC5/j^��<�J��7i໮�n��)IS�Lu�O�o
��x^�Dˬn93���Pw˵�j�'r �EN�������DUF0VEW�I��/�G�R1j�O�]j����/��$U��_gK�V䧽�ҥ�4`6��}e�m�t�DLht�3Z���pko�pO���"�
r��
��Y�w��ɯ�*�Cbi���j\滓���Ci��ſr"S����Mr=G���#��znx�50���]���.E��s6c)]�Hk��;�<�渮ﵰ���Z$q=��&���!�w�mL����F�f]
nWH�.��[��*ő�����4�(�]�-���}N��N�YX���z5��x��Od�C�N�������6�9ʴ�j�ŚyC۽���D(:��e�iL���N�ሷ���A�E��;������O~�ꎤ�[�_X�p�����WBj��\g�-�u���ז;��m
���m�zb{̛�����Z �}"ŉ��}��;�F:(�Yڑ�pG�w[��yy�"�m��{5����%���m�#�$���]xS��C�_C,�X�d��b�8� ���3�J�����jܐ�Pdk!�.��kb��9V9SnV�],�����c	�0��]��Π��˹7ֲ'�M�f䩇�+s�43MD�M3k\#\Xi��m�^�u�3F�Ý>2��E8ޱ����Wse��j`�����]�zI=s;.��Һ��zN���)��Ա��7�Pg>V�3c%��Q@��u����I���[��ft3���=}��h�r�7ղ):m�7�� ��=w6j���6)��k!��D��kx���n�Ռ؃^��*b�uʛ��l�oQb����E@k�(�j�-q;�t�]YUb��B�o!6΋i6F��/c�jo��de��X�܇)�%�`�E���[+&um��£`8v�q�Ed3m]5iR�w�P��Q��uk}���HC�T�,!�g]n����7��ud�,��->���f�V�%2����β�9����tgکYb�uA�U�p�;��_k*��of�ڡ���|��7i"BW��Y�I��*B;O;��T�{�M�VQ�t�pK�XL��Y��Vs���nT,�u�3uf�6�c<���	�w;'�3��^��\3�-���Ok� �UC��:����*�������`�wN�lpz���]Y��[�l���X�ۧ�u�D|�)��F�bY%N�v�f�Q��۩��>����64N2���f�=�"5�_
I	s��U�F��ky��Iv�Yu�Eam�;�|]���P�}LE��XB��H�m�u��-���e�w�a����������߯��?]2Y'u�BaL4eI�IR5%2���w\�u
3b��Ɓ6d@���"F%)CN\���##ssn��))��(@�L��JAE1s����`���!DBh�hɢ�dܸbFƈaD`#(J�(24 b�Ȅ	]�aL�,��F���C�(���eAf�R�$�b�)"HD� h��4���eD
��F�
RHي0bH) I�d�A�.F����c0ƙ��(�@�"2	�4��J!D�f#4�(SH!LĄ��$�!���7wB!&HH�b� �
�
 }B�(G#��,}��V;p��Qѣ�e��'��|���^hy7+�Z@���'{����u�Ú���t�Mftr��˹YJ����=}Tt��	��C�3��W��p�D�qq1��׏H}`��l]����s�^�ԅ�nڏu��B�t ~�Q��W�b�EF��̮
�̝�f�[��o��������/3��7���Z_����~ntN�Z�Yqjm�٬�8��e��]��ߦ$���kj�yʠ�ړ���Omsޣ�=Xx��qA����}�:��������DM�T�2�A�z�[,�w��������u[%>��~��������g����ƕ&�5�2l���8�f��Uʺ���?3|65���W�f�{'
���1�Ys����zn1����j���|����P3�'�D'�=�!s�j�y�9R��e]���G����<W*�R�����	�'�}n� �n-�̞�����W|���Pq�QW��U�)	�^�=;�FW�*j�ah>�T���Q)D��>����ƞ�V�0Z�
$��W�)xPy���Y�f�H{���;��h�w�S�j���XГV�tU�v��1�����$��2��N�բ���̼���u�%��J��dh{�_�w�awu�����<5�\dm�"e�ǢW=���V��)�=�^��a�+(�+���Gh����3��_6�f�cXuw7��l.�����gll��nR���>�'c�w�XD�*�iL�Ѫ�\NR�\���U�d�"�T�K�&�ǯ�or�X-	P��⺜f�e�M1~QS�\x��1+LLO��TO,���X*\�o��Xx�!���N?����B.��{����Vۻ��ȓH_�EL�q�fx�Z*y<�'�A%���U��=V_������,�;;<��*�`[n�bn!�;�t�����eLeF�=M\�=�ﰇ3r�{�I�R@��_�J�X�I��t�)���2~O��/院�W�����
�ry�Hd����z�����Ԙ��le�<a`�t�;h�1��p���ȹ�v���6J�o;so�Q�p�2�Z�UY��>�EU��q,���6a^�p�?oow�P�P�7�<�׼1����������Y���N|׈a	��|x���xd`Lc2�Vq����ݲ�{$Z�z+0E�tcш�5��������;��C��E���/��Ĺ�d�׸h_bN~Y���E��*s5�ێ�����ޱ��c{5ߧ����JyXFf�0=�|����(�@��:]�y�lo	Ɂ������9\i��x�X�9*��{�jl�M���1�	��X�����Gd�,'����l�+9^u�H���2�,R�Y�Qە36�C`>���4��Ρ�7��3�ɺ�i���f�W��z����q��h�]ۅL��GdN�F$u/:5^��Yν=�e��˸V .�d���/���ª��Z��xO
Be��s3�1��Uk]K�
��l1�<��T�^jh�m��h.�[fx�T
��N���^�d(�C s�R�-��݃ڜ�R���,����6�w�ҧ�O/f����R ]�3��ǳ�Uu�lX�u�;xQ��E�n�����Ӟ΀�/�t�T�*�3�W}�A�v�i�U!1]2�F�"���*�ᙦ-�C;�n��n��k�O�:��F&��dB���+-��!���4Ŭ����]2�}X�v�Ŝ~�NZ����X&XTЫ�����rЮ��߂gg=	�y���pm:4Ć�6mfLϵi�{��r�ȯS��N<ʒ���z+"$9[�S��&��GXx�l��ɚ���O�u�S#U�>pv���ҫ�쪞>5&+ԴU�#%1q욅�N�Gs;!oF��p�K!M�~���r�}#\C&Lr��
�٨Ȯ$.�:�����5X��ǣ�`1�j�r���E�3�6i�pr
z����Y����S|;*�xr�� v��MI�˞�0{�.�̕����[%�f��V�o����Ѵ�ACo�wS�݂z���h��bÂL��tT�����۱D�&�iMѫ7H�0�Q��_G�Uv"�4�(ut�#-٣��zZ� �ʯ���W��v���V�.933���1�τ�F}]d1�����Un�AL�}/���cs��b��,?�l��-&��иJ�Hێvg/Y�'�~"���D��/#w��0�@�z�{����/��n��z�ʞ�yq{Y�UyU�[������N��C[�42�jQ5x+_�u�z����h+�/9����*\�m)��:;��^�te�W�קv~��M��(�>�'>���{k0�cT`x�n*ω�pB`u��L�}���V�7\T�x=w��'�Ŗ;��y�}=x�xF�#�6u�{��FD'��_��x�،̫�,���~�{��,�/����=�;.sq�R~�G��Z�\�99l�(ꌂ�WR���y�"U����o7��N#����e!Sp�)�E;*_`Gx\'OAC�ѩ
�J��P�;ƣ���[�y��e^-�Mju�/�1�\��������7�8�~��4��J�r�TM�m�b��]A��h��j�� ���<���\�h����6���ݻ��2���2t�?lR�X���]՜�ý3���U��JH=Φ+�����]��h�UǾP������n��Z�5��L��q̕�[/.��]�]'(��r�Tл��u
.e<!Œ�Y gh�X&<��|)��䧽skfvG�Θ:������ܞ���"#��*Ҽ��7_���yB%;�FI��oᔼ.WJ�苺r� ��!S��Gq�i�jx-Y��{[ʺ�������O�I�Ӎdӫ�ʦg�_�O�ZbO��LU��Z<FJ�,tz�.꓇S�Fnς�v<�Pƃ�ë�&�o�vm�h�AM�VCU�Bx��b��j*�C}\�>��s���2�j��g{1��p}��U-B�����)�0f�Yĉ\��ĺ��8��oz��_`~]��8rſ����m	F#��~�N���!3>&9��.+����UV�0*j����/Mˈ�&�k��S�1��\�v�RoQ�UiS���.�\a��O3��^�. "�ۤ���項k�N��
3��k�B��ѥNI��7��k�B�Q�Y[׳�!Qܥ�zo��՞]��f�ϣ..��F�H��7L:�{à��`�	��*o��	�6yo�,� ����{u�g���]��~���y>�s:`�2G
��>'��.0(��fQ�%���xV.�1�z+�L�RGn��oDk�O\c>���Ov΍ʧ>?1Ǥ��5UXϻ<f~J�=�48�QjTkKƩ^���kbh��-��~K��'��e��32i�H,��q�ti�|�>y[X�γ�i�Nuw#�����	���)�b"�J���`Ls�{��yυ�k".�jQT��/�R���C:t;f}F��yΆ.���)J�ym�1�u���V��+1��V����j���|����k{ ރC�Č�
�j���{>e. �(\�c��/���G�����ʺ�\���W�"�7�x^S~q^Y�1u
J�O(Ǹ1H�p�{��u3�(OOyў�EM_�A�2���d�|Hx)Ȋ��������w)�a�-�@*0�gu�HV6S�C�Uҳ��}�Iu0�S���u�;�q6�����T��~����3ʭ�S&4j�9K�\��(�.���1�o|�ɧ���O�^�S�nq��b���Li�V��k�B�h��w����v��ɦ9���g���x�(����%O@���ⵒX3��H_�EL�q�f{5�[�"������܋�勥�#�Y5�k�(�3��q����U�ٌ�ul�QJ��nf�m���t+��_�����O�RGq�AϮ�q�D�?f3Rc��{�)���!q�-�Xd\O{qU��>�T�ֈ���D��`��MI�+)1���Ҝ��4^��Q���i�����j�br�B����,2-�x�p���2���Y�ǲ�����%^J��E��c���Aq.q�R'���Jhas�7}f�,�Orw#��·�д�c�!5�V_\����+{��&/���W����%M�4����Þ���<�w��$u���7��l/�Q��q�R>uW��>�EU�聧0T�����Yʚ�p)ɸ���5�~W�~覰7�fz�����ݙ��5��w��%���PӲ���4�㊐\p�U���מ�%,X��hW`���:�*�5��Y�����O��i=�j@��N��t�,8��~��6kF���R���s�e���w�k�n3s���*׿M�$�Տ�������Q-��UK�ޚ�j�x3��u�3Q�vD��bw��׾�����#�zx�Ox�^���z8�
3�:�o`���A��e�T{�pk*�R/{�.f{L��q�.���nv?f<>�l{�Y�������g���8$k�\:*�=W�\A
'�����\F#2��"�N_�-��g�/�=�Mi�Hz���{}7����� %T�r4j���uE�� �ϫ���}�P;��w��� ��Ո�����@g~���B�g���3�4�2&w�{�T3����vvWo��ʇj�:�X�J����6�`Z�o:�Ỷ!���4Ŭ���.����}�u'�m;�?��+m_BjZ�ʯ8�BP]��Q�j�]4�	fv=�΂,
�l����a��Vz���Wlַc�G���P���=E�Vg���D�{�2�;�iesF��h�w���[2��Z��`���\�����(v�e�M��K-g�Ӝ����$z�H�6��U�B�iٰ���D$^�y�����b�  _��U`՛�v�
u��:��W�fzHZfLR�W���@��N��R:�r2|j��
(�|7������y2���UT�>J��<7��ԟ�ԴUČ���욄~�.����ؗמ�ݼǤ��%�q����ɒ��ȸ�O����$.���|b�Uc��������f;���w;۫�ˊf�@㤀�|����@���g�Ls>�E�Yw��ە[�'m��9��e��?IѾ��W��hA��д�č��fr���2u�������L����;y�#QѪ����KM���7�Np�7*o��{Y�UyU�[���w�s�]�X��[��_�W!���ָ�wDw��e�Hˌ*\�m)��:;��Z�K�����fC��u�=k�<�8k���u�k3aс�B��V����¦g�i�uV�;=c\�����}�|R����Z;#���;>#v;Cg|����7	�pB�|/��;.{<�"١u��,$�_8���+��_�]4=��J�F���dj��Y9;��抑����������N�Rj�{w�
<�AΛ�[��{x:a�ۉ��z�S<�fWZ�E��f;]�/���oae	�^v��ţN�T��v��蚋����hX���R��7!�R��#�����D��������:��H
��q��[���������בLT��2��;*_`Gx_���P��jBB�VN�@,�3��@�uj���|��[,��U�=��ϼ������wͫ����q��Ai���Y󺻷&�/Q*�좦L��2hcWO?}f琳�rq��n.!��xzkG�wO��~Ї�_W_x�+��q�%a�/�"y\:0�H��3c)x\����]ӕ]Y9Qz3n�dy!^=��[Dw�=���[v=����v�2i��T���T�j�_�w����e·8�N��a����9�I`����T�H�����6��I���A��;Ҹ������_8��g��k�����j��fMC9��_U=B���&S�`�"K"���C�%���o�K�����/w�t����~�@�m	f;	�7S�����@�ALτ�;�B���>����.��m�����
?ׂR���e����}.n#����˪�J�ο!pp,���HF����0e�X��+&Ѿ�N3-�&�dh�®Nc�#w"�D뾃;��W��)���d��Bv�&̂٤$@Ux��T���ą�4Z\�zV�ض�3^�(R=n��T��f��ɽn1y|)��W����{þy���]�>Ν��H<��r���OzȠ㗈��|�~�9��X�4��1�ʛ�G��fP�3��y��:�t��\�N?������pUj�"���0��d,Jcc�)P
�2&e�͇�Y��{��L���]�gx{�d���2���k�cR�����2^��V��L����J�>�;���K���![�f��=�.w�]�z�`�O0�����Gg!22�ǏZ���Ǚ�z_xd�9S�W���ym��Z�N�+Lz��9���zn1�����(.��f=
g��{o����O��
B��7�(��W5������ʺ)U�}�^��]y��oس,�u��ގ5�Pw���E������
Bg�����nLG�*j�XZ�/gL�Mg|=&�����Œ�vç���D�b�� W�
$�7U�x�^�s�z�U���r���T��?Eݝ���������{�\ﾊyj_�k(+�a<�٥2tj�9K�EpL-gαz���ʱ[�yܷ��ߧkh�`\7]C���r�ٴ��M1q�<���2�������W�г�������Y�R.�<ٍ`HR�a:恴��I�V�E�°��5z�|��ř@�
��r�R��V��u)�n�Rp�M��s�QR��ܔΚ[-���kvta�S���x�����!���A�a![������]%zX`^ޭ�//�1hT���Y�%X�����I�33^�To�A�˧r���5ugDj��u>��O�@��h��3*S՟wMQb�B���%�A;P#��fC�l���y�R�}&T=��θ��[y-7�0�-�����{@	0� ��n(��`!��J��nY��� ��	�Pv̅�΋ ��׻j�l���i��e]i�-t��uYRF��Œ���w,cd�x#�L9����ʵ)?��쌗�Y�\�a`h���IVd��.���`ZY]W3{�-&��z̦.�n����q5z��v�� ���t�Ml��ж�vn�/�f�G_uƫ+@Ԩ�k��qgddUˎ�4Hv����i�E�i#rV>y�Cϵ� F��nB�)���Ǌ�=i����/��h`�-�k�<˄u���an:K̊V�W2d�:�z�N��1k�M�^[	b�WwjV�%̉5�|R$�O�a0_�
z�ս�HsW�c�ğ��W*4�K�y�':[-�[8w.cp���8˶#�����S���Of�{���Y3�jG�aF"hV�PX����h.��:$H���vwY��U�N,�]k���W��V�Woe�F������	u��v�ڛW�͜=�1���ӆZ���[�[Av�)l�%��; A�3t�S�A���[�,��O���t6�^W$]Lw37���\��pe��z�K�L��wWe���(���Q���%��|:�x,�0+�%r���Ù+���n����U�Ը��̺���An�۔+p��K����%]�%�#�ǗP<�x��畔� �f��3i�����Y+�7�=�*�cfr��ɴ�=|dZ��\0-`(flS�L�vο��W�jm�ӳ��xt��3�p��;^���F�v�I�*�t֙�)�ۺ�}����Ç�k*�Z�4W:�P��8�D��x�J�J��]q��S/�1�}أ7��ˮ�X}�;�w��!@K���I�p�`��W�d�X2`zgn�����>�n�z��6iM�Es�J�2�W��U�+�F�h �s�����P�V��)�����u^Bֹ�����V��l%���F���7x�`&�z�pV����o.q������f�;��9=��/|�͘h���iذ-��n�SA��V��ΠޝzZ�M޷-o�en���W�f���Y��H1F�m�Z]e�6�g�3{�Y���;���zP�o]���xi\9�8�edE]V��˨4���\�A��M�	�Is>��À�v��o �V�١��qP�)���s�B���hJ��_�����߯��0�k�I�B%(�"D�d�`�2CH ��E1�XDbF�A�h�P�$s�%( �$h���f�hK�K��,�H��lєH���������&BGw݁0l0]�ܸ�"��Ff�# �@��\�12�Ai&H�I�'v;�cC���Fe(,��H1�S2$X"IeH$�I!�)%J��!e0�"Ē�s�dL��L�XL�I�˴�&���c) 
!@C�cC�d!�Q#J��s��1�Ld�##$�ِ�e ėw(	�i�H�јQ���C{��O<��[w@��-
��Zk �wJ�F*�sF,��]̀5	����O�TxJӷ��Ҝg�Ju�)����b��_��K�@�yJ��G�tE�X^��;�����n!i���ZӐf�֮����֡��Ù�/I�"����uǰ�G�پ���������|�{�V�"7���է*А���"qy3�C�RkԴ����D�9���:�B�u����W��8h���ft���Q��>4?}�G��D��ZjMe&2��;�9�F��%23��XY�n��՞�[��rgR*|�\eğ�>uWJ�C��UQ�~s��2/��ǐ�|\-��k;ozE8.=�࿼�̺L̍���^�8.�Y�*L5�Bv�_|x���U~ʊ1�˹��e;�z5��uƊX"�����߿Y�������i=q�L���8*Kg֏�^�tYJq�i`�*���m�=Բ�\w;�=豽�k�OM���~�G�^�`k��P�3��l�D��h�����Q�L9�S6�$Jת�n+��M��R�����6�e�~~�G������|xz-�P[�tc0[���'��S/�0�����j�b��r)f�d{*�l����_��J^��޷��x�`,j��g���xj?��C�#�N�yC���{c2M��sHB��Tg;wL>�~���c'�������P�j�{��g�V��Zh6�$g�Ū���Р6�.=�ը�[Z�b�E��%r�U51��o�5�u7�ݾ��\0m��	����ol�z�Tאb��T���y��s����+�y���g�/
q��Lz)�L,�{}7�>GH^�� ��D���U�zW��zlzts�����z���s�q<�Ë��9�I
��b4��W|�����B�g��!�S4�V�E�:�V������[=`�޵_��]ߓw���cj�F.����:�Ỷ!�w0�=~]�o=���f/a݁����2���*d�z&gÐ����z�Z�[;���z/@�����m�Q�'���၍߫���m�8-*5���bZ���I���ς�Y!����1�l�u#�'��"�����l�3˶ul���gf]Z�9�J���C��I�R�W#%1{&�B�%���~��#k孳����;!z9.C���Nˑ���5ą��3������e��ܩ�J&�8�պ/����y��zj0�&��L
�&fu��&5����Y�C�gT{4sz�*���n�M>�sKk�_ѕ�2�C��ɡ/TB�J�H�f�����?k�1-Y0��u���J^���҆7sm�0�0��\���M}tif�j��"W�j(T�9R��s+4��-��O�Qv�'�g�1��������*��hӽO�����ӆnBv�eD:kO�i*�IL�e]!�ik�/���_n�t2�"{AЏI�#�1�m��׮¾��9�4�1�Np�7*oi��ǵ�UW�V�o������X�v��Uz������iB�5����p�*�Fe)s��J���rE�����ۑl���?h�K��r9��qn#��5�����!v�U���0;p���=.}�H��A�v;ٛ�~藈K����G?��9�Oc��7R;Cg|���eV
��=+�'��!�=�@�Y���J˩�	����ӟf�ڕcw�t��C����`�8j=�^��{��u�ה��P�T���C���"���I��f����N�����5!S�\3�n%�U�P~�q>�^*n �\�Ȟ���ɏ$�*�N��ڸ{��}�^����uyQ>�_�6��*��S��*d��j>�T�. �t��Y��. �\����nB����(S1ՅTQ�9����R�}5a���U!�(D�b�Dν3<2�����Z=wNU�x��pɚ9��V����,'�DN1q戜�.�M'UN�	��K�B!�����>">�9G(�!�כ R�J
GI/��=y�l���x�p:(V��!N��*�3�{�u������eN(�.�܁k]*�@�6�>ղ�:�9�l�Qι��M1���Ac�W���˞5,R`��Y����3�E���&��.xGs/�s)U�N����Y�5���޻~�pt���yS9"�wS��;6��D�
m�!����W���
�酯ٔ��/_�)�#uU�{&����_U=*�`/C&Jg�UT�Ȯ$J���"�E<��4N\�wvPY6�+���X��v�m	F;	����!�T�u��d'Sbfr����ݝ��Ⱥ�d��!�U	�q"����$c��{�S����Gi5&�uW	S���ڧ���Ɍ�Y���{s{<�a�1��(�D��Fv_���
����T�6T�F�8�67"���k�1Ί�9YN�;|�..��pU4.Euc�ۇ�8sJ�<3cyx}�&*���/;����j�%S8�c%�w��u;>��g@��U�d��vI�(�ԉ����K4^�����Ң_��1�µ	��g�6K���s�<����ݳ�r"}�B�e����{��/�ũ.22l�K��S9� Ƴ�D�r�Ǣ��9���zn#�<3ݜף�֎�>�iX/h%��>lQ�f�Q�pUJ��������]�Y�W�U�}�"���=]K�ĉj�V\N��zm\�!�dMP4����C�7�ks���z��fVuC��6�fWJ�Z�r��'"\��A\%�zr̛X�֣�X�����d��b�Y����EKg9tw:��;tu�2�W�W�]����"�lc��r�t]½;W쬳�ݡ��6����J�HTZ����*�y^���Fr<�S^����{]�v�ݳk�f3�Ґ�S�����A���Q'���<E/�5Ny�߿'�yo�E4��Mq�B��W���ў�*����s���};YAZ�&yU��)��U��ý�>�++��N��w�3V�(fw[.������`v�]N\;6����&�������3�{��)�?u�����=����'��2������%O@x�VlC�����y��ͯJ��NV��+�C����Q/EO�����huǰ�G�پ���*�`\6�6&�зa�Oz��Y�ݱ���]EP�D�}��I���ԏ��� �#4�Rs�=��޼8߸ylw��K���Ѩ����\d�����Z>�E�Q��U�p���e&2����z19A�ٱ�U�ǆ�$5A���;"����Ѕˍq�~h���� ���4�
���^�(��3��*����r���ӵ�v����̺N�Fkvg.5��w��-]����ǂ���|$��c�}��-U�������껓���}�C;�X+D[[���;9Jj����
Y�}�:�_����}ܢ���]B����We<�w���p5t��
�P�c�ڵ��*ڼ
Q�R ��IgJ���6���.$��e��]#:��e��&'Ƣ�����N����h/�c�W�����C�.k�~59��1���B���o[��������Ƕ_-ǃf�V�Ng�L)Ϻ�\��zǢ5�c{5ߧ���#:=�j���y�ޟg����N����@�7}G�T�u�3Q�vD��z�&��[��ϙ���y�^ńvJ��z��x���(z���ь��#�U�J���\���fv�LT��s:��c�����)���;�����u�����=�eP_Ѝy��WR/�J��=Q�3� �vΊ}ٸ�?Jv��:HU�\�=O�ae=���#�/C�R V�S&4j�Ö�LrW�xv��o�K�u��ݨ��:_����Fr#ʒ7��i�my.��FMp�mT�8�9<��1����e�ҤD��F�ʽ.yY닓ھѐ��p�+%�j���� N��u���U`o&�S�Q��d�W1W#��-=�f�	���BE�[�0\�rW��{<�٥F���뼸7��1q�Sצ�zp-3&�h��+w�g1�N��#|���Ш��5s�2��h��<�@6�����~��_�$���3~�/x+��<��}�hGC�,8)�W]��e�l���خs��*ƺ]Щ�+����ЅT]���J�L�Վ��9��5����d�����HP�
�c�Z�ںl��=3�ٹ���M=��
��-6vf�g��UUR����hxe>5&�KE\H�LTj�3����=2��%�r��9@�kGd/|��r�@���?[�h�3QWW�U�\�1U�^�}.:/�g�b�q����x8Κ�{	����&fu��'Y�	?s>�E�t�v;��Ƥ��yݕK�q�|=.��7K�6a^�hA�P]�*r6�ٜ�fpL｣=�������/�W��(;^"{�����]�&��7�Np�7*oi��ǵ�UW�V�m���L��_1���v�86>�_���H�ao���5�!��h��$e�.LF*o��>��f�����W��׷_-�p�����8*���s*s�6z
[)O���S>�p�c4W���Ij��/c�+˰j^�v���T��<���z���}	����N`�tU������̻Ue��Zw}�Ү&�� �b35�X�ԧ��e�n7jU�s�O��C����H	�����UＹ����f�ʢ�T���c��'��b��e1�eK���:z

;�js�׶k�'�su�n3q���Y�Iw���\�5iŝ9�b��t�w(�1���M��'�92<�bp%Ģb&k7��ZL���"Gl���#�u�i�������N;���:M�P�fؕÑ�Ơi((�]��~��A�>{�M�w��6K�}<��DwD9o.�_~@/
��"���5��T*رS�q����#��[�m\=擾�3�f�'n�p�Ւ�b9�a�-:T�EL��kP��^j�y�,�����4W��uzu����g�=����[�;5��fD�A`<�х`k뙱��,�t��+32�����vﳶ�٧锫�<�8���')���&�_�L�*���`-1&}I���C �n[3O;���Js���˸<wE���T�H�m�N�E���AM�VCU�Bx{}�hc�<7�fk�������*)Ą���5�az8�!ʫ��ɒ��o�IdO��ȉ�����ә_,���{MXv� ��y�z�6���Ѓ���'B2/4	�ғ��߃���D�bY�τ���t���Fvemzs��^��ٌ�X�v���!�!��bʉo~�g����r�3i��1&9z�x�}�(���V��pB���T䘌6T�y�Frn�z�^{��ߺ),!���Wf��כ�;�<`���
��Ȯ�u�p�+�+�xh���e�ߩ�K��P�j�U��H�����sZ[@w��Lڳ�S
����9:�g>�ɽ�WKW��s�j�i�ŒV��SWgN�
"�fm��E������|��}�Sr��Xە�9ա���TL�,�B���I%>H��CUJQvTZr^o�������X�T深ߧm?^O�΁X3̑��Ӳ]m�3+��p)�Ef{,;�Z�<����`���j#�L;�Z���s8�uNszi�����~���+�逑�Lז-�%z��R���*M���S�Y.g<���u���i�E+.ss����KS��Z��^{��~�P^�Pk����HÔx\AU(u�Q���&k�-wg��CT�6���^��-�f�Ҏ!��ۥ@+�Q�!n���A����g�������ۢ�/��?ˢk���M8Zy�]�h{觇�����n�\*0�gu�HV6S�COm]{O���/;�{^O4���-�A�Ox���T����
�XD�*�iL��0.��AE>��U䊬�n���p2+G1��J�<nLf�c�g˨`o��4P��&���Y��.��1;��l��i�3�&�Ę��*'���\�pz�D_�ax=	S�/�����ME�=Kš�{�����U�y�/���#TΫ�3�+EO�����hu��c�ٸ�{aB���	�v����6Ǒ�W}�Ԍ;���r���D��XBԖ'��n���l3���_�p��΢ݽjyK��}��� �7 �rZS�я,owE�S8�X��Sছ�����
���V���<��7WU����!�轝Sed��Gܲ^�,�MI!�s�*����֟��z��q"Wz!�3�/��XZ	A��4�Rc1��W92|�zcs:�]�s��w��\!]3����L����["먀�z�����Ԛ�Le�B��S������#᝻��5H��6��R*�J�·9k����󪿩U�}^��3��u��ԫ��˘����9��Z>��q�0�Ux^��t�3#m�3�����p
��^!��>���ք�ã���Xjr��>q��%����+�E<�qX�G؉s]ￇ�3��[=����q2�2�#$1C\y�4��7����j<��O���aƺ,o90pq�R�z�v�y9?������?�t�܏�`x�����࿊�#���y�'�z�&��j3|׎��I7=�����M*����u�����U��ь��#>8O��e��3=_H����is�yyn �_�n
�Ǹ?R7/��u����eP*��{��p��{��o=U�����D݇T��1���<�!W	)�E>)��|����H*�3_}әY�"��	�]�t5Ėe���e,S9�gkthV�u�����&>s,����T�SF�֝r��(�/��b4�o'EE��Jj�pܮ��{�"��X�����w��Wu{K��2uq�70�g.�"u�/Ut�7���&�Tl̺��=�\��V��C6b6\IX���S}�� j�;{�x��t��+��K(�p��"�uJJf����vGl��ۙj�֎�����n��N��gM��5��^�La����辙Q�Ub��J�31�7X�U��&�xh
�kf��̴��8�3����,�����ݰ�MY�%l�2͓�\�/�3�=�g�;�51�Fu�+9LJ��pR�*}�͗ J�qS#�jA�d��l�и�!iZ��l�g����
�����]K�n��ͳN�;o�J`�C	����ݩu��%zX�;k�-��K3 9D9#��iU�|�K)N{��J�����x�cщ��mbW��\��X��T���V��8!��E՗�7�3��z�%]�^<@�VN��)]�9�{N�-��ط7(�ׄ�PN��J��)�ف_,��D�����=�JW^�H��YC��ZN2�:=u�q��7Bo#��F�b5ǐ�(��jU��ܡ�k�|r�@�:�u{�%�y�ڑR&�C�J�&�n:Їkɉ��\Ыy��{��L��*�Cd&�1��v�vۊ쮢+h��7�2��:��.�K�e���Q�A�ցǤO.u`���Q��%K�]}Kh�P�K�	Y����d���Æ�V.5���T��Y9J]E&���-�q����<[��%�pۗ6B� ]<�rv��K/9�î!����-	�g����3����1��3s������,˦�y�V�m:LԷ�o���ò���+;���|,m����]���ӹ�n�eP�R�-�+*Exá�A.]ܾ�έ&g)W;�5G�R,�Z�'yp�9!�h;do'�j����vQ�k���M	Ԅ[��D�$�iˏ|�+��@��g�+5��۝w�i�k7J�]�hС,�ui�	6-g!��^�hwjL�y�j��W[n��QN����z&������F]٩]VfS��)�8j�ļ�%])�vY�m���]��jR��v{B����)�:9���Y��Z���	���bc��(e[���M��$zoe�tCt��7 ]��>���/H����+V%��	*yr����l�����U����ev'����A�N��4\.�㛗�Ot�)�Η��wF`=k9��.�݇���҂���n�5��f`be��:VwtF������p��;��]3{sp�/)�F�C��cS�7���qZ8�s�B3�l���UĎ�S��\�E�a��һ��9xP�ګ6+�[kw��u9Q�h�����J����4LOrLZz�s�/1K̥hv������-Pcѕ�k���}��|:��+ʜ;���3]�F��p���z�.�7���q���Cgg;�C�}���R�!k��������Mf C_���1�1D��F��,��d���`�4�!�Iw]$�L�f�̉���
 ��h���d�#"1b#c$RQ����4��3"̌@���@��IH��Y0��c��,�9�,�� ��A�$��	�a��3Q�hPѢ ��
M3��&%FD�D�$%�SK�"I�9]�"��4A�$�"̒F� S% �0LH���"C`$sW4İ���,b+��(2A��4�	4dfJ(�� "��b�M�f@���2E$n�������c�XBV7��t�sqP��+8D�1��f��eH��O0��ǖ��>��e�ZwD��	��0ǹ�G��PeNS.�{����D�U��������1T���������|��v�i�&^iQ[Wv�ȬV��Τy�2b8iR.F,��U���X��g�.q�{|��p�+�B�����ZǶ�����q+p��S<�+�r$-&����Cv=W-=�fS��tٲ:�s��2�|��K���lb00"Q��U!|&%ú��� �����}��8���m[ζv��P}n�����(�y.!�;��>a�vf����I�V�X}(p!�1^�����F.�}�ǋ�����jj��3&��WP�u�9 r\��@��O��\"|�@꠺�U�f-1�⑴�������z��\��Ǿ�X)�f;	�~��L
��֦�3��τ�g����g:�3f���n_�H��ў���n2���+�dЃz��	S�q����F5����Ó�}���
lL�Y�(��D�x
���v�C��i�&�Y���*~��f���߿Y]�Ķ?(8����wE�'�N��A�К�`�~8sE�Y#/
�&0�R�F/+�f'�4~'�^�=l�,Z�SK7��7=:ً��d��5y�„��ӂ!���4��;-
��1n_G8�u��M�e����.k��T���o��D׏�z�9Z�P���eJ]��:�8��52�<̧,�(��Uҥ�*��j����g)!|������l����������W�������ɹ#�ٴ��kV�pY	���6��>��V��������e���7����N1��^��W;�c���;Cg}�'0[��B��W��N�^T_'��d��F�����{L�5ֱ7�qS�z��9�ݩW�ޑ�跆���ԩ���<��,��Ĥ���C>�T�9���WVM1���בLT�$�c��}��{Яn�-t7Q\��^W���4A�^#R:�Q���E���&�*2'�c���J�S�X�v���������1d덷�b�p��*�ʊ����R�5]<�f琿�U��V��TU�;3��3br�/^�&�m����n����B�P��n�(�_\��V0�t�p6��b��=�ؽ�~����x��t�{a"'�4D�v��>L�u�&g�tx��0��1KrW+K�ƌv�kY���ľ�4�;�~�� 4��z3�.wS����&��j�j���H5PM\̝���]�}�hN���j��ED��߽�P�م迺��zV0�`�ɄϘ2·m4d�TI;o_fx&��	�#�Й��Q\��k/kԋ�75�:PQΣAέI�[�Ľ�0!Cr�w]oIP��1��"=����woPQ��6����p���wtT9�BV�8���wX9���O��\{I�˷\Y�<�������w8N�����:{ƆU�p���8�H�Jh�l��5����1����hA�u;yU8�z����Żks}�...3�2y�����ؑFvo��T�.y�˗�MH�GK�9�Q�����=��9Tҭ���.�q�$�?X�Z���Q���Ә.X�J���R���g<�W��R����̿m��X���7.��ѝ��qw��h\���[����s4����E����-�S��CѨ�:zn:�`�u3�w��s]�w���?^O��^uCG�����"ѭ5�4}�e������xM}za_�1	��k-����F����>��z��}V����4ߠszw2�y����ȿ\U5l��5R��0)��ۀ~�u���i�R��7S�-���omQ㶷C����'AC�;_ΎN\|���<)	C�(��W>Z�U\<����3~�l�u���]��N+��d@w�!7���t��E�������|e? ;��hp���P���y�������5��W�R��- �]/���H6r�
$��q���^�w�'��.���Y���Uz�j���\�n{j����U�䢹��J"�sެ�|r5د�Nq
��g�_��{8�B^�za��a��(�q
c�:k:Ƨ87�;:�R�*R�B���Cg8g݀"s1�`�Y�g*6[5�iU�\n�ݻ�ƚ������y��Ǖ$3ш��C�.w�O-K��ek��V�)�rۛ�5E֢c��{��n�԰_�WǮ�Y�rsi1�3��0;x��.�Az]d�[>��nF]\;õn�o���(yǉ�F"^��=ʢ�ymo��w�tE����T�x�+l�C��12�J����ߺ��l��e�$��J*e��3=�T����\Hhw����ggg����눭��P�V�tj�u`5��bm+�R����X3=2��}^����!�f�<?Sf]+>�]�a�O/�ݎ�+�K���)gB2�������q�@|<(��MH�Lz�˩�x9t�������a��96���ר�%ngC�!Fr��\Ih���յTg^L�a�V��:���v��q���v��������P��d�j3.�Ǔ3#m�3�~�`���`e��S��8�ڱ^&��4q���	�PGez ��˃K �����Ѣ��k��{�D���~�fw����U��;��^�J=���ˈ]�P����PӲ����u�e�)�=0�#�e�����3�K���w���6"eDq귢n9*�A�y2��X��>#�P��q
���0���������@�Z��V��ۮ�)�EbKU4��l�/,�1"�4��ȷz��:��;+8=<X���tp7�<{^*�,M��]2֐�K�����/�w�b��R)]�}c1�~����O�Ӥn�:0<P=�������T�y�-�����_�RܤeuZ�U�����*�د��}��=�e�j���:1�.pn�|�UK����)����<�V�fS�����z�n^Ȇ�����ٞ��ʠ�k�[��10��Tsl��!5��s�eyn����U9�fg�$+!"�1��0���M��t��~*@
�u���[���lV�fW[��\p�q�5^U��{��c�9T���X�1����A�6�?(�^���d+C��Xo���S;;JFD�YQ@w:رs����Ɍm_hϗP��ٯiTؗ>��K��[:��s����4��<�=G�O�!h�?W1W9�2��=�f�q��/^D����y���D��N/@������F
b��U1-\G���!i�#ԴTK����[Т�Y��^�k����3����u��V�m��6ϟ��$ҫj���4>56��&���'zl��i�]��
r6u�MÇC>��vB� r\��L��nE�"|�E�R��Y�n�?o�/3q)��$>1*����X�ޞ��A�
�3�rʫ�S~q#n;E��z�1#Uc���[6��3��3&o&���B�-;��ɺZ��ue��sg���e��Yg���i#�0���1�6��7��nP��n�������y6�x����e�x<�sP�a47B`P߹33�Ёɓ�τ�ϱ ����se���I"���z(Q���[�&��I��X2�B�k&��P]�J�H�oo���T��������fm�3�d���x�}��u�v����7ѵ�ݙ�����@j�-fN">�ع^d❪\
��wE�?e�}��`�u��Ud��R�M��a�T֚�����]�y���9"��V���2�ю�;i�=�s;��X�6�>'�G6��(����7pf�������Ϻ�X����~/Gg3�����7����d�.q��K��F����7/�(. �p\�/�����5��⧐�R��5���F7zGL�cúf����u�ᗧ]��H'NN\0ONP�UJ����bj<�b�'I��}�ر]T�>���J�����a�KAC�[F�)^NǥiO��o��m~�+�韥@�����Luz�H��^��wqY��l���y�w\-����7�Hl'J�w�L�j8-��3��u��w�L,9�O�,MI]�o����5�3�����쥰g��N��^��s��+�C�Ң-Y�M�?J�E;#���u$+7]���z�[�2������}�<ڶ���k�ڜ�99�e3)i]����p�=������Ap�z]!�S0�I3�Ö�3;8z�{۷���\F�u]A�OM`���?N�Ɋ��_}s&�<�wk��w�lՌ�G�B>I�]59���L��05�2"q��4D�2T�uT�}�S3ʽBx������tI~|�����h�#��]d�u�&W���פ6���6�UUAO9�9C6{���3�_�_�!��@��K���VHo��"���ꧠ!�U��`����pX	�F����_�;�2��%P��%��7=r릤�b=����0c6���Ѝ��@m�i�s�J߯՛~Gcx��IN1�c��	��őq\H��"�gӓu����)�ϥ�J<�������+�n/Y�Υo�r��*s:����k�1<�k�K�|�ck�+����(�P���;=E��؛��gf����X��7.���tgo�e����
��U��n�n��ӕ/D��~�^^�޹ׄ?����X8t���x;�L���5���v�����s:`ŋ��U����s���ר�R;&�>'����j>��
'�鰕R�����&ǽ�z?m�h�백4�֑ϥ�T�Y��>{x"��u�h<�73X��k�	���I�=��E�:�9OvSWf��)���ʖ��QA;H�bRP�;�w�OLa9;�*G*'L�Ê_CW�+D��l��G9�)'{���C���-�o��A/M��~����>S��rx������`S5� �:�H�Sb����k-�s�,#�C����ߧ��-���Z����:99p���<.
�C�(���1\L� ���U�B�1߻���tk��VnӧW-�@W�"�7�xz-ҙW
�Z���ƫ�,�����<6��^��c��/gҟi�>h��������-}OK��B�n�\*0�H�W�NuTt���z�5�9����VJc�uJU���I�b(��=��}O-K����L�:G��=�a>��8�靜��S�Rlm�t��3�ͤ�h�]C�x��/�f�^�eq�k���������8�6LΙhę�QW9m\G��u�tF�X^%Ng~���̩g�K�3�Ei�o��X�W|6��m�����@m����;-ٞ�r�.*�����g��i>V�� ��7q�7�>w!N�Eq"Wy�3�`>5&+Դ����c��߮}��M�&^v�j��S��ɒ���*��Ϣ�����+j�Ƀ���G��v=7�[u�z}앻IIڮ���I�ѫ�i�<^��;R���:��:�����%�wg��8�����k۲��cu�yd4�z2����Ƀ�C��:��n�"�ц�0݆c�\�U5�ή��;����Qu�܂O�gU�4��s��>і��7��7�F��"�+s:�B��Ƹˉ-:��W!�f{��ӳF�I�W=���~��Y_�k`�q�P��xl{Q�t/�&fF�7fr���w����ئ�7։�>s��]R�x��v{ǎN\A��`���1��+�O_���=�s]�f��U�����b��v���o�~��=>_����@��i�~��`٦0g�Jf���M�,�⢵����³�]uּ�ڣ�{Y���~���Ӥn�P/~�p3^�
�#�
��:�3��=�xo3��+ϰ�'�pĺEc�|�z^�g:���c[���Z�����x1H��8Oï�_l(�<��oR��]6�O����ff�5V�W�� ����k�M�7�g����.�!w����<9FV�9إ�����~���*�ʦz�~2�*��*��*HRT�0���ϩ����t�~����JS�ȯU�jn�)�4Ԁ�%L�5�g��{�,�yE��1���I
�X�1�m\=���u��\�����_]��^��z9ʬ�a�UH]詓�J�q#TPΌ��\\�m_h��[���l`�=�!o3�	�9Cx����g�Y2o�v⤈�w�3/�_��������ĳ�qX
���*�K�.As�NmC�ꬮ�	J��Oa���(�lB\��~n������W���T�{e%C5�
Wek�]�ۢ�3��Cu���_���IqY|�؇��4Ŭ���~��&$-$z�����mǪ���㪐�]L��.�9����\�_����G"��wE��pm:4ǐ���#�����̑�Z(Tw��[�y�g�9�{���i��3��w�a9>~m�������iU�VAU���׳���zg'x����{,@��2y�d�^�:���9.C���?'�r.>f�k�E�]��a�_W��CʘʹW=�(�U�Ֆ=�5�@��`P��g���{"�����<�{�����lK�>�E�R�8w��ە[�&��I�^l¸�M1z��~3R�"e�����잹^��N���#8&LF�@��%����~�]�&ʬc}��2�ʛ�܌QZP���YYiyVyEw�8}�z���ح�wE��_��k�(�"k���!�W�l|Ud����n��c'F�wsKs��d��\rE�qZ��k�.���:���~�G�����с�`.ۊ��#��"��֩���K���*w ǅ��}Z\�Ujq\T���^��W;��xF�;CgLDc�Jb�]vx��Xۤ�����p�sq�lB��r�ĕړ]jS6���QLn<��d���.	�A�J�Rո%CZtÔz�0X�=Z.�Y�jsV�0s����i$�
��oX���:�̘�S�o���c��"�'d>6�����Ú*5��
�좹�k\b�eq�㕚{3�S���)ΰ$�j ����4n.��v��S����N�;���ͷ���S��N�n��Ǣ+o�"�)��ۘ8��;�W[K�b޻�(�c���yh���4Yٍ�6smk���]R�=��YF���]��wjbK,�P�얮Y�	��W�M�6��ۗ�{^�.@U,�ۇ{�¡�82:�D����C��ت�!07-�*�����X0i l���G��_QE��TŎ��>I/�A���]ľ ����)��6�h/�p=�Y�!
R����u����z/���%ӱiu?����̬Oj� J�ʆt�ǎ�tƎ�ٍ�Q����p+ʷɉ��%�*ܧ�v���v;�y��k1��i:���I*f�^U��mfvk��R��`����n�5����L�+�]ѝ�v�x$�nTE�<~	�.�5efhZ�i��,Yc�n���X���A�4���i��hJ��J�ށ�����%�0�i�:��knt���� ��A��m���[[}Y�Ղ8�S�mwpf5@Y�����}��<��d��Ed�ζ�Y��/��Lh�ޜ�n9N��W �6����vؙ�2����]ABƹ]PUɲ���һ�N�����3V�BL���h-���>�J��+�]ow�=�7�!�`׹BT�wV�n���T6M�R.3qe���-�g0\]����R��p���3D��xTz��|�b�ܫV�D�V���k`�3P��cд���hbt��+jj�ـ;�=I�O��f�oKts�Ӣ�:��:�ĵ+ѓs��p)�nqLg_vR�x-��Ob� �������Ý/)Nި�:	EJ�6�z�ji�fe�x^�s<�o-m_s�T��;(�9f��X�봁����)yq�·�m+��o�r3�����k�Y	UX��桮�9�@���9/�t���]i������H&��Ļ���A3j���T��ckS�{wS�̓��.^gN�]��>�E�X�Qr�)ʤ4��\����1!�n�X�إ�vg����sl��/�a��Y�9x��W@�b��aWo�ɚ�ƥ��]�)+l��|����+���g`��ðXpMFj�p[�ptCk�:�RI�����WJ�;�r�wmoh�5O/�&��h+C�9X��-6��w\za�]A)��Wrt�����0P|)l!�v;�b�ۚ�D��V�费[]���e�Yu���]:��X�S�R��(�� �v�<�t6�57�;�J�/F�[�1S!DX�8R�t>+x96ƌ���@��#c��J�qT^crl�����Ǿ?{��8]�}��﫾�~�>��-�\�Ĉ��2LS�mŅ��)(x�L�
REhؒ )�s���!�b�%��m�b�O:�)��ذ��II	�2�E&Ja2CdQ�"�wtD�h��yӻ2�E"jM"���d��Fs�+�b"n�u&:��fBA�J,Y��y�%��ut<�l�';���xܮ�i"��1\��1$@W�	�Ewt�DK��1.�uv�@�ByۤL��т5��n!a�q)�P���$�s�Ex��� ������cQa��:��L0�^-tûs��I���q]���b,�Y��t�2��]ݣ��������g��u�8��Ҡ��^���7�s�F�+���\:�f�0	Wp�4U� Q�;����1�gK]Wk���U��)�S��>�پ5���~���i��<c��u�M��qS�{�V\��v��me^�-�#�V�K{�}�����a:�O�%N{�U�WU��b����)��I���V:Z�n1U뽼�<�v�;���	����ѩ
�T}*�E2}���&�*�����qsa�L!�[�N�{=�}uE?�����j��9��w!p�*�**d�֡��T�.WO;b�0M�K4[����,�hpz�L.Ep�������0�w ��LTtJ���f��Z\
wX�=�<)��g�$)Zx�Ϊz=���_�h�˂�����4���fyT����`K�$m�l��i�:�1&"}I
�+E��%_ŝ�`,��!�jq�6��n�4�����Z-��QN�d��Y��2��\b�UymED�վɨF3�}T�=
�
��xh�=>F/��w{t;�ޫ@ˊD���D�sF{e�MI���~�R`�m	F#��]�f茺�͹�l�+s���cG�8�0c �ə��t�Ȋ�D��;8�������S�<�xr^�u�)��p	�0�)�� ���s4'�.��f�w7H��_[/F�S(RWR���rč=�,��)2�d�o�Y5�� ��g�c%n<%YO�5�n�j���p�%S�[9v@4��s�V#3���%�6�N���Kj��P/o/;��dAWC}�^���`?�c�i56��UjT�u����\a�<�b���d~�
?o�^a�f��E��)'���Þ������l��+�=��qF��ס�3��..��E�������]nP�}�͌��ɺ�]^����b0�S}T�\w33�z1���c�N�g�{�tϤ���A٩~E�� ��焄*Ӳk�X2%�0Q���Bf��<�.w��9sY���� ���J�_v�s�`��{�tk�nv�O�4���J���:�=�z�`�a�q����˰:�=9����ƶ���.b�>LQ@�`�UJq�e�n��2}K�>�{�۠(�~{�=ν���
��\Bol���T��F<��.�}j���J�����򭙷�/�ÿL��Bv_���T��a���.Դ=OK��R� �TaD�Du��;>���}���0ۍ�����c�]WJ��7'Β����s��yj_�k( �1J�w;�"�[����xiL��02r�
��0H�K�����I�и�x��6k���9��bJ�T,��E�昕���f�+q���ѻ]ΰݦ��u��
��۬��<b�R϶�2Od��B�����%aZ��o�ī[�<7�=W�T�{�J���Yl���`�D�]|6�j�]XT)	j�{�8��Nƙ�;'� ^�1�Η�ݒ���,���~,w�N�F�1Ą]�U �����~>�����׺"�,/���7�M����c]�K6��q[;�@���H\52�ǁ��!h�5�vj%���%f<�I��Ëc��ݤ�E59/�[��B����6&�g���E*.��%w�3=$>5&+Դ��+�+�3-϶�V[T-�a�3��;���B�οD!q�&��VY]D��(��ݥP7�'�?M��.��R�p˺�ᘼ\�m/Qr*ҷ3��>��q-U���ڍ�[�b�=1A[��X����T ��p4�����q�P����f]�fdm�vg��W�	��u]��t}ѽ�ly���&#��Az(i�~<rr���0\`L�f观/���}��m�nk�^/h^�w5����ۏ�>�==�(P���@��i�t3�gK�.#)L��=�taz ?#D罛����P˶���Lf�7;*1�/������p3^� �r;�dH��-��������2��$IKz�o���B��ֱs���U���諃����sQ�ݼ�Y�g۽�����z�Π�c�Nˡ�hQv�#7Ӈ�i>*�d�ɬ����;P�=u�@�X�_>Oy���}km�zU������`5x��s��_�| ��0.����߬	+H\�t��у�Y3V�	�N��{�G}.�2{F���{���:���L�~���8��}�����p^��n^ƺ��7�g�ʠ�剣X)�}�o��M�2���?!���8"���
'���s��#3Q�I
�H�LԿ��*{�z��j"^)������g��Z%L��j���� �y#���nLyRB�b�c
W�x��U�v���^�h���n9����d���5!1Jgg)H葋*.Ws�}.y_Ǯ._[��3}�~������T07�b�����n5�ʯ`@w���0}�mw�=�1����3z�k�O�)���v��O�3�T�U�턋�<ف�~�v���b��j��L����Zd�C|�!n?!��=E߅?�l��L����R:��b�p��ٛ�|�UU*ƪ�hv�e���n��N�w��X���RkԐ��FKB�=�P�atw3��9.C� rd��r<���N��s�b�
Uת�p���C�����=j+������X9�F;	����&fu��:���8�e*�|�
����s-q�	?s>�"��c�B��!��)��q���f���o2��ݩG������Q�a�l���m ���JA�@9Y������ҧ`J�|p_^�Y�Vmҡ��V���%5�إ��i��卜��|�%:�-��֌�u��q�N�j��Ԭ�k�[���d���;�c�vb�-fd1n�N�2_�������wI\�u���^U�#o���\k3�dƿ@�^"_z ��~�W`ɸ*���m9��ICj������HW9/k2��ˌ�� X�ߛ�:/���>�zE��Mu�tC�Ú�g(��P�S��7v���n�^VOK���
�#��:q�����:����{���܇F�����+	]g�	+ϫ���'E��xT��y�sq�Z���>a���uUθ�~�#|B�ԏ���]0�罷�����^��.�5�X3�K�q�����Z��W<���e�lَܯ�J���~���n�g��#�����NN9�S�5^�*�ud��b15E1S���X01,��Z���������zWdw��OAC�m�����(���^=5A�S���h\S��z���k3�]�)�aT�[F(��p���H& �2bv��X
xm]a��߼��y��ۦ��������$Wϗ��<=5�۷p�;���YB'�ã
'˞��J�UA�g}�IoVw�ˀ��5J^�}wNUudΪx<�"'�4D�2T�BdӥI�o�]`���&�dץ�Ue_���V�t�%=�n�MZ-�����v��I�& Ծ�!*�f��["��\;��R�o����N۝�
�eA�͢�p;��{�z�� jiL #��O�j��)w�[��{����8.�v��=�-�P�ګ�r��?]��8�B^�O�}I���Ҵx�����p��z3�f�7@�
�����g�w�~�;��p�42o��'�mEuW��U�Ho��=�P�f��z���t�ћ�UX�^�s>@��H�B��$J�|���u�Rb��~�Ra�/�K�jXȅ��J^ɨ�^\�f����۶�*��Ё���lL�dtW%��Q��NH�O���y��O5�ܼ��!6��>���ZMI��e�\%NgZ���I��5�%���;.̨s��Go�����.��\��~���I�j�3e�룃��P��7.���tgn9�\]�8*������x*����}�{�e�U���88sJ�<3`��J�꧂����1�9���~���g�@��b���֣�q��\t
���p�U�d��8.%00^|a_
�&n+��,�t�S�ٽ�?v�)�q��?��O\F3�>��l�܆H�8���x��B_V�`S>Z`2c|ǹ)�u������^�u��^p�Ӻ;.sr�ON5���U�y��ˆ(�f�Q�R�,��pk³p��{��	���'���8�E�]|�bV���uE�>�f���MSܽ]�m��{�3�������ʔ����F��;Jmd�"��\����㹔*�޵�*ޔ��(>5ڱ�!w����yU��-�h.B=�{�&�R�a.^�u�����[��}�5�qW���W��Ur�`W�!7���t�p�ǐ�E�M�mxQ4�b�:�*��pv�S��Թ�f�ǒ*j�ah>�.Դ=OK��R� r�"<��uJǻϫ;��tK��q�"��T����t���r|�!��@=
�N��徿�:�s��(�D4��C�_�S�h[��L�N������,#�cn�Y�rsi1���ӛ'�n�=y�W��+�yT��7�a�M1�QS�_���+LI�G��U���2����ڪ�;*�l����[���(6����q[n��3"M!mEL�q�fx�Z*O��vj�48�mz��޷ony�+�[���,Iy�%��Զ��U�m�lM��pn�@uP��jgg��R2{}���d���D��
/V�*�W��.�t,���uS����S��ɒ���Z>�E�WQ�չ���TZ�>SN�bq��^w,o�^������S}�h�Qr*�J�·9q�.&��N^�4�z���T�)U�ޠN��9��!`dd��f���S.��&fF����go҉����;�WX����k��WP��D���ͻ�������v��w0;��P�F'jh�#%�lvo���:޼��욹�)؊�����1��_Ʀ]y��g�{��5f�Z�g�17)�I|�M�w���<aΒ<��d9o��ϸ�c�W��H��������&���*L%�^�v]uz}�i`/`�
�E<7S��n�>��ۗ۝���VC��]������=>���P���L���Ӳ�g�ΗX`S<f�fU��*2Y�UG{���.�1�K�̸�^���c{Y���~����ON������p�5Z�XJ�)��`������!�៍��s5GdI��q7\V:h\���.uF5�<=j���*=�=�S����[5��6�z��e���U2���.f{L�5V�Vx�*2�1�=*1��=m�eܐd���}�Y*P����A�B��/*���35T�����Ǣ)�L.���Ǟ[����ٷr��/|�T���S;:�{ �{�,�yE����	
��������T����k���n���A�v�i�g��2tiR.F,��;�m��W��4g�!�w�-�=��Pz\k{kFD.���<���bN�.�;�M (�
��_+�x�~�C.�������K8���b��������BE����(�����S��x����#X��Tj���}��a�c�{՝	kJy��_��G]7\}<�e���t��˾�������Z�vD����'<'o7Xe���a6���z;K��|�;Z�o�k�	���x���K����*$a��n��[�]�u�PG}x��뗕ef����F�����4U�#�����1�پ�u���l���7���M*�J���R�v5��{�_��S bP@��5&�JA���������gd/|��r�93��K�u��;_�[�����D����_�U�Ֆ=��5Ǫ�ݤ����Ju��f�I�9�^���3|დ'��	1��Y]d1ޡFv��[���}�]���ߞ��^Q<?U���z�z�d��B�EeʜH�f�٬�	���P0׈���u��]�&ʬcv�GbC��z�b�~��?�U[pX���*��]W�,Vl7pt_?e�}�H���"k���!��p��V3�������s�4?�WḪ�;t����rE�qz�Ѯ����.q;�Ũ�wMn����s�s'ݛ�x�{z�@��)m��>'��e9��=.o��	�������ϧ�DLV>Z���w�3&벽�b��(ZD�⪹�W:M�vP�g�k�`,��)s��S�/��S�V{7$��W>�v�\cw�t���S�(`�9�W����ոx�_*_g���^	��P�9�_0�^ܨ�^��'�ki��CY5�����]pf�e헾��/[a�P�K�6sJ�\�5��j`w���/C=|��H�]��u�%7������\z���N��*��V�xA,�ɹ�vm�2�XWP_@p��Uw�2�wD�~���O�[�!�vT������(z�5!_ʏ�\h��O�׏M�4�VFZ�l��.�߼�y����n�3k��w�R�m�����q��CS�@;��2gkP�Y���7�3$�����9�����d��ܤ,�\�T�gB�ו�^۸~��HZ�<�6!۸؏{�k���b_ѵ칛�e<j���+O��OG�䈜b��DNS%M^-T0L��Y�ҫ�����fS�P��1>��D��묕e��2�>
���r�z�R+;C[���O~����m�"M7���W�ʩ���芯-�����=�P�)�]�bzt!F���<�4���ց�����~�L��3��ԉt.+���툗]5&+��I��P�H;��η~��(M8�&�cH�;�T�u�1�~Lτ�;�FW%��Q���NL�w:���������1�?F�Y-�>�~���l��]U��9�jLW�k�1'���^"_w��];��{(�X���L��\sN���ҧ$ᲧX���(U��n]my�3�Ι�*��W�u�':�L~{�R�(&�f�q5�In���#mN�����d���/��h����v�+o���)��$V�hk,��:[��d��t�K��.4V\�r��D�oh�#W-�uBۭ uӷ�w 2q��=ܵJ�~��p��-(j�.�{z��Q�Ӳ�� 9֮��C�9
�x9>p!0"���	�5�n�X�pF��1Dۛ��w�y��-4O-3���Gkɼ��ܻ�ֶ9��C��h%5�Q��Y�+�5��dˢ����#�i<�������eC�]9Gʕ�wj�T^�m#�DL4��C@�zlZ��N��@y��}�v\;^��Z�[�"��4�\��uwu�F����ưU��h�TbJ<�딊f։s��-����S"�͊۶��^#���"k�J�c$u�,Z�ʩ��{�Wu�0 ��4q�9ƞf�9q��r(/�
�NeJkVm����pe�bT���]kr7wb]��uN�^�٭q(9pv��s�e5}�j�tq�\�s�%+���W�v�}��[*�d�!��L����N�SYAVg?�8�_���
�c}.t�v���;WJ��Zdt�'��T6�-I�rÌ�UhֻYٝ�yg�[�uwH����U4m���q])�����%�Ԇg!�����:���ͫW�V��e��� Jnr�q�x���f�2�u�V�]R�k��VM�'X����*#IY���s)&l���	86�$�.�K��p�"2ɖ�b��}�ؾt��t�K��]�oH��]Xw1;w�5qk(el}�{�L-M�z�KC�̈́s�y.��3��#[���>�[ƨ�`vZ�O�eeC������ʉDu#������[Ϲ^N��w�y>ލ����B���Z�@�u�;��z����{����Z��������'�b�yJ�f���m���h$��U6[#��L[k2�dҽb���(2\�[q�%�^uOm���;Õ`N`��s���r��:j����K_%"/;\Ƀ�5�e�ss���s�"��v9�'-�����/�7�����c�W Eg�>�Z8j�r�Śo���,�5t�	vv��5�W9\1������|Om
ͭ�k%�o.�����I\cvJ�u|*�[n�W=}���Ƙ��,�w	����L���.ڸ�_�՞�6�]�,�}�w�qM�Tk�f؟����Y�;���a�y�6��oF�I:3���6��7$`	켅d�j��@����{`m.{נo˱NWN�ә7I:[�ݐACR��NZ�ڽ���J�6thVT[Z:�B/z�P�ҩ��w\j:��Y�I�|;J�ke���|�:�i�L�V���*�!��U�
�Q����JY�Z�9[vEYV*�����r�ʢ�E+��R�B�6�eY�j�\/��0�ToJ�F�A%~+$t������@l2�/Ź��)w �q�h��y�EQ,� �89��QSr���L�$��������wt(DRi�PQob���1	n�λW,�ۛ��sI�H��DRE;�!##(2b��y��F���$�32#b�.�p�b����ƌQ��h�.����Gttx܇��tn	��\���cEMݷ(�wv��p@m���0%# ��/0&��	�F�˜HD�v�5&��rܘN�u�ww��u�tPdMr�s	�P�>�
��W�|~Öɺ���X����#�Wda���M�Z2 ����݁Sz(����9��:�u-��nE�m]�]��%�Nź�g\�I�B��Z�H���:�^��!�2S�J��:�࿻���=�s]5�a�g١�[����z�}�΁X3Χ�['�|N�!00_�O��,��L���x�X�	���ý\�H����~���}�g�'�gF�2D��zM��6UK��S9&;f'���=>�6s��o�pp<�pD�J�s��n�=7�5�x{�U�1^�cP3g(�R��+.��Pz��������$c�Q��c������U��W�)U�}�^���7�xz�*\*1�8�5N_��9��~��>�-��8=S<�OO_����EM\,-�]�hz)��~��4���	���]����V�i�q�ağ�k��K �۪�W��ǝ$3 ��.v�uyv�x�YGݾ�ײ_O8�YA��&yU�Jd��U���)`�+�c�uҮ��I������f�ޕ\���G,ս^�[��wS��alK��b������L���$ďs���G-��n�)�t6M�H��v��4�aa���:;�ۇwl�D�B�j*e��3<bB�Rk��Ӌ(u9\aӥF��up:G��<0Vohܝ�(o��%�{���v�M�e��B'�Ȭa >�ƶ��S�)��jgm�qb}Β�z��{��-���7�j1�)s�)�pDǸFʥ-L
dW���s��(�f�/N`���sX.�e*�׎Z-I���	��϶\����<���m����|�B��$J�53Ӟ�sY([BI�X}�7۸�}ʥ�Vh$g��J��Ԟ�t�)��Rc�9	���>�A_^�w�h�M�}��eP	],n��^��_����M�vѠ~�EȫJ�·8�K:0�4�l��:�D�a�5R���^��:�N`��Xl��U��f]ngV�דӗ�ֽ�%\�2-�����#8.��p
��^!�������<rr���0^�Q�Y;/����ű^�����閰C��xc�s[����1��~�({����/��lK5����]�׏I�J	s��s.2��f�v\�q�b��z���q�?e�}��#w!с��fJ�Y_7��ܝK35zy��ղ6𹚈�;"Lk�q7\V:h\���ק�����;%��kPR������ ��x�g3.1�8O��evS����fkUk+��#r�n5֧��9�yx:ü���u3)��tא�E\g�"���Q<��S��S9�I
������U~��~̰o��g�(s��Q���o�\�SK��^�7�����<���u|
�.��͊�u��pǏ7�u��t@��w�ɖ�Нx���+�3�Y���,�d�����rɌ��6%�w�_��5.��<����."�6��Lx�Ы��gPr�Κ�aq��z����{nm�:BwJ@�*dƍW�U�g��E����\-UF�{���rQ}~�����EK�w�M\=�g� t�^��Z��L,�u�Ē���^��'K�	��/���?O��닓Z�ы�`o8�{~n�~��4Ŭ����M *|@�u���˘#��9���ݞ��8��ߪ�!]���;9��<ف�]ڸ7�ti��k.�{�]K1�K��w�b�?���*���fq���u#�,����u�:ϟ��}^; �Ub�t[�UYN#X��e��I�+ԴUČ�ǲD/z���vB�%�i�u7�^�&�F:��w����w3�eH��P�����\�1F*���Ǿ�Xюj�&���ho�g#2Gh�?n��S��A��g_�93�������p�S��xzz �rM�����P�W�/H��;�sW�S��3I�"�At/�J�H����ˍfpL�������d������I؀!�+����䁂Z��M���y�S�_�9{�T7pt\s�_�^P��=�]X��`��<��+iہ����7)j|/D�<v�C�b��+��Z�kyi���Md�<O3[;�Ղ7�cKW��ͨ�8�W�,7{�'`��ulڻ8y�����b�\�_n葈�s����;�V�Ԗ��ÝBXJ����w�����&�P�Iћ��m���9�ʬ��\�1�J��G$_���F�2���ӷ����񮾊��:�G���e�Z׻
���������
���=.o��	J|�wO��#^(u�,�B��۾��ϜC^�#S������諃YU�Q/��Q<c���Z��܁�Q�!�G������{ �[>�	ڕx��>��C����5J}@_To�UJ��X�~����$ҷ��x�@q.1����R)�E;*_J�����P��ѩ	
�Y�h��O�x��r}��r� w�N��)o
k=O�)^+��I\R�t�;����s�?};��L*�NyH1�U�ylM��{��ݔ���R�U���ny
�gэ�qqm�<=5��w7�H_�N��³���9iж"W�Q�~�}s3�xa��Z=wNUud�E�̄��b���9w�>3�\��~����=�W����_�&���*��U~5<�i�3�LUĎ���u����. Xԧ��EM�{�$ޒL��n�v�+���wS���UU-�eT�B���TK{W��#0���3�U6�����v�^Y�%�3(�ć�ڬ����nVY��@fTB�ů!Kޞ�M�K���D	!�Z+}ja�n����|D�.�]㩥�g\�J�e5�6�s�W3�]qs�f�۫�r�����ұ�R������u��M`n�t`.`��ul
��T%j��C59X�`����o�(��7��^��?z����4 ����<��N�B2ə�1�Ő:�K�S��\�7�@QV}1s�[�fo1�t�3.��v�>�}.o���z�������!pp_Ѯ0��W~D`�E��9�F��$�l����*W�N`��x�J��l��+�=���F]el7Ftm��/z���{Ϩ�z�E8�Q��zEuZ�ۇ�8s� �x0�S}T�_s3:Ƿ�-���ni�����(<�~7���p��ȻK�g@��u<+�ZvM�|N�!00^Q�)������חm�ɗ�L��Ú=̗;ٮ�=c>���Ov΍�H�8�����UK��]��37=�F[Hx�I�{�u�L���\�����i�E+.sr!����c[g���e�trrآ��'�|������]����JyF_\b����-wpx�U�U�}�{�xO�J�S=��fm�u���aw�Aǐ}E^MhaU3���S���3r|�SV��av�����}v� �4�$��ᙦ{�ۄq�2�K�4��^U����a�#��wI�[�G�!p̭�x]���u��̋��+6m-�g"�5MրT��7R�v�:41\�k��mM�Qe^�(�䷢,�3��iv��f0�땛�ɲ�tv�Lw�N��Fnq�tv߻��z�X~t�*0�Lmj��A�_Ʃ�!ﮫ�\g�t��F"�z�`~�m�&c���w�+�ul�����};YAZ�&yU�4�N�W�)`�+�c�uҫ��ˁr��fEy��?m��X<���`w��u9;6���ɦ/�$"�2�A�@����S�J��zWI>|D��f���ݽo��>��K��O@x�Vk���"M!mEL�~g�HZ*la�_v��{4���1��=D�M8��Ǫe��NNF��z!Uc�wC>w�QtU	]�7^¦����������}. {�I�R@��]c
�4�R~�f��3�%!���.2e;w�p��,]��f�YAU��^���Q��vn�R<�����M�Ѡb�"��3���-!�U9�n+�͵����F\I�|�\R����UFu�i�,����fƲpL?`�"�W���	�=����9����253S��Y�z�Ra���P��}�'.,Jbr�(�D=��ݺ���"�c�Y�.<����K��~�fv���=>��E_��L�ߧke����yW��`�ty���߷OVQ9Co�q�X�d:N�	V�y�h��m{�~U^�E�!~��Ɗ��c��Z�r�	�gMWۑ:&�u���-�
�4U���/��ب�`v�E�FT��X���oMK��e��lU���;w��FZ�v���\�nE�� ����yK����g����zǾ�E���~��w�s���#w!с�=W��,ېa�F�z��ՠe�tt_�ґׅL�Vȝx�OEqX��5^��Yν=x����,�H~7�Ѣ�}����k�1�/�G���xYU2����#3_j�b��pAQ������s�0l�]��|����hfV���[=@!p�y)�^��y�*��*���b�E;.�V7P�=�Οu�y8w��]��t��� �R���c��GA,��\y�j�w�V<:��N{��;K�F��ч����v�iYƤ+�EL��`��fA���[�����]e��;:���&15}�pCθ�l�!�Ӹi��&yw���7T=�	���4��R���.��\��ߪ�g�$��O�������wj��'F����V7}Q�-�����)����̩!陟��\����cӳ}H����vg˻T��y���۱��;�cz�8/�5�BU`4<2���TO�1�ɨF#0�����,繃x=�8}�yW0�\�����).��5��dy�sX�7���`��V�������Ժ��Q=���Kv0���\�n&0�d�c�ǹ�T�c|�,�I�b&��\��|gs=��C�j\f��EU�N!�-�Z�;3c���&ƴ��o\��H��<�jB��j2�����=���������`1�j�>�����}\���|�5A���@�|����L�f|$�>�E�WYw�j��ʭ���\����æ�:]�ڗ����,?�l�-��\S���6�ٜ�S�3��P�k�K�Y:��m�E�z[��~���}��.���6�p�r��6�\\G��UWUlV�!�����/��zE[}U#c�ϳ��]c�3>bi8�V�U��VHˌ*\�m)��G$_���F�2���ӷ����
�ޠ«����L��S��dܑ£�������|N!0:𩙯�������&늜a��y��~�{���WzC�4ϧ�Y���G(d�9��F'�
%�
'�b37Eq�<��-�c�{7��8K����=N˜�nԫ���H�/�Hr���|�*s�j��UJ����ةs�P�N��ε�	��b|�!R��a�Nʗ��	����m���TlzUiO� ���F�w_�.���\�����W�e�5�׬T���qs䑊Յӭ�ͫ����p���H_�Ҡ|��~��U˭���u?o
�j�[X�<"}Ո�-�l��Y�M��m,=�.(d�����*0�т���q���qO>T�f�6X�ܠ�κ��5ٱ��x: \�L�D�k��U�2����8�U愊���m�#�%���k��y�Þ����nnmE֊9�3��A�ˉ��2|j����O#Fy
�g����c�������5��lS^�s��n�X^%'�(�O�f�R�f��h��9UՓ:���H�������j�{�y^m(�b|�]��Ʋiא��U�5<%mD�}I���Z7�Y*೺_��!蘾��ύM�����8c���������UU9YW�*�x�+�Q��-����s����B���(7x�}����e�y����hzV0�92S>`��"]�BWl0nz��MK%_>;2}3�L�{ٛHw���u�e	K*�G�u;yU8�~@�ALτ�;�FEq"_N�Ζ'�$\ۥ�;��)zn\�u�{�s�:�sݤԟ�Q�U%Ng_����\a��A^a�u7���N���ޚP=t'5���V��R�<�S��6T޺8=��
��7.��E�\�"qO����ǹ���#6�}q|�«>���+��n�:���D�)���<��1�:UW���y�~��3����nq;>��XM�A�92���C�ވr���Y��.ưh�B���R�3���\.R]ǆd��^�B<��n�b��PBxZ�ƛ�os�r�X�$��^�b8�$���ۉi��=nPUlN0����y׍��m9�̝��u�u`q1��v���Pqv�y��\�vtO��fj:&2ws�v�;�p���ٺH���\�dk�Oc�����l��d�󞮓��#�e�m]{3��p*o)�g�Lob&�Zc����ϡ����g�C�c��_�]�ҋ-�U���u$�������\%���2�����qW��^�Ur�d{�xO	.J�0! �[���Z��1�-�w�@_.�y^����f��y"����S=/�}���P}L+��{��6�S��L\Ct�
�Q:5�JMe9�=u]*�ϘHzs����}�w?A|��ݾ�����<�/ӵ�ʁʹ�S;:������ps���Tb�f<���w��y�ݭ��������'�6��=4Ũ�(�1�V��=΢�:��t<b��k����;}��z�L�e{�e��T���ⵒf��U ����f{	�z7�N�ېW�b�kD8�\D�co�2������XZ06wpϝ��T`DA-BޙK�$�ۗ3��7MI�Wi��?��8:���U[�xOp5���Vֶ����ֶ��m����Z�k[n��ֶ��նֶ��km�m����Z�������������孶���+[mkm���������Z�u�����ڶ����-m����Z�k[o���ֶ��km�m����Z���������ֶ��1AY&SY?����Y�`P��3'� bI���B%D�J* �A!��U%T)T�)IU"UD�m�*%QJH��*BJJ*Q�D�%T�UT$R%Bf=r�mm,E�*hl���̚�6�5CT�4��M۸�5�"kZkZi�tCa��ee}���P�umiVkij�m�U��+f�m�nꐾ��2��-��Rūf6���ږ�0ز�1kZ��&���kl����)S(�6��ե�4m�ff����2ڵM�h���l��}k�6��5|   �xi^�|��<(�ӽpЪ6uN��֝Uw��A^��騡�+˞ƽuҹ�7�����Ou���9o�m�V�自3Y���,���ic|   ���R"�瓚PM��(��(���{^=QEQE�q�E�P ��{�QE=�N(���/}��GGE�Eܽ�Ǡ>�4Ak���z�����զ��ju�ڛB���V�b�O�   O�֛�F���W�l�5NW�/z�J�-�w��Qt��]�k��U�9ɺq��wv��^ܼ��N�t�gw�MR4�s����k�wb8=���kg�Ս�km2՘��4�i5UO�   �ך��n�jS������l�e3�Wt�W�vۃۥ��]����l�U�Y�-����T���{���z��E�.wmҷd���;�{,��d���y���v�����*3i�����eU+�    8�-�}w��kz��uf�)�۵���y���e�U{Ǽ^��a5�z���z׭��nw���Q��˒7U��W)w��=��wJ������f��1��׽�;;�L�]��-
�ml++�R�\��   Y�����t��]�:��Ӵ�COw]�v'L5�����m��ݞ��-�[u�ӹ���x��w^��އ�z7n�v�w;/[��/Kۮ�Ώ{�x��մ���Ǧ�Ɯv�e�%Ym%�6�ʦ��n�  >��(��wj�5V��h��Z��sU��f����^���]w=q���%$n�.;�o8U-�Oy�ڝ��]m���R�w-��ٞ�{v޺�7��;�ʮݥ]�5-�!�l��*j�bm��  ,���gm�z��7��k�Rn=ozN�vqՖ���%=��WM=�׻���v�Pܻ۸�{S�����xzUzZ�֓��=��y�������׽Gz^�64��u���^��Su�+Y�X�O� ������v�={����uj]�s@�ݻjk<x���s�WN�+���ݞ�Meg��Ou�֕ޫòz�:��u;�^���W�^�C^�7{�TJ���oyҹ������� �{�PSŇA��6s�׭���t$u��<���u�oW��n�^�ހUʫ�ـuowzmz�vcy+z�(;��RT��d ��a%)P  "l!�R�  )� �*   "y�*Hz� iI���@A�����?���������T_gg��3+�����w����ַ�~`IO9��H@�y!���H@�B���$ I�HHd����w'�X�ϸ�uWaݕB����b���J;n�u��uQx���#��3�i�4-��V��J\Ô�sv�9Y[��&:j[v��26Ɔټɒ�	�(��[b�&X�3-Tk\۠y�Y�*-h�����N+��^��^��o m���J�k	��QH`��n�B��yL�4�PhP��j�;����)ӊ�ɬ�)4�J��K�1�жfM��n��[�O zY	,-ɑ�V�b�=�D�L���z#���
�+euGi�l�WI<=H�걒)�!�+D�ʲ,V��t��B+�p�9(:�7��eEI��oM+���`�j�l�����	~�r�3�����ۚ���؆�B��ؠ"�TѴ��݉A@	t���m2rf�(Cr�6�j��,�c#x�^�e]И�����e�Bl�7+J,���]^2m�A3���f�
��l�R܋K�5�e��:���K)[1d�iY�򞌔/*l2�@�yP-���U����h���yjʫ�/Ya�4\՛�-k.o�^=
�7L��N6��Y�L�fDN�n�*��h%�#���qˑҫV��X^��G�Z��z��3�{N<"�gЖ&`wz�qcīm��
ћD�h<�.�<�3q�x�i�T�H�E�F�bݓ{E�T&Jb���f��U��x�ϣh�R�H�ѡJ��s/�ƛT`&����.�A#�՗�]�2��=*�"%�d[�fS�o&��U�c6C�`ĀE=�YW,
�X\���n�W"�w*�I�qMԕ
��5M5��:i�z�T�̦��� �U&��.�4j�n�6��ʹ������C�b�,L]�7�A�Waީ���i�%�0��披�`	*�Q*��n,�*9�M]mG������DVV%b��kOC���M����Q�eGR�k�f�2ťu��ۻnSY`j�r��Jf,���cqUַ��[L��J�p�t؛����yV�v@h��k�]�WN'�:CG�ْ�
d�R��s �3
�+s�h�#Ӥ7��	r]�m��'Ζ��岪RP'�Q9�[�ۢ���It�a:�@�/)$ɹY2����e$�{cͥ����@^'�:j�z%Đ���	��:�-����:\1U�Z�ۣrj9�-h0�Ia�bm��f�[��=Wˊ��	�Пjkúi���qՃ��wX,�vc>*ƶe2���S�v�z�GA�%�([�dt��F��	w�� `Y���C+A�)��i�i�X����e���+%HJT�*�Z�F�-v�Iڰ�o!ăyn��q����m^gon�0�-n���Q��h�r]w/7VFMl�C70(�]-t�P�u�S"u�P�/4Q�CX�rᤥe�3Zj�6��O2���ҵr��q�d��'��Pw
�ӏj��8�B䫌d4��X�/妴�k)��?+���Գ��%K\t�T�����rm�0�+;w�kP�}���H��/0����1+6&�v�9w0;���w��Xe���HP׵�Yp�R�`�*�6�0���^�Ą�6�Vљ��쫛g�̩yt��չM�ԯZm��C!&�dK~�4���Y"�4b��s�iK�F*KD��H��-��I��).�m�v��
(�^��PU
�A�C�ލV���]X	��+4̽
N�"N���g ���kuԚ
�)�kVG3&Y��,�`Q�ڻBAF2�A����V՝�[ֻ9���x�Z�`�L*Z�^9Pk2�uGI{Ei�p��`��X7��qf#S��ԦK,*�Plҥ�M71M��V�Z�֓p,�ͼ�t��W��ɸ$KM!鳸�Y�%3�!�Em=C 4k!B�0�*;�BT��������Q�M�K]�Ϣwn�̼֎CXb[��YM`RknK	����i&<�Vsi좨��we($���s$�򂩹����,�YƩZ�[�6*e]X@���8�r;37l��/(�cj,�֐G��:���Ҭ1e��J3~�s�4\�N�f�>���=�m�ksj����4H�iV���^q��fJ�J���/�z�[@![{��FHr�,�!4U��?JwB�3�V��`���5�2�)rU���k%�B �4'��Z�:t�����)jr�x	u���� 8wV
��:{P�cP_&��֕�+i-��V��DQo��V#0��n�BSWMf٠#{Ij���n��AjM�^m+$@WM�H�{)��X�l�.�A�{ I�(�'�Y�y�����'�敘�vTv,���jɎ��^;���)�8Q�j6�(�*)�6e��S�u�6����!�a�QJuh�����*JB�m�����B�el�!�&V��a,���Sp�F�T����:�6m�IѢ���f�zH�ȍ�ݨĩ0��ab�tN[FF��S �P�Y�j�t���l;ٲ馜��m��*"�v�33-[d[F�
�5(晟+�7����S!z��7���;v��*����f�A����׮�^��-˷�R�I����Rj�i����f����+�t�F���ϣ,V]��d����VZP��p��!��(��P�DՈ���
f��TSޜ��h*˹��tA�b˪`B�ed���-w���/��,��p�bf�A��q׊�j ѬT�]��%>��a�.�3
�ٺ0��m����OpT��L�;���en�_8�ĴRzu�B�&�������݊ke��*��!�d�u3z4��P"̴2,��d�x��0�t^V� "��y�m�$�9����B���SL����#v:5)]KUq�q��n�0����ZڌL�=`��m�̻UвD��퇘MđJ����2���opkͶ�@^��&��XR;�f�v6��~�D
l��
'(n�В-VH4�R��ѫ9�Yq=��CD��zmT��Zw4G�	r�Ze��*��cu���&ՙvE��0A���
i��@IQ۱�5i=�-	��a����Īd�v��&��`ˤ�%Ք�+8.�)��iuE��:�N�^��-C+���%e$5�1�;b�ѕe`�**m9ʔ+׺t���T�e��̵z��R����7P�.<b�V�ŕ20mm�ӈ�oB���v3��v��u���SoY4+]1M<���Z�5�;����j��Ŕ޼�U�j�M�X�[Zm���M�����-՗�f���-ubnID��wn��L��e���F�Cj�Q@��AX��N^�%c ��͡�;+�و��!n�`ȭˬ�Y�c��=��.]˨�n�ؐ
��":�*dؕHȀ�Ɍa��1������w�jPzM�ڌ5[���y�`ooSl�.��B�˼u��P¨Є�*Է]ã/��e>�F�d6�u���:��êe��C�!bȾĬ�|�,�"�2�s[{NnӭY� kZjiēb����)<��"*Y�V Q˺`n�T��V�GiԈ���z�[SIC#T�F���*���:�c[k0jW����餒�Tm���m;q�{#.|6��
ʍ}���-׬�V�)�tk1R��t���jK����R#��V�����L��]ળ���Jɺ��(�������l��7����v@���5P��p�p�k8�����M�X�N�=���m*�U���� 7-�
��eaL�E��@2�o.�ښ��h��{��ݳ�]m0G�Fn�X�L�pP�t�S�RNL84�N���:��3�(��+�ٸ��O�+$�/Vj�5K�W�p�Ĉv��GQ����I�]J2��VH�J�'�c݈�jPj�U޹Jn��70��ʵ6�[2i�K�"J�	��{�np�8�=�u9	���+a4�6����͍U.P�1Q[6�J�r�e���2�q�JgQh�)h��L{J��w�v Z�=�&�r�DՉ�M U�:��E��v^^e�fDk4{O�i��\#TzBr�AS[B͕Y�F��L�i��#���F�
�!�f��D�)�$��O����&4v���3E*,���,:"V�6A��
�@�#��DV�(�n�Z��TM�܁L*��AԬ�F�b�˻e�j�k�N��-���V�lɉҭ&=Ii�wD�%շ�+%�RR1)���+, Ò"���YE==�63%0�u�6�:4K��ь��r�
��^�[5nސc�7qћ��� pIB�����e�F���*FJ�WW����kq 6�6B��n����pƝ��#!���;jlG/&2���Y�9Kg�퍧�+��͙0*I�M���2�D�l+x(��U.=b����v��K@�:4@;��*Y�U��F<-�.�a6�R��+qcv՜�x�J��+$R�5�I:�NnK�haTo�i��x�#B4�ɨ�����9u�3F�X�5�b��Xr��>���&�X���jҗ𨦱�-��Vf�饳kf�Dn�� &kl�;Zv�ޅ��&I78��:+oa����6������ss.�0m��r�J��]ؔ��p��SԱhHe�pX�����u*knX[mH�,,�ͳj���ZڣXMfK��Ҩ�D�e�8�T�i�vP�����^d��Lܭe+�q^�\��y6�[�b:�)�H]8]`�A͚wj=�e]eA�N��c$�T�3c�l��ӳ[�%�F�7>��A����ф���ɕu��4�<Ie=H�J���m`��Dt�h�IM�X�R�wKb��mU�HF��U�$c�mq�N�U��RwR^��.�ڸ�Ǘ���l� �	�m�B\m�$��VǇs2a�n8����� ��=9��(+l�F!����utunhi|MYH�MklRL̔�[����\��J��$�c��""	W��b�+֡��ܱ)�t��w��{)���`:i���E�ЉZ�2'��KO
�A��[��-��f5��0v��4��ֵ�KA�v���!�[��tQ�DaT�off���,�b}Bd�&Û[�݇�KIUԦ	":v.:9���;!��iճ5��Y�Ҟ��5�� V��`��ƈ���E	�ҞآX��O-���4�5�2�af�)��F��"�m�	�.���R!��Qj�R�÷u�^hW����.�dw�L�e��SɥT��tۥ��ʻ'�.�Ҭhh��^G�4��0T����塍�SW�lj�:�G��h7a���u�&$$���T��`�7�}���ڒ�� �0n��]J�yy��ю���/�u)� �[�q�P��tL"w��b�Ce���_]l�oN��q�����\�&��S�t1@�C*V������;�c2�ʹkI' [V�yI��m"���*�� ��孒C��n���eG��,��JĳxM1�c�]��`���d��%�#R�Y�MM�d�0^�\?�f��t��4(�i�&�XʺgQ5�a�fQCgsBj��-���j���r�!m�Z�c�SH��[1�p�ئVdYw�B�m<����ۛu��,|́�%��ZI�-Q�ٶ�pJX�8pi����Z�Ū�������U�3c�Y�Z��l�r�s�A*�I"���7���r�\љ�m�q!9q�m-�����h��KT�n�%A�I����vl�dF�a�Z�J���F鬎ZT2�.jjb X�)Ŕ��¶���3m1j�DP˖3BN,�a��2�{�9SP�U��qV}x�1��x�v�9O�4��b,�P��NN J!�ťYG��m^D�*b�+��)(�fܺ�F�&������q�Z-kj�4��C(S��1W4]P%ve�Z��k��@֋z�����7I��"	u��R���C嬊�l7�ȋ�lU�MN�`�njĄ,Dю�VkRe��K� �7^b�[)��)e7�Z6(�٠�o��3	h䥊�j�4#�
�F�@�-ʈ�x"%[[!����ƕfݾג26��^�'T�+rm�E:�����ut��آhLP��W��a1�i*z3Xih�VAe�����4�a���3��J��L�a�2бi�F�
��-:��<7�,�T��-G�Z�=.�,Z*�E�[x��R��YG��[��j�iag5�x�T�9f�K6S&��(D��ha.�Ff�D -�"��7
�
�����gt72n��ר�2�؂
W��ki#���b�e��H�.�a��5���v���R�k��`wsM5��fH5fl�1�j�,ȃ����F%n��gF�`�Q�T�H�K�Bfi�t:��e��/p-�x^hd��O���Z k7HQ�-֊����ӧ-U�B۔C��<�ӳ��Y��U۫�5���!�v}���`����++ڳ��v+IZp�,`���p:�6���d���ѤIb]2���`Q�OW0R�N�q�4�a�	w�L��  !��f�9BB�$�J��tqڠ.�M `m��@�ʻ5z4|ޛhcZX��KGqIj��T�Yk?)�V��X��F�/N��6�sn�ǬtĴ��������cv}���[p;LQ�w/bxI����ٍe
p�%�͔�[�I�E!�n)�Y��9nZג��V�1Re�63spA�,�.]ejj�[�i�x���N���1�⻳@�چmh	P�O`���i��44��ûFh27t��M�!#W.G����v;�VB�4M��3u�kJ��aőn�t����p�:�Y�{��d s�F���0[WQN���t�au{�`v�gE�,�;�]r`Kı�}��:����N��c�T;�5}�^̢�)c��خ.���n�8';/qa��<!���>ЪI�^C��m����:��:��Zw�r��7��3�*ʐ�����<vu  �y�v�lxWv�'VJ�H�4U���X�]O{a�!�r��4��6�/"-��tE��
"�78�YL�&p�'B�����i��=����or�p.xSY��y3j9�B��)-6��Ϸ�Y
�����̶�:��<�(��k��T�-{�#:��^sybv�]�]m�4b9�ɪ��N,wejlVK����0wS�0�u�e��-Zz2Uu�t�\Q�:�ѓt�>��=��=��ҩ�[n9n�U�Äب:�u�|��a��"��7
�����ks]ቋo2ۧ�c�����_v���MAm�ftA���%�1q�w5���k���Xڬ�u�`భV5�q�J���smS̛VL��ꆸ����-S�+yKUSu7���խ�z���j����p�fٳ�t4Hc�&��aM`���sI��i7O��&��sc��w������Z\+.m7�DҊHᩀ�����2,��l�����}��g��dc '(�W]��3oe��O()���T.E��h[wׇ��J�*��G��*����#㐌<��v{9ꇍ��w�Gn�t��+��XjfN/2�}����"�+�F�*Ji{�� �+2E7#	ֽ�0V�R�������� �8qp�ٷ��!�R��.!f�R�l��g�7s��疫^��Y�{Z9�#���M!�\��o���uӫ g������G0U�,V!K_R�D�TN�z��bC�.�G���zu��= Q��Kc���C�7�iI�7���mWm�(N��o˓l=^�����[����$�%;#9�S�YJ��.��0�y��9��eR�̎S}�.��j�Ww�(R��{HT�h�YR�2U���ZVv>�����\�4ރS�Gb�fzΦoD�"P�]��_t"���nQ뼦w9gt9�=ݡ��ӊ�/%�&Q�X�rI��|����Нa���&��E<tP�.���e�m�����H��Β�|iw��l�z��s���"uve�3}��ݖ�
F�@��fdU��M`��m�HR�Gx� ��#�c'j��u�&���
]y� �zi4*��9P��֢�e.�K�s�P��vi�͇c�����xb�/]��ֺ@�^��:���Xn������O+t�Ӵr��OGMx��9�bS�Ŏ�.c����|2����#J��
I+��Y#��o�f�͙��oP�5�!n�2���*���7�+rg
[y�u�c[�Wt�)�T9t�9]7��ʺ�/���Y�p�f��SA�N�U�t��C�6�(�����1�=���Ь���h�P�{n����l�@��
�e]YE��\qm��N��S��(]���[��4�mi�B���Vԫ�[3�����Z�OE1Ԧ�[D&��@���w�l�Y2�^����8�y2_*���4[��qn��dViV	뇻9�
�����t��Ȧe�S�3s�����Wd���oVl@J���Nͧ��(V� �����bmFB �z���E�K����+6�91k�ko#�8�����*d-�zRܺwN�*�%Jó��ٍm�[�i�'^]L�w��.Z�vF��U+�g��>�=�>.���d�\�uw�R���F�V�]]X�}ռ/�_1���v�<��l�%�˄�:�������;�L:��s�)nJ$��j�nW4P�i�r�� +z�u���[pf�z{#�;�!0�f��9�SZ:R[kr��Q�X[��gaP���d�N`�̥�
¨��yl(8Z�y��[jU�]�x%�.F�E���7p��a]-����Ds�Vt�L�Ͱ�J�����]�4\(�;4V�^�u@-�w�Ct�E�l�t����b?�[&gY|.�j����yR\��{R�%1�Osَ�<���Ms�8������p�n�x%�ے����N��8Eu�n��I�uq���LB�嵪T7�J�Hd{�1�&�;u���Vʘs	;�]f��V�<e�$Vu`Rثt��x�O��F��hKj]�B�13m�m[�x:�,�I	u%��������&�u��i :�9i]�@wtv�Y������1�*M<)��mov+p�K�ҭr0G^���={�h(^�ĸ�2�6�4��5���2	I:I_Vc�C݄���}�Ȗ�#O������]
�U;|�`��n�TPF���ʁ�R�ur�u�l���tiͶ�;�Ҳ�@�M�575Q[0�r�\�՛yX�Nѣ�
�c��.����8���]����5���h,h�Wu<q�����Q�c�f�R���mXߊ��r�@)��4��؍(��������t�����W*k�ۃ����)��.���|���q��S��H�Q�+�QcPx{�T���Z�`�ˀ�c�l���}�:���)�8z����k(NJ��a7�����SVlӼ��R�
�ywo+d�c��Zi&|Tp\c���{��}vт�1=�89e�+s�\Ӂ��%������Kv6�6]��j>ō��Y��H��Vn�!�L�������N�4�˰Q��v��cR�������m�\s,S���:�S-�2��ݭ��E����7��tK-�_`�
N��d2n+�3�,�M1�Wjx(ˊ��w^���q3d�e�	)��&lq��0+��M�3Y�����>PV�����.����ے(�Z:��4P���wK���J���N��s���Ǚ�(�\�����B�X:ѹu���cMM����Y��,��TOl�K�a���Y��W!la�c���B�X�o��#ےƌN�4��ɗ���)fl}�L��J�{N�a��	a�sV7��ˋ�w��;�ٜq�@��C�h��}�t��.�]��p�%���0^��ʟ:+'�wbU����%r�2����x���ֵ%[Ys�ת��7�Y/�;�|�[�qo.!�
$�|ΕWBs�/�p�ֹ"ctd���}��deҗkRH��W0��Z�
Ŷ"�kZ�/�MN�J=��Sv^^��:�<rĻO�Tں�
����9CL{�Y2�[CW�(�X:,hGa��eCi<db�$B��]9��h��1ou$�A���(�8��eI�@���bY=S���K��
��s2�1NWk��Pc֖,U#M�M�R���ŝ���fx�+���j�M��K��%u�B!
���mݹK��r!M�7�Ы�zʠY����.Sp� A
�PG�h��*��W� �o;6�h�!�J(�(�M:���\U�ø����E�H���g���]��g��u]n��jkb	Л�7*�X�:Fh0|ի��V��)n���g�eo(�P�6ve�.*utL7��������ىXƝ�������ؼ�6t�-m6�E�tb�z�EGZ�p��9�b&����0�F��rIv���e$7Ҭ�J�bk�:�]���Uׄ]\�6�;FiCSa0ޮT��i�C
��ff�7A��m�h�/���O�Z�Tͺ�I��J�)�̞ܮbf3r��J�j�³7�n��/����Ԗ��G7�P�� �����EC������^L��۳X�m͋�@\6��ܒy��̮�&�lk���Jͬ�[��+��j� P�_Lsf]��\��� !޸�S����w�DzR׃���\�S&��;Ή�J{g��&��:�o[1��V���hfH,�]1��,2Yv+u��mc��u��֢�fd��,3�9{�L}�l_f]�HJN̤��U����{
���������x�[)���ɤQr��,n�WKO�GY�db�}ؗ�U�9��q�^��(�O�d���=V:xѸS�0g.{�����º���n�J��W��s)k4]��+gΦ��^��:��^�����kL��$�m�M^�aV��7����r[���f��աR�+^�rq�Q�i.�L%Q�}��1p����H�[Հ��k;qB��J-��75���Zp+aU���;���Q+�Tɾ=t�Y���m
6�h[l_WM�ډp .e�@Gх˳�7�=��ř5�"�����7�JZD���7��	��s�wf֯��� �ǷS6�P[�q<�t��P��T4Ә) ��KK	]^Q��v�=C��֦���]�b�s�f��.��U���%#�#��#}���a�5	d�o*���ZŲ��(T�+��֢c'T3t�T���A5="k�S��6���_���=�Y37��,a���/�rj�I����ѳ�ڰ���ֺ�)1��m���(]�7J��O����"U|r(f�P�H�/��`9A�$E\⃁X�����]�K��5�Ә����4o�M�r�V/���n��\ue�.����+�ªVc4��V�d�.Ռ���S��	D1G�'UAJ�u��L�[�C�.2sr��ۄ#:,�VJ0K�+7��[���\R����l,����F"��J�p3�(o�	8I/3#ɣ�^����^J��݂�Eǳ��JhqW@� f;�鋩�JҲ.��w��v���/'uL�!�}�e�=hQ�m�^gT�9�)�6Wp���2F�8V�h�:*-���i�扸���E�j�N����T��>�ɲ4Ep
�V<�������ٯ��2��S1s��U��frre]5�1����M��j�����NW#,���zh˵�&c���6�Y�X�L�}u���M8�e�$�yK�wh幂�C�x�e�73�{uSDD�jmVU'W�]agK����^4�_=���Yp�k�WOs; y�q�f�ڽ��+�Alu�	��v�>��!�el��7Uګ��6�!��&f���!u�P�6���"㽪hbu��|����Q��c���^$��<QO5��z��I�0�	�tDu�0��V�F�+63���GPIya*�O��w�s1�����}R�<!&:���)k����n�m�"�v��`��F-��t���%�T"ǜm �����Kn�\�`gi�ml���s�y.�\ ��{Q�S:� ㊟c���P9�iat�mV�ĸ�ٕf������i�uN�!���}�ep��̙jਁI`7$В��`Jݱ�;�u0J�\'`��9�W� XO-�a++6�b6P��g��>�������I�d����Dl�t��sr�f^�T����:k�3�{�m�
2���p���hwu5�q��7&�Ď�:r��i��y8c�囙�V9:��p\�n�v�J����dܮ��F���(�й�Bf�9ՠ����&\� �5�a�X%��,����n��[��z��^
s�A�������mU�}Qn^i��ƙ�BM�6�A�׈\Y�v�ܬׂrv��zk��ɧ��C����fؙy��-��٢`������P�׼��Ѷ�:�a�cx�̷�� �β�[�nr���&��l̾��5����%ǽ��М�R�L$��,�z�n��HYj�F��:Ox"@�JF���t�&����2q�B����X�z�{%p�S���(U���j�o��㧽��j���x�-+�H	��M1��u�h��`P����p#�
��b���e��33f-��N�ކn�@�W]�Z�|Ѻ�#�;1�0�L_�qS$���3:����5�`���]1�r�.�m�<�r��"6���b��')l��v�-�x1� vi����}2λ�i����L殦�x���\�l����s|�mt�.?B��ܱ�(�E+gb�d�m��޴���u X���*�c���۠*��}cX!��cI�9�!���j�WY�Z�f�����P[�d�)�����Vt�K׈Y�tQ��ε2��M@u!Yd��wboe*��������]|�]J�q2�q�rv�{�`� r����mW���=+A�5�,�3�v��+�̮��F-o�pi׫��г���ɍ�����!O%�w�M=�y���[����d��Ř��M�
�����x%֔ʸ΃��NX�P�W�!�4�!�������JԹ^�?H�]��D�t��%��*�7�G��}<���b��RbU��&�4,[�H� �F�+«��ï��@ӛdej�����)�;�Hk�Y���a��
ۓ���Er�@�;6�s��b�y���M���+39����Ki[���.P@�#9�e�f�9�ރ�ت�9�f��\MH���)���@��h�&���S�Dy�靯$���FN�SJ���5�����W�7	�mVܵ�� 0�ǖ7Ҟa�Yt�M	`.g�t9�$z�e�����Դ��=f�h��k���biX9=,�vkp.z��me�h�
[ԇK��5�<���w����<���Ռ�P�yw��ȡO�J-6��B�N,��盕s�w�Nm��ĺ��+�x�����hd�Yс[ӌ�R�Ҳ��uܮ��,v��*u��[ؕo3+��^ˁ>�ש�tM�YJձQf�ɵc���J�#E�8K����d�u�1��yO�uN���PN9��.���%E}v�T�'t�1�ӥl�'z�eIus"n����������wg$Y����!�����$ֳ��{sؽ��~\��Z˖����#���8���ƅ�1
z.;��R��3jv=��-�X������sX�8m�����LSӒ�S���Dor��ҕf��R�r"���YX��Yb�b��A��*wES���(Z&�,���rnC}�よ��vk�L��J��]��Ԩ'v��GX<t\Q�Ոf�=�l )�
�D��!v(U�&kwC2����f��-7\�`�Z�*�r�]l#����Ge��d"*��t_]'��G��A`ћB�3zA�G�!��$}JiqK�+�\t��A��䃕92�.*���e�.�\�L���j�mu�.r���/,&kƹ�L��
{^Ѐb��,5}�j�X���"�4/3��Xw.j��F�5���P�ǵ�m�,�K�s.��p�$�	q�]s�HDm�VM�9hP�m��Ӎ�j�˫��:knV�_]��'��ʸYN�B�Bmf�/��me�f����}��Q���z��љ���xu����)]��Ho0\ 2���ð()U�1{��,
۶�'��Y�z,�ň�o=[WPw���M%���i'KS&��������V]��J�;N]��}�ҢkY);hN=K�ĵ,n���ݺ"H1�L�i �Da���f-�X���.����1&���]��g�vC�,��OBCP� �k�/�}S��YJ�v�W�d�#K)����h�^�|(kGC��_ �������Q7V�m���A����u�e�K&�rӝ,M�sr�a����(R�/u�-���G.7�:8C�+�J�:�pi�jչ��� ��,�vehU�l�e')"(��b�����.競LA4��
�jjh�����K�|���I�;&C.Q�����),ҟ0��(���t�w0&���������w6tn�X����wɊ�@�����,(N]`p}- [9�5������ӗ��gT/Y�L5a�l1�Mm���#v��x�-�9M�Ĳ���=\�6Lb�[�0��m��A4E�ú��F:���Y԰���\��H|���7�[θ�^��yIݼHى�nGIv$,��iО]1:�ͩ�"a��4VG݊���g[�8l�:��x5�G�tyu�4Њq������/�78YVWƃʗ]i�p��C8gQ�-���k���o~�9�Ui4I�`j��>+�a�;KZ��<QL��]e����Foݫ�G�9q�h9�^�R��0c)IX�Z��7i�[n�E:��路8�\��W*F��C^50�1AlEt��n%�F�p�\��"�<�19�fϏGf��b]��lg��o.�<؜y
�t�B�,m��ޟ�u���F7v�f���I�|�Jr�Źr],�$�V��]+9-���5��R�EC\7}�Z�'�փ�{�,��d��Y�nIӝ>>�[�*�VIr#�iX������Q92`7�@�{7^X)�H�a|�OFo`��/�#P<��j[\Mu�i��i�:b�!���3.��Ǯ8:�_=�-#�K!��^�v���E�ޮ隇3Թp��]��g0�τM�xӬ��B��T�;N���6P��d���7u!�t�[}�w\��v^�pn'�m;sg*O�lNu^n��1m�{w+����m�t]�Y�/���2"nJy��7�j��Rշ5[�z��CY9K}Y+~dcXLr��n�Y����bZ�E`K��Eʺ"-�E�,�r�!��#���9r�Y��x
'�mv��A��ɣ+�x��D����t�$���ԫ���U�7��툞Z[�\�܆Bv����4H/Lmk5��,�ʧےBK<��Hc�2�C���ԉ�@�5��Ayb�n��1qפv��]�x2��µ7�-���cɓS�Ur�-�o1�`��R4V�u����`�*^�)>5x{��zOU�%��z墤�X��h$.�k��w��X+q��:(�T��N]�{F$�]v]��;o��]�c@�|��cV*�D.l�b�)��n�ټ�e֥6'],K{+�.R�FR��1$0���Ɛ���N�3,����M5�Q��4��X���ȂזJ�QSh<gN� �0��U�Tҥ��\9SY�wXÑ��������+��"5���wn@��@�anh�t�;,�@�f�7�����4�p#=ē[�1� �)�q���vAI�s{�j�3ص3�'���h`PvF{:��u��9���c(q���}��tP�i_R{6To����hR�1<�k�������;��
k��j2��Z���=WDW:�s̡W��7�[�@���s)4I莮�*���Dt�ZM	��X��Ti�^�v�Тՙ��;��+��v
b�""���y�F�L�],!�sP�A�'Ǥ�QP��Wl�����j��{�Ah��K�N�˙"�Y	�̼t��tm�/(5�(�0C{[�F��w����ܔ�uIL�L��,�R�S�A,.�Sm��gj�i�-�.7}'wV���U����Se�z9]��j�r��FG��ED�Te��mR�c]{�N��ԧ^G���%��;�ŋ���gs]�v*YE�����D���n�.#�Ϯ%�W	6��xtm�'�w��������(��M���>v���l�<7���\u�f^�(e4{Z�y�3��D���v-�/���q#���_`h�S�5	|SS<N!���!o�9�bB�b:d[�Q�%"�&v�1ku�,��^�GE�� ևAZ�fQ�ëyt6� �ǽؓ�غ�}u��QGD�޼
f*z�/s�54��`8�ͧg�]�3�����.=گT2�,:��Y:�q��ڍ`Vz��S�R�]�3��EЪ�1�9���-ۭ���y��0`䳷�j��*��b��W)��c��P,݁�Vbz��U�jvڥ�����S�[��ev;K(�œ�|����dKU��Q��X*��j�&w=�Yj�`��:䀕L�+� �{��ۮ�-�Ύ��:^�R2�U���ܢ�;X�;��]��+�Q��ٴMY��u�'���]J�bT�DM[a�X*u��C���!�Tnh��S�^D�G�̢�^L]X�!�����9L�ޒ�ۖ�EdBe��o�{t��L�օo�����T_ "����6#����Y�DI�����$�7v=)�Ҟ��.@�!JN�����ڳ��F�A������i�[I��@�XW��2f�K;��J�Pu�a�����;�t�� �K��kXڒ�a34V豌��3A�cۺ�$ā}9��Uz��S�Pm�4r����l̮�qԊ���ouZ5���cB�X��1;�^ɢ��ln-��q�F2�۳����uڂ��N�����H��#1`#F΄EyF>�ɪ K0��
׎h���Dq(JZ��әHr��
����Z;*W1�SKLܝ	x��Բ7ذF��Y=wV�GLǜ�(vQ�,���9
��-�g]�ù0lV�E�+�����`��.�u[��#"��ޝ7F^���Lsՙ�m�O�|���-<#��L�U+��ugkrPf)��+w�ܳKxg#bQ�w�`�x��L&Ҍސ4��.N�*تG!;����-��q��@Q���t�؋Dn:.��r쾫Zq6�H��_	���fq��`�ë#���u�9�5T���TdXW\b���{9U�ڲ�Y$v��1Q�j�c�j験K��Q=����B���Uҥ�&�eT�*T�֦�[�� �oL��]v֡vK��W-]!XU�R�	lQ͕m�j+���v&E�۪��nAu�7���H��M�F��0^�����o�=e��eE��9���xkuwR��a̴soh���S2��8��!���^�\�|�9?������6F�ou�uh�ʘ����!��]oQ��)�Ev�d�F=��y�����PX(�wU�-���w)鱮���k��f��b����F,\oF�L�g0��-KN9S�.��)+�Њ�rb�S�2����Wb��)<��n��p5����U�)��-ZxTW
U��v򲊳u���.K�tK�9m�+�n���F��N��k�AMXX,��0��I�ɀ���e(���E+�*�0�����,�v2%Ag��x\�f�EE�ֵ�U�{�����p�%���J�}��
���1�o'.�R�����7�o�c�J���J�[�0�}t��u,��$T����4�9��#�w,�U��H*�λ�p󂘻���4��E�ڵ��o��(�k�`��N�ݙ���1π���:X�<�L����Į��~�3�ky� z�9�T��*��n��(J��nT3E$�R[@Q2�ov	JjU*ط\eG�MC��[��mF.�#@�טE-��ZB]��]�y,H��[�j�F-�6V��jP�\7�̊�66�Mf�շh%C��:S��}��(G���{+I��k�b4'C,26������^Hq]Y�Qt�C�*�ݾ'V	�Õ��!}e��r�n�D;d�[9���u��!���GjgPf�L�� wv��/��I��6n16�i���C��ho9o;�����HQ6�Tv��Ɵu�D ��������r�/-��Ȳ&U� ����9�z�:1\C�v�n�a���C9$A�q\�Z�ws1m����Q��Vt��(鏶 ���@�j����Rr��ޝzS<F�� ����BWPa�	fyZ0M*�3l�G@�8��ˡ��j�/)�klU��}��@��XԜ��j�.��Ƕk%�i�� r����u�l��h*�۾�Z�i�Z�5�i1Bc�[� R�A����a9�
̠��"�ɪk<p)W���o��
��s����9��Zy�Y���
����'xmy�b��	���`	�����
��%��¼C�����;�lNv!W�]	����) ;$�:q2�a=�(�X{,P� ��k�"��
P��H�%�
��e%�<���ͳ�ml{���H�ǋf�{���/%2`���khc�fE�U�ѳO��ŎL�ʺ�� oKEI�&Cw3�75s뾼P�����6R�T���}��z��6���i��C�o,���D]Ӗ�h�M��u-��[k����7�l8�" ���s���Ĺ��Q�X�ht�,m�������r^!u���"�B,�o��T�������PL���|x��)�o&[��2󥊹��<��>ok����Pn�.���j�=�,e�N2���`�;��LwE���x������g>T	u��%n�����YUA���ח���nne����V�{�,��l��m5σEp���/[�BSM3w �U�7w�Cɡ;T��k.����C�v����e�aah�κ�Zch�-K��6�Ê���aC���_Ů�e��UʝA�e�����l�\s��*�N��B�,��!�Wx������R�P���#�c{}��S:��U��)vK�RיB�wKYg��W,�B�)�7�29�%��:՝���,4�P�3��EI�ɽ�h+O��0�vk���՟*
U�x9�w;�5��":3�K@w�]�1�N��@r����l�|�4_KŇ���	�oR�G��/�qޜ�eYu����@i-[A�8�ǝ�G6���[U��ɼN<z���\���|�˕��u&�4~��
J�B���转��ԺYI��Vl'�k����d�j�1Hm�s��0V3�4�����U�("�X:E_�f�5�Ӫ1�Z����Y��\�����d�V/���WP��fIU�Eu��Y�ǨBe�C����*�ok�������Z����Y���2k���X�j��
�����0�EW+ӏ�)q��uu%f\��iԟ-�@�B�J�h�Ս�IYr���-�ܐ�y�q�Ƒ�B3���M]�z��H���|�ڙ�{Gj&ܫ������Y���=wtjG��{����o;��락��� �*��;�Z�fAg`���j�|VT��
w��#�C`Ú�v	1R*��v��t�f��Q��DEj�9�����Cj�C��bT��WD.@&�����Xm8F�'�p�8(?�%je4HSt�Ԯ2��W�z�l��vթ�;�3XFK��R.��Eֹ��ff�6"p�V\R���;$�&�LC��X���ء��K�빼��!���DW�Hm��%��Q��x\�uj�b��!���L٩V�䐑��I��૭wY	�gp��
Y��M��k^4�aD+��3I��ģ[h&
��2�ѓ�jb���Z6��7Y������@��jp�E:�Z���s(yL�h���U���Dl��M�e벜b���E�fòdpJ����O
[��P`W�����3��]�O�Q�ȍz��;�`���R�e�1MD��VSi�u�v6  e�Ɲ�҆�P5��e%�]���yj������@p �u�X�֞�`��+�_tpT�J�dY�x�w1�5ngMw�g�Ln��5w��J�k�<�^e�^NC:�V�)^�֧%�W�C,˺���"OJ�eu��՝��38nu]��ʰj�W�A(ɮ���$�f�+�J���34�Oz݁�]R&++�[�<���*ц�g�1JJm�1+\�-�[m֕	��=�Ś�.j�}xjޏ\�x63G<IJ*�V��*û2�Z�Ӳ7`�;Ge`�����K��˦ �]�X���\��Ԡ��o�x{��{ޏ���V���|���3Q¹�n����S�-$������n9��t�z,zO� �K�<_K�V`W�j,������l�afSC�އ���N2r�*[X�X��_�iݮaIse�P`8!VP���2��=I�fN�4o���������P�|�"E7u{H4E��w�,pX���ՠQ���v�"��m���W[H������.�kO�n�A��GK0쨺v���޾Q�8�T9u�%�yuI��MѹWS n�ꅌ�9�s/��V]��O��#���߀l#J�{JU�˦��yu�Y��)2jF���F�S��T�	�.��zY�8qٷCÄ�7�^хi�lf���z�W���[�%\{Qʜ�:�M�l^�ဠ]h���*�ڍ!Nhz�X�ZZ�n�OX̬a[��n�ɪ�9�/��ո���LsV�۽����Wu+7��iWF������lc���L�����n���cS�8ͬa���\z������FZb9�'܋2������[8+�VX�+�F��nT���]��s^0e�)Ci���2�4���R^��k�.#�K
 �E��U6G�F�gkP����v\��ĚݾOm�Xq�.��:-��^��Uĵ��b>�uy@���]@pd��6d�_��oQ8�U�Hː$D�m�+Ν�Z���[arh��\�6�O�������P�(���%��*Z���Z�[�V�Օ1h��F�Т%�BҖ�����Q�QB����Q��F1U�ʡV��VV��b1��ijհF�kPiQF�U��X��E"¢���Tm[T�Dj"4�B���D�V8Th�Z��آ%m��J$ŴT���F��kQR�YF�DD�`����XZ%Ҋ�m"��R�*PH�b�kJV�m,V���m�j0J[j�ҵm�#mj���(҂ԩD*ڵ�V���p�Q)R�Z�jX�������j��h��QDU�R���U��V*���Z�U�mԱ�U)h�T-X��-[R�-��"5j��1�-R�F�#P���e-*�QiFV*[)�c�l�b� �֨(�+j�Ҷ�b����,��I[el��j)mF�R�ZR�kBĶ�[KEEB�-KjZ��YF%n`����w�w��tgQ`�AZij�:��U�76�1��&���n9�	�j]�]nm�$НNZGl:��)+���t��s����B
�9rΉ����q]?.��$"�\^㛛3����=�f�>ח��{�Ct��gԕܫ�EoF�k�Ȓd�\g(��5���b�P*��ŘȖtJ=�-����;Vx�d��:�<'�F7r��Qn�?]�iex���d�b{�Hr�yM�.��n�Lv�;e���`Go�
u��uqGΗ������FQx�I��]�o:�!�c�	��k#�p��V�<�߹Իd�zBڞ�z_��'�$:a�"�_�2�j6���	de[C6���c13�����J�J��|��_���#1kN�
/u��Ϫ��٭��OoO+��-pZ
��K��'�=�گ���{9P�F�7����!�ި��H�a�9�$�bm��e��+�75u����g)�R��[����6r�.d��w�]�6�>Պ�o0��:�N��������1���hD+2�%�ԥne�;V��8`ś�<:#i�[V�G��w�1�x�;�{&;�5e����QA�4S�[���X�u;u��m�YO��e�Evf�E��
�����)bN�W��F�����{Jߧ�/G]�=
��qǒ�ϖv�0��÷*f�n�7z���y�6�UZQJJl;�%��V:�th�N<�0r�M�9�U$�I彯��x�8�c:�e��=N�h[��#Y�5o���m��i�������^j������3��M�B��f���b˼�3����"���w��I���ך�z��S�%����_�D��$�qe�����Z�vz2+��ז!��%�ڽF�&�Uui`e��;nA�Y�J�����c���쒯-�5�'��`JnK{΋���;q�Z��9O��y��	��8��غζ7max)P��^GmQ�ϑ���m��m��]�0�C�G6%�۞�N�J�#��o�<�>�}8�[��������Dp�:�o_,��n��`�����3���4��Sʵ[O7|���֞aĳc�ux��;I��sQY2@��N�jȷ]���h�x����`m^�a:��;F;�Q�eѶ�)�Y��qhPR71�\.7�Vd�ɫ� R��y���9��[���J���t�65ӗ/M�R�=�j5@>�n*�������٨k>8
�cr8V�p���Z�3���,/-��k��Q{���EY�E�\�)T���5c�ͷ1�����B�42�k�~:�h�m��{YWUWzJޝKf��s��Pf�ʧm_�`yVL�ֻ״�*�x�n뾍�"�"�Ζ���J�ֻy����N��u؄R��5��h젗b�
�)��9��v(o6��b9<!�=X-�ү��8[|}*�� gW����;mf��6q�<�H��ο|{���X�[�؃�>ֵ����-ɕ����m���~�~9��ɴ:^Q�r8��-I�>�9-`�dW�9T�_S��n���P��	-28��u��;-+�V��}��=|�X���%���oN7ѝ��g�!�^e��+��ה[4;��1�QX�m���LZ:eԭ�Q��9N�h��f ��\�	�0�گ+�$��U�E�.A���u��.���w���B��b�Ʌn'��I5U�ۖ��GM]������r��
,�]���[�A�*��9X��0+N��'�k���n��;��N��o"�~
֛5ˋd.�N:4U.�k�?T�_���֧c��w}^�u��a�AR~	���w����:��&"��_e\��u�r�T��;X&z��*�n;!W��GtE*���%�*�F"��.�a���u
��v�ξ�b�(�g!��9���P�A�5A�mm�[�)���W�Wm<M��vo^���2�=��e拼Vs.�Nf��D��/�{X�%���t-ju�-T���tV�qח(ׯ�s-/}�D۾=p��wq�5}3,�J�����s@|z�nFU�3l9��㚷��}��%�H�v!@���֋-��'�o����o��[G��%r���L<⺮z��Z�J�G��l>q����ʇ*+�ǜ�;�y���03�:�`�ǔW{մ��;�L�f����q�9򕞍O
i�v�Y�����-�d߽��ߣg�Pϼ�:����#�8����q��U�$�u:k$�4mGԨ+�+)��k�!,�M�1K*z{2i�TJۉ�=�l�rv��W���:���V�����4l�SM�u�8��=�K�Uǖ�R@qb�l��4+�_M=�v�-�
]3evtE��6��T�Պ����S�Dr�>�wOqb�z2�L��VW'��0��Sjp�J��t����F�a�[�/��5�}C���Ǝ�w����u��t�2��[Ĭ<x>�Z�a�o��/F����Y���14w�����'Xμfy�_KZd,�/�<�=~���J �c5�b<@��ݚ��^�r���x��^�������Q+z��Ԓ�aQ�|ȣ�H���v�n�Z��J�ҬjT6@�v���*q�A��mb���Ṣ�yE«����v�R���obm�o]{l:��ly~�-U�`,��O��R�7�ˍ��5��E �^��"ow�	Nh�թn���FW�A\C�G6�ٲ�����~�f\��H����Ը�ɹ]��`c��ņ�(6n��dc#��M�p�F�̎�*6f4���QJ�	�>괴ۇ#}\w���hޞ��ۡ�y�U݀�:܈#�Ƹ�e�*�l �a�G&_u����ױN�nu)c�����=����xL�ս��Rbɛٴ`e�p�k�3I�qq;�8�R�o]�-\�(/TJ+�8D�52�Q���XK#*��Ţ��n�;���v?��s�-�����f:��hJ/����毫^��t{`�!��T��5��s\�kǶH�7��x�B���s�k������n��+i��f����Y����p�^p��9����5���T9R���u���*ӄ���.�s_�}�+9m�:C��`B=����(@��yo%��nr�pI}��N��u�6�HVU��8[�2�bj:ip�J����U������4��+�[�y����?)�(��!�Y�9�f�ɼ��kI������y�·����X��p1�k����;}��7i�{�ŉׯ�X���.�q:��j�;4���a�o��U8�m���_su�!�j"�i��\���@}{e��n½F�FCo:2kD�k`i��S}�q�ON.R�y�W`Py�K]���ն���Rxc�;��v1|�+V��fM��Z�rr������#���"iH�����Wg%�:#�{՚e���f(@�O�S��ą�xiq�sgQփ�7
�c޾R��ѽ(w(�XĢ�FZq�~�]�(�«���i���qD����j��H'79gv.���>�.��8���dg,:���>�k����fH��u��zg'��b��b��=�ۗv��C:�}�r��=X�Ɂ��xIT��'-�s��fqA�7����n��#�8�^h�<�p�teq������+M�,9�`��z�H�lXH���^S�=aE������d�����_W<tc4�u����t�N�
/c7&wr��Tc��1�M�?y=~�^li�߻�?]��#yH`8б�k������<�g/5�ޠ����y��f��3P�9W���Y⣠n'	mQ咧�9�k:�q4����淯S�v�Vr�g�J���:*���b��Ɯy@�foB����b�9�բ9<!�=T��x�M���V�Gz�B��B�Y�3t_G�QSiy�:q�J���2B�ueaX6�K5��\*�[���Wh��4z�W� �d�֓�"*��ɊPyy{�����uԾuٰ��@��+B�yl��OvC�#ǜ�gB��	��k�J�p�2���$�a��#J�R�3]���-Z��b�mJ5R�z�彈3�5�D;-�U	�l�|���+V�B��
{]t.�)�ī
A'����k�+y+���l��R��KH�ƅ�u�K�;-+�Q�Kw7�M��`ׅ����6��gX+�3�(�a�ZD�[/�k���X��c�G�3�=t	���'�u���nS���+�`U�T�P�Ȏ�\ȳE�9!2�R�j1�Y�J;p�Z���X�c�͘��q�s��]k[��Ԉ��D�=�
V�[ֳ��.��6����J��o��W�	X��/,� ��ٶ�����ya��U�d�{���|��mF'"�j�uF�\�jz�1`��ת���{^�ť-�=�1uX����jQn�J#c	K[�r	F�#sidc/w��R5xՀe�}��\��E��|�A���l�:�q���8�^�{���v+m=�����K�CGVB��H�Ҿ���(��s�o9�/K�a{Y�8t�8�X9!V/����YmM�uس�O���qۥu�j���:��o
��Y���rB��h�U��S�C��x��!�y�{���oϏU�-��hp&Y���^$2	�3�չ�emz��%7z�qE���~h�����V�b�C8���x½�rLU����/U3�����c9׹Q�����ֻ�����qt��\��^E]n'�p\�a��V&���y8���J�F��4�c/���Y�]��8�v����(U�$\��ռ%�٠kS�<��g #�f�f0ѩ�}5WN�����C"�\B����#H�;���'�ǥ��{�]�q��#"Zi�}��|��;8��.�۔:�+.��=6<wR�p��un���-<����ϯ�|������6��KZd,q[����:�v�.ÏӬߣQ�O{5_��vE=������iGC�M.��T�*�ݭ�}������U��&t�Q��Z��˹�U���)����0�oN���Pd)E����u6��^���]N�����'3@�ok2�'�z�B��A9Jzvr���%OMe�;dn�k���INh�<3h
5���Ӥ����z`sBu&�v�Y ����kw���*Vgv��Z�ӽ���;��� T��D�s���ԥ�<:��W�~��\���q�tđ���PX�xU&!���{N�]�:��Z8ώ���xy���y�x���H
�Ĝ�\8�c��n�F!�y-�nR����6k_���f�g!�Z��_�@1��W(z����r��W)�P������Z{�~�ߒwy�v�ߏ���D��Q|��>hl���J��y����][�̭�sE�i�G^�W��em����R�����l̩Y�؝{gt>����Ryr�;A�#�'���!�3�tmsq~>�G��T�[��cw��Nz-}�y=���W�z�#�&�MkB�'��JX�%+BJP���[�lk�x�sj�i����!Y���hz:¾�V+S�����U!]�.y�rN�hR~{�q��0���{�e_�ڜ>l;�.��V9�U.웿��`y���<�J�8�g�VV�U�nd�W�hiU�[(%�eXⲰ������Z����$�n�Ί`Z�$*�]`���WG
i��Rv�"������e)Xn���l���4:���AZ�QS/+��k�)9�\��Q���X.��+x�q� �&qm`���`�u�7�N�=�Z��VmN���wOL�B��]s���v�h0|�z4[9f�vp�ЄV�ʴ�s��f���!8��K�:�*�O�v��j����"$G�}���Z�p��sjf�[��H
X�wFf��>K��3u�h�����9�m̫�b��2mN�ғ��%]t��
]|�tG�-�F�ť�6�f�`�ג�Q�H��bʀc���}!T����gT�2զVN]K�2P�u�x�!���2f���3�U�{A����\;����e2e��3�c�mL	#uvs��K�s��ᄰ��a���+�Bc��\�u=V����:Q1I%J��2�K8
p�w��'� �osĮ8��(G�Wo��Y�k�di�zK7؝�W�{f9/؊Q�|�F�'��&1c'�<�T��\��|*��ᯓX�KUl�fd)Ty�uyQ>G�,9�!Dl<�f�z�Z��e�zHS��#eB� Ŝ��qm�{j���5�o�`�r���2�	q��#P{�٢F�A���u�X[*05C�n�f�W�{uS�M�Cu!t��[����kȘ������yQ3.��B�w���L�SD	��������'���tV�7��jaU�xbzS�QO�n���Fc%��U{�J;9A��tP�	���[��N6����H��&��T�vh����AS������ņ�o+"�S��W{Pi���}4�Q�!�i�=)t:��.��ܱ�n6��q]3�4�ec�i�Op�.��=�Q���!Z��(H���KaS��Vo0_�Zb���������9���Yr�J����S4��8���\�2��^�2�c"����6�ڙ{��)����M�/��n)�-*�U��Ŏ?Z=wAxm�.���G�T)�OA���vE�tM,��k�*�T��9��Š��!лD.�p�|��GL�7]L÷�05�=Ԡ�*V��22N7d�X샇�ᤨvh������6��̡MaB���.�C����<cn���/���1Mɦ�ƫ��O8(Uf�1켭�,^SB�Uqk��)��!���hp��L;kV�!5�%�:�4��Uqo7�.�j�}a�Pf`b��*r��^�}Ӕ��]|�:E��|z8�D4&iAQc3�h��` ���}}D��uƗU�K�t�. ���et�B�//��޴+��\�\�E[Ww(fB�'#�(&+N5��,<j�kDnaY������>���t��(��rӜ��g�S��Sf�A��N�ʘ�9EV�n�lޗǃX=!������v
|������Z�@T ��|*��[AZQjZ�[h��k*�mZ���Qp�chT���h�F-�1��J��e��EZ6ҕ�0�hʔKJ�ډKjѬ���U���
!mjV�V�����mFW
�YF�*�Q�
ŔF�D��J2�[V*����p5�\W�����6��FԶ%mZ�)[--X�k--c)c[mj*�TQ�X�ьD��KX�-)Q
-kR֖�l��Zc��ڱm-F5���ؖ�Dim�EF1�%�J�*5J*(���V��mZі�Z��E�h�Ym���J֖[l�F�Ѷ�2��j��KmV�J*a�Q��mUVV�[U�U��#F��jڨ����µ[kkh�H�EV �[[`��Ԭ�Ԫ����cխ-,P�&�".-Z�DJ�R��Fڱ�J[Qm�ml�VV�m!b*#�jU�+TUQ����X�"��[lie[cj[YJ1+l�*�+*�DDT*�TX�T�Z+R�V)n2���eu�M�pԫ�� �ZY+>z�]�'I�Ԯ�3Qࣔ�&���u��Y�>�}r8L)R�21��fK�N�\7˰�g*�+�[؃;�X�n��M��0wF-���sF{]�67<A��(��1*8���[��u�f�H�40��e[�T�d?�l�\�J��e�߯5_��vE=�v�tr0�X��s�����U��->���^��w�\�7��L�Eb��F��q�X�[�4ɖG7p2ӎ��]�iex�U}@by��o)t�A����L�[��3��Qu��'Ϙ�F_e\����6G`J��e�Uu�sC=g�5��q\��T6���p�����[���dQ�#Ds��'s�ōZvs����C��ذ�e6m�FDDG_]Y%�|��B��,S5v��X
{:�e�b�E���#�gI�Ɖ�C�j��x�53�������cl�#y]�/-/}���xU�玘�Y�V��I��2���wZ���Av�.�������9W�e��	�0fR����rq�����Z�3��ܓ��9��	, k�Ҿ��͉&���&�
T]�f��#3�NIMY���V�ە��X��q.R�2��N��{�w.�$F�d����)�n���f��=KN�h�s�i��q��aG��7�t�uT�hhE����_w6��=�k~��eCNm_��W�0��4Ӗb.���Ҏ8�TV��穭���>Vr�=:B��p�SSЦC�v�����n8�sUꧯեνSӟ;��^�Ղ��!^+SjrT$tNU����N��������C�֜Q䠥��X�[�b8�Z��4�� ����P���]9�JP~Sˈ�KM]u�]SXq*��`$���O//����q�(�=�c*ܸB��K`u��t>��.d�irwIG9���y��w���}|���u���BҎ���P��z��SXij�̮�Mí�P����+�l�|O���_���1.ەF����J{o
���v1����K;~��-E��_����B���	�{��}�ҏ�ۙ<��Ŭm����=�m]�cm�GwE��a�w\{�{[�(oJ��V���m����h�����|n��C��I�Mc6��zs5M|�;䷊i݇:�
3�-K���7��L��f�/*f.]R�F�
�d����M�|�:ya8��i���uL��J����q��gP���ԇ�>�i��'��<I�d9��2f��{�����T��
"�ۼ�S���Ϸԕ��H�pN m'�S^Y�=O&�e�$�a�
�	����ahd:�O{��N �7����lz#�֡5qQ�/�ټ&V����Vd�~׆Y'�4_��VI��"ɷHy�u�=~OO,�X'�he�	Ěa�O�x��f�Ϝ=�^J���V?�M���Y��H)�fRq�Ԭ;�+�<=�2�a�=�I}�N�.�E&�����i�4yd8��<����'d���c��B~�X�����u+ﻳ��0�i�
IS>ٴ�ed=��&�u��4w��O�2޼�$�<��$��O=������aX�������xdx����1��b�Nd_��ƽ����	�M�i$��&��9N���Lξ��N2��14���?$�}� m'y�m����w�ۄ��gވ��q� �L�w`��g7�t=H|�Y��'���M��d��8��.Ol&�q�����i�9�N�w�	�����d��ON� |��=ы�tx�Koﲲ��毱��X�!=C{�(|�$;y�����Mya��ϰd�
ua��d�T�����q0�m�!~��N�a59�=�{�Ǽl?�>�'(�3�M������0=Iǽμ�����^C��'�k�bE�)6�Ls2N!�jXe$ǟbI�V�m'8�2�q��>E��xC�l}}l�Xsh�����ς�{�XNr�I��N�wu��f��x�_1&�C�RCğ3��<d�C�זO&ܘ��M��<Ն�v=��/(}b�__�K��95���{ʷArU�:`'\/�%-����j�q��Rwa��M��ob�)��EZ��x��=B4+�ծ�/�J}�yV�r�sµ��.��x�zS�"�U���-Q�N
qV	(���(N��u��+t�ސ�9�!�=�۠�O���d��`�M�a>�Xa��O{H�4�������d3�gèa��,4o!�8ɴ�I8�L��O#�򏵃��FVg�����\���zݐ��N�q��6��7�z��q�<����)�����i�G����m��8���=�pu
����<���=���l�+���t>��i�7Ci�I��,:��Y��Y6�O�+���z��q��S�N�2�<� |�٤���d�C'���� ����na�'���H�����z¤��%��ğ2z��a:ɦy�k$�y3a�'���� u&��hŁ���0l��Ns�8�Ben��o�����Nj~9�:��I�9��J�$�gx�J�l��<�q&�=|u<��@�<5C�a8����J��y�`z�׬5�RC�P� (1"�u���>rl�g%���T2��;�`'P�&q����3y�$�RO�IY7�|��&�=r�<��@�<�����2j�RW�C�W���TxZ���L}��Ǯ��w���<Hq>�xɴO��(u��w��I�O{�xe�u��5�*I�vE�y�=�pN�m'�Ʉ'O��xyǅ_��f�7�35wf*u������z�m�!�0�!�i�ISS��A`o�����T��w���	�'y�I]2N��$Y>Ձ��b
@�Fǫ��^Ҿnc.w�r��f>Y�����=g�I�P����&u�z�C��q�T�}��N%Bo�e'RzʇyHT��rw�y�I�9��`����7�ۙqG3Wؾ���:<��1
����Y���OsOY�'i�S�<d���I�C���b�i�k�d�T&u�M$�'�Rz� |ɷ�U���0��T��x\�j�Ts�v���>�Lŕ��y{��2�Q���i��פ.kp	\V5�0�I�����!r�mve��t�8�Nv.5���/ͼ���m��M!��ƺN��'�VP5�D�p��%<�AC�\5;Z=������ٺ4F�ӷ���I<@��=�8a<M�Ȥ���{��C�>L3G��O3OY�N �i��:��HO�qnΧ��L�7��{�@��GDXs��InD��I��u-p�'���I��d�'�M��	>`fwz�p�x��Ȱ�6��y��C�>fx��4y���Adɫ'�8����P<������F(�=�����?�������a{�l�}a9�q�����úĝ@�O�s:��{�xf�!��`��X�M$�B���h��{�@��Wrj&k����zuG,c�'�8ʝ;Bz��N?$�`��$�\,$��'9d���9�y	ĆNc>�'�jw��N��M���}��Z*o獲���J?��:ڎ2Z�����a��owC�N�`i&�q�����C��a�u�$�vq'��Mp�:�O̝�wYP�w��'RNQ�z��pG�srx���}[y4^.�Z���&���N��3��I�8��M�Hxj�6��hh��q��<���$�'<�R|��zb�q8ɯw����z���5�3�F뺋Gs{�>�IPP������,XaĞ��$�M'���x�q���m�!�C��d�T4{Hq�<���$�{Ś 8���o��Q��ڧW���{��}���=d��
I�5��J���3�M�Y>Jɞ��8��>f�
IĞ����RN3,>I�L���XI��51Hq��1�{�6�w���>4g?w�o]�����!�4�ˣ����i��8�m��y%b��3�aY6��'�`$�'�SG�������RN3�3a����r���|��s�3�s^c&s��Y���L04�oVO����<a8�����q�d�=��d�� ��I��|��I<;�u�d�VL��u�l��<��d����ڜ�>��q���I�A��|	Ue�O�K� I+�w@"�ҝ�x��`�6X����t�=T�o!�e�i�@�	f1Y����$Y���*�47p�C&�s+]ƂAAv��׍�����WSN�}bf&J�i\�)�yw8�>WFZ!�F	���޵�Uڹ+�����>�S�Xa:�?Y:�z�ٛ��I���`��OPY�{���&Lw>L��I��^IR��r]��&� *kc�K?-��in��~�yG��G|�6��<5f_RN���P��d3=�H|�	��q$�����N �2}�AC��%a�s*ORy��ɔ��>����5lӑF�ʹ��+R�Oޘ�z�_�"�n�7�
��L�O|�:��y�2����Xz���!�W��S�0�!�8��*g�u��R�0�'�Xs�ۯ�o��o]_=�7^����*OY:}�o2L2d���J��q��$Ri���{�XI��ה�'��=L��I�T:���'u�	=C�<���"<=��䆷�oD|��ʼ\�>
=═��4ì�%a��=d��'w��I�&N}���I�w�E&��w
�����jyHq��y�z̤�
L�{`��p]��n������殘%>[:IXq����$�׸:�Ԭ��N2u��Ԝ́�OY8w��I>@����6�$�39�$P�8��{����>J�P<>�|w����?�6�n.�69G��M��q�Hq�iY��i8��t�<I4�>�Y:��nw�q�8����u��O]�g^z��{�!�'��ϫވG�xI�|�d�����b����׿s�vz�|�C�����<���N1@ɪM��'��&�u���&�r]��'_XN�v�Ԟ�I��u��{�;`yǼ��EЖ��P���~���zL0�gNs(m�d�h�0x�q��<Aa6�Ì�J��O�q�iY�Cl�C����I���ğ;I5��>���1wMs��3�DG�e�|�_�˻�yG�1��|�Xq�7@8�I�M�8�6���I��ǔ2�M�Ň6���q���}C�C��a���i'yqu�2�;��c�K�_�IvX��ʥϺ���:u��7@��lT'�Ļ�Q�`ob�ហ6�Bpwf!tb�Y�Ϫ�4�:�sn��[��C:�Qcf��:��<5���e���CF]D����C�T���#r�ӕ/ra]\��Vh�J-�/mV�+�F�=���z� {͉� q���>� �=a�Ͻׁ8�f�'P�8��7x��8��k�m&����ēi��dۤ�B���u�z8#~��>C9`��hY�}�>�
<����$�L�8�0��	�G{�C��&���C�����J���<���lRg��a�O�F$�OS�6�O8�Q��z-�gǢ,fF}����x����Ӵ+��ۧ�'P8s8�!��	��:�ٖM���I8�}��<��:��m+&|� q��=M�Yu���c�{�u�7��:I�&���>�I�xf�RW�C�l��=~B�8���u	�����4��,���'P�%�$��8%ea5}��0r��s�{�q����_wI+'�Y;1�	�OY=r�a8ɤ�V�I�<&hu%}By�8��3�g�R��-<Bq����q��	�=dB=�5[��?Mi��򮯅ǽ��O�c���x}�q%d�����I�זC�S�P��I�35a�
�	���aP8�u0���2q!�^��_,��t��s�����@�D{�HV�o���$�Oo5�VI��"ɷH��u�=~O|�`|�f�_P�I����	�ćP�0�;�1u�;�.u�8Ϙ���n�q$���p|ɴ�O����d�+�V2x�^I0ə�{��$뫼I��e� �6�O��C���4�:��N��OBUhܬ��������6 ��� ]��C�>�RJ�3�'Ru����14���%a��`Y>d�w�6�<d�Ͻ�K�$�3�`�O_�;�B�=@Q��7�!����/R?������2��&MP=CĜAt�e0���x�4�}gq��ٮbi'Y>~I���6���6�z�����m�I�\oR��I�h�D�]8�I%؈���ƥ��@֑�jQ,h���w�vB;�����,
+f�����÷�;:�N�к�3��V����fwV:���BQ[|I�T��'�p�_$]�ki=��YX����Z��$7���̺��(DY�;4����8h��>_���GA���4��3	�)�O��N �gTP�'X�=��a�n�O&����:�߬&��2u���=;�� �虵ַ�f��sG�[�_x{c�����>p���(m2���&�C�a0���P��Y8���I�N�M�a6ì<Ӊ�I��`��}���8A��	:��:3�����2=�쏙7�'$��O�u�'���^C��'�k��$P�2�l�9�'�0���G�bI�Vua��d�Tɫ!��_�&��9$	����,�to���p�=a���;��u@�M?2nw�����4w:�'R��|�OP���!��f�w2N!�k����b���!�=_S+��}��L�Y�;���i=d�q����f�}a:��S�6������]�h��"�����u��s��d��qy ����`�}ا�`\�m�fV�[��4�6�2wVC2�����t�� qO�'9���O��2��qhq4ɯ��)P�3�u�	�ӨVN ���{�n��=��3�w߻���6ɤ�$�3�hm<I8�������-2m&��h1`q��<7O_�N2g���'P�Lv���)7>�l�{� ��I�L}��N�ǅ�Y\�X�	����*N2���u'=O�XN�i�hm����2{�!�l�Ri���X`i�6u	�9�@0��wD�����x}�=�N!���0$��z�J�$���ĕ&�Y3瘓�6����L�ְ�a�46���Ol���a���:(�}�	�&d����Y�g�@h�q8��q��0�m�8�|�I�/3�*I�ޤ��Ձ��pN�m��.��	�SHx��q�P�I��xL�VR!���Ѧ5gͭ饋�s�vqժ��X�jt�[�L�)247L)�[�����;�v
�۞��K��nȾ3�j�nX���������W�ӯ�����ὦ��e!֚��&���(d���v��R�8�п1�ݷ�,i�o�S�����{����廿y���!�L0���6��97�d�3|�:��;�B��'{�2N��y�$�RN��$Y7�����B=�Du�1��Ts�����'+;��ΆXM0����=N����3y=�PY%Lo�d�3|�I�*�0B�����^a<d��=�J��;��,�j��O�s���3̺Ƴ�k�޾����;������=fМI�T=a�e	�s��P�8��*hϸ6�ĨM�̤�OYP�)
�����[޸ m�M��Yv��U_o%����;��"��l�
���]3�)�4�OY�i=���|�Y8����z�P��:�$�<5�2q* c�d}�t�o���*D�C{:�E^�������'̛�q�I�w���'���1"���{�M2��a�<�8��<3OY�N �dՓ�:��3�ly��G���{����"��P!ع�'�y�{�=�L�Bt9�d�&�����O�|��}��C�ׄۆ���q"���%�&�P��MyC(,����q�L���N����w<����g*�g�ɜ���ݝ	��a��0�i�o�:���G{���d��ON�u�:�3�	=`g�ׁ�a	�;���e���M$�B�NP�$��xo^{�e�����Y�:����ǀ�{�p=ԝeL��N��t��I����N���=�I�M�$��:�u�'��|3OP�l�u>G>l��|憐��}�{s��I�>N��b�|�f�8���6��������#�3��!>X��xo�:�.�n�F��AB�Wu�5*��p�]pJʉs�W
s��^j�ox�9)U�2n�̍n"��rv�.�->[nu�+-����a�����0�=�6�S�X���j��w�V�� ��^���-^9�m_����,���ξ��]�uu[qWv,���ŭ�<�T��u�U�+�/5�=�l�0Ù�buce��ޮ��F�uWr����2��s9;�K�f{��,��Ԭ	|oлI���Q=Է���U��݆�t���s�[�D�[��he,�0�k��w���<�qt8²j����D�Z��&�ծ�i6O��uy�I����Y>�%����8�jq�v#3���kVt;��R��)��.��8��M>�6(�Q�ד�ǡ7��d�ת�q�{%�כ}6���=��އ2����.��U�����z��q�5�Xuv�K˘����+���F�h�΍nLܵ���Rqx4m��l��&��]���au�A�[��P�[��#t�6��kˋ]�׫�^�c�
F�/����6Mj7�&�:q��3��!%�x��ͷǪ��٧^�~"�'Ժ'o�1�'�ǹ�rF�w�-K&����ߎ�R}��qpb����L����򷌸�7:*�4��V=��Y�#b�G�1W�\��I�ʎ�{ϓ����qdԙ}�>J��S�7N΀�c�E!X�({m��:f�`��iC{��51l�9n�0����&E�.zHΛ�����8j�i��]�j�X�^�V9I����
�k����wR�ǋ���ؒG\;:�2:O�z���s-.�+6����.���S�P����B�LX����̻�j��Ŗ��x�pԧP'�y�1�k��o,�ww�*JWF�j�,q̑fZ���5��u�w(�\<��W�JεS�o�h��9u��V�5���S��1M�5��fg����QI�٨ݩ	0pGc�O)�(l:d�4��`�+O^�fʲ��+dSm�Tu���l#B;�4$��JP�����%����aC��t�w;c�2r.�SR8�%�^�#�(.-��k8���~~�U���vM��."ɒ�s욧Jt�=���l�9S!�Y|,�ay6�[1$]����{6�\���d�O�Uu�F�9a���)ue��h���C��E��"�(��6�����}�Mt{nqE��X���r�#*ʭ�%�9��)��^њ�}�Zh���g��N�*v�[�feN�m�E�<h�9�
&,�mEb
�A������ow���a�q���JU���`ya̻\��4���,lv��v 42V����(��J��ӗS��r���ݲ�ȴ�@7P��٘���m=����G����s'7lF@����%Ow.{s
}Ms�AYHE4������
��-d�m���L'�Uy�� @E%ľF�Oml��<��0�GVƹ�Zsb}�}­�0F����9Kp��S}Z.�l���L
	l��@�irF	�5{&/*/׻B��=u�9 ��+ 3�]it�(�hl�݊۳���7�g/.��K��ǘ�����.�@ĝ�����}y���k���KQV�Y3To�����X�������s&V�Ȗ���ux��Sc��b��L���C[|�Wqy'1��]�<Ok�.�O�A*�M�Z-X�X�\�/X��C���^,�s{V�Q7�s;W-�5�F����o�4�v��$1Q;;���b�aW���g	�����]9lPI��Т���9t���1-�*�,��vv�X�(4�57{/]&�JZ4�����jd�8�m\�w�T)�S
å�T{j��ZfI���M3%Y�0{y�D�����gC�����EB�J�&4N�� ����5�1T{�Jw��i2�dq�dl�z08Nٮɕy.K3uj��uqs��N�"ٰ0"Ǥ�"��I�Y���ܘ��ƞ�z��Vu{��`I�bM_���kA�}�֫5Չ��d�p
����.+�qmYr�\o3r������Cf��Wm��q|�Gc-[��X�E]�bV1UEX��V�"�#Q�T��UL4Ū�Т+h��Q��Qm*ZR�5��P�ie-X�"*���D-������ZV�È�-ص����TF0ejF#�T�E�ZJ�b�R��TU��Z���E���J2�E�
ZR�UEpʣ�T��[AF
��(�EV�`�X����Z��X�0m�F��R�UV��TT��FҊ �����L �Q-��P�A��"�֪�T���-�1�6`�m(����!mV�Tk*����-��V�6�UVT��6�[lQ�KaUEQE[j��)TW��X֍-�T-��8jbʨ�KT`��U-�+��*��V��+*(�D[ERڵ��TX�,���Q�R�-�+m*"���4m�+m��DF��4��*��"*"�j*���)��U��QYR�dUDc��ڭ��,cmDDX0EX�D��U�T��1Em�������X��}������ߵ��=ߖ˵�{�oE֡���y�i�
Q%x�ީNk.��.�'}Ka�^wWg�˄z`�t����DIZ{���S�*�SO;G�ni�jt {\��/й��N��!�������ׁ�t��1ކ��:i�.k`�,�W#9Sp&�S _�Ks$m(9m�:S�+|��8ܰ������q4����H��}�x�0�}W�zԲj1K�e0эl	�˾�i��v��'����Ty��ᾺN������j\+G����7[�&���6�bA�جLv]Z����U�i_���&n5��+9��Ƽ�,OƮ%Q�Z#��5��y횲ks&z�WSY/)�ʳ+e�N�8��_@���Ñ�'Q�yF[tQ 	�c_l�}��n��kʿL�,ژP�o3\�`�C����xdE�S��3B���s��1��O^�w�dц���g	�t8z�O�Q�a�v%F�LF[��.ŎBT+T"���֌E>���
�I/xY�޶S~���
n������f�|F�=rR�ZԷwY����K�|r ���}��q�����?	�^")}9XI���D�ns�.��+C����^�R�t��m�<�d�f�V�]�l��R���ҡ�g1�^�^:\���뺻�[��7"��U,8E�����)S!yAd�e�n�|�5�V@[b�n΄�u�_��p��36ęZ��v1Y���X��]1����x{�+��x
�����p?�^�|���6(0C1�����ު������5ûh���=A�I��$�<������#a�>�E���Ȅ�V=�J���t��t�5���J��2�_9��槶�@�:"}�&֫d�)�x�����5��c|*�	�Nxy�������W��y��c��Z��D�c����^,w�u9�l+��OlLGs��@��,Y�&��Q:"���f⩌��
�6��#iCN�5a���[]W#t�P�+^��Gos���7�,u�f:�e�d�P�k]��P�iC��c�*�!�1|���u �Wr�Ψ��j�����.�s�O�ѱU�)U�
�Ҥ3��p�;ε�3�Ք���2K��F6j�!:Y=�b��[.5�3����f�ps�NT�(�uP:9=�S��5����X���xy�{n�生b�6�+#�x\)�tr2�Fr�}��Pz�I���z���Z���
�`�\�@P�ךB(��F1��h��c&DU��G�X���ZX' ڥ�esy��1�d������+q{�S���s����'Ӗ�����{*$(��ȯ�S�<Y,*���ݝ�O�o�^g*%�+�I�
 c������d��P��v��V�t�3��Q]e"�m����T~���Ɣ����'`~����Cl�/fxE�����D��sL!J�<��*�@���N:��3:�-�ZQ}2E:j{(S��踟5f^?LtW	����絛e�����m�d��&�۳���0K8��j7[e��f��X�B��m�f'��e٣9���'���b�8�,1�.��$0�m��Ա�s����ä%�YBn1]�䉦�c�Q���9��s��T�_)�7$`��X
��t�(6{���SG�{n�w���Q�"�g+uP>�S3X�	��a���!�%�p�ywB�,'h�;�O\/	v��zb/%��W�Ppo)C�����y������}��#�ңE��|�Ծ[̩�~kl�p�^�"p`!
�1�xU��
4�}���n��Kۇ8���Uf�O5۱��npl��+���N{�f��0�┟��hA�r�������V�;d�g�V������b�K��������q���$Y{qʈ�Y2x�/�!��������a#.�
Q:+4Y��A-4S��Owz�xg�S+��K.J�_�^W��z@�@�>;Wc��	� e�b�t�oD�l��R�K�P����Jk,k���Կ��k���/6'��ӷ3V��쾓���\p(T\2�g}��<��ȋ��ky�ʙ���%v���oe�<.=�+' ��3Q���6,����L��P��3WK=�� W����a�k�i�C�=9�%�G<�6��!P��I���ra."���ݙ5��}��~U4�dVP
�Z$Tb��NJ�e�@[�;��Y�b����Ӻ�՘�ꑷ����4�D��e#�e��tP,�v1��(*��hB�[�SZtr�qN������ы��YM�Dj:�$@p�!=IN�Ae��YB���~.P���c��Ő�=�+��M�kv�`��-��r9���B@���@� �A�g=|&E�=8��Y1���Ea�y6c��ӌ�h8��>~�k�O���	���co�Z2�Q�c���D��
�rj���w�C�Vʫ.�e:�.�ZT�0[��O��S]�&�2G��i�mB:y���ǭ�Vp�q2�W��Yي�S����$�� h���˻��-���7ޞ>�Ɂ��yL ~� pu�zk_�/�vxAv|_,Ea�l�|@u�K��I��$%�OtnyտM�-V�nZ[Z����,���Ex���Mr�t��ްD�{(sò��,r���]a״Y�M
�r��3''w)L��D��ŉ����lg�L]���Gǵ4��Ya���)��Q�
�DQ����g�{��{����n^�=���ܭ���]�:�Y�ap�K��W/���m<�o�ļ��G��7}Y��J�N�1�ْ9\��gH�-lir� :��O­̓��V�W� [@�v�V�6�p�,F0qR�,Ӎ+Σ�Ǆ����"���<�H���,\�	���;Wՙ�32�{�8+iڨ�k����5�J��:�k��|t_�Lp�.����pd�1�;��C��F�)g�2�l�5�=O���������usй��Beiv�F����B���nje!o\أT�o�#J'�߼VRFr舡}M�A�*nd�(�l#��Oh`|����:�Z *pM*�ַ��&�Pڛ�q���*����`Nf����S�Ƅ(MS�5�����H�Q�a�OUg:q�Y���%�K�l>F�
iV�礻���yJ�Y�Ѯ����V��l(`4����'X�R���F�^S�Y(��҂`�Lv����w1��U/`dr᫜ɔY-��5��L:���n�,9�uw&7'�D��8�.�Fq�n^�,�A S����r���K`��h�s;��ek��7��b�+��ƫ���>{��(�f��Us�Co�yE8����B�E�lԃ�E�:.�8����))���Y���*�ž.�h's]�;@�}6b��nHmu�s�~�{���7�:k��1HGh1�x�y5�X���R���.5�(�[��Kx,#��!˅�#��S��=��4�N�nLKf rt�y�~��m�P衪���~^	�=u�+q7�bQ�ju�yj�O��\$ӛ���I���m�c�XO(Y��V���a1�Z�nS�ڹ�*GK�%<In�����]�Pe���pT�=f�v�ژ<UdL�<d<��GWQ����PR_����V���А�"�;�#�\�9<���7�Y���i�E��EL�����>$�gD���v�!A�:Ց��^]�+��X���C������(T��]M�ĖZ�c��V�#���b�нG�N��*�{��5]�7��4O,�b|�f6�Df� �u<2�l�>[���V���H��NyȜ��[��g5�eJ�-��B�lN����ٙB���a@��l�(>�uC���E.}49Z��S�N�Ee���\�\��iܸ`�|�����0~ʱ|+]�gR�$���u5lN:�8�ã[r�嗨�n+��9xV���W����}�c��n٩O�����w�}��w��YR��W�)u��!�ٝ-b�f����p����bW]�.�йrS�ـ�_�Qv5Sk�_Y�0d�Q�kc%%xNLb}O��Ч<{�{�{���Gf$�WOGޖ�d$���-���9�`�����u��ru¥'J��>$P��YaWz�2*���v�\:C�y��.
t��{\O���5��-ͻ��Θ�H!뱓!{�����}���f?X�p���7���NyI�tl�VG�yQf��U��'eY�[]֦����v;%��q���o���U�+��!#o�p9]c�\�U/&�#s�����ŲV�}U"�)� ��ێ��L���] �ʮ3�*�8͐�B:�2���W-��s|2k��n�k�t(R}��%���,Z��KӺn�^��h������f��7ybA��b�+��*�U� )�#��ͮӎۮ���x?�I�0RlJ�3�X�e��+%�W5e`A���T�^�b�81�.����W���7=q���S�I��#�Ӗ[�	[}��N���>N���N���z](�3�p��L��e]��,��_����;�"�;[�k���P:몫X�9����P�fHj�f��n��C55�����ƞV��̶�4���m2�ޖ�\�I�J��멺7��xaT���7zBۚrVj%������9s���o��ܤ;��kB�w��bwi��t��ǡ�r���N���2��$q_d���\��MrzU_�x <%�˩�z��fjw�F�Gd�]K�r�xD��p�^c�U��s���w;���8���fC����=ܯ���Wu��;�,A�/� �X�#�?�[:�8:���y���'ݥ�Luo]bjs���s��mbȡosL�=�3T�j����B�Ǫ�g,�J]ڻ��Z�(]���!7;G�e�^����Sc0���mb7�G*^�Y�X,�E�M�5)e����!�u�@p�2�����2�A�ON2�Y��
��l���}p���/W�U���s-������ ����o3Ai�C�=9�q,j9�Xѷ�u7���أA��s��4�L4��ո����3HFW�T+�zB1!oP8�=�]��N���D�.yÅ��aE����R�;"�d������W�®Z�Vr�m0�ʡ���z.j�c�̒��E�s�^B�z�#x�̑À�h�����vh�C�{:⪸� �*�u�7����E��w��x��H�H|� ��L,7�¶�`� ��m��8��ŠN=!6H���A��o���.�X����^��/H03cC���A9�*nb'�W�H�兖�s�<�^��d -
,өb*a;uݭӨ��^+Cl�-4���:�&w��}�z2���Nܫ�+;�=��/H�7�q6i~���,�,`��b�m,7��������y'>m�G���W�]��Qx�"��ر�9ڰ6z�`�C8��0���S�|n%�S]�&mё<x`�,����Ӕ [ c�u���Zh`���;1������N�rlǐ)d�<�!b9#�1Wz�����eR>1�o�*���(]�}�kαn���$Cـ��14�܋�i"�,���(ᇐJ�n��K��pr��a^Wsނ�̺�%;��r$�(8ǽ`X�/I��`V3�T�4���3�˨�������d��m�F�0�Vk��9*%{�������&�S\Ō�xH������c5O�������o]ὡ�b�u��t� �'`1y@��wcR�3`�LwY����|�c��`gT��Eت�IsK<�\g"*P�e��ӡ�+�x.Fb�;|cBg��x�f��q�q6&�+U�jr��?)1�6��aJk�tDP��� ����#i@��l"#�=�G�ӿ:9�3T-��* �.rj77H�Q���J�|pS����b�VC�A��]r�]I!u0=�wc��o7Y�h-p��Ә�����7�nE���uqs���K�O;WIݍ,�K�͓�Ke�b9�ŊK�s��B�ӗ��1#M�u\Y����x���^a(ak��qί���Y*���;��sƕX[�dGE�U9��*p��-�g�Z�;�H��Z<&2!oZ��Vt�(jsVa��6��2�u�&��ʋ;`[��I�׵��nqد��
=����Ru��+;��$k�b�d�+å.�n�;�i�@��s.����>�
�Տ @���z���=}ϛ�����j�5�ȋ��1�I�ӃҨyC�O\���׺��R��=�X��&A�y5�ٳ�Puz�ty��t8�వ�ց���˅���ݩ��.�!2�ىcj� S:NA��^pu!����f��`-�5Z��6���;QQ���LU���r�T��:Jf�9%ߌ1�m����zӻ�ʑk�<<8>q5�\GL1�L�@*c_1KI��SV^���"*0��䕵S�!�PǼ�^����Q�Á^��j��sb�F��nz��u��6]k;1P_9��	����#���#�M�0w8��cM�FcbƼ&���a��v�=���cIثe�9]+/���� ��pb�Y����_%���:�=HN�;J%�ww���kҤ��F]'*�Tj��3�n���@���c@�l��8��}B���v���b���H�]n���Ƭ�1Z8�����\�w��`͋1xyF)����ka ��ռ�Wш.�� �89�3��+�BO��[������K.����+��e�6֋G�˻��KT�\�]-�gcx���ΘCV+�Պ�v���t@���G1[�c�*�[C��H��$\
�Gr�N�_vH���6��,�L�e^
|���ܛ��_3:��EJ��f��8����sE��7g�d����]Z��ˍw��5ڽ�I܎�tvfU�,[2��Pj�V�nеQ;{�)`�ڷJ'�����SnnM����41f�����4��#��a�[�s�&pܳ����g+Z���M�2��=P��wԥ�o��ձQ�)��v���vCw����ʷ(�����n��^���目�K�s
I��N��f0�5\��g�R�]-ON�@�c��� �f=�:�;���Hr٣���4��'%v�4��M�h��&�4�p�흥��oa+��-�m��[�ӥ��@���i���.���� �&��dw)�X{롍�ˋ�P3����h��|�]_t�#l�c�N����C%���SRpz���)o�N�uy���O6Fvq�tn�RE5ຒ���*���Q���=)eAyN�"[ю��žS���M^��r���5GV�8+}n(ڡ��1���7�[�d:���K`dL�p�܊�bFe�	���SJ��`���l�ފ��+_*�QT�57s�u���G)��K'V���XH˨�m
�O�an;x�xGf;��j��8�(�]NX�3.�w:�k��y( �m��/u�%���о��#��t1v���I&�͌͠yQ��;�)V2ˢjCkf�Be���˚^Ҳ+Zi5�A	G�q}��$xV�Y<�zE�FS��F�փ�Cn������@P6��|o4^��h��m&&T�֮'E
�>ޮ�_2��P�v�X�Z6�C��!Q�8\�9�w�N��2*kvkiQ�̾��cE��H̛<=���@�4�M.���]#H��"�o3Ԩs[ ��S�St�41ۼ�����A��/���Y6�m�,:J�O\��������٣)��EI��rV��� :�qY��7���g7��H�މt�k;�d���&!r���.bKچp�[L̊-�:�7��[�����r�J��VT���)����j�Kq���7�t�p��a���8�*�+�0u�:	���%u�)��V�R��Tj�K���×�1��GK�-J�p���h���lTK���{Ko�6�\Om�/�1��Z�ZFLO�;�>�׺�<6y��ᡈ)�EY�TDDQBҋZUA�U�b*("��1p)Z �#c�Ԥ`�EQPP�* ��0�APR�DPF"�n.b#��V*+��ŕ��V�*#�P�QEb""1E+UQ"������DRL7��#i,���cEQU����Pkb�Q��-�Uf����R�mik
��
�X*"�U	"����F��,`�R�6�m���1�#�U��EEd��+j$��1-�ڴ�b�b�T�mm��EE-���5Z�ʈ�*�B�T�#hPPUX�TPZ�E�m�*�((�X�e�Yj�UQEF�kEF(��J��AQQh��VZ�����a**���1j"�W	`����IKekP��2�A��YX5� �QUF"���b��UZ��lTDX���hU���!b(�L%Y�)�X�F#iQqeQY�b�m��b*�����ER1QY��b��EDъ�����|ּ�(����ڷO�%�,��z���l���^�pSS(�
�Z:U�f�rL�0��U��r�]�.�R�}_W�<!�3�g6zb8�Tdͱ�en�b��OՔ3_ gb��+�o�f�d��VJ�[	9y�ΐ��U�����A^����-�pt���O�X�^HTsm(�}����uM�V�]���n��c�,w�Į�X)��61O��sSB�B����P�D�z��8=*f���+��{�,�'yw*���i�a�*t(����p��\�����He�j��`�;5oe3N;Pe*v{���A���8eu��Z��1�B��TN_bP��.L�yH1I�1	���b��|�q�p3���E���s���N�]���-���Ky��[�lȍ����2��aHս�.g��q<6�+#�x\p)�����GKLX�Y�9U�F�fXh�X�S!/L�Y����V@P��HE|��9�^�H��Ua8���/8���y1̙|�̡ʝ�쉉cj�Qd������0��w,a7--\k9ֹ��n���8 +�@�^���d�t��
�,S.,�n����e�^��I��~��1Ъ᰸�J(Z���CE\ݻq�#9;�O�(ڻ\�n�˦��o�T�c,\��yM�C~͓QܲEi�.��&�k\B���(��k�s�8\͚��7Jp�R"hƒ�i���.�rѓ
����ُbq&d el�Z�ݍ۵]�o������]�U�n�.`pJ4b4*zxQ����� )�#��k��J��_��J[�0� �L�^HO�5s'�u�cbJ��*À�]P2�Q�\�5t���z�.8y����x���V$�g�١.�u���Ԇ��e��YD��ou��F{i��,m�<n�_���ks���k�,o�E�陨�WT8�g	֤��+��v7}P�E^Ş'��G�3��W3z��3��_K�R����y�	W�y��� �6(�o�3Z�ܔz��<绫�ܞ5��*έ��(�\����2��ʞ� ��`��Ì1����r6tJ�g�'+@��^�"�Tn�ntu�X�����)�y��(j�JO�����/V#SN���soGw,R��6�+����ߋV�no#vq����$Y�C�Ԇ���-��>w�]Iܼ�01��c:\�s���F�y<�����U��@o�����.�*댚���ox3�L�;�'���8${3L-�T����cF��^�o��j�{#���v'G"pF�����Q1T���uҡ;a�ޚ�����!C;[kۙ� ��o<���Y�P'�Qi⤙�͋&)Ad�j E�d��i�yrS櫇I��Ֆ�hN�ZQ���w��n�9۰����+�ҷ�7�xx>�ʆ^%�:�F�R���8Uad:�c�Ք��#b1L,7�~�����\���1W���ݓ]�W8���M�CYvaŪ��P��IO`4�HN�A�L�:P0��	3��8��֮�'9"�F���>B7�������L���=IN�
,�\�"�,�1X��-��|���ޥb�mA
�[.yE���b���@� ��L,6G=\c:f�ef槺[ݧ�2��x�*;f�[K�R���y���T���=�gOx��ӏۛ�ݱX���p�8:�Qi����j��W��~��T�)�{=L�p�KGT���T�^��z�BO�a#I+��v�tX��\��[N��q�T���D��o�77�s�ި���}Y	5��:�Q�]f#�o�(]�]�W�O�H��cTUm�u�¹��
�Ɯ�� 1�S���Le���x!e�HyR�!��^[~��:������c��z�ː�e�C�N����&�"$c:ECYa��Q�F]D,ܫp1�����W�lذօ(_9�x��c�j��Za�Y3����:q�]nk���{��=Xd�����ek�g�����-ت��қ�*u�;�Zp���bާ��w��ƺ�2S�pݼi'��8Yr��v��C�*E��� =�f��<=���:a��^_F�5:>ɌF�z��q�)�9�u4><$o���Qe���Z�7I��p�	x��鎾�.Te�%#'`1~�N��r#%MZT�qW�����uklñ�<�F�f��˕pZ�C��3��f�.:t0}�j2�;|cBg���^Z����0�����W;�.��˧n��P(���*��Av�� ���ͩkP�����"�7}�
؎T�h
5�%@�EI��>�>�V�Ȏ���:�����Nn�%t�{�%?wV����Py����J�,s�MY�)M�}B�.��>F�
iV��Cm�)���[4	�Yǥfۖ��U����9���Eds�5�yLX,�E���:ߟH���𰷓���Z�	��������9�r�^�0맄Ss�����?l��{}�iMx�Y���o(4��C���W	�F5䀅a�(:�|\3\�g���<�f��j��%fjU�=��C;�S5N�f��l *:NA�OD�3l:����E\^ O2����7�~����[ߐOP�Wk�W�[� �h���uoa;˜f�w��b`=�"EydW1�M�d��n5�'��i+���P�7�+	�mK[-gB������K�; b�L��9B� NXf42�����a�Ծ��q]��� �f���[�ڳ	eh���Ӂ`K�c�xfdX���j�(�۷cذ�P�u|�`N���2	͕~��H$��b�6&��aD�AAVEy���}�&�~-���;#�x��pE�(�����
�.2�Rk����kTF?��c�UB���m�U�;5`��񨾽���~e�'t���3C�5��@Ra���FcbƼ&������r�a�g�u+3�I�6�^��]��l����C9[�����vb�ޫs;�T� 
�d}!����.�ټ�s��yu��v3��UW����˦�[���8�V�s�B����/j������٩uT��G����\Cs��}:b�X�쥂������o��*�{��)�r�y�_g���"�:W�_��{ ����fv7x�@�鬍[Q�C���:�˨'S�c��Q��u_rΫ�u���],��i�zV��c9�`�'�H��u�XPA�!�-��V���̌���jβ�JtB}L\�i�׼ݱ�㼦�R18Gd����;����}u�j�N�Z���>�\�ĩ��
���F^��tl��"�6���vw]O��Mpy�Ed���9���B%~�����mҳ>��Y��j-�������9ip�
Cr\�j���g�9z�M�Ռ�>�R!p�ں��U���{� /��M������H#�I"4��}����R5�{LBg��b�6�&;8[���E).�	���`p���q�fXh�̱�J�+���f��Q��6�Q��4�("D]N��m��1ѳ���O�:����
�c�&%������*
�����U�gP�u(����~�����V8 +�`P�������o�K��E��:���
8؅�]��G0�y'ܜӂĸq�N�\�<] ' �Oy�Sk���i�:Ӭs�� �bg+����J5�F��P��%�sa�ꈗpzC�������^��P)��Z5�[Ϋ��N�F�!�e9�c��Uq�}�&TD3�ԑ��u,GL�m��pP�mL�J�;���N�q�t�+Ñ�;��q�	���t5�UWk&�Xb/�_� ���^���[�j<�w������\�J��M��@e��K�r�p����>���X�`��ח��m;�r�%9< ����<��ϳ�)����P���b���j�����Q��+�bg�46z�'���Zٛю�,�MԚ�HZ۠»��g<6wO}g�n6hY���T��J�ܖGs�����gի�u��Bd�1���9�ǝ��3��m!����νļ��t�L�KH��m���T�vݑجt�]���b*�e����,��������5��u#ɴ.a|��2/5�1��̝n�8��`�>}�$Y�w�}df�ҏ`���Gm��գ�u'YQ����	HK�3���̲jڦ#r���N�����{C�l۱��M��(#OU���B�
t��,����UHY�ONC(0�!��>VNDXXxS��ڪQv�����lYyHRWK U�	xy��Zc��~�����nlR��+�|�rwo-�a?+�B���I��9���������/Wer��>f�qW�&�6=�S"Y��::�ا�X9
�va��UB%@�锏d�Cd�(l�D�c�#3 �ǆ�9��E�k�!5��AE����rT@�Q���$@�.bz���X��D�Im��nC�-|ꍩ~�L,ͦ=5�HZ�V��:�s<X	�������\;_7��ǝ�u;�{����蠬�{0�A�i�E�v�p�eY��T�����HXv�=�{8�0��w2�z���⪘��~�LE�P�x�N��{Ք�g
��e��a��9S{[�+_�IIR�EJIs:�I�N��Hc�*e����җxN�)j�R�vvP�w��t7ǚc,�8��i�"�����$o`�&�^�ޭp��g9��e<K�a��6S���ھ�\ڷo8:Hf���,�H\ yEuoU�.�u)�=�c�x�������S��Gђ]�F����N|�tX�����N�b�i�͟q��-*]XjQ���R�5�d��������>��.�WX�d��R�3�|4c�M�P�f�!�ߗc����,���iuW��3/w����Z@�͉�%$eCyW[6k�:�Y��ļ ʑW�RΝ���w�[�|���a��S�[@�1�����TDc����hۇ�
Ftߋ�n^��'wW����bo�˽�2F\�FP�!�� �2qe����L����3��Z&N^�m�r�f��oWF�0��ug�Te�%�9;Txk��#�,��4�o�@�=�����[���ˊ.�keJ8r��f�P⅗��fK���t0a�������gT�.�S�w}��2�ip���+����d��VRFr*nql�h�K�B/���9aiƤ[��u�cXu�hg��o�hC�Ҏb�B���c�s;)ruؓ��*r�#,�����*��9�����H*s��o�j�z�9ӎyVd8���(FuR����B١h��=�])��Yֹ�'.����q={"U;s,\�"���g�����ܬ���-�b��qiB���.��ϭe~�P⻌�Ws��E��Fj�;g��eDMM�MY�oT��U�x& ����a�u*�]�%��wQ%�[4Z����x{КS7M�Ol��[nf������a���Ȭ�t���������h���ђ�<Y��s6�R���X�c�����k�*/z��}\"����5��'u��JsS���j�h�{��"����q0P���0�Ƽ�%͜��yo[�y���{i(/�L��ue�,+�މ�ᬇ]+:��y�ĥ���/TT&�g"�(y�}R�6&��lB�%���A:�vr�i�#-S���7�fE��/�����S~����)U�����=�I�=�S1�	��F�M".���T�����-��cG�J����=�	W{��M���E*��$���ɯq��Tr�zE�TFӛ�0�.eŚ���S)ze�#�{�+�3գ�X'K�2wMc�LΌB���e�*L8�5^�F�m'�����������gAHg�!���WL�[��zW�ֳ"���S�e���ؼ 	(r�5֊�b{Ϩ Μ�q��m�o�*� ޛG�َ��>"U���
�������rkT�W^R�y��D��畽��Ƃ�(ئ��R@΅�%u^g=<�zP�bXiQ����oi��s��|^̐�Z%����89�(>8�{�9�.��tu6�F�ڄ�uCU+�n��x��(j&��0}}�ws� {���LOa������Jg4���n=E��6+(z���S��Fm71�3��a���w��&]��d=T�i<���Opt��V��Ärߘ5��t�?A�`����{t&�wz띀����A�)tX�t��	�z{|�]��#Bv�F����=�c�llGn#�h��9�V(P�R�l�*H�P��}n��l�^�!��\�9n\�32��v�Ŋ�W%j�Tc�%LZ9&B~��J�rs+���NyI�+�`^'f�+���ى��2���.۹,>$�1ҪM�vO,����k�e�E'ޫ���U����X�9��
WLk�dȋ�r�P-K�;"bXڋ�E�L����N��^e�f��Q�
/$l>:�N�pDc�+֔_L�t��P�`��	��h��U�m,��A�3�,pyG��E�a���E��}� )|��ؒ.�t��h�͚�w'w5�f�w+�V}��\�8^r��Q>d��[�a�Aa�.�2
�Dg��ZS2K�8�����G*dށk7G!܀����T�[;x{e����r]@f�yb#��r�wM�k ;E�.�q>���6��ڳ7��Zbғ�U�(���r쫌K�K��[�-v�	O7�:��J@swR�v��ŋ�ݑ�D,�oE�(�Up=YKu�҉^��`Μ2�>��fգ���Y�=	�ox�r�*��&;�Uv:�Tb��!��#�R���}�e���2�0���9���V�3]��,ew.�b�vr;�8�V\�z����y[����֥�ihu�m�՗��moĂ5+eH�u��%2��&��v�m]�����В�`hn3��Ҝ����\�`�%�%!��^܎��{��������51��v֞5ŭ��&:�H]۲�<���k�i��LR���9�8���{*t�̃wd�B:��i�CU��TU���E�P�#f��v���ջ��<��r�V�"��Z)U�P�_ˡ�kM1w.�i_7'T��,����Z9���D5�{�`��O*hk/��G3��-�v�]�ߧӜL;2%y����ol�(��\��ہbr�T��+��S;y9��\2k�u�;�����^q,wm5�&u�3ju\nVէ6���֊�8��-M��(�^��f�иM�N�/��]�A����[\l&��+���؂W���f���r�8ecoE��K��2#D�jE��g\��
S��w[���J�]rtUט�cV�\˨1pwrژ��1V٧W���V��4#���Yz$��+i�I��P��0�9�������V;.�Τ�m�8l�xm�ܛo6��'L��wJ�,!�y�STu�\�%%�\�l���x�Wً2�!BL��H�x��n8���B��9rK
ip����|+z�����5�#�d�N^r��	&��YXB���:d&����΁�vec�]��_!h���Z��i��_
rP׭FM(�Xʗ�*���o�]5�7$���%fT&������8���!]grp2�J�*�b��홸-��;�-���K�#-�VDU���i8�b�R�5m���6��n�ΐ-TB���ܣ[S+�ֱ� ��;r�zBmkZ�)���r��rsE#�f�P�0Y�,�,��e����^�;>@G/�HgIt4N�ҵ�Z.��Z)\�F�u)*���6⦪�0��}�kNaU� �B�Wڧ:.Ҿ�l�xb�֏"�'���1��ڷҸ��t3ឹ�hM"�:��7�Y��Rs�������9IC�ߖ��f�c�Ѓ����X�W.p�ǀ���!����b޷���(�R�[Σ�t�99WPV_oY�i��a�k:�3$��Ԕ��N���:$��Im�3ul=k�������GwA�·��
��-9�u�ܺ�.2�ڷ���$���TMn	�l�q"b�RL;�a7�N�a.����`�-*��J؊�UF�R+ib����E�T0Z1n11��b�jх\.*"V�F���QXUQDADQ�#Lb�ACE-��-kT*"(�QAX"1X��J�e�ETB�X"�`�TU����LR�m�`�Tqe��Eb�ְTb(�QQV`�TeJŌb�؊�X[`��EF#QUDTF"��E�qJ��(�X	m�lV(,EQڈ�B��*��E�Ů0Q�UDF,T*[Ep�����-(�-Ub,TX���AV �4�YX+�iT���#[�����Ub"�J�+�����QH���a �jR)�X��F(����VhUQ�V�b�DUAX���Te��ca�QDT�H���%�
")Z�(�"�����c�0Ŋ�Tb�#�`� ��LX������a��"a��QU ���DQV(��R+!l�A�T�Y

�j�h�T��Z��0�eV���EQQTŢ���#l�V$F**2��h��&c\�0�Ö��n%l�Fl�9cw�ƭ_؛!gu�̾(�i�R���C^�z%��tH�F����xx=��e#���?�]tn��Q�0���=V1�ڪ�k�m�ݡ�C��d`����w��O)],K�����.���NV�)��r�Ꭴ�]*�k�u�UU�&���7�'ǥg,�-r��� z�`bq��U|�CƮe�Y�.���J�D��p���_,�;�Z�bObл�q�+@/]h+z��8Ԟ5���~ol�q@�5��p`�H�ЬC��M'C���f=�h�����7�d��85�*{9�"��t�po��������S'���d��)��cW�������D�b�WC��s�p9�M�,F*�����F���9����@����v�ڽG�ԓ�KMz�E�E��r<�P��Q���yl{XǨ��t�t�j���wr
gCK�����|WK X��=y�L*�饫)�c���e��QZ��ct�XѶ��
�'Cp���SLvVP
�r�#�gb0��Zݜ�{o"��Q�G7y�4@�T!Oz�����0��L"T��H�I�6�R�YD�di}6h���a�T��u��,��� h��.EB�^&��P���J�cN�]��������l;Bk��0����o�1W[q9��}���D "���;��۔&��U�c"��$SM�6�O��u�m룵����9���+G�%o|< ����d&ͬ��J�ЇB��# 8�� gtk�0"�̱
�:��]*U�Ssxn-//���{�ۇC���7����c�Y����l^E7�nπ�	ڈ�L��&���ޛKR��H��o�E`���.�g`N2,�-^��9�V��`���X�<�10]ȣ5���@��:K��b2I��(����NՍ�z�S��D]�JB�bP�qRȸ�����>'�>_F�y?Wz%��[č'>O�E9Ip�X��/��v\�7����_t<�ŗ�ʴ���)����@��^�/IuUB�$���ю}M���}�>��ߗ�e�C�k�ɖ�'�2oD�%$cw5`,����͊�0Int-*�}��rvک~��o�1���P"��B�������{{qB�ѷ�S7U/6��4fz�S@����3.�^��~:J��2�2�9�A������c�:�*!��ң^�H9�'6��>��tփ�k�}����u2OP����T��v3%B��R���N���`��)���dB�G��������8g)Sᩅ��tH��Tz�i8����k�z�wǍxy��u]���������^sDu�2����d�]��*Of�E⢶wf�T�!z/5������/N[k@ΊÃ��db����	���{�&���AbOv�c��r>���S��4�[�*��T�?5`�ƎϷ���.�KL�@~�6���K�p�0�Zq����3c�h��؞�ee$g"*n�t�@�R�=�I
�ЙWs�A\��h�o(w��o�h2v�ܺ�B�{_���UM�I���(�9�4蛽�e�v�a��AהƄ,	姣�OU`�N9�2Z����J]����*�W�yI�e�7cM+D�,<�m0�_m0َEk��W9_?-�Ąp��uՙ�{9 ����	:�����.�e��Y޷���g��B�Φ%�k����NrU�]�W&%'�d�����Wkɯ�f�z$���1��J��R2+r���&�-��2�k�",�s
dݷ�/�K�E@r���p�����l�GL�심��	?�uxk�p3��gΝl�z�&��|��/ʵ��f�!\�H�F��U@��ʓ��^�1�}�I��Wk��Q����)i4Z;`��o���c#s��1�Wwx��;��)�V��^�T~�r��Ή���<��=�DX��q%V]�0��L��`��b�+;Bw�s����Z*ַw�TId�Cf� �A;r����5��|"�b�9���u�1p�����xzq�����}L^l��8&k�L95�\�^�ԑ���,�a�ͽJ�v��`�ˀv��V�^K������,uz�m�N风�35�P��e�>
L8�-���3�J��I}�f���TXC8�i�w*2β���4�ld��BoU��VU;4V=/A�N�%�g>�_ �jE���1��T���^(���Z^�����+N��X��Y��k���)�Q �X�t�u�HRzv�bWe,ǡ��S|.jc�
�˿��jۙ��(��or��D7::��PƦ�����;��6;�Ǧ���q���l�hP���;��y5�[�u6��x0@5��1�]
Nڇ`*w.�v2T�u<������9#����L�.��^����zj�������k�yo))>�r����g7Lc*�h}�%�掷�x�L���X�V��w���Ԋ6�Dq+����xR5oi�L�7�נ��Qu#o9^��\�E�l
�E<��Rtya�Ic6�PD�Q�*y��AW�6Yy���k�Kd�]����\W���1��b`��N�W�ѱ7N�s�t9+;�"̇.�@"�xs:�Jއ�R�G}woPfr�}�vs<D�����%��'��vE�0nA�vV��0��ݡC�L"M��	c���p�tMw[�������8�녞Z�J��q�N�g��F��{�c&D[t�P��ێ��lW,�t�P/����a�����\�^gJb�¹͐�����V9�^PbZQ\M�Դ{&%��;�
�)���]s֭�6=���U/�J+�d�����)m��������踅�v�䅴j��k��ś�۪i����ᓑ��5΍�co¥�&����Q.����ܭ֤ty���Y׻5#�˺7�%��%�%�p�e<��c���	����B��r�&��O�����D`~u:,�Q%\�"��aܩV��k�k�R��ff�VPĒ��k=p�f�7�s��ظ�G	|��o.�O�Y6}(j,�Ծ�p�����!.�8ِ_��[�{b� �t\��OK��/Czgf�!gD�Y
/t�M�"�v�!�E��B�v̫�+�_��FE�������盭�!�X.gM���7����U��D28o^�_<mv䍺u}�yw���X���qrlG2�^����Sc0���)�eo
	�Bzv}abB�K��+��Aㇺ�l�)<���Z;+.¨]v���~��uy�����V��sf�|��nR�hq��5lr�
�)gB�;����[Ii�}���Aι���N1/�Z�W��גR�U��_Y�/5�'q��v�_{ȫ�������9їY�YdP�}A1�Y�r3�UH\A�ONy�Zz��]dp���k]���ë��\�}!
�@ۺ}],Qg�@�f��P,N	�ҔZ�++0d��|s���S�2ƍU0���Rpcp���u4�dVP
�Z$TF)���(�c��L��]f�ԓ����>Dp���w�
{՜�FXa�}�) ��R��E����ٝ-D�ek�Ufe��8�и�_�[呁����@޽y�0�(zR;bgg٢;8�pJ�����o���}N�I�J;3mǨ^m�(�.w�s`&-ؠ�ݸ�S�����x���@�;l��a��0�/��Ar�p,X�0�U���R��
�+Ǟ��Zs����yj���:��gI��h�֏�+��k~s{)C����7vb*�J��ԓ��ҽA�]Al�
d[�,�K�F��O�E9Ip�E����;S�昝a�<��Fykgh$�8ݸ��5�zn]��Ȁ��,_��Xl/�|)}��U�c�jg^C���7�7��)m�����4�H�}e͇w�UyŮ��*��qBa��;�׀-��sA�`���HnԫBƍ;������J�e��X{�}������e�\ܢ���$���J��T8�b��CSɎ�;3����;>�t�U��\�Dq�|�廒��X��w�N��y.L�`���P%$eCyV.rC�B�I��5[z��QYa����s�CCW1¢�r� ��"c��b�y2�L�"����!�|����ڣ&dUM@�M�X�ݗ���Z|*��<%��z���=B��~'�y�`уL�7}�����{ȩBC�Y�"�HΖI�*�{T�la�
+&�Y���Z�ī�|e;�S�J�s=�2ݸ=��Y���ٯL�oܶ��E�V�ׂ�����j���Ύ��� }9��r&��MJ�|��Й�.����s�4V�:Ξ��U�R������s�8+�.�Wi��.l
m�}I���u�;J9�TT��}�=*h,�=��_D��B�'������ p�(����S�<��j�s���qaQRP�#7!ʼ\��J]u3�^�ٽ\�H[$7c�*�k��e�����W���+9��+�V
˓�wؒ�����Q�e�xzLuK��q�W�#\�^���+�^�w��@���MJ�ҷ>)���P��ζ.ƩQ{�.�lp�S�g%�KD�x�[������UK.�:r�T�t�l�qµ�+,tN�1���7#0��;���ݳϝA��L��4���MJ9"�Wr"Wi�ZيIvx��ײ�l���6H���{�v� *W���1s�ދ��µI��E��/Ć���0�Ƽ���ؒ��i�hWU��-L�T?#K��e�d����nDiN��n�nP�f�B�u�9PǯRk�4^,��L((u�*5b2�8�8���������t߆a�P�SSD�����*8M�`#�䗦ͨ�N�M"-L!�*�BP��Znb�b����\�rs�Q�!�۽n�����=�$���.�LA��/a�̌~P1�*��N⡾z=�3�I�e�H[8�ٴ�\m�t�9;���צf�
]��PcnN��ŷ<�N�8��$X~Ǘ�A�CP� �o�<-�L��Y˩p:4�p`�V�S\]Y�$�:h��q�'â��:�\.�:j��#4ל��8��1������۾�7��WNn{P�s".�Z;;�:��7�o���:��e,ǡ��.�}���m��:�P���=��҃�N�e�P�ŽT�N����Opt��[�j8հ��uH�Xs0٭�c[��%K�,D[��,�Y�s�ܴv��kw��
(jq��\�����լS�V�C�b�@ȑֻXm�����i�)@��~;sS%�����ھ�w�$n���1	��3>��G����b�u���5��o�<#y�Oco37�dP�'kD~ΥNڇj�˃��d������v3�6��<�i6z-�puy��^Όs�uƜ�!5Qd��Q�A�[(8)�ӕO՟('\���osVX�zws���(#J�f�B��D�m�TȎ%p9��d����{n+��ý�ʉ�e&w�l�n%������F�Hq�FXh�K�$;)*�i�徵؟/�>��kD��v�����d.���t���r9#X�u���mәB��n;
q�+�LL�]��#:�pщr�"88.���p�Nl�����|��9�_��)|���g��Ѻ���	ks5$썞�mLuq
x�-�åO�o�P��,x:�`q��"� �*��{,
�Yw�L�-�V�Jy���ޜ��fAo���bX�Z���\��pK6�T����qņ:֠���hʺXӞ�@�u��m���܊���J���N��O<��Z[�MOQ�}feAj-{&n'n�vd��k#�Ѯ���c� \`��w �Q�	�[���*��M{!.˧i�TW�o�2`���6
T's����xr�hc��ʐ�eyh����=��P�m�j�7̊�ۍ+y��	���PB]�fK*�Q]F�jY�u��hu,pVn<�2]�T%�&V��5�/kjqYX3$#V����b�]���b�Q�k�ǿ�0��떷(X���c�XިS�%�p�Ѷ,u�g�j,�Ծ�p���Mƚ��e��	��e��x7� {L�I�P�:��8ho�͛�+# �c���aTv ���GV��ñ�H˝������#"��٘�hfN�[@k�oI�
g\X��Ln��4�I����U�*<9��ՙ�#Q���t�8,s,��j���u�t�Z�8�V�����Z�R�>Y����P�X�I:5S�]A���?o�mA�뷲�/��F���U�%ڊ0Fo]!�骰�w#�HF�w<�cfz���%�X(OL����mt~�n�o+�c��zr;����2ƍ�uW��)82!�ua92��e ��-:ĹU}R�]ᘻE坁t�9P��!��Sެ�(j ;0��PS(GL�0g[Z���í�~s�%�&9��Χ�P���((�X0C�Q�#x�̑À�F�ew�[�ǖ��=Ot�0a[��(\K���\�ٛLz`^m�!E��w�s��Pǆ�U\;�@��^32��/EKug&�ŎI[\\k�a��g��ut��s�ڡʤPb���C�-<7�G;Qe����7b��E/u�&s����4ڮ�����2�ÇG_n�7YXD(g"���F�t5�
��L�z3Vz�+癰^���wC�1�j_B�������޺�������d��r��Pe��j�s�/�ڜ"I�(�d���AC�����L\#e]S���d���N�{$cv�]� �P4�:�h�	�"�Y��ݭ���ԆN�6����qG��X�)ZN���ul ���TBv���'�[��"��5�D�i��%wc���W�2rz��	�v;Gm�j�a���w�Jƀ�0��;�M�+����r����ѽ��s���I:lT��r�Ij��,�e�jY�Gz���,�9VQU����_e����C!��2��rnc7��*��l]*���[�h��u�s�Cѱ6��a��76⽕�KuvuSEEY�����$�ɴ{.���WWZs�l.�,��:�E�u�#S�緃h�!:8ceT+��7�.U̡<T��V-f�x��OtZ�ٷ��5q<�6W���^͗A�jJ6�ν�
�D�����ͪ��ɋk������2�ɩ�t6ɷ2Ը��e�pn�!VmY/	�\.���0�jб�#��E�0"�y��^��,�.�����c�2=i���K$M	&慯g<��:������䉚��1��3+�y%-}��ޔvç-�s:V$ޫ��c�B�r[k+�v� ,��nv�"]m4�j�+���3:s2�6K�]�1�%h�7����\�XpsY�# �$[�8ŨꑙxS2�dԪ 橼�8X��s�и�n�Н�Oܠq�q0R�5�yQ'�Wr�DR�K�o����T�E��+ى�]2^l�wZ�YP���E������{]�Й��+<F[ u�L( �X/���Z�&�VSV���.�p G5uث�}}W��s������s�j;�)[q���v:��VuS�.���#(м����1�7{"D'G�1N�.���<Ýż8I�)s��V�	�(��r���g�`ݳ/6Bӹd���w��U�WGA�3o�J2�vm��ֈ���oX��Nm�[�gx���"�m,�,v�
�iYv�*e�Ve���]�{���!�	Q�m^[��ي�rh�_1���%� �*^Ju��]	��C���5���GL[�PT���`� 7��[���B ���Ӭ��R�9���X[�Ӿ�������s	ݣ�xd�0�Q� c���:���`Wu�P��Y��jT�.��л��N�T�{�p�T�<�6��F��/sU�Mr�f�2����r {�\u�%�s�P� u�RO=LօF����w"�m�e�_Q�����m�3�}2lɓ{��
�7x�D���E�QEPDUQ+,TDL5���j*�ZUb1`*����iTAb%�UT���B,Q����EU0�"�*�`�E1j�
�iE#�
�Q"�1X�1Db��X���EQ�1UUPQT[K�V"�,Db�����"�QQX(��A����������X�E`���0b*1@U�"� ��""�DQ@E��U����Ed���**0EH���1"�0R(��Q�b`��F��Q��X��
���*"�U���PQ�*�QQ�*����TcEX�PDP`����FT*�*�"��1b��1DEEEX��
��*��#Z �EQX�
�T1�Z��UPTDVE"�Fڊ��+b��b�X� �,�U�b��QUX""1Q��(���X�(�QQ"�Wwt\�~{�I����o%Y�pǗ����1$��r��f��k(m34܇(����e1�
��{xx���vM.�Wb����s9�l���FD~��",!��"�ɰEz�N�.�g`�q�c���򽵒lm��[A2z��8��6<����� *}�t���V��\.x*�G y�u��U��P� �ޮ�f]���Y���:e
T�S"�,ܒ�o�K���S�Ip�E�����'g��1	�MG��N��u?=�F�i��*!�zK��zQ%��*'�떵�n�׺��W�F�L`�ָ ߳}�+6=B��:�X�u��%fԠy)#)����e0��D�8xc��|��FW�m���;U�a�AE���B�P�n�p��ߚ�"a���	�3kw�a��w�*fk�'�Ĩ��b��/>O­̓��5l�KU~,z�
g?}��)�V��\���%�N�u�1�ݫr� ����j�H��W�3�n��\����(7��e�T܌���G%��j�v�z�����=�~�0;��ZJu]li�(��iV׃�E���!F:�b�OI��d�Ma0��a�e��@ЙZq���/C8F[�o�U��t9�x$����i5�۪�L.:�گs< B�+�����J��6l�U�%oн��Yʜ�L%z++qT�ͽ�o]Gcr����I0;�5w3���t���#̦����i���R���Ze)T�e���c�S�:��.���Z��o���}q7��z��G��nd�i@�[aGR{C+|�b�1�j��i�������=}�U�U�0�ڜ��Z�ȍ�*�͌T᜖)�T[|25D�S��X�Va����jW��Y�U�u;V��0����.L-3S1����b���_l�܍�~�+����@��o1e�����Z/^S%^�(!~�8eG�I�������J~�^�7�H}�ߖlE��|�gV;�g:������'�5"�n�d����B&�L*��@C�g]p�6��ٻ�K��/�0���s�1��q��axdE���)�.ݨ���*��������ze	Z��{�Y:г��J��:(j�bYb:����\$����~|1�A�(�z�nؕ������-'���W�z�J5�x�&ރ(�SiS"�*��K����7ƀ~)�l7Da�ε~E�0.��=���Q���5�#rEu�ԃS�ݗ4{��zD��f68��ؕ,s��G��{�h6p�g��Ք2���Z�����Tg0+��RٛX��-����{X���"����j6�bj�{wLlf1B�4ia�'hД릜#*R��tQl�z�㳰j��O�N�����������[��<��7��3�C�(�(����t�X+8(�<�L��n���)j�B[�%t���O<Fn��������4j�����j���ć	�3ҽ*�d^�Z.ov�N�&� �sd<Iʍ��^�$��� W�;�3v��l�U&6�����F_��0�v
t�R%4z"��OE��U��Tgm��F,g�u:�$):pOn=E��K:��)m�Y�]&�ma��r�8�̋�A�'T2ڨzAU�վy]؞��"8��ƃ3y���tb��}�q��k�/ޡb���gR�'�mC��ܸ#���)�{<�8�M)��CTu���Vnk��h�j5��CSF�MD�Qd�E��A�O�١��`�LOA�ҼZ�ϧ����WKcY�;�b�۹�Θ�H!ة�S+��̬7R<7uz�J��\VĜ��T��9#X���u�����,�0�\>�*�Ɛ-]�"�q��jw4��.�d�Y{���@P��HE|��x9�k��dȋ�n��B�n;(S��Ι�A�ubs![�}��Nh?fK�'iܪP�Nl�����啁�@N�΅
O�=$��׹�}�.܂/�/JӬ]��tU��R�[�N�ɢs�q�8�F����Ek^�o,� �靎n��Wp��8o]%���*S_�&��'���a8�0��������
f��g/wI��e.K�F�9P6;Z�+��|�×3r�uZ�1�8���f��|�������{��S��NeŝY�/�J+��Axx>9�>.��1�:�v���7�@�۴xM�i�t�v~��G����Q>d����BP�$�ᖥ���w��$9!��[d��3�/���s�~�Cj��׶\eO0�wv�ՄM<IM���r���KU�O�@T{�l��I��Z��
��hS��V��b��᷉/}�TVk�P�C8N�'MD7�t,,'��7ʉ����Aƫ
z�O��;�����j�|pߨ{(�wOA�5'�>�5��y��پ�L. ��`�+)$��8Xq'�׌e*�Շ���csfc��-�F��`��9:v��I��S�����)�������O��N�(1���W�]̲i���;�*lnjU�r]������K��{C�~��sɚ>\jU��>���K&0�W[���P�|x�jJ��e��i
��-�5���2��I������ڱm�;�������A�����:��edw�lFf#k�߃P�9:��?L��d�vH��Ƙ��\�=��x���d���v��s��̈́qH
�R��v�9�S�Q�"�p�'MJ� Y����X9²*��]�U�� =z�:nII�:Ԍ��9���3�e�p��fT��nXY���v���[��bM?U]�93F�935C�H��V^���z��=��pU�<��|�q=Bj]�aN߱z�A7��孛ԇ8��<,�e������
�"1�u�@י0/$VaW��f��FG�gs���U�vtVVT���A�:Y&](�ͷ�y���uߞ񷎺*>�<��<}/����b@qiQ 1,��Xj�L*��zC(\��7��z�:�QC��"�����[�t����)�}I��fe�8!�&z��iA�N�=��Od���Po�[�Гv��;�3,`�a��:^}%��#Ii��>K���ō���^c�gP[�`�A�U�yb|X޸F�N@��^n^����Ib��H��n�v��m	���{=�Ӆ{���W���S��U��ip򩌰�Y�e�HdNv�p%co!c�g���i�|���j�}j��r�zV", ��FʀE�t�+/I�5DE{Ц'Ё(���wa����ъ1�������T�٭�/�6���-�e#��#k��0nn�W�bnn��wR�n"H�w[�둘i'#a,�y;�-��q$��8�A&\��'����T씓���`+�+b��0ʕ�lXf�V�� u2Dͧڜ��5��vU�e�B�ʷ,�*H˔C߄1(V�V_\�t�����:﹭��vҷr	yo�g/}�jd�frb����~!�ul�<��[���|�Y��w)\���x2k֕1�vmpb����L��P���KJi�X�F4v�� M�xV���� 4pjFb�;|s�Beiǎ�vB��P�6�q�F���֢zz�h���Y��h�ƹ�AΤ�vT��1Ԟ���[�Z��c�K��mW��F���}�N�B}y�n����N�5q.�W ���s�O�L�^�Dj�9���^�Ә���H�c����P8˩�E��EO����L1Q��/��r-Q���[���,���+B��ݾ��.d�+����1�*I��K��d����]8M�۫�Wi࣫R),��j���N�,9�q:���0*-�(�g)Q�K�W:5��n`��BXd���y���ʝK�{�㙮yF3��q���xdE���)��J3hS�)ۋ/�)���,�×mk�W�4���-��L&Qw���4[�r�G5�k��T�#z����۫��}�а�ƍ]��Mv��ի���w�}t�Ѭ�m�״��Sv�.�N��M�;z\��.��ۜz�����n\�\.���r�3Ֆ����:t�*6n$��a�5\���,EQQ����1^�b�=ht�Tmb.zj�=O���ӪCk'IaЩe_+G�ׅ�	��W���:\�]޼I�)�n��ETE�_lڋ���0:���^")}9XJ�#�Z`�z���Nl�oU�g]L��q����q�=�'���P�6ԥ�óT�3�����S��ę�Q0Vc����F]e��5����b|���[�Z����+��X��9>���V�u3ҽg-ӋsR#+q�n�I����
W����x@+�V�;f�=i�U&7�"s��B�+�a�gO1��/u��ß�����?f]�/{�Q���A�	z��Ǩ�+��
7�l'WdOG�(:}����qU�*��t�l�E�eP�P�V�/U�կ+��{��T띡�^�[���n���n��z�[��N�V�Bu(rFڇ~�r����d���5%�]7HĨ$F�����;}�M+���n;��5*�"�5ᨲj,�(��y>�$��U��U��c��#	ІU��o�s~�J:�+CI�n�%ص,�vv�@�h�T_1U�K���=p�%�7=�O�E���ʾ�j���-�`��M��LsrD�Xԕ�h˃Z��u�s�
�����g�L\MX�:�Y����t�箷9�oc�Ɉ�����t*6Gu��x�k9�f�H��LZ9d!�S":�2����|&0�eD���������Z�!9�'X����I���ʭ܇���cn)U~c&BÒL�S{w�]R!J�L@�U��!��Tc�F��^�wr#t�P�;q�1^5�\�:}�Й7���R����j�����x�AV�q}N�d�bct(R�G�^���c�&:-�{�Ͱ��s�ǌ3}r�b��t�}[�e��j4*T�NJ�0�k�x�L�o;���,z�`��3���i�t�vW�ӑ��?c�dY�X:��v����QN�+�:�%݀ŕb��X��q5.;MT(� a�K���:UJ�A��Atru&sw�����(���7$`�z�'դ
bǼv�[\2<u�[iC-�֑�$�oe�[;0���z���p+ܤ3��Rt�uT2�p����R����l+[��͠^��u��-%�a����3{H�jO���5�2۠�ZTF �ސ]�֋��Ѥ�ѥ�Y*U��" <�-�ɗj&w�H̷�-;O&�f�g�ԭ1uX	֒�˙�(Wq�эS��8\���C�5�L��l�A��z��Dk��u�xE��l�V��+Gt��J%�/�;�q=���Փ�6L�y�]z���g���U���`XuW���t盝f�}q"H��*��Z�R�Pm���N������Hzk*��ʌ<��8/Ùd�	�����օ{=�1䄞�r%]?}�U�'�8��$Yn9Q�Y�Yf�_PB,�.H�Su�'z��P�؍8ҥ������R���x\{HVNCe�F���&��|�`'��QY�v�8�C}7<��p��¯T��>ƣ���O�6Z��S���f ��
(͉u]T�t��jR{�n��<��¡YzB1!oP8�=���P���
g�ψ�*�Su��0��'��پ��pܨ4�L�:P0���Y��P|��=\��O�v�Jyڃ�M�#�uk-t�L$C�(B�EJGLW�u�P�K��2��q���ڂ:��P���*��EM+�z���Ԩ��j�Qk���0��_	�W���r�vchڅ�uz�X�g�R)]Xd�}i�FS�j8
����co�Z2��炮gM��_��-'{�1�������v�$�<�oX�Co�ԑ�Y�£������eSh!Z�fV��w]�5U���..�6t�6�؏�(p!v�%j��`:�ףo�:�`T,�9�xa��\�K��D7*�Ck4G.ou+�p��L�.�����d�^�L$aQq.a�q.☸.�^�I�<"�&P�)�i�'ie�u�������H�zl���9�s|X޴n�L����>�!���3.�,��#+3Xr�y�<�6�W��5����X�vL�l�f�D
މ@
JH�o*��L�������'�ܦA����g!�c����ÑWU-\0p���u3ހA����.�%�w^�z�̓��u�^��j����Z�~|P�]E��i
Z:�����Vng�.@+�s��� B��3��~��U4Tk�R�ۑW�oM�̑�Ӟ��^�1c(J��n�6��32���j[ڨ�,"zڦ;��ǢW�ӂ{Ui)����>��U�^�.�Z셖 GN��Y�1ӜB8Ǝq��:zW���ӏp�W���#V��6�a-��،*��gs�9��i�tDU�%1ة��6�
��O(s�o�h2v��b�g��Z�z��>��^o��05r�x�*/V���QjY5�Xf�t�4!^<��j��S��?��܃\��r�`]���E��^���D��ԧhzCu�����D�J�yfR�u���
l}��� Wn�@��R�YFT8� �Zt�iq���n��)��d��0���M�v��z�`��$�P���ݹ]֫���^�����T�Jv[�ް9q���@U�# ����ҷD3�Lx��	\u�fe�,|��d��%=�8(�&��sM�6��[�Z��i�ؠ����e�"#�f�"��j�n���ʉ���aM�ii��Wu2��1'�2VH�Eᡚd̲�m�K5�FX��\��r�+_�ܧ���z�}X���R�(+�8=�۠��9Z��-��aMʾ�Wԓ��j��M̴�$�v���b��d��%�k�
�%8,��W>���8� ��U�}ܧX}���Y�zJu�q��R�n=G��5|�k��EeWi�]Y���Wń�o-�2
��{�2�)0��5�����!�kF�x|Ps. ��߯9�n�@��A���]2���n��YG.i��n�,M�ؕ�U��G�*V��-,���V�V��W4�h�lfAEc\�Q�å�8md���X\�y�[��B��l����ٹZ�L�)8� P��/qn���:��e�v8�e���b��Z��u
�ے�<�!��v�R��mu���FN%6�����m�ɸ�c-��ͣ"��f9�Սy�����a��� r���(2�"�kx/2�`�M�j��ج1�F�\���VÙ�PʇN�p�J�۹��=�!R43�c�L�
�g_-��Ӕ�[MZ
Q��8c�nn�ȕB��܊K�{3|��k��wm�3��q�Ѱ��n����.��-��u��+�ɇ�D&���
;V�m�Wv��ŵtI�3!�m�f�h���B�lZ���z-E9�&/��+!0�4˿L�}��,���Y�3�1T��^��Y�Y}���+�h�⯔עar��u�!,W[�C�[�'��)�uwA*ݝ,�{�Z2a|�a���}��r��y��u
����+��l�Y@mE�|�H��k�)���k�S���|��;�����v���:�.��;�;Cq�
��mKv�i5+��j��_B���M�d`m^b�fB.��&ά����,�um�z��6D;�!\�}�*�/.]���)�.���esZ�%j�Q7o5L13e7�Ȣ�!��hnd����_\,Htz� �͍Ǖ
'��99�����f�P@(��/�^ِ�:��Ɂ�N��r�p���#M�!W!<3{�����Jb_Q��ZloK8[a
y��<h�s�Yng�%M���0G���ڻN��-o��լg
7$��Ιj)�hh�����Jގ��Nz�ܽ��.Hb�=�BL��e�w6�[&��<���I?K+�CB�����t�w0�7��n�u],�c����v/G1���]_@�=zۯ<���}�ɟ�~.52������*�"��E���1$Q��Ub�"��*�EE+UQUEQUUAA`��F"���UF���V*�*�`��(�X�b�EF1�b"*�0QQU"Ȋ��1�"������T��TkF(-J1Q�X����E ��"�"�,UT�UEUF#�EP���F+AEEX���X���YmTX�("�(�
������F (1EH(��EQ��	i*,TA-� "F*��� � �F ��
"
DQ�����F����TdPU�,��
�b���1`��1V�}��;˿�]�n�+5�|vSb��8�i\��+�"��>j���1p��{
ԫ��-��p�Qg]]WN�wݵ���:E-w�4�������:����;Q�*��E����}��j�c�)�͸q5���th�G8Q���<��F��i��O��PB�`�Lvz]vd�s��y�w�ͽ|�Cy֠���,��Ú�u�yFz-�(��!���0P��a�b��ھ�@8n1o*���K:�T�v�pY�yF)��o�u�i����Hh.�B�ܧ�޷�C�Xڸ��`��N
lܔ3a�=Tj4��p!С͛������S��j�9���aq.)N���SY:J`a�b���1{�h![�4��Sk��
R�	��(&���X�OL�A�`TW�x>�j/q�t߆��~�8�J���:�|�i�Ԉ��62Y
�3sݙX�����<yk�jjR���1֏[�%�Z����X�.�O��
���Ǝ-H��.1���a-Q2��"Tφ�J���l�3�8���P����D�[��Q������Ք2�����^
���;g�g�yU^��W��ڂ��R�y5�5m�S�oB�S2����g�5@�"��]V>�q&p��d[Z���;<�x�d�]���,�c��5��!㼸���-��۔�"�HV��r�\�	LV+z���+˱�U�.=r��x�v�k[���J �=pt�DΜm��Zm�����o��̺%�u��׌��$5������YY6mpu���F�QΝM��C���vZ�4�}�M�m(v��aX{ ��[]L˶贺L�I~�\s�b�t�W��8����"�Z�#:�9�P�*w.��m+G;}EMG��z�z~�����-���6
x䎍����hH g��x�[���S���S��V�[��M�0%����{9�q�W���*���u�~�p�i
�Iv�hmȅݹKk��W�;�Ga\\2�������Ru���X��!�.TY�aD�����7�&2�f&�5�]�nU�b�3"�;M�yB��!��Tc�F�����v`Sr�P9d�{E%owW]Sz���E�R��3�T�������\<�i�jwާ\�X�M^� Gr��(�^�t�}�R&��Z=���D�\sgՊ�{bXaF�*
�ؗN%��׭����a�<�@4J� ��3�̕�+j�i�bX�Rt�:0lō<�vb'��۞+]E��8;�Ŧ�;�gJ��W�*:ܷt��%[}�p�ͩG���@�*�֖��ST�Pv\V:���HVÛ���m���zog�L��񭸙�]�>��b� -�u�ݨ�M-Z��C�=��
&�uʊ����\&�C�A��K����Q��nj]�qV����\��ʗ��>�V��u-�mG���s�6��}^W�v�Uxݑ��F�%�I����*
���x�����p��Q���e��r�`mn�UuUW���r�Β�8[���a8\ql���Gi��t�e	X*]��5�;կ�X#���U�8%U��]g0
��N����q�<jg\PW�.�V�Zv[�3R�}0�ǆP�,�+���V·=��������/��t�x8��:�JOjL��k5���pG�oI@~c5J�Q>;K�]
��kG:��p
o^��!��]Sv�sY��x�.�p7 F�7g�� 5�H���u���ӊ��]A�||g�;5��fv)D�� -Kn��v�s�T8[��i
��!�f��>�R`�yj$�q4a57
� ə�TM'�� 6Pl�f�-0�*zr	cQ�΍�u#2��ޯ&5�Ok��\(��듽�跔u��i���1PY'�*��bBޘ�Q/zq�1������=���E	�A8+��k#�Z]��c����!_b2��R�����bp�8y�ە�8�F �]b�KeM��������uD�T�ó/�*������/s��9Z��rt���ܚ�*0��h=��b��PtA���g�r�] e�nEQpgo�*U����G�2��M�@��w(FR�~���PB/��#���]���aBƬ�:��sW�i�<ɀ��P��&T]u.\�7�����Z����A<c���˲mȏk�%:+.�6s ��H�HY�ى���hU�k�|�^��"��[�����L1][O�R���%�i6t���V��#�Uښ�'�/w��e,���M�WF�gS��T�)
��vL^��!�d�7č%�碘�fw}��Hۥ��l�f��^�gf+:v\߸���S���ܽ7�wp�\�X��N���\��Ac����Hz�Kv�3�J��8Av|��S�\
8m. :�D_�������hk��&d��pN�G��.�M�XH���j����7���wϝ:E=ctȧ�6
�wh��gH�!-�!��Q�P�!�V�e���(R��VR�[ǜo)��ެXE�糨��q7��8�:�+\�!m�H��Lf���#7U�>�d��(�'XY�eߩ6���R�6�9�G[c^�%2=�EL��	��h߭��n��X���
��/�Z�GYЧnv��ZՖ6	ӬK�u%�8��W��2iڕʄD@]��1+�fR��ֻ��d�F�&rDb�5;�1=hr��)���R�)�6L&�W�=
����5iS�^N�f���L���/+x�*���K4Ft�MR��;CۚdZ���؎SQ����=�ڜ��s���vU�d �[Ʉ\����V�w;�\T�	����d����!ҞP�>V�֙;s�b��S�\鋽yϘS�#�#X>�=q.j���,��R�7�èS��o��j��{w�u���0Iݧຜs�Vd8�%F�P8˩dٻ*�g|1S���-�)�Uk�vv�+g��=t7�'�Y�F��)����2�`�Lqs�w[�C�=se>W�'lT]���eY��ӧ޷���d7}F��F�^Q�V�E�!���
�С�ou'��9��.�q�1\�t,��(;[��f���[��Kx,-f�F��aL�9B6tc�W�n��v����X)F ):M�A�J��m�:�^(j�c)���A��uy7�(�,m�I���"n"���2�o�t�*�3�S�]��3_�1��m'�m��{q��fhG\��xUb��+�:{c���qe��ԙ��1Z���`t��c��'��vf�Y��Ԧ������������fԈ�{����K#�"�$��P2�����*BFr���2��w&q�x.�V�k�'P�)�7 T��2�o�RҒ�!���������;����h�̱�e�1�H�F��FRMO>vWu�<��Ngr��p���_�QNlPb��נ�6�^^�������e�ȠM�&��靶�ܓ��4(7���C�VF�חr.���v;*�ּ�,��Lks����f�S��ε����}�T�^
����r�=i��T����$J׬�-{�泈������?*Վu�GSp ��{�Bt��}Y�f��pn�:�bj��fuM�	
�#9F��Y�0�^l�F�s"�5P�ŽT�J���ȪOT���Ƌ��˲hjK.48|gE��spVW���@���JqA���E�a���E��j�]��j��ז�v3�6
x��;�P�}V+ڋ',�(��VZn�Q�/����ID��~��N�α>:ݨ�-��:,�ns�-C$����M��}F��a.aV�G#�o#oe����u��;X��-�pUj�ӆ�����${K
����cW&�5ʅ�gm���@߷ހ��=�7�Xo�
�k-�I��qWk;&r�(�f����Χ�d�aT���{[;�
����,�Quճ١�,;N:]+j���ȱ3{׏r��v
]҂bf8˄��s� ٭Z��ᮕP�aQ����V
^XJ��Q�����{�2!�w�ȑͶ/e'(M��[�:!�*����E��%��g�×T�?���P�S ӭ�Yn8'����3�:�lr���fú}+
q��JeŞ������z�z�~p�8�Y�s��a������D�0Oy)��^�ݮcW�=g�a��;w^Xӝ��&����|�{{���|��1����z@<0����^�!��U�,���s\�ON�/
�=����9.�uU~�^��b�P���ňf����I���������pM��9ַ���)�r�Q��K!�J�+�ԫ���We}�������e5�0�S��O�����>�0�ee ��nՋ�Ky��c�?����r:Mf.�rX��7E=JglS����!�`������gD�&:�:�0,;�;"%t f��n���K�v5�q	b�p|�x�-�gQ$�Σ��yv�}~=P��A��t���q�nݣ��{U��F�M��}~�L�5�n���Ic�0��VUwr�4;�g6�v�S37گ��/�i�,���C�/����O�9dK�2� ���F���;Vĕs��16�|z�{���P��ն��%��](r���C����wCk��[*e�����7��8��Ab�,��P�X�J�T��� �[�:�xe:�*���y�e>�3	U!pu�Ӟe��c�~Uw��u#{Ϩ#b��@�R���v'k&jw1����: qgG n0�4�Q�^���W�gFߡ]B�����yB�K5������n{ݕ��u�@o���ʺ̳Ü�J�vjb�����D�*/���2�mF�֏H���%@p�R=�.i�ʛ���K�f�:P0���X9{
�DJ������*���8������@�z��e�P+ǥ#�10�����d2��K#z�5yU�.�/�2�d4W��s �n�Qk��+��o�baa�/+���1�j����k�#�1 �J��ZOX�
ن�7*[6��>z��gI���V��\.��%�7�i����`ul�����T���v��T�)�{=L�pD�s3b9�IU�Å�	��:KY������z)�&P����;1����j�nش���=�)�Ct���TVNP�9�n�G�~� ذaK�v�&|ld��{\�U#gQ���xN�6�)��YS!���j�.��`�$�wg<���3�N�ʙE;��.��z���Ej^dCy��K]K8D@�v���-Q�Y��X!8b������;�ċ�$���	0x�-����)T.�.σ�X�u��Tp> :ͥ�\�n���YZ��#>ʸ��p���Q*���.�߅�"�Z�eb�3��hڐ��νٖ�A�y��6���'��
zt����Ɛ=\%�Bƫ7�H�޷T�-M)c[�{6v��SmGAF.
��%��c����c\�!�e�A��1��I���|,[�����0�q�j�v��[W-]:�R�<5�v��("j"Ҧ;��ͮ�f���L��%�&�C4ҟr���j�c��G�;'���D_N� �<{��e��o�z���n�~z6��s����@~�n�Z�a��h���3&�O�Ţ^ҁC��C�<����qu,i��x��o��	��xtba�� �*N�>�1*j���R��Xg�)��h@��W7W��bM<��9�9�OUs�3�N�u�q�/R�[���)��O-'c��hh����9��ό��r�]�mF�Ar����n5��+9���^S%Q�PB����>P�6nF���}�RUW����A<��j���13�򮌭ę�݃s3�Q�����u�É]�ƶ9�j�������T�f+�2ے��/,[�[��LLv�sŮ]j�W�k��3dI]�i�ػ�	29}E����6�ʄn�+�I�@H���X�ަ.�p�nx++\N�����n�  �Ú��A����r�9��Bw	�Fɯ�f�IP�����s�1��q�Ƞ���gz"�f�\�����e����o�[=g}s 9�N���y�q%���ACU�NX�8/_d�lPs�K��nzbb�넚u7��+ǅ�S~����pв��V��xL���8�?)�Xg��sLs79,���8�r��!pU�QP��Zs�k�v]7��/��K���Ho����qw��jȭ�������6l�?4����f�ZFE���;5e3��q�\@�V*�孙��wk�n��l��1�0gݮ�F�Z�0lk˹ºW��̲p��a;�G��T��z����-F�u�c+tӌ��5�B� ��^|��C7m�zٜ�^Z����b����I�}2��䵵E�A�)�Y
�T`��B��vy:JN8�J�6���Z1H�gb�Wsكo�u��g#h��z��6�� m(v����^�]_
�7��^k����@#5Otx��/�/���|n����i�EӮ<�*�����1ycHa�舠����ѝ�7iw����JX�i��q�2����vA	�e2��)� $.����7!sL��zנ�S�l�$�`AGk���1 2v��󃞱0�$�2؇�*��b��Mlq�Io-[�-��^�����,���S��v����)�L[�a�/,M�ݴ,��*�J�]�gS�� �=c�E��H.�C�bN�%���kJ5j0��sV��]�-�j�;�7��sK�.b��,�|��:Ɯ2d��i����w�����#�aR�����%�m<���ΰkζ���m۫wy3GYwu��ԝtg	4��B�U�3]��o�r��޾�eҥ��Sw)�.-�z; ��*����#z9�of�y���\_mo��[����u:����#��Yn�����Ī�do��� |A��y2ڠE�Iv�|�ٛ�g�V׸�5�&��j�_ك["�������ӊ�����X�����+�2��;A;w7O9G�v�Sf��[m��:�Z��@�'S�ʌ�d-GS��.a�4�3h.�t�ӡ4Y;@.����v]�a��f�l�q�Beʚ{]At�C��I��]ݩ��t ���J����C�����t��4C��UX�[WV9��N�ʓAЏi6/tI���㴥�bPc㊴����5�(�ᗌ	K��;��� +oPJD�Y絽�d�r�;̤�yl�� w��Ō�5ӬVuYZ���r���=t`.�]3+�'2!��0�x���E��:�X���J'3�U
��Bs�J[���pG6�ȕ��� ���G����kb���l L.��N�䑔z�L�OZ#����x�UJ�np�g	�P���]YGgFT���4eb�{wf+�8�u���h�^s%�X�\u���LQ��ҳm�����������ڗ� 'nͪP���n��a�}�}�mep����5sBwZ\[�acr�V��[��8��+(���v�x[�)�wۇ�
��Kg�u�-��ky����v���4�wX�d�(��cle-[�uZ��L�
U�ɞ�y�3Ir3|`���I�[�,K�:�k�X�Ho�2�o
����<j�?OM|��LṴ8eu.(Tљ�*+�)>�����L�u��5;��C2_M�5:���f�'sVAe� -�,IT�췴=�5��X72Sn#�"|_v����:j\��w���ܽ�Ν�`��2ZWB�Ԯ�bkC7�8',���x�Y��e�b��띡Wb�?���D��"
Lj4�Iօc�]�w��:w��� )��>�b��y]�k��g'�v8/���q�i�T�U�|� ;�Nl�aM"=�Pʴ��rX��K��K���S�@�Mճs�."��y.�^�������>�"�p�o*�ae`ِ^��fV���ˍ��FDX,Fm�U�����*EF(�**����b�+1QEAPX����EAAX��"��J�U���DU����""�*�*�����D�`�����UA�������"5(��1cU�����E��1PQU�B��X*��V*,D�EX�PcEQ����E��X��(��TDTEUU�TDV,QE�DPAA�TTV(���b�R1�V
*��(�cZ �������DUQb����""����`�bV�bb�b������R�Pb�%�-
��*�QX�*QV0D""�4 �� �P�
�c4�z�36�V�l�l�F��B�"\��|SPuco��KW���2��ݾ}5d�u�U����{t 4"u�)�8��}�lsf��Y.E]�Y��1��_���V�ѝt�gQ���f���\��)�ڈg5�����+$�����]�����àuMAJ��MD���Y*l�6�Tڙq��"���KiEä87��	N��k���q�s��!�f�pv��A,��-�m���#�Ij_�}�b9���G"���E��!3Ȩ��@:�dqo�6F�����f祛ɢ޷�v;%��q���"*������P���|��G#Z�������K�K=QzVku�R!�ҙBT��`)���E��(aS�w"ePsL!J�<��)�Oimeҍ[�mul�gu{@�I
�nKG�bXڋ�K�p�s��W	����K�^��=��}Æ���X�?R� ���*��3�ϛ]�U�]/^z��`b�S,�m�GӯN��Ȭ8'��p*P��*Ì,1���b�=!��V�(�mŌ�����N�5���w"j�w%tP���W���V����P.9Hg��#Eu,YYD�@����8���S}��z�W�
��Vf]�Y{QS��NT9��Z�i]u�V2��� �K0\8Pz�����e1٦��&W'Ei�	�^Q�?_p��Z��l6�4|�Y\n4nj�(t�t��\S(	;Mμ�l �v�ֆ'/��3��Z�q����������n�窫�^]a��0�&u����&��3�Ԝ�1e�M_.n��xbl�a},׃�v�8K�p_cU f��*9�=��u��w{gx����1�$3kdZ��_U�/��_IB�d�oj��������O8�6��js�M��]��U;�^��L{oK��!x�5x�R|>_;o�Jl�C�k��a^��}��9&Á��m�b3���n��tsX��[����s1i��C�n*{۽<���}�G!����q>�gܪ������Pan<.=�+' ����
LD�������� ��62��59��p���(C�@�a�j�
�*zr	cQ���B�g�_�����|��$�Y����T\�H�S[ۅ~�1
{�ܠe.Uow*�yI�xVw>��Kf�
f*�����;*n��r���(FaAu�hC&c;K��v�,��x9�7���(?bU�b3�k̘�E�RS�B��]R�@�K$�t�,���ʞGFn���둍�1g��⻢i_���S��@�y�VQѾq�I��d��p�:�M\Y����d�'�؋�� �;�E�����);qPW��E�k��Bhۋ6�x�v޵N��
�+d-AR�V�𬼣�؅
��7^v�ӮI��{��V��S�G2 !6�P�HY��!��A;b6�pœ�#H�bz�b�cv�1J���-�
"^E!~�����U!%�����*�Y����MPX�`ӝ���Cީrp���e��a��)�n�nfb/ �ޚ�~�&̢T��z�0�'��8�e�GX4�hX�[N�K����9�#Cr��w��^�x,��[2��kS�9	ǃ�I�>=K����U7T.�.σ�X�b�Q������� {w�T��*F��7Gn�0,��-5���
���@�Д3r��비/���by`*`�StE[������ ��{�����\���H�-li*��>�Q7=V�e�%A����|��l`�8�8&�PΛ�!+�]���-�K�c#F���]��>�1��y"3u/=	+��"4��f�72�A���(65݌9Hq3�xf�ǣ�鱕�U��P��y�M�59��r��w)q�(m)�E�:t0F
�MF\.v��ЙZr:��z�x9��=.�>k X���a��uH�ʽ�A	dlN�D=��Z2E���a5̙������e��c��
CwV�\sSF�[�ž�r�M�L$�|�Bt�R������f�����!T�]���]��y;Y�W�� 6�)"�v������z&�ц5H;y7��4v��=e$fM@�WKf#�2�ҁ\��1ԞЭ&:�畢��$�$��-��:����� �QSz3����ʚ��5�"�^�,3q�ù r �/v��޽J���_+cT�+�8炬�qj���U(d,�n�\J�&G\Q���
�P�����ev�0����r7�'�\�Ek�bP>'�uZW�h��*�0�n֗����7��ַ>����LF�?�t��;����_@���d��+T��.D_�w<.^-��=Y�ӞF�n��y���p�V�:�0�k�������l[��c�d���F�I�uR)�����U���7N���� .��' �gjTf�ð%F�N��ދ�'9^�� ���!������Y&/��OU:Ck!�u��'������}(ׅ��e_��ڄ�n�EZ�燇��\E��ڕT! �	��OaQ7-��0o����͒A>��x*�;Uu�n�<v*�v���Dr�zE��#jؠ��R,Î#�v\���h�����L��#�D�I�L�J���0>���Eꗒ�\��\EUf:�Xc�5Ϧ�C�`M���y��P�"�<�g�Ub��s�͙<0�@�Zu�u�՗Ύ�^"�!åd4 x��FЊ�/��{ǩ�<*\Zڔ�ve��o3o��9gI��~;��O�gF1Bh�X��q�E{�Vz�BW������!ɣte (޵}�1������=����+9�QtD뉃Z�����s�a�P�:�hM���7�OR<����\�76��:^��N#�2c���\Fի��
�鏺�k�A`�u�<�*�ʼ�\�rp��LX&�=E��6+���7��:���eI��6v��'��Vis4�:�d0ڶ���tw`Opt��[-���a4�TY��%^�,���J����xy��];S��S��SV�{^[����$vN�u�%A@ڱC;�{QtJn���N��%��f�))>�Jv�u������p]j79ۂ�T�wL���0m��udp4SԤ�!��2#IH��ea�)��ń�#�'� v�Y[��m��z4�v�!4�7�+*�Ci�S�T�H�w���E�U�+
����6�Q�G#]�pR\O���N�W��2dG9s(GN�t�𼨹�O��P:<���x^�}s�R�v���tX�1̼Z�����GU�x{��=��ڵ��)^�v"*��B����k"U��%����JK����)=��-�򣛕h�Q��P�}W]���8��G{S�(d�
�o1g_!pV���Է�Z��@�'i�?){�w�
m�WoN*r4}T�,��pB�uRBx��R�옖6�.Q,U��ϫh�d������7܀�������ةR�lJ���6 �����6�N;���.��x(�%�ԛW+�\M��s'�����,Xؒ�sA�Ar��b�U�"��#��MK��vD��gnxv8��t�g�5��=V1�ڪ����HG)�:w1�L��e_�y.�;�4�X6I��k"C���ܝ�t�l�"2�]����������-�R����V�OnMJ��T�'��pڡ>�0�Qxp�i��X�`1��qz��j'ٺgs�M�v=^�7�C[�-1��^}Jň��[:�����c�lLo1dC�Z���)Y��|�tEC^�1��̝n�8������"�w�"�^,��|��}C��~� �xFK�]�{ydL���R��̲jڦ#r�Ӑ����y#zQs�zfs�����g:�U�Z�f�4�3�.H�s����og���i
��!�f���v����~8�بq��Y�GBmY�;�ɒ`p7]1T�oJU�2��!����݂oQ�9�ǖi�����bpų$���偁K��t6�Fx^>�w'k��c�Kr1,�%��V�珿�����I
�A���橚	,k{�%���Aܦ�=],^�� ps=i�C�=9��X�a��:�uV���7\��aL`jj���XNL��������+6K���"Bޠ���Yn�`�E�d����;{���Ն+�f*��̱�*n��N�#/ђ��ǎ��c�����,��*Tl1Ǔ���rTu�F��f#Yb
=)0a]OIAz\�0�^�*���5lX�++��х�[�^m(�u)�#���LE��� �a�+/���0-�/k��{�>��Q�7�b˖3��;L1���ȊT��]ġ�� M'G�iy�O+���eM*q�������Z=y]������e(*�`J�2�[��eا�Fv����L��ֱ͗Z4���؀���ol��T�uE����N��/)U��7�~�@VP�o�x�u%���{=��N6�+"$�Ga�>1��R��vxJ�v|U��S���������2 ׯ;���(( 㔑��U����yD�3�.��~H�����_���P���p��)��^ɂ�x�,���i��B��y�}�v%or��P�uF��:�R�, ���DYq3I�w�l�mv�^E������Y�h����y}��ǭ���t�Z�<P��0�op����f�a�#�5o&Z��DŴ��V^�~j��zt���2��B�΢%�B��V�fu\��[���d�/W:����jt����TɸŔ�1c3����ۑW�7���ލ��RD��q���}L\�� �*��_��Sc]��2�)���n���z'�3N	׷�wy�	<�OG-u(\��g=R��R�dq���<q���v��	��7*zj�ٹ�y�v��J��0��@�!�2ee$g"��Mt�@�['\��V[�����ύ�B�,�M�k�_A�5o�lq�Q�P��o �϶�ʚ6��
�M{�ɖ\Kq�TC�S�DݭIE`�c�y���Q/T�s�9�՘aF�gڗ
�|�vҭ5�Y�ݠj�$z���H�vuƞ��1�>��Ւ�}�j�:勸/)��-�&x��`�g)-H�G E�U�߉\^e��L:���n�,9�q:���0*q��H���3���,�?�70xD�	�F5�X�Qٵ�*�ok�Q��C����H�Q�>o��/����{L�u�n�����9��9�C�{f3ke�xs������cE�ZU�(��⭐�:xG�����:�ZV�;�f��;{��m���G�r��F����9U��u4�(�Q
RZeM�|�E��d�7mhM';&Q�ﻑ+֝���HnzbX�0ʝ' �gjTf�A�hQJ�ښ��̝��MY���?S�"����$��J&e��T��N���s�WGŀ��[=.�5Tg��1!(2q�\B0�l��YVE>b��E��2�{LBGX�����z�����qe�����G(��5$f�9�A���Y�~#�K,,ٰ!���JA\Emv4����nиûs���j�v�_��Ɩ���.�_����'w��}D�&�7�;#'m]��h���k�cg=i�u�Ք2���gI��F�[��%�����N�U,����9t�s-`|D�c�y!{)��
�q��Ftj�p{UURM�=[��X�R�dk��!h��~��$�K���*�{�L\=D��U,Vh���t���v�#���<���	��#�Ml�h�Y~�"����}B�s:Sq�� �m^o^�8�yTŇ��==�)���24_��n; ��=θVv��)a����=1�̊�՞�V��vz�NI��]�12Iz�M5���GJF�[��$��]�)#a��K֒��I��#��-�\c߳i�E5���5�0�
���)��[w�,���I���V��#ئY�崸���4���P���:��,�����RW��b�S��5��:۷�٧j7P�q���5��x�M�z�mp�.$�Cd��+����xR5oi��L�7�'���k���Z}�I��'�jsԶTQ�cӆ�U8�i�ҩ*�i�徵t+�;�]����ęN&d�Mݦ�w8ᕔފ�d�ܲT\��1,m�%�xE�*zΒ���x�q��<�xQOy�~{^��|���; ZQ]3����8��2���ݔ���R���C���rsN>NXS�LY�j	�����*��:mv�v�v�����Vmv�<�L�f�u�0>�(�F�Ѣ��cnJ�MXc�%݀�T$��X��\0�P޼���<2z瞷�hvܱr�la��s�~�Cj������v�r��E�tF���'�`��>�s�%�kYӤ�~ E���#�w*Xڂt�r�]s�U�D����C���#��^Ue#��P�&=��5V��i!ϼ��Y�����>����`8�"P���+���[�Iyp̮��.-�Y����e3�M*�G�46�:;��d\����֑�����u[7ؤ���frnuS�QT��ȪTl��K`��9O��!WR$�ϣ���Z�,�pup�A˻܊˼�I�g#(���u���S(p�_oյ���G�AX���d ��TSy�Q8�7�:��[��9t�j1Vw��UG2(��0���,ejKk 3x ڮ_`-�V�ԣ(�]����;t�Zn�6�l��.V�ѵ�����we��!��*��x"�X�x�ե���ʑ��t:6���U�B'u�_����K�t��t��̾��V���f)lx�=�
Ov���ET+$�9p���A�!��|��$FQXq\�Gu\��w1_L]��I{D���ݒ܁����(�̑)g��͋����� �	�g|D�$2�S��Y���1��Z3��ƞKD6�Ø�`�~Z�`����u�g�Q�9S�/!�Cs��&�m�Zh�N�ܺ���je.V*�����bZ��G�)`l�% si��y!���7M%&���Y{%��.F`�;Æ� ����ر���ɨB�����F�E�eQ��e͎.�}�9�-���/nnɘ����zd���oUTd>�_ƨ�3�W1��\U��y�]F<�V23E)��8�).�(K��m��01[]��l�6{#���\���;ȍ��\8�9X�QU#��PCT2Ʃ�)6�2�w�,�m���{r���4�7m���[�s8���`��PvY%W7�3��B��ܴ��+p���v5�(�2.����T�,����FpKȶ���U-�p~¹wvЯV�L�N�m�6����@5dv�]L��t�tfnك�Č
:�N�0���h���`����x��pd���0���4�N�s��o��֌v�!B�`�6��X��Rֻ��&^2���X����	�/���}����S���(���ioNyB�N��j
�Z��踌C:��Zm��J�y'����ʳ#}X�mH�n�n���jN��6��2؍vm'��J�K���A�Z���ZDEt�~�*�*ohJ9��mA�q؛8�M�*R����j35]���hZ��IPga�Dμ�]r��_2vu�8�v���9K�Y�[��l����Z�T���һk]�2�G�7�vrB�����3;6=|`�{ab7��z�d���-�a%Rz���|��׺S�ʕ�Ύ���;AA0��M�w�E£�����f��t��)��hNyҵؠ���r���6@�M<B>�t1o�93`�4� �m�YZ��p��{t��q�0#*�㒵^�IYK�V�,\�P,����M�y�uqr��R ,]e��m�֮��nwl�r����Z�V*�Ɋ�{;������n��V�z�֗�|�߻�.0U`���(�",X���� &����#mEX���1R��V"�(�$Q`�DDDb)-,EB��Ԫ1*�)mm�eL5X�Z�����Q��X��Q��؋P��Kj����U����UamU��UT�AZ�TD,�E����iU-,Ũ)0�²(���ETTPih��YDP�p�%�X����A�e�UV5(��++-h�c���QT0fTkb1`�EFJ �VXVc[KJ��"����FF"��EE�e���ƥV0X%�X��E0���V�TYR���bZT�+[+AQ�sHT��	3i��M��/y^.~�i�Yo �AC��jf��Z�����t[�.�j[CE�&�ؘi�L!3s�u���b�wu�����S�A�衭?W���b�x]R�bR<#�V·=���_���d��&�o�K���#��b2/٩��ycvq����`�/���!��`ٌ�2��3���V����s�����=|vO].��&��b7�m��=��<6�y��� �N�ߔ�Vt!8sGNF�ShP���,�.H�r3���t��A���b���f���XT2���k�Q�7p������t�t��	�y�L*�ʞ�|%�G&�N$1�x:�5;|�էp��
�5JN�p���sLvE] ��EF*'!B�^��������x�䎎�A�)�V����q~UAL�2��
un;ѹPiҙ�1ҁ�uj521m��lY���re�PB/��#��rwk�"*b
=)ɉ��=%o���؂7��Ψڗ.�,ͷ�y����l^z)�#�X	�b���@� �3}n�z���eh�V���!k��.����a��1^U���R���y���3�).�(kN0��6d]�p���@�:�ƚ[|�:+��}J�1i��Dn݋�,6�_^�#�(�pV�6�T�se�}Ch(�
7iqv�uw^�m��sWZ\%��J���u ��q��s�!U��c�
��
��:$��!�
.�*%jZ��:��X��D�i�K{.vg�p2���.(<񮝫�P��)��>���#,e��٦��ǜչꌫٮ6����j�Y%��F�����S��X�|mV_,�G����\M�y���9����{P"�}�}+IUUB�$�. ����8ek|*g�H|2�b*���⺕M�}q�����f�
�FlO +�I��Cв�yD�.AB�}T�
��CC4��޴�����1�Z�c�b�:و"��$5s��"൱�0�Ox�f��5�l��k*^cK��2僔1��b��s'[������C�켈<՞9�h���U�V�5����2B�]eS�D(����k]Te�J��J��:�k�k��� �"�ނ2��C\S��>ż	,m)�E�N� �<r���.v�ܴ5R�����	.p~=iǪ�{e�].`�0h����>=o��]z�����>�»Рo&v%���O"h_P��J�tk�\��yr�δA��� �8�^?k;>\�v$�hϧ/}�z8}x��n�ۘ��;hW8��W�����A(�NJ�8�t������Z� �u�Y[z[[iY�$�X�N��F��D�Ό�\����S,T�6wY�@9��}9�E��`o��r��>涮����Z3uX�� �ܮ�cǈޚeg�tJhҍͽ�e 9B'{���+B?:AS�ЅA��T�*9��"j�1^Sh��(GYrai�蓼�rq�K&���˩�s���r����_l���r7�'�Y�t����,�F�ɖ�g1ʷ���a\��c�wW]f���e�����F�b����]<"��F�Z�T�p���P�����S%.W�r!�(��CI��O�Ƽ��(vl���l\;�y6%�8�I���L)wzo61��Y,5���nDh)�>~|2�R��E@rk	��p��#���4������SԳ�s�M(�Z���ӭ��$�M�|Loφ;��v��b��"RP����)%g�Jf8gQC���O����5͊�9������M�G�"��`[�:{����6�o�>�"&����A��A@Q�%�QN`c�B���m�n;�d�Ի��/'�S��-{�Y��8�> ?�VP��v�\#a�7Y+���F��|$,(��kE9��ʲ�@m�g������t�����P��E���fp$�kh�`Ľ�8:�d�`�|���O$mz�f݌��Y��<�~۬a��u+XwZ�H��*�Dl�&�4�d�{+ºfOn�:Nfc��[;R��-�#���)�w���3��x�h�G����I��S��������|�M땅u������4�%\�9:q�+�WEّ�cOeRc�`�2��|ic��h��ˣ�u����li�B�X�;��0�{�9�!����}SpV�����S\B���v��h"y\%j̵pN4�ۄ����$v5muk�ؓ��;���<�p�[�+j�u�Y����2�U^wpG�z�R�;(>�N���v2
j��k�p�9�`�<rF�R��#㵕�e�r���^N�*�c�G��b�>�.
t����:۶5�3��*���#��L�D��j�H�䩋G$�Cd��+����~��"�RF�]5�O4�1�]\QQ��n`�Nf��&�1�
�6SN�T�O�]�"�q�
y��B��e1D9O���^��3��g7�(��Lֱ>���L�n\��S���N6��}>KE@�-�+شH�ew.[��L���М���c����啎r�v���:�Z=��ע���=�v����2�#[�/����	�LS�ņ�p}K�G ��{��3��i���uw���}�m1���n�q:wM�Hv配+�\�Y�!��Y�*�DĎ� ��`x\��1�=��[d,S.����p��p�g�&e���ڽ����ZD� �7�Z���UZ.G[(�n�'���4ﲲ$x�ģC Z�t'-��j��qU�}[�ps��u��`�O�\�c{���bʱDIe�W�w�	��{�7IUf��/�u��k��>^�i'Y��:��P�������hk��5��j�v�s��K�؉7ꡨ
���a�J6�:B#+u�:몪�Е���Diŝx�Zj{����遍��F%P�&ϫH}�/�ϕp�ׇ�Ǧ�˱�~�w��l�Gv���w���Jtz��9Ԟ4�:⭽����P3M��IB�d�e��ؤh;Ou�E�Ajy�WU��9\FE�g6f1�����ł�ޒ-����D�����W/��#]��t�>�V[~�D�b�WC��s�@�r�KT�gy�ݜoo���ŝ�pBdV��B8��ՑwX�rJ�u9����f��E��.O�܌�*�,맧A������ݴ�Y5H�N�.�J��~K��]p������;�&+��,pH�<��T��{���0�i����K�^��^m�#���]B�5JN��Q.i�Ȋ�Yh�h²����B 7QӖ7Dܛ� \ݐ�k۳�Ŕ��Q4;v\�!�)W%���G!������q飜�A��R�D5���j��dk^�w�#�/��ն�I�}%��.��D
��fӺ���Ѯ�
����>���{q�2��͠�ݯ��M�5:�Cw��:��`�ut�eyug��=�yҫ�\�q=BV��t���I����$��YBǒ^^J�ve��Z��;���R�~5��'Ȅ!�䨍u���k���L�eeE������/����0�˳pvXy�Lz�eW��[u�� 8*����������Y��ٹ��ǭg���QAX=of#��@�P��0�f�Ky������Q�i5jA��&⪘���S"�gj����T����XJ�2�VѪ<���_�~7����ʘ?<yҥ��
��4����r�.�ՍT׍��8��O�{QmkB����f*�֤�S��Od�D��в�d[B�I�K������:�Z�X���`���$:��M����e�@����"��2�ʸx:ٳ^����W��x���2���ʽ�����r�ZTr8>��7c%�"}�݁
��w�Q>{u*!�p�H���ͅ�������f]½Y��P�1�\_�c��A��L�W,i�u4:�-^-��0;��a����7VZ�K趆V�}S-��\2X���Vwqr��!tA5b
�"2��ށ���*��e�5��޳8t��`�e_3Qe_^ ��e�]������n�hs�P��Y�	;�����Wj�S$�~�W�_/{��`�"�g p���wc�P�l�ct��l�:i�VWCĖ�f���Ui)����<��H�ߞ��i��P`J9MFa[��;oX��rj�Z��X\+Ny��ۈ痡�#���7e o3j��p�t�w�b;:�yr��ܢJ\�W��0l�hjj�:�A����ǁv�>�!����M]:u��{�t�^ʢn��.k���\FR�LhB��1
yՀ'N9�5QRA�@�	��uP���{�N�[/�nƙT��½�A
���-��F��'�\k�j�-��e���������fD��r �����c���]��\^�҅fʍE�@����ʁ5��'x�,�m�B���
�n�"�-&<aq�w5�P���(:�[�>VWn`��*�i�|���h���d��XZ�ȍT&�-��1,e\�
������Om�FF��z�TB;�o���ᎼΌ�U2�P��k����Y�6�&[�~�����Ҽ���{��s���+�m!:��D;�sa��*�$b;�`@�:ܧ����N��p`? ��1���M��bM�q� ��)ID���oD}BдYup	I�oZЇv�7�H�Ze�������kֻ��v$�u!�u���9K=����\�L/�e�b��&���DZ�CO/�]`:��-������AD���r�ǫc�������")}<�$��1QƂ�\�^�p����,�ɗ��)η����R/%�N�ޝ���:E�g1��^���(M�X��N�H�{N\R�Q:��5�k}39!���b����p�U��m�\icg(����]YC5C�:����'5���W��ܐ�>0*ܙ�݌�s�*�����q.�Kpl���`�����햧��t��t�%VlH�={���%$B=A�E���X)��61%�\Lu"�� ����fC�Y;H��GSuC.�b-�md��;�{�T�W[�-�#��ý4d����������Ч+���<�]F��1Υ��W��j7H0:^t��⎺2k5jK@[#p�
�b|5M�E�c{'���ON�>�n����t���5�=y��X�j��e�LZ9�2ۊ�t�J�js+�Hռt���>��d�(��!m��}L����=b�B7� �Ʊ`�ːE�z%�5ч���!6�\�ם���w�<YA�h�o!pF*�eGc�Q՜�>Y�w\�I��x����d�͎��o��́N�$��4a��A��	�I��ru�*��:����_���D̡��B&8E#���
o*ت��Y*���V4�V1�q�N�9��W���L�n\��U(�B���*����H�p�(l�b�YM<��LK��$䎋㼰u��s�^.��+ft;���H:n������f�M;Y����#�^��s��2��a��`v��Rۣ��p;���P'd\:��rNRko�={پ�SN?7]���'b�4Y,X�(Ws�3ņ:�.�1��������K�/�[qK��,5��.6��C��/�z6� ���2�7u��9=�o �1���>�(ׅ�Vc�bٚ.�k;o�R�؋�ƕf���=��(6m��{6>Ce�]�'#���Y�y:_�F˾��""oj��WF�Zv���\\ Nͽ��E��xB��<|�R!W���yŔ^�s_�[�4�;�ͻ�Ll5�>�6Xv����D���^�Qs�!����ܠ�ê��MV�{��
[�.�'Qw�90�0��ְf���V�ٸj���9�Vr/�ܵ;�Jh3�����aSݙ��)�?F�gYc�a�T���sl\��K��[]FK�B�%[�s'.ͭ`We^_�8�Ś��(�R}���{�������|�@�y��__�W��亁:б��^r�ʩkxCi���y�5xC�F�/{�o�^Ҷq��T���]bEkvy(��^�ty:����k�v[�o8���TV�6�lVؕ]�U���y���G��3��u$��s|���{؃;�^sv�R�t��]dL��Fײ_�?4�r�3ff�J������^I��%�.�m�#�ޝ��k:DT��˃L��1r��q�3*���'՚���շ�[
�@�>�;�Dr����gU�\�����k�u�ˍ��<�n7��tw��3xuF��qք|��V�F�K��ʷ
�c13��X�)�l�I�[���Y��o�K�M�	��p�/����ئ2maq�Y�G��A�w��b����&�'P����W_p��ˍ����N��/?+ԳR�u#\�KS�t�oW.��j����:��S�w���d�u��Ega�&3��e���Z]L9ո��}���o#�"f����7E�f'](n�˥&�\y��/Xu{{+�&��R�-�&�u�aT|	�ɑU�^�͢67�ư��)t�!�BsJ�-,��f�8�eu>��%`Ŕuu\���s��&n_Zv&��k�DPǱwQ�����f(��m����lї��l\�X�aY��_AB ���R�����ζ�i�I^���Q�F�N�s�p��"L�`���ỡ��u6�J���B���Snj]��[ǰ�7��Y���b-�t��(��eZT�b�T�}D���uX��W-��� ��b˥0S�w�lN��P��\2�V����t��t�>�t�z�����f�5@v�+�����M˲`��S�NW(�qS�nYq�� 4�f�䬲b[:�����	|���h�w!<N�*�%�U�Y��Ԭ�
=a^<v�l<�y:�yj��D�i`�&�U�w6k�J��kzS�}n�:+ �Z��h���O���rS�b��&�ڙ�N��Ϫ'�L�+�f�l�Qp��l9{�b����P��86��zr3����Ώ*&x�0�y簑ם��O�b��B��G�˅�KKF�CoF�����yQn��d�&̥�+�T��
�­n�}��"ؼK;�f�om���pk�w��5������r�R�tU_����Mw�fw˶)X���� �;�f�ͧ�^��Lc��0k� ��k�9i����K*an�7Qvt�v�`���U������8U��\�K�C��t��ĵ�������0Мe�KO�VjK{F�uQ��\�����G$�e̩sxҰ��@�AM=j�9�sv��\�t�e<�V�(nJ�n�L�n@k���8.��9kF��iSW9���{
�1�W=��ւ��gT�qWt63L\Փ0��e����v�Ը����]�x�]N�c��53K�h�Ue��{CtA38W^��bNiV���U��Ǽ���D
7k�&qu�32�r��1=�w)�0�U�#�|:��BU��5���3*`fJ0m�c*��s�s�#+N�d�HK{}� v]�K`C+��]�̸�9[Vۺ�hT�[��u�.�ViΏ/��(�*bU�۫���rݬ�Ncچ�b�fM{͉y˙�Y*�aV��zJ��ٹ����er0�/����殌������oTsF�
6w�=�2D�;���&���L٘����W[�0s���<�p�����C��φ�����w�����yn�G(A�Z�Cp�D�Ej2�|n�V�e�WwV�Y	6h���0I{XZee\2�+H� ڗ��]�E(@��Z��\�Yf�{��Dsh��)��AZ ��v�0^R��̌���<ۮr�q�|�6،E��g�\�6�1�U*6���1���T,UQ��L8PZ�UQ�%��QUT-jʥ�[aDbE��1�-�fL5�Z�B��*��m
���Kj6ʂ�(*(�XVڑclV[QSa�R"�[h��(UQ��dQEb1�,b��Ŋ*�p�BƉF.�T`����D+
���V��P�TX0U��J�R҆)ADAk
*����K,��PQ��c+am"֢��0qj�PX��ڨ���ѴURڢ-��YQYX*��J�Qb���[TEe�jˋ�XTDem���[P�e�Ub1E�4$�@��[���[�����j��l�C�E{�8e�j�X�������Y�1��I�X#&l�" ȖSR�sB�B��k��L��1��3��1����XImʻGЌE>lK}�ia�R&C����-U3R�-Nc�<d�[��`���eͳ�f8q��>�K1��m�����KVmv�4�N1=�� $^�j5���Fu=�Kp��W)�RTV�x�`�l�:<������1Q��n�7A%09dˊ���ښR�k"hr/�c7Mq�^]ep�z��u(��]5��UҺ�ԧR�)��c��>}�5k��I�5����n�<C�[����4V��X�R�z������9���l������ɡ>�򮧵�/E�:�r�E�P�v(a�ךT#S'��Ռ�Ҭ�'c���n��jh�g�՜9���{�,�z�9u��:SZ��v�ԍ�O�͌��u3gV��ݮz������^/���B�+I��9��/on	|���]��/R�FT�ttlfA��"	A]��r��_:&+��w
W�VN�#��7=w��f���s�c�m��=��!�{��>@�&Qy���$�!$���\�D�!�c!�6U�"�Y��W��85v��(L��gSOd�oce�Nd�x��r�ù�lɣ��_OaSf��j�!w��1��8�.q�X�хTQ�Ö��/�z�����W"bgˮQ{�����vEr������R�a��[�{�ֲb#���:�&�����N�������Ԩ�r*gl���}�m\�&������y����;qK�J[`J�p�"���da�97n�IkY��l
3tYP����N��� �[q�6��[3.��%;�]*���O:��#G]��ٹ�yu��K�S����UG�T�+��s� �=	ѝ��4I��&�mb���"��\�o�9_Pey2�V�܂�s�CU,���l�������.��{,�s`�����p�Wz,�w(���@�Q`^�7�a��of�!��3�'8����f�eE��0���������溵%`
��^�3d��
}���+:�7�D8`Ŕ3�5�+x�tA{5v|� ��쒺T���7,Q�ww�C�'u(x
�%56�*�����8��$4�gI��fٛg�X�Ol�����ev�\��a��7���-=<��Ǿ��NOZ�K��7r�M){�Rdz�H���uV�u�e�M=C����8k�L�8y��X�,W�;�e��P�'S�<�X/{;#y���uU�scz�:-�l/���c����G��ɝ.��X�x���4)+$OYq(�m�-���l�Sq���v�3�b�u���\̊�Mr-l�UNسy��bh�_[�!�H��gc�������荛;�K��!��5r��᾿cu٪��v}Ox���Z�طIiݫ8�r�]na�M�/ݱ��k,G3�ҍkuRli�ȗ�U�Gr���un�Ѷ�n�E�Z�6&V�X.+`�,dK;qJ��v�������k�ν3D�b�]A1�7�v�)�Y������ë�c�/��`�<��_i{�L���N�I�DַS�(h�Vl���2�C��݅��=9�Wg����e�[�Q�]n�p"�!ψUn�Ylp<�����+#S�1�m�a�0�;PJy�A�sE��3�e�K;M���d��2)	�:n%�\F�^���4&�R�a�nr�A\C�8ܷ�}(��Vs�[27y+����&B=sU�S��Y��GlZQ�ٻ��z�8��z��e�����/	��W��X�^��^�F�N�F�ۆ8��Ԝe�'%�E��y��콰~��������E�o6��nl�O��Nɻ瘡��٭���벯-�8а1H�W}�^��F��I�;[����0^l��sñz�,f�Nm�L��Mw�)�S��dv��o�2��̻�,��YXsz�cVr�f1`�y�+[�J�rs4˧�Q| ���N8z��՜|��TV�/����c�<��'X�{ẏ<��)j6�b�y؛��_�����#^u�m	EGڽ�(8��y94Mef�=����[ÉP�U����5��w�m����ᵄ��:�h5��D�JpYܥەs�^�D��']��`<���_Ue,�=̨<��QcU��!���-:���X$�ݥ˸r�2f��]=ܤ���j�:#�C}L83���nh���cV��]��eͼa�\���m���]�Nٻ1�v_Q��,���!��B݈�d�uy���][{Ķj5�1ї*6�'�ĕ����c0�k���yCk(��n�j7Rrۑ�s.�+�	�^�Œ���a��Q��M&8��aMh��'�pkD]����z�9�On%���֔3ԟX�a��>|���}�(�9��)t`wݓ �C㕼�L����o�%��Wh�F"�0�e�g.B�x��|k�&r�y+�,n*+&h���|7���Q��ٶa,�(i����R�­4�����[��#��8(B�kb�E��m=2�`I�ը��Z�37�O>7��[�*WY��Eu��������/cw�oN���i:�νaq�ۑ4�9nc7H�5yt���=@7F���Js/d�[��� W�k�~��4jr{��c5���
���>�[<�p���D�s��❸� ��dV�u�GywP)� �l�]#nom�E<����3��$G
�F����fᒐ78��;��a����k�>���
`��R����\�PaF�cg��h�la�hJ�53l��+�&������OrHRkh�kz@z�����r��ӓ���8M��k��z���z:�n3���P�L��=Y�_i
���y�Wr1���C��q�Z�#��Չ�^��<�z�.��>�a�7ux�{ـ���՘��&Aꓤ��nt.�/����$�/kˎUvRb�ز{3[���]��(t%�+/��_2@Κ9�92a�1zF�ͼh�i��gX6�y�/�Z�!e|�^�^ީ�b*]��6�s�L3��������,w-��� +�[�5˱��a��#G3��]ν��b���D��*��F"��tX��<d6˼��ݍmb�_hSLfv=�w��*{����.�)弁�����\��=����c���jk��׊ɜO;����sW:P#�{�@�{���E��2���)'(f����l�(I���Y�{�(�:��Ckջyo�f�ӼI�G���w��9�F�L�,�o�'79Ȁ<�$aw+{Sse�����S�[�s��M$8�"sb�S-���(�}]a�hj�԰��H���1����s��O��6�]�}�����YNgF!;[��ђ�D��<���Y�nՆ�bUR���8mC�ʼ��ㆰ���,S��� @�^!.�c1r�!�y�{�������y,�����f_�]Y�w��V�u��0�R؋���,ʾ�:��GZ�(���{�_hzvj�C�͔�kL�1y4�]-\�3%
�A��\��\݂��Vs47�a���y	�z���K�5�s��f���N4T7���u4��bͭ�����w�s�Z��s�h�}����䣁r7��F���gv��Q�>Z#����{ٽ/ >AV�.��W��k��y�#{[\*��yk��{̩ż� 󏵌����p�$d���6���0��Ŝ*�<�[��&��֒��J��y�H�c;���*ۑo¦�9��߄b��X��$�km#�����D�Hm�7"��]}�-�p)�\w����mr���x�뀜�9CI�n6ZRWb�v���D�Y7��Hrn�7l�/n��:�l��.�ѭ��4�0�
\�t$����U�<����ۮ8��J&�t���yΈ��o��:��v>���Ms�t"� ���콺�T޷���-���Yb:@�k��Z��Rl�f�:����O�L�����{s�I{mt��t\�<w��]�\�h�+�I�z��U�1���ځ��w!��/�ȥ��X.6��^��1Kݛ�M=���Y���1���ݳ�;�����H����1�;<�b���2�F�Z�Gl��S���/�FPlݴ`������8��Ta�3�t��^�ԜO��4�;M���ٽ�D���	�Z��=;V�FXh�rH�Y\�"�g�����+��V
�,�X��w�X(�-�ߟ�4)vr{˶�5G9�=Uҗo٬��^Zq�x�k��J-s�Lv��K;gr+ѯ�N�_�����r�6��S쿎�����\�ꍓ�C!ڻ8�/�]��J����Y2�`\kr7���`��B��.�5.@�P���r�]�Ŕf9�'UއZ��0��	���n�W���y2���Ϋ��LNt���T��e&�D���~�(��NB���3j!ے�]���b����w�#�v��kp^�
�[d[�n�l�1:+=����zL����Z�2N�HRo{n9�!��)�ү#H��Oe��o!�0z�����ֹ̲Uf�ʀ���� �ל�=�i�.Ә^����Ğ�����);�2X�'��x^�	=���$u��ʌ��ٹƹMcJ�F!.�$q�}Un�v�}�ׯ5XW����ˮ�����`�|qr�o��V�u��[�\/^\m�<�R	��Z���+q�x�[���du���8躥�e,�}}��.�ns�Y{R�CNL�����S�ݸ�o���7 [�8��%d��a��n��ɚ�p�r�UY�^��7[�`�$��]��P|8�}��]+���㎃52VjX��i�΢�d�9�P�A�^l�"���f"�D�x{,Z�6�Y&��PV�4�lT5��n���Ùnd0���F�s����ܬ���ʨ)(�2��F��n�ș}7_B��:�l6�G�cFހ؂=�H��y��ݫ�׬a��M�Q;÷�Nh�W�«�����:�4�k0���t�z���P�B�;�9�e8�B'ݭ�	��c��n���V�� ���ڐ�a߾SV˔�h���@�=`ާ�Q�"���|L���Wﻓ�f>jǺ�/M��r�n���&
� ��g�:YS�:b�!���~�����VP��R7��w*u��\ѱh&�"�hO�U&m%F����Mns/����+G]�*5R<mK#�m��g%�1�ذw�s�U�9�����UeEN�kU���'h2|F��c�w:��&s?f��޽3���u�P�ĠΦ޺�Ms��ܻY'
چ^-jz�b��]Z��KM]u���a�[�a������_
����.�i���i�aM�@���!��%�\�ď�̃�v���Tn�YkU�\ս��Y)��wFN�Z'c�´�����$�$�	'� IO��$ I,	!I��$$ � !?hB����$��	!I� IO�H@��	!I�@�$��$ I,	!I���$�`IO���$�`IO���$��IO�H@�z��$��(+$�k,��+ b�K0
 ��d��H�w��*���F�2���i�iE 4j��*�AU�U�(ҁ-���m��ъ�TUD�m$�[hj�*UT��X�+fHQBM[kT+M&P��Se���3-�+#fz7E2֍�JZ�l(�kT����;jj�,��$��%3U-�V�MUU��,m�K3M6U����ff�����,6�4�ʶ�5���ek1���֪٭�3Z�Q3am���Mj--�-�Y��Zر����Hճfm�&��T6&��� Uj%���m�E�)  �w�M�
��]�R�U�:��6��7q�J�T��;�R���ՃVյ;S�IJv3�����\m�m��4��wcm��iVum��v�&��5�Ғ^   ;��ꂪ�Y�]խ��Cf��C�6lˉ�Ƃ��+4�[m����A@wp:�1ӕ]5l��0iT���0{�P�(� �ƃH�ml�mkM��[�تo   kB�
(P�q{�  �  ��0�=(P��S����B�(=�{Ɔ��� (P�nyx�z(Zu�M�Ыb�L��:����3Nn�clԪ�1wj�6��n�-��ӓ[J�Uf��5U�   n����Cu-�"��u���J�U5
��SuӃ*��N�հ��53�qBh4,�����6.Р�UWj��ڠ3�T,�ٵ��Zi ڪ�<  �<��Ml�ݦkTڰ�E��j�Xn�EAJu��j��AV9��m�ln�5J�f��չt]X��#8JN;*Ͷ�m.��ʬ�����4M�*^  ���Z�Z��H���8���V��40�R9ۖƁ��t��e�e��i�dR�  ]��� n�0�,��2�e��ڭc,�!V��^  �^ 6�M� Q��� m���An�� ܸ݃���U�'pt�5�4 uյ�U�ƨՓd�md�j��  ��(zpF�W@jB�;n�3�Z-*�ta������P�۪B�ض�cM2i��X^  ���w M�9�
a�
 [����� h7vn@�0 �-�n uU �g��TX�:hV���4�331k'�  ���B�Z�3v���E���� �C���m��nUƪ���۱P�����H�kaeʵ�m��B뵆Z�jwuB���S�)P  "�ф����`4�S�<FUJ����� j��	JT   a�`L4d�&�x�� �x��������x���ۃ�=���?�F�����F��o��!����Kb';�_����I�d�i!!I�@�HH����$�!!I�d��	#$����~�?��������wrO�q����s!>9�L��/i��j����!�)�'��w�[B�'7 ��7]3a9��ؓwq�n���$P�[�bח�V��J�/pVf&1F��S@��Fe�X�z+C	L(++�x�7��^hzH٠ni,@�'
Ĩ���8do(ރ�'-�(P�ԥ�*�3�Tq�B�,(�
�[B3v�}�Xջ�/5�{g�N���oF�gn�r�B
�4-���/J���2�Y�1R%�ګc4ːle�����ld{��Sb:�8����X.ƹ)��w�q�.и�wc��Z�-�Y)mJqX�p�`KoX�z���S�k�
��[�t�D(�fQ4���']���I&�M^,f�W(X7�t,D��"KW*ꥻcF����<���� �'Suv�}.���edfQI�R�vXX��� �_�.���������]W;�EK6q*%�x�dBB5��77J�2^n[Tp
�T���M�-$mm�7
֛b�ѶH7/2ٴC����;8�1�l�Ț��Z��Mgێ�+#1I��i3*���h:�v�e�26VSv�17��sX�6g2��{��4��c����D6��̢pT	�c�-dͻ�o×Qte	�/`�R�z��8��Y��{�f^	klǢAUD����ؔºt�6�wh޲�9y�n�����5��5�D��F������ge��S+D%�u�s��Bb��u|ᛂ��A���sl,�G�����f�"Z��gB%�Sj���w�-�ŵ��v蚹��yjこ�X5:K(5��N݄��*$+	�h�96�$�	���{Cb���0�5��(��CD!)h0����F��a4���7�L;�0lsUY:ĭ������A�a8f����ct��zc�s�fխ���MCuG��Ҟ��7����ۚ�a1dM�U�	�J�h޺h���Z��� hW��֕6	���I�4�-_(�Y1,(���T�%�/�����@UM��a�KJ�郰��?J60��-۳�Qg�{N�&��֖k*B��,B���;I��9Umf�3],�r��6��#S+u��ej��Ŏ,ut���zqiǪT��v�|o>�%�bTB��H�1��G��Ga�Y5��R�m|��N&��2��z���a�6�z����6v��Z�lɨ	l��C����Alɹ�ZH�-kųqijYe�ƥ�t�,Ф��4��B/G֚��-�cj�;X'��e�苻t�����0��R+0[T�Y�٤h��N�Vr7eJ5��0��*�aղ��Z�oj�bɍ
���O�ن�b
��2>Vr�hU���7)��uҧ�6̷ȷs0�p�F:�͟d�P��jPx�'m�Y��q-Gzi=�U��-(��-6򉹓v��Z�a�]���w�naA� a֝Ҩ���ʽc .�⑤vԹ(3��:R�V:7����rm��jX�lQT���K�i���I��:[7S+]�����B]Jz�:��,��7ma�A�De[
dCl޶����s\�o(�9�Ue��WJ�-D	3&*��(!��&���u���c[82ɤ�� ��BmC�>#��y���zqa"�J�,h�d�.�B@#�л7y[)�1�
ۈcz�q�,����v���l�]�[kĭ$�����j�Q�(����6C��:�^�I�����X^ػ�5ޑQ]��^����j�LL-�6Uн�e����H�^�k��1�$�-��?^E�ԋD���-{t%��DK@��5�X��f�
�Fh�%��Ӳ�d�.�������Y`�w��F�U*l��
���'��c��^Uܔe&�ұ�/X!LV��V.�cV��1���s@�ؤ�ma�͛��#�׮SY��KR�M5��m7�p�VSj�oR2f��y�Ե����,�H[PDI���o+6���Dw#�Pm�� �:A�-�*�[U���� ���nV�s9w6h)�J.(�Y.�
uf	Z�씆�{6CClMl1o�y��90��݈ZF��\T�8���v�t���5���av�Ob��p]�c��6c�+E�A��������<���wuO��-F�n���u��t�]��Ï. �Hd�.��ios2��t�4m�a6.-y�q%(�9c)a1�s)�潲�%A�w�\�e�E��{%���(iB�it���x�[�b�֒s	�]n*"F0�K�w��Cj�Ŵ
�n�[�G>tm���CPI�X�f�Ը�:4Q;�[ϴ�E���:y�ɒ�����Q�x�5�!��q1�w�z�dS��p�#�|�c\�V(�,�R�mJ�Y)�(�^Tʼ e+q҄�N��%�ѓt��8�r�Z�KJ��%auz��Ggi6��Z�^[�Y
�+.K��N�����b�۟B��n�X����!)�LcZ"ժ-�M3��I���v�;�w�����Y֎ĽS�L�64�
��h�,%3�i*�8I5�R�蓃S�xB�[��<�ctx�p?C�^�ri%c��l�GCu�5���-�Y3-�ۤ%e4�Vl�x�3	2O�R)�7�y(�(O.���6��E�)3v��j�kB/k(�̳3'�a�-ٶn�,��i��M�����^�����,��.�tK.�W�.Be-��EK���N�qB�N��څ3�I��Y�G7'd�HmFZ�O.��=����~XvTS^�T7�ݗV��E7�Sv�J�Լ�D�ƶ���	P�#�L��GVAM��7��L�/��ֶ^RS��4�s�+5�M�ݢ�}aij�u."CN�s(�[/(��V�ڔ�:6aTQmX��`RZusj�P�o�[���4/b��t��9��Sd����d����wy��:��"���v=Zi�,�*�a˺��	^�!v�Mw�Œ�ѓD�Xs�����ǁ�Ӗbj.h��oB	 ����<�f���e���wVmCtI�D����7��R�t��w5�˅j[�l2�j�֊�S˃J�j��FLh=�/(R1�#E����%]V�,��!��9��h$FY���v#D�z³�����n��"���m2*d�n�T�%��2Q UL�h�R���7�'���;� z�!����l��9���n�%�EC�fGt��9g�71��(�*:"�1f��t���\�]i��^R�.�Si^B"�Q�RI74L��;�A��͠t�5Z5 i�ܞx� k�m��l�-�^{��Ly�W� H8#

r�5oE��eŦ�)�.��f������Q^ #k!Ê;2��=��n�`��`���6CT�ǚ��E�TcR#.iGf*���{�lUZwN1�DAyK�7F�ޜ��j�n������yY�!�>�4.��T �GtL���
1a��.l�bӷ[];��#6\�v�Q`���.��*e]�­7�-a�ޔn:�4n�Axq,pj4�3&Qm�n�H,޳�#��E�f�o.�V5��:|��aލp�P1P���4��*�qR&�J�MN���l\y�٧���æ����7��`p��UV��,���4^��i#hXě��1%jjÕ���\9eV�>a���VjI��:������е)t˘�l��b��2�e�4Q��-��VW�ţ�b�Q�����h���;y��S��C&�pkM�,z$�k��#�n�8��C(A�{��m.����⸒n�(��2
�,ՓPh��eKH���2��Z����;T����I�J��bRٴ/r���C"jŶ���ˉ�
m�5�@�k5AS0�gV�krC�8��R��K+Z�Y;Wv�l�zhU�B$FQ�v��`T��fu�d�je��+�]l�S�j����W�O�-!��3M�ɸ�g�f�oUk�(*)�xRC���̻�ZL�_e=��]�f�4�",˷Z�1:��8�X����To)����Ij	ba�X��(�:Hl�{/Vɴ�Y0hݩ�L�E�,�n^%wV��� ;c>�2�'/76�d�ņ����Q�AkjaE��w�AF#��h�Xb��3镦�f�!-�黂�۱j�2�"�zDĪ���cw^�j��亍�*�u-����(6�k���n�Ym�М˵�H>8*�aҮÛ� ��G-�54 ["-^���zi���<�=M�oc6���,Ewkaؤ�f|�܍&�e]ٻ?9.��M����DL�C-I^Y
�MZ��ZLUy���R�.�,�I"�E�Ke1sj��`9�:�w�i��e�h桮J��Yu6��A�5e����ɵ��X�zr
���n�x��m4�i7�*3nV�F�.�1��E�Nf4��ͻ��F� -�'L�c(<�r1�\�0�-+��h�ʂ}QZ�&�h��6Rp���V����&�6܏rMH<��̌D�1"n�� ���&0�<���*�M\/3�ٸի�f 	UٳX�\�bbzQ�.bEf���3尷�̀���*��YN��Ôbr�*���p�DPS�����L����k
�ѫP��h��r=cVt��D�;e���uM�P���f+�W��G!9eX��E?�Aj���iҪO��	zZ�B�݌�u+��we�S�0����l����s-�;��qdO{C� I�FK��ͥ�i��є�7{�j:����c`2��~���=&y֫[y�Ɂ�Y*���V�Q�x�)4����!c�.�T.,5gX��ͪ�Y����L�W���Qv���#i�L���'Z���u�kԧ�[��4����[@�,S�\X��2�+@�ޛ���&�U��%�Bj[&���wr#oIMah�Y0�or
i�E,7*̛�X�W.�;DG5�ɸ�Gu�͕v�����6�ǯZ{�I^兴$��%I`� �ޛrȭN^�P����#�������Ԭ(g�n�FQn�3R�
]�ӏ(�Oo#�z�lݶ�������eVZ�T��j7��kz�
	�0�:rC��*�]�i;���h��&+���E�!P	MZWn����M���A�o7d��(��Km�-�XOl���n��K@�/S�셪HS�/uf�q���Ե&�E�u`�sWƳH+>՛ɇ纣;Y�U���'y����n�^AhV* ݦJ��kne�;z�02&��������b�K��B��b�Zy��`f�a�-��i	Q���
�&����A��&l�`�L:q%�y����� m��;�[8ia�G0�Z$0�̦(D�o�&CJt�@.��<��\A�j	����47n]�vN�R7NlMU@�������`��b�ML�$�Y ��F:9@�5D�%G`�L�/v��j�e3� �ne��rbJ=X���u�/Ǣa���Or��f��I�`���%F��B���ق1���H匧q#�cI��EIi�M��	��t�kJ562���ҔѦY
	t���)-�U��v�Q�l\{c���d6Ѱ7i��^�h��ZFv���4���Rxgw`�82 �!�fD!2"q��@�)��T
z���ͧ�rƗ�[�DؾГ�j#X���"[�H@��Zp6��T����T�qؒ�n`���W��)�Qt�z"WV�,+G,Y̫'��lc�A��R����������r^�:��䂓U(�*�������ÖVo0�m����Yz�Z�21� �NhF��D[�u�JrCh�z,f�Y��ua�vY;��*k�c�X�A	E(^lyR�)��jbq���m˚wf���q4�_as&]
�Ԩ<ƕ`	:���6�WGHãR�hn�7�VA��0#.����;Se�r�14Yv.�J&�!r*E�����c��O0�0`��ɷ�-:q�F2��ù)L/�o k@Dk�K4a��%�]���y��H��7f�-c�F�7��������A���斶��H�̖�B�-���Znˢ��]=Ӎ��pM���%Y�B)R�L������w[���v�u
Vtʶ7uˡ�GW�8.�(�n�6H�Ӕ��![�o$m�8z��ƽ��ށ[�Q.��Eٔ�:øR�+X&�@C���E��Ɲeljs]�H�=�a�v�1Y[���L5�Y(]ju3q-h$�g4;H��U�'sULR�'瑮Lk��C/�=�$9p~4dj�onrH���Y;�`�ؐ:,��r��F���Zɦ��6����U,&>ܷGK�[�3j�員E>A���Ȏ)�f7���`��KvB�nBr�Z�&���ҭ�V�l�RV�
=���V�OM5	*�ǻ�sYuw�e\,����k(��30��kS4pZn�f՛��)P�r-���w5(�bq�û����kH�2JL
w�tp�)dUw�X��7����D�=�!��t��ctp��ɑ�Ǵrs�u�aEV���Y7*�&X{#�ϵ�� ���z���r�l���,��6�/LVn�
��L�ӥ�b��F�l�fd�F�lQ���
p�n�f5��L�U��:Ajȯ�[Q�(G��j��8�{[��
���W(���ˉ16TYh����j�ف��PCFӸ��X�������T�2�%�p<��H��E;W�&�:h����U�h`��C܈,�̰����{G3R�3d�M������LJU��X��L�v��p�EL$r�&ź�!}1�ZFn��PÒ����;i�Sw�rk٣��<�F&�g�۪C�w.�
Ė��z�.W��B��F��	N.�Ƀ��Z�Y����Ko6�#�-�`�<7+�1.guwd��U�WjKŭ�Oy�Sw�@28�ɯk�!4��ԏ��_�m�*|�$�l�O����k�u3d皂�����B�v�gPx��]4bi8�7f�j
�O�ٮ��g^蒔N.g��6����<��ቼ}q5,������]�7��5�Yȍm(]�@r���8y��_W]9%J�w�c�T�[���GvG���6dr��tT��t|Ay+ᦰ�҄b �h]ڴ)e������Bᨯc]�X_s�C�����d���:*��+��)��<��a����x���
 ͆��hG�g#Ϥjwv^�u�2��%�,�-�Ba���k��0�|;��7�`f�����}�)Qj����{ݾ�s�S�>Ȉ��
�H�#ur����f�=ɧ"�����i�8Uk�;�L�,qZV��߰��:e��5�]�7�a�:���Ԅم�k_i��E5�Q��+E�k�Imyu*�Wu��m�q�M��7~Ujw^�����>:4��9pwϮH&� �*�q�.ܘ
�s뮄�bb�4#ɜﰾ��˪f#;B5#�sT��B������>W�Q����ȵ��ǲ�c�]���O6-�nq�Y�N� �Ϊ*���Y�SkM�����<Gb(��x�8;�pY��k�
����}�V�@D:doSɖE�}��H�9B��,���D�m�IAy���ܾJ��3l�]��r�I�p(�#;��L>�&*J��[lΟ�}����E#�n�ܞ}D\_2�F��zaEu�A���C�L���s�� 6�_.U;��vo���8�_(q����<4�݃�RC�#e>����AG+m�#qhN��o\I������9��ˊgܚI�
�����z�%��Y��N���mv>�Y�|1:���79$%�v��J�"
��Jȱw�;}��b$�}_�ЎvZ9�$]��[��Dp {n�%��,p�kTk�&2��c"w�4��}؉U��d��m1:��ب8L�&{��9���݈l�u`Wf2�>s��x)D^Y��3隍�ʂ4A���vM-��攣X����X-63�l�-">��rYT;��q�&��T��D���s�q���{�2w�Jz	�5���6��}'^ݱ�4e��/�2��y���Ћ�B��rx֕�G������W�pq�k%�נF���(�^;f�d�9����W*#0�k��|��	��[���gW?u��~$[���ƻ��@4���g9%��_V�/E��Z�`���s�M�16OER�egWbF.]d>��WjR�}մ1���t��wC�כsX�S��G�-I��1�ke�a^��UF{\�7HX�Xw5�"1!�0��(��P�۬���;KqL�2����a�{�l<���t����岧ss�ֺ�;��ǧ��XJu��<�K7h��� ��V	f$U��Epu�|ڊ��υ�׽������j�:3��R'i�;f�^��{v�X�����L��v�]�[H�a�_;�����H	��8�YlgN�t�O����{��p�y�C�8F���g�M�+���E��r����;5]��Dڴ�Pw]�(ͣ��ۉ'XaC[ )�*-뱲�m�M�f����7jb��s�k�S+�'8Ƹ��`N����M�B.�^��2��(&m}ǣ�C���"Κ���w�cAs�,,yb�p����_3�b��ɽ�(re�j�ϡAv=����@�sb��_-�;��:K)N9w�8Ζ���oh�8��2CW;���\ ��z�,)۩w"�w�]t�����굏���u6�9�if�����N��Ɨ1�:���p�TX����P��mG��*Ôz�2���[�26�K�r+�v��w>�o|�c��j5�������|�����۷��w�&����k�t��y��'�IL�ҕ\�il��5�0�97�#*��*`J�L<���hT�Eˤ����{N{�3�Mg�Dhm�Ȉ�4½w#;��Kj�o���U���n^u��.���j,�O�l�Puܒ��|� ��ɿ-5�]�.�;]�y*�ׇ$X�i"�7��R�#7|$ݡ���/�&�51�V�j�t�ExS�/M�}9�bl'�"�p��G��+D�c�㘫F.9�ܬX�٠d�z2K���9:�K������niկ84z�=�����T�#�e����0z����������4�W;.���r��k+��X���{�O�뮨|�	���9���*:��`�N�oi�1�B�=G`�a\[LY|[�P�	�3�f�]{ג�q���t�{jS�V��e_f�4��h�IL��!Y]�:�	n�����N�@�.�g���8Q��`� PkK�vmG�N�����cޚҩ��驄��k1e��T�#) ����/ ���^$��Hl�X��E^[+tW9��#�yc	�i��x�Q.���ݔ����S�z3�n����3.l�����sn�}�:� 6�3��B��4-w��8}���c�'���{�Lm�JT�c_(����[��k)������/`������v@����;��2�.]KSn�wJ�b�Ï�R9�Ņ�*����tY���Ř����SR^[����'�yY��O�͚ʝ�J�d��ފ;Û�C�݋��%��������_��ti�9s�ok�m��M�+�v�A���N_^���v����~3�5��r��__�p���ɫ+i�'u����F��>!n/gX��z콀oA����>}�kק����g�����<���3�xAY��5e�`UNp�}tqݿ3K�.�SC��\�Py�lCj�Bۆ����9_k���w����+ao۩�xo���`C��R�b���w�v�W׉�4x�Ċܲ1���O��ޣJC��/��u���):�<={M�j�hj��Ҡo���73\R���������D�/�^��ں9P���%�͈��H%8���/{5v�v>K��{6�����{����;���&؂���T���z/^7k#uY;���C����A�u�
�̸�><s�Tk7|m�7�AcϷY��I.����T����� �[z��ŏ�$\�`l��wk`�h3���K����X�a�%= ��d��Y[2h�b��R�[X���ƴ��oh�<6L�sG�V�IU^��#�F=�۝�v���Xpz�z\�-r]��Z���(~�2$3%�V+ڹ�d-Y].�C��ǰK�\���������;��M���Z�U��"�B�ؙB�'�6���ո�z�5���6�#[�c��I�k}[q��5H�8x6�yzt'BU���>�1`�ㅵu�;���i�Evz������̲{S�����r;˹����ˮ�r�2*��p;�tUr��R��|pKʈ�v_4��_I��=�@^�gN��-=�Fyky=ۊ��Gy�$:�׀���ĺ�K�� ������5C������p�1����� E梗��{xz�rc��g^�C��
������k�}|5�5�aW�h^I2�ĨW�d�e'��j��W8�����tb���c���٪��w��;T���ը�XmU�u}t��4�nRR�l�!\�،n��#���s�P6������{F<<_e]5;u��/s��zۘN$�=y@q��K���Z����5�뤦�s(�h����鶟�ꖱ����%�jk���_��4�ۧh��;��u����4��f����fg��$E�.�n��9!��0�ei�]��)�.ⱈ���8��1C��۝�,�����Q��P�3���q�&ɑz��T����q��oN�Vq�2�� �J43z��4M�@���p��VxgR���t�ߤ䳖*Xr�s��e9�9�a8�熖qۍS���0����w ٲd]�@�-���LLb�+���ɏ��W�Vn@Ր��!�>��kz�a���e��4@�ܼ�*��k��pR]��$�?lږZ���oC<=�l-��rܨKFga�MfR�v��n��Ƴ��MZ1����gi�p^.�|+>���σ�3�c��;�}�*����S2;��I��+�*>AU������`�	��a�әr�u��#�]�����E��Xo��+;V���/��eZ��1�&��,DO]�n��"�J��/�0J��×m�uم�	�Ye0��ҷ؀��V�����%\bB���a�ɸU+C9_S�.�m���E�Y�F`��+��D/ �yB�E��g�����i��0�҃^E.�`Y�\����ݽ��]Xx�$Yfپ�uz���|�0*��gpTzҸv���i��Sį*q����.�����X�)��8�-�r�5^W=�w&�[�:OO|1�=V��L<�e�z+�I�r�;jc ؾ�=��H��I��OÊ�冱W����)���i�1~й�r�X�f�"r�;,0���I��uM���+v���9�H��]/�P�c��\k05��)܇lև�ZjT���򣗂	Oy�s�����5�SU�\�'���<���2ş;F,籷q��[��8�A!��K�=}|YK�[7jnSo'(�*҇JL�]kP��9++��r��=[�s�9�dt�����΃|���x�āeK��b��0��(nnm������K���&�c/���t3Ԅ���s��Y!p�jg�t�0�����ûz��4��>��IfL��@�
��]i�a�Z���M>�8:�p\]�8Mtw���E�[/`Դ��}��.D�-�"7Nf�sK
�-�t��גډ�`6����r���2�u:G� U�Ky�=N�Y���P��l��s��x�;�̭�ݖ �ʶ� ����܍����ׁ��9��c�x#��$�{�U��Ɗ�)k�D�9��
�/^��yN�]�N���y6m�{izO1�r�W1m^2�;��Yb��{��M���F��Ι]����r��<9z+3u�5�+�n��-�
G��n�����ynF�w�p���j]Hi�pV�+mw�����B��yb P��
��Cr�{��ެvn��G.%>��QH��?{��[�
�{��.��<S:���WC�����D��V^!tm��>v��z`f���Y������3w,*�t��}�n�k���p�Z�P�N��	e液U�QN���%��%��%	�
p.���Lx���a��)9aC ھ#���j�M��7��7�:r�ͨ/y����V.�M&�ַL��c��^ޡegO�'wǭ�GvVg�0�)��l�ጲ�F>��C���zgh彚�EjN�1u�/NA�����7{)#x��G�v�p|�	ӛt��Ԉ�Y��/{f��+u/I����<�{��I2�[�Qx�4���p���X�~�vAv�e�V[!֦��.q���*3(�!�2舾�{��;+_��D�޸����y�j�sY��r�Կ�u���BerW,�����r�dTgm�^pa&7K���!S\��r{��Q�r��ed�"g��
å�˳{�ىJԉl�;ř,Kh=��Ӧ_#��밺�uf�ae`�M�*�JY�\�Y���Ŗ��h����{�z��W�O.ğ�"�Ѱ�_Hn��&oϺ�	������N�V��*�X�Z{KQk��9v5ZW�wY씏]��pܽ�{�X�"���޷�P�'d�QH�#���ه0�8->H]l�{;�/A�u֭��R^�ma�ιɁ�����93�㻋�W�(E-�ܱ[튑���q��/�r6"Η�|��N1F��%�v��{�x�{yک�k0e�-*�hJ�%���o�'9
[3�Zu؉��T�
is��d�������~+��
��	��3��ҧ �5��K�.�8��a�Gf���1sz�8���{V�"�V��rK��z;���*2�J�j�ѽ	�l��ե�W�L�/��\�k��6��/j�Di羇}9ظn��Ѽ��w�D�L����ȴ�k�;�*[�:�-��F?y���!+Ê�0;����FaT&Jս��T�ΛP�)��Nj0�7�:ɸ��z��M�d�w:�伧R �_A�9����-��S���8��dYᅅ��#����\�3V�uR��qR��[�W�9���.N��h�wm@-s�a�{��V��V��h��y�vL�טA�՗7�~OQL�y�^ȫr�Fe���)9�p���^%QNT=�c��帨��ns$^�ğ֬�C�0U��u>xr�{}�ܘ��͘�0��D�ԟ�=�R'��=)пw�����t�����G��26�u罞�z)i�^Q��{�� 5n<�ϞaԆ���l	��Ev)�؏7�&�n�����4/q�͚������}�)�M�]ڶ���B���b؟׭�m�kL������L�鮆%�����;a�7@6��Z.+�!����":ӡJN��T���]��	�<䆣��Q�'`t�m{
O0o@7�<9=�|̋��l[d���;Y��L���	�y��IFw6���8X�Q�\�33��FM��ΰ�&���e1�3vFm�k�r���;��D��d]�u�i�Z�Ŵg��.t�.!4ǜ�_%��}	�F�r�a�Y��Wd���瘝-�W�r��f��e�k�}���Cx&y���x/�M�����;{w�͏W(�WR��cb�~ ��z�$���η�9��@�HH IO����������"����Y�7^'(���;r�o�%����.<��2WPB'+�k��hn���Y{�Z��2vf]S#U����ER���.�\�h�Y@��:�����-z�o$���	��}z�����dV�k����Ã����,����dl�ig ��k]_s��&�Y��a�I�X}�0Nۅ����}{����OG�23���)��ٚ��돮��R���0�¬����[\hY��wE���F<��ucr���Y�n��'�h��*���}���G�
��ƋCbV
�7��ӽ��{��A.�/*p��	7�z`�yL��[5�����~[��r<�-�P�㫟2~�o#����Ɋ�4ܝ�qW�2Ov�|�+�i0w'R�/Z�Z��.�K�	��aS߱�K���s_k��wΐKR�b>���m��{����y]3c�����{e�a`��P�g�tS����p�Ya��;2*x2��G�D��A��뚏��8cu�.Z�K_wpؓ17�����c:�����,4�,��3/�g&�p���M���x�׮���н�Жrg��ݡ����%�X8���-�f햂)��M��Z`�5"�^�d�.���0���v��v�e�ҙ�ҵ�"���bw�[8˧1.ʹ\���+�<.� {��_|G_v���$�0� �w����9KnVFi� o4�F�4�I��3��\��>�����.�2���F��u���%�T���[f�Qwo]����;x	\pe�h��0�K�Y�%��	$Dt�V���q�G}a�d4�[Be1m�����&
���8Y����8r��3y��gcK�*`޵GV�O,ؘ��?:����T�Kwc�]g�õ`|nQ�q���m4��y�I�	w|����Ic=�\,j��5��y%�K;n:9ƈP2u`B��!��եK\{ƧY)=֑\A�u�¼q�^�0�[��;t�M�\/U�渓ő��B����R��9�7^�z����;��C���V���=��[HT��U^��N�A!Z1���ǽ�:r��cqd����b%(+��ιn�}b��.�D���.^I�n��܄�e2Kyח��jtqf�̝;'�&��s4E��A�uUy���"f4��ts���O9U6pu����õ Fh3lڱK~J�rnn׿D�ٶ?y�ܘ�N���k��Q\��:��;��w"�o��8�#�dwkzB��v�K�1:��pHr��p'hѸ'+�O=�`�s�� �J�α���Ƣ�n���f��"������g��7�9;ݧ}q_h�nF,1݌Bf>
�}��w)[v[5d����7C�Q6��䎷D����DeS�5��F]�\���J��W*��璎������������l-�@�w���>����o�8�X�Y�g��ɫO�[c�p��v9��8M�6��/�	��nE�M-л�����5�,��jK%����n��Bړ�G�ҝ��j]��w,�L ���9��&����Wx�.v>��;whC'.��,���ˡ�YnP)�^�P7[��d��+�zBE��L1
|������Z���zs�BVj�F]���׏�^I�^݅�Ca��yr���vrؤ��[�sYw7x��ӄf�cZtT܅�Ǽ!�>���W��s)B~[���4�'��e]�.�bֵ{wd!!׆���lG��fsf)��d������_<%\PR��{���mΈQ���L|������~$虼,���L[r�ɀ�`��%����uB�x)����,R�=̴;U�ܻI'��K$�s���ݫ�PN)]�`�����ut��]�!ϟbܬ��i^�c�r�y��r{���	��|�q�������h\�Jp�볊�vʬ!6t�e溿�]��lq�(j�D��+�hc�Ә�f�_i��35Q�UfY�����k{�Þ��� :��M�Q�4��V:�ɰ�����w�~�z�izڼ�������<���t;�c/:��N�œ8d�aݎ�jg��m�6�=)N���˝�춥�-E��v	΢���/�C��=',�ٗ�v2�cJ�0RsJ�
Ʉ��`�s�3ɜ�z;i�m@L2�N��j�3��)���J�/����6�H:�� 1��#�c��^����̌Oe�i񻐰'}I��s�r��&�j�Y���XE��ܱ�i]29�{Ȟ",�|/��{��jf�/�V]���]��2��SR΀m�F�K��3����ºk��f(����ؑr��i��.h�)R���ح��!f7�Nz�l�ݴ���g���gD�%Q�&n��7&�	�_������>ĳ.�Yz�j���g6�WAr��+��S���K)�Fة���v7��J�QA�c+%;�F���7R�S;�GM+�������I��<&_�uF�v]�z��u�B-��e���
��^:�s��k׶G2��K1ӷg�ۓ�-���hP��$�[�G�;f��p;&��s�`���`[�<��S.-��ȏi�úĲu�qgR�ik�����k%�Z�.��f�O�\��L{�WNVG&>7ɧ�Ɲ���^6!���N�4b��{&�a�Q����Ah���aR�֘Q��M2�cGX��q��|q�7���go��f.<�91*M��۶]�^�Z"�E����r� OVeLb��)svm��8�Qt4E:�S� �^���]a��Ok�����u&
ŝ�kvu�7�(�`~�ח���ƍoS�^�Hw`��3ןC��������������}��&'��0zI��jNl*�oV�������z���(�����n1��r�T���cH�;�ݝyi��u\8ұ2����Z!�s���)4��cn՛�XQ�y�*�޾���]��w6X(�y�%g*L�5�����0zy��+rP4���v�W.�V�����MWt���a��ѹJ\P�ُ\9�Mj�..���@�Z:�ê��U�n����W9$����ȯr*InhR�QZ����45I�Up�s)wp�����c]K�>~�[Gv�RZ�n5����ݺ�r����'�9�B������\�s��K�f���sq�}��.���GV.�'�␣�`�����%���R]M�{4��DS!���zj��"b��R��kVlW��*\�R
:6�����lF��*���1�ٚ���Zɋ嚹�#�'R<��ھ�Y��x����wu�ƶ�8�����t1����w��u�qf�"A3��б�dS�[�e��0�y��Ax�Q������P������Bڴ5����o�!��V^h���tgg���@Q���u����V&����\��ё�8(<9��NL-����O��%����w�P�a֥�oh4���a"��5�>ޡ�aY;e��F[��Q<�S����B�ٝ��rԛ�WK�Ҡ87mDz�y!�^��Z��B��W<����ӧ8��r9���6��������/��� �Sgr��^�;��<�߷n{I#�pj=g6u8v��pG��Xd�@X��n�$��4-ݻ��S/ ����o�C�c.L�Ư,�9���!-��� L��&�:Wr�Kr�MEu]��JP�t�^N�52���{��ઞm০�����8ҧ�UaH��w�W�:���0i1�B`cJ�ː���f��9'i���3�����.,ݥ��5�:a���70.�i7��q�'�p��N�u��@u������%�˰-Q�v�-����e%%���6�vL<6N�lb�{��вU�8M�Չ�Ss���U�}1ҋ�|m�B`��|8>�Wl��z����.�]�1�"�����j�A�Zr��#7�3���LY�uڝq�A$�\��W��qeb�������۫���{!�J�ObK��֗^x~a�yV_�����V�q��
��f�߂��娆�wX���(�4+۟i�{��[�澕�M�UC��)^NӧOp��+��(��k@�B}£G�ە�������*e0��/�-@0 ��д鷂X��ɕQ�x��`���Z���/X�����O����y)
����.���XX��{�i\��*�f�UYD���!M�+�R�ÔE�q���h0^����>4���v�1�k��m��qR�4�g\4ƸSS��l%���	}3٥�c�i�l52�e���P���c��!�rA��*����ڳ[S��\l4p���Q�Mf�o.����\��u�ƥ@-n5a0t��.�ˎ��:n�G#�������ޘ�xn[ݴ�C�iw�d0V���w�IeGԺ�D`��v��3�v.c��颈�:pf�.�s:�y�pi)���"�BG�����i�bK�ӱ�o��߸��X��O��}���2p�QQA�ᛃ�s�M�7`�=�p�o�ƻ�ȱ��D�X�6�Uꌈ6�ґѧ�Ab��o*������';��1�V(���k��l���4���ࠞݬ�U�	�+���e�L�ۧ����eˉt7���\)�&r#.����*��
�#����Bv�2�h�SmVqT����ۗQ��ni����{u[u�B�MLi��LR�Q��a��b�gw
k��=7��c�\)W}��R��kH��Rɉd)�u���_6��3�V��T��BQJ��9>���]�̛�����j�9Sȸ3��q1�e^���� �����=�;ʅ��=��.f�E�K{-��*L��K�s�ߙ���הH��]��Fv�5�z�V�U"Z���n�D(����E�evYOh��|�54��)k^rR:�lU�SCb���a0��1��A���ɪt�z(��_
.��W���:���������z�D��������W�*��e�U�+7�)��0�2��RԺ�/�O���<*���m���V[�ƞ�Z8|�'��IcB! *�E�밷k�N�����)��t��(��&�͓�Re�@�r�&^H���.�wrq��}�����vm{[վQ͐g.�n@�6{�����L��gU�|�v�"�����E�~����n=}z��e�=�-�uP=��+�Mi�]�穰xǏ�NTx-�W�w|�#�B-�"su�g{���f�`���]�a2�b�YV����1��M��m�PWk�jgƊ'�N,f^4[���9#��ʽ���˰i�@�Q�Lk�z,ۏt��:����F�u޸#Vu<U��Q���gPv{��3h�3-�8�aY���ͱ+46c�y��U�ġ���+���m'�>�Z�
�>r�
��Ф$�1�(����	�� ���#r����+��=���R��6rZz�n��
 _nҶ�w���](�k�ѸB��y;���lٚ�R&ԃ�B֜ᔐΪ�{6�^��QhWp�Y��z�]��!uv/Q�<Z��'\pIV���颤�v�RF.T�;�Ԯ�2z�FeL�x�\B�Mۖ���A`�Vj洋�ɧ��"����W:���k��߬�m6w�]٤�r��c�{sb��K�f��Ѿ\��h�=�a�`/�1�{�W�*�tFh,H�JL3{�c>�糽X�x']�j�DXV)=ڏ ӥ^��~���c�p���>�lbA�DQs=�#l�g
dF��G����
��mJ�e(*>����J��ٌ��8
n�t}��y	�'L�Ӳ���W
ܸ��G�!]��RZV��ڝ+�q�I�0�.���3٬ފ�YU%�VM����\+u>Xv"�f����������
�2�4Yʚ�U���+ .�ɹ���]soR#���W{e~X�ܹ#����̺�}饆�����֍�e���S���zA58e�z��-C6ۥ�T���}��]WfL=$.,C�[E}�(�����:F��(S1Q��f�e+�X�!A�N|�s
�@+9u�n����R7��;h�ŪW���.��RӊX��HbƩYo�0E�Y:���b�7�$�e��`:r�dmũE|*����1:DU�}��.{PL�{:��]|5i�; D�����y8N���s��ؽ̈e�\�%v������-	U,�c�M=xB�^���&bO7��b�a�A��[:w2��j�V$L[�lN�������ry�<�e�Ls��onҥ��ΞB��Y�ݎ!�i^��-�,���)��]�m�3�:a�J�ĥ�U�7eo.���q�Ձ�;nZ<б��e:��2,v0�.�P���eWi���:h���."��6��a0�J�(�z	|[�ҋM�i.X�!�v$V�.��SH�0����>��2�_d΁}�[DP����:3r�"� �Vդ�ȭ(��DO����z�[uϞ^�U��""� ��M��|��ƎS]�R��۱Ba4U,:�f��|µty��Ί�����{�B�.���5bUg(`y��lJ��0���o��_1�w���M�WW�����bg�g4��a��e/�}Ho3�%�٫����ru�}Y|!Z��1Y�ǻmn���J����-λ�FK҂���h���H�'�B8T��Z��h|\�����հ�Xﻣ�Q(<�b\ ^��Й����&����éL~
���bXh�	���"��O!������ի���{��E+^�1.�~��
�`�X]LMKgrz�G�� fl���i�s5�}�Ry��-߶������ǣ��6b�d���OK���B�%���Z}c�utgz�us�$��	&���eh*u}�����q:�L�>�	���b���u*aH�F(����+�'N�����0S���s���h.��݄��:��u����+x���U�l�<�ݕ�M	n���u3sS\-j��qB�)�vj�[��� 
�X����O�:_��-rm�T}�:��7@ה.x��/�9b+^vT��4k.�>�S��͆�������W<&>q��|��!Gڸɹ�
��iAwN!e��~/�c7\��,U������9�"���m�`�;��k���f�\��P�8Vt4�Oe�N0��I�]0�9�q��	�����$:�"�c�<(�=�Eˍ���C3w4��EMԔX�]ٛ]Y�.BG)%�^�כ��Knǳ���R�{���k��X���t����9gz�#�E�Lj��i 0=g^��j�SRh�2����sx�$�����f�����-��})�r�a\k��-����/g:�3�+H|)��G|n>\=t�5H�ٖGd�L���tJ�F>=%0T�	T��F����א�����,S-w!����zG�gA�҃�� �f�]��ݕu�	��� ��$���>t�a�n��)ͥfs��/��W(���S֝=�f�i���f���u���4�p>��s�mo���	a��8����dh�=j�C��>�# *�V�k*�j�ʅ`X��((�X"(
VEm���"��
֪Ņ�)[��,�
�"�m5TE��Z0P�hT�J¡Z��j��²�%eDT�d�j�E�R����°-�(�U"�D*X�U��-��1eX��)Y��ث�TYB�*��)�bl�DV��h�R���X��T*U@Eb0k,���Q�[iiU#m��J,J��X��aP��TZԍ�YU��+�
�eIY*B�F�(1+*(�EKJʒ��ȌkcPX#-�*�DXV��R���(��D�¥mh�Ub�%JʱF���Ak+IPE`���0*J�EDAIZ�X�$���䙫�F��cǚU��u�ù�k�D<�؝ܺq�v���ܧlc�G��f���]�(�Ac!]�ˊ`;��ݗ]�|�b�۽�V����&r�����?����:����C�ϯ f��;�#��F�jK���*婾/
,��w�}C��p�4�K)b�2߇��;j��crE��z�I8k�Yp�1.�y*��̟~�����6�^��c����� ���^���5OZ�d(M���3|h_�\�|��>���̍W�b6�Տ�V}��=m�ż����T�1�s%�]�>����Ù��a��<�=Q
W���^7Ϥ�.�Vz31C��s����YZ��b��D��c���x���7��p{�����{E*����w�Ȏ,�6:�\tn�ř�mu	C�$�����	Ƃ�6���X��O7s��}	O�]��$&q1�V}�v��1�Pl��X��1���F'B�:�
��hwm��Z�I�R�6KLu$��h�!����.2(]��.�����B6-[�٫g����t.J�LZ����Q&ܫP��Kj{�cb�t��7��4����� ��X;�U�1�ru�N�A���7�σ��{�����	��e�A�M��>շ�RQ�R�V�ua~xd/�]s���Ї�Qb=�t;��ы�o	� *����M���b*r�>��h�`���<�i�;�r=�K�����}�X.RNuiuu���bͧ��!�4227]��-��~���EM�^���m��{�	��4�17�P9D���p�*�'d(�E(jA��p�M3}�㣪XLE��VM�j�R�><on�˃��Xdu�){�
Ю�x��X�%W@�`]��
��7�b��kl�D��a�B��607���o����Ք�9^�e�/��8H�c);`��g��1�&5)��k��"szl|�+�,�
w��ށ#�{���u�Nz�T'��1�i�U��N8ȵ#�V/PE�t����A�D���]�ѧvs�Uvo3օ�A(��24����VL��A���*�Ωğmx+Ud-�'�ʥ�/�j�kk����rN��5(o����K�rc`R�rH�[�tʇ4��K`�8ʚ��������J�w͘�޷����~"b�C��c$�W7}ݝ�E�
�ȫ�ޞ6���v�4�9�YQ�13��� 6`���l�C>�}�a_��a��Mb��h%l��+7��m����"��m
���f���^=��K��]^أQU|�Lm�Ia�j�!�6�]JSvh45�!u����'��|�Iwh���DY;�;4�}o8�kN���o��\FV�"o�v	{$�ÊdT�ۇ���[x�=�L�(�uk�����{=4�� I<�jnZm�e���b[��[�.�����t͍�QŘ�dF�P�c�Dh�h:��'����Ed?��2<_ ������h�m�-)��R�jc�!W�ޢT�@,��5 ������Z��Yt/Hk�3���׹�dm�9�ݺÙ�qP�df��W�*)�A�QG����9{a��wls<V�f]�tU������%���q�>ː����(�G+�5y��_H�l�U�1[�t'b2�W<;���*|ơF��q��7�5�M�aE�4��l ����K]��P�ׂ�,zTI�Ω�^�C_���u
�h}�X��f�ɦ�i�y��m �+`��;f��Py�54��7���ԡ�����%&���d��(|�=�l��ꑐ��tj��gT�y׮��"��*��֮$@Q�>O�� �WKȑѵ�c�(�����^��Z�91]�3��ǜ��C�|��Z_r��`lېuQ��-.��E��	l񗞙���8������p�q=�Y������!��Et��jbQ=;��;r�<�A2M��r���wC�F0��;���䮷lZ��{vI���J��*6s��7��"=z��{WB<�J�����V� fZ��.k#�$y+��m\��U?Ttr��=���9$�/¥Ńh�#��QNq��5VL�XZ����Iq8�d�$�s[���+[����la�n���:����C� ������]q�'L�¤�]��v3]1w��ѻ�!�gĻ�ψ�N.����b�@ח��{j�t7MY�g��w�V$�jW���;�J�b�=�`�f �ք�ͺ���`V��G�/������y�����Q��[��}Tԇa���i/���z:ՄXh�s=7뼱��;�$�^o(��_�����[�"����>�L�|��e��a񯓛W�Y���BԆ�=׺�-��J},�a-�蚄��LDŎL������}��j�]�^/b\��f�=<��R/eo�di�v6/�VHB0d�,^��y}c�����ػT�w<���y/7_G�?��Yc|5 �cu�0��aQ�cv;:�{"�)NC���0]�V�l��e��NMK���+3y�j{E��<��s�������=8.>+�����V��c��F�v=��T�0�(d���귩G�E7��!$i���̉A.�l^��_����ɜڶF���fKї�u��o���'���|Wc�M�+��pO�\{��������n'K�^�����d�|,���VqE.���׋�܅H	�f�^����}/���I�����b����nc&��΋6Y�����רe!�lB�7��ԑQbU���Me>���!�z_O���<|��]��T$^��������pŪ�>#B�cY��=�}*�Eu�j$�pT(иL�ݬ�wi�Ә/4���J�=�q�ʋҠt5=�jU�x���H�L�sr����%�P��3��[�}&c����>(�#a� MZ>vz)����Jz>�r%��h�H��ѳE�(F4�������E�ߟ�w�}]&��q�l��\���FƹqFM�P����9��(��N¹e( ��9�~��Tj��6�נ��q�$�+87��Z/'��P�`���ૡ����L��ǥJ�3����8f2p�r�q��VM��H�������Js%�}g�@OCr���|��1`�q��!E�ڎ��ƃ��O��֡3Q�WȊ���AAɊ��q�$q,G���������r%�y�͛X�����s�B��oF	�o��VF�������q�ϟu�4��'���ܞ��L��Wv����8������r53Q�M\�◕+gw<���W�/Up�Ӂ]w�>��U����)�V���@VS`O�-�*9��3���+����㮵��o���
#�&����F�OkgA3)܂6b"��`��uD]%0[�s��FTaϲ"k����-
6f�"�}�v����Poh�WӐc��N���w�d�FVm�-TDk{J��ȡ��m����G�W[l�U��K�
���4��pf7�^U���3���x�󔡖3�ڞ�X��t�+��p-
m߸}�X���\��fj�B��Bͧ�yۢ660k��4E��D6GX�f���0�R�f�����h䮐�S�8����p�dUv�R���v65�w�}~���Q�����j��}**Tj���YM�,�/���A�����&�2�_NL�jXͧ�'���������W`���Na��p��ޛ�o��Ƴ`wR��u��3�p2_�:�Şt�'}�!�l�jht��z	B�U֪�v+���z�;�dL�7⨫�Ư�*Xj��q1�==��K�dXR4����s|M�D%P>�D���{�C׊5R�]�x��b��t������M_j���U(�Yu�%�(�f)�يȈ��j���sUc�7��<e��<�������A8v�W�ܵ��e�]�isب�p�9|;I������K�ܜ�iVj�4!(�*74J!�}�J��槣6u�e��--�;�����imcԙ�u����ߊ���t#�ڣ�m&Άͽ���rJP�b���.u���U���R:���o�\�@(������sFH.�[�o�NR@ى���Ոu�F���wd;���l�w���9�xǥ+�Qm��v�=���,�x�D��=	zE�� \�**�.,p�*�f!�#�l{��A�{zm�7Ommlء�yz`4=�M&*�`���P&���6X>���s��~��s�ε/)^f����ȉYM�ESDT�<�#N��W��M?�O&h�����%�>bly��u���4������Z��/�D� dsjH|*`��󛚮��;�Z����v1�v�z�j���t��>,�-3e����3+� e���{CE����v�и�zY�X���Yǝ}L�GfW� �@�1� ��������6w���E.."e���w����Qs昣RY��7��	��(�4�<��<9TTB����^����9k�
<�ڔw]9�6�V�u
ớfV�·�{'�}'+�V�:���ٺj��Kl�V3S=tL�c7�[��o��>k�3å�Y|}��-���Mvwc���;���'L����T���l��dy�p�8_d��o98En����_I�g���YȰث�u"���&�z���^�'���:�W<��,�����cj����R����K��q:	��zl���(�R{������e�tsp�Xu�����mۅ��]/ �[WʔIx����ׂ':�nS�J��O�]\B��.��s�6�Tcl-.�'*�n��s1,bꆺ�Ŭ�eЫG�z����u��K��4+^����"��NY�cN���,5��qWy�_��5ϊ��K�PW�����=�oh�ăg¸d'k�H��P:��鼮���b�w?���.ם�Y+��֝ΞU����"۟����8����DQ��b��~N��:�%i�ݳG����P�]>s
9��_��F�>�Of�YH�AN�Z��$���>V��s�v�e�������̦�zbu�b�aWA5M�v���:U8�}H�������2r�;6X�ywy��{���VȮ�0K���za�����X��#1@My���R�һT4���}����t�:+\o�v�Ӽ[T�
��N�+�k���ĵ���gN�}�^1�Sd��Z���%ƽ��G,z��������Ԏ�Ow�8�q����if�Ey �|��r���������/;e�PZ������&�H�S7���r�W��|�d!�~��	�����Lɘ�E�]��j�֬fV�?s	X�+%[�[���}C_�|���O/
��0b~_@��K.�[i'z ���=�
�'������,�`x�hl[�N��R��[���c�9�}���nª2#��[�=��q�D:L��1MO������>�0�\�2�g��B7f)j��/�v뗗��G����8s/f�ޗ�Edb[�}}�0]��`:�����pX�)���g>��+�m�tB��L@4�Q~�A��g�EO�D��r4�1s�p�9�9V�m<�r�����0C��<nk`ۨs�1T)z��7a����T��ݨ�c-����a_�Q9�nʷt(���q�o�K5Fx��E잞��B�U#��\�od����j�_^&�v��W���)qc�=�3��� 9�L�~�0��N���̄�>C-#�#���N�*U�컏��ب>n��/"�&3�>hK�'�6��
Xx�)b��xT�49j�;U���F�Ϯ���+�C����X7ǵf4n�z��_�RG��+ Iiu��U��s[/+�N�ag�h+�V�����U��Y7�.��ܳQ���^w����*��П��b��Y�R��_��M
�f9�=��۹4z�
{;e��N�9�k
J�D����B!��
6C[�3�~J_�|o�:���ih��z�ZP�Y.#�o�O\��N�^�wX���#v�3|hX�rcƕ(�|�!�*(�ۊ�fFg*X��oԷb���*Jo& S��N-��=ύy�`��#�1��s��p��8҅�8^]�����?�-���may��RE�L���O�yC��S˝����[��˕��_��⁁���&������������%~�&"G5��钗1�Բw�l��̣/�^�m�x|�Ǻ��<t$͚����U��_�q�>�[�6��=D�}� ��%b���B��Θ�����#�O�ڒ��<�(ڼ'��c<;ď�6F�aE�Q����a>ۦ�/͝�uPq6�ܘ9����Xش#��B�%��%�:9؟,U�����}f��@�P�f҈vU�;n����t:����G̓���U�f�*�d���3��/��
��#�&2	P�dUH�
!PԂ%c���;<f���e�Xԙ�U"��:��w˸�b�Q#���ޗ�ԉp�X�p��{՜^壡^I�̣�7Aޕ�3'#�m�j�|Fӗu�l�|���!����Օk��)q]6�e�`��]��[q>v_6V_U�%9����n�Ӡ�L�v�g1�-�1L��83���J�mi�7p*�׬-ɘ�*\�
{�S�L}��uG;�Sl�>�����2Dޯp��8�T]qnhw\����
��q�+	u�^�>�йH��|E6689՜2�IFT0��/(2xw\�SOR	�sn���O,ҝ�zF��u��p�G ]ä����<�>��amX����~�/�9q:���Z��p!״��E�s��Έ��7� ��y����:�r�_K�l�+�%���>�ht�����	k|�zo��I��W#�[���ݑ�@��m;n�����q��i��{��R����Q�(03؞��9��Az���j(��6�R'�.�%Mµ%�~��ĳ�֮P�䍊$ꈓ�nC�����L�E�^��P�/39:���%�.�4kY̤$1Ӳ`i�8c��\z4�[��]Y�/\ܨsb�lr)D)�El��[�gkC�睻��9��Ư��:ͬ�>�.&=���-�ð�jjoqٌe�n�|����,��_z�CW:�C����\N/��m��)����
����:ќ�u�����-p�nD�Xɓ�[�8fM��q���-w��$����P�k���So�hnv^�Wã�Rɍ��/���LEh���q3Țo�{U�m��Vü�ո���r`,l�z|��F�<��=o_|2)_� Jn�"���hVt2qӦ�����f�H��4����މD%PΈ���;3������rYn^��;��r�q�K �N���B�M���͢����4�Y�lT)�Ѻ]��ҝ����W��\ͻ�H*ܰ��Ul�s:�6��(�V�Ë�Z���\[�N��\�8����J�n5u1R��+�p[���yv��Q�ժ�)Ԫ86LeTCr8�U�o ]V��8��YZ�syCޭ׫�Fk����Hc����N�gycP#- %N��ַs1p3%�c���6+̝k.�N�2A1�D>�����\�{j�`��:&]�Ζ��ꋣTW3D[/�e�x����joZ�L�D�	u˚��m7W37l�9B��i��,�C��~9�0k1(z������m��y}�y�ei�u8�f�6�H���L�x���MUq�J��_Ld��h�~��9����+��ls�1f����_���LO�v�6@��@9|��iow���3[��Ov���0hE��U��7�%ù�ʄ�]�U�t��eoe������:�t�F��u(v\���3�؉xN�J؝>�1MnpZVӗ�Γ������[8�Q��֭�a�F"�E�,c�Y*%�E
�#�����2,K��@QH��
�T#F��emKE��QU�%�Q[h�E�DY[E���X���@UF*��0UQlYZ#(
�"1ZՑV*����b�[h((�� �ETEAEEX�+J�+D-��ee`Ĉ �V*��¡[h�����DE%j�"���*"�-��[V(#+U������lb�EF
Ub�TE�(���E*2�m�AV-h��*��UQ#l�P����U,@bj0��AQҵ��Ȉ��lDE���i���Kh�j��b��b�D�����(�J��
2�EQE(1U�"
aV"��5��"Ȫ"�"R(���KlU�((�+(������TP�(�#��r��w��?�w�o���S	̫
����{9y��^c>ѓ}���_Ϟ��5:�8L4��(�q�c������ׯ�ۖ�]����ɘ���d*Tr�P`��`��v����l5	���}u��7v��o1����ޖ'�@�l�Lpx�T+�S5��חo����sV'�9s���ylF����Ȏt�����3�~4��'�ޛ�;&
��_����6MD���.��Ø�¢����j���*q1�k�WK�dZ��(b�@���TF�D���r�dE���|��?4Z�6�(�k!�G�CQɞR��X��X�q'�^���^���Wݼ���7�'�%�;>zDT��+��Ed�4�\���mK��ˎ�#˵���X����R�����@a�f*���C�R4l�=��!����l�.�0�xD��W,[�f�>�,�zLFRA�k�2���QPoq�9��D�+�-���Η�|�i����f[�M&*�`�x�ܴ:�' 7>�����][ٞ��Q�5`ծ���]��~��K}��)X�2p5d\�]bb�m��ɞ19y#���h���p9�$�?$�ANq����W�ֺ��d���Mqp�M�͸QkJ��}���ٳo��:Ow��(�i.�n28��©FZ1�}3�����)3�y��	]�R;_@g@FӺ9SI<�1JO����۽��YP2+�}�P��ܣ_TC��D�Nf�q�hH��7�����M2�O=��$���}���D�[�����
�^K;@ �;�3�ʤ���s�7�R��.�b�v�{�6'Z�q�>ː��c(A�
!�>q��)�=���v"�.c�ɓ�XB����Gt6����6m�k���q�q�r�''a,���Z�.�����Y������^+��읟d�ȿ6*�l3@�'�¿d����Bڽw��^w.��1�x��*����;ݲ� �6vw(G�j^#H�a�.��e�B�uvW�5VS�����jqt7�z��:5O�����et��[\�D���!W�@[���E���{f�.�s�V��k���edA�>.aKs�lڐ}��m��Ԃ��Ĥt��3'#&����T���z��C��\��܆�W�\hV�#M�C/�w���9�X{<�+i�k=�����q%�����Y}�iS��A�b�d'��G����g���[�Ƣ���ǅ�UoI��BeԳ�8�P+��{���tv�z��:Ƿ�%��X�C��(�\<���p��ʕ��\%TWn5�FѼ��zO7���d�����]Ã��{�ae�Ly���șhm]�Tf��]d��!Y����k�o(�[�oR̽�����Q�"�>��c�8Dl��t@"M(��=�`�r��U�����xn�gF�=J���ӹp�g/ܝ��=�`�f ���Q��=�V����P�Bz}��ܧ<Z%������+H�̫]�7!ۚ0�΃6U8�(R�n��`u�ɦ����M�7}���d��F��0J�����q���qb��y1��&�..��ݛ�k]���߳��\a�Nu_,��O��Ɂ2Da-��D� d#��ܙ��|�)Uu�/#�h�=�����g�D0;�丱�;���F��cb���e"�K�,o�Tt�;+�����z�ɟ0�1�M����Ϣ*(=�$3Cb�v�Y֭�K}�R���\�%�on����{G�|.�����]�%�s�F��P��I����ğ2�4�v�j3�h�^M7��8�k�����J��|e�S�p�
`g�:���yFׅMF]�ֹ�1�`�=��P^���������h|O��~G�8��=�{�ż=��4"���	h�m�f˓K7<��(p�볃6W�:	�0d�^��',��ݾ2���a�^Wx�]���n��'�Z���9�8iު׷R�;�g�z�g��H�Ĉ>1�n�0��bec��g#�J
���F�ۊ�/�-��ٜo��.w/�ޭ�#XJ75�m�9����E���>���C˿>�=�#��wf'�[q-�.:/�C���+7"g��8A�'��k���H��'�3m�i7kXu�f�A��'�^l�zv�����k������:��a[+�+i\W�/�]�d�����pM�)=ڽ^�خ�Ȟ�ۚQ�.6f�6x�l]���<�_g���#�9v.�4�ذ�Ӱ�AYJ-ә#�A����6�����ݪ�yT�gq�C���pp�Cs�#`���Hݸ�L�c�4�D��!��YX��h��I�=�1s^{^!Ωѓ)Nd�/���z�j�G7Zf/m=�Ò�bݍ��=�P��Q19�F�_2(����1�0E�z�a�d�?;z߾uI�s�q|(epa�!CdE��H�|JB�뎍�~�,����?R#�{F��e'LĕV9�W�N|����9�U��%1�� �&l׬I��U��_�q�&�TQam譪�C�)�CB݇g����/'Mlt���f�͗w|`�)������"ͫݿI���n��Q��]9xs9up�#tM���k0��W��U;\m��&˔��wt���8�3����M�=Ǵ=y)��G}f�7{6)�
�)3���� ���[!�;�<���
��D��~�+zxj��#P��^�wG�eW�5��{���+3f.M��	�?eS���0��nb���j��H��7��I��O�<���X݂�yJ77s}���C�!��ب��d�Bm(�e^C�����]���gb��T��#�M����;����7T /V��=E���ـ_3�1'�(jA�������-o�w�U�^}�-:3o'��z�����*a��.�|"�Ƕ)CzB
hf�<ݵ1S����Y�	���䶖ǘ���N	u�+���>v:}9���ǪQ�A�7�B��)}�rĲb�;��?
O�!oϸ���+�|�֬,��_��l�aM� 6�('7�����'U�����Z�����'b
�Щq��}O�\��'��؄�q�E����l��nuU�v�ѼI%�#e��\At�w&܅Md7�uj93�sPV#eS�q7��jW&�b7��1�̳$7U�'iP&t�\뜹�X'!�Z����2�ө����V/#��x��n%t(��Y�GW��P��J�W{�!���*�}���Ѹ���&��%�ʮbU+�[�M�1:z�=S4o�	h���S3�e}\�˘�}wO��l���[�EEX����k=�k;��tigRN������ڽ҇ZV��l¼K��� Y؞b�8��hl����缅�DŘ��g�%R�Nz���s)�,j���??T�hcX�q�D��N0{�bϨ )K�Y�~�5�l�v�˙l��y�z3�g*1�@�
P��
Y�͞�3`�	,.<�M�C��l�}���\)Ţ�Z��kp���d��\��"��sT "�69�F��d]����\��uNwV�%s�����m�P:)ȸ�nr����'q|� �jH|*`��m�@�fk�72k�v�(Z����XB2�:EeI�P�,�.����x�+���|�������y�&���u^�cS���3Ǳփ=Fa�.�0�BQ��ѫ��δc6�H����,GE�F+1���Q�>���[�!Ga�0� �GvDR�\*�ev�Fw!�()`��������yt
X��~lU��4a��W��W�����Pc[��Ǒ�XΨ�~t�el���=�2t%II"��R�y#`�&ڡ鲎�|m)���D^*�$��bL����1�ݼ{3*;���^+vo�Fٞ���R��{���U}�ܴ��C�4y��x9G��S��n�:�a��(����K�G�D�ƁM��ǔg$�7u�4�.`_.���`W���b"�����s���"�C��bGj�3�ݸX2�^z$tmm_�R�x+�)�m!qn���M�iNyt��~�Y}h���R��#�Q��-.�'*���,#��Y��ŋ2�lpթ�Q�,&��L@�C�I*,V�"TلP�rοA���ia���λ��/�c:̰����r\I�!EZ	��\C���鼬R�^?pKn;�'b�`�s���u���ޙZ����F?K��"6Q�����Q�eEc�b�jԊ�
�C��A(�:í�j�硖r�����T�hE�����Z6�#'7/�h��wuyoZ#��T܁�+F�e���&������:�*�H4�Q�T��v�ip���Z9ǥ@u1�@�"��*O�K�����1C��
��<���b���4����Tn=���\)��`M�sQy;��5�(p���MB@r;�0�d��a�)Iс�
sS�6X�� Щ!����_'�1y�7��a�~����l�/�1�Wj��X��׳/ll-݌��-Y�!�[��d�]�K2�}C�@��N3ɜϦMN�xzf���n�&��q��ٽx�ڳi�����BQ;�&&ѻnȧ�g�rH촙Ü�M��h�	.ſL��i�6-ҋ1ԕ���\����9�Y�Y��[�q���GG�4��\cd��;N�0�NT�46-����­��{i��zNya�;���7vX����R����ʝ�d
���t.����>�v�v�g�σ�O�7���>��q(�W�1{I�A�� ��#p{�_Gn��R*�$���&x�g ��'��w�U�w$F)�,�y5���)D9ޖ m$TX�=���h�+iL��35�^s̶aNx�@T��>ߦM�Qp;%�\�����U
^��nÈy����x��Lg���b������ҥx�<h���P�~'L�����E잞��$oe.Z���b"�Z��^�T�`6E��|v
�'�A�
\Xd=����1� 15��>x{�W���v���߱+��L��6!ǵ�Q�r�jz��4�3�?x=�I��'��,��X����I�F>S���*Ʃk�[ylXV'a܂R�Bn����Q�Lt�~�d�4Eu�;ť��*Q/�h���a���.F�WCaב�qؙ�5�sQ��D��p�-�����j�f��9�p�p�e�YN	v�,d��R�Z���58ئ�z�4���<�*1�An�ѷ���MtmLtGZ�{&�iq-���<tv�;�2�n�R�cjw���>��7�՞��ݤ'SF�gn��3�׭6'l�x=��YK����[0:T]L\׻k�9�;영JNe8��Ϫ:��l�s嶟�]P����;KL���C���^���j6h_"*��{}�AAɊ���v{�lX/�J��/h����#�ˌ��s�ux�`ha�t����ϭ��Ճ�̊ډ���=V����V�lf�r舀�t#�����S1�aO�"k�E!'�A�f�z���],�|�W'*Y1��l�m��s/S��G�X6a�I={o�&��ţ�,F�:��4�rCԶ��V.���,�>"�N��0��nb�; �TI��5�z[^�P�=���f7N�;�H��P��5qCڬʏ��^<�|O���g���Æ��1�3��n�������vj)�B���P Et�ȱS����f}|ϔ�z ���Gb�#�lr��&�f����To��v^������ņŝ�eg�ǲ=��C�rD�%M$���)? T�h,���)�,�a�>�}y���ݽ��>������� ��:�=��:�E ��3(m:�p�q��X�)�{��C��W���&�Y���)ϨIߏo!�aQdٛ�aP�'�w�q,�%C����\{�1˜��m%$׸2bt3.M����Ӕr1ف4u�w;,L��](�1L��ԛ|֪U�6nڄ3+�@�
����˦%�;bC�Z��t��dȝ<V��u�����S1�kc\$�MO�uJ�Y/���t�^ou^����{��ɡP����L!��Sy6{�xo�J9���x�����=fRi����b��+0�)���u�Y�Ǩy�O�Qd�ĩ�O�/P�;���׽�톒��L����=�>�L�=17�Ø3r�/�Q�_˕zC�&�m��,?0�=�`ز~�u&�\�(��8���	8�N';�C��!Xq=�̼d�w6��<�_̚��)��<}�*̤߾X�vM�g}���������$D7�}�j����a��l0�mJ�똆��y |�Va�Y��8����{�q&�P�g�p~p���f�s��d�3��~�u���Mv0Aa��Gw�����>����"�y���S��T~p�yM�XOY�0�;�AfX=���c�y�C�y3L����fS�P�Cv���S,��L (���<�y�ݜߝ\}������Mꁄ<{<�a�4P��0a�0�����g�*j}�

/�N��I��b���1�B�����q�S���J��'�O�/���0�w{)XNg��:鿟��� ޿�>��C��w؆�L��*O~�d��2���'���e��ɖaP���Psb���̨(
)�M��i:�Re
����>�*��c�n�Ns���ߵ�����nY2��d�++%zɜS��0AO�L�g�f�l;l=��
��s�=��ef���쁔X�\�?!�0�X�:���gP�7)h|��u���/�ϵ�}�Z�Z�߸g�Y0����~�2��i��̛̳Ǳs�,+
̲{���P0��S,�{��T��a����y�8Hl�� �)�k�Ğ� �i�>�SHq
����;�����9���Ƶ�o�~�����f�m9`]�+x��y������
�zɄ������P0�~�����)���aXT<̇����`Va&��i�Ms� �M!�X~��r����Oۿ�ޤ���R<&<�:�\��b��3��$ㄟ��ϳd�m��4o� �@�ްi��a���ݲe+:�+2}a�Y<ʞE5?s��!Y:�1�\��L0�
�������hY{���~/���8U-r��x���kq����ĕf��mL8�ڬ]����E�O!�����{Ջb�M���-w�����5m�r�D���D%Ʒ#^����&u�Nt5��o�	Y�Ǳط�X~_5ϧ������׍��zzt.�~䯷FZ ��vi��%���1nl7�I�6LlK�N��I4L�a����փ�[���mx̾���7r83�o>o�4U��.�����%9���Ƀ��c�K���?p����L�Me�y�t9����Y�R�R��@q��ۣ�U�Oˬ����^-��m�G��}wv���|��q���B�;I:�w�2K0��ٽT�>�������1�T��)�'[�����!��Z��hM���2��2��`b^��;XRR�x٤�g_ܲ�N&^�]�����9Uvs5��Bjh|t��sk
ʵ<x�y	۫�˝�9��z9$�:1�"+���HU�7�:�QdM�'ϋ/�]|���*�����6��j#Ѽ�ɖps77W*M��b���Y%��ʢGJ\�CY�d�{I�6�luu�m\�.�:��iZ���>:�$p���݁7��') /n�w&��=�F�@}�x,��nb�:a��VȤ�^
m���@�1}��d�X|�Y4RҘ�3>��ɦ��nvV:wEW��U8������;-@_{|�b��\��:ұj�O��zۖS����'yA;]-��ّ�@oZ��t��˼6���Y-)�Qs�%�z���㉚u�yH�gU`�����xwi3B�#k4S3�.�@�� {=V��=ހ�w��N��%�i2�;� Uʷ��z��m�|\��權����xߣ�"�΁�MN����`eHyM�t�~�c���=�ׯ7)��m��vq_|w2�Z�ͮ�O<� �(.?f����A�
�ζ(�&��V-�/�+�9��VQ����rYIў;�9�����F�쨩-o��H���}�e�^��̈��,��^E����ݝ{e�s���yB�*��R�U�u���\ܥqQx#&�<}����U��c�k�.�����`wK^Ǡl��b�8�&5$�}`���Y��z,�<�����j�D�bs(ͪQ�V�C^��R]���,GU��U�>����b�m��U^�'2�;���,7�	؊�����g�;�qs��[̒��!�N��ˤン�8����ʙ���VZ��!/D�%�-��%m��O\Z� �B�%�ȹ
��R��vf4�K�{�]����0��Ƽ�n-0ݧ�v:��� �hFs]8�f3EĈ��mw�������a��z�{��$3������yp8i�ˢd����#�A��ώ�4�ٝ�7ꖃ�������ܥk�j�;�ӆ��ib���;tO�l����6��xZq�,��<��AE�q�����VM�6f�/��϶c���:�*4�	K��[:��[���Q�*��#EŤQUdU�(�,�Ȣ��Q-�R(���FҢ�1QPYQF�R"
�aR�bȬAU���QUV1QAE�-�6؈((,��EdEb���Db�F,EAA��QTdF1AEV1b*(#QEX��,�X��X*�,Q�#U"��"*�%k*��Ƞ�1Em�DPb�AU�P��ň��E`��`1X�UR,Y��ZTX���,Y(�`��#dDQ*��X�+X�UF0X�EX�V��őQ�(�H�TA���(�UQ
��V"�!i*�0EUUb(��F#"*EQAUEA�
*0A�
�ł��UEEEU`����dUEUPQDT�(��"����AY���m���b����*�(�m�PEb ���H�UE@X��AE-�PV" �X���*0U��YEX�0EEC��cY����ː��W@��:¤��6;��G�o�Y�+9r��=�&�"e��2ͩ�M����{&�m.]?�����IR�~��y���a���2��&PS?����L T���3��q�i
���N0��O�ٰ��3���&��Y�� ky0N�*A���'�a�B�Դ��&=1�s��l� g쏕#���[��>2����_��3�6�!�!�����"̺7���2�G��5>d��{�Ra˔!�ӈe��7��L�>aY�N���:�Q�G�""�@��7�qč����y"�|�Af\ zr��HW�,�csW7i�9ϳ����E'���2�a�a'���yd�^�i�R�;=�
f�Y0�~���L*}�&S� ��1�.E��L��X'���ۻ���a�s����Y�6��

/X�g�
�Hs��13\�+�f�'�?b��{�,�N�I����a8ɇ��`^�R);� ǂ������q���ҕ��K����:��*JᒢɶT��&�e'��߱3l�&q��I�Hr�_�Y2���f�{�i�
���>��u��=H4��
�ɔ�6s�L1G�1P�u�\�M@��Y����!H)�'����eH>��� sv*�3d�l�����PXMwJΰ�y!���ì0�p�z�)Z�������&G}��ԕ�� �)�Qp"�XUgoa.�%��4ϙ5�b1�B��³d���7�:ɹ�k%IUR
u���E8�Ϝ0��B�Af��Hr���&P��E��d�i�Y�?'}C))��]����ܻ��Ԟ|��Y��ؘa����;�C�i�jɄ7�`2�0��Xl�14��VCF=�h�VaS;�'�Z���{6AAE�'�S�&P��s'�^��Q�����H��I�A�0���.�4'�{���y�Yęp��sJ�Sl�p�9�_!Rhl�0M���$���ꁴ�Ұ��PY+*~>�I��B���E����:�������m!�k9�d�
)���7�߽�'�k���}�{�]�I���X{�C	�O8�|�Xq�xɴ�~�Ha�d��^�!�����>VT�}��R�a�B��� wV����(iE&w�E�V~a��3������7ӨY�ˎ�V��<2�-���s���Y&*�mm��볺�ÛH]K(���MG�HqI�b��+�t��A�L
���١n�[+1�q24�Ěהo&8
}s�ͮ�a �f�N�� �7�]m�ϊԒؖ����  f�����ַ��{��|�	�gT�m��pL�N�a�TP�%p���X%B�̚ǰl�,8³I�g8���Y��0e4����O i? �N���L���[�����h��]����5���|)����~��m�S~B���	X|�!�~��4�sd�o8�4�a���)<�f�d�l��,0§�f�,4��Xe3�bk�P+��1��b�f�o��Mw�3�o��������6����=>�!��I��ϰ:�~e�![�a�Rmb�Ƭ�g�?8I���e��dɯ��� ��ɔ�z�|��%gU���@Qd�|\w��{��{�s=����r��M"���;��6ϙ0���T� �&}�G6a��)�w9+'�	�
��g�O̟�z���2��������2W���&�E �_�0$겤�;�{�ƹ�k}�����?{���Ԇqa�g���$-�<�_��,�@QCS��8�+?0�i;9�M��2��TYXT�-7���&Y0�A�be?$��0�2���2~��wD+�+?x����=g:�x��߹���_{�}'��,��v�SI*�C�a4�S�,뇽�1�!_3�;��ɴ�m&���,��e
������a�a?z�6�R���E�.G�G�|#� L{r}�|w�ʷ�~D��GSX�Y "G�G��o( `{`������a���L�ԞŬ����AAE�k=ĚM�T��?d;�'y@�s�4���&��.�� ,���;�L��S����񿩾���F{�~�;�ҽ`�B�=�a�I�j�	�P>�IY��I�O��L�QIRq�d�-�̘N~��2��6�Y�!�Y�J����"�d��? _���:����q�>���o=�0<ۼ[���{|�}'e�p�����H,�������oR�^ dI�eC�iRbî�$?[]�eg���s�'\�gXa<͟���A݇�޳H��*C����z�.k˖�x��q��������q%'0�Lw�(q%r�=�Ci:�fh߰]w+��˜'>�,���2i6����T�M �f=��yHW3]�,�i!�C�J̰�a2�Mgﻏ��u��V��Ի�m0��t�ޒ�����f������iָM/��h�ɷČه�؈JQ�ކ�0�ߎi��;��.:E[�Β~tW��F^o��g�1?u��}F˷�Ms���d����$��U�_L��䈎���F�m�	9�ONu�4�/���!�Z��W�W��a�}^��t�%H)���籴:�C	�߽�i�6�a�Ǳj�����2�XV���K�y
�f�r�a�Lg0�q'ص�S4�:�PQ�2��#��~�ɯ��
j��[��vu�ɖ]�zn�Xm�qI�y�i�I�Nc� �G�bv�r�d��bg��k�;nR�%O�UI��þ��N"����O���3�z�������8�}}��	��C,��,��'Y�&f�:��8���|�׮�I>I�3?s�V���d�!�o�&�{@�B����G�q��Mk�a&w��e��f��	�+8��9�5+>a�ٝ�8���Xay�@�>��C��y�o0����y�)?!Y�d�߰B��>�i�d泂
�O2a2�b ꏻ���0o��vz~�������}�f.���r�q0��42��a�?`�H)�/�2���Hn}�V,�u�G��I�+7�i�R3�sOz���B�����~�N�Ņ��#��:Џ�.</TP+==��i$�-a�Y�,�%AC3���*u�톐��'̾���aX}�N���e&��I�*AM�'�,�T5�&-)���)��1/����;��R������V����k3���k��q�>E%a��Y>e�e�����aRa�g����Jˋ&�M8N�����>d���ש
�,+��m;�A}q���c���j�r��~pc�0*=�OY��I�L�� �C��d�1<�i!�a���<镟��&öa��R�=�`�a$ٳ����,�
�X�!�C��y�S)����k]��	[j.�3w�-��z�	�}�Ro]�
�N�P�4��g7ˆ|�SL�]NXJ�S��}�,󴃫';f_ ��a����� �L2�M^`RT��f}�4���d�0���ӟc���~�߾������%b�'�<d�7i>B�&��ɤ��x��{�$�?~�Xi��
����I�Z�=�I�~d�)���e��5�cI6�زi��������4�~�J���Oe�a���o/qx�h��n�-�V��݉x��������dӖ>Z�֟��늽�������{m�:yβ�k\��z��v;ݔ��V���z�)M똰��|�g��Y����B�Vax�yS�����; �l�����_������u��� ��^QjM�E!�C��O̟�0]!S�S>/��a!��hްe�T�O��̩�RV~>��d�-���k����I�߽�:�?[?2WXιk\�~#A�w�`w�%��P"G�b�d�I�2���E�ԅa�6s�ӆM�sH)��q�7�(nf�	�u�񉔃���c�!�B�>����Y�0���0��Jβ�����sܹ�ؽ�>���;�S�~C	�=���E��V};�I�P�J�8Ͻ��P�fwx4�hI�
���,����l���f�?o8'�T0βT�J�� ��
��g�$P���u�����`���w��{����@'�C?}�j�3H,�&��y�QH)���ì�'P��r�X�)���4��i0�}=��M (�Gs�a���$���CL6���ɼܰ�
��=�þ�Or�"��N�;ֳ7y)��{�ޘ��(�`T���a&P�,���+�B�����P���O�}��J�&��J�d�����rA�	�{�{a��-�sb�g%@y׻�]�*�|������Iw���q遰��l:�Y>e�h�q&�u�I�� ��l�O�S̜p�?^�e'�����n)
É�~���O���>Ǳ�y��d�(��q��w�U�����*`���o;��"#���ޟ{Շ�B�;��֠u������"��R�:�!��C�S��"ΰ��X��W�ﻉ4���'��4��	8͝�y�x�W�9�|��{���׾��c>��?2k��x9�,�%L0��8UR
y&�����$�g��4���73a��4�W�2���4s4�����a�d����2�y�H}i�l��C/���OaU���k/�q���� (����}���0y
�L.h��w�aP��Z���%Mc����S��4�IP�,����+0����8�qH)��T����TXoW������}}�o���:�dˆ�=�e ���ƌ�0��6����6�g�IRo߰eO̩�P�;������Y2ì*�p(9�>�y�1A@QM�k��I�C�=���~9��J��)�پ׵�-���f�0�i���.�e`�Y��|f�;��)�{9v 3��A��l�W���J�~c�����!�p�@��f#�'Dݨ�;o�]�1������1��`����']���yp�Ϫ�Ͼ�|>p�ն�/[���QnG��"<&:=�����+%|ɬS��S����fRl9l=��
��{�`q����ײQ`V�s��XT����>M ��a�2	���5����߳+�k��������B��W��8Ʉ3s˧�I�g�e�d�;�9r°��'��@���0ϻ�M*���&S�,��C|�\���e0��^��#�#�,�n�D�{J���_-:��E0���x��S,:�!��?j���Jř��q������Vk�L .��a�=���!�a{E7�L��*gݳڵ�Y��}�	 �N�DXl�Y7�.0S��w��r�:e��Ӟ��8�+'}c�N!�R�s�Ĝp��TY�l�M�|ᆃx�P���L���0�տ��)Y�IY�
�'�Sȧ߹��l1�8��<�>��}Bl�\w�V]�5����i�2¾��!�R�e�;�iE0�>��a������J��g=�8�/6�͆XV~d��M�8��@Ἐ'U� �f��z���@��>���O
�������V��YY���mE�ƺ���3�6�!�!�/�K�0�,˩�`4�ݡ�=�i��&SS���˧(CGu��i�d�ęf~aY�O����:�SX?gǮ�|{�x~�m�ڽ����3�uU �����S�,�}L~�+�u1��դns�fM��
�O���e6Ì�N'�� ��X���6�I��{�Y��L$��`�,4§ڲ}Ͽu�?^�JGռ#37{��`{�	������*���`Vu���

/X>��&��)�\�8�r��7c�ø����P>;�gRu�M%G~��N2a�4{�T��O��s���T!����#��|�g� lx7>஺�J�ʒ��aO�S��I��B�|oؙ�y�8���):�iZh�zɔ�5{�i�
���}���'z����8¿�2��g>�z���*_UE��N��r���=��LT�������k���8���Gu�݇ʅf��9�河[�H
,��2��a��C߬nì0�k���5h~fÿ�4�2Ʉ���{�����>�7��ג�gU�3)& GY�46�O;/�-G[Eb��v���\�=l����E�<hP޸�8��c���ܕ�k��%9�@]/���VoL�X�M��aj��S���5]}����I�=�*7�'��c��<J�ۆP�dvɰ����ﾯ�����W߳�w�}����Wo�O�c�!�q�X�!��1
Ì+0�~�#���βl������:��q"�Ag�k6�!]��D�0i!�H.��L8�C�lՓ	�f���8��K�{�ޞ��~{���>$Y*w�~L0�C�����u3�Y0�}C��
���!�bi'��0���[E��
�&��I�V�+:��� ���ɠ��I�3y������f7����5��ucH���sz4���|xvH��R'�C�N�I�`�AO̟�:���T��=��l?j�	7��ꁴ�Ұ��PY+*~>�I��B��{���?2a�SSz��O�5��{x:
��S=E���~U3s���%@QO^�O8N�V*>d�P?&~a_̚N�X!Y���O{X�ۢ�S�w�2$�YP?o�3�C�,2�Ws]����Y]� (�!��Gc3�_Vsi��c�N��x��A�0�d�1:¤5hh1�	���L2l�E�W/P5��J�g�5�`��Xq�f�����<���0e4���s�<�������ڟ����fVk��_��G��@ϰ)���_��,�&��E�́��>f��u��>��"�'Xa���O!Y��0��"�0��Y�IP�0�9�Mz�a�ǽ��a7۱x>س�R�=u3c�}�$�

.�y�i<�Rm7��ud���B���L9�O��,�%f�|�'��`�)0ɯ�,�T�����I�����H⁔��Wz�����:o.f؆sv��h��� ���Lo�͡�hh��g�'�1y�7�]����g�Y��FmF�P�7-��D�}%K7�B��s�	�o��eϢ2�α�߽�Nϖ�[�$�!cԘp�l�:{��Z����c��ǲ*s�V�P�~�hZ�3<�53�����r�q�޼��:�*<}�&aͣіtU��T�EC��<w�^��#8l�W�c�)@��L��mU��1Cf�-xkᎁ��<���N��z�\ ����1!w5��s���u�.�HoB��;RyDX�D�UjLS̝>S:�H]�#<���������ky�>&�+����=4���r�?y���}(���ӹ��\7AB����ǯ3��yf��|�O���2�gߎQ�~5��mq>[��}Ӎ�{L%��o/k]�N��_e�Q:��a2�O�عG#>!��,@�q;j�ώ*�.���ryC�1J��t�㻇9���/S�9x\k�r6+{�ډ6�P$u�[�G��B|�F�'�z-Z3�ݢ$	a�ݑ��׉]�Jj�Y��u#�2-�/l�:�)�`{�������m�"�Nr��x�X��V��s��~�u�����K�q{�*�d��0�z�؞���e��Q�o��q�M%�#\ӌm�A�e\��r��� rذ�Ӱȭ��u�U���|���K4
���3���4���K�נ�:�jϼ�RH�z�q����r�Wp�3�R�V<J�c������yӭ�s#���Qt�-��Y�D��w�oƽ�u���J���(�MOA��SUbU�a��q���TB����ƣf�P��.<G�m��Q�һ��dcj,@���n� ��YK��i0oFEf�"f1�YY�i��O��o"�q�0�y���c�6!�c�p�gi���J�5��%Ӳ]��[bWk<7e6�[���eR�CLP��ŋ;Mڥs=�����V�!�r���Wר����� x����z�\L����T�{<���&�+<ո��a�	�t��j��Y�z��|0N~��\��Ἵ�/�år�@��!M�0T)tmq��[���BOp��$͚��N�o�M���)������ȼ�.��j��I��~�(oO^�A���??��/�nR��LHW{)dʫ�z�#UK��+�1F˪��%�W�c���e?yl����6��9p$���TfM�<��_O^z��Ƽ=���x!���!��I�� �4���͕�����L��u��w�R�����5�h�!�?}^�_���T؅��B�j��)1�z��^���;�]�=#�&NU�(����N�wH2�X��������
��g�v,2���xP`������1y
u$/<&��NOR�ԽB�p�O+a�/�ث��]��w�0|�#��B�%g���5�]���MjfM���Ȟ��a�t\���zv���T�H��7}q�!pSC�Hl#�T�`��m�1�o"�r�8Iq�|��0
٦W����?��g=;@s�G`�M�v��؇�ʣn��{����i�-��|���2�L��:��k0@s�~�F�cڟ�c8����z�2�lG�ez��Oot����#t�	|;�}�>�kJ,��֒<��hEt��נ��Om���CD��q�]3�n��I}�r�
�¬LT'���=��<<�h]�ov�@�?P���R�������*�\�����t�XΖ���O3T�h�T����zm3�Ε5�o�LWB1�z-c�$��>�<��!�oX�i�x��ă��c�2�|���(QQ%�bd��UA����C�Rv��:��7�u\%��gSP+j�R44����������,E���	�w�ϩC1�'�%k�x�����sա�_����2�ޫوfH���+�R��l�A�.�DW��(I�ݤvT��cW�N>z��5�l�,��[��[�.����?U�����ɱ΢4T�7/���|��j�O�a^*�qY��3��9	��}�Yn5��/�D�[~��Gz$�-`y]�N��
5%�S�h����j�O�qI�(k��dx�y�[�<#��bW?�y]�ߧ�5Wh��7����#��u3�zl��ȴ���ߖ���G5�S�z�}�������h@���5ߜE���8��G���7Qk����6m��r5����b������NJ��R���vnv�TClM��V:
����Е��K{����Z�f͑���	��\���wK8�=q���Y����v�?�ş5Ñ�m-��dz.�ۮ�Ѭ����E}�c��Vo�����RyQ��DW��������:ڛ�R����X|9W�Qv����9֩���!��S"�{<.Mm��ܫ䙬<��:q���z��+ބ�`s��j�7f�J�f%ݝ�n��@=���w<xg�`���^oMB��}�K�_l�G���JOL���i��>m������ۺ¹�+#;���ًŕ������ƪ��>U��G�_��"��*�Ks�lڑ�2����Q	١`�4���+
��=��x��3X�XW�L@�2H�J�_�l����Mcr�E���x��ԭT6�ɝ�Z����jK�2������H��K�bᘉ���en�{mt�I[�}�7�
��z��)��ʜ~}w�mj7X�DP��pa����Ʀ����>��oU���W�KUiK��ҩz硐�_��L�mS١
FbZ��"�u��kc8�����,Tj�� 6�Ը�>V��@�e��|װk�����9� CĮ�1;���p�N9b/	���'=�Z����jg�wL'�%�Sq���O�9�ĵ�H2�����R�M�xf����"��u)���`�
�>�ɧ@����U�|r8����f���$�(�t۽daDƽ?%B��"���$.G��S�7�b�u��Jn�pY�B�|���wK]�9�ȣN�?`[6�u��ˈ�7�#�)����o���v�����%��&��M;�+U�,�K�۾v��w�l�tBqx�c	o���8�ʆTG9�3g�� ���vD�w�*��+z6�.ƨ5g4(��͛ʹr(ܔ`�و�Wj�Խf���*:��أw�[�u��Lgn��W��x��^Z�zد'��+G��Y/���`��jqT�g�R����Pt�ϯz�1m��ͱ�ve�m�e�5�uCB�ܕ�;f*��J6���\�WL�5���Wө,�9�U��B�+m��W�Z�=@�V%D:��E�:a�J��ԧ�R�ڵ4����f8	�(3�:T2����p�F3�k���F�z��Z�T�U�Dc&�;�vU�tE����G����xy��tw4�㱡��� n�
)���Ӈ��uѳ�����"7*mr^��&��2FGQ�gw���ۋF�-�|�J��^��ga�%>�}�Bă�V^�������������H��/l�3:�"+�V��ޝ����x��F�ԦKT��ڙsz�$���&4ҝE��|̺c��m��R�x�怚���|o.�]���|�is׉8/xT�5k��T�*љҪGQ��e��ӡ��֎vV=N)�M�u�)�C��ݔ��������PX�����w����B�r?4��WL�7��kEo�����Sw/wJ�X-��`.[���MKi�X�<�@���Mu��w7F�&���b�xieS�<���G��0x�������h:�\,��6�K�"��ƞ�':Y�1}��sx��]�@��`�F�q���*kr�[�Y�
YT��$:p�F��}\�ˮƷk�M�Rngѥkd�8;�;v�=�F#��=Z�Ulu�^���f�B�#��
�h\5n��AI����Z�)�){�(:^�|kL�7s۸Ve�rX4۪���h��c�\�� ��A�$�t��RgV�ʋ�1�J�9�T{U���վ��H�p�����di}Fɾ���+�[F]�;�U��Kw��]vs��@GIn��&�9��8j��qWNe"�k����9q
z�;n�	�N�Wb�ԙ�؝'�lo����ϒp��S2��r�#%eѻ�W��k?����:m�)�2��B�i.HXK��suY��T���`O��1q��f�+�K�oa�7.�ڶ�`w:r=�3�C1�7id��G���m!6�Y���z���8��I�I)��t��aK�ˊ����[�d�pd�V�� zX�����#3Y��2��g:�y�`UX�F*�"��Ȩ��DAAEDA�AU�(�UAEPUQcD(������Ȥb�����*(��;�X�Qb�0`�QQc"�D@X(�Tb���`��T
$cl��UE����"�"������$QEE����@U�*0UH�EDDb�
*�AV(�1X�cAX��b�#���EX�E�1QV"�-@�UQb�("
�TJ�ETPYEQH�(�"*"��������(
,PQDQD��PEbȈ�AQ����U"1b��
�Tb�*#TAUUU��U�Q�"�Q,D+X1�b"��Q��X*��UFE�(�"�"��bUTE��*

�U�V+,UU�"(����`�-
���TEPV"�-�,X�T�Q����TPDQ��PPX*������b� �����ʃ�<�9ܥ�|W:j���t��1]�eNxY�F�zx7ӹ�/����RX��{dL�z���«�.�ڳ��� N3Kt�Z�V!~��<���E�� v_��^)�͜s����QKr����Mk�x�ˠt�@��e��<ٍ��#�"({���_'�1{vrw�0����Ꮍє
=���̽�_��"�Is�z�p4����ls�����ڒ��uw	��E���ܹfTk	�8j�z�޸~v���C���o?S4-	j��]�>�F��~�<�,f��F�Z�K�\���ğ2��j��r�?y���}(���ӻεH�]��^�;�v%��3/Ɋ�>�Tٜ��0��ɯ(Go�R�rF�1 ��*8�vbŞ����bT`ܓ&��M��4E=��G��J��D8�v�e�|�_d�0I���Gf^B�ʾ��P���P}/F���i{�N+~�8�lu�G��@��7����~���Yꧺ7���x���׋!m��֙����)Ez7͘R��"�B����s8�q
/m�tL ���?�;.��_̄��O��{�ThN��j+�c��W��^��;���r��K�V�֚���piX.�7��Wo�vJ0E�)�Kíj�������hm��G�^���.E�Ly-�xX�d��:�.���[c�mf�/ɥ6x����}
��&�P<}�^e�?d�X��v��G/�O��UP��m�|����6�0A��fR���s��OM�48��C[�3m��F���yٽ��K{�g��3�y-&����U u�2��+��:���qЧX���u��c2�8��h0yC�z���=�Ѝ\i�Kq|���D����^����F�񝵑nK龮�?OB�Q
��g6t�_���Ц!CGC����DU�8 �K-��z�b�vO5"dt0�JJ�+G�x�q`���p{��C�	�t�������=�1���i5~,��ի�/�!�~�&"G@�P��hs�8���Jc��d�!��/j0�u��7��ynLt+~'��r/���n�.*=�1
�)�<����RBk��vf�7]h���J�z^p9R@�[�z��Eۯg�����2���za9�xux�a���9�&n7{�(g[���C=��t���!
6՟yY��v�xx��&5�}L� ��*u%�==�Nݪ��Zӯ</=�,�}����j؅�Ցғ|x*���강HL�*�*Y2o�2����(����M�\E�̜/���ؘ���m(�j�BP9��ʄMJ�/����^�7����$�;V�j���^����I�j���qtذ�P�	�T��$��R]Ҭ������R�񑫪귖_lV>����xot5��挘���!�2)�R�v61;=�G ���Ŷ,�X�{u�Pb��'��*H��&��{�~�Si�R�;�&��io�r��H{�M(�t��P�������Y�x�p}#�u��voUm����欠�����oޭ"���C�rcR~F�E�}g�fnvjg�b�~DV�Ut`��*ȃ�g��!��}�]���s�Gg�m�v���W�=��]��V��qJ���������z��8�TТX�=�B�rjGgް��J�B�
6�[��Άu���8��;��m�Y�T�Nׂ�F�V��b�|y��S�<�yW��k�at}aV��J�+~'!��>���3`)pb�=8�=�	��ѳ�|h�)еN��Yه���ʹ��6CAS�@�ݐ����$W7}	������P�b%
Qmz�C�	�RHڽ�]7ٚ��l&TTZT��	����C2}�6O0BP��o6x���$���I������҃:�����	��u�ɲ�;��%��U�R��K��y�t���-x|�b�I�^��a"�w+���(��Z��t)�8ࣷL��q��e�O�#.;���:���Y5[����6[�0�:e���c��\i<("~�ssdb�M֡����&kX�8X�n�5�Bu���x_r�(�MU�y�}ǟꪡ����]{�|�ɠ��1?�4�Qx�����3񜄴ϼ��=���W"��.��z;����rk"'�� dB�P{CF@=�o����,5V���\��nL\T!$���}�J�/��&~�r�\R��o�}��kρ���u��끞�>�>�����qQ�S@������G�~Pu�9��&�E��m};C�@��+bJ�`�'���<��KHؘ �t���Ђ��TCݾ�#9LS9��p�,�c+3^��R�`�JZ4a�K��V�l�ڀ�V^���M��b��ܡ
��3�N��7`�Ռ�S,9��8��8
"�gԞ��s>[_c�F�3�ރ�ۅ�e��r9]�v9�+C����4��]ϊ��'���w<��vL��*�Ks�fԂ���FtbVjB+c�ʩ�QnpKg����tM{�
����cE�x�@V�#���y���kP��BX`3%KX5VL�XZ����~R\I���Q^�4�+d�������^����w�l�ŷ,WEn�N��0-��:yOzD�[ќC ���W:���w۶�˔��i�1���ص�Aܰ���iXjl���!�wm��d������`�(>|.EܩSM�A�Γ�"�����m�[U�7�g����������{���T���S��\X27d�N|Nе�,6}^��qhC��%$�cj�4���vKk��C�ppN9w�F:3����Z��B2�z�z��]-Qr��{���|�x3��Ā�t�a�+~�~���>k�5�{�:��scV�k�&2Rb&���l��B|�N3�y֬!J��@��Ņ�*lG��/^�{��LLQE�)�*��9�8��;h��0��<j��0���ͫ�+�/����8�O��_�=
$j:gvSjdҖ�� D��w"Lއ`�=����^4ɘ���kr��㻘�%��8T����`�u�Q�Ed�,X�1
�iϓꌒw���>��z'jr^8��}nR���ϳ��	���£b����F=�P���!�ʝ�d
�����Ե�dK�{uӕ��J��ϫ�f���^�-���B3?yk�8h��Ӯa�|�j�A=cC�iE�&[��4��.1��8f�Q�c&�E��2�C���b<�[$j���{��G'�U�ɶ�!ٙ{i�:�tn_YTMV@�r��b�p< �L�P�"/)����B��3)�pISx'c˅�۽L^�J�޾�z�]~)P�?qs�v�2�`��9�fT�gq
��z��L]K�Hf��k�f���W�����kw)�zq�9ձ�A��bh�+ |TI�#O#>!����F��I�G��잏"�^v�g*�ݩ\�T��"ݧa���j����=��x�<BLvuJ?@��d����W�+�Lo���W��S]�7��)iU#��T�/��J+ѭ�R���.�+lfB��g�+��
�&v `�l��������Jo�?G���b���ܗ�Rz&'8�Jl���x���w���WI��'���R��R��a�/p��&�_�Ԃi��>�!/��[�x�"s P�1�L����b �U��|��Uc��y]!�r|q�aU-<J�s���̔����7>^`/6g،�*b�kĈu�o�1���Y���v���<�(�ZşUzT5./���͝3�AǡLB�j����lоDV�,��Z���V��7�V(�!CɊ�V8�ı*\`�9�Ȋ-[�ha�&������n?R[�)�f{R���T��ڵ`�#F�@C�C��`�9�\~�U���!�՝,�'f��[up{-z�rЗO�t}�F�����l��|R!p�S�s,+ޛ�q7��Oɪ�ƫ��z���E��;�ha�є:�z���:v�����Ypu����Z)�c�0k� ��H�t��,�{TT�̄��򵴳��=�<[Q;IWkb
��3P��>ȫ�r/6����{�M~�On��	Czxj�f��	3GE�t�ɾ��HpF��?7��	�OG�WXb��*�}7�,�p�3.�����9T�:jr ��m�ծŊL�W��U�fs��{�cg�A�9,�!���>>�*>Y��fl�K|g��q^i���9�=Vv����yi�zapxK;�f7�Ցj���&1B���NK�&em�u�^�.��T)#d8�iCR����������f.v-�e����r��������긔~������ ��v�C
k6��뾏��NzUt
��D�>u�	��MwC�ֵ5)��n4_�S�syT���G�zvE)X��B���~��,�����l�e��Y\��h���G��"��BoM��Q6+�MpCh���L�k��=����Q/Prn� �'M���(�!���! �<!_�*#f`�����M�
,��nE��0.��(�wy�{���-�Fj6�7J�:���с��xl���|y��:��0��.]�떁�;�!�U��3nG}OUu�k�� c�@��d�v��������"J��⑵���[�Z�m�Xfդ��o���-����Jȳ���.o	��	Ji.4�ۆ��G7��J*����2z�L�n�O���|%�ѧ��Q����\�_�9�uϭ�^0�'N+�� Y���z��
󲍙ٳ�ZY�*jF�����hcV�ޭ6;�0�1��K�Pb�ss|��ú��#��9�\�̫����>�H��1�|�9��j�s�Sֶ�ؼY9�5�b"�� M�C�F����[���E۬��[��J�Amv>D�sb��;�����6���U�4�J�<�+!�tdxґq0��ܣq�/:Ց�O�]7yԓD�v�W�ހY�ڱ��|�Y� w�M䛕�ܘ�R�,v��n^�ILĈ}!Co�
%�F�[�EC�?�����u3=6m���,�z�uy�W��ì��׭A>���yň!�J��U3�:!��6���d���S���U.%���>&�����li�Qxh>�A�;)�7��^��ƾϝ�Fw=96����I��e7�hu��1�����ϫބ�`u�/U��4�|��h7�M�*~�ј}u�=zU��a�=}��9U�me�M��M�]���̎�l�L��{]��l/�/^���u	c͆a���]ʝc�\��n��p#�n���`V��tQ`��
�׆N��ǣ�կH�pb��H�� �[���#�v���x <�pC�:��OnɁ��R�p΂m��e�B�JOL��m}������^D�Lh���@�i��9��Ve��)��$tmm_*Q%�>�{�������.��*�Ks��z���M	�Q�\��+J�6�ÿ-.�'J-�/�b�������6H���j5ƅXȨ����˻�F���yFg
�`�s�5VL�XY�6��%ğK�����!k�n�}
W4��{��H~��ЩGG\���fF씩�V�2�Q��DN0ć1cGd���J}�~VGmo�L���\v¿/PקmVs��9~�L�R�{'&޷����V�=3[4!��b0}hLl��DdХ���ʁ���d��j���U��D�	���GM������4`�:ߏ?�Ǽ�Va�i����LNS��&�da��]=[�z8�w�G��8Kc�x}H��t����Uq�;�9�qץI�L9�,:����5u�´Qä�,���Q��6�C�>0)���5�vZn4�������T:`[`Ԣ��+�J�2�ww!W�ڝF�[$�AI�Ú���V�9���cf��M��9p]ϋӹ�R���Fk����A�{��i�K�^Y{�t+,K(�ƹ�u��N�5o�Lx������}gMv%E�KY�W�>�٣
��Y���j���b��#(1�\�cx�(ؗ>����7�v2�g��/y\��X�#��VҘ<�+���m,�g.w�m�p�Ũxyw+>�^���=��
��;�+�����|x����^�μfh3�c/	�E��a�#o�Oș����Q�o_�O&o5��13�d�m������$͌��5�W��pFC��TW-��-?��|��|��>�ۼ�����(��!J�)��*�����(�}J%M������\F�\��<N���{ZE�ݎ�2�O��t���w��82��j��C���v�m�(Q�C�����n�!�,�1���9���%#�d2�=������U#�&E��/��X��)�
\on��-���q\5���"ؐ�bg`z������=2������T',�c,�m(�F%SɎ:��{�Y?W�r����4�\l(�\���Fƹv.�7��Bjf#����d��7�4���|Cܼ�_�|o�:����Tz
��q���+�0�?��\WШIY��=�L��,d�������q�ۙ7��� ���*�f�m���ii���vQ㾜����v�8(u�t�:;�w}unė}p�+�k�A�����h�Y�l���nmi{/�Sބ�S�u8F�g7xz�a����ى�&�b����.;	��ҨuK�j�c7����]]�nA�' �m�{��4k����	�� 	�l*<�������ˉ�� ��Z�E���͸(^,�\3	���c�4��o3�� ����=�ۨ�r����N��g�烸l�P����Q�@��=�c]�Z&5����q>��+�G�o���{c�wL��\ڭ:�l��J�e�2gq�f
�dCx<oonB���`0��9N��Q�Jt.�sY�/ 1����o4�e�,c�w]�/�������+��
t�غ�q!�@ͤ�������y2��2��n,��� Ɉ��r�p^K�
�2����Ѱ�#���Վ�2rF�p��|�\\Zq�N�Z�L��U��i&�Щ�$��F�<\�Gz��w,$���mkw�Eh��;9DS����W��n=���Q�Y�����L��+xu��T�]`VM)�lp����l{^u�fOi��&!B{�7n��J>4/�V���Fս`�͘����jSXU�j�E��z��݈�s����LՆR��\ri�B��v��H��VX;�>4r�w;�:%��<��<���P����7M�FJ*ͨX~�"�M஛(p�c�,���kD��ֺ�,�������%d��&Z+���ٲ�����#v�i��t���x��� ������O&FDr���zʅM
)WnF�f%f��;��Щ'F=��ti���Lr��1C�T;���;�-����ˣ·���wzG���]d]ˇis��ˑCR>{ȜKK�ͲO
�ptYe�M��t'�ض�:פ_F�)k؈�+u↺ 11���U:ʷb�C�FEJ�i�6�)���z�:�?r4tL�y;�Q�ޔY�x\}І�ξ�|(+�ތ+^�� Qw.�;�m�Ȳ�m
�d��ӫ�߀ Yet��7ë��rJq���{0�G!U¦tk-��	f0'	�9З�ye�Q���ش[�	׳Tt�JJ-��e7A��ô��%�ָN��P;����m����^d�^��Q��/p��}l&���,TmH���sF��V�Mv�Q�D��tM������{^)���w��M���p�+�3 ��˓A�']Ǧ�+	�:�1��v>�5�} ��u�%3����ߍ@*���a����Z�u�n6��g!�H;���w�j��
�]Љ����a/3�V�.7D=:�.<�ɕ���e��.����A6���p�M�{���=����������vǲ�7[�čs���Z�u�<��cU��QAV(,QS�� Ȣ"�@E`��DEQ`��,� �T���AUH�����TE����UQUX�����**(��E"�b�DU���V�X�@ATDF���e�b��QT��,AA���""�EAR ��DAPb�1X��UA�TQU��Q`�J��(�AQX��#X�H��("��b0UEQUTb�����01U�*��"ȱb�(��������(�2"
�*-J�b�[EDb�E*�(�F**��,U� �(1EQAB(�#�`�
ȰYZ����HTP��*�Q�*(�E �,��0b
""�`�*1DEX ���H$ �>ꙉUIx2:�Z���Չ�\|bp� \T^���|�y[OaXz�n�ۘ_f��
���I�h� ����酫��ꪪJ��	�9�rw󊼇���B����Q#`�F#�E���v׉�:�2�N_�L��'B�̖�L@���qlק �����Y8"�͝3h8�J���^���j6S��;�N��4�dUs�M���v��`h�Ɋ����#�� �b��=�⁍>>�U��5�A^{���S�0�4��"�Ճ�̍وP����QaS1�j}�_����Kĸ����L�y���隌�X	�Ev�E����uc� ǏLB�A=�r&�\<A��<+��Ѳ�9�Ra�~�1�����!�
��Jo�Y���1��0c�j��:�9T���Q|H�CJ��ҭC3Κ��pZ����LeNCs�E�B��}���fqw,������fR�v�������#jk��L.{�Y��i�z��F��x�sǛq�\����J���B2����B�H�%c�����=���)Y����b˿t'Ao��Ժ�C���V�s/�-�����#�HANl��w����U�a-!��ե�������Ϣz��Äkդ���t_r����{��TE��/��&Z��is�b�����ǘ#K{S�w@�%r�Պ�#!�sΎ��v6�qi�O����w�a�s���Ϗ8�NU�$Y�Uz,S�̒���6"�r���6��iA-�_�¹���Y��^}��Xwk�8l%�����)}�e���/xo>�\��2됝�mgݖ���r����J{æ�ap#>���4��2�4����{T�9��0���
�܍:M}�Z����i��	t㌋
G@��<�<!XD����H�����ߐ<+�-��P�����*@��gqy���gε��T�E�F�s�q'k�P�`b_zM� �*�[iq:�������^��쾜�`d�2:���P���~����&z�ITF�*j�)��;��r.Zt��C��XѴ���!�44����`N�����*M�Q!-^�ݖ�L>~��~�ﲕ�-��/��t-��ሟE�a|���Us�
LB^����y�x=n�G��`�|yXM�C��6Y���[��[w*��)��1�(򫵺�dƣ�Oq�474�M�Q*Hi�v)��LV͹����)HY5�8U���x��Y��.�����X��Jt��8���3��hM�!J�Ը�Ӻo��9�V�w�p�,:Y{���S3��mr�gE�%
���5��e�^���/�*VM��f�Ɖ�i	�F�ش�;IO=��yΑa�J�%t��Ԙ+^@�U����鈈TҬk�R_.��?��[�����&f\5�g�	�V�ѭ��)#z�.�xs<��o/W�͵�thx�f�=K��f}^�.��{CG=��g�W�ކڣb�$�����1�&}��p��b�
!�|�F��vv_H��f⏛1��z�4�V���j����(R�cK/&�ƶ	=ƺ�
�GW��A�W��d���O���bnM��fw�-��w��bʋLU�ߙ�c��aXɭ�-��h��&K2nD��{����g^ew��R��k�)0/�k�HB��ȃ�.���s慞���>�g�hc�F��G��r��'iu�ئ�On��O��)���CN<t7�+�}��h#�6�]�6ϻ2(]MⁱL���6��3c��9� �Tcl-.��E���L�&c�k�
�& |�p�|w�@�:$�Mr��������/�J�Y���U�;�p��:)�R\I�(Y��$�cx��ݴ�p����0�ت�a����LwK���)*p��ޙ���:��%��6��VK��ֵ�G�'�pa�ql���DQ���q�XW��Zvs�Z}��~�ѻ���@tԶ�(�j:�ުiM; u$\��뺺^�'K�'þ��u����o��u ��mw����f�������K:�|:���3!d���Y�p��%�w]��F��l�>6��\�uqP�ڦ����
/��[���Z���<�!���� ��������'=�>u��W��@mQ��d�=Ȥp�3-�v.+y��jѦ�us��鞹�5 ?sgA�S�RA~u�����aئ'.���{�6�~�[�r���~G���7g��H��3��`/s�	�Ɠ�Wɚ�k��i\�]�:�֜m�[\�^���
8Ks``L��n���C���6~��ʣe�h~h�Ǖ�zuvo>�ħY�� f;�Ϩ���%�����ӟ���69�ʛBb����"��J��沕z"b�MԿi��o;�N2.�#vj<�I�ߒ���Y�N=i�*����R#�n�:~�+L�����^D������}QE��xiݖ�#6@K��m�&&v�\��j71�U�v���$�}hbOx?�<X�y��n�-?����k�&��UN��j<�ꈩc���E6T\�gcEXf����>��M�Vn�����z���șz�d�W1��P��ȷ`7a����y`\Ɨ���W��ƀ,m���kP��Iѽ��j�J��i������b1S;����	��Fۋ{C��9�O1V�n�v�ꐍ��}��2����!���2/v5�;�N�
R��w+/)���5Lt�RH:-+x6�/��'w�mqYl��)c� ���֑@���n,�����na��k���ޙ��D���z/d���mx�嶪GZd[���`�V�:�Lu���g����gzj��N0��gm�j �z��v][��>d%6:~�q{��u��im9�*����ʵ;/O����ODm�� ����=���{�8�h��v�oK=x���C!B2�P(Cr�m�T/b ��tE�<İu�2��#�Y�v��V�>�v���B7�q��J�9��F4h�J��K�A��-|�qA������˴�]��1�Ḩ�Y�W��7.!�X���1f��W���P�Ӑ��'uy�3FQÒK�ݙ�l���h�6���h(91R��q�=T�{<��<�Y.ux�Z��cB�:ʸ���v�#�>	�Ժ�w��9���^�`�H�������\�+�uMﬂ��a~����f��d����BO��`I�5���W:2�S��s�zh���z�f��߳;D�ŏQ�<�:S*�c�z�ρڗK���6_�]>�߼�������_�����\;�j��[��>@�K�y"	��$~�z�Z93`�]�b]�A�)֝�Q�z���\����R�SB�;���׺��B�\qD�oi~걓�{E����0����G���8'Z'��L��)�㲻���Tz�J���Bko��+}�9���t���v�8�zU�e�����X���t�;1�[gѷ�o�>�;+�N�[@��Csi�+^Cnhddh�C�h�gb��#��TWO\�Ζ����!X���	v�oz�w��3Єd����Q@�H2���������f.vnK��ĝ�[N3�Y׼�>�+)؋�?a~c4!Õ�lmV����\�Yܹ�o���C�~��P�P{{�ٚ���g�D���f�E���s_[|`����a_.�vwP�N}]㧲6��n���b6;du���$6辁�"szl�>vL�4�\��1�� �<���v��jylmD�D��/�R�&8���Vz]8�"��t
�A6+�%U�*�\E-�_��>��}'1N7/���]#!�iCX>����=aPw5�UΩğmx*�����g�]�}2���.ꕂl��8��*pS�rc RD�>U�}�|N��1B�(��`�8�٭�3_1��4��Ϊ����뜋Ѵ����mN-�F'g�=�)|��?D�^�kp��5���GW�j�b�L=�5�fư�v�!t����$�˂�v�P��;��a�[��S0��3��y=�9h"=<�&y^>w�gw!�Z�[�d,��L��7��Gu�G��QT}�!v�N��1����zU�ˋ��Բ�%6�x�ӹ[�5�(R����� R�\�f���~жs���E��0���K#0e=��`�`�|�/H��� ��s���);C�&��y|���([w*�TE7E�܍g\��o�Q��uβ#s�c�k�M�s��'�2.���ٞW��WF`>3��;,����J�����E)o(����38 dA�5=��'�M�)n�!K�����1w��+�wV����%��F�φk�ظ�&`�h���|����=���ǲ�W@�Xȍ�.�
]z�K����t����DQ���5S9��]�f�R���^����wՑS�jlٶ��xd�z�-��Ӿ���n��\]�yF{َ����J�#C[mAU�u��@���E�*�m�0�tT-ɭ��b�r�NG*�-��7�&�F/z�7�DE�̖�%&���A�8��ҿM�phY�I邹�.���5{WY�k��q"C��͗	S+���[\�D���>�{�����Q/ޕ<��f7{�˶�\�0�*�d,��\
F������K���֌��SM������4���b;#ws�F���:�������^7*k����L�α2��Q*>�L�P��3^�89��>pF��R�����N���/��W���Δ�U�dӃ߶}�k��w�����)Nlۑ�j7B��A	ҋs�/zl^��������9	"�5�^�{w��A�R���@ YG`TR�\��gak�3�'@�;��]Ld������|�1���������P:���缡�^,�����:����͋�馡��ck��-N��%^׆z|M����<	��T��G��}����=&K��/�8��k;��M��aF�����Of�YH�AlZ6�\�P`�Ss~�dR0w������(؉S�҂j���M@9���)q#~���)��ƍ��@�́�2F�lM�e�kqAl���R���x�Uw!XH��3|	�=�Ɨ��S�W�����U���˻�6��>[y�ۯI�`�[�&���,D�'Q���)�ʆ�^����]wS|��)0�z��7U�,����[�<�3Y<l�/���i�,EƫQy©�O���W�&1[R�F�Z	���£b�c��ǫ֡��ܬ���=OSr�];I��k�W}²ۀ��p�.��b&
2��3�Ce���|�=�4�2b���J��K�{�d�6ѽ��:E{���x4w,5���b���]k�#��mچ���}J� ��N�F�|Y6z�>Yή�#��\�o���Z�39�j�2��}.a��>e�zi��>+����֏f�g�*�rÕ�s����ƽ㱼9�RL�HٚJ+�@�d8Sfp�a_�k�0�NS����)���&2P�n�!N��E$T\�gch�+@�#H�b��z�����ʬ�p�7H����ѽ:�sY�C�c�R�Y���pD�=�����=G׽}n��:w%�bxJ+��pC���T��	q�x�6'�M8^�я�Ӳ����z
�>�fv<����x(���kY8z�v�d�o3�����gm(�WA�Ga.{�d%7��{�X���W7}�)&��uEC��O`jiF���Z�t�NPO��)a�>�ʱ#c\�b/aoj��V�D�'6���&'a\���
Ct�q�Tn Ρ �zM��נ�:�v׺��	3M�8�a(Y�T���6n�v��b1ɏ
T�Cb��FJ��L\���f��/v�oo� s��*no& R��N-�UOCr�ĲpE�gLŚ=S̞=�t����ȡ8s����QTf$E���zr7ܨN���~�F���^�Ae��<};�����B�T��e�ȑ�\c�݅�֮��U!^Iv.����;��W0�I܆oF�k*51����ԣ�[r�c�ņR}B��thq�ے��t�WNwv͇��Z�Ȋ7�ǈѴd�K}[��b<B��d�\�͖+��v7����}E��g�غ^j�~�,����?Rl�+�B�sAв��XA[:�	�b��_Y)�h�$�<IF�����U����eA��[���1�K� �S��x�U�{J��Hl�$UK�p�U��If��.2+�h���nu�����v"�T�N]�붫*(Ct������8��*�3<�p(g��sy�CM\]�ev1���������X%]w*�I�#p�7Dll`�C�h��أ������@+���K��w�M&��7+�:VF�)1�x�3��|�؇�>>�'×�;]��zo�0C�|����x��zTT�c���~E۬2�����#i��hmV��;|�R��
B�Y4�a�Y�D�@�~�j&������T����~Um���Մi|��K���"c�m��=�V�ѓ��!�l����ƥ�zw�|���`�TM���+�y -�r�x���B���u��ʵ$�z���m��R�@3��\k �N)ў�W��Xn(S��z6���Sgh�����ژ��T�Qsoiq�Y���o=�[��&F�v�d e'�X���g����Wh����kV^�^�%g����!��ɇ)�(� ߅6r^������m���s��gG�^�w��"UY�[�;�O��l�j#���.������8��Z�]he	����Ӗ������8�����*Gy_L�n��ɮ;�O:�n��!�b�[�(������X���Z��/$�'��5�*j�lwi�LK��X���	���Y��B�p�C^�����NY-R�V�� ]��,�޻o(0'R�7R��wS�W-C�\��\��QA�7�.�=39���7�ذ)*mlQEw׵����~z�s��8r��h&L�c�0F�'<Xy�ֹj!�a���.���B����t���/=#:u�X�IS��k�����������ʅA61�k�*�O�C%gsDU�G���A�ֵ���E�/L�E�b�OA�����{�[QgtU4�؃���´(G�V�z��f�4����q��}�����J���Ҋ��\��W��L{���nW����J�6`�A���dU�z�f�yY#�n�����Z���$ZU�(w�w(b�}*�-�Wk�`(e1d>��G:fh�����{�9ø��!�{=��[��֮��-��n]v�f�W�8���qy})���s.�hw�˅nj�/���]�B�:�=�\��K0t�|(V!]EIB��ά�wOu��Gy6���Ulʞ]�|9��0Wg�u�1���2`����]�V,�Νĕ��+8 ���{<˧��kOu�j�[z��Jf�.���}��7}�YEd�R��I��C��J��aΊ���j�dJIFV^	�u�ݬz���\�X�XOp3�1�)
S��1]�r�U�����"&G�J�������y�O�3أ�hoD��k��l��Ou��u443�*n�������{ Q+�)!C�P�W]�J�Y��UXS��U�}~�8�.�aJ���B=z���ZIJдR��b�{q_ ���0��{9MT�:�%LyZ_�\�*8���̢]�/1!�K�G�>2��g-���sȺL�a�v�����ա�=��2�1�z��֐��&��gF0#z�3��[՘8�|[v3Oc��'��9����ۛ��q��_b6�eC��'1fZ�����7�}��}9���;��z'F�ٰ7˻e�E��N������f#�a*VHt�JE�v�ӧ�'_X��^��`���^��tރ*�'MA9凯���b���~mR����Py�\ *�j
;Սd
��к���GpJ&�㦀�n�8�JI���iA*Ə�`Ll�&Z�_m��ׯt~��;p��c�ɵjQ�QQUV(�QQTb2�E��*(����X�"��
�#V��D��(���EA�YEQim�T���i+ETPX�b�DQU[l
�R"����@UDU�QEDQDTb"�b*"Ŋ��b���
*�1R((""��A,Kj�X(� ��1E�0EH�(���1DDUb0F$VE�����"#b�1TUEP��F)�1��PTAV"� ���"��*�(����UUU��"�T�`�-�H�UX(�Vb�U@UPV`�U��H��ݿ��s7Yލ��>���p���/���v�u�P��L���|�����q���:yu۵��8z�W7��ܩ�;�޻k�z�t�/�8����*�.4��t
�/PM�������A�D�T���^j�+Ҷv�y��Û�
,��O G�Z�L��A��H�*��I^
��d(��`�w�:��W$��N�
zE9�(\����ʵϸ>'߂�(QQ-=�N�-;���y�|���~�aL�I��(��\�h�p;gvC�hi�Ż�L֋�;�����}��j�'=�V*���C��>K�2�'
��xˋ�<UX�O��0�	�o��;P^<�*�Q�;�Zj4�᳂-�v ͂�DD!����UDdW���ɥ&�C0^�s��K##�rM�׼�dD��<�"��>SLb��'S�w�����J�<�謊�l��.b6�^��=��ZQ}�n^��e�
�p衬�c��K�w�g��hh����C2@~�#>m��ޓ}�{5{�ȺoyC��dx�f�=�q~L�^�.o���DG&�WE�wCkg.f�]����π����E�`��\�8@�1� ���W�j.�ga���`���n�5�^N��i�8�
�$�=�u;��)<A���N�X+מHN�͘\^����ȷ�?���bb��B��cX���C��ԧg}�A�����Xw�f	����? d�(��:�G��SIx����f�\�.m\�J�^\��j�gS	���LQ�!�;j����j��R���v��uUQ�Ǖ��:�U5�r	U��������k��y��Ki����{О�`t�A7����E=���;{��L[E��g��y�JL{]2�(�Vܺ�1�H�D��asѕ�s)�|1�
u�ֈ��m�	S+�����.+~���9����tڰt$W��Qɸ4�Х�|����0����86mH j�kK�'J-�Kg������C�$�&:��S�1��ȥ�qDl]��a�>��D��������ic9����k8fӠb�:lD3>/"��e��]����� �u�!;���8ǟ�x��l���#vJT�-��|�0���*&��R�E�2�#pE�����p��Z,��J<D=��}]j�=j	�k���
aΜ/�zo�{�N�Og�0h	�3��\�~� 6���`����p�h�8�:j-verQ���f]��3-�n&�n��� T?:ՄXhګ.;�>���x�{���W��ȱP �����;�J6�48,�
@��"��K��[`��ZF�YN�mc�c����K���{~q(	η}��d�t��5�myv�<4Nˊ�L�Q�/�v �����yk�J$�rz&��.a[�$��)>sd����)X��
��\6#��q���,B�3& ��PMt��p;i�
*�`��Ǽ�'�)fsd�gW���
#	noD� D��w"`��1�c��`���z�ܾE�]lo�ݔד�A��1vGg%�P�B�S�hp7jyxV�x��i����\/��7�q�¹��$���Qg��ړ�hl[�	���£c)�7�:�z�L �'))2)�mF*\�3x\�}�y�3d:L���)�3�����J�ñ���TQl�^B7/�.�]5�VZ]m����:f��K�(Z9�EB�Ę�/�g�|F�Q_��<��r���"���{��ȇV�K%�s=V�"��P{;�(�}J&21r1s��;m�{���N��:�U�Bm�ȷP��B�cY�7a�<��SޕC�!��X�g�׌��]��(��m�Vρb펯���KM�4؜:i��m���峅C�{h�`�6�I�e{��vfYz^>ah=���c|@��0}���{uJ�̄��Y�[�{�?eD�|��;�8ܧ�	6����<K�]�&�֖~=E9��^�{���m-NA��,���ʼK2N�w<�\����ge6;�*�}�Ew���!�ۛn��U3��&���M1rv*�v�E39Ϲ�4�'
�����eǏÛ�P|�}rZ������,��i9A>6��=����
c	����,-����Bk`��Ae( ��s'�F!1�7Ϋ�2o�l����ͫ��tm�����ʧ~�n;}9r6
�����4:1ɏJ�3͂�`t���/�`Tl���kv.Zu�D*Jo& S��N-�UOCr�哂/�:f,AǊ���q8�m>Sa��;��N��8+'��1�Z-{��o��×���m��~y/�cgwf�X6�wӊ����غ^���<Y�����腒G���24X��}��/��}:f6o�}�A���Hh�����x	�Eګ��;*�7J��t�ؘM��X*la�	>]b��"9��Bo��-�#S�����W����Q��U�u��#��T�qUmmyz�5�8�B�70�d�Ađl�m\]������,lZ����!���{=g���o�*�p�r���P�fʈ|U�6�FF��4m��!�r:��܀��sIܷ��+&�!�w��C�e̢�;>bvY�'0�Z��e�&�w�T�>�����yD����/^����0f�.�'���)�]�0��(�6�^@�t��[�a�>�i}����X�m���������Ψ����2�;��͏��B�VGO�1�ЄdUH��Q҆�X�lbvzF�]�4�ok��z�[��CL��G0k#T�YM�,�Ծ��A�p嗌M����2H5�
~�M�"�=V:c��	�u�ם�L<���+��=�r�A>Q��N�t9sIuf������-ֽ�/�v
n�<�B�4:d��E!��@��dמ�;���G<��:�R��!��E�^NN���T�c��Z��N8ȿ)�z� 6J�Dd�b��ʼ�B:�N����m��m�Qd�Cx�j���
���>��ҬuN$�x,��egFU�b��V�Nݥʻ l�cIcf�!�@=%ι˝�U����uϽ��Y���OXUR�g�+��z�����>�Ku-��缅`�� Ř��F2)�ޭ#(���"��P7R���6���0��K�g���>���,Ϫ�<k�g:�O�����r�T�ߔs�q=^��u.��ʕ��o�0��O0I<yZnZ�4o��/����&�F#����z�����n��"ZHL��׊h�f�rjX����"�6-\��$"�kF�}qʪ�si��Y���^g�+r�l�V�V��F�Y�#��ְ[�|f�N
S�)O\X�9u�|)�=���w��E3�wQ�q��wu�_���=&�o��%1�(�����ɰ9�F���O�i^*���z��y�u���ٻ�%�"�Cɨnor�1��k��)�29��k�S�
rtߡūs6�߳{m�-!J"�*OyB�n�p��9
K���I�}'��bx�1�7�:r7o5�T6c�#5#Ǳփ=Fa�t��B�e+�5[p���%�A�ɓ�,!Y�~���S��Q�U��7���"۰���������:�[�{���Z�a���KYc�V�"�KS ���:3�:�C�ܪ����i�]>q|�U�9��q�@�����l���9��RR`=����qA6מ�l<��o�L�^�ԗy�����oj��1�U�*��bFVW)��p}�W�@Y�!�.�8.�/mRY�.G?VVD^װ��-��R;ڨ�ߖ�R��	l���u���:�d��)�*��r�@̟����q�Z􌩳���4�s�������6��b��R�}vq̨����޹����R!�]sN���ބÐ{}ʡ����8���K��F��F�ǏV3#���!��ݨ�X�����Z�whI�A��r��|v�l���T�^�+�wAU�^J�LL��wfA�o:��y�q�:'ӓ���b�Tx�|k�2{��jmU�w�Q��
���֊lJ�9Mk<Q�ʼ�7�f^���ޙz��>������N.�T��G�b�XW��o/�ا�$�$#4k��UtR�0�6r��#DT�hE�������B�gUY����GP��7�'*)�D��*p�yEi�̫��$U7!�sF ���R�B�
��_NǠ;α��1��w���gv3k�w�H=V��r�����U�X�s0�b��k�x��E>�'��q��|\�.�^߆o�ք���ǔ�W%��l������ɘ����Vq�]z�"�Wo.P���w���V<��Q����}~��8����d����ʤ3��,Z�ɟ6���o���^���=�%�� f0�c�u�A�RB3ɚ����C.(t���;|��hKL琍g�1{�?�O��7N�1��z .�b�)�fB=Z�)�fk`��<�!�z�R��K]�r	�RL������g�g�خ-}�`�-�)�1�NF�����E幭?c�(IGwb˩h��S���/�t�,���mgc��]�>w���I����� �N�!ʺ-�R�9�,��.�QS�y��L�h(� ����){`�Gݽ���-U{�ÁI۹����8�[�Sb�_u�O����{3ѿ9�P=HG_��C��b�IBǻ�4�_�އ`�Omٱ��s_n�ν\��L�8,K�EΖo� ����l;������S�$�\�-A��{d�n��C��D��"���+�:��9wIPb9�#MX�7i �4�����碃a2�W`�E����������b��7c��D��G���M�w�=�^T��U����)f��0�n�&�X�P���M�ݡ�#��t�U�1�ʅ�js��gb��r�]��qev���&�n�wJ�z[��gh�f���Sa���W9�;��:�4�^�r�D�z�d�1�[9<�H�syB�¬�#��gn�m��MB��K�0w
'\��ϴm,����XP����ȥCGU�F4�]��p0Jȉ��&�[rv�f2ΉC�*��2N�=���t��W&��#��]S.�MtX��773��œ`Y�:R�j\�5Anٗ{��f�Ռ�,�h����E�	+h0ǝz��<b�j�_ey 2��Ȣ�=���6���o/��w5YC�N�/W�E��D�WEu�EP�1 ��C9�Љ���bk-�^P�XE����}CN*�jf�W�\�̤e�)��ƞb����)��6xi�=yuc�5��n��d�m���4�m��+`�,gک��פ�;�hFן���R�kg��\�-#7,�.X�ƅ����S������l.i������9���e�}Z2�wY�VS7:Z��f���4}�E>'x�"vW�/V�Pf�^�E;�6\p߫�\�x���T3k����t9��sx�uY;�9���'�x�d>���;�P�N��O[��(.��t^���*#7�C�z�+���I�kj�w�}��OE6C�S�0J�u�d�[6��Q�ގJ��#Wq��{֬C{N���@68#}��Qze�v��I$1˱@��OUU��u�#�Z�*���ɧd���=C�3�x�\q�vD�95Z8�!zZn�
�u�Ks܎��x�J�U���}Np�*�қ��q�_�R���*���sּ/��çF!\&2K�c���1ysod}c��WF���E:1�[�:�=e��y��Y싪�z���Y�e67]S��)P��z�u��U��Dqz��X�[��c��oy���x����5{���Dzv.�b$C�pc{�O��z��3l)F��__N,k��m�[{ �N�V��>8��6F����ޫ��}�+G7o��X�X��>��sv+E'�b'
�CryYX�NH�{��r�R�YMqz#��!=�,R�c��=(k:]��w�Gi#������׏Y-�ۤ8<�bhrc�!���H�����L�9��b�/�<�`�˾�)��+u���}�})�=L{w�
�E��
�ToR(�KHF�Lt��m�v��t�he Ҷ����]���l��SRnߟ_Uj�b�������U���8�Ti�C�Nu�]c-(��T���Yۺ���ފ*/�u���F�Xxm�4^��xT�ś�~�*Ewg�Y���i�5$t�`-vni�k�4snE�Kq����[��D[n�4Ov��-��x5Ĕ�>��,���z��1Okի3L%��
��`5�]��s����Y��{yqy�͑ӷ�^�ag�Ȇ��(�V��srXڴ�9g�C+S��E[ܬ%�D^���+��Ay��/n����r��be�W��(�b��Y�A�����\�I8v�����{ET�k��5s����]e��|�p���;���C;c�Е��/�*��Mq�K1�;,��{�f�9_m���a[��"�߅-G=!|M�
��Ϲ��V� v��ݬ���;�|K�����r�}�tFf<XюX���霶-�vr��s�S�Fr}�oH��Le�S�H�\tc�vE_��3Y�u������Qg+�r����0����$dổfg0�ck���lσ޻A�Ӝ3r���)lo��mUr	J�t��)�<W��ee�gJ�h\��j�F��v����ݛ(u`����o������v]�0���F��/��� ��x��8 "��>��冶D\T���X��v�0�_���/`��k�|�.ۣq�v�_u��	�>ѡ�ٿF9��ρ�M�1�R\خxna=��v6�ζ��;l.����Y�ӥ#cN[F
E]�;��q;�k��Vf�#:#�g�`)�ʸ�}�G��sY��C)��{Ưd3_�Esy}9��F/(������0 ��Q�h�C$���bp];��.�ev��w��,nOY|�j%�t:_�ņ(�A>�
mmՋ}�<O��{��ǒy������ 3�N,�{�^�ܾ8��c�h4?Jǽ�{���k��cjL
���#�\7�J���1-`�A�����W����j��*�l�P��aM����w�K�;�n��hjQ���2V�-n���5����(>�#��`*��N�_^�����-��of�0g|���6?w"�,7<�+/>uKa� w�7V2��Xf�1w���*�}����Y��[�n���T��:�]e�c���v�Ӟ�Wqkw<���]�{�t��O��7V�p���O�׻9�.\zކ��'��"C�HͬoU8�׮�R��k�:��N����|�V�l�G�ׯC�[ٰ�!nK�Ӭ�Ѽ���j4�4aim��|3������-���-�Wm!9�A����N2� �Km�Nn�զ�-\aC}_�צ�r���A���T&	$;��#tEP�$�)���z��ʥ�H��y|���M�"���[��(�����@ȵ*�Z�WNn�h6ǥ�S,��Px�����=�aC�;��ۼ�=}R��2� ����5
xco��⹗�`��rj���܀њ��"�	��!u*VD���ݻZ��U��I�RHN�����C��gOl�&[w�D�`���Y�s���3
��'ѳ}&�>�3 `,V"��x�eD�mTP�*X��PPc"�QY#R��
�����Q+*""�$b"�"�F,�n�R��J�Pb��Z�Uc%J�DQQ���E�(+UH���V�UDUQ���)m� �#UUX�1AE��QT\!bQPQp�QPQUDV
�TQQTQ�� ��R� �Ȉ�(�U[j��DUU�6�-�X,�#Z�ATQp��A��X�Q���+X�J�*N/뿱�������p���x�Y��ب�l�(���^�X+�}�v̹w6\ﴊ|��`ȱ�ja�R���㳽�MEn.���Vk*�A[�~i*W���P�.���o�v�ޜHF�=|�{[����av*l�V%�v>��J;����Ƒ��'����3�5�$��S�eX+�w�qQ����հ�S�f]U�}�W-�0��G�E�c+d�܊�y����[X���;�x)���ع����4�ڍs��ʭ�ᐍ\v�,�V�z�)4r�#+��A��k�v&��,UC[qX��{V��d�a�T�M�Ш��]�Q�
�	@��ʺ�5V�:����A�
��^�rw�1����V����h�����v�zy�nj���D
NJ
�2Dp*{M��{x2��֏W%"��p:X!���s�x���V�φ[}�N�[F)��D���U�[rv�\����=��\!�N+�RX�n����� =�j9��7�����/l:)�C�'�h��@W/���e��� ǝ#˾���D��t��J��e�+PY�0��) j3�⬲����u5OY���Y�����9l���ᇯ?g:WIo`������95�3i�ˤ��r����&��hk1;��U�ڼ���%�؛�;���[���F�5ғ���g�OF�:ݷ;�v���Pj��������x�봪d<(3��s��r�빠5���R�𝬪#�[F��.T1����vֵK�C�C5���l���g��Uof�Qz@���t`��/�&���#����7;E��tk�I�&�'��7���4����7���5�=V3��ȹ��O]6�~���(�LDNC��E��[n�%{\�tW���P�V��|'�Q}^(.9]���B#n0έ��wrq�곩^ܕȧ�����nG�lB!�@}�|�}��4�.�Q\��WҘk#S�!�]�٧`)��华�*�U��k�(�t�I_����u���s;��;�9dr�k|���c�_|�,�7�ֈv�z�|���z;���l��gI7 v�Dk4>�I����L�^����j��j�X���I���7���n��}�P�DV��8��R7��i�{�9Vi{��-��Jz��+:�W^�'��`>��-Y<���\��#q���;����I!nJ!wo�n��V�Uo���c4%(	!���͌�I��~�d�D={�)�]��By�~�V#-����*4��U��\�k(1M@�,rB������47�eh�-��aF��3�����sh�%�c�����h4�P�5�Yk*򭹠t�>�\ V����W_Vu�Xz��@����eKy�M���eɾk��G	ʋ�[Ou�9���뮝O�uÂ=.u1���K�`>5�[���َ�9���
�\�eko0������BX�K����L��b=��#����1�:���2�Y�YU��Cƅ��l����ꭢ۵�0L�tfn�;��b�b���6=YH��kš�t3PDRk%���a��jb��k}8^6�����]b���p��zQ���AlaJ�ǜX'����\���g׌њ�����u�X^O0�Kot��k8�{v^r-򃭮��kU�M�cs�;��m��'B3/s��K��5��ւ��u�FR<�]�5t�y�g%\&KA�� �(�s��������Q��K;��M�G�<X!wWX�S���P�V��g���/�i�5��f�2�8�0-o
v5C�Ձ-k������jT8"vzK"����)
)�\��~}�Xz�/���W9����v�����sڋs1��C;�.U�wLa��y�K']ݫ#��tB�i.������y&���z��i�j׷��p�*�j�{��gt�8�,i=��p�캸z��k�cT�,�Y�k�S~t-{Q��\�����%��C^�|�SQ�V�*\�Ա�	�Z{ �N�V׷� ��8�Tst #��1�fSjDΰæ�ry�D'`�x(�NJ�Me�23r���;ԯó���T��]e��!3��*X��`�i�C|;;fs8Z��s�Hȼ�D'V�O�]��� x9�cɋ�c`�0Ben}�K���nݥ���dɻ�Kyl�� �˶s��u���T���k���?4�A��OE�]�G"_�䧕����p��1��v9�zX毮�}��Nu8��R�|����q�p`|���fjd[�F%��{'gM\u�����ʱ���Q/�tr����w�j�2��M����cr'�p�BleS}sA�A��s�[��-9Ե{�>[��`%u㠹X��73���Sٌj��"�����2�����[�t�rs��Z�H�헗��FD���~�Ż��}]~[�^*/��3�a�:����^��ْ�v���}r�_9�f�Z
H�=�%J�{��>ʋ����g'���89#�F�W��7=@����.�OCm�k}��9(J����N�_��D��Bŋ5��"�j���@�(&�GHZ珓V�eJ�N���}�ū��⧺�Xի�.�E����b��]�d�V��ى�*J��<��iMjY��wD6�;
\P��Z�}*�;Q����0tо9����vJ�U�T9�O�+B�hۊ�?:���]h�%51]���)dT�����ğ���`���D��8*Ό�w�m�i��1ۗ#��,�z��;��tD+{7�Yٝ�i�R�v N�	l���ҹR�$"<��n}���5\�n�}������3DF��cK������dV�}�H���A}]���.#[#I��)���5��g]yU��&t-=�)@�'׶�a�Kd�(m�[��Yz֋k�BKF�p:}��~sV��Q�'�*/:gC�39p��9�Yg���I�5�`t�	l��%�6%��V��ܩ����N�'�Ʊ�ɼ��5�t�#)���p}�f-I��|wp����$��r&��^hk"'wz�.�筗Y(lt坙޹��X7����aH�I�ڮfp>T�lӭ�x+v��YU�J���ٸd�'ooS/R0��XϵS�l�V�:���S�xNf}C��î�I,�m�t�Lf������`�}UogR��R-�w]<ݦ�D$äp߫)s�
C��{5�)-��u5�¤����41d�pW��1�|��=V2{��(> b	�5�[m2h+Y��9و�G�����'(��kak���7�g�'C�oҽ��'��kPz�+nVQ���q�=4K�;K��z5;%�g��7ޱ_]�.H�]�>,��ik�w[��.��y;fq�Q]~28��un��Z����d��o����D�v�]]~mAp�U�h�z�}�(.9]��{�uR�{U�!f�#y�R�E�>�V�W��^T4qO�b���7u�v���˹|��pk�6w�K�_v?�Vi�f��=�^T��ʮ\��_f*oxM���MX`4Ѳ�_��vwhr����F���c�W��)o����������2+�������t�ת���v�:��A�*��q'l�ܬ摳P9W�X�gq�������j��l
w�eW�2���u�Z������5�C��fw�殾;{sLx-�>�Q�;�b8�w?u ���X����g�5���zۚJ��]4H�ݕl�h�ir�mL�B8?p]�%_s&�Њ����ɽW�z��Ck�;y�����D����r�ɍ#����*�����x���8rqP]�CF���y�Vt���Ňg-r��}�];�K��������x�+Ԏ�hq.L�3�ݝٻT�s��eQ��	�(�;�c/)�4u�����U�7w�-�a+(��H�v�*P�}@#cH$���W�2C�s�]�U����������R�F�rm��<��9�c4)�}�+7�*�Pɡջfrp���8Ь��6җy�+r�j���Ѷ�(����4��N:�~��@��м�f���r�|ֳ�s��J3��=�N����R�z[�8g�m��oW�Luu�z�&C�;��汔W�k�����Ey�\|�v+�|q��/.�ơ���pO�ʹ����E�=m_��w����l.*�یV�츘5�K;R\�?J�Eu�����!s�!�Z�>򞈕cT���S30��������1l`EW2�P<�V��k����+]��2�l�L`,TEV��^��&�=?:��E�2�v��o�����>N���3˺�{/��z�]�?6v�x�%���{V�v.qPz�`�ƌuv`���M;�tve����Vr�CWs �t��r�mL�E����A�v�>�<���Ţ��6�\v��D����<�_>��F�����琎r�כLAr�]�&�@�6�"
Řm�w��{0�������$b�q�)ԙ��go���Wb��Ĕ��e�*o�΃i�N�]潸�8��z�1��)��2�yE�~*�H��zy�a;��G�R����u=5ޛb9)[�kF?'�G�Q�Q�-�!2;�D,a�1�1�����:���Z�gx����Ֆ�+�}4
.�Sdm�ps��&�1�TV7'r�:��x��Q�X��&9���x*���联�-���P��.0D�;U���Rd�pڣ�W4����v��m���0�h5����������#���k���]�Q�h6-�V��Y��B�5t-H�oxd����0�:�k�W^�Ż��}]kz+���lU�u�/kcun<�'^v�-�����1�^�eRK�,{�撥~{�^vDa��N1v�0v�Ɣ`I�k�����.�OCm�k}���t�_��둷[�&]���9�g�N������S+��=�#�
o��馰����(����:-"����d/�<;ϜC6���ʕX���Smy��7u�7�+f�F��C�j�H+��[}�.�l9�A�a����hnmN{�ܣ7Ht82v=b��ݍ+��t�k��f�J�_O�}�/��������z1NF����=�vu��+L�Ҫ�/a�92����{4��Ny6i�R���hhZp�*�;V�<V����ܗ��a(]X�&��גƬ>;KP��P��kڶ�Fe�zf��i���frl��8��!6@���n�V�
���tOdI@��ŵ�lZ]�r�֒=�\�Y�W����L���O6�I�oE^�l�1uV�pȣ݅�k� 1,*���P�:���ʱ��g��#���t�D���rc���!���|���N¯+�ܝ�X2�>�(n�t��@T�]Nq��:k]�eP׉�Ha�0M>M{��yW���-�Fg{LOT������̆8�௥��cj��s^|"��F�:ݷ��G��;�����Xi]��T�U9���Tq�i�B~�j��J@�S@��4�tyy��W}Q�F<�>n�=���!��l"�k2a��v0,d����<E�����Qa��ݑUK�@��`���Պ+;�%;-���w��og!Zl�xu��;j��;%�\�Θ���q����EpS���GS�� }\�n��iI&��]��7���	�ș�	��y���y�[��֐˵����OzS��{�ֳ6:=s�Y�T�<�#�`q�Q�>��ڦ�}�������V�|m!nXfA�7T����)�,<���Q=vlVԝf��%�w�������]RzLj���q
�f��vn-�l۴�w`n��[�Ǫ�.K�x�U����8���M�*3�������p����ngjE�gp�����b��K��A�L�W՜�����&g�=E���d^�$�1����u��w��l�u���薋N����e����v�F(��.�t8\���w��Z[�L�w��E��`η��C"m�m��8���.͖�Z�2����dY�lw��,��o���~�����e�~��M�mi?<�NM�^}Yگ<ZZ�5��"�=UO�3,��(�L�-*�U���,�7�&���`��˪e5
$xzj�,}��>��y����.�˅fĲ¶=4��;�-"�1����SxU%���J���L<�5~p�h͹�r�3�0&Q�OgVX}:� a�2ܦ�e�i�lXĞ{(w��띈��o��<�|���r�UhG���(t��7��T���*�hT�6)�=�2Շ6�˂nc�p��3�����p�D�V��j���N�4�����)�0.�:=j�K:mUa��NU/��Y(t_,�º�Na�E�\��7uf-yw��r{m�,���y{�����Z��x�[��x�Wf���R�s��OHٴ��	��C����.�=5Zᝰ,���|�Z�V\y�t��}�û6rH��C�v�p�ViAf�r���=�~����o�D�Y�S�8}7f�@w�Y�'�a�ێӪa���
��9ZrKH�3M��B�:�u�'1(���e��F�C�m�[pnU�������K�8�q�J1Uo�G��`g��q��>0_jǴ��7����^^�.D��6�PՎ0b����e���^���o,�,�{L�}:o�(x�u��U52\��mr�un� �λM�&�%�Z���״��$���&�D;TڏrV+���vk���	g��L�ZC���w�R�tU�>��`�CJ-�;S��M�q���-�}���=�u�o	��CM�|��#B1ɭr�9M��Hf�0^sږc��{{�Y�Ӯ�`i��[bύ�z���W^B�]#��d��n���Rwx��o���\��QF1X�R�"��r����ej�"�UQUTJب֌���Z�TejKL8UTX��R���+iF��TbV��U���Y+(�(ĴR��D��������b�+im�[QV	F�DVW	����Ū��F�%A-Jb�TqT�1QT����ZVQ�2��K�+R��(��hUTm����UKj�D�ZũjPUX�QV5����TTKE����+R�X����UH�(lQb�B�R6�Em���V�VEH�+%`T��c���
DkA"���*ZZ�aX�U�TURLc���"ZB��J�� �B�T�X��V��g�e�5Ͽ}��־�qMЍR�>5^f��:Ⅰ�.���c����>4�<������q>N�r�1ٻ۠�˖x�I2D�s�5��}��m1��ı����g*�����p2������u�󬫞:���~�����>����+d%���ڮ�$��Y'ʽ�����-s���^���8l
�d\��A׳XGԒ"=�S���X+�xtH�Ҕ�(�׍dr[v/H�\p\�"��A��dk.��S�ڎ9����sS����^}����W�p��C�Z'��@��P]s"�me�$�]��<V�j�S	|��Mk�!�ҿ)�
��GV��"�l+���:C4�y�Խ��{��IU�}C޲{N��V/*lpu#��-F���b�oI!����l�U����{�G��F��pG^Ȩt�C��T��s�|�*�s��D��F�]6��`����v�srA�ְ�tƔ�*5�=�«^�} ��D�{V-��˭���wZ��՗��,	쫙��z�<��������&	��e������p���9�=*5����mI�{!w�-��g���6��8-�aºѭ���W���L���s@�3إ=՟���yY0Wj�Y~s}AxA<�gOd�;6N�k/|��F���Q|uF,J��N��P��`���qM��dh�����]f��sתD+W,:a���#�	��
�5��+anv�Ü�n���Ofk`�S�#D�
{�G�X�1�h4*�hk:^�к���Q�ӽisKs[j�=N�M��@�o�rb��i�h-�=2r�N�.z�s��
[��W�.��L�V[ַU9��T�z����7Ċ��k֭Y�i�	��;��P�"�8ЬA�+u4F\�wm���x8qW��57v���-�b��Ы���U�C1|���\�k�׊qs!?S��w��������d:Ҵ�<�C}!@�z^��x����ԡ�{͞�=�Gb�	wW_��;���|�]5W&�Xit���q��{�FW��T����Z���h���]�dG9��(��Y�6�0��8�a��B�坨)q�b�܅��2���W�u ���Y���*��.��u�*������X���m}�_8o��3Bhm�_e>8F�흒�'�=r��}
[ZKúcOe�5���szPʹ�д�IN-�<I+����}�V9�}jὧ7]Ɩl<�m�p�Mkv�9`r
�a�b��F�:�-���VD3�8ag��s��UE��eS�F�×�ʽhj :ᐦ��U7�%���$t�l�Cw���65��e+��Po΀��Q�1V��HȻj�I�/3*9�c��T�z��c�o��֞� R��^kێAk��4:���5
��RM�H�����A20sx*S���7gmc��2�0IǫZ9Z�����(�"0Kdp��a/9�ےF��I��1��ɧ(n��ۊ4��*�Sg�(W o1*qM��[�z�a�jB0b�r�T��#vފ����[tFR0�-X�VSĔ:륓����8��~�'ܸmQ�}sA��x11�w^YxW\�b��u�7�Y�MoX\{GV;�!�>a�����)K�Q�
�ȳ��{R���G^h�\�iͭ:�[+�*op�����R1X�GHz�Me�pu'�ؚ�ݖiV'��GW�#5�؎l��3kJٳ32|�(�5fkq�/�}��Ki����5`�y�ǷU�S#�F�dj��3�Ds��ؽ/��
�ѫ����i=H����p9�yԔ柫���"纎�yf� �^6*�
'�:٭�.�Cf��)�$uq��g+ű�8:�RH�ǻ��J�ވ�Cnb��SX����zG=C0�q�s�ȹ����F��l=��5���2D�о�1{�`������p�H�W`"z���	��Ӝ]B�O8+j��v]�o�^\�v�y(��b�C����U��=��k��72��WXn�ڝ�x��玆r�Z�hM�w�"E�u44"p�F�Fm��Uu�7,\�/[:Ճ��n�z���#@��?�q�[!Lv�:����Dwvb}��V�%�L��A��Y�1ܴ�!�݆�,��L[�p�2*��	�0e"1�>�m�sVa<�v�wr"$�:;��3o��f!1_���N���9�������t��H+)Hxr�����Z�tfddt�w���$Oyw�r���z�7���B�&#�u4BiY�`Śr�������U[�l�M>N]�,�I[|���32�:H\�k+�)�,u4wP��ؑV��H���MH�ѡVY�vqҽK$�n^��i�P�"p�yBۚ��5m��`�)݊����M��ܺ ��1\���`��M�5���tn��͠��-Y�zs8���`��UՅ�>����Lm��h-�p���̯c�o(E^4fem*>U�+����wf�챣
d��T��9Tu�ָܨ�P5q�8��MR6�B�M��,VU���,�B����R�R{�ڳ+�`����Q�b�#����w^0�a��D\�h`��:y�������ll�X�=�}�:�lW����8��{��(>�����@��TofR��91�����B6'v������@��/��b�܎�[���w2�q�`�n�#d-\@Mk����� �:�U1���2�nw� ,��x���拡��]@��[����L�Vک�u,D�9kO��|�^��n�CB��ݽ�r�Q�ap�ԟ�S3*f^��o���y�#��#bfjq]X��������k\����R4�Zr�(���w�~S`<=��Cvq�;��2o3�5�#�|����F��r�#��C��cO�F������&����^]oΑ0�'�s�>T��e�3�7���X!n�,�Z�o�#[<��o9��RQɎ=9��n�r�1k���"MTnq��y�������M*k4�v��w���=��+�W�׵h�gq�{Bŵ����K[rf�.<�����'-��[���I�����k���j�����o[�IH�`0�>[U��c=���B�&��
�6$YsKD�/��]��
�7K���4J����a��#��-	���~�+#��mvv�ܞW&�ۢ���z6��o�W&0������Ou�ɍ-ƟgvU�)K>a���+	�7M����c����ײ�	�Ȗ�MG�sX�	��a��4#h>4�v�Ne�-��KW��uyx3'2מ��^ ѼH��!�g^�/s�Wp�����������9�`R>�qG�3o],��m"�r�y���w^S�ܻ���H�H��jKo}/f�+y��s/��}3���T���.�HEGT��G}ׯ�x�ݧ6�����u�V&9.�=�H�=�1V%���+�O^1����n'̓��3AWu�����vL�xBYU	�Q�ihȗ؃4����w������9�V�cա�=�� [��~8�R&�Z�d��`g^ͮ#�p�W�wW7���t�쨟H<
g=o�AG��%��,>#��E��j��ol>es�0��\%�٭����Uv$�����X��V��:�o/-�H�g��<�(���6v(b
�c�*�a�u=}T�k�c�{&��.`^'J��s��f\4٢�4�ˊ��ֆ��*�;Q^���]���	9𶯥[sƭ��!eH��W���Q�}8��mn�=YS�����f�ʹ��XA>����C��N�m���{�+kێQ{;&����WY�/Z�m4RZ0e3������F�G7��' �v�O6.�gM��W�Y���ff.�|�!Qv�}��Z�vE�2w�_r�� }{�7F=���{.Z=gV݁w0�)�om�z@���h,*���3s�ex~����R�k���S�c2��r�Oc:2`���rw9R��ѷa$q��/Wh\��9gqQ�I�뽣8��[8b�nR��/��T��P���t�˩�w��N%�d�cX��~�e)�YTFS{`��6���7N���g��B>���Ðɠ�EW�ȉ�Ǖy^���-��o��9�0�n��w��7Ɨ^��JO��\��|"^��u�o+v��nL�Ln�]��1Νh������5S��v���� r��5�i�s�BoeI��GW	�y��G6�O���1<���طpj��lRQx����w	失n��8/D$�q�u*������h�H�Ǻ�����Xշ�qb��pv��jcxZ�dl��χ�F��(��].J���[�|1���
�|-��q�5��E��Jz�	��9]����0��N\�M�5!Ϛ��/��ӱA�ȇC�>U�eX�{�Ϋf+(#uXu�f��-�is�>ל�e�F��AF�dF����K_�4��v̑��Ja���[^^Z�e,�Ɔ��0�V�pm����kހbҽIe$���T�al�6�J5�>��#
<��6�{�-^^	�[vM@��	�"N��w�D�Z�
̛4WI���(J��S{��1yk�)�N"׹��o��ju[Xrލ�n����h���[��wk�g���͸�~�d��:�og��g��+��)�2x��s;�UkՇ��{^�{�P��j_d'[h�Og���p�A�U�D6����:dv�xO6�̞�gZ���i<�|�S���ASGqࡒĊ��H����C��٤�:�V�H"��G1�Zq���"k-I�ܝ���w�t�k�]��\�SjfSJ�Os���	hD�CY��wF鸒D�Vv"x�<���`�ct��x0�"���ɍ�u/�O��P�eo���R��ż�1v1Y ��t�߶�V�	c#U9"�ʣ�w%��<�?`K՞���eO>�2bgMV*�te"�3x9E�Ov2��m�&���8��.��8�Q�مJ�1�y4{�l���_-=Y�c]�c1��_F26��4m��1w�� � A��f�w��l5Ҋ�a�mV��Z����ϓ���b��ɕ��!5�xOG���FG��3�S��۽�S��ތŋ�F��௱(����{�����-s�!�o��W��� �MZ�x�N��Ĕgk��w����u�,Ob7;@!��҃�w��wkW"y�:�����]���=�7:�'q��
�⫾̻{�)�a`�#)�u-j��e.S�M�AH��,D��Ǣ3�f2��ӕz��ޙ����������q{�@M�;S�dJ]99+b�yx-�^.+#�ű��N��"δE����[�9dr�i�"��c���2�\ü�țʵ�k�����d����ۦ��c䱀C��=�^/܉k�z�3@����@Z�� ��!�X��ha��׺�m܌���t�`U�M�$`���W�B���qO�%	�b��SoM�y��$�Ua�>�L"�؛�	��C\3�������&�x^����cWٔ�{C� �
��|ĊF�gd�͟/]*y��kį��W���L�ڧt�9��E��\�l^��@&<�`�us�2��J��W�m��LWY�#ڲq[S�L]R����yf�ou���zx2�li�Շ�Dx%���~3������*��"�=yFO��v��^��<�`�{i=]'��#�r��|�|z`�-L��.�|�;�5RC�z��-BZ�|zٹdF�֛�W]�@���&���W㾦��`{ң���	ռ��nk�UuX�,o���ɽ�N;y!�v�FN��$���o{�󊧡�#֪ᆑܷ���lJ���m�w1 ��lmmüO-����v�����|���gm[�o3Q�W�H��uY��[�O]��
�.eIݸ.AH��Oit[�ۂ]�K��B���������e�Ki��nҚ�q�$�e^��½�`�ݫp�(��i#��k���¢d�A%J*`�k{�fu�;4Z�Ocpr[3]!�����~���d��t>1���'Mm�|�;a��2�fĭ��O:<zH��'�i9:��89�v��I���װ�i��s�������B8��V`����65H"�t�	�9/�v��Oϻ�)`t_�����Ռ�E=O�M|Q��;$�x����qPR����V�]��KN�sY�]�Ab�C�_
��ã���"Q��������2��!�o��*pH<���1�e�t�y�(�/��AX.���� �W�f�$b�TϹν�yٗ��l�S�_d� ]뽇�;��3�S`\���8�m@wR*�'[:s;5����G�N�����t3݀']��l(�g��D���8u>*��w0^�c@4p*�n|hd�uv�.$ٱ��-�u�F�Դ��pO��&
�3�̔yt<��������ڄ���z�`R��:���6(/j��#bF��ܼ�[:�
���AoYH�����+kwlc6$h��f���Wt��9Gw�O

����C+b��q�h�Ωn3�����p�yC/00r0hl���qLhiVdٹ1����:Ja��<�)�6��v��i�Of�����)����(�ټ#h���SZ��(�8���Vr;8������zU4�]���Ⱦ b��v����t�
a%��YÉ'ֲ��l��w�2�!��K� ��V���`{��'o������v!9�֝����c��i+}~��/�Ϋ(f���z�bҎ�y#]�|LL5������3�f�ӗ�)����CLe�D�%���G�\Q�ޘ\�)=�Y�]��+x*�!g��HP����X<%Z�'r�+ �-���-��Z�.�+��βŢ���76]w:���(f�U�{!��,���_^轩�e����W._N��9�y��6�{�z���{��U��o��ڿy����J �6�����҂�#mTF*���0mmE�X%�QUF�"#2�
�D�k�5,�TX
Im�VXUE��["�1bV��Qk(�E��Z�IP���T*�(��`,�(�[B�U����FQ�(�k(��Ym+*X�J�B��e�Y*R�(,�R�"��h��i�e�kbJ�J*�aJ5h��E�Ԋ�P��ZPY+F�RT��ֲ*��`�R-@RTYD
�DDF�T��T�dD
�P�b�jU����b�j,�EF�T+kdU"+
�T��ѣA��D
�¡Dm�b��b0�(�ek+m�DQT�+*��+aZ���[F�F�6�+"�X��Ь�YKe�T��$R)R�R�Z@ ��$%3_@�W�$�:7��/=��ʱ睜cڍN\��<k�T-�+��aWӀ�qW��yC4\��뾽7�އ�-d���jt�ٳ7؊#D��=�%^s%�!D���K���[�u���Ҽ�W�k
�W-�� x9�qC�.���`�S]QU��Ӣ*u�ch9��&���aM��(Yn�E�:ٗ��7���\�h���G�G+���A��:ݸ��xE�}�T9����л����c�,��}TmĶ=*{I��/F��W��;͹j��Z�7�W�XGԝ���w��z9X���;VMK׸�39�lC��\�{_��)���mwWv��-.��o��\�������RK��xڌ	=��eZ7:X}�㨶�JZ�bmuvjFM�r���{�a��i�Uv$��=�Ú�}�V��:�a�;W�dӬM�އQ�؍[]a�EAPlpEW>�Bo�G���ޏ��!ݵ�3\̵,��
5��uŔ�\OK�tf�۫W��C-��	F�>�£���tզE��A�-��ѭ��A�h�r�Hqp�.V�vA��[��լ�jT�;n����1V:�wq�Rd�m�Z��Oe��K:y����8ko��_Fb�Ў�Q\����q��hҰ��{�z��C�
lGjܞ!��*�uN�C�턡m1\���,k��BʑA��ߝ�j��yp�	�j&yt��Ǽ��G.�i1��q��o�3��i�)zG8C!2��NՌ�z�G��: �8���G�{j��0���o{f�BҘ�{���
=6�>ʸP�5���Inh�Dt�Cz8L�0���۞��ƥ/y�����	CY��������eQM�����;��꣙U��k�$"�!��ɠ�EW��N�<�ʻ��Y"b���{��u��U;��ǥ%3!�L��b�'��ڣ�w4��l�u�nw��^�}&�x�n>���<��=X���XΪ{cڣ��l^���Y��o�6�N&����5ܑJ����L�}���z�_̛{��3.�yqqL�ߞf�&������(2Q��.�c0���1���Ԧ4^>s���B�͟����7y��1���@�� ��25�p����5���׹�e�[_���E������X�:��)��]�Ӕ-��ю���xl�A��HbxF��:_sg�=�"�����[��Ժ3�CH���jRZ!cݾ�kͽs��P˃�-5�\�䢼�m{�� :�:��� ��s�E�H�T�C�{īދ�J��b�m�4����ʇ#૰OX/���������L�FO��_J�ֹ��ջ���N��#�C�!Wd#鉸�ݨh�M�|��[��ߝZڧ��hg8ҵ��4�)k�M	��yyZ�oWMU�k�Ի�?Ju�ˮ���n�Y�-{KPm��e�&�,]����$�}�G���������X:�*���K38��ꝗ{Ja+���d�O`W0�ֽ�} Ϫ����R#3�IH���;3
p���2�S�y���Ѥ�P�U��^��5m��ף�+�X8G���P![s .a���<�	�ӊ�5�Yk*��#}�ϊ������!������Y=L�E�,�_U�Q�����nv�{5�~��nq�*^+��y�-���$�ٲ��A����� d,{�W�Z�ۈ�^�N����$�:���P����1�V���F
^�GɊJ�C��g�-���Iҋ�F�z�	Y�c���	�4"��dD���:p�l��4�����"���y��x)����DfkτT/eu3�t3ĺ��St��V�°�&S���K}����������F��`�gn����ְ԰�I����3�M� K��x3J�Ȧ��g���1�,i)r�5wm��Q��s��=�=�lVR7;@�-�p]�3Q�ۭn)��T��>�fo����b�V/K@����b"�YQ��V�&��������������F=Y�����v��������P���Ꙝ{}��e�κ�{@�����3�+W&�؇�J�l*̧u�]�mF�E�SJp!w*Ý�@�W�>{_w]�G����ӥus���d=묘����ݬ�^�9�@��GR6^���9\��l3R����fY���,ݳT4^�cޔQ�G_eVm?7�yx\�Z��jA��.��:�As�>��k'u`�X�Ȭ��B}���Е����[��~���-���گ$5�!h�j[�a�zh�'p423	ʹ%�}���xD8�,�
��ʤ���z��G���	T]SZ��W��P��Nx^	5Q���n�iB�J#v��{��fo����O͝������V���H3����V�}��s*�kD�u��:�z˳�S͟7V��L.hn;�}*E���Ruvjb�X\�6�Xm��u0�
^��i��CY�Qνmz%h��v�r�&+��*�������"����5�FF�eR�m�Ѻ�H�/���Mm��+�j��D]6v���8P����'�,`|��|���
�hEP|5��ʻXn�>�B�w���	����A�|����OG���gޕ{A��s�sә@���**b�������#2 �>�R����Wn��4����Q��Fe�R{��ӭ���������%�u3��68�В�u-�3m��}�q��v���@T�}"՚܊����L�����$_�	q���P�*U�
�^=9��M���i���(������v�]J�un,;aٜ���NI���_�y��mS݃�#�;Vf+-�(e�2��̏"�fEb�u)[�wi]�5z�˞1���1Y��q�";n��ozʣ�DK��X�'ݰRlQ,<5������� ����m�rֺ}���*�Y�j��:�o+Q;��j�aqT8"v=`��PM�Ҹ�G}��	(Ef�u�3Z���~i۸oi�Sшr�C�S��U� �F��V�ꮧ&�;q��*�=�J�U��֬�+]�	�N������е�"U
qs��o�73Y�Xc4�f�z�:՝��w|�5o��X���P��B׵E:��:��S���sU��-�l�������㮂�}~L�"��ԔO9<�w��f>���L}��!=-���e"0:gݵ^�m�:�Y7sϥ�c�u��q�:j	cy�m���\�8Q�K7��<��	Ǳչܲ/�uv�Fhr�a�!�h4���[k*򭹣�QM�	=ݮ#fv�m�#7^�u�i(�_;pe;D옑���m O=��u2���̀M+�j�5��9��^#����-�E}�[6e��s1���tz�u��X�pJE��%`u�f>a��Z4���m	&G	�o5Z�U��̖v�3.v��(ܫ�mबi���@�c�y6#���	��*�CY��ǕyWk�˂7b�P�Y{u��7���릫�{�@��OFUw;��Sѳ���b���׏{.�2%.��'_��"����BXΪ{W������,�-]o:5�Uwx�:X��frp�E�}���j�H�H�����w����_F��E�^�­���+)s����:5�E$���W�2;R�9�4�B%-�����Pv/O p���\n��'V�����)+�F���ƾa�bv���ʇb�N=b�}�U�[Ig2�㻦�!��Xe25^���|>�V�Pl&|�pGʻ٧ۀ�W)ذgk��o��>��u�V�����޺M�>Sы������g9#b�6ݧʐ��K��V�,�Vw[��	d�Z��~-e9���xn<�d��%�Ŋ�����,���"�	������ō4���o�N��yڧ�T�o����wۼ�>����٬n������B-6��y{��R6�'���t�~bҲ>RM�\}��b�̌KDlͯ��!����Z8U+�J6�~���Kn�0���{x��Idv�Íߎ�Vu�Uo��ȑ�6"��b��,�ِk���^�V8���#R f2���YP��F
�ўGr��<�XSV7���W��m����������㌙���ي�ܖԉ�a�H�-��)x1�i��dD�ZʼƆ� �e;�{���,n�G��>�(P�繄����`��M�5����q�\�ZыķynJV��v��:є�ۦ"���ɍ�0fu�j�s�J�����IP��,mn�ʼ�v��7�6��-���g?!\�N���Z�!	��c���+�a��4#h>*wI�� ���Ha3Ps�T�',���8s���j2��c�����I����:�u����-�[��.ml3K�vm���f�F=������W������q�b������7�<#*틷���Ʀǳ�<����u#P�v��v�H���G������o���0�v��:�N�R�#I]V�$2j���\74��p�e���݄��B�*ooo���X��[*_o1���WZ�`2wys�:��v�� �����魿T}�N�齳y�aaX�#8&w����ǫ!wW[}��P�Tc-�99�7��w�R�V����a�{/�vr�%�v!�ҿ)�;]=���ݫ�w_^$vF��v*����z~㫸��9�1�͸ɍ�{g&z��n�FC����J�G�>��Y8�����*R�;��*w7��K2��n��\��~T�j.�a��Gjх�P}8�cM�QlN��x�=![�"��>}U�t.P N�W�>8�0�l��o�2��{L��ƺ.O;�mvnY���6CAS�uf!�ȣ�z�߽S���Yb.>(��0T���2c�[�!��,�K@�祟Wt�Z�<$���0�5�A�:Y��lA���/Vؑ0�ʤ���Jd�f���7�Q_����([�[Z�|�"P�`l�]~W/h�~�%���.���ʬ�x��A�M?�NVVC]��Ai�yV[���|�̺;�3ʒ+��+.��ż���t�V)��͌��7�}��Ɇ��sX�o���2@}���g�"osOp͔5�62P�;qg:��p4F��s�h�2^�\�R�ɮ�#�fڥ͔�,o�(��n;��{�E���.���6�RY+����jhh��|�7���U�K���I�(k���t�Py��4Q�ҹ("al�+�����EEg�O�����MA�=���G�}���`M'���gFK�z�#a�bC�X+�T��dWzٸ��ٌ��7d�A���ш��hw�߽����6����Ô��N�
o�^H)k�����O:�@D��,�͢����uo E$��F!�Rx�����^�'��ᚫk�DF)����Ld=W�W�q�o��:%�!�2z	����8
"�B��G�.x@�~�^d6�����/c:�1�2K��6�B�;s�$tmmXj�I��}�}�U��N��^@��-��R�T+/S��Y&fƤ%�򈭎|ʩʂ然z/ZGJb�m�HH9���V�r��]���/q��,0�������,=�u��b����/\2N���-8��z��;��Bp��E�g���dn��T�'��Z���Ϣ1�\H�M�;{7�D�1��뙘5P�|���p���]hl˾�NBIO�����\�����_Qv���:��\7��V����u�.3��۩n<	h�+9s��tf�r�6�0���;l���M��²t��uUoA۹�������ΞwQ��/ y�^z�ڼЍ��X^>��4���c{��2�ge�/6�=��������Rx�xV]�.���/��kU����k��/�1}
;���׽�ϹZ釷�U�X�$��k<yN<�����$ 	p�VKn�A���HI�^p�1p�HA��8��.pU��o�n��`��u�����82�8�WkFIK,q�{�b�6�0[�`���ĸ:�;dr�GJZ��N�i�󛢛��c@��)9�������v�Z���7�ɢ���)��4F]-�T����aXl������H��ڳ��a7A���+��j�
��ɓR����'N �}���X=�x��t����Q�]�0�'�+>��.� �n�2�Y407����m�I�����y͡��0����G��Rt5�l�S��|��@��ʛjZAܡ�V�+�4U����I��D2\���S�qd=���RA�<ी�ԩ��^gt��^Ҥk��x(��V���u�q��L0FZ/.�a�h�JT��Wξ'_�()q��E�0]�U��b�Tfh}�V&�ơ�&L-03(a���@�˶I+�:n�A���e��lF2O��wt!?w׭���������A�9��z���UH�r���x�i�y������L�r{⚅�hJ�9����~	�;b۬
��X��o��w�EC�ﭑ�#��y��5�6�h�~=zR�=�X�\�9e._u����{��7Yi�' ���ffDF�ͦ�b�E����T����A�t�+��.���f���77�U�n
�KǜպƜ߀��z�p�kt��	�K	���pKo��.#�5��M��Z���7�L�#�Ԣ6�ZOzD��p�+��|Xyo�<V5[<���R9!:g�ʀ����H����
Kql�t�D�f�W.���[��^��6��SN:ԳK�]��b���g-~9z��Ю&��ث�����t������yƁ��)p܎9�,��$f�Yf��Q�o]iGp�%�m�M#m�ޣ��4r���wA}>�4�m_J�Z�� ��B�r����ДrS�CE���鞜�޵����V��/�	>�p�Pe�oأS�]���ܹ��B'��=έ����:��Ȯ�L��d5�Eu�#��f�=%�2w�[+i�c�7�����,)��PĜ�G/o�����н)2}!�t]����I�ĺ�xS:�Zz���4d��U��7[�1@^:lqx���I�6�4_��)�m�'���ŊCh����b��*�F1-�k
���b�%�XER�Z�-�-dmRVe�VR�J��U�m+Т-Th��J�V�IV�+Ym��Q`�*"�P�"2F%k"�VT*F��ȂB)Z�
���
����A`"�
�E"�E�iFE�j��k"�m�E�(T*EP�V-Bօdm��[J$X���E�
��)P��ʋ
!Z$T��
,Z�-�jT���X��`�e
�ch(�AelH-B�6�-*E[mH�T��,-�D��m��`5�lPPb�J5�@Qm(����b�k�V�ab��`�"�ID*+jԨ�-�YZ��,*�DbȌ�����[B�#X�`V��!D�YUJʨ,[������$��2���|���8W
�'�'ǌ�8��=�wĈ��DV�[;gVW7�A�:V��I2�m�2�$����U1�+��z˃��]����F:3��N��j���~�{�����{�X����V[�H�K��yP�/�	�^���
��0���mϫ0lF íb1s7 us����P���U��VmS<ú�T�੸��i��sD�j6�#Kˣ��W:��cQB��옃�b��h���È��jt�l���5�(�v<}�lNi���O%2iJ1��H�,D�������!�CD?s8�Jǖ��;8���i�F�Z�0�ێuo:����5e12K�7�!G�s��$�;E�Ae�Ƶ��T>�=�Je��v��m`Q�����Q���ݎΣȨA�S�קg�Ъ���^�=�p����75�y���	�>����^��l�_������2��;M��]�Xn�Ĺ���u�J(��2�8ٞQ>��d�خ'i��O�<��|O��~=���Wk���Ou�f9��js�a�t��y4Q��|TIb�i�b��:�0E��H�g��|��:m��G�F�zQ�^��1,~����V���լ�Z�{���H9������>���������M�;��~�r/y�u-Z�v+Nü���kR�Q��: ��]�kI+,�$X��<�Wwv�7ɛ��n�'�[3��-�=�����[Ǔዺ>����wm2w����:%P记ݨ�n
���AZ�q�3�bi�Gd[]�m d5���Λr��^,���"����)Ezf�t'�'X�OL�ҳ�:��9$�dêpSт)NGX��:��t��=�:w%�ؘ�N����;���x�6!4ODm�(�\�(���)���8��1�����V(f�f�[�q%�t¾�Ȝ�!㮙 c�8>��'��mW�נ� �g��yB0�C!�wqw�w$�Y}�.�͍a�[�k��.({��u�#Vr����~&k�& R�td��[8�	��Į֣��k��*��/�<f,�q�S�ڽ����f��"�ȵ�i���|�2�5��Q�Pprb���;�,G��l7��.{��>ha�6.�B0ƻ�E-��ֹldk	�_Z�lm;�vb"��`�R�2Tz�'����-������Oi�!#�C��Q{r}e�t�W�<ec���E��Q<���go�`�|#��~�4���Lg]�b�U��j��2bў���|=�7�K��{�Q4y�x~޵�ѩ�Ǯ�"��ZL�lx��
?S}֨Dnozӓ�_i鴵VZ�yb� _]Y�.�ĲL�CɹXQ-#�?r��wX��rN�:����'WN���������\�4n��қ��X��n�����#H���a@�e���wk}94!]�R�{:[S���?���!���>>�>���e�_��U�TAq�z����fe���o�ٴ��~cZpW��%������m!_5du1��8�.���-\ž�y}�g����)�!h��J�cc��{_���;�YF��\��y�Ž�oc�G�A��!�,�x�W�v��B�X����w�0^}K�=���c�S���J0jS�h�*�c�T���(�zv�t'�R�����8쐄�fP��3q��wp�{���XL#�l�B����U���A��P�w�}�uWGG�$t���kgI��d��AJU_p�VJoޝ�d_���C�"�<!XD����\E-��&ԅ	���:vc2� ����S^���˰�+����U��8���֌��2xl�TS�"Һ7!�Z��yF���]%K.V	�e#�}a�:fԸ1@���K`�8#$�EQ�Sp�in�u��M:��J�_�s�T���i���%��h��4hJ���,�ٛ~��k�����v��o4n=U޺�ぇ����qmh����q�V��ߺF���o<��p�<iַ�(���N����yK�<꫁(ӭ���(��[s����p�Lz�b�C�j��էގ��cX<|Q<��{T��o���[�#��9��Y����xI�X5#W�c�����yp��ER��C�S�Z[DDC^mO�r���ɲϼ�b[��oԻQ+�z<�o�� �h���:8o�����-�Dh�h:X��DNIr��!�Uј|g!�}�_e�{�ҡ�`�֛�^��_�sD�v�W�ހY������=�o����,5V�Ը�����6�v���e�궪bDd���><W�9^�.}��'���u3�m���2��O���թE�VHB��0��~p}��͝��Ef⛨��>jbk"�H�b��R&�]�Ū����}q�p[��-a�ɟR;��@�5����Ϻ\D��Tz=׵y�Z�vo����nT�a�Zxk�d���\���T3e����K[�:tO*�j'�d�z�L��!@�=�a�7�,����+����4����{	~���Ȉc��5���Mꀛr�����≵���լj��D��6�:�ҕ�c�8�]������p�7l9��Vo��W�U���\�WK�_U.��.^豻�����4l>��Ń�v�֒���1�v�(Ng��t�r�6���v.|���ƏZ�go���4��Cy�^��������j����"��x��-κ��塇a,�ˍ�KV%iT��P�)T���=-�2�L�D�p����s-F�Э��rc2��7�˕�]�aޕ̗:��C9�Xhvz\T;�B�\���x�x��!)t(����R6f%�{�njI 5�*�*Q�c��S�\�K� �ݒ�>'��n���@�4)�}�A�9:�K.�Ǣ�yo�h.��e�׎M�}��~zv��Դ�K���Ń�z�8�p�3�1�����}m����\��b�g�[�� ~����/j��^L�侄��U�����P�΃6U8�<��GZ��Ng�pS���g+�ںݝw����y�G���E.�!�R'F�0�O\Nm_,^)~~�VS�Prn�����������t`@r���7�*��#�"���qbkN칡^�1gwdt҇�3���c[j��q�U�b.)�����N~�k6����nz|K'��".�|�/;�nQqJ��en;'$��&����0�KesԨ2�&|ь��;=x�.�H-_Q[#������[b�t��yb�Ú�κŸ���V�MٛoD1���w�q|�B�	r��j��A`]��L�l�:�=j�f�I� ��pйޡ��~��ݎ�jvx�
��,e�u� �$���{��Vt����׌ˬ��� �Tޜ���D�����Q�wK�|sY��wo����o�֩��Kx/���3�lWKp�O���v��'ʳ*�j	8��f�>B�S��r�-��Mg�{g�Hdކ���`�k�6�QXl��r���9��>c.���
]�d[��8"^�S��tWXډ"�
,E�
���yn4����O2��K�t�AR�~�+����֙�VA\��/ݗ�.^=9gk�l�w+��&z�K&�0�Vv�:�=�w->>��ޱP|�r[{��F3l�^>;�eYG�w�f��{:M')>6<s�C�8�v�<N;{9ٮ�B�]y7��<lS6�9�Eԇ��(A�s'�F!1�<�KC�AT>:�jϼ�_<{{��7A�����*�|�(�7	�o��pc�ԩD��!�����9�1�{>���c��}�Ę�M72�)���mS;�OZr��ķ�����\i��)ü�&��-��j<oo���s�v�7�\syP�]���mEEh�d�͢��5��0(5���3eV�=���;��zuݶr�J�z�w�:�@���lm����1OG�Onf�9qĄ�'e���Ϫ���q`:'X��-�s'��VVdg�����Q�̓I,��v��cF�prb���z�����`�d����P(�>#��Q�r6�U�����ynH�=Rb�iqQ|Q}��A1
��sE�L���O��AJ�,T�r?rFg����Y�Lٮ�'�]WK5~��V9�:�U�~�j'��~�&����-�0��h���_!=�d��"�B鶁ڒ��o(Y�������嗎e?yn�x�p{!��c���6�p�cǴ����p{�C�p����\C�Tc\6�(Y�Y���9u�MEcr�C��!ߛpaÞCz+���w|�o�"��rb�V��o�!{���z�ʣ�FAΨRvC�R��+��;=�ϯ�C��\�_�v3:����QK��q�O;�͵�L=.=���G@AK�7��a]�񅎱NJ��]m�D��k4�5�������O�('���̖�
��/��5e!�r��a�nP�&R�9�\�p,�>S:���
�?(�0����I�(v�����үg���Y����8o% �6���sw\�I�^��L�
�ѾI*<��G�*IS!����u(�����%2��ς�X��{#V��W����ǥ��[g�N�Ц�R��;�}�Y����h>vMy�Ͽx1������S��?6R�� {�߳~(ؽ�=�^���d(^��`��h��u"�Sr�<+�{� �����43*�����V�>u���XT�AX��Ne����F�W�O��D\�͑�����cq�֥����}8.vV	�g�k��2*�abN�W�>4@�۩��3a�6�a'�{��sVD�׾��{�:�p23$:��(
����/�hdP2�����9��r"I�<�f�j����g�U�xօ��|�C}L�K: ���9h����A�KzT��&/	�	,�sȤ�Xl�,���%��P��]Z�~󯼉}��Io�	�nm��ެX�M��1�a*��RCA�s�� ��W����Uј��,��,�U^�9�M`o��eT �#���"Jd;��^Б{�|�&�V5V�."�2h1/���粮��v�>����hx��t{�����^����"9=��g�^ט��v�[�<̗9�����{;�ML8ː��s"�s�� ���^��8���zW �����"�ӯ2���o5k*(�}������un��� J��2hs�p�s��GGf�}�e�6m~ħ\E%���{��\.��v��.u�E�"G;�Dƥ^��Bb,AaD>G�4j.�d8;"���ٌ�;�+&�B�.�g�ڕU]�>b�*����u;���0�r�rrvS~2�AK]��W�z�����ʭ���Ӧ����q%�-\�f���P��ϫބ�c��3V��l*�qp�}�y���#��;�#ص/�g�m�=p�(�=�RziL9� l7єJj���w)���#|�qQҫ�P�����R�/�^�����G��!f�I���u��J���rXsnA�F5m:��N�[���v�Ҙ�C�� w!��.�s�צ8��<D�o��E�E�l�
�s�P�������Qh�1��x�� �W�W��%IY�	ǵ�3=8J}w�2�{�0�y��鼬R�^5�Pw?��ޙ����wFW`R�:����ũ���G/J�1��Uh�S�����Q�XW����s�KO��}��u���l�������Lz"gxϝpg�����>V��G�/��O��{T>C�ܓ���O20E�.�;vv�0�Z��"/w���BE{�<,��\�2����~��s9�gwn��αVV=��Ѫ���t>�p^D���k��6Ud��|��{���'%oD��	x����S\�C��?nt�0meN۝�.8��_G1T�BQ5 g6t���	��7�}��Va�i�3�8)�����at����gesR:���G�L��~���x0��U��0�К=x���R��2�k��-j@�K�!@�0��DL1 >�qb&9:���X��L�MTl���c$(�ս���Kw�e�S�Ys���g�FPB2)�̞=��}>������Y��ޣ�V��p��Z�^��c4VT�i��o	�ӘTl^�v	���BR���*w�j�/z��aw�4�|V���1Mw
c3��;xj��ޚhZ�s����c�3�h�&Y!�>sWu���~|e�:_)C`o�L��Cb��[��&�\�Cz�B�c��GH�ETEK��	n�o�P{;EY��D�6.F�F.|�X�u���s��;<��o��m�7&YQ��1�9w��v݇K�ѪvU���Q'��Q~���n�l̵ü�����z~�5dYs�o@�75�ݕ�f
fv��C�y%����$ I?����$�y$$ I?�$$ I(B���$ I?����$��$�	'�H@��HH@��B���BB��I	N�$ I(B�rHH@�Y!!I�䄄	'��$��HH@�y!!I� �$�$ I?�b��L��B��
(� � ���fO� č���ҭ-���� R�%$AJi���JE�P�T�T�$ZֆR�
�UT��JPJ*���R��+d���5m)��e�ZZhm[Vح_vW,�[UeE�m�l+J�`�V�Z���Ԋd,�қJ��l@�i�Y�`��i�]_{��i[6��Z�ZV-�E�m�U��+JmmFͬE�-[M4T͙��ɍV̳Q�)3[-+(ڣm�m�*��X�
mRl�f�2��L�}���Z���  ;q�_vj�t^�=����m0��^�GH�vzu:�U���8��k�wv��;/mޚ�ʴۻ`����Z۸�{���-�U]n�{��uݻ�V�\��J��iިb&�h��k;�5�6��ӗ�  }��׻6����uW{{���۹V��<����wWOM׭-�n橺�ޗ�Z�z�]���^�wtwmvۻz��l�[�o^;�k��[uz�㷮�����������ջ�۶�m�(�kJZ[6ab�-j1�   v����[��bw^���mUJ�2����ܴ+wt���tҥ�W���W�K��n�&t�v|QFz}�QEQE^y\t(��(��/q��@PQEnqEQEQ�w�4m��T�ڶ��Pa�\   ]�=$��Ep���EQE��QER>�[�*��ݧ6��}��QT��ڪ@]��V¶�� =how����h.�MMm��cV�ibZ֖M�h��   ���>۵���T)��yp�j��y=p^��kV[Jv0��T�ָ�U{����@��������JT��im]wlUmT��*�6���   ����T7G�����MK��a�=M���:�Ox�۞�����Z�.��כڙ��W�޽���wSQWv�ճm�����青[4��)����|  �꽾��wm�k�yw�f�u+��q�u������;�*طs��;\Ҷ�n�;ך�^���wu�������[�����;zm�۔�szq״�ֹf�N�.���gr^��R�iI��v��6  j�>4�kna���aUu�o�*��k=���aO,��yW��f�v���T��Egw]�뽭Z���/]����cv]�޼������k��ow��몽��+��X[j��Al*�  7W��j����N}�WU����=w����]��s޵K�R�s[k��I9Ǜqm��Uֳޮ��W����u)˷vں�\�����5���f�ݫ\�w:������Ņ��*хmm��  ���Z�W�ڽ�;�j�+]���ֳ��zk��wj�Wm�V��u5Z�q��5{��wi��^�:�J��t���;���Cm�wmݴZ�����������_ "l��%J2 S�0��5M�h���{&I�T�M�  E?�SL  �~"cUU 0  !IT��� h�O��������k����?6{�SԌ����=�5��z}��:�/2��Q{>�y�QW�QE?�"�
��ED��* �
 (���2���#���k������ۃ}I����	�(`X1���%q �K��[��2�F�`�nM��r^�#+5ް�Q锝Z��]P+��%�2#��W8<����ѣ�8K.lw���P5Z�V�gF��a�kĺ�y���0���=.=��l#\�,0n�O��,�ù��S�V�db]���Jq�݃2lL5�^�<���M��l�rCf4p6}٭`���	t:@hui�Z�
軻2RN��v-�k2���R�r����Zk�Pь��, Z��*�0�nC[���4%Ք�Jl�Yzq�6� 	�r�ǿB��`8w(��N]{V>ķ(�;a	0k�<�/I�����`��Op� �(Ƈ�Kף��f�0�q��l�i)1J���8HO�+Ȱ,3>��J�u���"s���f(�4%�����.3/)PZ��)#�Oӭ!W� b�X�1R����DۥZtF��-�úk�H(���)iq��
�f9��2�K��b�W(h�$�
P*����G��yG�S�p�.��B�Xr���l�GH��b�be8������C*��H���E\Јi*9�FlHݻ�NZ�&]JC@�v�n���Wx�N����苃q�v�rӗv����B-�����*�Io0*	��X�e�c�j�E��Zn�ڳ�%7�
r�����r�XtU���qX,��{��.U�ab��$�T�/*�.é�ڔ��+��]<c6n�׀�(��E�-����%�9p��Cgv��Mf���!�E����h�Aln;�.��w��4���J��mLʆ��V�+"w@x�Yu4��$Dk�gv�#�y�h�C�P�Zf���W��
l2jQ�Z�H؊�$���Ъ�;8.6���n��L[ra���C�ᘤB��N��N�gv��hy��hE^�� #�P�X�e�¼�&Ÿڇ#v�hf�F��]m˦,eɎ��b9�U��J��5�N��9{6�U��ӱh�8��,��H�4��^-�6=CU��&�E݈�.B��[AD#Ӯ�ܒ��d�n�0S��9Ja43/0b{�l���âG�4������f�Ku������JV��/,ŦyY ���ꔀ$:��6�[�2a��[�q�I%M
�a�`Hs�+1e7�� V �$X�mT���f��,R ƑH��{��� �!�`�h����s;+[��:F��@IeX�\�˔�4Z�-��I�g�MML{7�e^ͬ� �5�������p��G�^1�b�܏�LЩKsI�R^h�&L���ޫ�f��;ZV@�"A�ݨ���m6��lWhٛx��������i��U��``	��ԭK(gH�Z�
7zp��u�S`�����-��aL�0r�&�Bk�UW[�j�ai�ҫ\ؠIE����Z(}(mkH[ܢ��J�4���&YwR���װ�+PJ��v�c�s�-4�K/7w�5�Jֳx�'b��Z��dD��V��)*�ƣ�q̘3k6�X��iB�cŀn��mhR*Q���Ԧh�͒b�2�U��C�Ne��ie��-��;&��4ӣs6(	���!8mn���5vC�p8D�PȔ�C������QVhB�1��X1�b�6�V-������eAؙ�S��(T.P��㒆�͓�Y6�+�Q�-f�[�Do�-�b��N�h�r�S��U�\�e�a2%� �ܩ���f�-Y��b[wX�r��ò�E��tP�M��I�&&(d�8��v��#��/� V�i��5D)( �:&���ս��f2b����,��r8�!�t(ؖ졙Z��T��j3,B�ѐ�+!�eiz.��h
��T5��]�A>+B�'®�қz�)����r �ȱ�Dh���?`^CY*��hU�B��5o4�[x�Ey��3.���'�Pt�6^<�H4�0�U�g�z�c���v�u#D�=��v������34]���;O-d��P'� o5"�Rp�]*�@]] �4`�.�kr7t�Z����V�TpڥV�5��.�S73�i�V�' ��u��D��������S�Ŷ*+GeV`��Mg�Prpд�k��ZG�w�u��j�n���� ���UJ�;��zʏk�ԻC�,D�I�9�&�V���X��.J"d�mV�F�<����րQ�4��7uo�z�#"dcB�B����R�sa��ũz��u�4�J�3$е&&T66� ��j�͍�0-�`���aͣnѬ�Oh�yt��4�S�lb������6���^�xB��>�Y�B�5qԓa0e�;SNQ�������:[���eJz@�v���-��J�ED�VU�(��D�p*F��L���\Lŏd����%Gq-g�ʧ�l|O#�+3�a���(�g�N�Q.�e�4�Ȃ=�wY�4*$�P�zr��r�
;Q_����⢶���
[��nn��ڎͨ��Y��ӟL��B��哵W�� �*�L��2�a�8�f��n��I��8�`�DU.��h��5BmX�d��X��.�y���,�]��H�*���W��3�؛I[YHS5n�X܀�F�'����[$�J�Ά̄Q���8)���E�³ebw�d�E�%���7�XU�p��ҫ4V\'�If�`�@��^�V�ɂ� "�֌q�3X�v`�Y��D�Iԟ\��*j�E��L���$�mP�oK���
��%X㹙AT�Sn��?mH�Fe��XJ+��I[j��ds6��/�\wA����{�)1��YH���h�f1 y���.���e1%*�vK�c-VJz�ܒAt�)L���q3��^��^��ӿ�cg��C�ںO/6���b�pJ%�R�^#x�T�ݩl6���g�1�'�1��Gn\r��8�(�ʆM4��J3mu�#��6�ǀ�nF�mmҧwY ���Y)��n���׮��n�Yb`��l�ؖ�S��NY+m�r����zqP˪��$ ֱ��D4����̆�n!*˸�v�^�U)n�JP���*2�Ѡ#Obr�N
����j��-�z���h�lа�Le<�F�Z���L=͗���Y�L�����S-����h�i�YJ9Kbn� ��	J�����4C!G]�k2�C+I�������7e�.��b�}��J�E�ܰ�C^V�P��$sw<w�闯j�d�e�5 ����,��^��V�����b�F�.����=�Ӎ��G�B�̼yu1��rn�	��E�.��%��`��T����Y{Yzu�1fhA�H�Wn d��]SJ2�Y[2�j�3B�-Ɏ�J�v�n}�E*�0,����
V�� ��,�ۺ�R�{.���S�ؚ�Q,%wkFƌ��˺�}0ʔ[��(�+�[�e��O�i���Om�m3[JfL�;��T�^XR�k@��IB j�'"��7wq1�i�a�))��Rl�Uay*Ig �]���(�bl���4�F>h9S�%V� #i��i�Y�CfSBt�
ٷv!Wp���GwV��a�8j��RT�ܔ����Q��%^��@���ӻ��k�8����z���.�n�M��4��p9,iL�2i7�q �7m�	ѯ)�t5��c��q�AS� !7w)^��`�R�wN��jrV�,�A-��V�]��Qր��8�3R5Fw&�X��˫a%�5��*5j�����U��J��K�Ӱ�t�Yw��4/c��ǈfXL��V��ә��V5�Y�,$#F$kRb�JX���Y�]�9�l��=� K�Ǚ
��R�3(�ð:��-��8�eǪjҶ��X7z���c �ĵ�EAVV��Orm���ԙm��a�v�]�����t�+�W��;W%�yF��nCM��g`��5��a6���$�2[T����bE.�T�}���6�5��P���!6!<�r�t����gr.A0n�&1�uj�H;6c�D��ES
�d�nI�9�QC����˥lf�=PPԍ�@��B{��_�!�s�6�O@��������.!�ə���CL�Zf{N��������ks�Q�/A+۬���8,,x�@��Ѧ񚗂�]��۫�2��c�Q5��h�'�,T��+u���Zw����h&�X5d�%�P<�@�h!����)E�D�mdE�RmL�rcd���>-�%�y�{^Ӯ�]�q	1����XE�������J)E2�h��wfn١B��c��R�\�8b�)�*�w���d������­<�gKVa�A����2+�b��oN�n��WZ�������y=t��g,��܄��Vƽ��I:[���vfTn�SeebE^��Rue���ԛ�4@��2A7zB#-+KVV���g"�f�[ڑ��X���	��D���/-hĎ��+e��B�ʁ`����d#�`РCd�,h`&�1�e�@��Нu������� 4v�%�Z5j�@�lM�p͖.n�
�&�������
�Bx79B�*���ǘ2�I�U6���:B���;Ε��M�X��}L�`ہGbV]�j�ۦ(S!�z:Ԙ����
�Í�Sn�$������9L�h���9Vi�P��hń�U�������1*q�?\k.� ��߂(X�ˀ*f��dؓf7OS���e;�*�����H�Sc%MZf #�2�U*��w�R)_�.�\,sC�Rr~h!�Lu���)��]ҥ%��V��n�a�� ƛ��[��׸J�~'.n��E&n5i=87Zjn�d����M���\�jS�D�Vf[-�����w�ݣ�S4VF��:S�Bv�	�W�n�����ICZ�n� �//sL�ک)�)i3�I��x(���E�{L⦠�IV��N���2T�+c���VP�����]4*zٺ 3z�����b����+�j�v�];66]����7ύJʻ�d�k��6����#JseC#��[���aԫ ๵�Z����m��4�Y�Ӵ���=�t���̒1V20�U����0
8ļ,:��f���Pl_BjQ�-yw%
��0�Ǚ�j*��'������!��ͧL�H��u��1Xيژ��T�!̌�2`��Q�
�n��$Q��)��sr��>#"oQ���b�ne[vh�5�1�7y�6V1�8���m��Le���ߔܖ��v�T
������S�/%�6��t��f��4V"Jx2�I��ٛC12�KjSI���حS�S�Z�Aֽ�����Gs(=����-�zS�j+� !b�̧�.�N�w�I5���v�"�����dI/���h�Z��	Fhu*\8���>�ٜZP&�
��ni��VB/!�E�AR�V��!�%�$p42��\ƫ�R���&ҳ
5�V���	�׮��4�u���R�ҒJF�6 -7S0GC jy��njFVĩ�ֻF}�S�)��*0���!���օ{�,p���v���
�ER�F?��{#̙{k]є�9Z�ʚW>x�
���*Xz�H,e0�4��D6�7a�W�I������]Z����t��xvS@)�������%ԵLŬ�*m��Q�%.L7EҘ]j�f6��'J.<��B��CuX���p֗-5���oF�2S�kE��P����LK���Pe��{�7xq(j�ri�BV:����@��L�dc͖��v���!�3(��G�ۼ�)"�kZ�*�b�$�ZY��]�˺m�LA
 �Z��zu،X-@`y`S�Y@�Ҵ8�պ���#/$DR�x�����6�<�U7@L���[r�8�٢�ITM�d2%���`����5���k.��2�����[�cɢ�Yt�퇲�i6K��EIy�Bm%�֓�b�B��Y��i�¶Ҙ	����jR�ۧPX�
EFC����t+#��r�Y�A���Q�*�c&�"�Ң5�=�@��d�זҠ�Y����eM7���0��W��^Æ@�BnٳaV����y.���M"��"اCp��L�܀ֶ\۩E-��(s&�J:�%NRf��.���W�[Q�ť�RHhh֬�W*��wC.;� ��ąՑ,br�Q]�0�^C�F�0�8��r��.���hZ7 �-і�*�֙-�.
Yy����'�SG^
�!7t�Sn��-,7�5߾�u+NS�+-�����@ �\h���7M�V�b�r�<Mcٟb����mRu�-!wi��JcnGB��̭�
A$�l�u-�T��(���[m�v�{ �n�
DDU�lJ�h�cwA`���� :ܑ��f��#`f�(����#���4s��N��M(Z����V�1dK(3Bmn���A,Q��n�1��0�1�aV�Z����DH���.Sd1F�ډ%�t��C_>�8`k�D[����=���%D�!���m٢^m���9���d��h��x)�ibY�; C	[jje�f���z�
��Ok�ԓ��e`uh�]�wrܫ#m�+]`e�	3;{h�7u$p�xё$��9����.,�Z������Z[xs��/�����f͵a:�𭚰+�0Lq]Ay�y�]�p�[��D��A,�G�%0Z�hϋ�+l�wX�Ea,�B�^��N�l�],��ŴZI�W�<͵SR��[�0��T����Ք��ȅ+z� 0���4��A�^�ۺ���H^7|x�
�S��:�Uɳ�ɒ> ��M�;�r��;2<���}j���B��U�>�2wz���ʝ�^S��VӮ�l�sm�o�mB��F�9�����-��5���!t��wF�����<�qAn��;~�r�Ƒu�1R�TzY��D8x���W�Ѵ����)a��k߷��j똓�k:j�Ŵ�,�-��:(�Ι�	�ѕΫ)�Zw�)go�*�kx0?{�Pt�u�sv�L[�!ǋ�MN5�ٯ�I�/p��~f(��Vh�rЬȷ{�ų���ʼj���oA7x�U�f<��`�T �Evc3k�xUci����.�����ۄ?ox��#��U��R�(��D+=�[Ri�nNy�ڳ�{F��[a�j��:�6�=���L�]Cݞ"��u��	�7*��v�WIx��]e��Rm��[@`���=Յm�wY�Ӳb37�M��.�c��\��onjs�*+��[�˜E\�����f���g_6nV������5��Z���ok�����$62{��2�6g>��G	WBm��D�XBTL8�'3�g�r;s.����\$*�hd��J�jΫZ"�Z5�� U��*���ؔxQ�4nS��s&�w/���l^�8�g���q���eoN)d3$B��I�N
6��')X_���S�~ɦv�Y�)�7oD8"�Z%dpcD�E-2�gp����ҍ�C'�6��'q`���޼��aq:Dv"�Qض��%
U�2��	�ԓ��9W{u�Α@�����}zy�ۺC9�CUJ��ؐ���s��^X�\b�ی\uj����}�|�s�.�93�7��3(�e�K�J%��DK��M�Tl���ېMUnt���֒f�����x���3�S��t���ۺ,�yvT�Y�����P0�:0Y;_+n�򳋧f�IX�ipn])l�.q�}�潵&ʕ:��c�`�a�B�Q���J��Y�n]/8Ȗ�0��4�w�yY�s��}}��@�!�x^��W�qW�|�pffg]9!l{3t�,T�`� �Vg��}�.�5W��`����`D�؂�L'��N��|��V��lWH1���IP��67y��Z��[TXA�<�afm�ƶд/H�o��%�lJ��w2�<ͦe�o)�}��\����o�?oE'|�<`�
�׷qBy՚ �£��He7��zH-ofiJ��7$�x���kw��=d���O,.��l8��l���Y����unvM�F��#z�x����aݐ1��׽�!��ݻ�!���{��+�;3&eGܷ�`��.���{�?Vl��R�1��k�("�4 �:�V3E��T}�0yW�:��]��S#6��0�Y��Ax�)2�5YԽ���8nl��[J���6�&��®-��$�o)�,�S*vp�QY_.�hvU�3��U��L,N�3Q�B7���P�z6��[zm�L*�n�E�;�Q��+��*�&�X�'&���[�х��NrW;���vw(����e�}���]v�����ʘ-�^+�x�������&SQLC�'٬m�����`_��*�M�1�X<�J�+��<���r]�uf���9:��F^2Q�nP9�-�M��ͳ��{��Uӕ���iʻ'�%��Hһ��BX�G�`�v�\�a��[|�cG2l<!d|��B{���l�g٧��U��>���|,�)��eA�&bV�"-�N���^����}�I�8S&^j$N��H�R�t��Χ�T��n�Jf=����-�F�p��v��sR���ѹ}���uTz��]�H�����sˣ}�&\�66��3���=:ډ0䙃��y*'��l�3&�V��x��i�ƂC��3�Cܒ{�pظ^kx{�j	Ӕ��YS�y���
\�w�I�a�SWwWmt�-q��9���Vi�Mt\,u�<.��ti���J%X�%�;f�3����ـR�CH��ӵL��i�;��B���}P�5�u�o����T�8Ş���M;� �4��,�kӪ�����dӖҍ�:��|{�)�u��z���ⳉ-�C:/^>��K��2�,_)|��ͣ׌\��
�2hネ>��10Ӽ=�+;�&|d��뮩˴m��t"�Mh�:ɨ:�s8n�3�ݚ�L���P�w��֣4�������(U�5�Ⳗ9*{ܣw����3f�!Ϋ6k��c��._[�E
��ؐ32�E7�s���:�!���&e��D� ���f�[�-:mX�2�Cݐ��$50p�k2��n�������p�Q��c6n0MQ��B3	�fL�f�ÊB�{�V�[a��:%�R�Q���
��eئ����q��0e6Y�S�1��*���V`�u�M� �s�=J���ugU���We|E͡��7dd���N�j/{q>�f��G#�6���z߽t!��:���[��!G��'9�h�5�ǻ;%��Ju�*Ro���9��Ov�u=�)����L��}���y�]]p�;���
�>��dC���-���x3�.�i��}}E�lS2�f'F�b�ƨc1�h�r� zY1��8��f����sf!���:��c�=�}-��;��u��\aG5��2������UWj�8��0��{9�S�n��N�:���̎����3vU�s�*g���H�Mya�����e��������vm=�	���x��,w��$�Т�V�Vj�; ��{].�rד�r�ن�dNZ���&Z$u�񮘩i��ţ]_3N�tފ��Ө��ϒ�K2ȧ�uF���y���&u7�Ki�.}�:�_"��f�j�d�\�ΰ�lO�V����Gծ��4U�<��/m���xɪ�����l,��W-����=�V�,\���Aq3}R�z8"�T��-��w�V��2qO�!�LRe�4�]X��R{�f��GAf��1}�i���P�Ó��d�w�V�\�=�#M�Q�Վ��(A�%b�+���U���Vʋw����LY�1-&�zقk̜	�;w6�&;9�� ��x ۴\6[���ͮ+s���ʹw�BⶁbҌ:��9��ns��v�2�Ro���xLW�Vk�԰�y5CU��F���!w#�m���hPͮ,���1^��:�^9k�$�:4��Q�{o9V�fuL�8�Y���?�1��m�֯��gv�%e�2̫*���5&i��ެ��i�k�rf����a���b3��ư����vƃ��M�T�S��O���8F.ԣ�\BV���j�B��i=�l�'v��%&L}E�ڛ�I���z�=]�AyY�Gl��P�aKmEs�
g��Π�{�g{/$�����4<���{���ѕ��Ҫ���ѕe�-���Z�g-r��D&�b�Ҽ�s��yu4��(E��¢�,��۶�u��\�t�r��D����m���)�X�ps���ћч��D�b�nu5t�*$�1?3g�-@a�f�ۿ8�r���	�<0ޞ�}�ᱶ�bI>بIw!y�д�cː��/o�y��|5�p�l�ב�Vݰ�7�7���vI�5-�)g��i�;��B��������Q#�y띚8��K��Dm�ȟat�l�'��9n �Wi��)�����T��-D��]����/k��.]Z��	4���:,f��W6�Y��RN딢�#���GݛG�r�(N����6�upU*��d
�J��V��� �X7�JM�|T���%Z.]�x�<(��+����P둉�ͮW��"=O���qot���%�F�1� ^9n��4
gh���aVz��TZ���]U�ˁq�\4�)��s��©��k��u�r?#V���=�4&��j�;I�0I�&��%����p�������R��չF�dm]n�I�M�D(��xSжMy.�*n"&�*x�n1�L��6�N��Q�O�[��6����s�d�fd�|�aMv��"Z�٦�)���u��&���H�\[��*|k�j���˲j�љ�o����ͨWb�r��uC�oc]
��V�b�t�-��1ӫ2'���&�u����
J��z�3�R:��8�s�WI�ucpf۞�R������r��6���ܗ6/���a�)��w}�f��	D0~�����/�w�+��s���R�F%Q)n-�8��qq�2�p��;dhX���eȲ�r&��ޜ><����F���F>�VI�܊�(�`즆ee�O�;8����VGDޙ����Ξ�	3SK0��� u��~�o�X�ڕ�hu�2*혍f-m�f ݖa�Wtě~ �+�._Oq,��ˎ��������*dY�cvz{	޸0�̫s1+���X^J�����)RAai2J��Z�-�4�i�vYįK(+<��R@�av�C��6e��k%q���7�c<��e��5�s�oɭ=7kkY<��4w�=�֔��P���
�=L�=l67z70Tx�l¸�����w�kLɰR��.��o+�h�c�rԕ����L;�A��坷�@1�(�����@$J���/�gG/y�>ߐ�p�7B��0+WIHJ�Ҫ�ł����N�p�����r*^8�9p�]�=�xb)�g)q5�h���r�X|���r7	�m_��� �mM�/��n�O.�\�:GXw����K��|�� z���{=m�c���A��Ghr���o���De��ڧ��®A�K+>gIJ�n�}�_X����,��(Oz�ZYkN���3���D�9�R�q�n��>|��ۑI�{=HZ��-����T��>���h�`�!��97�Ef���4���O3�J�K6�\#�F�>�FI��Miޮ�	��V�Էt��'�e�5�hX�
�����Z��l���^į�^���� ��}�R9K���\Dd9ܝ�w���c�S�Tvq@S���f�B�J3�ye��dmǷ3/���ͬX�<z U_3KUh{�=��ˢ?{E~U�MuG+Y�2&7��B�t�v^g�6�tdsZ�4�8���@"�i��Jk�w��(V�!]�.�*��;�K9��Z$s�y���gC�E�čNR������4A��m���:�,,lL����d�D�=�;S���t��y컥�7cp���keo^ͦ�*�����sGA��6���M9%3t垚w���\ݹ��hd%�ɢ/�V��fi��e�j��J�87��XF�sR�-����h���T��ع�4h���cK��V��m�M|��ʎ&�S9:(��S �N��!��d�U��:��[�9b}A�C�0�d7c�	l�pjV'�Xgx뮗�խ��h��v��p.���7�[}b���?��X�⃷��7��+Qд�l82PO���)�%����r��쎻�d�Z�{��em��6r!%|㗲��J�|	֮đ��H�ӯ�)���kAW˥�}��c�	�x����
�Y$�Y��鮨��b��=��}��sN�:����=�Y��r�cWu_۰%�[�]�a ��LJ�VuPS�;��q�op�ý��Hw`b�`G�3~te�3��!:g���g%�����a�����HY���yy��#�t���QAKӵ�� P�����+�tnk$�WWe�r�+��o��I�k�o��nE`�I����h"��8��yYy-���R�"M�����[.cz�>���<٬v�v��*J]����mh��"��y�L����Ց�k�+������:��Sjv�8�����"��h-{|�а�N��ƈ�U�&Kٚ���]mC�����m�]�nQ��F�_N��<��f�
�bzwB4��ӂ��{���(����إ���4L� �p����D���� ,���1��8�y�aX�Q����T{OK�A=Y��B]�w��l�y�.��1��p�m�x���@�X�+Ȭ۝|b��}�+��e�Ñ�(��$P�'<�m���G"͜k�:�5�\�;lum���kn��ز\����P;���F�<���9uۨ�Dץ#מi�(��Dc��/� V�,'���e��jE==��j~�����;ϝ�����e��h6
ζ�tu@2�-�[���VF���ќڟ�s��M�7pb�M��R�U�7_ �"���8���n�����"�9�ir�'8bO����M�dUj��W-扇�c��U⬳�܈�(V[�Cq���ܷ���s��
�xr�+KE<���R�7�$v���KUv�%�\���7]`�~�;����j�FE�@��I-t���+��؃:�/z�%��������v���)8�9�w(N�#�|���+��g�`�P�:B��?3�p���v#[Fv�5ۊ^ç+��2�>��g�Z��2������G�Mb_k�s����P!�7	�nN�r�ku�sE,Q�A�l�<�Ҏ9���ܗ�Y:-3�V(ۯ�S~E�y�I)Ѡ�U�{��R�a���K��Ѷ�T���R��B�ju��d֚����+�����{w��Y9�K(@Y��Eպ�g0FZ�1MHݫ��ӛIto�X�.6Uزư3�{]e��N/Op}�(-���	����Du���JӨ��K�=��=�WY���8������r��
:ڗ���`=w�@�;1�%Nb�u��gy��E֊zl�L��v�E��fӺ�K�	��A=�s{�߻z>��ܮ;44�@��C��%��P�o�]�JpS���%�>s)]c���c�L���j��*��O.Yq*R+�b��ڞIM!�g>��^o����n��Ms�a���� #�yҗH�ؐm%��=�z"=����D�s�5�﮻ݟr�s�t}����ߙrD֠v^���᫟m���%:�_;��KN�ܮ)�&����l�sl|^[�����_h���zr&9��-�R�����{�7d'�,a�8��r7�ۉ�J��Q�ov$��KQ��}�nBvѷ9������U�F���5Ϸ��Хfr�pe��d^\�� �g>����.�>iw�Ed�eĽ��R��0cd��!��2GE�������D\�;L,tX2�'f��|;���J�`�;�ǾsIvܱȺ�-�wG�E�M��t×odnq�fi���0⺬�iv�w{W�ѱZ;>��h]�CNg�v��z3i��L��Mۥz���N��f-
�GFA�� J.:�� ��6������`7�x{�=�C�75A�혖`�vT}e|�L��!&p>xc,Wm^	7ݕ�GQ)3��er���{WE�ږ4�1�#J�]�n�7 4
�8d]�ͷ/�3T�1�R��e�x3�=|�oeΒ�UW���i�v!���j��X�[;A��;�/��x��^qv;����G���ԇ�ܩ6��o-MO䩂Ʋ��5+���*�^�zP�:�g�f8��6{j�BGRZ�G�\ZvL�F��<Yt.�p�VZ]��pL�h�6G�ֽo�l���:��W��%�s��8��Ǒ���;�-4���!��]v�ib����&���-f�|�H7�tM�o3e�P�l�Ϋ����Y<s)�'ԝ�	�;Y%����7����Y-�%�@�<�1{���지������ہ	b��/K��3g	�!��xdA��+��s�;}�
n�l�V%������UH���}��k%�&�t��N��L��ĻV�=�]�i�az��4{���L{����\g_\:�Ӵ�����d��-��x{Xz$�f�\*��Z���&e��y5���)��*W^7�Y<z�]���u������� ����uѾ�NۙV�u;��Blٔ���a� rcz]2DB�H�	�z���9�Y.�S)���e���B��k�M�s%����LU����Rz���_9 �-b�K�I�b@�sv���k6�Ez0�Z�T�iҀh����`���j����z��Ͼ���5q#+dv��2�5�汣D0j&zFz���Y71s������xh���E}��0���s��<�;\(��Vq��4/R�b��N�n��l���h�p���x���'�\�͏\�%�I��[��U]<�p����g���V(��R���:�B�/�6���L�0w?�QQ�� ���j��� �VmJ�ݢ2�>��8c{+�,�gu/)m&i�i���ˠ�e�Fz������x��܀��QV3\.�{�$iT��E�xcEL0�/s]}
�땞���[��
�D�s���p�ky�+��WZ�l����r�����ZuMT����֊�dr,q�\U����n͜�K���I�q�G�@2S1�g
u^̊���ֻ\��r�<��a�{p\;�s�g�nXwL�)yΫ���b�r.KG�I4��7���,S�fk�vb�}Q���<|���NB)�=���"�*F��Q����Ι��Z�����wm�̀�#R]���"َQ�5�Ù5ʀ�%N����U��z^��i�F�:S���Y}�H��0ď� 8�̌�eb�����uw
�T�;˥�V����G
���w�g�̋[�/�q��Z���;�v��U)6"�]ov0��d���>J�-�4������/h`�Һ������:��	�����{5Y������y�Yn�E�2F�C%��TR�E]�w��xC�]�W���Q��k�W2��^���v���lg#� ֫�����\va<�ӻi�\�����[G��]�y�%�r����ۚ�wH �x�=F;��Otcڻ|��c��.��r��j��6)�bjt�n�f�OB�hŇ yEG���_Q�)��ԉb��j��+H��HU��7���Q��mՃ�a^���=����>K��]hйe�>.���}3M�Ѿ�jH���� �l@|��<엒'`SgXa2������׊�V�i�I��{R��m�����c��2�w^��4>���TvS��o���[�5`�Ω7Э���>۝��gA�ޚ�>v�&e�Q\�஭����Jdv,��E�f�n��k$s��esЁ���d������w�wsmc��)��9����?�1V�t�$sCS	�7��R���P����6����􂁨�gnJnt2
em?��*�����qA*ܩ���X��!��A�;[�XT�3�b��3)�8�ގ�2q����J_<��Act�a�[O$��m>���ry�.��Fo���i͈����zqn�E�$x��Ua4�&�d�v�'lM ��K��is�0�XT���ء�,�wA���k�xx��C�Ö���5^y'�txk�J��sj�*v���Nl������X^
�s�錇bR����C�V��YBoXWtW�*�6�"��w�A0M�����P�8*�ap��f�R����]�@c�*mJ�չ��w1�������J��N��}unڰ�[ս͑��!3I�����
l����ڳA�v�� z�;p�DS�T՛͹�6L�e&:�Y���zK�"=��%*1�R��DY�[�]b�Lɡ��h��
�2ڷcυ#�9�#�'e|���V�=��r�>5ʬ�2ɕӖ���(�
�P|��`�����LC*Z��e'��|�ڎV���,}�S
nMrsk�G�S��&K����Y��w1^�{��#K��$�3fnܓdN���{�I�����vr&�캗hᙣp�4�dЕ��7�x�.�/M5����C��w�D����;{w8u��� �K�/\4�G1n�����wQ�,q��݉�\��.����hl�ԯ�����Jp�=��\(�5X��{�Q[������v<��L<�ˠD<�uދY�ح�Qq��ւ"`�)��pX�W'g8�O��틋�b��v]J�Q]Tdc�k��=��	��@����8_»s���sh��p�,V�9��J�(���ӏN[7����j�㚹[������ó�2�;\�HLv�1	�R��c�p�>Rop!8i�q�dL�zΝ��n�и��\1�*��;�Պn^�1���b��Ck0��x��w9�3��khŞ��
���V9֐#F�2V.�[�����6��Gp\}A�c+��I�/���r�nl���$%6���F����|s�
g���+:^㦨G}�6���pՙK;�_���̤θ;rX��m4n��1�����EX��,b(nh��då���wJ��44��8N�O0l;k���ص��܉Kh�[�R�@���Z�7ֲ�S�϶���nD��K۪>�q��奧&��ï�^O�VopQ�y-��^iy���Oc9+qvk��#��Q[9��h�BĻ�s��y�>*!��^�<$�_]=J����y[w$���/�@xO���"#o5G����f�<kq�1�x�n�	yt���yQгBW"����7�{t���)ޢ�R�=j^�1�؂�4�w�x�L�b�+;�@���de�"�	�����_IJB���֍-�ɩ��Ϡ�L��$2X�!�:����[�4]��B��XZi&3BT�=�<��;3D�Z��P2D:�՝�
e��T9:a���z�#�sO�����V)�|�Wc�Q��|�nY<UXL�&�O�<��9T�g�/��r	��4����YAh�N�{N���\���6y͌dƷ(]>��/jJ:�����n��!��2=���s�:.+��ד�jc���VY��Y���Q}�:�C.S��.+�2��)S)�����*c6�V����,^b:׆,�J(��d]z�9���I�.��]���1v�+�ˬ��7xa�m5����D�Q���j+�L;�r��³�K<uVF[��\
�ՓɅ��N(Wٷ�PR˺��Lǀ�+N�6�6�No�Qȹ��.�Z'�xvJ�͸yM��fZ]���7@���k[�'\����ӡ�>�bnS�ý3u����%�r;�;�'�n��`Ի���V�����ur�p4�x:�Ȑ�=a�Ќ����/�!��l�ޱ��Y�T���g1t�ͽ�Zh�4:^h����29�<��/I�\ɴd�v�����g�C)��ǩ:5CO��5��`�o��3���U'�b�RZ��r�ܨ9�!n]|֌�^,t,��w*-���]jnj�(��ۑ�eV��&n�`鏌Ȫ�|ꦭ��(�`Y��)�$ټ�$\m���*`_c�F3u��:ne��#��\Q+2B�j�خ��� �B�.ۘ-ὁ�7+�˅�M��;v�l�糫K�cz=I�^��:�{�Լ��&��U�����P��̳đ�Ga䎫yKkR�f��@\��Gňâ����V_�r��D'���â�[����B�Y���a�{y��dҶ�i� _R��F�{0C0:sn�#*�2�Xm�?����7�bP�:0/g^s*<�ֆ-��^+[:T��+z����Zع�-��R����#g6�!ZNC��X���+e�g�Ġ+��H)���#�Y�l����|�u�v�+����dF���陾�C�45�?gFGϣi�}�Ң�*�'��ɘ质U���C�]p����"zB��\���K�t3�9s;I�j쬔�����c�O;l��m�s��)��:�^�n�_:3��D�ȅ��O�e�6�eed��8�,��N�W9C^DζݍNv��RY;�t�Υ2/G}=������N�E��3�%�{C7��)�
t������ۅ⚨`_'�7i�r��u����u��H|�;��Բ��zK��f�Bő�4UV((<x��]v\�T�����C�=��8�n�����5�AXo\ڸa+�Sov��R��T)鷶�{���]i���y�{�a[#������jEM"v����o\�(+���7utgY�r��y��Y���<8�:�r�ۃ���Y�r������ّdT9��UXͷH��8H��ِ��g-�%�壽�[�;����|���o�!���ĕ�-���"��#$���۔�`=/E��#5�Fu�t��ԃYȞ�,X�c���Qع3�o�f鎵��yL����Y�w$�WlS��+Fu0*�5�ꦢ�F��2f.�\^^��W	@u�z鬏%86�77`O��O{�Yy���ϒ�M.����pcH:�e5p:�j&��\J`5��W�"�郲���go]��+��Ԙ��r{Q'Zݎ'�7n�ˇ�hxa�*r�d^ҏ	��p�E7��7q꿬�-�b��wS��Phկ��)�Z���G�.��.噹��A1Nbw3���j�kf�g`�6���~�7���4�Wf3�B-�c���^�)~��ȥ�֧�4���tB����t��~R<�+��l;a�cdX'q�Ҡ&�Tv�n*����3��z�t�茚��vRϡ��\4sv�^��զq�պn_4��&;ۦ���z,I\���O�X�mR}��w�{p�j �y;�˝˔���erdk���~M]6�-Ȭ�M����n�A��B�&��ǐ���!QK;Z+��SM;�֜+���rw���3)�D�8��
��M�H���X��Y�
���ۉ���^�ᛕ�ǵJxH��!�&gbi(i�����W}C�akQ��gN��8�]�-�;��,!5��=hak[���SD<�̫��v������z�vGux��3+��Mh[�N����r��0sK����Vp��ts#l���N�Bô�s�Y;p����W��|��]�sW
CZ��A��=��;�n�!j�-A��ha���r��ڧ��3�'h>�,�)�7�o�`���7��)��V�X]�ၼ�}���&'�r��E"j6]ù���γ�P��4���a蝶gM?�k���6y��<����̜�E�<��3��}�����U�we@��a�1k�R�k![#R���x�rޖn��.��G�[�Ut�I�W��#|{�0sʎQ�Q¶�;[j�S[U��Hv�v�U�G��w�b���#s\�Qu<yխf�fw7ؑ�n��0�Sw�T�i{M`	dv`�ʾ�V�q!��ܣ�P�.-B:c7vms<*��Y�n�vK#�	�C�QJ�R�yg��}�a1�bF�+������Y3�}�z�|����C�,ܪ��ݯHݛl��+#��r�j�&oR�Z]�-ud��"I�-ଘY�������1R�w����f"�����[��uʤ���g����s��F�NxN�2&r�+Uj�!4sP����ҫ�N�6яYɛ�Kt;4>׷G���e�O[��@��t�dkm]K�fө
�V[�u�dsp��%@���}�3(WE�ݠ�ȥBe��TX�̠�k}ٜ鴥�r�Ӵ�uZ�]x6�����F��h[,�zݶw�����/\�sD�f���<��j{E�C�Aď�s\Ι�0�6��n�{*�h�l�\�0⫼>���k����Փp^Դ��HV��j�-�� �B����晋'�z�z�u��xH �ŪJ�v���	�6�EK���;s$��Vaww��]�
Omb�HR\�Eիo`|4�]s6�L�3]
ܲ�_v�մkH�BT��hhj������X���q�������ڇGn��ם��`��v���:�����{	S��+4���7k!�uu�^�P���$k��,�%v������ƥF�u�Q�6ʬ�R��^<S���Y�<�)gZ���V�J��4���9㒈ȝp}��֨`�t)���x���I:U��5mb��9�(-�D�fh�%b/�����cX��1ΰ�z�W���$88zj���/\�Og�z����k���Y�46��}�x�F�U��j\[�,L���ղ����'TcLjcT����8���#}�L��uppH.��.�I�G��1=���9�G��G$�y�_o]{��s}G��SO0��o�>��yz�-�zmRR�=��h������f� ̈*H��(�lvY�>j�W�)�;���e�7j	�N���)���W����Zej�j�hQ7��yB>���΍�䀗o��up�IC��т;=z�pa�,m
`t.��+��:�9I僗�ڏʸ��L����4�KMu-�)m���8E��:�GY�7).��e�꥗,@�X;��..�P�ԥ(�îdn����)�}������F:���kV�vҝ�X):ĝ�V,1#���Il�*��d�3��pǣ��o�r杭�It�ܨJ[���9.�X��<VJ}��C���,*�^����yӎ�`�>��R�e!�PdTZ�
}��>' � �RIVX�f�ae�QUE��ED�Ve��Y�U�e��PQDE��DPUQNe�MUDC��E��NYU��UZ����8FUe�E�AQ��V8A�kY@F9eee�feMYe��k3,#��,���"�
�,�2̪�#''12�
�h�k+��,̌�"�,2�1�k*�� �*�++�����0p�+3(�+,�"H���#̊�)r�r��ch��
l�՚�,�332	�s0*��5jRՈS�E�fY)e�e�`VfeIXff�Y�YJ�dU��T��XkZtFSYaVE�)A�����Y!Va��AI�dU�YU�%��a�49IE-dY�f9dY��Ve��fd�͙���KI�ePd�0e��Z,�&���h� >��"��W�t�Fެ�h�2�)�wd��l���*_?o���d���Yn�hŕ���`�r���¬����g5grvd*W�R:��ˋ2����wf��2���p���X�T���f����{l���핑.1Wp6��5�y_�*sm�|�?x��P��ѱ\;��,��e�t�Me�d�/�Q��/H��rGbV�
w�Fm,V��U�)��=�B���<&��w=��s WX��s��=P��׭�q��<����鍨�Qd1���y���ہf���T��V�G>׵54�Ô�鯃��݌Cbv�ʼ͕��q%�q�ջ3��U�7CU}|�=��@ꯄs���P�̡�������ծ�qC6(�%��ޞu�FG��@��� z;͓�{h<�[5��>���a���nl������{���K������Q��>]�&5m3�t,��R��U���e�r���sw���F#3�]�RZc˼�V�wbb�Ĺ�xƬ=�F	ra皷���c�L�}쮤��Xo귑g�έ2��&kc-0�N����1VG!���e-Z��D{PozV��s��Å�Ss6�9���aw�ۼ	�͏F̭y�N}M��K��S��kڌ��\]U	��h�r��32y�ϳj�/�m�FM�j�2'un;���B�r=0�V��˝iiV䩷���kH��)���F��,��;zk��:���33 �.dO*���r�cL��0�F���q�{���ƈt�c�
�}ȗ+w��q�Ľ��=��8��˫�f�m2)1\w]=��z�f�R��9�I5�Ǥo�'%�፝��(�D�[�5urK`�.�:�7W.����tvu���NVy�E�<����e�A�*SW�S�6蹫�)D{-i\=�P�8Y���2M�/�cX�.\���y/D,*���Uӹ,�fÎ� ���f�<�oUm3����t�oJ�<�f��S���u��P�>�$�Y��׈��Hf�ug^r��Te�*���uZ��2�1ַ�4/���Bw:�xw�)c��F,��^YmY,�zs0R���=ö��̝q΁�:�䷗FT�35h���&��jHyє=�����鑞��P����K3�+��*�E�o�8��o�S�*T��)]Z4soy_G!�1��W�:ٿ��\�z�K�I#��cIqM�o���H�v��*g���n��fu7��`ee.��j%�keq����h;5�c��Mκ��2E�N׼�]�'�}r�Z����(C��w�;H@A�gzi�z�7}���_��ՠ�G�y?8H/6�V1'�ĥ6L�/l>�u��ݭ��[�7�;gl��(���a��g���<A���w�3ȕ��%�Q!��u�ό�V����Wk��M�P1�cȜ��c(<�	KY�(M��^�xC9X��@Kx�ص��ljk��|qv�[`,ED�ќ}-��x���cĶʄ1�J��dAi'(�%���;�T����{��z�,��4-Ͷm�<�>=v�\tf:j��q'���3ȑ��[M/y���w��r��v�}�Y���eN%�w��m�&�R���6U5�LK�l������q�융��=\IO��jk
ѡ6�Ӝ�ǁ;<�Q��]���v/!D�Ɔ㼀��.�I��:�:�.�8Isex�`M��}3Ԛ�V؋�[ד:�����Ȫ4�+׮�%$q�L`�8�/�%�b���,w�h9�m�C�'U�;òxC�j�<�ǽ�1����y.߱�X�eky�X��#��T�ϛ.��a���N�Q"�t��ws���sziN�'�ht��,&&r8F�\JA"j^�1�q�29m��՛��\z����r6��Hk�yݶ2�
�'�;feM�o9���7�Q��Y�c��β�iۉ��Ȏ�͇+�>1;B�&T��[�h�.r���Χ
�З9T͠��ή�z8�	�g�ȣ�z�8��V�zk��ەֳ�]wV���s���S��tUWG�Ӯ:*��'�Yu�<�l�鍏U}���Q|:|��D����LqƮS�S3����)ɋ�ҕg�S�S.�q��q����G�e�J]<��lypi�)nQ����9r |���zt�F�+U�B���c+E�W�⪺�.�ʣ���6�J��ȫ�AP2�W��Ģ�@ɒ�g�R��d\-�Ξc��yBZ�DL��f̧�c��c���HK��!'�Qh�VwV�W�.���i�ZK�f'����${H�ŏ¢�d�T���,3�����y;�&NԲ�.fM.�©3�;+7P��x�y�R{ʅ��͂�LL���>=@/����H;:�0g��!��÷45C��2''4�R�Դ�-L�y(:Y�JQ-�(���R��*95E�P� Whܻԯ5Z!�>h�Icr*�����ju}-�*-���Gm��7 �|c��b�\��;n�)�����dt�k5�@V�*F�d���U`��4G����:R�S�ٕ�*��#0CBJ́�/4Do}�����wՐ�ƫfc;֌��r�!��f������}�����s���Jt;۩1���{��2� ��%�i��/lB؇��od��7f�%����/Y�DQ�q�p%&��m>|��sk�
s��W.�`���P�4�t@�6[�f���ڞ�=+�����ۨ��������~၄­�V2��oL<����wɞ}�bΎC�jbhgYͫm�u=���/�kI5��5�x�7�X��S�\O����R�/�пAN-�e�q��SE�����pi:ɷ��#�9�%��60P�:�W������ p�߳��N���wϔ���b7F��/�gJÜ%�i^48ؙC��S����Ct��/�?o�_E-��Go�UQ���p���4~�c��uMU�=p���f`)�s�ͽ�/��Lw|�s����`3
~�-��HGX�b�����;�H�J��<"cN14�� .:b`.w}�.�,j֭�W��&E���S��7�sh�\tѫi\ni����nt�Le�W�a�b�7ݷ7�j}��;.:P��$lkښ�ұ�cC�����6�g�Z�K����w�^y��򧥔q�0������=�����s�:�-�P^3|��1�+�o���kͅ���bw���y����]���ޮ��V�t�ۥ�ư�����y�¥�X�����ֲ�Y���`��H�m,�tݛ��Zt������-���ZGX8�4��s-U��]� 5�κ���m9�aC��uM	�ɮi�9�C}�eo.�����{l��P�D���I��3�au��:�|r��4lq����i߻�۱a�laie����Gj8l9U�[&4�?v���jV���r~�}�J�@L嚛��͙^Ӌ�����lм�<�+�.��BXQ�D�>���і8;ڬJr��O��U���3��5��ռ��Zf�i���I���9PU��艤��X��s#���%r��u��=Kc#�����#�����d���������� u�K�e1;�]�qR�;N��G"e�)˃��&ԇ�$;'�AU�T+�3w���n��5x͢���DZ�֊S*ߕ�*�̴�^}:��S^���(����a���<�l�;Q1J�42��:1�]��`;���K��{QsQn����3~iQF�9pzX�s�����ٮw��Z��ώb	��ȬO�E�Va�aV|�k�׃�����AstWZ�nZv�msܢ�~�]a�EY���as&�\vFk��}N��mCƾ��aOt�zf�<ut3a��iaΥ��Y��C[X�KY���#�=4�X��V嗚zEJ��pe�s�YEV�E��	�t�p���髩�ͺk�eBkX���t����ik�+��2a�8XS8@��IYM3+���Wnn&�zR`[�.N�����כ�ɊC�@}��]qo�E�7�6��b"����s�i�Gg�곝xr�M���oj2\G�ÜvXOQ;�<�;!٭c*�KtD��f*j�H]�*�(UA��e�l86g_^ڸdQo��@�����Tn��9�(�ӯ��a��p,�?x���ɒ3��6sc�;�IK��������N�l�U�Ǡx��d�;E�������>�꽕j���tC�f��RO��n�}�5�0C� �V�B�L������J���%��D���p�*�q����ȧ��R��p;[At�wo��2�ٌi&R����:�B+�0պt������y���#7�X�Z(�,u�PW�_�9��&plx��*�m*��EQ4�Z�/�.罒
�h�1rd�ֈcC����zˠŎ�o���n�"�Q`^%���7&�m��:�h&}�A֮����݇�ʝ��Gl%5��P���Z]��t#���o1����ξj�Lu��$��,�k
ѩ����$4p��J��5ٌ�R+Vȁ��}��
���QV`5b8�+�\�h��ۼ�?E��Mԥ_jv��^�6��\�[=f��P��9�.��u�
���7�w/Q7u66i0W-=�;p��vw�����B���S�0,<�y��_��O��v=ɨ�dSa���.Y��\�,�u��U`����Q�E�A��>u���d��G��G���C���/%�?>f���:lzz`�ڇ|
��ű��@��y6���f�1�B!ƕԤS̽�UMY{ؒ�\$�I���և�t��،����1|J�r"\ܾ�>y6��n-Z4��r/2��}��]oI�ҫ��*�RXfZ��v0�&k�#X�% ��u[��C|�ޱ����Mh����qTx뙔xu�@׳a����*Ъ�����_y�vz�1G���$��n��d(1�q՝��><��Kp����L_�J1��� d�H9�"s{��g25��}����U��-���O�K�aV�����kzL8�-�sH�|���w}]�l���G"��	TV{Km��P���t˽Y��(��@ɓ
�j���&���]��dL�`�	R<�`(�,�ve>�l-�c��c�G�*�L�ܕϑ�}���c'�t2�1���=<�=�#5�#
�e�G�UNrj���C�x�B�Zɸ��糮��Q<2����L�K�4��m����e�3=۾�I�p�c���o�������
+���[kӚ���o��0�=��QSW�ub�D5�8wyn�X����άD	�fYT��6�ڠ�=!�KV��.���*��0�D��}�op�]�����:kD\q����f�o+����J��G�k����}����&�l�{ݬ��@��fؾ�F�'������q*;g�����b��Y�wӽ�vR��eV��7y=eST�%(	,nEP�L�#9�-�*-� �����71.ji���2�k}T��AV���b�%fU5C5D@V�C��XD�ʬK��q
�����՚���9������g���I�3�����>j��Q:�͖���X��)'�:�仫p���φT���ZQ�xo��`��<oG���x��G_&�)V�+�o!Lb̨.9<I:��!ƬQU�0�>�r}��_Y|ߑ<�Le�h��<���|�����_��Y7WvGo���i���ziq����{-WPY&Q�о��Qg�侉ĭm�v��q�.P\�n�_��zw��N/|W,>�/:�W.��f���Pfi<��[��7���ڽ��o0m-�uu���O6��ז�H�e���84?���s&lyŜ�Ξ��#�đ]j��f�ǜCM\��-"���ۻ�땂�f�L��-Ȧ������� u��������|�f��F��WR���Ͱo�{�NS��np<��@fw{��zR���7e�1^��Nl[�72Ƙ�w���������y�z���F36��N`w�NUkr��6�X��Aҙ���t���Q>J��x)驨����L߰F�8Dw�#c�m��d���D��z�V=��ObF��M^��a�Tt�}�dg(oE�$�&�����MF�,�����3pF�� `�W���T#�`����}@+�?-7��μ���5�SZ;';6�}�f!�W^�7��w��Hꒉ2;͓�{h<�Ul��ވE��݈;3����Mf��C+�cĞ���8�ʯE�ޢcW�L��'L�b�&�����_v��SmW�W�+���J!�y,V���T!�\K }^1��Q䝒A�wYr�˰�������ed~9�[�Yᒴ��^�f���I�P�� �dXqd�y��cQڗR���9gQk�#��L}�0�t�u�\�� �^\oeV���3�âʪ{n�<�٤��op�JW��I�ucyV>�K����㏀��zl�|P7�4k�zt��]5X��VGWT�&]kBJ��}Q� P��{�������=�T��+�q��"���*ʖn�s�8y8�T��zqAw�gbME�g����%u�O�MiRQ��˔��Rf�ٝ)�9Vsvh*ж!$f_vL��Ljev c`�Ӎ��ĥ��X�a��Mh��+z4�Rt*�[w9�I�εSE���`���-hV�d��tj���9B�+"��S6�TX�h͞F?z�OWKw��-�9b�A��qʕ	pf]t��������f�*�ˮ�J��&�tz��N�G�5�gs7�x��F�x��ݙޱ���o~1�EW�o�_��,�^�f]�����+�@�:�f^{�6�b��q|���|�*U0)N��x��)���;��n��9����A�(f�y�yzf�g�&�s��:dk�Q�o>QFtX|s��R���������3�]�:�>=�c$�Ce�!\��A[��L�؃�)v�uV�ؖ���v=���Uk�.v�*9ԯ�L>D#�^�<	���:c��m/��W6��T���9K�x8��e�;������MPZ뾮#znp��.���R�"�ҙ�j-8]�V������!-3H�;@fK|])�`uNז��Gu���3��-.���t�wג���t5�<�Lfnڛ۽j�uNۙ)<���ə����+ �+6��a�#J�v9^��ۧ_<m���W��L/<mT��uE��O�/�`u�oC���Z0�r��m(-Y�:�N�&�Q&�~��Ż<�hg��L�it"[v�h��C�q[Xjw�]���hIS���2����Ԇ�J.� R�hs2v�Z6v��M�g{u�qvγ��]h!���T�Y��sᆴi'�A}q���ʮ����5�o�^�g{%f��0S[`�TΏ�
yP2���	^���`׌u�S�Xj�.t���O7{�!����w$����A˹�e�΢4��7�Z�t���T��8WqW�b��י�<.x����_X$L���ӵB�6���	ٻ��]�������|��*.�kl���,���C4ڝ��X��9,R��	�),����\��&�����$c#�K	\��6mb/z��Z{��;��̿`7��?3w�����.�#�t5VQtq��i�ze�*���¸.f-d֪;mh������pT��p �ײ���&�"�&&��Ʈ��q7�7�����b=��xmLx�J�a���H^*ܜi;��q_jwN�Ev)���m)��ksq��*��.m7W7u����b�XT*8��g��m�5�2��l�&�72���t  �=G{=\�Sΐ��{ؔQQ�ܺ	 !�j
�%j�N�mN�W�\��j4-[��zt�g=��7���vwt���tA�5�'�`p</h�\_y�u�"WG���K����:�������.te���ʉȲ�ķ�.+�z3{��d��\��"ܢٕf����YdXaA�8XFD��ddN�j-CM�Y�XUY�љ�j��F6Xfc�fEfe�TٙQ�eXE��afEQfdVa�M9Sfa1Y�fVEF`ddaY�9-���6M9��k2kDY�f�VVI����ffRe��̰Y��XeEPd�e��4VQ�fX���Pj+
�����0+"�U���	"�+"����c�Y����Cc�FN��5a��ѕQ���k0f
�f9&U�ƴfE�ek2-5fk3VFY�4Ue�Uc�SVde�VYK�����"%�jՙ�a8de��6fe�Y%&jէ"��-h�VK�Y�dM�2rɠ��5�5SDe�f`b啓�Dk���e���c�9�`Y�نLE�U�96�Ye�YR�Ye��Y�c��X�u%��!�� ��7�Ǯ�e��v��W5�v�<��O�z,4k�k�W%�v��9�6����v�#����p�V޵fk2]�Uw=�(�qZLX�hX&q}�ς�S8���9V�i��@E�u�-���7<^zZu���g���mW�%������_Qs�c%�[�k�+1?IY���Ԛ��W�H\�Er=�~��	�κ���/����u�\G���B��_�;�z!`�Ug��}�c;.�;�K;�j��r�0n�+�D���ĻްH�<����S�3\����i���L�Nr�a���W�"Jb�"��O������L���v��5�)6!�s�%���&ru�ׂ�;Wf�P�1oce(���hp7���)?E�U?<.��Cъ>vF�-�U�a˕vRƞ�9�L\3�jr#`x�X�Aꎇ@,ΰ��[]��i0�%�W'`�b�M�K;�	ʗ�n�oDr�e`�MY��� }��faW��L�a���6�����U_[�*��8)��+2��xN�E�-U��g���x&C�pf[iFFi�KV�rB��r���At��~4���Ɵ%-oVК�D �Uݽ����
�㩃X󴜒.�1vg����,t�fI�W��vb�6����od�S�q�F�.2�|�V�z��u��+�܂�齙V�x���|��Ӡ����z)[ȼ	�k����<%��,�s/�T�� �u�F�.��oz���<fI�%I~����a�
���ۣ8�}V��u�<����B8|%Q�77�4RN�߇�r^o-�A�/GQ`"���8;��	H�Yt��*�K�Fw�ʳ$�ƱӚs���pp�
�>J�J�}C.&ڬ��|�İ��S_��p��:c�]��Πص����kF3�#�U�L���S�ɡ5�h�;����S��o'��Q��fnX�+��K2�|�v��>��Θ�L���(���.��L��Q�k��~�e��>���`�rfۻ�I�۽�a��[�hi箲�=��9
~��1~@�V:���"q��@�ң����˫b�q	u	9~B��\+��Ⴃĺ�8Kc����5.�za�4�%N}���:,�3yw�o<F���˿W)׷]e����+�I����>����G�1�)�g����/��R����Wg�b�On7��o���uy�D�t5ծ������/f9��3.-������3ɕ5�i�g��o����Pb�Y*��+�,�&�Y�ט��[w��+ɨ�z�C7g=��-����WVP��^�O�\�N�u�]nSp�u�Y%��l'M�e\��|�\��}�`po]�������v�wý}m���Vh<Gr�w�lڦ*$��4��K;^��t�ݧ��U�|�!\���V�ޥ�{o046�IU��-�~��B}J^y�Z�s���.@�R�v�-���78V��Zw3w�7�s�s�4�c�j��Ϻ���$x}�k�P��}�.�{9�J+�o��mˮ�4��&��˪6g)��钁|'dy`��C;�n]�69;��y�eL���͒36�V��V֥��ؠ�ǣ �~tORFj&�<�B�f1G�B��M@�Z�+\'��ش�j���f���W�0=u��ا��v��X<�M�*$�z."�y�]L���k�,(����}���z�
>+�3�tQ���B�e���HH�7*�5pn	��T�mB�^���x䞼�&9�wT�������"�lD��3��g�mQQo�N���Ze��0���v��E��t���ER�Y���
�u��/�=C����8�+�]p�d��#�ɐq���ڗbdK�)��B�bR�;�ܪ����P~B�@��.'���ZyA���z�G�ǚ�������.%���p7�U}����/b|��y�2�L<��ᑟG���v���M��2k�Ĥf�ES�S��=w�H�2��\[�}����x��9�8Y����%c]��mbz�v�^&.�S�p�,^[������	.R����o��g-��빗���n�p\� �ww����v[C����c�g��)'��ٜ������J[�ڭ$��$��� ��]��R��eq,y�Pпd�{��YVDǛ9��l�P~d�te��|�&����sR~ՠ�S�h��Xxc2����&��uc�X���~�J��#�_�.\�	��:K�3���O؜\
��7�����T5�]�ܨ�&�77Z�F
��W�W
��Q5���~E�b�]y�pu�ĝSUl���Ś���ލ�UY���f�b�'��ѱ\"�w((�_Mw�$`�i�K�t�վ����ӝ\;f�s����PE *!�Nf�x�ZCJZ�M��c�t��υ���1�y.��B�rnK<�������Q�Ĥ����~���g���7�r�:i�y�s����3�ܤo�����Y��R�H1W��ǝ��s�յ5xP^3gP^��m��:.�����(O��U�^�w��W�;�p���:�Q&G�ܵ�a�mѽY{��ȍi㵕OW-�7����(��,�JZ^tX�p��ŋ�DƬ4���;ѷ�6�b�#^1�u���8�4}w�ͻ�/z���u�T����{Wpr���9�"�6p�������yA���Y�y/r��Ψ��
qb�N�8<�;�fIn]�e^s��9o��^՛.O��Ҝ�Хb^`���w��yU��{���m���%'���oz�.]X[o'�t���'$̰����h�Os�F0*�=Q��4�d�xWod��Z�j��HG<59��%a�V�{앦j֙͌��D�#�#��Vp����ˠ`?Gb��&z�G)td{l����a���}�-��_bvx�ʬ,�ۑS�֙�z�LطąkIS{�	���ñ:��_6T�*�p؆d�ML*�jVa�-��!Zf_0rd}�� �{��FNH��uJ'D闁{����pj�1׈�X<j]uɩ��U{[2_֖@������X��+�p��s�j.V3��u��J���]���N�z,���vu��ōg%5���P��A1������ȼ9Y�lM����s�E�>Y��O�K��D�`�JӞ��\��R��>�d���ı{�@�����=
����M��m�W�]��mmd��T�6r S�-o��c������W�2X�d1kyB����P&�E�>Yj��mv����ˈ�.SȄ��7�{�)D��[C�սC%'���Dp�'3Ƕ0����oxcι��<ٵ	E0+���uR���;��y��Щ׼t��]�q�+@�jw`�C�0���`^N<{3`0���u��S\��ͷ��*2��X�IM��kB�o��@ɋ�N�4Y�{�*&!׸7���_m�,�B�ܣ��Z�:��zSvR��px��B�ˣ�Q�{����yY(c�l&3F�W��t7��.j*�ن��x{�t�f������%,zQ$��ʗu��ӇO�6�$�O(�j�\2zb Nն`��{�uxT���钔���v&CH���v\��z�<K�*gv}ʉR�O"���׾D�d��
�yR�#gk�j�|i��7f�}�wz��P�|)j�ԑ�œ���F�^=�b��R��Ρ��3[%��[�ٝD=��S0쳄L�T2�]dAx>�Ƨ˓'޺D1��^؄F�e�b�\�~!NŢ6oؔo.�;�V�q̠{�%��Fiz���VF�**q,3���bR��V;¸��*b�ˎ��o{�:�S��	C����ɏ�$��d�AR>�Ճ7ݪǻ,sS�Ɲ����|�~~�Փ.*��v˫qס#�_�}C����u�8Ibl��mx��޺jU��c.w���\0/A���a�&� �9�õ
�Z"��X�.(X�%q�L��S],'Ԫ���g�Ά6�.�����I"T�N�x�4��M�ׁ<Ѵ6�\�Rg�9�R2�%٦��WO���Г��We\J����ò����ۅ�Ї��s}���\�1[�&��}�7zg-9Ó��Ꙫ^��i����%��\˽�/��+	{��W>��K�z<M�,'�/ ��[/��cx���b��bj�qu�� �������NT�����r��e"��7��>o��@{�? ��x��0gk���*��Pz�򞀆��9R���)x��k��L(���f��U�w��D�Ga���x�f����9./]L�2�qr����Eқ�i����9ISs��5w�*g�԰o�f>İU �B�6*B����2�7|ШO�KȆj��Wː�-͋�x��{�e�d��܂��M���gi�X��$xsT"��S�w�N�U�z���f�n.�ٓ�`iA�Nɕ2cA|&�g���g�5G�s��dN񤫲y�5 ��i��6�g�n����]0>7�hG,Eq{��z�Fj&�<�E���[�/���X���a-[��t�=�7k�di���6��;�X��R{�T+S��/�b��m�v��<�^{e���v"N>=�-~+�g:(�^n��u,�<jBG7*����B�Qz�l��᫺=��\��g_M���b�칖���S�l�˳�ҋN�˫@�"��m�ř��5g�cuX�|�n�'Z�q'�^eN:��s8�΅w�bgD���ǽH����8���ň��j�ԛl�K��b��uqa������{g6���YS�_�����|GD�\I܉�
*��>A����Z�'zji,I���qT��%6�x7��][ɏ�b�%fU5C�D�j&��:%k�3����{Y�Ԗ���.���k�3m���Z���xGT�ӵ�| X����o��D�ft�y�=ٍ5�P�n4�>;^P{Mb�'����2�Ui����"5c����Z�6�w�[=E�,�w0�eAMV�i�P�4�d�>}�z3���JgU��Y}X�J���Z%x�)xK�~d��'u/�C�Y/V��˜�W��p�'�y��쮫�iwn�R�_]�U�N��*e��#��.J0n�9��ngKӹ.�S���X}nC�`�O���2{{,������(v�X)���Q5��7�l[��;��m�O�v�
�m�M� 9*�Iv��#(3���%tlW	J!ܥ
#UM��=�$`�m��K�(��p&(��3��K���ͥ���*�*{���Ɨ�Ѵ5�ᡇ��t��?{�8	�~���2�%d�w����u���mXw��ޡ@�hd�hwSڄ�JՖm����Pɚ�s�t��n��׫.��m�hNEOx�/���i@�&d�(�t.0�5u�r�����.�S᜹=S��R\�˷��u���z.�
\��]vvaJ_y��S��G��{���ACSؑ�{SSJ�,���3l�-��]�c2��Onux�g.>�<��\,�k)i� `�B�5}�f������PM�j-��D��k0�ݾa\#)?u\��rpiz�9&+��%.��L W?�� ����ۨ\�!r�^>�坅Aq�W�3��ec/䥥���k���*��d�!(�]���;�9�����iu���p�Чͼ�Ut�����2Q
��4\ �{�0�Y�MT�*D�.xwxw�er�Iy�ƣ�x��D�l���Y��2V��Zg60R�O�sa�yS���[��yhT
IY�a`dTAWD{n������T�u�]K|3
��J�>�٧ͧG���<�wK��]���	[��>�l^��?6��YU�"j�̙��F�g{��Onz�o�Vp~ʺ���fg]�џ���4��N5ZIs���9;�(Ry/%�k=N�]��ɓl�4��Z^��{�Oj}���9��÷��hw�f'�$����K��Hݬǎ7)^��hL�-��M�v`AN�y��N�.�_z�|��X��,o��3}˽b����v�ۃG]^�7�Z�w�ӗ��x����S�:S�Εs�����$C�h�z\l�uϑM>it��TcЩqtua��!G,�����=C��Χ�.�������s�ų��4�=A�Eg�q�W�����pys*��LJy��o"�)p�+H�t�D�H�V�2F���]�X4�da���ϋʔ���G��]J�t�8�R�*s9� P�=�UE��]VE��&K�)��o#(���ñ�x���*�c���q�%�#�%<;���6-�c�����[C���Ƨ�b𛸯ޒvNن�ɪ��J��뛗��5�`�A�sҘc��Ѱ<K��z&4Y�ao�ea˘Wy>GJ�vyrZp~�p&2침-U�Ȝ�|��+�N�l��X��R�(�G|��eN��W���NN�߾�h՞���/�K0y��L��4y��2R�<��P��}q�H[�R��288���[5�C��8-Ѿ�,����{V'�T�_���(�~-���oo�n��]{P=a���)#%�*'jӂ�t������α�:/��qYg�ӻsY�����*
�5�@�}�.M)44h�6��ОTh������p-��cW��b����j�U�nWxDB�[�d��5�Ӭg,$���xU:X54��J���WI����j�@���V�����ԦO�<�$_Y�2��=�#[)�G VR�qU�4��k�yy�u
���"��NSW�e�[х�WXw}@��%p�g\�<�r6�S�&Q��_�5��Ca{�9��]�$�I�E`�}���H�ʑ+#��J�#C�#��*d��/��r��ؾز*�Z�a�M�8A=��㍋F��Zw�}��ѐ��׳mQ��}K�:˗)�N���ӏ�,y�\��tv�Ӄ�^�/w�\y0�@7���:坹���	��w]E2<ǒ���G�C��
���g)�R#��S�Gvj ��o儬އu��%/t�]��2�k���in|��+z;#�l��z����C)kմ���rW��@�´EA�3�3h�z?Q�q�FywU�V�����"���;��k��4ExOA�uyr����l���{�O)�4��pI��[�" ���GR��QV/ݫ�gn����G�����`Q��A�ai��:9&��h����ʆe����1�&sQ�w��<�\�T�Z�b�,Ruf���яPH&�ؖ��G���uc��C��Y��}�F2�6���,�Wl9���pY���qt�� �*�X�$�W��N�Nn�5Y3�=��\Dݲ��J9*%l�]�
,��3n.�{�	ぴ0�e"0l�}՗``�Yj���.ty�t��ܤ��`Qس�W5�md���u�{{ŎWfβ_s���I�d���g��u�6n���^ձ�3�"�{}4<��M�o�.�s�
���dl׀�GT��7fEaSJ�J�'4=�+���4�#��vv��&�n�Iѽ�}2�˃�"rV�}��>�6!�m٨�cj;�Ë�o���V�R��n�sM���%]f�M�d���5a���m
�{�3c/ILa����S�����+Z{��_��Jh^0?b��tҫ���+��E��z';�7�W�n�Ţ�$gd���cy��xm����/-�K
C����?�xOa,����r`^|;tˡ9���
��e&��tA�}����&�U�b-l}e�;�heb�9][f:�㖁f�U��n��.��ic+Yj�\��!��}u)�T���NYy�;��u�4�ك���݅��l�Yz���a>㖵�j�#r��BK�����M��.��7������Z/�%DdS/vr:͙}�)��p�kh�w��t5[�9\���Fe�oi\����$}�k 4i�n�<���o>x�Z������v8>�)���%�b�6f!q��K�%�N�k9�];��3u��k��De�HQ��v������^�����c@��غNx�l���=S�j�4��d�/b�J�M�����E��t]�(F nګZ�Z�̋*�J�ŤՖ�Ģ�&r�1*�(3h���*�(����2�3��

��"!��̬��3i��-��1��9j�)�����*L���2+*�2�,�"��2ª��$p�H��Ȭ��Z4k �#&��"�Ʀ��"�5�F�����#kU�Ȳ1���',�+#$�00�"3,+(Ƞ���)� �&�ș��
̈�̜2(Ț��3(�&*��2�
���ֲ�2��dMQU�dDQLTUL�Y���̢&�K�9fbd���c�j1��cQ��ɵdTZ���1V��沖��2\"�Xa��TTa��ֱ������2�eLE&�3�*��"��
��#Zֆ��*�3#2�ʊ�Y�MKjʉh�9Qj�L�j ����PeD�BӖA��&b*j���&
"*�+R�AD�T%,�E����U�ul�>}8�d쾙���m�������G��>_B�!x]�g�B���h�GT���\�;�n=_a�1*����Ε�V.����'�_#uD�p��Ajm/X3��z��S�T(�5��^�P�sg�k$櫈MR�hJ�J��쌘��IO�Y55�bi�a���ъ�ѹ]e���)�����m^��\�g1��v�� �r�P�6���\�/��%͕��մ�ѓj*���Ǻ�0z�yh�:ù8^6"��Z,c�1�:��b��X��8��,�cv��ҽJ���*_�9�n9Ԧ�E�r��R�յ%���	c�a���0*i�	�]ّ�-ss�q*�=&S��~��f�ϤR�r�k�m4�y�4��|T {z�����{�.����n��]&�s�m!2�F��ZU��ȇ���K���#ֳ��l5�5�IO�Z��3Ș�~�ò�T�z��_{���P���N�j�r��13�<� R�&:���̭����I �����ti�j�bM�C�13S��`��C�>�/<­C9��
hA��S�"�7{��e���uW@�}`c���w���jή��rG�5B8\�	���X@[<}o�W,
)h�r��`�"n��@'紹f^�&4��#*�ex�"��&C�e�4Z��y�׷3��6i�x��}�g7j����p�Q������ ��:GH�78;�]�E2G��Rp�j^���M��r�������]�u��������o��z��������pf[�eIc���O��e�-ٕ���J<��I��[���������z�d�O��P�����FA�ɓę��Ǖ���9[k�9�F�HO��^U����%���L-��);�&C�B��fғبUnu�`�SZ�`5���uYv��~ʙr��%�rFܕ.�:(�_IT!�����箊�q*=~����쇽���o����Ad�i46\ł&�����)@�$��CD��5W���S\�U��5��ջ���k�ԋ^�:=c�u�Kf1�������T�}���P"��*F�Ply����^�K�ԕ�<%�"`�� 5;pĞ>6uz-ϼ��Ufj
��@���p�J�����oF��pV���-��Y���n4����c'�(�+������!A� o{�=���O3���L�ޖ,�=3(;�ucn�ݤY��#&�ѱA�zgMeV��N�^�n̺)�D���4���ϝd���ḡ�n��)�؍������=r�\Yr����H�BY�}�u�lQ.�&��������8�7���)U��꼎Y��/!oh:�d�^�z��k6z�+�/u��'�����s�Z<�c�
��<�]1�45F��5���4��gxɒ���Vjw.x o�W�}���n����������J�j:$��$�:�����R�q7y7��Ok����V�4��)�t������`~���S����*����^�؝�E?���������ۡyNɬ�|�&�M�d���`�V��ح��R�~yζ��ea����Y������HP�8���������XnG�*��M�{�H`;O�$O`S�S������y[��v��,��U�(�Rg&6y�1�
b��=KW�{�GB
Sؑ��jj������i���sʔ���F)'���Y�f�}c�9e���͆����0b������ՑΰRZ��}��{e����u�PP^2X�?J{^4��)�Cgk�m���>6IĔI��7:^l��Xy���9'"n��#5��<�V�}9��Xec��������Pj8mʬB�����6'wI��ͽ<�_\��J^����<�,m�b�����7�0м�<�b���7���1Z}�ѱc^Ĭ=�ikhÁ �TNjf�?k����_�ɣ-��;�t7��WW���n}}��L��w\�=�͌
�>�m�=j���)d���2ΚU�d�@̜�[�Ѣh�gS����z�A�S�ul�2��G�-�M���&�g��s�����Wݾ\�����O���F(o��G-]�]u`>��D��K�z"""2�&�J�ֆtH`Q&9p���2�27�]	}� �����+�^R��y��� 9U��.:�X2\c�ü� �	OzxSb��buclq�}�<A�C��n�I+�ͷ���F$���W�W\u)�9,Jg��*d�O-I�5ZI�|zAGj�i�:a#Ϗ�\�9�W��6�����V����V��Qs�d2\���E�,u�X�����}BX���aZֹu��e�]@�����ժ>��B�<��+9^�� �B��oS$5���t�Ɣu-9�Z�F�y^V�����,��Ұ�ؙ�y�/�ްH�=b�ɠ��Y�U����uV�nV��K�*c%â�mw���O��d^�2dƈ�6���˩��ɦ.��.D�����'s�:�X��S��)t��
&���@�8J�s��n�y��[Dh�ת��)чPw�Jb��ڜ�pt�ĩ��곜�`�;�ؒ����4%��=@�Le�R59�������Vf�/�o�͸�p���lP�oNWB8�vU�E��Gc�G�g��m����VY�$����_F�q��N�]GFe��E�CvF�︚lc,��и]=�@ٍ��˾�1oi �����5�(��Nކò�Ը�B�N��f%��a������v����{���-s�|��ff�c�J��v�
D�����Ák�Y��X��{pk�79�J����[���r=�mnn(wȕ���&K�ʉ��F�x��B����i��/ӘA������,_B��g���{q�Q�b0<�\2G�,�5�+t������ئ��Ҏ�i�]�+�ā���$9���*`�8��E�h�����/�W����˭�^�_�n�Ͻ�'�Q(k��MVs�:�/��0ЛK�p�k$!R�����$�رgv,���s��pp�1F�+&�:�愈�Ff:ꄔ��L�#����f��R�\��w.���H�/���p���]��FZ�Lw$g�b��U��t9�O��
�}�Q>qɾe�t=�=W�7�֌�w=vnz����+��Q�c�x��:᮪Gw�fqs�4]�;MY=��SB�/ޏ�o�	�'�a���F�m�.1r�s���ia�'u���}q�FM���ΝCgE?n�˱��ҝ:N6��V��ׁeU��'ow`�]�0�pJ����w@��k�e���f_|	�JK;Z�����N��/#�dz6t�¶a~��V��Lwz�#nHk�;9us�ܧPd�ةMH���݈l}]���c�j'�.�[3��Ь�9�t�\�Ҹ9�\&�;x�t�ع=Hr;���G�ڰ���j�s&~��L�Ʊ�JAg�U���lB�����5�c��Vu�1+��Ε�ޥ4a��-j��x�� �dKwU*k؝L�`o)\#W<�B.�ܴ��X�dr�w+GF��[�ֽ�w��O�F3���B�$*B�\����	�R����*
���U+nݻb�;���z=:RR�W@�}x��1S7����J��4�NhS�����A���ݼ��*x��ȍft/���,+�D¾�3�D㌱���l�7�n�M_r���-i�������)Ecѐd��D���M�*n��a�W[WϷN�Q�]��Rp�O�i��vz]�r��q*�U7R���4�ɫv��m��緕X�.�s���1Bw>����ZS�7yK�=��䟥��
Srr^?o��+�{yκ_#������;u����{��<�9څ�M��㋷�S���=1�#�q쎤���r<�����9�1i���.�P���ܜ�'�w�������R�����ט�y��Oƾ��X�qY��}K��yO���G�ELDd����hN�=�ϵ������5���`{:�Jy;��?�r}�������S�pܴ<�I��'!���U�������%���g�{�4x26�����kX˨�����v��'Ea�Y��Tn�㔶�t(*۾=�)�X�p�y)o�Qork*����N>�ۧi�jR{�hc�}�6���Kn��k7��z=Nn��L�fUeю��;t���B0B����z".�j�v�Y�_�H䇿����+^{��MF�?����	�r�ք���fA�r䟧sܼ�#��#�<���z��w=�#���v}���*����Nl���Чޙ_-I�Pˮ}����9�˸O��K䚍Ht�zЙ:���!䧱��'����_��w'�r|���\�>��1�c�&�i�}�:���O�pw/���a�h|�a�P�[�Α��o�'�쎣���|�Q���`ru����<��ϰ<���LDWɸ�\��e�ߵڏ��A��tq�䴚?a��]��d����5�|�/��4�@rO��=�H���}�{�{'���>�Hwϴ�)�������-�����|���r�� Ϝ�ީ�#��>����X����>� y'��7{#���<��ཟf�7&��X=BrO/]�#��y�N��S�7�������Ʊ.Ͻ�>��{�>d�+�E�MOк��z���'�����_O~`�@rN�a��ZOӸ}����ܛ������	����}`1�rs8��]6���{�ޏ���s�z��O���%��7�}+�M��擫�����Խ��=z��-��ߘ&�>��}�G��nM��u���H�bJ�;�Efqo�]}�>�������w;���Δ�S�9����>��b�!���\��Gy��r����:��`?����w������a����d��RcE}���}}SsxrNF�<�$=�s�v~��O��~y��'r>�
O������ihw�u�w��{nG ��Z�tǟ�_e���\~���}x��}똈�M��s�C�NA���=@~|�����?y�{;�%��iܮ��\���~���h��\����ZZ]ۻ?u�=3
a-�ϧ蟯�"�78&��z��YʣHb���_��Qߋ��y���ř��]XV>�[w��jҼ�wC:w��F�}�}�
;���i&!��]��N[�����}��i�\�Y��+���CQ��a�ٚ�D�O9�����4����i.���:�Y_�UUU}9��/>~������V���wy)�z����d���''�}a��f���^A���	�<�����]I�����Tzg�}�/���	��?�Vq@�����}���ih}��ց�7==�A�qI��=��䧯XR��}'�h'wG��S���䟥���ܜ��߻��%������=�ֻ���߭Z��,���R�����Ͻ�z#��z������h��h�}#�5�O$�~��X�pny'Ϙ�����1�N�:p9'���;���}y���,uǕ�{��}�>��{��U}�tǮ9u��rG#��C�b��P'#q��j�����GRv���Jvw�|�ϒ~<Ó��v~�:��|{N�����"7z�ӽJ�~�>��GЀrO��P�!�i��H�[��.��k���-Hf��$�{���<�fd�ܼ5�����9~��ʓN���v�����Yz<�Ч��{�S�W���ܽ^@�<����=w�rZ��4-�9�:]~�u<����Hsx�d���nkHy�w߮a�#����#S�V��ו�>�l��~��r{�B�'�~�OR;���yy��_�����K���hs|�?F�u?�}��MF�;���}�g0q{}U�4�~�>�	�3��#Ѳ�GkY��>�j�ܹ?�0�A���ewa�wy#��ZC���_��@nOc�ߜ�Й�~�t���?̺G���b���S��-O�jC�}���O��`}?J��;�<�����$�\���M�A�����={�%�x/�@n�!ν��CϦgf2oj���Z����c�S�鏒�H���ߟt�}�����gR�?֏�}����4OҺ��}'��n��'�iyO������}n�9�Nr�����v�\�>��1*��͵����t�|����d�}gv���fX�ݙ{SE�4}�����"_4�x�K�Ξ��[2�S+U�ޝ��ܠ89%����vY�X��Y�T-�؞���-(+x,��M���][��*�&���̅j�����z<z�)Q���}����_ϱd�n�֗�I�~=�:Sp=��}<��O`��zCrd�ֽ��&㙁�䏑���>�˘�eFLzg�lz5������M��k��w������8w���hz��$�rGW��q�w�%=��ٽs�~���t�a�w/;�9&K��k��G~�A�nW�ߞtf�s�{�Z��{�?~�~������&�R���8���ܝ~ގH�/a�ɻr:�?b��但���s��}��;���h�����L{��>�>�*���ǹ�f�tf��|���=����Դs9��rG �7����S�X�������'�tkz>��^�Ǔ�����C�7>K�|�}#�>wϺ^�r=���ֵ����{�}�;�����
O���ޖ������_������Zs�w�)�XP���{��9'�ޏ�<��1�w/z2c<��O�'��͆tG�|O�o}��_~��3�?J�Nk��s����ː�斆��ǿ��4��޴����`{'#�C��?I���ش���f>��l�#ݡơO>�'���5O�nϰs1Od�/F��O�<����C�9�7������'r9����GY�#�I��ZO$��DP��FO��}1��/$�CS��,�c�@�;����ԧO�I�>�y�nNK��֥y/�9�K���x���b��C�C�q��Н�}����>��W�#Nv���X�U��Ϝ���)�7>A����<��0�^�R�y��9.Z���Cp���yѨ^K�Ϻ�uyGa��|���;�ڈ��@�G�
c�L�/��'}5�����{~��Hu<�Z7�y/�b{?A�g]�I�N��u?�w�c�z�Ju��������4����j���~P��[t���z�2��i��G��Z{o
�TA`��_l�GR9m~��t���kOgy��f���l���v}f��v�95������Z&�)oeAp2�}}m��{,���X�[ ����Xi�#�9�hG"ݮ�v%i\۩�SA,U����G�#޼������_���j5!�w���&I��?f�����ٙ?@���by;��<�c�؏$�N�é�Gpv{���y��<��v��xϢ>��1�#k��Y�m>[����2>�}'�䎧߱I�R��L�A�}�i }���d�/���w'�r|��ܜ���:�����������*��G�oku|~و�>����x�9�������Γ��GS����O��N}�ҙ���޴�A�Wc��K��!��I�}>A�1�E��쎋�&~T�m��h�c�w'?a�w{#��P��b��C��}��s�Hw�>�=�e=���z_g�5!�ϴ}#�G�9��~��c��)�\�O�2��跂�%|vZ�����d���O0CI��������1ϳP�q��C�'$�?o��M�v����`}�Ý�|�`�yϘg��ϣ&ws�ĳN�Z�ݿ�^|����9ޓ�|�B~z��.刺0N�9G�>�+C��ɸ䎻�BrMۗz�����k�)�9�{��ϽS�1��}�e�ɺ�_��~�E�d�>ֹ�M���Aչ_c�[�u/�p�����w�O������a���;?a�7���C��ܿ�O�b>�eF/���o������[{���#��T�K��{7�!�2\�vo��i�=�{��?>����J~�@~��b~;�;���Y��G�{}>�0�ލ�^�}v�3l�N���<�}=��<��'$rN���K��#��z)<�'��~ޖ��v��u�w=�AϱZ{}֓�w�)����K��Tn���U�ΰ+�+��!��+�{��!�0�������=���?��;�ԟk�����<��-G >��-.�ݟ��4���5��حs2�_���_�U�A�(��w��4��TVJ��Vt���� hU	�P��z�u>�=o�N�9a�,�%�pߚ���΅g;�	�JɇY\�[���#�^�P�!��^e�m�5��ƿR�/ƞ�k	�]�V���ȕ�Yp��������K�!)���2��9���n���d�Y���ݺVN�[*�c{�ѯM%��7��d�����hTCNd���t�w��qr8��gV곒�1��攳6�N�ל�f۵���ӷ�(寧U(TS�p�@�h�R�::�^�(r����lz����d�G���;թ4�賹��Ӧ���Ҡ�wG�$�Av�vL���D�]��SW�pT^�����f!LfMA�7�P�,J����`�f���ֻ�������g�ukA,�׏7��$�z$ g>��z�����^����,�)�3���y�P�t��fC��mJ�4l����/{3`�U}2�W9N@X�V�5B��#�İ�Y�U >��*�n�޶�IQ��&������n��t/c��RWd�fLC��uF9}��Y�7Q�P�p�|����~�w!�1���Hi�>kz|ޘ�{rX{+u ���&�9���UW����wś�3z^��#�tq��(]�Fl�s_t����ul9<��A��@���M�=�ݭ�!�b��쏡ݾ����z����k�̧v୔�p՗���>�Q�]ϐ�;����铬����>�\�j��'@_b�N�#Y����?wu�B���f�����fH�E�pR��?^gG��@�Ԯ�I�;w��U����v��{� �FOzS3Rjs�
�۳#�n>�#�,!��v�-�w�����N˹I�9�gnM�1�5х�|()�ՂN�4�'2�Rmf9t��L�������u�Q�͇��ymw��9�q���*��']'o,�beJ��NܽȬ����D~9�^=p:�-��>�1�3�����t��pc��vC"5��W������IX��ն2���Sx���,54�ب�R�gNVs�c�k&L�}]#[Z�S��+zhI��;�쐒�4�X����if��AHF=S�����h��X;.hI������Q�gG�#�-]�]�se�YZw��>͏zѸ+��)�����5�y\�.�����#�@cɩ�^�5��imn�݊M���w>��8BoT[ս��k�p�i3�u��Σx�!�)Myj#���N�备�+�p�ߦ'ǮIj���@��-ɳ;n&wY�Z4G��kvx�J�v�[�$@�%S�2�:�v>*�w,U���3Qp%|�����t��ꈈP�)t��ۙ�X�4ã��i}���/7��jG@^E����Iz�Ȑ��I����q��^K�F��;���X�}����L�X858jls��;I^��y����hkk�x���;�3���ujɪ���ATe�AEU$�̢�jgX�A�9��d�f$TDLS�5Qj3VTQD0EDI���	�p�X�5NYd�df4Fc����PRjr�'	*�eD�Ue�T�TT��E�9�ATVa��SFI�dd9Y�٘Ր�Q-T�bMQ�,AD�ECj������K��Q�LRC�d�aACE-NcA�D�FFCAA%T�U��I��h�&2�iՓU1U1DUTU4�M4QMRTAM�!�U%EMAE��Y�1UPSӐd��I��T�-D�UPQE�MYY�Y94��)�-fKED%S$�eAU-41,jʦ����d�TЙ&@S�`U�QMTPC@MQSAf.fSQ��MD�EP�eE4D5T{j�����W���G�w�=��w�L+�V/�u��I��K_w�]���枬xv=��७s�pu�V�nX�Jer�:��}��U_w�;����~�o��P����?��p��GoXnS��1�y>K��3䟥��}���;o�/w%��-.[��9�'p/9����G}����\Ϝ�b]ܱ8�����""2}1��G�"��<�����Jy���y��$�\�`��Srr_�ֵ+�|�*���c������g�i�S���ݽ�x������S}�B>D��s�1g�i�>�ԝ��7Jv�ށ�w ��-#���?K��������#��C�zg�+��>����|���Q�c�F<d��ݼ;�_{�{�+G���q:ޓ��q��ִ'P��3Gҟ��X���]b�N�����+���=��ԧO�nZF�ϼ��_���\�^w�_}�>��2^��Z��}�C�1Z�9�/�j5!��zЙ'/�3�'���k �S�����w?�����O�zy�S�.��Ͻ�2�����{����~uߚ��������䴼�'_`@r]t}�v���9���S�s�/�j5!���?Bd�~����S��ѓ俠�_�X;���>U��F�y����6�F4b�8���_��U���W�8����y�{�%���=��5�uѿ��Н�7Γ��GQ����I�ԇ\�G�9:���bLx�o�EJ��f[�[��u��>�O��G��ryO��y�{-'���W�x����x/g٨K�1;旨I�s�i�>y��'�짲s�>A��C 悇@f�eg�7|4���z��~�kA��W����<����X����}=���Oѻ����<���Y�7�z���yq�9�?��U�yaJ�ټ(�f���盙��b���7�/��u/��k[��O#��u?B���z���'�?KK����	�$�o��w� u}�!�7����� !����+?��給��C�wp��dŃ��6��A��i�!#�0e��r�zu���w��
o*;xZE~�l�ƳN�W2�ڇ+��A8̖{ʻ��LWqd��8t�U��d��s��6�����=f�$�t|jT���0��%BGd���G�5|����������������@�S��}'�z��<���2\���_J��q�9��䯱��5/q�MAܴ;������>������DT%��ǇG�A�Y������?o�w���7#�{�=���y�`~�����S���\�!��iɐ�����;���Om��� Ͻ��𘈹��9'쥂�]b��������؝�w';���=�w���䧑䇰ny.�sI���9�hN�~��)<�'�{?oKKC���δ.ᣠ�ZOm����?}�^��s;����~�]�~�����q5��:���M����!�&��Y���;<�����?`����{o�;�ԝ�����?���I�r��4����^�����~��i�Y��w=Ϣ=3c��v�-=�֓�w{)�:����d���w	������7>K�<��NI�ﾟ�u'n�Η����f����5hb��Z_.��=3�	�>�����|��n?f@}>w���u'5�윏%=�
C����������Jy!�`rO���nb�����oz��~��S�m4���.�_yO��>��������gߺ]����=@d����@}=�G#�I�u֓�7Jk�S�7<���ZS����>C�ԧ��_QUqX�e}7y_A�h���S�	��RKC�{��R�������G�[�����3�@d��Ǯ��:��9���GR{�Og�y)��'s�C��ћ��i�}Y{Z�y�϶}�l��:]N�8}����-C��!�it}��Ԏ@o�iu��9�/��ԇzޞ�2NGљ�j��浓��w��]�?�)��s)r\��1}s�)����<�<������'�p�^@�{�!��jN��rZ���дG=�K�؎��}��MF�9��2NF㣿����
��.���7*K������b��t�%���!�1�vZaռ,�W�)�������՛x5F �W�non��(wk�d����]�k=��p. <�=̵�,�8^r��;1�jWw5��@���Op�ȳS�^drlg����o*�=�z���o�w���z��2%?K�`�'r���=�y' �����߸j^^@�{�!��x���@r]u���Z�o�'�>��;G>��u�Z��{��r����욍Hq��>��5?Ga�hO%=���Y��>�~��~�'���A��G�����5.�$}�!�s�D	��>��P�]و���^9���V��|Gp�>�'��:����|�R��G�9:��ٽh>��z�9�I�ϰ��y'����b���_��수�L}>�1���
����tt剾߳߾�y�~��������G�s�Bw�>����;�K�Υ�s0�G�?O��S���֓�z�	�;���:}��C�zf#�����~v>W�9��V�hy���q_HrM���}i{��G��s�7�<�O �S�<�zCrd���W�75��y#�~7g�S�l��E�򴟍;:�����/�g���4����&�9O�w����rM��u}!�7�����S�7?�g�Sq�'����˞Po��7Ԥ������n�y���VM��-}V���y>N��Z��"�ɍ���7�ٜ�Q����0{4�ŝ�^��X��'^�9m�D�ޱ��Y�&���^�����}ѓ���z�Aa�Thբ)n���վ���Vg�ˬ�p��'�Z�#����y�ߛ���b�׷���1/�O3�5��WN���՜s��t�"�ʱ^�	��NF�S��څ�&��`�&
���Y����}h��} �-RV.��DL�s�Qɐ;�>䯩�+�e-��M1�vPe�W�R�՝�a��N����2��z����� �Jw.z������U^�k��<�U���d�1ʹ�mߥ\J�n���R�j�,bu"���*���I�Q���`Ƭ��L���8��+b�8�V��AO^c����49�s���Z��إ��' ��ï>#"�����T��������Y\M�l��A�PU��_�rcx78{Vx�s��>�&�]���<%B@�w�j�{^���OZ�O�z^z��SdX����3��s^h������ۑ�f���
��13�:�!@cuށ�W�f]�Isgqߐ`�wQ�足E>�P�ig�j�r��h)=G�!�jX��k՝��;����wO;wsܷ�C�ܿK< ���N��saȧ�}Ϸ2z��v�)@�5�	+F��&�<Ou����ۉȼMf��w�i�r�7M��B��p��-&7�T�r����n;*	9z�^�湥�2<�W+��M6���^�ЗY��� �m�˼>�YA�gu�b/[��T�{�#St���]��ӥ#�����
]��yl^�O���[�&ϧM�	�}���^�Q����e�����)c���.{�u�P�r����磌��L,��}3�w�p���Z��M%qC�󪴐���V׫,��Fر�P�-+����T�v;�=M�<�R���1����J��Wǵ� -�׼����VY[ϸ���rv����z���w&Tl���ѫD�ڼuԤwn�����Ʋ�wrX�����j�Mk�ȗV��Y�0��Vg]��u��Z��-|��h�J��V��Տ������;�W�!���j�t+:���[x�ye�<����/��ze<r��ԑwf`������{�q�eAlY^��a�V��
�
��.�*����]���(̘-L��-�MeP��.3o���/� ;P��{^5�.1�� ��(��p���:�:0<Q˄��2)� �W/� :�v�b������g3�H�Yٛ�QY���W(@���N�6*`��؛��=��-'-H���Wgu%Ɔ�١Vp�5aK�9�@�6`sh
8��Ho�΅�zn	�I��FͰYZ'Z�9�c�ǨM,�\�3��e����Sz��*xN_t�h$�gb����N;�3�V�wK�NAǻ�V�vl�����ӫ�2q��v3�KQ�Į���G���Z���ֺxM^���5ŽA��O0kXݑ�9���U�����U��	�*99�=�q��dV�uz�8j�v�_���yۺ;i�"_-��yΝ�ﻥ��&?�V����b�kg^��	;F����X	]��JN�|�u-8�c[��4'+/X<ju+&�Cʌ����Ǐ��5����Y%g6�U��i�W��m=;�v�T�,�^ڣhT%���b�3�v�� ��r/:V��K�E����+�Tc�����KP���׷<�{^V��8��7廒7�U�ifjj"��;댞��䩞����i�jm�͉x��߸O3��'�q����3VU���=��d���[ML��r�}X�u{��a�Q�V��n�ｵ�e�^J���A�NTW*��BbFV�Z�b[[�Q8㗛��}Ah�3�nZ��c�s�\j9��pO�GeܧW�w�>��6���E�j[�c�6=9P[� ��k{�/��R����t��\>�p~��_]Q*�-����ز�rq�/;^l���rî>�{���uf�-��C'.�=fB�c{�oD�V�׷�;����������JgFQ������U�����q��A8��jӼ�Zf��Ďm�2�:1��W��q���J�G�o��:��I����?/s��v��p[�!=�N�>~l��X>��M�k�1^
����0woO��y绒��~j�����<�{T0�M�p^�a��WZv^��a2�Bx=��^�mW�Gm��k7��y^���0�����N��3�ce->��R97�{��ʍ؛U�=���f�<mm.�|�`�<����ն�,x�Y��*�?�W��~���f��h}�)N�f�(/'�[6�9�ْTd��tw9c1�Oy�y�wf���Y�J���|'b�Sp^!�R���nPb7���ITB4���O��Jd��V�z%e`&�&n�(��{���S7�`�|��HTsJ��V��|��v�ea�r<=��Ǘ!�TU;�_]��$�f2S�}n|)��'���v*�Oc�k�tt57[R����Z��O�C6�e	��T�X��b�n���g+k��t���zŮ�O��]��A�y���Z��j���[�� 9�Q3�	�����L�7��ꯪ��)�����I�6��G�i]1iդ�E�t�'xEڻ���%�д5/.��Գ��&[ۊz4j�5�b����ck.3VG!g9ޔ��u"���x����ԯ�s�귡�����ؾ��0�|�ۛ��L������@�Qi��\��*�AoT�'��s�*��)v
�&_�_g1QP�'@ܾ;vonw!�)l7��]��[-Gpu�%<F�1e��#Ez7J���Q�Ќ^�3Ɨ����.�y��l+b�I��7�W$U<:����K�TX+��+0����<��2;�VO`n7f��i�t�����+�F��p5�xҺ�6���:��S�y��E5��"/<s�ݯT\k�J��Čچ'��+{���
�:���h���&�����Z)A�S{��=�}{b/���c���^u�7c%�0�����d�~�&Vj��q���&�܂�_3�_y��p���1�mP�5�.-�7m���%�5����J	���^1��;J��ܱ�9���o9CF,ژv5�b����"��C��f!��n(��ff�{����e.t�J��DDG�δe�]�YI}cr��W a[���E��+ϺE�!�i�V�u�2Y�j�O�/=T�E���~�9x�x����|�mT��F�����6��%V-<�M]��δ"�uh���p=|��^����i�m;��<��xV]gU=k5[]�c_�{��j"֛��,�(>����#\��OZx	�p0��������KK�;s%�o�6��H�d_:�I�"���M^U�$�G����N7[wvu댞�6�Zۊ�6�˂/�{�r*F�C!`,y��	����6N��5:�����⌗k�t2�e�dhեT�z�+���/Й�M��Ƿs��}n%z��jʋM	z{a��u��DY������k9��ygi������-���uc�u����^�UĪ��'�tGlJI=����[fw�!�P|*׶b�U�#�x�|zo5-�,����P��Ij:q򾽳�R!�v��j}�wQt(�P���	��mjˎV��k2;���Ѣb9ξ����7������Vq˕;�y���r���'-���]t���z^�]��B&�l�M�ޅ�Xٞ�Y���YB⪃��~@  �(��s�ߖ���2ձ]^��T@Քk���.ȴ�ˉ��w�3O��tuƵ�2�eF��1<%�������b�ǭ�Qt+�x��4ԃ툞A��Ɓ;�9�f�O(DrϺ��Y=�*���w?a�]�*5�91�2Cjm�:��3٦����Yx��Nm����/d6�I����ڧ�^��ƞ踆� 8I�Wc�/s1��m%ܤ[Ѡ���d�F(�W].ަ_[�g�6'R��U�Vk��[{\���C�J�w_;~�bm�_ay3�j�u����Nt7���Z��:����[����ܸ�x�7Յ�_(
�b��YGE*Nr'���T�7~�����;S*z�K/n!Q�f�)Y5SY՗���9���B��.-6*�U�+A�z9BN'L��YؾO%��H��j:u�~�XtNC<{���T�>�k�X;�n��ե}j<KGS5q��r���^g��s�xO��V,A��*��
��F �%Mս`l��vV�%H0�yb�+����[���#.
L�"�|Vr�<��=ᦘB1�@���*Z����3�A뺗��K�ԩ����rJkcZ�S*�&�a��P�*f�״AF�u�[�����YU\.!9��#�:pI��3pm�cf��O�1��ǵ>���V�hB0�lZGG\�0+��)�����;�F��ǁ�ٺ�h�q6-?�&Y��o�X��yַÖ��<؜y�*��Fxy)���f��U/{���ы�k��w+�`��EpU�d�+�{�-ˆCoJc�iDo�2�d̓,��=�n�s~O��d��S��t4��n�R�EN��������dv[�l=�r����N�L�>�N:;�� �x8e�ݳ����α|+�T|%D����xf����4%{��8�]�����.�'z-�;�������`}�[��P���U�y��>u��MWL��Ł�Z�G��F򯼗�T����[sO}P��5~H�̚�Ԕ��dۚ5��0��3&$K�����[{K��[���e���'��sW�?o7��A�C2�O71d)tV���;38���`�;h��hv��-�p9v�P��Rޫ`���w�ۃ��'j2���3�ouGr��væ��B�V���{Z��.��v��!�tP��Q]$&-�����k����&'���WP$L%Ư�ӵ6�k��r��[�}qD�����'�t�e�Vs�],@��`�ީ��soC~{�QB��2IF�#�wQo�^c�w��Ȑ���i�!��c�=�g�0_g�Z9��1�M�l�Sg��\����Ne���_R��r��ryO6����&J�:��ٜ��*��^�˃�X�:�������SО�'%�N�ʮ�L��Ӊ�35N�c�G���h��K6H��ǚ�u������������˛��o�Gq�S�P -PY�9�/S�ɵ
Z�7���fK]�k�k9B�6��i*n�:�9��x�M�_��L~�r��[/�}�<7���+��!���ON���=�Kk��n�3cq��޻�DM�V��y��`��q˚D.R�x��9�2�L����"�Rl`5Rfw|5��tx��d˹y�Wo��P�1���#����w������+��J�Mv����+�Q��v�jL	vtd�R.9�W��UyH�����Q�T>�����q.��X�5Ի�w�]����u9��#דfv���w�Gh���Ux�Li˥�#2ay.��D1�>�i��Ϧ�e�&}%#��h}ٛ�&���ڦ���&()�����WEax�����=M�];۫����&wF,�wY��3(�� �
���/, ��"��X%SLJP�TAQT�D�MQ%LZ�"�*�(��
B��*�"���j(�"����)"���)(�""P���J��"���(�2�*!"+#	�����(��Y�:��
�)�(f���DD�P��U������(����*i)b�j�����5&F�""�Չ�	����*l����&��9�2�!��
� Ȧ*b��(��Q�EF�Z	��2J0����(�*��))��`���j-a�LTQ%T����UIE1D�4QM&bbL4TQ4PPQ�f9%4QCCDRQAUD�T1%P�LEMQ�ML�TT%RALQAUVfY��P5AC�UAMU4T�%�Y�L�e�TEAM%P�R�ETMf&ENYEAED�DKDL�Q1Tdee������^��חWtn{�@�����K �S���T��C����ĩ[�|Gc����ٕ�bp��-�ܷ�c������o$����謁�q�]�O���&���PF�Uz�Y~�N�>s����R�������qj籔T�9f�pŹ��5�oj���^�O.#5eZhP{]kbGD���4��z��F�>�r�1Ň�^ѫo�-m��_D�Ǚ�y��Y�o؛�Kz>y�z����W�{�׬G��S:��b�U�,y�(z��H��Iy��d�J�M?M��J��)¨aDe+�ƃ�D��5i�v֍z���ή�#��`�vNË��y��o�[�Z��|&kAm7=�NfR���PZu�b׺{S�c�v�+X��CX�R��0@W8�������ϰ����͵uo*#�b�T0|�H�N�B.O�ո����i�5����+nFmz8OeF�������=�9Ef�֭�=��9��{޷��i=���iHL����M���3����b�oUpYD�7��D�����(�.������}��z�2�l�x�L��:s9J��-�ɵ���ս�Mfjjܩ��۲D]�����u�>̚�)�n#�u̬�6�7*����5w M��=�t+9Wo�	|o�Ψ��i�S+
��\p�za㸥s��ڤ��{��z�u<����W���Ĵͺ����ұ_W���E>�c�;�ם���c_��y�����p�]�]��1�[.���:{���C�[��4+�;r��]Jv�����i^U��Ɨ�p"-tj�7�Hy�x�g=뼪��C��&we�k��M'ųӊ��B�y�>�Pb�B��P��A�>�|g�U!�X��,�����=մ��j�+&�3�iդ�^�I�wb4כǮ����[{��)ŵ2�P};�k�5`�羪�UF6��N ���txZݕ�/��v�*�W�%տ%c��u)���g=���g�2AV+gC�;��p����U��:v�D����c��ئ5�=Cu)l���EMoj�wog��ރ����D�ղ�w,���$�'����Ř���]-g.�X��M�\��.1f1��v�S0��l[�
���X6x��)O�bU��6v)����$fF���W�o��aD\��rL��T.D�y�Y���U�@H�\�e���0�A�s$��C��5ܐb��A�z���Mue�H��׳��+ys�ݯ�͉e��݇�Ga�C3��v�l�XJ����A��˔������E��C^W�b��9G0���>��0����E��*�ns�ƺ��ks��+���츁�kƕ՛U̍P����n0U-5uPV�w�4�fb�>���u��W��������w�R�n}}��K�>���`�98�>y��`���c6�����e��0g0�S��3<�{����{�4;z���r{�����E�!�kcr�ԭ��g��F�~�d�՜����Ty�j�Pr��C^�;�j�83FZZ�f��O;�r�Rp뫅B���F�{W��M�,��S�Gn�;��rw��jbh׆Fk��5&����LsJ]g+=r�5�P��=�WM΍n�~A4�;s%�) d�(�n>0��t�<!OOl���W����vv�����AFD�+,���9�f�;��E4�Oq?�-�u��h��)��!�5ԃ�C�iY̓hv]wH�8;q��P�C:�>S-)4n�қgZ�k�}�@��m���S�@C*7�j��k��
��d�뛹b� ��$�V���x�Uꔚ�9g�Z�*�mLr&��s������x�L)gv�'�N����juod����%�Z�TʃD���m��'�
ƹ+��[wT�]�����eE��@{]p�D����]��kU�O�S����[�1�k�1kj�y�:��K�ʸT�UDT����euk��N�U����3GEB<��M�}���<s =b��D`Y���=������x����h�}����Yη�'}�W\dD;�8��o^�+��V6�tۈ�.
��2+�c8�� ��8�b�{!�Ny\�_��ϧ�Y�-}�<�	Z��y� �W/�F��6q,��uW3�9Zܦ�Hz���N���k�
,��[�� -\��-���MCݵ���rͲ�	���뜨��UW��:A��4�C�l=���n���$�힝:k�wK�.�ۈ/'*1@������oa2��R;���ЇJ�z`��Ǽ/�zs�;���9�x�Fl��3V�#m6U_vr4�
T���T@���	ϻ%�,݋�d�uw]��f�Ko;q����=��T\�|�e6(��3Y����x��:��ZyS�oxJI���b�>�H\iv,�S�z�(���胝y&��	�x{�E���'����w�L�լ�D�=kdƽ]5'�!H���[��5�U�4���n�r��Y�[r���P��_�ԛ��m��{���V�ъK��l�J��7|TCi��v�T�,�e�6����T��f^�D-��iUz�J���\�{���rN'���	�jB��ItP�����|t<2n���O���b�6��n�YI��2��=�s���� u-;�S���:ݙC���1j����ފ���\]1ܵmo[����c��}���Z�-���ns�5c!��m@_��w��Lm�D���UĪ�����Ƞ�S:��Z�TɁ��n�M�:��*�ٷ�x�,S^�p�e+��(>N,��y�VN1����Ƶwu�6>�`���Q��P��6�^��Z��F |0
p���͚�p�O}i���t�����/��Qg���910y�mb�Qo	}����$]Aw��Z:NiӜ�ɻ��wg��w����ic�F=�̀,�;��7��q-�VecW���sښ�{�9��9Q�\��)Χ�ʔד��+��ꪜ�L�?C���Z���W?6}����IZ�ECX·D��Qpi���б��sַ�L�~Bv�c�qk0R�g+T0�M�'T��ݚ3���kt�WÃ����R����z� *����iV���p�҂+�C b�89� �V���H� O7bmW�{^�5Y�kWQ���Ъ�.^f輫j���;��u��k�LmzKxI��Z�g��ɗ�/k�z*�+�\�qݮ���v��;y�3�VhW�;r�Y��Ѓڹ�{=�ɢu��ԵQ(Tv����b�$�w�ڨx��C�3q>�ݍ�C���%��4�? V�-lA�J����-$+�Ҥw���@۩���	�����3�w��~a�.�+�m+��Ӫ���N/�C��(gVu�<^��u���qñ^�����2����/����F��"�����(|
�u��Ec=װ��D_W`����`|�+N��f_7/����N����&E�߯}��axi`�{��pU�M�hz��N��!�w>��3hJW�ࢫfu��s��<�͂�р��uԳdC	<<$4�\]��zi�Ϛ��5��9K[���Dj��r}K\��~J�g���+F�Ky����w[�9��疯����,�η��U��:w�K����c���Ƕ.�s6:�42�Z�[�[ܺ�c�n���x}:��DK����ND��n�����ho ������*�W�Ǘ��\b9�k�ڔ��V�p.v�� �dǭZ����Rz��v��,�c�c0���=�5S���J�� �Hq���#�z��U^��+ê_L��a�N�Wzͪ�B�����j��i���C��K��^�p��U�7�V��𸶂��>[�U�R��Ba�]��v�����(A'Ϟ }�lOZ~�%XMߊ������y��p�~��p�+Kƥ�u�OX���v�z��=����*?NH,p��l�OTb�o]p�Q;N�\>wMF�mz<�������bخ��ۗ���ҋI�&#G�'nt��;��;����\���QeY��w���Qun�t���y8�������J������g{��)�畳v�=�t�y��[8Z�+Rb%�s2u����t��#(L��/��v�Bq^�y;og:�������Q0r��:��ws]bc��l5��7������Z����S--ڣ�oh�8�!8�֮�[Y��-܅Y�_��l�TqY��,��A�����4��,ܩ�5�{��U�n4�+Auy���Ng��Pb��q+�)�Zo��'��qN$���L��Z��p���D'ɹ�������ߧݝYm�/s�riw���" x'Ts_��Ս+�Fjv�u=��Q��ג��T+��z�l�*���b�坆�M-ڦ|eN�wڲ�4*���%��m�W����9���Iu���1�}�^ً[gw�:��:�r���V �d�ҫx�5��ѕ��Ky1�Ap�3�lž���G1�<�*4���ⱋ�5n���Ck��*�4q����X|*����v'{U����.B��J�R�}�OHׅ;�R�f���)����1��zu���]>ž�G��H��9��(S�4k����#^sw9�&bo��}��)z��J&Q��y�͎t���+�Z��h�D�3���]8���|7!w;u�1"W�J!�:���u��>��iA����8a7�YϢ!�X{w�I������F���qcs�}�xP��Q��<8�iǼEv�ǹ��nE��[�}�*�r��`���nhc�f��[sM�W[�K��\fkBr�ʹʌL��^��\[� ��O�U`��ץH��e���#v'Z
���e.�|�`}/�ّ��z��g��g���m��r���8=%�~gb��p�R��Hg!:Ǵ��O�l<{�q���X���y�u��[���P��\A��t����2�(m��Z���X��k�*F���ON�C�2a�r��tyY����{_�w?�a+�p�`�|��i!^��y�h>�qs�ڙ��M�tz���ս���61�/n �J�q��m+��N��P�b�ov��
���{���[쎛p���F��a�5Xx����v��$���SwŋC ���Um[�� .��{�jWOP�<�삮�����>O�"�ZJT�m"�_�~ܳ)-�/�6�זul��ڙp돕�hN����\	</^�5P�t�s�����.�p�8��4z����}{�Gj�!fO~��u�o�p�炸}����d�����q�E{F�Kw�M�̬֊�j�v3���'q��Wܗ?we3�S-zUĪ�>���6�b��&_�_mo�y�uP�\���nvw!�Դ�v�*R>��n�3n��R�{�D5Қ��}��U��{�ʬZ��8�_;��G1��'kҠGk�8��+b�8�H�ě��UlˮV�v��[d��W���5�1��� �S�}�9�~��R�d����dmu�v����*{굕�6���V�`����.x7^\�Ώr��Bd	6�z$f�1=�M�jg*��`��E	�����í�L����Tu�G
���.@y�ׂ{_xZL獥Ոc�u�S��"ӽs��RJ�-�x�!�jǺ/�抇�"��^u���eK9���ؗ��D�j{��x��T[���������v��;���qVhV�n��M:��:&�l�ԖuÃ�+���F�qcu<ĉ�/���	���FuR�"�!�[c̍\��% j�p^Y�y��/��}e�+v��=�p��::���_Ξ7|SN�>��Ӗ�A����(�R�{�Ց��=_��yo�rL�M���ޅ7���B�F��o2�c�vU�p�4�z�y�߃���]��k�[��묋�6�Qm&L�w��t��W�XˤCw���s�;�{7'���a�+�U%�X��g:�>v�݂�/}Ў[|F8u�>~���Ǖ�=��)��3�1c�e��N]��V�U�!��^�	����nM/�xa�	u�H&�+���PS|'d�pZp ݰ�GFr�r�qnuZ��;R�r��k�Up&���)U��74�m�yը��b��7�%��k®�/�$�]�r)8�X�˅��ͨ=��ĝ�W��z����G��TYK����A��&��D̊nW.�u&�C1��ӵِVƒ��gn�G27��<��,����"��j�fZ��G7�ujv���=/p��X��I[S[���u��']����7�0#Z�ί,���^\�[�w��N�92�u`�@-E,�ͬ,�Y{ �g-��9#�u�9|�;
��۹+�&�|��@}�F�[ns���/q�F0��1�	��iY9 �҂��n������B�Y>�-�#��:� ��9��Y����QWV0fե���	"�ES��;k4󫢓� {٤�ץ�W��_��-29HĝӲ���\�f�C����f��,ӂl}�EwL�^k/sӍC���/V��GQ�\����p�Tn�k�ؼr<��
���>�!�m�M�مh~G��eǜ��"�U�u��/Op]&�K3Q�y8�:n�({�ⶰ�3<B;	F�{����`�ʭ�=��h�����u���:�d��u=��ЪE�$E��$P�:������t�w�����5vo*RpCp'��殛�mv���'.T �#]ç^��3��pk@Q�5�Mc�nu�.���4���*�[���.�y��G�y�����uv������X�V�v���5�+�˛&z�q�UZ}�`�u[�z���g�R���/i��=5��M�=gj�k�]b8ְ����Rmܭ_�C���Iu!e��n�t��L�tA��� �׹K3R�f5,\{���<=�R<;:u����X�3���Ö]��S�U�c�8�{�IۅJ�����l��[9���Ӹ�k��70ILiZܳC_tX��md���+�#��t�ڱR�R�V%;sLr�1��u���[�%����f[J�C7��c��ɺ3:�G���ᕲ��ri����rQU���,᭝%:��wk.��g'��[~��U�:��%V��3�ׄ]�WbK�u��S|:�hD�����y��R`�>Fl�O]�{yR;�>B�|��a&�9��e�W��Tg6���☣�;��[w+�	]�YSS^�40MPLTT�TS$SL�D�fd��UY�IVF4d�YUBQAUM1PUQ0Se�D�U34�$AY�$VXFFM�ITYaQP�1T�FDMAKAEDE4�fdLQ5BNNSL��Y�EQ4�9�UD�D�D�5UTUTU$SfdIFY�E�c1TDEDD�UDE4�UAEPQMCMDT��QCMD�%A4P0S6a�TEUY�PDDU5TUATAMUM4���QE5T�D�E,D�M5daD�$e�5UVX�E5TPI�HD�%DDQQETSE�feQF!MC��	M%32U&fD�E31TEUE5I1��PK1ETISPSQ1PUR�EPDMRQT5T�PSDDSD�H$A�H$�	e^w��é?p��lo�qp���1�����k��4^��tw6��=\��r_ZG[]t,��ճo��R=z���%��1���?�]N����8�j�+�T�<�mT<Ou��S�xsP���x��칗��/mQ�pn��E$��#��\S{ư�B� ��'�z>�U��C�Thլ�[�WC��U��M,ٴ��9�k��N7[nz�k���JeT2���#F��/��q��RJ�ȶ{cm;�\�ZYy�+�i�O�^8�uo�X�����a�/��Y��7�Z���T����3{#S��;4�D�/a��u�~l�A�rw}:�dY��G9G�-5��<���c��X�lr�v�q*�UN��d��@��J}���Kl����{��LZu�F3ד�����}��H9�ȭC�-��3���#-[���xӾ�~��E}}�H�v%�2��Y���͞"V�f�bu�q��'�"���>��j�m�����Ɵ�W{c�6׮�1~B�^�0W<�S�AXb�w�¸��]��M�V�*@e�{
�2y�Ҳ\�㗖 ]ZQ������k�b��P���k�n��A�,��>��ҹ]�%P�;r�}�%6����;Z�Eʺ��5���}]|��x��>Yk���p����5w�l'��qh\|��hz��Wy5�Z�����U��E���|���=�P�h��ʖ����sP�Y�w5�ːy�����>î��eF���@·u�Ot\CY���Y4i)Z���Rx��R-�p�,��+'�1E�y��U���|μ�z�H���6���r/2�w��]ێGU�¡��_(1�]pIH�,��idjųu�w4k�Tx��M�y�
\G�2>�y���C�:���� zp�%܇36k�����ұۙ0�Z��Ҷ��@�t(êX�ﺣ9��݈]:�Ui�Vڤ�;c����'�s.�Pguf-�3S�4�h�K̾��kFc�/��R0UcK.3S���X�%�Z�T�Z�pXW9�W�������)՛�-m�S!vF�[ڲ�4*��
xO�>�,�E彧4m�2{C
��ʦ�H�>���Q�l���6����Ƅ�:�����o����p���a�ͧ�x��e�CN.��+q�}�n��1.�s6W{Y�����@מ�(e8�	|3tDxp@�,��V�wwR%�z{B���e�>u�\��'~]��,��Eh׷-mz��uc�u�S;{�<�9ŭ��̓�Mf��{�~}��+�C:��[��}��\�W2&䪣5�N2�U�i�mJ��l㸕p�2�����A:��է�F<�y��a��^j�܄`�b�R�Gk��c8�鑮^��q�2�0{r��9�*]�wzǻ%f4��"`lnr=�X�����}I�uA�D�dU��ޖ�^��%��C:��>�KX�p�E���~��,�/�\����v�Ƿ��I�t22�%f��U�w9^��U�+\cR�W8��*�F������G����v&�=7Y�kiu������o��՝��o_$1v�\_[�t�u���{��^;��;y�k��x��q����fD�v�Ovt�O��ۈM�C�[��4')^3k�o*kk���l��X���O"�?>C���s};��O=$���gѼݺy�:����8�c\�8gT��rƥG�@��Hn9�%�po]��'�8�!��G�v�O�s����U�$�ö!}�M����r�1.��Cn�YC�
��u~���ή˴���(��A���TrI��|�xq�L�:ԁ����^]�:ǫ9�F����^��/�U��E���p���;+�%j:���\�ڼ<�쩖�QQ�V�*/o�ZF{=k�����ս�U�F���'iZ������u�~I�8��F��-2{ .��O>��R�J5ͥ����p�k���^��[�SE}�;,1}�u#��ҙ�/�BfE�e���N%���G��\uD�I����{�y2�f�s}�Yw�,Vl�#�y��}@�fԖw,���#��9�$}�=.���k��˦Va�kr5f0u��D��æ�9�
�2��\�+j����?{���v�[�U����mSx2�z����Z�)w(MpY�=�u!��z��]`s;Y��s�ڜ�<�:�w�$Ђ�&<�f5q��m��kN��ͦ�*�N�Ҵ�����"�=��z�c�+w��KC����W˶�	3n䫛}K3�ɥ47ue���v7"���^����Njݑ�f�tYC�����T�'��i��R���}�a��G(���9�r���֖r͕�}�u{��cG2M��eu�72�N��z
/���b��;�o��\��瑎�0U�0��� 0�ds��bRg<mNJpq�A{���L(?v����ix��-���<��抇�"��)M�����!��W�|���g+�R��yO϶���S�����S�U]��D���7؞�a��h�Q�Rt|�����l�~7�_(:��I ]�m)�����SUyך�nQ���L1�����H�%Q��(��Q�)��w:at�K���Ew+T�8s���J�neO(�Ŝ��o��G������MHp�?a	����������=QiL���h�F��W�@��A ����)'��Vw,��YV�
�O�^8�u��G��D��D*��ኛ5��Vs\�(]s]���.�[��Gc�'��Ϥ�Ro�����O/��Sb�g�۴����٥D�Q�I 7[��	
%�Ne�$�*ݓ�zq݊ls�� �>�"�Z��T:G�}}EC�w���}r�ѷ�u	�3�S7�9^u�Z^��*��ryijzq};:��!�[���$�{�*߸?3�{(X�1���e���a���zf�A����f^9�����w��!�
SU�.Zuq��f0b5��D�9U�Ƌ=y��F�Ʒ�T5�9�q�
��R�+��
�W��f;ubQ�<o����rG:C�P��q�ۯ�|@Ǿ��~{����1�6ǻ�Ob-[|9�H��}��Q�}��_\XO�p��a�Z�v�vK�9$q�L���f�����9Ք�����͍Y�k�~L��y[ޑ-I����p��~=s��l��\V���@�w\���9|��a�6��ON��H�l��ݫXw=��E�}:�U���ʭ݊�*M� ��ᚓ�狽Qy�����H��ɚ���C��/�z����Y�YO��o�G�k�On!6�'��u�����j����)}���ń��U��E�Y7���)0y��Aݰ¤��2��1I�������G%+��R��Ls�h"A-����< �ew<�<7����=.e󮰯bݛ1"s6?P�?i��ٽ��{�YaUe�:�Ì����ˑ}���˶TWn	�H�+���zo��L�pɲ��d^S��Ƌ��Mo$3Qsn{z��1iU[H[�Y���z�'��w��9��r������JyN�3��yd_;���1����ƞ�\b���ea%ݗ{�Kx,\��e��;�;,��K��3S��jʋM�T�9����v�\�mo[�wd��%B5����b+��.�#U��HI��z.p��}�	��g7�W�X(wS�J���7Se`L��^:�6���K�˭�����p'�ʛb�ǥ\1(JZ���Q8�v`MwT5V�������!�R��\(�a�l�SV�D2Հw��^��M��J=^ȼ�g�?����^�|��T�
����5�7ήY�~8^��f��~��~ ��'nq�إf,Ҭg5C��q���x�����B��'3R�S�}[`N"vε@c��:��V�)	J5�6�*,���X�6*�Ų��o
��{�cۂ_a��W��m�b���V��Єv	��a*Aw��2�D#N��tL�ei�y�J�mJ]�ĩ}yż1�s{c�=�$WCso��1=y~0���LW����%��fu���ݙ�>�0�ll�&�ܿ���O�W���ۘ���fM�6�K��
2�B�7�yܓU��ҹq�F�qN����5:�F6w��}���	�r��l�k�i��m���w�=�%j	��ȯS�,���/����b��+G���)�|�!R�+�t���{9�R�y�6�ƻްi�ï��s��P��:����+�?� �w���\��^�<Ң�˪��I����ј69��J���#^Tvyd �ˊuW�2�����h�ˡ�r�ߺd mp�1oJۯD�D��_*a�.�,�`I��ܖ�����z�gڷ'�x<K�����hcΰ�j��^����Q��L��;h	W��8�Z��CX��q_��h��X�<J_ޔI#��O_�կ������(�z��!�NJ5�݋���#���Z/�l;}.͞�J�B@ɒ������n��]~e�Ǭż�h�g���3�O^c^��D�Yq�����vn�`g����}��O�L���o�d��xD��F�Ws���뽻r�7��ܢv+xk��-{�'w�&�G��e%jt��nt�:��]��Y�I $+����ó�=l���2��o�M�Я*�vy���2��<i.�6�	��^�xG�L����8��N�ܿb���[`/i\(�T���t����NuedL�ǉm�W�nEB_�5�@��$�Z��囻SZ���j�_n�N�$!�֯lB#^��1c�[���n�#P`�.f��#V(E��ಱ�	n�me�	��Q/z�e�� 鍟�g�y5]�s�67�uH9�q��a�?8�lZ��z�����&��µBk�N�W���Xwb=CdQ�I�ڶ`�@�U8�U�؝�ea�39a��x���.��	,N�����ژ�[�^������IL�S%r�3�=�>=	I�#�Zadp/G���
��W6(s7#�	�H�g�O^�O��U~z�ry.��W�e��`B��x�����5.�plͰ&�;/�Cfʵ�DW�Hi>��;ۧ.e#��v
�\z@Y۟[����5�:;�o7��#���-�ݰ+q��{X#e�%�����W�����q�n�;Hx9ʦkS�ԶEP�o�E���yӚc��b�i���<��չ��D�h�,TOfM9��Md��S�k2{u�'�r�zz-���l��r�eWuT���R��>n��W��a��+"���rCrs˨�f*��<����t�u��W�:��ҳ�B$+p����䲒��j�������)�
J�m���U�P���l��Fl�"p��\V�]-2�7�͊�}J^C
�ld�m�ǊK�Uq4q�8Fu���Z�(3�0A��\���q�/}P��yӺ����
b�ڂ��2#Y�j����.]��9W
���njXb�����9?�+"�e[�m8���Tp
�
���Ȇ�(0�u��du���ݷ���'i#1_kʄ h�c���NrgQ��r��S�M�<�teWwW��E���+������@��W�NM@�.�`�ҙ6xه�?����u��^<[su-/ɔ|`�Bs�݀xԄ�y�r�#W�� ��1��®n!|�ѝ�cj�Mɝ�>]��]{R�	7�Cq2����X���QL�}q������ЕvGwy����L�dJ�MV(j�����M�O��F�����S�����ݭ�=K����W���p�g[�{�����՜�U�� \�~(؛�m?���_��k+���4��w�����qğ8�3�nj������^Y�X5�:��_�3����h+.d޴���g���y���B�0��U�OkNZ���n ƋXGm����te�{Y���;u��wR�cw��_7�jB&�v���Řp����V�	OI�>�
��.E{"�,R4��5��hүTy�5	Q�<g0�g���l�
��q4nbQ���7�����+��ӱq뙪�����לg�n��H%��oGL��r�(QK�\�ym��l}�oě���c���湙*�y�=/-=;ғ�˘�[�7hRth_f@�\�r�s^�SZW5���O.�cע��ӮX�OV��q����{�yW3A,0PO�a���)d��yB3c�4^i���iخ;h�V��^�$rնo�m;�+�.vW�7\� U���^.�
�n ]=�������Op9{ؾ�Z�Q���"���0����%�LX����k��\2+�:�0�#�t���drAdu�ȱ.��-�D�� �5Q�_P��.\�ݧ2u��;&j�G��=u�1J�\����2�p�L�vĬ������;�j�ⓛ]����Z�5LR�2��iv�8���������"I�1��S	�z������Y�xJ�Gd��"ݝ�]�p�!��B۟d��X-�Б4mJ�Co&r�b9��L��U�u������Ϩ������ݦٔc�r�A�v�Ʃ���sB;�{����q�۲{�(�ٵ���R@�y�GQ{��p�y�}�&�n�)�c�Lڷ����	.����s�9+����э���J��Q�ݹ���.S�ɵg�:0d�3��ze���5���f��v��Ao�eYٽ\�v���ZV�e��ڠ-��*3=}��_x��e6�����)UtJ�+.N���]z�Cn�l�:eT]M7u�e�4.kxǵ�H���α%����׌uSpO�с���Ɩ��xEgF6���{.�mΊ#�ERν7aWV�V��jH�+�*5����л�wv)j"���Pv��b�#iљ��r���^ �2�gs,�A�uڟ��;�Y�n;w\��R��p�5�N��n��]�B[o
�w�\{�}m�[{_X�t�,|&jZ��p����m�B��&7�a��`��QٺX�˨L���tr�t�<&�s����0�S}ȉ��U����n��l��cP͇)j��I�μ��u�����B�7T�:d�v�N�FT��4>�Ý�;��::���D}�کtq)�����@,k�x�͗��]'B>��8�z��^W\"�8�](m�r�FL�k�f�� �����:�u�Wn�hr�iwִ���f=���x`�;9�x��ǋ(�WW�-����w��XU�P�3:o��.����V�	(�"������"������i�(�����bJ�����Z
(
****)�*�����f�j�����,�� �
"*(#3
�	(���h$���()bb"������$�*������������3���)i ������"�"J� ���J
��"����(����*�(�&h�)
&",�&�
b"��3"��h���� ������(j"�������h"J�j��H���&�� ��"hi����
�����j�J�����
�JJ�������*0�(�*H��"d��
J��*B���J	��be�*Y������
�(��)*"	����h
���(P�W�P��ǖrf�y����<�^>5�|<}GL��P�3��MY#�4&tK�d�;�drI�!tD�q�5r̀c�a�������ϸ��\�7k����rUa���p7����J�Әw2�ҬsxW��>e��^���.�u���5�i:��0�>�_�iL�z���D�J��\Q�ȭw����p��V1�;U��$Uí�ͯL������=5���`ͼ����̐�-���fj����(u�y�YC���l�0�K�+����O�<�o"��c���j��\�
��{/K�=>�s��/�����MF*r*8�H#G�x:��>.����c���m���X�"���z�Z&aH��qx�;��)#C���
tz3ib�rH@��O�V̫��>�qk.�ர# ��n��r�q�Q���7�6LB{Q��bC{J�v��.-�����Z����& ��h.��ұ�2ǁ�_gի8�s��O4y��{9`��e���#�}q�{�:U�X65ma��V{,y��:^vOsq�
�iz����
�K�et��R�H�P2;�d�]a�۳�����+i�K�8�n�_��ub�e����W�
�k�[��o=
r�)�4�m6ش��=���2M��̔��J�I�e���'@��a����ޣ�-|3����hxc���#���Bq�W�}Urg8�;��@���-�T��TQI����
�掽�z���LkZg��X�1�i�3'�,!n3Ko^ƹm�0��g4L��LXL&TNw1P�22f���@�D�K/._�8f(�]�/=snb���\��d�2��&kP�1��9PT;e�Q=�x�¾�8�y+��%��� 5>�p�4p����h)�u[<���0�J����ުĽ-��?s{���Ju�Xky�I���<�`���\Ɏ��x���[�^�W�C�ٜ+y"��23y[��U�F|���i���U���Ǌ|�����e�k�l@��޹�g�9ќ�v�x�Ͱ�.y�ꋚyպ1����c�Tԙ�1�R/YZ�;/��gx�����f ���ȬO�<Ys�����C�F�y^V��!���$]+u��T~�F6d�{�7�;��uɈ�z���da������ve�M}'T���]7��R���v�s]�`��gW$,eW6��h�
U�ӝς�(���7�){��ז��KN�۔G���A�C�i���]Z|V���%j��DL��{^�1���h�uJ�a��LJ�t�:�I2"�O��\ة*�9@�n��Ur	s��n&_l��d&�E�/���#F{[�<�z�Mǽ4�Qw
�}w]մ�&������?�j�!�\��R��z�o��a�v{�.��_{��Wru����y�8�9��+:ſ�-�g���%�u}��XZu�-��7T���뻳[+�
�}�w[�����ثU�%/҉$u[�_�M�lby��M��y_{s�;������P<�.�@^�Xw�޻6z�+��&��D�x,b�4�Q�f�{&��hƠ����L(]���Oj��W��N�k�g"��z -�vN�Tǯ�3WowcD��i`s�V�!����)���I�ѕ�3CcĶ�+�7"�>\E��ꇢi�V���m#� ��F�W	p�6�Ϛ�3��n;���a*fV�]�U�>뭣2w�>��D1����Ց��>vT��Q�qQ�~|ELm���Cgi�� �:׷�{3:���Lz�%xoK&j
����ө��2���a�"���|K;%Q�'1?V����S�t2�FyV(�.�8Ibt���-�KhD�s�v�'���ã +8m)"���5]
F�Ԁ��K7]�����۫��ż�5{D�H�����X��#���%s�uw��{.`3g�^�T�i֣��]38S���P�nP���R,��D�v�K�R͑�f��j����x�̠k��@@�ȒJ4��7��{s� �<�^�	z�b��_ܟ*�*��13pٍJ�#2ZU�����k,���ܸ~�/�y��XN��2�`U��ʧ��sR�븹�hҜ�����������-�ε.�ي���s=.��� � =��gx�i��i�=�����3���8�����Mh���<O�9��X����~��ʾ;L�v��sy�z��o�Ɗ����ۼ���1�b:�B�u�r����)�
J�g�F�p�� d�H5��V�c�j���w݈
��ѩ�E�o�	�)y�l޸9#�����16�g����c29�v��vQ�U��W�t�1{��Ux�S�<���d���[��V]�z�'ay��;�w�X�w,�/��*G�R�f��:9;�B�i��S���B��oZ~�ǝ6�ZŸ�;E�#؉�T"�aY�_{�T>4ud]����g��~�k:tY�]z���h�RRp�U���h��WA}Ү���.W-�z�����Պ��er�)�[��b�����p�
���5Oؒ�d���q�TV��ZW�P�5�� ���e�J�r�RVpH8D�r��0����-���d�y���Mv���A�a.iܠ�n����Brd6�r7� �Mv�S�o'}�q\س`���'<ʨF�J�n��m�8	�&�_�{�"vMX�\�Iw�^���M1��V��F�A�Jʦ��rLG	/r*��L�#_N�����-�ӣ�"�c'��J��k�5��{[F�����X��M�5_P�Cs�����B�#Ӯ����7Fə�=�vVXzJ�>~��;c��mU��;��
"�
`ׂ`��~(�Zc�߈7�{��eM�۵�h��|]��QÀ��e�[��Xގ�����"QQ+3�Y���NZ����w��L�y�,v�f�!���0�3�%ծE�>N�O"L�~U�j>l�5|�������>u�o{��\s[����ސ�s�Z��V��/}R�YSkR�|�@��V�˶����F.#�r��R�q7p�:��G4
B9~b���Q�C+�����f��2�>� D��!Q��X�Ȩ��!p������M���t�H�:�QV���r��f>���p���ҋ���X������T:mq�1����FLUs�l�C�y��n�)�z+^ժ�@��ݲ�a([����7��1g-0ҳݏ�bh�O>�aˡ�Q&�[������uFs
�';���yN�����y��6��G!5�L�̊���$b�.�GJ�t2�-W�|��#6m$�mޫyF��*�4����@=0���A��mRKJ�aǚ���Zi}��Pָ�Q�+��ɗ�6xU���rq���9�j���FඹO�� �X��V�|1�viX�c�����|%�%K�=�A"���2w�����|Y��R�r0b�q�ҭ:]W��P�u�����-��P�rȨ;��c*Z����*e���6X޽�l����:F�|�;V�e)��ڨ��lm���=;[��]���}���,%���7�ָ���vٖC� ϒ��*9j����îʓ�X���r����U�l扑�O�&V�^�T%��4'W�ju��=��JW/9�]��@eW�=�/�]l���%i���t��P79PW���tKw�.��t<�
�Phϧ��e�x�0:�k���.�8xL�x%o�e�<�C�QX�f�
�[����3��:Y���I�8@u�<�`�^AU�+��w�{�{!C�˷Դ��-'����'��n᧕�v�$� ��,/m��>G�M�ΏrL^���>��$��7%�0�ɝ��{v&���[Feu�wR"�((u=^�����}x+Y�]��4d[yu��Z=�֍����.��b�~��wr*x�G;���1ss�s�&�y:�«��wuK�=)7,�w'h�ל�9P���D����q.q��N���}Qr�`���3{�1�*SX�Uu�=RN��^���$s�>HV�2�@>�Z��(9Rf/��.�Z6s��2J����o��{q@�\S��t{�h
�j��׽`�C�0�k��`u;2�æ�_�Y��с��j��y�z��tx^cj3���'�ۜn��;�WP�:�ς"�ݚ6�zjL��x�l�Az���9#�}�P�o�{�7�[�)*=�tΜB��9+%�0�@$�dY�\벒��WXP�خ=����]`y��Q��Ӫ�_�u.=�H�����.�M�Y�����!O�!\@��n�����|����k�l�Ŗ�۽��^MO����H;���:�<)��B��Xv��̓։\�@ɒ��u?u�<�sNI�E�z�TC{1�;U[At��$NvJ�dx��.��m���^�Zni�=���m�E7zW*�2�:@��,����^=�b��D�y�&x�����,�ME�wET����W^��0�T����loc9�u�vF�~�>5�r�I�W"7U�o�:.�����k*ļ���ސ���ft�w�"g=D6髩�Վ�X����:$�R�ڊEA�����n���&4`����J͙y~�Y�h��r����s2�t���S�zf�(*�G�g&O �~^؄F�e�b�]��bh��uu�����5����/�T�J�LL���Ѿ|��J���+4������TOY����ZS�u�1��T�r3(ҧ3 �����|p�ѹ���9�uy&�4���{FHA|bll�#<��P5���s�����kő^zd$;�Q7���fn�=�٦������oO�[څq��q%�aHCac�}~��^�G�6�%I^�t1�N�֓���=��N��
�v��j�/��F.#�Z�K��ٛ7��\����S�q��/�x���C<#z�޾�6�f��q,y�"t��T�eC�Ց��Y5qH�B�mU�nD�)�x�dv��C�_+Ա�n���x�6a�A�}���k%#�[]ه�2��
���h�r�]tܾGh,yN@�B���j��5p
E(�]�zm����Ʀ�l����R��*ٸ�$u��R U�L�.�S�x%��*��2���63٭��&m�EH99�8�aԡ����M��u(���{���Ͻ�[:���Bu��7����z�Vm�%��g�l��'C�F��]��� ��x�����`Q|��H]�]G;���k�ʳ]���)cK���B�\Q7�勞����ihd߳J��[P*9m���:�B�V����qʬ�.]Q�;O��L�����-��Z핀oy���|�`���S�� K��Ǟ��K8kb��ĺ�3��"j<�E���/���}��miBwNZ�����3�'�z�$�P�49�\�GiI���m�"�Z��B�;�ؕ«6����v�v_����K�#R%�y��s~�&����M��j��=���J��K�sS��^��`C��STF�LGė��U���3��`Ŝӣ�+�1�3.qCӻ+�;"�o����O՘�L�Ѷj�7^ڟ�qP��ƨ�
�nu��s�Ǌ!��hq�nm�P�W/5$�*��8�aT ^�ҽڇ��ʫ5�O!@d��O��N��eHi 6~��Oof����춑z`��.�Op���@nWC*��lx�)�օ$;!>�X�u;���\n,����j���)�P�5�#&���FPz3A�sT_i�})d��P�N��v����o��.��kZu��6N��Z]CN�tB�`�=�tۃ�iR�����_p�V�8�E�]Xx�>��r��y�it����ˏsOQ����q�ݷZ/���n�	YϠ�2�6���`m�%�o��_r6w(�'ؓ�z;鲼fne�и�@Mz|bZCϹ�H:�}^Kw��z�7��2k�y���?R3&7��qĩS~DԹ܄����'9�o�J7�Ut�h�+��n��z��A�b�R��W��DױS�^�.R
���8:�6��t�H�1�U�Uwy�3=��1l�
6+��_r�0'��Ef��xZ�����`�M+�,�I��u{��.�ڥ�p��L��8࿃G�ʦ���l������+.�N�%sl���\k��d	2�l�+/�T)��(�_��J��C���3�J��ұ�2ǃ���C�,\ ~�[�_di��
u�hn7NL��6W�1,W���\~Y�po��j��V�hv��}\S*l�n{v+G쏫��CG ޽�l>�p�D��0g9��ڵ�a�\���5�t:����7}���@�B�e����2��!Q=AM7U�`YS,� ϒ��݀F�v� i=8�ye;<rK��zǪߺ?b%�v�%���b�,(׉����}���P��]ܸVb[�TsoEE�0LE�Wt�gX��ΖR�l�n�:(O;��٘�ޒݏ�)�[�tW�l״w�(e��EM��{^�vYGm��W��c�|�5�I��K�U��
��JA�+N�J���fj�9[�-iFolH<ي�e��O���N�����6�}��y����y۩g"�s��­��j�9��J��\V9}{b���������o��^��ҡ����C�^�t�{�ǖkb
z�1{4��%6m6�����N�c� ��ǫ1Z��0]6.��;R�>z���2Ԯ�d"=��q��G�)w7l�듟	��F"Ԗ1x2�飝��K�tz≑����o_{ޓ�=wR�Q�]�;���@��g�NMڝ�O��z���M�[0c��)Ի+7;C��k,aT������J��a/��}D2V������p�5�p�̷���>�lb�Î�����{;[�S��f�=�7�9p������
la������Cu�ۥqb#[�]|��ũZN��Pxq����n��h'L"�&ZT1�f<T��?>��R���-nl�MN��yl�z6Wv�ChRډX��-�+���ﻏwtT��9[���Q��i�ٖ(C�1Cz���+%�e{���Q�L�N�G�(�\7�L|1�����E
`�Ӭ	ks^gn�]Լ��榞�"�:ܼ{uv5̗�w�sSJE�x���[yt=A>W	ڎ14�K�b�ֽ��º�*�/L�g2d����'���Im7U��Cg��1�����`\q����sF3}�t�ɳ�vj��[Ű$�����vz���-��H��$Ƿ5�3;u�eur�-�\R8,����^�A�ۓ!H�2<�U�s8���iwh���&\)�F���#:���O��ҮSJ΍��@��{2�Rge���X�xG]����%Ċ���Q�,��ْ��I�yVV<���C�]1&��PR��2��f��-Νc�=�wR�;��r:2���dޡ���ܭ�5��h����p���������l@�:[���b��G�E�G]Ӣ)���n������]t�B���B�<;mK+G+�չ��\n�w��N������K�v�	=��5�]���>�lZ~�5x`��:Vn���(fήᵂ����8��9���[ɗ�%�âosa]ܢ�T��s���A�:���<�-��V���gn�� ܵ��BP�fC�Xϡ]wu��x/[ɲ��Jл�}Ж��Bƾ�7l��}ц�s�^�0y���d��B��}:�JY���Y;��N�mi�C��6j:(65Τ�%�Vq�=�o6똕u���)���y�Wb�1�."bǶw�e[�^���=���oN��1]��Θ6 ��vɯX��6�a5��,�Wo�$�78=�KSu���*�ݻ6p�y4��r��r�T\��n�L�?C����+�:C}`�`�7�
��wp��|u��EC�d�Nf%��UL�LHSHUABU�AUST�R4�ŐP4ĭPMAAADT�M���Q���`�RT�QMHU!E4#E4�Y.Y4RSMRPS-�PP�$�!EPDEVX�1UD0D1UQI4�515AHUNX�DTR�TDAU5D�5�fA�Q��R�RPU�aMU4d�a��U5��Qj2��X���%Q��2\��
X�"�i)
i�kX�X�$�Y��UM5�PTTD�Fe9FM�ՄITRe��M-$E1 }D  P U3��o�Px�C/�N������3�wY����<Ĭ@�Y��1K�H��[��Rn�x��B���*��\]	�zɊ�.s���s�[#�&�����5>9�8��^y���@��`&����k�ѣg;-�)���>�����wFG���^#�k���*Ӈ���7������J8�l���fl[�B�c���h��Ü��h����cƀ#�+��:.�m��:x9�V�r���x�-��2qZ�>
�F4��KG	/F�<W�NI}�0�W�( 0a��뼬���x������P���ԡ���T=�Q`u�LR$�_���ȁ������{�&}<��{���= �(��J�W��Ƚ\��|�&�酣eٹǏnx�5���î��0i
��t�96&c�
��U�!k0x$�B�r�2��u��.� ��,��~��z�ڮ���{K�\��L��-�L��S!�-o"h_uqc7i�uc7�QJn�WQ�gSɠ���CN�|���s^�����ڧ�'��_Z��V��@��sEZ7�>^2uI~L�A˝�A��js�`�1+���uX���X����PX�����$g5�
%\��Q�i�́��ES�+��y���g����^��ȪbJ�����|e�a+~N��ӣ�e�޹��̷7�BLC��v8�+����wwV�����IfP��Fu�kU�.��/u�pW7l�c���w�Z",�˷����X��9!���;+E�Vf�_
B����<���U�e�wkuit��c�b��^�{q�3�ٯԉ�k��fS�xl|��,ީj��,;�컋�y���W7��rd˹����D��TH`R���XX7��Ȝ��%��T�I���r��0�4�3{����N�m��
z�4���D�i��׏y0k��O�r�#5΁�9��f�B�g�
ke+��� �=�Z��Yl�(��S�Qe���MNJˌ���V�� �p�W��j�C�2�5\��\��q7V�m��:L�g@x�%�6��3z�42����Q��؇Q	U�L���Wl�|&���^i�vT穼;��	숪�d��/1�n�YR:1�;b2o�y��-gؠ<���u�8I`M����MW����g���O��;'wG�Mz���J�-�p�,����^��j|��ϫ��u�X��Ԙ�5���G5�^�"�]�~�yL	&���*S�Z����	~c�o9�K�'½���[�|�D�%چg�����S�Ahw׽��w��]c��T-5��~WFYr���A�����"3uu������<w9�HXw<+��Y�-�$�O�/��S�f}M��
d�>��.�Ͷ{�zL�R�O�י%��Zɲ�&WQ��ܣ;#�v�㨭0��9'n�^6���H���wS�m4��۰Q�V����2��9��13�2e�� XƮ\��c�!�gp�_�)O��w\T!���w�VkP�PȔ��8Cxm��+;V^L��pX�L��~^*8�Jѫ�Ct��%�v��yN@�B���Ƃ�mH%�-�ry@Mf�Y��,H:���`�Q�\�2�7|Ю�\d<�ˆ���%(0�uY���ge̙�׍� 1�a�1b����j���v1����.��đ&��	!k��Z���0?%e;�eIx��o�O��`�|�Ż2������;�iۥM�Y�۽X�s)�=��۾C{���ѐd�d�|������B/�Fȩ��M�X��)���/׉l�=�}Ԑ�#�+Нړ6Y�"��-�`I�P<�N�p�LWA}7�̶��ӻ��׾ME'�wޠ��o�b��םs�(��*�'���=tWs�����`�Su��*�{dU'��rT��ueJ#���uMQ�q&�܊���^Fs���e�@�<��Q�����h�C��
�8 A�N��������G�Z��&��/f,d��;o/dށ���p~[�.#���=���1�x�r���*�Q��,��M��C7���6ȑ�x:=���:q֥�,��z�1?�T������ى\�#�m�{J7��Xnyx�>�j�p1�"��&��:':J@�VT�!u󹼽����(�;n����:9cQzp�y��<���*��X~B�@����D�n�\�/~y6�M�o4U�.8�Y�q�`߫�����s>��Y�¹�����Pʭ0�6<E�v�8��#��$���糝��b�8��3��2������	�H�\��LM�ތ����S6�x*��l;�o@�w���hl�c�'u/�D>u��n�l��%>='�'�B95�Wgw�2��j��6�pD�?mC�9�Bk܏1p�r��taΒ��Η�p	u��^+�5����,ek��o��4��S���}����UQ�U�E�a�>{��M�6��s%ծ=)�����ng�{���P(p�ѱ\'�!ܥ
#f�Ӈ��.���7�uԥ�5�f�zr֠7hV��3�6�W��%�8HՑa�5<�_w`�giq�F���.�k8�
<ݕ�.���W�ڎ��Q��&'��t �ObF��M^��a�J��2�+�e$3TXG�I���0Vľ�ھ�ͫ�r��;���&���:�=��urC��|�a����-�\�&]��*T�b�ڜ�NN��kC�����"�8U��˒�`Ĕ�p�\�'G���u&��M��^���9�X���r篫)C3yG�o�~���,���K�������� �_�¼�W~���z��R��"�Ϊ����3��\��U�P4�tÜ��W�;�p�䬒:��I��l���/yr�Byϻ�,*���(L�F���<|���e����p��ŋ�DƇ��ceE��l�Y�wlC��i`s�u�R��j�g9�,�e@� �ʉ��*:)�ԕ���-pk8�c���;�,v5������P՞x#�8���Ze��L���Kr�?���zk����R�"\FZ�	+:"n�Ȩ*�K�����J�Y�Է�&'g��wk�C)#�;ұ�������&2Bc\%1�<	���ð'V6��_�W��~D
�XS���Ƕ���K.7��ʺ�z��cc'%�g��\�jt���'V6�	�J|�|NY�YY�fm��gd�)�1���a���ܡ/�O�X�p�^����%^��[9����_"7ouvE9I��$��1���X��B���=�'������Ƚ��;M���ӷm =j�wPU�m���>EkM����!��Hp��a:�xm`�9BԈ/2�9�ٝ�%���X��A�-�)9���[�A��Cx�XJ���C���/�s���b]X3��A��i��{�e'F���F�+���X²6�W1T\��R_e멽k���+�;��1�S����+����0��rY�úV�V2Fן�����:�_w<\�Wƅ�J�e�5u:5�X�K�x��l㢂T>�=�2�->�U蝢dє�v���k�r�uN��lv�g��/�5�^tvy)u
W�,�� ���Q<9To;5�z���!z�V.����un�.�f_��V�`߰�Þ���=��9���SC�y:��t��{����0˷�'6��h[������w�Z�����ç�X�N�o�5W+���H�tg�nߣ��פ�j�߼5g�>��]��G��Aμ6��z��ז�UE�����f.����ޢV��;�<��Dv#
�^:(/v�s��2��T����/�^���\������lѳ箽�xs��#%�Nh�!�����Z��gV�`���*�C��Pv5�����@[���P��Z���<�\�>���cC���׬��:��Xn*$5(}��9���;7�W�3qWۮ$�p��AhM���VF����ܻ��k���l���E]~k*i�qJ��8pd�����ʕT����rV�}�������W��޳V�+���;Y�4�:n���d��^J�`3��X�}w�i�}b���B�tWŻ;t����h�n����~�V�k�=�7�D0��ý-CR�Vt��i�|��d�f�.�H����؇^n���fe�p���,�XV��m9�ʚ�]{յ˞�Ȍ��I�ҽ�p���fq�_��Lv��3ʀ����p����	��Q�ICޚ��mos��[$��(��O�+<�E8|�_���(v��C��
����X(��^']OM�.89le��e06�&��j�l�O��0*��0Ɨ2}�6_����[X+Bw=��2�������J�y�_Z�u=&���2�Pw��|�^d��	S^ L�,��C�y���i	�b7E{�h,UW/��q�=�|7%֤8�j'({z�g,0�G0/9�Z}�#��*��bU3X˘��W�F�yS���S��71�n��WI���[���4E�
�bB�r`���Sl6��B}J^y�Z�s��J��q��ɾ��0�%{�o�cUh�4z*�iM�`�K�������p�2����6fv,%]��C2gec�P�q(��2d���'5���k�`�ݘ�haŽ,{��#}s.�S?j��ڎ���oZ�IWe�+�Z�w�X�7�3��~��6�Ձ��M>Z��(]γ�Ɠ|3pQ�ۜ���*������D+�u8�Ÿ��D��3x=���Wb��"�{�g��x޴�^�x��Ե��үI�yWv��Ew'���9�I�U�J����*��(�2p�z���?
�*0vJT���)h�Y�����8)�a�L-��+�ݩ3e�h_��S�bGiIኁ�B��f�/���P�n22mi}+��ܕ��y�L����.~+,�3�(��*�6����=tWs����Ѧ��	yԳ}��s���σ~�wV��,x!��k�L�%�EP؉��g?�̽G�j��l��g��u�U+�:;cV��Kf1�nyX^"WeSU���W�B��*G��K�x/bc�RF'q��.
6.��t�S9�D^�6uz-�8r�ʫ2ư�E{\Dkp�s�9շ��j�d\���Z%%g���D��.|:���r����rF�R�j�\�G�)C��˻�N1�;��O��9g��}�q�n�,�]��N�1����Պ*���-��RL�̼+�n̿E�M�y�D��;�|2:ɷ��#�9�&���8-���#��`ґ�3�y�gD�S6u�/ݴ�űo769�0��/�pӭ��;���ƪT:藫޺iT�/Y�=�7��,�i�5{�ưh��i��NmF�����i��.��s֖:/v��=.��G	h��(g�#LJ�{��s��}��t��._+��r��kΕ���/c0$}n��t�o]�zA:�����l+g홙x�\ν��F�7�N�����qx{z�����ī��ꕳ�]��*��%{hڵ���E_
O�-H*vf�9��U#��';��b�ϻ���bz jFlmվ�
�X9s{"8ޣIy@$|���T$jذ馧�K䶨�J��=�p������=L͜z�uw����<�@E�4���Q_��{���AZ�č�ښ�M����_C��gZכ4b�p�{~�>�f��z����\,�k)i�*��=�LQM�H�S<�.���&�-��]B�A��I�8>�Z�=�״�����oþ& +���{�¨Ox��՚Sk������a�ꭚ�)��ǂ�(c,%-/X,tC\p�r��x�C{Dt�3ۜ���vͰ5R(}{8�6-yت��~��4z�/�y(��h���y��Rk�v�n�S��LY5_`5��m �P��L��%a�V�{%i����]ccq���F��AkC:$�D�����6[���Q��ћ�:?P����u�\��;|Ϡ"�>\�Y�v���;{Yxz㳣�0��#�NT��j�Z(�R���}5�A�����}��w�^�՘K��֟�����t����e��_KR=ΣR�&_v��
V�m>�b����b�f�C���/ipI8��_��Y���EWIfVw���@�[Ƙ�j:/��c���d��U��L��"�C����$>��uclq��aU��e���bhA=te	1kySO�k�4Lz�Ŏ���W���Ħ~O�d��^�'V6�MzS�5�(i��U��R����_����vpBuZ��ש�+N��mT=�3�yS�{�̕������ӡF_�������CmR��U|<�؂����j|�/r�.q��T�7�poOuM��:�W�yZB�t�zY�úV��u{
��oJ�g�,�E�=�d��o��%��GUaq�nV�*R���1���W,���2�->�U��y�%��F^M���f�D���̼�L�ԫ�؆��T��{����.�e.If�C��{�7�Y�`��*yJ`�s��s�ƭQ���t�������<�:z(�զ��5����G�h�'��U����+����z��:V"� �vT�j�n4CC/�щ�2��1����e�z�D�{.v�ok� ��U�.>�B}�gj�d�v��̠�^�G5KU}ya��{�� 2J�5I6�m����]�K�v���I�]3]F�e^ӳ
g31����.� �ث�;{n����%��X��8I��ЉN���ʺ��sJgc�|����XS�)+&z��C؉����Ř��.�')=�Y�8ϖ��;��U.��$�V9��ᤁ�|�	>5��t5�0���Ϥ����X�f�p6�(�
`?X�B������d-�n�jH��;�1*Z6� ��+� �3�Gc(�n���V���3��[uk�;闭�|2����k6n�Z��a�A�Ƀ>�<rh���C�U����#U׽`ެ��3m�Z�b�X���oVI��y�����±�E1b���/��F��]�нBLB�7��ݓ��+��]t0�Z2�r�x�|R^�BJ{l��w�}�8��B"D��3���fK[��q^�f�g�ͨ���5�%�Y����s���1+9��p=l�'�̻E�c�$�SD�c�	��*�p}�/P�<��҄�co)�\9���/�U���q���JU��v�cǓ��w�=]e����7~|�L.�����޷��]w:��[-Ç�=��9Ȧ��>�;�_iA*
��]�nV�"������(f����Y�v	�2��_;\ħ�ӮQ,�kB�7:�&����e*`Ea��ې���d�fڵ+�5,Q�omI-�%r�޽�{[j�N��Ud��WB�Dk{6q��5��p�csJ����e;��ŷ�[��z��*y�5��J���57z%�a)�Meb6��zkbLev3��n���3�_�ȗj�
�ئ�ң���y\W���kM��*��	�j�B.,_[�U��f����3���\��Y��ˋ�JͿ��h'`M�O=x�R�oWd�63KQ��RT \����k�v�o_D7.H���jI����c+�,!rJr�����b�nȤ�P:U�>{�>jb<A�
�_�����f�3%�ܒ�m��GW\���}�}�qU�BKf�ʹ�A�w�&&��Q�b��͡�3�L�]w}��8PgC-Seg�=��{�5����{��&�Kb]7��jt�d�Y�15Ҳ7E�Ofؖ3.�<x��n��t�5��h�;�5���73��u+y� f
'c�*��ǎ���(�t�f䷇�Z<k6;i��Q֪���}�%�E���:)����8���f��U��l̬͒��2M��FM7Jtb��5�҃X��_;��C���C1��/L�I8�k:�Op�G֚{�e��;F\No_`]�d��Nűc�˷	��V�;��V���>^T�i3�l�;YL��2�	w!h��#aoj�����u��wK���G�Ui�*�)ud�pXќ����>����{���¶wD��ƭ��ˡÂ�s���+air���]��My��3�j}G\#Fљ��ܽZR�TI��ETI����5Y�LFA�Mق�UTU$IE%&Xd9DRU���P��PS�`ffTRP�SQTI����LD��]f��E4�M#EL��3(����2"��)��#0Ɉ"f,��b�i�H����,b	������"��"g#"�,̠����22���Jmba%D�ǰ
�+�VQY4DQ��D�Z�(���JR��h������(���%�����i*h(�+&�����#
ij!�5dQ0STSM5AD�4�CM�	ՅD�LDEI��UQ�QI��!3��޻���}ϯ�s�q�[�4�l�^	ݛu5����qv�tm��W�0$��*E�&�7�#z��j�9�#�� N�S�}x��-��y���T�@{Ҭ�)R��O"����d�wd���!�������i�{=�M��6�*5��X�d3��V�����-8B4��&r�e���Qy�\���DL�S]�/�?\Hs˨T6�� w��d����6�DKB�\��9�ˬ��ڭ��\������DW�A��.��}6���udn��eN%�vn�3����.ś�^����GP�6!W��SU�s&:P���L�#�6�����J��շ�s��%�*Fa�2y�*�,7-2�}�a#<�b��\�/ó�w��Yio0�%����M�.��z�0oѭ!����U��@3O=0c�.��x1l.������6uUa�]ސVu\�G;�ʹc@}�I�B�����M7���z}��/�VT	���r�{��O=9�>bF�#��ٲŝ:E/�[���i�~݂���xa~�?܊R���=|�����w�?����Ur� �!M<O�;b��:c0_���VpbY}W�QW��WP�T������OoY���m����i�Sk��̴�є�޺����/+Ѕ��r�`b��z�K���c�g�����LDp�:�������K���*�{ �,�Y��-�p���M���Z��>=�]sϺ�b�ұ�K	���fm04)�p�\��])����	�r ��,����9ڝ�[��A��~`�p��!��X`�Q���0�+�|�O���U�h|M�"�qU��g��nҽӥ%*Uq#�~�y���c�gh>�x�j�);�񫣪��:�]�w��P�R5���@ɒ�<K��p���
7�.ݙ_�ӻ)��=��ƽG����=S"����]�<$�J+�d,y�=I�����B�o���:����9���Wi��x�2<��
����6u�A�R*I���P��ՙ��H�[�6��&t�I�AA}���'Ǐ�ŀ(�VY|g&Q��IT!�������d`�c󘷓B.�sշ��:�Y���w��suMQ�_^�U�+����7gB����n�K�������g�5;cT��٬X�s�Ǘ���T�b�cT��^�;�����=U�Ofet�V��9�#M@E]wFG��Ld��`�9�[���2�̽a����9�d�{/.`��]ky��!�S��^�)�����,�1X����=r��;�����`.�={d��ĂQ�c�{�F_m�k�-9���c�!_N��[V��p��=��s�e�50�r��݅4Xo)=��`}%T���S����(���dH"D9s�I�V�
��_�<ql	�M�h���E^9b&�f/\�VcRƹ.*��PU��'V���K�&2j9��o�F�c�ɸ��j�ZI�}�B�X���&6��y��1���Q���s&0�6��.>�~N�_|�&������s�M>=' +��n��p�������
^�����fPݘ����(l{�no��{���+X��ٳ���"���� b|��8�A�Ѿ����|��ux��=�@׺�'s�D�8�k��<f&���5�����ֺ��rz�EC���:�#�l�; O_;��0u�T�s1����Ẻz�ݹ�*
wћK�$��	ë|tXh�����tmJ�|���{[=/p��I�3��w���(E�4��R�ǹ�{�GB
��$o^�����K�[�>{��ӛ�8y�<�5�Y��C�^��(�Zd���=��@��ҡ��8�g&��(����M�h+�?-#�5��8��xXO��'Ի�x_��v*Ν�#o�Z�y�����zR��n�kEմ�oA~>�%!�~�wk�U�E^o�I��G�l��Y�Wק�ܷM�!���+���@�{1����G%w�S�wf[�n�{=t�7��\�\��{�������ڦ����J���{��s��)�%���s�I�psd�Sl;��k�ԉ���p��iKK�X��;ϸ]�̠��c5Q�ܲ��Բ�;��2��g�]x�5�C�F�v*��W�W�<������if�dOc4^w��lkyH��U�����f5�j���H3�|�g$��3�mC�y1��4�F����}ɜ�
PP��T�o6`dTt%� j}^bt\�+s���l]W<	����4�)���f`r��ޞ���;�ucn�*u�Ux��%F�5^���oϖإ~���CuPʺ����+���r��1�,�����5ZI<ck�S*���.Ivڐp�.C�o�����s(u����1Ϫ���ꋘ��1�`�Ec[ݏoU�pM����u&�b.�4Y�X� �����b#�ZW/D{�����K|��ǵ�<��*=&u�+�Z!`��W��,�9�ˡ���^���P�[��SzPr�3��j�r��]�G`��:�dT���<T�6q�@:b���c�<�X�^d�����J�tVoH��G������ڝ�Aie�uϩl�]��>�xn��Nѡ<�	���E�Y�V�-� +u|V5%.^9u;3ܫ��6���󺽸����K�9���Q��1��n��tG屋&��<���Wt�yh��%&NP�ꝯ�o1"g�л�t1���N������*;<�p���T�^9���]Vjd�R��;�H5�y;���ow����ި��~�b��Hè;zS�ڜ�ptk+������F��ZW"�ɚʻ��C�J��	����4jva�k��~�ղ&��ݜl�˅�	��U�b��ۛ��,��I"P�4������R'ݮǕ�Aμ6�E���]��4�5N�V�Wg=���3ҰL�*���G��;�Ȱ���k��Nu�3�@*���Y�3t���m^jr�XJ�	��^�Ea��i�*'jӄ#A�������r�D=�6i��2g�����x����B\�� �]F�&��K8e���{s��tS`ǧ�{�U�ڡC��R��kt�� ��s˪�|E�KG*
7!��UN���3&����v?�Hϝ1-Yv�P*���Lu�	+�Q>�´jv��GU�k+�%��\5Y!�6yL�^%،��{*��	x6\J#|��*U�� �
��jI����y��Q�;Lk����`xv*��V,U.�y�7�A�*�5���d�L
��Φ{R�IAp�ɭѫ�+��+�3���Rtѕ.�����+)Ȑ%t޴=b��Xzz�bC]r{�u�}�]��.�zK���m�wϱ���׹n`�}���Y��E�e������kրf�z�)c��c��H_v�|�Y����;�⫝A��2Ќbu	8��
�w[7�)�^�3���Eq>���x'j6U�c�X��sr�󸹕��)}j����MW� ��x��|�l��=�&���d@1��=Uk���McAr��|�C��#���Lb��Ǌ�փz��ų���^����/ݍ�p{�^��\=�9՝��n�ܴ��X��H�ٳ�.v�\�2����(Fߕ���	�P��N�olhr}JY�܂�c.�MiW�y[j�𨡅%7������y���c��;O�����XZ�v<���g�e���r۾��,a�%���^'5���VQ�YJ�9.�ɠ����[�t��v����۸�e௮=!S컈zL��FA��螯�Fi�b��S�n���w����o�63}�do���JȻP��K�,��C>�qE�f�o#ED���gA�6�
{m�WW�R��=��ӜƼ�N���lz䌉VI���gq[ǘ� Ld#��A�'����g<�X�Pu�)���	���<mjI���#�;���9����۹Y0�,�M4v�w���Iz�=��/Z�Ѝ��m�o���ў���mD�I˖L�}x�`��>��;v��x�F/�q�9�F�]tc{��ml���|��Z��R�������E�9��5DtJP/�;�*�b5I���Ѹ��5Ԥp���*�vA�m��7<O>1q��_�d�ZI�D�"�@D���d��{j�m���j�wu�#����H�3�</%�5��xF�����zi[��g�����j���D?B�,���L�	�����7��D�5>��d�F�є�HۜV4ʝ�5CSvO+���JyT���ǎDn>(������2��:��Bn�,��<B��s�s3v��rm�WAh��w
���<���w	�K����3�|79�஦�H}�e�m�\{�{�ݜ>�):���f�c(p/ݴ�l{�p�|�sä�N��Q�c�-n����9қ���6%y,����J��~.�y�u|�Ġ���3��Z1Nq�;�4kTx��pT�4^����H�d��.uQ28�v�s���b[Y�ׄ@�6,6P8ʐ�c�Kl��"�^�;���NCx�B^Ni��l�k�ڂ�T�mj-{Gƙ�)/ynx����٪�/BL�3��}������\ބj��Co-���DL��+j���}����N̳�v�F[�@&�w!j��wk��*�(�q�[7���Dƚ��X�G�*�*g^ŧ��S�MiwL���tky՝���ӈVa�B�K�z9���*,��_�z�V=̃�b:P��$t�R3]��Bk2��w5����'%ɓ*r
깍A���1}�6�R�rT.2p��L �I����3�R=��[SS���Y�5����}z���}6!zO�WD2T^���,y�w�h�q 3W� 6�K*Ul��H�Nw���c$�K�,tG>ڮ�#�n{�WOE�1ߪ���m���P��W�_���R�yت�W��L��P%�N\��6��V4�������BZ�z%o��5a�R0�H1��W��)g��q�]u��g���.��JW��O"�g\aT�F$�$�g*
�e�@��(�>�Fi)��G�%��b0Y�e_e6�@�C���?i���*���HO�%1�<	��y:��U}fǺq죈��K���I�NOM�e�m%u�$X�����cc'�3�U��i�d�Dj�{�FFe��d7N���䢃b�k*/`.��Vꬎ�<��,�U�N���Hj��S�A쩾�@X�;�߉J��aNE�ZΣoR�ʙ� ���w�U�ɹ��V�� &�0�o_e���o,$��b�ѵّMg���Ƌ]��kn��O���{\ė���JXU�-�<ɖ��
�P�+��)�"�ڨx��d�3�89>�I>OM�sq�x��2|h�m{i���� ��Y��+c,GcTTf�X���4!�:jT�|�&�酣g�i!�];����3XT˃g-�������4�Ҫ��a��;������ڇ��8G�kL�6�y��:]�
.�������o�n�KI�L�=ȟs����·Sý�9Koy7-�J�J
��I��j��X$����{�5�*��)�]S�A�A lg�9�L[=���m�F).��ەy�u�LIh�(�[��J����E�SE���h��`�X;Vd�d���ZT1"�C�kڛ��[|�$u!�؊K
�Ǣ��.7�.�W�<�H���٩��?�s}��۹JRݓ��d|���@��5�C�X�	�� ^��ǫN~r�)�I�N�}���N�F�|kʳ٫½��W�2�2_��i���{����T�jFs��U�v֪Z��"�]������3��ܜ���j	�Iڸ��P����5�vG��[��l��CR�M7i�
��؞���>��7]rˍm����d�۽j��mn��aq�nWu���ٱ�u5���ֻ�\��ƶ�L���]Į+f�%��4N��c&uedL���-���>�T%��"<V["�4bd�L�z���i8����f���M*��bǮU�'��&���t9�X�3Z�ӫ#t��;��{3x��}�=���ko�&+8��M5]���o�E� <�x {|����(.����ξi�b{�P���V}���W�K���%%�j���.��]i��D<��s���U��of����{��3���	�Q�^+�$��Qs�n�1��j]�{[Y6�4�>���|�rB��؅��o�����c�7i�/uV�.�ޯ
����%^&���z��)5,s�+�nT9�dc ��G���&��L��i���u��Yw��zi c��=�ڶӘ�w��*�q�e��ҙ8S5��Tq)��{ű
j'��w\�o���x��Z^�No.��Wf��B�J��R����2�Dqr��5s�b>޵�V��?N�/Cу�B�r�`m;r`|U#��5��4�6�ʧe�k�l�>hg�P\�*ܝ�9£Fި7����z�ͼ�@�l�Q.1}�@�2��\���-`�9��;D��{�sޞ^�CK�ꀭ���)r�Ǖ�E0�b�\�+ʱ>X�b�s:T���h�p����g�=*<���yZ���͹�aq��Az�<�[/�&�_L0��[{F�s���H�]�(Eo��N��ѣ�fJe�]vV����3�E�umdҞ�#
i���[�ypG˜9f�R0��u�|,��h�.�N���si�'�G�V����~�=+x�,�A�I�5g9�g�����ׂ��7C��eEwo���+�~V��܅���}ǈ��X&��p;���G�3���sA �����H��0���T+�"�M۲<���mi$N���	*-�R�rP��@��&_�U��؈��+8��:���gE��ߙ��`t!���ۂ��rCn'�%Iz���R6��z����_Z{^�
����W�j*�okh��������S�z���H�����n���m����+>����&�/�<s89^w&f��[�1��|"�.�6.�=�+�O�pb�a���i'ˬ��(�ʣ��)2_׶���8{EmНN�	k=Ea�O�=A�e�s�豫1jo��s-��W7�&F�B������V�Y��f��%?S2D=\B�X�o�j�z�[ߓ�es
�:j����<���ȭ|�K�X�I�m�n�n븋�x�O¯�c���t�'8�}J-���.]�y	2V���RF���s.�����g�ʹ87��g�\i��{��1��y򵀞q[��5 �Hc�6U�F�TI��E��h���ǛN�U�Ut��2d�����Y`K�kyr{mZ���X��^m_˂7���P�f�om�|��:��O4�|1iݦ��V���Q�#�ó�q��)�M;�`n!��5~����#�y�ݏ��,fݘ0�%�4���u����:]f��!���w^�k�@�yxDi�w���/z�{zÁ&|�Y�N����`L�����kY"eo�5.� �qS��b�M�żu�ؙ$�u+]�������e�$�*���WE�rM�雾��fmj�k��{@�:wIS;�!�& iM�w���1��)xP�P�;F�a�5g~�,����&���k����m]>�QV�b����gc"�munjzr�f���^�`���(��'7ҫ.�v�2���NmV�7�Ū��fE��.R)�Y�	{��wo$�����6nE݅��}�}��[�nentlLz����_U���a�F���f�����1dv�b�D������@�a�Tάy;&m�U" w8��7�[G�x:�;�1�<q�ǂ�|y���}��=���s��i��T׼�u.ɕn�>vy�eZ���v�_�k�;���s�$�"���ɤ��,�Ƞ��"�,*�1�*f*�3��¦�3	�"�2�b�'3��j���&2)ɩ����Y�Y�9e��9�Uf`Q�aF��4ASQ�8Q��LQUD�eD��D�a�9d�ME50ED���V:�r�"*!�̳�)��5�5j�*���Ɍ�&��j��0�3�r�(�
h���2"r0���ՖY��	�� �b���
"+,���+0ʦ�+2&��)�՚��b�R���*s0H+"k00"��"�b��ʪ�2�2u9&�Ʀ��,�iɊfը5��hɣ3!��"̋�Iu��E-Ud�RA2Q5TVa���u�Z-��ն���s��r�\(�k�yv/M��T.����m�VhC�
xwd�������٣����5��LĶ�*�`���*�9��9R MU)��\�r
�;���^{@V�����p����qp�K����w�:���Qw�d�m�%�sQ���جo�xL�MV�%��ɾ��݋���ٰܸӸ�E�[=0ڦ#[ؠ�����0�ʯ/��޴�L�0�w]k�UK&������܃7����.�.��a�Q�S�r;JCV��vj�YL��yl�����r�^1�2��Fv�Ǩ/����e��W:(�BJ�
հmd�Ӌiý�8��k��x����/ɻ=~S�;��uo"��.ꚠG@IS2�v͎��0R����Bk.�q��^F�k�Tڢ��|ӣ����1�V^��k	"�(�)���(��rz����T�|&Jx���D9�H��N�BV�+��,�8qi�E�A����v�}أ�j	l��r���)�At@͔�37͵�+?-���!K�y�MXW�޿>�N��������r�����8͠eX�2n%=ڃp�i&�u	2�0D���p�#�������@�c�s5-�+cO��M�[nr񼘓O˼%[����|A�M��t��h�kx���އ�P,��^D��'աj��ݨ���;���^�E*fvx��������4��>��ˎ�W(�.���V��q�7ׯOaOJo�%J�{�0���e�]��=��vda�z�Ծ��y۷t&��S�in����r띢_�='�z`��x���aD�b�^�y��(.s;Z��ʖl����Ok5K��臨��,D�b`�z���*P�/�/�������xui����sr>����j����N�$ꚫs��Qux�Q���]Q"�w)T(���Nc���n���=u��4������$q���Dƚ��X�H�%C��M�{�|i��ݣ��N:�-E��/b�>�~�2�g��[J�s����!�P�(i�����& ��jS�q�n�,���;�-O���cC]�
�>~��rU���gDnK���Z�sb���iuT��h ��X7��������?J{^4>�3�Ŋ��f�uP�!�z��g=�vVm�%d���D��'r�m�ُiƍ�@�uc$���g�:X�ml�Xn��3�ƴ)���W��]�&4�wg�\>z��v*��W�W�VncJO!�n����~x#L���h�] �@�6q�P[k
�Vu�}ʯ+��ɧ4��j��2AwOO��O	Qq�C�����o�q��QJ�����t�eʁ��@�ΰ	x�5]gj�RP��_K�s��-��˩����)GT����Y�`!�=W�$T%�עVW�j��#��9Q9��U��ﭓ��r�H5ݡCZA�1c���ֳ5��5�&hl`�ƨ��AWk��&�,�*�K� ����&d���e��|�̀o�aći�i��:��=���2B�	W���&�C������������ݗ�ivM�̉9;.�5#�+���PW\o�nb��2r\�~Lu�ݻ��A)]���~�;�}#�y����۟v�)󲏋�i�"RW��s�,�V����X�SI�V����Kzk�Y{ֲ��y�*����[��Cu���Fmx���-��ׅ.�P��E;r����u+<�r��EaA�F��\��|�&�酣g�iUӰ�@�;}�����v���D)�2[�y��\ˏV+�����6�ܽ�u9SO9��tP���brK-*:��3����w/�a�C��2ޑ1�9	�H�3��*;<�p�eX���;( ]E�*2�r��w��ب�1TkvkX$\�DJ���M��61*vy�m�����~���/��t:�-�kx{[ء�]�?U�\��3�����T�z,��g�S<���Ƃl��l�;�[8���'N��<�[�p��e�c{��|a��p{v��*�����Ϩ$i`�$��ۘ�uG��Ζ�ֺ, K�p��y�J)GF ��u}��u��3��_a�eY��pk������X��l'�\}�=��˟��KUZ�>�\�{�ĥ�Q$��-�&���9�8���E��ݖ��.`�u�I��7�q��N�#Okd�|+���p2d�*$0)�aY�
ݯ�����=��?v�e�jN�OQ�N��!��K�Vm�D�!�?
qY�����X��xQ��x����K�@}y�U���8�P/���3��kX3\΁�
�?�m*�u�������RE=�(���f�W���{Rd��q[fl�X����yĸ�َ����N��/��0濾j��R=���E����oB$��f�+���	M~6��)�j�.���ch���O��3��^r�H��fVǧZ��.�&��5�d��Bo�����r��yP�]$�D���̽�$1�e���s�l�#��G�/鲼B���ڡ3Ԛ�V؋�[��@3��]+u�G��K���n����=�.K��^���T��v'1�M֋���n��.�ޢPg{7wg��PZ{���w��~��=W|����ɟ�A���7��u4�$��<����MѼ��$��1�{�(�ړW\���6Ӓ������{}�d=yK�����rpj$WU��y;��3�w+�V�`Y����w͵�G��)��u˸�le�]ǩ���z�)e;��f���6f��g�����i��hf�B�5X��o����L�̼�Y���4۴t��,������]Ǯ��=��
i�}�áR��7]fM�NZ�ֻnBk
���?J��q�f�wJ�ǅbu3^�\��.R�j���\_�y&&��ں^mn�Ԏ�x�P�)ɋ�N�cm٬C(V�X(Tbusx�`�ɸ�Ӑ�&vNÃ����U��Ng���^���%(uW17�>��&���<�q��-���zc�����{�cf�#����̠��]��G�E�zL�'؜�o��ؖ����qy�[뗼��\w�A��,�X!����-o���>˸���(�z2��Dq���uͼ����^����ш��� ���A��*��Y`*W�.��m�b-�(F��8�x��im���@�nu�e☮��m]���b1X7�p����������5^p�Kitt���$ d4{̛���A�y�V��,9�����:%LL�$r��c|{I2���1��_]E�5,��1&��K:@F��n_
��>,l0�<��N�� ��Z����}4-���j`�n0��Wg|2�x{gnW��5�IM��OZA�*��O�nl����l�W�}g+���]���'6Δ�$.�����ey�_EKj��|tr�S�g�٬�F�n���v��ɻ�3t�,j�9sS�Xj�"��T��O��(�:��'G/���`<��[�3k���^A����%�U-�~3+��\�;2l��͉�M����hE^-�1ny���w��y���`��{{����<oG�P]g��)�O��V%�j�U��tl�6N�@ �Y{m%ܬI��6`��FE�mǶ����͢y�D��u/��nk �^�l�1{R{�|�\��+��	nft����u��Ƶ]+m��8=�H����Cg躃Q�w���nw^ۓ�߼��\Ͻi^6>oB�tt���n���s����û��A���8������*��z�i�'T�[.�Et]^0a�tlW	J!܃�'�͡ۂ�qS�ˬ��!f��
���8��ܭ�24�6�+>IW)P�:�-:�Ǐm�d|���ٔ�,0:'܉�OI����71�G�0�,��_�z�W�d���(,��v�-��S.���F�+�ְgE�v=LZKE����}���|C� -������x]�w�m��/��bO��z*=��$k��s���T�<�D�}���7v:ݮ$n���_�by�d~ݖ�F���������?D����奔lR���mA(g�k8�����3�:��b<���/:��ƃ�w2K�y�:��@�յ5xP^3o�g�OkƂ�ئ`bl|]����[#�_��	��7w^�d��6N��l;�[5��D�s��]i����h8 ��Gl��-5W����U��r��x.�����Oo�:�7UZ��EY��f'������z�ޛ�w�Ҷ�/y(�%cv*�Q�D�>�����l$�T�Ο;z������Q{���q4�*�~�)�xg{I�)1���*
���(��"�td{c]7rF��u�=m؞n9�_��h�Y�9�Har{u��d���S����$>��y�{���Qu��鳳ku��+��QB΂%%t2�E��}��V62r\�~A����hR+��b��4ҙ}�od�V�_��h"���u�Bm����{]t�+��{w�$ֳxv���3��40)�U9X����:�A��x��2�T���5��8A�_yp&_ҵf�F��\$4Ȼ�_ֈh9��]�e�mM�.s�WQ��+N�o+>�߬�|�-1M��y�� IV,�X��K
�d"#'��F=K�R����-�O��r��o�ؼ��TS|�a!�1*4��v��E֮��1����;����]}B�}{9Z�ҥ��Ʊ��˞���m酣g�i!�];�� o��Xr�~�M��ڛ�6[���FK�k�S����da���N�����B{��`����8|E��x�&��Sc~S�-q��+��v��LhR�x��w>
�F��Y;�7�`���6���\�kp�k�� �u&�w�vkXȊ���z�ʚ�f*k֊@�A�sҘ�=V;�Nd��CPp�K�ҵm�nK�J��)�U�(���W���ފc.ʑ�͵LW�(� 鈴�ݓ��(���gMR�nt�l�U��ĥ��D�:����"�`�����>�v<��U�	�Z$�u�_�;<`Q�,��-U��oe�^��"TT.L��ԇb4"y�fzP�y�bhg�ͻ��҃�~$�A�c+�T�m)j�m��8��G�N+2�2X�t�����fu�v�q��ۻ=�HF���WX�':�VD���Bm*Ď� ���\kX�T��R��y["��<nG������v!�Yt��>��xf����N��	}����Ce�i������wnX#%r�p���F�[�&��E_+|��[��K�o�k��)��5�Ӧ�_=Mΰ�c�vOw��2.땋��kRԹ��k�\��VcM��[b��kL�y\�:y3�;�iv��А.<]qa�^��N�css�9;�a賥MR����.�9D����w�����vq�WΘ�ARᲩ�̘�#�?,���V��������M�n�,Ny�a���������Ud��q��m-;\K�t}}���9������{���ƫi��s��&��
��^-���u�g��;����q4vgNe94�&fqI	8�u�ܛL�y�7�ìp:��J�9���F4�D��!]�����:+������fk��R:�*d�a���j1�J�r\ܾ�>y6�wgN�r�3���z���x��):N4��۾A��[^d��	�>��PȨk}˽]�o�g�+�U�Hߧ����̮ҙ^��Y���pLt�`�f���+5�e�KI�6��X˘\�/e��/R�Z�U���֨�M���K�i���S��7>Ќc�o��
���
�N�u-�]�1yu�0��|몐.4�P����k�9xl
���
Js|H�8ߐ]lu|͚��y���n���Y��X�f���=����B�PU�.�{��q(�zL���^'5_cUZ�ޞS.�<n� n��q��X.�k��-p��kS�e)�U�(֥e�mVW�}�r�vƆ��틮�ՙ�s>��]*����(>��zC�c]�yR6{B�ȴ�k�-���:Y�׉"�n&�e�Ahw���>���y�$8�5>IY�h��A}nUA]q�~���fB/\zB��.�L��FA�K��6׎fͽ���]����X�*R�d�Lb%�L�8�(���Rg|Y�#mO"v����ȧOJ�]Њ�`'�*%
�s��/4_L�6���^3��`\c���]��[/�����C�b�����1�9(�0{��^J��t���b�S�e�^@�@X�bn�Z��ޔ�NYݜI1x��������q2��N����EE� �떪0zaEYxv�+�W��Y��N��#��SZxk��*F�d���,�=:���'G,D^��{3�jSJ�^�s|�J���T�mU˸�0����T9TN�D�N�>nS0����ێ�CwKڗ�'��{�၄��q�{N]{j�\ߑ1��M����ic�ɿJ{�SJֺ:���A�>\���Z]BL�B� �˽A�{Jd�|�9�D��wR�w�b�̈́[.��I�]O9a�}K�4�Z�W�+���۝��~��h��:˯>׿gTA\�tW�J
�+�qWTA_�
��W�h* ��AQ�"�
��
�+��W����AQqD������ED�"* ��Q���+�DTA_�D�D���
�2��a۟@�>�������>�������UUP���UP�w:k6��[lD��B��r�I�5Q�UT�ۛ�u�kl���kl�(���È��cf�l�[m�l�7rٍ��V��@�P�8h� 4  �@�l��.��U���l���6��ĭ���ش�T���Y�kZQfN�l�ڊ��,B�Tmf�F�	ݦ6Ƭ���k+ZVP�n��l͙���j�)*�����[Ɗ�[k4�    O5JR��A�G�2bhd4���$�I@M`	�da0i�2ѓ �`A��2`�S�A)T�I�L   L �101��&$Ԁ)L# 4SѤ�Sjz��O�d�����{���ׇΊC=@������G�I IY��($�� ��$������HB�F�����?�4��$��\��$����BHm$�!h2E	�BHeo�>��|b\g���RB�@�4U�R�����I�Y���2�PQB/~><ύ�+o,a�*���,�Ɗ{Y��1�.��1��Ch�@uXmni���X�y+^Օ)mh�314��D����RT��Y2��* �T(�\�"L�#n��
i��C3���SXn�x�#Eɖ��e�4+#�K)m,@����rTZBV�U�WC��R��
^WlC�Omn$�l��4]�X�d<��������n;�;Q�B0���	.�iO3��F�V�Ѩ:I��p�0�:܊�9�v��/�Ѓ�jQ�i�6��@�
���:���[�VՋ�Ec�N�Lv�虭b�w(�r���m�YL�G/[�����%����ة �����ay$��&�+��V":\��cuul�Y!�j7b'��m�%�8`�B�2��:�6'�,�Z�KdYB㻲en�V�P-eZ��u�+Cr�T����ئ���DB #�֝X^4@R�31$Е`���0>�@y�2�
N�-��S*]-L)S�cOi��l�X�5�i���"E��Q�t���l�TI���ekC�&��*�ۻ`�#.U�y�.���;��8ۙQw��n3V��:�{���Z�ّL�H%�jɴ7]e��VG�����Sto.�BV�6"j�����Ś�Ѵe�1�nIxn�O^��n��[��7�x3&4��`,v��t��Ԡ�8ضE����"�McM2��W�X\J����Kq��1^lf�7:q�����_2��RV�Ì�x����Ԑ�s)ՋU�,�y.;{j¦�F�4㈫xs^P�+�~f�5:���16)�㭒�l5��.�OH���B���6%���aik7oKv�閊f��*[�j5�]�FȬ�ӓ$@À}�Li�kn�yzZ�;-`u-;������E-��%�CJì֨����qn�����շ[�+�e�\*A6$�ǔ�۔;��MWoz�PGQc�,:u��@M��V�J�)<N�f4�p�F���`t��:S���t�3� ��ÛR�R�v ��@XW�� ѬU��ʋ�_k0[@���1�w�vjAV���eA0bF�ɰ]���-���� ��v�$&��(��6������>M�mnl��Z����̊V�1P��I�r�dj�Sw6����+��n�b&Bq�z�C�C��VM���Xj�`Si��be����[�H5L���Y1=���\��)���/d�슗h^�А�V,��5�<݋����K�RKY��J���f�C.%kv��軘L�e�ܿ� mJ��v �f�.�ݡw��7�[1e)5���&���D�+`�r��Գ)IC+t��~��_�z�s��}��ȑ=g�� oTz(1��=&�����_�ɚ̾Cvnt�wJc����ʸ;���b�:u��7����L�l�*���O���B��k6e�,������TX4zW�>uci>�n��c9�^G�#tT�s5�ַFv%��t�P�i���8�g= �e%�����۔��,�5Թ��[��\�U��� r-��ԃ�ԉ�+��kn�������Rf�I�A�^���кѺ��(v7��w�կ�����i�*Nz�/�+�F��ݬ�%Tѵ���
�`vt�}���,�cx�"(��L�S#R�1Na^�O�e�j����������oQ��fY�W�irJ"c�o���F����;U�]*3�1�G&؀�Ӷ�
�
��Eq�DLh�����e�>�����x�JL|��`f�q�$���R�	���eZ�w`;�A���.��d�a�0�o%7@�v�]\y�v]����4sZ�fk����.W&�����%�o��9��-_�+o2J�Ц�p�49�j��i[nR��|A������G���Ay|��b"
�2�:%J������D>+U�'M�5�3{�×k��V۷�(��"�Y��}+09m��q\r�D_[�9�{U�9��d	��M�c�M�A�1gf�M�ӽ��!k�G�Y�����x��z�����A8|��v'�\Ku��^��p���uh�nu	��\�rd.���7�}�BZ9�ۼO�;�*ͲHR�n�w�{;l�EW&�s����y�X���w�����]�c�E��E�0�X��1�7��vF����'T��K����.�J�ln��x\:��$���]�J4d���
��X��}M1h��kB���z���vQ�3��{xޫ�Xc�<�m�aθ$Ѧ�u�����յ>Z��X���1%��j��곹�7W8�+�yYW�^G,�+E�	��^�l
�`snh�M��I2�k;���sʻ0�J�	���}B-1�ܟ3�"�y�{RvJ{1Jdc���"]:6T��s�OVP��<����ls��+��1�a�X�@d�{ܻ��O'��`�t+&8�nQ	Ʋ2�4�&��_0w��n�vI��٦c\�r7�w� ��f��8��98hӚ�Lo�X;��y�6�V��/Q_{�hX7zh��
aV!͞�9��]��Nh�Y%�Pm�q��3�Cl$sݡfY����01WSR�\ھ���v�����5�ȧr�����&Yc��)d{ҹ>���YB��a+:�Ճ�5F��F���[kti{��m�F��T�����y��"Q.knz��aj���}>����a�����BHCːNb��I$<gv	�&Ϥ8X��$?�������P@�8�!;�ٙF�a��a��1����tX7_��m����`�G�*f���ݹ�v��`P��=��"�}�ӡ+c��NS����v�t����n�9%�n��׽9s����d�ɰ���X��C(b�w�X˷�F:5'�����YN��Th�Y{��7q^KjS��p$,�[ZL&a�R&9�	�n��[۫��A�P>[����x_vQS�*ZsX:n�[���t@V�*�V�9A�q뭥��^�7=���r���Z#vk/�ۤް��a�Y��ڷ,�uj�����6Mw�Ÿ��90�&v���]6�7wO�����j���)�ТC��K�T�^e,�3 %#l$�����2��x%M�2�V�����o7VWQ	�uB��HW]�y}�>z@�K/X؟Qn�)�/M��-�W�o7J�>K5�@a��Q<���,���ԥ�qʲ��Ʋ�V~�X���e��q�(+x��I_�._f��i�:o˒�W�!�Z�NX�t
2�ݪ]�m�&�n)��+MJ�6���;�Vт=���{kjS��&?�+�u�o���)�"9Tܭz��c~��GX�8�D���s(��4�4�.L�#(XQ�YM��9I���2�ok:�l�A4���E�Go�<
�Y �+�%��>����ɕ��v�;sY�0���Z�>\Z�M� |��E��[]�ę�Ub��@L��������UA�K�6^���B����S�4� !���y��f��,��Θ�뫗q3�+��&**����������M;��{����]u��\d��9��ie��j�:��c ��I��J�Y����X���/1oV%$�(�L|,��7���#����|�w��iA��oBح�o1���*�ѮJ�/9��J.����D�6	A�<�e�H�о��^�b��wP�\�U.V��HM��oj�$�l����κښ�.��,���j�en�T�2�L�Ʀ#���Ӎ+j�G����6����O�?;�}����qH�pL�p������ȝ�r��a��._X 3��0�c3*�)U��7sZ��C�r����K.����}ڠ�o4*rd
�S(�k�B@6�C���#�d��1�ӇiQ�T��2X@ٹ��W5vF<��f<sFbD��]Q�<�ۭ��I�q���ja�� �<q��� U�T�$�/$���
B�}!v�k�rJLpE�ֲ��ʂ����$���eX!�t��6�^
:���F�֌ `/�8/��6�-���m��6�q[��y$�
ȿ���X�<�A�n�EN�&�|[�ݮ˷�a3��v�	�u`�k�w�� ��#ST���	�ͮ�{��Y���w;�u��OH�v��1����oBw9<�;���y�oL��Y͞O���ɥƦb�!%kk���]Yr��(���PX�EE��TcX�*�QTE""�"�U�R,Y�AH�X`((,�A@U�$P�"f3���3Į��Uڿ9�!1��������P5�h��|O�iu�ߝV`���OG��y/�w/�[��:I����.�vnQ�Rc��q7��=Ż����?���oF�߲��E��Ȳ��blK��22�Lz���q��ʿg�h3�?��דE���(���-��ܩ�����;|���-#���r�;�i%����u]�]���~�
�3gm/iV���Ǔ��i��b���{�a=�e�;ִ�����[XP����� 4R�o+G�)_'��y��Al5{z�������0��N�1���eO2�%���EB Ǳ�.���9���6���w�������F�F�lP�׈]T<��L�V�(=�F�VQ0g����ZOy�����oC�O���Bo�^�z�����$y�k�ޮ��o�b��Bټm�M�r�i� К�������{�&Y���@�mχ��2��s��.�D6;`��=�<��zj�ʿdK�����kyz�ݠ)��J��^=��q�vz�t��ɻ����}P!�&���R����:�J1�c�=�|���ud�����j��;tQk[�-uq^6?j�y�].����c"�_�O�������!�i[�y�J�������W�cX2Un��g��ʪ$!�t{���~Y���������x�0y��#�\�����^K"����ϡ�dx�.w��f1n�6��c���dO�y{��[:j��	ypI��G�[��C���(����~��}P���T��.۝��i?K��xU�f�!{$ô���,��\M̽����5���'b�z'��~�zOA�	����ޫ!�Ko-�@L@Uވ��3ޭ^��>�S	��㙺}5��\��:=������^�c�l�����^N�����"b��U��j�c��Ʌ�)�>��{��2_�,�~��oy��}�H��n�����j��w�_�o��n�߹��%"�1g;Sy�){�?^�-�����@27�l'�4�8��AqZ+�=�����|�����3����j�?��0���Օ���Nì��/sHn��աǣ�'��CO{�|oṰ̀���_mY�E�}z�V�+�%��%2��SJui�6K�Q���!Ss���8sͩ�R�l$�k0?���M<�UXy�L��R>	>o�)�uմ{�g|gVʹuv땩Ӱ��?~e.��4z�x[,����t��q���m�Ρz�4��;4�Ro_u
i=�{Z��[��J��}dF�tW���w������UL��,�}}6&�ݒ8�<�On���v�Z���JW:H����ᩮ}�o2�����-"�A}��u�TPL !�d �"���"ȰX�`�RDdDP
bȲ)h��|��<�oZ�����������*����q߯��%
f��F��Vd~fmn:�r�Dt��~�4����fF6�e�Mn{��[�z�L�o���+U�kP���*�M�ǩ��ʈM���x����:�ƒ@�ʗu��k�Q痷A��t�0}��(b���o�r�9��<�{<�%X�g��//��G������ws�{��V��3��ܻ�[���yx�՗!s�N�����6`����VU~��v��q~.�p�[ei��U��E��Quͨȉ�=���l�kv�sR��o�Ecu�nB��,�Y�-ͺ��^�MrG���ߢ�~V��t�/@��W��j��O?m4َ�0����U�j�����t6d]��-n�,�E0\�Bvp�i��,,��P����&�{��s��,�/B�ٲ��xY�l?g�L��u���Qq��ӫ3³#\Ç���yۮqF�Iɋ��z_�N��x}c�g�g��������F�E�h/N4׌�"\s�8��Ol9V(��s���_�Y����l^���Ɇ��zl^�	�ȇ��$��f����"8����J>�۩5Y����[���4�x�� �%��Ä�p� ��n�{;%�>��;�ּU���pv�ӈ)�W�(9r��Jro�i FU�Ւ56��.���y�WkwgG�	
ƶ�*�֦Ά�Y�n��K��H5Xm�Ą�R���cz+(Y*��hM�wo��??O�I�왜��:;`������Ѕ}��G�j/��Y��S)��b�o<;&�b�+��9	ٞ��=�(p@��Bk`6��m�Y���5uo�}N}��W��B:��5W�}z�`10qu~WR��[ q%ۮ��v!F�z�>�]�%��K�P��t�g���K%]Q}��z����V���5�n^s�]��'�Ʀ�{T�W�P����5�a�y<��9>�P�����-ʝ���l�RbXR;��+��S�����wq�u�a�+�ed�W�0�hy�y�5@�C������ߥ�������Z�u4M�1��C^0Vת5n]nI�'Xֱ^���-��m���s'r���,ˮrQu�(��{�Vp����e�­c�T�*���WL�����Ⱥ�so��]��t�-��Q���Q㲩$;Nؘ�g��4�V�wvh 5u�w%W�=����6����p;|�7�d���v��R`6'4�A�l��;Yw��Q
ӽʭv��S���tn�+��91�GgJ��g�K[OM+`��1BLڌ>��S��S-�2��g&*��_{�3m��<��ryY((#PE��1dQUF*�EX,1E�1b
�*�#b�`�dUDDUUF"bb"bb&~������=�H�y�d�\�������Z���<���=���T�{�\��˞�hp_����lK����k�cnq��f�� ��e=��/Aܶ��������R9�^�4��u���������o�׮���h����Z^���)��d��C�1on��F�ט&c�$�p��e������d�W'��r��x[��ZQ0RԶ�^�͒�yvoN�O��:-�8���g�Ɠ*�`��n�P��!=��˟��x��e��GO����/�aU�oV���U�����e���T�}=Z̘/��/)���,��20�^�Iʮ�� !qUw^�]�JyX���ܯ<���5��7���j�)-�-#�J�_���ҽU���b�|@��tA�Ob<��ys��<wD �����[ab-	)�K{T�[�h�ռ灭��U���f̾o�����8a��|�=ٗ�c�0U���?��[��^�3��g��\ޜ�7 ��ɩ����w���G�ٞ�k}d����'��{��,���ฏ�%8:�bt��ъU�]^D������4���?ukq�o�{���aqZT>��2�����L�ZTK�e�c>�h��K��kC�S=�����g{��y�,�/�/�2�2Z����0�L��#דt�b���U�y�m�?)1 T։�m�Գ6���幋�ݪL�`�isu�oxަ�G�,��N ���!�u,���-&��u�V&�%r�2�iūi:��kV%�Y�u�E��x�l��c�C)��JDI\�kX�YÓTU�S"�&m��&����f��9N,/�Y��w{����2_�ws���`��Ȫ���u1>xͰ9��ֲE�0�{F޹N��ms�̆Y�w��(�9|Z�Ӿ`�(g�,�Z��}fS6��%�ַ��	��V��ԚgoQt����p��]8�ᛯ�Yfq��d�\�1����m�PQ��(:_6���M�Ng%ԥ<�*�J����C��D0�8��8��e�3, �ع|�T�m���2�\���6Ø��Sid�y��Lj�r�f��Z��^�w�2����m��j�0�%f��nkw
I4:e�2�ų�&:�M����̦P���QNU��]Pۡ6˧��
,����K=}�+d�U��"���k\�8^�,�6�Q��N��.ӈu,�I]�����P- �j�jݶ��^n�:�����'Y���e��])�f\�ŝػe&��K!��f�,]��ۆi������P6�^3(���l���j�u�[��z�M�ӆ@R�1�V�w|��2e�SqqA�7��q��q�r0;�՟	����]w�����@e#��+h�`�5�e�����WE��w���|Z�+��4qZI�W[��.�B���g �.�úl�1>�"V���$���.u36��ih*��!��p��md�?��m�N̗���m%�yf�-/���+����k!l�%t�3��4Y-5IԲJ��1��C��c��]j
��&K���#������x�Lܞ2ȱ���\�P�+Ó	���q��=���ҷ�nIw�sC�[���gY�9]9�b�
�E��1c)�
�`⊥�E))X�K�� ���o������يN]��y��f}.];��_����u�ilT�[TA�j��N2�Y�_�u2ΰ���zY�l�B�m�X�\���&R�#�!d�/�Y�%'l0�f�3���\�l��)�m�i~<��e'q�z����,��kT��c�,�M�j���[����s:�*��3����k-
@LL�>���LG�);�[iv�!LNL��u:��Y&R(r۶л5z�z�TB�w���-��.˥��.٦i�lsol�Afل3�4��q��rV��N�0P�I��X����x��Ri3(]��o85j�f�Iv��:�Z����&�T�s�[�hP�M�������։���dg��\�/��ifS
Nޤӌ�b�ȳ�,Ʉ�o��'[!�K	4�g7�q���HE�ձ���lf����]�����n���+N��!I2��H) ���q��W!d��PR) ���Z`r�Af)�ƐS�RA`l�Y ��
H) �wǏ<fi"�R
AH)��RAd�RAAH�P) ��%$aI�'R� �e$R1�{��H) �2�AH)"�R
AH,4
AL'Y ��aHu%2u��Y�J����H,�%$���@����R
AH) ��Ad�),�I
��I��<s>9�/�V��|�-�\�櫘��S<��D0sg�������1��EI�R
u�
AH(bRAH) ���R
AHf��فL��Vu��&|�a�A`*�R
m�
��Y ���R
AK RAH) ��) ��g�����i ��فI[�� �`RAB�DR'I ���R
AH,4�k[��$���I.�Y �I.�d��Z�����H,�e$O6RAH,�e$���RAH)B�.�I�RA@�RAH.u���
H) ��*�)�v�
A`xi ���R
AN�RAaV�Y �c�ƳnjY ���,�Y�JH))�
AH) ��R
AH) ���o���D�Ad�jY �-�� ��′Aak�,�P,��RRAH(u%2씐Y�JH(JH)�[{���AH)&P����I ��) ����Y,�H,��/�col������Ŗ��ҟ���m�='wL{ku/�1�4�0?�}�D��G鏦~��.o�m��mm���0�Y���s�N;�K$�q�5\CM�ԡ��e��_t��N;M0�E�x�!��2˦.�{U͌�6ٙe�F���j���[2e��Ыє�������.�GI/��5iL�m���6�����k���i}���I1?n\���<N�.l�#C�$��Z�L�.�1K�i��<vύw�5������K�X��5� ��(�T͵|����'R`��W�E����9��v���v�0X^�����o\&�A7��V�i�*ݴ�ǩ����4�f��gXk����q�]�&�½}n�P�V���>�A*C��U�n����� ����菧/+���ߦ��+]�c4֬S3�	^(�]��Ti8��K����계�%&�m�5�n�/v�T��q&���8β�8�*��w�ݹ�gP��"�I�_[�
B�Y�HZ״�(�i�Y�r�2�N��8UZ64Sg�}�=�'��r�Vi��@]UԹ�ӵBb��|h��#��"v��}�Q���4U�m8�&:�Kn����X���Goi��yW�,i��) ��i�o��5j�c�K"�aV�{]�9�%�F�G+x�TІ*�!�@�/{�XY��e��K�f�b�C��g����.�I��O7�o�T2Ρ���ժ�K���5!���GT;Q竖9���������ٿ���
M W<_��xgYd�u8�i9Te��ߘ�b�3l�S0��*�bK��g������&PX���nQ�r۫Za�e�R���Y�xv�Ci�5���[��
�9s����׈�|���I�J�M��rr�_uf�49�|� �D}G���V\����>���$&���/ϸ>�N�uǘ%ޗ��?ݮ��m��T�x.��U����5�#L5^y~��VioMu�2���P��������H嵴���4�l���Y�2��O��Gʆ
��|˱�ꮳ�"F��cVl�:�wK�i�r��i�*�l�T0U��m,rˇ��G ai����NۙƦ�<r�cYµȂ�n��$2kNk�Ε��:���>J+v�������p&2#��+���40��;��(��Í�U����R�ń�x>=|�����r`�Qv�8�o+
��*��/�#�����S����ރY8}��V�ްam����RnF�H�s�q��=�[&��\_5�'tG(��**"f&��>�PUD��aCV"�4�%4�QU
��MJ�P�)J�
�JcT�)CT4
-4�Ai�(�0X��e*E"�T�}3��S3�Rd�7Se����>���R5��Y��F�_^Z�oo��9A�)e5���錞�i�Z����x��l�}�+��:އV�bi���\+�ټ(���*����/m����j��i;K6e�C{5��*�u؇ !q���直$�Y�����C�t��m�ލN��׍Pkń��`�3�M6�iWA��0������������:�_�	�r̡]5�����4U�������&ƚ4gﾈ�"r�ʪ_�ҧJ���>�Ǘ07YqFf6*q}��J����1i�s=2]�a����5�g�\�20,Ra"�ګ�^�+�1�k���2tz�0L_����9�q�_�7S�7��4;����Y��lE��z�ԫ���
�+s��DV�h�OA�Kآ�xL�+U��'G1�v��<Ǣ%�ڿLV-���/��zkR�1)�a�$��c8m����1�������X��3�f�נ�ěZ�[]�b�ɟ3�������e�y.5����ݐ���*˞m,�0x�Y��(���+�pݬ��^w_����<�N]�2�Ͼ����n�B��+��,��1շ�5�����x���=%e�V��gW��ųH�N�o(�N�z��V����ӛ�
Jzk��o*��,@f���y�r��w��N~ܴ�2�F�b�0�?�}�DM^{�ʘ��v�3����p���;���z�YY�޼&� �~�C��/$9=���3B��=���,,]�Pu�D�c�s�d�u&��g���]O��9��|2���g���r���ݗ�ؙ�[W���Ռow.�dod��~>�r�\��y����5�5��ڱk��V�T�
�׎j��6b+�g��<��˔By�yk�Tx�ƴ�듭(b��F���꯬h�[��[��!�LW��<8���G���5w�]h;�u�~��X�+,v�QX��rWW���0�Q;�=+�s����S�g(���A�-��)1 ~������K����XΜB����z��y�JR`��}��gY�[:����XcU����vΙ�R�=_Ï�����c8�k�T���}�ȉ����\����=����U�U �����h�if�y�����wc h���^�X���d���ݢ�=�3(�.�n,`�3rf�6 ��R�A�ŉ�bج�ϲ�9�luҝIK�������D(�^u*�Ù�Xj6=���%��W�q�}�)0�jV�5s*1��ޱ�n�}��PbM���g��ݔ��f%mb+�j���[��7m�:��o	��i���Dv�6��y@Ƣ���D���]��7(��pa|�!�`�Zގ���i
��7&�4놊���IIL���1*�)*�AH�2��UUB��EP��j���1��B��*�P�(Je"�MP%�CUH�TPJ(��U��eQj���R�R�Ai�R"E������H"5T!T�P��Ti
���TP��4�U�M,Eb,��IT�1i�*���!L�EB�PQhV2��Q*�����{���|��%�e������'/���'[�J���LΎ""b��E�ё���.k����LEz�^�;�`�$ci�/ƺh���Oxႆ���[�w[ړJ������k��5��7[6����@ �n���)�|�?�}��W��T?ۙ���Ǽnv�K��o<��}��U\8���i�^k/���/i����s�f.C�ϭ��\N�<Z=s�q�(-����Tڡƨ+mte����{����]��߾����_�|�^��%8��j�$~g�S��y{�~�dT��Q3ip�����X����f�V�	Uo({�:���'��b�^W����e��8�xu�y�9�f�璼x�t�R����X)l��\قF���D}v�=u���g�*��Ƕ..��(^M����}��׳��Z���ˋ��z�h���WV�o��S�=
��;���m��&soʏ���s��ĭWZ뮅;s;~t�5��� ����ꯪ�5���ȠoV�����?Kq�`%�X�ǜyr>�X������|����G#�Y�c�x�������iH��tk��d��ـ{���(Q���ӎ
i�0g��#�.	��j�Ai�X��0���j��gηD,���ͥ���������xV��5��G��^�*R����8/x�v1�u���������-]������p=���6����Gӛ��yϛ���[�F��`t:XpS۰�g���R,47��7w����sG��J=�Kӎ��� ^�%�/ρ�n�����D�Y݋�%��T޿=Jp/D��rQ��r ����nj�ܼA����.��B�\~q]�V�]{��kCMv��Gr$5GuH-�ەk�w���IW�a�8����Kk2`�(�y��X�\.���ufaۦ���N���l� ⪳y��ZZ��=�W�yۅ	�����-�fEQb��a���µ�S����>�2a�sk������r2�KvD_�s���]�C|2Ǝ^wƺ�ዅ!E�Σ�-*�y45#�ר�W�}^�ޯ5�-[��ݻ^��aw �fˈ��ز��L�>}� {yV2T��=��Ǩ��ݜ��k�i9�7�x=�l�'Ig��/{l�m6���4l�t�lr?K4;��q��{7�T%\��RdpG����p�W�fP�Vh�ͅ��u���Cԋ���I�x^֢B�W�O}k��狰���]���Cq��!�Ÿ����� 5K3��3�
�VS�3n��| ���3;��B��#�֪rqgD��|Lܔ��R��Ag)5N-m�\��om�F�!ךia�oo���)̂�KEø��k�d�-E�����#@���k��\n�ֵ�f�(}�H:�]��ܲVu���1N�T��TT*��ZZ*������S��-UU"��T-T��R�!J�(�S)��%%*2#	B�QTUª�)!LU"�TTDX�E"bb&f~��b�]+Y4ĸ�DeR�%j�u�X���	��~�w�5Ҳ���@�i��췬�K���k.ݥgU�i���7�=ٙP_bk}Ad:mP�x?xƔ+��G�A5���nOL0]-Z>v� W%����s2����lq�K^��M&��|���r��v��-��T�k)v����ս��fyk�-֖�km=�2uQ�YRf�Ou��o��׳���Dw�&׊�2'���!�V�x�c�'�ԍ��>�d}������}�-��*�M�:{�6��8I95s1�Q�#}�W�vM�V�8bs�Ǯ��6=��z;g}�/�C�r?����J��^��pو�M��U�U�Ӯ(Ls�>��`M���s���D����-�g��:���Qլ5�Ĺ��
�Jf����hs7wyl}êy-�.�|o�2W{c�a���'�3_u2��G�Jddq0�8v�6�wvs�^����`|���^��u�j���G���5vfn{�Q�B�;������G0��l$k|��������J:�C�ni�ˈ�)h�	X�^ۏC�k+�}<dӅ��[9����bf%��&�@ІE���k��gKz�G��[�av�xk�����p���*o7'�}7�T��~k/739õjy(��]��	�8h�۩�����L�����OdG�u�'�m%����0��x�����C��79�ž�՝��Z1n�n^�����,�ӆi	��	�ʭ��~~��C��'x�o z���V���H ʓZ�d΍.o3�R���+�̽6��w���Σu�j�m+#^����SÖ�[���"��6U[�^�<8%f�b8]pޫ�Sצּ��Œ:���)�r�7x�~�J���	��Uy�\fO���ټ�y���;<��Dye�}�W�g3
.&��~ݴɖ���K �ET{Ҧ��3b��u��0{���~���Ǖ��;���L������=j,غN㍒xA�G�x]����P��� >߯���y���{(
�֏���6� ������W#5�sT�Q>}[�ޅ�v;��J��x�.��^����� �����p� P��RmX�� ���'���7`�H�����yyG5.�Gy��q�dmLn���/��j�B�p<�$����ֵaKiՌTAŪ
����)R��&�+��[�FY��=i���
sw�F%����SMΝB�M���Y�]��Ԧj���gJ�P�jq7|Jˮ1�ڗ��gN�f]n�k���^��d5�/���:�:os5�\J�p��61^+Ӡ6ʸ��:h.{���㵽���(�3.)�:C:�Q)GgA��j�kv�j���cSd�Ri-K1����\
�����7�-�W�-�v��
DT�"�#"����RE���V,V,F
��b � �b* ������
��+8���ｓ���HA}��*���8�/f�7��nu�Ui�=P%0��;fds
m�@>��0��51���ޥ#%�+�0S�:(�2;$b��'�%�w�k��W.Y�
|�mK�y�g6[:�k�'���k�s$�D�D���e��>�Nξ�`��O|٫<�n��Z�M޾�ƨ��t�Bv��B��ѧ&š�#�׵�n?�'?�C>?��B��t��ĳ��z��]�k��w�+�y�����#Yk�10"��"�wnW9��Hm�k��Qb�E,8q��0��b��"<e�^Ɖ���w&�$��VM���,����:HHR�o��Ƈ�	9��oJ�u��ms�%G5*�"�5�e�n;� �޶`�h=og��OV��m�s*u�03<Kѷԗ�]Yk+5%V7N	�^U�Q雌���so2�n���C�_g�a�n�y&�&<�q����Dԯފ�n�m�v����3�vR!���8�˵x}T�Q�ωw�%B������;������z�h���,l�ڹ�f����I��ٓC�Ǹ�����O�����z1b<��9���m
���3�j���ߵxe��H�I<��#� ʿ{�[p���u��Jʌ�.�q�k֩�4���_�YX�=~Y�2p���sS�o��l��I���\d�O=�'k�a�Ǯӭ��j��[��n#x�VJ��ςΣS�%	�i���W{����0HК���=���s�K=S0+��Cp���
���QӮ�X�f!%�������F�H������*�����X�e��Cd-��T�H8$Ͷ��L��:������ʴve�{R����Q&.��UWU5{�g`j�uq�0$s.YՇ;8�'������b���Jl�-�e�GB�'+u��зC������{zG�F�m�^<�CޭȝfSY�$��J��f�rT6��,Y�sq�w�%��ʘi�u>��3+-$v�,�K6
%6^��d��x*�=^�&�c�4A�Aj��O$�p�N��#M�ڵ 6�I3}���(�=��Wޱ�P��"�n�*{l�eKBm��7't���@�we���=�l^��s�y�_�3��Q��.�ɠH��������nTѷCΗ��e�k㱵���{�f1�yr�Zj��?FkW�9���V�>��1�eM��`L]���A�t[����iZ��oEh�T�T�,�EFw�d�A�wrs�x���]�X���)u�G#�;�/�������ST�#"V�\��$wp�l�Eڼ5��Ѫ�4��;-V&ʎ[x�D�J��H�$���z�]V�v_lqn<��r���2����R���|U'���k�LYFf���`�!<7�'LjL;V֬j�^��#�,gVm@.$�8�ǰ�������Il�8H��Z���kb�EQTX��PEX �X"�cV
�(�����V1��PX�Y* 
(EY"f>�=Ξ`����c֐mL��]n}�t����������{s��
K*L2gQ.�^�߄�&E���x��$�/t���`<��1��fs���'q��L����	������uN\W�P��U��:��6_К�����Z�j1X��Z_{K��#�\sM?B��#��s���B�mkۘ���h I�K�י¹�{GS�]�)&�y�g	}���wGW��v�"�t���n��F�X͙*�� n*�<�hkHDߐ���J� l���@o��R~@��g�,��.�IEa�2�% �$����W`�&��/؉���P���d�,h{v����R�'����E�����I��ȑ6ѣ"�Y���?B��08���PwK^�N��g_=���u��	�l^=�9�c!�Z����#hR�O�Y�=�W��ln��>.���]�m�[�:=�'e��uE��j�Z��n�]�!���(���:���q
<�u��$����6�R�{DY�HX5����{�޸M�Y�S��]���b�2�b� Cؒ�ܬ�?�C���O�G�����r��1�CHo�*cL@@_�p<�m]���q�ȁB��n֤`^�(��������rg\��`�b��?qR�{nm\�C��/+CT'/6�*!mg{�9J���A�CH��� ��J����ՙk����~~���v��E�G]�ǃ=��);q4�flx�W@���	��-g�����s��}�{Ƽ�u�����>츪�.���|�b^��\��wJٞNw�!�&���^ب�g����VǒN�c*�K�+��yfHP^IJ����v�{��9�1��dc63�nޛ�T�c�B�QA�.�U��@��d�u�vu�Q�Hh"�1����x\�~��){�SZJ�R��4��{�����^ש���Y��fkt=�{�*�Y��-X��4}��%���D@���dU��� [bキ܊z��J��ѳ�C`:=��u
�ߢ�+����]]7��_�m�žK��/�r�>X���$��Ppr�O �zy�y�{H�ygiO˫@���G��O�����:��;V�xMC}p�s��. `!�fr���uG~|WHlu9[Qks;���0n�#t��T�����s�U�,"��4��#1v���;��R�uS����Owq��P����6�#Xy��gL��;j�8�fNwP�u�	*�> �⤮���̃�>;ݲ��Ib��u���9��h��̾q��J�n�a$��&�[�5�{-�&�c�|�KL�ƒ���Q�����Q�\��L枏h���r�1-�q�q+XgV�w����I�gX�mn�幞� �ȉa�d�Y���H*��E��X�*!�UU��UUTESZ��o����]Ԁ��tlW�[���_K���Nd��|�Y.����j�#m�^B��.�t^��:J����gV�zj�k��Ƕ]r�W�u	.���>���J$f5g2�`˚��>��^YQ��,Ŝ�˯$�<)�*y�e��y�ǙR�3�w��)�����{_�=��!yd�,�[N�ow�j^LV��׀=�uv$�
�����U��6|�p����ɬ�Y�N�:R�r6k�U�m;�Y�53��Vp�A�x��Y�쭃_w��u��/n�shi�Ybl�g��W��jwK��E���WPV�R�w��2M��Qa��lܤ�.LʏUG�Qg�>�*���+-n� &��w<=��AR��|=��N�i�����WD�j&¹�핷��vڄ���������v�/������n�.Vk!�]ku�	�͘r5�U�o�g=���;`�A��g1�c��Lؽ�y�G<�^,�d	爕d� �׾�YzV�X�y��_���������^�Ьv�Tʫ�V�9�z� ���^�f[2��}�u�J��:7��j�G5������Q�C��TL��=/�u�e�
��x����6���E�@������5zQ�*�l���>]]�EǱwo0a�Y/މ�����ʻ�n��6�����xu��������.���~[�Ηm�AX|�xeI6��R��y����[;kL���WV��|i[�eW�嵩�rU��G���CVܭ�~���<Ny����!�j�[�n��{��b��.����&�^��&�1o��]�V�9�L)h~��1."�����7J�}�f�"�]CѾ��ϐe*�=�ݺ����e����M�w��/�{S~�H�?^(FB2\�M�&u�ŜJn? ��PO9gY����p�@7k�V�l|�U�Ç�~X$gӷK_����-�hMT<�c*�k�ױˢ�{WӱX�Zs����c�9<}�lÌ�hm���W^���|��Ȏ��[��hv9����l[\�w6M�C�=�����U'�E4���h4H@�h�~rB���RT䐁$<~��ĭX(-b�>Z�[���,_����B�������$4��
�`�~;�f�T��p�+��z��n���N>�ҿw3��'�z�����j�a�z�6=������7�k7񰱞x\��	�15�� �$�򓿏��/o�~A
����$�����$����XE�Ic�<�s��A��@ğT�����������D�G��$��@>U�X?��@�[_!�OwЖC%�����bGr�Y����*��fD3������c���`0��I�ωRB�ww�/�W�ϕ�l[�B��{��8U��IE�ϕi�V��X4a�yt?���$ I)�e!^�?zg��򟴒��=H��-<�=>$8y�����c�������?`a<��ʒ$�����zg�Y�9?�����-_���Sd�(2I���?A����' ���>��)>&~����I�$ ID=�A���"���=�������""��!$,�>2B��������I�h*O]����+��6bBy����!$32zl�1��=?��y� ��d�I�B�>i���ÄLb�J��9�9��i3�>�e�P�4\��P�,�0�$:X>���t懰��$/�G�!���g���'�~�(~�� ?�����K�O��/Q������<��~�}��������n���$ Ia�/��HE������$=�}���tX���?S���'��<�[�}:���#a>���Ϯ�����s?XC��OW���3|I�+��	C�z�K�a��z��ʽ���i�Ԥ��zH~Ψ"�{q^�Q����� 8l�@��$����,}~��~G��5�{|�HC�'���0�_�C��d1��T�cV��U�O!��"�9�z��rE8P��:I{