BZh91AY&SY]$|��߀@qc���"� ����bA��    �/���fk"�f��(Am�Q l[fi�����[2��Ell�U"���P��H�[T���*��3lѵ�dֶ�l}jNڃZ�[,�Md����eM��km�[5*�c6��KY���F�cZ0�����[R�-�+k+m�I�,U֊�ͶV�mx>���T��[��#j�6��V��32�6�#Z�Ķ�ʉ[F[MV�a�ա"ړ5Um�$T#Vօ��-�D�V�4�,�kdٙ�l�ՖJ�w�s�Z�i��@�   c'�jkӓ�͵uV��4W ��[��jm�u���UtqS����j�V��tݴ�\�Ջ����UZ����:ڶ�k,hF������6�   ��t ��l�;��� ����  1�u��g' u@
�rݡAAAqX� �9��R���h s�R��&�ʭVl��V��a�  d�ڀi���.  ѮΜ[P�[�`���5� UM���� Q��w����� kF�yu �{t:s��zPP{ݱ�e�mUc[mVmY�-  u�  =.Uq�A�:�{�J����P�Q��)Jw��� {<7�f���  Ѯuw (;��@�7;akk5,���m���ke�W� �< 
�m�ܠ  �,t: �c �
W;�-��� �ha�4�f��ipuC�m�u��۶h���� (Pw.,5�#����Z��  � 6�k<� �;�S���Q�� `Ƃ���ji�v��*�;�ڸ  ��(Pb�Nht pd��6�ֲ��m��3Z
�  f�� {�\�U.��` w`.�@
���B���� ��s\�l 
ػ� hѺF F� .eSf�������1�  P�` 4^��@���B�j�� ���P��F ��8 mv�t:5TsK�2Fi�+bժ�fՕ�*-X^  T��]܎� wZ� 4��(n� D9� ��ݳp$:����ʷ �7\:�gI�%�[,�Fښ�P��  7^ ��` Q��v��I� ;@ .�  mE�C@�梀Q�� PL� hx   � PPCS eJR���`LLL�i���i�RT� 2h    S�2�Jh��    j��	JR�р� �4� ���M�L���CA� ��IR���OS$�&@ ё���t��d��9�M�ǆ2R�%L_P�64�Բ}-������>�/����~w����j�������e�Ukm~�֪�o��￪�;�UU���_5������^����mƪ��eÀ~�+UV�{�����cmV������_�����k�sZ��ֿ�[_Ym,���,ڿ�[^f��6׼�^�m{ʷ�ս�k�5�-oyk{ʷ�־3Z��׼����-�y|f��-�y�{�k�[^�Z��k�k^��+y����5�ym{ʷ�����-���������6��m{�k�U��[�k^�m{�k�[_�m{�k^�Z��׼������k�[oyj���y[�*���ͫ�Z��k�m^�j��W��{�W�ڽ��/y�vj���j����-^���5^�j�����Z��V��U��5mo��k}�m��V�y���y����ַ��[{ʭ�򵷼�Z�����5koym���[[�mV������[�mmoy[}e�����{�Z��Z�޲�k{�[[�Z����k{ͪ��kkoym[�5Z��j���W�֭��m����V�^���km�6����{ͫm�-V����Z���V�{��W�U�����{�V��[oy�[{�UW��m����kkoy������W�U{�ek�V���+^��6�yZ���y�{ͫ�m^�m�+^��6�y�{͵�-�y���k�k^�j������-�ym{ʷ����[�[^�����3W��+Lֽ��W����ǿ��һ��z�?fP�ߵW���b,
)0�����ݛ���l˩r#�r�u5[��� )����wvé�Gt2Km_�(1�㡦��+w�/).mo��{�],��1Z�
Y��(��1SC(��ܫB�V4�Ԭe+��k"�mWVb|ަgH��D5j�U��z�LF�� �f�cb�L��mj:60nK˸�xt���I�����bw�.U�^��b��<�c�(�^ݨN^6lP�0֖���[up�Cl�V	��s ���X����IP��H���i�s7Qe��߷#;W��U�e�F�ܘ.v�N�bS@Ր�Giʻ�(��Y�TIY-b�`�x��-Y��/��Z1S\�r�oQt�4v	�tf�tt����01��BVG�,<�ݳ	�/YF���V�Y
ݳtJ�V���
tM�jΛ�.[��,J���P��E�O��H�khh�X3%�EM0�S�1��Ѩ���!Z�=3^�7q�IӅ�7mLA�ZYW3q�sr8�ȮF�]�zӘwjP�9�.���h�6
A2��敝E>���{�:�]֭�oc�ͤ�S;2���3I�*"Eek�5o�#��ʡt��b�ZD�ye�vM�,,u1��`;���2�e�+c�F*��Z�[cX Y˛��ĕn�Mch2L��Ey�(�T5�ۭDIy�Jr��v��z�AJU-�'C�M+B��	@����e�p�Nl�*�![�5�vrn�Z4/�+l[���ŉ�N�"�ڟj�r�����k^��� ��t��B��ԒJ�C�f�ff7�mL�͋qÆ���6t��v�>C���8V�tu�7��A%�q�a"m���M)u.鉃.�b�ZX*D�G��e�V�-E7F�bY���/(���uT�&S�6lT׆���J����O�,PƐ����a��`֫��0���d2��YW�Ͱ�;�]Tψ�Q���b�3^�^�sE��j)�u�+^�����ƨ�"8v��LZ��Z:ͫ��� zp5"�.�,+�ٺ��M(�
ź����SP���v���Vitr�Ctب4:��]��1^(�NJ�*�S��kf�?����3.k������~t�v&�PZ@^�_>�9�K|z�)є`h���ij2�ei�3E�i��@ںݶ��F�M��l��:�H%���6�<��;b�I��&�7m��E�����'b��� �LV�[e7��efC�X�(4�]�H]�
�w�L�*��ƥ4h�U�������F0\v�+0:u�4�%�ݏl�\�6)����!����N	�0[�f*�����[�[���X�c$j�Q�f���%;JmG�&�ʪ�st��VӁ͵���(Cn0�74<ke�Lۛ-��Xb0���2{kBC�l��խ��A�W.���b���&�����-e�J������9�x�m˓1	������1u	I�ս-B��(�u$E=8���N�
��*TR��i�#����6��M �����Q�ܛ.�
ٶ�X�Ш��4��-��ے��L{N�K�`�)ZS&�p=��m��a-\�D�p�G31��&�Ô�,a���MN�	/V�;�@fM�k\&1��z��c �%@��@�Q���X���YMV���2��Q�������I31���P(m�����MJ�K�2#��(��/]�oo7Q�$$1��]K[(�g6�`��0n��U=�F�I-�s$m��9B#cM˫ �R���uJLәb��l�l�z
J�[f�Q'2��eA���ܲX8>���n&����r*�bL��n�h��ef&����gZܵɁkDf�*�孛�,zY�#S�F�����ϦV␬"^���d�S*wBSH��+wBB��BɵT
*��V��i��+�p_ٜʱ�;�y^��S��5�q
M=x��t`@ʼq�B�!w6V[��^8�Õk��fdl�ػ�U��j��L��3���4CA��;����z�tb������h�[BXY�keaI�x	A�5���wh	�2�S��Gh��a�Z">��;巣�C�B5�nƌ��̎�Q�t��+K3���8���O*��(��6�W�'B���'L.��d�(�wm��sz���6eLS^eb�Fd��%�m5t�T]`Ƴ8om����1�i��2��/[ũ,iKb1E6	R��!@�Rd�4t����弔B�3M�+�6�b����}�{��@3�I1LƁm�A�ٚ���(��W�;�vj��l��L�[G.'7����k���=r��	pMn���mې���7^���6ێ��tA��mJxlk͹X���[.6K@e�U։�9b�I�Чi�1gi��!md.���rٶ�`�Ă�{6�Ӳ��ҙ��!���Ib0aV���r+X+)�ߠx�Q�0nݛ����i��ћyKV�Xd�b���	�}٤R�@zw��� v��Vgۯhq2�!ŖA�fmf����9���nM�r�d i�̻��V���[HMxf+�O"+$�T��mfmp�o���XdoS��;�iP���54��c��Z])�h�R�;���;�=6h(!��ܩ��Y��֫J�:�.�)(��8J�ԙuv� .��j���ى��J��DUbB�D7n��12�����U�Z�i4��x�Y=i͏%������ᇏ0yZ�CWx��Xt8�8^�����k�sq��[F:��bT2��٣+�1�"IM�
Ɯ����<S�v�.�̳l�Q�;�C��,�����ޝ�����=т���B`�M���ӳ����"P������K����p��6��TU�p��)]B�J4$x ��5�ٸ�WԂ0\2�nB�P��;���7�v�S3[F��T�R��2jeX�2Ԭ��e^��6�Z��2�A��,F]�h5p���I����q�b�aq�&⫀�����^�ߢ�� \��$ն��lA�"���1w����V�i�'Y�%��i=����j��$��� f�Lk��6�,���̆����lp5�h���u�`a/^YXBd��Z���li{�oH�ʔ�\�g.��x�tV�7f�vY�=�x������9��������0��ԛ��hjr�@�+f��@���zH���TN͡ �/���-6�a��[�g��xd�)^�
�7o2�f��f�7%J�դ������ꎹ1H�v�N��24��F�_^6䬃$6^&+��9����[��Tu,������7k��Rd��i��hE��5�����*@��"A�1Pِf+حL��Mf�u�4��Ke˺9��&�����0��&��U��2b�A�W�GX,݊[��gsV4��sn�-!�ٹ��Ğԧ S�P�U�V�[a��!	�����`����cw)�1��������9X��t�n�,jͣq�o3�y�AKV���Ƨ7�wW�g��9MG�7yA�S�r�$e�5ˤ3P���{�k4�^�P�q-ݚ����ӑ�d��Y#�̡!5r�r���#��`���F�uV�M6�mk%�Fj��2I���
1C�;z&��!�2�8 h�۬ń�щ��B�شp��ͩ��-���N\��j$��m�؀"�n�M�P�Ւ�31�m�f�%��?��$�XeU�q��y��vT�&nJ8kM�mAM�50�$���ɎԹyR���sM�r���ˁ�r*�OEֺ��S��a��S���:��W.]w[��(�R���R+)r[Y}��\����ckz�Kb{�J��v�sx��-�;6Ei"X9I��E;��B�����oT��(j�A�g$�Ӷ�|��>lQ�h%g���dQ��NU�?m��3N�)�^AS�kǳN�l3+�Z�a��H����j-bK��V��;�r`ӲZ�ӡ�"Ռ7aX�t�s";N�X2�Gb�v6*��,�#��6�E&��!�n�f�JV��	�%R!�kp��V�4�KP�v>��ݵ+o%n����*LU-������1��ffl�m�Z�Z�sE��EG3P�3t�oPn��r�!!!L*��d�fΘN,�
�v�v=�1��^$�V�f�~U���͛�ݘ1+v
��F��<��h�q�����t������%����u��U�EǸ�ul�-�́�M�;�,�K2��[h!��Ɋ�*�M�a�=���|��$m��îQɊf�cV�Oc�4�M)r�h9.m�v�fR�3E�"Ӆ2���,Ӣ�a�c�)��Zk/�!�����U�O4�ʐڛRS�h��/f`�5'���d�e�Xk.VT˵Q�Z�����sv�k7hi�^�3(d�U�jl�?�ʣH7I�pϊ���J9�0�m��2<{1A����[�5�h���'�.-�a۽��r���?�œ	.،j����1�j�.@�V�إ�X/H4tI6�*ׂܻ��z�j�̄���e,b�Y�,K�cj(膵�l�,�66�r̵�El��5n�AC+H���Dyk�O=�Y��ź��ѮÕ��{�h�a�� �Q�C12v1%-j�*����&��LY�F2P.�����O~I��W�����ot���h�R�F�Sdѡ�8/�ϕU�J���ǯL�8��uႲ� I��/N�4]�l8�)iǑJ��Z�/� ���+KNnڹ��3j�;k�$PՊ����`��eZV�ē8�p�v^x��2���1�|�cJ�V�\��a�������vC��e�T�a�#ߘ�U�;�R�׵gw�����Qd=�0,PF�TM�'ײ��f��^�z��N�mk	b@YKu<H��Ƕ��r�ot����� ���v攎'MS�v�����m𰲆�o��.b�r�k2�����JMi���\�cq��m�ZD�c�;e+ ����ˉʉ9T*���F2�"��F(���8%6���ݬub�+=o,�
��CGo����;���8�FL�6�S��)i!�h�V�-"�.�с-M��4��l�:��ӷ�uۡ�������MsL�k��m�4����y�a5j#�� ���S�N:��ܽ����w"��vV�
��Y�h�����Q�ں��bc3��N}x��2��g�N�E�y�������c�,n[��A�Tq\�t����{@��,|�8t1�(*�(e�up�8�2swBǴ����x��/V�d�f�C��p�H v����dCl�n�� 첥9Tw�҆ah'6ɫ��%�~[��i��j\gpu�i^eӛ&c�_K�jзSSb]�@����ԎP�Ŭ�/m�N�Xc�BVbu�RmU�H(�����n��EF��O%(�fmm�K,;5UN}Y��bvO� ����UuN(��	�I37a�>�2�,�7!��pP��\���>ՠF��F<lGz�!+D��v��XmVi�I��TI��n��Mϛ^�������Rǚd�oU�3%�ଌJ^�݁Y¦��s^y�;%eӠdD=Ko�-+J�j:Z	��f�1K�bsfZ#lM�j@r��FXe��퐯4H�ĳ+t��w�
��{�NK4���~�Gj��)�bѵ��$�,�Ygvc!�Mu���l�-�0$�{k�xu��kF��;���6�Xb�V/ Op�&�ث�~*ɰ��5j�t��Ș�㒃N+������E�{�fQ�c���a/Qܦ���Р�T�T�@�Ӕ5D�S�wS3B�_�_l��݅��/Q�l�V�v�{�.M3�;:��v;��wSPVV�j� �պ��s.����
�wR�͘ձ�'�o Le� �ݙ�:�e��Ұ�f�m%M�Wqjz�:-�l)�3/q!WE�� ��-�㚻X/:l�d����ʔ仭��m�-"Pn�p�&d�[�%����e�%�-����B��F%K\��������m�M @I�ioh���Ǖ��h���b| �2�zsol:	C,l#opUܐ�r�DQBI��D��Q��wP�h
��x�����Ӑ桕�Vm
:q�d	V�a��U�����]a�Ct��U/�az�9�&$�V��T�wD�N�L�r��@�0����A݌��qc*��j���x"�b	
qνӲ�F���+-3����g0*.�v\X&h�$��	����4��r�VfU��st�(usEլ�e�[mb�X)�J��D��+b#5=�p�x��wm����#�%���vފ7s$�7� ܥB� ��Æ���v��J�(�ZS�mWV�ikAm�d]"���#a��AV+.;�*n���-�T�˧�V�j����
v�r�$�T���z����, p�N�����[6�kd<�7Pgn�Dvv^�N�Y��ct�O`T�̟���iw�,��^�qn�5t�%,+^jxF��lp*jڠ�`G$sUJ�t�L��w0���+v�[+Y!ـտ���8��5�Xq��q֊��-Ǐ,���X�Y�S3H�RP�Ԙ�f�L��P�7e�	������V^�����S(Co$���Hʺ͠ꤼ��3$������0/��%fZ�e��%++v�^����8�ͦ���� ;S%H#�ܨ�9��zF��ש*dz��fC��� ����� ��o��1N�>DA�� �4V�xV�� ���/ �bqG����L�F��zn�
H覊��(戃�+ua��V�Nq�48�kl��U�
"��&^�sr.ĸ�dG�RqMGQ4��H�A�F6����D��&���$�,��V���l����Z�����i/o�g�ʻ A*�`����D$"m��F	�����>���`�3o�|�/jr`������7����}�����{?@?��zT/_��o�D<'ׯ�}�~���Sz�PS�LF7O����f���q�G&�:�ΰ�ϯ��K"�I��.F ZP�cc�X�1�fW��5��\�ٱ�U��w'v�.'�w�@Ars�,j���ջ(�ݸ�����{5=G(�W�f�T�7��T敟j�`�q��^C-Rtyr����q}�ں�0lP�U�����˪t)vwm u>Ձ��jH�7��J�w7\�(�\0�ڵ�6���G����%����M�%E�Y�3���)�T��)�m�[مj��'a�mG�$�V�|��mH�U�wo�pN�|�����\��8e�x�췛�s S]�[�M����t����u���WRYC��]ϪΤ�U�R��X���!�]ըn�
ҭ�R��ZlUA��/�JGk��][Z�-[���M���jt�Tw�n\W��OUe�,�Ӑ���H�:�ݻ�j�2������N��el��M�Tm�#�Jq��'p]���\����Kf��Mg��pZS{	}�]��2����+��kig�.�.��g{-�z��6h��֛˳(F���9�y����I���\2�)�k�mtK���ke��6���1^��M�1\:;��l��In�������2��4������e8k�[gd�jL+"EE��K�:m���dqwy��J-�ٜ6@�s�J�5>y����Q��Vc[o�����r�0�ũ��HE�q��S���~WUڰJ���F�@[f���ÆV�u��;3�t�l��H!1�����W��޺��zP�k�Y�[�z��0[�}ݹ_)�����Rv�4�r&�_"��@��unlͰZB���l;h���*����ZS����9f���g+��م����P]�m[f�w1ak%;sU�b������ҭT; f5�5�k�k��|Lyb}S�f-�4WPN�v81.��|�r��d�W�4E�½��+_���JP8UO�h���ϯ/���YΑ�ٹ{;t��>��]w.���ےJ�+g:ɭg\��->(��e��GY�����ǱU���Ғ�@v��8��.��f�G��q���\j>�y
��im*_c���;�&_t����\�W6�J�3�9+��y�U�ަ���|�[:�l�ՠ�t`�=U*�|���[.�f��Yys�|u2I
f���C�����������$�:ɻpu���EB��K�#e$����`����l�ه�T	�fV��d�,�͛{m����� �yb�P�	�i�����;"߯��	�v��8/��Go5�؎��X	���b}�	sE�wZ-�hz�}�_ �.W>C���sc�*�i��S�> Ư{��4�Yå=����u����Z�5�0Pw��إ֬����E<t#���9聻�o��`�C�vn]H9B64����/7���ؘ(,%��3�j���NǎS�|���Z��eaV@ufd�//���uQ�#�˥�#W�\4)(�7{��1�I}�\�ϰh�VR?u}B��9j���	�eXnD���|���Q��[v� �Eթ(M �B+�Q#z+��s,�gG1��˜ �;�u�s ���N�֖0��������駳I��������-1U=���Ηp�vf���e�+8]�3i������5M0����\���+6�B�(@^�
�fV��boëV��$Q|	|�2_]2�VҮ�|�b��j�s��� -Al*��c(uU�;���i����UD��c����؆hKF;�ڱd�Qvg`���Ov�B��/6��:�첍�e
�ek��E�I��3�*�=���&��y�\OP�u��� A�D�N!ٛ��T:�щ��d*m�\%��xʉi�l��=�rT!�C��q>mmEN�wh��sk�)�`��ޖY2�NR�{��M=�h&�!�h-�e�͹όo����y�P����tj,45���3K�7�y�����w݂���)ۤ��VH;��[o�˭���	��x�	;57�lJ���η]n7�|X���\F���������՚�I�Y��_Wb��ۭ]�PZ3��={:0���.�&�|�1��� ���ϝ�DV鿋�{���)=�-(�ƻ�s���5��>�������Pf�|��ԃY{ym�����ꩻ3
+�U-��ю���]ֈ��E�}r!�dV��V��p"�ܙ��ʁ0U�)s��ut���I�S�[���:��WPwEKz2�E0��h`xq�^�P�x�T�c[v��y�6ҍ��N%\�֖�2�^�d��op�J�-��&��ys��m���c���E��������l̗5c���v�c8�5���)/��F̗ }����Ni�RM�̦�m���VK⃅>R�Z�	b�v6)�E�Ż�6K�W��L��Tڢ}*V�0܅bc<��^n��}]�]���F'M��N	��3^�P��/�����՜v	�,/��L���)>�����Q=�y�F�,>+w�]�݁U��I�\���2�4 7��ls��E.��'�P�=;f�獫z-�`�GE��̤*u�op�y(����m�3��s�s�߭]�i��t[�S���	��l �޳��P��E��kʝ=�^��̱�?
�ཱུ=ض#�����7��s�0���0�;����R�.�\�&HM}�t�l��`�� �m��wis]v���<�K땋�־L��JI`���5��b^ʵ���y��:�Y�Y���&�� �Gw\��u�s���hA�QO:E���B���t�x����"B��&:�zuᬸ���Eݚ�*YI���1<;�lin��x�\���ˬ`�!�6+l�C�V�4�����4���nP0�fv���M�6G*v4>x�~gG�ʿn�K�*졊�ƋLC�hf�QmF�P��.V�����ow]w��ްo�h�8:�4�� E�:Ώ1,���n[���d��_-�j�N�ûb��k��W#�ݘ�ݓp�oI��c{"����pv��Ddw-뤑F�$\���/�˚�鍢�fV��m����,������P�$�;n]�Y�01�Y&^�X5�����{gV��E*�Ӛ�e����*5��f`w\4�٘��*��a �ñ�s�s�wg6.�30V��Ke�/5�igk凞��wJ5��8�I
�F-_Lbet�4��X�ՙ�w��)f����9rjl�q�kb��>F�t�U���n(��j]A�� 9|�A5�m��t���:��~��R˶*�H�5��H�x�f�[ӵ:�(�V�Uz,�
���|u7y+���R�Y;���[��!4��m�	M�2�0� �++k!���w�E!aLp�}�]�Wִ�l8�rv�T�+3r�����M�" ��[ڃ�/%FV�X�y�;CV�F�]kk�^��x䮔d'�]�̵c��U,ͫ�/�Ĥ�¤	f��@��6f�����'�E�c��wi{��/�B;�ڗ���ʓ/��zX 3+(闀��G�/��-�Y�'ԭ��d݁wr�pL�*�����8���iK@t{��Ee���v�AO��I\]������h�J��R0<�3��{u��h<W��n�Ew2> �*�+�ۺ��V���i�-�Y�t5�;��C��D��A�}Ն-ֹ�Ke�"�����f��vF�'h]���y�Y��I��8�c�_sj��=:�op���}V��gkj��.�$��C��p:��v���m"�v+�I7$=�w�m��L�ﶦ_mo
�+����>)0N2<E��Z6�v����ޥ]��X���1�Y].���'K@@]6��H��uvVG�6+��#(�;Ya$W$�k�,�wk�F��]����P:��ܝ���ґ����w1�N��C��b�$Z���v�����@�e#�E��F�	�]�1R#�v��P5�Z&��e��@��b)�^ʓ�RX�mS�QR8K)�	��^ժ��pf�� X8x�U�C�/����ۂbY�W�,T�V��Z9�z��3v����J�A����`Q���T�������j0�h�r
H���u�:�jhq!�3�l�O4a5<]i��#�wL��h��;ww�� cvI�K{�瓣��fF��ׯ���)t�hM��QpQ�[����Z=�U�>��۶Es��Й]9E�ȷK�#z\�(�k1�b��ݫ���&R x�h��;�a��Pd˜:��g~X��%S}՘�E*��DHo%�t��)ǽ��\��h�KHtt��_�f�tT���s�X��+���Y�Y��L���Mj����<����P%K֭C+�ѧ���\r�8u�TR�g�:UzV�y��V�'�h���6w���� j�4w���+w�]G0s�}f̳P�>����\o�ۘwE8A�Q�:'g8 5�u�M��E�w̙'^�4@D����i�U���mUJ˱�Ƣ[,����v<+J�I�o����(4�1c+0���x�,�M)�w���m2����?<֍0��h���qօ��u�ڻnH�TU���p��Ϧ�-Y`�ً���G\�NhX�����֥�l�u��
1�i`yG�"�bR���5ӊZ�����v�x(�W	�g<�Љxq�OVob5��no�`F�J2���Z��5g��m]��ӥ�6j#X��c�9s������X�����Yp��,;yu�ek�����=�|���6y6"=����m�?V��}�f4�ؤ���o>����g*^�j�V���\���Ъd�ż"�֮���������qg��ܻ��h
�GrW�/��n��T�wK��Zr�&��R��[�بw'b(oZ2�Z]tF�$<YMRc����g���\Bff�	`�.٘R�Ď���n�G���N̽�!��ajeᎎ�;9V8��9t]�
�-.u�0+�^�[�7n^M��Y2�AQr�a<���Y�]	-��fڷ{K5��g�����N7��s6��{��Ep�lq���B���%۰�:ܹc����@��
�l�rJ�pAƭLg�w4�V�.m��Zv9tӱ	������r&=��>��+�:	�e��!��k�.1���b��sY��J�L<5b6��kz�*��&���$��y��]㒗.�}[� �i��q�̣���������V;k{N�(艴1bB�N��c�nvQF�:�t�J��Ls�}f�Lk6�tՍu��ݿ�ٙ���ט_ ��ړ�*�P��w��/�5q�&H}���a�:&��6�s.˻Ѳ5�l�]k����i�]O&���ˮ�kQ:j�Z"\���|z��AvS��a��j��@u�D|��0�x)_f��/g\鎲ۿ�vP�D:V ��,\T�Z,�$�1��8��fMd�SBR�U3hA3+R�c�nh�f��.�3M�	=�S�؃{�z�� ��ؤO���0��m�xSfQ���P}�8�6EK�ɚ�,fU�����ʒ���0g;Ղ�DcGYn�XV�d���HʒZ��b�ݮ��=u�,]� Z�n=�KSB��ݱǴ�*Q{*"T�M���*d(q]%�n�pŵ̝��{U�	�d��#ڒoՂV�Ʈ�(	��]n�K%+��jL����� �l�A�X*tË��6���Ҧ��Y+���e�D��uX:4��E7�Lr�"L���ӾO��"\�EM\�}�)�|�c�W^M_�rnT׸���Xr�yCI4"r�e��{V����b�;kD:]{�{O�ֽ����C�
����]�>�Kxf���K�3��*���f�	Ug`G���y��+GDs1�HwY��됮6QT�h�2٘qv���\�0��h���]L�vǶ�C�"��ԫym+���W]D���e@�:3`�f���3P�|͌?R�h�p�'&1gU*m,���zƤXR�P�s�Y,z������pR�r'�b���2�9�ݵ}YH����Cz����v+��$Kb���6u*�9����tf���;�X�8�f�{~�s��4����Cn�S�q��k0��B����ji�o\5o �C"��Bm[˙{6_U&ts�ک���C��|i��/C��2���+VF��8FL���Ѩ�n�9�jI�oS�`��qv9���q�����Bκ���Xv;r8�����`��:f��2]�����O0�M���"��F���!������0
�r��)r���ـq*��߈윏q�M��ֶ��;b�Cn�6pU8<e��8�����y+l���[:i��ա��l�4.��ܬv�rSܠ�j'S56Ƽ��c(<8VX��Q������t+e6~i�zKB_t�.�9��%Z�V{{rpz�vt.��ٵ{"w[m
|�)}zs2�7p�A֚U��ϻ��[�O}�E�Vr�c��/u6�^�X���[L�%�-��q�n�5ݮ�N�/M�����t����H>ɯ;.�5po]�Aiq�)�	Ӫ�`K-f�u+r���.y_�k"Z�J��L�S�	ٸ�c2�F"sm�٭\�eY�|�:Y�8�j Ta38��7��G�rmC��ȇ�/*Ї�U�����r2+[*c�V�f�u|�Y"�=�hʽ��<�LEZ��t�Zh ����li���WǇL3������cFMF�r�t.2�����%K��K���A 2!�����򯶾�����������[���j�ܯϾ��x��7�-��|�o�r�9���x����mߝW��-��ֹ__]����_~m\��(-��Ϯ�*��/�[V����������mj�U�������$k�0+ HI	j���+Ŏ��[m��8O��U���̺)��/w��x0�E���A	���Y�s/rH�R�C��^����fh�����C��rLͨ�緩f˜��Q���S�0;�[��JfZ�b���&۬l�wƓo�v,�˙/�N���&*�m�5����y�=���le��P�YXxK}�C;e;��;��ƈKi��#I36���͎�ur���ݡd䙺����>;���(k�(�[;O:�X��N�|3jʰ3��\��$}"m�ݝ�D�����H�JG�PCW��h�W]�엝�+�.v�XXI��X�lɥ��$�)|�saʺ�2ve�2�y����,�[Y/�}݀S][��g5$��g^=Pr���u�s�0I-]�����^	��g..�5�廍?�k�ٖ�q%N��U|��OJɒ%:�k}����<��lsG��#Ӏ�q뷡:��bu��f�؛)��S[;n��m'�-Ѡ&��}��k$Hpqz�Ž��Љ�Cqݹ*]bV���<�ވ:P���ҕ�������(�Y��Nn��²DjV�:WU���F$"�-��Ă���l��z�Y5LK|�u�f�Zt�����*ڽ��8������2�j�r����k*�~;����i��׀5��L�x[�;b�����E��ξ�n�e뵘�,���#���X�U�tn'Ԣ��]x�.�]�,2oN����}zh�Js��6f'�hDv��JY�դi�`�y#l�O5� znAҩ�u΂Y��a��v���s�����޷"�{4���.�|*��D��:?�r0����ި!���ͽh�K�zF�w/0��p�����Gy̅�b����]sn���#�	��}1oG�A�u:����m!9�h�c�+x�\]�7ܦ�AJ�깘��]xS���V���"���8Ar��k�1j]�δ�f�6����
D&+��c+p��YV���S3뺺�!����ltE}A��Tu�w�)��j��7�gN\֒���A¥�1X��Nϗu�*��4࡝����P��O���u����:![�m0����.�>6�vv���d�C�9Hԅ��9�.��CX�5RM3yY��g>y��xDb�w��x�j�� X�Ψ-r���������W@�z(Y�o`�h��_2��ݤ�E�\�V�����"tR.���b�3���K�i>9)�Ts{ݪY8,�Z�B˻Ե .[��|[N�mԈ�&b��6Mn��檿�t-�3-�Z8(5�vM����.�*1D^�td�;P@<ߦm��X)���N��Z�P�W+i�-��8Z�cѽ��.�ɧ�<��H6m ��DpJW��iJ�'G�h�Jr���vY�#&��؝�.԰�=���J-3����ȝi���K���ZY!��иD��<F�٨'��Ա���n�)P�L2p2���1�tLc D�V��{VwiMd��N+��鲶����c�)RWᚖ�o�Mx�gfaWlr�Y{&�NHgV8N��G�[8r��F�+2]M�Ԩ�*]VS�Zf���.������A��9SU<X�E�=ʝ�r�����r��y�[\��PR{J�͌ѣp�vvӉ��ҫ^�X۰buݭş9���bܬZp��\�/W�2v�]��:]�"��/x}�����TL>ҷ6�iY�N�m���K���]Yo`6Ņr�����vT�I%�*2,C}��`���n�X
}�q�Y�U�8{�k�H�j��N��f�1b���Z[�d:f�wwEq�1�\��Zi���pK����973XM��.�¬͚����K;�9GK�6Rq�A�p�i!�}����9��4�����>D�E�PZ�a��K����͛�U#Y���2�2��I�[Oe�� ם��V�<�ܦ�8�f�p�xʭ(Q��9�X��S[�<)�rVk�\��Z�2��-�`�+6�F''f��v�AVt�A��h��{-��
�6���3�%�޾SJX�jIӟh&��uNXɶX���Ly��"��^��_.y��4m��n�B�Z��#�	���N]nr�#��ZY]G�8��K8'R��,���+�ۺԌ��6ʪ���l�(��.:��f�1�q�cUVn-����z�es�I�Hm#x���]m���=�r��Z�I'��.��+� T6netorޣh��D�p����ՠ�$xT��xݎ�����l�nf�����ց��� o��Z�	�Bm"2���.�t5�0��<7�,d.,tWus|.����^g@�d��
�e�;�4��tE(��wP_vh�stN܅�oh%G%Z9uⰳM���]F�ӵZ������I)Xwc��R.d�ָ�Fk���cBɕ3wA�45̀�K:Xwd���9���0G�=�*ח�{��e�Z�Jl
5��oʒ/M�+�8�9��ܴ4�?%s�(��A�w�5B��Jpq���dY�)�6�x>�gn7.��uH8� �m�OU7��t�h
n"s�-�2���wi ��8Φ���d���<�6Y��\k�$��w=ݾӔ�s��mot�$9��u��%
�tڜ�n���楷kq�l< ����,s��"{��}�թ�:���SC��s�c���[C&�3y�X�;.�)��5��d�so�Z�r�XC�y'b�Nl
��Y]z�,��%��g�9�m�vY4H5��6��F�ל���4�2�	I���ͧ]�ɷ�V��G�:@�!���t���%�n��H��m��nZۨZ��X�f�^�9�D0&U�b��k���mp����2�Y��uV,R33~�fZ3�m��k3QӮ�X�O�]�X�i/49��G��}�0�q
�L��ӏ��W��t�aۥhJV��E`D���'c魼��r,�n9S���)��櫜�sxh�R���.��h[)�dX��nb��^��d���6ĹIXv�+����F.�I���oVK=�>瀖�M�`�X9C�6��xw{��Q�B����F�|S���cC�~����7�YҺ��b��hM���L3%Ք�'�yJ����Cruru�bYq�Η��65�y�؅���f����]�/9U\y[i^��z�-WL��o��56P�O�z�*����2��i��K����0�WxiH����y��3�������>�]ӗ�����J�<���.���7D���y��cJ�݋q��C����͝�lvG7;U�2�"�*��G7X�On�l2��r�f?����Q�(%*�A:��9���#b���>K7v��{`���u�z֕/��t�w�4��~�eI�D�ߜ2�7[�A���B\�!�z^�\��s�!�x�m跊�K�ݱ{��Kܑ�P,�)�mɵ� �_}����P�^�ᕰ��ѱzK��a�Ă�ŁeV�����=�H�����=钦�湵*Rf7o9z.�`wx�Or���,J�������0�3�YA3n΢�bH�z����y%G���#N^K��P�]vh����)`��B���B]LB!�]qh�g�dM7�A�\ݥ ����n6�gq�K$϶�l;}����4�a���V*ӌhoS땻ú�^#��VL�xl��8V���gѫ���^�;&]҂R�`+��z��87��q>(M��:��/�_9T��X��S ��UHEEU�N���K��J��y��	��[�L�[+%��m��9�ؒT��PZ�e[��%tz��2��A;�z�"Z��m��Y!�;m��e��)L謘��"���k���}�;=��y�QT�԰�6T�1�	e�������CKoU!͡|�_U�n.gn�f\����ˁ|"� �X.�P�&_=0ޜr�آSoǽ.��L�R�]cv9�@��Ͳ�T�mrJU�ghS�ew���}��}q���ܶG�&tE�wt��sJ�f��V,3X}]�0�H2Cɳ&pGw�k隌��UNSx#Ț`HYy��,�l��bK-i{Fn�8�r�+a̛9U�ajmg'���T%C
���V���2�ژ{�-r��Cr���J�b7�T�U���,4ˬc�׫.�ĭ&���w]Z���zˌ�f�OTa���m��Ϧ�#�jb��xN��0T����Ԅ_��`$�y*�U��=�{�F�0��I�J@���3��먹wͽ׫���̋Z���4%!�ѽ�[�+��$��|��ӧ�6Z��Z�-�]#�1���8+^A}��2̘g�E;;�V��V�:�y1����3GY�x��l��+�+��gz-�Ӣ�1���v+ڽ�41�x���WS�^WU�͝;%��7Z]�%un������������m��46.ՙ��ݙ2�X�(ځM!ٻ3L�!���(q������z1�Wn.�Y3��,���%�ҐU��E��[��.ڮ�iu�m�u�fM�"}۔Rf*TF�zP�U�����ܢ�_wM� @�`+0���p7�$�ꕽ���h�|����X��Z�V)���s��]�)h�F��gT�׸ 
$.8��XD���};��N.��r�Kڄm��;-���q�h]���K��ػ�%M��V�Y���t^\3s^k�!��L�ݩP�x)��8{fM��6�z��9�Rv�h��08�c�A��]�kq!j�M�t6::�9�s�����}Z����񱎴k��_�ۛ�-q��+���K����zWs�xn#¡���(�8֌u㧷a��E���7C.͎��]x#uc꼮����yFp	E�K��W�&��K�ח�����j㾡4���!׼v�`�fj@�t[����f�SO;�FNJ��/i�Q�ʗ������ʚ������+iK�Ɯ��B�dLJ3��r�m��	]�J���G;k�����0L���@haQ)�N�km�c�Jރ�I���7"�*Vt���z���3TT�
e�B�ocz��V�īW��� �L��[,ǈX�-��5�l�9�c�հvQ�7pf�λ��A��48v@�J�T���;n:��SF��.z���vq�8*��̮�I��,*ŀ�UlW*�*��~���yQn���n�ܡّI.L;�E:֘�U��ޓ�4eћxD��Ri�7��d�B���q�n�ǽf�4j��s�j�$oG(n[�JJ��y9�M4�(i�в��A|+a1�9y´���Y�x^^�Jn�*��@ e�kE��_^�Q�y��h��������x� ��sS7S�fТ�WN����u�:ea8�M�(�^��	���S�V%nu�{�Υ��:Aa{ƴg4���������Hۙ���К�3g;�;v�t�|�=]�yj��	V�;�# 8�A���O��zf�鬻�8u������7jA����9�$�����*%i���,����u��[ʑ��[��pU���@Cg;Q�ve#��Jd:�Sb����D���>�X��G�/2;�9��t�c����eG���|����h2� ;� ԟu�������gm7�����^j�~�T�_Hx:�۴3��)���Ww�`��X784�=6lB��YV�k�s"� �ɥ���W����}u	=Cv�;JVѰʁ�Xu�E��>�?_ƅT���k8V�Ef���m++3AK�@�B�㛦l��]3��rmbW�|@��w�WhdV�u&{� n��m�wW����m��HV��3�L��!�od�}�(^ dVH�"+0]vi���-�sɦ�TU�;\�ehf��v��IZ��AS:y<�_=�t+{*����x�Y&�p���h�cqG�Q(��\�EV�yN��[J���X�ra�39��$�9�S�b�/����}j�ereQ;�*Ӊ�җ���UuÀK���]p�AKx[�3u^b�\胁�{�-�]/�\�٬;6��9Ysa�bG�&^Ye�Vy��v"WY2�ܰ��l�7Q��5��O)��剓�9}�x�A�.i�P+��Ep�kp��)�_v�r=ֺ}�s5}�*͹V�j�U�Z�
wXo��͟9��YD��g]�<��-�ۢ�Ű�P�Eq����-]�m��䙓7�ԝS6����U��#�o�C:.��#��n0�<��Ț������p{����)d�j'���P'�	�w7��͡��㡷��v%��Kgo(%��j���ժ������j֡�e���/���T]ƴvq��\,��,�+�7M��*��1P��#�JE�Ơ���:�i�@z��]v2o�+bҋ�D�4�=���^��s��AWZ�r��0�p�h�֦��ബXѴ��pY��n���|�9��C��������R��\����ɃM�*{hl���wzJx`\���h��	��m��<�}����)`�/�HKk��J�#n_�$�̣u7RDN5��2�f��w7����w�89���)앹66�oG1�X�2¾Õ���sWES�����`��h��h��P�3�W:═�;RF�>���N�Mct�=[��^F���h�i��G��
����\9 �O����þ��֥�Y��פg�ٕ�����qX���j�9U��`�����ܒ�$K#k2�=�:���W�%sdtZWwn?�W==kZ���]�L�e*�YK �X��3d��Yɦ^����HI���m]�HO1	w[��p4�����B_-E_=�k�O��Q���ǭ�;����KFm�pX�N��{�{.�g-�Y�2uڋ�}��ٵS�С���R�"S��H֕+�s?��si�1s�O5k�w_�4�J�n�"�ܭ��^�[��-��VS�����I�Q�z>�0��R�a����M<�tvޫ�/U���`�7Jft��P锏Tj�m���6$�\�n_���  I+�o�;�|Y��,j�r�cW�V{=��g�����y��s���@�@w�vxv�M1	# p��d2�jAH$5I�P�L��-;��|��&6���
@��i!@�YN�"E����&�c��B�-p��>�^����辋��x��b�~��kwi���OZc����y҂wX�q��96i����^�@�H������wY�.�Un_	I-}�8�X�}5|�8ȕG���6$���'�-v^g(�H��cn0�]&�3�#��,O/)s�I���{1�]�G��Y����e,L�*��c2�PQ���2�WM��J�Y����GC��kZoH�v6�ww��:1�Y�/3!�n>�s�Q��薎qn�[c ���g
Zڹ�\Y��6�o��yC_T�Y��'�p�ڶ)y�Yr_v,	��A�/;[ި��龮��Z�Av��U��)�m\�i�&�U*7���e�v����;�`�k|֠K���E�ҹ,�vj��Hn�ΑKJ42�X�V-�ĉ�WeT��Xt�SdW������}� �ᣦ��/W7ګ��$����]��M�>���M֏t�񻶘�:�{4�u���gW
�M��	Pk��˙tڪ斮����$�:�`�c�/^h�Y��}�	P,xu��^�2䜙��T󶄗�EI�����w�.��z����.AY#�e�c*�Z�+����1�]p7}K2�n�Ѕc:��{H�"C1������)���e�M���]��׹Nd܃�.���KgK��&\�u��� ¥�h�K�1�bI���"Q��D�%#
�YS�������dDNO��P!��eF��U@�&� ,'�b$'���q6�?Lb�fdhH�r5P@A��.'*b&�s�y�y�^��O���2��	�"�) y�!���suӉ	�c@��Q02坺11A$ĉL`L����D"!&.u�$L�:0˻���K"Fe	wqC(Q"�(�i�I��\�͌�8�
	"�d����iݺ����	�0��R`�(�]���M)��FQ�9��Q$�$� H��&K!�Ɇ16RfA!(@a��PI� �E��#��Ja�$Ě!Fh�S$2MLR�t$��w2MN�`�Pd�����Xar]�$CII�Qe0�4444��FK	�H�d��0"e9�%���������q��y�]�z�?V#��<bpt�:����:�GkM�a��B)�i�x6wR�NMv�Wi���Wub����o"��N�n��w��c�)�JbI ��a�c1�����e��WH�\��*?"��w_���"�}*N94�w����im�{�O*˘nOv��=�%w��/�4��\��4�>̚3�]�x�<���[7}�P��N='j;�/�+�*��+>.VP���Gu��@�e�5Q���L_z�_u7Ӵs�G��ZȞ=y�U][�'���k��pPV�ޖ=�k|.���o�nL^�t��|c{k^�d���]�=����Fz����Fy��'�^3������#c��gwOHa��� �mlF�n-���iv;�+��{wgx�2W��]{k��g�v�B�#Qά9ϲ<߽��';�V���(o��flS�sܧ�w��w~��χQp��Mf}d��g����7�euwޫ�]y@�@�������=&���iV�X4M�Z��ܳ���A�X�#M�8��ƛ��6�?�/�x��>n��Na9۔�T(饍���K��h�D2�':�a����T©�`�b��R5zAf�s��÷��8+{������2�h�!�9���59M��Ӎ7MLV���^
��P�N[V�LAn�h�������C��k-NR���Mu�`�4�fҎ�^Cj[K�L��%:����.�_���>�a�K�.,�����݂3nOG`���ݻ�/��Yʜ��>k&{��z1�~d�e�����>�͍$���@���Ǘ٪�Ꙟ��SB�59�T!]�w���=Xϋ��r�Vяx�� �x��^�8��Tȱ�E{�^��y\v��/Z�2+"紑�a�v{�{��f�vʦi�ɯ�j���k�<�LO�M�(��K��4tY;����2q���':��HjD��oo2&_�=�t��^��ĸ{�\~�m�-�t�{"业�V�u��{qהM�U7���{miS7����o�> kޛg�Z�l˄\��^>�z��>�19,zJ^�U����pt��p���R�����B�ާ��A�����ׂ����$�/1�cT�~݃��8�"��^�n7��K���K	j�w�v��ɥ�Y������sKǦ��%p'(��gzf���{t���kM$4 ��R�a�'�Owy�G.�nإU[͉k��K�۽���ݞ�u��J�sib��K�FXB�J�
]���8"��stjNC��X�b+�66��2pwWu��6�����Tʞ�K��>~��o���{s�V�_�*�pܽ=��-};�^�O(,��:��y���i���y�=�1���z��G���:h�҇�s�υyͬz�rl߄��S�s\�����A�|}��}}���7k��n�/�<�9���v���|����^�@A���SӶK�lD���w��`��`:��~�NįL��'.p�&Z����/���������6I�c�hqn��1��=!�]��5�P���s�\ɻcï�͉s�<^���t�t�Rl��˙RA�ES�xD��=��)E#��Hm���Ga?v>F&��Q��׼}K��;�J:�1jV^[��wD�<��m���eJ�'Ӿ�:�X�����r�V^�\6�#^y�.�=��r����]%{��~+��ī��?&e���Lqf9�F*�Y��p�G�w'�%k��H�8�o-yˬm*�/۔OV<>���^��-�u�6Z!�^U��x�8�DZ��O;N�%���c�F�Y1D�e�b�˸)�}�E:�{�_���4"��R�ў��:�㖹;���ָ<�-�s:�zo�����g���v���8@�22r��G[iY��^C�o.�S��:;f	�M����Ng�l�p�t��%�k5��#�5,A�x1[� k�k�W�0(�x�T��ܷ/<a�5�����7�$~�����ʸ:�>�X\�O}�t�w�T��<��˷�%='��C�ln{�*���v	^{�9S�����Li��:�,�����df�$�;��ѧo�)c��g�t}����k���!ֳ��H���<�s?I7�o�"(n`��G��oG�|=~;R��/A}��#3��I��~�ⲫ���n���'�t��8Ss��p�fvWo!䈳���F��{A����=�=�v��g���uʆx��v���7�`�G���+k~j=���CW�傩�{��O�;�aY��kO��f�/{���Z�_r�&�X~jPP5Pp&e��Lt�!��]��k����k�+����u���YC���2�dm!pta�'��=�Ҏ�/�b'(;��h�&X��y��&�!2-�Y.������qWFw���������Y���v��Yk=8�䫶�}�+G VV�=�vi��gJ�2Rr�z�nx�Ю]��ʟ��6}�����,@���eNEzY�=�4�ܺ��xp^��<I�����9�@�q])��3�R��ާ���r�q��y�g%��{:Y�s�H��=dw# =��*�����uz��hʵ�v"ko:��� �隗��71rw���aM���OK��L��im�S�X���F��4��}��pFC���&�cdk�9��]��։��=.�M�2+~�ű���U"�	�´�k�xs��I˃BV�T�OP���˃�=c�u����W�탩V�U���l����e��D=���4��1�~���Z���ڤ�T��y�*N��}�o�ѐ��G�0]ztN_��3���z�G]�ok�6o�HX������b�U�^�D��[�Y�l{w��5�3�崪ڎ�M+2��귌�y�6� i��g*!2��G��ڏ�6�Ʃ��Cq(��UطY#J7��1�)홊K��s����-7LA2б�K�ź����em��j��&�������Jx�{<���Y-2+�����	�'K�v���;�*�׎Q�]�7%x�J�Y�=��A6*�q4��s~Ӿok�^�tHq������v�K���v����@֯���*�������yR�9�v��讎�$��q'�M�`F���i��Z��c�=�o�y�1OZ��=�Y}�*Ȣ�ò�N�y�Gs	��X��*^7�]��U�A��66���V��o�QQ�L��yc��@���3�)����j�5�Ѻ���k�m��D���=+����F2���5�c�1��S=���{j�<z�m��y��ş��/�7���>�Ѻ��פ�|�xB+ۢ�<�w����kӯҷ3�^Wݞ��s�Y#���;2n�G��fO]�(��u��_^�����uˬ�M?^�e�Ɉ�V�{�o���]�IOk*9.](���=^v�s�ɝ�1�áFw�أ�7�i�	ap�I�ү5R��a��NN��u�(43�*fi�����O�d?>�]1M��+�No�]�j�*���-��&�Fm�.[M���n��U�܉)�|^���q�(	wZ���j�f�c�_�U,�z��$v��4歬�qb�"���~zz��{wף�i>�Y�~]:Wyv8uؓ&��5A����[LM4��+=I�OY��������4_I~�n�2�q�}z^ٿOOA��y�R�����I��5.��>碟���[\��g��O4$k�M����zƳm�Y��'���q>��Ͼ�J�����������0�铧���O��0�$_�����uF����g
�(���}9}�`0m��� �U=:�?2k��ߏ�] ��Ӭi{�'�9�]xm�`s!��6��o@�_��rn�uo����^-�q���&s��8|}�\��w�SR���6��U��P���F"��"�/\^��Q����cڶ�T�zhy��Ý���<%Fp�c;Պ�=��t�����h-� ��:,���]����w[]$}��줡Pi������}��h�gfG+���4��Bp��֟S�'L�6�H���N�������=
x&H�^�w�ڬ�:���J'�=/8;$w�}���N�P;h��g.�lBM���a�y����g�H�'jξ�9J��׶��%7r-���tV|3܍R�<�7UӦo�l��.g�A�Q����fJ'�piҢ��\|R�-U���=�_c�bl�Q�[�S-p<�;�uj���Gu�ry���K`
<߫�Y>�4�4�//z�d�|6�{��S��oW{����\���߲�٩����ɨ�%���I�&��^�����)�U^�OvM�j�3��D�W^�G�_�u��~�F�7����=�[���&�5�g�NU�٧2*�do^�ʊ�:�ٗp��sA��
���Y��{��;����F��}�j�ڎ�"�o����y�5�4o?b��Khd�%{�\���oڙ^���������ye�\<zG.f�Э{���㏬FVT�uGG��#Ѽ6}7�hv�V�1`샱�C�5:^�r�_zLK�i�v�z��A����z�����=�5��C��r;ޤ��eq�l�Ç7%�2SS��pǮ�����m婊3p�E��Ƿ������pxy[��
W�\��o�=t/P	�.�Zoy�z��l� X�H�,�JU �'~��.�R�ED�Wq�0!Mo'ƍK)��ۗ��ξ멼�2ͫ!gxP�ӛ8���l'������ܟ{��}�}�+`�T�+ڏ���a�-]Ysm���ܬ�"갹��:E�d�]�����Ţ\5�|�1mīG����5��_�[���5S���k��ڨh	�ģ���z�I�}nf������S��^
�MG�ޒ��y�U�y��E��m+��ϳ��|��'��׬�<<W�<�YZ����u�ˢA�\�\h�>U6�2jo���K��˲�e>���a��ʜ�+��9=�\{#�`�ُ���͡޸�(��_X�Mt�X�ǅsW~����
Y�.���uw�x��v}xH�$W�ƈ�Ұ��^�{b���U���ǘxy=�I������g+�7;^����v�3�n�z;�L��#Oq=����D�|��:Kc������k&6u���� ߷������4�������2�
e�G�4�X&=�J�Y���w�\�3)��%J�k�r]b�ð�^ţ-*B�3��Zѯ�r�廭��&���NG��
��$�$����gj��y[��:��ƠN�,jy���Z��5n�zyZ;Ҍ�f��[OM�*�c��"���=Zvu�=^���/j�)�_��<�P�G��yv�%�g�e1��^�\+�Wۇ����+�h�w�}�-1
عX}����Ա��=3-�{c��OK�Pr��xNH���\o1��g�xi���g�ζ���Sr)xxd�rf���-���;:��NM�I�-^����(�{Ot�/�0ܗ�!��a�W��U]v�>+�ȳ8��6*�8�=��ni�|�׸�ۛ�i.�J��E�&���=`�s���\���,�7ݚ�tF�ɹ��9\{��}��3徘B��\c�Qڞ�o���ƍ(xo?��0��ϲ��_.���iR���ߗ���a���g2�M�o���";�7X��G3���<e��ɩ�r	 ɉ��N��9Kx/l�2���s���+�m��gs��^�o����x�=��g����x������n�`�j�0��[w�M��>uGY�E�7�]�,���f^I���7YhoE�WS��38@{Rї��� {�p��ku�y�d"�d�H6�U��M�rW�N%�r�c������x�j*��S�k@2��$�C�IL[����n�*p�-_�(fܼ��?f!�0"���ê��Yp�^l�u��Ve6�XNn��%Am&������e:�[w�­����:�ݼS�hl�����ۭ]�����
Y)3�FI�Ӷ���ZCҩc���K�ݖ�U�whM��4ﵵk*�Dj�1����K�f���P��7PAKh��z��݌�ݱJ����g,��v���],�A�[�m����U��HV�p�s!P���{Q�uB[���H�n\[ZdIV�S�WSE������j�6wg�'�l%�L�Ֆ���]&�hޅ�V�q=�Y�`ۙ[\$=w77��X��$�f��]����{�B�M�j����; VQΆ�8w��-��,bF3h��l^?���\�;�z�"f�9�Vֲ������F��؂ٙcu�I���2�-S�d.�]g8պK2mn�:���gS1��+�kNx��O.r-r�ӕB%�b�����.��-<��%e-P8��99�v�6U]�<�T��@�Tp���s�~�)��Ʊ�,ѳ����S�a�k8
��Y�i0r���ݼ����R�Ph�V��<1��py�N�hM`�%Y=���&�J�,�X I���깁�ҕԃf����d�l L��*ԍ�Ɣ:�Z�Nf`$�NgT����$���͜��c�{�c��-���v/�ǃ����i���0�jQ�t��!l:�1�� �Lǖu��G-��e�m�@�B�������u��Bd|�in�3B{c����l���ڬk�i���٘Z�V �Iu�m^��:�8:"4}��:�s:��݋��T3^�%`�My���i�$֮/z�"G��W��V4�n�@��{��E�Lۻ6eL��]�:]e��I+c�:Y�O�[�]�A_���I�&<Xp�ŧ�뙭��A�X��=v�֫9���V��p���3�k9IC����26Η�.�zb�yD�u#>�}�y�����`�:�vM',N�˞�L�X�#�eu'D>w�c��RS�s{}������t����X��[������e���-�>�:��CK̳J̙�*.�PAm���éݓmN�f�e��I�Ya��m�Q�-��b3Qc��Ʀv��$�R)��\��Y����N��R8뀝�\*�6�j��R�H`�m��.��I"v��!;pƻ�.Ɍ���[�]�]*c�˰+�!L[�2�2E�P�wۮg)p��:B��V\.�,&���!�&���oWmA�t$/kW�e����j�D̕�lm���� �j�8/��e^;���{nB�]�,7r�r��r�6�뫚�78
����v�}��s����~$�I�idѡ3r�HRbH��JB2D�dL�Qs�幃LI���$�p�wur�D�B(����Iӑ&�FFN���$�$@hLMGu�F0X��t�CIE��!Π�!ݸ��I6�0��K���q$Jp��Q"����(�w"��Er��I�ܺb��dba�v��I$��h�M&!��<�ܮ;�λ�//$C$��1�&�s�;����t���I]�k�s7�ۀTH��5��1��3��ǁ�wM�s�����<�]x0O;���wuٓAd�:��y�ѽw��C79�0βwL�p"��30�<t���<��˼��T���N�4�Nnɹt7���;:F�tus��ݜ�xl�<I���r�B]�uqr��ו� �+�^g�t:��<��^m�t�"����w[�����$�`O����Hx���i݆�nx�/j�'z�mn;Q��&[WEL�h���)���,M���[Gd䁢��Nح��W�S@��`�� @Q����,�4�mc/\� �S@A{�9�����]C��ܛ��<��9��:�� �C/p�֟C�o=OE��ޑ��73M{�K����oC�ɴ�nw���p�r��̰ ����hܑt�l(~�Lpza�����&Z�}*}9P��
\�3u���*'{��$��ݼ�Cw㉕��v:��m1P��.���
f�$F�W�x�M�鋚~ȗ���2�B��hle����4gXzo[`��x/V��A@���dg�$D��!����R�J]�����g��c!q9�;��[ ��Z�e~U>,����� �t�)���$(����^5�˘��ʥ������v�o���#C�R���N�ሔ�t	bWIje��fǨu�%�1j�/3��mQ�%�E&nd"��*U�/�CDfE�N�F�T�ሤ�g<�oQ�9��s�Ԭ&I�:��jΙ}��^~���@}ͱ���s�ړ��^URa0C�Z~X�A.Z#Zኗw`qb27u�7���{4����#��i�s����u\�u�9W5ل^�7���-�<=�e����i{��$������\K�hV�S#�mG#�r��8����e�GO�����|�����5!$JQ��WsHU�{!�h��6g]d)�ử�n>�k&nK�#�2�)��س%���%��Q���N�R�gq��hÊ_���͗������m��rz	��t��v��v7��h`�����`Ȓ�	c���,��Sp��NI^ūs;G�żtJ����s��^n�3e������C�<����K�Jb�R�(v^F�1�c�Y���	�8���}���ny����:�G�1Chp#�W�ʭy7�3w��J��X�L�ק����Mou{���bX.)����PO�5��w���!N�d�[Or�u�1�v�_��~���62��Y+���	�4]�q�b�L�z�J*�Z�N)�l�ꘌ��X���%��m�1����s������Ѧi��.��b��Bbљ�l�I�Ҭ��W�j��/r�՘%��|�� `0%�k|�eobj����ح`+���K�c�ȫ�}Y}h�q����Hj �:�={6m��l��sӼNI�1�oEWqb�f.��Lݾ����� ��Ƣ��nka�C�+�Y��C��cQ?�*�~5�z��.2��aٱ���/�;�č�æ��Z���-��-T))��[B����5C���)���?;�o6�d�+|���Uos�JY��eӵ̺|۝[�܏*�o��9�]��[�{���8���K����Sӎ���<[��A<�A�sm[ᵝi�5�l�q㱢ܫ��ƞ|�eA��0Al`;ك.]{M<�����_���߾�Z�#K���?k�W~�p^?���}�F�"<%��ŨtBd�����a%"ՉTS�oP�:��W�6DVB�s��6�0B�[B�8ށ#�cH�(8��2���=��4�R�ȳ��?�3)�`�]�
e����P�fwrn��PO�E��-ᄉѓ!�A֑�pNc�^ˈdA�P�5)*X�^��i�j}[�r��m�"��fۋ���1sO���z�3�Ϝ=�-y�!����Rrޝl�N�V�K����=�XjV���~�6�憫7(�����%<;�n;�lm�0t�ވ�h�݈���&ѽBZ��v)>؞�o�Ĝqw�QaB�O2�S�4'��C��>��U�|�\�.DJ��(e
`���ƽ=#�k8еn�c��2�Z�⠗��A.)u��-�ﱫnoʪ��J�Ⱦš�W�#�Ά�i��\קe�ol����aJ��˦��;N?��!�w�z����¾9�����R�e�ȗ~��t���Ӓ쓫ޗn;�[�Et�bp���]A[�nz�[���ؿy�p{C���Ey`�_��u��->0�s���<L�aW�ܵ&�|�KGv}��{$��nԯ+��b��x�9Y+pz�w�p~�����U���2W�u��g��Z�g	��}�dG&�+h����@��%-�-��]j/��u1x�J<BUz-egdrk�B�ƅ5<�ܔ��{�ԝ�-ˮ�V�Z�\��{���صۻ�B���>݌��B�P$=��B&a�l��n%��fq�_��Sl'/��_/ӏ���U��z=f����@�j�"gͷN��b��tS;yf��Z2z2�DI���Y{�s��B<Df��s\��ƥyU-�y@Z�(�B�����=�6�x�2�Am|QW���.�4�9F)�<Dkc`��v��vq����殂$�|�#�O�D�8�
ze�ᄼ7�";z􂷧5�Z�ہzmAĐ�B`$�n����O5t!)�y��c�%��{s��S��b6s[m�>��y�$8X��|�x'�g7�s;K滙י�Y���������Y'X9��(�oמp�Q	�k�D��"!0\�Z���+s�3}��1^�'hZ��6b�ɓ�R��n�c^������� �^<��{T��C�E��5�í^�L��(Bc^�>�H��'qUeWC�ȴ����t(~d�8uX0T�h6�Q���Ѓ�a���,�X��E���	��I�V���&F뷛�2�ni��.���'�éd`�2�to�Q��x�M��#�-��]��ͬ��mR�9!�lg ����tf�+�~5��Y]T��@6M�&��եsmt�����L���Y{OtaI�K�=M�1�nK��x�k�i&d�G��5x��z�_�����X�e�.���8�����8�#�:=k�	٦�%���6�r�k�|���1[���s5Wh�R_%~���Ͽ]�v���@A_p���T!�]0#a�1�nt�&�oR1^۱��#v������������ݖkϴ�W�����'����|�E'���~٦z��V��#��vk�p��B̆�>�)V�~c��ŠvW���-�C�C��zA�xf4�b�s?1�jݺ�M|��'u�o�S�=����|M3�X�K�( �S@BYRŴ[�=���j�s5�u.�ە6�w+g@����8�՞��Nv~�~��C���Q2�d�A,��#&;{���1��Ч�ݭE�pô��4S�"�� ����g��s�}�8Թ*f�ftޙ樦8�I�����X`�O��Yio�?R{���S��a�y��O
��	XڊL0�o�ޙ�9���]�z��� vTpb�b�N��o��z�o�[�y'K�&|��p�T�r{��~�^��M^1'8Ĳ.��dB�Hݷְ�ܬ��)�+J!����\������=����a4Onm��z���9=�VseY}��ޣk=��wiD���$��DM�DCeK�[�J��z��s^�&^��KpϵK8�[Ke�eJ͔����͊.k�[ �r�4:���,n�&j^��+�����Sr2�TE}������[^-]/ͽ/������H�K�DJt�����O�1�Q�����"��{!P�4P�N�������/!�ᛙ�C7`��ha�`��	�`�J�| �Rr�sȣ^�\Ø�Ɍ��z�]>�,�\�7�\�muR�����-�y z�M����}�6�_
�n�	��(����p��/K�OL2�y���1o!���y�"bXF���!�c>#����#��V:�Q�ί�_?<i�s˕�fF�fiڥ���kt=�@~X��&��ׅ�jd.� h�]�B��{1ss4�DC	Sn�e��w!,P�ʶ�L��،yUAUK6kӻ6�b[üC�p'q�y���,i������x�r����:��^cYc��V�y�A}�����=ڭ��f���D���rI�Щ��c!�ƻ��h?VI�İ\SH;IE���:`5����,�F��Sy'p����#Y�<��i���lmH�o%�A��L%ڽ�iذ�=3L�0E�a����e筡�u�|�R���$���h��"`�\��m���>��4�9��3�-���f�z����B�:NP�q��}/��$0B�K��f�.}U�-XOm�7���A��%�~�&�J&��l��Z76�����Ryf�U2������M+��9�+��8I�s���NQ�:T�v��+�_t\�﹚�]�����c�ݤ�w�����u'�62����41�B�)\�k��OM�^�f�����m��ȧx�`L��2.#���\��}v�Q�1~����Χ��2=_�¼B���!���z͛e�)�?4����������q�-�ug���������l�B~c��r���T��Yܰ���ʨ��B�$����)�m9߶����VX��B"u�T�����3�l1���2׾QIՅ��+�,)��[yI�u�`�LpW�^1]^��g���Cd��SzB�k�t��r]�H��ŨtBd��c� R�@�UO��p�|�eG���_�B[\7��~��'�v_P��<�� ˲�m�a�iޥI�z&n!�m��g �kymů"��q&���˳e<0�ǡ�O�'�^�ɽ�+:�*�����W�C!�S��c��"��摋�F׏Ms�w�D_���H��ew��t�-��=��؀���O]
��I�P�+��\��̈́���9m;	O�ѹ�!��kyuL1�m�]��m�&���6��b�,���s�Q�bN8�*K�<ʮ�k	Otj��o�U�6����k1�8��v��z���UL��x92VBv���v,`GW�_\�S��S$ݯ�|���2�NZ�u$�2�-�2�JZ8�-�{��_Y͓V�W7�f���$giL-]����Urt'���Z���P�qsc��{3y%5�o�j�g�����{kn��i������`�L�eBzG6�����t�{*	{k����p!�1���i�D��
�[�w2:G�f69��s^��e��E�5aJ��˦����yh^��U�F_7s�X�j[�@��3�%"]�NC��o׵�쓬�.ż�^�c\̳Рm��+mw��';�^�.ܡ���&e�;>�b���J�3��<�S��x*�����G[�[���c�v/"�y= ��8!�&a���e�P��r����f=�Q��ʸ��.�F�w��앯bj/��c��f�A���,��r8R&��q����z������'�d���j<��"�Xe�/�w4���cWXʩlj<�.s��"e
6Up������Q�~ɚ���WW����=|S<�sc`���C��e���mT�5t)���7���a)����+Z帆��h{�����zǫxi��v�[&C�L����CHΧ��@��暆ͼ��/V^�Z׹�K��0L}��o�_q�P����8X��|�pBx���`����k����p�
�����y��y��^ߙ�پ�g���0��?����X���L�L�{ +6�m��J�%Ҿ��֛���$�t��V�=[R-Ȟbu� 0W)|��(��i���4�����o�Sz���P�l˗��v��x ���m��,�5�#�̯N���`/ɼ�`�cEL)�+�5�G�t]x���vZ����˽	�5ߠ�VM�΀��k�*��N�f):ac�J.���Lqt�wx���y�6�qn�o2��[��w]�S!�!���F��= ��S�&̧q&ʮ��E���ƗJ�����tn����e5j#�ALAo�C��-:`|�z���D��+����)������Y�i�Fz�e�l{�P�o��glGc�2�v���5����qDG0>��8u��'f�U��-l��o��͊�?=��d�o{�:�g:���+���;ʈ]�t8s	�����2�I镻�e6:9y{,��R�(Gm&6�:�/�gӏC��5�O���@O0J���Z� ;�Dv�n�*��]��W/X���n�fپ�_�AŜm�������%�Ш�p�_e��e��]��[�c�2��Si�N�k��&�g���
_���hH�CH/��{:ٙ��-ەuM-uYu՘����x�kKO��L�l���^=���X��4�4ru�PK( ����R���T��y���R��u���НHv6�Ø�a5�.���&:�����~��m<���L�j���3|;���E����u�Q�Aވ4�v9oG#5��m"/Fq��{�V�3I;�'��[���_��_-Ў�Y���`ܖ�x�=��W���{�]oYdY�R��M��u��Z��t����x~�x�MO���c:gZ�F���vVq�uv���Z���Z�Vݜa�C���{Ә��V�S�{�k��\zxW�V0I����o8�!�������q���[�ǥMK�{
��:��ݾz���o��P2pD�X��&�*�f0���ۅ�f���{ `^����'�%�{	)�JL����|j�t�On�e��Fr�!�)�z����m�C!�lJvl�%�u7cH"������'�)��ǁF�[X���Z�{⫘�g{��ع�w��C��Ǡs�[ToK6קg�*�,�M�N�tҤ���r��O?�Ȯ�Um��(�k`|���ʘc!{^�#ϲ�-�w��1�cc�u�SIs�K�ل�;)sb�OPSt��g:v��S���d"�����f�D��w���G��B�z��˥Wҏ�|�ʁ���ӑ�=�.jC#KĊR1���%�lw�K�s�;�����<�v��Ԟ�Ax��r�ۯm>��T����SMY�2��X�d�ͫ��
�Y�^�ٷ�����߉i�}������߭������{�}��~��y}4h7�C��EE{��p��jTg �����C����=+�vf@U���}+���F�{g��7�n�ժ�qqK6����JC!Mu-�уX3�J]MMwY�£n�7u��v�Tv")��-�*�4�W�S�-m�T����I��ݲ���2��.Z�4%�N�2gb�G���6X���n�]�Ŭ����g$Wº�^ѫ��$��1h��V-n���+��`�.��c��-ְ�cs,��m�G��p�lm��k��Ja[�g8I�gj��u�%t#	�b��ǔ�2��fV#du��V�ˈ�3�T6��8֊�����n:���̣8`[��m���v��5�Z&��;���W�x�v��3�J�x����XW5���y���SB�Gי}�c�l#�w;�>u��m���7���/�|sqڗJ��)pł���$q\���X+:��;9\��{�KHZ��yݻ�%_K��ۺ�+�	х�Γ���u��uq�f���r}ʔڳ�Fj>H\Vx�}[ԩR=�Mi�-J��Y�.��Z^��(k�ʋk�A>���k:�9���]m�=�w紨�߹�/�$Y�m���u�D�'�`+���ꋠf����h)zj%/��o���Yb�2���Ʃ�%��ò���jμ4�4T��9�Sjc/�\�������F��B����Et���ε�h�Q���j��e�ctӄ��j&��4'e:W���V&��Z>�s8lf�lb=��ٰ�uh#o�Jc�<D��8�2�J?b��][��5��}�!������kshK�xk���I��{A�n�tj[����%u��s�EWyAVk	�_�wҏx�E>��+��c�v3�y��-ڪ�e���nŸ��F�k��0e��Ű�Nԯ3Hx�XyS��0+A�q��Z�Pz�K�=�ָ�3B��a��Tp�s=x�4Un4y�V��!WA�w��X����K�岮J���d�I�P%�:ԭ�t8s8NjC��N��W�fǙ/o�T�֚���ۗ�U�ۄY��z�T;����[x�Dp��w�SmĎ-%���2�@���S�K��܌q-��T�c(q���o�
u�����U�HG]�eZ�&�6
'���x�[�����b�q.C� &���x���'"z����+j0�I��Mɬ�T(Q(��Ӽk���͊,f���zL�p��@��U���MI�;�f�kr���Yy��	��^l۬���>YvHy��Kv�h3��2��i0�Y�M�Eo7�/s$9��g�d��A�����h[@)��Mĥ����P$)����[+5��S�/�6��V�YN�2=lm�A	��Ѻ�Y͢�2+S���+��z��vF����q���9�y�I�Ȕ�UF��[�.��,KV��^�5�А���,�;h���(|	�i������`�9�[��R:c-&'9��ty�����e�;�e��K����3~<����])$d"o;��[�����yy'w�9�aI,���x�]�R�x񼓮�c��'v�D&�ȉy��k�$Sws(�����n\�ݗv�.��i(����t����/uݏ���<s��޼����9$n;�:�7'Qt�
=;d����]��y�QwrhȚ����W����� �f9./:�$�F�cw�;�=y�^�\NS�\��&����:�^�M;�8h6�lIdb#;�(��$�����v�D���Xf��k�û�Ǟ\�ȋҸc.F�\�"��bNnx�6y׫˷��6�L�$�p�'u=v�lF"�lZ3��Xآɹ\��eAWw[�7�颍m�9�a1�sG�?��0aB�`M���O[�ts]�`�>w3�m��n�l��U�K������ٙ��VV<n= nI��=���b(t@�60A�7sbߍՁ�Zi��l��N5#��Q����}�*��~������u4����?�H�Y���~}��Bպ�ë�cYc��������j��}�CX.iI��é{_��ƺҹ�d�A��W|��C��c\wU	�ym�P]_4���`�h��E7��`ʌ�,(���o���c��C��VS+�_�40-10���vF�V;�7<�gX�bK��"i�w�Q����)�q�|=��YVFÃ��y��["]�Ѣ���u�Ӎ��;�Ǆ-���Scao[F��:7���I�S^�jM���m�ƴ��6�kdS��B1�y�-�{����YX8�&n�c��ƐΊ�Z�rd�VIE�|ئZ2����N��;�%k��V�)��g����X=�]�(o^�V6�@n;'�,�,J��r�Om�ʋ�7J9hvX�n��]�vx�e�c��5��T�F�\����T9���{��Z�B��U<���]���~<�&��d��5�B�[Q��1����9�k�K�Nչ.�$�L[��$�D�0���ա*oz��V-�C�NWs������z1��A�>�H8�2�vK�1{r������u,�+���9Ym�>v�1a�·�R�v�ۻN	9N���޺�m{1b'���'�D�eS�8v�=s&�3mK��ޝc5/���q�g{Tcݚ9��,K��1��iN�r_1����î����W�5Ul
����0͎ܾ�W=Nu8u���������{��wM�?J��{#�5����h_J�@�E�|��1�� �cO��O�����kyi��A�����-=ۨS7v���IO6)�E�.9�b摴�z���!��@A��UCK�l+�b�4�B{:�Ph�y/�I���i0��+��B/<�ǖ˰О٣r��g宖S�ݚ�E]
S�3耛Sק����D�qG��t�*�U�$'�����\:��]ѫ�z��qán3�r�|���L	�yQ�[�J�}~u+u��Z�9/L��W&8`ӂ�Zb�q݊���,�9�;�0G�4��i���קe�m�,9��R�v�>�#��V�y��*�j�t7��9L76��e���h�D��.C���L��\�$�Z]��6�b����sS1]�E�)�G���^�H�������������24FJ���[&b�
Ƈ7��)��u�m���#בh<����� ҉�c��{�mᎸf��e��h�7���������R�1[U�k�4�������W��諐�&|��.��y�)�ާ���VK7��l��[���i��K��T����J~>��7�����x�z���e��0����jyI;P���y��gx��ڝ$5�ZOM��ܮ�\���v)�-0,���I������᳢��WҮ�`��v`[!�噘5�o.�~��<<� �� �+7���^uݛ&���)�<DsK�^��O��{*���yH\�vd��I�7����~=�G���s?%�u��pC��S��pϰG�A�0~ه���j��C����xtI*a㭺�*m7�ƴ0Ȟz�����;��(���Ǉ;3�Nڏpi���h;��J�e�(�j�A�G1��)�ɔ�ɜEP�����o	������cϡ���Iʋ��OMn]х�]�E�qh+{LBN��K$�=R�5lp�I�>�s���/����q�U ���R�-٢7;�]zLpe�@��i;Ϭ�'L/�J.��)�]N�F9l�8މ{d�5ٻ�Hnt�K�#DC1i4An�'������Q�����Ut=Z�O�iAb��v���h3���߭�?��L{�-���2����%�ɛ`Z���|T�s7a���t�1pb�p��l�
u�׫�"����On;XC�\h#���\�ÿ�I�G��2�w������E��ݞ����;�u�yT_�i�S'?}��]:
��'���7mt���j��ҋ�yڈ!���:/��w.�Z��85�{0��ʛC����K^Boa�5_��+��b�b�He�2vPh���H�h˕�g/�˃��ct�6����_*]л���m�s��k�H�%��uѠ#&����%nS'���wu���M8"t.�������� ���t�ѝϝ��v�6�	Rca�u>XE/_�����j���ɀ�぀�խ;�E�^ܰs��۫'�T�m�{��??Pݐͳ}(���G���&+�C���!�����a(��ۓ�2m��u��y��E��:};Τ�o&�)t(H=���T7a�:�3W�!���j�4�ؤK�dEC�tK<y--$d�F���=��9/{�z�4��4�49o��(x����u�~m�m���$�WQO�ʾ�-3>�
���C���cǄ{����{���o�	CG�b����&�_Zf+ݲC*Y8��Q�Y�i���i���RL`B��(��832z��}ۇwc�0Gm��R��Kϐ)	M��Pd�)��z1���^ ��z��E�K�	��0�%N�0f:�a:���$�5�A8�q�d^�SL�Q��~��|j�=��h�Re��-�C��ݳ9S�8�tB����͔%�*�cH"E���:"S��D�6�E1��&�҅?n�S���M+5ڈٕ,���uF<��kg*�682>�,�O��w��$�E'*��gD1������t�Xj�XB.䦛)ΧR���!�(����U���}/"�/�a�c�r��� ���v����T��2Y3��u�p^KO��~�Qܝ���`r�`��X��y�4&���ZJ��6^�'B�ug���4�kB��m�\��mv�КQ|H�2�}����������f����nY���Ecp��+�Zٚ"j9�R`Ys�}����-�?��M�;<���K�.�{�{��h�0a�n���\�.�lYu��A/^�Z$r1L"�H~���Q��G8�v\�=�C3�.Ʒ3�=����wus]�^-E����y(%��H1.����q�����J㭓�n���u4����
O�'�S�j��L��׉̛z�+�@UR͚��͸66i��yb���o!�Fuưe��p$C�~/Bz�{L�\�L:�Ʋǰ8���Ĝ��5�B��������Mc.���Oj�̺����\0g���G1i��������}8i'Ǚ�
Ǌij���ZA��h�޴ƚ$�Z���o��XHqEM�/�~08�b���i�������7[����ж.���l���7"<{��C=�ߕ�Z~�V?F��i&u~��m�1��@hb�A�e�oy����w6�����	M�H���o�i�m�׶E;ǰ(F0�N�gV~=����畑�Hd~����k\��۠őY$1F1�/&������@@���o{���?۝��J�.�[�CY)�������V��1�lW�ß�O)+��\���̙j��d���k���64��:�W��~n6vK��z���Ы	��p����tmȺ�wXj��s0�vk\p��\a����8���ڶ�ʫlV�ŵ|z������~��_�89�F�f<����P*���������	�,�,s�
��r�Om�Oq]I�ٵn�틮�3P0�6͈�q�1<�>=:ɲs�����(��*�;XɑNϗ��v�kOT�,`Z���Qmu�+�����	�&���4xh���P�'��3����ES��Qwv.��P�bU���ӌ;��oD�#� ���eݒ�C6�^c?n��H��Z�mwv�W��̳��&*��Qz+�q�eٲ�h� ��B~:.����X;Q�Ѡ�wr���Ab�i�R�́�m�t�n���#h��f�~|p��u���AٺI���V���	1E��MУ�S	�2��֮Qy�%%�-�`��ٹ5�d9��"gg0�l�t����g�������yց&�Y�bN8�⨰��<ʮ�k��Y:V�&(�p��z:n��VZ��W���O���1��ͻ�hZ��V8�=um�Jb���ɵ]���j�{e;�(�`�j�;���5�69��sBv]��m���-�����k��?u�|�87�:*J�*�ᶄsJ�ݖ�hX�ؐՒn�.���iC����
�ǫk��5��҈�Ik���&�Gyqm�^���v��wo��E�n�8��F��	�	����Ǉ
m(1��H��o{D��6����f�sV���� |�����f���X�[h�VJ��ϟ��kj��{w߃gMc�(v��q�nc�(����dȗ~���<�DLn?_r�Dt���c�M����Mۉ�K�e���v�a~*%;W��c�LC��D[G�-���˼ ��.�� �R���x��w���ׄ<ۦ�V�fyC��Ht� �3 ��e����Y�ٚ����5m�[���ތ<�1��Z�c2t��5�mc6=�	��f/@���&|�O��<�m1Lya���u]9lj���Ίc�X?~B�ԯ'ەR�˯�B��ve��(�rv��E)�����{��a��Czm��mM��tS:��L&v��k�l����x���Y=���Lq�>��7�+��� sfD�J�h]���z���)흡Ʉ��R��5sq���T�]�A~�^!���L]Lx�Nl%)�j�U�9�}c���={]�0�y��F�]Y��n�W��>)xc׻3�E�^��2��/�:�x�%L8>�s�{���h��J���]�we��"!0���C�"U�N�f):a|�Qu�7E1�]Nݟ��+(E?
����ҭ��gb?��8�Ɨ�g{��Ŵd�����8�G�e8�5��r�툗��x�V/�W`'�z��A�zdhS�z���,��@��.uy��N���|��Qch�=� r��ە���k��E]��m�yko)��� ���F��Km��6�F��[^ff���]��\'mQO,������p��S�n�(��I�Uzʮ��j-?48����8 ����9�Z֎Næ�\K�����=���kH��ѱ%�ɛ`Z��,oRM��f�5�,���Ȇ�؞|?WvOǨ�����[�h&;XA�����4�\�%��U���1�U�C�wjmB;k�_�t�r���uO��ܳmt[���à<]��7���"ʇB�SC�/FC�ǠqM��*�eO�c�o�fy��nY�xņv2l����e>K4Da��y����+^a�>'�N���{vC6Ⱦ�_�1�I\Zeb�>:"رܛ�;D�e��uk���c

VĀ�C�A�8�"L�{���K �Xw���
^�BA��B�m�l�XH��w��xg2�6�
!�hdK<X4���P�-"_�� (7K�Mx�����o��k�x���0�72�)0��^M���-3�U�Ś�??�<yK�?�#�n	��S�A��;��q��ޖmo#��%�lh(���6����W0�p��4`t^��R�juU��UP�!U��Q�63�SNk�w��^� i����ӧJv����UJh��݊.�i�:�6�ɦv�V�.f�S���)V/��d�`�x�d��9K���%��!K��b�r��흙1,KmK�_�-������~�W�Ui5��Fڱ�Y5Q�RmV-Z���}�}?{�-N�e�2s&)�Va��Ic�������j+�7���~�(2jX���UӬ}霁��xg�������C=�iςg�;��l��j��ezdw�͐�d�殈A8�8Ĳ/`�4��Mn�Ol�.1�`�T����;T���s�2Aa]�!��\3A��%��)�r�	�]"��%:o_%lݞu�'�v)b�ѷ)��.�ã� �5���m����3�Y��'�z�$�Vvt�U&�����1��p�^1{^Eu5�9�=�����R?�^�݇����K5�T�:�s.B�W�i���ټ���a�����R	z�A����Q{�]4!4�}�x�k �غ�|������g.���O��E��5߱J/-H�0�䣹�>;���y��b�+�<��_X�<z{�$%w"J��!��*U
.l	2)�A5mw�2��_�-�i��|�a�/��ͦ��ݰ����i�&�=���ȇm~O@OC���Bպ�é�k,{z}[bLW1=p��+�5�Hv�ϻ�}����A��̂�A�</Ҙ�C�az��O�;M�2��Y�
<�`z�w{T�3Ku�
����;���ZH�k&wVO����	B���VD���K50,�J>5^�O����=]�����Ui�6�!ѧ��*���o�9�u�#�]�Ø�4U+%L֥͙�y��C�!M�[�ٍ5ݳ�|sq۞? ^S�{�ߌ<��=EY�Q[R��d�Q[f�Ƶ4�Elmi�� <��3{����{y]�e}��V~{r+Z���,Z���xg��9��'-q0�����J�u�HnXt�pW�fe���BU��G�4|t{��hU圥��I�� ��	:�N8𭦧�Ȼe�Gon/�c���3M�]��e�ډ�kljO�r���킒c����Kz�V~�����;���lq�j=:�b��v�A�x� Ũ�CQFu�6+|��Ξ9�u%[W蘚7�[�+�;�P:pB�C�=06=5����j�B~c��s�%������ݞfX�*���=�\�	B�����me�M�Ø�a��e�#>��Y5���D �_��uS�&g:�\���Y��b�gK v��T\9��|��
�]K�N՛��\���͆}��z�k*�FZ쾲[)׶"y�JE#�TP-�-�ȶ�э�DcL:A�����5��rr!�_�p��K�ǾvA��!���4�g��LU�y^��@؎�.͔��ƌ�!���,E1~y�L�v�B�����{�C2�����jRy�Sl�����0���t�T��@�����g���x�}��o�����|�DMe[�T؇|��$7�7G��,GPӡ�3{:�s���d�Ւ�7��A���A3�� ��r�"k1�m���s������o�"����U�S2�ȴ�F���
	�`�zn�[�[5ي��뿱�"��)�X�N�)r�'�7��j�%�Ӵ�o��)/�-��(���ۍΙ�r��\�8�5��=��V�o-��ը�ŻzX���9��Cy��s§.A��&�tnف�|�|�_\3�:��|I�jN�[7+w��%A �S�%Z|c�:,�����w�V=F5n�U��m����B
�N���Y͕�&���[0:�)n��oT��':]a}���-�=},�o���u.-�eE�ne��}�@�ż%ܱ�Nb��ǚ^.s���4l[܎�oN�Mf5@�]/���
�/�t\����x�Žy]m
d\m�2��k{�u�ͷ���\8�� s.�U	�n��}'����9\����LY �O���凼�M�mK��B�IL��r�Ѵ|2s ,�*��`�G�E1���^,$7�1����p)CJ��]�A�ݖ$�;��UB�]<n����b��]�T����
j3}|ѡ]]��ݤ4aq�}[=݀Ռxl�ʩ�O�cw8�cRfp^�*|DS.\=���}F�F]��\ז.��Y��JHUbY�RUE!�CV4Q�Z��v��2fb�Ꜯn@�u��T�q�D���\r1���-��i���k�'�0�3B�oo��VK��z�l�l,�&��� �&T��..���-ة+�[[�nR��!E,_H5�	vnT��6��|NY�'W�:&s��3��+'S����w.0C�3����X-j�(I���]2���|-�vf�F�uUW�jT1�J;�=�n����.!��)��[Q�h���<z�R��l^�{0�+�wV��}��l��x��\��I*�E� )�q�c������p�񬶭U� �8{KCI��Mc5��!)�Z.KA�7N��"�3��d��y�v��M��6_Z��LR:v�8W2U���GW�a��oT،x5���v��c-k<���ά}��9RU�$̇��}���5���򜚆<F��Au�B9��f��/��Ѱ��>�՚ �G֤��yp<�\�ԕ���`�0^{"��'~񂲲��u����q�$@O-�CsQXk�52�ϕ�]\��/yeY.���xөE��7�T�)!c&�����fK����J�;<�$�f<y��gr�
�$��s���4͐��5�Y�uσЕ��w��
��H��9�8�:7�uЦb�69�3fL�m5+�&��n-'	��N��F�f6�7J�</&��Qkt���᤻��&��0Y���2���PY���੗�R�q*���w��C�\��}�N!i۹3n#��ׇw�Μ��!��>ʙ�<EA�B+�a
��E��$;�����4�}5�fC���l=a�����_������*
co��&��Nv�P��=�51�b̤�H�,Q�:
�\(
�K��n0�I�p��sn\�B��X�s�h��ѹlhؒK4T`,�K�B��HFX�盪5dʊ^.$[!�	A�KA�-rs��n���DjM�[�H(�wXش`�&���҉.\�1�05i,y�!F�5�D�I�a��˜�#b��vPTd���"Qy�b��4F ��Rx�Kή�Iwnc9�d��*7��y�)L�'�vH4^���"l�o�^������}��*�ZV�Gf���ᄪX!��r��c�{��|����`�u%�\N�&���Eѽ���ο�W����|����Q�5mB�UT��Ue-j0ҍ�_?�[�SE�-
�C���6��y.t�Уxi0�0��Y�E��RX���b�|1\��ؗNmJ:��-wfW�����)��� ���ubMг`Ĝqv8�,(,��U�X�t��b���n��c��ؖ�����{p��3������p�1���Yƅ�u+v��Yv_�,�ǭ��Qת��Ǡ��X����'��{�aC�y������l;-���B6ԴK�C�Q�����|���or���U���8ô�i�nj��^��g&;��`<{D&
�C�X,��	��6j�u<z�������K7�,4q�.�8˱ǯ}UBtE��S9|ח}V�>������-];��֩�f��h��BS�
��m9�L��쇜= ��8A�0��#֯���=K[v�b�WWF�m�5!p�p�(E��	>�5�my���f�A��0�z\�"(���t-�.���k�<~����UEg��T*�����sE�j1��f�<)��4�ԃ�`�=��ï��l���r��z)�z�*�X��`��4#?l����fM]�~>?���W{O�߮�^�3^��[a[3�R[;�^�|��D�Ev=��_^����k��@�	n_m�M$���������pb��MT�Nnaڇ���Vk}z6����l{�g<�!����E�f̢��du�
`��٘�yD������������م�j-�-QTh��l�mS6֋mbKj�մ[k�����������������F�~�BeAb�I�*�w�Ӛ��z����v�[&C��E�cmN��kDMB�^�^�צ9�t)��^%9���5Y�|�O��q�=|w�nV�Tb��f_)�xf�/�C��%�h����v����w�ĲN��)�i0�خqP(-,Țw:74n����Z�O�oC�;���1#�*̧}��0�ʥX�ǡ��5�Kv5��m�<�~���|�:�AG��8m��P�����F�N⬩�w��$�+TV'.�{��� 7a1��a��p�;`>��y�kP���;4]X�6���tw�2LTsjn�3��Y�w!kˍ(z���Sa�8���P.A{p��R���8u�˻Z<j�j�|�q�-�k�qciS��mΔ��V�NKԹWҮ�;C���� ��9���R�������]�
�Їjt�ۏ��LxA�*Lq�u>��>�z�3�v���,3��p���sod�_s�A���P<,AO0��mC�ݐͲ/��c�C׸��&+����E���]x6KT��d������9f�g	�۝�kd�@wQ�\n�]���	P�l�2���l+��حv��ѹ��DVpJ�v�0[D.��a����@�+v�s#��`}�J��=K���dX&WU���5>z�@�ώ��n����ϟ�������_�kF�+m�[�Y-lZ�����׫��_�~y矬�Q ~�g�6�G���W����!���DJ�/���t��X�K��	�<+�����U���H,)%����^�>�H؊�X��C��Bܱ��=	�{87�sV�!�OBX��j2�[}�I�W�'�e)0��z�m=sͼ4��<z�sKO�P�}Np��Yռ�٦��k�c�ݼ|e�ܙƠRT���vP`��P��3f��=[���c�c�k��&�Uk���{QE��+�}E����/>Cy	M��LB�4��t�
=�Bޭິٛ����{�0�~�.,7"�ٲ��\��q�bY�R�ej�&�4Y�rH�tM�ڌ�w���KO�1Y_��iA�e�D�xSs������%�tD�I��Js�x�&uj�K��XGA��]�e���Y�涿E{�q����s�1�M��~�������$~�e;����ҹ���~�u;f��x�x9n��(�Y�yksj����y�E8�a!#��Bn�;'����-�c�n&��LGa�m��;�Zˡ���"�&�z�(���̤��E�u#4�@~�ь��5T~~��Y2<�^~�Y�7[���u�<'6_;k�<U�t�꓿�9��ݕYo8/��R��=���C���6<g�G5��[�����^>�d��o^!et���gs�4�Y}�q���0�'4;�%�Ez,�� ����;+�f �>�/����>>'�V�[l��z�����}��^��_��οu���X��5�w�;�E��)�����ܿ����$XׅY��%�uQq2۬:�7]�����ò}U=B�͉2)��4զ}d16�=��Y�'�㩡
>\nn��ƾ���J�`��X@A�<�v�E�z�hv��:�è15�=�=>� �����Z�ۇW�j����_@6�E�����p^<l4/��l���3��C��ߞ�����u�������[S��M@��q�ϡ�������5��P�:oD�9��O�F��G���ga�49o�˵ɗb��c�hU���~�D���ǳ�fԭX�M:�u���󪷠��+~��>�e)f�=$�W��d�&a�����x4ȧx!��&���ͣӃ������sW!�ʳbq��! ⼲b�VI^(γ�l�.l;���-�.簉g.�=;����7�D>c��[Q�H��[W��	��� ��@�*�"g��+\��Lf3is:o�^ʋ�5p�V"K����i���M��z!Z���N̈́�;�f�-��.�w� 󓙍on����n�؋/~{]r��;O~�cd?��������`T̮�L�s�fiǧ'/����)���\ow���z�n�|v̩�yv�&Td��V���t�N^ZCzm:5��gq�np���}�����lT[b5F�k�������T ��w>�~
��������S�>	[��Y��I��pF���@���"Z�.2nԿFwr�^��n/f"S�	*�Ҩ�qӌ$ȶ�@t�z�#a��^�]�y�Ź�x�a���:�2X�F�T�`�&+���W�t�z�o'F@��jE��k�;Ovh������P�#�z�YU�Nۆ�'�;6Ⱥ��4�4���\��gYQ��Y��^��Xh�N4y�9��'���5t(�L+p�/Fe�/)A>�F>}�S������ȈRD�R���d0t�17�=ά	7B�x6⸩������o�s�qp����[*l���t��ƠAC�i�B���t�>��R��WQ+��i�ֽ�w�gOF����zN������%A.(.�8ו���!�W����~^��[�;�wm5-5te�(l+sj��m�Mc�v��0��z��k�a��2%'��,/^�-ut��8w�^����AJK����o:�n�E�� ��C��rb��D[qL�����5̌�b�#_
{x�)�NԷ\ ���g�T��5հig��U~�s�p=�
SSxcs�]��ʹ��������믤r���J.x~��7z��UʛJk3v�Cs��f�������*�}��q�S�ɍԐ^<��X��:4��-q�����Z����5[V������������Z�n����3�<�y����e<;��/f�'�4��4�0���2w�=����1ij͖�9!K6&�h�ѡH���:����ٰ��6-Va���\9��͙���fE^�pk�.+��!�{;��+'����\:/,�0Ba��8�E��{P�Ǯ�����O;��@�~��εӝ|�]�C%�"d��e�/z૖�>z�+�/�R>\Bx�8�VK�;��'�Y��yK[U,���%6��&T*�Od�;��ǫxjkgk@Ų��T�l� ᵪ���b���C >�L�NW�k���Bn@�Jr�&	y��T.�f��_q�>�Q�A�L��ξ���Q�C�iy��3����6���I��d�s<��p(�a�%(m��5���seV��&�#]T�n�����9٭X.z���"U�N�f):a`r�E��Vi����6]�:���hf-�u�.�4�;�6�y�� ���#�&���t(��I�Q�S���)�gwmu��t7"��XJ���Rq.ka�d/�J��M����_v����?v�����-M#{>����F�2<�H�RPbe~3�to������Z"�w}�c{:��%M|��4����fS7"��r�>u8N��H �ݨ^�dRh.[���R�Ĭރ���*��%ݤ[̲��y�v˖-F�z����������������vו���9�j|�Zi��`[���c��V����*�K _=��*f����A�a*��q\��D�)ɦ[`I���қa�ac���q_�|`�w	�TB�יj���K�y�E�����P��9�������jM��*����xϧ��g���1�K=��7�w]�M]l�Z�P���`<y��:�_e�tn�Pv��)9��=(9��ʋFM⭭��즭���L |>��̽�!�O�&������D��{v3]"d1��`�˳wV;�4��隚�n4'��i�}����~��g�����Ai��I�OE��811�udf��Zx�q�bj~��p��}u?~�?��'�
��R�3T*����(M�E6n��䨪)�cp��ץ�'ӯW�8�:��u�מ��%T�m�j�=��^���Tߨ��͂�.?_��y͹��#X1��ע�Ӣ���Xڊ��)��)A�,Q)�WN��E㰭j��j(�'�U��g'�x.�t���,�L���l4d���t��Ƚ���?���SOC�1.���Ɩyi:p��$�A��gp_rvelCİ5���ˊZiK�v��W��34�@�ʪ���Xv���Ư�T(��V��ծI����.��d��)�nӨ��as�V��qp�g!��ám7��`�����)�T�Z�.�����er�i\�G������<#�v4�/��ވ��=R	��.�|T_;nd��SQ��؏>����Q���s�@>EîX�a��a)f�ڞ�a�`���ޫ�Ƣwg"�*�'K��NVyhb�a�G�˶?�q�[A�yȄ۷[7��jT�=Z��wr��oM�_�0BR�6a7C�(���[��,h�7.�a��O�N���5���*&��m�����A�n�騖��@W5�E��c�(�zO��Ļ�އ�h�0���9�Nw�j<���2K%�C�?�+�\�Ơ���0��FM���Q�lQ��y�R?4�ѻ���wfR��8�?0!�����z������4-_��L:�Ʋ�ūX��+��*�]\/��z�	����m��Ρ�>�`ϡ���L[�;^���?�ˀ��~��[�n6LOj�q����rg{�b���1�P/a�G<3ƈ�v���ër��ՅPWr���r���5�/i���1gP�����G�y�B{C�*���I��m�{p��,��.Ɖ�爩�6^���3��:�����q�>c5U��(f�8攡d�¶c2�+Q�� ��v�ޭ&��_Q�x��+Z�Jf��w%��D���-��u&e'�y���'��,i�ݷ�7Ɯ��:�f#ϥ�q����>��\�\��9�S��3��{��gm�{�}���h�]�)�A�0��|kO^�x(ntac9޻����k���L =Ŷ�������6������*�"��9��L���,n��z(�c�)��}#@� ��|Ǧ蛐NKͶ�B~k;'g����:w��S���{�-��8Όu�5{*.[�k( X�.2��󴮝dՓ����u<�]��ЯN[�\@f�!��_Ec�Z�R�TXS-���T��������t"�"��N���V�V�޼����B�����	�{1�X)P�~�E8��/uk
c�]ޏH"1�^��ʚ� �L��ݵ���8Q�CexnK��b4Ҥ�<^b�sȢ�q�Lt�vl��v��S�|&��Vkl�B�Ap���C\��/C6��*���JO69M�.���-Z�H�IZQ:�v��jޤ�8�S�K>��A^|!�n�t]tZsf��u�ª̮xj��//����kcrVv\>�:�X֯���H�7��B���c��'�r��PW�>�+��g��_�,B�h�S�S�M���n�ܶdYǺʴ�ӵ䂵�%�3�����!���/m�o@�f�qP�ӈ[Ӷ�ϵT�|��7H�ҡ�����wu��zrV�!#���H��,�"��[�5l+��D�]}��Z��nq��2��� ?���7���!+k�|����g����V�����\��W�/���g��?��'H���iR�*i�n�C�wY�?M�Y�[.��S���Ts	hN�{�=��4�̨cO��
j�d9+�(��'e�mx�&�0�@��k��E�Է5�y��g7��G;�W$�+�w.Ǟ�H:���պ��m.�t�t�w(��1%ی;} ��i��Ʀ�G[�^�k�#��3(����F����V��)��F6��wK0�{!����J�4K��i��.!�d��;�����Z؛xc^���
�eā��ؚS�V��ޣa^�+���SUpc�
��X1���9�H��t�P�E3���zä���K���j����S5e݇���ӜKsv��^aU�B�Ru���l'��*��:���9m�Z�E���{��<��34y	.�oN����soA�o��ʀX�R{U�B�E����i흷A��;	�\����Sf�:�\J�0;�d��_)��B�	�y)LPRU�7��?�������^>�o�����~߷����u�A@��<�@i�Sg��%�Vq`�$܁�wM��:@KFi��֙B�+�ME�:Ǽ����w(!���UV�Cv�eC*]���Q�_/��}k�h�;y��i�y�asY���ηn�]�g�v����՛���yI��@�����Z�?F��6h�ҳ��Q�$�dlݴ����Ttj����7�r��;�l׉Ҹĝ�0t�A�ÕVe��[��ׇC�Z�}d;h�w]k�w2��ð%��*��T�S:�����A����v���{�A��Z��`+�;�ѻiإI��v�д�ݓ��_"� �]�]�S���Ƭ�ј�T�*¬��,R�钐��"n�X�b�q�{�����J���5�O�$Pf�pf�0�Ɂ}�d��6yw���F��+�����M��%k�:��2��)$�<s\p�*�٪]�uڴ�$����o�6�%�1����{�.�u9]�9��,c����0ɚk�8����*9�Ւ`��M�c�4w	�œn��	js�1��gEN�u����-��[5��E�5���xֺ���PR���;E^]G���6���	�3me )$�Y��\p�����q:7���ar�tj�w�:���V��W4�[�1��,i�È�@D&�z' �z�em*J#��9����D*�Q۾�L�b*X�7\���cM�$;y|�42��0)���ZLƃ�\'Raݎft���Ե�����4�d�m^�����\���]���أw�%�"��>٪���;�+����V�=]�y.�������O�AM撄�e��S�u��}A����ؖ� e��q'>9۫^S����b+D�P-�1�V��j��N�'�*�kES������kw�J��ٛ(�X`�^��ػ�[��;��[Aض���vQ��}2�r��W¹�c2<;�R�-�����dQnp�6<�R�ϵ�כzq��t���4���V�qr��
�^��Z�o����2�뮁���[YNA�q�<6����wkꣂ·eM���z�,�w�%�(G��l�jj3Jʐe'��v�7V;�GJ�0��<Z�O=U�2.2��O�>m���׶����s
�7�F�n�,u* [ZH�k\�5;G�)'qְ\Ѥ�(��2T?�����3���7�E��\�n�j2�X�yu2*4�q;�-8* $9�s`�5)�'��ɸ��U�����3-�ޝ��q�����mFEd��Wػ�,ە%�V����"�{W@.��P��:z�6��k'}�H�S�]���7bj0暫c��ٗ'�"�4������
/�N�P���r�cj�V��Ŵ,	��.R��vԽ�+��\��' ���ڷ�-�]�>ۧ��>M�t���A����o7q7pG1H��Z��X5�S{yX� o� ����;���	�&-a��665ʸE�E$lf�v�(64,PjHۜ��B�X��0��#s\�"�MEF��]��2QFMb��F���4���6�����wqb�r;�,��r�W9�\��.EAnj�A�Y�nTb��F�1�\ۚ���ы!r��h��nnQ�Z�ss-�4nF*,lm�N�-�\���\ƹ��F4X�-����5���F+����(#G7 у�r]ۛ�c�cÛa�ڎW;���cs��v����������<��q�2���*J�
:��Muf��vUd�����.w�W9}�H�qT=����!�O��nK!� ����b����9�2���ZA6�%�[!��6�L �%��&!��ﾏ���q#gs`���x���:w�Hqm	����O]� ��5�L�N�^�gN��XΜN�����dZQإ�[�8@=�ƽ{_ZG;6X�,<s��ȁ�4���Rtµ���bVP�^v�l6.�[���)���n�4��6�M(fƘ�	��=!1�a�Zf���
�a�ak��/�z{uq+ۛ]BmL'�҂ƀ]&���p���XG�M�1�5�Z5�{����XW/�l�q��s�Yb�v8�0�j;��ҡ��sh/N=���:�ll�3���л��0i.T���OQkeb�a\�V����߂�搮�ht[��Kr���S�֜F��K�� ����>h��Ǝ⡹�l��U&7�Q���=��3<�[s�dI8����y}�����3�`�����<h�^D<��{��2~���>��_�1�Iy��PI1k��'��̅b܊���N2k6!�'��~�!�����E�;��A����;�6�^.�U���se�[C�&�D�MC_��4c�}Q�k	�����2L=�N|ޞ]R�z�8~l�ݝ"�j6�[Ƹ�d�\<�ۗT<9ZɊ���ٮ!ق������OS�����k�o��Ծ��,�S�ݮ��{6w�]-m%��f�c��겥jX(���ܝ�?��p|��ՇSF�X0Vi��a�Y,^��aM�v��<={uz25�������P���,Ӿ�XrW!�2a�ȼ�OC���T;�����g�L��}_�j6c	1O��2��}�5>�{؋l�S7_���,�`Z�;A�6m>0O��j�w+.�rgŵ�������t88��Ƚ����U��mEzF��lr�2�����Xd^�m�q��ij3X'�vҬ}i��w��t�#K��`�*���N+�K"��I�֮�K*�q�%�b��Z�V�k���Ơ9휼��FC���S�d3����}��Y7L�k�H̋ɭ�
v���R_-��O9]X��4���y�ϑp�� �5���m�mOY�m˧�J:s�Lu�fʗ=����U�㸝Ti�I��'�W0��e�>G�e�[!��hސ�_�k���H��[!Cr����C�R{
�ia7C׹E�偔�_y@��,=�!�s,]C�����M5u�0�d�t5��ķs��Kv�*滼4���̡����M��؋e��r�>���!�>�v�\c;���<����Π��.L�Vt"��z:�k��Hw�"*��W�2�Puơ��-_�F��	n�,���F�P֚X�@`��g�ɼsE<9�u��k��ܘ�Q[Z�5������c�z�/\�wG�jJW׼���v��J��$�l�x2e
]��n�abv.���@�A(�;�����U|���y������e�2/N��:2�n/��mpz�����4-Xu)�vf�h��m��G���5�����O<�<������T�C��x?��5�<�Nç܁W�����t[.�/87GgRsg�L��
Za/<���,Z���xg������n��ɎRq���U��s�Ҧ��������3��Α;�3Eی;���k�E��q�W��Y/5�#J��jw�M�զ0 킞�D���Tk[�ւ{���n*f��%ۼ�� ��L�M�5�N����k�7�����x��.�p�!��ؗ����حj[	BX��Μ���-v��|�%�f��t7&�k Y\��I;��0?ߒ9�a˃�ȥ�.��"ؓD���3־��7U�ˮ}'F:�%��ˀ�g�o�^ʋ�6��
�+�"��W�'��˧Y4Ц�cIcNA���z���8G]dF�<�TQt�H�UQaM@-�Ưs��Y�:owA�k��񘓶�E�&�j��L3`Ad��
��>�O�R�j�QN.�l��'ݑm
����y��ǮA{t��K���Զ`����ʺ�o�Z�s���[�+�DM����ۑg#;3�6�5��:��7���=�yʵX��i���9j>r��5��uRT֓�4�ޫu9X<0��F&�0n��Ε�@l��Yp�mԏl��yv��@���% ��D�����F���x,|��C�&247vC��v��4Ҥ�<^b�sȢ���6#�˞�%�@��a�J��Zw{TS��h"1�C�/�= ��\C-�|��^�Si�S"�09�2U��<nD��p|�%����{4]�3�ㇶ�p����z�I͚�o&f<5�w����_�4˼�tו�)�-�`��ٻr\>6��t����_��x��t��#o���1��;
z��qH�,(,��Ut�XHOtZ�+A05
OB�01���ԯ=���=��Y��i���7�;��/��4'�㎶\}K��%�	Q�%m	֡�aߠ�_pèN�,]�?K�U���5)gEʓ.�k��j�>J��q�i�i�3�����轆}
��U�Fb�^�/S��u��<`��#m��NK�N��Y�Aܢ¸ėj�.���jl��5�����+�������_��+T�.���24F�)�z6��u3ǲsǤ�v���oe[(����A�m�����r�?�X%��I�;�1��5�mc65��_���e�i��=����o3KD��8�=$c�z����npރ��X�zЫk�켣���jYD�۶Or�`�3�*������_s�<E����>�-�u4�� 1��ԫ�C+��\�]��#��n�V��[y�sG%MMN����� X*U���ݷ���7�ۀ�����{諐�"k�7N��L\:��g�`���$���h��#�i�T)��o!�n��R��┅�gaT�(Q*N�~�l$\�1��g�HBSsS�U+�l4�U�{QK��E;Hޜm�کnnt!6r����P��vл=9�C��3�>�SJ��n\Ou���d������|���vO�l�S�΄&<^%9��0MAIT-x:�}	;5����D��&����*��{0R�����WQ1�ʅ�������}�r���^~�ƣ�t��呙�ȵ�=\�Y�~|ɋ}mhٯDB`��zcXD�Ve;��S�{~a5,����5ό�<��m�i�K��4��6�8zh�
��G[���L���V�n�'_yU��䴞���aC���UZU��-E�洠�]���p�����0t����q��F��n����-q1%�zzm�jNP���B�w9��w= �4�>���O� 8L�*S�غT�N�0�]v�1���zvi����IE��]+^�(%�^��2��m�?��\�?~��$�c��}W�ͬ�rU�Q���5j��{��Q��6�B!�<�Np�jO�̸�a1e�s)er�Z)��ɳ<����4��Vb�L��\= ��J�*�;�&+����k6⮍.�7��ǵ�C�[�y�{1_������ �a?��O"��H�����l�
���GS��N<ZǤ��yh}���[��Ы��2�	�T
?��0J��Z�+��<�j?V�m��_��l�k�j|��kR���^����;)�ߨ�bՖ!��D�ǐr�����E��N�k���rw��vW��٘��GONjV�ki]���'���o�؊��xgA�ChC ��UOԡ�"�	uxyS\���O}�z�6n)f��Xu���0��^M��y��ֆ}�Z�W6��۲뷯�-��q�"22��j})�׳8�y*f㰃%ql9�Gh=�6�1lE��|Q1���m�v.����N�C�k��.=<(U����O����c��ɩb�O��\�b��s]���/��ڙ�.�SY��x�� `�an���5l�(d���t���q�*ű�|5�1ó�|Y�]�4�£I��F��P�t��{w� ��Q%ڼ�b�C�����A�QB��]Xe�4�#n������b%9��E1��)��G\sk�\:��<��	K6��̚�A��ٴ���{g��V�q��gw�Z��)�)�C2�65`��Y"��M�w��ڍ��&Z�; �7x��V�f�p�ؚ|�T�1���3jЩ�r�v���,N6��W�ŷZႝ���7.��Su�^�,j+RnN��h�[��9�j�;�+�wK���;��R��yO�{�E�@sc�E��Ϛ�-�Fb�1Q"ޫ`��h��D��!1�ON���mE�v�Y����?"H%�o)�B2��7{ͻ���*���-�9g�:��ÜLlK{�U�7X�U�xa��)\����E1�^0-*���ɳ�����s;Cs���ݙ?��\�	b��52��t+�d�{꫺^�ݫ�b��\��9��'tk �<D?vmt_'����i�kң�#3��0A\3g�{O0����{�}[瘶Pp��A��~��GNy`�r�9Mi��N�v��'�(=A��RN�3L(w���:�Cˆ/�re1��E�D��=��^G.%S�:��X��Rm(�χ:D���\eش�$e����@b����V��о�-� C�]�>1Ǽ�X�0�gú|�/�L��I.�/M��G������`�6��`�wզ���������<�����1 ����Ƚ���W^lV��H8�rb���߫�G'���o�6�z��q7�osHL6)�}B�F�y���������%&�oA��V�9f��o�]�:���uѹ�DvӬ3e1{�������9{�m";f�$�7cB���sX{��8�6��Cp���'],��7	�Ube֪(
�irA�+����W7���g�cW���$�y��`�)�Y���D܂r^m�/wczj�DU��]9ֈocsn?�,�,h��g��|j�T\9������Iq�Ꙏv�E���{�x��<��u�yKC&19wA�?'��-T))��[@[s�]Qp���D��W=��wOb�K�t��N����C�V�Â��=�)�M�"�)�◽8�GdX_��*�|��c��A��96uĻ�sy0Age�ň��ʻ%؆�1��J�,�&*�<�/@�4�o3Ӊz�M�3��u'muR��O�A�v!?g���q��v��E�LSs}�DٳtU74�b�RSd��1�W�zi�?,s�p�Ѓ���Cw>OE'7&�Q���
ޠM.V���L\�gv�Y�xe�s��('��i��%���(�ð����6?�~ن�'/�n��Oߎ�����~�+����ܕ:9�U�%=�}j��Lj��-<u����T�:���_f�Y�"�N�Rԧ$&��B��Ԭq�˥kߊ�^��G0��'Z���;�þ~�z�jρc�t��:� �:����׶���7Ǻ�֤y�E����J����Lɇ�#t�Z�X��%rW6���N�S��ū�i�;�қ����nnW9��a�Y�<6V\d-�%I��V��0N����������t��E+-�{j
��}������S[ꌜ�n�����	J�`�|H��-�;7�~��u���K.��o_v��q�F8Or���5*<D;M�����<�������
���"O����omu�2]�uc�Y�|w(���]���y��V����{$?/��4�Ug\/+�x;iP��B�,O���0��t$p�w���Nܥ��4�n�z�TW$ہ� ܌Cp8"�Pok`3`.!����'�s��^TM��X�%��bTIy5O6C�7��_9���B�5���M]1p��x ���;y�i�BJ���/��G_t��u�ƭ��*[7Μ�Z�vd�f:~����h�޸*�Zh�֦����B�0�o^�}Н��C�;�d�q���R���D���!2�,T)=�Wm��5H%���@��	L&���ד�ފB{�������ӊ��^��|������ħ7�0M�ݓ]�:��M���Ɵ�����#g5�>��=[�	-�'H>T���hO�_�W�Ԥ�P)�2�g�q��a-���&3ՍEL�Q
{����}iٱ�0\���!��%G��,�����r���|b�f�]��;��-���?n겤A�T��l�`�]N�����k�Ћ�pu�I�bw�2.���+������Y�y쓴D�jJ����g`�t�,!u0l�T*��n��b���$h�zÊ�1�ə��`��Ys�͐�Y͑�u�r.�o8��r�E�7E1���ۋ�/	���~d���U/^e!�����իo_���B���[�S��Ut=���ܔ4I�栜K�����=�K��4��0����A3�����T���ę��	�`qTa��w9��C��,��Z\=�.vu�DH�fP��~�s΃�l- �G�8}�1�-�D��W	V0�r�Z�T�/j㘇cl��*5E;f�^�:�Z#6]3R�Űs#�0gC�9����>;����M�r�1>eO�_GZ֐��ݦ-fD�[n�}ܽX�^��P��5����(�y�V0�/�H�W�l:~��!�G73��<�����e���X.��#�C�&�r�����Ű��z%�<������%M�.��(�'�^�w�|��]v��f�0���C�gh��L����A��)�k�c�0��a��}ɩ�ʪɳ��M�-C!l��I�ǵ��9�f�i�ø%��#&<�M��sE<6]KGs*���F.:΁M-6k>>K���O=z�g�䩛��ʂ���������yz=>>^�w����{}��o����Aeh�} ����٘:�#������L�g9����I��)Fa��-q��`�`�)�u�H7��y}&.M��P5d�Z�� ��C��[�����d�Y:H��S8X�����Uɻu������n~�C���C E�����v�ܣ5s8���E
����Q��O�v��7f�_m[r<4%+FD�b�p�n���v�
��0!8�jQ�|�]�e�E�n�y�ӛ�5/�PY��KR;�e�A׭��Q���MC��;�>�*�J��|o �TaY�JΘ(�.��?��0���zP�4s�i���d.i�~��$v�*�h,�6X[m"�&�	��Ѿ�S4�J���K�A٩�w~$u�,��g5��Bj0���A�0�ǖ�Y5�!�l}ِ^�h^<����2]�%�3B�JG�	�)/C(*ξ�2�Sw��:�7�lP��5.�=zcG���N��d�27I��(�J������@����zF���K��5���f��� �E9��w�f����4�]��%e�f��9��6�h�1+�痹�ةiԸ�aIu.�(++�d5��L���-��e�erDn���o��z�,�ފ�^~��{����}���5�z��L>mg��jh�Y��Yx��f>V9�4���:�O'32��hdtwd�N�%\�9��,��������is�n>Ѷ텗�P�ٙRKsF!��^ )�p��j̷*��v`x���ݹ�}�*{}�wTd���I~���/Q���<�L��j��p�w��8Ͳ8�:3K�Mn��I)CW�QY����"a��_�G�)VP�Ĭ�,t)V�*e�_T&G\�M�ƎDخ=��`�	��me^�nٿ��El�ִ���uc�
mlʾD������e:�R���p�JgETW������*H�iq�+9�a�ՔE�R7;��{�2O��S
+w�j��r�c+O\�M�&jĭ��
Ő�d�5�Du�w��|�U�NPH&���xx����ą���1�lp��L�{�8���s��^�
^���!�r[5�h�Ѭ�N�4��M���x�ⰶ��ڼ��}bn��.�J���:ܙ%,m�ap�&.�Y��I�ff V���I��m��Բ1Yv�$[�����LqUu��U��\�{��$�nN�h��eu�O8<����A�vL����V�[��ס]���naL6��cy7��y��o8�q=�9ޚq�}W���M��ʭ�y|ݘһ,g��u)=�G����gp{���U+/�^�:/�6��R��ʸ�Iٮ��i��$zsPA5�{�Zxkyg H�Pm�A7F���(�ޚ�\�dWd��USin�\eM���j<"�E��қ�5�{՝Fs�k%ш�޸�*��o�n�re�r��:_*Ҫ�g�Խv�}�����5�/����������h޻���;�4�ߎm�k��Ÿk�9�b9n���űwu�4Q��(�-��.h�+���r+�m͋F��(�u������rwU����s[��ӕ�;m�V��6�;����\���F��wv��$���M;���n�nn'1\ۚ.RF��(�[�pƻ�r�]ݴk���Ewuȭ�܍�sss���ɮR��w7gu:��Eʒ���u�q.:u���y�˺�7,h+���x�󣦱�7,p�Q[���э]�nk�ss�2��y�k����r������\���您ũ��n��A]ݍ��#kr��$@$��=�m��{�L�
����}��v1�����c�bl�oo8�l��	�%��%�*f=^\LcN�j�~1���6��yQ��V�dS�`qm���b��V0J����D&��(2c�*:�0�۩ƽ�����{��a��n�-��վ;�
N� l{�M��xVO��;^�X���_w�1�6�e��1��-��Q,��I��Ѷ��ό��Sۼ	�vl�xL��7��M����l^�d��l�s���̜O��'�)ͮ�Lh�I��:皟"��{���[e��-����7َٵ�:¡3r���e�+P��oR�����s@�ju��=^�#Ͻ�;ҥ������s�.��*`��y�|n��ݝ6Ԟ�v�n�S����P	|\��%���D7P)��Gi�U���!ko���l0�`�01���C�dLK~��nќ���{�0��~�D<��<�I5�$?9�p�\�!�&��xQxk��W�G��P�B��ɐ��4�Ƹ7�����fe[V��9�w��}�?�_������fgv��
����(:�yP��-���/�G+zBK�gS���B��1��Q�����gO:�ym�����(h\S���}~f����3�P��2���iN{�٧�k�\w��Է�=:�1]gL̜V.�ki�歇�G�!vr�;�V��%&�`x�m��,��wGr��w����4�e�gTs�Pp�6۷è֫���N�xT��y�x�ۙ���Ɉ�vZӭ*�]�uc%鈴������w�CN:���� uX~�f�pl23L+�@�b���Z�{�<9ុ!*H����;�f;�vZ*1�&:���wHn~��C��v�2�ZI������h��;�7�W�ח�n<J$K���2�&
ubzq���G���3M�I.�E�b��v]im-����:$nچT�׏Z�o�E;ǆP|a`=Ų/Q���Z��A�-�����0������`le����r3��3f�V@�t��N�����f<�x��\&z���y�j��s�p�th/�~;'X��]Z�_��*-�U�J��.�~CNa,�O��ﻯ�y��T]��mj�Lw={�e�|���U
V��
e��/P��3�M`���q�L�*"ow��Bv��R�t%�uڀ��d'�K��	�{1��R"U��b�goq�W�r2�.Ej����R�K�%��i�?0ѰC.�v!��C4�2��c�E�Dܰ�[�dv�<�6�A�g�w˿D��l��p"1���S�/C	eeK��5)<ϟ��眞�uM��!��۫���{�XoH�����lRˣ�3�]��L�c���J�k�k^�)���m�G����g-ݐ�E��ɣ���E	�+�md�����z�{zg�L}G���t�Hv�J�ݾ�1��h�e�W�#��S-#Α��;9��0���5���m*�Z�2�����B�c>�{K�����L�ߙ��8{h8Z�Cw=OE'7&�QSأ�Gf�{|��Qa+ۓ��֪yJ9�{�Ӱ��٣ې��m���	��Í�#S���bZ����r�5t/S·�O07��i
U�%=�}njp��1�ԩ�+�8�8���ҽ};N`T��)���#�hg�Ԭq�˥k�PH����|���W=�~�U��)=Emf�tk��5y���6��@}�U;.�hv�a�^l�k���+�Ks+�J�6�U'��h#{�#�P�uoa���K� �<h����߬NK�N��=�ە�+��G�L>�j��+�P/��o�h��w�xr$G�m(<��P��ٟB�ء^a�>0�ۜds���
��[�Ql�����ֺ����!�p�j&a���e]ok�����q�Fd���W(-7P�f��cy��r�
�֑y	x<��#�(�HA�1�i�P3���,͊�+��g�md�F�_��=4�է�ԉ�Vd������%�"N�G�>�S��P�<��v�a�?u�Z\��iJ��d�T��H&�LYz�W�vRӀ�t��Ԃ�ȕ��.�/����馀^�����`nf��qJX!ٻ�c���w����A34�Ӝi!�w��ҭ:ù�f.��|��ѭ��8����V��ǣ�c?���H&9�C�.�c.کnj��"�]�R%�D��]�,���+)�3f�Sz�e�Wj�5c�sռ55�����{3!=���1ͽJce�S��M�9��b��}v�n�������K\5ݓyC<VЮd���O|�gh�5�|(vT\��z�YN_vOd#�޴��qu��LJ2�容
Wq�U�LD�_��˧?�<x���xSL�s1�~[�(��y�]0�U(��7E1�]N�F9j��54���oeT��u���Ѻ��;��B����CХ�S��Ut=Qi��(,kˤ��&����ޗjf-�V�:�5U�0н�0{b΃�,���6$Ͱ-C	��I�6����*�AdmD'��<V���ŋ\:��C�
�tz�:�^��mV'����J��]+^ʂ^��庁؝�6�dm�]�,ʺ-����8yGvmtώ��7:@�NT�'M0��1�f�l^�}讴|r
ϧ\�G��p�P�Q����y�Ƈ��55a{��O�7��c�Y99����s���U_�̚�ۏ����{~W���~��n�m�n�?<�t�=�GyK�����0]6�N�֘�wQ̌۝:Ĩ,��Ԝ��Keb��/u��+�}˱|�X�3�W/
�7�n�Z���Cƕ�3������$��w��:s����}�@�b�t=1l�C���w�/,46�qn�r��.�yc;�gs¼t'���M3����A!��K�{����k��Muc�9�'��=䝝D��ֶf֘��C.�m��=�g ޡ�>��L���p	e(#&<�y6��4�ưRO[��wx��S�<p�iiC���FS����y�ٜj\�3u���*'w�-���^��j�|�?<���~ܗ���AI<YX^�V�k
+%{Q^��%6Ǹ��j˽��kY�/��Z�4\�F0�z/���վ;ǐP2F��8$=����/|����]��u*��5;���K"�
SL�Q��qo��L����� ���]����3]	��"*6M��4�5ݪ�ɤh��;�t]x�Jsat�c^(�kk���lz�\����;}ϫ�'��Z��3s/�,ʺ��4˰R,�w�ޕ)?�NVxsȣX�Y�_0�<�]�n6<�Oi�y��s����F#�����g�vtSJ{*��au�-? ���O�Օ?����2�����Y�Orm����k��3��|}�Rǰ c�y�C+\�M�4�Je�2Tw���4�`[)��F��#�X�ϔ�����H�o�qݖLZ�Et�b������V�d�W��٧�9ܵl�.�Xiӻ��Nݶ`3i��t�z��Ub�k�d^m�R��`K�ߘE�3�
5����˞��-���w��g��w�9�e��%B�)��Jwo��k-{����H�xQ��: B�Q��w�N�\�\���ʦO���ȱ�oP�6(���\���̱6���s�?UBr��i�Yx.!��Q�k��]�������n'�(Y��Ja�ƲǱǧշ&+����Hwn�����M�V�ry�Fbp���^�4����~}��A����Fi�qפ�s�ncϾ�0{o;��ɘ��z����?��E��Lq�.����۬U����\��G������?9���߽M�����jZyL>O�A�4[��)�t[m9����f�3�z�v��]�;�&���5d�q���_l�[cW>y��C`��/��g�4�����r�}^���L�C�h�����{�g��yt_��R��墲Hb�c=�S.���K�X02pBO~������_uMO'S����@��Ư'�:�7x�Ɓ]Z�^1���=�m�5���g���a��U�	�<�����eg'��2��^1���MoKVRm�T:�����ڲL������C���X6���ϓ��m��(�b��Eq��,\_o'�ɧ�c�1s�K92셰^pp��f���
�߆�'�+��n�[
���޷]�lw]���5�"స0�˔�&��\��2ױ�):��P�aU���j5����Cu��)�N��S�'�g�彏p�K��گe���Jb�:!2Of"S�*�J��]˦j~,�n�ù�����r�0>�Ш)��H��Pp��2��.�4��ftҤ��LR��ʑ���P�3;��G;�+�t�zw�xa����i�!?P�/^�YP�����v�p-䖫��W��+��2)���^4�\`��+�%�r�+,}�!�T�5�{���a��L��=^�TY̷Q��(�oW0��s�U��^m),hr�vâX�k����?>O|�_��a�%�^�-�v)>��з�4q�/���^�>��~��Zhr��P �R�wdk�\��k���b�Z| (�5=#�s��\�V8��V�����Ts	[Bu�y�2��0kzef=�-�#�Ά�g��N˲��m�
V2�H=K��Fh����m�����ۇh�]�Yw@�z�ԃ"]�CD&�o�9.�:�n�w(�>o5cl��c�ڻZ?~`����Ԇ�I���M��tw�k�&��=���|#C�(Ǝ������4ZjQ+jYID{�L�����Ɋ�S+�K���IXgm���1�t��ղ���׮�-����)f�N��;B�	�&žq%�S���He��=r��(
�B��Q�w���G���U���������+�j����3����S�
�8ȗ��M¡17�n6�S�^kA���݌��@�C�J2X$����؛xcC`3>d!\1ea��>��9�ү]-��z/L�cZo#�yj�G=y+��My��]6��u]�Z�a�,�9WA���^!�\=�O>MF5,���<�-~�!��D�*�_�E�N0t���;;)^�ۚ9�a�)��ll�8�v�N�W���b�0���K��
OOI6F4
���nix���
Ӛ��z���Ol�����v�'�!>���nt �m�"e��l�Wf�p9ػ�W��0MAIT.�7�^��xOV��C�d��^	���z���MYq]��[eww//^L�9,��:\�Lk�L^y�>{2�=��@�a��ώ�oWY�u��Jè��;@Z��6b��9T�����.�n���;�׀����{����*2��`�ע6��r܀�#���F��wVUt=Z�O�~J���Rq.|޼��f!�n�?��9���T+
����M	�
�Ґ+�o�Kc&�p�@*o
�r���rq�tӥ4�Ū�H{���ht�tgI�D�G9�d��*Ûځ;M�č,��6-�ĺC�M����:u1�r�!����Ja�ڷ8�������<�9 G�����B�����Ꝛ.�	3la7"���@Z��3t�w;Iu{��ٵ��-�/����Ѹ!�����ֿFĶ������%YN�J���-�0������}ڣ���[��N�;!t�t��yg�_����7:m�����2�"�N�PNOn�mA�:�,r�N={��1چ�9�c;0���|�<��7�P�Ru��E�*3]���d3lڔ_�1�!�c���_Ohv|z�G��$����+)	P�m<�
����XU�nQ{њ��A��6��1�$?q��.��n=n��%���k�eM�����M-`�6t��gOS�Ӛ��4Nn*f���è%��#&>��x��������5h�0�*.�כxi/,�bw���&||�1 G��E��5x.J���vPdr�~Ⱥp����X���d���_��٠��[���s�:I�Yb���_�N���`��j+ѧ��k2��^&����M�p8ܻd�MAb�O~UӬ=[�M<��}A@�"X\� ��U!�{��L�$bݴ�ӻ?�����h�cM���
+�pC�n���}�$������kֱ�A�Vj�%m=�6�d$�N�:�6���ָ�r�4x�"�\^_X��x�0J�%J�ɝw7�\�.�
�r$�0mnL���Iy���-�!yYV�:��qr[��.�Ƚ���Z�I������l���� ���.�M{��Y�R�/����ў�F+��t�_}��'�b%9�.�Li#I��P�M��a�.j�]����I����͛��}����r�{jHe^;.�M�N�zT��b)9\��)���+��a��P��L^��v�5.����l!#��Bm�;<���K�.�ɵ?'��Gj�}��wQw����۫<�4�O@~�b�xEօ�>�4t���s��L�τ.L��o��2���;]k��nH�0��w=~X���,k�����˽S�W:���&�V1��Y��������� �������E�y�ѓo*���U,�[�Ͳ63�����Jw`�)�ԩ_C�d^~$�hy�Br>��BՇR�u1���q��l�b�A��B�@�`����w�]y�B���:��h�mi�M��	�~}��h?a���Fi�qh��b���Z�ͻ�p[:�3=�Y��7��`wk�<{Dk;@Ca4���6'dk%`wPnys�Mq�.�8˱n g��������^^�o�����}��/P6��o�ч}��bi��r��iT ��E	��%\V�Y�	�Q׫���jയ|�k�!�iui+��;����u�:�ܹ��M=�y�.d:�-	M����2�q5�3�nd+l�� 77�M��Z(�xu�/�6���0CL>x��{����w7D�64-h����n�M���ht
<mԠK�@u��ꩼN�[�f�+A�����f�G�{Zx ;(��6n〙s#t2,\�k]b�b�e�V��e��;��,�I�2���+��\n�j�t�8��h�o�z�y��.�]�e��SC;�ٲ��bbA$�;`�8eZz���b(�+
w �,}Q��0�YK��
��/3^��;OoB�gh	CH���"逊K�.�� ���#yl�{c��sLw2�s��k�9u�"�YE�x�)���0��KQ2��K/-�l+�p�4(a�}�y����H��	�:U��z�����tT�7i���V>o^�in+��96t^��d�D,�q����Q����|{��c����%r�"�[�� 6J̬}%��o-}q����S��L�ei��e�O�X��c��:��<��Yٍ��环�6ۻ�浄����gq�E'6n�Ji(�M�Ԗ�]��^f��%��V�:�����'�)fS6�`�Z#.��78�0!����ą�Mf�{|��@�v9� �Վ�d��5��W������G�O�qV�Ѧ΢�������*����v�2�]c���I�#�ɸ�����1������N�� %�8���N��4��'X	��`g!yX��\D����0������
���x�#d�u�`뺍�5w�$��J�ȤGl�l�AmgWw��|���<��g{|�"���j�t0s���ݧ�r���f�v�qoӶ�lZ�J|���!�V#�A�șG/T��ޫ�NI����[��P�'8�"#�A�!J%y�*���v>�;f�TУ5��)��/���[u���b��P��yd,�e%(�����A-�-��y�nd�λ�A3��k�ǐc3���J�� j�;��|n����욝0��K[v�6o<�̲JʍV��=T������#� .J����VT|�/J<����=�y�JB��e�q]�Kt)�xU񛊴�t})�g*�3�4��ͺgX��i�x�i�16�28m��
>�[�'
$�//����x�C "��NsL���tNK9���<w%4�s*;��a͆�Oz�s����ČY�V������ԝ�6CKL�ͺ���Z���֕mO%��]��:5ر�@A�N�Di�p�Է#ő�z�V`�%�̣��Į����Ԝ�&��@����\�AP��3�<����J���K%)�;���򇷻1��v8	XGKi���ج+�r���՝u�XjH+�fyCk�l��9��ܹ!�}�̴��2��ȸ����
���/뺮�\�����\���h˻\ܢ��-�u��3�W���S�F��ZS�͂�5��9�ME�mr;��lQEq�m�5�q;����r��mݝwv�r����s�(���(�nV4@w\�U���9ݮW0ƷwE�q���s\�r��Ts�4k����r���6��#���s�d�wv�+��7廮�.;�ۤt5���㮍�ݴt�U�\���wQ�+���WCѵMrӝ�;�+����+��sn\ɮTd�����X6*-�W#��r�Lj7;���5ˑ�Xwncw]��u��wW:f��Ͽ��������=(�7\��=��)5���]3{-��%���(ܻ��4oAiE&�H�i�K	V��6�V�Ԕ|�m��{�n�V�G?�vA JD�dĄ`���{/T��f��Z�$�SC�=��*�->�6��<����>q����Eo���u�r�m��uVS`�-�V���ȹ��Y��qLCi�B��׹��{dS�{�3�#C�["��ϫ�����2�D�3}�C���̼z8�BZ��!��:ϛ�r���zw�,8!'���/�+�Lk>�ig�e}ʩ�9#6򢱨�B~ka����
��z1���2��=3f�	~�x(d�\�:�>��gCp<c�S���Ӭ��as����RukU
V��
jnq�{�pnu������;�a�{����ހ�K5�:N�/e����S��	�{"S� �B���1.H����C9������'O�E�u{���F4�C�>���]�i�3�T�W����\�z��{��������W=o�lS���-��@� �cO��O���I��YF;e[:�����0�h]]ù���fT�<�d]"�9��{��{��Yzw,��5�y^D9��g(m��Bql��}\χ�e����&B̮xj�r��PX��i�O�û4ƱO�Xu��=����q�d�&�M�e�Our�����f߼���%�e$�\���`�C�i���O�v[O$\� �DKg������֋.�^�Hn��:�dKV�w8�n�x9���[�-5G}p?]�	�x�����EHi��yr}}0K��K��{��^Vsn6�N`�[~��=zTRsrn��1']�TXPY�̪��Z�5�}l���zZz�+��֦^�[)~����pVr�t� ls*�9���L�[��]+^�T��%G0y�Q
S��vU2��{ܕ�:/i¶B�ù�t�#��ن�3��秥�m��sPl�kv��cuU^D�4��u����X�j[Z�=ʡ�`�O�K��T4?�0{k�4~Kv�r���!ҫ�B�����X!�����b�zD`���}_t�--*��yO�3��(�ּB�W:�����yT� ȴh�Ht� ��f`vW9i�j�����$�rݻ��|�����_�]�����'ۡh������zJ�!H��M�Nۦ�E�NK˝f�Q��r�F�w�k(�Wr�~,(1��w4���cW_��[��!s��A�,�J��s�i�?M����¾�T���C����cX�1�;�j[8�^�KsWA^O�9HL��^�6�M���i���A~��W�~E�]�zj`��ᗴ���A�iN$��`$;'�6z�O2�z5ƛK&�5�l�ͻsC�`�F��vwF��yy��@����9M1�1�Ʋs�S���r:W}�g��{eKZ��K���X2�c�b(Iw�r���۾�����s�5g�$��ShM=�LWn�v�
�`'7UμѰ�w���.Nf��%ۦ�>qt�_����D󔀄�1RU�ټz��	���Hql� ���N�b�i�0��ڭ�cE���{Y�2�:�Ju��Y'X9��b�&b��=ǭ�>��	��'�ڪge>�,�#'��΄� ۜ B�,�w�Y�N�X�R���Lhb�v��\���\���X���=՘����TˆC1gA��t��Уc'qT,��{OI��(,it�~mE�8EF��[�YmD���`?y�����#�ku	٤��&m�l&�V���B�w9��m��;o�ĸH������C-��ZAzp��PF��:<���X��mQ�Z�t%X·{I�!�Z��m�M��U׋9�˞8����|g߮�;\�Ӡ ��s	����44�	���رV�ϕ��Oe��*w�N�ԥ����(�|�r�N?�c�Āb�;d3G��"���n�u�W*���`�����:~���7�K���I�z��;(��O���-���%ާ%*3�}�w%E�,1�(����a4�mci ���A&a���o���I��(pRj�P���4ٛW����d1#�M���F����R���Q���S�ˮ�:���[^9������[�b�qZ�zu��ź,�V!��<�+�6u,��&�,��-v.�5�%.c���F�-.�1ê����Uo�I�QlP�M4��y��GF�m��ˮ���5_�n��?���==�g=�C�7�N��K��PAC���[�{r�k&��w3t�F�p�^*��f�U���C���`x��W�T��н�Ư.J���Պsl�F
ر�oV7����lCvq�7#��)?cռ*��E�E�EG��U���x{;�#\�s�gq�e����2� �)��z1���x�-ϯ"e����<0��Γ=	��;}��34y
!����OW5tA	��Z`���Mw荷ơ�э�On�����r�ħ{��C!�bS�ez^9�WcH"@k�%�tD�I��N[˜K	Mm~���BLk�4�F-"��/w�H�U�_�1̛0=�N��S��Ge�)��N�zVRO1���F����2k��S�m�L1��{]�����[�1�lLpm�^�5�*]��n�hdFG=Lc(����k��:�� u����f�I��E�3�
5�C��s�c�n[]�]����ԇ�k��n���<^-@�0��w=X�:|b]�=���!������vO��7udʵq�W�	b�r:�r\�s��3xZ��*�l�V�9ۊ���s��R�� y)q����K��f��7���}t���4�iܠ��Bh�`�J��ݛ��f��s���n�^��k4��QR�Xi���]Χ��څ�W:tuuyY�b:���dSmt���0���|h�ͫ�@UR͚��ͻ�1��+2������=+��e�0*�>S���D�<�^۩L:�c��ǧն$�s����ێ.�+t�O4l��by�<�2��� �i�؞5ܾ��a��df�P��;	y�xO���ڍI��n�臅�D�����#^�L���X��dW�����[ײ �3E��m���lƜl4q�C>wsy3K*��q'DYz���V���������	�����A�5�5�4^(���ٴY�z�x��6�0��ԟ=�6�kdS�{�2��ql�Ӗ�Q��n�)�ٺ�[ڼi{�+Z��A����Hj�Fu��f�W��+�r����1g��G�m����k���g:�<����ohʊƮ�A?5���z K+�Y��=�eEØ��8&]�B��s/s.?;�B��8���d<s����MC&{��D ���O�����R�*����y�P��In��i#�ac 8
��V�Ϟ�ގ�,�R��3p�})�WD&I��N{��L&�=S���7����♭|��=�����V�����Y8��QR������lg*)u�n�n��UUd}��)<&ok��D�I�`(v���6c����[;s)N�ѳ(t���V�QW&���ύg6Ö��-]��e�2�BxbĻ��{��L[�G��K�N�&Wr`=�D�v_���~���!��v!�Cr�U��,�?k����m�׽��q�x�X�E�ܓ��,��:���[��8!�B~����G��Duv�ڶn�};�[���6�Jy�Sl���Ӌ�F׏Ms�w�~yp�Ѓ����h	NՎB{:�Ph�L��|BMХ~Τª̮xkU��ܹm;	O���>;���Z�3p�j��С�y��6��y�;�7B͘��.��Qa^Y�̪�J�����q�ރ����V�jg�ᝋ=0`���0}d� �bީ�ۜdRe
�j�eҵ�%�V&"r[9uSp�{[^�g�S2,J<h%��#G�(~��~^�6#�h�,'��@�K�`a����
:�~讽Y΀��ʥ��ǠYz/a��0D����
[k�dG����5_�0ԋ������v(���$�Wv8�	�v��-�8�r�5��0&@�]*d�Y�=R6�&V�C���)��)����w�"�y= ����O�3'[*�m�ll o����eҎ�҆���qN���Jz��HP�^f���5��p��b�$k%;�X����Ӳ�lM��f���r���/��ވF���uc�W��wܷj�t� Bc|{>�ncu���&b\N��Mwų(Y�X�ݤ[hF;�����c:��k�Ke�'���s�b~���Y��Kg�i�Ƕ��~�l�D<���#���"g͢�)�K���e��7��.���9@�����{�[���bS�]�3{��|?I���� �eȒ+�fݣ(k^%��P�����Mٗ\��穂����)�|�����j��!��;��Ϋ �ݔrT�Ԇ�!��G������5��ᦞ��-�8��>mo�oo<�&8ȣG2]��g8�}�G	,���uͥ)�`()*�؍����xOMn�Sh�	�>�g��Uk���[�k���]-B�>�3��xd�h�cEL(y�+�S��'��`؜��P�MJ��~����"��'��_z��%�3���Ƴdl��nn�cy���6�\�n���j���/`P�Y�9n�= ��R$ٔ�$�U�����$��[97��J2Xr[d3�s��K�kwI@~���`嵦8F�T��urf�����*�=�d
g�j�z/���{�F�ʭ�����q�*�?�t#���WW�e6��Z�W�ѻjn�X�UUT8l��ws-m��݇s�d<�+�]:��ޛxO]g��f
^�@��l�Y��m�Yj��Z�Jsb9
�����~)ޫɭ�L�}���Up/H���Nx8�l���&����=��I�� q�U���:]y��n��J,�N�t���!�zo��t�ov��>;Ҽ�0*�^��q�*�I��d.���S掯��VZ1[�kzr�wz�w&ۮ���(�|��}8��3<�ܳ1a����fp0zn����W�C�z�d݅T�C�:/bz��`3mt.}!�zHzZex��I�Ũu�v/Uw:$��|v ��,�sm=������<�DOM��;��`�6�լ!���H��h$�̽�ym�ȸ���]�/FH��)�G_��/@�0�iP���y���"F����3��c��Y=�T&��U���:�j��$�pFL��#C՞��/���Qp�D**��a�GAG[6VsN���qv�/�'�Pɹ�%I���� ��v�t��^�^)�
!HVdѝ�G�&��[ �ͩuJE|x^��{��~�����.κP�(�)JQ�Z�j�X��3L�ĭ�[3�K���w��^�Ѳ!�*��'Y�;�x<uI�$O������x��ϖ	����/�u��5Ժ���2[�����IEM6j:R�ۼ:Ƙ/T/,��p�����}����[�}C��仱1|����<+y)�)!�@A�(�[OM��h���MU� j�����kD;SA'��/��;�[3F��=̳4s�{)�Iq�M������t��pY��*E��В�w�Ĝ���=���ۅ��ʝ�Q�21�X[��ǜ��#����ŧa��7>��m���'/�nBܮ(.������<��4�l9�ޟF�웲#9S4�1��K�f�����Y<�(�0�wX�&>�dx!�a�ͯ�`��=��&ѽ�c$���59�O�\.� Ҁ��l���ZW�cb�f��pl�ν�����nɽ4��J��YC�um�1�dk�Uq����h�!�2�/��2h����#y��=�gð����z�ǹ�qnÌ+`Zm�u��KX�D�ۃ��{�X�gG3��xVj0�W�:,�E���;�B����.z��C�0��3�'�y���3����$�W'ze糯���i�4�GNj̼���|� �=,��t[�,�@Yo7�بvfFD�xYL�y9L\�~��43�T��*�9 �j�O�X�7]�F���ͻ�x���eC�x�Ķ�G�}(����}+zlGWVgU�nJ:w��7��7���3[gD�t�\X��/	Fb�p�fefm�z��.a�HV�M��i�R�d�_5=nwT�J�^ݍ��qUp@�Ƽ���n�%F�_Kt��*����8;�f��ʡeVLY�y'k��_�dRJ�m �Z��9��]�3�v�n��f���&pF݇븎q��΂��(вd����@��M�{�D�P������U��r!�+G��WH����m���9��E�ýj.���a��z��S�n�2�
|�K݌D�!�n�v��q�B�ݼ��s�o�"��L���mv �Ng���!��!u��h��v{btXѳk�G�;^���%�o�Ӌ�OGcko�(��[c;`��ЫZA��3���e�Ues�Fh%�>q���B�wXZ�kZ����y�
�wS��Q�ʄ�F:�w`o+T��M	[�8ʵ�K�~�N_8��2�Sޏ0�`��{hgU�J��j��g�����=~�w�����<���o���bj���{1�A�'�`���q&�����
]����|�:ϜM�j �{�f^�b'm�R5�3v���.�z,2y�:~�ςQe�k�=�H �c$%�E]�Z�bN��6C{7dmB�����BP���	�0L��%Tp����!����ˤ�(�T��v��fb�8�@�wkS�]T# E䷙��@�cU���lޥv}����<��tz��ݑ9�Λ��%��6�i.m؅óq�;����n��s$�'��z�w�2ّTܸ��U�Y7a��Jaͫ,݊���k�=0C�ǃok��D-r��\�����h�e+�U�v�4�a/Mk��]ha}�N)r:��[eq���r��l��JS�&`��}7����!}7fӼQf�>�R�c�/8�]��B)�gܠE򥛹AE���q!p�%J�N	n����5��
򶊉5q3j����=�4�	�S���Z�ͨ�Q����T�tz�f�B���`[�h�j`�$QJV��5�����g&mfn<%�QwNC�� [����2j^m���e4y<Ӫ���"�J\�;zc�m`J��m�����5u��w��x�0�<��cr�w����3wt��X���Qꆐ��uoŻ�G]v�6�ܸKZ;7!�kQ���bŋ��v�îP�᪓�eUY�Q!�kb��1�x��A6--F��(��n�d4L�h8�N��n�y��W��*�|d�s�^�xQ���ѣ���"�=l�
ka[N\�h;0��;�̼��!�/K8�w]�����M\�z���ɿs��f{Q��k@��tU�3��w+<,�:��.�RsO��fs���q��h�e�Ss>ê,7��e,��9k�Q�`�ݗҵU����bI�.�U�-8�'QaAo�`�l#Y��oQ�O�C4p�Ғ4q�X}���b.�]��{�^���ǉU�]a�׋��/���g�J Iǽj�U�L�=gL�&\�M.��*e�Cz
ѿm��G��6�G-��v�M�0H�ƨ�E͌ҧ=�I})&��� d��{��w��r^��9���-`�u� �:��Ƥ�䵶��ٹ]�[b�o:f�]�J���n�IL�sq��܂�]����i2�@���Ү�K,̽�*LF����>\'V`4�<;������q^ F葑�hn�,�5�:yRu,ۗ����u�d���y��Ã�Bg�ؔv���On��y��I������y�捰�xS�R��v�ꎃ+�hQ�y-�-h���ي�̝"&�/��^����r՚�@��8�J�K4�����٬V#|�_+}�k[���� �e�*c�V����.�,z��s8�Q�T���ӻ��{���c�&t���-��]tnv�f8���`Q����\z������f��	k*a�qš���۝��&E J�¾��WÈnnN���効s��r6��-�s����ሱs]B�\��n�]�n��r�ō�I�u�Hы	n�$FI+���.N�`���7er�CF�t�w�Pwv:㨪79�\��&���\(��v�˺N+�u��4H`w\��\�%1�I��ݺn[t�ݫsnj�s����wsW!�r�\�p�)9���t��J9&���2��]݈�lM΢˻�P$n�r�s��.t�5�cE�*w\ع���W#BQ����T���\��w]����!9]:n݋�N�PQ�QWw\�c���u�M�����}z��2���V��E���1��i��E��p9:����t�5
���� {���IsEJs/{��`��v���Ɋ_��ky���Χ�����4)~3�3t���Y��D�e�Q7=���׳u���z7�Q>�5�1������F��J�����Y�]ozW�{1��Eꮔ��-d��7>&;t���gAC�r#��1>��9��g�	vu�.�W�tj�� �!$A�tpR�tS�\�r��5��0Q�ڳ��6Fw �y	����UW]y����#t#DH=ɧ�L�qq����SM_d�!��<r)�}����S���9B&��.|�����j��]�6���;cd�/tyL&����_���Bf�p[�pɎ���Ю�}�7uo�ݔ㯅�Z⼱JQ�8�H��3� nIB
���	��_3*s���#��Qfb��#C�W�)(*[&��u5l�:�_I.�3!��ކؾ���?��r$v�2�,�#�y���6�__��|���<�R���]\���)�"�!w���� �!�61�ݟ�>����|ӄl�뀫�Q=�-b=ͽ^\�����݁C� "� ��`4[�ϕ^뫶�ۜ�a��֭ ��s)�yRU��(��/����l��6�JസG��V�}!�_K�wE���cm\�wz�n`�:C�i�����4z�I\�ԊLf�Z�Y�"�s�����K����wm�����o#^nM)�h�y�GT�>�&����w�����^���\@�m�� �l�>���t�5�ji���\f�Cr3s��k����d�;��i��%���z�l��t+�4M48޻�+{�mg3��u�ܵ^�m
q~UѵC'i?H�7gq���/O1{�*#�C�'KD��e�eR���1ٺҧ(q���d�n�Ŗӳ�cR�)XU��B�w���ki��|m���E�=A�I[����Άm�k0�]n�ث���n�-/!���B6�+à^Y�č��e�4��ur�9pr����4m<#�K,T�ٔ��m(�	�ɲ���τF��Y�ƫ����f��z���!��O"����S���?����	G��M���G�����߹ƿܺ���D�;�usZĶ�!Siέ'�k �t�)�K�io3.|�α�����s��}^W3[�e9M)���В��%5:۠i���;q��{Vs	� ���"X��)�H-rX������y�vP4v�%2��"l	�U�ͺ���wo#�TJS=��i���4�a�X7a���EE�GV����Ԭ�6�z�2cgx��9 �+2h��(�����9��j�������J�<��
�F�j�'�dk�Uq�JP��x�y�`��C�gy���w{Z0ꗴ4��q�\�rUv1/��t���I��oz�9b�Ѝ6�8;����>Y��O�yD�1��໱��e4oJJ-6 �����r��e�y�ں��2ُ��� �Ð�Do��5�C�J��$ut�]O��R��a���2�1sl������.�d0Z�u���Ǟ�l'����w|�jr����_z+Tp	wHՍ�a��q���'��N�ΜnL\�`ч�(��<���0n�iK�ZP��HL6]�s��j���9���x`I��ݗ�V�%u1���w=^<�;�ԶQ'�o\����Wb���./V�����'WC����޲�x�R��+�.�ֲlOI��_*�W��چ��$!8�\1�黋����SB�3m�߸�n�oCZ;^7}�/�����'*��Y��5����o>C4�
	)����b�^�Jx˨�a���*�{�?VS��t�y�L��c�w����l���"y�F���Vm��.�~�����u�a���-�i�fσ�˨�^԰un�b������(��q�&nxN��>'��G�\߲�1/������ٱ��c^x-���ԯ-�ǂRA�~������5'=�x([_���$<����_��4�oj@�8��dHv4��K��{uQ�b������?8ъ̝n�����"�������� �Ԛ+��e8vg���4�讙�p�Xvm�i1�,c���Dp��Q���΂���b"Y�?lޱ�͇{'���P=y#���W��A�
�e��xEj�n됭�p��g}���1׽�֎R�ƊJC�5A��j��n�vdHY�1�#��}[Kk�y�2\���^��c���W��\%�d톪s>�t�/�1�s��p�*��,p;n���(�8���m=[��*Z�9�P���E��3zz.2��;by����ֹ'����k�5��+}���E����69gq5��=���;84͚.;�:�Fvv���,��S�6Q��.���=qX�[h7;b�Ǔ=r_Pi���l�ײ�cHɾR�YMF�x����OOO�dJQQ��qz���h���'�t4��i�=^�J�YE�+�i.��YF��ϢD\��k�\�m}mٌ��`0.f2��1�(�4d�u����ܩ�j�s�ص3/����&�?��L7�s�j��J�+��Y�gI�q��h����"���4�{�l������F�T����n�V(�ϭ�<�����C;Q�˦�i��}�4I����`Eֶ�g=
v�M�4�C�OwP6�X��0d{o�P�$qcX<Lv	��ng��b��aWu9��nN���&���^��q����f$$HI!>D����2Uk�^������.k.��e�L��!j��ں���\v|�6��v;^޲�q�rz3e2�]d�S봁Aq	[�ɡX�kQ\}��,�0���֓S�����5�gK��]������Φ��=ru]xNW���^@��A5	ܮI՗�$.�R��t�f����#�Ф�.%�+v��0WnC���f�qÖ��.����\�n�oX)6�G�>�+>��6hgI���Պ�ל��z��%�i�+�G����?Q#��>q'��g[�w��i�5gq���^�IR�)G^���s>�gY��������n�4�ey�ʶ��o9
@����x)*�ڹ�e4��������m���ƈ����"�G[|g�e%`Y���<w�����(uP$���/�^7ѾV)���f����B�)�gI*�%�b��L1���0�]�3G��k��?Sim�-Y}>d�������]�:�ׅ��(�|�n�`�m��r�y�ڻ�3a���(��������=���#�)�c����͂������y����鴼h+`�Y���7�-ꃑ6ݐ-S0�}����W>��=E�t��)mx�j)S��s�^�}��`G=4f���f��(�ٻ�8���G6��}��X���7@o)�&8����0���g��j���m՜�#��r_��2g��A����*3us#�v�@�\�Z����C�u��j�ػ�s���u䳴29<2f�ƶoK�aM�b���\ٚn�f�;�L��p�)�����f%'�ha�) ɽ��-I	2v�)-6R�lv����@NM��W����w��*��e��[d_#�Ǥ׸�a/ֹX��J��6&&5r��9"d1�AU��
��{�6��gq"D��x-k�Oyn����h3x���Jv)�;Q�
��~IP���~����Q��w��� �=U���m#/Q��O�/t�lS���ϞA;U"�����)���7u�o#+ۑ�
HOZ#��El�U,��-@�p~����J/�b6�E�Ϫn����ɍ����䂐�:G�@��sNf5�M��]{�O�����7�������{Ud.�΂��(�)J:��y�錆2���:�Gfp�V�E[@��S�+77��!�g=OL��Y�vz��휎v����֎wUy���t�t�.<����>�����7��
�u����;�[�tF>�=#���z��}�A�!l���<��D���i�-�^5�C�"��r:� �!�d����{X6�^��?J%�V���o�ҽ*��J���5���	�o`�kC)`����'/g��5�[�#���K��vj㋺f�]�v��K�����{�d�K9�:f�σ*o?�2�����>(𹷮7�ݘ��(��+M � :�+eOst0�-�}�O����{Eh����B/�	�[C&���+���b]ӫ�	�kױ4AO�Ywy��g��#|#a|�M�:hG*%�NiJin�2�ʨd�F��V�(j�=����r�^l��n
3�����Į�Z��t�\nO�̌���yڱ���c���r�@�c��|�!t ������;6Q�V�-w&1�F䈉��׸���#'lϺ��C8����u]@E�Iڰ���ҩ�Ԭ���ḁsц4N�*x���G���� ^}��+1fl�©��W�����ʱ�^Y;� �<;Y��ط�.xR���݊��]��ps���=��G�j꽘��@�8�����\#�r�DUP���ֹn+ʜ]���SlJc�N`'a��{���:W%��Ԝ�{-��NL��&��0�?���8�ٵp[�B�Fj����2t�\�9�׳�!W�۬�#R�ܖ�9��\I�֘_nכ뛨PT^��тS����1О�nL����n3{4hk��H����ƒ�F�;�g0\��-�o.<W|��W�+xA[����f���˜Z�k�ꑲ���:���YhײWH�!du������+�[�آ9��N]佰�5�&�9mT�3M��'�u	��[D
1@�ۥ�ӓr\�v��K��E�)&<g�H�� +�:B$�Za[9������H�� ُgA&��I+�)q��[>5K���m��|ֹk��t��н�o�K����E�*���FR�R��j8��A��x�i;���+Ob^��������y��jz��UB�琮�������Y���:�ӷ1����l��C�ޡ%9�o�xo.QsВY�Q��k�X>P%��~��~���MXpF��]"3�PƖѻ�E�?�+Q������'�������i�-��������]���ߧ*e�[dR�3tgq��6y��W�~eՕ�/�oa�f��`8z���S����C��ݬ��,t�i.�]���Of�`t�حWY���Ҟ�(�FiS8��j�<'�EM�dt:W$4��_�z�~'J�����{���K���+J�k 7�L�z˨�Y��`Y�Dw*�b�Fj��.P�'R��;���%J�a�I}/��|��`ݽU�'�������zf�\t{��<X܂b=�+�M���riFk��1a��k=LGx��/j���G	��$$���0�\�S\�}y{�MZ��8c	m��F� b��)�u�3v=xH��:�ni�wa�e;���l�Mx�����S�y`ԙ^�߯�=�f��*}����{K��T�"�q��9�����3�@��N�F���y�8uq��Z����MYyWO�{m�z:n��4��X�R��j榜Ϫ�� b�&��D�ߔ�����周A� �p�_�t�Ĕ������Ǒ��z��E,�l���?NwF�Tv�f pF5h��?.�#k�t"P/	V)����vml�0���u�~2��5�\~=K��?!~I��;�N��h�J�T�nU
���u���;�G��g�>���&��aNA�pX�����&���?����������|�_/������_�j��Z�fY�1/�o7&>�������NF�wQ���D��E�٤w;�Nrq�.(�kz�f�:5|����'T,��e�wy��vc͎�
E1���D��jn�31'��P���Ȉ[o69%���;o���l�<�"����,���V=��fa
�E>���j��P�˙R��,��jv��X����t��ɨ��[����g#��Qi� X���H>Ta�����7��x﫮	A?�Ma�<��cf��J�v��Hw�A�yR�ݐ�M�of0��\��d�7%�Jn㥃x�wm.AE0�ԛT����˛P�h#��.]ٓw�,٪N�0i[G��BX��s5n��j�Ť�s�`��B_Aݵ�Q �*�u�-'3U�B�9����I�O�TZ�U��"({�H����i�Wp�ҐD8�O�iP�Mޕ�+���-�S5�;�5���� �d`9�� �{r��� �vrWE�8/�^�����ȲI�]A�Q���qj�/eJ9�N���t�u_`P��NQ����R|�����-hC]V�+�	}�t����|�9�ۣI��'	�y��>��8:��bJx�ah�J��2�X,��\#;�s�S���F/%襶u�v!�8��%Fm[�;�H���k/~�]9���L�-��&v*���Z6Uv���b��y��λ{4�:�+�kK9�����3��:TXV�R����Y���Q\�P��+�g�]߅K�;M�&��F全���gM�Y�+�+8j	Ӄx�歹�V$��'wl�,�fƝKڈN+�y]:��Iн����I��cF,��Ռ��|1�eh;����	kM�7�B��*��H�Ow^��+�-K��Ȗ�Ϧb*��8tru��p��f�[4\|��*���4�'����Om	�4,��9�Nå���ŃF�N���5xyv�O ���N�qi���G\3p��t�n��&t�D�ח/����ڃ���s�=�������w�h��s1S���
�c(���o�O2�1&{%	j���;=���_R|9�C׈��w�R��
�a�o�r��Ȉ{υ�Z�#���c�����c!�V�óI]�1D�(�w��w���w��\�T'�n�<����y���N��2��w/�C�s�e.��@������Y.����=���^bɻc�1�F�(�!]�^��lM�I�tq����T}-�7F��l?�xm��J��ٗs�up�P�����Rl*W@�Ը���&Tɤ��gŹtf��ݜis�3��c�rcnc,���←5�(�������	R��ѢX�ÅW\�ke��Ь�fb����@���(�+ ���%�Ӥ�k_oE�l]���%ֵFmp4�����=�ȳ:�s˽��}@ݹ -I'�bA?^�wQ�D˝�m�wn�u݆;����Ǝ�\�R��.nk��w].��gv� �G9��uٹ\d�esF�]�GN.�8�]wr�v+���b6DJ(�����v�ۜ��M�t]��4!sN�nEt���H�
4b��r�rܗ:˺5̛F��D�cBh�t���Gw@��9wv܊�뻺v��,X�%�����������ww;��ƓAh��A�(�6(�v��(�)9˷s�v�RM��q��Y�BBD���l�;�\�!r�E
�����~�"��A��H�#u�G~��������˨n��N�ZJ�6���Y{�:���-��5;te*��Q�i�%�Y���i��EJ��'Aq��d�LϜ((�"��_�k����I��e��ogvom%�4C���^V򴉐��HF_�������[��;�ew�M��3q�x;��nd�H������t���v4�!���sw'x6�e��s
꟟��R��-�ҳ�R�Q^T�d^J}�;�l
)S�s>����:3�CX�A��qTknN�Rb�[��r��1�v�k��&�v��eev`c-�M�Z@C�>����-�����|Ǥ׸�b-ojvH�}�j��;E��5��wG� <+46q*���E�D3���j�WMMu�^�n�<�;)ا��g;�]�ܒ�#�h��@��zw�\E���?R\�69���Z�K���;�rYŎ�+�96���T{���)�ӏ�'��:�^@?qC��6�GsiH�e-|�åޚ-����x�t�N�
�ّV�+!��kܐR�:G�@������hM�r���;����V"}@\E�m<8�;���H�U�}y_�o�����}�d:ĳ۵qQ����xOPd����Ͻ�N�E&é�#�\��mb�=X��=�H�X-H�:{���.��͎�t���1Ey�(a�*٘�,�i�MVf��״w���	�W�QB�wO�Oj�]��\�)V�&;2�+��X��;��q���y�>�\�Tâ����u�8�cǦ�����ca��7p�4*�Ϟ��n�\L��
}�ܢ3��RvQwLOl�j ���i���n�:��uw�Fcދp��-�Y.�+�bnl㶎���sc&�h�IET�Xe�k[$v��n�T�2��)�ٛnt��8C�*Dt�WMO_(�X�#Wt�X���0���s'o��n��)��t����`?q�:�G5�`�V����+h���n��f�3�?��)��S�/0pg��y���we镠9+�����*,�v��Hl��k�^�ݐ;hl�����R��VTk-�v����Ⲙ�k�=3۹�5�Mנ����3��Ǻ�sW� ʺ�~כ�	�U�3�;�+�U�)����s�aA�`�!�r׳7L�f/�}Wf�ȩ��ev�J�)x���-A��C#D˷Dыw1��|�{E7N I�nT4�A�xxۣ�j���0H�;�»�1a�V�i�kf-�%�e.o%S�۱u��p��WP�k�����L��h�'�Ì��<g��{!� b��-��(��[7u:�.C��xo٪/,�<xjD�Yk���-L�	���8���=�n�zԾf�z&��HrPR
�'�py��{���֋��;*-S�2�`�*��{�p���\��k݄,8�9�z��d�k�w#��ۭ �ED��-�� �0E3p��Ѭ���+#Ӵ�M�e�� nq�Dɣ:��z�zi�M3��r! �ͳCK�gx��Vz�o^z;;��ݙ��I+/�IK�5^{�#r�OfHY>��d���0��v�vѽ�	�7�}��\�K����el��Nn�X]p��F�0�����Y�#xt�)U�)���CT�#Q�\��2��^��YB��zz;]轮vר,1�K��~��f�OP�d����*��}�o���R2�$3�����el~љ�):A�u�f#�i�yb����(XY��^�c�nQ05sd���|�H�=��vڶ^��b2�Q�n=������F�,���-5��"Ջ��p�w��/n̔�}!Y�w�k4i�e[7�p�cb���}Tb���,#ۭ����V�z6J������^kˋ�̺�ㇶ���foJ�d+������ކ�`WLgj�[\�Z���2��������>ӧ+Ïu%=�hl����:��z��or�m~뮝����:;&��I�[��R�Ie�u�1s��h�6�!�T����w'��S�T�j�L�7�6�d�X܂b;p�h���=y��v{�!��x��t13�댼G�<���b}�HI!��)�tX��kX[^�2��X��V��yY�=%7����7k��H��Jd<�� &m��!;����_���G?]L#)嚐���=ܚ��:�(K�7���A�g;��v�ۨ����
�i��>��26Y�As�[Σ����l����� ���$/on�d�g���%Ab��� ��s�s.�����C��Z�Y�K)��5����'N�SWUF���.ʩV��� I�{6U�qWC[��M-���)�[+��K~9L��Z:��+�Fu�0�%ڼ3\��wr��Ƭ�%'���M�h�J���_hQ.��w��z5%�r[̼�F	���Cۘ�>�ɍ�lf��0(J��xg��	����AO����%*
J����9��d��h567�kNv�Q�s?�+��d�r��lF�e%`�)M�x�v�{}�s������=û!'�3�}��8T�%loD"(���%e!E�s�5,�5�n�[���.0�nϻ��m��8n&3WgT�T�M���x�|}�ۼ�/5�i���&W/('��yx����-��7�Y�̪�X�/�,�U�4��յ��R���t���8�gCy��~���Pv��w0JN))�=�б���Җ׊&���0.���Kޡ���BV*r�uߦ����S�`���>�m���4*
��kG8�������JY�0�~ͤ�^���Iٜ0���1�A}�1��wl�#�ǤۘofLf�.�d���q]��wN���3��5��і����N.�Ѡ{�����{2��2�6�
L��ö��zw��/�Ś�bj��V-��mP������X)�9:C%�oyo{d`������{4�6	}N����8B�������p2ѝ����ޝ��R�7&Hա�>�W��r�#o��j�֛�|�I�r��������v
3�~���;�] ?$��nM��g`[ֱ��\:9䃽��|y���"{yu%h"^jV��s#%��E�­�.�&�ߵt�����yݙ����*M{ �B@�C���Q��>�U춷��k��Y9}�=��p@t`]w$�%�&7x���H)W#��ܢ��y�.+���	�K*l��{�@���
�p�.�"�n�?�J� O2)�)Qw�`�v��Ϊ����5[��[8�]9"���\����λ�묘�R��.�N�%�z�*�$US�Ǻ���x\Hc�BoZu+l�o�mn��#j\��E/nkH꒗2�}�=�Wp=fCf8��B�r�7V����ݶ�+:�C�#&����P�K��ZxZ������3��.����^1���L��k�f���Muylo��QH�N�`ң�G���h7����P�g�߮�����L�Q���z+%�Q�>��Tc�W0��4��c�����1�Fd7$����&M��f�	��g�;�wr�Z�a��<��&�B5��d���=ғ3W)���S�Q�5y����A��jn��d]��.�ț����c�/%u��Á��x�l�~2t꽥)��n���i��r���c��"�/vPRi���b3c��8H�ݓziS��79�(k��f��nVrz����;��w���������B0���ZnĚۧؕ�խσ��}��^����ź�����3_��K
�g~*�ٿ��q��%���O�\���]���==�:>�X㷢k�m�n�5ָ��Ƕ��x'Z/!�kl��=ydD���)��Z��V>��k��۷W=Y����=�4"j�a�Z�5f�����vX�F�*9j�����z�`�Թ��t����PJ<�S�g�����a'^���w��DQz�[�.0Y�S�1v�麉s#?�W �w�-9y9���ڬ�vS�j��6�7+x��d�3��ם�4΁�
���4bjG*d�!��e(�O�6H6,�t}��gv�co��n��V��CQ���#Zsұ�B��w|.
Am��А3��s�W���r:�2�{]���;�72���6���lk%H0�� ��H��9���Z�H�Yӯ��YȕDUwW���{��\��RR�L���n�vd�gd�"]�n��=j˕�Fh�/$)�:Gc��΄M�Β\�t%�Cem4���ɦg���<;7�7N^�w�r�(��s����e5]弨
�5���Mmn�_\�`}�\���7�!��G�����0����粹�M)�R�5��rw����Fa�=>�YJ���5���ޯF�U�4d�v��ijۯ����흼Ԃ��0�tu�:�n0�7����1I�Zn�2"�-������ʝN���g�Gʺ�sW����[����~ݞ�yy��l���8������2�4��>��$k/�.r��B�P�շ���Th�z��,����^��C��>O��J<�{�gW�J�w8+��m�0ߩ[��3��h� <*/���p��1��p}�U������z���%�"x��bS�\��E)�oe�0Q�E^�+na��7Vj�G~h�қ������}i�d�鵖ъG��M�����Y5x�NK��Q��b�:�gΦ%®��J.mG��Z�R��}�l!�e�)��8��S;��������ͧ:9a�V�Ɛj�a8�?�.�m��T_��_xy�?0�����X���0��p����|諞��:�Voq�3��&�yJGE<l3��$�PkTtg: ��v۷�\\�)u��)Wd���^R��s#e�
��y/ߤ��C?�.��g�~�N'%-�����|rdў�j�TӘx5�y�2dH�����Ʌ\Ü��r��(uY�|���L.�w��2UOu�]�����C���A4�'fp��17�y,o����#n����RV^yt-N�2y7�6%����|+�U��k�25��5ө[S��Y
(�Ǌ��m��/s��g�z���qC��]fp-����?d7�p��}8����G���3V_��W%y�5~u�?���pM��dv��`ޭ���j�1ʍ�=��C����4�aɑ���'��vA��i��3z�_���Ɉ�l����=�&��V{e9�����qG+,\.wBN��� �����K��G��M�a��c����i&0��aH
���k~2�[�ܽTci������s;=���-��)����:@�w�5fuK��(��bA�����W���3�^�ܛ�������|+��l�*C�Q�4��
&���0-�o1rX�g�N{w��|�D��?�_]J.��q��knN�R�+g��n�򜖾x�����kQ�*ֶ�GU���#�!�1��sI�}�1��G�m�<S�骘��h��D�a�䒷ށ����X��:с���a�ujƍC����/=�0A3�c���HILcǹ�Q��~��p�����Ua�eEE��iuxyU�֫���yhA��+BQ/t�����uð;�z�����~nt�WW�tE���B����h�h�G[6S�ξ\[�o&��ݍ˚X��l����]��ĸd���h{�
U�M��q���]K�I~�ͭHf^O�i�s�#�D�ڧ�u�+Qa��9Jv��̨Agf��$�A���Y
��<�:0��n>��z�^^>�/g����{=~^�/ka�Z�K��߶����ܽ�Eo �h��wقK[���j�����ּ��@��]t�^7�Iܹ4f�s9E}v{���i��(im��}fJ�9D+�����D�z�M3�ķ�,�m��}�=#�p��x[��K 	�Z��-\�r�}4V�vW&<��=9�(�1�x�7As���`��]�v�pv�Zo�s��\��^l�(a�b�\K��o����C�U�-�.qoyK��L�[�����ct�n�p��#ף��e�=u`�FA�2�������yN�Yh6G� L�zz��R=y��w|���,D�����FخxS�i��s=��_<�G����\#y��]�+Cݼ`Mrb�����;7[Db�bM�^ӻp�Q?7V;�:�XO�ԝu��|y]�b�Tᦱ5�(n�ghL����GY�4J/b�r��.���/�.�h�A�&�s5�W��pj�.�< 
X�|I�Xv�Al�����c�:UR
�Ky��|����ٶ�9�bu��(	3�����	�铛,�+��%���p�ƺM�`��4l�o'nJ�PZ����$$��peK�3P\�F��m��X��pǗs��]�y��R�@P�8��k��foZ	.���gk
�V
q����-�07�U\��!pU��%X��OnI*V��ƥ�n\�W�Y��q�%UYC�g��)_wV�q��R7��=�,���\CF?��zX�B2&
�n�gO�q���u��@j�.H�}��3���}v�u[��VR�-`��Ū�n�S3+��.��R*�B$5�͇C�қb�:@�ӧv�ls���\
��GD�9��\�b�g��.�Q��r�F���ӣ�n	�1Ze��e���:�w�j§&]tГӚ���m�[��-�x���<jЛ�����`� ���Jt�r9w"������O��'Yߨ�d�	��ݻ2��q}d�ͬ4�H�]0h�a��:���ݺw�8��}���W,^�N.�zq��(�W�^{ޜ:�a����Q�Cw��-�Ɉ�Z��T\��P+דP.���SH�<t��֯;�j�n������e��S�{�������l�sYu�kS�ǳ� F ڲ������v��ӫ��1vd��]�^V��F�>�
�\,A��qWY�pd�0Z�?���m�,X.��4�[�(V��xet�WXD/.�� �L"9V��ͮv�s��+����^��@�K�+�s����:Ҍ��(۾��׹�^�' �0P�4ѱ]�3�Q琝���ѕ��o�RP���Q�˙�Os���ѝ������6�7���	�Ѡ7�]�rb�V�5vi���V��������{p�m/�1֕�u���޾��乗ȑ��c�=#��M��g#ʙ]��ٝ��L���p̐A0DoKw8ř �3D&ҕ�PRDd��+�W;��l��)�F�D�L��wtQ�] �Ww�(�����f�P�2cF�p(L�M�	����L�s�B]���1�!�n�㻡����m�� �dRb�ܹ�r䤘��:����q�NvcH�##;��!F,����K��QI��wj�깁��wt�b����)�˝(�$L�JWu��6C3��!�;�24�ˬ&�	#%��N�a�r���%��Q��f�	��.v�o=|}~~}����߯~~}y��9�D��q�x҆JX�0t�؂��؅
�ne�ƮF�y9��ާ���ك#joc�ۮ��:����D�w���>oW<�	��$U7U�ө^���i�A��*������Q�׌�I��%̷�מ�8��=fCf<x6�k�H�i羽O����I9�L�������5rJ4r��-�k[;aU֙�5L�n�=i�lA�q��}�`�t���}U�+�h�1A.��x��x�,ϛ��Q�B]��k�3c�G�q�:���0n�JL���閳w��-����� ������3g�Y����";�F�mr���Dwfn�p9�a�۫E���.�sݠ��Pn�H���B�؊�w�I����V7wv5��3���Wn͒z���v�r��Xs=�9�?4�餩�p�����:��Ig��#V���/�}���˞��W�l7�Ž�ܒ��Qz/��Bz��y�m�1��"$��) �>y{%7B��;Ni�g1������'T��E��lTW�_m=����됦�Ru��du�\�9�G���)�
�MQ�/�)�{�����T��n���<�f��D੽z��P%T�gj��˹D����i�m`Ed"c�C��z���L�1�~�RVž�5�|(��zѡWT3�Z�5eˢ�&:��/oTs�e�pj���7s�/s�����g�	C�OP���E��S����y�����H\�,�%v6����20�
�X�����W͇�&�K���qey:(HȢd׌����4�&��=�H=΍^5;��`Jh��ʆb�D���$���IHrMs��Z;q�ʩ��Z��'[zr#�R#:�ro��g��gB&��I.h;�W���5�V�k��<�Z6��碤m:C�1�	����:���e4Q��T�-W}�ޥݘ���/�go*Tu���zCv���H�F��gcy~ �H~T�콪�8��~^��|7�S��'�p��y7�yK��s����Q��\�YF��Tf�r�x���3r�I�@Yܦ�nʺުp��������y(�ʜ����ὠ��KӮ�/�x�6o�}^�g��0fƐ��@�]eg�Gd�S~5���>�0)t�§i���D�B�x�M���c��d�{�f_X��E��$�����O5�f v�oeNq�����+���^����99u�2��r�I$�Ɉ�K��F�g�1�©S�s�Z��t�ૡW��ب�BO�L���g~�_q�=�u��n �l�ۑ����B�/Y���l�I�ƃw2�rw��6o#�E�0c?��ϗό�ؼ��@㞢(qj��g"����r#ZU�s��nQ������C8 ��<����~�}�\��<���^ܴ�b`\��SP:�]���π���|����������c�(LZd����4��73DH��DH=ɦ򔎊x�t ��tU�fk����y���rLK�8������w-��UD�ݖW�ތf����z��O7F��6|�4-»&#8��4��zX�(�õhM�@sG�1��E������0��#n�J�H`��$���,L.�R��[˄����}T��C�\�m�M3�WH�vT�u�+x鄓z��k�I�=9��.���B�3�Y�T���<�E��jY�y_f"f�M-3'��wHW���׌��]���>�6;U���(R0zW�G�ګ���+M�FWR{���`�_��I-���C�Ӹ��� i�jgV�Js�A���jL̝J��􇲺�o�Bcv�v�͞�<~���k�\-�T �Н�Yn��Zʼע:����s��r�U��3�[�;���l��"�=��k��U��A���E띠-&�QZ�4��i!q~�����a}d�I�m���9c4�ơ�?F�l���mP����s:���j~����wu;�5wC4]�a�<�_y�gS�,�S��R�(��7;o���юf��DɆ�;�1�.$���K0`�9c�1�m���Rb�u�6���]�uFI�|��U�r6|v�t��3���ٰ#d���Ǥs�k�ݷ�۹�5�<��|Lt��=A�k���t`F�.]�(�w�i.�����<�W�r�b�D�8ϛ�p�<�G^_�K ����Z��m�Tw\ML�s�����]b����[�yHD�'�%hJ%��t�b���*07s��B�ʬ~;��ฬ<s&�������y-�*$de!�T��B�$_��.����ԯ�F�ܪ����|�{r�s�S�w�g�{Tr�|׾���=Ǘ�)jw�J���͝;��S���zzَ'w3{����{����)�7��bX
!���hԕ�ZΝ�yқ.�����z�p�Zk���������D�Ƶ~Ȱ`Ҙ���_Y�b;?3}�l��ꟛ�ɥX����r@�@�1�ڄF�CQ����8�=�3�ix�䋚u"�� �(G\��]��L.j�ކ`�����f�GY�ξ�ܞ4
R�vK����H�ǀ$�UC�۲���G��'k]�.ۧ��5�z8!9�q�5����ESuX�R4��i�l.2׭'k5۶�����"�-����7�%`s�5�y�uu�>l�䇍�5 ��k�.��I,&C:�ï�`�M\���K��[ֶ[��7
�c�W�*����q��@��b6WWMOP�S\��
�r�E-99���c�u���v6��f�<{C�3^�W�&�9��o��X:�{=97����������JP�i��g��}����ݕ��`В���x��M����J�7QTY��̒������V�Y�,��56;,��u��ϲ��4�W:#���t���o�G����%ǱTW�gN0�~�m�ڌo=} ��';tf3xE��3*+O,�+�γzCn�%�6�[�>���\[wW��;W�C��~��'=&י��J��a�b	�;�t^֫��ؾ���j�u &�#YiŴWic���^�'l��c��%ރF]�#$����`�����{\Q���_i~7����^��ZP76����U��yu�,��p(BՇ�2�Z9��ydA��|�&��k�����j��k:7)Ϋ���ngCXQB�]��&��f�� y8��e@�����:Š2�D�O��:�����X4����g����-��z�Z$�?Nwi���� ɵ&��i�<*%̌,�+�,Aܨ��F辩w�/�!�&���{uX�&Ato��V�-�4z�M<zi���P���-�c�9l��d!o�.��;:�%l{Ҟ��S�$�>Z3�C��댠� ��[g�<���ު���)�d#�f3�~�I+�N�=�֪���fZ���b��8��R�ց�4ʊ("�p�h�b��s��(��)q�3,&Gp~Ð���K8����ɧ����=o/�7�R0�b#�%�t�B�rҩ��Di�&Oe����5�Jx���f��)�
�j�m�0�%w@1A�.��.�;S]Գ���nB[�-S��Ԍ��+�4���*���FRyhx1e�0l�ɶ��0�{�2�l]���zzC�����t��g�jy�a�q��N�S�����3ۼ�/5ו�4]�0�R����mz�,���C?V����=��'_�==X����NT��M	[���z�>�����*�{0I'��9wP�4�:W�U���J�t ��Ϻ��L��,���{Wct�A��3�I�m=�\��ܨaH��n��.o=��*��^��<޵��e���O�b�]#�	�h[|��h��\k�d��c��Q�Y1�q�.�����\G`����z�2�a��j�o4��7*[	�\�x]�}�S���:�m�Vh qHJ<�ּ�O���1YjH(W������*+[����ۼ�=~��BB&��2A�L}yJy2�N������Q�},��5�?7��X+aW�#���\����I>����Yg\Af1ՓU��Vg:����Ic�a����x�@�)��n��R6�g��6C��[CwT��ͼ�s�Jf����c�M���s6��	��L�y)1¯��A�{���/S��<>߫"�ۥ.�AJ�2=�+志n|sͻ1�f��S���u����� �%�& �PRT�J�=��.�5�"�*ڈ��*o"]*�t:�NP��u�|�G:
F�\cL������)�9pB�ԣ���]��7�}��`M3�\FL:]lFV�EdT-�=sB-_,��룏�0�O*�k���O���R�7���3�/U-%��_{tq���V�ʕx��=�d�u3�}��!e�5;45W��ղH�Kkʫ)��ם4u_�&W�~�׽z1~��F�+�M]v����t2#z��]��ڶ�qE�R��8�ɵ�4���3W���t:F�/��(�ר��U=�cTzcgUGJ��ZR�(���i���`�ݮۤx�H��f6_o�ڐg�>�
����q�#Q����I����C�,���Р��6|#I�W�]�����,���ۜr+�}h��KڱWga �2z�O+�7r����{s�k�T���Nz����;�u��W�Gk<�9&u������az�JSB9���vM:�L̾ε�1f�T�j���ti8�&���*�YzT�0��N��?k~�l@���Z9��#�dz1�)z�8+�M�n�g��~��_�����5Ż$c��E����·t`F�BC�0X��q���Qg�"l��ѻ��Q=Ď,p�<v
:��yR�*��uնۛZ��#E�y���>����WDA�w��JДKǪ�D��x�gɫ��۫�y��a����C��%㣶��rB@�� ��у��Y�qOm�,j�ћV�e�M�n�O�+�`�w%N%�&7x����mܧ�<͜ݙ�\�o����N��W�N\K��H���һ��w��h��k����d��bC��@�*�����V�}V� �"��Tl4`���μث��x���EM��85�5����l%J����֖�%��]J�����cK�q���ŷ�%��k�O\z��UU�fņ#k^T��ك3�*a�,���o=���7�Uw�j�e9{�j�o��[��zy{r���=�4k�� 1d�M��U\��Џ^�9�����}ǔ�m�����5h���u}BW*�{ӧn�I�|�sx%ەg�����u��������Y֞=��P�K���wS�{n��7g�6[im�k>�� ���pB�F���S�MOP�P=5�]{Fė�Ƌ�[�1�;���H_-�X�v6����̸؍�Uh�}�.��D�g�>��ݒ;7�Q�1@�U#,��#6����+�+]�X�
j[���=χ(�ngͭ�%u2Օ˺�A�;#pu���V̻�h��q�޽oUؘ!�#^��=�f�<��-� ��;s�^�r�*��%�&�s����K��:)��9�>WP�E+�n�9�E�F��^�����+ŉ��N��Ԓ����k��pB��}H}�F��0/,����n��{�]vu�·���t�V_sӭ`�!F��M]P�:|*���tZv�vtf��HG/GO��	:	�2>����W�|_��~޽y������;�o�U[m��m�m��ۿ�}�ڍ��mm�����+�o;⵷Ym�[3[2�elͶf�2�f�f�Ym�[2�f�f�3k3[3[3k3m�V����fV����L������[,����U2�el�ٚٛY�ٛl�m�[2�f�el�ٛY�ٖ��Yel�l�ٕ�5�6ٕS+fm�+e�ٖٕٚ�5S5�5�6ٛY�R�l�^�U٫3[3Vf��Y��M�k3VY��k2�f��Y��*̵�k2��Vf�f��Y��*���ՙmo��y�Ŗ�|�ݶ�fUU2�m�۲�m�Z�f�T�Z��ک�ک��T�
�Z��U��j��j��Z��j�m��mUL��g��m�y�7�m�f�m��U2�W���v[UL����U3[m�j�f�m��uUS6�ٖ��j��UTͶ�3m���m�6�lͶ�7�v��m�UT�US-�ٛm�eUS6�l�V��̭���lͶf�el�ٖٖٚٚٛm�o�lͶel�ٕ�5�+fm�6ٕ�sul�l�ٛl�ٕٚ�5S+fU_��_�W�Һ�~���m��mm��3V�mfk��⊖�뎋;N6j;p����U��!�̠ӑi������G�������UU[m���W�����6�խ���UU[l���V���J�W�k����_��>�񪪶���࿍?���y�]�������u�;_~����k�W�?~V�U�km���i��cm�ɭ�ٚ��6�lԪ�m-UJ�UR�[m�kKm�Z�USR�m�*������UR��m�UT��lZڭ^�V�Z޺��o��_����U���6��Z��QUg�oʻ�����o���\���+�*��S�  I*-��z�b��!ZH�����_�ח���y��/ݯ��w�UUm�꿫W�k��[�^��_mj��o說����L����km�[n���[ϚkUV�|ԫ��������o�m����W�������_�ޫʽUꪪ�g�j����G��U[%0��!��
�	�LUahg�b?�������Z���������������m��������W����^_�S��_��������[��_�}��_����j������f�����j��z���^W���[{߭y�o�kmZ�~�z�����խ�km�w���~|o�?�v��b��L��n@�d/O� � ���fO� �~3�yR�%T��@�����F�)T��B�J��T� J@�P�2Q	Z�T���*Q"�"JRJ�I%6Ս�[MV��m�l��)jU6l�ժ���f�+afښ������ml��ɴƖ��f��S,e�e(V�V���el����[-�kl��P���Mel�f�f٭�m6��ɶ����bl5����e�b���jR���̴V���ҭ)m�Sj�MX�mikE5�m[U������a�T��سmVp  �רin��, �ЧZ��u��@����CB�-�;�T��J�g: i�W]n0�.�ݹEm�T�jn�����CWm֧M}��б��3��*����0�o�  q��>�
(}���СCCB���}G��hP�
x��
(P鷕�����P=-к��4�VK�v(3y�t즕��Z�4�c;s��������3
ѱQ`��jm�m+l�   ��A�Y)V�\�J�*��[:l��ۧC���������K�vV���y�+mJu��]�K��`�v]*��n�ن[i4�3J��ҡ��Vڦ�6�M6ѭZ*E3�  ���͵A�����@PXy��m*u��u�����l]·AUUjt�4�n�ڲ���db��n4u��mv�Pj��-��4ʣSf��Z�[-�  ;w��(3��]��Zv�je� 1�*7m��A��� 4�Ê�t����n�m��j�ѳjV�Z�Ѧ�Y� <��W ��et㦀k�����\F�4Uf%� ]�;kCR��. k�u�e����[�PsWl�ٶ6�Tֵ�g
��m�� <
�h6=7 ��e��X:qlԭ� �1ZQ����Xl]�TP��{�*�E)�^^��&�E=�I�Zkm��h�+J��&�� ϾE�J>�Ե�
G�y��6�+p���$Vr����PR^q8�Rvw�gE$*R��q�4޼w��iQUu���R$�E��j��64�jj����� �R���Mݵ�UV�r���'�������n��I("w<������Gz=��5�J�n�w�f�	Jޣ�4�(���oX�P)Wmg^��֦�Yu�kk6-��   Y}�U-���z�w<y�%N������7���T���W��Rh=��U�KgI*��R�{=�JPU�nz]���)���P��S�0��� ���hj�Uy@ O��*   "��j�� JD��R�  1??��� ���'}���]����#�3a�*�>�r����h����x{ݸ�����
�+�DEQO�APE܂������+(��)��?�~����,�[�ӆ�;�/[�
��(Y�d5�:5��ܰ!�*� 0h��ܓ%i�of��{v*Hl:z�U���w�r��7W�6oha�.VQaM�S6I�����
�ϙ�w㦮��{C�bZpMJ9GC�P5��ekݙF�c���h��t�����mP���Y��Ͱ�v�A	l�ۢs�a�w�U���`�HP�/1QǎY���hѺ�N�	�p���B����! ��eDUɭt���)edm[:��vV�A9�>�V�z�Rt7J�a�ދ�-�uKV6�*�B-w�T��װ�X��.���0H�.�+Rl]��޹l=���mT��U���:�i=A�e�oᙛ��b�{I�2�3���a�c&4�1Rtw
�P��#�%�Uc��F	LI%�4k�����𷈋�f��u$]�$(�D���ZJ	�.܃jZ�Q�^�WWF p��LJzl'�S�)ZB�m�,Y���m�����2�[e�ո�^Q�]�$���SmkmYa1�� y�Q8��;,���	�dD(g�Mz7Lc6�y��4�l�F�|6At+N�z�*���`*[Z�ֲ�Q��x�mc�t��_aŉ�Xw��mؖN�7�4~��@3��efn ������Tr���e�aT�Q]���h,��u���j�|��Li�p1Z���6��Ca�w� �^,����M}�%Q�Napn����WV=0�;�eu"ʺi�xtc�~(�z���];�s@`�-,|�K�H�6�4aj�D�>
�!spne��
�Ϛ�w����۫-�1ثu(Ә���f,*e;�h6[�.V��1�l�%n�v,*D4=j*^`���D!��$���	�!l;t���xa�Х�bPۙZ3+^��W%Z��Eh44�j�x��a�0 X�No��*3i�WB����SF#�Ytj���hh�*�wV��W�fSҫ"��a�ް�T�4�FjldD�����sEfc�3,ս��cP�n�kB�H�<E+�Go�
�8�2�搓W��u�!���6�5�R���^�^��4��(��UA�4��ǃ3����Ux���(R��⠘�Ba;�T;`�OJ�HT�v�.��T�Z;�VJ7�E���q*�˵�N�6�Z>F͑9���afl�x�k�	�Qْ��hڌ�6�WOn�vN2$ьP���(���*�U�E��*����q��o)��N!�U�Ǵd��,<`B�1�V��f8W�f��[��F�ȼ��'Z1B
͸@��N��I�Ss ��|j
u	����.q�V�%F��6][6sQ�cq4�7����UN���b���L#������+0ۦ*��T�&��i	��X[��e�=vT��\�P��d�{1M����@}��k�=����m�Q�#� -Hb����xF
�Փ��C��Anӱ�VV�l��n3!9[F����Gq���6%m��7�)*ڻ�*8�9y@��zM�Є��eX1A��K
�r'H����Gh�{.�x��P�h�l�M���h�����b�af�Gn'��T�#*:2�Tȃ&���ZVmPY�F��Q��c�-ʆf"�b�ߴ��(=:<r�qR9���D{�lʱR�+���b�MT-S���J��X_m)i�X��TU�DPɮ�^�J��JSo�(L!�Ӣ��]i��A�vEe��F��)�R�ÿd��Պ�XayF��۹"Z44R
Yɺ������=�����.
��;�m"w�Ռ�>t���M�A�S�ئ�ٺ�/*������˧�U����.HM�7�<S�%&l�n��jT�X�E�t��jj��H�K�Ӱ,u�n�E�-�楫���Q�U(��H��g�c��� J3jѦ�A�8�K�H6k�t�c�r�e�YA�Sq���^Q�d�>eԽ���#.#ug)zr�������h��/.�u�/j�ue�M`?+R�3H%�eâƐN`��'��Ҡ�M� ��\�N����5��4�%v�i��յx�KA�#l�蘩�x��P�/M��N�ۦ�*��Ä�U�Z%�ib��hI����.Xh����uj\N���#��x�N��Đ`�XF��ȶ)P���uR�_(���@�!�W¬�\�	of��2��-�cq�Q��b����@1J���f�.���F��8�ɳ����J�0P5�L."H�t�����Л��r���i&�Ila"�]��P�ٲ�Ď�,�6�m*Kk��:���6x�v��'wW0�[�|޴�5̈4��В�ǩ�5��h�a��m����
�i���u���ǐJ�>��ZZ�J;�ו���V��+{�w
Vf9q�.|�
Ѹo�6�,�ؐ�x wP��wh���Ѽ
��mݥe-�f+��ge0�cT��I�Ӗ�U�H����J`Ϧ-��ñ|��t��Y�AL���۳8��ּ�I�B�C#�<ٸ�@��F�{���crS̸�I�n��6���
�	��&����2���5�> 30�, ,��Uv�PeK]24�6�v��|�$��\Ƥ�K���㩠N�S6cw�e�ޙN���n�ٕ )��QX�[���޳��x�LJ�*��6�e��vn���B�1���J�[�.w�f�x�w*Y�)�N v��mւ�Q �c��Dѵ��V3C>�՗Ki���џ^�-��Zr�R�ЧX��2�J��,̪��Q�+N�5kX�b�d���8�"jl-R�
�'�`z`�Wj��%����7�3T�Ɣ U���V��f�
�ujS�˟HN��	��6�Q�$�o6<4�H�@]1@��P��&��i�����K 8�N�-a	 �vnaH�N�� i��f�ecIU�D�۫�wv�iUcnj��bi�.�۪7T�����`"͇L�U���mMb�/c�P`��p�����i:�o&SE^P�o74��f�)fҧ42��25�JG)Kt������d2��+c=�p
X�)t�;�eIl�Z�r:�CMֻxl����ˇ,b؃�\fӑ`uu �/[�A��s,��
����(Ꙥ$/7)����
���0��@���ˢuaT3)��n�I���7D�[ZF��
B�Y{��ɶ�A|�4\Í��A��J�*[*�KU���x��n�U�����o4��߆TܹA�r�hN��y���/v:e��+�����Ǜ+i�"mI�kX ^P(�ڽ�KB�)5��uOk5 �Yͳf��*P����gBk]���n"��\{7D�q��Z�Լ8�J¬�= )�X�e5�:���8���dߣx Ɏ�[�C�5�6�b�!��0���ͻ&v��]���cn��Q��1f�D� ܭI���	�Ђ�ح���n1VF���m�f
-�*�1v�f�Z@�,�2B��F~�r�����
����j8���8�,GuZ Ǵ��&�'��"M�nƉ���Ns���[�v���M?&�u[��)B�?[*l4�\�$�.2	�H�Z�Lɺ��e��@ј�&��BZ�	1�n���û6���i�&SՉE[�*�&С+Ne���ͧY
�R��#����Ev���O�2d�(f%�O+Ǚ�z�e�Ւ�rE%5�9B^�D]�J�³!��	�'�7f��T��n�j��^�S���(u���;WJ�t�jQcobܤ�f�Vl��(����fCe���R�X���jU�bګ�5�B�R��e�w�Q�bś�7n ���j�$4K��{�m�@���7���
�򔴴*�ݧO��x�T�[&��K�{ efĵ��j�ĕ��0�;d�}�L��
���`a��m���b'J���L��ۉ��VJM^l�
LB�يM#>�A�3�����Fc��6�_ ǐ�ЯWW��9�!��ʇi���a<.m=Y����L�e^�-��!�s�T[��1�ۭ�r�����`��Q�,,IӼ�O)E5x��4]����R�S[�j�2��l��k�M��Z�^�q+��TB8%��X�dU,�$��4�:���z)AX6䡮�J,P�X�R;��X�̵v��I���VqZ��HDsib���Q���e^\������78�N�n�Ҧ���hh��|O��|C"���ҲH�+չ��r�[Q̒���Tth"B�h^�XrF2�Pܺw��f��8�@�y�)�Df8&���є��]���#oU('w��	ث�6�ܙ�VR����ST�b.�f�kmA�k7f�3�����R�u�kpS�t���H��-X��h�f��V�b<�u��Z�ف
z����+�ZJx�2����\5�A� k� �tC��xIO��b��m,�,P�֤Pݬ2�Z�ab�fR�2�A+2�Ǹ)���ztY��DM㧕�nI6c�;CNc���[iSl@UՁ��@;�w.����ژ嘲n�m��H� �%�n��!XT�:ͼ]�J-��@bV�v��i�+$;qRp��9z�+��O,�Y��`жp��T�����0��ج��.��"ѵj࿘J'�e��o^���Y��r�r蠳N�(nʖ]�.7Ar;y��m�F*):�QB�,?7X��j�r9
Q��^[�5��@)+i��{EZd�B�ǰS�$��:t�fZ�;��.�1y7ceY�dW�LJt���$"3*:�8Eꚠ���B�H�f|�Z�$��Q;�5�a��]@��V�a�Ug�E�BhR��ɺ�+Hx�����ja�6i j�ɍ��d-ܑVSi���Y��4���񙩂�O�T�v+(��D@��Ch�@�����N����)[g(��Мt#��e[����<.',�7S�v^U�����u��B��Bh��0=(�8�n\�wB�!��l�Sk����.rםn�;i$��P:r*&�k$����򮚙[�TN���`p�аF��8-�64R�*���B�{�cJUlsZ2��}^��3 ��Y��G5�è~������vQ�D2����¨-��=��;�D�X�A����VȂ�7D8(��.���ݏiN�j��e�a�Sn9��D��Bv6�:�N�2�an]�RF�)9Q�X���k,K ���5f;aV�ON���4۳6�n����T�j�5��I^ҕ���Rˠ�;���F�IM@jR�䒉�Κ��ڕ&$�̛4�/C.@s�x�:�CsV^�;�2�GZ�J�h��3)ڤ6�+XXx��U㤱��%:e��rLƦ�/oGR	������uC5H�Z����/�GaI��Z� ��e
����Ookc؞D6��T�*G,,�7&'hR�yj�H�ov�1� c9��۴�Lp+6��5�baL9���9�HU��E��2f؊���f����"�j틙e
Nƛװ�o9�m���P���f�QU�[��	f����y��w3�\:e��⥶�:�jP
jb̻��T���V�|�5����D{�@ˣ����3^�Z7�Ԙn�7�҂�z�e ��m�̫E\��m"_�m�9��g�YM�[��aђ��1�	�L�Dn"70M[�k{O72�0ޤ�nn�y�jP��̏,6��^X�$���R�X-͠7u/���2��`����A݆XʱA�Yi��;��Nլ��/r5���9W�%����j�ѧV喀*�Ype��i޳!�b .�6)��"	&ʀ�E�eO��
�7�R�e-A�c�$�WnKR6��K���ZXF�+#���2i"�iMVg��k���dX�ߖ�0��n^F�v����5)u��X��Ԕ���#O�$vZt�m�Q=8��^N�Un�u5���S�72lE��(`.&�\�e�Yc!lZ��7H^��Y`=8%��!�a)uY���1j�F��U�}j�Qk)=�!��hCBܻ�j|L�i�"�����&eG��kY�ku�k�u�HuweM�#�	.�i�x+[�ݠ�@i�ʰ�gu��y@�ܬ�I�P@TF��7�֝x+0�Q����l3[!��ëȚH6u�(-���G,�а�T-U�OX�ZA�>�r����[���X��-�
�pl9W`�h��i�XK)�Z�7����`yt�?n�W����K�T �< ��e�⩅�-�!��ݦ��mI2H2�G�rB�Bݩo�YNdnk0U�r�sոĢ�����*�{���
��������tH�e2��S.�|�ݙ��aCm�$ٓ^e�1kGCJt���[v�唎(-nQ(�!/[�d,n�2֢�ʄb¼@��bO�~F]�)!*��n�-�V�|�$���ȷME�$��&.m��L��4�ĝ�cq�{%hZ�!ʼ��$�Q4��!;l�W�]��lj�u0R��w�偕�`����MK��+�R��m,�R,Ã,i}�����e����@��JG&:��i^���dj��@���5����n�EE�7��n�N[�eҰ�*�O��+��k *���ʐYu`���ܽanPd�Z��*�H��l��Ӏ	A��d�Pue�6��P�_7X��˼m���b�٫f3OiJ�X�wkI�UmK7%L�rfܢ��R
ٹ�Qq�+��\�[�9���3�
�?D�5�y�x�����t�CV��Xo��K�㵟fP��.�(�چ�����Ea�%ک�V�����l�Ce]c�1^�)j-L��t�,6���:�כ3n��E�*���g�mB$
䶲�T�i�����&��"*�(��6רo,X��/X+�vo���vf�S��={�m��*�*���R���n�3�;�pr��D��Q��t⍉Ji���.�B���v�W[��|5��-7G����m�l=��h<�ޕ����*�#O%໎a�t3m�hfL�}o_,+��[F�����/weV.��-Nۖ7S����l(>��w�Ę|$�+9	ԷN��gf6��n��Ouey��Rr���[�Ǟ`���kf�ީ�@���QF��g'�Z`Z��\'�����$X�کݜy����t�Ո��ť�7;�f����F΄b(�yU(L�1ʜf�r�yA�N�tU{b�&����M钻Yer�¦7y��,}n�&�\a����.�II����Vu˭��фUd��B��W�%���j��7�gVe8�I�fz��OLҖŹ�0�i��N��Q*0u���(�f����ق��&����_X���m^%�j6���3�u��q&�hR=�ZB�yP�䬻�)!��]`�CQ�͐b�꾚]^98u&Z�W�m�a[��+%e��vaj�u�3�Mɫ�Xvc%V�e>�jc{v���Ry�V˯df�s�.��x��w��7��H�L��mԬkN��6���%i�;X����l��\�w&r�!���k�nJ�i������5NՉ����%�N�w�G)EB��r�9�ל��+�\�f���y�f\Q�1�Y���G�%�U�瑼��gu5n+����Xy�����bo��;Z�����!s6\��K�(V���ms@���mp�����6�%���11}���Ruf��<�Q�|�J����H5�y'^3��\�w*�*����DF��O3�����]V��S�۶*�◹]Af��{x�I��v�:�u�락z�໣�"��l5״P�F������Y�o}bH���E�w:_aϙ
AU���o�VԺ�G6k�6�&rIn�lD���u��yN�Xnn���AYd����&���Ɲ�ov�Atú{J�P�v�/j��Ow:���=�pKRn��m3Ze��lN�:�V���6T�S���N��d�4�&L�\t;��q5�1,�ܭ��8�k��+�� W��[�jb �8�tb���hm+gr��,Z�(��r�mA.��#6��sG'+��w��-Z-X��������V�N\��{$��&��Ƹn���0RqЬ��Ӱ����A2Ɯ"�r
͖��wI���;��Kg#�r��KW�p�*C�K;��A+Պ�����&�;
81��q����@;�	�;�.���.�S�M���3
�[��//��F._CWMC��z��-[�W��.�K�m�"���*�gm�ǜ�>��n9n7�/4+b�g1�9�Aw�����j��P�>��\��;���܋!@D١Shcb��Y��Z۸W��זB~ypuew�:���M�p�r����\��lQ[�ucVD�j-��	՝�-ɓU$w'��Z�24�g3B���[�#P؊�7��e���%�o>��	N��5̚�zn�.�Xyd�a[�9��R�M�X��K劺�j%�۾�{�o��ʒ	ns�%5`��m�0�EK�Ğ���	�y�I�L�̺���b��w{�2|/�s�Ԥ�Z���]�$w�Y�v��g�n��k���X��˺�spW��"ai���:,S�]��Kb�vV>�܋^��p	��U�������jS��c�q�Io,�ѱt�}�R�L�'O�Ob���+%�SvK�p��C}׹}J�j�֋���9�HP�"z���r��S��R�^��M"�Z%�n&_3�1������g]jHX� �3G��r�'J�$��X`k�m�$��4��]8/,w"~{4�B
��|�]��am7Z���\��Y���]��o�\�׹W�`�����{q/r�ɵ#��R�����Al5�>��2lKVA`d��m�x�ϻ���777:�kZS��Z4LJЧ&ޝֶ�`먗TI���B�H�}�k�lB������/k�I��3g��.�3GS��,{k7��f��<2�"�+��6oE]�a�0�>��KXm����h��(�e��LN�}4sb�h1�\2�uvֆ{� �	��\�%����)t��oD{�k���
�K�a� B�H(�7��0jϮ���'=h�u멕b���,r��,��Uݔ�4�<z�Hu�fmi����C�yF��]�^q2�G�7���h���ͭP��D�Ƒ���k��eH�/"lm-�&�<E�&��٤�����4Q�8%�ቃ���	K��ˠ�M��L�]^.�z3mǀ�L�Ǹ�$���af<�D�eК.�n�`@VE�V��\��B��x.�;�ؓ�ڱv-=�ڝ���b�y
=2��H�[o��Eew�4�ݭM��lZ!�ޒ,B�������F^���a?k�\]���Q�_��R�7{����lk��{|���D;pdA����q�X/:ŧ��nt?1h���¡�f��.4��v`����f��[�w��NA����-���SÝI^�.�O��،N,%�Vީ��E�mfF�ɫP��qoM�/:�h�G��ww�����6i912�P|Vj��^���M]���nVT�z��$r�;�lT��d/�\�����ܺ3��=1�l�&cҰM�n��2d5"gW����CG���J�G.1��]>ݾ�0�{N:�P�eZL둷��Ka*���%�fnQ��dn�ѡ|n��qh��:]���Qw:����l�uR����R)ޓfϪsDj�w���a�\8f�os[�J�f8fI�{��]�X� ����|��m��Ry�G.�D-��7�귚��a�F�hqd;��g��l�ț�Z"d��z�So+��i�®���8�Z7 �O�LcƲ�MV�=��R����	�n嬝}���tHn���b�;lW�U���L�O�L⎮�W+ �Z ���eu�Mmk�nf1OlP�݅8�؀�u_�����ta{��+�w��M��ʺ		}���4m�"=|��b��w1^����Zu����;j�>iZF�t���@� ��u)����V�ܴ��K�c�6�˱�Di���U(��L1�K=�90�dJ|�B���rK%;ye������6�j�'
%
���*�O�s�^E2�:C(^�/���B���c�I���7�}kc])���^Ͷ�,s�F+_ILV�s�n�Ї8�q���W��yk켻%��([�b��f�SOqU�G��ʗ�U����^h���s����OJ�1J�^�yR]x�9�z���$�؇Dh�i=��U��X���ܑ5N�F���zEN��}��ʌ�UkF���%X��pP�a.��8\ܾ�dL��Q[��}�G��
���3�k�:oU����;z`��T�ܒq����=Pv��qW=PQ����&�3qC�B�Cm����]��w&��f�ӻ&s�[Ev[Œ��2ɥG�K8�g��nR�
{�r�@��z�[����������ܴԓo)p��`y�Q�9�l�D�\0ӧumucqδ��]j���\�љu�R�
��#��l܅f�&s<��5^��nd��s��i���`����b6��A�aܶ$��fc%���d��/�-�n�'f���2Ú��Rݬ�Bv�������:�����3h1�[��� [z�N�k^��0>�C�t��<49���,[ŗԞ�=�(���+Bn3�76�|���kLyEu�4Y��zm5-�t�-j���'t&��!�'Yz�g_L�'��IA�g��BS��	UŚv﷧7�RK���M�B���q�\��{csf�X:M�Znj�~�
B�d|;�بv��
�N�(�k%�ÌWmŭU�=gye�Y�fAy��RBs���NJ�s�H�zw^��i�H/�Ϙv�U����JM���;�`BB;���Zb6Y솺��+����*ylM�Μ�Eݘ�^s����	�� ��yv�����y�(�Ӯ�C���a�h�Ⅷv��}N�-L�(W;�k�t�26b�b�oj�;�Ӣܛ�j����:��Ol��N��(!�:yY��gct�t��j�3�I��eɿ*��/1�\��V��ŵ��'E��j�G��&�Νa!!Y�r�Sr��o!���e�:-��o��2Rw�,�Z�-�䀼�����sVaê^���jJJzd{.��Y�{��^�0Z*�WX��[����D�H��c%��2�n�î��y}�W��Al�ų5�ʃ;%���"jb�s.=��p[�V&���X��r���J�\�.�tfIo/8�c.Ur��-W�Ag0ԙT���
�·�J�v)6����ʓ6�.B�Q.�Ʉd��{ruMXv��2��zf.�t��$���]����ka�ymg[��tD6�G�>�R��T�\��.�lJ���MK���GS�V�ȵ�s�3�ZI�aΓ(D�k�Jj�C+�~��ŦyA��?�V���X�7d��E�|� ����F���7x\� sph+e�v���yJ��J��$j���]�>Wxm<�Z�~�-e�nkX��#|�8VՀ���d��|%d����˿������+�M��H^7�P5|jc]Sc˩�Ϣ��S�ˑ~��u;���[oQ
уɛݺ��`d�a5ٝX]쳩�
��T{T�5iN�����˲��s˧.i��l����L<ō�ghd�m��8�۴��zY�3~��(i�������d7��DX�*՛�Xg=�Z�%VxwkQm]�T&�
�]n(j�/�$]�؏[��s�]b��D�;�^�D�]��"����UM��I�'���)K[�+�_,�A[�i:�V�����NX۱.�tD�^d�l*{u�M]j2|�כY��[���p5�y^`�����S@ e�u8AD^�MY��éY��Vm!µ��u���b��֖(0#8���zq���(!x�Ҩ��Mږ�YdZ{[��V2��P��[:�S�1�I�RY�$��{|:�;���r`�AV�3�/�$���}�o��͐ED��(����6T"˝�
���Ogb�֖�g����]��ύn�	rY��Ks�{�F4�M=r�ev���Ǯv�W��>�*�uYs�)��
G:�<%YA{}8��]k��v� teұhv�����e{Xt��GMڿ��>�Wp=���F�<,�n����y��o}N�I�֗�r�a��Fk�\�S����}���#\ԑw�;ם�����P	̽���7N�PN�@Y���G����L��mt���V{zޙ����
�)22fWG[;M�GIú4��'�R=]t\�E�wM�.tY��;֬��i�,�j���P��ї�C"tB�)�.�Tv��k84"��p�����	�Z�Sλʷ�m�`�Qm��vNK�JhsR�]yCv�	@��Ɣ�cP�lBQ`�16&X��k��Տ�bgSSm�L��:]bx��XAp$�5��'��We<S�վ�wc��&1w�o0`�w���}�'ZJ��ln�9aw��9^��w�T*�6ahad;��Q;�A��Uԉ�ޣњ4pL�EX��8�9�Y@<yγ7&{�;NWVNĹ;�����j��,ը�`$T���w�f��Ҏf�gk�;u�րo)nQ��R=eC{R���0U����lV�,�� q���ז-
��jyjV�y��R�%�I�f���Jv�P}iv:��8��6U����J��$�`�W��s�&��D莚���]���ec̶o8rn��v��N���z�-sEdfT<)��E}+-��h=N�����c� VKb�W!�e�M6ʼ���ƾEZ��Bm�0X� �>>Vm��n�1nf6s�Հ7Y��� �mq�N�ă�.��G+�CsD/�̛ �=e跪<�y]rY��z��b#N`-־����C�Z'Laٺ�����d�V������Rcn�,��M����N��;�0�~�ݐq�m۹�cg��G��������*X�^�J�y@s^p���e+L�����Fht;h���d������0[h����y�
J�^����X嶩�M�Vg����:��]T��Z���6�Ԩ�B���T�xɭ�pc�@7�$�;b:0����� A�@G�21�-�6O%�[� ��`U�V��4!|�J:��;o	�bv3m8r���Z6//�ZB��`P.��QGZYaSn��{E����V��q�$9i�����Y,�S^E��5x9�3�bv�.�[qu{M�WO&�`[̏���g���I�1�T-�{��:;ᜬI� z@�ֲ��r�p�ΛsV�푥��X�V��n���N�Iv�;��|��w��6_jQ�YnnW_U�Ί�k2�Y+��V�4g^�
;�h�46��)m����,�9���Dh�9a��&�PbHf������n���Fδy9-}�g��[ڰ��_u�����.u�5CMV=�W4�;��w�XAcz��ظ�^�7p�P�lt2����uh����;j����=����X�N� "5o9Nj%d
��c.M[mI��ۻ}^̉kd ���� �\[)w7���ͽ&kw�e��-l+�*��M�^o���p�y[Iq-�Cr��Wqt�XTo��[Aٚ�v�㚲^_a���w���Y��o�l��Tġ��0^U�^}�bɧy�{�����Q�b�v��<����g6�o{c&��*��F6��͉nS�� ���Z���g��ߺ��tf�[.;�8�<	+���L�<�4���r��v�n
�dI�M<5��vZU��Gx�ٜne�wZ\�5v�5J=ε�`�A��2�YBc�g��C8PQ*�D��P��{�EWz�C0d�.9Ә��r�yķ*�y?j�=���E�9]ČBw9ӿ�T�*��A���μ�_-������i�
�և���&��`�I�������y5]����
}؃�`l��P�=oz,�1�]�M�v�;P��Q�ơ%�x��k'De��%�&��"�=(�(S��z�ғ7|�+����a���>ww���w��Ξ��5����P��+p8H$�íh˧�!���i�d�*�+&�og5+R���XD����H �f�X6I�L����x3��Q�01V'H"FY"݀s�!�/-��5�=�P��Ŷ+Yˆ��*�;�0�x�PE���9r���Gֶ��X8��*��7ءu�zv1�����%֐�i��ܔoq
<��Q]��F����_FM��0�oS�f1Y�5��Z��v���(�H_
Y�:�7(mf�Tr�T+1�E,���{��[�=���u6��v��8��s�vLj]+�����F �G:,����M�oE%�}���}���e�.�a�Z����0�a�fe�呥G��70\�]�����ʧoD�)��t8mI�^�3�u����f�u����	�M�T�K�:��#�WWZ�s�D�j�l=�L��:kO�Ni�u*b�9�<F��-���)��%�V�7t��=R_�(*rdkZ�r��� �i�V���$�jU��mr6���2�-M"R�]���R]6���N�+S�����YR�o
�c]�����C������sX�c6֜��U«wj���i^m	�k��o��u�V�o\�!���m��ؾ�E �=bU�E^�*��="�c:���{���.�Cک��Tz��+�:n�ѥ|,8U��;��Yt(�kE3����uo�.ƪ�;ʎ.�P�sm�G|k4��VP������M,��{BT�#�v�k3��`�۳��V�����s�Q��/�[R��{6�C
{$]��sf��;��ѻ�5X�b���xbǕ9k�]EIv
����7y�4X�=7+.h-w*V���5�^��F�H����UC7���pWC!����x`�X�4r�SM��s2'��P\c*���[���*ur�c�*�퍣&���\!)0ᛴz)�5��YR���x��r��������8�߳�U���Q�p����'�n�:Iѹskr���F��4,�=�%�ڗG�V��h�LDУK�׶ȲrA�w�������(;�Y�-=�n\�1��ζ���h� �Ʒ��U����1Z�u��+bo)�^�� �Ze۩R
�
P��LN���/���e-t&͐��V ��fu;�ɑ����^�N�7y�ֆ+�J�TQ_;�؜lu��F���X���?R"�Dusɠ�ϖZy�@IC,�w.wsN�
�c݃8+i���X[(Wp�sVa���x�'6ľ�ܲ��/e4;E�v�M[.d�Ў�;��i�\�Y场���%[�`�>��j=%l���B��ir�{N��Ww`P��Ρ�*�xe����w�b����8�������ƶ����p�ŉp�E\�촍h~�߁�`��ތ���*�`�<r�W%w�����U�xE�9]k(a���2���O,��YU��kܻLU-���;]]aZ�����"U�N"Cm)[�j��:�5C�K�hv^K�ݡ�&]��mVΡY�� :��q��<a�ϲ�l���/^|�2��������Sq�,xN������e:
�VnnjTO0~�3� d���f
m���u�G' 򵥵ʚ�=&�^�ۅ١�|���/I�k��%�خH5�)*�#�xM7)�1	�^�T֓s~���ƕ��w����_-%�b5��_$�W|��%>��}K�C�R
�Y��( �n���+s�c���6�ra����_vd@V��/�j6�N���LZ��ۙ����<��uuc�Ֆ f\�oxDY�v3g=J����,�f�f�� �Gp����	��M��G-��
��\n>��B+���b��'��A�u��@$Y3���jT\��r�V�����#'Qޕ�[ñ3WR���Gtx��z��Y$��-�W=v��D5���7�.���8,��g�>W�9Ͷ�KP5���/R�V��G\�19�}�W%HLi���W�.�^Ɩ��ԩ�CL4hԷ�ɴ�bn;�g��;�5۱;��9_s#��V�Tz-�7
��<N��<�li2z��*}z]m�|ҏi��
n9�x���۫`
:�]��GbhQ�7�0��²Z��8���,ӑ�,�%�Z�����}�r�]�KR�8d��W�Nn������lR�ZQV�k�F��0o
QDw]�b�rl=,����]S3�j]$�� /0��l�-Av�H�Lv��D�
���N�w:�=�)��F��a&"}���{/-�{m����l�bSˑs��nᣝ�1�3WB��=�Fְ���Ϭ �<��|���gt�ck�����γ��\/a�l�[X�^ժ̳.;�I�]f`[Aͤ��rI�a�b��DyM��
�F���*
�Znf�1"E`H���-��<�/	L��}˖�nl�-Dq�tD�`����71>�Tc]4����/ �as*� ���[��q��4�7�+��BҘ�uV�,��u�e��P��6��e^B>[��aw�"�O2��p60�wM=t}Q�4�V���:�xf�'NUq��7s/m�s��]1U����(�_)�ٸ�"}��,j`Y�@�v�L�k7q�T�!�x�g�받�vtZ����W��NN�3B�\t��"�Q�}�b1�^���գ��V��K)��w4!�,�VA\B��+{�f���0%��p`���E��Q!q$fXd�am&&l�� ,�+�u�}�C������U���@�9wq�j�dǛ3��m�ycN��-dQ<��.Y��#��_Z�MiZ�J��Fȏ�!o:�]L|�ջg�sC��:\PК��[(f�%���X��֪7�B�ҫ�O���&�������{�!3��Q=���c�r=�l�615��gh�jYX
�3�\h�7Ko�k�	I�CF.�sV`Y� v���!9m�1�Wq"��z�%�v9��c��ܗl�V��V��D�]=�M��
X��wnL�Y���q�HVv�wwGc��gE��P���[������{4WV\�`�G2.��Ǜ�h���e�*�hgmJ��i�e����Z"�_.��/1�ܜ�A��ove�o[#p�;/*G�N�w՝��%ΩS��_#1�����.�w:y(�N	��@�tm7Yo�-��{:;V��L�K�IV;&WWV�.,]�1b'��\�7�X��������eڵ�-�sC"@s���>K��D(9��ћi藼 � /��	��ogEWw�M՘�W5�q-��hj*�WCF�vw�\v�� �@u�B묙Y+�dK��V����Mi[�iE�%@�W#�%��܋�vElJ��VX�2jփ{r歹q�֥���6�r8��Iz�$��Lʱ+�.7�+����˥�#i�6���9uk��d�U5�rO���$�v���L�-�X%�,�J�ۛO5�!V�s�o�)A@��`����b�ZNH^�ث{��м�-�8ݮ��aWR�E)��ʙ�B}{@�ٲ�i`u�/Y��/*W�kS#4<��`���h�h�oI���pƵ�������9�(��TvҒ�ջ`ʹqߝ%��٤`��/
<��F����|2���IaIt��aJZ��1����T��ה����B����:
Z2�a6�;���}xw7J�WVt`���^ �)��"�FJu����o�ao&ΤK5�<?;�D�x�^%��R�MQ�F�{y��G��F�Z���էܘ�[�Z5']x��3�Ժ��J��fW�,ͮ�p�� �۷�XU��i��k:�
�4��صt��U��h��5K%w���i�'b��P������[,��t�ñƥ$i\W��%d�3����e�L��j1�Vh�[���5tޘ,h˳��n����AF���ڼkt�r�x�;ʞ{�葠V�A�b�[�~�*h���G:֞�M����]��X��C������/r�m�CE`ު�����Ll,�%!�ڨ��X�@�}ʹ�ï�<��<j��̴Yil%�����\.��Y��H���!�nIsL�p2�p|�k\�۬p�G��b��U[͢s�Vw�많�iWbLh�UXw[�j�*d��N�cc��yeE�4͓�����U��E{F�!TN��6 )�m��Ŋf\�,C^5�8�Y]*TysyJ� �l�\�)�)�*P�NN�R���ϪiVqNP�|Xˍ��nrѰ�]B�5�@��)|^���a@q��%��v���pvu>-vb��p�6�wl��x&)�i8�*#�n2{�����5ۣd�}/I��=U�_�)Y���k�o�����:ZV�,)t�Y��5{h���/3����(��Rȓ|�D�5ګ��_IF�$���]=2T���탯��Q��Yq�M��H�ͽ���Î
�<ΪT���;r��j٧�pY���wpqd�ėR᤹(�G��M�*X�X�K�3d�l��N��2�C2kR���V�<M�!0F��P9%XhZ����7��o����æ+]Ŷ�Uf����o�7��P���88#�&��s1�/y�R��Yi�ͺ�f^�L�ӵ8/&5��`�E����������k4��`�c�ȺIBgۂ���I��	LJ
�b��-z f���P�5�� 5�թk�Pv��e���r���j��V]��<g�9#dG�b�ɽ��]�9���34,��͈-�}!],Ԫ�>%ι|ìY�6�n�`�Dم<��i�j�Y��\X=�`�҃��]�������a:5�����؝�a!m��	-hj��艨�7�:�+����v� J���\U0���0e"��N֗�k�텫=.9��G�΍p���=A�u^��b��(�I 3�Q��}j�:�,7Ɨ1xW
��H�]�M�6�+`����+r&�o�S���ҍ�*]���swR���5]�;sX�aH�ڔ��Qro���C�!���7���
�������yv��+o��b�hw`�Qy�$�������:���e&���3 �T��M�D�
DP��6�VM+�ۡsr"LA@��=c%���y��_i�r�R���xf��9�b�\+�����|�][�Cb���������ݽ��[Mi��͂W^Q��#�4���������Y鴃���V�/�̎���֩^�h-��ѻ��@qph;6(�,�c�z�æ�q��K��-�=]�����PO27������^CN���v+��[�e�F�����6���@�il:�i�����xv�]���ԧ����s��-:��h*�C-�#h�V���;�-�`t�NmKy�k�зw��s�2�4✛�܌�Eu��f�fc��dQ�-H�{�-B7���a���E�u��Sy��M__Q�/ʍ����didVn	4��;ypB����\�
�6��㾅�n�Ҍ���H�׵{cT=*�N�Jڙ]� T�=�&��FA�h�|��l��2sN[�1�b�cQ6;+NU���n�]�k�l�|������J�l�5e��_�3f���1�j�bi�H�]X�+�*�����9&Psh��]�w���<�c_c6��^�A���Ս=�"	�u�-W1���w~SE۳�(���F�ls*�{�3�V�:��\�rJx6�h�3wP�Bf�޳X2wN�}xv_>gk�9��sb!D��[О<�f|(쵗��չ�[�S&����� �yhe�h2��N�3��L��^��RXU<�(NśBF��p"��ͫ2uKU��[F�Ưeˁ~7�Nj � �54�]{�.Mp��&�`��Ʈ�p���ȀD*��u��i:�eەwʱ}{Kw�s}��v$�\��pr˭�i����4RYIm��˽.J��E��@g'���M'r�[U��[WCS]s{w�yӐASƾބ�mjk �����s6�L-9u�-Hs�eo7����T,W2�rh��}1����v�>�*v�L����L���3sd��X��t�!����5|���������T�v��k���XRG1�&��0I1T��6 �vN�Er\��R�SoZ)�<���'��ΐ�m�M�2��YRN�z�I��oC��Zʲ��lՒ�B�>��9K�k�qjy���gD����x�ߐ9w�J�������]�3w�h��|��/!��j	|�46�!�
�M'�����kj�$5C�)=���ݘF�j�nZ:|d6���{�(u�nc��3�]JVl.���:���,�۝b.�(�B�+�j�W�{Z1k�����s#��c,^+ؘ`vд���B�����n�e���ql�-L��"[e4���rm^�U+�A���o&�5.f��5]=�gw�x�J��U�U��؉��1�D�7��(����*�]��G]���Vrnb���2G:���5�2��n�t2�7&[�u��Z÷�vg�SR�����S���������G����e���4 �l�Q[T/����m���b�{af���f� nŭ8��ǩ�G�!�bL;<�fa%k7YvLGX��\�r�"7�j���7��1�L=v�\� +���)�M�rXe��Vd�V%��M�bR�s�qi����"��+S����24����t������EV�����	Y���+YW��뛂Ev��084^����{������Ŏ_N2��pgq�[��t���v.O����,���5��9<�SOUĜ�]�� ��B��x^ɷ\sG��v�n�gsx�/��X�\F��д�^�[2*�S��:DѲ8u���Y2{����ܮ�/y����g�����j���2���mD�W���e��u��[��1�v��}�6�W���`σ�n�r�r��7ttw7Soo5�R9��iQj:l\}�9�y�QNs,�|�����3�Vl3X���U����x�'�,��٭%G�mG�I8��\�Ō5�s�θ��i�R4�K{9�Һ��t0�a���N��X�XZ2޹�kO���}l�A`އ��6;����	�񞦢�7&��SErwW�����%�v�0u�������{(���J�/�E#��6n	�Ż;Y�j��Z����j�h�Y��]�V9�#b��:�rR��X��=��2�n�&7z�u*�^9Ͷ�@�o)�z�n<�\�X��a�
���E��N��9�#��X˥���5&0QBK3�5b���z�3�����ڜ�G�kx:^
�m��_r��xr��(������xr�/`���D�e5h5\o=�����kj_^#k~N�롵�kB��i�L-&eU�ujB�C�5�LN[��?>���q��F�ѽ;�geV]j���6f��#�$[c�d�{���=�:��w�+2E�p������}���Ѵ�J*�ѫmPLRD%PRSDѭ�6�LD�)��TPEE3�T�ED�AA3EPQT�P1U5STD5JD��RUm�Z��A�� �*"$�((b
��f��6�[B&�����TPPR�1A4Q��ڍ`��h�65-QQL�11%4@D�4QMQT4�E4CE	LE5!T�Q�ERUh4SM4PE4$�SN�DQSQP�CE�5UAMh�CMkI-4CDԵ15DEUL�@U!K�UDQ���(
M�@QQ5��QJit@E2�3J�%AMW�G�|7�A�a�MO��v�(X`grub Ѯ��֣��0Ը6�ly$�ë�|׆R<�E��@�{��J��O���}������N�4?�Y��Q��`��y��+�c�Xޘ�N�A�U�#l���� �ѕ�A�r\:���i�P�?<N����Pl��c��}�+�XN��t��g3��缮(��ߞ(ȓ��g��=�yf���F�xV�bᲅ�����k��"�?N�\ǹ[��u���_ݶ��3\4�d.��ұ�Ơ0��j
��j�/;�����M>�v-��ҏ�$�����LƮ.z�q�����GVq����N�F �Ρ��6�R��gC�a1a����E\��tc�ZfF+L�c��
W�0x㹇�t��:u[H�7;''M'�3���tB��ȭTX9ݏ�7$[<�ꇔ�p���j�U�{!j��E+V��~ϛ;��p��qtW?�5^E�0p!}��+�yz̶��F��ʙo���\.IK=�7��q/�1�::��bx�I�P�atu�#*0Y����`;7uI�֩`B\^+|y��ƈCi�\!d�*��x�A�:y��.aU����Er���)���r�s�SW�Go��*�1���؇���'o��.a$J����9�ر�;�1�HyB/��W>�w霞��e�!��ux����̧[����˗5�םM��l�F�c"yh��)ۗ��*��iń��rPj7�yQ���%n���??�Uc9�'_-�.9봎�9xc?^��!T@�(�A���>*����QP�� �ZHg%�;�N����hȖ��{,nCu�M�w��K?I%�.��gEQ�������KL\Y2���nz�}]1��@U�u�j�Q�D��1a���-�м��E^l�3��<c�����&%m:7ґ�į�+�!Q��1q�����ʠ�W����
�: ��o�N�q? Gx�����vj��h���=�fT�FX�A�u�a˰��W|�*�2h�n���݋��a&za��Y�[������C�\k�L,y�k�oxO-��[��K꺅�;�1�F���QnP;m�ٸ���l�]��N2�X8�����ڌ!i��i1y���;F���FB�AY��4$_�帇O.τ�*ח1��ש��	�g�su���@����� V�bіu��뙋�47N;ƺ{�PL��q�4h�V���ڦ�q;���l�~��D���0��<���'��#+��),��i3������t3"˝����dI�v���%�^���)ќN��t��5�Է[�kBi�o+c��Z�	J0bZ�K�P=���UY���A���S|L6M��e%���xRnnk^ռy��3��	��HԌD�ԴW-������\�J�q����m��+F��|%��Yec����߫�!�ge�W�=�&T֨3��l2Қ���tu�~��	t���R��^�$�=�,>xߒ��;FP���7���*�@�W��?��`�/
e������L+N
:[�A�Epw����E�S"j��3�2��F$Njv�σ�-;Pڸ}��b$G	�1\�����l�=�l,(� ���@�U0[�o8P�u,`��ь���9+ʴ0L�ցU��dG�p���z.UQD�c��0f	N���ef_p���{�n��]�㧳w�$���&�wH-������2�:�����S\@��c��J�Ҹ�QDg��*#1��N�#Z�9ѯB���\9���/k���pAD���)& 0<"�zWu+�>��!Fjy=�_�P1�u�)��(���/��ڙ�H��0fc�����}.�_T8��]����|���e��+M��D6xL��i٢����p�Lx�}-��b�6��"-�z!r��S��θ��v�n%�vz��-
:G5m�A��kHc���q�$��@�Օ�|���پ8�ŏfz���!���.��//;��Fӏ�o
	��[����L�H7.r�w6C�+���zqDy��;x���u�"&=�/�G�E�t��r/��"VO.�����E��k�nX�9��rܵ@y��+�ץA�b���ڵ�%��˜�q҄>�0(�XX��T�\-t�W@^4`�deQ���G�p2^��dv�eq/]�;�#����Q�0_ݲ�ݮ�6��R���Әݚ��U�2�|�j�'6=����Lu,1P��dVUi��������]��yc��순ݨ�깖N
�����@XuW^"����ε����}<ϻ-*Kvց�G���PJs��V6����O2�ȧI��\c6�U�b��`ᯄ!��#�S����U��oi`�</�RP��C+����4��p���V�e�X0Rv�KB��S���N��ϡ�+������Jxޯ+�H~�\�X�����\L1���ZMV�=�	Z>h®p\�P��������QŒU�@|aUm$V��,�Og�Ի;Q�H8ݒ5�dn6���@�/�R6�W����Pښ<��=*���w���{:�%$��R�6]�KC�39gQ�uI+�i�x��5�s&͗�xj5KK���ww��`]���N[�|�XgQa��*v�\NJ���N�wv�uÃ��s��c8�t���Pj�_j��+���]��XU�b���W�n�zw�E����DAB�W>�zf��Ng�f˘c��' F�<w#.�3Q
P"��u�2r�*�{��ۙ=iEN-�5��<!�c[��z;l��Z8�cT6�'m�3"�L���O���� ��y~w�f�{�oX����l�\7 )a�9��W�u��9j�9 �d�f��ϝ/m���;6?+Y�z�~�K��*ہm�t�"�E�iL��ҽ����~߹�d��9`k��J��@s�,��b�^������]�0�4�OFm�P��ښ��r�us��Ƅq]l��Q� pq������3������Prlt��;���v��\�����p�����0v4n��]İ�:Ҝ�M�������9f������Q�_�������f<wZ��Y�'q�\gZ��0��Nup��J���MB1`٨҉��0�t4_G10eZ�}h5��{/��I��#����nV����cR�b8��'V7����N�n��EQ�2&�:A�z�T<��!���DU�a��@1�I��+N�.�;�+��Ok�y�� ��Dl�0h7@�ٶ3��F=���pb���ݭ�f���X��խ;Q���jW�>Ba}��e�X&tp-�V��ණ�qgǺ�]Ɛ|��û7n�w���m��Q].-W�d7�L��/o��u��6�+�Q��#w}:�d˫J����8	�Ѱ�Rଭ�*Y�,���?X���
�X�5Z�����DcrE3�N�Y�zm�o�H�2-��1umg�e�{��FQd�;y�T��a�߆�
+UT#}SJ�spqQ�-�kz�x�?0�CfD�LnNV��l����I�PT+��F�8���%e[���50p�X�4��Ǚ�1�8b���ɴU�6�����(T����U�WD�����5&�p�?_ت�����P[<0s�K��#Og�f�_
��\�4�^���/��`�6��$ƢEF��S���宸hϥ�Xw�����q6��Og��04�@9�A[rpV�ޢ*��,oP�&)�3�8<_Q��u�)&���"~�!P�Z�s;8�U�"_��`9�<k6����D�������;/������Cp6��!�np9���=m�a9�(æ ЄP
�I���O� �xm	�_<W��*x=���vgIFz!��Uv��u�m��2h�6�leP�#	+�������!)�nH��*v+i��Zm�K�b�!1n���|�k�iʀ�t�F�3R.u� +�j��2�w�p�b��
�{(@��Av❃"���<���>S�b�2�^��鴏F2�gre��8��0<f��}�S�,�+'mԅaT��^Qb�YG��������;��������!'w�3�s�&��r�ۆ�l��^��|`��;#���s[
�O�1����W:�b�3e6M7�t�#!s��,��|w&��J	���ۺf���w�:��Q;�~P3<��zhp��@
��P��#,�3��s?M����$м���yȢ��V_l�?[��w����>��Xi.�;aW 6����x�W���OS��!��@=���o&������9�ѧ�<O�ϒ�,�u�g��kfU{�D
���S�~�"k�z�W��x�[<����c��<#v�G�RpdZ�LI<@�Ф��5.s������vvf%t�a�u򿴺`�/�-������E��Ѓw�XvM6JC&޿v����"$æUR;�R���b�֧l}p�:C0�چ���8��u�����ZzI�P��Aś$��&�s q��F+�.ݼ�B�Ա��KB��0 �|G�&��{+s���S͙��QG᷶5��<n�' P�����F���W�1>���n》��3��tk��mqˆt�ɽ��e�KKtf\묖f�7A6�O[�Gkd��Ϊ��9)�r�@�܀����Û�/U��L[�swo�yA�ZtZ�!�����c�3*K�^i::�g *7r��ѝV18۫�,b�#f���`9�ܩ9���N��*�)�uÉz`��uHM|�J�� G�>��h1�qx�H��c�i���iT�!ӣ6�%�p���g ���w�3b
$���JF�� ���a���U�-N�o�a:�a�f7���}n����`3L���k�d/�U��P̩�%��Q>�|j����[�P8cD�/�����7���2cy�e��UY�
����L^��-���97�^�^���XdV�d�J�b�����K��B�wt.`9���Nq�b��Kv%�Զ�GK�>�Ջ�����x��sؐ5[3��H}n��j�=��X|>��8��Q�����G/��ϴ�
�ѡV8�A���9��|����nR�W�X��U�r��5u�+��PH�jW]����tt�W���Q֯f�B��c����a`��p/�s݃�;r�b앨�F�����B��Y9mpf��?C11�^"�� AY�jwAhY��6���|�#��c{ �r㉀��1�y�S��gƸ�j��(E�yf��)����u���1o���f����J�4QK"x�um)KuP�*V��\6�u��eF�H��+f:8E�6���S�ZS��ON��*��s��)��d��GX�{g���b`�	���g�v&��n���ѹ�n%.�*g�6gc
�Jt�!�"��t�p*JuHEtuag�]|G����l�дX�z��6�`ʞ����j�z��Xd"�j�B���{w�����K�И8�z2#\L1���eB���2�m���~�-5��SG��?e��}�K�!�К�W�yU� Պ�k<"�G����]��V�<k'��a��ֆNo�u@�w���#F�H��+Q�H\��g�Ng[<�Ԋ���i\Q,w.a�Ӊ���~�\�|S����^dM��=�[u7f�i;����8y#>g[�ñS��g�斎C��ۘ�s,��Ot��]w��K�\�Qþ�D�I��B��C�,;�����[c�����Jb~����ęvN֋;	���&a9��db;_#~mN!1�r��VC����K=�̫F��Ψ-b�n��I�`O����,��B�e�A];�cna���ۄ"�<�+f���5d3��*�,����2	�O���UY�*��u��af�)���V����6o+@�a;��%'��Bcx�W�$N޻����l^_h�\�3��pޫ=̵G�me�k�n{�v+��tT�H���8�ֶ1�V���d��7�x���Jv��г�&��o��WV�wiL�y�l�˃��WuD�}�rӭ�ȾY��0��SAL�#bW���vN֝V\�JsM����.���Tk´*1p�-}�[gTa�͇o_d��v
�]w�;�3y֯�S0���N�����J���4�X6j4�a%*��{b�u�I���د�qQ���d���H
�k!��T���s��Buc{>��02��I}SP���|��Z��@]����]��q;(� �7��V���:�(�I����sV ��z��n�_).2��+Q�_�
��'s���4]<�uo�m��	�| i�Ǘ�u�6k:u��#��u��7?gmԌ��I�G2
��jaɡ��
�e�L��Y���B��vs������c�\c�l��Tƛ���P$�(]zev��t��Z+"�� }y3E+�(��b��T��s���!�u�M���������soxzm�v4�oL�@�l�q��Ȧ��P[<0_=v��r4��g쯜��U�y�;E�|Ҋ/`��EQ&�4�js�
xEB�\4d����X�n��}Ʈ]ܐ+�y��f�
�8v%F�=�6K��i�£��˵E�)�E �O�Sً��sz�QWs�xyFێ,Ҳ_q���I�.�x�<U�S�Ko6�I�Q�Egw�^�jq�&))�A�չ�V��!aA�'sk])�]XO9 �L\�����k\܇j�cUf��P��i۹Rr۶��2L4����Г�w�{$��XuW�w��B��C�X�͕y����EY�SrO +gb�K"Ꜽ9��R{f��%��̧�}���u�l���omT|;�����ӡ�лu�T�f�nN�W�x*T�F�[2J���jP��C^�W�k:�K;PU��`�q��]#�"��/�����z�=n�C����E�>�m�u+����;J5����\��V�W���k
�	�N�����ƂW����+0`�����Wgm-"�,�S�S��-;�V��e��[�u���u���fv�w��K�V�T���>
�Q���鷹<㒦]޵�ۢ��"V��*��{+w9��'>jv��,���u��c"��#iC�W%X��q�uv�a�/AU���`��
��b�L�Q��v��$h-��ǜɱ��
�̭��^�8j4v��r�q�.���wZ�M
a �'oa������4�ɳ�kc ��O�_�(jL
Qf���v�C�Gl1�V�[�Gq>�Nn��[���u_:�d(ۜY����/^��;�br�nt6ơQ�<��D3P����\�..�m�5ˮ�46����9��5�ж�%��e7��[�~Uz�am�E��>��&EoY;�Kbkek���m9�;Hu�@_	VS��R�N�P�#��Uf�[��;�d�+l��/�����v�#�#�s�b��wZ��2�d�[�h�2j˗�I��=���=�tm&o-���y��/,�`��G�Gβ]�T�c0�Wl ��ң�s@�$Θ*��ټ���U�Y�Ņy�l��wE�ux��,����OVы	;L��� .���I<��_��1���w2���e��oZ�ה.ı�X�4O�̓$ВJg9�������{i�'^gjt���X�1[Y��/bs�s;2���ѶT\E�6�6zM���V�Z���M%�w��2Md����+D�<�)���먞  Fa�S3���^���ش����v/����`�.���]�PΜ�Z�H2�e���!qwZ��2�d:'Ep6"w҆=׺!@�x�	bk2e�� �^T
���V�D�i����&���ƶ򶮍>�6�j�օ��p���.�<��k]���m3ۏ�m�}�<�Q+=����Q̖��
��5��\�92�܁����mE����s7k��0��eJw@[�i�(�����e	���r��&�rm
�;��EH��,J��1�|:R���ʽ2a��B�q��XB��ay�
�佒�5:�����*��UT ��(J�()"
H��h�*@�������*R�*@���"(����(4.��(�iB�J��*���SZJV &JV�Y"Zh��������j��B���B�*����
V�)(����
�"F�*�����h������i*%��X���R����ih
b�j�����������)H�*�JX����
j��)
(j����
)h(
b��)i)���������)*"$���"*i�(������F���"�"� "���$)
@�
"�J
bfhj�*��h����*d�����Z
)(����")(
�)("*�
��J���hZZP�!*�����1+#���p+�&��zB�ۯ;{P��́�ף���c(Mu���r��,��T닄��6}	z�Ɂ�2;v7f�.������<*�u�s�N� �%Q�ܜ�A�z���	���;v:����%tc��{���9��pz��.����w	c�~~��:]�;|�ޗ���.��'{z�+rF�V�z�
L�Q7���}��C�f��5�/#���}�N��g�?�c�%=Gg2\��ɧ���r�(|�.�c�s	���8}���������<�������|��X���q��מ�{�e���b>/�=������K�}�{O�w3�7��|�N�mz>s�P��F��0ww�������.IIt��#����~�������>�pC�1��3���߱�+���ͫ�N �DO �q����C�����~�ޟ�|��O}��=A�?s��}��˹y|��/�ܚM�o�y��|��_�������<��n�/7%�F����C�׼�>=�!���ݥ�ê^�i�]��y�ܾO*B�:��O��>��g��x�|���<����%>I��=��'��������A�rOg�x�y����|����#�?nO�r�h��'��vl��۹���۽o3�Tiwx=���/q�'�c���t���%��?������;����A����� ײ�9���|�i�]���}����������/{�&�'���"�DO��e'�s��]eǚ;��y.�	���?��:��9��O��9`����J��:ۗ���r�;�Pױ�^A�����K���>~���>A�K��{�R>����:�|'�}�#�خ�������dn���p�\��O�xu=ˡ�c���'�:�
z��c�wP�~�u>���`����)������*��|������\����_���p
��>�>�+vr�؀\���`�u��~?w��>C��Ph=>���^��9-�t%�{/�u�=��{����|�O�t�~o�u����K�h|�\��7��u��|��������)�?���#�0},DH�#w�^0f��r'_�[�Ͽ�翪Z(<� ����!טM>_sއ���9/g�x�?���p��~n�*�e�q�0}�B_���}��O�t�/���^�O�����:�/#�s/}�C#�\�M�ڛ�U�'0��H�w8T��P���6�w�9��9�SW;fR��f�V8�/u�����M�(bFn���R�l[�NƯULĭ�N�9�����o]�����;������>I�:�e�����̰�B���6)��Ni�}��G�a4���Ϝ;�/�q�%|;���{�yri���/p�>|>�z��w2��N�d�{�r�܇'��NG���������f�I�HtB��hz�P��*��6�V��K�R����{��z�K����C��<6~�A��\:�˨|��}�^_��~�u#�����K����&�!��������#�Ǉ�}�#g1�'re�m���S�/�/��������`��4?�y� �r����=�&���~�ۨz�G�����|�I��� ���_���z?��������Ο������E���H���z0ʂ�3W�vfn����<��|��{���&�C�r�?`�|��)���#�9y!�`�(��?OG7P��M�^C��^G �npt��/<���=�S�]�k���D`��Q�s�:#�
3���/�V����_�?��=�~Gq�\��}=��p��_��s��ބ�A����'qߘM=Oo�:�//#�ѧK�.Ml{.���sy���.��K��"<#�5����yz�v���W�#��䜏~�4�Pw��z�$�K�3���=��sހ��������_���N���:��hyc��^\��9|�;��/.N�%:\#�9�8�~��P�r[[��8�D!��M!�׼�#��a�w�y�:� �y�}��h�%?�w���?'��H|��u�4>���=�|���^Ǜ'P#I���>^C��=A��h���>��ٗj����^L��􈌄����ϑ��K�;���}�=K���'�s�_����/!��C����|�i�y��N���%}���Oc䜻��|��PP}�o����%��ːch�-�/dZ�Ox����X��P^G#��9���=���)�f�=��B\���z��.���'��{/ۓ�>�%�k�_ϟ�t|���|��z_��&������/�Q�=w��<1�	UŹ����<��Bx}�&>Aq�:��t%v}����w0w�S�rNG�;��:����'�u��`�%�c�z�����|���0hk��'���>@{~˾۾��y�i��}��tq�MR暷zk);����n��-n$�;�ك����׃:�+έ�<�L_�뺒�HCú�]o���`vt�2G����ju��SU�Kc�aJiPÌ_`�.�h=��+햝�����qg�"�N
���:t�����SV~{ׄ׀��~���4�\���:�����_n]���SԺ���>Gru&�?����A�O�۟0�A��>s`��S���?���>A�~�U'�����
O�Y�{/���z]��?�����r=���^K���n��9�a�������U�_#�=��p�[�|��w?��z>��藓�䝟q�>A���y]�����r�c�:���G�}>H�����i�.�ŝ���������u>��9'/`�s� ꥢ����������;��������9���M?�e��|���|��?G��N��������/*�ݟ�U~�!��������?�,�	����������a������:�
'�[��{�}�k���{/{/����O�������}�T�7!��O��cÿxs�{'#��<���%?�8F3����D���_6ʽ���V���~����<�\���v[�G������>�?e�>����R�ݤ)��� �4�\���Sܺ���=�))���(�:��0��H���"DG���H���&�fǫ��_O������O������~�BQ����z�`�_�9Rh4?n�f����������i��:���w�R~w�|���y���������q�k`��>�v�y�4�p�1~��9���Ͽ�|�(�%�t��G�8à߲������HP�?n_�� ��O��|����9/���NG$�����%R�G�c�������'c���1���YQ�>�>���[�ST*��������R����DP�� #�8����������e�O�>{ø<������������y���(|��˹y������.�}�GQ�u���.�:���i�]P����<LD��Y�#�[���������k��M?c�9w�����î��4~�����xuS�:�'�9��	���������/��O��=��y�^C�w�:����B�������s��G�>�T�b���nϭ�>C������C뿹�?c��I��w�C���v}����	��ϝ���`�9	���<�g�9�ʓ�O����;����>���^@t ���Eص�#m`�z։3Q#�k$st'^#w�������>u9�6�p�!��'�CU���zͼ���(�3���z	���f#�]s�)��4�XV^I*.9��t8�[͘��i����9u��A�.�Ω�����_t�;;�6b�7���R�#ﾜ}�)�s-�:����?.��s=��%_�;��C�4#{���u=˯��_#�_gO��!��_9��T�����w�o0�=���rr|�I����'�H�$1O��g����v�Z%�y�BU-��q��]g������/�w��u	O�䣟��������e���OoϜ^���yS�����#G����;�K��{�?t��*B�����5�X�Wf�.�㥱Y�B��9�_M����e�{���펏0{w4�]P~�C�0r~���ΰ�|��s�8{�w	Oaל?I�}�������O���G����>��A��u�)�z�ޭ2�5{�;��#O��}�{����?7��'K���}�P��/۞�6O�:���}�=��IIN���z���rO�w�*B�������z����>�ٱ�#�H��M!n9���k�e{�8=�O��?Ǟ�'U'�4������/�~?����/������M&�n��ul���*�ϯ��?��? ��?`��GS�ǚ��1/�����~�1Q��s����1~�������s��(\�.������\|���9?c������Oc�|��� �	T�s�(=��r�{罉��������8�#�%=y����~���1ʏ��򺬾����O�Ȓ8�Q��_���C�1�yS���hѣ�l�]O��g����G*B����{,��1���|�<3�J��s��sC5�tL�2�{Bw�WT浊�(�<%��*��
�W��n'f|�0< ��-���>��:���~�9y%G�u�z��"���x�Ƀ�8�S[�#���|o(�b�h��v��H>d�~����E��˺�H�8�u��b8�����r4.}p�w�_Lj���v�Y�yA�x����Zv�{ܴ��ƒ��L)�Ix���;��������	q[��թ�E�ʒN)b�ѧ�h�fEjE��)�d���p�%�ef�T��-��e����҆UЋ5����j�]����.��Ͼ���%��sM]`������qt���~a��;��\R�?�V�mMJ������>r�[Xl�"$�/:�m�&z�uZaW0Ya��S�㜆_�g<�/�mq �t��#B�]�w&.��H �+�1�Q��ڬg"���l𱼵�Gy��x|�O^S&�y��v�6�w�H�}WD������$<K}�2�-K]pђڿ�;�cT_]�I{ZFWr�yt�D�n�x��Q�~F3@J�	��ZͽU��\�wc� �d� ��MAܻ9�qB����2bً�mր��H��oD�F��+iѸ���^B���ξ������'~�֡Q�T9)��\9@�&R�<Q1 &{����7e�I��a]�H��
qS�z�q�O�����Y<ɣp۠9���!�x�y���U}t�x�s�*����*^�qm�xt-+������}�~d������R���X��pRmp�f����iZ�4;��2����{�	�Ux�zf��J��k[1^��
F�=�QS���v2ITq�,kh���h��V�70��X"�y<13/��Hƀ��YO�F��k=��hz������F�n먧xF8^,��+agh=<5ev���).�z;;�7�9�O�݉gJ�"#kgB�/eQ�iR%@�ƣ��G��N�&�>�齽�r�@��Ϻ�!\�r�����h���11��D�@ػ�6f6��p�+��k|P�9�b�y����B���>���Ea�K�N�>�)�j�ju�[�(�`��r��a�l�U��s�R��U1Z4��|.R]e�ǵ&�\˦=퓍�~>���*�@2���<��u�������p���nN�$�ɇi�	�}9�<{�*��c��N��2�cb��&)k������,^�9l��n��1zt�oR�O�<��I�]�p!E�8�<�+ _¼c{�GfT�j�(MF�l}o��3W�<\���Wcbۀ�5/f.��1|Y'�@\@=�d0���u�wC�cd����)�ske���)�Ӻ�4�ð���˖#��7^r	U"�EW2�@U�
k%�k�b�ca^�-f�tK�W\t����p�o�c�BQ'�֐U������u�@�㖲�夸n��đ�����#�gD6p���w�3bB�%q��JE.�Ó��Oޟ]V��S�l�y<ˬOS�,e)cs/��jv��������ؘ���6氪mOL�߮�b��ɭ�B�*{j�pӐƫB�8�FǛ�à��*�L�$�; �u���H����<�N�Ï��#ll�2T�K���ﾼ­��bZ� E����gF�����2����c�
�d��]���9$ �L�^ǽ7=�o�`O}2�>)V�1�:k��<wO�Wa��d;s¤�DsN��9�ע\THGn/���7G����-m�L��Iس�@�1��Չ�~�/�U�;[��Ww�aL�`@��vo�N<@�E����\��w���� p������~t���z�W�;��U��s4CI�ц�J�V�*e��ؘ����8�����u�H/�ѡV8�t�c�������Rr2з��=��=U-_���[0��ט<�������LNo�X'\�[(1PJ��:]J[�,Tí[Y��������W���G ��_5P�W2�υG[U���9�j��R�=�+�E�3xk���"�� �?:��vtgƕ� �l���(S��5�3\!�\Wڰ�[��͘qf�F�!�e����(D��dꠊ�sAF9����)H�58�b�y��)�죏�t����q�]�(ݘd��W�k�-~[P��r��vMbz��e&�zfs��A��|&�8����OޟNƕx`����V"��5"�ǑS��Q��Ϛ�Ⱥ��'@D�7J�շ�i��xk�R�n=�d��Λo:�m�x0�\(��k":��eA0�C��f�dB�)p(E����v:��ё�I��H�G�DE�����׽Z��(�c1�9��鿢ntu��<x"J�?A��vֽ���]t5�a�qh�����=���r��5%��r��=ꑷ
��P�@�bJXΩǂ�њ�b���f8Cf1�q��oMTR�c��0�i�N@����e��f��#�}w������%�3�����G\K�'�ޯ�@�L��C8�ޮ���f �-�`��u��r��'�N����R9��t�q�'vl���6H#�M��P��R��׿>��ֽ��<B}�����8(�>�'�/�Տ]'��'�}>���8�:������ �+!��x��c�r3�9����;%���^Q`JuR���P�2��ӥ����W�#T�a)����QY��s�!�Yhd6���@�@b��`iy�X����OP?&6��p�<�27�����̅�dBҘ�Q{�q����΀t�E����/fr���ʃ8�����*�a�*��}�s����@ Rgx�vey
0ӮekWq*���0y�b�Y�`�N�Z��T�eV���-�B�SU��c�Ҷ�t[��|�h3�6Ƴ�MS������hd���x���k���o�����P�o����te��ؐep�*[��]2�cs��w������໶i]�� Q���\�]X{�R�}�G�]ŭ4ݣhi1��p,����}'�'/����C�\1���{^h�	j��"�y���sE[����yS�� �!"�N̦����o�x�&�^	��bc+°�o����y�O�v6�w��h����8�v���x�-�0;�\��u�a��o3lvb8��Q盝ʯ[𭔼�xe�+*܍�q'	�eW��wU.�3W���_S4cd�p,�B�w8�zsO�<�Pق�P�s�X0�U��';����P֡�ڞ�x�a�B�uL��`�L�BkR��#��_��םP�h��n6]��n@� ^kw4\d0L�Gfr l�~�[U��s��-�/��H�9z���.���k�����,}�+�������TDɅ���ٞjv���\4dKj�kN�����q�Ipl��\�t���-0/�q��V�;���[�Ϟ����iu�ok8��=Q�ui�F��ߚ�lg���&-��ɨmց<wF1��������� YZW�AIO.�a�v)�ُ�)|�*Q�������
�dx7�a����Q}�v۶����*4����i�-L��,�V�o�Z�{j��]�Huo���5�n�l�X�+�	lh��
� w�R��x�1R4��tc��oo�o��n���fHKB��ވ��>��r��g-�X�ު��&/�T95�n��� h�b�S*N��}�/���������5klŮ)O��T�I�g(�oK�|�_���K'�4nt8yT68ŒC�p�d�&�{k�"�u��׌^� ��[g�T��xt-5�.$���F���l�q������2�'!��wyԎ�l����U�U�uF�fç��x�xb.�n���P�ޕ���3�ֶgb=hU���8����[Vpq7yE}�@ݚ�k�;�~���Ǧ�b���S*�]�g�5Jk��N��x81{�<(��m�y��z4$���J*������EcԛrU3=��s�o���z Z�r��ɲ�cٸiW�����DQD��+	�}YWZ)�>�=!�2��'A��h��a_�K,��s̾w_1���j�d���ׄ|� l�`��x��K|2&I�c�z}Y�=�	��/�p�`�.�e#�"���N]���սz�Ҋ�a�.��8gIs�<!ڮ�g��Q�s'S�>z���Lpq]�u�r��a"1��/s��zV�<0lqw�:�w
D�:]��*�@����(V��X��(�t�D,��3p�yqr�/��k�s3�{o(�r��[�ͪbZ�H*8�۬J����C�W��'���xj�nc~��b���+T��Թ�u�\K�%=�,*Z�$}P֭��H�D��.�+$̒�.(�oG,wkHb�� �X���d�돝,�M�ǵ���؜�e��]̈́Y�dh�u��	cqА�u�T��^qR�q�H4{&<�gS��S�])yvq�Rh]Qs�Z�.�5V Eaw
:����V����w� ��	���Ig�o�C]��['u�G�Z��v���\ �cTaT�v13b�<�zs:՜�)���.��hu+((E��nۡ�O�gla�E�p�q��޾��I)�xP�����XiDň��.��f�o�%us�З*�������>�p��$�����J�w�o���``�=-�\�卝NR@�}R.���muv��5J��2M�f�Q�OXo9p��&��,�V�s��wǶ�.�g�n�[��R�}�C9a�vĴ�D.���;��S �ۭQu%��U�)wQ��U�,v,��l�';�ՙc�v��w�X���L���T�k!�����(��\̢7�/ghua1�ӐN��:� ���o��BKH��F�lJ��[��@.��5�Uݕ8)ɼA�zQ���.*�,�V6��o�͏;����C3��.�ضb��{:��Ta^�CY���d���"�
t-U��n0���Y��|��^�S[���:���V����5��/W�zh8+�:ǔ�o���m�G�!�,��3�04����`�M�uv}|/)��kq�b' !MZF�KכA�pUh�0�|�V�I����+K��v�'�.����-w�W������`^*Ǫ(6��K솴F��0Rhߵg7�T��*B�a쒨��f��hl[}&��F�y|p֔Uh���j�^�b+��&���4�Ku��3-�Qa�:�d;wܷ��	��.���p0*VZx����^�r��f��D!��Ϻ��0�����v&zVT�����e/��&��q��g:r���4 �$�����y��&f�2���B<s�Z�]��`K�������te ���Ų����)�Z�<��9��K._Vor%�}D��I�yZ�
��oJKB�\���f���ۻ��0e��ٚ"^��Z;;P{+U��f�؆kĬQ���΄0OBE�ֶ�7l�ۜp:���אs�eݭ9�f��yVuG���v+��#��]trg�]I�,�\Ypr{Im�j�eA���,���F����^��;��$���7�m���v�d�+)!fm�+�1�͜=�+-{{2и5Z�����;�5�N��p�5T 	Y����7l+�ra�Nev��� ��!Kk�/��x�^N*�p:�L���:�fݬ��U@
��UU���S%-15M$EԕI@�BAL�4�-P��IE!T���UQU41P�UESIMR%%,AJIU%MTHCA@�RQ4UDQHPSE5M%)LCE%U,��SE)M%I0�4PPREJRP�T%-4D�BDD���H�%1!IAH�E4�%TU-%%MD5A@QCPEMR��RP%	E�P��-RD1Q5P4��̅%BDU#ECT R�CBLACI�P�PDD���T�4�)R4�P�$M4TQE)C�0�$T�TUUU�(�ƾ멌�2zn��;�9D0P�)ܚ"Ppw�'۪��ʺi�Yq�Y������C��ə:�sJ�w@o�P� {�x���~�M}�������q��<Y'�� w9���E}���v� :}z�(�G$�Ny���r�Y�+�z`A�eKoj�V.J5>��f	N���eb�����<�C�Π�Q��8�J�Ju: ���S�J{0FS�BiL�5� �L>����z9��s��.XzkAa�"�d��5���BN�9Έl�s`�n�	���*�"{Kf ������}]��* @w"�z_��3cx�}N�|��`3L�Ѝ`�;$Ց[2_Tzak<:�rHABMn�k��^U���Z=�.7�i\�Ή��Q��Xʫ�S{=xk&�+�,�z�{��ל�/�GV��X�:eX�|�_<���	�+'v�y5���;��-�͠�8��e�N�9��kʐt�{~0���b3ؐ5�:�ӧ�x���tU�|L�Z���k
̱�k_�Ń������Q�� ��F��l��;4�p};�>W��to��x�>�VC�37_4o殢v������]t�p��b��Y�����{�R靲�TF2���2$U�b����ub]��XX� 4:�/x܅ܼtI���n�Ӷ�Քo%�:-�u�$������������J'�PUۑ��uk��2Kܜh�z����u]�*��iW�c"�UuQ�>�">��HQ�C��'��93�b�y������|���LH�s~~�􀱻�A�/>��rY�@
�ꖍ��h�A/��pa|ǹ_��Wj�G�`��I��&�wa�/�R��P�i?[�4��l��V��ep��V��𣜇ўpug��T�{eĜN��{{"RBr3���{"�p}�^��q�h
�T~��Z�J�޿&��r0����Un�*<�m��q�;њ�a����[�����Ƹ�J�3��"ĳ��rx�v��E�;�]���
����xs椳c����C%ss��@�F<�C�v^��y�oH]�Q����l��Ucxⶮ*�X�7\���#i�nixR1�
����A���5+�DC�Q��?�iL��+zxj�I�.��<FK��x^���>��Jz���Z�����l�1'�M��P��Rÿ���S]l �S�bv5M��T�ސ�en�F �%?���aR��(��3����:�':
�No_�}]i�۞ؒ�Wi:����a(#�'*�n��B�X�:&gz��ڗ�e�6S�.ٖ-]��ɤ�5�t���j�oJ{ߥj}>O��ݵ*�yC��js.��Q���ŕ��OKn���_��S}h�͌�]��'�(,;F"��ֽ3eP��qS��K`G���ﾅ/�a�����!�uO�*d��9`k�",	�����@��G��]��im6M��>����^�.���屐ګ�d)�`iy�X�g�,��姣�֓uP���f���7��|��]���&��wX�uP�Y�͌��`s�t���:$:�]��1��=m;s*���+�)�\���=�;�Ss�I3�
��ǳ+�Q���s+Z��K��EV��m]	q�=���P]U�&�V��`�j�������v��d1����lhX��\��\}�0�rK`^�M6��J^Z��U�P�i����Ϛ���c�����S��%&���2�|��K���߳K�kj�nZ��0���^t����&����e�瑱ϖgg*������ny��LG<ޜ����Z4s�m`�
l����"'���Tg~{S'�;�]�ϸ�zsO�<��pً���Ȝ�`�?�[��0�չ��^�$�<�ʡ��uH�
�zb��ڕ�<�g#�,ڎY~��� �����2Yc�&���Hj�T�j���p��"~�3w�;�ў�݉r�	���<�+x�P1��7sq�%#HW�7�F�۠�?�3��(���\u��֓�:a�邍�x%\�5.��J�ٷbR�[a��u��5_GK��z�t�k��<-��;�����P0/(��U�[��q�Wc�f[��Al��|��Gt�� �١�"p�}�GR!�������_t;��艓I3�N��OZ��O�_7�ϔT�h�j1�}W�����wp��O��@F��Pt���]D�ʗ�imt2������Z��
�yP���2�D�ņN��@���h�f:��5d�x"��{)���93te���1P�
������-@t�/�b��UJL�D��{�Ɋģ0o ��$q�f͊T�3�ozW�O��mTH�Y<ɢې5���Uƨq��I��Uw�XEnĒ]�3�G'DT,)=��X��YUA�1�t(�/��L���tÑ���1ymICeu%�����7�O�&V�¬�4�v�
�s5�6�y�4Sο��o��eo�'VŇ��y8��{�֜r�[�c�u�_�[������҉����ژzjG�˂��M٪u[�^�����ިBٖu�Nu�Q�Lf���	+W�(��,���K�卩�{�xKޥ��0�\Cr1��M)e�b��ól(.M`�3_^��G4�4���Վ�-V��m�1vT�f��t�uK��,�<�cȯ$u�IR��c7e]Q���w�K���ۇ�>�Ѹ�ċ����TG�>�#�-K�Ln��aB3)�� L_>y#�6M�b1l�J�E��:/MɌ�(�2�?*��[�<�n��)���J����U{�8�8Y;�s�e���������ۇQ��m�g�[CgTK��㋒6=��I�4t	`{S.�6"�P&)k���,��e�L�x��T�p�M�a�C����V� ��?"2�@�WX���{v�]0��ޞy\x��yP^�^����p^p��iƚ�}�q��P�Œz��A��*c�2;��s��]�Ou5}�B���Æ�0��9�c��J�B���F���B��ZO9�@�6���\�������1>���nㅗt��s�I�b�-��	��O� 5t�;�/֬n�}*+���Wz��,���7��CP��}I:H�s�9�yXn�s�&���f6�E�W=2�^�S�j�VY�l���W8K����;n�w�9b����c�0�J�ѝFkcVb'���Ia��QJ��5�<k���b�9�����~5^�{����u��`OGn�����G2�'ˈm1��`^��2,�È�*¯�o�R=�r2)�w١��w��i��3f.�hэK�Y��f�}�v����c6s
`Xw�#|D��;I�s�p۬��(��k �V�3�!I��
疙�"3Өk�W� �ڇ�� �9|x��^�.3�FuDx�\�.�����v~�ɀ]���]Q���T��l����֨�q��v������W�%wB���nX����[@�^'X�]��,���y]����B�<F��[���)!��ab��1\�kTD�`�bD뺑Q9�3Dsk��w#��U�X�Ǹ��&ʚ�ݎqN�6jc`������� <s=�u�E���߿e��"�P�W�N����tf_x=��^����uX�v�M/x�p��_5P�Us,��Cۆ���y��f+���Vc��e���&3�ٲ	t�^7�pY|ǹ]^��^��2�[j�s�r�/9Eܼv%���pO��ޚufe�
�^�Ep��Xx@�:�"�k��˦�@�A	�Ȗ�]տ �͇HE�r��u��|g8�B�k��h
����QZ�J�޿!��5o�n��tvqw�yR�#�n�؎�E�џk��2��@-������q���2�W���������[r�N��ۑc�R�e.��e
{?WŪxq�,��c�;�f�3���"t4۶���bؐn,��`�\AQ#,˧�&�^1.g>(��϶�H;�z0P�|�v�5�����j�+��;��e:�M��ޟ��'m�h�J������u�.�o6d؄�8�+���3Dv[^9Vp�i��ގ�Q���=SX�Y(^]���#�!)ԛ�n�X�}Xf��1̬SC8�*��c��0�i�N@����%1{V^T�Y����=� ��]��Ȉ����I�>B��-���
��c"	�-�;��=�Dn�p��!�u�T���${����XH��1)�:�ˡ����|}�mV�����Y �&�޵:�:�:���c%\3_B�17(��1Ύ�V�"�]���Y���ׯ��A�iü�WZ��}S�sT�x�5��E@y���8�C��>�]�o]�m<Ƶ��y����sl�f�!�屐ګ�d,/����Lt�zm�W"��[�:���-ZrJ��d�.l;�u�n+eqh�S*�pG_'w�>\�Jr4��[��T]�H��"�A��r�z�y��#@��d��M�}t��9�)�ε"aٍ��s*�r�)�UKRn�Π���M>�f�ŃgB&/>0�����\T��$�d���H
��k!�����ת��ޏ7���W]{��8%��83o]��Kq�.�U�P�i����ƹ��pzp��/��j�5xvu�jk+{����O�z�khLC=��,�O����}�sV��Ɇtu�݁�N���'oBR�p��J������z�����S��6�EŞwGY��ĳ�T8B��B�oJ2��c:��u����TB<�%�Y}�=��Y�T���x`���dc���r�3�w��hv�Mn0H�=�>�4��u/F�&��"�&S���o�zm�J�ݿ��rEE����1r�����mԌ��Ĝ"Hޫ�a嶯��t>����L)5�ЁF�Z��g�]=9~a�:��҆8��򮬮B�y�&�.Gh��O4�;]zlo�x_EG���0�*zz9�e�φ�C_Q=��^#\�uQM�K��޺��Q3O��������PǙ��l�~�[U��7_�-�7���+7fp�����'NR�ۑ���?e|��P*J= �艉0��Q�<���<#y���Fjq��i��iX��S��;�c[��z���bY�a�����:�7�}1B�2ʼ��;�i.,q�c]P����3�.�?1a���������$n���訕)�nȾp\���}�Hs���+����W���˄��M��� Є0/�o�\5^����8TRV{~�p��!٣����0��7�+��}[j�E|�y�F�t4*�7�M�eH�Q<
��S罖�W��2=9u��iHE�����2]�_|	�u��NVu��V�Bz���˞�W��RYJVd�kz�p�oyã��g��ӆepr�����"q����o.Z���J��Ի;]dtW���z�U�1�< ����L2�'x~�1d��f8���>b�ȍȇ�s�Y�|�t(�/��L�Zh�XZ�Ze��Z�s��"^��v��پ/J����Wm�½�=�����Q��J�W�b �_��ފ�ޞ��]�)i�������8���a!\va��"AzeFW<�<���.� ��P��f{�뙋�sCt���6�]�t�wo�0���oLN5U�d����Ʀ�|�'�0['�� LE��3�V��&||*����EM���1Z5� �m��OT9��|.�%���m�V:��g��q]1�;,+%�MDs�e�����y.��:�/9"f�w���]��~�Py��&"M"|<�X:}��5Q�0LR�_+�K��`2���R�J�S>�ĸ�W��>�TjaZpQ���p�\1-o�6�2�*a���)`��e������}��l��m\>ό�?P�'�,��e�̌��+�lo��
�#:��(�/6a���Pu�x��7�SF2Iì�gaR�W�>�3��$f��me����m[�٨���M��G��fTε;���(�rչ��M�C��&�ڪ_�r�]7�����s��j��dƁ�$�D��ӫj97x��r#Gu��zOL����Z3�[,O���J�"1�]�������Ӡv�3˪DǢ>���1k��b�xvR'��e�D_p��O�$�Q�:��9N�%�=�#y�	��Wջ� EX�T��S��P�?��\����/�-�_T$�"��^Vm��$����^KU[!��0�>�ve�L�h
���F��:S7x�����'1�����c�صj>������ޭ.�u�rH>40��o��]���^:��ᩚ���#�+�g�u�!�F���i��2�d�z�٣'1����xd��(�_c�ӥ����_?a�����V��%\)ڕ�zu➋����4�� �s=ܰ	��8>�s �l�z����N����1�7�^��ts]��FA�Q���cE���9�#�k��qb�����B��x�WW����y�}]�:�g�_T;��h�1�,gl�sk��x�[��)�����z;?V��Gn�n�~�L��+��G9D��K|O8���}�W2��1���ĩ�����h�U*��м�������_��W����l�K��	}���8�=ˎ/Ҩc�
UU����kg��y|ԏP<�����E���R���N�X0��ӓ�ӶZ���(��g^�:�5)W��:�z�����s1���۲#��%�G��[���GkT:󩢚�.d�CwF�w��r�S
�e���J�!�u���ί�ü97����&�gj�Շx+=Tr��Tе�$;��A/�i;Q��%��W�c�]q��]J�ywEi��_�-�r��N�gE�e��U�۝	��N,��HV"9Ac�u�v������{���]�`�v5��Q�HB�W}.AW�,X������p�U����H���v-�a���fF�ܥ4�WB���'\3]��,��mc�(�6�MeSǀ�y���w)�L�`���6��H\��+-��5!{�	R٠/j�]H��V,���%*� ;]�hrO5���GwslT�&����i�h^X��-د,ru�۸���^LI��&KX��,�t6x��{ջ]�;�p%�qRI͖�p�9�Z��/pBD�DA,�k�Y�9�s2�%(�j�v��e���2즲9\����6P��� |%�Xѣ��q�}�ö΢�n���VfN\�Rz��0��m��Gƃ���v
�� �r�Yݑ�z�]�ъ��k�d�H�ͽ�{�s�ђ%=]ǘ)��ֺT�[���,�L�p�g<����]M�W+鬍z5��.n@�g�Gת��UK��U����/_i2�E�oP�{�jSO:�4o1��Wt��BA�Q�v�&����N6s��<(�� v��n�V$:�un楏%�����p-UF���5)���I��o��d���}4���'R�����wO����V����\H1�yY�m�$�Uoy��4�l�[�4�v�6�\X�%-u���d���5WZYx fi�j��.���	�h����<���=���+9ɠi�Tt�j�gj9c:�W�n���ݍ��ͬ����+Mu�Hr��y��=I���r�ӲU�F;�1�z��+�sM��t]���F&�e �jض���B�G/�*N.�Q���+���7��r�C]L
V�M>Ey-�5�Vi��U���o�`BZ{ډW��7s��nbR���Mv(3,����Pd��� ��I���>�b�ʹ��E��Q��v�Jѱe�(.�	��3@�SiB�[`_>�Jm�1�ǳO+�{|�\:�EX�N��Cc��\o�gf�(nU�������CLN�Af��E콌^v�A��n���}��Jn�2���6�v��X5av]}�b���}�~*?z	�[�wLzj��%
��y$��tm�Q��PͳI\��̡�iVp*�'U�q8�E��R�L��]V�o3�\�|;YA���e���U:����d�C����F�[Iۥ5υ�Z�c��һQ�r]�;�n�hsĳE�"	Zb��q
�ǌ�V�����ŒDs������^���K��*��)����))�c EDE�CVΨ((�*

i���i�(�a��R�!(*��b���mE5CM4��UBDR�SMi-5T!4Q%-)UE����J�Ԕ&�4%)m��4�����ZTkT�QMF�$Ӥi*��E�5J��AT�iLT4P15�M4��TEUPZ]ɤ"�J�j6�QF�AT�Z��A�ƍ�E�EEEkM�j-���j

X���"�ul�M,DSP�Q5�F��A�����Ѥ��B���bu@:(-��UV�UP��8�B�*�6p�8����(+Hj"����h���$�URIQQ�kCF�_�������y������)�A�l`�~�B��K��baT�|2�,���WRd��^D���CILb`���:{�� {����^��^��?�}��*'�`�T��½�����>�g1Ǟo��.$-�&u
\����tb��[�LBe3�)��g8�.ʔo�0l�~Lɞ�B���9֡�i����wS2{�eٱ�R�.��a�� ,�L��n;��@� r�: �����w�Y?C�mWSe�븖b^���v[RY�� ,=�ީ�~F�!�nўcD�@[�[|
ݒi�H:jO�q�*��V7�+j�c����1�S F)����_���e�����OUjzSԁ�h�:�2����<*���5ˊ�|}�Y�S)�o�W���6�˔c�
�=��S!717�ꙑ_)���Ƨ�co�0��x_^�%�%Q�xb�8x���;�㳭�2�e��F2z}����>t�j�q��}(-�N���y		��{'�|6�X��b^�A��d1a�O��5L��1�",����-56�k��^P�G�5�jꥧ#na��چ#�<�STb��
p�Ոv~���:�a��x��ؚ�׉������g)|=���3s�r��z�7����R�nEYl֍�s���y�̻����RuE,u���wfN�����h8hl9�����ٖB�<�rj��	���M��x͵�{1ݗ#u�}U��L~ԃ���>�����=�f����Y�6�ý���=�?����x���w�aWO0<�]a��{c}I�m�����å���U�Į}F�+B��-}�/	o_i0)3�
����E)�sԎ���%e��>�D����Mg����k*0����_�9G�82o�PAm
�Q�Rj�����GT���:�bucz�ޚ�D���\½������֔Ł57����R��V;L�T�|�G+��M���3�b�%�~�]r����t.�t���}e�"��<*MV�����1�"���T[�#��oD�}1�u#*����n���<�ҢM�w�.~���&�h`�P�]��.���?0�CfKT��wK�wؾwI{G�p?|&�Y�I�Ih{]t��F�s�e�Z��<�e��'w�0*A.��۠�=�[��.	�U�6� 10J8�3R?%�X̷?T�cr6[�QYϤk޳Ã�V�h���i냌���B|*J= ��!i"Qž�6�`OVI�������+�7�@k&��+���U���y��p�˧Wc�FS��Ȥ�:�Ygm,�F���g���-���F��ݷ�T`�FI3I��2�r��*S����Qk|�+�ΔΡ��]�pe�q�����i<D���B�����O`�ۖ���;���G���Y���MP�ﯺ��SU��e�븛���x�	g���T}�x��,��p��b=��'��^�Na�F+�u�)&�\�a@c&�mր��H��k�����Y�x���]���1��!��S�u����_0��p�C�_Bn��� h�F,��pbi��&�5�d��qr��Aƾ=?I{X*�9��q�+��O���D�Y)�E��V��3�
y�c8�+�<����&�i�IZ��S6�}��#��g[����ﻯ.Y��s����{"�V���l��?q.yp9+ޙ��*��M��U����^A^����F$���b������}�]�T���Q�ŷO�9c����-7��<�,p��{,$+��2���X�O)ϼ<�G�u�z�}wr�:�.!gY��뙋�47Nn�����~��7In5��^�Sh����z��Aj���� ���?E��2�6Hb-d�4��\Gd譨��.)���s�m��H���:NV4����?q�/��ѳ���O3��<��숋"���[S�Ϧ�E^E-�0z�,�Oewy�ZzW+<1$M-e���eN���s�P{���=Х�)ٞdc���0�߈�!^f���4syOe+,AvۄngUK�O,d����6�؎�w*>(�9����G��Y|ڱ���'3{�*��K����}�$���< �6���v�'���U1DlIȓH��X:VF��J{�]�_v���9��2��N����N]����V�	JE[���)��b���ȃ��@�WX�;�%���i�N����;!��A�o:�_�����\!��:ڨ{�q��P�Ov~+� wy " eѻ�v�tt�h�W�F��`��gU���{.q�Qưn�뭕B"���>�*�B�Ô�Xp��!�t|l�
~�щ������.����F����ꐖ����]��#�U+A*^�>0[��l�/H|ywWԓ��g6W��`7"������x˟^oXVP(H�Ńk��EQ�O�P�.S���@�L��1{�>�G;ML��u5,�#�Nlh��S��*!M��@�	����a�U��6�fj�&�����tGfg�Cb���!<�&*!���L�g�W�ǈ�Pp���"���ҳ{2Q��5�ء5GS��u���h�����$�wȰ�7,y�k��{e��&K5�#���#\Q�,}<7,��(OI�wyo5��m��:Uי�z�Q�����Z)�囻5��Lr�ˬ�5��n�vФ�,W�a�����f�\�g��1�j�7'��[�_+����n]]�[6���/$0ڶc�|&?}�x #��}>�~7%��G�Ξ��w[/ac���]k�X�t�1#]L��\�pr�$o0�����ojվ�J�ڨ�
fZ���Cu�F�j�'i.�٩�N��moY�����/L^�e�(�f����"��M��x�r�D��W>U\�%6�܊ã%EoT��޺Nve�Ȟ6ޫ��ڦ��X��#f�R\-���Xߡ�tiPjr�(�Y�pb�*څ/��D8��e��3�x���*�1��Â��e���(_�*K����d��j��[�u�*���cUXY]|�r�t')��<�3�aụ�f ��?&[�먖���{M�f��2��Udo_��{�U[[���n@�Bw��qS����]�e�]�~�o����	���U}�a�ms+]ĳ|)���gZ��m�����g�Z��p��d�d���:�\���D�d�9�����]�*��o��N%�g�ʼ7	Es~6B���%��@FZU"��4�ҙD��F�t��K��+x�/Of�nL��姺Fu��/۬{��˽��.�,h��,"�h��&�)��@��._��J���s��MwO)����;����/Ozg6��8�=��W�%��>�꺮\��Df��UX���lm��;���W9�.��G�&$#�eܮ�����&�=3ՏC���1�q��As!�17�ꙑJQ�A��b!}H�1>{μ3d�o<����`�f�<-�H��u0��-Yg	�D�'��J�j:Q;Bf9�	�0X[{�� 	{X1Q^�lc���G�t[ƔΤ�D0�>����KP�5�@d'PDON��LA:��7�'Q��
9 �du^T��;sl�f�!��ښ��2ܰ4��v�S#U	�k��w�����0}~9�-��͍�þ���\_�ƊܜܝV��@U�Mv�Y�>qMEC��s����V]�Ҷg/�]u.�늭gݿa�Z?lހ@���*��<^j��}�g�f�"��pOW�����7�C�́�2ȕ�Õ2�Y��/�/������{Q���c�w��P8uJ�ϥΣ؝X����1Q�*t�#@]�*�*�<)��<�G�({�x�>�R)"�z�B��c�̌V��.}���qߓ�;ڤ���ݧ����Z������'�]�|Ǩ�
狃F���G:��nH�y����b:��"��&A�"쭩�Ɂ�z+�yMFj,���QZ6�%�^r�efG`(8�u&eN��xw�?�u��P�<��k��sט�|����@]c�Wk���؆Xiؗ�Ɋ7iwV���w�j��F����Օ��ۂ�:��
��s@���\/BY�Ӹ�?�{�
�Kb�\&��R3�s��jJf�ʯ�6��(�B�w���i����0&ĝΪ��`�ҡe�ю')�ɉ��'j&P���eaQ��e�Z��1�աiy�m۠m�l��V�¸��pڅ�p��߁�x�A���q�g"�G�[U��OF��/,���W��o��K��r4��g쯜��T�g���zH"=���r���}wr*����Z��Έ��N�h�m_�졭��/D�	g�F3�%3��z�&��S��p�)�89�5;�l+K4ZI�l��۸C�i�ˣ!�!��y�e-�4���h0{\�]�����K��&�;�9�/�Ut�A���e�rzU�y�%{6�
=,
�3q�e�L����j�hHQW=��j����,���8�.�s��^N��Y�^�U�-�?i�O�X�"�d�;���X���V�pʋhm|�V�5�F��k�f*���U�S�j�gu�˃�rx"��;��>�w��eؿ��<�V��v��B7@�m��'P�,��fn�m��a
`���6��0��3n��2�ɛ���S\ǋd�V�9���p��Z��8���s��K�+vԮ��;��U����<��9or��.N�i�9z�ƾ{'\�s�u�ed�ñ�2_q�o9J���q/��$�q��r�w
e�9	�q��l�O(��M�䫫�7~~���D[Z�P�pU���nr��:�b��\�®l\�[m-�b��^��Bp"��;A����qH,�onө��PՍk��?r�'.>Ù��l�{�J��R�N�zrۿl���m�O�b�;�sƼ�Ρ�������rY8�Y4Ug��9���5��}r��7��m����%|�\��r���;!�T�-n��:�:��om�k.#-m<�
�¢�V�U�O��5&x�G�TD:{!'{���6�y�+�R�
,�K몬�r��e��ۂ��cG5j�Z�z}��v�r���q@W-87��t9���Y1���P��3�s��ԚJ��?]�𻌝�֎YMɝ�{�9��N��hPo�Z��:�>��p;	TUu�8����J{J�Gn�\$�ha�L�I�FH���$T$�*�:��ݱKGfw��6����N!5$%;U2�N�k7iN�x�\5�2j��#�\<����-�	�N;���>����-�b�sԇ����FQ��_
}5<�w&�����YȚPTZ»�eѵ����k0�!�T�U�1P;��ت�g��>�Y��m���z�ꅝ�'Z�����Ꚉ昚Mƻ�G#]q��[�1a�wmbh+W�f�c�涯5�饩:�X��6���-ߟ������c��&Z2��;�:�%�T����sڽ�w����[*�y���'-�ѕ�4�F֯p'^�qۡ�;ؕ�+�:���je�8�5�.�]n�"miL3;�_����f�3(��b4l����o�y���<'m�ie�5Y���[�[���1w�p7�i�ؕ=R~��h}�*��������*��]�^�ʤW�\B��j��wY
s{'-h����;\t�6+�p�\&�\�{q��=(�
A^��l
�/��(�6�Mep��E+}��hGM�u��q��:x8l�go�(�ޘ�K�->�W�Eu�@u���O�dM���#Wb�:�2��u���7C���JIF�l[2��[�������癪!VZ
�}$-�GU[m͹�Z���{�H��T2� �}q�*U�u�Q
�+�-�8n�8[I���ㆣU���f�&{r�`_�}��vRJ����٨-<h5��[]N�F�GJ�Fk<Xn��\�[ycu��S�L䘱�+�U����o��o`��f�s���J/�r��(�!O��wI`�Ko~�}�K��7�m�'��p�	2!��O-ڬg9���Z��l޹fa���|4Ϧ�2�W4iu�c��q�i%�R��X��s�|;��T?�#1����Ӂ���G��b��w�%��/�{7��>A�}S�0������vBu��QB�k��_R}�xF2*���e7�y�k��jg�8s_6�_VJ6�-j���������k��=�xj�=�or%�TD����nVw';+�ְ�$�)�0/.���_A���[u��xj���\���%�u�qRܽ��8�JR�&�h8���T|��*�)��,u��;EXkkav�`k��y:��r�S[k�5b���B�s(=D�s�����|�"ܶ��ک�%˾�w�v�n��^#Sb����v�ڨ7�4�נ�)�(U.ۚ*��Inϒ�(�f�V{�{�ld`��DJ��<��X۱��hj+zf]�.�T�uV��mk�)5�u��h�4�̒�پ�j��Av�R��[�¡�QP�s��V4�����Ҏ��M���:Nr�w��vy��
�#�&q��7�����`5a�v6]� z�I�B�.�9w`��c��98U�`.�:&agoT��H��;OǴ�讑̻���MkQ���:N���Y@�]��a;�Z��\>����d�Ru��s$'�j�Nu��K)b�������M`�@p�9�:�PP��]v�ݗ��]#�k�<U�W����)��ӧ�^[�D5cЇM�րI�bV�,��V5��UL�b
wP{�ՙ�GN*؆�Ƙ���W��󜇂�\���1�fʏo�ʒq���Z�V�5r��@�O0A�h�����R=��l��a^ܪ���;dn�ǚ�JLa,�*qu��n��A�w�,�+�˕�q�S��-�%�K0,IN�H���ojm`�qn�<��R���%�������D�>��'˦_(�!Hv	3�[�2ƭ��	��djWʇ#�c���R�B�}h������)���U��K&��[�\�w�S8D8�Pɑ�#��A1d�x���l��4^S��K���7}}e�h�T��f)#�.%���4��T�F��f]�ec��AE)�҂�Z��Z1m]e0�"���������k(��tK�@=��l�Eqzj=gQF�c�V�f���u$�}�j�Ɉ��:�i9g�[Q����7���j�[��)U��[>���{����L�`{��k5S#iT�"z
G'f��0�,���h;A�[O�z�A��v.�fϞ�չ���1����dP�e[�>��B�'�ι�K�q�-��\��;�o�>��9B�޻R�ڕ=���d�n&rZ}��br��N��ӼȪ��\eSV�����0�&m�JU�|��2�N��df��R�hhއ�;X�nI+�tۙ�<j������Z�ʙp2�y��r���,f���8�m<�A���Y�7��ݗ�(�X�LWN��=�T��k
�I�O@s"Z,���ۘ�.�ΰ� ��cnp� ��6��"Y�V��Joe�]���m�0�����W�r��d&�:ҥN�8�	��@��� �3&Y/c�[�����������|ˍ��ס�<��x��yA�� �j�qu�����f݄SP�S���p�x��v��{���cA	1�P]��wR:-�������k�O&���	��S�Z7�-�k�׃��1<�N-!&��br��Cw{���^�p����ZGF��*� �ZѠ�b
j���Rњ����B!�(*��bJb�!1mA�i�Mj��(�4i(�-	���MSF�)�j�cEbh
���Ѥ4���M4D�EQ1	��+H�ME:H�Q5@RRU�R�]!��[�Ѧ�Zh*��*�����J)�hh��hM�T6�4bP�&)Mh�h)-j
(Z(-�4���P�6Ƃ��(+cB��B��:CTҚ4�SACKTi4U4Ӡ5CUQ4�)M��4��P�N�iM3SSJ�U  h
� N­j���æ �q�c�ae-��f�������l�[r6�wr-0�¦�lU�JAM��܁Ae�T:��@G���햬����&V\&���{+29ٺ�C2�s1T��R'�fb��V�g8c\�-��r{�<���jg�^||B�֖�8��O
����������sw&�N�W�T>��&.��=�9���v�Y��ä6�R�4��(ޛ[����n��-�x���V���m�|����G�������\�U�U�l���yVԹ���R�KCw�ἥqqqs�d)�0�*�iV��m�މ|�Т���I���ΝH�\.���P��m=��̈́��k眶ͥP(t�Ϥ�1����)�\���bt�����&xh�2L���r�E�6�x�T9J�PS�w:f�K�����|���a�y�v'��[J�;ո��x�l9fa�fͩ�orS�z��_�����W=�if�P�J�|��T6���3��v$
Ö��T;>1�4bR�V��Vt%&�5d�n��a�{�ޏu�6^K�*�'���>����WR���Dz_$녠�!���.��� [���ΪG*�<��M$8txQ\W�"\�7m���U���X�Zy��וj���\���
�B_��n��	�gO���*����뚞]�{���2��4����M���o!�p-��J��g;���`S����Ô9�yk�9�Ws�j�n�"륾q)U�Ck�^�bk��k����Dr�-mDj���ʜZ�T�C=['5�w��hf��ٮ;���u��2�����{�v��/��g�ե��&b6R��H}���߈��*{�z|~��3U��=ʽ4=G2��;K�'��}e܂ɽЎ\���Q6��;TN[N���r��=Ƨ��Ӂ�7	��O���G�}4��	=T}�(��Aw�υ�)����\ظ��lOv:��k�ZOw�Ѥ�w���m���g��X��Y��=\�޹٧]��3{\ۚ�t�Ӫ?C����n���9(�<�j�.vu@Ẑ(V_v����G���lv-q�1V����떞�|of>�Ҁ���!���Ղ�q���>�F��R+��S�Z�G��o�uw��z���S���݅�� �2$%]k�0P���ə�����0�v�����!��[T��&�˹�( ���}��*%{��5���ؗ	���;�Zy8��z��s.H�F�-�f��x\�;�T���u
�Mjon���[O:�_
<��:�F���u'z��:N1Pn^��I��<k��ͨy�)JKs�e\]��(���zBq�^�Ǡ��h毂ޥ���}���O0+��2��yo+����,+տw/�x�E|5s�G:�o��Bw8����R98�P���jaf�ƻf~�B��Ou;4;�6�tm}s�w愙H�q�����v��}�[|��#q*�3�l�:��1k�z��:�6�1Z�^���m�ήBy(��G"c]�<��[['���w��oyª��Ks���[Q���	:�X�MCn�G<�~B��~Jm3y�T�6�.F����қ+2����yY6�s��\9�v4O*+c�f�r�~�����y�.p�|�]��%`���:��v�^2���vx��\�g�d��~����L�\$�Rު����ZM\��gq����j�ôqf�+���0���KY>�<�S饈�~�r��t3g(��� {&�4��L�Cx�j��� ��C�C#-Zw,�m�5��⮮�,!�6'�����fs��e�n�br9����~+'�j��KG�U_�ۇ���R�ZCY"ft�9
���W�N�%���5�}{�|B��U9a�{�oi����(Nq�o��k�(��6*9sb�Z{p��n+�ʢ�Y���V�b��⎭[��D�Y{D���zj'T5c]+����妟�gGm���e\���:��%< P�`�Q�.]�XT�R�-���,o�A�y*H�2��d<\�H�aٹb�f��
��e%��t�h��������]��/`�]��=��ž9])P���>
*LTIb��O�)n�2+\.��(q����mn7��r��!LG}�	h߆��m[Uv��vuZ���-*�;9m�SJýj��m��,�!u|%*��v����	O���w��9�zzr\�����Q��Ts��_3�&.3�H�w#�|��3�]Tu�	�d*��n�wn!X�m�ʖ�s��(w5����".�ۼn������|�Ō��K�_]�b���
�g<�L�`�@Q�s%�:�/����%YX�9���N�`w9d+�LMâ�MU@u��H:�h����n�vvz��	0���sWO�oy7�>��������7�A�n��]E�](�ܑH\���f��vjڅ��6�k�����V�G4���Am���r����*��x������Xa�/%\�i|��;�ķ�z�!��o}��j���U���:��9���~m������e�[�Ԗ�=�d�\�Mj_N ��P�e�+���Ww&�R�|���1���r�h�l(���:��ݷg*9̥ݾ�/R�J��窭�n[X=^��obLڮl\��O^o���^���Ve6V=�J�I�Z1�WU���j'T%p5Ҹ�د��{-���#��bc{���t,�@�ِ�|*;ʁ�u�y:Y�;��a�a~�=A�J�e��Qa�N�N`KOl��|(t�rf
��|�jRy
�t3*݊�5�"�k���J=~HA7�����F����j�8�13)�wgr���p��B�����F��W�P��{�J�=gwtc��%%��S�6�����r]X�"|��]��=)*`���DH&EhfT��4��2
��[��nr� ���{vxl�3��'���z��9h���C���A��ͨ��L�]y�(����c�mc�T�h����ծ3^3z�*�PS�w!ٷ�^��\��Q�K pq�������}��Z�`�x��9f�{;��VH{�]S�ϳ#E|[٨�\� ,U��RM&��)���7�q��z|}y�2��ǲ (�ek�˲�����|�R\棤A�w��Y�^J��!�9��}�X^�	]+Pg�\�n,>�oyem5q� d�\5��7+�.������k�s����;���}=�[�:��2��{�Sܮ[K�-�擭��N���M�Tk�z�l]!���%5u�8���k�9�쨞z755��[�r�����zhz�eOs3����<�!xO�
�<����6�~��e����iڙzʮ���no��<�PٻEJ՗h��&�$�kf��N�@�V�MԻ�$����8J�MEyo2���d�Y�h���9x�iMT�o!uyd(���O�Uj'�d��0L`a��s*�A&_`��>��K�M�F�����hs]�G�ku�a�����x�TYs�`갹TM�T	Lu��˙S�S.QU1��Ir�_
�}Ze,�V���ݽ��� �*�w�#iԝP�p�����x�X�ˁ�zgk[���]�n�o!��e�� s�5���{׭���޾U77��Ɩ�[��6�}-=��{�G��T
F{6V0���iQ�t��Ю˥J�Sx�>���i����P�ę�)�';K�V.@�����j��A�:{5�����6��8�{"keYv6�T�PɌ���%����f�P������w8X��^���Uf���B�6㥙��;䡊�����@YԷ�a�_B9bUS��r���z��8y�
�m�S�e����w}�'F������֚��)�V8�n篳����Bo��톅B�OG!�:��-	��,8�K���W�?��7�ʖ:�/�vmq���Ő,Gϭ�B�Iq�h�4�{]s*A)�t��fٛLZB;w��+�s(8ӫ�r���j5���n��ήh����̀�ݹ�l
eU���Gw^,�4��R�H^V�E6���'pܘ�g�imB�7�5�P��h\k�:9�M�\]d�K*y�C��a���q8��j��V�!'SK)���yCU��{Kƶ�U9^3��Zʲ�%�䶧����{{6���k�==�[�bl�������3��. ꖲ�Τ����o9Z�N�u��E�{!
W6���U]��9�V��fw���3(���Q78Gxt����sαգj^X�ޗ=�ⷹ_�g��u�&���fݜ��3+�A�{hSz����:���}h���]qulWܹ�r�ۅ]�j�b��TR�T���Ncӵ7�'syX��/�J��p���J�ط�|�|_<�{��[�@[G�M�&��4��RWL΢vx�����R�|[���ㅮ(�۬'aVX*C�y{v��m
c�?��TN�K�u�_�s���i502�o�h�&�VS��kO��t(&�����3X�z2��A�īP-{x�.C���Y'psV�+��o_���R�4�ЎJ�7�+V1B�oseN�5+��q�+f�B,�r(�3�V��4!�����X�{�Ok�)���W�6�t��+sK}�t��Yө�����@��)WO|�(�	1CRW�8�hE
=�����RZͺ�o�����'��r���}�	h3N1�!�^=wgm��km��ovtAM+��k��l��v����v%\�0\q����S�����鯧u����1����\2�;�q3�*�r��/4�;r��s[�e<�4��r{\�E�훎�� ��o�j9&���7�de���.�a�X�N�U���C�G�ҟ=��^?{ݹ��7)s�Cƕ��w#��&�k���Q�ћ�H.~m���=N��{>9��î����L~���솗�����<���z*��k��uyU�֫�wU8Iu�p�����L��I�5�>���^Ls�z��AL���ڎ��=�g:Sw{n>�;Q%1��2�|�y��/W'7�{1n�EіȾ�]���� ����efvf-��ga�*�U� EH���>}n,�q�5��Z�%� �N�^�N=�UeٰT�=]�}t>�a1k7�t�Mj�2�7݊�i���EW҈��e��%�hS����w��	��T���wۏFGo��t6N(00��Ԉ��r��`-us����b��I�U͋�iꞼy��n�ʊ��B�lRa��WeTE!�E܃���u'T%�t���د��z��v9a�H���=�Џ����to��2z������{*u@KT���*szl>w�3�9�V�ކ��|Zy�oz�:~�@l�Wϕ���g�Dvg<kȃk�5G3�n��.on5�Z�,眶ͥP(w|�>*1V�
���+I{�;���`�*~�z�}O�7���k�\f��r�r�

�M
�YC�Þz�[��M�0!�Cy��}�b}����[�7�)�;346E3R7bK4��۠�84�#&#>ލ��us�|��T$Ҹe�{��;/��%fc5����WZ3�,�D�}A+\��j��r�vaK;k�i�^�p�X}�{/V��q�Ѹ�T�����ua[iқ�g�W��8^��ct��]�����@�nÆ�����u�tsk-�[v�+ʏ:��s��m��5�j-w|�XQ�^ZԜ��^u��7��V=a[�;t���;I̹��)�;k��^����2��[�GiJJ�;"��T��ْ`��9�ѻ��[qGV���yMp�̺9sHV���b�����z�oS�(�HF�b��
�Y�_j���p�b�t&6�" �٘c'%�ǝO�-����i�(
]�5M�/��[���f�a�I� �!��J�9!��v��1���)�N�w.�	�x(qG�7�X�A���ݔ�0oMe��⒮k�)�x'�i�ӗ������.&)�r�Ia<y�� Wh�n�.�Đ{ʴ�iS�\�w��9G}�Oo鼘+و���v��z�6X�xcM�{2��MrGn�d:��=�t�5c ��IݝW/�,���NxH�ș'gIMj�},��T��8�ؔ�T�Z�_s�3G.1��d���𻹅,��RA_Fk���Ďv�L��{�`�ӱ\@��x�C��S���XV2X�TH)K�Wh���).͊�7i�SR�98��fe��ۧ�m6.G ��b�eb�X_0��c��\'2�;;|ȡ��1B�(��=ɍ	|�B�+'IB$u���WǫT#v���F��Y(��'RJ��DW;V3�04n���Vv�<�^�H��@%�.�c/oW[\91�!�3�
���+�N��tL�r��'¹)�4��oko�ݖD��c�D>rD1�_�]��\���s����Ե���o�ݑ�����N�-V�`�iǶ8W\`�?���~/�eE�#"9�e�e{�aQ�j����IU��3a�r�7cz����K~����QTn�(�L=���7l龳E�U��}�`·l�Qn�A�%t8ʸ�g^e��o��5t��պ��k��u�/LH�+NeXoz��^K�)8%���hy}SH�r�f'�8M�R��3k�~@1�ǀ�Q�����-���鄅9Z^���:V�_W*4@ʘ=#n��:��x�wwٱ����3��m��8!O�C�ы(N��sk2��]��Y2D��&XD���܏�Mvk�q;ǜsH��,�C��̼[���Dipa�	�!�J�(9;�$`�P�EG�C��]��N	�.�]3��?,U��c�[5��ԗ1}��8����J"Xx�ŗ�٣��*`��\x��o-0&��M&��{`�T��Ǝ֋���v��T���{I78�S�5��C\o�i`�5iv���ّ�hot�Q��MW�^*ͼXVQih�148�u!l��Nd�j���͵���]D�"�e�͕�v��:�l��"�.C�}�qC�e��U�u�3l͔�0yOv��h��8q��I5��߫ewa;}B�jQr6��;u��]`fm;Є�D]@ik������߽o�n�}��TR)�4R:t)ER� R�@PRPP�@�Hi4�it�kA��"h������!��J	AV�4R�-!N�#�44km��A��Ef��4�F����Dذ�[g�:4��H� ք��T�tR�R�T����ֈ���Ũ���)"�(t��a5@�ڂ�@��-�ց��t�4��Ѡh
ZM�*��y��}���	�c^�������[kU�3�ز�ɷ�5�Z���:zp؀������U�VΩ�TzC@��o%�e.��DBթ�3б1-�����5���y�[���-By9�[4�V�VyoS�׫���N��8fځ�ܭxn�X��FOT���vy<I+*��B��a㨉y��F�Y4�9{p��4�4=G0�x�)�G�k��V�%L���f�f:�m�IX2�TLe��L�g!�j�`nѐ��؝�e��i�ۍOCo��=��Q[���eP����р��ȓF�z���rk1/7n9�������U �*���m:��#�0�5�X+*�]#�Cx8o�܇m���n�,��o]��=�U�ڜ�m����<^��Q�r���KCc��y&��t���� 6U���0�tJ�\�%���À�V�vU|�T֦��j�c���{qڥ!��6�z��kc��T8;w	��H}�:{4Zy��ע����x)Vl�
��q<A&�Y�0�Ҏw/k��%�;d�=�t��w
���j�L��x��=\벒������]+KJ���C;���c����Ɯٻ�\i(gVd����끃:� û:Jw�`�骷���B��XR�]��y��{"��u�z�7�C�;��T�Z4sW�oT-}!���28+��ˇ"ڙ�����96�E<g)�2�S�S�-���0,��t��˽q|hS�q�S�"��[�0So!�8�]_@��h%>��$������{Ź�Mp���N��ʎ|�7��vôn&!1�l�ύ�����MD��,�髮{;�;��:o�j9�&�M��W�U��t~Xֽ�8z�?;wԦ�`��Pۓݙq8��j��V�s<���OA#c8��q�:�.�SńN��|�ZSk<����'�Qz�j���Dz��o�/=ѻ��Y+����%Y�c�C&󡘪&�AX/�;}$��
�ݼhiW܇S���g�ϡ��Ԫ{�߹�ʂ�G�9�=P��*��i+�x�'8s��-4�!L�c"^��Mo\u⪞����v�=:�7/_07��(�k���iq�ޭ�������a��]��9Hh�,�m��
��L0��\%QEg�����\��D3�zb��r������ڹ�0�עњ֜�Yz,�&�b[�c��L�#���T�W�.=3���'U�Vð����C��εb�*ٜ�]��+/^u{�^8���-h?���
�6�W�{g*��
����L��f
��9��*k��	F�]n�M>�|�9�f/9]�ú�=P���m6g����P;�b�q����e������!S�X��C�����g�l+v���7�;�(�N�\�������z�Z�y�u�����c����zs�9P�(����*�&#RSvjҫX��y��*&m¤��}��v�r�ڇ��9FQ
{��,�O�ލ�MCy��-�,;<��y�uB��)����
���r�E�n��tfk8�g�!��01��|�@M�>9\���_3�+g#fj�\v�<�̵d�.
Ηe��yF՗�M��߾�N�|���ꚎI��긞����I��<�qҪ��T=vG1�
ڈ��2�9�^j���ﺇ`��7�@�]�6��{�D�Q؞w�-,�h�Ֆ�Eruʘ�yβ�3<���%N��+M��k�����ա�l�;hk�.��s6��,��JYҁ&��p!1����_	�2�(vU�%�=�wx#�Ë�L���j䣝/ U��u��䧝�$2{%�o8��k�G*���s?[_Z3s�n.~�ն�c��
	c����y�:�nu���j����V�BeY�Ip��������H��gIl���e>S/-'�C�=Qy1���j��X�-�/X���pt�pg=U~^�È_1y�'-�jg���N�n6�^'�̱��d����� zl�������$�}��s=:�q��{vo&�H���[���ĥ�S_Ee����O�����Ӫ�=�R	��k.�̵y2�^Q�H�Y��z�ѐ�z��	�;^˓�,�sY�p�
�vy
�V���o7����i�މ|�Т��Ѵv.3k�*P���w���X�=�!]J�N��\5��-y�;�iD���L&�̥g�����kL8��Lso��;t�Y}n�?t~������w�~1^��J?5�S�8ƞH%f�2xSG����!gw(ը����ڮ.M��M�ŕs�t��aZ�@���:��wS����]�^�`��u𮡸5t�]OR����5~�z��+���l\��oWu��ښ�0ݹ|����D>������oDg>��YՉ��҇Y��otD��Ȭw�	=t�ts�b��]�R4�f�W=�k���I�5kX/�eM��:��(���	��*y��Y�	g�A+\�]��o&��Y�5��=g%��q,�����o����	R&~�_x�89��|y��8�-��u:~+�umj��X�6�V&%����6/�~�:�N��*�bp���r�TNv��յ���N��8f���m|�V�5,�VU7�;e�����m)�����m>�ڷ|���\sO��u!Gdf�ˋ+�|�z��
����Z\���я�[O�L�d�1Ȝ�ϧ2�Ȫ/`n��.��;̙�=u�l�T=��V��6P���IVY��Q�ޮ�m�=U{D���3�w8j�yE����U9��5���)�{�;FЇV�ě�][N�Z�[�k��|{ˠ�z(J��nE��F�^B�lS3iRޖrVY�Y�tٖ/�=s^���:���70�!D[�/���-g�w$u��V�p��z�1�ŎنUjd�+��t4{9M������u�ڕw�&5w7U=	1�F�G>o]7�v���9���<�bs�����o�z��'6Nˉ��B�J��+�p�Zm�Ĵ�V�Gm�Ʌ�&�Û�}#yV2��v�+���C��_N�.��*g57��5���6��<�w1Z7E�;�!pVT��Cg��Iw
�gw5!�y,���5��j�h��h5ˤ+q��WJT()��}%A	h�<�d�K_I�9�" �/�A�ǥ/\=�rW�qර Ϯ?�7���f�[�o*��6z'3�k��sշ�+�J��o���v���]BR����j]K'�B���"^��������o�P���T��)b��Ud)���fY�zi��,+����v��-\������&�q���т�=kT�E;�e�����^�r_fO+�6m����V&|"\������2+϶w��)2�2;�ͭ��de��⫭ϳq����c��1�"�L묒Uɼ�fU�ͬ�wvnD����ٺV�����َ��W6�2��b-�"�]��^��.ﷄ�%�PIw:E������q�g�@@���u_s�2�t4�=���x��ϐ���̫<�қ�y!9��<��^�l� ��9���ķ�R8S��k�q���؆E�i�	X2V[�O/`�������4�Ml�fyY����]Gk�^O4n��̢�~�F�}��������x9+G_�O�|ӿ��62#<��95�>!o�֓+���X���C�Ɂ�'�P�-F��69�aKOT��¾�sW�P�vΌj��q�x�9�'gE�\��d���	_�]+ب����}%Va��ݹ��]������7��]Sd� �:x������[��h�WZi�����b֔v�&�ٽ��P�@pQ�򨝔�+��R���jع�tOBJ�L�|�����X�M��_
=�邠��&&X��q�2�]�Gvg��j_OAo��;}��q���r�_��uah��k5�d��k��K�S7��(`ۣ���[g祥���\���J�S���)D�c��"�݅5�*�I�^a��~�3:��+j�֚�W�ȃ�㽨$�Y㏷4��Ԏ��9��w��ZՂ�)��F�p���u:!\Z���U�9:�՛d���8���z�;���8�1y?T��h���z2U-!;�������ro�|����شL�V����y1S���N�-�ے��D���N����ov�8+�e\c�Ç�!Y���1�Q�'dLr ���
�˜�y�yc�E}���yMd�b�eXJ�+�ؕMC�i��ʭxG1����ꗘyl�)��W;�����I�{�okr�������[��\�j�u�O��7{yʷ�J�;@r>��תz��o�<ퟩ>��Iڙyp��kQ����f�i��n��~��Dɛ��[��~uJ+��[�'-�3͌�^����4kb�h���r6���+8]����D��
h��3�
����i�۝�c�O)m�i���L�/(��_���V�����:�݊�Ƈ��b��U��ۦ��t\�;�^f�q5o��Jvo����]eu�K�7̯|�%v�+�0�E݀2�x�z�ƥ�ƴ��ʛ�����g7�U�jJ �� �'��C�8���[Ag\��i�S�j��H/h3Ҹ�0�v��m�e+�C����lY�Kz�8��kr�}r��֪2�]��bv��'ӄ'������yڣp�ꥡ��p�^6��%�3@��^�ʩ�o>J] �'xz+[�>�Z-*2�����n\Τ�놶�z���ݷ�6J�4�$�fz_+ϪYo3qy�����t�j�����ٮ3^3v�\�W���Mq��U�Ca��LPɌ���-���b}���z�EYBx^l��M��[�cgk�(CQ�V� �ڬ-����ͧK+z�����^J�+�b�[{��y�a���v��,����V���]�3z���=��tf����Z�TG>e7���;F�aR'�����e�J+a�K+�V��OK�'Z�Գ�s�pک�X����k�g]q�j{f_Xs3����s��IW�,;u�*"qk��Z�i$�bp�E�jʱJ�Ѻu�{b�*N�}�����M�\5�`��N��K�=���u�hEkּ��C�2��Y����ܦGmNlN4J�n՗2e�ƙmPongPI��.]1]�9�ZA�9U��]a�Ry�"ٽ�}��֣:G}�,���4iź����)��Ì����yVdڴ�~�%�d�6�S���w�^���];u�&4bo+�N�) ���_{Z^�˿gVet�7����/�F[N�^�.�F&�O��q1;���T��?Ojl�����-r�;~Ê
c��2�ܲwn����K��Eopa�\��Q�rs�|Ykz��qʫl���%#UDLۧ�	*_�+�tk�х�_s�����]ueؤì��_�9����6�T��DuJ��u�u]+�د��x�z�Z{q���ݷ
�B�';4�6�&vI��U���|:��.��R�u7��k1����s�[$%/nٽ���⠎���HjVH\��D���s*Ȫ���j�\�9�څ�r��_
�}�A	h��_|���0���7S躭�ɝ��;��܄�EC�r��?"|�@`�KC��5�ڲ�!bͷ3}]��٘F���\�^�&��*�v,v���	�|�֠@�q؏Q���;�V�����|U%�B�g�]�WaJi�ݰ��wz2_<�k�ф��ڣ kdĆI�t�c�ۓn���$�CJݖ�z��2Q��q�3g"����
�&�r����F�K���of�Q�V�S�������.7�p�����x��0���.Z��3�h�Պ5��t㤎��u�[�rF�CVvCy��'!zj�zn��|�Mw2!��J��F� 7U�Ӻ�v��jmM����U!��K��c4�$Ѭ��O{mnL$t
�O\7b���}����xpss�f�l�Ո��s�H,J�FtZY�)�v[�D7e�蔬�E��d����P�;���R9B��S��N����O����9y���;�Me�Zw�>����9�WbS�V�Z�(e�:q�2�h���ҷ�#��9��4�ɸ����62�8��b���|�W����1MV��҃	�y�7f9O#�:z�%��^NU�h(��o���>���ә��R����WuG$�
쿜�[�m̛W-�=7r��O��*t��aZ0�k@�����<_t�m�k�;
h�]-#�*m��oiMP��sis�Ë{�.{�N++4V�}�[gBYQom� PI��.�ᱰ��=xc6խ<�^��L����̀��|��a*�*{ �+�>�s��#7�l+�m�ɱ�gg'Z�D�%i�����]2�<{Kyꍩ�v�wo%���|�]sH0�F��)k"��V;�7�Lvvs�8�me�%���ؓ),�E;���ƚW}�I;�Ց#/9D�-�x����j}�u5��-�{st)�ީv󴤥+�p���/T���B�;l昺Cf' I��R���@�;s���݁Ǡ����@��}�4�w���ܦ����>�{����^�q�[����X6�Te-&K���XW3E�v��W�G*��Xs�U��כd�U����W<�Se�V�H�gc���u���x6�v����GDӊ��k�vh�̔�U���҇���e�׮P�eJNޞ���x�A=�q�jY�I^Y���D�n����+/4��m)�p4����ۊveb�}�g(���g#�]��8Se�u9v�d�8U���y���jӽ�7n��Էh�� ��
�O2%�yI|w�F���pTjw���ݾ�4�ބU�����P%��[��.ehʚ�C�c�S+���_H��1J�*�UrH
�[%t��̝Z��vNU|D����B�;��.6��[[���[0:��t3L�0�X&Kܙ�; 9+4�_V�ZB��� �ƒ��i:;M;ȼ��P(���4���]��T/�D��P�*���}#K#�*Iˣ84ˡ+���5�������:���s2���#�*��>��#E1i����ch�h�'F؉4h��5����SK�4cKZ6)Ѥ)!IT�ht��R[U�"*C�ѣl�t�i�d�	A�IAI�HRS���(t���hХ%·.��4��)4j�ұk[d� kJb-�����ѪB���V�+Z4�������h])��F�JPi���RkM���RB�T;`�E&��h����E���4R�Ѫ*�)�h�t��h����lL!����;����Oo��[��G<�=�lk"��8SZ��D���O&�H������]�Ĩr��Y;)B��b���x��I�pky�y��p锈]_	H��/"�i��]M	kpqt�N�����=�Ϝ�o���p��¤ۣmO���nΙ�W�\�CnOk���;��s���昞�7�+��f�:�.l3�{5�0�ϓ��f=���#����|�f�'3����9p�\�-�<���.#_E��yn�����̫<��)�䶫'?ERy���*NU���Y��g����h��\��d�/��z��Z�M��]��Hq�|6�$�	�j��|s8c\�}{\��9�g��=4=��Op�=ih񘊽�E��չ޵7w���;_Ilu���>S<�ȗ��5�}{n�P�d]@ܵ}O�ВӔ+��z�c��[rT5��9�`��N�O�d�+���1�5�;75G�R�]����.ruBW](��}n�J���W�tjԴ ^]{�ឋ)�Έ�y�m��U�D�`�]n�����J��U�ul�Ǖ�}���Z�:��3��1&���v1f��b@�U����,K9A��K�7�ʣ�L�=7I�{V�*�Y����&Ԝ-� b��]��j�=+D�c���tdL_V�:����;؎�Xƿ�����mArb���c�ޭ���8[M��oz$u�����TN�JZ������ͷ{�����IMAM���kn���^�)J$w|����� �DU.��s����J<j��Y�_Hou��܄�5�7�Q�D)pfQ}��,VGfIp�O��,�/ᩬ���ov�M+��0T6��J�و]�)u�ԍ�piqFNN�|4˦��=������5p���f|a�{I��x�򮢂zr6x������P6�sSk���{�|'(�>�ez�+	�S/޴��_Wu�7	��!�ì��2���=pF��6b�����ZՊ�U4�Ö�c�r�^1�tZ��e�g4	<���v��A6��b�����)���r���N���g���:�y�vf���S�]Ӄ��snX�t��&��q��}L�	D�y ��7V�Ou�u2��`�T�3����ޔ����X5�E.�6��,9נ�D�5�`	I���<�kKl���sw�t���m��䡹*N��v����[�n���|��UF���P�BŒ�M���sS��n��I�4�N�_<]0�U���	j�k� J_�����h�	�2��Q9o�'�
%��ӪrxY�ix͛Z�!ml�Zqn�W��`Up*������Wճ�ǢmOՍiW9�,Y�	����=#>ؙ���,����8�X|�ي'T$of����� U4%4mYC�ZԷ"�}p�\َ�9(ȃ�A�ZtT�������=)w�齸�g�_��n�Ɩ�7v�ҹc���@�܀�9wDM�+X�*<�
fu�R�ϕ�u�MjOu�X����ٴ��wM�,�K����&�0�@�^��#����+������/���Z�g��6�*�bUĪb���z���+س)���4;���f|�F'�J�F�u��J�j��D��K�g9?����v��3�!O��S@�7����}�q���	g؎������TT��n�p{��x���P��`�a��eY���/K/ZU�ׂDI�xw��[ͭ)"|�U�y����ܓ�9�Z����ݷN��WM'չ.ʣR��l��(���x%)��^!ţ/���d�̝Ԝ(H���u.��3��e�w���L�B,�|
Q��sNj9e:�.a�TVcZrֺ:��rp��\�&�;�7���R'��	�s��ٲ�p�}b�`=f�(�<d_t����o<Z�6�MB���6�\�z9�}�Z��0�O�z��	��E?���j�'�*q뫌մ��$�:18f�ځ�W��Ʀ�"\$䧋�S�����R\��%�9�4�{h�>3��w/�.ve�zP�%x�G�fyi����nmR9���u��	�K��:������;�,�݊o&��[7�d�ip�5u�w�3>��=�v�D=��ExWbI^n�ڟ.��r�W��z^���f��f���^����m71xM]1� �_��]�v���k�j'T5p5����c�o��cf�f|Y
Qoɭ�[|���F@�sg�]mJ���R�J�Kb�7}�m��Oyd�\���ڣ�a�;//����n�h2VP�m�z���H5��䬵y��L�:�U��"Mdgi�TBO��^سM﹎=�?�ʸ�t]s�Q��C�.�ZP��k��J�ŉ���BK��^�󈥝�Ya5j��z��(�Exe3�
}�/u쩽[�3<�6�����k�M��|�w�s��1\EL9P�;v̷[
������U���0:J����ݭPu��(�b�����Jr9{ս�ik��ͯ�qʅ)T

{���P~	h���g����)����.Tj�v%5�O���jy��3��D)#�d�sH´��e>���������Ψ[�)&����@y��q�����IX�Um1�˻��	G��`��槟n�N�{�9�M�v���A*��:m��,�6���@۟��s_].��Y˘t�T�����P�Ӊ�s{��+�E'Uc�/'����>?b�=)�ߟi�-�7��=��9I�ǡl�K��p�79ܨׄLk?[P3:�^eD���Ϝ�$���7�(8��y���[r�ָs׌��yxe�ٞګK��s����x�̰����֞�nPf�@�t�ZJ],�F8S��E�GkE�:�O@���y�Y����x4f��w"��/���/ͧ�g�� 2�1e�Z���mJ�xǛ�b���.���e [z�,��N&�����lS�)T�'8d�j��B�ї��׵���ƱoB�;��hҎ��V(@�+3��]xty�q��ˀ����D�b��Q|�D�AĽ\�K%ȹ2	l�Y�, �EZZ4_oVҭ�*��&;�>l_���OS����S͛G�����hţ�>;8��Nk��	X�J�cbN���J�[!V�I��Nb��Iu�K���q(���k�����I��X�떫�ι�5+{\aO/�P�^5�����;�������,�������&{:����i�A�OBڋ}��*:~�M'{yjW#ع[>��u�;��s�5x§�_�������3��Nd�p��j�Q���/H��������u�Gk�V븄�͝rgh%�u1ٳ�ȝ�]�y(�
��h?{5�����.�6�}ְM��E�4�ꍬƷfM
4��˅v�Lܕa_��`^�Y4uj��a�m������gZEc�0�Ì��7��vz��n�N\���y�������ں���b[����"�8���"y;�l��[%NB��C�.ubn�^��O*��U�X��\���'G���3r�Ͱ�X�ڡQ�/aFF;盡�k����}�J��ɀy����[��a��������j�u:��Kk�v�靎�����xD�i�]�jk�ҁ+�܁α�4�S�Rʈ��w�+g\G']��*�d�WU���U(��j��u�5y�\
�yS�+��sS_^��]�rq�c�;T���瑂�h�;�霓.�̣�`fOƖP�c.;TN[�je���6�tH�^�.��x���
Է�>��!ʾsiEdvSڃ�-���VƷs�o;k��4�q��g��z&~��!mo_��s�
Te:�T��T���O=t^�n��SГ�����jԷ>�m��:�[1��T����ɔ��fķsܳ\ZTu�zx�O(��ҽ-ոn�o�%�����`��_�{��az��-�t���TRt��Z��t�Ճ2i����'q:~��c�Y���ܻ�Q�/f�`E�o ��c	Μ�<�k���N��5�p�į��l��Ҫαk8M��5B����9������8O@���J���#y�mK}2V�U5��Ƹj��YP�-�$Oq�Ъ��t:��.��aYR�P܎Y����DIZ�l���r�_ܵ��wz�� �y�m���It�n1�����LoϤ�ih��\,��'�d%-1�u���N9a�^��{�Ի��x�Ӑ~�:c~����OKGۥl{�F{���_ofv)���_�0�jB~��DzgCd;Lm�M[*y"tIK�5qV=β�i>�X��6'W$v^
���l���\�=��ޖ����Y�-1���8˙�����y�S��^Y%��D�����4.+{��r����G������^~�F����me;��M焯P|X�J%�e��-F�F/�6*&�<�\gSm]�a�UB�����䉜��E�:JT��W����"��%P���'tº�n��:=��ǅ�^߀�ͯM��5�r��Y9��^���M���M	�;�.�����6n�9ZzvR����oԖe_%X��u�o[����)�漵E�\���o/��'�A�9���0f����+�v��[��B>oU�%WE�;@|v'�:���z�^�9�é�����L�����Cxr��.���ɒ���P�%룼emM�.q sKUMw|��k�H#ګ}�������ǂsvx73/ZX�ǟ/9Q��8&7Ӓr�R�ӷ2���á��8����rj{ݱ��U�6D�Ģ0���qq
g�d���Q��F�U�j0�8+��У����\�ޡ�=
o�*	AmJ�\���Յ���2Ò��GV�n��7�]�	�yR�9i��z;��>�4 ��(8K�2��8�ݮhu�r�n���?W�T���C2&b��\虸�25��qT���)���C�O
�ٟ'92�]�;yb/��zq~��M�Q�UuL�uj+!�=����l{�D�¨�(�<I�c�+��0p�����"��7/�K����\<�d�+ӊޜ�����HzW�T��uL;ɞ tԔ%>oϮ};AE�JY<Q���k����ꉤ�{��l�O3c<��P��R�Af�A����3��4��`���H<��:��1���0=�^g�Y��n�)�e��kp���Q��';�*e=�r$�g�Q>2'��:�)c��dm���~��}8�|�i�;�S�ɬr{L����H��N\��Q�4�:S���#f�<��MTV�.{���V�iM�34̊
�Wt��tz�Vn���W�] �v�ԣ�F�����q�Cn�N�M�cU�y�3�Vc�yl�Od:��}3�I���&�E�now�v]� ���z���E�LO�t���P���eɫ��Vj�i�Y�+��wTZ����ŔΑ��7�I�8��Q�O;��q;0tC��ڬ���ם�B�pӴv�n[�����T���v�{�^C��]���u~��4מM
ג��&O�X�"�{a9�>�{;��0�x���[�r��p�4��^�TV���|��u(h�g"ׁf���w3�ya�xB^7���SW^��W�
U>�t�ڥ��gZ��D:�����g�ބ�C_�6�~������o0w�����XG��l�<�:�rpT�,��.c�G�r�~�^�ec�F�^�b*�U���������i�ۙ�Љ��b��P��U��5k�R�_���~8i�] �4��=��ye�Y�R�i��&'�۩�tx���Q�3l��K�&�z@��]���=��z��{vs�y��ˆ��ĺ�cM-���	�Ĝ2���+f=�g�]X��}[Z��N�~�T��>��uTz����ƃ//�u��o����s���4O�xn	�6"�8�PR�'��R�Rc�s�6������eKI��Oy܁�d�]�;�*�v�2ܡ@jв� �4[�6��b(>-y\\�
̮�����oN����^Tz�7�4Đ�r��hTO�f�G-W��rv���Bh,ѤZ��r�ѽ�H�4M����]R,PL���+��$U�e�b%
|��P����!�u�=Տk3o���0<�0h$��c��=�++*�*�����{C+�{.��f��Xb�Z{���N�|J���-���4��� ��n���E�f0:�	�j��rhU����kX6�h�q!�Ht��j�Lz�l �(��;s��6G4�y�x�%aI[�q��e�h�
��$��!F���V܂ż�	PZ~�]���%��w�n�JE�\f#ռu��
�PW����w�|�qV�i��Leb�.��Q��-	8�"�z���$I��8����v��
�4�j8�;wR$�*���1ѕ��5|��Ő�e��NS_G�[�'n��JB�h˱8*K���j��iW%�j���z����㡤Qp)[��آ��,5�1	�Z�����S��bZ�ڽ��H�^�m��L�"�-wF�*�)z�T��(`�A1(��O����*�/r����qՊ�Uc����P�RQ[}%k��6���\\,pf��vqt��Au����K�y�N��P-���xP]t;c�!�eҾ��8>n�9 �Q�nZ�����0�O_*{�� �H�$ 셍���e����Tpx����/zG!����9�k݃;KR�`�,�ǲ���,����3,D��pg��pI�X��O�7I�x䕎q����_@�SNv5�ɽ-��8
I�#��5~�~[իR�H������IW�o[�u��6��4jq�b�@N�W�fwC�_C�ST��v�F8i`��CC�;�pn����i؎�O7NҸ��;jv�����wV�=�m	��e��0>t0�:�\��nd���o7��*pD( ������윶v�o������I��9k�^�z)eB�>fԾ"�.�/��6�V2���՘Xvb�_T����qL씞�����5T�Oz�=�{�/���up�W��U\6���q
�҆7���lJ����k�v��+���5�@[�]�Qp�$�@�t��F��c���m)��-�"���a�-m��W}n+9	R�	��������܃�p�Pd�x�@(Ճ�PXG�:ЋZ���e�W
�a��槣�	��}���A����]�d{��e���!)��`�V>��r1M�h|�wϢ��SQ��8^�ٺ��x�Z��1�cK�8n\��ؒm٨4 /�u[�4j&�{S�N�v��=�*�8����F,�Wg���M<�+�W�N����Q�gxU
���$CƀA�Rm���'AM�Z1��kKE1����4bt&�f�ւ�tQH�EV���j���h��s;mEtQ�I�Hj�Q�4��*��V ��&��h��H�֒�R[&ر�I�h�
(ъ�CCA�Z
"��EE:4�������T�"�"�̕TEHD6��� ѭ	������jX��hi)):�]QE�%;f�JM4�PTF�m�6��it�D��M�;	�R��#gT�M��V�*tf��ڊ�1�V��m�AMZ�V�TB�� 
�P�>�}����9�:����V��es+��Y�`���h��^*�Kg\�&�go4�w��_Y4��9�n���Tgd�t���rG�n)3�J�q�����߯�Q�ߴ������x�E�TeG*�� �>%ɨ[�7�563'mo��\0*�L50db�|.3�:�D;�!W>������_�i����w�M;���U�PP��f.������r[�"����s>
pu����%����Ƹ�b_�8�5\t��� ��]q7�0�����2Y�a���įWQ���h����=�#���]�N5o�ߐ�
����d�Dx�~���q5
e���!3_P�=�����W�ͫ̌3�+���n��c�SG~�t�\4��f�u��*�q8K�+YÝ�n���}z=Wܑ���>gl�ϥ������Ԟ��I�n@�q�*�F��������|=2UT��S�h��z%�jè��࿫__�wK�p���g���f�EzM�z`o�]�lL�陗�U�Z
}�Te}��فj6,����Q>��v�͞���<��qП�/Kt�fs������+:{�3τ�͈������&�N銛�i�4���|��sʼ�^����y�꯲`�q)�A��.�MZ�����w���ͪs�XQ���f2����UmtF	�uHeͺy0!5���#��'���:�]c�'�.�/	��p:��p�ë��rz�ޢ�͔���8��̨d gU�E���M���4�Ԛ�l/W"���i��Z&����vu��c�73��&����# {շ9��{iz �݉<��z�ͣr�����ޥ���7�K�b~�z�8�ܨ��C���}��#:�"�K��4s��
���s�e�߮=�֮:��v^�Ł�����!Nok�_�l����=���/�&c�z���ֺͮua�ir�E�vy�Χ��kϫ�{�!�uĚq�㌃E�v�=1h�{ō�U���n�U���p�G�����l����J�xf�f��-�;�qva���[X ��g��9�������~�*=�]j.e���(āN�k+��t���8\���.J<-���nx���^/v��F���⓳�p�:e<ۯC7�,���s�s�I�x��3y#�Q� ����D��p��JU�u(z��"VNG{-5����x�o���*:���s�:6^K��X5l�$��K�=��Fd�W�;Q�9[8�v�d8Y��5��迷ɳO|&2����̿���q��O$�W��/׳���ݽ!cx��n�_h���60��T���;�{�J���U0F��J�9�{)}�\�ɧ�7ݗ׹|\z�k�V�ؚ�7���Γ��t;i=�V���c���7qYz��[�s�nK�nr�O{3%ٵ/���}��9����L�(�����X̅m<5����Q�s��UI��ϝ5�p5���9��C.�ѧ�:E�QD�Y�r`Z�m��Oe`��^��c����|߮��ߘׂ�鹗�*/g<Ϣ9� ���h�q�%�`��s{b%�a�����k�e��jvs����OYT�^��.1���p�"|�P���y�6��kV���ӱ0�~��y�X��y?�}��>���sʼ��w�wި^s��Q�s��nM�R�ӷ2��^�{�+�Vﮖ�bSw^��K��pj}�x��e���@��KG��q�>U�k��d���G�L�����pi|2�>'E0��Q�.�T-���LTat���9�,\:M������]�n��`T�O+0��W���SAZxV�˓S�#�Gk�x\�E[�,c߽�#�in����|�5��D��ʂ�nRZr(�N�AQ�|_��N��4��%���X����	ǻ�.g��k���е���!�Q>�܍� �ަ=�DNL*�4t���N�*���ʥR��y�������2%�P�]^a�R�ٶ�u���C��8Ol���'j���b:���P�9����
�3�m�U�J�L�֏\
c�Ƥ#e��[��rC
(�:�t1�r�	ݷi�}�v�Ů��r��ӗ����>ۥ�d
����8��7�1׼�e��-��Aҩ*���_��/K��H�5=(eGL��h�� ��+֌�4�=�uyw��'�\2��q�7ƣ���j!7^�ճ�<͌v�mO<�<i�zd��{�S���kWS��(�H�������݀�Q|�1�O�a�y����	m�]��+<6a���L�7xߎ�?ZG1J-V��_#�2*+�w�o�K�*#:��E�yY�E¹\��b�f{��|����~�Q�+�:u���	W~�Y��_�ʸ�
�f�����?v�n�{��r��Y�fnz����&��`c���`�3����1�d��*"_V�ȭ�����2Yx5E�e�r�9[�\h�ڝ9�5���n�k�^ڱ}��O�T��;0����ͪ����<2���!)���ۋ��/Ok@9���`�B��֕�b�Y�v�.{ٸ�r8���.X���z��<r;���u��c��i���/�Uߦ���?Z�{��eO�Ze;^�2ϣ
;;q3�l�wS�t_�R����`-�<����l�9��_�NH�KnQF��e��J�,�	�,����17�ˆS���y$U	��7[��nr8:��o���T����e�j ���٣M�:�{���N��\�/�����]:���kZ9o7�՞ �g ����կ��ҝo=y��ѝs+��{_B�1Qu�Cv]��g�$��+lU^��,z&�Fͳn�a�NeDs�"�½��T��׀�[�~2*���M1�M�T����y	�� e�q�z�����z��`��?q���7�kơuRjw��Jr�3n'^	��^|�tbtG��J���=�ǖEz��윮�dmI��W�*a��A�Uɚ��1���w�ǳ�K�+�A���uQ�v}�^\}���+�},m¹��O�ˁ's]w8D�bj����{�
�@C���+��������:sBk{���Y�/I㞷���/:�nd��1�*�	@��
w�7 ��!�<e���}^�)}>���!{}m�w:���S���5��]뉿uW�%P@J��&K}$Y�^s��V�և�}�lVĩ�sd̕>#��C�ѷ�͹�&�:�����<Q��{x�+��g�G�è�9�S�%�׭�Q�j}��8{������|�g�������I��w���ڜ��ϐ��>f�v����%���Q����&6�5~�p��@�=> g�3X|�R���^�B�[�_禱T��h�
���L���y�7��g4@���B�4`��!)���N�^��J����Cy]}�
0^8o9Ass�]�u2,�-]�Z;W(,R#x��jr�cV8�p�ŻR�b�����	6�v��M)M�7BGF��i`ҋ�ާ�K���𚛟3�o|���������^dɨm��U�>�k5�Ì��k=�32��n4�A��P��+�pT����|n��y��f�EzM祃Χ	����{f�	��y�g�6}�Ī�dǔl�}�O����ަ=�Uc×��q9O�����R̹՚�n�_,p�4�M���ʳQ��̨*<��쉹zhӭs��������N�����m贺sJq�|�_���7���n���݃G��c����L�Lb6�Y77}ڕ��J������$c�^����{g�y����TgNI��.Y>L�6⸠�eo��J��6gr��~���x��g��:����^k̽ȧP����Fm��	�V�?wfO[��b���G�2�i�X6	��vg�����kR;L�2����g�/��,�D�R��5h]M�Y��V\Q�+V���(�¾ڟT���Y�v��\s��p��z�կ�L(�=�\�J��r����{|�a�f�.J5�>$���`�2ܭwP}z��(%�ړ�����w��v�g(%����V�y,���+P�ڊh�A��r��1]�A٠T��pt8/��bZ^p��V�ªS�(��ozt��(�M0<�E����	���9��.�9���u�$܊���Z�n%������;�/*� t�N�b6՝��J���և��{�o�=q�'K�0�\�P<��11�t�Լ�`���z��+ݽT�n�O���wr�������?N�%D{}R6�T���9��sG�F�����Χ��@��RvW-=>�|=)�o��"�!Q��s��p��-���pm�Pղ��Z%^� �d�73�ٱ�pj�����j�*T��{���5^��~�"|C4�~�3`UpZ㗵���{C�
�5�����,��u�=6%5�ȩ��i��O���#����f�t��|���X�W�����Z���ofI�|OT�}	�����ek�q�ަ9��ug2#5Fzƛ��_wH�ţ�;���K�ͿO�;^w��k�@�jd�`Z���,���9���/����V�#���<jojW�=���ṗ��9�ez�X:iڑ:�P��\NH6<�Ɏ.J�h����e��#ڰ6��Oq:s���{iW�uU��X�ǟ+�Φ�e�f��<�ʳ�������9qq�qܖZ��&�pѕ�J9e����q�{Œ��������,����/�2�7������C�6w��)Y՜�[~�����ֱ�l>��
 V֕��O{�yf�ZU��[5(կ_�i[�}��C�#����1���||��΀����w�N=���F[+2�&�!��d�����=]���̗�L0:ʼ�|kjz���WH|�㉁���G�������^g�Y����dΝ�Fn�^X���N~��{ma�P�>��^�Z|&�ܕ����4:�`���)�y�kE7�s�8�؜���鲲�H{���]�(ݖQ�~5U1q�J}9�̨��ۍ]�=����y�+�Z��B;�i~��t&�_ю@���p�h�@�|f<x��*:/�6��o
�T(ۍQ֞le龒��uTj:��MB}O���n{���ڦFs�a�6JD�58�9�����Ѻdv糈|��6]��47��^�:M׼C4ϰ�������W�G�:{3�����V�Ag�l���.}��lt�7~u�P���ٌ��z���}:���֞��^~ڎ�#g��W��g�⃪Ԏ��J�ub"�����ï����հ��w��jF(��=�9���,���'��F@�v�%Oh����1+�\����9����l'��'8�t���(��s�1�j����>�><�F ��.A��,��C�q�QR��JC����^P[s���+o����G��ծ��`��B��->�eC����Iȯ�B�
���KM�6�X�]�G�!��2�%9��mv��t��6���T���xB��U����V���Kb��Pu8^�j���U:�}�>�Xzb lu\o��Kn_3���=���yL7�d��� t�t���Z���)�*�19æ$ ����mO�?}^���W#���7�{p�>O�|q��>W���yt*#��W��쓌�(i}[Y�׭S�d�K�+���r�TG��Ǹ��j���k�c>��/�Wq+��D�r�!EG��u	P�_�N�FeY�i�qdK���b��ճ�_�o;_�q����{<���
�[���V�^t�j;�>7ؤ^?�oLL[�Xkǉ�:�O�b��_��@y��|�C�]uVV�@�^�wW���F���r�Oǲ!�!�n:֋�KDQ�_�
��%l�T�F��Ƣ%���o{�Vr��~�k��7DW�כ[��x?\K�4�ў۔2�)q'L��n=n��z��ܝΊ�����+d��&5��Q�\�7�e�����W�xvNWp��oz	5�PW\���S�I�� ��Q�3���L߯�b����R|_�t�z����{#Q�k�z�e��t��@�)�!J����X�w]�G�ԅz����ނ{7ڏ�x�����5�K[��B�d=+���3G5�����ɋd�W�(����P٘3�-�n���©�!�W]��ӆ�yw�Zjr���X�*��g���Z�\9UMDn9:���ub̜7�TXuL���1г!��s�b��[��o2M��@�������B�;��x�B���,�P�xϠ����{�PzW��:��և
�#��s���(�E�٫x�\5��O�:����g,� 7P'���=G>��h����e�.�����8�q��������\�ĻeXd�6�@����?rM/@#��$3�A�5�]�n(�sF��DS��[U�Ǔp��I��R���<���93JY<2�;�.��c=��#�"��T|��Չ���Q7>gh�o�i��{P��Qؼɓ_6�wr�W<�;^M��.��VF��ʦM�g'��������rV�����j���7�1���'.���]ꘘ���,��e�VQ�/L�,�_�j�ևu>Ӣ�):�{#z���u���O�}��]{�^R�rj�Ѽ�r��*�+fą뙳�Y;�az�,�Q7/MD��r-����L�᜜�9��ǀ��p�s.���7>g�!z�o��)d������C��xy��_�i̴�oT��Ϣ�[%��k�
[���zK��To�s���-���̊\K1�X1:FMJ�sw���\-i�y]P⢸���u��j0N��b�}�����H"�=��<m�wU���z�#]m�VXx@�m�|����w>�K
�IL�z{y[�k��a\���_-o*��&�®��t+c�HmX���T" ��y�]�����]bVH��p@E�1fh7N��`-l.
u��X?�guuÀѭ����V�i}�Ԁx8]�]������砭�m�Mn1�ժ�z����	ՠ�f'`iI�l� K�Q�N��>����9r,e�r�M��P�r��rC{LWY�"��q��F5�쇄�:�^����K+�0���C��}�X���`�/��ӊ�j��l�R��{5I��c�qY�:�{�{�J�Om�(��_�>4&>��Xܩ6�.ʜ��GT��
�o� |����^�n'�r�ˤFF�ЈÖŒ��ݵ�-�0�VB��]��_8��m�^Uc���a�nO��x� C���u��.T��ku�аl��'kF�c�퇵�2�R�D����Zt�1&]뿀��+�$�,�5�^R��k�L��i;Am��t�n�V�Ho�v�GѸɈ���@j�P��b�y;����F
���Z˷W���*n��O{"�(c2pYOX�Y0�L�,���EG���P�ъw�4�ܕ�k%��"x5��5�7a�g�3�wp=�Y���g�f�n�X��7�;z�]�x�WgRξ��k��]��e��QB��t���b�]�ݤ�����
���"�ɧ[{��iƨ�J_���Z�s�5C��+��՘��ŧV��Y)lu�־g��z�e2��Piu�J�����`E����wZ�Ǐh�ٸ/��EWZ�,�61�%ْRzX��:Y��;q�[���!p�RZ�i2����X]r�ս4s�*�2�p���TB��p�/0�u6��A�H5I�V�e̗�Ĥ[DE�dx�+���֪��s&"�$YѪ'W�;�d�����0��-)����\���7ٔ�AH��՚��2e���&���8�빲E�t ���!-�i=�՚�#;4�z T�R*�<�\6��ۖ�+)���Ӫ�]ܶm_*�\��v5�Ⱥy,*M��*g�y�l�ά�ݴ��7+]-U3p7��Е������3Mp�ϓ�,�����Փ+J��擛՗��
��p�w5p5¦�F�Ʒn��f�ⱘ�N<V�C&0��,O�2��[�t��t3�سp��3���:�f7vZ��EZ�sp\�5$ܓ�kz�t�R��Yw��9�S{-���ؽ�	]���v�3�M�^3�������p�rٳ��6�٠)4�����愇:os�l��݋�[|!����Y	���Ր��qjUM�M��k������.����-{�v�8�y�TH.���R�{�UpѪ.��Kz�&o��+���ykOA|�i/�&��ev�Fd9Sn�r׈Ӎ)}����⺗T�GT�w���8��#<�����	�KZ���`5m�6�U�4V��$S$E�(��"�4hb�*Ս4�%-1	$�UN�b
R��A�QLAIMTڵ�4UQZ�5h�1MMl
��j�ld�EDU4m�-jX��&�gM4ԴRU�Q�[� �Ѩ��(�b֡����PmFi"+mDLU����$L�DT���)�*kF64Q1Q��Z�1$lӨ�i�	��A��l�M�M��H�ALQZ�U$DVڨi�蚭���U���֪�]�>߯�W�t��/llD�&�|��Y$޻��̬Ȑ���\�eLC��X�M(�њh������^���HHM�vAS�[��<}̯�O��>�~k̽�wP��������6��L:*mwz�R^��8�F��*�%���-���iE}� ��sC�4��E��7���v�A�������˸D-^�7=_���l�j)���p
~<+j}R�B̩f�v��\G?_�~�P6R;��������c��Q���ǻ�;%GĕQX ��q��9���>���*M(��Q;��e�Ϻ�[{/��ʎ��m!:mӨw���" yW�a���\Nd�?(�S���}�;g3mL�C=l�1��s�B��M��.�~;�`�|��#o�LM9�� 77z*�=��i
y`��T��<��&1�
�o��Y7����`�m�_5l��'�z��FUj���h����v|j{H�FD�HU�R��Х��{����W�7��O�����O�ߋ������� Q�3#��L7�K��qX�q��T��5�#����������ٔ�c�{�I^�2\F��5����;(�'r���1��ތ��^�y�Lw3Y0fʉ�}3݉8T��YX����{���y��ƹ���Tf�l����wab�e����[�iŐrb�`iWfoóWb��wB3�-eɰ��{i�O`��.�%LB���)9�i�CU���l�s��#x�E��C����Ʋ�e.�R�OM�䶑����z����T<r��� �y�
����d�E��5xخ5�����O\�|����]�nW�+|�~3�+áz��s_�x����:j!ڑ1������c���3ކp�Ӝ�͕7w����$l��IҸ��~�/�&�k��:�;Q�X&#Z�l����ʆ7[9�`�nq�@��K�������� 6O��]b/Ϫ�L��Må�v�o�=�o���2O.�����?��v��o�Ñ/��KGJ��C� �x�`z�c�G����%l{�n��Z�α<�=,�Q��X�g\Ν���Ep�i�Q�2��N�=sC�.�'�*A�lr��[��z7����-�_����zc�Ix�Q�N�Q̃��+���T�?#K�Tr�In�R>�^�N�G��-��	���@���h�]�(��+LÁ�G�r��S���ml�J�y]>�)ǜ��=q�U�/f'W��N/H�Ͻ�C�~�R6�uL;�l�վ��5�;�c��s���R?����9�W��uc�u�QJ}�H��ZW͡�j:C��������Q6
j5h]	{F̷�U�m1+l`�aLL�zoj����˘�uL0p.�V 1�8�Se��ki"3T$�����;�<׃o/��M�թ�K��=�J]��At��</B�g���{�����sek4�N�1��';nu����i�c �)��h75s<28ߏ��R��m�����)*zu�^�"��|�l�F���
���KSpja�D���Rt�{C�\{����1�=�GA��W4�����=�tY����=q�3c��Ǘ��J<�-��99���j��'�I��,����jz5��¾o�R+ϥ��,~�5���1
Y=P��z����{�^��Mj���Jn|��ϙ������o��sTT<rM|�04���M
ג���d��ea��)�E�ֺ7L����\�4�Y߫e��;	K�y׷!?]��ޠ=Jr5��چ��{8�u5.�O�"�QE-4>�*�XP:|r|�6tz�+�m]>'�}�/��:�ǲM{Ldy�����U�>���3W���=����~?����NlL�~��·u9GEԪ�N��`V�G�����[�H�	)3�/�������W�43voL_�g
E����|�
�k�}R�0�2vF5��CsrT�e3��6����Θ7.y�����7ִL^ܬ5G�~:���l�5�|n��:~ƒ*����4���2�EWMȳi��2D5g��!��IÚ�l�|;���;θ��{��F�OB���qy!n:fj��/^L�ڙ��{A߬���vo(�εk�S�ۂ�5�J�hV;�/�-�n�]z��9f��k�:!j|�-�U'����@5��؇�Q
>�J���rǹ�^�<;>����mܲO�(����e��8��h���Ǵ�����x�oUG_�\�8�e�F:����},m����)�TXمu�Y�D��<�2M8�V	=0����6�{��]Jf�ӚQ�OMƴ�/I㗀�#%*ށ�-B�������l�*��$)^3��X_k��W�
Q>���ʼ��A�a;�)窎�ZBq8s�{�4��=���Ǫ��b�J	Q�1%���8���B��t9��=�o�rff�K2z��{���w�����t����a�����d����c�z����(�+��s��w��\=����F��,#C~t��%�U�Km`�B�I��P�.zYo����NM���_q���J��Ox��BW񿼘��M_��zP>�K c���P�y�Tḩ��,]�SZ{����
N�V%{g��r��7�]����6�fO��2jr�gc}�b���b�7<W��=��ɮ�EH��lNu+N��}~��O��yp�����ǽ��Ш=l���*`��v�b˓�j��}�dk}�B�N�����9�[_eok�7v_\o o�}���4����4�mZU�&^P�l�R����j &�Tf�)�h$4�d�3+�7��!�/N��MWU��A6oz��|�i���D2�kLH���j��:<��sv&wcۇȽ��}u�j4�*�F�O�Z����}�E�'\OdoS��gj\n�{s�p޺���Քv��O�=ޑޕ���!�IQqx��*<�,�Sr��r8m�< ����={�Nw�q��WS ev��.���ϙ�5"��n���n�⣬��jÚ��[k;����������>�+�m0D-o�!�^���z�}Ӟn�%�ó�$�ɑ�_������a��x0��Y4<���+fDm:�+O@|}�Luar��>e㩎�ת7x�qp��7�kH�UP*�'�*��C�_"N��0���&�,�.��4:�K�[��íj�!Уo����Bޜk��ٍ��W�|v��h��W ��¶��,���\zyH�~ �VKf��h�NP���<��x8�C�2����C�3�0��F��%T`@K� qmϻ!���.4����ol����hP�:��FD/uy��yQ���Bt�ΝC�%��D那�w��zf�f��˾�vq?᥌���7�9�a{�߯�˹~;�s�L���+�~	�䏖[�>NG�ӧ-�g�~Eך`7}]��Җq]�*� ]"Yڜ/>4�ԥ��yPPG �Q����p;$�w�[3D��4�����uӝf�w�%^��%t"L���RwN�lt7R�i��b�4hl˗Ï�4�k�:�636NB�@���zը� W>�>�&"wԁ�-bf�Q��_w:�6��-�����6�<��ܴ٧^���{�i�*�&츃+|h�"e�����4xv�R�o܅F�y������uz���Ħ Y$�_Zޙָ�z]���H_L�]�P�a�-�X���M�*|n>k�G����7�펎��
Ww�X�L8��td�4�k��1���O�'�L>��0Z��8��n
�LpG�����,{}�{�;Е�3��t-�z��� �}�x(Tk�@�d�"�탘c��n�Ğ58�{�����t?{�s���z��Q{YLy���48μu`�tP��eH��d�F]&"���z/��}Y�<x2K��a�O�L�����f�+��$���^�B��=n^��ͪE��vM�ԙ�ǒ�ե�yŬ��僪&�p��O�A��&�����3�Y6�g��ҋ}T���a�.�8�q���Yv�
�#�).���mK��A�X�5}���*���~�(Dz�"�֮;��X�VvT鸲��2�P3ŋ���ti�]j˵%��p��V��Ik�y�S=q��v�]�ew�O&�������j�A7���4��}�逸M�՜�7����O����u���#gv�Wv�hԩ�f�I��*W&��i���6�KmP{Z`�@ޕ��d.�#��3��9��9w0wP�h�V�mxm����E_C�3�l�K��U��ܯ�ĝ���ˆ��[���Y؞~X�u��}.�Go�-�p[7��ڈn�=6�h�I>7�ğ0.O�yP�W�Een�\��Y������~�Ϊ�˗��	�</�|�����G�T���Slٽ�y39QW�}�I�d�3��$��n����45���}�H�A����F�z�v,���3��\��L�
¿Uj@�u�Gr艉n��t�7C�F�*C�z�1��w�&oL �25��4o����a5��-i2�{W�2����
��Q)���g��%C���P;_�s�w�1+�b�~���j���f.O(^<NA1��{W���Ee�= bI��s�tmvz���烯����*!�UH�>�K�e01�q��&9� f<���Gi��Ĕ`�[���;'e��+���z'�=;Ex�-뇦�7�S�MI�� t�t���8�о�ԃM?\�W�r�X�����~�p{M��
�����#�K�YP��V�|��|�1���Uj�<TPlN�wH�3R܂��mJ�˭����i���{���I�؜��,�B�HOp�љ"$��dI��Ӈ��}��I-�n�Q7Ӫ���J'Bz}�~W�L�.R���w ��6K��R��MG$�)B���-�]l�B���)p��d�cɛ�>�䰬l�w�ᶮ����\�}{^�w�J��6�벦"J��B���O�]����Q=��Y��g�3�W����t1`�j��>���	ˮ��3�s���eq�ad��W����45��|
j����Zcmܬ>M�p_��{W�(�Z�l����g}��o:�������u̡q��L�s���T�f��Z&/nV�ĿW�GY��9:��չ㹫;���\g��]ɞr��޻�o�d^zW�=��c�"�hxvNW
��R79���B�y̓�.I4_��yC�)�؝L5��Q�v}�e��o��_K��s��'�`}<��Eؗ�4NN-���?(��jg�1�u)�-H��{�鸍h3�kż�s�0׋�y���6˰lj!Aʠ�B��7�[,f���ϫޤ%�{]G�<����ɬ��̍���~F�:~:ȳ����e|晇p.K5���DQ7�F��;�<,{�K�z��_���X�-V��y�p�X�Cs�MC�P�ӗ0������1�}>=ix�G� .�H����=M�L���6o�	�Э���E�Ou]�=C	mqk��Z���d�s���b��l��b��s;s	�c�TW��n.Bk�A�����G[�,l:�n��lf�L�qf��V=99N�Ke�R��)�`mh����{D�9����L��?���� 9��������W-ωvʰɦ���B�I��w�\���K�=�9������H����n)O��uC�~Bc|��I��R�=^ o���%w�9�lg��! ��&}>'ED�D#c"}բ�+)x���R��s�\{!��{+��B)x��}t�]��`f��ٞ�7ɓ��<T��c�zp;���D����z\5yp���~��$f��^�Αt�C�ǔa��q<�E���7YF�K¬�id��L5:T�N����a�}��[���ּ�*�1pܽ���#�vC�ؕ{X(T/eN�,n���9���\�̹ѯx����h���s˯�
���b��Z�������xr����Q�����~�ߦ�=�oє|R���Ν�*e���i��됾w+ޓ���NG��>������i�ظ�'��̧���G=-��U��'H�x�������yU0�ҙ�Ƴ��3n8�x8N��s�\���V�	��$�<=uA-Z�J��Gk�q��,o$�Z�:��l��|m¥��J���:bu%*�̸nur#�ۄ�}��rS*K��o j8w�T6F�-�Ǆ��H4-���xqҗ��gEV�7::#��U��2p�뫡ZdD�z�Φ~�"&�G��3\}n�E�Y�B�����2f�����;Gz�Ĥ�熗��ܶVEy�{��9��(� �`L�X��u㐳*Y����4��{�T�jT��K�Φ4oC\.�8�ꇷ[1��QCĕ�e�/L����>��\TU�������*�-S�=����d/uy��Tt�Ƕ��7�C��rY@@���O�ذ�,�X�7eۂ�>&�ě/0:�F��\M�����#��\8�����m��������s�7#�iUK\�>�HvB$\�����h�u��E�ߩ#�3�}�uh+Q] �s�����Ҧ}<]������35�$�n ��f�I��R*Z:7����Bc:<��I��d۪X��,��ot�,�%��f���\��= �^��K��8�i��O�1�sEA��n��7X�}�nx��j�_�o�d�sN��1���L�x�;?Q�ٌ���_�ޢqы�F߻GR�o�������U�ΪEv9UCi�v���A>���.�~'��^�7?/T
)r�˙���O��^�0��ze���^u��_�����fw��V��jDƻ�/>�<W��P�<-�����|DN�nWu[!p���{%��<}!6ν��S�.�-t��Xh��
�ؕ
Vb�r \W:	[���U��{���P�-�2�O��pf��(��=V�5���ܹ�hXޠI�RŴ�"�TC�NV%D':��P6�2KZ����h�Dr�f�:K��\�]��çgob�vʾ2� �{��Ŕ�}N���,=�,J����q�Qj���z���>1�B��g�!��e
јd6�lIWAʛ�J�ֹS��'�[��H�������H�D��W^1�e���}J�,+y��E���X8�����r��|l�B�M�%�(���j�)埦+Ռ[�^�ӖD�W4d��[�\s�R��FIn��:�3v��- ��q�e��Y�<��.m�vx�4"扮�э�歛t1�J���ĺ�1��Me�΄h�{�����7.Q����\�ܱn����N3�5Irݲ�]V�*���|h���ݝ��&p��ǚ���u�i��z�\�Z��F���#����]F�nT|.̂����;��JK��54�f�yOU���2����<�h��T�U�-���$�x#
`���T���ܢ�Cm�
�Yb�&!�[b�Ov�(mC����.��JE F��gw�]_)�.��gK#(LJI��t��R�2�������R�=��sk�GH!�y���DB,I���Y��>��x��k0����NY�+p�����蘭�ҭ�v��6�{�D�cj��}-����c���h�uus�t�-�������j���2�=b6-=��m@��
k�)L��M�c�2��)���T��Jb��;o�|�ВN�W��+
�[�eu��c׸����$�"�����9`:���S}˶�V9�t�;�D�lY��$&�]���}����7G�r�&QC#�6[��z�l�Y�Ya3F���;{|��������Npq s�/A7B�$�9��K5��K�{����L����^�V�U(xy��+E��sa"z��Ǐ2���j	L�
�F32��w1��N�V���Y�P���@�Fo�wQ^U�Ӷ;,lH��b$,gV�:n���i<q��,���. "�1�)�+_;u��^�]H�A�������`�"W����u�����Ra�E��/�v��Fx�����vmsj��d�}�}v�EJz�k:�d�����{f�J�q��N ��n��ײ��MB�^�1���"8�sj_fִ%e
T���=+]����NV,8fmS��`�ν�t3���W0����Jwr��V��ۙ�8��,���9a�����Y|��ص�%8^�J��3eu��Btx������G���oh1��RxMM8�G3���t�M��8����Ȃ�೩�v�kk���7n�m����u���1f�A�<֋8i�\���@����w�o����_����jJ�Y�"�����E���Z��d�6)�L���U0I11UkV�1Q��(*j�*h��Vڊ����E���Q�Z(���Mb ������b'E�T�D4�Qj�N�����cDQDPUQMV��bJ#ji�������-9&"��-�DD횪"j�������cTDMD�TM��T�h�f��щ	����"*�ְkU3kRQ���IkS�I�����mN�QFڤ������TV�h����i���`���l�P4�1)�1RQCUQD�QQ�(4��"�(��*�("�����0@UQ�T�1D��D�m�(� ���-��[i"5��SA4T�Q�%QLT��1l����C�ot�z󶹙a[5�z�H���3��o.ι8Uǂɶ9��T�Ӻ�Ku�ٙ
�ݎ��t�{�\gzg�n�'�d����h�5Z~!�l�=�����1}3/ZY�/9���}i��t��g3"���zQ�������Μ����ӶV������^%���V/+�gΩx���r�d�:�:{�D��閯=H羍�Ko���h��K��KG�S��A�q��Y�:�/��띘cc����~�}��Ń������v:�b���MO�,Z�x��3�!x(�`p��Q+�?f�g*��e�9��9`�Fz=^��^�Y^��AW�'�r�k�<Iُ��g���g =5��7��MQ�1;2�ϞeD�Ӻ����8M��� v�u�鿕��'Ɯ���vԛ��'�+�@Á�<�=u��z󪠳N��M'���ϑ|������o�����v���P��I� �;��`!�,һ�\gM��~��M׼o�ճ�5�5��� ��ɩ��'��q�t�W����xߠ�TD����끎/ŌP�7�!ƫ���!;��ܛ�yz-���3��ϚY��n�m|�YBc�=�_Q�P6HH���)����˘��"yvQ�Uc iە�v�����t�o,\�S�L���{Dq�ܩ����j!�(�1uA"����4�2�2�;��B��ɳ��ە�
9S�5���[���Vst�U�x�v��Тh.�L��)ʨ�p{w�S���VH�t��Xs�������Z�Q�5~a����L�%�*�^�t�r�:�Uߧ�m���e]j�׳��^�6��S��r�M�:c�����o�R*<�Y.`[�q��'��cɓ�~��)��u�jϡp�!Q�eEOzs�e/3�q�Q�ky�1q�Ԟƀ�_{��8���]�.�}�O\s��>�\Z�r~�飊Ǫ\��]���{˴�g^�,O�|rz��)�c�1�1x*2RQ���A�sܱ����K�䰮·qY^+������y֮=�`��DWt*�~ʼLT׳z#��2���{����g�>;:O�큳���:6*U~'fvxOr׫���کN�@��Yg�ϝ�SW�}�9��F�鉷r�׏�;τ�2��[9q4&��u�˾=l�Ͼ�Ty���}o�F|�z�W���C�Cx�</ng}e��G>���٫u��Lӎ��1�;�H�hށ��GX�����kq��~�u��ڹ�o�X���7Y���^�?E�n��x�=�J�í�.MDN��v�TuƗ/�4yc�o˝�B3`h�}뽛���%������.	:rq7v��t�!���t˘� Sȇe�����i��n�O�|�}$�\�kڰ�G�V"F�nPݝT��y [���W���C�t��m蛼/"�8d	�L�Tɹ���ɄҒ-�DCU��(I["����������ў��C� '�
|	=Q2��)��uMφ������W���s=�`�+H�@�q��\,cx����׍\>ȃ6˰lj!Aʠ�`)^3c���F���QY��i�דOd{���kv�bM�!��t���#O\G����aع,�( %G�DĖ�H��ϸ���6G*:����[��g�>�������xcnwIx��˘S�x�x�ܨ�`ڃIF����d�5�d���_o��k��,#C~t�>�"}�3���|۝����G�>��s���A'��fo������?J���-�����1Qɪ��ޤ�z� �
��C.�c���@.�]/��"�V-'C��x�*pTK��WYKǬ�)|y�j<��wtvn)ܝ�w�=��I���L�����v�\q�̚�L2�ac�>��i�:��/6^���,��.�^��U�^�����7ѫk��n���eQ�,�E�k~Z�O��ǀ���K�}��+'|�1�λ��/W�#!��/K����^��币�<g�ߝl�9x��t��6��S��1
͉�$��kܸ-d 8�SgR�ܸ£�eH���~Wfx��<4+�Tt{8>��X��N���黲���#h ��uI|�4�=�t	�b�3�3��c��u�aI:����x��p�Rmu�]%o,�Jn��aK����h;���
�����L��Vs�3�����7��LE��/g�hڭu(�=:/��]DϜf~=���pԤ�>�\ �gs�:O�G��7\��dMԥ��}~]aaxZ�zO��tt���m:�5:��4�����|���������n=gڏB;~ز��Y�z��v,�3��ѷ�$�����tu�;2Ҋ����v��ɚ�I�[�G��C��{��oP�zr=����:�j�9ƾG��4��`w��/��׈A_zjL��ʬ�v*�;�]M�t�O��R%�w:cEƸs�/�;P�T=�����ǋ$�`��X��h�W=3{�yԔ��2=��NF��>�z�P��7X<�>:�8�y>}��Q��=¼��@�Of��l)Y�2�C< V{�1�0w���+�������\M���Ϗ���?N�%{}R5 �BD��}C���#&N�}��h� �<���Y��_!1�߭�����7�WL��V�~��"ծ��O�>���@�S��C�%�f���&_�
��M�o	��ȱ��uӑ���=vu��]�J��C��uVUmH���fi�*t�:!)�bf5��ș�bK��]t�sʒ��!5��
�����3 �b��;�m�W| �${��0gM{t!���ьF�Q�[�`�Z���{|�,��)n��'Q[�0b��w]j��ӝ-��ev���Z�f�l�|f��U�!1��H&��}.{Ƅ㕦�S��a{�ײz��w�O���|��*�1��ѓ\Ӂ��1�\�MǏ�-Gm@N�d�~�(��9ٮή�g��jٹ^����M^l���7��H��r�� �X�ѯ%:�>��ۙ����|I��=^#�_z:��i�]z�M����ԯÆuexo���q��3>�u`鯝��XU�-3x*&z���{��<�q9 �l�Ɇ�?�+��7�\�}�^�9$�ڍ�*�j�Wƭ�!Nxo+1�LLkV�֦F�X9ZZQ>d����&1y�z����)E���;��W��<�&��x��f��>���Ӛl:Ky��	�PO�u�<0ӡ�*����ܯ9}9]�u����n|��O3�^�ݸ����Xj��Ep�Oeĕ���1�E�W'Y�����\K�>��hu�r�n���gz\�=���11�^5G�=˺�P�;�ҳQB��#���������S�8�*%���X���ף}�7m���խ�f�{�U	�Mѷ=��?��=�V�&���u��hQR���*d�$6������yLn��z��vgl/K���Ѫ���V�Y������g��U�a��e.3�^wӵ�5�eè@`�Gp�����Q�}��<�c \4qe���s��F�ލ���*������y`f�
$ィ`(��L:���=�3�|��D�����_-�������Y �NST���u�	l΍�h�� ~Dp�X5�w���r8������#�s(��>����LTة�X�߈}
���=�Y���ʏM35�� "�}DLKu����(u�S�W�]PO��=���k�7Ѵ��^m>8��%�0�a̲��rG��L7�^SB�9a")]�#�棹��0�O}Dgw���o�Yd�'��l
�n�iK'��^�*{#o�9��=8�w�]���zuңqY=��>~N����̍��d����Ƣ��wH��G������T��I� ���ۘ>Ֆs��M���ڎ�Q���jM}����遥ϧ�L�jedd'��U���P:Y>XW�T+㿵�u����g�5Jab~��/�Ex�s���ʉ�5�\�������ι��wR3��]F��������'�5]>'�DwK�?*��x9�t��[�-�Q����3��R�~UQ<��f�g�3���'�����(�N?Z=��lnp��U�lQޕ3uN�չ~s�]���^�U���7!�yw����TY��U��gE���5������s��͹��֊h�XıI����T���3D�%쩽�R<Z͕gg_ee=�gV���J����˱��1D���+�i��3��R�]��DQ����t��5|w��m��鉷r��,��a�e�����6{^,�MߪM�R��u.��ȁ���Z����k��g��u���*·�vT齆��qt��c9����y�1�h�T+��w&y��>�u�n������K���]x1�R�'
}S��Fw(�m�R}�יRܢN��E�%zc��.MN��}��Qץ�Ӿ#���a^Y�=fǏ>�3ʷ�/'��Hq���l�_)�$�L�&�C�n|�.����N5t�5�e���ͧ��|^��7Q��Q�eW�h�*�,	��x��:[,,�����}����O����$�R;����w�#OS�P���;b#�}zK�1�Xuy!
�vnc�X_R�=�����N�p�ֆ�M�p���i���t���Zi˘S�,��{h���g/�d��z����R�WKGݿ@u�,#E�~v��[��a�Q��'�n5N�"EC����=G'�K(=�i"�=�FQh�~/���&��n�H?*�d�n�q�*Z�w�|(9�[�7�x��JZ��	�l���Le KV��;ww��n/�az��3�V�]�����6ẑ��U9���{��C�x�ޠ���%<���j��0J79�f[\��͙G��-��.�ʼ����\K�(�}�s�b�U�`
~��*:�I�R��	~8Tਗբ����Y�^���q뜈�+�F��̚�����/|��&����C;v/��d��a�5%����V�����x�� �y�=�y�F$���/�z��_9�1��q-���v���5���Y�����ꁓ����l��f��2�U��	]<N����x<2�ݑ��Az_�Н[X(/\͜����:񩕒�	��֝B�t�;c�\��ꛗ��t�;���*7<��!�z��v�x��z�w��1�G�$J�':���i-qk	̣1�!����Zd��W|6���쑐�Shܹ�z��f���2p���z�~�?�G�תb��Q��[5��4d��P��S��>7u1�d�~�x�_'9��b�ץw��\6VDz��v{-
�:rN	�I�K��::�ve�� �8�*��\�]K��:��>�K�����q�6}Kꇠ֜���+Ƣ�v~+�P�a�v����s7W�=~�}�̞�iq�r��jD�9c�\9��q��a砫f:�#�?G�$�7^x\��z*sw��>��+��C.=��K��G.'.��H(F���y�+���C|V<xlϣ��5* �����;�qh^�hP��*�`�>4��c Yճ�bв��p�h�+w�(hX��@��}W׊�l-,��I�d���z�/z���H��gT�n]h���h��2��*:z���鿝:�!(��v+���WE��g���{0Tx"��72�^Ø�W���$���P}��{a��i5��4�%���̡���P�hS�Q�%M" �>�&[��KG���"��m��7RTcY�u�l៎d8ǞG��Xw��+���M[*~�h�����"e����M��WF���J:Fd|�,8����Ѩm?�f�/�f���U�!?x��0R�:���Y��9�6������לj�u:�M8��_w���UI���FO2�c���N�&cǉفj;D�.�����ɮ\��w��J�z+U{��oSm]�b��uR;W�m0�G��Z�P;�p�F]��*O{�2����N(yPa�TONa^/K��cdܰ��^���r�^:�t����fr\㻊)��v��~�B�o��h�Lr��w�+��7���J���w�H�̺څqWv|�l��>�֛ژ[�83Z�oK���*�C����qS+ģ�e�ߢ���I{�E���{�<�!9��,�f�R�ְ8�Dy^),���n�{}��H�u�oq�[�m.��[N˅׽�嬆%��:�+H�������mo���Y:.D��M*��;R��K/I����h\�r���u�Q^��}n6�� �U��6�p�|��:��-?�~�j�^9��{�u�o�>ɝ���;q2�P�௮�g�7Xy��ƍ�E��_{3�xαܙ��tc��k<�s��õq������vY>Ve����^�q��̻>�Աu���N�|��Q��C��sC�0�`���9c.9�g����5���m�,�e����
p�v�m���=�7D���h˯�����U�ľv��<�[��8M��� v�7\�+oE�F�Ѹ[�������}%G@_A~�嫇��0Yn��MD'����_-3c}��=��ޚ�q�0ZY�i����#:e�l���v$�!��<e��uc��~W9 \�,:j��tj�}g�9��Cr4��}r6��L�9�Y�"�'�Dķ\q~,fb� �ad�^_�ԭ~���zxm���1p^m>9,�[s6�(O${ʢ�l����h7C���(w=>U�AҔ��z|=�TF7�ǃ���,�K=C3z�aO�\5}pכ��$�V,�6�k���]F'�.��Ed��y�|�Y'2F�T�y��W�o��� �"��APE�"��APEr
�+��*���"��APE�A����+��W��*�� �"� �"�A���"��� �D�TW��T_�PE�EA�$W�
�+���e5� '� %�!�?���}����W�|��H��@)R��$	PP(������I
U��� ��U
�BP�R��"�D�P%P�J��PT��
4�;���U
��TJ�R��HUD�*�QEQDTR�(�	���(Q� ����A6�	A�m5����hU�jT� U�H� �Ҁ�lS4�pa@  �� A5�  f � �Zi[��Kl�*��L*J8 N\�(�T�V!mHڴm���Td�%1��2��Fʐ����$P� suh���hȵ�)l�%&�Y���m� (��L6[U)"Rb2�;���[-l�e�IV�VcmP�J��m��R���[
14V��ճj�(�1��UV�8�*R�-����m���SJ�T���jY`kh�*�Zm����@�[XT*JũR�n �Je�4�)J+fR�f�Em��hhm�m kZ���6	�m��cV �+i
��ö�ʕMj�+`k&Ԍ��R�E�d�V�
�d+"���J�6�T[�i`�j�h4�j��)Q���UI-Qc"���U,!6B�7 t���@�P&�ZcE��*��Y$ha�l0(�w��@( E<&m*�"��h��a4��0�%JD�	� ��	� IM�mF)�Sh�L�4hf�jB)� �%5#jz�@     T{*<��  � h  ��B����چ�h�A������c�����x�苿���o��{��_e��*�TY�ޒH�4ȴS�"D!��RY�$��$!r0�)�U�rI�)���_Ο����Z�!�Q�����S�QBL <�AA�M$������ 
uH��.6َ#��Wg�"!9$שr��^��'�9Ѯ�Kά����פcrŖ�J��=��+^����ՎY�c��2*�ѷs>P�;A��O�n�ø�U�[t��V�J|,����ʆ}t�j��koC�l�ne�*�����\Xɠ�kw�R���H���yj���?e&TJ��WE�����/ᖒ��({����M;����C8�w��,u)����/�u&��S���K�h�f%,�v�볃#8�ޑ��[6OSR��՘��g嶵��B1��7,��H���	�ٸ3bPB["�ź�cKK�n5�۴n�x3r^M�Pތְ�aF]l�]f���k6�a֚����j���*�8W�hP���42�<z�;ԕ���%�1T���Qj���t�zu�'����y�˭,���c��<U���H�i�����k4��wɻ
��L��\c-b�m"5��Z�ݷ/q��yf-7j!RM�j۬T(⊈o-@����s5j�o��w�<�{�Y[L�;D�I'��w�H�͘�AmM��f��Ě�K'f��3�u��VK��i�F
En<ͱ.�4�r�ߢ�A�M4*��'W��	u3�t�6p�;9\]������V����4*��ַ)��v,��V &�3,w��j.[�+3%0� 0jS/���/Ne��T��0��Z-�Z�D�N;��K��t�Z��(+�}z@�x��CW٬�K-�w�3cǆ�ե��g-��M�(��vZ��0n&�\��<��-PʷYj2��ơP�\��t�em����ˤ�XV�چ���D�ӛ�VI�f�6������Z�۠m���J�����_�:�eZMMhe�ʆlLh���R�K��+vĠ��Ù�a��;���%��G��\PV<۸෗E��`�V釅�k�]\�F�*)]��R�ܫ
"�]��j �A�Xp��u��+��3P�9-��|�GF�QM�x%�W���f:����Id�q]����XV��A�h���J	J�o0�V�����۔��;H��m6�x����-�l�wo�/Yŕ,�ܲ`#1
�	*���R�P�=5m���v��ct�C��ջ�0�.e��:+�31��z�i�^*eU�n��P�Z��V�I��J-^�ҷ7y��rՄ� wm��Fr- ��P5�q��U��l��l�ض7�u��a�v�{�4��ݫ"���<t�i�;�]hWt����(�,��թS0�KT�e�.�f	3q��C���Ř�/)S	^'�Ŕ����\�����ף�����o6֛f�s�Oe��۠d�Jܼ��$`Ӆ2)Z�$�拔�ݺ��R��J��*��H�R�b���R�n�)yLG�:ݚB�h<�A�B��&V��n�t�Q�~�W�t�wʯxV���E��%V���EK4� �+H�,�x�0�`	jZoI����Ԇ^ɪ�#S	��B-�̶B���m.>�z%Z����ԇ�`�v���Z�Qf��Zw�M���Yʂ�,�%����h�sm����4�
�]�ʴ�sU�r�N���%=f�k]���Bٶ�F]�eP���5�Sɇi��L�V��w�.�YQf��ݛ�t�ٗ�3i�[m�=�S3j�Ļ�4����|^5��b6E��o���d���>Ё�j�Q"�ܻ�@^ u�v��K'^�xI�3�B���5� �X���(�E�q`�tcDemD��ެ�ЫT5bk�R��T�5����O�V��+�:�Hu�$^�N
Mo�L�~��yvUm^}4f��C�@U��ӭSF�V��@Vj]�Ŕ��;St��B�m"ؠ�n�e���_;Hf#p5J�l#��3LV�Τ���#�W�,e��E�5+-�yzf0o.�9�,�,]]"#n�v�9j���h1b�|�F0�׮���Y`V摌y��a�sT,`�m����Ũ�Iyu����Gn�ds�����,Vl:"��V�H2'���K*�n�d�&n�p�8��!�D��`�Z{$����<:,��2`תR���M�pS���=�]�܍���ଅV�م�ǊdKH+ݶ�Ua@-4%Y�ge;85����^�2YӀ��n�l`�R'�Ug��Ŝo3B�k0V.}��W`0Z�J Z:�ҵ�U��Vٙi؛�J:J�܆�vjI`u-��ӎ��J�11�V3R�h�-��mV�8Fiu{��Jˀ�`I@�r�a^Be�C���%����n�VuU�y��h��x�����SA���W��פ�3Y� �
5f�*U��h㵗!��%X,i�l��� ����"��*A�Z�Z�ͽt�_\4�7C�=ĚF�cFX���00,z�eS��Ę �V���5a����-����,f�}�WF��ۮ$�AT� x�`����:��,��K[osT��͕��Se�W��-�iT����(�҂FQ�%	ӏM�݁.�$�L
 �@'�vC9�ﴇ�-vS���7{17X&���t1iL]<3T��')�-Tʷ��� ��@�ѧ���λf��.�if��\�w�Ԑ{����t�H<����}�̀���!5��ƒ�@�;)@�[�t+�t�%Ru���{�\��z�QZJ�	k>7�e�^sl0Տ#ۤ,!IP�sUܭ'U:�#��J�-��+��,Df5���x�W��o%���)��ԔX4H�Ǚ��G%�wwYMX�����e3���-լ�m��&U�Bj���&7j�!�_�^j�1M�q3un[q���ɴ�x���+卾�tf6�i�S�k1+�;"�p�Ú�;/X]\�n�#ݰ򄛍i�iH��V����;ua��M�{j^ܣV yuPO�7KuQGq[�e���"V�I%�t+i�F�2ɺ:�+LSJ�]�2�bTbQ��R�
�#�1%���|Fgǆ�`���{���5�8��y+�B�wե�e�0�� B�<�]����l�F�J<�V�ԹW�/�!�A�@����Z����0\ڽ4/V�E�+q�,L��1��h�a�$�|���ay�UӠ��+7f��a�I�c�8��E�B�m�Uye��RJ`�
���Ȯ��Nރ��|�[��)�{�Ɨ%}G��4@�p���,k�(FR�b�M�ʲ@+A�#tHa��h�#�Ԗ��)�Ţ���YŖC�Z��Q�"�)ʽd�N5Z)�+��:�a��YOuf�;���!;r���K4�̧�4ROh"j<��AM�Al ����e����
�K"�+����e��OU2l�\)�J�,tޖ�]Y�&�$��#��b�m��hF��j�X�,���Cw/6��7�X�������F��-����z�MC�X�a��.�bL˷zPn�-h�F���4�&�W1m��o�/���.���7��^r�e�GG3�h<,��Sws	uP��{�s#50�BN;-j:�n̧i�hx���D��r
���+S� �Xu÷�+V޲2�ې^e����Pf�ec���$�^G�7
{��?jR���Uj�Y`j��V�(�`���0w�*<0a@�2�Iy�yzk�K{�;A^g7�tՆSB���C�cG�^�8�(ʺ9����"7Uѣu2;����`	qEӈ�gp⽆�G%LݼD�x�Y�B�,Vh�vh��a��d�;��`��櫠Q����3i���Mq9ԞkzNq|������s�w8�]o3��κ�[����PW�O���{�iʜ�:+���,�)*^u��Å�]R��Q�D	@���4 ha����@�3DDD        z<���G��V��ګ	���PVv�                                                                           @  `                                                                                                                                                              �  >Z�eZ��N-�tp�M���˱�Fm}��`G��:�5.�ޏ,ޚ�C�q����Ζ���f0�3��$�)�9�����:�����ҷ��їWQ���m,QЭ­�9��wX;�C������a���۠��Δ1�[̲��i>)�yP�;���^�ou���rpFve���Ϯ�ۆ�i��U}�C���<�Ov�YFwc��ٵk!4J�jb[x��Ηz�Fr�]N��f.��Y�[���\잘��"�ufΐQ�G3�c@!f͈os;:����zm�����n6r�@�h�ω�����B�nũ�zmKX�u(��h�3kN�H�\���L�ʒ�}6��oAK5��T�d�6ù���>�#.\Y�-�i�l��ܥ���M6��]eT7#�����L̮'q�*��P��.n�����ʖ��3*�&}��1c�^��6�@��K��6��Z��JݫJ(�tS3�mW�za��^r��%["��b��N��M���f��!�H��f�b���D5Yi;��o>zwz&�]�tk�he��k�Փv�4S��U)��U��:)WU�#�+/*��n��J�J��_�3���wvS��0���٦f�ܦ��'%<4[���y2��D ����`9fr�qe��+�]ݹ�gGC1�B=���5Q�ͺ�!�]��0q����vVVTP��2d��Af�X.)�;JW�c�/4c�ݪ0�����o]B�©�����oVP��N��
�d�F}��y�������9lʐٖ{T�-�T/Z�	QU�p��aok�EX
�I�G��B��p>��a�W^:�7 �h�cf�;����֥C]8�y���+R���H}�:j�Inoeu�M�y�q��n-��g��9�r�[s���3'v,�\-+��"�)׏z�|I�ൖui�k�������`�ׁ�9R!��τCEO���v�4Ԛ�{�g�2�V��&��,G�;�� 7�j:q��[����s%Yw� �ƙ:UŻt-�yAvfw9��Ġ��j��xyW���t�x��7�5�m &]�v��x�p�Y�pahب����e�r�ڦ�����׶e���&ScC�u�,w��T]���,������,J�p���GC���n}}���S������!�3ut�8����7T��;=1]�ۖ��e�p_|v�E��U����C��	��n�	�̽Pg@idV��ؾ�c,Ζ�W�װ-���t��pd��}=�Q<ʔ���Wol�<UN:vR������7g��R�k&U��r�ѕ��Ōp{�z,�Ͷ�h�q��2p��Lhz�������� �>=wڝ�4	�rnݲ���Jp�nM��}�X���aUg@��������3Wmm�]�2����f�����|kN���X����we������r�AM:�a�r�Qs��jh;e�ᕌ췈��:4w�[�e���Ի͹GN\=|�ћm�'X(�Rü�(���l��9��EC:�Y�����tyr(`�|.�_|��OY���){&9:�wVs	�$�k�3��тu����q���Xv���w]!�J��n;���KXTk0�H>�^��
9��HJ¯���U�cW�3���Q��Y�l��W$ǹϧn���F�3�5��9��Z���7�3��Ao�U�e�]��LzkB̚kw�#�	�
�w�`S��K�x��n:��f�C��MZ���6u���"NX�k.�W����^�E�ڇnW²"x��M*�JM��L
���_>��-��;iW��>���O+]0��޶�7׵r�B��V�fq �lPM��v)�n�/-ue�׹�QԲ��`��S�AOj�;�I�s+!�p�6�\�[t��;���o���5}]���ËN7Qy�ݓ�Xo(��j,�m���϶�K�wX�F��Z�t����Ϯ�n�n��ZX���-
��a]{7v�1�S��-<�/Gj7��1�	�\۲�+nT��P� ]X���__q���D���I�z-��mY������3D�T&/h� m���Jx�,Ӵ�-�#o0W2]���.��Em`�A٭�*�S�8�N��kr��D\,4��u����ԝ��M�Wx7�7T�j�Z����+M�7����'���S������J6���՞�@6"�S�����zi��P��5�d�SI۵�E��L5G{۲�����ej67x�ؕy�I=4'wV�[**�֋��8<ޔu��� ­qI�-o1}\�s6�{�U�3h%+	��v��Fߺ��8t>���'C%�T��2��+�W ӁN����^��_m����z7�rWV7���-v)v�p`�������,���w2,*��d�(H��m�jiթ_XVj�¾�
��Jk:�d 2�a�]��d���#њ�H�n�m�xTbp����]l�0��u��&����F_1�5s��6�u�I�\K��<��w�fc�t��س���Zյ���9�̡֖ALM�tx]p�Pc��m�Q��zP]���5\"�d�<��o(-�.���+W*�Xk �o3Qv�)��|��"��^�#�}B�4���8�!�_�w��-95v�<���� ��4��Jf�oHE�9�u����0��*0�s-�I�o��Kα����eZ�x_k_lu|�+}��P��:&�R�72��!ȹ>.������[qR�x�;��sc�d�j2U�/5�a��N��C4�i�G0�ʏ@o�0#+ri�&b[CEv���c�k-nd�n�[G�OJo�1 y7��Q�f����,���Τ@�Qy�*�s�ޖ�ۣ�[��ii�ill���%:d3��oY�+�'W|*Ѩ4v��XY�G,���]���;��S�A����
��YҕXj�j�z(��u#�n]d�U�WoN�p�cˌ8x01����7���Yՠ?�oZ�K�U� �f]��U�U�Hw�\'�T
�7:�vosf�6�K�At����Eg��H(���)��&f^L5���cU��(���^wEN���w+HUd�;-��v�lX�k4{�k��mȹ%M�Qꇻrv�Ѽ �dM�X�
�6��$���cr�-Ǧ9���Z��V�R�#���[��'���%R��{c�h�mk�ܙ��	Z�:+�Ԓv��Y3�GG>��;{�e�Շ�Z�2�FG�-����`�a�:��[���M}���Y�B�e�lʳ\~�&GK;6)����2*j k�nZH��o6�1W�<<�Wa���7��B���|��rQ����fSfA���5�[�Fk16d�;�v�n7��Pݍ&ɚ˭�굷�������k���nuX�O�����u���5xx\�����m�����3,���¯�e�>�DOhRW*��tc�݅ˋ�������n����D�*U��5�G)��r�l��V������L
�;k�����8Ε��Sv���7-
�L�qaPƱvΙ�T�V�j�Tz���&��WK#K�\���TY����7�*D���l1�            s���nNO�ll)S-t� U���#����h�H�!K�Qw���c�tnH/|���O��A~��Z#�x9]���  ��            ��z�;��k�kݵ�ܷT��H�_dS,o����촺H�h�M����0��	U������w�w�#��Y��Ѡ�����\�G	�E��y�^,Á�\[x7�(���F�-���֩�FI����.Z3��w6����J�r��U��w�b`��@wl��.��]��]���,��n�r���34�T�:�b��ͺ�Im��MS�s��u�b��++��:J!����[F�@���j��s�a>�cE���hpUW-m<�)_K�Q:�Ǵ�v�����ʆT�M�9��Ei��,)����	�3�ٗ�h�%����_]�O��*$+�c;�A��2��R����3�Bp;!v_��iq��R�����e����^T43�3�f�E�/��X���Ӟ���ae�q�3���0D4f 3���Y*�=�[�\2��k��'.�S���'��M鼔��J�S����-��Ь�4���;9��B�CY��#vĻ;f�z�VKH@AYBS7B�����������P��S��@-��6�ehǈX-g2����0�)�� �;w<.�N�Ic�� \���l=�[h`O��C*��MCO�S�>TrG+`��Z��N8�t4��޲���[����I����x��-<(]�U�lq�wxa�^t��4o�M:P'S��s���ҙ7-���q:�J��$_n��|���d�N���Q3R'p�
�:[u9ػZ��`��5��m*���0���r�s�Q��U�*f�&H��8w��`�aL�C�l�i�����mҜ68Q)h�)љ�����H�qֵW
�o4$k��:�����d�b�V���^R��Qs�����n�v ���	��q��r��%T,��1k�&n;��B�W��լ��=y��$i҉@Pm���|]b8�I�vm�mr@�ʁ�I�[�[R�V��
�j�P��,v|l�"����Yj�ծ>+35������K���É��H��7u���l]@o�5ծٵ�5��c�T�A��:�J�*���ǔ��ڷkxn^3׎ct~HX�R��P��i������>�9[�-n��X��e�8��+gj�śYI��Q��2�:zY
�H�Y�kO!IZ�����#�0[ܾÀ��ZTKGi��
wV�Z2�+�CN�&�$%t�i�lvk?�PJ���9��oa�q�K.^	�;����H����{�VK<oN�l��e���Y�*£Q�d0��/żæ���5yװi�JvwT��К�l*3�ޭ�>��	�YnW@1$ƍ�e(p<YHf�ls���� 9}�f�e���,��l�X����K.� �w��w��)Խuv�Kpv,HX���1��(9)��$�Jm�9��kP!LHZ[O�W!ݰ�٘�����zi�ov�[5�ӏni�����D�9������D�
�U�1��i6�����jη�t���8%*�A��<�Ob�X����Ɩ��Xt^�g<�Ӌ'Z#0�8E,Y6����,صwU�dި��Ǚ���V�Xv�Uޔ���[9�8�"���E��:w�u7]J�8��u6�Y��������S��(���Ls�D�0(���Jh-(�]�iir\��{���1e,�g��Ek3�v�*'Pޱ"�{Х����l^�`��3)�����[���"�k,լsLĦR]�|�,�s1Ŏe;�u*ڼ�$��3���X�%��m6D�n�]Zv��W�O�P��֢k{
u�K]V]֮S�88�p�\�����5�n�=F�K���4�U��&ࠞӸ�/~��E��I]�]ӫ�&}-g=7cS��j�t���}4��K�;�+i�V���c�u�X�VU�W�5XfvR3b�+�GJ�Y�hdݝ��!]f+6�e��G������%c�4ڜ�-�V�����u�H8d�u��hE.�꾒к�)���:̐�4��p�w��)�#��O_'�6L��ٵ��Y����(��Nf�[\�+���%覧<�7���6:�N<ޭ��X��Q�o>���dUn���n�M{7�뫨�a��4���Ks���I�;ePC9Ag*:�N�fWث�[uǒې�ZI��+Pp�y�9�� 3�j��B�ʱ��n ��\s�xȮ�Z�`楜��.�V��ٵg��@��Ҳ�5��a\sr���A7eR�.���\Zw^`W���L�(����h�-鏝���s�Rچ����b���\�:�J侃r�M{�!߬���T� �����L+UWS�۳�{��z����x2�9�Y��|	�u���d�'ƴ�.#-꭫V���o��	j������˩�wbL5.�����E�Z�ki!ʍ��F&��v���+j�M��٣�q���`A�f�������*�F�4jv��f"v�����|Q��X/�rXY��U���r�n�eQ��8ȜN<r�ܳ���'Rd�Lef�dZt���)�M��gl�N������I	�R�R���I4�n�ǰo	�[���A�Y�,���<A<�J`,K���`��q�c2^��LsN�uT���*gQ�����2>�`�m�Fe�:	PLU��)�Ų�t#<6��R
��s��\_m_Q��W�)�W����������B�+EAw39Z�P�K�����o�$��t|�T�xI0�{}\M�2]0`=P��"0F_�K�mD�J��x�"��=�f�gm$�:2��1v�J��t0� Y{�0�Z�uԮ��҈x�]�����m�K�5a�������ɪ��Ҷi�(/N���g<�� ��ʩ��%۠�e�1
�we�r]�MG�a"�R���X�S8�h�wݯ�mVMޫ�S2;Q�B�'-���׎U]tyV�x�V����q����Y�z�Rt1�w�����֕].�}�Я���k�r^�xɝ�R Qۃf��բ�3&*�kfr���G
��[���u����I�k.���6�4�j���_PJ40؀�Y�j����V���y�&kg�uP��B���
�"gb9Fw��-�\zI�t�C�1�Ծ�fMr��D���u��>G$(�A��*�{f�r���jGz
��)*''_#����w\_iU̇z�aH�!���cL�d��NTYH�S)d]��fȗ)�r�r�I�W��]�ҝB����fh���at��Gc������-�CB��=[�T��o4��J� �t�Uo_B*��v�U 4�W�ǌXi�B;����k�����-�ׂ\�y�Qqv�(|_��!Xt��:csy�0�Қ�r�b�q�ugh��� ��v�lT�V	")\%<c�Pޕvmi��Y�|4t�M�!��(34[5>���S~笻���2OeF�V,���I���J��JÏU�6�5��zvj�^�y,"8(5b��M��,�1��fj�~|v�oP$_<껗B���١ �Q�T2\q�r�[�]��'.�P]9��*h�)h8�����J_Z�)1�Te�u�r�:���CV]���2�Hر.��rt�I����i� �W�����|.�n+ݙ�ip�Uyʄ��{�d{��TU,'.c�D���#�}��#ul?�Fv�Tj�e��x�{�C�f�;��tr��ѳ��י�-N���:NM-뻺�|M�ۗש�N��[��ȸ(аr�������W3f=��]P�Ь�8�iiڎ�3Lz�~��Gـ+m����=%s�X�0��w
A�N�o� ��]\�Gm�L�-O�Mf�7��� � �H��!ؚ�/��!�(+��hp��Z����Q�g������                    5ݗ�]�L.�ƻ�Tkf�|Y�]=���Q넓��#���̬�:A[i^��oOunQ�����Y)>�8�6�r !���&����U1E�Ԯtl'.�W�s��խH��+X<2�t�D/�cR�J�)�gk�u��D��s�����-���%���EP�Q�sS�hr�
`������ttj9Ga�7LJ\�ur�6Ui��I-�o��t{+�N�d��φ�tֺG�ݻ�v���wOYU��ui�}�����X����F�J.����GVX��C, ���}>�;%lF�']*��ȄN�[:�b�0��:5����M��dr@�'O���oL\�M�������wE��2�ѻ��ٽ�ML�m{A$�9�<�کѨ���ֈ�'�p��)��F-1DRP�@��ADyU[!ɤ�L� �.�(�F��#, ����"�����J��AQ	R����'"�
i
�N��Ms45��3@�U%w�q'��4P��#M$I]�$KM%4�Ap8K�8����i��
_,�j��&~�bc�O�Uf'���!�T��^�t��/���%|��T1Tw��&�Թk��>�]�����_�}K�/M����܍���,nƑ���o}:����+�V�/+s��F�{�a���4Ð��_[UUu���Ъ%k����F�AL��+�t׼߫��?w&�6o.u�9�T�wѿ]��|��T	�9x���6_�`}����������Ab�1y{���Nھ�x����E7�����X�7��#��,�B���~횼Z�3��lX9)rI��jr⺼!GFi��j��_�������������=V�m�cT���V{��ζg�%�4�ނ����YNn��	���V	=}�R�p֐7�wi���=NHM�S�s*�6!�)^�oV�}o���I�7"��T�,���www�����&q5�ٷE���t���X1���>��;�]�r�2c3�v��]���8�'���[�}�E�s������-��ks��ϗ����Kخf�r�\������Kb䧴zx5t���z�eh�.�$U5^�m���8:b�ӱ̽������l�BRE�C�wPu�/ݚRf�};<�����)���|��4��>62�^���g�^]A�ҭ�m�+�!<:V���|�\eN�YΕ�����t�y���nĪVM��u���V�f�N�Y}h}�jT��F�X�ٱ315̸�����X���]�nm��T�2�Ă��Y��c���]�U�����i魉��޹��b��uw��)"����[����6d�Kȯ��S�?J��w	s���Ź��!Y�Oj1�D7G�k��O7�K}E�����(�v��`ZL�CG8�3�kh�=ڷ���Fyo�&��{���Y�}�$����V�񶅙�.�fkm�'���nO���o2%;�O��-)=([���_x��{�+.�������	z�ޡ�y��o_���Xx����`&�~�~W:��w�=��tc<�7dI�N���׎� %�n�QJ�i���#Rh��7�8�nI�c%����W��'��?E|Ϸ�3]hأ������4ܲ��Ь*�[�����N�`�2y��*x㝕aSi�����Z�y�v����[jf���f���:MGS˽U�����d�f��P[�=�|5
�Lnu���g��'7������t����Wu�O�]
��1c�\w�%������#�/3��V�����=y�/F��V�,<��=)8��ﴫ��X�ءS��jǂW�N���G�6+_���U~,�=�Թ�ņNS��羿)j����{cV�}[[��lh������݊Y��-���]g-��<�ܞ�������	B�T�dйׅv��`���7�ǕgT��3{ݲI&[�*����;c�7��13�h���米���9��F�=���x�}J�?;��.-�S/�����^�G�g&|ߒ�<�%c��!t_�鎅���aw�����cW+�ũN�GլBTlB�٧���}�9�<�пn{w&7݆o1��gާ}Y�\3�i�"v�̵��I��w
=R���o|<��*�5^ƕ`�3�৐g/�i�(t�ek�t#ߵF�g5�EV���F��k�W��+����v9�zU�S��[�C���#G0m��P$���}kd����=R<��-�v��9yAbӹ쫏J��!W�l=k3��ya��c�vz���)ω��t�)�usW����>�����PM��vԻR����L��p�����յx��a>ޛ�Z43_)����b��5��V�Y��n��}�IAwz�����5�aJ�K�O���]��O�|���ޫ][q���=X��+�}���o��R�����g嶞U���yh��)y�S}�ȸ�?���ګ�)/y�u�؞u��4�}B��.f:��M��#{�c��W����~B\�C��=>6{0��gt�ɓ�Yg�����/c�
9��Vr�,]�se�k;n����Bhv��y���T�l���a��"���O6��NI]	|�>�
��S�)y��C��6ѿ9��Vz���X�η�ѕ!�^n�~�%8�Ae-��-y?|x ^������lRr�×���喧��͵�������T��v�e����h�oޝ}�ٖ��o���fW����l��4��~��������(}X<{��uj��Mo&-�yy�a4ͭ�h��K�w����`�ߟ)I�)�Ý�0�����B��N}و��-�|W��x���-L\5�T�����/�丶�f�V����ߙ�3�;�H΍7'�C]A���{Fad���|bn�EAO!v��w��;4aQǳG��^1mr�<Q�No�Z��ߐ0藶���[tm���T��mŵ����~m���>8��~�[T�e\����|�)+(y����OTy��t�W}t��j�����K��9?G�t$�J[��~��dR1���w<ǻ[�6�$�^{�SMR�*�[�6�5�����z2�߮j��K����g(����L����M�f)�b�B�E\7��ܘiS��r���
j0��5��Yq�k\&ECou�d���=o
�X��邌f���Ek�7X�d������sٔ9���w��E�,��'��;vu[���正��R���6��9��q"�y�̯<�ׯ_*b�����ZNM�h�r^ ��>���d���S�˾5�8|	���͵�Ǐ���45�+��
Q��=���PPV�j�Yމ'x��<b�'�N����Ҏ�;�y˞,Q���ױ���old��	���ͱ�#�OF��)މ	b(��X!V�_){p����Fѯ=9�cy��>F�r���ܖ�/y��ljv�
�9̠c������ݔwS'��������$t~"�+=Y�/z�=ݮ�k��_ȃ�2�b,���ce����E,����|�K8n�Q۳���D����<;ǻ5]@���;��^����qZ�=ѕ|3v,zM�������7�S>|(�F�x��ì����J���km�}�׹={Nf�E۳n��W��椒�N��
�dXF��7a���g�aɹ��=8�I�^]��D����k�e���fM*�j���E�j�[�M��*�r5�eN��Q���)8�Ǻ�y�!��M^;��Z�Vi�y�/g=��c�^�Ͻ���f��F2)\�����%�}����~�VJa��f���J����>��W�xc=�Y�<�J������:K	�+�Ϸ��7.��1E�ܺm)N���J�͝��TC;2p����^���_=!P����HX�mf�I��)Q�Y���	B�]�a��*��Y�LA�[7�+9i��V�^��4�3�1+s=�y֟g.���A���!�8м
5�шq0V<�X:�uz

�Y'�9�P�ޗX\���,�7��d�x�&φ��e۴:X/��1�LB��;ث]K�d�v�X���e�RI�W��6�\�z�	�]�F莾����*�sn�<}b�W7/Q���(Lu3�̚%�׺+L�y'��$���r�-����Y�t`خb��-�1���3��&��8��1�,e�4�`�"��;���e��� �Hf:�k��u�����8���_�߁                      �쵕���E�F)lZ��:grs%�Nr:tW�v`��#��r$oK5�Ia}jl�]�2����}y�_L����'(���1���	��'�r dE �>�L����A
ُ���ŭ�og5*u�wt���Ʋ���@!1*�9�����Wm
��+3���e��9k�{��*�n���u��n=�ֶ�i��L{����</#�u��Ş�)��:X��أ%��^b�P�h���
�+����c�o_�-�Ow-�3�c�������(v�ֲ���V��8ʸ�4Z�aF&_q��.�WRZ�HSfh{�r�=��OWu�-��&������;;%g��!����G$��q��W}��SQRD5�QT����)E49�ETJET�T4�Q]��I@��/�h�R%(k�r�h�"��+X�������e4��q:J�hij��H��9�*(�&%����,�J�J(�$iZH�H���Y�d9'�)IK��w�%'q�I��4�Ov@S@RQEU5�|��)hJ))*"�F"�' ��!�/:�
"�,�T���S��;�������²5%�\��8tOE�[O%�e��c���v��{����ڧ����S5�Yˤ*���z�!֊>��~ ߓ��l#��\��X�(W�X�Z���e��O����5s��}���gg��/Ȕ��ॺ���W�g�y��.ς��z펩�nU�#�;$��oLb:�m㜭�� E�3�7"oߦVx�~���C��O�����{�D�ΏVl�p��&J��T�}.2,[������5�8���a��Iv�\9����s���}��SX�0�l+���~���;��?o�|ͣ[�>�U�ݜb��W����F��n(.+��	su7f�=f�ڻ�T��V��S���R~��������U�б]�X���HS�"�u�;m�[M7��d����Y�����]���}}�(VS�g_�a/?M��kk��Ī-M[�����sU����q�"��|�l���ޏa�sr��W�EI��؅MJ���uQS��M.�^{kݧ�n~����`U��[�������bjOe�)�����o�6*�����[\h���ˀ�+��S��1W�W~(7���q��ͼ��S'����5^�����'�����ġo߾���8?�[d���J�Q+�&W����ꪂ��o�~�����e5�
�;��!m`����ުhֵnxoJ暭4y�����To�	g���{ޢ��I��ܟ�j�+��؇7SZ���ٚd@��F��>��S��G���f�b����� =qЕ�*vO3�ٓ/в⓾���b�v.POz�����LC%r�S̋O/*}F�Gj�lЗ�{���5\�����!6_ü��V�6��w�<�S#ٯZ��.���y6�o��Z�m���x+��o�ך�-K�.[~)7��B��J��^*we���z�s��[��q�W�+p�U՜�H0�����!��k����aQj*���=�l�K��T���Q��ju[�B7��C�v��,'F��}m;Awi�;��]���w3��4��/xanv�^��y9�gf�X��6�k,��+r�,b���p�۫�;����|������ǌ��?-�s����X(��r��/�m������CynA���򽨰���8o<�r��>��k���p��v�U}����m�����_��Lx/tT�V��C���[�s[�];7MU<�*ъz�f��m��I���>�s���}��X4��ڂ�zA�cS�ť^{���G\~.@���1���ƻ�w)���97�}�xy������}��ԧW0�R%�����By!A�J%��Ц��K����B�!�������\y�?o��)︝@�X�1�0�A�`� k�=�5�<C�>NA��Ϛ��w�A���E�w�����r~��U�9����7��us)�����`'3��܅��K�<K��ʶfu��+ߝ�+���~���>�vt�Ex��S�\��٠��k��ܐ�z3�
��-q���!b���.�3
��o1Ģ��h�}U�;���ﵯ8߻��|��aOaݒ>G����#��:�7ę)�y��=���7��ԯ�8y/p�w��z���>�׿{��̼K�x?���/���%u�{!�c�B�}����O%���}T(j��_x}\�R��_E��~��W�'��̾���;��p�]k�*h����9�Hrf u���䮸��ם�{���;�������'#�C�;�.�w'��>��W۩z%�V�#�'`s9 h��CFa�]��k>��<�����|���)�����p=��s�n]���{w(nC���w�%��;����ܚ�{�������������>�D�w.J�rkr�ǸK��u��x��è]����=�����y��y��|��|q��o�7��c�)�f܄B���7j���S�0<��:�=��y�܉���{���f�����7����(u��2]��{�w���=�q�퐾O8��=H��!7#�zw�w�w��<���w:��� y.�ܯ�h��
i�ɒ���]��|�����$%+�K�>�y���믻��<ߦ@I�)׶���qJ{<�<��|�7����nL��3r����jS?}�>�0���d��~���K����J�����*�� �O}��[���G�ޑ/zx�w�:�5��d�9]�����;4� :ڟ<��`&n�5 �g}y���� �]A��)^�k� ��7/�����M�A䧓��voB���]`��\@u�<w��;�����]����=Jk�x��8�䦸�%r2Mȕ��	�O�=���p�o�<@�s�~�{������<�˗0��H�!@�j;��S�0>�ܜ}�s<Jps�ɮ�|���=�9~��O$)6��>��9�����׾��2���W�x7Η.e{���C��� �8=�MG1��)����d��T�����ߚ�������7!J}�n_�%�^���N:šw|�{�������܎�15k�^`�Sι�;�/s�Z��|ߛ�C�>�P�A�{/�=��{/�0�!�.w����l�8��B���J�냿x�7�|�����8���S�s���w�B���s#��/��
{y��'x4��\b��u�W>{���{߀��N�au�y����'��{��^��;�ۙ����_���>��3��^�:Dؓ��V�d������P������&�)y�ܞ˹:�ܾ������x�p��zW��~��߼{׼��|��s�ܥ-+�X'�}!��y(y.B�d��ܧgا��s'X��}�h��_}/�M���>_�ZL�d�˛��X�zg�߸�r�U���cIG��Zf����o��ߟ+��P���3l�z�'Y�1���6�_3k+9��_4���B� �;�>y�� �P��y��=���::��2p���P�>�s����_�a93�_��<8���k�8߻�{�S�w�éd|���u/Ч[�2]c�2 ��ܛ�����M��:�\�ߗ�o=�~w��K��O��.��!y:��Gؽǲ>\��Py�����HR���=�q�w������w���~���9�y���S�qܯ��rk:Շ�>Hp}�jGGx��]�䡽b��}�����ל���{�9/2f#ܽڎ8�w!��M�����\���}�]XjD��(<��w y.�לᫎ<�}����w�����K��C�/s�)�e�^����O9�.NA��S��S�N����q�{��o����|��(5#��)I���H��.J��ZZ]��pk8��e7)�>�;}�8��x9�d
s]{������߫�.G��̉����y/}�@K����8�x�R����s�*j:��w��}�{����瞻���N�u{����)OgP�/����Ϛ�W�y�-�k�wRf"}�g_}w�9�?k���~o~�ԏ��j��:����O%O�X��%7!����0������!|���\|y�ݙ�wƞ:�<[�����.��8�{@�O�����Lǚ����e(�����Vo%Iǘü�v�"�*Q��'X�����ݝ����䈅 ���|����:������=�MAܧ����u�R=ɹ;����w#��˹}��u{�;מs�u��{�|��>�- f�N#�N3�
=��]�}(vs�nB�$z��:�����������̵��Ͼ������W�:�Oα:������]HPp}H{��'���1;��w'X!���B�U�ߢ��~�f���R����O�wu/��w������M���<�=�`�v���=�H{Ǽ}�q������R�s;���0�D�˩���|���ޱS��SrP���s�M�rn>��|�w�� |f'��)��7.�����L��H�^x�<�܏Q�C�;֔�u�����ι�޽�{�^�=��N��>�<�d�_y�;��M<�H�^��k����� 5���<�y�����{��<תd�X���<��~��`'��0>�W���Mu���]�ΰS:�� 8��*��}2/�����f��~�o�ʴb��\y�#	��~r$�xѤ}���m�y�tG����������t؋\@�*Q'7Q�V\� yԫnj���Κ���,�[�2+0���J�̽���J��͍�N�5���R��}^���������������rz:e�!��:�#��L��l3vML���yl͔�c����z�� ��^g����Ěw7'
�Jv)=���5{��ȭ�:���|6�,ݞ�*�ɹ���A���g�S�Q�Ny�O�鹻�l�~ɫ��S�Z�����oq�뇋~|��{a�PFh�f;�Z����MP������޾��M%7L[���kW����;�{��O9u�u�<�d�=+i*� ����F�r��36���q�튽�%��n��U��^����{VUآ����ry/OwW�p�ވ���%��o�>�#�pPs|�l�*�8vU��7����@�HB- ��P-(�H�-!JRSIM$E1RZ�wמ��c�z"4*r�]��N7�v�(��Ȼ�����7�+{�*[��;,�'#]���t^��/����/��e]�X�׷+�_�/>|�te�G���'2��Ǻw���콝������/g��܆�Z��h,�m��:����I(u�x�����U�^���q&�q�72�j���^��ux���-�7p�ݻa�9Y�\(�m���߅�d����P��[��uu(}[�P��;Gه{�5ȃiU���fhfo"{%}�9ϖ�O���'�����y#.v'/�g�黹
s�ʺy!wD
�)V^r�Y%B���5yB)p�I����ԯ$'�VX�U���`J��ۃ`)	��ڼ=g��T�I	�ڡ��Ns���.��TFJ��8�i�5M�T�"����ι����d9����}4�E�|�8	W�]6o+���%��Q�'���l���i/H�l���;��I�V;��%kj�u�4� ��rs�H1��6���5�VY�x@����&в�Aq&�u��	�ۜYķ#i��lC�i�ah,$�#�(<Fɔ�v<gB��qԧח/^�m�$���]KUJ{��ʂ�^EZ���e�����pf��=��k黗vt�{����Vl���=�&���X5b!��b}���ڑz{7ՇF�'������u?��                     )��U�G�����n�o��|,5���o�#�m��vL���|s��se���¢|+U���Bh{\u���#MEf]�HKT_Q�цs�@X�ƗT[5�pOroL�b��T�P�����@�:�%�+�;����CƱkȬ���օ:�Y��r$����{ٶs&*H����Q�[J�۵m��)�+�)�[�Ӗ.�؅��-�.sK	X��t���Z\�u�rR���"�>�G�=0
���t�<�J[�c����$�[�1��(�,~�\�5�`�钌��N�]�^��wk����+9���KB�	Y}�`����;��(1�t�V�E[���E�9�*E�	,_|cNI'G�y��ߞy�������������2�h���j�(R�h���5%)Y�:�-@�RPBd�A��,���%8���\���.$�^&���G$rI����� )��2ud��-�6��"����SI�9%�\ε��R� �B94%)���qB��rR����5%.�$$u4�� ���pYR�bj��wI�
!�y�.tW�U}���>�sޣyթVI�ns���Q�KwF�����Գ�Ѯ�qͱ9�4W󈏢>�-{�p(K7�ޯ3�P�c1�B}_�����L���^���^3�x��v���O����'Pr��~74g���U���]�SAc&8뉆��EqU���x�˛�=w�$�\�-#+���b�~��߿k8@��C|���Jv_=���ܯ��+���Z�����Y{�ι���l�	u�F/;9�VV��݊m���M5��{	)�~���^��7
g�z�N�z��}R� z�s�̮���v���g=��vZ�~�LJ�T����pA�.����kIEYs�~��Ts��p�@�n�>�NЬ,�7Z�Wl$'}`Ǆg��ܮ%N7�_v��}�֯�M���AN����9�7(f�?A�����~$�6�T��J���m��=<�и��<^i,���8��z
��t#s��w���&0J|���jԛ��hD�'�����>�u�Xk'N(��x���\�V��\Ri��C=R�1�ej�������m5��:�TT{Ӥƭ
��K�\�[Ѭ����_�,���)�t��	G�X��o!�݉7�HZy�F�4���3��Ô��7��\������ǻ�'�~��=���ׄn�&yY:g�43a'�w�0\����?���c��iu���=L:�����ܣ��jPk5��$`��(���}��}_|7S����]��{]�b��1��E(��{ux���%}�}%9�k���������l�%��88ټ ��*��;�}��G{��*����6�4��"E޽͔^Z��ύo{x{>�AI�G-^���:�������n:�T�"�^nq�36E=���h�3�n+j�ҝ�OW�S$����v�4�к,ݞ����v_vE6���<WeH7���3ϝ�O�IMc���6�ՙ�'g�������=��/T=S^���<E,��L]��l��>���ݚ������_§�ޏ�=.0����=[9�}X�:|����=�+��j[�3,�cS���UW�}�`q�<���vRB����:���4m�אy�~lk��xU{ׯ<_E+"�1���9�����җ˗F�3����g+����Ѷ,sV�-�P��9�7��4y�����U����$v�ǋ:�~�S���6d�;bOч(82U�P��)����KV|��r=^Nw�`b��YW["�|og�M׋��xS*���aG#T�TW�uǫ&n����[�Ơ��(==	r�ҩ)����2n=N��:��)������fq��S̙p#j��}�c����Xf��(�A[M��լq���P{��;���^�}�9Y6|
�'a��ʛ�P�e����[�}�u����Xy6���]����u5iz,뇗{w��<W��S�I����/o}jeK�)��>�����u&E�V�$̮��Y���{ĕ
l.}�X���g�F銾��/[N�j��zg��/ow�Y����C����y~�W��c�{���e_�C�*��D���^� 4ֿ"��C�:�i=��b\�{�l��Ay���S�N�}i"���|Ǐ"O&˞��Z��z���A�V��b���;~{�ht*/0��ޮ�r�)���c�Û:_����{�(*���b9����Es�c6�<7�6�#�외�����Ɯ�p��]V$ �Gݷ�Mv�|�R�3e�hC���ʄ����_}�/�y���ho���Ǹ6(���<sl�Ǟ짿b����"��U7�Ƭ��s�+�ݚ�w�p�)����^�}�o�քuL�+���U}��S&y�҇^kͥU�(}:�S��yux���saB���;�=�V�ט�i2�-�=Hz���oО7ٞ~*�F,]69��S��>�2��PmE���`�)I����z�>�Ljߩ�}{�����Ϋ����ԋSո��˥�V�ǟZ���C[�����r��@#�S���S�-�&��z�y�ڤ��w���%��r�*pmC�:�h��+\��,���l� ���UU_U`1'<��G�m2[ݲ|(�8؎{W�������ǖG:�nF������q�]����K�~	q���i����i-��z���W����jw�q�|�[�-�Й
r�k��
���Y�N������df8�k�I��z�W���܊ͅ�B�|%�5\�|�����v���V�E{<X7Q^v�(��9�������������`,�8�1��
�]]{�װ��'qʁ(�H���+]*�o<�*i�u��\�c]*T*���렢Y�ڀ�IcH,t/o�Y3�πu��ӑT8�u�8�� �<���t�*a��+7Ռ�ὅ��gj��3��������ޛ{?S����y��;Ѧd�3y)���v��u�O��D���t��ђғ�h������v�|���R�J�aGzvx~���$,{W����Dw��o����wǔeU����3OoTkx���Nz7�_F�ef�E�v�/N��P=Y��uZ��JL�g�oO����Aũ��.9��:�����s��_u{��`ɾ��?W�F>v֦�&�ϳ���mc7�y��lC�>U��i���՛/��H�5⒡O=nz�
��a�\��L)�z+YH�T�E%s#2�Wc)�Z�Rq���QMȍZ咎_6���ܲ�=Q[�q�S�ih�.n��pn76���}��}��$�]�k�W~y��[���*�W��u�<o4���J�b��}���-[��#�7ѷ=��h	�9�u���{!�̯WB\�.���λh3K�\<<�;��X��ʯ�in�L�A8�"�mz�Ǫ���V��.�H��;tCJn��uoz���֊Ƽu8������|�=�}Ec[��uu&eo����F���{�̚��f��:��;ٻɫq'M�^�N��z�1�G���Wy�Ϻ��P���]���S���˗�0^�y��3xs��}�)�j���3�2a��=�<��X��'vh���ъ����yќ��"ʾ��C����a�=?��������X�+�;l��JnXT*���b��\m���Jqe]]G2�< �;���M/f��G�,Ϳt��UD����č/~M[r�������W+�g�_��PE7�fU��K�kZ�[l�9�x�=3����B���F.y^�9�/us�����Zƪ/\��uqkQ��C=*v��s֗t&-�s5�y<��U}��Cn����ƛ��w���en�\�Os��^��q#���<�[(/X��#���x��>=��^��~�ׯo~��'��g�kG��fY��VSd��w���瑸�
��ˬ1CF���S/kY��g��q��jNK�x/GcqIKkw��ۡ����3lҲ�#�%yW{{�k��6�m�i�9'9k.���й�v�.���ҝ��a�|�r�E"�aF�T�k�%gn��.�N�)��\0J�X�n��޸��R�t-����`P��],o:·g�m���HP&��t."�v9[�+����i_`Y%�>fsp��5������t(s��f_v��}��45��I�
wY3@���y$�Zt�*�37:g@�WY��wK���"�V����z�C��a�uy�hK�XoQ<Gw(,S���a�Y	[ڍ�;m�������c�9c�+i"N}�|�HO�� k�����7�Ѱ^�~d�H�۳�'                      ��[��f��nI/+V�*�G�>s;��D����V��ﱥy֨Ic{ʻ^����t�o9�4FW.7�)'lQ�ζ��&رg1����n���j���.t�'(5�;���y��5_3l�Y[J����
�����ΙB����̓�s(�):��ew7�ps0ù��wc��ޠm��)ur�b}9u2b2ͱS�V����n�=�vtuU�/���Ǝ.b��4�#��{��ʹĭE�ХY����*Z�+��G����s{���tT�o*:ѷ�	��x����z��%�çI�P]<M�9�!���|o�З��c���j|6��R띚��z����n�=��TZ��)���7$� @B8����1q1�O�?}1�	�q�d�B�TڱZ)�SĴ�MI��v��kX���L��j�5)�`�R䆭k2,Π����Q�2ɸ��(x�12J22��!/{��ԙ=�udK�d�Y0���0�$��J\�q��q+�y��;̂�SY�E+�bOQ�9�$>�ˋ�V�MPudf%d�Y&�	b�d䎉�-U�֍W�0r+�2�wdo2�'3 3>ѫD���TU�@ �);��ˬws�]���nYh�=�����r�#�dR��<�����}f�c���J~�_Vd����8u��H+و��J��L*��_��ߗO�=��*�o�;q�
�h����*�ӊW�v�fu�NNm%�&L��!�MU�>+Օ�t����Ms\�2������1]�e헕'��5�����MP�3������w��U튊U�{o�(����!���Ǚ��7�o�[:���##��󾪓l\���u5�����u�Jzm�;�x}tcL��v���W�Gc��U���T�>&����(z��te�����
b�zx�5C%Oz{O�����IG7(�{�\�ѹ��%4���nb1e�:lٸjV36r�*,���5�(ۚ�ꪯ���'�����_&�j��w�*�kl�:=���X�8i��4��+�!��<���"��+�S�V�Z8���D���F	��/>_=���}���S���E����;��v�J�=u�]�bkѡr��Or�Y�/}�RV9[�Ue
��7��TK�܄p�;WI�A���&�啄�֧�ﳐ�[�6�{��S�)O�������Gx�&���Aݝ>�����v��k��~z*�F�E�S�:���j5:Pc�+���Y^�ۧ��r��HS��Cؔ��O&��Ym�����KF��ż-RdJI!+˾G��˵q�Ғ(	QY�p�xpڳ�{��O!	�4}_}����z3R�B*�{�}���ԛ�����zu�2�������}F�<������|�o�ZϺ��G}�����̠�y�ݥ{ϱB�����U��+���m	����w���`�E��抺�%��Ϲ���_k����'u���E����>d?zUĮw�7�q�\}�,�Ҷf�G�������W!�ˢ�,ujf�5
0���%��A���ޭ0X̨�y{ 8�?o7��_&/e��yu�mw����U��7UM����՝�f ��o&쭻C��n��/�Ү��Z��Vٔ���r7�l_JVoL9|�)�zf��[h�X:��p~�����$���9[�)�H5��.�O�Y�d��ĉ��ab�)��g�;��'Cv�K�o&\�r�ok��{k�ǦDv��)7�h�L�=yw3�Q�~5ըD��IH֮�⟣:}7�n��RLpU��Z�||�R���ިL=��ڷ�+����-�F��q�b��Y�*q��*���^�
�Ny�x�����^���9�������=�?v���u���U=v;'�����t�^��~7���_Zy���"T.�К��n���WW��h !�1�1��/��C؊p��X4"�!���7F�j�W�LR{��s�x����5t9S�E?���U����zg�Ă�Zˎ�-V5(�a�I��f4Қs[��"�k���
�R�����˽�%3K��=^��iF�6I������P>�Қ�Y��'-z<�f�G)˳6~�i�Uv[7�к�.�ֻ{;�fu��]�o���g���x��k��9z���n�zn=1G[�~��&i��1v�+q.��qт��:�ˎ�-��Xנ��Ie/N�& ���re�2��lM+���gy�x{�׎�t�[b�աԌ�V���3-�����1r7��Gf��o�j���Om�Y}M��d��"E!�+.L{\��QY0ve�%;��p��W��%]L9��t�~���y��|�l����s�wRM��i�k�	F����F����|϶|F�ֆ/��-ʾ�Wc���2'��/������o7�f�N�
}׹���� W9y�O�����Kj��p��&y�B�#�&��$�E�k���O��5��U6���%(7��D׈ZZ|��'�R��~'����h�
{��I�N���\i?�ƿT��!�a1O���4V�������s����/<�r�Sk�������v��ͱR�%�4OR�A.��U�l+$��^bO������8Pgm�^i/�\{��3�/g)��-�/nZ��J�%�������zT�awu�^���c�k�#���s62��)9l2�z���r�~��n@Ef���ǯ��Οt0��sL!8޻��/{��~�v��zE�.H�/��JE��1P�j^�r
��ǜI�7H��x|�pXUD���@��F���-�z�_z�Nb4F�ϧS�s��T�N��ڲ(W?b��=��65p�<��������@"�f��Խso=�t��5�lA]<V��Z'e�Z�
�U[㣳;���d~��XU�dB����ա˃�C�k�R�)���K��^k-F��&�\5�rO�R�f`f�ѪN>N	�+��)٦��N�IrEĉ�F��7r��tc:Q�br�Pw��6�\efo�>DƷ�	��{��_�H�E���DS��<j�Ä&�sB�<����� U�i�Mv4E]��Z�^z�*e�LW�Z�9ڒ�^_{eP��> 鼝<��[1xE�p�f�x?�.�w��Ckƹ��`\ևd�|�d���ޮ�v0���߇�� ��,AL�;5�����{��>&�K���M:�k��x�N�
���eCKyz{"�r��܄�:Jf�04a���0viU~>���5��Ƿ��!��돇Հ��&�W-	��Nb�_yQ͜����f��r��
Հ����vB�O�w�B�>�t��?e�k�(�+7�8>曭�><>�Z,��
���"k�禰�ׯ�	��ͱ��j2}�>��+�^#!NQ�˖���t{D�J����X��%	��T��NRe��}��'�C���R��c��8��I��ˋ/�9VV�t����X�Y�e�'GVh����Uj�e�W�����h�ďi�P��kEO4&w�p*�T�s����R���
�ʬ ���ĸy�@!L:3ţR�ߌV���M�Լ�.���YI�bܻ��+5@;��/���^�@��_AN�v�rG���@�]CG^*�5�kU��H��?G���uy�����6e �[��K���� U����{�������}\l/��./�x�����Ϋ@4L:849y̾��AL1[��h��ηI���\oTϡ��_Mj�����*����
&�E��7j�w�)������o�g�d���/��M�^ ���usY�]�C:7Hmz�緪�wcfHFq��m�ۭ�[��E��* ެ��r���]�I��%�{̣b�I����)��<��
�uî=D��=�t����{X�O5w*a�9�|�-և�h��_�UZ*��>�g#��o)^��5c|th��<*�u|�f��wޑʼXw��T9�%���`\r����}Lz�
�%1]ör,��_���8��*���.�p�.yU���!�yU�0�w���G�v�p�� ���^Ӟ�����H{�&zM˧f|� ���4#Gx�� dԶEP�w��ڠ���y֢G�uj��@ӄ��^'�ܬϯ��F۸�RV(߮]u�x�X��)^#������Q�on�z�xk�D/O��®����v�Ѩ�+�k>]��ܤ�`
�\۵X1�5vO�<V��Ø�#�'w%�pM��m�X�0uvB���v�^.U���s3-=�Wo,,��G��𮾅+�0�»/�]ˍ��H���=�r��c�Ü�\ݐ��Ǖv]]��]���G�9�i�y��H�u�dmk\hͭ�i���(f�kW�W'�0�B��X�V_w7g�Nz:ƫ��͒�o�n-͜OP롸�#WwD�E��5;��������Ci+�bE�ޙ[WS�㍗r6����t���UK�n�b�G�U���WF2�.�g56���O������A���cXU���P��{6�Ы&�ޮf�o3��}�׮5D�7��z�0Y�O���Z�{S��ז�9u/z�T�+n-=!��I�㘞=V�;Pn[|�L0cuh�B��)h_m�Z��]5�ovtpV�g�������t`�h           ��        �vf����+��L���S��X䯧dʏT���]+6t}��Y�oB�.��/w.�.�n���8"]��6�v���.���v�[!����VX�ç$Y�����ǯ�;�t�H�^\�ɤ�t��4�D�]�<΁К������z���y���(��K�>P��� X��&����O&|�}ӎ��6�I��5�v4c*$ee݈o�%e%xB/6��#�j�m5ϧT%	[Ԃ�z]�|��w|h�cw��Epk�+���>��7;{�&�W	|���H**N;�[u�1	|�c�7�E���.]a������t2钮O��J�pʵLa��A����u�yi{��ݕ�"����yj$� Bџ�*���D��P�aC�E��F9&CK�V�Aŭe-Y�yh���͖�3*ɬ�*����Y������α���2���tA�x�MQ�V`P�&k2�n����EU5FBeLIYfv�VM%8��&@ff%SfdA�QfCY�FA�9��q�EE1+��YԜɩ��
b���R�Ȩ�y��QEɒ���AT'S�UI��x�C~�|���H�]�a���5���9���5W	T��5_ #(RHK!���T7��w�� �����b������Y<8\�	O����6el���S1s��+�X~u����@-4U�o��nw�� h}��V4Y�ᇕ9)|	��l�*6V��뙻�zb�h>��u�L�:�VQ[�7��O��F�.�U�����P,�Eh�.���ή¬u���jz�qf���L�KG���HC*<W�Z��K�Z�*K�^���E4{H �^V�Ӡ����_.�U{<�0��9i����ӐnC����Ӓ��\�C�0xW���ؼ3�ߺ���w���Lx�M.8mV&�.���jI�w�'�F����y/��� �?Gx�[�Hh>8Q���BS��/d��/��0���'a�j������"�Ԉ��κ7�2M�&M�xo���IoLw����:�0���/*os{;������~W>�:�VЫ�h8�ʆ��B���3�R�2Wq��s�ʞ�N#m�\s쌺ro.���.�4�׌��n��]
7��j�Vkm���V�D�у2//i^o:<�w�l�=���\|0!c�Q�Q.j_g����d-��}w3�T�˅"i�cb4�W�
6V߷۹��@��yt<�����pTˆ��VV��;ޗ��A�C�p�~>H���Y��b�D�n��V�`g���w��Z=ųU��
r��h�f�]����D��gƐ~-�{y����V/�+`�ee�����(��<Ӥrb~=���������<4�x�[`��U�-Y�%��u�")o_��:.(G���: k/����A�45�|�mI�:��n�X���m�9@K�ƇJQ�0�J��&��i��>�Cq��cF�b�~���@n��neuVL.�kK��%�W�l܉���W����F�2ĺW�����	+x�狅L:r�/�w���3�؞�!�j�y��W�B�
O3�U%���#�M�w�ֈw<+����x��g5ևF�p�Lb`->�v�Hi�Pui��-���h��< �*��5�[��'�� ����nhX*ؚ8~�t_c������h�S�^^D*�D/���th��kE_��9H�W��y=3��M��u�<#�k��S v�'��* �LV���u^q���������*W
U�����.��(|8.�����ﴋ=Xj#^^��p��е��]��:=��zP�����,_]���ᅝ�艹:�����;�ݛ�9e�Q�1�I�}�um��s��#��G�-��3�vJI���a������͉���G#�w�㝦��w�Pʮ.���F�� �a�ǝ3�݁Z�#O������4�**��
�	V�Ɔ ���^�S/׷[yHWeX��t0ͦ��:6��QB�x7]pɽ�V�pxxM�E���!DהX(xA-���]��jy���Q�|=}a%Q.b�R�E]���S�g��ڎݛ(����9�.�v�
7Ք�'c�u�������ܽ���J�Td���=��٨�l�:Z���e]��C�wr�Ez׼v[�Z����)towEu��ĺ\E;��D��y^��Z�n���[�����i�X�ۀ�S	�ȸڙw]$�V�*�f6b�ڳ֪�}n����1���~T��0�5��-جW��(���¦X*��1&�:V�f:���*�7Ir�uᦫ�,��{,�5!�1��U`���<�~�WR��/��O��P��:Rw��z��^7�3���/�ǿ+�0�}���Z�`�*�Q���[��ޗ��7� �A,�TV+�\�f�ūh;����È��W�rff{V�MՅ5V�
���u�?	sE;�S���F}d)�NJ6�>��JU&-P�>�Phu�q�ʇ���_^�_�}յ�d��!T�k��Ӯ3Ɯ��@OT�M���{�)q��#���X�Gf*�8҇�O���ٷ'4JWD�g�ŷ2�a�A�g��T<'Z��ex�.�/�x�)V��y��G����i���U��*Z����M�&=z��J �W�U��˭_U�Ҫ�$ �ڸT�~�xV?Q�%��ZhWo��L$;�����9#�;�¬��۾��!��;�e1ͤ�}Րvc5w���W���&TT�}S����R�ofw{�;T��3�T8����"W�T9��> -4U��뎀>�2�R����W�EG�v�x����^���Aw�0 �q���&pn�>��^�Z��~��~>�����C�+� �+�h+v�bk@ưR�"n=��]���/ۙ*������T4tX  f��k�	��_<A�]t�D�z��u�����Ъ%�+@-��~�)y��ݥQ��
O��><��|+=j����a�5�4�b����\���w���
�w��M�E3�V�/j�:쪘S�c�Yۃbx�_yR��@Z����^
��88?�9p�{�]!�IS�m�+����,Vh��MR1�q]�7|�������- V�Bī1�*]2�j�i�t��V��[3������%oU2ƨ֠�sm��e��2�Z�#�k5�7�Vл4RH�T��!���u�1�ח���z�ƧsWX\V�ΖJ=��"�Z�>�j󻽕D��ȿ�� vqU)v�g�(
�h�^J8��uҺ��-�>��NU�t~
�`��w�oFk��7�ݭ�8w�W�j�xP�i��]��X�:ݥs���褚�ݴ8�0��M?+\U���0쫺'���RB����|Jf�#��QZ��\ɇ��\��l׾'!t�^]{b��`�[ V��<\*jJQ��u��G��<�RyKh�+�9�Wl}�z�^�t.Ф�%D�_��Q?>�t˼��[�8��n����'��hP��S��nn�1V9%\�;�����˃����wD�v(T�����q�Ԩ��@5cY�iQ��0�*�-}�9�@3[�j�[W-�`*V� n��+�=�� �]�~�Ӗ]��pł��'fw�p/���5� ��7�<���ײfN���Bj��uD�U�I�z�?���
���C4~=��ѫ�@R���+���0vg��{=��M�+�F8 D�]��a i��K��T�c�6l>�sw���j�Ml�*â�j�D
w�`d��K�Z=�o0�����4�5¸IE
�6b��Z5 jꮏ�׋|*�A����z���3w��|6e�M�%N|���S1��&sc.f��I�8z��p^2yP
���+@�~�=���ox �㢐� �����W�[5!I�+�hIhRu�go;ٻ�
χ�p������k���&��
�<ڲXsIl[ی�����2{��L�<<>�4T*:'gS�s��~�m��n.�z�Vk.��j�<�Z6��z�j�L7��NK����In"	���{m>��7+���l�2�a�$jz��4�_�w�b:֏]���ɘ�&�vcj�q9w��?���)�y��+E~�o:��F�Z4=�P~
�_Y����;H��U� ���*_ !|r���op�*s~.8ye�?n�7���Y�E�<�Β�T��,WC��K����}����U�57J���0p�� 
����yG%,u�o��߮ҫ�^��ޚ8�
��4��B����:8#�ͣ�7ݸ�04pV��ԯ�j$AH����b�:5n����W�Vp@@ŉ���UX���85�-��HD�{���6	-%X�V����	th
�	sE;�R�mY�rI�o����x��Uw�x����*�zNi�:����D�WL�:�OeT����T���ߝp~5sP _����H�rϊ�z�
:��Νf <g�J��X����R�8�M7%�O���Wl�4�@G�+����6�2R������i���(ڿ]ڻC����J;��0�"�|O�j�"�����i��0[ša����^:�t��q�=���'��{ۻc�Z4�͏��+m1v��yW�r�=��M�"�`�{;��ܐ�z��S'�P�⡬V�a�_NCVLz~�Ou�˽�a��jT����5j�? }|e^*Wˡh�z��E�f5߲6fy�M�ϥ�&��Y��x�Y�t������R�,��H�*ɨ,��a����Z ���;���ۦ4h���4���� �sk*��~{t����$�n��@Y1��j�����3�t�oV�FOD�f&��1���*�s��ȋ���S���_�kM(/�Z�����`����Yz#��O2��\�L޾{dń��W1����5�.,<�s��[�@d:{D�U�
�͛n�\,����F;,$5�[��p�a6+Jru�o�� �O 
�-ɕk��,�Z�#ז��7(���P��qX	�+9��R�m�s��s���z��&�����,k���e��Z`�!�����ەhf96�t�B�gh����]dpjw��N��i�m�@͵�z�i�71�֐��5���}���l��{�m�]����㳺[���E�cip-,�I&S�8Y6i���E,���֢1�� �7 �*sA���<1R�EdPWj��V�f�ooT�5n��Fm�Nk����B���� 1r�o0j��%�盷�iʓ5�;��g@��8gb)��wƠv��P��\�g{?m/=f׋���                      �oڟb��J���L����w�I�ŕ��(�U�9c;��t���uU�jlk)rƎ�F�����^��B�����q�ɯM�U{Ǩ�-��?߹)J���tݲ�f�F������kwk�A��[M�E�6�뗂P�t>Vice�F���he��dfTs0!��D��z,Й|1�;�4���k��/����c�8$d�'Y�0���4��&
U�,�;
��ɽ�[��X��z�<A�����զ_q^�4;1_֍�&)JL(+E؆����í0i�;f�4-��!J댸�7��;Ϋ���P��,t2��r�*�՞w#"pq��֚`�㡏��_��r��v��'� �  ��s3I-PPPURQo ��0�&�݄��U'��Z�g"�����Z8�:�2Z7�DRL>�1q����j��$���q�%LTD�UQDH]�LUD�AMR�Qk0�b"�"�b� ��#"�02��c	s ��&����2�j"j�� �d:�yΰ���"��r��������1""M��ȡWWWWU]���}�I襔��]��ʘ��+��	/\�8k6�q�z1m�ֳٱn_��[��}�s� ��Z/��Z?Z�?��kG�#���	���wP�8X�5zH���-x*�dB�t��7����4i4�����T7D��RU�#:�Rt�S�x��vi�^���c�K@V�wR�v��˴]��1^O%���1V�\}�*]K��hH�`����y:y��}��5� YMs���ۥ��n�EKʃtUN��ũʗ�k@5�O�ࣴ)�gv��	u��/���xP�OC�x�X֌׻Q,����&ٿ ���]�XX���5�^V��V����<����{��C!�CF�8��x0��+<6�ʽv�6�_��;�3��k\��t���7���}X"-�D֮Z'ɬ _��H
[۰2$)�3P=�M�Z�u����*�IQ8a����S��� �V�Zs:b<:a��g�:��]��Sn��`0�<�v됗�>YKN/����u|���#�1'Mn6�����%�� ���t{|��`�>x���U�w[K%��(�Z���X�<����Ɏ�d�}\T:ٌ��.شNI�{�Y���^�Սg�yzN���WY-�W�oߠ�ze=u�0v���P�{h��WDӇyd^���ۃ�T�N��@�ƹ}��a i��x{b�J�ۻ\^^ow�ՏP�vH��k�$)a�K5V":�'G����[��7ݺCX���C^�(YCF�ثt֍@Ʊ�������Fa�I|�\<>Zh����8h�0��GJ�������PW )����#N\p>5+��u<�����U�KEgg��c�[�sW���<M<���5s�5�Y��]9�k<����ٹ���w��s�ַ-Z����,��Ղ���wM6����¤���4p���`a�aU��0/\h���E\��~����8�-�ʙp��a2�H>�@�3�2�V��<e�����+V�L��L�#��?p�B9��8	{��=Y/�ˏ^����#��vz_+��)]B��#��]
^�ZG�p��I����ʂ5R�u5c�th��P?�lq��B�]�oݛ��_��|�D�
U�*C@_��{�h��L53��DӃc�/�J�g�S�JI���Gte���R��x67�6W�Ƚu+�b1Uu���n��1�C��ĈMX��ubG}�5�i�]�ے�Y`�Af�-�

��C�,�|�o/�WLx���o��D��>�T�@�<��+�i�|�`٨���yE��[�K�����޲���Be@Iq�"EZ),1�;Q���3���Ɋw4p��?��L��w�r��>��Y��Ӯ��"�jk�������fV<8U�.����h��;����w!M���M��7Ɛ����p�܉��tI~�7k�Ø���������D�j3E���/+�T&K׾Y&��m��8�5�jZDBι�Ɉͮ��q�y�^��<��`�S:(z*�^> `g٪���yS�|E�1�=1Iמ؆�WDè`�>�
�K���Qv�^h�'ks�S>��<�Ƙ���5����������Ø�om����^��SָR'GϏW
Xs/o�W�%֪C�yC��R_��^LN x�ƕ��<t��5=77#��񋼓^�m.�n)L:����k�NK&�:��ǂ7A�<��V�ѯ`��dt���=O���\���TX[$�w�"Y�yO���O#�S���=N��{�m�s ��L����I>��i��MK��aO���7�����zEm�1	d�Ӡa���rӊ�a\���f�Y�����U,�ãhT,:�]�`��O�a��>q���s,��Vg��K5h����B��hu�|��ľ��.z�� n�赊�k�Ä���4���#�ϕ�w"����|��HU�c�J�*~
��~�ӰtT�Z B���K��L��ׂ�>9Vi J��B�[�T�e����܊��{;r�#��(o��q�$z��4�M]
c!�95�vC��jkՄB�υ�O���&�>�ȫ��Ū���g`bNy{�Givj�E�A�B8p���u�O�ٳ?��4�aS3�jb�:\:̬��:s�y��K��SH*kҚjL�y������H���f���Q����h[��`}c��r.�`����. �r�	nK�k��4D\Ŝ�շW�8v���D}Cb��.?O�3�mL�^?b�|&6~6>�Kٗۻy�Rl_�
� �8�S��+��εX<p���w3}���B��бPp����d,������OyJvsWE�$n���^]�^��i��Kb�(U`4�e�O*��Og{>ne�%׫�;�w�YH�;)xrj�1��
��Y]�j���ɪ6�OŐ=��:�ps�Ubg4�S�ݭ�g6
��ꢕt���Tn�͗$���c��U�0�yK�&ȘS���R����k�5cY�hq�2��>�O����>��������d��V�,����=��$Ҝg���\�RyRׄ��/ ��R���瞶�21Tkx�#��4�á�;�yA���u�\��e&���3��u1Չnݰ��D��+4D���mnO��&`1R�+��������A1�G[Q�w*f]+wI�Kr�W�Xs�G�F60$��C�º�¸=
�7n�Ѣ���;����+�Ga#p�>K�I7�W��%��GC���U�[���T
����I�a����O*g*'4���;ݙ��Z����\��aY��
���m6�Tu��|��KEu�q|tW�p� r?d W��`3ܔ�y�Zd�)K��ۇn�.6�5��0M+��J���u��Ȼ���G��G��ִ;85�B�`�C�Ч��B�G������B��G�W�^�p�ݸ�neu�^Vx�,��~�g����k�Z��S�_h�|rZ�޷��}�v�x GF��I��5�5�SI����E�׬��./���%8Ev��&ũLuvԝ�,-���˥�F���|Fp�b��"�磌9�y�l�~?^�?8��g�y�X��7������1��F����È���Y��HC�,ny m���㽼��V
���p��7��t��lPY���Kw�%�PT=�we�m8=�*D�gEo�د�j$}��p�2��/��P:��RUɭ'���_�vRχ
�DG��y_�v�}݂�A
;��-IV�4�е���.�K���ّ&˞����ߚ���}`搨�u||3�hq�aO���R�ꔅK����T���WuȦ�����<y�����s���@���^: U�iU��V4Yي�Ru�r���oo�C�L:�i��¼��u�툏�Ż�d�U�~�����rɯ��gi�4t��[U(.�\��`�O�䤈񥼕'f�O}{�Y]B�i���*�G����('m�����I{ދt[~�p���߻:Lw��W3j�M���|��Jù3��^u��SִR'FP��CX� �ҬY��Y�4[~�;t|>\%�X���@j�h��,�|p��^�3ۮ�"�sh�^�+ g�c���*g�c+ŷ=#bY�=P+ϮM<��+H7\u���;��.�liES=\}4W����n�*Y��E��� �~�����^y�z����a�j��]qS��ڌ�ҷ�S��O�#�֓bȂc��`P���V?/B8ײׅg�U���dX������
`�w{tm-�/e�,�r��3r*��&�nf�����5���W������V�O��^��=�f+F��*r���8�{et�霢�r�9Hxf���ůd�d����YlY[.�2���m������+�֨w3S��p<G������ŷ<�/�
���C�<�Wx���Ԁ_^�0<)ZU��@�v�7�@#M04���J��+F�u��WC���EKh*3=��ܔ���f��A�P�F	^<i�o'Xn�g�^�Y��Ք�"i7��
L��q���ƥy�T������3��hy�w�N\l�e�E�Q~o��
����P�ȫ�������c�`�b
����W�ꉫ�xt2k��ڷ͒N^s��6�2Ir��+&�I��*�*�W��@v���L��ؓ��q�(ps�N�������l|>��l�-�Do����vK�y.��K�tYH�:��m(���W��>ʔ�Ehp����w�>]��[�8�xQ�4��A��Ux�����(mV��%�B�xX�ܡ-En��ӻ8NL��XrCd��,�\փ(h�Ұ+ˡ����\p���J���Z;=�\�c�S��^d��rq�$Ǩ}o��2Yt�P�;�$�]0Ll�춳S9�]0���j���W���2�"V.+R��Q�7�M�5�^�F���%��9���+N�|��GQc6�Ҝ�!v�S�����w�1��B�IqA,�+:�\�ᛂ*SQ9Ndc������5	�(�� _P������s��!JnCG�l�0�����r��q�,��,u{@�;��|5R��ˬ9M��/Zz�dM%4�L��X���R��!M⇻kP�8;�#ޔ�R���V�^ʙ��`��K}�ܠ�=���7��H4�r�z0+=(��/#��mL�Uyy]�                      �j�t5z����v����e�ĸ�9�@��ڗb�C8�;iۼ!j$Q ,�l�j��W&2R��[�������2�Ulʹ{F�.�QXr�(��F��I�pG2
C���*�M������Y�X�ʠ��Ղ�%��� zY�vmHFb4JO(��5�H������P�~v��'I���L�{+n��-��Z�M�THv�\�w��7��%&�S9��Z��`�K����p����j��L�&z_�wʣ�72��w�xC���;V�b�7d#^5�,p����]]&]8�Ɔ�3�B�������{e�G+fp\BK!�x�T�%7��l��z���
I�C��l	s-aKUD�.�$� �  �zj��J�h���3�(�ʚ"����8�`�����)"9��kVT�LS�a�I��T��c|&sT�C�UU�eSUdf�k�ʊ)%���
������)���Շ3�U4�Q9e�TU%Q�s��dS=YT�DUDTE<g�;�z��.�݃�Lǔ%�U��F�WT{��;������Lk���j֧��Fr��~�υ!��$�Y�cÇ�[�I�p�h�y,v��l(����#W~Dk�kʁ��#C���N��	ߧ�ٞ�W�z=���գL$^'����kn1����ݣ�uN4J�*��$�ԓ���ff��r���nUr�����f�"�ჼZ5�~HV�j���z�R�����ihcG�,�a�T뚹��R��B��X`��3�����n����/�kG��OU���F�7��w{���픈�4E W�B�t�8]q��k��ʞT��3���G�:_P� ~<4+š�)�VjP��z����N�o6y�i��Rt���v��`wR�N�}L]��p�+Թ8�
��v'L7mB���M�f���+�-n�O��ur�}�w��n�sy IԸ�7k��>=�i:f�cslMNȃ��c�\�h�#,�Y�½g�ا[��4��o*P�x,������W
���G���$K5���gZ�Nisxw�l�m�)蘩�T�D��1W�#��x:گc�n
�4����?�Q���b߰����/��u�+����9R��-�h��iy��9�Wގ/�+�Sp�K�yW���n��6�V{��ځ��=���Z%��UKMEX�X%�C&ƭka>���۔K�K8oὔ�;��cX�K0^Q
ڂ�^Jwzy��߱xs��T T�hT7��_:��g_^�po^_w�P�D���j���#����5.IQ;77J�e-��8�;�������F�+��pߍ["���­s瀵ǭm^^JF`hH�3e�g,P��;y=�"�W܊�����Bu*�X��p����WT��w�]��3���Nk�y&ɉ�U��罻u����]V�е���'���3\��25�=���COg*�|<�	���LU7k�z�����_���̮�3�9���B�: U�i�)`Y^�r��	�Ҥ�U.J\����-8T�^�`�j�|��ْ�)o^����aq~���Mz⃷�]i����w�G3�Oq���a߼M�n�MO;z)4�}8�Y�i9u~F7;��{gX�:)���hy�S����mV�{���o&nM�<��"yYT�{��U�tW�T쁞0 ���
s/6o�q0m��<+�kn�_��N͊���ii�.c��_{\�<�bk@����UqkV;ۮ�f�lP�\�#9��m�ـŢ7n��q(�ONn��n�̩t�/D^��L#���dn���٠=���"8����^u,�|0��+(�����v�=�Gw��	�{�e�8;��8k����N�_,��������	��E@�4jv�o��k��U��Z��^�^\a^]K�-]��KE*П����,R��Evg�y��+��u��hZt,�Y��<������t�2`g�V��f�ѯ	o�/��
�� ����\)?+�4ד�{vW
��օ�U�^>
ҥ�
уDīg��	O-�k<�/j��v�q���ɂF<���j��%���'t������v�,���hD�oυ*f�*�l�t���Ƴ��37Թ����Xwt��YU�����	�YQ��O�l�t�ƾ�Hmx`cق� b�W�_�ҭ]W]�8ʻ@���F�Cݍ+B�������lxhg�`�~��T���ywGR%�z\b3ז�ֲ��si^u��4�)Vʛ�m4 q�:vb�w?WۍB�WM��`V~�~�j����	�%��X/��8*S����k�v�+UhUf�Y��xVi�t)l\%
�X�lѝ%��;���i�<Z)�Ţ�}��(r��9
Wg�.�|}�$����Xb�4|�5/�/ظm���V#�f㧕���Z�0qp�bcΉ��v �k&�������hb3��c��(��ꇴ�5�G��;�F�k�U���=�%j�.�%�����u��e�h��Ul�B�"׈�4
N��yŗ��6��gD(b<��8�@��ʬ g:x4�3�fM�f��4�p�$V��{2�wX�V��x��OLwu�o81�ͷ����Y�k���B�eVG݅s�]r�]���QT�t�'$�����!�M�L�|n��R[�uc�J��W9+c	
N]ŚD�nD�F[uB�y]���?Gնp�q�3MAh_�e���y��5MG��妉�>rq�Joo۶�4�h� ���Dѧ�	yVW�=�'�;�{��@wEE_?� ��+5pa�c^*9a��S2(�6��{����î���+����0p3��@�G�w�AԦ]���.�}��v��c�����QUb��w���ӽj�ٙ%���C��G�B���'�k������`��[֯�d٧ck�Q��G�9M�O�lS���c/^K6���+WG���n��1��6ȩf���������~��;Mv� {�׽�T�H�`��NU�,O,�eʗ;E���.4��5Q'��v_M\.�9���:zo���T�݆H��K�*P<��F`o���߱lK��J��GxC��!���iK.5���nƟ	���7�7�*Ⱦ�aS{��w�r-���u1�}R��w��	���E�y�z@��2�Ӂ�쪼Uf8)[�AA��9�÷��nG�u���t��T^<���]�r�֭���%1�޶kcQN���3^�u�庢s�S�uM����]��I��������Y���(棠�|16�p��T��M_d�b��f�{�������
tkÕj��hT4VN��Q�-*͵-x�s�I��llPg������<}Ƽ/���"9��CEM���ƈ��k�ٸ��U�2�N$��S�}�]�h +Nഓ#w1T#˗����L�=Gʞ�px<��P����p�#�jӪ��ns�F�M�2��+j3�Y?p��'FՔ2:��� �᷽�t�ެ�7꽿er=�"���P��
��B��Y�z�u���CIc�i6��x��Zx3;�:�.�Wش�"��
V��Q͹�b�Y%zљ�aӹ]}"��1iVu�{ʔ�̩�P���3'#����)<�__pW���u�:�#��X���T��V!N��r�j�x��M۰<~������u�^�^gEy(�0�6����������˅佮ܰo֭�M<��H7H
��4z3��ߨ��n��@f�z��3�i�`�z�S�����s�������h��H �0�$��{��IV�&lhy��a;S���w�`�V7�+�'B4jc��3L�~�*Fۘ��-g��riR�7=(��p+�>S�)��V�Щk�W����Sč���C=t������a�b�g�,�S�=��Z���I�3pʒ�.G]Q��ur�\�Q�e��R��|��K�n�����!*�q\x[�̬b����uI�/�*� fs���(��Ao�-�a�8����z�\��j��=P�bҬ��r�ȪT7��ɫ+/���ƛ�5�TT���#�OS1e����g����{p_�����W�
+�� �"����u�o�g���@?_��Y��e/Y#Nr�W�
\��I1;JjZ�Ǒ�~9�wC�2��E� ���fY���.ZP�0�>���3��FQ�@.k��0pV`�쁪�e�D���:]��秼�m��;=pM�]�J���$���'2��>�Ò������M>��NV��w�;��m/	�]&<G]k9/���^^a��o������AZ����S�͊�\,��p�:��#1��>Dl��\�A:�:7�P
�.-h��V:�f�9;=9��Z!x}�Oi���db�&��7"�6���C�صj|,.��j��2��Y����\�Uѷh
�r��v� ̦�+_S��з��n���h�rB��G���nNq���
�sjm�6��$�.1���vGy�L��l~��I�9p���
�8�/��
�.a#��}ku3��_w��0�
�k�ӄ��Έ�<2�C�t��Fzg�rǹ�� ��d��TT��+��E8*9C�ʊ�0�d�rl܂�fSxK:%�T>qg��k��Ntׅ�'���W�*�K��؝ʩ[O�߆�k���X�;=K�Y^���R����������e��4᱂�:�;ѹ�gnc�p���}~~W 4py��S�U�С~9���O\����z�����j႖�R�� ����eC�����:���䚒}�=�Sjb�eh�`��wO��f	�߮�g^�w��Oq��
��0FC���X���ݩ�S^͆��h����y1�EF�>CV����Z�)����#*4��9l���W�ı�xJ��l\ۜ{�Ǵ�^��n:�K(�2&�^��Щ�Z
�znu�ʏ6���
�Tf<��֚�F����7�ɴ�E+��-�� y�g���y])�r5$�?N��Պ�&m3il�Z��7s����rI�,K�,h@����א�Ϯ�&w:D�'7������vS�f�F#q��m�9-���񗧲9raX�-��ݵń��;@Bi��ِv�wO4n�d�M۾����k� �<yERb�6�l�����Fslgr<�:cxP�I��<�A۬�:���
h��(r��IWU��CX\�f�g������Of�&Ԥ��G�L��|cd`ܵ�˽�uiѬ"J

&1�[B��,���;�  Ȇv�d��w���N����t�4     �I$              %���_t���.Q��P�qZ�[U�"P
ي�Ǌ��N��7�j-;�wX����ѫ���x/c���tOXj��y�(�Kj�+9�yG���u��'J�6�h0Y��(Lڼ٬�GCv5�����[��8��4�7�bEe����n����j?��Ea4����.�>Rd�!v��SUc�dͱx;��)oWô*8!jj��1[AX2�ND%�ư�M������9*�ux��Z����K&���d��s�c�G�I�ƈ�u!j��Ե�Kڝ�eX={4��)��7��ܾv��l�]���z�
�̻�/���]oK)�z���"��{fQ̼�]�]�x6j
]T�  @~~�AT�G��]A�G[ޓ�Jj��9EfTk2��ʩ���ewe�y�S�eTUUCQ��2***b(�j*�"
&�3=�1��qi�2����*(���f9eCS3MDTQQVa��VFC�9Q��9̪Ս4F`gvUy���a����SQ�d��T�4UHT�Dk�{q)`ܬ]*<����+�A]g�PSGv��ӣ�kJ;e�}A%�{ާ�1|�*����T���8���t�l��/���h�p��U��%��*��l�kw�8�ɽ��^������|&�9W�,h��!"x�s%�k�Wl�<��P?[sY/��l*趝�5���v-�wwiP^�Z�}�ץ��B�3ؐ�5���}P�.��k
���RY�QOG���
�D�0l��G8�*yU����u������[[����]K*�]ܲ�YYSDY���>ʊĸm���u���kE��G#ßشpt�����ቷ[���*`CWޜ�Ү�7�7�*�����֎Z�F�h� h�5��Sg�3ɦ��gT��S��L�j�6]��H��1x7�`J��֍mK� U��t��I���rl��Iれ9�ʺ�O�5��q�۔QW��"����r��˙K6�\'N-)˕��nG��s�Ղ�=��ֱי�_��)��I�A�Z?�&�f�D��9��}�=�܉g�j��NJU�i�& ۈ;K�`���2i7��G���^{S�ٳOL�<~���P���VP�X�c}���Sޑ�n�
�Yk�s=��yK^o�&��
d�*x�qm���9������|3up��x>�~ h�����^�&��I�t��3?i^�̍t�Ͻ��4W�^ �X@qzv�N���8(xz�/�p2��/�٭u���a���?P{}��iX�^�}��������c: �5�aѯ��LT�I��5�v<^���*�> O�F��H�x��1�l���Sѯ-�����&��:��	�|ǅh@�S/��G����{ޤ�xV\��IG9.�Kl�Rڕ�5u��3�z%]���� ��䳗����i��{�|�76̗dn�nvr��eo�ie�����I<��~p쾭��
�����n���
ʗ��=���M����F��x�:�>ӡf�Y����V��k���{�n��T�e��ԍ]x�({Mw���ܻi�~/��?$�/n�u� o�B��"`x��<.�� V��:�c˩D�/I�G���c��n{*1//4K���ق�Sʾݣ�X�-4g��/́嚝<��^�=R4�
B�ex�_Åԏf���7;7V�="�G�C�>�#�͓�{��yp�cG����o�T��h��@*ָl0p�����F�|5^��==�ͻ��i�TU���0�:>ѣ��z�}����[i�b��}5���t�l�[JLE�/	�]&<G��H�#��<�J��n��x��ʜ5�ڊ��^�=ӟhvK�˫�j�黼�5$��J�W�(uj�r��˽�nf�0�B����&SG��{��<����?P9W�1ޡ����+�1M;(�]��dNJ|�`Ë���	�Y�p�z�xxl:;5z���u���K�
菓�w��A$ǢI�n.�6�����9���bOg<��1�9R���p�쫨���H�\M+�LW����?~��¿g�]�'t�8���ǔt+�9���Y���&y�G����J�ʴVs@Rd�{Ν#�xFT�nxt�n�j��32�}.����9cG�Ѩ�*�F�R�j�cDyL��ƹ���R�Fa7�rI3��C�s�S++��IOL=�%�nYPM�0,���w�_F����Wv�����۪������ �@X� VY����7}=z�]3�����mt���ʖi]��X�twB���tm�i8o;�)�jb�+E읲����\�V�#���EW�Re����m��e�5��PP�����v�Z�<���[m
%�/�#�Q��g��(a�S�xtW^�H+������0p3�����{�������5�k�;L?���`�{X�����	y,�E?- Õ� ��i��_��Q�L����75! ��ϰt��w�]AYz/
g-և�*���8Д`���xNʙ���G\�sy4�S�d���@�����+��+e�X+�״��㷌�%S2򸭯nB�����*���t(LW��_�߮C���<�M�{g��ap�=����4�]i��X���7}�	�thG���IR��1��U��%[�
v��Oy��Jm�ݕ�H�M�<0����-���xWC������F�7[<MX�e��|�ީ[ע�6���7"rBc'1)�o��$f�ݫ�X��E��]Ջa_�U`.N59�S���[���O�ֲ�x�(��Æ�m��xA�<k��Pm���C�xv+.���v7�����X���> ���>mݑ�s�~�&����B��)��v~�t������Yb��jFh��2�Zu.���'
�L�s�]���u!ݦͷ���;��Px1V�pj*�|i�$ࡵh^: XF�Ɲ�)$���n�s%��*Ш�S�W���e�Z
�¸�t	���=X�X���3��`�F�8�y|�x!Qˊ�������}��A����H\�s�k8�W�\(�d���p%$Ҟe���;lK�T:�/�^Vh����5��'ͺhS�f��>>En֙��1^a�x��0���xv3g�?>!�ܼ�ql����F����莚9馎69�a���^��ȹ%�����lVU�g��s*ݔK��Nڧ�WS
c��7��n���rL������d�HMl��[P�=�
�P7]V3���Q�P�`˸0m�X΀'�V�U�u�d��j�u㹾i&��+�螛��sqT��.UJ����z��*�6��~~|�_��ګ�+��Z �f�L��hq�<~(<�����b��^�;χ�p+�R���V��/��=؎��)�w�ި�!�V�.�Ӿ�hx([�i<�� ���D*Ky=��)���W2!_J'����,��W-T�w��=ܣ�{7��]�8:)Z\
�t�i���x[	R� V�	� a�3{پ��M8�&�tz��Oe��P�ă������5�MNK��9���Z*㲫*�z)=�>��ЫŲ>�e��=U�	�6�sy������e]_g>)c���1��dYt�t����y�6B�inl���[up"J��ySl̰lDzPѮ��Rg��p���"��WW��ؿ�WF���љt��,��Õӣ�.��֞�W1�U8ׅJ�@-k��8A����x�D���kty�zs+��^qV��SNp�;/�o;ݬ��h`0ч�{�������:�T�������\{K��	qu�N�*V��p�1h����(�����t\�^�����?����GUgF�Rz�Ol��sݛ��i�0{�5{�Vs]huF®>�\	5�rB�H���=�Y,`��o'ʖ��k��.:fTJ���<�����=Ѭ��(�oH��حRވ�ڵU����Fv8���{SeK�˾��s͛��*�!�"���ͷ���|����9ޣ^^��ą��2��B���'hk4�Q�#Iȉ6%�1��y��<S��}4�/]�.o7��1�&5��d������_N�ҍ�%�z�����0�fa� �u��w����G^�XסG�z=��K�ī�yc�m�����n^[�:�w���}�{.��rS4�H#��{����#]���1�ç7Խ}"�JsS�/��GcZT~��쇨q�Gn�j��b��][k�R<�F�B���,ggtJ���Kw(���X�r�^��Y���O�A2R9��/2���|q���?I��=�!Y9g��k�g��l-f�����$ǰ��4wY��E�����[�u��:a�7�l���H_ rڥ����5�^�jɃq>���e�=[̈�ň�]�l?�.�o����%���jM���D�7"ry�հV�{��Y�᳻mvU���ڋܡ�f^�'V'y<�[^+yjy��M_j�7���c���S�=���['��8\�:�O�OO}��ߢS�Qk���X��*��b�B�P�����<�_���Wި<��,��k	W.��={k�J���yݪ~�{'�ʂbq���\�K7�>�+p��$�*m>Az���u���u��q��q\���.jg:1s.L�f���Ǯ�skѮ&ң�=���s��z� ��6��|cO]J历;���,����Aܘ���}R�Z0�f.]܌�vř��P���c��#�u��1m�;z[��b��(��>�}�k{Y�5PN=n�Q�}� ]|]`wI%�_���
h.K+�A�3�;��ܨ)Q҅��y�W�	������,�Oi��:�V&�\Yyh�9@˷Y1�#�Va��.Ggڇ{t�e.I.����΂��X66�&mH;WK�"�>�w%�r��:�-Y��y�d{,�&V�qM6��{���fK��U�Ō�L��^c`�3s���3�f�Hx+�𨚈h�������VP��2�'|g������Jp��+�sjX�&B�-Fv��I(3�G�o'n�u��`�N�5s�s�yx@o9 @��������_�                      �ۖ
gn�Kd�����fVZ'�ɄS�]��S��H�������=V����^.�S�k�Ȟ��K-j��Zh�V��]B�.��We���ÁV<{�u�n��ז���::�
�*DD��Kp,�/e�/k~V��W$�3[u�/w]�s�=b�_:����Vצ�M� 7v#cʜn�iKN̢�ٝM�ʈ������A�*�v�v�!B(Q#a�m4"�������/�pXYI��֟�s��	+8v��$�n�v �Ph8�Zr��憇g_3"�{wΞ������j̰�8��>�w�Em�˸��W�[Nݙ��FD7p͝P��)ڗC��o�IZJi�0����:&��UB��[���	�����bb&Hb|�H��k���
�ʢ`��5���FYAË́�A3V��Q-�.YQT�deTOX!C@ЕF�(��a���
��a5TXb�	TEESC՛̚J(*�*R���(j��
��)(�k#%�ɪ����:�
*��ɂ(*��&9̨*���0���ˉȊ*�h����7��P�*�H��xۻG���Z�NYZf��yt��z�{K�q�oO��Yɷܫ\�~��p�zy���=��\v?z/;��ȷ�|�i>���E^z<�F�b33LgD��[td��b����/"�c��ګ���{k�<��`��Fg�Hi�d'�7�/U�o9����j~/L�����RO_��M��{�OA�sF�j�ow��jO���ovLJD
gv��c���q�yI��m���m�"g��<�\9���8���S�˲<g2�_+�{�遠[��x�o����]��K��v?o���Ip�T�f�D�m�v����A3�1�[9}��[���J��{���|/�ym� ���2�"���O�	�ߙ������N�1M^b�9N�y{�y�P�z״A��T%;q"��Q�(��g�4�^����ߓ�����}��ו�Sخ�b�W3!�ˡ�?f7^�M0r�0��.�fA�R7#,5���A���h�m��a��F/zp�T]���n�އBb�Э]^E�UͭC-Vz��it�s���;�nW��߽�3��ƅ[�α���(8�D�Q�رq��[�aը�����y=2$[�k�zs��b
=k?Vg�u�7���Խ,�{61wxt$���`�˙�EAw��Karط4G�&;Q���;���q����ѕ�:���8\�FJy]�;Jtݱ�J�OO��q���>��=��Z�ߋ9{b)NfQ����'�ߒ��y�2�,�\r$����%�G{��q��x�A���~sP����͟Wؼ�V�%�<w 揽+w�X��R�d��o�tf��s:�#��6څ��ɡ�Z�p�5o+%^N4��5+VĂ/�iR���ڞ>�s��H����C�F�ӜS�)0�9k�{l�f{����կ]*:ߔ{�!5��;� �Ӄ�
�z)��^>�dw��Qh4�<6n���+qvY:���ޫ1XӅ(0^���� �����
#S �.���^�vS�n���]%�Z��\5������ͷ�5t~��o�_�<u��'��i�n����.ΒA��C�Ȏzp���|�X���k�:;��7���N.~=չ8�|��k�8�7��P��G��ό��:*���$�/÷W�Nx�燽��z]���0փ������������8��J{�Ʊ�a�c�#�S�{����R��ߥ�E�WHw��Z\�����z=Dm�z��j�����Oѽ"�x��)��IF��Io�2y�G�(1�y�o��~�����'�x㋃g�nb����в&*x�(�M�m���[d�+]부��9��Uˮ�T޳Ө�%݀�
ިL�WCzq���IX���".��SW�Q��?zZ�E�!t�l[.�=|� M��۬��qв7�QЕ�=���q��5�p�j��>��l��v�Z�벉{�OPu��ͽ]5b������z���4���mJ�]�9fz9��5��e�M	y,���A��9vu!�3/�c��oD�w�B^S��y��]�����м&a�s�&��U�y.��´��;|��tȀ:vy9
U��̲#��*[�<���v��眔~�^�ug��AIN���L��tb]�΀�c�t�}&����}�*�x=�V���Ӱ�� I�X=���:V�r�lX3$���(��m;i��u�h��C�}��s����(z�-eU�sn;��u:������7�qB��pr�Oo��7�Pگ9��q���e���t������؝�aA�i���C� �cЖf�rl-�留r�o3<�T��9xnZ��'P�*5�Bu赍(��T>i��L[�S9���5��gH���q�8}9^���}yg*[g*̊F<�f�^��:L�����v���Qz-;�:E`IT=��z��(��j�}���=:~�D\˹*ǅ� $@8��i(�F
ۡu3@ah����+��D�{:���:���_VĴΧ�Z-r�y��Yغs���w6��ȟ�u����~}�)ߗOj����x!�6{�+�g�EPx�g��$}˹��.��W��*�>�M_	+C��`�1�g ��K%���[���'�+K'�~[α��nrh�8h�vc|,�^�o��s餧O�,�Y�(����[t�U'�k^�cymc��ed~^��A�)~u1�r��b�#��NEu�͇`���n=�iފV�{x[�^_%��ny����C�>���W��Uc��~����X��w�If"�<�kZs(��m������I�FN�=RԄ�6L���
:������10�͖�����'?U`��<����?��9�T�f�6���s�����^��H��{���)0�ώ�9��F86ͿIC�0f/d�EV��E:�xT<6��߻vK��G\n^Z�ZTt��)����%c��fT���OiQ/�b���׻pڼ�5W{.9��Y�=�:�w����^������v
���~���8'�2��u��_��v�wEf��~n8���nW����osi���ݳ�tެ燱g{��v�p\K��`��ڋ�m�q�Vz�d���#��F��D�$�գ�8���+� �� |\�U��-�gg)���f��P�s�ϐE%Ǫ��7Rl����<(Q
�k�xU/���xߞO�������uo'翿4�ƞ���Q�*��}�c�Nzs���qM��x��X��`�)]2G�d��H��n��N}��!���-*�z"�h˃$����Y�����Rsh��W,`�!ǽ*�s���ο�
����Mr	��~���J�y�{L^���w{�w������i5*����*j�O�����i�;�$��F�n��[{�z��z� ¹ȷ��K��'\��uS3pZ������f�{��t�U�k�@�7��Z6�
\aS�f�&�*�-䜢�Z'��������:�m��Jq8�Q^qc��ݝ�=_��\��{R��]�gqW~:�34�uNrca����mx�tf����|��N�<�8>yj�g�%Z_���R]�}z��:}7�i�.��{�W�X�������<�ۃo�͍]s"3�d�o�u�����r�59|�zFr���V������v�-�$~�/vZKk�{�&�����!�^�ޡLb�}���c8.�P��j}(�sQyX��z���X�n>��ޞ����Ɣf�%�#�����VT��w�X��=�ȴt�+���
u���#X�|�˹�Cjdt��X���Ly��LW�J�hN��
�{>�%Oh�PW#����mX�(��oP���N^���[�`����d�c��"ޤ�E{{��y�U�j��e!�{��=��9��\w\���.V�%�r��.�ز��_Мwl��󙰈�V4G˴�q�:�$���4��e*bzh
V�טwt� �u�]nt�R}|�>�B�(����e:\pPf�&��tvk��S;�4���뺺�S�M$P�+�C�e+0�gF�\(�ݻn]!�'<��uu�Oe�

YN,�'p����ӚvMt��SZx�A)1+ŶƘYۻ�m���$�o��;7<_ag��5�ؗ�G�F!V:vn�d���祥����Fr-jU�>��� 8                      +W��ȝ�*m ˂���m��GW�Q">��%�q�P�+\�p"��5�6`$�ٍ��<���hJ��5��j�	�ĩ� :�J�Mx'P�X-PᖶL�i5՝6�V��|+_{�3y�E��>���\�c����v�kM5����yƇNh0���#uT�v'�l��-<�`^�;Y�%\ꕨ�hdx�ٻ0.����Z����[w�E�+�+td�ғk]Z�,�UY�IcK��0n�s��*��e;α�)�@᜝Y�wjkUțP��u�׍�e�O#�.	��;#̒�B�s74K��T��GǠ�7���#	|3[�V
�@�"����f*�.轾�DʯM/h$4�~o����6h)"�Wj*���(�&���q��"(�)��+y�PE%n�*����2(�f��*���ݢ$�%�9̊I��2�j�()��"
���"j���7�(�)
j�;̐�"�������"��JJh����1�%1M�SAM!UݒU�Pu	��¢�bR��*���������;�)$$�m�<�Z��I�Od���\�*�jM����m�G�}���yث�����.����iX�఻������`��Wem�Dڕ�|Z�Ƽ�o�Q��p���>���΂e5��6Fe?�M9�=~ɦ��}QP�Y]��=j�5�ζ�]�Y�yv�w��u]0�j�u�%�fx��n���r7'Q��{�4�nq�	q��Y�5\3�V�Txdz���)��wI'3�kIW�N��^^*q^p���F{�|�,��F#r5m�N{�ȕ�]�4�U|�n#s��k<줛�:��e��<��.�~ګ	���-X�w��n)׮�/L{��^ƺ<<M� ��V822"Og*�Nu��o����~�<�É�4|���z?�]D}h��w��潽y�c��-x;Ą���B{��D����٩��H��.{k�r�ƭJީ!L{���I����^��M�z1#�
��ܢ�T9�<����V�߇cT]�%w�bI5"���nj��BJ���I��o�&��˛�y���Ҕ�z�+$�����;'3]]�߱GF%��ؽ&g��0A����F��2 ��uv��%�^%����H\�\��8��\&������5Ъ���ښq��5��֍8/}�N#��ـ����͑fv���}`��,�]�;�객��ŝ��y���<^c~����Ʈfˆ�oU
*�<�j�j+�
�ݑ�.Rf�%/�NYzU��[5xi�������ݞ�	�#�����Ǯ���¶W��y�!8޸.���+�k�/W�ΥYWQ�B��N���U���8�dZ���JJ��`�`.�q�]*Sm
����{N!^����
�,����}h]s��x�����΃����e"�_�F�u������ZG{�w��-�o>���7%c^�����
c���e�fp���ȝ�'M�=�k{�	��>����.��̯Q=�����k-.�VXB'��Y�(8��`��%��s%zםg�Nk�U�{�~=�+�2��0[e��m�_[[	v �оƄ޹m6��[�����b,��^��l�wn�x���0������ӷ�h�}c2��Zi��뜻7��VK��x�-�Z��ָ�z�������o�?n~���Ac[Z�wu,�$�v琿2�Ϋ}r�[�s^;x32�ʷ�w����_��[r���9J+�h2lRӐ�i��{�!��pG�aU����/����mv���iuvٗ�V�߰*Y���a�~]!�>G�K_ds,S�^y�^����������5����}0fĹWj-��4�sH�rvo8�uћ��U�]�i@�(>��3��Ɉ��8ےD�@���1�������]M:����'ʘ�i<�bt�VvOG<���L�+s�� ٦s+7�u�ޤ̗���;取k͛��W��G��g%r�w�A��ɮ���o�f�k�C��/���t~�.�|��M
�*�8;���;Q�$��fU�R�O� ��WTܮ}��ݿO��*��V5
cj�xLB�ygCg���ݶ��㫓"�Mxj9n�Nі�C�3��cg��+����wC���c�@UxG���h����п|��!U���x.�쬠=iw���3U�(~�^�eo�s����UG��5%m�!c]��T�U;4�oiop�S�.�v-�^�p����I�f����܉v���{˷�<��"��:��K�a��?y�l�~eN��ʷ(~�m��m;�+9��o����~��5��y���i���V�N�<�v�B��N��ۜ�Y�B6���V==��ֶ�D��o��8��Pk\��2W�!�u'>/�a�:[[Uu��+��=��.%����%����d]R�}��(1Y�hytO��^�R�&�����.]^�ٔ�Ƣ��膤ͨ�e�o�TÐ�T���cΥC[�EEf]T�8��g�(7�ZS������證/BGu�[49A�{iv�!z]$���s2H���Rŷ��L;�0�D-	����nՎZ��Zj�&5��N������<ŭ�h�xR���je
{�`��.z�{��~�M��1W�~Xw7u�L!�]�mJ�ؼ�=��v���L�z�����y^k��w�2y��Z�4D��S�9�63Y�M;��L��Kz<�6�~��
C�n��ř7||��e��w}��v�43\te|�����t�xoV�﯎�˘��|�g}'Gh��R,J��V>%��r^�3l���Z��<ü����G�;��s.>�� 9��_s����V%��P�9���Fw��6z��#]w�y��]@�=��h��%�3I)(�V\LX���܋H)h�9��5�v���}s9ɘA����&\�a�V����\o�;���䧼۳��KY��Z���YoKyj�1N��-��_�m���f}�[�H���<ށ�$����j+��$]m�_C����Jb��w%����>�Y��U�mM^�~��j��C�~�U���ѕaG�5a���{��a�`��t���°��΢���[����nGcc�=�!�����X����|_��V��.���T:����u��Y�Iߦz�X� �m�藠�,�&?=���N�]��͖#}Y�H���!�6���ˎy�C���&N;Q��\�kӛ}YI%w�ˮ�\�<�\v�0���4.p$iِ<i'�]�{ϸ������H`�j1�iT�n���w�M�ϙn{Lӆ�v��`ZOq�Ygxc�n9��������ϑ������o��-�OG� 녿c�y�ԡq�9+)Fy>.z�P�/VbT7��ٍn��M{�h0��m=R��s���^lߧ��,��T�yl�]k��q�H�>������96%QG��|��z{e:��X�޷�������~~��p�/GwT���z4��2�yO��t������F�e�W�Nm%}���_���đ��^l�y��l�ok��r�	�>T���$�x�.12������yR��x��0q�����!��^䟽(u��`�=�6P.�O:O+'�s����dpfӇ����� ���>�V�ޅ�^<"�'��>�^�J���*��`�t[��{;y7����n���o��D�j(O���~i.��/5V].yJ�z��^���ᾭ�͏7��b{ZJ�zv^���z5\yLU���xW��~^���N�{�Tkcl[��!;��,y�V�4�P��0�=�n�+��G�J�r^�9�y�˙�_S�D��(�z�M�?w~u�|o���A�'�~����Y�UA�V�^���D��<�Qd�$D!����*)S#�,��b�ey|�-VV����kS]4��D��X��*(%UQ��\k�x�=������u��~,w	�������:r�1C��1s�_Jo��x�*�VtM+��n:eі�����\��hz,�/2�',^r%�cSfY�e�<���]��ɔ���׿�LѠ������PA�F����~��4��$���b!Щ3$�~H�i.�_��捫��O�"{���m�_�x�~Ӝ��7�gg�H�CQ����Iڤ�(l�E��j�]$b�z�����,����1Eh�z�W��~a�r�I(�:7��Q����wbSiw�I�1Z$D!L۱Zi)1�{]�/_6)L	a��w
��P��:09��3B�<ޚ�`���b~�^����2&JUUIgG|8.�I��|�-zT����D��=�f��M��~��/q��ϱ៑���wjT�H�1�KISE��󑹓��;yã�vL�w�t��c"<����˗luʬS|���;�C��_l��e�vy<��ޢDB�RQZ�yu%x�L6feԧ�,4��z�eKZFRBBR�$D!������1{��iUdp\a�ږ6��W���1bF�!�FMׅQ:��mD�C�t_���ũ7J��$!h�1ZLS1I\���a�^�^�jK
%f���a4�]8��!�9�x�<�t|�`}L�DB��S���lH�#���`W��'�RIG	��R����O�����zkc�:�.H��8ɵ����U(��;	հ���{cډ�#��lj�>��bDB.s�;�+�J�$Z� ����+�H�B�{q2�+T��=!�48�9�u�B6�]����6CR��x����)E�z��ܡ���s�Ѷ����kQ��zj������g;���"�_Z9#(ö3��*�vc��5=�Sq�����UGME�mY�^Vᩊ0�ǵ1H��蔄�C�%I<�瘸��(��^s���4�v�BD!�'K�p�L�i�vvY21�VC�!�z�ZC���N�����"G�,��cj&�9��ܑN$:4��