BZh91AY&SY�Jm�J߀@qg���c� ����b@}@    <=
$@(P�� �U P*
PPH �   	  @P��@ �� (JQOF�UTUHJT��HBEQT�UBR�
$J�JUU*�T��)Q*���JJ�E
EP��T�%J�D  �2U��EH�B�)B�A$�T��!D��!P��T�)JPJHIP��(�R�E%I��T��)
�&��IE%U�  �=D��hH��Y ��� VQ �"ؖ�
X�֒ b���hP��I�R��J���UIJ�IQU�  �� `3m�U4I�[h MF  ��l����
b�@ 4�sJP�h��4 ��h �ꞷE *�	R���O   M�J�� 4�'pt ��P �S� �\�p  �s� �J�GB�2�: 
Q���h@v8�T�T��%*$*�R� �8i@E��A��� `�h((b����`ʀ�K� ,� h -L �U`
 P���I$� �@-J *ڠ�-FP��,J ZV � ($� � 6�h �� �����T�& 9@�љ5�VQmP�e`� j`
�Mh����  f� h MU��������"�$T��B���T� �  eB� l�4$�`P ʱA���  �
�a�PҰ 4l�  w8�U*A�*�E� 6p����@��� �j Pc(� j�  Z $f�  � P-E	P�	@R�G   6�  �0P �� # ���
4*�i�D 
YS (�j2���*)B��HR�T��V  �� f(��,  �S 
$� �� b�S��͘ 3K x    �AB�S eIT�  �  �{A�RJ�L� �  ���i3#I��OSM!�� 3Dz���D��*`�  �&0a0�` 2i�a	Jԥ*2��0C��L d�@��q��tK-�������]\�u�Y�M��m[��ҭ�)|]Y�}]��l@^J��� @U��B� ���2�Oy��O�����S�Q `<�U}��� *�a?�t%O� ZX���8����N�&�'&?����`O���L	��D�L��T�
u�zʝe�'YS���D�	�dN��Y���� ��z�=dO���z��`^��Y���T�*u�:��:�=`^�/�A���:½aO�e�YG�����a�XS��:�=`^�X���A� �`��� ��:dN�'YC���@����	��"u�:ȝdN�'YS���'Y����	0�e��Y������D�u�<�XG�)��	��*u�:��dN�'XC�u�:��ex���(u�:��e�'YS�
u�:��=eN��Y���T�
u�>�'XI��
u�z½e�Y�#�W�u�z�<a��X�#�Q�(����=e^�/YW�yaN��Y3 u�:xex�(�~���ePs
+����Y�(=az���Q� �@S��XP0 =eEzȈ������"�XA��|`U� ��@�(�XUN� =ePz� ���#�US�(��� �U���eP|�">Y,(/�AG��X�)�G�"�YN��XS����
}eN�'\�N��X����
u�:�=`O�)�Ve� ��:��eN��X����"u�:�
u�ze�'Y�	�D�"u�:��n������φA�=����[_�ڶJ�'����N��V��T;#�5�rvS���ښף;-��{5v���Ԓ%���vdGS��ݹ��a�Px)ք�Q/]�K�]n�V�=��ϫ,�9N�K�M��S����gA�E*nv����)9���9D��ˋ/1G���;�Q����{�ֶ]'8w(y�ɗj�rm{'&��f���-���]%I��gh
d�r�띚r�Vm�ܓ�+Ӏ�?<� d��/�/�X!_^�c��KkD�3_+�pq�Ͷ�asJ��>3g��t�d#�N|2ۖ��=p*�7�E�@��ˎ�ۻ�Mt��2jsZ��tq�������5��)���DLptۄm]�nm�଺ù�����=�(�.���5�ow��H_wg"N0�����R�����E,��
�yغ�w�vf|ju�K���]&��ɝ���$CM� Y8���[��.�\{C��-Ӵ�,��V(
ưh�TJ�i��XV����j�<H�8�x�/}��:�ΧI����;���)U��j��m�5�)OJ��	{y�Ւ�kԊʍZCY���4�x��ac��k�V�{���8��i]����͝��*����ƱJF ��;uN�\]��Iz��S��]��vv<x��l�B�wx#�.��᫗H��9;*��f�9�����[d:�{�ٻG{��$a�Cyi����uu��4��Yhu��O��{�sX��p�7D#�KUR�.�	�f��g�M�{��wYk�
����hȝ��8#A@AP���Lo����Y��0I�>Z�HY�r�l��՝x;l����/�G���^ܒ>Y(\ڬθcs�.�Yy�J�E#���Q`����&1k��I
�7��(ֆ\*ԉ[�*�f.�2o��ck��*�ڭ�N���:�[k0�����Ű�Z8��Z�f�v�x�U��[�#h]"m򦡦n�&���UY���kMp��f��7H�܆@i��z�HN��K�EyN^-�y|��$�J[�����7��QN%��7 ���F�t�52�sz�+������W8 uj�s��kN��쇆����Ѽ䵴��6��c�;�S��9cI�d=V�U �p�wjH��n��DˑP��>goeT*���3�eX@�o�F�����l�^�`�w*�cpN\�4m��ޣ����t�@e��������T���(њ�U�T#i@ƻ�bv�]A��'D8���A��z2%�;�,e�f�<J���Sw�6l@�-k彇�V�M�c7��׶-g0�Z[��t�=x��E=c1�|�U��Ej�U5����-�S	ͨa%��4�OVr�MP������C��HQ�6��-�7By��4�j�_lE�`�i�Bn霕��9��R"MC�Y��;�D�[�M��n��܇�!��sr��b�2b��F-���?����/�4ul�"}Q��6��u��v-��4����z��wj�6^���a�K;���z�M]�65ʷ�݁�K���X������h��f�,M@�jvpД��(=N�K}<}���
8f�r���i2|�55�hM�F�a*�s�ˋ��q^B�s{�z
v�e1�hYc�����d;��#�u�V�ǂ܌�o����=S�r��c�;����q>�So(as'��j���rf�ϗLӣU��V%�^>e��f�4�����%{f��{���Ds�X�/:�x^.C�u�ڼ:��ҵ�ǇV��]Tk'L�wk@�x�:w7�'��	��>[İ �Q�v�ϵ����:%
<��QǃP�^�����t�0\�=WK,iI{y��T��լ]u�_�٦��d-c��V��;Uu��gn+�.�9��I�l�N	�ʫ�.���P�n��A�uR&:���o0sZ�VK���e�޽�3^-M*4N7�ݻ���y%������H>jCЫv�w{	Żl�v3�������5؛>��Þ1�xe���n�����E���9]˲��8�1n5��4<�%P]�;��N�k�F^p,o���O���w97�Qۮ�����B�cS������Z7��]��m�"�x�.�g\� spA�`��b��9�tX�
�֎�ۅ���=�y��ǹ���&�a#ȡx���8A~G8��zT�4(�ݸ�ej�:	�j@�ӆ�&�H�0�$ig5Vi�Ӈ!�����ޫ��1���Z�uG�U$�%Č��͹&�o+9f�V]z�CE�v�Q8�m�V�[���C00�J���m�n�ёe��)Ի_v�gwFk'H���8�au�Q�j.K��w��B�p3��>y.�ŉM�CۍQ^ì�ֲ���T����8�"�u���D�])�ި����y�ݮ�2�u[������$i5��]TCW[9�u�oi�y�
���,OU�%J%���0q��㻌r��cx�w
w��k����Z5���5�{�L珏�<ؗ,�cV �u�ژn�	��`��t�����H7�m P�����D���]8�ϋ����vBp�ȹ���L\���=���t��p��;������k��4��d�M>(<�).Xhn�wnŸv���ңׅ�d�R&ϫ?1��SJV;�5��ˆn4�E�0�bݩ�����^驎&Y:�qt<�j�"�ã	��1�@�_:�n��xS#����+��s������&��4�i�*���b�ػ�궒�I!�Ň��֞t����Ő/(�1��bh9��ΊY�Ijp�l��{�D=�G^l����zI��<x(u�%�����yZ�L_rw5ʝ�&�w�m�F�+#�!S9�,�^L��J���Y�"<����D���U�կrvᛷ-�6��W'|q��hm��I�K�����7N>�[�e�
k���E6q/�{d@�t�����+�4�4���U��I�I0��=�3�^]r���tӽw��vv	����R
R�[�sKN��%e��coG5����}Fv��!��A���Ou��H�AYY��j�Xv��Py�n;]���]�]
�iл�ۦ2�zwE��3�f�̻�v��C1�9*�-��^��(���К��XQ��ս�R��ڴM�\� ]���5Gi�z�-X��W�3�.Ih��SZ�LF[CQ�B��2@a�7���k�Vѯt�>�(I�ε$�1<�>�t��ߡ�5e��
��ʟ5c��=��$�U�v��;5�2UƱկX�p ����N�Ճ�N9TZS�E9>紡��X��'��i����ΫxXN��K3�%�����^�ߔ���C�S����T�u��w{*N)�$��jTq��`�n��a<P�_>��/-����0��Kݻ��Gh3�����ђ��;w��Ď�@/���Ji��7nvWG��`"�Ôl	�YyV7B[{��Iݍ=���� �&9����X%(]/�oN�����vmB�Ƴ�wa�42�Q�l��oF�ߝ:P��9�������{eb���o" ��Ӟ���;,L�薨��vv:��-�1�7�96fM�Txn-�-6QfjZa����S��̎���5�]0��[�}�8��e$�����G{I�>�;69vX���m8G�k˽k:�n��2��&� ���+�����Zm'hڦ7�&�����x�=J�^P=�^v����7�w9u���]%h���-�L|2f�عךdTqMh<z�]���2��v�VU�rXk�<�Ց]��y����ܬ�l!�%l7u��6��Ay��:�>7D�j�8(�4&42n!,0<��dj�n��n
�M;�f�)-[n���No���a\�ˎ��7&��u�J�-c�!nQ֝�摷�V׺�SL0"�#�X&&����	-y��C��7R5j�d�V-ݖh����u`<�:�������5�6�珱���r,4�u]e��^\��1��2����r�*!���R��Hܒ�>�7�ѥ��짓D��k1ا5ݳ��a��[jW��%�.��#�����'��5�=����7N�:е
{�ݜ��vq�nލ�9��p9pC���n���r��sQ���0�z����W/?�p��B�X�6�0�H�u�vb�_��:�$�4/� ��	yy������_�,o:`�[�K�w��H!K5��m3h�r�E�rOLy�P�,<K`�4�[�GK�)�s�Y�,���4N���q�8�[Äx�8*���u�lY5�2{�:&������p�F��!��vk����|G8����I���#0��X]7(�g�/;�������<k�' �)�h�땠���E�8lnJ���ݒv�v������j�W}��46�<9�h1̀X��1ni8B�I^�h/`κ1�4��8���j�oY��֨+5�n��#��&m�P�nH `��V,�oQ'b�b�t΢�� <��F�7�Zm1�W�g%�rk�s[�����6������Y� �+flGj�A�dѼ�t*"-�X���Ǟv�O�uy�=Qهz\:s��Z�b��������4�Pv78\�u�!�Yd��إ�#��ݺS�T+�'J۝��e{�oA�[
��2�{c���M�28n��4���6�;:C�I�r�v{���5���g�`�)��v��ob�/��jBrԱ�sj�XI;%�UWIi[�p�ޫa  �kna���m�=�d�ҵk!�E�+;M�9���č�24�X�n�#�w�8	7#tbHO��ݎI�޾̬cE> d��Mc6G;�c��;�Br�z�/�o��\�t�e�X�6�GMg��˜���3Q��휀�wx�J�	�;o�s��蛫r$^�+d!�T|��R@0��	�'� `';gk�x������=�q&yU�)�+�{�[��4�	�9�u-D��IڇU�1�Bj�9�}��'��'����%�2p��W��?jk����z8�
���3N�8���pSF�p�IZOv�-�%��y!�����k:=��:i!k֎ra���
��J#�E5guf�%�k��綠n�yG���k`}_���jȞ�=R�4w��eO�V`K����#��t]���jx;]y2����<���1�� �#��¤�QI�5X,J�Nn����w�.�j��J�;$<0�74�Qp��B�1�`��;�
Z���q�*����5�}Y�X�8͛N�.L
]���81�Ew�7uS�C�xq����K
��0#��s�^Ż6%�id��>�;��owx��\;�%��Ӵ�8�D[y���a��Nh�������6�\ݓF�����x�צw�	v��Ԓ��N�,��uW��E7j�g1�X��($�.����Рǂ[�"���ڣ}ɛ�)<n��U�u;|�Q���`8�Ҵ�{%��9=�k��.�{� Q;��r��#m-I�ؕ�P�u�c8蒢���[�P����Em�IN���q��"�����a5v��V3qY�x���rg=�C���GhʟȞ��~V��j�ш���5tbp	ɍ˭�m&��KY%�ޗ����kmB;�	���맳]#*!�q!���#;����3{�����Ӵc�b:�xI.�G)�V���o:5�ݏ���Z9݄patCn�^tcRQ".Cǻ!�����q�3h �Nܩ�.���p
��9�+'`�]#pf"�&\t!âo4O��V��-����P�9n旝6���Z��^-��ml��CZ�'�.�T�<�'��ש#h=�V˓��^;Tò,��u�&��m#�:�.����`u��˙J�k�fN	��m�hw�� q)ɛx���C��6쐘z�i�ښ��e���VŖ�,��ϱg$;!`���_2�\�G����vw+�P:Zۛ�P��.G�s(XV�t�ӣx;;q�gd�Ǫ4Z_GVF�n)���G8�'�"TҦ��sx3N���0g.Ǽ���;���)�pQ����@��Yk�lx8q2>����ϻ5d�|��I.B�e9x}�9������1��-��z,컭�w!�hj�d}�4�V�.�褨��Uf*Z;����gs�̳F�7�5!EɃ�ך����"�N�j��-�hwk�KZ���n�:@w({#W��ϵX��]9��@��g`�>�C����7q�`��	�	�>y��gqGq1�9�@�-��շ\���GX�[�%F#5���
�p�^�`�n����n���坷E���1� 9A��$v-��q)��-��#�%/B��pa�>x�_ ���U�d�E��	u����ӼH:⶙��ռ�|�-���;N���r\	5�S�r�kX�a�����F<�d폼[��O�u3�.���ɚ����"�<v�K��/?t�}���Q(y8J$��Ox��j��Ǩ`��d�_0|�<�u<�`�tՍ��!Gf�>=�5O�����ݾA^�������� Y�5}�2���>+Myz�+���������P�G���=<�����\�Or����9K>i@��.tv�<��MlR&
���`𬦳0��u�!��V2����J�+h�|�&j��0��8z���Ft=�s,��F�J�SA��O������OeɏC��+"�F�/Fl�6s�p+.Gq����b-�l?���?{�+~I����Oн~������\���I$�I$�I$�ITdؤo5)���]�:��v廘�\���j��J���L�&6@���k.:EW�yH��s���}�t;�9-��l8JgU�K��K�/'KZgJ\��I��tv��o><Q��k*1?9�r���9&����n<ݲ���n�g���,�^�v
�P���On4	Zg��C��(ǋoA�*:�J�2��3]r�j�w�����	�*?nh�,�X^�)�h�����vv�ޙc ��d]�T�c����۾ۺ�'�$�:�}<�����I8wv���44+�N�N|L�ӫt�}�m����z���!�T�}���,������Gj��:�|��B����b!M�tx.	p����U�*DL���ٷSA�Qb}R������������B`y6��!��u��%�xA������<.����e����fs+�y<��ܻ�%�u�3]C�bߕ�6�U���3��������1��,�yuq�gA}��>긽���}\�ؗO����>Oȝ.M6ݚ��G�"�j�����ڹ����<��fX����$wb̕J��I�s6 Q,W+�K��p��Ӵou�wa�H��ݒ�^d��b�qxhz%�@�5x�&�x\>�S�l~ƞ�٠��j������>��+�2���"��������������j�3��'o�=7��SJI>�z˱	�$�p~������yS�
�3I�ۙۡr˽���)���(l6��Lۑ���^E�v�����$�2ʼx�wXͲ�)�N�#�H�����A�����#�%�_U�R	*�k뻧�jx��f�M� �<t�d?}O?1�УF*�@��W����z��,#D��
t�9lٛ���e����4����H�>��(,��7���ஜ�`�g�����}p����"�Ή;Q���y�ػ��ɴ�ҢV����I��p�I��"ו�{�������J�����Ru:�V�y�,o�7�yr�,��w���o�G�u�Л��[�*��
֞��9d]�.�s��r9�YK��Z;�p�ԡ�^��n��zA�U�G�ᶞ��{�k-G�M��r�$6N���W���Y��Q�-+(L�����z�Z#xRj�˭M��!�Uґ�?h��ҳ's���Od���I��O��4^:�K%�*>��j�
��v�hТ�2�U�tS{1��<�C[����׹�|u��*�O>~�[[���g7�x ���K:��o���;X����4:��/�z��yM�񷒩i9�d���v$r��C�>�K�֎���H`�VlY�����eS)�P��]�Ӫnz����rq��U��iQ��=��y6oL �Z~�Pn��E�kڳ��l;�(��"�Sϼ?	S��_M�9��
;U3rt\(`}AjzZ�Yuԭ���|�'�;ۡ�0^g��t��vq�)��,���*S����,A��E^���g�]�(c��8-|y�4c�/�7ςȇ��-z��K��lF���zf�'��>�z���*�3T��*
ǽD���UN�ޑAl������ğ�}��M���a�k�Er�)U�x������֞�6�b�O�}���Ξ��0��D��߽�.�3�i������C��u���"�d��3�fY��.h�GNG]츴nX|6,io6`�ώ&:��t�	0b��<��l��-%�-�μR^��k..�'�ђ��`���[��mo��¤��7�r������5:���f�r���"-�/Ki��#�ыS���5�R��L����ia�h�yM�}��g�in��Ѩ�{T�%U2��S:[5��2��]|yo]��.�ܷ+:�-�$S�h��V�TW.d�G�U�T�?���P�d>_:�;Jʱi<6PT�I ��3k[��Cu!;�����������)c��f��X�w-����j{�G����L~�b�:׬�QM�͎�3���#]�ܱ[�V��Gn�,d�ә�ϙ��������(��旧���ky���ݹ���U��J���!�tg	C&�a
�5���ǒ�ݏ3}���������0�n���c�@���Z�*�8Z��q:3�]=�B�T�a̽08�+_fR^o�0�#�}�� ۞J{�Ԅ9���V{guLr��ç:c�R�͝#LĆ=
۝���U/pX�`Ϳ^�2���"�{zl�(�=���t��7�י�$�VQA`�'[�U�D	z�͜s�\��_I{�xAg7������D�[�<5a�p�hh��|w�@�o���f7�|A���`��=|���\�s�w׹Ўα��#K�*�;\�1�!�|uR���U�k�%�ݖ�㝰I|�.u$�\�	��wِ��l��3}LQZ�v�'��u\�+M�wJq�K��8�%9�P�T������C�W肢m^����P]u�5};���ʰT��޽R�m��c�w���{B�; {;�ќAG��n�x]p��ܭ�VmӴ��/��r�Hg]�==0'zׄp�����=`N/u�G�V���OM��e��D�N�a*��^�kי�ս+]:��[{2��l|EȘ��2�Yw@��E��HUaN��)Q��^�݂i��0�%���l`�y޷~~��y��=u"B���"��x�����@�ϕ3�ϴ�u5�r�r��Y=�Y�j�;& �Z1>��W����Y�Ӫ�n�9�.�$U�ElM�<$�����U����ηRV��C�W�.v�o�����pG~����O��X75��Z�T]ܴ�aZjK��^[::�{�	�ݽ4�ê���MS.[�uئw�bmW#��!�
���s@�S�����6T���)9���i����4zo��Ap�cs�y\�b��� ��LԺo����H�oT����s�H�������{U���K)��{�vp�,m�[z���r�`�Rն:�2�L��l�O���C �LI1��;���r���ؠ�Yщn(���f�o�������t�W޲�L��s\m�p���nڮji�}.�6��^����r����A7<�s�Һ��]/Q��gZz �;	&N[����Lyݢn�5�إ�2T;��U[y�9��L��;k�j���f�
�X4��7N��ٰg����z84�3}�uuI�jGw��*K��sR�Z:�5���c�s����dzHȷxz�X�hAzY����1eA��fj�=��a��<.�)3Wr�� � G�N���p��8�:_GnW.O,;٨��e��k�x�=�Ô �v`�YuT�-���1۽�.�Y��?��xWs��½����Cv�t�k�Q����W���d�}1Q1�6����x����'�ȃj�n��۷\�"�{ܣ2�u0�;�d�|�1�mK!K�ޡUle!4A)r��N땁�Z{E-\�7ž�rn̪���W�m�o�*�������(�����k��/��5v3�{}󜫭1Ub��n�ѥ��7!��)��|���!�i�a�rgc���Y�S�q��.2nl���ùt����!n
q:�}�7��ZWy[��S��me��U�s'o�2��P[��d�����ny��}�r_o�#bԀ�������P����04�jY��'�6�ϙz)����3��U1���v7�n���/��!�v:u�õ�k���J��&��h�=����>߀o��z�+wެ�=h��~c�7�z����q�C�^���N�<4�<8l���Q��l��<9�u�F�����-�{9V%-��X`]]��pM��暦yP�c�h]v�ڂ����nm�:XJ-s��Bz��'Ko������1ur��{z�n8���
�>��9�6ڤgbs;<�AQ���:�������d��=z3r�b�ƛr��p9G��D�Q��A"շs�nM[LsPn=�!86*�OnG�C8�2��T{����øg�"E�ź�i�{�

��g}ى����d"�+ų[X�G�mc��WUƫj��w�����H��#�� �S��{��N��<9@B��&ԕʃJX��;�7�fwr͛AV��
&v�����K+����Wn������F �h"̻�r!ڶfKI���Lܯb�u�� �L�`�,U�Cd���ޚ�Z��4���v?c�}Ŝz�ٝ9�_Tr8��j��/�����z��y�ty��0���e���ֈ������M���Ժ�эh�(��u���{�{O뮋�C'n��Y=�`�j�*8��v�LW�y���*�^}��(0#�ß��ɸ���M�U����<��3�t(���TJq���4�]A���Z�����㺹a/ڟJ��UH����n��b�k�t��;�m״�u92m�"��Fi�*��鎶q91�R�
O8)z��=��"�8�T<�%����6=���x�zW�Gh�l흕ǲ=�"x�=Y�۹�g`"I�j����S�3����a����V��{�?`r�V�	å]c|A��ﲝ s��Q4���7�^Xbdؑ�jwN�z�ogs�,��/v�\;�Fܕ֟���<Y���K�I���H��u<��q�T�1�^>����/�хh�1yڎ/j���j6���G�qD8��ƕ���	Yc �Q�S=�o�w��}1�5jYg[=�1b�\ h��>�B.A���1�܌[���
ud���*K���n�4��*�M$2(���^>��|=O72�ka��#ӌ�aջ==�Q��>�֞��Wje��r���ٱo����N���D�_�+~�^4�Ѓ�m�kC�Ӗq�%⧢_]�:��+���zづ�_���>2㜎=h����o*9[&yڶɳ���%�ą�����(��o%��+B9֣����t��9���zM�ھ��Dw����`ݍ�F���\�Ms*��m�v=���ryK�j���Eu�R;a�5]u*��]���jDrj�z�2}g s�^ո���`|���Z���d<Qٛ�&-�s���S���y͙�flޠ�����A�S�ݭ��+S�xQ���^��6'w�Z�{u,�p�ƹ����+!�X�u�x��kǀ��gEĭ���Dǻ�T�ݹ�bꧻ}��H2d�v� �!!��&jY�OX ���T�7�o+�2*�ݾGd����3}n��)۽~�����f�#!;g��=�9�w<=�^b����G���+y�T!�����lTC]r���g0l�ۂ�FF�>w}�za����(E������|㺵K����gp4:�a���]��� �],d-dO��E��Vkh�k���r��7#��T�\�\($'1Gk����S�v��y�^�ski�ḨJwÞ:�x1-�M�Q�<�}�g�z֦�хb�z�.vG�����N�!��̼o'�9J ���߆3��;Q��o7�V�6e�|�`P79�EG����K�09�{�wF����qH�m Gjh8�-���]_]=�sFzۀjʃ<���Ywҹ�G�6>>��o{˱�"�g�.��7�˶���C���f��u�+�4'sJ1�����7�Ae薹�z�nnL�QGB������Z��˝��7���3D)���gV�lU�[AƤ#l��6��_ZMf�t{���%����I��2xj�W�㪕��R�YҌ��,�Wd�F�d�_.)L�r<x�Y����0�Fw<�ݓlՌۙQ��cglq��P���c�=ÞZ���'�ޣ:>U�'<і��p��������o��T��ٗ��`�i)��F�Q��|����c]�mYǻ�V��z�9EJ#���<#�#[.�:�n0��4�%�Yn/nT�T����2��Т���E�"y�ޱ���������clA2��؛'�a{�e#~�c1�tŠU\[�������A#7���ܚ�C��!��\y}R�Τ+����+���5B���j��q���r�z�]}��}���[\��nr[��6��R�N��%,Q/ 8^v	���,�/�����[R:��?�]��slV8X��Yj>�}�G�0Gq+���6U�6��F��/q���J}��e�8S��*�Q�����Lˣ�<��D!�ѯ {̾C��T��vzN�.=�yj<.�'{˂�x1�����Q��5?"`��pz1~�]�cFv�8��l�{�&�f�4��jm��UL�T���4�p��|U��V;Dq����1�1_b[�70��Q�kq)1R�3�x�sQݜ�|��G��=�맞������)�jOr����.��Y��;0�E��,�V߿��Ai����^�"��V1k���t$έă]�5�Kb�bs��ufb��L2�(�֪א��TW�S�3.sU�S:�1�X����أ���;c���)�2���k��r;�����ڱ�p�\�\g���Ѹ�M�T���&�$��j7ݽ����V��s$��rmAu���|��T=;ξ�ض6t�׶�75le����
���bQν�ܤ�I$�I$�I$�I$�I$�I$�I$�I$ݚ�o��I��#�I$�I$�I$�I$�I'3�7�0�T��8���~(�3�et
{��l�u���x�$�p�2�i�q/�Qjm��S!��ǃ����lD�q�Z����`1i	4��� O��9�"�$Q� ��Kb��M���/��Ug�A�h"�4����lP�2�0$'���x�7��Ɩ3��Rl�p�6���e�~@8�s�����aE��	�/���"'!C(0	�����(��Y��DTU5Auj����dvH "/(����1�1Å�%2�W�l���l��+>�&��>��2-Ծ*�T.� D�׻nE]מ�h=���e�vu���:Ɛ�;c�![�[�~�Pk=UY��7s"��q2�;� ����e����b�A�{%ޖ<x{�l�f�H�D��/��6�^Ǎ(;��]�m-�4�����M��w��-�&������¼��?7J��}�_o� {����MſI7d�d��U�'���Ɇ������x`�eU��^u���_j�ϰܴ�d*㏾���l��[t��YU��E|y�����/�|xSזŘ�r��`B�\�nD�����S_y?Wc }9;��3���?{5h�E6z��=�j~3g��7.1͛��um�O'�:�+�s�2����X~��f{/�l�f��;5޼Ԯ���Cv.�	>�*���w��K��Э�f}�F�k��(��L�q��H��7.���{;�QO]�|Ǧ:�u^�^��z����O�<��k~�b��k��b�{+v����U��X�iJ�h">�^^��j��!�r:U�WΤ��r�um)4t�r�F5#�k�U)�\p�wAB��b���3U9.��8/PF�H�V�ۚ��̚'�����c�(|�p������%Ś����S>�d���p���x�=��|����̈́7��_�r��{f,�½�.�e=���'��y��R��t��$mV�N,�rU�8�mbFc�*�[K���b
l�쫘7,8�X����fy)����e+~���"<Oa�|w��%΅��6�����$�h�Q?S�gxϐ1�grA�H���g��<{���Kcaoo6������#�K�xrbOIg/g6X{x�3i�:
���]��hn�w]��lY9P9#GK��K��맴֪_rޕj�U5.�IӲw���{����hFB�=��7i>������[sû<���׽ǭ@�"A��[}�y-�{�o�j|�1}�W�~�����������hL{�Gk����a^�>by�q������{]فjpw�*��Ա˦čΡ��t�W��m��c�飖(����,gj,ȏj�x��r�xx\�<���ݾ�������:��-C9	�ⰺ�X�������lGh&���΂��_C��;z	"X�����V�.k5lW���ƣ��p���hèJj��_�ȿI'��H�Qܶr�<�^�崆p���$+MRg�}����遼x�����U��,\XgI���,=̿.�|�[�r��}ݹfڕ@��Nqv����$��8g\�5���C��^��g7������{�:u�8e�ݕ�s������_�bF�\܈�nn����6�[J9��
c��١�WJ�hX�=�
�7FЬ�j-�Pቕ�F����ܺ�&!w�h�����L=3���T��omq�B�%����ᅈ� 'pR����7NSĽ�뿻͔䨰GF���[=)e����o)�.u���[�;h���r�N��YZ\�6�h=�V �����@�~Y�P�H��z���Z~�cg�e��`���۫��<�%�9~�a�ר��F1 p���޵y���#�����rYv5S}����h7�Va:~ڕǻ�1x-�!�|�-�g�1Gey4 �Oz�?=Oo���3��3�KN5��w����-���Dfk�����=�={�s����.���S	���/����q���^>K���O�_��ͭ�=D�Rw�ۼi�x�8��Һ��%A�єkɹ�=�W��j��,YZ�1���9�:��Y�
�`rƮ�F-&�C5�Wwr�A׸����=��Q=wI�AA����ְ	r#�G��W6a5���%�6���pFr͐mT��>.��˻4�ok�rgZ����e噩��;����Wo��g&���r� �@9���}�61�˽�yfg4�×P�w��E�և9Brz��*�'��re�%�iQ�z�4D���眵Ǝ��_��H�x�gS�m\�I��llO�'o���#(�Z�v%䛼+���Uj�bf�u����r�M3�x��Y��F��h
�kc���=m�ޭ��>�� �V0���#7�2rX�3w�HDQ�\ٷ�j�n�����B���|o�3HLYîa��`5�⾠�r����0O-�ߌ�I���+ѽϳG�����E��T�N�}�>��!ˀ�����j~�}��� �ۖƫ�w�*�uǫD����x�=�ݓC�$+��n���q+���v0����=��R��0{���C��@ǯ&>��Vx��[ʥW3B"�P���n�'��2�I�����p�Q���@�젹���[��wo<c������ӽ-U0w�Ȯ�!�8�EȊ��l�<j�Ol����Γ�(\����i}���i�1�Q8���JOF��8�띀[��e�F+���v��9�H�y!�땩�=�{�k%�kV�����c��p�F���4ʓ��
\6�L޹�J�j�˱T$��`J�u����>I^.��5]��h�K�o�zyn/`�p)�J��X�A<B�0��J�]f'�ǻ�m;�b��w�5`��Lv�B.��ۭN%K7�Ӂ���{���ӏ��fѩ� �R.�)p_���������؈G�o	ڡx�w�{���g�э�'��U1�S�v��7�M]��&*�?n6 �2�<u��{C%^��=�^�Ԉ%���0v�W�������ld��[�A�*/_J5�]�=g�qh-H=/���9[K��d��2���W02ިwM^�j�N}�����\��'f]wC���%�݌!�@n�d�&]Չ����p�_���8�E�J�[�#x?K���7گ�W��[{VC;t���(�_t�8E�S������{|X��G9�uZ�uXZ���t�"��{����ʲ��P�n�[i��Ԟ����\#��e�A��w^_ Ec̳��TB8k��x"�|���R}X<l|���<}��	��-|�K���vl|�/		Noz�9�X����̚��kr���Aѳp�u℮c�e�[��:ls�ZN[��Z��L�Y�'��lpW 缽'"H~��[�{i�-�l���[v�i�=���{3:<�	�9�����Z�Z'Fޤ��\h&�5��4�Jˏ�W\�;A�qi��7#O�ڳ���V&�{^\���ʻ=����������s��>�`��ǎ�;z�I\ꂑKW�]�u+q�Uݷ&r#wt�"�qM[�,�r��&=��X���>O�^U	p���`غ���\of��YE^5T�Դa���OhΪ�b !���}����p��M�{}/��j�v�Ϛ��:��F��<9S;�
V�,��͠�C�w*�[�G��]�\�b>��X�˕��냼�T��{���Q7�{u����s�&�'��8��C�	a�< ��#\�s�s�]ķR�X��s�<������x����
;.[��Ǝ�)$;@=W}*��I��	R��\˽�F�A�uZ���Y�|�
�>�"I�{wE��V��d���\���b��Cf�&A��+�f�l���o2�Ef3Gei�.���%%O^��Jɔ{	ӣq�F��l\��]b���a�]�b�Nۺ2k`�}���ש�)
W�x�kʗ�)��-��U� q��Ƙ2�ĳ��|<��pS�	_���ka��<�Wv`Շ��#��y��ڵ����hG��[�[W5#�LFG�
�H�����n�8zv��p���\�<���s��YvQE^!	��N�P�$�t>rm��<ٮ�6��Ʒp���{q<�=j,�4K�ң���`��;ϕFo&��Q�yA�������gK�U���S����� �s8.�<�wM<���ݼ���|<R�8}���wrp���ԧ.7�H��ZCgp���kdpV�G:�JV�F<�h.w2��:L��=uq�/x��	y�
T����c�H��\(��Ǿ�A���������{�w�S�U���"��Y�
����ġ{��@�Q��l�v��mܣ���,�d��@u��s�3/S��������h�hW6}n����P	��Y"����W9� .��b�tg��� ��d�h��9�ѣ���x�>5�!Ɋ������$j�#��u}��:&��j1��X\�Wt����T�}`�%`�|�:p�K�z,J<q۸�p��U7w�b�;-���E_Cxv:�Ӽy���ʱ�t�,����8��$y�{�qy.-csU`^���)��t��v���hק���e�C������j�եM٤�`�Zn'�i�R�Ҵ���T�RI놅��eD�P[X\��k$�8!W�u"�]P�A�VY��`�i���7��.�q\N{]ެ7�Ș0!�9����.;��)�oP�����'��^Y�s/E�Mq��Dj�O��Ꝫ���1i�c.O�Ƕ�J#L���tM��.��5ŽM�{`�N�#��uu�+8mFm��]U�UJ���yn$��Z�!������87�_l�u;���+o�����3���	d�
>2.�|J�F��'���{Js�#��7m"�锷����>>Wf=-�k�_�-.s�Z�|�����Z�<�˛���
���%������y)���X��.����t$���������c)��|�/�����+�=Oe��oBC���u��h�;�XEf�)���ɉ�
��u&Nz�ˎc����x 2��Cx�n��6�YhƵe�W6�����+�EU;x�[�vQ�d(���%��-��-t��סŋ��+��FJ�������r�"�#+:��ѫ�"F�N&w�����X;��f�����g�|�r��n��T:+0j`��)Bv�)b��7u{Ս�X�	���B���I�z�L��7���z����[�=��q�ڊ��x��>�ǳI�΄��g� �/1���sJ�噒Y'�x-nq)Р�i�H�{���vw'�K��q�;F����*fv:�NWtO����v&�^�뵹��1��+s�������Th8��2��W۞���P���qx�r����XK�i����B{z�&4���Cźx�e���Ť�ncHe��;p�P��wC�z�:tRGB�q�����uZGᲜ49]�f�#�ٳ��=;<,K�{�Q=�u�\�c�x�Wy]��NC=�2g(=8 ��p��ٽR�qa���3���|%3f��d!�{��vʮOn��R��2ku�{'�7�(�r���c{���j'n=�H�ۚ�/ޱldop8cްb�M�Urp�{��˸yT޹{��w]֘[�+���1�V�Va_=�ҧ�pc�.vpx7h��7�bɸ�����ucwh�1v�2v�n�s�7P[�hP\��4!�ؗ-BV
T�����:d���Npw�>ĻsY�xf=6֩%�[G�[��.����sȗ/Y�C=�痝��mї�k���D�<�7�s���_QD>���)p�|�wc�w/nM\Å�!�5�\��(w�i�iWє�O��&�8#%��[���i�Ym5�kLS���a�[(ݮj�^UW�����(�3ҕ�>����z�-+|�i�h���~̾�~�<���u	��N�;���<=u�>u2��\T͖ꪖ��a�6�)qK;}��w\�*D����0��C{�"G^�/	3F�ĭ�SNk޻���r��u��'��P����ҵPHUn��^
�C�l�rSYYGMPE*�~/(��f��O��}�A>�ɚ��2���`�"s��d��1�@���.Q���n����xs��G�W}��R�6+��ƪm�R"���'�����:��K[�U����n�mMA�8o\2�7�r�[SU�ف�v2�ki�߰�$�/�������M;3g�Q�Q_WEǚ��w��fm^�]'�3�0l�u9]�-�.�Yb��8g�:���Lt5�Ǽ�sٗ&�Om���q��%̠ygAOs]�4^�<���
���K��"��t�%	+��=�s/�[�x��l�k��b��UL_,�Y�*�ۗ��|wr��A<�c�T]��Z*�t�Ӹ檃�<��/8s����PY'�]Ϩ������W�Z����S�S�4����5�|���/iI����=/E��D�4���cY����u嚃�X<������ݻ(XXK���x��\�/O<}�~W�ޣ���ً_b򸳽���Rܾ�]$&���e�1�t^�c2I��?�0��y��x��&�Ӷv\[�M=��+6zr7�o%j!ش������8�iۏ���V+�\��Lm��́p�&8��M�[�sH��{���O�xP\�oۅ>rb�7�����6Ԛ�%E u�ʄ��FɁ���;�=	g�⳹��t1e��R_���h����>�x|��|�<�v>��W��s�ym�=� #E�ecg������`���5�Sɏzw* �_Y�*k��X�HqWf*i*i� OB��Kt}�\_o��g�,bx�7td�����Q,��݄��~A���ys�xwb��.h٬�*1ǩ��4�mfșפZr��dB��$�^����f�(->ѯ���;�0�<ej�f�R�Пy�s�rPo(ZB��mQ�k���ˋv�˳��Sq�x,�m�$c%uv�&:}5�{:iw�zf�:��)]�n{�"ie���T��oLJ����� Opt��SƳ�=����r�&A�`��Զ�k5�c�rg33���S������1�Ȓ~�a���5��jU%�u��)�-��U��@��9��g�2�wi��&ޭ/��}�:����;�}�.%���ǁ�� ��wxn�����S77{7{�͓�f͛6}�����|������}��W>� h~�����U,���>Ο���}6U�É����N+�y�e��i�zܸs����i�r��K���3f#��ӗ;H�j�l�Yeپn��i��t�_D���wz5�C��;w8�%1��w���K�1�~8�Ow�f�W��M�	k�y�c������w�2�^��c�-�������-8e/��ot/t3O��\Ѹ���l��'rt��t�v��s�b�\���
��r�m��hB��:�_E��a���ާ���$���.�_'���E��j�\��\�]�w��c�0�%���SR�O�3����4�g/�.�����mq͉�9�n�Ӷ_a7�:<*�Gs���L�P�^�5���p��\�Ms�Ѳ�+��uCB����Nk���>�]����\%Ͻ�$ޫ���Gk���M�VWk��㍾��G�Al�elo<�2���N���g���y�a�{U�(i>����� fU;s\I�=�#Rs��ylt�O�jҖt�o��.H��Q��ʟJ��1��,<�^ԉl���(������(����g��=[�V��N=�v���*e�;*o�+��	&�:����.��X�.	2�$R�R�D{.0�I���>�x`�?MIGz�V�㧴ۍy�Z�=hL7�P�/7�_P1iؘĚn�����|/�iI$�;�l���{{t(o�С���'�2
,��p�P0$�7>~�QESET�0RP�UT��4�z�Ss:(�
��*)�q�����(�*%�ɨ�Zbb��<��3I$�e�*���
�	"*�����LQTQEQH{�^�h�֒-8��glF��G �¶�h5E���6T'�`9�cNf ���+�h�������U(���a��(bX�b"J64JET���SITU41U�U4�\�IAKF���S�4�UR���4PUQLMؠ�5�������+�j��CAAC04UA^%�IM!�qSCTPRDQT4h�^��Zf �b�"��^;�^���S�y��~��>}�L�N�n��'�R]�'Qm7v'xB��{�\ү���I	>G/N��t��������y�3N-��@�,]ؕc)F�A;��/s����	�f��"�	퍼3>XJ
�վ�wg���EI$�}L�e��dh�gq�?#�{G�-�y�Y��V��|�WJ�r�
� ��.cH��r���� '��&����a����o:vx�ި�]o�L,�$[�H�����݂M���o�fא/=���n>~u�O}a��$��Y�����c�i��W��ԽM���/L���d�޾w����"�?���Xg����d#5����ѷe��d��AgbG]�Oq���`Z�PdP�U7{��V\��W�ؙJ�o�cz��-������ﵼ��̠����3��ީ�ˣU~��a�
z��A�Ř���o�|���G�~^��fV�E��ϣW��}:�*_���JC�A��\��3ޚ+�;D����:�[�U@��͜rl8�VУ6k��Ǌ�7��i�1�g���x��ҡ|�ui�����z͙�@jDq e�,=󚯼Tp+,Ł���V{�i|T�|׷��T�`�������L����+�Nq��͔������ǫ�n�ԋ7^���&���A�D!�f�M`��ʐ���o�VvM콽U�k�9�x&�뿢1�n�P�G�;&𜆓��-9���szs5��ua�H �!�f���tG����o��7�E�=��o���YM�v��L�����[�p�)^3�뉍�
���"��`�o{�݋s���෸�FO�����杘�6�yf��g�����b}P��=<ly�9�hFD��|�ϗL�ܩ%׶zX����~�,��Q�W��������N���=��=Ŭ��G�V$:O�5�$��d��W�n�i�M3Ǉ\x��&6ۇk�T�Ms�M8[��׆Wt�cz�'@��O{��z��ȃk�
�\�R�{+ԋ{i��fM����l7���S<��3���N�]K�����X6��0�Ozd��4<��h隇*'�v�uӅ����0�|�/͑���%m��j�tp�5���:r7xr�L�xI�E�:�ʙp����/9w���/��j�nr���6��Hн��ݾ��|���"c��g��X�c8p,H�����	k�M=W;���tߘ�M�q��2�1M\F�E���o��G��V\���;�1�g'l�k׃�n*�k͝��cf�Z�g���J,)b�t<�o��3�'n��>�����Wv�u��%�-3[���d�;�V��}���r���i57�*V�3�Y缲�	2�'��Ǣ�[�G<�?�upz��tɗ�L�MVKr��nx<����Z��y�0V�G�/��s��=*��p1�be���=�ӿ��s�2T�$0!��w�l�H�/}�z�A���^�����o}�9l��v�[�I��ϟ�%]V�B�!�U��~��%�m�Y��#�����ٛx�J�{���С�S�� T}ֶ���U���mV���o(�p���a;"����jo`][���O�&]߶�7x���:�/P����"tXz<��44~L�S�ū��b��'^ۍ�������V������{�Pݩ��xs�2W�fb�=^}���K���w.ɗ��.��r�݇7�q���ɹ�*���|�w���Íd	����=M���	��\u3�j���]����xw��Z�~.~�;������8�y��&�t��G�mDA�iKWn�}̏�-{=ժUT�tw���𾳣I#�׻�'��j�knc�q����/U�uf�ƞ~-H���G������z�$�n<h6�r\wq��{Lg�:����ST�S��SM�A��|<�\�_�>��}���zy.�S4����kM\X������<�ء�A�P7�~y�ɓb�g�)���>�����d�//�=���`~Ux�!uu���t�wo��r-�~�y�s�w���秹�d�spZ����P�BwA2�Ene��^��x�$���K�{}����~�=����|Z�O>�?�|�o�!�u	ʓ7l]�����e��'s�Ga=M�d���c���1������o{��������77��J�Ġ���;9v��2��	�{��xp�{���:�������n
�Uui�'9xڱ� �`_����X_�o5^/�M���s�<��[�z�i���!��&yv5z��}�� 0 R ��IZ��bg�
��!	H{@����Oy:n.�$�3�Z�s:o(��J{ܳ]{4l�6��tD�!ҫ���}ޜwl��ɦ�k��]��<��$jcqҬD7��L��p�᳁����v�
c'7}`o��)�s|f�L���>�}����H,Y�w�����=�o�ǨΊ����t-���^�����ѩ�z��^ͺx~���`8=�+md[O���ނ�Tӟ�-S�ݿI�`鞡띨G�r�[��=��ݰ\]��GEm���|�X��^�<m �s��'�mX�x� �a}Ug����G���O�-�}V�*I"������@n��xOY�勅����e�z�����
��z{=y[�ؑ �>��p7�}6���X�ڤ����/ӯ����{߄�6d �>����a."�3��v|>�4��<�52��^���O�g�U!����5�(
��vX�D��6.�Aq���4��x%��$�w:�������i-J���2E%����z¬��:�}���S��X �S_%9�%���ئ���ضn��u�Y�lXE����k��-����#�����/�a����4cY/�ۺ{���ޤ�(o�Y��3��-�$�����`{��k�]�Z�ǳՊ*��5t8��|�-��&�G���;\c��'b.D�����#3N��nX��^_Pa�9~��6z�b�{L��מqk=j�V�u*>�H�d��P�%~�&�O��*�
J(zY��V>U�R^�*��8߼�zׄ�-GG��~g�]�6g�EKwDxD:o����3��y��N���)��w-����wL�����m���t|'�Ƚ!�܈�r�r<��<��sj�K�k� ���zCW�}�;�
uy�d=ٓ7ok�1W�������{��ƉB��4h��k�1l��o�{�o�����,��'�K~�{m]���l���z����v$Sq��q9��40��8���k��v6�.6��e0��c/6�jw{�y��p����ݓ˯ʼ�N8������M��'/C�'�u����,���
H���50����I����}��}.��9���뤩�w�o���5}�&�%���n����@fÜ΂n�V8���
�u��V��X�K��~������g�@����f~�<8����o�3m�ҕ9qՎ���3=��K����5^}�.oX)�k�a����ו����T�
mO>���󩞞����'LԒ��WuVW���5W�r����
��v`��4/�GY�ޓ���|�;�.�Uw���A�QMDP�b�V`h�>�v)��}���w�/=��*�K�LƠ�W6W�s"�����x;�WT	�݂<�x��2a��{��u]��z��w�)�O�9y�n{o~�L#�mkꁘ��9�j5�
Va�m�ͮO`ɱ���;���y8�12��[�N�R���Oz��.�>����d���y�T��~������<fdB,?��1�`���>�9�O�ٓ��S���>f]`��*vSף������<6�C�~+t�n~�=�6��F==�j���Y�b�E��zn�N��x\�H�^ƻ�w�����Y5Lf�g^�l�]*��:���M�۴��Y�e�Rl8b�D#q�������2�.�>
{�q�~�J}C%����.Db8L^���o���Zó�\ڛfxz��%��{��=Y��g�`8�Og������[wWS����:u<�kܵc�/Q����8n�p��z�����9Y�[�	�y��[N=�}�X$����R�F�P�N���&:��5Owg����wǀ_���߅���t��i��E�?O�P~����Z�]��ś 휇���<��P�Nt��lӚ����S��Nf��o7�@/��3����;!��A�xߜ��pM�Ok�E����tq�k���Ӎz�`���+�=��An��I#�{��mw���pl��n������s?}]���_�<��v_����}����̦��K��^���Sv"e`�
t�P�@�.��ˏ�V��شv�ٗ_~q6(��c����R��So	UW�Ώ@��#��pL#�}��g�6�=�`;��t�y��{�����[]�$5n��f��u��G�L�[���M�4Ofh���3��\.���:t����%g��7����ҧ��~�Vo9}v�>++����f`�]��_Z�_jR��y�tL�݆�����k����y��ϸq���\�o���fz�I�靳@�������|�ٹ�bn������oD�Yj
�"\���<D׳�y=�-���{��'�����/=�g��K�y��ޑF|�ONH9#s�|;	�vr�;�^9m���MO�g��Wz��Խ+N����N��z�C��{�N����%�zߍ	�rS�3�����Cc�������uY��͏��#-Vp�}����E>��'�x����$��?4�k���d��`��y�7I,�v��r-O|w�:�����Ͻ/�3V���	�xO[~����r�ޚ`LRW+�}����ts�GOf�rh���'������}�y8�����������r,F3"�ɨ��;kfn0w>6d������ߣ�E���I�*q$���q]��1Tp4�T[8�4U��p���ؙ�g5��ׅXfe�eRHC^��{�١������b�����-�`�&�r�`V7�G-�:`�ȮlX^칮�1TE��]�ruΔ�-�fY���MH���Mj�ɻɉs4�4m�v �|"���������ϭd������������.�季7��i��ð\���ӽ�Q���K���u;����&��^�I㡶�
�>K�A��>��p5B�v�����񞅺��~f�g��������T�&
��<<:�h��K~���5A��ܿm��ŧ��OIa'��G��A���·�d@��>�Ճm��q�-c:��$צt�;���پn^�l���=����M-�̏�����Sh{�T�9���M���z�;���� ƶT�Up�R�z��p�^{��mz��è���Թs�?��P�͘2ߝ=}ݸ՜�j{d��|ٯ��ol���>6�0�������`���k�L�:��� ��ĽY�?�~ߺ���6`����EKwD~=���Bg>߯_������z�z��ׯ���o���߾�_���pN�NzxC}�`����Jz���yC�������k��2�QX�y	z��	�N�u�ȱ��J����n/R1e�|�'��٭�E��w�=�6�1ãH��ͼ�5��'o���g��2�t�sZ"�;%�ǬxA������ W2��T>B+��"��@��
'(�
�3aBi4aڛD�v3����t�2Q��
�8/�b�n�vT��Y'��H���P�?M~�w��m�P>w}7��P�e�ՄeI��qZ�:eA�.Zh����C�Q��}1Ң�Dn�o��&)�"�ỗ�̽�Yn�#�L=�����`�_����;E���]Nꚗ\e�\��s�u�!��G��h߈�j���z{��:��-*j����zԺG�_}\-��c�s���Z+f̫řt�Z��q�[��-Sih8Q\��ˡkI��\���/�n/���<W)21�
�!���4)��A��X�GU�t��:�Г���X*U�(k9j]�Ir���B�_�5����~@y%u�w�n��T�KEBo7�:�It����,:���12�9b�I}�C�4�V91g=��(ͫQLƮXti`���>�=�݌�EY洂_U�ˠ�G#���P���o����p��
����P�y�;�����#A|qk�z�n�IdO5s��(Y�s��DS���"�'v����ϙ�za� ���塐����1���Y��!%��uD�������Xi�c�t
grF�mrp88b�A߽N�l�2�;��;��6�B|-?{���xN=�o��];��N ��[w�s��3OQo���v�ݓ�T��-+�4�iӋ������;�$4��^u��a��X��l�ϡ��U��r�ҷ����Q	7�se���"�K���!N�驤lrZ���ɤ�8��x���]���a���+�ж{ƦcPo�L9G��{�����������C���x"�v��f��N�ّ��Z�߾�k�8�㲱wm�y�e�tWa��r;�=����#ؔ��m�ݫac	��dŽ��j�B��.��:y�Fz��٭�z��s~��|M��k���x��c��C7d���b&�wow��Wݴ4�ZΌ��NdF3��.�h���@@�|z��67�9�Zm�(��K#�;�!%.nB~��vK�N[�:�X��ʷ�'F��
{��`6�{�M2�;���nvn���<86m 2����}�S���=O"	N�]�x�(�	����j��S ����foSS#��!.�ZwΆ��Y��+xw$k2���d��r���=����W�sN��~Ib*��{c|���i(M���"�5�Z�i�5C-U�\����(i��n���̎]�e
�,,��,�[|�Aj����������vo�>����?3�R]b�]�L�ܼ!etk��H�?��4�ADTPw(��	�*��gMi:T2ET��`4W-Q�QR3a4�AME%A:],BD+CE45E4��E�ꐂj&��j��i�t/�yLIAU��sf�((&Z(��*$J��EH�I$4PW��li�����Z)���j�"~��E)F�Jj�)��8�(y&#�b���X��4DE��K�լi<�q��AZ9���a��i�`��S��VUkm��Y58��mA9-���9i��8$�Hղ�l���V�ImgV�P���9'���ՒM9ڇX�E���<1V�i���i4ju���gZ�\��܃�Rf�f�8�TA��B0}����g߼?~[�ɟ�9n��_t�P{p�ݝu��O�^}�~.�d!Ҡ}�[�ڂ��/$t*U��<��X�|��&,���y�����C!�d�c���D'Ě���-Ǧ���ϯ&������Q��b����F�{g�$*jo��M C����k<;�Y���+��X?]�E��p+��h�J�k.K���h�p�ȼ������dFT��O=ɛj��m�2�+QL �ձ�D�Ũ'�bv����t�{��5N?�e�'��焙� �?~>�U��BUc�N�?����ޜ��!�[9��Z;/���R�#���gXP���[ռ�|w>
N
���	"�����%k�5;�UӔد9��t�dA	�x��E�#4�%*SS���s����)���'�$�67���	�}�s!p��l1Zi�����]'�9�N�t�eE*Mmq�<���tx����'�Y �WLw;!�����̛�9,ʽT�x7ݰ��2L8��5�|��ct�O�Xs{�"�����A���'�y�0����smzc�l�O5��H�㐛������r�5�%�a�ۢv��7
�p�Ӎu���M0�T�=����Xb9��Ĳ羬�n�Q��~ �/�?����?xz~�d�_��_������ض?m⡏��%�%��f��U>�ǬQ*
��'�'���Fʼ���,ʧ#�S��f���`��Bl#8l9�i:A��#[ƨ�<j!��U�[�Fnj���AMĖjɒ":����sz�De�z����LK���}��+����i�*�[1�¼����0���n��~����y�;s��άy��7����M
T�xnbڞ�Ή�:�2�>�o�<��O��D�ۆ���c����r�C� ��W�nt��_c�%r��� p��4�z�]c����^5���������S�g�ۇ���"<���|�N����ve@�pk�7�|���0��5_k�P~;?'7C�\"D��(��nZ�{�o�=i��M]K��?C=����v�h�M10��f�ȁ�A���	�.W�˱i&?���8�ຎi���:u���
��1��:�,(T<�!�4�������}�Q���l� S����߽�-:��M�_W-k���]����qt��2nn�o?�=�51��ܒ��^�V0n��
�U�������<����b����E�b�n@�t�9�����$���q��0W[�r�O�C3��j��M�/�	S6Ԕ|>}k ���Ɗ5�������ﭠ;:
<-��/�r�L�.�y���[��p�c��ėiβj�L.z~��-{&):ZdJ*�0��Qm=�p釧��p�߹Aש��]Ö��xo��4/t�WN}�;�
GF��E����|v��K;ql&��]J���w�8����:���a�94UnT7G`KS�^%��tb�9BM��8I��W���r�u���WY��}.����d>�xwbղ�޾!����g�^�1���ȣ��O��}謭h��l��u�����C5|&9;N�p��%���$��%:��Q�	�'�ǫ6�sfQ<�WY�����R�y�P���HB1�C�H�!��˷���#��&@�LS��:��p9�t�r��[�p�at�PWp�;�0���%#Y�ρ?` �y�%�5�,x��3��/�m�=�jޛ��E�09�o<����'ȯpг�q3���{�_��6r�k��7���=2!�Jۍ����C�G%s��I�RX�-�a)�" Yڎ��G|?��ӥ:�K�:xOژL�]��kz�eEs���(Y�I�`���,��U~�Z���}l�� �v����3�5��Y���N�1��̠��R9��MVJ�[�c���Le����W6nĝ������/��� ;ָaA�̂���0�ږe�;h��u*�tֽ�&Y�_��ԫ�\��w�z;e�Q&2�5���^��3�2%� �`<h��<�o�0̏�9ޗn��F��[�zl,��^l�v�ռ�� 7��נT˴�lk�[9yחx@��#�<���s���|���o�5r����)�����5�]�{��{���%�4�{�}����\s��4��իe+��Ƹ���L��WH�i=B���͡/H}����p �|�=�o��5Wml�ٵ�{���#�˺fvdwIg��͗&�B���8�5��������1_��}���s�w�*;���G �C��_��TB&f]Έ�T:&����d!_��^��P"�����+x7N��B�/�ٷy����݋A���/~�x������덧M^鋇TE3���}�0EY�/}����)`�C渑sX�_�TcR����\�-~aK*D� �<��zm�O6g�&����}�O��D=/ρ����h��v��1N2V'j[���D���L�x,4)8q뮛����A���NT�by ^:�o"���Ʉ��`$$vW�k����ż�����x_bk�ᝦ��ځ2X�)*���X�����Hqm:A��;<of�����U�>A]���!�t!��NS<ht�O����vT�����5TB}�֐]��L8�q7n%aTޗ;:E�+�M"{�L>��(�ahԢ�tS*��P�F9j�����Zp?X�)���`r����,�h�cB`k�"N��(➗�1i���Ac^]&���p�bƪ�Y��vˆ������!.����F�WT�uf��'h��ʓ.E��s6��s��o6
��fH܅T&tƶ��7��'i�������7�_�%���=�O`�'���9]Θ�����O��WA�j��&Jc$����ކu���9^u6tkz�0%\ik�c��-���sw=2:C�槴E�/�ؖ���h��g���߽�o�c�i�B���)����h`8�p�`}��k�{ji�_U�V#S��W�,I�\���������Q�b��9/պ��e�t&A��:g�|��`9��¾���Ţ8��QL��_P\s����SN�z��?I���z��(s�q���G����Q�cF,3�.�p0�Eݣ_�f�!*��Ҕn&`�}�����q�E��D��{	h�:"����GD��9o��{�a���[�~E�o;;�S��z{��j3\��^gv�����	@� ����_E���a������+���٪>�S���hC�.�x4k�����5�w3Ez�K@���#&;y�b�ڃ�qm;���Vw)�V](<��Yq~<����:���g��*m��m�i�[�`�.qUg]JUo�X*�kAN�>GxߴLM�ê��Q{�Kǧ�J�id�N�+j����r���¼k�ݷ�5�̂�4�£:�üP�o�G7�~���Em�Z����E,ݓ���3�y�0%]E��A1,��Fi��R��]���ơ�l���� ������v�+P5%�2ښ�����q���b��؃��VR���Ŷ��Y�a�@GC���.��f���w�z��)�d��"����{�u�`��x{���ZhX���Ϋ���؉���o�y�/yd��1�㻅:g!Ӟ�n#�1�����Y\���#�]�o�懫�7���>��v��������<nG�~��v4�$vI���'��=>fN�@�\
T�����|"��{�z)�8�E�|���h>A	�ni{,����v
@�ކ;��O�s���t�T�a��͹���q�D��~���t�.[�;Gb�t����� ��}!�Bn�& !�}�%�=�R� �&�~/I��z�CS��'�,��%u����3��_?n<�L�	�?K�X(ZD�wf�:���\�7ݣ�W5��Ψ�ЯO�ĕ���������z���!�����% S�H���E�����������U
�M��d�5g���Q��&;-J7���O�Vǋz�S�Q�{�ͺ���#�?)vg�[4f�:��-��K�mCs�{�P���)�Ë>����������K�_i�ˍL�`�}��y8�W�m��ˁvt�kkH������M�;M4���Nf�Q"8y�y��_��`34�|�:�Z��:�c�Y�D�R�/>���s;hNX0���H�J��?<��hEf��q�b�>���]��e�fN��]'�{�������<;�E�4��I��N6۞��fY�d>߇߿��?������MFp?�!f��M� ��-N�6�fa(ct��Q�]}b�ms��������6��[�j�J���R�0Vɂ_ɬ8��|���;簍��W�9Yg�ߋ��+����]�u�m��֡����خ�����h+	��*���}��C�}�x?�������+y�k�o�Ͷ��eç3��3<]+�琕�n~X��-�5P�ߪ�}\�;��A\�[��{��}��=����G �jdA+��3���6ʲ���z�`���A?��w\pϊg]�\�_�)���br)y��h��ׇ}('�P%�����c��*.=�4�f�j��{a��M�^��$"y���]�i�b����Ѓ ��yN�t�&d��Am�0��1M�׶�V����j��c��D&��,�S	;N�p��M�OЙ'��%:��m��VF��C8]��Pɼ�S�r�Q���`�E�y1Ӎ萃z1���!�e#n]�4�t�H��dɼ�-14��1�/iF�i�C���&����D���>����"��n��G<���o5���j��Qu��d_u(k3�I)�E�y�h����l:	Q�=V??2k¤ wl��6����-]Eo���6�
'e0�9+�Z�˔�MV�ƹm;	O����|y[�J��C޳��B�Y�m�@ƴ����YB̓u�߉TX<���8|�ϕ�a!=�}b����<�{_�!νS�m���+�ɂ��pgq
�7�O�{�Uhhd&�n�o-7�s6��]���:��3�F����q���<��f��W�H��N�zr�/o�P�u�&c�{}�˟#@�x�����7��wR��t<�:4%9��ktߏ���TB��P�>������7����|7�[%��&p�1Ω��dRej�V��^���9�3F΃.�O;}B����8��߇�xYx����U���`&�s� 3-��X�J����Mk��K����Ct�������e{2��t#|_�
>���a0x���B�zd�ψ�e�oK�7��-F!�(e�/=t���7�X!������Ş�L˴��-�	c�����6?X�
�Vs�U𱒃��-�����Ʋ�*��Ȳ+��	ZS�5&a�l��mᎿ�6��J���A��6m��6��ˌ.����n�4�BA�_A諟+�^i��t��������VGk=\	aQz�Gw���_�3��
z�xE��{�1��*�����B籆eAeЪ�<���zn��=�g��v���},#�
��u�,�� �ӂa3�~v��♒��nm�Jl�2&����yU�������r��~��Y���beVi�᧩�1>���Qt&B}�^!��s ��x2�7A����k]��0�x���8�`�G�f��k�<'�o��[A:A�ǁ	��=q#���a򆫧���<i]܄2�C���S��w|�C���������<ܝ���<
�ʾ��<�yL.��/q~/�M�N�-�Ru��llx�I�M>=||"^�$=�R���N���������/{w~7��o{Ф���]Q��wW%��  �Th@Q��_�|�������}�t�0���3):��d�`n�eIL(?E�{�־�H0͑���,��;U1*w.�~����K�c#��J��F{"���E�Y��U妡���-�w�R�B]�6um:��a[/!p�ZcDsu	����hQ�4��S��޳��R��td>��`m�;��0¬.�ɫެ70E�������֡#[�b[ɖ��a�/cd�%I����K�����sz��>�Sɹb��D:�!���7�G0�:=p�\�����%��)U��b:�3�������Si��UN�t�/`R�i7R͵�E�~���:ǈ�/"��H��m��a�_�Cq�9��ʴA��E��\��(�|&=�_��ݵ�LXgc �f~ƈE���V���
^��g__4���ν�\׳d;od�w�IHps�Ϗ���-@u�v3�.�h����[��Mb9�l}�
X���	Mw��K�9Hr��[v����A!�'���o�23����v�_;-���SPQ,�Kp�L�L��Tel�H��Y����
��� ���f�<ec���_�xQ	'���bei�r��������oo��	yl͵y��=~&ݽ���\�n_'�$��V�`�����uM[���@�����onc�٤z��5Y1X==ݢu�۽��^���|�z1^��=����T�7��'�����e����g�}�1��}���%
� 4�R%�4�4��CHQL���� ��l-�z��=n+�����a��/�֭��k��v��V���[�SX]4�3�\>e���xķ���VW�M�֤�Pz�o�1���N�F���Ϣ���X�'�G2�=Z��'�Y�g��os�^[<%_�9B�xf�u&1���[{��[�z��;�
H��������'3��W��gx\��՝�� �3{@n���Ƚ���+
�&�o�C���ȧ�p*V���x�먩�щ�L�9��W��0S�����<��	��@�):�#"�$�57s�r{�n:a����fTg�~_�������^����e���&wI������g��O����4%\��U�Ù��^�����\N0�G�Ȅ�Sgry���y3����.mfD�����wMƞi�D�+�d"����3L$��,"���mi�#�N��~���ڕ�y��R/K?�oe��'���T�{����F1��c��t����'޼&�j���2����g��˅w�+�<��t8g m��L[�=N5��֙6�b��L�el[�6��IZ�$ZZ�7�ppf����fm�6{����{�>>>�_��g:��O�a��pɽ�=�*"�9W�݅���S���Q'�f���χO��K�N�ev���潿�VG����r۾	��/��t��)�{�"O����k�c�3�Ɗ3��3Z�媈v���E5��q�G{ZL�^�L�St��5���.��'Ȼ�[�^�gV=#"�C�{l����	���y
�Em~lp%�}ӳZ��-��u%ۚ�B�R�}YtJi�#��m��EL��ع�ic.�ZU��g#Yw�ۼ/����}w]�=\�x��kɏ����lfud:�`"i-����'�냞ت�0UBX�ݹ9�))��e��ä
�c��y�I��oW�y�x��3�n��D�c��!��-˯�㜷�e^ּQ���{7}g���z9�û���G��O��s%Y���V�m����xu�����*����̳��<\��zba��v<^z���ke��IkM⦑8Scs���w���g�A9a{�{C`�2֋c��5�4�<����];D���׳��N6�׶�!"��S�K7���{V��1*z��(��w���nzנ�ڎ���o��==�R��l��WAϾrܘ��z�^���*���:����T��{�n�����t]��\�-�t�޷Z{���t����dW�Z{`���7��7(}�"�=��l�n����ɥ��=uK��/�� �=�v��b����;Vo�M<��
ݱ� �ٱ�0!�$�Uj�Q�1z6=`m7�p�|~Z���Hd;2m����L �Y��7*�b $354�ω�ߒó{���ZC�,w�;c��nZ�ݒ��Ay�mM���Guk�]l�]]	���X����*����W���{��s�L;�p9xqY��Ϭs���Vi�&�Q����n+;]����M��P�6[��_X�]�̬1������}��+r���uS�+Z{]X�w"D����v�Za�P�+S�ET�oe����.�����$��N�Nbms���iS�{Zo�y6�����
��p#כ��|�(����k��+�k�/6�JN��l^M��`�Ž����3�.��v�%
��Pon�����۾[�z�9�V��^�O7��]���)X�5PT��u�[Vs;��t!G9znrC����q^� ��K��&�~:*B�J�_!�ݜk��-b��V���u6YԺH�ʤ�\��cX� �{t]5
�6��N�쒕��4�"]�;ơy��݈�aΑ�l�k.�2���ю{o�sܔL�Wh�Q+��X�}/p�bp�c�Y�f�(qP�����j�M�7�=��1�*s}�����y����^��w��D���>�g1�ά��dX��ꯨ��R�X���z�{��W��G�W���Q�Cg�K�\�-pWwS��l���Tp�lRW7��&u$ǯ�ǺP����>4�.�p7�9k�&WH�I$��MU�ß��?:��L��#񏑶<# d����8� aj"1�ZD��x������*����5���E�-h�F�$�l፛g8��+���\|Ж�Ω�m���y��͑ӣE�V�hq�6MEit鍂m��
��ɣ����l޲�95����q��\vF�y��.�<��V�s*^HPi�-f�<ƃ�D~��"�)�|˧��<`�d͈44i��HL�a�� 䛆CC�6؆��J �J�+�:���rJ������TPm�j�� ������E$HҔUC��rKE44R��$�ғ:48&B$)�h��*�<Z��
Ji((��������h��&���Z)����Bh�����x����t{�SEP'�qQ%A6ɤ*�КJiӦ�Z�&�fj
�)* (J))���K�����������a���!L�y��������;�+�"��^�#�u1�#��Sv��v��j�H�c$�}��蚖�������^�!�S:M���C�>'��b�C�_�2O	�p�Yk�����k��Ŷ��P�non̓S`�^�~,pr��ɦ����{cŃϸ������4"�c}@r�e�r��������2�<	1᝽ �L퀹k���lmH�J��瓸hE QvoY����V�"B���<�~4W�V���t=#~��a7�8���"a'V:��8;�{f_9�EeW'�=Saם��r���Sl��#.�-��=sͼ�υ;�."��a =Ų.U��]+/�V��;�˧{���m�H8�fd�T �h(�3�͛e3VP��J�럖h��q���� a3"�M\(#n�>c�
��[�'"���� �[����P%��c=2��Օ[�[(��-�B����ཋDb�fHT�8�(LJv��:ū&=?B�오�֚�j�0�]f4\6�d�y{�w������) �?p���Q��Z
x���Х���v��.�;!70�	�{󘕞����b�̲\�6j�\&7u�[�r��Cj��]�:m��ȶ�э�DcO��H8v!��n\�ӹ�C�<�T9n��(�^K���Y5�������J�\i	9��I���h���(ʘ�/�{Ӊ~��`^���'�{`�O�� ^n ���q���@J�3�sW�=��{']���x)7�R���[=�Q.�i���}��֒����ԇ��Џ%1�H O�*4�!H�O>y�������I�ϼ�b��E'��-�Yp�� a��!#a�O�&�L���WQw�w����ݺ�4�9uCHӮ.�{�6��,�1�i�������z�3�ˇ������qg�0D,1����
�CYt%������@��,r�'�I䱎[N�B�ݛq��i0�˟"Re��;/u���Յ�|������u@άYB͘��.�TXRΞeV�����m[�f0�g�Aڱ��\8ˇ�C [`�L	� n�n�ʅ�(X��Z������m>��uooʏC���~�b�g�?�^}D\�Q�`�ZrN˲��m��J���	K8-42�����r;�]�Άi�f�O@��^�90!އ�����߲a�'J�69$�II�|��s9;V��a������1נL˴�������[9|חx�΋��~�oN�kǩ�0wyߌk�M�7wt��h<P�C�Pi�&a��D[*��xc[�j'���pר��'y��y������|�B��z���T�A!အ}��B��4�m:m G��=�{��hEw�LF��:�mgm�Ɨj�08�p�Rd��].��q5);[}jw�پx痪�kV�%�����x�s�����Ǐ��f�g��B���uY�iǗ�M�:
�A�*�Ռ]�M���َee���;.��!�0��}���O�� $V��>|������gڿ���S ���02.:.���Q�]�0�عH\�0���B���nv��۩S�������:��a>���46)��-�c�i���1N2W;R���D��R�9�<�T�ޘ����:�W���'��=�-��h`���o�����C���C�	�cn}��+��ƆlR�{�|����*�?,P/_���2�2)z6o��վ;ć��6��6֋5.��0�Kod�&D���1д�:{Ot�N��K$���PH�aO�|��s	�2蠏W&�~)��1t%��?1?U{��|�ˁ��{��I���(�av���]���MCux�>�v�
Df��P��il�˼�:FխA�Ӊ�s/W�T��1B9���	�{
7�4��W��]/e�?7��#Yq-L����B*+y�j�F�z�K��q��#�M��[��SEՍ7Z���r<u��%Q�de���ޘ�R�K�F��1��8�+�t=��%��Ƿ 8��o�`�_�.�m�ZY,�=f����-͓y:b�eK+����QE�^�Go��C7mŰ~����qà9����@��;�T�����Ծ��6K�q�Q��!/�G�Yץ�oe�4�Y�2��n�nӃ�/����qq�`u�L� ���_�Z{<	��1�)ob�v��_Sw�x59�b�!�/vܢ'V%�� �����U��������9,T�P��+�S[��|=�� �'5�Y�$;��S��fۮ
���(�|�LC5����j�r��a����v���x�k��1�BcBF��jއ���#0�2'�ӊ�x��g����}b���DS��U���yݞ{2k��r[#9����*P������gx��f�Yƃ�ݬ`�=�K���"�.j�u�1q �񖎮x�\%��"��D�ǸG4���ZD=�O]Qx�s��5�p�4h����*x���ګ���ˣ�EnawO/L����y���yg�,Aii(M FFS���G���&m�m���c�ts!��Z��}~�ؤ�j9Ql!��6�5INP|ؤ�1��t�w�`qma�p��eGAPy�kOqf&{���^���%6_��5ya�Oj��
=�V�o�[�xfL�:C�~�=�ػ�΄Xjx?v���(�5?Bo2p��"�3L�*T����ۚ���L��gnj�k�wh,�^B�ȝvl�1���y��
e�1<�>9�N�ˤS"���~��t<9����ر�r�~�����qC5��Rʹ&82��v�R;$É�I>9�NU��h�vHkn���� g���E�#��L��^��}�X8�ID>Ǚ�jX
�=�-�V�<��P|R��C�Oql���T�WWi"��p+52����<;7�e�!Gۓݻrq��W���J���	b�_����A��:d�������|	�n�vh�g������W�x
E���}�������� !� (P�P 0a���^V�J��u��f�wL�� Laz�������D&��a<���c�ˌ���7�0q�o��<���ǫ�KT��/�)�./#�#4�|@~��~`�ZD9�F�2�;�i�H'"�_Srר��@sU��j��&�G��:J;^�e�����f1��6H`��ik�45�g�>�^������ʡ\�}R)�z	�kX�2m��)5͖Ż�l�0j�k%�V�����u���������^�����i�j��Sxqg�X�ǧ��$�sW���
hy�Ȁ�n8�����k��Z����LX	��^��3y6�i��@��	��C���zr�^�9f�U���YU��qC��@��_��.Q�<}\//�'f�D�� �%o;E�GM�k�P�z׽[Ƌ���v����E���o`C��h��xt�gT�m�y�A�;uC)�*��Y���p���T���n*n<�5r2�>�֞�<����{	��c�Yմ�i�dV�8x7J��y��O.جj��0�&��Pj(�3�͛eY����s��$�n6Yu����Y��-��+0a�^˧�I.*��R�`�3���Q~�y�����}鹡���wܫ~$u����Ѿ����������s��G�0Q�^�4�}�\8�p+v�Mv��<X�S��_��3�=� ���ɜ���5]T�yeJ���P���$B	B�@"D*( "��߮w������ß�������a3�)l�U�.��X�ބеX��l�c��H�m�^��*�&��u3��P����,D�LO;N��M��_�Z�	�N�i�I�g����H�gɓ�H�ƢÙ^\�t�C�p�� ��A�k����ے���]���0���.tKL��ۗ�h��\��&���IſE0��к1���i�H@�/���.��9���.�;ml���)e*��<��	O�K��,���0����i�'陳.�.{��4�c�J6ըX�A�8��݆a������6Ⱥ�7 ��e��Msӿ3�ˇ�c�}���"c��	������S�C�l/��F�i0�9+�X�Dy(�	IcC�ӰL����;0i����u����͞c�s� &)��/�nE0�N8�J�gO2�
�XT��j0t`W5ۨu4�2��\�t>�H[�D	�Lm��Bպ��|�!�V��o�<��lhzliE�j~�]~��zꪪh�K�xӛ!�xp�38C���}N�Ӳ�v������y�b��������k��8����q�y玶����`5���f�=��:�=��{}8L�f��u?�;��h�<��x<=��x>�eOj:w�5 /��L��7}8�ye�&���7�����j��x���519}���ouƨ��+������?�}��}J�P�� 4�4�" 
R��'�?;���>�ޟ�|����5�`���>W�Է5�,�1��תD��.5�B`��oJ�Nq/��s�o���y3]9H���a^&$�Q2�u虗iD[�}(yw^.#a��/շV2�j��iЇ�|a^ٹ�K;��@�oW��{���t=D�6x�e���i�C��O�BkOu}Y�ߐf^C L߄f�|� ��U�m~��>̂C�P���P�My����v��)z��j����y���!s����Ô�b�h��F5u�T�� �H\��e�{+Y�U0�k\��<j�!�z��={zm���:��g�!64��,����%s�-��[ָE\�te����]��5��AcK
OaQ�z/q��E=����Đ�B`$�̭�]��X��7tv�Pdl�W��)���)̈́��MJJ�v#f��_q�=|w�	�knx��iv
�Դ:�u�H�p>)�c�Gc@#�ϳ�e'XĲN��)�y#I|G����h�C�8��=��՘��iZ�K�k���xn�ñ�J�vQ��y.�#0Q�-�L�����-�â۲�]P���]ڌQ=rn�{�yi킳��Fe��M�=�ɇ����?������������!!ng&��
��<�������!�-�)��|�"�v��&�v�Oˢ���iu^��}��e�E�Z].���JgmI��y{��I����A?��,B��L*+@!B��L�D�"-���=����;���;����~������Hp���fƑ�$��0�D��I�U��^�I��Z祪n*6r.��훬4ܼNæ��\<���=�d��p�n�;4]�`[F>�����!����L���{���r~�}�>���K sH��Ƿ 8�H^�'��������s{�E��N�ou3��_�讉˘���Z�t-~A/r�J9��K6�	�"�����B��X7��ı�}왑���k"щ��>;��ئ�\I���u>X&}8�8��Q�c^1a����A�K*�seZ\+#q����t�טy���6�����=���1x���H�w~���<��z��j��}a]j��7����p]�
%�,9a���Y|ڌ�K��'v����w��z$@#�j�]�mMw|����w=���'!��vi�}�>�ɂ��KHd�{d������um�2���32�{�3n�S�N\��ʘr�t|�,)�of��<��O������҂��No�S����Ή�֦V�-C��|�9=����lX�V��&+�C�fͧ��V����,:/~a�<�}yg��{��Ȩ]N�nl�w�3c �UCU��w4���d�M]3Ǧ�����9s��#�`zg�?=SL+<��{t�o[�����Ӳ� �#~��n��IYc"[���/�i����g���#�P�M�f:`��W|�h�b\:q��3�����OT�"<Ɯ�QH�}���D�T((B�TZ�B�i)T�D�%�=�� r���ɵ�C�W�G�MklN�z@�"S����a�O~Tg[��=�L�Gx�;�N�Œ^�{=�&v$;:�[5�\�1!�0D!��zF�*���Ђq@��E�#4���Rk����;NCQ��D�E�+�{���k���d�Jvl�L[@#���A�%:O�s�Sud��2J��=^u���[YF\�6=C���
��(fܘ��{%�)�;��O"�ȣU���s������9ȗ%x1�]Gh��c��y�|�-� �z�	��86�ܞj/usFa�=�E��9oܶ/z������	E�匤�������	�?H��y��^z���0`��83��ڕ�!��|��m��֤�Qy��F������-g<;��1��!�a=O�����K&�����F�p�L\����֙0q�4�-�*�f����ʲ��fF�����^�gg>Lf�6}B����@g�jߌ�P�#�V�@L:�x�Z�z=;�b���얡�w��I�&C�d;�-��3ǐ�ŧ���^��{�.�����NF%��������<��=��h<�=����g��)A��ۃc��f��)���zm�3�e��rejJ�c�'Oj�[�@�C��\��-����[�I�{�3L�rM3)aΨL^���͘cʳ��s��F�u+�M,�gt�A�7/�3�L[ޅ���w1��|?�}� D�̍"�(Ћ@�J�B�-"�*7�=Z�ER~�Є��Ȥ�9�[����s�>��>��
O�b���H�J��?9����g:�{шB�)�v@ñm�.�N����<�����j��CE�i���e����n6�t��ܾqF�Y��ռ�e�EO�,�4`�]���A�z�?����a�7��h�8��b��32"��H��`�|����1>���V��o�� �ˠɹ+��(�/<^��]dgN�����Q[8c*w��;�:���>��zaS7 �r*ڗA	���	ͨƼQ�g7��L���l�[�/yzd.���\g@��"S��LO;j�dۓ���Z�LRu��bU757j貜;�L�����K�U�)�ۜj�TO��^����0&������v�=�;%76��tBh�v˴��pY�T�n�D��(еaU$��:m���-�WN7�A��qp�2{�NL͆�f���s��C|��n2��;��x�LU�H���@��/��o,�r ��9uK m��Vªo�	"qNT��^Nv"�Y�P�,Ԯy��m�t�ny�i�}������/�����������~�_������������������Ǹ��t>�I�p����'oj/�y�����bI�׳�}�vh@|�� �iY<�%XF�!b�JoV�17�_A�^�F.�Z;Mն�Z�J���ͦ�5�wwy��]6VL�V����]Txȩ��s/��u�1L|�S����:E��7�[@����&�a�[hn�K��ܧi���oqT&i�TD��oW�*��%��5&oO�6*�]��0����F��C����y����x��;���R��}�z�|����jՃ��9�%�;_�N�!������c��{���6�F�H�E}�^�]C�1|���2Z� �ˣ�w	VXWz�dm�T�j��w#p�%G�Q|�ˇ�ʌ�����;���v_P=���i�w���O�����>�k���u���������O���O
�A�/�\}�^x��[5��q^ͽ���*�ugu삆�d<��uqe2��x�Dr�&��D`M�'.�zqB�EP!Y3��}�zju;�Qn`���m��ڟ�(z�d��9T��+�^]��B㴿-����?E?]�-�����PU�H�N���¹\o�3ga,<�p�땜#�Pշ��1�F���ا`���N��B��[<�_!p���%*��<	�O�ύ��x_t6_�amI�� �vQI�u��!�7ڰjǦ�7���8p�+���TENE�ݪuW��6ò6�(j��u��}J��r�v딯���c�:����:dV���Ե�����'�A��c=W�󛡉�\�\���y��vN�({Ϡ��/b�C����^�E�j=��E�wL1j��WL���)�֩u��e2y�{���r��s��o}yt�
_y�5���ねC���i�	8tʻ�O6]�v���c:��Yhj��0rE�`�S�P��'d�1�euw�~���2���w�d{�7�G��N��+����b��ǐU��2��U��Y��}���a��CE>���6����_��4mR�C���9*n{���Gj��̕[�z�3�Vv�zn�,1Ǻ-݇g�4���
�_l��24S4b��cj�1�ɲc	Ǟ�Ϥ���N�w�9�ճ�7���Gʯ9{�7ڵ8�=�e�	;#��ʿ�J��n��z��2�J�8��s�u�*������5���v�^`�.�TrRj���j�X�k��ʋbmzC�-�K Ux�S��{�8ϓO9��Ÿ7�oP�!x��]�Kdʳpƒ�S�j�Eb	��{LI'F�>�ݽ0j�����y����L��mhK���b�����c��fs���V:������/k��SV��0v=�3�������Û��w�M���k���
Ã���t�����.�V�i�A�w�g4-��J"��xS��k�W�r�o����A����ӂ����'	s��&�7ݳZډ9.��q����Zݬ�<��v���n�0�:["�$���o?q��K��0KS��AA��T�mC�A͊�*�Z��������[��KUT�)G�E&��a|M@L�HU40JP�Dh�CPTP����{ P�ƪO0b奫��LE	3G���dӧE�QE�it�"
�IC�(#dM/9�3!Hh5BPP��%(r}|�<MR�z��ri�j�
H��褣l�P!�I�M4����'&�����*�Ӡ�)J]�V-i|[�B�)� 8E!@�AC@�^���J(��R���JJ
Ŧ�cBz���|�!1(PP>�E�dy'%<�����)
��G=���ݼ�=z����/��>��?^<�f��j�dj�{[C����7MB��.´�������}}��s�ߞ��w�|�����d��H��f��
V�h�	�	��=��~wǟ�?z�~��q�ݴ7s伧��4(���{�%s�W�\��iIc�e�N�3�B�N�U49�}{$g+wf�w�N7y�u��[����5�,���+|J�ΞeY�n�3�+5��I�Y���P��p*�3���B�[��[�`(Lk�R9��MV�V��z��R�Lm=��26��ǯzS��)�~۔0zp�[�<	���T|�ϬNjv]���r��'�\�-{��
�@aڡ��ԍa�Mk�L�Fq�nc�(��{�`�hȗx�`<�66�I<��gT���,��}���o�z]�|w(��LIv�L�zK��j:#���_Z�'#6��.�ÇX�G+�Z���xBC�9��ºnu��;��G�dZ�x�� ��8A�0�C�,�B|d�V��K��}�nW/R��;G�(#�Zq>��c$�꨼{k��9�Hxj���W!�U}W�B�в&��I����Y�̪2�D�5Q�<�+���0}p�2'��D������B���,�n���7nq�ܑ���p��6�����>!	��C�v�֢� y�3s���۾��C�֬�=��㿧����´7�dD�Rc�D.�E�Ʈ��+QÓ+x��+�f�{��õ���{1	fCa�{qnK���M�B�+��A�~��L<c�-v);�.�Hu�LEx�5Tč;i�N]K�޷:Eu���[z�����P$�E
D�C0R�0AB3
�"R��Q@�3{��&�z�eq�i�� �M��Be@,4)_����.�Nk�M<5�S�;B-�'C�֭�q��W�Ѽ.y��׸4���5?)���JsiI`�AR)�+�e�������n��'���ǿ=1a�ff�`���j`�#�� _�锝ax�E��\4�/X�8\qaŢ���p��{��I��'-6�DB`y�\���i���<�EL,#R���n�d�l��^�3�I��䇿��|&��8`���{��k?���У~i;����}OF�7��U궉�3�4��4��Y	�u"��_���K��p�~#�6����S�E՚�`[t��@��)�7N]�j�ޘC��J^�Gs�mf�e��Z�K�ך'r��u��3��v�Ƹo��Y��u�e�q-X�V���%V�&=ұ��+�E�J߼�*���U�
0KG��K�T�ddt%H�G��yЇl|i������6���p�1�Qt�dϧ���Q�cF,3���"
���ʆ����Ԏ� ̇��by����_e�?p͐����ID�h1^>a����#jH�����&-U=f�w嗣���#�'&x��t�C�+�f����?���_<)p��q!�ߘ[�K�{Kǉ���Z�ݎګw�����v����/E�`��xN_u!w,q���8ǎp�#��c綵�<�-���+�]���ߛ���o�x<x���ZY�R��Q�
)I$X%ZUf���ު��gl�P��+b�Aݯ�:%�8:ap�N*&���Q��g��s>ݬ`����Ffh��w�m��]����HC3*[E?�lEC�ȖxBK!�[=�O�x�{8;�kv��|�)�z˓5�u�E&h@�,:��#��5O��](?��V\^?��_��ߘ�;��ǫ����ks�zw����E2�)S7X�(2�Z�`��rsf��M<,�h�_~���л�j���r��&����t�W�w!)��A��i=�Fu��Nk߱��CF:�6�m����t���X�p<7���A�i�P*���ЂpK�%�B3L�*T����"�NJű[�/yl�w�c�?<��H02|�S�eL
GcH#�>��%:N��:1p-7\}$:�o�\��;\��s�O�`C�q �5��JZ��/���y.�Od�q8��v�t�Y77ss���Ϻ�)F:u���%r�,9�c��y�XE�����	���>�?�8b-ڶk׮������#��>!7K��?"�A.��ᮙٍ[������k�8�WV�0��&nS=�nM�/$8���W�s'��~����'��l{,w���6H;5mJ�>�������r}W��_h8�E����wZ��d�ݪ��17�\���z����uZN���Y9-��3]<����5���E}S��ġg{T�c�}�
�b�V�%��J�R�D�X�Ͼ��w�ߏ�o}�������{Y4��i�k�vQy��F�yT_�*�W�DL��4ʣB�R�-`�X+ϓB��A�Yu����ά�Lh&����)?5�i�oV�W�J��m���V���^��1U���#;�JŇ-~ivnu������"����E�Yk�����P�e���{{5Z��+��&�4�bF��T��:��}��hv�.Vڨ�Ԫ�&�6���L�~mz�s�NX�qß=/4G3�hQ�"&9��#Y%�ݲ�W�Ռ�Ef^[����jN�vЊ���\eش�0]���/\�o�D�ǐq�q�s����T���.9	"�;�n*�b���Rʹ;��b�����M�I��x5�)�WLoULU����l����BE����|��u��^퉶�j+֡L�B��8�Y���W)���@�!XG=����;Ŏ��v�ya�7 ��VԺO���NE���Ng��,;��/��ǧyk:o�C*.и����\f	��i�Y5d��nt�H�g����ܿ�LL�����0 !���}M���Ӈk���W�s��K;�Υ#�F$iv�:�*��EmC%��A^��NڣW>;�qX(.x�޾��wuO���c>�[�O&���J��7�#���	�r]�S)-?~s�χ��=������%H��|��<�<��p�6ۼ��t�L)�m�5uEë|g�[��3]�a'i�����w!��ȡUi��k��r��A�9`轺�N�S>j�RK�3%N0Z�Ѹ ���H"1�C�tn5�N���>gN�L�حK��1�&S�0�Bb���O@b�@��avm��/ =v
�ɶ*��CN���?u^���,k��4�T��c��"���ˋ���}��h<�J��I����[ʚ5�p�hq���w=	y/��hQ���U��,r�'�	IcLVt�͏a����9���8�5V��
U��q�W��j/���W�YB̀bN��%Qaq7�^i_f�"�uNgS)ͅ�ԇ]��D<A�ȡG�.�
Ԭ�ǯ�{f����i�j4����U�ym��/՜�\��u�����Q�P�l��|:��1�k�����A�^:�Uc����'��N�Hr�a�@J��]5�K�E�Է5x�e���3�끀�8��v��X�̓��pE�v�~ږm.�����w(��bK�,�\��l:"��g/�a���S�C��k(NGK��Ϫ���a���n�Nk�K��zvb����:w8F�����W�ygpr��H��<&�ǦN'������Q��7i�8	w��N�7yE;b����~�1���w+�N����s��m��\���>��|ޓ;?� ?� ���B��{��ى�QZ����@���^a�0����2=r�;2,����!��2&!����I�hvY*�<�pJ����o`38��%��fJO2��M�v1�2	B�/�H��o)��g���/��i d��~?��|4�>�?��P���1e���pڟ�-�6F(����1���Lz]��м�/xb��Yt(��3;Όu����c ��_����~�t>�4J�i9��Oq���*U,Z���,�	�,4)=�Gh]�ǧ5���S�;B-��m�ɫP�3�,����j����'{\_�l3����6^%9����2kT����x����u��㏆ٚy��[7SB�rs/[�� �����|k��2���x�E���S(�$m0N�l�6y�%���$�Υ2�9���5��HP͒B`��n�h��Ñ�]0��J.�8�y�Z0�5�f뜜X܎�C*�NZ��kǜ=O�PP͌�6g�n�2$ٔ�&��.bXЧ��[�{NUwF+�Bz,�1NX��a��?��+ܯ�w��Q��x<[���>s������C;��Vr���0�nz��/UY��7��٦x�=�qo?e5���۳z�>�����W~O"�~ʖ�e8����|��w��s����ރ��g1ZT�%ã��y�������ט3�y�׹W�fГ����˱�������1�xO���}��>�ẅ́�.����f��aM�4���{O��UH�sn5��á��!ï��>wV,��cWUPsi�cp���ʚn�����%Z�Z�9/R�m��nb��}@�
��?D���_�4�n�BK���?���P��j�4tXjl�r�1,��Ta1����ǮY�ntKeN��/�r��Z�B�����v�:3�7���S�<��{چO�l�m��(�A� �+����h�3��/��wu�V�*�ōp��x!���ĩ��6�5��4�ݬ`�/�c���4ܗ�Y����"����O�P�^ȖxAid1�;S$���g9w�c(�>�(��%�.T���<
�R2a�ϯf���xmhg��->ABf��y(��YϱJb���]ϊ�}%���6�J�m�2�*������6�i�t	wln�{���.L�M���!�>�5���y��I'ks�^��%6_��5,3I�ʌ�
�����h�mLQټ�Z�x���Ƕcqk�"X\�Cέ�E{%W5y�N+���E�#4����z~������z�k�T/Y��/��|v��m5?�����{�{O-fF��}��7ǎE���yӀ���w�'#�a7�04�f\#���loDl~�O�����6soa�l�(+|W#oO_d�_�ͣ&��|�M��ɝ���L�6Ewn}�ުe{8���[>��|j�=���[��A���]�*a0]� ��d�z~�N��՜Ѳr�����z�k^�p��|��2)��Jjn���>Eê�G�f��!)f���S��v����q�j�kG�/�\8^�]H�:�Nw�@g��2���j�1��>G�e�[Pr!6��s���N���Zb�Ki�&ڵXlX�5��K��M���1i�c)�./#�#4������ܨ�u�c=MX:����_È�]�p���jw���]����5�����3����Q���wUSj�,mf�Xm��q~k�P쟏L��[�7B��X�~&R~e�=J�-���U#j!��h��]�����d�v�����x��7�C��/C��hv���%0��Yk�socC�΍��u�W��P���I�6G��wn�����P�ŧ���^��2}�v��L4�V��ع5uq��)�y��a@� �{�W5�nZ��w9�4G3�{�����N�V�@j�cr�\��j'�?:��`���G�ش�0]����NC�<����h8��0�;{/�!ڧ!4c$d1�b*:�^��^W�z�%J-˝�V��Hvol�9'������}2�^+Z�몦5}l'tsw\_CZ~�������tZ=�S�V���v�9�W�R/NH�-`���6�w���$��|[��m���T�<�+���	-C����c��j1����}���+�Iv�T� ��F]�U��lOc�q��(��..y��PY]��34����a����ܞ�Uϫ�۱X��P�qB� ɒ�A��~��g|\����O�Q��`T�6��$�s���L*f�br*ڂ�!>��0�w��=�P��Ji�ܷ����:�%�`��'V"K��1<�>�Y6C�s�険7�^��^c��X��j�CTQ}��Ф�S	mw�Z�����H�oB�,�ީt��թr6���nMD�s.���Aj�n^{�(�I��bS�	�*��]�M��ȶ�޶����C�lq��]P�e��^�FÅ��}�.�4�t�Ou*L���Xn�I�.4�3����-�v��;�Ҩ;�MI�����!!B9��s�L9�v@�]�a��
yC��"�ܷ�F�|���fm]m^R��k�7.��3���88Z��7s��?W�Q�F���«�%s��I��B�S�q}[Y�b�4�Eb��$Xh~�&��Q�*�
�3�7���tf�Q�u��z�)߶x�O.����9���B�[�-�%�����G��7iG}�;��:U{���Y�Ä���)mf���SS�qnkV{�y%2Hvy���$$Ic{�l�6]��bo����-����	�腰���jMe�}�<K��������O_Lzj���[�Ki*��U�n�����}�e1�����a��sۇ��CsO�[��Lk�R9���L����7�]�!&;5h?J�
���{�PK�Z��z��W=�~��?�3���ikY�[1��kh�Y,tf�8���t?)�v&�v�j:�a�Mk�&�+�KsP/�ae���d"]�Y,S�<tR��,]�;� �!��e�Ɇd]�o;�ܒ�@&$�P&Y��2�%���m9|Ϩx��uY{�����?�\�;��|�d�'��s���f3"��wH$9Nb.�/p��N�S�ξjz=�z���m���`38��Je�Fd��*���n�4�A!��GV���R�knWnr�ν��<�)#^iN���`�x3�XH��8�˖�d_���B��j4�B��={�+9SK$zB���2>Yt(�Q�����W�b��tS<!	���d�p���3��j/)p��7]����~�-�O�Jlr\HL�t�.���.��s^���i흵�5�xa����U�
8�8�}�G\���_)��%1�ħ)A`��)*���[����=}?�~�z�~�_������z�~������K��,�;��_ʙ��a�~�vw�t>��;{uڭ��Rж�y����^�o�wu��"x���Y�����믜\紟>2���"��{^���5+�pK3�q9��^%��L�B�������;�hl��s��)&a��9���㕒u�[!�����:d�6��=�ؗ�lɻӳ�e.*7����ؓ+i
'�.j{I{���cN�sЖ�]�m��N`BU���CZP���a~K��E���}��F�n[�2 ��/y�`�g����9�Қ�y�ũ�:,�M��-{����-^~Zȃ���<�9���o�}��=^cQĎ��2���u�鲝��X(�`�Dպ�RX�f������C�mH(��6�(-4�o�7��G�Ǔ8�vU���wkX��w�a>z����#��`^��g�X^�9�v-([�Q��D�iX�[Kd�l�k�<1����LX�n����h��cr���u�� �sFQY|�-��� [��5{�fn𳟽��1up��~���-���냢"�����(S]��^v��Ve�	�mv�O[�D�=a��f�\�����DUA#Y�;E�h�cbI'�������M�{��{\
�ق�]nz_s��٧{i����s�� ,OY�t�3���ޢ��J���
86uvVB���m��W9[W�3�<u�xᜢ��So��wP� 2�H�g;wF�_A�.��ە�g�ݞ������K�𾧭��7�鵻Ԋ�i�h Rw���ݥ�eAek��e�=�	3����~�|���ߨ�+α��ӽ��}鯈~�y�;���RX�r�uj�?G��/>��*āe���h����#�u��+Ɛ�k6�:gwLy~�{���ң��9�����C���t��^�%>�i�G���,׳2m݆��3z��������1��o˞�M_Zꌝ#U90_���!;"݉}�@�[��,C���}��BF���#��p�.�����]8T���K�9w(�U�`�t��=�|�҂&��:�=w�Ƿ"�y1��4�͢�G@�(i;cIH�A<������.�i�64�a^>}�,��v���m��MW]b���=��*�;e<ǰ��� 1fz�2'��r�]2�{�U�����,#�B���aRޞj�Wa��w<cQha��)�#wu{��Zv��`��5�%��p=�efH�I��}_K�ޱn���ܬ^��=��W\O=����O0hB�W>?ub>V7t��Y).�GY�|��6����&�A3|j�K�x����\t\̠lg���Ƿ�[�]C9M�(F�+��P�^��>L =�aD��2\�h� ��@�ݷZ�%b^']�&��˨����ٍr<��j�>ɗ�d�������3�啰{�j��QtC�WsΝ�87;��n�k��A!�$˼:=�w�l�����{͔2�'������e��_�%<%Q`����٘|�Q�'���(���!�9#�&����5��?!@�ATIK!4��p�P��("Z(
B%QmJ��AB{�4��HP-%�%%A�RH�� P�>\�Bi����
JJh)�R���P�((2&���J hV��^Z��R:P�&��4��i�B�����/ 4+�R�O�����JR�t��ޟ��<�{����O^wxy�{��{B����{,*�"�Vh|���=3f�ͦ�w��9,L!lIf��p����ٗ{Q]�w.�١��j��� ^fġ����*2l
?�=����oV#��0O#��|g��	9@�K"�tS,��*D
DM�,�~뽎2��^���.a=s�@�a�$DO�������;ncH�^@�AlR}`��(��oO&A�'�n���$��r%�c�t�7q�NY�6�Y���!7P7H�4(�e�q���,��V�9j4��֢��ZPX�_��Z�C����u0t��#[�2��DS��d?y�����/~�`�F^���s7�t;��@����us8m�"��s��A6����w����0�;S����ْ��J��ҵ�%�^S�h7R͵�l��]�x����&0�? �����bwfN�ǣ!�q�:)�AT��(�|�gӏ^�3̵a���/@��XKSԌ�Lܽ�a��z3���D"�:�_e�?p���~���/p���Cm6�����KtͰf�
����=�PxO\D~y������`��9J�/{Q��gJ�S�1.��6��fL��z�
���v�����	3[?��a�q�KGy���2H��c����Ycpd��s��5(f������v��ZL�3�"�>s)c��4V���E
B�z~����JA�ڎ�'j`�������n�=���XH~�DŁ����*��m��p��{1����uy��3.���ZD�_r�zm�S�2�n����5������>�]E6w��������7p�4P�X*�!Hɇ{�9��Z�?40���*[Fd���(r�B22�X��^�{�t�7jRͼ0��E6��qKh=�7�X�oph�
3+=U_v��InO��O���W��f.=*�&��V=;��!5�1d��'�Fu��l/#S<e�b���+{���H�^���@��.�@D<�[^�E��\��A8�bY��	cV�4NRֳ'���m l��R�G[�P�r�َ�������S�d?0Y�� ݒy���v]��c�sݛ/���ڵ����D�6�E2)Jjn�u�5ȸu]@0�m>���a�2Ùo�g�����CZ�aāƕ$�����+�[E�1/e��Ϛ-��\d��w��L��$��
��&81��%�=�*]���/��? ��;�O)A�^jF�������ܪy���밭���gl�{f%�=���n�ګ���e�Y#YK�����3�B����N8]�Uss����?S�|vc�X8sȇb�zdO?�jE1�&����'�Z`��yǚ�ó"�.���aFg�t(��p���νh�-������3-���'�c/�`�Cu����Iu�-v"P"t����+"bė���S�y�Oߞ��y��Z89n�<��ĨK�:�bb���
����Q��7V-���'�L���;�O>K�7�������2+c�\/d�3W�"�ٔ���CG��&��,��P���"��Y��:��O[�͵�jX��R�޸ٗ�?�g�V�4�jpwB�F�-1gml/�P��H��i�5�6���Z�ގ�A���°��0� ��+��
r�sтs;=
��mOvݕ�e��>��w�\}�z�%i������6"�L�v�q�b���:��<����%ާ�n�k�\������&�sB�cH1�́�8�n��}ٖi�+�Iv�6�5r2�m�I�础���d��ۊ�L�+����w�0(��ű/uW>���X؝ �E�A�P�Mm�R^
�?���ϯ�7���^tzf�Ta_��ƒ�P2pBN����nA+�l�5z�O��9���TY�ց��]x��R����g/���hʋ�5p��X�.2�1<�#T�&a�6��F�|��|�Ƶ{��3�[��e���:�-yL�a,�ۜn��uOl�T�ސ��6W6�=J:3;�SNU�����t;h^�����v/	�bF�+�I�tt�	�m
�N7��=�)��m5�&��)E�w��{��3��vr�����u����p����ah����r�.�Y��}�yV�>��~���������?g	��T�%��$޽�:q��Ӫ�{R��E�u�b��c�o<��v9�՜���y:�r��3`א���>�3�D1�ѿ&��8v����.�����*Sx	��7H��\h�8_�1�5W5a�)�����I�А��1j��?�����q���?�o�H	��Ͳ.��i���յ�^��j�a~Ⱥ�����Ȟvmg�`�� �kȇ!���/)��Q�F��aTrW<�;l�i:o%��"�wO&��\^�&S�����vm�|v����!7T@Lm�^yրk(YO9��<pr����=ڪ\r�&V�-Uj�X�}iZAa�B�)��@���ǯ�zb�l��0�N��9CE�k��cR�,�0ޕ�:�_�k�P/mj��N�\��{�=���h���(WB�&
���q�^����;.ݵ��,9��Y�<�f��f��5-� ���|�+��f(�D�c�M���;�`���n�ʥ��V��t��Q`K�v�L�rb����:��_P�*��;����/�r:�8������W�����y��(��� ����3=���]Wki���$5��2��eC�m�����2eĈ̔��T^=���5�j�C�ҡlB��9�~��ʆ����k��~��6<��Q?~U��5�:��{����&�~k�x�Ob��̋���+mx�z��>���{(Ɵ�����jޥK�¼�M M8c��,�G˔��T�<��id�wK�&Pft'��UZ��X��z���7g��ۑ欋!&3�ϾǑ{k��n��8�}�[�R��W!
Dך�e�g�b���g�`���$��K��݈}��c��+�6�ռ�����57q�u�A��L$IҨ��,obY��Bmi�WQ�M�N�+E�i����C��m����ږ�����&Bd�Ȕ����z@�z�=[�uĒa݂^Z�$+b���c�������"�<�<���6ħ6��5)*���O)���N�!Ok��9��M��ჩC�CI_0�$=���^m��^�ْ\�c���«ˢ��!C����M���Z�ۯ�a�?_,��xpߞ~@i?�?�P!��D�����,kl�=O�s{t�=�^�R�[lg�͏��U���;�ׇM� ��Z�p��&98�SV�cRZ�\�h羍~݄2��;����^������Ƽ�L?5�]���:mi9��2n�
&Y��-��!95��1LhNл�2�-Gs��t;���4�����'��P�&�y�ݍ�.`W��#�q͍���~����S�$x���c��/)���K6ǜz�1�����r{�ǸS�[=Pw8b��;n����j��]�&w2�c�������hܧ����q�O����n��{&��	m�p�� ̞O/ޛ��gL!wk�z�0Ѻ�lb�y3��[6uB6� ��GNu� �ɞ���Uzj'Ή��!�ه�ܛ���|��QA�0y����:!�C��i����Λe~��1�TI��J}:��g^y�Z	v�G�j�c]� ��Ia6����;�c�:{u���lE��`>�Cg�'�἗_mv5j���E֑v�Q^��+Y���\؇c��������f�[�մ@�z[W��{ә�=!ʹ���C׉�MC�O�P�YϞ�!%��!���v�"�H��lP&��qw�-m�C�/��;�kH��L�W�`h���0a��oM��X�xi��iռ��ʖ��s͛'���DdkO�#)��T�Sׯfm�jJ����A���	���fͧxi�ZUQ���{��H?�a��=�]�0���Ϣ����U��y��D��&Pd�h�'W�9���� d��^Lf�;�XU�[�z���-��8���
{�bN8�lL�h��(�e�9)3޲�g��M��f��R����۹�<����	J�.͐��ƐFNWk�\�<����O]ƭӨ�t_D�V�|)���:��������<�����m8��h띂���l��hz^����Sag�\3ޏdb��y��g��a�=�a\癷�y�Q+�jcZ�?ߢ�����t�+e&c����Kz	����
�{y紽���� g�L
<z���7���N*NOht�16�>�V�;yuJY� �s���m�vx��}a��;��L8�)?9�NVy�E*[E�5 Lav����a�g�c��޵��/G������"���27$�¡ۼrt�1i�`e ���#��bͤ]�&-}��ݍCk���/�PV�п��/+�<&�_qr~�T}�8��[#�K֨�~���qE9�@\���Э�qg�%ݣ ����c�ƃ%�vNUx�?����Ơ�ƻ�'���<�dkqe�7U�]�J��8�S6��vn�����?0���;k��T7>׻MWy�e"��^O:��,
��u쮟W\���A�=B�v��73������֦Ǹl������9�MoHr���% �#4qy���-���,s�<��cX��q<�,�\��Jb{_��i�s/�+ߛ�8=�hEx���C�����:��<��`հ�ك��OSx*V�� ��0|�X�昘���[m:��>��4��K�)�� �9v�]�8N�]�j����z*��zh����P|`��Ⱦ�����7k}�,�[|��7Y�{.��vM�CK��3�!�۶�7�C�ڽEB|�ɕY6��r'��Fr�֫:����$����I�-�c7v�&Q�z���^�[gIj����'��������-�=��"�^�/V��>��eRt�g�\�����y{;��\����j��|p�p���!'�C�=0�3r	�9m�������|˸Yw���b�Ol��/B�	cE�r�Om���K����A@��\e	��mn,	matɞ�ʈn���[��fr��^S�NaZ伧Ei�JªL)��[g����z��9of��<��B���~͕m[ҙ�Lo;H�b'ݒ[���$�6�uhȤ|��qv#��Od[B�շ�}������m��u��Agl���C)r���s��T�]��a�E'�\h"��0�j�W]j٢m��T�w6��E�z�c;!Q�P��YQ�P��<��Eӌ�ct]ܜy1�
�3+8㜜C� c�U��z�3�kj!�טr��Lz%?t�x�&l��黝�ǅ�Oƻ���/o\�z�⤱��4'�vm�|{e��� &��/<�O2�;Fd_]�����@��D����&�<ʭ]k/t��m�A�S(R�������c�[�A���Pڑ��;UVJ�e�V��(%�Ts7�A���A߳�0�8��{u��p8����c�^�D=7[��K}�=�RMz�"٦=�*B�f�}]n�3:p�͒�_�*�:�Bl�DVZ��r�J�A�T)����Fuu�yf![�Y���<fݛ[�M]>��D������V��^ `Gv��fj�q"h!qH����U���>�i�6�n`����65�6뜝�e��E�1Ԥ�'a�s��sh=��N;��}[��ӾV��>�f|�����4Ba����:͇m'r�
ėj�2�u�#���������y5��U��%�3�ևr�:#�B|a�Ql��f3"��J�K�R�$�d�Ov�\y��\t�#�1�z�ͼ7P����p�p��T^=��]�}6(��ݷ���ڡ��G �֜��U�B�&����Bh鋇TE3�Aax'v&�N�.�h)m�}��}=|#�Wc��֣�0���!s��2���Q*N�~�l&�*��3�U�xޘ���t�/����s�ü������j�8���KsS�N��!2���'����zs_E�E�øS:�p�]!�i�~ghТ�G8��S!=��o��S���x��Ғ�4�)v�z�w[���ͼO<�u]Po���x�o�~≿�8��H>T�!?c8#�wD$�#V%B�FR�f��q�-\q��m����7P*L��0���s��}h�fY����sԹg�D��n��.�깝��G���/ � �ې��ݓ�[1sC2vn��]ԟe%*�k@��œ�����8��3ܑ��6���m�3�������b�ge��Z�#����5�%R����N��"T����v=H5_��9o�Ǜϋ���?���Q\兂�Qu�_�L��MCu������ 4?��fs����$!l�A�.�M~�+P��&D��N�⮗�f-?5�(,j���?5�� ��?��30�7S�h�d656��D[*�\��M�-^�v��*��Z��3a]砲4��8y�Ee�k7CU���U�0� ������Z�����Ʃ5�:S�4ҵ�%�^�J9�G#��q����A���LԮ-����:�`�����H��nǯn�7�*�������:b�r��MX��Z��j�ˡy2���r�1�ؗ�8!�y����d�S�i�����z/q �Ց�_�=�~�� ^=:�����+�tE1n���=�.�1aZ��Se�-��!�{��ݤ�?v=�f��~���wA!�'���o�w�~��,�9hmG��v�`x�X��(r�P�؞����` n�h�_I`h���#%�}{6��)�Z$����跞�jS���r�u�#�ZpdsH����U+�(��ٜnԥ�,�h��v������_������g������~����������}����~3��"�J���{����v�8�&���9#VVwj3���5'�,gj��a�L�s�D�ޮr
�"��݃U�k��R���|`��ߌ ���|i��\7��)J����Yǂ�Dr{�CZV't#�}�=\c�co�3w����H�&Z�'}�o@�v���3����J��]o��`Ʋs�SF��ޜ�3��,��Ț��9���О�]<f^���}�R�(�uO�"�cۓ���p�����V�Ւ@3��h��`�v6
W�y�L/,��,P�z�_)̤��q�>-0u�F��>yDjT-����	��Z����9��.4\��1P-�B������t��7s=�=h���N�����"�|
~y_�ڡhZ��+�Û��
\Z�H����ǩv�Z�	�����ĥ�u�v�弗P�k��{I�K�;�RSm &�5���;R���9���m7GG�n�����3�!��H������@[9q{~S�}=����lQ�/��-8�[X�ׇ�~(�R�˥����*�sR�8_��������V����K�e���d7�Kk����ux��g}�0���ޱ�������NGfy���=�����U�
Jz���A�K�}U�cJYDp}UcFi��3�'_�'�ў'�����.���|���L>�Hf��zp�1鞹4G�x�8<��ǔ�˲
F���a>�D��hI�:c�Љ��p��;����l�cs{�op�p�x+����L��<���?C�q�Y���:�XH�oQ����,yӨ#�oM��>�e�P��z��+��<�����0�u1`/hA��L�o�$gn��d^�Ԛ�(����Q�t�̷:�\M�'���&�C�:�O�E��X����]���v�&ͫ͏!��1s:�1u/��ئ�3n�D�ۗ�������eT=���c2�{'0����F�S�WU>=�9%��5�hut�"۳ĳa"ܣm̪�@�a�N�\���_�ރ��|�p�e�Y�<|�����A{�������(�N�,�ɡ�u5��u4��ַ��(���e`�� �
�ۥU^e�9D�Ӂq�=m�Q���l�i,�i�׉pl�{��G>�|3��=�W�u3�b`�y�D���3͑��Y��ms�����%rO�l�ӷ�2�q��"ss	X��	��3�l�޽�m��x,�?,�[E9��j�4�
j �vlM�)��j�P0�qbs��ܽw�==
�lS���ڴ��nx��j����^{s�v	vg'��k��VMK-��cqn���u�� �����'�Oo�6����ʵ���$�8.��З|��z��T�]�L��T�5�������>����}�:砏����跼}�Γ$�=��A��#��­���BnO���U���}|&�Q��+7��U�"�$�~���o��%/�T�4�AHz�̎�@/�]%�
�E�d�CB�J��҇�4!�M	�H����H�TҚGJ4�����4��C�
�b*��<�h�����T4rG%itDkJ�	M:Ѕ-W!9�ĭrOR�A�ҍP��hZ�=O/V��@1>m��4���:[��%9M g�����[��>}�:�Ά��~���3f���w�����O'7���}}�mWˠ�V�\�к�ҥ9U{nݴԋ�/{m����S�M5>�?�ȷx���,9O1q��X�+�����;�I�/�TM�MJ��۹����#��f���?�׊��%�=[�Ѵ�o��'x"X\�,�]�����mR����ًġ���e���v�IM2��Rkۗp�����l��Sۼ���vk����	��K0�̾�������zs�'b�.�L��5��\�S�\:�:<�3[B�]�	��y{v(J��r+�I��1����.�I�0�{��O��Rr�@��h��IF'l>�Y��Mm�2�9:�zV�(G��A�;��T�m�nO5'¡ۅ�mOC�Z~XH%�./#��4��kJ�/U��}j�!Y�<]�_�>�����x��~��&������k���^id�k)~���5;<�+�yEi�7�𨨇��C6�d�F��:�y�C�~4:�W:�R)��6պ���w�M�)��>��SOL���z��Ѱ6}ʒq?`���=��Dq��g�}�98�S���g��k̤'��P6�%0TƲײz}]rk�|����C�O�3����!1`3���z)k��3][Ml<�Z峓(�cB!4������k�-��	���SuR�S���}��ɺ&�<�w�9-�i�}P��~��~�|��i_vP�5/x����Z�b��z��(u�䓜x��(<̭��b�H��{�J	=E~����m�sBN��z�p�1,4 �1\�������h$p��Q5%unI{��g��N�6O�c�=
��k�!��_H�	�.�aط�pA�^$�=�U]s@J�r���4ծ�e�R
D����8\�tԤ�c�q���t�e�f��]�6�5jv�ds���VƳm]ާd>5��P�o���?�?�:2����+�{�Ѹ� �U1RY��E(�u���9Pne��CPH�3�l�*�ΞG=;Ń'$��|Ǧ����5/`�����<���Wl�d�8'ֱX�?��1@��+�A�}�G��*��,���l���QUV��B�벳:�Փ��:Heρ(�ukM
VRaMKnq�uEêϑ���\����im�
��F�6TƗm�v�vJnj�~��=�1)դhZ�RN.���a�MJ���{��fN�vOB�V�]�^���0�!�e#n]�4�t�H�I�x���)�W���)0O�7D�[���_��(c�;V@@�ƑB~�s��,��P�}RQc����#��[�?y�0����A�>��=�8f�o+K��F�J�V�"�|5����1ܖ���ټ��j��2�ϖ~��d\�st{ʏhǉ�G�B-|�r3�4�O6�ֳX�k��}	��7�gi�|ŠS�(C"���)��ׯY�Vn�у�C]jLK�wҟ�-2[$����z������9��?���`�w�F�=9��f�y|󇶄#���!_9��}�}���~��[.u�wwE�a�ڤ���\�L"�),qn�j�欣�O������?��"7���C"9}C�(Y/V�U���U�]k�O�<���\0b[��wz��tóc6Cb�u��sk(ʳ���tj�H������ ��<'%銨�X�j���GJ)����Nt?^�?�#���	������-��,9�aJ��m��f��5-�bm�6�;L�����Z�o��u�{�#�K�	��0����ږd�X�.ܷ$��LIv7��$2�>Ѕ�2]�����{��﮹v���^��^F���:#ȇ�U;~�j���
�������&g)���A���*BH�������xl���`0&P�.&3%'Q�B�U+��e15{���^*5�fF���/���
�"gͷN���s�>�X]S��#+j�2�k��PF�=�Iu�ƭɘjl�B籆e�\]
�U�p���.b��z<ޅ�������l�Z1=�0�E�.v�4�<��t�$TKD� ���C�8�������'U�w�vk�W30��]����egT�~<8�ւmb��ܥPK/a]�pP4t��糳l�s�$�T�k+R��Ϥ�.�nMs�qi*��>��mA�u���"v/A1|[~��m�#ƴ�q	�F�J6a���%6Y2*XhRu'$R���,$3BVd3a�o�zZ��M:#"��|gh��m)ė�!=��@��&��߄r��ǉND��m���q��S�ě��)_<��r;�-�@��[At��L�7��/�{���?]D��&���j�U�&Q,���tS*IRaO�|��a=k�H.͗�.xb����܆t��.�3��1���������Rt�ѩE��m���P�\˖��^=2	ٱ��&|ݺ-c<�b�;����lT��3�hR�4��Q�]/B�Z�C5���]���w�p�ܰ�9�k�݄�t=�2�=m��/����E��4=;4�X56��h�z�fF^���eT���,��k*���H3�N�Y��9K��p�z�&>`���οW���j��ޢ��ҏM��OJ�>��R|��c�^$��ފ�y��u,�[����@xG�v�M"2���M��*��z9pf�H��F��w��ռ�����u��fy���K0���g�7��h�^D<���~����|>��{H_������y�T?w�����7���@E��� U:neɜB6�����<QL���N�������+ڍx�^m��wb�zr1��M�\����Ag�lu���β�m��\�g��qB�Īw���KKX�s�O��x�+W��;#�Na�����:��;Ǥ� ��({�@mMC�C�����h|."#7P�&%.��ۨ�'���o:5\�2������$=D	3��[�}��2%�%��.��M����
��Gg����̡������uiw3Ez�KUL���9Iw#:m>.]��S+��O?e?�WR�%�/L�9��`PO��cm�f=�q�5%LۆdE��	����Zs��q�V�3���#�?����Q�xށ.�08��a�y��OP�X�+����%6Ki�.!s�Y�7+��塵��N�
��
=�^��x =�;�A@�����DC�ղ���+��8��/����s�t�d�N(Ƚ���Z�I��K��3ƃ�^CIX����:|��@����/�h���1��b����D�8��o�%�>9�N�˥y���)��:癱�gG��+��+�ou��K����Ó1er�a�2�`{�L8��F�|���+��,9�^�-�f���+Z�!�=ڼ��, y�~m�����%�
�g�>�1i��2�K�oO��64���,C���h~�ǹC%s�s)Q�|�Ü䒟Q��,����֪�q-�28&�)J!ېs�$Ɇ����ҧ:����gN0˰�SKMI���d�],�6��}z�M}�g(�8��r�Zo��åLK���U�#����1Q:������3.�&��y�긖{��=�W�
5�C��2#�sߺ�i��Us]��^_(�eb��O��������5�]t�C�����ׇ~��ڣB��0P2���<�|H�7{\LUQ��T���5j��D����z��r�Lz>�>�c`oH���<1�����#���>S�uH�6��
L_�o&Ǥ9m^X!U0������3흞�Y�4�h�Q�����b(�l��pP��[�C�f=�n}��A��;I86��0�H�r��sP/�ܵ����Y����F9�M=[��W�3�u�G\����1�^�<����T��և0Ԭ�P��|���0�w��+���;�����8�ͱp��"�Ƌ�f����N7[���{2�3E�$��g�?_�u���˛�ʴW�xkW�g��L�> ���cشb5Q����z���{N���潟���LΓ�p!�����@A�g�ٳl� [:y�=;��`d���f<�W.�ft��G<Y*���B�zLU�x�A>�A��MȣX�_��^��8fЂ�m���X��l�Dy���+UG.��?���a�e�4�c�~ �o������#x��� �e�T�>�ׂ �|F:�{��{b�L���N׏c�u[t��$����K�Z#;��}�y���qb��|��vF�z���Ѓپ)�}���qZo(K"����8�ٝX�<8�U��'�1<� wN�j0y�?B�오�֚��a-�nq�uEãl����ߞTZ���%�GY"�3���W,�^���>ܗnЛ���"��bS�	�U$��1��Y��ae��i�FX/R�h�8މ
1� �}C)r���nt�O�I���d�KdS��Q�J[�k���N!�׎�PWp�|����9	�σ����P�o0<�ǘ)g*n"���*���E�.9�o<��zk�����z4cJ;;A�|�_�"�&#E��w���+:y�`��ʋ
����T$��Ic@r�v	�ݛq�����2n��}[��UT���f�P؁m�C*+���YC��='\]�.
z9�u�$q���-N8`�3e�bz����na;���gؓ�s>74�^s~r;��q����k�-б�(%픿0���i�l�\���c&�۲���yHw�p�{y���p醑���N˲��,9��R�m�Mc߉�i�{�lT��즨�k�J2�s[U��t�gF;��:`]�G[�R̵��z]�Aܢ�������gv��U�ꦼ�<)�&c�<�A�����ݺ�|.s������)��#��W�$~9:eFn��ڹ��ōQ'b^�?����/���1W��G���6���9�Y�X�McȘ:��}�Ž�b*�_+E��55�����ev!1������'c,m���]�a�1�x��i: c]�����  `L��:]��78�k$�o�9C<Μ[e�p�f�f_K�� ��8A�� �eC�m�lg�`L�"ˆ�N��n��̙kH�e���!�un:Qc�=���5������W!
DךE�Ӧ� XT�׺)�,"� Q�P�k�>A��/�r�)`���b�k�TcRɘ�=6�B/y��%�"N��<����;!�T�E6{���m�w�QK�)�3���q����$N�|?���1�0��M��L��B��;Qӭ�Zp�d��S��u�^:�=[�S[;_��L �d�HvO�l�S�܄&7����i���ݼ/7�÷�3�&�����)J�؍�ǭ}Ǆ��|w�	-��:A�	籠�*5�y��eu�V"���^C�'8�%�u�7E2������fT������b�G.:c&��Sl�ΡS��b���=C��?c�t���StS%�a��`Ӗf������:=jK��r/[C�����YF��9, k vpУ�S��jv]Y�O�iAcAt�~jN$�������P&��M����}����☿^�iµ����F�����C���ћۣSY}��e����_�&h�o�cY<O�d��X�wzfR�RL�C�̳yT��&��;!�E&S�w��k�zW���A&��6c�gfՉX��\/9��Ε̞��MZȣG��ZK�xr>�y�z�0{li�!�Bvh��SlPNл%Q��Q��UH�z�>�m��w��T���8D�\9���?o�f�WL��]	V��zV���l����a]�%��T����Л=ەOD��fL*A��_Y�VV��7:m��
7�;�����y��� T�uɈ���,Ɓ��d���x���&y�<��}��z�q�,�ʺ艌�}���2�A�E���`ҟ�B⟽^��-����@�t�ʋ׋֮����
m���i���ۭ��r��rF�ci�C��$�4�_E��b*�e�#��曲M��z��o���{hec#�a�zQx�{�cp�i�/��<
�W�Iw�{yGl�Kk���S]����yз�xi��������Lgzv�箧�_�"��R͈a�q[�(O�=�q����~�6�O:Gx߶`�|-�2/�.==ҜV�Q�v+әu�|�uq�w��
��i���@bS\��z/���з�xA@����� ��_�ϲ�_@��<ב�P�.�gVs��/�w��-�z�%�x���o���IfF�oup͗	�	��w��K��T��?e�f�޹�^X�����jяT��F�'V�������Og�^��%"�[o�}v�x緺1�;c_������L�_���S��]�N4Ƚ�?��+�I��i����|gOm���
��jxp�y|�{F��j4������i�����>y�J~L1�@�I����<��ȸu[��d�&��R�gS�[��� L3sH��f���`� Ì�i'��'(t	\�aͳY��r�oj�*9;m\/�T�s��E����i� �ņ�����*]��j}��Q��m8��v�qk�u���NN!|���17�z�W�,aq��|!	��~G�՛R?��}���}���}�g��}Uܦ�s`�t|��z��t���ч��>f�9/"����6���q�T,ޙ韕5�fK��ժ�[V���i�oOt��̳el[�6��t�4S�6�]3/�=?`�щ��K����B�(L;�x�X�OO��Ms�����64��8S�3���g!񱝱����2}��A���I��Fi�D�^y��rУvwy٬��P��'%��d�P� �3����0(昘X��ԍd���w��L�v��|k��>�s���|������~�_������}�~Ͽ}~�O�{��iً���w)��s��le=9]�5q�U&����.8�{z}		\�U�}�S��TJ�6]cyk:���1!�C��@Z�c�^��_3�0J��:^1l�:�V�%ƴW8.Uh@�W2��InGK�tS9��x��ׂĨ�:d��%��y�;����EyX��U*�Q��T0b��r��u��Q}%1�����~��TΞZ>�1���P�+h��@��������2\��Z9Mq�kz����(h�/m�|[
g���)=���*z���`�k�� ���!^;���b8.��(=�5瓘hgn~�{}d�Mc���S]���R�ψ��DIf�x��5�4n,�N��#N�s��J�o��x^�����£[5{/�.Čhd�q��#��R�����ɂ���b�]��a�����юT�v`�uڮӮ���oT�uo1�ej��ŵoo�-g}Ѵ>�ZFx6X�]�k=ԲM�Ɩ⮦�W�G?>~���>�ʮ&_��fWUhV��F�:�ɉ�kfa{�ދ����}��:s�EهQ@�iAE��Q{"{�.��i�D���6y�#�rxO�Mg;�W�\H��A->��9Մ$��țhR��Ro`���n�T��tvNn
5Ӎ�|��7Nzz��f%�/W3��^0���;�rvm�>)p��\��0�9jK���������	�!s�ZM2ˁ�\���Fj�Y}5l���hE�����<�{+����>H#0"0�c�{�ˣ6���o �.q[�"��M:���sr�r�����#8Ҁ�s%��[Q��m�����_{���Ǿ��g����ԾV�I4�z�R��64�qw�G��]���˼�Z]��猍��uUt������qm��b����~�ǡ��7g0�}NJ���T!�;�O����Wܒk�-����tz��)����'[t_!�v\��Sq�cn3��t�Gi�<M-x�G�^�:T�mG���zjۚ9_S�����1����I�5��}mfW�Q��q���7Ń�N���N��yc`�d]�G��>�;�]iIÛc
޻I6�uj޷L8M�6`�;�n �,���"dΘ������A�un=�Ht"���{;+t�;���͡��A�|��&v�Gb�28w;2�%SW��f��IΞ�"O�j�nE�]��!~eM3}.-]V�=��|<�����gt�v�ﺶ��>T�|	+���d�P�Gi��WM���z�⒕��\*С�ގ�!�^�o��/��������	�������AS���p��H���������n��
�5�75�zg��,�W]��UD��������G��-�<2]u����QA���a�:���@ztu4�,Q�j�����u���v����1�ˇI���%)%���U�v��x�>�c�/�]V
ܻ2�R�3�T��9$�M1 �����d����%�� ��D��� �J&�&�s���CZ
 )V�SHiA����1�(J<H�&�4��9�\Α����#jZ�k67�������06��N��8�M X��r9	���.cBb(4QCIBi���t풜N��
4h����hhZh!��(Q��6��j��ѡ4h5A���IL��u�qR	sP����=Jc��<�ː!�G0�G�$t�t�-�Ei�4�!AJдi�<���8��R��@�I�%---!����UG'IT�J
C@PP~s?=#�ȵ|}�r���7��9�+��xr�Jξ���5����������iN�Q�.L��w��U�r#�/w%�ԗ���H��>o*�x+3�)�^s4��("��0��=��m���^j��!�6�~g�I�uN6ۜ��̳L��mF�d� �\�Ov��e�m�5e�m��={�m��ȧx	�#@ql�ت��um���f��/<"�w[��فڥ�rp�N��PC�U�Q�g��e��Ξy��=`��!'}�����^:MFfҾ�u���3�7�i�Ǡ���]�֠K�z1��Օm�1�"����Y�i�5�g����q�ėi�:ū&8�2װLRuai�IL����O�nlp���ЌYQ{f�;-T= c��H�ގ�,�Ba'i��%ۄ�Jnf�L��s��F��S&�UH���=�n�.�}&\r�d�	"�:�q�!>3�A���S�.�F�L4��J�(��KCӵ5]�-��<��G7r�Ek��Ɓ�p�y�-ᄍ���i&O�&�7 L�@�Ix��q��ܣqo���C/+���iM�.��i�[�#h��= �����l���C4�8n���fM���!�O��j8��ҡF��L*�9+�X�BO\�ƫ���aA<;�@�ח����z2u]JC-6'�!Q��q�����(�X�D��vs����ͫ�k�u"�r�Kz�b�B|�˺|��\p^��N��k��q�Y���۫c·���P�=�3�pV�wƛS�vH�J�N4��n�9'y0VGՋjH��P��=6���]޲u4j�c=s��������!��V��� kZ}��s����d닰J�¿������p���xOp�t��6�Lq�'(�g&�:��0e�͓��wfy�-p[e���dRej�V�������9�^I:�%)��槝��{�#a����38lsH���קe�m�E�4������~�?��'Y�o��q3���>Tޝn����2�eK&����/a���.�����#m�&�tGt�p�3�I�z�˸Du�A��N�W)f:��;`��D���^y���4>�)��y�"9L��ܒ�L�jƲ�T�#ّe�� ��E� �3=�-�<S���0n�o��y)�.Bjѓ�*ٛ�p�����U�m{��#2@_A�r�My�\m:j1p����̋�ɣ�i��Xΐ�a��8�sI�1��f�z�@o+ϔaT��Q�Up����KY�H������E��XL<ß�E3�[pL&�#���%s�-�O�Jl�L���ǔ���z�ѽ4[�sL�͠y�s�Z+ʸ���<4�{gl	���B`$$vP�1ڢ���mg�y1K��'`�O�_[��,v��O��&uC痟�L�+o�������.�19�~.�̸=�
z��:k��6&>�C�-����ܸ���h�Ğ���o%]j��^
��Y官#���x��q�[h>P依�����Ul�ڳ%#�L|��Y��+�����e_�%�jR�}����xO���C�d��U!w0̢ݎ�'aw���ki��BB��O��c�E�y�)�JSW���\s��'�}h�a�>3��x8V�6�Eb,,����}���*��F;_�(�a�*�.��)�yi�n���E2߿v�Oei��O�8��ܾ>�ŗ�D0�1���B�������z^��}d�4I�溎�/�MP���[G�^�7���V�������0�x5ظyr��A���F�3<J�/^��g������iMM��k�[''�m�]�5���<� å�G�8u���ئ������"�_0���'*�f���r�+ރT��_��f��^短�u����`>�,?���G��;HK?���9���o�!�u��:���"gӮLG6��,Ƽb�;3�0=�uޡיɚ�&K�����y��q\��v��_�?��!�a��,ZG0�xw����9�e馺m�v�ف�S��q>96����uߖ{�;���wA4��$@"I5)Gq��{5��J�[�h�wh��oDQvk{� ��j��v
���Q��n
�ko�r�8�s�)H'�^���&�{�{^�^?��mU��](3�: �m�����P&CQQ�_F�7�.��î{��/g�`hL�^�k9��*�#��x�;0>�P~�/�{w����۔���ri��L9��Y�&���!3��O��/�t�`8n�h����ߊ�DV����舖�zemux�j��;�U�z�<��kC=�Z|��Ϗ��*��ϹM���m9k:oLm'ŵ�f�����+�Ô��=�����3L�L��!+7P��Ū�~��hı�:������ҫ��9T;iyDJl�L�ɭ���z����/K߱��q��,.�o<��&eU^U".�����vG
&��܄���\�4�¥I��F��sS:|��w��1s!�2�_7WO
#�Q<��Bc�)�i�1�&ހ~�N��s�Z�ʁJ�[_��fc�Z�Чa�]K�mF>mOf*��q^d��li�%,�S�C�Y�&H�uI��Rr�@����Q��]�����"�Y��z|�>�E���1�nc�l�O5�*]��&�wynЖ�4�2;�Ni%�M�u��r���"����G8�xeϞ�ɦ�u��D2M�]W<�{�E�R��5IO+ k)~�Q��<��#��ݱ흅!�7̹ݓqW�ӎ��b���P�{{�A�ܸO�B}�YI�sE�����s+��Hׇ��`8h���dY�XK��*�D�G�9?�*Ok [���c��N�Ԛ���f��[U)���3�p��r++;;�b�~��Ǝ��jk��ڶ�^ƹ+�SZ�8p�_�7J�0x)�=�L�ާ��ƾ�O�^Ɨ�1��2͚���x��C���jw����6,g���P평�{�m�Bպ�Ë>���OO۷�u)�?s�f������t�kg?���2�ង[&�̋�'��#H;)87�]4"��1\�A��޾4�Sn���gqjz�e����q���� �L�B����2DoP~y;��bK��N����WB��sin���,�y�;���g<d��� �*�i���9�lNs������>nt��T��:�4.Ryڊ��H�e�@/�i�m�������[��E�-;ڂ�h��)��}ܽKL�H��}1b�b�/f�P�Ξy���-��[֔fc�~�P��L+EVP=�M�Г�at�P%�k��[�1P�j��Vv)f��2��cPދ�5b!�-X��	�}�8ŨFB�nr[ʂ�B����
g��d5j�9�
�����l*e머y���ޅY���I�}�#��Ny?3C�E��Jr��7�l��H�"eڮ��6���vءՃG~�U�S��L���3GN��U 6{4f�G�l������+Q��	V���!��~|=�~F1��[º���]�}�#B�:W!��#�^�)�P2?k�򟜺/;aaTں����|�?o��!�z�濄��	�-���8މlY ��W����505�m���}Ko�r��V�|�<�Xn�֞��^w�xa9�!�~�G:!�Ð�Lρ���קD��ԹuCO�Ԥ��1L��n�ZB�y^�z�^��k�ji�9���v�P�/�Kd�Z�#�b!��6�!�hR��¨�}�nr<�5�S�����܇ǝʁal��(���[�U�
L@���6���m�@�:��Ī,(Z��2�u��^�Y�/�ϏU�6S�mR�͊��\:�=M���G�t&��ԍe@v��:���c�k��1�6��<���٧�S��=p�[�Bq�^������� >'�,V�s�R�z�#M�����۔�_t*�^�'(j[�}z���̙���}�S�e�^T�$�o�Z��/B��`�m�9ڙ�r5�(q�.�	�c�D̉D[�@�r��.�4>J�kK`�����G��(��æ}u���,ý��#vGpz� ��	3�tE����u��̀�����E��6�g�������Xı��߳����%�rw�mm�^�$��DX����n}P�<�+�n(y;�t�<>,�1`W|�/�̊�p=Cף�:���9É+��k��m�̜��=!,]q��yi��0S�V��o�v�r��)6��7��C�<���[����vm�=\�X�x�,���Bɝ��p��tԐ{�\�D���ѕ�ɣh�:�yg�b9�{C��}sE��^Ե�JB籆eC�.�2+��4���o��n�G\:{VLT9זrSe������.�,$"[����;�\wT��+G^rڼ4+���G����흐/miĵ�@$j�EKK��WI��ow���SLݷ���'���T�Tj�i�	�p uŤF����a�؏�f�h�[�Gt��t{�eyW�J���F��u� �W\Vw.�҈0�_���jk�m[�����t����Z�S�D7^��6�6�0��`�!���ղ�w�߲S[7��H�Ģ��!�o;��k�M)�-�0Y�l>AU�]���J13K*Z�R�g�_G�����=��{h��a���6uWL���V]�/k[.�?
�cX�e-�[0gc�z�K�z��^7�A쒲�:D�b��t��{8�Sk�LG7'��tT�ۭ�{7lQ�t6�wj��;5W��Vf��+�ã{�iR����T��T�
��M�_#��zjK����=�����?v����5}y��zv�g�Nt��;���Q
�L�O�7�o�H2�c2:s*K*��I��o�4�m��χ+��v�	�;B��w�G3�>���Z�,����N�p��s�~k_�/ޛ�3$c�Ԡ2 &���.篖$S�?[<̪��~���١��Vkl#�؞�)	H(�=�@-�c��c�]?)%^�/��6��k`+�B�JU��7��tC���b94��<̟��w���=sqvrUz����,�÷��!`l�QnE�k�\��mu��^O�q�����+.�F�P7@f0d[2%�n����=��-6u���T��]�b��%"��֏e㋚s>��AR�x)�kD�.9r7�v��;>�@��%(\���s��X�sݣNPh2�E��M6����aD^�J�c�t��#M�Mx�J�J���`�3������D�La�=�g<FOca������#�&��y�<���^����\U]&[�����i���#��������u�L\L��G��{(竨��6�uB����<o(��CÌ�n�sUȨ�N�AnZ���X�/S+*x��^l»��o��e����+��j}��nq��E��z�>��d�x?)�H��>�iR�ܸ�I���.�	z�Ӻ�'/H�Ĩ�|ُo��!�!k�;��ѷo��}�=<�fۺ{�ԝ��A��Y��;eOst���#zvcҹ�>�s�l�(U��v2H��>�;:�SA'�5c@.�-�����웏v`#g1������$\��l�4`�P�JU^F�f���O���=^r��hܾw~��RB��>q�g��p�bV�a�OuW��v��
.ŋ�J�n��8k����y��va5�χa��vUx�s(�rqZ�.����KQ��]���h���GPe���X�uYq�#��9~Y��S�=����;������56��lRQh:(�S�g�0_3��b��9/k��f��szc�R��NHr����<9m��"�ϴ7����y�֭�������ɇ��.)�φs��v�B���ۚ`^젺�\b�>��=U��Ѭ��N�XQw�;�"��L�)C��|���z������V�V�vp���E�H����7�1� WA�ȸX�s)3�X�;�L71�eέ��x��칳�,��w�3_V�e�!���C
��T�R:Y�	����f:���ޒ͏d0˥s9zxFEO�%�|A�*Mq������+Z ��.z�aDV���rh�в0A��E������WD���7�_�0�޵��a���\�;ٵ�x�g�y9p���:�|�R;,,4�,j�B�
��W�ػ���5O��n[���)!nB���iMm�\<���r�EwI�z�]$��R\t6��j�5������v��ޯ�ޭ�Z���mWl���_�r9�J��W�������?�J���p���X6�u�҃�"4Ǻ��xv%VYtq�J��%��`��ׁ�+�s6!��][wSn,��S�p-�ْ�Q��=ܹW�w��v�,{J��ӽ1�4g@a��t�'�Wi�A��=�:��������~�~�_������~?���|������v�_���=p��+Ƙ>l��
�7ˀ��k7B��j굇�&Y��har��m51�o�%wF����8��fq��7�6�D���<�X:�$���ek�ŭnF��ߙY�r�F���$9��j�ɼ��L�E��Q����&�U���̶I��Sz�h�m��_�lW{(mJ�4�R<}��v���
��.n���۠R�X39�:2cj�);���C��[�=u��W]*�u��� ro�:=��M��ۧ� = ���u^����n�Y�`0���}g�^�int�kt��R��z�҄G�ޞIo���o��I�ߨ�M�T�O�'#����jBc�����..��^��Qw�Dv��3��Y�
iY��B��R�����e:�}ݭG���/a��3p!2���eq\D��U��H3K��';z�ص��6N�=�=��'����3կ]�p3��X�#�t���q�Ѭ���'�kb��ջN��5Ki�����>O��yE5N^�����4��u��aDu�i��P7��@��ga��SD!.�H�}_��(=�;�����o���Uz��I܆n�[(��oɄtt���w[����60��(���/	4�pw1ɗ]��@��iT-]i�i�e�c�c��Lnj���&��R2w3L�].�A��� :-�T\���mdiuCz��.��F�?{٠!���i��� ��e��rcsV���{�Ξ͠��}-d�x9L#��֞�aI��� +����w��+M"E7	꒜����{��-){�p��(m��O�p�Y�`�d��	N�i4�n�m�{R+���<ğy��R�}�t�
�}<�v�"�g�{_�/6"��f/����������Ӥ�$g�ۛV��k�������<��8�|fG,b{����Vp��+Ex��ft�\�b`M�
`Ti�8D{�<(�֨�=�P6�wS2�7n�~��ar.��_������ѓ���6�lɫ5𣷰 \�z��$w�y�cWH�}�m�kfs�2�:JO�酽����_<���(�^+����1�:n�o��齋v�(~�ū 8Q���Ϛw�����cn����d�I�h8�B�=�s}�K��|1���<�&��T��2<�N�c�M�RX(;��Bn�t���:�û�<�X[�>�$�Ђ�z)����1�`�Uk�90���	ƁX�arH�B�:R�b��q�b����]Q9��y�N�u!���F�"B�v�j���)wyG����l��7�n�U"�H�x_:���91���0]���gzV�ڻ֚Ǣd�+\����Q}{�{�^��u�����6�uW|}l.��_��l1���wFE��L�N�p ��7B��O��q�I;~���T>����TU�M"P�@��1!T�EAE1w`����h("B��䁡(b�$���5M$ETIEQH�L�P��5s���-ID�E--4� D�ݖ&��
�0`�b�J��"
���
j���� ���R�����b�<X���
J�؉h*���$����h�>N������&�b��))
�����i�&��U^,TDP�R�P��}�����(�������
B���j�H��?|��ϒ���N]���Hu�Z��Z/5���v��3a���5X��t4��x�pJ�5�w�ه��i���%-�v?H���'%�n���<��dGKv�|���3��q��p�r_r�	v��D8]Y˪�K���n����l��4l1�/��C����hЉmA�,[���ḒO�*H�6Y�D�	$���]:m�;P@�r]�Oݍz#Ij$<]ǕmN%~���7{��$�0$�Ί�y~�y.�\΋���ݬ�����:CcE��S�ht�Q���H>W�ʈ�ܛ�C�A���F�w���6^\��@�Q�
�=ܚ�����Ċ�/bt� ��ޭ��Ԭ���g�Ϙ��G�������qbU�ڛ3����t+�ݵ�&�M�§�'$���s5l���nC��cP�-�߶���Sܵ�]���ռ
�F��JUO�s�m2�L-��A�y�m�����_���0i'�h�5��	W�2��Iw$����g���԰�������+�"g:����:��be�p.krB�ި�P����v�V2}��E8Oo+&��B��6�s����*m�Ͼ�c���w{����j\`�^<;Yx ����_P_}�=���%H�&���H�,cC�v�:i?K���:���j�'�z�������zx�W�_v9"���*Vv���X���<����s�>��Ӷ����}C��91�gs�в�����GSbڌ��׺j���Nd)�ў�?e�;���~V��>��$�O�e�]�ҫ���n��V�Lӯ>� ] �ƒ�7q��"6uC,fB3�gmkwhΎ�+����m��[@�j*WK������Y^�8�e34C��u���8���ţ y����8cJ�al���T� Lt���w�1��p+���$���fCs�3F+�����h�s�[�����Ϥg�[��Ɔ{=����l��ly"�!�����Y��J����e��	���Eџ�}�C����q��rx�8j�f 1 Et?$��������)�!��}�ï�z�{s�r�� ��x��b��K8��A;U#S=<��>�:�������u��x��ܒ3~2���r4�`��ڱ�J��4����K��ѹ�����=���C�U����ROb�n�38���Bi���̾�7t��8�W��46�kY(_X� WN<j-�1���Y��^�MmAM$6��VN�U�n���C˗��0G���xl���5�q�eT��l������:/�w11(�M4���۾йzw=�`�B� �҃#�a֏]��9�^�*�n�e���O	�D,�D{N��[:����J%�2ror0�i��{��}��d�Gb���pq��r��C��@�] 6�a�	��J�������Í���VLe�oe��o=���GV���2�O�G��V�>wJI��u�A���}����i���g4���ųm+ r�p�l��.�F�E7���2ߵl_u9���h%K���Y��;eO���rZ�o9O��f۸�&-���#7�W����]�]o��]��V=D����&uc�bn�h{�p �:;�u���d�>��<ht�%�����*�#i���̻sB��Ɣ�2�q�x���j$dt�H�4�8,
�/�h�Tf=����w��Je�P��]���pgi��w��8ͦs:�b����#̄��X'��,	���7G� ��QΚ��߹��;��}���vO���5v'��v��Y�4p�g8�籔��ќ��K�H�7k������p:������6|<͞��WU�jF��	#���i�,f
_�?�O�=0�#Cd-�ò<���c���$E-b�u5
��p�񖘻�u�?=�'
�`c~�0'�:��\�Ky�e�7=�T�&�g��n�tu�F ��	<ܤ��㢈,o��@ц<�~ԍ���kʎg�ץӽ��#���!�ǉ�y�m,�E'-�!�SS��j�ʸP�}�U3W���W�RW��:��c�ڧ:ݲ�#'v2��u�#_����w5g�FEO�%��}EI�q����k3_Z�JE���^��vgî�^��v3p�K�֍�iQ��z�|��y����m+�r��G��~��>Y3M�� xzX
����+V��LKݰ��������ʵUh2��_�K�)��GfD�$�Ȃ5�8w4����6�W�˚|�=Z@��I1|�$�7J���ml�S��a� ���LX��u}!�0�y��w�=���_��ိ��/L6^���w����;�M��<k����6��`Ȩ^:; X0M�O:�W���vMʗ�C���n����;��6�Ȃ��V��]1��V�˫wAv�˟���}ڧ𥎷�ެ��2~����ϥP9��/o*�6ڔ�o>�==!�c=�4ų)�Rj�oT��Ah�u��o���ԫ1tq�I.�K.[S�Φ-�U����s3S6����u�ٳ)W����9;�Q5�]�*7H�ؚ���[��t�,����|�;���	3���=���gԙ,YM�BZ�rp[�k�1�c����q�W+�-��:���h��q��+4e�;�_�e�=��kDu�꣧J�n�z.}�#�٣a���8��\O>�t�k2��7 κ|<��٤l����6��$�1��i�xt7RܳF`oMߣv��k���8^�<m*ɼ�}àf[F�p�D������bC[�P�ܾ�����M�<�Ԕ���k�w#ل���H�D3��S�����>����u���+�3?��0�P2Uzf����Ek��rM�!����6�����M�۠��0&�\%:�+�^u�Vq,ײ�#kY�!�X����_F����f�q�GY�u/!S����]����v�8�jZ�WM��4Z�3&S���|�U�X^���&}¢���]�KdwP�Wk.46=����b�.W��5��+�N~�շ?TK�,�z��0�$bĢ��s����v�{u�l�h��D��U)9>;WQ.lU��p�n�d�+3+�g�Ƚ��s��B���<9��'�P���s��=4��*��D��}�x���0�˭����wJJ�c��3�$���s����a��MmomT��y>-�*�c��u����<��imҡ��U-؆"�z���U���V30O��!ۂ��]c��PS@����n���Ζ���]ǎ���C��
���l��6�[5�71��!�ҳuݽ�1��Ш�<��&�O����ހ�z-�*�g�hv��[��c�C���#K�G��(��V:`\���#|�0�����#K>��ڼ�fL��� n4al�χ7�f�c�������50|꽈I����k4�����Ni����޿W?b��<G��t�G�gm>�3�I��$Tb���x�%�%�ޝ�� �jxD~��^�k �����LH�ЦE�ಲi�������w67q���FWCz�,[\���cp��;��=8����D�_�24��}�̪B��?���6�A�>�b��}�_tv#�����&�qu-�;� Һ�2���q�Pkf�U�& xG���%C5� ����$6kb�}e=�9����)����JǗ�΃�B��]�tv�0�R�qI��"���6n���o:(>v��D!��M�)�S�{ �᪑�Xsr��9E�'��SY�1h�B���J�(�fʬ��8�mc�kARW�L�*_L��,G���;�����������֏U๧1A0��T���s�7&����(B��b��u���D�JJL��7f\kUeUKv�������&��M[8����*�"�n7��.�ܒ�0�dp����'^-��4���n��p����Ƿ��5���x\H@`��e6��w/��n����z��&�wo �&A<���-��6� ��lG#���n$�TNİ�,o-��d��E���8�T��չ�( W'RY\צ<{��<��{Z�ӓ��D� o�4v>��s�XP�d�l���%�+2ȗy��u��0c�Z�(�M|���{�I�]s��mA�D�f���>=ʺ��ݱw&3��m�Ў�+�Y�8��7�S@�oi�/���2�S��������3��'f��ضtp���gv��rk����lOZJh%�:��v)� kCY4v�C�PYgKI����,�鱳:hҨу�]�H
�L�p�݊a�m�*a��gE�h9�1�o�H��Ћ��Od�T��_VP'���tF���*�����,vy�z�b��PQ�+�0�f����G�[>�; G�/;m�3��
:�MyM���Vh�@vNu1��4s`S�u]W<��ǾMa���8gnߞ��z3\:�������K�KG��2����q@��z��`����32!����@�%�~����9�=���k�3�G��ߠ����=J\Y���s"&�f]�GWW��U�>[²^�ߚMXf%�0�[Vϩ�z���z�꙳�#"��e��*K�@�
��L�;?�ʵ0�Iz��-������z5#�6��o=�^���{G>G��X15���
;��o���A���|�OM�6˶�غòm����_�����=�m�a�Iȷ���<'����2��'�R?�c}0�<�U�����8 �z�n��b��*ʁ�-eC�=�zC�sfv�vF�T�H�=l"}V΅t("��|�A�G<w4<WՙT�����zh�F|���h��	�}�>�Rd	i!jr{���J�3�-
-�o�_�s����Iq�6֊�7��o.Ȅ���]g�����Ë����`��ڂ���% ��d�r�pl�����Xtaa�(+���>��f;��J�m�I�J�-Z(I�gO7cV�:Uow�d0b�a+�":w��*��3g���˖>����$#����1��̓����a��-����
�գ��+��P##�Y��7{'�����Jhdl�������X6��ƢP��8�Y��:qv��.���s��'�F�4�0��������A[�ʭ�Y<��7�mR/x{��$�0=Wg��x�:��Ucn."��p*+z&r�R��[��Mi�lZb�'�O�"��K�U�sk�����w%b|cx�v�%�n�����{�b�۶��CWmJ�|�j��A�΍S��7^g<����s�C�ި'�;��[CMѱ���i"�ZI���}���&��pǨˣr��h�~���}�dV#øt�h��}ȑ$�P2���.m�a����]�3�0�^_�5�A�"�=%;.���k3	\y?N\�K��nFs�ˑWi��w<�l5�>����^f:v⧱��'�nk��~��Whr ʺS�E�+�s��N�E��+Рcj���dC`<�-=x��=�4D��A��I,0��N��SNf���AYuy��1s�2MOC^o[N�����o�D��O��Rz�<�)J���miѪ�ne��do�_T��Ʌ�?\���t$Pc��7��TM�B]N�붘:��S��^uD7S�o8"�<R�m�e�c�H�*m���/a�wDC���rr�ن}ݾί2n�Z$ �Lj���5e6�v�=ޟ_��<�|���w�����}��W����ṷ��r�����*�3*.XG���p]�sIu��^�d滶ap�_Eͱ�u�y�^��"y��.������j�miv[ӈ�����3�]�ߏ��
8s�����Iy��b���B���R��d{A_6.q���j�_�Owl�S�T0�e��mry&�p*j͇���m�Xd�E�ο	����+e��ۈ8d��ބo�?/��xy���X�ڇ_�Cy�aݎ�'vtLY���GtgBd�ݡ"�^r���(����͕�'��5z��,� �9��,���=.u�ﲈ�����t���١��sܣHwmA�H�U[�3�.t-z+I��2�/O?<�|��!�Ȗ��m���zf�*��"�//���i�%$�GԧtV{������yzu�q��x���HO�����=Ͱ3�4�y��X�4q_��y#z�|VN�+,��:(�N(̳�֎��G���:�.��ǥ�܋΀���Y�}�t3t�C�у�L�Gm�:_s��N�:n��7�|B-{�W�8,���6Є�ZEp�ӎ��O_V���}maAB�iK�bt�xn
�]:ڰ�U�!�k��q�Z�g>���{B�!Z��agI$7��x��;M�^�W��MG�����ݕ��UgQy��|���b�P����y{����K��Y�DwLMW;г�1�����zq��,���:Գ�lBt�8uT�C*iK�WN�ER�O��FŇ�ǭC��5���JncE�J�Ǜ��**��G&��*�����\s�J��|�R^��rzt�z��jS���\��#זG_�Y�3I�yg�WI��w-7O���^5��"|�d��>�-Ӵ@<�����*��V������җ8�<�`�ZD�:�5�WYլ��8�#��0]�uK�]��b����p�u�#��d�;��lU�3���\���o`[�|���s�u]�'`�y�\���G�~�+�>yz�dޫ;���3NST��Σ��U�S��p�5t-w�	����-��Δ�����J�#C����h9�-K���;����*ݮ=i�;�{���'Z]���Kȶ��]7������wu���$�v~ɜ��ه���ܘ�����W�B�z��W[Xa��3,I�oruq���=9/\��h�W/|��v��6rMM7E���Y-�̲x`����%��􍧺b츺��K7z@�p��;꾻y�W7b7gEQwog]��	2������#_�����0�d�����r���?_{7�b��ڣ����P��%1e��Y�eJ���`9ڼ�s��^��X��v��<��]S�#'��Z�A�y��z��|�hX|x'��M~;�w]@;�~���e�O/���/f�Rȟj� ��y��o�Ī�u�j�f��;]�8G����� � �R�5/{��g�^�]���x�ќ5�� <%�P-��|N�H0R� 4H�ܪ���ֿ���G�h��������!KDAK	@��4��Q4�EE1UUD4Md(�&����EQM%�T�K�8I����(���K3�S1P�ЕA@Q0�TME)MD�MU�1LL�U�DEDATTE4�Qx�AT�P�5D�QU4�S+T4�L�STQETSALEU:TL�QA�ࠢ*��"j*b*�bh���|F������j������������L�DDSDKIDLU1TRTU0ن��&b��&�����i����* *&�i�I�)�������1AR�D�QM4�UDIQTUDT�i�����*H� ���"���wk����ǟG-���]X;�o�۴�}�z�ڛu].�3�"�����rk���ѫ���[{5�d�θV���R�%%i��	����ca���)ɨ���ב�����D���fv�ϘWC��5��H��I/;�"�kh���;������Y�$���H<��[�gC�@�2��)s7��1���/Q�vg���W�%�Q5)�`\���g}�6l(7��/g1���F�a���F��s�Q��9��{yH@�� �nk�*�r:�-�-?p�u3��hF<�g ,���#�-ў����(T��-���|�q�yU�
�D�j����wP�L<+46q*���e�9s/���yq�Z��d޵���{[ �x��lS��3�!]�*�N{��ł���r�����G��O��#O#@�By���5�M��|�بȉ���6���&�ns�>Pn��"eI�z8�+�2M%Eiͥ>�ee�⺞���SY���Gl�X�އ���u꨸�D+�PS�Pk�8�"j����搩�V[X����"���G�����V����_k��ƀ/5&8�l�w�s�w�v�'�k"k��]x=F p��5���έ)tO`��*��2yKD�U���������u\��N�K��G��N�FtW�Ҽk������o����&�^>��#��4�Z�!v�	i2��;T[l�B������{.7�jh�U�U���C
tV{q�Gb�mH�֡�$�U>��{�}�+:w�U�䒦龺u#�^��?M�Z�8���FsGҷ�{Ǔ�}&��c��{����ދ����x�t�Bپ �e����>�s�N��m�{H�;+���Tׁ+e���;ag������(����ٵ^��8�s>
[��Q���R�lu���]��X�\�;�7�y�W�k���2�-�2Xg2�}3қäѯ9T;���t�P�}h��/b���[N�	"�����1p޾�R�d��E�]���ۇMPf��P٪��*�aZ*;hd����w�
���6B�Úzu[>S���s�n�3�^�/i^L���/�ў�ǝ�s_�'껽���M.�E�s��KK�u���!�y�f��+�W�C�Ҫ�]8	>p��nn�^5�/5v-�2�Y��#w�Ї0U�MF��r4�]uT��]�b0���\�_{��C}�~(�Q��z���8���-%j���u5�?�jW����r�?"�Y���F�q�Z�3��/7������L��D��h�MC���d۪߫F� �H�Q������r�P����w]N�S>R�/Å9-C��N/.�9p,�:�|D�*����G��`��;�7�6���K~��T��qc��P�S�3g�2(�^��4�e���vM����Q�㝌zn�]H��+�b~���,g3�%2�;Fs�Y"h��}&��o:%�i�B�.a!�],��U7{Q��̺;dw4rH�F�EI�j�)HܷR/�#�.�r�&��ⶲ�E�vK��A>�nm��w�$�BԸ�m���r�2ŐfB�W��x0D�V�M�G��f8t��P�/��WE�)[ϸ�Q4�&�3(�^F롯���C	з�qȞ���vv%TqtI�K��R��A���n�-L(��h�q[x�2�\�{�E�sT0�˞���=&�M���[�D^�LEA��f����k�p��C��{)���p*���-�=O4E�a7�x�!|(��}job����E�qd��/�����-��;���i�s��?�#��]�+�ȡ�e�q����w�ӳ�5����$��������J�d��0��Fh�\0+�d���iʖ����9[��@�޲�'�t��DJ���#�����g#{0���"k����7�0픰�He�u�z.w�d�g=~$���Ρ�_-ɘ�b��x3F(x��-����8��d�A�_�s�GSBh��.vl��$r��v��E�<*5�>�Gstf[F�p�H/?2�몟~���TG$]������+�p8(�,�%cf���n����$<��*H�m��Wg�51��C=����翤tS��g��  �]��3��͙��μȡ{�y�Wl�N��1G�U
����yJE�9��΅8���e����z�5r��@FDv���ܒ�T��c����뒅���ÿpn�	�?2��5�^�;}��<�.�.��C4p�}�P�y�-�wh�J�p'U����o�ڹ���<��׊T9��=ޜJB��P8�W�r�������z ���]���N�+��WԜ�|Ku]NRv鷛��=�����<�9&ڂ���N�w���� ��Y�ov���~��3�hG�5�|#N��t�����%AJT�5N�u���l��rN<ڃ��{�q��!(lEo�H����H5�r�mG���U���З��d5ө�@"�䭩��X�/��E�}I�c�ީRuŧ;��la����]��`�0O�V���5�=Q�8c�S��ݷ'�/z����O����I������~k=Ö���a�rO�  Z�L�0�RC���4�F���]��J����2�8C_ñ�74�;p|}�Fo,�r[��EF�?�J�-rq#�
�Y���lv��P�F8~ߎl���~�^P�4cس��#r}�Ԩ[#�P�S�LszkC�^r*N0�U��Z^�7�A��-3�	��#�̌�������|4�c'�-���;���D+�S�+��6�G���³��w�ki�{[YC�4w:z��iډ��SK���g���u"�^���<�O
׻ݵ�s��1+y�U��,W36��U������,R�\N�w�'gV,N�N��bq�q�Ꝃg�Pȴfv��
���3���|rfL�y�Ggv�+|�/�#;j��;�������X��x�gb��d3�p�t?$��}��&6�������#��c����hH�g�5��b��YG����(UYGޤ��A�����D�UY�Q�7"�o$+�:<M%@��3i^W�V��Dזy��)�x1������D�C�q��W�����֭�mp�$�dN���LV��74�B����p�[�U��G:�(���$5]�KgO-譫�#g&w*�U��k�@p��tV�������^�]�t��Nȫ���;�Ê�E%T�P:�ԍ.-��^Z�������4�3y�YJ�㌤��ˍ6ɒyu�؆���u�y��玧��#V5Q�j�$��σN��獴TЁ��+e��|{ew73ݦ΃-5���uؤE�>R6eut��{��gf������IMy.����ꄹLZ���NfdLcy��ÖH��A���%�2#�	ë6��N=�o��S�y�B�{�+b�?+�[�	Y#��|$,�9z
�����Ӂ��}�w[G�bL��bgL��t�חbZL��lc�Uj/�>s�ݽ��#Q��s��K�m���g��7[��_�4�L>�o������ٝ���.nH�I^鞭��ͷ��;n�;���Y����"�X,�p������%>2rw*J�]�M�M�[��D����g`{��Os��^s��؍l����c�2�������Z�x_M��4�4�eW�$1��>4�t3��u���j�~ܦK���~}�f��I�7����='y��%��6:��ݖ2���42�\�O!������b��c2�y�$H(����-��AN4���c*3Z��N���t�T?�fdR��&�j�.-:��J�(Н��Cv]Fl���D��s��a8��UG_�l����z��Ѽw��k�}���:��;2��,��q߄Z�[Hw:!���қ��v�z��;f�x�4��po���:�?�s��5 y9>>7�,�~���_�(i�xaݚL91�5k}��()�b�q\�S���α���xk�A�Ow:�ah8��bߺ됵�I�b�_���7�H��,_�=�f�ZdFo3]��ӢX9Z�U�c���S㩡Wݽ�P�\Ab=&��!��U|��w\���%�W*~�����5Ʃ�m��0*LT�JF���q/���G-����]�P;aH�
=���7:+a#~�I+��IY���S�x��2ٽ}��R{-�E�h���F�Y�^=�%V�\oͩx���&.�97��y�\��0��ꐅnp<0]=&z�|�W��Ѣ��.��A0�d�Noo�zN�R���6@a��cj�؂�*�׏�'a����F+:�}u�$�U���b�n�7�:Xe�#7<�_�
�ٻ9K66[Z�ہ���g+�9<�,�ڶ��R�] 썞���G6D��Nˮ���]���E���
F�t���ѳ�l�6��ʦ(nУ+�_�b(Z����3�$���\	��;��������[�_%�+}�b�@xV��7�w��ٖѻ� {}��8!O,��b��K�<l]
Z�^�<%�?����Oi�������0։�g����=�/Ώ�����Ś瞵������<�A������N������9��ӌ<X��;Z�rלHH�D�cJ�9������z[&��ԩ�&᪊�����7$��3��
l�9c�;������#�G��Ǐn���.d_3�G��zJv^��F���T��N�h�e{�A���#�"Orj���
�E��O�s��=ܞ.����^tDm>ֱ֞�z&����]��AR��+��^R��s;,�
6�:��gڇW�Z_S'����FD��G���^3�>j榜���U��X�d��e�lH��Sm�^�"Gb��r�D�*�*!M=����u=}S����&e��3�V��m1V����Ғ�f���3aϳGM|۩ؔ����6g��|��;"�D�P:�u�{a����G��,Ӝ�;�4��E_��,����[l0�A�d�պ<�͗R��Ò5��c�Q�����>sW����{��;6]�=����Y���8u6p����H���tO���:��PY= ���_��y�;aa�y�.��|?�z�����M��}�~������"p�I8'���g�)MJվĺ�]7�/j�D+0W۝3��^4�O������<��3�޷j�'�:_ �C:�o�ܹk�7SjW+8�Hc���w�ɓC���M��X�����Ps����C~�o�f~�d�K8�j+ҟ���;�[4A��F��᎞Wy��1���dnH��Tal�-����Wjr�/aY]~4��f���� l�1���9�u�[l�HY[��Z�ە�A�|�ZT�����P%��cf}(3�v݁uGF�$6�u+����l���|{�9��F�O#�"G1����M�P���?�{FR^į���� �>��y�q\�V��E� ��״�B����S�Ng�-7�n1��̤1�����l{Zd� |�'��i�I���;Uy��	�@�5�J�#��3ib�Q��Y�ق͢�c64^�l�}��а���%���Q()��*���O^�e4��Q�慵.{�D�bB���P`Poj����U���ҳu��*��$R-�[w�l�t��U���x1��V��~\�}�|>߯Y��~�_������~?�����}>3�ļ����[9i���ۆ�Or��3Z]��_Cupon_d ���������[��YK���pH���@4]1�*���(�#_2���1�Jr6{�^���K
��ehf��f�ᬹ&�ʣ�L58�f�#����t���0?>[k/���IpG&(D�{�� `q^�=%^�P\ۧ<�gJp���&�KZ��B�!����A��i�C��"��Ɵ�|�r�~b	�Q�yzJ�kCׅ��r#/���f���q��G���-z�B��ޘe�X�agE����طL�}�=�;E"�8\�Ć_01p�����{s����3vx[b�jF���x%�q|)b�˗�R˗�1���_�s�uҎ�P}�)�k�Ӳ�9��C�g�:/�0�!�R�]���v�גN�M��˱��a�I����5Rm�
��P!�C��]�x5�Z��hj���f�㾃��q��/�%��=Us<(��9�����Ya��6��m���/y!�%򎭑�e��k�������{z�އ;ʎ�p(���s���N����tI}ñ���"O�Tl��ԍ�!��糹�d�;uug2��D��:�]:CX�K���r��J�C%�s�g��C�A�g�!=զ+�@�us�sY��R��te�X{঵����ͣ$IhsH�2�D!S����������:�E�S�5��pW�w�f���aٻ؃�F��wg:􉙘�M�r�h�h_Lеm
z]�;�Y�*U�s�p�i���A}�wxtΝ��_ ~�I6׾j� ��]�>\m���A9ֿ3O3�F��v>T9��p��/]�9��ˠ�=�WV�N3uKa'�ΥN��h�=w��:=�pc��T�gp�����m�&,E-]�z�i��%tڠAHS��[����[�p��3�S����A�yP<��|Y7v���b�z�vbb���9vm�x���)،u��z	�b��=|'�?M������mMF�s5�6u�M�Z9Z�uΖ�'����j�7���L����(��C�7�F1�Kp����&� |x���p�ңزw[��T�������H6�}�w_C�ϙ�����`y���L]�u.õ{��
$I���w��)�/�{��N�%�1;Ï���3E��4;4��=��.��kE�X}��$�;o3�}:��t^O#/bg�'�>�x��&h�r�w�2 ��(�
(f���*��!SCe&1m��+}�;�ݎs����~����q�΂��K�]Ǡ�Rz=�������XŎ�*��"</k:��k�[t3���9>���jt�el��e��]�ߖ0�T�I�M���&=fur`e�SD��.���gn�+�ӎ
�]�w���GW�T�'dy��M��?n	�m�
��<G�8^���w���i���q+ɱ\�W�{lb���GDu�6lhq^Bj�&�t`4��W1KQd�>RI"�Te�*����"���kĘh�a���������(�b���bX���"�&��(�"d���b� ���x�PUz����DA�RMT4E3D�TEI�RQ4�EQ7�x�PDE5$�4�1EP_1�������
����J����*o1�����3TL�PD�$�RCSUQ1DMUD�1@�l��4Em����&�&���j��"��bb ��
(��������� )��h((�vMTK�AQQDD�DSTԔPA3UQ�CMT��EQLEA1G�j*�^cS%K��D�3UU5USPP�QTE12Q���L��CU�g��~���w�����uNّ��=���������ȏAV���ˡM5i�Ʌg2�S���oN}X�6�4�8���?�k��R�vI��x�.N��ԫ�%T�]r�K�+� Ѭ�S�\�R�n���L�4Yt���)Xn\kͲd�]D��{|�9:F>NU��=��8)�f(.:}��6�SC�)��k��R7S�x889���wF�(-e��̧#T��.�t��{�L������K�%�'Y�TS��Ux�v5�� %�8�k���Pu�F��:M0r�w%U��V���g:���67$�.�~�`�'��d���8(Ϻcۛ�Tf]�kDi7�Vg\�t"�?oQ]�Fvm�6�=����n��E��R{��n�|��y��7���{��u1�D�{�1�d�Pc��s8;�SP�P�t[u�>��8��Ud�*����='���|Ih��F}��ꁱ����u�Gw5N�k�1�
"��<i���wM��,���H���7��/o��=�l]=gw���{�P1�q�
��
>�3s�0��Å����fһJ�xyK=�|1�3�dy~�g�����%�=y����1�G����u���룬�o�1�mŶ$�R��V�k�Mv�e�	a���fV���1��Vم�Q�o-���r�krz���O����c�
`֥�,צj�.�#���<��ѐ�KL6;���,�n���n����V硪���=T�xL�����2��~�=�b����v(�{dvp颤�m��ED���� �,A�~��[�ћLf�^l�NL�\�zX���D�A�<����'�4�4΁ov�W;�N_�������V��{�lX}��4���4<�RT)N�0�z�F�s�)��7��Qb�y�E��t\�
6ۆ�X݅>E��oG���Ԥy5�m�&�����;��m�s��O����t�ƍ�0���\����G{���杌��u�N.G1��OHa�����]c��U�T��9�S�ɭ��YNz��`�6�x�q��;
�� >��2U�,yyc��Lr���خ�׃�o���O+]�U� ��{|�+q��7�P���1J�a`��}xn��R�O��_^�;6q��t�e��m��Ήws��*�L}s�;r�����o��Z������̳�HaY�Yd����*+k>/���1亼����T"��+G�"���T���w�;@��k�sZl��S�J|{r��,�S�G7!X�?6�����;L����b3`쯆��ݪW(X{Vh��JĮ�vF��o�cotޡͧp_��"r�������q�{es��9>��.�����=�=�Q
C���i��T*f�]pԴ0���
�2��AW��KI�H8m᜾�[檺�1���z�kO��t�� �C�,�£^7�����w����h<�����˝�Νo-/��S�/�3��@�!f<�����A򼋛���ٺu\c�`�:C��h�<&��S�O��{8�L´ɘn�1�.�o�ti�z�{q그��ҥ ���yJ}sNdl�Um{���Q�(�M�i��Ѿ�����8Ü��i
���U)9>;V�Ib�&�\ٳ׽�n�A�f�wKǛB��r�V=�� ��7B$�O���X6�FV��i]$��ˍ趩����g�Dc���eq=ө�[��Sf��e��M���kv���n6��u�1\��73غ�/{��2��q��������;?I[��q������d����g�i?E|wy��v�c�8
�����1.,o�ŗ������Y�t=�{;�p��qjz(�/OX8�U��LLi/���!�{ժk_�c�����͒���8"�:+h	��Ǘx��*1fwm�q}��3��E�b+Z�fv��_S�aO�v�6,L�p*c�Ϧ�����%&�e1���oQ�~H����0:���_T�흠�r��hP���C���.sj�WjڢQ�W�'��\e��r��Tϳv�VpÔ�ϮXZ�
�#\g���S�T��䳁D�P���E;<�pk�	 �F�	�O�}È�`8�g�#rF�R�al�|9}3/���[����$A��kyL�fB���cy�sH!}�#$,�-�m�Sb��ʩu�j�$�-Od�' ��>�t٢�j��#�,����35��#_;��jy����q"x�����(�ا��o ���.�i}f�m�٭���]f*����mT��7x�*Пr- VR��N@�gtX�7�J �K�u73�g?�}Ѕ��[sL*�SE�u3e�&�ٍvu�qQI4h��,��ْ���������Ð����sTQy|��~ۿ���lh�7|C=�o�_g������{�o��eV@n�j9��E���2dg��ҧ���'T��5i���_�o�x���x+�CV���=����+�$�ZG�K]�v����ý�Ѧ���}���
��
k��
ɡ��D-��(� Z�z6�1T3�I�}�^[ەC��ˉu`W�
��uȃ��R.��~��C�d7o@�{$g[�����I�.
L�ʹ�!8m���9"U���ʒ��ne��z0s4�Ě�	��P)*��P=�N�ix[<8��wf[,���+:��>�d�v��)[r�T��i7����>k��|0�-��r˺����"ݺ��m>�*w�.W�@l��y{��Ϧ���	����k�6ּ[�a�ޘ��힞��3ֶ:�S!�Y�"r\��.�79ZWcs0���#6�댍��^��͘;Cm��ć�6�v�����=4i����#4��pQ�t�����^��l���f���A�חm(��^�Ƅ���J���&�y�/qřt�{�Y���~�[-i7n�k������io���z����N~ޖ�H��O\yh����됩��L���������OR�Hw 4�ۺsB�Y���]6��1[�Rl2'ԟH*>��{��g`v�������a�yik���MW�nOKv��o.�L�[ G�1�TH9<b9�ё���C;��:���b����T� 5��gړr�9��r��L��d��D�#5N�#��Z��_,V���@0�((����S�V����C�4Dq�{c*H<�,r����J��z~�haaD!F<�h�M��2�9^S(��~�3>�{��[qݹ�5�� ��	��<��zY���=T�E�2f:���9׷�gL�v�d�4T�ל�uĹ��ԝ�9���.�.�&�A�����]v`��Kч���+�J3�}&�����4��Bɧ��Z�.|�Ά�c�<)�j4����F��.��(�5O��]j���%Qy���юh�Gd��y=�="��R"�)m��v�F�"St�����ưm㹞��UƯ0X�ty���&�A�bU'fk�ER�N�4n�玲,���.^.H{d��A�W���y��°f�,0��~=���^U�O�O�V�^�0뗙���`k�>�� ����װ�D���K{��9:�����.�O�[}�vў���H�!/��y�{t����A��m�g�'���e��l�+����@\b�Zok'%�4d;dl^I|%�����.��� ��W�K�L1��[��=�Sڡ��&��n�Om���H��TO��4�{���R��ce�G�i޵���[��^m�Y�6w^�}7�*�=�+��S�������\S=����Hb�)'E���v����j�J՚8�R�] 썞��z;M[����������hMB��pS[+��ܨaH�.��z/y�秗N�n���o��=g)���$�����_W�BW��6�`���|�k�\��o�ٽU��[>�ng�� w�Y^�hd�O�q�>4�n������ݹ��=��7�p(�K玊��EGO5�G�a����f���{��{��i�ރd�'o�9@���|vG*"A�M"�����6�wS{=��ޜ�*MP�0�Lt��t�v��֣ٯ��>�͍s{�1T��5��#/	�Uբ��g��������h�'��	�{����.��gzd�f�Ob��~n�O|ɔ�/G9=��q8���g(Q3�c/���#�M�,(s/�{9�������w�D�����\��Fi�m�AO�R+���m�9�t�M\�n�Ph�%��ȫ>uHÉW������IW�T��5�1�9v��=��{�H��Um~uǖM�tDj�'�p��]�Ǐ��}���1��\GuN�峝T�^�u����@�2@������ķ�h�l�]�^yٜ�?�y���z�7��$���k�R$k�"�Euzx"���Q5���9=9��Zx�����P�)gouvy�l�A���<�N��5fm7
��и竴Ҭ��l�t��K��&B��!���Z�ƽ9S<�Zՠ���1C��|�h��ڶ��bB�1$�ύ�t��7u3W֢/�C��@�� 8;ϑ�=�*_���lx�j3wws u]tN�<�tTr/pFL
�����<G5 v�{p��W�-^�n	�����n���7��m.�%�L}o���
ۃ)�0����{.~�����W@Nq{M���iT���Rau��#��~!�sK?o�^�w��9׹�z�O���:�\�3�x�傀Ϸ�o=�-�@�o�z<�_NN��.�Y��e9�^g����L�j9��c��6�@T6:yNYʠ��.;M�ߌ僿5�:�l}���#z6Gh��� ��=�������p^h~a�"?��c�����I5:w���w���P��ezǤ1�;�3�u�^��}�h�#�v^������rFt:����l�m臝�&��9�VRֺw���oo��>�T�_[�i��w��p�u�HD��â�᪑���܊�֤���	)Jۺ˵��K�"��N��59��VVϮ��XK�p,{��
ɨ��D+J��a5nm�K.�yDα�1�OZ�z�ni�
*��>��5j�ю�f�+��ce�/�'��ǃ��*Q)AQ�NUΫuV��
b%舖���^����m��EOR�i�vW�&�T��%T�Q�N�i=}��IŻ�O�����]w_h5�^�e�79��$9o�&I��N�����M���Ӫk�f�����~5/��p�;0
�Z�On���ּ�-ȝ��/mi>Hu�����-e�N�EB����+�s�@�$�g���x��N�y�x>�z<�/���=�!�L��G�����V+v5$�N�[��Df��(�{���ᇰ�i�ܓ���Nd�����6���x��*x��Yl�4����[tݛ�=o{<�i�.Tqn�������B�==أ�c�&������K5�gh��-��yq�J���l.�}m̀�t\dlΪ�4U��>ئ��9uwD��nv�7�f���f�
�1�F���Ͷ֖�i;�����\��s�m����W���'��od��m��g��&�fg��b�H}-õyz3(l���dG��sԭ �|Tt��>�w��E��mo����.�%�q��׿vx�cy�Y��#ti���I�m�'6�Ӑ�|#�M��#���}x*}�V��̲��@��Cڶz۰�3�������S�]��l�ӥ�3��B��e�҈��̳����C+0���Y���x�����{9y�w��K]������r�JH�
 *��*
"��s�@	�䊂"П����ǡϩ�sxQC!(�2,ʳ�2��� (�B��00,�3"� L+0,�0���̣0�ʳ(̋0,��2�ȳ�2���3�!�0,ȳ̫2�³̣!̋0,�� ̋0,���L�2�ȳ*�+2,ȳ̣2,4�³̋2����2,���2,��"�0�ȳ (�L2,��̫0�³�0��#�x��2�ʳ �0,��3"�3̨��P0�(�(�aB%*�
�������@�T�A@�U@�E � � �4 �VU_|C�Ua� !� !�U�P �D �@ �EVUXa t� UXeUa� !� !�U�V@UXeUa�0�UX` eUa� !�U�  �f�`XtV`Y�	�f�VdY�fQ��y<E�@�`Y�fE�`Y�8��a��Y�f�eY�f�F`Y��oQ�8<�����T�RPD��PӢv�T��%u���|�t��$� �3��	<�GZJO��x_�j�B �Y�9���MQT�B� ��z0�@0�q�8B�S�݈w��
��r8���y�!e�)�J�?q+0%��6A'�b�E�P�E�
(BDY@Be	�P)R@��U��U�a 	B �aUaBVT  	FVU� !eUd� " �4�T�p"C���p��?��"�"-@+B��`�G,��@j��&��)� PVA�A����~&�	�i@O������ *�6��7�`�=�XU u�
��d@���(LЂ�
ݬ7��  
� ��D�y�|�p{���yO�|z��	��
���y�P��x��
��i)L�eu����l@0O�X}AA�( ����@]`N����.�ܳ�$dH(�$�^�:��+P���T@_)�g����2���6R@}(�]Im+�T�f�H0n��QT���l.}ل�ܟ��
�2��/l��2�����9�>�����UJ%)H�R��%$*T% �"U(��"��QB�P�J$�*�J������P*UQ	@�U$�m�TҶͭ6�j^�+��B�V��4D)�[4�j�@Ԓ-��BZ[R�V�&��
�����J��2)���-l٤�:B��"�	ڰ�Sc%UY���$l2�Y�M�UEd�&Ke+HS`��T�i�j*)m�ִ������5Rh�Y�l�D҄�*�^   sxkj�V�Ϯ���Z��������-SVҧ��;ټ��V��V��v��[3�koM]�x�GݧC�ݸn��]{�Ҩj�=9�zʚWp�^̬�T[P՚�5���  oq}��cldo���>>�
P�C�P�CC��(hz(P�C���СB�=�Wl���*�zݍ��\���C��ӛݺٽe�oTf�۶�ݳ����jWm%!�+BlS��%
�6����Ҫ�T��   f��}-��{��cKf�n�lW���V�թ���ӡ�N�]��޷v�:ӷ
�ۥr^ս�ع�V��i�:�4r���4��{���Ξ�J���:s�UJQ�d�V�� (�&�  ׽s�U���u���g\������N�Mn��X���W-چ�{��N^�;��h,��
�m!�^`y]gv(HT�i�R�lʴ"��j�T_   L�UF�}z�;�^��3v���꽃U^��G^��^�ha�v��׭jimdӮ�{�W=��7�=z��� �v�I
�٭[*Սmݐw� � ��j���_f}{]ֽ����Z����,*�!��뽭������8�B�5���C ;Uz���Gv���ѳ!UT�-�(� ו���Z�1�4��6aT����:^��]�TuW�B�z�&����  �s����r��]��Z#VʦFUM� %��  �
�}���@)�h�@�4U�� 7$�� ��`( Հ i�}n��-ٷ : 
t����D���T�B*T��  9χ� wO���(oR΂����i�� �K��� �+� Ѯ�9�N� ��8�z� 9�9�A^��� ѡM�AKѕ$[�ګhо   }��
P�p��P�� @f�� 3E�@st� HϷtz  �/n 
t�� ��r� t�S�T�@4@��a%%* @Sh��*P�   �~%)P   ��*J�4 2%"LʩM  ����_��?���������I���E�c4ʩR�۝�곐6L�Ol���������ۗky�4UWꢊ���EPE܊����*�+ ��)����?�����鉻k4���^�)�1ZJ��;�t����лWr��[y�)�Ie�	LZ�̰㳉֗E\�ж��b�Ucčc��$��m@�c�&��8Umf���5b׹��֫Ԯ�t�U�B�l
[ʈ�m��Yn�(SLTw�F�צi��S�����lOܼ�S�v8�CP�Â���X�fX�(�)/��-��!`��u�i,��o�Vo-3u��J�a�X5�e^�aU���P^h��n�ɹ7uc�PHڭs~	�����E-,��U�ed�e�64�2��h#�aӦ,�l/�q}��yxr�SEս�@��QX�R6���%���E)���J�i^�{Q���^n�S 1�h��v>Y"�>���,�k�NR��gt�y1f�2t��(樠�ɻ 䠐�k[��-B�^���k�b�64hg#x�@�s�*���`�W6Gy� RXu�F�,���Jl�$�?j��Df�$�(I"��7�O@^�`�w5	scnm�2T������̔oh%-n��%��kM�����b�PˡFm6�D�0 � [�6�^��t�3���J=�{�g�*-ڸ��݋;�b�E��]�X�����0)�*A1���K``;���	j�"� ����w���c�.ѭ�2Sw&�M9��J����M�x�jM^;��j��j3������x�t�X��'�j$��6��;qdK و1���SQ��ba	%��vLY��x�(�j�ٯ^ͽT"�hcVhV[CM������{��`�5Y�"潤q�x�]�ͬ�r���&�b��.�\��׵��:
V�o_��
�ҫ�A����՚��Te���p+��&vX��5>M�"�g'ֳE�)/ٖ�{H+O7c�D�(��٩3�%���qj���Ķ�V�Y-3e�xے��IB��7�{�St)����{QU�`bLڭFO4٥(<�[(�M��`EWy�Bh�Z��<@L�K@�f$�궭�� �q��c`ÏSav��j2w��Fc�QH�'e��R�VI�mim��Ѓj�V<�/T0�8�lJy{-Gw� �2fńS��T��J���#JkoS���T�cJ����REԖn]huP6�i˚Sײ@6Y���7f	�-9���R�KtlՙG6ݙXce�� ��L�
.�`B���3,�3�4
ѹf����f�ϴ*L���9��x�ώnϭ<��\4(轻i�a�r1�@mn�ę�,�[�\N�l�Z�H�+ri�Թ�oD6��r����,PZ,�m`�a��n /)�ؔ�`֐m�J�jz�T�Ju^����Ƨ�M� Pєɐ�*���`�N.���!�g)ǩ:�b��P�j	�0��O2��nث�۫�������(�ӱ�ksD�D�Ƴe�L5��]Ɯgg�t*�%�h�Km��լ�N���H
���"/1˕q��ۺȯ6�����SyZ&�f�N�/M-U,Ҫ�VU�� SDc����^��+U(�� @����9��"d��3qf�8.▯qd�Y���C�t��r�Z�WI\����n���iY���M�M�1�/e�Y�нP� �Z3jPz��c�d)�fá��I��TI�M�m=t��-� 37F���f�qkTf^��M2Csic�/*]%(��X����W���Z�ں��Z��;I�ЙF��VA�+`l���A�f$���X�g��Ɔ\zis5hSW����1���B��3dV��!6��)��gm�hZ�GB�ҵ�k��KWq8qк����*}&���[Y5�dz��e
��:Z�4���1����v�"��=���xM�@,W�d1�Uap��a�4,�Zj�;Jk7�SB^l��`�py�bcZ�M�qޢݛR�K��Z�Yx(�LYr[(K�gK2�Y	��Y��Ҏ�U��la�BFZ,�"=�l�Z��ЮL��7�-�#�YNƝ	'3A�2�Z m
1�ٻA�e�p��`e�<�Xm��N�+ٖ�F��;��6.��C:�v��[5 �+s^�b��GCg^��*`�Y�Ɍ�:�p,;GU��E#u+iY/X�q`i`zs����S`{)�����6�U�n�̣�Tu�ML�����` SR4]!5�
�[�k�i��H�ʛj�Q�̨��t��i��� ݪ�{0۫��Z쫩-�Scj�C��prl.�ISѢ�
V��W1�)s ��3pla޹�V�ܬv�{�u�Ydͭ��h�Jn-�,f|�SA;ؖ�̅ZjPۛ��Z�͘�����c���ð�\.��B�L;P�P�g���כ�u-YīD�Xr���u��l�0j��(�B�{)ͱx��ıl�a∕��${vj�R�X�W�E���QX��IA��j���wV�u�j+U)�#V���O�K�;X�dI,{x�Pv�Q�a��b�	�7b7�^Z��Zh*ShH��]+
�9�Qz2���2��/*�n�Ŏ�קp˼_V�:��eA�'lV�;� ����Fmޭp��͗R�a+*�=iM���BA�Dc2��	�
��oo�2������Ն�n*�-]+3F��w�q�"r��yIJ�d���tc+kDu���z������ծ�e�Ű"���7nޥ�m`��Z�ś�@�R*Zb�Ji�.H���kS��`%�8��mGw�,:� 7.�]�mT0g�7cS9QDۊM`;wQ�[��ˇ@v� ���Y{h�mPn��1�$Jr�h؍�!�-$�+0"f�Nͳ���jĬ�x�˒唭'tՑ�
i�m5 ���;����nݍ���hҬ���	Q��f]�*冪�ԗ�=5�ݨ�i�卛��{�jl Qp5��b�RKf��@ʆY�ͬ�E`�ǔ��tK�fb,�9+8F�% !��Lf��XB#hId��3� �Ր��+���� .^�m���(�I���
'�1Sun�wlH�*I�EL��9��b���x��+�X~�����=�v�;�J/N�A��h�B�Y�u0��u�:u3
"�(h�r�a^i�8úG�(^jXo^d�Ы���c�w5��z�&Ii���/�B��{�K��^لjX۫������V�b,v��jlV�P��Ǒ+��4�ujJ0����*9PV��)M$�Õ����[5���0k�B��vLml8��F9&ʽ�)M6]����Z�66Ԧ3U��^�O*���V\�5�l)f����M�7�F�Z���iz�ݢ 9�+q[���qO��oH 8U0���^�O1���Y�Fv)v�V
����@�r�I�խG��R4�w���}��`�
�4��7{�1
�^⣴v=�ۄ�'tY��tܴ�8��ܵ1�A��ˤ ��Q��n��6��y(���B�Rk,*ʛ&��	��v@�՝�+ �oh���&PM�qY
��>�]�M[%k�������^i�����%hHJj�3���F2�b��5Pk%LrIy��^;XM]Y�t�ا1<�-j@H�ʂMY��*ڤ��
ףu��+1�)N�^�`��u�L�/5��54+��M��-��v�4	 Í�'&�m$ m�Х(�>�g\4b�+5 ,-٪�^=W*�'m�M�J��Xm)�ѸV�YH6����s+R:�E�z�oA�AAR���|��mU�E�Z������ظ2���A�3���N
\6�]�i����k�����Y�U`淔P�sMM�����k4�m�E��.Sֵ̎�/��4�N=��l�m%z�mD�i�i1�Jfʱ�[e	��1T�,�Pݼ����v�347*�7Q�����N!ur5��"��	CMùLRxkw[lY9��m�5�MA�e]��J��׹k"PK�6�*:iP"�SV��u(��r���%�$�VC�],���ї�VG `�YP�6ܪ/$[w�4�mF+tR�K�J՜��FY�%��\/mT�z�pr�7N���-���ZC=4�f`5pÈ���*���($�Y�)A�/1V7���4hKw��X�5�;ًU"#x�b�%�3�5e�͏Ch�Sl�0����41,+Ҙ�m+BR�V)h? �����3+my-aeй����œv 2���S��z�u�mj
�r^��� ���6�l�w�[v\T1X�7C��ǩ�#!e�o/h����Z@%*@fU��Ȉ�j�q9����)viH�7�)���n� ����]`*�q�#����g -i40]���&֘q,đ�`���J�d�.��e��&�1�k `�L��1�W �{�QEh8RZ��T#�Z��tQ�C��7�u���~t����:�i��	B*x�&�m��c^<�x0|��(0��Jr 2U�(e�D�P=��ԭ��-hL%iz�-Z���^��.��p,n�wq]���I����6uPP��7cx[U�Nn�Ld$���!Z2�9we��1#��a�a�Nj�h���	*jmi�P�����������g.�qS�I�J�or���z��b��"�����04,�X�"��e7C]����	!�E	��uhw 9�fAZQ\�4�t�� m�):�vCs.�\e�MJ�V[є���hP�sr�ܼIKۚ�}v7vJ��1Y�K� 7j����ۺ�t��wJl�%�ݡ���.ی�d�Yf�a��Me�N (EJ�	Z�-n�����6qm#�V�C-̩u�������z0$���@n'��V�ft1�4�>�9��t�Z]����Ɉ���Bݨ��.���IT��m����f�n����m�L�hn���ŵni�kh���VkE�qU�v��+c	4B�"ТfK�ծ=W��gP�V7)C��V r��;�=�[�ȴ���JU�^�����Jc+H�`VB�-�e�DQ�`�aͷ�����;�T���h�L�`9��	a#h��KSUa�-�B�)&�
�$i]�X;*�8��n�W���X
͋̕uY`�{Q kN�"Ҭ���0kL=8Ɗ�fcc��"�7SKAU�-�0i�����X�ѓ*��?n�ӥi;�6آ6-�b�{hl���\�#x��ˡy�"�W݄��<�U%��CsD��͉R.� �.�pҫ �z����3oJ�R��S��]�$���,"�̋즖���&~ݬp��2mlgt,c5�[��N����Mgm=׊"v�����9J�6"{X5�Y���mL(F����7j��/i=jJVT�k#���ɤ*v��9�� Q��̆���O�Z���Z)5�(ŧF�D2��ec��X�͘FGsCS^��oHN��I���@�Xo(މ�ɒ��F��E��"�.��&EJL���lѶĠ�Y���
�V�)�gv�zR˖1Z��mmur�5f� m�dӻvF�t�֫�l��]X+�N�U���v��i�4s*�*�f�PeA��IڽrV�c���I'�h�Р�Kf����#	�����f]���/jax��9�dC�Q�JB�t��/6��8]�o.�zUۋY"Y£�R�1i�۽Ս�bP9���TN:x^��WR���;q�4�c����)�5�6�pf�gڀ0(R�[x�K�ͭ���2�$ǯY����J�Е�40Dkv�ƷI�QlV ����[ʸHX���A.����v�b�D%k��T���3N㕷�	�!SE��I���9/-m�o�SNm�V���X�:N-vm[�f�����F�˶����vC���Ⅴm"i.����	�4[:`_-:`ӻ��	�3{G\��{��S�Lh�zŶt��Mܕv7,��Bge��v�JY1��;X[50� ��Ůfj��o*��x�����p���G�^n/��j\chlSE�*��f�Ĳ�wD.�%E�Q�Bj��T������sZ��B�`�������CfenѢ!I�z ��+7)����-��#t^�I�r����V�l��X�˭@�|p��AJ[feɲV�	�B]H5�v�]a/�9EV]���@�(%֤��6�F���e6N�V\�.;�kH����nV�c`�������R��m]EZv�P����ڕ��Y+B�!Цk�ux��H�K?Z��3T��Ӕ��%�eY
ѨX��Qi:�
Ym�yV��yBô�.�J�`m̲�1aS��)�#WP[��e/��+3w�u�|ANH�V-�zCf\�+��%h����:˫؞�3r���)�4m�B�x�ܰ%����դ��5��y3PH�|��m�c*Á�����dD:��8��\[��6P6��K�u����Ѹ��M����ڽfr���+A���*n�S��n�h����l�>fiSvS6�ek�鹬h��[���+�[�5�z�CXڗ�h�D�x�Z�X�K�S��c�w����Uܽ�`�^'�&7`B��ʫAŃaU�Q8;E��mc᫂p��,:��(�7]Y�Ӓ�"��',���Bp�U�IO��G&�;��Ҹ�a왫�i7#�Y	hqjɤR2��z\HC5�������-ʕ�WAZE�U@�2Bob��aF�+���R���Z��֐E�e�J�r'���a�ћmk���'1hi�#
�AON��YDj+{�:��״�����5�ҭ��	�gU�vkc���Ƶ��7V��:a�i'H�ܱQ
��QJ�X�0�T"��=D���2�Tr���WNU�r��dֺ(�Ӊ�����f�v����Ǆ6�^��f [*F�H��凅Vhי��6���Ϥ�I�c	�(���w"��ʕ��!���D�>]�j���SO�=h��G��6Ĕ�]�e\��D�_\��������vk�p肩p=u9[6M�%7r	Wݢ�=�����.�0ȍq5�;�)ܬ-�iC(�F�Dq��9m��ۍ�6�fTg�6Nâ�*|�:�-X��������YX5�����Bq�㓈�݋_K�e��}�,A�p8�;]����3.a��XN��$�6�1s�9����+�}�5��\�V�ur�B9�{�ή��;3�����̶/�3)4:�.B����ih��+���B�HYκ}�\7�ډ��S�C���e�;Khuf�����R�+�S1BײV�U_����_��t?�JdDv���WV<Gl1˻kG(�K��5.�.u)V������~v���;9��үUʇ�'�^Ǣ��{�c����Q�a���`�XRŎ��,A���mҼ;�2
=��9%��-n�a�����U��e�x4��vf-x�N�r���J]��@Y��k�}ۤ4λ��{��}�a�S���/,�Έ���>s����oX��B32��\����\m�g�V��ϭ�>�M!��w��k�z�(��pP�Ĵ%;Zc��a�?%�ei��WlGZ���a��b�簓�����h#Ru�8Ұb���*N�^��]-�����l�Z=�74Q�˂�^W�*����r���k��w�:bޛ���;����OT�+^,�h_#�-	�un�љ�<�ޅa�X�j-��xZ.8�ɯ�ɺ�Y�4��!�V��Gv�^��6j��V�h����skzW%� �l�H�5�F�4��z]v>�ܢ�娎,���b���
|�3�[X��w����K���ew^����W��9^�;.-x�G3`�Gf��˗eWX��7*:ܤ�~9e����ѭkiLZ�Y1��-����"b�q{@-ի�X�����dU�Eo��wƅ
X�Y�������݇yG;�]D�m����8Ln�0k��Z�xS�-ܩ3%�8��Yv;��5��)V�C��q���TVv���J&�Ι\:E�4�3�p�f���쓆b�k�5-�u�J�n-�X�[��H�I�k$V쐙-����l�/U�� �D�QI	#sX`��;X����B�za������*�H���㲋])%���-�8B�-�/Z\<��{5e�;���io�8Q"�H&�u�������:�ء����פ����/h�� Ԣ�eh	^h�YR� 5����/.G�-S�a���^���]	ۖ&r-Hu���Ts;4Ky[��pT9�}�:on6^�f��՚w�f�i�X{M�$���Ьr��)I�\�-�+�K�ՕPW�����h��c��	�����N�a�/Z��+�Z��nRÙQ�;YI���o�̣[(�z�������#9�6�嵋�-�i�:��%u��ۂ�f�6�m�t�7��94����+F6榦���G �dk5K8j@$(m��ͷO���T��<�c�+�<eM�*�]�Z�n�T�R����J��mJR��y�!K��7��Z�y��VB��z�eg�Mҝ��eFɕi��;\Ǜ�6lS��`����eM$�޺�i��RWpc2K��/WU�De�n=i��A��gd��~Q���s�,�d4͓�Z�6�1>�3FܙҶfa]���v�Ze\y���9���p�;4,��:��L�r�Y��5-�����S9�ATbH9��Z�G8fagy 2JPgC5T\Z�e��l�u��a��+�k��$�PG�F�}Ȏx퇐6
�����aV3��-^Τ�Ƿ2�����,����]�Oe�ɴQ|��eu�ɛ��/+ڷ�@�`��-|/��QT�gN�N̄�Z��=��6p���0!�b��#��um�"�^9���Tp)�����8��εz	ʺ%8Kܜ��u-8pr��\�Dku�y"/�֙��^Mf.$+Q�^��� v'ˆay���qow�e;��K�v���������Ĝ9��n��t^]���h�������]hVR�S�g�P��&�Ce��M�\�o	*M�.��b��v5�{u��R�U�d��@��6��
cj�hes�V:S|,Y�9P2��nm�1�o�~eZ
�r,�M�ƞ�x�U�놎V���*kh΋�N`����!���Â�Քn�u����E2]�h�w|D�eDD���'���S,̦���+��w���sR�JѹKM��� 1YiAE+Kr�1�[�� q�F[���RV�3�ie`�>5a)��~�;W!�n�G�ǿGv�:�K[�oo&k�X8��-��U�n�����):F�����dꚖusZ�U2�S����v���k���,��]ZvF�qw��́X~�ӫ�ܫ������vD�t�ı�d�jv��m�\oO�M�lR[�j���:P�2��M���z�P�;8�ܰvʴi��]e�d��^�1�4㠈�_>�cJ�β!�s&aМ�CwVgu����3Φ,Y-�_$��K����[�r��Q&��q�;)[�dfn���B���yqfv�E�*01?S��Ag�M�V%�o@�a��2�op�ӊw=�KD�<w,����������ݽ�h��Ѣr�u	�z �{��`wñ��w��{�JCwq�I�TV�ٜ��n���j���i㗴{��Ϫ.:�͢A@P�Q�o�Wo����v�-�x��L� ��Aņ�5��Wp�I��S�g�\�U��X���
`����)�Aj��`XѝN��]���D�s������Ġ�2��u:��C��J��*vctN�r����9
Q��o��a�v�����eI\�͸Egf��s��-ţ���]����[���J%�H�ќ�Q:��Aϩ^���p+1;}w�V]�vvilx���]�Q���N�(gQ�ܼ��is�t���G(�L�٠uC(G�|5ܾ�[��ᮭʉ!9D-�Y��jt����	����Ж�Rr�t�I�cx7/��R�7$t��W�f2��L�r��<&s���-��f�<�B���-yؙ�R��C\-��wm��-Vs�����,�Z�s$+�8K�)�i��YX@�Gd0��C��gm�����v*�.�.Ɇ��*�D�X�%<��� ���i���'%�4!��b�El/(̂gh��,�������t����LJ���5�
���f�IG�#/��>�OEke5g�ѹ��gN�0dz�y����yy�fF�dw$��%����yM�삡�о�C+��Vc��*�(+\�k�瓹޺]++/���R]R�%6E��\n�w5������:^.�Ȗ�oiT�w�T�;�zc��Jq+G{^3!�s��8�(Z�ǯo2��ԗl�S���۷�@{]����0�)cm*&��cv�M:l�*=�E.ݻ:��]������-��m��E�(��h����������9���PWt���Λ�ݬ���vŁGvʌ�X�u�id�N-�ݱ�V��ꥮ�6b�ه��=���*[�#!����[>/b�.I��|v�'+Y39n�c�U���ճ�Ed:J��W�Y/X��j��"�!Y�Ԥ�ӌ6k�K5�&���d�.�p�m����-Y�F�)M��Ü���SrkN�Vus�H+��/��w)-��Ē�6�H_LW۬�����!n�5��������ZO	M�,����)-O1ME���,E�PVb�V*�rU�+�m���K'���7V��N���D����o�ܔ�f��7�����h֢	�w��t�c�&�̙8e����&jü�z�[�gC�+}���4W
5��[J��Z2�#�g��Lu:gnqY�J�GU��ף���[/�3R�Xw3X�+�b��WS�@�D�^*���K �C-����:n�M���ԅ���˖]\�4�V��GP�Y��Ԑ�5VJ΍�a3��.w(z=�^�i81�[�q9ٸ�]�J�ʱ&���<��5>qFk���6/.+D�&����>��4H$���ԥdf��:�5�nJ��r3Q쨪��lW8�ࣧ.�)��F�\�]�;閶�թ����9:l$�oC����k��P�B<Nnv�<��S�7�;�X�8S(�ZFfo/+�����=.XE�Ta�@t7U,��p���p�lv���Udv_l�N�I��h�����S��MV�S^k�^����,�<�lv�n��շř�] ��ykb4��=wkk�]uj�X7Q�ٛ��^�Z3K��oD�^�ݮ�̳����6L�at-�\�q��3�,��:}l%��d�� ����M�e#��:89l# 8ޛ��,��A��a�� �xSn��ѦX�&
��U��e�
NŞ�=��^�rxi�5��ޣIR�9��k��s�6���{���yQ� t�?M�ND���[=���CR��,��g�����#(㝷C�@��ʕ�6��)E	�R�����S{b�k�u:c/��*�j�<	R+)go:����+(H��U�M��P���05B�N�:�r��;}N]
NczvK��n;��Y�����(�^m��j�$r�׷�EF6��\2����]��G̙���g+�b�B*�U�B������Hfv[r���z7$���{�Hn�ai8�+ ���ŗ�����qit*d�]8���a�uk�<HЩ�n@��M�I>0_+�C*�w9�#0wm�UΗG]�m��^����9^�j�d�B#Xc�h9��پ���Z�o�.-��48��"��ܜ�5����V��MF��B�Y��Sy���l�kj�C��Le�[��E@�s����H�,��o^g,��l�Q�|2)�j�em��'ԉ7� (J���υ_.��D/�6i]V��V�8������[�Z��Գ28��+uM�;b@ƷFuj���-Ȕk�mWom₲�����R��U4~��J>��b�wR�|3�s.]`��TZ2fb��V���.�|Ś�L��zn�B��w5׎�8Qt낓;�Ů'(�@N�u$tmQ��ގѡ��Բ1�� \g&����z�ێ���7����M/:X��Y{�(!������ )H�jװrM�Ѵ���ɸ�$4:�ƾ�"D=p��	�1y�ذ�l�}�{�bn�3������G�L�S����.�v�v�A�(�Uٚ� ��Y}(�[&�Ɛ+7v�W��N������1�]���k*J�p��}�9!V��]��G��bn�V�[�EGg*��$�HGD�����=t^���-Q�����D�\�n�9�Ĭ��-뺜zu�z �`�M�s�Iloq������n	��=�����*����#�O'����5�2Sbbq�8��u�Z$��)I.Ү�E� �ktL� ���pH�\��:S[�^vfS�J/+���`Т	N=�-���v���( &v�q��Ț#]�������(MZ�)���ч���9��J�@��H}-�[���k/�Ayyϵd�9z{4=�~U.��x�]	�O�lT�'{f���8��Y�V5���]��������U�{���mV��N=�♚��o8�Bl=U}�W_)R�LB4����f,8����ɱ�s�q��i{�q�/��-�3Ǻ^"��T���k+�M���=�׮�f�����=rv�]Q���=�w��
p㰼�o���W�4_�J����,�|�����:�E��'R�	I�}Af�љ��[��:7Y���Q����׻������DA���U�����˅[|�:���V+G5�.̬�}�uNX�QG����cB��xH&k��@�uK�5���^z�`nV �������Nֺ[���]l ���;�mU��p��
����gk*�I�����6kx�3��X%�B"F�=]S���K�`:�
	�Ρ�Q���3�O2(���n��{(�e8Np]2�S��d��h��l���*-�=ғ��Y����W+s�'sF��ެۂ���YV&��7j���,��J����e�6��7:�gb�����0��L��[�l�9�p�}f�bXܕ��ի��V�-p�����xÛ��k&Ϙ�h[jM2�~�6���v�O_e��ۡ���pd��s�����kh� �0��wU�!N	D8K6���.>FkoT{5�r-��4�����*�l�ܔt��/���w]{����ڵ\�u���@.���F��M��#�v� ՜��,�V��B�&�+�eMZa���R��'j�%�SR�d�J��d�*m�r��D䆺�元��-�v��:#�}5st6hN��Cmh�����7�_�����b�p��yJ2���\����e�\��>ZWݝ7�ǛƔ&��8J��%��GfU)��=f�H2Uf8��z'Y�k�O6��{��J%�[��vYY��<{n�٤<�n���K�l ^�'D��^c4�VA��� Lڶ9�" :�*]=����Y�ä5;`u����Z%�����_Wa��u��3E�Z�z�.*K��+Q3�	�a���֝��I�PY�.��8��T��&��#�މ7g�4�L����XU���q�1�=��v]�UNBf�d��t��4�U+�4�.z.P�Ő���;cl�{�Kqu�W��4-�M�%�_5�����M��BG��.�S%�r졒:���B�w\$��gMv-�V���ۇ_j?K�� Hv����;z��Z�Y#�����@��yy��t;JH�[�F��F�C���z�WM�A�M�)Hf��4n����ˆJX�)+�(=t��]ۧ���H������)��GZ5�u��Lvc�����[�;F9)�J�d��)4�]i[7���M��7�t���������x~�{����O�����2��Q%��l���)��vԒ*�]1<���b�b��JW�`�}mȕ��N�.�j���w���������e��싨�����]:u�!�u������ϝ%�X��k�9��z*�\+2_vu՛����c�jW$?���e��6�p�U��r\�N��)��ۑ7W��u{�*��e� *-Gh^�W��]n�vm&(�s�h<$�.�+�&0s��ۡjhn�,�t�\�5����7#UҮ`\�a{�;��	խ���͢gK kE>�[���[�e^�/�T�*�mV*�;�M����[3u�=e��@���2�fu���������T*�]'��C��a:�p��{t�w���:����&^l˻�T<��z0)�U�K�d�Lm�Q�@����G{��j7�_֝���+=��=ԶKu|���q�9�^�)KWE���M�Y�ɐ���t�����Fg#��%��ZOax�ju>9����%���v�7J�R�ITb�K�.��/�Z�n)�	��.�Vrr���=(@T�R�;��yor�+�D�KRyJ�΋ഫ|M��ާ;Ij��Xrw����T�iP��j��o/��v��Ū�D�K�>6����܁[�N:<���{.�C���7iEs��EVZu�M�h�T�ù�9Cv��֤v 蚬��1!���a��.�X`�}1l8^�pԤ����Էe �N���hG�����nd���+\ڲX�3�N��v�F�*Ӯ�Υ���eǛ�TN��{���Q�[�GVR��#�q9ص[r�dUԱ�Գ�4�Dl�W(�Qd_m_Ae)m��%G5���5��|��=��\����N��"��Y�/i+����tX��iS�����T+��μ�#�ך�6�T��F�S�G�͒�p��n�U��Z:�Zuݝ[�f�Z�|�[w�w!�]��R�����q��,׏4«�w-z��ܲ5���B�b�L�b���̮�U��z>Ou��ɵ@����s�!X&f���y;��:�skz�C����ұ��8>s����@�%mՍ�Wb���G�lĶ��z���(p&�Q���5�vh��nUGMI�٨�u�j�)y��k�t'R��˜2���
��l��,b	J�Y�4�S��^Ӯ6�
��OU�uk���d˱\�Z�.dݠ"M5ӻ�p׽�'6��(J��vb�*��x�z6>$,z��m;��V�F*E�}�p��f��p�w�.�s�}0�6P�ƛ7���n)�Ta�5��^�K�~��gR��
m�aY�&�P�u��{ai&�5n���wC��k:,��W0v���5_o\5�E)�����r��(i>�Z�����X�[�o>�-��K���X����Ȟ_��mvǜ�s��ݝ7Ц潧�Hܩ����Y��=pv�o`E*R)�����.�t�_coY�J��S���	7�Z[��I���8~维+�Pyӯl9�4vX]t�&$��I�;�7��w��%���9�])|e�����:�8)$h�K��'K}��Y��q�̻���4�,�ѷ����k�yhj�ui�!�$�A�W.-��j�~ćgV���)4���REǮc4���x�Y0��I�����:�;5��t�tC�ok�D�$O`��Y�.�ٶ�a��L��5[N�jч���mv��Z�بh�۳`D�mv��gZ�8�}N�u��pv��ʒ�Y������=�Ku�����<���.��A���R��[u���
�xVz��3٬ҁyX�T5:CN��8�Y���3� [K�V���Zۨ+*Dʍ�4X���k&�2�jvc���]�.)�W���p�	�FoLe'?n��{�އ�s��q\d��E����>Ò
�2�����G�J��<�>c��HY��m_Z��n��oSI�t���L�6��\�ы��J��G�-a݇[�}�Ϲ�6�"�f�Ӿ,�
E;0޹k�5ˏZ�R>�hӮy��вf�-�yҖ��T�� &�q�$w�+pS��K�K_-Aٓ�ڨZyް+-c��|3���qkdC&Lӫ�7��H��5�'��x8J���;�"9!$��&;A��bg�Eueh��7:X}�3x$=��&�ld�
� .��(���=hwwH�*t%u#�y�oa���2t�w���{6(f�x���H�9t�z�^����B�ǐmvP�]��n�oj\q�Օ���J�8gEO�r.�����p��6�o/�֜��˭��8�$�Ģr�=�[Iû�fs�׳-,-r�),"�ٺ�w�jf��T�N�y)��n��e�}u�]Q*�e6��/6c�+�]�U�C��.*t����k���[3�`Ua	���Ւ+q7Q�4��0HH+���1V�:�//wC���%"{����"���gc�2^s/B�G$��p���w~�Sd��޼�j�I%͗�l��BF��1ȑ2�S9�T��w��z�.$,�t$����  ۅ��;jS�#�z�q�RN箅K�0)6���x������2��]:�}T�
u��mZ֞�M�}��:��g�R=J/wz^�Q۔��|���R=�oKN�2���(�K�Թ�4I�S˷.B�[�����yD'N�9b�m�}�S�b�O7+w����sD��S %�����L�;["ϝa�j��4op�X�p-�Mb�6vݣ+#|�u|��Ma���T�	�m�M�����A�� ZO5��j[�ӵ�4p��jn�m�%l��_m�`=Z�Y�b�=�c�C�暻0�in6/�Mo+�6*���98�K�9�̻[ƶ��+$l4FSt�:�����o�W�g���1rY+�e�J�S��sZ���GmsvB�cQ�Մ;FdJ�ˈ֧�k&=ʛS�=�N�c_m�ݡkOr�Wa8��q���Y`]�WWt�|����.�"�C�ϻ7S�R<*�%Ӎ�3�}y��n�]��
�m�y���]D�
���P�؂+�D#����Z:����i-��OX�g�*�wpjF��Khfw^��
� z:�R��4���\�uN��gl���(]�d&Waff�6sѴm+�t�A��Ⱦ6�yJ�#W{j���KQ�ІA�0K����x�ą4e\�J��Dh�z`f���j�HU��v�)7r�[궭f�a��\��M�p���Z���ub�f��o�w}݅�&V�u0����Hf.J�XT��[t�V�Ì�J���]X�z�x���Kcߜ�Cw�.$���G�(b���v��uF�p�;��[q�e�zb�8�u�+�'dޏ6�]��_r|TԦe�t�?��0���A�+�����&;���b���Y]y��đ(�2��Q�q*R��[��_Z���MO�P��J�0�
5���D�-d�U��#%=]���ފ�]jw�=%N�E�QϮ��Rˊ-��4�uַ+�+�����A�-�t�:��r��;+Q���n���t��b�,��˴����Z��E������r��n��q�2�T��h�}FݽQ��X���f���:�H�,gC��H�r�ܣ����[�;�b�#���--��u9r϶�K�>����a�v�ʣSnwV3��󔲹v⌔��J�Z�6^m�u��v����Pݣh�h0��U�������3�GkB�+:�]՚y��:)���#k8�2n�s�*��ʭBζ�D��9��=F�7�9���ww[��$h�LH�r���XT1%���3(��;�{N)2
8�B���9�<{7n����9��8��];�GV8q�Umd�y!̹�єۈ���_e˳�v�ۛbP�����J��D�ק����v�c.���_W<W!�����->�BP����G]˱;�*��l�2��J�����[�=�u|�I�ڃ�Īq;�k;hnmIV9̶����9��ּ�ʢta���5�i,� ���MT�]sJ��K�va�ו�K��k��7J���2�V�ˌW207s���45�� 3�\�����Su,���}�3"'���=;�+�	V�r/�Et���w�Ի��OQu'����o6���a³�ۥ�
�c�Wws	��-�8��s�n��8^��5z"�
�Z_I�<����n�r��b��ܧ�PӔ3�̘Zʎ�Y���[�^y��R��*�[��gb#0@�D�X�-��p5a�c*C�a��ƍ]�s�X.�cx^G�OT�/[���wWf%�:�R��m
V���E:���P��y�⅊Z�]��!½`Yaҗ���_e��v	)��z�S+F�(�m���Ö�
�1/�ˮ�0a_��xAʵ�C� ���;�7��y������Of�)�a��̮�C=�&���b弋�Z��NHqo��O.�t�Q�]���lHV;^��/���jWf�n��6n�/��Ӊ��"l�"���_�r1n *LrN3gC#�a|�������(9�{���)�|�i����s��.��N�K�RQ��V3յ���ȶx��+�i��:uC(^��W�KJ���MV�;%�#��+�`���1���}�LOs^��j�;:�b��j�H	��G��0���v9�,�n�
��h�s�]{L4Y7C�8�Y}E�lYijm�3��k�2A�av$Ӽ�Yr9l�r��t��%�Ry{���u:nK���Γy;{v�d{�� v�ج#�l�Z�ZK�6�T�y6�z�͂�l��,i��z໹A���k��9��f�7אI���ɺ�93Z7��O�L�W���>��,uX��$�G�C�]1����БX9�eG<�GmU��NTz���u!�I�Xp���a���闎��J��U�Ӛ���E���;���//M��I�.4#�V��|�V*�!�BY�W@SُpӖ�(v9�f���Paf<SGzB������#8w��Xj�6���I�zv����o��βMgع�ȷ�U��Q˝;n��3��uqd���ѥ�7Ԟ˾uv�TW}�H�Hu�%�=W{Դ�{��.4�ό#�+�:��Z:/r�����+[=�t� ����x���a��p6�r��	��n����h_����RȾvJ�F7ͭ�[��B�j���RfU�`w]�On��7&�]�!:��Y�����*7I���`TW��s�0��������R�*�)��t�cUqt��ņ�&��o8J9:����v�Fk�t|MlB@G
�k�7����(m�ґ ��L�����E���ۚ���4�c�������jG2���q�G����Vs�3���)mvf�%n\�yJՈw��lE,^WU���
���Q�3�k�,9F�9�t�J��J��^�,�o����
�D�BMd�+H:���BهzˌE�ڧ���r��æ���X��{�\����[l%�T"%em�C1��K��(��-_�j�Ծi@(�´ݦ#�tsu��ݜ�k2T;r�W�ܜ�� y��*���
r�Rt�U�D�jPU3˫��l5ώ+�q�,ͲJ�V����Yܫ.۷G`�D7N�Y���{1v� �9�cӭA
ĺ�3�ne�,���\6(AB�;1H)w��s�L�y�j%�|��t8��[��j�!(���@p߭�T��r�N��C��bw��KڰH]'x:d6��Nbn`�@K��X�9��+n��`�*����ҜQ����V]�8�A��e��q˵��er�yX�Lr���NL�r����a{w�/J�<�}�r[a��qr믷�Gtκo���ܩ��V�|>��n�TzV�oF�=]c+�$F�{��v٩�����pe,��wP��B�dū�����*������gi�ng-LM�.��w�J�4�)���r�w*�69!�FR<�[Ht���q�p�%7�غ�(u�p�[ٷc2�
ް�H"�N��}��<�:�� �eդ����J�q@:�j�J�h̢$�%��+h�{���&�4QY�9MC���sbV��:����#{�Ǻ��ƾ���zqک��b�{pr/n��l���4�W���u[�b�����"3u=bg:eK�#��5T�MWt�wlhv��vA�[�RYr;�Q6�њD�X�4I�h�y/�sp��;&n�E�F21�a��4�Jgъ����}����nʩ4[�|�ձ� پ�Wu���`����&�:kr�{�ƹ*L���yZ(bU���3�֚�:���q했�W�T=�(�D����d��n"0;X��ֵP�MWU�hX�T�dabg�ò�3�`8v�Z�N|T�5=�h�V��u������!r��,���;WK6G��]�v�ItB�cæ��PJOY�<w�;�]��+��k8e��:Z�&|75#T�X�BLU�ci��ל��SL��;3�xv3S� �LYY)'S;��v��8镧�,��	�'�S�;�ٸs���ɒ{p�����������2#�Y��7G�k�-rj����C���b���]h֋�k&E&J�΅��I|hݳ󙎵�+H<1c��WYQ<�@�����ü����V�6�;�G�S��$j�rFC���e^U�i���9}
+^���3��Oce�>�H՜g3�N�g{w��V_g;�6a̢�#���>��%�N�����l� bӒv�"�ؑ�|�E����+�oP�5pit�$IY��C��u���דr�}���[zSL_c�ʂvI�,�& k�;j�,�Wt�n^�6}�3e��n��X�f�8�l���'G�p�d�yМ|g)k�0]� ͣ�RC[F�t:�*�5G�pW�d��ht�!1�䑣pBie�S]��	8`1_Q��Z���(�/�ngM®�k�f:��=�x{����(ԗ1|ٷ�f��k��*��c��Yw��Tf���/���,�����y�yJ���[�:����>�ʺǠ�f�"k��� ��˭ �8VYgE���𣹯6��x�U�9�b�j��9Fp��f:��3�ju�Kh��B<���S��*u/xod�I�5�A7�=�So9'�s���I\����0S��FU��3(\�VH�CE�TSG=]\�[��	;K�ep�L%\;�s��#&^� �����Fv��/���=Еm���*�7"���K�b�(��S]��\ۭ|�F;�%w
8��h�x�w��*ŨGQ��k��єẕ�o��2��ܶ�N�`�*k���k���& ,^f� ��@�n��;	|�@��x$��Md��K�8䛸,�>�+*e�T�J�����4h�F=�*�"H��e:y����/�^�*VfXP���`��]q�n�ܝ�u�*��"J�(<]�,
|�v'`e[�T^h�r���L�ťG������7T��y��E�Í��e�f�-��s=������C�N��`,�Ȗ�}y�s(!{B]vs��G����5We�qx�U�6��ͣIs��n�
oo�d�j^����Pd��7���_f��9�����J��@r���Ec�U�̮�Lp�v��1�'73/�L�a�OPވe��ʖ1�oV�(���μWõ�Q����_߿}���~�s�:��4�M�5u�s&i�&bb�`���gM$CZ�AMQm���֘�*�l�TUT�CW6"b��MMD��4M3D�1<�SUCELU2D��F6�j�����
�j ���9�4Q5Z�����%�cM�5V�E%D4��UU4�U3DZ�LU�r��*(���)����������m��*��h�kcEMDE�Q55A1UUm�8�\�
��g5QKEU5EF܎T�؈����5L�Dl��(�X���"�(���kX���*&&�-�S0�7#AUL��s4UUE!F�)�5�d����D�AT�֍m�.�������(�����"`���m�� �䠡�1��EZ1$��b�&"h�A�����

 ��(*�-i��gU�k��?|���:R���P�6���u��d�|�'�An;|�/&��L��J��9m��'V:v�C6��\͔i^���{:{�sd�"��"��*�(�`���D��mK��3G�n^��w-��h�����	��WV������?_����}c�cB�pﵰu�A��R�G����43U뛗��� NM9�@r>�������%b�V�1p���5�ϜހAd[�ƶ���(�NqU�:=������<!�'#{S�U�hf�D\44�F@P�ѓ����k������J��5����Nb����0	t�8.�K=����wȍ��Ӡ""3��A��;i�y��o�����8��U.�^�'݊�3��B�3��U��{�e�[�=�+����sK8�a"��J���Q8+���io9��z[?���z{'vGG��E�>�(�N����'��6B	�V�[��r-$�h+��H|j6�}������rX0DM�ŦݧXm��+��HB���һ�J^��k�ɭ	9ip{]t��\k�>��|���/^h�xŒz%��ŢYz_�lO:&�W�7��'�_[�7���S����}�w��ܬ"7Z��5����e�x��0�颺����e$�^{���*�\�4M��:��qfo��*�ƈ�D9��09�K���S/�aV�5>�;���Qt�#G������e�{!�cc�l��S[�թ�q\�Wp����V����@��|��c8):�.:29c��sz�q�e!@U�(����.���z�{�_�E�Lu�(�S���61:���-��ʌ��wo]��q,�]/'u���L����z��RW��B'�-�Q�u��{�Z��I�hӤb�$�o�A�Q�ʖ6��|*�"�v&�<GP�&.Vӣb�R=|���he�ɮtg���o�YV��u���ΰw�_ 0xT�Rg�'��0�����[Yb�s;F���9�;���
�H�Nm������z���[�d�m�F��j���$��Gf�Ų�߬�mnr{��ۊ�Z�H�ͧ��+�aHzhj���rwh��>dз.�3^�d<� j
��Et�p���\Ď&�o��Z������E���B��>����8��]z;\Tb���9�Ϣ.�oD�J��ya&X?m	_�H�r�֢"�z�8��g��ds(K>>��)X�l'۾[��Ye}������EV���f��Iw����S{����%��ސ��Q���f�F	�
�,�b5�c����<��n�1��m��Z��Y�^#ٳ��s���]K=L��9G�R]�X�7�ţ����k39�H�uf��̒:�7n}�Tj��<'���iϮ�Ǥ�]�����,��i������W��Vu���b4���]dU����U{��K�:���I�y�j/���yF$�7���E���/<�FLQ�"M*'G��t���Q�f�`�N�l{_��8���K�}<ǩ��\C+�岰Sw�E����
�A�W�Y6�0��q]���p)��ꙺl嬢͊R*N�z��t�3�D#�ڰ��>�"�t�c5���ғ1hd͒m�*"@����C��t%ئ�b�K���=����sv܎��'��R�$N���䦮�!pN.N��x'>2�)V�pc�Y�F��X�X�t�tXe>ZRcpb9�k^���$-{�n��IS����>*�7�W��8��ׯ�/�c����1��tY5\X3�,���lCs���W���Eث�	t ���.�Y������9H���ܛ	��,3l��F�!�Hq���};	b�i�Xϯ�-nU��Am`�N�j���\�÷=$W4�Ѵ�j$X͗�I�D�d Ʌ�[^L������W.f��.�t>���,}���ծ��T�R���Iv��6�z��͗v%G�cn�w��WiN�tN��n��zd�Z㗆P�]�١�o$���S1`*Vv��k;U��+��Wܶ;��/�ز��YcL��ۜdi���|ӌ�����CMn����gy�}�wzF ��)�ˈ&��G�zĝ�nk�Fv�}��e }�	��vPY���p�=]��q�caqmU8��3*5���1R�s}������Af���B���&���c�V��ZUb�^����gx���U�<z�&����� <�v��?5F�{/D計�x4��|+�,s'�8,�Ԡ�=}���{9��rz� 0�]����,��5��ڿu�u�nCV�7�n�_h��˺DU�NV�oeF��M�=T�CS����h8�2��I��=5:�G� ���U�6�PG�2�w-y���+��'�_�<�+=������l:P,7)��N��QW���.?s�K��/�+�ż��#�g�^_����~�[�|�k[�
���ƋP���=�+��Yܺ���w+w��s��.K48�J��@C�
٤��j�n���T�9K��P��н{��y��!gA�`��'�k�uW�P�@g"O0:a�����Uۀ\<= ����ʸX�̾���JۼSwF��0��+K ���6錩F��ڲX�k;#����S]t7nS����IL�����腪����ՠs�l�y���êcָ�h�<yQ�C8��df0�s���1�WC��,ӹ���C�#ͧ1��]9�r{����OU��(c���4u�px{+�^����Bg��W$�[Di���!.����(l��ǝ��A��p8�qt�o	N�#	�)̌�ۑ9��31AL�iT�o����]f��	��
BŨ�o�P͎�҂�+Oޮ�8��0q:���W>t�]o������xM���߾	Vm�'��N6WZ7�C��Y�=G��j�/≮�mS���]�+K]������ڢ+E�t�>��t�k�3�8���
j{n3ͪ�1��ۊ����Q�� XQ�t�{��X��~���@��Y�ϩ���v�q��U��Y-j�;Պ���l��}�|u��r}��>�]� �֔�\+B1p�B���S}iӏ}� ��Y,�|��~���w� ����eo�݂��C4�cA������YHG�z���M�����UT����J"�z�.��}���{�m�U<g
zs��>B�JQn��:���.�/|UpT+8�7�)�Q/Q��i����Ar�ޥ^�"n[E6^ln�p{��Z�*��V��;��f���rt++o��[3�C���tC+��v��܋��d�C*�£��Z�D,�p�~&A�2��Ͱ�\܌�=�7����S�6�S{//��8��	���ͧ�҃���_�#��}\���{�׌�������-.�s�BC�
K5�
_I|��k�7l�|�O�=�@��Vu`ў�o�Ɛ��/p��6W?�4��� �����	ܕ|+�3F��b�Y�=\F���~{a�R�zr�8E/ONTL��u��Cʭe�wEڥ�}��#&�Ip��My�o�5%��lP��/�o�_��:k`����������6�w�J'.ї{��-��e���.:2,r�i�4��g�^r_��^\�Ѹ��{jz�P�@�q���Jt#�8buѱ�[W���{*5��'���ƪ��-�[y��6��X��4!U\E�K�z��b�˪Q��PE�嵠wN���`�)��㐺+�k��.���wT�C�����%m:3�#�Õ��h�ȹ
;V�{�E�ׯ����O�u�=~/��Հ��E:����w�:�G��s�|�vc�E���,<�d^��:=K�>��	����L�m�G<�EqI���'񵢝8YC������A���������otʃ�j�#C-hJ�^�7�|.��T�h��o�gK^��R�R��_TY3�7�H\��]����)Z�MGx�reky�+�֤��ҥ��",n]�M}����%p��UѣIJw���c�}�t�X&gn��K�$���=!�,W����\�x�#=�|ɫr���l��p�DGlߞl9�\�h����}RP�}�D��ZH��P�d�8����G�]z:���V2�-u���^_��y"�d��3�9�+!�(���j"*��qp��#9��6��A��3x��6�`�U\��c�W�jf*�Y;�d,4����X$����7���YkT�-�/R��H�n�Z�w�e���qj�i��tY=���y.8�U{�y�W�wK�{���.nDs����r�}����g��j�ʴd��*r$�=>���˥|3�q�Z��+��Kj	�|��G�l���_b1xf4������)��]�o�W�2T�W�י��N���*g+8�ܞ;�}����</��Gkͫ��3����uT5��w9�.^�b��$�+@Ti!��V�o��wM�DŅR�"���5�aٝ��l[�V�ۼ9Mdࠠ�~u�:����]&B%*�lA�ef#^������;�w�օ;	_�.�YK� 搩K�n���"p�8��_����څX�i�<K>�8���U��m>I������G�^U�����O�v ~�����+`��n����
��Ρ2(9��r�s}}�5N$�s^�9m�0�$OH]){܂�s�=�0F)�Ğ�� 10�wNxg�����1�t�5�}�\c5/nb]7ɢg�ֶ�.rg s��m�}a�@2�I�6j{�r:#lv�>���Z���ҵ���3�n9�r��<H��]nM��t�d���R�D�Di���v���;5���r�2%�q&�AJ��X�W�K�~\�÷=$sN�N@�`#C��I.f�nM���l��+I�����E�u��^�vmW~Qa'wP0�y�q�O�M��n
��\ǟ�[@���:���>0��o�ُW
���ؼ5�ŵT�Z95i�K�e�hj��[�YVx0l��yS�B�Y�m��Q����Ь������H�R�k⢇�|��Ά���0D��s����Ps4C�^��fQ��r�����^����zz���e��;<J/�d	XՆ��e����������xߠU��C��9s*1\�I���ȭ�[ou�3u�be�غ�P�t��m�R�ppS��ʞ��k��°�.�%�X� �7%>��`�y1��%���GC2�&���j�~iY�
E7���]�ﻶ�t��}׫uԭ���d���g;絼�Q���٢e1��y��~cޣ���O���\�Lc�t����p�Q)��Ef�BN�B�]C��MS�T�C��pѭ4�s��2��1���peK|`�pW],�� ��Dip�K9�=x|�롞 ���Je3��t5^�W�s�j���v9=mk�%g������QZ�O�[�>ӻT#5��c��W���p:v�fW�yl��O�P���8 ߠ���0��B�i"�Uʢ���i��5����L��(r���{F��T������,�z�����^����'&�UUk.���#�e��bl�=�ʐ��r`k�S�sH�)�0$p#N�^do��F��7]�_�\���7�������b�����DEiH�9����^y�W$x��o;eM��,����8��91"Nj����tnB���젗[�[VY�-���ׁ؄�*�UI�}��U5�"�OARS�����BNÓ^���U��P�>VaÎ��},�u�햕#�%����^O��ַJ�/�`dBr�Nh�0��yB���ӂ�C���5�[��3��o���Mm���},����Ӡ	����x�'e� ��Y��,��i�7�#��BU"�t�т���M���`�m��o:	�e�H�1�s����pa'ԕ���l{��>V��b�ăB��6�0��㪎�[�T���v-�30I��7�����s�A�:��곿n=[
�8���f�=�%ؼ=��U��Бҏo�37;�7r��چ)p�:�J�Y~�9�i��9��C�cG��Yw4��DW]K�s�Y�
+��1(2.PfTc�>'�wKf�߬�����u@�hf�D\4�H�*�q�~(Q��ݓu��C����}�z9c:�Eְ8�.��=.q����{=���jS��CN��8\��.�{qrI�a�.�\>�<-����5�)�;�c$��\�w׍�#��.|���6}�.5e!y�S��{��bI�E	�U���5Q�JL@ע�Wuݘ�}��~���l���o�V�[��l�'R;�������0u��f�Yon�Wd'H����9�*���+A��-/1X�KON4��k�� �O2輫�F9^�Uq��X��D�ԭ�h�^���
6�u�	�U�7�{`��`;�$�;��7�}�fs_��0͈�h���c8)����FG,t��1�Y�}��Td�ʈ����N��M\Va�<v �d�+㓫�0t���:���m_�w��p븘����P�q�b8��������p����n��o
ͦç�6E�(S������`���C|R�ʼ}{��bƷc���[0��kU� ��vn-/���ek�t�Yv��}׵����s	mކ��IP�&�umc���<��Ϧ�=�&��G&WCİ��$6Q�B*�kR�)�Q�ݻ��Y2Th�F����c����6�U�a�mu��n��ƕ�'P�M��u��㢒��|�d������ﹸ����c�c_`Ң�X/rQ���Z��L�i�̔e��G����V�ڥ*b-�4�U|2�Q�f�/��4��SP8ٮV��d^&�P[�#�J�39����^���.�`�|hP��!pٙ�S�Pī9'Yܷn�=�"�Zv�Y��Ec&*����j��2�Ɏ%��%���*�I|zf���q�j�vu��$t{s2jz��3ZW؀U�b�ͅ��N&s�c����E�΢l:�3�.��w)��Od1e�Fk�gJ�9񅑘h�����r�Z���{����<�VW�P�E�}ي�+`�����ս��Lh>n��/�����仡��,F��;w�S�0Q��\��Js7q���%U�#&E�(MvX�:M�n��������20�ā��%l,��o�i}�we��#�Dj޸���7�|��c�Ss	T����5Ԉ4[�����D)Zn�����m2�y�s��WG׹`�b	:fD���n��9Z�(�}	|#K����y�3��!O�	�&�gS���ϳb�T�sC�]ʈ/y ��q"p{5���U�r� {;�]��}V̎�[z��-�i^���Yw���5���@�9%:_R���+(� B���t�T17��ձ��36��y�l��q\
��)���p�I�X�nͫ�tyU�=�mn)���v�K	׶�+�Oz ����p�il�Ȥ��p��z>��\+:�m�nf>�A�]��.��cRj `�b�����mLJr<�ti���oN�T�J��Q]��T�A�P�J]17�Y%���}�`]B+Zf���Q��������9�bUv+j�)��)q��;87�5.�y��b
-�+R�R�ޭjs,)6�I-]�R�-\e%�bi`�yNܹ���a<!kk.������lPq�?�%�Cx!���4u3�}"D�WR(�Y�2�,��o��t�Q��].���]<��y+��T�<�1��T]��w
ڽs �k#�M��3k���EWPHs����T{q����b���"��.�ȔJ��B�� 5+N���,��@]��k{s�oǢ��HW&֛ͦOMdS�<
u�FP�6�1w4S�:6�	h�7�g.�P�;d���dX�a<%�m����e��a.�{@D۴�- 䪸]L��¬��I�ㇶa�8�y��*��q[ȣl�^b1�)��Z1X��Uܫ�s�ms�U�[����=����U
�MQDUUUUMEQT�ES]�5cURE�j��`�X�cUQHTD�b�J��T3e)(�����b�J�"���AQ5UT�AO6���jh�J+Z"���.AˑE3QDk2V�I���EEEICSl�4h�����d(����fJ	�:j
�X��mb����	"
bi

)�*�����"&"�f(��E���AQUM4EH�m��'��͛m�RPkM�AD�TE4�M5P��UTUUEQɢ��Zb4��$�  ��JJ9h�������b��Z��kK�`-��0V�4�i��&(���V��X�����5kUF�5AD��l`��͈�*�h��%9�EZE��*��e�����*�*�j*�"������X��#}J*պͮ�oV�_t�����v��Sם���lnQ�℃N���$�R������.� =�u������A@���G����A��BUy��A��9G��i����u}���J������=��?w��������p;����~?|��zc�0 ���{�2<��0N1��yj��	S�G�q�#F��� ����}�~����=��;���`�{�S�}9��nM?��c�!C�9v�e�M=y��ǰ�����S�y'#�'���>BU>î�|��:�ٻ���=����5G�	�.�a���z#�r^K���;���g���;��4�wݯ�s�P�A�O�uu�������˗$��,�]��rt~�&"<G�Ip:���w�7�:����^�Š� }���",D��~������?y�O�>BU'�������yοa�G.�����/�ܚM�o�y�������+�^G!���u	�{��X���T #õQ�~>5���`��~�0|G�>����O�`�E!s���]���?��O��I��ϝ?���$���$�y!+��t�P{����x�{��<����x/��	���{�>���`�ç�x�i9x>),߯Z%b�� Ǽp�. ��y'��U?��ш�_��]��A��^G*�~�:��5�9���a4�.�������BS���z^�����\�X�#��=����:�NwiVfv�,V_����f��8Tc�b�?#�z����rNG�>���}��n_�A�K�u�����`�9?%���??߸���4�w>��r} ]W��V�� Lz�=��a
����ߚ����p��$���rz�C�?���}�?I�HS�����wP�~~���'�}���!)�����=� ���|���A���^a�)�|�"��(�����������?bɻk�xj�����9��}�a�΄�ߥ�����z���������O��:����K��9�ː��o�d:�!��=��S�;����_�1�1�T��Qt�K�&��h��k���{��{������_y�����z�{���y�����|�/=��{�w	T{.��9������~����^���u%���K�8>A��y��>���} =�m*"H�b�*{v����ȁ�8��wih��r�[~�{C~��z�s��Q'�.�o��T�����/��rsօ�ط�=5��2Mc�G!��QE�:��ZtX�
B܇n�EWR�Aμޙ�>2�S	�o׮�Yٙ��+�ڋq�#��9�F�87���� &U9\������q��YG���u	_����<�4���/p�>|���;�e��|9�4��NG��G/���:�c�9G^��;���?�f�I�Ht~���C\���%~{���>���年)R�i�{#�Ǽc��>�CO������?��w��J��=���u#�����K��ܚ<��=ǐdxD ���܅���6�iV����?}����?�|�O�r�������?a��^�����i4����y ��޸W�G$����.�����z?�����;�K�������`
���=0==�G}8ށ�^�����o�:~܇�{���&�C�r��s�w	O���>GRr�CA@QA�~�r�-:>��^C��^G �����ܼ����P���~?���� �D}�H���S��xk�'���O�t�������\��}=��p��_��s�{��:��k�w�N�0�z� �2��:��?c����&���]	A��0u?e�����S�~��G�;�v��G6o��+8��ˑ@QԜ�O���9p���w�y%�{ǯ��=����]������{�=��?�ӣ�N|�hy�c��^\��9|y����˓��9%$}��Փ����}ٯ��[�r�DH�8&����u��9�w��y�:� �y��?t�BS�o�~��>�PrC��A��޸_0�#����8��}�&����/%�<�w��#�D��W�鮉^U��o�:_��o�=��;��t}~��/���u����~��y?e�>O��~���M>��=��ZN��%w��I�|��pr=��
(?������%�����s���x��`���۳]��}�B>��y��s/<����u	O�;vy��r�?K�O�t�_�O#��_�'���������>t|���|<�ޗ�|�	��o=�y��uC�h���7��%�bkj����$zbc��s���BW~d��sԻ�>���9'#��v���)�?I�u��`�%�c�z�����|�q:������p��i�.�n���>���������F�<t���v
ns+ZQ
9Vs���VkF�b�Ovݛ�����!�a9]2z���4FV�@�(�W"D:��Z��Ttؼ��Y���w�[w(���W�;n��<]V��/��m���M4�H�{{�	ͯ�곟R�`����c�C�?y�A�i|��#��xi�.����߾�:����w����N��'g�C�r9���a4����}y��}��)��w���}� ����I� � ���R.�k�Z��؉�x,#�����:�_�Ɠ�u�I������=�BU�_���8=��%��d����]o�|��y:~I��C������!�|�� �y�`��	���!�Q��u��9�����b���$=�u>��9'/ �z�T�P~����w	{�������{/e�s�	O��y�����!*�����N��� >x�/*�����Q��a�0���5��U��f����#�"�'�GU!C�{�uK�s�	���\=�����u���S�a�����O�����u����.�?���w>G�r<�羸��	O�}�=�q��r>��o��)؂\SǗ���w�^�G�����e�`�ב�vs'PF��Q����`���:��v�������K��0��{�w?%�W�yԔ��u��J=���MS��x=C�D��;�����8.%�j��WB��&��>G����}�BQ�����z� ��NT�ۣ��/0�:9ë���y~w���?_��;�;�BU�/g_�t|������?1h��>��J*l���S��Xnz�>��=Ͽ�p;��o�~���y�(}��.I�������䜟��~Ο$�rN_��n�*��8���9	y����:����yy/ߞ|�<#��g�8�#���"j���~賽��%Q����/��A��}�u�{/*~�����9=�����������������탗r�9�!����v���:�ΰ�%�FǗC�>c�>]�#�nV<�l��+���Or��������{'#���z#�%=GÝ{�r?A�@o1ʟa��?���}�N��C_c��x��u~O�pu�|���G'��m!_�(9�DBXK��l�7�f��Ϻ/��O%���>�]�IN���9�?c�rO$�o8��~�A����M?����z~A��!/㛏�>�'��G��p�O�4����`������PT��!ULQ�6��)��.�D�VW�e7;���K3��������b��t�-����$̔�;3f��c܏g<���{x��q�b��^Q�kZ<.�jΩjg�S96ea�-\;F6̾zh���=�9b��� �m�ZC/q�1��4�j���6T[{���-N��4������u����TwP�~�����A�9�쿣��]�_#�_gO��y��`����t�(���?u�`�a4s�{��9>�$�M=��rN^^���y����Dn���/�{��@ }��E�pw	u��prz��P��͞��J}�%������p�.�Pr{���1�^T�?���y=�翼���]�k��?t��*B��ϝ��:���w6iWQ��#�F��^q������y�=O�������������<�T�r9���͞u���}��9����J{����>��I�w���O����Ͽx|��������z�ձ��Wox�=����� ����:^�g�y����t�͠;��u�h������O�w?%�|6o�RS���z���rO�v�ʐ��>�#������M?���=���������t�k�?�w�J��'��>������A��~�	�I�=����p��?�=�>G�������ɤ��Լ���w���=��p?��? ��>���GS��j�Ŀ�G\�%�(��!0;ةN�[T�W�����}��?ׯX���7��ߝ���rG#�����'��>~�װ|��_�� �d`��+�/G}v
��Q�y�ۻ~�Sj�����&-���D�
�ޡk!�NQ�zOB'3�Dp�k��NÁ���v��pf����߳����V��k�-�3ƀ��A^��Ӊٟ5�	VB��|�31���EȲ*��Cmc�R��ٿS����Ǣf�ZeC�{����; �:j+:���2".�t�6���֦�Ț3&�KJ{mӁ�.�vzr�5�>��8]#�,�^Ӷʈ�_Zu{�~^�Ԇr����c���؁.�0��km���[{�F���;�J��D�_ѭ�����V�'z��zJK\�օ���|��4�o���qw�B��*^L��l���X`��^j�YۻRR��ѱt��H���w�����3��p�n�`]7j;��?U[��e����-S�����H��A'hL�s�sPȵ$��^��MT�/�g�4N�pw�԰�%ᔽ�R(EA�.֋�a��a�cS�8["�XPO?J�62y�&mJ~+�(h�厗9�i��8ϲd6����d���7w�{�\���P �#�H�;<���^��c=-���w��dM	V��N���Lg�tq`I�X�>�Q�bw1��y�Q��#��R1v�Xo�gj�RdW�v��!SG���C�P��ۭ�������=�;&2���Aٝ�$��F��P��^bg>�{�b�ܪ5�h+�� `�1�$*�&k��	��=>Z#7���5��iWcauZ���v��Ǔ���LZ<ɓ��Q�L����L���҆�\��#;v59��N����V�C��Qy��Ut�wh��>d�,A��w�U'1Jt�쫜���%K��8]ɝ/��r"�.������:H�*h�8�t��1�wy��z1f������%��˫T�TUnfL����#�̚���*u²c��Ed�����W^\NgN�a�81�h����ȇ-�ۏ�o���O�3��"&/��@����g��D3��[��m���Uw��1iz���Y9X��m%��Ꞹ3F��8���į� ��¿}�,A�%�'2��7f�|�{*�UJ��/�^��
�E3�����z�b�W�y��%��/�i���͂�-W�M�E	�L�3u�ϩ��{|��$����Z��d$O�f�U�,o�藫�<N�t�Y��~�U9ŏV�c���	���r�~ٖ!\��2��yƢ���#�of��]�$P��p��E׎IӘ~Dw=W��.�R�~�u����ƗN��Xl%)���^3ܨ@�T:�q��Ӌ���PQ���|�P<+��Z���m���(�H}�-
�{Ц�� f�rY�ݥ;���c3�}QP㡒{�����&ct�ڮ�T�z$t�,{T��=�eεu,8qn�Ҙö���J���G��B%*�ns+1�DFD�>�=��Ou=sO����m��_nv4���R���J�b!0���k��k݋U)�Wv�r��U��C���\k��N�0��l��+ �m�D[��d)�W5)�A(�e��8�p(���nY��ޝ�|��刦�oz���r0L�2���@��3np�5]~"��z�������J'I��n�y�p4��!�h�Hd�h@�V���;�U��Ng������Dt����S���gT�Ӧ o1նV���9���;4���Sx">�r9���;�GKf��Č�5��GC��m��؊
m�L��r�F{{�=q�>�)Vmb��&8H�h����7ڨ�����Y�k��O�3�� '�yI�|̭�ځ���s�-}�CMv��>W��e�39הo�N�U�`�M�"��F7Rдȴ�Y�@%׼�|���/��T-WJ��V{��^��>�n�(�`ҳJ���{�\�j;&z�C2�\\-�1���`VN��c2B��h�4����z�lr��5��o�x�����G�JL��,W�[Y�V,r�#<OC^=�HzZt�M��Ң�֥�Ȟ,l�cV*�L�f3�����s��~�VFDL��'ʓX^�
aOCg|�uA/�O��5�=���:�R��<��U:#�tV��à{���'z"y�*cWS�d0�AG�v�qut��\���K����u�aʁjp��+o��F�	�:q�t��s��qʆ�����U������k�l&�I�/	;��g�[�7�Ֆ�V�ќ�3e+w�h��Ūܥ^�W��7+�
Rt�t^;jP�A�k��8�<����d=�Φ�f���M-��ֻyHNKN�:�FAu0tܓ��W%�ۡF�;�n9�r�Z�G#N�/eU
���]�'�%,�q3� ���҃�3&s��%e��[�<=�w�mA���m�
�כ�9k�l����R��t�5�ј�}�J��RY��<Y�+�f�2ss��� =���V�ε�zN������ZA���ۇ&�L{� T���`c�S��O�U�н>��ڗ���zǵ��5bϗӴD�>��`)��i�v֍���zR8�FE6�N�.��3]�쓲N��qu�,���u��	��&�A���.���Iu�Q�-�,�Ѥ�Z=F�绥Ψ�xM�K��s�I��r9U��m�#�ȷi�3_{y��m�!0��]t�{�M��&Oۙ8N�FP�Q����8�v��-6�+�t�ו�{R:����]���=�՘(�/-���K��ߊ p���{�U�V~,���Mx��w(S-�n��s�=�ܫ��UZ��r�h�R6+ۙC�$��������y�*ZfݴD�ԌE�X3%��<��ge�4�h_���j?����9��L�����<"�����x�~{I���V������Ҕ�Y�����y!��ؘUC���=�}O���1j<�IwKl��\�v\���&o!xg���E�!%���2��+G;V���r����u��	�UT��0�Ϻ�Yu-���Ո�JZ��7jf���7{�� �|{����(<{�$ex�"2r����z9~ͮ�u��\!G/,�<X(J�ς1;R�;N���s:tDFe!^�����T�0<,W �����א٪�=3�8���r�����op�}�&'{���i�P����_@��g�i<U�;#mJ�(<�4�8)�b�z<�w��}�:���l���m[�V�h\�(���3�ʯoF�cu�T]<���E�Q����Y�.�����e������m[��5��&�	ՋP\�,��v����r-��d8�]"�!#Bs��]%���){n8Y7Ǹ���+,l���U�����մ@о'DO�O3#JG�&m�M׍ ��FE�Z�qϷ�a����	<��1�/�Ó�t��z�X����@�uE |k���-�-���c%�~�����5�� �8k'!1ʻ���؞7�}!�����K|���V�e��Y�PܥC�ם�ٷW��L��5$�af���[�Hp*:ۭ��<v&���<�òbem:$��ࡇqn�+^7�ʲI���IX���E\�-�jt����6�h�Vz�t2��q�j�R���s��@iс�]��J�J[z�p��F�p�Q�L�&-mՉ>����ά���e)���g���Pw�7��'�%[/&��\F�����꾤U�� =�+j��Z��`��7'~q���2h&렼f�DlZ#"%U)3^�D�G��ذ���/ݫ�~��s�Q�z��Q�67��O����LZ<ɓ����n����-�u�v�b3�I��x�v\{��I�>�8��^��׵^X\�W��>dչbҙ��:�����^9�2�El�a��pߙ1r\H�P�ʴ�~ݕ�v�C��O�������+
��w)��iW7���/f����+zU��q�ܯ1�c�����©�����/w�zYl�1�U�^��B�4����L�wJ'v����-W�znr��z�A�7��ks���E�%90�"}i�1~���6
�}�����sע��4���7��;|�j�&&�f$�Z�7\*T��RGIb��9�e�ۿ8�|E�C�E�ܜ�T���x�u,��	X��$�PMBg�=�+�A"�'^W���ʳ��L����+2���&�f����1��"J��l�Z�8��(p�����g��|����v�ϡʋc�YKORW9YPz�a�ǲ��������]]�eೈ4mg�[�ۻ �Rf7S�M��7]���Ţ�L����tڬF�ْhg�usV�����׹ث��q\����0ܠ��t�9O!v���f�=.|�������pԨ�5B��s�N����3��W�H6�!�M->R��|2���<���RѳY��'
�s�uL[!U�"w̌�y��r�nYY��ˇ�6�o.�4���>����=��{-�����Kmc s��.��&��
.�:��p��rI�7���BO�����zi]���hW��nĊR�h�!)��[ �8
�Y�{a�����-���y�̱4]�C��NŇ���큥�i�˒T:�w���k��z�&K=V�	�Ӆ�~�[r7Η��(�܍`��
�p��y�2.{R[���� �j6�zs�4�m/F���Ϛ��6�L[�^���T��}k�^�;�]��"�v��@�#=UN�# ��c��Օ/h:nY�|�3���J��Q��-�=�V�ө;���>��ѽe��OP�DԬjK���joq�z2�	b�(;Ś&�t�S��&>��Z���u�n��5�+U*U�VE7B[12t�\��[]+���xQ��t�!/f�|�X#�8�)�c��a��(���b�G;q�ţ(��ܰ�AK}Z�,����`��-'�T�m(��Vv�@%DͰ�-b��e+69�7;�V�"Q�I���p���n�'�V!���yJz�8.�=��(.Ծ�O�Z����4)�aI�XyAu��WM@�{qq�˕i���\�4�1�Mb��˹�Ms
]����[Lf�Uz�Ґ�Z�������s7�4ʔ�j����F�̈�X��_a�����߸�x���ٷ�B�.�fD�X���*�Yh��
%]
�@2��Ǫv�2^։w-mZUpɬ��8���-�u.v^f�%��G+6�\=�5�e���%��)�8G>��m�憓��1cUيV#b+�1�8^�Α餚�Ӆ���f���y�rX�m��_�EM���Vm�#�9��kU��靱K�8�v.���wM87*�:�5Υ��H�ʦW6��W&QW�ј��L�O��yt��ճe��)�
�ypiXb��\Ų�\���w��.��kw��Q�n�s{R�)i�4��}uJRz'��0��K�	���=�h^`��ӷV�֩�=]�
2:���f\ɍ���9r���~#�0���%l^R6ME�P4*���Sǻp'^��sa0��`Շ���:.w��?
�wz�5��i]'�;x6��T5�t��oT���8^ӝh5�l��4s/����S�p����.;�}�Y��mYf
5�n	�F��a��F$Y���e�%_F��R��z�v-�[�]��P0�`/���#\2�:n􅩍^.���B��W�Ъ&���k.�ɂM����������{�!�c�6�b")4��KmE%V�6�LZ��IEr1QIE-%ڒ" i
b`���!$PUISA�S�%ET4�TEh�:ySEQIQ!�1���N!�A�I�"4i֢��4��h)
�+Y���U4�D�4D��EM�S%$UTQ)T��ZX�����*��g4�V���&�Z�����:U�US'6���
h6�IEDQ1Z��B��"��"�	���(�-"H��
5�#F�5��*������&�$)nnTr�
�4Ѩ��d�&���* �1TL[m�AM)II5�*�MSSV٪�ֶ��)��M�&���)+Z"��f�F��
)�l1%D�P5V�A��b6�QUD�ѥ�����pe�b<��Q ���[�Ji�֭�3sw��5q�l�J{y��PS�b�ӅA��IP;��n]d�b��������Oܕ��}�2��?�3]����b�h�'n����%[�}[��z|��Ѕw:ͦ7f�3�]��P��ݮD`�1�Y΅J���(�>�!��i"#�VyW��˶yj���L1o]��*v:!\�8��i,=�ci�(�
d��q��DÏM������.�.V��˵���t2���ǆ.5��$a���Nr����C7 �
d�Ǧ�v�ULW���-�+��o����<_��GJf��#)��%2:�ͲZ�Ȏ ���рb�7�n>j��6H\`"	��^���$T�b�͞�}�dzyhh��w�f,�����V�w
���+X�vd��N�d�D: ���E��iL�+plKҲ�6�g:�'enZ�I�PCt�����:���\�;������~uK��ǫ�{R�C.�'�*�_�oru c��։�o§��c�u������!k�
ug���0o�Ǖ��ў�<E3x�.�:������J�!MW�����/��訉���X�^���$V��3�����6�C;RU��U=jPŇ��XF2�	(�ȷ-�
�iM�AVm�j�D@��&��P��H�v:���P�z$��A���^HY]��'��ɤ�N���W�������� nLr�ʯ{w0�� =�{��$��� �?�#lVUi�y�v5a��4�d�g[���u�r�˺I(��V�9�w�ˊ�cՖ��'D����.f�<���ٕ�F�p+�Je��t�W�5ڜ=��soRn�ʙ06ޫ�"�Ӑt��^���+�𦳘��X|���߷뼮%h�Z�$}���ދ,V���=�]:�k�K��D@� �3>z�I=�h�{�M�sc�������VX�v=�
�\�2;%{��a�,�Ƹ�J�g������l���i�z�w�����`��g)�����r��h���2=�W�Z9���,�� ������1*��yn�w��Y�!�"��_e\oMP���o�Hq�p7&מ;�������Z���+��BS܆�!�t��d��u�i�ʏ(�<1utvJv�M�H�s# r�AS%uF���rS9�jM�~��P~H�������A�L]m�7!K���B]nd�b:�z��q���2s�I ǪŘ�xoՕ��KA�sU���գ�Ⱥqv�s����_T�E+��ױJ������(gJEh�f��R�'U�����4�1Վ�X��^�ϲ���K���Be=�������]��ĭ�m����иmlLR¡�|ꔖn���E���p�û�ѸV�ȲEo�o������N�c���uU����{��ko��\�"�����R%y@b�"��0DlGN����^P+��D��*,��=���-�h�Z�8Eg,�=�]WF�P�7.#K���ňx}����-<<.�%�r_�b�-]���8o��@֬�Ľ�L@�e���	W���`C��l:�;iky�7&�z��'s�x��tE@���'�^��uԸ�9�)���ЈvF��+Y\�ꚭ'tC��9Q��d��P_�V�h��t��g�H��7+:�E�V!.����{��<7�N݌�.��n��?i��(�+]��@H�*�}�</������\3lIOoʱ��=�ۻw���٘u�_���gW/����=�q�3�|Ot����� n�栐G��^�43w��ݿ�Ϲ8�r��y�Vϗ��1}{��r��C�xQoX
������w�����/�Bf�%vC���=��+��v��Ů�@��q��Y�s�Sw �/�."@�t��!���H�Jԭ��Ԗv.2FRͱ�D"uW��F���o����Ę����n0���n6��syDr-�t��u\����I�Ksk*��yRB�e���*q�C �_Pܿஷ�U�+���ݎ�Bǔb��%=ѻ`ǁ�Otxd����ZqR��憟k��p5�*��΅����oW~�����gvw&�]S��"����B�%�Lt�24�}�j��n|{�r����}��z�ڥ>=V�^_X�c����EIF��"�!i1@��S���buѱ)T,����Qv/5��b�D�<�N�6븗���� �+H����iR�=gY��`Iн�7�	�ZV����Lc�c"�6�Fx�
�N��b,<v&��� �#^/��6Wz��y���|�/u�[4z�����;�hȽ�2kɺ�/<�8��P.# UJL׺Q>�"U��jUcǜ������s���*H�r���\y=�7�&��Mm�G<�G�c�yc�#���yN�'ګ�����v��~~�m���ZuU�Z'v��s�J��+w�����U���5`�����C��8Y��$d* ��"��i#t�h��빪�D��s�K�2{zs� xקv�
���ܥ���,p��{*�$+�*aa������:�v-ޮK7֠NH�u\�3���E�Ӄ_W��WSc��~2��
�m��2g��k���F�tU|�G
C���j <׀ӕ�WH�K���)�$9�����Ҍ�'!�N�K�]�U��Л�Rgz���̕�M�yv摨W9�Z�#V:�ʏ�i����{��pT���[�g ��h�p��d�_}�D};I�w<�L�hs2�N�/WYj��G
{k;��[�z'׫�ω��vh���7=0��v���?n�3b�@h�ٖ!X��C��_o�ߝ��S�mKu}�dMT��e�g�����tF}<�4��%�Қ^�Q�0M;�_tb�@#�W�O#���e��\��!�V)w����!�Y�S�hQ�-{�sm�2�*`���<>��pe���4��[�[�-ቊ�{"8�&�{A�?ePb�->$���P;���V�]�N$�۩���z�Msزn�a����O%���;a��8h*T�.J4#�����BS����VK�Kʸ�\�e<� ��Q>Q|���T6+)���cIxA�S=��S^���l�r/�����F��]P���j�j��:({�rt��� 6p9Y�n�"��QT��|j���=�ޙw	D��M�D@�z��`ҙ��E��ܛNG@q`9�d�Ʌ|��W���R��FbM�B0�a-^=0���_��=�}��G�t$i��d@�����u1:h��v\Xc{�+ g�w��F
���-Wz�r���9)�a���<er;BΜ-;�J�Q�����n�me�T\�ے�Vy!}��u�z�P�V鿢	_ז��rc������q���I)d���ԋEMKx��z�=ُ`՗��� >�w�/������ j�h]?�z�%��u�_c�ӥ��ĪW��
���;�K�f�#��83��"�I��`�eU�H���� Mj���^�K'�2B�'t���\-�a��E<N[�󝠝�N_=<-����*��x��^.��L?�ƅ?��l7ǖWf����N]n��]ſ.Χ����s@ȼ�L�͵n0A���>\{U�;��GQ�*��Vi�홽>�|Mt������w�YU��g�(�2�5a���,��1�mW���xI��546v��ׯ)�L���U��Pԟ\L��'�be�Ȓ�O�Q
�A��Ԧ\��ԼOBݯtr��v֯S�穭y;�8Ԭ6+·Y\#a�^�j�Ef�W
d���S��NF򁻨��Ћy��!��ut�r���:�k��m�2�}�0�|%4�K���]�ꓟ��^�72��I���J;5�ۿ=6��u��<k�$�>1Y-�DV���umvG�Tء��%�m��(�,ߨ�>��SÍIdm��a鷽Sj��t'W��7f����r��3�6�z�R��_�Ҵ&cͺq\��T�D��i��%b.�=Y�����jԺpgС\z�$��V��M2�]U(� Hb���2��jY�uGV��օ���DO6��r�x&��M�U�v�t����8a}22+h&�Φ��<����xx �Ju�Bع1w?zJ��#$t
69am\o�Չ�e��~*C�ǼҞ^9i�,���jsƺw���X<eGL�"T�TOQ�_
�<���kWG�&��r��^<S��q�ۦ*e>n�غ42ʄ�f)L�h*�!���O>��j���h��ѣ�Ŋzv�@��8/�]e-���˕)�r9>	V��i��Ȩ{M5T���V.�ɊA�zn������G	��}�K%�2�5�"%:B'p@��-�?D���~;����]4��t�(ڿn�P+ڞی��6=��B�ˈ��v�.D��{�xԊz{a��ҼaR/L~�����7�[ā�A)7' rN�ON����^��e��Q�e���of{�z��;ڍ%�#�8�.8Y�ٺq�]K���S/�����xCLN��ҡK2��Z�ԜD�U�=���/�@axx��k���c�V��I�d��R��jÍ%`�D�MV(z�A`F��d�U�i��(���c��I\
����ƹ��O���T,��M����&jT����Ay�P=�o��WK]ٓ���$��F���w�VG2�j�S\�l��o"��!��V�>#5��7YVb�Go��y+@cv���ފ'��P�U=��M���O����p��2�=}�M��`��$Ƕ�mɞYz0�͡9�x =�x�����c �}�[m�ӿE˦�g�W�M���{�֙P����_@��]a�멵�([^K�Ь��Τ�3�~�m�l|��D:���nUO?
�K�G�ڷ��йQq'�i��
�ɖ�?sָص��pT`l!J�r������_��l����g�+c�8W&;MNNҖй�f���$���mB���\V�1�dO��֜�RY|p�
7{��8ӻ���ȭ�Р�����'��:��d�Zڬg7^4���85-�:��^�渓�a���E�1�Y�}��(
�T�hl7h���E�]9�:pGj�ۓ5�IT�h���bW+�ý����&޻��K>���z BY���u�{,S�9T{�y"ԍ�bS�~�m?|hZ�	5j!�D�ȸdכu�;��%l∕rlWoj��c��-�ѿR�g�=��↴he�ɤ�t�f�
�]s|��Gm2=���o�;���k�a5@n�_*9�ÍW�q�Y������ڑ1�Y<ɣa�Q�z"hC��Y���*�i5�=�/{��*�IS ���qTsz�*&��SPI�Nd��+�"���\��7T�=6��֛�)z���I��:�b3������7=�}W�6���V�L�p�Ώw�!�]�Jr�Z{T�Ot����E������=��v����X�^G���L�#��aP0C��B�����qxB�yag'v�W#z3b]�2�Cs��d߰���[��������!u�$d* אW�;X���,��nי
cO�N�9�Z�Tl<T�ku�������U���iD�ٟ9a
�HzV�L0�W,�d��ު�(�N�J5Z U�B�K�F[�d!�j3N}^��u1|Q9�du�<a���[-{73���.U�һ�O;5*��H�"BxAvڒgU�{-@�W�ޫ�����q"G�ʾ��D�&&wx�PwN���:K�Apɡ�S/����C�/%r��*�s]��A]@�\jOC��H�p�;EL��uʠ��ϗF�pl��g=Y���Ǘm���ue�a{z��Qb[�[� ����\%�|n�m��S�L��zqot�ճ��D�Ua(T�1Ȅr�K��h��(F��(��g��wIH�6y��7
bD�
�\�6R�h�����ŇR�"��4FsvÑ�pו*Q(���BiԊ�1��Kز��rj�}\U0A��v�,uu��ح��]�O*G�f��[��.����u�)mm=�a�AT���c5d��ή�s^��۔�kv�L��Y���Lp�]k9
��������F��ceI���"�i�{f(3Us���JN#������������[Q[���=�'��������r�� �tq7�my�	�$y[������w�7Y��C�(�7��ߴ���}��X�רN�8\��9��6w�;*Q&u�/�W/I���]2(��&q���>&�#�v��f�:S7���S������ԗUޕ�v��Fk	����C�C
)V�P�a��W����Y���\�Ì9���X�e.�LT�����l��D�]�%�D����dT���R�~�3�&V�͖��o�!aNo�	*���	�S4ܸ�hs��V���^,�HWJ	��R�a�����uv�r.����n6.2�\_��p,bu��..���C
'������<V��t؜/��b��7�"�3�3~͵n2<&��yq����?=΅5�I�Kg]vm�U�zx��g�����.r�ʭ2O2Q�@�}A�	SI�L��v�ky�P�1�e&�'jg}{Ӝ}B�5c|L2��n�_kK�ؔ�1�W�pX�|#[�OQ>�9.�b�B���U�ű���(����ρ)a���AYc��B��W�d�6.g��Zkgv+�K�ֆ�����͙�R�ҫjv�zf��>E{|�!�rrݜv�Z��1�Y�9^&�(뿷��4
u�����uu)�ԓF���Q�(�]5GgX��jN}��ﭑ�XTGL鄥���ʋ�]fe�����[����0=�a՜�Ud[��}�I`��/E�vhDi�V�3Km,C�ؗZ攁��0.�7�A	^޲
���j�]�ۅ���w6�ɩ�5)n]FR��m�{�ݧ[���]���anPx�w�W!��onwlb�6�sg(܉�Pr�*7�w���u,����!v��3[Wuo�B���J�Ʋ���[z���a{SR�9l�`;Z���ޕ�����+Ub��n��{��2�����ݨ��;�l0{��NLy�d�2 Lwr��ʸ4nff�v��zֺ�ʦ|s�����a�.iŊECq�۲�)yd1�{��8�|�@'g
s�mQ��T�`�1�[� NW�6��s�4�6�^�+5h�4(Z�i�<����=�K=z���9I���L�y����f�b�!��w�֭�}J����gJ�J5�F���nf����w�»�kCS�σ ��F���TWuګeN�t�u?��tt�����:����a��c�p���.��RuJ���6{nM��o��eL.�fŗ"��V�n�1!�����]Hl��8�|�j�f�R���m�zP�,�2���y�*�[�K3z=��*�D��,Sy���wڷ�[ �O�*]M�ޤ)����2�zJT$��}{U�Uʁ*��qPnMpd5+n���h-榀aۈ^P˾�yN]\�AD+O��<u`�y��u�r�$ɚ�6+��D��x%|dC"G{�b�=�Ƌ
,����mrM�8�cJ�;:�ń����1eA�d���kF������
����`��+���]H�Q�/�|ڒ�}7�wo^.��vj�O�o8u�o-�-48̻�h6h�1�(�'O�e`8��z�Ӻ��(^]'x6[[�2�9+ہ�ƍ�k�ftM������#HDH�m#"FX�x9����G�T��0v��4��"�M�U��C�A�),[(U�BK���Z��t8�˗r�5���4y�n�K�e�-Wv_T��\gu��UF�;a�B����i9�ko���h[�p"�\j�i}:)��u�\�Z�$�صL1����wti}oz�#6iޙ���Q��]]�.�<��m�6z���Æ�K`�:����݃6�Q6�Pn����bf��w��b�K�(:
���+w���tR����y;\ܡ;/tj�'U͡�	�������p��(���]�{N�6�#Fnt�����:��F������p�����z�cAg4S����Y��˧G�K]nEC�Fr��K��ꪨx
����b����a���(�(J���.**���QU4QQI5T%Qm�����(*�AM5kV�%DDDPPUT�MLSTDE�:%AHRE4QQCSDRi4�T�DCQ�d-�RUD�U3D5KQTQ4�M1RW#QPIDE0E!͢&Z��5�&�i*"�t�*"��$����F��
�
h�"
)("((��*f��������(�

"
it訪��c4�A4UA�)J
-��UDl�:��c`�4F���*�b&�$��ґ�4�IAM,KZ�h�m�CDS�M�*
if#lIT�L튪�F�h""��Β�bJ��ѶJ��3G>���o�dR�@*����Mu��5R��}��R���cX�"���S���Z�7�7�{[2�66��w�:�`"�o�_}���v�r{��Xr�)SeI��s8��`�b�+u�\#a�*�^�gT"��ڶ����9�;�\����J�B�t�XnS=��]A�#WeJ7dD�&d�R����"�a�7��H�q�ְg����c����w���B���c����`�w�o� :�-�1�=Iec�9��'�������/��f���R���Y���-/zf1L���Nƙ�ޜG9���g��aLD.����ǯ��f����Q�#�!�:����P�v��+���n��;�ܞ�ԁ��ӭy�{��a]�¯�3F��.*����:Z(�.�:����:����ÚX鑐(&�N�uL�W��F�/��D$wژ�9׆X�����:������T�n9�'��m�(��,��OO�.|�:ҹ����-�MG��#fg�\_u��kouOa�t�-�!Gh�_j�D�
�@�T���v��-7|�y�w��%x�-̠ĥ]�l�W�a��Om��]\D(���{�U���~:|4i��i�i���:W���C��ڼ->��S��4�����{*��K���d@�f�w � %�;����X�<]7Zh UJ����.�Q;�1�����i�Z���^S�Αv�ט)ʆ#�l�!��k�D�"�l��a���f������7����+zfI����S9W*s��|Z:��CrrZN�ju���Q�⍸��'r�v�.s̓{�Ed:��J�xV���k�j?�_i:n�W3c:����xFy��
�
������a� ��hOS�Lo
6w�Q�����tj�����ܽ|ӏd�d�f{;ێ���p��;
z\�=�����s�F�Kk��vp�+�x:q;=չ�\`{7�N����;�P_i���FG����/���J��m=���S����J��\c{�ܦN^n�n�fn�K���@.�2>��$_��T�mĪЄU�~ʌ�Z�#��S�,����u���.M�@˯P���tbWa`������Xl6Aj\m�=1����x�n�=9d;��ii�I��Z����D8�"	�Z��9椲��
v2yJ�/Wu�,Z����o�\`�� !�x	:�����dͣ�IWǺwyh,h_��WN���༹j'���Ҭ��(9
J68��3|k���-�,ԭ��Y��	��U��H���yE��c4���+Y�5v�۶v+��Zc�Y;&�K뵴s;G"�d�2�x�O�|���c��隨Mh��J���u��[|�='=��Hz�����˔R�r�W,���$��@9�$�[W��M�O�ճ�UW� ��iONѲf��Ӎ���!�Tn �w~z�O,�@�o�`BU��靪Wy-i<�$|������w�T:�P1q�5j0�/̋�M�lC�Bt�����m	�*o�uo݅�&'��J���h���~qZѡ�9Pd�砷�#!�FDQ<3�I�t(�;�ݱIt6"��������u|���q��v���\o�����	�'�4{��1�1<�a�}��U�U��M��IX���kE?��魳�W�<%���^XR07�t�G�v����բ�Țܱl7{f��3���":b�.�2��+�i#��Uv�Y�M<�"U�FI��~n�`���"{]z:��E��^T��D�A�vBĄi�)��og�{.������rX�j"/\�
\�3��2,s��Ӄ_W�jf*�:Q;������D�}�n�؊ �^�	�.�|O;5*���Di}bBW���mI�EJ��=v��$]{���]��4�'bؙ�5�;C�R�Fx���X�P\2k��_m����8�nN���g�h��_c��6���m�Q�"�
l��֫?w$��eWt\�Ob��-h� ��-;\s��t0Jj�'-+T,뫘;+ �=;F�J��[��^vN��\����!�)c�Мv�y:��2�Ν�]�B��Won�\p��^  ;��M:���$e�6�ċٹ9-�M��%��4���=�	��/�����h[����:��j�a��&"��~Δ��n��+N; �L�����(&d��p�������B�@�a�;�G��:Q��B;M���3ꊁ�>��N��
��_��*Z	W/�����Lu�����4.�����j�# ��:��
&��u�`p��G(W�x�.�P�"3�!�0�k�tV'�%ˡ�O[���y��e{���\̓�Y��G��^x�� 0�h����{J�"}�Wt����˜��f����]FJ=7ߞml]��{>f:d��pj_���L�
Ҹ�n�Jgc��5���\t��\�kT�ؽ�ڵ{��+�)����xċ��C
)V�P�a�U���N;��٫�����o�u�Eⵜ7:��Q��v*H�ӳFӐ5�F�
/E{�'��nz�
�1)wkf����i��B�����?u���;!3
f�r�	�s��V���[,�B���E�=;���é�4u�٭<*�XiL־�"ݍT��{{QƂ���	�g&Lxv7��IXt��8��::�ma��a���Ա��0m�z���N��5\B�):b��շw1
������Z�sY����y�Nޓ�]�#^J�Ƨ�s�9�_UUUVv�:g��#����*s����ú�l\ed�����fVK�����Q]WSG'#�fR����N��v� �·�j�{R�e4n��=�)����"d�%��ӹ�Pqv�՝�b���c�~�T��-���A=f�����Xd�d�ܙ��%A�g�D�ΗOv�El�/��fF�jM�����n��W�=�Y_^g�~��6�=�k�;�n�7���s��*"`>�h�9�t�XO@ʹ�QN
��x9�+	�KԺԫ���+�[o:���4v��|U\,�k�DU��@�7)��u���"�]�(ز"��ds⢖L^m�ml���5��:��lQ��=�p;n�3ϢB���am׼~���Z;�|7nod��0�$�3�@�d*�)��_]�͊+Oùz�#�Y�Du��kC$�NU˛כ�{*���4M�HT�I@GB.+jC�U�n}0\�=ơW3��I��ӸTefk�u`[�W1��3�dJ�h�:י	w?��+�xU�����8r9�Z$�%yEf�{�<�N��!3Tzz����T5ض���<�æt�2x�I��Ʋ����a�R�
�5˜^<%�wx{]�2G/we����O6�$ԪwN^��I�ښRu��/s(YWsU8�1L���r��3�� Z�k���$�qoJG��t'l:�f%U>T���zfه��m�;ϣA��	��=+p��
G���[hp��Q�#ȞB~��Γ�J�r�}�4<mm<���.�T�(���.��"��](v�Y��z��sT�x̸�yFDHN��>��3�Tz�ǽ漻�Bm!�嵹&�k�C*�̸�����%�tn<P�|��0�5hݜ�9�-��Ȧ+��c�@�Տ���h=y�{�p�|�+�~��I�;�#�R��c�^]�u�2>^�6~�瘯�:��m.�>[U����|�^�y�:��i�ow�;9A&��rX3�k�^re�	2�y�(��;�`�U
�]c��o����!�ԡ��/K���f޽�ʳ�9Fes��^��j�nS�ID���6^$_4��M��o�J���ga���Q/� ,�xӽ8�#�B���U����z�Ҋ��nz�}){}����C<�1�J� ��Z�ڶeZ�;��QUs�g�]xQ{gh3Y}&�,հ���d�r8q`�}.W��.E�%�Y���tL��X=�÷����R��ͻΑI� 䝡x�;(.sWE��ˮ�1T�Mc����_9ղ�8ʼs���I�QnM��}_W����R����.�?A�U}%mNt�%J���cZ[���FF��5:�ܸ��mΡALj|���J��TOv���y��	��x�P�|3܅���>�o9gx�TTt��I@�s#R\�3V��m��x���*�زd�ӝ�޵٬gS�r��^P����@ilm��W��7i]ms�y�yX����rҸy�p�b��v��g��H�n�@�z�=Ҁ�[ӡ!z�W��o�\毟m%�)&���w�m�6�S�fF���9=Y8m���LG1���K">��'G���ִr�.e7��,c��71Kr�Sk��^��<���'o�k7��9J�_�uO����[1G��p���ќٙ]��j���P���'��k�[�b�A߯�C�ci��P�r�������4-�^�V�7C\tŮ�}/3sΊ��-��œ�ҝCxdt���=��:eүZ��.�nNa
PEzid�@�Fe�%&�X��J�)��hY]�E"f��ͺ�[�R�4�]G��d�E�m�%�,�8i%;���s>���RXiɝ�������Yo{ �"rfP��o'T�,�Ǽ���ŵiU��'�����m�j^�c-{sW����A�֖��Y����g�{�G�y��լ	X�<���+}��8�t���ͥ�o&߱d��V{�ON��O�1X��[�>�L�at�]�WzU��Ky��(R=���o!ɓ-�*�(����R玠�iaTcq^��'O=���H��/y�y��o�gD�r�/l�
q'���_B�N�g\tZ͹W�ZM�ā��h�<C�-�����Hș�m�W���	=a�Z}�^ȼ�%�����b\J�4�Y-�ke%�.��7P�=T�a�E���U�7P�9����-頥<����c:��9AJBa�P���:�w����[<�Ί��K1�O�/��c���b��w�Ȝ��ɣ���Ԓ��bh��~�0��Rؠ4�y��.7��V;��֑㉜�dL�hnvr�䔒�ή��_VZ�o[��ڪ�������-��W��H�.��Bq�ƶ�;�%���W�=�t�W7��۰vϛ#��V+5���O Õ9f�SP᧸�v�iM7����[���c����[��/��c��:=GyE�,���������su��Ѭ����v���%!�	��[����c㗮iw*,�ԪU��FJ��p���8�&#������ڶo��V�id9�+�T��񾷞�����[���T�4�kɱ���	�f9F�X�)h�9�E�b���Am���ڽ׵��ZN��i�i�#hsʭxbC�˩�^��A6��?k�����D�����;���c�5/���q��T����̇���q�O#/�'���[T#1P�|VE��N��s�2�-�\��1uYv���&���1���:f�����#F�	��C�"�{��y���U����i���~�"�׽��sV��z��r��K��IA����e�B���O��ة#��ފm7%���ʹ�gY�㺁V#T�g��MR��P�TU�ץR�S���\�}f�{l�R����Ȗ��
>"^��ќnmʈk-ۦ�mJQJCh'�lv7�/t=�Rkjp��j-��׳�P9�h��7�+`\2�~�����S�a:��JK[V0Q�r#�ä닠Ѷ"�H��0�M����+B�c[��IS}�+�S��l�z����6��<�z�W�W�k�{���aO�ԝӳ��������{k����%�7��N���z��l������:������u)i�RymC[oam�JZR��ᩬ���)Ψ�r=�}�8�ԕ�����Ɯ�蝥%T��.�n����[�x��q�p#�݅�%�cJk0B�R_y*�ø��]]V����ⷕýK̆��r̄aq��6	���&c7�	�ʷ��3P��Z���>7�.j�/��8�[8'ʑ�GDs�R=^�x�o���	^���B��w<ڬ�[[ͧ�}'y��c��	N�+	Z�y�j	����G]����Ȩ��\�{V������Za��f�͈�U=�9|ڄbqm�a8��[ڴf�y-�\�$����CQ^�^���}1�FU�/Uq��W<7�8S������:o�>�[�Q�F�mf�S�N��mW J݅��%���6�@�����vi�ė�>�]��\��3��M9t6�`u����t�/�i�[k�PC��ʺ�a�/$�*�gB���c*7y��\*S��Y�2��kV�he1Gzvb��F�\�w�M�>#2�CW���5BX�����eYYvױ2bΩ�fŢ��}	T����|��^n�I�t�A��%Iqe���R͎�l��W>�6 ��Kj�v��;S2�2�7%oZ�a�/%��RF�&��t�z:JT-N��X�Kl��M`��%��)���Sn�V�j^�Út)�9����k��XT�
�s{R��4G �R}f��X�nuA����Kz��}�J�a��t�{�cgޔ��镣WA�#�]"f�w��fb4!��U�����v��"ѭ4G^���x�Ejc���r$-�\5����-����
ix�p{�q��F�%����UAWE��V���qʛ�#q��d��J���r�A�g`*@l�؎��!렯�lN���y��f�<� 1i�4�-͝u�} RnT������:6z˵����wj���5�.*f��-V_]��#�#:֠�agVut��h�}��vld�Ř��.gj��S��ٻ�8��6�\��* ���-JӮ8���f�leI�xh��o`�L��>�"F�$�k��B70�ށ��T9~�@�^��Ze�F�l-���s�#y����n9J��v�uՌ���Z���K�i������М�{�V�C$��Fl�{��\tq>��R���8'!�w��#:����jd�x��4��6.Q�:3{ڮJ��
g�RK�n����_����E�������{�V�9�})}�n����psו{�]Ϡ�C��mf������0:��[KJq
6����|�;��S���+�՚�]Y«kX���KL��Գ������'\��/�fG����h�8�[��,���*ݒf�+fܧAL��e�N
2Ό�fF�[�Ɨ�VÜoԵ�rClзS��TH��Y�Э����QUbͻ��x�I����� ;�\������Or���wW^��{���y԰��!)�_�'jf���X�KnlVq�2�$��[Vm���jX��馪�'7댪���IO�"��m���x�9W��]��H��:%N�c)�':�b�a�2��z��fWe�1�T��%gJ��٦�!�h�$pJ߄Kq�ns=(,�n������X�͛XU�{�Y��=΁� Q�.�HH�-;t�$�ĺ� 9M7�\2�S����L���U�� �e��V���R ��՗�3��P��C�Uu�Ծ�0���9\zA��B�3�}Z����q� u�lP�-�^�4�kҹۄ";��׷w�p�uS�i}�=i�ud�N*yD 'm(2T���my�j�A�(�*��(�d��3x;}�z
�y�7���� @QLQm��A��"�"64�DT6Í�DMU�%kE$UE��ADAD�E,S)TU6H��#mQEI�N'�I4�EI�i�j�*j�%����������JӨ��*��Jh ��+Y��[�!��Q4QMREE%4�AU$�E��IID�U���1A4MUAPDTUN٤����*��&��f�)j*64I%AA%QL@DSICh1SZ4T�QT�SRS4CAKP1%UIAM�T�̔���T�KCV��P�	CQIAN��QEACT5�-f���Q@�E)UH�QP\�4UU4�ST�UIA2�0AMQPP�ˣl�*> P�U�W��s'vh�DY1|^���q�W�Z�Χ�hn���iu���u�μ�q��Pfhӵ���s�r�}�,��=�����o�.�����{�L�6Ƶ��:�<�Uf�j��)�œs��Ԩ��bƖ;Nj�'�� ��i�R�����7Y�5�VU��r��*�"�L�xy�۩Y��~�:a��0�|�=)7�m�����;���1j݉	m�����"�%���U*z��	^�hcq�ƛ�����}q��o���}��Hi�]�u}ZIJA�!o�:W��^��j�Li�o`Z,��&��{;n�č�@d����vGw��G*s��%���7n3P�12e4���{i{{,�u
1�-��`n�P3��!��{=[����*F*���f��ı��/U�m�Ba_{�HwS�#-�v�T�ێ���r�(�އw�!�b}���<չ�7{U���<�q�SUI���cn&J}��8>7�ki�܅���V!-
�B�Y��$����홡YWu`���r�)�z(�C�$ЭD�-�35M�U�*F^d�AU]L��}�(�2�Kݼ-�k��W��"{�������pάy�M�M������>I���u5v���]+q��H�P:�:u�]�{j���'�^�[��Ǉ�����m]V`�?2ˡ��>/\О]�~�N���˙M�;݉��y��\�ow��:r�
�8��\L��4Bwp����c��yye�����~RG��@I�[��RQ��ߕ��xl�젭TN��8��M�����c�ݷ9�I�x�6�M�^&�m���s^��k�bZ�I����U2���w�}�
���y�ˌĪ��R��1�`�QՏ*�Y�����$�F��W_-}{�j?h"�=~jv4z�ʾBEcNʗ��z���y�̓s:�;�]�d�)�Fes��	�ʒ�vB�䢼y��%�坑�9�p&�1����Iʩ;oڵgY���V#z��W�Pj���Cэ�����p�vdw=�n���3�2�!g]�B{*�>�T"{n���Tj�{i���=�7��]oͧ��i���ϻl�z�F�(��ݡ Ӈ�"0�
��Y�����P�._������M| x��h���&�ܷ���;�v0���:n^�<Mc�]O:d�塻+V��c�7ljxR��̢����(j��1;6��Z�-�a-��	2��9��"�����K؆�X2��Toޔ��Ԗ(к׆�B\�����P���2t�ؼ5	���U�-��U����1�ޚ
S�kZ�b��q�
R�Rx�km&hgo*��Sp�����cc���W�'ŗ�����8��:���|����Vm�8dq���S	Kb��xw\r�4���fi���l�q�Y��v%��G�B{�`?[5�����x���-��ٗ�樛k7��C����!R��GhA�:��v���}s!�Y�ݛ��yT����7�44�Sc#�uى�f-oMZ�`t<�����u5���׭��Cvnl���S�lFs�C^p����Z{m"V*1o�i�fuJ̡<��絹X�5/�����j�[~��ҭ���1��}�E�Q��f-���"�W�����	ۋ:����m��+��9Xt�-m���X��(�q�;
����9e%&�LT,^Y�S"ƥ�:���Z'���R�l���lߺ��:�\/I	��Wz]�L	lR��kiC��voS�or�8>��7�7�.�wZ�b�{��+�d�+f�ﾯ��r�u���a��������x��-��_�,8����}EԂߦ�7�EX.�ZY�����Ҍ�����sV�����uaͬ�(�ަ� &�VV����'���Q��4�����tO��(����}��N��W��ZI��V�f�97�'�j��V#�a�=��5Y��j�y���]k���Һ��4�R
���=�]��R�����,�6��Y��}�Fm'ݜ���'�
��I���"'��W����ή�=z��d��gm��>�[��S}��
�N���α)�f���&�F�0�LI�q������Q��)���.�[	�ƙ읻Ӧ+e�*�;��ѣ2����M+%ޥ��Ƞ�;A�2�=0�{p`�=�w�i��X�f��Y�O�%�Xe�;�a��H��������n)�k<��%��)�6<��r�5���f�W���'y����"aǈZ���dG�S\�9.*�i��k�_N�����f�+�'D�r�]���uiQ�u���+��'�Q�],U�Su+�,l�0�lu�9�.�2)O7�����ΞP��nv�vnG�7�|��o�hsN��1��wں��.���n�Y0���ۅr{�s���3���+K�j�G�v�셈/b��b�j�_08�RxbZ�Z2� ��S�\Rs�kT��i�w�3T�M��� ��5n���{T9��1o�Fb�6��`�_��1�bӶ�޼{@��fq�w�R�mͥ��Wi_Z[C�1�r�v*���r�M�Ҧ�L�~��2�!5�;Jn0	x�۬�y�U��s��F�24��ʎ{m����s�$��!�I�RnozWf���\�7�6�9��~ލ�ڴZcxk��s�^Z�g��L�b1�ƛ�M>�e�m�OU�Y���Un�7��rz#4�A�BK��B�����]Ixp�.�+`�UL4�\��+{b��Dn P"*���ɗ�:��+go.%��d�ȜNS��lG��rI���I��k���Ղí�{t�<��
B�����t��B������O�JK��L��Ť]�rA�Mފ��/L�١�Z��mV���X����I�z�L�yُ�M˝9�ͅ����0��JP�Z���{��Rp�xœ���m�5����K�Tt�>���>�<�Q�KԾ��C�7�ogg1z�{Z�S�A�촵��/x<g)�ue�I��c�������[O���kN�ub}��-+�<չ��b���f-O�rk�3�N6��1�ޑY9=�Ѿ��i�w.�KBB�N�W�������G�{w-�j}C`��hO.ڽ��Z9C�3�ݕvk}���[�q�q���	R&y[������o�g��ˮc��������\���e_(���������t=<v�(<n����6�v�5�}T�7��U��:���5m��o*��:�s,���6xb���d���ߗ���S���N�kE�LkX5�u{7�~6��)��o{��DL��]�{^��2�i�*^#��k��_L�+�@x�8������,b��^�y=�����E���U��ϼ�� ��[
�&|�C�`k���K������h�˰9��|+%��Ӫ�2Ƥ:[�\��Q���7q�y�j��۔q��	ݢ����ϩn�$n�7��f�����R+�,�f������<��-7�+�8c�p�tv*�t���xl�=H_%4�:]	eC�4�a��;�H��y�o}qm9��6��7W��ǫ�UqŘ�vb��]�s��F_��%�M>�/�l<��휪Q rU%��"�75%��u4믖q��'O8��l5��}bZ}`�����
av�;w87��)8����wJ�Д��o;ϡ�����i�j����K��{3���/Y�����P1�'
M`�KziJya�k�XΠ�U�{�$�(��0Z�ƒG.�!'/��(Kb��Y�G{��_u�X�U�t��}Te�W�9VyP�Vn��R��;�t!G�F��2���T1ٓ7���Dș�����&y�^���Co�z#���Ѡ�G���-��8�1Z$�����y�=�����7�Q��p��D������½���p34-��V1)���Ռ�ar�r�+)o��Q��=~��'f����)�C���o'31�q�l:�ST.�U����w)�1�Ø�P^�Ąq�}���oZc;s�wQ`,t���D��nh�e�g��0�s�uK�������l-���_v��jZ����Ӊ���a�ŎQ�;�S[DJ�ո��m�ۮ�	?b�z�)T�W�ni����9�J9T�&��9����X�Z�;�U���(<��'?ERy�5�����Vх5N^ul@�pv�v�B*y2�:�����E�?����$��UL}ᇧ��k�ꅠ�M�y��g}����T7�SƱ��\?q�dk
���g��̮չ����J���~s�{�3�j�����9a̧��Hv���eݢ��&W1&����P�n(�qbZ}r�6�z�gaڧ÷���ū��j�onL�����H�d9�mC�Y~m>�|�+h*�n J�ÙU�����@��_�t�륏ǧϹ���[�k-�-�S=)qQ9����ܬ�lޡ0�GH>F�t%-5�΂Ÿ���2�Ȍ�[�ś����nZ�7�����Y\m��(����\�!Z��T�ݓ�G����r4a/|������c�>�؆T_{�Xν"t��3����EwU�-J�3�j�$�&x���&��.f�eso/qu�xQ���zs�@�y6O)q~���&z����u�'Օ�E��T�%mt�H�ު�T�"gV&N�P��B��r�����t�����W��V���b�`X�.�������;NY��)�L$#��zc&*�s1��8�^D_\���6���K����n-��3�y��7�૔�+~��y�3dkм��=�k�k��y:|��}S\ӆ�b���=;ũ;�|ܭ��d_;uq:���2�9�j�����mTȘ9Ad�3��-��eP��p�l�P��8�[Q������̖ܵ%�ȁ�m���kx�+V��~�L���s�z�-���OXb5�>��~㞾k�����߱�{I�*^X1�f���c͠��׆�o<g�,]W_՘�ڒ=ߧ�lJ��$�c9	�i�R����7Y�5������𬘥$��屭֡sݢol�n&�=\)8��҆��w��}����4T����2�n;�*�tݝYd�6̻��$hЖr93��I��(ʔ�Y��ۧE-���7�:wQ�i��L�˙CA�xS�}�9��ӻ����Omӏ�쓪�\���cS�����X�$�I�^��)���f�E�#w�[�C�d��T)Gu�`�.z�'PJ��Z��P�z�s.��'e����1q9�ҹu����m���9yP_W�P��J6[����Ue��R�5&u�	e��}r�����_(����II����`���=��n��Q._Q�4޾��=���ߍ�B*:{Ϥ-��U|{*+o���v���E���-�w�o�/��Z�`�u��)o�����`��bNP�)�܆�����8�/:69+�[؟c/���[���<gj�vv����j��=��%Y*�I|b�{zDl�f���U\q&���;�n�(�^˼��)�Y���FB,�*6!k�˲����s5���*�t��DI����V�����*D��:�%nMM��`F�\�3e����j�ݖKW�Қ�1Z;�R���/f��k����]	��I%a̛��K�t�N͍���]�i�ضq���0�w�O#A�lﳵh]]C;��j�v7c��B��Y��Եv��&0��h�40.��c���[�o,Ӈ`�q�
��Ɓ[��7a�3��� V�ծ�w����Vw�TI����8+_L/�����+3�]řf�U�-�K�۝xqa�Z7�44w3iɻR�	��kJ���4�5�wW��r�5(r��:�۝�� ��t�T�y$��s��2��b���O�n���V�Һ�"�e��Y�S�v����oMz����%K�f0��*,y�w���Q��L�_%�$�`�QBtײ�Z����Px�{gP���B��e#�V�t���o�Cc�����_c��|;@�Tf�&ǘ3-��k��=�̉�/o��}��jVz��.1�tu�F6�t�rT���#��`<bp�֞q�s��t#��UK�v:qG5ٽ�N������\�%�S4eN
WC�'u3�|��n�GWua6M3L�ŋ�V�J�"*�Ґp����ᠾ���-e�a���	q�w0�6�ΊNb.�Z�ϗg�}k����]'�ɥ[(�_���X?��]F��+�5�/�����J������*�< ��J�R6�8��l�.yu����U�LV�g7�ʹlш3{��V���wgnSUy���Au'�sR�:����q�Ue�`P:�"�r.�4瓧L��g^j�P�i��[�t�{vm:�����vs�zD����a�C�ey���6��GI9[�����������c�s��V|�m�o��qk��s�Lɣ �5��f��ݒ�c���(m=೔�n˝��5���Ø3nCۖ��&�b-��{%T{�.�	Y���7.s�6�^���%�n}7%-AH�t]� ܣ)4�i����E�r������8�"��mU��i�����ɵu��{CT��r���r	:p5NO�m�Xްl��+t�:o^t��t�K��t�p�n9vf�K�Y�PT�_nK�]����;�j�bty�e_U�xRW1����n�đ�C�luI��,Ӌ����#A���V���G�C�En`ý]q��V�����ش
|��t h�����q�}�$O�[�o��
#�Ճegx��	 ��U�l��|4��=�9t暢[CcC%S{�r��"�9�:��$<���>C���ն쑏����Mr�fwZ-Δ��;�d�:��#��CF���<��@��F���7+��5\ yX�q�7�N�&r��b�!ɽ״��.H��ϛ]=�2�x�r�Ј[C�J�[�v�c�u�<큍���~3��m"����ur��)�X� ��QrY�D��J��t�,d7�7gNƄ���,I�/�AZ�����|F*"�d��5�b*b
�lƐ�AA�()b
JJJi��mPEE4��������*��UT�!H�RLJ�PQC�4RP��Ĵ5U��R4�+UR��[`���h֒����#�Il袒�i
i��'!tEO!4� rLW,U<�h*��LHP�CCM�PPi�i��'�JRDr��R���h4�J@�C�����"
�4�LA�"����J�@h)�-�ru�CAQ�4�;��q�n��nhjaW��k���Tޫ]Gif�9�+]�c]�p8:u���=] �Dp�`��������x��m��]H䮝�&n~{z�کX�O6ƻ�3�5�Qh�nad�f�e�S��j�n� ��X�ܪ�����']c�B3[ʠ5��=�w=�D��v��'wX�ׄ�a籛�����y��k��Ǖ�z^���z��N��B'�(̆��ٷ�%de�9	�;*^#��kNj�/OEF��!5�F���OZZ8�_�maŸ;�!Քgu�B�%���GI�&,F��E!�v��ެ�;T㲀*�AޯK��N��tl]a�/�5&�,�ո*RN�N�9�=5�3��[����=�u����+-5���-BeS��՜�\kqB�kOP��X7��g��F�����f�q<���y��t$�T%*5�M��j�{i��͵�v����شj3����y��[�'���#Ie*�Rޚ��kV���5w~�;=s7����}�U����������m���l0���qìv�Yf���I4��[��=3szM���?�K�Y[!��Kg�۞)�Ƴ�{��󚃫����8���wJ�Y��5˼vd��̋�:72�Ӯo�e�ޜ.��훿n��T�Ňu)S�V��݊V\�]��-���k1���ӗ�ө��Z�;h�Æ���(��}�_s�Lt�W�#3+r��U�{��;JUD�v��u����z)�3��.,��
}*��"!a����3P'���t1��k���CqN#�B�(�A���QR����d�}���H�w<߰�{cy����T�4�Sc�k�P&º�aQ�)zx+�U�uM4$H/yl�uM������؍2�N13�L��p�U|(��ķ1ohFgT�ʞZ���ܬw�������Q��4�*�c]��o*����b��Σ1}�H�iN�P�T(�1Kd'϶c�g�|�w��Z�T�����׵�z�����7>b2�ܫ���M�����X�zBk�*Sq���k7�=�*�P��U�lv-��|���E^\�x3���qXk��֝�6 �����ݲ<ǥ紲��b��7#�������y�0��sy�5K޴u�ܓ�3���mʃI*�t�,���������]��)d�2���;���Xr��ܒ&rY����Ճo�Dy.;���Ш׾^X�a��C�F'M��O�Wfߓ�Y�v+0�R4�I=}ǅ���Y�NXspt�ƂV4�W�W����i����Zg��p�he���经��������1��I��e_�*V���{b�Sx�Fv��]��F@�Q{���bF�jd��K�����h+�F<W[�rd̙�9m����r���*:Gy�W�qb5%z��g���vF޻��ʑ���%�4���7���9F|�)�{�Aq-]�VC�f�%9v�V�Cej��v�i!�,�Ƞ�;NY�aQ�CV'�Ky7����n�Tmz�`'�^O��&����\�e�;�8�[9�鱎7hp�1uYϒ���zB7���/\���y:�:�}SC�p�D)���'��V�M�\�[WO=��w�|1A[^�p�/'9�n��뚜�-��Q�;����<�K�O�C��琯4����x�}��Lk���K�뢥��N̋��E����
 �ee'[^��*��yڕ�)�
{@h�wm�!����e|�!kc6�Hc��$=:n��(*ή��бw6=�J�nr۲m��	���;�k��A&��k��5�3�E�����уȪ���}��+��Z]�,ζ Լu�i����4-�;a���f:�T'���"����z���9'Nj&�9Ocou��O�����k���w����)R$��Vl���_�Z��M�����q�3��V4��)x���f޽�H�<���j�OE�<v#��}�V��WS�Z�j�Y���J��%!rN9�kPݘ�IywG|���Q���cw �Ϡ�%�A.��hcqY\�$�s����տz!c	>��zz\z�뷔'�9X���P����]����6_!t{X��,ce�o�Ob�z*:G(��
{z`r�:.X��]��QY���s�n�I����Z�p6�EGw�F�v������ꇅ�ʵؖ�ӗ�~KZ�b���)c�1��*�B�IԻJ��4ZwOE7�b��k\���.i�R��Ӊ�y���)����:�n�4���/�f�0\Yh��{�`���y��u`�W�]��� QX�-W5&n�,8�K,u#b�C{o3�'���갍qx��v
������Q9�]g�uu�A�c�q��ݷ������X)�C{ը;{�-+�V�{��y���C���7:�����ۋ�l)fB0�w���'����g,\r�iJ�����s;cfm(�̍ȭ�z3�E��+�݁�ٵ����x�����������'��}y���L2�;G�Q<�j��پk߽���^$�D[��
����K���j����h��a����u̳΁���<�"��s|��K�OnT�j�՝��XI�X��6Ќ��k�lNY�}sn�bV���ű�z3:�+2��[cu:��w����k��kr�:��R�,�X7�lI܊7�F�Q�^)Ȍ�m�+#,g!5�;*^E��o�]Ae����O���k�������ZA�֖�5��A_`�\(uH*�چ��.�3�#��w���x��s��O�A�8�7=�Ut��Ώo��9���V��uy�)��mS���㺛��f�ᅞ�6�Wu5i���a���3��^!�iMfc�R���X�7D'���d���H��L��*�D��:�f�S4�{��\���U�n�A�J�4��LG��j�7��qtQ�)�ATcqC�or�}��z�T�m����n9���[�'��M��H��1ZuO�`F�l4�����z�yQ�;i����R@�u{Ƕy��(�?]Q%mNPڝ�5����ǰ���{)�"s���.Ju�x��~#��S�I����讠�%,5��}��/G��"Ni��t)|�9JR�{'����W��1>$��yO^b�[�����i8�K��j�2#��i��܌�J��fqb�z�wzwa+F�˷�A����,�Ƞ{Nٟ#
GJCc�>H��n�@U����F���v����:M�;�f�+��K�Rp;����h�7���Q��;�{�Лܜ�]�� �T�ӊM�w�pZv��۬��o��b�E�ܡȍ��K�˜絻{��ZN��Cs�b|)Vֶ�[��%r�B0�(���e`p��{��6M������mF���:�|�,7 0�8���n�V*��<����c�e�������T}�EW<�s�5�Sxb�\w*m�R�<��W�n� m���:iH����g+v�d�}��]I�r�ܲ�<1<�E���wu:����������<n�{��O��A6�$�_��讲��b�M�T.���w�^2h�vdfՕ�՛��lD԰����^Xi�Y���?�h;F�ܕ����.����k�ڪt����Iy-!#��~*Sv<|缞�'�HO����٘���=9.Fo�Dc�'������Xbq�&��=ރ�O�΋>OM�.�Z�)����4�W	�W0vAo�u�lZQ@Z]��|Ƀ!����Ӹ�W��V�6�e��!K@�Tw��sZ>ֳï�wio��V����`�oLL]����\�m�͡Cf7�0:@Y�'u]mC=j���k�ݦ'��a��{/��kl=��睔�QQ���
�8�Q�5�;{��٬�O�kO�y��号q�@<g(9RB��t,�p1n�3�TV��7ж�Ď��"jee��@v�'ӇG.SG9{u���@��!5-s��K�إF�R�+*ί^�{����7����F�]k�4�8�']�Ӥ�R�e
��ݒ���)�<J�L�Bwl4b[�C�Q�����r���r����U��S�=Ln�/����������%{�΂��Wqٹ˳�M+�z�7�<�;A����yu�	/�KR9�e!�=)̹w糲�Ω֛��Ն_C��8��#�w�=;��'��U�d#�D7���<�+@�N�(����u�$P�k�,�2�+.�v4_6pHUw�'�yס��sZ��T�?EJܷsW�x)�^ޙ4V���j�F�c]��k����*���{�N��8���_?b�Mm8�kՊ��s�10�[q�ʭxn��ۺK�'�r�޽ר��?J̯J{cu:��MK�i�k\��ǒ��F��_k�A���X�=�{��=I�[X'Z+��V4�j-�|���E��Ԭ�\�{�*�+S>�p���b��֢�����:���߄��zD���8��z&��l�iz���w��y��j�5�Ǹ�{��)���^��a�O�:7�h�(;|b�{�wy���j��Q����SC-׮�r�C�ǲ@:N�=\�'�眜z��­�xn����$�n��B�S������D9T�'Vk�-�kof]�w`��9���i��Ʒ�w3k'Y����v��r�ї�4�4�ľ�w�;l�
Q><�
�^���E#�������q��%}��[��]i%�ob�y�6���Т�/�V�uf�\&���ډ�_N���B�^�����*8��S5nY�j�2E�#O�����oJ)ބ���c:�E��� �E�_]�Ȫ�Q�Q����	lV�k0#�X�P�녍nX�9n�}��C�c^�Ѫ�'��\�I�_]�2�r��t5�B���7yY��;��]fy��Jٷ��TFߠ�W� �nO.��jq(�3���_rP�[;/���M�;�v�*/�h�B2��$�aD;SuZ�6r��augK�ݵz���龩��8�m�v�N�1�4!;pVE�պ2Χm-�QgwX�rݛ֫����Nz��hu�[G�7�5<��D���[�:ӳHP�Uɭ�]ImհO�ۭ���Fy_/H��z.<�=����K����4:ug(�����'Yj���nv�b�(/GT�\%��e#���ɷ۷ǥ!W���C������8s�(��nm���ӌ�s�2�G~ʽ�m)��HE���o�^�j^���Y��s���|����[�˗��}���:Gl\��'~�e�P��V�ic�/��(,��.��[���U����v��UCܨ�;����V���QG3_<7�I!��M�{��򒑵����a��R����Z��12��v^8cqϚ+���W)�Y+Ͻ�Z}{�P���\�N���Aw^���Xt1:C�a���_���Yyu]�֌����3���6�(�'��΄����T�ya�5�������^�;�:��ϱ�U�P=�DÑ�#c�� �i)S������ol���u�8b�y$���]<��R����Dw8�4�V�%HR�|�^=�0�t�2_Nr�kw�3�������vB��;��;N7��Z���v�^{�T�jӖ:�&��fE�{�SN��U����	�1 �$��x0`�Y[4��6qe�яM�gѫ_݁>���}D*�
[���U%�0m�4EZ��jޭ���+��9U��5��W��{�6��i{%��ڮV�h1PA�o�H�imK$���P�t��N��'n�%����9�ێ�y�κx��l�&X��W���Zo)��+kΧ��nP�e<to��)��.�7QN{d�\]��{i���YZY3�Q5��J��B�����̴�d���^"1}a՜�
�y�ݛͮ��i�\�7��\�ʆ���(d糑;7o<O������d�9+p��Ʈvr�͵�EL:�C&����P%��r��9�a枟b���z���oZ���\4o�f�dF�����u�l4��WJ�<4��Nn�ka����ˣ �0�S�8�at�Tͤ���;�(fC�!���y�/�=]��0+�[\7p�3Sp�Ք��5�X�z��աU��C��ӎ��YtGvp��z�U�R�����ʹuT-u8U��Z�pY`�7E�����5��G�ɨdA���<h�yB ǯ�$ȻB�f,oS�[���VP��դJ�>c��l��4%<�C��=Y��ً��̋��Al�@&�}ݮWu{}Cn�X��5zN�сZ����.�Pp�N��WYb�J;�d�N�����w�D��mұ�7o@�r�K�-��wf��/n=�[�|��.����K���3�cO>��3�'�\4	x#:u^�[R��OE���^�k�Ϋz��¶#JTf�is�G8f�Wd�}]�q@z�F)|�>4�n�8��VN}�[�䎎���k�ĭb}��v��[�Է����"��NfgV8j8Vօ�\��V�h>ӷ)KÑ}�%�]��]R� �pZu�mky�A�۲[��BH��t>T:��D�F��ŕz��[��'�����"�^R����Ys��tp<v�kz�#5ɻ��9j#�jY%Z�[񣙧IL.|x&pz�)ݦ��u�\��t��+s�w-	P�&�6�wI�.��m�b�����vT�����oc|��[����^U�P���݃�P���Xm�,N��՘��5�eik+�k��\���\W��5��@�'n�)�E!ꗽ��S�M�x�TƎ�:� ��/�#�����2�+�٩����K`�jcD��^�l�u�:���m����j^`��L���+n�I��.3OMr�𹓊�Q���V��$J`v�ׂ���[�Q�_����KT��P�R�YՏkK:k)�V��U�.YF�[P�o�wz�P5��-�P�6�k9�=�]"��˓9���N\���n��*�T˷F��M]rנ>�L�Z��'��զ{���������./yo`OѤ*.�$p��"�T�Z�.�➺��^La��ٗCZ�;2��q�����?�_��ς�U7�IԺR������"(hB��#�4��֔������;�@�l�4�EQZtr\��S̀����t�����KUTahJ�%1U	l����s���������+N� rl�)���jF�F���@r^A�еH�Q�tV��1R�劦�i�C����M#�HP�Q&�\��1��*�����(h�&)�*�170Dr)y5˖����s&�W�i���F����G "5�
I�5���`*��ŝ:+Ins쿪�u��}1�-�EM���fөu���YŨ�;(D�G��\'A�N�]H�m$Omf������<X�5��E�&z'�U���� ��~��.�M$;Ա�Ƞ���g���n�0�t�����+[����~F}�Nj��C�5Γ}�6�8��T�� [�H���w�5��@汰nr�S-;�k�6�gW(a61�{������w�f-@v{b�e�?v���Y�^����Nf��t3��\�,����1���QeglbW8���6`_ehWW9��T�����}�F��ʄF���7��6�n��ډ���|�Fb��ꆶW$�-R�{��|�ׯi;
e�Z�بm'�W��6.�=�;D\z��&�ٺ��.T�In/��|�*Sq�<�=��z���F�T���2i�a�)Q���Υ�a������!��CU��x�l)����Ck[��V���۲��n׋���[�%��<-(}�=�s{TMi����qVSל��s<"�6h5�j�D��P^xZyb��A�ʏ"��C�Wr�|Jö�Nٌ�2��CSflQ'�7)�y/8��n�:|o����{;8Y�����S`��Vf��i�B�:=Qٮ�t�cUHʙW�^�KSOg7H��]�:tV��2�29��_P�p�J��9;5e�X���I�at%��m6�Y�6��N�}��8$��R޴ ���^�S�d�I�o-�kl=��睔�^����}>(,Q6�9�#^�4��5�<ΰ��������>��m<gXB�������܍b���["^tW���ٵ��a4�;�a�Ȧ��31j	���܍��mU��_����#`�y��K��%6��w6������f�����Y�t�[�tk�H��Pp{b{~�*���ӝ����Zo���ؖ�-���L���h���q�� �@�b�+r/�ԻYKF؅=ԥ��bf��o_�j��4i�5�3>�f$h�[�!�q1.[<杣w��v�
����W�ט��Ruؘe[q���X�f*j���ݺ��%3I�F����<�M���;��u����\�9@�������x���/,�}��n�\J�L���շȕ!ߍ/�:k����uv8���ð�[�2uZ8�v9`ǣ�]���Ay�%ՎpM�B�qd�����������m��0�����:� �{{�н��v��Ƽy���}U���>�:�̄O>Q�E�̳O(I���z��~*Z��|�TP�j��x�7�BƎOV�s��·�A�UP������;���Hy��|���������߫$~�)���{���ۖ�.t���\��fܠY������b����a4�����h;���Q><�
(N[�A����P2��V�ĩX��[]�����񽞨��F�����{�ė��v7g��^����;0�{���om�5O!e7�b��2c�̝�=��QJp�>u	B���!$�_��
Sı�CX�����p:���a9���Q�7��	lX��b�y���v������z_>��VN��b|�b�3��Dv��D8><��W<�������Q�8�H2Zܻ2���g;ue҃j��0i\�����uG�Z�?ݾ����Ź�wj�nVچ�)a��S����)]r��f�
y8*֎�-��X�TP�E���y©od\��́���%�r�{|��X�)�;���Ų��_)�}�Z7�%�T�G��;�<	Ԧp̹�p̵Zݽ��	�i�>9A�f���w�^;G�J9F砽��J�wSk���/�-��jo���=�.n�o�k�q5���^k�$��5��n��rG8�xs�}k�ۆ��U������5X��P��4����0��̶��:�Ecϰ�q�"����y�'����x|��桺�����$��}^�e\�B���8e�7�IΔ�4v��������ϲ]�&��ry���"�zvmg<u}x��o��r���U��D�h�S�:�-tQ=�ƫ�Zn0K��[��͛��P�WmDwq�w/����Xf�\���>���o4݉i��V��:��]V3�[��;�c����0w��WT�	^�J���X�z��|#�К�f5���o���Y�j^]�uj��>[=�ɔ�p��گ�z7�E��Gq������m=5�hüE���-�G����c�"��ы{��d���-oN��"����v2åv�k7�8M;�{P��r�7��iu��k�]Ғ�2�֧_u[�av3=O �G���Gu�cN�ܯz�`]�J�����Uxv��Y�.׷;,��EGO��t�����%��P�zHv�s*���M���{$ɞcz9m�h�r��B*:Gy��$�jJؓ:�+3���o;��������z5M�m��9FQ�>�wH.+Ff�DÃ.n�d{��{��/��ϕyCͫ����c9�A�u�TB����pj-1\x�mob�R��b�����!7Ck�l&͸V�A�[���^^�j��Qa]A�B6�sSk����� �Q�i��7vj{��[�P�ʫ�q�>N�H�dA[^�p�/�=����������7K,����M���4��#�^��8�K4F_P�(N-}����M�N��RK;m��Sx�n����t�mmw-|F��*�JK��R��6�%��g��k"�+��J��� �0N`-��B�P��UOy]�N��_�A��;(aZ�z�N^���u(:�U�Z���y�*[`�CYҭ�ӝ�3�֊�q��l�v%��������Ӻ���d�׶B��:������J�s�cln�W�����1����u�mh�s��b>ϩ��|z{�>���Qˮ`�8y�=79@I�c9	�i�*Sq�^>�����ễ��8�y���z�*�˕&��킮D.F�`����$͉I��KO��gy�ˌ*6!˶��r�N�ի:��Ъ��K��:�W�3���
9�S.i�����EV5|�tYc4�l�==/#!mo]��=� �0�'P��Tt܎�j���W6_!t{^X���k����oxLu�QP��e�o�.��K���u���}P�[�CR{~}m���眶���EGO��G3}���c;����7ծ���B1󰶱ܷŗ׼����3h<g+�{���Z�P9\*{�{Ƴ[��Lob�����-���a���;խ�DJ�W�c����[���y)�jC4��7>���ges��P�.9I4���t'�ô�p��	�{����Ҟ��,�l+`�G@A�����vZ��c�RG%�%�������� [�G�K ��I���W.�����7�!�8��.�L�RO.G8��\U�o��o;
�9�ʈ��g�(����Z�i��Ύ�$O=�d������/k��Pvʆ{ �6!k����ɓ�1�G'��!�ݘ��s4b�Y�S}2�;G�D�(�SVV代5����I�殂oj��]��e|������i���1��Э�9��˃I�bs�U�յ��X��շM�V��������T��LMnR�+�%b���8�N�e`���a�W*�wѻH;�m�<�=�z1:�f��{Ф�'e�fv�����}4�x?������Q9��y��
���=7�J�3� :/�
�^FW�7����q�&�p�0��&/����ƃ��݃]�k���2�^`����ho��繛���8�q�ғ.b�'�N����>���O����t��7����O�em瞊/`R.#�PW2n9�e�}n�3ާ���y|+M��qjI;S<{�B
� ���~�gˁ�A?�g�1u΁sbua{�.�7�A���Cr��j��D���3� �_~��"����)}��kY����j)m���6�w3Hj߫vx�͕-��:uz>����XC�-�$OV�ͽW��7���zG�ާ����:�z�K�)��5��/�븮v��y���%rM�ka����e[�֙�d�\��흞#��2��̡qR�����)M	�N���9C�$��ڸz�q�c)l �ǯ۝�s�0�����ė�e���y3����D�����
��ki���#w�;���޷��V ���oV��q�B�rQ������?�I�ٞef#Q�n1>��O#��vB��V�&^��Niħ�:��e	�2T�q %5\�1)V�qeqy�(�^�T��w����O{��F��8i�D3z[+�9X�n�m�ȅ2J�pjR7��#n�`�c3fr7U<�z����>��ӣr����Q�u�7����Y�9�2_���Sh�\Q�>�)Y�t^x�w�^�t0ێ��u�x�43���{Ұ�rBq���i٣q	ˁ�ЍF}Q#WH+m\�}V�n]��w&IqD��܁+�*"_e��Eb���e�Wx�BN��:
g<�_Z^Vsǝ
*�����j��T�[,��酰svӬ�uҴ��0(��[�s�땑7Yg/�ךA/ȸ�J�2���鸆�__�G��N��_̐���F�L�'Lm���*�e��~�DtۥJ����u)�����H�j|�V�f��H
U�����m)���Ѥ�lVLñ�<�x\ْ��5��Ti�]�!�6PC63Ι�����®��bv�,Mv7�pn�Yxi	��c�AYݍ֠�<��]�6qB��5���\ïT�#�%��ա�uO	��Tb����;�ףz+F�ڼ�%�.��Γ��u�^˩$�F�U����\_�2�p�b;�~U4�d�E9�{�ڸ�����|:9�Å���J�|gՏ��M�x�X�coꜣ��]��ɔF*`�e�)�g}�.��S�0_�5"�ӑC�<J���S�.ωL/��b�e��A������0E�ä3��g��rSB�cr������&��l������s�o��e&h�R3�n��]wz�w���_�j�*(�O��<���7�7v��l��'�I�3
�_T+ۚH����n�ַ��|LʼX��υ�?	���?�;��@=6�FZ�A_��=_t�MD���Ǡ�T!puUh��~�%�p��c>���n;�>�*q�Ӑܜ;o����#5
dk��=q�_���Ҳ�xlyeg�ؿ(��!�����C2�㋧�t�i�~�H��%�Q8�Y�W'��n�`ks\��,��1��u2[�<����ेq��e�]l!�-��}��%8���P��ӂ�&bs�+����s�1Iח���'Wf)�Q9hHmv= �5��l��E\B�In���h,<i�րǬRd�:�Ɏ���AL�|,ͥN�b�:����&y��֘�q�����^��Qm��38�**����OH%Һ�2�W�)�]��G�g����j��+?W��a��;����J�ޔ|��->'-/H��Gq�>�;c��S�T/Q���@�6n0
��rDt�v�B�pZ�߳�[
��~�z���W�t���Rٛ<�=}WF�� ��`a}�#�b��@�_���i�V:|�<�wqv<ԃ�e_����/�o�뗧r�Q�:�/�N�rn<��^��dϯeƏ��}��c����E�m�,��Y�����_ԩ�:}���m���SO{�W2�]���^i�|�����E�����/l����K���<����zQ>��@^5p�S��2���n�f��A��=�{$l?���}�3�h���<�6~���BqB��Xn�P�iQح3"Rt�K���	~��������:U�4�=���:n,�{��/3�
��q��@%�dG>Y�[��}��ٲ�&��j���[�z��c���Q�ꑗr�:jO2L)�̨ԗ3z�zOWm��)�%�EƵw�it��!�Vz�7�-K���� �=_t�I�Po=�j���xx��{;�_;�l�kT��5hrP@��|M�8u��!���jT��U��@_ly$�}N�U�,ܴmr��)ou�)1-�smeWm�.s#"Υb_�uU��/%Ӆ�"&r�fdPM�n��6��@�iG%\�p�,M��u=���v�A+N��DV�s��IZ��V-������d�ى��-�x�}"���1aZ.�m�a�g{9Djls+���חW�<��g3�m�
t� BQ	Ɋ��7
;�!�S[P��ٙ|����l�n��Z����l�[ە�c�$aX5�B���_3݆Y��K[W��z��O���oc�庫�1�����?^[#y�+�t9�˫����VŦ��ʠjV�]g�=V�>�1��d,��Wl�]V�Y7��|���lfIf���.e���J���������HR,	�u��u��˛St�اe��Wn�]n�R��srQuL�}�92oq�q� )�N��=�ڸ�D��ee������:W$w-����yӔ-^�Y�X8w]�}��p �H�)����dxe5	M`�.�N�n^f��K�(c�u�)MT���r���*\��4�N��:4JC>:�evq3z�	'֘�.�側K�Ŋ���X�m�ܱ���ӷ�c{U<<��܄nΙ�k)0���m��́Ӯ��j�Υ�p�2�n:`�n�J)�&L8�ܳ�K7�_s�	_������©�y��mY���A�e���ı��<��F��q�)ރ�;����N�vS���)����݉��6>u�Z[(uvd���s��T��b�V^\�/��ŀڻcAj�
�Iӑ���!��@ᶊ������F�e�i6ʉʙ������z �M�vu��d������T,fѣ��кoj�B�.t�Nl��� :�,�[Wxo8.��j�7���Pr��1��2�������_R�V�n�B���s6��U�qr�݂#�-��44X}�RO�	�X���w��=uۅ�U(8��v����t��Wuԉ�Κ
ǌ,���+)���Ʈ�&lc"�����ׯ��uH�vV-�H��ٵ�!5��`z�n�O���?>��J����� �v�`g�vebV��Σs3�X�Q$�Ԝ�ο�_`���P��t�=��]�[C/,wC'^�W�0��$��t΀��q dߒʒثԙ����̎�������B�wfV�֌���B@4u�o��Km���Z�z���ݘ�]iVN^��ND_*���+`J��[���n���C 5��L+�X˵��括W�G8y�e�ز�wp�Ce�0}�u��ՊKx���P��
�X��q(l���'^��hi�U֔.;ήnG3�����(Qlc�&];�{�^ԩKj��q�}.�p:G�}Bk�|T��� -�a��Z�w)t	�X�u-�t�w{�r�����א�f��Q�A�}�%P��D���&�Ls���mN�lr�cbZhh
NTh7.p9
���F �tr�1�O'�y'"��-<�s��争v9�lgc�(�2j�rnp�s���y�9��9����3����s���И���ܹ����gc��NESI��[#F�R����9cX�I���(�������6��A����j�s�
"X�Zj��b"�Z�f��MRQT�3�H��Z5�ŉ1�� ����:Z
����%4��t��1E�v0qT�-%����hJb�**j��kC��4LQZ�ڊt:"j�:
j��栶f����X�0$rtT��gl5Mlf"��ED�d�M%F�5����j֨�ݷ��z���GRh�����t)�|t��{i*�K���[
��ƍ緆eq��z!����s+����'o7�7:��S���̞�%�J�M�V��%��C�(��θ[��`�<Zճ�._�.o�S��=0��������L��XϾ�n�K�\<7��\�����mb�<rQ�S���GL	����Upe��>4��Π�Kd����3�G\bw�G�[V�����W=`嘥	e��՗�t]�;�Q8_ΕD�|��k���	�bg�m��\^�Q��3�h`0(ʑ��wvl�������'�>�ۭ���J%��!#�y���A���q��j:�&��H�l	tL��=�&<�O�ɴ�p/�3L�Ѝ`�����N��2�lݎ���=��^W{�;j֊�;�,��R��j{p�UTmd�IH���
�K�ɨلv_z�fD�K�����x�z5�>�w�]n/;��������h����ϥ�;m�Y5
y���-�;Y��+��Ηǉu���끕�\T�8.+�i;�ݤ���ǡ�{���c���=�;�j�C~G��ټ��r�]x,Z�T��a�s,�s�9�ש麕X{:�������Z38���5|32��T��F�eǢ�d1����A�=��q��+F[�,ٺ�*����:��Q�E���T9��%�걆�eM���Eu*�<��_��l��c �}�+�X<]�aW4Duu��"_s��|�t�0�:Mygbtc߷�VR��| OWcG�s����Q\懰�k��q��뎔Ne���P_T+�Ua�����"�]�S��;�眶��D� �]�q.y)>��Q����t,_m��S�z��Ĩ�e������u��g��L�fY���t���,��)���=�}q��y|=���ȵ$��[S3����\�=�哞���%qS+�.+]����]0o�:�>n[=����|�
7�@ݷ��蹽�g��I��_��,_�S���/�EJhN�L`o��1�s���K&�5��Ώ���M�%m��`��-��sHW�,�I�(	��Q�=�>�wQ.�h�p�;�����o�W�x=�ݢ�j����+�G�8y\'�U
�\�k���P/�i7�<��F�x�y--� ^�퐫�h�q.gy �/�su�I��:��ꐚS%O S��)V����O����#��~�����b�_i�Q��b�Q���|\�Kg"�`7��.!ϙ��2KF�5-�a��G
��W����^Rx�=��N+�Qѹ��q��e����'/�e�l��#X)�H�|���y7����l�Vp�eoJ-d"�2�>����̒�s��rn��HamjӆM>T@����X7�����ߙ(�i�9V�Z�=׸�[���N�gI
�D�Al�J��{*^���v�ڧ:��][,MT92,��E!hn�<;��������x=q�Ӌ�J���a��o��:�7�z���H|�]ы��vh�r�k�b�Yhe�[ۺ��ا�&��xa�D��T���:��6�u8��w��U����RtN'����=+���ɗ����~�b�ו ��'�zam��1��<r+�i}�L`Uᰶ ��j���u�,�vڥ��ct���;�X��T�^J'*��Fd�دS��G=����v����K�&ˎr��Ҧ:V�����~�ܠ��R�X����9+�RC�}4�c0k�������3m
q���-��re@���~�<�'����m\o{�w�o�7��"33i�܁�0�
GO3�8����L�r\���.���d��b���2����3���ذ�X�:'cNn��]!�u�>��o�(��e�@:P�_�T^�.�(�,�yä2i�+�(����7��p�Ү��i���T��;�a2K��L�lW]�
K.��R��~���k�Q}Bd���	H�{D-������B�G<�$�!��~T��6Y��)����Wu���3�PywXrW,ׯ��A)ٺ.���ܓ.��"EiҎ�y<��W�+�6ӹOv�.E�F�&�n��te�ɪ��4Ù�]�&��^�0���;�74���et�W&K�Z�Y�]G�XU��a���z'+����#��n=�����|���E�ϻҔ��CRZ��c����T��UH+�l�����!�
~u��:��ֹʷ³Ý��{V3���뉸t��
�g��7'�<w#�g"�(��X���7��_��0ş8��'��WF�l��N����
u�`+��-��m���f�6��n|���������8\��t��	<�h]r�gp)a��톺�@7�Y�\�WIU/{v�n*��'��J��x'r�s��1_J�tn�+�ozPi��ϗN�:/���{��u�2�>�%0X}�`	��(�ρ���~��[Y�Փ�퀅,F���okvw�&Tz�����Cj���:Kt����r�\kʐk����������nc�ğ'����%T��9�/�Gt�;��ߒw|q9�Q�u.�X�+&}l�x��(j��y��y]��龽'�a·q�c.+��:}���m���SOzq\��wpz����?E������_�{
�*�Mf��U�zZ�<_rr�X�8�S�8.����Τ^5�cҩ?0eϙ�mIvF�������חP9u-Dd���`���d"8	��ѭ}Kf7����*�V`���+�\�v�w��8�{�٠6�Z�O�.���9�W���V�v�V����k���wJX�Yֻ,����j�`�i�K��Gu�����YO.�\���9�һ/�츿w�����Ñœ�pf��(\W���R�	@w݊�2=��J�\њ�v'��ل���]u${��iO'�geN����3ƌ�B�u\o��@$�r�p%�ݽ�ѳ��r�G8�ܬ��9�r-���7����hd�ĝ.��ŕν��r�ALȡt�8�c�)YqJr�bWp������W�T%�+�q>�`�=](v��6�Y*<�3u߯�|�ި��T��c�}tY�J�M�V���}%���d��:�h6���\M[�q����c׼W��}�3�HS����H��XϾ��ۧ|0r�KN2<p��*����ћK��5��q>j�u��<z �d��F��O��bw�G��ա[�{�[���Oz�l��FV�>����ܫt�x�'M�uP��k���@�&9�>�nW�F��;�j��L��ܙw�jK���oZr�~���ɶ�h��iL�����F��~e����u����r_��{���K�7m;���&=�˭ɴ�p-�`>F�
�])3�� ̦}�_�O�>:.^j��YX��:��H:�P����-1H�N�����Y���
�O{��i�I���m{���<�^�ټ	=��[�YO&�8�Z�ȼ�\9*]�:Hd�t�[8Ю6mj��?�J��)S�9��q�`q�'�V�uJ87��
�\��c�%���Kө�Co����dɶ��ЍP���2w
��B��J��.��^j'�e��rXw���R{�V=�/ѻKM����{����N)ɸ� �e��(�;����'�=y����G�ύ�,��}�+��xp_�\�I�}�H;���c�5O}���٩�~1!�;g\s���h��1��]��B�+V�����j� {Y�(���js�ُ:��vD�u�nq�_G:��}���W2/�(����/�aez�	>�<�<��說v�.�W��\�)�#L_y5d\D��R}�=�>�Gz#�_Μ��r��2�EMi�/�ڴ����ٝ�3t�L�*��f\p1�&��e�}n�3ާ��y|+�>��ٶ��*o,fP�D�L�pN��L����T
�Nh.��y�ea���g�M\>�1�����ץN��f��{�p֒��&\P����f�䣱IU�������b�ur:���%fC>>q��}|�+�rx�I���~�{��=�>���K�o�$Er���D�~we_#�#@��<���-49_P��k3?]�;�?�A�o��N2QP�-Fي��w}�����iBv��r��̑A�2c�1��X.��ҽ���-v�3��H;���d>ָq�ԡ����h�]��j0��q��ɳ=}y��ϻ��{sc�&_�.��{\�~��R�W�\D�a@�)V�q�<�ɂ������vȼ����w�[���<��M�}��+)��n�i7�ԍ��RP�J� ��6d����FwU��k�o1�-�zV`u����N�>.}���9��m�zß34�I\LN;&_�FJ;��u�T4��,�"g�����|tn|:S7�>5mu�6��%�C��%�>^/(�P>�{m�ߡ$hEK�31��^�f�W�v�ޕ�k������;4g=�GnU�o3�B�*�����A��d���2C�~�0K[{+]}��u�w{Y�U�rǐ�g�3��K/�m�ou��nXo��X�yRl�z��؜�t�0�t�/�gzr�����Ү{����Pp���y:��؝ez1߁�7�b���H��J'*��Fd�y��_`�zn��wp�KK��xNF)l���V�S/�O��~�U<v�~F\���K,�d��z�38���p�����^��$�'��ʁ��C��2��[;ͫ��s������[s��wK��]���|�U����e�}�N���wN��Ļ`�>|�k5�[�F�oN��A�ʸM�ܵN �h�m��&�2X���v�}�0�����\�VGSx�5O��Lg6r8�E���S�.ݼ�u���Y[���S����=Zܛ�$���5����h�7��K���%��5�p#�?r߱/Պ�;Γ,}N�;�0����y�DƑ�Y��w��U�t+��P+O����:�"�4���1�z-�Ϥ�]49��1K����u�:������9�����|g���{���A�;�}�R�?NWS�A�ދ��F��<��Z>Oh��ݠ��:;E��\Q'��0����}	�������� ��}J�
.�ۉ��+x|Ԗ�}�:�y�#�
�p��� }>z��� �{m��w��K�p5W��-�h{�Sڇp��q�S������ۇ��eÚF\�!X�������x���#�T�[��e2�d;��up�Jv���9�#��1�u'���!o�jMŎ���� ꩙_��Qj2.w�Q��ԏb��˄���i��O��s�I~@��f� R�Q5�T��3��;�+iѿ��+�oѽH?L8R���Q���j�#ý�Rj�/�̰1���?\��X����=1����S�?L�W�S�O�ՉwgW��:P�5���E�X�Xn��E<��D�n�3T�5��IS#-�F'5�EQm�1�2���xP���E���*ԣ/Ơ���V`�n��v��V1Q�>ޤur$�2`}\�����Y����J�9�P�c5���s573����gh%����p��yLsj���:M�l/ЎU��yRGK'��|���c'2��5�y��9�:��7Y=�q��Zw+��;�>���:�>ĳ�.4����Z����N
>�uv�� ��88:���OJ�p�n�f�����4�ǚqZ�ϵ���aH�0(݂{Ӝ���|3=�Q�~�4P�3e�}>����d�W�O�ช����:�^5�c�*���������R�h�����q��6⟌�E������l��-����kVV*@}�(��vt��Z�7���f��2��Z��3ޥ\3O�=���:h2{�����+�UưK�w8ؘ/Z�svu+��4q�KDȍq�YS�N�A�������Wݾ�w(����<��2�4��3w/3l���
A�.+��,�UP�K���=���Cۆ�}�1��'գ�Q=^�ø����vԩ_�&_�,	��P�*e9c��EJhNDjV��Iei�=���<녬۵�Ob�{q��=�S��S�l yX���f��E�>g���p������+u��ۤ)O]�V*:�*(6ɭ��C|�페����1ь��{���7:Z:�:��{fu�ҨA��sC&�F=(�G��A9]<��ei�X�bQR��H=S�@�����䧖��V�{Ÿ�,wd��;��
��7;u�M��2qg��z�?�w�N[�f���}�@�
�Kd�ٞjr����й��K��칭�{B��I2�?�{o��7[��<w��Ө�FJ5D��0y���m�����L���+[�f��f\U?-�ͫC�]q/��Knp��q5
e���!#pvHg����d��ܮ�חO�Qt������7Ѩˎ]nM�n��i�1��)^�og���YS'�y�<��i�㡂��.|+��u��v��X{�On�m]Ѹ�d�m�Йиpz��An���j%�۰>���$��U��:6�mx�YS�p]b�b��KM꼸^�N�bq.L�s�22o�Wɮ�g&��ͯQp��>:=���ᕁ_�/�U��ݤ�n�1�g���맏|�;�H&�F��Ξq���w�«���(�˃1ΠNa�>��jU`9w��k�^�����Բ��7֠K����T��7Z��4=�N���ʘ�R�ݰd<5�������3�jn��O��m��L���L�'�i�*=�Y=<��S�<�pn�V��t䝻��Q� �����Id9Dg�(�Fܩ��++�p�Kw:--�x�o2�4�2�]Z��볖aʛ�Kq�[�Ӷ��t��jw���n�/	�6�N8V�/˃�	x����#��C}:+��%d�����Cp��;Tù� ��u���,(8\T�^���`Ԭ�K���|��5�WF��jU�C�io*\fAY�-�	��c�䊂���]��B];Η]x�ԥ
�K&]\�d�4^�����R?l]Ȥ��sv��0W\�RC3���l��P=*+�z�4�� /n4m|��.���X�ST3�p�svc�/�7V��:�v�VurBg-����I.&<�����5�Y�N隫{)���Xl���k��1���`hΤ6���.�|�r��z�c�Ӌ��λ� �%BoZq�������ܝ��R�����Vh4b�$(��&���
�ʞP:ƙ�E�򫊲u`z�P��LwT6�p��'ΚX~�U2��۰_K�e� R��xD���x����s7���.jo�c�>ܙ���Xm������y�`�ǰ�Î�;�Ԛ�OmG�#��Ww��Q.���uo��\Ƥ�E�m���ά�D��GL�Y���R�Rqca��u ��ДWX��Y8�Y�����[�5[�u#�����#Die�N�S\Z;�"���ܨJ�c:f=ɺ��H�y�Ⱦ�%�6�	ոeY�)��vU��g��h3�
���܌�k�.Q�f=#�5�.�iE}ԜڻW0������T*Nk�m]S<Έ; 5{�իL��[\�8�b�������V�'WK�p�Z�*�ҧ%���LԶ��VN��	��}6T\Z5\�Ȭo�
�R���F��۹����K��8ԙ�LT�P
�3�q����m+�+�mè;]*%et��36��U_5/yA֧ywX�RG�Phv�tḩJˋl�T�
F�(�(��C456��=�G�R]%C�u��"�f�� �;��/u�!ѵ�4���M5��tP�J}7�2��)��͖,��Uǂ,ֺ�T�$���'9u���^wT���7d�(��n쫺{�X�Iv�i2�v��5qY:�TI-8/@��ºm��	䠡Hf��!q�N�M�]f\c�v�lc�E�u3��CVL��t��㼣�QV{�u�^,�7+:߈t^��Y+r�afn�]M۶;3)ʽ[Hk�UwC+v;��L.P���:�w�-�lذJ	���3��mwq�]��Q:��nV���d
K��eLP�!>�P�랈ISU�:7�E�[Ī�VYR:on�u!�;��ZUھj�.mմ��Ȫ�<ѩ�����*EϹGh���2r����q�i�[�	�CvM�}��˪%�*u�zT�3'j��#�0ݸ/`�mu�����ev�)��c����p��:�'��͹��E����.���5�e��93���c#��X��;�ْ�2�Q���|t�����W[*ۙ+H暗P�seN���!X4P$��llEƣX�6q�[9�#c4��E�[`�(����EG6b�(���ii"�( ���j\ΐ��i�LAk%�I�4A��)J�V����A�i�9��Z����(�A�[`4PSMR[m�1L��������
�����$DT4�lDQVڪ�����#F���lQ�1h�lm��kT�IQ\Vق�1E5�i�s�Mls�#�cTZ1V�5MIDQTEbĔD��J ��ڱ5QU�(���ET�mQ�
��nlQrb4�j�I���C���:��bm��k7.G*�4[Q����j��h��*�b5��i�PRTED�IU�T�V��h�TDMIEL�8�h��� P�>�$P�u7��s��K[ѹm4\�nP{�	�0m8�ih��g-���tX�����ZPc���T��v��v�v�*������۲.��w���A�Qӓ(�l�F̸
�c�M�9L��P����5��fL+/d�,��
ޮ�;�w�mܛĒ��(uD	��_L]j�T�buaz4�`��tX}�7?|PM?�p��s3�_rub�>3�\m�g"ܐt���OW3��QF�)*�7��=1l�t.D�^ec��$S�����5p���0���QY'��(	�{��=�>���K��������gdUo`�]	:����h�k��^O	��J�\��}�@}Pf	��ZK�S9O���9[�~� �i�l�k7����:}�+)��n�i/�͇T�ҙ*x ��F|on��ae�{y���2N��n4��Y�Q�o���;H� ����C���X����M���lY���8��}{�YtOaq�x��&"yW
��\tlqL���ˆ�ܛN_Ϝϙ-�IΛC}F�M�T����t�ٶH��Ӳ	��f�DJ�f��W�v���-+����0�Ѯ�����������8�wl�{��5z�ȭ��$�Nǌ-�/�
��T�߷ik�XngW�$?�C�����%xf�
�1�v�1Ov^��g_������X��p"s{t�B�/��JM���p�ocE�u�����G� ��@p뭚��>t�l��ȳ��D:�f t4aʆ�-9�׫�*����.Gzy.[5Π�$Ƈr��������+��
fۖ�w�C5�H5,��[�su�:�8}�:�^ۂ�}&���^ڵ���7����SU=8��g�����o�C:�R=d�r�Ù�H6,��#���y�Q�LwާZ͊��IӀj��n��Ҫ��j�O�]AیY�F�ܴ<�ݿ��Qc˅���;����h<�W��}3�>'�<n=2�v5P�T�e���Y�|ڸޏ/;�� � ��V�:+�.h�o�<.��	b�gG_�.���A��&Pp1[����j�;�[�ǥa���5Y�+�o�p�D�(]L�3�B+�V���7;^��׻�������\3�7I����G�<g8��2�C$�x�U8�S)�W�"�Ղ ��[���)�&�A�[t!������Z9��m�A������rQ�d�^2�����5}�_V��8N���Yj�7��M�V�KS�r���T��T��D�gP.�_��48�� ���@Lep7g�^[V3��)>��t︄|�a�nN���e[���e�a��~v1pw�ۡz�&!Dʡv���B�q{"�q���A7w�&��Ub���%Xo�]�UΏg�ȯ�F��ӿB�݌�;�t�A^J�w1���`�e�U�f!ou�%|�"���y�����;pT��[w��;�՘`��=շx�3{��]q��<H6T�~�TD��h7��L���S�qt�w�����;)?���?�VZG��~�N��êFEB�(�T�W�� �}4=ʹ��
Xw��b�"�ϓB����h]
]e9�2W����Q<
��&c�����Vӣu�]�u�rV�)��z�����&^
kz��i�܋�j�/�3,y�llEy��0k�Y=B��~?eS���	�ɵՂ��5�m��.)�Go۷M�{lzUto��
n���G*ƿL�œ�=��*蚞�����ӎ�KѺ\9]un��l�?"�z_m텞o�pn�r|�`�!,������]|1���s}����u3:�xk��c��^�2�+�i:}��o�m��Q��ӊ�Q�nƵ�sRvU���5�E���������N���d�WS�8.���9�Τ^5�`����LeU��=V�{˞�M���v��~�n)��j�[���42�����<1�0?w~���Tn��޷w�&ۊ� 8[�ё�i��N�=�U�4��J,jڞ6,�JW�!�g�5��ʻ���?�s���R����]���f �sRW����x�6�������K�}����kr��5�||��r�TC<����ǚR�)�볤ذ�V�{��=;t2���|�cT�Sv��֊�ڻ+�p� �e�W��f;�{�D�H:�'CN9��۫93�l�k�O;H���>���Y�O(�}��G\5d\yO%;�E�A����?�V�>�hd�ĝ �qI'�h�ٟt��/Q��P��g�� ���G(����=���Cۆ�}MSntvw���}�W/:.oYvO���'����L�,{�뢌�4'5+z}����%�|�"�b1#!��^�\yq�W���c3�=p��@�A�q�g�e"�ڟ3�M�	�N�`{ޛ���]T�}�qw����	Hö��N\:�aX�(�t;���H�ٞjs )��n����θo�+q���%��r��A~�Cr��n;����N#%Y�&&y����2��g5�s��B\o����dƋI�C�����3��ۜa��J%��} �H��}ǐ������_����6��q�e�����f��Q��ܛ�7\�4���`
�I��b.7v��m7�ur�t�̤o��wgez�;g�Ҵ�yP�Wto�y�&�@k����2����*�+폃+&K!�9.8|n���b��}E����;�'w�7e�4���p9V0�F;��5���`9�U|��wa�<�
�	4N�]e�Q#/;"�b� f�/��ǕK�F[d\��w�/��+.K�+�̋I�l�Q�Ѳ�h�/n��ï;��rT���'�e��}���u����<ns\Kv������5j��{����vۼ�q�����ѓ�o�/�U��v�u9:*gf�>�Y�'k�����hXq�o��F7C\��Vc�
�W3g!���d/�'t�`VW�NS|o��\&*f�U��I|��� T^5l.���8�>uc4�#^��2�R=��g�ax����.��W����;��ҊqJ�M��"{�ǹ+ ��ʘ��I*�ގ{|/:rN�$�+��v�)[���l�-����p"}e���wN���[.Gѳ.���7�S/r-�&{���6}y���t��ｊz<㮃��ܞ�I;Q2á3�_�2�b�U��1:��]0|�2�}>5+c�'�:�ڕ�g�����Kn{�>�\w�x�$�(	�����f�䣴�X��7��n}�����P�*�! ��=���j����V.O��=_@@�$\d�wL�&�9���X���'UqN&����HR�xs�|w�p�NT��.J5D����߫�t����k�f>%���ٟ3Q�o�O�%����e>;��h�o玤m��M �K����p~6���7��l�V�WG�=����;w����s�&�z�)A���HC6v5�� �E!w��.��8*�1��[wơjJ�����%��fZ�	*��-Lc�����ש�(9�l�IҮ����wL8g@.����h���e�yx�|�z�k=X}#�}����/�̀�7����Frt�P\�Ke�O�ߛw�E�7U�|9V?c�3f[�'ȉ;�i#bS�q]K���ҙ�|j1��'�9|K>Ʉ֮~���k(�zN��XC��EqGf��s��ׅJ�f��yWi�}�KM�tCZ,m*^�����^��IwF7sh�mˁ�ЍFEDl�&��v�zalf
�W��b���8u6��=�\.��u��O��J��;�uT:<�3m� ��s���d�@��ۈ�c���Ug5��={�ª����S�vGu�����ǡ�������~M��U�����v+"���{��7]����^�;��>7�L�'qL�����D*�xO����硫Ѕ��h{��߳����Mo"�x��Vs�)�Ӏ�ˉ����+�X@�O�ʁQ����B���'>�:�z�����ۙ���\���O�e���F�ߦps'��	x[	h���pJk�~�b^���
�Mʗh�^&����5�$���.��=�W���D^��Y?+\ez�qa�������\��Z~|!�CY�������mrX}+e�����N�������0 ��>�L��^0T�Ջ���9�:��᷎�X���@� ��C�;��uz�27P��*��<�e	`��P�2x�k�]���P`v�,�Y������n8�n����; ��Ή�i9�쁹�sԁp�t7I���������T�(��a3Pg�c.q�K��m��ؠ�VeT����Gy��Z>Oh��ݠ��'�ЬE�F�,��'3K�5�\���y��{;D���Tz�+&��j�7�7��S�֤�;��@=7:�e���)J��3�U���.o���� �_��ýL)�h{�E'�p��q�8�i����
y90|w����3YYnG�ό��x�Az��DOҕh7�S(f;��up�D�i��t-��d(ʤǦ��K��s	M�N9�d%2Q�����mG>���W3����_�l)�g��2��j����o���Ye�l��C5�V�&�ʓ�&c���+e�U�A�&�d�����y��ۛi���O��o��2_��?D#q�R~�����2��~x�k<S������ݞ��;��y�ڇ��=�=��>N@S�7l-M�^T�s�S��D;��\O{e�>`�6F�J��K����Ҵ�W�;Rw|q9ɷS�wG;��G�l�Ǯ�=�Q^���D��j���mVG�0-C����i�[�"�o�i�n�"u�8۞Kt��T��-lSgV�n�Ӳ��S�p4�k��e�Q=â��w1)f��ӝ�[����hӛʂ���X�m9�h�{�v�Ҍn�u����5�(�������9`񯏥���_��c'�i8s
e{m\?}*i��=w�Tg��Gt<������U_���2����m^R_��X=�pJk��|�}v��5@I+3'<�}��_��XN�^@�S�g��X����1y~��~E��~2�.&��_B�|b��8����z։:���P��2%'LN�+<)ҍ��Ԣƭ��~��)Y�𼏴�����8.�[�v,��f��J��� ׾�T#�y+"��Jw>�t��E;��z'բ���Hˀ�*޺��/x<�!��@i~$�q&٨2��|n�T��%w�it�%���ᾙjX�V�(�>�
�絎�>��d��tt���qS)K���)M	�ԭ�|K+������mm+ޭt$3��nTv83�U�`�� >�2����������XϢ���;#������\�fF=p�%���oZ㑮F���q̣`\�k���Pd�[$^��S�����u�d�%�9�]��S��cG�SV������n�p��N�t�&���}�@J�N��#w�+�,,
b�l�����{u{A�3�FuJC����^ogrX��z4]X�lp��|`��60.ӷw��+�O�-�+N��mf(�Σʂ5�*�<��-��5��Ls��z���r~��;j	{�9���;:��f�$Z䰰����*S�=��b�˒�����MG{?u��^���j��ޑ��j��C�\K�C3��ۜb����e��4�W3��oF��Y�֩TqyO��&$JT����ckz�2�F�9u9=�n��f��F�	�j+�k������n�ܙ},�(��6z|*^�
�O3�v7�i��=�k�Y�u�'gގ�w���S�U����U�=���H�L���Gf�>�>
Oa��Ŷ��7ii��yp���N@4Gh:��^��Z/�ÎJ)I�� �yf��3�q�����VT�8.+�i;�soGgK��]K����%اn�p����G���k�����^2����ݰd/��!�xe�5u�:�Q��N��V��L���| �J��N�nq�Qάf�k��y~���Nd%uL��F&��1gi��P.uq�7S)���H^䬋��JO�T{�|���+�����C$Ƨq7x�gf}f�ɥrIQ�鞉;#�L��+eq~��*��tɽS��Tr;~1@�C~�zޮ���G�m��U��}9u�Ip�D������.+U����it��A�+=��x)i~�-�P]Hi��Q�w���#
���M+!슞ۛ�s���u7p�
_�����TtsP�hf��9��0���݉�<�&�6�vN�칷/�V9S�����:�_6����bf�a���'xW1+
ҷ��T�d�Ös�G��v>Xg8�G��7���e�C�=\Ͼ��uLZ��9u��4��O_�,��}�\07����GnW}|�+'�qd��2��{�Θ3���uw��T��@+z彺�r�葪�����G�#];q+��T���(�qx!�h�L���߳��l��^&�fZ/2��8�TO|���x���r�M��R6�uHOW��${s0W3���^x�=.#�zh��1-փi���DQ�o���;H�oKe|��<�j���ďk����_�����Q?��35
d��I��}d���\WR�r t�n1�ˆ�ܝxV׾�v
～�lv��~y�t�����`�D���Mx̅��VAg�5+.7��O�n���	�����,�?-��	�f��.�#Q�_l�&��v��ؗ�+��{5t�q�|��v�{������6��z��!�I�п'AL�7,���,^���C��P�|y�c^�϶{�R�^q��c'��/�R���0/m������#=�V�U���H�DGh�����Π�����bTfj�N�f�f����HEc�R�°MKA��/���G2���c{:�ZApN�1\�S�}�}���f�̵�ĭFM��6�����z�Y�u�Pyӓ�1��܈�P�J�����xP�+���� ��ݔ����F�m���S�h�tZ|�Vg[� V�묮��L���L��uP[}���*� Z&�@��]�r,Y,�����W�H8�1R����޹6�_
_'On��[�Z�
Ѣl�+i]`1˗Wa��Q2F�)t��E�D�.�ڄ��e��I��~c�YX���kfS�2�u�*�_�p<�r�E*mTGJ�u�A���P +����ݓ�f)�-���s�ɏ�쭂:�^nAfɮ�y�!���bI*n��k��F�k��l����\6�t�Yz�X{U�r��3Qyw�$ސ��͜��Ŋ���4&XH<�8��{g�wJ ��+E��[Y�o����w#�&�]��j�����-�f��o<BR�t]�¥��9��{����&�H�E�0��	�+3S#.|�\������,]֛k����*� �j<��O j��=l���IJ����7�z��[��6#���,�{�Fh�V��t�e�콭R<�w�O�|�gG�>�&����,X5�:���f�'2�;�⯹�𥻁��)��]��m
4$�����ŀ���2�	���-�i;N��풘�̕yB\���S��сU��G^�=�&�m�6L_Y�(�ƾap���8�����@:��L���XEl�u]�@R)u�3-|;���JN�YϦ`��������N��3x�潍�̙���x�r��ܰ�n�:�U����X�R�i�ˎe�-"�+�V�|�Z�FDc�4�Ed���p�]���:��3�-�e�Ǹ��#�.�
X��]c��N��&հy��4)���Q�Ŷk��I�$�ygx�=O	*r���v�-�n�=u�2ƻ���/�{���5��T�9��!��3�q��g��T���N���K���\r�u������.o\�JE�Ih`����v�T�z����[�}����4e��!̝�38U\٨)��Iuuv���8E`��
W�ʬ�._r=e��3M,�n#���@kwR�%Ֆlw�v²�$�Z�QgZj�F�ئ�-����5G- '_-��j��+���'X�2�+��J��*�*t� ����Q[��Ԍ����˺�ն;{4�+|�f�{�\S��p�۸��N�H�4�b{ײ��8��7H��,@����C�칑��N�7�#��ծ|z*c�b�"��Fs�ҭ�&��;tfۛ8�(�ˑ8?���̔v|�V0K�&H��O��ȵ��+�IV�J'S�\�VZ=ۖ�C`�,vJϮlV�Ӻmn�b��epU;2T0۶S�a���@��!u��+pΨ^��Q �Pn6�ӡL�ꨍ>Цā�<��;�8��{�P�U
�Z4pCM6ɂ64h�͌kF�F��ӂ��mU����(("������"����(��h���H��M�SFڨKY")4�V��Ej�l�TEMZ�ATն!��4Dh38�kѶ
��Q5CQ��1Um�5����"�"�Ӛ4i�������(�&�i�[�"�&#Z#	6LALN�*����"���[���"��61cbт�b��S����؂66��lV"-�F,�V6J()��V�h�� ��F��(�����S11UT�ljZb"���*���ӈ#lX�Mi�Z5�QAU�T홧��&��4j���3$5CTUUDQh�m����[Mrs�QAs��7-͹�r���g\ڭ��E�nF�k�����O,T�*ĂLG� G��+у&��릣UV�R��tf�fR�mY\�Y���N�ح�t�o\���/�(��f��O�r�kZ9��X���lMi�rLs���`������Ą���;2��p��ҙ�Ҧ���p�js��=��h+U�^�ܽhNN.�W>��r�Ö{�`���+�Zo��OFL��T>�U4�d�y֋I�7�3����N�Ԯ7�������d��"&P���.�	*C��(�
���U����]/	���M��?��j�� �Q3��M�,����gJS/�l����ɟE��D�{�k�{�h�V���c���Hg��L����,3�EyvT�b�$��.]f137O<{ٻ'ρ�H8��#u�PT�]�e���Z9�{D-�n�z}��tu�����i�v������q���I�3
�u
�f�*�Tz)���*���RZ��c����T�S[Yb�K����uO�@h'�d�9 '5X��cJ])l��9I�Ĺu�z
�g�����-�C���>���P�Ϗ����e�i��2
5�G.H��*�oL�P����x��m剾~w�C�Pl�'�7:�hD��qng0��m�N��dd)��I��m?I��B��U��D�;w��b��>�����)nad�O1Xʔp5�9%�JHV����4�QE�T3��	�Y�G�X�)�l�YM�c���jId���2��b�pQ�-��F��V��+qL������n}���nh|2e�-�+7���������-�O��=��Ϣϙ+�C5�Z��I�&9�	�
��f���(oչW�}�2�����&�k��VC�]ȿ��w2��4*<|��A��D�Fg�X�P�i��o�ʕ�B���Y�Փ���7n�����Cj����N�Sm�K�ڸ������H_�әk�B�Qs��.��g'î)�a�����Ȏ�Zw+��$������}>��9J�a57oy@�٢��o���^L��P<k��C���c.+�i:}��o�j��d0���E�e�Z�tA/&�s/{�{��^Ӱͣ>7Y��X���
��p_�=_�͜�����G�˫��� ���W��;`��X�z���8�e���D�_�az⇭��لG���f�y�S���e..��D��,v;L��$�.S;*t{
�=���:o�,���+���c�f����&W�q�Y�Q��H�k���j�u�<��~S�N�[�{�w��7:��e�IV��X��)M�a�r*�Qq%q�3�⌾7��n1+�^�����,�{P��\=��ٺ���T��h�tvȖ�um�B��'(T���˦'TW�\�or�������s����'�.��zI^|�݌N��jړ�Pu���le)ֺ�I���I���2��������H����#B�+�+�����kD<6:�ݵ���k�pkUl�ց�}���]���(}0�S)K�뢌�4'>ԭ��Ó�췌>�]��m��"���/T�v��\-��|��l= �P:y����Cж�WYyQ�]'�\��.����<��\r5�ö��N\C�F�.J5�@�
e-�c �kb㇣�7�Y�~�t��9�O�=-�C�_����0��x�'M�:uP��x	aqٗ� M�3���}^ƺ��F��a�8�(����F��ޑ��&�D9uĿ386ۭߝĤ,،�4�8�{���}r�fq�#x�$�Tz�W�}�p����Q�r�rSs���0;{�>;^z\�n�������6)�#n�����:*�#g����7<�Y﷥i�On��wD��(ֻ�;���qk���� g8f�hw2}������l9�W=��-�/ѻKOe/
�O�t����oY���g�k��w�=�S�~r���,�ixg��K'��`������h	%[ŀ�4���j�X	/���:��=�x�5O}��k��h�
	_�|n#
'2��=��^����g��j���̱6� �'�*� ���sX%�)Z�r����U�ՈZžF����J�od��dzh��]��������[��;2�#��mjE�/5!e־�:��fms�ٖ���՟1Z�t@р��)\���^t:�]�R��wg�2>M�A���G����Fu�}�[�U;�g!��W9��;�k�����}�.ۥ7�;zs��3�ۙ�fax�S+�Xd����H^䬋��JO�T{�RS�V��X;~�P�V�����,�����<4s�u�2�h��t��9[*GIp|1�&��e�s���funG�Qqa�a���w�G��h���$�K��A-�SK�*�=�M��Մ�e�����y����W�jK�^*{��l����xϴ�G�4�r� >(z*z���G�b��_;{���&٢�U��i�<�:C�G9�p�f��Ƹ�O�~�z�޶�ݞ�}Jq_~�C�3����D����E¤����G�5�ï'���P��DU�R��Jʁ�~��ط� _���}�����+��=�\K��Ê�|u����<u#log��*n,�Ow�;{����<I�@�#��p�W�F���cܝwg�[$�/a����>�ŵ��4�ܯ@����S$�6jR7��"e:�WԸ���t�o�|j1��������p`5�Ǘd�̱A��ɣmƤGE�;ţi2�6{�8�Վ�Ffp�X�u�>���d�s�,��\\�:�8�E{�C6�S��қ�A\b��vb���8 %*�[g��s�z�.�1v��	I�k���e�Q�h��-��>=����>h���.�Qd�%�#XB�D����|fc���
�S�к��z ���'�0}Gz��ݟ{�e����Du��tb��f�e�Ƅǣ�$���'j�ؗ�)�W�ˎ6��Wgn��Z�SR��d����I���r�7,���,^��K'�b���/{6�ga8�u�%�q]Y������Dw[/�yl{檞�F'A�X��Ι���0��������V}�\�}(��|6s*�_��V�8�o+��
���Ӳ���|�����(�ʢ�ۈ��p��Ϥ���`���
��Ss:r*g�<p�{�z��y"�Ͻ���f�G�/a$���]t��6�7�����i`��9)/t�ѯ����^c�&�کߺe/e����{}.@�7o��n�,}N�=����#�vT鸲��(z҇��}\�:��Q��e�.�P��Ҫ���LG�:C<�&{��������O�����4���ǽY�~�qq}^3�n��OuЎ�[���h�{D-����D�tuCv �����ي�Yt9<D��g����NB�ۣf*������-%��W8�v�M�6�������;.���͚�k�Z���w�gw\��2L��[� ���(NvJ�W�3l�ۺ]�����`f�U1;6�PbL����Q���������k��Œz�2�}0�[4�Yj�7M���:V���-N���hn ��g%�Ѫk��r=�>��u �QP��}e"���gR}q7�}�޷1;�ʳ*�5�/�|_�q�N���e��f��(�tǪ%�)V�ze2�`S�v�.ɩ�u0.��sY�v����C�"V�#����d���ͻ����3!Q�T�Wh��O>�ػ��s �r�+�{��N�����>�mu��o���ϙ+��d
V�&�ʓ��|w�1OM��5��+o<a�*�7�ճ~�7��o�����]Ⱦj�/�3,~���?\�ztl��P�����������_����Ml-r���n�-7����]�t��큥�8?z}�ut1�wy��|Tu_E�o�AjY=_����'ï�u�n+%i|s��Zor��	;�7�sl�Q�P��Ya�|=V��8�`����zVL��eƾ>�:PŃҝ��%>~�t�������q\w����u�����q;5�c�6ⵕ��������fџ��N����[S�8=�������c���ʩsW찯��/���9J��w��4{d��w�Z���R��_6���f�i�|�*+�L���zk7fN�s.���eK
/��6JK�6%3O])�s�n��͂�ġ��S����glf�ا[jS4#ˎ������v�;E�>����s՛w�K�|�0*�C�I���W��/ߴۊ��8SӘê��#+�+vҕקs71��~�BQ�."�������2:)'l}N�=�U�4�=��S���=��
<Bʞ�����|C�?2v�23=AاT���Q��
�<��q�<��[�z)�9+���,QQ(������AXo�R�\�'MDIl���F_��� �bWp�9~/	g�'�T���E��^��$8�z\R�C�Ύ�l���`����C�u2���뢌�4&�&Lz1N`���"d�E���+O�{%�y�}��*��x�A�|e#���)*�EO:�N`�V[�;��U+������*w�,t���#��q9n�V.J5�@��5��sg�Ϯ��=ޒ���̀�G^'|4z[V�������7[���q:\���d����Q��3ظz=���R�K7��,���R�m����Ջ�G��ա�r�lN��@��w<2����9b�-z8�e̸r8vH�{N��\r���������u�6����:�t���tb�L���x���Dn�D���w{��r��i!��[��IG�1��/�����bu=\i��+V.�ŁN���U�rf����Ne�c�fd��;x�P�ՋE>�,=��u��sz��Z�����+p��#��m�y���{Z?;�2^+��;�3c���3)����Q+kO���;Ҵ�F��؊^v�M^yl�[�I^�����&M��hL��/�&�fٯ����>
�{��m�w+>��m=p�NUR���j�_��w������\��.ۆ�,�F��|o�,��]��
b���=΃������op�h�t�i;�ݦ�{n�0Լ��N��Y���^2����0�s�}\,G�Y��z�� K��Դ�S��3� +�ƭ�D�w��Cu��sC�w�{\=����-��J�3�~�w����	��9�f�}0��|r*e2{�a� �%D:�J�U힫}����VђN��gH�����C���x!9�%Yf;b�W�������f�mV�8�ͯ'�����y�\${�O�3n�d���Z8$�$�K��_�zW�/�1qZ�7���T�מp^{���g�~tX}�g���������D��� =(V���r6�=5�t����t�v_��G��%V'S�0s����h������>f��ǃ$�&j��J�'�4k�y�V��vZ-�:�m�m��8u�Ĩ%��ԉGa�uU�����K�d(P�lO`�NR����T�@׌��J|;���mn�YF���ʧ ѩ���Rγ�@�ȝ@(�t��5�p�f��z��{���1+�f�`�y��� ;�b�9|���}w��u/��x�Y2�Ϣ9]D�n�H�I�s�h�k��^O	��J�v.�I
��OB�{B��6�.���1�i7�l�2�	�����[���ⲟ��F�50����榵L�勷#�U`�$��8���.H���A�����>
�x�b�Q��'id��ߏf�7�bf���ߎiq;X����ϙ��2J�$�p�1)�
���l��1��6���������j�q��;�p��%�9�2_��*�$TqGf��s��f�V��
+����}6��9z�;A6�;u�o�Έv�]ы�i٣p��И�f��k�(��!�4"Kwȉ�j�F�����>����՝KM�v��U^l$��y9
e��8���~��}w�f◺��|O{i�>p=0���J��t�/���
>��[L�=�ez1߁�/ܽbkbr�(5��;;��NxQ~��z��'(f�9�
�����2��>��L߶ձ�UO	���vˇ��p��Qے�5�A�~��Z7>��p����?�Jvޘ����͙b4 �,�wӷ1 Ċ{��+����y��m���QD��@���^A���]�q$h�ʮ2����Oz{@��}�z�P]�6�Ec��|�Z�w�*!Z�Ƭ9��Pv�z���vik�fu9�#��E��������R�ы�p��\P��^Cx��:�zW�����~��q�N��=BgG\EK��k�W�u���;�-u�R�e �c��T�`��&{�K�3}	ޣ��:n�'��2�������2��n{�;�s:���L������/�:`��Hg�n�=�u����Lv����ʧ'��e�����i^$˃1l�A�H]L�7�m����X�A��x����[pݠ���z2t��^�SX�;��7��\�Iya@���N�C��\n)���*��D��p8Q96m�7��A`g��&G��A@�{�� }5%0���l���Q�+�Z��T˹C3P��:G���-�8v�x�F3(�)�Q��8�K�&%*�o�2�C21�U3��4*�����uE��1���#�����3�M�n�v�S2)L�j:���G��όp'iV>�������)Nq����}r1��_��>������F@�V�&��Q��.L�Bm]�J��G`*��	�F�d��x9Po�q�����y��[�|�����*�+��UW�*�+�A�T_�EPE�A�Ȫ�+������T_�
�"��EPE�A�UAª��A�4UW�QT_�EPE�A�TUW��T_�UW��(+$�k ��`1[�0
 ��d��H�|p y
��UJ"�)IQ)UT�P��U)
E	DE��*�))�I"%R%HI$��P��P��BEJ%A$R*�RR����%JP�T�UJ"
{V�I)T���R�����R$���$T��R*	T�%U*$J��*� UD%AUD��$�!)B�@PT(V��� �)J���*T%T�UTBE��@����  jsG�+m�6��ٮ�U�ݶ��%u���@�WN�Ұu��G+b���n�R�ET�20AI��ճ��H+F��
�JRP�   ӪT��(��Y��+j�hwF�(ۚ� � �Gwm\Q� 9�k�(�@h���.�GF�(��Ft1�E E�# �  �JH$B��E��-��  �b���`���[��̘v�h
ء�@*HAUUE�*���4iUhaU@�6�٨P��L���
IW�  ��
mUa��Q�0 m��V��^�;Z+�����Z�ӱ������kt�)N�pkr:(S�i��U�a�)B%$��	D����  ���J�����lJ�%gT��l��۪3)�Ф*U��Ҏ�$�l���m��m�d���N���u�9� �1��P*�KX�*Dx  �Aңm6�0�li\�eN�B\ͥ+��0�h:Wv�6��m�����X;aJm9ֶ���@n��Z�4�cD�J�U���  ��(ւU2V�^�(�Sm��[M�����N��Χ]�� K)+m�Aњ[��c��lcN�MuCR�l�u��;��P���!�
�EPD�  b�쮚讍��.��MeV���G[;�݊i��lj��u�Z+7w����uF u��ȦԺm��n�km]ۦ�������Am�$(%E�*�[� vh{a��U��Wm�20
(we�����wr����4U�ҁ&�����PQ��aJ��5��wn��)F�dZ!$��)`�Ѣ�   �+�����P�tҺ�j�¸�:UYm��N�� jQ��t���փ�W[@��ҙ��4��V�kA� j����J*	�4)�IJR   �~�M'�hz� )� ��A�F�"��UT�L��iJz`�IFO��s<�`g��E�I�ЕP*�@�ބ�#x�3�&?o9��k�}��g�!$ I;���$�$�BC��$��BH@�rB���BC���K�b�o߿�����PC���P�[�[���B��8N�H�W��Fa�Nx�𝵳"x�Tı�j���v��G��cUL
QZ�5g.	��Sk^�t���d�sks�1k�
n;��lJq�Ԇᡩ�ǻYV,8�Al�:����X��ݸ�U���&A�+JU��F�1�ԩ�llTE4�U��[m]�蝣�4��e&��iEJ��1���H�i�k6����0l1��;E�Ð)dա�=f�C%C��8�*�F�=�ҁ�R%����B]�nU��ID�!�$ۿ��ޝȪ�mf��*1@,щ�c1�rU��[%���5{�+4
�T�j��P���b;vr�*lV��AGW��ǂ}��؀��[�ͣ��W%� ]](�77�*��b�eE�$̻â+,��5ZX96�!X!�s1�j�˻�^1X,*��0V7�;Y���EL�[ړ�g�m�t���S,�B�96�S���J��[0��;��ں� ,���+p<y����E`���֒������oj�ݣ#[n�b{�;��5�a
x^aÀVFn�Z�F3��Ma8��S0��u���$�v֊�H��B��� -�UZ�b �Hjf�nQ	�K@-䛅�Iz��5>ʴ�N+8�4H.f*QE�M��U�aR�ՕM�
�"-�A7u`������:�������1GZs�e\�P�9Z�`Gj+AEdG�a�v���MhYEk[�+у6��6�Ƅ��!+MX�OP5n�SQJ&�9�<y���k�D�Q|#v�,�5	:I˲�2�ɑ-�Ww�'n'��vK l���I��ઐ��S,��-��i,G(-bb�Y��5�Fh���Z4�����Z�SH��)S��0��˗d�Mu��/���E����r�7Vb���;Wx]{�ah��eշomX(�c�G�/HyJ�m��6�7[S��[Hc.�D���a�h<���TS2��1�c"���^;��2�K�?vIL|h�bk���hYYl��bб5Q��lܱ�qj�"�u��"�Z��i.Nk�X�te����@ҥghfJ�zGٷjB�8�U��鹣P�*t���gsnk4�\�54�`ع
��M��J<�@ꕈ(r`;͉̦Ϊ�f�N��0��Oa�q�kno�[:�ׂ�%���Py�3ř�Ct��+(�=�4K��fX�K(9n���R�@�����3mV]kh�u�p��8���n��� �Y��V2VV%��Tn�4����H(���-tt��)YI0�
`��s4��ʼ̇;\�m�TjWX�o%X��A专Y��)�&��Yga� da���y�d�h+��)4�!a��60m��|貶��Z��w�U��6�@)=���3r\�8DN�l�d�t�%�)�EY�&�*n�����e��,<*
n:��E��&���[�h2�ۙO*�������^J���(X�[+D�	CN�W�a%l�u�dgP$a���,7e�;J^��7ڑ�J�������tf�5�,�+)Ԥ�C�<�T[�m��cpJ�`�k0�im	�4%e���x�nͦ��1�4ǟ�v���U;�ҽ��c쵳f(�U��9����u�H���4����V	��Ml�#!�m�@4�A���i6{hbLe�ݺɔR��^Z�3Z�ь^ �nmX��%�����e	��5��%!lY�vdJ����dL<v2(�9DX�U�2:4��L��飅f�LA�ff=�-Z� 0����*�B�WR�AZ�+q�qec���:�	�v�9p�(]��:'!MS����/(�;AmY;Q]Z�+㽺�I��ec�ʘ첵h�
�!�t���7KsP;yn�1S"`RR��񘚸6��Ƕ���L"�S��i�N��x���	u��6L�{{5�"�VCe��uJY7W36��e�[���y��jeb�P��%u��������­d`�yla�3��D� 4�(o��]�q����:7�V0���]�Yx kEx�0�T!lj�Z�[Vc�&�KkY����^��h�)�.���΋*��#�K~�F��M9�أb@�;+aH��!�`t��^�Ӹ�ff�R���@�;r���w�-���N|�7A*y#��ɏV���Z#xΥD���/.嫡�Tx�İ��9�3��
g���[����!Ǔ�h��(�^*iy+&��ut��9���kb"7�`?��5ʁ�فɄ
{D]��Y*��ijb��D�c���˄�Ѹ�
͐R�^n����dY�Eޱ3Z��D����n�b�I-�ɢv�3sB�Z%b���"��賬%&^� �$�k)��w���W�Ղ�gEf�Be5�5xun�6!aڄf6���޺��` �p�p����j����o ӱͳ�$jJ*�vK٘� ���f,��˙{���A�V�Y���J�_\Q,$ln�
eb��$�n��ܲ(0o)<��h�r����m��̴��ٍGu�����4u�$�n6��3����ZFԺςN��6�nEY��4��m�曬��L��lKgi��Z6%�;�ln[�T�v��d+��O2P�)x ݢj;��Ʌ#��VM����=ZoV���D]�N��e�1��y�����.u�wK:�C�^UMN��ww�m�72ѩc-���#6:�W�i͑�ӗb,���oS�L�H�/Zկ�s�1���YYf"0nGv����8-	�,ˀ�2b����KE���mmi�e0�l��2��ǔViyI\�dY*��n���ח��+��j���� m^�&5YN���o'!�W˼aݺu���-���j	6��;��^r�v4#7^+�)E�/��8E�WJlT�a�h�p�p:X��ڢ�����%v��Sj�Sס��l�I�Y�f�'\
���M��X6��Usul-�o�Y�rV�3,8V�fq��,�R嬤U��;[8,��Ö��f�t�����?���9�8��t�5o(n� v��jRG�M��fM����-[��*�r�U�5/^������Z��)-[��t�T�0�mc�ݡ�f�d�r�-ܮ󍣔�bO@l���*/rO��	D-�kY�7䚳6|�Xnh ������ܔ�*F�u{�;��s+/R�� ��z�k��L�bދ��	��Az�*F�8�Sv��3GΥ
ԅ�P��HT��E䭱iT��%���h(F�S6��4Q9���b����f
x�����%�n4ov/��#V:�ņ����C#@�ҭ�[4���&޷�֦r�%�d�Xv$�da�ś��4���1��1d�Cj���m8�/t7�Z���ؘ�J��J���#��{7���� SN��{��QZL�j+p�bd$����Ui�R�����D(Ջv�T5����Kj�v𛒥���Y��[��{���JEQ�݆��f���-�Siqa��p`�˘�ak#��Yf���\;��jd�[�0�mn���^�Ul\ ����U�`k6��6�����І4�(����k%���g2�kA�j��sc#+aګ��=`�4�{y��֛	�e�ix���$.�c	wL
6��.�*�h�n�D�6N�����CWW4���/t�X�u�r�@�m���r��6��޻4ڸ��+z �-;mɣ.R��`�32�T�)�/�n;��B�b��h��o(�1K�:���B�3i(ݠ.��?)��Z�z���U�����Cv�P`�&PV<�
��?�wtP���N)��ϵZ�r�,�h֣Z���w���t���SD���ٴ�+�Y/f����+K6��Q��d�u��m�-P�[��P�$���8�w��PRԞ��CՓv�_e\�M%3azFک���Mi��Y��OUi�ӕ���F�ˬ-l���КUcV%�f-gBW�a�e�t;L��.����M�U�R*n8v�oU��:9r6w�R����Q�@�F��C��4��F�x�	�jk��UY�ϖo�V��J�S%�۔^]ۢ ���r�m9�-n�����Y�S�51���h`��ꙕ�e�ʺJ�����`���1]: U�R�z�d)��3i�t�jw��j8�]cc�)f��C�;4�4R[�.˳i�t	��p��x[�փl��n���тT`ѡz����f��Q��7��R��!@-�d��4C��Xģ����j^T���On���v��3+U�x��(�s|35#�)k����}�ցJ�*d{�Cv�"V����M)id����z�5����(�e��U��{���+n��Fb����Wu��Tf	��X�����ʬ�)�)�լ̘�f��l�;Ւ\b��)k��*�n 2��i�i"�b�I\�?^ݙt��ز�5x+�VZ�B\ݓ-������Q�ˬ�⧄3���gqStԗz�p�,ݳ��j=�/ڔ4T�`5�ItV��%ދ�Yowi4�16�<8�������&�,L���Tҭ{�+*��,kt=�sX �S�-[�.k��z���7���WR��kX�L�ʗ`�2��C���Sd�z�Հd��8�Jf����^��ִ������6���Q��C3>�n4�-��ؓQu2�{ZVm�I�ۊ��ˢf
8�"#պ�SH1�0fAkc!Ӛ3p$��.��m�1 �U�̣��1X�FnmوY*«�/f [��;il̩Aj���~���N�9���(��1+F�B"��iQ���	��=:���/��+��T[ڳh@�Ԉ�@��� Y31�qf�*1��LS?Yɷ�XNH4�m����j��O��Hb�T¬��#��"��d���
!�� f�d������6T�x3�@\�����.�����xN]r˲𐆕	��Y
;�O9z���:vȵtM+�kNV:�B�U�\Q^�@bT6e�ĢD�A�sVd/p�:�0즍m*U�����{�U`��hu�7��R��		4�M�����ۨ�]�x�WNf��73����
�k�x���S5	-!�{w��f4V금v�,S�����"v�`�֘��/�{.��h� ���"Ci�3�o\���f��I��Z�)&���F�ю� !B�c�g��s5Y����{Y�X6e�S/r0�I�_'�i�k�Z��&����J[Fk65����<�a�K+l���B`q�Z���a-��=A2osv�m�Tm�Y&�)j�qfh�pc�1� x��P�v�z¶����e��%�(�6.�c̴���:Ѳ��Cc��ZKld!34�I�a��q�n!Ah
	���2�b <v6Iwr�ˍm���ԭJ��Wuq鿵��B��y�h�(�sSvf\Rѡq�(������f���I�6���ZV����eb������#��z"�j�=�-�H_f��Y��y]�FC{J<9E���JD�x6�m�A��o@wR���z"h���Ze�O$�Г��$�1v�#4�5�`l��Q�E����
X��vӛ�"{D�-�f�1ә�	[{xU#�`4b�.��N)�2�e�����Cr+�S��kzw(E��鶖q�.��׉�gt�J5{"ɳ���5��gK���-�b�2��V.:b���T�_�3Uj�K���W�J
j�.�� �00��v�dR�X'u:R�<ȢMd����(=���$ٶ�w�0�"�D��U�W���U����a(o�j��k%�L��{9���>bf�Iax�e�
:��.m^Joi�ч.ީ �2m�&M'1�;�#Gs�af!�+2�{ka�CtZ
)ZW������r��%ef�1��}�])cR�AdȰ�VbyVq��T�b٪��$f͙x��i��$��Y�B�jL�!�e�on^�A6y-d��� �ؼ75B�$ŦK`�N�ZLjO-f���.ZS�5V�J�n-ƒQ� �W��S6n�1��÷DPӘ-끬wBi28��m��U�wj)Z���t��t��P�_� ����ͭ{��/�X�l��%�yV�I�@�:+[;�T��
�s-T(^���7.��k]�/-����[Vv�1x�&Dl��[�!�f�֫X�\�E�p2/+��4��2y X�*�l�O7i�yS7j
�!]+3
�<9�բ�e8��+-��!�(Ł���j��Y v��%�b7kuդvä�[�N�Q3sr�٘B��kQj�j��[Xs4V-ߺ5u5���񼙐3y]����.��S▅�s&|�!	�LҠ��l0�bd�k��GD�G`���N�Pi	Wtu¢��J��� ����j5C��%k�+�)k:&葹����h�L5��J�"`����EЦh�@�.�T�Gw�Mnlkl	W.|o�4�����r1��-E�n	�xج�x	�n�6��;�7Hz��*��v�2��X����U�D-�&�Vt
%-K�7R��L��
�kofe�x�Eo#�U�H6ˏ����QBf�K
�X�ʶ�Q3���RS�������Q��
��6�R� r�3�Q�-+�s.Gaa-]���d;v��4I)�sm�q��V0��g-2�PÔ�9R"���ޝ7K�ٍ�b�	�4�E�c4�M�K�/n�=�K8�X�f�%Z��j�O`�yy@�p��ԡX�b̒�'�^�ͫ�B6�Q���R�f��ӛ�v��J<J������ݖ����{�)ò�ά��բ�����Xw\B����g5ܲ���O��2;���;�bϟt����/�A�)��j �v"�����e�f�C]��G̬�ˏ�X�X)*N�AhOtT��POW.a]��yS5g �}7V��Dfۤܡr�;vx�9�D,\�;:�yHb���}-���'2�sjS�;kY9� ����s�s1��u9��T���α�;��DV�c6���1ZN�����%wQ}W��wwrY�Qe2�؄1�-�b׫Keq��\ջ-��&YBc�2\��4��D�򂋄�CeT�)Ɩvr�ݷ|e���E�Հ�\�����W��� �BF-ma�Yd���#���� ����-*�}����Jae�ֲx��EK��48�u´a�+&�T����%gP�D��k'�7�$��^��[8r�׬�Q�7,�/skE�j�f��������T^uf'�n�jo���¶���eq�[�k��=GV�{*e�}�텫9�55���o�=�L�_d¾ե	S�}�����W-.#��՝}���Wz؝���̜rD�js����:kw~Z�S`̂����e]���E��>�Rc��w�9].�;,��ޢ�D����K�C	b|�i�I���~�m���$�> d�2D��J���<�ԍK��ũn^c<��[-�����Wj�w>��{Q��^����n,��Vz�m�ٚ�.���:ܙ�5�OT�0�}O0��f- &��-jn�lK#w�k(�L�t�AqP���!��gv0��9Tx��G�eRc�E��sY�e�����_hڽ�a�����a�;;Q�3[����P�t�"�sI�Cz޴��
t�u�^��<�t)2��}���gQ�n���ڙҺ��uci�D����q[b�45�O�<Υ����b�!�Y���:�|yP������ajZ�zz;�x������Qfaǅj������x��M^�L�b]���2Za�[���w�8��l�l]]˚�6v���M��<�Ru:���\�
���^�"Y��k {&�ʒ姎K|��Q{�:����闚��2���=̡7
b����u��iR���
`�1��塖v�s#�y7RW��78^�]S	�5^b� �,�u�2�*(Wrj�LB��x���9c�r�v�v</o2����]��m�r��Oq:u����0���1���p��{�&��rt+
V�u�gSlJ�����ws��+#<1�}۟9�)�k���5�ϼ�m���v|�@ȍ�)���U-��wN�t��L�f�NsO��������'�I��ݬ�ŖF��nSQ�Q{�D�����%{�a׆��f�w�����UϝJ�PU�shw�oC�:m<^�X��f��������f�mM6��P�[�	�s�$hU��,m��Wq�*2w�FS�y}�̴��ZS+��v ��a|���Е�Zrd��ۇft���y|�\Km�Ӓ�j�K2�u���V�X3�Q����o�.�q�t���A:�V�L©�7�:�S���QN��V�Y��w�v���e�<g�:Ȟ ��0_�����;�:�2���L�k	��į�N�k{U-��n�F]WQx��݃�:���y�}����{��j�U=��D!Du���\��]n	Ax�ލ9$���C�@vA�Y�cݼ��싙�c]v�5�.ӻbu]�`�L���N4��k�kʽ�i{r�;5aQ�j�Ran����N�O�5��W������m-F���z�8���_,[��ub�i��uC["QE�c�W]VfT�����
�9�rEI� �R�4�*�[��̸���]�.
�.�"^[��b�I)��o����P�
��o�p���L�fsњ��wY��\��˔o-E�U�Q��9[�Ga��tØ�^(J3Ep��|�{i�����z���{)�-���ޙ��J �:����Π͊���0ur)�u
�.�y��z�e8�p$�=�`M�ŏ�b�uv���`�yo;��#�n��o[Wkbv�:u�ٝJw��˱�s�нQ*�UK���mD9��@
�Kz��ӣi�jOʑ]�9:x��ߐ���HvtUuڵ�:A��_p����o.��V��T�7F[gd�u��Sw8m��5��4 mh/p���f�+S�r��G!yg�àZ�+�3�.�I���=�u�Ii���s�uj=�g\�u��q�U��v�#L��#o��1X��ᰆ;qvtPffCr��G�]�����J��mPK��=.��w}v�zt��cޭ0e:I�bQ�4e�Ϙ�|/S8���WoH������e�̣� �>w�\Zn��b-�n]�p����Z��4/_u�ٝ�B�9��˩�:Öw>c�J77Z�Re��ht��]���rՈ�]YKdK�@#T�x#�
ה�w|���U���ޚ��q$Nα���f�I��=u�Eˉ�H�/6]��ٖ9q��3��V.X��N�ș	��+0Հ�r��ۤ�tY��ާ�0�uc�6_h����� ��FP��MG0�a�(��i���뿯`b��^C�J�.�&}�9(�[k�tdlk�U7T��w�b���2=�*� O=���u>6J�����T�|5!`Ӷ��Pn��qɧ�*�e�K��B�Ѷ齵og F�[��vU %onf��[�+bBya�Y�.�����v�%n^P��5M,}�W]O6;	���m�ثGvȴ8��z��8�c< �8�1�b�ն����!�)0.뻱�@e�奝<A<Μ��:S-��1�ݺS1���mR���ଷ[OB�&o�C�n��W�CGM�]*�]qFQf�}��iԐ�AdU{�Ɗh��np����z�bB�W�q915ꙋ;ki��l�h���6�����K 
����&45����t�ٙAf�	s5ո��}[�A���&Z����e@�`��[93�wͧ2q�]qմ�R�7��,mv>��2�aȃ�ǥ��[n�������md�k_Nq��[�6��˦�d$p�+�y\fk%Z�c��k<�/I�;��e��Oe�M�9W��e�1��p*F��b�Su�k�5ޭ� 8$pT���4~�x�ݙ���9�t�8�=@}9T�[�:�oc�q���S�4JJmwi��8Zƻ�9��w�S���\�m�:C�*����% ��m�3�e賀��nW��<��q'��¶�x'5a҄�U1q�y�v��Z���U�ehć��&y>:�*{�����WT�o�$
�ZRX��k-ee����j�
	֓���3�C��Wk�͊㝕'o^q*�v�K�z���v�L��r�$��,��4�q��e�v�U�毤��g+��#r�\ ��������z;�;�n�����(����ѥĲ_EvOp�J�<��:�>y�IP}a�������n��	9�W������)żs�ngϺs��\h/G1�v�� չG-�8+8Z4ZyB/��&+s�BwZ8:�s7��(+���(��I��3���JO_.лQ��8��-��]���x��2|�F�\ ���p��9������]�v��Œ���6ܔ�Vp�R��%��c�Ek�\��0���}F�qY�+k;^�2��x��+�Ubmwk�}\�i�:�N�!���c�M�J���(�����FF
�x!\i<̃����	��VZύ���\���ܭ�Qw:RI�;���Wr���L��Jɑ���nb�h#]"n�Xa͊��7��R̂�'y��Ύg�����Yn��;�7�V>f݉E��� L���m̃uZ�N�m<���$] G^p�(Q�F�r<�]��Ә�)9����P\'ƶn��T�9�E�Tx��d��e`��8��l�7�N��/�5\�sD%�%�،�t��o,��*���.6�bj���z��蕃�ꮮ5|�f��ɯ�J�1��V����0Kw��P����#���Y�9�\2c�� q96�=�L��h���Q�םP���u���2[:��iZl-��;�k:Z����ʾ��Cz�unn�O��X%R�-��t��X�N�ۓkfM�vd� ��W:��	��VnT=e����#GZ�������3M��[p%��w+��Y
�����P��\���9�7,Q�w��(����S����3qڭ��������=U"�{�c�� !�h[�6V5�<��K�70�����X4xu61�s���g!Ә���O9�����YE`�Gu-Uc �x=�E��VuA=�M�)gEtE�t7�5P�z���5�;+�_+[���]J1w��j��� �R`�f�{����jԶ+CkRt'[�����5\TyMa�����i�gV+�'r]�[[@�����6���r|A8疫 ^/Wr��X}�,�9S*����sqt���`s�XÝ
{iܜ�򬽵�/(lq��<k"|���G�� ������kA$=չa�i�oF��_βj�M�Sm-�:���"`��u�_n.��0My�LӃbA�	�R����2�����/�:y�����Gs�)�Z&�δ��mo{v	yɦ;���/����k��ϰ5���ȥܲ�H'|�Tʸ7�A��C��V��GM]�{ר%(�4��ъ�z�uu.�e�	���-�Y��l��3�����F�iZ7{ͣ`�{d*`ϯ.���:u��mse<jU�#n˭wW�&�U�R�͢�E;�ԫ�Xq�)��yO�����)��)܄a�5[�cnZ��ɕ�@��+n[ж��t�tw���ün�1ֻ8;+�R�̂F+��#K�����r�5V�,%�-V�����N�u2���] �YH���u������e��rq�ѽ!S����N-��*y���^
O�V�-�	�X���Y-�B[kS�Gu.l�6-[��'{���l���_^5d��3c(���T6��|Ұ� %^�y/6��R�:�2���Ly��.oKں<����M�
���/k۵��p����ҕ/�N�mm֌8g�"�40�^�K\�.�<"���b�1���#خG�2º�8�����{��ߧl[����#�H�6�>��l�P���{fsz� �����fn1�.d:�wrV��G|�!�v��f�yCS���l�V�J������9��Z�&�/~.�{��3)ꫝ��Ujw~�~�O��嬫�6;��jǍ�V��^]^s�I��ϗ*�l���V�\�%#��_h�ag�s�l3�j�M��Ǝ>�j#�vȘm��L�o4����Ὑ�3�Drٜ���{��J��V)w�)ɛ�.�٫:I��k�t՚�j	���9�
��F��8�b���\���7K�Jȏ%r�W7������5J.X�Es�[����o�y���!]� f>e�U'6�nmEID�����t�/s�7�'�7g4K��.���]N
>Z,X��(�Ql"��7�C��:�4��g5%�5�U��F��J�xy�B�G��`�g�h<��b쨆x;kk��v���v�(D�oo[7�8���%�۶�b�H��f�ķt�{,#`KQ�ho��!��q�M�u�Cvw���&������z�R�M��Z!{7�,��,^�{�ܝۛO�-%�����o?�5��n�j�*{���8坖�񔷺�K����1-�,���tB�Ң�,4��ݧR�2O�:�q�$4r5ׂ[��5�ӇS�T�/�0-8�JD�#!\h��TWz���t7~vDksn+����c85v��E��̦�@F�������7U�6�O��|}j��Y[O%���=MM����Ufl�3�B'+ ���c씴��{\���[a��4n�p� =`Q�7��-�u[�x��-}���'0~4�hwq�f�xf��;��\U�H򤡀@��xh���3�WM�&V�����zFnт�#[$;�>��-\"b��r�p�q�9	DX�6tX�\�nn��NY��V�D�yK��򷭄��,_!�ܛs�<HuCWk�iaξ�uԓD0�`MW9��R�gN�5���Ф�ӝ:�BG�#O��Q���++���W��I�&�9L�O/�"w�>��k�ܮVhm�A1D��Ig��+���>*z^���^�� �׭��,��j���t6m1Oy�h��]����@m�!|�h�Q^�4�u� ��<C�vk�T�*ᗬ�X���+5b�t}{��j�L,�J:�]Z9�m��`p�s����/,��L�J���m,��|�1}�.�{�wIlom��j�j\��]m=lU�K	�ѽ��ܟ(��M�̝�T
����
�zI��}���G��䏀�Ld짵j�P���*�XG���Φv>��,��8;6���@�֫�Ǯ���p��E�X婋���x����m��eTwz�]���S�Ȏ��Y4��_Z�C�c[}��ғdk�w	�u��>�zo
J�b5���:F;B�:+�ulm���s����qV0k���pV2xi�ݬZ
��T��*�w��P;��v:��1�����������@�ec�o�Z[N:��eh�VD�Z:��i䞕բ��ڼJr&��tMż8�e�(�
�ƍ�|i�s;�L���$����]Z!��y�AU�K�oklU��7d���Jom��5����K�=YjQ2�]�����R���Y*3�rq�͢��f[�i���T&־��RX��Z����6�(����b����k��`�rK����'7jWOXKpt���vj�V�I�:����Wp�v�W�g9�����ﾯ�I�!$ I)	!Iߵ�y�{�����k�>e_���0,��=j�iuys���凪n1Y��s�H��;���:���f�z3�,ԣ�L�:=0�U�i����vf��x�7}H0�B��Q�	U�}Ԅ�3;��P�g+M�Sʇ�L�2Қ�&�v�()\�	�w"⮙����5�R�{x��.c^>��*NX�1v�9̮[;iWx0W�w�1ʒZ�`��s���k�N��*���a�ͽ��N�Z{�����\뵍U�C������G}0�ȴq�7q�!�q��hz>Gk3^qiu����7;�P�������]�RjL�Wy��$F�U�!��t^h���1���%���ݧI���X0Q���eu-k;��M��Q�	`�U�
1�kg�|�/��\���3�"��@l��eY���Q�݄���l��Q��9��-7�_�ZB�[���X:�;�]��JI�Es��sD}]�a�3%]��-�G����V��R��dQo�\��#U;x���@�(��Uɮao�	���8��hh��OA ��os��Qػ6Յ�6�ms��yW�L��m���oc?e9{ �#����ˡ������1:���b�2�.�ZZn�3�D��xoq���h����(+�<�hբ������J��̉|�{���\PWh���س�3ʘ�lW��1.���ί�wn-̳ƒ���M���=�3x�h�����(+�2����̝�YҖhY6nW`�o�ͨ&��<���!ʑ)��9p�`�3!9�Sitq�Y�� P���[�R��N�9)�G,� ��0�^�s�Y6"�*s(�h�P����6���S��}�l�VZ���W!�ڱ�P��h��໺�$�Έ!�}���r�U�oP�@�V���0(�V�7�M�>ZO*��_Ex���$�ӯ[2�ά:�J'�ƞ�F�xͣ%�lG0YCrW��%�_�t&Kd��z��2I�Y|²�3��$�1�Te��'s��F@��d��V��e�x��rVo#|nr��٢�bF9�hp�ejHu�d5n�4�� q�wC,3��t�N>f���y��f��
�y��hh��Ko�n��y=����|b��:�w�3��M�
���OwM:�31�x�y�1IbAX��=)v`ө7e�-��;:4�Lٹ>����⁢��I�F��Z�8cM��e�J)l�}ؙַ�9h}�6��]������S=�s��Ε��F̓�˶J�E���kv�VeѼX
Gj�<lgN|J2���+G�T�&�cR;�x�:�y&w!z�FV*��K��HA��|:v�ţ.�Ҡ�xp��z�H�v�n�#)r%Bx�`�ML�lZu齁\/x+���F*6c��!������d v�8����R�]R�"����ڰ�A�cwt��RYV�^�q��f���G���
	�Rf�N�1�W�@�� h퇝*�ۃ�(��s�����NX/�
�ĸm%����Q�t3U�T��Lt��m>ރ`wn�Y��د*�gn�] �7c�f�
9���J���<VK%��3j]�	�3U\�d��ӽCL��:�j�6�%n)S�e]�[�gM�J�,ē���\�cޜ�C ���S{�V��N|�"�]��
zx�M�W��J%S�J��z�C�����R����D�5]�h���#����'ZZjĵ�r\�t����@%uҤ�IX�q<�}Mws��=��(p-U���:��
�ڷ�U��X��s-'�{��D�S�ȇ�&r���v�"	�쥛��Q�[zy���҈ Mb��ɖ�pK]�0�m�]N)\!Z��:#��e�#�ee�ީu���ǁ�c��87ki�`��k�K@y�����P��������y�6���������c�Ⱥ�z�9��)���7��	
"Jx��bֲ���V��b���:�O{��Z9�u0�զ�� j���j���=�����Ћk]�N]����gQ�ڟ�6�ͱ�1�5Y4��1T�
Ar���Y��[����N7D*���^�C����>4��kp�޲`��,N������(<Z��un�)_YԦk���Ki�М<r<�]sז����l:���o��@��+x*UȲ����;n����*U�񚦾:�a�9�6^�-��Mr)�v;۸u��]ͦ�4�����r�o}md�*��PO��6mKY۳_�Si�5��K]S+����Þ�#]63ӻ�+ǃ(҆����,]x��	m�����3Y�&�-�0�to+�P}�7ƻ; ȵ+����T-�,��W���2�u�u�O#��c� +�Ƕr,s2�J�/x��y��P��(<�g��NK�콍;.[�Xŕ0��V8S	�^c���M
�.-�6ŅQK��ar�W�ӕ�
/��qM�����;u*97� �_:!�ClY��>��et�	�<;~�˦�������3�>���)c�l�dTX��4�q�H��>����o�ɴ��ݖ�؈P�.=�U��zR�ܝ`c��K!��F�r��5۾�:��K��j#�H�6���r�����Pj���eM��F�T9}-��0��)�5kCĻ�Sꈛ�������rQ'�ǻզ����џ,ܦ����u�W�L�g(a�X�ć�R�;&��`I�ԸB��h�w�+ Пf0�F���d��WbT�aI�@�\eP���6w9���^pw+��yNVi�lN9ל͎�
�qs]����X$U+.�s�s*r�I/�[���h�^P�P*�X>�w��� ���ᘦ	m;�vޱ��M������׵�+��[�@w:Wp%"�u����wp��s��uϥt��CSu�nk���Uw���W<������$����r=�%]v��F�����n�6�6������B�0_q��e��bu�����p�瀤+��'�D���c���ռ\̚ݣS�0�u�g�lW:�V�e�a�Hc!��靤r�Yӏ;�[��C��n�ъ�[k#�9�t��4ovr��"YNװ�Ģ>��F�;"ot���+o��;��@��La��>"KT����7Yۥ�ۇ4qj�3.�_%��$ِa<���VL���jltu
6XV�&�U�����</�#k�T����U��E9E��08�T��{*G���,U��!s�t��Q���{��1�(.ڙ�hp�'-C�o��C�@�;'���p^s�]Y�<(^4�e^�5�U�wi����S���$���u�b�U�	̠8t�oy�������,.{�)S��@䔤��]�9g�7l���Ұ"�+��7z����<�m���@k��S�����B�V��x��d}�+Aqb$��j��v1�v��*]��zT3d�YB� � �MӠ�FXв��<�d�F�ӷ��c4��JJL��T��M�]C1kԬS�P����umfӤ�x����k�@o�2*��
�+��4���$�u�KyK1]gw\Ǖ�]w)��sڭ�'voZ�׊,�:�K��׽ֵiz3�{����їW�f&Е3�q���J9�w1/��l�.޶4!0��(g7�Vr�D�]�Y����۫;[`+���d����ֵݣÌ=7s�H�ͱ�"�ǻ%)���1�V�rE��ˊ������,.�L��p��\[��S�P_M�$�u�ד��E�z�qW�m�c#��Y�p��&��� ������v5�ٗ�Vs��Jx�O�e�X�����6�� �l�tUA]��{�u!��Ƌ��kB����ܴ\�>5��w�����e��3����H���$v\T�^^d�He�<�Mv�r�7�7����� 2��(|�3[]]�R��twu^��N!<�i-���$�(�L�c�U�#���m�i�fŴ�t��l��G>{W��-�c>(ۄ�:�&[�dK���.E�q���b�j�,����G5�doc������U5��wwʠ�ooXV=i;lOI���H�ܘ��m��n��v���Vw��H���r>�*k�]0�ڇoe�k��rW�tլ0�p��0��F�b��oVpYh ��Չ|��u�:+w-�-C[Nj�įD�h�U�b��LT5�Y���䶅C�6T�b`�M�NgiZc�j�Ƙ����U�s��W�ܬn��<to;L�WM����/��%���lB��u�J�pB=
�^��i�����Z�)<�Cc}t���:ְ��	�fΕ��t���D�'-��`���c0
7�������,31�bj�q�a��f벒b�m�Czt"�m�^�����#qV�Z@�ٿvIwSH!q35I(�,�B�5�d��̓��e��Rl����j#�'w"���Iѥ�9�M������VX�o��i��}�m4��*Fy@�o���0b�ĎrbAAt��XX�ppq�Ke�:#���'$[B	�6Z��E�Ǯ�2�5|0-��M��"y��]|��9ɋWL�s�f�J���$�5c&Z��cT�$T�"�֝��jV�k+�c���>���J{N#'T�;#�2�O�E��FV�=�+���kٰ�l �9dT���R��8�-Y��/r��qY�u,��;R�2AE�{���d��Wf����Ow1]����Lv\c�%��}+�XƂN�r���$�N�U��)xZ�����[� A�]-*g����h�(�l�\����l���%̭���R��{X�wb����˕�'є�)�vz�Sɡ�4^b�>Y����$��s:k���}7�����K+;
\z�][�٠ӍL.�=u����P9:�
g�_K���yJ�ò��	��c�>���{�/�9���tK��L3��n�ӭƪ4��z��*�����n�3KWe�.��:�d�c�{�ȍr>X�IWD�U���r�;Hѳ[�N�KӅ�\�w�5�Z�V!�]`B�cUd�\R�J�y}˺��|7�
��[Ζ���̾\�7NQ�ɝ[�$��P�+����5:Jhw]B���#"tEZ9:�)�04�I9� Q˾eR�����y��V�:��{����bn�4����Pn�|.Wb]���e����͐7�Sy�yл�5"4�4��}���Ⱦ�Ҷ�.��}�h�0�]g��k��%�F r�My�\�y��w[�.�طV�<2}�"�[O9hnj�ˮ���YCKCL&Q��'�Y�n=㳺�Z��T�w�"�>Δ��T��۹څ���*U1n�\�6@�p��r���q�}�������o�]�)���E���э\�je6�u��5��V�LhV�U-�R�Ý�Tkvs�ʳ�Ծ��k��|������ɰD6aw�VZ)L�65��|�f�*�h<��62W�͎�J���*:���15��՛��om���'�ݝ�&��� �ޕ*�W:�����2k�����Τpw��mʟ>Kd�V;_KR�2����u�e^Oi��֊���db�:�^�5u*�:J��}4V�Ք+^֍4�݃#|�i6�"�������Ȍ{���N��n���t�pD��q����Rbq�Ginc�O�=r	���E-f�]Xi��5��(ڷh���%��3~�!�	�[ͨ,�3U�]1�y��I�A+�04�����%��Z	���h��G>�J�ox�sdm!�<���+���_I�1J� � �9�m��8rT��U�U���!�4�w����ȫ�o�S�ph��Җ����w �nW.n5��T��V�;�o��R�J�[K.�sYbR�ٷV;�Us\չ���>=�WV���0IM6W=�q� ��b�]b^p�պLSSu૷'+��
�WR��g�M�������.9V�� 9)����t�Ȫ�[��R�ɗs��>Y����c��řv
��z��.F�L�9�ϯ7�t�zS���R�0��M�
.����I婼�f������Vg�N��',��.=T�7�N�K���z��UAV���9�$�ދ9��k��;���:#��1�{+[	�R;�V1�4a�������4d��ұjv��Y�����k��y�k�m�/pbtS��������ٶW*Ŋ�[s"��f��И��\f�cn�ކ�=�����p�1QN�Ṭ��2GJx2��ū)��u2�$�-7����	=�ݰ�d�j���T�޾Kn���TY�5Lۘ�F��K9m���`�n(gsy�hd� S�
���%Νh�pFWf�|���VҀ�x�"����?|Rd��m��m�u	�]	����'j�0���l�@뻆�B�A��=�f���@�CW��bX���e�7�pu�^wYb��,=��S�B:�B��N^v�g�.w��d�mI��uoc�ˠ+y����շ/1����1�Xc)�&9V>�$E-}�	LF.���,����fwV�u�;��&�y%9�r��{9v��jJ��y��?���pQ�w�gH�u��2>O��݊	��v�V�ض
���� j;8n��ֺX���*-���W(/��w��%QZ�z�����X����� ��ea���wZW�#�G4��v�揱��kRS����Vr�:<q �]!�k8��Z�a�u����-�J������:�޼η���nS�÷��u�Ot��*�]�G�J�٥���+h��>ǀI� ���K#6�n��vؕ���ʋ��wn����7��M�np"�Lʘ�2�<x�n�|���CwZjG�.�أJ��Z���E`cP�B�lW���s�������됷�2ČMgL�WG:�b2��H��s�!f'13`	���Y���ީP�y5����ﾯ�>����N�E�rR��5m��.$����D����bZ$����p�İ�܇�y�Ad;��o6=�͑�ӡ]��n]��Z�m-5
�m�Ee0Ĵ��S��9���EK͊���V^\��è���o�@�Z�U� T%g�kM�y"��b�I�Q'�Q�b-���:#0�)n��é�R��*uum<yԗH��/:�K��2
y�Ul�v0E�N�MFn���N�,���Z��d�Gc�ud�U�9��a�9����ӥ!MwA�bvuZ���j�ӫp�&gY.�	�(���[��`M��8lp-E������L���Z�2բ��7�+a]��em����]��I��SN�F۽}�ɇ�͉����f�^���Ի"��w����F��M���je�+�ͭy���ZݸoIn�N|/H�3B��h[�67t��P4��I��[[R�7%����(d����� �v����������[4�Y)�յ�p�m ���K�]��v����r��C,�z)毐q=�mmw�B�Y(s�)^�X��y���j���b�H�����v��PוtU�0�7(j���bzOMMQ·Rs]̤+	y9v0lvw,��oiL\v�;ZYK�JK��J�wkmVfp[�ꜩR�q��QދV��g6�jSF�Rr�c�4A��x�����~]E���#�4�c����QDQ��
�����ڨ�m*�+QJ�("��ŬU+R���V(�Jň�
-j �UE���R���m���Ŭ���b"%��*���lQb�R�Ab��X�-�,X�X�T�V[QQ)E�ieh�#���TkX�1UeUQb�,V[Qb�Jʌ�EQUUX�T,J�PETDF+
�UkU��+m"�*(1UZ�#j��e-�RŴ����,��
��[FjE�c"´�����JQ�+EX�1�PU+m�Vұ-�mV����Z��V�6�V(��m����Т�j,���b�J��0QX���TKh�Ҫ ��E�*"�@�1V(��AX�EAQQ�����X�DX�KT�Um*-�Ec-���lEUF�!P��TDb�B�0H�--��V�U�U���c5�EE�}�c���ֺK�w�m@	��_Ö}���ɕ�۔�͹t�������Q����ܺ�ӻ��v	�w����I�Ubu;�r=6]��%�7�K7]k��'ϓ�*ױ���@�<5��z��X�ѽ�9r�w��S�
yp����|���j�L%����g �>��ՙi>��Wi�Sֽ�Y��.����B}E�g������*�������ؕDB�Tú���΍�e��'����-��n �:�.n�������%l2�B�q=��FLmM�!p�c� ����ޝd/|XBŀ�u�k2�j���fd�E�7]�`�5,\�Z�+��W��geʹ�~�cXt�����ɏ�*���
�2�.��Hf�^��>���fs6���\#��������p<-��X��Z�$v���x��\| �eM����L����OS�Tт���Gò�d�D{Cی�����Ҿ}�8z#
g�$�鷙�6��w���k�O���)G�^XLm=�D�r٘�þ�;P�=%��sju�<e�j'��'u�y0��{֧ԥ�.�����fT�S-1���ѭ9�Z�ͫ[��D�=��U6��I���XX[�u'��
y�	�[�O\Տ_i��n��>��Ɩ'YH��R��w�K8�ɹN��85���8��,t�C�T�+F8��B��W=��/����w���#��.�N�ۼճ9w%VέyM��4�n)��,l��<����.VZ:l(j��mL�q1C�3���Q`��a��T;�M��Lº��,���l�YJ'�Y�*u,�S`�Tʍ���G�\���$��>�%���[�Y���y�{�D���ݭV��b���@�7�۷��G,�XZT�O.B���޾�Ať�s��kؼ"��H�͚
��>��:�u�̯�D-/E�Lܷ/�l�ډK�di/*��t�,Ƭ�������`8t�@f�m뺬��E���zvz�bR�jx(T=}�C�e��|:K̻�̩k�7�˨|-�$0f�Y��ժw\g�р�$ 3i2��I��T-��r)ȵlt�(�� �+�����KRʭ;Ot��ތf�C���^�dm�Y�������Pu��&o�"E�����<����'n���4��d�����~�ѳ�Z���817��In��
Ü"������SǓ|�
�qP9A��V5�x�r��wıMD�P���-#�g��R����[��X�"ڕc�\)�[;B,pe_ZbQ�|�j��KJ�<6-�p�Qn��[�h|	�|V�GEW��PL�uw��vm.�pB�onk�ȟ�+��-��l�s*�b�1�if�g�uoQ6�2�-�]ݚj;�QM���Gb�M�:dў��yq���gs	V<�E�2ޕ僳�Lo�ytJ$#�<=[�\�����в����m��z���Xg⳥�v�����{����m�?�]�Òr�yf��3V^}U�J�,2+�ݰs�ؠ϶>����c�{'k�S�o���dS_vb�[�|�X�aXuz�}>K�	�!��h0o:�Q`�qm߰b�z�O���7^�ݯ8�u�P�:�#6��7��,���>$�����x�}\`:�ʘ9wp�Oz��*t��:��\���4=ɛh;@ꯒ�R,�e�ԫ�@�DQ��脫�}�m{}�{OO�]Ƒ�b��Ͻ(�oӼ�D9�,lܲa�����3i�
V^ixf����9�%�]�rO'��9{���Ǟ��?e���mW/qVP�����mB�=�}�J�ט�5�B�	��)�]�(s����;w5x)��RƑbN~F��^�@�Әp��������w"o|����C�"M|G� ���q�Ϛ�(���^y������U���?m��"=.�6���k�Ø(����/��3�W�Ů�S�� �Ի��n�E����b R
�ػ���maN*����Z�u(9�(��#������zy�DO71J���2����%�+��V̽�Op@��e�׽u��mgS}�֣uػ<1�8s邡�0�5ғJ�J�!��C|_�Z�lR��Y�S���]N��0�U�v��(�ђX��	������ґ~YR��I���6�6�ӎ�͍E�M8喰�J����y�D��;%/+���x;֒f�)�ő(S��~�2��}Oqἂ�3Y���C����zU�\�Qf4K�q%�҉���b\&�h��lf��=l�h@�JƇ��->���<�{^�=�t�uG|��p�OR��(���\��c�~�c�]y�m;f�;����9�k�i�I�]k^B:��	�����j�bEsZ��S�y�F���<�n��{�X�̌:�����(O��׵�A��*T��)g�ꩽC�-��q�^}Mn�ו�n(�6YS�iѢ�iW�;%�v9�ޛ�;;3i��O�i�;��9[L���~.\�胉�|�%(ϋ���6Ϥ�sk��X�h����}6�qPz�;�tH�zjD����s�O�=�z�O�`��P���;ۋ�R���,��Wj�Eԗ��-ݏz#�QkG�&_a�5�mp3yEG�V�:����l�K���X�X�;�˂f��ݽ��+������v����.��V���$����v��W:�SI*�gG�8�q�<M����h��E�K��Va��T7�]�x�ƚV��3|�&\��0�{}��t��еґ*�R��}]{��}��`�����
��:�7��7���� �5yQ�n9�W�v� ��G|�XîXC��v:��B��q]x��n�y�.�3/���%���/���u:/���Ϭ!Ҿ�����B^Þ��b����ȍz�r�Ӵۙ��d���.X~vB�k<it�y/+֏��x��}��f��盪�e��·��bw+�~r_	S�&����x��c��u7�S|����%ٹ��_WJ��j\������{���r��W��};WT��a>�+�7�cꎻٸ��-�����RS����޾��]�/2[����J`�%��fا������g���wmzv`��:kW%I]Q�����=1�h��_a�}��Z���+}�?��m�*�4���+or5�v�Z/{�)3W�P�G�{K�ű\u�x[�ڶ�ܖvK��{xЕ��@�lZzx���yE�UF�1�_b��u�M�Fi�Zl3�n�y���F�����t�C\��x�#�5���w��blmΖ�on����x���[��N������3b{�N7u��>��߇/Oc�bb�D��������ɭtq>�F��o���y����������8�Bl䨟��B�g�-�����LX�k�>�r�u/�G��#���
�x>aJ�}�RiO��=J^u�	ƅ��d�ٿ7,':g��ꕻe���[�7��}y�W���b��\�:�P�p��!���=yo��ٻJ�v�^�q���y��6u�|h�(���u+���/&���w�aj{��)��3Xs靮��~��	gh:;@�b�����kfվJ��|$ȟ^r_gY^��=�=�k�����x��	fT�f����2}]�һn��V<��+��(Λ����t��o��}x&u�x�^�]�������~��"{��ZhnBߙ��Mx��K�	%�H��e�c<�=��3ւ� �����;ٔJ��]1�H��E�Q��ʲͫ�Q�us�FPYy�.�!=q��'����(՝�mN��g9�^(4���. w�E�U�hj��U�A+274�U{g���ޜ�؂e# �6�
�ܝD�fMeܝ�����O7���V������}��=w����.޺�6:ܩ��6�b�[se����XOe]k��n?�/�z?h=�8�k�ޙ�h����vŸ�3��>�o�D��;�$z�,k,��#/j�����|;�5���n1`9�NFv�u:ͽ��O8N�m�]����_fx��%Cʵ��>>��W��/���׹7��+�V�кcv2/?A����+w��;��yV�������b}���=�*�)������>>��u����{�n��v񫎇a�,��3m�N_�l�)������kʝ��F��\��a��4ϔ�~6��c�.��B��*��7���>M��[�`q���\��߲;δ9 �;��*32��绖��♃x�61�Q΁Ǜ�N>���w�|d<�kh<���A`�l�ƱF��t�I��v;^��w�8	YU	;3���Z��Au�P��ka��ȗ1�zU�[�γ!��{ս���B��xռ����E�+x����*�����L<rգ�ü�i	�n�s(T�S2�2m.��]S���uGoz�ן���J�6��{>��y5�ON%���[_v[\��.S�&z��M�V�?q��=ۓ&�3܍_.�T�C�����t׽�4�&S�4׽�M��;6�C�_�O!ί��]=�������N:k7ޑf�}�	�Ż�ïz�`����\��r�8�����|�]	C��rJ�<o�%���8���MF9}yr]�a�vJ��t꿩��yz#�XFL���˹}����g�\y�U�p/�m���V��^�=����Y��̮�y��޸ߛ����p�$=���w�K#���{GvW�<��\�J�ɟV�e�ށݳ0oDhy�h7���d�Wc�,���xN��_N6T����w�����zWO;ߟz�{��)x{���!�2>�J��>$�z=�=Y�[�{�J2����>U%�u��lg�y��;uP�3Q���W���t�X��)u廳�|\ w1�<s�.��׬V��\RjF� [yF�Rr��0�]7Sǰ>���ގYp�j]�;�:0i��	!��gb�i��s���9�u�D�s\:��6'T`�]���M�8$��M���)��:�#�Q�ͪ��ߦ�jV��-���~��c�q�Y�&�ѻ\�u��nZr��2�����n���4�z]��C��ɾk�����,�d^��}���r�r���=�?XVew~��Xx�l��OW/dS��Hh[fC��-���:ol�Oh�����ٕ���}��_��>�������l�zd����lϋ���^v/�arUt�y��g�1��{�������u6ly����%Nz��S�������y���z�y;1��ĳ���u�C��vT����7�.]����v��<�q3�'X�痓#�˝v��x�_.}`!�H<w�"S��zԬh���=ϋy����3e���2]�0:��g����q���H��빨���eԭ�7�]�������w+�C��g��ؘ%���,���<���n�)tz�L����� ��Qs��HϷ��?d���#�y��z,�;o&FYޗ)�KOUv^���u���g�=jCy�+B�U��N��6zE��̺����c[t�X�[�ݲ;�7y��?�E�}���J5�铫s�z�rtS|�ff�Ww�f��o��=��l~����Թ28S�2�ߠ���\+c���T�����=*m��y�ȋ<�~'�</)w� [7��5ҷ�Iu��N��>ln�ϫ�t����N�pv���﷜�}��[Q��ξ�	1�������ؿ�ǧgh[�:�'=��G��|���9���|����s���pz �3b{�N7^L�g:n0�_��`T}<s���Nk�-x��G�Qz}�w{Y������❇z���Ѽ�<���H֧�Ϻ=w���+���p��GR����I;�x3Hyײ�ڛ���pR��S�\�Utd�w�f��rӝ��m{ӽ/�����[�s��Ϥ���j��>1��;	l�c�v8l=2tsB�y�]!�2߸d�0'7�{�[�
���Ŋ;���^[���;����bh�'t����g��fڙ(o6�\�������*���������+�U������t�ֻ�H���;g��U�6]m��jF5LP=*j�;��ER7+k��`�X�n�;f���G�Ë�6�������b�D��p�礼xc�w˄Ź���K��]���-�,��x�u.�H卍u���;��"�AT�Z�Ǘ���̂�y��F��Q�Sy��(�I��EͶ+ī%3����ն�33�B��7D�쾊ԏ,�TW�׎vE��`����{�3�����i䡛hsFR6w�G��4EÔ��/��gPk��|��s2��0�ߐ�Rc\�AKQ���m�#ʇ�u�\z��t[�fF�0PV��.�zU�(��kZ�#/8X�c�w��\f]*�
�o1f<)Y�V�*z����(1d��̬wx�.��Qm��o�V�a��p�4հt`�i�
5c��Q{���ˮƎ�M��o$�3rն�����r�jО6#J9��:��[<��=n�����K&��G���vWcƼ}OUgD񳙀gn:�%��/;[]� �8�Bћ�ppӮ�P��.f����h����-�2��ٌ		eį+�7)"���6f�#T�I�ڼ�`ˬ����8v��[A®��`���#ܶkg��O1v��M��XX��!�v��T�Iv�/��8��"ޫ��R�Ei��ZkJޓ5��v�~	����heY���b?eCo���T�ۛ1н��������t�0k����J���@���;�2�u��i�x��|�m���«mi�F4��hu'gunoe�XU��0v�I�j�a�z�W,6��1	��ObwjӔ�R !�;��b��Gz�!v{hE��v���U�:�K=��W(jܭ�s~���kzvBZ/c{����/lw���4%ҚНwN���f��Ժ�lv��|�T	���h�i[�2n0����++L��ޠ��c��}�qh!��EnE���r��D��1��:�S��Z�Ϲ��B��e�3U��u����%whΫ�fƒ4�+x�p�`�|)�X����[�;e���E	�H��w��Rh�WU�=z�ü4Ʈ�s���"ﳹf(��c�,�'�;Ҿh#�I��+J�����{Y��Y�vX������Oo�u04���3h�9]K�����`\on�u4�Ns��r�`�}ˎ�umZ�fgG�'��Q���(W,�;�۶�6��.���zG��k�3����d��-���^�91l�s�M��/V�4�
u��O7�,.��eP��Ů��ooM<Ƥ�.�R��ʙzf;��}��L�2=u
^m*��R�c��*�k��%s��J^�Y�Ct�UbC��R�K����*>����w#���{�{X����i���	�9�K�߹��>^}c<~ �ڡPej�*�T�X�J�X��#+e[ATV*���ŋl�QU�TUQQ�(�F2�ETE��������Q�ب�,QQ�Ŋ1V��4�m�J�*�-��m��cR�+H�U���#m�*������Zؕ�YKUJ�X�+P�+l���Eb"����lb������QU���e���"��1E���E*UEckQ����Km��U
Ѭm��R�m���V2Ւ��*"�EH���(�ZUUERD*�ʭUQ"������(��,*[m��j��cEJإe��*��Q�[T�h� �Q�����"(��YE���b��J�(��e��-JU���T�"1-�bEQQ�m�,b��i!YU-���U-��b����6�[J���e���J�(�Qb-J,FTU%EQT�RڬQU���U�*��+���ܧ�\��'oh�o����P1V�c9�@�ۧ}ڸ�Dw-�{;9ԍ	@�'�+/�=��\�/$�j�&뫒��K7$��\G_�S�S���}��6�%��Gh�b��/M��.N����Č{��5��}��'#���%���. <���Gv%�BQ
���Ve{0��,�~����5)�5�k�Wvl��yWR��߻�ů�}�O�ߓ�_W��M���wsd/Q4�@(��A�}����L���=��C1�C��$�vGy�.2����c�:vJ�Nu'��1�]����x�~#.�������lj����rzL�`<%k=��V)��/��c�UR+���r�_�t}v�<�-ȶKbą�ϫ�t��('x�����]٪[Qq�=���Ov��q�s��3�=u,va�(�A�k�Ʒ��R���|va+��k[�_/m>�^Q�K���~�g�fI�������O�}�,��O^S�fܞ�pm\���~�u���G�1�����Fn���)Х�i�u���dZ��f,T������WpP�VL�1����s���R�T9Id��1����&�]kJ!���z�+w�3�W��T��EID�p�yo��v��A�����Q��=�����˙�R �����Nk�pg;;���ӜߪkIX��d�u�Oܶ��o=���_62K�l8+��q�͘z�=��H����c����|�l9T|_S���o��Ct�{���N�9����aY�;Nv�Y���D�erC�Sq߳���x�����#�0�����ö�+;_ �����;�d×KkFԕ��u���Y�?g�tM����bu�,��h��U#^�5��׾����_;rd�<���6~޷sn�w���g�[���}���Q�6�_l,Wǜ�9��;]=������Av������S�{Gro�z��n�y�o�d!�a���փ�78�~}���B��c޾��:�Sv���N�4�������Xt�g�|�uX����&L��t�z]��^�|"�G�lu߻�2�諽�
�`I6P����}p�C����gȅs܅',��X{�*"��N;��z���y�����KVTEx�3���g�2j\U5�N�LIY(X�����w^p"(򲷕��mY*2q�uv��N�&���gx[��]��,�d}.J��gr̮ޜԲ�v�l����c���0����߶#���詋��>�t�+��V���[�Ox��a�h]�Q8;�ϫ���>�K��`��n1n�x�U��Z��xg�d�L��C���gΖƺ[��T���O-�v�w�	$~�VCǏ�����q��t��ኪ����9��Yw=���\~��c<�b���p_���j{�#�6��͌�{��z�^���{����\~�з�k����pw��أ|�<�ao����'/��3c#��ٮ6�+ε���+���e6�xvl��3�z����V�a9o>�� �}����VfgYJ�5���N��yp=��ˠ]ƅ��\>��[61�iΙW��W��b��B;!d�~�2'����[�]L������ν2{>��M�K��N�D)>���c�V�������0��vu����v\�]����Ǣ�̄p�����N	����+`�&ʞ��q����'���v?��Ѽ���z��-��({����(^'����^#¼�m����Ʊ���|��S�h_ow1Y�8�rv`�Y�d
�F]�M<ih=��	Ք]JV�u�ԕch���+���#�r��]l��u���}����Ϥ��gk�D-��r����k�>mU�k�����nk�s�=�.\wu6����ois�3�z��;�*�{;)��J��9�<��;��7�%���w0:Ȫ�-�k���tI��~�>Y{~v5Mu�T��N.�Aw������6���<�g�W���ɲ/�L��k����{������r�L�"�U����Σ�zO}����~eПon�)����I���q��6r���������|���0��O���1��B����������]���2חv��l&���M �<s���Y6��}��4���p~d�a��+�I�ċ'��*d����d�!��>I�B>��'3?�{�j�c[*W���Y:��=�y��
�w�Ad�>�<��}C)8�L�t=��6ɯ�ē̚�ؒ�2N��e�'�x��I����M���~?����wqկ݅��?a=���2ɶI��4�d���pI�<�w�Aa6�{�d�T&OkI:�l�|w؁�M�o7i'�6k���G��� �����K�w�}퇿oКt��+�O����2��N}M��'X�c�&��'�]~��C�x�q<�d�g��2u*?{@�&�I�����}�����}揌Q1#ٱ��+&w�����!�'9i&�d�^����
��b�̛!����>[���I?z�.�N?&}�94�#b-g���m���8��rq��X���Y����1s%�qm]�U�v����}Y��7\�\�X�X�,��F�-���M���kX��s����ߟ�Ra�,��:ԟ�8�Ő�<ɔ�ŝd�J̡�Bh9�*�:�ɓ�ěC��JϷ��O!�Y���>f��d��c���﹞��箹������5�l�d��=3�I�I�8�$��`~���R~I�T&��Mbΰ�aS�Ad��\�<�ɞk�:����НI�|�ׯߵ�oZc��{�Y&�z�Y8��wx8�i�'߾ĜI:��q%a�C�-2�y�P�Ő�~d�g�$�L!���s�Y<��ο{�=�뿮����~5ǜ��O�S�=���?�<I<���O0��N�k~1$��L�8��'8�$�6�P�+'X�����'Hϩ
?}�!�ߗ��?�޳i�0��¦�&�b�Y6����|��Nꇍ�'�{�q�N�e''��z��O���g3=�B�M�㿱%I���!Y:���߯7x��k]u��k���ށ�2e<`�N��e���1C��~dP�������`i$�߱���2e��`<I�L��$�~d��q
�y�n{���{���������w�j��	�u
ɔ�$�N38)'u?��N��s�<��^�4�|���O2i�����Y>a���	�e��2�s.�2����������~��$�~d�߰$���T&ޤ��J����:���	�M�鿱5$�;���<ü�2M�C�{,�0�_��Y_��'�Ŗ�J�?/ݿ��h�������fY8ŝ�By�7�$���T�&Ӭ+'�~�'P<������u�i�Xm�<��8�$�}��6W�m���V��9�~�W�}b�p|Ì���?2u&�>�� ���h,﬇��'�L2O$�~ĕ*I�ް��~@�,�d�'�S!��u	���~}�z��+n<5	6�G�_��W��3j׬�ˇMNS&An{�F�8m�^����
�{�>1�-T����eӣ\K��ݞ��qG}C[�i1���)�=���O���җ�e�d�b\��4+7.�u0a&ro����W<�����|-�!{��͟���� �I��ڽd�JÜ�Xu��^�&Ru!�XT:ɤo��
�I;��$�I��.l���,�r���Wz9�_��߳��U�Ms�{�_c���0�'��<��C�˦L��M󘁶e��}�c̒�a��py�W���y'PR�>I�M�a����I����O�'�5��IV��گ�~�vͬ��_��#�����|铉�Xq�|�3��Y<�~��O2|��4gx��e��_��i0�i�ISs���N%d2w�0�&Ұ!3Бٓ���Vw�{�vn��� ?}�翤�d�l��M�q+	�䟙P�	�y;��Xu��s�L�y'�h��'�'�~�|��d�py2�6���fs!�
1^�~OfS��~����Pa�M�I��ql�d�s;�	�MRi���:�ń��fLY�I���a�G>q�:����&��'���R�?�݄�h�a�_�}_p���:N3�I�;�d��'���y���hϱL&���IY>@�'ɆCF,����ɓu�i*~͇PRLSܞ�n;�{�7�>�>�C	:�����d�Vg]�N��1�fXO0yO2q���:�O<gX���Nq�IY<���J��'Y�CL��Խ��u�'~�?b�s��w�?{_���q�����RLk8�m��X�Jì�J���P<�����,���̝~I�Om�O����'N3��$�6�^�4��^�5~��}������%d�&Y�RC�'S3�I�8̟�u?2N9���u��X�"�̞~C�^Ă��?N����O̙=����2}5�O<I�g&}F�O��~��+v6���ﴏ�u��#��!�ӌ*N���-!�:����0�q'S'�g䓎y��'ud>/pd�'�!�~Ă����N�8ɔ�\��1��/x,q]�b��Y�������gzX[M�Omf[�f�n>C�Z�ʠp����n�'|�j&X
dcfm9��S.MN� 0��@�)�s��n����g�i���f�T+m�9���^n���/mbE��/�^�s��~��濿�\s�f�ɻ� a�'�2���q	�e���+$�wJ�����'PR~�N$�'����:��3�	�d��<�!�^�4��������C�����~=�w�7�����y�=d��)>�ؓ��O�e�l'��s�b,��~;�IPP�g��J��(a�N&L�O���['����}�o^T�����k��������P�c��d�|����O�N?N��2�HN�y2�ę~ϰ�e�>�I:���T�&7z��q+'�P8���1��Wq�@�3ڪ~��)[6iڛ�kěd�}��	�9�]�e����I��}1�I�Iߏ\�8�L�� ���h,��`'��&Og ��k���>#��oꟷ��%*qW�{�:�_���Jɟ�I�'̜'����P�铬�C|�/Y2�3[��&P�l�2N�z�����O{�u&�Y���
�L��ںǿw��}��Mo�r��o��L��J��k��"���
��a�L��d�!���Ι>d�9�@�y���<�a�v�1d�6J��B#�����W}�!
�u������~J���H,4��s8?0�@�l�6I��O���p�a�I����u���i�d���������1��������~Ce���6WS}>�"J���d�T'9fRq�IX{��
�l��gd�d�ϱ%��u�9B|�)�Xu�|�3>���a?}�I�O0�>W���C.��<_�u����B>�?���'�y�{�Aa6̝�'�u������N�ovOz��M�p�q�I�L�Md�'�8�8�)��:�4ʝ�:k_�Þ���ϵ����z�XOkx4�d�'ߵ�6��y���<���O̓�x�q<����ާY<ɧI8w�����߱%d�I4�L2u>��;�_��G�ۃ�ӧ-�?{v���,�[>oxa\���L��6�ԠL�{��cW#�V�F@5��P�.����2վ�Ӗ�*d���և��{�O�l�?���ݍ�Lr;y(S�s&c�x"�Aʮ�bt�� ��m&2�Ʈ�1����������Œ��Hq4ɔ��C�&�S�l6Œ`�\Y:�ɓ��C��J�~�!:��/i���u���'�;�	�}���d��P��_�|�~ʗI�9%XOκiO��+'���ed���gCI���ɋ8�q
�a���d�T�9�B��'R�O��N����<d�a�?���X�U�l0�Y������������I�,���Ěd��!���&�%d��Ł��u���$���� ��s�C�:���w�T�d��}���P}�}Kc+o�v��G�����ݿ�FY&�z� y�'}5�)'�2f{8�d�g㿱%a���IY:����C�:̘�a8���L2N:9��}��п��Ǚ+����O� ����>~g��H(C�����N�e��}�6��{�XN�2�	RM���V,&Ct���,?ZChu�ɓ�3�����L��w�c.���?�"<~y�9��'5d>��i�̜t��O2m�﵃�R|ɖOf���&Xe93�Bq2ɞ��'P���*
���!��*�k�Ygc���������2��d�a�~��5�y;��{VC��Y'�}1�d����`��$��}�<�d����bC�2�>� �}��H탽����_��g�" }�V�T�2��I�N~�����&��7���:�9�H.�<�f��ԓ�X}1�a�Iߏ\O̜a���I��'���I����Y�0��N;��~��]V�}���a6���*I��ԕ'Y*O2m���_�'P6����l�d��^�~C�Y�	��2��'��u�����yǯ��^�<�߇��q������!�M��!��'��&Og�I���T�'�ӖE��X'Y6ɧ����:�~�;I�'Xk��g�>C:ݮ�����^-�SU<�7dU����޺f<��/f��ko����U�Q�,5��h}�	������6JWܻF��\d�y��G3aT���d�SO+Ʋ�J����q��o�Ԙ�ظXóx_e'�$K��x�o�]��3q�y����Нk'_�꯾��]g�ؽ�����$�V��Rq��w������AC��J�>�T�d��a�u���W�I��,����u�~~O�/������,x��u�9�0�m=���:�I7�I���x�1�l*�� �J�v�d�����I�T;���I�M~�$�d�ϱ%~d��1	���߈���m墪�������������fP��L'��`�2��I���I�O ��$�!�o�<��m���:�	��bi'Rm���6ɶ}ظ���@��}+�B��l�W鸿|u�&�8�XO�2e2bÌ&�������ϰm�d���ěC̞A~��	>C�g���e�m�N��:�	��c�d��1�G'�u_����{���w?o�o�2����a���T�jƠL��m�d�d1g�&���hy'����b����,��&��'����:��wy?2O�}�^�3�����7�sW��q���Y:����`�'Y;�M�$�$ә1�IY2���N5'�fC&��'�8��'T��Ad��\�<�ɞk�:�����[Ûɴ���ZǸ�<��k~	ęa�w}d�a��2u�	����	����ĜI:�c8���!���+'�u
�i0���)�I��`� ���km���(t?z���>�﹟:����T�I�T�,����:�$��u��2q�],��l�=�I�����J�iš�VN�G�� ~?}j��>��p��hm_�y߳����q�������yɿ�2y+:�Hd��k~Ă����v���I�{8�'̟o�!:�2d=�B�M�qd�6���{���\��7߮��w�\���+'�,=l!�N�pY'�u?fÉ��q�s�̝t�|^�4��Oj���@�I߮�2e�,�;� �ğ5����>�/�N>�x�1��TY}NYY��%.^f[�\1G)�Tb��ޗ�%��ٸü3u0(���8kz��MU�HvǤ9]i A:>�n�V�w��Wg��y�ӹh��M��j��>��lu(����8�˻6Ƹ8�|��A�t��i&n.�#��W�UD��}�c��q�o�}
�a��_�J����B�u��hIԜff
IĞO�l9l����8��L��pa>v��d������Y>a��k�b�x��<����w��7�k_����|�2e�_s�y2əϰ$����(Ln�%d�VO�(IԜfL��O���5$�3;�C�+�O0����I��~����c���s���<�[�s[��'�~���L��ӽ�<̲q�>�p�i�>� �N���q%J�ct�
�Ĭ��I�2s�3��u�i�ޱ�'�:��~���yc��^�M��w3���ax�?w��a�a���<�;��̝I���AC�&�Y��Cl���?2O$�l�*I���
������M�{�?k��~��u]�w8ϳ̼�w��=��e�'̜C��ԟ�w[Ǚ&��w�<��&>�&Ru!�{�u�h,�{�!Ri'���Iԙ�ؒ�d�u��><�_�th��>�y�p��k�Y?8@��0�����6��C��b|��I��bٖO!�_2J��5�Ad��w��I��N��d�V{�!Rm&x�{�f����9y��y���������	�O>ĕ�$ӞY:d�gd�:L�a�N������'�:�Y� i�d��}�&�����Y%O��2q+!�������������o^��&R��` m�;��I8ɬ�+��d�o�I2��P�	�y3��Xu��s�L�y'�h��'�'�~�|��o�'1ﷴ�����f����m:�>C��2u+!��|�̚t�s���q�'3�К`i&�ɆN��XM�I�Vu�i*h3a�a?N|��u���\���?��wf���z��C��A�����O!{O3�I�;�d��'�^��O2u�M� i�ӟ}�+'���8�O�:�I�!�~d�d1gY&������^͸����f�֩�a���u8�U�. {�!�ݻ'fe�-�[������W(Luf��B!8�{%��p!��gP�57I�_ټ�CT6�ݍֺ�!�.Ey���㦯^sS5i��e
5|)o)�w�#�_:�V:�'vM����M�:���,hӃSȕM�p�-88��G�·[}���w�)w\�R]�.�'h�׼A@�Ab��r���V̶�L#u�K�]�@�mwqr����6��WK�Ib�����֯��q��9	g�m_k�M2v+�rXb�w%��'�me����[��J�Yh��G��R�k�s����jMC-���n�CRpe�ѩ�3��r��Ւ�^E?�*>�S��$*4�׬Ω�:�c^�[���t��\�u��W�H<7G�R��`��e�Ѵ:8���n]K�8�
����`PV�w�pgUH�������o����!����M���݃�=��0|E���o�WW�	pAV���e�:���}����(^�]tZ��]�i�M;;���8��<�j������쎢��V��	'v�T��gNS��{"�j�#q���<R,BnjX�*WX��Ѧb�u�Az�wϲ#��U��a���mŚC�2�\���c4��K�:����/�u�ı	�iQ�}y��,��h�2�v�(9';]:�0�a�����LY�;�b�m�b�Kެ��%�����2� �:h�|)7���[Y����:�Z-Ҷ�RüR���cp���MЗ�K�|���I�z#�	}q��0F
��wv)v���;��9�V�����!.��D����"���`E���|+Aĩ�Ok/Vi]cŮ�K�v�LsR��
��F�1�ʊƜ���1��:քi-����`�yU���+�<e̋h�4���D��d�i�`rھ�x�Nj�t4�܅���_�Y�*�)��k3���e84��|kzc�:Tt��4�o�{�-ݽT{Ow���X�.� Dw�t,3ԇ,��ĸS��\W�T9��㮤F;���7����A�"6��E�U�`�ܓ�dK�w�ݫ6�;EV�s�U�ZU�t�!J�����A�_c�t!`̹]y�Ι��k{�2���wj�K��à@V4,�!���^`/������$O��vQ+E7�w����9Z�n`�V�Kk�H�՜�Ǜ�\{5��:E����e
�:9���0_a��^��5���d�$���,�����f��Ԕ9����>�{�k!����,\Ӌ���\�f��K�v��U/3o���4�Y�1��]|-��r������k���m��h�[�%�=]��#N[,t�R�G�7GL�QAÊ�'h�<��F�f3yjA9Д��7n bE��rb�y��۩Zc�2�q��ۺ+O ��Î�}O���+z�V�8�+ʄs�ogT��d�2�a�W_U��Ak��Qh�U�"Ȋ+�J�+X)F*�*�X(E�Q`1-��Pc)kj4E�
Ո�J�)j"�FڰH�ej��"�b$X+FT�iDEQ�VDjҩPYb"*�H�`�iJʕYQb� �kAQ-(,YQJ�ڪ�YFJ����UEZ��J�U�����P����@��Z�-J�T�
�X�QZ���PT�ER���[e��"ƱZ4*��`֬�
*"�"��j���c�PZd��PZʪ�"��"�%-hQ"��-�%J֨�U�T����E�-�klm��"+����-�B�#Q@�Ɩ(ѥb[DR�AV�U�Yjь�
Z�B�TYF[DT�H��**��X-B�|J |BD���,�
�L;^��V����<�����Cݘd|l��*�J�^b�uP=�V|���p�.�ku�;ܟ���G�|�lo�y�<e?�*
I�}�T8�h(>� ��'R�:�u'��;���	�^`�'0��:��zɣ:ĝd�rc8��y���B?}d}�H��/��W��W_�>��L��p�:�������7�T<����	Xu��Y��pA@��wܲO0����N�I�M�&�$�s�:�u�1����T��������ݟk���+��<��I<����:��0�m�'�O̓�g?bd�Vu�a�O:C�bAd���'�a?2g��x��&7��y�p�s�}��ٯ�˿g���$�����u7�%a�C���*O ��ZChy�ɐ�0�q'S'�g䓏1a�N�d7{��'Y<�M�
���~��b������rz�Q������	���?J���Ӣ�Օs�h��)����=ܯUra�s�������ܙ^L��7D^��փ��:��I�Z�I�����{��x��K�9/�.K�,:;%k<^��oj�ݽ�Ow�T~R��U>����,w�����
\x"��|�$�`K}h�>7�/mT��v�M�U~~$囸��kr�'@��b5�r<����*Ԃj�L���竇L{s��<��w2�C�̣��$�ʤ~%�]��գ<�cib�F���yX�;ѕ��k�d���m��L��}�Qa�m�U��W۹�)e`��yK;p��\=�(lV�'��5�w����Fמq�M����"[N���7�c��V�M�϶��5˨Gl�����T$7�k�yՎ�g���}�|^t�K��'u������u:Ϳh�K��O�3��}q˻M��=\,�;½�f&d�����g6l9�Lg�Y8v}~��v[{����V��{���)�}s���7)�.�^����{�mM~ڤ��~m����E�n>�=�)�L�Fߠ�|2����`'/��8͌�n���Ǉ�}WS�f���W��-Oq�tS�{���f1}�p�k������w��fQ�{]��~���
�P�i�^�aN6�m���-�ܴ�N�^�tC�i���ts�9��/��gh�.�N�wcfޙ<�7�*�G��>6ߺ���9��bk�������~�]��=���W�^���x�����%	���L���@�Q�:!���>��T��t����{�/i������r�=������/&G��:��D?��K�]��+���m�U��
�z���R���ܺx��C�����)��N�T�7���k6�r�J��m�	R�+ N�{}=�{ݖ�0{��뚩�965[��q���F�_.�X�oL�X��Ώ<���Qv2f�����G��'J}K�w~���}�ָNw�}6{��vn�8��n��,wI��2_^	������w���>�FB�m��Y1�w��}��/���N�2�'�D�f<�x�y��:�u�Uj��uڀw��;���U�\1��*��)G� �\W��F\+ø���m˩a�2�vP	��G_�n0��yWt�ܯ9�w3z�M��\�Ÿ����wN�;D��7�Et&e��������/<��G�jO;������gk��c�㊻����y�q���9n�@fzܭ�c��Mp{{*�wعݹɲ�����V�o��ڷ��ț�z�)�yn�����=϶��r���n=�E�D=�4�[����t�|�۪���l���������w���)|��[��j�wnn�����7礏}rz³u��|���B�[fA����WF�t�E��25j%�Iǥ��{�xpŧ�v�p-I����)RY�;|A�.z�{�ɵ��2�x�.��׋����	����cj�Dwi^m$ո�7nK�����6V;�}�h�z��㤸e-�ϻUbݾt�e�Ky������ lWT�2T���?���s��	���Y�՝���v��KgwD��K�o�:��S#`��6;L��	M΁�|�u�}aY�ō�
�,�U�ȱK���.���Y���r��w�c��x��~��O��k�n!���.���;�w.�='г��7!��w�T~��޻�b��ls���Q�YOq�[ $����c�����!��G�XC�|/�ϡ�f��g��g0��o��u���}��ξ�:݇��5�O>�kr��FL澙b�b�r��|z���ӿI+GK������(k<i9�t��)�*�����7��܋s���Է28S���Z,&��*X	Z�b�8��J��bc��[wU+����?l�{b-ȶKbB�63�wM#S��q����x_�yy�k|��{���yT�}$'��-�41��f����A��¬u�n���c]mq6Q�i�Z����ʹ;"����R�)7s�m�Ի��Q�2i���e���OM>�^"��FN]/�4YS5��Q��@S��m����-l��N�nua���C.`��k�*�[�o���ʉ�1'g������{����3�XX�l�]6��w�^ޕ�oQ��ϽW�Y%� Oo��r�/�ɻ5S�x��F��
ݪ���nO}{��wn9u��>]��QB}];Y��z|���r�����[�*�q�W���Wv^C��3����☛��fۖ��`ǹ���|.{�0�qL��ɔ��զ�Od�k��߾>�Km��08o���9pt��s_��֬�m՞�a����9��7<r��Ӵ���[e�}�ٿ��B9�q��8���^~3&�U�OB�$�N7��O�g�Yn��v��{��~bOg��&�mf�L��7��n���\�Xvu��(얗;����y��<����V2sF��	��	��=��}��;�,�:!�����_S�p�>��]���C��!��^T;�}����w/i����>.]����)���j�\s3w8%x�x���Պ�I��g�t�v��W�Pl���v O��w�~Ӹ	��c��&v޺����>K��.k���Vm.��ye�!Oܥ��q�x*Y|�aZ(Rs���N)�E�K�tj�FNT2p7f�9��Ii��og_89����꯾���d��?��?~�L$����������ڋ����A�$z���j�9lz���,~�f-󫩴7������ R��"��xl�\�6%k�\��a�&Ȩ=d�iyi����:O���y1{���7�������w<ˡ�9>�}���:��̣��J<�~&��T,!�{n����x��M����c�zo��|Cg��>��r����¹Oqޞ+�����Tu+�O$sM��_c��s���-^چ�mB�~|_��]z/�Y\=rW��\�n��������~q�3����5�R���{�yFy����|g�ީ�5�믻6����6�+'8���y�\SyzyI�q�v��gC��Y�Ҽs��4-��c�{\9Z��=�S�fU	��W^yW�����{>�w���Ӱ�R�S�l-�Ώųxߧ-z�:�;�,m�t�Z�v���ޅ\�k����%�)�-�y�����U��J8E_\�{�z3��R?vz����@+u�v�x�LNW��w� 9�a�FR��ʏ>/i��u���;�η\�SM�ϻjΣ{[�-ѷ/�0������>���ﾸc����#O�Έ��/f�Ѷ�_�����C�{�dki��Fz���+'s�{�/2t�ɰ=���'\������v;	s��-���fen�W���>��8��Oz	>���^���������b-o����7�3,�Z��I�2�U�K���~}�s\�<�q��ηE��@�u���p���E��^߾��M;)�}�\���~��;'�Z���6'm,:$9�b��\�OG�0u��x���t�}��/[��κ���F`)n��+��Q���o��;�stM���ʺo>h�r��ڷ�/��
&���<{|�d���e1�H^�I�.������Ug�a?Ir�k���d��Uӯ�������yȬ	-��ߣ>��ӱ�q�<Txnw���}���f1���T��������N����1���Z�W����x���*�L���&�����ݢ�o.W��O#�O'^�ԚJ^d��o��Y�GHVmr�5��Ύ��r�F �x�nV��=�1Bн�d�R'yb��t�E���]|�v�4k��i�c���1�=�fo
�s�fJ��@6� #���|�u�s��ܿ}U��_UJ����>�Z��2�Ѕ�}������~�����c6'���l��<�W�����B�����y�"�����5gT���4��{��k���j�zxG�<�����}�?�XZ��m.�~7'YLw{\=�V�b�j�Ӧ�R��p.w����q�I����N��K�>���i��|����������h����Nt���7����>���Sj�O`��\�>���RaϷ:�C�d�ntϋ�߶u�-��gKO�۝O{]V}���|����v������t��݂9���I�3`|v��g-���)��V�����h��(�v�W����r7˼���.�������>3��.r�;2"7�y��:P�/����,������Vs�=��Z��fu��;!k0����kr����$"(Y�d��j��P��Y��5��O����S����-Q�Wp�Yj�NPȌw�~|e�m�4�^W��~fݕ��ŹBubOx�e/.!3�4�� ���*���/c� �B��h��H��K��GJ�Gη+�<�ã�6kю#�l����m��>����Vw$��r�Qy�s{1K�fVl��g�祇�d�<q9��9��5ʭ6=���[����[z:�kjXs#ȩ��
�aɷ�ʗ��l]"���ݥ���os��܃�uO�۩�nEIl\���	���e?g�^u���/��H�Z�P����a%c�v�ϻ�5���axl��Z=�����gOG���-�ܛ��E{j�������/}lk�~E��&��љu��h0c�6~zs���6�_�Ú����yn�6���wUA��la���r�y�Iy,7/p|�3d���7��}~�`-�_�@w�s�}�;�(�e�i�7� ͷ��n=�G�\����)����޵�=�w{޸�ж�b�Ǜ�����{s_�����vׂ>�²F�w��/3��S����[�Pm��x�o�#�0���V�����I2�qУ�o��쒰�盻�z������.��Qvc<!Ю��3qNSm�&�v��.�P|u�fq��h� �L���t�����1䔦��G��Bc;����\R�U�Z.����[Rx�#۲Hۙ�9���Wst�V�w�2�~�����t}$���ǯ�w��l�|��+��͏1'�z����t����������m���<��GZ>�Ŋ;%���Z���Z��)��c���ט3����'@��ס��;�wΈ_o�8G1ˏ\�E4yN��ߺ�g����#q~R��p��^	����:�<���\Ɯ�L@̡6�{��]�6P�����<�fU�2����RV�S��Yuy9O
��ͫ���� T}ڟ˱}�������s��ǑW{���B*��+���8�ӓO<ySD��{-M�t���Ot��lF���9���=�of���Svp����s��;�%։����:�J="����N�w���� ����`�/��zo�ϝ)����D��Mԁw�:{�h��l��{�\}<{\�8͇1�ϣ;C��c�����m�E߅{eu�N��i��B�Elm�,Ǌ�s+���O�����G:��a]���pG�>�o>�u�u�xN>����M�`e�i�N�,W�]�B��6���wm:�e.
Z�^�i�=�����U�j�i�,R��U����b�sy�gV����7��	�(:6�P>����g[<��e0���n�+W/l��C�{*Q��p��u9[��)��^����ITy�����"ȏ�V�J�oM$.���e�'m
�u���k:�q��VC6��d�z�*�:��5�De�ֳ�a�V:Oν�h��k)�+eG�_�x��H1²��M��ɮot4r�-&��,���]�8W�$�"�H;�dy�������ą
���eo۽��l��vpǗ,�]43+i>�C%Z{5�R��!x4�v��;t���]s�����Z���wi��甀�y5�5�Xq�f%�u�ڹ	U�_�!�~#�gZ$�F�={�����^v� I�;v���d�Jƨ,�8dʒ��i�aM�[%��ۨ�ա`��6�5��S���h�Ѳ_r
�2�]���&U��������4p�Қ�5��tz������-�峲V�I�!�G�;j�LaD�[C:���w,���n1f����^Y�y��e��N���jر}¯��v0r"�2+�V�0���|w��p��)u��WqvqI�]�X�9���Rb��ќ0�%��f���d>�.�O*Gv�s�W�z����,R��=J�-aL�%^�w�:c�i�>���e��Zv�~��퍎�/�����x�>x��4�;���Q�G��A����.V��tM^bwJK����*���M�.(6�+�G{�%L�����J
c��u��8v� �-Wsqom��bw�k8�F��K{��Q�|y�8]j	u�1�Z@ᣗ4�^k��Ǒ�냱	�v���Ch	���؀��{hc�_^R�3
[Fig����u�ϒT;��Wn���M��Ԑ����Q\Y��{Lԃp�wdeL�{���2!N�P�@A�7M�h�[Ž`Y�A� ��Ҁ���zN�k=��M5S(F�\)��y�E��%��Ṽ:S�:j��'g"Nu�րs���;Ә�w6-�c�������"�&��iuorO{s__P\�-1@���W`h�S/s�[H�ṵ5�1/�U29Ք��9iV^��wxGJݣ\9H$ЏY�ot��8��c/t�K���r���34���:��ʼ�^��`ɧ���Y\r�o����S��4|{��;k�A�M 1���N�8*�ˮZ:�d��ܫmMø_;!�j�꾍Xu���f��{���F�VJr�����Ua������a.��ۇEՙBS�H���7B�îL���ռ,��M�XF_�A���۫��oP꽎.�����t��.����5��<��������)e �J�R�֊PPmX[d*��Z�+VE*B�R�A�mD-�l�j���IPh������J�P�"�E�F��F
��Eb���U��B�R�%-V�Y(�YFV*�����HT�%B�ڈ
%B,,PQ�kZ�XQQm�[EX"*�mB��eAAjQF���QB���*X��X,+d�B�!Z��V����TJōhEU����eIEE"ѭDJ���kR�*A`�0QA@R))Z�T�*,F�ЕU(أ
EXT*�J�H�"6�J¢¥`���!YET��-�
%�l��UV*����@DF*�"�-�KIX���H֬�Z�k��3�z(P�����da+���jdꛝ������FU٘Wl��xMTm���ü{ǹWN�31���W��}U���+�{0��8���s}G���~q����o_ݛ�X����Q��t����=�Kt5y[=�ޣ���i�B�g�����׈�k}�]{�ts�Jy�3��^���%x����<�z�S�����)�s__���=t}���n˩�m�#{S�ܰ�}�i�)���p�x�rl^e��gRBmz���V��"nL2?g��f�_;
��>1�˩�Ke��S�X�{SF��Ԟ�y�&f���b<�����K;N��>,P;o����\��e�sg����)5�k��������w�f�d���gi��i~�qުΔU���{�_����;B:��g���D�ϼ����eV�m!��I���]����Pm�qf���!҆�o�n|c�.�úL�֥�F��W�>�t�ɭ㵎�P�}�4#���b��qS���Y�*z�@���%�����] �6>i���oz��O��^��X��}`���ͼ��n���Cjwj��R��υ5�H�gn��G����й��f�.�XwuowQ�`6�R������B�]2�S���=�]�Z���o�b�`N�p�?�����g�@��{���}���=,N�^�Ɠ�WOk}�]>��
���ͺq��y�y���#�1H^�M��Կ�8u���U��N�#����{8߼e�>1H���qƠ[㱟S�v;1&�;s�p��}mts�(\�^�fvO}ݷ3�i���1��1���v��*��{��c�����rz��]�:V��V{����������{�`���$���3)�s���8��sQA��+o��9�ή�������`���n���;N�o�^A�3��{��m����vW��J��~7�òT�N;]3��0Kr�r�����=���
���Ɲ�T��sF�~�K|�j�rc;��7#},����}�o{���v��||cy=�Y)}��V�އS��$�c�����Cc �Μ\���{�[�xw(%�"��o�v+�Mn���&�\X��6m�g�8�8v�m���T	�$\��#&ֺDe�~�n��	��E]�ueo�嗸�턎�r���%X�ҥ�Z��&u��s'N���Jxa��gz��IuY�pY������G���4N�.A�矾����$l{s'���}�6N�+�����M��$��|��}��������غ�g�h�_����������٧�dW������OT}{����ؖeJ!o(��t������L�Oc�x,a�>}i����M����2_^|&u������K�_�==��o�{��d��%���=3�׊^v����g�祇�d�g���J���|�uI��j꠭�7�zc�׭��dx"��
�96��Q=�d4׷aےsc����ę�9���Q��?}�K�lF��\�Ł!z3[�����Rl�ptǷ��S����h�����Vf{��۝О�����������x���6W��w:�[�ߡ���oÊ+��}�-�N�ަ�*,�/�g?.�<��C��s��������׀,��Of�ޕO��c���5,Q�֪QpM�3�V!0й������r���@)�8WKj�h�u�έm#]��U��&ܺ�e�w�DV���^A�'�� ]ٕ].�͘�dT��{$n�WC{> ��ɕj�u���3R��C[��9�k�����^̣��(��9~�龢��{����^�/6��ښ�V���C�^�5��ѭ�V�~~�Fd���X�k�ۖ��ǹ���\��x�J�����r�cjG�������@[f1|,y�'.`=;��k�^Z����Of��\�Pۘ����oY�u6�ogrփ4�d�ۜ������%���֢�M�bLə�/��n���-���|�_�og���δw+�Z\�
��O���N>���cy��s^@5�����u�	ܳ�腼_������E�!�Y^w�^s���>�����<��ܙ8���\��ۭ�!d���oh�y����8`[�`!�����'�/;��%m��j*cm����{���ӻ!O��C4�_U���(�w�����*>��ShL�E���\*ԼQ�:�N@��������o�����A�m����)��j.�q+��X_5��&�jY���{LE�F_mÉ��#��up\�ԋ; u�B�T���9��w%�f����f�3Uε���ѽހ..����͢�p��}��|6�56��H�un��������^�zڞ�uj�מ +��R�����>q����/E�!�tﰗCD��s(縝[˩I��4gg��#�¹緎�<�"5��pv�|�Y���b�{jw*���j��I��߫�������3�{�xM7��3�cӑ��_����;��R;�,4�Y%�Q�z�>���=Nw׽l`y/���q����=��\Nxn��-�ogjݭ��wQ�T�>ͦzA��r���f��e�|����z��|�\��Ak��ߛ=�l`�1��k�k�<�ܳ��܉vOn����_@N�{S����i����Ln�p��\�b�f�	���O|{�e�p����6�_;�Y����d��h��ͬ�]t�:=;K�F��o���A8�f ^�y��%��,4֑���p��pߡ�T��A�T��̋���R��;�O<�n����-���#k�����ҹMI�v��i��J��Z�,b����+#��@�Vkw/d�
������� �'nb�E��R�vU�R	���b�kK��gTޔ�Rŝ;�}_W��kزx�g���A8�w��7��7�lf��L�̐>�,��C3۝�;r��ܺ���>�pQ��u}N�T~�_�{\ٛ�s����i<��gz��<zc��;6�[4>�k|�h�����6Q�(6���jO�(�g&�7��kn��`u�vB�x�˽3k9�5�����^���}��7؞�N��]�J���0GD޳Ɠ�WOR�V�{,��T�0�o��M��w~֥���?��9!�xg�v��vaxR3~_v*�)����lI��U���r���k�0R[!l����+�<߅������6�D�ݽ�N�$��Lx`b:��]ߥ��:1�s�_%�
�,0l9X֥��o�[��f�<�3'�#َ�<{)1[�)C<����ș��[E���/\�u
Ӛn�o��p���OL���$���x�2�aߦ��9/cDx�5FI�oS�_�޵dv�J�����2�e�)o���Gv��꺔�
E��'�XΊn���f2����fAbL�q�ڿ-㽕�_ӯ7v��\���<"=�|l^S.�i����"��7�KN�����Δ�nl	�qs���p�"���a��ٚ��
��q���W�}_Wɭ�޿fyH�~�8m�<�������
���.�C�-񒗝auQׅm����=ޏw��)OJ�rɬ�s�>�s���2���²���X�(�Bc�X��+�*`�~�����}Nj�ܴy(=
�p�`�z�M`�C��9��r�|\�ݩu�/����*�����-�y�וʨn,��/.Y.���M��d+����L��ACܷ>�y���ZZ�ckP�@�PJ$������*��U.���c��f��Ru���������3rJ۷7E� �*rǆ�_�Qi.I�`%�D�)�g>w.j3������Z�t�u�Bu�m�'s����oǕ����\u�;uD(��)�@�M��۩�K�7{���~�-�P'�=��hn?{N�KƳ�O[9��L70�4:R$�q|�X�,�`��gg��\�BK�� ^�r��`�e^ ��_�IS	��¡��E?6R�'����6u�Y$�Z��W�,��}E�}A����ǎ9Fև(F5��z��+G����õ���ii�p�7�O,�@t=� ��j+h��Sa��ރI7=Az�ƶ���`��<k��"莅���'�����i�r�L
钂�[gnw<�Q�p��XlA�`���t����Ƴ����uw^�V�1��y��� ��2�;�ug��@����<�
W���L��s!�����L�k�Z����3�Iy��o戠�^W�eؘ;ּ��f-�C=�7^qp��N�7|�;d|oz�֫������uo��& ߭�r:Gn���Bƥbc�=��Z|)'��oxK�7٩ʕ����%k�
6����{	�炞<u�*�[�֕���Z+�=�����W��I��z�q����=2����[K��=��i�����g�[�Ԗ��]��%���j�U�����wǵ�A�m�q`�3�P�Y���rm�U�;!�W�ޭ�3:��=Vt��+L����`lDq�0���br�@�w�����X|}K�{��ލi�g���e���SI\�rN'�o��Zn��������/}��W�m�� j��g~����=gM:��U��j<�U��:'ƚi=��X8�ewV����:���2�	����4c��]�Tk&R=r�%���q�#�̽�μ�$ޏp m�������qK+�����6u����}�8O6�&�gZ�6��ɲ�P�z�t��r=lE�R��-��R��#��^��'�u%]ȇ���9ȹ���Y���n�D��H2��]r�f�1�7�A�ᎮA���:���o����p=������E+ѳ�^ε��M���6a"�o`���;՞Kg2e�UGΔ��Q��&��9EE��`�I�G'F����<����rs�b��B2�L�ر�S5�������g:�W���4�zRԬUC�
_nq���A���K�Z�L���W�/CL@xʵ;��wW�`ޝ�Ԙ(;��]-/
u�����`�ޢv֞��ʙp��jpH=*�u���,��{���R�3�B/�b����Y�m��h�K�avk�<F�����bU��8��>��y�~������[D䆟#��>��Q�a4��t�/o��C����0�a�N��n̽���r����0R��l��7�pSԳ����H���k�Ypa��k���e��f�A�o�מ��z�{(y(�,+��"�ά��{�p�v�_+}��4�B�[��h��KP�s�i&O�o���@|;+�[pX�9m'�^��C7{�~��ZTRZo�������?0����>6����������������#\z*KG]�,��X���,�;ٯdl�YD^�;��7u
�ͤ�\�N�=ż� 8��0�2�9oD��%R����d�� eΤ��Sz�<���r���%���r��bŬu��������D�0�-��#����L�YW�+3�`n�X�l��������V���甇�W�{�d�����;��
��P����x{��s���w0+�u��:��\nW<��]�08�>���3�VȰ��	��q�Q�-WP�.��T�g>�UUqƵL~*�Sx����N�(K�0���;����e��֚�$�N=:�)��W�����ק���86�į索��a0�96���o!�y��L�t۳\v��X�F�~�v]�b���L�O�2�j6�����xdF'��<���ü�>�Xd%�!HV��i=z��3Y��ܙ!8��?���1�����?!�'�}������瞳����Q�i��ǣjG��h�v'�����D���x(S3�M)�m����pY�=��Xs�oo�;��o%ޜ�똅��_f�+��Eן�z�mġP����ޞ����t��B}����d/�U���(o�ɗ������$��:MEI�:&j�q�푢��5ؾ��p���:���-ы7��<��8j�=!�xg�v�˳|�iJ��;��綑����* 'MO�p��Wh������X�*����ɽw�.Vx�u"nӴ�ud��5��V	R�l�]�K��0��t�9��]�fb��"��sy	����O����uH�{u��)n�Pƺ�R��FAS��wQ���z{��Y�u5�vL�!��G9�7�7W���|Y,*G��vn���]���їc�u�d�2����rV#j�un�bQ�ݧ�v,�X���q�8�
0u���TX ��W,:�_7��ȃZ���D��2��f�%�-̗�1�e�%�0�������
YOsv1��4r��<R�+"�c��J4M\�����b�!�3�@R���V��c8�SԫYYd���d �JLwHkow�א������g,Щm�5��ak��ӱ`�@�;s�]ʳ�GL�n��������U3]c�K��O��kx�/�`��Qv3��2�j�r˥G$��,���p0�۳�W)F����3T��˓S��mG�v�d��!Fov1�����_7;S�t��8�ËM�ٷBb��,l�ع�����khEWǬ���kO5���Vp�nw}�f�f����VAx�*Z�ͅM"�}6�;	*��)���6oX�.����]Ǹ�u��2���[�
����y ϯl
���1���j�o����  OI|�#);sm&��T�wT�`5�46�\���v�7lS�90l�b٢X�h���J�[�-r�,F�j&�H�Y:���f����@��+b�m.u�v]���{a�3*��చIgǻ���Au3�lɮ��h��T��A:Z���9�_t��es@��*�-�쭮U����v����x��:�B�(`���@�Y�-��^%;����!֤B�X��k!3����4oku�)gS�ݙ����fg'��T�R��={�o���Kr�(R��-�w��`�����.c�&C��ޢOY\�ʥ-�}D^�6��2�N�%SE�(n�>�p�C`�JH��J`fv-u��ԕc[�#f1�*3�ϒ�+_�����q~�Ċ��R�X�j�2m
7����2آ����V������fV�6�Ek�h���,�;�Y��t�E/�A��l�w9X4>/�]���tu^�N�$�gEJb��X꾠m�x������ݹrN�r����c- �_M2�;���ٝ@�]գ��Wu�>ǳ�]�w�1��@����&b��߳L����|y��{n��TU�[ܮ*[�4�W.���G|r)����pff��nL٨L-C_C�$�b�U�*U�����\�;���껾�"E\�����a��Ƨ ��Z%��_mC�^M��N���e��'[2��Us����&:R�`�Ue�&�&\X�*NH�>n-Dî�L0\r�Y�lT�ۛ�������΍7�Ӯ`W"�J�Veۢjֺ�o��>vze�K�C6w�6RY��9��3l��R�
�e@Q����KV��m(
)*��,PR,�%B�[kP,XT+
ъ�D��,��
��me�m�H�-Z�!mFDT�D��m(VT
�mDcA�Qb�b1P��J�[b�Em��Q�
J�d"�2(��#m��Ȱ��Tc�(,R���
�Qm�Qd�E�EX,�(,,�X�l��V�U�("�*�F������e-�TJ��J�D*�,+b��R,R�YU��b�(���b1"�U��QE ��`��Z#m��EX�ؕ���b�H���D#,X�,�PX"AJ��"�`���EQ`� �Ņp�����J�ʐ�qeaR�)[B��(F'<'��U:�]G>X((8\ץ*��$2���2�wf'�ͼ[_k��;v��u���A@�	��[���}jط�������0�5�G�{�I7�_���={V^��}��`��l�B�&c�Z��LGJ�ů/���9�.S��0e�g4�LWV���ߥ�ʣ��/���҃y�UQ��=��;/!���@�N��/z��G�ݔ���J�1�Inx�{i�Z�Ƿ<�[�<X�{"bw,}�D�]�H���ޕ�+yu�	�}{K�G5Z�<xb������*�}�Yy����uҷz��&_�.*>;��t"��Wgk����lC�	��o����A_KW�u��l׆{��r��G���9�lM`��bu-x�=Ճ��#n�����P<И��QF����m��f���d��%x��w�4�}L��s���Cyڡ�1�����e�c�ώg���a�R�0Ui��\^�r�v�p�oi
Ͻ(���r���О��CY2��U����iC[�b'�0p���U��v^;�9�����]������j�!����8.�>��9��`�6%�Q8����[Ĵs�.g�//Y�&61y��V0-(4�U��$���mo��,L�}�q�-��P�[��Z-^E�~��o�X�:���b���%��f�������s=�3k���WYX劉�s�/�8��]hJ�kkT�xE���$����^��i�^��� ����d�<ղ3��b��={�����P�W2����@�:C��S(P�R�����&Ǡ����Ѷ�}������a{J �x����.S�O[92��D�D��I5n>;yP��e��q����a��
���a��\f�� ��~�*g1ю��M�KBݼ��������c��XG�Ѳ]%�����	��]����Pfd���Wc��mhyGw�����U����KG��s@ ��E�`�\EX�ʎD�5ً�t���ў�Ez{|�w�}0��ݕ��t�e��6_��؈�GПw��l�%��a_�6���;Q�/rܵ^�flw��焫�h�r�&������L�^A�
��~��"�3$�J���(��}t�n��{�C�k�
:�E���5�߲�-�Y��k�U��>~Y����:D���W����`���5׌u�ܱ豨t����M�{��cO������F��=�/��r<����5�d:��u�T^���9v=�Y���~'��R�����ȫ��&�Pa2,�۽o׵��E.�t�eP�Q)5gNWҳ�]�D�*�%��b�	�U�'*R7[Kt���ϲ��/_R=Ļ��m#���;u�3�@13Wu7E��5�sp�t�pĻ����3��i��z�"�=ܬ�^�qܝ��ꪪ��Z��1M����1�-?��t�倹�¤G|�BO�fu9x"��}S��x�g�o]=��j�i��v=�VZ��Q�'A\�1=��з��#�Ka�3�����%=/Ǯogѷ0OEQ�3��掆��0�-Lr�Q�m}$�?U5ƎcJA2���������4�p�3}�	�=cH�#��^�X��}2���$%�1��HX�ή�VOc���De(.]����}�ř�l�E��,�S��Je��h�%�%',R�.ߖekU���������r�0<i�[Hu���j��ִχ)�I�����L�س��xunWs���k$Jv�g(�7$�1{'L���L]b��#]��t��<u]w��hc t"�^��Y;�g!f|/��u��G��-+�y��[_nT%��b�9��ڍ���ecW���5����W|t���߄��b��&���hg��4�.���\堧��>t3�z�ۯ#�5����^T�H�u/�h����s�_y�C9�Mz*y]Ӟ��o����y�8`��f����� ����$�{J������ܾt�!����N�]g~ʹ�� �3u��9�7�S7��1W,�WY�F����leN�r�e_Pk�!Z��]�xkh�M�-� ��Q���y5�C�h������o`�].s�_/��W�U��z�G����Cw�/�n���邗���`ۂ���Gh颈�i��O�OV��<�C�$׺5�p4���~3�E�y�E�ո� �XԱ�+�\=�XY`׸�wS6:�����vkz+���LSy�_qpuw�x{*kc�'����7�[J��r��8}ޝ]�*=�fi����މ�&���m:F?�y��p��]���;^��=ř�ٚ������ݬ����PϽ��ռ�L�⬰�M��ɪjs�Z�S���
s;ڝ��i�)nٙNf�x�8���<���n�k��.���0�[^6)��p�.=�Ҽ����=^3t�-`���r���<pJù�|^VZ<N��zvK=���tĺ��T��)Pd]p���ik�QOJ&.mC�����+�ӵM}fv6t2��N�������@��W����f
3ѕ[���U��c��}.��5�z�(���&�۷�x�ً�����j����b����	�x���P�Cz�mo��� ���B��>�ȹ�vy<lIb4�K�mU,��Aᩈ�w���%v{�y%��}���^�w(��Y2��7������;�.��$���4P�3����<�65��irl�o��nL�2!ogR�p���k�r�A1�uLζ���ힿ�}_}E��{..Y��9�����֬4Ht��45rP���EK���o���?
��5M�1o�%v!��c9%��ZrSy�5"ç�zfq�O]���#�!��qQ,�.Ϫ��y,�]���o����%�hX��G�3`j�Z}7��ˇfQ?"H�刁���]�oz����!o��x���qxN��`&
6�dA�T�Hi���lL�0���5w�=�<��Ȫ"�d=����	-A�x)|��]�ໞ��#M�k�R�3v<������C�do�F�J�@�R}��?����g�F3�+w��w��<�":�V��\����f�K�Z�j�)>�W��U.&)����~��qKHו�N��=�S�E��1�~�'Ϟ=�I��5�+yggX�7֏E���0�XB���.�x�%����yt��	��������⳧ǈ����.��}�b3C��N�4G���-ulζ:�e��x�j=�fe;���՞���r�eY����uS������=�U�g7*��'�c�p�i�o+E,n4�ì��SՕ�;�X�֊7�gd�m�����ӦN�e��m��4���0�9Yv{�V�Ֆ����L������w�0̮Ԓ�Gq׀6��Za�%]�R�Y�Ww|)���}�}��r8�7ޘf�;�i:M.$��(P�4;�E+���s��ߗ����ߜ�5U�턣�3��yA�繲
�b�)4�Ui����0\�{$��H�V:1_�Ρ!7�q��wvCvw��[��ٌ���X�,��T�	y&l-���*���e���D��"�_�J�Rp���S.׾��]e{*rßl�ĳCmQ4ԸKb�*���v���7a��kLl{�쓽y<���=�G����׼��|�x�P�W2�i E��0h��[��j���_L���ש�`�;�����x'c�[q���L��2��[�'���� �4���e���A����ӯ�I0��Br��6�\c�0k�A��_�9SK�t��J������-�~�M`���_�}�}���n��-fua��Ɂ�+�������;�W��Ut{��7a����L��t�_�|*WIn'��3�5̅�VB�k��q���2Z�N�t}�L��ނ�DxR���<��hpV��-yT�U��H]�C�F[�{W5�nm�R��>���>
�T�NS'�

����&��wx\�+WMw������D+���Ս���-�}�^���ԭ�ڭ�tj�F͜�Y̤�&s.���)5�,�������ّr�������PS�*������K��E���U�s	V1�m�d�:G�U��w�y��i�*X��	�����ɻ׉�)M�C��
��M�w1i�K�.��.N���ϫ��b����k��s--�o�ć���7�Zf*h{������v&=�c�`j6�igޛl�h�4�7j�G�"�pw�'��䜯����~�g[ �z�-�|���6�t]Nf�N&v��_�K�Fx��Y���c9�c��ap�&ˋi֕c�hv��	6�32U������ޣ��{M�GݯGO�rޯ����v=����4��t�j%�o�L�)�
tP�d�iD1��ޓ��m����BI�'������o,*
�j�~Թ=0�/�_V��6i��0�����T3vY1�X�.=���Tk>)�v���_s>}��?5Sل\�"V������9�ř�}�	7�Yו;�臘^L�xߞ\��|1����uy�6L)yC$��m!�6�M^N��|9MBNw��z�}�J������㵒�V������q�FC�g	*(�9��Ϛ��.���L��Ý�MNo�i��K�2/v�&��tƀʜP�6OᔟOY>t8�߫9��Mᝣ3f���KsC�bD��w(�x�'»�r_c��x�o����;�͸��~і��?S=i�r0O��>".�To�c^K�|w���O ��M1�&���'-�,Ǖ1L=yh�H��)�.�]ïq�"�h���A��M�Y��zr�վK������t��%B,	b����B��k��댼���HLFyy�a�lM{���(��jFs�ay��h�
~F/����lvA��S���,�*y��*l����h�}����I���8�ޖ)w�B���`���OR���f�邶�*,��Ǚ��s&�B�E,�%�#�����:c"��=��==[Y��}g��[{���u������Nq��s��,M�W�Ww�C/���m�ccĘ�Z��^�QÜ��@Xw,ڿ2��j�`Wm�i��O>L/���x���*5Q���o4-���ٜ�&e�s$�^���:���=���/�#��:*�o�v_�9�A���7��ӔX#|���W)�������p��֏��Eb����2xKԇ&LkE�z��AP�Yn��h�{G�{E,=�Z�(%���z�Թ�7:۽i�.�L�B4.h�y�g�9��}�=]��$�G������٘�P9or�9[�9��ABK�� "9Jf!��K��,7������8^�Sb��49(@B�z��9�i�Z϶�2����NX���XrVǣ�(����O܃���u�<���:����+rLb��z&2���ð�-�0�sj	���(N�k�^���S�m�;ex��(���E����������G�j�<1����[Q����:��e��m�\{��dňE�46�wh�ޤX�WPL��vo��b���jM�_�^�'P��%�!�����'g�3v�!֬��wh<�>�u2�u�b����5��Ի��H��f�je֘�3+�x�)3%ޜ�TY�Gr�*$�E��J'�x��z��t�.y����z�P�{G��n�~S0s*5���9��^H��6±�;[����8=�=�YS�^�w��N]�N&'Qk3�`�a�ȃ��휐�<0(a���R�tv�׆���^W�	��#^wYr���/~�szX��J�+f0ұ5�P��<���M}��x����߄�Fϥj����σ�����E���w�aF�4��uf��S59!��5��
4�e)��5��{7@��h�4�
ŗ&;�B����w��;�v������3��.Ց��jݩ1�4,�S�����1uj��l��y\")�i�<�/K�?���'[m���iEb��2����I��nR��Y�&wGF�YJ�A� ?U{�A��x�#�e&+S��TF]�ș����΍�dMԯms�3�C�^����I�oJ𒷖vk�J�do�FY�y�H[J{�c�-�����۴��P��9~�g��3�qY��;G"�Z����:wJ��1Y5��޽�d>�>�7KW��n��6)�rٙ�;����z���#|.X�ձ���7�LUM�'^n�������OS$и(P�47���,�C���.�.����[��U'��~��P�cH�*͊�Q<��meUq��&�*{��ƌC%�}��]ng/e7�r��������+��Q>J�ԫ��T^��=7޻�w�|�eG�z��ᘧJ&\��3��P���ZlK3PJ�I`l$��1v9�K�NwT����b�u�z��{p�{e�={����0�]��E���:C��Ye��jV�i�|��Z�(Pr�|a���^�M���v<E�����O�1=l�=d�>��w3�}T0�z�f���m���{��$R^�`�q��T��Y�3�ڨ�ܜ�ea���u��r������|�yCdն�{ѳ>�-�J_u�݁� 8�f`F���(.��70�T �on��5���L:PR��N7j+��:^b����Wf��v��PT��h£����U�V�586tC��;�݃ ���Cy��.�VI�A�t��
=���b�9a�sd������\����𱷃7����z�������[����:�1ӁMd�VN�[7k���B�NK5n��,UO��ʳ6Uš^L�sL��	Qˮ�Ų-#y6�J�a��ܫ}
qܐ_1\:��Ƚ����(�_)��Ɵ�l`�Hk5v���R�}N�qb��W�U�>�Uܦ����]�p�W{��}�N[!M��J.�N���5�W+1�:�}�M�С����
��t|����{Z�T/���(6���3@���;��� �-2oxT�x���|��^��t9����
�k�Yzh�}ل�ԥ�+8oG�j��W�Vk���ޏA�t�u��\]����1���[��o��w�M��-��ѵ���솟@`��5O���V������B��Z���m�&hu����
���ڵ`�m��!,�b���aT�dz��IJͶ���ǯI�	��%�Hp�=}L�]Ky]v* j�D�u�Ul��եǠ��3=ޣFN+������Į{u�e�^d�� ��
�h�+O���`Z�I��
��
W.wa�IˠM$I{�r'@b}�����gMn龅�]ǅ�2�K_*�ڈ�*,"�V�և9�\7�:Y�Y闽��
i�):q��&�Z]��[w}�9tX�Q��؍;\�ۺ5s)r�@�W�_Y�kpÀΥX/xo�a��p�(��ؤ�ν�uq����Wz��o��w���Ү�)�\o�'�����+7����[�N��Y���-�-��[�z�_�^��n5�����^���8�W�|*i6�{���F�ʱ�&�>�N���q7�c렋k��}y�T��n^�V9��#�/* Y��a��xtY�c̕�=[2�D,�g|>�?>�|�!F�hn���qf,K���CV�%�`��(���mK�o���l^!@���Gcc��t�=�t�YV��|D�1��On�-�q�J���Xz2�c罷�7�͡I^H��C`3:p��@P:jZAn�j��H�ggm5o!7�b{J]�ۋ:�օ�����Lr�a��gGAJtEv��QӮ�2�al����:4j����d�]M�����������%��Y����^����ө���Uׁ����790�\vgP����7�:��᳙H�\�����Ea8�f*U����:G�t56�uu�Ij��T$yx`�(�n��R��}����tM�5��ۺ:��m8�r�}[��,�٩�ً��������U���¾�������bՑ`����ZQ��(��EH���VDT
����QQ�"(�E�0�X�0�E��,���TUE0ы��1�a���mQŶ�DW)V#ذ��-�K�E[l,0��&-�*4e���-�)b�X���UKJDQ �cY�QL&14Q��*����TZV��`��j�E��DE�Tek���3�j
��Z�T�*KZ����eV�*�QU���EQŪ�AF5
�H�U�-Qb���mAb�E1iEb�E�Y
�b�[eJ����PETUĭ+�""��ڶ�ETaR���"�+`V���b�,TdPVҢᨠ����R��R�U�UcF*�����YO���qr�>�ǽ��밷�U{˻E��ݧFN��j%sm_>��C�P;�@^
D�V]����m����χ�5�4O��I(��m{ᾆ�>k�}&~
^y�_�9SJzy,�j� p�~��(����Z�4�U}�}����B�Qj�Pf�̘��+:��iz�oV�L��E��kF�NS2�K�R/� �\E]P^Tr'�vbÌ���t�FJ����w�y�RP�\l7v�Ϥ�F�bJ^V]��h���<F���(�6�����~�'[�[��Ov�П5����h���3&ܦI�#�yV&�� ���{;2Y ��Su���ޤ�_*�9�W�I�c^��b����5�c�p��(��mz��ʢu�e���i腮w=Y��_?�o�mTL��U�!K�v�������?o iy�\�w�X-R�r�:^�t]�^�{O
U"6r%�d��0����p{\D�c��Nf�-^��#̘�9MrLv�ز���n��nY�"Mx�tK��Ԉ睈I�]��J���M��i�6r
��O%�^8.s��3�����-ZX<���Va�~������xr4��H�.�����g.]�YAG�-ǔ��<�
��1v�#�+/]{f��ɒ�(>��̺'�wXw}�
l��h����}��5�v h��47ovX�=�.�o��.��K���҃Y�@5S�72�f��C�G�|T��[���i�o8�s5�,�����`����i����ʆ���,/��v���'�+O�;�zן��u�w6s�J��C7�l�d�#c��^�F�	��X�h��y\�=��G�����`ϒ�;	9X�v;:�3��Y���$Py���|�z�$�]зl����YڹO��w�)3l�>�>i4������nd���kL���$�y�ө9f]-�N�^o�k�e�>���قb�P��)C�(���cY@����lƼ�9j�:m�a%��fe�p�7��ϋ�~X9��,�R��
����$q6�xs��k��@Wh�䝚�f�V��F�9~���U�.�h7�����B;���f��N��=�u`ͺ�k�vn����z� �-�0=���P����'$4���:�� �fո��Ŏ�|���֏����Zа���ZE�邕�<�.&�?%��:�k���t��Obt};��X+�d3Q�kQ�0����w�<o�����ƥ���V<�C^И��{���C+ja¨ye,<γr�AW�C�8MX:ʨ)�D,Y�N��y<��&~�`<�s�Q>Z���TMÍ�������
[��JPW�8_4�[,�
��K�W�q��e*���i�IBNI]�QW3�d	��ݬZ8P���s��83��F��Gæ�O|��E�L���2�g]���,\�|��G�^n7ݡ��I�,��t_�60:�o�V&��~�i��O6l�m���z�_����{���]�m����P���w-���-,^��WR�.��e,�6s�۴Fؼ�f[H��t �Ti`��fS��#�����m<�p��G�U<b���l%���S˼�h4� f\8;M2��fp�r��9c�=+��e�G�n�Z�z���ΰHc�|�D�抭"�
��K^Ҋg�����8�o!�{}�9�W�v�50��w&`��q�2F*�� �s2�*2�u���𿟲�!50���[��Ë�x)��74zќ���Co�v�oR,Y\\X(.�̵S2��J�+i�=�J74���Z��E�{��ɕ��8�Z��!�������S/>�L�z�0��^N���wId��Z��\��9H�����3�L�;�GP��*%�ǵ��/�|��Sb����ɯu�tS��.aߎ�Ŕ^�2�()֤;�6�;T��6��]XU�u`d=V��ҥ�i�>�-��'1��b�g_��7���3z𭬙����
Z\�p�������o ��aBMw �;�Y�KN�u1;��@���~ߢ�׀M���X��`�j�Z|"���O����|͸y��{�{9�D���[]{v+��NE�cd�E�q�Ev�8)�'�z�5��U��'`�>/}ѱ� $X�T���R��}�X_�uÙ�0RR(B���=$ӹ���2wc`Ϥ�˳�-2�x�>�@TRVy�ww�c�����q�B���L��{=�& ��
۰���ϸ��}&��k�(w������T���ڮ�;�w������c�Oc�'��8k�O����2ޕ�+yu�	�oþ�x�K��^��J�K��Ĵ,��z�P�\p_�كݗ�18���߸�^HOb�xÖ���Ӛ�3�$[Sq���U�k�y{,2(�w��{��ϩ�ŧ����GP�x�gFy]�6z�9����c�X{J���'�P�B�Cp�`��R�S!�b��Z�BFs�n���{��'ul�}���mq���p�i�Yd��|��$�zS�l^ =�Gp<�}+M�e,�Q������8�v�wZ�oT�Z���x���)^��z�*���M�=�qJJ�(��w�w}�0u���d5̆��s��V��Z-V�>z�SO d%G|��U�:uo�]5(���o��=ܺMJ�),���u�ȯ����@[� ����,{��:�P:��P��j��qx.]����I��ݡ��]4�����ϼ�oӼ�xJ��`�6%�j�񠖥��Kb�؎?<��;�9�/Z�>�|��zׅN,P={�����
j�R5�@�ޡ�1�*�KW�~�낥Q9e�
�qg~~w5yM�u��KE�'?z�}���}^[�w2����*���.nelԧo6x�0�D��M�m�C�����g�q���*��*�n�M�_���sk�T���dyl�ϟ�Cs#])4�U}�P#��{��-�������ee{rb���X��WcǚR\ds�zyܵO��]�f����VD�#u��{R����gu����%`���.�9%"4����>�E��R�U�n�+�bU�X�N9D�s��=�ŵ��Z*ƹ��	��7��.�ȋ}�M�l�b�g��9|���9>�
Z��R��{���i��'�|��<z����1w�q����d��<;����6��Wa����o��b�8�@��E�[n�j�Ȫ�A�9�c1�Yۤ1��{��0s`a`�Ht\�@���͑>lgU��f�޽�a=ǚZ���ʾ"���t�[�E�3���LƩ)� �[ש|F��.�f��G��F�5�y\���zſ���xy�Oƶ����dc�g�C���io������3�eJ�o��O��<o��C2��Kb�L�W����P��qg��tS2����"k�����:y�=lf�H�Ҿ�/zg[C�{�lث�6Zd���倹�[���r��`��=�ޛ�f\�u��3��9x'���B]���;���VGM]/Z�R��ẕu�4>��?TRjt��+�#i��=.\��;���^� �P���-i��}�wuz�J��<+��0*�6�\���g���κ���y�hv�̬̯%ܔY,*�~oN�玣�)Z���#��T��4�W�3|�&{�92���ڞ��Oes�/C�ط�U��Ѣ���&��J#`�0�!��]H>�|��\"�����+�5q-�>0wI�a�u�������h�U���i3�	�[�l6���ܻ׻лS�{����7i���)���rVj���fZ��;��3�t�I5�������fp�~�y�zr��ܗ���{:X�t7`��Pk4b�'8��q�8�:^D°V��I�ǖs�0G���̼�`�@n��s�hQ���ƴ�D6	�p���	o����#��g!f����Е�@��9ڨ:��c�@;$Qk�N�'�~�7�[g N@���j4�����]��KA��0P���IerS�=F,esk-�t^�>u��n��;k9y�yY����_��'$4��!ەDB���L�5�{�do.�Xw�j�P${p{��뚅yo�����JǞH��2���)�o/��]=k<//z��^,!a�םb�����Ls�#�>��T��@O�xX��'��?Wl�r�v߸çV}����*u��+��ˋ����!��{���[�U	^0=��-Ou��(zy�iz,�R���sn��A����Պu�3�l��cu�ή����Jy��0_^�h��%Q�=��=�����n0큞�K��q�ꕶ�Ͳ�f���g��Je�V7Ƭ�8}�Ĳ�٘)����=C �wV��p��GF'I�~WA�O�2L�f�=�PR���9 ��*�M2��fp�s�>	�iY^��@߳�J���8�w��p_�e2��Q8��é�����Q`��a���P�K�����]���B�}�%Ʈ���Nn��ܪf�m<����h�
��̧V���t�`���+u�����ۥ���/���rĶ�s�rY|��\/m�*d���-�E���XrW;)ΔVR����cie=��W9�)E��x�b�ls�4;�wŌ��[m��V���P�c�g����崚6
��,U�RDw����ռ}��1�	��Y�>s/y��(28	f�ۻZ�$X��qq`���ꋿjY��Ўw��Q�����!z�miqr���z׭�o��E|ġ˪!b�p�s���Xߧ5M_��l距�0�uĦ=�F�Sׇ}�s�9�Q�:|'�g�NаC:�W�a��d�zr��|vz�bR�jx(T=ި�=6Zh`�,k�<ʖ�a��&\;�4C��p$w�T�7wWp��`
51�<�]P|�v���E�Γ��ȃ���)㞳�eEo}Y�ٚ�ǣ��6<%u�B+ah��5>x�?��X_u���0RJ���T���e��N�����f��s��	)�w�^S�"�f���p����<^��"��Bm�cQӭ�Ma��Ik��ߤ�����kQp�M2�Z���픯\E^�j�Z�w{����l�AˀC�v�gFT�s�^��,k�J�I�oJ�{V�Џ���5�-�!�{i���^Y�]��dx��K7g�Y�����:H|+�֑��|�
�B�⫽��J�!�q<�Bס3.�p����Rg���î��w8�rHq�Y��*
;���l��Σ2億��kU�^�/��i��L��f�sz���w�u4u��}[cM⶯��N/f�ხ���� {�"��K�i���ܾ��[X&OC����B}��>^u��\)V��P�6(��N����/	u�f�
�1�������
�S�b��
ý	���ژ*�Ԭd(v�w�5d8�=�����*����\�qwH����e�|5�~��J��NٜU��}Nɡ�jc����s�
��1]�Gؓ���kE��Barޮ�({�ٮt� Y>񵩎��Z���|�[����o�:g����H�Byg�-�w��	C�Ã`��(�8�9�0k�U��6��s��yvyē��Ꞵ�|�\��6��,������Ó�v��v��e�S����uy'���R.�B�<��˧S�6�תX�,	9��}=-�`ڭ�v[������秣�a��'L�4M��?q|B.�6�TRX�j^y����={U+%G�j�vy�!ÂxT70�5ҏ��Z��2���CKq`F禮��7�G�d����6���mj�@g#�\�NRț��0�Eu�@��gjwKj�/-��x7�BR���n�Cj�kky��U����r�У1v����t�`�c���K�j��ɋp�]7o�P��\Q�ƅީ�Ȫ����bu�ĺxN�/�j�v��gj.c��kF|��'�Cs)%])�T�"�dYڭl�[~�W�OW]�4��4�ZÃz]$�0��탒R#A�,^.��޴�68)��Ɨ�qd溝0{FZ��VH����8=o���%XLƉ�2Liv�L�605�V�{��'���cC���9�z1�^ױOP�W��(�{#��'�p�5VФx��ꅾ���)_���k���LY�k�7L��UZ�ԩ���5��,xc�^)��5�?m�J}��\��������K?Vd`�ζ����̀�^�>�fi�1�ѝ�)v��M��W<��M�����=�_���b��6Z�ly�\�9��� ���
~yל9�t�v�1���9��32����oW�A��x��e���8�ţl����u쩔��)����bhS���k�G��,��E��`������i��6(ΚV|�ԋ���|��ƿx��K�*�����4Ұ��3}��&X�4Ã������*5U�{��y�Eh
ΤvsѼ�t�Z/!�[% ���e֊w���FI&�x�R��̳ �K�|�%���J��ܧ�.M���u��L���q�-U��~y��J��t�m�.�	�Xs�1:�X�w[�2p�T�qS �sYШ�64�c��ҮKǄ+F��T��e�_vT�K^�ޱ��_z��YL^���c�+k��Q�����F��}{�HGҀ�6��K�y���>�6�Xw�j���ڴ�f��9w�J��[�*��)�	��
: ��z��:�;��I�S)t*�.�̎K�o/����\�PIK�K�H���ǁ>
�um�%�Ͱ�a���݆����u�&V�*r�U};$�o�؏eY���s}[0Dַw�+����ӡ�Y�pv�`]1dPI���9�GB$J
<�z���ս	]7�}P��$z,��ރn���,Q�Ѳb�&���]:vs��M7W�y�*kz�
d�&p� �w�n�I"��z��ǭ�6�z��r+|���r�C`n"��	E��/��t;�Ȣ�}���#ժ���9[J���̣l���CI�R�({�7�9{l��ȡ�oru�h]YWkqU�fZ�kkGt%\R�3GkT�W^����Zr��.W�\E�;4P��r�Y�I�K�� �a�U�aCgx�g��f)n��p�Gj�H�أ�W�@���n��S>��X��p2�Q��:�ƹe���RŒ�]�p���(�
��D����0�x&n��2F�˖(�Xݞ��{��.��Nd��1���ʘ(��yyFM�EJ�u
�.�<`7���;�X<��X�Z�I��Y4[�7i�ǒwQՊ|�n�Qj�Od�K���`n�֡G*P�E�}\�t�x��w�̩���a�m*ŏ��Bp��G^�٣L����9O�`��3���t:�9 
�-U�^jkZ�v_�����T#� �Y}ɗ�_	}�tm[����ܙеY򲦒��n�rڭ���N��,B0� �.U։�f��)RAi�;s%�ec&������yJ�hqK��Q��]}�Y��4lV�T���k�
.���vZ�����C{,
�x��x��Vsn�������TΜ;x�ر��t�n�ףAz9�³EXP'#!�3*=��e����7ψd�f��Ɖ�I�㦌��̛c�d��(1Ժ՝. ��Y��u#�qz��P����ʧbd���1����|��R��R�@X���>�y1����4���{��U����4�V�P�
�V^�%����wʚ�mu8�p%�����m�k�:��llgvg"1��u�N��Vi�M�G�_tT:mkF�VR}�!�(��X(�v��'v&���;�I6ތ�&�X�V&-^<�[���x1�p�J�CN��Em� �<�0f�F�Kю�TzLՏd7A:]�Rӄ�n��_-���$Z��߭��3��g��O���kj��ZTR[TT��)�
b�h�!l��"�
�%UEX",E�a���qe#�*�����V(���%JE�(�b"��Q�""
�a(�ATQ�a+b)kB��b��EAdb�
�,DbV(2��Cd�f��TšF[ekQkX�� #
�H,QADTT�V���b���F�b��YRH�m[B��(�QQ�B�D�QP
��Y%jb�A-���D�E��ŀ�
�"����X���D`��aD���+a+H�a�����*Lb�
)1�aUUEp�X
[AH�(�����`Y�`��1d���acY*��b�ዅb���Á����1�`��*�0��QA1d�Q�E����YE`����E�MR|G�Wnǹol��w����7�;:."��{�*�:BsA�Z�w}*���l5l�{,�骭���^v��tj����\f�|��wqd]�G�ࡨ��2H�U�w�1�ř���׿yN5�K�Y�����|1��m���w3�S��^}2��(�y��Wm8���-�ju�=ZØ���5��y�Q�t�Q�Y룧�� ��ڮ�@�:Q+LƲ�dWۜl:݋��}����s�Tx��������2�p�+5zz�!fZ����A��}Αi]:��,o�ؚ:��&�����y��D�\[Q������0�Z��`����@��h�E��6����)������`�����!�]��tf|�(^}[D����pJ��{RYU.���ݫ��dY��MX�O��on�B�{��E���7�
^w"���L�z�q���o�fK��ݥ����2��Y�/����s�~Ix���WT��`o��W��~���Zz�ɜ��
�ϳ�g>[���{�p����v^43֘Z:�$����>���p��o?����^9ZE�����ϗ�x@x+w������4>+sk;�v\ͼZ>8s���ۅݧ8Q�vQk)u�m�����63NRA�t�xt��=+-�Œ�+���������@��/ſ-�9�jX�*�d�i�����|3�	u���	�����繏F1�oU޾�t|Y�.���0�t;B�@C��q��v��7���7���.ٶ`;�z�z�����2K�5�FUr�x��8=�1L07�����駖��s8�8��B<��j�Ƭ�p�S�g׶��NfxGa���>��P�p��s��wCw���hـ{�[Y�-�,.���0B�lˀ�i�ZͰ̱N�(|��J�� �����ϕI7���Y���w�]#��i�eVژ)P�w��f%a�e�I�e��?vI�7�oS/��۹Zb�q�킇��g�V�`-�ѰWK�����ʷ2�����)L�Z���sϲb�0�Y�`�ȿ��ꖯ|��b�\\X>���=���[�q�,]�e2�v|��y]�kA�q��y�+��N �_�%K�\��h�6u�`�����n����ｇ\\�m)�n����W<��jϏ	��==o������W3�����]]��P��ڟ ���j6�^���CIc_���=���L0֢Gq{��Iƶ'J5���~�7 �Y<EE��])^]�����r)ȵlt�(ؓ�sS+H�;{%�:�Xh>��0T�S�"���}&)����m�y<����1^X�׾ȩp0P;��t��z3��wv�>�"���ڳ�5�z�(
YSc����Je��.T�ut��!c8`YX�]�.=P*Xv=����� �j�n2:�_�nWc���P6*�	�u�6<'XD/�p���#�<ԧ���\�o�I��V��Ю�祔����X���wl�9E�%���˸q�����H�����T�_eb��J/ýگ3�3����-%k�¿��6�N8M����#~�>�V�/J��"/�Ƽ�Y%%ڻkte��8ȗ�z|-u�Y+BHne�+�����7�uto��Gy��<�~��ǫ`��\o�V���W�0>���qY��;G�y�67'����,���>kd����������W�J^u��u¶�}�lPm�3�;���ent�ܕjw�M��i������x׍��5e�VډC�\p�47�z�Qd����r��GN���֧��c>7oP�C�e�G��Vnԩ=��m$�ʔO�ٺ%��72�u�[r����?D���#��4b�d�9O�{���a��iP���Z����l��������՜n}r���;DL�Ӽ�D9�/�WrɆ�F���ŀ�=�v��s�!�n*�{�\Y��Af���O:+��)����3X�5�ܳuՖ̀ݹ�ثqܢ{4��ɷ�	�Ы�5�tf�k:��W�
����CP��H�1�uu͛��3�h�XKޮty�.�t���f���_cg�"�)�.��Ȣ����Yּ����%�����T�/����&�z��|�x�.��j�.��:�w�4�ͻ@��`�JE0P�����8�����:�,i����=�yG6:��g��#����M�d\�������
���*�o��x��j�&{U�vGco"����w�J�7�m�P�,�L]���p���4���W�S#�Y����O�/�~�����o�wG����eL��Wc��mh��9`��� k�/�s�%�����t�.�ϩ�/��r�~�k�.�f_��9%"4�J^V]���I2^KN��]�fZ��y�u�~�mR�b�mօ%g�L����*ƹ��LƉ�2M�#�+�੹���Gd}ǲ��aƴ!L�V4;=�[Z|+R{G�׈�.�*��{"�2���sy%v�7�nG�ی�'٬�_[�Z'�b�ZW�JK�x���[I2k�k�GRgix=F�-��kw�7��l�n�,��g�e�<ybk>������>󖫯}�
GמJg�b	�ыh��8Wq�C2�AkZ���8�����r=������2ȥ���:Ϡ�pk�{6���ր���1yȵpos�Vk,��㖀#����O�+A0���핣8`=3[��3l�o�q�ö�h�uۓ�E؅��\�w�P�9�7������lqX��t�Cs�W�;��f����#)=kzӞV���N�gSH��L���9OɁq=^�;��_q	�!Cǻ�]��e@�`�Z�puu����h��=
c|��]�l:-�QC��{�=�tFkyKP��"��T�}��s_�+B(hC�;�C^�^セ�����|�^;+t��> ������hw,��/�O�R.��'J`��>	�]˱�N�^8Y��l�w:�g�̐�����p�/;Lؤ��;����2��K4O4�>q��8�ԃ���=^��4ud�}��\�v�7jy�5�)�'��b��e����m� hs��*��`��|X/�=n����N�;jz�íz�_�ܬ���LB�L��'�a�k�t�JΉ��t��������7r�L�K�}�R��+�w�C-p2�#~�(I[V1Vj��.�=���UW����������T��ەzG+�ޛΙO�s��4O	6���Q9mJٻ�
�-ҳv�U����d��G��d�";d�8��B���2���v����R��p�H�����n��K��`�s[~5\w<��7}��GV�������G��4�%�gX���3��9Eڋ���-E/�-���Vg3�lbN�c�1�o����ڢ4�ۄ���]�巢�D-�=��q�z`�~y"��EF�g^*9��tמ��oZ�`lV�X9�谇�i�?�Z�Mp�2�.��=��v/��ƣ���%���:{ly-lP��2�|�<GN��"Ȳ��7�W��xL���-K������֭��%�(E�<���cK&���xE��Y{�4�<���[�j�]�c�ʷ��<{<�NL8Տ|&�Jv�w�����.�׵A�G3�h���:�U��}~�7:�u��Y�g���j*�5*�q_��VX#ڜI��3>�a����Q�{��3�p��5���/l�����G�Zv
���n��X)m�jP�b�!�e�s��-mgS��6�޽Kv�v�}[}s�83���u��e���P�[je*E�b�rf%�iEb~����C�)�9[�q>#��0)/��({��p�X:/���-�!Z�e��g}S�D�?<�2���MZщ�>ɈC�_���If��wkU�ԋ�\\V>��;o��[�E�͋���M�g&Fo6�5�hk=Z���7f���R9�^�B�WN�9��'m�ft��NB Z�ƻ0'�n'�gf}i����Օ�s>��&V�,QO2�롰 j������ge��2�&G]8���2���]&k��T�NHv��es�C"�b{���{�ؼ��%~uD/V�VdϺ]8�-�V�k��ξ��N ���{��}s�-*&�Oz����U��e��D�yQL�ֺމ>팂���4ҺQ���\m�����ks����[qĿ��x��A��x:��/wd��lz2m�8:Ik��_Ԝ]x.��c��Ƚ��-f��	P�T[��:�z��t]�/8*�Pò�>��!�ְRgf�1���̳����眓w����n�$�d&���Z�Z:lL���/)����3G�I��7:����v5&�0欄+F����d�Yԃhp>�Y�R�U�lvR.z�n�������=x �k�F�N��
Ko��x��P�a*��E����v872�R�/�(=4������*�xd�s��֚�}�s5��֠���gN|�<G��!_]C�ܧ���?[��ؾPs�=���t�۵f%�J�e�Ga�`��ؠ��f����������r%U�/_8��,���%,���U{*:���K^!�����Cɖ9�kS��SmdI������zf�7�ߌ�O�YG�T}�uv�:�ku�h:r��D欼�܄���hu%k]I���`�����Y�9�w�����z���vt�8�����SQ��կC�6��M.��[jeT:��(v}�����0�� �N��\��BV9���oW�g�:�:�V�L?��=>K�>Ih���]��TP�rï-�]3D��3}H�V:1X2u	��z����B�H&���~��J/����d9w;k�5s��/܉�(O,�҉��;��klܰL4:�L�!�s���צ�<g�4�y��R�/>�v��r�)���
�[�0]u���]��_��3)ߦ.��Ҁ<�]��Q�0h%�L�C�WRg]�����:�KE�[�[�����8��0wB��2}�d��~6&&��$�_ZW��a�5�Ry��Wjf���6�>���i�U҅E�j��8��Ξ�p�
e#å&���GR��\t�K�dn�����z.ؑ����.	,���Pg�ʙ0?}����Z0,NX�lL��D���\�G鷙�0_�[;���X��+,^��,��7��V�0�j�:���nJ^/�uɭ�܍]��']%馁T]^��KJ��,�e��.���]�ez��=����3̌}��֣��2���D&���v��6��}����1J����B����e����Y���2��������Ig5��t`�-|����3��������,z�ݖ�p��n��)v�e}���7��Z咴&cD�pS$�{5�����޼>S�ԙ���C�P��
񪕍?o��Y��{G�׈�p����`�t�y�J��{^s��z����6��.�j����ֻ��3�x���[I2k�}�!A,�^v�C��cw��l����0t��m,��g�D���Ƙ����Xƶ|��i�<?LM�R�ec_W��
s0iq2z�{���μz41P]�-t��z�Q����<;}��OY�*K&��5��0��m�3)��<\�������D���\�xC'3��bn��'i�u�X�>�4�G>zjD�z\"ӝ�y��i�t��S����Ѯ��c'�m�2���CA�����Cg��<o�4�=5ݖL�CřV�US�8��z����mԝ��(��L�z��h񵦠6��G5R�w��4��^,��&ʕ#h_
/7����-��>0>ׂ�<��W��Ͼ�h�f��t� �� �.��d���A|Y1�ו`�n:�� �Q{�čt�άF���ԡ�������w�׵3�*��r��N��h�!�	��1�N��d��]u�[K0)DŇ�ՔK؃��|DDw'|�wh�mӧv��IW�ݽ�����mAo�u�iM�vI�O.C8�P����S���y�^��ɘ;�L�wH��(�Lƌ���n�m/�;;����������9�o���*e��-��S�,�*b�0Pn�9��#8e���>�Ո�R����wX�K�;�Nŀ��X*e��"�gL2��-B-b��g{�6�b�ӹGE]H�5K
f��p���� Ͼ}E�{]Q�Yg�Umagv�x+gK��g�ѝCN��!��BX�]�b�巂�D�^D�i��
^��T6���}�v����Tav��=J:Gڬ�g���2�I��c�L����z'��5ʕ�`��S"�N����%��
�v��E��X#�t���8�0���|�jt�R	j{S:��؛���]~�2�њ��Z��upX�f4�ml\���N��p��c�]X3�}.�>'�oz�r�O���bV=*���L/���x���ǥ{͊��q�3���S�U6�o����_k�n�A�%me."�#���Ew�Y`���S�e�0S����;P|F��%�Z��E�j5����O�J�&Z���v^ౙ�U�=�+��b/p^_Q$k.��I�[�9��Т���w�QT��ў�%��9C�a�y�ܖZ��9Zk-$#V��Ǖ�rU��#b�`�H�΃v6P$�R���6�feb�2��z� �n��vK"HgG�x�8t�yy��y��Mol�Ii[2���*s-��X��\�W�G�U7���kGuҤ��\��s:���J:�3Nl��b	Γh�['��wi��$Ih�vhƈ۝�k�j�B���W�\���6e�:<CY�̻�eEXFԋ)Y㯂ˤ0��[�luf���d�C�J��0Ī��:��N����I�+̻������kt�]��k��֦�M}a͚k�e���>�xz�rÕҢT����X�^����0�,�&0��&�S��e�B��� ��j�N�q-,d�Ao:�e�O ��h�S��F�$�˧��2���ލ�S{'oGg��.��\��P�u�N޳�����+t�65񍃸9bٵz��6��TgP}���]5x��C; ��Pa����vۭWn�}��!�CD;1��M�d>������mh,��Zt�6�d��g4W��nV��,�[�}|/�g^�<b�em����pa�6dx,?=V@46�j���0�:���DA�E9u
�f��	#���Ҿ�ǚZ
��z�ǰkbVimM�)�e _Q��mR�"�����7#���e<�uum*h5���v���8us�gbN���wf���hH�u��V��J�+luj�pǮ�����	�01�G�hv�hbN����t7��0rw	j�or�7�A��h��Y��F�я�����f�=}���	���5�IIW\FB��m2�i�f�ݽ%v�j��
�����,5�С��I�6�6ڗ��xw��Q� �!�̆����,Ǘs��Pr��(�hn�-L�7��4
a�_M���dZuq41��;bjɴ�ݼΛA�b;�S}���y��9�]Bz.�dxH����g!/	���X�� _f�X�H�B�G{����V'����{��v�T�V��NQ����s��.܉��ٷ�9�X+e�ɮᮍ�B�z��e*����%�=�N�ыz9� �����5x���#,`'���|��Ҷ*��(o��yg�[S/"r��;�p�8�s���j1MO�2����];��k����7��Ɍ�������V��3i	X$�^Y��m��Iȷ����d�8!��@�)VZt&�y�x��c����|��:{�溵dǈ�6ɰ�h��Y���G�a^\M�7�J�P�}���:S��s�v�δ�%q�Hw�� �
�KTV2N�=�:�ob�)<�`J\v�S"S{��^�u4��uY"���6ۻ��h,��;��V�s9ю^rEyB��jV"D[iT�E#��j����-�h��+)l�X�%V5������0C	U��%��,RV���B�-���X\U��YZ���*-�pȥJ�f!1jᶐ��[b�T��d�3	%B�	l[�\Akj� �T�J��D(����-+
��a�a�AEd�EŢ1W���dm�)�
�@Z*![i�A`1KLR�"�DRa�1C	P�¡FD���D�����ڥ��L5m%`HT"2(V�,���1 ���1fJ�Q�U�a�ֱ*J��\&,�2a�ńqJ��(��BVa�S�R,0����j�,V�
��TĶ,0��""��
ԋ"�k�$�J�3	�XVB��H?R ��2s��u��a;�M��)x{{^��M�-h3fub<B�Zne�ڵ�^�5��F�ʹk��ʹ�"7Nj/'��s�{{�oM_���m���a��eR8�3ʴ��`��ٗ��L���z�9�7��S+=��cqOH�𝴬�9���V��-Vb��d�"$��A�&K=!��t*��)�bk�t�a���P�r���!��1�9Xk���h��E�U�uȧo�.�j���u��cʧ��^c��b���1x��fl��v�_�QB\�~������冸�݄��ǱJ	�c�x�~C~�6�"�=�����Y��v�"D;�0��sK9��>���^!<\*��\A��m�
dۄiϔ���}\�N �k���N{ԏ��
/=��{o��r�Em]?V� �5�i].k�P�z���l��c����)��ܳEQ>�̷�z�k%G��Xg�q�Gˇrz�f��H֗���net9{�^�|
pͼ���/[X��K��g��9�j��p*:8(a�ѱ�:�!|8V���jS��U�-5�)�������_�^�S/��oL��P�%�\��Z:e�CyL�$aQ83�˘C��s��`�"�-�2{햱���.��.��czV����Zhq�
�w^]�	�E)��XB�m��1���@4��yy��N[�����g-8W%k#�j)�wM=������f���|�L�>Ǡ�(��Z�V&�9���:���j�C;��eK�Mg3b���/j�L��B[��ؒ�
J��L�r��w�c��(b�%��Ǆ�A��e�b����Ta����&w;o>C�X��;��`9���в��n���;3�X��9ۣ�����N
�`��mK�%qQ�e���k�����?Ḁ�,���oQ�jw{Ü9���\�)!Ꝏ�D0J�	��_��ΰ����%�4U�������x應�'��T��9+����ǰϯ��+/��b���aބ�JK�P�W"m��O�l����2���K�YL�ә������C��e�G����u��=���l�t�ŵ|kv��ϧ����,����c��"�X<��$��rޮނƵ��A�P:�k#(�zF����9��>Q���՞Ϳ��^}r���ȑ���"d~��r!�Yl܇y�ݡ��~�G.}�{]����ތ��Q5�\��֞
U��t���\�g��6Y4z��"����֔��:���ɻ]��3-XyH���Q�5�\��9�_Zeө��M�u�}u��u����*�PN[�;YcE��Nv/�p�4����F2�N�괳-�<�����f���>W]E�}/eH������]��u��A�ך�7���j�����O@�`"�;����c4̈́�#���=G����t��
��v�9�v�Cm!}�e��mK=\�'8�����}�~����z�ɔL:&&��$�_XPqX�q���Z�EV�c��_d�Ԟ�.�p)y�(V'��2d8r`�o醑�ғJ��du-|����:�鲱��dZ/�hҠ�C��|��Y�A��*d��"�.#K��S����!ͥz�EC#��{��5��"3�[ZEX����g�Ot��ޗI[P��+�	)���R�5y;���S;�v�.PA�|��� ;�C���KO2��F�L�-3�tU�J,Ɖ��w�x�U���t�����I�kaͩ+��hx��i2��V�Oh�Z��]��`�X�w+p*>M�>�����HE��C��N���Y�ֻ��3�x���{s#xY��e����-ܭ��xu�Ƹ�|{ι(=6��<t��r`�3�x9`ݵZx�\�-[�)�<Ϸ�zyiO��tX)���N&��}��qX��n��Rnw�Mk��o�Hm���R�iW�u�C�Ԉ��t�NU����x�{;	~Q�����۾Aߪ����i�A��i���z�V�&�Sn�ǂ��]s����Zk��]?H��9�j�Ým�c�W]G8⥘�
����9oo��ˆ]�;�trݵ���7ܛo!z&`�piE���}�P=����ze;�����yQCP�K*K�}����m#��ԉ`��E��`�.��gS�uא�~�jn1��>yZf}Yk����6GRw�*0�8�J��P���&,��z�PۯA�:�����,�-�ܽ�Tk�G�K�x�M@l%�;	�]˱�[ƕ�9��C����/���E���	���<e��AL�-6#��>!��F�h�3�N�$9���߯�z�3���Bc�9��+~�=�b�]˱���ƙ�t��J��vN�+MzUS���d>S^����Bk���R��LT���[���)hY�r�A���=fu$R��,K��V�B�*uP���%�����-��T˅�+�t�)h;+�^�]�oq��������ق��V���ig�����9M�k�q��gϨ�����"�b�wcyy�N�n��۩���Q;�n��3�*���xM	��!�:��}�[�B���.�A�}�e7l�`��v�`�t=]v�}=J:G��,�� �m��L�R��Cܐ,���l~Y[�q��n�$��ȿ^:�m�/�dh2d7�Ջ+�۷@|��{XŵӱȖ�V�BZ�6���A5X�ִ��x��E�����
�=����{+�5�z��Ś�����M�IW�4;u���o�h��}��sk9�:ʿ,�͗�\�G+���XԱ�*ǜ����>�:osndY~���M{<�ݚ�7ܶJ+�s�tyw��&_?��G��T�;�n�[Iͭ���Zt��� ��k7�K���n7�W2`���[�q�7��m�zdGò�f}%��n2�^�u�x���g��9Btz��g���=j�ME�-����B�Øue�0S���wy4��P{�ܞ����I-��'\<����UE�R�@�9xP`��e�{Je��Z�Q�U|�n�i�K��8����RX�Շz�|^VZ<l-5�U��(q���ɮ����_W��?<��Z^Լ��y�0�.uB\�h?�
�v����[I��йv ��R;`��ٮu���4�y�{�p�覯l��똄;���,2/讀��5\u��ӗ$7��"����k>���1ݗ��?!�����"�=�͙^[8"xWhW��t{��Vy���q$(6�_b�7���̱޶�ϣ�];?-6��W+��w�F���}���YB��ڼo�A��������T��uT�S'�O�OzW{�.���BqK�mԷ��3�@�������a�9V���|eD'T�fG�5�Ŵn�Y]��x�k������0��͗c���v�nc��'f)��Ă�Þ`�k|{nw���z�,��"W΁-f�V.k�P�z�z�P��-43������-`��d�k(�vv[��6=�V�Եy�K�B���j+�9�^���c������0��$�۾2;ൻg�VD�WoS�Q�a��L�0�)��H���m�]�a7*JǖÙ�0ù+{��Y�z`��J�).�;�Z�%#�.�x�)����7��׮��O%(X�;�Ցwy�OYC^�tFs�����\���>��h�/u>S��M�h�n)�s���yn}�O�S<�\Lp�ס����;UX��;���p� �������1mX��wveK�����ӱ�j�ŭOX��ږn��=JD�o^:��=]�6�����N[�#f�=�"���l*��p�0��+0&:RW�'�ΰ����`o�]�P���+Eo��m7����L�bu-x���g��F�����+qT_}U��T��7�.�7r�lݞ�؜��c!X�R���C�9w��ޯ�_��U����"�+�!�\����ծ5�O��������yV�Y���ib�x��Z�97����4u�k2��PJ�,��ʷ9I�L�W{�uz��b^��m����}�GL7�c��nc������N�����p
���gXy���Uj�8���R̾��3��k��ʜ���˭h�RK�� /�xw����F+2u	��oWh��m<���s�GMsc�����z$���عv^;�9�P�X=(�oӼ�zP��Ϫl��]K�z�a�lVڏQI�@I�QҮ/Ӵ˩S˂�p�xl�m2o9ྥS{����(�E5�凱���.��2��whG�`��sS
�e��]:�^��ֵ�oG��7i��3��4��N~�OK~Y2����a����Α&���С�i�dť���=iWGk��b٬��Ǚ�x�2�b杭ɓ!ÓC,�&�&JTT�[��ڽ�y[��>�V��q�}e�Π�E�2`~]����	��L���?�3�̩�U_���wr+��OO(��W���җDf��f_��9%"42zz��ޣ�;��x��[�Kn�z���68'�㚕p��\2���37���� ���VE}/�j��H�r�D��oB�V4<k}��Z|+i'�x-x����+@W�2�g�ey�&qn�<ߺ�KD[kp�)K�1#�mw��9��\q���M9��9��K��+W=�6���d>g2�*��W�[��wؾw�qZ�����n��{4wVD�Mw9���L���s�^��Ƀ��&>�5��ݑ�	�Qk��K��g>�A����F޷��3��X#�G��!������� u�?��
%/\�����
��G�lM?e1���P{rǢf�e��/=�׶�����,x�d`�3֌��ະ��>�\���QBz�� cn�D��ߓ��y�ܴ?m��A�����hFƎ����.t9]vt��d��5"9�|a'i38S��}�A��i�\rS�)WV>���S׵1��se��+-r��>��*_����iĎ}�R%���α)�66ޭsɯ���o��;Π��ln*Պ�IإCf]�x�ƚV��mVJ�]ل�o'璏[�i>��ß)��g@���Ӫ�1K�A�9%�Ӫ�>�Y���Z6��(�2����|�6�f�����3��Z6td`|�i��,�ul�^�'��1��/�5D:�z�:"ך~O��.{�{���F\����+ν��V����~�"3��6�l�ZĠ�ӭg�"�8�x6��\:җXCr��	ꘅ��S5����z>��!F+4i�	��c=:���������[��3q�X����3N�5�����u��o��|S�����D^�ȷz�v;��X�v��:�9G���U�w�5V`�:q]	҇d�����C�>׮�j��N�KսO{^3����w�#EA�hrE������h�(�D�mF��\/�Ev�ֻ9��1���u����V�"�!+���k5�_�댺�{Gm��g�����;)%�V�Y�c�o��N�U�%���҄;r��m�4%�Ck@���¶��W��r�{����3Ҳn˹���ɲ`�y䊎i�n
zL��p�D5��Cֱ�٧7�!ܺz��!��[��6�Wݐ�5:X԰>��yˀ��:��|tnmßY�7�vǹ~a�M���ů����b>�=���ۘ̾�Z��:V�pX���f,V�W����fz�Ow�w�6h��k��J?Ki���z��&�ϯצDz��%��n2����^5,�� �w�fw5���X�5�n0~a�qe."�2<��Ec��,�N$�m���9����M�Ym�o3�%��g���eOk���["î����q�g�it����*6�av9�	���R�ų���N�(y9c�&���eq}�x��MA�Ic>���2r��R���j�@�[e/����`���m��Lh�O�{ONT �2�<|
���/���N�����y\Er���d�]�� $$Whm�ʋ+W5ys��:��j��K=ߠ�=B���}�h+���?g��mnG5s���X�9�{�-Zh��z]2<7�ڇ���m(����eΨs���C`C7����VW-���s6�:W�[���^�ć�$�z4�k�]�Pg"�]��SϮb�+�`�ȔP��YѼq��q�i��.�=<�@�#�`̋�2��v^;���yNz����<'���)Z��[r��vm}�]1��đ��@�0O&[)����o��V�ü�G$�:�b�ɹ�9G٫��fq�?[ŀ�!ӠAʉe.k���X�\Je����n�y���ýr���ئg�xES�E�8ˇpOY,�$��K��I�ן]������ąY�^�Ma�r8ځ�1f}�`�a�ȃ�������0�̻0��h�;;Y�"���핳8_,,6ת��.b�׺ǌ��%rT!\��r�\0Ih�2����j�������d�M��@T�	��6=�nx��q�P�JIp��rX`�+�vm��Dn���=���FV���'��+->�Z��4��s��%�ZgFv�4}�P�a*|�_��.��wد3D76Xo=�9�)�#]�oP.�V����E� �Ǽ�]m��)w�9҂��Ƃ�����⿖<!�{}����) 5�zN@�ۖ�|�ɝ���e]����꒱S����]i	������53��یam��8v��]E�`Ѯ�E�m��u ��{����3y���7Jd�{�z�VZV6o$35�b�0Y�Œ������g�{I?sN�{E�z��ׂLҋ2S��wG�>�����_f����-/f�LƢѬY�L��k%^�yawcv���5�c�\���Cn�[��T����wP��R�dQ�؄A��}v�U�
TO-��q�Y[J�&K�[��v��kC�u�烹nM���]�}!�X��9��{δ�g���}��åeŇ_6d�h ��;h
p|c�����d�i�Iui����d�P���6��(`1�Q.@T��w#�R�I��y�5�q5�7�˘ˍ��x�:G*ZJ��3V �Y���e�'���u���7���h��%����t�B�.��*t��d=�Z�	���:���L�u�F="���*�nQ��x;�|E�rJ�.��8ɺ��Wb'77�S���q��u�Y���-\�k'G��ŃC��]�Ү^l����;��؆�$��Q�W��]}KP�B�WTD��}!��>�d�Yt$t|�;wd)m��1ܙD�yQ�Bp��t+����d6�ӧ��w.*�WqzU��2T���VӋ��U�`U9퓝��[�b��왙�:-����ׯ2�yo���Mf�t�܀(1��_�5wr�}������,�©��vZ�}lj��ɾ�e*9Ա�Ql�������x1r�\���T�AWt��t��l{	^�{��n�osh=kS���
ݞl\ѱ���.RB�l)��{�eţu(�ek����e>�ήҫ2f�J^�2*#ol���8AM���1(���˨XWh�dU�=�B`�����$bcaAl�w��=oS��P���A�ş���:X���� f��M���tǁ��z�T-뼚l�X.j���r�lab�ٚ��k�g@E��V6�7�~c[���A�7�wc�c�y9L�X�|����9m�����ep¥ޕ��9�"�`�];�^V^h�ʼT�y��|�t���%7�"��G%]�t��^�Vr4T�Y�%u�7;�PE�Ե�RV�P�`����S]3yb&�ic�xo�-�¯6�6JRY=�NR#%���ž3�,��qƧ������|����q���K[��^����@t�d��a�k�� �9_\����'���X�kYL�m�qk�1��޼����}}�'ŕ�sk�������x&��;RXI�ѻ$�dE�K�)Ӯ��;0+[�+p��dZA73im�M��-c�H�N�i��/v�o�͎��߂i�|H��Pm���!m�`����0�0�լD��#lR�jT��QL2(�ժ�0��0��0�"�U�kTU+0�fa�&1$��ÇU*E*��kڥIAB�RV�-�"��ȭ��,�j��aXkeii
��T*
P�h�A`��j

�������"�`�h�RQ��ib��V*�d�l���ҕ�E(Ȍ�ĭ(�E�!F�������(�!R�J�ڰ�J-���,m��h�b�eP��B��Te`�EQ`�P�Q�*��m���D�,�KUEYX(�$���߾7�ι����@��G��N�r��}���J�����~Q�#�K���kx��n�U�DGD���Yٴ��Su��j�Ỻ��u����5��8��`�*X�x�����R/f���v��ӏ���WvR+^�۳ϸ�5K�i����օ��P��*Ñ�
>���z���'c��R���}�o&3rٙN�->��`�w�\�x׍��Ƭ��z<�����P#K�Ό.GE�<�T+p��{�5
d8�S�������C��,2=uf��˱��t�8��޸&��*���}U\^�M}�jo�H�V:1Y��L�z�Dfƴ�����ʩBy�o
��m�CҨ*J$����\^�r��D�l'�J&_/E�V���i�����ǻ::�6���Qs�&��L��˧i���^Sn�<==��^�Og��̙;nr���x�.Չ��ۻ@�<��Ho�11���9lؗ_J(��&�'yr��{���{i�m{Ӓ6�����e3}=d�s�"N8�����D��Ov���3����m)�t6&/Eڧ�I�_���Ab�*b�p�邡�0�8�5+�S��p9b]Wl4��u�|�Vlg�u�6�����hx��eƲ�oU�)�c���֪Vv�ϞoM��{qM�}�U�#fkY,�4J3|XN��28-\�}���v�Czo7�.�ή߯��j�ǂVD�%4Ufn�0z
�D��[ǺWl��NpY���U�:VD;[�s��������0?Ev<p9F֌���S�h�V]�Oo�^���ᚻ�#$�^":̥�E$���Ϣ�(�e��.�����+���ɍ�;�ϯ�E*�Q��*��J��<�
�����b�e3�r�1g��ܱ�M7[�h���]E.���s�9vDdwR�� -�D���l�M��})���sƟ�w����V!�Rr���O�oK�ۮ-Ö���;x^N��g��E/�ۯ�,���.�8��1-z	w귚���xת�2J�t�lPx���鷲�Y��v�cOpx;�p�1�<��ʻ���	y�׻�W*�Գ�:�2Z��ݎ�9�M���=m���N<8���7OnM�=��u�HA�+��X�e-X�sl5"8<�$��33�r�O-���I����f�:|5�/)���]g }JxT�*�4;8�Ǧ�K��+� �לּy=۪��>�1�Q�3�kX&T<��!妃7�I���]�x�Ƹ��ޯ���-^��"` G �tm�x2�V֡u�۠�8�8.�8)PX7b�v��X��ks5Gs�>}�J��^z�+�~���iߐ�|[��%e6�9C��k��H��x���ol.��e`�,��ː���ofWbU_t� �h�]��ǏL��s��z�s'�0�`OX�'�ܼ�Q�)�.��-5��\C���y맘Q�^vil�����g%�3�6a0��<e����L�xܳD�:Q���
~�Ω�2��Χ��Ae��%���Qk�?-3Py�y�OT#.������d^o{|�8n^,����g=6��e-J���5�"��6���b�v%�)����a�������ױu�,]z=<���I����@�JE�����w_m�_z�ظ��J]BŮ��yXń����[��ost��q�P*s�$��8-%�Z<�~���s�n�n�_G�>�3k���v���<{�h����rP�bDC�B_
�+�-�r!�\��<���^�g�4v��/j���#0oL�y䊎|e��;�]%�R�ʣE�:�S�˾n�7^�۰��.�SY�u惢_�%�x?����5'�P�s 0�g�Dx��sn�z)dL0L��sj�w�76����KL�νI���3Y�U=��~}���Gc��y8�P�4�F\.Z����%ϰ��w1R���"9�!t"�@���o��ۋ�v4�Ve*V��k�C���Kv��m��Fn1n��\mv������{xx�zH�ƍҷ��."!��WN�k�q��7�vk���1���2���wJ��6���Ʒ$�����KI��y~�����X�h��WT�X�����0�"����%���'���dV�����R�^���@������S�&��MSem��м�`���P��0m��u:Syq�\��A���>�:�唎 ��ł���H0Ee]�;y{k�f�Ωo�S�k�Y��������޿_���Zj�ҝ�3�?Hy��
������Hqꂄ�6�Ğ�]��eΨp'/��({�L�x�5��R���g�d�x=��~��6E�Ԓ��搭z�9��b�}s0�Y�`��k}l�%�w}+d����c�뵨����2$3qݖ��4'�sk@2.3������^C�qq�����������@���@O&Z	���ҙ�ۄi�=xt�c/|Yu�yow��������M�:|����z�, �!�΁k*"F�ݥK����|*4���?�q����M�� S3ǽ�U1i��e�V��\�RJ3�Q��m��D�󬻩u{[������{uio�؟�ۙ�Z���a�Xk�ʉ�бM�ʘe��T��^����>t)��da򚶉1G���y����Wu*S��P���S�37�;m�W+R��V�S��q�ٮ�͛Η.����Zw��+כlSy�:���Z��I���+"�Ev�y�Vxg�vč�	]a�[\��a5j�3�k�b�>K����q��/��W�))%B�38��d�����oN��^�9�I}���32�ׯ,��{}{�I�|�\v�8;���\�%�	��ގ併��W0�p� 8��޾ �Qxi�U.&8)-���������z��[����O�h���"�y|�{�bC6��'��`��Խ#xlmH��{ې֋[�z��t�޶tA2�f⳥�v���ln�t�=���t�E�W��,j��Y�gWt��ؑܢ�ȃ�n��6&3��fe;�����+��?
�~v,J��a��Lt�𰌺��w�����Չ3�Bew�5S!�t�d>t���5�����~#���c^=��{g����J�ʭ/��Ih�O�[���#���.��B`.[���w.�,������Gc+Y�i4,��'��Z�����������~7�r�W5X�e�+�����5ɫm��P�P�胹�R�vgf��T7J�s+���t�������樄}ڂf�b���0�����U���g���`����+����G�	�|�`<b�b�����n�Sm��a�� �\T�^����W����:�;�\�C�Qh%�Ш1�F�ʞ����<�I�ٛRU��:���'歑���A�ya���<���be#��0�y��B�?V�Zm;��[�9̅�W����Z{N��P�����\���>�z[��O[9��L70�<�$��[J��kGu����4x����}ƃ��]�xT�5�K� �"�~X�L]�29��P�{(��6>�1�?��ħ�P��d3������Y�A��K��ǎ9F֍ΐ�W8S�|Y�/fͺ�K�ů����A����&#zE���
V�z�q�>ޗIXj\���-F�^��T�ݕ��t��o�/+yv����
y(���k�(�)g[�߈��Q�Li2�޿C<���>xJ��6�6:U�߸�׍TZ�2����L�>������Z��2�(=U�-8�+]@H��t"C�L�2*ժ��"���/������'������}OL�RL��ƺ�nX�X�鷲�X=6���cOZpxu%���ek�ŋK�IG��W������;u��m�ٕ���KQ�P��8�ald][8�[��;\��'{ �z����;���ݸ����.�����(�ƴ>V�Wof���.YΪl<#�mqE<�6����B�V�y�4S8<\r����g�swz\�����Of6	��l=���	�Z�y,A�m�貜��`dwrf�w9��ȸ�wس�1M��lg�aY��JU�ز�iX�v�{|a'�30S����j���M�Hk�l����ԈF{��YgŊ�K��g�y�..���ӉMH��S3�̬�.��Y�����s���::
ְL�{+-r��A�u'R��.�<s=rn<�K��h�L�ĚP�Zf�k�d�0���Lk�&R=*��t�	:C��wGй<_�K�+e���]�Q|��vW[K��f��L7��<p	���&z]#��D��c�/9Vʣ����g�W���t�D,�A�s��Zz�r�V��8��z����5�\�{=��z2r�ۤ�&�PƐ<G�Ma�~y�=���}�:���{
����<���:�j�B�j���`���y�Z^�P�˸z��K����amF���5�Eu��5�x0��{xvU�ظ�P*L#�Ier]N���wv�i�G��&ZOF�V-�~˽��#	T}+�w��w(XX���o���］k��^�3+�i˛XV�p�ÆX�2��)GC�ݷ]��"f�C9��rj�{5/t�_h��)`�V��αpa�}�v�{q��굽#��wk}7H�Pl�F`���EV�8$4��;J�!vJ��\)>[^���u4<��X����V!;�3�o������JǞH��Z`�pSԺQ>Ь�f�#�<͝	��e���xk���~��_�������z-���C�P�]��,U�9��:�<GO�����Ү�&p\pMk'�f�*u��Ep�6���<<�[>��J�/�pXײ�^Fi#$�/}��R��x=�o^KD,�C�7;���*a\F;x=�/c��۝��Ʀ�HD�����;���t��=��ռ�	�u��J��K��	��u"�*�����3d�a6��u��i�([3�þ���0Iq�\ڇVR8[�WKm���8�}�[*��X�Y�\���`�/W��n����l3��NX��u�����iْ���Z��R�luO7�A�)�}Pį索���:����h{`��ɘ�y�zMW����=��}io��*G&�.3~TG_�v�A��yv�1O>���a�|&s5�L�����<w���t�E�.�2
�Y����E4� �����6���N�;��eS��vR�-�������CD:�ڶc�[7�{���^�y�o'D�ĺ��C���{_{�:N���6���t��nGz�$��ռ֣�:v����1^�k��e"��
���A3,c�-����|d\Fޓ^�v�b���T}{�9>~�ױB.�"D�H��@mu2�P�f&�ߟ����GQ9�ҽ^�x63�Z�j��ޛ���>�3�L�hY���j%`R�>�L�j+����z������%���:K̻���%���S�u-[wIr�T��3����I>�O6ن�������4�'W��Y���Fܬ�?Ev�x8*�>������O�ޤѧ��}�)~�!T�b�/��T#/�e��b��b��%CC~�����sAA��j���ҹ�ɽ:���\&�1�M��˻¯���z̞����2�|�q�`Ů2;7�ڕ~���};���,x��/3ʥ��R[�����Ul����+�|��3i�ۛ 7���y��Ut��f�3��n�(oò��אy?e��M��w ��*���7�P��w�۳�?qW��aT�;�rݖ�1���l\���f��Ƒ�x�̧oiu���r�g��[�v��cS4+`=&XU֨Љ^�<R(�s�n8�!�ӻ��k\���]�:��{�sj�n�9;�b�ڵk������vP�&�t���=:	�B��p�(1^�����eHW*���K�uq\���A�E�n���֠��l��b���������~>8'�x��U[Ǻ��b�ɾ�3q���T�0
�u+
��`���ME�S!Ĝ��B�oW�j}�9��޴�Kή�;=ѐ��*��g�g�XN�e?0�� m�;��:1Y��E��|%�㗋zvZ��n~��^�$65� �A�¨T�R%ʋ�)W�.����H�LQ4<�ꙭ��#m���^M��ר�v������ZÃ`��a�֨�$�Lv)ԫ���:Ր�Pϓ�����,>\��.,�d]�A�ya��y�
j�R;v�x�|�5=\C�OC��Sٝ����6�z�O.Sn{�RƑ`I�����o�=����=d�ba�R���g���s�����D��|�
��6�TRX�)y���~X�������h��\-���^^�}� D/��]%�Z��2����8ɪ��Y�L��Wc�Y��/+�c�>���q�V#v'�C-$�${�\E$Κ9���Xs��t���ys��Ѻ`k�:�~kE��Մ̒��6):fEٵ���6�t����eoh
��}��v]�k�ؘ+�*X/���}�G$���`�W���_�.�I�K��I��V��P���{�gJ�3�eZ�k�X�0�Q���@����f;����T]mgf�U:�7\�+p����%|�8jSU}\Wsw�tStO>�s�ݼ��Z�����n-��u3�Nʹ��Y�-u�9s�8s+�*�}t��	�:��wR	8��sMS�N��rw��I]�Za;�o[$n�̀�[�`�2�:w��u�Yf�:7�����w������{k����~M�h��]��GI�]�G,��`�yM��ͩ3P����B���jcf��Y�v�n��û��M,�
PUy��aͬf��*�U ���C����.�*U����/�{��K0�a��\����
��,�E�x{�w�ɺh+Z�gPb8+��+v�*�8[��r��Q:�e�k3��Wxi7�<ʜ]�Z`U�G�]a��|f��<a�}ۘr�S{�����8�5~��& c\����8���Y�E���͕��W�S�j�6��ѹ�s�l>F�A�#���%�N\��V�а��9��#im�s*����	��-��b(�cK�˓���-J>�۱vEm<�h��]����.H÷v��pVV�o���Z֞���!�m�$7sN�Li	e�=�k��I�����G�e��9����6ֺ'Ւ�p�ۮ7�m����4G�	6��8�]�.�-�M�F92�ƺ�+���d��a˽Ox}osz�V���:v[7�x#17�?�K��.�fob��^nVКi��
�Z��f`�	����b�����\m-�༬x�Z�ma����qca�+��S(����}UٖR�]y�ȝ<�� wh�m5��f�HU��_>�ۊ��&<r慼E\����t��r�)o�͏�އ������(�8e��	�st�|��_1W�sb;���(�0\������/P��s���o�ciU�-�=�i�.[L�ƥlj��y[bI.Zf�Ao9��4z���MTbf�8u��nn��.u��	;[��x�H��w���\���o�Í�23�{R���XJ�3�0ݪ�9�ӧ�IіN��5�f�l�er����eoa������K,0�(��U��<l�h̜H�;B=���Im`d��l�G˗n�n�)j�q��e�J��Fݽ;�8ћy�Mt�5�#o�;Z��%է]}�����
�p�'G7���4�Q�D��C J��ῤ�u���&^�Z����Qi��j=�(��t��4�̥F�;��ζ�.v���� i�����i9z�x܀���̛����V"���y͖���>�t5�)
��h��W69n쑚}�%���ƶ����ee��Tj��Um)[h,",H�-B�J��[J�UV5��R���)Y[*�(��R�j
b��mZ�FШT��m**�j����h6������"�ZP��Tm�m-i[j�e���5j�ZYU�YmYZ�Z�A�BڌF��[+E�eKJ[e�EX�"�,F"*#DTmZR�+k�h[R�R�,F[B�YX2�icJKm��l�ŋR�aZ��R�IQ[E��D�l�b����Yj�Q�F�b(�m�����
��U���T��b*�P�B���J�V��V�mTXTP�#*TmZ��`�hԥV�dU��E`��)m���%F��6��*�#Y*J�ih ��
�b���EAE����VU�V҈��U��F��1�����z����U�����Lk0��67t�uj���&-�ݺ��Gή�	厧�JdW�"k̮*o5hDhrbR�V�_+�
=zp����Dh7%/+.��޴�7�O%��3Y���34��[��g�}Q�Թ{�^)�ItU��a*�1�\	�w�O�<�zאx8V�L�a8-�oR�*�g/z)�=�w��z�����{�P�W��(��q�8��r"���2�p��^rqI����OC{��C@Vx��D������ԙ�虀���e��zm�ݲƞ/�z���V����ɳ����O`�Ƴ#�u��d�l?vd����3�c��s0o���gk�OI�)�;���_[{�g9O����0U�R�0y�\�S�
�`^����N�f_u����{o���U��k��-���8���C�Yj/��ׅ/3����a���5V�����+�N)�zR���r��O ]G�Ύ����P�Yk����?rO�
T64Z�G.�v�#e^�.��&�������2��1=��﵊�g�)�v��i�ALj�!ו/e�7��^�0oU_]��v��^,���0�g�س-{r��AL��h�v�����>��֯��YķX.���϶��|����("���{E_��#��oW��Vny�J�C�7����g�L󕉼&�M������ �ă���\��}�x�����$N�س�fu^,�>CM1b�R��gV��b�l3���.|��=&ɛ)yx��qg�îc���i���r��1LP��U5w�gj��wW3:��<���P<4͎�@�J%滋�eȭ�6:m?
���S/ĚfL��>�k/{���}�]�|�]�Yϭ�œ���Αi_��y��=c��/>�����1���{y��(>��ǼWl�R�e�D�(K��@Fr4/�����T֐��HV$��g��l��wh3 r���k�2+0�U�N	>F!�U�&���Wy��3��;���&�^��F�w�*nu�O��o�邕�<�QϢ���=Kv��(��o�Rv,h��=�d�#���-,�rZah��}�û�F���Ab���xE��[K�U�iUG|��k&�f��d�| �<�TЯ�l���e�z�t�"��cf.����b��l��l�Ü����`z�;v�c�k��~����+�&�G��":t*c'��z��˪~�����L��{�Q�{�d���|f�����]��Uw"B|��,���U���opg-�='�eڷ�4�H_5AS)Ѭ�υ�y���j}m��C_-\��-�:�٭6ٜ�ZڽA1R0�py����-�Km\��Z��;HVu1��I�m:}�	��"��v:�f�Ⱥ�x ԥ�n3S4,w�\}W��κ˿?S|]=9E�7�y(�3�s0�v��zK��ru���G��M\H�!ͼ����oC{��W���B����P��a�t�r��9c�&�Wڶ_â康�s�gU�M��S���x��N��J�b��ܙ�hdc-�Mj�׎u�E㉋܊��-�YY�\�7�;(3s;��X�E�9�jlə��n��"5y�c�)����a�D��#���g=�ڷ7M��A��n�j�ԋ�+�� ������݇�0'�skw�k;����F5�U'�Us����^��v�������@mu2�3/)�7ޞ{�˙9��6e�n�� O׆z�f�j5�O��g���X�C��Ak5�K��o�����]b��~�3Ei��q(p=���X�e�eK^0E�8&\;��K0e`�����`���`���}v'+�m��Qk:Kx+"���
��0�:>x�(���Tf���)x���(v]g״���Yzu��7�
JĕV$�`�],w��Vk�.Ǎ�Ѿ]���z;CW��v��C1�&��sM3m��7ҷ��;-K����Ǜ��fڞ9K8gr9��S�y�a�R�)\j�!����hZ�*u�u� 3ws�;|t8�ͦ��>���t��{ػUYW���|�lO��/g�����ϷP���c��]h���@46r�K�ǽ��x��/�ZJ����+ñÞ:�>����X֥�:]do�u�gҵxi�U,���K~����7���|�e�(w��L���0�5�%X�I�zTkڻ�α0F]k.$�<9�U�K������3f!��?U1KC���o�(u_���g���+�i���ܛ7-[��6���O�g%����5���xN�0�/:��:�K`�`�܆��fe;������GP�T�8G�8�7�
��י�e���.ϸ�-/R�*�ԯ삅v�Rj,�C�uK�'��wϰą��w���Ia]�w^��k�0��m0�7	G�,�&��N����ZJ��]���ҙ.n�8jL[o�����Pѽ[�6lkXm����l4��N��2�>��S���u�G�\	=�\�3Æb�(�sӼ�{�C�Àlܰ	��_�Qh%�0m-�"����U;k����N�-3�oW�{p�xl�k瞽������.�����@�<C�U�����R�~�9Ow9r�-�Ѱ�ɦQPݮL'�uiM
�q<7�M�ƈ�*�+�(�v�t�Q�)e?���I�VfݫƲR�;oRzvu����S*Ʉ��*ΰ��� ����4�|,.w��Vm#Wb��h��y3���8ܔ�0��Z�(Ps+�B���/�ϸ�"	9��}=-�g���s ��a�UOէӭ��1���&JD�C8�$^�q��/5ڧ��0k��^y
�\��c�/5� �=�C����%��Ӝx	�����t�WT��W���9��>��r�LTɁ�
�~���Z5��ٻ+�7��f|�Z1��O
���I*�t�_�}R���*���Ϣ�,��<v�y��T�eM�e��?L󾤠����0t	)�ܔ����y޴�7�৕����ToB�{\��a�e�ݺfE�b��tU�J��1�\	�z"q��b`��k�<+|���i�|�P��SY�ʳ}KL���<1��ӳ��>�
8�Z,�OR�����oIʜx�W�i>�{S��w1��\�{���?fu�Y��d�Z�y�T�����Z�^�M�{��X�({O��Lo'���f��:��X��̌=lT}���	�Z�y.�E���9�&��А�Q�������8	&;lz�=���+�A�&Ǚ��s�`^��ǣ��g��{�uښ,��"�xC��@���{ wkD�1S� �>3H$O	���Kȅ>Fr���㕥�v�b�<]���`)]����'�<{5�C�]J�R�<��ں�^Zу�j9ڷ��r�ͨ���cY&m ���Gtү�e��m��{w�O|��W���<-���.=}Q����T\�C%qV�-�+.C�SmŮ���4�����`��E�;�.��g�^��T=�VZ����u'X�|,wG9�Ɨ	���/?]P�pl����3|6a2�i�����b�Y2��h�챋��;y�����_�k�(C����v;[Ɩ�,�v�&���2��J�ެ��1�4\gW*��ͣ���qH�f�����>�8��W�u�=\f���o��|�����F�S��/y�����&.��t�=�:Q+LƐ,��4!�������v����}�
�{��gŷY����!g.T�, �疁�ΑiX�P��w_m�;/��B����j.�b������8)���"�g|����P�	o-$(k5�]:�,�����������57��|�����wF`���*���!����!ەDCo	�1��y��[�buI�G�hwJ}K|���4�^D�i���J��EGVX6৩`ط�uxw��*p[!܀t�Tr����X���kR�a㆟�+i���b��}�ț.^�WцŅE���x,Er�+�ê�v,�i2�mc�r2��5���tz��[���f��F�l���׭Ț�d��u�P\)��}���9�z.5�:�9\���o�RE&/�7��Z`�9״��^���<��X����=ݵ��5oM����c�7���`������g�0Qν�I���5��஦Tc�|A}"���>�z&4��E�tZt���e�F�|�+\�zU\|�_{ˣܬȬ���nӗ�|^�&_��.���}�(��x��8��`��|�%���R�R8����w~�n̶�)�5gA�L�fg���;��=C>��V�뇖R8|�����}�x������:ߗy�j
�e@}�i�ZͰ̿�;���rǎM�����o���ʞ�G����z��Ʀ���Q��(q
;é����Y��`�� ��k��+eH�ｑ9�9\1�ə�eq�[J"�W�]Q}v�X>�j��1wu5��Ԅ��n�u5�O_nob�1�͂�"ĳCmݭG�,x����	�c�x�~C3��f����UӪ�Zޑ��r�6j�{޵�w[Ǳ{�v�}"J��5rP�u2�P\=�y��ڠ�*AKJ�U��H��愮�Ƀ(�]��
/��C��#l�<fs���o-/�6|�+,����E�w�r��}�J[�[;s���kj餆0dKFZ������0�h_��M����=������[����×"K�ۏ°��Ž0�j5�O����re;B���B�Y� �zk�;{o����h��~�(�"��;�҇�i��%�~S3ǽ�U1i��x	����Yp��-%�<�H���x�D�r�
M����o�9�ZΒ��9Yp�?'���z[y������m�OG�u�7Ƒ�#�#˭�������;�Ř7�
J�@��b
���ļӋ]d>��U��˃� 壦]T>Լ�"E�͜���&U�ޏYmy1�.
8�?u�?�{i(�,+�`�r��K���{�p��h���&�ʥϓ-�n̫�����=^�^��v׌�d�ȏ�����a+Ρ$k�oJ����α0o�ytH��l�y��b����hY�y^�#isW�00;/�bqYӟ=���M��ʆ�w�=g�|Ҽ�Eo�U6�*�$;O��x�[�0}]cU��Ȯ�v��6(���N�-!����w~:�o��9�0�}�a��w��x�i3V^Um��P�V2
�a���3��d8�S����/��M=Ҭ]V��u��GL��T:/� ۶"JŘF���&Զ�5}Eod��v��`��"���
���m���3T���ͽ}m���'�������k(�4�xz�`�����lmH6n��!�z���2�V"�E�+�Ey���X�l���p{�O����ș���Vn�i�V�k*��˖M}�jlw��,��H��޽�D��쭅����>P�$����g���P:�%�Y�uYh��͎�ف�w�qy�1>�V���k�;��9�~��s�J�`����Ĩ�!�В�5v��v�҉'��-�"���3᫗���?
��0:Z�Xx?G�9��be#��?=Wg��X�״�q�~�0�'�(7e��p;w5yM�u�RƑrs���OK~Y��gם��{������Fv&��I�D/�������QIc����~���kB:�y	���u�*N��/����T2�G�M$�I������Qj�Pg�B��b�.�5^���׹ccWc�:6�g�X��邡�2�N�Y�:�jg��aJ���wE���+�]����u�͎�+���x"�`����)y_���y޴�<Ģ�-�M{Z]t��P����������Kś��r�Zf4M�)�o���:���l�]}G�;�ӜH&���-�ω`r��d�e��$���BZ���K4�K���&�Я�a�+��I��.WEtS�Zy�|��r8���8�����ӢՈ0.P�G�/��s-��7�@���J��V�OG�^�p�j9G����#��WG��;nI������7իix�0V���>^"<�<t�uG�E�f'�`�����J�(]�ر���<}p�U{U�M��o�����֘{�=�:l=��̶�
��xv^�g���uG��s�v4�Z8:��>�%�d��a.yx:��=Aa� cn�Ef�6�ꂪ��fw���ݯE������kt���շ����ʞ�͏C,rX>�:�:ٻ�8��=a��ܺ���,�:f`�/�.\�胉��y�����VGMX��S*_�ߟ�۱���®H���_����f�K�E'7��oi��+Zȡ���Κp�	Ń揳�&����+W]V+���w��4�zT3ݳ	�=a߬�{ T���=�\Vփ����k;=5�;��u0(kA%��#���˱�:�4�j�fn�&��<reoz�m
�����{�-�Y�7۹Q��p��6Y�ht��Wm8��W��i��5ﺖ&ʽ�����MB=��o!�~Kծ���-��C����Li�M7�汿�$���$ I?��$��!$ I,	!I�HIO�BH@��	!I�HIO��$��H@�脐�$�$�	'`IKH@�|�$�܄��$�$$�	'�!$ I?�	!I�HIO�BH@�h���$���
�2����`���������>����� ��      �   @(  @�  �  U  >�j���-�ʲ�)�$�U�ڭ��AkM���4mmQ�۩][6��[4�ʚZ���{��V�Mf�U�e[Kmj�km�L�b�ƶ6�0̭�-�)(�&�k-jJ���{׆Vl��  �� D {օgw����f���Ji��8�n��h��z�g�� ���gz"��i�ܑ��7x �Gn��V��s[ۻ-�3I��w�;���ܯv��b��m��sע��=rk^��CKwk���m��"��)]� ��   ���   �Պ P �]�  (�([�: (  ۙ��zuͷ��4�˽+�A��E�U�� �r/e�Zݰ�me� t=��^�����
�n����ިT�;��(=u�:ݽ��{���p:P7� ){�i�Z����E]���Sx ޴֨��&�FȣB�ݵɡ���{t����ocDB�հ���z�ǫV�In��r�"ڕb��Kmw� �� 3��kj�һ��R�l(�� ��WXu�w��-���Ѷ̰�x wz@Ʈ�����5A�NML�5Z�Yl`4n���gkYm�lM��V�c� �9�@k5���ܒ�ةPw7m�@,��B��8U�HƓ�L1��F6< z���k�Uki`�چլ`���@�VP@����aJ�P6֍�x 	��M,�����Jfb�m0�u��6��4�
�e�C��ĭ|}     L*R)@ h    "��Q�&�    �L�J�SL       "���Th h      �$�@45����	�b"l�I��lJ�@M0�� 1Ǐ��C�n�ߧ.���e{i$2���P��/3ҭ+J��P���X%�j *�A�A�E�TT,	��"T,"�\Ra������g�~4~x�5���K��*(�h	��(��"&	.0D�PC('W�5�� ��ʹww|�QTT3�,K6��|�yL����UC����F��<�P��E�����k��
n�5���Kwrf���G;ם�c[���r��{h���źլ�����S�iOfr�)�i�,R��w*O��k�f�7u��>C�������kΨ�J�ր���FY�h��s��\O"-3���xs��Ի�ֽW���b��$r1�1�3��f��ac��!�51u��l(��M��T��vӝ��_4
/�UI�X�L
�R���(غ�Z�7�.��y>ũ��o=��k��w�R���yn�� :��m��ː�F���[�&Π�ŷz� ������3�#��	P���z,� ܉=X3������c(b�H\���u��U�Ýz ��Pj��ެ��znÊ�'h��������U�ǎ��x�t���ڻn���8����TTGz< ��%�<��������0����Eì
/� ������d��lɬ|�H�L���p��F�`u�E�b�ugTw������.rZ���N����<�v:k?`D7�0NVS��}0E�grQ�T�3�0����ܱh�5��\<�S�.�hW�6m��#k4�æ�	N�v#�pV{�nKya�M��f���h�6!t�<�g)��U�� �oť��<{�r��/.��j*8b���6�5Hy�P�ŅM�����{��u�{s��)9�&�^�j�E�ܺ^tt�bQ����zh�]�x�Und�uǺ$9� ���ѓ��Ø9ǎ��[�ݓ�ed=c��8��(`8������:f��wjf����2�ƵE�s�Z��t����k=�Ϻ}���w���g=�7$0iZ��y����p7
�ӆ2����ӼH�������������^���`B�I�bh�9ǹ�'�8��UT������������Pص���t�ܜ�$�׻�8�Lު%K���ಳ�K��6�>+{���4ӎ�˃D3ѭL�f>u�N]˒�����̛ns�8g�q����Xxn܏�A�^sTLh��x���ˡ
�t!w�ݹ#Q)�--qu{nSu�\��^p������Ik9Q�o%۱��&��������r%*8�dR!��646¹T{[�{7�<M`\SL�a�/:�ٮ�F�7J]	͟u!�i��f"�G��{��5��,���Ye�8/�����n��mŚ(@��.�{v[Ԥ��������g�	{6��B�
R�M�Ǫ3��ŵ�C I�����t?�Bs��C����\������;"��228��{j�J��,3Mٽ�)U�~l�]<�9�pl���l|T��[DY�G�:m��vpX��;!e-�5���xu��{o,��dֻ����p���bƳgXL<����^a����'y+�����!��\)� �)�hsq�缤Y"*mq'�{�����9����ǜ��i�1���(.�t��9�̀#�=x�x���9�V�+�L�)�! `R�˂.fq�ŋmS\2n��#N�S������mYzl��mr��|�-0�ӊ��a�{���8k�aq�T���r,g.�6�gI�m⒮/�=�35�LV���U�]Vu�w���+�Wҧ�tɅ�8��IH���	éf��qw �g5�]MR�|v[׬�Z$Lд�M
�A��|�N"�R�F���n&:��P���㯞��A3׆�A��Lr��1�T]Ů����m;չ9��c��
8;���T���ά���S��˒=����7����;f��k�p��m�����A�sF<��0p`���trn)��d��H�;:uۻ<���v��
7D����36��n�kZ
`!�ۙf��ާr�:60���7��V��306���𰶮G*�!e�fN��6�)�0���$܋D�Di�����Z����CXE-(������a���>'C思�n##��)WO�!�\ӓOW��<��F�kz����t,��pm�0��6]x��bi�U7a�eJõ.�w��S@�Cؤx��-3N��c;�@ף,�&���H��	T�n���$Z����D5rV��LG+��2�:��� [r`C��.1�C�����G}��B׫:���TZ4p�i��.��dէit��j����뺻�����T��J�ns+�x��m�o3���)�v��<�����,��8o'������wl�f�(�D�f���.}�RZ�q����`s�<��v-�	[i��v���\<�EA�"���L�s�H�hoGP�p���3�mN���v���vf�qX87�'ri�K��s����f��SF� "�u�lZ{�U��<n�׬�'J����+�f��t)�\���ǹ����/��\ +&_���T�zt��ȫ����R,�0F�M`�א��}���fn�����pa��[2�śr���n��@��pL�vs����;HB�DQ
k{�nB��ƻ�I�(ޥߖdM�ԉ>�-ndF�ᇡ*8�J�)�nY��|spu�3�a�NK���]�qd}vҞ��K��
[V�LX�dߦn��n� ����3�ޯ:l��c	�wT��bcz���6��w�M�V|6�����y[wgc�&ɨi�sH�&���ĨD�qA����BG�O�	7hВ���jZ�G�p§w}7��`|	���yEy�h��x4�H��4r}�z�o�k��7-������۹��Pw ���B'�q�n�����`�k����}�-{zje}�=�u3�w�c�8�V�f�� �QaM��[�Mz��� �h��Z����;�zMQ�ȕ���w:��u� �x���t�p(�u�R�+�]Lf$tVeY���s)$�ݐ�QU����t��)i�VQ��1�7�Au]Q:�v�|kRegf�����,؎�a��K���a81�<n@g���d"fՊ�q	s~�
�ky�MLaٸ�ޝX��pW� �s�a�X@pdr)�����8eM�����Lx��e���68�|�"����x�v�K�ql�a9��j9�A\a���a���^ż��ٕ��s����q��-�rc���y��z7jڑ������.���d�6W�x�#��錤�A��� ��m얌���5}�V�۶!2y��.�:�\��:�L%�I�+R��ˈL��ss��pb#��vds&��e�_b���׽:�����ª<�vGҌ��aL�[����~n
;|�}��ܮ,�ɧz]DQ���Ӳj緻����s�`{k hՌ�������2�.���:j�]����xh_P�H[��n�r=�R=7.��C:��r��f��	��]��N��q�����ԜC	�L�eܮ2�M (���v�ŷ-ˮ�6|��-�w39M�[��e�^_h2=�F�qǚA⤽˔=��X����ȷv.�>[�j�ĵ�w<�[�{�<{G`�g�ͭ���uL�r,��E�����)o�����N�j+4ɂC�������B��vVW'd]Ki���}M@YR�jTz �ۜ��d ��x�d��ޡ�*��fnh�ݛ�fm�F�����R=mu\�b�n⶚��0���eR��;� n�N�j�˰�s�z�w�����r0sC)�֮��,V1\S}�i��;���������b��ӇZpp�c���Ժ^6D�EC��pw]C�9,�V��J��XZ��n���h�xn�V�כY�6t�Q�rn�l�pYS��omr}V+�&v�c+B�M+�E����&<�a��[���sPzYJJ��ؘ�*<��}Ο�P�z��
��P��K�u��oqiv�y�=�Z����B�0�x6v�{(A
0.����f��y���;&�Ǧ7/LD��;�Ӊ�
:0a�_�N��Ǜ�{-��Xyfv�Bzh��>n���{�/od���@bo�Σ�R�	�wwN���!���r7�cB�(t�i�_=|k[����;*8�6z�I�8�sѴڱj8(r��_hX�G�H�0�FA�I��ί;:H�K4n�[`�8n��ޓe�E�����5���,�oX�e���:]�ɍ�seX�Ib��T�Û9v��ѫX�۝��8�{�����F�q����)�U���i��F��nmG�`�ec��\K���^��[V�����jLέ;�m�)��d.��n=7{!�>p�|+;���	�&��ĥ�&mO&E�;�c�6���QY"v�˲�u,se�*J���Eh���� ��5Ε{c�Fx�g�W���'�xG���0�9�l�ђA����;�m�� ʩ7����q��׫���S�i�&�o���7u��Q����ʦ]8���A�a����eM��
�\qR`�ۻ�dz�+&�DgWF!��`W��Lu�y��+�<���ؒ P���W��^S
lT�����)$���>]hv˓�C{ײZF�����q�H�4Gn�����Δ��S9a�7(5k!�u��mY�
V�=O�7�fK)�7����Eb�L��[�ܲ�q�@˕�bV����61�K��ĵxL�e���y:2�ݚ�����+��zf���O@��y���7�ܔM/e��g�=-�Ƶ����
ɏ*�Y+5D��.ɞ���u rx����t��G�,����C�K�0ѥD<�I�?���~y��b>�����<>c�r{.ֽ�J�H���r�ܶ^��u�]�^���ٵ�W�:[��� Qw�z������s���y{�O�a��kk�1�F��e?w���H�G���QtH�x�x[���X�!��W �����L���]�f2�k���o*�JKZ�4�͹e�s%�K&�j2�{[]7�:�V�[���9l=��:G�$��e��C5"D�ԁ�&dկ7(��޹��iI�ޭ��h�"׊����"�W��o^W.���d��\��
�_H:�+K�s�U���&�x�m�]�u�X�RQ�Hө;IH
w����ި,o�/[�^:a��gB�q%��f���WFK
�ηEe���/D�yP���}���KyH>�8$�^��wY�v|iqsw*c�Wu�\���gf	������-T�miff
ѝV��j�ُ�px	�,�@�s;JZ���7���r3&�6����=��ź
!��x$�0E-x��We(8���>+���mZj�9�PI�3f�̻L�`���]���=� ]�CQ��;���_�+:�n�l���10��q�W��v�v�Z9�4��DV�%F1��Ah�nv#D�٦-ꑭ=M�Q>�/6폚��̖H�j�[���w���Mg+dI�����V�7w7��p�1��2<bV
��rjt�m�[&,�=ZWK:��Dx( ��
�&b}ԏ��G��Pˉ�/�y������lh:|D��Mi}�����\�m�4&dV����뫙f-Yܢ����@S;o�B����N��g��"���o���K�ek��5`NK�1G�2K����Sx�Ӛ6�P�4sC�a�d�ط�y��yX�F��U�v�==qލ����ֺuտ���Gv�H�J�tt���̽��J�m>U{�6f3�����Haͤ�R�J6D׋C���f����s#A��h;|��HL�y|�%B���r�����U�̦ŖƂJ"�QB�Ռ4��ot�(��4W$�Jm�͜�g+[��`R�e]۫vз�&q�@9`{(�Zo{C������]���������u�j�\��o{���n_&w	����xY����Y)\�E�[�b��.]�o(Zw��Ń�>����|�[۶m�cVR�ќ(�1��`.�C�n����S�v"}����0gI����6�!LĨ��}p��(��]S`!K�x7����ʙ�g,���������)��J�±H1(�rʸ�3lK(X�kw9�	�}�j˃twej���c���% ���v��5���0q6�B%���ݾ[��r�9�>]�)�:�U�ͱҠun6�f�b��{�=6���Ӕ�-���I@c�X.�iN�ڷ\;��a���))dk\,8s��>U��Vhw�Dr�V#��⭳�$g�^����'�������jʰf�,��F�$1�D4����nR�u֎��Kqh3&�S�QNl�k�S}w� +.P<�^���;��(\sD��+��X"���x�vVڙ���:�)W��R��n�y�w�2�s�9�G���Ybh]���t�:KB橘J��Vo���tƺ�>H���:��2k� `|ݶ��A�*�ͻ�	��j�W�5@�r�Śf��=�kA�R�a��/�f�*՛[�]m0{�$��^�8��}v�m�tР��29k���}܏[o��X�K3��Q��*_[��k�fe�P�B�v��;���5RIہN��%�^"���t+n�N����%��ʯ����Wv���*���*]n�Mҫ{ĩg}mE�]3�X�u�`bU:����	�t�1�︴�]}�p{��5+�]��J��$�W#� ,��kw��n���WP���x��@|��	h��kt3Y]B�����s�ZJ�q����=Ϋ��6b���rT��P_]r��ͥX^�ԫh
-�0"+Fm
�eA���QY�ȭ=|�1��بvޢ~�!ՙ֐�0G�ʺ�P4p�p������K��9�ӹ��*�<-�o ��Ձ�+�^Ю�+����Li2���}�����}��V��<P~ejb�ʙ|�Wn��s�c]���p;���O��z�W���vj9��VPcʰ�ں����9l�N^���j��
U��j}��߹�����5wQ��Dr0<ҭ�њ�۾��*�ğ:\�(V���i6ls�ٝ!H���Wu�Mw,bG�"��/T�0!��rۧf�k��t�I
�F����p�thVb{'rݻ��tL��Q��JQ9���y����/�1p�t�hF�/9�����^N&|.3��r�um�D����d�L�M6I��W(q=��]��+B*s��!��kt#�)�a{t^�8����'D'��Neķ�"S|o�dˊ�dh�8�b��!f�@IJ�]�vdG6g�}sU^w%���;(��/���h.'��̏�;����b�q5�s�_A+��ڦnMp ��ϓ�	�2�s��##��V�
�`�$݁+fw>�����ɡ��E�x/�����r3��rdP9��R�7���x�q���wV�ҽ�8cd���(���_��)h����C�ڙ�ǗR���1wJ�ʹc������5�BU���3h��� x9�2�mp���;��a�&7�"�Hx�WN.:6�=���׌7Ϸm	������eDg�<�=�X鞞|5	��az����<�MA�Xqa�Q��� ���I�I�1�y{U�i@�{�9�^E��.h	�`U���&]�#_��gj�V5��OxC�{��<v��8֞>��]T~ڜՍm��)�m�7E0�����t&�"��w"� u�s�:���t�|���sJt�&��S�Թ�D)���\d*����F�قHN.���Z�>���F�h(��m\<6��%s�V$�H�W�nqbۻ���v�:_����o<c�u������L���O`�wroô��p�Rf0|q�Hu��G��6Ě\���rW*��r�q�s:�����3�W�y<݋�=.��z��Ǐ��|�q
���Űb���u`���{�����<N�GZ�y�*����B�I˷�kU�ϑ<�"�^�r��4Ơ,�\�-��A�r���W¯@�Q��.�T9x1^,��Q���Q���4�)�Ԯ/�`H�׾U�z�VHޘ�k�'S�Y��]��!a�c#]I5��z��4��"g��i�F�_8'5�zG���}ת���*�q-BFk]�t��f��X��U�Ι75t�7sL��=��ٌ?�N�Z������AQz�#���.������EQZQ�w�䖝
�2�	�s���Bu'+�Æ��Vn��
C�z��F�3�\�'��OЊ�>e������:�<�Z��m���gN8��b�K#m��i\��I�=�������f,�n�:zN�]WS�h��r ��
�#q��f���9	|�k=����%�9r�%B�<��8�E��q拭���y=�I�j^�y�R+����&�Xk���N��0�b<%�^1 ��I�-�u�Dvt\��Vn�
g{6%�:�Zѹ��[HR3�pZ�*#x˾�=�jڑ��j9�vxuoKkj[hT�7��S�n���??4ǧ�ڜo����	���3$�R7��>��V�d멪��խp��jX�
���C��٨��V�z�ֿ^����v�قH�v�d�nNd�5۠���6�NԟH�Q�2��]��-5��������ݕ��mc�pZh����+ �t�AY�)3�(��ۛ-��C���1�*
v�Y��,�Ǽ��X�Me����/��w�4�_����a)�Yȧ�f-O+B<yӔJ�wO?=g*�ýtz:�K]��0�݁q���0���}vu�/�;}��l>�R���L����vYns7��´�VڌtAs5:$"�2 ��o-�dt<61�1��S��TJ\QL��9b=�d�
U�X�^Yl�/X��А��ID蛒�|Lr�7Q�RU��K�RJU����ɉP�w:̊=ح).��͹V&�[��En�NQ���W�D��/�m��1݆��r��Mi�l�
�m�K
�P���$��D� P�<H�~�D�1#�M]��}�??VX@�e�,Q�,�#�yO��n�IujhH�|�L�v���nC�O��_U�*� �q_H�H����%Z��Lf]��9�r����k9�{IXp�p�v����)ۨ'X&=��Z��8�i��F��N���X3_'���6jf�³n
���.�f"WT���Cu*��tfޞ��9-@/9D�!�}TQa�%`A�r��!��l�lŜ�O:�1��"��2�y�oW�Hgj��>���H[�9����[8!��V�C���[�۶�X�V��'8v�N>���[�N> ����5���X�ޖj8�sr�'1!��|]`�+���Qu�v��*����7F�n>�vMaֽ橈l�ej�ʸ6�d�qXe�3K9��ĵ�u#ȇbH����_7gMM��U���{���o��/ie��&������Q��j��(f��\���VwJ��)=GVʛ�r��)�A934�	>ѵ��oj���GZMO����
�c�jG�`zAxdX*�<����aj[3���p������r��S�-��E��6IܟM(\Ґ�o|D\:6�\��Cb�'��y܀�2ı�r�V��gT�J��v�̦�@��؉�hE{��6���&k��b�x�]��� )�(`{tR�5���q�w#T��¯�#]���6��A���#ʼ�jrX�{�+jd↔2�wc�O��Ti8l����IZD�V;kkX���A��r2)�4�TZ��ǈb���͉��{c��2=�����Y�K�d�������.��60����w���pZ��-����3�'��g	ha�T&�d8��.p=Q#,J���ܿ���Zf����I�oN�1NaM84ӓJ��r�6�رKnX�߻m쑵PI����ĘR��A�ˈ���s����X8k"�ЧWڀ�뙹yaݣ2&Ќѭ�ۊ��u�w��K�);s<2�\yc�N�+���4a�D�fx7")�c��;ok�m��nc��7DZ8�N���$5tA�ώ��א�)F��)F�R���C�%��e��^>9��<�*ԤK�
^-h^5e���%��e�`-[׵�	�	�UĞ�b��N���b�qm*�2=v��06�����R�B�m���YLVL���w*�W�v�T�]��~�>�x�ǃ�4��nk^�>!{�$��!�}�X���ʎN��`�&t��F�*�`Ʋ��G�7](
�,�z�[aP5�t��]m�{���9iSY��\+<����O��ܚ7�L�6̆�W��N̈���.��uNѹ��vXB!�Ғ�g�+Ѧ�B��>b�B���nQZc��'ul��j]��ȏX�)r��w� �Z��2d����Q���ͮ//�*�kh(s��I���[��c뛨� @NPw�� ϯ]J{9�טi8�:qp �g4�3��M4�7���&�p{9�s˪V��ٖ������зt�i��Ze��mb�E�wn�m77Z����#��O'@���D:�����T���von����y�����<�5�F�U���X[��]LPɏ�"Č�ֶ��u�c���
�&��mZ��;���Aj�@SL�Ռ���s��X ��=�<&,IqG6g*W��N٣D��t�3�9U��w�8>�h"���7ޏ�^f'�Ź����̭�#�9���.���G9��h���t�Ӈ�b�vз�-�	X��x�n����O��GGY���E:{�Mk�h���+�
M嗪Ö�&
�~��q�j[�+>���D^;���W�Ч� ���ټ��3e0�3ٷg�d̨�hvܚx���M'���yaW�J��Q��a_��`Py���<c�����<�x2����7������,H��/QX�S�B�u:�7��ÝM�Ԏ��M�૟wJo�rʎU�r�R�������1rYB�άn�x�����V� �X�����@��;����)���:3�s��qS5`G�R�]��Q���C�2ܳ�/��u`�y+(�+ao᝹[�(uPW�L��{�n����y=��m�Lt�l���5��<�o��őM٤�%f����J�;ކ�Ӊ��vL1
 ���ފ�[_;��D��&�ml̩��b��[��A,��q�E��맾�|}5�t7�M��f�y��&�]KM�iˉ:U�-f�fi�wn����h$�f���yɁ�F�SR�2��g&\���@���G�t�[��nй�3fq����t��p�{R=�b��>��཭�@�v�"�t�9�U9wyE����g{'R�4�.Z]��=Z[�f�;�\8hM��!ub7WEm�����$����SDehF�o�7g5���%�iw��E�Duv�6�Ôs�e,��޽�g=�*=�&�M8��h�ViQS�*uN�)��H�hqp�N��r�~q��ۤ�j�s�]�u܁l�4��}�<&澺�>s#�9�w��s��^Q���<���cz���������ˎ���,�x���S�&��R�v&n�5G��0�Jz^�X\�w�7{�A�%��ӺD,ӵ���O��;C�c��^�(Q�^�������_.���<Z�� l�]��;����,e��!�54�\�q̾�*���b+옥C�6�uY9��9y@�!X�rq��Tk]���zp��5N�%=�p�U���i��o=s}��q顭��-|;4dʍ�����D��N�K�ޚ+pV=��{;7���. �0UZ�>��һW^��"���t����ޯy�s]�א��PBh=�Iw�c���j������M���G�����^�Ns��:�۳ۀ1���ܴ!�`�}��qX[�o���ݜ.��6��s�+1������E�ԳH7y��т�S�bG�9��
Ŷ[���ÌY��2�M��3�������YǢO�����g��O5��C.���wGw��Ly���M��Az^�޶�З�v�r����� @1���[�s��)�q�*�X�(],{��VU����.�rK�Iu���%�L�۲o����o[5������9�<�ppug�>�e-��V�0'�+�+���OkY{X��hA����ڭ�(�JR'؈�U����G��Mu���t{������^e�]��������x^���&9f���muv=�֎�\X6E$h�3��ў�;�v^�'����-VV2A���iXtm�����Sv��$�c[���Y�8g��7��І�]y��8���}�8;P>&�ސLӸ1oA.��rJX��cP��5˗7������qwZ_=,X�hS����\�mNaXf�]l�`�r�z_;��uӮr�ut�4iN(�=Hoe���b�H�[A9o����3o�d^.״{����|z���ܑ�ր����D6�#�W�7W;y[\5�e�'F;m����ϵ����W܄�]�PMsoϘb�8�_�ǅ�L<��Cd�gk��*�v�ISK7(��cX-'[OC	�yP�G1��I��O��e�;��a��d�m���z6�1��>2���@m�xz5�U\�X�}�xK�}V��^�~�G)�0S��2�^���*M����T=����Յ��Wס�>^�p �˂��ՍaJ&���l��Xv@��Ӯ�Y�)(��Y.��N�s�pB�Y��;��^��_����̲<v�z��5r�7�]֥&g��Nn�]-����U	ӕ�$�f�5.�n0��<����VCc����2�+�3%���E�sV"���E�JЯ:��ݞ�����%��=����:䯼�`&���{�JM���u�n:w7p�$7�h�z��2�'�"���J\�%ҼU�<��U��'0�ߘW�L�R�>1�p�*�7/`�g�վZy�c�f|u9�:
�`I������7���
��2Y�W��<hB5s�|=���[�n�'�}����� c�8\y9���e�d�]�@�����c�J2��:��\�`v�ww�dx��xt��Z1����ù�dz��A[3�٭22�u'Q|AS�|�^)y��^��=`ǩ�C{��6����Ce��|)��B�aB�q䢋Z7q�Y�[ƭ�8����,��A+y�mHb� �6��W��L�rs�N�\&k�ŌO�`��3MS�Y�����ڗ�$�4�<��J�����?^l���ߘ�v(R����>��<_e�fo�f�ۯ���W�,�Ǒ�󡶍7W]��Uەn^�VDƲ30�7uw3:*����F���B��]�X�8�;|}כ����7.�ڒL��{�=U�6v�v���=�*�]	��[=ޅ�}�f�r&T��-c�gV$���%�u$)-J���EQP�	�܆"XB'�8� �#�c�#�\	};������6n�M�6Cw��K��8�On�(����`@��ݲ`�����e�²;�q���lR�#��+;b4�;k�7΢1[���:�r���S;M�"�ڮ'/�N��Qe�l�v潡L����49uc����1[�,j�)��ț�[HQ����߉gۻ���р�J�L�mOw��\�n{������3���u��3X=:��w�z�V6�m��v^N�2
jK]��T�#���`;�0=�su���$ĸ��r�e>�WeVMJ�)��ú�&N3��uI�<9{\�rSwZy����d+�14]Ԗ��/�t�]]��}Pxw�է7J���<�sRO=�x)�9��w|���ݤ�#�j�rn���Z�][�f�`��Hv��h�Q� �GMj2��<��j�vB���x��>�����gki
ɘI%`�UKQL(���@� ����mQ���QT��˂�
%3+��l�d�5�X��L�0n�̭���iED��Ԥj���+DP�,b�iKj���X֍[�.F��B�R��(���l��*��5�kj�VԺ3�Z��E��ѩV-Ԫ�`�D�-�Z�[Q��Tt�\��QZ6�-F���SQ)�[Pn&9V�LL�(T���ҲіFҢ��TV�ƕ�[J1�Eˎ��Fځ�W"���j��֭�(��
QX�˕V�����e���`��-����~7��y��~˫�q�ܜm��J����R*k4|p�2��v1���g�IF�I>�ׇ�{��\ݿ�$�?�����?��LU�kcrq� /.`���+z��Sh��Y���*�s:�|�Aejc3ނF_�ϡu6ٞlf�d�1�ӟ>]i�*�<7Ƃ1�o�'��T^�μTmt�rP��7�Aޡ$����L��[���"x�S�v0lB���Ȼ���J��-y@}.��_M������P�*�R�Q�i�5�1�H�ۺ�̔�[Ch�����6*ni���!���'��8)M��z3����W�<J�/->&;�Q�x�76���[ܿ�C�s�=��=�*�6^��9��Z;?E�C����za�5
��F-�`n5MV��$���D�s�9K[f�azg7Vܢ5΃�j�yJ�u��S������Sz�Ws-EΨvDs�z���iP�~�tV%��h��3X[�h����7~�z�����?V���Z��p�푫x��l;����1AuNO�	f���gO��i$���e�ru�N�-��m	L�>��F��G�	O
i�Q�z�.P��w=5�W<�nsb�z˪�b�u��M��L�@�wa%��E���Im
k+mu'ֹ���:4��Keuvy��,G!hۗ�Ki��*�k5��|Ӏ�9� ˉ���U��f9�����܊�3W�6r�+��jk�kI�ϱK������zop}-P��^��}�QP9۽\W[>�
�i��\]�-�C4�b�E�Sk{0���s�&aeG u�~��HFks{Y����_v=���N�X�s�z:uLMSj�Ү-m=���FR����N�i?:�^���HNJ40�=Bׇ���S�7J��v�EŇʓ��S}�⫰n,���tT�� ���U����OELjs�okxM���tyҶc6��<��י��v'�8��r�]����t�9���y��ӼD���ղ)�e�l�mF98���J~ݥnD�@ͪ5�y��&�x����ڼw=K�2���.�ѳ�B���(Y�k,E:�>�N*J8S��U��@�e9y�ƻ�u��D.�}K�����כx;-6���q�{�Ly�zv$�m�.�ޓ(�x:��ӧo>}5�bC���U����mJ���tK�_6_[�u3�e�G �#�kͶ2�l�=.�p���"�1m��r���u�Y��&�i.����O� Ȥ�0TH��s-�sn4�LG�$�����pp��%pWԳ^�Tz�<�F��gԩ�`�HQ�۱>���qX��Z�I�ڷSV��4����Q�p�WvP^lZ��'�|��I�1�R0V�Ҥ�62��\�'x��Ŷ7���������H^x�����sL�\��i���o8U��u(0�i��c��i��������3۠�첥Wo.U��ӔQ���養Z��E��z�&��6�Yy-��)�J0Q�r�%�9}D��}�o�B��j���,��>~�;�|�%�dd�;>}=�1fs�Q��#zaϺe��M�T�Ԓ����M
��C�௮��:o � �R��Z���+
���k��M|MP�E
��w��JÛ�#��N��2�ys�&�&�ԭ�S��D@���	ɏe��h*���>ϊ6�3o{1����#�s�� ��ן�g�-7������N8�r�5M�7c���+�߹�7�T�#��@�0�D�r()����N�"���dj��b��)�n;8�;GTl��3g���SH�t��Kf=Y!���䘷�ߦ�a��BhH�{AW��	hB�Fʁ�cڕ{"����b=b����2<�B�#�V�oL��pI}*�&7'(nl��7��]��|{7u˥sE-�/Ng[ta�}�-�[׉N|`B�g;�O`X��!���=�� ^�`B̝ҹ$/�0#����P����GY��eh�5v�X-�<-Ve^�|ʝJv=ת�Q�8k@��Fd�N�YN:* MW%���F����ta'i���Ō�L_x7����w ��e�Q=��d3�L	驛��\���224��,���N� �S���x�ƌ��~��n�����A���rhU��b�Mu�#�	��*=�:�;f�3�&	��aSf�U>$������yGOZ��7T��4�C�3r�8i��J�"����Q�'�؈���.";��8OG�%Lt!�V��Y��6�OS�S��E:���u圜u�5�x��HQ��꧓`0�b����
���,���{G�ܿ�Q����Ǉ �K)Vb/fT��	�xyպ}e,k/��>"�Ixȵ���j�_V��S��KmZ%�Pm�W��[���X*n�2K/r!�Ij27'd<��qP`���F�(@n\X&��1��ˀ��ތ	����qhT캑AO�&�]�ӊ|��2 H��ۄ�vm'ġ�<�!�B��U�.����(b%�$�\��)����4+��}�s��[��s{1͙���)ڦ�T�a՟�+���
D��Ϫ��/%�S�fF����ʊ]��[��x���_R�zd���jw�+abk�9�.LvP�So(�U���R��>w�]��
�MeG���4��lw7�-�P�}v�T��"FO�Ƚ�����3���O0�<��VZ�Tx����^�P/���9u���4ԻV2B�I�$�W����Jy�a���e .8�==$ē	Pwj�^L]�����{S7kܖ�qb�����,���sL̴��2�U;׽˵P�p�G,2�`�gd�ܴ���v�F3"��*v!F�:�WS�aN�#F�x��ۖ���>�iTR󾮽����	��/dW���� ^�jr��!ў������Qٽ�-O��	
qODB�RcbI��"(.zƺ��%䠰ת2����JRlTt)�b'c������W'���0��;�z�ߦ`rP�FE�UjLz;f�^V�rp��u{g�����>��m��L�bY���|�@�]t��*z��"�+�$J�s�U� PS�v�<��$A�w�W7�;����o>���Jr�Twu9�5���r3�)2�2T����'�*���;@`�bL� �v�@���=MtP��{,9�>z���P�^�� Хc�����1�2�j�m��㞂�sN�vN��;�2`D��j���$���qP�fu]����H��YZ0\N�h���9�&l�jM�������u��U��C��4ܔ���(>6�	�M��@�
BRy�]k�n�w�{��i�X�@�����!���i'dA6��%�1�&d!�ꂷJ21��@tӴ�3w�KN
�9�T���:���
���	�dp����m�����rs��k�á)л թ�fk���xY���A�Z}�{�KO���>�0�>�E���ͪB�Ӿc��c6���b{��8ZM�0���j�(Ϭd�d	;Y�
	��¬젮x���I>�f�=�5A
���oh؀��ev|��Q�S"��]��hvD��J��#e�ِT��9�&��l��=�u�=���?�ϳ����=�9)��z�i������v�^��^9�Y�.� �C��3i�nH�T���@�5'/#3�4����E����ji鮗T����z�C�]���m!Y�%1F�9w)r� �t=(���f�r�l�NB��Ɋ�!Ȉ����}oyD��1�,t���.t�T��D��GPꍟZ��ؘ��iN.:^O���)���TZ�~���B7�L�N��R�"��29�C�,VY�7>ѓ[4:�QM!SS�p����#�'�8���T[�F�r/�:4"&�������@����~X�?Cm]K�'�i#Y<e���ǯ=�%�-�<�Z��{EB(jƂ� w�zF��s���`;�b���sǿ�˝����Y��q�Ç352U9�4S����ZR��%��fkT�t�_D��m��������p��t��׷�ZY�&0��;�/Z�{�(�7$@��6�����7����,p?����Q����.�������[��Wb��=��3u�z���K۳�¨�b;�w��	����&#_ry���VSe��X&uJ7k�{RvL:�v�8��9kc�g�k8VA吰�o�^�-t�yqq���Ƥ΂��z,�����ʺ[�\|�Z�L4��\����w�t���ݦ��q �Z�s`���zT�Θ��9\h���sp<�*��1\ӱq;���3Eo�s��#7�R�����=ۓcKn�A�:	�jV]q�G)M��A���j�3�Xx~�t�tə��tt�p]���{��
� ĭ�{2�v�5}��_}�����|���s�'p�XV��,Or�.����mJz��6�	]����]n��%#}����45e�NMgr���7�B9q�q���yQѸ������'��%:}���6v���Np{6ދ���{�R����-�S���A�b"k��w;n�}�!���J��<��'9M�ѻ�pc�����������́����� ��1y{+J��S�k}�{N,�b�nj�rZ����.zp�O%o�p��|����W�9oO]�����0T����*�� ��Ww36���츶a�Zċ^@�M-�<�^W{u�Bc�f�=)�H�#�̸to�Қ�9R�ڗ2�7�W�t�X���a,�2��D�b�u:7/E\Ժ:p�q7�,��S�FYٝ�n�n�j��&��P��br�)�q����ѹ�>�,	��z}�����:��g��N)��5���p��Wiٌ�yyz^"Wi���Ig!�x�/�{[	��]�%��Z蜫���ޠ�5Y\U ��e����wlÛm��L�Î��GWA�Mr�Rݥ�q,�V�lf�*·g��C�v07V��/L�Q�ܾ�k)E2Ԯ��͝]�N�4����$��iJ�K��籠W�j�}er��m��R"�ĸY*!l����1�R��iE�Z�-ekb*���؅�FҸш�AC-�++X�ielUDV4�X�-m�a�V*�UQr�F"�e��@���Z&Z�J"��p-�6�̫������(����Y��F+hQ2�U"0F*�*��E�ƵPDL�(**#V�F�3.m��m��h��j�-*(�#h���V"�R%B�*���X"
�4,H����B��#V֡VV�KjEY���%QQQ���Q�m��b"Th#Xe�����]���?w�߷���.�2���=�L{�:���ݴ�+�A&��0U划��}�B������EL@����vTnO@��$�bGt�r)u}J�HO�YI\H흁9�"$d�ȕ�����c��>��b��^��-K�Sp9��̇ �$uI"!�#��W��N�ߢ�>�x�U~��d5#*z:����2a��X�#h:B"s��ARץ7�~���Q���X��F�<ܸ�j`��y
U��q`�~�]7R(��P.x]�ӊ|�\t8R��d�g���t��x���ݺ�y�������r�����I)�8Dlz�F	qn}��^�t�|D����Cs���2cIZK���A_�H�!����K��&��������,�eO>�G�i����[�]����_R�Y���z}����?5�uz8u��p\*v�џ��;��-}=J{V�8����9�V��A������>A�[Oq�u�+A���;
U��q:�S������p�}�-��Ez��6��|���t;�e���}m��yE���f��*<w�^�"�O�'��.�w��B3�24�0�H����g��`����ט|�1���v�<[��5�!��>Ș�nb��}�J��U�;���6��X �,vu'���LT{�H�hh�3��g�Q7��"2w�s)��=����S[���s~�O7V�k�{�Sc�Չ�Ͷ�ػ����N3T�}�ZjZ�]ܹ�Y��g®�tr�+U��z<w��!��h[�UʁW4e􅒔�a�s=q*�xI��ӌ�~�y>@qС`�ϰx���f�+����X��&ۅyU��,�4lNH1l(���:-۱b�"_V���U%�3׆�]�Z\N�A�{�nu`ϛ�׳����-Xh��F������Vr�J��U��"#U�W']�Sw��s�C�,�x3W�L����;���;�9���sL��/*���3
z�W�ɏP�ŹQʍr��q�oSJnc���ߩK��#=�"F����V�G���3��w>s-JǸԂ.=w�R��H]�����x}m2�u;��=�1�"d^K
TZ��L>�{(G\H1�}9�1Î��.k5�C�v,L�N���Tիns�!^�6
�Ji�x4]�6��������B��cc�d8��C'�1�T���m�Ӽ��3�Aȩ�P00B3�#"��@ջQ��F쁁љ���FN^$�X�c&�� K�@t�����gEJ�Y�T[�ey�7r�m�EWh������jEX5jE�`*��P���@,a�m;�z}�t|F}��EF6�ϱx�;��9����(����	��k-���Wc
�*��D��K	�Zle]�Mu;)n��{'`�:���X���sԓ�Ѣ�씳���+1.�"Z���SΒ�.���"�5]�IN�}w��^�z�h���v�(FPUC�Ì��j:u�sQ��JX��f@�>p6-�b��0}̐5��í�醹��������1��*tc��~̃sN{�e�Ȟ���N�1�kճ�h�^�G�8ɐ]���p:�&�1WY,�T.{��P��{M�P"�ޑ&aȡ22ҵ$KJ��KjŌ���9�:.��G;��=t�]P���]B�1Z�R�����\��=�j���yz��̔�m��ޡ'��jޭ�J���H٘3��D�[�[u�r�G��V�oq#�T�$\׍�xt(
4L��J*4c��܎!�n�:�
�DCET��o�c�;ں됟��H�Oy�B�W���/�a�ծ�Ӵ"�h@�-)�t�M���T�TY��.��Ȯ~���z
�}��j}(���tbx��W.^���	��>�~�˾5h��Z�2�b�9%�}yu_����`�B���f|�tʞ�7�o�M�.�>�豂����ױ�f
���Ai��������2QJ���Cj<�_M�R*��l�V:�z��H1B�F3�(�[|��㰘ꋑ^�E�ʑNF�nyM���?���s����Y��d��g^ߢj���Nʋ��� 5#`wK�(ګ��g�t���xhP*�	��6}bD����Ð��.�ir�	�܋�P�lQ�r�̅�dl�p�&H�Bd8� ��X�A�ɝ�Ǥ�;�W>�P-ˎ�n�M�&O��P��!�LRy��"zf<�*$�F��c�uY 7.	����f����Α��ǞJ�s8�jEP��Q��Lp]�C��̸�+^�,<㻔k�ﾫ7H�+uѽgQ>0�So/<U����,�郳`���t���_���a�Ѵ(�TDk"�ؐkmNt{#&u����ɤ9�k�ӱ��Ρ�rOX���?3���]��ܞ�^&�'�S�o�3y���wy:��тzW�pVÏvz@2��V�Fx�w)���^�Ww2�Dj�Yg}�z���9n���9w�q�Ϻ9ׁ��\�a�et�Q@љ���<9�����7��~�"�r����.�v},A^�,�:4���)񍈋��κ5�b*r�U�K~!��;�5��9����!�4�:}^ޫ0:*-�ޔ��|�-xQ�
�w�W�\�yDE�*���Em�ľ\݇�+�G� �<���i�,���4���U�Fܸ�P���3C��Y~�6�xRQO3�,�=<�{�,�N�y{�I�]&.��i��ӫW5o��WVs[(;����3#����҇Fv2�[N/!	u��R.�ƛ����]���sjI�����=��z3o����#�DwO��S�S��M�]vOd��f������UcM?{� }��+<��C�E:��Ww.��lu�w'tv��o�����9Vi
���-]�eB$�����T�Δ�*�H��W��P����~��~�R�������a�SK���s�&%�#aC�3�}>���eD���pz�����Ƶ�ttU
T(0�}aɏP��<�A�o
I���,p�r��;�:LH��D�(ر2 �V�{�u�Y{���3�=�U����C��D�NLD��M`���*�a%��68�����DMP.\8� D=�F�V��S������h�}Wp�i�T��+�A0�l\��>� O[��HB��P�UM��|K�J\(�� \S�Sp�(dN�`l����&3��*cU\}1�=��I�,f�%D>�_cXj4�h�/�Fm�VnY���؛�T1����-U7�	��=%�]����J��h��N(y��������qG�b,~{�oQm��7�ߞC��A5.��8a� �0�V�)�ѕ�
��I���p⣸�dl�6GP�35R��W���{Ƕ6��Έ�(�z���vjԋ�35�}#hU_���鼵�����򽵂���͛�t��R�aW���`�=t0�!��<�V2�x���,8��G�)�*���n��,lMȆ����t���lS&��Ҝ�+�j��q��fw�r�m�C���R��k0�nٖ�W��/��_'֣i/��ĥ�S~3��~,8���8=wu�@��4]m<�9�S�dtTz�U�R�gl��w���2b�ޑ>�r7��w%������E~�ҬŇ.Ӄ�t\{���i�P��eWj�{�˰���\��3���i�vo.�6�^�����z�/&݋�br�P%K���?8��s���`�w�������t"�����N�R�}���K���G*B��x�+<�m��~�
ELÚ}>�C� 3;���;�T�L��h�gIe��K��K��#۴:�M��������7��޷V糹5["<��i�{f��z��8��;�q����5����yui�id��]Ј��P��Tߺ~�>���w黿u�v}�ݎ@|S��{꧊�۪WZ��h��(��X�7����i��(�k�eV�@�2�;��P0'��s;���ľ{���<N��]�yLv&��\�Oy��s�i��u�F�#�Rz�"��i��	�dWV
�t��(7��r��;5���z�ʔa�=�ߢ� V�J.��ZtpUz
hV���=~{���I��T]Cz\	Ρ�6�R%�28R��V�ۗW�x��y�Wk���.8���;������&a�/^�+az��Ād��w�Y�1{\�y��,�,^��d�a��LP7�/��b�}�fj�k�S�:�gP��  �RtF����(�����u�Ѻq3t�nz~�%�-:������� ���^O�ex�#*Ttt�lɇR,G���O� ^*/u�?!X��C���>�Sї?B_W��dT�œSw+�M>MD�b< �
e������묾����P֕�x��%���Ԓ������	��rb`ᔠd(-ft�_c%ƍ�b��P��l�{J���EW~9�.�f�?D�OR����w۩�=�7����r{g�8�,��һ:7����ᗷ�2.�31 WI���zEW
�P�9f'_s������st�����l��/�m��؈����:��n6y�2���t.^���L��+��}4)��߼=�uٲº���L͠�6��]�۴F*�)V��������]A���B�ѐ���y)Ҕ�ޝ���=�m	.Q��ܞ}�!�{���d���g�AK�R~a!�r�2�kyd���nl�P�GrA�휻���6�|1\ҭml��<׬He�Lm}�����^]m�y���U'<���ԫ�P2V��$и��b���W3m�7iE��ψ���2�X6��Wye��w���؈PS,���m.�����3�(�N�oe,��:�i�q�vR4���`��v�6<���;#J�uxDV�ݫ�mu��.�Ky�v1�t��rl�0{�%8���^�jr��>���^�(o�kur�s��j1X���=շ	Z��kl\�f�o����Ja�ϱLy����f�;qh@�w��2��+�,�Rܺ����)�-��k�(J��B�ݘءmnr櫖��Ҭ�n9ju�ۼ�(�����f5g3-]��e�ϕ�"�=�mn3hv�G��)R�5��d��_�>�����wڷ&v'�ů�s�I���^�<�vO=x8`�K;��wq�4>{�9�g�B�y؍�˥�����*GU9qJ�шx�U�����Z�����l��eKo�SJ�ڍ/�7��%J���S/q`����7%gp���rd�0����.Ό�4��s�O݊��׽�ۻȖ.�wS9����Ұ�\�ِ�X{Z |���s��+�ukJ4�l��R�ʰ5�A�dVp]XL��lAy��rÇ��v;�`V����	a-%d�R�ЎIY`�	 ��<���R�ḯ�cm"�]U�v�YW��R�qIKp��Ƭ�]�ԡ�>��w��e�.�j��Lx֝������eF�#@��嶨��Q�e���b]���$�զ��.Wl[J���4͙$-�+���5NDǋ��L��=M�2��Ye"cP)d-&a�_�Ky/�?��n=� *�Zʨ"�յʵb�QR" �ee��m��m*��e-���-(�(%h��*����� ��ZVĥ*%�fP�eTU�ذbE"��*b�DkYm�0��e��[j�*�\ˊ���$Ę�H��TDE""
�,Q�-��TQUb ��Db������*���J��Ub�m�,PLh��1QTEX���"�`�1���UQQLeL����X����`�	��1km���*"8�DE���1X9J��%_��~������^7�nzp�R/��[	�G�u�xD��6d��f.L��Eh���� �o���G�mz����E�W�9S��o�b��oi��\�������K��AD���0g�"b!9(]lV:���Ǩ��J䤨}&�3ʝ���ЭFf��*��w��Z�Ӎ��C���N���`~8�uv�2fq ��f���.T��x��y��g�2TR
�I�������hoۤ��S?]�iE8��i �u�?2u���a^�i1�d������������>Ŀ�����p�>QH(�'���a�Y�옐Y�<� (�4�aR�jÌ1�a��~٧��L@_�!���S<�3>��������~d�����c0��1��ϙ?sX��Y��,��O�3��a�y�xx�R�c��Y�VLd�*M}C,�������oq��i�$�l8���,���TXc
�ÌĂ���Z(��*k�?0+8�����%E �4g��t�gɦj�Rz}������3_o���Ğ���uJ�Xk�+ ���(u<a����T�ʬ=9t���StRbAC�-��La��5f�
C�g*�k���5�5�s�{�>��H,?0��'�~�|{M0�
���g�0�3l��y����Rh�d��[�r��1P��`bAer�CH
)0�a�ǀd�	�͚B�@ɚ��|ch�g`�m�GXM%\�ø������8q�̬1.G�n2~�[𕞉��'�61�\���A_T!֩Q����+Ixnՠ�f�/�J>��L�(����a�����ǩ�Ldݪ(z��`~�AgY>ϰ�(a�����R:�J���ԅ`V���ɞ��?s[�|�������O
��L@Qk�u�RT�l�kYm:�\I��vɉ���,1�O���i �z��(��6�^0+?~|���]������{Ώ�z�����A@�6�yHW�hx��)�d�x��>���A`k�
A˿,�'�>����LH,�S,PX��>���k��5��s�ޡ�*AO�@Ϭ�&0�����7f3��M�*H,��LO>s�����+�O}�Ă�Y+���yE ��l���*Ms��]~�~���>�=Vx�AH/ŧ������I�6²j{f$Xb�Xm�H)��)1�8Ɍ<Y���%|I�Ă�2~<���B���g<�=��9w��w��}�}'�u�n��T����{`g��C]�gĂ���Y�8���jAd�����V,Y�q�2c*N�Y��-�������k�;�sw��(��
��@Ă�L/�(���1 ��/�ɶM (�'��M$�!ܤP8��L;���~�1�I�!�R��Ry����<�Z�s��=�E����������a���$u��0�@Qd�ʇT��3;��LO>�l4�Xm�f�*��H<�*xɷ?Y�{߿�}��<���_��0�0�Ă�0��i���)�X��*����a�G������Y�|� (����l+~�ă�'��x��	��)Lu<�_e]0*��z��;�i6����톒+�{�+XW�Xj�Y�5�iUI�PĂ��ܩ�B�!�q4�P��Lf�u1�!9�s��_��R�{�t���gs{�C�;�[A���&�%A]��PL�q����VlC���O��O9[�d:��� Թ�iA]����d��S�ʃJflB@�ٸ*qv������"�4��Ăɉ�
A�?�Xi�8�a�+
��+3t=�i ��3�aP*AgY/(�V��CI��_SL�{��"����#����W__|�k�{2�uI��a�r��R8�n;�Èi ����0X,��fn����Ă�S�LH,3���+%eH<��L!5��?s�|g�ߞ{���}��凨�N���I�kt?2M�_�:��C\���i'��!�}��l��y�og'̬���30���
�@�,�c��ϩ�u%~O�3�!�m%|O2Ȥ|����VgSZAvZu��C_kYӘ��������4�R|yb�A����Vz��R�VVLCϩ1 �f��I!��+u8��
��Vk����gL�� L�3>�u�W�m�?7?R" +>�8�I�2��2T=�5�R��H;��1�aܤ�t1 ���~�u
�SϬ�:`�P���L�>�Q���6����u+$���(>�2uRT��ȡ���� �f0�4ì*A}�ͲVgl�� T�2�$�_��;HVa_?}����������d�IY��G��6=�{f$O�]�H6�����CI��a���C<ݘ�XV�AH9f���L6°հP�J��a�� ��%uܺ��5����ߞ}��~�$ߛ�����$;l��d�_7`bAC7a�I,�f0�6����Ă�0���{@Ă�=��H,�g��|>�\���o߸}/,��=N0�4R
N!Y��wRx�X~�N TO�ă�(���bAx��c<d�=���X�Ƥ9i)�a��5ߗ]����5�o|4R�������~[Zv���*T0��1���ȷ*���ΖJ_�d��4b�7Y+i曕1t���`���o��Ea�`D���<"o�=��wI����H,���I:���́��X)����c/��1 �h��*J���fP�J�Y*Aݝg����*����2U��k߳�y�^������)�
�� �C�غ�!Xm�5��Ă���&��>�(~�&$L��4�}�(Ê�H)�
ͳ�cϬ�R��}�}yy�������� ���C�<a��g�LC�+��?Ohx���CI�`T���'s�B�4���y?P�m��.��R
AL���I���{����zE�3���{f$i�Sϼ�R
g�f�wa��V,���wO
J�sT}�iE�>@�<2�$�d�=aR�����������}���g���T_X���bC��ծ�
�L>�z�R8�C�I:�N̋�`��h��ۣ톒e�3���'}�������~���ACi+�큉vjyܓ�0�<?PĂͤ���E8�]}`bAO�Xu��+'��i���c�g+�&��(
xDxn��v��+��?1����>�ǩ��
��3,�>C�E �ɯrH(��j���l+�C�+���M (��w�4�`V�{�����xLJ}qKE�8{W�|G��hz���%d��U �=��H=� c3��¤co�iE!��d�2�x�yd�Y���$�N��^�}�~��o���3�L@Qx�0���P�����n��m�`h�ư+6�SR�(�`T0�LH~�N��4���ֈ)�`�@����0"<>�K&���_V����m`�IR(L�Y��Ă�;d�|�*MNSH(T0�4�R��d���u%H,�=2����d��$����xg{��d��';z�Fо���3��	��ODoi�&X�ƛ�������a�)�ǶdWޞMM�ܲӕ��[���A�.�!��8�i��I���_}UT��|������6��!P�7V���O'�c+%z�ܧ- ��7a�4�ya�l1�U
���bAgY�f���=��
L�ՇXc!��ܽ������f����� �	t6=�@QC^w	��d���βs;�?n�aRZh�Y+ݘ��Y3vc�Hh?g4B��4��7dĂ�'���nk>���{�?{���N�(�}7Ld�*Au�j�X�G�a�$�������aS�
�큉�SF�4°��{f<`VbMn�E��?s�}�y�����-��=�ϩ
�����T������O\IԨ�+�a�`�P5�i��XbAVͪJ�TR �?t�p<"<���X� ˿������d�a_�`bAep��H
)Xg�i �3�²w7�1��c�O{�g���'﵂�R��'̩��~�i�
��}������}�3�R=f'��� (�'(z�I��a��O�bAB��ۦ�1E5��Lt��T��d�;�i���
����=d�������߹�s�~UH,?0�5�|�+3�φ�R)�d>ORq
��T��%b��q�$9�1��y�b,4§̚���ޯ�yu��o����� �O�s ���|��`Vm���wXAHr�[�g��`�aܤ����8�n$�Tsc��-
A�ӿ\�������ߏ�8���c�W=T���Ɉ�0�0�H,����d�C�
AOO�l�A9�~���߅������3���֑^������]t@B-�6��nh;��m% �1��r�<�d�ˤ�hy����vAہ��ٵy�:+'��]wǬ9�.OdVv�G��K�r���Arg��Wa����Wގ
���d\������]sd��d(�ٕb'c��^��_��~��	Qf���T��y(ȿ	��3� W,�0P�i}�|�՚8�w��&x������q����m'm�*�<�*�e���k�9� ��ٗ�JN\�9u�K��#:DN��o�Pz
l���9�4v�Y��{b�Cr�1B�q>��OQEE�tSm�����s�뷮�A{��/��H�U�{�)�b��L�4H衶�\���u��@M[��!;U�q��w%�f1�8:r��F~�_�"ǤYȝ�:�T1xk�s5۫���cf�T�d��)]u_�[x3���9Iq\�j�}�ʥu��6�yF���� i�G��C�.Y��p�^�i%�8�ˇpet�a��r���33�a�KC$+�����6�o��t���Ց���w��υa8��/�U��(Ž���WU�n���x{���z�m�Q�U鏅�.xFd����А��jԌ�3Q�x���I�-?o�G���%M@W��q^�J���AZ�w�k� ���n�����z
Ò���8}��V~��aвF/"�����l�[eF���D١N�ĩ¨�@�dе	Vc�o�r���>�>��,-��Ȼ��Y�:0	�BL�ƹ)�T�J��8��z�O)�'�;��:O�f	�}��"LM�w;� [���;l��(ɊqZ:��rL� <�R"��B:�(nO�GE����S��|a�ξ���P�Bd�Hbfל�iP�����J�N�=O�"�3�]�Z�6(;�?'��;�tf;���8�;ܚ��O%���0�!�5��n������r5��F�v	7����jV�2]�]6
��o[\[2ƾ����򰜨vm���R�t�wJ@���%��DO�� +9&�qQ�W�a���g�a�^�C4�� 1���!�Y4�N���:�Tt��;#`��(WJS}>���h��h𽫪���W�=u����9W��3��8^�ӣ	3)��{3&�i�M{F�@���$]���R�#��
dm�
���wa�n{՜�sB�C�DR�܎$@�
6#אuFt�@�{̵P0�dUȌ�红�T�#H�N�ߤE�)����W3��s��/���G�l_H���>U~�@���d�9�w�eV`��Ԋ6X5Э�0's�DP����G���@�8<h��ٺ��u(ph��@�; �}j��h26f��<�"mY�G�L�%�"�������R3�ok����I�X��=j�K��������L̉oQ�q��{���k5���#Q�Y]����yh���6Tm-����qH�q�V�����V/,А⫌�*�DF*�,�� v�"�q徭3ZU]�{�_ȳG��lܹ;����
�n�]:�o�T0�C����7TvlT�
}~r�\�^'EgFn�\�o�+4> ���AZ��f��w�-�>]P���g4];����N#L�'��8+b��� �ª��3O�el;޳�s�����F�@��
^�oGjD�g�Z�?fR���L<�ߏ���p������"���td�붸����f�W�v.R�y5/dC�#`��"�aX72�涩x�و�*/D�s�.T���]�n@".<�n��c�4��J(<�3P�FϢ�TA4|�k�����;9�������n���tI���#f��	��*V����B���çD� ���˛:�Ky=�{۸�gG�aK=����A;��u>�.�f�ȯ�8d��ִ��ҭ���)M�C�q���p��[}� =�(�S�aA�>**�W4+�~���\h��T[�J�v_Z|�*:g���d_�z:�ו*(t�R3��M@1O^pÜq���/� C�[�0��eu
R\�m{:|zC�S�Ĳ�����"�jX�Q4�LfH� �~�s�*��}AL�T�G{�-	U# �B�3�'b�H�׼����:�B�_���j��^kEOt<��A�)��NxȨ�#�lhR��W�	��F�	擘���ck�1R�T`!�G��nR�A�$p�b�B@��L�U���Ǫ	
o��w5
w�R�Ĉ�s\�7��j�o���Hb�'*��e
����Y�x��Q{t����k��
�;n�x�Y�x�i�ww�\��G�u�~�������$GNt�^V�)�Y]2���DWVU����4����l�bں����یAȇt;����Uudt���I���LS�sz�	�vEQXX��kq�u�WL+P��!]� &��r�:��r�f�d�Mx4�3D�o�U��e������{��4l�I_r��;�GAD�c���p������^�d6��� 5(�u*�b�a;��n%t��ڷ��ND�Ԡ����)�35h�H�Wm�٥q
�y��i�lm؉)�-���T�c�7(%%=�u(V=���3Mxu�5*3gbNv�u��|m(����,�j���A��ƽ�����OA���'�}�!W8��>{ʜw����u(�K�K�Z`�碵!V�Z��;˲r'�yS]�x�qp��}��-�L|1>,�;�V�X�=Z�$;�ɇ׬f�9�l�-ͮ���7C�E���Jn����72&Dă�S�0^[�(ov	�fJM^v��X[��:��Ny{׻6��$�p�a��c��I+q�6h�V셀��N��3�v֧Bs�-D�\�W�VR��iɜwkX��p�[���W��IHft�Ԅ��w1R4咽�{�r�-�ReZ�6�7��W�n�}V�Ή�x2m�.b��3F�j�(�H��-��uXf����_�ΐ���J�|QK��j���5�7�$�!`������������J�։���\5����H[���PI]�j8�;�Vfǽ��4̀��˷g6��j�lJ��8%ȗ�w((��h}���4w6hZ�rmWݹU�&f�2nl�V�x��}�q�zipl&�8�<A��w^+:�\�lٝO/��*{av�t��C���ab��ꁹ�v������OV��-'�z�G�v��)��ƹ"�ذN��k6Ep��
H"�g5���|$���u\��De���*�+J��0m�J��"��4V"�,EE��Z�(*�*��AV*������*)QPEF"�"���-��b�AQ�(�"�Q�����(��1�Lh���dAKJ
�EDKkX�E��#UF

�X�W�,c���EY�cb�"�Q�E��i�*1U1`�8�D2��Eb"�dEDEb�U�b(�B���U�.��)����,��m-U�����DD���"+"z"?r������lM���n��S�U�0mԤ�|tl�:Wn�T#���B�f9�� <�y>i�ȍ�č�W��^�F�E\�>� I�m�㱴lNmd����� (��(�{�����96���B��cbT�qw}NﴵG{���}�*���~ᢌ&��f�Z9�u��B\�
������eP�+�o/jG�V�rv>"��7��	��W	u=���-и��e����]�V�(��/[�yj�2�t�����>�@�$�z�&�^�QW#���tlEB������ ����Pޘs�qB����>����Y{�wde1�⃞��Mm�k��w�|k@��
.���.��*�|���lOMǹ�y��Dʉ��l�

H��Hu9��f:�y���r<��
��yV�Ð�o]z�׫���ȯ���*��s�^Xh�CEc�M�y�W�jt�-��ާ����n��3*�:\���)�]��9�����$��Q梨�9�.��G���J��~�}�{�}��m���d�M(F!@��P�(r��r/�DE<���<�r��������s��t]Ϝ��u+4l�k�Nm@q��0HtF���ϼ>�)]�F	{f�=��&�)����aS�����=ј��k)ǭZʻ�J8�E�7�{0e�CGJ��M��
�RD����G��/a-���X���"�C�B"F�C� i�|��4�`����.�~��)/��"�ܸ=��ZX�Zp������^�S4�ʷ���ma���ПP���g�����}j�j��]��>.��$��-�l	yW3FF�&\z"Ԇ�u�(d�6G#��be�Rcr��Q�2=P�Գ��P�զ�Q���DP>4�WU��0)f���*!�zA	hᓌ��mӼx3	w���yQz�T�g��nj|���q�R�]ӘE�4�*�y���nm�m�:����qJ�ĬX^K��S��b����5&���;?:�ګ��0N�EL@��]m8���*FV6Ӎ2G1#LґN���#zL	��(mz�K���#NL<Ǥ���:��q�B�=��`}j�!@06dJ��f<QOփ����q�'l�}#��+�Z���޳}tL)1YR��������T�zvF9�;j�K�{>ܴ$~E���2n����\�:�2�n��z���Jr�{z��nÛK��.v`waӬS�
���ȁ�֮�]T���j��h"���0ȧ���4��h��0�?r���F�/G��܏��ߔ��9���Ҁ9��O���b�of!91���B6�Οw������k�2$αTg�{W	�=Q(�G@3O���S�BWb��ìo�#�z�i�჎��R���^�v�1���5�L�2�K\�a7�����r�{9�r�y:���9��3�Z���d����{��=z�m��ڟ��*��^��ý�A뜦�����o'��I���0�~c�o��.���Ѭ�^�J��Ϯ�7 ,��څz��*O�9�<iA��ʾ�`~:"����c�}�u�Z�X�Y��6,@P�T�{c�B�}�������~����{u�����1���~���sSF���dڗK�vo�{3c&}��Y��{=��7�{bX�˫�v.!lǽȗ�
�7R���9�%�f�9g�
����Ÿ\�V@��X6cW���*��A�^˞�B��SDud�g*�<�dX
z.,s&�N�p��xH��@r`�u��*6��i*��:���c`�1թ�dTI�}1�.�Ͻ�o���lze���v�®^a��6c5�d#�\+"'8��P���њ)��jR�����6r��6�`��<M�{���㮴	�)�/�R;g� ����{^���E�{b�Ol��rt{p7mʁM���2qD,Wۉ�**m��I��:�R��JMGC�^!K��1"&�z1)ծdX���2!My������d���.���b��E9>t�M`��T�!G@��PF\8� D6rsl�ʣ�Z$�C �N$�>���$tm:&o%��9q�#.�./t�!���KR{:L���ʰ��%V͛g����pV߾]��8\��������qв�E,ѓ�7����}�c1M����[��V�S�4:�ٸ���G@�3�E�.2.�t�((��b���]���n����)uyX4%�5�=̞�w��[�!���B=|'� [���42k�2�r����54�Ȁ��B���c�k��o�7��ù����Y�D�2eZ����%^Ȥ���~�[����ՠ�iv'����;�A�n�Y�oE��dv�����z�m��}�
3�w��Б��
}S.=�p\Ч%Ϣ&����6�ʆ6E+w�]&�2:'�"v60S�� _��xl��U�QnvE���h�����⪈]��^}d]�}�#�|���0�'-�統�B�yV�Ð�uϭϻ��������5s�ih
���25�ҁW#�@q��Rm҇~;`�"�7�Ec��)l�/@؇#@��UC��\79�:.�>t#j�Ʋ�$�9���z����������r��=XȖtm=e���h��.G@�,Eӄf����NlHqсO���M8���Eў�?q�VL)K��#�F@S{�Vܺ����Ϝ%7$`�y�vo�"AF���v��r�և�[�=�盭X�p�Lu�G��j��V	�w�
�t�2�S�~����?���E�a�+��D5��'u7�}��W�����g�>�$t*eY��%�GmR���[T�� x5�������ww������^��Z���B�'�hF;�6�o|����t��'�sSS�ξ'��Xk��v��m�A����Wtx����q�\���i�����q<=���ٓ�(��ڿ���K۫��Yzl�"`h�CcmP�}�bzJT0@{;O�ۧ�&;O��
@a̹�x5W��:���M{g�f�ԅW���v�\(ŕ\fQA�+j�(������x�'��s#J���tXrVOG�%N�h֠Y��=Ǧ���iqqb�_� \�QNA�Z��>�^1A�������h����y�0�`���]����>�[Aĩ�P�]3�T�Im"�}9&2��50`��)p����H���Nj�~)u��o7���-59T�`
��Rve��5�ͼWN����wJ&G�W�G~,�[��{�r��r]�;��s:VsN�h)-�;ؤd�S:sp���D(t/���{��i%�[�>�ˀ�.��uc�XuN/�D	�讘���B�!+Y����f-���2��T�st݋
X���E��
�νxy���}5�a�*��b��s�o�(E��ne�������&������r�xEZn�g���T����&���R\'�
D�MW�I��j^�>��[��Ӫ�(����bL?m��W�U
plK�DK?`��3�nr�<�Nmu��`��&�I�3Pcћ^��sz'$��d^��L��<�,�F@�����hЮ�3["0mA�`��訶�Ck5��N�;�dtt�.d��t��eEG�	��B�k�����Ɖ��"��W��Ȱ��l�h�����R"��8����ݾ\
S�����U!���.�K��$"���wO���bY�[N�+���)ȩ�;�>*�c�eg,��4:���)�cY5L�0f����Xw�����M��͚O��j��9�Sc欹�:��`_=��7�WgsN4<���!é1�$���Ժd��>Ƴ��^�S�Wz�eA|�rR�d���Ù=�C���^D�0^�z�������S��;^u&()(l�"�U�0&'@4: Fũpb�X���B����X�s�Cb��bal�됢�}��s�D	4�AdVMV�Z����W�z�
-��P�O�z�w�&btd��m�$�*$F���H�؈f١B�7 lM�nZ4ct����X��$h��NOD�
�� �@��ˇ�F�5;��.EG�H6�߬T����?i��[l�!����&���"���w���D[.��(���L@ȷ&�\Hy��Wܢ���ˑS�JZ��\��u�rݢ��+�h`�U�oR;z͐���"p�X��ݕ�)e��]Ce�;���qݼr�T��xk� {պYM=�0�Pȵ��d�!{^�O���7��$�oF���m���ԃ2:q�|�^�ç8P���x�9Y*�OU�͂"�1��qG��QV�\p�̠b�W��C��Ӕ��$�4�W�/'�祔�����y|�7�\�<�p5OyulV��_�'���(���15c(�p}w����DU�k�g��l�����X�鼦=r+U�Xl�粖���]Ky5�^�]b����:�W�At�ʉ��Hڈv�����悡ڧ�T?:AѕO�Ok�V:���gQX�m��o�����7��+ް�T�B�-Ir��P�5�{��S�������]�����{E<tv��3װ�#�tXV��ڪw�vt�X��p�D��\9��'üMf��b�s�S:���̦iWd	E]�~ot�9�k�X��8��'m�x.J�ln̢)�!���Dbh����ћW�f V�ew8[��māxp�vp����8AH�ˆ���R0 ��K+�ͣ���Kݺ�7zyEv2��.���c��ǤIJ�B�ß/b��n���ogT���p��덝����
V)0]Mx�qRRV�]���l�ڇ�i+Tinw]v�&��Wa���E`�i����0�W� ����o�b�,/sZ{w�td;ލ0�+;҇xo��a��Ko9찥3�-�e�d8���_q}�3���O�nfVy�Pe a�t���͝k+�_0�֠{��8��5�w��y��[��\}D�Sn��l���@�������b�yn���VU�Xۛ���,}�nkm�K�WR �V�F<׵h�d��_�]P�i��6~�hk�c3�T�n.3r8V7���ҽ2,��B�������}�<�YB�u%ֺ̳�/R�!�F���5Wo>;R�$Ь�AbJpZQ&����\F��t׼�#�By�]'��.'|UbXqd��*�DaƷ��	���u�v���'u������"�[K��+��.��̮����wɝO7�.Y�.�Wn�T*�Z�����V��7��`kU�c�>��6���8)�\r�WVGd7��6GǮ��f�#bP����6��w��h�� sY�����a^�X�я5ժfXC{���n�����+v�c��N�I˛�9���m@;k��ܔ{E�z���w���s���X���(̻�������e_�����@Gs��|�D���x��)�r�ZY��ޏ\l��m��8S�z�1;{47�;T=7<�m���
��)�x��n�&���mC��d{kIP<R��[(;c�������#iaI{�#==#Цb QDm*�XȬEE�(�;lV"
��"1Dm��,U��(�(�j(�c�A��)IY`��FE�e���Q`����H�QD����[b��X�ĈQB�J(��#j�D����e�-�#r�E�X��eKiX�E"*�D*Kme��el�adDjJ���j���eV�[F�kj���5
�6���Z
1K���1���*�m����X�b�-b�\k�ڥ��PZ�ŶYm\���~׾q�~���w��m�T��|~8Q��cߎj�E)0�ؤLI��*V�������rm����1[P��.�8P�B�֛b����0ш9�0����\@�,t����@0�B��
W@��dR�̶5�R����$�F����-�\GJL؞�#�F@S{}���L�_���)���D�@�4ي��(�<)�{��ا(Ѫ� �^Q�h�T-��wQc�x$ǲ	b���2ӵ�=j��
LPBr�	\}��6<�dˏh��n9^q7j�`eS��"��A#F�A���e�
���b���R�S.=S6�7#}rD
�'dBK�jht1��y
=Q�Tт�u����T��]*��>\�
��T�S���כjݴ��c2ଥY���Y]+H�7�Nt!��\{`��	�Nw�^�v.��tM���I=7�	�gEb��˺	v0��'hN'$u�mں")W��Ƴ÷�£�P[\"�OoW2]�*�I��
���)�0˹�/�'h%le��S5�;h͑0�W�{�ÒG[o�>��R��A\���
�V�T��_��M�M���=wY�����b �w�~��VW�S44����I��-ɅR�p����	�ǎ�ܣX|̬�FNıl��g�}u�l�œSdxt�N�T�lT��ھ�o����hȱR�T�b�[�np)$ъ3b��Y��3Y�q.M �\lS�^c$��nA�k���Z�"��@�uz*�m���<�ix�f|`e@�T�ڜ����l1.��+[ھ�O鞏CB��ӓ2��^թ�u(���"�ڙ��:y ��zF��~v8VPtg�}�S����5=d���^S�.�ݏi�Y��,�כB��=t/ ��{����^��%y��	����n�Mͳ�>=ɳAT��׼o�O�`4�%���9�-J[��"B!���nI�+#�fJJ�5\��,�d#U����G]��d�Z��o:�k�P���{O.g�����DNO�VПl�5�6}=�LN���7J�ekm�̈́�߶�W@ݒ#c��XڰbT��n�T�[2���/�t�"=Dn*�����T�#�>����a�+���;K��)�J=�(T��ә�0MW�d�ō�{^U�],�=n*�����u2���e��g	nz�!9sB������v�Ǭ�����/�>����Mx��ԇ�����*�~�סgJ���E���M�c��i):(�L��q; v:��[hT�+�,�����ٸ��a�t�p�WA�;�a:��wQ�e�S�a�;VY�,�u^�
$�Q�۱0�\p�	͙�c�炑;f�鬽�� +���J�U� Pc\���ܛ��.��mu޸�VWG0t�M���BJ���r�/#�LL����\N�:Ÿb�{"���@��W�1��#��f�R�#�X�g���v�)}� ���&��t��
^��ٹ��{���
�vc5�=t����y�<{w�r�����Í��w}F����}C'0�ɳ|�%5q�@�ZՉ%_UԵN��O^��ZܙWe	u�ꉋ=�$�z^m�43l��t�(@��һ�p��ά�z�@�[�kI�7��ب�(��[�υ�>�b1�
�20	wb�[Z�?LbI��s�aVe���#xu=5,���	��^is+�t �
w���O��{�J��6B���\��I�#�ޖTI�2-��# ���Ez`b��.B��^��#-���C�y��,q�Ps��\`3�{d��Ck��6\{���w�4���D��z�����
����j��lOj�VQC_�nfZ���եg�ǄeM'��Իh]�HG	��C�Qi �+�`��+���j�E+������O3fn�����]���V�ޜ�+Xձ���̵�3߼ �k�m�F@0}�݋5�y>��㮂3�{k����{��;W�澎��������_G�_�c��,�r$>��y�߬�b'#j9UgSC�f�O������2
�5�(\��[4>�'�����	�78��SA�];z׏7)�����)��=u�׽���9�\��-]�� ҁB<#���
�Zn�Z��⼊��ϧ�:wwX�^���^�܊
X��BjA�;1��&��yԺ\�q�p!�Y�Z
�Y0��Cxz��u*�;t�G��x��ͭ�z��:C�uC9ъ���Iȿt�:4"'P�Д�)i���b=���\'� (N�o�'�G��9~K�� 0��	-�ЮN�İil�r*gcӢF9��yDݬ���+�ο/��f��T�!�i�"�d׫�9��~�3��6{���*(����_>F:Sm�k����]���9�8�%��=�6���5�ت�f���{Ԋd�衙7#�hс5�8�+M:>� (>πPW�>kŊ��qyԪ��&U-6�Pm\(�C ��Љ�F:���F�r,�c�p7)�̣i��p��-M��6o�j�0ʄv��D�������������W.��Pj�@&t9o�	�V/z�	�yj�⛩��"�^��f;��r����bu��Na�s�����N�^�=�6{��MZlp�7�]׮���,�8�Qwښ��NTt+
�$��R:��������>4/�C+AuXt��m��Tlw*��k�R����&*<9ˊ��%���j'コֳ���+p+��}8��ꛜ
D	4`�A���f�̄�H�E��tdS��C)@�ND��&��jX�}��]1.L!�lYFͪ�sq���Mn�ۗb��V���*#E�RXs
rI�v�[6cJm�H�Z���(Ԛ;-�J7P�f��FQ���Z�:�0�Lf���~x�[ɧ�;�� �P,^;p�uO{f!�0:4K�mO��Y{9��戆6FL�z4HQ*L�P����ҝ�w+:�>-��݌��>��߾"�e�y\���>g��3p)�b��)7]�c䋎��;+�7cG���� ��^fѠ�c�B�N\�±���q+�{_��� b��ۃ/�c�>�
���;!��/� �$�R�X�~�J��B<U{�	�ki���L!2�'9��B��,���p�������T�#�-�pڿ�a��Ē���m2�������.pT���]�ײkb�ˎ����ü�HvԚ+��<S��~�2(O��S= d���"��E��LĬ�WzIr�{���j�P-`v�u�륙��+¢�Ӌe/�'�O���.f��/8{@�=sG�i�PɨO3��e��Ku��N�Ի�t�*8�+���w��j5|I�<�Ub��.qέ�s�v)6wN�]+��| ���s��WH��3y��5"Þ�3�.d���:�u��ф`����ߺ..5�W�7멣7� �B27Z�bO!d��w��&T\ldϓWH1�[�0�\p�	��ϻ77�����b����Hɇ*�.Lz���s�^u895csi��J��>�w���ݴrn��d�������o�M�z=�H���t��i�84�ci�O,��3Q
����i��F���q|���`��
���W��*^QU鮣�A��Z��$"1���l��J_:�з`M{�=�#eҔ�Γ��<�Qo	d�*!C�].��u��jC��}f�˕�~_A��J����W6$d�Pbw�`dS�vfZ�i��暡Z��0�'���ۄR�\����=�ڬuk�7#2;)s��뎤� u�+�,�S�8�؛�		#�F����a�t[snI��qTE�V

]��B
S�� y��g����S; ���Yw�n��$���
r�6�7���A��թ�3�<p^����rd׎�-W�O�/��E"6�ϲ�W�W���`���У�/��#ֵ�'��"��p���>5��n�4�^}HK�uL�V=�4���1�����D&j��ɣ�j�!/-�+��D�C��v���Q�XG}t��b��ץ��2"0F�PT�ǭI��T�[��C�7�󣶎I���.�SJ��crk�������㦷�#b�#	C��\q�Ӏ�3�OIrk��W�|�* 0jo�ig�zf�1�ƲT�Zح��\l��g2��k/�)��b��-�-דc�`툣��,Tdl��g��SSĝ;��6��^�]�T�#Ǹ��u.n"|w�[G�Z���eN��ݾz��C�k��pa��������z�rv*�o�;B�Z!�߾��}"lG}�$D�4�m���BqF�+��^��n�m��sX�����Nm_>j����)�Xr[�ƶ�U��V�U�r6��ѻɞE��oXى�U��G=JE���lp=.��E�h������OAQ7Ӂ��X'�F�2:W����;FP�'K��(�u���	R*��9|e��Ъ�b���:˯=D��We.��{{4�p1��=�e�竸�v�fvy6N/oK�CU],��,F���|�@g��EeL;��q5�Z��t�2D�"�_u/��BW�Љφl˿�)�݂"�&���0��j�6����]MY5�U��(��X�#��4L��jA�ƥtd:+�1�ݑi)�7`{4;��RS��YǑ�����i�aq9O��%��8��'���ӯe$�^p)�:O���ɏ�<��IW���5j�.�N��j��\u�4��.��	�)� ��o����GS~�=]�OC�N�7��e�Y�����7h}���1S�N,�����(;}�v�Qz��Þ��v��z��p�~����s$4t�K�M+��K�R��*�O̗�H�x�o���,V�������^KD�r����[�:�m���
�|�����c�C9޷v[Q��n��5�#�N	ws�	X�<�_c�]����˴,7�\g��v6���ֻڊ�7R��iDq�f���ۘt�,iN�hXj�edR腌m[��^��8����Y?.�j&�ח���^�h�{��ֈ�mٙ�H��4����w��t`���{ďFx��+�������x��l�{p�����T��ˊ�R��B꼺奂�F�L��S~���v�y9͕��.C��d������T�vh�ɨ�������Κ�Nոw_�W.Ɋ�#���,�kfE ����<qv�~W�-w���%�F�{3����a餜��n�Ķnf��"�9��\���̗�n�d�
#�$�$ u�w۸���d�rȜ�|jW+2���J��oa�_��I�:�]
�5C��X�)T�s:�x�י�������}��:ƙT�E��гZ��u�Vw0��RJ��2M����(W=w}��e��z��y�ui)f��V��[�]�Z<-�v�� ���ФC�.	]Vo��'�QV�UE,\FZ�R{�<�F�1F�ZԶ��JР���Z ��UPU��EX�[am��UV,UT`�b�YX���`Ub�"��S2�Z�#R��(�1dQ���+" ���A2��1TT�
��W-�b�"(��UX���Z� ���EUJ¡P���b�EA�T�"�R,X)+
�b�("�F�����pb����AER �*��E`����DQAa����b(*��*��11(ł8�b"1X���V*�Q`��2
ց�U�8�UE �EH�U[k"�**��-�b�U@QE�����.��a�P�^l��T�+�I)�����p/�C����aKL*�+�b^����i�	~�r�3�}ZK�~��ä���'��ȸG������)�O���n_tw�mLn��8��Ѝ��R���=k��k��[5��"r��Z<_��!��AY��wb�Է@&u����Y�;�
 !۽�Aj�Xݡ�^�۳�-*���^�j�E�$i��X9��{jƺU�W�ʡ���P��BѡtaR��n}�B�J���{���:��i�-Q�tvf3�c*����z��+�|�P��(liSG�F�H�d��{y����ie��;���t)9��PmQ�*1��Ŭ��T㫔�F�	:���:�M����'�6��׭<����m�	��e�W,RGbsB�5d��8�pN�z������^ep��@bh��1Q2�T`�� io�������Ȭ�Oi.^}��<��^�9.)�O5[n3��8I��k��c�ʪ�y�Vv^��%�}@���D�����$V���Pq�I��):;O���Z��+��A�/�O���^Ix]]�p_:���o��ף'�6oED�d�BD���=�Ot�g-q�_��3���qiԜO�o���f�ҧ�Zg:�gI��2�L��[�z{�}l�B/�}uTE��{���%f�D�F��^Fi6���؞g���y�"��O6�:���Z5l�)��1^"P4r��c:z%��΢���U��_\w4F-�R<����9��
��n�m,�0M��ֲ����t��jaì��3g+�rM�mڧ �?xG�֛�W�o�މn�`s�aS��<:"2�j/���2&���5�W8���CP��P���>�Ѫt�e	���Y�i%�����zg��,>nt�ņ�7��g9�Y�3�u���1���nԨ*huD�`G=.���}dd@~���3	I�=��<N��Q��*}��|o��ɷ�9n#^�/!X�ׯ�U�$z�HЖ@�}�uճ��P��!֟�LD��ζ��<��?}���_t�=@4�;/�ax������(��ű$!�l\m����O�a6�!�b�P�K?�V��>~"�L)����L����-�zlϺ��������j/�~���N�ir;A�8��t%�`�H��3���,QČtF~{�{���Lt��n��q�ߗ�A+=��J���,������,��v�%`����ɾ�j�ȫ�}���ĭ1o�ƞ�O���4ä0y��:K.VH��w����-�bxĎ1����L ��W7�|�F	��X|c�5Z��O^��Z
z�������1�c��Er�G��OMv�-����l�3��oj��U������i��\��6�$X�Y���w�dݚQk�e�E�=�X+`ݿi��U�C�����x���D�b��1�W�ե��B2�KG��Ң�Ry���8V���M8}dYV�|kq-��r�؁�E;6�.�R����ƶ�1ҁ7Y�Dt�O�*��Rr���:T�2�x�����vޭ�s�5ړm����+d_�B���6D�NE��w�ڜ�-G��ͭusj�LҳAq����"���Sd�黣UuX���C�|X���e�`�����J����&̧+��a�$34�q�z�ou�suus��������Ú!7�b]����{�*uIk��9z	�Ϗ�����krHM��&dG*t�I�pSֺ�7k�D*�W�.%¡�0�#,C�E�x�ν��jn'EkT�iIz���ހ��V6�͆ښ����űTp���4@R��������ș��
!Ì]>�p9��=erbW+�ϝ�I���E(5c�o�,�ڈ���,d�v�+�Hj�ѕ�`EV�9����iy�-�SB��|�m��?hbUӕ����@�Z�Vq�����9��q{��8�M�u)nr�Z&Ї��)����1����.P��=��ڎfv�5;)���s�q�E���Ґ��Sws�Mg����[������Ne���^��,,��,��a���{/lR�A^��_h9��
�������cy>�]�v(d�n��U}W����s��/�r�#:'����<�:�8z��VΫ�l�CޟRum��U|�O����7�vA���iX��U�0�n��Ou��A��1R��Y�� qHU��L����2����IV�<�qY7k�d���\��w�(h�[%F��:��7\��h�{���+UVV��C&4�T��W}��orm��9�B����*�r̬k��J�����Y9ۤ���Z���	�Q�rC5B�������b���)��ɕ �p���緗���tz�t��o�.P�V
�j�+���k������nX��&K%���5
��sU��
g{�?'��*���M���9([�έu�����C�Hv�sVFfZj�k�)%u�̾v�yrs��'��_T~��۵��w��V�R2��E���i�3C�'{9�T�VU�Şج��Gx���d���Ʈ�*��(blM���V�e�e�0��D8m����^q?1���u(�t+OPq͋ɪ�B�ֱ��\���2����=�
��t(���y��S�R�8�Qe3{���9������p��B�<�bAk�e��y]��H�����Zĝ�ZT.e��O{eU"��@��J[M���Q_.�JY��6�5��g�������f�ת���clJ����Ie?���oa_���[6x�6K��#��И.:w��w{��*��Z��7��iBG�3���LyؙE�S����ֳ��|���H'ALCT�4�W��n\t�h�Ϫ����0���\�:;�^�nX'6`��h�;��y��;n�K�N�RCˉ=#G)J/[���6���&*;&�݅\���x3�˂��hc��RN{+��˛��c���T�m��4\efռ��i]8�������Ve�K��or>WX\)����6�2�'�w�+$�0�Y��Lp�u7�y��[�VOVdnb��i�\�ú��c:��C�fVJ;� Ow$V��s]��#%�iRI��TM�Z�s�=��:y�5�n��"w��>f�L�[f�.,�߱`��T�-cH�*��ҫ�����,��9�#�	u�8���7�K������r.1��E>��DH܀�	"Em=��9����D�'	�ѿ6u�����8!�FV+�v�<��^'�i��e>��V#xu�����{��s��S������t��Ē:��o������s���yN�{���6����Y"�,�n1k�^�ˌB]�f��C��O����od X��t�� D��6�#�4�0�{���W��Y���I%Q�����c���M���M�X������۲�Ά�m�ȶ���/B��G;�:��`?p�/zKkCf籜�L�6ҁ�<c��c^�h����ܡ3�a���u�EaA�?R�>���sc) i�L4�y���׵n�X�N�	"���j�N7�~Ey�{D����yDW�$�z{������8yQ!Kwޥ~��Om#i�#֑�g��z+M���*�z.\�u!�Q�!�E�{X��HX9'�7y�ƚ�J�����k��Ρ�������kӴh�?p�	�1�ig)��V(�T��	�c�6���з��+�p긞�&�\E���y3�؎��Ξ`>����[t1-QKY�˻��j�����sVo+�&%���.3zwS��c��Ʋ�2�U�� ���폣u�� [:i�M4:���j���K�1�1:�U���� ��X��|b��g��{����k�+VՖ�1)��mu�5�Υ.���M��S#k�%���C�
����VQ;Q]�u�]�Z�EM��S9"���������Y��o|[KKǽ�} ��#���4�����݅%X8��i�N|�%�ro�_7�*0\(p5}s/ai�>-���Ή�n_X�ޖ��� 5��&��B0����R��4�gC�,�fsEjm��:hOAW6��b��(^�3��;�٤�c�e�߻n��{���}��(^�nØ;j��X]D�D�c�_cRQS�a=�mM�8��WY�].�K��O��<i^:sm���^�;)�|d�^0��uR��R�k�jԾA�r���OV�ZY�����Y�=�E ��Q�ζ��MXi�∲+	s*�:�Au16���MS���D�űh[�O�IU�z3�3�c[�F�.b���Q�8�x� A]X��^��=�GN6kV�H���ש^���b]�(�J����&,���i�Y��� (��s��'/ĺ���&��X
�����V�,�[��7�����ˑ��)�`�8��A��7�ZɔN��g���I\���L7(�[j�vZw!|��]Jܵf�2,ە�ۀ���h~�;��9LO��4n���ü�n�YpL*�9�UF t&e�|������D�N���RL�n�T��Y[�Ѣ.�����A��rW�Z7N���Y�kX�E�칄�fjq��-e���(���'$�<�)��������
��E�Wv�DcEKJ""���DUQQD`�)ƥJ�R(
�,X��`�V
������2

�,��AE�1PX��"��+�lPY`,*��"��"��ciF �*���)d�H"�AHbV���Q�AF
�`)��E�H�"�"
"�J�+Qq�Uf)j���-�m�F�QKJ&YPX��JŶ�R,Qj��[mU"�KR�+P������E�,EdR(�Ȉ*��� �EA`�U~@����.b*��{�T��}��Ž.�Z*R[���e�Q�+g� �M��7�fW��D���D�Y�Ej�*(e�Ԡ�7wp;33�{3��<�Թd�DC�֬S�l�)�8o�NXA{��f����o��{��7[ؙQN����)���"���R�v���U�[���a�;jM��j}�\�5�N�c\�2�3�t��k��k��x�ј���]w ��R�)�Uxu�,J}i�P$��pـn�v\F�4��+f�C�7ک��d!`gD���s��Ÿ����`�~��T�v�-���R0��bhfQƹ65�N�U�sJ�����P�!��s�R*��dlΤ�k<��yn�E�^��ݨJ�`�駒��R�X }e�3Os�LXR�õ�(�\7�-
8`��\0l�CP��M��p*���N�ݒROڡ��q����MR�m!�m�}+�������]ߩA�K9|fd�T��T!�;�+��-�����\���2f�e���L���*=4E��}�k��֍ iZ�Љ��'Ed�+�b�rO�AϹP�2���e�v���8z�4�v7+�Ư���n��7R-m��E8�w|Iq��DHܡ/c���ҡ����V�����y�%��pc�E�
D�._�~K����
���<�$�Ug'��ĹW;�-	��xΞ^N��eN�N�X[}�;iB	I����d�o�b�ϫ��+�z�.c�]Y���|e��y�Q�v�d�"�n�u��5��	h���4����Z��!߆YnV�k��.Z�a���_k�Yl���P$t��J����E�ե�s��T
g�*O�L"�9�dM�X�0��`��4$)M��:���aј�"9j��@�A��7����[�ڜ���4���5 �B�嚔��wSsYv���yc��&��WfN��H���Hέ�����c5�_5���c+V��Oj��Mx���}��];Uט��d�&��nм�7�u�V:��w �^��/H�a
�ɝ�}�`���6u��Ӝ���YS�ou�qA���q��\n����JTڜ��^#�Fy<r�W�̬&����V�Ĩ#����N�h6�"��ٱ��oQSK���)�3"Z]��B
��\
�K�u˥�AV���%[�n��ؘ\.9�6z��+�'W]�^�:�4�W7kn���to��f̷6�$��C`��٘ׯh�qy&�1z�(׃;X�}D�#4jS�m��&А��	N�ȩ=b�W���,rɍC|��oWM¯c:��	��J�I�pZ�ֹf�sS;�V�rUo�tka��j�C"��Nˋ��;`ݛn��\eA��L����A�����9˻6f�jE��Y��"��'z'B�nUj�:���M�,���7�X��u20��d�$6�R�Z@ˊ�KE�Uc)��!$F��e�}�]�'������:L�e��+Rm#׺���Z��߇��S��4�jD1ZN+�շ���Db�nn��`�}�ڳa˜)���R�5��b|~�"��đ�s���^�K��Y=���6��\��q�k��"롌�k]9�bqP����iR���Dv�:��ORp�8F�pI�*n�f�; ��2[���=�Lvi�T��d���u��kmG.�zX|h�Zµv�����Ͳ���{���^޸�-A�p��!�=$�&j�FTڶy�\��s��d�,�U�EX}gT�kMy�Z���Ŏh)�W�HiU�=�+<���lK��M��e�������$�f�ם<�Ž��TΛ�J��L/@&{�>��e����t���c/���ygp��s+i-�*}�x�� Y�RM�M�V��%^�鏶�ˋ3=�=�Q��{�ڥ��Y|��l����˝���d��܌6�:dQ�kԙZb�a�r�:xk�vVJ�������ՌW�|6��/�lB3�w�n_(�������]bC��|�+��n�`�{2��S/{Ib6X䂾�&��u81�|����B����\�ekq�{��n5uy^��MW{Z�R���q.�.}%��C��G���ȟ�k�A�������*{�9�ixuD�NhJ�ۨ��-QhΧ���27y�ƪ�*�4#3kY^��=e	�ƹ��W��$��d��yJ���t1`��']�ۙ	>���T�7R�Gl�T�u���������
�Jmi��Q,kr�HP�W�id!le8q��]kW:�2I�a,��{���"���W�b����f+���*^ToPV%Zw�rᐸ��z�6����К��E{�!���xIM\�_0t��FF�bڗ/���P�%�U�O&�2�+����o�D�B��и,t�F�f�3��im]�5\�oP9��J	G���R�͢'��W6�7���L�I���l[�.��*.��&��Fߠd�j�H�h��I���Εc�F-�.���/KU>�c�Q�"5!Sf�Ua%U�]dIg����{C��u�KO�~b�e�nzn��!��jSFg��J��[��W��7;xv{��\�����@������O�*��KwggZ99�atb`�aldfN%�rG.#�y��0�!���z���l(�q��_JOz��Q|o��w�^�qή�2�vrg��&�k�܇��Dܔ�az�god�E��[ZT�1����`fr���L`*�n`^9�k%#K�|�i�v%�c�aj���>�mN���"l���s[��{�Ew����V2��z;�V_O8�����p�/x	�'�Qׅ4�+r�5RD��{���"�|�qs�gKՆ_'����t��CjUuE��șӭ�8^�N�nQ���)�w9*4�q����q��{��*}rb8<�gЮf�d�w]OQ��\X�y���7R�"��^'�zp`��Mۨ�g
�s��B1�N�d[V�o��N�h����sv���>�7y�P�v��n��SWb�������o��7��Qs8��3^݋K˃w��u)�XN`QJ�7ֹ�De��E��ndÕ]�[��/���y&0q�°l���}�n&(M�ƹ�=Lp5XG��BqD�D��3�Aʇ\�s+d���Q���^�<#P��&pt�oHyeb%�>�B*�_Z�[�F��:;.�Z�[S319�w{i�C}��hę'd�wŔ]��!�Y��Ne�ᶲ�v�Od�]ϖ�B��nm[�U� �Y瘥�Zr`�����c�^�sΕ�[f$G	59M����֮e$g.v�����]�E�M�z�ԟ�\��F�d9�������{8Q�ǝ�f�˫W�6���}:P���P�Qb{o�v
�mZ��L\�s����)No��u}Iwj�ÉI��/T\W�qk��W�3������j*�jw�jE>�d�*��8�b<��N,m�vt\p��gɎ�M,���L�$��j�?x�{�{[���|g���qx⁞mnqI�\Z����V6�/޲T�J��5���ڊl<.�u�k��|���I����r�z���~�W[�T�8�p|�H�:Ҟ�9���j1��܃<"m�ҽ���0aCP�+3[|T�1d�G��[t1��w8��$M*�����uoG�\Ԏ�"�5����G���z{�Z�A���F�bp��d<�2���������b�!.�;�ׁ�'��o���y���ц6o�FF_&�Y�^v�r�s1Yw--�FaL`��tr����&'v#R�]�5lz1�Vm���p�W8�;��ݔ���QD${X@�ݼ���5�ޱ���6X<�-{��]F�:{��,rx�!β��&+e�P��e3Z�u�D�.f��$w4ĆݭUZ[J�����|Es�3|Կu�r��M�}��O�=wQ�p*�U`�<�y����;����Nβۤ�/��#5e������ݚ��R���VL�c9{�(�6im7`�R�=��0���.�	�`=�b�����e]6b�̽|�f����f�ӕ�S�����w}�"Kۧ�ȍ-c�T��g ��� �v5�oa�q���77��X]�.{{/����+b.�5mT�w�i�t��.Jb��|�Q�0	���3qv˸�qh�y�Кg��`G ���n�g�m��c��,�-�U������vz�lU�'@�&���U��{ Pw:�*�'C����@3�١v�2�l�r���:�_G�JH��M`WZ&u�`�l����Y�6���/���#W��OJF�tJz��/x�w�8�Ձ��7@ܞ/яC��h����n��s87��o�K8⊧<�u�"����y�ܩ\�6�Q*̿�Ax�`}�����-v�=G���9��+�hљZ��XPwl=j]��P9t:W[�2����<��fK;*�ޅ�p�vy]tq��j�}Vg�wIМa@��V�:\��o75W^_+�z=�L���V��ux���;@�S��Z��p�L�����@T[�/��3l�hS[R�Sb��zn��j�sw�j�7�mY!]��oV�h�.M:�B=e�1��=U?sh�)�2�^��R=PJ|���K�����ǡ^k�s�����|�Z���ԥS&V,[�!E���@9�m+�Ҋۅ���s��t�,�q�ݭ�.���b�����fR2Ֆ��Vm��D�FZ�F����m-,QB��H�h�����h�-*F�EaV,PDX���5DkAQ�,BҦ4TQ�ƨ1X����"�DE�R�j����ȰUDDAb��ES-���"U�[m�DKJT��Z(�2آ��&V�,[J�DA����8�b*��X�iJ���-J�S-Qq���T��h�KX���2�PS
ZJ1U+3*�Rշ�Lj&Z[�QEҨ�� �-QL��j�ڢ����j�F��[B��j�K[b���-�jYT����[e"�۫�2zu@}v]*|̒�`��r);�h�r�J��˜�@�[o�s0�6��GNEp�{���,�<a���;����[L㞓�fV&���յD]�7yX8�X�Z��f�Z�wȵ�5�Ҟ��m�tkT�F�Z�uƭ��l^^$�q��v&�N��V_�����WF�����Ÿ��Խ��$nW�mxO	}"�SJ��"H"�RG�pSԯ�vuFD�Sm	o��#4�P��rS��Ք���Ϸ��X����F���֚b9�n}Kh�7Xշ�um����dDU�iL0+��B;��,[F�������7͠�n�;�_�c2p�o+}E�8���7��LuD]l����:��0���>eA��G��������D�%��$���r��ݭ���'�1��7�.�&'�3�+B!�Wr^V�M;0ȣ��g���1����m暎���T*��j��4r��ru��$g��Ym�c �~�Q��r��
�Jܐ�o�|W4�Rz��ӫ�>�#��1ǳf3��*NyZ�kq����X�7o/)=#r�m�Ҧ��j�K�^'�!�\Fk���v���7���0�����a>�%;���&�{LaJwm�{H���D���X��k���c`�VىF�5��B��5&�3�Xy7YLor�����a�UЦ�½�+*�$O9���ia�t�w�^�a���>#��3Z?ityMz�6����*��]�6��U��yv3�y
�U���5sV�oT{*��#����%�wE$�R�8b*����$�}����=	��r�LP|�_v�)R;��}d�C���i2�U}�}פ���R�����~̖0ޞ%V}�M��Md����Г��U�*��A����ހk�AG�^T��<Z��S�_T�څ�e��^�]��	����>�e
}����d������g�7b���N�Cy�vSI�%��b�-�+шh��&g�+ ������1�)�5i;r�}�ݎ@���͝s]u^^�J�cTKu\ fc3os2����2���v=[��knq�F6`��R�ƂY�q���.�3�W��l%2��]㡪/�TSD�A��Xԫ��&A�݊\	����6����u���!�u�C�vH����ٕ1X��9�3�5E��ĺ�[Z���r����S�Qႍ	T��oz�সf%��
��4�Y��	;�3��ow�IY����W#���Զ8aT��Ы��tvNdE�AW��(�c��3�!�!GY���J���1B��!�}�Md��B�V��m�K�j��P��(��rҳ������I�i�7��,R���q����@I/��c[���:����t��m�^�#�C����J�6�Gk���k�z�ɕ �,�Ƀ�u7��|�O�7����!�.������^ݯ]��C+�T(PR�$�u��׷�y{���]��{�~u�w�_M���f�Sy%ױ�=�6ea�����)��ƬdנԞ��Wv�"�AG�ፍ��D�-�����jȕ��uE#��p=+b��u6�}�72ު�\[J8Hah�Y�$q��WW����lE�YZ��Gz�;#k�X��Gn�\+�g{3|�Ey���z���D{�4����5�ww3�zF��}S��FV=�Fڮ��[�uV�_P�\�1����k�E�y��;T���]�<���c�����|w�2k�<xM>y�����D�yU�+r��p]/wn�µ�|��:��[�m��vkn������`jKo�~8N:�P=���3|i�����yk@}�r��t-�c�Yk�n�%+�]}�� en���mּ�Am�]d�<v3!jS�8`�o.)-�,o:��^�u��Ͼw�]�\G{D�U�5��[���QT�ě޽��Jؐ��9��;����=m���-�],�ƽ�Ԋr��	 ��lw��5B�o!�v�F�y�*2ؕ���cGj�X"m���m�f���^=���5b��Ѣ0(��1W�~��GqRx
}쭯FV)����ak=Q�)7�᝙g'˓��]��7����H�f r������7c������-����oJ��{���v�u��A���q�m�B�EG���K�hb���%��.C�D�X�����Ŝ�KB@� 3bV���1wIvޒ�񵙦tne�	��9(���iv+32�(�x�5;on�ºt��L��ʵ]�Qjz#��H��q]�cE9�����݂����@Ή1� ��U9�8W}�2�S<��S+��r"�	�{(W�v&w����Z`��I�h�da�c���ٖ����F��^o'�~��+kw��#��{]E�ܾ[yw����Z�p�I5��](�Z�:,�y��q��Ѷ�I>����31�N���ۃ��71�ݹ�XT��z<:�f�e�����t�E����Ψl�'�	�AoLv��0�Me�2�s�k�ZU�7`��!Q��>��L5~9IQ������[W]��M2'�=Ƣ�b�e��p�h��,U����]���y��,��^Z&.�}�yN�>��B �w�Ut�m�[�S�c2I'ޢ"�rV+-7+��#��p77���Ѝ��$�utګt�%�����N�q���h��#ⲇ�$j����V*�i�AL��J�1�k���9Q�ǫ��63B�hNe�ᶲq;<�si�-��g��F��h`�R�<�Ȼ�O�3�
��f���U�Vc8�^f^oӎv��Q�0�szH=ְ���v!�i�)�n�V�8��}������kf�y�p��e�-aOt�]���!�����<+�=��G4ixέ�Z��F:]C��I�)7>әlz�t��\Z%��#�{�ʽ�܍g\4z��[���\�0.�V��B�^<*�pI�Ԣ��\�;3��cy���*Q֥p��'���Z�u�+zk)G37|*��;�۔A5$_�ڟd�����o#f�������8�i�άmߗ��*nz�柦ߧ$�Trx�=�+]K}~L�@Z���L�3��t7�\��Dd�R�|+��'Gd���RFt0LhQ�w�FۥcD��*��d�\<!Tvs��<�:������Ӫ��v��;x�./��!�5�8q�L������qw��}��qz���E��1C���Q�dh!E�t˼���o���cݛ���PX�0�R��k�G��ɤ��x9P��b����Y�*=���[����%��}ӄ���-"����R�i�i`��+��0(�m{s�z�9����}���.�.�P[�l�����:�	E�,���h[N���SjI��Mʏ�ew����a|���Op�vQ��e�[��׆&��I�P>�O+G���-b��=9� �"eW��� �<���Tb��go���-)ڳ�d��vyj!Gldh@�Ok%h��8���<ΫN�k%��������X����p�s;��)�8H�u*��ʙ�Ĭ7�:�}3
#_njH�ј}�'jd>��b�8-B�#r�.:y�ij���0	�t��#!p�ݽ�2r�;5M6��V����8���\`+(�b��rN�S�U�%`�!j7�ӣ�ʒ�1t>yw}�:p=9q�m
����4��p�rז��uR���ebˑN�ƯNk�*4s���/^��vnri6��O���"��9�����!V�;j�CY�F���*}�vQ��ܵP|ns�Vk[u w6*���C�v�6����F��k���ta�g>U0��%�:h��i�vR�nݮ4���e%:U�����]fݸһW��[�K�b� ���c��$�zw��|�p������'�G��T7R�k��.Gq��8>ک�h���I�Š��c&@��*=V_H+#X�2��+�aزҲ����vN�u�hQW�3g�Q=�vt}5��xv�xŝN�?�����vwq��ݴ:���gG� �I�}Ft�1v���x'X¹��[��S-Ѡ6�dv��rr|hw�q��Zn��B��:�v@�pA��l��`N;2��׬Ŷ�vf�'���Ե��
<6sh��R��eF�V2�IT�j�V���ʇ�Wv|� �;��V�o��c���iM�9���Pf�r��g%�P�.][�_�ѕ��W�l�(��}f99.�sXڴ�ǏKݠ�O�!ͧq?vⷹ%�Ǫops��-y��_���ɯX���y�BER0;�{�Q�T��u��l����j� �#q���ʶ.�D!3ۃ����BNP�t40�ӟ�č����G١�Y������Ts^!���.���5G4t�an���#�����"�Ϸ�W�S*�JPL	wK	p��ѳ*![W�˰�����n��9��sd�q7���ۤ���fUB�=qf�6n�AzP�@ b�Q�Y���Q򳪋#W��8ga������K�̃bg�Ny��GY�ɼ=��Á���{&��(Ky(���T�������)ɸ���d�Y�7ܭX�*�Ĥ��}hn�kSR�ܾ�Y@���'qϧ;rܓ��FȤ�P�@ U
Z�i`����h�32�mص����j�ֹ�k*6�*ٌ�U�*5�1�8�J�Ѳł�T��F�ZѨ*��TF�
 �Ar�r�6��[R �ֵ��ی��K�����Z�ЪT��(�2��1*%m,Q1�3,X��T���[b�imZ0��0�Jµ�*[E��RU �TT-���-�����"�
�����"ʈԢ��ʪ�Q��"�(����3
�Da���c
�������k�3�ݯf=s��K�<�1�E��]B�Rj���rI�vn\�-竳�RHC��f���1ڇ%�OB#hT����j�%�1��ծY������]'a4�{�s�q�|�ba�uLnar��fK}�d�y��2�D�ٞ�n��=8��8���C+�0��z/%��j�^\���Sb���`����l��n�e��O.�f����:+(�
tI�{JΞ�ȗə�c%S�=�K���� e�v(od�g�~�bpR�:�8H�J�=d�s�ѫ)�+R���mA}F�o�ȳR����q�{�V巬�����F�����I4/��u���oc�Z�^C�ʎ.Cia�g^a���7�Խ'ۢ��;��Y��������"F���S�6�bM�R`Tm������+͈��VK62�J�\���uyQ��#���?7m�?���D�.lp3KYJ�ؖ_Q޷�[��k�I���R%�VZ-5�1�,�J��Ж�Ɏ08fL�Ș���}Ŵ�k�����2����h�����!������S���mɟQ5�[����7SZ��	�Ig`�֏�����z��*�o��ӝL����_CY�њj���Jr*�����$�غ�����]�y����P��#j/�1�Y��v�?e��Ľ�d�*.��`ר���9�Br��m	ܔ����#hg���s��<���j%��b���J�YQ�gS��8�){��5D�E���K}� �U�/	f���F���=]��o�[� S{�����bL5��eX�g�g9`e]�fs����rrI��u�h81�r���Rݩ>��T%w��sa���(H�5s>e��Nu��B��ђ���W�/��i��֩��v����;K�	1��7��!G�!��^���Ż�μ�w�L�3��Y8ݯ��y��`��_�Z��z�<���co���������q��L�\=3�	�����~�p�&8����'IA@c�Z7Ŝ���o+�\eb���YxO'Q��cz,h��ză<"m�h�����bO!�5
�g��0�½�ێ�wt۫K�Y#��\���R^i�mlb唜�t3�˨36�5eq��E5��O1�H�r��q�8mZ[+[�X�Au��.an�̠�Q�Y�9��Rf'N��Ԙe�>�K+���{T��M��{'%-���!c�xZ��ߧ��c�z��b����7��0f�d��-{]��t�՜*S�<`@�ǫ9F�vZ�f��y�U��q��EM��s��M��6���6�{����A3Vs��]b� �B�S��AX �c{��Lg
^�Rb����ں���M�^3�ԡ�3���.�S'#���xyB��#"t'��y���iiĉ�e:�h~%^���{Y����\��W�c�(��f�~��{M'��o����#�1M��f��n�e?^�9�X����h�ʘ��4�K�>�nms
��H�YJ��=�P>X��nM���H����E&��`[8d��jQԟ\����V;0JB�칀�J���M�}`�L�.��{ٞ��F��|��2�,�tI�o�t���Bf��5S�%>i*�zyl�N�c�`�\jB�yS�;�ml	��6^����BF(��::��r�iL.v~Rӣ���7Ve)�I��zi�cb���i����ەZ1��/�&�Wc4�t�D?5Z-�3��]�����F	� ��ő��.rcޖ��]Q��n�*ݡy8�,���it쪱�f�F��1�)��
"�9A��Ȩ)�T4�cdL���}����5+30�]�rL}�E����Ǫ��ɚ۾=gٔ�d�ʮ�`oڭJ��A����ElHY��hU��K{��wc�<:�p��glg5�y�Ao��h9T��o*����Mο#�39����z�������'(<|߷�t#�L�J"�o��:a���O��r�:ȇ�x���zm�+�g�4.�&�&�$�%
<H��{��o<�L�J�0M�t��J����êN�6��O?J���Z�-��#�H!������9��оv1����8q�#�;�3aEr����1�ԇ ����a�ڄ3P���F�ʺʓy�̴64���n_(��-������
��$��Ƹm��g�����G޲(�R�v��H�tJhyjχ��AE��{��5�\�:����\�%:�xh�Qǎ-�p==ϑm@�]�����v���n�LJ�6����(ky�f��W`>}t�^5q�ث�,>'j�%�TT)r5&<����r{^�k��%�5d��^js,)�
�4��8�ֶ�H��[k�5�QH�8o�q��]ȧ�'��e���2���:]*�iZ��ؾ��.:(SB\d�'�s�1nrz{bث������K[���
#�t%V��^��Ln�r�w�����+�0�xܰ%�p�V�U��ѝ3�����6z���<]p��2F�Dl5Yb��o"ލ|}�en8���%��5p3��o��-�HK������T�6�9�1�hN���h
�����)�ջx�Ac�W��:2�rފ>W-*���ul�u8Yk0qē��;cm�Ԛ���u�F?���xE��҆�.V�fsYws��M�.{~�]0p�Wy�����}>����T��a0�Ȁ�3J�Z7�����S���o7DH��'D-��M��*�e'|_ʛǡ3a� j�Q;�4r�*m�uF%sB��^j+ad�ۜ��� By-Q�tΎ���+Ӎ�E�ޚ˶(�W�{.�]'a5�[Q;��ezz�W��bf=�>TC��^r�Iwy{�)/?i���0%B]E�o���[�k�����Zڄ�Z���`=C�O�YQOk���E���ML����m+�'�P���;�~9W�iy�y�GC�:�N��䢻�~���[Os��t7wO�b���y3��nT�lͶ�.t��5��#	�Y�F�w7��p���\y�HIb��p򴼃�H�
dqU7(K�x>�(Q�ϻ�����MoEu,GŽb^3y�:��'�W����LQcW�42�}�m�}un�X���͌�����*:�e�뤕����];�p�m��YSY���$��f����m錍����9�6�˵��>����8!���0�&���X�*86��Z��b�F���`�`�w�g�o�s�O�P��<ɉAK����g�f��T�5�QK���I������#Ԁt���g�x¼��i����j�C�^�z��Vg�q�,��x�>9�;���aE�\9^b��Y�'"��J�f.q�#��WC3�(��cKq�Ԭ�K�.�{��ܸE�	mG2�=��x׻�R���ޑ����\��m5F�'�g�f(]��F�΋k.��9O��x���K��>�:/�B�GT��i����o��Xz�+���c��P�8cM�\�a�sX��gW��'g$�\g'޽�]=&��.�"Ӕ&�iϑ}y�3��wy\T6b��.n�k
{��D��jHgs�5�?z1V���[��)��ڋp�5#F�"D)�ǥe�N6�W'Uv�l��N�t��ă����*YR2s9�{N�)���3��u�m��5�~
�t�ȍY�?G\��;r�A޹���խ�##G�
����,u�w2�C��\��\��b}���Ul�K6��O�!��쁼n��7����.N��tK݇t�����ud��t�m�VK�oE��y��&8e�A�f�^���"=�m}�Tzñ�����&Ԯ�3�qp�8Ns�\^���0{ü��}�ױ�`�8wi�P�\��hۮ|��3��J�ֶP��ۘbÛ������KE32�\�Kjn��e��YD���y�TO�\�V�Kmm�}W�nKz{%��U��݅.,�iZ����MC��ΓoB�R���b��h,���Gpnd������� ܡhujxXjn�h0�`U�7h�1�f������7���+�����
﬷�ÛO!���+^
9/����׼]6�v�ue+�cK}Nl��yz-%:d�5, ����w7�����+�c��z�:ʍ)��ױ�cy���5��\��J��[.M[|c�:$uF��ܥ��Q����17�*�(ܥ�J��t$�X�Z�"��ݱOek�Bd����"_�ø�Q�ɺ�,�-A������c5���5:ն�K{�2��ע�i����SxS%�V}x��WO{��8�4���:Ǒ����k6�k�g,8��ű�9fT��W0�	�c3c�wҦn��ymr��=�ڈ�����b�r�*W�]\Z�zJ�}�c�$��q������{��4�5�[��l�S[��[1n0O�Z����o$p������$ۡGu�7��ZǽS�E�!���<�i��W��Wr����*�ɩ�-S7J�;�ź�HԂ�*�������s�8w��ld��+.�Rr�]>U�W0ғ��s�ꈪ�����?4�=��c�8����}��[�垏k���U5.���Iwa�"E���ۚ�������w���~���P�R�2�(V)h�Z
((�ڍH�iB�Qq�Z+Z�Q�VKZ�T��ĵj�Bڵ%TUm*�ZV��*J�*�1Į"�(ն�W,*(�0�1�[j������ƙj���*%�(�J�%�a���q�ʲƶ"�J�����F�Z�J��s-��+lj�Ke����b�*�V5l�%�ֲ�µZ�*�.12ږ���*ҥ��)ir��F��Ҹ�VʉZ���ej����(�+Kj)E��s9��vn�פ���{p��Xu�6��ܣ�%���u��V]��"Z!��crO��T���Ts��؝�k�%��s��Ѫ�N�Ӽ�C{<q���:1�`��5��S�9��ZRC��,)]8D�6�+��
:��k�ҋ�_�vs��[N�U��x��K3<���r�����媭�\#-�jLWݮZ�}o�X�9Lip&�ޮ��2}G*wA�|Q����PB�N��J���#V��c�v�mJ����~��:\�;�]eo--Nf;��,�d�N��݉)�	ړ�;C�y�YV�ba��%�]����:��
/���z��[����2��)�5ua◩Ɗҷ*��/��R;%��.��7��ષ���1�Q��8A����b4"�q�w��8ee�%0��SkjT!JU.X��ҷ���:��My���t{h=��U��FD���S����d��xU�
4^�ѝw*r�:����3:��=��(�F��T;��7r��"�oo<�Ī���ţ�3�m�#P�`�9�/1�����!�6���)��c7���\�G��CpۀQ�S�Ѫ��}����s�w�?Wr�U�WOz�-�8b���)�IQ�|kK�s.t�(҂V�c�o=�5��p��8f�]��FR��j�Yd�3����yC�����!֫��&�4���������z�Sg�ԥp��E���p��ɍ�X"���0�U�{�p떡6���c��9��+�i��	�{�ø���w�����
�������2�ܱv^R�v���ybw$wnM&Rw��D��ӁS�j��#+سi���I��c�<:a�UۛDU��Fϟ�9�ޗ�V�������;�H����B�7�oZN���|��Lҙ�U�=ⰴ���=��r��{AA�i��]+��Q�*+u���J\K��`��K��rV}�m���{�+s;��~��t�����#��$��x��[���/K�bA'����30�&^���3ɮN��e�Y�������`��t����	B��Hn�׹�N�9-+��g��o���Y�B�fr�uU��X*��&�g�ZBa����,��)�"������H�|�RQ�r��6C]�5Ak�n�c�#cr�j���H��a��U��`ǹ��$b����'����A�b�Z�ེ�5��2�c�=��Z|��z�;�>2�(&��*ǺGV�Q�/��yܜ�1!f�V��\��fa3޹3ì��ի���p��M0Ցg���yÜ�
�r�~�On��~ϖ���khw��{�G�slN�gw�=X���B�]LzVAi����Oʂ��(���"�����A^�h�iD^O1�$\�J�[J�}c:FuM�9���q�
{5l�F���u���=Av�eO��ٶ��j݃}�TR�Uս�i���rk{���,�f1���Ε-���p=���hO�v��&rE%ͫR��=�8-�"Y�O����htw��%�oJ[\��f��|�+��7cR���s���[�b�`������_)�ך���mF��g �׸�v��Q,j������/L��1;�+\6��FNײ^v�A@І�8��ݡ�Cvx�Kv�3�Ą3b�B��&x@�E�[�nsi�]��J��x���ѴhE]ՙ�<77��<������Dk�KTg�2�nEo(��x��^�Lkʷ�Ƭ�/t���|��'k�n�;V)�Eh0 �~>���N{�ɦ�7g-���6��=ő뻧f��N��||�<������S�Y���%a.��(M{�3������K.	7_{�&z5le��I��be�\��C:�����V,����b�+;�\�*�N��*,��f�k�u�x�V��Jw�e��8w�nWR`���BP��n�t�����!U�a����ut����Tl?zv�Ӑ�t@�9�5����)�-�럕ךrٺ�[bD�M��ԁ]�t��mNꞹ����FG5������`n;=[�Vzm�L�G Mbʦu6�U>z{�}S��m�}N�IB6Ƶx�5�,�J�N��H�3fI�aڅ�\:�$P[����f-V�^+u*�6;p�,�H5�ꛌ�:�3�!�*K�:�(<u3%"����U���V��ԁ���L�f-���M`���Ά�w��g���V��VkWM��~�|QM�]Mf������X����둵/�,�S��o$=[4et����̡�����F�y�搧�O�%uy���Ux�m�b'��+�o;:��/f�Ꙗ��X�#8N�Lqm���/1�˅���/
��ٕ��k��G�͜F�4c�Y�S*���{D�(�Q�Ւ�zd�Zܷ�iy
�g�mo��(ԇ�3���dSGȧ��ty�h�J\=�QL������"ph���G��˝�N���r?g!�&�E�� �N�R���v�����Q�ݢFm�e]�di�ޫ~��y԰X.���U�V�"�yO���:ᔞ�D�v���h|��yX�e�Γg>�`���Xv�� �RIwp��%�cjL�4��&�����o�wr~��/��Υ���=�~B�^�����A��.J��W2T���H�݂`�>��ɛ�ڼ[Se9<�ͬ.�R���v�����%�8��ڡ!�x���n��83��f��i����M�~!��d!8(��ڗ>,lia�a�5{u��xe��b�����l5�C�tv���t�����Q��eN��#yhѝ5�f3+��nL]"�qk^f�v,7E�cV>9c�,��ٹy�6e�/"�ASz�׶��]l�ѵ�]���`��1���$��85�Y��t
`>W�=� ϳǬݹ�;w�w .�E��%8J��'ZYO���w;@�JI3��V��\W�l��gE���1#�,)��i�H����tJ��p�q�x�j:�B�ë�v8yC��a�6�5�&�d�|��VR�P,
�{V��H��-K��w7O �wBsǠ��`�w��d�Q1��"�e��	v��5�l2'Уn7��jƨ������n/�	�ӜiB������8�2b5q��bm�ء<iҩ8�Z�׭���ѰU�^E�v�s��h+����и�kmg���`x�`)�3I�mV6�u�����~�1��ك���pb�>�x.�jaݓ�-������a��J�_�� �6�w�b.A�ެ�B��:�Zڮ� V�[[V���2��3+'u�Ra-���䒌pUႆ���<"�ʾ����\^�Tj6�����Z�b~7;x��:�)0��e*k2x;�\�YC��>�ޟ�GK�)�D[w��G�[lK8М˅��c��&��ȹDڎe"�_N̈́���ɷ9�����A4T.>�~�k�}��AP�~���cȼ�˪8�Ss+4��֨���:���+Z��MY�g��}�!��H��d�lAq��lM[�Dpy'L3�K�-�v0ʴ�y̌=g��zA=���EJ��I"��%(�*�s�(�*�!(tTT5��F$#�y���{�P,4����?��y��D�i,�>6���lr0EPL *(�(�H(x��%$�!�a��P�'�Plc�-M���])ke'�7�AEC��&ٔI��\t�v:��&�8�� �Т��ܸt`@��hD3E�!��߾҇��&|a��]5�Y.\��,�%�+��jUTT?5}����]��}`�\�;U�E�DP��D�)lrN��0�&�?�?� �D�\�����N��y���ಎ�%EC0��쯝��9a��`�=dR¥�úL�F?���.$�OiE�AJ�p�*�Kb���s���$��l��wbūBw��"��C3u�u0z�Յ`cOV��EBxK�t	��gq���aF��X,�}3��N(m�?����(�*Wq!$�G�C�7�n0����]*Ќ��i�n����K�����5�=����Q��L��΍��4*��_�ic��C�M�'!?Q9sCw��&G���
,:��(2��+���ǧ�;.<����7f�6��+���9z�hdo;�U�u�`L�=]C�z�����X�=�P�!ט�F�L6���!`�QTT>����	\��=�(N%��C�40?0�eҁM��<���aC���	@Y�7а>Fc��!TB�-�[�@AN'@b�=XMHD��* �	���A�Y\qi���j�����ͰI�� �LAUM���;�X�B�"*���'��/�+�߸���>����W`�����x	`S�pq]�3�uB����Xrus��OX��Sz�|8�L���(EQP�9�/��8 2y	TP����	�O@���K�c�6��D>�hX}a�רw	��ch���	� f@�6Hz�с@�6���� ~ b��@�>��6x������_n��EB�}bt	�a�2��I`�]�܉�NAD7���;�ȝ1(���.�k�e����7�֛�1UQP�A���|��<D��3���8:u�*�*���	�6)��C�^��(\؅��z-k���$arH|
��#�����ܑN$)��