BZh91AY&SYC僦 �UߔRyg����߰����  `_>>'�B �H[x@U%Ff��T��4�)u�zH�ܨ���vh�������@���Oa�E^(��g@i͔8\]tt�1�$��$]@twaK���W���m�\��{;�!]2m���\vU�'GIXp.P�;nfU{� py
:em�VU    (*�2��H�%�(|%4�O�U)��� `M4`L��I)&@4 h     ��hdhd4hɄ`!������*2b04Ʉ �!��� T��0#	�zM�jz��@z�<H���HҨ���jz��i=M��420O�풪S��� ΂��"����Pi�"�/��*A����	TQVAC��������������6��~r����������c��(�U��NJO�|��#���X���Xfxv�$�bv��JRO
=d)LB$�I$�S�`=��� 
��'����������/�!����3�?��O�\�>����ځ��[�V������;�G!}��A�N���]4��n嵃"M��7��q8���<�Ι؈�'�gD�%���^��:^ҭ�o�p�g���^f���NӐ��.�w��z'��:yӽ<�秞�s����N�z<ﭨv��0�Oúw������[�x2�,��}���9<�_�q��&�K�Ic��gN2�V˱�KdFO	piܴ�&����h�#؞ȏ�^e�|e���vq���Y���&\��G���5업�%��_$���6˳�D��7�bH4ܴ�R�~Դn#�K=�Nd�~�6��i������K4�Z<��xG�2��Ìٽ7}��l����ʂ2��Dwc'8��Ru#�	�H�O3�ه-�[ela��&dz�龙��Ì��[e�zsl��Jِ�˸�5�y�<�落gd��IѮI4,Ԓ��[r�N妛��w-<�Z/��D�;�}^���O<�7*S��L����%�����zusu�	���O:s�o:Μ��yN��,O��w��ܘ�u0y�u�L!��N�3��}�o�m����}��zx��u�С�xwý+�>���{������
��v�zL�Nxw�W�^��>:��L�%�VWrl'Y&�"ZlM�RvΝ����I�-5�w���jS�6w���#�;���$�F�% ɜ�^��	6��E��MH�#�������'zC���u�N���x��}b�����&�Fv���Kr�ܾ7/��i�D�7/�Ǳ��{&jw���3�3,��VY�&L��l��7����6ե�k�?Q<Nx���iָç�"}9�;�wɾM-�ٗ7|e��aٝ�&h���PU�S�~+�>�������e'��f�/��%�/F�A�JdH��G��ǲ��O�����2󣫗�k�Ý�w�_:>��Ώxi�n��<^o����7���:�;�s���O�|;�xkm�����龓�oO:po�<'��i4���[�8ͳ�Y�Lä�2���g�n�A���.f*���Z�����[K��ǟ"��9�q�5�X��5��pfܟ�c��T��KxV���_���mC����M����ԍ���9��a���H/kh#��0]��{+���B�}ｴ��uJy��Se3R5�l��O��
�q�qC�XA�s7��7���A>�>��c���I��PG&�$-s�1H�Y9y��a�/g�wp���T	^q��g�1�� ��or#��£]����FمZ�*P��gL/�o�������d��6���h���x2 r�iC������c��6|~�{�)3��BU���N>�G
��ǹ�P�Iq�I)�0@ǹ��!'�Qke����>m�ݠS�s�R�'%�,ɻZ���$�j�O��uq�|�L��ٞW����K
	0�.~�5���	(�,�h��L���af/���N�ڕC�ǰ� B���NF�+�8R���x���ޅ�|���y���8�^x��0�߾�`g�����9����D��8�f�'QM���mǊ6FG���
�T:SHU���(�LUh!5[OH3Fh�dwa��Rw����<n�]��M�[q��׳{��x8i$����';��Ji�D�ice�ݐ���&螏�g �l�'��	YHC@�2��{��4����|�V�B�\i��Q�CFY���Þ��<�<)�m��[y�@@f�X�[�.Z_�U�hLG�#t�9����oz��o�I����s jqZQ��A����;^����)�k��_P(�SI� <��phP�{{n;����'	^v��7A�)������沔~oO5i��k�HQy��M(��������qU�+�oZ��FՖ�l��Y�t����|*n[��,�M,�R	����MB8ӊ,D5��w8U(��-}�DJ���Ιه��F�%��<�+�멎);%y-�v�!6	0V��<u�,'3�T�E+)��BR'�'(ɩ�-y���q�믛r����}m�|�m�]=�"�U�!NE5��3$��(7���y����v��������}�����HZ���1�������%����6�Y����|�N��'�����|R�s�O��-��|��n�Q������-r0%�c`�d�WsF#j��-ʛT���'�H�Jc�n����(`-�O�D��I[�P��ٝ����n}b�*���Wy� ��.(�⍨�#fDK���e �D���J�65�kTp!��h��-bd�b��P�l%���cR���GA*����B1��gěQ5YZr�q�i[Q=G4U���$)��m�w�k�2�	�T�
��Z��<��%݂r��)e��1I��ɓX�8�:(ώDP���4���pO8)����*�mU)@@��g��J�I���ڌ��Uz��y���A]��x��H�P�a�M����$!$��qB���m�`(��U��������c��X+���1�/o� ����?�aڠ��5��{�|�������椩D?Z?w�iw��f������#�>�����X\
��|�/�|�"�U_1U^��n�EUW�]��|�Q�z���ܩJ���TUUTUUŵn�X���UUT�\6J�P�URn<U��b�+�UUTV��mU\X���tU���v���!A�h�eV����EHU/U�y�mU\X��|��ߕt��V��{�;`�(��@�4��m<H�Cd.Q�oWB���Uv��[UWWZ֕]��Uv���K�@�.��4�)r�-�̴wYxɐ�&K+Ѿ��]��v��U��ӭZ��Wj��]���+WE�X�*ID�Uc{�tT�x�sΕU�Uv��[u�QU^��Uz��ٸYg�ֱImXZ���b�p��}��UqmUx��]kZEU\[UUŽUV�CE�J����2Y]X����q��/�����Ӄ�x�?�}�� ��eKmQb��>������!����}o�����} ��>3��DN��	� �DM	�6hM	М,���p�Y�'����"x�ӂpKĳ�UXJ��eQ�ܹ!٫< &K_������SI������12dH�`�X�B����m�*_nl��n�5���`��@"���4��k��-�+d3"r3��e	QQ?B)�ʊ�LlҜ�D ��E�(� ?	qa��=G=|��ߪ�`�MW�PA�����"v��� Q�$Q���.Ǣ�P�n
���D�J�$X�jB��§�*�Eb���W=�s�����Q����UUfffeP�Y���������
����ʤMkZֵ�Dx%6l���lO�툽��M�&�	l �Y&FӷńU����4�$Bbz�Iy��/⻋i�-�ni�I�ᠫ��F�tQ�瘼��b��#R8��g���4CВF/�tѲ���K��Վ��m�LoMcn۹�+���Ra2�I�1�4K�pQrŌ��;K�I�*9�O�����瘹�%�� �c1�L*@��Y���w���d�zI:ݣ�Qz�Z��Py���s����{�حF�%�i:����<L�LL�M'sq{�Li���(��z��*������ڭ�8�Z5��'�W��"0T�
F�y#��Z���ZD4e6�&K�4�:]y���Kg��ƾ>���=�H���
�D�}��Ȳb�g��b8�xwsۗ@?x:K=ĨUz�$�������Ō�.-y{'Zre)Ī���ȻgrvYwfI�5���=L�Va�I;���3��� ��ի��*�[���]�j�/Y����]��)�� Ն.2�ĥ0���&
23lU�w�@T��V53H�M�[�u�%$�Gi�Yt�ݚD����+dP��V�c�	L\\F�&�����ێ�ҙxVffeZ�M<4��sm��ow-�N��u�24�>*�|�Mq*��9 ,�~`�B=#|o3��@E�GG��8�u
�F�mh��1�OSw�pw8-���ol��b�k�Ux�����/��ٷ�l۷��b�|]�p֛em��m�v�\<g����//Y��_W��q�^�˦t����m��]�3j�l�]�ͮ����Ǎi�;_Zb�<�����ļ�7���9�dk�~i�����"�y/|�ӻ��x>���,���,s����kߥ���9����6�l��l�� 6�lǞ��0 �u���M)iӦ8rW.�U��X]���,x�8��	��D
�d�F#��G
K�B����%Ġ1�����S{�	R鉇�˷(�Q��
.`!����R���&�Iz,^�v/�9��Scz�"HX�Ro�r��i���_%��ub�H��%7�60i"t�r-�5t���0C/�Zo�,�<)&Y!Ɯ�8rxU�E�c��# ��J8$�%5P���o�����HC�Z#v�-�QK����J]�h@��<n�0�$x���-�2�p8kꪩ�ZӅ��Dpܦ�
A��i�sFJ00B���u��a�&�M���$�t�q��ˡ����f������ԨT�F鈼b`��	
O0�/@"r�YMXq+O�,���O^��Ó��0��.Dc�:JO�"�/Rs�r��B���ZP�I�$M ��%�ݨ��zO�ٓFJ62�g$���"SZ�p��Q����˶��@�%�u""q�Y��п	֍��0�v��Ʉ��\��Q���s�G��z�ʚ���z��n_�p�?u���T�D�kUDV�*��j(�Y|!Ba��p?(�@��T�ʒ�#��)�&�R�撅��|@9�z�L0w��5 :�i2�z�$Ku(���n��������jK�EQ]t�H�Y�䉈6p�F��e�Ӕ���� ���o��l�d�G�L��L��Җ�SV�J$�+m�.���_&��f��N�8i(htR_��%E,�)�����_����5]����FY q�$�I&p����ާ-�bZ�z��_4�˦��<09��S�+�/'��E�6W�B��(����o���%Q�8��	Sj.�=j&��C�Uu�cM5�<J�Y)�WXCmӑn�Z#%�!�� �mN�a�'RX�2��zĒ�%@=R��L���6^��	p���+%]����6�]�n���v�6�m��핶m�v�\;c�����k���v��/L��;v�޲z��_�W��m_cj��6����t�z�*�|��`o�G����w��1����L��f�X��m[�g4���.X�n�]�(�j�x �P���H���e<}��N7��ND�o�!fH�Ci�؏]����@S$ydٗ=/qhy���DD((D�$ �JMi����=��8G�)�'v�ǮEuR@i���1z-ՏSRb0�Q�� ��!�5��Q����m�[m6^��/<�i�m����!��M� �`���}VH�����""�� T��V(���a�$lCa�XA��+��\V���.���nf��+�$`Bd���m+񖗷j������7%8H�Z���Q��.X�`��V�ZMި�K�h8�6��Y�\�s;�|�M������0����2#��mV���Ѥ�����2\���j�*�2,����,Jz���g��$$�]v�9��Қ��z�Ǟ��5�������+���'.�,�ho��|n����~zβ��x�.᧥�!�MÆ�L�±�����Q��/Ir�I}92�V?_�S_!z��-^�����UV�F_�A"EH!B2	�8L�Q���r�x"�pŎF Ѧ�$��M9_�l���M8�Β��}�y�`�զ���}p��(8��`�9y-E���[�����b;�O�9i�rr�	r�������᳧S,.c�,x��.蠹�z��Hq��y(0��Âapof�0x����;��\B�(���v˄l���	"PVx�5�QU�,Ql�p�-gw:���2�h9�$�bX.>n�7P�(��Ō	��%^_��,����%�(��E�r��㍧�y���퐳E�e�]:!7`띻N@�0/�ý�J�{	�l%=<Q�%�>��q�|��ʗ���OP�r1K�T���X�Y2���Q2�n!�c�%���L�@Q�q )�x��0��tuv&�7�c��Py,V�Pw%[�JK��e����ȾMj�ER��I�b���(*�(��V�S~�k$d�|��t2�d$nqC�G��Tl�����0������2k���I!ćo�ٓRX�*��C̪�k�U��}o.ٷ��=_^�5����̾�[t�6񭵗n��.ܳ����\]�eu��t�=v�oX��=W����z���_����٢�+�,\���1��j�ݼ��s�Pth��#�h��ooh�������F?h��{=���\@�mq�m��Ͷ���k��k��l|A��(!�a���A�u��A��m��_�r�����1
5��F����g�}��f��㗽�ĵ,Q𘠺d��M:|c��1��Įxb�ȩë��.�-kB���[W����t��4�����u2o�[��J��m:�p�C�ߝ�(����7��Z��,���k8��(ʤ��ĵL;��*C`\0�i0;↮%!Ԥ�`��a�8X��!An�!�X�6d�,�週�s��%&�E�6/T+�4�)
�\9D%�/��:�����%�l6�np��I�J{���෸p�b�)�v��BCyJvh�e�2w�OC �t�y=�Ip�^����`��q/s�dK��s�ے�2�u�+V5�C\�d����J�vᤸ���7.���4h����R�sq�W^w�P9Mp� 6��!9۝:n�[ɂHX�6og4@�:n��8xّ68��<C������Qʬ�l��_	r��"j0֚�Z�:�m���E�LS����Q+dC��*|��!M��;e�K�.b�������T�����9h�b:cXlk�Y�.e0�lot�<�=�%7�!$vdѓ��.Q�����w�3����X�B�Y�'�ٓL�ne�����L�͌g��f���,�*=��<`��۫���3	.�����`��7��P$ɮ��{܊*��˙��Ⱦ~�b�j�����QcUg���_��rd۔�J0�0�K�4lє��&Rݗ2tɒ�8;�Q#ޖ+�ca�!M�Q_V-�����e�^9��s��q�F\m5�$�q<�.����<`a�M�Ƣ�ϓ�0�Ƥ�71�Í�.�4k�U'�R�Z��C�em|\\/�m�mmvᶶ�m�[o/��6��+n���]��X�y^^����\/�����/L�ztΞ��{m��ǭz�=V���v��_י{O�|�E>U�GȨk��=�;�BϜ6��օf�h/�R�l��F�wZ.�j[͆�X��[x�I�!�4"28 #q�[j�D�yR;���
Ȭ�dV5Q��<,5�nd�n�M�Y�Ɵ OS|~GX]t!6�}v�Y	���tY��a��m��aGM��
�!MDYFCFԵ�aH�-��NI�SmE�e��A7F���Ms�s�oH�mq�m��m��m��m��l6�k�a�@�Q�C��E8!�!�M�>D�p���QB;
Bl���腫�G��5e�V�\Ta�q���hΉ3V4|h�b��T�['f���bթ�Q_�{�uGe�ϝL%&l���6X�p�a�9-֌	���2`���J6d�Hz�|�޴^�H`rX˃��RUQ�D���`�|�h�&{s��jXۆ�u��]+;6t�c!���J1U�0��M�k�<-D$:7\���6�A�2�)ܘ6d�x݉��-5R֣0�X6�p�[�GDӶܾ4����]#���-@�$n�!Xh����)��-�H�h�u�f�Ӧ�f�b�����$�Ir�t��4�7�m���ZW��%��a%3��)�!U(��b�]�F!�(���b�փ��݄�\��^͒e0o�O=$�E�xQ��f��[�����		%SL���R�dfJ�a��X��ƃa��*\K�8دl�i���/��]�?,�2�U�f�m�S9�_g��E����<:p�c!���s>�RT�4%:ny2����ŋ��F;<��>�ZE-�sp��o�Ϊ�|�,y+8��F��;y�_4���*�\��w�b�E�������KZеE񣻞eQ�t`�d��Bƌwɏ5���nqD�л�%�<j�EľKW>�3���9��QI esl��&�P)Y��fF�q�bml�=X��Q��!n{���.��Ml�D�qM\��%��1�Q�!lYU_f���nE~>�7����0��y�x'	Z=�2X�`0k.-%��f�����O������S�M�4e�6M�����m�\����l�E�@�]^�q����}�3s�i���Q��q˗;y�L�1}Z���qqv�z�m6�m�vͶ�Η�����[co����[���8m�^�m�z�;��;^�����^޴��g������������]��?-N/�SQ|�FK��O�~�]��/�ޘ=�/��7s�F�{�G;�$Ͻ��ϛ�>k��m��m��m��m��m��:뮺WNZtrr���"�+#���\pwM�ܖ�����ō�1$$����5�3����q*���Lu�-Å�m�!,d2�b��i�6ܻ�r޴�%���L���.�{��X���a�x�Qܞe��b�'P�uER�[��lcc@2	��Ȇ,u���$pL��?�$�Z��\]��1\�ߞN��z���۩��O�2�ŉt�y��1\ȯPH��[�J���<[2<��x�N����#O�7���.
MnH�q��y,��F�ϼIM�O�ܫ��A�O�F��MC;�qEs��pa��ۭ!b�C���v4釶l	b��Vycؑ��!t�{�[���Ա����c��ld���!��a� XH�γ/R��/l�u�ҭ
�8.m����.K���(ه�G&[>4x�h�K�l�m��q�����x����/����bm
�0��p�%�h6fpD���"M(�RG��t�kN/(��>#m���IT���D��%�b���n���Ҥ����M�:����:q�d,x�p9�ө�;�@y.Qf�i�Χ�t�B�I�I�UPݪ�-E[��8Y4o/K�4�h�m�U�GG.m���Y��33�ga|�U:Y�w+�ܴv挷9��9�B�W�W&<S5r)���_�h�)�;W^:C�p07�x�f�.I[�Ss e��p锏D3�I�J��8x�/��I���x��m�N�<jI|x��h��b�bT'�Bx!�x����6��k����v�k��fmn���6��M��+�L�q�p�6�.�m�r����;^��׌z��O_�m�=_W��v��^ݽ�흫�_�N��U���%毜k�G�W6�l�&]�y���0�X�f�I�;��R��ĥ��8�B�|���%H�D`�a��	�����Zm�l2��Hߓ����+��rSb��pC��aEN�ϊ�KH$O�Z���86��$����j)SNVK;u��֤b�V�ǣ��lx����U��p�]��cNe��Jl�D�MqE6�mv��Q��	�o�ݶ�mv�m��m�{g��m��m��
>�S�		@�08���	N� ��m&���$�wRWjm���&&�L\��J���<-R���R]8��2y�7z�2�a-E��r���<`41*X
i�G�ng��č�'?����.(�K@���n@;��/p���OB�E�4h�:l0sP�Iy���؏hs*��%γ� �HJ��׮���E���!�&�M��Kg�����Jӗ'3X9�����s<a,Ԓ1���)gB�rI�=.�5c���]&R���٢0�����N��q�d�9���ڛc[Z��Zꌃ���z���TBC,L&�{�˶�)|�M�m���pQ���T���n����d��ܫ�M����q#��m����X�B�>��s��3�δ�S��p�Ե���n�,�`礯;2Y��V����a���K&S�׷N��0�$�q=��I*hyM�<M=M<MjIw�6�2�p�Ҍ��j��#gx
���}��UM5$ �ld��5Ze��g��	��MF�:i��n�f7<���Ե{�σ\D9��8��V�I�)Zjv��ܖkڡ�O�(��X��M��ܓ7<O>��^8�5�m��F�L62�߻T�<�)� _z���us:!x�c����j׎6���T�����m�c�R�߻�㸘�` �+*��h]^ĭ&��ɶ�M������__��(����UVnN��<��<x�D9A��َ�b��U�[+�W�U��ͮ��t�[xͮצ�k��fmkl��m�M��s-�xm�rͯY��p��徼gkӶz�oY�궻z�W��v��_+Ɗ�<\�Ŋ:L+�߽�z���cؽ}Rc޲��=�twв\͍���W���e_t��m��m����M��M��M��lA`�
>�@�
8H!�|W/����'������r2���qr���5�C��rt�M�%U���`�`��U|��&��y	��Jݶ*7�=��3�x�ϲd�P���p�)��e����(��k�`�m�l��$�;%N����2d�
�Mxy<P�a�H�T�D��&�����]]ӳF�N.��[��i���Mg��	]�L�s�84`�FL�nr6K������O14Z-Ғǌใ�3UUUU
��*�h8�p��a���$�(�ͽ�c�J<d0QֈD�6�f�wx�L�ٰ���-���&�T@�FM%�Ϥې��ٳ���d	�����ަKh���0;6��t��v������V�\N���Hpn𐏜�Bi2�u.X��	$����Ɗ<d
>�KE�Z�"of+*��:G$l��H�,�r��ޙU*��B�Jtd�����h�hߌy��d�L�Y�t�Y�5�i�v�/�x��N1�1�'.�d3W2JL8p�5�:&���)˃���j���b�ݤ�͔P�K�dC��Θ<rQ⌔t�`���6�)�V[cLB���'�uL_���	JjR���SI�۽��h�̈l�}v�J���|%S����ɳFN&�q-\�'��A�2(�C-1n+�����C`!#5�^☼Fp��ضL��_>rQ���ڪ���i�̏�~\^§O��0h��-B�����Mm��f�<m���m���6��]�m�p�o3&r�6͹f�Öښ^��L�}^�����<z�Wk��_^����m|x�{^�o�1�L�	c���'*O�>X��E9�˽�O��yW�r����	�Q����Ǯk�c�UM�Pp�#��rǜ�硠��]c݌=O{�=��Q�>v����=����ם����ȷ��������[��x}~�.ps��a��Ԣ�Z�"l���{��UU�)S�#��6ɛ6+�+֗,%Oc���Q��z�f�@����4�EL�c�6=��� ���l[ѻ�&d���'�sn)/��^�z�g�f\�/\��A��|,TLP��A�F�Bi���e2bv�U0v2Ƌ�JK\�E�M�^(��[h�	YI�#-�a�g�����m��m��m��m��m��m� �0C
n{��u�	���S�'�0�1(�VJ�*�����%FHXKJ&K�J��B�R��P�����S��\�p�gɉW�lv�g����3����FG��Q�?o����{������3f�����J����0���9#&6�-ܝ�V�Z�Ъ�V͏%Χc�'��1Yz����
:l0g��	l���m4������g#�8�[�-bKU�����D:�oު%R`,a�ziR狖(����9��%�}�%��u"�K�N���Q9�|\�^��B�O�!��[m�[{���p�M�(���f�j�����T-GF����
۶�Sצ�I�c�%�*�4L��dPp#�eE3Wc���D�>a
�M�Ͷ�q�3����ɴ��pM��T�0u8׌�c'Mt�`�����x��Y(���k�z�0{�d ��*UT�8��t�9��Q�{[fÀ�l\�����Y��&�z�
���|��s$�4t�6n3m�� i���p�����˷-���]�⹞�k���g3�@��9#jM��~�s���%�:���wŌ�5���9,��X:0����>�E�锛�jE!a#n�A	��`�)l#BB=�(-\��(IeU7q�"��`���1�\�������5�c�Ƽ�F�Sg��OrBB.u߬��|bc6���(�J���x�)�0�>Mx�(�J�~����`܍3-V�s� ��K%�Rq�=�qp���2�~'��'b������{��#�e�Zbq:�����(�P�:tK:"!�8A ��4��Z||i��,r�˖�t۶ݶ��om���rۖ��dӎ�Oxu�Nd�0Q���TX���8�t��e����g�<��yǯ�ȼ����6|)}S���"w���6�w{.�{��7�G����q�Z�n>�y8�H�<K������{����{ﷃ��m��qoV�آ�>�g�p�-����{��[b=K�[����^۽<}������Q�t9�_��N�i�:�X�_��(����i��m��m��m��m��m���,\.^��A�w�� �.}6�&����Oef%�&b[~|q�|�#�6�̛,p.{â���2ZHy��I�*�r�i��[w;#l4a�L�l�-��!���νzx�x�˪�5�7rGId���I5��NV����F�m���x��vm�l�q�K�OXӤ�y٦N��.M66�K�(�oS��ZH^�Z�J��y
��O:x�L�.x�car��-i���^HV�L��i<��t���6���q.�����l����lx̕F�g�t��؛���#��,\.e߄�ӌ�]<6٪��UR�]����Cؕ�� l��o0t>w�Q����OŹ��7��#�v�"y�2��h�`�8b��қl`�������U*�������j`I[�5�DF�����ST�$<i�y$�Iӎ�o{�L�Ytٻ8k������?0 �G� J���Ǒc�r�Uz����Ǒ\1���b�U�:�J���̑�4�M��a���g3�K�<��:�s�o����2�=8�������u�{$
�'(m��qy�o����x}����5���=*ؖ�-i|V�nz��F<W$%y�c.�u3�h����.paPe1C�Q80L�z߸�,�/�|m��I$���6�����K��ct��M-��6�rv4�m�}�����}�ʢY���ԯ�1Rܩjն�j̩� �bQ�����~�?�^�"ɋ����,Һ1�i�MPj�I9Y	��.3���殖`�%�l
TE$�Z�Z�S�2��'�d��IK
P��R�*��1
Y
TJT)aK�����K
��IK)aJ)IJ�XR�a)R�%(R�,)d���)H�Rd�,�R�R�K$��R��JY
e':,�)�R���T��R��ST�JX�Y
Q)bR��"���JT��LIJ)IK$R�R�R�)��S���)E,�QJ��%,)H�H�RdJX)��RȥE*���I�z:㎸x�Vb��jZ�-E4��I�JYK�KK"�E*R�j�##�Qe3&R2P����Z�iIe%RҬ2��B���R�Q�a�,RdP���iZ�T�EKEQb�T�)*��MFFU��m-��Rڲ���-E�UKLRb��E�Q,RU-,R��Q,����K)%�*���X�R�)U%�T�R�ʪ��,�e"�KeJ��-UU��r��E���)T�UK�,�*��K,R�ʪ�*�K(��b�X�QeBʖQeB�,�Ub��� ă����$$�&a�R�ʪ��,T��eK*ʅ�YE�"�KH��K(Z-K�RʖRQN��Ֆ����IbRY�E$R�� 0XFA�$��*JY%*E(��R�K,E,IBȥJX��E,��R�,)��Ȳ)d��,����*R�,)R<ױ��ReE5{���ჶa�)��Be�;k�?�~���%�"D�"����y~)*����5����9��߿�?Ç�>��o�����A>#��C�9BD�n����HC{�|�61P9A��/�!�;��$�������:>���_+�B���w2��	?:]?:O�����|���~�`����?ނ��
�����O����$?�	���D?�AE�R���QK	?�%Rʡi���'�I�'�}�t�_���O�p}��aZ���J�2��`�g����s����G��}��}[�?�Y��ߨ}j�����bA!N����4����q������86a�q�R��l��&&I���b~T��6'��dJJK%ς�@��.��w��mHk�P}�~c�O�W��LYp���F����[+��>_��Â����*����CQ'E�}���4P���ʖEX�G�X�JF��Ő��HL�&X���3:�j���CY
�S`����F����������K):Q"e*�J�%�P��Q$L��Z�"d�%��~��~���������t>���������"d.�,zQ��'�#�~������ �а����������%������cH(Y?"�0�d>�����O�M?�~�}�~-��� 7������[���e�_��m?����.���§좏�}E}�?O�PU��?K�����8~�h�4P>A�C�ԧ��H��?wW��?X}
��4=z��?8��}���"��}���ȅ!����$W�>O��?	D������6��^`��!c�=+i K����EE����)S�ҮM3�1'��p�f2Ē$0�������|}:$�#��d�iNYS21,?�2��W��sJ��2��Ӕ"؍�Z.���\��&�I���\8'�)	#ｶ�m�m?O��_���>�P?0��Q��������_�}XC������o��O���}��Ŭ'����}��p\l%�O���?�3��?@Ġ>��a����C��H�\�o̗O�~������������؊��\KG���}j�d��A(`����6?:(
k���K��Z��~�? ���?A�?o�?������g|��b�J�+����)�5U)\�V�Æ4�%�>��-�����0���Q�>^�FB	�.��|o�ؙ0}������D��	�l��z�6���H���`�2�)%>Io�>�>��E-�0��K��$ ������t:��C0:=O�J�H�ß���r�$�}4y��R������/�����O�A��m�[����	��,~	?��;���tAE���ϴ� �� x2��K���3E��r!���}��Y��#ڔt���H��~a��V�w$S�	>X:`