BZh91AY&SY6>f��M߀`q���b� ����bG/�                  ��&��m��6�[(l��M-��[5ZT͕E��Z�JZ���ō�6�-�6�Qf�YR��Ԣ�-`�@�V�CU���QG66�F�CF�Xj@K@���UE�K#m,��Z��'j�"�DZ��f*��km�:4��>��ݘ��z�R�' �ZL�n ���PY� u�5�i��� Z��j�mP���6�l�S��ZԬim���B��U���n��RD����:��!@
E<�$�  7�TN�>5A|��������Wn�������kV��r��Z[�Ǟ��'{����H��ݝr)>�3�C^�������ѯ{�>��Q
�٭V��я��% ����;�t���{�Y]�+��������7����ݪ}�x}�W��:�=罧�zצ��ٻ¾��=>p�����קU;��
z5ҩ��E}5@��65��*���ʹ��=�p��b�����{O}����aϻ}�Zd�4��>�����=��]��yE�}�oK�z�R�Xu���_}>��N�<���������B���3��j�^ڥi�t��5�K*��kU�ҕ �7�Wֹ��&�5�CD����|�i�{����}��j�Z���x4�{��}y�;�ԅ�}y����N���|ޠ
UN��Jz��/;OO]k��8uـjD�Π	�ط�%)&�5xϽ j_G{�������U*������w�}��ӭ[��ƨ��o�q�|��TR�}�^�� {5^��{T�(v}�y�^��������P����MIkm��B��'��JH s{��( �.�� �� ^����} �����z� 
;���N���: ��}� wo_| }䪵`fJ�U1�>I$� �^��
�� d�� �	�� K�� ���wx a�  �W���]{w��<�}�x i���LkT�kj����f�}�RE 7� =��Ɓ����P ���}���������(p � 2'�� �]�`q�B�6el�Չ��-��|�II I�d�;�PQ���@;�� �3����� 
#���P{϶��@W�Ǡ�zN *��:ù�b�,���'M\���I% }���� ��ݻ�:��>��'{���3@ [���@)n^�� ^���G����ϒ����   
R� P  �JR�4� � 2b "zhĤ��0�� &!���2	J�~� �    �*jU(�� 24@ i�P&�	��� 4 D�Q��J�	0j`��2h�D�O���g�O����w��s�i��ٴnT��MX�m$�ɾ�޸��{�W��PT]

����D@��N�!������?��C�O� 
�?�$�s�_���Љ��� �D���-�/��_��~������Lbcl�&����.11��b����&3l\b`���&1q��\q�F11�c���&0q��c8��.0q��`c���&1���L`c��0q��L`ct��bc��&0q��`i������&1q��b��21q��Lbc8��&0q������8��0q��`�F11��`�8�1��bi�0`m��b����.01���`����.01��`��㤌bc8��0q��\bc����11��`c��&01��`��11��0q��Lbc���.0c�����11��Lbc���&21q��`����&11��t�������&0q��C�01q�c���.14����8��0q�c8����\b� ��\bc�1q�c���1q���`�&0`�1�i�0Lb`��.11�c:\`�l`�8��.14�`�l`�11��38�����.0`�a�]11�c8��&1q�bcL\`�8��.0a�1t��.11�c8��.3���\`�8�1��Lb�#8��11��L`����1q�c�\bc �1q��`��0q�c�1q��.11�c �&11��v���8��1q��\b��I��1�c8���a�0t��11��L`�8��11��`�8��0�1��b�8��&11��bc1����11��\c�L`�a�`퉌`c���&16�`郌`�8��&11�1�`��&11��bc1�C�Lbc���1q��\`c`F0q��L`����&1q��8�1��a�\bc���i��L`퉌\bc8��i��Lb퉌`�8��0��1q�c`� �&0q���bc���&0q�c��.����&0q��\bc���&1q��`��11��Lb����0q��bc�q��11��Lb��0q��0q��`�8�lbi�c �.0q�����8㤌\b�8��.1q�m��4��1q��`��b�c8��.0q�b��b����.11������Lb�����1q��`����f1q��L`����0q�bc;bc���&0�Lbc8���Lb�1�C�`����.01���\b�8��.16�����&0#`�;q�i��`�8��&1q���q��L`����0q��t�8��8��&01��f�8�����	�C���1��]�q��L`�8��`c �8��11��4�8�����&0q��t��0v���L`c��LbclLbc8��01ۥ�.�8��11��a�11��&0q��Lbc�0q�3�`����&11��L���&11��L`c���&;t������01��01���1��`����m��11��`� �01��a���.11��Lbc����� �ئ0`�l`郌b�8Ď:`�8��&1q��f�8���.0q��`���1q��`��f0t��.0`��1�bc�1q��v�q�i��`�8��&��b퉌\`�8��.1q��#���0`��t:b����.1q��\c���.0q��\`� �&11�bc���.1q�c �&1q�`��b� �.1q��8�1�c:\`�l\`�8��.0bm��4��1��1q��`���t�q��lb��0q�bc �!�b�8��8�1q��b����.1p`����0q��b���.1q��b�����b����1�:b�1�c0#`�8�1��b��F1q��\`�1��6�Glc 6� �(8�G � ���G��b��D6�`�� ��G��C(��*�l(`#�Pq��0U�8��\`��U1�b��Uq�� �\b��Tq��1E� ���ccq��1�(8��L`��Qq��U1��0�+�cb)�Tq�1A� 8��01���:`c��0q��`������`��&0q��`����0���`����11��L`�l�����&0q��L`� ���1b퉌`����N�8��8�1��\`�01��]�`��.0q���&1t��&1q����K���1�c�)�CF.0b����.1q���\`����&1q��Lb�C�`틌\bc���!�`c���\bc���1q���b�8�1��\`�16�``���1q��\`� �.1#���&0q��\`��.0�b�8��0`����&1q��0`����.11�ŌL`��0q�9�-X���z�
���	S��n�-���טe[������,J�k���Aa��#oq;��tn��n�W7��4�϶�-VY�:��X�^��2�V������gt�i:8,��T��-5^�-*R:N:�t���(f��`�	w��\Yj��zIt�9�(������B�Y�c~�2Ҭv��HR4�ե�)�0�<���p !w�m�w,/3*�z��<4�-�,��2mR�m�y-�#}f݈.�ڤ���ܨu[�c�a�$X��aj��	�vT�ɕ{��:fֆ�5Ĵ�z�*�VZ�v��A��A����D��@ʦ�O�h�a��(���ޫ�I��U�E]Ps��fL�4V�N��Ẵ�9!ƭ^e���U�p�7j3���ۋf�%��L�p�BhBXL��Z��љ�H�4ѩW��㴢�0͢P+�j�W19.����h�p�v��^����)m��L
��+X@Y��ӊ�׌^F%��tc#j3@i&#�¥�E�5Ռ���5���(����E6+��+nl8���ҴԵ���a�S���x��۶� ����4L (NC���u��L���ֶ��r��]���k �N��N�hc����c^�t�	n.��f��0��h���a6pޅY���/^�D�+R��Pjt��/5��7���䀭rZUW4��.�⡊,��vA���%�n�[˺��r8#n +���cZ�]Mץ�f7R�����vPJaL�����y��ǣu��g���nf]1�b"�[�i
�r�V%ܗ50�V�`\F���յ��dR�e8-J�7&�1+���@)��N*uwC%q̂�22n�<�A�JOd[���㻲��T��Â�I��;�kQf���T��#��0��W�cW��i�lr�v�M���t�AJI�)]��3<u�G���{<�F�S"�JD;�JdE!uv:�m�b���W5P�!V֍ޣu�A��l��Z�m�/m�.1�L4�%Zۗ*�Lzޭ�^õ.����#���h'dY��2Bm���WOm�,(�a6AD���r��mpd
B�&�"[Њţ5^`���|کA༧��ԥw�M����ef,(\z������ȵ�"�Rj�W/wo%�W*wi�f:u2��蠮��x��[��p���aY0%r��#$�#x���nX�6"���Ә��,�qf��wQU=̛�^��kR�h�lO$��	���)�FoKچ��0\Y3omţV�Ihc2��1*nX���q����j{��3�4�yI�U��ɴvĬ8�ZlCW��"�sp7Z�7kQ��]E��s&(�-V⼧s�&S�7-S��2����l,�
{+d�Q�틍X�r���Pٙ�`�_b�매X�]���Бe*w.��LԤ(X���wCsE��a�kDtr�&Bʘ���k]����xI�Մ�VI68��7��G)]`I�%�>�ʚ�����up���b�Bna
���:YY��Y�u-�:DB
�ڽб� �j���	�`ˬ���j6�*��MX/owr�̺��e �I����I^�-�)v�H��t�n���'��&I�x&cj�5-�#W���������+�W�툯e��jW�м�Yb7���۬te=8��V�,�X+Zzf�`7�K۷���%�v��]U�D�M��`;�]��đl�#.����
�,�V(b��!Sp%�ɣi,դ�I�G�0�34a�/IcVM����F�LU�lKK%J�ȇI��XKM�F�V$��3F�nS�4.�^[��ݥm��Me^�4�Ğސ㷔c-d�9{Sv� ���ڏ1�y&��9Gcv�����n͚gҥ�M,��b�&��
�.�
�݋.�;"�/ZES��R�Q=�,�#M��i�32�޵���F�^"�8���;u�th��]��n�ܛ7�a[�e�z��wVG�(`���2�#�J1\mV�^y���wN��1�8�%r]D`�3)��Y�^��V�v��$ѯ\����l$B��;�B�wSR��Y7I ����f���y")wJ�F$%E.DsY��yX���txJ�B�e0�a� �:���,4�L
H�j�L�h�ᙪ�!����{�5�!t5L�.�:̤*��ɶ��zUہ�.&!A
5x�4��/3b;ڧ!�z�xƑ�I;����	m�d*ǸUip��cmYZ
	#n�J��N�mш�#ƈ�e�3le(�(������7|�&x�`�f5[wG![y`����L�]�&�ݖh�m��ۛ�"�nlϫe����:�{D'A(wDn$| *f]��B����+��n^b�NS���t1<��w����Sn6�$v�V(=�F�ե��5����O^�k/��ݷ��]�(M��
n1��v����D�*UD�6�҉�y�P��ڏhZ���Ӓ^��eD�ִ�[Xl㭌Z�5E*�2�^n��k��=�8�۸��Y&�W�鱴���,���j��W��,�~�1V]`���nl��=7R����JgSv�G%0��f����oFm6��B�P�a�wX[�V	E֛��"u�͙�!a�ꀽ�&�7l��$�ٖ�c��4M	醴��f!o &�TR^+Υnm�)�m̒䩗�.c�6��	֜[�Ԯ�+e(4��� �q�6Hp��I��.x��׸�\�KdhPxE�L:,�kYݲ#�B�����jk�p *;����>�C *�\��w��f���^@Nm�(f�'Z�V���6�F��V{(���U�U��[1�ҢD�M��<VX�l��#���x�0�pj``��������Z��&UI���C����\vҝ�Rʷ�Y�Q�4T���E:@9t�
�+lȵ��a�{V��s^���U0u%�C�Y�Oyv�7�hB��U&^�N&�0P��GI����j��v�Q9JZ���h�^�N����R�hɐ�H�L�/!F�vb�I'.�9��:2�$	�eI���ޭ�A����������L�u	��J���:Op-�cI��@`P�{i�WVVk�0�j���T�6eH��h�A�ض����2�r7@ͭ�D�Y�v��l�ɑڡ�1���1�&��0���C����q�«%���������lݶ������C�F�w6�څm�N9a�R�e����)o�0�5�Z�&��\����j��g�ɧ�)��yhc��)+���r�<�f���i�n��̕��i vm�Ф�6�b�#�S���p4��m���a�k]��ff^U� �\v[�`Stŭ�"[�qD����dmnc�Y@�򖃂�+��c�)�B���w�2襯0�,9�=�D���;��F�-C��o\ͤ��Љ�E髼~��G[kA��h�#����l8f����y�k��:A��hL��:jLU\�K��Z�f�8F���a����,�ɔ�{�y{K	T1"2�L�����;75��x��
$HnFSulӂ�:��.�9�w���[�	��v�܃9��:�!�)�bLF���"���ɲ��B�@V��:������Ekb��y���:�d���I�^kf��rཡz4�t�$�˺w$�L�c7V�r�͂h���x��j��DPl����ܶ�40Jko2*[)M�R�֝y��(�w�dLh�M����Ul�`��M:�)�N�&i���ݺ��YXs{���a���J9�n:�S����v��ܚ���������HH�3v�Iaȫc���h[��J�j��2��l�h3�<��I�������0�j�ݺ.j�����{Np=�I��Qdլ�C�얡���lgi�h��/aS������2��P���ũ��7	�+Ey�:d�h�2O7&@lٷGF)��K/��KY�lIP�ս���ػEV�*��А��.M�%�M�[�ܕu��a�x!
�a���n��r�R�
�6GO*H�4	R���1��$�ZƮ�2V?8-cƚw�7k�x� r���˨IÅ=M�ƔE�%���("vZ��j([�Tf���0��'5�iRW��+M���ɢΧ��ʹ͢F��Q�f�76�扺���Jb��t4e�X(�JJ�HD��U�˪�d8j�0�ʠ��-��h��d�n�
�����(�4E�۸:r0K��;r�o"BE �3U�U0˅�V��8�eI�����zq�PF4lV	X!YV0۲����C4[���!���iI6��(��LHh��Z|�N�q��ѭPզ�pP�"t��v,aɭ\�l촄�v����P���ے�2�U̫3NK����X�qE�ԓf�r��v��A�ReA����8�eG��^PI/M��X�Uf�F�{*M'-��Sq�l��ԋMY!Vm��{a�2=�I�zC�4����ג��7��n�tB�Ȥz�xͻ%�uB�$���|ǲ��WU������t7x��4ELS��n�m�n�G�4VT�mU�B$�6�1\D��hͥ�/]�ϝ
���-K��ب%�mҲe��E�Ѳȱ�Ӻ�c�����^�iL�ba�rMwH0�T�7��˒�㈖u`���AcҺ�vk�*�^�'yH�WxR��u�m��*SY��Mo#x�C%�D6=��Y�1ap�f�/)Ԋ�Z�d�V�JŌ�aS�LoJ�ګň�nUV6������7F)E�fA��+%�f#���[� cYD,[�l�J���X���q�m�[z�J��ۏ뫧v�w�cR��%�i���O.(���L+#t��N;E��~��eCc^�1Xv��Z�+6�ʎ�a:��t�H�m�mbr�٭E�h%�Q��ͻ�`�m���D�x�L1#�-�˙OT���F��;�n�$ցn�L�"B[�ћ{��-+�tF����E0]A�)��:��η����Uv�H�\��HSB��H�������D����Tԃ�T��E%X��Z�z�WoQԂ�f�j��[k��I����^+h�v%�1z��A�Tگ&�h�cE�ԏ+�ؑ�x��V�N���IKV�ԁ�o)��]-��x�.ĹRާ�]��ibƴI�eXs�LY��\�*��I*�#�ڹ�IE1RT�R��(s����Aȹ��$�.o%���OEݔ�Z<��Z�J�b�R���Q+S�y9ڷ�9&��Ok���W�ĭg.#�[��Ȏ.Ě�y,�m`9�jԞ��mW,��-�I�K��9,\I��]�Z�K��iU&5IlGV�ch�y��ؕ-�-^$�%��\��Qo'���Q$���D�qcy&�8�$��v�)�Y��t����ؔ\6��͐ŀ�J��5KW�a�U�%I^,�X�.��h%ƹ-U��@�o7�Yv�`��ԏ�	��%�gj��wk�LJ�j��o+[Ԗ�q�]%k�V�Q����幣[I%i6�V5���I�|#ĭN,�b�aܝ[�����9X3,��ܖ�� ��{o+2��b&�����ر)� �㽗�r]�]�n�2̾�Ģ�km���,ղ`�z��k-H���G�ڬK���3�B�74ԹX��{w}q^&�Զ[���|+]�i_+�Qڷ�.��q&�Uj����Z6�T�JL�wkZ�F^Ժ�Iri�'j���-JRme��b�.�rF����X�w2ܱAe�o,F���3vX-F��d��Z�M��X���ڠkDҖ�.�w&�RT�(����]�X5D�r9I��6:u�2�v��&�n<�n*դ�\_��,-$�R&�򀔯�y-J�$x���5z��i-N��x�-k�T�����m��i%y��$��\�Z�2�T��%�LW)��[ӔL9b�T���yr�Qz�#L�z���9^-Ԓ|�E���4�]�EIV���!R�D�]�K�.o��x�F.՜��Id-�M��$AȤT��m$�ZT�c[jiV���5LO�mkTF�.B�*�b\����)c�\~�k\v��p�Ɠ�g�b[�:��4qTYjRMRW]�S]v.Zx�%Z�\����4�X�I&k��I$�R)KM��qo,J�H��b�Z���52�j5"�`4��i&�R"�%5w.�X�ӍR�M)��0v-J��_*�4��I��j�(����0LK�w"�Rf�����i�{M�yY��N�ĩ/+�*����9y60ݭպ����i�	�ԔR*U�5-����:#�5;F��֜�+1b[�A�W�:�I�ae^b���WZq+\�yHj%Z���E��N��]ʒ`�.�b�����T��b�HԒ�I(	�mj�]��rOR�$�T�K"�ܸ�G7�Ԣ�*�-[j�F�I�Z�4�喕�I5���1 wS]�;��1TH��K]h��N-�b�KR�=&�GK56�����'H┫�|�-;�zE�KQ�q,T������Y1���bKՊZ���5W.�-��JbmF�I��Ke#O���Z�v�CjmL�|�JO�.Mwq\�-L[bv���\�&��赣��؟"�j���Z�[�Z�1fg���kH�v|���m=z +�"lB�%�+Fh˴�ֵ��bFә)�K���I)�Ҁ�L\��V���ܾ���F�W��Ԥ�Il[K��Uǹլ��S����Հݮ�Ʒ%�ĳ���kYZ��%��إ$)���[ԹZQ)�i��՜���4��w>�mh;I�Ǝ'�uǛ�W-�A\�H��/v�R�O�פ�8���x��iLV��Ά�y�-.T�K�F-j�b�W8�9@ZH�$�v�j��I���ݩmlK��軕�R-*SW%@�'�bMbSR��:��U��<�{��X��j,��1ՆZ�S���0r�nG,k�?�o�h+�֧*J�D�M��)W&
�"I8�T��KN-K`���N���T����.�V"�m�U�E���qKOR��=R$�B���u��}>��ݾk�9{��в;������r����/�~o}��ߤ��^��)0��Ҍ_�w���Lwwv������{��y@���aw)�K&ȓ��]�9㪛�;�͵y��,uU�N��C\���w��Wl� ��\7{�:�L1ڥ��}��{�W)��4��ł��r�.ۦBé��<j��\�i��[�ݵg��9ZEܦڭ39�E�L���al��붼u
̢�vE�ʲ����:�=���Ց�N�H�v����1S�_-@�n����wt�	-�R�[׫��	����B��qm.�T3}ҥ�5�(�2^��])8�S��{��_��T�}GL� ӓz���9;��,��\�d�v��ͧ:�F+�*����3s���jq5�L�Mǖ�v�2����t筢U�^DS�����҇3-5̷����3t��E��-^sb`�f��oiW˲s���Ps�ZFTqe.s:�޻;��`V��hZ�U��a���Nt�wm�-�3,���[ks%��4��7L���yD�0Bjkǐ�1ʷ{����(E���#�3�����u�N��0�j@z�u��o-�dy>���2p<Ӝ��t}5Y����4�y�pH�^��O�Cb��c;7��1�5���1F���ν�MH�
�V5O��Z��ͤ7��r��b���jPڢjWN���N;�d�Ax�|�����w��Ife���1� ���6  ���%Vn�!��kR�z�wd�&���k"��ier����-�{���v0b��Av���I���Bm�k��{U�.U�TY�)��h]ۺ�L��"=RC��Ju0�t��R0������W�f�ԝi5/U!{ϑ� �J���!�G�e���v2{tXwȂ�㵻S2�.衇Jt�N27m���&!
�C�ã��#����_#�܁�uSz����)s�]�;Y�D�W[�٣��)U��\���t�f�Ƃ�zC2�,ۘd�;)'t�-Y����%Nrq���o76gXβ�'�r���*1�)�[�EVu �����=�"F6�n���\��.���`u=��W���ދfB�,8�6�L�n��n�oݫ�o*|�LSbߌ�.^�����8C��\5K+�d��.-=�<�z�[F{;Z٘oj+��܊'�~�{d��_ϱ�j=���饓6�q���J�]�Y�0=�pv�gW �Έ4��`)Y�Yj:��s�*)t�]�;�)�t��և^����bݕ+5Η�8�{��t���c\֎��m��\'�l����^SY���u�^���c�NY����w���aX�K�72����#Wb��R�'��E�wӨ^U��^��ySt�˜3�m�_�t�����N'����z�ٔ�t9`����7��*3{�Uy(V�������,�-v���[�&-�iB�َ��#e�:���-�;ؔ��S!ȑs3�9�}I[���i#�kxOp���06��Zv���#(�oqr� ��`p��tU�J�uyڢz��d�r�b��S�z�]����Wd�uW�Ȭ�팙|nF�K���Vlu��[%�{�륩ڑ��9��4�ߝsׅ��g��컥���WWsܮ��k�@���i�#������Yɖ�דi�Z�%X61T�Vyt�� `6G������W��h���ƦM��Y\u^*�1xTF�ɫs^ ����]��V�8z������o=˥s�eK���3�c�*�٨�����[�,�Uك�jc�0Oն��N��vk��#z����6��`�I�XO��V<��C�U��׍˜�s}{C91�:]�=�u*��__��P������æ�� nѲO��Ĩ���k��oL;nڪ��]Yu +���S6`K�e+]agc��^����ݹ�muo��2�0\ub8	[J��/�6��u�Q��vD���8���(�@�CH>ޑ���7��6����Υ�Sz�/��p��P]��Q�	�ssKb�2�1hR�i�=����y#�zЦ3Ov�_�l�}��#v��}�Nw��7}�^e����ՠ�AS��7�r�ܛb�+�Ƹg������6��B����:�Va�̩�鈹.�rn�۸���8��5������0V	�	��wM�ܒ�lB�hVu����^��&`v�[oM�g�%9uh��2�T��!����}%r��,�weG��'�^�'rqR�F�:��yu�[ұ��\�+_YM�dq؛��k)#f���I��ݻ}Iբ+0�)q��5%�4n���um�S�Kb*�ȝ��qr���F�W����f���&+��jtT�պ.��a�Et�+/2�V�P�"2Ԋ� (�6��[fI�LiY�v�[�ֳZ�ؤg^s[��d�u������S��ȕ���K�b͹�Y�3lS���@�J��]ҋJ��j�)g��5�;��=��36�y8�n���"�ȉ��W��tm�3Y�X�nھN�D�������o��拼,��@�mi4��/FaQQ]-�y	h�T7Am��|Wۖ���Y;n��iT8;y�X�����=J��N�N�/t�b�{�VP.��y�(��ɜ��鶦��:e��a��y��yX�&^�pF/1t}��H�b���:��֥`<e�p�"�b7����,v��Y��"�]�'n���3A�|�*���f��b�E1MՄ��#�^�����6���v���ˢ��ob��K{5ٺ����je�P���2��rK9j�V�]-}�m���mgs��2�H4��e]kiV�ڶ��<���Kgi��o7]#���m��f݉���E����&�%tRd!�Z�����\��c8�C3zMlXb��.�d�͎�%���M�[[�ř+�ξqr�M���LT�`/�ۋm�[���w����9x��L9�
����]"U"��3]463��m,���|�]�c[�Ϋy���u7(�ooq;w�[�7�i:=�5��h�/i%��;m��ǃY�Ү���G:�aB���\�߅f-�h��	Y'0���)ia���Vzq���Ψ��WU��v�I_nIf�M�}cmb�`�|Y�X�Qn�2Pԏ����{��Xl���?p���uE��r{H���3Q�I��S�N��k׹�\�nJFx�q� �a�Rw>�k&R�8��Fʼ�G1D�Ft���r�t':6dQ"�:�/*�RP�����.N��],���F'��'���T�۪i7�dQ�i� ��D�Fû;Us-�;뽒s���&��zճ��&:��7�ԗuᇜd��B�s���n�9Or�t�㔩��ԭ��b��%ٷ{��6K��y0�!,���tθ+�jsN�m�ޝ�"�#_iH�%J�C}y
�Wc�	@��#���e��u����o�f�x�I�SSEX�/����D5G�������+;Qf��;��<�*�8z��Y����swxm�+NdK���Jn0Ʋ����j����+����vOa���&e_#���p���M�)�[���đ%ɦk��*�#eɸG( �^���ü�f�ϒ@Փ4u1�)N��d{��:�V�V�xqo���
�v�o!9�0u���rs�ś�T��t�L���t�"�XC�d<D��K�9�M�t��B��M[Y�	�S��[|�ԁ2��ːq���3Rb��y?6�`wY:���e	����S}gf5��jt7\	��)L����1N��}��h5ܦ\�S�z�f�R�K�aՌm�u|�y�'��.²��^�o����K�/��>�Kkl�u�W�8�s��r�%�ՓD��>���ow]�9"��FeoPT |3 ����j��s���\�]��l���/�V�>�����k��:�l�H�8!��D0*5[Z^�Xi�1E����(����Y`h���b@\d�z�γx�������eW�AOj�����z2�E�UEku��A��|����z�IŒ���w:9�Lk!򳼸MњF�J�fQ'��:��Oo�U��6K�y۸j<�BR����`i���l�j��A�,ru��㿞�ڊ�t�g���3��ʅ�|��S5At���J8v�Q�4v�o��n)H���E<]}�\��Uum� �0��rv���٪`���d,}�e/�����4�^X9���tn��z.Г�pN�Z�/xofщ�}��wi t6�mu
�qj��6��n�A�ٗݫX��WL���we��6v��5/��g%m �X\t�/8�2�0��W�<�S�s�d�����.:W]͞�
��ڶ_YՔ�w_�كme���,�4�Ʃ��Mm��f5Uy+kw*��^�$ y,%!Y�HW:jЛ�%8��ı�o2��,]��֍C�6�bʇup��_b�#��LUg&�#�C�u�=]Eө��8���)/9՗�FH }���mjŔ��r��k�N���iVE�ˤ"e�t�)��W
U(�6��3��zt���,�ok�:'�AZ�g0�ӆf�ƹ
`���z�w\{�g��p���*>	f�A��ם�N�-�@��C��4��P�������O9��=
;4�+�O	Ny!�kE�o$���me����7���֍�VL�zMُ+�\C�����wPn�ơ�Z^�y~�Ċ���TYD���a��V��=E���H��ϸ��^Խw��|���I<��U�o5t`�V6���5O�@��}]6����I5��s�9�_N�y�x� �C��.�t3�L�|����y3�����H��t�*7�?���]ո���og0�u7c7/�Y�{�Ӫ�f���e��:�c��4^�	�&h^�p�E��/O�ֺg{��v^��q��eC6ov�Ǹ�}�ˇ�a���9K�;|9�i�o�|�u�{�{R�>��N�Jp>�η�.ם"�-N��M[���7�_n���r�H��������Ꙏ�7�̝B��#��I���6���i�$�I$�I$�$����9�I˵�9պc��3��֠�2�Wv��:��}��Wf�P�o�� ������`��P�uE�[�iS��r��Os�(����ܐ����kfs8Ǘ6�G���z�o8�6w�Z����
9��Z�8�zuצB����!G��j��D�9f4��(�����Q����1C�߽0��8����:I	�]�I�9�{a�HNuךw���N�_@����\1�@�z�/�Ht�$��ܰ��� |ϗ����|����a8���y�=[&}��C�u�<N��J����-�Đ4{Ω	���rx� {�=��2ϓ�wo�$��/4�;��N������,��Ȑ���C���R�N��{��<{��jq��?_�׷��W�}���=�!S=�}Y�O9H�e;�����v�sZx�z�ny|@��I�] �λԻ� �p��7����
ٹC�K^ !t�=벴��=�����T7��j�t��=���w�i�e���h'�:� �l|��n,߾�{�#��؏��AAO�����v �(���|�?��O������?@� ��" ���?�~���߲��������8�E?���ڏ&!���ؓn����:��j*9ZM��8l˳�7�S�a�}L/sR��2.��%����0MGA�P����y���2�I�ҏ����-]�ئ|T�{!q|Y�k\=R.�=i�Ha�B�&S�!���Y*吥N
_*ZZZ0���� w�{���ʛ�u~�4Bkrv�]��R�k)������	>�aos��:�����f,�%���R�ZZ�N��p��Cln�n���IQ45���Rl�u�Ɋ�9��LQь4��û%��o�˖�gn[��\�t���\y�F4;I��c�`9�3
�c�]u�>(�6�bV�3�q�m��2���KQwSp�����S�u�k��ȁ�����Zį��6.G��\u.�ۅs�<9�Ӄ6Ri�g( TQ.��{B%ٮ�3w����JQ�-m-�w�Q&�^���,hD�-��fپ�،�=9���}�A�L�j��83wWד�r�ʛ݇5T���u,��78Ќ�sgIAܒ:2	�Q��b������t7�Sw�y���]﮻���N�\k�Z鯭kZּk]5�kZֵ�kZֵ�kZ5�kZֵ�ֵ�kZ֍kZֵ�k���k�kZצ��k^�ֵƵ�vֵ�k�ZֻkZֵ�k]�Ƶ�kǶ��kZֵ�Zֵ�k_Ƶ�kZ�ֵ�ZֵƵ�k�Z�MkZֵ�F��kZ־5�kZֵ��MkZֵ�k���vֵ�k���kZ׍k���kZ־5�kZֵ�k���v�q�_Ƶ�kZֵ�Zֵ�kZֱ�kZֵ�Zֵ�kƵ�Zֵ�kƵ�[��Q��-���K���b��Y���<��G�̂��f;AWW�������w%�� ����x�����
��z��Dj��ٲV�޷!�҆qK�qg�|>��lË����%N��\[��j�9��{^����U3I�i�Z��o�[�xr��n�k-��0,����������(��Ȳ��4e8���vM�7�Ԫ�Z�6�:�ꬓ}�mmN�9�En^L����C����	���<�#���t���f	N�0B5r�@�.»���b�9(k�8�]��tm�$�;i��b�؛7qy���č�"R�c�s�K�ݭ���e5�&�u^�vJF�o!їp�{��(�ٹF��f�qo�'a6'!h�����[���0�C",������ɸ����O�k�Wod��e�no`��P��!{˨����W.�ˠ��3V��}ͅ��Yۯ �ɩE�#��詪�ŭ��q���Cն�w�e�Gjnb2Dú����Q��Nc�6���.}G�hQ���r���NǇ�o���m��n5���kZֵ�hֵ�kZִkZֵ�kZֺkZֵ�ֺkZֵ�5�kZֵ�kZֵ�mk]��kZּk]5�kZ׶���ֵ�zkZ�ֵ�zkZ�ֵ�Zֵ�mk]5�kƵ�ƍkZֵ�|kֵ�zkZ�ֵ�5�k^�ֺkZֵ�5�kZֵ�ֵ�k^5��ֵ�5�k^�ֺkZֵ�5�kZ�t֍kZֵ��MkZ�q�ֵ�kZֵ��k]5�kZ׍kZ�kZ׶��kZֵ��ֵ�kZ֍k^rs�^k���
sM����ۺ�Kr=Q59vx��m�&<{n�ۺG8��3cb�X��d�(�/��f�ӣ$�NZ{#��as�{Y�/jw*<��Q�k74X�b�X$��lSm��ru�\9^cg�����0�f.�Q�(eɻ���a�������V��ː`-3��m`��:�
�n�ooA#�ν=Ut�n]�w�N��V2�L�F^��i<N����Pv�'��m赽F�]7�e��]o����9v�\�^T徧z`��C�t����\�U\`D]dT�s��l:T4����*w+�)���/�C>ݎ��YR-6��v���Y[C�ReL82��m�E�1@�ݕ�1ZV�۽��|���3��B�YF�!4��E�)^���5����eX�r��m�dʧ��]uM�D�t�r�NѪۧ؅T�bopJu�ɘ
f����M9��t٫o��*p�˿MB�4*�bQl���]�E�;��;us�󐷈�,{*m�яh�:-P]4O0�5r�=5j"�g��������5�k^5�k���k^�ֺkZֵ�ֵ�zkZ�ֵ�5�k^�ֺkZֵ�5�kZֵ�ֵ�kZ֍kZֵ�|kֵ�kZ��5�kZּk]5�kZ�ֵ�5�k\kZֽ5�tֵ�k^4kZֵ�xָ�kZ�׶���ֵ�5�k^�ֺkZֵ��5�kZ־4kZֵ�mk]��k���k^�ֵ�Zֵ�mkֵ�k_5�k\|zzzzk�ZֵƵ�k�Zֵ�MkZ�Zֵ�MkZ�Z�MkZֵ�Z�MkZֵ�}��w�n�!��t�<�t���옲�d�N{x�#��J�ul�^�P�5 swƒl�<����XzG�J���zJ�%u�2��y	��z���qs��2U�s2�!rN�u�-�I;Ŝ2,�&e6H��#*��������3T�zu�^CI<��ܫ���V�m�N�=�<���F�׊�	�Ճ�rA��kaۿ�7�"i�}��r�8j:�_�%K&��Y�H̓l�R�
((m,�v��c�n��n�S$3G�}�˫��g� ��V�)��psͦ��I�W+F[6�h`ܾ*X�ٽ5e(؊�4�7:)2洴�Z���s��A %<��*idczfm^�k���1�}��;�M,���s�GL�Y�b>�v��ٙ�Q�O]��I]j-(T�E�=�ut�U���m�2�cy��ܚ樁�6�c7��~}ª�U\�]�SN���{ۥ3Zh^��<�tm�t�#��w�č,G�Tj���pr�9�9��ae�nޫ׽�G*Жq�_M����[訨(U�.�[��0����������Z�ֵ�MkZֽ5�k�kZֽ5�k�kZֵ��MkZֵ�k���k�kZצ���ֵ�kƵ��ֵ�kƵ�kZֵ��kֵ�k_5�kZֵ�ֵ�kZ��5�kZ׶���ֵ�5�k^�ֺkZֵ�5�kZֵ�kZֵ�mk]��hֽ5�k�kZ�kZ׶��kZֵ�tֵ�k�Zֵָ�k�Zֵָ�q�kZ�ֱ�k^�q����ֵ�k^5��ֵ�kZ��5�kZּk]5�kZ�ֵ�5�kZ�ֵ�5�k�lu7�)\9u���`��tԎn����Y;s6��e)Q3n���Sx��rd�*����p������]s3o�J�.7���i$󚳣�����R�ޖ[�[�SѮ��i\���8��skLGe"�Ҏl�zN���֫�m#=���R;m���ew�9Pς����+�z6����+S�c��"�ǁV�G�� j�i��׻���H�Dl���ѽClJB�RYr�{ޮ51�٘��[�T��1[BVa=x�b�0��{M���h>

(�d}�Th{���k�X9C/gv>�HH a"��n�܂C	��i�����V�tU^�l�|t�#8ieZ��v{�ٻ�{�%-LH�t��U�8�e*��]AY�3�M�y�p&���o\VܱMfL�*�׼G�^��0��gY�4r���Tw��Á.qv�j� ',:İj�-�h�A����M�
�X���!Վf�6��LK�]sx<�"�`��^@跲�fӪ3��Z {�q����1P��ţܭ�K��o@�Ƥ�w�0�_`d��B��[{N���iCyagt��7��yj�8RK�G�U#���Y���̢*'��Rt�L���v홺pi�CH }��9$FVo-���W��{؆�k�ʤ��@�OTfN���I�ы��U�p5��G{Z�z�DЉ�ԇ@�!/����q���A��t��'�S�[.�ݨ*�+�����9�1�ԁ	�<7"��3��r{V����1�$�3�</
zwWfE���t�Y��	��g,�h��U�=�m�����n�Ry�ꢺw�S(�\�)U/��Vv��\f�ԥ��S��_�qI�@s3hx3�-�|�K�`ѓ��؈4I�sX8��Fƚy��w�fv��Qd쥫�҄[�b�Em����-ڙvw-�΁j>�ȹ�:������8E��H�bJX�EҞ y[֝�-TL_T�ǣgn�s�s�݈�m�i�-����Pȶeo8wj������Q�W���5�vK�	]Ee���c��Ȑ��2U��|{u�魫���בн�xr�%mWr�̅ ��6�_���B���AԧXn�L����{�:��-]nZ*i�W�0>��׵J��ٸ�juh�|Rw�(�ë�V{2� t���a�v�m@��n�<b�c�# =B�66�e�
6�ӎrp=�'F�|3K`*���?rj��)ѷԴq���߀^�=0m��ّ�L1�[HZ�k��;/���a���m��TH������$�Q����v��Ї�}�u��c�6]��;g)�BP�󕐑IR��_�^FE�e{��с�N�B��N�V�Ars�}O�&��c/���xz��y.�W�� �X�L:)��<�XR6���d��[Gw;�3J�m,  {N�9xB0Ql�)k�����T�v�)�uB�>�Z��{�A�;2�Z� ���ݾӞ�V�ɍ3o�M���W3�_Y�[OY��=-�X6P}��d̶�^�6�?z��:��H�mr���4n�f*��u��6����s�u���;�(�p��9	�$]8������ʉ�:4��u`:�j�wi�j��r�ロ����^#� �L'�U@u�-j���E�-<�t&��
�YB�ʒ��'��F�YV̡�q
ؕJ>�����u���c�Qǐ�zJW�1AM@�m>b�>���xa{J����ËOru �� <N�Ůzj�5ss��^��(�P�M���{��m�ۘ�l�&� ݗ�jܖ��+�+4-��3�Ud�B�֕\��ƻth�$��/��_Vl����,�ss��^{�����\}G��t���*�]f.�
f��꠵��%��|ox7ev���F�3Ut~��gX�5(޷7{51��$7��̪����UL'''Zc��i݂��v2F8�e�׽�J7����!�W��%����@� ���,Y��+/,"�	RQ�Em^�� �`���g��ko�9��ܐm�է����b�m�|2�0�r�i��|>��Nr�u�5.�F���Q�c|��zm�;�PB+��6��kM=�tG#���{��0`�أg��#/] �K��"��t��o�V�f�]���V!⋁XZ��U��/#�ӱYj�o�-%�z�O���w���E��C$�,�	�#sw�87T�<�'Z<�D�*������÷��U��qs�y�@�Up(��s��B�%�c���ε[j٭Դ�^��#o2\eb��nw���6�������{���@��t������)�\��v	��j��9 v�3��DB(m�LyJ�;�F5��6nY̼�S��`I\�v���/����Gs�,Ȕ�$�R�7:����;7���oN�!��1�x�>�z�#�[��r�.`Ɔ�50��9��U���oQ�уW:����-���^���(���+ {v�X�׬�b�V��1���3 o�������5��� ; =Ϻ�feǜR"�ڞ&C;J	6w�Ԡ���9{g6��}���v�!���\p��#˦�uuA�;-�ovES�-����ި%٭1��ͰZ��{t��
�>;˲��O����oi�^�R
���I`�s(�#Y�5(��Gle��9l[�_e�zM��;�c�����Jo▊�.��
�;�:t�M�ͺ&��Aɇ.���Z8n�s.پ{R%�Ź�oY�8g5�*l��#U�)8���W�.��.��Q���u�L&�H{76���p�E�$��[�.�˻,v�w�������]��);#9Ķwa�6��A�F�/�2��n"5�(���"�\j��rguX���N�ב2���&�D��9M��˵k���9�[��^�Ǽ텻/���pd�k���g�M
4 ]2�.�t+�d�Dem��pU�ѥe�뻉�Rn5���X�bv��Z�ዚԯ���[�q�<rd该��$n�q�5:�Az����e�s���N�\��v�O �EZ����4jrk<���F��R���^�j�H�kZخ�XdSo]�mn���]մ�W.���I����׃�ѬYW�񗇀Kmh��^�6�y�lq�w��E��O�0_cI9j>�K�N�ΰVب����+Uk���鹪N�8Z늡�kD��bڛ]Ȣ�:�j�r��#���y���lc��1���{�!eJ�� _
ugX���h��xL.>��@�NIf�`�y�	<D��5�8L����檲��J'`�7\��w\�Q�}x���kc�L|U1R���HnЫu�g>��lݫ�����(Ծ��b}�n�j�{dGx��-e���*v�4fu��D���`�G�����ଷMV?Z#��]�]>�gjZ�_Q�A�{���R�4^V�e�YU�=)�	�@��9̤ɪl�c�Cw0/s�r�ܺ۝q���V]�t���v��hEh*P���� ��	�f�dЂ�z����݇��#����l�e>��q��C;�����  =�{�)�������/���b'��k�S?tه��y��7��H
i���"nHp�2�q"^m��LĤS�H�"ٹ����qF���;����n�2H��	$���!�QPE3q,���QԴĻi��.����6�m4��\�tq9�q�Lsh���Az'�nF�hD`5,�����u���5��n�2�.�T��LAD�z&Kl�R��u��Z�㙸敮���۸4�M.��|���M��2�ѹv�vʚ>D�-��Rl�S���e��h�
L%�B&�0�r/(�/�A�A�a>i�b2Pڢ�H�i�%�FSL3?��tX	:�]p���s2�ff��ݥ�9rV����kp�s��q��ƥ��Ќ��##BHbRLe"In؄0��)!c~��*4X�n7����p�7M^:"�7]ۃSn[�<�\�<ʩf��nTݩ�\�Tpv�nlܵ+�m�un]�f�-D?�RU6B��eTmQ�6�a�#d�\q"Ï�Q�_��t�R>[7x�TJ��ح��x�e;,g
�z�e���Y��\.^�Q�%�5#���E.<(;�Hnٲ.�5���O���Cu��:R�\��o���#T�}�hc�� �t�X�TҮ�51f��Wk�>X����JqS��5(���T	X�,��x�M�/<}"��,{(�9ً/ov-���-����g�L�J��3��j��	�{)���C�0�Ι�.��3��:�x;�&��Ÿ���I<���9\t�[Wru�1���}���~�(�\�͙$VƇp�;65�NM��i��7<�+��L�ޓ�A��Vٛ��Z����%�z��!q���"����t]�v�*�b'�`m���LR��U��z��@�u��00uG\z�k�S�]{tC���F��e�Ns�+�%�.S`�K�
ۄ��Ǚ�N��ƽGgu<�j��]NƬ1���9��om-�C{p�ʗn��� �U^N{+�����os�6�SG������N��m�8ҩWd��}*�nFcM�lDCh2b�IoР�-�R��b$�'󨩐負^f�e2S0H&��2ӈ�������dL�p���&&mV݆��L(�ͮ��v�47-�3���mA>��q8���E(4ā�Q�I�g���~mHς��m��,����E6��@N�pH�h��	-�d��L�[f$�$�J!7Rԑ�˒&�i��D�l���L��i��J�FeY�B2F���$��w����R���mr�2�[��a%G!�F$�q�� �R�@d�b��xp-�ʩ����uۆ��uϹA�&��M�!I��e��0�%�!@�m�Q�DSq��d�zDH^"�q�'�@��["	.EG��sK�\���滦jn�6��юo5ۺ�k��u˦��HJ�B#�X2'1F�(c������\�f��k�B��J���1��3а��5�2�f����]�4��e�b�k�lqr��.�r�j���w����f��`��"�� ���D�F�M�!I��m�0�%�*&�m�(0��K
-C��0�	^���q��$�Z�h��s�i�S�sv�۬˱lf�
�"B+2��a���!fp�,SF$Q\ H�M�!�i��M �%�I��CR!
8��$M1ԍ<[��L2XUfل�l�6�J(JiSi8D��f@dp��i6��P��ũ�R#�⪁�R�YR3#�0J0�1,*Q5!�eI6�*�!���	} ��E-�(G$� �
Hm6���Ke5��t�2���~K�[w8)3�e�
R��i��D6�)�~b�E�����,4��0˘��cM�F�7k�m��ʥ��[uv��v����]ˮ��-�[w3]-�sm��pS\5�6 ezC	`��!�B�F��ǚf��si�1Z�zΒb,/�&X���*t���u,Ƿ���ƾ5�kZֵ�|hֵ�q�q����R!`h֋�F�D�OSRc5Q���R��3GLx���|kƵ�kZֵ��ֵ�8�5�� �=C�ܐ!<7	�Ξ�P8�QVA`Ƥ�6A�M@��zkƵ��5�kZ־4kZָ�8�ǜ�H�v�gHc�5��)�{�}d�ulC�s�	�+(�hlg�=<k�_^5�kZֵ�|hֵ�q�q���|:��	HY��`�m�.0
*�u2"�
5��ۑ�$�����鐘��J�X�@Ub1REBl�V;lR,Y>ڱ�2�#āk*�c!Qb�°|�q8�CE~�A��B���RH(��I̡ ��+
0�HLa��;��(����w�	QEDDc%NYDB�U\T���!P�Z-�Q#��"*�3���Զ��\kx��Ih��d�) s�0����Ke+P�l��+͹eTe����$*�%�U�0z�/�̓KYm 5s��)a�x��42��q�}��rn���J�V+ʹN�Lj�2�2T(��Ш�(T�S-�Q`�V�-��zB�JݥT�;g{Qz~��g�Q��fs݄=����J"\��f;���R㖪���V�n�w1J廉�M�vk��ۙ�h�]5J��j��er�m�ܫ]3L���Z7E��1��_�)������X�q>h֎��ĺ����7w{��ej{�vS\B{��ۮ��T���'��g;���[8j��m��hNy�!K�U.�kj��eS.����˅��V�GaR晕�p�L�� ID�$�dF�r3#0�B�.�n[�SsL�Q�f�:�扰�g�bB��6�FB�f�l�ȑFg��Ĕ,�"A�blGqx"���P��g�9b4Dl��&��V�]��5��&f幺TZ;n�4�.�sqmtK�`��L�f�sǦ$bFb	��}sv�S������� j�0Jiu=�N�4^���5WB�KMP���F�Zʛ&��[=S�۫�i��T�4	���\9ޅ�tfV��~��!�6�M`ӈ�Z�X�R�޴�E����eh�.ג̟Tӱ�k����WGoS�Sה���@�>W+D���7���}�{���S}ɻy��׮F�Ĳ�Nt��p'4FS�����9S�%���N�ټ�UF�v�gx��2���g� ���C����tF��r�梳LL�PG�F+T�['l�p��A/�+�^7=�J�������8�%��-l�, ��u=j�����3��U��E�}�Q:h�0Mi��,3V���g��=F}���+e���y2{3��y�7FϨz��Gƾ�{�f{:_L�K��wb���k�VW��NKن�����K����wl*N?�[}��u�!�/4�k_���r
c}ܘ�a^εdf���uͺ�H���u����}{	](,`����B'pvuM���W���;r@�W�I\�{�:�kƻ{:J��t鋬=��������z\�ٵ� ��q�u��k��d��N�&�����H�-���kv��d����/s�e�Myf@�p�	�&fW�E2)#`�Pҧ^GS=2���u��=������ -;��'��&"e�"X�����F`1���I6ybC��	�y�y*�L�n�F\�9jB�`�Vڃ�.`a>k��ڍ�x��R�I�Q�x�sĜ��a��#QT>Dߩ%~�4�x��z��m�r��Y��i�RϢ=T/Ś�{4v�֜Eh��U	��V���NJ�UMS��3qdcEւ��萩A�e���JQE�;u�6�/��"��n��J�.�Rۻ��"*����[� ?����7�^�.�M#X��ޜ�W�d�R�U^}�ۧ[NC�r���}���Nk�B�ej��3Hm�)���{�6�1Bn��`Zd����P+�OJ�Nݧ�A��/b���푭�\�{�%�FQgFw��a��H�^�N�%�Ԫ��&
��G=q�Q:�z�,_C�ʥ9��g`o�M뀑��rt�3#��u�/��?�����ƪm�������Zq
#�G3; �����3����r|�ӇbIv,'�"E�Q� ��1�Hq��d9;5�S5�sI+�y(�����e��0�����S�y�3��-oq��Y�I7�?z����\�߉�Q��t���(�>{`��\@.B��v'?1��~�z���,Y�	1Gb����w�Z���5����Tj.�t>��ѣr���5CU�����ΡGr|���黷�c�Bך�4����;��-.T[0���x���H��@,`�0{tp�J	`���m�ڬ:mX�����Ϥ�MWQ��U���\z4+�Nj�!�7�΄�UN[4_t�\��+��v���ˡ��׺}R�����A�Pm�n-<��+K+R�k�aY���^����!,c�-�s6O��t��>Ʌ�b1,���0߶ʩۻB�)����T��^�ԭ�0���l���mβY-ɃW̄�M��1^b�|;���|8����_�N���EO�ZHv�����Tq}�Pv�~���:����r��c�@�y�=��6n�1�VpRхH�H��%̍xt�H��ir�]����W�?gz�B�~K��7a�g���G�+8�%~�mf��A�h'��Rﻵw�iD��w�	�N���"�)IKX�˧V���ж��,6V��3V����|�f�:������Q�H�� ��J�w���K)3P��ǲ�WNw�/��$���FS��-��^Z�ԃ��c��"�*��b����N설5ڂ�s(��Vmgw�W��?{t*����H$U��}Hl"] �R������ET�ʹhdi;�~魥1}��R˿v�B�d���a;����++	F����P)H�Q�*ґ�6���r��6���Me	WE����}��b+�*�P��O�=rk���{�����)xs.��r�v�SD� 2K~����H����6��:�ͬ�����1�������iV>���Wo<��0�.`J>�M����Ux�f�ꥁ�o9ckd}����Vx�|@>>�����ۣ"��/խ��8yG�hq���1�uψ姻��s��^u�V��Ӝ:�5Ӡ�n�HJ��Sf�{��W�mE���5�]���kP��jg�[0�w� j�)G���ok�Ǽ"[�7�šm�yɅ��ZT`>Y�}�`��[%�����&��
�?qѯ�$Q ^��#t>�q`T�X�6�9紤D��1k�3XN(��E�n㬪��O��V��5/� �{!]�?���v������{JIq�H��Y���)uQ���'E�o$Mӗ1��s}�V�ΫU�DJB����^��Y�/��܃�s��6�41Me�Kk_PU2��zO���׫jx��;gӒت\r��'9��޾K"��B�U�ZQ��1�&���<%`�;SH�[g}��uQ�����q����ٲ��O��YN����9��ҒVQ:Kz�j����g�� Kp҂�`.��hu�^[�l��)�'�z9,��D��˝F�����ʕ��7��q����s�u};�YMvE������j�����f�c�iP2��)Wvqǖ�8�9n^֙ o�뽡�Ƕ�&��lH�Aݜ�n\�u������T<=�O����x���ݰϢ��O�O��I�O���ϱ�Ci*Й�I�U^��������s�))���}V���ޑ�ޣ���7ҥ���zr�m4ۢ2<�3H7�"�����w����驗�c�ENڗ����He�I�8�=���2�@���5��ɗW� 0� ��A��F^jY���V�`m�������f�2ɻ�Ov�r�3Qi1z��p-cw~_ٳ�'���X��|��N^�H#D�F0���v��IBBz�[�4�lXYb0
��{��T���=�/��
}�.|��B��}C=���e�[K"�c"I��hD��p��=��w��hXb��L�)>�&�̶�>�����	����v�k�Y��^7���[�S�ٰ-�[��H�{�}o)Ԫm���4L⢉L���ql��^����I���r�>L{j	Մ�z�]��m�j2�:�\�Pd�Ż�FC{�(+KNL�YO�s��:��kT���y�\�k2�xk^��$c�η�K��a��c4ޓ�,gwܷ��Z5�\���Q�!��~z�:�M�]į �ݒ�Пxy� 7�<��QS!�4�^��
cU
.�3�^�/�
6�׈�Q��JI$�����g�۸�TNhȻ����
:�:}�g�Z�P�����Zc׵�W�ݶ�Pڄ�h��ͽ&t�<@�����-�^ï�BV�M�R*��myI���f�Ո@�kp�TU�ґn]
pt;'@ܐ)B���RI����MVM��m�_���E\+oē�m)0��@Bog+Z&+EF*Ո��"N�2��[@�zD{%�[�Eh(�e�YGa�A��9��ϻ��S�ތ�UQ����l�T�����E�]海��mϔ1�f5N�l�#(���^R��ٷ��&�@���Ts"���ʻ�6�T��M8i��Y��c)�Z���}�f�R�_:�f�CTAu��$�=nY�5¶v*ɛ�j�p��L��;�U����m���=�άx��p�h����T<<<=���[��N����і
|h_�8���`�IuD�N�u�6�W!����L�����Z#Գ0����fq�m*�ĽJW�����ُSd"���)�g'�[���S�u�*���q����i�+llu ���r|����R/,�^�i�Y��Oq>MI/�NrwT�GSXc[����Y6d�h֜���Nyb�*�U��/LC�2�L�T֜$��P UXx��Vt���1�*�©J��:�Y�����ӵ��	S�W����h��<�2���3�P��U8s쩫���6��Y�C �"�� �6 S��/������(5/���!�k�n�K�O���YU�ãa���w���z�ɑ�fNX���R%�d]�Ňkp0�1�3�-_�=�tFȀ��q�.hM�lZ$�*��8�j���Y�������Vo�6%���!�rX�xi��R�ሮҊ)���b�w�}�=|�ݬI��lTb�����I�q�������H�;7�5���˧'3�=��dc1�C{��Y�/K�w�w��2l�vf"��M�<�������iR��gY�ޑQk3\�x�磕�6+6��HQ�PK=��o_�۾���P�r($���Ô���'�c�}�[����J̒��v/m	�F{��<� ���H:��}�_Kʕs�6>����f�8
Ja(}%��o-)�ɝ��79Y�b5T� i��)��������kC�d��J&gs�����1YR]�K��8Q�.����A���ϛ#Գ�z���6NPEf�$-o�Y�k��m��kz�וrՙ�~ݪ�{��C]-`����;��[������ʁ
�m����Nÿ�RX��sZ�e�Y.V�K3�bR��'�T�yt����zq�=������{O{�8P$���;./�Y_L��(�'&}��gƆ��r��VR���y���"1��;8e���Қ�"$Yp�N�5��>`9��!�Ü���+7�[��>7�0
�*��x>(v��zYcSץK�����̡[��r�\����2k���۠Vv�s��B�u�q�}d�K��1
���6��������#�$`�b��{��e�ת��^�^�<k�qw�Wg��5L��[���mYEh�}�[>}�r�g���O!�
w�/@��^ߩݴۆ����:I�� *RDG������γ�P��`���F:�g��=�e�v�CQť{l��p�b���Ӑ�g�lҴ�0b(�zܿ�g�`?��2z������9�Ay�.+�����K6�>�A�%O�tb��IjY�iW�H�[O�n6�r1��PZ�7�.^��{:ǯu���D&��K�v��9KZ�@|��ouK��&T������1�����C��-�1v��Kq�0�"_Y�^����ޚ����0h�I�g�l{'��웥7rQ\F���3݅�7sѻ	��=<����tb� ~���u�L����{�㒝"$?�<�!-Z�D٥�Wy:����5�e�0ݮ��K�C$�n�ǒG�r\�P�:*���I62p�9�L�}kjfD��;A�	T�}x��So�w�����Hv��Hqc��7BEh�2c]������)/^!�)jخdݹ#�܂���՚��=fT��"��ܩ�!'�l����$�����R.�<�o���'R7o{o��IR���y�QV�`�j]�[��n6�V���-S�Ӂ��+���bڅO�9 {�����Q��ܒ�b�2�
�,f�+���oD�V��E�Թ��4Iy��C��;��Z�j���LY&��������.��58�A��Xp�8��/�^̻���.<w��xյ�'ebE��0Zγ�9ns$�N��F��pf\��&^�`��&fT�s#��T�����k'X�;{\����aĪ�c!�9�����ũVŋm�[�s�VLB��u	�D�v�j����t�y���E�����b�nf	o7��Jy�HAgt����+u���K	��R�ׯ�olV��ڌB"�����ͳ����m�\;b���D$�9*��v��yg^��Ψ������c!�2�@)1ٖ�Y�a5�?��������ˬz���3@ѝV�gm>�L������Q����,��b:���$�8�;��&�j ��4jTN�N�s��.�;e�;d1�m��*����%ٲF!
�(����m.�ʓ�٪����P�LK��z�63��n��V�K4w�YE�ek�9��l�5qԑVel���{�K��!�[�U[j�3Gu�س�kZǻ+NJl�[�)�v$]�vMUĕ���njw2�=1G}����Z����d�)�wu�� vi]�-L�h*�r���co�1N�(�<Hn�p��WԷ�}��[��Bp`���	�+ZC�)��W���v��Yd�;R�Ķ��L������>��VJ ��p���l9�����o�:�&�^GB���ς���o��nz�R�Y��V��}������ͷ�Y�-/�i�X���V���v��9�_S{���P4[7]ID��ȃ�Ɲ���M�S���^s��&wKY,��wG��V����E��!yHMAfBݱJ_�)���T+�Xa��S��ͷ��z5bYF�_���,���s�d�	޿.�
�9kr-�Y{6�!Iʫ!��D��jvسy��t����>�������F0��.��ܻ��m�;�ӺN�NW���{St���Ԅ�j&m�׿��Z����x��U��йB��b�gTԄ`���F�Clzv���>�?<k__]��������}ֵ۷n����ߌ|�S>���T]��OTRҊ�t*
��C5c,���^�ֺk�����������ֻw2d�}<��{D�,E�J���7�h��.�!$!X����Z�׶���ֵ������}}}}v�۷����<z�Gi,O}���/�r�_�9�.N��&�NP�3%�l���}<k�Z�MkZ־��>�����ݻw>�O'^�_WܬW�
*��E�lU;�U�%A:��&82�5����2�Us)ƨ��u�n���+<��]<�:�����Rkz�� �Vr��3!X�TT�r���"'2�c�J�s%��(,� �\c��W(���0�}Lx���r�6�h��>XV{�%�'�E"i���{c�U���qJ:0���\�	���{�MӚ�����T�g	����<������:t�i���}�{�� ��W�)�r��� "�����p�-}�ux���ג�{�(v�?��x��t��f�jy��������g�-(�
1/��zcb��kѾO��Txh^�^Y��L�/���ꦺ��b��<j��N ",��69|90��_I��B�R�[�<x��;��QM����Z��N�j��{ym��ȸ��e���s&E;����$�TO=�GE�A��@k�V�r��-�x{���<;��aӑ��-s�½��.����z�(~�}����00������w�������d��IR�D�������<�{���C瓫���`�7�1����̡t���[��ũ�7Ѷ������Ӎ8�=fUfgr �<�v@��~|�=�\_�t�GwE�u�A�l��>���}W�1I�-�׽���7R ��W��M>7��G�<^Ƹ��2+���Hŗ5役m��giЀ�]♙h�e���NY��8z��w���jy��Ii�=76{�P����~m�/B���D����x{�;���&��u`������;z��<�9�� ����^��<6P�OU�~��8��o-�`��,��X�$�-]uk5;Z���$��xZ|�S/s'R�YkXy�`s��%�ݽ�fޑ�$�=E����6YZ�A������>�1�;CZl�'!Ϯ��Fw,�e�c,���e�>�����xy*͞��������9˸L�g̲/�5�����n�b���/���z3���7����������3���]�>�B� 
+���'� ���5ظ	�o;Vlu@�(�{�����!�k��}��������V|k@�l�szx�!��c=���j�4����.(  �>|ln�À��5�	�.�Â[bXN��t�}f���~�8	�'�ns��~t�NWEfj��&�֖v��}�o�__��@���J���0��wYd�ǀ�ˡ���,���[Q���.���)Q��1M{<s߂�x���*j��q#�*�<���6��B��%%��$��R�<U���=����_Xx��9�j��`9�H>iQ�U)�J�)��_�i78�_{�ɦ�w8��^��d�בM�x[8^]Ϭ3�pn�C�]��|aԶ_�����΍  G��?_3;̂�|���g���a~0]8�m?'�P嫌���q�3�qfim2���<=��?�x�{c�1z��@����ߏ�}�w�&W�ߢ�yh�Y���uZ�m�~7�J����ud�l�z�iA�i��آ�Ck*Ʈ�W���� ������� E�Y�#�_H�F��^���\���[��<�m��5�c���q��%dǧ���g7�J��$�Ik|nK6��xzx]xz�R2Ĥe�:�ξ{�}���3���|�{8��t��u���S����`N�o��̆���/�d�{a�47͑4t͇O vw�o2�s� u�n�*�s65��	�#¤D/>�N��L�#�ڱ�8^������z�z ��yj�*�Ol8S�:���������%���N#�	��-�a��,�wY�����v�H 3@q��כ}�����.�k��pϐ�Ќ���a��k���2L'>���ky�@���b⺡�v.9�=�i�E��'����E}��4�{��o%�\��g��ɇ�A�֟�̥cu�(�Ȼ7<L�=�旄�I3t/�O���b�Co�?|l%	�=0��x`ې�۸�0��J/(fym�j=� ���f�s��m�s.'T�:�تK��¹��<���� K�f��z{��n4�wx��o�7�����S^��hd	L����ٓ��O���Tki���P-I�ܕ�׼�q��`�w2M?>/P��g]Ng��_8�k�Nk�7��q\���{�j�2�']>|�ƷJ��>ɞ���`��O�OM^gm�˘<�황�}]�m;�Q��f��M��ǀ�M�M� �z������&0�a�P�P4tz t��E�@ϼ�ҝ��%U}3���mԱf��X�l�9���Ƀ�ɚ<y���ڻ��;��kJ��ՃR����T�^#���JUzϒ��z|�t�粫��uM�b[���==��ڊn��z5��������|��'h���C:%�RYc�a�~�:��߿>;Q�=� V�~Y�����d��C�gh~�<y��|�W��[��fq�xx*xOޗ�zj�����7�X�,�����w}��vG����7�p���֜}��"��>��&o4�NC���g��Y���8���WՈ�͌t����S�ׄ*��w;��ZӴ{���`-�'�}`��C����������0�1$<9�j{233�W�on�p�(3�aX�k�t}k��+�1���'�!���^���h^�`&��0lު�W}����ۮxY��ss\��л��m��L#ո�����9�>C�k��#er�RS7��/��({�5EC̻�?���p9�L }�98�{�ƹ���XT��s���\�sxcT��6Ga1��[��w������xl�&�J�N0�s��4`	nK��p�x����!l~\�[�~����}�V䇛~5����{۠�t{s��fj�qB�����z�>0���zj	Ĵپ�:��]���� ������ǿ|'y��#N�?	3霪����}��蓞շX��'ɇUKXuI�W��z�үMy���f����4�V�X�
���-"ff�r�����S�}���gu�����Wʋʉ����}ڦo.BRW��hm�':�҇vA/1��������:���.�W���^�Ĥe��X�Cߞ��9י��u��I�s[̶��CI}���şA���C��7����I��_����K���?q�+s]�,�w5�bX���^�N{.�c�U�� AC����\@�/��2�F)��t(}U��ָ{�����̀�s�ז�~�ᚬ�$�jk��	�� r��>�k�]k߻�{���n���Y��{�(�E���z3h�7�[��q�����&{�Wٙ���x��\���r�d~U�@��~`�^�m��`|�1��y�8���^���y�
cu<�a]C��Fg�� ,�o�#�iё��lk��ұ�<�&k�-��0���#3*����E�v:FW�����<7k�c��������|���=�T'�ve���xM\	�̙�.�ǃt������yojN7�{6hz�:�����ul��,����9�Y�czڙn�r'�u�o�Q4����)�3������o
F1�S�<'��3��<0�q>F��m&)�޸��<�\�-�F�c�o`���Kx��%W�P
>5u)�ڀ��x��Um��"��H������]O{�Z�9&�+ǜ��joi��72��z�b�L)Lb��̹8v_/
t\Y��3П>���D��7A��ϊ������޾
�|�(�_O?<}cH�FX�d���y���|���Ls
o*`
h����T>�.�t���� Y��%���cƾS��o{���tI��{Ň�aM[��N:Fy��S��;\��LdWp�7��w.�G����ߟ�W�����+7M`Ãљs֏�y�G����S�߈�oA/�J���0�A5���^�s�>��w��~S?+�ک��L�if~�5�7�y�x�|�C�j��oA�Ѓoj����1���ق�b������<�i�����-G`�v8r�����:jr��da��!i>��� ~N?Hh}B&MtT�]z{�ż{��Ū�q5��bt�=��`��=C����A�#n��n/��i���);�D�~��;���
�� ���nW�~�� =F������C�\V+�?������������`}�^8�1��MkO��L�2v3p5���*���O�F�gHW$�}�%��o�n��. �3��W*��f�0	�뛝��:������y'�zЍi1�V@�t�0[�<���0����?��a�*��VC�^�V���I��ۮ�v���a�@+���Y0��-���vn3@��U_���D(�Gz��6�EF�nv���s��*��:>V�s� �j�^W6/3b��܋�������9d��䆛��FX�2�K,���I�w�����:~f��%�IIn��[f�3{�!�՛�k4�ҡ�!��%����
�N�h�vo_��Y�Weh�H���������"m3@Z_{�?�@����ZF��)�e�
�v� �O�Ҽ��_��%�~�g97��]��j(&��浃�<+���]Ju����c����T2�����#"�qf�ɧU���T��q�1h 15�v뇳��������`!�s��x)t�l���:��7�u�7~�Ho��r����[�[hhjb�=��`{*��*�2ݱ��I��k�G����xo;�K���{���<�n�m������� &��:\d ��a�qE�YtM�<Rȇ����9z�l���x��i��CZ�� ���t������3o��K�Y���<�c��Z�OO�
b����^?���!�������q�Bѹn���,�pL����������oO�{Q��f��^�o_�c��s�����`��̵Ƴ-�zư��ln����aL�M�����iޘ�8M8��k[��9o�Qت��P��;`SxD��g���R2}q��Czu���E�'�N_�7�(� �ӁN�a����i��Abz�m=�׎��0���k��d��o9C9���wv�M7t�{�g?U�]�sw�p�e��E�R$��5]J��J����q(w^>㨓SGX��Cݭ���4�i[:uN�J���n�#>�#,JFX�2ć��{�_w�����*~O�&~3=sr������tw=��ŵ�p<B�Â�Vk���³��jj�>p���8����i!�;�7]����[9��l�?������ט� <�'����ޡ�����;�j�y�)�7�z�\Fy 7z�K7Sר��SQ	�BY�g�/������e��r����I@���f�!� `~ <�>�����ڝ�`�+��=��Β�aM�G�ǜ��]�Ǻxm����>���]�]�xqtt�2<�6'������[߱��4�B�3�P��3��@��!4�� �Aظu+s�Ul]�V��ȫ�2Z <��zh��X_����DD�ߕ�+�ш@�?����[�_�S���cL�>�����_�L>��wR6)��@�c�!���K.Fy�r�-�Z��mUWJ27*R��ܽ��=��~��^���[ռ0~u��ã@��p��<�/F2�
cY\��YK)Y3�����] _��ӬP�� �[9�Z������$?��Op��r�ҋ�3fa����><z�/0%�b�$�^މ��u�ШvĐ��T��k_�*�^? ���'�f��J���1�x�A�b��A�4sWf�Y�w�0�M�"��W\݅5+�Z�vv=��ޯ��6�|FyFX�FX��Ya<�f����N���������쀼�_[�-����E7O����������9ָx
<.h��k��z�gq��ɵ��߃{�����卺.0���:�ڛ�LW�L:�Ni�y��p�@�%�T����x��*'��< 77����G�59�9=�}j	G�j3�垫�ٞ]܎[M <XSӷ���\c���L�~�}�����s���]~Ǯ�C#����yW�Y�\�o�$܁�(F����I�m�|�a���ż�Z� Cs����6skhF��������'����^¸,���4������xEM �'��к��6v�
��d�쉾��\��;3� �:��UϽ]��rk���o���j�C��&m�gp�@	�����پ3
j�J�=���U�%��Ƽ�b���B�EQN�Nm&<%���Ӹ��:�����M�K�H�I�C;���Xu����bz����߫ٞ����Dy�_�A����O=��K�\�v�3��kdx�=3���e��ok�����߰�{-���}��c�F�ָ��:�Umż�ne[�YBı-�v�vU���t���d&5`.gu�6�T�����;��;`�ˇo��O���{�Η�g2�6�.�.d��B��o�h��v�r���wa�����gp��ފ�O�?o���Ycc,e����޽���'�U3�������P+�R�C���������YQ�!����'�lKfЦv�A5vV���.Y�`�Y�ڷcä^����u&E;�oM��iQ�:/|�	��pu����x��z�gf�p��ӎC�ܻ��L>U��)?ʂ�/�H��}c0X�o�Y��F��3�Ʉc��j��}�Zuφ����A;8�ĝ��5�?i���h5��ٗ$��^���׿���!��OG�T�0��* �������@��uϹwO0ϗ�w�f���l8�9��%���_���@��C���@����Z@��[��6�p��{c�[�1^j��AgU0p��}�͎[�z�҉�3��wΙ|�'�����" �1:�Ҙ
�Mo�U�ML�w�Nv�y����Y�� [���%<G�G8�?v(ghm����m>}v'/+Ѷ�yv���xϱ�X��;v}y�s���l;>�ooHT������?�����{Bz.�Mv��a��{z�SUd�aX�Ε@��y\���
�`��D�� h�s���w�ξ�]o�7��=iLF~�.����-��d��Vփ��Z�/���8�	�H;4tYV[A�u��s�����5Yq���p&�w:PRwZ��>�����=�r�%gf��gdQgt�r��6�7���q�=��r�L
�'[S�����໌yj Nt�f[����i�>��A$A�K��zf�6"�����1��"�Ciח�28S�/]�ޱ?r��gk8M�4|������V�2`�¬T.�Xۙ}C2s*��FI\ ��^�cG&j���o_b"�(b[R��t��9��l�t�VK/9��G��+8c���L�Z9���������.wguA��`!�0ݸ�	��z��>;SD���(֛��IJ��N
��н�2�u�	��X��4�j��W����ݞ|�G���.�V}��3�vT�k��H��h{���[��+���E��^	�WS�Yٽ��������+H0m���Z�6��K9�4+�7��iS;�5�Ł�s�������EV]ƪ7�5v���C�2��6	&:�˭��K�D"�&lDoJb���a]��R�\DIL��ΦO��i#����b��+��¸ئ�oi,~r$74znֻeФ�j6�a��XN�.<��[P�Q�"D�!�q���kWQW!�*9��!qI�%'�8rYvӴ6���T��J�V�ճ�^d�YR��=��Φ{��{3,X�x"oҞ�)Q��/O^�Q8�V��|���v�) ��:G2	V�^P�����9ʰ;)��=5�a]��⹧��ѣ0�c��779�F!��%k�+�Oi4�!������L[2�ni���[ܴ�C��X�K|mu:ִ����y�G�c��X﫮IF�[���vbs���������,������s6�i���c^kF�f��Ãvk�yn��g�f�6v�5�Hٻ�����];���Y�9��냇�Z\��,h���G���ݧӺL��ϸ��X��R�>�y��%=yC��2�+��b��J(���U=�=[Ztؕr@���n�I�t�:uT�,�&�0;	;�;�u�=�9RK28I#����ns�����KV։0��3s��w�P�E�[؋��鋛&C�Ԭ�k,�F�m��>�uU�u��.�"��W�:���(q��4��:��S���8L3f�1�>7�.�;�ww9ݩ&۝S�y�#-N#��:*:����E�?��hd��v�p��6�V�v�W�`�	���ɨ���ӷoO��׶��vֵ�k�_X�����۷o�od8N!�|JHe�Yʍ��Q%Z�,ѡ���ɩ���WԽ͙2u6t����MkZ�kZ׶��}}}z�2d�rt;�dz��+
��㙡�Z����{j:�:��Y��1ӷ�><||}zkZ�mkZֽ����g��ɳfϧ'S�X�Z��X6�
����N�x�fdUP0��Π�{qǎ=�>>��k]��kZ�ֱ�k�ӎ8����\�Wxŏ��3D��3D<�O;�2�o2���fY�ɔ�P���1�ÞSyo#e����/.�c�Zܲ��N!���k�Q/VuB�YP�[��ј�#���S{�+e�E ��gmG��<�l"��OY��r��;�;n�*��i��Z7�ʣc;eb��TZ%2�i�Vv�8��f6��hUwR�W2��޹�����Θ&4�GB��Cf4�L%-��M�!d@�������<�	bE���SFۡm�(�L6�LÆ�J�\��@��%�9q
�t�g�s"W��.�J����0tҵ;s9Z�<V���:�ճ������S-���~�M\ح�Թ�ܦ��k��tr���51�#BPM�LF�/�G�j*�"[e�����S1�LB	0��T�u�p�:�F���SDTI���*B�1��Q��}P1b2p8�l�R.(�"n��!^L�$Zqȋ�^7Z�B�Kv㉃*(�b�j�6���˺�_��y?��3&LrX̙��c2``b1a���?�(���~� ���"�s�]��y�=D紵5��5��K`wY���/\�{i`q.�+uՙ{+.��>�Ya���) f@���+iQ {�����?
�g�S������Ɲ���ަ�4�+��&�{ƾ��<�D?�iϔߟA
�~{2�[:�}^����wx��H��߽Z@�uL���j�o�Scu=��pΣ�l�``4:�\kzX&�ǃ[�^�vرO�gu�t3�)ƛ�=��p�w�G�<�Zb��p0/ƚ��$[~�	y=0϶2=K���z��3D�n�,�=ӗ��@��@ ����{��������қ��9�4_����"�|I��ۺ��2�W��R�=��Z��u��C]z��`Ԡ�L޻�E��`a�j@R#������)�O�>W7>Џ�`mN}���CT�K�sSX�5���T=����B�zk�Vk���켽(�f� �#���a�s�q`Z�.�H|p?��u��#���ezǕ�e�ޟ��e�I�R����m5g�	J�c��#ܕx�o��	o�P���õ��~Wv�mM��E���u�\�� ���L�qo���ze�v�����X:s��W�kL;�@ oԃ�T<5�}�v�25��b�kq���p˂��K%�w��B��ZӼ�3��o^u��� {H��`૧a}���=X;���3��7�m%o	1�ͽ쵎'�t��&d��w��w�ߝt[���,gS12X̌��f3%�۰�@	�Iw����������X�2)��]�P�1e����kxa8���i�a٪\O�
��ѣ����<�<�<:��_5�{Xߛc�Wg�~����yh�r���u��������%���<�m�<�3<= �Kp�惐������1׿=B�%�}=ߝ�U�K'�ƽu�|9R��o�ָ&��<2akz�5����O>ԙ�5y��'�Ӭ'���rJ�Z��О�	��B������ܸ\����z��OQ��pͬ��z�������<5�E�����i�jߣ�
	�zf��v��`ϙ����8-p�Rj/l0n�`0o<�����!ٺ�x&�qv�_Ui�X���H���N��
��o|}|�=0?x���0�/���=�-^�1~wM�j�3�֧�b��pL�{�p�f`$�q�O�-��=�������D�P00g�2��ZM�oH�y7{��=㘙� 8��l����~����x���U�r������V�@��s�c��#��"��w�A�p���"/�Q{i�Vo��W�|}J��/�	���| �?�����;���,��h~��O�-:�ە�P�X��v]�kv��˽��G����R�vķ�+5XƲ�/�&,F(��E#����6[�cǴȓ���v���g�۳��w�1�%���\�W��e�qN�EOqh�`<�����N����y��N��;�=���:�fFd�1�3&fFdɌ�B,���K�߯��=Z�u����95��>�*�� :@~*��w/�����@h3�6���g�Pv8Ht�۶wI�Ƚ0�/�l:ޝ/n�y�C�]���@�O��߫�;�@� Sy�<�(9)���<w�1���q��g�����@F��<2��p �r ��Ǔ2�]���lWKMa��+��kn��^{>0��l��X��C�s@���Y��{���w;�[['���3>��<Ɛ��1���9�-���$xyDSw�9�;�d�	��İ�ʞԎ�\�����_����l�~��9��}}��a���k�r]>�,t�<�Q�g!�$s[lNq�y_�;��?���0��0j	�x��q��syG�����>��(�1}�z�¢����8"�d<�q9瑼�7��>sh0g����O�� �#�؜��f�dN���K p�d��l�gp�`;�[���@�4�zw��\��I�O������dds_{�r�|zc�}s�e�m��(M>��p;�R��LM��g��g�O�~�]�Y�E?6Pa���ŲP��:D:���/CUxXao�{o����2L�N���K�R��]O�̒,��OK�_�hL��,Yգv}��tL�I��C[�6�Y��J�<�.m����a�{+�j����1��l��1۳rGn��۽��ݻ� ȀH
���s�|�x:sO-�S�^��]m���m�r'^�xl�xm�C��f�n�z�ʹ���.�@j��C�z�� ��]�훊���r��LM��+ԫ�Zv �ɡ�7���Ԭ�����&�8��~��I�`i>���	,�ﺠ6��#�Z���qO��0��Ih����K���k�۽NL��Q�[���u{B��7%e�ܮG�I��&H9���캨<����W�O���_��i�/��e{��W6=>��X�p�KEa��䫭�h)��|^XsY+���/e�U��������Ơ�yP_iT��O��t��]��S"w����xm`���=L����n��� D�LY=:��aD�����F�\r�yi�OuN�>�c��Xs�����
�����p[Ac�U�k���Z��%j�4K7n�z��Uǀ�`)܄�榄��`a���&���ͭ��}	tO{����*eJ�n寻�����c���:��8C���jRtf���n����;5�r�М�Tb��Ζ�Q&���Щ�ă�0Q��[E���˷��t�O<%]R�I���l2I *T�m`�ʖJ|;pwub��gmr�/M[Z�$U���l�I#Μ�����y���e�ju�W�k���5��6���&K�c d��0�@) �2 �
Ȅ���2��g[C05��Zn��Cop}q��Kܜ�v�1���м�jJ	b��T4ʺA��Tr��kԫkGl�w���c�C���d�eIC������/W���AcOC��4���<��j"=>"+�SȮ�h�ڃ��z�yf�L1n�<��S�̷�=/�w��D��x_��_�����ۇb7.��/�O.�^�����3P���M>	W�u�?;�G�(�y׶�G8�`��Ii���qӢ<��UK����~JW�W|%�� �{(�/���6s�W��J����E;��`�gg�>d��==={ۋ��N�xfx��q-����=��+�t�os�`}�m���L��:i1$EA^�TX�Xy�r�ëjyؙX�����tn���n*]�uߣ��p�ɤ@���n|�w7���7s�X��0�k�%����n�n=O\fa=\߯o�׷O,�Q�wG�<Uߝ}�3�S�5>ƀ��\��4�*v�uy�}����7�c��3?���L��S�-�{��K��3�E�8)׿ %(o���R@w~��>���{+���
�A^��,��ϟ��|�k�;��"߼����D���~:<%��-�H��v�S[�V�r�<��ĸ�uE4s�q7�a uT�Ā�a�,��[�l�I��~=��"�_��-���^����� ��|fe�!J��@c?����S��/�~?c�4A�ĐO��u���1{}����/`��g�뢉�����r]>�
ٻKz���g���81�c�S.C��L}v"i��E4�݈�v�n�Wp	EP���������E���Ʀ5q�4�VȀ��-��{�ݔz��/	�>�l~���aY��t�pX�� C���z����>^f|��p�PŠ�(|B���
GoYq�6q8À���QW"���L�W�5���)��z��{g�������F��Cu�/�h>���@����=2���zՄ�&�r���p�'O�x�} �8¾��Yăf�>_~^C�Kch`&M�B�ҟٝ3�Z{��aǔ�n�o'���t�����]tI���/w���P�8|d�w{~�ee}Y\U��Cw�Ƕ&B�)��yn�6��~ߠ�����{��T�kjraM�������^��H*%N����R����������x���w:Nb�e�7�T��]E��+)��6��P�o��ݚN9�p
|�N�ٸ�ޏ��a"�۫��WM�v2V���]����<���@7[۽D���_�o��S��9�<p�:�9��/��9�����LCw1��D�h�<�y~7��������B��8��g�~>�����P�����Ʊ��L���_��ɮ��WIy
���]"s�-֎�H@�����v��1��u��9���l^`���H�R�Ԟ�A.���:R\�F��ó�� �_]^�j��Q/t��<���^^^����OH�����dfL�����d�!2Gn�M�b$dD$S�y�u��u���~0��X�=���ߊ/9��~$O��~kq f�m
d�!�c(gNN���<Y�NY���I�?�k�g�^�=>�	}�A���c������2k�e��yUi<�pM��W/����uo�̡���u�q�/v��8�� 0o���ަ�=�8�]���&��M��x�h�?	�޽$'�/˼���gւg (�kƆ~�7�1�7C��ѥ9���,��J�h�\��[(~<���������UG7�C:*E0y�Hf�r%��({�u��4z�����</�/��Gôv��� / q����Zp~a�}ͭbCDs�+>y�ę�묚��~����8*��5��\O��ie
G��{Zi�S�[�p@E�0���G�]%�ۣ����miTO�o&[@`)�0�:�zK�P�c�U]���y`)��k���y�fJ�-�%nYs�p}%���n��!��+5�-�t=�o��G� ����1>}ǆ��bz)�����)׻�Z��n���;r԰��~4�l�{䧧)�+��a�f���>�gN�z�P�:�lM��K�h����ڲl�[tQ<메�BM�/��S�C{k�0�ܟ�3q[��x�V�C�_���<?eB��>�����@V��z�Gr���-oV_rE�u�fcCGn^��9��4�# 3{I�'r�;�Z��\�k{�QǶ=�D;c�i��*���Q;c�j��2�"H��{���}����w:����w��8^OM�|�??���8
,T�{�Ps $��>�&jě_g��r�w������P�%���[^J<_��l�������~�Cz���x��R_	��I��Z���fd4FX�Q����yH���6}��gz܏��a�����j ��gCs�MF�z�v�.łe�Ӭ'u�'��/�*�E7��h�^5?q�Ʃ�f����{���mp!�y�LW�|he0y����ou�z��V����~ܓ�ކ�ۨ�pL��p$C�qz]��"���Q�3��=,D؀U%@/0f��-Щ��p�l�;�m�w���U�<����:�DK��a!M���E�	~`;�@l�\��f���eJ!eoc���ɻ��Z��"��p��ތymo[K=2��:Q��Q����<�t�r�����[;|�u$x&�O�2�nG5�e(ma'�O�x����A�c��er#��o-���]jp�@y4z��k�9�A���75��9-|���Ӎ<�Ky�0?�y��z;�v�:�� ����Iէ�7i!+)n%-�"����!j��n��*��A�m_WΌ#ś[���*�ʪj��� {�Eu	g1`3��9w��J̼��-��Q�#��"�G���������bB����d�H�c2dTt�݀�n*+"wק]g���F�������w�t���������*泺3���9�o���1�W�ndZլвw�]7�jP���9�I
�%FS`��߸��.#r�����EX�9>�5=��X$��Q�p%=�^w3�v��ٳu[�d�Ԙ5�����|Ƚ��R.5�Cx[&M`ol��N�WP��8�� ��/v�5���� �=�ht{O��9�u06}J����οBli���*]>�b��S�Ͻ����M����	�H�~���q�7���"a�.��7�9l�|��Z�6��g#�D�<@>E�81�z|�Q��)E��,G��}I�_�w~��z�Oy�5�/]e;���{œpOͭ>�y��6����a&��4�F�vE����v@���G�8�e���xy� ���<���-�鷭HL��?U��ssP����_����A�����> g�M�Z)j�̎X9۶= Suz/�ޯ?s�L$z���V�os	����/*��6 �p`�kݓn"�<^��5{����ýa�#�a��)�@p-�ڑ]^x���{nO[^����oKy̋M�;�gu�'9���ߠ���/�����E���-HSq��1�}C[%Ʃ��1�코����6��LϡG!�N��b��Nyu_�K�'�up�Oהm�������pE�����@�8����G��u`��u�G{�7%���{X�s�&`�U�w��wS�՗C��F�q��y؜��xxQ��������	"��1۴Ӷ;v�v�n�M�A�@	@�Y�G%�f�f��|��kH���@�k�@Z�y3��ቿ�e��������><�Ƚ���J�Ea��O䟬i��;������+;�xF�����q���\� �X�ig��;I2������*Z�ŏq穏�P���4;��DcZ|��^����Nx3�}~{W�N�3�[�.�[U���ޛ��'|������[sw?�[��2#��@A��y��xȆvk��#AyOG��唶�`I?d_���1�o�7j���u::<�@��|����mC�G��E+Ӟ�n��*OQq����sC{���O#�������+?���|�ڠ4@�\f��ؖv�W_Y9��/����2���[���g���w���q�8Q�����I�U��,
�h�v��M�-9=�S���A������y�+cgN�/;�z�gē��������/��}�_�)}��?����[�������U��w��e�(��WBAN�w~�cv��B)n���{g�z`p`#3��"�i���5��r4�M�zF�3��fV������Z���c[�+d�;�����(��hFv�9Q���;U�Yj2��=�I� ��uda"�A����*���w����X�L�ub�ڣ/;n��6�f��T�̹Ӵ#0�4ƶ��8����`rr�������� �#����c���ǭ�%���Ns�aLM8/����ng.&�SV��\�]��7/$#���u�*�x>�9�#Q�5�������b�t8�)M������S��>�2�f�Vnoe��
�:�AͩrT}{���U����T,���0�o��.������!<( ��ZӮ�+:i2Z���Sa��U�R� �)�NX��z�T��%?+Wݝ$7��
���[�w����ˋx)�b%oI��N9MGnQ��8�:����L�/69BTD0�FwF2�v��'<�Kc/���a��ԶZ��P����ۺ-���)�D��HY��I)��݉���eU�l��S@��C��[�gi��:��=�ktR}��H�-����z��r�tj��z#[�B�y{�#T�'s�嫎o]���#Q�[�V���`�+b�&���7�x�i�2��=�-�Ck����-�b�q� �-��:zleAVf6°�YB}n�%Zf�+��qOb�e*Mz[�jmfu��+y Ar�N6���^�t"��T�L7��aU+6���2���.�YH�8�K�s�Z-����,^��m�)c�VXr�`��gjwX^��-b����p҅���4�pK�R��q��T��:f�"*f|3s��c�N�[�|Z�n�{�b�ൖSVi�ݓ�����|7OӲ\{c.\�vʜ���OSŲ:�S>:L����<Up�%�o�{jY��ܧG7
�Yöc����u�G��}�N'���+�9��2�-���T�{V����s��p��1
������:˕�E��s:̾!�ƴ��՗ٍڬ���,غ�����d��/�.�;',��(M��x�;�S|���d����iM���gtk��2�!���us�R#э��桽�����r���(���Dv��
z5�q^t��l��1UӢ��33���,�I���wh��~r����э-I�{1��a����uۮS)�}0�٤5�#��ۙ����B��vd���Μ���'>����Ԓmέ�p��X� 8���՜��ڍj���o�υ�x��`�~���<���Vbo��mB��B�JԩVZu�n��ٓf�N>>�5Ƶ�vֵ�k�ZƵ��Sf͟NN�ִNr�*�P�w�"�D�gN#��aӊ;�i��Y�ͼx�����kZ�ֵ�Mk]>�fϧ&͟M�I��*�
T�-j��eE�ŕ%dW����fO'��o���5�k\kZֽ5�tָ�96l�l�N�Y;A=KS�t�P�P��t�����_Z�ZֵƵ�k�Z�Mk��N8��߰�lw�'x\�"���b��Q2ҰU9��x�]��Nr��L{J���f!�s9�	h�QS-�AR�4�<�)�L�&`%T�U$�e+h��8�%�!������6���j�Gݦ��m�Z�Zܵ�jB�Y[����DJ֌���u�c�fE)e-���P�S˸����m�Z����yt}�妥}�.U�������ȇT�|��=��c�p;���y��KO3�l�8�巆��>MuY��h������-��9չ��"Ub��U^����&��۱Spۦ;v(�v�ӱ 7AVE���~�>����Yd�Yn���?�PC|ZS�d�qm�"���'�朰/�����-��8Fc�"b-\-5���1��w������y
^6�S�N�:�i�$��fO�:�VN����aԾ?4ī%rð�<�����O�Q����'9xL�G|J�/���u�
⟩0�=�K�T��Z�=��7�}<�!��y���Ł,�2U��x����:���k���Ii)*���ϱ
�y���}�(i�w�<�(b�}�w�'�K�Cv]�n���I/��O|��H릑�5�>�n�z����|6�.Ρ�޵�w΋�]���b<�s�:���.�a!>l8�N�����b���/(-��_D��N�{��������N��m<DO�w�z���N8�� ��
 �>�A���� .*4-?%���nhީO�~�^���'��;�T
4��y:~�v������E&�oC�[?��X9ڑLgG�Or�72#�9��<\���w�.E����.φT�MtS��s-����N���A�������j^�ҥ:���y���vHzQ�w�)�ծi�>]�e��R�k��ڽ$�V)\86l��ЁX�'˾*]X�B;�ʟ��Pj�ҧ;�-���(��o>��J�ُ<V{���O��O��jb�i��2|���=�{������YfK0	���B�2Y� ̙,��b��$��u������5���j�Ć� ��]F7^�Q��~�' ��fZܬ����8�9�6s38���g�sS[^���n���X&u��=�v����@��cz�8vօ7J�U��N#"��]5ۊ����{�ʘ�E^�m.}>,�[�1��9��SwwJ`�u���ܐ��~ ��[z%�:@����}q�]/H�9�?0�k�sM�7]��
*���#{N�^m�ϼ��-��o��6%g�wi��:g��8��fܢ�U���}2.�Q4
��0f�����Ը�����I*�����pqm�;����w�y�Q/��﷽"�ح�T�$k|��Uuf�黗O�.@�&�p$e�~|o�������������xi��Y=���Ȗ/��0�y���t�T�g�h`ٙ�_[��p���=�\T�A�Y~88l&.ߗ����ц@�~��P��=u񀱻���e�0���� ��<d0�n�:���y�]����z��7�7���m��0���,�\j�����C�Ր��n���Q�&�JcqMr�J��E�7:Q�-Ez
���A7L�4���h��Hv�����V��]��F�q�f�S�`����c�﫜�v��Nx�(���ځ��;t�Q�ݺv�۷N��D�PY!$�}�ߚs��r�ߟ�5���s;����)�m�[�p�ty�Z�!{S��+�m*ch��e�A���2����%=4w���}A���M'�sz�Ce�0�[���	t��m՚B	�%ٻ�6͌g�`��0�L��?6C�=�'�|�0��p`A3�s*���J,�p��7���0��p�זap[w���g��>�ZH��-�U�S�H��է�"�n����ݯ-�>�+�cT[�\�m��NZ�я	w�b=�Ž��j�}�fa�-&�B>i �y�~�/>A�Ξ��g��Y��.tD�u�������� ���/	�^\1�c܊��o1�}����0��r��x����5��>�뀚=��m�$�
-�T�۞��;:oU[�w���z����}�<Nc�#�f g��%6���������}��Ok`����oyN�����=�,�&��>�pu�j���H���v!�_Z�\�^t��zf�[�ݚi˼˻�0�V�1����P���j1-����ȉ���@��`}��{�fَ���\��������-6�N���dx�#�U����#9�~�|���P�����6*zt]��Y�%����=�2���+��7y�T�}��8��w�
�Q�n��y��-�Њ#���{�jg��K���C	<�)c����"���|9��D�����[{��1��������뎝��۷N��@t�ۧb���̖\��ER@d# 	�����O�ݼCx|�j.�Q�	��K3y�Z�m�77yu�s����c�;	%C����_$5�=�����j������%5U�d���k�f�M�c����o���&ֿ�����6�H$BY���r���=�rR�?=���w�ooM��g֟6WΜ���xu6�SN���L������;K߆�Qy�Q �\t�^��4(��ey�꿎�2���^��k����	V�^<�5��W���|�����q]�>��n/�9�NƬ�x3y7쑌��n�0���;!"qi
�4"X?����ƣu�^.�.k���v��<�^��9�q�����M����o2X�	�+���	;0hp;w���_t���;�=|
�
�Cߐ��B��܃��5����P&��Z�y�왍��a�һN�߼,����E?>�旕�d#����4~ji�C��-�hg#�OSw���$�o����`��L
��M�:P���x�ţ�@C��/�Q����T9��MYOh�t7Q��Un�6P,����7|��[�z=����b��à���.��,�l�����T�a(	�C�e��m�R�pլ����s:I�h+�x�����d�f�2d� 2YfK0��$� ,s���������Y���u)p��A��2�S��o��Qp���=�����	<�;+���l�W���qr�-�4B�;�]�ǧV�F0ԧzC[W8]�͍��i� &V��Y��lli-�`ߟz �[�#"��4>���~4;�sȟQg�q�R���;r��q�9�\��"!y�4�x��qs���Sv���Ӟ`5DYz��Z�����b���jw�tAŪ�5N���+_y ?�y{��0��o���y�׮y��v	���^����Q��"���}*_:/0�B[ ��3��[�o�~���ݥ�]O����.�g�;��E��V��x8��q�=�^�X{�2�w��4�Q,"�H	�:�_�G���8�'كb�����s����/_s�]k���=d�n9%�nz�}okSQ���`,k���w�XQ�:��>󁓨�G���ʟ��;ʳ^�w�@�����O�G��	�dǅHk��C\B&|5��Tz�`��Cip��K�03rΫ��a�U���P�� 0���K! ��#'�i�@��!���V���\u]Q��Z��DZ,��$�k�q�����g�<�M+��r3{q�;5`����H��>�aTUt�n�ѝ�-��J�SR-W9�6�qe��H��x���Ϗ�^�����;�~u����"?���N�H�ۧ`,v�ӰR;v��"�� ����wer<}��.�!� h~/0�\"
V}�-��Q2~T#���� NE���g��}T_�����K�Wdh��(E��^��N��V8K�p!�[�B˩�y4{&��F��C{�*=���T|��XZ|(~��T��g�vz�S wQ���O9��Y6��yy���f���;�{W��ޚD�,���>:�����A���ź����;~��}�������ۄя����/v��N6
p��SvW>�Ej蹛��_O��<p� w?�yǹ����q,�[��f���Q싷�x��by��>��}ە�K��i������^T�U�> _�ǅ�??0�	�;+q�~��9�gd%-R�]������W1�@�xD��s��a�{�4����Ɓ�[ɹ��u�� ���0������x}ŀ6T���1˯������>����/�g�z�|��5�S������a=��y�ע[��k��5���^�ac|X�/xa~4�?t �-�0��������⧜J\�}P�>�W��14�FJLd�G>�ʶ�K�zn��0��)���v��F'��ShB�����|���W:�Aߤک�mw1ڜ�yc�}D7�Pz`ѝ]�[��ݡ�ήk���fJ�=��||t�v�4�ۧ`�v�ӱM�,�f@1�X��w�zf_���Y�j���P*�����ۼy�c	��ڛ��8���r+��Pc@i�F�o ��\�g�fa�C��TMC<OKo�0&{�зL����K��G�˼��4s�	�0a����Uu���i�b�����52ؙL7�,#u��:�uL�O�N�o1pz�\{f�/8�-���������b<�o5�L�����?��n�4�7"K,�|�jx�u[���@��OW�p|{�Q�?�TG�[�~O�������1�kË������*�ȸ^���4<��Ԝ&�U����>^���> *��Q�����;vC��M����|�'�-�I�׺a>�{��H�yo����n�c�a��ޙ�i��~U�����Tg"�����pp����H½N��-��ێ�&��C�q��5�V��z����sQ��u�	��ӁM%�/;T�x_���h������3M��x/L��w��R��4��o�7��ލ����`��E��dwW�yw�&�M0�NF��T�
F1�Ƚ���b��ܜ��i8=z�;6�X�aa�|�ʇ�N�1_`!�Tx��@�q�&3�eo��
�8������8u�do����Y��X�+�^�'��X�;$U�Ya1�w~㇎7��r�P�ݧ�_WgH����7�7uv�<+*;E�Wmے�^J���OS��R�|��M~"~5�N�c�n���n�;7M:v��(��^O/�s�Ϗz��5�O���,EI?~��@�'�N!u�?R%髝66n��3{-�r$�랳>4��W����]�k3�s�~�Q�}�	�!�eF�]%�8�̮����w��1x����2+���zQ�N'��f`ν ΰ�N;�����[[TV3kH��:G�l^o��E�ߝ5{^��6�i�Eb�����&�_m5v&�ǎ��ՃGC��O�;jFe�5�k���nd�u�k�瀥�޼�X��Y�e�%C;��h`�>����&��>���Mw�|��+�w�j�vv,�9��+$�PE2���}�$"
,!������e��z<ݘ�_S�a�61�>��*�[yc�i9��{�3m����^�Cmt����>(Ǟd�Q?+�����O����F�Վ/8k�P����������1�G�Ro��;���K�	�x�$��(^##����������ᾜxї�R_�Éߩ?�b)8,`<����p7��1�q	wzo���Zn��t˷���f{qL���o�
9�7��w䱂g����7C�N ��.z�V���y��f�B�.>��1m�[�G}�y�
m��]�]�5��Ǎt�;v��v�ӱX�ۧ`.�1����ڿ|�	Ͽ��F~������S��/���L3A|a�OG 7V@�}չݿ~����&����n�Z�O�S��u�'0���035����Rk�qL�����>����s0��0�ޟ��D߅ߟ��	~z7��߻��䆮�����޾�i�/���a�o�y�qT��f�^y��d$����o;f~��ƌ��f�&yE�?�퐺�{|���n2��>��r�B"S�W�ԃ�j�o��f���@;��ɸK��ז�
�)�qo�l3^�g������D���j�Q(÷����|b}@8S���i�nA�]�P�1f"����5�S/K�,�u%���G���ƾ�<���o��@Q��qN=:-\�4��xy�}U�O߶�Q��,��M���q|�<�TX�//���G�_����B��:�0�_��4�)۩'5�'v�7�󥲱L0���7!�ټ7�-P�`͉�J�f��~�N���tV��V��؎�cѕd�5Ė"�۸n��v�i��ƻ㽝�t{��ӂ�h�x�͔f:�| �%}���D|�z�DY
v��%�M�oU��8t�%K�ش�G���K�[��ǚ��T��y������w<��k_�K?N��;@#�n��۷N�c�n����2,��u�o������s�\�}@9m4�������1
�\�����1�
�
�8~�ˢ����<v���9lǖ �x��k}ƌx0p�?���Y�0�5���x<��H�S�P�ߩ�}7)����������!H&���s���ދE�3�46v�<���}�b;���F0�~�0��^�1��Gb���他oP��(w��PH���7*��{��0�/.��� p��=���~^<)����z+߽`�<^}t'�&TC�:�ے�ϗ���>�f�8(a�ҙ����/
�A�^���*.�7�p��1��6��m��Us{��8O59
E����k����==���~2w���}1����$��Q����GbD��)�Ru#�1�>���ڄu�Y��+�(Y��x����N=;/[�aE���rܨ\��DxL��8~���T��*���=U"���-3d��C>���ևR�˽(�u?����ـ ##�w���|lA�Xǎ|�)�3��=�9�<Ǽ<< i=L��|�I��(]���Wʷ��x"N�}����x����C��H�7oRv�\(�.�\����!ޗH�wkKI���3t,oGKxٙL�s�Ke.�nGo!�C�v�Z��Y�^J��$��䉛CZ��y��*:Ę#���յ�q���'�9�ڑ�$�)S��j~������YN�ȵ�s��9��d]�s1��Ó�P�t����gX8��f�B�,�$�8%�N�d��h{F�d;��Z���]l�av�#"�=��|}��Mѽ�|�{fxt�3�:]مScJ�)����I����^ݎ\�����% �
hgn�n������J�1�;%���Kk�E���Xx5���7֌�Դw��9��|�U��6��J�^�Gt�n�뷢����`�.�<��M��h�.�.�:/����۫��ޘp�8�b���V�)1���2Ccsw+'v��a�j�}+�������;���q��-��=�J5ԩu�!��Ҥ����R4�m��o��n����rZ8��S��ה���Ȫ[T�:#��^��9Ҿ3V�\���(�܄S�0z���ZR���g7(�%Ƿ��Q�h�lex��F��h��
�K�TR*_)�Pw��Pc����7�g-��ۂS���V��e��>���h�iJ�r��ZQ���-�L�n7�������q_Q�o:��ՎJ���a[��s��.k���s0�sPƨ�V�N�88�pWUK�}�O{�ڄ6V)��-�טt��w�ނ0VZBR�*�\�p��g2n��/l��"�S}o��]2��No�%+����D`U�U���ݻ�t^�8���o.��Ok#q�5Z����#3���n����/ �婓1�tz�;���Y��{���әE�v�`B�j�|��՗�G+�n�Fx���};�p����'��o��
�L!�=���b>�[N���w�'
���],��]�l��{�'��XD�V"I۵yt��G�E�T��-1Qt�gy��"(�]]��C�\�$��lBܭ]��o�U)6c�ns*�v�i�YV�5�2w�*�Q����-�{��5��B�v;kB��X�S%a41-�k9
]��m��&7:�R��wC����|1I���qNձG%Ǚs�;=.E���N	��v�owwo9$��F#������]"��Q�_���1�ty�������U`���v���J�5���7	乛�{�X��^��>>5Ƶ�k�kZצ������q�ǾN�miӃ2�i1�nA[�T����Kh�0���&M��ϧS���d��k\kZֽ5�k����ӏ����{e�~�\r��v��2�#V��*e6Q�*��R��Gf�6�����ֻkZֵ�k\kZ�'�fϧ&ϦN���8gXa��}J�6�KO0���Q(�i^lܛ�n;;ѽ�z�۷׷�o�k���k^�ֵƵ�v�}zq���2g��5�l-m���`��TL�XQ��0��8M��2�¤f6S@���6�vÐ�RH�&R���*�T��ip���"�.i]�ʢ� �3.*�Z�Z�[u�V�b��n��-R��"\1L.\k�Ҋ��m7w��2�Z�;�k�%>���/]b��*&9�B�1���+�f\��P���
��[aZ�ǉ�B�s,P\M�,��3�A�)�v�Ye�%r�;�����vх��ٖ��.Z#�(���S�3�
��M\��ۉ��ܢ�J�N!G*Q��4=��r�z3f��PD��t���X�b	�[���P��fD���!�!*�� �m5#P��3"'�8�.2�IF�h#e�
"B���pH"Au�'��K/��/�t(�`�=N�gR��iXu�s=�#&�:K����V�uҖ�j��X��J�JT@j�IDBl2:c��k�Z�f���.�f��$NF����E�#r!h�!)"&�
aWp�66�[.ѻ�E�ˍnm(�4�n��%܎n�ku�mu�����9�v����7��r�� ��c!���C�e(NFܢra�d㹢יJ���nm��]R��˙i�h�0�2�!?N�%� fL�a ̙,��2d�$�ƽ^����x��O�#��~�m���jl�Ś�Ymv�I����A�3#��C�q���G�,��e����v�Ӑ���h��,uQan���-J���b���b7՞�c���o���T���)�T�f�z�)������-��#k� ���̃�Լ~'��(~c�����?0��q�9/Z��v$Qp@�/\��@��k�:f^q>��^Z8\z�""|ɤ�@e��|C�[]�J�J%i�p�;�]	=�='�ԯ�6��C�&>{�e���1�܄�-zϤ�^ڼ��buÆ��ku�	���7wwP%�v@�y=z�=8~}c�kW�҃�2Tr�>�ݯM����I�
d��4�qy�ZA{����W!\��za�ۡ���.D�`q�@����q��\��|��*�_��0ĸ��b(�Hzka�kj�Y��Ն6�Z�GOg���lѿ�+���4������A��⿑��/�y�]I���:IgI�8n����n��]^=�{��y�g�=	�q�p�vwѳz�
�@x>���zn�؉��j�=�s���ß��BO��h�0�ym��z�<�Ƴ�n�:��g~u_��!�/6e�m��y
�"*���aMp�J�b�M�~� ʵ��]Ж"%bGc��Iy�n��k;ei����5�ܖlשL���<�7��^�+7�����;0�I�E�.�����ӴX�ۧb��;t�M�ӧn��&�'G�9��}�N}�j���~�&�6��|F~C���Q5���#�ϴ�׮�����RUգ�,3�h��M��w3>E�^�O���cOoD���K�ĸ�sk3�/�_�ֽ��{�ˌU����2y dM������y���6-�7˞|�Mb`�N"}�3ĩ,!J�]M,�d�֖�x��C� `T�p�g�ܯ�c�-�c������Хw�mu�p8�F��>5�v��tP�ɴ._�����Pwz��o�]��p�4o���?'U�"��޾�<���X��G��h��C@�e�"��9H�ٝ������v
�=ٝ)=���B�a���;�7��8^�#�b����n���Y�����s����8�y.X��ng���m��H�0�`9���M�W6gX.�6���X�4P[j�F�������9��>c���g��(��W��AJ��ߧ�40�A������~~�L{k �zo'�Ċ��u���=��Zk�����Ws�-Nޠ#NT	�H��|ql��t���>�͖�5;�z���U8Z�	�S��]�;)#�G����}��˽�__Yo4-PP�w�ϳ)u��'p݊��P� [i�D�x���v�ӵ�N��v!�t�w@�^��w����˼ɭ|����I���gL$@�O��W��ffT/���{i����<OS��?��f�Xծr zo�~��0b�^�v�MId��O���;���st�S�=�Է��8��Ƶ���$���b?��ʁ��p����g��e?F���9�ƻ%������� ��|���Fwo��1p��5錌�
wn��U�]�!0�ޭ%b�f𙆓��M]ѣ�԰�v
�08��A�7��~��=�*_�XϘ�w�6{�aytr��u��Ĵɽ�Ǎ�\�e���/��,�l���S����$>_�!-�L7�l-�Գ�������{�N�����!E�t��A�W�'�}��\8554�9�|����6ь�ܽ$��������s�K�[\��|���L<y���g�Uu�^m����Q��H�J�g���^������}���_��\��W��R��E|�ڿ4���~���`?  |!G���9@�կ��S��yw�-���ʇ!;�-�-�k�?g��x�ۇ��+z���W��R@NϫPh�4ܲ:��r�	��Z��[��XX\P9C\�J���|+C2������Nr�;��w%V$Ҙ:��@�P�@�;��H�2�����,io0�w)����r7:ny����͟��<k�`1۷N�#�n��fL�a$��:���}��m�o�� �ۚ���=]zr��6`kt�ey�x�ffd�X���~�Na�[��������ǜ�0�k�:+��/�S聡�	n��֮P����ݮF��V���Re�Z�΁���w�u�4:��}r��/W��}�wO���C�]ϋ$
}�-Ϗ�a�ƌƃV��),/�_����=��f�~?�ζ�D�?����H���U��:8k�_Ue��'�YN'����g������H/HhĮ�%ycl�8У��/���ޗ�k<��>J�zN&�l������O�.����m���3�:@l�>N�t�f=.D>^T]Y��T/�~����4w-����d�9>�u���<��^�A��8�'g�q��ݷ�:aN�o�1�w9�����o
U,�!�����K��g����2\Kn��t�C0�^����x_���S$m(U!ڧ� �C>��q^��x&��ݸ F=��v8f����O��/��~U��w���^�4</s⾙�z���4�y?gW�X,�������t��m��x�X��@�Xnܓ*L�X�9(1�R/�#�4G�!�!���#��������1
��U䢀T��"ة�Z5R�#��/h=�-Ve�]��.��^\�}�������c�`t�ӴH�ۧj1۷N�W���~I�������D1��xd�;Ͽ�ۜ��<cMK1�������;��h$;�w������v�T���b�@[aﾬz�?�?O��P�S��ɷ��}b5yĨf���w�c3��ʮ�N��p�y�[�ȶ��z=�=�S,�u�>�5<!Z���*�(Y�5�7��0��]}���I����E?��\j}5^�ā��x��gw�'��y�XKTzh�:�͂��f�o!��t �@��" -���h��oE͆f"�6�W�Xsp��)t��b.�:�I�l�wh�!�3��֬������YeІ�C �����3�_f8x����[_�O~{}?t��l�3�d���l1e�c�o�qz#}1��hӐ: ����K��f��,�X���zi��>����S�#���Z��!�B��B�̶>�Z�o�

�����#�a�F�9�.'֠��z��4�@+���'�q�gu�_��!w�Η�������j�����7I��1�~	6��Q|�N���~n��	z��&n]�}aI���r�y�{�	!���廫߯���C�!yg�f��!��s�y�K)�Aa��O5{-�B��
�F~�:�&]�53�_��Zst�nK���[m��B�hӮ�Μ3N��p�u�BԪ�c{g$�E��Ԫ}�)��F��M��l`��¾�����[�t0orm[_E�Ggc�&�c&fڜ�Ʉ���cۯ�1�����x�v���R��[&�J��n���t�H�ۧk��N�;E�T�G�y���~��}L>��@��-��O��3K�'�+����]l�%W���k'0yiUcw��_?�Zt���Z�y1�O��$��X"?.�����|��2u}�̔{���e�u��5v��O=��������y���<덆(��n� h_WιX�M�'�3 �rm)�I#�>x�<ތ|���}t'�����y���e;2�o�/`L4ը6�d�=-�i����S�2�=8����>��[3��hWs���wyI��Ux��@�~�H��u�n��i���z���\~e���á�|�ޛ`��JD^��l��ˉz�G�z�<�v��IQ�UQ���]����/
, �򎟧�}��~��ߘ�1-`"�O�SϺ����+�ͅ|��l+��z<�HI0Қ�Q+��.~D��������#���3i����8�/5z��7�Z��|k/l�KӼpP#����aL'F`�s�qt2�?fmΒz�[[�5�.���wWw�$��1ظ}��O1���A|yǣ���P,cHؗ�o�=�ͺ�5�C{�^U���,�5��j�iE5z���Y"x�L<X|8*�x���](Nʶ��c�I�fL��_[p*7���W��������#�u�-[C�Ȁ>������n�;;v���n�;u��}����!�����ۨ7�_X)�怸�v>x�	�Pc"��Skŗ����ȶ
9]��j�o$��iq]�<��WAkb��5��2#���葮�aZ�*�a?T�7��w�����>������||`"�y�-��;�B/�=�|���# ssH�ר���43rήF	���|��yw����9�:�Ə'�2/H\��VIj��A�Y�>F'���/F���pJ���U�˞{Ld��Hf}�� �@�~]<��v�e���K>����5���-��Ʒj�Z'݌#��:9���g�bǀ�����j�m�Z���71�Ut�-u�fv���낹
n1����"f�ם2d��y�>w,����*����(æ&h����5����,�/"o|��ޯ��x�Ԣ����|mr4���'�߿r\i���}��l��'�����4�ߛQ���1�*�'O�9Og�1Za�����{|�����e��S�_L��r��@���	���!y,k�R=Q驊h��
���3��Ae��ˋ��P�+���Ӌ�u��ln^��N�v���hn涳�[��m�ce�I�X���dv����TUb��:�F�ɨ���I�&:��*�a��l@u��Oj��}ʔ�v\8�v^[����Y�g�|��Ӵ�ݺvv�ף���?�xt����ۦ;|-W���o�tQ��T����(�ڢ�Knnku=�:�����l�6�l�^��	�۔{��1qS]c[�E������憂퍲���v����%`���7c&���CH�Ng�o?�*�J^ݞ������||���\^���w��gz#����]�1h�f�ޯD�_�	�8��ȶ��g彦�K4D��V���z}O�A屻��,L�9�}��)`������\�[�@5σ�ev��9�]��3�/���H�ٸt[;&��@�ܼ�<�b�[��w�{b��x�$8�ι\��>�������	���Wl������a!<�ĥ��ON�Y�7'����Sݮ�=�z���ʣy���X���MK
�<0�w�e�X<��}��l�����v�ZQ�!Tѳ�� ~o4x�O�5��4�i풤�[�]E��m
'�'��������ߞ������c�֏��	�!|��P庨�Ꞟ��~�)�4s5�݈�_�Uz����ut�It�plSW+���zn���uT�
��w���f�f�L{e�Ө�>��'\N�/�HI{��>���(.]�k�x��P� ݄1d��rԺ1u������sY��Bwuh�O�,r�_g�S:뜹�y�d�?:v�۷N�;v���n�;o���r���>�:���X ��nd�,�}ϳfw�>�~x��*��RVڤj�|在��t��w�PͶ��}��	W$�ur��Y+1?4O�����{?1�[���4�3�g�ؕ�6"�h�=y��TO^P_�lg���~�m�*�h ����*�5�1ْ}���2��ջ�N{��^��⛙�yw�h���<<��>hln��f�g����R]�T�r*�r�D�6���	��f8=�̾��W������	N�+�����
��m{?q�[Vo3陿O-�j��}����^koF8L��6{˱]-�W}hL��h%�I�3�G��Ҟ}��`M���q�|ӹ�!��jE���`׭l��Ң=��&Mr�9�(�;���eY�G��{��K���9����+�^�M��H�py�됂/���"������V������Z�v}�t�Mz�0�ݟ�~s���x����u^=)����͚�+��"~��y�
ߗ����+Wԭ)�!
'���G5��,�#�I��[��Z�r$�,�E��)t�ŷ�����i�9��}�[3?&@"�:��ya�ҁ�~�"O��j���ӈ�J�a�o��8���/�~P������j9��� �S�^e�D����,�߉�{��ٓPZ��]p{{}E�ob���xIۇ:���η\��N��_nIX4��:Vxk�c��p��[�y��^0?�?�~�/???'lv�Ӵ�ݺv+y����w��=�Y�{����o�V�S�6� ʒ��aJ�MNᘵ4�1�D�|�S;j�-�p���)�'�ŗI���3�^�P6V/WK��9���T�L����4�� �3Gv?~���%5��z �S�~N����-�:4���~n.���~Q�Nޖ��Ǖ���E�?�a�oI~e1 �!��d�1�9����4��؂���9i�u܋a��`�	�P� �T4;'�.�h�2���4_:֮<�ЧvU_]�6�;��f1���|P`I�U�w��c<�>��pE��Dqd������f�(�b��r��w��׎y�cKI��B5⼠&�+#\�'�@��F��z��m�O�j����թ-�dL</�Vޑ������`%Ļ9|����Gj:)�@��}��F2�Nn�k��`rn��M>��u�2}K��M�Y�C�g2E}��N>���gұ3�Y�KY�ڬ�� �n��zj���1�c`LC@���#�P�����	�0�`��/�ҷ�^��i^!��5c?[� �,���r�����O�y+��B�!�2�MU���kqei�E�W3���$�u�V�}��u��ˁ�lro/����Ư���k���rz���\o�ra���Șɺ��7%.�|�9M*H���:Z��B�͕o	#����q���9�}��.�+}���3qX���}��6:ļ=��6cX��T��d��Ny���Uh;U[ի�|WO��p꾐8.�(�
��u*"'M�σ±��K����v,Kº�%�N$�o����Fi]�)��
�ұ��o����9{;p�'��w�)�(��h���<90l�V�-j���|��Q[TqI�:M�4r�;�gF�F�TLo	{ׯwj��v�Z)��x'ڃC�_,��\�if�Ž��r^��h���	���[2��&�����A}�֖�ŵ�Px��J�Y(V^U\>�ʀj�㵐>�k�XD����j�ڗZ�۹���|E����W�c
���.�e�]BHn��}�0���ϺK�D�i�0�Yaɶm-I���k\�q!�4�&���v+C����=��#E�S�uyS�����G���1J��ω��ޙG䦃Uf����-�m!1cob"�e���n�����,��ɔ�yj�]C=affW;S팡�~���ז�\f���X{k�����{l�V�X��e>��Y)n)��W�O�uBW���ά��ՈF��K�z.�6�[�tA�4a�g��
x��
j�+N��_��M�1H������ؠ���[��O��QL5̺��"�7&pF�A4P9�rh��ZՌ�'K��5�Պ]��(c�n�4�͡�Q��	�.;���2��@{�W�΀�;�6��@]���7t�Q(.���&�J��|Ov�BEi�Ko,w�v䘔�@W2j�'N���Z�V�6lu����������Ó�ޜf�Q�m�;�[��w+4e����ft�pF�D菲���L���7OYw��E�O� ���4��"���2�N�n	p��`���9�ߠ�E?���6��'u���Z�[��f�f^	��^-�&s���4�X��2��bH��1���
o%��"i�J�-&i�
���-䅓Y9V��0cj�������'߬�]�U.�ꀛzr���O�(wc�Iݾ�F�ݍ�.�:3uu�t�P4d�OJ��֞�WXn��f�%���kM��+bL�e�4�vtFms��E�d=G�'�q���L����y�[fs��wt��w7WT��k��q�p æ;��߽�����:U|�_��jX�5ե��ϓJ���S����J���R�e-S/�%�;��N�Z�mkZֽ5�k�kZ�8��l�Y��8���,F}w"Ҳ�i⸾u�7�,�-��e1�$��8���]��kZ�ֵ�5�k��㏮>�{�$��B�ʡm��(�PDF"���R����TPm>q�K,���{+���MkZֽ5�k�kZ�8��l�Y�|a〯����#��.Z}�lf8�(�
�>o.��d���;}z}}xֺkZֵ�k\kZָ�>�>�{�<�!"hS�֨*��"��Zy�_���������TUT�I��v�R���U�R�����TPU��gMD�;&R�%�q�2��6֌EE��,E&�����h����,8��S)f%�\��x��+�E�
1�����9j��4��ҫC)F �1Y��̸O��1Ʌ�XS�!�c+:|͞!��Z�+��T�T���N[2"2�zJ!��wh��R��-��S�DU`�"�R����J���`��}J/���Xe���RA>D����Q��`������`���6M���ʔC��jX�)tv ��������Xq��U�߽޿2d�d�fA�2Y���yߗ���jw�d;���~^_���~k߿|�������Gޟ%Nߤ�W�s�?���U�gy����V�H*���{q�g�0��g�JS�*���5���w�p�c[8�v���S�p��>cK�����ߨV��C�VQb*I������,Ls���>��os/zW7]��靰��|WO�����cs=Cu�&:.=�6vQS��e��K�ى�w� ��G�#/���?~�H=�}��nT�EuwRo!,��Av��f��0�ҳo�z=9	�7;��	�84{�oMq@�=����y_=��i>��KRWj��5_u���m5X��#p?8�3\��hY\�M)���׻�����O^�����I��0moD{��r�a:�ȉOI�x]�N䒷6�3�(ekU���O^@A�t0gO�j����PƟi�bwr/t�I(:����ܿL����a�+\k0��G�e������V��>��G2%�C��M-��ۧglX:�b9&"z�v���ٿ=�Gw�Q�W�M���7��l��A9���I|L0c~� ��`�����������8�S�]V%�Q����ѹ���ݕ�a@�?�^��<����������ۧc���Y�y��]?s!��
@8���w0iV*��nI�j���Q��<>3���ob-�P�/��֬E�m�J-����;〵y�%��j�6�޼̻<W�ւ;}>�~�Jr*���g��g9� �S�Z���V�gy�Ld�}�l��A��A�o\v8����S�9o�H�"#��m�$��P�f?��MYK=[��a�[{��73y��kWU4�]'ݎD�(���{���s��Z��P9�T#Y��T9B.�w�!����bİ��z��Dz��@�+DR��Zj M1��*�����Z���~��[���������X�].�UF=�p:o�&�
�x���iB�zE��70�@lD�������F'��ry�$�A7���;��l�S�y�x���8�)���M���������{1UrME,�z����e��ݮtW|!A�sօOCfx�Ì��6�Ƴ�j����WfN0»2��9�M�_5�3�p�`r�]��:VD��[vw��˭;�����q�N�t�Ӳ;v��Gn���vg��r��/��85e��!"�*�M��ܘ���N�/I�x��:'F�RR�׍gl�xb"�i�e�w��g�ҙkd��cK��d�UTz���ﶀ��F��h�d3Cp\G{n�}5���J2^�{�y�ofq�T5�����˞%�'y�F�	����b�ǣ�yΤ�^� v1w���Ǳ���F/t�M�</�%�!^��|^ǈ�v���euU��p!��.��u\|o�ݻ��y�׶z۵�gξ��V^o @f�g��������'zo�_,�:�7h�k�����]�5=�!����tl��Y�:�����q�F)`���H���	�[|��� >�d5������T_)��d����wӕ54Ų�\�iXc��^;�k������F�ǵ�pwB������`6�ŵv�)z5�"<�``��٢�u���~w��V��3���[�f�ю^S�]�������6T��!����^���C7a$��_I.�3�oEV��q'��r[�C
����=�A��ZoS-�i��J�2z�����;������l�}Έ�I� r���-^K�B1pǮμ؞7E�r���G��ɍf)u5
�ݝ�z�v��RE�7�3co��,�e�e%�Y�ɒ�[�$Ʈ�݃O��5ŋ��E7:wwg~}�|�",�Q<+�5�Fy-������&6�E�OeY͓.eLK�
����s�u�S\zȘԣ��H�cدU�^��Q�R���T�>���m���?[@@`�V�G�}b��"kc7s�/vU��p˓y>@�R���cpn���� 7�+�LwG�C�t���̨�����\3�s�f��m<6��+��_�b�L�����"����wn#�1)�R1����n��~�J���j3�u�H��*;��K��-���Θ���'�b;,;_g�hj1{�o���<�쀯��o=�nJU{����l�ה�ó�=���������7��ײ���v�q	f�n�^�7j����1� ���k�c����yTt��4t��6��^�%�ToD�~++�|`�}����;oZ�8����X�uJX4��C�$�CA��i�ɖM4�IU]"�e˜zggm�����|\ށl0J���\�ru0��R����=F�9��S��5�e�U/�*��kU��
��2Z�]�ۭg��w4�t�3�>{x���ݺw�t:t��/�y�3��>�1<��;�w<m�5��n��|RP+پʍL�o���͚�T���;W؉��P��l\���{�޷8��,c\�WmkzY���KI�Dc�<u�������9p#���I�>ېhHU&�x�+6-�5���_��m�ӑ���1z:J��:�h���h��.F���<"ѵSWQy[�L�}�W����o/��O�7.�Mwqo3x���{�a{'����䶞/Y�w'gf>i�!Cڏu�|�ꖜ=��f��lc��3y����p��m��i�Q_e���^�����|�N���OT��~�&�U��7�$2���۶��-�KT�N����.�%��`���e�6�F���A�9�>���5<d6�HJ|z��#Z\4�9�#=+F�=�g��sf`�lƽ(|�ޢT���6����qQ�0��\�49�ڃ��M���s��j�f����6�lvx�f���:"q���yWXH�~4 �;��/4C���zfv�|��=���%���+���8^p���j�8D�幍�4A�v������<�8����������k���:>}F~�W�wN�\y��O�vk������e���ff������YӇ��w.�={��Pϖ����wG��Ό��'^��=e���DKL�8�[Z��*U�dl��~�?���)ϝrX&;�̰=U���;�4����*:`���Ip6Y�������@>`|˅�O�a�dU�vn�&�1���%�H�O�D蛞Q59���A��Oy��0W��2�0�s~1�}̦ ��K�ۓ<������8l��I3��~t���g�7��=�z��ɟ�3А�.��9�Kdi�փ�k#�t��ލ�f����&�i�W7��[�O�N%i���� �����1��D�)d�z@���D����1��?l�;փz<�}��e+��w�l��JV�</CVx���m�Pk�c���?*�k�Ό���7Í�Κ%l�9�>2�UΆ�۠�r5����{)�;����y����s̥��]�s�<Wh�&��-[�{w�f�{��.�jݮ6ۡ�Y�Ye��d�fac2Y��O�m���M���G����m�F#��5.K��#':c�>�3`sT���y��!��Ą�R]i���.Z.U9��eM�ľn=���/���o����x�k��Ҵ#vb_f��f��v�Tb�2�`���#����B1�<�\.�j��o�B�<��&�<�|����;�:�f�]��[�^�|�b������=9dY�\�z�t����ޫ̹ã%k ���F0A\�C���̌�{{��W՚{5ػ���5y���#��Q��[�^}�;��C�n
�ȍh�gi�T�Nr��@�u���n�]�n�����a��1�`c4�UU�s��j�x�i)Һ*�޻�Ʃ��n����L�zg1�n��~��ѼL+����T���P��ۙ|h�*c5��g�j�����g��+���E�L����¼�K�����L�Sz��Z�H�Ο7:kO-�j��եV���Q�K�g�#����;<_qW�����g!g0�Ų4���`���qD� �8Ϊ3�c�9L��Ό�(����Y\�r�m%VK|�iġg������'����w��0��)�6���ݘ_q}Vαȳ�eb�C3\n��;ӝ�|]�s�{�s<�f]\����·N��:w���=���ww�Ϧ�Zl���}Z���<u*�_)�L燁�����Gq:h�23��qP���u�=#^Xȳx��'�x��}��z��[���WBYL��LMԨ�=W/�e�&�Fi�����H�n�x�|����Y�����Q��ڇ���#4f���2/,�;Ժ{2-oi�i��S����r�-�L8����y�QLm�'�·I�׵��>̳�̞��!�=� \��Y�B]�5�drioD�����좑�cl��!��f��I�BS+n�>��ST� ��ʖ��N�!�Ԗf��ةz=����QTzyj\C��l��.7v��/�F=�T*����*�b��ӦCl��.^)Z���m&�U=��wbNufa�Z1�Q�^��X&�
<O� ���I�ڷ�����{�1�y�g�~������J��.W�7o{x]�a���R�9F�=���9���ҟ;�PPn>ڐ�l&����+�a��+.�,dqhz�Vw
�Der�zʹͮoB�=H�n�:uN�J�~�����Գ�%%�Y�2d���s~����QI#ro�����f|!�-��Ɲڵ;�P�.��RɽǓsj�0M���	����?�<�����y��7;�%�Z-�]:��pγ3^���U3�ўe�l�\{��;�j%�^5���4?V��*ѭLt�U��=A(���d7�g��;�ï��ŵ	*y{���]�g�W�	+ǔV#��Ɍ>g�q���%�S�� m:��*�X,~��r`u�g��x�V����n��C� d��躼�7-qJM�;-�=��X��~�O@Z����p)���8��!�G�<�*�<]j�[	Tt���ѡO��V� ؉o �%�9g��ۛ�wR��05F���/����V��=G}�F��0�S=d�z��Je�N!ӗ��fq,��v��@����C���}!\<�1�nЈ�>���t>[�aJ�ϕ����{��E7�R��[��r;z�QpҘo}�����!���OS����H���Z�}f�%8^M�^R�si��Yy	�6��wN:��j�U�ó�m�����m �����^^g�������t�ݺv�buzϾ�{���w������x�{�{|{k��4Öb4�;�x����G������L-�M�]X���v@���=^����*$���pV�,��[޶�w�EZMݝ����X
���^�1�XS�܊��/1���}�#5�I2{��{H��B�����[U,m!!:�t�aI����{a��Tog���/)�6v'���-O�+��W�'f��-S���9P�f��9f��@���ռ�-�9{������<]y�_8�nnfZ4��=��g�r��^l��}~W��e��E<4�윬<H��J��S�޻m��#�^p7"3gq�7x��T�&��k�<]��g�fg�7��8�^�.x��Orcґ;h���(KDma�7�	U�uF�;�y�*Tz��H9����"9-�]���é�+nNN�۫ɶ!u�miT�8����9%�9]|���$�"������4���*��ӇR]ܾ�Y�Yi��6Y�����c��f�C����s�j����C*� �J�D�͆�o����j5S����t��&��%wNYط;'��a%5�f��88�'onΦ���l�Td�d\`���ܧz:ʾ�+-A#X<<��	�,��W��-''L��Y��Y��lܭT�b�|ys����>�ʺ�N�d�i�ۍ�8�ye��gO!�4e'��N-�-���9�]%���۶�o!�U��2n^����=}���#��:�#���8�|�l�/�%����s�Y��FS��NwvD9u$.�^7%��nXԈg���AÔ���`x�DH�=��=�C��#�M�.�3�`�#8Φ�.�'=�@V1��223{_+��%��������*��s�̺�aC]�0�`��]4K�F�ې�	�K�ǹ6U���\�z��x+N���Q�Ӝ�sk�]��A����}z�_�8���k�����	N3�̜�q����Ѷ��5|@�9V�+��]J�슱�V���
|в�D�R��9�{@�!+�R_+�AS%ΌsTPЫO];��W��d��f�˸��ȑY|4��.���E�A�	(�W[�0dqV�?Z!3^�Dt�3�Ւ@�Sa*��u5�<fYv�-\b�bQۣ2�>֔�y��,-V�`�SC"i�tRW��Z�)gu@rq,��Z�-f�i�T��E��D�����]歛O;�;�JUPݺ\�������gtj�����x� ���Ǫ����6s�žy��-��dY��yr��6�xV$�0�[�Ut�r�ڼ�սj[�۲U��S�;M�o�9c�혯0����a�Z��uo)�����T�$]�T#�l)hf�fI��]��s �$/`8n]'O�� <�r���o.$��<���<5��cTy�>T:�Xo�U��}�\���]�e&c�GOs�E�z���c��K9v$]ӳT����9[�üQ��<�QC˕��������6:j��:U8uJdeu=aW��֛�2d���ir�m̶PCmtӜV�c��p�R�mW� ���XQ�,$1=ٷ�-��|���e�E#bh�ԻUG����u�����U��A��e�9�tFP���(����+���	��f����L��-;���39��;�t�;��=հk��`새���6�x�9c��;clUXz¸�V"�C�̬[[�Ub"�t������;v�m|xֺkZֵ�mk]��k\q���]<�95!��Y�"|�(�[��UF�������j���6n1�i���5�x���kZֽ��vֵ�q�q���|��/�dľ9�kE�Ɩ�����b�)���Y�Q���beyLa=ӨCZMBI=c����xֺkZֵ�mk]��k\q�}}cÃ;J��Va�J�5�Ŋ,DD���$t�T�+Z[Y�;q�������kZֵ�k���k�8㏯�xr�ZP��*EQ9i�E���,6�WZ��*ڡ[:�)F*0����*6��X�QUz$����+N��}i���D\�*��6�,Q@Z�AR�J���Q�.#ˈcU~�*
=Y��d�(�|J�Q��T�c(�-"*�P\hv��nHWv��!z���Aj*�i(ʕ��"�۟P��y���Y)��Q�
���1Ȃ�Mی5
��� ��ըF(�@�.7�`� R@�i��������&Cr�d��CQ��`�����b@�H��[�1��M����w3r���chH"�D�IAj#&@����H0�$�.Tg�OUB�/��n`Y�6m�����zH0{e�e;���S��}�]�*�Ï;����h�a���L��m�n��1k]]GM�˺��.�ũ�Ms[�����GJf���R�7���k+���D�a)�m�:J���%0D)H3 �)(�eE�r�D�"1��M�R?8%�̄�c.��Ti(Y�D�E�[���"�a0���l6�-�L�Ɇ9E������3v\5�T�GtM��8�a1!R&�m�(I@�s?�~�Oe�3&JK,��%�&�ϟ�0�����\������D��	��k���[rrYW�&kY�P��ڵ�|��yn��S��6��gsԫH�����4W�I��ω�}ц<�\�\�ױ�f��Ȩ6ͯ��+�u�(��:W�[�$%�h�#���8�� !��MMCq��mmu��y#;�ݚ�҄�~R.T���kL�S��ko5���=d�$�Gtq���4�$Fi��2�>�b���uϵ�{��cg��4D����^�cl�;J֧�@$j���J�]��#[_��>c0<}љ��*c��+U�sR\���wx.ݚ�&b�q>o\�/y����#ss��7˞߻ӤH��U;���Ү�,�K�x^��<��n���_����F���_#�7��h0���G��{�u�Gi�/�ս����i�^�!�g��))�x��+�rqz�En�@7 ��������|o� �(��C��i5d`(t$���M�+L�3�̮�oO)LF
v]b�ybf9�.F���UI�\��E+��5��u��9�M�&]���3!�ky�(a��vw�a��ӭ�>v���'#���c�S-ɀǿOe��%�3&K0fL�ds��>��v�������qj��h���T�������ksx�nٸ�G)}��}� l��O���ʣN����vs��a}:��WwO�8f�w����{c�P���?���ffz@���r���`�L�EhƗ��Glv�#����ku��p��� g�M�hT�s��B�j	+Y�H�-����h2,X����9C�V���m
y��d�����G8�<ݞ�}��8��	ʝ�z���R���3=�l�;��+�϶ؔ����D���'���m'����,.��Pv���s!�w6�q�k��\�G
��fe��y�=�&=�V�!Z��[Nv���w,���������i߅����)���{�)���1�/\���F�Q̊Ή[E+ӹ㖅r7n�%��Q�t�\�l�����r�ط��(�u.���F��˱���j店gV�^�ș�r���*�lRZm�;�gN鲙"S�4E{���U��<�N�wVc�oIԸP�Y;�Br+3�*K��"�.�
���l�::���Y޷�u5�o��k];�ۧq۷N�����xz�_{���e�������	cy,�l��� ۸�ϭ̊�x����w+�9�.⦞�-Z:*��\�; e�+�-�%������󅾷�3s�*V��,,���w?� Ǥ���4����%� ύ�Bhn�y�Mu�u��^��!����|��ƽ]������uy-[ϸ�"��{�eٔn��6K��W���h�m��v����G?�x���W7��"��-��+ko��Ժ6@gl��f�9���Sa<A�r�j3�m[�ܵ�j���ff��G��_�K��./�������Lv�f�Jt}��p57	��@F�C�kJ>������i�S��˼L���ۡ���Gg��yb���wZ������AR����؇�R�w	�;��g��f��o�qRbс���� �k??4Np���[�
Da�p��پ	���9�d�=.���QLy��?ed�ί,bY&�A������F�����.f�ZC����,ÖvBmD�),Z�U���&�Q�-2y���噶;�5��k�lv���ӧi�t�C��;��=���?&Y�0v���}�+z��+�a���ys��#�[���yn/��{N�{�����:4*e��O�i�Kӯm��i���/W"���q-""\c��i��W�S�kH�W���{���X��Q�i`�8̠x ����{�>����O��?/Yu8��z�\��n8+�j�wu�0���<O��Q�����@�@�v�U=��_vꁖ�����(,�������=��������M�$�7s�{9�0���U��!Dc3<;�4>�@�ff�1�i�7�5>u��������q�3<uEMj�-���t��c�S�[�{�1��W�z�V�ޭU���ܙ��g_�]�^�Sn@�O�vzA�3���\q >�`���,��v�F£��N��^ӹ5ǥ-�[�L���c��8a��Z՘���|�r%�U���5�MA�O��#������QG�+30���r檸Ff���w`{(!��O����^�ŷ+����.���+��=ز�rT��%�1��2�+�7C1J嬛����>{�o�j�d�$Y%�{������<fL�dfL�dfL�d�����_Ï\�:����-�r�_殹S�͛�[5G��uR~8
�u�[}P@fn�Q�]��G�u�cNsD�=#�
i%7"S2��6{�ޘ������黍/�IV_��/0� ���>�"#jU��X�IH��T`�v��̙9�r���\	�s&.^��3�����8�{��7�/z����hF�)�FK��;�kJ�;�x��&Gc��5��ff�z���Fy�� �y�j%�#�090!�<�.��l�"�����x��s��~��^wp�ex��*�w�+3�P3�t����,;sX?����#�|��}�Ѭ�@�����;<�{[�U�F��a6�b�T���P1��A�9�s<��7+x>g���l�T�s���R7s�I��D��h���m�j�:�����=�c������Q�}�':�{����<���(��9)N��ĺ��w�P���.ßsO0�w�]� :�J~� ���=�g�r��]��e�8��	�����\%�ߗ�e��&�P���{�}��{8t9}�S_C�!CӘH�>��'f,ʇ���Z����&�m�6��ԑ6v�����q=�s�h��5����jw>I{����;c�n��n�;`mۧi":���>����}����3tm|e�7r.���{"=����|#(�κ�-�5�I9�&^q�$��֊J��g`C���@��ƆX���۝3���;SB�j�ܽ�; ^vB͠�zV�{S�����#;< w�4�q���� L}�h綕OR>֝��)@ݣ<�#��/�U��*��]��Gan-��-�dA� 
�$���]�/!JK��ze<�����U첎j]L%������ϊ�vnd���1«l��(im����8���QY�/��(3��uO
`�ѯg�Y��l�K�gTj�l>��(�z̃�k�`�3�8�{������6s's��%��1�AՁ�6f���[�C�����qC��Ⱦ�d�F�9�g��wj;���i^h��Y��������wb�Y#�"���K3n�j7��X�δ���L�bl�ٙ�Prwz'A��F��9�,����:�n��dHZ��B�1��w�8-�K{fs�;ow6u�ߛ|�/�����K,�Ye%�Y���{�-�4�;�<4;����������B��w�$U�+zi�T��uE�i��[�p�m|�`hj�RW`�
��H4��S7��b[29��;`�J����3_�d.�ck�RR)��E��kw�E��{��D�p�[$��^��q긻;)�ٓOd�S�g��d;n�ڣ��wz,�x6Lșww��ft6����q�9��ca�V&�>����p�����9J��N@��=�I.�6n_�p۔晞�'i��|��ht,؜�
Y����H9���w=��Q�Jl���qd{����JG��?�=��t�"'�e.���|�ʭ���'Z�%��uU;���djN��$�U��3Ľ⾘̟9ᙢ��3܅��[�]>�]�+<�\��3N N�>ViXs٥W	������Հ?f�w8}���}F�wW�˳��Sݹ�enD��3�R8W;�f_D����w!��f�h��f��� I�I� ?�MC��b뵦W]�p���+����i�':��.��@_u����^�0�5�mc�V��U�1�A�=�:t:t��۷N���o�g����g�I�;���n�l��ݳ��	��ÏpUm��p*<J�;1�Dg�������zd����0��{~O>� 6�S�q�}�y��i�������+��o�k6G`\�'=~Rh9���6y�^�drČ�M{�'�y㫫Џuh�o{�m͊�y����m�C(��E���)U�w
�^H�g���R�sU� @zF �����U���~Ԗ�Є��x�2�}c_��z�����X&���[.�G�fu�5ԑ��2"^Y�Df�,�sz�=����=�C���n{�z"�����s��Sמ"��v����qOY�k�Q2�L��`���v�3�ΗNt
�Ѵ/��F9����ѭa��� �Z;G�[A�-�c�B��*�{'��XwOwu2�kY�m��C[?26�'��N�x=@��3<M2�Ή�i&��4�-^<pI�G
��G�E�.C{��9j��8���\s"9V�rظYi!}]��[ qk�}gZ���t��+����r*Õ\ ���d���%�̙),��P�p�|�k�,�TB�����
�p�r3��r�w�Ӻ�E�-��DK�u�yimw�B���[��:���EY;R氛�m�­:���&
�j��x�{w������u@|{�(�r�ծ)�0𦷸S[�M_�-Zz<�����<���\�vK��Jr��z����[W��Lwp�س�N�c�;����m��Wx<��ôC5I�m�_��Q�o:r��	��8�K�����-瀝�e��o�9��s_�w����n���;��q�-G7��E�(n��%O���=�i�Qq�o i�;���0wÞ�y�^_,���z�� N�7�*7�����Ţn�]{�0�^q�baٓ�1ݒ\Ĵ1nޮ����/;�l��H�!�z|�'��=��!��`˞X��9x�c�Q��!�f^&&}:�B��Xi�>{��W�^�暥�e����kL,�Ow�j�ͻ��^)�n��\M0cX�6Avʜ��L���~�n�x.2��Ζ����'C~:;1�QѶ�7���U�&�˭���$fm��B�C#z���vh��U4�����z�,7�Y�bF����s��e�6�]֚��j7�5��/V�����??_]�n��n�0�G����0l�G�gq�T��j{v�/��&)		��H�O�.}%>T��e�<tj�a꧟:`��m�){VSܕ��-Y���;�?M�����|ܐ�B��}����~>�^��񕞾ܱ�����쥸��/� I`���w�V�����歳���}�t{P�T���7�=���˹���/.���kb�u9YT�}>�,���T�E�+� s��vm �dNXΣ�c�rv�P�O�3�<D�z��Kh9����/��]y�:��f�{U�g�{�����+�����[����Ȝqy�p����ol�fXcy�U�	��۫��j�%h����˻)�=26S33sϒݓ����r�A�yz�zm��Eڳ������ꭊ��;@qoL�����Ƹ�8�׏ٹ�z�;�^�g���@S�s�]�j����驆�����_�c���7.������=U�^�˷v�f�w�$�S)n���{g�B�	���Nq�k)Ud���&2M�kmJB�r�>��ECG'�%FQ�%��ܓ�W;�\6��4�8���D7���:+jၒ�d+#6^M��Z�����z1e�kq�QK�p�B�B.u��P[�K6��V_C�ͪ�:㢇b,řMby"=�̨ٖ
��-R�+r�R�F�X:���g��b�|%�P{T���v7hݝ�<'.ص��p������L]��ܡT��u�c9X,<(���P�[C�ɖ$��Kܰ�x9໼jlW_0�;��	�)����n%�Q����ͩc5AHD&�zo�I�{94��n�X��Y�pX�KV�oz�8�h���Ln`L��	����e���P*��]�Ont�y1�Í1��fel��cL�j������a�u�ڔ.�'!����U�Yp���d��.��Eh��2�D�kŹ���#��pm}��ev�K�(9;z�<n��	3:�j���A\���vZ�;$�ѝ�u��0���vl�/�����y#hp�T��̵:��h��p�'��J�PG�Or*���+�!:,��*�Ȣ:��y	s�2FsLe<�O/;������X�Z*���:Y��8q3^�:C��d �!RE�*f�y�NL3n�ɉ8���-���2���4��J���(5u�ݭ���}�R<�\{���Ѷk�9�[tѫ������Ԧ����z{��x�j�7B�r�O/;z�9iC(UlxԸ�l�_�Z��v%Wo��xd��ʞԻ����,Qtq^Q}(�����pu7��6u^TQ�����%�U�mZ�d�:�Cj�Z��I��=F4�蛭�`07���S��r�}Smn0��m�]���c��k�sx�ÒK�����iA�p��8�D%.m_3LŮ�(v�.�{7�;Y�R�c`
dC,2Z���H�;yj4�`��e��uÖ��a�ܭ�mk��f��y��N��Ȼ��F���4��ک_�ͨ����d+t� �;��ʳ��W]�{'\�5�[��'���Ÿ&�6�
��S���⽫Eh�����s0�)�v����$w�4->�s�N)�K2|���`��1_}*�ܪ����z�����?/���ށJ�����ޔ�ktQ��]����۽ݽ��ܻ����JsK�$tr>kv��Lm*��ʯ��!���  ��EXr�mB"�֞�"�(H���n��������5�kZּk]5�k\q�}}cÓ��2"2
,��UH�QD����_��S�Y/%�d�}>�5�kZֵ�xֺkZָ�͞ω�w݁�ň��?Y��+X*/V���V"��٩75��Dd]Clv�|x���Ƶ�kZ׍k���k�8�}�YR/�fAD}ZX���`娢������È"�?D�Ĉ�����#�2̞N�S����Zֵ�kƵ�Zֵ�qƿ���Ŋ�
���V,F�m��P�DU��
��2�+P)״����>B�T���*���w��
z�DY��ŋ&2<��B�T��Q^4\ch+N��2�.�I��
��F�fQ�.Ҁ��TE���N$vʣ%J�繂���e�G,�X�ؤPY*Q�I�J��d��B�2�(���X�S�]LE�R����h�H��~�ޛ��ݼ�ρ�-�Ưzs�l���&��M���l�N��gh[ye�rr
.���~�{n�N�?�v��v�ӳ���'?<��󗾴iý������FQ��0y :��~�5D�V��0ĻW_����y���}��m���Vמow`Y�2��^xC�U��3���z���|8z ;��]�sr����&��<s�>������;��ⷪ/�E�z��ǫ� 1W��W�nr����D�5�ʓ�T�f�`�=��}m��30i�W�g=��ċ�,�]�OVO.�DɤXJ��L�"hoB	ګ�����c�h.6ilM�oz#2�_-�&q^_O�=n�N�
�d-Ŏ�}�U�Iſ�E�3�Ѩ���KsM�2-.���T��ji��a�T�6ڛ���??nmNn�Hհ��Huj�gg��O�Vz�(����i�鞲^�u>�L�o>�^P��"{��k�2uH�����P�VS�;^w�lI|���g�Vf��I����ڋ�d�L���38f�B�����ؖUY#G���<��6���nmf�<�������pl�gG?LٸЯ�{fUk��s�v)u��a�x�L��v�e�wW��4uVg5��������^^^� G���0j��o���v|�b� �G���sO�3���K�l���jRV�z��\��+�D�Ξ�5���ma=�~-���W�G��t���e�7R��Ve�+�I��/u�_���[�.NȬ�H*�)O����woR��s48�ݕ|�2}v7Y�W���l[*�%؛'�ü�)��P {X ��y0�������*+6z�y���LmV=�,���1���M׺����ӭ��;35�_�ӿaʽ����r�$@��}��`����R���뽷�+'mV�(K#Q���kV�qUr�*�.���wI1��~f�[I�w��9��LMN��Ī>�#�'`\�����!f���=^��T,ּ�����{Ye���cE`�7O�o��qk 	O��
����F�����!w��ڈ��Ua���5��	��c���U)�u���[�s��ݵ�;�_P�r���
T��]���l�鸟rJ�-D��$��'�q���:gq���/�>�ݩ��X�ҿ��K?��2Y��2Y�ɒ�$X_[2�P���B�^_�vᴃXgI:ggtν���>�B��/&T�;��Y/UF@�y"1���_OmC�W\/�z6�3C�:(b��ʉ�)}� �(�gl�w����OÉ���É��u�n)��
`��g�n*%́���L���ɛ��∉�q���b��F�0�?M��w�۴b۪O,Ѕ��|�8�<_���.�3�t�V�W��/r]զ��xxwUb��2��y`���r|�zs�������quW�ߛ��'��(�u�乎���(������v����!���r�~,���CtwhYH��f��$��vJ͠ܯ[���\	�k�p�.=#��6�"�+�=y� �i�D	�ٮ])n��p 'g�k�z<zE�[�}ƍ��N����&��L���lV����T(=m,�F9`�X�عfܠj�>C7�Ӕ�'�(vוMǔ���������8҃Qg#�������򻕉5-S8A���G�?*Ş���Nl�M����Sq��g�a���Ǽ^ �ݪ/>��!�����}��{Ӵ��#�F�^qZ{G�0�}��-fc�}�Ȭ޷@������^~>~~^g����ޏG����k3�v.�oNw�kc}���a��s8뒯m�{��t\1���sj"�v��Ѵ��Ǳ�`l7��`��}��w��0w�{�����m�cN���my����fA��->�	�����5���u*�!�V"�L�7Q^�L����NV]>n��0+1��������P��3M�T��;^οF�!�c����gS�8�S.��{�n�;-�{݃���~9[�Q�`+p#Jݜ�jh�����߯?<ίy�q�!-тRT�;�Z���'���G�>z׈��$��1~�o6��/�����f�L�+��[%�����%�3N�i���w"R<��T�A�c�mzߛ�7t-�C�\�8u��b��I�����i�`�<�v|rA��}I$zM��s�8+��|�r�YL���*��o;�T��O�N[�ػd�����ft�(���,�xlPP�F������K���_�u�fʓE�prC�)�h�^�<2���6L��0e���~^SY9��w�S�?_��t:t�:u���y��f�t��{X��S�����:�;v�a�����g�� �Ha�<5�ɘ�'+��d�S0n^n��K.�*�|���%�'y�y��7*���۹{�yV�����̜0\>�-�� ��d��Jaɮv�!I��͕����:�������c1�N���\����/�!����{#ygJ��UB�*s}���F}�皺\u�P�����7�,Ԭ�@�}��ں��F�5^��9���2��{U�C�\z���ʹ�jΨ�aT)���z��o^���Qs~v:��s�b��z�s��R�����iJv�ӵ��Q�h��:A�S� �X�S0M��+�f�%v1T���M�˳�?�+�p�i�Vx0nܸ��o���y5}$8ׅQ�bbZ�V��0�>;P�o���yP�0%��<C��z�+SV��O�C���.��9.}�6M���hK#�p[�ɩ���kk�x(@-��J���Dvǣd����\��b��\x(�U��t䫮��8�.�����Ɋ#��sU�<�}kv�z��ys2�D����;v�t�q����eR���Kz����d��y{7Y��*�gClO���uP�-Z//|)���o4����e���z�-��TӪ�5싫�zl�m�����8������z���ECiń��)�O��4*��ӽTk�9����ss��w�G�G�4L{s�L^��ކ�bIs<�;5���}�"�5��B�����u�C��oe=�Y^:i�{���ٜ��� N�N_BZv��P��ll<���SÝ�\������<��(1��"$��y�Q����rU� �T@����w�_�g�7~]���k00��9;y�\�F�����ն��j�)KvY_HO�x�-��`0��^��Ǽ���{2K�'Iuj������)S���J��f���z)tD��quՙ��_�݃Y���ȥ)��#�	��]q�#r`�	^���S�U���!w�tz�Ǩ@�}��j£G����E)�1�&\s��/Oܿs���F&�Pg֕*yՆ8�X��o�������jw����*�q�Z��⬞�����I�oZ�{E��]:������?��e%�Y�fL�c2d�?��3����%z�&O�2+�Iȅ���;��5����lI�۬��M��&���u-޵7;����͕bV>2��(�R�E�(/;�T�L32p������o
���dqYq\�����{|��|ut���g%�	���٨��2��u�A�
Ӯ�x�hxPH�n*T�-؍Fm�c���9dh`��(�}��k�%�pw�[��<���\�S��κw������R��¶�\�߆W���`�=��e��a=0�dN���ܹ^ڵ�N �ҽf��e,������Ѳ��;{8�+/A:0iA��,3y�+x���	ZO�N���K�5��N�7���h?s�n���V>_��O�@PT�7f4#�qKL齛�]m牦t5�̠Sg�\�0fNk���5(|�f���S/�Ul�ƺ��v����z��u/sCMI�X)��Xx�p�V�v�����W��ߩRU̘=�X��~
��{\��t���ﵯ�t�q�؋H�LB�K�h<W�oI9N��9f�q�m�.���zܹ*����@Qς"��zT�v3�U꺫�~iMԵs�o%q��jY޽�M�[��z7�i �=�K��s���y�|�ۡӧO�v��t��A���{�|����7���Ku���Ƿ}�=]^@�kt,W>��D�y���s3��s6��I��Cun���F��v�G�6��M�m:S����vl0�d:�u��n�ת�w@��T�k32��s����օ�9��ٸү���='�p<v3���boX��G6�%��A;���g�*N�k�mto���Οq�*wc�W�1=9�yP���K]�h�]�gww8������`,f��g���Ի��+k]���V�Y��fD�Mzbj�����\��\���}&�7��{Ч���[������g,����Ґ��E��gA�Q�ufVO�V�[~�ߺF���;ض4y��qx��*�wnNs�JJ�U{��8�Q��em��;��۴oc�.ރ�ot��q���'��t��9���C�� iE��n���J4,Y$X*�=�u�nU�~ ����[�؁/y� @щ���m:.�oWk���M�v��]��=��&�[��+�!%L�ߝ��{���s\��w~v�ӧO�w��?���f/�{�vwl�z��QT?�/8�7��۩"kك���>�۴����c���泊&ٙ��õ�\�
��4������*�,��Fp��e�ե�c��P|��n������y���Fg�$��6�oO@�W(D��ɾޝ%�*���۶>kwY�k���׶�o�LD;8�(=�>����A�~�k܀Qڍ}n���z�&z�6ޔ���c���c�Ur���)^�k=��ꜦG*ޣN�KN����`� �C�j���uB5��#{9l�~s���oJ�ҏ��4�ͯ0m`9�����\�)j�3�s����ٝ�����3'��o�2w<���H. gy��VE�Vh��<�g��7�"ϖ�b���(����t�Aky�P��Ov;��O%�#�̍<����r=|�*����	��C��e�c���֝�:I,l�ȣIH+�b�K��iP�S[����yrR���,�;0*Ӭ~�ǳ��6V��>O��]�e��q	�3\~#���v���ӧdv�Ӱ��}t�:��0z6㕊�5��r2 |�N��n��5*m���1W\��E�.��,,gS���-��Sٚ�ZC�A���]ټ��TƼ@g��a��l��8R���^-35&���}�'۾�B�;E��s�R��;�1>���E�@ܧ��=ՌÜ���9\8
&|��n/oggsv�Vc��:��ݣ7�ot35�ږ~C��󘎒�#;��STVE�������!�tf��G*���^�]��|E�(|{���Y����(> ;yy��t��T�Qu*��+"�}oz���jN�0-���L]M0U�Ӄi�wWuz㮫DJ0�}~����->^΍��[�qsݝ:��I���©z<�;w��q�OtrZ�pGF�I*t��1e��2�������������`��n�8���E�t����U���b���Kv�N�}�����VW ���Qti�y3f�`B�%��.��ղ��n�7*!6��쾍m���n�s��[;
�f�:p�D��#���狷���n��S	t�7�Atb�;n���'U8�vXV����3��v���݂c�*fȺ^뷳n
�6�����W|;VW4�9��s��QGv��v�vY�+*��Ɣ%]'�m��N�k���iS�u�+ś��qV��ٸ9)1\�B��% Uښ�ý,�#L�룦��x��+�ۮ�V�'��6�v�v�1���&�q�f��CO �ܮ�}n���5�
�Vl0Z�Iu�Q�%L�/#�ºP
���Զ������.[��<J��+��*Ilۺם�sm���ɯ\�e��:��w!�Z#��JYĉn�:��\)ps���=k/6���]w��ަ���s�[�`cMwAѼ�;��]��*��!��>K�x{|r̯��v�I�Ip�Xd���vٝ�k8%|Z���mAq����P�Л.�D�X�}j�n=}ӝD�v\,X��N��W��Q"�$aq?�LL_!VvΥ6h�*�d����u=7(lgK��%B;ݨNDp��ڪIoKb,�A�豯�yH��N����+i��m[��K����e�VД��I�3v����P/(�:Wk9�0��|���G��"Jl�!0��B�	��8����L��X�9�U���U�P�ⷽ��{1.��^P���4h���HR9P�ǩ��{f��9K�����j�ȝ�16)ZC��-=t��Y�;��O�9��ҤI�ޱ*��%�z�Tga�1u#�tm�OB�Wfl�j�~௲�ipٴ��3s3���o)L�����ޗ�D1p[׵s{Jx�J��WA�]�ٷO������X�V�,�G����qv�΄��i��ܪ>p�F�L��&�VZx�/����=�y��ef��\<��A�R�a���T���8s;�e@Ax�Jx%(���w5mC���D�f�3�]�A+]����ݙS�����çµK��x����{Q�sH�*"͙6�dܷ�D�Z.���������ot��=�т��Z��G-�E��^���gGqv�B������J;������־�&����Q>��U��g.��fY���9�o
�w_'�$��w^٦zf
O:��>}'wN�ۘ�NWZ��n�5
��@�,
ɱ���)�/�LH|O�u��T:J����5��t�U#��YB�C���Ӎ}kZѭkZֵ�Z�kZ�8�_��^u�Bd@�5�RE�|�k<��{���Ð�H�1��ǧ����ֵ�kZ��5�k\q�k���4j0g�{B��S�,1�U�+�y`��`�h� ęg'���_ZѭkZֵ��cZֵ�rl�|N��Y�Kh�wK D��`�`�X���xeI�&M�B�;t�mkZ�ѭkZֵ��cZֵ�qƾ�{�$��Ґ]��*�J�EATP�)�+���Tͦ1`��H��U�A���I�f�|nZ�@Q`�[�5����bLB[AT���Dd*�#���V*��*��YX� ��E��Z�C��
x���b�m�У
�d��2�%�̡�E�mU���IDia����E��$�QV�@X6R���3�"�.XV,A��Ӽ)3RB$�:L�A�Ad�����R�X�M�b;s6���iM�wUXcqe�Ĩ��b��D1(�1��d���(�C�x�Q'f0�v9W�םx:���Ŷ�gK9�k9⌎v�)��#ٙ4����̭{��vN��6|��"&�D�#I�ϛm2���N|S#�U�����i�TQ�
b6�%�R"�$3��",�	�B�F�.�mIC�7w0���6�w*`U&T�ݍ�w-]�u2�]ԴV�R�7�ȣa���0��Dy3	��l!(�%J�D �iۢ��PP33n覫n�n��n�nfc.�c7c1�¸i�u6RYe%�RYe���#�mο�n����11nʟ�X�;j��;��ڛ�k���'
�j֤d��\�X3�*�	�9dt`�4Q@��K���)o-��UY����~�_l��셑��m��#�;j�c��K���-���S����t�̼��5��-^�c�f�6�k���sY\��e=F���|=����4�J��T�������x�X�A��٠d�n�9��~����܁w<�v��N(���Fnb8u�4�=���n�b�#��UU�$�(b}<'��t>0:�ǫ�O���Lw]�8���Ȗl�1՚Uiw9���^��;�?���r�u%ﯶ"J����o�řlud�\�����������mz���;9�Hi����v�pl��eA͟6^�۷�O�7;���z"�M�[2����Q�M_���O��� ��*/ie{-&�B:�+kM�89	��aw]���*�1g����vNx�W� �ᩔ3��Ҋ�K�+���>�z ��J���e�~Yު�L�-�]�������&�X[g�)��'�)�X�A�nwv�W��*��h��U�u�x�a�(�s��*�w�v�Z=�U���O�������G���y���wy%\}x�s��y�B�d��n��}7�3FZ��Kf���層���N^�)Ӧr�h��&���@C�s�Lr��Af?�~"l�B������ުl���T������F��M�}��"�@P35e����̥��a�,�n������l���������5�]Ӄ78�S�gIށ�^�I����eг�����5lo�7K�d����}�Fϫ���}�����9���!�gU�]�wb�����1v�n���&��Guw���l� ��s�8�s�@�妓{2�4�f�:Ξ�Wf�����p�g$e{�@*;C⁗�.xV:�E��8@�=�Syӛ/���4�!�۽&W���R�%�*��޲b�1����x�fB�c7��h�p�����2e`�`�UpnX��u|���G��2Ϯ�s�J��mJ�K$��w�ו�8�T�y��Y�)������>U�;/�Z�&�e,�ΎЙ�G7R��z&�5�I�����뜷���񑌬��B�X0a��~�o�{����A����fy�JC~��O�����~8��.Y��]v���Z���G���=ꊦ`��n�,�m��#x#H�A[��K2�6Z���F����<TUS�^E�����MԹ�:Z2��۝RkO;� �窓B8��Gu@����x��6�+7��K��o����r4�TK�7��?�LǦ=�3d����:�Y�"�2׋W�OL�Z56f�$
g��=6�}��0��0紥IT������^�P:����*��@>�N���ݝω��%�sk�y���Lat/tV!3�2Σ���$�����uD4��3ӳ�;[�Ӷl����ζ<�.����tz�WnP����3&�1߂�N�ջ3R�C��w�Tsy�<J�<b�����y�c��*����M�6�fn��Q��ꋗ'5z���;=t���z��B�I#�"��X�a�͘hu�\@`�kZ�F�p)�x)w:
�8���goua}��N�m��('H���'�]Y��J��no3��K��{�|��0c1�I/�w��/�wx}9Y/.�5��M>�4.�a���_@�\�jwD��eP^�.����w���o3��
Y�/�}~#�������ӆ�!m��;8~�M�ֻ�^;��Ɋ��mnzQ@Ǘ;C�"��Z1�q��4��t�5�u�����*FT��ɞ�Ю֭X���}�\q�5D��EY���ݵ;<��RQ�հ-ς�G6�T�uԵ�H�ԬE��6]5�s��K�l�w��la�J�v0c�B� ��f����,���*��k_�Xv_��O�
2w=��;Z�"m��g`�:K�CWs��_��2�X�Yj��68��(�;�3t-٦ff7M���:n��@�����nf�/ce���(��{ğu�矐���D�������u"��27�~NS�d��N����Y�����x,%:e��(�ڛ���E�*�r���Y
H���;jlO�ku���F�L ��>=u{d`/Vd�e!�%�W�z+�����ޭ�eKطy�I��/1#1�#�3��;7߭����G�s1"��-r�s�tY��d��r,ꠄ鐜�:����:g��J�����Zn�tEEU<�M5���̸��V�YZ�;	�=����t�=4�!��+�rQ����9߹[����>#�,�yh=\�8\��~�
3^�ξ�gn;�W�r����܇I��ޞ�����s��L0ƈ��I�q���kd�A6e��i�Ý��{�چ6������:�K8l�t�0_#���ͻ��y�n�u"߯�Q��X�����-=�Y�3ӆ�v��U�,�;m�#��`�����r���ߺg����}+]��hotfgr�ޫ����[N���<|��7l�,���;���?X ���挎��(Y�P�]��Ii�LKw�gف�s�!�E���\R��Y-q��p�`к�	n��HN��[�Pd[�#�f�Ԟ��Vp�3�o_�w�����lc!����cvvm��1�_oV��sbJ�s�
�,p�ϔ+E1���*����^#�x�im�ݓ�:>�uٺ�x2��u`���{"OҸU��*=�aaS���[�˜�{���O�`�b���ݒ��Ӱf��yY�����s�}��El�cWoc��j���3ˑ��WG�[��?m�q^=2z�̵�E�K��;��'��պq���ų�y����eoz. ���z��pέЉ��K����=��a�Ge�⡘v��/__�M��uN �g۴o)s�I}���4��tr���h�\�0pق��z?����W�c47gmF;#���+:��/��a�r���PA8�S���hMk2e��NV�q�n��q10��%����}��Ton/�W���_�h\�}�i��coҪ���N<3�>RI)pm�>H���ǖ��C�pW5h*�/=�R�u�#������^F�g����CwO�s���WW�k~��k#u��Z����/kï�	�x+5븏L����;�Q�4���KC�!��wv��VΫN���=�S\'P��:�gT�Wun�7�B�)���q__kP����x �xRP1�O���9���|�gP̞����4���u�p��:��$�ģ���ic�0�����Ϲi���+1?#�b��_{����wߺ���Z�`���AU���3�����w��2�n��L�^�v��Z�X�b%���$���Otnz��g�f�Gv�'T�ߗ����Ξݭ���j	D�4�ntə�H�w뭶�ǫ��M�9^���w�Vl���<�3�,�%�w�s�'`� �)��8��4sPҲj�۹��7��"��Q�h�}��p���u�y��1�8�.�nlD;=$:U���ç�/k�����9��,�d0f��0��r�-��W:[��Ly�����}^������^�SS>�r98�}�@ֆ�{�X���o���uF�/p�����?�Ȫ�8)�B�h��~Ť��[Qy/�B��WE��ꇢ`��hK������^��ͼ�X��H�u+Y�/<��*�]!� �5�zj��ᆌS���W�w��\�5讬�;��_�w�>���3�ƑG9�1v����&�M�Sk��ŌJ��W�J���e�;b�)xc��9Y)�GZr<
���Va;#Vsfg@GN皺��?��F`�>���>�y۹��C���7��=�\��/�i���l߃�٬��E����<���d��� 줒��Zc�N��of�n���r�Q�I��'�s�����n����e'�ez{6��V�85��e]�F��v�ڪ��{�l5���X2?��"�@p���*��;�A�(�{��6�:���q����-����PM��l���\ ~���q�������+uY�mm>��a�hEn�N75M�Y�٣�˓�w]g���^�U�*�gp����9\l&}�l۵x�hS؝@8Ww�}}������< T ��� <�m䗍wm�]�����_q$�y������/\����b���`��˻��C��ͫi��k�l�SՕ�z����`<*O}���`�y�xY��:���-��r}�v�r5�P�k3'ʒpޖ���9�kQ,y����CXV�$
��3i<I$�O�,���Y�e���=4w�viU�:��&��4�#�À��I�QU֍�q�>��Υ'f�����<|}���G�eh���T�0�K~u�گ�ۧH�x;gNmWpW)s{N��!��pdr�۝ ��4�b�<��.����n<���rLE��UMC��yj���湊����Ye��=5FzNO쑐�A��[�K��M�Vܧ�j�O�Uo��3f_vch��8s#�I�ݚٲ����5�86Y
v��Y�ɞ�g\�P~��[U�!�������=]�Z���d�ぽwK�r�L5�ݜ3ߝ �>��a�T�z��X����>���jT!����ԗ,�7�U2�/�s9^"�O�=ݹ��[8�r6`�����ɫ̴+Q�so�7��~@K�n\osw�<�Qt��p�����bw���m�K�Nx�ɜ�Z��p�;b�gC-W�|rn؋-A!A0�Et���gu{+�	�M���RP�,��@v�V��|t&�m�:��h
�u�)h���e�����?/��d�J;���[����.�[%���Jy���
��l��d�5B���e4��@�^�|���sC\Ff�KQ�Uθ'����
�qzz��:yp=�05]���/�o&g5�y�$����1c � �:��ϯ��{7����2fO�ɜ�I,7}]6���o��=Th�Q��OG�Rq���q�F���r��q��̩���w�FIO�@�
!�����[ϊ<W���ɟ@�W��seɞ�F���OoX]�xhW����?��h�g�T.��d�Vv�ڋ�QE�0g+�z�^���'|���	;-�`���`P�7XOk�7�	=P|����c���b#6�����789��V�������Jޒ�I7�������T:W�����*�$�fچY<#~y���-�)K?�Þ���B�tV{#��e�Fh�T�EFv�h�y0����X�°���u�[��B��1�a�{z��o���J:V����oW��aY�c��k%��.g��O� �����-�sږ�$��ؑ,2m�" �L6�S���9���S|c})Z�;jl1r��VR��{�3{�yزY�Gm�	E�͕L5Ǝ�6�+���jh,I[�P
r�rt�,,rrոN���G����
{|x]B1f�v�e�B�E�{+��^F9���	C��.���ϑ��Q�Y�g'E�k:NuҪr;/b��$Ό켸z���}MKFs��f���ޛн�es�����F�fbA�n���Fw�3�+��B�\��%2��z�(r��<q���!t�K���g)�h�zZܒ�FIG�#��9�
�Cn�>�Dtb��Y��-��2��b^��Pƨ��i�i[������H'�r�᧯��!���/�%�{���7V��EWBS�3�L�OWv�<���4�M��u��$��Y�C/�;��eI�����7�W�F��:]�2�p���B��0��n���qt�6�`뙁l�.��F#j��*���5��'N�%C�%�Me��}P[1��%�zj�}`K�⩮��uy�f�|��Z�C���P�i�Ɗ��6���)pu��p�\D u�'f����C�WRWLP�Gb8&k��.э�����{�BUR\��m�� �@۳u��*B�˴�C��WT(��-~�VV\��e�V-ô.�U�֧��Hk�����$��u'�0Md$!{�UL��;����dF�P��8ѥ�j�]�F�=7l�)��I3AܐY��;����0:M�"��d�!��֕�������	ǹNGt��3)�HW]X�k�nķ���s5�}��j�G�M�Go�w���,v5�1+D����{�m�Y8��9�����Q�2K��T��=˻�8G����ùI�[��l�l[�r�*����~6��K�����t��5-�̘ad�_ ��W��[j��P<��ѕ1pe�a��de������A����6S�]�s��E�3�:�W-DrX�PK�l��pI���Fv"�![ӈ܋��W]���Xn�$�ڋ(u��CC֙�pPe�M'*
XΖͮ�Jn�6��#[[u�d�O\-:�o1%�f�ٚ��;��d���5��r�)�X��Y��^�.�w�U�&�+��+�M�:�9�3��15hQKZ���0\V�1�(��:�r��������x.L�3*�Ku��x���2K���/�+0�Es\�C�6��ћҍ�Yps�N󱉅Ƕ#c{[�&=uݲ�wts��>�ɭ�#*h�X#�j�|���'�7�]�\%�P�m��wje-J*��R�+"�E������`�H��L���֡D�>;v������֍kZֵ�|kֵ�8�5�� yՁ�bEU��_j��h�R>�PQb��c�AD�޴H2�۷>>5���Zֵ�k_Ƶ�k�8�}x,�#	>�')G�R�8ϰ�%qݪ�m
1�`�&,~���e�z��2rq������ֵ�kZִkZָ�8�ׇ!"rXozM�E!�6����]f
�2����
��#U�㜡U<�~�L�<�ϧ����}=cZֵ�k�F��k�8�}{�{j�bwJ[�0dX?R�j����*�,ğ$�C��|��C!�S��PX,1�%Ax�P����%d>�)U��b2qP3��ěF��;��Vz�ç$���AX�eQ�XVJ�c�ٔW2����'3���@F-�=�55Qq�I�*ȹ��*�KK1�!؆�2رbyj�J�<LN5"���&x�LeH�㊬7p����̻�Si�%��[��!���WsF��:v�F"+��˃ʫ
�>���e�o��&�`~��b���xeoF�u�D����12���&`+��$%�=��n��7O4�	�wvx��5�mEb���dw�#����ha�69,�`ǣ�K�oc/wn��5��s��竀�.����Fٮ�>�W8
ڒ�z���̅xN
{�����;�����C����9��;]P�f������Z�aGbEe��1�jb�S2)�"�@v;o1��(a���nat�S���Ӑ�_lPw�wk��9���-^��� =��
��������J;.L�޺͕Xf�Z3!�WpI�8Y�L���VѲG���}��c MD�g�H�% l���h��aor�>=M�4	��WC��=�7���m���056�������=>�/}��G+̞RXl��͜�nwOHNE��Ke��_����ޗ���G��hs���sQ�Mۑ�6:��\��叆o�o�L�[^S���<�C�^�������pc4�<7y�"g����W�D+=ԼTN��]q���n_=e�����]cc��fJ�Ѐ"�qڔ�����;u�[����y��o0v��� 8�/�կ�{�v���"8Mt���+}5W��ME�IuO�<��;�0p��Y>���x-@�Z�95�,�QR�5���(��㶮�ih��}��o*��O/u{�ԃ��pǞ
y���[���f�Ss�+��o���{ϩ$n�_�&���5`wa�qs�inӃZ�t��MG���;��@����Tަ��M���Z�5�Y�9\�{���weD��4G��G�έe$�ܷc2MM�I*���^ 3��v_���8+�܏>�q��ğu{g��S2���S���'L�Uc�;Ѫ}��S�h�A8����~q�T��Pi�ws��3����^��9�lFqJ[�S�>fx
pj<�h;��@��m\3s�!����O��,�-����I^����4���p�`0�5bX��\��O�Ȱ7�}�B},��R�nq����=�^�yl�̘�A��m�v�Ab �y�1R�L�/θT�DR�(����μ�ރ��*jc.�֫Yg�c�E�5�'�r8��i�9��ۆ�����wԻ���1����W�~�������\	����j+NM�~��#���2�����E����bXj�$"b��u��xS�ARH($Ro՟���㟨X��s%P4��'��3���٠K�l�������c�<���=g�����I+��.�p�y�9ԛޔU�z�*MO�K�l����X��g'����y|�k�o��O{���B0T]��bY�4�Ԟ�h�u-o��n��U���^U�w����3V޻W=��͝~�����Z����ӷt�K�	�.���̩�Y��w+9���=�!�N/�P���=+P�����I�W.r�%��ܔ!�&]oF�R���Uܖ&�p "r�'�ܖ��&�I6x������u/�Q��@�L�.^�7 �=+@��U[m�D˿�?G��T�)	`�����m1�ː�¾�*�lEj��&/ʳ�w7P{��٩f��,�l��%��r�o��v�Ư��G�jw�0�0���a��1��j�Z-3b����:'m\A��T��z��[�mgӫ���؝p���P�Ք���w:S9ikވ�E̶�4��`r�]ˍ��S�>=y�[��G��c��D�^������y���v|J]A��^�:�py�Ǫv��D�Z�8͏91�6��j2�ku�o�oݦ��M��ٖ6���b.﫧7���޽+i�Y���߻=��J�u������d�m�K��f�R�*r�^�)!e� �=����.ښ��Uq������-C�W%@�(�/i�\ǹK��J�:<��Fr�O�����k꫖��;�b�*��ҵ��!q|�7�M�[�iw�,"k�Nt҇�^:oN��3��02�W��-W��s�D�d��y4g.���	λ��^�����}۞ۨ�L	��8�87I[Z����~GQZ�Q���z��&��6���a���;V[1Y�ޅ/4���z�v�9�Бe��<�uæ������g��S��E�.��Կ�UbUl�l��^5Y7Ʋ`+6{C�r�$?�bX��9��Y�5-��-�,w��xb9~�q�C�s����U}n�d;V�0��\h�f���Ďn�/�5o��Y��u/��:�/a���U7��LA��:t����$��ι�__~P�yL��K��������O�Ͻ>�ݒ�Bãm[�Q�,��UU�JM7��*X���_��8���dJj߷�S��>�ҵ�D��7�t�U�vݫ�}����B�)�����g޺�1�
���QXo�:�Ë��ꂦ|v�uw�$U�z��έC���&����]ff��"�I$+� ��w�=�Ρy�����wXޫ�}���V�;mz}SB�k��܋3݌�:�΃��Utx��j�8�=sIW#G]�6LU���k�{��7�sΈ���~S;z2�uc���z}��OLsN{b� +�6���5�C5?p���`30;\�S[���qn+�y�9WL͎��ݣՖ��C��l9��r���
c^����jg\l�;JN��z��桵ʲ�Y���� �и�sG�-ߜU|j�}�R���NZ�߹ؾ8�{��eO�/ك��+n�{��M�5oL��I���<$na��^|��[��R�V��t�C�6[�jmwN:���z�|��!Xc!��;�e�N?6d���K#Yٿ�����`�����0`�mZ���Kx��*[�k�s*�;���(E�?e��V�޼y������2x�;�Q��q(��Ak�*:jr�#�:�U�������^O
ꣴȿ[�[���	�A��aڡ�.�nꧏN�˯d���Gz�_P��4�^Դ�03�#g�j`af�ݳ�_���=��Or01�a�)Zc;j&��>�������V��ޱ�`��6����  V,��xb�!�}!�K��E��]�#4s��x�l/��d�����o����CR��q.g?
~���P�}�<`�3s��Q}�=�����D͘�ŝ'=��U�i�zޅ'��yY\v�Eلq�%L����� P�`��#b��qE1�q�}��4�\x(�/t�օ[���K{���a��W���^+�9v�&�����:'���o��:��63���ѼCu�X����Ѕ,�;%ۮi��;�� w1sw<C��^�!�4~~�:��ƴ��L/9v��;�'�x;�R�	��C�7}�w���*b��W�y�_W5�\�����^^#����/ T#�g��#Y��=��Y�XOw#���_u䗸�*qSE�WCT��f'�VǮ��3EBs�e�� �[��AE.�Ő���̀��x�Ͻn�؊��8n�C�)z�G����`��j9TGo�/k����l�\7��'��Ճ)Ӂġ�[m��
�Ɖ�<���o��'����n��~���p��
{YQ$�~��|J��w_U]g�$���0��E7x��3j�=�ݦ��Sxgz��ո��&^FS�Sr�}"6�_wI̕@������R�U"2"Z;wR�}��,�b�ph�޾fff�\�8� ����'1���o	��ǧ���6r���#�>LM��U��*�����f!ْ�[��tm-��`�Ր����^x�T"�X���	�꒧�[��{Ȅ�������v2��{�L|2!s0��Tuk
U�_�%�DU�G%���]ko�#�R�{۟j1/Y@��򥆋�w��72���>�0�4z
Y��v첖K�����>�5��!au���t�ا[Cy��s�J4�~[O�١S�F��ܻ�0衊{[ f(hX[�]b(�o�t�>q�˪۵Ne��/_~����;�<�}�]Hs��U|�L�]�E{6N��[�ȸc�t����DB�*𝖟"1�*�莧�������V'5H%[(���V�\�1w[��h�W&��-ʿ}絞�j�p�l�j�?(�V(�! YW�ȁ��f괮���oIڠ/i�	��p��ds͑_�j/���έ8i��"�T��S����k����¨��[Eg><R�=;2���1 ً$���m��� �8M[N8uz�w,j˗z�ٜpm�xɖxxf�`�^$�n΢���5��6�O��u���[�z��x���f�!���'ld��d�c�8nؑ����K=*}�U��jݕ}����ԌWʶY	���+t�8�u�1d>������r����*��f��竻�9��z�8�����<[�t�?־������m�V�
��[�j������$�f�3֥,&��Jxf�&���Nh���
B�K��l_�a�c��dz�'�}���1�>�>�kqp�rc����qp�|��-v3%9�o�Sw����vM�f���`�/�?������Fޮ�ˍ)-�AUSm�K����Iݶ�>�-"�mF����o*�؞eiw��oe�?���ùy|5�`��'JX��6elF>l��k�؋������$�ž?�P�*z������T4��W��^��4�7M�����XH����MV\�y�s����+Q�;���v�'�^ ;�������Hp�(?�0IX�虨�u����~��ʓ2��#�t��������PJ��W��b5w�!�.�51g�'_�&�1�`Wd3���>w����jƆAUM���ϞS�>廡��Iz�GRJF���~0�^�.z7�݁ �p"h��8�S����5��;�ngz�[Ţ�M����AY]j���q��;Tm��ˈ�'�D���.ϱ\��"��`8�ٟ�1�"�����9S��FQ���nb��h8a�NcI����~-[Z*��v�Z�q�G�V���ד�s�'��d��nݦ��x��ޓ��%�:�Y2f��d��"4����O'J�J�GF0�3�3V��s����O-���������0����vWr,�1�|3�2g�ː�::2 Y���W���.��8��;��:v���'Fpt�����cm��9�Y��/t��%ݢ<q]��=���K>/c��v�9'Q�c���;�ܶ��=����W4��D�o�X]g�i���6� ^�%�9�4�5ӷ�(ܙu��eٻ��*#/Md����m\��ٜ�Gsa)�u�v$��z���C_(ڼ�HϤ'ֻ.ѹ��6#m�$@��P�̐v�B�"�j��A ����v<ov<���e
�Uћ�t."x\���4a���>�W�-�un���ڀ���uf�इ��e���bp��y��ۣ��V'1��T_i��D��B@Ӿ�Xv��Nh)�ۮ�����������ZG��
���@PS�/���O��E?�EO��h��$(q�:�R<���E�	#$�X�A�����F(�BF*�a
$d�	`�F1�b��"�2b1��ň��H�!H0�221�b�`H1b1b�X�1�	���Q�dd`*F$X�A"���b1cY��P��R �V �R1��B0�@
�0T�ĄH�,�,X�����$
�����$BF* �@B�d`��"E#FBB0 �X����`��, �"FD 	� @`��$B�� � !�IBHD !A��*(@`����@B
�@b!��"�@`	��
@B*(@`	��
�@b��0P��@D 0��BHT 1D��BMw��+�$*@b	�$"@b	����$ �@b	�� ��@`!�$"5�`!�$*�@b!�$"�@`	��"���*(@`	��"�@b!�$ ��� ��@`��� ��@`	�� 	�� ��@b�����@b!�$"��$ ��@b��$ �
@`	��"	�$�@b	�$�@`��� ��� b�iҪ��*��@� b���"�b��h���� b(� ����@� b��*�@ `� 
�@�� :D � � � �B ��D�1�1�0�� ��1P�1�1�1D�T 2 Ha!"�R$!l T"�A	 �
�`� `	 b�#
b@@�E 2��& D H�A�"�(�
�c ���@`)@�D$R)"��*E���dF
0 �`)
A��c ���dda�F�db�b	����@�����PF1 A$TQ$��x��w�����`�ǟ������k���_��?�����S����I�?�������>��  *�9���������@� �
�����A��؟�����?��
���_�����i_�N�?���_����$��EaH�Ab�H(@"HE@��b!�$ ��X�A �X�@F
�$R*�$V���"�$
�$"D��"DX�E��T"	 �$�EXE��P 	 ��$�$��P��B ��`A� �@D� ��$�$H ��(*(��"H�""�����"�� $� A�$`�E�$`��@ 	"`	��F 	�P�� �$P��"!�$��$�� �$��l�A	��?��?r��TI 	 	DI����o�����g����~��h�s�]��?�����?_��g�wI����'���� @U��P���?;��Ȉ *�  *�Z������i��� �~����AAV� �~�����v8���h?��t�~�G�D��m @U�����~��!���� 
��;*~�z���xp���~����C���?'����~� 
����!�s�?� @U��u�a��<C��4��C�l� M��=���^���y�D��� @U�;	 ���SH�����~<_�%�H(�/�`h?�����-���w�!����e5�B%>�9�� ?�s2}p$O��:���������q�m8�ε�9ggk����.�͹���u��-j��u�Uͭ�;E��v�Wj۷se�77L�������q�lK6�X����N���wk�9[t[9�M�t7v���;��Y�N[�u�WL����"��k�f�b��뻷F��m��EK��k�ڪ��M�Fmg:�\�[v�q�wl�uq�;��c]�n�:�]�m�s�`�nl�n�Ywkl��w]�n��έݵu�w'6vnmmݹ6*�v�3����
����nr�n�n��U�m���n�u�w.�kv�m���\�;�%�F'lֻ��wn�X�tx  ;o_oX]�����+jݕ�v�'Yݵ�V�o*��w]Rfͻv���J���ڭv�ӫk�k/Gy{kYm��m��or�JW�����kݬ�ض�ͯ]�c�YCw2�ն���Y����l����6*�  u�>��СB��.����$(P�B�
�>���u���[�����ۺ���շ:�7;�{�jޕ��R�p���oW\��r[p�m�k۹3ڦ�j��ɷ8�v۶�z���Vݛn��N����Wnw�  G|QM��}͹�G�����y���kw[�z
��c�ښz�s�J��nw�z!Gxv��=+mD:0u���vGJ�Z�w��+]���ms����t��   u���<쮵;�z��*����(�w#�L�U���𭆵�v�(�v�j���uTk=;�XG[��Z��n��V�ꊽ��6�r�;MS��2l���ngZ�n�   ��4ֆ�*����B�{n�^��N��u^�H1�\�E�*�8��Uw�l�{T(��y�Wm^��Y�ܻv�Q�;j�I���q�hl�Z�[�-�m��|   w�%k(�ޞ �;���@%@���A�t���4��<�P�z��4���N������:@��{��CwoL��aӪ�tݍ6�6δV�ws�   �Ц�n��xP�V���	� =
������(�F
:� ���x 5�)w^������8  x��(C��M���3�lm��;j�wws���   ��)@o:��( �Wr�
U�^�UJP����/`C��q@��uy���3y7B��5��+�@���iN��h�q�Uk���wKV����   ���B����] [޳ǡ����: �sݝ�E ��t�P�h��J W=�tj�p�i@��{� *��n���Yw[����gub�;�fπ  ^s� ��tР�k��� =��=z*�� �o[�  罻� (*=��<@ ��w�@Pto{gh�/�"m��� ё�E=��)*�h)���� 4 EO���U(��  ���T �� �)I4eT�  3S�J����P�X����͎���mk��	��YA�|}vͨ�g � \،#�f���7�������m�1��m�6��Cm�����m�����cg`� m�������Ǉ�&�@'�jҒŪ�o�5Qa���Ti��ju6�����.�][b^�LMj�-YA؂�v	R�8)褚�!1��RTVkQ�+	�v6��>��#̸�Zo��r�w���6������R������a*���TP�v��p:ۥD`���H6J0;e���S1$v�� ��M�lP��B�^�[�"B�Pc
�ڻ�i��ux�� ?n�Xf?�+���e>N�|���l��`��+fkM,[�Qȳre���NM�kC6r�����C�GnE���jE]lz�+�G.e32��C!�3K��]�-z���E[�0�KH/Dw�j��>��]J��ѱ1MFXh�8?<��1�ԳPIі����B��MK+���4@��IN��x�>g[�:ÚL@Зi�rY�������p�h�	ˢ�Ash�n۠Cj��-���C���G7�P�
�eeA�g�	�:�s�̓㰯�÷�+��
�KE��C-@!�2=��p�/�Kssc$`f�Yw�,v�;��3�,+�iwV���$�*,h��B�A��䍊A�D�X}f�jжӢ��hUe���)m�u�'��T�*�$�#�m��;>��KC>����B���:O9yQي��1	�����V'6�vtա�rӸm:�ݗ+�N�R�1*cwq�M;R�����]�>�nҚ4)����2a?G�	p�@�M%�ɒyՃD�(��n0fMZ].+��� ���C{u�{��6y궫�d��!J��FeM)]���J�mӤ���m��tn��@"ȘXЎ,���ܹ��;摄M^��d��1����ӥ�4n�\P��&%�j��V#Q\����*R8���݃f���wlcZ#Z �5��RHٲn��4�'R�X�̖�w1�ke��t��u�
�і��Q�&C(�)��:whU2���w���1[����vOlY8V����*�J��3Lgf���i꺺u�˕��SGT�YAAI�Z�[�������s^���&������&�'mlՓcN7%�� {
Z.]�,^��F'&����[��KI�
�Y��A�����f�{M�OmSˎ���T�y�D�P]5���~��7<�ˏ@pE�/���.�:H�na:����Jj]��çR�g��cb0@m�,�`
ec�f�����k��SkkQV��/U��m�P۬M��,4[fK�1���*(���8ް��a;+vm�ͳ�4l��*�杺_�!��汬��zL-ekk�����P+Y�QB� �8�*��Q�f=89�*q-uth��e�N��[1�b��o	��{�����GY�d�v��kL�S�t��Y�J�A|�l����@Ӕܛ��:(j�զr�:B���W!�Ĳ��<0?~L4c[�ϦS�
4D�栤n,�TЖ�۠7rF�3�4İ��+���c�D<���7]cF'n �f�ݽ�1mJuqTK��xh����	��Z�z�۴�x���V�r�A��r�0���� ��̖��A;���n	*�շ�-]\�:wTuIn�8�g��ְ8����B��2p�Yqm	n���D*��l�]Xs ��\Yw`f(�@[�O)9��@��-V�1�5Y�Ze���D0ɘh�94;���
���
6�G������E�,���Mr��8��b�{��	m�Aq<��^�x"C�N�ay\w�Ц�M"�
y�"���xY��h�&7g2	�[z�B�i֩��a?\�qb�c-�%�t�b��rF����ϭ�^_Skd�2)�&�4����� @	H�
cя��x�I��y=EVZ������8�@�.�$$�e���eZa�繨��x���ZI�zû[q(���raV%�۹"/�A�t�a[�b%�|�<3i��7\�	t~r�6�e�g�[���.��HÂ5Yf��*�����@�wW�!	�8���^i���$W(�A��ي⫢����ް�R�mhZ�3a�i�sVGx�����F��8�����X��A�v�LQR
M6.��ƣˬ[Ǳ�Ci������?�5�R k0[��r�r����J� �Q���i��)C�aFf�v�t�[��Gw��pۋ�7C	q��yQn#���r 54��fK�bJ��mC/{��@T��b�^�(Zpf�2�g f�7�6*���T5)YO�uSnkݶu���t�ay4c���3r��l-�h'ȼ^��y� E:t�7�r�6K�v:��Ǻ�ϴ�@-Y �i�PS��e�.�k�"�{>��n-���lӍ
̽�-Z94F]0^V6��Hd��0
'7Q�jo[���QԶZ�'��<�V�^ۓS�M��FM���_�r���R0h�Q�D	�Gr�}�\t%]@%a��7X�j�k�^��v�U�˗B^�q`���CTb�f;d�~�ɆnI'���P�&���N��ٺ�x��Y�;j2��cutQ)�< �3w��Xh�t�E�CtЌ�s(�ͫ#����Lx�N��u�N���.�nmV��M���*|5"3q��P¥�8�m�0U˛��YÅ:f�e䙦#q�V�j�hIB�]��S:���J;�c{(�x�ijּf�U���0U��e8��k4�
HɨT��"�U((���7K��B2t�r�.�,8�xM�ཀྵ�)��1��f�"~,���3i����h��5W�(5�]��7�l�'u;�q�M6��LG"�U�q�#�pm"���m���5�r���J��	��P�{w����y$[��z�#��� ��[+jfG�z畹�V_��ƴu�X��siaI�
I��
%RKj�2���Q�I��&�b��e�C��Ieމ3S�E�^MN��byX�÷�F�t�[1��1������NSEǹ�7�V�y�^ܔ�� ���"��Mw$oL��p�9�|��m��E��������`ܡW,SX�V��*��1�&e�-�N�
�U���mܪ<ٴ�y1����7l 	�Q�L�Xޫf�8Ѐ�U�{�][��̨��)��J[�`Z %Vf���>N�`�C=\m˅�!���~@�:5�6���i����.���Ɋkcc5���D��f8�jxe�UQ���J�%ܦ�ҥ]�'s&�D�4P��m�v��I �$�ةhB���4�cw0��Y�v��%�ޅ-�˩� �Zf0B���E�gۭ+M��I��L�O�*�@�i�Óf�ujݟ���C��0�g�E0��[��2@Em]-tA�j�2j*?��V���t�o!�х��S�;1��k-3�ܓ�̓bˬ=Q�Mi���f�=v��0��)��=�6�`+�RYb���:���i�8��׭I�֣Y$�x���i���H5�t+��dFË.;�v�U�Vc�˼Q���l3ޘ���l�9�+Ph^!��e����ٲ����w�NVSSAѥBֈ�]iCl\XH�dӴD7"*�T9��Zչ%ez��XsL��(�]l�L�&H1a�L�[�h��wF���{M����[Y��]-w� ���fH�
R�\;���V��f�S6vSbL����v�n�z����	 �5,]ٶӥ�d���0�X�`u��#x���l2�:(����Z;�O .aq�nf^T����X#�l���Ք���j+نA��x��6K�j�p#���]"�^�G�\�u���	}w.fT3	������yJ�7K[8����H8�_�l*������E�I�Y��8P����G�>�>b+"L�������2=�`˰��7�Lg��� ��<`˥��Ǡ����VqU��T2�	�ѩ[��bթRsD�����Qmkۊ��5�:M%�+6�J��ҥ�M=�V�db���ښ��b��R�̳��Z�Ik!��̖W�V*Sv6�Lz�׼�n�r�M��r�!�5�2�l]b��J:ek�]�ڔE-M�~wZ-y��q�1(��Y0l��I�%'��oG٘�c!t�3ecȽ�dO���2����rܗ��vʙwQh�[��u���d��QSv̺KSV����.k�g+1��L�K}�fa�.4Y�� �2��K�G�\� 3���.�il:�m�|�ۡ�$��!Ֆ�*ʽf^�D[I��/(m[�i�K]PY6/�cq��"�i7-��i�"�2�3a5�R��k�֍m$Y[�!���bv�<���ך� #���G��鰵�ı���[��%)�&��j��1���f�P��F��+D��)>�4�H�H���a��,u���{F�Ye�
�\2�>���I9�Cp(X�U�Y��V�9QM��yxC����X�zUєS����J���V]@��m���ŉ�z�A�e���W)H��DV�`�罳�z��R{7@"�f�%ր��n�f��#�f6@��9��/*�a�Z;(ˬ��=�����J5W*�7��yH~�^������5�]i�����t�*�W���%��(�@ⲷ��6�PP��"���D�ri<����M+J��K&� V���#7�Jǂ�^�ǖ��T�K��rW��ub�	nV2�ٖl�6�F��e�К�]��hR�F�[HSD&���ā�%�_�J��#������m���tL�f�m���DW�E�����՗YM�H5d�y[�UhЦs*n�Gcu'y�)�`6�q^a��n��	Ǜ�V��0ʩ|<��Q4�J�PƤ������ҴC��Z01wH5pU�Y���N�8���X�K;Xi�5�y-H�!�B��ERHP�wl�nޤt�7�Ž��e�W�u�X���h�Z/ְ�Q�5�5n�����	�h��:Tbc"���б.�œou���Tx��֭��`nEe�qɱ��6ZLF��/��x�U�,Rm�"�i� � �E�H��	�b�W�'=7[�(̉RQd���N�^>t�-d�(=y�$P�$B�/-%리OM?zA���,��C�U�#b:/���n�0�.o�,6Tݶ��{�8�\��*|!k0�	36VR#�'F�+n|�f�!�kܠ:8�˗q���֪�)��H��r���M�z�0<����[4�@� Y�SB�;u1�-fƈ��jz�g�x�y9�x��-�V3���(,��,��_�Q˩j�G���L��*�	�D0驵�vȿ�H�RVPAh֗����e[�SN�����KSu.F�m�@`��F*���YE��ܠ��8���"�T���Zd?�X���&��K^�x�3c���N{X��L5�b����S�Z0U��0�o$w��+U,̱)H���X����.�:l�%��U�A4�
ܑ����3�le�NFp�4i���^�%n��^:Y(eǪR)<�t�nKAI�\�-��Y(7wq�oJ�{dqS/�5��$f�5��Vl�b׳6Y����"�1I�v�f2�]Iw0�)h��ʐD)I��\�7yz �ⰶ�)Ad'@�D$�.�"hB�M�RQG5
�;���)G��Z-�'�F��@Vky��hX�3I�i����,l���h�=�S��"�#���E��f�$)p��oK�9��8i�9�[�#�U�9�E��yQ
��M_�;�E��|����kM�^�о�H�U��Ik#Y���Ǆ0��9Ot8䌆�ur��v(<�O"O�yv�ǅ�ʓ��۴5��[�A�݂�s��Uœ�K��nSDs�CQ�>����)l�&� ��	x�� �rD,:��{�_zy�0�Ű<9*Cf��o�J���5�y(k�*���-f=f�*S�B[�o�A�1QQ�Ir
L��6Ve�`^�Ib�Ť8kL�p8XOule뻰M���bfD���ix���Oh��fc�#�)������e�����\�Ц��):�l̆����}�q]أ%�|m�{>V��Z��	^���;)�ԳU��P5n���j�-� ��Ʊ�,jù��6`���Œ�w��-L�1Z��������R�d�uۭ%�	�;Q�lYX+6Ӛu,ga:�^�`�F�!��ͱP����r<�-̈́$���J7ȭ��f�\,66)���ʣ�l�l�Qb��y�D��Ϯ��e �)�Ƥm�NT�.c;���PҴ%!�U������LM������&nf=Yp�1^�6-����;���.IHp
Ym�'4�==���L� XG5"ǹw"A�n擃)M��j��n;�9��Ռً,i�,Y.�oD����\J�/��kl��LՙRSUy1?�@#�P��u�qn᠘�b'O��(�N��A�*�[2Jc �f�JG^�[��[,�$֘��`2���[2���kb�suĕ`.ʲڎ:X��&肾
��/�7F8�{Â�I��%.�t�=Sm�l��[P�F�Ѕ!����C[���/���kH�^��2&�A���"�����{v�vk�2��f^
VYGE� ������D��
0n��75�Y�mqd��b��d����M[ܗ���!br�[%l�)��hMX�y�u�J�9�݆Scl ��̧u�Ί.d��h���A$�j��Vhy5����=��q�Mvm����d
�[�Sj�Tf�R�T�Y�_V3�S����ٍL�� ռ"�ѷ�j*�H�/���ل��-�1t����.�o}�BN�Ͱ	+��z˻6�w�r[���o�軸��?B��suov���cȇN��6]݂C� pi�����]>z3D�^#�.�����p�u��5-��坱�|���j[��	B�`#��b�zo���Q���E)�pV0䥄[*>:{09=��/�� ��L9J�0�u`pf��n���D1baZ�^�xI����t�(]pa���q�I���*)�C�x$��("���"���ynN!Ke�$�l���}Ư0��[;;��6�b�+�R�8X|&uq]��ї(t�&�g��3{������DP�Hu�sد<U�I<P|v�mpx�[�x4b�EFi�5� WTo�����V;ŭ*��{S��\@e�&�k���	Ӕ/zM"�:�o:(��Tצ#�$l ���U��'�S����	����\�X��d��@2+��[4'۱w�,��ʶR�W��g3�u��1%�n.��ռ�]�u*��tt��u���pÉ��Ƣ�9z���>��؍�|�.�n��䋱��:�xi�
�8������S�G�V4K9���k�@,���ler3������R��C��4�5��`�SB�\��ls�b���Xv�ݹ6ų�F�-�v���8b�|��Lm���.���ݗ�~ǡ��Lʬ@�c���O.�� �MWr��a��A���C���X���6��#{�(e9�s{1"֎ rO�V�i������b�׼K�z4��g�E�St�����Y�{\�n醮!
1u`B�]k4���aͰ�G��V;.$������v�4��P"����M�k��xfK��t��~�Q��Qy[[�s2�hU��
�Ȯ����y^�{&�ξtS jv;�m>�tW΁�H�S^��2�Q�����D��>�mfDv�|�`��v��Ȕ��5�{5��|�����{���􉫱�B�_Q�;Ԁ�7��V�)��q��c�E�d�Fk�:l��t��峕����[�/m��7`�yq��M)Ǚ���K�}��^vt#`��}n�75sb��t��+�
Z�G����G��
�_Q���s�r��7-��cR@��}S�ȯqp�3�]��mH-t��J���-��'�O��LK��n���Ov� zַ�����.�N9��X��1�Ѧ{}9��^�FF7���.�p%֗q[�pup��u�dB`Sggz�ӵ�	y�x��SLI��'�H�&;������ܖ�����w"5^}��1ˇ��!��ҰQ���"�o~q�7p�O���ow0�ɣ{!a���tN�!��u:��n�Ty*��%��č�hN�d�2j�/�vTYAH�[z�8��n�d7S{�u���Fp�t5�'�2>�آ�d�d�Xh2�Y��X.����
*��6�~ٰ�x�PQU��Ԭ��M�q7Y#|�u�p���]�;.Os[������#���G���:���}M��K]K���7%pԦY�Q�L��	`s�e�b�����<�q�)D���i�hfMg���� ����g:���sN���2��ޙ�ɌwG�����G��V��K���p\��{���.�����dh�g,�Z�Y�m��V�K&��V�+�e3��gZ��}��f���cM	�ս4��0[���v��t:��r�8����^�}s��D�ц���A'�[W]L��"�7\U��U��v&ۥ���Jugu��/\��-Ga����T����6[��>#��mf�]tW�Z;9�ݵ�O0{7,���l��Ʒ�wz���vK�-ۨ!b,�
�(��r�4�ys����w�rv��6��=}��Y�p�pҢjdq�ћ;����[x��-����(�r���":Δ�#�0X�K�ǖ{����8u���^�Q�eΨ�L�h��T�WF�*����!��5n�F�ˇ9�/3(�̓��p�1��w!��z�tz�L��'9��T��6Pw��Ҭ���Lf�])�(w.n��[t�]*T�Р�Wf]qޥ�0�ﲉy$|��tfL=O)@�s*:ccT�d���Ԇ��9�	D�qX`��k��Ȳ��Vܛ/�[}�6ϽS1�y�]㭼�}���w�NH@�2�X#ƺ�9�*86f~�_"��e�3��v�o
H�C���S�l�&��#�1�v�QH^cit��n��FuK]m�����ng��2]�զ[��|#���&w-�99]E':-'�w�^<6%F��i�S���ߣ���U'u�D4	�����Q���'6��s/3� Ew�qm���h;�ƨ�ݘ���ca,Q;�k�[�_P̬�[�%<���Ռ$U�ĆfWd|>�N0��=�4��]xpåw%.ФU+}K��:w�ɻ	�����,�8H��	�u��b���q�K:e�_k8�1�^36c�y5�/WX�"	+��'6X�ʅe嗃6֨��f�փ		�*۶���n<�����8:��]Z�b��Z�L���X����%�㻇D3�����P��댛r�`n����R�lM��I�m��W��Ʊ�I.��Y�jv�hK5v�A�W8�4s�8=��܋��b���Φ.�<�+�k�>"�糀�sx�_>K�v�U�����6�[���S���	!f)]���l�x�]��rQ�4�q���|�䎆WZ��qi��2D���`�ԉ{t�6&n�g�ddꐾ�قK�[B�t��* ��1���=K�9������FY�a��Ι��e.����e�r �ȑ�" �*�����]ݛ��ΠH���u�K��]��zl��Z����|)U�O�(����wpށ�f#�ۮ��u'K�c�>�A0R�1��������4mŨ�Z�^9��3]�`q۰rW����ej�^w�����ܴ�����`���p2��ڞ�ٸ؝L�W��1OH�0�̙4��{��ɁgkԠmw`�m�#N�m17���1X��k�r��Na�@��z��J�-��U��:�G�큠,�B��]2��wM�.���g�� :rB���p��g,%�jm�Cdٌa���.-���Y"�!���}{����ۼ9ߝ\�ol<�g �(��{��Mu%�ts�C(9�0n�VS��������m�e�-�{��W-1b��k�VI~͇[c�w�]#{'6�&,a��c�I���ѡ���vl+��îwfďI���f���`� �����2��7:ӧ���Tj��E�j�<^�#������/��e[8e��z,������l�w�vz]f�5�t�F*aե(�І�o��7�_}�.y�Au9�vW�Ay7X���U��]��T���Ǚ;�w|�;�q����Uc�|3�Y��c�)��N��gӟq;k�3�ĩ�"�0���Sj*5�[Q�80�g�O�r>�J������Gg'���[��^�}�ԣˢ-[N'Qq���I�M�욻Y��c��a��b����D��5�7�v���&C*��:��m !��F;E��I@e[�Y�����}���R��L�k��Z��ՈJ��hW��^�s��t������1�]n^�n��%%�H�M�Eq�Ƿ��)%:,^��R��-19�g�#�)_�����Uѽۦs�B5���jl��u���W)��^�����ȱ���3Leݾ�E�:�ː4q�S8�K���
��;C��b�{�ƾ�;^����:^;�_+J��=�]�	@�X�-1q�$��������D��&�Å!:�5:�A��vL�b�,S�V��:�Ä�
Ь�b�q@v[L��
Lml��!�:I�3Z��nﾏzպ{�wTK��:��2 �)[:��[V0%4�;�tZ[:�
�u�,��$�ڝ�.C��t�[[oqhg�j1[6�%��p�J�t�f׻��j;���V*q��%nȠ�v1��N���j=��"�����X*t����ʯΌ��v��F[���������R�R�};KF;׮�VZ�nnA�P�%�h��sYװ�F�����m��U��R�I�nҦ�cV>L)X�:(�����Zk�no��#&"gi�#;�٦��ӛ7��r����j��Z4�gT
 N��c�P�pXj�c%�t^V*?N[�@N�<9������������&�;hӎ٨8��c��4丙�Ֆwm�\k���V�u�+^:�[����6�3=�b�B�'���[��6�JŜ�a�[�OFm<��XC��� ��=o0�
rd���N����xStY9�����GW���z�[�R��}#�j�ƻ
��<dP�ݐ�3������b�Pkto=�Q��֐��A+ć	���b�:Ggshn��SUvH٭���keX?�F��!�ժ����C�E>C����Iw�]�ނPl��E�S)wv���Z/#��{�˴� ���Y� {m&��*�u�)Mt��pw]4gG�-抒�l_we?�_oo�D^���~�'v� �F��)?av�ao��4ˠ���@L�Z�WR	T!�K���C���Z�Rk���kV�����e��º��ʰ@��j��;F��5ђeu�km����.��݁ػPU�M]ţ�櫺)��˕��֦nr���Ʀ
uD�ˁ�_S�.�u��y�tq�n�'.[���N����B����ud�>�d�C���^�/`T!��<��)�K%���z������M����(�d��V�b���l�8����{�z�d��/qd�X�{zP�e&^�O�'ؿz/`��M����O8��$�� ]cEeu�v�d�ܮ: ���ʘ�b�]v'peu4���8Н���8�}���ϭ�ӷ�ؽ��q��f��ћ�����ܛXW�CN������V��1�e�^P����_�Ѵ���se��[c}���9|���|R�n��V2���;��{��ɦv�.J�x_i��W)� ��J�
S;�V&�Ϯ�4�8�2t!U�`��+x�������;7�]+X��lJC:=�=e�Y�ʆ]>���MY� Z���o�ol<F�"|tQڌ�[�ᎥQ�7%]��f��1>XXɫ�o����r� 	�����he/������'5�qq�B��5�n��[��fs�m�q4#�<���,�����x��=c�}Q�w݆�K���3�V�����]Nӱa�q�5�t�B٫�ֱgq��n��!�Y��j�w@N�c��FzcM��ܽ6 X�'��Mk�Ի���kVr�V��Uu�f,="z|�r�o��)-�΍��cQ�܍]n�y�T�(>�\O/8�{D\��9��ϦP�*
��R������Ɔ�Q�v]3]w(7��-�g�`p�bai
�Nc �E��;l�u�#N<b��zt�M�q�vs�m���B�{f�u	M�0�u��Z0.�A���o���@,�*�e�r��N["�TG�h��OweG��A��6��^`e�vҋ`�޹���}Zr��g80�,:ww���9N ��[��n���}��Q��u��!]NJK�=�߅��DP?y��:��:���	���z��%�Z�Y�mmp��K#��ʮ�����v�ݮD�
c(�F��l�
_����4xE4W�J���l�>�7�q\߱kK�\x8��dc��q�ø�ε����Zv�
r��kB��.p �OSVhu�t:���o?�JSj��SԲ�L =-|��D3m>��'nh�����z��w͙`��8͞���Gf.}��U��$}���޾����]ޞ�r�ɀO"�������%��1U�vu�kR��8�C� K�)7��)�3����t{w5����+��*���;w�vc�¬���k4��E2��{[�1�L[��*B���B�ux�wF�ph��+�|�s{/j�L�ga�ep~5��w:�ym�j|��7�ns4�}�×������Ȥ׏%��t±:�wI�g�GxG�5���ʯx���+��o�#��<=����5#Z�J�}B�&�l.�iƋ��k�j��� l�n==V��Õ�:��p�QZ����EI�8�\p��1�乴 ���ݚݽ�����D�E$j9B�Tb�I�l���%|Lw��ɠe�t�Yݼ7=ޚ��+��%�Lw\�r��\3�澮
	kX���.s��c�v�7V{���{`���*�>w�^P���BĚzh�����GG:ԅ�c�8��yOi�_p@F��[��������F����u-x��-�gϸn�=6�r��.��.c��y�&��
�z�j��\��5Ի�Dkł��:��6�]NʏVP��6���x�d
���N�n���v�eC���|n�o�Q���B��	|�:��F�c���1{��-��ғ�8�vp�3].�k��{@,vLu�:e8h��c��f|�^���W%C�'f���|�JS ��,��c췮(�覇��ṝOhĥݷ���Ʒ��Q��f+��!����.�
-5��p].��{���l�ֳ��z9\n��0LO�ـ���A�֕R��h��ϯ��f4��_$�U�0s���G.�ms�)�ƀ<T;+zp������][K���7�8�K���$Y�V_U�!��&���|��Z�utoʮ����^]so�Ν�4���,[�nEV�D��]�X7���J4�;�pw�_}���r�/�m�|�z�f�l9Ղ>%v��'u��U(�'oS1�����G=^yF����M��w8�[���Gb�]C�@���k��b̆�lvP�3���%�&	:�,�Kg�;xX���dz�F�t����,h��^Z�6,�X�]n��F���%�}��h��wIl�������������6�c��6���׳��?(���_K��]`�>�Yi�E��A].������S����C�+1�[��=����K��=�᠎ӝ;ټv亳����� ��'��X�J�B�َ�h�\ ��9{#i��)��P���O���m"��6�1��7�>�k��qS]RN�����h�y��������Y�$�S*��[b�z����u.�-����Ч�"Hw�,B�̜o6+�Ά]��22���ח|��\�Ws
�"ܰ9�`J��((<g{*�֊|S�:��u��"V�(���%��U�.^�L�Δ�<�lj*̨�����kwS�w�e9�kR�1>��|����g&$Km����|'�!�����J3l��Z�S���	�ˠX�B���D!��Z�V�<j���;sj1�=v�m�NU�7GFtdA�2M������ѓ��L*��[�M�W[�>os�7z�u�V��z�w�9��̀]C�KvW;ޑa��f\H������c׀��kw/�I{w&����=��М4�dl��W������N���˭<���'9b;�ɕ7�gj�� ��]���%�u��.�Z�<��`8:�0ܾ��3����5z�!���yz'n��=�e���p���ô�tT"}��c�}Ӎ_V`��q^q����]LZf uГ��eE��.6NT,M���}z�+o�̎��]��p����on�����	�S�v��7�/W�N�#�{cd��i�CCjesȻqv���Ur�����ٗ�6�m�@#����y��M��f�230h}}hR]�����3:�3NL��\�9;e�]L�7����v[�{�1,�@#��\��f"���3�{;�'�yv���RK� n��k������}}!�&	ד�[�U94Y�ٞ|OY��瓉�y���b��ah�y�S\��_eI�ZX1���Ւ���z��g��q�����TKAA�<�G�	`�=\(�[u�0NMlǞ�x2�<;�Z��\�V]���^�WP�6�*UoU�!�rj@iN���h}ulR����h�R8���Wk��U��hJ�hھ�W>S��R沮d����t.G1tM�C���VS�zp�xu���s�?�$;��8v2��D� =��:�o�n���	�r�O��v^�Ǹ0����F�Վ6�bdo]cO��k#tʫ��Ke�Mt*\J�2o=�/��0��i�-u��ql�jc�J�oh�g.t�K��)�y���C��:g6T(6�ͥ�Aዹ�G�Zx9W8�E���}����m��C��h�=��[�4C�+��H�*�*ֹ�[*�-WW3�Oi�� �͘{�"���D�mX���q�M�c�LĴ�/0��;B�ٕ������^&ΣDY��C����W�81l�/���|�Х����̝ݎ��;b]�����կ4�uqE�ؠ�p¦K0M�gZ��9=�z���1l�J�ᬝcT��Z͌�Rqw v���{�Z���i;�T�S��&�i��g�y�o;C����_gJ=��K(�J��Ɔ�C�#�Wv�϶�����8��9���l�Y��8v��뜶��^vTfl�<n0����U�l�y��� p����9��ދFء�<Kŗ5[�tr��)4�[����l�{uϻ1�{�/��K�6^3��Lv��Ӎ6�hU�^�e����T�ξ�L��)݅���^[^�����8\Jo�����Z�Ȁ_6�vY�@�H[�������F+��$�=�l�1v�(B�oݸ��\�`���f������F�2�<p�uŮ/Tt���r�I�&��c�����ͬ#�k�������)������lJ߇j;��.R�j^�.���Y��*��������-'�T|y�b�1}�;+�;�yΓ
��M��gw,�R���셋:�6Y����t�&%p��4�Y�C{��U�5u� �H�x��J��
N'i��Xt�令�o)�Ք��|�TF3�|����("ew���-vWu��+ "��ȄN�sT�3�Ӑi�3����ɓ-@�7�щ��}~�Χ��;p�x>��<1��e�� �N�_�'�ѐUm��c���O�N]�������t�a�xa�o2�F�]�9 f��w��,�,G;,Z]]�.�mt�EgV�J�YJ"o
=H/�㲡��E�>g�S����iCxLt�d�����=�юu.�����s�l�Z�L!hX曾��(X�������#A<65gG�JaWu(������B�N���;�i�����x,yx0�޸��hT�V;{��e���s�BV�7x��^*�]03�m�����'w�Wt,��x$t���S�� ����4)�1��{v�Z[0c�}�����pŮ�O�.쬐�y#qЩǮ+ʷ�2ú�Ei	5��Nn��MKf]�u̲d�_O0
lwu)��ܵ�6��:Y�7��k�E�0�A�d�֒['��.D!���+�AJﻳ�������9�j�-1��E1�7V�x���q��X*%v�`O�3CB&�'�ʱ^ٿ� ��HҚiה�S!��|���0r�2���A@�YTSv��.��WW�Ӕo�&�oE�+�:�)��F^�A�΢�^Vc����I���Y9jυ��Y�.���V���3e��8�+P�3]a���d%^�:�r�n}{���P���h��9gA\�Ӵ�(s�ㆌ;+-�:r7�V.���4�v�tӦ&^p��lZ�ຬQ�Jo`2`�= l��[<��Qv��n��mB�LY2�#:�����L��|�wu�[LeY���J�����hk�D�S��]^��%u6qfYf�D9�J9K�p	ܬ��Ѫ�,�-�u����g_
�9��̻y��H��.Y�#lMН-'\)�����U�媸�Vn�X��m+І�&�=;A:]��	��
��v�NHJ����Օ/U?��͓�E���ȗDh�-�u��IZ�Mn䧪ġ��K��20�(Z˫��ƅҸ�9nt�pzb��k,�K�eX��Z�����
`�A|B�&hn����J^�۸LomTm<���h+���]��:H�K����6&����y�����ΰ�[�#ڄ��33q��A� `�S�|[$���X�'��Wp���7{M�F���&��t���M�cu`�)N���*�!`�y�oU��D��o�-�퇏d�k��T�p��	�+<r�0c�4壙yw���;kq������)���#�#-u<���uZ݉�W�yÓpķ���D���P��露�>�U����	1:�g�4DH�4e�U �r��$�(�D���YÒy0�-iF�ݦ��QxT�{s.����4�:��;%V͠���u�t��K�Ve�������yV�Z�$�A�mR�`�Ik3�v1x��x5��݋���5�+u��hN��<|�TU���@~�a�'��<GSҤ3t<s[Y3Y��eo*l�o3�!���w]�"98��)c%]�ʞw����2V�^Da��P&�W�|���f\6(D�V��a�4��݊E]�6�gw����'+�'u3��l
��S��x����OG,�������S��2��6��r3ƍ�r`�&n� �����.^�2�8�ˎo�d�.n�y��J�4Mv�����1��t��`�i=�S����Il�%J�`<����N:��R��|򹹵�:�5�������At��b���f�"�&�q��}/��}Y*i\���F�7�nqCJy5署��#Y��>��̺|�\W}1숁�zM�=���u��8L��`��"|�q�Y��Ɯ���*�)ZçC�GN�ǔ��v��z�9#ͅW�n&���걤R6g%If���k��k�XN�ل5bX�ؔA��[�û]0u�7��1���P�e��'z=B:a�y�
�Μ����͞����w0cY��&�����5k��d������F��)4֮eJK8�ڝ]Bqu���tߏ�԰(e�S����p�3��덉ó���Վ�,�iMM��r-궽����-n��PI��c{�F^�� vO�i��P�G9�4��;��U�!�\뺰�T�N���:��N�R�K�$F4���^#����ܢ+m��e9Vi��Rl
�I>7}��o2����!F�Z���+W��(p9J3DxXU���`7���oC+�'g=�${���3ӭ����i�Fr��xc��U��-A*2���yj	�\1V\��ȱN�'h'A�c{e��;3L��K.w��k���;�c����
f�}5��	{c����@v" �p���Л�z�櫆�- ��2�T����i�Yݺ0�[�	\�$O6j0_i���Y�Q���u֥�ὪPƝZ+�9�����C.�)^�ʹ��뻈�q�2�4��8�����Ok��.:O>K������׆A�h���x���qɯ�̅�,�W�k}uzNY���Qb�:�w]�c���c8��Մ�ќ������+O�FJ/r=*��b�t�ٌ��|�MYaA�*#n�g��OLU3j�UѤ�xF�ASl�PjU�=ܥ��F+�(�d��r'���*��=��2�^k8|����Sm�݋T�����������|��q�݈�=�������u�f����Q[/�8,˦�����f�E��˖�m����G��}����;�E�k[\�fǝ��Ѱ�dH-!�xq����]�_'M�.%���]�l�.sf���䑺�v����� z��D������������L����#��D�=[Ji��6���=�N�K�LZ#��N76Jx,hՖG�)����]��u�އ�g�s/1Lrg�])VSȜ�i���[�38mI����)��8�@�˫��C�=ʞ��xqs"�ۨ���W9���}�pi�E�Rb�]b�P���K��� P�j�ٵ��gI�va�L�ؔ#,R赡Y[�/,�H��awMɕ�q.O���Fm�_<TJ��7�4>�%�9���-N�4m~��Ο;z�k�Z�Q�%�2�;�)<!�P����Lfix�;s���A�bw%�f�+]�Ո�Ƅ}O1��(P�,��j�>cx
��U��!.�������MkR��nn(*l�3�V���`4�8���ӹG5���۬g4y�M�V��ɡ�6"���N�ڽb�%�[{����}�5��{.�`�<d:2�%�k�t�dq\^Sy��.���8�l�U��7XV�ݑO/�Nu�o�7H��8�ǻ;�������
�2-��5(�e�ř����n	R��Rt��9%�Yi�C��}��,��}Ҧ��`��&Է�AQ�5�<@)��
ͣP����g�Mn�p�qQ�pW�7��� r�	��Q��j�=��[ud�=&7]�&LSz�ا�`��.{�P��k�z��8qO��v�|L�1�+5=�Yn��޺vZ��b���5����閕j�o�CY�T�C�89�S��
��;�tr޹+wƨ��VN��:Ѝ���Q�g4q��I���Iu��8j��e����ic^���B��6 R��lom���f꓉0�=,U����0WJLeL�c�����)����iV�eqR�ypJ���Z!F�t��=s��
g���!	�f��s�i
�b�kNY5�u^7'A���;:U���h��e��D���}�.��)��N�=�12�e�ALW��<;B�{/0�Eo� E�Kj��H>o:���a�B0�vJH�-������9��X�#S��\6�n����rs\��en�t�[��Z	ʼ���u#�]�O��s�Sm�|�u#w��u�Q��J�֑�}�vB/m�����S�)�G,HtJg��ϡ��=�*,�tZ�[uw6�����ɻϦ<�:W
{{e��o�}]�+/v��7/�/�2nך��*���s��Q����m:�W#��8'�=���/���!��_+f�:fb�KPM���lX�[�J֨�jNg����^ja3�N���i$a��� �g(��B'�̂�:m��܏��ik��ev(��s1�m�FTu��]��wf�ys����Dc!wj�K�l��,�<t���m��޻�-x6��lp]��g��P9�����@��˔�(����v�u�&Kە��@ �{�.��7�H��>�.ʡu�}O��Y� n�8)�����.�3�E�������3C�w���9����0'�B<qu;�۔,��s���&��}�f�ق�s�o�֣�o&5.��W��y���33\�ӊÝd��m�0�S
N��ݶ��X�$u�y�m+Ÿ�T�I�Ÿ�RR]8�}���R٢�M`�P�C3x�k��TԺo�v	����
;'s�ڋ �)�\��j��=�Zn�;�wΞge(���QZ�fb���b��!��:�Ǵ�.]LIu�[J�m.�[v^�1��D태]e���C/1�P/U�ͷ3���3D��i��e��@��'u�j|Q�z�v�G��c�F�(����d��B�E�e
|,��� t�I�(�u�L7z���lɩ�!�t��3��fR�ܼ��\�i�*s�M0�tI9�X�)�����/K�-��^8J|
��S ��L	i.`o�9������I�n�VV�����eЮWO/O\Tx�����ჂEG�p*7GR-�`���l��-ڜ�J�q����"��U:YWY�j�pڍf,�;��פ��sNs�3_d�V���񓫯ݟ��������}�����9�ixu �̨�
čF�o:p��q]#�^���J����}�U�!�ƚ�NM�6�ؐf\9�����0%=�$a��W:��I�[�b_C�+@l��*x�f+y��P����A#��s�F�]oȳ��*��ͦ�gv�_u��Ns�s�Ish�{�3��y��CK�4��b��^FnL�k���T�o�8�cW+=����v_)� ��ն;�Йq��^X�QT�����Q-�v��+���^:��<V� �%	����3�rr����f˼׉
�8b�DاsPf�nM���F�� 'U�[�����.����FD��St_)X)>�e��:9�^Ȼr�}��&%^F-Ѝ����X����H0j���L���<{)��o��� ��]g�����)r���P��E�bq�
��v�5�}�~)4ބ��@�&�:�y/kșyo�����^j��gK�v!CX`ZT�:�m��f�9�>�'k
wF��ء�>�X����,���1(�vGa���:k�m�}�itk�v9]��l�|3��)�w8w {]@�K�Y)sa�fN��^��$�I�ޞ���& �g<4��q
vSx�1v	q<K��!�u0ml:S4,Y�d�%
�j�.�S�˛�m;�&jJ!G��S�b�G���"���嶅���gd��0� f�i�#*�%U¢������
�X�*(���gYʹUW(.pE�T.�W&p���(""-B��Mt6�9U]�
"�UT�ǅ�*��]1�J�L�J�")�8�t
��N�N㹵�� �T��\���f��U�OQ2좪�B9ww�I�3�wR.DEDU���*�QTȸ����ǄG*y@��D=Nu$.\�`� ����(�ȥD�ʨ�Q�DNf�,��.L�D�<l�(EB� r��I>8�PP��^Z��S�y��+VTU�9���5(�պ��2� 9G'(�x����:��9Z�QQA��QUr�G��"�-��\���9���̧2v�E]���>�g��s<%o4_O?oe���/��,����º�i��V8	s�u2����A@�,��Ϥ�˫�j�i:�U17\zc�w����.@X��!��y5��}�b�|�d�B�h�B����W$���(��?G{:f`����m��^�^?_��$�ʁ�)��:*�ab��y%�m�enO_Ncxa� &A;�d�2���y�P�#R�b�[�\#/�1�^��8/y�0�{�=��|�W�R�ԫ'Ysʍ����m���!x}w�����N�K�W��7pNdy4lX^�eki��)����X�P8�_��K�K%��`���%���E�sai�,2�=B�&��	ޔc��-4�L�e�
�Q��ž�Z/D��G�ף���f=}p�^+�j���I�*\���c�/�
��|o��;+�gU
ۃTsI�/$�Ϗޜټ�n��^+�̊z]u]��o#Pl�r-ೠ�o�`�`����p����Č�J�� ��.�a�Zb]�}"��60�!��o%m�H�	\K�V�B��d�L��N��X�"�����!�.�i�ã+
t��ݬ��_���v���'Y{٤­HA��Є�{�1+�h��S�n�3��&�����w'W��	���"�/x3t-ou�'Ev���dՒ�� ƤK���P��p��D3�l[����9��ٍ��S�2c��u�|�|�~�#ݾ}�]�98٢=C�r��ҽ�/C�������z�эB�P�qn��XM��&p�awN�<*-
��i�	tE4�z��o[�n��h��I����}�@^��s�+�}܅	`��{qW��������9���{����N�N�l���y+lFѦ�J��u]ʀ��!�:�_���P�v+��k�b�귩�o�d�;���||m-&r.��'�zd�ҙOlR�j��A�>���QX�7�tM2�H���Mn�0����&
��w�Qz>`/s��mD<i�4����nj��nI��͑���˞F�o�"��[@I0��T��##���ԇ[U)4��KV9Jo7w�a���B�|��xS��I�*��t�o�صO�z�:���#�N�=��%�m�xѳZ�c3y}����Z�V驍VT8X6�U�Z�px��<�w��}�s��y�o,Py/d�݈��Uݛ��^��ox���ʍ��Gx�\ ��|/R�?l�=��&�\��ku�ԁ�~��)��g��O� z��)l0��Ŝ�*�� ڽ�*��dI����x��^=<�+��p(�ߛ���v�6��R�:�C+!�������R�E�`tR�S��Q�������+W��ÊV��'5�C��U�>�ܰ!�}R.��|]���]?q�%�䥪��t�,KB��%�\�[�F��O��{���C�:�)�=3�	�-��B�5��L�ˏ��K��4���l��B������a���� �X7՞t�����*e��/
#�"ڨ�y��4�S����c����~'�R<r�;l��f�L�g�2C)#L��S�z�
�� �Ufߞ\��:�x����[��Mm��=s�X�p_1J�o�u�s#�/�h�D�4�������jL�..k��xD8?�����WU���ЇXh�+��^n:Zx{N"�����-3�����j�{��C�
At�r���Џk��Z�44M;Yk¡��<��A�Y{��Zm��n��Sn)���}�SOE�Z��P��?_`���R��giA�,���^��Y�HJ�%�J�_�*�\/��u�=�W��TD��!-�2����B��ͩTf�1����:fx�2�.F�I޳��j�Ҹ���ws�s^"���^Gt7k-�*Tm�X&~Wz$�M�b�껠�e��D1���S����8�N���=�-�D��Y;x#�76f�`o6�;���� (k��oo	u/W��n���uP��O��]mp��U��y�|�(�vy��-aH[R�"����s�X��|��C��@u�^^�֧��rfY�҈�&��"=o���HsJH�j�l�&e���WD{�#�Q)�(i�8�
����	����O9_�wn��CĮ��3���9�n�3��W�z�_z$���v����^<d�K�k�;�Dz��X<6��cUbV��;�
�K�k�Z�O}���3��,�u���?�R��a��K��}lfRՊr0MY+-�4���;�h/h?��u���޺�/x�I�ν?7��◫��f_��{�k
���/w���lQ�3�i��{�b��^�l[��5��.Um� �S��7qO����&Uң�~>�^��]���F�v�����*pW�>x����ː���|9-�`�CWu���U⓷�%�-�vٸ�O�֥��L�K(�)ȬŃ@��}�T\�I����M�zgT��g�;|+7�Z���p %��~��'���/g'����h^�뽯�e/m���XO]Q�Br~k��xUX�.�0z�
OXLw:Q�u�*;T�S�Yy�;M����p�^�7��7�N��4�nht^�y@�Ou�Iyf�F�^7�+��s�=�;�ʹ{ ��t={ٹ����g?ggW��n�:a*����F�y���<����'%p}�e
L<��܇��휜Z3������zM74�>�����=K4A���N����2�k��d��*{������M�U�}�8���ZlVUe`�J��h��*�xydfA�C�K칌)d�E��z�r�������3�1َ�����FJ!���*�KJ�(g��R	���ĬG`�]�^;,�����ɀ��v��k���#�g����� 7�!��`�+�2n��טܤڍ�PN~�&�&N���G�A��^��
_�˃�14ju��xr�$�f��8����Dk��.ה=xFY a�=��ۡ�0�<|�
��g�v���־�iY�]�2ɗ�j*]������L��)|�P�jBp#�wf��,��ۚt+s�=��ݲ\����&�U�����M%���x�҆��+nb���7� �q)ݾލon\�-���\2�����[�[uN!x�P8�_o�~����홴���k{;ա�B�=����@BM;6��u� �_���NUr�*����p߳e���{;'Hr�Z:㴎SP-|%3g6�o�˨wpg��ƺ4K��j���u�	�X�w'����gs`������ }�]���#2}[�՗Mo�AN,�E�}]tj&����	�:��`��CW�g7���.��P�k�쾨(�����ڭ��3�Ib(��dn�Ξ�;�X�%�p �r�����[��$+�6Ĳ�'l�Ǝ
���sFg��B�U���P,��D��^��բ]�9xj�O�X=5N1!���DحūM�C[�FS�-�C'�8�����ʗO]su�o*�i(�b��縆\�F$H�z���`�!�n�z{!��$i�҈�T�"�hD�p�� ��̙Pz�uT��Y��:\ޗ�'a�T���m#�f5�^��X��*az=s䥓������*�my�sz�)�����uu� �x�Jq��e�q��;�������M"��9�}��������.�"��8����(N�������k���`�]u���	�xQ5�2F���'i���Bd�2����#l�{(�&����r�=��bBz4�Ъ�k��R2yQ�~E^�kr�Ӑ��zg���E�x��7ಗ7��+���_���7��y�Pw)�*���?z� ��z<�<fA f��O�	ڝ��r��<)�F�!��ߝ��Y4m�C�$��s����ܭNЂ������[��C-WK�U��;��9c�T]]j�,��Mmud�
��6k�������Ӛ#
ws��W�nl��uO���ӵ�	�4�m�N��[�ğwX;���N�9�we�i357�c�ǲo_�Ы^�y�����tH�U�<��	��2�L����h0}(�5��y��*#v�g��&���P]y��%�^3`늢N��yc�7��Z|k�2�*i�.��i ���D�f^��6���d���O�Vac���Z�u��w>���G�[�<ߘ�=:ǦM��{���XW�씪����Df!����jZ�;�G񮻷�=t�m��o.�u��Ӷ�� �b��K��qc}�.�{� �%y!��%���W�z7$�J���D�W/
�f��gh�{LbM%�=ȳ���ݥ�����G
u�e���ZdG�3�/:���{;z�.=U��P:�^�xo��s��Jv��D�	�h�Td8-$��K�5��9y���^w����{���n�kl���[;l��f��M4Q�EFܣL�������gȖ��G��&��"��夞��O�uP��F~iV�%�9�s��)Y��.��dxn�򩡼[�k"��f3wIv����ez.A��҄1��wz�z��4�W����qطRPY�z��:ǂ����lKP����
�<eQz=Ǫ
c�:��|��"��.��r�5^�x�H��7�'�Y=�J���S(+�J�K�$��o�&宕ؑ<p68��웍	[3�+q����]$���B�u��*��Op/֚X�����͠9���v��h�C�̲=�R��c�8�	V@���Z�*�C3jH�޾��f(�N�R1^�X��WY��T�e�����i�'�� ^Qhtb�w����V>:��z�|[W��3�������P�^��^<1��;��Cc�z�2J���(Z�tEBH��(YU t�����bÑ�ܱ��N��5	���NJ���V�B���S-m,���2�D��5/{;'.Y;���͑P F��{Z�N�K�z�Z�܈�����a;�W������
�b+K�f/��Kܳ�WF.�G��0ݔ8W�V>L��*Ԙ�zݹZ�a)<b�$��=L�q�{�]*��_{C$�q�=����r����o>ka��imf�d�&Q+p١��8sbkT��z�������>��/B��c��z���z>�k��y��ӓWG	&lhfrYV�X�hO�b�Nپ�4��M	t���z�d=�LL�3=ų���g?����[�^>]`��5�?�!�i�A!N�6��[��-�q�?z�_a�2t�d�sts��[�&��QzM#>�����B���s^��}�w�c&�*^�8��J(2=���@�Ϩ�Q�k���ng'Zw�з�p��1�R�^�V9��:@�l
�s��&���VTY�q&�.�ʅ��Tɘ�S�|mк��̬~)����)��<e���#��;��0�㧎_�}�t(�GO7�ڲU�pRsR����Tl�݌�����D����U	�^��+�;��_T�\�'�����ss���?F=��_M'�� s�+�83�GH��}{��H��yE�Z5�lʊۥ��v�1����X:����ZW�6��� ��Lp�J�����}&�\}1���ܯ����ړ4���:�*��A\+}DCҊ�'���4ˬ�d�qr��wI�j��A���ۅ|ÿsZ�E0T��P��>V��+̪��zd�Bц"Cc�²,�H���V�w�q��^τ��FPf4���� �$1�倒�Q�����^q�w'������D��l�{?i`ptL/��iVp�ds�=���� Νڙ�UE�W�n6��RR�������^A�Ҁ�Ů���4-U;�\+<}|/�$^��<��s��6�c=U�/����,U�r� �0�~�(���3�!����Y��u���k'M�M�u�ѱ>���a4ZKH�<mKFX�ysx�H����^>�c��.���)S"�����H�*r���М�B����WWZz�V�y����v���dzL�9��=4���|��U��g_Q�cU0&�����oRe�$�t/�º�]���F~��k�le��yU��{��@��I)�E,��xÕ��4j��n�hX'&�Ӂ���M��Jx���EV�^zj$n��c�G���t/����R-���n��F�W^W�N�ʤ�~T�W��~͹`*K� ���Y���.�CB��h_��V�6�*K��Z��/�/��Ӽ��Q�S��]��-M�����݇��}^�3��oLW��m׊�Z�=tP�`T���^.��?N7rK�va��鷧��|+��ho�����tX�K7 _x�:"�����ZKϫՆ��]Me�S�oH�Ǭ�'L�(\*�O�g+^�%9����T�`50*Ջ�v���{��N�o]�{�N���4�A"�Oi#L��D^�x"�^IHp��n%���Ve�uh��5��y�� m�d�6�M#�e�]��։�ьL5�G�)d�N���{������&�ǒl!%�8��� {�]�8ֲǸ�8�!�8.�Ft�����xS�z��wf̢�9|�H�}{DK^P�1�gsvv�Y���
vGʸ�A��fr��FT�F]�"�7d�+��9C4��Q����_F��Y��u�M�W�G���yt��7�(p\{�ա-8ѡԻ�M�M(��;j�%r����8>8Ji.�|)Vv\ܮ�aj�+��Z*bjQ�+r�^Mϱ��΄�v��cL�E�|��Uc���%+�s��k���K��Щ^Bl���;Wx�E�u���3�N�N�Em�֝iF�f0�����q��`�:����5?E��D�9Lj������Ӌ{�z�x����L-�YN�R�+�H�bEu���sL�IC~�=i�{g�;��xQ�fv�v�T��$����7J��c�p��M��q����1;� �R��lq��=���+f0F1VV�J�J��������Z��::5�
���(Pk�2�=U�d����}����<��9K��.�t���N���n�9��ɸ���e�v�E�Z2[ �0�hՃK&�@���E#\��k�X�-�+U���4m�Y�����b�;"�x7<�c��%�x`�j�Tϐ�5����m�B�^o�wxe��6щs]���F�b���:�G�2���R�Zku�$G�x�5��f7���z>���:�Ynj��[H�>w7\e�L���S]pv9�ҵ��R�]�t���l���w�RR���e_f�k� ��\�,����8�MytG�	��u9]Ǝu�-��/6ߗ�\��k��è5.�.��T`�v4�SaAH[	ܭ���ݼ1Ф i��WKt��E���mv�r�<,��>��o�sGs;�|�㈔�ӽ���W<ISWwO/���Ҁh볃���i�l���;��9[�r
��V����:~�OE�9Ӝ�v�s�w��|��Z�5H��3:4H��g}���=7�@���z�{��=���!��Z�l��O;��w=�����6�a�W��Z鐢.�w���"'x��W�A��\<���D���k�:�hMX�A�;���t��z=�]ݮ�؂W��^4z�7�s�c�{=00|�{`��gv�Ǳ��W)�y�+fa��D;@]r��u� �Ka��r�k{VZ7W��~�����5C�j��4jS/�wq�������������Ƞ|�.��x�ָ��4_e�݂�
�=ccZ�֤��U�t�v�ά��fAD�9��i\�s��<�Aci���Loװ�>�����}	^s ��ӏa6�iζ�5J����Ȧ���G��-�Άe[n���mq �94sU5}>��BR�v^�`�Jb�G\�������M�a�Q�z�;�9S�=���z9�Yg1��o����7�<퀠�H�xX�#�9ZQ��yi�A�+���I�Fl��|�8���+e_S�uƗQÝ��J���9:��4�gL����~�<4"��qЮ\�QgNG
�E򲣺��<.Q�܍*�]ۺաD��H�9��.y�EwW=q�]*��8���+��w�xs�e\��� �.��U�iet�C�Kx�q�������1��v���;/:�2,6�P:�'�G�<�Z��gNZ�I*���Ykws�Q|����BTR�C	s��Ի���=JR���t�;��Ne(�\��rC���j�\+=ҏ"B:2��TB绞�c�<{�.\�TN��YUU��"�)�Ok���&Q�E�I�Es�Џ>w�����Q���O��\��s�jD��M2ԭD�חSs�3�B�J�B����&��rx��D^pI�,��@�0� Nc��gz���Z��j�wwhh$.�Z��2�F����Uhy�:�1z�I�/���K��vđ6T�6�]Yn^d֚y}�t��a��]㏉�6<w��©�G߽�BO�roG��+e���~�������G��oHHz�hx���Mޘ97���v��zq��p��KT�{�������sU.с����(MU��߿�ߞ����v�NTߵ�߈O�'}����x��������=�x���v-��H~G*ɾ����~v+������ǤM��9��� x�ġU_
 �+�r�gu׺��dIK�|������0�A�/�s����}ON�v��{����'}v�����	'{�~�~?�c����oI�7��������i]�G;�}��\�����]�����5W?Z���z7y}{f���ۼC�����;���}?�x�Uǟ��<M�N?{ϱ������<���?���7��Bw��{K�`�N�>��H~&��89?	1�5?�����iiR퍢���۝��>�w�i��W���bW��7󾾓~!z�������?^q���oi�0��ϟ�zq��'&����(��9w����϶ˤ?_���= zI��?>��N��;3`���®��YP�Z#*�p1���C�9�C�����=&�/����<q8]�����v��I�o�Ϸo�ʇ�o�O��{�ǯ�����~��oO�~&~������y$ߟ �wfnp����r(�M0���5X��ra��{y�>p_�= ~$�����zw��M�/�~' rJ�����?�?P���=�Q�e������;۵����v��'}v�~�����ڼf=�z��`�h�s�l�`��v15m��i���c�v�|yvf⡥�O�w�����|1��>����O�����<�c���!��|���]�|w>�����x�U޼��<M�	7���7�99�ݚ�;�2v���c�pơ��ڮ�7cwV�fjv̠7�܏3o�=�>���\�}��=8��?�������;�?�������bWo�c�{w<�����}vN9o;�G�'���N����jk�?���(u�w��k2�q������(��<C�����[.�����;~oߝ�w��n@��?��o�J�]��/����P�������q���OX����{v��;^��߀~��������1�K��ك��z�D7=���`{�!���N�`9�p��/���t��;z��w �mIv�`�:��4�*�O.��]:�j-Fr����3c;˭��6쳨���4��i6kK<�C��׵e�G'L�]b�$-�$:ʾ�NM������x�i�.�:��;�'M=�����`�ju��>�K�_�Q�����w�i���~���zL5��N?~��}���'�'��|��x��$?]���i�q��8=�<����ً������Ů�g�dT�����~|7��w���ǧ������[���?�7���vS~�ɽ{��olڟ{�j1�.�ٽ���1vO�k���b����h�{���gq�=t�s"�_�y�۽����S��=�&�BC����7!����:� $�q�����~;r�I��&����z������;{��N<q;�����ی.��;���(7�;xL�U���敛��뙱���o&�O��?щ��?^>������]�����ӎw��ߛ�p(
('�z�w����t�������I	߮�|���o�z�O|Bw�k����.�.�g�e��{�ٻ���a���@�Ƿ��{��I����~�����H����;���<M�O����c�w�������<�m������N�m?��v���xt|���a�z����<<���.�1��]�+f�y��:���I������߉��Hz��������u��e����|��Sӿ]�����oH$����Ǟ�o��'��������q�I�������O��̦���r�Fe�V�X/x�FR5\~��L.	�'�x�|����~��>�������z?~������Ϟw��P�|BOϞp{��Nw�߿|���N$��?�܁�_��|I�<?���U�5|S�8%��:rO��{C������{����w�E����v�
?|N��N��[ro���o_��<����������NL/ϑ���zq����Ͼq�@QC�>�+x�{�.uc^�@�`��:�UH�������}�}�~;Ӿ�m�?<���=&�'!���I�BM���x~�zq�޷����}v��'���>ݼ���I�7�'���m�=y��x������.��B�X���fTԞ�3y�o���ݪ����w����G߽���ߖ?N>�c��|�߉��w�������=$���~n���>�{C�x���~��}Ǥ�;۴u�v�z��{Ƣz���S�ѳ�>�����H"�zb�=X���^k�eh���rH��Ore�]�(�ښ���� 2͌3��Q͛w�����^	4�����#���;��ck��Nuzc㳁�f�ن�kޡ2i#\}J�.KV�-f̉����Q�
�I�ֻ��v�wS����c�W�_k������&+�Z��^�J��X�N�E�0?�
�-��z���Yk�$�ҏ���`�a��p���)�����ٸ�>YD���I��S��@��M�RH8
l�ԲYk�`>3hO�W�L�m�lSO�4ЗH[��ѐ%^h��ݧ�����*�hm��c�gK��?¯�~^~�3�x ���y�@�a�l����CX*o��|
��z��K��|�tC�#N>�2��w�\1�^1��&�s��=iLƛHiX��E��w3��%�I�r�3C\n�&�z�+�텡���s�����M[8A��>Z)���ڈC� w�;|+7�A�\���0x��B�R������cbV�B+�%�����p����E�i�}pK)��8 ���c���a[��׷g)iR�>�^�4��P�����|�j��T�
�,S��!��s%�&���ۇ6�^�6��ypև����N�l��T�oxӿo�u��௟��΅-�V�\�?zl��'��3����(|�K��r���E�i��D�������i�v�)�*��ZjU�g^�B�p���ZY)����5gy�:7�i�R�gqǽj<�v��=���ٯTO��!Dc��m8��+jvt׸���.ݡ�rN���>�H
��0}�s��C�3(Us�.}���®���~�\@{"0��Fş3�hP�A�jC����Q0�Z�*�p��28Vx�����T����nwrì��_��R�����)yGJ�J�k���#cm�>�]u�SSu��N7�QY'>"�o�Ӈ���\[�eA��@KFǝiω*�s;�Y�^�S�<���i��{��
�R)ڞ�5��Ն]�
f!;�f��~� ��������74���V7�OFߞ5���m�#�z��e�z
y�<F�k�v}�F�W�T�us�$�0]��Aǋ�I&3b"�����sQl|�r����������'��G��Ww�hM������������=C�.���T/2qT,�
��e@�X�U��W��ꢝt=�O^�:���F,}�x��tT�����qۙ^��~��2�O��h{qb�ú��.��ȔUVKed��7d�S�fWC�D5x��fw���Nl�J��m���"�5�ɟ��/i�PT��YG�{+�l&gW^ݫ����CN�J���W���yΒ�+�Ϥ��}�7&�ej۝�ë=G&Li=�:�n!�=\��童��]�9�B�k��L�P��I�\�g���l���J���5Ն�u�c/���%;��i9;�ԫy��V)w�P�ı2��p�Y>ٜ�t�\�U��fm��U~u2���³qS�j��4�
h�O�F��ì��P������OL�/B�`�pE��)=��~Y��}��z�#ږ ��\��*D���C��˥{����G����ֶ)ok��ؽ���5�ڐ�W��;�B�=K����'xS������}�-����]Z�~�/d�C�w��{;Ύ����4<v���;
ڀ�qW��m�+���MxfRPPOt������u�Ӛ2o`K$�)U+i���/(�;�*ɸ/�7�=�>���Y�Ƨ��<��ΐqڜӆ��X%��lD�H5�ǒ�O�fTCS@�c��G��"�l�w��.�<��y�r�4@[�1��U�/�	�uw��\���ʯ�
`]{��"�s�+����M��7ӽ��V�W��z�/�ye��y�������[@I0��Y/�U�K(3�V�<�w��p���h�U�l�2�LW��l��<)��$�<b��7bޱf����w��6��ho"���F}���Ŷv�S!{�u��@�\���WF�9�:gzmt9ث����8�����a�� ��}������۝WsYܤ��Z���L��d:�
����7�Gn-��7:B���1����9ର�*:=��me繢B���u��`�M�}r�Qu��b4]-�y�KN�֝Y�t�<�t�v_Lbt0l�����0�'����C�e�� ���L���+���:S��ʗw��/Lb;�r��2S+Cb��Yu�ԑ�%���y�Q如,n\���驲�V��a�=��[�E��W��g�_ye���K��hp�����b5x�lK��t];30w�?SZ�~@@�a��9�G����)�R�~2���ơ�{ҡ�'R ����pk�&�א�u-��ۥ����n�}<��>�t]WEF�4�I�i��b��I��҂�C��N��������S��iVI/	�8��Lv\t��U�x��ܒ�N�M;/Y�E�����R�6��E3X�i�I�Pu�zȺ:�M��W��5F$_G�Bn��ܳ;����z��z��yd0{u ��B,(����懵��0�x�s��G��s���gT0l>��N�捌�^ �+�T�X�i�M;C���׺��.j8��m��׸�2-h]�V�t��.�
�{�y\�J=�L�=M_Jev�SJ��}���0Qo/]���I���K>��Sԕ�&��:�]�NT7(����1u:��)D�Aτ�	
���#D�Ƞy@�;=ֆ#a��z����"�)��syu`�i��Qwd����+L4S8Kb���;������Z�%Z�P�Ї��������^����(��H�������$c�4���\2rT%l�W���
��YU�}��ҩ^�y�E��|��l��D�4:=��avk�N�}־�#~5��y�;�c���@��j��B=o>Z�,�ҁPjC�~&���6"u�.�x_�CGs�ǎPݷ̊ņ�1�,�v��R�E��dJ�WK�q|��a%}�2Ǹ�'uץ.Y�g�mK���� �?zGyy���18�ꉯ]]��y]�[����#x�ޏ���E���D+�J����*6�r����ky��&�~`h۪u�j�*��	�
�2���M>ה5X�j�T�uఠ�TZ��5X�����/��q�����w����b�!�i�CY
t����������ߖή6����~5��n�������YT���L�@uT/���h���>�!������|a��<��oj,v
��|��x�ͽD����@/׵��̟�V	ۢX��nG�c	���}� =�v]��s�᤽��1n8ec$�⢆��W$��/�/Q�<�<	���F`��M�h�dE.1W\'.�dc�Ώ.<��P�3'o+wYܪ��N����D���]*�:#٭89M��o`�- :��Mi�5��y5�t�o.�]τ�D+c���qg//������q_Q��*:@�xa���4wק8��w]���kB�A")�KX)#)�+�-�+	�< '��\�V�U���o��`Ƀ��X�P>3�j�A˓[�\&��]�얆]w���`�Q�Fi9�o��r�����V8�"���B�N?�B�lO�S�S��ʍ���6<�Rї"k+��^����n�y�W��9#��*0@�}����������Soo^�;I	�m�\���<;٭d�2ށ���|�QF���i`pd�B�k���z���;�P��t޶Lmi�ɨ���Z<}�Ȭ{����ߙ�Q2z�+|,��j�1��c����t�C7g�����&��0p!����p8��*�Ƽ�����D�xq�y�OJw&�c��'v��=���1[f����D,|��F}��wMO%{��1~�������v���}틓D`�~��v�R>c�la�~�+�)c�.#yYsʍ�r�ҙ�|�Lg�w��6|.B�'h�t���S
y�V�u1���H�����%�k��Ú�޼��Z�{�I�P������S-:<��ڠᇪ�x{�X;��[����X��[AS��g�m����9�r�LM񷯕)_�U_i���}�C؍m����D�^t..;��-��ǌ:�����|L��|g�G����S�E꘱���f��ɩ�_��oݮ���TG
�(Gi������U~z<"�;9*��L
�M��ۀ�C�:�+��b�i��\h�9|2��}o*
��K0%���6{�'Li�k��3�f]ݕ�;�lbQ�Hj`b]X�*}ef������x�L'��]3h;�{����FS=���;�0��0��aT�}�9Z��)�^U�!ƍ�y6Z.J>�/��s�y,w�QV_搂���1�hٵ4��0H��{A��FY9�>�W�s��w�����<��Y���!}�z�|�]oQ<�gȚ��ӄ�7��M���<!y^��g�/ZQ�H�'���M�u�S`�W��;�Q)�|��އp N>A_�g���o��.n���紓w"��R0�Z,l�#��C:�a�N�h�`:8��Ѓ�U�d���-����2k	� �k������������o��4D��T��bB�!S�X,u?�Tx���1�x�iݽ�լ�i8*�m��vC��>�G~Y-�;�mښ�r�*u��e�'�����mf��D[$ E.J¯H}��uo;I]�7��E�+:^nu�4ۭ=l��A��|Nϳ��������m��`HOB:͊�������z^{�OOvC��b]zӖkT5��,�Ҹ,_���w��%�"�t ��6�%#�F����8r2|S������(]���z6�<6d���!8���]�M�y�z���q�;�<��.��
π�mU__�U��y����В)�?x�}V�IIeg��m-w;����3�=f�]����S�5�p7��j�^��i�⋟"�k���NT��KqW2��6���4�"�4��D2�j�@j�~g/n.Z�|%���B��M�3(�@4:�zZ��E�v��=��9�XI̕�p_X�?"̿g�k<L�W+���Y�{�zL5�z�Jz؆N�5�����؄�+��b�`�����.�C%\^�̾�k}��d�p��s��z���yT�_�1u�zs!=�V�+�{�p�)Pң�2���ۜo+�i2��K֝#�U]S��xG�9�Txo����jS���בh�5ʘ0QsR�1��`C��,s�����Z�ս�X3mT�9�þ�<}�����=��������Yg��,h3�cV��$]!r'Q۶@F���EI�P�/;�f.��2��o9�c���-�p֍��:�ݿ�\�ԝGg;nWlȆK�U)�B	iV�R��Nxc��6<|�ͫ�(�{ñ� �p�S� ��r�u�Ⱥ�fd���*�N5u���V����r� �P �[ݨU��fU�t\��z�]�h�����3����ԁ¹/hr�&m1�q�p��u��c;����Wjk��W.9o:��{y8�ob�ש�z۠�;L��ҋ6Ty�z�P�<WW�jX����.g=���G2���[��ծs��l�%x��p�0b���[�A�h������:��zP��vf[��T(JΝ��-QL
�VVS����ߞ���Jt3�uO���n^+ d��Gd~;y��r�p)���A�������MG��z�e��C]Ԋ�yk�����YN���y��k����6���4�cC�:�>�G��(�n�oފ����|)�[}��6�*�Bx�F�I���g�N����I��כ2X�e�=m���pjM��c�&������ V���g����Y��쬺r�"P<=n�s-�HQ���#a���orub�/���L�0ݼ�˖s��`|���5S/x�1��֖��MU�f�E��	]�`؜���p�g��ѯ���C�X� j9� ���l�.շi̤h�zq)���hI]�7՝yԱ��3)nM�Lx�Q��(���ö�^ǆ���|2���R�%����<�L�&VwHR�e���,uHH��ޜ�5r�Ч�z�Vp��b;��^���D�{�?y}0p��v���9X�a�G��1�A�khuM��]����:��!u��9�4�[��f�\�֚�7�]u�������16��bmu\g�;O�LĢڝW���7ݝ>�4+ՅK�˹SaqM��b�J�7AhN��"XכR�dN��^V�����IO'Ne����jڴ�DJ��eξ���#5�\�Wp=��x��F����r�	Σ�U˫�x�qd�,���c�K�bN	���������Y�������9&d�����vI�&5���]�Rj#ۘIsu��w8Xݝﮭ<F3����Jn��Zv�:�J<�{�핃�V�ջ��!��-v�P�����)S���w�L`��U�(SI����O�oV� �!Ψ��9v�]�F�ג��pa�[�����쁃{�;�I��-�X2���I@�S,c��%��ǅf'�jWej���N\�U#�h-p��!��A�vZ�k��S�+��oĈ{-�h$��xN4z`�_G�1m�m��w�xJ�O39�FP�|�S�v.U�I6^UB�3�7i�3���/��*��
�'������Seu�{��!��Mi!�͕+о����We�β�4��ˍ�����y���@~�h*!�T���S����]g��s+�y�Wx�ˊ�H�[�S��y�Z<��_<��%^��r� ���"��҂��Z�%��E�<�<'t�G=B�ϗ�^pUu�E2��+�R���9:]>]�H-d\�,朷��i�盥B,�@�R'YF�����<|��8��"L3xuЎ_�V�j%DbK>2>7s��R�UEʃ�^wx'�wp�-UQB�URSG��Ւ�U�Cj�C�S�:�rȋ,�e�ʫ;����E=�V|��J/aUȨ�wYW<��sڴO:�V�j�8��G�&DP]��MG1�w�u�K1e6�:<y�:���bRC�;�n�=Z��Z ��w�b�ܜ$L�"YYm�(�h2�7����۩�:�Z���(��� ����<�w�)�Us�\��.&]Gͬ�	X so.e�<:�*�Jඕ ����y�M�ꪯ��:���rz�EgѺM0W�����X�l|5p�ZrF��ћ	�DaY�5��I���W�Kټ7�bү`�2�}�T�]��������g��Mi~ļm�N<�<�h�kKl��Jȹ�$�2�}G�e�LL[A��N�ss�@���L�&�5����O�nMJRѹ����+U���eD�v�k��qhx}�k��/�ި+M\`��*����[�kY����5�l��+��
�Z�X��V �����D0��>}�x;��O`��>\9�œ��w�C�:nT��6���ڡ���Fj��7��+;wˋ��k�Ћ!�-vɵ5����'1��$ة���Z����˭�!��T{|{�@�I3Ź���I�c��2����j��QL��E�׹��24�������iL�Tn��h�/Bǹ���T�W5��՘C~�x��J���V��T�;�)��r�\�n���8m���&�S�Q�>����L}�5��S巗K5�?i�����>�z=q#D�Ec�1l��|n��14�fg]'�B�)�"�p�D�`�j�71)]��82�e�Y�ױ�y��b"gw@m���o4�ޅ�-�3Nx��Qw����R�:��Tءf�b��L9�{��M���Ig��_Fq�8$�k_2EE��>���q����ɺ�L6E���Z�go5�$����chչ�*�����[i�,��ޓ�Aبi�Dl�'m��ɦ
U�%b�����1EUx����ռ:���GmK*{\O��6a2��(K���i��gl*T]���hlns)�(@Vϓ�'��,IlY���D]�t��Lz�"X�*�V�������CrrF�!S��L����}^��k��\�#Nz6b�;�u�J�%JR�(ՋVM��|���T�r�����֏_��ྐྵ�b�*1��<u��b��L�l�6����ك��n�z2�ȖJKQ�2�a��G��	gG)�һ��P�_"kq �eNf����L�Քͣ-䥍,�R9�F]v�X4Q�,�V��P�Ž��@���L���1�(�Ph�w��òѢ�R�~F���� P�H-8TY�{v�tt�䷢O�3�ŭV⇌��շ;_H+ͺgg����Ӓ4sdo�'e��1�_qy*�i췵Ӌy���l����[?37���en�٢U��z ��i��ꈶJSىQ,6�x�u�FC�U3�� ��M{��mė���[��SHo��{JlT�[C-zhdi	.�y��������s}�b�{��#*��>65T�
�\�\5�Mv[����Ģ��}"�z�y��|S�S�~�{���������<�p||'�-�[���kYg+�|\�w8߽ �V6xfy�1Q�q};�a�h6�`l9�YUc��0AV�V��1K��4��S�{�7�3<-ep�(�Q�\ޤ�gq|z�g��Nl�{ӟ`�Y�RJU�dkee��m8��U_�<Q�t.���<&�|�,�{=ǩ{1�Za�>�.aU��+42�վ�1w�)yW���Rvϴ���v��x�ǩl����Yj%V������ұ͙�K牤��Oc�u>�~��U�f�4A�^��>�4Im��X�wM�`{h%�P74*�է�ۗO4返b[%�5��vP�Y���$�����6D�'
�\w���Vz�h�2�y��W5Q���q�r�;a�k�a���)��Wf�$3�Vm��WPp�:<,v<=9�6c�p
��%ڙjz�t�N��w>6���o35��H:P15^_>dK����a��n`n��ΙhٴLޠ�z欓k���'[W=�'n^OV�,��M���Q��_�cC=Ng�Q�}ɩN�,�y��w�+$�ϔj�{Rm�RD�P�Z���T6ǜ�C�A��^�id��hÈ�e&S�-2[B�m��yIQ
,s,�ˣ^���J�-�5�OH��K��9v>���E�~;��m���yd�!	v�����h�T�{m�{��Y^�퉾���`efw��Vy�	��-HIq�|S���{�4�ȪB|�a�i��g9R
��7�O�)�x`�h�r������tܧ=LI��[^1S���a�Z�anMC�ת��j*��e䦣���!x�s�l���{��^�td���8���c��A�w^[�;,��f�'��|���Ħ����#2�yRk$(lL]�ҽ���j��j0�t��m.�,+z� z������7�G�2=t��/Z�(}��	�˥v�O�d�����X��vN5e�a�h�k��`��:(8;8[�g}�'	 NWd�/wYo�}x����g꯫���o5�jՁَ���f�)��-,�U�Jn)�e�yL�=݈3Wv5<���ջ��Ԇ�LT\�-���q�ai�%P2�,��Q4ۖ���¨C�,���n��r���2z�a�Tz�T>�Ի|!�9������	�w$s�k��R��K�"t�
���Am3cv}jM,��{�6��p��闈'�?Q�{���,zs�H���у�a֖��[=Rrɓ�4�k%�i,�ҫ:��Õ��x��o/�X3���]��So3	�i9�f�T�M2�ث·,�ڕd\i
u,�}��e��Wjg,nR�8E1Lγ�h27�)��sj蕏*��S*-]	�Nd�<`Ѳ�8չ�����=��չ�����α��&(�N��6fD+/d�Y04��Q�FíN۞u�QȟIQV��5��h��/T�1}a����4�Vc���F������Q~|�p�&WMic��1݋B�.s�u�ʔ~͚�5]��fP�\rL��3����C�������-�,�F���&;�:�n��@�g��RE�͢2�� �� S�J�ה��b' ������y�����HlY�L�K���^B����,6m.pG�YW5��Չy�����~v��+���}�F�S,�JpJkZDZצFP,��1S0˳�hISVe+��I6���5uԮ=q98b氲S=�Qr��e��˝��*lE�w٫7ۓ;s�Q�Ku�Z�L�sX�5�Ck�td�R�������1�ş'��8��֧�d3xɈ�\_N�������γ�٫���[���U��k�y*��7�0��b7``����������r�|z!/�7.jgt���G6ّ����ѫs���81~����l��m�Q��(Vf�#rɕ,j�U��V����*.�Y�Q�B������5�V{7��R2�{���H�%Aj�c�v��*.��Df�}.���o{6y�ԼC��}�7�����l��̑YL�YU��ЏL��J2v��4���x=F���M<z�QW����r��}�]��E&Ҹ�+�i�N�'=��<=�O����r��ܘ����(��R�w]�;�ޑ��*���
��ʗ.U��,�Z����������S�C�fK;L�w<��TW����;{��jH*U}U_}[���G6z�l�d��l��`n��91洎����l6߽�w�m���9p�s�o'���|��OW9���F7]盵�;=�(��d����{���\RP�Z����q����G)�� 8�g��įS­��^
�����yfIcKHKQ�F��YֈpU:�@R�M4i�U�,��my��ݡ{���SmJ���W���_�pv���vy�
F�[v����)ĳiM�����L��b���/%4�ǭY�l��|)���ܻTcY������n�{^��Р+�s������&��[^��UW���@O*ݐt���5
�8���l�z�z0�NM�콜���cg��s�MJ��=����3&#���0�.����I�5����oc���}�����_����~�a�O�e:���d���9�&���d"�G<��;�{����7l�.ώ�첺����*��M�0���E7p��W��D׻�i!���_f�7n�Hhr���E#�>���&���u���<�վ�ON�����=����r�Uv���x�������;zN�銹�y���l�Y�&�J�n�N�����&M�dkee��m8��UZN��K�mW�J����餅YVz�b���N�U�aY���V���Z��R��:n�"�VL&[,�l���%�
�f1�Z���A�.�k�j͖���% ^�w|�s���j2}8܏�SD���X�$��4�.+Y���F�$�ҌYU���E�I���j���gJ�ġu����>^����m�������YP��
s4}�T�X��H}8�ʝ��W��tPA�������=�o�<">\���wӦ����ox@���c�Ź�,ܚZSTޅ��mjC-�$2|�����}�W��^�ඤE�	1Ί�E�e�+Hdw��ݬ�V�H��=5�T��Vc�b�l�*+�Иl=�x�8�TΥx�n{0�%�Z�OyF��/�r먵+}y��x�C�멝Khi=�z��|���(��r����-6����M��������\���z�u��]�]{�3�˴��wra.p�Y��f����[��dc�X�a��:�-�|涷�wv��0�w�}��!.c����r������7�DG�_{���T����L �涇{
�����yUL�zJ�&^��Xb�-���L䴊:ש�e�mF��i����2�W���q,	ܔ3��6hK"�2aģ%���2�q��3���aY!j�9����Z��]Y$�>�*�+ЯuT������3�q��@$~7�Z8r��.6�Q��[sf`H�K�T�Ό-#U�x{\~ȼ�X��ٵӵ���(�?t���#I�@�W�,�l����`�U*�0�l
O�&3S���v�SNw|�E^����ܨ}�u��g�[#�D֥(�,d���T�N�u{�,^T^�W���:!�ռ����۬y�^�lU�1yjh��M��w�Z+"�(�X�}��u�/���gGDtiй��K�lLAj$f\�i��1H��8���"�߰;����^=Nv;���D�.���
Vt�I�t�����+����3@������i�l�&���e���~��d��yP=˳����]�j�4�)�o.�����gw?2��!��,j|��3�\#��_Wُ;z�
<��>��AM�<i��ӫ���{�S�iK��������o��}��{6�<�#����}����ږVEϡI5�)�z"�r�䄧o"Z3�92}��V���g��:5W��S�>����}��۟{|�-7R
�H���¤����C��o��m�s�Q�,κ/�o���Py�o�鷪y�Dn{Ǉ�ŵ���Ɩ
���v�m�u�<(�KIQ�-qm���d�Ue�U��!5�4�lTE�R���%�í�2_�������)��6���qIL�NipJk[�"ֽ5�4��.��g��-�;7as_�s�=���s�W*���>�	Yޫj�㪫��*��2#�5�{�Rf�b���z���; �nN񪸓8�bl5�0�����u�Ŗ��<��F?}��5^��\3<̘��\S�?g-�wV!���5d�ئ7q��Nn��]�VtMw8$�����>,���^��P}��V� ���S�1	�q4�h�`oCS�F�<�ѹ�E�zi�e�1���o7�|C�Ns@��%w�Z�������u�Yn4�N�����w׻ێK�]��'࠘�l�5�����C	,��N�W�0�k��`�T#���d���Q������ƪ�dP8�h�h���o��1+�َ�A��y�Wn�0.N��X��w����^s6�<��c�:6���:�}��3��*t(1�^�i��V�ktv�>c�W��v���B��U�M��B릎L����-N8.���U'l@�v�G����ldVg\j�sxع�`e�ni[\�M�^�7���^݇�j��u��D�Ѭ��:�K�w�������VbȔS0��0�������G�6�����eq,�٘ڵs)COb��M)�A\$�I��#�*ϻ��٣�6��2�j	szgJ�9GX�7�0�h�|�Ea����!w���ˋE�6;w\����.����
l"y����3�	$Lݬ �]t��G��L>�/���
�Vp�qĽ�,WA�b{�鏻��[Z����zs5�p]u����ӄ�+S�8:�B�t�{��K��N,OH�緾�<��� �P���L'nv�;��*m�\��sl�U���P�J�:a����[hN-u�ӎދ��>��ʉ�PP3vȥ�򝋪z�곉6S<�iLμᫎ�#�q;MW���|�>��2��z\�1!�I�ջt�?�\3�.�Q�A����}����A�cL�^!��f�`�鸐��u�}����s �{�g���Ϊ��w;'L�;��9���;�xK1Ĉ�}1��{{��m��<̪y7���A�ȇ=K.+�W]���۱�T\K��8��N�	W��3��X.�BKY��ftYxa����{Y^�O`�S����k��ם&�1,,DON��GY��J劦�o�FI\r�]61&��4����}��ې�V���'оy5T������o�4\N{��rZ+���뉡v���l�O-�^{]��Mjzn���l?��nO�B&�.���ɗ+H]{�
7�h�%��<���df.ٗW��HS����)���t;�5�%$2�d2�ų��ɲ�q{\�ʄ��K��g)[I^Ç��s;�{�=ӝ���P�<su�<�xfLbo0�� 	H��g *ټ��|�e�n���_���1�g�J���{�(г|ǋ��uq��C��)�gn<��N��rӨGh��n���iG}�']cw8�)/�RxäV�of�ڻ`��{[Ƹ�̓����2e�q�U/�h�Jx�ӐA�����W�R����^����P��}R�=X�:������3i[�`���&,c3i<ﲎ��w�\(�`�so��gD�|;Rvݩ&X
�8S����[����u&|xr�윦μ��FG0�t�M0���39�-^xy���D+Ed��")C��������rS+B�RMJ3,��$�$L�^4�v[K)C���2�Qԣ"��Q'�s�\�3�y�1e��S�TT��+�L�VI	�S��F�y�p�x�EZ�y��E���r��Nek&X�ԫB�TujR�edQ���$'�N��2�%�S��.�h��a�F!Zh�U��N]�,$�Xl��El���DFW���I�TQ$P��BE*R� �'s^'
T.D�"�y�N�4,�P�0�),��hi [M�GQfqS$7R=M6�r�U�ez�Jrچ"��:Xh�,�:WICB(�Ԉ�S"�i��y�9��)idU���%����RBӄͥ����ʻ�V��"$&�L��D{��Hb��J9UEX������W�+2��$�R*<�樒D�
W���!+|�T�v1��}�kXΦ2ghu��5�Jy�T���Ux�m���4�����gս�*cG���3y�1�д�Ӷ�[���*�o�f׳��U�_c�x(è�{Q�=�L��7�z��R�^�G�����*��V����*.�7� �2.�*�wWY��}װ�gztӁӞ�ڧ�>�
�ES�h����
�Qw4���ٛ�.vMiS�h�C6���B�M#L�Z��H6B�d��f
�/�.��HiQ!�nЍ�ޜy����;����H��ns�{�3�_��s̓<�{lΓ�4��yOc~Y�NXg��/'���b�*1��P:M�E�MZ�uw5�	ǖV�KB�%�(u>��e�6ǜ�C3��,��fig��o2��[d̝�Ɵ���ʼ#��wO�,i`�	`a��tj�l3�+��޻�����G�f� �=V���/L�F��4�ZuLE�%Iȅ��<���+���1�G�̵ޫ���ؗfz���[)��M��5�צ}x�
��cT�ټBbIG���8�z���7��zG����Z-W��U��w;����+�w��R����f�3���=3)<��tz�H��8��L�����<F��p��u!�?j>�y���^��ڂ��o"��xe卵���N���s��[{�o3{�sp@Yd�1;����[@W� ��|��\���Y�໽W��5J�U]�a�ט�)�3��L��	�[������z������^��5J�m�ʹMԴ���i���#WKhe��ğbY����Sl'1F�U�<�^d�8h/��̵b��mZ���꼻Xo~�<#(�ӎ�u��&���p���'#,��nх�i�^J�m�5��c+N>e2���Β�}qw�S�*�4,�	��Ym��k,1bi�Ӧ�W��2�C)2�6C���t2�T������ܡ
�l��k��Zډ@�Q�RV��Ԋ���M���zP17�X�%���L�#"�'ӱ	o���g0E�挘/���W`V&�Ӕ�/V<��H��Ǩ���TD�ϒ�Է���9�dأ���{J�[-u��QP����j>�>PZ<��-���	��c�$Qۀޏrs��C�V�n��oZWXGk��'5n�a��j�[%Y�[R�j/
�iVC�D�+-3�z�n�|A��J�ȷa3ݺ��8�S���`�y�w9k��4]��>CKK�����|gV<�e���B���P�g��������Ve��9+L5�3�-
�Һ�zF���
H�%����m�B���j�9:i7Y����e��6�d���ߐ�yI�yL��h�eo��=l`F4��x�S ��E0��]-��sk���Nk�TB�a�3�/V9C���"�xx�!�epQ}~���w���M �}���h˶�ܟ���fΛ�'��?{ו�!>����9R
��7jQ�K,��媚r��/6�駐��`�d�b.*�k�# #.�@�T2�}�[��b^��btИH�p��T�>�,Dє2�(j�שW��kݖ'��W7�r �����Gp#FiBǹ�����j�kU��U�4U9�S�ilg���n)��2p(]�5=�kjXgF��RGٳ<���(�����.���͜~ՏwJ��0(]�-���q�alJ�PD��=2+��S�EB�r�x�5�1��Hrf��w�y��߼ǠFԱ~#e���7��m��}W;�w'{>-f��\"����5'J���a�-Sgw���g��A]�wS��
���}/F:+���Z��uN��B��wr��*�:�����W�U�9`���S��ke�a��ƭ�ҋ�BL\h,w=p�Z�9)�D(��`����u'�q mn��-�6RX6����ceWP+e����{;�3�p٪6_�~]��8MZP6��Њ4�/U6
s,�w2�`�^sR�1���V篜�ɸO|Dx��SS���l�i�ΰ;��﷯����c������W��r�^i�ħ*�����K�/o_.��u��\Q��&&3	�3nR>�5��Ө6��۹sj���*웥mj�f"��V�2�Q!C�b}�Z�l9��	�V��a(Un5���y�$�L�Ӕ�/^Y�X��	`a	a��i���r ���ޤ�"V2�-�\\lB����\��T��%�Z�-������a��0�p�|��)n!�>�[���$�g'��3�8�%6*b"喽�#HK.��
t��+�9��x��x*�s��ۃ�;�z~�73�Ѯ񯑤�$��<��6��ns�ص�G�yl� q���b�`s�X&�S��S������*Ɗb�vۧJ�r�ӱ�;��E]_vWM�ٮ2�.Xa�c|!�p�k��֩�a����\�������V��ޣ�;.��	"���yʨW,��^
����{�{m�IJ2����Q�U�3��,��~�f�;"������
�X=S�Vs�|5� ID'OI��yQ�/��G��UwX+c�bY�hV�6Xy�9V��Ӆ�_���������?f�ɯ�<�-���a��5�B�8u|{��A}��ݦ'`'U�k^`�j�:�j��,�dkg����8�U�bb�b�,^���ycue5D�N�-�1�z�X�ӧ|��mZe�+^T]̱�2�+�k~��"���x�V� ���������i�r�׸���'�9u�
g�f?W����;G����Ӳ�	ʷ��$K!e$Vad�ZڷE�\��%S{=ワ�����i��yH���:Q���<~�fVV�g�W�Nܼ����ܼ�)�����TkC9Ɔz�Nc5J!�b�����+˿��)�t�K��uI��G%_v���+i�V��j>��h,z����V ��z:�T��k�7rQ����h�qU���fS�²Fz_v��Ve\�MJ}oV�y����P�c�}�.��<Uǡ���;���\:v`i�g`e��Ӥ����o{��0F�O���8�y��גX����f�$JP�Z��/�CWΏלƧu��K�jy<)r�b��m�w~���C-�X�!>�22�۶�r�7S�h�k(l2gHB��{�-V��Վw�E�T�[C%Iȏ�w�ʱp%�a�n��{�e{D��ɫ��0�p#م8�)�Sl�^��ɞ������ߌb@���]�N�;Mi\������O�Ob~y�\�ܫj�\����hF�mjwn��y���Lz�%YG"�;#�g/��~����V3�3<�2b=.bx�tϞ;�0�gjU,'�ƙ�
�wV*f�m��o{73ݬ7��y��HW��@����	��Q��6�R�>х�M$�^�7T-T�mތ逊��]��I�}ݛ��J���hL�Z�lz�b��4�s
���)��>d.��!~�kB�T��u�� ��'�;��'�Κ2X���uef���S�k��>>{�=Ȳ$���9���~�B[���q��LQ�G�:ga�#��n�9�;�z'+�H�m�4�Yls����	\̻\����\��<����o�꯾��`����蟫����"�=�=G��}�z�j%	%�J,�85�lh�:���)Fl��%��8�ճ@�����F�ߗ5[���&vь
m��\�t��V�ܦb��+V�2�wR`�`�u �$�R����s�s1�ǎ3��<va���uՖez.X�K\��L�����g�!<@|�
�WzM嘽�v}I$6휫����6�d)"R�SG�q���hK[/e�H,"��:Ɔz�%�,�����-��6�e��Hd��ʇ�f[n�	��%"��s�x��lyֈpK:[5na��K6��i��NA�3Y��4Rlx�2 Ɽ�,���cC�u���-�gbt��e��A���s������84È�ȗ+l)魒zh�4���Z�2ܼT;�UN�9w����$p����	���@��SYLD\�{hdhfF�m0���������)����q+M>ǣs_h �D)�hZ���{�#W��*�uҴFC���.m	9�_pR�)f]�������]GoU��5�.�p���E1'.K;om\��>cXn,��uZ���{��vNd��i���G��"^��������f�+v��ef%��y�\5����E�bb%��IFO�{�[�{���3�z���mþՎy����e/B��՞��-�\��V��U�MKC�}0�4+mX��~�A�?}�筳�EE�BOr�XR�:0��j�IB�ݹyY"��ǖ����,�w9Ϋ�ˑ׍�U�Ub=^��>}��Υe�Ƭ���-]����E*=��灿[2W��{:s����}�x���ڪo�����C&�k����KY7d�PV��2���Ԗ�E���(B��Z��nM�ĺl5#>+��i���S}0�ăh�-�J/V;ހN��սӱ`TU6Mq�k�$�ǽ���-T�4����7G\���1kΰ;��+�Vp@��e��=��~������r��\�;�F�����{�U��X��\�0.;��\��W|�Ԯu��§7��Tcj����a���yr�]',\�|op��_��Z�~�Ypo��h��[����AH*��L��ow���Xo	�/��D{7^X�=1�x�`������+z+���X�*aVQ��z�.,�Y�u�ܞ�����Q���j�� !WI�8�CK���Ys-k�Y��Ok�W�_U{6X�&A�Օ��e�)�9G����`�a_�,��O��5'z�ZU���Yo�Ιx)�n9�B��KԠ�!�`t��5�*�����:.�ݸ�+�P���)̦�{�hCn�r]5�"����W���`�Gϱ�d�c�0��8�NR75[p֨����N'Ħ�\U�{hF�ʰ1۲�CmY`���wP˹hV�l݈5�.}XY	j)�%�����	z�%�&�M�A�z�4F��f13�*=.*��P�X=�Vw��Q�~��k�t��fډoue
�Q���ƀ������My0��l����h��m��xuIӔ�G3i�BͿb��YWT��̕�o�t�,�G�{a�~�w���<�n^.j�Wl�KǴ�g�KY��j�CL��r�A�F��QN�$�ɽ�^�m�kM�֘a�%�N�U��V�e��Ү��������dm�woK�Y�E­��=۴[yc7���|l`��l�8ɓ�Y]J���,�\|˰j�}��o'�.]�7���T�HDE�9%ޭ�IeN�}N�z�h�m��c	 s��i���������a��d�� ��_}U_}Sc~Nt>�������Y,ЛT����X5D�(�a���fg��ꦞ��l���9)�c�2�c᫁[-�פi�D�l�y{�
 9���j����%�vw�X�f��z�g
��FO[s��Ռ����	0�֘ZN���X^��^���*�N���N�+o���sj/3Z���E���6)z/�>��U���2Z�,�:�>\��P�:��6���I�
e��O>|�M��i����8����IcHT������"��&nf�w%a�3�z�����۫׈�ꈶ��=6�����r��q����7�+�EW�G����7i���S�)�A��-��c��O�����>����.�� �W�tw����+�x��z�G�=�����T��	3r�Z,����M���F]k�,ʠiZ�+M�ʉ$��3��j&k��R(�x��T�΃�"GR�Bsc��V���hJ1R��9�k�Z��G�w 
բ�:���,mjq�ulF7:VT"s��@���@:4�+�م���rť����|t�zk�jee	��j��
͡d6��K_,U�
�Dc��R���w#ǎE{�������3��Y�[3{��	E�.V��z���˰�P 2��w��A�����u��r=��qRFuH��lu�]L+��e�wz��4�Ͻ��$]8�靵[c����k�����~���ۼu���6cTPNY�0΃�VW	Ki��xpv�}���i�vK)�(n�p�;<r�c��'q�N�`�z��k0��Ko���ʹ�5J��b-<╂�,�9��i�Wn��D�v�Գ*"�\X�#Ȯ�t��o(�q����+�K�oe�G�d�zG&5$�)�����{�v�tT�x�z*�v9C��O.��a{�n^8z����c�}'/����V��X�"R��b+Tn�Q�:��Ҝ���7|����{��K[���Q���l����I`˓����C8�`�;9��7K���%���g�%���AN��7�T��%`�;�}ƭ�qy��o\d��{�܃��� ɜ��d��MWĲ[����wc���>�i�6+Q���3�>����y:F�:�z���z<؆仜�h}o����F�U����Z�o��.�Ѭm�7Y�7|��f�r���a߅���&�M��j�\��=����띵�vX���o����'\ũ]���k���
�\zoG(��l|�m�k/w��c5�Wg�V3�Y7�xQ{u���h�[w�"m�� �T���n{����J�ӈl-hz�(�Nb�V����z��gO9B2�hp@��H���Xt�v��3v���M=Ko$!��8������׭���:ȓ���/q�5��yog�I!E��X�5�++����2�m���Y�)��r��ͼɬ;}ģ[Ҋa�Q�i�1�;E*�Ng;�j��=P��[�}��˚�gf3�`I$xL�����rB�$ܹq�u:l�Y�w̮��� �iE|�����pX�3/�K]렺�=/�%�E`��2�񧂭������G{Q��y��gm#{q�&�>`OWX*ӷ5�ޙ�_m9�f��[���� ܝ�mӜ�0KYY"N��'A�MG��]�V���'f���K4���t"L1�pe��\jVa�]������v�t��JG+Z����\�H�u_%��؜�p?.��'�2�c��]/�}�gB���Zg��t�w;h���䠻�Z�ګ��I��j��߻�B�P���,�U:\�_˭އ�R��\�3��6���.�ˎ���	](]�7��5��@��oa�ث�(�>(�[����.�hf�L ;�\ஈYw�g2��cu�#� �"C*��Q�s�E4���͆��h��QyDA�%t4�;:�Ֆ)��NZ�iݑ\�Y���j*XD�%Z��gJ4�QU�A �w:{2"�	$
%#hm�Gvf�2*H�b)�`Jj'	ws	T9a��iI��-P��N��&W(#3 �Wil)-
4�"1-C�#�9z!U3$��6d�XD����u4�V���Y��aYi%�$H��Ş RQ����¾wq(�E���\L�A�dHb��F�w2�¨�H��8i�I�,�Q5V��8�J*��Z�a!sjU%jW"3eish��J�s�Q����=wH�D�"�*(���Ii��LA29�^G;�%IY��Ӥ�2��nB�M*UK5�T�Z��Ĥ*�E��աT�is��af��(�BU��*թ���9D!����W9z�SCiFdW$�ev[˸KQU�%VH�:CN�֢l����]�̖%��������&B*�;�V���D9��κ���)��NWF8��ND�k��9k/+�\o0d�]���l~����3^�����?�sZ�	j2�$/���ye8�d3��1��U���l*W��WW���ՅX�z��ug�x�k�犽��t��<m�ڹ�8��-��ͣ�I��0��'Г�����[F�mS%K6��Yv1���b����L��O9�/����:u��e��ŉ�i�@ʼ��j�x���-M�Qz�1���	e��Uo���ܲ��C�G��T>��)�x��czeV�cl�y��U!��m�f�J��*.�x�/�=�FDO���6���/��x����M��Wx��Y"���^��NR.�|`�>�@7�DL64><k�B1K�D�˕3�-
a��;�u�J�T%����5i�P|}*�v����;�E��Lֳ�%�'�}��V��*���੒�U�%n+�q�9y�Xg�/l5��S=j�r��zf��Jo)!�s�:o{�F�kf�'fC���1�+o�� ̉��|�� ��� z��%�neJ��J���y�#�:�'���qh�L\'Uu�`��/����S�y7~!�9��Z����7m7J�m=�]uՂ+��/�,1T�;R8b���&_�+N�u;&�R-2gM4��W���T�����B����
�ã�X�aG%��sn����s̕��x�w�u�&9�s�u���Ş^.�C���ꇡ��ڊ�r��������mJY�Bj��4�lTE�O-L���ֻ��9R
����,*Wz�GK�����3�`X���S+^����[@F&�yE�W��9ft��}�۞1��?n���2�竂|�1׼qU{�%�?:�����w����93c��3��$-ϧxÜ�+��M��j��Z������qd>$�Y'����8��g�?����0�,�G�r|�Z��h�Ϫ��/�,
˻�	�;u��f�B�Z�VMf%�wL��>���Yn3Yj8���Ph�bM�uS!�Y
JӶ�Y06M*�ʭ��ƙ�;���k��Ta�G��Ν�b���a\ޖ�{T�Jcl=[�KF�4��Z��RX6�������<����o�}�t>4aw��vb�}/w%rUO�Gk�{�fwS�|��"���r��x��L���\�陳j��	'�Y�%���5�e����������l��Ρ�󣹎�|��yӟ(���ڎ^��ݢ�r���Λrj��-�c�Y�����g��o7��7�W��p��vkcz-�'��Z��D�Em�(ה^��NR.�C]n޸ru�V�2�*�g�d̆m�@˖��T�3�يD�ur���{�-)r�Y�܋w5����9g�t����i�֪��#{�-�GQ�g{s�߽*h9�ח�';�<y>��*��r�5_:?^OW9���ڻ=K�����t�����X�<��1D(�ạ�g�a�`���l���{�eK����L}����̯T�����4�H9[�;H�T=z�f���Jg��xnu̙;p���T5[�m��X昄ة����9��7�1;��D��^x�����-uv�2U�Z�-�p��JlT�E�׶�N�*J�r�q�g�?yq�Ǩr�L��d���'CP�U�1Sίޫ��kr[3m�`�'�f+V����&�`3|vEG����W*�� �!4=�K�j�v'�.��>��4�2g��^�>e����J��������T����R�c���v\�]���+x�L�(�a�o�!�0�x��ͩ��2pm)N�'G/D8�E�zǗ���a4̧���KSkhv�ѭ�[(nm��f���^ieW��3Rƹ�B_�3�T�������7죺�m�ޠ�إr��h-�Z����Z�n(Y���|����o��C�;<Z�rh�P�{�i׋�m��SV����M��4�m�e������?�d�O7�MSy��;�Ϩ���֛a��oa��:�ʼ�j�+�>�:�O�Q�]ğ_{O.�I�o�߾�5R�<��m3�f�
$�%^V�;Ml��+#uUS�x�H���ciQw3��������Za�婢HK[;d>`ݩF>rv�񹾪��1�ʳ��/�T��W���=�%;w糰����5�vp�&�ҽÖ�^ҽ�T��.��	�F�9�V���6*mQ*X@�s*�/eyNd�,�gK.����ƅ$JP�}G���j����jMN74͍���k'��]nKS*Wx��He�J�ԠXsM���)�@ �0#U�ؖO]���+	�k������9*wo�n����=;G��m�(r�݂�k-G�a�6��Jt� ��Lr��n��O�iA�S�)�=]�ֆպ8q����{z�o*�,R�uA��o��NO��ui�|,v���l6���o7�j�F�)�����6G�h�
8%�ʖ�sv���;�/���n�jelm���Ok�vw�Q*'�a����C�ڛ��Ncnfb�3;���5'��T��ܩ=Lm���BW�.��e����*�Z�؂�2���_5���Y����i����`��>jm�m���i���j��-�W��zվ���~V0�\0�-�C�{��Gc���?t��5E��z=�#}�4fm�Ϭ��A���X��Bjo��F�fI,n� 3^o�Ea1vQ�6�T	�
}�L)b�х��M�J�m�Z���X��u��L��U��KV>e#'X�(���έϪu�z����wM�<�w�޸٥��̒��0�����:�"�=Wǫ�P�����ur�nlF�m<���YO0#�ׂ���fϒPs��U��X�>!�'��Ҧӓ;B{D�$��Hzu�4P�j��NN������U5L�ƶ͖M93�O��1�$�=;��*���(O:7�{��Y������s�F(���O�g�jf.s��$�y:Nǆ.X�VW{�ћՍ�S��z�K��d�
.K\�i&����������ۚ2�s1�W0ե	6��H��
�Vs)tGV�0�I���T��ٯ��o-K�C���e�l�Z'rκ�W���JU��h�K�c��	f%���ZT�>�d�jZ,�s3k��~��ʫ��G��[�jz�i/gM>�M�FLM�H�L�6ìhg����k�ż��Ps�o��pd��k�U�&DU�?o@�Q!C�&_��n3�G����nc�k���fk elK�ܒt�ȧ)���֕!,!>u<n3:�����5�	)�-R���5���z^�Ĕ�k[�-�'��i	�o�(����%���~���7��y͘��j�}�'!>%6*f".|��u���2��ٓ�5h�-��:�.�Z��b�i�E�V&"h���fE�i6�j�*�V]e�2�sGc3`&�N2P���/�K��z��V�<�x�n�lp�����?5`]R�1���΁=��&|!L���voe�f.s(W�Y{Tg�;��]]]\>"��K�RƑ�L4����ۜ|�/6��0�4oH��rcٗO��d��;OnVqT� �o
X�얄 �I ���KΦhB�L}4e���_W�}����s޿sG?w8ߺ#�7��fĔ{���ʴgQ�Gw�nE�75�w=��9����c{��|-z����Q����@K����#y��ϥ�Y���z�iL��b�e�Lj��2��B8�:c�����첹�ӌ�|��[�K�F�5�e-�se%�i�s,b��&[�Qj-�gN��k�Fj�=]�}����$��Em�(ה^��Nn2�d��m$U������/l[C!�u�
�-0�kcit�\��i�;{U,E�>	L�[���^B��j�PZ�0��^��'{>Jr1��ތKaa�����@:���T���RhRM!N��G�e�a�z��{ꔂrϭ���ݨ1���ͳ��
|��Ic�B�L����u�45|��g1�C�Ǖ�<��R��{�{ֳ'A�%�>$����$BXl9��52��Qa�}�nP�
�&�:�wa��ګ��M#���0,2b�/�����m�������쉵ё���n��u9j�ky���Sq�鼞�凹�Ay�:Z�8�SoA��.�����gt��ۛ۶����q�����4�n��Tᄔ�_{��ﾘ���*L��j�u�ІmՎi�M��E��y��YRᛒ���4総{48_���p@��dյ�3�p��Sb�B܈V:p�r}��]��.�� ���+��
�1�W�\����.��b�F��j˦|Vb�z�[`"�ݟ��Gd_�'{!])�P[���:�W�Ν�����f�Z�6����S��l�u���;������`5�}��h%���W�e2i�%�>鴙�BͶ�[>X�u�L��m��n��ă̅6[�X	��^����Z`Ա�ala��y���{�/>�3�o��w��'j�K�E5�M���y�0&Y��a��ÈLi��^6�2.�Z�63(<�Ĉ3;�׍k��ee7^�[-�ͅ�Z٨�%�GѶe:U/����p�b���p����T�rF�ln��V�D-5#L�Ա���G�׫}ۤ�IX;�Q���t0�斈'bڲo
�'*���ҝp������u�I�
���;G���:�����-����T�t�]�ū<n�9"]ˁ���h�murDLs��z�nbYxku��������{9��2�կ�y��-�mv�dsV�ܢ��TU�9-G]̨-0��ٹ���a��]7=�p��}�qg�:���{U�痦�����ߓ﷗����v�b�P�>���f��&|�5)K4nc��Jǟ+C&�>JM#�E�2�N"�>�k�Q��)��C֑.�O��+�f�q+C-�V����܉k���:Y���V�}������*�9v�n�sDZuk ى�ט�m�6ezu�>N'F!�~.W��n_fxt�e�7�[wvK����}��}ܙV=Z�a�B���4yBXl��2Y�]��~X������/Llx͞��nt�%2Jg�f�+^�<���di�׀�;�f����w��o�f��S��We��bb'�e������e8�zmy|��|��]��V�M��U����YQq�[A��Պ�BMj�R��Q�a�wYk=�9#�k��[i���5���O?�wu��e������������V�I����R��잻R��qR�ݑ��y#��9\@��@�7x�[G%�ۨ��^�Y�t�'�+"����l�Y;	^���}s4tj�n�����{������oY�m�%bM��A�cP��KEE�$�6X5,S�>�X�R���؈�7��3���9������z\��"��b=^�:��:���ʘ=���g��-tv�U`�{��L�Vdf��\dU�zZ:�7�}���hz�h�^�ԅn�nyUXEX)+H��IX4�λ��9S�(��<�.��9���d�$�ʔ�3g֦�%��)"���^��ng�u>c��]T�v8��c2�swk��J��jɝ30�h�î��^��zS}-��lW�c���7'-���M�m�����*e��*��u�K1�.��Y
i�9ٯ��M�n��"�w�6�d�r�P��W��S���>m}?v�'�6�������O<{~�{����ÙfF]k���DxQ�,�l�[��n���1��%�v��X�r���B��$B|6�!;,�D;sfي{L�<܂��׾H��x#U/4b�YRw�_cS�u��W�4�ܕ�0yZ�#�RÕ�&���*A�X�N��e�R%
n�����)D��v��| ���E�t�L�p_*�G�̻�6<me�3����O	���n��1���s+�8�_]m����,�6n�Ʒ���܃��d���jn2��3R�	��tZ�a)U��^��$)���*�e�į�v�^n7��	]-7���>�U�����/Vްk*Lt��&�9��)�x�B3�f-h.=0W�,A:K0���M�pb�H��'u��ƃX�kl�@��L=�5oj-Ł����2�*i��"�T%c��v���CHX����Ѵ/��u��h�*�f�v�z-��][�������eK�W��lꏞ��2�F��6�[���K����p7xf��J�(����˃�����������M���$x�^�tu�xT��{��1�;=)a�xє9Y�����:��)�z������$��{%b��hT	�l����w6Nۉ�^��OW�;T՚$>��]uś��h��<�C�X���uФyy;�-;�	!�:V��^M�lJ���N� =��`2��c�c�dc��������^Z�r�Yv█�!ؔQ��c�7�B�'���B�k���c��h�!�����2�'fQ�V\�8���j�uŒ�b����2s�JZ�M�:�MR��FƊ(�f]��{�x���..t+�v��/T�8���]�pl���2>��1��9�ݙ˺c����t�+s�w�}LZ������n�w��ȑdw�Dv�	\]�)��k� �ja��Ni�嫕w6��%eG�Ύ��BO-q�'΅t{�R\֖��6��k+]
b�D�4\��Q�F{������\v`Ȉ��������d�q�Znܔ1<�#�,V���f1q;�ԨE����#��l�����䫲lff,�]�4a{��G��5ۃ:O{�u����ܷ3L�jr�}��R�)���ꊇ^���S�h�y+W[{���Ӻa��F���WO$!`]m28�Z�hp��7�tˢ.+&lY�v�Q\xK�4�����w=�f�=�1��{n�G(��*�<��h��W_)uj'p|��r[�%��sƺ��%�e��4���2�Dih��}-Yt��	~^�L��.�VNƴ��]��Lu�f\�O���!_a�����9ۉ��n�X3p��1DU��40i���<��7��/�}���4g����Pۻ\8t���ܤ �8?�	���>YZ�>ޛ~r�1�|.p�ƈ�Q�:ԕ�5ƃp�óL۸rJ���X���IFJ�V�ʝ-���mؼ����>�&��Ɋ��q���{7V�u!����Ŵfq�X��dD��yN��n* ؆�wy!��",���9�Kc�rM��ot�?�g�H#��(4��R�E�[B� ��!(Q�M{�#�Qr��#�<9ʒJ���JE�-j�Ȉ�%I*/u��3�/1

��):efeXI5B9|��֦�Ft�*�D-YU��E�J�Qz.dEQ*�V�9�+D�VHuR�%���]41d��Q���-T�e$��b$,�iJ��xUfN`Ο;�R�P����TuR�DU�b[O]�.VsY�*���0S�'+�FJp�åVUa%F��F��ap���N�Ye,���	��sb�eʪ�TI
�$��A$�RPaY�i���*�|���@ʊ3*eY,��֠fhIU�rvB� �QSİ���i(q3Q��\��6Jٲ�4��q��$�4H)��� ��!$��j\*�f��DW-H�$ ��T�I�0��Y�7w=H�CH,�*��V%t��)2��T�F�V��.�I���*�nw*��������׮C�C������v�tL�q�ҹ��;3�tcKv�����y��\����ܥG��������<�������۔�;�g
s�����\��l��#(>X@�l��/-�.q�3�i���m7j���	��g�M��9^۔k��V^<��f(�͸z����yEyޠy�2E�OcΆ�\���Mbb%�����B�i�7FF�aD�o�g������{~2ETz\US�j�U�T������T�����ez.�;p1=5���o�tG^7��fE��z�,)a8��j@�0!�3�-�t�9N%����36�l�ʼ�/��#[Ds����O�bmx��1�;�������9��X��J���'�3	�9u[���YPE����n�������و����TېsN�7�pt�9?fΦw���MaS�S�1n�ڂ:� '<�7�5�7������w�hwD�ǹ��+���z�a˚Κy��)�O!�z��Ӓ_�S
�Э�Du��x��H3���Q�]ɞ[cU6_�B� s�$�6�����FG�{ή��wp&�ĕn��)/]��>�]� 	:fGmS�-��n%�sVGP���BӘ�r��W7��}*>�����ٖ���<we���X�o/$ �y����GKi�	um��c�h�GnF]ې�����Fr��/�ꪬo������^|]|̧(�[h�SZ�w*)�a;΍T�pBᾪ��K�a�*����uG�dn����-���U��(-�ㅦB-s.�Y��;=����K�˘��5n�5�h��:�p9+C�ݝMM�U�^�L�)�4;�s��z�s־�:2߶��+;�*�9�YMy!̳gN��1��[(��+��M�����h���)�̇E�;f��fl�hE,Xr3�������\&���Ht�|ON���}����=���n��kb�m��_Y0ns���m3�L�<�dw�k�X%��S׎���j�<��w�����T$�s�A�t��c�f)����FB�q�-�"_z��`�H����^ڟ�a��7)~=��L�6���&�yޠw�����{��#W����pV�6u���>SL,3`\+�^�y,��m�.�f�[bub�Cy���,Vy�xb��,߾�}����L@�o�C��K��H�%��Y��(c���#��[�̓`m�w���1�L)����~މ�z���v�U��wd���D��=ͩ��)f�S�fR���J����T�۟�!�Mv�­�R���_i�e.��m{o"*��=��ʙ2����֗�i
C(�IY���;�������#([�p��AP޷� 'WI�6{�vd�����#ȩ[�)��o��[FV��Yp`��j.Y��oy���V�����K��q:)����O;�5����Y��Vt[r�~��-�v��"�Plw��5�i��9;�p�� +�1-�+�z�jrd�iP�ƛ'��ϱK�j��&Q
���L��|V��'�ᑼ]8r��{��:�� B��š]���E�^�����4إ��BB"n"���c]�όd��U�V;���ߛ�+^���	��)��-�U6@a��zJޡ,��5��<Tu5�Ud�gon���3D=7gLp�n�M������d8\!;捔�b�g�s�X՝�2��A�ʎj��*��}�ʎ�@�˰�FR���.G�;�Ta�P�ֆ�wi�vdr;�ݙ��ߍ�
�~�.�X���G ������M��Ѣ��SEwD���lB�$<�/����P�}UŁ�t@e]
�p�mz��<5�N=6����5��w��=�P��X5\¡e�y�228���C��:���)�c�׏�2z���p�����q���}�^��/�6��yf���S5�^�2�\�l4��B���>�xe̻pb��n�/PH��g��ڒ���Ǵ�렀%�r�.%�����u4ӷ�inAk�+��{{v�|�0{)�9V�];�y;������fu���|��$R��v��x�{�0p\�i���N�s�*K�mt}=�8������w=�~2����Q�� WwK���8���>G�[?�S�fT����^o��iK��I�wzx@Șc�]3��4��s8��x�d`w�Q-�\��`F?C��:6����8�r�o�cxm�c�'&i��c���z]DU�����Ӣ�^U�����,�j�ם<N͙���	���Ӄ)x�)�_�ME�ϸ�;ܿO�j��_��p�·�k����ܕ�m4�v�؋�[��~N#��T4/�K��!��������jPe>pU�o(+��J��.6M�QԂ�c�nk�� m�:��E�ΉT��$&~"��3�f�.�ڮΉN���չ�6t��u�$tuO>n2�Oآ�k�+�u�����2�/�f�T:1��O^ݫW=3�WSYkT�خY,�ap�ĺWoGT��'H����R��Q6�D��=c��F���Sf�8�4�fl_�C��jy�����OGF�7r��ӄ7^���wB u�k�����+�2�d�oV�N��#Hǹ����z٪i�D�r��##��d����οwu����~V������¥m�h=��I#{���.�μ��-~0*%;�c�\������`�t$�Ri�X�X�31�S�J�/�%��Bz�`�d���׫�ۣ�{�Û�O/y@e.�S����;�9��W3�5��_J��_oo1䓝��?���ó�tK&y��N�2
i�.�]Ts��8�`�f&C�	
^�:a�v�������뙧��⛺dtSZ�w*)�aȐ��t1{�p�3-h������r_z�tM��T��U�I�챈w���8��P�]S\&�L���T�Ql��e�і�-l4c8�0���K��\D]g01��<+�;@B�Dg �����o�=B���d:6�&��?Ax}5��x�Z��LC�Tm^��z�W5��-�Ԝ���۽�@s>q����(;�r���fC���G��?E鬚��;��u:~�oPc�M1��-�6���;35�_��Y
i�M��Y�g��F�����K��;�\����)�8Řw�?i�d~�~S���5�K��_�#/��;�j�u�*���f:�8��j��ȈHS�1���lӓ�!�c�.�����vk¬��[C��A:Ư��3S���oL���gU��w]c���d�G	^1KY�Ԙ�=�1�U���"{ab�0wN4�7�����<�sz��7l�{n�ڍ�h�{�����gB�U.���_�jW�P]'/ݛ�L�{�6z�U���V��A4z񵝕o��qw)]ޭ3���5d
ζ��%Ƞ�=0Z[�����Y�]/��zҐ�U�[��>�6^���;ݣ�gP����jd�y�X����R�W1��`����w'|^�~��jݶ��FO�S���;L%�N��MR�p�Z�ت�/]�*�W6�����3��5;�3�j��{JļP�*���}���-oSEzL���S�`�Hjn�ڂ6���R����ۓ�ug�$��k�L�Mc��Y�ܫ�������}iJx�Y<��O����St�XΫ�d,D��|�.A�P�
�D�g���M��!`���([TAu�%�!����u����η4���n� ^�l&S�NR~��R��E7L'ym��`V1�A��C%�g��'�}�5�7�:*�V���/+��pg�{
Y����Q$g��e4Z_A�����P�sƌ�|>\�P�Þ�yJN����O���t50��m䣴
��hޙ���2��ߕ<;�,NHd�z�m��40�F��~�R^)�q�$?gF��� _��M���}M�Q=t�scS�w35��cvJ/9��n�>fZ.����:�d:y�gL9=(G;�[!M��u�&d�֖�3���2��z��V�n���Pb@$\D�j؇�4d.U�cg\����-Z��C�3��rî�קY��yѹ��&l<��3�بn�Gx��=�7[L����r����o� �<p���ݣ\klf�ؼ�D�!�^� �k+u�n%�}�轂��}�yg�nW<�"�/Lq�mn�M��M7n��ApZ�)�`hծٍ���t��3Y�o���?�D�w=�>{��DW�E�,I1>f=��{��iz�ל�*����k#5����i�!�ke����w��R����3�!���pV�6u��L��4��0TD����p\AUBcI�5�6MK$�6^��B��<��K�7�M����FO���9U����G���wȊ�p|�K���3;�_m7=YL)����~m�sz�����?u�@̚����������Xa7�7	8%��q8+ޕ��d�z����,��+:/�[���)���٨q�׵;՛�fwz0s+� ��:�7��t��|o��� 9��0Q�"�&Q	��ۼe19���eV�=OH.�#I�{*�\�̦-
n�T�m",���P���8�ު3�j;': {��+��=��]�:��q��g��h�y���~��L�e;΍T�sq�T�����'��o:'~_����E�/޳�:��w*n�8�[h�p�y�N��)�~�i��r ��s��-�3�U����B��i{l�Ttg�;��E����.G
���Wtb���u�����X�]NvP9�$���jE�u���g���H_���c:�%՝�kX����)�\��4	1�=��!D��(�Ӎo��<r�/���Z���N�+�S����O1ϡ��oa,\��]H��06�9�n�r"�4�L�K���)����l��Q�T,"�'vs����\g����?!Rvu��t�巒��)�:�4SOR��U\�q�X���,i糾�����Њ>����р�%�)�s���w�';g^�)�=�5��]�0�g���"6ޣb�;��_[EGL�䢀�0!�b����1�
���)l��޲�ORu�J��"�"g#����8���w��qJf�a��F/�C����:K~�r��H�~��M��.	�7�]��q;�.x��}�o�:���!���o��g�؊b])����<MQ�~Yw�jο��X�&��z"N����(�q�Ǫ_+���h�?{��^W���R��u��<~�G�fz��t'��Lӧ��-�{��"�֢�F�KF�yV�����҄�w��
iiLfo�x��x�x�b��B��J~yl���aN8�=���1 ��z��0�{#&r�Y�/���W{��#��Pо��K��|���׮���<��#Pz5�zjhY9]�OFOf���67j�1�=�7u��_z"�gD�i����?M�3���Fc���r�:Eg/�{���f�獍�UflS�ۻ�K�:9�#Jjw�����b�p%�g��W�Qa�|�-�0�pw�.�܍�P��*�e��μ��"QI��7;�h�}�Pv^،��;˺��
a����.N[�l{��@sA�s�r�m�f����ܥh�|��\qP���4*�|�f]I�7oV@/~��.e~	z����}'�a��W��Z[��cy�c�D�5��g��\!��\-�:�?��)���B֤8T�m�U�\T�g�=�r�s3�o�s��w���-�G��~�MgSSϭ%M�z:6��7m�D���Rٛ����Ҩ�W�u�b@��z����B'�;��þʷc�n�+͜���������u4(	ŗ7UQ�����Ly�\�)�C���n�dϣ���B�^���D��Z�gF���Jy�&�P���O;[�+���.�|��O��#��֡�ʊ��"X-�v��F8.�S]F:�`K��y9�=�Z��o�����p/�8⛻�k�k��)��7*��3�&���TQ3�h���l~��.l��v<1����!hZ��_	�yf��LЦz4���Ĺ�|���=v�
�4dƤ���૸<'6�93�WH@�Ds>��-�=�,;����L�����*ՑWW�����ף�
���:m����<�j��J8	�W����<�B�o��x�.�l����W_^�����#��&z���v�~ͩ-U�͵#,�q�L�Q>�-�>o��M�����{k�<�G|D��ߘ���.�^
��Q@�T��[x���j>h�b��t9wPP�0g;�9�1���o*R��Ur�W���d̽s?̺� O��߀�}~����fB{s�R��z'5�K�y��s��+��a�7��]q�dC�3w>SUy��DD�q8n�qf���M!`1�����)�|κ���i�ݳ�)�����;:g��u[�7u�=�)��-�d>Q�Zũ1��� �u_�wp�����CYq�j���g�j�,����*s��L��ޚ}-�7�_��c�E�/3��δ%���ᨭ�o�	~oMÝ�l���a-�:�=AT�_�T���U�zf�YPE����	v�Kڅ�'���w��D����==��D�lT��kz� �*�E?q�QZCL�<��%�L�e�xS{���FC@j#��'��"Ȧ��W�a˚Κ{J��d�m�����f��u�Ê"�ug���9)��E�C� *%�<��M��!X�LG9B�Qz���WkF+�_ X�������Ͼ�&�}�y���?`*�.�TW�����a��y�A�B8�8a6��t��F�j�_z^�ӓO��,wv*���8�Zhr\˹e�όͯ�r��?�$6x?L(��4��{vB���#�b�{5�!ޢ#�I�fY5A^̲ܺ)]Æ�Z���ňQ���M�ۘ9�v�]�Ң�{�"������4��yu��j�\K�h��(�P��/����ՠ��'����81Z{lΦ�ֵ�O=5�1mՍ(\������SO��׫Kж�\���o)�7����{U�D�D�rϚv�Yw�[;����ЏY�kA~	˭�Q�?f�<�����egv_�r���|����/����q�+pp�b�+"��lݓܦE�����3�̙�bL�A����$뵯	O�Z�y?���}���wY)��¹���^����G�qo�gE3�ruA�<�.��%ȡB�H�����e,�Ӝj	0�xtbPx,�͎�]�u��
uZ�7a�:�2��9���Ϻ�� $s�`X������Т�gn�E�o�/��~Wj8�&�d9�m]�r�7#�ݙ�61l�/mT/:FQ���@��.p/z8��{�[ۖ4�pk|!���G8 ����R���8��\��f��;��(o���y�/͟CD�)3��^��L�Mk��	iI<���A�Wɻ{}�x�N�,��� ��XԲ�<�z�(7� ��*��͔9��hܦ]Vo�L�&iW���OM�{��p�L��<���l|�!ި��P�4�dyhp�[��UO����a�+�ԼI\�\,q�MM�Z.-��,y�<�G5�h#� W�A=���)m~4��O�zK�}n{��B��24��	W5m�����K���.)<�WS�l�T�����O@W�
`�n��N�8fON��cb��W��������0"�y
��58����yqNT�y��efACzI��(�O6u؅9|#|�f��~x��Ms<�K����ѓ6p�L�n��N��GRN��ńm^,zB����;O6L����ޤX����Ѥܩ��̇��K��9Srqy�ܣ��J&��� ���F���"N��[��Yq�b��$Xk.k��C��Җ�/�����XÖ���Y��9#Kh]��j@��h���m�c�d�I-L!���\�>��s���;��eKx���\�&�t�[X��ɾ,���zS�ly(��a�BiT���3|Q8n��oR�죠�Awh�亍���*��ti���ǫ��:���� ���ʝ�4F��
e˫��K��o��^�& Wrm)�G�ƨh˺٪/������$O���;�44]6�s��V㍼�YO6���ea��o�-��g^R���*ˉsa�`x2�ȬLR�C (8��j���0�j���#����p{�!iV^h�2��wdel�C�����q��R���;�*jLb����o�5��gzR!�|'q�5$�p�P�h��b�;�O1Wd���`�N$*'+PU�
*�(�)	V�3�$�!�!e�D�
�PL��9r$"-H)�ÔQPPz�+6W*͕Td�����kA$��U�A9ȫ���ԙvJ&e&\�Z�r�Q"�ND�Z�I%Q�i[T��В"�%$QK$�+����(�FT�"ds���YY�IiS8eHs2��ª��u�$���iT��:Rl̊�eU�)4T��]��zh����abdu�����0,馆er��\��L���z%U���;�&Z�Gj�jQJ��F�Vbj��QQ�˦����"�R#��Tt�I"֘KбJ��e�(��i�!��h�c�4�\IJ�"I"T4�P�"��VA�X�d�q �(��!�"4�%��Y.,����4�a%�kD�(�At��㬈���e�!:t������J�UVI&�J�&jV&��J����E2�0��5�-��~+���߾����6p�WP0�g:;�L+�ˋy�����S$t�/O9ak��Ɨ0N5�z�孭i�L�=z������9�~��B�7�����8Ң�S�5��GX�J;@��h���/P�Bܚ�7-��T��F\A��a�����2�)�w^���}�:��c���#8��}h��hN�;��{xWjj'�-�5|`s4l�3���������[;��j#ÿn��d��
Ўw�us�U�\�N�mk�d�6�#���}l)��$E�Dλ��|�d.Wr��u�s� F���t��UQ�-�_a&r:�G6u'}
��%�S;����yX?rē��C�~fi������\c����f���nٜg�ߠU��q���/����*��@��r���ڹ;mO��-�ư��L��ُ5���`h永NMKu6�X�y�P�b��m����}��{��& ]}��m����,��8mnM��=1�ק� ��]���+�	�����sz�����?��`�j�1ӓ�����Pr�ar�$�/Sq8#�8;���\>��g�s7(��1�g���;��vL��X��}�N\!�,��-�+�U4���*��O�{��<��f�q�1\^ׇ���j{���&+����on�ǫf�O7b����x������s��'�ǃ+���8wn�Υon帼Z������~v�Wz�����v�ð��ɜ�\�Lt��دn�=�!h,P9-��Є�|c(��-l��fB;Em7�{�a6�Kd��Y�,_捚s�s��z��s~� B�LZ�T�r"ȩ	��M��WV.腹X8��Vbզ�;�u���nSθ_���:v��򜀯�r���~	�Y�M,�[�n��{�RFg]�7:%��А��,S6��7m��C��F8B�7D�vUl���5��l��Y���n9Ŝ��8�m
r��M5<�;�����݆�2�uW�m#�]}8o��Y�W�rz�W��°��@g�Ey�Ci�)�
i;:�N�[%=�WgSF�ݾ��U�m�;p�1���h=�V}���U�?K�`o��#_L)�
xlQ^�}��g��~��!V���|ʌw掾����nQ@r�r$q�y�\-N1�
���)��a��p�|�c(�0�09�ѝp��ߜqBq�}�u�)L�L01�%����Fq��}Yv�����\â��1�3K��3vL��J�w޴'�����m�A�{LG;åa�/�@q{��\�u�z��<gi�;�Բ��5���S%�%�}lm������$��K��/3��>=:��w�T�ژԋmrz��
��Yh�f�½3�f�d]�&s��ա׏/+CN���{�8�|���QS2�'C�EL��Y�Cn�AJƧ��zر�`�0����Θu���/�v��f�@��J�'�ܝ�S�5ј���~���9Vڒ+n��}_0���ط���>Kd�:zm��kއQ�Ep���i�݆���'Ȩ�捤� ����Ꟛ$/�P����i4�ϗ�����:���/=��>Miw�=���V����u��͆-���-�۔��n�tK��4���
��^�N�}�όe��E=�6n��)�(?A�|�~]s�1�5�۬���N��������2#zBg�.��9NԞ�ћ�ʹx���k���.]��cx=z�(\*�|�eԝS7oV@/l�y!jg+��|��ԏ-��y��h��E�ݎo`����Ԯ��Wh��P� �G`�:�
��݆u]6��P������F<
�����.�Φ��ZJ�)�OGF߻���+���|�� &{]|��@yB����[�g�����
�:2���6��z�i�&)�9J#q���a�C�����ɼ������^��i��\�+֡�ʦ�L�Ɲ���]h���u1��nl�`d ��`�v�m���R��S��)��dtU�wr��aȐ�Y�����
����7����aW1���[�P�*���:��6:���r"��j`�ڶs����������������0��t��z������&[�J[��^��ۭei΃��2WRS��q����͐�qgg�Σs�r�tȝcy�wQӕ����z���f�T`�.~��� �������5�i�L����H��呆��Y���~�9tw,��*ᣙŮ�f�xc9��)��v���xN;�t�zhS=��tva��'aN���z/8�Ñ��s?F<<�t�
�5��9�Iɘ;��!j#���	li�aߺ�k����}�������V��
d?�/�^fޣ:{_���M�9؈|�j��d������l��l��/�h����rL�6�>K<�����{������b�t��}���hz��]V�N�7z�Bjw��q���W<�#��4�6/�%��ܴ񋈃�-��-ŧ'0C��`\^iBZ�;���1:p٠�tA�^n=.���y��gU��w]c��X�Ó���z�=O�"g�K>�ɋ��ON�Gh�{[��F�w�A����3ϧf�VGX���ͨѸ�2�v�噜�B�Ulq=RQ�����1r5�ҡ��`�{[,-��:�=z
���
��7U�~�sZj�QHT왼[� �����p��/M9D �ȗ�Y�=kz�)��*-�E?qE��i���|h۱B�6L�����oP�%[*OU�#˦}q����jA\[��g�%�u��N��t��@��I���l�=����
�:���ȩ����ԫ���l}�pds�T�����f��{!/A���^$;NȮ����"S����8 �lÇpS�o��f��0Js�Ho�ʄ-�� yD��M�=X�鈲)�C�T�0��{:i�)O#��:��;��ȷ-+Vf�����h�Bۧ$�[h�W�� ɟn�l�
�LG9B@.�s��7�����3;n;�d��h��[�v�@���<�mӔ��DX
�Ի�Q^��>Ѫ�6c���5��8
ܫ�R��LrЬL�|�����(���ت#�P[�-�
���!S\˹<�jt��k�[f<Sfh�w����+6)��k��&�CS��/�Gh��Ѵ��U�^��Cn����u�:�*�Y$�cs�Z���=
�g8����dy�ߜq�d TFp�-���q�NT8����d��y���=�̇�l����fb�h��F!՛!��6gL<�=:��u�1��1�����QW�o�ܞm��-�}l)MWH@F�"g^�-�yh�\2����ͽ�[N늊�j�<wL�Tj;:�+���GZ/��_)�yM�EB�q�bI���0�>��)g�^�{�|������< dL2��8/T;��K���|�ޗ�U�r<�+��\�~a9��2�L2������;O{�T�Iv�Lk��v�r*ѹ�g��M�]��cu�>�-�3K&f�g����%�o�U��~���ss�n�@n����Y9m�)�z���.�EZ;�ԝ(��tgUM�>��L�����Yu�.�0��lF��^f�:���=�X���0�z#�5^�N�m�g�������o����b��V��3n/*l]��3I�\��?\�`צiQ�e6G;�l�|0��Q=[��z'��m�/Q�b��x�yjr�֙���E����O�B$~*���pV�iLe/pr�(����L��egDe]*�,j]�j�fF�8���&�^��E>�7Q��\`o�[0StJ����"�C��ws��.�VZ��L�(�
�͇��ޘ>VR�O3GM?`�cƓ�oeC�� A@�8BU;���U���#���U�}R���Q�c:�{�%��.IO:�mepYӴ^��� +��L�S���T�VW���Y'��ՙ�[4o�&�L��B8ugM<ڄ�=,S6۹Svߺ'�qNִd8V�^�S�tt��N�Ww�V�N��6K��8��ji�G�^\��MO-�ʎ�F�2�z˪�7�h���/3ה�y��0J0fo�ɡܫ]�v�y�S8(m5�?!L�vu��t��S� ���On\�`j�)��twV=sB=[M�8SZ�g�V%ܼ������=/��o��j�U���]��}M��;��qb��UaOVNlQ�b�֌��)C��@5={'^_J-!�
7W��uÐ+Y��B:�ゼ:�We�Lw�ӭ�,�iHu�~o���@ݜY��[�n�z�Q�ap��o{ӋWh�c�w�"����w�æ�+t�7}x1��S.��q��ўhS!E7(�9l�r�C�\-N1���C)�#-����Mw0��vI���\"���'��y�)�醨3!�tE9�~2�)�n`��h�׫����W��U��g8e�93[v;��Et��Z��`P{f�6��@�nv���b=>�y7S��n��u�ј1��'�i�;�&��oL�i�M=��q������e�b��X�c����SD]f��': q��m��}6�z��g�ls���:z�즫ޗQj+�nwvm��Wm�&٦ˊ��I�Mx9���{n영>[r7	��ɧR�v}Mz�[0���|��UZ�߂���U7x�9�sbz��m�6-
t����	���@���O�Q,^���+�e�Wj�#���N���'N���9��<��ۺ���5���T`���9��)i����݁hͤ��aa�p�1ɞ�s2�;�oF�z�NP
c��Yu']�D-ג6�q���w�ѯ�ݏh��݅Os^�w;����39P�b�O^�,�jWt�R��3(�"��;!- i�=fe���Z��0o�uFTt����G����!�͸h���HW���1i����7��VS�Kp\�ԗ�dU�Xҫ]��X�L�i����G�,X�� ����5-^�H��\oz��|+��NaŐ*7��m�*�����&G�.�;��Իpf�oC|�[�Ʀ<ƚ��WS�����|�E�
���EE��99���i*h���ѽ�[�%L*�+:e�V�!"A����.Aܡ :�D�y��< �cLAs��4�"^�����v�D���+-C��R����녃��%�wWSu����5�vr��%�<�q�zLAu�٪��'�ss"Z7gv�>��q�?��3�C�
�b�|���L��#���;�QW0�O��g�{��92wp�cM�,vq-�+2g7qV��uF�����v"���WwT>�uMp��)��*��0r�Z�z�s��o�(^OU��:"����F*��s'�W�Gh /�E�N���(%�?:|@W��믜��>}�M�W{���3����'P\76�93�WHA����[S�.��s��Ҭ�5<,;�.���3!ɶ%��-�s�_a�>տ<����\�$��Ît��t�om����mӂ��%�[��@�������)�>��C�~���Mxa�FJj94ّ�bvޖ��դ��!�keȊ��~���wD��'�j�3�-�-��"���i����\t'�U��a�{���aIĪw����S(e)�����ds��EҜ��E优z��}�=����Y������aw'g��'hFOwG�K�jno�6��K�7���:t�Z���=�|E�E�KD�G�~��^���i��'_sp��̊9Bb�wM!�����	�w���<�m��V�M�u�|��E��n�K(�ל�:��v�y�|��M� �)�s<z�e�����zs�tG>i��>ϖO`׾�ڍ�J�c=93k6�v	5|��ǘ'���6w�[L%��Pg���p�U<��˪ܼ�,���+�&�C�^g3;�0s� �ox�"P��Ȓ)�C�i�%��b�w�Zަ��(���oj����{�]nj2�����vT�Q-hW�'��b,���w*�a˚fΚ}$.l����v���:���4�'�:.��r�� T�Y3��T�m"���g�k�m蹬���Eʧ��/�f[
`��O�.K����.�TW�a;�6�T�3cm��tE��\:9�F����9��L��f��tb00u7b�|��8�)0}
�"�.糶+E�v��+��?l�ˋΆ�q�b�_��>'�[%�Svu4muUp�!�y�tÛ�m2��;�`3W�E��M5�w,��R�x�������_^�v�A|6+�1���r�7=s{�8iT,Q���/vZV���[� �C(��`�/d�I���p�Ն���	:�p��ö�Jz�:�l��Yy9��>۹�.wr����WA|S[s(>j�nfq� 	*3m�W&w�!ݦm�9�u�qD۽�D�ق�5��Df�M��L�
��)��L
��v|X���/B������2<7~P�ū��u�Se��^��8I��@.m��[p��y�j�E4�8��D΋>�KW�;yX��K��xL��:��MX`oc�v�����F�U��:��K�q|�y�7�	q�5�"_z�6s���i�x��ދ��ū8�c�dL6ߵL�P����q��R�M�/�������r8&����ެ����9�s0�a�s�98�S�`���Բ�a�׼Өb��-��߾��O�c���1�����#^6i��_D���um1�5�y����i�х�¼OV���6)�79�IB�霯��������yV��,����%�?�XXV����ڼ�y�D�y��ݧ�L(�zJwi��9�3��w��u�9
}�7Q�а&���*�i�&H���k�<�� �Z�rΪ��Q��&�;�u�h��<G�c4���sKu�  �����:�H������R�rrZ��&�Ԏ؍sY��}	�d��p�4q��ct���S���S�yL�x��g�1z_�[Y���;�v�Ǡ���ۮi�l�_C]z��欖�.�7����U맰�t
����-��<��҃���{!	bޝ��3΋�-�\3V������o^�W7������h�4< ����!��ڻ�:\
���i�A�Z*2�Ivl����tYz���֝FV!ܳ�
|Y��JDޱ;w\#��o8�6�HC��e���A�xWA���0WR�w;Ŗ�������Ƞ��h:�b�]��!Pf�
���n4Ո�7��V;�O�\
����7��'4<!-��l����i���Kɘ���NqH4<��E94W�v���;'����_��7_w:�s-nj����h�u6��\}���;��vW�_��Τ��7�i�t:Qu6/��	ӟ_':����c���Z������7�ۏ�a3�j��*��υ��M��sq�ؖ��v�S�1���+�T�g��nOxi5�g!&��SiY��������H��P�˙��r�=W��ir̳��y�f��ӓ�x�X8j=�s.ݚIT����Os�-X�+5s��9��).`f����+B��iݕ�m�g��&��뱩�/f.���V�Ox��ק#I��n^��HE7�|�p*L5�9�9'[��6�[(�M�A3:[80&߷�.�;��C� �&�9�-�)�`ٻN�<��
j�I��+�Eh���Nm����%�:�耇�	�;wȍttwٸ�"�]-]��$ᘷs�âXH��}c�MYݜ���]��_-�{�sQ��v�|�����v+0m��U*h�9"w�× �C五%���¹��Ru:y�}���W4�Ծ�h�k��7��:Y���݄�+��W�Xś��A\�l�&�C�AC�����e�`\��#���I9ic@pz:���Z�u�̮E�5Ǫej7ӻ�b�@��#��p��� �Z���[y��Μxv6��p
��'�S�Lt_-��R���;�P�E�c��ʴ�7��5y{�N�\�d0�k)溍��]ٓ�5�%���fuel��q>��X�d	��˼lBCzl:��h9ouR��K�[�v����7�"�i]0�֙;�:d>!��\�;��(�����c8qN�j��t2��6+D��jY��7 Qu��s���*㣵iә-h�Y7�.2l�v���<�(�H\؟�w�X��ޢR^���k7ա6�J��q�m�����#ؼ��Zs:��=\��k���I�ăqU�f� ��m%H-�8���ooH��\�*�q�=���n�,P
�^3m���g* JW.y��Nʛ5��zOWh��t7�@���K�	����1�I�*��SoP����CRT�V�f�o:�� �ܮ�zr�uم�w/qg��y�_J}=�iF���E�Й%�X��G��g�R��g.>;�_iB�n�";'c{�:R�Z˼0( G9A��:��N-~ޏǿ������\�5�D�PE��Gdh�H�UWejUE��B"���p�2���rH������%2��yU�5����UuB�ŖpJ�ST �U�ՕrL���N&̬TBAI�Թ)��0̨(��u/,�
�PJ�JIg4��b��G,D����S(��F�fg��-H9&�22�Y$QG"	2�(�"�G�"EI,�VbH�UQy$F��$�DAg�U�U�C�"L".Z!Ȣ*���h	U\���
A8�r"*"��V�s"9We�P� ��\��DUUb�&DNBÜ'! ��֒�c�",P��Q˄�Q*�DWn�dQ�)·+�Qʭ�r.G*"��r�.W�7Z�Y'J����Qz'(���~������=�b�\�tw��#c�)�ucc�lVE|����uI���ذe[�Gf�N��A��pX͡�@컾��sl�ٟ��i��������A
�:i�BB�)�ܥ�8E���E�AKj�A�(�c��Rq�a���bq�[��q^q����1�[P�*���w*:1�:�4gLl�0�H�sU5��H���fΤ}�p��8��w���|�I�נ�u�p�9wκ��(-��;�n����u4h���M��#�z�;?*���=G�V���.3Ё�VSE���/��Y�o�����k��Ӯ㫩��Q\���-�!ȑ�a��h��ʘ�Z�a��K�b/����͙=IS��	���-ߺ��%3]0��2��sQ9��"���T�Ξh��B����Rrf��� W��w�O�dXynSo�5�hC�z�<�ʇa9Nt�dM��K�9�����u�	ɩe[�0�4tfJ9�m1�����I����F��&g��~�똁-��97�#y��o�ң8m�c��nǅ���d�$��.�|�}k�t�(�ة�E7u�[��r{����&��]��ׯ����dw��ө���ð��=g`�	7!Dt1(�Ï�1����/�F�Ob�+��̂n�W`.�T̜jp�{+Z��:�bu�ۭqA=C9$ۥl���<W�A�=q���I�o���3p�qZWO�K�5"F���nVN�avּ��u�Η�OVKN�:r�Rq޵;�.|��r��`�}yu{_y�JM�:8_�K�o҇�'�
��,����jw�����FS�(���S�n��OE>�۬���@����]����-;F��Ž&��GH�s��s9·{m��'(1�y̺������$ oC���Ҟ�{�$��ٟ`���n4�*��r�����K=�\!�.���S�B0�ҫu�A�|���x���"�2���p�u��"PǶ��/8����u5<�J�)d�tl��!t`�����t�11\�'n�h�w ����ơo��S4�=1.P֓�6_��ݓ+�呉����HCkݒ^0.����!h;9G�ɞF�w��cLAu���07=v�U�lA.h�F7��ryܘ��JC����=T�+�dtW��;�Qp�fe��Rw,�S�U��xp�a�J�s�u®����u��,�:q�wuC�3uMp�� O��R9C��V�D�#�ޤ��z�u�vZ%�"ʆ�q��^<2����b;@B��3�W����\!���F,�Q̞��v�R�:S�fn2(�ݭ�p���ggn�[nY'�����y���D��t��ή}嵎V�E3��&Nr���ǚ1���l�|(���c"<���0��3S�-�YӁǝ1�/��P�ל�g��B�a�N�Sl��\��c�/gE�3܉Ԉ���.�_�����k��[6�c�0wWPB�G3�H����v�"Q�v�fv�Fc��6�@u_{#�6G�(��G��[������ߞ��fa��U�ޓJ��/s�����Н�_
i�^��,�ܮ��+���Jb��{��i�eG���ڞ!vr~�9jk&���6h����Mg��E�����wD��{��1q�S��MѻM�99�sK��.謝FI�ɫ��OU�Gh\''g���v
�=.����3���i������r`�n����*�>M����m�ɳ���73��Gp)�s<z�e�y�"�>|~�/�Ο^�+� �/Jo� ����P�;$�&�W=g2�r���%C�t�KoN��PU.Щ�6|sy�%���6�������X�wn`�n���n���n(K�#%C��P��o��Y���ND�xXǞWc��:�Mb��捊r��!������n�@J%�
螬{i��)�T;����s(J l��٭��M����fN�Wd�rz��Ӓ_��.B� ��K&w�R״���{�KN����N
�#h�'c�Fqa^�.W|�Ό髂�vS���޳}����G���K�H�լ~���V�!�����B���r���S4s����3����q���͝uΡzlw�v�B�i��"��.V���;�H�X�x�����R"I$gk�	9���Z�l�e@��9�7NR~�m`*kR��G@N��Jƞ�=�Od�ٽ6���9�
����K߳ap:1�����C�zzi�)����a��223oS=�t7b�쳳��h�lSX��I����{��vt�g9����ƴ +:�";4K�GL��-���K��D<�Z�x����dy������Ϗ�����f�g��f���3b�mg�G_S@B:7�̇F�,���uK�l�٨�.K~-�`���1�N����`��G;�ZZ���(ߝ�������RM�=KW�et��>G�P� I�����s)n瞙�b`KV�N"�*�}�C�q|�ynO>H��~�)$��b�߸�	e[�/^�^�h�`�tt���95,���8+ת]�Z�wL��/���|\g C�l{i�1��hn�O�>v�a�Ԍp}��>@X���O�jYSh���{�:��)�x?}0��*�L���֌����R��ͽ�.���p�:�,k泥 ��Bw��d��)�1=[�.P������7�Z��h�Qo��}tM�f��K1�3�<���}�2�j�]4�!�ty!�4k�y�gf9Y82�k:�7�pϬ^���Pr��dڊ*N̩��� .�}����a�/, �{��^�/1��os�i�A�TqRov%�t����Ȱ�:у�n:X�ڷ�99���ڪܽv�U��wd���D��BI�b0c4���S�5��̹�!*�tk�{��Zr�O3���f��t[���Qnk�=<7�X�U��l~ʓM.T�n�rx�}���>��sٳ�� _ی�>+i�D �_�f��I�{*�u� !^S�R�9�{m��;�"�s��::F3�l��9��kP��d��p��2�,n����� +������H��Utk;��'~ni��"�5zg��*ΚykP���X�8or��]�u*`���5j�lȾ���9��y�%;�h�N)�,����z/�)ʩ4��ܤ�(���Ղ#��Q�"�jf3wI|M��U�~�r8U��r��]�-�`��g��~B�����D��u���UU����[�f�+@���h�M=J�;����������`>�h?G�/�z��v�XL�N񣙻��t)�=�5�
n�w���h�4)����P��D9Ìé��^��"��۬�6oNX�b;�-��wْ�ѮBq��'�w����y'�g��?��\g�]2�^J���I{�K�.�(���#����l--�6ƶdː�#Htͬ��
�`�5�R��z)P�6��'���Ou��q�;�a�Րh��d��9�)�Cz���b�+�2��Le%�'�;���KOWn�V���YW��˫�p��Χ\����>�£([XX'9ᔳ��;��WK��x�~0(9%���e$ ^^wI����H�m�D�t<��Oz��ֻu��hӫ����s8���0����$�#1�犑��[�� %P�����<!�3[c�'&i�׶;)�ymdNN���|M\��Gb�B6ۺ�tW+ʷ�91}�rp���m99��F8̄���1�� *,fugY�:]�p�(�oD�A�l����������UǦR:K�GJ{�m��]�F��ߺ|�/�� *����S�Z2�8_u�h8Ǧ��v�d*0|�t�`��)�DMʋ�jI5i4�D`搙�����;��o��)�Ls�o�Ru]�Y ����ϋ�t��I��P�8!��3���&y� ���ьx�u�K<5�\!��\.:�?�&L(��-��P1=�9�E��Hp��u�"PǶi������rk:��m%M���#e=4%���}q��,s��p��m!
� ��N��#PǿLB� =�SNPy�(G�v�2\�~�l���\{ܾ=�t�/��n's��8V�����<v�
��g���\pξ��T��
���{㶠v��-�����=�֐�\����8�����_p�>���};�YzB�p\+Ij�W����p�Ϡ��=��!�Zl�m��ob�i6���{:���vIx�K������!V��ʮ�d�,7�;��b1VٵT;��d�q� �r��=��L�|�ON;�Gh��=���0�2�1��GEZ�w*.��v�qOoM�f�Fr2�7Y�����9Ίk����ON� �qt[�f�����4Ц@O*^B�>a���/�
�fQ�,Ό�KDZ�h�q�b����Oh v��Q�+�8�]�R�jhʚa���Q����3�)�̇�~Bi�y���4b���.ٰ��۫�;���WB�|q5f7��N�[9=�[�{�+��PfC� ��G��������ߞ��tl���2svq��On�y�y7�������SN
n/��<���+��m��}~����Rc��}.�L���0^�~_��횞z���-ji�6/�%������G!N#`��v��C�6���λn�a|F�]�u�X�l�F�>��D���Ι�y�o��6���r`�6vk��;n��тx����tl��4��
i��^l�}�ʼ�w�ޞ��ϛ�4�>��>�w�ؗ��U�����sI��h^��mf��fh9|�W:��� &�5�����5�ʸ����>K�_)�r�>��:��Gi]xaY��J�˾�����殣o�w;���wgٵ݉T�����9^��m����+G�q������m��2�ݎ����;s�G���P���1׏>�gE��r�	������
���pVؾ��Y�:v�x��:\ܪܽv��"�� ��N>W�%�r$����ȗ�X���5��nC��]���'m�&��8���X*������n�N�KZ�Տ Q*�T׳������h��e�#���{�i�ʞxY�ji�O�t\�z���t ��z��z�m�#o��ﾆg\����#���T�f��$/Yl����>&��O��# T֥�ʊl��0����t��N��e�3�np��2��f�[6�����޴��k#�n�[�w���&��������]DCέ�#��<��=୊��~�3�X,��l�s���{9O�8�d�n|m�ʪ���S!�W��u�@J��F���^2;|��~�;7t{p옐�9����L��0�9���Y�WK@B:����7	w!����/B������P���2泺�_����[!�hSc��_[
򚮑M$ �|`�a�my4�W��d���WES�_�s���>~�ĥo5Pd��]�[��K�zGv4�`,�_�Y�uGΰf�@S=d�+��ͣ��ح�j���f�ŗG��}�%�s���G�c}�d!θ��q\�ަ�w|�tY�����Ź��|n����>��Rs��|�m�4*��,�Nu�z�ؘս<�)��w���D�Sq|�~Q]�
)��ѵp��:"��z�Z��gS��'0W�B��+�;�&��3oL�P��Z�w�0��ޗ�W1fIü��U'����TILb{`C��\��l�i3��0���Բ�a�y�Lئy��]�,�B���Ƽ���t~��߻��[��d��� ����[���yL������>yA�+�sA��'"�-��j����<�si�CN�����ͼ���2m|�u^/��oҼy��d�|]��� Ѷ(�^���8ht8~f��L�
{:-�E�i��(�5�՗[(pl�Uf_���%�&���\�+l�ƨ���`�Od뻩l�w��3�e��~���K���sm�( �2��9�����EX�]RuSٮj�x*Bg<)�#��b�xkP���Sθ[G\{�h�o)�
���'�ݤ��F��l���3���M6@a�P�gM<ڄ�=3,S6۹Sv�P����JޣPa�"A�� ��SZ2utJw�)�>+�Ƙ�z%�ʃ-.s�Q�XcUYF[D+˪w���u���4�A@Do�lT�,s�,c�~ʊ��\�Q��x?7~;G��]"N�ҙ�+8����F>��[uy���D��|�K�����;0sΊvVY����jr��\���KI�y�1�i�'w��7j�3`�Ķ�����)q[�����G~}�E�uW����­4;�W]�և{apxE3���\S�i���Tm�󬓏	?�O��=�vt�`��T�^�*�;?*���ϣ�^�>��!~�����&��t�����:w����7wN�����f�2r r!�ض)����ξ��d�5������1���������l���'廮��yL�L4�ex�P��u�nz�@��n�����c([5��9�,93}���Et��x,�L
zȭ�n���>���8GyX��=�p�`�u~1�z��;Y�>a5��6���V���k�v�%�u�9Fo7�����*���t���71[��~6�F>��81�ᛱϙ.�Gk�\ĉ���Zt�y<�ke�E5�W�n�i�M����i�錅�!����m�h;�exW����¥�W��T짥8☙����1�)�}�ymw�sb7xC
����"�5ϩ=�Y��i�駻'��	���w�����=4O�-��s�1�5�۬��F���eW(�W�i�ۂ�rU�G�w��
[���AԩΘ��J�I9�.������6t�����"�Ńw���n �h�Ϯ�W���ރo����k�,Uߜ,pYx�;Ekx���g&�TV�B��|K �F�٫=��tӽϋc$6H�YR;�%)��˗v���p�8�V19Ht +k����'Y�d�C)��^���,���N���l]�[ܙ{f�<��{es�ir�x�������a,-oO�cK4��a�*����"�TU�jf�ήk;�pS�����dp�1`.��Lv�s����>k���i�0�g��:��!�X�p�3��c��x�k���A/
��g�Ö������!�)�^���w:K��l��L!��wNr���¯�c.������O�`�L`Nȁ1�c|mk;|XZϵ�|B��S{pl�}�9�^�Ѹ�zȷ��乤��ɓ}Y�oI�{\+
u�E���P�M��)5zxm[����&0�O�0֜� wM�h���о��Q3oE�h�=��t�Ν��7)��S-w��a�ˏq����9�]�l���qi�S�	�a<ԡ	��۾���"��b9�k�x;��4�V���ER%h:W��r��Dx���FZv^oË����Q�״#�v·�Ve��.�c�I�F#���\~�r�!�HF�@vȻI�Ώ1�;� ��1䝣3�SyP*}E�s5��L� �(<u�q�K�7n��ϼ{OI-9�j��W�=Pn���R����9'�
��}�YҶ����	���P���»�+�p`̾��q<���]�sR}���G+h���)MyW��b�(�E���k'O�����H�ޏ���F5u,Q�V�;|q�dΖ���t�
f(8�K�n�=@s#�3�<��S]�WL�g;�S�1nP=xk��� &tk���:�r4�:�Y[ �7-���[���j�����_��,+t$X��YE�b�tm.h�A�(kml!e�#��a���&��2���+'��&W_MgY�3g:�kJ�8W��]��x�Hd��I�z�ɸ���o��r�_v�c=��ni�ca�]����9l!�N�S��y�*6B�M�k��^荾˼ew�ׅ�^/{�����f�EOp3�y|ѡ0��zM�Ş���yw%eB�h��LhtQ"a@_t�{�t�@3�ep�K2�l��T����/'(T��3V�.6���6Z�� �ŵ���so+&��	�$��]���p��'�^Pf��u!�zQ����c�{I�r��fذ��m}��w���IH���*�^��|��ݸ��跏��������s�	�Z�8�7��d��[ZC�&v�C�L��-u�(�|=���x�eb&R�`8)�"`���Ѷg���;<��T��T�j��:B�r����BL��U�w�K���c�存w��������"*�8\���Y�˧J�����C5�E�����Uh%@p��
��i�p�W=T�(�u�H����s�;���r�Y��Ǖ��|��E\(�"�/;��Q$�"*�y�H�
ySdA��>G�B)�J�J��ְ��J9�AS:@r�9ώ���Q˔|�\*��2S9G
�U���Օ���T��J�-"��QQDgS
�B ����EADY��r��s�i�F���2��UDGU�Q�UUQ�q�]��ds�Pz!p.�DTQ��N!A\��(�̮�
$Q�
��Au���"*�UwC@��������Ԋ>[�Ȫ���kH��GUU�#���

�p��2��
������
���QQ)�B�� ��(��EE�+� (hW�C��{�]w뭬ھi�^g�OL�Pm�/��CL�W�oWY�����o���Ƌ�w���C�v6u��d��|��wf�o��S�����M#���l�gإ�7�x=z�(\*�|�]I��a6�bT[}�X����9ss�GG^#}�z6��߆�SK:�C��x�,��jWt�&�Y� �2'*�ۮ�L�K���S2����Z��!��D����@�\>�l�5�_$3��.?���;��~����-�.Tݷ�8Cv�@C[��D�ym�c�LB� =sr�4�9N�1FJ/���4�S�<F��.�/)uu7^���5�vr��%�;�w��6B��鱕��6n��l�w��D�~�_��ǖa�{Fc%!�v)��i��M�2:+֡�ʁ4��������k��{Gc���C�l�Ϟ���g����SON� �q�:q�{��zbxN�<����2�؆��$�3K O�ԍ1~ȇs,�e�[�;�U��)l��b;@B�Fp
�;9�Cvj�����F�'}1HC��9�̇�m�i�?Axq���k��s`:��0-��v&�xe���E�D�D�C�!3�熶�wH��ʣ�d��l�צf���nφ|>�
����u�Z�>���v���5���[�Mi?~��9�8�V�\2
�A��-��)�Z�M_S�t�e��
�u���a�	��ߊ�E�=�l�y�۵FK
t6Xw5�0�y� I���&{m���Y��ⳑ�����Fho��Ob��5GV�dŸ��8dq|u��Ժ_�)��w޴)�7�g�S/ܮC�"__�6s��Vs��T��{2�V^f����O><�&��oDঽ�t"�ji�6-��_y=�Nq����(�a'�fN��!3��_<}���I��}H~`1�1߂j/=3��LOK��gL���Ϋ}��ǽ��O�Q��o;��N�Kڊ񜑃�ѳ�573��������*��;�A�����Zp�0�/����5=O��X.���Q���y����ǦiP�b�w����[zup�y���ϯH��ֺ�;�pvX�ڒ���V��VTj� G�[�7�%��ҡ�5�/Ų�H�؞��W�ny��,��iSǢ�E?q��Hjn�ڂ/�p�
�KZ��ǀ(��xط��5ɷTs��R��<�g��;��͟M<��R�)d�rz���9%��E�C� *%�<\RTlZu,���ݳo{<�6�zb9�	 ��寡!�a@�	�L���e'�q`,��*��|�m����e�sGV� �/�Z�s�Xz��D�[UAuM&i�6�<�]��7?w���a�AI��l�t@s�E�td���=!/z�� �t����f_�-w4xw�3�ǤH��VX�;�4��Yx���d
����GN��zMYCO�F��%��������A'��j����K�ID���5���-�DK�b�ȵ����eB��f�����^�2Evh\�"�h�k-B�\˹�[,���CE8+b��)����gWc.�*����sk1��d�[�+� ���Ѽ�������H�xX�B���p*q����4'�E�msēgL��OcrA��wu6��G_SEzO@�4���	w.�bPZ'�������@�՝Oچw�$>�gD9*0\s�.d)��~�?J����<P�BR�-�j����F�Υ��?z.9��c�s�S׎���Q�#R�w�քK��g��0���a�-�#��S�Q����g0C�����dL2�ޙ�z�ߠZ�wM�R�n[0�Of{���Mgq1\�/�� C�+���:�rg*a`)�.�^ߠ?�����O�\��"/PReF�u��;�uK��E|)�W��p7�:�m1�5�v�vK'��#X�xSY]s�����O;�9�mi��<4�oU�zn�ʷ�읁��V�H���=*9���:���毑��~f�����g��+:-�E�i�B�Kv��"�\`x*�;_'��3�Hh|_ǉ/vtL~�\ ��� ��۸u��4&�nL����Β�*�oQ��
ꕼ�����=��	��~;E��+��qZ���tv�Xu��������.S4�(>�nm�jRԯ�_Hjޮ�1��r�2*�c�q-�l]��M�N����'���gK�{To��(�K���<i=7oeC�n�@�[���5lW'���9�������蜦ˑ��#��
l��5�]��$"�)�\.8�೧h�Ǎ*�C+��.sy3�`Q�� n�N��5Se�E�h����!gD�Z��=3,S6v�~6�5��K&�b��Q#9��(�#��"�!V��
�%;�1�}�����a����V�#	�g��(���'m�V!����M�g�v=@�4;�b�:�����pP�<z��9�0H�s[ƌqy�������d��Ζ�=J�;�֡��U�w.�a���1lɧj�A@���8sY��b���w�';g^�S�p�|���������Q\���*�뿱u�����#����E�f�1pxC>9�x��2:1=:�Z��:ِ�w�������=�Z�=��_�|�/���\�س��-��2�:���xdr"��� Q].��Oz��3p��1��
#ܬDLh�"���yM:�X���[dԲ�ޙ�ܲZ��ڨ��|�C���L�읹HZ���m�^ �e1�D7ܯ�+�}H`����]�HJƞ��B��9�6�]���)k��goF3};�i�7���(k7#�͕ � J��ϗ�(�c��6��S)=_y	�
Fz�����˰�y���'����U�,�9��_)�����nb*��Е�}�Wiмw�/��|
pZ�<n�>En�Y�����SU��芵�6ۺ�tW�^U�����r{���i�������­�����g���6�~y�������oE�oD�A�΋}���k�S����tp�ҮG/>��E#������?��ޛ���ܞwxk�z1��	��\������v�d�i�����n#�b��yL�
螦�������l	��b��O���ür���6u��V�o����OBI�WC�ܛ�]U�#y��>Sp�O�鈳:1��xlR�֥p��|n�X���=�ѭ���U`�ѵ%���#�u�@��yD۪m(c��/��1�EЇ%��nj�vo�8��o͏ݙ���[�Svߺ'n�!��YD�ym�c��,o���v��vFr$gk�uM>覞�|��,��M�%�2��n�h�SZ�g*�%�?]��nCʎg����M^�����.���ڨ�U&q�Tv��%!�3v)�ʞ�O�2: ������L���V��^�1�w��S�K}b�9b��]@Mq��i��w ˩�X[T=�b��~������ن�4v�=��n�}$D����Ҧ=y.���׍���!�"Ն�f��}��&]��WK�]>��.Q���V�LN�ɶ�b��2{������F�T�<��N�#GF`,�,B㻦t>X�/,@��Z�\t,�d����l��[?yeV�W�R�K=+�q�kǆS����#�Ō��W@���
�N� �h�w���P�z3.l�w�1҇˂�����^��؈�]���{�uT[�0���u�������*�]m:��g�c�\�pȧ�F)���FS��$rzT�q���9<��Ϳ?lD>V�uL�s���M8.�ᮃ��i���� P��3'ѿ��k���%�Q�قp,�l���MJzm��{��E5���ؾ����MU�r"#/w���bqNyf��3]N!G(ݦ뜜����N�z������Ι����M��[�͔��}�u���O��X{�!�x�-%�~�
�z����W���A޽�8L ��>
�q�l��;A[��z��7�f�k�^L`��L���d��5��~C�WZ|z:)^��,��k�n�'��E~�����|�e�n_�\�\`ߺ'+�"P��Ȓ*T:3SZ�n�̛+���HS�w =�Ej|���޳�<=�K��I�SN�nߍz�c���K�`�R�Y����Iy�A�.��|�t���C#�â���!d�bL��el��>��:���xev.4��do
�uH���d����l���O5[�c�����i�Yy�{�S;�z��4T�EE~�V����ڂ:� $!���޴�qWBu���a�`�f��GNC�md���t��ZR�)�d�c�?�q���.B�� �n!ɖ²��S�d��S�k�3��-p�,sLG9�mQ�a�y���_�ʁ�-�L����u/�MNjSӃfea ��%�@�����5{J��2�U�3O>ͅ��DY��l(h4�=-��ɑ��K҇]=5�_�E��i���c`s���wʕ�=�1�ҟ\���z��W�C�t���:����;z�M��ѵ��S!
������8Z!����y� C`UD<FP�U���A�\k������Fp����M}M
'�SA���r�Ìûۄ�)��Z�3{c���7�,r�=�C�ٲ��1L<�=:�!�hSc��u���SU�)�ā�^ctq���&�"E��a9�n2y?xvL<�2
Wr��g\�:"V����(D�W�g�'�;�d<B���wgzy?�K��`��LN�1����~f�J�95,�zg�~�mt��v�r�Ww	{R5����{�����_"�߾�A��m����C� Fk$,�V��=F����\�<C�G�B����i��Y:�6����V�H+���}c
mP8;�oo��i���|3F.��`ɸ��3�Z۽{�ı,�o���5��0c5�����̔�
�����\�߈�_���ϑ���c߂��W��=���W4�fV��1�޲MT�+��<�m��_i��o����& ]}��o�οA�0O���֯.�7�TC��u���-Xhi~f�9L+�V�މ�7�ܻ�����-#w*�B/�pV�+~�Xi�Cmh�7��0��\Oy��5��>ժ���}�-�Lg�E��՗[2���D�`u��Zu�oD�؉W3��H�������o���� �[��S�$B>�4��sǍ'��ʇ-zEl6J�M�sy|�}��߼I���M���Z��(s9B���0��jIO:�mepM��x�Mh]��m]r�ؐ17���vr�u�pQ	�<�5Se��Y���(kP�gM��<���o���R��%-�l�f�{��;�q���
��!¦��-�e8���� ���NU�1h���֊�ǻ3�Y��M�l~�;KF7:�݆�2����u���­4;�W]�-��.����b�<#�F��C�:c��B_0B���ӯ��OhݝM#�KGp��Z�g�Mb]�Ǚ�q�2\&������+ܦ��¬��J��˨��cŸ�ø�߮�������U;ԕ�'���$:�a�N�罰��}]J�辛��`�MYm���>���1�{�W,)��cb��}m�}:������{�{łs���͊ᝦ�~w��B")�9ۇ|��:��T���1�
���z�u��Tf�R�8�K<�!��x��
���C�\'�-�
�ǆS�=|ON�V���Bq߯WK����٭�Fb���t�t�T��-DS�g�- g�a`��xe7F�\<��^pQW��kT��{�㼷t��}��mu���
G�ӣ)��ޯh���B{��s	��e}�sM:�ޥ�;�������0,;���<�C�w�Ɗ�:-�o�}����k{Ϭ�>�L�x�l��OJ;)�ת]DU����M:+��[��ڐ�i���扼�p �y�SQ��	��#�Tc������;<��aN8�&{z/z%�_�:-����-�۔��nѶ}-#�d��n�,Jt��;���Ss8*B�6O;���>�A��|�~��C��>�T�gz�G�)���/��?j7���~oT��g*��:���أPpa���R ������q�[��g��FK��oV@/up�3<�\&S��K9R��4��]o�=}�+iQ�|�)��]m^�Rn~���K�[�3)#z����i�fUk��)��7{"� ������y�C��Jx쑺UL�A y�d9�����Z6>�W���Zx1�z�s/��*�s�1Sc6��X�ww��X�:�s��S�4կB��/��N��t!�������O�D����P"�m�y�D����L��0���=^(]sY:���=�MO,�WSB�����,��t��ͣ$!�'�'� 3�9�%I�M6�W&7��T:b5�]M?!M&)峔�7��{ �X�]]Mע�!^��T�f?<�հ3�;���p�s&~a�i��m��s�U�c��=�1)�+�ئ*z�<Qv��t:}�{Q1��'�(�r�w)b#�����/|U��xzgG�S��l���Qӎ&�g��b�b17������S\&�:dt��D;�F ����ݰ�O�'���\L	����,�ZL�M��lF<[�tWu
g�T���p�s^~������e�;����y���5Ǭ����"s$��g�>d%���Pw�Q�A���C���n�\�iˑQb�e��}�]p�%��ܽ����/�	w�O-�g�r����?����;������-��Y��ȸ��>��ʏ�ֻ~�|����*����,f�}�O�վ����7�� M�b7����_�P�ǵU����.�t�q�B.8텡ھ�n�7pL5���u>X��I��<�ū��-��m-L3u>y�p<�=ٛ�+�w�W����1������|,k������Q�ۭ:s��I�V4�IΨ����,��7���y_�*wVfkO[a`�����Mt��v=�V�i�&��-���V�Zf9�bT��9�"ضC�*���B�^y|�ٝ��4���AtM��Wh2ه�.��l xe����גL�n��km��/wnv��9��q�t{����1ml�WJ��c�=�H�q�%x�~�[�B7p�7���ep���Ex�Ul*� \M�ÌN�m^X��k�Q�P�,�v�0���o A���MY�d6���ܗ�lr��	�N�KK���y��vΌ�/�r��ܟ]i�b(+ʛfT�}�,��Z>O���aw-��u�-���3�)݈7<��:w��t��2n����8E^��G�����8$�kGQ��ec&Vs��#f��C�A#u����U�����i*\�	�{���l�r��x ]����5��-ӹ��l�Ҕ�.�--�I����D����Y��r�z�T�STW��#<��Bz
�n=7��#���s�,i�s,IxD��w]�*�}ҥ��(��t�y�Й̎]��A���_Nr�ҳ��)u��[��I�2��C�F.��E u
�8�Gón!]O��&B֎!�.VɌ�;�x�k7'����@0�J���uX���uh�uV>=c�_u��.t����t��"��3;�[ɩt����t����u���{�N+d�m
���)�wJܱ�ƞ����:"L���,Q��k^�ol�ݼa�E���@��z�a�|=n�N�.����Ő#�;�m��Ҋ�B�4�Lʇ^3w����_S�\:�у#�B�ᶹ���+�%ހ���"�� �����ɜ�*7S+�k� �����ܴ`feJ��`�6�����;
Z5�.����{Q��ZfFQD�O����_6{���#lJ�����-'sI=�W'�Q�{�᝔�@�t̸l����6K���9�q�>#s7@���β{�u�KdY@�h��W,'�����Fe��(*D3��j��3��7�n�
����V�V�1�Y�1s�c`��Z���bC�ih^�u����%`�E�7L��\zr����z�4�M�/�%����{����_�S��(^���W��	�;�Kw��x�	C��b�*���}�O�M%�u��Mї�������3D��h��+wv�fi���6���E���*��Fվ�5J�5m��|Ў_:��ST{뉣믞�3�K���GC��A��o�O��  ��&��;۴���*�I:�i諷+����oouq�*�C
��U���jN�0�.7��]���y���l���O` ;��,��U�UQʯ&,�<��r���!p���(�P"�Q��&p�����XDW�p*��Dr("�#��B�PEs�����8UAr �6y���"�AW(���z�E�i�.�D���"PC�.U��UQY���r�G((.wV��Ĩ(5�DTe�(9rQt"��J9S"e�QDr�EDU|�\��y�UÅr"�9��;�TDR�*�̥Gu�Ȋ�$G"���(��Ј���	��A�G#���5ar�"(��>=ЎR�"UTQ�K�2��Ȃ�wD�)�"T\=S
#�C�r#�WL"�̊�"�9^I��_p�a�s�Q�.s��"-�p�r��B�"�� �Xq���/0S:��y݇mp�2�p��S�}�J�D\{��[��달$�]�	v3y�5�� ��S͇5��Rc{D�9�\��$��Y���L���c��c߂����Dv
bz]���L���67���E���D������rWX�~�90e�r�כ�����	��a�1�;ĤgRa�k� ��[��LT�ͦe>�ޫs]�x5��ٵ7�C��2^`\|��~1^���E�u��6�g=Aβj0���R��=��/^�YPB�`"z'9�!/��$gA|E9z��;�O����y��������z� �*�E?qu8C��"�� (����
P�MGZ�:i�⧀*�J�u�˝fΚy��<S,�C�3OR~B�rK��@@ig���^g:�+�t����b[�i�����b9�Q�a�yk�He���_i�}������ڦ�D�L��H57��q`kR�磠'|Ѫ�S3�,"\-�������\�w�8K���S�"��+�5\,���=4���ㅦB>��r�a����CE3��)��?s���c#�^L�[�f�'�|�����{���i���,Z�g���R�`@v�>�K<�Y;�g�*��:��ċ|�|C{�mͅg0{���(��GF������֦�+�tܭ�J;��T��#��Z��)�m��||������|��'Z�i|u�����dVԦy�5���h��;;m�u�s��
�Χ}S��1�Vf>ClQ����3��t�s���|ݒ�F����� /���lg�G_SEB��d:<��_2ݎX��o_P0R�:z����#�6C�ϳ:a����	8�|��Sc��_[
SU�ve�<{�<��D��/t���&x��ڐ��l.Wr��\��;Z�O8�J��G_��|����\`���K�gt�2j^���r���ǎX�:IW?o�&��1�	Ly��K*ޙ�W�]�ҹ��'Q����q��U/��_W����pA�5��������0S`\'&���Vj�L�ci�:��2�n��:E�L�����}���������E/��-�x�7����p]f���P����':��vX�
�1*���oD�Ӎ�V�零��v�tKO�yh���4n����vv�F��GzLc���z��������΋���3ܢ��v��"�� ��O��1s6Eӯ=Y��ۧ�����^����ƨ�^�(�p���n4���Dc�^ T��O.@���>s+� B�bЮ�T�r"Ȧ�����i�K�Z��%����]te>f����9*�!V;E�]cZ�WJ�wp`Hf�FF��*e:j���+�H PB�G6
5)��vs�7Z���%��v�m��on;6gG��e�P�-tt�H�����c~��pBVѼ�f2N58��]�a�g����'+˒��N�忓�r_��� +�\� *S)�Y�j��i��M3�P�P�gM<�m9�t^OpQ���~���v`��\��m�'�mn�`8E�%;�h�N)�b�j��Ь�8|Ow15���/Wޜ���zN����݆�2����u���½i�ܪ�ėygC��V�7*�U&���ykiݳU�B;�4�b_�kI�צ`�u�Ҟ�)�:�4GJ���+֡��C:e�i��]؍��p�N��v˻�(F8��|B}����F�K�c���:�L���Ц�gum��Ց��k�(�q�H��f�<�\-^q��^8e��=X��p���~q��D`��]�*r�Fw[�lrw�*�SB�1@������D�g�ް�Kg<2�93��t����M���9�@@�g)w����E��So�)�Ԏ�U̫�;>�vԦ|���R�3٦sb.�{�M��3��4�
d��ƞ�{��#���m��?1���\a���sp�U��N���#�2"_�B�j·Q
�W������.���][�\���6[�Y�$.�&�ytr�e�u����^H�_g��s���|�;��>aq�u� ���s���lÍ���]�c1i��p�����s����A,[�8[PmEf���GP�F����u�.�&��9��LgUd��d��b��ss��O7�`�(߷���ϕ�?4���ю3!?>�d�!E�&;:;��/�b���^n��k�6��*c�����R�vs1�]����XX��;M1q1�w k%;���>�A����s�[p�͢�t�RI��S�#u��N�����9��)i�NL�	���	��U>S�,���/7w����9��o��·�&5�;�������$ m$��~	zޢw�g����)��shS���^D�G73��3�\�z�.���R��(�#�u�@�Z��R��U�(c���zLu셽oWq/]#cw��uBM{:��}|�4,���-ܩ�oçn�h�Wt R�N�Π>D{���S��\��;���
~i�8 s��4�"^�7<��M�%�2��nר�㡸�S.G��[�C٥VP��}g�ip�9v���C3��w�Dg��o�\�K�����
��-�RD�����鑰pr��C�>�����`��7��z���6O���������D>�I�/պr���b�B]}n�,�"|6�����V�:�I�ka���w��xe����X�=VTC��r�̖̯f���Ӫ�o���HL!�s���͆��r�
����v9aT��"�T���#�Gm�pB.]dl�>�{6OK��s��/mbp����{���G�B��/g.Lm�::�WL��/S�`�k�ZE�k�ps�ճC�����:e�P�dA��/�E�N;�t�zhS=�̇G�%�pׇ1�N
�����jzw��ƣw���ɷ�(�*��:�ɘ-��-Ds>��-�=�,;Ϲ\�
f�2�����6ƼL��C��ҕB&�����ҰU��|�gM�=1٘yf�R�IG;�_�����Y囕�@�����k/�fr������}~�F�`����e><�&�=6�N
��t"����l[wD���:�T��l�k�h��D�2����ӑ�S�1��7i��99��B�0W�.읔���'��x��b=��ּu=y��u�g{U[�w]c��2���!��773��B�0c�|���&�&9�U�9v�f#=�)�(;����]3ϧ7�}��ZӾ��#Wǟmc:��el��=V:��윩x��⯱ߚ�S�x3�K��*�|��O�}ڲ��B�D�D��p�B_�	��6�euOMg�t0��F��X}�ȗ�^Φw�Zަ��(��4(��8i��0A�\ M�yNv�^�ǉ�Ț���Ű���Z�&��b,�i�w=M�\׳��҄�'��=I����{��ۣ���To������s�4�p�:��!��H:u-�b�\�9�++Y
����\��gL�"�C.���`��=&X���{/�Õb�n��;jGr>���:N�k6܂U�k�0�j�h=ݘR;-�C�����U5{{Ů��=�p[�|�Aw����#�� *n�d�;��+ޘ�r��AuXf�o�!�a@��A-3-mv��%���@����R��Et�w�h�L)�!`�.�P]W��>ڵ��=LFe��;n����Y�{枚A_�E��V��L�2�e�l��8���N
؜��0�_-�*.h�^ONQ����	�7gSF׺��K�B�W&�~V��s��ym���Oݵ��=o�,�����1������������:�����ߋ�`���h�R�ÖbӺ~�>���i���͐��3�X��'�Y���y�u������)dE\ڙ����q��b@�."g^��<�Gpʨec:�=x�L	�S�"��W;����¥C�V��޼�i.x�v9��L��J#=
)��4DK�_��`�HX:E`X%�&��3oL��S�{�e��Y7]�f��g)w]�/��/������W#����LL��4��0V��h�����:�M\�!`j��i��S<�m�������[��& ]}����g_�f��[���XZ�T��[N���v�r�r�:�s�0{��$<�Vdȩ�:�ӥĮ�_H���e���"�9�ټo���Y�wa�)w{��KG�6v�ϟu��BC�z���N��h�ǃ5gWrͻ�H�\�}�	gz}ט����'N_�c�y�O�;)�=9��z'��m�/M�yV��3Y�%���b�v����n��兏�'����ֿ�Y���z�].~ދnQo�c=�-�v��#�I���C�RE�rOa:t ��Kf
�D�4���ҡߍd�lR�mQ�"��![B�~���̶�%�S��3����t?-˨um�$¼�bЦ�M�",������K�5�HA�?.�b�Gn�]?6�Y�k:�tn�Act���9[u�pQ	�F�l���0�3�P��!N���dngt�Ũ�~�����ݝ1�o�Sv�7D�~��
�d8\!;�l�����Rj�C��?Mܲ��;��w鶘cuy�~�gr��:�4e2���#�5��r��$�����O>G2����w�C�
����k�~B�&1�tc�=�RΦ��ԩ���8B�jSI�sSS����s���D��Ϙ�y���ӭֹ|w蠇�����Z4�������C���`���y�22)���^D?T~惪X�
��t{�u�yu����Ե���v>�ٙ�(�?@�;���$��<uԐʽ�zu��NY}Sy��f��vam����i�鞚�>�<���FU4����J�]���ColZ7נ��%p֔��z�c�c�lT��Ӕ�<�Q�\bb�3��&)��Q�h᢯n�q�3�8����A,qu��;|_�8��S�1�MtCSA���E9��-��B����qלns�
I���������(��@o��z���!��x>D�G�ҩĺP`�^��i��\n��K/>\{d��Q��w���Z�4��G3�=0��d`w��s%�\��~1����-� S+8V�&�`��I����-�4����MW�.�+֢�F�wSN��+ʷ��zj�3�.F=�}���6f����!;���rsD!�.�?9�N�z0�Q3�Ѽ!�6gE���!�E�t�m�Ym3��욘�k�ޜ؍��;M4�s8*B�{%;�5��=x�j'��ԢV�w����d���QԂ�=6�ݷX�lT��m�9���*�c"0C�~�[g8��Fi	���,����Җ���
q���<��˩:�v�d��y!jg+��|�LE�hAф�	s�"k戮���gT�خfY,��fWz�%Ҹ\uJ~8�t�f��_Z��R��U�%{bѷm�ꃜY9���7���f36/�!��u5<�ZJ�)�d�tor��~��˴d�;� s+�����m���P���Tu��ɵ�0O�P�\����%��������<D��%Fy2���GI	��i�]Ƀ.��X�˩�'|�^��̶>βeʟJ��%ԭ��X�4M��4���ؠU۰+�
gf�,�kž��^�)f��,�9�;��}�S�����m/�}���(A����-��)d��
*���KuɊd�퍍�^ة��&�!#��a:�N�A��XO��K��ʻ_]>z�5Oh�d�>p�2�׳'��f�P��0_�{���
��?+��yb#���b\"�Z+�Q����t^��ni�;�.D�eC�`�8��P�L�S\&�L���T�Q~ȇs>gFZ&"��E8�1��sp�d�'l�FVr���vI�^����������
g�SA���r�������]��?j�{zr��y�\&��93��{�!l�9�y<5�7t� }�_#��#����q�Q.[�e1�*2���q�N��vM�F�mp�%��ߞ���=j���Q��օ4�q|�~���:��t<R�FLVt@�C�%��ػ#�v߶S��L'�c}{��Ez���llm��:�*+���p�Y#1���;��ߎ�]{�l9�ɕ�i4��C�1��#a>1���UdY�O��75�Z�D�O;��3�:i�Y����ٹN@���r#�2q��P�\����ވ�ǈX	�I���iO_ �Q�/3p@*=��Y{Q��y��O%�ʳ��-9ynuMZj#.[w;~1p�~u��m˖�U#������l�8�}��ec��*�*�"��g��I�C+xŬgA��Ǳu�H����{�ke��8��p���#�=A���3�;g׃����>�e�f���<�;k����1�C:��û7q<�1��'{;,-�N��PU.Ъy�q�u[��W0AW6���,�Йi0��J��/|�K��N
���dK�T���[��P��i^��#z�&M�_)ɼ��9 7�bZ�p�6��dB�k6L9sL��OiBxՓ�u�I~"����B��\+KЗ�/+R&�_9��r ��,�����D'9��]V��5�$23��l!�����'�~H�?os��Oע0V��ʊ��-�U0�>B�^�s�s4��0��k�6��V���h�q��Wd���(-��y�49
�s,e��;=����<6�5�W��x��9GLv��
}������;��[%�WgSF�uU<<���C�~G�%��]cϱ,4)�ؾ���(����)Ix�8�6���1��c'��e�wKc>�u�4SB�a�e]8q����]�n���̄��t}b�m�ux���<�Ry�=�q��������m�1���m�1�����co���ch6�����1��P�lcm���lcm�66����������������������Cm�����lcm�coͱ��6��m�m��m�1��@�lcm��������co���co{lcm���e5��W�5 E� ?�s2}p$��;�U(�*��(PT�����D�U)B��"�J�P�����UUR�	QRU ���I(UITU�**�DR����3eU*)�6i"RJ#l�D���T��T�[h�HQB���)$Kc���$E$@*�R@�.᪎�U	���Z0J(U(B*�$����	A"I�T$�*��� P*T�B% �J
�}��(4d!   �
�UQ��U[ �h��5��D,�������X�]��L�	���AeL���- !@U)UT	�� k� P��� QQ� 
)D�(��QEQEq� �(��9���EQEQn+qEQ@QE�QEP��(��(��ƨ��⪊)J��@(�+� j����j�v��+Zkl�3Z�Jn��n�pU��nk]7m�a��l+4gC�la7i]� �Y��J.��0�t�*%DITQ) Wm*�  	��L{9�ٻ�l��]��(��m2�ɚ�Z�:9f��
��0��+C�t��CA�����F�nQ�fYӪ�kgpmA����@H����I �   1˽n�vV�������b���ݝڛ��n�妁�+�uF�����JUv��E��m��Xۦ�juSbcJj�ֻY��A��IUJD�-�iHx   �s�ݜ��b��k�)��GZU]�-��`n��:�Wm)���9S���J����]��ҝ��ʰ4+Z�ln�����V�S���J�%TQJUU�   1�=P�S��SP�U�Gcv���JUݸ�vv�1�m�m����uͩfQ��us�\�.����:�I6��	Ek�J��*��   C�m�2�J�Vզ�k����N�f�2��N�V��i�Xvf�۵�MYT;�g\��n:�� (Qr[AE[%JR�)%-f���<   3.SZ�zh�ʚw4��խ��ջ�$Ԇ֗a��]�e��J��p�(���]l�BK�����+f�m�ZRln�*�*�	*�	AT	B^   GUu�[A �i�m@GLU(m���(��԰S!�eڐ:�K�;7e0 (�-��x��T�Pd21�{FR��  *l#(�  "��	J��@���UT�L��iD�ʥ4 hJ��H&��&�"c()��D�Q�DQ��?o[߾��<־����$�BB�2�HH~P$�	'�!$ I?HB�$�BCo��L�?����ox�|��bKfLgn�'�z�ק[`]Y7��X@i�f���x�\4�u�q�v)�'%n ��⬎�)R儨e��J�ok35(����t�T�PK2-V���N�h�H�h]�m�/�������1�3]��m	C�h�n̵o5K���yZ��4��e`Z�˴�m;�p^=��v��eH�P��yp䭵aJr�ur\�5E��v̔��/�U���t2�YE]�B�;6M��Te<u�J�`^��X���Yc(��6�)�(N6V�7cJmleG����Z��J��J��wwa:�`��ZM1�hhAX�Z@7"��
�Ňz֨܍?�C�oY�Hv�d���L�#4,[X�U�E4��F�b&4ktc�w��.�Y�՚�n�aia��ⱸ���$���,��3�I�)�k2�K;�!���W�(�k"�W��5�L��^���إ6�!�je@�[u�B�r�M��9Kf8dT	ȳ���U�؀O��@�ԦvѭH��՛���a¨�Њ��]W�P��D>�N,CMi�B�FL&*���w�,X��e� �΍�v��V/�㵈�PVOFi��{)ު���KE�/V�CZ�sv�C5� �F�/u�E��y�K�f��=[p2�s�X�/s�Zt�巰�@*Րbֽ��J?6����WV�-ekE<0GH�jX�1��ٴ�־����j���Ġ���Ť2�U�Xbԥ�f�ܬPSsX�ɲ�e;���@�%H� �f9��ڎS���$:�W�`��i�
zbs��0��� �4�j6��@ދ;@�w��6:�`�%t���e$B�[)��1Q�r^�5�ccv��`��~ct�\�b���M��X��GCX�޳/2�:�0�Mh�Lu��7M�zrV�׎��e��bHh�к[E��3LM�R��n��Ǣ�i=�i@���ڝ)[�0FX&3)�ܓZ+m��M���E[fT��L��&f����ą˕W"��M&��J�e�!�q:�tZ4�kKj����]��f8�`nm����юS��j�j�����iۉe\lD�r1Jn�T�F�T�t��*[�-�
��`ݫ���UDKu�dA2�N�w��n�X�R�EJ�{҉+��M0ԥ+�b'�V�ۢ.�T-���O.+.�:�6M��P���V>�  [�,ڣ���kDW�O��]*Xf\9�Ƣ�fJ��N�1�(�J�j䙂�-�7jL��Yh[�١���ו[�0\�-a�G�j
j�v�)�	�N��*ׁkcȶ��DL���-�k�L+TFmf�Ĥ���0֪�t�d��b�.٠�0t�Ck��nT�jdsucGsq��u�������p�ki�V*�G&���V�z�6ƑYl^�:2D#	E[�̥H�2�<�8.���7D������Á���bnX���]<����w���+��a��#t1�2��飨N#�4*`$D��(D	%��rIf�ڧbZ]'%nH��өl�����`�Q;���ǒ�K�nST6�����6����ڀ�͙��f�w)����ˡ���f�צ�4m.-:ĺ�716ĭE�ۭ���6#̠q<i=��k��t+v�coe���-DQ��T/B�[+��gP5�;���0:j�,�#h�e^�Edf�Z�Z��h�d��[�E�W�֐�JՍ
���yfk�n8�:
��Ć�x�CqP���ZUbkY2 ����OQu�����6���#����M 2j��ach�����6K�Q�Ț9c�)C����`;�d4D{Z���h�ʖ-ہ�4	��6X�C�֫r��.��1�;C?b��^j�R%�͍���)�3)҈,ɉͷUy�c6�|�m�(�^��P9��:�IYr���n��U��s.�z ��aP-3p��Źr�,Խd����%@�H�Lbu���z�ɰ�W���\(��fjSQf�2�H2���T��x]e�+m h���F9�۬1�5[Dx���)�z^f�1�2�)�ֆ��<�+i+ْ�hjC.VKSu4H3�8�u� p�o�ũU��A5��)!>%J+io�h-)/���$����X��L�p��wSdN,N��NqV��{t,mB+v�vŦ�,���ӲջCa"�8Q���(cx��9�u����V�'j��:�f���b��S�X���E�����'s*�ea[��!;��qE�Qs	W�#��V-@�5hաg)�u����ŀ��CɁ�b����/@��I����V��Zn�x�^���Q�*6.�hL�H��X1QY�$������ �V)�j`�/���d�A��P�	k��r������թ�Dwif+��Y[m�Soq���ؠ��xmZ����V��eKXwo��y�ɲ�Ť����<�� N�\�*�w�c��e-x@���I��q���ˢt����ؙ���dۣ�عv�V�դZY�$�X0���XZ)e�#��0��D����-�-�]�%�˘u�d�(Q����-�U�Z�l֪m
���37qL���o繶�e���a<�MR�Zi�g@��	�E���Fׂ�F�Mz���YS�*��6���̵X��Ϋ�7��j�<J�I�7:�{���ut�j��۱���m͢���F�6����I$�di�',��_	V���ͥNZB@Ej�.�,͉��ڡZ&G��@G-�g!*IM`�x�=�Z��eb�x�8��q�Io�H]��O��ʰm+P��銮k�'m��71��pbȒٺ�2� �i��`y7ZOA��lZ��nҬZ�j��&<���SEެ�WL��N<9*���PdÚ6)4�1�V���kp+�Ñ�t�:��J���PVv�せ�[&R;�k�q�6lf�	2Y�BU�b�J�)n@����;J���!��7ոQj�ҵ���8B)En���b��(72hB��%``L˵�+�h�ݍ�2g�f	Y�Y'7n��`7#[z�[i�eo
��9��7,��e����TcvG#��ڧ�L�W�\�����B�S��H�Y�bש|Ue���X�a����-;ľ��7+`շ[y�V�U�Ô�-@���M�&X��J���Fô�d��3s�W��/#�r,�n�F�؎2v�;������W�vp����uB�̷M�72���cR�&Z�x��Me/�I)�Z�`�����Q��΢�^}����J�,�*5����+P�*��ؔ7r.�K�.cXEL�&�XYV�k&tZ(l�6�C�m����`�O���а��uk�*���ø�էp��%\T��jPժ�2���҅��/d������ŎE�Y��$i:�0�KϋM�UѶ,�f��v���u�����V;ϔ�CQ6kF���Te;��r�d4ݺ��#�J�W{��H+O3�t��6Z� n�
|R��
�1;Ÿ0
Cw��]埖5$��h:�[��1AubQjL[ze�Mo5!%DA�)^��xq�<�Lir�v��(cY���W�1����Ů�ڐɢ� &�v�t��ʒ�U���.U�)��e�l]�Zd���f���P��B �
����7�hӁ		F��eݪs�얝<GlU��	#�y�W�쎵�S�r�� .�ff�ïHL��DV�)Y@JH����xELٕ��lFrMi�B�$��ϢzL6��8�SZ^�,����������06+ImųvT���!�%�-<��C��zCvu)�3[*cC�	L���,U	q�4bٓA��^��H�P;���d�U��4#�{���6�+�A���*�]�;�R҄ʹe,�(����� �{PS2lSh��c�KB��K���kYYs�9��q�o�-����#r�ْҭ�%)�+M�72��hq#p���P˼�MᎦ��InV�m�;�n��In&�h��n�K1�J�"�⩸7����*�ct��KK"D�Ud�6�C�l�K�E!���J�p�Q53rkn\�e�t����^̺M���l4/[@ޓ�X�r���h1a��L=�W"�m*����I�f鳲��@|Ņ^V�j�f�,^.�h���.��̨�&]:g+LTٚ� �4ÍeH�]07YHےczpi�I�b�&�0�6�Y�E�HAa��X���N����י���G�bMQ��Ko�͇0�0]��jݴ᚝�*���K@�Ь�b����a�]��=P$!ǘՐ2�r���x��z(��eb�8��+
�v�E�2�H��S�MaW�"��b�.&�|�ը��5y�=	�wJ�������n�\+)��b�սKm�SR�z��eZ�J����yh��cU'����m�4-zS�-�so0���Qa�1�A|*�kÄ��n[W�@mѓ 7"9���U1T� ��8)�Z���$��f�YEEunn���VC����n�0�L�i\u*l�.��ާQ����1�N�]4lQ�5��Ȩ�e�ͭkrbv2�4�0U��i$�IЬRf̑��vR�kD����+*j���n���	GA5dQy[B�@,�X�oE�N(�M
ƥ���w[nE�|�'�,�nH�o]�#b޺�0:�#5�Z���n�ɔF�j��A �m���Ej[QVh�-�]�T����p�:RJR��`���7s5j��V�L	��	V��BR�l�v���o�k^c�N���T�X�W9�&	X�%^�W�v~�v�iW��Tv�)f��`7��fV*�ɡđp��WxBv�f;ɺ��:9��C�;���Fl���:G5��#^��q{H�,�q,@�Ӎ�l�����)b,�4�d�[�M��4e6���4KOb8&V��f�m,d��n��GVD�ڎsv�cbm��a�2����$�8�����K�5d�O#o�Jc�������5�8eH�=��<M]*CZ3bzV�J��걹�u��u�"ث������R.�4���"&�S��Q�:*$�FVSD�6�v�̻h[�qb��pS��B2�3�ڶ���Hd���;+6�j�M�`�q;�2�2)������J�XE��4 ��L�d˫�N��*b`I	6͖�w�[d��[,�B͠�_дh�˱%gV7��3��I���$Fe�̱��l��@�H�Z�Zt�pw�/ �;�G5���Ct@���Y[�VkRY� ���t����w��P���Fi՜TMI��Mב3u����Đ��Ҭ��TA�7b�L:�L��/m'Jd.a�,�E��lif@�#b�cmӥt�Â���\yW[�h��6�����)X��<��̕���ZU"-MY��i�����U���(�+1�j*K�V�k����)>���*�4ޑ�������X.� M-����"6� ���Y���8cPX�[��Xt��G�Wdl'!�b�n��*���q�ܽ%[E7�D�B-�g��η(e����1�o�:��m�QZ���[hV�^�ܵ{I��Q9�yf�N����F�Jh����J��ЫVjG�r;Ѐ-Xb�Ո���n�T�.<���!��Tl���.�J�^��yd��q��i����
[x+H*ñY�-\�)X�����[Aۥ�h��wkb�X��]'JJ���7�fn�3<C�)�k�@"�@)�����tC$�b��i�go]fVj6��q ��1����'&]�l9bQ���* Sз!k#�u����f0�,�f^�\p�Vt�Z,k*ږqƶ��k�.�����:��c)P��e�tS��n��Ӈ6��a�Ŭ�B�X�ڭc��PU��EYj�UY�W�Lǵ !��d�Sl7�U�j�M��7�u�Ӎ�i)le��L�K�n��1l�l�IRN0h:ˈ1����Hڤ1X��7`X,V[�3�Y�Y"������D��,�dV�DSoWY[d�@���!�{�;�$�ϢB��C]O��$���qJc	Ok#��*��v��l-*��/v[���@SP�/c�[`LaxE�oDֶ�m(Ą�Ǣ(Ƨ�;]�����GuVkC��9y�޵S߰,���GC�t6�j�P�W��U<�m�p�ˬ��*eL.:��S{�PM�w����dm�Ϳ��,��eY.T�XTˁ_���T����.D&�/H�Y6�^T���@�7h&�YV��[�P4.��՚z@ue���b�r\r�C�f�����y!�(�y0�-�2�R������[ņF��L����4i�Y�[��ï6�,K�����"8�ia]��h+f��k5�8���F*=+jf�Z,�D8���i�*]&/Q�ȧ�n�[�H�nf�\�G>V�Rs1*��:��m\�R���֖�����]</����P��+4�-�OH����Z�	����f��`��e]�a�n�D��Q��C��Z.4%[���T:�^,��Y���˻&������f��Z�,@\r�B�j���rm��:(J�TB�U°^1F7��}��X����75�^�pU���q�F�-B����.7�(e���pTU���J��bnm9�LRP��r�5���ݡt�+��&M��$�Eb�CQ-�m�`V�^�D+WO(�[sV�L���D�kl��C�0.�6Ӭux1m٬cl`1d��;Va�j�!Gv�!@qk�6h�5<gZ�GTi��{}��R�#�x� �y���(�T1'��w�j�vU����"�q-�1�5ϏwWEp��=��ӫ�@9����fQ�b���f\�I�����)����&�7��6o�z�I�����U�q��K��=�t�� \4s����i�y�y����5��X��*!�҉Wڕ��Y��9��9n��ZU��4�6��YV��Ӯ�0�_G��;U�c������zV!�����xNz{E�~|��UG�e��:�O.T�c��Wt0�_e�Lݶ�캻@KG����J&=3/�����p��=�ħ[y����^��4[X`�4WWoS̷�û�ʆ�*����x�2�O���B�˜q��c��f>�ǽ���&l��l/u����ah4�\��Z9>Es5����������3w,[7�Lb+�k�3�.��Z���u0z�^���'s�9���dn�i��ˢ�eBP�`c�������gS�w��К1M�k���6��r�e�)Ӣ�����fۓ6�b�MX�� F�O�Ineg
j���������ѳ�:���C	O�ݭu
C��bz^���|�1&̍����:��p��"*��kV<!�P�u(�Wk�A�`���p3,9�u��S6݌63o�t^�.�5`uV��%�f,�w�볛h��gr�|�m���&Xz�'�oDı�����
sȱ.�!� F[�d�dr�o��):���:E's�t�o�F��r��7hc�M7���wk��7�kU}�8��UJ�Ҁ����/®�`�������|+U�"tr��J#�*D.yM��%���:da�����Y���H�r�C�-:Շ�x]�Z1N�j9���V�j��|0��;V�LN���o�>-k��0Ⱦ��n��x���(�e�r�ɶ�85ub1�"N�i�v݋�a����	6(X�+�jZ�S���bT��]ʤ�M�^P Vv �f�}���w~J�2�\�*DX��:x����e	xY[f�ڷJ^�Q�g8�ɯN��(ǧv��ѝ��:��|n�5���,���eg-*e^�oNcyгw�2�n�<���9��g᪒���>}�
�Dk�tufN㬎��p[Yz��0��In�(�O�Ys;��'��gn�$#�W:�ʾ�i�;��u����J(�N�J'Y4��8;�Uµ*�OmRicڙjI��Kʑ�or
7����**���q���	�����s�)��ռ�5�Ѐ�\�e�����^՗,QvE�5����c�U�v���#�Toe�N�Bc�.�9�Mǖ��{#�����K�����<l��s:�.B��q��^�ĝa�)�����Z:�=Ã�S`R�727��c\`v�:�2��C��+��8�2��c���j��A`���C��훢�e��(�'֝�=-���y�D��VU>���i�վ{��[E�՚X�Y��u�F�y {�r��v&��u��ݳ`������8*dd�"���)� �9��qz�Aew-Ji�i�k���	�X��~[P8�
����7�����<��;=#���7�����`���E�(��	.����\�U�o'-�+jڜh#���DI5vv��t�2�Ҷ�n�� �����[�5+�(똼�MM9Z�
clr�flxњjNp�z8�0�.C��f�r&uLku�;[]Veeq��T�ۚ�pt���\5!��P���r!:b�p��pXI��g�4qG��̊2�^R`=�������g#[�*
�)3zbK�v�ؖ��.M�E�:��AZ��J�x��L���8'.7ҁ��{+�T��ȉ��[\���@p}�����5��nV�X|'b�r������y���%sܲ5w�J`i�jKe�G9����\!����N��g����*�޺}}Qmbeu����G�5QlI��0P��舾�U�V�u�oZ
����q�����"z�|�����\���2�W�����7%ҍ��c�]/ ����c�Q��C����;{hN���e��;D�Ð���Z��7����2�����C��ΌZ����L�#W�B��7�)ͽ\"3t�)�D2�Ia�u�n��e�����|�_%���縩�ACU�ieb諳�U�T�.��ܼ3]��b�LVw�mG��_ʍ*�<�ݫ�X99�pv��6e*���<ƽ����J=/V*���k�سJCw�{�8���FT�]�)\�9��b�[�j}�t����1ע�vM�=��E��Q����f�*ͧ�2`�H5=���j�J�ov��\l�WI)X�N˽8�w�wt�}l;��6���9r&a��I���AfdE>��<k�i��ȩ�sz�YmZ�ի䃈�ZT�w"�s�R�2�ŉ�b_,�tO<�._kȡӥ�3&ܕ��C8�.�h�X����]�9��j����ef��R��e�����)�;y+�n ��ڕ��� J��沦�k�t(:v��yl#�d�v��hq�ե��-�PI����^�(ӌ���,���a�˝�BΠY���j^)�c��������;���klTW�N���"9u����t2�Z��)�k&�/^�# ���e�pd|R8c E�ZZ�A'P�0��F�u)�*��0�Ӣ��z�������-h�s7�D��
�����Eo:�q��SvC��e�wp���.#�d8n��'�vj)Jr������*ȝ�r��ՋO��ؒyt[�|���n��[W�{V].�^ξ���V���׌�օ{z����u��>1�Ii���Gf�qj^���MNgf�R��֙���*H�ξqn�d�4D�]b�ـu��Æ|���xF�Y�me>�����rW�Es\R򙵌�%d�}\4�@�N�;�pv�#��[E���ͺB�.8��6�$�;euoT]A�����$�a��]r����-Ѧ�v0p�
���e{sjh�N&�;�e��s9�-0�ہ�轚5�O�x�﷕KN*��*�p�ݹ&�g^س�|tҤW1[or�k�OS�2z�۫���	��ۤއSgV\壻Q���]��/�%��P�����1�;:��}H�E���.�⻑囎͙L��9�	�dޖE�,�.�����ۥ��<��:�O�d�����2�=hC����/j�e��ZWid1 ���ޚޠ���꽷K9��DM���w:Η-$����8�V�Ƶ�-��b�Z��X�r亷�1����݀F���g�ڳ3�Y��a�u��WA��h�z���p�s������i��ͷ�td's�I���.u���,�G2l�hq��W\$�����8���d�O%c�.�u+N<n�#�}	{�=�M\�"����+#�����T�k)��}�>��R7��Bv)]��T/i!��F�`ɔ�� �s��;���m��3���Ǖ�cS� %i�����%��SsC�gnP���"�c�K;��r�,qs���"�� �%!��*L��Wz�oPsze�.
�@}�VF� ��ύ��lld�\�λ�r�\U�P��ް��Xz�x�
��R�V���Y�Q"����V'4�Qw�M�����h�70pW��4��|�ή�T�7�f�oL,8+���d�K�B��ź�w�?<Y�`��	�����(;���:7Fp�Ifޤ���v]wu�����讜�5{mX���)�P��V������Ow�%��I>�+vc�|��������^�mԥ���q�}�0�a�]i�A㹂#���Ls�+���*���k^�P��AҖRMۂ�@��n������ܵ�/*w
`%��3n��FZk����PCܜU�?<���빜p-� �:�_ti��`���`�P� ��0c��	g1��km5�Ϧ�ӭ���oy/����d7�:�@&�=WM-.����Xޒ­����7�;{X��:��()fY�βcG�V�|���x�j�]C�Z��Y�%�l�Ww!���*��sX�pҧ�C�����!��P�*�yک5�6�^A���b������mVg���&�޼�S��m���+����XN�3-�Kg,������x�\ ǔ���Tzqw��WX�\���9�u�n!,Rc�kB�=�V&�va|�7s��V`����g�56�z��m�䄱�ŗQ�SԭW&��Z�D�o��.<��Z#���b/����]&f�����9�4����:��&�k����El��4x��D�Y�C4Õe���u0�|�c��Й�;jʼ�ZF�6�z��%'X�|{Qwҝj��:P�@���"R닁�����j�:a~ʛ�,h�*	������nu���%�yc���tlnq�R�	�ncYf�c�r �4z�3G�4�1�n�U���s�^8h��%��	)W][[��J��u+����Qm;�A[��>��i�.VD����w�� ]�r�DЗ���dn)󶺲���-R��@��ڧ���RZ���2�}��ܝ���l[����J�C4:���lg�V�`MV�N�p%�Tܮ����(���q.��O�id�_Hf�&�<�Eޱ�7ר�2�`E+���p���F+,���I��Xqpʺ���w��vXI�tjn���`�4Э�����X��Jແ����PC|�b��u	�8�f�'� �t�Yb�Q6����9��. ���I�p��v�d�}�r|���u#��T�_��:��n���!C;o�5�M��KUv�-K�k�x�����B��s�r���hf���Ӷ:P�55���7:S�\7�����X��(b��o�J�V���܉k����b�U*���΋��fv&�Y�*>9{z����B0ұ�V�Gz�ݬ�����4AR��*ӗ�I0�+�\yI���j��'΍�lW�S�hV�x���1w��oL��c�qo>9CAǣX�Q�����0�8�un��6��>*��Ҷl�N���Y�Y-I�lY���<�{�V</6r�O��ֹ���.cL+��'���U�-Kc�xpt��g����i�y��E�xjJH`ʒnS�%���(�p�㱩R
:J��Tr0�;�נ����0�*��tF���ޜg3a�������ܫG4c�l���VR:���XeG6v���Ȇ�AY��s~�ə������Ĥ���lo
'nm͛ҙZ3TB�]��KA�V�/���.�y��P�oqn�uX�%Fk��i����)�א���I�r���֘*����tC��ﲭ˰ge
��0 N,U�9r�d*�a��fv�<� ��X�-��#�j�7���4oEP	<L�K���vqBJ��^.�g�Vzm4��3����9ʺ�n�!3X�-�E�*��1}��iͽ_p;;�l�n�rB͗nK��YWL��C�ۧڕ�ޭ���Z�6>������f�pL�F�[��	`�[��je,��-����X&*vVh�r��!�|�:u�0<a�U�ay[OlE�F4Y�Vq�MAI���J����v`ћ;ݍ�a�{ú����N'�#9�㷙#/e��Y�è�u�x��<�l+��Mj�Ԩ27u��^��udŲБid�^���x���Т�Հܬ�q�\ɽ��_G�9A]$[;>z�;�eSYa�1�n���Z�\h��M\�VC��J-�z�ع���-��spd���u�ĉ�گ����=g<��F��b����[3��׵n�j����������b&i��0N��t�VL�{8(/k��[���ȥr���h�hH{��]�3T���b��7Q�6��۠��g;�+�%b�3��)VT��0In���8k����ۂ���D +gd�f��x��/)]�tj���|�3��9��.T����ư�Kg]�6�w�[|��v�rF�t6���A�r���o��a�V>�#�mQ�o)��KI"��@�se�6��m��Οev��N���������,>��9�k�����:�EJ8�BvuӾ�Z8NS��U���ո0Ӵ]��V�s"�,�\\Χ+��br�Wj�݌�H**N|$r��+�@ϓ	���U,�)��_u^[x�E..	��W}gK�:��xM#�;�!���[������1��o�n��{����]�|��hee�����+�j5g9��]�r�[���g��ӽ�_���\��'���϶Ӵ�,��C�p4Y|�c�Ż�[kizh�7~�ں�¸v����[y���]�pP��+�R:�h�2���{y�c�,euI����ԃ������1�ø�1�9����&n�V���^9ú�lH�5����m���b�i�c�96�b���'�E}to8V�iE8̸e�+��Tޒ؄P0����A]Ejn&����Gf��I+Χ�*vޚR���w16���<kzt8�f�Z��l�3�:��w���hG�#�,<��U��5Ɨm�����`�D��Yfp쭋u�q��vd�G%�o�y[��C����W�/�V�y�o��*� ���-8l)X���`�M���ك2�|��R�,�1

�H�wd�z�쬤/1Ϸ�o6�뻻yӲg.�� s��jq�v��k�lA������+z�!2�髐����N#���ԺŬ��%��Χ�9�M�>|�o=j[<n�<Ɂ��f�Wji�:t\S�����iK����	�$N$J)%
Uڴ�%�%�+�*\ �#r�$�-H�{kie! �������G�˔�=�mΦ,�:�,(�:������u����9����o�?�$ ����$��Ѫ��W��U'��[�RV2`죹�cn��Gm,3��ܢF.��T�K�V0NLޡ�Z�o=Dm;[��n�����tj���q�, 1�R�U}���
j�ǯ�"h�1Z���JN��X�F����ɑ��e�{�K��pT��쭼�nl�j�Z�i��X�ݼ���03َ|�6�"�2&��#��B�0�Τ���7uDr�.!��w��y�ɚ{L��u��:��,� t��r�"]�1s��P�̕19\�Ud�g�;$|�.�V����w�o�u�T�9��6�4��t#c����W[���Z}��o�kܔ/W�bv�L�L=�a��c�η��n��n�,�yx�8��M���d�r���Z�
�3
��(�4�`
-�\��i��*7�y�zF�͆;pe93e��� m��\�wu��$CZw��vܛ2�^�֪�9$\3�:uf�X��e�(�h�iԄZ�]ڗ�%sm��҂v��R���u���c�+��$�[�5X%�y�q�U,�|�=q�Ǹ�Pw�D֍�ά}��P��c�����%�K�U;��*Pb}�oy�*V�I<��Ϭ�y#�/,�O����]}�`<�L�_�wmw.��e��;|.�Vx��j-���z�w�V�C�2�`R��<�x��$���P��O���ofh�n�:�X��՝�����opO��6��$��>��-��^�$'eU�H�Xz�fm+:s���B�oN�U�s;n=h�ѽ��� ���xրiÈ=*��B��S�N�OJ�L�_-t��f�<ï�����P��X:�Uм�J])�֮OtLS��@�
�PգQk��j��ʊ*2�q0u*T�qbkd�7N���Mx���M���Xȫ5��y{�"�n�f�>�f���Cp�!�&.I�����ǃ��T�c��O^����W���	>�m5=R���w�xT�%f����e4t3��i��ty��bc���^���U4�x�j�o��
�����]ݷ\���q�r���Z��c��/{���+������oq�"�սu�Gn4!N��%�+��f%zѕ�U*&�[�|8Ձ�N'��m���-���He:��@����Yq����>�>�[�c���&L�)��sh��4Q��v�e�*nn��F,T�$��3�:���.���Z���&vRҸ��eӻ�[�LR0����!4�p�4ǖ��d�̥��cTb�Y�hAF��[>�%��$Qyt_3�.�c�:gl��Ab�݊c��:��	u�w�$���/\�KB�ޮ���c۴�P�G�5ϡ�{)���X*��IƻwVM[nLW@.9�ue[ۻ ���bӋb8]�{����8��н�t^��yg9 Mjc#��v}?��4X�F�
�ã8�ӓ�ʎ��N-����c���]��P�m�C��p��Y�-[��+����<ۚ�n��|OKP�}��+\4^�m>.�l�3�z1�v���YϾ��6��Ơ�(��>;�tۘ*�D0�z���lH쮧�^����-e�r�!����Y���X����l#��}���\ig*ÄE�2""R��ܱ;D^o`������O)���X��M!�C/����32��b|Sy}��s�9]j�5J��T'bP�cN���[�N
K���ڀ�diVuP'�D��"B�"zU��՚��d�a9V � ��%հ9�^8�o�-f�u��g�%y�nc�W�����U��@��v�ql�|n�E�'
�g�Q�p�r����A4NH��T�	��=K+']��Ȗ�G�-�>F���ur�C@)��»�`����c�[vSf���rm�e�uk%б�]�XG�٣��#@��� ]���	h���H����[ƈ��sV ���b��V�[�,:MB�,���kr��kV�It���A<F����+1�Y�M��Of����j�����K���; ����i�u����c�kg���G�W��c�X��!��i�W���pH`Yɤo,�h4x��!Ŕ��"�t�굌L�lev�0+�O��vՉFȾU�'S��dxl�>����{sF�Q�7e�� �(�0�G���+T �n�s�[3�
���e1z�#7�FegsT��\��4ZԲV���+����:���f/>����y��h~8�V��A�<�[�C���x��F� ��{n"1�:<��}b���wo,�8BX�'1�crj[F���:>��H�f�d_m./��-��[���v*:�#\���6^�d��zH�q��}��أ�}�-2�:۱�I�Ea�����B�/tv�1����`��4�c����Yo��y2�5vW;�!WY&�כ���Xp��g2��2^�u�!��q�.md�w1o���(.�J$����nUÝ:5G$䫝ǒ������Ʃ����~9oI�o��o��쿆]q�N�B�R�tb4c�N��7u�r��߷����˴H#��K6^�u(u�b|ܷ����knb�uւ=�v��9��&(/h�9�Ģ��(p�۸���nQ��.p{ˀҎfoƝ��W�Jm��j!����ǹ[W�Ҥ&ӹ��<*e��'���I��:ͼ" �z<10�jپ��U���uO���n݁,ư��F�����6w�����	����I�G
�_d������Y��ͫ�jm+&���;�6��V�(5��-��m�*�0����Clos�t����Vy*9�c\}��Mwk�DT�ϖt�crq��w͑ ����L�X�[>]����%��Lu���|��{�zs��c�(��sIu��Dψ��'k���܅-�X���,PTOm6~[����>Ѹ�#�,cO6.9���n��Ġl).w.�˸��\A�
�M)Q#�55U,�����ѹ�޽��U���#��s���n�o+Q���h�����#�[�~e����2`	y�x)e���kK�
��(4���{��J�ܽa�H�V�'4��Z��rnl�M��U��1�#2ͽ'Y�)G����kOwf��-ԃ��c�����D��c�ǒ�,1�6��d�
���F���خi䭊K�k;��sr�`�5Y|4�	����.�]�}*X���NK\P�E�֌�ͥ�1ѵ&U���e`Y��P
�{9K�[r9��ʑT��r�e]e����]�+�jSf��k���{!�˹e�|�iUsNgX�Lc|��·mC%�2H���aU��>W*�V��t=Z�����*.|+3OX���v|[���۷��w1�,�|�6��L�ܼ��]��Dn.��4J{�U��k2��M��P8�R-����u�Z!����K�t�r�[V�f�E���[���MU�t:U�fs��DT�l�X�B>}q}T$��h
�������S,�)��r��/��;dT��L+�U�RU�㭸u����6� ^х��o^qiM:=��Nk���_bS�*u�u�r��al�����]Zb��X�9��v��0v=��}��*]��*�'��:*S7�Xu4�݁@Q=n��n뫔�r�Ky/8T�3�u2���J��=�0<��)�B�{yۡ�r�L.�Ѝb�Muoͦ��� �'��7����S��;�F��o�Ǘ��C٘��������ܕҵ	Ϋ���wn���z3϶h��gA�03%@�O��}��u��+p�ڹGJ����1�g�1ĝ�v��/Lw\8���ΜBF�
�Hsrn�'R�VVAw�9h\�0��ݼ�p,��7`�#�N�u;{����y}ƅ��K��8u�Z�p0@b���WO�p�jr��h;�R=�5�y��Ζ�I���D0��,{J�c
��I2�)=B�r��ܺ�)�of�Lǽ��c�N�Z4e�{�P��b�:�.���������L1�ox��C��`B�J�N�[��v\��1���������*'q�1mˁ���u״�N�q��)�X�g-���z����q���z�-M���tac8f����n����1��j��A��sf�����̥V�-�x�����}o����G~��_t0�EsF��A�v镚�Y)�y\�N�_f�$f��h��L���^@���[�y��wG9�������Z
Gf�C�x�N��K�����J�ks^�Z��G[�l@������/t���;�Ӱۭ��n��
 %���S��c{.%�oX��P�4U�}�3(�]�ä �2�6����6����z�֭ǔ{�u�b���[����櫷��#[�P�`Ɇa{���csGk�ϧۛ(	����{����%_v�CC�ࡎ�M�Y��4���I
i`
c��:,�eT�W)�`����u�:�`��¹����;;��CVV��xKK&gl]C�����uu�-ڷ����X�]���_Q�I����Or��*Wn�*��%�nY[.dҨ\i�*���P��F�ջ�V�A(4q���86��#����}�HbQ	�3:qf[�ҫO�*���G.���wta�D��F�Y{Dg>�D�����X���� �ź��M8��˜_]`�N��;Xۖ�s/��#T5M��W\!5nO��B.�.��̮�C�A�ݼ0���/RU�e^�m�łôMW&
��<��r�h�sqk�r��x�1v����$T�i(����?�;s�[D-�f������]̪m3\&�N�ݬ�2�#\y<�m�j��P�ᕄS�W�OP�ŕ�-�J���aS�P����f�j$CYJ���ֲʼ�-(����of:��B:�~s��ߐw�2cZ\s�<D�ݴ-�B����D��]v�!��L猜��A��Z6k;��N�.�X��A �Q�����s+v�O�QY���V^�e]�]��ȶ�]��*9j�6���yuq3Au��ݝ.���f�Z��)�F�IȦa�Sj�L�Ԍ��M��em)B�Z!5�XJ��$ṫ#yy�����3��>̽�q.��Sְ��h���i� 3mV�J�0Kˤ�(�/3q�t�z�.F�Wmҏ����1�7�X��0��=M��[��]��%���R&�\0-<���z)Z�P��e��D�ݍ���>4�	����m#�]4=�L�}l]�{:���@`�֠�Oo)%�9�TO2�'W56��ym#�W]�xb�N�R�V�7]�.�E!Kv�"�gY��ሀ:�4n�&���fXr"��Ya�d��HG7��tΒ���WTǊ�b���§"��5i V�B�Wuyb��$<�.�*N��D;/B��`�� ��*:Yg'+�����Ýg8��L��;��S/zc��t2g!0�I��{[�
��3�D�Lf.޲R�֥�!��n�.QT0�M���ig7S9Z��&�6)���WmM�:Ӳ���%�є�{ҏ%�2nd�"4)ީ����{Y�7���JDQ��,���L*=X녡�۠.�I&�:N!�6��������Xsm��K��6�1R/�C�L��Z�d9Y���c���N����7�:�m���"�g٬\l�߯?k�,t&VfсLo��Qq����.��W��x����Ք�:���ԵY�[Y�����Q���l�sMgo3�ś.��ѣ�}{S#�.��Q�s�;;d��{��Rd�j�.ỡ��=,��Q��f.�7rK�M��Uc��)��+ށ�����]6�:9����qr;r���,M��3�I���O.O��O�ZF���C�B��LOV��si�۸�����������K.��b��"���g�� S�i�������������'o/���ڷ�fjne��bHm@J���
��U)rO{� B�c�Qʰ��T�
[8�*P��f�B��p�0�솟:}��7������#�-]��6c���4�������+�;!Y�Z�N=當7���x���]�$�����Pff��݊��V�����6P�k;�n�� �4�RUn��`���3Vb;2��]���U[����'wk	�s��ٌ���@3w4ە��"��ӹ�x�Ư`7�0��|t�����t�y��T.�:2���6̳���^�
��]@Wj ���ʷPc0�5��N����=1D�*��GX�1�b��ls�՗�-u2C�j�G:�U�n�a&�'B��e5ȌI`wX�YnV���i|S6�I7e
� ����B�7�I�BrP&�S �����T�u��1��
��
�raTƧτ�{��y(�2�fr�6��	\P�5�T���"��w��K&̬�E���U���;�j�$G/��i��*�NQ�N&��q�y�7�T�+;yê�2��=фa�3�,���h�.��}�Ҟ,˝���@K��z��)�Z+{���Y� �)���[����]<�{��=�H�=�9:%�x���F����G�9�;�SU�������ыf����;��r)�S�-Q���k�:����t�{ee�t��;#��#s�#D}V���u�����"/����J��v�4�X4�,�Ys8�ɹvT=�r���ۛ6й���ݱ����`0���F��JO�U��=�l��=���r�V�\zd�*r<�����\ˏ�W]�Y���Q�ŝ���Y67B��NE#�I�A���3W�K;h+�&%�yʺZs�]w�_0�P��Ɔ�K�����n,ù�PݳeM�\�u����vX��{\�J-5cj	����MӬ2�$���Kr�Yf�q��`�<P?k�xm���S�:�᫩�I��sq���9j���l�J��x{����X���R��|�ӄ����!Y�;�v��M�N��r����B��jC�U�Ɗ���p0�\�8�wΡW}�.dN�n�a>G\�eA�5/
��xBݖm�Q�GnW�}�6ˍ��"��B���<o��ޥ:�V��;��p�*ovoYv{���o��cj�;��I��+�����A��0Cf�E��B��rM̦w�*�l�T�/oI���Jѐ��K.��C���k�ެ�ޮ t�WҹLbm̹�Lxښe��=�p�6+F�U�j*��Q���U��!��򮰢�l-�~�܊�vҲ�'o��>���eG�n���i��9�caZ@��+w�CtjqSR.E�윿PyAu=��%)�H��H����gV�}���P�;[���%b���*	�.�J��Y���;��q��f	�5�/����y��.YM�2*h���}�Q$j.�}��o�|m�m���d� =����A�N��
�8oK�ch|�<�iv��48Tu/��uv��wH��M�oM�.�u�ͬ��L�C�|�j���K��A;/�r+O67;5
�������fN�U�j��db�v��>ج=ߐ���F��N��)s^]�c dG�u�VR[��s2k���P���j>���	�h��c��,E�):4P;ҹ��8�l��Ӡ[�':�n=ͺ��:R��n��9�%|�d[�6NW���U]��X�Qv�����E��J�mm�O�c	QEAA���QcmaYQQ�Ef)TEX�͖�Ush���� �b��a����+L�KeS�-iEb1�A-�ȱ��hڊ�ƥZ6ԋKEX.+����Z��Q-�*��J�Z�hQT �m5-�Aqk�b�ŗ �*5��.1�F
8�Em�R�����T`��d�*���,c���-TsJ��j1Qp�UUX��qE�	��UK*�e���h��G���UJ�F6�3J�*"�"L�"� ��ڢ�8���k�-����a
��p��b�䵈��
�A3�L��0����QQ��ڪ�0V�1KhֱX1Z�A���QQQ�,qe�#\b��b�ciU-(�mAD��V֢�,E�i[+ZᨸU�}5���߳�Ը�A3��KEj�FL�s'�	}�٦�.����gY	v���rcb.u��wlE��ݖ��M�3�����.=1U���1�*nE;���q��Q�u���@W��o!�|����0N7����[�}{~�{E�����*C���:x��C{@����B�5�f�˝�E�q��,�p�k�T�y�1~m�t��XZen�[E1�G�f˿T�[X$X:���l��ȉ��
�E��Z�ۜ�`�Hmêt�3�'�ٻ�J������b���e�	__P,:Ik4nB2{e�{n��TMpi����d��Եb{�G�l�K�w�r��)�
|ݪ34����\:��<�Q���hއ����{�����D�a�C����s֫1��\2��>�Hזc�ǻ>[�N���>�0��T�K���1�w*�Y��Y:2�Y�y�֦�<Ow-ݰ��������v��������i��qy�#Z/5��<�W��m>Е>�I}�O"A=�gۙh�v����L�*�k�kUp��Cbgk�e���I]��.o��kZ��bsY�}���P��r��P�f��[a�G��m�փUݼ����J�Y��r:�*�mo7Θ��E��M���)V˩ngj}}��3���Z��{�+��88v�k.;8f��eV7W���m��uR��J�	�����S��z:���r-RKV�#9��6��ݿ*�J)FXl:��f�ht�R�|յo=�՘��[�/�쳶ƭ�
��y���t��R�/�.�"mg�6 �Y��$�Y!$rw,�{�%
�T%=��lr��3��-��t%�&uV9y;�#"�d^��-<�B]x�۱�NEf��9��M�~�DF��[B�5X8�ܗ|�U�_���G^z���(׷
����Jn�	�`�#-s��s.��X�dH�G�B�W�[*Eq�Ϳw�B�N���+��+i���ZڅA�$��xЙ}�
��Y�l�<����u9&��ü:i���Ԯ�^���&��;�`d��]9}�r��N.8��k���'��u��^�Jo�w��!���
�1�k��ט:�9��7ݪV��+�xz֤�#�/�$�gch��{�d@Z��,B �A���8�;"N�K��n������~�3d�:��32��8�8����7qol�H��[�=7;�.���
?oM�;��ԧ�<}Vآ��K����ީq�*�g}������H��z�j�*��ưp��{�=<���٠�c^م��۲�7D�x�f�T�\MտO]d����/1����,ǥ<��[fO7�74n�.��Z��3{-<q-���ەr+)
��B���\�ď�|�;-���ɥc%g��]���k�_k��*qy�~�zP���rQ�Ž���oW=�S��r�R�a�}��ov«��F�(�t/M��lMW�XJ�c���o�E�,-R���By��j�j�W��krA����2�l�hS+��^���cϸ��#^��s�]{w�5�V��JP瓦��ۆv�6V*l��)����;�P�B�i���n.O��9u��$���(�;x�}���ۭ���@������s�k�5P�\�bAL:��6��,�۴��x����
��,�\T�הW^؄�)�[��rW����ȇr�7�d�y�UX8�ef[�Ί���M���CY5���tYJ���a�oL�B�u#���i�U��(p<�ΗVy۾�jT�*鼳ĩŎ���1l��Z����"�^@M������[L@<�qfh�c�.d���K�8���|���oS�f=k��ݹ�z^�^�dH���]�e2�M���+tm]v5���ebq֨�Z������Sv���ԥ��."���n�O*ljU9��Lv�x�j͠z�$f�y%�Nr�7y��妐[pF�L�M��~���e�ܛ�uxzE����7�
H���wM:U;'�,H���fښ�Z�Xۥ)f���*�W�2�ӈ��6(%�O	]�=.j�x|WG����z�կ���!V
ƫיH^c��z�f�������|u�׆\��y��S6���н���m�W"�����D�7�s�8m@;�z(Xk�k˰�W)���)��5�z(3�x��O��W�إ�N�I.�����{�n�7��>��=�百}}�tۋ�R����>�B��Z���p��N�|����Bҝ������5�W5��B��Bf�+U��o����� 3���2�ҙ��=��� �V���M�/%ߑi�kݧۙ�v�6]�R*=i�=�/�"Jsd30m��+H�W���Ղz���犅���u�����>]`sYJ}itY3����h��GRP�Ɏ��<ȷmU�E4�WXS+nlN�p_$hZr9j��y��T
B�]aǪ�L�ŨʮSXʥ9`jU��2����@ĩ��L�F��$M�E4�-���bw�a�7��J)�R��B���!��+��˗M駳ۘ�gF�9oy:��ޛo�ߵ�������|t��v�Dv.u��3�,�`��p�f��9�{�a�
����Z���N���k̜ջ3uڟh�a�r)��tB��j���@�Ch%d̕���_l2r�+���ҌGe˗�-�5�'س�C��eO��S���W�<�E�	X���ǝ�x�ˠvhەM{qJ]k��OS��}�ci	mi��kԣu�=a�1uK߶�C�{=Y�7Wm������JA���5j0|+ˋ��^7u4�w��n��א�=X��AL�vner��
G�2�p���qu>��;�ݱ/��GE"�u���r���T�3cX����/�oV!������U�ѐ�42��i�7YA#%s���G�m���<� 7o뾥���M����nr�=y6��<�(�s4NV��}��ϲwbj���-T�+���nN�y��5x�\e�h5�M���kg KKB��uaOF��/��4�C��n�����:��5�{�y��I�ٞE?j��\-�Q�c�J�Bc��E�++%�hP�S�su��^x���Q�9Qg���)�h�4�VE�������@(�ع��hP�L��S�U{a����9=צM6��cY�׏��l*��ݸף����AX���_$h�x�z�؍	Ԯ�ي��Q����~�5���U�
)FXl:��f�4:�����)�ܶTd+i����з�b}�3��2[V�ɾ�{���E�
���=����N\�@Ħ�UJ{�����tCl��-��K�rje�XB�Q�]�n�:�[�Z������R�1�/ds˸���DZÅ�K[`@Y"���y^/�o���ԭW)�#gE�������u?�+!���,9��wF`z ̡P־��F�-d�a��G5��P�[\��	�a�޸���;7����n�Ox��g.
��$��0u��iF�_.��u�D{���3Ȅ�!Ҭ�ܥ���*�R�+
��=¶�]n�bFw.���mQ)3Ƅ��VM��W�O6�;�<��S��z�n��7���O��h:�vL��<hL�ɹY7Y�έ�X7Fd�f�;��vիѕ	��C����oj�
�zxuӗ�0�A�e�3���\��w=���7�h�s��+r!������:8P�Kî�����y�Puc��O��*���Z����rǦ��2C�����|�\����%v��l͚��cPz�ī���-�!c1��.}�����돜r�^�d+�o2�eO(R�/3=o:^���HfӃ��%\�R���+B���=a����y�m?^�~�8ߵ/K�����V���Y�J.Lp�p����һr{��Ovv�X���z�ߞ�۞��f�J�x����n��V<_R֥�w��J���k��%��g9��)ތ|���ݵV�E(������=��F��%�zhO�̆hhmv�]Դ|�;
f��f[7u���G�ݺ��:Yl�4<�zB�ّ;Mq�d�+7V��eǒ.3K����ic�*��V�N�wk���e^��^%���t|���X�����IY�6�Ί�b���Wy�m�$s�>2/�5�J@窼:� �8kZ�շpz�)��	�-�u���]T��p��̭�7=^��m5��J|+qr|��˶x}�UJʉ{٪ V��k�B�����t�}as�ƫ5�P��Ԛ�x��ފv4���s==�T��C�"�<)�[~��EqSZ�
��nvm�z�=x�d��d�ׯ7��nG�0�Sv9�)3�D�� ,�L��n硫�:��rZm�ss�� [��U����:A�&Es<je�JGN3f��2On����4��Svzi�{C�y�R�3b�[^�T�d��b�K&����ӹұ�SݳbVH��B�Y��޴)"�s��,��-WuVrŽ'/��\�u�-f佩ŗ�Ui�b�RUٳwS9l���2:��-��a�nQ{��G8�v���{s���옚�@v۸;�6�,�o,�ǖ�M�RJ�X���<�'��n�/V��r��CI�:��XD�$�18� .T*�ޜ�AXr�-�¡fnj}���Ku����'$V2rg.�W�Q���/i�wK�Goe�97.������4�02{U_���}�����L߹�YM�ps�ī��YZ�r����������WN��t��G�Y�w ���vh��VZ^lir�\�Q{5{id���^��+9��7CS{oS��Owo��i��oTM��&.э��O�/\E����g9�*����Oy�̈��+v�r�����������l�9<5���_$hZ|�oB�Y컸��͕w-��oq�pޭ[�ët
�9z�u�2�����\d_5��J5�j�>٥ʮm樉�ͧz�f���j)�RވYS��#��'��l�4�'}�z�X���}�����-�gW��e
�C[`@X]��i��z�K��F3��ծ�׶!9��BV�7/z�
���)#��l�O1�� ���c���eas�]n`N�a^�nG-W6�U
���DM�g-ov�ʕ그r�t'5K��O�w�\�A{yo�.t���Mc��L�a��L�{��������@�=��F�xbHۧ�U�WP՗�ؔ����ņ���cG"/U�ͫV��[)��.���;�u�ۺ��s��A�w�Z(��cO�K�����=���k>K1�;��#y�1tr�[&b�ԧ���ykX��*G?�d>G�a�L+�]b�e�ǐ�����q����D�,�ٻ�V
�KwNʲ]x��9}����9ʊ^y2�5�0�X�X�l^N����.�($^�2CwSA�8��۠����H�r<�������/��/=K����pc2�k�h佽��Xri��jc�U#,MvN�wJ�o�6U[�{/�����X��H�Y�w<�ux5}7��]� ���q�H?r������R{��LJ��e!W�
�}�oSg��=�љ���L�{"��׃��ok���ʜ߸^l\؏N�*�3^�S�R�� �K�iM�,����g[	��t�8*��ݸף��_
�	��_$V��ټuXD�S�Oge�o��i�y~�m��oʭ#*/a�X�+nhs�6��U�-���#sT�V��w�v�s�n[���hTw�ҭ�]���U��E�2�%R:e?z'\���亵^�O�Y8�t�]�t���d��}˩��p��v�����m���!��7g�unu{cI��̴P�Vv�f�n�X6�*�>����l��E��!'�v�
ָ��\Z	�V�L��>�������h����qm�ͷxsI����M�K����z$�޴A5��qy�[��cu���� Nd4�ڪ�l#	3l��)J��^��BӼ�����emo��&��cfX�Ȫ�Yf�4��Ld��EoO�]�&�7ז�3���'`"Q���ε\��%�c��ux7���v�k1�[Z��hށ���c.���t�8�E�ö�X�;2>�3kBm;݇��;��j|�-nR������*��KKb��lJ��&�@�ӾU v�_Y��ws
A���*��{&�<�[P{y�fH�U6W/�9�q�6�u1��rI
��NEt`G
Fcp�{��L ~۳��k��L!��ũ]�M��KK)��v;%]>Ě��|3Ĳ��d�j�^��D�C񧵇W_�^bы.���
���Xb�dQ�����&U�$���n6xL���)%�Z�'�Ns�<�,�ub�9t���ڞy��*�{ed�Q�oi�{�	�F�v�3Λ`Mo.f��.j���\w9�K�L�V�k6���`�����_:��Nq}0VqU���e_�����u�r�)�& ����;�Xص��M��]�廱i�]]S7�;a��tM�\�:�QX��FV���\N>�3Y��z���!�Uk'HQ����l3�5���,���`(R�P���[zཬ��(Q<á0I���{s*�Gד�p:'r6�4��]+90)�����C0gN8-�Y݁�����8�:0��ΰ͛�HNu#@��Bؔ���Z|�lVqμ��[���_�0����{i�������;��L�z�U�,�1
o#���!�P�)=��ىx�C\pl ܕ�QZf���Z7z�͋�`�3�a�� �髚&oO�p]}���\μ�[�;lÁt�+z��Y�5�U�cC<7f-1�
⥬�|��=K:Nކ�c���v�f.�ssz9�!�:�Lk��C��_:��blΠ��P ��2����V�e6��[(���f+,�|��ug�V5����::���k�U�lg%j���V;{��Ϛ�%�T;I�G'$ǖ��*�<�(n��Ǵ��r�"%p����F�k�78X3&Ԭ�{C"��dΧR8N��Fٱ��ɽ�m ]�3�* ̹�3S`�hB�[3ZJ�NNؤ�@�b�}�EDcR�r�[�r�[�c:CW��f��[@�:2�!��b�r�T�w�u���
N�K[.�Eܖ��2i�	�u�J����L�p��\��7�ɳ�ob`#@P �� �	�l�0�(a��H�l�(��5qJ#�\Ҍ�RV��f1�U%�+R�5�����m�G4���Dr�p ڢj�#����-��Y��J����F"����Tb(��*1VĶ����X���m�1�"�VƲ����(#RT3j��f-d0��&e�Ԙh��cp��*�
9aP����8V������1��a�
����qjڵ%�ܸqZ
�La�r�J̸ŅbDQ0YP�,G(�V���9Lc(W#�F�[Z�*�m����V�S�-�,Ub�fs3�TT��"�e-�,
�b��b%�qAb����J"��m�0�
��[aQ-+�c.1�[sj�B���eE"���oN��1��ǽZ_W�ȟ:�F�^��B�}�����D���GZ�2bŬ�w��3;tкw���G�63�Ʃ�NM�����KkVg.�*�[؃��/Pn�(�qKa1{۱�
i�\�ۦ�b���7;@B�>��/��P��69u�
mR��|��
%��Þw-W��=��t���@�ۼNEf����=��q��ٌ��V��UKqb�#tD�3����d����yE��½��TShVdM3{��o_p���\��J�t��BevM�Y"�S\s��V����$e,���w�{����*c��.C�D�g����0�.��]���^�����w%������h����I��!�0����]y��QB�us�f���ø�Ϣk���1��>]aM�ڒ�^�8d��ӿf��ͱ�t��Cy	�U�zU�ӪN�2����m�(X�߹���hf��J��ʄޮ��~O+ �{J^\����w(nc��\�q;Vs��^,T�N����t�_$��$����<4�����.�M�P<����yTWLX��ZB�cw@���W�9[sC��wq�}H#K�v��Y�C���ia��'Wu�}�Ԓ��.�s����o4�\�xy�;���˟Mk��M���e��v1S���>�� ��yvt�{�M����U�e!B_�����s�^R���==���������-�v����ʆ������:�i��AfVdĝ����;RK!J/�zCSx�ǜ���~UyM�F�Z:��-(�J"��%�EAj�j���mw�G����C�<�c罞v�l*����Ý��*�����yGXv3�@���$m-窽з�y�ֵ.Z]R�:9P綳�ƭ��m��C|�l��B�"�Y�w�qW'���ZU(�������1=��v��*�j��(t%� vWG`��{]/rŮ,���a����|[�z�%�sa�WcX�C� RG�y�[b�ⲵ���F�T�����V�vs�o�k��p�T�{K��X��<jev_¹lz�׹%�k5c&Y��ΰΞ.ג;8�6��7�0ķ���螮g����ݘ?zt���?'�a(9��m�)����܉P�ԷJw�x҂M������H�j�MW����-̦�ᘆ �+���s�*I�n�f֔Y�Q�1�
ggC����Ẋ�%p!�:�>}���wo�G0J��\��]=hp�o�ᆞ+d�ӝ��9/�����9L0�d�x�V�q��I]�37N06��<��Ԇ�{�?`�	���!P�M ��s8���Ԋ>����g����?I_v����Nw�VV�wIY=v���pO�>I��l�XM!�i'�j�l+�&M^$6��2n��C��Ͽ`�'R�!P�&س��:]��L��lq��۟s���1��,0��<��IĎ�ė�$��d������@�M���d:��3<��'y����	�5x��f���
IQ�ך�?v��;���;���s��|���'�)��&�q�Ԭ;�B��'�}�OL�xw�̗vI�P�`�M>�<�1
��&��0<f��ӨN$�VCl�'\_}�s���z������oQcނ>G	��y>�ed<�16����a��p���w�c�I�OC��2]�L��y�)6�����6��4�c����w��h�I��.La@��ﾀ(�"6RM!�N�'�׻��N2�sx�I�O_Ro���>I�y��M�=����d�z���}�|4���I���.\ً�úν���e!�=f	�'O>�x��'��m2u���'�8�?S��I�y�1:��l'}�:�봜���{� ����
w8*�X�>���E�[��7ly z�?��$E��cI!�0�3a����N �xj��d�T�݄��Xg�q2�q���;�	����'Rz���O3v�s��˄{M��q�k;~3��π�=��+��`yߵ�q0���dP��I�>9�e�qSFl4��bg�C�:����q��S�Y2u����I����{�˃�u���������<<� D{�s�N06���5��Hx�fL�6���q|��2�8���&'�ağ2�<a�N�|����s���?T7�����e_�ƺ���g���BWvm]�V��b�VD�S�WGMN�&�yX���z�M[�e�3��e��aS͚e_�iYf�ZWF��k��\#�9i�[�su�>C��䩲�r㧥�F��n��*�7�ܥ:_v�p���3�N�?{�H{���	�O;�I��G������Y5�pE!�>g����.pu2q��c8�>Mb�$��|�d�?y���ϣ`�{ysʖ�$�8����z ��'!���C)�l'8g�:���&S��>C��''�������%ABfw�:�d�'��I���*^�5�xp���c�����}�{���i0�q:��'ڲZd�&�XVC�Ӷ���0zÉ�&S�=C�x���Ad�C}�T&���S3K�q�E_%����y�BN�8�>d�5��u�l���d�L�Xzɽ��@�OXzb��H{���'P2}���i	�ў`'�=?1ʾ���л��ܾ��{�� �{�C�wY��I2y�8�����ɜ�N$��n]��@�fj�Z�q�O(|��d2n�06�oXh��!��Py��_za�rUK��}񕵯�}�"H>d�;=�q�<�9�b�u��癒�I3;�:��}�^g�'̞�u�	���˶�7�I_Y�^3�HD����Պ��N��Z7Y�]yӚ��=Hm���<d���>�*d�<�pAI�L����$�K�fJ�$�ؑd�V���:��M���Bq�qp�>gùVj�ti��ϧ:2�7����=a�x�t>��!�a��,������N��9�
é4ʇ���&�3�Y<a2���o2Wl���D��q�9��A "=�O�B�������7Y�����Cl'gi�6��&��&P���	6�C;�PY%L���N%Bxw��IԞ�����
�l�ﺮ#ޢ ����>�j��`r/��&��q��x���V�x��!�CI��m�!:��VOP�.�I6�P��b�i�=�2q*���m'Y=��}� |��&8z���|_1�����D(J�Y��<7�M.�:n'��x�R�VM��?fp0���9�e����Zaw��7yd��yyx��|F>�e�\�в�,���P�ۍ^�i䖻��k"���	�u�Z����p٬�Syq�')fs�:��J�)�uhe����{�8󾤙@�;���L���$Rm����14�mSњC��|���'Y4ɴ:���t'�8�~��G��_9{� ��%Ѯ�S�4�e�c&���w�ޜd��{��b������=�'�;��O�0�NnȰ�>`}�bi���	���$��pd�'�Փl8����'�8��>���|��{y�o}�0���|zx�a8ü��|��y���d��&��I�Rz���&�w��u�Bz��}�'�9�M$�!S�r��Y&}��N�`_��W�l��u�|����}zM��N2�yBz��3�q�$���ĝv�h�L@�M��h�q'X���s�f�ċ�&���q"�C�O�F;�,��z�o�|�y����"��9{X���ďy�� �����z��Nj���!�N0ϔ봓�<�c�=~a4o� u&�Y5=� �C��w��'Rsd8�2q�7���[~t�����y�q���d�T�'i;�&Y'Z�Y>J�ިq��N��2q�����$�'�������ޘ��'̚����m��o������F|��.���ݻ{���� {�o�� C'�,<���I�50RN$�x���	�o:��C�C��2{���8��;}I8���0z��&^d�]�sWJ��v#~��Y~�|8�>����I�35�2J��Ϝ��
��VO;�ĜI�4`��I�ϖ5$�3凩:����}CF)04���=�A�o�y�R���?q��� �}#���Beџ�C��4�{�d�!���2V(L��aY>J��s�8��M�̈́�&�&�:ԓ�ϖ$��z��ێ�ng3n������V���d{K>zbM�C�2�u?}��q�d�1�!�=d�c�d�<��fJ�$�~�XVO��y3�I�O�7�a��&����?�?~�M�>�̜c�z�`
�u�D`�n�c���s��Ĥ��l˿%)�be\셪�s=�HS�u	!�AqJ+�������S������h��&o"N��:�e��P�����`[�H�j�r���mJ�����9ޫ��[X-�P�z�S����z~�������J��d5N�6�	��u������N �<�1
�Y6��';���'��<I:�R�Y��a:�_�D}�U�	�+Ҍ�H�&�6?u���='̜d�4�hfug��N��6���!��R��a�wd�I\o�Oq!��b2m+��
M��>�+�G���B��r��c~�7��Ͻ���|��)=t���q
��&���4'XL�Y���<���g����d:���{N �J�=��u�B�N@������>���.���M|��y�{�Ra����I�O;��%v�uydRx�����V�4�5�C���>Si�	�O5C�m�2q[�&������O������ĹU��o�޺��q�L�%d:s���'�Xk�����y߷��L�xs�䞸I2�w��I���q����=Mf��!��6̤��4d{�@��̀bGgYo�#_ڹ�϶�Ϟ�VC���e$�7��N%d<o:���M�k=d��ý��z������	&S��(|�0>�14�i��$��N߳�P�\�a�����}�~CԙA@��'�z��Vy��C��0�x���d��	��� u'ϩ6wX��Rz�s�d�l'{�����|�=�@G�|�~�N���g�?[��l�fY'�;�AI2��Y>b���O�q��Y��O�u�g=�N0�ӌ�t�zo���=~I��u����Pg��ٔ�d}&��];��-���	�;9�H��<d�5�`�I�=f�C��3�2u+:���8���d�>���'xcz���5���<G��u}L��e_��-ߛ�8���Ӿk!=d<��!�e'Xj}��d�;�a$���I>~1a�O��35C��d�6�q�����dz+LT�uW�u�V���o�� ~N�m�x���g�G]g(����՝��"b�����eV��V��xi��yk	d��#U<�o3~��o�.�f꾩�ӌe��:�-�^䮡 u�1e)x���ͥ|�,���+�ݳ)��/�\�.Ӎ�4��P�|���7��G���'�|@��{��Ra�}��!8�xw�B��
O>� q2z��,��L�P��I>O&(u��IC�$�=��s=�oE]�v�N�?x
>χáG�������XL�w���f�5�q��q7�fJ��Ϝ����);ha�M��$�M�O,>�I�;ǘ�o_�����Ր�gr_��äx|" d ��!X`u��]��:��bz�L&\r��3�O��y$�o�̕	�9����%d��p|ɴ�5㋤��H�T�퉺ėpc޳�Q�\G��}�(u%v�gvq�ԛ}CX�8��|u	�O���8�$�7��'P���� ��0�w��++	�w�w��O�ٙq�lp��s����y�ޙ��>��4�;�	�M��n�O���RWhM�C���:��|e	�I�؅C)8��s8���Ͼ{��=�w�/^��u�>���}eA�S�IY8�S���@�'�SS6C��f�x�$�MXm�z�ɫĆ��0�w@�!��g߰i��)>�Ϛ�}�1�����K�}��]v�4ŝ�1 ��&g>�O'Rh/5�.���~ċ'ΐ<�pN�q&�Sy�`z��МI����	����a����7=��LS��_/�:��}� =�#����'�)9�&�u�Ԭ;�B��'�}�OL�xw�̗vI�E�Ri����b��M;Ml�g����.�38<'DP���M�n���ߚU���,�ěA{>��C��� ��1�:����9f�u�iXz}��'���y��e��{��wI2�w�"�o�;�B� #�#l}����fɧ+�\%x��HT�Y��2��N��m���T�Hu�NS��I�y��8�����7���d��&�� ��y���z��V��2G�DP߸_�vXW�jɭ�Ո^�ڊ�b���%F���|�݃��M�d��TinL;ݗI�{=a�)n������mg%�1s��'*��ܖ���an��CEg��4mt��x5#ɢ9=��+z.�]XH�[��U�G��/d�i��;EZU?��|$��?2Hm3	�4��O>�x��OT��N�v�|Ì=��L�M3��bu���Mw�d�'ϩ7�p�����Y���c��'ޚ����3�Q���������q"���C�cI!�0����
I��pd�
�Շ�8�ԩ��'�:�'��e$�ِϽ�Ǉ���ߊ���#����~���ǿ2|���?�$���O_�|�&����8�Bz���$P��$����$�OC6AI13�!ĝe`i��8�Ĩ�=�Ͻ���f���bb~��M�,�	r�8ó���O�a7�P:�N�>�q'X��k�k!:����É�&�����OY�;��N!�jf���$��Ň�>��&�n��8C�|��k����I�N;ġ8�S�L':}�I��G������Y5�pE!�>g�����Ǚ:�8��G��!�O�X�#�g�O�~��_	��?D�3����l]y��k��q�q�8���C���O�:��8��3<��XN2y3�I��)����q4ɯ{�)��<�u�*
=��Y8�ý���sX��k����I�M�'i��P�e$�<1a�'5d<-2|�O�+����6��q��<��'P�M� z�>�=�ﶀ'�� o�_|���~�Q���������\k�T'}�XT�����pRq���	�M�'�>k$�d���M��x[8�Ԛ}a�Cџ=� jr8�20��!�sځB�C7ty�;��1�����d�C�ߵ�*T�'�c�*O�Y<�q'|ɷ.N i7�k	�<��J��8������� �� i��3��Y'V��ͮkz�z�:e	��ge��s��z��w��$��ĕ*I߯RVOu`}�pN�|��S6�L����<�����;�g|<�KN�.����y.�<!y1�E^�,Kq��Z��uʖ�.��Aུ��%���v�#��y6��**����YX{�7��4�^T
�u��7�d�T��1��_-U3?��/��O_6� ݝ|�5��E�+�3��:��ʱևd�H�)O-�J4L�r�W��>��'��� H|��8����1
�Y6��9�Rm�'{��2N�Լ�d�RN���O�`xw8'Y>I���hN0=I���a�kE[���>���$�����m>d<��!�f��:��*o�u��,��!Xu&�P�����l���x�e���y��d�>�,��|�Ef���;\Me:9��]�_�@��w6Cl&O)�u	�O5Cl6�!5�I�*ӈ,��7�2q*��16��=eC��*M2zw�gԒ��K��!�C#;��m��������q"�o�9�B�6�N٣4�Ol��0�m�q��$�C>��)&��w���J����6����=�>s����惡r�s3u���$��}���Y�I�;��O\0�O'9��}`xw�d6���h�!Ć���2��M�ɴ:���t'�8�~���Oa���t/�����O��w��7��sY���|�	ӝ��'̞�I�;��z��]�$��߼�>p�e<咰�z���14�mY�њAd�&}�u��,�{#�������E����q�ٳ����I�=�,&�vӌ�t�zw�8��O��o�ĝ@�'��<�I6���C���;�"������I�8��	��_W��Q�?e�l�ռ��>��:v��>I�T��a����I�}�N$�F�bRm����u��y�1	�C���Hrw��N����ժ�Y'����\}y�=��g�� �:f��)'�C��%`i'�:�̀0���y����j+�ٻ��>v���`.�aOWd�/i;��A���B��и��v��r�����X�Z��r���[ۣh�CU�u/��έ� w30�k���f��WbZ]}o��M���y�-眞��Lwr�@�o
5�8�r���I�0�52�Y5uat���c/V��i�˳�]�{f�y��t�.����[�Z����P�7�uf�@�r�[��4����>�B�Ж��вX]�����V�@̓h�w.�Z�s[����Kһ�6艥�K��`,�⦵���c 7莏;7��dֽy�I쏎�������"E&x��웕�l�Ob����x�^�������������q�=��	o���:.����52�'EbZ�s:I��Y�|�eR��-��Z�t��=HRE�&���0��`���ݻ0^�Z�g�W/vH��r8�|R��`b�
oV�|�ju+��h�~�3J��\�Z;��'Aձ��l��5m���@�lEּ�;i^>1<��;e��-���8�����W5���yH_��m�v�5gy�Fպ�sz^[é��}�4�6&�����ʺ�B.�H�L�=L^e��zx0�t�n4ib{��v�wѦ�P���<��+ܪ�U���Z1����V�6��k��-��@H��M�NyU�Cq� �a�Pv��R���WVVSb�lG;32���])j������Z6�4pM�'k�M��F*r3oe�+n��JJ�#�e*]gn�[����5�]M��W&�����K��WIg8��B�s�+�5j��ř���	��;\�eL�����[��K�D�v���`�cÓ�vF�/�Q�]L&���Ï5Φ�W��&5P����Vr��Uɮu�����Qƅ���'͆�u�W,&�e�4��^�T���]��R�T���v���*^
�;���4�C&�J���:Җ�����>��!=`f4��RWd0�b�f�ipc�s��4
zK�G욁�����C0���-L�V�ws`uN2����XGfh��YS ��ƅk�(F�Y���7A���׽i�<:�B1g2��oF��^c��{���B�%�k37S)|�G5���0�,2=8�E��f[U�e��)��s.;m��L��<J!f޲���gXF5\0Y�����!Տ���W�&[���-N�EDv��؜�
6�itF��('`�1Lv�1W�$ΧA0`S��L�;:N�ZU��4��k0��s�&���C�*t&iWC�������؜�B��F�u�h\#X�ra�o��X���b�x�
�Q0R��������X`}��q�wb» $k�(�ow�G��ۧϐ����d�]�Ki��E���!�_bW��z�\�mZ�ە���3}f�s�c,_���
gt���>^$�"�u�E�ëk�n���Ţ�8����4��>���#�2��eTrc�дSǁ:������8���YaŚ�};��]j�AhT�ь�z%0e�[)|cbNv�ݬ�)b��������۱�S�J�����"1̠��o�\�Z�����!3�p
wk5�+`�]\�*�9c:��b��$W{X!�R4�Et���3]'����kps�gYV��GV������N���Vl��{c9�-u7M��k�;��9[����jt���q@v�{J�K/K"d4[R�ͦ�eya��C���ϴ�3�̓,�8�k{�YL���e��M�j���L#N�xY��,�q?��u�է[�唻�}CH#��H��{7P�e?�-�y|,mL��|��փ�-2�Ǧ�Na%OT����+�Z�!NYys��+熻�5�a'�i�#x>j�&ꭼW[��)��q�єIb_t6�K��T����l]�w%���Xv�ܔ�*?x;�<��Պ��˷m�x�BlWL�n�bڍ��y��[��i��5kP���΂�[���-%q�� L�����S1:=[�)�R5��!b��G��T�F��VquWo1�u�1ś��}�P���N$��evP��ݵN�B%!�m����jSrwn�A������5ipw>�}�q����׿
�¢�TPiB�5��Y*(�h��*T}��$��)�-��h��1�����qG��)V�KcKj�(Q+*�����B�l�-F��h��F�A��ܤ�f�+R��%�e`ĵT��J��ʖ�R��m�m���UW4.���5�-B�mG��RکYb9C���-Rѵ�Kd���aj�*E�--[lTE[l�˚X�j
����F�e��6�j4�1�E���EmR���-��P���En)��V1Qb%+@��TZ�KR���U(��ҋ�kJm�kUB�J�Kj�DF�D5b�������[�8��d��m�mG4�
[V4��k*P�6��Z��P�h���*����|� ��>#�F���svMrs���q1.�kw�q;��ۡ�l��;�\x��}ٗ��M�i��W1�kb��{v�^���U��|���j�̣����Ǻt�N/yM��ہU[���*��ˋ�(�?x�N�dz��S��{|�f����ҭ����pM��ce<����Odg��|�A������䬭̦����O�,�L=� Q��4�U���8��,���^�S���g3."x�����^\�����;����s�8�bj�3^�jm��Qa̐�.��uʮ���Y{�L�T���T�{˪��j����r��'�v����^�P�Q&��T�8�v��C���<�euĚ�}	�����|5#�}�ozY�}\Dߛ�+#�:�]���G(���e*<+$~�/��Ί��;T�>wǆ�rk��l��[�́NzmY߮P�X$�a���@��-�VL��w=+����{C��z��KFC@�;��E�͉�sl���W,p�A����.������TO�� ������m�e�'�T4,��h�Ug4D�{�J�M�̧duN�{ykX�f�_�l�#Kc<&���S(�L~�����N�"|o|��F��g+�\^��還H3��N����v�lK.�ee�\J鎷ӎ+�\�����M�j�oe/��ް�f*�\~�u�O���nfsOo{^v��q���5սu���67В���ݯ���v���n��׊��pmܬ)�q���| sVr[w�������fV��Ή�d�������6�Y[ӠT3�뽶p���}���{���P� .�}\�o���v,5pt�}�tm��ߏI��\Qx��+�L�wH���\T�kī4ks�r��li5�;j�E�:�_0�};g����U"�5p)��(��zi&��+c�Q��eX��N��)�V7)#����')@UӅ:j��!�;�3nѺf�{nxH�=�xN��;3(�_U���pl�]'Tp�my�?y��LWdD�o����ư�38-A��J��J�>�!�J�o�1T�P'] l�E��"�K�fb�6����Q���[����}Kc��;��`�b���+l���i�
�R���>%�;Ǣ���D��gdd��p�}\m˥����5�g:�D�UG�Lڈ0Q�2GR1%�ޚꊹ��W.;��%�a�C�Y�QV�����QcX�:E�bp����QN���2�6"P=1�^Y�a^�׎Wi�+*�\��Ts��)Vm�~�O����α��w ���t�;pfb����6�n�pS�4�b�Y2r�Q�{�J��f���x<��v�B��-����u*к&�u��2l�̗7�<p�1c��Vo�;Z��/���[,|U� ��H����6��o=Րc�8|YLu-��^�X�]Y�n��򪾪�9�g���y[��ˮ=�H�v�ʨqE��3�Qt#62�;+��F�%z��ǋ��#5H ��gb�KQ�!��r���݆}Za�2�(xVf�%�u��8�A��P��'J4I�Y�e6�Z���w�pp�*�X��aN.���;b���v��Q�6y�ԣ^\�����=R��f�+5�G\mT��Sl��W2Wx0Z�m����Eߜ��{��F�K�:fk���:e��)�-:'Mx��d���{��H�^p�dm�����,y���lc���W�4�jeG� /�GJ-K �G���s,���Z�'�r������l��Sy�a�0���re"�nM�:b�����D�����*�`c'g���L]!W�3���>�wO���&���j���{�3�:]s�p�kwUE�N޽�7"B�M-�z4]��9��]A��B��� ��sH�k*�6F8B�x��ͷO;2�U}u��nE(�C26T��^�N�1�V/��\�%V�K;E
����-�h(�O�vQ�a�t��r���=�|?A�{`�28�v��:_���X��9ڬ�x�����淋��N3؃����m�5��lu��T��qB�;�q;u؍�ؼ��H�A��E����s�A�y;VVv�͠��DAp.�wg\���d�%�ʓ� ���9�����#z�G��Q!��v��g�[>�5Vs��<�J�..x��'����&���kۢXOj�O#y����Oc�,�F8gN�WA
j�����F�.����0�CQC9r���
�%׮Z�8�+�(�ol+�+zE���=�H��*�Ia[���dv,�sQ`l�Q�2�vLJ;b��#~�*"��#2]yZQ�I��Lj��z+]�M���[�ݩ`k�uj��F�d kæR��$H[C�]P��r�,r�I��Bz�&������}79k~ǻfR�F��\�0C$�6��4-uA&��dVW e���)ֶ�Ub��Z�g*ёG9��8k�d3BV�Ȭ���})p����y�&So�Z?p�/��n^�P�V�y��N���ca��0�_	�{��PK�',���ς�i!�#�?{�����b��c���D��8d�yr�dP�;.lt3�~*�a��0	�غ��'m.�s���-��_�%�>^��e�F4�*�vxJ�v|��O�S��< ۤ�F����t��\L�'� K�ݸ��ت��Ga\��Ct�
/����Oe\ߛ�)���+&��-'n�u���ή��^D���t�ar�N����)[�35X�F]�	� |��2e��L���Y=z;H+՘gR��ct�_I����;7:+���5d���<=��!\s�(�窙�B�B4/'./"tl�`�r�7�+����u�D�g�!�D���6֝�}<���L��^ݣ~�P�v��Gf�֛43k1SJ�oY�A��ͥ~v���gN�}<d���5�Qهقܘ�z��Kh7k��x�����W�@��H�)Fk�`d��+�3�{��Y��r�<���ٗb>R�w��<��u���3ˢ]K2)M(6�K$ײ8��42����å8��<��z���D�u��v�ڛ��Qa1*�Ü��s�8t7��-�X�DH��,�����h��~
ָ39���h��J5�;��/�mE����Q�%M�U`�R�(b�\X�e�
F�wcjv^E<O^�3�ǐ��,s�y����JiP�ԸVϼ���n���g\q�)�vwc�i-=ON�3�����p9B�'�vs�uE�^S ���#Ă4��t���vQK��=�����Rw `�	>OV�T9�z�_RW�`[�zm@5m�(6"+c�'X7��`���-���e	��Gk �CZ�FO�{ӔcW
}FZz!g(�X2ǄG�bux�y�X��z��W��kUҝ��zӓqEmȀ}JC���.�}�ĴX �}�n�^f���p��Էk��ע�8wR&ɠo+�q	��L]�S�W�_}_4�����OA�>��!��4"��ɄZަeƻ�2�mC�x(+��M�ލx�P=G�R�܂�R�;�%���K����^(�ٹ�sC���F��S�D�u���S�K����j�?T� 
�8>&7����p�7���	{@�ikZ�����VC�Nck�,�Ԅv:d�sЬ���[&��L�Y{L�l���El��y7a���(�;0˸�h.2��u�,�)7��6��^���ͩ2x{�p�',8���2��Ƚ8����������x�X\/���F:Fꉃٲ���M�x�L<:ak^�q�趟�cg9��N�"'m[���뎈�����Qtzطע`�Ѵ*#����ܪ=�+��LpzU���g�[�`_�����(\f.�]���n�W�u\�M�sm�"��8vn��}VP7�-���Zs&�s���f�9p�ՂV�����y%�=q�u,���viX'b�����R��y�	z�x̤\�3���J�W����e$� ��MVa<]Gӄ�p媝�u�j�1[]���܁�����9R̝�+g.*�V�JPX մy��Y]\�Wv����"��>6Vm��}�i��#]kz�Z�s�A���Ԗ�fw7�Gdw6�r�,�gV�v8������C��7��xz7�֩+w5���~R�a�ҧ��S=ή��x��di=S��SA���\�@U��O&��|��j����Qa��T9Y�b}�a�g\:�g������Lڌ����u�Q��L��1��X��!9���7�dX�J*��6��QcX�:E����g�۹,���4�u����|���}�$�2>lx��!O<�!Y��J�)��+����Osq���F���Pݼ�S5��I����ڥᎢ�})-���r�R�9��KS�Wf�k�]�q	��ζ��vT堉��h���R�k�B����|MY�Q��d+�ÝXE�zm�dy~X���S��J] %W �Oy�Sk�㿛����x?�#��	�r�{��V�Vt��ʰjY��⬱�g���B�Ph8dvE��g�� �Gf�&D�/�B�-	��.q���)�q�C�����@�RҘq�Ӣt�F�DI�i�򣞭6�X�e	��Gǚ��sGY�5�I��*�g*�Il'�ba�QjY/)2����o�]t!X��하�I��d�.	b�G-���M�<t7�{��tE!]���e�#PWB��Xf�Ws��}��U*M�M=�odsmZ�oS��d7`\���k���	��g*]���f-���VU��g'��xʲM��ph<W�orv~���F���{j٫%��<��3�a}.R����1�*�t�TLHܤI\�0�ucB�*P���d�]&0z��5���cl�U�7�x��Q���20��tN��͞���m-��fo�	��Ƨ�5j���B���,��sH�}YT��1��d�ftRt�:�vv�(�B��\Ey�F�Zwc}\Z�+�:�Sa�幘�VRei��=z���wH�*���v:.}�$r�F�]=�p�=�[>�5V[�Ru>��̱x�Vݚ�k$�oR�3<a\��l�M�)��������gzgpWA�]D	������ݺ˻��������{*�p�A�RE��U{aV�Bl�	�nc����\���k�W0�Κ�
!}2�vzbQ�.�p�4c�Fd"�^V�gU:Ő1Ěӭ�������bw�0X-�޹'z��@"�ᐁ脣7�$-�u�ߥ�ȱQ슷F�;��lK�{�m��#T|��lWj�k)�(��(�O@�s�����*�/�Wfv�6ְA�f�OZ�R�X��(v����ܸ�_7F�6���|C�jQ�ȍbB�2:n�Rk�"��ns�9D�|��Y:뻱�ٝ�9hSx����f�9u֒o�b���Nݰ��m�j�tv��N����p�ͤ�e��a,��f��x =�W���gsYٱ��l�ł%�=��[K"�ԩ�Ò�R!� ]>�:Lm�G�`�.���7��w
2ݚ
��q�[���K��f��JC�J˾0\8�ZK������tpb���E��%,V)y/,k��:�Y.l�w��]�l70FA9{�B-ZQF���n��ռN]�`���D�
�E���R�]�]����S��E(%l�o󸝚�#��k�+`�avU��eF@xBVE�2�n
�p��u-\0p�%{J�V_��l�NrF��ɷ^�X�D���(�Zv�¤�M��+6%�z/n�E�`d�#�Z������IU���������R�7�v��k���hA�e�AϽ�f�U��Ճ}icٮ���l�y�*��V������TB�,�� ����Ѧ�H�.�E�y5\��218��t�&`u��0ΊSN���428��42�;}Ҝv�<uǧ�����kz��5:�j��E����kD�ũ�J' ��dWKpM�����r�
�D��&�YB�*��|�9׋X�I���껦4`�#}�wSz�f2�W��<x'm�Q��<��4�D�#�F{|M�9�j�ى������7P���:�ۺ�O�ۡ]��A$x:��U�:p��A�mL+�_)�Tꏜ�ngE�b����U}���Ղ�o[܇����������V��Q����U�ƭK��Rˋ��e�������W�-gM�,�$����G=�Kޜ�,�ɫ��V��8:e�B��������o�OTCu>y7�1�+T�5}�̈́�r���<����fz߄��J��P��q5�B����9j#/�Y�@_K��J�w�Y�ަlS��&ۮ+#=�N��kʀh[u
��&�s/EĊ넢:vqJ�x�%d9ȑL��5d�B=�8&kz��S�y4pS��x()S��8S����ks|U�C��di)yp��K�!�9&��/6o��ߋ��H�r����7D�i���X�۷�
�dB���B󙶖
�H�L��2v! �`�90�f�{3���,�^�����rd�~��A�!�UD#b�A�2�;�GU�2�xe�3y�v]Z����y���w�u��ՅLW�\ k�{��;A͚,�)7߮eŞ����V�\��a����I(Ԟ7㵧���r�%>�(*� !�W���vv-#L��X �db�
c��Z\!ǉ�O�/T�	��L�v��b�E�r��;����q�ׂ�ꇵh���u-y˂SF�N��Z���Ŷ6N��a���V-;YY���A�=Y$zoU@��*k�nuc�b����\�iଛ��:���M'x�s*LrՆ�k�W���R3�)��bv�K)��LQ�� uR��x.�u&n��ϋ.�QT
��v'�D�9���B>��ެ��B��m�\��.m7X;{s���H�����g`�i̵�a!�ϭ��7`2e�P߯���3��ERv[��l�w���&F��k�Hi7]�9��̛X�c�_u8P���f����E�®������WBM5v�bM�v���C�GN��Ě�˷{*�����r펥����͗��7}L>;���e
g�g������1�}{n���}ܢ�k۬}'u�M�)ۭ���ÿm����$d���q7L�u��\,�q\����}�����hޤ� &i���i	���zh8'h ��k���c����۫8)Ez��t64̵�3@V��˕�/�=�p�Bpa*jg*ʖbe��v��f���Ha�hk��8���G�n�g#�L��w-�`�WD�Z��1�u��p�k��cs���,ÝumG�d�Of�#�ٜ�u�����|3�LB��O0pY�!���Ҏvb¤���q�J�knd���)3����`�t��h��su�FR��s����1���hf�2n�3M	�yo6S[e����>��JGx��e�=[��Ԁ]*�0�c��]8Q�Uc����8�����!xw1M"T�S7w���r&�r��*�$����}5E�+�� X�c�`PA{�f��Uu$��s�OR��;O���]����t.k[�XU6m]�9[>��$^�c.�D�V�&͠Rɖ�.��DFAL�юJF�ձ��y������op\z�L|�mj�s���idh�7�'�����n,�
#d\��q�QZ��u�ܗ���ɴ��wT�2��K�aЅut��Qe1a���$��%zo.P�IoH��blD�Q�dq�sj#]ZX���:B�S���]Q:J�f���F�v�E��yǯ�k1<�.���P�Zj�J6�y�n'������:�|�	x�x������%�՗�af�y�;&nT��m,�6E������^���{�g�:Եc����R�<��;�;�����|�;y��y��E�����|I����[@;���u�{�5�؈�>�2�]���ubӂ�%̚ʾooV��7z+U����c�n[������N��S$=]ve���I��H����/�h�2Cb��[�	a�J���T�n��L�͏f���s�Wz�,z�ٵ�.()VW;F�evqY9���XC��<Z�v��4�ttrk��hCvȩt�YM���ێԌ�sf9�1�7��L�o�=�3�}���m���h�)DU��UUJXՂآ��LV��5�qemm�J����Q�ZZ������,�im��҈���m[Fʩm�,(�[iKj����T���[-�U��ZR�J+��J�hX�S�(5��-JQƉKF���h�pf�9B�YZ[mh�T��mmA�V���� �EQf-�im�*)UEbƭmm���h֥U�&GR��*UR�5K��DV��ˆ8����E�X�1V�QKqnH�B�8��+
YE�U* �Քch���D�
Ԣ���0P��)Yh�l0ʬU��Q����K1��E-X�-m�jPciTU
�U����-lU���ej����Em��.18�J��6��e�j�(ѥ�V�TX6�Q����Um�h�J�1�T[@���q���-���B�έ�c�`\:�:8Nt��1X�H�l>��ӳS�;����`�޼��qWꊰ�����{����5�v��o ����N^�
�2���Ƒ#X�6ո��r�&�a���{LC�	C	�\g��Nq�骖}U�+ӈ�����>"��HTu�������)�6��;�	�'�^����,��ǱٯG�ٮu�S��(�s\BU�����{����z"#>lN�7��=��ת�9�o=U��]�Y��vy�Æ��o���:�c:Qq�wnKW��i��'ٳ�Σ��*�M�ˡ��/#]�;����8��OT����bF�O!��؍�٥G5oj]�Q��q`e"�'�ͅ.��b}��3�w��÷tw9�6�+u����r�����4�d�S/�{�+�)B��ͅ�X�:E�X�=~o-��0#���֗r���d��e(əgl
UEX�p
�w>E!Y�ҧ�h�8��3p�3<�b|������q���p��B���;Q."�k�o
�]Fly�T�[�kwu����N������RF�"�KQ�"Y�*#��Y�x����LaPݶ��'���X|��k92q�v�(.M�~˾��|n��5�z螾U5]
�H�rf`�is��Z��<��~^�캈�b{�3��b�ʎ�����p�HoWw�5+vc��͕�i���wT@��;��Ȍ����ţ��[F���:���^g�bg�pt79@���J] %q�
T���R=��U�w��^W}���x����}�މI��A�a]�^ފ\w�U�"�R�u<6��#�`��{jte\�G��=|�̻m�e�~��d8��c��3^�>����)�/��P�k�Q�d�G#[�9�b�ߧ;�H��N�c��]�y;�F���=�B��QjQ�������|��o����.k��&�A��+�_K�*�;~%^c���9��+��
Ҙ�5��/��=�a��cb�gX��"�@�G&pႍ`2��[ڲ���p5$y�C�V�cٓ���l=[�l%�H̆�N��,m��X�n��ً���7����n�^�RMk�u8���5������r�0��e�Px���*��-���G�`�-s��uWE�v��JҮ�:�ZYCjGg:G����6]=�p�=����ګ�6�;��JM���ϰ��Kp�w��������ޤI�q�#�q@����
��bYތ���m�X#�c[J����2��͒+�D����P+X�o)D�:���B
����lS��f�w���+kT\z�M��B=��ֈ���3�_'3%��Π`+R�4H��3S֪X�mn�L�˻�k9���W�NAPxʾ?���������䟰*G��T�0�����.i��*�W-D�!d^B*��b ���1�(Qb��ײxN���$j�VYQD tt�Q�&%��P�8Q1�#/%TyV�j;�5ܒN��f�ۣ���O.������W�24:e(�D��u�:�g��a�۽T8�35�|9�Yq����F�j�k:��%��5k�	4�"��
�=λaA���9���%]�c���,�����Em��i�SE��aDз-rY�E#)������g��+��pu��N'Xx=��.Fp�g���N��.�3�ڷ���;�J��2���}�}��P�K����o�ōqx���t�f�]�l70F2;��+-3���q���M�vRJ	�z��\}yvȯ�^�6d3^�;15��:'���C���On�qT��'Q�$�rNP�XxVTdt:�Y�y���/3�pr���2#y��ƞ{��'eh��U��G^�>�c�b��"C��o�i�Rs�����k®��ġ�V����+`kj����.�e�C�LWv��U�%r���x~ٷ;����dWi���xNί��~93��{/�he�p�ŧN's��T��Wa�4*��whYO0��OD���ZHV��^��ԫ{eCH5D��;�t���<�����}O2��:��
_{��V���z�eaD\Ə�H�`ّ���Zݦz!�8^ƙ=�6 ��^�.�u�V߾�OfP����HJݖ*�����Hc��-F��y�������:�6Y��O��=�=�:�˜�p�����tO+y�#Ꮣ�p�OxdqU�SC/ڝ��Jq��ݛ��P�~���e���u1x���� �f�ݐ��f�#σ�j���nD���{ޱ�2�){j��^C4Q�a^b"QzY�LoJ�fh:-K��(e��D���l%���q��4�)[|sP��9�Y�P*���.�$WY���~�{���$Z��.���JǴ�4��6��Q�G(�rNt1�)�0�0�/��b}q9Aڬs^4��e!�}�O�գҡ�3�p���'��+#5��5�@1#y���܌Vg$�Բ�aAb ����B#]�(���"��3��M�u��y[O��'sw�/���68s	��5�|�
��r�h�,�z���b0�]���9�t;������K�����2%G#{g=�NpY��x�Ɨfn��ڹ|u;������8���A]����B�e0��;9��v��::���8��αhw]�ٙ�zhB_w=4�(�j���a�WCZM���K�E�����N���*�W3�P���[��� x�m�A]k�"�p�NQH���\D
�҈��>�v����eU�}�/U�c�(��{��[�fP˗��pT����+&�����u-GVU3��^�.�2z��[�6*�19���-�!��<fk)�����<����(�g)6k҆���������7�� �x���#
׫�f�l��� �^���)���VC;���^}�tl8�0����t�|H�ǣ�-���p�'�sg�8��a��ݹ`��7X����XJu�D`+cN���p��3�2du�X�z�3;~���1���1�=ε��Q�T�N@9�.�)#&�Tce�ao�*��T}p4�|$5�W�كl��P,�ٙF���e����͜zOC�x�����4ӡ���O�t<�r*�5R�\0c�\���>a������L�/�6z��Ϗg_oYz�y�U�.���K���j��;�wP��独ߎ�l��p��ߠFj)�_�OV<��x���P�FJ,���B��z��6۶u�y�S7��۠�EI�)�F�w8��K4'(gu����E7�=/�*�n���h�����|��
ó��ϭ�؍l��f�q�jĈI�q>s�3�M�k"����=aXf�9N`�B�P����;;{��MwuͶKީ0s��	]X���{[��� =��Ƽ��o
��bN��T�
�2�ǹ¸ѐ�U��o���q�K���涡�c�d�M�fο}0˓�e�/L�;cԪ��2:�T)瓀�T�Ͱ�ԩ�#Hu��D<��ۛ��b�K`�ݩcX�*�+��qQ��?\��s<E��=q��.��U���r�z�;UGen�ځe��O`�\�q�t"i#]~u-G`�,�\��Cn������=S͊'ot��t:�FW����hGt�Sf�
T�ߥ]��q�
{��9M�ӎۮ÷�w�w����2��7%��6+�\��J4wMJ5�⬱��=B]�,؅f��p��F�������l�SQ�mK�Ӵ2�ñ�����ٙ��}��P)D8���t�uP���]ղ%|e{�z�^�K��(��xu�����Y�+�Q~ə��(*}��IL8Ȁ��n�N�5�w���[��t��6ǆY6}>��3�0��)W�S(�n՛���*z���㖭�W���Y$?'���51����o�ۍ�7C�^lAh��ճ�{��)�ג/m��-�j�� }�r�Cy{r9��J'_<2r�^̱����f�28��v�k�`��rS772��3,M�Ì4���B��]NۚA�R����}�	7�qf7��u��o)US\
+)oAԳ���Z�HFvn�UuUܲ�/� ���u^⶯v����D�=�pl=������`�~}�e9�1����W�|����#�96��r:4^�Ϻ�P>��'��t��<Yq犙*p�F��Wb�x�9JΔ��0JU(h޽ְN�]36 :��P�ܢyU#���s�Y������Uw��h��߼�m�3u1i��ǰ�yfv\[��b�Q3],�g�F8�q^+`*�T�3X�w�s纖�Wd+pg�-F����4��La�ë+��{]�\�hb��,d"���N��:�{�'������&%�O!��AL��MK��dk��Kˉw�¯u���j�$E�N�Qִ�3o6x��'�<�岵�;ׯ2ᐁ�t�Q�"Bں�w{�s���;'�n>Rw,0xvK�Ϧ�QT�[5��\�0C$�6��4-uA%���[Ê�S�ڶf��v�Z(d�xd:�lX�(�g�Y�^��J�Y���ÀK�Hߋ��n*��Ș���{;�<g��6�U�xZ���Ӊ��^���j���+�0S��#٩�������˽vggW
n�M��i�*(3sO�]�$��S�Z��	�u���������70�h�B�T�R��ZxzH0E�4��)��OXκCn�����K���R
2��m
�j���£n�.�B߹�R�q4�*t�vYI�%I���ﾨ
��.~z�`�Gђ_�4�����R�p�E��/T��X������C2F�O��������R�,��z{.��\�Cz�Y�x��*��P+<,]����R�H��J�	g���l�'<{A�yS��2�5�I��h=eF@aWG7*��B�B!���<�j�_%��p��������ݒ�����<Ӷk��-L>���J���.���ewG����<pCmp��6+05�w��?6�0`u�Z��f`�Q�L������y���"3ڭ�s$�	����(��~ݤig_��}r�l����27��V�k5d_E��/$�#��V�L�:)M8*4�O�*�)���}��`;�<ǥut�����
��˘��6Y�4��=q`)�J&b���n	��[���C��B.F�OF�7�|�)^�1X]��*|�Qg3��",)�3�ڎj���nP����M�y�>�sKS�Q�%CTˠ�(�J�㚄����Y瞚�Ѕjm��Qnd��o��{�k/y*r�(�T`���yJ��fl�7�ӄB�5�F�_Z��y�*��)�=�Q⻸=�+ԝ���KX�X$�vT[3"���s�6E��7�-���^�s!m8�W>/y/�ǵvr��,�nb���	�(9���<��okg��ﾡ䬫�Ս�*�����,��}���9�X�Q�s�uE��d����#�b�ֶ=F�A�	�J�Z��5z(U�S2�x���qY5���Z�1Uq�k7\�l��GA�Y[
"x�]��@pً���~�=�iPm��������)���k�A�՗ е�G�������Q��H�̈�#Gd���on��Ԇ�:��Z�,vI��t6��w-�4�/-a<CB����V��^��q�<���
�o��c���O����:�pg�����k�u�S~8�U���l����^6=܈�S�����y6����y�8���J�P�;r�X�|��{�����s4u��:5�&N2�xl��Z�7�@p�P�`�>6'ne�7�":����e�喭��(�.Mƣz�tT3���a�nT�{�D�"v���v?��/3/w	��ɉzL���c�h�yʪ��
�����KX*Վu�Kgz���I�U�H�Gr�^�"��䇟1j*��V E�mfT#�g�ʃ5����4��)����FP{�F�r��6�yJ�i��{9:��U�rt��/:W�=ZҬ�ι-�M�(�K{�jruDV�\T-��D�f����[����<&3��{{���y=W���(�U�����F�ux�co����x}�}L	ݫ<�A�7�z�z��m�O`=R�e�ǻ{���z�'M��z�ϘyF��M�\�}���e3�;���[S�E�"�.��.��Oc�<�{��`�a<qc�4����n����-�v�����6$H:�,���4�fKc�>�n��	�S9����C�oO�'��]�Q�R�t11%��#���Y՚�Y=P�jk�.8E@����h�Ml���}���֞_
mܖ�_B��v�*��du�*9�����
�kb,U���U�֧sw�\����͍b}Վ��ܸ��t��*^�.g�-��a�j{~OҞ<彫k�q��lG(�v����+��
�� ������Z����(�S��gչ�WH���Rw-(x<��C=e��<<+��r��t�h�� )S�gAH���q`��ޡQ̂߂|N���F���qŋs�NY��a�⬱��=��DO�z�.�jأ37k$צ��w��&+��3�W��A��ۓ*`�q�<5ͫS��r��c�i�eѹ�:�O�q�۲�������^o:\Z�
,h��������=RwQ:��L�:�v�^�Q<���w�M�Zv3�غ;4#(�y8����DT7�҉�3�ԳZ$�v�Ḣ{;~��Gۜs�#;0ӀLB�ޫ�Z&^f!!�T�7`���m�em*r�w5���5��wJǸK�9ͩy���t�0����,�W,v��k�}��z�N�=J���tu+t���m]�a��zq<�Ҹ�%��_0�'wf%a^��m�Ǻ�-�M����Z����vq���;�����kk*h�V�]:�I��p���7rs���)éh�6�w%�i���{[�]�N�Y�z�,��`��L����j�{�}�[�ω�Fɶ҉)�/R��J�=u�%
8����;	���ڱ�
���H�ĵb����X��^"�����%Zjd�|K��h�t
���]���Ѽ�ͬ75�Ɠ&��X`���\k�#6���7׉�:�oL�n�܍`l�9�����-��w�U���(%�:l��R��j����ښەܙl�)��X�JT��Wgb���Ahvc��K�hmlt�
��F$6�I%}�0���J��OU��f���;f��)�=���W3D�(�Z�������9�w<	�5h1�n7o,�r�H�.�UѼ��˾�<M��aq��Xҵ�)A�p*`c��WS=e.��L��I�ns�B����evժ��P�[�a��=�ouV�WGe0�Pt�pn]^�7[u��y�,���η�u(�P�

΁�7�ێ��;�Q�X�<%s��ǥ���7�����x�֣R�Y�ei��gR��\+5�������-ࡎ������V0{�M3z5Bbq��ݲg9̮��3k��>�Q��A�vr��4lo^p�!b�ʒ5	�x�%��I��R���X�!��:�w���=]��wgiW��Ӝ�p����8i v�:D�K���l�Y��]��¼�x�r�H��W��ӛ�����@7w��HJ��+�-����WWV���c;�;��e&�F�	4��Q��8�n�hP�|�r��\�fU_q�st[Ow�L�0�s���gm�t7 Y73�� �g_<Գl�\�ŵ&�9�X�Jٷ���5�.m2����\�P1�kxQ�Wi�ŦN��9LL|��}/�������������Υy	[ �����wn�S��Z�]O���Vf5ua�Q�+��/�����{��r�6��î�+}�On*r�]��9q�K��Ѧ�.���X���ة�sQ&�Z�%97̫��'S�����N�e^8z�N�.}{2h��V��Y�5�G�L��ͭl�o:�3��s�Nc�G��a�����euk�)��*e�H�i�ݒ�rZ��v�>�h@j�	��a*T�[E(,k
�cŢ#jYX�k
Z��p�*T�K��*\S�.Z�� ��U�ծ
5-�A��iiTKJ5�h6�Z�j��*��m�akD�TQ
��R��e1������5���-T+*�"\8��qB�X-h1"
T��Qb�[jT��X�jTFR�¥��[IY[j�Q�ڍ�EUFҩ��EDX�0�"Ե���E%Kl�F�QPU
�V[Z�ѩQ�EQ)h�U���(�Zi[J��X�b	Dm���#+F[R��kJ�((��X�*%�Х�B�*�k*,Z��Ua)���bZ6�(���1�&)qlEF#m�(��h�*�(��(��b�X�+(�iV��1(��R(��[cP���Q-�l���"EVUUQbZ���-b�#�Q*-��VЪ#mF���V���h�*�����db�mPQQ}��|������ɝ8�{��O�W��-m+���h�t9�h2u����Q��緹�"-V���Їs?Ͼ�����u�xW,n�HY�T���P����
��q�X�l���>��(JaƋN�Ҳ����npgZy��)���<����]q��9mp�Rd��Z��Z�y�TW��
H�$�ˍ��z�⫘�E�\�/w����r1(u�g҆�2����*�r�o�����k��Y�:�(w��c��NQ0��$��짦051�A�u�o(�c(u���
ŉH���VΌ�6q�م�2;n��ݮl�+�僝o0,:�n�ߞ������k
7���b���3�RyFȮ���%瞓"�\%����&��9�#|�X��/�ZӃ�1+]�7)V������kX���-e�*�C���/9��r��p��V	]!�g8�j�*�oe�������H��.�;���zjw^j�̢��<�J�(9�F�3��=�q�#y���Ob�C��.T���`����}�[�|v���MR�Í�VT8�w�]��;�RE�Hu��2�B�^~��M;�O��]�-�"�	{Ӄ����uL���t�Q�J��)I�T���Fe[^l��6�9T�}{tr���5y=�E�'C(�@8�z�83q�N��^3Z$Fpo��\��qy�N��p�`4�-��m�eI+s�9ȩ���M�9ק��V
pV'�=]BQ���vr7�k:g<�ٕ֨db΄i+���J�$sV��w�����w��\�3���^V�n��<X<�lk�w���#@p�@�L��D��O.�"Ch����Q��\���(�`�g�Y�����f���fC$�3�0ӵ� �_o��0�o5��4
C��CȠ-�B���p���p�l�hJ�Y��7r^
D��)x��V��vwmnj����TlE��dd���rِ��f��/zpK��f���+� (y�e#S�?�1�}�X؛�uz~�L؎�I��F�����l�c]E㊯�/c�Zp���l���'�L���2��=����S�*n`��/m%&)��j.;WT��9�̆y�є��/'���T�ļ�1!H��h�,�\����<�YQ�%d90��T��;w%���]��Ӄy9qeؚ�`���ݓ~Q��G9$h{{b��֝��':oN�+�����
�ڌ�X��:�ڽ�o����񼁕dq��gqK�Y�������jЀ�}Y��=n�|�'6 ����`�t�C9W�l:B�-uT��:���o�A��*�z�)�7��k��x�R)�L�bw��N�r*��Mh��f�8���������Ŭ��_���ס.��R����z'�/c�u���:c3�B�VC�w���q(��kB�\p4����q���U���΍�*gҕ� :�In���h*sP��xxۗ�Օo\�*?�Q����W[xxŚV�^����U���2�jvm'ƽ���_��Lq����ש�=~��0���ˋ�.�W��t��p4ڮZ��H��<p�ǇVہ_l�H��hm���Fj�)Y��y|*}�q�<>�sW']�M�6K�wPj.)�w�eռ�oLBQ�CH�
F�k�m��j��9g�M@d�S\
�QpL�6��2�ʷ�h�B�����Db�^w��f�����r�b9F�s�uE�^S5��&�fR[�q��Ie�&�T>$�j�C�T�՟$�MZ=+ץ����M�X~��_ �h����B�ut��S/!�� ��PI,���DH�2�r!͜��.������j{�����yy�J��ǟ�t3޺u�zn q�E�U+���ٔ	tג�^l��j.�d��'���Q2kGH��y�@w��,X�q$/:i`�t��U3�2v!�+U���ӗ�����kA�crvc��͉(�q�Pl)�.lW�^��Z>ӏw�0�9����y��-R��bYF;�K��p��C�C�MVfZy��3:�pI9�2�wP �JMG,�d�dJ���(�hx���ܚ�I�)ŬZS'l�N�M.�>VV�C���0J�_7�z�g
3-<����l��5eˢ5w�O���{�N�*'o��6~w���f�np���E�P=p�H��:9�;A͚,�)7�+N��K�y;J�
�aT���u���}j��> %.���x����v,5pt��t�T�v�o��v���E��0��Rn5�ד���^�����`�W�4w'O�mk]�(yF;��ז�>3���}��pN��+��~��U�ִ�7�;�A���e+umdS\�\��N�Nڬ�%�O����0tՂW���쥂�x�c���sS@j��[�ǦuF�W�os��Oet�<U7Tr�:`_��}ӡ�����]M��yp��[�'<��{�c���nj鵂5��߳g���EҗP�C�g|ڧ�����6�:&1�S�>zS��`����W�i�
�T�;Т+��FJ,���B��~�'ٶ�u�Q[���V�:<�sH���8ҦmFzbJ;~��:���G8YR����l(g�o-
�25MD���<#O��¬7�ͅ6�KK-FL�;b�QW2:�W�O<�!^�tn�s��d�k�cG���%]ȕ
9ڌs]-M�2� g���zU��d���Yr�qC��ض韭���uYQ0�S\�et9�u)J�Pg����7{��\���ĵ7�.���P��)w�ٔ�t���ڷ(t��ޗ|��+r"�*6��  �ͭ��^k������4p�����ܸ�
�,�zD�dv.�ӵ�ص�}B��v�Q��t�����Flk���S�Y8`!�M��\%�k�P��C�����S+J�s���@��j�P�Yg�<+��)��6�� ���S7�hf���3Y��5L]��uC�(b2͢p�g��2�?�|\�>|�,׽աB��;/fk[��[����5�pe���r\����wʱ$��j�-��OO��r�/8��~�~�����C�Ѯ"$�(j�u\|6�#���\~X߲��L�ߟ�(,Œ&�������{7=�Uc��)5�g�:^V$��8Ԭ�@e��0��k��oÄ����(-��=�3'em�}��*�ހ)�w[��ا��*�ۍ�7�͊L��rxK�Δ;��� /!�S�۝����fM�rM�ƪ{�7c�=mb�E�tP��ޜ{sQ��^�JT����Uh6F(b�x��1g=�ˈ�<T�ܥZwc}\H����,T��ti���6�zv:��h�lI��6�T��Q����D�+wGC�g�՜U�.�),�˄���.�m���{4˺
��{��^.��b�2�Q����ӣ#��ݺ�wֲ���g*�-c9�3B;��ҩ�:nb<�
1�Y���Tk1b�����&]�<�xɦ���Jm��ޙ�3��5�P����r�Ga��Ng����r���Wl8���bQ�7Wxl>�r{ }EE�s��_�Q3��d�<R1���
�^�=S4�,�'�����Y�BZc��l������Ss͇VVz\�=�tJ�.Z�41HXp޼�+-#�������N׾�B ���Kޜ�1#U�VY�B��7�+��R+�J��� ����n��c�5��fTB��-��T/+J6)>X0.��$�k��F�d k�2�jk��8�1A��N}�zT��^xτ^]fQ�᷉�w�6��Z���N�Fd2J3n�f�-��rO�����ieZ�K
;�kl��W?��a�˅�>m�����˶���ʜ�k��,���A��X.�GIʦ�
�e
�j���qiŃ�Ξ\����Gp�R���M����P�Z �a�e<|�ZJ�D�����WIp��bƸ�qS��ʳ��ҘS�`�,�[yպ�i�~.�a��0T�ʛ� yI(y1OVQq��h�3���\�h�8x\��5�̔*��>ƹ}}�F�^<3v����x�@����V���"˹��EŨ��x�a�s�����nt�&1Ys��l�T�/Go�-�Y�%�Wj�@�x�Θ�usj����ԑ�c Y�;�E�p	)ٗ���tS�����U_U,RhY�۾��X�U���xU�����(�\���ʰ��eF@x
�-єS63W�m-#�9X�;�;Vo���J�q`��������6a{|�>{{t��`�^J��d�$�
�7�Oy�&�`�nMq{T΁�2��H���� n*q�3ђΝ*��C�K��=���3{���SӚ��c5O�����r�n�7��!@d�Q^�T2�J*"	G�Z��ӧ6T}s�ZC�M�x�EZJ}li�+��iVׂ����\�xg�Y!��O.�U[���W�{�r�S�7k�<���Ӫ���x�7�z���)(���f�[�m�'B�"Z;�9E��ڸ���dVR�jx�Kh+��Fj�)��e����E���^�q������Op�ڧ�rN_V'���mJ�΄\p�eґ��[|sP��89�<�j�ǧ)�.,�R��|J�%�pY�}░��H݋��
�F�^��e���f���QcX�Q�9�:��_���f�����s9�|<�=+�B�K��ֺ^{d��w���s5�J~ע�i����m0f���ᛨ�`��6�\@Gx��X�J�Zƕv�ɱs^��k\᭿x_�,)ln�ɗ����:�>���*,�:�WT��v��N��H����>�{F֐��'�e��M'��HVL�2t��=�밹l���L�����7�7��=zv��s�,kʀm�M�#�@�+��C�j�L����L��Fe�Hd[y$�V㝫��N[ɣ������AXח էPTE�:GrB��QP��&���/�y���;�9\���V�5�\�C�=H�r��S�EG�:�z2MeT�����c���˵��\��vt�+���I���Ɓ�C|���^8J�	�k��˛�s���orUUnK{�{Qk6y���8�M������^"*x�J���5��	{���(�dT_T�{*��.5=�Nk@����J�Ef�T3�.�ٱ���K��u
�<}W\G�'o^w��r����x�j&�WUE�����$3��x�u���kƖ6s�j��u��Y@-��p��_U�͞��������\��^����TP��P5���T�J���V�?1p�s8�cfH����`X[���S���
��>�Z��K:��$�@�3K�0�P�}��wf�����/�uG,s�����.�N�y=�����6�=s=hdKٺ����=SS`�l��x3�q�W��^:��w!2�N�Wm�2��OgcG۔��4�yn�_�3�]V���2�pw�&M䯹wh�b�uNNRN�W}�w��f=�7Fu4�j�.�I���oB�:�U������{t�]<�Qjn��"�?{��s�V���e{#�`��U�߳����.���t0�mS��yL�c���맚%�&�'�y���T��k[<Ӯ�Hg�Qr�,'�ʇ+#��'٭i2Nӕ��oQ�F���q�����Lڌ���O�B��]���=fU����4������Om��3w��1,�5	���fw%�a�Цe��UE_�G\
���"Wڶ�h�Q���z�Y�kƶS�4q��s~�'�^�w כ����Ӹ�����v�'�Z�	�2�4�`�Yܕi_�O\,,������T�޹N0�c�A�H�D[�j;d�wR&��B'3u��єe�9�[�ظs��+��Axx:���>.��0Y%Ǻ8������e�*�w�ܻ���/	�������Jpu����Ye�-�	�R��ӊ��׼NI8\;4C㢶�G�m�8^��]-x�Ėg��sw���1��ǈ���0=�;�6�dt`~j��:�Y�YQ���,��\,jQ,� ײ���31��x���ϋ�"�3E	���~����@+�z�Xb�+i���V���2�o���h�c�۰(Oh�pW>K;I^nE�ߓ�e�:G�np��*j�4�ή�7֏Q��ٓc���'`R�j�=Mܛ[�&.����/ǎ[Z�54�'����]a7�vi�T�N�uq����;�����Dd1�N�j�>���d��H�|pjl�m�z�A�ܞ�y��;T�݆�DySJ���'o`�6֫>��W�g�	���Z�IV��n�?�\�Ta�٣��?w�M���v��7w�ł���P�#��B�xki�ᔼ5|����|�_�S���j�6'C."��L��U�v+�f7�uj�U�欋�,'�,U��6�p�L�`�>����q�_�ܢ}ʩ.�ǲ�Ii�cO4XƳcQ�x�1�|}�]��;�Ϥ���r��yD�t�M\qHŌ�qo�_����TO�fw:W3|ҴK�,��w�<�:�B:�)�8�ueg��3�RJ�\�_F%sڜ��M�)�\�Tdp�2�Z����w�	{Ӄ����ue��)���Q�1(��VyVm�b귎�ܗ��j�X�*#"/FJ*�t���N�';���S�Bj{'��p�
&��F&_A�Q��$=��P�8WQ�ͦ}Y����l�
u�3#���L��ܢw'�,X��Q\���18�C�]�U�ʕ2��5mN�9�ɗ�//:��/*=Q=�)C/[���G�QKuw`"Ӳ�)g_q-#�fa�
��Nd[���m�U^pW��,e�ӂX!441�#�q�p�*���m˕�-QW)�eG2p��o�r(�����.���F���*h����-�&z�U&i)N�7���6)�Kj��������I$�2�������\/7���T�@�ݝ����炊r�7*�g�gϸ����oqn[W�Um_hÊ��V
!ځ�U�] ��\;F�vP�-nЛ�Mz<��ܫ<ܾ��c�-��\�r��z�\nZz��r�'�'!V6��ej�=�)J�\�T0���hP�}Lw^<�]54:ٚ2�$�]���;���0��;��FV���V"Nus�ȫnX�ԣ�)�ޏ���fB��5u�K�Uܺĵ�.��U�'{��-j�օj�Sf6��6��mm�ZK	p�]�m��b^����3QPs��4�5Vu��ɻX����ڥ�1���QL��Q`�m���n�;H�mQ�Ԙ�N�n������9����[t���N̈́�����rv��dv+���Y}��.Le���Z*.��.���
�3Z5oJ�iݥ'ܒ��.�@�������Twsĺ-}
|��܅�d�q-ձ��V��V�)q۶ʣ���ƻz�Eg�U�8f)p\[�a��XE�t(�|i��z�����:+�(�z�n����F�[���"�{��n'������L�u�ָʓ�]$�#(�YG+��"8��	�3j�3�v�����	�xs��3"�B�3\R�D<�b���}�mW�Fej5F1�eNZ��fu�c����sl>�J���VRtJ{�f��c���Y�f�cə���͎��Ȼ����]`��}�}}���Xʼ2�sSFh�fH�h��em(�]��A�X�1��.�h}�#�OY�2�w`�ޕ|9O�5ɜ��	�<��b��-���@�cj��n�%�[d���*�Ϯ�ÔOHc� N׈�J��wW�����	<M��#{[���(��i[5�v�3i�\��wn�^���}/W0ơ\֞�q�)�o���O��:��u�f��wh�u��'�5J�K�ul���5iQI�u`�2N��	̽���Z��sQ�� 6���"�P�4M0G����5-p�
�!���L���kp-����.���aJ�)�n��e>Aժ����#*V4I�k��4Q�-���W}+]�wC�>O�c��~H���A���9�[��/r�N���E�H����d�=m=�U�%��n^�J˖�����i`�����b3�w)*�	ݼm�8��#W�.�/���z]��n�F͙�J�ou���^v�&j=����b��%��ʢ�,Q+R�����K�"AVT(��`����V0J�QUUZ�X�UIQkcXV6�T,Umc"0UUR1c�p����""+�dUm�al*��J�X�Z���[h��QEP���E�m��c"��V����X(*6���ԬH#J�P�R\\*(���T��"�(��Q�V���UUQX�DEb �-b��[TE�X�5+-�iZ"�Qb�������Q�(�#�X�)F������#b-Lb���QEb�b*(���*��ED��Ŋ�(ŕ�j(�ZX��U���m�*���iU�	b�
���cmQUUY-*�DPQUض0EUb
!mE�*�E�m,b�L8Db,Dp%QQUTX���mP`�E+*(2�֑QQEX�,TX��1���A"��lQ�QF6���,���(��T����Z�Klb��$PTFb��(���w������g�xG�bu^r��{s��5�\E{�j�ݎ��X��[$@��e�CwEb����\Փ����L��������{��h�?�=�$�P[b��|`s������Q��ڏ+�9���N���yWck�2�1��X������
����e6�U�p���u�-8��x{5Z�މ��=:Z�{��L�Ka�t�1A�݉�T�p�i!�#�zߞ�D�TX��������)�μݫW�:�KQ�]�U���,	�ر3s��IC�1OVQq��2�+����z�t�;-��t�V`X3�:�`J�l�(�C���ʰ¹���%dM'�Ve�&�&�2��Ug��uZl9hu-\2�aXz���@%q��&o���%0��edX�����}<2��M��+6%�z��62T!~#W�̍�N"��3Ѹ�8��yT��&[KW<��]�L�.��OsnM_���frb��ZY>�(;��+x'��C�E���ֈB�~{o�+�{���@������ʯj�%:�cO	^V�JG�)�~"W, M�}+VT��.wzq��6a�-���F�8�x�b��7�`�X'e-�r��U�t;��{���|B�3:�i��H@ͼ�FRq2Q�b�f�*4y���eht��E�Wy{Z؂��,ξ�̛'�u�zz�w
ޫvƳ��`9�Q�*��[�8�]N+�Up֫��]B��J��ٱq[�s���7#yQR)| Y�ع���~�N"��DO�mc�S�Խ�f�;�����^��uG� �u��W�6�5�U��UX(չQ�Rˋ�eה�(�J��P��89�<��j�3{A���:��t�u����
�Dk�!l_��\���)e��,�/��N(Z��V8\�]��iV��ia9��+��M��s�㮎�Z�y�;O���/3_�+��A8�W�������f{��9�/#5�Խ2�>�-4q#��	�B��v�ں�'��Q��C����5�_m��"�)�G=NG\[x(+^\V�AQ�H�	�׮A*�9{���į+a,��"0��s��0�m�A�
F��j(G)b�I���:i`r�����v���gsg���g��@u�]��9��G�Ĩ;�!�J�!����n���h�\����q��=Gs�MU���\��*�J�+	;|<�Pw�"Uo�us�	k�Ļs��{ݛ�X�G����|9�+���՟S>���*�dR��$��To|�A�<@U��!<,�1+����#�&�·��&��vV:��A�ɗ��5Յ,<�׷K��-k)ίZk̼�W�5�*�ff9sed"�/WG�r���g*盲L��*��t����[�'vl�y�9��;�����\����C�Qu �sJ'������깚㱓ԟ�Y�^�]�tl8�0��j7TL͙(ށz�x�l�0�Їgb!�Ù��r���;�aN�9,ע���`N��8��~rlPL�F�G*���.�1`̓㍛oT~�r���\�.�������]�F��(�U��>��6��)Ŝ;7"��ڰvxN���[Xd�U��l�~�E�N�����/�U>���x�'�4�����b0�b��A�Zî0����+� P"���J.6Q|��3��Yo��k��g��JnI���w�;.m��L_N.�� ֟.u¢�"A�"��(QyH�A>�o�]-��Վ�1��J�y_n)��U�:��n���Ι�&$��Gg�W�G8Z�jm9E��j��}/2���O��n5��cgPo-�
mܖ3�%��<������*�k��j`�l���2{�#+e�ˬ�E*|������wp7.!j]3�"Y��O����/b�a��/4�ދ8��P?�-�	��3`#T�<��Ny��c�A) ��C"��A{����*zw�7:�h2���۳��Wq�H�����1�ƞX՚�)Vw�Ѵs�m<�%v���-�=�Ƭ��Y�1c��[��3Fy���tR0v���!x���àZ(�S?h4d�l���Zc7�vnVr߷���43o�<y/kx��Κg���?�*Z1��x:��0Ϗ��!\&Q��L5�C�H����_�yB�ۧ��樝$�5��13�+@�b�����T��ݚ�m��熛�"�!�	ޯ-�3��gRa�^����^<+l�|6��g�;�+��N��N�ϷQ�pl\
궻���W����)��t�׆9d��uP��=���v({cf����V2w\���:��G��%n7}�|9]UA�AWϬ0[J,K������d��i!�a},��l��޼�G�o�~��,�j0���VoاLP蘐7)Ey���1�����+|ۍ�6P9���p�M�qէ&�Nʾ���F˘f�Ɏ9��,fΗC���kw�ݡ�sǬ5�б���ޱ�-0����������6ni�MeR���Ràr�%5�#r��������<\X֘��e���,��[��:�a�UA{B��Z�X+�j���ͤ��V �S�0��=o׫��|w�g�~Uw��x�Oc�*,ߜ�#�OW��Gp=�G���d��<���v`�5h��+���������2�{��vv,��簅�G�4.���>ݗ��Ե+�\κ+h�t�g�U���e��jF�a|
zU\�G�Qm��[�U��I��g��{@�:���1�&Z�\O.����Cy�>��ǑT�"f���%��B������f�G���p��`�%����:�B;�5Jc6YX��{=WD�Og;�G���j���59Q��,�<W[�
�A[�1y��čV��%@S2�q�]�VI1�SZ��\i��G�*"�9De��U��G�'���Ӯ	��k̂)�շxյ�r��Y��n�ur^×J�vE��+"��=�,����FV�f��\�%lQ�՝ffq���׋��p���&�A%��́!dU񐯥�l9G;"Y�ڏ+ֆ�=��~��;�����)Ӥ�	x)�v`��GDXT�ɏ#t̅��f��E�M�]��̞�󷳮��u�|��F�HWe:b�ئmL���z$y+���VU3������hse���{�;#.2vt���Wlߜ�F�⚼*n`��IC�1OPQq�Cn�WE��G/g���z�4�t��<m���_b��� V�����^U|�!^�p��Ve3��;�=ٔ���Z/-��"�-\2�aN� `��vM���#��'ޞ�S�w�e��w���ֺVdm]cƤqq�!G�)j�ő�~�q��u�c� �-v8�Q�%ؾ��ċN6}��k���>���]��gp��Z	A���^4.>g/�Cpv茼4�m�b�ne��t͗V���fe�uG:=�:��Fj�Q���܎hs��`��o�w��^@�9�nf
��4�ʽ�F�T!`d�q@�lϷ8��.��;7�Qx09�;Q�\r��4�xɧ��&�5Gz\D�,�d�G��E��ٺ�J����C��6S=�ϵ[í������)�O�f����������,ҵ�O��+��fP���:�v�w�[�[�=MM�jv�0)�l;s�x+��aŞ#M�R�er��V`:��o;�t���Y�;a�J	��N"�Q9m���S�:l��ae�()����V͆Җ�)�a���{m 2��Q��h҉�r����26{/N�f��Q�0��ƶ�E��	�f������zp2��s$vŊ���UtF(e�m2���*!�Z�Lp
�Ӊ��<��Y�}M�p��F�*e�㇒�T�՟(]#�dO8ف���M�ħgt�n��_�G��5��h%���/�Deq����;s�"�ښڪ��cU�`���1��o[7Ny���NG\7bB���A��#��M���T�2;��m��-�Κ��ĕ��S(݂�Zr�0�8VY3|V�W��(7~��F�T�����fW��^���f��^��y���Z7�Z.�:c覰e��O"������Y�O9է��ؖ�wEk2[��[�'�J�ՉWKi=4�uf�����]��8�;�N|�Di�Y�ق��Aה�W,�9d"G7u��4����_D�n��4�y,�5���a>K7|�J5�x�	��B|D�\1�TB'V;cEn�E��T�ov)e�s\M׷��h�{M�`us��DR�r��{)1@���2����9�E[����|�}�>z(�C5��ڞkóVS>?.��������,�f!��S�۔����[���ض����Ǆ��j���ć�ν�k2&m����F�|�.w�z�Ag	!^�I��y �is���>��+�@o��(����Z=o��.�@�z��ޜc��L��)DLnRF���7��Pt���]1F։�6�59��x��J��:E�*�ʾ�<�6S�����_:`[�O�v�����`��+Ψ3��E����RiLz��lS���gԪP��ϨA�LŃ��jR��RƜ;�]�Vb�'�/S�-gk3�޷y�M��qc���=�*�"�ĉ��"�(Q�e"� �S=���9�S����]E�i�(Ӣ\�D�u��2��uҜ:�����w���+pnJ�[$�Tq�'p�0;q%�x�Ӿ�G&du;ɥ��Q��ʽm:�sz}pZ�h�z�ҽ�V�4�>�[��f^V�
juw>�R�:�t=�'V�u]m�� g7^�*�q��쏂b}�m�:��3aͻ��9�6� ����L��2�ǹ¸�j�k�ݕ/�r���N�?j�f��Q`k�H�bp���ͅ6�K�Yj0L�;`R�*$X[{����knuS��R�z3�XqSY�ҧ�h�9T�k����P�-��b���{˽���O{$�VjJ�S*�k��7�.�f�F�-Oe:品����D��tZ�8�q�s��G�5���P;�ːP�7庌_^�3��e�h�Sf�R�o8�Va:�μY�|�^��3��{M����.��x;S�t鸆l�G��Ka���v�[Z�d�����Ъ�g+5��GdXmxn5t����[W�X���Ԯ͝km\sw�;��{�.��]�'D���J���:	Ygn2c�0.��oii�E[�_�<|�/'=�:��ٙ�΂�<�@l7J-K>����$��!�P���p�0��B��d-��q���y���m��aӛ�GqΘ�tLnJ$��^A�����SyQ�EL�3�4�5�3��DOt���n��Z�|3'<swGYat��l�{��;h����b�n5��t ��J����ՋcK���$�56C��.��C�eL�0������K�P� Uҡ�5;闥o-,�h�ᵝZ14f������{'r��ഔͷR(�1f��n��f�mYC6t���D�������i��l]t�܇��T'�u��آ����V�� �ىG��ʤ�����WK��}����o6G��;z�j<���+�N�b]\Z�)��@9�;�*��������_oh�f�	��;��};��.QaK����ہ��������TY�9Hż�k��Z���CruN��l5i���2�0��P+`.*^F1���:vº��Spë+%�3�N.�u+�r�)�}Y�nI��@-A\C�:�O�� _9�WVy̞�X��E�6ó��u�*Q���f1F?���T�����\E{>�FX�EW�+J6)>X0.��$�[�x4�qJӌ�o7���u�ӫٙ��D��.���+"�9G��>�Y���O��Uv�:��ӽ�|Dܗ޲5�8�u%��M��E�!U�6��֢���|��݊{�sgzM�z�����y�WSq������2)y�%%¢?p��O\�ӊ��ܩ���r��U�l]����!��*�(�]e�핣B�b�Y�"�T��g�]ބ��=r���Ǡ`N/�������Տ��z$s�ʊjmMD���"����T�����Drd3�lG��GKXW�k���$\�s;��*��sڷZ+⟄�W�T�R���*`�qL����J����VT���m�[;�[��iT��xt�R�dV9�sc��ઙ�70FM�؇UA�YQ͈BVE��O-i���yn�솷�i��݊P�>�����O�\
�$R�kø�$�m�����0w;r�{W�% �g�^����d@�]��i��g�p^N\^D��@��n��^��
1xd��w�o��
�/E�z��5F��;a�Rs�Ù��ri��/n��.GSYK½W�#��eq�/8u��Ò#�O�%�:kϧ����ۓV��6`�&*���Y>�����R�]���8�s!����=O�i!/��3��ً�f�����뭍<'��Ү��8�l�p�������4[��!z/�^�p�Y]SC,jv�3�8�x�*����
��vR�u�-��I['��]?�Z�3ID�T�3��j	��/l�9l����V��e��
�	s��u����y��A��G<�:캦���V)e��2�Hҍ����/zk��=������"��^�Tۍ!tXU;�4�V�q�V��1�w���<<�o�h|����
�:��هe�R��n���=�FX�7n�uU��%U�]�ܴ���ӉQ� �T�B���$�U����t��fGy�^Pϔ�q�-1��ӎ!�%�x�KUufs|4�x���y7{��������F�>e�4�[�֐3��s
�f�&��ᗜ��T���[�Ԯuf�J�-�g��H�nx�)k�G�ԍJ�FQxk�s��T�t�Uȣ��`v^���:��$^T��l�C�"���ی���lj�Uq��R�=�.�gK�]l׸E�N�J\7��Z��[�LV��ST�d�U�c�1�+���V$Dҭe'l�S�-���A��X���B�Y��.�,��)i;Έ��n�k�eV�b�.�R���K����8����eѷ���M� �Iw��X{�.=�Ѕ@�h��^����w�;���ޡw���
�T�Y���\ܾj��f�q�m�7Blb�t�":�;��G�se�n�_hl�"����e��4+k>V�W
h�^coPN�)��; ;����`�̾]q�&���ou���;��&��o��ԤE���$���|N%īc7w2�X�4ә���*���]��Z�̦��D�56-��yA��7Z�5
�q��v�c\��X��`s��u#��P�&���y���*<F��	r�a�,���lh�)v�M7ʚia��HBS蹍�/�흓B��ӆ�wءt��/�Jʴ�P�T�f���Y�����X��B��/��5W[���9��jb�gOD�=R
�vvl��	�� ��KHW�.|���|@��*�E����LD��v�p[����Q��b�Y����[�2V=ϞZ{���F�u�ߧI:��!����/�Wr+�R;�k�r��1�h��Nݻ1����9��0���R;�z���+F��qT X�p��̥��)����GZ� u
���s
�BÄ���ZIԊ�+;\�t�)��W�[B���AH�N�&������eW-�V��ضW�g�L
uX���)B�M�޻�zݫ�l�9�C`;-�1��DS1\1��P�FM�{%�l���KК��&�j�y&���S)�
ӻ� ��,��N�i�i՝=iNB_Oc�};�̘�It�ޕ�����gn�s�w�y�;鴷e
���0;��QN[�^]��=��U�� .*��|Si�/�}Ү�\È�֭Cgw/��
P�t�̴�x��C��uEmwj�2��zڻ�K���m.5��v�\�;wJU��b�`՗,��.��	�UzJ�	Ke��m���(� ���y*�!c5:U9����xk��6�l�̠�V"��%`W��IGuY��ʩ�o�E+���=f�<��q7xT�&�n���5�j*�ǲ��ہ���������&vIe�a�Ӯ��Z�����߳w��Ʊ���1Q�F1i)KV"���EF1k*�"�A�*�TEb*0����QDPF֩V"���TX"�����X���	m�Ȋ��k�`H�QV(���PPU�*��bEIZ���V*"*���%JEAe�QF"#��ĵIc-���(�DT��A��T�1���A��1TEU�Y(������
�"�ETUTT�UDF����F(��[A�X�-��"��AX�����1���B�b�J�0�Tm�`������b*������Q��
1aR�"�TX�UE�PZ�"1EcR�X���`��QZآ����(��W��TAb*0(֢�A���*U���(��EEm��TPR(1k*����*�V1b��V�FZTTb",PQX�Ɂ�Ŋ�b�Q�Z�*���"�ee�#F&,�[�1
�kR*�E��,E���b�-���  T`�m� r�z�*��k����9�*�}��GEk�Cm'�c0�&��hF�9�}���tV���1�
r���������F��y�X�g�f�=9NZ�
�U�vN7[>\�#2�f�����h�ɐ�G6���շ���Hކ�v���r�xÈH���q8��h�}�|��;;���w$�:w����3t�����/V�A^k=6�62KM	_�
	�|` �#,ث�+�t��7�ܐ��'��K��.���b��ɣ��uŷ���u �PTE��H�a��8��s}3u�>�h�r	s�R�0�E���#�~.��C�**`)b�d�� �s��ឮ.��*M��]i��O�L�d�<4,��h�W��	�t'�J�\0]�ӥF���YWx���'l�.�B����}��߆s��"��+	;|=1G�;����8�j�ވT�u1���'h)�E��&�;��K�ef�
�f�Ϭ������{�Y�M�;)��;�Un0X�����ga���_e�q�avzM��Q0{6pT#���y��Zz��6�o��"��ݺ��U@����>> �c��/���{���!��eRe�^A^�) �e�LfVK��=z��-�y��M9n�}ӧ�}[�rK�ѾS>�u��;;��$5�VǓ���[����ױ���e=�XnE�6)���ٻ���6q�=�$k;(@�+�Bvh�\�����Vp :`j\�nn)1�J^g}��W�T<u����5�Ugr4�A�d�n ��nRF��}Ѡ')@UӇ|�k�(�	�Gb,W^�Zu!ItY¦�T�U�Y@�l��Qu��_:`[�O�t[�=Û���Ζ����{םfe1���`�#Z��o�$X"'] o�ҋ�iAK�f�K��Kk�����u�G~���y_(�R=�>�����;=OT�R6$H�D�b��fՌ�����YW7�"q�KcP�^pn���2�I�}��ƴR�ϲ��Fԏo��n�ޔ��s�P2!\5ŭ�{���bx�5����[6۹,b�e��3,�����Ú�K����ַu:�1
y�����
T�SE �r��k�w���L�z�UZ~��cW��^����ʗ�:�����T���T�3xB5KS�X)�,��!h;,\LO:�{�5��Y��'<zkb/ʥ���eE��9�0��a\&J����P?sF�.u��Or��;4i˻%�ŒB{��2�]��u�]U�/S�����@zͱ�7�W\Ƣ�	�w���x����u,*Z�{C�^�d�r����;�M)crm܄KT�uT�(�B�}n��x�F��yLt}��	�B!�yd�؇j�x���������/��}�lg���U���S4>�=�����ѭ��x���W�k���E��?n*���%ݒ�Tf�����k>g�:���ώ����3�]�V�B�s2�'ʏU o�L8�i�:hu,�st(�p�dn
�vnЍ��V�����ئ�ޑ�:f{��D���ۥ�������gԵL=D��H�Q�w~jc�Vo��*���}y�	|���+��
u�����~��N5����V�f�q����Pc���7^2����(vΗ\�ڽ��"ϛ�lvƺ�G�^�$�3-���_]1=��S���^)I��ڔ����WK�¨n:�=z�*����m?^��NX�v+H{�zl��\i��yM�3�zfnWH@ׅ�(q���Ko�[���
���gi,����T�E�����ګ�6�r{QQf��#�L�h�͹޺�=g��K�8��:�1���}Щ�k�l'��WAST�0�l:��d���gdލ��|���rjI�.Z�4)#
+��I[�;��89��Ֆw&�i�XT➬̜��w �0e훃9�ٝ]�P=f R�Q;�z�T�k�І�JZ�*vf��E�}��D���!������&L��|�\����{0q��;�y�>�픪��
m�૕�Ďk������S�����R2�i��*cY2~���غ��k�H���8�ß��?�j��)yq.��U�\9�xQ��_�;�4فJ��N�{�k��kXO2E��ޙJ7$H[W]P��r�.�ٲϦ�Q��+Tdҥm����foxԩJ-�%��4MZ�M8�� HY��!_K�.�{Z�/hDR�ս����6_�HF���Ee*n0���� '�gI���V���O]���^��Y�ٽ��-�9x��h�C{���:.X�Y/�fRKOD�%b�^�T,��f�&��=���A<X�\^8��N˛�C;�U2�A
n^��]݇�eDC1dB.--����۹��ӣo�*�����8������	� w".
�\/&�
ܽ{��F�{�r�pW1p�YG7*��tk�Եp�=�?�u2�� ���:�P��L��y��ڼ�dl'��.ɒ��5�l<IΛs0VlK"�^ݣy*KU~#cm6��alMɧ$�t����=�gbÅ��Mynmɦ��O8-ə~��,�\|�UxקY��ʐ�z�{C1J�>�;/݂�J�Mݵ��f��T�-Ȃg$+2:-����)z�6��oW0�p5.e�vl�y2���k���v[��)�[O��V�P�-���e�\�����-+����*Gm#�!.(V��ھ����-kk�8�
l|��fC*#��L�B��=�`w�*���f��\�Kϼ��|uO��o2��SJF�I����he�S�ћ8�x�g���6�<F�f��=�`bF4[�T7�79]�3WJpM��/e>�O$v�O�w|(�����$x���͹מg
���0�{�:ĩ��*�5�R�1C..YmHҍ���F,+g�!�ĐL��ղxf���r�<��סZ�G:e�<�H[WT:Ī����,�P�kQ��Nm8v��7WO3\Ev�P9C����|צT=�Q&��>8������+�zI����FI�r��`�=��j���}<D�u�dk���@5m�($�VF��ʹ.����Yʨ.�ϕ�CH�q�l�t���q��z�����
]����
��Wg2���>ɡ��w�����Rю*U5��~(�ٿL#�`���W,�9dT:;z^�W&,������o��䐝!�K-�9��~��������V����A1��Iy�/�!�i����g͵��q#w�V�)�#-z��*�7��������;}�+<Wo6+�V�t�1b6�2�7L��(F�~rc8�Q��ku�����䶧��7��
��G;\�;*�p�ޝ�}r�n�լ)p�x�rîe-ژ��ss�:A{���p�Ua�4�0]KQՂ��9[,�l���{)1Ϛ��7+���ۭ�uU�3+`�:'h9�E������ɷR�ޝ�w6�g�Pl������ޝ�Y�P�g	+z�6
�gc��C컣~q��zP�!�����L�3}�*n�+n#f��՚5��m�:p�be*q�c��+��W��l�z�^ʤ�\=�ZdM���S��x@����s>����+C�"�r�0/�n��NR���un����y.��r=zr`��LN�^qg��7����o6[�{(�����!SϷ�gʑ�w7�3$y�����w��D��J�;ظ���V��H�t����-C�dh��s��F����(���r���7�����'��V��;=OTҕAblH��E�P��'��!�تVw5��,�8_>�6�[5��m��q�;�e�:�N���x,}o ��zn�9�E�=!��y�sKh�=��c#�P��ͅ�X�:E�bp���ʊu%�Q,���j���d���2{+2��:H�Z�]2랛���󄻳����=�輟��Z�ؽ�AU�X��͚�t2�3n,7����8N58���W���1D���9l�7��B��S����G1J%X��/e����MV_mmb����t^:J�m_!NtB�)�\Uԙ���Wi�+*�X�p+Ч�N��VPT%Sޚ(�u(k�wpDH�=��w��TX���$�i׏�\v�j%�Q�
z�reQ����N��V��N�'�nȹz7I�U���:�РC9��D3Wӻ!ϯL#[��,!@&T|�p��rS;v�kC\�3����� )S�gA��ӎۮ�����o���i�=E������y��óqR��E��Y���d�32;"�s������s���!���*�%g4���ة}�:fk\�h�`��y:'Mu,�s|zIh8g�5{§e�+�̤�)4(�ݤ�+�<�뭽U�n����!��m
�H��ܴC"�y�7~.o$��>���R�����Vo���&'r�$W��zcS�<���xmV������<��"���/lAh���V·S���Ń�]��������o�:d����h��9��%����ܛ��b�gM�iH��@߈�P��F;JWva����k�Sq��JT����Υ���)�u�D�v����u޻��$��y��-�׬{-@+��-]��%X�^�����ެ�F x��;N���1�V������74FRZ�i��+�1�4ec�r����sǇ���[�ȱ���0(fc]�����=p.�])�*ӻ��~kX�h�gzg�$W@@�[wF�H�Qgz�5Z\�5T(b}�檑��Oc"�nzݳ�/v�N�}EE��s��O�K�gf	����V5�D��$��<�X�[P�T�3X�w��t�t�5Jc�1�k��:�%3���:�]��-D�)"�B*�ol+ ��1	{ӜčJ���$ŒS�*Ujq�ٚ�(��d)���Z�s��\�*\���(��El����oJa8�����=cN�߽�h;�:����!��t�Q�"B�]P�8W!�=��ϯi���w�g���Tڽ�;U��m[5.yE�d�mђlZ�M8��E_
�^D���F6��o/wo|�{�Xuث����^
T�a�K�H�قdRub��1d#�kVj3� ��/D�.W�0�GM�V���j��R��<�ub����J�D�%.����2�ڽ�~�_����wQ��Q���*6Eb��<Y�����o�*y)wb$\$-�Q��'F*���}����V
J2N�Mފ��2�l��v�U�xɈ��4�]�]���@��2E��A%<�ptB���7�a�s3��t͑�ۣO�7�T��x���/�N�V��-k���
x�:n�[8�>
f �V�Y���E4o�l]���V4���o.�.υ��Vb�Wة�5d��o.�Ú�Em<}5XǕa��� (JȰ��9�T�r�Z�A��1����*rU�y�s�EH�N�5Ȗa[|�!��6֝�5o�#�-?
�2N��[=N��pGC�{���3&ptt�� _u��gf?6�0`��u�h?j�������Ƴ���+��-O��QaƑ²F5`z]���K�z������,��9N[pu�~=WR�:��Z�lu*zֵ�g�D�"�M(6�K$�ⷔ������8܇jt�
��ˌŚuW�pVe��Svt�-1*���%���f�[�oإ���DO-��tJ{#�O��\�eto-������2Q�n�4�Sh�����ru�tܡ�q�9|�<e�>�w�}��tS�vj�ܠ)��Q���	{Ӄ���&�4!Z�G:e��2Bغ���*�"��Y{yy"_1S(���Y��;H�9�(�܎Qz��j`Ⅿ**$ѱʙgq��^B�⯻�<�>�m^d=�vNĞ�V�.�%Rs˵�kOV�X�.�	� �-��[,�q�P|>Jq�4"��a�F���f�+=��hu�7��:�sǓ#���j�V�U�Ng��ۮ-}�9Zym������,O.�U�&dZJ�6���E-�ޣ٨����D-����������nx���bw��墬��8\�|���	��V��[z���O�d�B=�0Q|��~�<�h�#�,7���u ���κ��g'H��#=�o,�'��і�xc��r*v#^lؘG6�tyH�r�
r�jI�t��Ɇ���ռN�<���Sx>&U?.�M�c���pв�������'V��q��z��ǝ��,��8㞪!��dР��[u-GVz��42���f�6�ˈ(���ӂ��I�/U����;A�����`c�	G��������^-��u&O/!嗯�>������d�π�3�9���gc��_e�����6��`��8v�޺�'�-�~�;]����u��wY��eg��5ݏ� ��w�f�=h�o%ӧ�@x)Bz��sy���܂�8�	�1��k�%���@nRF���7��Qv(^sܞhH���Ίbc����X�Q�Y^0Xɺ�r���(�l��Qu��s����h����>s�ҳ�8f�V/Z![�(m-,�u��f-����e�Ǩ|�o"Щ8j�_3�jX��u����T�hړD����2�f�k:�;�)�;#I����2���n�m�{�C�Сu1�zf;�E����R�'l�0#�R���t�Y��9+������B�c;B}�S���S����ͧY�n�e.9�p�����"^�#;�!�7J� �l��5w{`��A�\��2Cݠ<�T�'Z�\��r�����%w�-ט��Uh9E}��T��r��޽\E<f	���M�l�U��e�~��v^����@�]���u.��oEgJ�*�dt�+�fH.�*
[�v��@�s���.�)���O^e���5^�]`p��ݪ�e�pu�6;���C����/��ns�S@��;�`��Aas��sy�u��,Yʕ8�+uVhM�y��0'B�5�E�� oM�6��ҷ�q*��<����-�N&�͖+]$JK���r�0����Um��v\2���n�Ў$1ky��wc�H��#kqb��M��V��7.o�.�u7�c�ϟ5X�"���y��C ���}�D��Nm�E�ͮs��D��N;��j�cĜ�8B	���o։�{
��7Q�3�5�Xk���򆤔�p��3I�x�*3��*���@Pˇ���_N�m��ڕ'!��<�����f�P��Q���%Cz�l���I>�]={S&��U5�j(� �z2��K�,���s�3W���\W��a��ڇ�5uKh��Ӓk)Q�I`Z�+\u�_�gaר�um<������7��mM��*P�]��97�Җ��&�/QN훑�4t8̼�6
��F��b��iT�%p�W3"̎C5�]X��8��̭��1�c���eW(Jݩ��� 
e>�=]�_!�*V�!Vn�
c���/���1YgB|�J�]������3��< ��D�e���0=ں���k��}��_!�����c�_��ú4�LH�A"oX	4��=JHE��[u6�f��g��n"]8�"��lt=���������^4�{%�a�dq
k-���t��C>��&�iW[���˫�ҝ�Q�-Z�+7���m���xkw��mU�%����m��(�6��z�����bU�n��/.x3�u-}��$E�$+�Q���]����z�׀�{��	Ϟ��r!���*�&���	])vvw�$�5֡</v�}��癙'������U�s����m�yt7PN�j�]���Y�n�P���.���G;zX%2��eBZ��ֻ�YD�l�]��[bwj��7M�Mu�J�+vf8�"m9A@�x^.����ף$�+5�������	�*����םz��v�}�~�����*�*:�����E����U-�0�X*[UQ��"������b�E����cH�j��"1b,E�����UEE����E��UL2�m�APTQm(��Z���Um(�1�"
��X�U� �TQTb�����2��+�1D�$DX����Z�@��U��Q�Z�Ԫ�Kj�6�B��	D���"�*"*+Q���UF�#iA�1����(�DD*�" �X��*" ��Z��F,AUV8R�TTB�
���E��EQR"���TTEX0R��b�F
Ƞ�F ����1TDQ����֋QV*
��[h���F�	l*�*�*���0Q��"�eDb�`��`�
*0PTUD��Ukb*(�,X�����EĩA�EU`�""()iD�1h[QJ��J�gq�����Uf��_q}\D�wع����]�Z���;�Դ�ݖw�_ǰs����%ͭ\��ގ�*t���wsy��d���U,�0N�['�T\�cdX"u�3�6�nf�z�%��㕹�d��k1Y�)t0�iS��yL�`w�4�OX��i=S^R���m���t)"�O.����j'&5L�^o��R�lf�>Ͱݳ�1�S7�6�N�k�zbJ;י"��D�q�˾�Om���1��W2�����b8��bp�����M���Y���jj�뽚��݇�[|���}�K�#UEߦG\��ΐ��Y��T�MGv������d�#���R��}��U����v����J��8��O�- ��L��lebv+OqWU��8�ꉕ�u+�n#Wu�C���M$k�/Υ�������p��1�~kt3����sTu��~�>�����+���_	H�\`��:Sk��J��_��s�Ⱥ<����M9L<���n�b���a��Գ^�qVX,��.�J�0s��^�]3��eW���v�����P���Mc��3Z��@�R��Í��F�!�d�V�)�>�6��l�Z; ���l�����\u�M�YU��f�;�C��mf���d�8�Q9���#�^P�&��א=����ajp�װp�r�q�\��:]�0����\utWV���N���5�O�ۥ�*Ʈu�p�,��G+e*�Y��+g�v
x��Vḻw���s�`ڻ�����k�����>�A�IL8ȋ��W�˺:�BV�n�k���ñ���ɳ��Y�|<��3�_K�J�"v�8J��pK倿��e� S��o�<�qP��r����M��c�3�a�αMc6X��,�yb�G�h躞�U�'~��VϔC^ְ�{�yy��o׆!o�=��F��`�a��X��ޛ1qI����5n�_�èf���?{Z���m"Qǲ�0�p����S#r�i݌�^�t��ﱍ�+�X�ICB�wJF�l�̶ќ��]�$n�EϹ��F����c�Y�L�9V^�ԝ�>��˅��Iu�a>ɟ:Tq�=h�9�fK��[,�B�F/#�Q[qR�1�g6�3�l+���L��Et��e��Yi�VVK�g��tJ�r�A�1HYQ]�{a_�
ޑc��=�lƃ�r��t��[��B�����HS锣�Φ���*�
#q�#,�Uz�R<�65⠥X��7[k[���F'{�,�u�9ݯ2�8d z!(͑!m]uG���>\6����2^��^"��"���W`Y�U��{US��`^��|H�s&�z�0݉���{�	�'�~0��(kĸ^��@Y'��F��y�Y,��J���ʂ�gk�ӭ����&v�)�����*s�G.��SCGs[���S7��m�˱]dwvf��31������L�j�i
u�3 �IF�&�s ^5ò|iWYsB�y�1�Ez���(��y-r��z��+���{�j������g�)r^���KTR��U�/f�1����a{�:��'���U�R���ls��AR����\&e$��D�t�ҌQY�Ύ݉��AQUs�J%�l�c]E㊯�/-�O�ms~�s`4��v�g.�\(����ռN�C6�L�b��������z��s!��f&�Q������D�;b�gc��u�5ė�`�yvU��\�	V|��/*����W	f3c���^�b�5"cP����Z���~M��~q��E��$��(�kN�aA��f
��;륥���{�NDc�黧;c~��B�07#:(�6gqS��-�g���M>Z��y�{��S�$Fn�}������b����2e�ԭ��|7���G�|����r�,��`v}2�N�6�J�1�u0z~S��'*Y�SN�N�I��+�H����`:S���:Ѱ�1����sHk�ˎ,��=���u���p.�'#��0�x�<Z,ԃ��J�I����
��Ub�4+kz�e&2����lQ`6'�i�Hݡ/�F%��a��";Kh��4]	��bEV�X���ǥ����]|:���X�Nv�O/W���8� ���#M��z���r��+��&�Kq�Y#���Db������`�>hxNS�z��l׊]tk��.�x}4K
��ٛ��R�+إ�,�b�ɗ�]g.����$�Եh�	{Ӝ�e3^�'��R�[<���)��O-'��)���ڵR��Nt�kG����S,�l��'#�k�5����)�\B���Q��V֒������#/yf�}.�E�!t<�\�{��z�W6�/V�
�X=6�9%&��^Vt��''�j�#�G�2VC��̎�VM�{6raAo[7Ny���r:���AH�qb�Ⱦ���� ��T��U:GrD��.A*EN�a�Qy�ba�.��#U�5hel���� �"kxf_eg19A��v�I3���T�v�w��$͌B�\]z��� aP��׶�=ܚ-t�4^�5�mHGaL��VM
��ilU(ׯ����o���R!D�����J[�p+6�.�w�u��ՅLQ�
FA�Ή�sf�7
M�c��κ�V��g{zǕ^M�p�o�~�v��ʍZ:��"l�4B)�E�.���Vt�bv�}��7*#�FWs��K�n#�v_�6<���%�\W-Y�Eשn�d�0c�(7���g��;[��]L_q�F�,Ӎ�rń+�LQ�|o(N�j�ΫJ��ޤ#����byy9i����v��O�"q�>�v���ؾ��܌J�V=(j��9���%MGB�.�oK7�U캍9z�.;�,��)���3��w����;�E�˶�z��[Ͻ�S���ecX�|��h��x�u1���X>�c��[��7� �&գ}mk�>-$��f�U�������e,���7��Mpu3e�7����v]uz.�է��sY���z��zLg�.Eފ���1_!orv*��
\��J.TV�Kk�j�Pi���:�?t��6���m�{�Y�A�e`���pi��\(�5 ������Y%�or]�Q��e"�y>�T9Y�O�o��:��3nmܝ�tͨ��gw�Γ!��y��8p~��B��%���E�!(�-�3j�5��X�'Xo-��&�Wk�"wJ�-W;�˒��e(�3,�UED�!O<� �T�m�t��9��r��Kjdc�U�g�B��s1o�$��R��;�j`��0�uؼ�3�� Τ~"��/]R�:]U�ȳ%��^��ݸ�,����+�7�!sU�;�����;��%�2�zF���p��==���R�\��Ά3�l���uj̽��P"/����\Qw���P��e��.�[�NQ<�;K�V��;.\Q�Wc\�fs��K�t|����Ff��1N���B���M$k��Q�$K;^*!������C�^����=�׶��k���L��p���(���.����:mv�iWYϯ�x]�/�m���|T����<���͝�R�o8�,YޗvK%Q�9��Ȱ*��ڜ Ό�#of�)޳4�]�f�w�:�K�����������0�BrN�e��YQΙw��D�=��%���r�x�ی����l+�N졃Һ��^t ,7J-K:Q�&���o�s���ޞ^�3o�~@!��.�<���U�;^3��p_� v�� >����1�7���NzU�T�:>V��S�{�%�x]ybĤxFj��|�o�|�ߛ�f{}(<#vc>Oj6d�o���������,_gE
���@�W�'��T�����Ώ21b�B��Ý=NUF�C."��L��8s!��(5�,U���m��ޙ��j��f��,�C+��W�B��ϧ�};w���Oc<�{p[�}��/��w'�VObu�{�{��쑭 =�c9i���"��(���)��t�l5���[����7����%5Ü 7ܚA�s]���N�����2����]}L^�y�a��E�"�B�'�[%"�����9���Lۣ�=��y}���̀_Sי]�x�[z��������o�lOW C��g|k��f�oc=�K;юӻ�4pJpV,�P��k����Ss˃�+=.i���UCQb��/!oh.oH�y ���[�<+����s�@�`:��R�����O�m�g����ߏ
�k��7q�g\��W�;j�fk��:e.W����$�_��A24:e(�$-�u��g���Onx���t_?Wo_٩�6)j�j\�^�(ȷf��Z�M��Bړ�ڞ�Ù�g9r�41���,C�s�%�4l�jV�Ȭ�E�L�0�k�r�%<������=�E��g����V#�`��W\Zq:ޘp/��3@r���N�ذ��2.�׌�<"%]��8B�?���l��7�E)Ip�TX��/U|qymi�͔:O	^�"����f����i=�'f�|j��AS3�{m%	a<^��S|)B�����"��5��LB^�W������K�ek�L��0�b�> �+"ã(�窙�^���J�E��4���\�d�m�:n�
��ׂ�_l����	6�퉣�NtK�
�Թ�	��m�t��f���m�����y��#Y��Z��/5h-ٔ��~�UX}xȸf��wtZ��;��u!ې�;E��k��gWe�ܡ�D��O���{���؝���^����aF�:$K��l5�l<IΛf
��&�{��)�k��w	��0��>ī+�/$b��fw8��,�w��:i��KsnM_�1��﷋��b�l+ޡ����HGf$x�eV�ᑤ1C$Z��T3!����k:��q}e��=]���$
�n]�v:"Ztz8ۜ��,҉pp)��40K�2����x*�}�9g@�(��
8�ًV�L)��yzmŞ#M��z�E�Q<*p�n	ъ[��l�$r�
�L)W�4g�y��9��f��CMS�:�wl+�DX��6{j���EV��8��,�[qQR������g��#N�k�j��9�<��W��+Sh�L�wҨ����rn�K�ʋ��7�:���Oe��jp�]Y-�DM7�h�HXV�W[=DeZ���{7��cM@�N����MZ�Cy�n�W-�p��:���@3/���ۊ�l�I�䲯aA~�(���g�q���s�!͜aAo[69�G �#��s����F�/jg+�(��6��[�T2�>��,�,nʝפEO
U5L��e�{Ij���'_�lK:�zTKv�A��I��h�[�<+�V�{��/����c��Hvu_]���}��z+E�[�rc�V,��M
����Z����uZF�	���Y�3���zY�yD���O.�|�
���H�	�׮hMa6+��,G��u�<i̹Nv��N�_V�r�=��I�7��3���c����8O(C����p<e9�c�Ei��ګ�V��Yo�3E�%��)�)��
ɡ^���SF�TΚ��g�F"�V謘�X#wsKjc�x���\0i#/`�:'h9�E������ɷR�ޘ�Gq��:��SK�c7y|p�T�9�DHĈ��l ��v/Ý���컣n0�/
C��k"6�C[SmT�\b^K�G�T{'v�D�"vո�Ju�D����Jh��J�j�]3{tX��9U^�+Ӗ�sg�!��A�)#{�_G��k
y��z73!�*���'f(�Z'Hf��H�z���o6[���YV0j�̼X���S���t;`Xz��N�sǻ�l��X%v!�NV��iУ�]A[��^����oc�]EB�<×P���l6��v��{����OX�4����PD�R�{e�q��lUJ=�U<�3�c��L]�W�৐�qKEX�]���T��rwʺN�E�kF��#9�J��k�Rw�MA0}�ߢٳN��]���]��q�}ä�9��H��5�;'3�v��;�;�Iŀ�ā]31�m�]<����]���h�S���0���H�A>�o�K���X�f�n���)�_�$^c�>�,���N�r�a �8�S$*�\c��\nBQV��E�P��'���E����̕UO;T,y��+Q~龹<�_B2�ߩUbdu��
y��7��O�ћ�̷�^]��-�z��xnԽb|�U@8ܸ��t�ڥᎢ�}�P3�a��.���6���*����j�M���O+�l�x�E$g�4:���C9��D3B�wc�N�J�M���׮�e{9��6��k�jP9T�����q�
Oy�#�m㠶3<�Mt���XXV��\�M�iLlV�Ӧ����8�,Q�%ݒ́
�A���.Th4�B�����������ת����d�K\u;�I:�O��z��C���4]Բ��X�i�J{��b��>�N�'<<��g���l,��#�5�L��DN�Ja�+���Ł�>����+�����/)��l�P�Y�y���T��v�8K��U��^s �Uq����	�/cCU蠸rj�W�۲nZO]�]f��jq
6�Ժ��h��V�eovV�= <���LD3�FNowih�۶��,��̥-)�uy[�y�Yō�\��>Fuj�K�����d9k�j|�s�GC���K�b�޶s����V5�SE�9쩽�E!�ಜ�$=;(q�]��1)��l޻gs<D��x%	N�9,S�Q
�	��B#�� !�n�1�S�YҝM/���u1�H#4����_�)���촌{��[��L=�l.t՚��l�X��#9j��ǥa-�ˠ�\v���-�����X��9S����-p��t���x@�����\�,Q�Jޭ�������l�}��i�ٹ�nQɣQw�8�/�p!uti������1�MQ��u���b�=6W:�k;:n��oKr��k7���t��]���q�Se�ɛ�;���]��I����Z���ҕ1\���G�tW#��복�T0�uxstdl�J�]j�=�f�ս[���1Wi�f���j�i�r�$+�fR�}��+X6��&�Ǯq��QH�|8JS�"b�x
�k�:]�GwԂ����1m�6�f�Ӄcxӝt�'��x�Xq��w=]l�e�x�mn ���WJ6�Y�)�;Zi���鏵r��K���p�VO�:�Q���&�������k���,l��e��[o$\��.M��O�;Wc�E=�o&� �듚��
C�zf�+�W�?�p�ݫ�:��uAv^�m �BJ0�o(,뾾��a���[Ci���۠ ����\�#�B�~9�( �:��1�����flB�ʁݧ�.�<�S��'2a7��HΕt��Y�N������{�N-���uKR5��4�g>��O��"��.�ܻ����&\�;�����%q���瘁0���AK0�\��]d�jvn����h�8��Dڳi�v�%O�0��9[�)[��B-
�����V�D�������z�X����4q�-�VEf��+kF�J��N���F�r��jx"���x_v��0s~�M����]xZ���f6E+:m[��[E�[f�ǆkQ��ي\��]�ql1�o ��컥XFge+�3I��b
���nv[�*�TȷnR�}�R��4����c\ޝ�c!�]	��&m��]hZr3C}Wv�z�������pmu�]k;t/4]�PBL�۹6�j@ҵ*q�WGM]n�\{��}�v��,G)Z�S\Ó��K�9y�8ż�ï)J~F�+%a#�T���h�6<��"��`͵�ٷ37%b�A���	�}�`��Q鰫Dz	`�u��79�I;���k�9�rV+a՘��-Ue�U�r����֑��O��".����Y�Ύ��&����0��:ۢ�G�m�T�|�1�q�����Wq�/�c��Qv��"��]��3�ů��w��վ��X��A�
���UR0b��A��PEEb*
���DX�e���2**�Q�*�J(��`�X������"*(�Y���b�""�R"1D��`��R�� �Ec�AAS(��TQ��Db(���TX��
�ETX0QV��D���Q���DX�E���Q+Q���2(��Db)F,CW���(��ATQPU!DDjUDEb5R��F"�Q�0AUE����KlDYm�
�F,EU�m`"��(*�[�b��#ūR�T��-�QbQD"���U��Qp5Aqj1X��UDA"H��1A`����X��V(�b"�1DTb��Tb,QDT��(*
�b+f��*�AA���*�E
���Q
�#Z�C�QcA"yR�:��V�so�E��F��tg�dΕľE>t�k�α~�� �ۧZf�gx�#y���V��	��p��Q�-���������OBz(i���,WP�|A�G�f������:xnW$T&DZ�O�v�=TN���Cv1���Z�G���V������}�ta��ܾ��r<�i�]x�͎��W�]F�e�Px����dh�q��E�{'�芉�~�Z�
ȫiq�r�{}3=�����Z!t8��(�UH��t�0��N��p
��6�h=E<#Ӧ?NR<Bz��q�9�F,<�f�Y&�8�c8��/���[�#�/WW�N�<��[�9��]a�*&TŜl:����쫢U�P,�#����k��:�X�������0o:CLKޞB%�VY�B��=	��Wm��eD���do2��iս�]-;H�~ޤY�O�,]7�I޽y�Ey�!]2�nH������԰�J�;5��nO)=���/�{��*�m#b��f�r�����[�Dծ�$�pZ.2�����V��0���[Q�Ȗp��gD���X)Sq��¼�j+�y{��bڿsi!b�bY�������_��2+�<�]���}ˠ{�gz(�GB����5���{��q��PwW=%�k|r��}�z8��O:ab�U���iT���`P�`��o�j�l>���i�6�}�pYo~��Ys8!�L,Ս�N���u��UH���7�٠�:6p��eK��f��PC)�{���;���x�jޡu�DI��F���R�p�E��/T��X��V��:O���B�c�.=ߋ��J�~�l\�݇�+*"�K���F9M��.�.σ�X��sLg�(�hU�sX�q��V�4;L�Mr�r�ʰ��eF@x
�,:2�nUz������t|Ojf���
}=��\;�9�ݓj0���Ή緶(߃Zv�¤�M���Y��g�3�9�K��oN�".|'fx��6�C"������f?'�Ō�jЇdƃ崵Dv�vl>�������#=��g��T���!�J3]P���EDW�*g����@�+�u��w3��X�yW�^�4��+y�_�x*|�����Ύ�*��̜�/#�TOʗ��:L>�<_-�9M��Qv~�7.��u��]�{�*�Ur+��'7��"r��t'u�3]��,��f�&K[#5*|�Qg3�W�������G7�uؔ����+�+Mva��P��Wʥjb�Ԋ��[l�=*�&)k��������hq�ޕ�n�|��_��S���]Gғ�Q�ԌC�Jd*�Y:(�V'T]4����v��ۅ.Ūtz��C���:��y^WS��_`\7z8����k�i:�����+o�B^���,�ɫ��U���K�o��i?^���wL�G�AY7�/�tl�E���2�x_m3~NG(��+���i�M�p��G�k��Uꗰ\[|o���7����HK/�bK��g��7�,���M��qY�b�fXQ� 쇗/a+y��k`[1�I(�C���`��$�z�tL"�-�f�Ng�m��՞���8�}��z���X��
��r�l�gj���b0�������t�rS�t�ߏ�-{)����P�P�
X��&�HXΆ�R���/�XOPгM��XM�̈́,l-�kj�h̹�E��Q}�iA��#��HD�&F�f��L5]�t�C��`�=��P��s�ڢ�����3����z�I{��;Nl�f�)7��\X�Wtͭ��4l�{X{�紹|�z�K�K=e�^π�P?)�����vN���TV�_]4��7-�5dQ��q�����^��N�����>~������x0��]��*���Cmђ�n��v︻��������Q'��+h�S�/����5�y�m,�@w�sƅ��{����!7�˨�a�V/pq�3�:�z�c�j���1��5��e��d�Ƈs;��3r�A�8�h��m��c�j���w�
��e�E�z�0`���go�`CxU'��@��Z��� �8\X��ֿ{/��q��C=7:���0��}Ѿ�Qe_N�}��l-�x1cS|-�pu	�^/x��"X��L��vv��q�9k�=�oU>��[�=��iܫ�w�\ܝ�~`���{���SЌ���������QciJ]C6K���T�;C�g���é�����H���\��iZ-��gmu׾�(W��rV1sMf�0۝p�)��٭�g\c��c(�mP�k-�λU�Y&�tͨ�LIGf ��2�� G8Y��P����(g�^�<t�1�o_���bW,�&���_Sn䱊%��=3,d|��l4���Z�\9}N�WM��L����ܝnf�0������#�j��`�* ��]JAU�a��v&��J�8����>��kֶ͸+�ճS�YN�d��!V:"�5�a�ެ���8[��W1\i�X~JOr҇��ϯ�3[��,�+T٫�H��J�'��`�=�tM�ӍL#�;i�gX��}�,��i� �vE����^3�d��.�<�WsCy݋S�M]��K�=�wVW}fE۠{a���r�n H�ǘ��c��{e�����!c���u%�~�Z+;WQ�rm�$�A�����;�/㫾J#C���ʌ��aps��g����F�7�U�2g�]�,�F`���D�W�P�_86),N�HY�x�����c���ώ��*ē�/��o�w�u+��n�'M�4zrq��9���r���*"�$�5��F�#�.�¼��"��zfu���0O+�#�ˁ'���po��.Z���.쇉b�z�����\�U�'oÄ���X�N
!�蝋�W�of��Q0��$��S��.�����{!�ġ�/�6 �G�h�4��,���g�=��6A���J�TN�kw�ݡ�����X�P���)�y����)��J���X�m�L�7�����(:�,���
̆\Ey�F�ӻ{\m�Qb�֤(�!QٻFN�V���h����gd��5�P��ܢyU#~�t�08E��tϰ�Nve6��f7����Y�_��<�J�)�R1a�"�Y&�q�"
�o�����N$guh?S��|Ҙห��t���SSaՕ�\�=���x�H�k��f�\���Cb zˀf�"�S�V�y}�R�O+W^J����}ʇz��l���:7���bBoFm��ѣ�G�Xs�Q����A,�@��W2�����7�F��6s�y>z�g"^wb�8�D#{:>y��d�T"�ӉU��*�%�Du�R���δ�\�wb|:�~�ʼB^��1 ��4)
ac�R���?F#�)yq2Ť�_.Ǔ=�|"-�,�����`�X<�o\��c^g�8d k�R��"Gm�y��V�8`7;}7x�㬍8:{�ʝ��cfm���%td����[e����5y�9:�S<H�����([2:��-�olD���Е��+<)S6m������ƷQ�osTN%�j�b,US#��H�h*��١��ޜ����]3��b�L��L�c~}���7��>U�N���/�H�_����lՍg�е.xt3�X(cJcpH�B|y�z�v��X`k�"��JعWvx���W�.8�X�DY��p�f�:����V�>�W�MLK���"�	�0��RNPo*��VTd�	Y�Q͙g3-M �&Vbb:ks���X[9q`��20o9�&�a{|�>{t$�Xr���s�sD+�l�\���-k�n ��&���8桶���6!���q&���ߗ�ڴ!j�'@�J���w{0ё�)Q69n+[�T�񳋜t�̬���4��"��[�b�Dv��!�^�.�3^u��	�[/���0�BB�m��\cS"2y�9r��K�G��t�l��^G�D7�aLY�� �3�U��m՝�p�k[)#L����[�/Fn-�x[�%8lV�4�߼�\�\8�]k�0���8���}I>�;o�ϦT7����n&'@�Fk��Y�+�H��ym4�I:y�e�^�����>�l�O2�����vQ�w��U%(*x����%����n���a%�;H�#6�8��Fy�O���꫿g+Qzp8�Tu�*�fl��Q�˭��<��{ږ�D0��qyH�R4�]*��!/6s��<�	���B�6/T�:๑CgbU��:v���(�Q52:�C�ee�)j��6��Qc=KFOk"��z߄*��s�
i�eN{��FEP��H3��C����_C�ᰌ�m#t�q`7\VEV�7������l��j��w�4v��"Q#ð�G�'��Ѭ�L�x�vl�����O<��8�t���}4]9
���

���5jI��t���й��N�4
.�[�����}�P��V�)un�dְU�j�*Q�T(m��\D
�E�)%�e��yi"��Y�Y���/;��R�	`���d�Y�\zvlO*��<���Ǚ/<�t�+"��qss\��f
=�d-Eq[�u�,��u���g�!�'i;��@�&�&_L8��jU��3�!Eη���'�4H�����I��YP�6":�����ì@f�D�ox�(6�v���5
��^|�v�]KQ�LX7��n�ۦ=�	~DT�\<4k=F�䌽�����6h�T�����'ӛ��2���DGZ�5�sVS<5ԙ*�;�}�BDO���l��Es�pխ̍>Z�����7����\�=^6*�W��`�V*�ִ��ܦ��ϗVP�F�� �_�$(ռ�������vd�ǺѲ򼪯� �\��G-�����E�z�1d��Jf�|��v�g��t������47)@U�4�[1F�?���|-��P�u�M���V̌YܗJ��*4�S&��A�O=��k%Ƚ�Y������[�pvs������gTիO���ldqQ^���T#}.��L�g3��/���znm8�E�5�f�`o/}�U�u��*��x���-׆�.���5���t��&v�V�'����X�5Lc��S�w?	��C�F���h.���C�i��ڃ��ꪰ>����
� ��K7�uG�V}��e�⺥�����0x�Z�����n<3n���<5G)26؎�Rq�T��Š�[���y{�$�6�u
2�Q5JY#����L��H�h�y� ����7�q�mѦ�����=GgB6��e��B��g7���4����V�[2��duJҸv�Ip����kE]N[�XB(��ڭ��i7��WJ�\����t����Ճ�W�cfbE`����?��z%�P{w��4�������Q�8��輁ƽ]��V
u�'y[�AK�X۝�/���SN�����Urc����F���q����Y�
�6j�J�Ć�8��{��77�|��WC�Qnû�7���q��n���S�l��^lD3glR�������f�㭈�pQ�����r~/�˗KՂE�J�Y����x��=H$]���5�ݔ�of���m�5Q*���%׏�R�o��=�/j�*}���wo�7�2�nf�1̬41�wT�n���^Rz�ī�SSWu�m�^�$�I6j����L^*��fT����Բ���P���Eo�,�������c�M;���#�OW,u�1ujz�'�y��D�y�3k�I��>��}Dv�-O�n������d���W��<�Ύ����X5L��(��Qq��#i�8.�0U矲GxW�.�'�߳�$���)��g��:^�Xn�|�7�G�NJ�F��de��x@�y��a z��l�qOw�6L���*Ս.�[}��)nG\��w����5������7{���̝��w���C�ʧ��7�hp���}�g؛�m>�36U�MxZ>c��`�^�i[����yS���j��/�=9�"Y���)��nkiζY�{���(�a�;P���46}��f����;�&�;�,ls�6Ӳ���Q[��A�޼�n�JP�t%�"��e8�"��vO9=�/����)��=��Xlr����^�@m�(����FKoj*U��Oo����͕��>��R��7�m�NH�.�	V�k�r�yVS
��+��Z��Ts�n7C9��Y�׺��mn �j�zr\��uQ�t�L�˅���Zr}���VO��ގ�%��H~h�[�}% b�V{�B�-�2��52�&�+&�ɵ��`�O���ߊ2���1�O��~x5=t���n�魗�}P��:�́[	u�'NTwٖE�:�Ru�'�]�&�܇3dh��:��Aj��`�f5v��μ(j�����]��"��53{2�m}�NMV>{9���Un��9�c%rJGDdޕ�@����n*�/��m��L�&ӥ�A)&�S(���X�-L��6�9�ײ��6�Tx�q)I[��ԉ�z:$����{tӫ��Ѝv�d�D$G��]eQ�!�v�(�u���e\Ÿ*T��d
�9�D�?j��`D�'dN�'�uk^�kt���n�զ �i��JqJ��>|P����R�6Nq8�v�/v�;$yE�7lL3l�r�dԦ�4������ͥd.2��O��}��}�����38-�-�`E@\740 �V'G,LƑ�!�A��w6 #WA���"#�����B�n>�|z�m�ͥp��A	���.�C��+a��f>�gd=g�˩Kx���1BĖ����F��l���,��uA�6��F�V����䢹U�b;�#]�J�Q�u=\b29҉|�}��Q6��c��umfv�t8[���ç*�,G"���do�4��|GM�߆r���$���e�K���tb�γ`[RV:�g_a��Z{D�J�f��xR���tx]g7�ɖpf ��ēQ�u9_@��iu2��*w]KXq]�ՂRx�]N�;�s9���o��i�8�Y��WfRR�Y��`��t%�F-��o��M�gY\�w��m����C�/n�CtW^e�]�L>���e9o��O�M�i�F��d�Uւ/4���/���Vƺ���m�-���7z��Ϋ����goV�H�YnRI%Y��g;5���<�4bW��w����gg�u�h��]�O*����}�4
�ӧ�r%��;�(�������7�͵�v-Ne5\�i�X�fp��� �n�|�����e_T����!��0h!��a
��r�owp�7Iw�y��jr!R��j#���u2K�Ő��� �J9ŀ����K[�=I7eƲ�Q��Z�5"���P�8�����u�p��e�T�y�5b���)خ�Mͩ�ˢ��A;a7N۷d� b�{�l��ʴsj[O��p��iw.�X��icϋ����Jo^]�.+[�Ģ���:1���I��R���`�3�͂e�EY�WΕ-���ձ�psgFd�z8d�]���!p��+ir��Y������_4�^���97:t�w!�;Oae.˼ъ} �w+��O���ьf�`}5��0uf�n��G���c�41˸�OgΠʾ#�t ˷���ޘ�3d���X�mj�	j�����&�l�)S)���Re{�� +��	5���3`���=��1&S�G �t�:އ�����۝�!�N�������R������9kG���y�oߴ�~ɖ,YQETL�X��U��b#D� ���[JAQAUQUb���"1��t��,ETDAU��"�"("��E���ڢ$�PPQEQ��TEUQ�"��ŌUTW�Tb#cES������UUQAE�֪*�
��`ԕQ�QX��TPb�ZQX֢��Z�-
���+"����0�� ���PEDb"�"��#l��E�(�Pb�(�**�P��*�A,��U��DTb�
�(" ��c�
��*��*��b"b�F*��R�E`����	QQTDEL4�1F0Dc+#A1DX��QTAA��`��Y�
(�PDDU�����TV,AV**��Աb��X�"�ŬUMҤK}��k�v���\
y�k7�j9"����ptgR�x��e<grW�_saK��ܩs���g^w̗�]A�˴d��h�m�V�;��u>Z]�	-*eaVK�Ձ���rʣ��R���ô�ɠ����z����l���/(r!��c��0�t�������&��{�4��/J[�_�0s��X��G�X�Vm�r!��b#)�����j�{��q3���ue۟k���Ǧ�{�fН��j��5���^z���eWJ+k���C�����noq"���������p�G��m�q�ע�9W?(�X�T^�S�C�:����x|y�Oak�}�r�׾�%�ș�o�GU(�hE	Ƅm\5�ZY��W�>Y(����%>	���{��R��c��B��ug����B�W������3Y�j����j��֫�t9� W����.��%���U��7e�~��}o���
x���cX����=
!��h��ڙY��cfy�%b�]Ae>9�;�g�( &�с��A���D��"T�ø�@�B��rM���#ˤx�ǄV!��j���r���L%[�G��bneD �-Sgf�h_��枃�:E;7�E��u�l��Eak��fozn��;��E�E������4��*nO?`;C`�U�d�%�^'�{v����/��i᭸+�
�tW^؄�u�[}{:}7k{j;+uN��ssϮ���vD�e��!\���%n�0��G7;R��Z2�8�T9�]���m%dȮG�F�X��U�Q8�ns��i��N<U�����a%�J
I����is�3 و���v�.���76��q��ԂE���O��a�-�]����fG-��iMaЅ�R�7��U�Wn�8�@߳��øh��;�Ե����hC�u4�8�!�껕sX���U��@����nV嫍�
��Fk��x��o����{���\��8�Ե��+_5X�������N�땚� ��7�M_W����C8�عY������y# �`�h�1&{W�|`����V��9�^����7٣�}}��]�[��]q�Z-]�hN.�j�'�ү׺Pҫ}ù���T����Mn�����0�¸ȷgV��[�����u_7v8���1�(ɱA_ac�õIdH��{�˻ *�٪@�7Z�x�_
[�~�ן_E,�2��kˬ<w�r����[M��� �̋�;�����O2��y�q1�z�;��w)[���i��
;(+'S4/�5n�u�yx���<a�Q�'V�v=�*�k4��5��]m*��m�t�\f���bR)�#�<���ܮo����1{�0�lj�$�mY�c˻��K�E��@c鞯>=S���j@v=�������G��{~�{���u��1���(P�� u���)ր�e۱�4�4y��);�~��c}��J����]���4��p�N��Y�u�Y3.���>�Z��Or�N��\�r-W7�J�Шm��V�wv�L�C�;M]iF#�����N������2�o:b�oB��p%F5x���'?D�[Ǫa�M�Ys�����s��ԃB�M�b��fV�4de�uG]��dÆ<]uN�C2�I��m��b
n�u����� 0�W\�78�a�$���T�^�/c���te̔��swr��3�uA�Tg�΁���)�"���h�YZ���wݫ���hӨ�Sq���1��o�\��d��v
�X�Վ_m�ʛY��u�b)�[��ڦhb��s�ո&�v�g���j�=�Z��y*��5�]�W�c��0�'��/7��N�R>��c�|�H{{-Y��OU�g���[�.�?�����~����մO�_���3Af=�ݧٳKsbj�;H;T3k
�V�H�����VR/���S���y�ԇ?k/U.������>Qr�ډX7�(�ع"5�C�3Y�yN&�Ni�՘Rjs'( ۽�G�^?u�ꚼ�8�l��=B��w��o+:+8�������يW��)0��g+��c	�|_�{Ա�ym���"���i��Z�M9��M��N��T��uy3�9�z
�(qKy��gtMlNcI�����N;��\��K�ް��׬gl�B�U
������Jƫ�4���g���o:)�@���h|��æ5��Y;2�Tj�X�ڍع�5�Y��s����2L��G31>�O�`���^�����\���������*����Yr���[��Ds��k�5�gk����2c���k���ڣڮ���j��{�m�&�ysw9\s���&�x��(ko�,��ٯ�m��׽�ώvj�UfJ8�AW<{�cr_��t�&�<jev_�d��SZr}���V-ɪ��!�T��w7ٷ{�f�%H9Oj	n����5��7)aS7ֻ��`�6t������y��t�v��=]��Ib�T��&|�uל�ٹY,���R1��ca�<��sg���-X�OemI|�u,����>7*g��sԣjV�U�әR�/2�֙�@�sb�c�a����Li��ɫ�9��h՚����ɨmu��71��#m3A,zq�1ӑՉ��dխof.����~�wT�yy�؝��m95W����{�x��c-����rF���w�o��h�O�U�_�@����òˎ��"��0U���af��]'R�l\j�aF���<u6��ދ��ͬ���B2;<^H��1j�B�s,[ V�UӴ1|���;�����*�I��eZa��E��홛:9p���X8�<��۾ۡ���R͏�n^����6{�Mf]�;H�z���S�z�nS��v�lgyh�Z4"�ݗFt6�J�h��仺C�F��璑���o��y�ݵW<�F_�]��la�s�X��;y�褭�lD�3��Ƽ/��z��uxZ��y�N%:��_�1u<�k�m����K�����\d[��O��c�Y�I���쮪��u��Y�Z�w�������V̛T=���4��
�po��/ѺU�.��
.�ƛ]y�g�{�%��QtD��
��,�S������}��ͬ���ո���?F�)�����Re��d��N�6��8j���ۭ�ٝ�e������nyj���*IY3���d>7%�l"����Kg�Ɵ�>ږ��)�ŏuވV=�e
�KJ��Q:�&��]!'[]����s�c��ٿMǪo�Z.�Df'�(bE࠘��y��+P=4]����oB������n��S����ïE	��������ݐ�m�3Z�E����0%��w���ܻq��l���Wx[��ذ�b�z���̊2aƇNw5�C�ɇf� �ڮ��+q�U��V5s�4a�=��u�5�.N�M���RV2��I�Ah�}~7��3��R�9��ӾEĨk�;�1-��K&x��7�oYm��S^k;<6B��w*�Տ��+h�oOW:��",���Oj����}o����Vnp�m2�T�W]��ʹ��,�/5�m�o��k�yv8q�u�%�׽&��3�X��u.������;�ȧ7j�ɕ&�C�s�n���x��
[�m����q٬D�����G&���͈�LP����O���a���}~t�^إ�vӮ��v�]F��;q��ԏ^b=:���[���^�t&�)��vʃ����kqLpަ9��O���纹�>]��=UO�)��ݐX����Uu]��%�i^ �oXΦ��Y�yw{�R���c��M����M���8�Bƛ�Y����a�]z�u�z�;g�C���[ǵ��zc���$��dx�g�Ry���Q;����JC�pfX�5��ڲݥ$�]��n�]�9&h�$�בWc\�ܛ��M ��՝�X��U�q`�܋�(Ak��+��mn7WO9�o�k�FSF�N��������&�͈]tWn'��T-Na�����.:O�;|l�e��U�rrkUw#��� \xJ;Yׅ;ۅs��-W7)���8�H�X����\��>�t�~�3�a��)���7"��w��ܐ�*�gdo$;v�!5RT�gh�|�P�}�~�N�����R�5�<5=�RE�Y��櫆����U��nf�YSj��o�������֝v+Ъ!�[�;����1��jͻ<:�'�!T���I�c��[�O>��vu�x�1]OֻcX;M�X�߹����A�9M�1Z�S�T�Q���r++��X�v��f�c��5�l�*8���%��Ʃ�s�
�U po���S6�ؼ�ō���nҝ׵˼��	ec�t-��{���O��Xͨ�ͮ0r�?uE�ޤ)R�:������U�"͛���e+�)T2��y�h ���z{���$[[y�Ty��ڴ#	Lzf��N�K}��r�@M�չL
J0r��&X&�WX[2�o=�L������ce�-��YM�|2�.���o;�������r����Mp���[/��[��u��.��퀪�7�����D��A䩔���fogeoV�	�7x����=��
{,M��۪����{Z�,�U�狊�X�ͽy���U)B�B]��&^�r�]๭Z�R�j��O,JkT�{���׬gc�����{ӽ-�����VP�nɮ��Gk���Vj�+\W�޶�|LN���KW��[	�Z�W�5��\T�Z��W�����ء�VPg�՛�'s_	��r�SV:�vD�g�B��B��2�V��by�D�����kEb����O�u�
S�[�ohC�>n��>g�ze�L+�^s��x��#r���3��I�v|�~~N��K�[�΄*�`�&@|:�9}�qȞ����e��D�z�;u{y�o"&Ӎ�C<�y�[u-x�6��b��"�jWNM���Y�^*j��EUo��TFd�Y� �u�T��._ݮ;��Z�;Ԭ�
�F��9u��w.�eq���_�1��;���Щ��ͮqE�Q���85��,ٝ�:���,Zј��ъx�Lh�����ݹKS���e:����@�sb�c�m�3ީ(��d���s�Qgy�����.k4a��>[�R��{�*gQ�[�9�pZ�F�]��gK�1�h^Ppst�9���ҙ3�q^ԫ��v3}n3�͵Yr�����_=��w�~}��-*�/Ҳkk��.�8�{)u��Z�]
R�a��������e����tf�T�ѝ�����[b�etݦ�C�
��k�]��'�5��`*��J3g**v�0;lòښ�����lD�#B�#i�媺f �86��_-�w,��u�7f��L�9k�u�2����_5��<|���bQ�����Rג�b�9�����^QN�t%ī�����\��+ Mk���C�����NM�%.SaoUC7�K��.�d��P�����	'�!$ I?9H@�bB���$��	!I���$�䄐�$��IO�H@��B��$ I?XB��$�	%!$ I5 IO���$��IO���$�`IO���$��IM��$���d�MgƄg_�f�A@��̟\�,{�7�H�!JU�T�T$��R�QJ**��� �JIRDJ*������Q(�U%*��P����T��E@�T�J"��OMR�ZԨ��"T�� �TR�@�PJE)�JR���T��HEEU	*��+�J��!P:�
�����RB��*"�AH���Q@B��*�IERT��D��U���� ��R���"\   #�j���l-P[RҤ���&�eUi-M6�[jʢ�T�-�4�l�KE3��m�5��mKb�HɆ�d���%��*R)���h�T��   6\�Ak)��I�5@�QbZf��M����4YX��U��*��Cehm���[F�R$���j�T��t`�P�hP�B�t*�vi@�D&̩p   ](Q@
(]�� :AE� E� (P�@P���(P�B�
(n�
(P�	�aC��B��]#)V�J&6٦�jѪ����km1��l5Cj�(PEE!T��
\  �
i�-Z���V�L��&+Ydm�[J%����bV�ڴci��ʦ��Ś����Sh4�mi T�c,Mi����*kP�RJQQI   ��ST�!���Ji��ZVʰ�����Hi��2�2����
XmJښ6�cK�Ҥ�j6�V���S*��Uh��UJ*��TJ�DU   ���*+mePkiRԂ��iZ�B��ie��McV�֕
��Kj��CH�� j�@Vc  F�U
�*���TT�� �@�`TZ� ���@ چ-X��j�P�T6�()A�2���mh �`�DJ��"�@�*p  n�Բ���MYf4 3X
���m�H��3�Ua-@ �T����QI�J@N  ����h ���	�b��KP
�)�
P�A[&)AAXM��[5M�i���hI%�J!@�JR�S�  �v�ڦ�cmUUZ̶�c!EZ�aP�XS��Mmlڛd�R�6��[V�e1��DSZ�jPblm��d-����eIJ� ���$�*   0�0&2i��J�Q��ѐ*~�m(�S�= �M$I�U( ��Z*TY���+\ٹ��,��/�8��J�-�\-�>��{�8u�3yP����M�G�I	M����HH@�����$�`IF %#�Vs�Q�b]�@�V��PT IXR�Q��\{�$�M�lT1��\�c��-V=��*bT�X{P]�@�QM mi5�Йj�5�ʔN�E�:���e� ��8��ڶ7�(��Z�&�o~�u$����61�T�5Sp#c�)P3��sLM+�.ō��y�,�
T|,�X���R��8�IN�K@�E�,���KФ˔
6��n�2"qŀM�Y�B8��N��u�D��	i�(��cŸ��%72V�ԳFk�(���j�IP͸�Gh����<�y���ܔ�h8��Od�m\� x�
�X7,�ݳv�4�DU�R�[�o!��7Z鲱�lQ۽�#T�h�5��G��\8��w�2���F�Tؽ�B��N�҉��Ⱥ�e@�B�Y��mmd7�0%���
m�:
[qѣ(��q��I�e;wa�j�B�Lů�� RR�;r��Md����+��FV�W>*����uxʳPlk5��j�t���AE���BJ�a�%QV]�8:�`#a�̇]K�,X�H^n�;	�� sh��ӄFP:�˄˺Y������1���
b0��0U�,�����r�[�������������P��5w�0T7a��T��ٺ<���&j�6����-��f�jaTpD��2��/~;	7�ӋSt�Bmn��xȨ��:��FU����z����pKy^8�j���*�A5X�d&��cu�\X6�9 Cp!6-
�Z.�Y�)�KT��@!��ţ�ӱO]�*�F����N�Jc���s3عEG�$�du*�k�(T�*�F��Խc#�w�V�0����P��dL�NC�ݧNnC�h���i��*[9�=z�U���	°:�yM
�[��;-��ѣw�
��!�25�a��E�M�^�0�,�wK��MƎ��J�[IՀt���Pܧ[�7j��-^�^k���i��P�ۍ˺EФZD��pXdk�z�n��$��YD�Y4�f+�������9Y˱�tX�r5�kR��ZIG��CR6�=ӭ�*ې�\/�q�Ȋc�ܽ�S]	>T2�fޥ��X�M�E4����\�j�xԔ��B��G�"WL9�����a���VR�9l���A�Ӥ�k�M�ź�+fRg-Hֱ>U̉e����D+o�I�Y2֗fj�#A��x���O�ܢ�5��ZED��Ө��	�t�?'���]c��im	q`�09 v��ö��a�k$$���~�Tq�]���������˕6��<��Ӣ��\0�f�mt�A+2r��q��X�������l�Ӡ��&(�*�&���jjK�YJf��{�%$�k?=@$3��J��.0j4�l��Ov���d�1�)큖Au �T5#+�xL�R[��y#�{%㖶P������jQu
��p@��ʊf��8e��j\
Q�V�*ST�׃5ҫ�nƅH���5���n�(j��z,��)1d�$^���R,ŏ";r��WJJ��x-�X���X��^j�;�f��o�q� ���.��7iY����ch�7�;¾$�4(�4��b�ej�:�(����9��,PU�bu�j���i�dŁysL3ik{gCm+ӧ �q� �����3�{XL�2��Ȩ�4Z`��2��t!��V��ډ�+)ͼOu�Cu�#��j4����x\˙C`��k���G,;Z�uY:�I���ӫ�t�n��ɎL��[.�6Bz)����ؗ��f�KF��1R��%��kFVS��j+u3N�̓L�m!�s%��R�&m���rܺZ�hӹN�I(]�t�*������n��i��	�f�<12v�LtfL���S���6��U`J�w%�x�C�(��Vl,�ȴ���͡OPse��ů�=R�5W�-�������m�,*��]=T�������㷐ۛ&v�z�2�u��l��+iF�W��RS��4CE��[��O͔��dL�3Dt`�M��Q���CZf���r�+F8�����
7z̻�,�b&;jVc����N���W)��/���[-��l��e\J���'�+q��غ��eg�C���c�v�Br��*�#N���!͢.|ܻ:�ܕ,6��L��c{Gn��/B����b�n���.��2H�{J� M��."�{��^��-�D팣q* 4�@�nݛr��׊���J��S��2�<���hҳv�컡
��n���o5�d�'�bp�%0��A�P�ݬ���7��HV1�r0�hi����Q]Q0*� 85��.�&��i���re��5�U��0��a��n�8�,b�Qn���O&ٹFR�J���EhWK u��K��l�i�75$�x2�ԍhʖ��u+p�E]B��0�r��^+���s	T����=T�-���T�!�c�4���f='m���p�9���ʴ7F��i̥�%@^=.V���n�U;��D�)Kb��h���G2P�^�?j��(�9c1&\�Y��>���\�,є�&"V̺0&�V�E��­e�j�ݙ	�Zp#�V���I��츣�e�t
�N���.Ñ�`�
�C,͡Yy��%�\���H��vq���{q�"��ABq�ê�;zڗu0d��d;7E�����{�+ø��[�)Q���;W6n�	6.�rP�6��j�)h��u���t��
HdV9FZi�����ޕ�Gj��*����,�wujtֵ�ʭ�l�[��K�!�͹�Y��¶��Ua��K��h��ɗ�N��]����G7k	����S�f�d�)��ϐ骖&\� ]�7VZFh?,��*V[Z26�;�ё��N��V[���ç�-�QQ��3bj�Y pn�,S���(��tf�o�q�U/q�[K�Fe����(�D�df�v�4m�0�X�0�*5��-��i ��Wx٢*Bt9[�Y�f�V��G^�B}����7��L�v�ͼ ��	�T�X���-���D�7/BN�̫�tζUFw���w"�
Tn�S6�z�u��k��L"��W�rdX�ǵ2�C�+����s� ������[��h��MBf��CC�ujP�u�ַJ*ܡ�0��C���^ ��n1��S��`\�Ф#5��q���j�����$Te�90�m����Z��Q�ް��u��ɶP�[j�R���EB�ؕtw
���

�YqS)DPv�dyW*k��Q�ᱮ�Kf�2��j�����X�z��n�����<w�'- hn`mİ�يQ`����	���̥{��X�d$,(l�Z�����LX�Cu���Z�W�҄�uf�6��7�5I1��˙���7��r7������7����[r��
� �f��V�g�B�f�]7/)�.�6���1�H���ok�j�H� 6v��I{P��Ո4�E�Z��b�:9J��S5�W�;w*̄ڔi�yW��[q0�b�N���y�V܁�tffcK�/f�NSs[�@���d�ɶ-T�j����o 8�PCa�cyw{�����j��Ӳ��ki�z�0V�2�ȣA#�r�R΋�M�W��an�m4B.Pss]�ט��������%uwcw��@�R��CU�ȴ�����$E�jB�KX���I�k
wv)�5�"��"G4%�)ѭ:�a�e�[�t��|�s-��)�D��u;R�{��k��h�v�ݻV���M6,vqJT D��C�}�Ѣ�O�;��UO�iIAnǎ�Vj��b�𬔤���;�"�rM��ބnhx_�tް����+s.�m�l����B�:���*�㎛�>��d#^T�U�5�r5,l@�ؚ�̠�Z� AKf
�mkVƼ��Y��㸂50����kNظ�j"6n�A�^�a �+Z�6���˓i���}wm̑|��;uj��<S�l�@�i\tUZ
ޢ6Y"�)m��h����j­	�j��j�f
�@�B'��bѦ��؞5M�%�$nd?fL[��wG�G]�@����j/�R��y�ej�Ԡ)�϶�F��&���M�nhF=������#hX�L�кI`)����6)����@�8*Sx�(��:�������T�nK������u�$=�T��C(��tk-l�2n
!�Sa@P,5B۫5�k)}��7��[�#[R��D�ԛOi�-�yW{d�ӊݣ���Rx4�VN\ըt��
��VR�7,%��kU*��A-ƞ��,n ��J��bܛ�3nYA�AL۴�KH�ݭ��"ǉ���l�ьN��m"!+t�Z[�T���5�f2ʨ5�"�)1�������e��XE���	ϩ8�M����y�p��"Y0��f�t�BƲe5%�W�b�eYi�:��+(s�j�˳4)�[W#����A�`d(M/�E���`����AJ�i�mL�jr�S1wyJ1N�6��ي���l����b��[�Q�^�Ni��hH��-,#z��nQ���eKC����2�kT�`i��J�v���+0ʗ/6 �����G&�Y�^85�t�VԹ�u���R�)����0QpA�����_�bz�Ve(V3�퇖�y����i�rf#S�V;� ����%b��$�i�	��5-�V��];�n�LV+��*�GJE�v�V�kōڐ-�&�a�*�c��#i�����CYOBG
�E�Q7�6y�Y͖�㷆�N�]֢��v���r�Q��ƭXe�(��,�#h�+^ݖ֡[t*:s�(:R��K�k�F�(tf b(g�3��4����I�d,4�]�N1���y,jX�	�yRi��xL5Ȝ�vֱa�i�,,�۬�ͣ�N���%n�q�;z��ܱ,�4�L�SO� ӷVlR޻Z�:���HǢ��me��׉�i�s"��1oB��;)j1��nʼ�7�ŗ�Zሜ�^�N�*X
�"@�Ew2�UХ�qAI�6�S�V'V��ÄS�P��	)��7�&!%
���f�Ғx�B��I��-�M@u��$L�,�]m�Jl�&k��0j�V$ѷ+p���*+��ht�L���S[��td��VA���ih+,E{-֊�e$�:��7�L��5��,b�p�J���E[��)�e�IԻ��� ����@.�}X�IJ�ŇYD�.�BmMu���aV×w�,!(��+)���n�@`"�״r�AĤ�5JdՖ�����S�v����zUm�:P��#�����ݬ�Z�Ћ.��&@���@��5�7�%���j'�v�FJnlx�G.�B������Ĥ��z5=�9�e�(T{[�S�Nc�n�[Ԥ��<��ˊ�e�f��RXʊ�a�Ri{X�a���G���/n��긱	{����	-�w:�)��.��+�YVB4c���"=�����Wk)*dKt�oTS#�H�ʳ�՚`��+qf�؁ع�h���ˉ�hn�q�S�*��J�\̢x@�0�4�6�j �CV��5ᵤP���<���J=����ֱҘn�%Ze�z�4U�A�^�F;y@�*c�Vf����Y�W.���6
��F��]�v��Ֆ��)h��H�A�R�c\X0��AaM4���vj�31)�	�r�m<��f^�1�G�m��mZ� �s�YB���hL�W1�v��	�H���#"^���6ap)y��2�A��ܥa��`��;��h�[ce���OX�F+�:A�%��T7gM44|��Z���Nf��Ꮅ���;z�#
J�!^�I�����х"�ZN�?@�(�[��`
{�c���u+)n�q�@YZk,&�V3�E��I2������b�X���i{m�͸�6Խ����f��Y�"�]F��TKM�9[k������[q�4��cH�j�Zr���Q4�`��ؼVK��뮛՗t%�w)���� �5�Se��YB�Y��M� he:q�^E1�|�-Aq�iP0�X��yM[�:4Coc���(�7Bt**�`JA�DZ���N�&j�XL�(ފ��˥�i:�'�C/'H4����	�.�8���\9N�P��+b;�.z�� )a�y�X���v��p��;R�)N����M2�?B��Щ�.`:ag��۶V滗W@�3T[-Z��.w�vR�El��لmb�H�m�7-?�{��P�X�;\�&�&����fv�~��AS�Hd��i��1F���.�Zx 쿱e�OP�A��eܡ�+S��4;�������5d0Fae�ϱT^1,G^�x\�f����owE�y�]ԉݪ��)Q��`�*A��]�U-h��5f9zDW6�b\hH"��͙6LdJW��5�(��Kn�]j5aq�B�n��2+J�c]��	J�d1�ڷcr��$[�*�Xm��jqE+@+@�:��Ț�8�
�yZ�ᚊQkg5
��
d��ut��05$q�b�m���Tr�3e��Me��r����X�-�u�mӽemeԐ2 ӗ�D,hߖ��XsH�P&V\�Ʈ��YH;�l���u�u�њ�T��+i=w���MpʗDdgJ�lVM��Tl�G���j䫦p�ј6��
��[�T� ڔ�XC{���vX_2�jI�H5]M���2�jBC>�:�0`E���+N,��:����t+\�0cBS۽�k�X ��WޱR��q#��v)�eYi�1<G);��kH�\ځԖ�#/hTSVPM�y�o�T�����Ө������lm���ҺS'
��G��I��9�|�����U�·=Fn�9lD�\��7$U[�}��q*�w]W0Gb����ϖ!7�����B�&fě��s�2��/~�b�W����78�y&dØFuF!Κ�98H��_��ptu�1�Ω�&ͫ�a�/�g���G2���$��w������8��8��r�C�.&�'�Џ2�p�J�-��-h`�XI�l^�7������eJ�'���ȸV����&^�ļ�rQ�����)��grͱΡ��MQN��w鏯ȸ�#k·��[U��c�]X-gqm�j���2�LK��8��Κ�a9hA�侮��:1�)��z��T�g��\2��cg7�B�{�r�3�MV5�ʱWt��^�1 ]��NTݥh��@�4�0��a�!f�]����-I�QDd��m��݋�U4�ʈ����s;��:+��J��x����-��D��Wn�J��p�t�Z�HS�x���.�]��U�����V,�N�o�M^׶��o9��N�h�qc�O�%y�I��xKD���]9wQ��Z�G��L�e'�M��%���/$��D��r���z�a!1�]��E�N�K�+�ˎ��WYyE���7���+Y�Y�R�K��r.�ԅ�®�zWTEX���c8�&f�ep�=M��],Ds�!h����Gm�6���/-̈́��|0�޿��7���%��t����ؓD�j��Ki(��w��h� >�X������e�>tB9��G�X��n�5�x���ӏ_M=X�A�)f���C�a.����K:����KYS��ױ�0�� 5����V`�b��)��OI�5R��[��ɩ���w�ms��uke�k�L�!�����'[����o%�4{#t�l^���՝�ႍ��������Z�I;�Czpp�C��V\xUZ��+9����Ѯ�ͫg�Ly}�W3B2s���C�� �>�K��{�w'��#eҎ�w��\ɧ�J�U��5��8�K����_$o6�7O�:�ͳ����=���y�tۼ�<�T@��:���7y]tX�W�2�6��gh�DJ{
Y]�,�*٦�Y�v.;.�k:��O����Zz+uԠ���w�����%�7,2��"��׬�:(7�SwN���1�\�V)�k[�Ň7m�y	Y݀ш�Xp��kr�Zt��uD/z=y�qo�%(O(Iu`�u}КpT�u����R��m�m��{�����:2o�w�'Y��!6m��9�qЬV���+�^���k��u�g+��� ��ok�Qχ}��շ�2�r��g��dV�v^�s��d(<��^����i�M�L���9��&�^��醢}z����J��s�h���cUr�'U�dU���vrd�5}���h:kkyf�麸<�R���0��+S����QTɻ�^��WY�N���욯��u�S��Í��-���+�o)�g]B/��b�J����IY7���.K��#C���mv_=���k���u��]e����)K�jܽ�|G�_U��.��yH"_d\1oD���������4��:p��Po��L9Y�Y��S��u{%'Y �B��r��Uθ�ӛ�[���N���;�	x,�W�B�C"o�/���֎w�5��*=�{(f�<+#�f܍�6��g��y�j7��/��V��/�1�W��-����}LJ]J��&�*j@�ۻ�t���������.�U���|�Fr�Y"�;��$�G�ݺ{|䡲e|����v18�P)�Mm����%�
����D���3r`�Z�ڜ��dw4�z>����ll����ќOM����᩺nR�yYWKV舒�o2�݀��4�P����+���ݱ�7f�݊�w�nq戢i��^���׵���u\�W5q�jԲ�Ky������4�u(���]%-��\t>��>4{`�-��΀�3̅�T��V^�q�V�n�u���a[�������u���:u�����9��2]��cc�\5S���u��#++��G��8�I]T�����ɺ���y7�DK�a\5{���S�Xՙ�
xt��$��tɏ%洔�tm>X�vn�ƚ])���|��w��M�������2�
�[��F�V65aú���I��
cU���][ה���g]�sŲw2/6�(Z���m��h����֧dX�s׹ݏ`�FZ���ZV.�A�\W"�5`�\(��Yk^����xj-�D�g;1s^�:�WA�s�\��:��D"������j�g�_JrX<�fJ��Rʟ	�o@�Ѽ-��|yΣb�@V]����^�܆��sl��ò�;��że � z�o'c��vV�]�����!jn�GW[���P�3����4a�T�N�r^@���a��V�6�� �Eq2�p_W;ke�tq��Z��u�Y2�Ό�txT(b9�05����j��W�]�L�B�g���l��lBճ��=��Pq�;A��swʊ�q1,9M�w��̱��\���.��L�u�1�����Wx�3wk�w�H�M�S�n��Yq_� ;*Ŧp}}�ӽ�'���y<���ʱ��f�WiN�4���s�TǶ�A�c��ճkL�jm��fu1��kH��U4�]KR�Y�}�:�_ku�5c�m�<%</�2(�L���f�6v���*�7q#el9Ih#{�ggrk����b���4WVV<�KubAʭm]Ka ����.�;�u�a������&�u�h���\��{!�o,�����b��N�*�nZMuD&���:D7�@�;�����LJ�}����mn�WG��� ��ʱS�`�,A���q3u�L����ݏ23�d�-�N���EY�N��:h�@*��s��ER�q�;&�a�L��,r}��T5(oTz��������:R���!L��h�]	W��7Y��"N�P�ȁVZ�~�V��*�+��"�+([�'�Q��}��g�;�HU]�w6:��	��S�U3V�:�ķ�wV�^N4$�A	�}������+�����oZ�\�����������q*�H��#�ؠ*m�|�1*�=�:��=�+q�t��\�vծ��K�7�(U�M�,UҭG�Ԑf�.�*H�f���	��拂�pc��Qj�gC��+W'��!yxc�2����<�
�{6�h��	CFh����bms�;n�b���6�ߖ��\��9�m�x�HK�O+�-��Z��:�J��A�*}��:[x�c7�}��^���W��kGh�X��SÕ�yZ���*�t{espM���b냴8��RZ����m�
7��No���zN���,�r�qG*�)��v,}V2�c��tl�]X���!@A �{o��Lh\�ͭl�>�y*t3�v�vjs��4�5�x�.N�3�Bo�sܩq�l�z�T�c&5(��q����#�H�����պ���v��Xs>q��9n�wC�N���:��;����(X����Ŗ��W��r��d*��f�u��L6�nR|��:Qc���pW1����t�����ֲSg������'�P����=׫`ik��M ��wR�З�U`��3��=V��ڜM�=P��;4=���V�.�y�U�SNnY4η�P�s��.�$1_wm �@���"U�����������&��Wڭ��Csyi9-�E�i�# �+9��%Y��{�eoW]��H|�'.��}��ǲ�]���T���0,���u�u��s9m�SV���@��1�\��C �_R�máܵ6�!k�GMo[X��\�۷i1έ)�2M]ZΡ\LnL{��z@�לb�n�^]\F��Ճ�j� �v�J�!i�_S��P�e]��Uˍ�1ѥ�;)�P]�kI[�R;�a����I��:�Pr�=����s�
��}��Ќ.�iU<ix�����J�!ni�P?���� &�K���:��h��s,]��j�1z���(�S�b�%6����*�����F�8.�ϡ��R�6bT�Ո�l�B�ECIJt,)n�̕Y.���}E�x�sf��]�7�+�6���b4>��uo����S2mΒZ3�n����3�"�=��F��,;
�:�����"{�[����lY}�Y�9�<�Q�wC�8�F�����Fmli�ۭ�{)YF���^R ��VY�`Ic�[+1�k��@cۇ��ncz����כ�`�Ҝ�Y�R}���	g�8r�bPl�a.V�>��3��hI��9��`���vՙ�+J+���ݧ"�6�Fp��*�8MEÕ�2���#0ww�[�9r=B���Dg9j�TO+���+��WPV�0[O^Y}���
#�̑��|� /�)�Q���AT�ν���Ixs�J�ֳE]u-.�5|g+�!�:���2h�}�:���l.�:�Jn��oc���RE���� �WՊ�r�L {[V���n�]�K9�GeǦ�V"��g0]��]�wu��k*� +YCl彰zRX�|��]}>�B��Se��$��a���s�3��}�P�01֞�]E�V�|�a�pU��g*�-���ƙn��_V�x�;ޚ;Z��*�;it�^V	���fr�y��t ����f�*���s��)�5�.+se�1�1���9!��-:	�X�J;��Z53�=	�H�;�� ��G�N��Y�D3���6SLi�;��Y�[��d[��,�):�R�-����1c��#��]����V���S��.k�iw?��)9�^�YYG٥��Bd�Q$; OGK<-b���B�����VaE�-X��Q9v�Q�����i��/�u0�gs*`�5��6ծ�0�	kJM�5����� ���<E�s�"�$��M��fu�)4�c�pɷ��Cm�7+ם��ԫ~n 6�h�^�+8����Y(�X`�w�F{�A�U�t����[�����j�'2��G������_�o>�'v+k2v��З�	�휃�*��h�Y�9��b�d�[:�ӝlt�ܬD�쏌�e��Q>��KR�Gz�[�����4��͍��N����s��!�]E���7n��j�e��:�;�cY	t2��^�lЈ��N���9��\��0�5Ӟ��m��C6*Y}���`mb�r���[g�e��mCd�����k�rڹ\���Ѕ�������0v�-��j<�6����� v��\��ʺ���G���յ�0ѫ��B��8KZ.�Mw5I��.4�{��;j��y׌n\�띗Wc[F�a�Rk�^��)���b�&v�mI��RS�G8�D�T�wu��.U��L�w|��is��/{�κ&�)�#ĎF�:Vr��#��&�]���Q5�����;*��G3�͢�ε\f�]���4���v���4�w%,(r� ����[|�
�hR����s��
�n�m=���~{���s��;����GWwWvZ�f����\)���)8�T��E�
ˑ1��љ0����H�׺�Uͫc�M<B_ֻ6����Fc ؆k0�݇(�ivm4n��sBq�Yz4�cU2�V�w���2vc��ϻ{ =����Lh@m��]]��M���I��hi괵�h(g֚��K�*�}V,�W�u9S;LV��G:��mSJ�����E�+2�)�s1f;�5����u����8B����Y�1.�Xe� ,�P��LǙ5�/�Q����=M�O�r�����.�T]�[4�"�����݄�B�:��F��mk��|nn�+��Z:���x�^�����DJbkB�eiZ���� ��B���;�z�|kI�ǲ�Hf=�"�k����\1-@s�*a�3& ��%��0�	'`�b!I"����@b��I�u�p�#Ou�@v �p�3����/��&���ھcUv'���.fJ�݉Qְf��#ޤ��ޚ6]�ܦ�'���CV;0�*�u��K���H��޾���o���
Ⱥ��*f=��rgp�.�_v��@�ݒ�p��!�&ORKmvg��J�b�}��W26k����׃f�Z�Kkc�)v��*^W�=XxGFᩝ�r�a��-[ԦmMU%��l4%����7�aN���`�����ĠÂ�ui��h]79ewZԲ�f��e�p�c�洜]�:��[�t��Ts>�����1�z��|h���Fw�a�g7t�J[��$Lż��Pu��c�Fի��*%�7��p 7v��S�_o7k�XI����=�}W{-Σ]��h���O-�(���!{� J�
۲����_pΑ��Jv7eZ����_kpE]2��+0ek�X�(Ӄoy]@�eq�6�Px&�0���SPغ��J�$�^{xh���m*d���������}���"v�O,�&nվ)�C�j�9q���6�u�=�3i�|�M���O��:�2(͊��-#��t}w��u���;m<����E��6�⑋RK����B���u��X�M0l��ً���}f���7K��YZ�gm��V�7xm��^6ZQ������z���	]î�d/�4wU�W���96G�Z�^dީ-�>b�:����A����ӎ�Dzʩ����x�Ը!i�W�i��nBS�ދ�4���F�2ӹ�.�^ �}e�WG���UwR�E�p�(cf�Ur������Wԕ�P��uib���75c�����s�n�|X�\s��� 4��=���d��Q��:�-7�Yx��А��íŗY�(gs�?y�Ё ���$��	&{�3=��_9�^u����V��oj5���Ӂ�����𩵰��]Kj��\Uح�T�R��p�F�ެV�$t�t�lA=SV�ֹ�q��3� �s�t�_<[cK��mZ�pw�EZ4�i����sj�d��q�l%58�㊃��ψ��]s�Ӹ,��ZT��EJJb�͌=����KܭW��h���	��k�м'^ �1�ms�� �YLk9w2t�[ �)��|��]�!���K��
�u�Lں�[%�7%�b��P�u�����C�f-շ�4̑Ū��ًcBhZ��Βe��q����)⥦ؘ�U���SKF_l�))M�Y������}o�}�;U�����*��]�:C�w[�pE͘�Jydڽo�
�3S/1�0WI��)�ZP>Ǫ�r�#7���P�z5P��ms	�Le��9e�����g��� ܊���_=����t��b��!#����8��k]d�I_PP[G<�2:�T�õ����
��+(p$1;��Ԧ&KWyL<�p]����t�ij��T�U�죽������ ����]e�A�qTz"�7O�>�j��C \5N4���<E�.��ܱ�s6����f⥝r�sYל:�G�u��]jH93+K�;��
ӗ��/I�<�్��m�<�:�s�ܓ՜�7E���\I�y��*SF��+�u7��t��gn[���d�(�޸�j�Ƶ�"\��@�o5�R��(�E�bμu��e-��w<�[�SÝ�R�m��ܪ�d�:��of�����WL]�� �Wr�f�.�[��p�fU�eh��c�Cw}�u_7�<�Gn䘷�)Q�3��v�;w�/����Y,��r���0���t*�,͝�,�V��XΫT���%�� �X��Ii^1Ww���2�Qѱ!�$�n��%I�f�����Q�o,Ҹ�o`�բ��������R�)
��#��n��0'� �đv�N�e9L�O0`�e�镻������靤 t��Y*e�͇c�����Cˬ���E��|���-Sv�b5����j}�W]�i_TU�"�� ��ۣ�m^�kWg
��\N��s�}�'@]�9;�-��1×�OVP���U�;@��]�@�1�����r�dL�C�r�{`��ˤ�z��z0ero�Κ�+;��u�R+��]�+2���M�\����Y�{�֬�;i v|��ݼ�`	��J�dk7��s%iè'f�0Wj�#�[����Ug7����ʹN�44�w���Eu�L�y��(��Wy۴��/]V�P�e��]�&�Pk���\�ʟV�u���n�Z]�I���r����65�.XiU�;��kI�	;7$i��w�h�r	�ηv)J�����wvx����v��oz��Z���n��ͨ���N�3s���r��k�f��4_$��dꗂ^��0N|����hN�ĝ�P���!��v���-��@���l��͕������Wp��k����+{��k\0`�ځ��W��6�p�q����2�C�p'�ъ�eKt4G���}�m'���:��j�˜�ģ�[f�:�P��x��G ���BR�����7�������&�{5�ѻ���c?N�ؓw�ü9��`�>�޹&�EV�w�r��X�h�v]ܚ/zk/6�LR�`8�v13�+(�|�$d}�J��ӛr���R�#��n���q!gc�P��Mf���/�w�K!]��y��k6���qՂ�t͕�G0��N����۽aM���c	��j;��\9t]�}Řv5׀�h�͍���҂Ckl��Kj�%xk*[(=������S�B��|rAf����	��7.����Ζb\y��+iP�u�^�5�Əf���e�^ٷ�>�U���hK�Ť�
�u	��_g`��#�֯��r�u����.��f�lH�Ƅ��\���s���獪��Wm_^�5���
�(v��v�l�gG���$����C��si�w
}����H���1���;�����條Dp�ԇ8�J�H;�M��ݚX����Eʮf^+xE�WCC��>]!V�⬚�)R�:�nn#�pa�s,�)��܃���_!�2:��u�[���%9TR��Z;����"�.}����p�n1XG	m��F�	V�}I��]S3U��%fk�:�k��:��)X'��92��ԟ�,Cy�/����rR���7���Ʊ�y�/����������4Q��;�6.��; ����v�r�l�,V�X����B��V ��+��ծ=[�x�Vj�m4i���Z�B�,�\��f�t�meot�&�C��(��^Ȧ��r�j��T�`Z@�8aÕ9p���jص`��y=�%C3��A�]WL��&0�uzM����b*�W.��M(�����ȥ�ܘ���%fѧS2%	����/��ޡ׮�vO`�Ndg��!���;xc�\�$D�!@���j�=���Yɬ�e��P�j*�����x1�j��#��5a�'��wWG�qee��뻕ܜ��=r 0v�CGI�"7�����' �)�QT{�G�e�׋J��Zr.���&����.I�J��t4�r�Sl�{*|G=�ܒY�V���˽W4��:�iqV�ϵ�]���������G�ˮx8|9_ȸ����r}�k�������vÞ��nh��t����RM/)-gi�p�=1k���ARۓ�ֺ0�_r��E��GhN0Y�Ba��)t|�%����мꆧ�
�(Y;��Gn�v�j�0��f�㒇@fN��G�̜�څ��U�O�jA�К��颐�ۗC�r�S<X�2���x�ؓ�:�b��W��E�ڜs9�vC1�)�A�8�6X#8����I��:��Y�v*&-�=b>y+n�����ב�C�Nw�k>���D�+pE�;�7�8�bp{�`2kmq�Ӛ��e�T�%�d�w�W��j�pa�x��Dҳ�Ԥ�	/-�x�%�m�;3;�_˕:��V�[�i���++(��wC�3�����J�����5�&��A"���!����R�ټJ;��[�
�M��8���[j��1v;�f�c2ڗı�L'��>I����^!Vv�o�}��;2��J�zuj�,>OU��+"l1Q�S�E����i�( 4���d�}���W�bGb��0�3�X���͌3�\����O"a�a>	�eރ�x���pO�i��on(��.\�H�Uݭ�LF�%\a�nb8':�0H�7�o��Ae*`�
&�k@�o�C���;j���U��p'4��]��y�%Ҭc+�}F��%�ѹHm�h]��z��W�M"�hfXt�/�	�왋��9�qڅ�8*A[�;�N�����O��t"�]�6�G480�4=7]�ը�@W�2�r�X�h���u;�����u�.��p�7}��l�nF���J�XtN_o�c0oT�1P9�JCR�w2�Q��f�\E����l*ĥm;v{�Z�������|Ř�,��������C��t�eNиv����gXB��+���Ǒo� ��XR����Ra*��]HݓH�Qf�J�M+Z������H'�6��^]�w��+���w��j������`�l�0�Jh�Sr����ٻ+r\��;�����ɍ�@��[�P�Ӌ�Nݬ]4ZT\qT�]�z!Xii���f�)�P�7���KZ�X�,���n�'J�̖����������C���x^��㴥�c=3����y��.�V61d��Y�F�
=�.ƃ�ܫv8V O,'N��[k�>D�v��ͭ�ܗ>��+���~�eݩ�2�4�V�����uesNn���J6����47�E�P�/�G���<����JL�uƻ�)��o��׻��Q�X�+ip��a.�\@;ݬI]��ϛ��ָiŇ��s[[��;t\������7V8�hR<DwY �fݼ���,��Gt*%)�&��^f���H�=��kkwm�|*;A@���1����a���n�H��H��=���`��v�K�_݆B��Y\F��:�"}{�
!I��+���8Vi�Q���#jlW{`eMջS*�#ևb����Y1��t�ܩ�7�V��<�V���׮����/��蘛4�U`)s��ǻ���ֵ�m&ֽVvD6+����Y&��\�.�[j��\�4Vk0��$92�K]ڠ���H;�8�n�u!�|i��C}����]S�Y�hF+:^q���H�R^j��m:�Nf*us���'+��fuc
�i��S)�[�uib\���f��e4�GT��n�:�^e�v��h�no��SF6gn�XO法��\�zkI�ƅ�{�������t�Ҭ��P��hm��X3;��g\eD:�����m��qN�Т4v�ᇲ��n%B՘���vF��(}��xkK}�������撄��\Ԛ��Y�P�1�6�'L�YW��D�����:Wu�=�ym�j"�׈B��(��V�5��{�����܋�\��'�#�� юݰ��#����6��T'L[���0���BǄE�p�Z�ϳ)�5��F��y�25���N_U����l��"�Ywf*i�9�v�z��q��lZ��/2��I>F'����m8Z�[ϖ��'g�/�w1��Uּ��7���� �C�hG���z�۳��pU�n�t�ѭ�r�\�6e��;�@=��J��u7��x�1i
�/�5�$w��y;�����L�o��T�)n��K���#�I�2*2��j�Lx�1�^ٺiߍ)�9��RV�eҼz��^�*谇>O�tn�m<)4�]���KU4�k|u�ۜ�u���[*7f%>��a�r��f�}�µ�5���WLҐ��o,C��R�t�BRN�G+86�}*fLp�}[���j���O6�3\��,ڍ`C�t=MW_i�����	���
"�!�r���fi��63wa��iG�ܼt����7�k]Ϗ_@ e���Ʋ�G�=ӻ	{�L����t���ݍ�yS�A�3j�oV9���4qV�&���h�.�C�T�sj�fM�����H�<i���c&qL�F:����k�{�F����X\�>��=����W!ӻ�h���U��-���!]�z�&_'C`yKb�p�ύm_�E5�W+�����gi�fL�, sF[��^=�Y�Q����* (����kO6���_s���Ү�fN�uJ-TV>H7�֣�w1��4T�������x�3ZBu/>�ܣե݁��V�ܘ�"��9���t;������Ot��f]v�²76͉D�w�pw�[ ��-�{e�|E=`s�X���P�׬�B�]��;r�-)�ge�:��O]ZQ�V�>�\V�d)�p�v��B�˭3WHt]Y/�fj��
lF�&���e�0�I�������slƲ�̶F�T$m��Ȍo�B=f\y�Q|N�7�:�J��}��^Ωk]�C5	F�9��Sζ�� q\���K��N}VL}X��r��.th�{�	�zڲ�l0�6�bG�0��=O]�_ܷx��'r�/U��7,*�*cF��PO/4k2�2�DT�0��do[s)غ�Y %��U�]���a�E`w�����Aa���m�j�oz��J����O�:�X�f�6��b�J�H�䢮{g+ʾ�yI6`�QQ�L�rƽt�s��.� ��8�.{:� +qGm�ζ�����cO9^����z���՝���ʛl�D<x0 �;��f��
yz\Y�/�ѬjS·�*�9=;���f��%tK]�ʋ�r��W��:�t�8���M�++Q����mvop�'a��+:�=l��Rox$>;�wS ��YƗCO��9a�&��A:�%�
��7N��=�̔�����^�� e���Z�J�uۋS���z�
�����)`�\1�qW-V�ɫ���T�ĳ��k�Υ}�P+�걭�Dk� ���R���v�X�Z���ļF��;N]P�:1՛�;���G/��� %,:�� B����m��H/�'w��K��.o9qr�U���[K��d�;�&Q�l\;��yբ� ��d�2�\�+���j�5�0�premfi9������X��|i-r�G��5�w��sT��aKy��I�:��u+��B°�
PTb�C�MU���*�2�k�]]>�
7�ʸ��\j\ TkEѶG
#�Ko&
�t݃6m�Yx��rrW@M�C�V!y�A�ѐ�	C0��o5i���ͭS+8 ��MT��o:��Zu�{�����m̚P,@wt��3����p�Ю��S���n�S��hQ���g8Ρ����@M.YJ�mA*ݺ%�̵�1X��>��m;��b�#�w��LB��]yO����,����0&l
�Mڽ�ħ�*�[8uEW-�Չn�ź`��v�sŀ�I��L�&����os�{���yWNak%��t	���nI�NR�H��d�c�$\˫��9�tѣ�,s[���a��0ni��m�r��khobݼ��
�o��4����N�hs��G���ACX]��������o֯+M����Lx�`x�*s���7�jQ�$�Zqm��	�R��
I�+2�Jf�R��^��hŝ�ڮ��  �h`ܮDl��3/�rv��|��5+�` ��/�陕�frMU���*+���Ӷ�A�s�
i�lA|yɎ0;7M7����@���ʏj��#�
8fe3W������]}@����vMl���._�}_}_U}���Y�Vy�U����u+F;���2��r���i�Dw`i�mn�}Z�|huN�H[[}�Yg�j��*b�Tm�����!SEK�1d[ќ�y�J5�d��1�ܻU�����cU�r�]�i�K���hb5�Y}X�+ ���UĊ��'M�T�ŦѼ��@+.�GL�HJ`32nKg���B��2(�&��llei�(���t@Sq2V�{ʯ'<�6�A'�W6�x	�����V��lS�ō�y�FBvs��ۜ�R�o]����>ݸ5�8� Z��ڨg ];����J��@+��ؔ�wV̊����K���}�%Jv)$4�y��*�iV���JÚ�]�ܶP87E��S�˷�*�m�zK��ɬX
˾ݜt���4�]*� ���%�^d�z"�]k��ir�ݿ]�@���k��R��;��]�u7�&m�GA��-���,�/t��f�T���\�qT�O����n�7r��1Sʖ����uO�!��ao]�wR�)�Du&02v�.��>�A>�v�������q����[�W�t�����f��H�R��Z���ޓb��\U�������5`�-=Ma4qr"��11y�k�N�j�Qn�r����u���6��(��M��Yƶ��;����G�7�����ѕ����V�߮;~[�<�i��19nv���,c�U�X�(�Օ��J#R���Q-��D�Z�J�e,QQ��DYX�����h�Ҫ6�%��
�e�jհQ��*Kmcj�V�EJ��j�%Z�Z,m��U��YmE[b�ch[YJ,���Z�6�Q�6�*�Yj�*�mQ��V�H��UX�hV��2ڢ���[Q���FT��lV���+*
�*���Ymb��*(�TQQij�X�iF-([B�[kcZ[lc*UV�(�mj���(5Km*b����Q���jT+
�j�+U,hň��E5F��TU�V�5�(��Q��ĭb�����������������B�F�AUm���!Z։Z�D��%-Z�h�(��Э��l�Uh��V����U��6���ZZYZ�6�� �[j����[A�[K
�mb��b�Ҫ��F�cYm��Pm��
[EP�"����*-�F"#kE�յZX[bԭ��eX� }-<Gr�����h���S��7���f��KSMI��Xp�㭓Tn��66�)h�VS��]'��NmoV}�.L嫯qQ����������
�O/Ů��E8�r��+��v:"j��%�ϡ��L{�v󖰩�X�^��=�'�6%E�˝��!쫑��Y��]f"��<4w/#����,T�_F����8 ��s'�A�*:A�2�����ڱ�(Ew�l��\���k�]����ݨ���P�qQ�)R�6d-2:uMD\཯r���Rԛd�w�hG�����a!��C�f}=ˋ���:���AǨOTB����<�z�M��]�"e�9�a�<y�f��Q�!F���n��Eqb<D'6 ���q"!�:�ڭ��-a;9['{�U�ǾIVC��V-��Ѓ�l��+�����!��
��.T@u�y�ngQ��=�Њ���&���h �%�_I�ī�|�O�Z C��Bk�vn���n��+[r�,̼mp٦�.�����%����Eگ`T���]C�>N)��?XL�k;~=������
)����� 4"��Q�i������8>�7�"���ߺ���uB���3b�j�u��F��yu*9��r�7�Ƀu�œ�B�ʾ��"���j56�}P�(f#]��+a�6��� ;n�|4n��(=ξ�HE���������c��".�Jn�|dR]��#�N�ɏZF������&[uu�W�i�]�q*�@N�����6f�xv$������P"�����ᗢP�0�Y'{7�Z 5��v��1T9#d(�|�jB�ddkvv+n���1�}�������:�A݉T�щͣ��2��Ƕ)C`!�߷��~Wj<B�s�p*��<m����۞���SI��hG�OEvKf�`�Uюo�T���G�Ӷ$t8�!t��Oc'"����zҺ5���C���L�7\��VrZ.�\�S�C�J�t�_zŵ�x�Cf�È��p�m�-�{f*s.2�w���X�A���h��b�\E-�t'����k��鞊&�o
��d䌆	���#��Y3��P�j�b�~K��_WNB��b���2�Aj�q��VrV�Q9cX���rJ�Rc`R����uϵ�]N�rb�*Q8�1\;gu���l|����A~� ������ ����hi�+����`��C"EoL�=p�]����c�b�A݁Uca����A�����ma��g}[]�=堭������^]�;F=��%���z@m��F��Y�d�Tk��h�=5qF��%X����m�(��G]�����_�5C���v��,����`B-�Mh�@��&�����k§l�t�;ݽ1�kT� �Ys
�8��t���Wd뻧f�*��+��ʀ��tRvk��������Z�=5 �����֗T�7#�ۗ�xdE���2���%�Ȼ�G�'d��9�UFC��׋8rxfYS�fS��AU����A���Ak��-�2QF���!��S��Kt�FYꛗ�	<��E�F�,�]�e�Lq=�`L1Hp���9
�
sP�E	�֏��1�Y�����)���=�'�֌���~2�+�d!�e0aD>G��7����^�=ƒ��%ʘ�s��e�5�������{$��V�v^�A�F�
xAy@��}�36�Ϡoy5���=�b#Ϻ��Ǝ�5޼,
B+��1Ҭ�{��U�V�=#���}��.��`�d8�u�9�t��	_{��k�k�p{fR��2��d+`�Uz;hEç9h�d��̺ĘS< tnϓ�7n2V�ɘ����*'��~�?m
��.��j�=;#����p�pZs�G��GKS�ٷ �Tcos �J-�y�;R�L�D��:±L� ��X6�Σ�{�9�f˷�2ʭjN���feoV����4���Lu���6�yj��-Ճ���ol �=�-�:o0�#�7hڅ`�8[����uٝu���:�8�!�n\Y�z�����0�:p�u�+�t\�3�V���$D�{`��[W�@������"���X�I��z�%μ��Ud�ŌL�M���aIq.�nl�g^��:���=S+5���`Ճ���8m�=yt�pz�y���.�A)���m��7V{�3�f?����_�:���,�H����<]���Z6r������F�f��S	]�҃���B�;t�hE��������Q��"2h\�0D�76>���򮶧�Bɏ������ JS��)D:0�LੰU8�(Wq�/��DYT�Β&3�^?I�8��G9�Uԑ
+%���28�U{x�:|z=���?	)u<�����
��ČM�ܕ�k7Ϣ���:��<B�YT����8HF�b*I�ٷ1 S�S���Ɇt�U����v���Ӱ��+g�Ʋ4���l^;>�전P�.X��f�^�7�6h��ƣ����_o[U��X�]�b:�`}���v�`�����1�&s|�a��tMr�'�/'��5�ws%�zݖ2�{(���������a�}Q@�z/!~�nb������-�ˆps�	��3z� qP4\����czolVb��op���y�����VQ�䕝�j�˝l����+TDY��f�ܳ&���rϱN���'W1Hs��R�Ę���C�fmi�L;�͠3z!R�_rW��j�q��D�#IֵoR����ꛦ��p��ݪ�J��V|����ׯQ����`�=ǭTV�otw�;5�0E��F���1 ���2�F�����<eCX귘��G����}���1s �n�m>��v�a�{4���>>�P�޲-�NÂ�F)�T6'��Q$<GZ��'��<�=%zp�{�=P�&\X"zEjptڕ~��dc�29��y��Q{*l�y7t�mF��qw��m��D��mO�dª|�hu�{]�����`�E�3�����Y4Ƅ��H��o)\�ȭ��ޯP��;�biF"�aA�e\��rڛ����{�ʒ�ƫw��F�[�X{!��T�H��9��Ԡ����뀳�>��T�Ƚ���l���vd,\��P�R���l���K�4�X��ޭ�ms�P>
�Z`
x��XFm������E�lGL���G�_�q`K'[L�LY���*�S�\El;!��L�voX�p=}��M*o:N�K�h�
4d�K}[�ň�����/=;�Ð�`wYP�ZoUrb���M�lŀR1+E��[�U��zy�Q/>W��ܡ���u	��wwN�f�ӭ(�P��Z��u�^�p�==vO����j��$�(�˅!��3��N
�j�(p����;n��iOq��{��ՖZ���!i�cj`�ܨ�&-;��k�,z��R��)�ˤH�b�ٰ�[����QP}}j���r�@B�P�4�Gm��48{}�c�D�;s��J�nǜ72	���xO�(]��x�7��_NA�cu(�������=����&"�ܥ`ߵ�:jۂ.�p�M��ڒ����U�'?�K�9��K����۳�n�aM\.��_��|���>xo&���;%��*�Tv��G�a�%#l�z���]wK��jJ��5���b�i�4M�Nh\d ����Ė�����J�ww�{�'������Fkԏ�+��z��1T9;!D"H!V;��\��㧪vlF���4����f���v�S<uP��S��!,��-Z�Q��8��8��ӳ{yH�j�r���L�B����Դ_���:���=9h|[G���K\n�N�Y���VC)��WR�S�0t�aWGz�RU]"T�Fg��B��F�D�[��z��e[z��ܿn҇��v3ث<�mH�#�P����w%�Y�j�1�y�v(��L梷�(�P�=rL�y�p��N�jm���-�h�&��9���۸ �N�W����	Ve���E���bT�u	z�ǖ;��;4]��p���\��0�r\�e�z,�[g/ �˥�ZgT,ή���sԓB`��L�\J*^M�
,��O G�CQɞ�*�A��Ҭ�ĝ�Bс���C��������=g�U;`���0�@;%N�1�)q9�G\����6!91@�TN�CZu ����#��w{~�W��H2�-p���xԬ�^�a�#X�W7}��(���i�^��D��x��U$dHbr2&"�L�
� \�q�A����'�G_)�2�M`�X�^Uj_�ָGu�s�W���r8"���e?* #�3���]R@XC�?*�i�7��WBo7� �q0�у���ײ���]J"%� 2!S6�L`�!�EاOG�/��f�*����=����[�_�f�o/z=�Ue�6�j�<�Vd��Q�!�Юsޚ����̵���}��H��<��t}�ݜ6��1�0@�9	H�5�P���G�O����w]K�GU�80�Įnzj��gV��GfW� �@Ì�(�@�~��M�L:��eX4�^�k� ��+��މc��O�lQ�4��I�[�m�Qc�(9ܝ��3������z/=�v�:�H��m]!#q�1h����`Q+�u��K�l��f@�w6y�$0^e��#5���d��Fr�L岅̩5P@q�X��dڏ{��P�Cj�)%�Q�������'*N���.u��n�۠*�9�r��}��mNİ�v�wt$��^���E����Gb}�
a�Kʘ�)�u��*�1
��U���l��:E��N��6/e�e��'f�{�%5�����q��혽��h��Z;����������-����S��okD��Bn�,���L�FV�)Q<�*��"�^�� �>��7��Þћ�&����q�ٵ �U��"�Cr���L�K�3�q
�D����3���Ģ�`�WP���֫���κ���d���Ɛ=�S��$]���q����@�ՠ7���[5�!�~�ê��z�h����]u����d���G�ݩ+�[Sب���E~���D%�)}F�������jѳ���S</N���ӥb�Jź޿+���<�e#1��,���y�H��*�nsI���}�;q���όC3���H�NC�� ZgM�N$RAn��`g�c'�U��vn���,�y�
��T��;�O�"lo!�F������+!�{��wEA�@fJ��Be��ݔݶ�.7�E�Ӹa����wB;��^�fy�"��8�=��UCX�F���t�8�R���tiF;f��Id��:�-�nu�Ui��T/s̄D��[�Q74���\��6�I���u�e�b���;GT�­䧕��/�sd��^�:B�G	noD� D��o"��&cfØ�2j*�5�x�x�1�v�S�Q��bkN�5��1Xؼv}G�A�����("6���K&��L�����NY�����e���,G����e��b/25u��9�Kg�3�/��wv��n�3�r�6<,;(?r�K�պ�xS%xRñ�>��[=R�e��j�	�vg90���Fl����{]�v�$s�3(X�w�����1��*��x��fw��$����{'u��jߩg]�m>� �*�w9��ꕏ��3b�i�\��&Y�Qy���*�v���z��m�75�E�B�b�R��/�v9��<%WfS�W�z�Qb�n���b�1i����ۺ��`�".�t�����S���(#�cd����F+S#�͑nzķ���f��MrTL�WjU7��t���c���;C��d:K�R�������FK��|�JD�15�7竊�=����z�������y�1^��z�8�!�D�
�t88A^�؇��ה�a�����o�&x�s� +~��6^�ѤS��a[B��
�//p��
���tX��]����f����|;i5Ѓj�a�ϸ�])\4\i�b��=�6b*�A���Z$�sY��4�꒓���/��ؙO5Ջo/9|�efwu�-$��өr�.'g>��G��,+A܋R�H��t�H��P|1
��e�Dd�Y5�ѮG'f��Mq�:N��b�lt6z�ێ���P���Ǐ�R��|������ ��%pW�%#}4^�c��*Jo& S��p_zϪ:�,�m3�1~4zju<�w�R�νSJ ��;W��F�z��D^�:6���-�㷻�}W��}�j��߶�/"\�.�Vgo���۳�ѬRJ��j�c.*��X7�r�b"��f
�\���צ��7��^X�O#6!���{�&��u:�d�by/��9ؿ5��b~��miv#���r�}��ܞ �h��m�R8G��h�,����PX���'��v��;��}��6g^ц ��nb�; �u^ɨ692CB(q�:zUnȨ��U��~*!s��#�i{GrU֡/�����+��a:##cPٚ>xv$����1�v�	}5�4y.\�r{���([�2��E�3ЄdUH!D"�N�_�`������
��BQy��l�k�~|���T6��w�Kz�=��sW[������������޾j�d��If����˛|�1����ı�Qc��<A)͑�|2�y���*�Q;Ϯ�g7;`G��5
j�I.kӢ٣�	1Ժ�fd��J^n�u$� _Y��G\m�\��ZdfU�N��ccwQR���U��h�VFe���L�xs&�4���.K���.�i���C���w+E�f:�$^q���H�Oi�rX:Lw����m�цu�gn�EN��(G:��N�ؕȧf��*�Ž�`��������i8x;�w;�^�I��t��L��׺�r#��3�!C/��XM���U�Z����,��1��t�`i����J�.f\veA՟m�y{ZG2o��S+qmV��1��Սf�K��x���!����$s����vu��llz��D�w��1�-ʰ؝'f��A�i`j�K�W�)�]\�ż��Cɗg����W�JCcp��e�9��d<�ӥqژr�G���s �d�K���3֨�+�+p�erǗW�ͧ��k)��G����\�I8A�ޛX������X.��|d�ɕ�pfPErwfrh��Ç[?ƍ*ac�H�6��|��w̉ǋ8]�2eB��i�R��*�,ix=V��\�΍5W����!lF����d��6;'bB��Д�Q��݂Kv.���zխ��a�C2���S���Iw�,�i
*;(-s��cK$�	�n`��Y��m�Ҩ��VŢv�R.ΊL`����Ş��(�P���U�ʏ ��ޙJv��U�!0��,�Q!Xv�����,&�sMe^r:��D57����k�*.�N����4?��k�Z�;1V�-�ój%�@�o+�ÓP�8�oL!��uk&5׬��Vg�]��,��Ib��8K ^����h5�YhC�`;O�9�i�����H*H��		�_�4tl�㫇M(�3��M�b�C�FE3\%K��@]�n��R�ʇp�y���0R�͗2�*bܢx]c��b��}��rg�5	����:�|3C�y��U|������1��Xu��6>4���C��@k����)��A�3�q%�̞>��⮲�=&�{��Iy����ǝ)�LJ�;�)_@�s&>Φ�/_k�;)cX�ۖGӕ��Э��e�A�ç�G[��1��.�сa���/zti�C\{�˹j���3ՙ�;�[�ܚ)���@�霰EyIL״7��	��m:��@�m.�;+eBXO��Gf#�+�����B<�ڿ����^:З����	��R�]�U��])-[0o�Jw�\�6�}CiP#2�U�,v��5�鯭�.K�x�u��$^nK��ə�!�o���h�m��+7P@�;�kϷ��U+b2�b"�B�Z�eDE�cE�kYF��dmD��#eKhTj��D���* ���R��R�����(�k*,��"�UV#XT�%@DQ�kT�e+m(��m��
��B��kj���D�ѢU�XV����H�j-��mQ�Z�`�Z�d�B���"�����DR�J�((Q��(�e���R)R���,�*�([k(�-�ZU�)UQh�iU��b�ň���mFR�"����EF�E+X*�[J*�*[j*��*,��Z*--e�Z�(��UF������E��(���-JŌ-�RŔ�� ���Tb��YIX�QV�QTYKc������R�U-�*)m��
YDh�b�ՊDTb-�*���жы"�PF���b�Vh ��IR�JֱeEUEm�ĩ`֢�����m��6Ե�*T���DA�,b[k(Ő�`��2h���R��DUV"�F6��T���>y����7��c�e��R�Y�����0�B@�Am��]s���{V�8,;�^��H5���ҽ�
�Bd6߆9����f����O�D��]�<�;il?`MG\��m���}����<�C63�rWws�,:�z���L�O�z�����~2������ONB}W}��]�U4sz�0nX�n��]��BইL�6�J)ʫ�X�"�z.#6�b�o�vZ�y;�"�������;ħ3q��XS�����ƺ������q��d��4�c��os�����6�8�Md7�u{Qɞ�P�j�n�g�S�>��VPz)�����n�駍T�#]q�~�@�
�d��9s�
�r�uϵ�]HNj+�eWsyw԰KejY7Q-`1FG�� ʬ�� ��5++�:ØkҚ�e��a�Ć�-*�&kT7��ٳ_�ʰi�	u>�F��Q��������c��U��n\<���v�Z�m������{Ab8!�YSNDD)B5�'f�������~vW��T{M��7�mܠ�&�U�O0�"��򘊮D@�L\�j�0T��t��D�lۜ�3�՗F����ӞW�sF#**ْ�o������LguP�1=��u�&����P�+S�8��Y�k/�O��R�TO���72�o����y����jz��,�8�����:�Ɩ]��Kp�_m$���p��-��b6�����Ц�BN�b��P�gT���:���ۚ�4uD:��qCd��Q�|&b��{�V0�q�M"��>�i�(�C��%��C\:�f;4��tD���*R̾�M{ܗ]�����MA�ǱV�g��a�] a�2�1�~ڜ~��t��|��n7��e��g����f8j�uښ'�l/���۰����rFN�
U�]7��H\m��u�;�=!��w�;����{`O��#��I��N����=�����b|{�=�Ɇ�.�޲��_	U�����b'f�ʒ��a�t�B��R���M6���(�qİL��͙���Ϣ���OX�bA�̄ݸX�[/�temX�*Q$<ܧ� (����ci���U4��YWm�W�T)nplڑ�j7}���|�����Y3&"���mf]�2��H�1�Zf ���$�R��Ǡ]ul2T��2:+U`�˽��ǽn�czp��"��AX><
uc��n��Ƹ$5`�>��Y��M���A,c��,�;X��3p�^4"��-�v�gL�/B�Q��\�+���o���u�qWzĒ�ϲoV�����{)Ҵ5_��X�ħ�R�˯R��CB�Ӌ�գ4>|��ξ��v�i��&]�E|JC�5w���s��=巐>��*��j�l>��5q��r ��;�`����T�tb�6}���!��Z P��0�T�]���L��tub|���)��a�y~�l�j]�ґ���?�u�0߭�T<ŝ6>��"���v	�o{���������Ϧ�����:0i�6U8�i����v����lyy��v���b�=�鵚p8!E)�G�ꈝ�b���.�[E���*K�	,�*�/�\���sG�:t͓�^��
��熉�@�w�PRf6a+g{�-�De*�9���+����h�R�[�<hvj%Ɲ��f�FE9c��XS
��tÈYz1Z��,���z�lѾv2K>���c�ڒ��o;|3
�����F=7Q�]�9�:]a�;���v	\sM��r�b�ܪ�0�J���[�o���*$̼z�ƌ'��<�|����޹�^߸�����;@H�M3���i\�=s�\37<��cܢ��-�}=�;_��P;LG^R�rF�1 �T)��r5�z�`|TIl\�M"�Ҏ�;L�É���[�N)�ԙS
G�K�&]j��'t�G3�7ZhЮ{������;���'��Y��@A0O����%Î����\;Rw� �!�O�nRn��X���᫡[�ٽ��:;wE7�aſ;���i�j����WW:��)~�{��!��Ú��A^�]B�:������t�'aÜ��S�UCb{!v�@Ac[���=8hV=Ul��wW�tp|�C´e>�z0-;�b��Mj�ڔ"���q=I��T���~R}�|%/�:QCl��\*�������a�L���ɍ������`U�R��Ŵ!�J�'�`��z����D�FؚQt ����lE����}8ʶlT�S�r1�ذ�C2
�D �9��~���K��ɜ�)<��p�ZT�Ԣ�?FP�ʜ�����*F��Wn;7�B�K�4�D�7)��r21�<��ή]אR�ބ��L(=�u�5,�[�,����q����;S�WKysU��CR.��5/�"�_�2˸�ܶ0�E����6����o}�`�\X�7���S��st�����5ȕ6!�ج��l�45������j�ߗ�_:}��A1y��}5=D���̵W��Q�2X�@�X��d� �N�&A-&j2-�'�j�-�Pj�XCB�"�{9�k�B!�{,隺�u��p�<Sթm^o�t%"���v�*�]���Ę�t���_6
�0�6�}33$�s�wF�YϮ=�OK]].�eCA�%)�9҂:������^xwI~�<��bevi�=�ԡH��9����6r2��
��_�rx��u�v
T��x7I��j]N�+h\d<���� ���k��':���#<��^�4�Ŧv�)������hD���p棄��i"Z:�ݑP�Y�Ӑ}f��r\!��y]�;	�Pٚ/ĪʍyY�GE�a�ܗQQlg3����R��\�U���P���I�
!�jAU���W�4iNj��z�N-��W�f.v-8��b�7��Tm϶
�h���͠y�y׵�v���j�➬�{����%�s�2��>"TWd���*�-͌�PEϔ@P��+��E���ib�z���B��ĕ��e����vHV��L�tp����%��J\���.4�m���^������!G?my��j���Js1��U���ԋR:^��pxB�Lq��2X.դ����!��)��jB� ��o<������X��ңJ�T�j�^�\T$���/�/n��j����
��.u�\�����_���u`ַ��|�a�Q��o|F_LL�]x�
��ZŽ�t�runΣD�Z��6�}}vw�rb����.���Z(����ͨ2�m���\�+y��u�7��ޘ8��&3�8��6�
����U4�Jm�[��MT3��b�M5�lc9D�N�ÿ����Kδ�Z2gb��p�I��pc#�	�A���H<��O��xSØkѪ�|���:�k�=ryo�;�����������g����
� \��EA���J�\�Df�X�	��R=JXR2	|w�L���L�EM��@J�O����]$�=��8=�*Ct3�6�y�j1ؤ��s�:�):q9Ȁ��L\�j�0T��"�S���\�K��#B ���g$wy��-@~����GARɨnv���������y��R|������	�����N����/i�YSy&�e�7&��!���!XT)��)�	f��{��?�bF��5�;ڰ��,T�o������|g��a���#B�
!�>q�kzt^f�s���[Im�Y],9�(�7[1���j�=K�d����m�Q`a�3%3e.��C����oR��]�cפV}J(]�酕�\��])��x)�/*b�Z첰g�⬳�����\^�N�h����V�N�	�%Ϭ.����e�}�𮺃�6�{\C�}ESk�����!��p]��{���)�+n���դ�H�Z����u��wR�H�2P9��&;x���j��V��9��S3V�]ҷ� q��k��S�\ҝa��]'��L��{Y��@S�t�ܛ�:ʊv�u�m:5�WQޥܝk�<}UU@$������b�5�{0��P������n��%�| ���\���Wi������-c���{z/��o�nK�)y@���)ns�6�TcqS���E�r�*[w^�(���,Uy�Rc"vƑ���`B��&aA/�@"��fJ�X���9!ۓש��u�N*�>~}ݸ[��<�N/���(p�X���uV���j��jlਉ�r��m7�'wR�a�֯%&����n�F$n(7^�я���*n�@�MR�ʊ�Kg�BYU��1v��m�L[�`=���7B�o�SɡR3[�EF�<�ɕ�y��o�G�V�sײ������_���!}=�M�a�@:�R���
��s���ȷ"*I��}���Y9��MDQ�'�%�Sq���&���f#Q@O/x�^��4o�Ɩ.��И����4z�N�͒1צ�t��Ks~�5$;ň�ʪ�	M�cވ����1��,�DR�܆ qe��k#Nb��c�VHB3$�b<�o�������{����'[�>l@�Qg>�VG
}�N������MR���y �O,Z]�{Wj��*5�CJ�dn��.`���d�C4]b�F��=`����rʭ�zM����:x�@gl������L*��#�	�_
��I���A=ZE��&|�塛��q��"��8��,�ط��i�*62�#e�6�s��r�.��h)��1�cC��a%,��FAɨ>j�̟>Fܨ���v��o-�������ݘ��NnC�Z#ok��7�B&�{Q��H��0�[Ծ�U��xm�a��s�/�+}�������c���z�CeZ�O���"��UA��`m�Xu���襩{�F�uM�K<�U����|��#\�W���C�b�R�Y�5�V�_�>Fp|��!ʲO.y����w۳�}t�p���]:8>C���(#�~'��}I��ݚv�SOO;/zڊ�25�E��\r)g��E6aK���*�d?��T�����nܫh 2c������o����]�^����j`�*W4�)=j�z����'�6�5��f���(���o��t�&罭����s�cT�9��b½��A�J�lx�_R�˂���n���qrf�lǽ�K �?P�Z-��X\jǽI]����P�<E*Q"�cU<����e�o�7�Iݺd����6���Gf]�PNޣ�_c�L��aU�1�Zf#B��e����(�2k<tB3t��=�V��#s�:+W�+k���*�rp:����-dGFq��:d��^�#���5q��k��ive�ٵHnH���æУÐ����_e�q�O]��~������Y�,�K��^�}1�ܸbY8!l�X��{���WC���g����A�����d�즆/�{N=�$(�-���E���V��w�ڬX#�9M��q�[�@�&da��5���ˊ�/�X66����i��`UVMl�k�Un�9�l�c$("Z12+�8���/>�Ϩ��~!^$����K,H�O�{:p�L��_NA���^�`�H��~n(��=6�;R|�lO9�yV6N;��g_S��~Qp��\�)̚�#��71~L���� <7�Pl4rd��9uړ��6x�֖��t�=�Q1�8#zr�b.��J!ߕ�CNh\d=��57�,1�0ۨ�p{�~~�p��u�t��f%Dh�j����� ��<X!D"�jD�wQ����$���=���]�x5c��}�>�c�~�g*m%w�b�S�
��0u�A���H�Ag6w�{�˷�(��̼������T��lxtw@8E ��̇��<O��e�{d�Y��;���C�I�W}���&�Y������I���l<a}��殘|¡�N������q���9~��f{�߬Y�OhLGE�N�Nsb٭u�ѕ���w6僂(�ު�m���*�bů1Զ�Ibn��]�XЈ��0��hw�WWk�0>]/�*��v�����Ӑh�Gq�c��������^M�b�K)�6v-�O	�u���>�����瞿s\�^��Q}`T���f�m����e{HVaܧ�P�� ��û���OR���b�2x��Nf�A�����{���>��J�g%@y�c'̩�)+�y߽��c>�\~g�v{Tw#��@
=�LϖO��~aRwϰX�{l�O\@QN�|��{x���!S��9��HV&�w&ߙ?'5`~��i�d����)�3 S�
0�ʫ1 �Ȟ���}~���y{?�J+�NO�D@�|����1�j�`xԬ�o�ӈu@🩞Xq�"�0����W��Y4�����y�����y3�Y�O3XB�r�i�d�5��{�����x5x��#^�w3�����)��  ��y��Tz�A�3�? ��ca̤i��y���
�C�M0�1S�c><�g�JśN:CI֓���0�=�]߿~�{�k{"��WtG<���D�G�@� 
�>v�P�auE��l:¡�;���gY*z_�T_X8����J��ɯd�)
����>C�H)��Rz�'R��~�bz�����s�#��{T����uo�Z��@�������P���~9܇��z�*Oݦ"��*b(zL�'P���n�s�l8¡���Pub����T�&�]'*M!S���']���Ñ?������\}��"�<d{����c+%zɼ�ϳ)�Y��H<���!��~T*�y�w`z�Vi�pE�Z��3�,*z�Pě�`kv�b,���������<W�G��~)��+�q�T "@w�0�v���6�~�L����@�}t°��';�<�Y*i�>�M�����4�Ag�$;̸B� �I��,�� �i��M!������gX�߳꿣+r���q���.��݁����4y�0�CV�r��Y�Y1w��0���1���c0����I��C��wv�+4�����PQ0*l�I6�������fq��Xz��_$���ʑ�1��}�Gt�!�R�j|��z�~Փ�O�0ߙ�B���o��l1!�|��i+8�+4~��Y:ʝE7��I�
���9�ugY1��U��ת_d>��y�eſ�.��,����|��R��:6;-�h,S,��U�4ՉNG�gb�՞`��������R�kAyř��s2]Z#M �x]'4s�z���$q5p5��گ���bɯd�f�]�<�:�Z\{���-}4]EM"����h˃D��1�f���1$D�3�r_A,0;�Ŭ�G;�ȳI���RPA��gK���V�H2����о�]�6-R��U#� TZGޑN�Jvf����ͽ�=q�0���� E�+O
(N]]��x����0k�qk��oJ�[G6@��5�e1Z����wk�5xyo�Rt�<�fa��6�Q�Պ��0uL���7�4��h���J{.�Tv��*lI��W#���d���DQ�1���R5-�fir8�uL�ُ#�بjڻ[�Y�<�2rB���V�"���S��xh�;�.#�4�(U��W$�p��r�U��кHg<�5�;��uh@�ʾHQ��]|�.�#����\u�H�:�/FH2dl�őpj1�ݙ�]wg@H�l� W������P�V3Q�άg(:��J,��V���KJ���4jT���5��X@�ս(���B5͋�W�_�fM=e5amn]^;�
�tB�&�+�n����h,f_e��o'Y��as�K:�a�s.8RJ�ʅ�a���4�y��h_Z��)x1�ۡ�e^eu*ŉ�F�q�5�իY�ש�{ϸ-j��q��Ӵ�{Y���0k�z�4��o$�F�"1��C$�b[�(�o7++�o`A��F�Xܣ!�j�����qcN(��m[�'��ܪbۭv��N�ܩofA���q.��@���Xbcg�[���h��l:�f���VA(t�L �+���s; �]`sOus���b$�x�WpN�u��ޖ�)�hǂ���Sʼq.�����KV�泲�p�,u���v:@���eI��X]�XڇP���20�x��8�,ʆO�������{���Btͺ�oE��\U�3���`�������;ܳ������?u�9�6G�5[�����:�A�W7�W��u�Ŏ
R<vL.+P�wXg[n�gX�u*$8�\[�9y��j�.�;s�����wEj1u1�0G����k:��� �����7�mgL���l���LU�����N�Iݖ(�,T�>�y�>B��u�IV�țSZ��L�gLLX�{89�3:����ڗ]�M,�(�.q۸�+���Q���f�4�wF��k(���6R�KN�TogS�$�YK��\����n���Qx>�m���I��g�[ [�Ļ(�G����Zs`z�T�*;�X�g�\W�U
G]@��op����mĒ�&*;܎u�{�VνYe�����3+۳�c9��8�4$0��y0���`�KE�Gh6xю��e���֟X�z!�E3Ao;g3���k�=�q��u\(P�*�   ���*�����Q*R�Աe�Dm�0��KcD�(�+mTd�Z(5(R�j"�D��X[J�KK[
�U��([kF(��TDE*J��-Y[mV�*֢+��Yh҈V[F
ʀ��*[e��V����iE�����c(ʊ�XVV6�m(�V[F�Tm�m�Z�1 �e�@X����R�J����[jեH�����+�*�l���[meF���Z�`�"*U�TTQb�U-iiB�"�U-�R�b�ԕ���E�
*�(��c+-J���iZ��*
5iX�cmPQe�"����ѶZ�+QTUQU��U���Th؊��+
6ҵcmR҉�Դ��A��!Z[K@�#Z֪�X�+l�Z"V6��1kQQ�elE��kD�-�,��6�Jضմ��ز�J�j��QE)P�[E[*��Z�Q`��D+�
+Z��m+jR��بPQb�ш�����j��V�2�Y� �cmm�DVQIUU*T׿~��#�O!�Il(���G�Ί=��^�q����E{�)�70��e�l7�6K܈�8Wj�$����� �CG�+֌�<#¦|c���M�(�a�{�i�'�l��ь�9�B���'�6���;�M�c>d�̛��z���7�'� ��p�d��8�T�-��egS���k�Z&�ةY�����+�"<����6ΰ�?!��֑݇��4���Hyhc��m���S�QI�� b����m�2~�䟷f�z³l���dq�����ҪAO�����������k�z���}y
�Af�@�/�B� ���w�<�Af�߿jO�
�N}Cl?3�z�No �d�]Ny��0�C���;�CL��&$��p�,6§�Y<7v��+���}�*��6a��+S}�(��
<2<& �)?j�g�v{f�PQz���a�I�>�y��|��HV���<C�P>�1�$�ĚJ�aOY1�w���
�~���0��~����_�	���]��~[ �1숁鏌�ԋ'�T�l�0�I�+&��M[:Ɍ>C�ۤ�A��֞�d��=�p:��@�8�;��N2z�i[�Ld{�����1���@�����V��Z�{�w�}�;�R
|�ܢ$�YR׺� }��B��Y>Ձ�YY�9�����Vq�'P��l�Ì1����=g�Y������w��8��=@�ћ<�ǽ�Z�����}sώ}��ft1��Y�C��
ì+1���� ����a�*�AN>��H��,���Xg)
�����H}i��a�mP��L�4Ì�=N|wi�%O��_������޳�]ڑSlǜ
�
��?x%^@�Y1	��iaS;a��ɴ�B��6gr�(�T��0R{�X�O;���PQ2o(�*M!���'���+<�S��'�s)<�[s��b~��|�Q��d���
|�������*A�=���ڰĞ~�7@�+4�<��mE�����)4��T6^dYm��c&�y�i=A���ֵ8�PS�.�?���F/���_�qP &<." ��s�~��|¿2x���4C�%z��r���S�<;��?+*�9��H~�*��27`cY]��
@QI���WIY�O�u���i��?�&��mS��w���f��Ŵ�@�0�:��x	����[ʛ��C�:W)X#��ނ�O8mk��S5J��b���n�p8^�y�|M-�ˣ2%x�f�O�X7�ou�-�O8����wr�x7r�+g�MfqP�3��T����}�o�������A�0��!�2~aR�7��i�8Ɍ�KTP���z����
βo;�����L��0�ΰ��I��U �����i�k�L�!\A}�i�����^���߽�������:)�����0�<a�b�Qj�Ĭ?3����6�ud��,�u�07��I�+7�&'��Qa�*w�o���VM�d�h�Va�p��O2�f���ǷY�u������o��}���>AAE�:{�Ci���<wvOY~�+�������r�CvLg䞸����H)��߹��*A���ɴ�����G(J�+72�E���~��&x}E�;�?-��j���DL`|>u��n��&0�}�B���5߲:�*���VO\N�Vy���OY=s���i������st��̕��rO7E ��̘$Ⲥ��Z�����]s�z��f����л�7�Vw�f�l5}�3�iE�{���Vz�Hm�,�A�����V!�M~�&�SL��s�ɤP�%|z�L�OP&=��pݷc�cã�cϔ(��E.Y�w��Ͻϱ�k� ��t���i*���bm�PY�>�@״�z���3��Cv����l?&!�+��f�
x����`��6�}��s%bͦ0�Mk�?n��+?n�w�������<3uf���ydS D��	�y� 0<����Ϩ�V���i$�Z��=��&�PQx�ՓI�
��~�A�,���@���l?0�)4���d
�RTT S���: [?oֆ���ܘ�0������QU~UG�U@c۰���i+=}��M (�jo�N"�����8�l�&&���I�a���svq��y�kB�d��z�w�'�|ɧ9ff�O�{͗���}��ߵs�{�~޻'�<a\a�?`��H,�yM5�yE ���	<VT>-#�!�Xqߙ������Y�1E=���t��a��z�$�u>9ܞ"ΰ�}�o���y�Z�n�����{��o{���%~O̘Ν�CH��J��9�����㿰w�!Xq�|��+'ߵ�s�y�6�$��72�'�<Af��T��!]o�8�H}hy=��m�Ɉ|�	3�o�����Z����7-�ӹ����q�R��L CEu�m)z���V��]�֩��-)���f��K�W�]��Y3�Wj�ɛ�;�&L�>�n6h�hom�]�&��en%g�2�Y��kqp��).W*�t�-]��@ַ��˚��>��H)�'�ݡ��1 �O�a�,�q�0�X{�O���?���i�a��z/(��Vy��Xk�(�<�j�~�Y7�i�=�"����Ƕ�n'F�{�����l���\�>�ǧd{�d�c�#�e'Y��R8��>��R
z��܇ό�����k�9n��%N{�U&�Nw
�'Ȥ�:�sy6��-��L��||���������￯!�!�,���=Bh̟݇���~I���$��~g�P�+	�>?Xq�l���O�J�5�`HT4x�" {�=���{��v�ݺ��ꟄC�LO�bC��֥g��kxCi�%�!�Y�s�7��W��L�!P�%t��VE'�Vu��0<�B�������Ou� �~�:�Sl�P|��ͱN;�Bsz�,��� 	�P����H?X��ۈ,�1!�L@��6���{��AM��{�Hz�C��+i8������>,6�Xi���;�$��xq��EU�;�*/�G�� 	�wH��(~I���f������4�N Wgy��|�z�����
�ܤ���n�Y�����N�R
o����*��2�4�ý�y����]�b�E�|sl�v ��xl� }��� � ��3h��?N�*d��l��a�& �� {l�%f���I����~�$��Ơ�����4»��d�'<�mw~yv�{��i�����y�ߏ�����i���Y�P(����� �C짿Y�CI[fs��Y�d�+mJ�a�;�4T1H;�s��a�Y���̆��+�u��IW�տ��t��s��9�rw�y � ���]^�Z��1�q��f�9�d���Sl�]�`bT
�M~�L��AݓÜɷ�,�1��۔��0�b{/�)*AM3G΄G� � ����]���#�}2�.>�\��ϲ�~��X�i��M�����<��I���~k!���I�~=��m��
�{C�C�;���;�m��T�>���M2l���O��M2nF� .<6<*�	빉���FF�q:7���g�Wݶ�
�TE�?�o�-��ogj�cf1$M딗�G"���ִ��ˍ�2��48!��L�*���吥��z�pp�f�j�)K7��2�mM;
�iף�8�إI}�:ں��7��	Ϧ�Lَ�c��/I���� U���|����%H����`�'�QHjg���'�0]!Sɪ~�m1���5H~���4�*J����2N��IY���P�'m�g�<���'S�wn��g���jߙ���۾F6�>�U?{� �M'�ԚI�*b>�E��B����q��֩75��%~d�(��LO�I�~fM$i�\�
��i�����Y�1���`q�c�<v��wT~��������� t��z{�w��z³��rO7Cԕ�|����*9�k�$�
�s�VO7��xk��g���XO��c8�Si+�AOP*~��η���3w��m<Oԕ��y��)�z�Y��N�����a����4!QH)��~�:�C�qa���k�%b�O���i�&!_���M�(�fs
�I��$��}�m��/�Y<��x(� {�}��G��m����+��>5�߽�v��J�O3E��S��f�m�ԫ�!Xi�2���甂�'����OR����ȧ̟�`�C�f�A������pya����`.�0y�@��'mN��y����>��ƠeM�����1��[f��i�T�<��C�gz��u����@�O���xg2s)
�������'����i�d����)��`@Dx�b����&�Mw�:�>���H?��~����B�>���p8�Vz�3�Ն"��Y�d6�C�b仰�E�a_����+���d�@QC���06�q|�&s+;�Q��1'6D�# ^�~I�+���3�My���&��%La�UU �?O9����yOw ��=La�9���0�y���
�C~�a�b�P�m��d�Y��4�����7��V9��o�:�SP~�z����`m�������!�6�����q�Cw�լ
βT|�AE����Ę����~���!Xm��h�!̤�ڤ��N�H��p�F�7ݘ~%�K�_�
Ǽb���;�i ��m3;��,6����w�l�RT����d�ʘ�3�T�B�c-�5�M��
���T��gY�����&��u������~��c�'`w�w-[��w}��V��=�зw�eZCL�K�����T�r����P�Wje��f
�[^ۗh��Ձ*u^��f�5�D�B��m0���;x��71�$��|�)�o�$w�,w�;gJ�)ڄS<pWh�quZR��p��?}UU���g���}Ͻ��6��B��O�a�Y6�j��++%xɬ��fS�
&���ͤXx����P<�0��Z��!����+R��XT��P���UN�ԅ��V�x��¥-�~\��o<��}�ą�?$�o0��P���i��I����3��g2�]0�+4���;@�VJ�f��dڪAN0��M'PY��.��,�c8�{�\��d��0��7V���_s�S�>B���T���m<C0/�Jŝ��8�iZM��f�d���q��T�h�=����m���}I��C��wv�+4������"Fǀ�{km��Sk�K��0�>CYa��fR�������9����j|��z�c%M�x�Ǚ�B�����l;�Hn�-�IY�IY���"��T�)��4��,{��dB�~w�9�����l�#ި�1
�����f���&�R���]& T���=��c'٬����'�6���;�f�1�2W�M���
AO�aI�eH>Y�~�wvT*O=��*,k�I���15? f|�Ǧ<�}�~������8�����b��#凬1i�`m!塌6w����L@QM��&��@�75�>Cl���o$�1��+4��y���8�`ET��0�S�;�����g�툈��N���~Ag@����!^����;�e �S߿jO�
�O��I�Y�i>Oӛ�H?Y+\�<a���C��C��LI��Xm�Oڟ{'Uu��ln�_r��`{�	��	�:}��u�C~}���`Vql�

/��=@�6��O�a�5�!X7̇5I������|��i*<�!���f��/��O=<������UU�y7/���&���Q�>�w <J�U%�b,��S���bO�����M[:Ɍ>C�n�q�Zo��M (�Y����IǇw�i�O\�!�1�|¿�4���p����}�{��w���y���߮�'���\C����H)ě�X"O�� ��\�ya�P��5d�V�ef�;����4��a��:�?��3�0�S׌1!�C�y�4�1�W�������ַsS��pݼ�#�R����z랒)k�X�2�l�#��"��Qq���!�Oz>��ӻdl����{/e��$ਉ�3h�A�����1u�;|��ѵ�NN���K,l�d�0p��[W]qo��r�f��!�Գb�yE��\�x{�������Ͼl���$������k�m��k9�����>aY�~���8ɝ������k$S�~q��V�B� �ϩ��֐_O)�&��
�4�SL9��0�$=���y�qeesS��*d����gɌ1!���a�4�5d�;��0�����ɴ�B��7��h�VaSG��I��`Vq<��AAE�ɼ��@�4���Ԟ����w����c`~�n��������;���O���B��O\IĽ��
z��Ϲ���T��{���a�<��n��ViXy���Y+*j~邓I:�Ce�E���&0�o^d��&G�}�1W?f7J�ɿ�8;��%@QN�̓��
��S�'�辶0�̞'5�!Y�%z��7E ��p�p6$����k���ҡ_7́���W����`{�䉝�.���v��1p&=��P<C�wwi�~a���!�C�����q�<-QC�J���RT+:ɬ���0��f�z�C�� ��<��i6�����GP6��Y��q}�[HK����{ٟ{֤xLT ����M�9h��4�|���T_�V%a�������AՓ̱f��1���N�Y�Y1>-"�aS��Xm%B��{���
Ì9��)s�O�}PN��W=ϑ#�eLǀ����$�

.!�߲N�T�&r���������`m��R~C�g��c?$�ě��H��Mo��� ����i��!�F�1+8��d�F��#�ϘJ>�@ F}�P����c����6���a�Y��c.����;>�y�64?SYx���g�X(C�=,^�0�l��{Q�G�Ռ�>�A_��Z��`�哵˿7k�g<����@�4���:�z�L0��5���{�B]{j�d�$H1
4�{^;�K�X�3#u�zcCa���A��m�@-m�1��Wv4�7�X����գ����4F�*pZ��^�~N��ҧ��1�9�N.7+cf�LY�tS��5�RQm�8[-�Yz����5e�l�:�éQ��Wh_�Ov�]��kb/����G9�*��:�,�	�E�ѕ(Fd�1oP����{󏋸�T�ڶ?4q�C�WM>qu��Q�͊Ѱ����0�'��#�TC�ަ ��*,*��v2`h������݂b�=&�������1s��|F�@�}s[Z�s��U
^�+|�� �R�+��]����ud�h��8����g�8�ÄDm�����鞋��ttEo�DLfbǙV��Fju�kşb�29��y��X��م.%����MGd��@��+�m�y�n����&���X��;~H���ǻ�����;�x��0}����xC�MrT�j��9�t�t�p{ `��=5p��et��r�]li�a^�w ��( ��s,Xz���L�U�Ķ=��cd?N�̪O�J�\"0{ǡ��`�R�=���H��.�dv�u�1����ؐ}��Zdt��S4mx�C�sy1���qo,��5�Ow���{Ƣ֗��'-�^R�=U�爉�U��<����&cC
�Γ���畊�#�(7ʹ6{�a#�Y�Ϋ:�:�q]񮍔U��wG�⧧B�Ǵ��OuL}��cU�s"c:�T�.=��
�����Ѥ5��K
B&,�/�Y6��)b���Ħ:��0*I�/�rǔ���=��<k�Z�!�z�� �M��ᡫ��+�����v�������<ֺF�/���"�B<D'6 �5�|��`�IU��Ջu~~wsW?,��U��֪�V���äB��)B����(-�a�C�&j2-�53�u�9t�r'W|�Ǧ�*��Ch�V:rx��!We;*ce��U#D|t�n�����l�pt�V5�S.�Aa}&��K�9x��"���+���y�F^��S�1���@����*UnȨ��2D79�! �=}W��]��*�Xg���x�([�9&��-GC}Cfh�;|�9Τ��ѰԤlW8Uc��u�Iҟd��2��;��ʶS��k��GV+��]��Ю���x'v/�ѽ5�2��>�u���dƔ�뛵�jFX>�O+a�/�k��>��t!��2Ő�#��*+�Vn4k�N�ZS��^!��}���! �o�o�6EK��ܬ'L�Gd�c�ht��z �����*����k���
�bX.��r�&����[
���N�����3}��*s.2���5Z�On�'KYlb�"NP]����� �B�r� �B��x�_l>5퇳�zc~Ք �i�<J�z/=���-����0#��h�'�jƻ�\Բ���f����-�lerS� �쇝�wMA1�v�Ǣ�t��x�����������8�|���P���ȕ�u"�Ss�ɴk���c޾j�vN���ܻ3�U��צ�;jH�fMC�U��đ��Z06B�L�ٱJ�
z�\��rW5��e�[�F���)��'*Br���ρ~�0<P��iUe�P��>��9
jn�V�\.Z°Q��N9
�3<������T8��� Ts�7 3�Jj5���%K��{��)tT0��x�؈u;�6sBg_�gb*o�Ј��k���^��_)�]�w�]���H�~��?-z���V�"��T�͵S*PX�A��g���5�K�w�'H�bb�mN�.�A�Ƭ��LuJ��g�
v���Y�Ea�[]��|���5RơS��� ��b�p�<*�^�c>u���aV�Nj�7�J/�;h�g����i�}�+�=��5^��|Ƒ��MA���z%ĳ��u]%���7�A�ۏEv�5uyZ�SvD81��W�..�g\����0}�!�k�I��k�-	Z���mM�m^�K���������h��iF��]I�f]����	�2�)�;�S�\��h��B�-���{�������ɳ����N�2^U�9�J9u�ذ*��lU-��u��>;�!�_���"#�[����9#o_Nθ�J{Yw�?j��uW�Sǧ���.>�@a��䌝��27���NMjG���g!8��R�n�ˣ<�5��Ep�4�;:��Z�y��WY���lע|�������L��%�������.�ظ������P������9���h:���7n2Vː�Wi׵��@���)����ݞ�~X���
W�W(�y���>�߰�4���kN���y�����k0�|t�{č���b�"��*ڲ��ע�z�V�Ҏ���<G|���=��i��O�mu���щ��nED�
K�"\@��CLB�H}!EH�Wu��a��y��ω�e�ܘ���\�]�T�$n([g�1��B#e,�ÜoU�m��^d��(e|R��;���|}�>]�:���6F�.�o�Fb/j��v�Qy�2�<�=/�0�J�>����2%n�e��V�7!ߡр/�UhX�Ou��}�u��rFotT�z�$L7WӰ0
�ɠu�F�$`�M��o�"X�9�h�Q8���k�35P�T�]Y�v���Ĩۮk^�w�#ge;/1�uE���]�ٍ��kki���ȷ�s �n��b�6/:������e����1��u'�C�JÙ�4+II#'/9�W��@�	wH(����H!w��A��|��Y��62b7*���[י��&��\�d6�"( ���mp�%͡��n�9� ��
���]� �@L8_�X�7FX�f�T���f�ה�Yu�F���q��YE��o6�3 (}c4wnL��[�Y��_ �����7pt�K��-h�ݷ|��3��EWa��w2���]}-Z��m�&S ��D��.��\h2��qvEޜժ����b��d[R��8�B���4Q<2����9��s{���:�2#ܪm)j*�SG��V�h��y}i^uL�Y�yiҾn���k��wib�L�y�_����I��12�JZgSs�B���ccz�.�
�Ӻ�b-:�6P�mr2�D��k��܈�Y�]�:/]g%YEjP�����j��,�GW<z*��j�^T�3-�!�.gp���%q@�;�o-W+v�]��3[����|S��)��X6�m�s:��Ḏ��%Jpj�e*�r��vK�tY����q��9Wu��5�|��q޳��%>�(��ף�W[���	�`�,p.��k�OO�b[j��%��]-w��[�Հ�����j�I�OT�b��[�.�&E��;L�W¹��{eT�,Ij*�`����Sfvt���k�P��.�-r�:�6%+[�y,+�K��.�GO 6��	��ЧL�@���2E:ݵY�s��y��)"��w�A���v�v[l����s�Y���G*7���8��lЗ��o��R�*6���Ϻ�R����uِ�Κ%�V��
Е��ހ��6-�-��F�������t�Ģ� 3�}�yu��{�ɬB=��%(R�!�xS6�ͪ�8������:�^d˫���J҅vJr: n[Ժ��(��x���V{�[��36f٪p�Β�2R�*gM��p�l�e-��ʗ/���$�{Ss��]9HW0�BM���:{PۣhR&Q�2�]
���;�wz��Z

$�:{i��չ/����Ns5�2�۪�[+I�m:�^Sj�ؑ2��ܻYK�O�����X�8��Ď�6��s=�3���z�Z��N�p01nֽ%wQ��F����1�:zu^��u��؊0.�p]�ԩ5-�����.�8&c}@ �s���s��ז�
�
WG�g�� ��L$=��Ycq3�sz�N۲^`]��U��f�=Zf)KE[��z�*�@��X�B�kɇ�k��`�[.�|����w7����M	0�s/B�F>LL�Z+!�t9Ԗ(���������v.��Ob#�G)�n�s{8]��if�����,�۹���ot|� |���W��+�T"���+�X�#ʌm�R��m�5��RR�(�[kZ�E�J�#e���*��mJ,1�e[T(����*TZ�(VڰD��T��������EEH���E���U�EjV%lDX�EVDeEE[h���Z��E��mE��
PQ��*"�* �*�ҬAb�x���P�Er�Am(,DA��U2�J��+Y�7,**��G
U��UD�UZ"�Q+QH�b"Ķ���bU�r��1TUhرF*���Z��[�D[jbQ�TQ�0��R ���*DD`�QC�U[lKaTE��
��TV�TZʊ����5+Z�U*
Z\�G)b
VPTe��faqQ�*
��1
�E��eU�kDQbe�rԨg�~���|{��o��}[1�������M�6��ɽ�ST�=���"�f��c���;�,��w\��t�ЗB�(X��=�=�㙘'�����@�1�@��~�Ë����:����^:B�Da-ʣ���Fmu_Q��n��C� �>�xEC^B�W��*��"��>�y��MXǘ�l50*#H�E����Q��d!�%J�f�u��4m�%�DTP�^<��v}��:�a���_N����G�3N�Ō<�v{�ǫ�&s~�[�T��ȫ��j�̗����-��9�xc][�&��Ei>�O=�O5��LF�1� �&��j��Ԏtљ]��V�+���n��|�]�̽�^G�C��fَ�>��_?.��x��b�E:\ً�sWT&O#�1�$�݋S��3�+�Lع|9��_:��l<�X�<~�#���T���x4fΩ���6��]�e��̧bzp>�\82*�����
ђ^�j�L�M�rq���7ݽ�N����F+S#��-ͺ�K�Ey�
\K�꾟
�X�{���,�<;����uOA�������z�̄��~�q��&n��{��F�|�����Yn���ը��s2�sEMN<�W�**�[��5���'����*�{W�=yq�H,hV����V'��S�%<�{;pͦ��z(�:��/l�ؠM�&Qtc�G�Hr�*S����BR�t�p��;"n;��9�� =�{�9xԫ��ED����D�C��
��5�<}"��{����Ӝ�Q�T��n���L�^�J�e��հq
��D�茛�Ȼ��\[V=�CXEX<�t��^ț�:˔�D��P�Ȩ�l��kO��p��,�9Wk�{ձv�.&�:�ه���o��-��7t'�������0{)��o!X/K�&4u�^Ğ,�˄����
銗�[����Z�Ȋh��0S�X���l���N§^=�V�}����]�P�mX;(�ѳ��ho0T_�3!@1�\L�C@��v�6��ӹ�1g�˹>����]�ָ=����+M�>i����;��O�$R)9����kz�G��WS�9 �q�B�uM��ф#L�1�&v��*�����m��J/
�R3דPX�92y���;CE9��"#c�6"=B�χP^҈xj3��\��*�R��%	��26/��XJ~�������[�bT�Ѱ�+�N�}Voܗ�� �Hd��^��	��űI��������ه\x:�E!F����)��b���zTZ��{0ŋ6��Y�{B��[u����&�AuNࢗ����3������n�cW:�u���&���+C+��Rw36R���u�g�W(�<  7g2��p�.�:B�}A)����dV��_�]A��	ŝ�j��QQL���݊l�w�����67j�ux&+$ݗ����ْ�C��e�/> J��[]ٖ����%>�˴�-�^��M2��u�5�zpV��/��Xw�,9��4:gn1�'2����rf��)9a�uu�-U���+���VS�c�A)�K�w����`���$F�v��`i�&�2�d��L=�ҹ��F�W�r��5�#c��o^��κ�b��ig^��/�c2��7J�ˉ�Bс��<6eH��*�l�:�t���MgF;:��<{��Uqp7=�k�w��r��'&(��lTC���l#�UhnR�j-Mm=a�5۱v��iq�=!��p�ݐ���3͞���1�ȑ
LF
@�>��CQ�X5��GqԻ�g�EE��8O[��d�(r���4��Tߋ��vnud'����	�o��e\C�3X�����i�S��\�ס��/ ���AKX���fe�� �V�Yq�ek��[��\�s�[�Mѹ��6���)V��]kl�m��P�␵�����K��K�f�I:�묀k�8پ�0�6��F��c�T������<MVumc��Mr�7�Ƞl��k6�6�2:�J����lw�{�����y��{�Dm#�����-����Dj�R3&���7(¾���̂�&�*}���Ϸ�w���� dk�5%�~�S�R�8*�e�­����u�;/᙮�h��J�0��B��Jj�LQEy�3F�=5�=�������0�9+I�Z�wdޖ��Z�]
��t�9�ϸ?�[�xTs���!��I�p�3��S�~�:��.��5��R��H��AM�"��\]�酌��K�\h�ւ���ѓߺy��b�o����*�y���ʮ�X�`0͗V�
��.���v�[p��1]��2��:5�{%WQ�0.\�A���=cij�2��MӞ��lh��#ӽ��M3�H��҉!�>�{�iu���1-�0���R.���L^f	�)(J��[��AN�[��t�Լ����ba]30*��R��ǠL�w���u���� ����hU����Q��0}+�q'��!ECLB�H����(��{aǤ�J?o��.=����������er���x�]��Ez��ц_:�٬��n��Į�X��B悗��Od� ���'�j9�`����;���nА�[�2���n��3�/���\���s��9��f�89=������Z����x  ���E:��FF�������8.{�ř�yS��������ע7�Ĩ�'����s�T".q���}5J<c�\�q������`S��Xl�mSɡ�L�˄����nbA�e�0��t,��^�{-��}�BĽ�^69N��Ғ̯oo&�U]ڔ�ӠחS���SN
��S�:P��t0K����L7�t+�+�7�Q�9�o:��l$xF�HW1D�9拋�@�8�Oe��o�/��\)c(�vb��,�悬��|&����x�$�lߜŚ��J�u�Ǯ�ć�ո�ʘ֩��؊=W�r_rd(c�Ϩ�(1Ir�n�8:��~���9�e��
��b2=P�Y�[9by��w��ߩ�y��c)27�Q�P�0���[)d�z25����D
w:C�1�>��X�\�D���[������V�P�X���7*��6ˏ��W��<��{��}Qwp2�}���UoR������xk6ʲ�nMz��#�TC�����F�GY���j��6߇�{2]����'�ޡ��-6�{�q�}�����S	U �^�F�Фכ"�4����umf�ڎ�+=�|��KΫZ,�Vpi�`�M.��s������@�'��v�.8�a�X{8J:�_ =�{޼̼;���`��j����h�{_%3Y{�C��ut'¶uP�Z�s��AJ�ܥ��3P���"ݧa���b���ݨ���(��9]�t���]�0]��:j)�j}�u00lqؽ��k�b*dst
�qȤ��0�Ŋq\!<���2WE4oc7�m����30�U�R���a�.{�C�X��=����n��<
OD�ܣQ��c^���>_{찲�Mo@�Ex]TC��"��N߇��og;5�W�T[�s��DaJ�l�zv�ˡVH@z�{���4ϖ�d�*v5WFǼX���l;sF�!�ev�\�e�iA��o͛ڡy*x�T�A�ڑң�L\����yg��..8\�N��G��Os�M�BLY�T�J\\�pCN��8�q�G�����7�#+��/.��wwF�AM��*�����<�q�3��{'6 ���q"4T��20�sP�����Q�����Q���=����ӹ�1�lo0T\�c&�(9�6o��/�C#�Q�6Yͤ� ��7ԋ\
�Ҋ���t���L���͡W}�d��s�_q7�[~V<(M��>QE{�A���ov ��=�l6nL�l�;J4X@wʱ�1(	�fU��r��ƒq�45V9�|���hdj��]��l�-�ld�&�p��ꪯ��+����mJW��e*��^ڬ�J��M���G��!vK �H�Ғ[�����Gl�T��˕���/т=T1�'�lX(\d]��ns��0��nb�.��lyKì�盒���8�F����vK��
������H_��5�.�]B���EfJR��+2t^��q����n9�TFF��3]�bK`�u��1*t����#b��
������v'c���ɭ�&cte�t��C>��Y�X/ޏۯl�*��8;��ܝ�+�޸�{��Tv22<����$0��h�z=�8��
��O6z&��JռoPȅ�$+�}��/YճM�5T���ʥ\�G�zv���T�bJ��]�r;$*���ͤZێ<�)(l�B.	B���*n ���Z6z	��P�pk��b%�;�����ۦ�Q�"�(b�|��.�#P���}fq���c���wpc������C�w�%��zzeܸW5�7J�:�v�Z06B�g��ҠH��tx�=���׉)�*��Z���w%fa��Hщ�u��v��v;q	;�"Od��]�u�@,����t�ݜ�i�r�,��Îp#���G2{��K9��'{N�m@3Uu^��A���/gwiQ��8uvi���;o��n>8ZΤG�<P������;�j��j{rmO޹����}��J�7hχx��r�n��`xU��v$M#.�%Ӽ����ntp�ݐ��i@;;�Hڜ�n�1�:#��%C���)Es�	2�Zs�sح��솔L ,�ب ^qQ|'����C3�6O0B�	�a�v"�r7Ux���|)����JM�q)Ww��J���C3P��.��>��T��epꈦ�Ø��DW����S��"u�;�cI��Ȼ�OE:,3��f�I��;({�VZc�.�~:���c����=Y� O<�{�H���D?u-��)n�#,�¥�o�,j#�lh;��ǽ����?j9
�
sP^h"b��F>cO���>g�c�3���D���=�ި������ibC�y���.�e�9"�Ḓ1���F��'jx;آs/h�J+�nK��V^�A�n��K�+>�t�ac"��]xZ��eESۼelM�iQ��E^͊�Z��c����=�a�����lעU�ؘ�N��:")�9�n'����\k��ަ��u��M�B����+�n� �sޝu��K�eݚ�_�-ST���yo���'�6K�K=�bPQ���Hqt��vA���{� �� ��cj��汪�܍I��G�Ż�{�����������S��P>��P��������\Bꑫ�ZNC�lm!�T������Z}�rZ����|�u\k��^L�FVՁʔI��}�r�hW:]��E�<�\Gx��r�gt��wc}y-M���We���k�<���v��GD��:¿S3 %#��
�.���Hޘr`�ȷ��7p�.�%μ��S�;�]KR*%5%�È�����ɭK*�p9e6��č�
zgZ<��t�C�F�9S��]�T�č������-z��==lc[,z��tŔ*�\>c��wF�}+V��Ys��<�u���Eƭ�F,�I*͝�r=4�
�3�}�fw��UC��g�8>���l3������!n��Psds��[8*iK��(A������2N��]�8�&q�R��1Jz��)v�G��f"���Hv@~એ�x;]O�+\�����8��$v���]׳V��TX�Œ�oD�p2ަ"�'Q���b,@��T��v[�1�c�l�:��=��.Z���o�i�*�s�L7Xw3�h�R���F0��kLhC�i���H��I�3��5:�]1�)�4;�u�H��q��.wYӊ���{��ۉ\x���ᡝ=����7��o��+h呶D�G+��� Ö�G�y�Q�����+>����.X��fN�|�٣mX�>g�����{bu���#0�L쌃���f���ݎ�u��a69Vð�f/ѐrj0�C#��UgO'��2��a:L�,;p�TP-��!���w��Q7 �tV�����<z��]wwj5���4L�X�w�����?���l�v��Ue|ܡ�)D9_$���1��3��j{�@aT_�U����z�>����Җ�>�鴪��;l+�����K�Vw[�55>y�.���i���F)�$���N����j�tp|v6WZ̐�j��Z�R9�b.�:�6OO^׋8�L�n�s�:�IEz5�
\c�1M����sO2M��o]\�
h^f(�=]�㰰]_��>d%7��{���&n��8<�:�C�sK�ڍ+��'"G�>_n��;+��2Q\.��5�<ƹh]li�a	8!!V_\�q��$hfHae( �ʜ�?J��!Q�!��~u'�UpvՏx����� ��?o��B�����^rDV��vҜl��('S�Q{S��q��.�]M�IjbL�<��)φ"�8�zmUMa��aY.����ֺy��F^�x��A��z{

�����]o���nY�E�r��u&��+/�So���i���D�j�ϔ\mfk�F8a�2Ҽ�:�����n�E�!���u+�i�N��+�R�ݻ+<����r��E|-^ё<ʺQ������pM.���D��%	[����[�_*�ۣJ��W\���h�۷��؃2����*��E���}ʻvp��u��� A�/��ʅ!���tN��+M=Q�����#P��| ]�/v� ��=������餎v��U:.s��L5�l��^#2WG��u����N��is�.b�YŜ���;�o�d�Je&�z(�z%���
Ӭ���hܤ�:��]"9Ij�Dq��ʇʒ����J}e(;�yre��e-g�`7��w�m]1�,5��c੫�z�m�LA��:T�Q�{����N��9T@!���3���\0f��[H[���7��Vb}{���Q4�c��fa��Xwн
�X����M�5��"˱·bb�0Ѩv�L+4����n��vW'z0���e-z�J��+bѳDķ�6N��Ӳ�W;�a�\�`�V�9|�����Pm��;���x����o7/9@�;�;�ɨeLIW.��tɃ�^���7\p��}�b&����HR���!z7J�b\ŁN^]!����z^�C摴�ͫh���Z�]!�[�\�rVc���U+��-�v$dϔh]ևP��]=}R��LT�V�MZ�L���vhvʭx��^��[��SCv��s	�#]b��z.�),�$�uJïm���9Rsd2��Q���Ӯ��rX�bN� T0R��N���s������:a:Y��oCc\7.������5�sF�Zk��P�j��j�D�#���ce����\����:6�9�K�/T�L�Sx.y�x/�E�iڗ���= �K�6�S�IA�O�
{�mL]Y|�V�uXE�8ؗ1��$�{	�/J��xl�hlň���n�o"51��r�zIs�;�խ��s8;�!̩)p�*L�mXy�u:��"9���+��q�O<���cWcF]�*����u2���ֳ�]J>���Yo+C����b���Ӈj���ۂI�K��!�u�</�$А��n\�O�(�_>�3��@�EA0�Y;��h�7[!�w�0AC����"&�����������n<Y�2����H�ch=B�\T"U��K۵�ْ2EnE��D⵮�7�p�`8������|y�ΖR��,��� p�ę����#���1i�F�U����/9�4�ɜԵ�:�ia�M��F�o2��8r��7��#��	hb��7d�W�&;�����~���^���*J*,PDZ�D�Uj
�E�T��m��cRҖ�j#����֙h������V""�$��S��,��6���ł6�
�%�-�b+Eh��Ŋ(�m�*�[cQ����B��%[�0�Vk*T
���J�h�e�1�mm
1aF*�R��m�4�UjUQ[Q�PA"�ETb���%�DE�V
**��-Z#�QL�EA��q
"�EPZ�R�b��m�-�(+h6���VT
�*(,-[�*"-���6�X����cX��eb���(+@X���Q�DQ�+1J�,A�*DQ*�B�T
�"�X�E� �ŀ�c�"��(�icPU�T�h��(*��R�(�%�UJ�X�Yj�kQQ�Ɣ�#-��B���Q�+�ZB�n�vvR��n�+���Ds/�u��		�G��C��כ�2��k]��8��n���BY��$�]r�SE~��Y�d�Ǻ������s��B��G�*Q ����GJ�������\�.���g�X1Zp��p�9�w+�nT5�sМ��d���eLp��P�Q
W����l�o�s�7n���d�ǚЭ�MaQ�!E�L����b=���M�V5n$A��ĥ�m����'N�z��VK��|kK�rوW��9���Qr����\D���[�㏆򶻷j&Ba�F���FE����Ĝ���G�ʬO�Z C� v����35�5sq�"�B=��Y\��>�
�,u���#�lS�LA�s���mBt���fL��#ٵ��p��-Grz�Q��j��L�4"�@h�'0������]B�<V��;���Ʌ;�D=�Q»�i�2�ګ	^���N���1*h��j#p�Y�3�]��Yw�O% ���gT9;!D%A�����خ�����ذ�Y�Z:Z���0k��U*V�VeƐ����'�ζ���Sٲh��Zo��KE��ME�H<B�wC�W��4��Y�����Խ�&��y���@�X�d6z	J����t7�xw�mع�ċ7KO�&ל���O!ŀ�.���w��{�2�*�J�dbT���T7x\��!�G;��s�������)�a&�ud�KG1����me�����?x{�3[���ն/}�z*���peD�N2������ONO�h|X���]�
�l%|h�\u���E�{4:d��XDRU]"�*Ȃ-��hP�W���uWG�i�ܭǲ�;�g-AS1{��S
��ԅ�h��������FN��qx�7�R	����>	,ku�ȣ�a-�r� 7*�E�F�puN$��^�`l�~�x0s���m�`���x��n��cc Rd�29s��NT�'&(QQ$7L,}�����K�!Z����������!J��6���!ԍ��l� ݝ�jXxx�<����㽜�[���
�)����|�&��� G:F��'�!\&pA�(+����X.�*�Ω�܌X*� =����N�u�����ʝ��ϭz�Z�^� -��vK�B�yx�2y><Q��\΢?`�H�w�IK��S��� ����x.5�gQ~Խ�d8�L��RA�����q@l���MT��L�ؚ�ӂ��e��<*�3A�o�Ot&f�na�T�{_�n��M�YH�ml����<��݋�1��u8��2�L����1MK�`�үy��9 �iv�9ř;��cr��o���;�R,�m.4�#k�i�F<��n�;�){�QÝ�쮶#��7���}�}`�G��sʢpɁ0�~!B��!XT)��yN�^����#g�҇���Fd]�Zyu*�-��{y�EE�/�����P� |��o�y��Ƚ�D;p��ş��پ�z�'�w	[��Z��8l|�(���Ô��ᓰ���)�ڮ�t��I�}��z�����yv�����>���Q�v�0�ʘ�)�t�����銫�U�LٯD15�s�xG~ދ �ۥ'N�I�c����Ob�]x�
ָ=�){\Bꑨ:-����u]K�\k��(�,�
���|�*���EBl���L�FVՎT�O��!W�@F�^�WU�l�٥���:��j��p�h��'e�ڑ�j6�9���*UeJbf:'��f`B��&����%¼a����I��{P����2\����U�;ቜ�nED���]C��3��������`g����GE��[<�.{�Ń#vH�N�k�ʜJ�PL��!��Փx��jaSz�L�!��Ր8Dl��Y� �S�<�[T���p�"%�s��)`�;rtϧ���x#�m���r���y8�{�oUrkfm��R�e��;彔j�h�TݡJfK�z�u�h��x�C�ru���6������������DD]m|�iF+v���lj"W���g��ô���`V���kNr�Zg>��y�+��TtX��ܭɡ31���!��7Bʨx0ͯx�X]h`��tM�yy�Rv�Y�
f�ٰi�6
� T��v
�ɣ�����W�MV�.�+���a�K�L><b*��BćsZ�h4\]�uk�Y��
��И���N�F<�ud�j~�7�F�lP���o"�����sb>0)���
"��N��:�r���:�di��ŌV}G(!���aA��^o�2h�E�m�\�l�c�(��/u���.��B�9�mI�6-g�;�N27v;Q�VI��*�vT�ü��5��a�[t��E�;�=�b�NmEY��2OZ�_���xi�M�F���ٔv����õn��=Z��9��?��A�)[Υ�<�ub�5ʅ���˨m_�Ӊ6�ph۽�����J�-u1 �EB��#Ch�J��D�6.F�$f��K�0G��T�[�v{Q�TK~�^%~�+.U]�d[�'a��=�L���ډ/P��LvP@yI5B����� �Z����;�V����iN}J����(^��6b���+H����9��eƷj��2R��W���Se����K\�u*�`�I��.i���|��f.4̊��H/�����w
'Wv�K�: )o<�c��Y\/�꯫�n�îO{�(}��6%3��=�z0-;���Db�2:�"�ۮ9�������ol�k�{�ɢ�W�w����= Y��#�Ga`V�|�Jo���c�&%�W��6zk�w>D�lձ�\L����[Cҹ�%Q\.��+�xU���
�S��sa��]��e��}2��6�@�7Nd��(8�GH"]tFM�>u �\-�}R@����/%��}�=��� �3�I�.��ĪUYB�i�BB����A�ܯ"fo^`������&��Z�2bl��qlק�7..Y8"��;Sh8�zUD(<�oa�i���U���m�A{Ϻ�2]�"��Tx�F�P@Ɋ��q�$W#�Bsbj+"+}��*�|d"��x�6IՕ-_�2���=���}����t��uAW�\�%38Hu�%�lV���`dD��	����hd�bz鿬*��s��s�E��ӐcǦ!N�1��u�D�7<�ff`-�C�ӊ��8G��[S�3[q� �9�	���bc�rd��~��Ϳx��04ی��eŌ��� �l;N@�u��L�N�1
�Q�Vٛ�{���.�X��|��r�Xxa�I�<��ru��)s�����a`������^Z�|u<��59��K��y��A��A�H���}��+z��{����Of�x��;jc��>�'
���~�
�֠4R�1�X󜊩�4���TW��z���Q� 1���fˈ|���Ddlc�3D�bH��������?�Ѱ�Lx%Ƽ�Γ�g��Ͼ\�0���ME�Uv�ZH!V;���Wg�_������9��
W�ӆA�}ȌLz�Y�cWL�0|.}�Pt;}!5�@���}#��U]{#���Cu���$ӫ�b�o���G��+��h�>��TKD�P��]��'ƴ>.��WR�z8��7�Sݑo��tk`(
�&��L�6�T%�Uт/ԫ"�z-	���dKΎzk�]1r�H�L�܏!<{���=�X�mH�)�/PE8<!*��0F�Ź�
�z�T������X�NH�c��CY�}ը��\�w5H�*s.'�ׂ�P6B�g��U(OVUrd�g�n��\]t�T�; � ��ys���r�����QQ'̓�L�B�#*��������8��HG�x�ICV�Ԭ�� ����hi�+���nΈ�"�B�cJ뜆1,��As������@iQ�{�Ծ2Bk�Q��b��^U)Fm�y(Ĝ6���*�ml�w���\i�款w�n���ل�һl�ؠ�X��\'ul�Wh vt�M�������5u-o��qݑD��E�f�_R��r�h]i��O��U؆�7��F��+����)U��������&��Ucf!�=#`T�"bn���@k��Y���m��n���>T G�g����]$�=�󲸻��zV�����S�f�*�e��[|����:B���t��ʞR�=��lR�Nh1��붭�.����!���U��6�:��b+ d5U/��W��7C2@���Q�s֍j�pƏd�Yp�nɆT12C��9
�T)�Ay���-E>cH�g��v������"鋞ygs8�ZC�H���Щ9m@������.�gC�{"�xn'M(�Z�lv�ǻGb֗Y�3��F�u�\���B�h9H9��AH�#�������^�XHi7)�{��F?}7�].���.��"K���`v��el�6�K���R�Rf*�;�k��9�1U�9�SP-�t�r4��M�}��X���FK�=��
��1�܏\qryu��S< t0;���v�c%l���h��o.����~�ܱ���U�e�����Ўjl�;��i�R���I����,ӂ�8�7�J�>r2�oq�łʗ7 �}K$Z����hn�^����ц�~��e��K:�${�~� ̬��S��f�2����v{IK:Ӝ�b-B}n�;�!����\/���1yDڭ���NU�r9��O��l���6�j�~�\�nT<3�/=3C�
陀��;�zu�v_5�u:%9�z�R�vםhY���}����jK���yEl��]�C�G�V0:UkuV�ׂT5`�6y��wG�֊lN����+䏩y8��N��z��57�A��}@b�8Dl��:2����x:�7��F�WP���p�S8�fu8�wz_#���H�nU��R3C`��Ȩ�ǀ#&�EE�Ss�g^3�T}���8�{s�<q�r�&���p���3��ʧ���W�!Y�Imn�����O�ݜEN>�|C�7�X	}��C�5�@�U8..���&�ژ5��;�v��t��x��E�Q�[�0�����b(>�1�x�(R��"�멪��yc������4��ꛌ��cb�;>���%��fN�[�4Y8�8'8\����w-���Z}�������9,*���>��J�����,ux���g.�n:x}�<�!-}r���r��f�qWce�H�̵*�p�09������¶���I�������&p���s���g&������貉س��C� �^n�}���d-�8&�.M���ʓ�5�\1��}���ԏ!�y���/�}&����̕�ە �=kv��/���Kk�d��@mV����I�])��?T�7�J8]�v1�0��K�u��1��2��:U���k�<v^R�o��u�5�.��,K��bEPy;�=R��Q&l\�!#7>2�����Mݦ:{����jF\�4��T9��P�޲-�v9��*ddN�ݨ��
 �),V�Z2c����Ir�hsf��eň�PG���==ck�V�G7@���E"�1�h���A)��'N��n	g%���12�=]�V�2\�2����$�.�{3%b��U�㏻��|DђZ�E���w���szJ��]�hS����ީ���$��oSg���[��(��C27֩@��ә��Q��F�-�OΤ���8�;o`�3���ɸ*]�pzFK�@6oj��%��T�A�`�|���Qb�.r{}��@��;��k�M����Y�J����]�@��,צ6����gjb��J��b�b�w�)�{�u	G��dV@��M�6�`�iu4 7ԑ8�%-��g�PlꙝO$�Q判��4#zko�X��}�w)ʻ�jm�t��Sf�"h�}W����Պ>�[p@��[�]���\!8�=�����jYew`���J�gl7�gW~�T-�9�Q+�|FM_"(����Ѵ�-��@�,G��؂�VDT����ځ"�<ʿw_n���)Uö��_Z�vY��f !]B�1J4�O���޻f����u�>���f�M2835���"�U�vT�-��@�o������2jz{��B���V����m�R8G��@�K��h��'?�>��`6�I�g���O�[
j���8�#��PqD<7�Pm��{��GS.�� ح��h�k�*א���ƅ���q��A�P���;A������и���6f�xv$�Gs�5B�*�4�:y�ڔWE�
�sCL�1��!D"H*������W>>���V��&��FI��Q1S��ދ;\�� ʃ\�`��t��@��|o�z������s~��o O>�q0|�#�Wd�,�h��.w*�8~��ON
и��la����?;�p���+���]��R;$%:g[�*��+>�]�Xy�F�q��*g��=	���K�Q�Հ(��2e�w����UYK�K���T�7�[�j�[�u�qYΌ8�����t*$������o`T����r�n*؎�w3x��WmI�إ|�L�L�b��*�kF&.Tӗ[¨t����`?;څf�	P�΄p8�h��+q�w�����A�U�O����h �ŻO�n��¬�0Նl����LK�2����s#B����6���QM�q�2�C+D�R]zW�P2E�jݫ[.<DS�e)��Ԭ�9��iԴ]�z2�M��;a8��,V.�d���n����
-�����������We
`tQoN*.�ӕ{��[�#�����W����,�]x�Բ]��Q�Ȋ��Hέǀ�z���D�5��`^��E�4*�o
;�V1C;��d;X�h��
c���F3��8V�ɡ�ohl-d�g��'�B�A}�ho8���eu��b�[�i^]�g�]����p�xv݄�F�|Z�/�<Th�j�oZGZc���J�Z�E.�t�ey���v��F`w6�m��M��oq'����|��-�D6��}/y����k��I��覟�_'���B���s���f��XI�����9�wSv3sn���-[Q��]�@qk"�i�3��3K.Z�k7���F�(��ud_������j��VPLwt7��Y��n�A�d�IէK�b�����>���S�����;��ƅ{.��%��6)��
����U��
�aU�m� )�#�!P.�0��ͬ	�	�a1XF��N��˥���!�E_d�r�9�w5�a$^�d��EXm��0VY��Q�,ų�X����]��Ѕ�n�X�ae^��uv��ڹdK��aW\t�Sê$�1��)�NS��eq�2�ԁ�n��
)�s�ÛD�V�̼x�7y�öE0&�<�^�p�]��!��%��ՙ\��hd������褞=����x+{e<|ڍ.΢!�K�'a��ਗ਼�k����{-*���r����GL��7X�H�G�y�T��j^ hI��n��A^e%ZYx�J�����eX�Q�͚�N���d�ͣ�Y*��MY]}f�N��J�#ȗV�ą�s�O��+u��d�مW`=��w`-��7�f�.RQ�K���,��=[������>5�2*}�� ��1��cӄ�V���;�ܘw%�p�J��$o�E�����4��\�୤�|�������r�Q�
]�K��<��\MV.���7>Z�.uc���N&�N�s�E\�:�۩�4��'p<Ϻ���㭬w�+6覆u�E\��j��+���st̐j��P��U�}J���D�E�I�b�`Ǣ_!�i�[�
e*�yW�I�*_7���@ʵ]��V�{��s���.+�hc�IL�ǭ-!�;��s���1%{!� i�!"��������?@*��E�J�6�QPb��J �A�UDEDAV
�X1U����*1*%��X�)���C��
�[�,1�[aj+k-m1j[`�"�H�������*+Ub�R,B�DPDU����Zȱ���V�Pb��EVcS-�R�-��b*�����������Qk���(,�8	��QEU\�&Q�j�e�����%�QTq�1*��A��8��X�*�2�\�ģ�X�E"��̩�01E1*�1q��Im��X�ЩXV��Tr�X��QIYUEf1IPm.Z��+2��b��(,APYZ*��Q2�33 �1���E����.%2�T�"�����(��R"��q�2#E(
E�EF(�J6�V(�H�"�DD9J�B�T��2+? >� I P R!��ʸ���{]�㳵���<7����>ɪ��P��"j)�}��cN�\�����eJ��8��p[{���啗�:.t�s-I�Ð�n~��(v%����g�V:�R,)�z�#���
�*#f�H��̅�F�'�ۋZ�����:&����Ud�o�C��#֑�U��8�6�F�Q\�N���d纻����U;`ˮ�O�R�F�S�s�; �'!�s���r��	Ɋ��
#+�*�.�cd��b��ߪ��/�����9�U�E��i�#gvC�d��X"�B�2춶c��T��"..&!�HܠP�v$��EA���s;��AN�-�O[����m�W8��jN9~���T�t""���	Vk� ,W�~VW��nL��\_{�w;�^�F�)u(��5���j��E���O����!a�7�6)I� EД9�}�weJ{���a�T({&���}Q
����<� ���I��R�S��Kt�n���4Ź�{u����&��Y�ޓac$8`���%"\�h41G�C�S3���G,Wv8���\��zY��������7A�F2�0��+����l�E�lӞ)x�����	�������L3LA��.'$��>�87��k!4�d{ =�%�<�5��e�'>7w֯�h���S�<��7or)�`7�G0�B@�K����yR���D��m��n�çRN�ұ�kx�rPރs��ٳ�-K(��>#X�R|�^�h�YSޕ�Ѫ����Vpuq��^�l�0'~i�-Owt$��^��;>�[ң�+��>��LZKB���d��Ҝ��3��ВsCjcb�_������Y���)�g�{�B�ƔɱO\BѨ9´<�X<�gl��On�96�ֈ5Ϟ���uK%����ھT�Hx��*��#ׂ*�	�s1�&[B76vu���ш`nP;P�9��jA�F6�"�A�t����ڗ��g��ꚧ�Z嵦��ـ9���ˤtJs^�u�~9��yօY��ذ13�6�b[�3�r4T�B��0���3�+�suV+�R��,��*�\Y��$r�e�d��B�[O��vW=Iյ,-f⅄Ϣ(c�8>�"6QgD&�G���#����V޼��cEI��X���u(;�z��s#Z��B,�f ���"�g#&�^Y�������0Iᖭe�m�N�?�~���������;��:�S��`��\/�SN
�E�[������o�V�����S7q�a+�b|�ŕ)�NvR�#N�b��'-��[}yc�6�ԵH	w��#�T�lu��`t���q���,MC����:�R�eb
�I����������]��-�]��-��.�Sx�]ȳ^؃jwDf�R�Rt)�@쑂T6#�	�DM�!�CQ K�q%�/a���QZ+�m��W���'f�iV��ҕ�t���ߴMB��o"��Ͱj�.�]C[���XJOq-ίw��^�e��z�縭�%Ɲ��f����.X��f�u������Y"����;z�hҟ�eYz�W���� f0�c��ǲ*r��X�N�W�m���F艹�y��a�A׹T'�QVa�L�K��t��'�=�B4�7�{P����YU�=�bޠ�p�ܹ�B��Κ3`FF��!^�qB� �g��0��Rv�
��]�'uesQ'��`�yJ!�z���R�UA��6�jy>*&,�$f��Q�/E� �����&��;���xVC��i}��P��ȷ~NÂ�F)S#"w��b��%�ٵ��0b�-���|�4����Eڮ֘����Z>�z%azvV/�8yH�l�r���nM(���֪e�W�����8��;Jd:��U*=]}���{uJ�s!)�F=6r~ҥ��+BT�K���/K��@��/���̲ �q��8��ڌ��Q�f�H˳Fw���i
�^�x�^Y���ٮ��}D-�7�1`ʃ;9,�]�Ժ�� ��yq�)}�;�؇۔i�flvxf�{vW!r�X��D뺂Jrc�vn����q��w}bc��������_.�[Cҹ��(_���y����pH��R�a�xzt��V^�{�r-J�"4�̟c�(΢4�Q��,ϓ�������1�~rSK��������r6
�(l:�v㱳{T/%��J�HlPz�*2�÷~B�GR��n%���`_W��*Jr"�љN-���Tt7.!�X�3�1Rzg��Ѹ��jϷ<W �Xz�b"��T��.<tmd�Kv�k��	͈�u�E]�vY���Gpջ0���R����.��ʛ:S���� +�
���9X/��3����x�Y��řT<* U{�&���xe��侑��G#�&�������;<3����u�yCT�.<��*ܮ�l�6�P5$G�S@�I�f��.2(]��:�tL��E=�}J��ch�v鹋L�PqE���1x�ɒ؊GTG@�U�V�c5�_�<��<�,a�����*=Aͥ�+��`'Ddl`}Cfh�;|�9�%-Y�o�<�)�3˴�W@�hu��{�s���9��#����������p:q�U0 �"(��y�;Tb�HQ���(�w�}�n�ኙ]��`���4�b�z2asPߔ��u')㈊=�:��緃S��j���;:6��WT.�l軺q*�Zv�#b�«��,;�<^�9�q�c���n��vin�k�r	̙�3��o7��O��؇ô5cs�ճ��P�����$ ��h�z=�2a�-�z�dg7�]��\��w�ؘ`<��B�'���TKD�xg���_ֽ9l������n���TQ�p�	�r����2�`Xr;$%:gCa��BU]"�IX�G��<a=~�:�)x=���
�B�׹��]r��q�b���ԋR:��NV%Dl�X�J�ʕc���ED1�w��2mHqd�Cx�P�L��J�sPm#t��q'k�B9+:o�ݫ�j��5R�l�uǆ�ҠB���%ι�\����G#�}cY9S~���YY�����\�����f vRǅ��s���ݯ	��>��0ףU��������~�M�K�V��N͘j��@h`�@�.��|(��U����\p��]�̎ra�<�uV"�v;�+�d=��U���;S`B"(J�H���UDdW����T� I0��*~��se���h���g;�Ω!�l���L���e��U�J�D��1.�_�z����p��+{�J��T<f�pi��3�.�f��0,��=]-١�����{"b��m����q�+y�ձg'��K��deC��5�Sh��;�'�r{�� %[Ϋ����5S*KL��`�z"vK�3��!�ۙ�cv.-́����V�X��2��B������ ����O��V�x�r��<��ыs���{�
�2ˇ`a�yI�P�VHp��9
�
sPC��CGѤ%�F�Xْsxa��u����1bɫ��۵�f��L�����0��~pWy�z��=7�;��)4�Cf���u�ş�ݴ�'�l-*{ҸKj���x�\r���ЊGH �%��3��K�b���W�)kP=॓Ɛ��C`6.�w07�S	�9��.�{�OOʶ��؊��N:͜�:Jj��i.�ƸV���O�1t2��9���(�%л]�բ�u��W^T)W��{���C�J�y���ڱʔI��}�}���ާמ�9cx�Ƣ�VVD[>��
[�ٵ ���m�.d�(�8מ#�$h:9ͤ�����s1?.��X�{���T�`��3%�;5�Ѽ*���d����7^��~jI$�skptg*�#�]�u��hZ�'�,�e^�C���"�g�������>�z��G/{Gq�L�㱪�+�N�h��.�+,�+K�Tx���ҐX�K{T���m� qS��O�Tu�%nbJ���AD��[҄�H��Lۼ��83{q��`�p:���S�����b��B��4�+�$2Y"8�(�e��r�t�Fk0ޠҝ~�R�^��0︼�	]�M�cfⅆϢ+����Sk(U��U{��~>�ݑhZ��Ǎr���ܧs��<�u�F�.�iI�{��]a7�n��8!۳ہd>5ۣ�Y����||>в����V��I��рL੿N$J�<�_N��Π$�,�QfV�
���1�=�Q@�>�*
��L7�7���!��j$	拉��Tb�o��W��ܴd��Pލ�4z�A��9��t���[�D� } =�b*u;�\^�����C����E۫�h�U/e�.�ƇM̍9���3^��E���aFqS]Z'�mD���R噗^a�1�F���I�"�N��Cb�v0�£c)�7f�Ӣhg��M��yҕuŅ,U��*q�Bò��*���պ�7K��tϪu�����r�_*vmj���DvN)�~ޠD�;���:���4f�##	U[ԾǞ�1��7\C��g�A�H����)��*���y�`:ήg^�@���w�;��J���I4롏h�W�\5�q'�jfR� e�{��o��]ʈ89Cc�2�]�O��I㦛l�Ѣ�<�u�:��RX{εr��|����Vqc:�B�eū��o��%lg�5�i���QHަ �*,*�����oz+�ؽ�{C����ƽYs�)�ՉTƗ;��.���h���A25�Bm��;=�����r�D�X�n\V��I�c�r3���"pG~��۝K}��.���ݼcBYڒ5zXr�U��6 K���U��/�W�I�3U�º�X�*�,>�㏮Kl˿)�1y'�\0�V+ǵN�ݹcn�V�j���X���9�v�dq�'rm# �⽏ʀ��F_:�;��T�4�K�N'���FJ�wJ����96�H��&�/*�Qj�T��u��QP/����H�2��G6�C�;�"Fffp�F:k�T�c���=�Cv�`��\ߎ6F��}�[�y�Q���W�O�)Ia5ȕc2��o8�CY�Me�yBۚ �U����T�Ѵ�\F���b���T �X;n�H�7;��]�+;=������>Cl1ڬ����<�)Q7c7�����n���YaK��wv�E|28��r���D�*ט0�m�g���/�t�*�j]���^]�jGˀ�@S��}F����$�ݫ���{�0�hYj,My���"l��^U��l��+�О����M>�3{���Y\��0tt�S����QSA����٧[���4n�������I���C1l�c�b���c+��6��F5�C\t�q���gW���u�;��N��7Ha��A�/z]���٢lFO�Aɭ�SK����3����Z.v�Z�;��|�iPb�\�vװ6�K��uڕNd��p���2��OJ�\�bq����=�n;1'���B�N�g���<���o��]�ʇb�L�"x�s�Ѯ�H��&!��fV&����;���@:X��{%XS��]�*����b����®A��|k�Ƌ�5cK㫸�S� c�V<��
z(b�'Q=7��ev��ݴ��LOX+����d�k���������n\���<�"�T��dvF'�A���כԅ��ka��Mue�=�n�¡"���PTo��V�`{�lx�o7��c�rd�\F5۸���s&�fH���df�2Z�*Hۉ��/`㹎虘���9C�l�Ou���*um�2{�:_�����BJZ=�q��?Moz�:���rN���ʑ���re�h��y���ֽ���׫0�`��2� �e��a�т�����A�,$p[W#E'�(*�n;�s�h�gF�~�9p"�,Vv�<N7���YU�/�>����$Rp!x"k-e-�؊¢lc�KUE�vΝȡ3��"Z�A�O�g�5��&Op��r�k�K���X{%��QM��HGcI1���D>]Bb���Cܷj�>��\��D���W�.��n��C)��؊�t^h٬g5�dC❙K
4���C���J�m�۷yt�hW��Ϲc�O,=y��[9�rKn��?>��+.)�z_5�]�S��-�C11hGt�_U	q��1�;c_�������͎ �8�~��OJ�\��y	cn&G(�oڦ�t��֛���p�X�7�Cu}Wa�ξ���=t���
A�lG�b�r+���4�
{�Q�ֹ��Lbc�M��.���J��V�l5�'b���zF���fk���k%�v%Z��udz���Ժ���NmoIY3d<�	��qZb�Ŗ��\s��W*R��ju�y�����m��NS�E6sZ{W^q�죨�t֢1
�[ޖ�y�E�k��`i���gs*:#�	��1�P���v��I�E{ђ��B�s6�����.�K���f�{Á�E��2�gp�ī�l�c&����q��Knq�v�)��ls�HWv*s�\�� ���hZ��00����:�ю���uj��.�v�S�3OkCV�u�u$-e�9�� ���j_*|4�V��n6��ű�)�^��[��ݹc�	���Ym��I���휡�����h��[rRu/ng!�� �]j��2r,Q����P�٣Z���ޘGg;(��L�mDr�o��t�(5��z0d�w�%��%�����0I�pfb�[-�^Nn��"v{.������2m��d�%�䷻Ѩ�����*����W0��� ��[ī}��vh�4&��
����6�e��u�h�I�Y�F8e���w*أ��Ȓ��q�-2*��fvlP>r�dk���G��G0��qbyX�FHrk�����v��}�`�V�
TGz^1��H<O��]\� ۋz��D�t�H���R���g9v��t����#�噘vW���ru�8����Yt���>n����v��yJo-&Vhʽ�ޛxe��wfչ`I�0�9\ԔI�&����Z�ǵ|t(�nL�OA~���Gxj֮=3ਜ਼��������`�uK�gr�v"��
T��z��"�es'��'iV�B�_,�"p]
�m��jld�O��r�_v^խX�N�:�W�RbN	M�b����i �X��9�"�%�`�p+�k7ԭ�i垕��,#*胛
�HA�w���A�fڙ�0,�;9��Ȳ��^�rZ�O�r���N.�=�}8>���{a����1#H�T^s|Z��zJ������{`ZÂ�t�<����q8e,��*kE���/�o~�z�u�6ŝ��L-J���vJ��c�)tu�V&*�n��d��b���9�M����r���<��3iY�Cj˳�9F�7)��A�s$5cv%C/r���)e`k^��ݦn�n��3a;J%ݲz���3�K�۵������ne�2��=�Xg��d�nu���:Wk3cz���Kn���)�0�]�m���yx)�����Z"��2pF���t�=\d�+hq�ݺ	���x���uh<#}.ތ�;�b��s��<��N�µY�q�ږ��+2b���Ƅ��o�ޗg���fې��uZ�"gz`�,�(���2�d�[�0c|1��qN�ʪ��CDT��UW�E�#"�ƢŊ��-b��"�H+eG�Q+TR�f!X���8ٌ��i*+Y�IE�L)+"1TE1
.&dP��DˎKe��Qd�Uckl-��
�AbfAm���B�E��"�AA��VDU �-Ɗ$QV�X����E�QJъ-j"�-j�Z�R�ЬTbAAUUEDE�j���+�U��$U��TJ�S,+XQf�����QE#iA2�F1�X�ej	i
�EX"("*"�+*h�B�KAE�ZX�ն�P��R�����KR�J�E��թDX�A\)Y*��W� (P�Њ��u �� ��}f�u�s����[����D��@oo:����J�̴���L��uKI����;z��%6CQ:��9�o�*�I��+H�Ǜ�s]*������TvK���p�e>���a����U����B�Av*m6ՇK���]���b�6�̪֮��#CG1ո�b�=�PMޕ�Q�N;�V�9y,��ۺ��˛��3Gj�|��1�;����W>�cd���Ͻ$��݌��}������jH����P��P�4"p��VLv�,�W���Pz��3��-_^v%X{��Y�6��Cn+��j�7��$C��fg�7�{��\&�`�c���uP�o��-<�i(�t@�w�OW^MR��_U�˛z��"�\p*g��O6�C�4�I��T��w�Qb���r�n�l�f[2A�4FH��xL�y�a;APm��iS�u�Wp��vgBb�n�D�ړe��Q�l��{���ĞQJ'S���Ui��79�e;q�ܔ������l5�neik)�䕠+<sՙ���r���@�Gq�����n�Z��hv�x��dł5��c�H�
=��h�A�N-�vM��,(+T�i��:�}�v#����ʵ�LNK��(uE��k��3ܹB� �z�SC^�'w
�����tFRᅱUx�Q6��qqn�~ǹJ���Z��>X�e�as���aM�gfu����W`�J��ʮ�悜�u�?j�WS��&�j��5A�Y�����IQ{��O{�{���f��pc5B6�k�����y�^�/u�^��ͺ�f�g:���WY�N�����:�a�J1�7�<�aΘ�}D[wU{���.TD��r5Ո�\���A>�M��v'3�2�H�S�yH�j��y��B��D��V��g�Q}E�253���_7������|g�:תGn���U�=��f\pJz�"7Ǻ������ܙ}�L�Z8s�۠�.�~O�Hm�v�W�y'�W>�~;���U
ޕ�Tf���o��b�5[���@r��L΋H�!�1�U�j{/��5�3%��❦�حj�.ܬ�r��v��U���2ѡ�v��W5���0��Qꫭ6@���J����	ځ�������#���3�8/��pL��wQ˟nd�1
�
#
���o�su��T0�\�.��G��l��aL,���
�\�Q�Ր��a��v�u�V����6��E%�����	]U��=yB�d� ��$B׃%h�eߎ�zy�p���
L[�'���s�Z����Y�+�îPwP�:��6tm#���*r�a�#k��	���v�,'�k�A������Zʼ�m�*�2�=���9K��]����qpa0Z�'�Mz"k-������G��_(39f�=������rT��{'&4�����hlםnڪ�v�X�yM��]��+b�0�r�Le60X�]N�y��l5qA�s'�[0]�cN����t���g'��t��
�3�m�9S��׳[8c�YV�9f�=J���itT��'�YH�����A��#�Z�N#�qk,�Ȍ�WwkV��kz+���qW�_��u#s�
���ǵ�^T̉*��/�k|PU�ܫ��]K���%KjP��6+M�f�2�[��T���o�a��JɌ���it��R�P˶w�J��;��} ��nMF�g�c�'Y����m��Q�̠�cj��l�
�b��}#	�b�:�E�KW4%���)I7��f�k3_T��qo����7�A�\@T;���ősדs�n��N�WT/0��O�6պX��{%(�lv�C�S��f�o:�
3*�U��xt�'��z�럞zO�I��[����j:4b�N����ͷH��Sƞ59�kF=b��Ȳ�Y8ݮ��Ց��6���}��6�t�Әg{R31���}��ᐤv����+��C�4���{�ܳy7��5�/�L���ߝ�j�;B��Vo3)��"/^`8�mO*�v����X��V9����I��As���P�8��q��dޭ�{�U�t-�W	bAu�pu�v�O �'`���H��P�5���X9Y\뙇��]�袱No!F_Y�>�(��cy�}	�j��L�%y�9�1�"�F�.�<���uy^���Q�l���&�cQf�kf�Ѯ�"�}�[>�Ǒ\�~]0���{�~��6�B����V���X:��%/(dj&4W(sz����[�n�}6

'֏-m5���)ɪѼ��
 �뫛z�&�m"��l6$g�L2��[i1�Ĺ2�����^a��^�:���\���F��R^��k�aUv��7G�HV��v%��7�w:E�[�qשd��[��#hk��;��fݼ7Ha�4+
����Lvj�]�3t����y5R3~�7���X÷b��/���ꋪ֎�6duJ�ckM���k���i�qy5бs�Ƶ*�l�]����P��*�u�ڟ�OrQ6���=�eXV��w�5ү�z���Q�A:��:��:�9w�L�!���.]��1�Qi�����N�V���c[^Ҭwd���m������WQA7cJ����E���"�;�M�|�UN�{=�s>��D���F�:�j�ݨ�\�71Z3��7U���6��Q�9�.Ը�c�CB�ڃ�������@��@��c���*7;����=g$�H�>m�?<��/E�H��e�=��bEѷX$�nB������Tٽu�I��}��2k�t魖���tf�3YS�}��,K�=餽�{'Jb�Zu�4��5I��q0e�ᕼ�Er��lpށV�Z4���3�pݮ�sV�1�S8�:�wIh��n�t�^G&f*��/y.2y��ۻK��
�o�8���(��Ym��ě��}g4V|�_K��GW�`t��m�$`<}K�)C�\����9�yi�����>��
'zNS���	l����N��Z0%yyګ�}�/9#1�X��&��15���*ۚJ���B�C{7�M���j�İ��K��hk>��ǂ��I��y�?�u8N���ь��c����%����>i��h�y���8n��ݡv���:��B�zo��Ԫ.���z�]N�ÓE���χ&s5ӫjz�L_C	]~��<���ȺC��jQ�yk�Ưf�6+܁k����za�FO�����-�5a��7:y�5�@E"�n6�Vi��j��:SZ��wp�`�B�8}+����h1β�	��7��YdM'4x����'�h�˔g9��kr�B#��u;Ӯ�x��y��p�I(�A��k;L���p��ѷ���]��l��]ۨ��Ը�t���u��l�d龣�aG9�gWT���;�da�y�F*3��t��o��[x.��)��u�`"'iD˴�t������5�u�W�.2��_�8#�������lˉ;��fl:G�h�t�RouG0��~s�*��UuNʡ��l�*��?V�2q��KFħT�%��_���į���w>�>m�w�=�^I��U�*���6'�]֕�ݮ����6V�u�;��;q;�i6⽏ʶ&ȜG�����cU>�s�0��H��Í��*��/Z��ʤf����XF�PR�@]z���j�$�V!�>����e�ڎm�n}�����j�.ޭ"��F�'�W�A�X2���W":�C�,#R�[�ε�xe�'�a��TӁBP�DMe��^U�4�]Kj됙ݭ�����Uu�p�+GH�aLY�j,M4"���D�rlT% ݮJs;`�ۺU��N�B�0;OQ)3�`�R;)�I�j&sτU46s�(����(���Q*�^)���*��&*�5f�S"i>wl�Q��ۛ��>D��Ѻ���
�|ą8����k��� ��j�6H.�R���	)��l�;�Y
�(V��{�_nʚ��1�o*�ľ͑=��^_K�gv�l�`�P��%�''�Ϊ���,eu:y�(�W&�3ѱ�d��C��K��[��٭��6+*�,>�C1�'����O�V�}�騂���kU9sY�7�ǮӮ�7YH���ZF �٨%��w��W=�[�-l�^F+�G'[ޅ`�����]u#s�P|{��x���쨽��+=�,���~�<X��z���.*�b�V3���h�r"�2n�.�Z�E��T����1��Ζ7r�OCav�n4S�m'�3��J��9�(�E�i�-�58�1���u��ZO�Y�'���k���;u6deأ��-\8݅�Z�;3*�j�H?#,[����/Շ��};��%���UQڶ��̤�8т]	���Y���Q�Դ��"�2%(�7�V��6�"a����EWu
QK:��ulS�\��<Ɛ����]j�⤕:�kh_.�҈gT;=!+Ղn9e��ʶ:w+��l�{�(5@^>}�\+�؆��RS�VA��i���r��l�%�$�[�F귻Hur�q�]�L�i�4�[��M�!��9��\��u?���l�"���R�U���J��>����i��ڞ*j6�K��ŅZFL�ک���4�N�z�(u?U���^�C�r����E8s�G��1tKhE���	��5&��0k�Z���n7�|��'�꼻S���2�#n�>�籉���Ğ��y.�s����.WQ�Ln��c��'wz�(]�"� e!@al�Q�/dG?^�zn�J\�WԚ嗗L�l�3�F��4n��V�ۼ�C1�l�o2ª
�����Ό榈����K7 }{4|��b��jWu������ٱJ�M�i� �v]��7������7^سp.��[��X�)��%�ʥp�����1.Q\���^�=����Tk)�)Ǜ�l�z)�\�4�JY�g�Ss�ꪍ.w��=E�؂�5Sm_�,n:�1��U1���<�I�^mͨ�����:��%��[�[ x�<�uԊ\���#{��[�`��b�޷G�Л��4�477���<��NI6�Aǅ�k�}V݂
5݃�[��.BwZ��fc�:�M
Y̱�1U�+z����U�#�w)VO<�)9����]��X��(&�J�5 bq�%t���=9Wc/���n���k4�>���)�C��>U�!]�vuR�8f0qV�W�D#�x��we����G��Т׹��Ћ�eY1ڐ���l'�s��KOk�7��j��,k��rO��dq��-{Q�ђR�����o���Z��݃�n�U�D�}a���y �J6��{T;�6�]nօ�E@�X�s�Fr�K��v�O6Ò1��d骖�+�~�{ßj��΀��T3N�g�d��
��n	o�^�����LE:�R�7�"U��"_��C^���YY�m�*�SgD�v�g4W<p.�l�<^��0�`n�Ɔ5&��Mg�;�����[.���b�Q�7L�E��V{�U��;�]$�M>c���a�~�Y���9�l
8d���2� l���ʋ�Z�&�D�*��l(K<�dZ5d�i@���j4��0�O
���r�lU�+Hrf����ـ��V�ӷu6���8��� � �v��N��D�l8����}������\;pkw�$W=�C����3éX���� ��7���TP\}͈�2�i��I���>��Vo%
wkk�1��D�e̛�F�6�ĈO����V���Csm'W��2�����%�?=��m$�Y�ܕç�oj�R	\�\��y훕��9���'EN� ��=<.8�;X�.{M�X��G�t�v�v�Gx���&`����G�я/�}5�1�\����h���tEYy,)�.�SD!Wp-[�$����]I�gB�8H�����)�23rpy���䵑׃���p���v���V�_�r���R��Y�Cz�7e��j�ԭ�۽J�)v��]�%ݒ�:\�E����@G)m��ͩ����e=j�\Cu���:�<�}�M�D򲱗ʮ���w���P!3H�,��܀���+z���:[����qT��Σݳ;F��Y�������#桼RΌ�`�L�.��hNqkCoi0z�`���b���8vCGig��V�-X����ᓻU��A��`�ќ��J�����L[�;(���T	�ܱՀl�9]�W�t<Gof��p����r�Ց[LW�ӡz�XG���sy�M#��Ÿ�	�9�YɁ�J�o�1�'I�VX�6���;�n��7�ޭ���7f��X
���h����+���K?gKb6���y~��4�hyT�o�7��][��xx-�aw=<	iS�δ�u�%���:����ԍ�w�\+��]A-k��:Ֆb͢*#�,W���ڙ/�ܝAEl<�ާw.1fՍ���ѦF�af�`	�����`�֣ʳ��ܢ�WV*C���̺�V}��������Յ�_u�+��/g)V�Sf�mm���>|2ٕji�u�
�/<�x�78��ù�ձ��q�'և��}t��@�ل�	Z#&Z:)k{`��U��l�0�.�V�"RQ�ݩl��&����ұ�]5|�J.K�J���,E����Wc�Wj_Y�E�:�V1)1�3/��*�L�u{w]K�v>umI+b}c�᪱.�����
vݮ�*�M�䬫]_L޶�.��j�F��[ҥ��lদ;���Ȏ��ݟ%Y�����f�����7��69�\x��1s|+�p���uf��tF^���}�
Y����e���] 7�RI�nnpׇkl%�{n͌cN��:�	�<��A�Kh�lu����ٌF�����;��W�mzO����1ʖ*sq�ܐf��k�+TY���vƫ8l����sn�3�4\n�L5�;����e��0�n�Zҷy�k��:�w}���-KQ�=�.���`��[B�j+ZT�-�ZьQ��CJUjU-�VTm�m�[Z��QaR�E��ar���D�(�B��VVc��)@YPT�e��lm��1���*��V�Z�\�jҢ�JV��%V+m"�iAb�K��kJUb���Ҷ�c�PQm%b�����R���*�*�KZ���Qj"�H�E��T��e��[B���F.8�**�m���PQTTU1[PQ����+l�Y�k**��T[j1��jU)Kj�F�2�����ZcKK��ne�mX�Z�J�d��"���j�b9j�cZ��Z���G.dQ�Y[+kKKjʰ�KJ+R�m��)PT��֑Gh)����IPS)U�Z�X�m����ҥ�X��T�QjV�S��5*e��2���J"EZ%J�2��\�����|�3�۴���ڽ���	A�vtL�P�p8[׽n���f]��^�ی+gb��J;7�8�w3%����o|���&�j��QS�F�fww�W�u(;��:����]!�����F�-y����6&x��zsv�%���)��E[�p��r�VR"�h�b5���@S�4��1l�p�T�,���T�O1�⼬^�x%��s֏�v�P|q�~����I�{�f_�L؏#��=Y-��ǃ�{g�ͨ�at(�Z��E��7��*�2y҆�6#~Kw_e���#� 6�۞�W�=a3.8"v%X��7<����*p���ė��/�����w��㏬����)�^I�u��}�����zն��Nv�����`�kwG,��̔�Sn(���+:�7�lg-�K�����>UQ���n��*�\�V��g'F!�P�Kct�R�*��f�k�@�D�#q�,[Df2�kƖ��B�6l�8k�ո�ڇ$����vv����\�sBL;�ӭ���{����d��uE���WY�4<A��b�)t5S=隯ow��3u9�][9X�e]-h�(G�y�����ҭ�ǋ���v��5�K�.��O�I"�'���S�m.��'����n;�g��΍�Uc��-��=�U"%%r��dBvV"�ӊ���V1_b��r��|�Ȧg�����TZ��GH'���0��Ŗ���B��f&��1ҕ�WZ����1kOJ�-�����Z��|"����	������p��s/�pU�z���B���ؗK�y�5�|��j�Pra-M���9l�5W���3��ݻ�E�7Ha�41��������q�]q͜�|�ۼ��׳D�@l�0�MueW����rXxv��̴p�)�5�.��Y������+^N*��,y7�������{;�Y8�<���~�C6��=�t����<�GaqT;�V:���_(�L��g�Z\Q�ll��q�����V�cq�;�]�PN���r옶r���g28o�aF����잾��2��lV.X��#�Y�Cz"����)۴�S�ݜnE�,X�:]&F�����±��Om	��V�[yjBG�{�N�{#�7>�w��@e��޳p��g�U䂶�w�N���i��t��xM�f�n�<9-���[C�-��^K����*�y>Tr�]���\0ʱ^����۵�Z�*t��U��n�ȍz�$j�U�Ot(��~�5%��*�9����Ľ�yX�\����9���y5[�宮J�J��^�}�۩�H��.��{���*�䫍oXV&c3�'��l�6�H4��W��e����訩t-[�]�ټ⹫�F�8>��<ф�x&S�e�ڄ��L^�f��Sʊ۷C��p�r���7�C�a��(�[�F6j��	;k�w�p�~5�rn�SE�G)���pr��	qX+=E��'��>�n���y��~"'wU�]�ۣ�(-��:���ǳ��C�o�m�w��۔���6h����H�4f[�V���]<�&�f�x!�|"x��t$�3�rʊn���RWXBҷ����Y���>gt����`ws�t0ig�)q!ԣ3��W7l�>=33Œ���W!�l��_QS�V-Du��4�Fn]������>�=r���H
��Q5ב�F%�T0+�Z0j���ir
n���Ո����{���{������F(�X&��������x܍��D�����?8�5�B��w�:��^p <f�1�kJ����i������4�^�*K|�n6�U��FY��nk\�ٶ\9��UX׽�zu�=j�Py��s�OBm�㳫���My��*ܚ���0�f�
��r!W`�"���A<���/E��S�A5�V�6Qz�QJ3u�Sp��ئ�#�q�vB"�u�ꅍ�������.��Z��,�C�>��Hm�v�M�u44'</�{�4��U��7���^�|Ms��X;��ݮY؝���2n+��uq�s�5����j��bj����v�u�V��l��H4�4K��vL�>����S�d� Ϫ�1ɜH��9<۸ua����&v��F��m���'*���h��*�}r�4;"Y�x.xT�����;Fa6׽2^R�6��&�B�j�5ef�2V«�^mq�wE�NU�p@T�
�.�<��b/,�tXS�z唳1��ʸ��L*�ţKհ������Ԍ�Oެ��a�Gq��������#�Ѧ-iV4\-�ș�'��n�e����,My��CY�����Bۚ:f���m�;������p���)P��S�\)�,�&�B*�CY'-�k*�!��>0�d�N�T{9k�Ui��XR��vS�cd��ߥX3��{>Β�>���G��VK[�ci
S>�t�ׇ&�0�-�7��rw-���Tه�������2��W��f����m�����ɭ�������t־Ԯ������u�����-
���8�j0����cu�,����ēϚ�
�q��z�_�z���A� �=�iu"f�A%&��l��,
{g�6%��|'�s�2p�_N�i���Ok\���.-P4��̌e�]�mc�=���z)������[g�}ዞ-��k�G�Don4۝�S��Q� �#��Jǫ7�히	������tz�2��΋�:6�j��ͩ��V�ݜkzh�$��}=����[�WL@t���M$�{[�e�~�_ n�2u���ٝ�83�yVcΰ�مu�*<��!��;^W�VU~���߸��:��8�ϛy.��V/!sd`�a�J��t�����ȝ�Gy�/U�mn���؝������bEA��7/z!�љ��[���+�MP��۳�VyN>�I:p��:��q��#����C�� ���� j H3����-��L	ލu���Շj�;R�����5Ղ����.q���.A�5�q�4�u;���0z���47Ƕ�yD'`�Ոi��(k15���L���#�'(�gln4(�g��8��Uw�DBb�QbZ�Ƿ�P�bOV-�:&5�.q�ڜ�Ei�W�.���Ur�C�=�h$�59E�Pƙ��9S���io]�Ly�����yv��g%
[�[�=�	��Ċ��ԅ��r���S귮:\����o�F41|�v�y����P��Sg�������p׾�� T6�˒�;4�=���ւm;��\fX*uNUc��U��6���0����)t����擥�3�ւ2Ղ,��V��v���[޵'j��rrWQ�5K{l�u���
�r��I�J�]'VH���3�yP�z�/^U+���*�^�-��Ŵ��u5
H��	�*��7��{Ј+�8���u����]�V.b����p�sQ%��8���ɳdځr3���K�齕w�X���v�8�DL�2���쭕��\u|�j��c��H��6��nuqs+-.���u�0#���f����<9�_j��i����U"���ѩ򪜒��� �8���U�����-��T�L�qTm˻U�z�;[*�C��֌�-��K�UP�մ����2�u�+s�!�8�N�CX秗��g$�U�ߝ^�D�ׄ�={y�w�T�L<�6�\d�9������7�8��A��W�㎭�QO�65���X=�r�L���h�	�>i���N�驡PK�l�dve��́�b����!���`����j�����܋���Q�d�N�#~ʹ�'z�?>fJ:�+9��W�U�P0�[�X\�;�Ҏ����Q�܏[�G*G!"�&#�L:n9�Q��<�XU��=Cew][$�:tSԆ2���')ە��G	�o0�'u۶��r_@2���M��t�,o�7&�SN�\�����{s�+џjo�v�n��!���������"wq�ʻ� ���!C�[Ws�.;r[椔��*�7�f����> c����y[�v�V���`�o�c�U�1
���>�t�����\W�9KA���2/	���Nm�#�5�<��/1�.��'Y�"�������;��V�I׽6�83V����l;r�1�WN�h9G�Ӝf�QIF;��g��]tc*/�ls�3NG7v����\V�չ����]>nooܒ�؅��#hF�'("�De�.J��~r�v�5��rЫ�OX�_��\\��#
s��ܥRo���M[���Ӱ���*��{����=A^{U�}ck�-����9-]�������!S���LT+DQ"��#E
���K8
�}1�Y����3e�^�)剡�KZ�'�f�&���aW\�t�s��PӁ��[�]zÀ�}�UI."I�2���pw�O�b�[p��CG �S�n-�2v�.�Z�<ǜ�H��n����^��\3N��,�^��+&��b�B���Z߽gv��;��H�!���.����Q�e�U>�s�0�i��f6wt���BU�n�}i��y��9f�=��+�[�d��mn@܁F��&��q����Ӄ�FP̪;�]«�ir����RP!a���^x�H�h��@�-�ɂ"qH���j�]V��0_v�0Ղ�X�8�CY5��ՙBۚ:d>11��Mr�2�NraVWh����($ş5&�Њ���#�$_r����U�Q��9/�����Q)װ�=��&,繅��a�\�g$2��z&>��T���~'n�h��CdX�K����O�t6'Ce��+�Zr�v�d�F�N��NNʁ�,�[B�oB6��,�~���F6n���h������9��:ξĝ2v"�*��s�B���w�V^��)V��ufm�H*�4:��7;���ݑ������tď%����nv^Qf,o=9�Ba�;�@�� .%�g�.$͝-��)�X����ޡmIH�]^nn�x&�bI���[�r�}��_�Q{O׹U~�aŝ�;E�V��x�G)���
�E�z�ڭ|'�Y�ɯ�y���w�h��¨zj4%�.v�A��s�1�WL��ԓ��m�*u�%�pS�=a�>dv�����d��"�_D^L�0�d����I`��#)��(�K�V��d�
z)��B��;[��˜ȥ��ä���OX���}φ��Wv?�mim����gdV��=Ek�%,�}�;#El�%أ�e�q���#��;��,,�B�ușٻ�x��Z��%�ș"78�m��.�f2�p���m����斑ɶ�F�P�x����D=��<c&���E;%�'ʮ�\�i�Xi܍��+�8�v(\�S۳��B��:�]RSU��{j9�!��p+҆�����%*��]��r�ur�j�m��!1���$T�-��pPW7�*4
�jc�� %��37�m�ޤ�j���&��Z�{�;�j
=+[r.�ˠ�h��h���(vDe�庫��b�V2V+����/�]��˝���"|2��g���3:�d�d�(
�Йʊ+ɴwQ��",�G7�oj�u�d���&��MNF�1؎�-���۵��;�	�8/�+�9D����`6��U'[���q�i��0�B!|�vnL��teF�Us�f��Nl[������\�t|�ٽ`�b݋� �Q4ZP���X����8V�;�%$3!g�e�o���[���s)��]�7w���[�y9�P�V�d+k�oe�q�N+����Kso���V󤹳o9Im����P���k���R�,6�7OaW�)i˭δE��e����ˎN�y\�����5f�!��8�U>X�j[z:�]��Z�[�Y��"ޘ��J	Iϋ�,H�x�"wf:X�o]e���Zi1L�;��WIugn��RG^��WN���u�F�&>��E�f�\�;-4��U��zm���|Ǖ�`�Gi�*��h�7�Vƴ����v�5
9>A�S��onWe������G�;�]�ݘժ��lL���i�!�"7�Ww�kv񰤃F
��T�xk��]w��ƴ/���Zz��_*�!�*�α��+�&�|}�`���u��2��(��m���]\S�����_�{V��ʈ�ǥ���U��SN�Xrڿ�cg"(Rǩ�H]oT��n<Y�r����p�?nh��v--:�JX�Xۂ��#��i��n� ���Z��{�2�;${CCH�����8*�=V�B�vi�:������4�����1޼m�ڻ��'���8��[MZ��{u�(��0���|�lf�kD C\�,�m�d4DXv�f�غ�|�����\�ոeIB�p�D7K����8M�Ɛ���_P�U��1��{�.Y]�v�J��Xׅ@��;�n8�޷��6�Ugw��z�z�^r�w�V�̦����7��HfY%�+N��ȝ׼ѭy|1*B�jL@�h��P�ͩ��q��M�F9���0h�8���]�������6'm����C�B��!�;S;�i���槕-r���p['b�1p��^�-�����R��[��©��$���=�Z�˩<�Y�c�����j$����:����F�CWusZ8��Z:����}�����2��P<5�F�V5 �᳏1��B���Ĳ{{	uu��g��4I��k���jN�7/<���9W[�-gl�����-���1Eج�5�v���i���_2j|��gQn
;�̛F�����}p:5�,C3\����*�Q@�-:��K�#��7zj�U�n��a�b����C��N;����lIV3p�]����ߵ�׿z��¢5l��bVY�)�EAmm�P��F�DV�e�KPZ�-�m�j��mURڢ��E��jԢ"&e1RʖKmQ�hĥ���QicE���#cj�Q-me�����R��q�neĪ%�)m����ۖ�ZXU�Ur奸a�mmb��[B�2��AZ"ڤ� �U���A�j[�,
�[m,V�mR�ED��A��Z(�e.f5���V�jJ¥(�V(�Umm�j��j#*
QR�PJYj�R���kKR��QYF���%����)AV�e���j҂�Qī�E�
ZT��h��"��
%�,)F���+Ur�e� �%Z,��-UU�cr�ҕU�X%b��Q[d�2�r�6�X�V��DU���,�[cm���30J�U��A�Rյ�Q�i\��(�H$�B�����c�^�H GS���KwL��s�=E�-
\3V�z�Z�9^��n�z���q�+�k�S�T����#��[�P<UE�pr7�DBb�Qbk�
c�o�OF���l�umE�c)}�eڣԨ���ۤ>�sI1���wwHtb�R��|����0EV!�:wq`yB�aM��(Ylob���cj����췊�2����.�׳Ds���6��:h:ݻ���"�8Ўot��f�ݸ`����pڞp���?B�o���տ_�(��R��T��]3�W=
��M��[��g1���X�47{<�����'f^����&Gzw�rQ�q�Y[��]|}�*ͮ#�{��Ŗ9v�X�W��ǆR=e��1(^�-�ܦ�U,NՂ%� \�x�Ƹ�E��j�,v�H���a=�<ڸ���I�~��G��BE=�Ú����յ��މ���\̑�f��	j֑��Õ��tZ	 �pEW�E�tk����pM7�Vp1�J����κm�;.m���)]�]{��s2gw\���YG���[�7�uZk6NWM�|Ap1�o�V��[��2�G������&�,�uŚ9J���g2�G`o�W#t��x��W�3�kI�����Y�W�S�-��I�m�Ԛ��E>-�1�KI(��a��-#*ܸ�~Uhj"_"{2���g�΅��y���ǂ:6s��9cZ��mT
iC~x-{Tigz��ooy��;��<T��p{��x1"7t�X�O7���-<�+����ݦr�3ٕ�Z��b��9�9o�e#�����DBv<!^�JbE��gu�73`)�2k/d^��,�����(Өӌ,�Ҕ���O�*��X��Y(k"&��I�-It�弅��&L�E;��o��P-��&�40�5�>T��}��*��n���pl�&����[aU�xy��Am:!�4CW�6f[�
�ꈕoq4�8nu��%��L���7��3����\ր����|�
�����բ^�u,S�;�|.�f7��#�n��f���#��m(��O@U��#�����Vm:�x�7�=���ɍn��P��N���s�(�zr��/zqD�݄?����6B��l�<��������6�n���^����V���w/�kN9�op�eEm> p)s"`R\�*��C8�p���ޥ�^����S��� N��b�W���Ӝf�|�]k�vs���- bC��݂!='�)X�	Ga���+}s4��|9�E��J��~'�.Ր�������k��Լv=b���A:S�Kս�y�V�B��ct��J8��ۛ�}ӱ^hr���2�+/n��)ጭ�NlC/u�$���/J��q����JaH�k�M	L�xa�jެ`�iQ�;u�W",�W�ݝ���;��2m�ʡշ�Ҏf��;Jy�ޢ�sDt�ghZ�ٍ�n�U�z�g12]���bk�oF�)z�I��`j��H3W��l�R8���;��,�7s��4�����ֲe8%Mǂ�H;V�)�V˖2�%�t�5OIk��"Rndc�Ȅ�5Nx4�ׂf��J����2���f�
�����&�t�]{a]�g@i��\dZ�AhΓFC�B
,��Y[Kve���d�ۗx���J�]e"nظkWq<�`��X}0��Tik�w9m�Uҍ�F�hyײ����u;"�̺z�u�.�#�ft!bղ�ؑ��= ��}�����tG�0�Qbh�U����(������ac��o��2�al�vK����4b��E%��2���<nݢ���B�b���&�al�ƺ]hxrj�"ι���5�5�C����^��uu�E�2��hP��ϑ�u'W-L��94��oo&�6�4!�e_�)�-���kc��=݇����7�=��{�瓷Ƌ��7�U{Hi����K��3=-o����̍�@rH��%����n7*���\���sS8o�g��r�B���s�#�շs�)��J�I�nP���U>/����mn%X��C�����]�_����m�{4 L�h�T��-�F�6���8th1�aԍ���6@[��Y��n�mc��&��f`6��$�5�,�kH%�Vì`$�y}�R-���e^3ۡ ��WD�w88�kk��H�����{�����D$��5�c�݄�舋m�(
���p�3J<�-4gȫ����Wې5�Lv�ڼn���V g$�U}�ڒ5�/�����ʭ{T>�j�F�e�~;�,�ȋ�O]9Y{G=֢�{ܬs9&�2%���$��{�(t����ڹ노�V.����v�O&|�X-<�i8(*�s�좳��v�6����5�O޼bl~����������CV"�NJ��s�SK�Ͱ������d���V{-���w�A0Z�%ښS+5ӳ1�aa���.�П��&��U�]��V���ۙ�:�rVEҍN�x�WHc݊���M�;���yB�e�{�(Yl@P-ttgj��[�˾Q܁�ܕ[y�L5qA���q��t��P-�C'X��C5�&�����M7A�CU��T�sϯf�x$6=0�Mp����+.CȁgP1j=糺��4}JW����k��X�p7{<����]'m�KH�^���;��$C���Z�ۛ���U���������E�iĳ/8����J�:��b�⾶N$3�,}��!K��`�4�5��V{�h{0u]��`J�uo6�cy}%jM�����#�D"��\ѽ�����t�L�{�G��*�Mٰg@�W�
Y|w����lh�w�l�]\�<�6Ik�����#�lvW9\��S���ω��2�߃�V�e��<c�j-6�󥎕�GR�Q�ǎ��og�r�VC�2���PMޕ�Q�{F����m(���PT[�ݩy.��9C�Up�%X<����se`G��[ɒ7����q�gl�6̵4c�4-���P�u��s�1u�����;<���gw�5��U�d�V?:��]Up	��TQ�3�跫1"D��!.у n�V����6p���뢢ǘYG��c'�~9Y�;6A�q���������<۱�u�R{��$qj7Fo�[�*X�Uǔ2|u������� ����*�^f����k]���!��,KN�|
��˞�O'kޤ,�i�C���^B��ܼ���dJw��N�ܣin��'�~8�u1zs�s��%R^�<�=~����W�	���l�&�ژTBB^9����ʉ\��0e����z�f�6���XWt���L�Y)�Z!<�[C���]����/ Q�<nSp��۪�f7.�BT)S��ךcj,M �EPhk1;���yB�d���o*F���Sʣ;�(aHwBж��l�\S�@c��;���"1���׋kV��7v����t�C�5��95�\P|/S�Q�.��d.A;V�Qc�
�OՕ@�q�c1���"���Ś���������f��m�cpZ!t��u�Ք���hq��E-q���l�GoY��&�q�i+�����W��b�(���c�=h��x��L0̬�ۻ���Y6(��ɶsj3�(ܝA��J�g��Nn���I�K4g�[�ѼR*�m0�:�ƣ�6��s�)GF��d	q����c�/�R�9�Яk)�Os;A���KSַP�q��̻OE{���bl)�&�'9)막T��������`�`����N��F����s=�^�2�nyRxLĠ�j�<���ٛ�T�'vn[�쪥G�r}V5�
�5��r��qC��Rni؈�M��i��gr�:~�vN��:KK�ƭ�!ֵ7]�=Ojƚ��<�s�E:n�Z=��C,����k7Mъe����"�:ݓ4�|�c�:�\��O�+����}�FW"i��+��U��V�c]�.���Jco�5����^T�� �YqH7㈇�F�Fc/z"�
7Ѷ�a����3~�^�O��@�(*�"�T�8�:.�1��;p�&I���ک�L�j,KNO�ao*Ġ���ʖVv\�g�7��=�z�qG�%
��y�@�Ŗ���B*�C^�.2)�:����Z���8����*����0G=�脘�-A�h��u���Ci��]�O�d��(]�7M����G,k��LD��UE3-=T�_�F�����o:TC�8~��-���}�
�A��T����n

�ޓ���B����׳D���5��}Ʋ��;E�����b�'�*�0���)�O�Ԓ�w�7{=oz)X�N*�K�=*=��@;F�N��D�)�m>�9
%e�1g�ة�b�k�+ftdo3d�klMtJ��XB��=̪LOA�J�+4��Pִ�X⹙��R�:=o�Fv��!��j	�n�����r�t�j��P�Y;d�M���zg��A��g;��k�qyTmN�ɽ����(�f���doQH�N<J;'y��v*;�c2�8�����3�c2�A���]4DfrR%a��a�d��1n��f4�|�*�{7hc~����d�����|��~����G}j�ژDg��\����\b���*�aU���Z����0�	�s3'��X�Uj)��\�mV��~Ukڌ�}4��WOt�n�]ɕ�l���U��3֏3�}cYv�w�
�.�H>�� �Y��@H%��orR�I�gwv����]j����mL�ga7gD^:!C���R�랱F��ͣ�3e8\��T}��W�k�F��t��̐:F���V!3�-�� �� O�;��n��j�>�u*����4/ʜO��k�� 9�T5W3��x�=��tǙf�Viv���De#���RR�= p�7Lإ����R0d�77�F�:��r̡UƠ������<㳶ra4����E�nWTW�a�Q�;�҆nr�6/t=��]Te��w�r�9ٓ����
��;�'u^ep,![��݁q���xkӹ5<��Z!���cmq�f�����v������N�%u-��Ě�em>}]�Զ�I�c�;36"�z@��U8
�'��o�U�:*�e�C­����u�u��t΅�_8j�0��\rH�5h"b�G�O��Ӭ�MA�<{h3��f`�)s�,�xg>�3�{!WB�E�)�O�v�7���^Ȣ��Ku>�I�ǐ�������{��?O+�o�&�z���RH��AH�t3�����f�<Ϻ+r%P���/�P�9�U1�r��S�~l��9�`t��U���V�=��g9RSP4h���Kzb���i2}ZkEs�]=�>]��t�A�L9ܔ l!��ϓv�oGeTQڃq�db��Y=���i����k���]z��^�]x"�u\E��P����jE�-�-[U�NV�p�M\[��'J-�L�K�L�D�B�S $��$��E��jEQ�l��+��+)"�*9���W0���93���ʛ�tK�_�g�P�V0:|�ꮠ.V�ư�[��dk�[Us���qP7g@�N�5��M�F�u��?S�����҃�Wr9&i��.�Z�cs-�[�l�JW}�e�-Ėv��=�yv���68r���e�%ڭ��c:P��xE�;��*��h��RJ��e,�5�u�)����f��n
xA��(�{���1���+�F��4�����I�;��sT8x<��1P���M[
&�κí!�f�4��	q�$N�|�`�6���-\�'p�o���q���to�U�S�.��I�"��Z���C;3���og�K'N�s�E@��me]:��u��,��B�3�o��C�S� n9�W1��Ѹ*я�ju��ga���Q�r�**T��&X��F���fY~�^��V��k�Pd����Yu*�����{o(�Kti
�{G*�K,f*X�B�#ӻ��c�����C��wtr�_{���?��1��;^�[� ;I�7�u㴒��X�g j����|�����A��3��y��D̒�e������/:0MkS��t��l�CNR6,�X�O�m
�Li��n�l��h}5�vf�h�B7�%8)���ad��򻹘^>���e�z�uv��n��/��j�:���Q�Wc�k.�*�mr}��Z[Y �Q�t��k�D���Y+�`n�=������ǲ�35q����T/J�}(U��G��b���R��|y�l�M�.� ��ܘ�>�A�0M�x����
�nDE��΢S�������M���j��鈚ŵ����-�+WY�fV�GL.�ʒ�uJl��8�X��15��K�W��[·3��v(�kr��X%tɵ����J��)��`B�u+�t��H��\%���rgޤ�T�ִ���qE�-ir�
d�v����1�鸭��s�3�-]��ݻ�ѶS��s�tq6�ƞ�}�B���c͚�
�4!ٍ�jļ.����Np���󰉸0�"۪E� ��t� ����
�X�IyHj�˦`�ȧ5D,�����]v�^��p�>��3�qV��t��[H<5�<Z�U�k+�Pt�N-$!�Z��%>C�Y�YS9�]Wy*�Y�;y���h�6��_�aH��/m�BC����c+SY��<���3+0ʙ����h�/�Z�v��^����	n��=8S�u��T�?[7�N^�uI �#>��uG���s���٣�kS�+Tz}jG8ř�)�K�&���v�ŭWJƺ���M \1�y3�<˸l8�\�1Z���� �9޼�ϴ�`�/'e���^�ZR�@SІJ�;�s껸{8��;No)����n.�/vd.�+�y�`*�V@�j�0���X�v��P&:,�K�mɀq�[r����*#���g.�f��r�&�F7`Z�i�����
���;�b�7r��"�'y�Q��j9+uw]��ZR�5�b�'J'Y�Ż��D�˷�y�_Ez���X�h@�h�Q������늮9(�����S�[�G�	�(U��9��UQ�E[QK*�RՋJ�Ԫ��*F��ڴ�(��Z��Ҍ��Qj�)څ�#իFŊQj�U�c�E��m-�-Z�L��J-�j��[ZZ���J��ՠ�mAdZ�QmcU*T�,�cQ�m�r�mhҢ�
֢�U�P���[�+h1m*�R�e�+D�k`���m�Ę�im%+m�km+U*fU�ZP��#kh

ګm*��m+QmceQlF���EKj��e�R�mJ؉m�Qj��¢V��UF�P`��(ґ[j�caZ� )U�F�֕T-�Ո�m��[mk)m-[A��ƶ��DUE�1��B�hآZ"��Q��-�J5*��-,����D����(�E�j�[��Qm�4h�8���S��X�L<�é�YzY���<&m�ϣ��9��aNT�݈�h��,\G��lGQcU^�d9x�WS2s�c{9*�J�R����#�\`�r��]j��=^v�F6��e^ wӯN$r'S$~q�B��\�~_e�0���г�ϼt}as������}T܇�ې�c�7Qۨ�Ar�D��wN
�*�H>�)�3WӰ0T�I�B�]���*n=0�[L�cA��P{��b�AD���HW1��&�E����qsG���>� �
e����2$u��t�AVMt艄��^��w�����K�H�U�C����?���EY}�dI��'DG��#�����9A��d�,wT��ž1�E�P�W�� ��#�N/G��x|�VwѰq��Fa�ؼ)�o�L ��,���!�&��P�gvB�&�sp��e}��Y��f�n�8O�+Ǒ豆���nb8oP	U�oj��y]L�(�����ܦ�p!�=���9
����"q�3~9F���r�v����b�)��1��Tb���w�\��p������=R��Q$	�r4�����_�=�Q��*aϲ='�,1Ty%���u�%�0����p��"�q픢�Y��t�ɗ���S[QѫG8؝`��v��[�����ή_�T�/z��aͮb�]���>B���0�M.����wV�t�jR��݄� �t��֧sN�ԧAY����9�fM���$�O3�q�;�=�L�7����t�p lU��G̝��*q�`L�f�s�[S ���X�+�����L��ȷ6�E,
O��0�ĸ���������5e޳�|2�-5�&v `�pb�r:�N�h���ǻ�>�0Ct�i�V��N��s��;*:�ˢ�>����ae���(��U{OH��,����#���8�4��
�N����iR�kj�~̭�#�F!1�!��\�Yb:����nx\���P�h�YʲH�mL\zL}����y�J�Ւ�ǈ�J$�mH��<f2j��H�Y�`
<o��;Eq�fޘ�o{y�������R�e��-�v�,=R�!Ajd�즆7�-�G�B,2����~�z�G��:&*y߸���� ���
�O��OA�X<$����L�;N`aBK7)��Q�[;� �ӹ��
��C�f���B�p�_{�&�JeUa��F��P�·��!�������Nv/Z��������m�R�6ksgi��ޝ���H�]��㥸��eu�[��m�8��F�������tXX'q\u!)�=�*�n�8	D�>�pv�x�#�V�oo��vf�y�TxeD�:`�i'�*���&������q�ڰl�ʢ\�ū.޳fܔp��s�ƻv�bV��C��z�
�j���v�����pmBۦ�����x�*:Z	c��q*�������ڀ߻�*���)Y������{���5�)_��������w�N�ݿBU�V0_�V���.��v7|�J�����N��{7h�����������B�����B�v61�;Ϗ��9��C�7��1j[�Y�p��>�W���|�G\���o�ڏ8��tQͯzh!׮����0�|��wZ��0��x����Q>�U���>Q�5Ӻ$t$bJ��˽�a�쐩h�
xEMF左4��ICfZЋ���3�b2�dE�����{�S��%�3�i�U�#1�ѯV��ۦR�N5��_|���m���2��zۛ&ԅ�k!�4��s�3�51D�Ge��mDx���˱.�E�F�w�S�;^
�h��
�L�ٺ(��!W@��G:�8k��O��9�Y�X�K�sU���NT�'&(��lTC���l#UG�����P�A�.m�����mZ7��R��g�����Z�/n�8z� skFQ����t�V��M��wz!C�q��:��n_}�WG6+=3�t���RU�BU���FE@�Gw[���Tg݌�̦_����tQo^�=-ȉ9W�\Uin͇9�Y�r�lW��m(�;��d��X"܋���b TL唢���;/[r��#���u񪆝�:���������u��R���]y�	���)ѽ(ޢQ��V��V���{gv��� e	�����@XC�����ʫ^��j{��u��*3ؤTHl�nvr���N����cO!�O������\��c��{�2��	ga���d�6sM���E�q���A�QF���|�<�櫺vz��H�P0�-ɋK�(� ,��
yTt�aM�c$l0u�aP�5<�D�����5��>g�c� �Ge�ٗ!f���=��o%<���3i�!�����qw�;�"�E<���> >	�Gw�Y��o�m?gp[��5������Ô��2vR)���@����E���tDx�x({2>R���ͥ�=[�L1j�-F�1����b��8��f��o��R`��� �$��kU=�5�S�*B��"d�>7#5?�Z�<vV.�Zr�ҍi`W�����[��]M.�䜗XǴ�B��]�����ķ���+��f=�Dؑ
2�4m6�U5���]J�����O���h�˳�^NW�n�2�L�hΗ)�՛\9���)�	�:��s��uj�G�Jvv��U�	���$�/��Ɇߪn�� .ZǑJ�����p��.�u�q����=J�8.���~�N�e[�
�jC�a��T�>n�[�.���3X�XV)�u]��)}{R�N����V�V[��l܇����%μ�DtW��ɝ���T����q~�C��uc�@mE�9	��)
VW5R@��WB�h�=��n�)p9�wySx���a��]��;�9\�:ryF'��a���"�D
��>���c�����U�=^v���"r�2k1�t�F<�Z�J����d������t,��m{��)1˰:��d3�\q�蔮����$p٨jgM�N$R��f��``�����e�*pC�S=õ���C�|�p��k�}0��U���q!���UQU�~|��S�|P�r���kt�:o���i���*���^Έ��@S�X��f6m�E��S���q`z����2�{��lq�>���iڛ���Ed�,_��N�@o�lѰ�eן�!d�[C��x��'y,�.y�Q�:�j�ȅ	g4s�wں���ȇsc:v�W�-�]P0l���$����;�dV����*�Vd�*��|�*6����N�Y����^c݅̔�R��CwUk�ڹ�D��&��˕5�lT�i���]]P��\�U/Í�� ��̮��_�m֦>VX��[��w/L��	���^;�Z���O:�,:�\0�bz��Xv0��An�.����s� -GM������S�M�Z����ВO[�{��L�0��K�u��?���l�h°2k�<]!���bSՇ�$��E`����;� 4YQ~꠲v06�T����*��s0���]]	B�p�1Ə�S<D�|$~��^�jE?HF�2-ߓ���ъuU��ʉ瀨Qb��U��L�,�J������JU�`���jU�x�1ڙa�-ͺ�]q^�|$���:�fNı{��(o���C�.J��t�ܪ�x纂R�K�q���n��:8h�S���nYy��
�>?z��9�%��8pppװ�5�<}>�=��\�qW��n�B�z�43$?,�Dr�2q��bi���Y+ʝi���c�7`}�d��B�`ˇ���;u����.tr�p�pcҥD��Zdt�34/k��<��:��t��-�>�@װ:D]z%��^��F��((�����չ�|醍Fl���.B�nn�A����X�-��M�r=�&�_)�a7�fvp�wN�-�M'ղ=�n�:�Ŵ�E��#W;��R0�r��OlI�:�є��L+��8C�ڛ@m�m5�\M�d��N/�Y�P��'.,K'Xi���4z�*������e2���̂�L���b��5���AFDL�Ց]���y��=��������k�U�/&�E0�.]g7<�Cnm���3J����v��4��]Zhx���>���(p���2��_6�i�+���.�ʉ��
�(X�SXRs�*���r�?yO��c��}�ּ(�J�Yy�}�ϑ~�Ӗ5�K�z��.�  ��x]��Ts=����_3��ۣ[�_��(�y�sz��(���hD��<�_Y����,{�è�P�򱻳me�*�.��S�Cޥ���!�N���Ͻ����XU{��l�3������خ�c��u�^F�6���4����v�ZH!V;�ȭ���+1s�a8�����q;IR����Q]�f�����GX���F��v��)�ْ�C^�.X��u��̉�y��3E���!ʡ�n�d���ν#N��;�bJ��w�*]ra.�tEڕ�b,���af���jX��Tr�o��ر�-�߳�c��c��N��n��ᚦ�WN4z��9�閦H����*��]��J��.c6��4���|��()��7l�Vf�g=����%���J@z��܉sٯg[+f�݂�U�`9S�bUԙرԫ"�z�����I����u�ҩ�Ɏ���k���3�q�>�
��ڑ`)�/PD'�+�%Dlةz��,�5ûD����=�qL�o&q�_o����G��Bw&�o��.�}\�1Xk�����Pi���}�K��]��\O\��}9s��NC>������	�E⊉lTC��d{aq}�4*(GN��O�z�{����{��O��!١�Mswу�����D�%G�K�F�>�µa�g%VǫpR�(�r��w	�Ƕb���2y��t#��Z��I��L�r1h�4 �P�,���_�b��򲸼�ס�Z�^�� ��;|Й����{�:t�A8�B����0T���= �&+f��3�*���
��0�֌���fN�˞��n����D*��(�@� 5�u�C~�{�>)n�uH�.x��'[0aUu#Ej�}J��Ɇ"���
�;�BR%�F��D�������SӖ��b�|��~��7���o�J�Ce�V�'�:}j��Rn�s9CŖ{�{�"��o��v�u�*��)v�<�im������k�[һ�ZHq��$>�+J��F�t��[i�˥36�s��rU��D�c=1��Vj7�����U�]��I{ǳs{@B{��E���(AaD3������͝񩆓���y�?:�:VDR�հze�j,wT��VI��$_+
/�)5}\+<r�N~2��j�՝�f8�4ו���ޓ�+�u�]��ʘ���;>��:���Պ��Z���ٯAݜ��e:%�lk��Wwu�+et���K�ƸV�t����.��0pmNC�ee!���v�� d���X���U'������+e�c�+j�*Q%�>�>�b�@�`\�������a�z��3�"�t��:mH:����\�!�Qnq�;R��1�41����@T8d�''sTZK�Rn{�]?,=�,e��/�K�x�ɝ��&r��tK�%�È�Ln9�j�{�k���T�1�HX����D��~�M�����T�J�~]�o(:)�I�ҷ��}����]����\��8WD,��y���/A.F6�>���DE��u[���I�G��~ܭɡ31̓�1�oA"2lpB^����|kＡ�t=��n�W�Ӹ��S�E՗)pbU�I���y��9��J��a��[Ê��4�`�`Y0ؼ���-`����]Z��� sH�X���g{�,«.�sx�����:DF��Vb����~;w2����-0�	���0U�)�{՝�P��	<Y�QΦ�z����۪�i�4�ĉB�K�;9b._��(�t
��؛=��GX����*X�L> q��oR���b���h���������	��YC�F�,o"�䛾J�u�~��F����0� ���T����E�
��Fˋ�S��/Zn6�S�D�uΰk#O���F�[���r�{��(.���1�F�V2cT��=b�)�5�~�P�8��:hl_g������b��vMG��<�!�\�2�H�����Kw;�=���ͫu��
d���[��A?y�g�fKs�u �dO���o_@��K'�tw0s���Ԏtё��:9
��pFA�g�9F�����R�Fv�U��Y���)D[(@���aU��ڬG}�A��T5�����}����[��ݱ\�N8�D����+�Yp}���<i�-ߓ���ъuU��ʉv+��z�m�쯾��C]d�H��+u���P��&�/����k�7�u��S��Y;�O���6�ۨ�	!I����	'�BB��䄄	%�$��HH@�I!!I����	'��$��$$ I?�HH@��B��$ I9$$ I,���$�$��	!I�@�$��	!I�䄄	'�H@�l���$�$$ I?��d�Mfzq��Uf�A@��̟\�"o�<�( 	((	IE(P
 /� $R�
)"� D� 

��
�IB�
���`�*�QTT�ԒT��6dP�T��� ��!J�U)$hj���Q*�KֈB�P�B!J�JR�$@G��(��
������!$�*�
�)BEI*$!URA
���$T@$RE
D�T(�)T(
Oa�D��*p  ���w4UJgI�*��$Vmi�E�N���qU)��k���QۢwM�[emݛ�p�F�bΕ�5��M��٤�ֺw[k�M2�nQ)(*�CH�D���A>  ����AҙÍ;EZNK۹���gJ�閶T��ʴ魫�.��s���ӥ-�rۦ��wA܉]+ �!�R���cwU8t�M������"(J�IBT ^  ��)ٵ�gFn��J�)ڋ���Wn��BJ%�:=ۨ��u���s]�k�<Q�{��GG�ޥ��F���{�E@ ;�aE  �PHT�IIB$�D��   �Ǝ��(�we�( 
 yÎ�=w����S-u�`GUλ�c���P��P;Z��8N���]�Ӱ�]i�C[7	�K�(���� ��lIE�   ,���V�uTpk�ѵ�N���(]wf���55n�T����-��Զ읎�gT�C��˔�V�i�9ҭ��D�)T�T���"*�H/    �輭R��]\Z�n�۪���ۤ�:H۹�6��u�ݓr��ژ�+���b��V���t;��͊k]������6S�*�* �AB���U�   1���z�u�L볪qNQۤ5ո�d549j�m;��u����s[��n�u�s�m�u�uv�]���ۥ:�䝮�YU�qѺN�]��ӹ$�*���PJ*$�$�   fv��&�;��]nڊV�mևg&�r�ej��4n*�֕ݣ-]*U-���Kk��I��Uu��`�t�*-���X3M3��ة$QJ/��*��  c��SZ�k̻�����Wk�n���Vc�i�]6�����]Pk�4Wmѧ;�nZP������Q�'k�a�ڲ�v:�ۭ�HJ�4ԄUT�J�   ���kI5�;!����Βqv�T;m��J��r�����Hv�V���֕wU[�[��w\��GmS�㫷[�ۭ���c���w�O�Lʥ*   "�ф����� S��L�SM4��)�A�J�4  T��j�H4 h I��2�L�0x�o7��}��֩��p�'ؙ��eE�BK��w�׏���H@�t}����$ I:		�	!I��IO�	!H��BC�͟���7N����tuN���V���H��ͺ��Q"N拻Kni;�AJ*�)i�c5�67W΃�Ⱥ��w�����ͷn�Me�[�se/�thV�#V�*�;�c�KE��yI[X/6�ocl�@��qY�Y�۫��Yyx�k,[4n�ff��yI�[��m��O�G��mf�²�Z���WQVd��-�+F]�b��۠a��G�n�����H��efU��:+	Ē�!Ya�5�v͋VVX�V�	#�$P����K<с��)�-n�f��46͍y�������ɢ�n�ɬL��Q#�-�٣�W��䧀Tڵ�� Q�%m=�%jaZw�UYW6j6������@e,�vU�W�p����9�K3Y;��MEr8T��V��sE�#@��%[�V�2��2�(����8I"��5^�x��,��C�%^�8,�YPim�!a�[��r��� �F�-w!z��$�6I�d��QQ˪Z��n^b,I��Z"��-Q��G&R���] ��f�d�Y�A 0V]*B��U*�׵�*\`SÖV�1����|��^ݔ�.n(K�m�� �hՃ#�ѡ��7�O6UZ�m�c42�2�;]N�i��G��k4EjӬ���a�وi��ۼW.�c��Q<1J�ڼh2F�Y����&�3kp̩��lbR����I�A8�\qau�8s2<Q��-�٥Q�qG�i�m�d��U�f�AoJ����!=[a
̶��#F�V�U�7L����0�	��ݶ��P�� �Սp��QF�^!���8.@Y4��y&ei4ཫ��*�4��dGu�`d�ZrL���.j�n�
���e�1�cE��5��nT4&�w��T��	�aL��KZ������Րhi��ٔk��d�y�;Wj;B˗�^Ci���H���*7�RX��$W�ŌG3��t;~�'y�#�
>���4�uq�b4�!�
h��X�������E�ٺ^�!�t�p42�m�n[��cH	���d��໫|SV*Ԋ�@cM oQ[h-ʽӦ�D!RR����ݨn��+���a���X,�B�����F�[h��a���-�H���r��E�;��\�	�m
	f���8^VG��	3owpl�Ě�՛���b!��r�#LG�-���}��aO@p5����.:��m��Ӣ�B��f6:,��nB�p�k��h�r槛O.^4�i*@��������XTzL�BغzcXÊ��p���wj�n�E�b)�+���&,�FlK]��iz�ƥ�.ʡV,ޓY�:��L؈�zU��SV,���"�3���(n��F�����g�;���I:>�h��ݱD��͖N�ś]W��+A��^���q�Y*VҌ�ST.��E�Vr�����©�x�OZA�9 ����kz�,��ݮV�"]:���rM�BD��N�0p��n��^�x�%n�Ͳv�ݵL��J ���J�^�]@m��kŴ��i��[D�u�����@�/Qɗx$9.�ܕ��
�IGZݪ`��e�231�/��:�+p��"��MX����S͵���޴5�T���m�j�����#�U�cSa��Q���c��b���{+u�� �M]��h1h����m�usg
uc��U�mm��;��B��i�ûvp�R�7�G�zv�R<����vN�����Ż�f��kV��ۭ��ݪ� D���2��bBj�n��U�(B���j�V,;`;J�&ͩx�l�.�*�Q��S��]�����B���ǃi�К�ܧ��)�N�����J�;J
y�w�[�����\J�[ɚ�zF�n��Ast�Λ�e۠1L+�4Z�)=DXG�Q���s\���J�����;W�ҷo)�Ĕ)e�c/��D���w&2jS��3��B,��w����iYZw�0�gFV�� ����;��d �U_��+ݻ�x8���g�5V�m��Ѐ��3tqлOB�[����X�8�zc[���ź^j�Jc���R% ~)�.�c�Y�J�l�F�ڻ��W��4�j���U/�Cr��ͷX�����-ٰ��0��,=;*I��[��J��5��4X���4!������c�eL�p�WZA�.����W+$X>f��K��)+.ܥG栻U`�y����]$�7��x���t�J��Vv�����O�u��{!E���MWy0]�����TE�a�[b�f�m�V�h�a
�Z<vV�����6��~�D�Β^�!ao�QU�i�U����x���K1��JF!�6��V�vVe]�k�ո�&2=�KN��o/kM^\l黦+)[�m��-m廥�f#�c���shH��B��Y!�qaA:=��ũ7��/�,ɮK{�� 8iD��N ��;b��31�H[��yC(�U��J�~�/f�B�Rʗ��2*����m&�k�N7&��1QXȉ�l�R�PhP�v@h���ͫ���$��<;-ah�7x1���e��a<�X��]�W�{�P�ҵZL6��)�[6�k2F�����MD���b��#�7I�s1ʺ��{�E�����]od�>�wRf]4��k2=�A6�nZm�ԄW�o^�˕� ���ա-.wiV��e�)��(�s&��·!@��ڨ�fԈ%��0F�  R��%U��x�Wێ�(b�R�&�7Y��+Y����b�(v�Vk��&0�Վ��U�Oy*����Ga�b�+#�n��雬Gm�YO3�ZE0���^�Tҧ�c�hK��)]��y�a �5��f ��S���$3`�1nɗ�h��E
wX�`Y���;�zӁ1zʍ�kr�U৉�R���$M�8��W�����9�Xee�\�gk�M�Z����y[��ma�R�wBZK��Km��tj��[J�*�`f,!Zi�eU𡕫��6�k����9G��b��O�i�	�n��輫$PMj��7��eޕ{�0��+y��p�n�A�����l'�zQ
��ݸɆ�84f�L�"B�/p
!�j,��j�;����B��ך�%���*�"Z�kv�U�O5n��=te�Wr�O�4��]�h��{�������PM[�Z�(!G�_-9w۔�j'�.fd������mhb��P6��V�l�9gT*^���KƧ�pm*e��x>y1�Y{+W�.�8��%�fE��Z��0����d�6���;)2].��n���L*ɚrb�+
����v�0����l2��S[�-b��vJ�R͂�d'lfV�Zm˖�7�n�5Ț�/����nmu�{���r��5�sie�J��!q�Wnڻ�7r�J�֒��O%��t�i����b�.�tu�j۫��cZj��7��sG����a����ib� ܫ���/P�����k,e�[������e*��-m�F�V �j(���L1�*���;h�vLt�����v�W]j�Oq�-Q�k7V��א�2��ajDb��Ҟ���Y�My*F�MXp�h�U��l2t�)�M��.��攘��M��lA���Y�R��_�rK.�Vf��m�s+����E�E
�(^
.�ө!�	;y��W� n�-�m�����r��Hec)��83k.�d;���6�fEa������k���'@�n�)��h[^����sb��qnj�#�p�O͓2m��7);�vS"�-�J5!�٣%Yj���ӫ�[T+0��2m����x�g�L��	�*ǗI��F%�;��Efe�73�.^i�Z,A��+c��g5R�i�o'G7���&�����m��ƭ@mݪK��|��[��Zޭ)��`%�P³X��ivn$B�\�<��w�F��Z���`��6�Z��J�%�[���<{��A�鎉�Rb��z�Z\�T��v�[���Un�s-�ݧ��7WZ�O �>x4)c�5k�-͑�J����V��Ʀ/'��cY�Յ,_X4�i�tɮ��9ZE��-�)hY�V�U��U�{����Kw.RDL�7sU
ݧhCG*I�wkk/^`KUt�bb��+�N=2T��cF��{�!��:&�ܡ���ސ6M۔�cb$6P:�n0���&�ݔ�U!�+'^�%�+]K�ܻ��ta�Mj[��'��Pyuy��
�I��ޠ
�np?�iS��ߋa^U�'tU�c��x2�ɔ��ޜֆ60C�U�H�`�s�{d��tT��w��ip-�Z�6���b�v�y�U���5��a�)A�W��K�����%3r���8ҷz� I��ҡD� �U�7����;��C�Ϸ1�`���7������ʛ����mkoI(���%���[P�n�f���nv�蜻{b�eˬ-�jO��X�E�f�] e��F�p��%�*�{P3�%)��XW����mӢ@٦�h��b�������ye�[P��5�0�
ρ#*�:]9��(EI�Tʱy�Pn���3�.}'
��)<jh��ʷ��-��*>gU�`J9c4�[�b;z7#��\R��C��q�g2�)*���I,�TA
��-�����C,���#d
�(R�*�� ����Ҙ�,��rn�5a�U��3D/�'i����ő�����kl�	?[P[��ܽ��V���+j�����~C
Y�ssh�8-�kYL�kkL�/q����EhŗN���nmitu�5�h�F�6�ӱ���X�;��o F���r
`��Tӑa�0"2)�E?�Ǘyr	!�e���fTw��n��B���#�����i��kV���Bl{��*F�k�i�5rnU�(u�r���WX�ͩ|/�鲉VCW�-�`�g��J5�k6����-5��7��
z.�:�́Iu��"��-���,����Y��]j�ʀ��<`k*]�f���象�.21^�I�w��[�ʉ�S����(t�E��i�˫;�fK�9z�Ф��^�phl�ĒT�O�� ����!�%�k�5ǆ1R�Փ	
��i]��E
YA�ҫ�⯫��3F��O.�(�P�-ڔ�7%�]e�������6�%�VJ�{f��X8�_5��	�p��ݭdw!�N�W�|�w`�F�=#�_l�F��SM9w`�骈Et��y�i5H4D��Y[��͋N��ׄTYI�vF�\�tn�B�^Y�X~Cw\"��D"V���ٽ�Æ][�N5fط���q��e�[� �Yu��cq��b��P C�����2f�=[�F^)�U����̴��G�MBA�qy������ A�^�^�7�)��+,�fC���53&�yV���62�ϋ �Br�dm��a��/c���^[��u�R�2���W��Ë'�f�1��uM��f�5�I�x�B?4��X��Yi�"���H`jn�b̹4[0��V�Ț�w�i:�;5�t:�l�u��Y�)x����0Mh,tjLU������Յ!��ܤ�WXi�{��]��Y�i�{�#�W���r_"7sp�����<yrlt&坠�i:.9`;WXAu��u�[��ДZ�(���wd��wU������V�f�%��]l&iˣI�J�ǷtXO 7�-*��oF<�*���w	;6�l1�ܽY�o�T�!ǳ(B �y�j0�ݡJaPIx)O]	_%�on�j�G��"�b[���š�c8;�5�"����hЇU��dJ̴-;�h�`�ܖ��@U����Y�n�g�V�N���՘Z�%d����L-pd��3o-)�i$�t$\L��d� pˊ�]��E�Z�Kp�ǹc)��c+I�q�q��0:�CVh�m��G��i���͆�m�㢒ʌ�(���i`Z�/(nA�U�חt�Q!.,��%�1<�K˭v�Л[�7����j9L�[\�B�UkW�bH�MNa�x�u�oU�Y�tҦ�i͚`�;3nV�n��T��Q�7��R{�Jw"X�A�P������Ù>[B�[%�X��kq-�D
�r�T�v�K#���Q�^�KL�B���"ӥ�yysCyA�C5�;�f彼�0-�4���ܣ�L�C�Z5����ߎ�z�ٰs%�PJ:��AX_b�km���h��:��6�k�M6��Y굠H����Ay3#0�0�KF�����amA��P ����49�̗lcǺ2k,�(�K[Nf9��Z��C	�ȳ��X�p�_)�L"ζ��b#W�^��f��ʲ�Y;XhI����� �ݺ�Edӂh45��.��r�)�&��(3��րӊF�u@R9�u4���Ѧ�oIhP5�������m�1=��Z��fn��u��{Z`���זk-]��p�z�H8B�j`�[���7N�⼊Z!I" u����Q��a����i:����	Ж]af4���&E�ƥmփw�wNT��$m�5e1sVR"��cS[�J�*���{���	���ΝD��U����ml��(�� V���Fn��ݰ��,��ø[���ʔ)U���W2I��
�8CA����xE��x���7W��n�R�5�e�O*@�{�#���Ǜ*aɫqcT@-D�m�j���9��5^�<�a�j�%���jI�OO���PN��W�:��)A�����b�m��Po)�ȥ6��YV��Z��u+b�%^�� �Ь��e:K	3�оu���t0�l�}�i��4�f��Lˀn<��G0�X8�)��a��TF�ڕ�%Pɨ+���ӭb��w�m�^��?�5oq��3&�dјT��(�x��	:X��"PD�9N�����ڶ�B���n��h�{t�j�rB�5b�\ؼ�[l�`L����}N��@�]�v�����m]�.Z�n�B�װ謑�����78>�f=��5[�AE�N\uyy���B�ϕ��@������N�f�3]�7#�zá٭.=��e.+��|
�e�x�P�̙7�a�ͤ���jқ�{�k�I�nԴ`�$`8u��+N���st;S�`R�YǓ����Vb\l��i<��A���)���G{OU��!έ��۬���x@�7w0�h���@o-�sM�=�S��X���=��0EG,�GWJ8��#x���qD�ޖ35���/��6��㙜rqN$C�UvƼN������Q��6�2/�d�M�������"�L��۠�-���I�]���s-�z���X��Y���~�)mCq�qN�����;s+�l=9@�^i�Z2�7q&GIɃV8������s���^�Y���ۡ{�n�:P�u��r�Z����)�����R�7]fMŏ��u�
�-���T�(2R�*����c�qU��2mn�:,<���1ch��2͚D�B�냡J�x(�з��R�e���P��Q�� SkM#���(٧Zr��MwZ�e��}���w#�W�f:�?��%�q!kqQ�0�˗�۫���`t;�������x�J��Hw��>�Ϧ�S�|Ue^;P¦4�1e�s2�@)��Q��ܩ�����f`���:�dv+R[iN�ކ�y�*t�G��p� ��4*8��2in�;�]�Y�&�t�d�O��m��++'�r�V�(�p��F�ݜ:��6�i!n���-mϵZ��׊T��ו�f��wpI�>�P�n�H�e0E�&��˥��-z���h�ޖ��`^��T%�Cq���X�7��WO����p�b9Mݼ�ī�����*� xv�T���b�twvFQzf�o:*�Vɖ��ÆKv:|Xx�ǒ@�n
A�|�SH�Q�/j����W�8	���	5ڹP�t�N��2�
�4�l������U#�W�oC$T�if�j�\瀍�����2�1�18��O�^ȣ�
V/�U�˽:��o�\o&Y�R��f�b���P�2�Xj��rej�f�̚.�<+0��h�z�) ������b�Iޣݢ�K��>K�P��m��9�m�ؔx�s��9�S��J��q'����)}vZS���!���6�LLM��I̽����ZЮھj�5�N��uÛu���9�j��+�J�w��%��=W�w�^��e�0�ը�㘜�>]y�l
�/^}k�d�*�4)>a���c�Gtp���ak��,f*�@fRŷ�j�V����,j�(o�u՝�=�
�ב6ϵ]-����ٶğ8��Ku�1}k]���e�]�A���|Y��m����"V>�x^���k��Y��=hк�q��*@p�O���9?�#��٘�h �xH�N���`��恰�4�2�Xjo3�[���g}mE����w+ν!mA�����9�\��N�-� d���]���,�u��v9nM��l��	��ҫ��&P\��C�R�ٵw���C��P�"��9����e;���<<}�}YCy�=88��+�{��fa���F:�i�IZׇ*v7�z��xM`fZT��8�_�]5�ST�h��8�@�w�jbԷf�5
43�հ�Vn�H<���	��:�K��5x.�M�h:�: �P5���;0�wJ��{��J����Ժ���-�|8uƾu��f�0�'\,�Y��k�5�A��\F��*ؗ�+U�^WW"��N�b�l���4�`���q�Ѷ}���c��Dq�d�{w9m�F�[{�s����X�F���s
��e�X4Y���r�w*g�c�x[պё��7�E�ʆr��ܵ,�z��'S̖4���Z��0&����؝�5�\owpdv�;���c/u�����9g\�ٛ���v��Z0�a[y�88�4�V�7wӌq��O���6������(U���J[\�� �]��k�j�3|^`Y�8�EŘ.��e>W}��탹��T��y�f�s\�!����B�	�Ve>�I]�Ɣ�*�U9���f�gM΅e֜�CF#4X��@v�1C|� C#_�p�̭Y��.vغR�n=�d�iF��&�ݲ��$�lx��U�gN�W{�[Qo�|[�5|�����>��wk�f$,�S�Y���Fג g]�M��S�.ff�KM�dYKo��7^�']nm��Q6l�7g��XS:tR���C�O*�A��#M��#w����L�(M۾��e��˸�N��l`�ЕK��CYv��Ji�6�u�@9_ܭ[��)��X�}S.V�2;`<�e��\iU2���q�������/6��i��d�x�d��Y�rR*K�o�:�XZڜ�'mn���Hj���҃��:,�������R��`��n^��,�w�#�p(越�4����բ-�H��\�b2�̐>�ۏ/G`�F�z.v9�����3Q��0ť�ͳ�esE�Ja��(:�<s��9��ѿE�Gק����Bo;�]CvaV�.Ou��"1���m��W\NH-WT_L�{���)sعP��'�t=�e��^����'�v<�H+o�p8�}p-c$��%u�{�4+��И�;��.�oVGӇVw#Kp�7bjl�5��qL����uvwU����LMy�mL��\v��a&�Vg(
T����Ĩ���+H�����]XAg�a^�k���%2��W/j�!���J֎Ѵ�G�vW\;����Gc�A���f�Z�M50�r��<�txX��5`��*�"i�zwp��T�ֱK� *-�;�,���5Jj��s�d�T�]-����yV��Y���BP������-�sݦk�on����I�jj�Z/��b�"dܝ�y�U�}*��M�L��(PgV��X�de�C�0�Sf�F���O��¨�z�tFv�K&â�[�b��cg�<ϳ�+���`�4E�,�̓����:��%a��<��h���
�F-�t��3A�S��ķh�٣��t���^��.��Ӧ�`+s���V���r�wv���7);7�^#(N��L&�y�0���g
�C4r�Q�j�fMV�Na�gb<�~4�A�ܾ��Ψ��A˹%�[ԝ�4;zr�X��$,�H4��Ɏ�F��tS3b;�l2��Qg
�×p��Wi������~�����W.���`t,ۏ6Jp4��@oj�����u��R�����ܨT�x�jW %D�B,Q�V7���n<���h�f`=3���!�3V��}��`�+�ATI�DbFfC�.�ۏ�Jq�d��t�H��^}��e�w/r�!P3��vY��+|9��d�p�]+$*�o;�cmk���(a�.DQǊ�]�2�&֢�YVVA�0�������܇Xˡ���G-�S0#9�� �!���fVZ��Eܜjѽ58#�)�c;2T��� �=�{�kXnk'^�tȐ5�|�z��ȍ&]@zk`Ō�������n��4W[�Vjr��q%'N�'�J��ഷ�,f�Qcw+,eb�P|�����c�:GS�t�e�e�oA�<�_���a�:Z��br����Sf���#v�z��{�wS��7P�����=DJo.�86�kي���1��[���gn�X���T�C��,:^eM�f��V������K2jB��Dgf�h���Z�� rݓ�/x���}L�}y�4�̶;Cᨀ.H�'#���3�����>{G4̏�uu�K�!��黤6�Uq�2��&m*��u�P��1WC��&~GW\����aֱ�v�]E@�.8HYO�^N]�%ݦ�^�'�/%\� ��]�Z93����Jhi�Z�j�E��!�.�6�d��xqP��ϠH���hcG��U�Yt`ӷ�na��ӌバ6�)��]�L�q�uШ]Gc�˂\9N�){Jũ���-��I�l�f��R�Q_X�覭U��4*���YYP:�K�]�)�̧/e�m��C�2�P_t]���CԲ�������%�tll�^�E�d��.���Ih]�6�W�-҄{[��;��V:{��v��������%K�L��ʇd0ɹL�u�4�ջ�$oEce嗚rԔq�o�W
����c��Y�r��a�5լb�RT���<Vł���n��"�+�Q`,,������]���E�z��Ÿ��s��Ԧ�j�D#|��ˌk�Ad�����)�y|�;z���$��r�@��guXc���1^��e�'�ܫ�Q��Z²6J�ˮF�Ǩ�1bog+L^(��%�uV���o��to,pŜ���M�d���'�E�r=��?9���Y��6O���f{�P9]6�u_$��]H��Pj�Kt���ٽ���&�1�p�e,s:�����`3�Y��;�OZ�ɚ���H*�wα����j4�Xf������n�Fӡ	��Öh� N���XJ�[ ���������.�ջ�{5���]C�:���0���ܥ�j�w�k]+\)�N�2󂡹�_F��Kh�r�ŋ��[n�Bd�:FV^r��0�&V�
�b��rr�]#E��+:7H-��,[����w�Wm�Q��)laq���=�ݴ��'J4)�C�����m;�W@k#F��ʗ$�*��c�9��b���Z�.��uKf�w4#��ɡ�Wmu��3��\�gtnآ\w�dV=[%�е�ػ�T���&�>R��!^��S/�j\dib��2܈/:��IT�b;G>-vJ��=���U~B���_��TU��Υ��8�8�ʓ���Չ��}�;��:n#��ŵ��K{�4
dKj^�fª=�ůo���aʇQ��NO�w<Xk����zv��7�Ag�ztTn�G�,����`�[�ԣ�8��B��7����/9��u�����.����k�� ��vei�J�@�sN8�˷�VL7��ZH����R��;�md}�4����{6���6$R���a�|�㌫�E�Bs�Α�r\�Uw:���]߯����d��B�j[P��wJK�MF�"�.�Ea�\�L7�s7� [�&x+ϱH�T����A��	t��M�_cAﶇ^�3*�dV�d��a'�
��43;9oeILk��H�l;���ܗuy��^:i8���Ԧ�A���V���HH⏴:���6���)��a`lc`�;'�ft�v��ʖ�^�B
$QgU3��(:j����(�컂�%RՋj�|�����S��p�7W�-��/E���D��W�X�ou�[zŦ��ߢ�ل����=�ؒ-�.w�M���W �a�7j�]71
��]R�$kx\�5�(�V]���<h�@c�2,; 5����M�UcqH0Qoӑ�
lwE�"m�+i6�ʾ�+{1��Guv���UȤj(pK�����L���
ݹy���iV�[+���U��1h;���5X��X6��2��ⵝyQӾV�m���l%�+(�JMy����m/�,z�-
�,����J����� f �t�9s���v\�.�WćdΰΛYI �;9n�b;LK/M�&LGD=nL�"��͹E.��]��UӮ890m�s�����N�z�4�$�(a�;R�tއ��o�F>��t�
��Ӷ�^�}Qm(y���'�q��'@g"�;HF��ӡY��8��h��Z�:>W�]픶���uAK3_*����0$�]��RjED+wi'�xPx%�j���gs���]H��]��I$�A����t'�~�]�7��k*�eY'Hy<�g�t�t.��"��=ە+]����-���r] �	������Kn�8@٣0���Q�������E`�lc�P(yS�nRӊ�뷙�5��;%WW6sm��\�cL���.&�7�w:�r&��f��Gk�=�%ҧ�x�6����c�*G�m@���4��3��s��}�'��B=�J��M�Qm�k2;J�7���M۾O�������Йoe�gFҚ)��H1A�@�l��Ű_Į���+�T$�PB��*J��v�ӊծ���1������N�L^gN�V9��95�:_���:��ܫ�:m@Q/h�f���ظD[�����|һy�s�7+ i����QA���:�V<��xm�I�|t�M���#�g%Ţn�Q-{saSz�h��"v<�O2�*
�ܠ:7�wp�����bӭ)��Bkd5p��Py؁�d_:Ho��u�7��������'�PwR�wr�l��m�����s#����w�K��}ڲ�j8X8��q��Ӽ���.%�ܮ�f;֜�&	c,l�@J(*5��)ό���t:�r��j�{�œn��X3N����;">&u��{�Y�ھ���z3�[��t�:L��Ħ
6�b+��L��mr��W|�F�B��]��\���rTc+V�E��\�iQ�+E[HӚ�M��櫡����m�"c�ܒ<�P��y^�2�*�8�*kge�z�Z��ǲc��x����䂘8gH��]W�q�6� 5�gl�٩��
��Ufu������yJ�Wo'Th��e�d�dl�S:�J�23Փ�VP��N�%����&zl|:t���-��s�nٓ��)-�&	E]��*�<����ܘ'
�t��6Vۍr+$٬����� ]ui��ܣ�8C��6]�iE�V���
����*�W�ЇL<^��~{��}�����2�HH~�$�	&k������x���옧Vk K�D�_�$8X���Y�"�b�dͽݼ��c���t��2T��ć_Y2e�9H�f����		"�\�3vL��4�S%�BM��uC;y&��n#dL�ދ�v���K��-�jںn!�.E�1�Δ`A*���{;^�K��z�1i�����&�����Ǧ��>��c��G�K�8Q��x� �nL�*��@N�������Y��iyʏ��{����^��v�;��v��^���2B2��$>�y�y�⦭gRל�nJ�U^�+w�'��l,xfY������6b�g�F��ͳ�evU��,��[�{n��.C5A���a��4]과JC[B��֧V�E���٭�@�Fa�4`-tv��o��JG4���f84�٧�\��!$Rd�t4���n��j`������;�����{NwMC�(�sOnH�w�f�v�Śj"����m��^�v���m���(E��P=8��j-��P�))Y�F�6$5]�=�D0�ڱ֔K6���R�v7�E7.Թ ��uݛ֓�WȞ�(35\[ƕ�֪�b��eL��#��WFV,�c3a�q��W�{�]�P����9#�ը�PMWdr�ƾ������B�@���CfN���9j�P�^,��9T��v��ü.���Y԰�����Z
�Mf��T��}�#cI�Hj�6˼K�I���|Q���¢�q�_\M3��Y���1{�}�)5C����H��{�\�nhomj7X[zY|�u�[�[G�[���i����hjx�V�E�	l޼�`'f�.��4�$��S�Q�3��̘~� ά��U��r�]�)ج�F7lt i5�4�y�%"X�6��@]dA7N��/]�r����8��M�Ҩ*�
�cl���	�F��䂾p�I��,�F[�7�V���Ѹέ�\�|9�Z7�y�6v�����
�nR��	kw�\7U�\ 0kZ����ݽ[��AE2'��X~j��VXW���MG6������b*D�*�k�w0(�j��Wȼ+��o;��s��q�nc����|�nZ����S��>I[ꔰ�y���Er�4z�	�$ ��N��G;8���%X�a�V�����6��e�}����V�35�rW+�HH�AA�Wnf��OlˎkGm�;�n�8�nf�����a�^��w��9D���(��(�r-J�������x���L�2��[���"ڌ���VV<�CiF;���L����I�9�4��]��w����p�`��T8��j��i*k�c��Q�A�J̇_,Fk�|DA�qP���V}�v(����+��İw�Y�>^�t7�b���h��v[�g�ǲ�)�v��ݽ���ڙ�l涕Ʈ�-7P�����[-&�i�ܫ:W�3���V 3wW�����yow5Z)�Ȭ��{WFT7��XU,�i�d�����Y�1Yo�(�����W��ی��wX]Mƙ�mNrb�NB,�+���g@�.]K��
����HV���evͧ ��E���s��"�A`L}�C_t���V���Ǽ��i�����R5�.��� j4�&�q�Ҫ�tX�������7�Zf��]P"�n;���]oS��P][�ômN����4��7 ��8,�wE�.X��SϪ�K[1��p� pD�$J[�QϞ�Ҽ ��32���XV�㘓�E�#ː��;��t��k����mcu����ӭ$:�VA�X46�<c_,Zp]s!�C�e�K�ft�q��?���q`�ȵ �s8�PB��ֱL��nh���"�sin�(�|o��9'7�� �9'u:�X�;�Y����*�8��,Q[�Z�����ӥ*.�Z�+Q�F�p�im�Y������l�ݷgkV%Wt���`D�����A��+pS��bƹ�I�A+�
�M6��{�h���
��*9�2Y�]��+n��Бh8,�E�1���i�P�W'}*��7ՀMQZ�,�$'�l%���;z��[���ra]�H�L�=��hB�� �����5�f���ט�ѓ�ރ�ם53�w�ѭ��^vlS�p435Ӏ�
��?,�/:�R���J�]˹�!=�iVe�,�d�{��J�d%��D�����B*6����X��b`���2�ҶMK�r�y#��נ����#���@�q�4p�u���3zh�H�W��\����#�j�@���U��@�����6r�-͜�9A˦�2��
���U�h*.LY6�yC�!��nh�v^�:�n��gvT�Y�bb�9��[X
��0f��0nS�j��F&��i�wviL�W���{|��m�OuT�X�u�Ժcv���\�L��I���2[w:ʕ9M��ϫ	ujjb���0i��1�V٣��/luG�kd�6Vo�5�r&�^]s����$�S�v�.�,x���\��U͐#J7t��,9�(#C��`�ؕpy��!j�|��6�Ə�w��a�V6�����Od���69F+lp��r��
���V9�UuEi,��[+�]l�3�U��:+��7�3f9V~�h�'NB��ce��//�\8��������2󢊞����+��D�\�*ۙ�vXPX���ә�FzF��;6w�s�r������[VK�Ӻ�t����}����]���|h����1�H�]׽܈9Eb�jf��#����4(
X������D+G�z�e��|x\	��i����K%�,X�;n�H�[γLn�����/h�g�
����9
=S#�9�u`ϓ���EuƯX��|�R��}�V2Ѥ����g�ȫ��J��`��a�>g5���:���v���
!7t��2�e�z�)Ԇt��: 6���H�2��/NU�ٸ��H4��L�:7[E��Y�D������"��W���c�,�ζ���0`��E�7���ْN���OI�����.�&r��h�������ua�߆��R�n�*�헑D�O�V���xMKR�˵9��,�_\Qf��*�L�{Cr�@��tvV��F�n�?��A�F�kmh�X���.)Ղ^P
$�*����B�Y�j��&�3p,U��|���V���3\�T9c��C�:�˹tkS�	�"�>rN��:ws���u*M�KXfV���I��$�,@P�T��ьn\�x�@]���$��ѵ��h�p�������v�Գv\w�n�rَ�{M�&Y����h勺8�,���rU���tF�X�s�x����]�8�.�Ds)����ұ���:�*��Q��+�{e��Q�?ofm���M2h<9u�[\�]�6��2nc��-a�� ���͘J�!,Sٮ�s��L�)t����;�^'l[x.�0pO�� ݫ�ۂ�sB��"�����;��ԹG���u��50#�S� �\�����M:�����D�A��wY%Z`ƅ;(j����ou>�!��8�<B��n��:�ϱ���O�S/-�����EЕ�����'
��_@����Rl��^������a�sZH��)�dAǳo|q�;Y��z�.��F�Υ&=�|WP�&�0(]���!Z�/���A�̂�k}Y���`k)E��;�$��u��7Z�kEL.�>���ve2����>o���(S+쭭�{���Z�5�,��$v:4�� �УRኢ/�"�#@:��gros4p��ς)V�% ����RLa��ºƱ�M`�g����bR��n�g5�����X�3k��շ�r���d��62��&��v�o���$����TOd�f�k(�G���y�v�\��>s+��{pݱ� nÙM����R��c*�IcP���C��'m�� ��u<�m��xbZ�-,ӉeO��]] U˽v���]�JO�Tr�;j����ᫎFr�H@с�c�mk�}�l{�f�2�ա(Z�#�������WJ�4nW9�Z�|qr8S�z1� �j�*��g���pq<���n���᳖�f2�-V�yxY���VN��cS'f���O�`�����onRѯ)r�N�2�#�U�)s ��	�*��IkoUk�p4������ ���9so�n�عg�`��W�mhkM9)�/X��3x[-�@�np�2��A�D��8N1u�WB�D��ѻ;��˷W�2e<G���Ơ�-i&��pDU�5ҝ�e��V�9ɻ���.3�Om��t������v�8��u���M�-K�0�Ą��9�����%�]�wZs�|H�um ��_2�P[��k�Y:^���\..j���7��ԧc���;��
�H#�ֲ��XV���Ŷ�M�����j�j
��rw"�	s*����4*<�G�ђ;{�5��(w2�h���s�EC�8�3]K�Z��
�t-�&�������
�G9*v���d�����=�d��Sb'��]1Jm;�o7;6����!tXwt��n������O\6Ě�{2f
Z����9��\s�J�D�m�o��fB��%�>љ�`Ibו)/D�!w��gp�X��{����y1#�V�&{U��^�`ʼV���E�K�[����&��YP%��\�}�v�rv��x6�$kܫ��ř���莹��t�ww�R��u�*M5[�u���Rjʧ@���t��w��uv�Sp\x� [fHs��Yl�PL6ڌb�f5gNl���Di�E%�t����x�����z��E�s{xn��Z�s��O�[��l.��2�E��*%�/�t.r�\��;6��LZ�%r�[7�4��`oWz�K���.�#&Ga�6�L��wu�6�!]X��fg[��m	��9{u�� 4m�����5lD]a�ՃqR�/`�,�K/�^)QZ�=�����ݾ��e؆'BROy�D����!,0��QK�Tnj��n�u����!&>�.�v�Г�M�����Z���neئ%������b!�A�8�ΤՌ2N�!GM#{)�ɂqǲ�*"�i˗bl99a&&[ɐ_nվYC��d�v�,n��Jed��K�ҝ�!]�n�=Zn�S��m�E�SBc��6�ZJ�@�iyܺ�v'��T�Fa*�v��i�7�S���t���62Ȉo8et�u'�)ZG]_�|]Aa݋�ҝq�7Y-NsԿ��{7�R��Z��u����Nhq���LN�1���Q�]1U�Y*C݌<�@��p_i�_z4Q\�a����h���.�4bJ��ܡ�����W-7z�+���q��-|��l���V�Ģ�ě��������Q|��,&]��S�S]��pf� �j��n�R��j�)�i_31��3�����FA�HU8w1���5�^b�']b����q�:��hn��Bq�:5�� �l�5�b}�Oh�䴉�[֓Ψ�t�]�H�P����A2;M��e�ӌ�,����i�Ap�b5��wpq�&�.��1�wh=�u�Ŗ��;z��՘9�I\���{qֹ�N�b�[�k�ŕ5��`v	�%��Ҭ��O�irbgJ��Dl�Y;]�Y�w,��!��aZ��_�;�j�Em���^4�.�o�ՖzD+�J�E:���Z�����a��L�k��\�'�Ɠ���yOMtL��=K4�/bzx�����{�{���m��9��sE駛o�e�֜��Uh{�'/����+d<��k����iCD�0I$�f������%K�)��(4�����w���j���}2����2�V�F0��Σ�U���!���r#��wW%X�)���t�)��,��2��ͮ4��2Puk�����: *j���V�k��Q�\b�����B�uz���T�5���P�r�Siw��/UUj��'Ο,��o<J���吭���F+՝eE+s�P�Қ|�˗�0�N����wa�J>Ty�3(M8�f��閩O�c/f�ei֣�gbNf�V�O�cs�q��a�+���[����Jz���=�����戵�d���m��i��w&���c�(ᨭ����*�ف��a�'m�m�`�ܩC��oLȰ0�Is�,�f��V[�*u^h�V�z��G��Cy�d�͵
w2:���K�@��M��G���W��f�-XI@
:;�i���;eJ���sx��8�n�vH�e�5�o��-�����ĻT��{��=gM�[܎�%j"V��+Z���N���OZ�7��#H	��l�Y۰gO�x6޿�ə�eI9����&���}��\�Κ�pn�t�Rpt��by��у�� ̫�G4��U9���3w`�\
���_r�I�x�;�AԖ-��Z�!��q��"à���7��]\��70s��ӧD4N�rV\�K �k�X��꧑���)wL���8^Zڃ�-6m�[l�]�Qܬͮz�w��7ǆ3\����]+{r�n�҆����9-'S��n5v:�d�_|�ƙS�����E����M��9�7!3���r�����T���* ����ڳ�{;�0o�DQ<��N��\DK�v��l�;)�W��sT�׼/(-gS�Z a�ڸg&��sdH���k��r�ư��ŕ:lvNs�y(�a����j��E�"���#pe��yn�4���:�f<�����o:��>߶
N� ]�[I1���Ǝ�t�WSB�{��%�,ӎ�DV������Y�UM�Z�X;�ۧ�t�KMՙ1�b���k�5��̃:�ѻ���Um2�Q��}���ǵ���%���(�ѡ�k� }���>��<Y�3<�A�[��7Hy��܊#�Xܜ5�]ɬ��XV2�:�:[��+eK�{�8�1�����7���IK�6�]ūr�ԅ�|e���ҏ#{X�U3.�1��^\��uaT��m17:�g&�ͼF�Bn�D	y��{���cv�:����MM�#>2���JCk���M����e�N0w�Tǖu���[!��FK��Zn�_[i%"�K����Q�,Ԃ������ս6A)�����l����-�3��5�r�D�'��ņ����*@竬Y�HG+>tn��}ɘ�����
��[{���=z�p�5�_r���$�����m+qi�7��#��=Q�n�P(r�U|� 1�4�����ӭ��0��2���^U�5���G���E�HA�;sT��&D���s<m������� �s��)�)F�L�˖n�r�%��V}�z{�t*d�0��8��p�SU�8&�8{L:ec}���i�3{�J+�c��*��gObb��[Hn�]	w���nS|1b�\�A>�����s�)����,�U��\W�9��u:K����{�jdt)�G/^�k�4*5r��_�ت^�-\qE�r�H'XwU��r'�oY�FVF�w�K�WhxiqvR��sw��䂯��R���� eN���NVzZ��R(˹��{��*e*�Ԉ�i��75�
�9��E"�j؋�n%X(���b�(�*1b�V�Z+X��,[e�e���S��F&R��T\J0#�QDVMZ"��2�uj:�(֬�Ŋ�-1�i,X�R�*�"��&�PuA�����E�Eb-d�(�h���Ee�r�0J��KlH��e�չb��U�UX�*��Q\����f:��EFE�ZʗM"8�!it�k*�1J.U-��X�R�.!�Pr��EU@Ut��6�U%��]5DFZ��1�Uek���IiV
����(2�+EJ��T@�֊�Qu�I�r�T�A���VD*��9j���U�*(��h崲�+A �j�Aֲ���+Tb�2�h�Mat�LeQJ�ARԱQ4�Ur�
�J,�gd�l.6�w֧'�X�f�|{0��P�,X;%Ň/�}���u-�dGnQ�eh������ŭ�A=p��;�+�Y�9�{�R��v�+O�M��8����ҡ��5p>�K��N��x\7�\�k�ڼ��]���)��3hJ�{_ҡ�����Ʈp��G<���	׌x=��ᱤ*����]Ds�[�bV#��_�:efW�mR�)"�}lHp�D0�2Ib&�׮3��}գ�r���	 o׸"s>�[���Ǝ\׺U��i�E�x���]:�q�f{gw��\�Ƈz3�\��K�����efg���3��Gzʏ�1-�:xw7g�阮��΂����{���
N�G�S�
�wL�k�uv��Kz�"�^z@V~�9{h~N�OK H�����;��=X�7:��1�e���Ӟy�!8�U���4��qA�J]�Xc&R��Q�����������	ᩋz��w�;]:S�*�)�q����
�g��	tt7SGВ��䑇�HQ��1�3.zܫ����edz2�o�V��8�(oE@�U�P�eQ�>����/�"��Ҿ�V���l�'ux��I�Ev�ȟ�z�㱣�ݛS�^��&I�dI�*x��x�z�#33��W�`L8/!)�Z9��ً�1/[��jٕ��>�&�=x$�ãzSړ�K�;IV��r�����p1���uh�޻�fS���]���i{�%|�dN�����6Ա{�z���U���/�
-�\�x�S�Һ���]W��ˣ�m��+iG/R�+��xt��AB��I;�D��㜔ӟt@l���^���ۿvgK��Z���)�`O_�ߣ�I_ӗ��G�OcM�-,_p6.y�S7�eS����;c���X�����Ps��X.���Ud�|�؝�R�.|]�q��P����J��/O>��X�]D()��c�������L�Ϧ�zt{瞽E�|7*�S��XN��׵��{�rY)��gB�n�]	F��J�6�|��7�p�bdp�8#�I5�0�s��\ΝJ�V�y��r[yZ&L�G��r&��T�N���T��c�Y�<̽7�o�0]��>x���*t6�s��LW���-����A�/��U�o)��4M����Y�dI��F��r�zw�b^�e �Jc�`-ް�/>ՍV.��ƨ����^���pݬ9W��&&��Ώ<�+ �J^FI#��:�XճV2�Ku���)�%�z��o��˼�\�WI��H�9ϣ;�)�ٽ���ʕ�.�x,�iի�I�p'tW%1���&�i��ͥ�g-���z2chm�;��ћl�f���huH��76H@z��t;���Kwk^N����ˊ��#��K@sV߶j�Ρ�ߖ����o��nR�]3!�*/pQ2X��=��5*k�F��;<��
����p{�G:+� o��cYS�a)k|�EW�`j!) 㾣��Ҵ9�nNtݓ���5B(���c
��D�={E�{���LK���޵2^�}V�=�	�6�Q�(�;��"����b��k�i��	ct�}�kP�m@��/�����8�ŭf�$�}�2�޴�6}D�g֔�aZ�)��Vj��=�LZ���7��t�]��&� >n���"��~E]G~5�Z:�5Y�%0׆Uq�=�+`���&W-��rr�=�z�|H����=I�u1�	3Ҭ��O<5I�Z0OXw%_�F#��e4�{��=R�zœ�X����vW��a�u�ʷ�xlr�uQ�����h�rxa9˝%�x��q���c>���^���Z%��kU��=�� �:t���_w�]����3"//;�@�m�+�ӝng�|i��asۀx�@�q����,�bo��jf����F�!�=)t�������e(��c����p�&�����?#K�X�g2.�{��������ܜwZG��+1zշ�k�g}�L��[�f���6�$nIñM���g8�I�sK�b���'k�;��O1ww ʦkc��i�\YӘ-j�N�hݱYs�f���W\�$*�o�5���V�W�~m�^td��QY9�sg���t����p���gb��3�k]�)1ɱ�X55[�1_�Aal������t���g$�x�,�p��/�6�[�ˮ������-ݰ,j�=�j��~��P��ju���-p��y��>u���RJӾP�5��[��G�����Q�e_�����d��r�M�;8"^�)���Ϩ��b�.�������ܯ�kq�CQ+2]Ǜ������V����@���PV�T��(�o��p���{iP��wƌٍ�2�'�];�^��y���5+�05�buZR`���nsgii�������xM:b�;]�{�~��&�h���K3Ő�@�䫄/,D�k�X:�N��Uzm[���Gw�3ݙ��!繽�P宻�F
�OQ`�T��������0��:���K������<�T���ӂ2�[�}U
�]�����R��f�{�xQ�"pxV�FѽV�y?��ζ"�.����{w�X��*�0$Iء�S�s�I�/%��:=�SA����:.e^HL�Kc�B���s���-�R@u3�P'a�{WG��ϏX�/��$���%������l0U<�ݼ1ԆH�Mŋ��VN;�N�,=K#���cu+�ʗ�^�M���];ְ��đ�MG���d�x�'���[��������U�����c[�X=�E��_����u�Ne9��9��_���])N^����Y_�ׅ;ٚP�'�U��^S�����N7��6�:Y^�/����t5\bt�|�f���WS��Q.��\w�9BvmӠ���"����2e��^+=�4�c)�b�93�&��;je�|3a���[���ť%��۽;!��XJW�,>|�OK�S0H])����/�UI.q��쀃p��P�x�9e��7�w���?Z�6tW��X���Ug<�ʯ&ڥ�$N���=
�^�a:r�L���k�vV��m����'��g���0�4���9�80��%�殞WXkG�5W
��{]�S�����V͙N!C�*�oБǔ��ix@�<�^��������V��)Aoc��f��1�4`��i�;���{�e0|������qѱ��c�X.D� ;C�	}\D�e�hԍDjE��=��"�+���S��ǀVX���|mZ�5��"��2���J�41�W��9Ndf;�R�����b=k��֤Pƴu(m�
Q����C��y�][(�At�,ݑ5D�9�ֳb�1����5���x
�Y���R�<��C���J�#���%bD�A���u���.5ܷk��Eis��-�[�5Z�O�ૡ��J]��#�"���;w6϶^�j��λ�'�Rw3�-�� yY�ZI��a�1(��sމ�aD}	���"y" z�{ů#�q�����U��S����z2�l;�h��YB���R�({y0��K�@���ݧ�NHfog�Х��]J
�ў��3����V)�=��75_���F}�E5 !}���Z���$�{��ʻ����T�uT�<l���;򂅖G4��c�c]�L��" nr��;;�7�P�N����x�74/Tw�+�ˁMe<hOcM�e����g4���w{=e�;e�9�Z�d*i�v��g%MUa�x����PϣvQ�B�y�[�;V���zД�B�\]Bi���aϫ�ga�8 ��t�	����S�^��P��v��XV�w�[K!�8����Wd���]���U��{+�M����7�<fJ�a�K��J뛓�e�Y�m^S�S��Mp.q蚹�=��N��ޫ��Wk<Gp��L-�+z�u�+����Cy����eueyG�6W<��\�M&���>	�\e��'oe>��J�T��vT�M���;y��.�fu��?]��BoF��w��շ~IN\�{n/�[y�z��J�� ;���zE���0s``,��=Wczt�������<`�Q$�/1��{��	t�*�fGH�ᒃ␡��b�%�fe<6�}7g�o^���`���޶;�-%��Et��txj~.��p�10f��c��&c�!頽�Ek9>����x�P�m��Җ�3�K 
w�*�	;(g�Z�vg{�5��챎M��Հ�X�|��E�^"όko�lUץ�BZ%E낉��&Mrv��2�Q����N�5��|����7=^�����+�hx�R������<�`SQ~��rx�̬����|�i����>`�x�,�)��a_)`e���yi=C²�2�ώ����9c��Ȝ�����F)��&��=H�{�W��c���`�)��ĩ�SszN�އ���gF���5��^ı5���n�v|L�ᔵAV�SÔoZ����x��{�[�G������
}0	ƍ�9b+���RU���id�koh��P�(/y�� �~�C�����iK�Vz�y�H[�+/e�9K���uFj85*��;��v�v;�%P4mX�F��wٛ�e���z��Ͷ�Q�+R��>�&��r�al������wL�ciz�[�P��U�l�S���r`�ZN�g%�"/{&�W��W��ə����?�۩7��(y����N��G'_�F�o���P���#U�Bj��?ow�����y,�â��S�S�X>�>e2���g�S0n�2�U��Ŋ�O�~.���8����B��7�/Fq�Ť��P^U�]rZ�g$�*����t�x'^7ޘ3鏫� l��}��]oޓi��oo]��~@G�� U���l<Ke�%�����f��j^t�O!�v����&�o������`����FVB���/�X�:�*�e����so�,v�V7���l`�-��S�6ͱ�W���r��*5k�D1:�ynk�r 7��%zԭ�Xg7x3�HW�ї5plz��x,+ҡ�%�����J7Z��M>ݫ��J)�c*�@Uά��+���ڒV��;��`tۿ,�u(�dL�n�Őd��G_�;}�]cfɟY�?L;@�gr�`��eh��e{��MY��b����h�{����<ݶ9�i�8}�
/P�q+V�
4���6���[�b���r.P+�U[�Ѭ~����}P.���ںڽ({K'0�Ч���ˉ]��J�����Y]�湌Xf�� %�(�q�g��<���QnÐl��0�t6k�jv�}�)g3�O�Ջ���~��=%?z7�����c>�v�ɷ2@L�{C8je��S2�)2;{o�TA�w.ƿt�V$�JL����W:ٺZf�/���<��Jg�ǯ}��J��q��w��Kt��]>�`�.���0���Ƀ"�%bVz:}Iw�]S��£U����/D=����WnPc`��L�K������h���L/6T^�T��<��_%o�/o5�zh=N�o�+9�Pj�9�I��_@o�ɢ�lu�ؔ0�(N��������<�oq�V�`�.Kz�myA����T�ke��p�.�1x���dw�{��:U��#�мCN�ϟ����ԸA�*�z,�Pk�3w6�]GK�ٻ#�ײ�����ۥ�%�Jw"ߙ�
*w�4�<O�m���`Ϛ]��+�	Ih�^�;�WQ�ً��n^�>��5��oQ�y)ǁX��\)[^M�7C�k�@�Vxs�ɹ��^�x�|D�5��`����L�Ϧ��}�	o|�,��Zr�o��[�"�xl��O}�o�������u�C�t)�%������RK�o�\�,S;�p�jhs�K) =�w���f
 v�r�u�X��v��7tr4]fQ`��rnl�g,@Xyx�e���>}Q��o��/}�OJ}+���;�䜥�{3���p6{Y��͙N�x��S�m.��A::�1�I���v�kP�ˇ6IՀ���n�zR8��n]��)bP�9gL��&ڥ�$O�}lHp��C	�ϝb*:)��s���g�2z����K��#�X�b�#y[���,�ƴt�6�ݦD������+Es�E���Ϣ��q]	yM=ixA�f��X��`�x�4���ݔu�o@.����=H�>7 �bb�{�e0|����sVG�^������~���i��N�����V�Nf@�)�I`	��c�1t�-�T�Jv;��^��=�t`k��u�Ǟ��L����3�*��E��ɔ�R��u��>M����L5��zF9d�{�?&�j�����N���bZ�%����LK
Rȕ�\��N���1h�׻ӏ'i�G� ����q��]�ʼZ��Z#��P���P��n��c�칹�r:�A�o9��1���M������{T��DuYXe�o׎Ҭ����w�y����={��_�O��2��C쥟Gz���͕:�xt�PP��ҷ�tO]�$|�W;�����zr�sjo:9�2>�F�S�e.���#M�g��6G���X�t�0�CoR��ao���v�K�ȨC�u�u]�'�v ؾ�����n�Ր�/�]����w.�^\2�z��������4�9�K�� /yq&���i�Ň�f�J�4�q w{���VIB�� �.n�����k��9y���f���fq=��-�j�|�"\���UbK��o�0�O���3LEZ!v��#x^�o�L�ᴘ����:���S�`y�T3���_I��ꙝ�\�9��XM(wnK�t@��[3fIJ�)&�B�_����n�m^�����Ό��'	\���n�a�Zka�r��Y3��9��K��Kp�X��ͽ�c嗉����@���.�[Wv��ƌ9���δ�p�@�Ź�iu�Y��m�b�2�=�L��&ު )�swm�O��$��ЫԵ�Mؗ���U�1���|Т���쾔�3�م��Z��f�wG�%���E��z��}��U����S�^c�1�{ P��L�Ϻ�f�ա�t"+�W�\Z�+K1&� {���d�X�kR8뱾/����Oz��}����k�鞤�P�gS�<���Cּ}��2EzzF�H&�uĺ�{*��n�m�X���f^r�w��"sL��d
�v1N=1��
H��diTk��/6��R�n0�{jm�W��p�6�;j�rO���uң�RJh��U��IM>�ڗ ��\,�ݵ�uu��n o��tn¸�u#9��w.JK�3��=��S�<�|�:���A��eK3�h��>r�Wu���O�GWi�\L����N�rߘ�g{{X<,����h[��}5ڤ�I����8��]�S%N��\w-�C�/�]���w�V(��J�P���A��nj�+�`<B�;�@|&�%�g�e���]�����,{Wr3+߅�Z9��\[��iՔn��c��&	cC�W�-x�:�2�\C:K׮`d�*�a˝'7V�ՠ��Z��c�fT"=����K�xt\p]ھ�JOy·��T}VEYr�Iv7�1�go�e���WOl���p���WWO&�f^ft���������y�/h���]Z��K�q���w�f4fG�{�L��>���-	�)��]�$J���	��ۿ�C�v��.�/�]Z��3|�.x��-�)*Gh�W�$'o��.��r(;�S�V��T�*w^͇��̵� �Z�<.ŝ|�����
�f��������4Md�u���F"���Vi����"�@cLฮ�̹���܈J�s�(�۲G��o�������tKim�ψ�|]f�_s�Ѽ��	���8GE��j����b>ý]��僆-oi:^����yN�V����ݮYF^hz�68��ml�v̂p|�904v����2�;����\�C =���eȠwsN�R߶�u	�A8s*���Z�Yr�Z�`���d��p\�*5
1��[U��DFBԥ�+Z5h���Jԭjօ*���Z����E�E��
�F���-�j�6V4hQ
��91�+V���-�+bV��(��Zڈ�5�UX-��lQe-�T���YDr6,mk[R�Ũ[m-V�֩D��-�c0e���ij��ֵ��ڨ�D)KV�TE�sm�J�2�ml*5M7I���Qlmm@AF�Z�J��Z��[F�Z�l��[��m���X��n*[��m*��Ȗ��-b���LEp���X�e��W.e�mR�������#�\��ZԪU�֖������\���ŵQ��)V����PU��mn4��(�a\bR�s;�5�s��Tf�l��^��"�v8� oy�n��ά sE:�*������w�M��^�l�hZ��M���ʶ��HR��x��@o_�/����[9�U8����p�cM�R����5u�r�pi�������O���������9(9��=׺W���F죖"���̩��B�xL�=+�-������P_���z�qL�>�gk��Y����+^�l���'��"�/w�GV�ⱱ�p�T�x`X@��&��,�ة_&���	���x[��_v�[�����#��`E�gg�7L��+um�K2�v�ύFտ�,�y��f%ٮ�9�e�r�P�{tǦ(I�z��ʣ�����	;-/�U���1��0l�9�՜XsJ��C..�c�Җ��ʘ���@n�G���2����.�2WF{c��)Z���bUq�ϲ��=9�!�q�sҖ�= S�U�*vP�����E��;�F��5��2tWXpKQ挣�
��f�nR�]3!��VJ@I�5�x�X�}���Wk	��g*�Zq��꿱����^�CĘ֏u��ʔ�!¹=W�{�؃g/Vv�U�M=Ǉ(�ڸ�ٕ�#��h[T�v&f�ds�ȁ�bsd��[:a����li�MWS�SX���0:�nӀ�4#���h=4�F��YP�z:�Ӳ��$�4W;��;�R�΅��l�kIw��͑��e��8��ۭ���ׅ�΅�)
8����Q;�^�E�JԽ`�G���ȶOgE;�%KG�ed�<�G)L��I��Ћ�lZ50�:�&�b#\@gaY�$G��~������%H��y�as�e�bs�Uu�eN����Jr��Z��V���[�'Y-l�Ir��$�F�ѽ��� ���h�U�!Q�5�-�%;�ngۮ�!^Yކ
኷n�-LO��	�ƨ
4=�t� N��G�o������>�o��;W����:[��V��;������<���������2�WT�3��t��[����8�+�Ӭ��q����8�|K�:��䵪����	�,��SF�Y�-�\ʑ���F��$�{<v->!��1��7�>o���&u��Y]/�l[�B̃���7���#/��z)x;�JCL_��w�������
�>+�ded1���`�\��}���nz=<�15�������x���\,:��\�,.)�MV��~g�e��>TU:u54@|�y�yxu��ú�|S����%u�+�Ú��]��v�)�q\6�L�³h�����Wzs+l0%��k:�ꋇuǷ�����SH�3~��Pn�{�;M��M��i:��z^ v���s!�\e#�^ދę�^����hz�
g�+�����/�7Nu�=�g��( $Ɠ�~�}��+�����rh����ܩw�g֖s^�Ã���Vi�V�}P���a?�mߖ�8�[�y�Z��~ޙ��31:�s$X��8��+�>c;��/��i�2�ꦺj�D����2�����}i���NhWȱ^顨��A��<�D��Z�AY�A���8Z�{���6��Y��s.o@U�#�9��M[5�^U�r�XL���&ζlR�5P?Oh���o�^�z���s����2�(`PK���wPayb$x�[]�K�Gu}Itԭ:�q�)��d���Nī*�1S�m}v�&D���C��⢱�����e�,e�c�;ͥ|�.��ְ��aޫ����Qӏ�&׶����uI�C�ɢ�펵�F�>|�~y��t:�[� P�%.�_��P���� �`���'5�Uv�f��'�/����
�6�7�������U���}��k~0�B�?e�c��zP�X�� Y�g+f��o�[�{����(���Af�ݣ�8�
5w�:�m���]%5*m�W�͍(�� x�\OG�h���Si�i�#�ٔrV"�<�8�Zeڬ��ʄI�2ݞv*������Z�-�RS��ͅw���u�y�5d��u!����M������\�T���4X��OeެMKo__eO(Dm�}��p������a����Кz�K�ʛ;��~>�?r�V+�\):��=7L�	����'�5���N��z���Y�E���( ϚV �W�L�ɮgڙ{�E��i�7��В<��}¹қ�ҫ80�V/�>�>��c=���_T2,S/��.$���e�Aʩp�+L���y���[<��8mԶ�At�	�w��VeW�mR�)"ʗ���Ъ�w9���|�ͯN�׍�%��jJ�I�9G �˼xe����/���C����%��j��a�ߟp�4���X�H�n[�$�zǈ��1�+�:�=�%1ʽ>\���i`�X��S��La����Z��[^.z�-��t�hإ�xؐP1;�A��@�o�N�ly�X³<4>�q{5�{SVug�N�.��4�5�y؁r� ,M�%�$Y���c쭉rz�j �ǹ��a9�jvAi��	KK,������G����GӖ��3sՔ���.kN�r}�E�S�����p:	��{�(9�%�[�;jt�IV�j��_o�h��r���	�S�IY��9:�)m�}lMǎ��V��J-���3ۄ�>��bm*���̣��.���qE��'����|�of�Ǖ�Vj'���F�LKQ<{�1F�Kb�7B��o�J#i�G�(�DnS���E�[�����\��E@�\e1J�x�g�0N{�i�2NŦ���"ԶG���^#M��L>��ާ���ލ�2ĭi������FJ�U}��	c�X���S<l��x4Y�*��FM��u<ap�/7;��y���SKdN�h|Sɀ\ssB���S�O���G��G�˥Rp\ʿ��ꕋn���з�[8����"�P���Ŗ;#�U�H�ʍ��b�}M*��,�)��bn��mh�:����tzh��z�}�3���v}:g��Sg*�P��{�=H�i�ު�>�x����g� +��2�]jlT���&�M�����2�F� Є�s_�ӑ�$�-c;���U��Q2f���Ս�
��&��%�-��%��T����R���c�	uLq�R��i�6�{�m&��-���Gu�mu�k�-/]�͙�>ܻZ3fY�t��rJ�G�5s7(��ʏ�s��m'��|$Z��c�敭]�*=��8=�ȶM��m1%��}����s�0�;�ѧ�N��W`a��S5f]A^cثl:�����@�kc������eyk3(��ßEی{�-%�yS�t�]הs�>}�A��8�ټ<�������WJg�9e�i�W�:�ٞO�@�)�2X S��Wy{�^ן
K�IKf�]�V����걊�b�^��g|��}{b��qx���X¹�ߦ���i�w��X14��+|tc����'y챠�m%-?���mp�z��f��&jvny��!ԑ��'��B(���c
�K(������������AVX�hj����%.�S�n�9��h���MY2yc���l_�װ�`�x�L@S�,�8��7�9i���>~P�m@Ϯ���u�e��%���c�7V8	��P|�s۹�/����oP5Z75hc��{�V� 
}0�ʎ9b+�G~5䖎�z��C���y���.���K�(iϭv'���H�OT�09�4��	�`�9`H�+�i�dw��5m��GgЦ	Kt�0a>��/-�x<��|����r������A�4�� { 隸�3]z��F�.�H�JOrޣKޗ��5�R
�/�a���P��Na�ܓ�)$�q�����6í��.͘�#�v
�����gsǌȜ��ԃx]�����	��i>�i<z�G;7p�oҹ�p	l��WEZM��!{*���y2�g\ZKϵ@yV�u�kU��آ���^���5�4wZ��^�s��~��)o��u�zM���-�nx���~V)���h̞��{��q�u�e4�=���|�4�$�h���B�.#q\����{�,��|��,��6�[�	J��0O�c�.�o��W����Kc(G�~��	p�0U�QV�h+���S_o�y�e�g��aPߜ��++��˜���w���R�^( $�G�`���y�1-��	C�p�5JyVZY�z���MػڒV��;����Gۍ��e�zܗm��ٜ��CT�3J���#�ł]R}��s�X��'W�CŦP}�^�ؙ�2AG��ٚk��Y���A��L�'�/k\!�n�c#��
��@�6��r����Uڵ�eρ���ce(��v�XL�����ζQ�1ha}<�V ko��s�Ui;<����!z�
�ׁ���b[V�仨0��<P-�M�cњݿp���@����sN1���&[}��y�n��aD��{O[ q܆��[�|�B�a|�H���Ф�o�S��`��Y趙�]z㏎kS�|��1�r��f�fޣ���2�߳o��Mc�z����D��z�j�^��p���bի�г�\��<�]@���n����@��Wl7B�����=v<��=@��U$�r�n��y/Z�7��K���ųk5i���&5p2�"���h���Q7���7��x�R��N�-i�QIm�UM�}[�"�����ٖ=B���-�n���x��GǞ���9!_�ޚ���7���gǠ^�B#�u`}XV޾3j�aުA�!���y-ǽ M���>e]畃C��K*G�/w"چ�Q�czP����^w��*��+q�gK�V��Ô���>s,N>���2���W=�uN\
��ͅ�{S����U�7���:�V������U��G3���( d����}5���-�D,7��͖�E9��m���2�R�����Ê�"��Lb|�{�/9�*f	�2���|2��8�<X݋�5����wt�k.��� ܧ�b��X�k*���镙^M�K+�H����2=�w9/i��yC�	N!��d�"`Aˡ�<Q?7�v�Yc���:�d�N���{�z���L+��|-�F� c���k'�6@q����ʲ�D̆�ʉ��]�'Y�m�٫ɫS;�)��s)v)���/a�(�r��[�:�>�2��\�n=j*<�L��o-��7L[;��C*v��]ִ�]W{X��&a���é�:1C����^I��V�C����
w<k���KDv
�Eu*��H��i�/2�͎o	�c)k�bQ~���X���}�22��<$�B�"�T8����sKs}��->����(��U�+����*<'Wj��B4_���].�ĬN��,"�$J;Ck��,c��>��.����D��L{C|������3�*ȱv2e't7xP�Ąޛю;��}�!�:�u�W{6� �f�}7XG5LKU���މ��P��K�v���Nz��b����]vCD�P�6��������g)�.xU��س�y)te?w[:V	W�ba?w]j�b��u�g�������)��W���O�NpLOy��o��	[�^��@QUɀUs��'C�U���S �ZO���sJϬ�j_p�Z��@��m�W;p_%�o�f}-��� ��nh^��%uP����:x�H���5M��ʲ5V�:�Ⱦ�v�L➜��A��%d۬O��U`=�MgFL�4�i�Ϋ�񱮛/�:*u��
�(r�� G�y�un[Ke�e�ۖ[d��N�r�xe�?]�T����p�< �:\'HR.S�nvm�H���^j|zT���+�[��q,s�Bv���])��ʷvgB y�;��'&_���}n��yZ��GC���c�j
_�e&�+|��)���oT��v1��Z>}���x�������Fz�|6��k����[+ɀ��yB�4�*\[j���s�X<�6�X�e��ִ0�+��ę\�������ϥ��g�(�6���r%N��W�C�����P���=�J5+���͉tá���T�	7L�ӡ���{%�Ȱ7Xd�:9����������������6V}���.�c�t�u� ���[�aw��������ǅfC�׃^��֚�9�Gb�t�fy>VAZ����H�eMܦ�E>��܎V6,���3�*ٵ��<�xX�����`ʮ3���G��&�y�5��vw�N� �q�@8}Ґ��"�fj,E[���d���c_���\<Lõ}��[���sd���^s��+��!��5���ؙ>�B�ֵ�|���ƽ��{|f�8p�fz��N�un���b����L�^�G�'����ґG�U�[7HLLp�|���j����˃O4�0�vi�y#(�"Yݲ�m���7��2e 7d�۠�!��
�u�n��!��]]֧�i�V���WD,
�U-*K�R��pf�)��s[\�md�Ґk��ja�*�nM�h���j�X	8ݺc\C9�e����W)���;uw4�֘���hR��u��M���@�w&��4u]˅C���اgH���H1���y�u��E��yZ;�tǫ����*���'����v@2D�>nc����B���:�Mu7mu/���J��ܡ�P�q_�ڸUt����`�:o��X�-��ɛo#���~���7��:��ٙ�/�4n8��x�Uʿ��Z�iԓi۩�S�rj��u�;Zd�;y����2]*���Ɩ�;ʒ͘P��ǭ�?��+*LPkV�k�t��
L�pi�SG|qV�Y�t�`vgC|�}y��̇��
9C08uNQuʔA�"��*tںT��a�b�:Re�z���ZG(=���.U���#��1��m��JH=�h��sV�y��En�Ӭ��]�mu��SpG�u����
�*��G4���S�����!0	��bu3F��wY�It:9���I�P���	�J:Eg'ZjR�Ov��UCb㛽����QG"�Q6��]�-��3�)R�y�<4�iu��{�j����<�^+
����&��Mf�ѫ[�S��1,�\��hX坁�E�/�.����<��z��q�y�.�N�6�?N��:fj�8�Dff|����$]��=l
�9���>�p��Ie-����H�C�k|��EW*V�W:��ڞ�{��q���$��L�X��Z��ĝ���γѠ��8��]� ��%���雊�\���Eiύ�3�H	Ļ76=�X��=[n��vK�.�z����Pa�S��I��X�*}���m⚩S�U�*�C����Q�ٜt36��g+�[�6��t�y�|^��#2v��-��y��wv	akV5
8ҕ��J]�N�Ko�ƙQgryx�)v�b([U��Q��g��Bd����n���bC|�M�+q�ɡ+e�
^,ku�x�v�b�F9P��Ccw�e�B�1�5i�Mz��mi�,>�fGx�"�H�ط�����q�V�(��
�T�m�e�$��sGwp;������V��k�e���s}7��p��,�k���ܲnN���n�`
�x5�Ӛ���9�k}WK��)�Pػm�o�Nk��e�����ހbE�(^T��r�n�,_�N��7�'X����R�t�>�z��Э}����S%C�����U+
���Ѷ͛�A>}l�fҷ���1�dÄ])�m�ͮ��{e�s#�܃\�%+�f����w��
�fᶈm�;O�3��ͮ�nu��K+�ЫT9!��wz���M�
��j̷ݏr��I�3c1f���XY'�LQ��Ps��.u�Y�e�b�QkV?[��d�cS--�m�����UFWMALV����M
4milE�8�Eƪ�Z��AfZ9E�Z�ե+)�[j���b���Z��Z���h�U��bV"��D�����	DQ�����QD�kq�b*T���)Z�S0�� ��d-JU(����c�Q��pQ[`�Kem�-J���ŅB�V�J[Q`�**ōV�Tk�f[E4�TAb(�i��E+l��
�Zа�c,U�QTX�*e3�E�m���L�b,���j�Q��s*�%D-Z�Z"WMō������ĭPH���ƍ�h��6���������%EE��Q1���cQdTT\�%��4I���mVUmj��"*[dUV��TX�h�����(�Eƿ}�����}����\�AW4���u㏖ʼ��/�cĺI#���J�L���3���妛�C���LΥ`��_=]~�Ԥ��"t>�Z<�%m5 O����Z��Ӟʫ��*v|���SՅ��{�Z�t��xA���AN��`ա�y�O�L��8I]����
�O<�LNxLiR+O���o6v�Zl8%uױ-�*�̵��֑���Rc�C\�&zU����3�͟aJ�d�*���R��k�;�ﯫ}��@2��Y�,{\j��U��e2�}8�ge��s��5�zN��U҄��L�D,an�u2�g�E�w��4P��V�x�T��\��[�]G�fF�W^�~���+>}"��i�{�nCU�����L�\&�k{�u:��<��w54c��x�!�C4�/��	�Rbꧤ�Wl��J��b�����i�9�����`�ٹY�ܤ`z�]]��<XΌ�2T!1ꇺ�S��Y�t�k�Lp��'��60V�C���@׸5n��n�E�<^��������B��/�7�lOB�Y�G��Y�v�/
龏d��cA%4�
f�d�U'�YV�tV,qn�ީ"���yAW�M�(��K�;�#ҵ{T�C��0�v{ka�ُ[.qKo2�蚲G���u�(�r[C7l�ܐ��4��%H��D�Y��4*o��_F��|�F�3/w�2��'I=��\"�r��Gb#S�=+x6�W����Y}Թ��=�����q��5\�[k��������義�E�A�i�G�g��`*�����Ϻ�`�I�V��:��;@��o�8\��B.�	����%5�!�hj+�%d��O2��%�6�}tj���g+mr>���C܁�KO�m�rӳcD��s��]9������\��*ғ50y5s����jͭZ�?zh'�R�������A}�k'�0��S
V�q�:�F$lByѕ[^���`}��^��Ӽe��wL��^�+�TwZx�����ۥ�D�\I܅@��GC��_��+ޮ��������oe�U����%�Ue�٫�tTcu�OW)}����!-�S£'�c�}%�^��Ց"�)}Y�J���oUž�*kve���06�	��ڦ��ԧ���kQa�3�<����N�H�C���/�G��S8�m�5.<��3w��+�oG
N�ǩ��(�?L�A�ۥ��J�v�����W�%�� �oG�i;D���FW�`�>,2y���ޙ�bq��~5�z�L�N<
�	�I�WzS~׼�/F�ZSM��� �7�O9����kqP�*��`y����S��U��6�.�/^G�� ����O6]Dh[ٷj��
g)�q֛�L� �Y;�Z_wu]�R{R�u�+v��]�ӗb�P�$�it\p�������K��i��:!�&̓c���'������ڼ�藥e_����P}�u(*�ȅ[Ü�e4�A�rg��/F���T"lc�ꔢqs�m^�%����.���VP�7^7׹��cPHs�2��"ફ\�]�
���^npY����q=bÇ�5yͱ\#�m
 ������H6���=�k_��*1��R��LO�ã$L�lˀ`����g�}i}%��:0pa�ϒ����[���C��,����ȳƴt�{)�͕�<s�
ªW���u�>�� �����E#⟦fu<����6j�í��5�s C�<2JT!�ȅ���q�#����l�ܗ���9�z���Ɩ��b��ڦ������t��2H{%�$[�k��u�����w9��7i���}�aʯM����x���I��4���ߙD�x]���ijI$�6�Gȡ�m��길=���U��`�O����LKU���<=Y�ɫ�b4�T�Y4�)u����_`+�ȃ	�6�N63��e��w�l��"����GŬy[}��ӷ/h-H]о�ҍ� �4R���lE[y�aON:�=�
V�>b��ݎ� _l�vu��ܝ��X�����h;�g� "`���N�[}H�7D	�7#U��X�7x�y+����hn�7Z�oV�:Wz�p�{}������9/dnQ�/h�P^�n�����Ϩ�>E�l�v����4�t�L>����Y~����e�Ē�F6����s(N��K*;ԕ��cxhߔ,�Q��;�Т��M�ۑAPbI\���7���9'�*� 6d�>*��G=�/Tw�+�r�SH�<��1�3��4��Hp����%��_:&�<➞FC������/x�]�������3�tEV�M�0zsT����&q���|���Cc�^+�E�Va�^�a���L����~EON�x���w�`)��[��v�0g<�;e
>�J0�=v��`��3}���,��*�X7|�'���"<It��y�J�˿C��MDVW??� "\oͿ3ޕ���@���6��;Z9��c��wݬq�%�I?�y��^�X�K��T�}���x���9��n��J�4�Y���2����z�ꮔ���T���J&6ו�<�,���_�#�(�vޟ}ex�}�bb�Q����Cӕ�!S�g�)i2��C,�۠�յ3O;�T�SqD��8�\	�XBo �����H��7��}�XJkt-�8��c�x1��n�X��;Ṋ�����1��tH�\���{ ]�K�m�N��ܬ��r�BFޙ[��t��/�!tv��:�(��]^AI�ھS�wxBI	�{מy��=��k�S8o����C>ҵ��YϖW�	j<єyAX3���,�ze��Y̸��[�x��@����u�W��L�h���ڌ+bá��0�o������ʖ{����R��7���,^S���g¥<�`
`j+1�d�L�3u��b�V¾R��6*]�*ng�9[�;�T`ʉu���LK+�h�?dG>MY2yc������it���;�ה���t�uej�tM�h�0��@Ϯ���u�e��%�Rk�Hv¥�v�Ml�_���d�tLՃ�,_�4�K7T���6��b�� ��=9Q�',E�e��wIC���+�I-;���[2���Z���$�Y�Ԙ�P�(I�,�b�P:���FM\�t'a����Z0N��Cn�`u%����u�Wj�&v��O+�i����ў�9���CcU�������y2�g�~05�ǳ����:I:��ګ����fz�6&���:9i�{�n`�v
�\x�V]��7��󼨔�d�u����� ��L�~y"D��>�]�u�D��V-��_e.sּ��p׊��u�W����>��Ky��ܨi��AC�N�}��+���]������}�8hPr�: �)�;�9�vS�1%�t��"vvAfW%!ʪ����=~͜�+�|�R/�o�,�bo)1u='z�~�{�V|��9�V��iK>Q����[��,��>�r���b��((�(eX�{楱�B9Z�`��J�N�C���^k��N7U��+�.U�-<�>e���T.�yؼ򐬯/�6�[л�Y�|&�f��zK֮[`�(4dJ�UA����H���M�fV�"���JF���'i%�SΝ���(=޻�φ�J���T�`!�qZW��(��V,�mVt4��{ܷ�&}�I��b��]6�%q	Mo�o�hj+�%d��O'�86��,PV{hV�7h�׹3�e��z���\<����6?P��_����<��BN�ƺ��:������R��g�����Rgl���!�tyO8��0��=�Cl8�����8��sZ���H﬑I���CB����I�1�o_�����-�>���8_rq>a4é�=a���P�3�q|�,&ٝӶM3��l8���ul�,�{��IĞ9�I�Y s?~��u�g���y=�PY����{��CH���w��4��:/�6�22w�=C��	Ѯ�C�m�<��$�=OY1��x{M�)8��Gԇ,�|w�ݳ���v����9�{����35��@��*�5r�N��m[������Y(�nv��H�n���1]ʈ(ecV_*�A�I�����v�Yx��p]�ͮ��ݳ.$&�J�3I�,;qwk�w��o8��rݾ�\�':�f�N�;�Y��Z!�N��BH }���~�f]w���c	X��{�g�H�o$�&057����ٙ�4��:/1C�C�N���gl�g��݄����3��l���d���}��������o���y������}��0��H2f�7�����扏hLg\�$�&05��v���|�[�C����g��!�'z���+<N��W޿���/߿ӿRݔ��)&�	�}��I���2q<Bu�m�I�ĝCt@�&k}�N��5S���v���P����Ѽ�0����2t�P-���n=���~u���/��ri��Vt���,9�8��>C䬞�{��2y�'{�I�0�;��'i��ڇ��!���z���\�'̔G�U`�k	K4�g�Z����i/�Z>�i��`x��>@�V�)6�3��iwM���&���=�$�}ql6�d�ް�$8�׽��!��>��W��QI�����W�����V�ﾱ���'��o3l��'|̆��I�z��&��=5a�"���:�R@����"öm'���}`m��l�o	�_W����8�O�������������q��	�C����<d�0�;�6²T��>d���w��i�$�;��L�&��l�M�C����j��XN������;kzP��r����N&��� x�i�&�hO�9��>d:<��+=I��d��+4}��&���=v�=N�:��'<�1��M�C>a���n�{=�Gbtk��z=����:a:@�=a�m��8y`z���N��d=d>g����6�{�,;d��'�{�E&�oG5��H����l%C�s!�M�Bs���׾��<�מ?{�~�����9<@�'Hs����h˷�'H'��d;O�)Y�x��{��&0��$�>B{9�2W��Ȳ,�v��"��d�{�{��u�]�~�1ЙE�}��똗n�P8��R�;F6eu����;�Tɸa���Pw�h�4�j���Qc�]����h�8�;��mL]$��to���&_mh����ݖ+aLwiwRs#yаt����!J�p˙�MZ������#���~{�o�W���~�Cě|d1Ra�����:Hq�z5O��05-=Cl�x��0�S����$�o������wވ�T��+c� r����߀������c��3(�E�~�M0��d=a�����l6�0��Bx;3���0钳�=��m�j�֧O����5R�3rV�O�v{4��?}�$���DY9�A�a4�Y9�vs0"��5zÉ�	�f�0�x�w��C�6�0�d=f߼�Ĝf2��x>���UvOw!!��ٯ��y���>�$��ތd�����Rx턩ٛ�;Ḭ:3�&�+&Ӽ̐�C���'�M0�e���2�xͳ��S��}��}k��O����ߜu
���X��!_W'�;a�J�MXdY3�y�a*���I�Y"�sy'�8���N����bC���eg�N�:�C�6��8�g���]�:t���~���W9	��r}M3�I�:��l�|Bt{f�,�La�v�Ϸ�(�ԙ݄�ts�����7����m;32�N��_o/��4���'���t3�\>��}*M��%gO)'�8�����	��8���{g,�n�����L���E'7�C��	��9�I�L`�d��	���7�_�ΞCV���}�U��8o0�̇ɻj$ힰ=����+<|Bm�C��8��M����M�0�� q'��m�m�����;O��\����T��\��^|\~�����˜��I�=C���������|�5�:�<d鞠bN0풿!�Cl�wf�XJ�G��'���O� m'����Y� �~�ퟃ�׾����_SW��o�j��F��Sl�	�o���=f2m;�a�	��3L��k�}j2t�!�:H�q>g��!�E���i��W����C����\3��ouQx�����k:�V���H�ɗ������gr��ˠλ�tJ��#wN�ݔ�NX��tgp.i{S�ȫ�˕�)R���C�vW%�Kʕ��I�ud���y:�J}��r5��ao1;|{6����G��S� �{�Ӡ�E�~B̟{a1�7`q���vM08ô���ԆНNy�N!�!�Ձ�����=d���wy��q��;7�CL��Hw��,�݇\�<��gw�ӟs�g�}�{s6y�������$Rh�a��	�G�m6�����!�gf�	�!�=�Shz��m��P8²T��g�&�}��m�x��M`�w�������]y�s�����N��`t�߬8uHbh�q�银m�ݰ����C��n��O��rs>Ԟ3l'��öJυ|��UTQ|D�>~6����~��O��y�p��E9/��J�F��Nyd;5C;I�;��C�3x|�t����3������6�:;�40�}S�_}c�>���K���B�mox����6y�_j�Xt�_9��E"��o��O�����H���`zɿ,�z�����:;�:`q��>d<`yl��C��i�����:������ַ��ל�~}�n�םu�&�&0�o��z�w���J��Y�'9g�y����~�E9���x��Ht�i�2,�mTM~_h����݊�g����ߝ�y���W�l�$�6�-���4}��>a8��g5�v�Iޒ,����C�I�Y��`E��z������Ym�	ު��C�;�����y��wߞ�����E	�1�)�N3}Cl<d���[!�d���X�8��fI�������Ne��}��I�i��a�'W��O�M0��Ϯu�\�e�����{���=gHN�$<C�x�g�m
�m�'���d;��q�����,���4bI�N�>։��"�No	�'2��>��!Xq>Oy��Ow�^<���߻�ϙ��9!��p�0�|�x��Xzϐ���k����u;���$�t}gi��z�dY8�O�$Y.O��RE[���;��:�6l�wW�zj�|����`���c���T��],g��H��]Ύ��t0�ټ���Y���"���9,Y����kY���=y�b�q}�ю�/��M
�gT�Q�����Ì�0>sr��t���%�fEt~�x��o����}���}�oZ��'L11����v��6�'y��C�t_�g�N�u�3hv���<��N0񆧔�:a6�^ى8�!:��$Y6�M�c�3���3΄?GR��\��;��2�-���U_���բ�a1���I�q���p;HVb'-�����Ş2x�P;��m�l��=ya6Ì4yM>�M��+&�Ўs߆��Hc�7� ����������x�R$�G��A;Hu���z�����o$���2gI��!���zu��'L���8öJ��ЛH��םrJ�|��b���ݽ����\+�}_��ǌ'Sw6��,��'I0�9�2�9�ڇ��!���zϐ�G>���'|̆��$�[�P�'L���u����ϼ��1���l1�d��8}Bm"���,�I��m��XO���M�}��t��S�o�Ԇ���4g�OP�d�3�1&���z�z���{����޸��3�y���g��y�	�{�I�m!�:H�m���R`mwO�d�MwM��q�Ώ��m�'F���!�6�g5!��sz�g��f�}�|�����ߞw�����϶:ε�@��d���$�0񜗘x�=N��CL��Hvj� vɽ�w:�1�4wO�!:@�;��m6�c�v�m�|����c�<���ֻ��u����y��]���:Bp�1a�%f�ts��+%x��a&�,}��m$�<=�!��|d;5f v��,;��C�+����'��M���}�yS��)z=�j~�%:���華}�U¾�S�%a���I�>a;�x,<IYĝ�$YM�y��iy}���H���d=dߖC��1�OXw����|��\:���q��{ϳ�4�z��i�3�NӸn���Cĝd�ã9��0��jE%N u;�H�Y6���X`|�(s�$P������A&V�v��I��~�]�]sE�O�PsP�Mu*J�l<\Z7_0�{bWuaJ7�-��w���f�"m�����'��8�i`m��Q|`\��W��*@��̲��x�dJ��A�3:�ތ�d�@�,�3��:N��G�k"U�]�Z"�.7W�N��uap��3on����kYUke�uV��3��[wxh��Mw%	�)�0�E�vp��)�QtEVW�Ul}�i��#f��T	�����(�f�g�<��3�D���s8���ħ2�2ƌ��R\��W��z�?�o=���>���&S�O�ӽ�t��Ӽua�j��>Ti��b����s��+��A%�r��2Ao�T��lv.�_T�ћZАĥ�N��i�\U�Ͱt�5;#8�w��Vo!WRM����u�I����saYarԓ�/Z�q��ux�+{�Kz�7����{���9�&�?f+u��B�4��}��Ȧ��q�8$�ٜ.��՝aţ�;�eҳ��t6�0��}V�A��-;��ל+: �󂓑=E%xd2nQc��)��U�kw�pԐ�c�I�w�ܺ�|���L���/Z��36>�I�cM,=*5��Ԗ��*� P���������2�޶;p)RU��ڳ6�����-�EB
�j�읕ڃ���*\Hp����wP4�kJ��,-uk<44x��n0ucS���C*��%C�J�u�Fjw�\l&gZ�T=�v���[��	A4(N���v,��3TIv�z�t�t�ϟ��LQ'F�-���&.mV���j��v&�-�,��X�Ջsvڻ1r�<���J�v6w~�!�K9K��q�NH���ׇ�E�\�a���ԝ�*V$�&����R�,d��ڽ��mr�O�3X��ڽ����7q*�
���X(jq�('�Ҟ��P���eu��s�����]u6����6e�i���0���|1��z�R�"����vV
O "�=b3��*�5v�m�Qw�fw]�k��%�[�w���a�n�����t宻�NӾX�(i�H�QB��+�V�Ǳ��wA��RZ\ rtJ��k7W�"�+�J�&�d��o�9�m�9��r}a��% ��y��Ւl�st�e,�_am<��?����祁���w�cJ
�rN�D��3GR܆�÷w�kldt���7�+�e5���U�j}zo<�D��[�;�3��N��cZ-�%mo��z�=n�Ө�+okt�֯8;+�K���Z�X�L.��7o�ۭM;�.�tI���֖9Ε����M�y��奉u
v��M�ۘ��ˮ�(�������E��8��nGȧ�B�J���q����-m�w��(��5jL��(�wݜ�,ݾ5�����F&��1��Z^��3����w�)�x*�SѺ�:�z�p���n���������	����H�$�2ŋ�uع�:���|+�>4I�
 Ae��A�
��ɒVEU���j��Q��Z��!���F�F(���+,�4̙j�c����QQF�D�2�*��Ub�E�UƠ�#jJ� ����J5Ve����EV#�����")Q�[*F(�j�J���*�Q�*���UF"*�)4�V"8��Eb�ԥh�TmY[J*�5��" ���J�QE� ���֌�D�QDb��b�����ңT�QQ�s1�%c�UY���+EE�J2��KB�m�m�kUQ�1��R�
ZT(��D���4��*����#4�*�2)m`�Պ,m
�m�Ų�*.*���J�҂ʕ���ʮP�!�,kAQ\J届���Q�S�pB�*��TTQXE�QPX�fRł�b��-+Y����b
�[h��B�-
�B���۩ۀ���K��>�$9����=˱(���Q�}s��
պ��*�L���Z�Q�t'79ܜ�Jz���?W���}F��ӜC���)a��#�I��tj�d<`j��6�8ϐ��0�_o�O�Law̓O'�}�E��@��t�Y9�v�>��ꫮ��v��������_��⺶�6���N�m=d;5E!�6ϘvȲ!��)�'���Za�%g�ul��q�P�}k'u�kRx�k����W߂U\�'tR�k7����R�������!�d��p�d�I���O��L:���x�u��'��C��a6�i����q%gXd��և�}�Wدߧ��u������;=Oܓ5d��|�<d�Xg� VO��f�C���'�C�N̡�g�N��Hx͡��S���q���M3{M�)8����{��<2�1�E��s�>�﮺�8C�'7���%`h�{�3�$^��������t��8��ff�C��^b���l����:d�<N�M�V
�!���wd�ZB�ø�ɿ���s_u��2x��m�d���P4��L�|ԑ@���c��}�x���i
�g���dS�^`��O�T�a�%g��h��s�k�o�����.|u����hp��>�M��>�2|�!=M�);x�hl���Ρ;Hts|�=OXLN�7�x��z�#�*���_Uh��Cw�<���y�����zɦz���0�%gi�,��6��8�S�c'���}q��r����i�>N��5	�C��}�z����|�_�U���w�?+�2s����������ɼ���d�z9���3��XvȤ�|Χ�&�,3�m���5�I��'_\@��;�	�C��-W�~߫�u�?w��zҞ����T��hv�|Ü�$�8��fm�z����d4ϒM;��4�!�;dY>~g�@�;�۲E���6�׈Lz�Xa��&�l�;�L����/�Νk��g����ۗL��:��Sö�M�R����(K����W"<*y��X�Ó� �p,���8�j�'u�R��%�s^�r��.�kk�/�)tkj;5��lN_i
e7׶��k@��񋜫r䥢�������NsfU��u�{�����Nw֯�1!�6��0&���9��=d���s�l+%M��$��Ù���I�w&���'���f�vȤ۴:<�1�;�ܰ� }{�^a�n��7���^����=a3���O�:��'������E�L��$��d��+>��M�)�}�z�z��d�t'����7��hY�v�ʟ���Z����!UX>��NU����������6�2u;�C�C�q_���l'��öJ�Ro��"�i����M�SG����	P�nh�����{���[��[��5�	ɫ1����I��]�0� x��hq��><�=f��']d�ã9��!;�0Xx�^ w�"Ȳm�����{�o[�}�/w:�p"��r_r�d�:�d=I��C!�OX{���ǭS�'�Zz���'�Ra�'[�O�&0���Rt�}ζ�ߦϽ�z5�y�o�s��ֵ�,�<d���E'���y���C��M0�sYXq=d;5E����:�Bxͺ��q��hq�l��!�l��q'��_=��}�E��2IQ2��{���}�~o�x}��}��ɼ�:��4�Y7�vs0"��4�8�0�ar��N���t����,��۳�<I�c ��/�?:�c{���;�~��|���m����C��;dRa��ь��:��'�J��������I��i陒Hz�,��	�������m��׆n�n��j�s����ό��󆙌��m6Ɍć�m��+�5>�8Ȳ}��J��y�gvH�No$�'`]٤�a��=��$=N�fVz��^�\�~�s���o�k���v|w�P��2v�']�'xé�4��&��|ɏhO=��N&0��2)+�o�$P4s�jL��c:��'�11����Xq6�}�[�y�]{�/��2�?l&��C��Ѵ��y���;-�^�-�ŗ�OR�d\iX�ܮ��z��}��ꬿ^׃+,nĤW\Ӏ�/A�����VEeq�*T׺�\�7�\��[�L���V0�d+�)S�pGR������b5�:N����ݱ�z_�}�U}T����N�_��PU}�~]⇌�l�I�2Vv�{I8�hx��0�aߴ�N>!:��$Y<ݓ�� q�7�4H�y��P�<a1�}b�_����ϗT�<秀����V]e����̅C�u��2��x��z���'v�Y���	�E�t�z�6�S�c&�N��@�O9d�����R����o	_��W��NQT�ᥑ~rć9ϵ_XLg|�I�=CN}��J�gl�o0>g̓]:�<d鞠vj��<d��tyd6ȡ�ٷ���\k���|s�^N,��_�jw��ξ���<I��No�N�0�7�2��;�'��	���$�Y��N�3�OXx��3L��k���|�Ӵ�0� }�Tv��������}��/��;z�����H���|��,&=n����tf�N�a�v{�jChN�y�N!�!�:�aY*jo3�I��e�����}d4�۴�5�w7�������~:��,��a��!�!��ϹI���m6�c�}`q��l�oX���*���E��y_�ι��~3Ε;��ݻo��O��!�Sp�9�~:&�������F:{��"�u������ὺ�m���g���T�Mb�N�}7�ك������+}�
~sҺ����>��2�͕NW���7b�BN�ӯ�J����_zƹ�����X�����;�%�ub���`1��Ghz�}��i�﮲J��,	�K؃E�w�s��HU��l�{[��T�H+���lm1g�ru�Ut�u���	�0��}H�H�g*�6un�Hu5��b�.�u�l���)�%q��,'�:̬ق��5��VN����`)7�lq3�<-�ɫ�'(U_}�}Ua7�HN]������Bb�w�Cr��o�,ɄxT��U��y�E靚g�=�8b��/=]����i��̹������� !ͺǝ�Zss�|y�����\"�����2NG�q�_Io�tdqT�ԛ뷧6\�@c��|`ɷ����p�WVܯ��𹰥���2��P��%_N�޴�X0z��:�{�����92{m�n�ϻ�1���.0WI�zy�k�:�"�q����,|�V�Gվ�
\�:�b�QOnU2ʧ�/�̓��1�^��߸G�ō���ITY�������
V'^��q�|fz���C^�>Q%91��>2��������{^uu~[S����s��͗\[v�ͱ�t�3<#�]���/څ��9�qz쭔ʛ�Rי���(�9��Ὼ6���qm���P�p�N��KՔwS}�Zݵ�W,]����Cdk�Y�e�aU.m��kD���z���Ռ��Fs���愒�:���!�� �F�9���[}�'/M�G�Ѯ�f	\+y):�`OjU����M���v"�`�"��q��n*�ﾪ�4�z~�s�8�x��S	��Z_�Zǉcy�Y��t��m��΁��T��K7��7��.r�͕��@'4�P�~ʭ����%�g<����h��6�kfܪ�%�М���μ%����ҡ��u�f��D���f�M��R�v{㽴㽮��q�3o��=Bd��5��#6v���ߺN<�b{�A�_@+��;�=�~������bFd���SZ�^��@;��i�P���o���d��u���j9+%�7���ˡ�=����ۭ>1ۅ�s�;1�y=��1pM�#�p��F�qʆ�5�s�+ݜ���ԫX2{/�<쿲lb��������d�)���U�ʂ�-�9^�Ĩ�N�V�	[�����,^�o�p.e6��!��[g'�wS*��s�:3�����ۢW����r�Qkpv0�_'��o/d�z5LV�gٰ���?Y�W>׷BUˤ��Ge�������(;��(5���6��w���)>�y ��To�J������.�+d��B�j�]��k�=����ِ��;5���ﾪ�屮{�	��Đ��E�y��W��L��L��n���� �v�Q������{���L8��7�yox˛ҧ�l����w��o�bϳ7'�*��jN*�^�?��۫�g}��o?��1�������-�}$��~�Ƽ9�^3k�o5&���uo/����YE?fl���Vw�Q�S��$��L`*�{UB���מR�o÷�U�\���k���Y�>���m�S[� �<�:��k�p`���Rᝏ/�W7�f�k^�2�y{ْ]�6���r�oL���W�^?���]�YN	�����hl��h���qĸ>]���{^w��6f�d��$�����{��2�I ܴ��ꊱN�7f_ʜ�o�t��b�_O,�킞3lK�W1�#��{�����|��Z��i�+fء}�.�b�ʿ^��{	�,�<v��Ĭt_F�E��vP�aL.!�ku���b�����JQ�y�lfj�1��C��<�����VMyF�]�eGA�Zv����$��Z
��)����)�T#��;��qּtP]s�l�Ǿ|�]LI��f�߻���1��K^K�G��������)y�fx�潿�-cʠ����9_�y�)f9��k|��/ �#�~W�.�����+�vA��;a�"�^Cg��	[t$�tvy����=�y����hJ����l��Ul���~�d/�����bvQ+Z���ooh6����wυ#���;�����xE]�J5��F�耓rC�-x;��N���z����`�����zP�|��1��9�Q<��������fzn8�o����T&�^|�X��m�R�g7�z�jd�C���o2b�{��1�ڏ����rA�ɏIc]W	3~�j�~�+��w�m]�K��;��W4��������~���)ͧ~���{}�֦�T�so
.�gl�PeX��l�&�s��d�&I��>&�m��SM�m��:�}����%-��g�]t�쪾��H_zG������y�2CN�S��΀�ÙlV��R�Ĥ�>�68����` }*m,��XClK8��gZ|�e�!��)�u��I�畍o $s�.�{�j��g99�ڊ''I�K%uvӗn�k�w'-�q��D�`�4�#'7�6.ff���Ñ�!ǋ���3�+�������n���-,h�~;n�W	ro�yV9wX�9�w�s�P����Ǜ����k7	���Hee��ve�H��dC������ �o���fd ���۱w~�vc��>�	���Ru]iٖ����Uآ[[�h��.�m-�If��[� �������r��eϤ���y��?#YG�It6�0�,:w�8��P��d�O`2���Ni��3&
��\�ߕ�t��=�y�e:Yk{���J̊�هY�]�VByŠ.BH�]Ob���	+i�d��;��?Og�j��EW�}�:5]�˜��s��/�1>���0��(���[c�{�]R��m��+]B���/�ӌ��;���U�MV�bU�fz�K5�={Aq�_,�f���f5�=���z�;�h�:�P��]阯��J��+�E���u�q�C�������)[�{����+F!DI�p��ԫr�=�P�s�2��T�{�W:xk��)ۥ0�
�ՌcvMv�X�;q#��n[7��4�G�U�2nt��|e�74Z�;t
��r�v�f�Νb6V�t�Z��cY�Nv��}U��T�gO\#����������Sɗ�n�������~��zv5[�9�=^���':?d޾;8<�Nd����{�w�����nyR��k�u��6Tt��A���]>�:�u�l�uŶ�ߜ����+�OAJߺ)�V�;��K�������#J/��,n��+�]�tǆ����_��sh��5G;�?}2 ��yT5=ϥ��I\��+�7W$>:� ��N=}��<�6���ٲ��P��+exu� ��LP;����.��[~=��߱�fG���B����k��dМ��:��n���գ^{\q�Փ�����:S����wȹ롮gk��dM]&P���Z#�Ɗ�<�\����^��w�VMv�5�_��=����^߄��gk��Ê{r>|���v;���*�Y{7(9���̚��tt��jvx'O�=����v�dݘ�����Gv&�{�;I�q;sm���d��[�ߒ���2�����^� �ZT�C��Z���ʽ���KW0S�M�SKȌ�?fR[옄���!���j�}�L�\���;����j7����r�m�PN +���Xw�w��ƚ�ev�?Ϗ!�d�tu���̯S�&�^=�ѿm���F���ǫ��O���o"��3�U�=�ٌS���&���m]l����u2�;^:���G��=���KӬ�ZU�xu� ��7��oh��7��׳J�^k׮�_59^��0'�*��0"�ř��Ń�Of_��<pW*Y�ٿeo?��?��yy�ˎn����:�ٞ냲�7P��mZ݃��x�1���d���c��/w����8�f��F{�+�5,F\�};�ˇ�];��}K*u��G�z6k��hAL����}�d>�������S���%>�Lq�Ú5�6�f�ڑ��Q�[Uެ&�秜A�x���_�ܙ\g\�j�}1����y
��י�o�b�uu����d�	J�99���ٺ�ݵ���S�du�8��p�ڀ��x��f�>[8���N9�}��av0�v#�{�1��gA��
��(Z̭���H�y;�t36��ޭ�߭���3��k6ɦ�盚r����΁�;5�N�ԯ7�D��E>�n+��OwHU����_
U&��ץ���-�NV��y�Z+�%��c[e;��4oכF�'-;��ֺ6��M�z���x=.��?m����q��9-�Z��ť(��}g�:Y��N!��v1B0�a&��淴�Ԭ,�خ]�]��k�Ł� ��[0Gn��J�!Z������ziU����,6��#��D���1�ǹ[)3���+���(_(rt�\��#n�����9��O�G��]���v��ޮ�3�*��*q���n��:t���>E@M�nM
 u�ܶ�u�z�v�Y�.l��[�hk�9�x�� {H�T��������c�\B]Z����/o-�������j�RjZ���=��p޻5�ұ+&�����ft�QT��25�
�s%os��[ x7k���Vj�X��7�-/,�+�3\dQ�G:�b �E�ٕ�_}hkV։]Ʒ���rfg:9N�9i�C�|S��F���S(��VdŖ󸁍$i�D�F���0���ڶ`����i�7�b����J5�Ԗ��N�F�7��:�B�����j��S��5����|�﷒��|��I$M-�ʎdX̮b옛�][+%nM4S.K(^�m^�P�6��ټ����[�r	W��0�m;�챱�i�n�9O'4V���vy�������RG����b:����u9Ԣ�����w�����WAì��R�W�Et����V�T��so$Q���'t���t�4@���� ̡�`�Y[w�;/��-���\�"�Z�*1R>�A�l�/ڿ^�9 �*��J�T�^m�&*�*����
`1ʲ�-,��J�.��z�}L�W�u�vR43n����U�C�k�i��
 ��w��C�*s�n�RR��]�-�]�q�3l��i��Σ���E��ٷ#��۸��v�fn+z�"]��wd�P@J�,s��M��eA���j�%�3��h���s�m
w]»u��'�A2��6AdZ<��{��A���ub���vEٚ*��B.6ie\���_t)�QLߔ��G�:��[.����r�
�Rn잖k\��Z���z���;�Vu�Zb_���5�%�`�D��J�-���r�U�3��'��em�>8��&�����$����l��쩿��xk.��R�݃��:�M�t�.���I�S}��3�Yf�L�y�-!�]w]��BV�� ��M�����E��/PxD����ȁ�4�	|F�!��8e�s�tu�.��Ύ��}��3s��1�s5;f>/C*�Ӱ��܍���{��ꂖY��Ub

F$�����V+�R�*ZU��Ջ��+-(�b��ph��+(¥�+*�b�UU(�X-؂�3�+�iEUdT`��Q`�mQ����l�V��p��X��1F���**+-��"*±�UR��AEF#�J-kTJ�%F�*�Th�h+��Kj*(�UE��([Q`�+J�b"(�r�1S,��KJ���QF��kZZ�b�*�m�&R�[m�)J*�QJ�Ոō�Յ���%kB�c	Qrؠ��,#�Z3
5��KK"����Y��+Z��LaZ�%j�AYZ��V
" ̵0�-M%H�X�TՕY��e�bIR(���,DF0V��D,�-��Z[Q,\F�,�Z2��+b�(��-bZ�",�*(���UZ��s3�m���k	�*#� n�O�&dΘ�u<s�wu���L���q�v	P]�}#�#�G^�{�-��Q�WF��u{㽍�}h�e���������o:C�.���#r_�J�l\���7�7��^ν����p�:o^�zzrN��j�;3i\��e�yO���{=�KX�M,�֌M�uM8+,��~��2��[V�#Tk�^�;�3>�����e}ss�d]�cdv���%���U��|-긶i�}�^~�5���D�3gJԷ��z����œʆ���~9瞪Y�2=3���ϳ_�q����*HUs���J=��A��7��# �v{�����z�RK뵭�REy��](�k!�9^����؝�u��w�(���E�y���-�n�o�&zþ�2�������6=�Tحs�f���k�̛̂�]�*<��}�C�����2�05L�/��W�W�������}7D�r�։�s�KGn��k��g<mj�|�`�؁~�ε�W���XTb��1w�<.��[W������Mx��G�P��Y�.#�n��)�W4���:=VR��q�Q�S(@�%���I��.=&��a�W/	�ϺČ�{nr�+r�dǘk���q��n'B�=[���~�����B���VwƟ���Qq߹y�k�Lo��w���լx�k�a�P��H���:�x�D����_�K�ӦOs���p��*ɮL>�Q�׺�ꕈ��\�:Vk�o�a���dwU=&殺��1>C�+�����8����]k&R�s�{9�6��F��|���o�Vv�h-h���Pk�z�f��lE�\��yV9w��y�]9�[����}�����tc��y�\(�,j��_���_���)h}v���~gt���_����`t���0�s��^d�`j��/����k^S�t��O%�:��i�{s��t=GҦ�&.}##|_hb-�^穲�����@�J�{&`;�=�]{���*��z��$fK�<���*:�)a2=���Dy�#Y[=��%������}f]T��g�^B�ح����Y�pvT+��ʌqM�S*Ĥ�v�eOTu���J�ϕ�b6Ӭ£�\7S����Cr,������=5��'p�x���΁q�gp�	=Ma���L}K�F7E�qn���i�u�ddĪlu��ӕ���5-���;ci���者����Hݴ�W�ͳ&m�sW%��ް�P��<u�L���\8��u���	�L��^g�iV�d�X[1�庵q�y��r���>ǎ�hO^�l�{35u	Ne.l�[����=�T%C�q�UG�o}�IŵϽ~~&?Nĭ�/&��4ʮr�����x��M�z���R��������)w�3&�(���>���©�/��+���${�^��c���5\+2L�Y7d�������u��?l�^=��k��|�mNpOi���>a�M@x��շy{Q]K���e>�:9Εl�����W7)���_����$�}� ��W�1�^����n.ϖWuה_}��}��uѿI�.�[��v��>�g��e�N9��d�������<����<������q!stm��Y�et��8��vl�� �^�n�e=�G������^[xM�R���:��y��@��뺺��f�r+�R����p�Եn���	{IM�W�n�d s|�[Mv.��h�X9��,�X�ܜy��h��?4�;�Q����ղ�%2Z��ؔF��}P!�L�/���}������k_���ko��r���S�}�u�1��}�6u]�S��;َ�� �o�dG5��w�oG����'��%�<.}�0i�]����)�Yᷔ�ٖ�溷��xk��P����(��;��l{�~q���;������}�\��Vf�4�megP�_�a�zN�<'j׶7^ͽ�Vm�q���PyL�ǐn�C'+:�j��W���UϮ_R�E���#�8�wڞ�WY�\��G��"k�Vԝ�_�+�4��bf�=��Ӥ���"+��Uҍv��}WQ��	��ū=�{���Џ�H%g����FO|�z�e2��W9Jt8nw����X�A�&�W���q�;�'������K܃���F9r�'Mԙ��^3o�7K��{�U����VȱP�{u0�8/�o1���N�k����Ve��i |/.��8TԆjM��#)VA�,f�ȬyzZR](qUضw�#�v���ʾ��©e����^�;��O�#u��K��I�����+9d��kݵ�ɩ[3�t®:��$��z/l.��5ЙQgN�~�����N��52-���m��~�����&oj�6�|���6k�u֯-��=X��{>��d��yNm}ژ�_"����ㆤ՞{��Þ�܇y=��c�̧�̦ۿ��2�ι$վ��0�~�5����+|}kY:D����%Z5o���$.��?��lN歷u#W��|�s깄t�߻h<�e��m���Cs��n�I��lNfζd}J�K�v��@ׂ����=$���mA+��{n���߫��>�I�ߏ{�m:І��a�Zeӧ$��A�Ϝ�����Uʄ����U}�R/]�왭����>��9��U_募꟯�ђ�PyA�~�I����ڋf�!}�c:��C�Mߕ�n�䜕���.����L1dσʆ��k����?/r�
��Z���Ӥ]YI䮦��f`��\;�뉯Q�a*ޒ����6���ډ�*�x���˱��ɰ"��I��7��٭�[�fmw�A�{%v]mq�K%ĩ�.��p�����I��ɧy]C)�i�M�3Z���5�w�͊�l�7�\���������\j˝�i�F�l�gd�0�!��}'tKq�7?�U_|���P������\���ޱ=Sꏅ�=��q��j��y��Y&�C�U��Q5��x�__��U��X�����
�S�Î��당��m��(��eTv{��X0z��m�J)��=�;��9�������9�L:L�by���M�O�h�Y�iu*>}�1qu���9�	/e�\�{s����e�Mӕ'��wn��O�<{/`�"��^N�ǯ�k�]y]JסV��/ӥ���.{��ߴ�;ٵP�[Ay�˱�܏t�5y���%��<Y�u9�z����|_IQ��i�ݵ��6���x�y#�Nq��NDqz쭔��-cϖSw^1Vs���}���|��½���^�M��m��^O�p�y���{�KX����*����^�~�p��!���n�tΜ�w�9{��ׇ_Ս��u�ƍy��L��E���{+��M�t���w,T(�X̌[hMT����Vj�n�t��9oeӮ5(�gv��.��vZ�K�![�^-�|��	[����'d�8�;p\p�z��uP��Kk�su�J�o��w%2/&�ؘx���mm\���>_���~�l��mY���9�s�9��+��s�]��^�ӯ�J���ۆ�'<�1?>y���+Mz���O�ƃ穯G/�0s�=�������wk}��)��˰�o{"��ezy�����	����όY2���'V�M�������˗��4���ͧ��A�b�ufE[0�����j9+!�SwHL&��������^�oO�C6��\����'���W��󀯹�d��7dNb���@qkY��H�����n�X��Jړ�~;=t����}.������6s�5U�.��~�
����'�U��k:���3c��P=:<뇠;�t|����L��\�)��9S�J�����^ͦ����OfF�ꕉ!r�5����=1�^K�9�r����w��hT�p5V�1��ӹ�g��l5Y�sWP>~����Ǽ}���Fߍ��|f<zm�u��B��]����M��R;��[���IyG��X;�iy�f��j��b�{[�x}�d>���8n4��y�&k�R��n��vn��j��*����c4�;�+{���C�wG�R��2^�so�0�i�7�M����lq�ޫ�wG�����ٰ���5u:�V͗��5sU`�zǽ�/t��8f�窻�7�(t��4|23ۋ��VL�^�ᤄ�4w�<��.rsל��5�S3���S�� 	�ǃS؍�KC��K���v��	�3�<�2}O�7U�;�9̇��+uI ����~ʹ�S s
�+�ܩ�Z�u���.���~���&���eyׄ�7uQ:r�M�Γq|{R���R97.�����3;_�f�;Ϥ�	��KѬ�U�U�I�l�+�T����U֝�ʥX��ҞC_�T�kNw��El�NU��[:f��z���ә��!�/�O�6j=�X�^�ڞ�᫲�q�6d����g]tY,K���$��|�_�?��i����h�z���]߲H9[�7�z���ؤ�XϧdL/Q���X2{��dH8_z䙺:�]� �H�b�u��)�-��y������8Vk�!{X��K����.&���#��6�=J��a��^䭽v4�f��] �s�]�[K��.v��ǔғ�]Ɵn�S�9�3�[̋Z�r�Q�^��_Q����FU��?s��'�k�WJ=����{��Lv'i+u`��W��ᗸmcz��{�+뛀_e}��+�ʺ���z&���%f͛�¤{o��K��`쇹�`����gL[��1�ܹu�3�{���l���~�ɦ	��+��6�%S���aǜ������<�Ok���3�~�c[�����v��m{����IO�=�V'�pW�{u���B�3_I)�7��e3cW7�s��}T��\U~�7�ټk�5 �{���j�LN{��N�g<��d�=��L�3�I5o�03��Sd�W�/k����=���4��T����*��ܐ��-�p����H�=2�����Û'8q/Z>�;ݸ�Oe#����]�o��M�y��v�������MXS�o]5)i�iٷH���ʨ�n�g��͘�a��{�ֳG������A��ޔ�ܮʃA����Ĕ���;���˞�0�RO��v7˳+�9D�s��u*4{7n�[��r;͖̤PfB����
�T�3��*��y>��d�y��7W,��о�C���=�:��䧔�YJ��ˬ*��s�y�O.���N{}�b���]PO�e�A��r?�ع�#2�9��g��K1bo$~V.`yA�I��+�-�[6�_zF�1��8[���w�}����k��}g������"au�T.rZ��eڭ�f.~|T��[�*�g���3"��u�{b�IY���>F4��ė`��^�ۼ�	/Z��6r��o٫������O�c*z��g�~
�x�G��ݞ�����N��Z���-�cW�핌o��&�0s�W�I��7�9�Ӈ���G��n��ˢ�e�����y�36=�P�{�p��I���=Y]�Hz�n�߼���<mj��#����+�|.q�o�[T��a���7N}'���.��W/ק�����Wg�_�����:Đ�\��M�8<��d쪝2{���x�ʾ�H�x$vG�J��B[<�Ůgb��V�gow���m�#I���^�q�o��7� ��[1I��udT�b�.�F��)!>y�g]NJ�ٸ���e��H"݌�\qC�}�5PS;��4���Ƅ�Zgr����=���yY* �o,��1�؝�1���B��9�s �/y��	�����2Eeq��-�t ��:��u�fٯ��w0�b,��>�ma�ݖ�ba\��.B�u���͋���}�ֽ"��=�6�u-�M.���N�%�؛�{��;&��� ��-,�n��CmE��Z���p,�����}��5S��N�إ����쌔�m��<�g+�#��
���Y��~����::�0����un(d�y�[u*�;�V��!��g^4Q6�u�w��@����&v����Ye�P�x�ъ�]�TB�Eff���G�N�%Z��,���%��Y���e(���@�I ���oCҲM�8ۮ��7l�yv%ɦoa��O^Ku��N�s00◙�zz�ց�S��&��R�:��ۼ�2Y���ծ�鉋���W3P�t�ޔ�Hh�����n�c���Y�O;�� �����ڝ��ͥM�X��Pu�],wAj�;���*uJ�����V�CD@��ӅN��n�ʴ��պ�f�����sm�"�)�X�B.�vX�0�+�QڂV�̽(�ĉʳ��l�=��Ӑ�Ы�z��gm 3���@��/�R�MU�ע+,ٜ!+d�7NtR\�������L��O�/\�P-���[�2�$�d�)t�%�������-ݳ�t	��͸K�G��`la��q�=�!�r��I��m�0r�*��K��"�'�c���-��v�v�8���s$���f9�rc* �mw-L(�0���V;�+���ؼ\�:ʚ4�N�[�1�⓱����ޘ�=���%��CB}to���v��#)��,|���4�q'�]���]������|R�s8��!.J�+_mh��W�I�`}�8�Ù:.ʷI�j���]��3��h��a`]9I'!���,S����!Z���o傺�X&"z�튁�`bJ��g[Fud�U�v����JqB>�!� ��
�I���4��ȍf�α���:�G<�6Wfq��zkgu����1]�ŧ'e֖�e�Iv����Q�!Ɣ	چ�u"i_D�2�7\�c�6�2��g��7`��g��A����Z��[B��@�>��v��c"��2>��"�u���Ҭ#�پ�ZXK3!fAِ�s0�ov�L�3O-����^γS�(:\��n֭9ni�p��T^U�V���G��ioBWKVwVa�8�w�_ROv�f}��c�o��[z):�қ��:�`D�)S�\�렃ۃY������}o�jv�wNڌpz�yТ�83�*f�yG����йjf^ԹD> 44@!"�D�U�+
R���K�c�QkX6�[h�1�Ŗ-��V(���Qr�q����mkm�ڥKB�����(��+`�����Y���Pa�i��X��chԭ
Q5�U`�UPPF���jՑQ���U�ب��1DTATX**��*-�iFDAUH�$kTX�E�"!XQ�UQ�E1U�""1E���(�V,U���*
*�����m�5�1��Uj*�31De�
��V��Tm�V
���V +kh�QA�",U�U���E�TQ���b���ZKKF2�P����V�Ub �%(�TATEF6�"�m+b��Tb��
����*TEb�1X���Ҋ,m�E`#X�
�QUX���"�0�,m��2(
��Q"��b
�X�Q#hTE"(*��Ĉ.ZAX+[eQQb�b��X�X��Q[h�2(�b�QQL�8

2*���*�DDKs%EDEPUQ����}�f��]�ޤ��ئ�[�7"+��l����,����f5Q�\.u���{}��{Q�]�r�TZ��f�H�,���f�N���H�X��,���Yγ^�;��{*�G~^�u��&�ҭ����G��чr]�e����m���I��cl�tn��z��o3eOsh����'v��� 	�ut7^�m�X�}g������rj،jwU�I��珄\_�\��w�J�@��z���_���B�7D�o=��6C�n�N�ze��?�������(���9+*��N�&�Dy�yF�\�A*�_�L��ޗA����r�� �>��r��ZK�w#ܾݘwΑ{S��b��b�u�7�xG���)W,��ފ��_n�~�o����l��P~�?�d�Gc:�dT6a�zP�5u�֞��q����];5<�� ��g��!����ٞ�_����{ȯ8U��^��u3gC��W�t��{�`!���{����r칬��<�H7�;s��{v�s|� �g=�6�U[�����*[�O��2��G`)$��ְ.���U}��B'�U�Ӗ�e}2w��٣�G1o"P�u ��c�u���ٖ�GCBR�WNzwXwKǉ��� yN�>���Ӕ?}�ǲwJ�[�^?���+��Oa�����NψOj�P���W��J=�oy��0�[���Ӿ��P�s��Ox�N�4&�^b,ָPc��.�����lmj�7 ͔2�x����c�*�Ǻn��R0�AY�x�%�U/������Y�Q߯s��:����|u�y6������`�[>���7+�5,6_���H���Vﯲ�T��YΖ͗Ŷ��p���S�z>	�^�:z1�Λ��y���5�>�\6�t��gRL�<�ωo�aG1fi����I59p�{OrZǉca��Vݜ�7��%+p�����������:������� �t����������mL��97�����w���w�̚7�so�����1���$���s'����1�4
W�a�{ـ�K���wӓ
k���QkpSTc��
��<���%�+(��w`�y�$���3M��ɏ���Y����%ɵj~�	����;��u$ȭC)�QT���v����w̚�v����j����XE\�o���``o��d�C%.zm�Ew<�7��-�6�UQ-������N�o}���U�=<ճ/������a�����s�h�{=�>f�.nuD.���y�yB\��x��ަٶ(9�,gVd޼_j��U ��N�-�z��V��u"���"az�u����穅���yҍǏ�K�[>~YsϽ��N���􈪮|�أ��'dL/Q�%n=��;��ǝ�[��Q:ǫԵ��f���ϛղ�UһYOa�\~%G�po�����a꫒t;U�����Y����)��~�L�j�R��3�-n��)��>����O����P�ՙ��cO,[뭕�uL��%�Y!��_s��t��.�S�C�{�7b:������+Z���(fj�ά��a���ս����{$?s���U�87�X;����v�gzo˩�;z&[�o�7��7�OL���˜�j��92����~��~͡�9mx#[Kq��r��y݈Ss�[�U�\�w��{.��Z�*c�5\l�!�����6��O��Vjg��zU��mh���l�}��ˋ���A�̔�d�["e��C��4k�����Y�\�k�8S�C.��ڐ�ճ�N�bV�k�����ݗ��8+#��z���߹�req�u$���1��[[�����p�}��,N�Ż縼6��R��6����w�|�멣�/Cf]Bl��$`]�B���6n}N����}����3z1s},�$�׵��OgwWz6�̡ٱ���?��׆�5�㫾_�u^�="��wj�t��:��񷳦�0k��0�s��.���'�;��A��-�O׹�=|�2x˧]Og���ާ=mq�r��ԟIxk��ޫ�-�2�U�9[+�GK��{�*���g���=t�Ri�%;�t�ϡ������+�yk}�b�h�<0�k	�?*}C2*0���rVCk�*�
>U鏏��z]��p=Bw&vc��ɗ�]��*�\t�]��\޺)};�o3��}�ó�U�6z��%lo�|�+eR����-�}^`���G��{0�y݌�`� ���^ԕ��I�"�B����ז3�{/f�+G�[I���\U6�n3�WZ��:�l�&�r�E� ������T�ͱ��;�]g�z�NQ�;�	9w�[�s���fo�Q�*7�.�
�H�8�g���q�2*�5�1"{�?W�y+������?|�R�l�}��ޖ=.�ͯW<1�l����^�3��AC���
V�ח:�Je���J9��Jf�f�r�EK9��Hܔ([�k���Ck�>}�A���Þ�����ę�;��;�yM�J8����k�0��+��� W�k��˲X������gMܨ�L�����������Zݽ�ʊ�_\�YS���g:Z���jg�dd���ea�}�7V�O=$�8�y��p��M�k�o|b��X�;�Fׇ�[��/ޏ]�}��9P�����~��T�:���%�y�X���/@-��|,�{����j�,�2�IS�刽�c`��}��W
;�_ڷ��AOz:�X�N���2/7_{�޿���y���`\����
���fR���߳64l<OԪ���'f��z]>z��rK9���,�U�"nhŌum�[��BRXS��*�Fm7ŝs2�r[������yfq��r�-
��O��W �i'�ܘ֬����݌]7�@�lQc\�t� �.��\[u� ��[Pd�\�˴��=�ڪ�(u�Dj�6n���FQ\z�f&�=����Ɨ?{����T�Կv~�V=��5����_�z��U��g�,����4Pn�<~��3�fsl�{��X�=E�����A�b�ufE_lì���s:8)�=�;z���y��E�]���_�����&w��O&]g�U�b1��
�^�:'oDG������;���Q�R���#^fz�U�=��ٌS��mb�-M�v\�ޤ\�DW����oؘ��J��fz��y���b��
5�a�+�:�KJ�<�f�����,�o:Z�����!��'E~�%d���۪����,�$����]��^5Æq�ߧy�$���Z}X=٪j��z�6��t�W�����L>`gq�j�}�r��Cp7}�sN�zkϼ12-�{Ѷ���^���xdͪ�,��uﳝ/�l[%;�I�û=�y���>�Q^�H�󛾩~��ʅv�;^x���}%�^K��B���5M�i���$`�N[O��W�����9��7�Ҕ��U��7t�l^MAT�	N��3��(����ji^�7:���lK
o�潳��_sֻe�}p�29mS�uc\�O3@ v���m+U�mb[è^lE�������C�}@��轂�Y������.���g]I&���cφ��R�;�o)�xz^G���X���l��w�����{͉��l�� :��g�Iď&���Az^�w�7"8����c�ޗ7~���
8�)3V���{с���ڤ^�Bm*��fV8�ﯡ�O�MG�j�{��{�w�W���?x�Pw��s������\�u^��~����f��A9��]�M�9��:>���#����o��J�u'�t<��V��3�Iqz����N�U���`7������X=b&��u��E�S;7c�X�f`����Y�����Cz�q�x/��F$�u�רδ����<���?����;��G[���Z�=���;!��(���}WQ�v?9/���^���|����Vؕ�=-�[�)�z/k�\��ս틝u��l�?��ڂ��c����MߦⒷ\㩷[�Vl�K��E6� @����3��I<��T}��c�S=�@�q ����M6y
娯�b���vC]O3�8`���
y���D9ǮW"���Wه�5{;R�#{M���_�������J���(��sĪ�3��������<��=uŏULV6Q;=6b`z�3�y�z�h�粮���z=I:�r�TT�c�������nk��R��n��e���Yl���sV}�nϧ���y�ʍ�y�Y`Eϋ��8���y]H�K;F=��7���N���=4V��9�3S6 ܧ&xeT�ON�<��/�B�z�\WO!R�|��*���֘Q#؄��X/��K�mrk�Pp�%�KO�&I�+"w�y���w�	���������o!�����)}���m0��Q�t�h�ĺ��¥���v��Ζ��C�夗�Υ��.�=iക�2�VEL?��w+��1{84�1�5}��/g�:oHa�z=])i2�UH��Ԡ7c��ǭ���W�	O��̉��:Zmڰ�����j�����X�V�/������	;(`կW��>XV���
�g�����QY�8x��PT��0�V<쥔��A� �%$��>��OO{խP��s:���5l^��-Ԝ!gzkY�&������Ȃn�G��Ԕ��Q�2!a���Ӎ����r]H��ү��1�\����)�r6�Zܽ�	��L���[φ��(1Е�vd=�]���w@��v����t��2�~��*w�z�����.g�b'f�7~YXK�`o�X��Jy�"���!�n]�F |��o9������B(�b�V��؉�������@�{a��U"��������k��K:�gL�ޠ�6�Q��&O_Ą4:==lؤ&!G^�;��g������]�J�6vzv�	�3�DS~9t%s{��鄺c���a�PW��n����u�le��0T�d��i�s���@"���>��U��bz����e*bs�cD��	N�ؕ��ip�rouy@�����}"r�=�z�Q"x����ҁ[P ���Fr��ߦ�O]B�7*�O�$^���{{����K�X�J�/�j���S�YAC�r�L�?K����P�i7S��^�o�D���Y��l�$��sx/���{V*д�b�����	�:z�2k��s�i�B�=�ҳow�X�,�@9y���Dߐw�_]�d	ؘ^\�\ka���x���ʲM���|��9׍�+/��r*��v�|�G,n|:��,��ʣ�`<�
0�0����M���%��
�s�����z;y��CJ>��O{��u�S�$�p�W����7c�=��+�[iÂ�V���V��熬6�0��&յWcx%����̈́�dI��j�C�EE[9�F�)9�c[;���
�U�wt�=R����@#�4�Y�ъ����1��w�!j�~�m?]Q��^�v	�������PۗO9eY�Ͼ�jOu��/4�!��9�J�f���p��/�.rb:�ތ���Z�L~n �j�i������ ��񪙞�j���L���X�ڜ���LU㝔��^�4�y) �$8˶��̇ms3����l��zD�W��d;u��O��r�9�
��mt̆�MD��cN\�sot���N'r���u��j%�V�B���W��1Å�}�Ý�Z�n���P���^������`��	�R�^S�JL4�+��,3�?O;``���[���շ��r�t�1fx���.���TZ�%k�E�Jı��N�K��M`��<;b��wq�z����]w����\�������"�n	;+}It��v�M�8�y�t��VW�O����t��Rd@W��,v�X��Q�^���a*���Zp����>���Y�!�����?�װ��R��_����b{R����,@��D;MZ�3VG�:��[c
�)V,�WJN�������i�Oq���tfE{r��ʃj�Ĕ3�6둜k�Ϧh�Wv�6J�2��1�]0¢�t;8��7fc���l���H�΅L����poe#S��o ��F�1�3&�_)]�B8����Bt�t(��vWJ�մ�X��RaӨ�����gV�L;;d�±�t��ec��j�t�R;;pU�ݣ�im��].�T����2�lLn����C;y�n�S���t����ڒ��^m��n�ӆ�m�-��4M��h����[XZ.��n�|.��NXT6b<���\��q=��n�!{�f]CF�B��%-궩Cu��Up�W5];v�B{K�_,�����U�W\�2�_^G@�A2Z�'* S�«��]�k6�m/�-��Y|��p��9�[S�f__Z�*������F�����X�l)����yH���j$�Yk��������MQ��d�=%�]I��n�'�,v�cچ�5�ǃ42����Z˹���m�ȕ,�q0��.��۹ �FVa�]�d6���m8q��Г��GtL���S��z&�R@el߃iQ콺��|U'�ʻ1T}��	oTYf����w\���Q���Z�>��-Q7X�#=o&
]-|��}�O��Z}]�H���v�L$V�ݻ`��7���7�\kL�u��YJo1�E�����Z����.�jX�ɮu[ϴv�T���¦YOb��:�9p��Rаq����/'U��!�R������A�~S������K�U�ޱ��k.�p���;�9��l�4jd�{���ʻ�o��%��YB7O�r�ϖn�x!�]�t0�J�-񦕮0�/{	1��ڬ+-�W�n����=�Ɖ{�(I�i��p;T�Ɠh�,nFAO��zw��WljU+#�ΟGR`�P����v��-�J2�whKg1R� �n�r.�if�����(�I��� �՘�e
�s��˗C�˺��2� �'�Qܰ�f���Փ7n�Hi��6��w��&�� Q���vGX�e۶���L���B�2ѶL�:Bq�3Ὓd�w
c\�Xm|�w��5]��SM����d?=��ׅ������g=`RW�V-���xn�%*�e��ni�ɛX	;�d)���B��c0�Ύ�>�9^�����^�
��ʄ�sN%�E�:�t���޴@o/7	ӊ�MRV.�h����]w.��à4+3�᳎&�?���2�%�J�[$�7���	��d=��DU���ԻY�;,�T9��0�8�ū���A�S5df���B�����Y-��˰Q�ڣ�#�u��v�*f����M�F���b��|s��8W�F��g�q�Ec����p��k���5F�l��+ �s�bջZq��U�Es���r�\1�4�����F��:�W�L)�̨�s1�K�r���>DA����DQ#���U��Q�X�QUR1U\�Db
DDU�E��̨,`�DYDDDX��-��F0H��!DĭB�QDkU����"-�Q�����Q���X�A��b"e��"DPDX�DQ@�QAD����",+b���*�iTUQ`���R*��Dbŋ��+X#QF
�1EPFZQQ�Qb5*�����"(����QT�(��mX+
 �1EX���lQTQ��b�1�(����PDEX,Kh���E�j�*(�PTX�F((�9mj�A
�-(��Y`"ȶ�T`��*"��Q���+H*��TE"�PEE"�"�X��DTEUJ�Q�b�DTEQ+-�A�b,UT���QPPUdEc"��������PL�ETTb(��DH��T��TDTD��2�Ub�X,����V1T�TK-d�9�D�ސ�;O�o�LY'���>��e"����e���=FZ��0����}z���vwEf�}��]��F��폎����v|"te&�y1:���J�.��D�<�F�j��i�m�yOW9���w������{P�/.�`jjX��ST7乜��ނ�]c�;_v�:��7]�S��g��TuC�����j����u�%��{hp:3��(dY���pŕw�e^f���^+=�4�c)�b�92�������p��Y�7e���\>ڹ�	W�A���3[�JW�,2�;�~���d�_s�/�I.q�j�s�Pcjv}�}��7���p��/yADE�s���m�Y^Q�91*��aO�$��m�Η������b[k�	T�tePh��K��uʌu���sW8�ƴ/�ۮ�_^��W3��I����Pt�������Ick_b�갱�lA'�V5�39k;�*.�$��M�I�G�ъ����".Ά�{�Pn�>L):���<7A3�x��Σ�=�������4界'�;�+��훖�7%d���#J�2��0o�aب�ܐ�<�0m{��-cz4.��9�Y1>���q��%������E�e�u�>���>N�m�ew���S ��`_#YLc�7+&6{vdڎ랋n��dS�8�:��X�s����p�L�d�� U� }�W��VNC��4�j��Ԕ��X���wϳ}8�����C��K�-��u(p	ȱv2e+���q1���\�����[��Y��R���hs��L :9�DĿ����9ᔮ��0�¤6�&����γ��+m��z
4�gN/��9u�/�BW�e��ѷ��K<{w	�8+�*�C�_N���vH�e�;(����Zl5��}��ǉك|���
*��f�KXəy�y�~Ӛ�	S�r�\�RN�x,4��Xb�&��8u8��IWy�������y�7�P�����ssB�Gz���ˁMep��1��)�e����2*�����WZ���*���\r,��O1e���X$��{����.|]�q��F��Y�k�tq	N��BP�h���a�)�3�lA�NL�ɪ��y��_�Z=�A��!�1�\�n�������O�^���\�K��e��I�+QX�����G�n��Ʈ���p.���Jr����Ƌ�6���Kօ*��4��
�zD�5���4-�Q����u��N�.�Ze��^�N�����ߏ/5����~i�g�zћV�39�襮���%]b���X�e��5������3�iL���凍��{�!qA5���s���WWK?	����Y���j��o���?���1���U���~���"�(s��1d�WPuG�]vW�<�Jęm"�U�H[�3#��Q�{��sؽ��:}�]�}]�ZL��UH��u(:��.���4�+���!�>����y�%�YbyE�2���Ѣ����AZ����G;��@������t�(|���x�;�eY5N���TxX[\E��֝���X�6z�+��Q2X�����N9Ϻ���"��K��T2r�5�l��daitO}r�QU��HӃ���;�;�1�zN�!�[}yv���x�/�X�+_)yD�05�T_�j^��6����?e�G��ȹI&�0}C�8є�����%�!N��O��	�� �u4]l^%m[�b�x�<�陞�1��8O:"�Hr�\�|�����7��6+)5]f�5�B�eI����gs���V���"W& <��*8nr�*���k�-�%;�e%b�ݓȿ;d���{60�Gpμ�`�ﴺ_�(� 
9~ru�,U�߼1[r�AW��Y�vY�JTa�]�X�xk�������R錦�u
���s(h�m����Pڻ6��,�Ѱ�=�35�9������r�t���	�l=I�C,F_h7+B��Kq��6G�$�9��3��]/���Xt�E��\��n��uϗ,;?}T$��ž��D�[��?<�;UOqOMg�C�q�ͿK������`5�z��d��u�q%��k���x�q��C|�.�3O��'��0�hZf�Y�=��P��=^
`&��?:n�e��p�x��N����x�ƞ<y��v&W�2�ƶ��{�f?=�rN�W�b:�izi�='z�fX����Es+|�^��PxH����X�5�{I���G1f�Q�W(cW\�)^>�E�Z�`��I�O�����.�r�x��9R�^��~�N��V�r�yex��sW�/	[)x�L0I�J�CUA@��=�~������S�K$^Â]&�5F|=����E�M�㕱$?�RM�H���������%���&��o�U��|���0��Ѵy̯y�Ί>�t̆��58�q�V��g.��Ɲ#�����{I/�Z��g�}������{h*G�0p�FM�Pt�����{x�������JL����W�E=j����l�,0����0ܻ��wu��@ئ��;�^DՔ�VH�\�����)9�r���]�**Т��2���nS�s�w���S$1e@;7q���n=i�6�٫3���Jw����>�R��+��i�*���V��M����T<���ާ����_ꠘ�V������D����n�UY�'Xiz�S�<F���un9~֝'�Uu��K�~|O�� �A��|Dk�G*��cjN��)������������T�X0X���o�2�F�T�{]�=��FE^R�,���=yQ�O0�\}��]]*���R�ߡ��*ڦo�BblԘ������3V�u��vb)�?kd���2B�m�CN��������!5c+L�L��,.�qu�[���̽'z�C=��X=I�=�9!T�Հ54��ɀ�M0gܗ2��-�]Z��@�3�W�����s�����g�9"��[������*%�\/�}g(N�ۧC{��e�S�S��#�^�x� ����i0��Lý#��A-�r�W-9q7�Ѭg^��<%��~�rR�Q���\g���g8W�=��W[��yG�I�x%�Q\}Vy��9��y��Ǚ�E{�,6.V�ب���;�ΙY�M�K+�3t��P�d�ij�ZZ�V}p�PV,�{�����f>��bL"�>=�0i�u�6M�ǈs8��+t��T�^VhX��s=׈�76�mYmY��kY銵R&l��j��5�]2N��7�'Ȅv(3�6WJ��sW�,Wն�p]�5����զ�V���Rʹ�&tm�����;����}�C�aє3�K����r����Y�.�5t��4�3�/��5Ԟ�����W`��"T�c>7Y�%�:�1ˀV��X �����>��yt\��<,��Ht��yj<$4!��
�W���tdyCu�=�������.�r��`x�5w�|yt=�5\�NfA�pN�,�@u�1�U�ԥ��s*v�u��:��Σ)�g�m&��O��e]�:�%��Q~�"8�7�C�=~�γ�Y�n3sV�%��1e@�`�J��6z%�����bZ�|�w��ɸ�Ч�}9����8Bib.�WTv<�d;�[���\��T�%����h;V�?.��:g�R���4�G�KdN�%1���`ᖦ��8�S��eV҉
Lzkk��y;dX��`�`'�V�h����<l�?�xt�PP��ҷ���m.'����CF����7
N���̧�����ʿ�����IN<
j��ӽu�)�UT�ښ�����	��F�����U��z�WU�'�n
�Ys�i[�V.`� GlKF+\��x
<�P��q�wW���pH8m�$�&+��y0( �n�m$r�E�l�g�;�2� b�K�FwPcw�fQk��e���V\��O�������.7"��].�`���u�W���\r,��=�O1e�3�uH�Unҋ/��s7Y�m;���ļ�*ƣ���p:���[/Y�*����_��{UM:#��Ɲ�Y����F�շe�A��K]e�� +���*�yB�=���ɶ��X&Ur����o8q�g���si�Z�D3��$�Z�&W�cDI\:�%�B�w�e��WF�k�~u�Y��]�3���м�3�kEș&댺t3�����g�+4Gȩ��3��iY��<lpǒlB+8���h�]Eیz�R�^�:��Jv:;\y�9�+�}�VK��(�{x��;��7\�w]�����FC�M/��8#����k�BN�cjf�Xx����v�|�KG,��S�7fv�~ɪ펺�Lqaf���l�Z%rbAD�͑��F�#���Z��^���ã)��� :��Z��0��D��\�3��!�2ymm���2w�����=�����Z��uAa~9g�����P�贞Ϩ�X�3��an�w����\X�v��eu>7u���H��[M�MIY�fA�]��`�C��	C�܌�Ē�2j��K�e:��)���vV<�*	/��	�f�&��݁��8�s��}����	��#N໏}O[���Z��r����+��I��{�*5�<ӵ��+�h���MY/	h����	�p�X��N�Ay1nz�ȳ^k}(��/�J��Z����w�,�5���8����j�
�O5��;#��)7�NIv.��_�� �����e*s�:�UV�X0s7p�W���}o��6L��p�TC3�rc�=i��@x���}P�S���N���5z�tN���<T�����Ip��[���	�֯�j��➚�
A�8>^�}~��^����"�{���� �M�'g"��/}�zq�i=��U�i��gܓؼ �8=����v�����q��Gla�I�za��h��ndM��x�,@N�[Ǚ�ƶ�-��C}����e�%�zR��w�)1s�w��	l�\���	NX�j���X1�B���5�s���&���n�a�Us,ŢC��Ꞹ	�f����U�P�Om]�Y�p��ף�r=��({l����nu�=�(�<X��}�vk�F�<4x�$$�;x�'v�d�Y���]A��R)WR}�˞�����y�j�m>|쭬L.9�S:�.p1�9�X��K��V����:�;�� ����C&spd���⨇�{�Y�l��W�<x��|�F�i��5sٰ$le�{�y��9ԥNs���:'�-�T�g��To�AJ,���ٷ�w&�{���u���7�Ɂ|�-�i&���l��nP����q!�����談_֬y��]h���Y���8�Q2E=;'x���{�A�4�sj�W��1�TO�C����t�ۯ��z���`��1`w�W��F�W�6GJs3�m��\�	�B��Q�:,R�ح��F-����ģ�%L�xEn���=u
��j��F#b�ĵr`ȼK�z];K��i]��*�W����j�<F�2��2'%R���A����]{V6{�Al��;y��8�e̷@����%��V^,�G��-<��@W��,v�X�B�?YZ�q'���N�:�[�BUuJ<,yz<�֡�kv^�1�u-�T��]�}6���Y���.t;��;0�FCc���ly:.�V]V8=�p�j%^Zg�-l�|�ܖ�6���o6<o4<>�vX����X��'=�#X~���4��`*���H�t�����}%�tVd��׼�L[|�$!wrr�p�ٜ��F��K��ZxMo��/�/%�T���V8��\FK�q�l�:���o� �^Z��������z�U��%9f�6��؝B�N�Ԣ�I���l��B�:)Po���>�\/
��{3��T�:_�����ǵ)�FN�R�����x�d3q��回wޗJ�����[��J2�V �S�*���2��g����%���^t��nG*�
�ya���@�9���ݣ�?G<�Kp��;|�:����ܒk<��8li
��"�(�W�+<[j��(�ӝlHp�]��No�=�����Ʈ��gx�'�B����E"e�O���r0pa�zK��]<��3�)\�zzGT�[w�C�K��A�u^N�O�ˀV��X �X�t�:Kϭw�HO��;����z�x���-k�D^(��e0|���>�����%�O�}�'<�а��=�~E��x�<�@�w  ����$U�t���Uq+w$+ԭ��k�2�`XXc�h%֖X4=ɟ5�J��K�� ����u+��#鱱9i���~.��V�J��M��]��K���蘖���>Ԋv,ۓm��yD�V%B�R�:�n�XF���0n�J9O8-�J��S�Vws���OKS]�XIS
�f� `ŦL�x
�=�s$�����մ��dʾW*�y�.P��o���y���}at�t7`�8�IJ�m��$]�:�ï&�S�7*T(��ݖx8o+w3�dU�HQ5zv�3Uo^��8����[R3.��e[���=tݚ���lZ&�D-V�:,s��!9��%fPLQp�u��n���Σ��W+3�������F+�JgFz5�B��u��[�'�ɶ�SI	&��腩̽ooG��r��I�O<���gdL��3&=�2�ƻng�%{�wő��w� �G*lz
�$�hk��j�ohr�o�_����ڇ�[�9�0�$�m(�3:�g=���҈8��`�a�8�'*��n�o=��c�)U�ejw��*�nA)����S� ً�˲���d"��
ȻY���n1���t!)89�X��©��txk	W#w�*���8�Tg��˥oj�@,�C���X�W�&v�
f�Ako�k��5��e�ˊ�+���2�X�U�!���h��Z!<:	Wn�lm�B�Uv^`镕d�{	<�k�Zo%k4/�]h��S�d�OjXl8&k�v�Էz��4�i�g��m���R�s�ʊh/J�%��v��P�d�˰3k]��w��9�^䱥dP��,���u-��%�ĊG!��.�R*�U���7����n-=W�&�w�`)FU�Jd���VBK��R��KY݆��t�놅4p�oE�����-�#를s��:��K�w[ˌǊ^�Y���霣̊4�-o[�5�H[5�n�0,�����]薹�Gm��	��ݙ ���X�^E��M�R�ޜ�M�6n������W�Uvl!u �����5����}��k���!�C���['P�<���ub9���6��˵�y2�oFr��_&\n�'[}:WIǛ��wK���f���Z�O4�����l˸��,մ��EӮUcIy��@�tf���Op�}�9̐��Z.�����^+�c�c
�ڹ>{ۃ2���J� I��C�x5�R;x��`e��;qLF�htD�))�]��"P@}�M�Y��Ehя���8+��K����G�@�RM*÷���k�q����I��tHv� �0+���T�a����������9g��U��3��ȡ���6;.�!�{��􌶕5F�?37_;«WY�����1#5��R|�68uu U���k�F8��ij*��O*�.�>=%����|qc���+��[��V���Oc�葌J��Cʏ����;�v颴d�����;)�^̼X�*U�E]���,����8t�U�ϫ�*���J�*���ލk��	@�*`Yv{X%���o�t��E�����gs��:3e�X�L� �7XΎ��t�g;ӧQצ�ؒ3�dʍ�/v̘T )*Db�(�T���#X�0UQ��"�U���ETDUc#�EEcdV�`�,aZ(*����ڊ�mZ�T�QUF*0b�҅b}qU�bB�U��E2�QX�P� ��
��QE��LB���`�,V*�����TD����TEX�#5�kT�UJ��E�D����QW���"eX��TQ�UUUm�,Q+b�2""����X��	Yb(��q
(V��*Z$F"�$QUDT`����TV$b���8ʨ��1��1�b����,TPTQ@U��*�� ��X(1Q��QDEQT���",QU`�"�e�2##1X**�kD������f5X�-(�"�ŋ"��(�"�Q ��,EHx��ˍ_r���1- �2��SOi$��˶ɹ�pGPd��k��|���67��m�\e�+&K�G��n�_^oJ#i�G�ԣdAuD��)ƭlxo�u����/�樿!�϶#�_%����u`�`����C�U�Ȑ��"w�V>�F���Xί+��ļ'`="e���{\�ú�U��2�s�r�_�ԕ@������gԪ��y�N��˿x�w���-�綽�|Ҟ9�h�N����*�9��z��I\����N�և:A����%�+��N��N�m�9)}�dۮ�)��JC�q�{�f���5H�UOy�Y�e���g ��Ξ~7i,�Ōg����L4w헬��!�ɞ5Sӣޕ�g��U��9��9�+-_���ᾡ¼�gþx��uX�
�]jo�'�H��V=�3L������;��ܰ4!><�F��$�-c;M��VE���zХVz\�Ͻq��SԆ�X̓��D)t�}��oˇ�u�|���.�$ǔc�������X�a��<EGr���/.̭����A��xy�<ʟyk3(��Õn1��KIy��1B?'R���ˣÔ�@�e?S�ŧ4����=�WQ��E�&e^����4����4M]�Xp�.�,�獹�0�}s��F��L�{�!�����ޥ*�uL�^�5�|����:mX���Q���]��Z��gvA�̔��<iI��͝�:�ۚ�E�m��3���,��x�]��',�����Νtl�'��AZ����H�.�����|�ރ����ע�ܡZ�z�9g�	j<�8�V6��7X�r�R��O,�E1��scw���"�=����lZq��걈��6X�c�S����y���B�DH�{ɍ�{s�E05��摒�2|��"�X�ʡl��]��(]tZO{��{R�6c�͐Zw���O2�z��2ߑ<Q3�"ϋ
答D�(��ю%�Df�����^�ʇ-;��{%q`J}tD����'=�W�*v�g֔�a��c�ed����FU���2��^֒>ր�� >�� �ʎs�ȫ�;�1�$�qG"y̮9���o�(]k��LC��؞;c�$f-0���CO�H�
3����w���J�D5m��GgЦB��`�}����O+�zk���2�O�� ����n���>����<7
�ZK�D,�f����ќT>%�ڠ5�{�֫+�{��̃�Bţ�3�i����v�y�K�_"g!�]�8�ޢ�u���%e65�sk�)�sru��a�,��@e<���~9@��%�n�Y�ij��nD�E٫2�gEs�ql�z�]�Pz�.u��$�N�kz8��j�+1nn��$s��W\��1�Q���3F�s���r��e"��v
��]Ô��u��a� hƽN�V=��=�*����iF{ԝ���!�.�I��o���f+��κ{��{�)�y�5���V�)3݁)Z�=�0=w��5x9�SR؁��-�\���YCTU�w����bw�H�Y����Y�gՅC���B���������gJZʥ�ǧu.�����q�k[Vi�ꨩ{[J�,�68���V��K��}6��U�<̮tw�;u��φfs�2C�T�2���Ş��~6��;ƒ���V�]�����<��rd]�cb��N��M���� �A���D�'>���AY�B�v�w���krz�&bO��,Ë�ˠ�O��a
����,�	�զ�3�,b:&����;*�1nl~�h^�>0>!��A1-�Ar]�^X�_˓E�^Jĺ�t�_V�Fݭۥ��fN+�8�}u֝"�!���t���k�5��
*�����eE�9��*ȧ���#��էG_��3�7de�%D��RH��Iً��{9�+���:/h;��V,�ౖz��Ls;��O��S�����H��M{�3#��諫j܆bQ�e�Cn���M�s�G�1|��8�iQ��Ơr-ꃭEٲ�(�y� Ա����7���.z�/��
�RG�]���M�U��`��P���(JrN�R��e��l	S:<����E��u+�\�x��-f�R�T,x�E�2l����/MT��Ԛ�.�Y�y���(��XV���zߌ<�X�Ɗ9��Sy9�'@�����C�d���'�]+�G�'��B��UN�f�'���m��{'�tVj��\Z^��D�i}��X�}S��M{�[��y'^��a�%��>8������={�ڄ�X�P��]C�7��PA����pt��oG�{�o|�,+������k[<탓cfj������W
���|�{�,g?EW�T2+�o�~Q���K�o�߶v�O%���%Yv� ���
n<��|��P�;:]_��hV)%t~|b����v�����ѝ�y�:��E��F�&ٗ �ˡ��h�7�K�-�9�`�ÿIu��o�=y�Xn�{���79AX$�E{알��"�o讥]]	ˮi�U��p�4ۖ��z���0��J�R���U�n'�S��^����@=���l�G���D{�=ͻ9��8ܕ�� ����s��������g���i��c����e_M��t[7�xyC���W`b�:�#�Ҳ6�&A���S�	m�I�n��3=��Mx�pV�c'����22�ּnA@��� �XL&�`�>󚲖r;h��
��G(��ms���u���SP��s�G���8VI���$Y^H�'��i�zR/}W)K��K�^����A)ie�C�g�T8�ߡ9�}޾齾��\w��vD��7���V̡�+:VD����%���EBt��K8�]���j���)Q��W^m7�HQ��<��lzm�o-�����5G�����������y��	Nx���i���v��a)���#M���0�/u�Ⴐ���˽��\�o1z�IW&U]�.z,�V'=��x�S�$��0 �|)�91WPʖ�N`X�nז�r]�>�ٟKC��X��nh^�;Ԕ�⫫���QVDY��
���n���)��҆=U=�=9֠�}:��U�����^��2�w@p�
#5���!�[�(������3�MAC��(S�G6^���3��b�t��vȕ	���g�cW�\ʲ��\��=Þv�a:��������XB��KP��i�/L�L[2r��+[��/z��	m!{��862��f�7�_m%g�^7���rp�������Nۼ�����G!�ޓ���VU���U��M�5��;O	S=z��B��)�-u�%���+�t��K��]
�3z߻�c�~�-��_'���:Zd����3�D�^8%��U�d����ș�����8-d݉�sg�)F��t�h��fe1Z�W���xEN���y]꘯�cu�Iv�;h�]�5���<�A�(�w*�x�eeyk3(��Ñv��KIw�8��Jc�;���z��ǃ���3;�$�c�EZ�P]�*u3�j�_�Z��τ�l�ޔ������M9"ڏ�{��b�t,������l�σ c��bmR�4ePV���u�7)e/K��}W~nI[�sT�����X��
'}c$Wř�¶,4�׆"w��cXLCM���ɋU��w��ɾ��-�߹����r��D%$d��'��E�]��W�^Q;�[~��Rb����d����Ժ���1,IOb+��+����H��¹�f�!12ǃ�p��'�N�Ԥ��"tO�V��4�W�P��.u�e�;ؖ&�)�У�fՑ~�����Q�[�u,�[�k�Ka�=�\-sh�>��Ҹ�f��7�M�8�VF��8st��"�f+ΉB	5EW�lͫ����}�&>��$��7��Y(��c�V�1'-����ئ!���3�8�vP�n�r�]r��'9؆v��HYxq�8emi
�桫C������D�|� ���r��\��*���k�c��c��E'�ӻ���Բ���!�����lu���ƨRs�i�BMOG�%�3wb����ގW����=e�V�����`�}���U�O+�zk((���+a�W>$;��N��:�sD����C*EZL�D,�o�ܵ���\ZK�P�Z%�%�|7f4g��d�>%��Q�ّ���Y�O*V|�E-��߈����&�������&u넂��1�bs_)��������/ԝ�ʑ.d�����|�Fb�NX�����bߪcS��4y	V�P}���'���PQ�|���}MKb��=ptͱ�]ZNX���<M��>O�Bܭ�P��h�'ྡྷ3�����?/g�Y^_Fmζ'�w���-ø�{7Q7C����~�	)��O�Tǳ��I�VZY�{��Vej�-��]d�G1`���Kٗu�I�ޟO!�ßzRLH0S��Ҿ~8�w+	'�Z2�9�ﾨiP�LұW�o��}*�[���t]�;�ӈspqk�w�E��(o����J������d��r��� ��۽�v0�����`}���p�5�ɮ|��V�;�s&'��0������VA��K���Ư��xò�o*��N�6&Dv�e��ʂ���orN��?)ҼBu�w�45��L����P�D���t����9���7���c��+u�3��9��0y˶��X^U�rE�ɡPf�;g���{K۝�8�:ZYVחNe@�_s�Y<y��ژR���k��E=R]��yb$x�[]�KF�zWu��@��|��}k���^z���+>�����0GD���^؜7�TV#:��-�q�o�_0:�݂˔���9��^�B���x���[��p2���W��"q��I��N63�7��׻=A�dH����(f�R��Ǟ=���^��er��W��Dx4�{�vw����ӻ�S�1]%�*6'��&"���<;fQպ������3j�ac��A�T���i���KnY�����b�:��+�')tř���AJ�g�,-
��\x�1���Ƒ������.g)���S�bq�N��5��o7����/�p���]�R��g4�+*��.�l���>D{��r�PA�M+o�ɞ�;�[�U:�]hز�
���~��`<m�
��gH��촶�n�æ��;gw�+��cZ{�S-7K6��I�\3�+��ټ�Ζ64�ǥN������֌D;��\����dsy��0��@��C[�J��� ���j+$�#�Ykv�ΑX�(o�q�\~t7N̯s�^wЦ`��2��\e���}�t��5������y��xo��.Ss�0�0���G����]g�mR�E�����;[�b�J�9
�.��t䉒X��]G�m�����ͻ�v�K&_ww��j��l^�wT�4���,gj+�cB�y���BF�.��֗�%��C˅b�s�;�䔭G����8X�}�ntp�G)i�(��yL#'0$�j�Ո�]�u������.�y�;?F+�k�M�(C���7%d��	&J�st���У��	-&���>ͰԯM����x���JZ^���\��T��'�1U�uN�#�7;vx���r>�P�6����\|����<��X5+��8f%<��ݻ���zKNG��ǝ���|`{;U�8��3�i��c>[/B���~�|&}ˬ����L�s7�٭�-o�meT>��eQ�Ϧ-4���ȝ凞c���,�<�޷�e���؞%�.Y�0�ӻ��r`&#��_S}ܟV؛ f>h2����2�wI��MІoTM�.>Ȥ�ђ����Y�螣�1)�N��.NR��jn��Y�Iof�`��șAbOk�t�{���g����� ��;yJ2j���y�M�(�j W9�t9t�;ԕ�c��~2�`��jt��3�:򤉹�]FuZ��I�ʮ����>/%������%s���P劽��#��ɛĐ�+���Fa>?:ɷO8��:���U��*y�4�TfT���dEV�M�3Ӛ��>.�8�ۨA�AU��Ŭ�����-��T�}ٽ:mv�� ��"��G����E�֏T+������
�&��/�Ob�Ffv\��$��;�g��-�+����d��<_�#�i��u�&9k�"n/��ŏ(�6��y��#�_s�n��X�Y���>�M���ϙ�LV�Uêbd��2�������vׅ�?p=���2�dcq�8{<��W�a�| ��Ϣ��:Q�/p��+�@�ʺ��z�u���1��gQ��(.��
����',����gNtx�'� X�=������[{���b� 
\k �#졃V�^���xX���yAX2��/뗷K+������t�����������2�<�4��o�r��0K�^P������]�ػ#�Q5���%ӳ(�y�q�4%o�z�8B╒�����h�y;(q'Q�\��-4L���*�,\��SUC&٣I�}Zsm�I�"eo�����ڳ�ۑp��[�t��GS��n)|o%�M`��o@����:tŁ��}	�Q�k2�*���[GF�L^!�ޅDf<K��]���� �!ר';������+0��&�k }�d�S���K�$4c��,!�$�+UcJ���3���{qv>�K	vn�7�Y��*�;Q����w�׶��D�T�L�k��1�Z-+M	�kIn9D�ֲ��oqެu�'u�ɘ c]��E	� ��[۷���f
�5�t���0���v����9�:}���U��å��p�	չ�C3���\�tw$�-��v��m>����[�����]�c��޴�r�"'�ͬ\&��ܥ�n�8ICV�Tl�[͂�ݩ�5��m�����:�JMvӭ|�$i�O4ʭ�{�g.�n. m��ި��+�o�i��NVd���Ѵ�DV��{�ܹ�3��Ղ�`��)�;D.������K����=ʺ�l��\�6���#��=�$��:��9W����I]��)�e��
��Nڮ��Z��˷��V�JoLg�iN�+�1e�&���XA��y�rb���ř���S�S��`��n�2���o{�a|��I:�z)�_�dO-`�Gs6��؍�"�Ce*弆XpsA�-��P[�-�X�eq��/o�T�B&*���u��5�Q����/A�#���|��"�7�b3K]G`)'���k�,��כ�y��|�	�б%;�R��Xn�*6�:Վ�<��#�al\�a�.�ѳ_Swr��^�4���f�C&��Ф P����
Q7z����
��pƨ�SHwt�"��)VhY����3��Z��_G2��k�J^+�i�[�Cl�:�M�ʃ"WvI:�;���GYt�>���s��{]gJ|�߲�I�E͡K�k���)
������;̻����G��n�F��{q��oOff�)
��M��G���2�5;�a�7/D}֮����B	����\�����&���Ut4>�� -<:VrҼօ�Z��pE�z�^+�O���Jɛ�9M���� �%_8�L�B��M�S�3, W$�'\�90L8��T�r�s}�����J��Cb4��
��_�MJ�t�:ف�w�I1:BZ%�wN��y��D5�[I0��NoH�>[e&eiq����nH���{��M��:���F�z�\��vX.�uӰ�����m��؂�Ɔ��-v#�B�G��N���5��2�b,v�贯r�Ed3�V_C�&m��;�� DDQb��`")��V*�,F(1�DcX"���PEb�PE��EX�-�Db#b���"�,r��j#EU�2,Dt�U��E����D4�(bJ$b
�2�b�����DUV1Q"���
���(,dH�b�(����S)DdUTU)��PDU")�WT*
1�*.61H(��`���Ŋ:h��T��2�DX�U(�E7(X,QX��bb��@�TD5J�TT`�TQ"���EEL��������-�(8�DF"�DAEU"��q(�Z3#��Q��VETQ¬"�jT*�� �)�",DDE��EQKL�������b�|�2U��Ȝ��fݮ��Q�&�,p���o�ÍN�{uܰ���9�[�й>�s�T��@��bm��̠�8�<@,�:@I�x����\+aШc�7�+l�Z87)J�&j�>�� �w�5ʳ٫�VcH�bd���E�u�a_)���ky�`��ܽ�]:�]� �TK���LK���
�J멥&
E�G'e�*a�$w���nv�4%YA���^/v�&6TJ���y�aO5���KX~���S
�wɿ/
���s3��/W����j�<9T�GխӸ *�L�*8D别Y���k�\�~�tz�Y`�S��)�{>JblyLO��Fbj��'Ρ��	���A{���<�]��:�Q�$_�vS+Ge	Kt������T������Q���8�9ƍw�Px�ރ���=�?���ʅ�҆F�I��d/g�?y;[�~X�j]cj�i�k�'�O/��nʄe�ڪU4�����zxѿ(�w�pw.��m5�̂�}\x�+�y�M���^�|��y��T�-�[ J�5�o���Չ�JCL]T�=��-� �/��JrƳ��{����u�n��ҵ��ʷ�s�Z��2Zր�I�Vc]\t଻��U:6�pXF�,r����k��Y�V��ց�����40ZZ/'�@�_c����̓�]5�Oz�ou�OI4��	W�B�rB���8�t���3�F�\[�F�tXzk�ǖ��N!o�rR��ze�PoRo�r��0Q�P7�������]����
^����9{�z���5�1^�*������2��rʆ��>�R�y}s���Y�N����I����w�f�5����/�R�A&8��5Tz�LUm+�&�%��j���o
o���ދV3�s�a��k(���8����Þ���*�T5N#*�ϹUb��oæұ��Qe��t�Y�wV����LW��-�w�&����QLTOh	�K��@���o���D�I&���W)vǅ�r����3CWt�;R,&M
�=G#�L���m���;���֎�.����8c�Ԭ+o�\g*(Ò6!�/,D����mM�2�Vsˏ��{����[��@vzñU�ڦ��4`C��L:%�$��؜7�ỻ�_���ݞ^���������Lm���pUzmwS�XD}��z�I���(��O�K�Ֆ��IH��zp�5,&��C��3��T�ق�pح�{B�[�{��fV!J oM�a�f���x{#��~B#���0�{u׳����)<�ꭁ`Ë��&n�}�y���`�,�O�9^����L�{l3<=�|r��bn���B�b�f'���T��f4o��?��P7E�ѝ�Rl���RV������k��.��j�o^ϋ%��R���}��O�/'y$w�p|z��ܯ�CN��}XV����{G{�'�5�6s�{��h�ɬ�C�g̠�����7n�F�$���A�`���w�	YY�òz��+9�z�b�rW[yN,cK�d��~s,N>�/�k���0o%s���������z?+i-�Kܰ>(:�]J9�iA4�A�rg�Ms8tF�i8'���$�ʶ��>u��r�|�`��~���u�g?EW�T2+����]�2�iǗl�l𛾔���gç>�~ٗ
)�<0a���8ث��_�����&ڤ^����"����ny�O;�#��0EC�"--Z$�Iq��9t<)0��yv�V��w�u���� !bw9����,��.��/8cQX΢u�b����Ok.=��fkݽޅ�.����4ϋ�;6�1o,�t�h��� @��q
��N�P[^��7���Gf�^�����P,�xc��^�8�j���8j��b�̀ S��P�%�=��ve��T�Fk5�����&v7���OV[�9�v�2�IK�,���L�mg�E3<K݆�ʑM���̸�i�%G�ܭŴsu���f�wM�3/fWm����jq��e.������t&tm�*�3z�i�r�Q :�>ʼ��/Y#^��x� %��*p�(��DoL����{�q�M�Y�<@4gԊG��c%�w��3畝+I2�>�1(�?H=5�o�,�{�t��}C�Oau�F#����x<�.�"��Co��c�ї�Y݋D�<�>�[y��)��۽(J~T	������w�֠mv)I�[F{>J���Ѝ8.�y?O��Xt���}�)V������藇B0+��:�[ԓX>�K���#���Z^���gjsƌ?u$��6-�\pUMV��>���<��74/Tw�/�hú��w�CV���Z�86<�F��,�+���Y]�iC"�n��,��gr�Pq�����ϋ�D��}��]���,�>,��[�� �a�Gbv=��dSz�΍e��ӏCor����Ϟ�zt;��\�y�"�Vx���.��p�5m���Υ���\内��T�5,��	��a���+NG\�|����&���%��`yD���K�b.����������㬶�$�qU��/Z �J᩵�*b�N��L�+���Uez�F-����;�Y��3j���9�Yi�
X޻Z'P��n�b�5;��2��p��`x�N0ev��u��&���լ��%6��׻�L�5�`�܆Y�{R�����+#�|j6������c�*�12M�t�eQ�y]�k���IH��]������L�������a�c�UEیt��[�*b���u�a�G�fm{gI�:�ذg���
�/9�,��cTw�>�Q�g����;AМ\*^��R��;&�y��w���t`N�W ���3�^�UY/Ty�Й�f+h��޿Z������{��{JRo3��� �y)&x��XzC�*ش�agz�;�l��N��;�#����-�֚b�n���OU(��ЙH��FK���7P�,�.�0����>n��F�R�>.T�
��{��"�zE{R~Ȏ&��pߎN��ޗ.�_.s��^�٤0fb�xM�h�0��@� ��g�B5�&���~�̵�{��j^����v��Z�QF��;��h���_�� �}0���
K��K��!�g���V�PH�՟UV�X�1�*�����&;c�$f'�Ԙ�Pԛ2<[�G_�<��x�9�f�U�^ɥ (x[V��oW����a��юVfý4�z8�Z���͂Rٸ�_V�b(c ^�X��$�e�̕%.܄�H�osԻ;6ᰘ��S��ًl_;�4˔�3�H��ܚ��f��z��]i��s��wk��@Ϳ
1�	�E�h����`�}���^[t�zk�'O��MN����bXc=QqV~f҆F�I���B�3}���C�{��z����E��B{&��7�u�dK�V}�I�^�`�����*k���gD�߽&�J�7`�?q�x��׺[<γ�����b$ӭ��Ё���ĶZ�fl�C�$�l����3����fy
�od�Ǹj�ы��*�sHA� �蠣|�m�c�楱��gc�-4]��}�=(5��	�.
τQV�+Aal�)�8�mz)
�/�6�[(����v�v�e�x�)h3)A&[�`V�c4�x���ΊŎ�]Ɖ��������{2��J�q+M
���6�}�&J H� ��3��V���-�߱`���zL��9Rc��_���ϥLL\��kq�ME�d���
ȝ[P�&�[R�(S>���m�0:F���p�ky�.���ce(��򬳕"�dШB�=�	_��BB�WT�ٽ��3�o�#qT�[�մ23��먮.=f�
��+�	E+����3���� Ȱ[��3��;D���Q�Y�+v�-f��]'Xz�gv�q�,e;��2Ab���`�,b��4�i@�d�a���or�"���6�N��;[��/U�k�f�<�	���?����Xf��a[f��TQ���l.�e%%zW�%e��K��c���`>�*%�כ��K����h���F�bH��3���v�p&�-�*v�=�דó�(�k�#R��P��#��R]5R�0��
�RGC��'P���C
t�ɽϜ^��U�'��"���iT�xQ�"u��N�Y-Y�j��z�{����j�.��}�:sI[�U�jIKQ�m�4=����F{*�h����D����Z��w�X&j��t�E/��+ᓮ�1��V�=2�W���xS���ߣ�IN�M������2{�y�H���z����͸�|`ƗC�/�3�2��:,���Wi�y/	�7��9:��`^1�+�����r��ۧAy����<҂iX�\����ֱt�� y�q;3{�����aї����
���nsT7�;�VSPH^�w��ˤ��7����,�����r\�}2� �����.�1�Km|z��Vyנ�V�GC��C&�s٢���c�4�W��a�7.ud�h�7�U��&��r�{V^,�Fi^[�����oR�Íce7��ڱ�QǼjPŢ����X��������O'�mYwq^�&��T�9]i�7��j���c��W�n������E;C1w�ʔjF���p��~�a:d,��3.��C��Bў9i|�q_gi�܃%�I�Tז����=�i����ƴH5W
�X�.�Р�Eu+��H���>�^��V6G;è��s��X8_��`�V=CY��^Z���s C)��J4<_������8D��͒*��|{6��{�jϘVg���my�kk�M��N_Zy�	�V����tt.6�7�IͫH���*?OV|�7:�3�x��Wx:c��J�I^�4��K8��#C���l���^+�z�a��1Q�>���j�7v��q�;�I�,�}Cy�Sh�}	ϓ��䈃h�ClE8�;��-gU�����������$:TR�\�Uq�k7F�LZh�#��;ī\#ND�^�̵;ˠ���d/}Eo���u��z3�����2���}��;ԕ�0�ϊ4U�9z|�{z?+�H���X>���Q�+L:䦜�����>)��$�<�Ҥ�H��M�>=;��g��Q���<%i�����{do5������t;x�-a�S��5"�f�N�3*
	?o;h.Ǚ� `Wm�+;]���k�|��NI�v�ŕ�[6<	mgr��#���> ��6���6�7d.��c!Tjüf�N���v�{�%iyi/T򀨮�Ꮄ�M���B���]��u�'���v��xR��x�^���_sĆwbc/�^�j�_�s����5���~���=�*�e�:2i��[�u�'�`u�ܝ��2��.�*��r
�qZ�r�ö[U~����>�\��H���휦���k�+i���X&������Z=���cUc�n���]�.�Ӽ�\�H��	X���u�K�=�aq�ڷkG?32���ʸg�$�q�N����W���vg7�Wz/Z��u��n�����ea�288r.�c��Wb���o�*N�vN�]�u���y:�&lao��j��]]�S��������<��8MG.�|���s��=�+�<�T�+R�D�9���I`�Z������x��;�8�V}��;�_S՚��;�!*�a=S�n����@!u;��P!�C��P`�}��d������EΙ�ٺ�9v��m3Z%Q2��\�2�<�b��JH�ቓ�n�X�v.��΅�%�wv蝔���`����E��o�H3#�չܪŞ4imy�غ�0'��i�_F�paR��o�(��0��4�2���ve���i�̩Kmp��v�y4�t;��,�+F���/(sr��y��e��rr�Bhsp29��Ve3I3��@7u�����=��K��n�}R'�4L��z�L�x��}��1vQ��5������|��`�&&Yùx�(^�n��J��
�]�r�z;ؗ�{��RX�/L�����P�i�OQ.��'�xg�Tt�SÁa�t�F�Z&�݅]<n��;��l�{gReU���T�����::�r�t��^&����	���ԙ՚.��BVz�$����RVk��
���T���R�+Gp��Oz�'s��x�%,���H:�N�w���ܰ�J
i��O��k0n�2�U�������r֋��qi.��x$@��ѵ����X.�� ��C�䷕erOb���L�S_w��ջ����ixn�[�|�@'y�$���w�ު�<Ǫ��Mp�]9�6/$�|���d4Þ��]-i4�d���zwl�X���'��Z{3�$����,��AF���^g�Kaw�ʬ��\x�q,v2fΝu��W�[W��%�.QV�W�<�>�^������R*����#�@�����2A�g�]G��/��ڕ�o5ଠ.:Ux(=�w������޻����gr�z:�8� �T�]��[,1	w�"�7)�>���ka8u�8����@�egKt_)����/�vu�/�Z��Ƭ������ұ!$�+TȂ�9��e�x�L3�Wni������[t����m��l�.�������14_�5��mڤ�e��J�A�z�E�-�*x1Q7��5ʫ�陸�Ҷ�I�S�_*V����>Qڱط�\\#�oGMb���*�YL���F��
�XBa�Xu�]/�]ˠ�f]j�f�!�y�S�墭�	MN�C�����Nq��h=�
Zt��ш;��te�]-�����S{v� ��<r�H_9 ɇ���A�5Zܥ.�5}8u��Q�̼!җN�靹��0;s��O��Ef��|�t��R
a7�ϤX���>(�-���*�*��v��DjYS+pWS��\\�>��q[���tv��΂/��,pu�otKe�'��.i����thۜ�u�����yI��Wj|��F��� 初�� 9ݮ��滻��L7w@����Lj���k ��Vv]�H��Yʇh��Vֱu,�]`a��EF��Gq�Չ:\��SwXJaDf���.s_oV
�y���6��gb[����T�!�4�]Nw�����b��H��Sf�u�&���sT(tE]��V�ӣ��=�����O�X�3RwJ*�ww�u�|2�������K*\iq]���X�z㵝��󰛍U�p^&x�p�e�V��#��Y�}�+yƎT��Ϟ����÷f)Y\�����h����C�ܵa82�$��w_a�s�4W�4ξ/3�e]���tU�m�l A���6ڶ�����D�U)��7�ݙ�杇H��2f�uC��Nμ�g�g.��z�ݬ��E)�f���fh8�_5%7���~��t�eS�iJdn'r����R�݈I+yVݨD�+��XW[��1�sG�Z��fJ8�`;�Τ��ۗw9�����]A�b�<�� ����z����xa��o˳�t�t�y�s;�$]4Ժ�ջch�2	O����šЩ�Uҹ\��I������z۳�c��hf�P,[�m�^�N��p��i1Q�ә�r�v�� �%�r����^u�㲒
@�^�F�8\]��.h�X�y��6��=-�Wk̀��6�޻*��hƩ�41m�k�V����Z"�Ѳ��`.V�i��r�Z�gKR��Y+U�m����0rV��Z��>,@n�ьNTUd�½�8%��S�#�\�Х�fWL���*P��G//��l��/�]gP�.3̋�������u����f����z��<��!����c~n�8�#S��Q�c<�=�&�{w�q�ޗ�;/�����?~u~=>�OmUJʱQ�,E_Z,���j�(��(�� �Zlb�U"�&��1TVcQ�+* ��R"��"*�
���V
���l� �"�(�E�uj��U�e�c`���[V*�E�,DR�VB��b��2
��*0b��*��D+[��ŌTDF��QTQDQX�f�UTT�$TT�*Ȋ(��GM"�"�������"���#�ӌQX�Ŏ�QELj��*�b�4�,Eb�(��*1(��J�",��V�"(���*++FDcV1X ��"1ƑTTcm����DEU-)Q-R�EcZ*���
%���5��(*&2����""��*1r���{{�n����/��yݛ ��B�%͸��y4n�V��A�+����͌�NJ
��D�cr��zƈ��n����T={J>��e��i�3کLUm+�&�#�li;2]�tW��Lݬ+3���L�to�73��<L9(��� ��3������F3������nt�����RR�.�K{+�Qre{�O��%��C����QK)�������L[��9=��aaz�W�Tlt��7��o=���q��|hةN!�^U�d6L�s��^���T�NZ`�;xٟR�ڨ��g��Ņn�k�}L��B8fs��7�&���=�c��+yz%�ף���.���Ţ
�Q��.ѱN/����àLl�]/2OOk��{EEb,{�ܘ^l�����s諾6���+���kt��uOY6+\*�:HD[fm��e���֣bP��ўĩ��`�7K]���d�OW�����c�����x��]Ԛ7�7
�ᠧL^(N�Hz��}�ٿe��������李.�y,�ru��.m4���!貙A�����σ��K#�I\��pE�ߏv�F.m]{k���[Oޝ �W�z��\Y��?i�}�����~v2 t����n��}�y�+B(��Vh���,��c*�I�Im�3*D'y���zn����&�e�HL��r}�"�g_v���!*q�S����O.�y��%\(��]�Bx�mm���U4���ޙNe����o���EQmp"�EY�di)=�c��^������雡��R���#��{�2P���t�}%8ן�can��9�^��/x�}�,��}�u-ӆ�U��.������؈��6}��l^r��2��̾$���~��7P��5�B�6Ck�5^�z�]{���ue�ˬ��)�$Qrb8Up���t䉒m�p���o�<�=u*����{�X���K�9������76�Ұ�2��p��Y��+�^ UԎ9����Cg �����8���2��;6�Ű�ל�#Q�%*�E�{v�u�^z���'�t���|:�:����y�^��8'yX�X;��jV�ѓg�7���n{ɾy�������u�v �g��c�1t��@��z��u���-,���W�>{��
��Z�1�p��D���P�K�`s�_�i���,�YZ@�j2�[� �{�� -Y�.�R��`J��n��}�e: fz�� *�Njͧ[b\�¶-�3>�jH�:��]�+���evv;&�k�F�:k~��/�t��H�F$y��B;��] �cM"e��N��k��	�I��B��Kp�w��t&�sݪ ^��J������:@����l��F.�"��Co��`�^\�4�<���.���>���><��P%}�P_v�t_K^4�=h����c�l�ܙN����r��)�����W������J$*P�^逗��Yag�ޤ����W�Y��sdt��X`���|mAB�sJ���D���z�j��2Z�`��wV�a=�k9��]y��^�y%'.5@x{���Z3�0�]/����W��u�6]n�8;g{y�7�GˆϜ��s�{�zK�(F�G ��|�ƶ�u>Lb�k�ڂf
�18;[�GO�W}�2��,X�{�L�k�a��Ǵ�>����S�V%���Ep�1�^�'r×�#x�u�p	�ǔM�K��N�X&�=.
�ꖙ%�U���~� ���?��Y��� 9�m
U�����*6���͉t�(r���9��Aڗ�����]��5X�p�g˷�{�y|�a�>�G�D���ex�1�88r.�`ȷ�
��ɱP��J魭;}Њ���2R����Ά2�j�r�7�yeh������K���ǒ�A7P�X�u+V�2srR��_m�octH9����:����l+�eE��ɒ%�8�s2uL؀�狩r������Y'#L�ܫ�D�����l�&��~��P��A�we���a�Xg�f^���C��D�e/#��u�S'l�y��]��T��%V�/쌒GZ$I�|v���4M��������f2FC�w�5�/u�Νi��*W��,3*'pQ2_ؘ���|7���Gz��#���E�2n��4�0ϒ�[����<�`z�ß	d�3��b���s��8x.��{
t�kOaT/O 6j�P�|N�`�T���ʑ^�G��"9I�&Ll�=~b��g@���Mly�4�	��\%���h޵	W�PO���r9td�Zwּ`�97�'tٶ�f�턺c������N�5Rͅf�y$s���3��=]�Z��E�/M�:R7��Y0IAZ,s�T��:�
���c,UKC�)��:�3Ub�#��<�����omG��SS *}/T��H��Q�V�ϨJ[��V��;�����x�����Tms��9�fS)�t�3��t����n�wY	 ����0{�B���__�:E%�;�.���=C�	�)�U��í:��ƴsO(�W,T�'v��yI#�a����,:�п2��]�u84H��m�Wײ����o.Ki�+�b�X:	`�j�2r8`��)�ӿ�j�?o�ë�7f	�C�l�gY�{��Jĝ���?W�h���ث9'�T&�N����>�K|˭��m4�W���6��ޏ=�KV�}��<��V#�?'+a��/ԝ��d4Þ��]�`�O�_T�Zx^zs�ee��j2�{�*+y[���2�~H@���`�������2�������]ӓ�/0�0�V��&8Rr|p���dj��4�[>�
g�+^�B�]>��&���Q��,�5A�_�Ϣ缰z
Һ�RQ��:���˭T�*D��߬�����砅^/)<��c��M���8�{yAY5Q�73��ZL9^���>H0�8Y�3�AX�ݭkϵtX�9�Ҧߨⴍ�Ń���Z0�^�S��.n���jOR0��B���`<���i��m����!ډ�u�J
��(�o�Å�簽_�f0�|��h;�Y�Wug+�_��rۊ͓�*��F7v7�tM6_O?�����a��XV��p�eg:��^���^��8l��N��1KfU_��eN��<.y��̪k`�K��0��0I�ҦL������.�0y��9�\u4)�s�4N#�����mZ8�������vs�]���S�{�]w(�P�m=Ϡ��Ռ�3y��RyA8�
�����m̷�e=�f�O:����]2��òV����'GdU�c�1�������!Ժu�ҁ�w>s��c(7Ctz�x���	ʯM�a�LXl���Nd:�U^?��nt�ʷv���.�#b��l6E��kI�C
"�[F{T��0W��W�� .0Jo�{��:�#���6��E*}Y�m��T�������ǠX=k~�P�{3!�P�^8����?��o����9*�*=O�`�:f0�$�VL��g��^ tnZ��<��n��=P�
2czu����,^��u�/�ttf�=�A��v%s�f�����ut��W9p^9�K�+��/�}g(N϶��U��E��t9T҂I�ɱ����7{�>��y���\��-�E�rӗ�M���a����-���S�����Фԅxx^o~�4�1����G_MQ�ܑ�'�.S��	�5�B��X�j{Q| <Zuǯ/2{�UA����s*wP�RJ����P�`d�ij�rKÔp�������W��׮�Ou���7��K����X;�n�t����X�3�Y�<Р����x�N;&mIVl�o���ON�アՖ]ݰ�#����Wֵ���)t��3r;[�������V<$X�+l�f�ŢvU�YŮ�Քʝ�Ͼ��a���.�u�3u$�����¢IDf-9���:]ة��V��r9��r�f�䐖��W^ҳ����M����efx�>�����3�Roo�k�y�:P{����X#ީ��fo}����^xZ��Sw����jQ�FSң�ݯ>����'�����=k���Dr2L�yTO�7ް���`h��¨;���}��XNM���4-�.|=7C��K!�/�GC��X���e-��^,�Q��{~�'�m�F�|tڢ%i~%�&P]��A	���<2�כF�!GDSɞ�5�܍��-�q���Z�7���/�Lo+�2��f辖�h�"�<�'oy�ϓ�.����z�}:�b�f���[?�-��3u<0]w��� Qߢ�t�	bz,�ZG*窳�����$�D�NZK�p�=J�1^d��S������F�����f����vmH��B�)��Ф^IM:
�@`u8zƛZX��s�u�*�Zn�iyrNu)7�^�i�*�]`��ҽR^�C�"��x���3�MxP����a�w���ĺf��C���]vnU�\<]���o�i��e����J�:Π������Gc�����Ɨ ���X��9w�����Le���r�[���/�x���c��s�� �k}�DժI Vs�vۮ�e���f���+Γ��r��Fr�}U
ga�8 ��<&�~>O=z��.�mB�]U2�����צ|����:�PӓgL�{+��E�ܠ����h�KL�ƪ��Kp�ɵ~��ﻈ3�K�pJ��}�� �*�2cv��5WN֎~fe1�_�p7[�$�6^<�{�X�䔋��6���O"ϝ�	=�����cM�����������^�5mg�D�e��Ώ�r����t�;ǭ�@�p�bb�w�>�Q�=�Bھ�N��q+�e��n_��o�bR�H�]$�����&��<pD%��O���I�a�о�L7�Z_^ث�w��%�L�@�ڋ*ش�UU��9y���C�N���A�ư
���cX7�,L�O"����#&'�+�U�}��M��edg��Z�*�MD�={=+R�0��w�b_�S؂��Ju�o�D�9������^ܽ�d;gr���8��N�ި�0:�4;�#D���~�X���'x�<l����>u瘏����/K12+��5�u�d�0:x�^a�.��)A�P1����f�e ����w�=�vMj�ԫ����Qe�9ѻ��tâ�v�q��k�۽�N�7]��v�yz�5���s�}h�i�Is^P�m�"_�M`1�����^�AV�SÁa�u���Z)P��'>.�'ks��fj\ 1�`\�!��W���KGg�Sc/�ha�����;c�3yW����2k��J�bF|̡��XL�UOG�+�y�L	��/\U��`�����(%g����^�R.�S�����&}2�W���f҆Tj����u�����us�%��-�۽�{���zW�TW�h�\��Y�=����sϤR�r�tӷ�~ x������{&����,yDο��h����$�~���)1{��\�\�LU�V���[�0�����+|%�C�#�t����ه:Q;����ב�}���;'�-!�Ϣ�(Gٙ^��K�\*ƨ�|ʸu��B���V[��vɅ��o9ŏ�Tk�Ɏ�|fE�y`��u�0���ƪ�/�T�*�i_y`.�ɜ���䔮M���VeW)"���PU�ۣnngkGR��ADȑ�p�O#��w�D��Lt~�ߺ�VN.��i˖�$_ѭe��T:��pR�Ask\i��Z)����*3!��DW�l(+���<8�eH2�g���:�3绽خŬ��J+�eN�ʰn�s�,G����8�Q��K�ܭ�����ʤ�6�2D��
>C�����]��+4�߭X���O�1|��.W�N�n�$��V2QD3s�9��{��ة��r��%�k�,PV{P���Å��v�����1Ep�F�6��۽�L9��G0��������y�M�ddw`�:�����ǌ^s���J$����+�ٻ)���8�*���T^Xib�`���/ភL��-���yF�iY��̹�Z�+H����:�LW0;�^���6���_ӟ�?��*/e*gD��%�*����tf:�i�f�n��I�H�s����z�� >�T���j7(aDT�h�`J��
����_6o*���\ؠ�1nӵ����kv{�+C6
�O�7
�ᠧL^(d�.��������ׄ�g8��J�t��ӺT8�n	�p�ZUᰌ�YA�~��
s޺S�o���9�cn_9��V�V�稄$5�E���홤�Um�yN02z��ޙ�;~�UT��3��r��|�Q����wD�v�ֈ0���BUr���������ru�>�~�H@��$�	'� IG�$ IB���$ I?xB��@�$��	!I��$�	'�@�$��	!I��$ I7H@�XB����$���$��B��H@���	!I�$ I?XB��B���PVI��c}C�@:�w��X���y�d���Wǀ��  �T� =h �@��C@R�((i��)Ѫ�-e��mkm����f�)Z�ٲ���5eSF�ֳi
U�v3m[[<���[5lmj��m��4��lSM`ҭm-��e���V��+-V���қY�Y��}�z��J� / l2�#Mvt`Q�Ҧ�3l-X��,b��Ҷ�Rt�[��  o o]�P��%AmC �����;�p�;`�s���&�c6ڴ��� �CI�@�bւɍ4V���VeZwp+]�6�K�����3vʞ���ɢ�uK��^ =@y��uEY�����  �X   �� :  ��   Ps   :��C�I�=:�=�:U٥�[����b� �z]gi�e)�t�]�1��v���y�Oct����u�#��j]�:�ۮB�ER��Z�U�lم� �k�i�v��Ү���]���(�JT��)�Gwn��7oLJ�Jt�7vzIz�oAu�洍f�֭Y �zt��C�#��Ҟ����V�q[[t�n�oN���\m��7m�;��	���6F��ͤZ�x v�٪j�2���m5Y��6�"��b����5haR��jU���`�ў �����-0/s�P��-�`$��U��C#[m,(1�5XƵ)���=֨���L�֒�0i��[
��:2������6l-m鸞 
 L*R���� ���� O�*��@�a hd�1������ @     E=����!#F���2 �a4�(��L@�5OSڌ��h�&OM��I �R��=bz� i�ɼ�˄�>t��ǟ;Z�2�o�0�6�ӕ1��0�)��  4a�.2w���G� �D@� �� ��V'����"B���x"A����|с  CFR��	�&  �q쾹��f�uq��U���ZY�5K�q0w�:��@�hU�����_��V�~�~�@����7 l��cn�51Hq]%.NaL$��W�7���pj3y=��iٌ��ַ�iؚN=���n������
H+�/r_�Qgl)�/�NS�!�	��KY*�,�L�!%\�vn<	M݌3�l�XE�7p�s�&�P7n���ъ�ˤUr��NMp^xʖ=����m�n�绝�x�6��#�rHF9�Ӥ�vE���f�A�R�I��&79�fήY;z�am�qp����聊s�+�D�eZp�ܱf�m�9�^w%��єgW�r�۬�a�H�C�l��>+�bc���goX�x�8���>��-[�/˙: ��9ƣA��,�=��遄�U��Y؁�q�3���sq�,�����e�9ot����j�ͦmW��AF^�w�Y0���n��	��`���z*u+;c��=�O_.�x��.�K1f��@ï6�օ�j³y	�
p��W�Ls�#;s�P3����V��ؖj�Q�J�_��/4k�Ɗ8Wq�!���W8�tKisf�4�\ܤ��,ws_n3t%0�w,4)��%Dx鐭m���XtuΆ���|�م��*���֎YXy��.D"�C�ۯ��!��<N���\(q{c�w��OU������%ờ�A
�NŮ}�[�1J��]��#I��`�_Q��.�}ٯD"�]]ԑq<���}QV��򻣁�^s¹>�3�=on[�w7|�\mil��]�{]��=��E�wk���@|�`q;�V�h�U���z�R5���ɵ�*��r`����W�n��`Q�-kh���$x �@�ج_Sn���\�e��7c�4,t�~�DV�*���5^֍oE�͗_-�S77��{(�6��C-S��v�҉�P�U;x;�F�.��Q>%G�b��^��\1
.>|����)ؚ]���"^'mXx�B��L�J����q�(o+rF�3�+��r�,��
n¸�ے�M����;�l�� K��7�$v���r ~x�|� ����gMɈ�=�w8�Yl�(&β�*J�Q�	��[�\��J-��8�^�Ѻj��'�W��{��{����ZYM��س�jʝU�0�!�]@;7������	2`�w��#�����4c�'��q(H
�Ĉuf�D��4.��1�ӏ�� c�79P���aһW�D�X}��*9��L�2�9\[�q�����Q��tkj�n���z� nզ�����������9M�Nڇv�4Q��3��ֱ��Ɠ:�چU�G�4E��� !��3z�>���	.�(����r�3���b�^�pW�j��۪��^B���7�k������8����أ�g�;w�n�+C�š�L�6�>��T���0�v�����k���	ԭ��(1�8��4���m�r�ܓp����9,?=��(��&��b�ř�*�Ɠ`V#�����)�f���9we�je̺�H!E��8��ˁ�X�
�<�Fr	���g`��h��F��N�.K�.�s;�C�6�eҝ#	F�ufG��âj`s�]OW�s�i�as��{^��4��n��j��N�8#pkL�>�7���\��`-�1�����f��i1�גY�[����*;�@6wu5G�ĊF�a#Q��ɫs����+4o7t"F,W[�,a��ޤi���Xiad(�M\
#l����ˊ3��o)��hlw(����eQ���x���F��S;Zw��c�EΚ��Kӄ+�X˺�Uۏ�ұ�4Wc�a�8&�AF#s�d��"{_c���;���bM8V<�	���[��[�!��N��t�5vP�xq v�y�/_}fӂӯ���aqq�|f.��k\�ѡʈ�檸�(��L�Z��{�X�U�7_}��a���n均p�S�,�s����]Y�v�7�Ca��z���{y�����VINe�z����������'xr\�)("�k[Y��njCH�52�P��Ɍ��K|��О�	u`ӓ8����oAL��8ѭez�a��Bv�͘;����
We�n%I�f���b�"�Ē7�;1�x�հ'f��h;�f�w���Fu]:�\�
%��s
[�;ܭ`p�[����:P�t��vQ
Wm�Uu�ӒR�b8Hh�)��a`iV���.Cabޱ׋�<��}��K�,�n�X��q�\u�5=-@V��;�8j&���{�c��L�ѪVs��=e�NT��t&��7�v�L���ƍ�4�t��P�ovLJ�O�d�C��6��D�_,���Ǌ�jӔ�x����q�U��,SR:y���##C+=�h':����K x��0ZVٲf��z������Pu����*�ƛ<��ڠ�G!�����i!���&�(a����At�u�Akӌ�$,quɅ2��� ���uK؊X~��&�K�i��z��������M9ˋ�|��ٹ$7��К����T��N`�4Ђ׃�뼎A5M@o^�WE��P-s�]Vm�ʈ`܄k{�����p�y0n;��$��.5��G�bcf�E]&32�Ӄ[��y��${��j�;���!�L�c���eH�K�/"�;UˮL�J�(�:���('y�Bfiwz���|f��h�K�ka��iI'4�+n�2<S���Y��E�����X�����ZV�Zx	�r
*�S:p�;��2d-���t��zߺҞ��#m�vBh[�f^KyR⻩��7)ҧ4��q$�(sp�Ѩ.I���!qS�:�e�{4��;Ih3�g/n���@�{��c̬t�ݠC�����:����]��Zx7�`uv��8�|�n9h�ջ�9T�������9GL����Ty���Ђ�jӯ����5Ux���wϭT�����5�J��8OB5��"7ñ�b�mz^�7���,�Q�N��໵iBnV��nP;q�嬈�p�J�;���čU5HE�C�����+m}K�k�/�V�̙	w�uIg����_P�> ��j'�ȩэ��G���ʧ1|'o	N(S����SR.h�f�YNv��J�`7FN��d��-�4m%��ђ�Ѯt0��(K�PR{f�x��(�;��_.�ΧnE;[:���n^GL�{���B��L!��,A��!!�\��g�߭�_B��e�f�2s:�v���^&6g
�|�֭�q�S�$�@,TZ�D M���NYIGtdt��x�1�B�Y�Df�ѧ6� �^˻�)�������AY�v=;�B�m,N/~�S��E�ڹ�jU���9n�q���C��q�Kq�����vL�7��	���lk.���22Q�3Tp֔7��0jSa��/Zd3"�Zv�Ǔ�;��P�Ƅe+�L�.�E�V��z��m�R����>��9�;KŜ���Ve'n�^]'A�y�����Ĉ��A���W�vp������8n�T�m��0L���sX<�X�:g-��T;�����Y�;���f�������5�kͯ�)�l�6�@�}tiS^��Tݸ���X���3\z�kv��]Rq(X8��W���M���YX�c��]k"�
:�X^��$�k4j-|�`�q2n���]Ҩ�5�t�X��tj|ᱥ�1�n'Iw������,K`h=�ۃw%	�����	��S�Yj
6S4L��7�Z�![��{��z�59@<%ǹ����X�%�4��:7�X�O�kL�VU��o݋4r8Z��P�J��-D��3���v<��mFm�t,5�qeBD���k�ӻ�^��:D�w,�)�F��l��sp�l&
#�p�����<��S8�,@���/��fM2�~���J_���~˲�wNI5�{������Ɏ��H���`}�:�*f���i��c��RG�&LWR�آ��[(}¹�#sn�����D���-V��(;�Ɩb� ���IO�!L@p܇!Z��t{'���WM��z	�� �f{� h�O{��;w����2\l8N�a���
l�b�N3E�.tt{V+����N�.�wBq������ƶ�\�oc�]�@s�����Y؜��1h��Yك���A�"��Ү��s.,�:U���7z��V����7�g"�NW*��<�ek�������z����#�Q�)�Kf]
�7(�&����l�y"���Z�!�Ώ��������nNY\���K�3��א_��1޲P_c���8��K0K|^�o�ծ���ԓ��ܕ*�T��	��r�[}P�+��J48�J��Z�t�����փw5V�1��d�V��Cz�lg9��՚��Y�|�Kg��vFxU�h�&![��x�#6Ws��ne�T3������@/RFlX+��7�Cw_|��(����a~Bm} �í�.�|'_U��'\�kx�Y@WV����#�%�
�J��k��-F���X(�+ZL�)c���Δ)�7���<Z��:�l����HIf��Yf�7���.��S��m�ڀ�}�])�3R���ºN�B�8��e�3C�����B%8��J���s�������x��Q�y�ѽ^�����Y�[6���u=�r�F�RN������r��|���mj��-��H�/4�7��u��M�u�z��,��VZ���Q�Y�K5g(��%�|��Ζ�jc��cn:nF�<eL<YsK�g:��9�m����y([�p��I�.�-#�Qn�[�y�Y�.�&&
)���!�ywK�;�K&�.�� {S��2�j�����q�f �!#|$qvK�G8���8)*G�u�ޒ�!���Qһ�w#�h!�L{���ϴw@I��I<ر׀%ͨwJ�&_��(���P�N�q�Ö�ʕ��wB�[���&����@�=�;юgc^z�{w�z�q���R���X�v1��m�M�;QE��B�&�%F����J
�L�'.���u	���D���[�a�S��E\Jc�O�ƫ�q���4�ӉCR�#����v��C��$���ң��d&�c�ɱ�n�]��&�)^Qw�k������}�ט�+Jv�U�R���A�W'v��wu��/(�e-�,u�>�ٶlY����}g�ނ�ۭԊ�K�!=�Wܩ�0_wFI��G%9\6At&�@�W����K�6�{���T�;���N�A0�8�qؕߋgAP�{mZ]��X��p���ݺ�%�g��6���zB�r�6�D�:��6��_!M�g9��8��D�b��p�� ��i�}��;�N���,����H��Z�b�q	���L�wY�E�{tI�j]l=�60��z��-U"�iL�(1�����Ƭ����kS-[joq��՗��{P_[��٫�q"����O��"RבQ��)ڮ=��K���!RGEF�Nb\B�g�zr^b|��V쏣�� ��E�w��2�Kr�uA�Y����S�u�S`
�1�ν��{~�&I�r�v�h�)Z�-ܕr�&�q�Uq�'LՎ��6�]N-��ѐH�]�/r^��r�`�l��I��/5k6U��.m$7K���t��&��^���j,��d���Ӫ������kۖ�����G��SA���SG00�-.Uw��ZjI�L~�����d�|w=��8<8t�ܞ�e<��Q\�G�U�KW����Y�HdmlE=WuzC�"0�ws��u��!��WX4��9ή]� �LD��;�������G���^����.����%���9�K�8Y�����p���N4�)��T�-����M��F��s�y���ȋ���p��NJ��{(D�qG ����=ۜ8u�V��]��":9ʹ�V�Yf�8��ȫ���O�؄�rV�6S��������k��'�Ӌjթ���Ř똑��[�_ql@���2.Vӽ���N��o+�WQf?��dp���U�eh������4;�P�S������0��**DЫ$�:�<���sa�FsVh��H4y�ۆ�������L���htA���g��Mɖ�˒�%�W��W,��WZ��
�5�����~����g�kq�}��W�^�R�<���T���f��f�6���G�np�p�=�iZ���Uz��#J*}�N��]����b����{xdƄ0֍��d`�'m����6L���l�_f(^��W����h�.o;�r�r�=�ˁ��'��E麼	D�@���s��z/�B��]v��U�p�M�᧵�[��I�e!�=�y�g���r0e:�V�!�����/z�8X��ʕ�uz��eq�&�<Us�y0M���G�1���=��Y�W*������,��qNU�;1)���C�RZ�z�ˣ���{MU�+s��)����`溵٥R����`wu�؎.��:�
��|�fT�Q\�E�X��J�>�5-t2�eB-jwv�$���n��;�I&!k��mi\KNL��&���¬r��� ��^�YO�XX���q�:��ֻI\˫N�l�1�Uu����C��E<�s���Ӏ���W4�]co�Et��+�pD��^v�J�h�9 �OT2�\pv��j�F�����<�����z����C�qLX�-x�&j*�e����e��S�6��uԥ���N��n�z��'�z%L ����՞�LV��F���L���εY.���]Ix�ؼ8X����2��0��-I+2�]ݽ��R�B���c��!}�P�8��W�^����9HB=B��镪Ä×Y��N�6�!5��qN��Y0��Ư|E'rA�v��Ԗ&�ɲڮC���M-4:��G�ѕ{�a�ȯPL����5��^�`|=mѝ�EU��o������X���9PXZg����7B�i�DU�*؅k�^3؜z p��]nIͨ����j�>�S9���|���q*�!+�,0S��R\ 3�[�5���M��9j��7���rZ�"� �^A%L��7�U�ץ�4S״2��6*��Է8��{�j~�:r�L�p�����o9�T�.K��r�V�YR�橁�M�088�K{w*�J4�S�
��9gt�A��XQ��y=&'f�n�T.Lr�VyQ�$�p}�4�wd#��p�';�(�@���0ٛ}�7��}��X�rwي��mMe���/��=�u`�����j�S[)�*&i�J�d�l��8o3q���;1��t��qɛ�'7M�b�m�N���63"�sk��jI�;Ơ{W���x.s�lH�EVδ���G��v���R�J�4���˾r"��c����;�}ރ3,��ʝh�Y�/oZ������<U�}"jE
��BI��#�`�#=��$�D�r �G$q�rRK�% e�:8�q�-H�٫IC$̭������/1�Ny7q<�1�p.�M�LK�/6Ey�K���G`�|�.�S��WTz�HI���N%63�wI��E�֋�z�2��8�F0�Lwr4��|ui��ObSE��{{�a�yl�ho��j��I(^�WñД�.ΫȪT��nفI��Gf�r�C�J�\��[�2:Kbլ9ҜV8:�1Ԭh��Ngo��f�
묚]�I�:�5l4�SF��鞠ݡ󮣕a�f:�rFB�g"Q�ge�Wke~��r=��󴸦���]F�0!Z{`;}2�hè�4oۚ�Ff�t����B���k�A�q��{;����U�H�z�}/���:BU��hdK�bX߹q��D��@�INǹ�F9��*�{_h�:�yd٧`����O���%����>L��M�V�GI�R|&�@Xrr��x�,� �����E\�a�ų:��w~�ve��"ٺ�W�]{��WfS.+����_���3#9�o|���	mL�]Ն�"��T������]�ڼ����)��:lL�wCY��l�K�I�ݦP�"	
B�y�-�B��eyy��M�~@��������dq;�v�ٗX��s��ũ��t�ݰ�	���?E��7/��8���l�*�������X̃�/;%�D�� ��H��\����E<�ӎU���X�_Kj�ql�ԡ���6��՗S\���m=�G������W %R�Ca*u�}.�N��5?%G�Nt;��@e����A��ْ���/�pQ�̄}:�v���D���O� F���1��jq��M�a�C���a^\3ްqjU�^织��������6����>�%A"q_���{(�҅?���s�آ�/�d�Z���\��A^��9��|��͐E�5���f�Ti�\x�Ӊy��3IH˼�J(9$�-Ys_�Oݺ��21S�0�׽��R&=�[G�b�!�r=��ryn�	�-u�lF�m��
�'^:F�4�gR�s�)p7j�%}����N��*��6m6��V�K��e�&Z��J5	�5�:tl1wc���ݴa�x�"�{��3c�V�ۣ�2�=�&.�\
�Ԯ�̂w]���E��ڔb�6�Ho7kA�stn��ޮ��8.�0��J�j={�	��#a��Sܫ�Y]��N0�����Γ�i�wR-�ޭ��kI1
��+��F�,ˌJ���+��~c���F�H�O*�ݲg'�2�� ~B?n9����v�Unύ�2fۭ0�^ճr�=�O�G��J���˷�Q�S����+��l��r}���JAp��8���9J���Iq����1MO�>	��d�f��l2�a��xI�ĕ/�"��2�&x�2��5{�y�I}.:��/��Rd��H�+RVJ���t��ȹ�.e]n���n403<�>�炑�����酋D���Ky
�k�(���d���Ѝ)1ڡ�����v��h�{�0��:�k��F��.TޖD�}&�]�8���!ٶ^֫�R|(�E!�(���W`gPўi�K�r+�,��_���UO}đt���6r��$8g�1�0s�C��mL�+E�q��cT����_˴B��0����Y=|�tb,�[�3�ff�(Z��+�����"�$����cnlЬ^�x�t�x��gl���m\�wu�"����R�&:�H���&�KT�mfM��.Rև� �͑}V�vZ�u��b��ٚ�#�� �N�`<����_hu��k)8��iU���e��`!�m�Du'��of����o�kw`+�ZQ���Jy�f��l�>�[[W
hX1�ս�a���.˓e�@qL��vnQ��q��eJf��j���-t��~YUx�����9��g����^C�;"Ù�sG��rPo�V�Z�4!�8�����I;a�֞����7gz�,�(x�:I�ՁD�����9T7c}M�Ĝ�7ۊ�O�mMGkc�;�_x���~�� ��!(qf��C�L���5;������xҥ�q�G<���sK�<"��M4�yס�g�{��=�,��]*��`���:v����(	�YDe�j_#C^�zd
.P�hf��<�n��{ՁJ�Y����f�t'*)S!ŕq��-��پF�H�u_!qX�_l�gls�� N}�+�rۺ�8um�IWI�]�ںa����\Z6�s�%C��1u��xq�آ[�%��$3�'��f%�.[���N����~�k4}��Ӳ��CoVܗ#q�+k�/�
��խ��e�8C��튙�3I̫yƻ܊�U[}�K¸]����\�V����NM�һ2m!3�G>��ڔ�1�T���_D�u�!I\����m���E�B|;~�V_�?o
��o�rF�#0̓���6A��tf��4M�BR�ۼ�V�7Kݥ>Y��_dս����8� �0�]�����\�:5�E��Kq[Y�Nq��7��բ�=�j����2YE�#�]/ڃH����V��}k�4�;��}����.�����S4䉹�v'-ۖ:�����$L��2۹����<��w%w�d��݇���>����zP1�_�)�O,<z,��:rO�c�8vń�t���g#�7�������*fU֜���T:�U�-��`QYe�}nlV�NO�(!�9��ꃨ��un��[����|��ߖ���fx������P;>��9��e֙�pf���R��h����ӞS��J�`��Z�N�⫓8�g{w#&�gB*�S�%f
Sv+qGl�EE��	�V6u��ńͧ�ѷL�7:r�"=��E��;V��7�9�=�Z�&MqW�/W���-�x`f��w���o3��R�v#Z�'�P�����Mvh������Ӵ���um����[�{���_�R��8��=�z���d�V��dcۊ�YckI;�w�9�3����)_h꿭�3%
s�۶{���$��{��DwPӑۡ{�2��9��a!��[6��R�xAϟb<ﳀ7[ҏTaB��X4Ա�[�?�v9y ���J̖��s~<����xd��I�Ww�f?BF�I�6QF��[wY�N�/6�"�M� ^�jB?|���D�ao��|P���^YdR�C7�fff�H��>ь��f��D�Զ��i5A�`l��ܐol�C{w�����	07J�Ua@5#�m%�9��]gn�l4@�&!�n92�J���nj�f�u�60V(=G�װY��VJ�qI��X�!�}Âw,p�'�d��-��Y<�9�Q7f�R�չ�tf�)	��thF�e{}`󛛫^k�64{�`��pZOL9�ۀ�/��������^i=;f�]�>����k(WQ���:����;%b��ӼN1�DÛJ�=l�a3N�^�wt���� ̜�չf]��-V)m�E{��QT1�Ն������\�84x�]�;��Թ=*e�fsu^|�
����fub"j�d;��.
9��s���sD��
�W��J�m�����1KA����pWЎ�U�`���Ac� ���"%!�jL�Y��N�<A}45˭��!�Ն�{տ�=OP⭂c>�8<2 �v��.�g�x����;|�S��6�8�Vgp짣"�(�����xM�u��9�
J���Ξ�:r=��]*�K93#���Z�L���-��-�̽#0�||�ѽj`�]w�[��R:;1M�M�Jw,;;����ڶ��5�5�+�R	Iy]�wnm^�B<�@oכ��1,x��˝�+~�qOp��U��m�I>�y��rD�t��G$�Pcup,��Zxd��u&�y�u���������i����� �E@i�R^��V'W�UΗ+�����@�1�k& �L�#������3����X�L�OW�u;��H&�Tu�{�ۢPZ�,�r�-*�3.[��x�M�v�8ɗY���Gԝ���9�5����RA��!�ڰ��G��g<��U9�ꏺ�X2����Hf��S]��P]�{/;�mY��������l�*��;���7l�93@���te!X4{Fz�-��Gϑ���'�ͷ�������3S����� 2�]v��#-jʢHx���7Wr8Ƶ����@���і���}�0;V�s�H�������9,\��u@��ؼ������vd��ۂu��`5�M�ʶ0@�=Ţj�W$��c3�x��b�;�������x��[�:�t��D�w)�38lClp���J ��U,�G9�p*�&d���b��ۼ湋��U���iN���s�`S]]�Wn���T��)��D�(��Znmohg�Y�zXA֯u�[]j4�m���V��Ý�
����]PЬ���!�#*���h4faf�vs�����f��Z�T�#�P�nƝ��v/A<.K�-m^,qJxܫ{}�-5d)��a��A)b�՜Ю`���4��@�'/d��,0]���� $�@T��h����,cWߟ(���ȱ&�&7��\Q��oH��+�Y���
�������I���8N4�u�ݢ5'{Wh]C�p��:�J��7��k�l�\���6�\�^�&��5HWe�=�=n�,�3��?��eE���=l�̣�����GW�^��Yr�L��b�:���.���5^�C���'N�� ʯ���n��y���C7�v�{����8[r��۹N��7��v�Xt��d���=QqЦ�.�j����\oӲ��هvv�rZ2D�a#8����mlX�/��[(��&�ި
ԇ����H��>�$'@�C[8Ĵ8�tu3IÆ'�q�Tj�c�0��H��D���19��ܢ�@�
�&.��p�WFY�:s�|�"SC �7�]q�w��v��oa1�t���>k����w�t1JŒ��IXV,��h�a+%gL0Fe��9�\i���c�`��T��L@R�m#[�%fE�B�(b)m(���")�
�2��`)(�j*�ʡc"���墕���@SHU@]R��T�j"�e���Q`�h����V
ږ�U+F����mJ+f5��UjTUJնT�5�Fб�Vc*օjVԥb���D�K"�墨�Z�X��qUUY[mJ���Qj$n��h���DΧ�	����5�Ypʍ��Q&����d�-��d���������z���t@�4FFUe}x1��c��uqe�ǹ� <�q���S�7�k�8�<Vmٌ�S�c{f���i@<����;R5
���6p[��:2�÷��ա�kK�i�@� 3�b��Nƶ��LӶ���cOB�s!���KN��/�[n;!�8���J2��d)蚦/X-]-[O9�cN,&0���wI�a�͚��kj+k��y�����۩�δ��̾���5��P�s��/�@?M|���b���۾�e�6B�kT�9݋z�(����t���x}(��-p�D6�)���;m6�+��.�A��Cd�M^T�`l�s�u�����0,����%��
Z..�ܝ�F�OCp�:�6�΂�j*	?!�B+�\q-N�d�7n�K\�B�r�.����t^>H��=�xJ���w���=<�*2v
ͳ�d�q�/���ۧY�"��p!��9�iVh�|�gu�o{9'�o��t-,V"r�Ե�
tgq�X�sϔ��'���w`m����Ӌ@h��a��m�k�,�������<Ad����,����5���[⼌�s�h��VbV��%�zϷ ��͐���������~��w7�R#,��U���`bVl��m���c��ӝcQ\�� �d��
J�����ED�����aetR��t2��g\5x  ���`*FC�vs��f��o6��QH��M���[��Z�x��WT5���J�M����IKv�+2phg:�Tv�;��9;�������:OIk���fM��5�h,�P�u���{j�l�xW��w]��D^�K�������`���M��9y[�Uq��B[Ł����fL��ʔ[;�w����{˖��BS;^zvJ�N�WE����kG��7ԏ��M'�9��fܶԺ��a  [�/w4�4��r�vo�J����qt�E�Kk,҃-nG�GW�*�ob� >�>F9#椖��+�8�*
H�c�����9��/	�����=���Z}˜/|RsӊZ���v�SI�!Xt9��N����\�1�c�a�'�8:���OeuN��Y��,�Z�/n�x1�6 �6���7Q����7���r���%T�..�Aqe�|
�HW��+�~k.
G�HO�6.ph���Jo5�ฤ��NY2C��t02��.�읫�v,tH2W>���fV4{C�6A��d'՝�#ֽPy�
�6����a�������&����$c*������AV�n����29Z�@VOrMlZ�F�%��L,��Tn-�*�mHc#p�ެ>�?J߰F�9��M1^[���Q����ԇ*(�=�(�w{�zPI��[�jŊ���$����h�R����T��J�� �(�W)ȽD4���D�j��1J0*
M�%��gۧ�7j6�,��X1�o�r|�+5ӭ��۷TCzl�M����p"��\A��y��P�4���6p\;αa�s{��@��P��C�pr�1 r3b��48l����q����a,W�Nc �_C��-�噾X�k+pPl�<�#}aT���"R���u�fȊ������i�2H˽P�X5��B�ې
��`oz�'��u�$��!�5�*eiZ�:����r;�-�[Zz@qW@�^hՔ��T7�B��;���|1�VG�tb^s�2^q鍟�1T4-�^p̞6睝�`<�]�5��iŵ�l�0dYf�_���o��t�Ti����T���lm}s���5{�߽w[�Y���RJ����O`���o� B� �}��Wp�y��Э��G[�z��V34��Q���fM�Z�������f7����w#Y�����^�̮�µ-�(*oN��1wn�mK�ȼ�1^h��7n��	zJ����9�ݴ���Gs���ŗ���)�\���gLJG��R+�g��Avs׆6k@����mie���}7���.T@;cj�Ő�.�� ����ӔT�)?`gC�vcH��<B�sK2x	�S�yvi[�!ҕzv�0��ۗ:���!�c�
`@ccx�}W|�-�96y��S�e$9V�	�"�޳�:���ed=���qJ��kM=�������v���S�t�U�V%���m<��RQ%m?Z��w&l��;���X.n�l�Q�9�8A��^��G�z2Xxu��Ι{S�d)����Yt��w$G]]�t:�ܗ;{�wk1���&�ө2]pݔ���H���XD
99�R��pJI���Ky�!����qr�h�}���2����ܙ�����|��E@�����;���;�o��"򗺻�vJsc;�4)���h��c��±�8��@�S���;�4����T�v� �v$c��o"�.6'��G{�;�1̛��6Ѿ%2��wh�P�y�Ӎ=㕝5\�5���ݍ[z��l�T]k��{]'ok)��|{F,� vTN�j�	�CV�MM�/���� �Cc�ؗ���l�W^Ok�@��[�YD��H�5��)�٘=ɾ����Z����r�xM��u�J��s)����D]�4��p'�h��E։}6���M�a���r:�~�'�>�/o.���t��'�_�ZJ^lUf��V$��R}�n�9�њ<��ϾK�st���8.$a�7z��K����Y��ƹ���"�����'��օZ���IE֢V��hK�X`ub����Z�Hy������W�9��}!�~3�5���4ܔ�G���Z�9�ǓE���d(�	\������ �p66�� ^ƮY)@]O/(���g9�6#tDŋ�k>����X���kG#�,��̞V/O��x��b^�Ŋ�{���eh�[HܥV4Q���X�u5[����>F�*L�)R��Z� �r.l���Ly���R��*u�m>)	�iҝ�!i em��8.�vW��w�	S�Ğ3kE�lmx�0o�2L�j�"�{n��q�+���y��$����.h7��%lR��5��FXŴ qL����A�i���(^{z��i��:��OI|���y�N�5�m��v�B6���z�H����Ա5�j����R/-^��u���SVPom(��&Dj-nU��vx�0�5>��|��S��S�0��KP�/WIؕ4n�;�6oh�Y��g�y�D�EC����wң�r�����$�[;N���-�3xI�
%R��-t[yp�0sn��[}�"�0�}3N�ogB�s�*��&<�[DD+&��6�����WXX�Ƭ�Աf���T^����Y}�e���,�oj�
�vW|�����
���۾0�u:{܅�1��/p���
�VW;YD]E��v�\�}&QO{i���/R����]}�w_jʎA���9���A��*vX+u��| i��Q��K���ٔT�A�1�=V��2S���(?l���L͏��o��n�hn�4bK7�1F��W�յ���^��Y��K�eMA��_>��S��s���zd�,��VVq x����Z�UV|Ζw��-q��T���6xt�[-��"�蝖���M����թl�R����BH��������ea�?}[$d��n�B��h��A�ͺ��k:7Fmm�Ḗry�tD:�2��n^27@=�X��qw��=�a�`��x�Z�
��eᏽj��e5�����B��@c�s�Y:7+���T-Ml_��\�^e'k�ݦ��B��,�x�.��#e�y���I.�RiKv/��T�e=9,-�5
��H1�U�A{ִyq�P'�t�y���#�ql�@�6��T8���&�Z�6��^)��>�$��1��X�N ���(�w�}D���$�|�ÔM*�=��(dɵ'jFe�2��`�g��LY]��=ёy��@�:��}v�'LᎯ{P��S�o����%���7J�E�&Z�r�qI,�r��R�V�Tɓ"9BQٕ|��W賷.���ޣ��έ�{�&Q1++�/W��׾���m��¨%m�Vڍ�ذ�7
ZQc-�32�7F(hfd��GpAQX(�q1��m�DVĥh�*�KQ����)�ʊ�(�(�T�Z*ԱEATe�j�V�UUU�5D��eJQ�K%iB���pPZңjԥ�����ڨ�5-�ƪ ���[j�Z�`���lER���mH��m* (���-�£Q�E�V�2����T����(�)V��6ʪ*l�Z��rڕX��(�YDe��9-�
�2����F����m)�q-V֕�meJ�Ej(%�j-B�D�Z�ƽO}���[���gD:m\h�b%��H���M*��{�g;�
 ��Bq���qN�����rk٪�_k��^Tg��)��4��%�<I��s2�4�o�������M�˖�|Ʀ�讗)|3#�\f��j��ٷS�ݮ�^^C�)�����wdݫa���3[�"��\vh�Fբ<�6���\=�C���s"���@;a��x/Sg��V��V�Vo��F���3��F<b�.��X��/���}Q���s���SZ/U�p� p���a�Q��[���SwO{p���|n� O1oY~���}���9�7Wv��=']����TA܇�vF��*��� "?+�{2�9�>���\�W6�X}s�E-�BsbF�Z!Q�9��𦇻^��ɦ��c��}av�zc9�J�'�2M�]Ӎ��[j)����o�pU�l�5NӢ֋0�[��􊆏'�p[��в(Gw�ݤWӓ1%]�%������I+UP��"�[�6�4����c��Uʆ	�N������2�O��,�Lɀjq��p�h���-w�"�j3z!�����:���V�lb�Y�s�0)�AI\^����1��m�x���xN���mO���ޯ>R��⮮��k5�A�ѵW��L��<�}Ě�)�]Pڲ�rA����s��edO��&�Ҋ����DZ:KM�A.����c�x1a�j��r�����A�����Li�gg��Y.��y��}[6ҧϴa���  ���
�����:	�l�hp��]�c$�#M,�1���	k��)Z��Ո.���_�G����t�����Ȋ�:4Չ*� �ҁ��7�_H}ؠXX҇�r�u�0�>fI���Q�����з1y�2cA̛�U��m]�w��q�fQnV�i(��D��z��`+����e���e2���l ޷�i�H�m������� 7L�3�뱽�b��:�yY���=bjr�P��=2B�,t�������R�[����N×���L�@+�EI��Em����m�C�[(й4c����h�Y�G���[xQ��ѐJ#V�쀣k�du��� Z�֗�fb��e�b��b�,��S\�R�r�,�#���\�f,��8Ɨ�#d;�x�߱86�Hw予�)d�~/�MNס�i�nנ�_�9*ɓ��-��)�M5�;���L�C���(��w��S��<�{���k��`Xj�R*LӬ弁]O3�� �XdoXR��\��;��o&l�2N�6��ڽ��0\�|Vf^�۵NN}�zE��9� ����$���R�J��ꋵ����f�����n7/���ji�.�^��o8�8x�|��dޅ���)�ACR��M�Uy°��uҟP��|����-(���ˉ֐���	� ��c��
�g!�R�UfZ�2����#u��U�Ni��8�Y7W8sR�Qs�;�|29��qF�s&�MWFMn��7��R�q���5&��s�D���l�Z�(k`Ď(Y��d���n�!oF'��ga���;8�L�yu� �ˎ��9�fޞg|0;?nl�2?g{uv�S��'�&�Γi�u�oF
T�w!�9B5W�Y..*���T�	sO�X�%C<v%	�;-��ʊ��y��^�+n>��s3SQ7'>�IP�Ǜ�,ށ�Z������ɻ��*���'���2 �2�T_���W*U�K���`�/���Ø��. ��{��ݓ�:0����Zj��Hq��,F�&0�����/<j/���QKA�zY���ssw��*��o��U	j��$�Y�Μ�i���ñ{R��x��������J�	�)�W�����F��b;=�㋫ͳ-�iJ�⹸���"n+��ʈ�0����Kc3�8�)׾�H�N�w8d����ˀ�Lų�;�{;�	́�T���X��ٻ� +���n�V�F���{�K�>�u+�Ő�odf��[i�R؊�q�N#Ct��PK-U6�f����l�[34�*Y`�d�=puN�T�q�Lq6��o#�Pow]��կ�1��AI9u��--�WB���Tu`g���3�F�D�,4�۾p�0�PՇ��*��\������o�3��a���W{}Og���6�RY��Y����#c��$�QPu���w�5Э�l\p��`�C��s'i��sg�9��o;�ד�X±m^;�ʾK�L��i`��EEL`ё���w���8��E�������Ģ�p�t�K�hi��L!J]9ܬF��y>͡eJ[vå'ix�n�0�贳3���C�&D�Zz3s�pQ��R9��b�����"�K�n����A���mbq�^��B���J��[^�(W�o��/O���<�AJ��%��]�i�vk/��a�8�$�tjTQ�{$��R��d�|;�'�o��e�g�I�7lS��-'o���ʊ�{�t�+l(�	f_GV�S|��Gs���:����8�'_B��d�,.��]T����-�_#���%���vV�fP'���vx�#�N6��@t(�&ŷ~�%B�Q�=���սw�h���q�ǚ �a'��W�w�pW��W��c��SO.L��32�umh�)b�}ӯR�n�ab�ƗI$u ���9��\��-�v�EI�2x
�E4�S	3�<S�C#E��0 -dƃ���,"�$	<A��C9���fH\����v��z��Ntt�[�"�V��$�#����9M��N1o����;X���Nob�J��^*���˧�k��{�eS����7)��Q� ���,�i��OUV��bi������t;���K]P�� �T���ܚ�i�wQ�Z�ccvo��5��S���~�i�JIP"�@-9Oz�!�y��	ó�/�'<�
�y��{����bv:��cv�ޒ�Hi,��9�y�Zu��$��	�&�����H��L�z�;"n5*N� :~�f)%���h���NG��\���gc��H�p�_�sf5�E��=M~��77�]o��|����jT(r��el8ʕ���M�dX"�V��c�U���kR���3���Z��B�N�G��#P�/���|����'JyKr�>#m[�=@��o=1y��[�s�x�P1a^�e4/�� 0�b��������b�Z�b��5�QKAt�L�i'7��Y^��:�IKJ-)����~�~?�Z�fm��-g��͹;��ٴgIx��|�gl���X�l���<�
���<V]�jmnȀ��`ަS�Oշ]�k)���5� B��,ʛ
[i2�����@��YK�X��,k��_z�j�Af�����c퇝T���H�]]��9r�8R��d���T��;&�:��KD�7sR��糓�&)`˼�vq��`g\}`I��.��:v#�Miu̓�E�u��!��<�&������΃*Y��=؁|�5��WD%z�Kk�� ���>ސVj�Pp�9�����.��gC�s��׽9\��b���ホ�/rW0#��ew+�쨶^X50�da�����˭��]��H)ꨈ��ʲD�� �Q�8B�4�U��nmp�{��a�qj)��F�^{Y��A!��s^T�fMd"����XxH�)��~9����d��[��|��k�2��a�sd�G/�_w.������C�w���e�nB��I��C8.ۺ�B NB����;g*)C yC���h|d��(8����aJ��G8e靆H���X�{HX�p��!r��z�LL�<To�0Z���\��^S:2�Z�.��)�Ѿ;�>˺<��oӕ+��Jb�b�� ^Ҏ�����
��V�������%
��h�3��nw+Cf��oF^�˺���n�@�[��s��u�z!���"�%N�}W.��Se�٢jK:��'x������м�-M�]r�����qK訍d╯J���j����U�8Z���6��RqH�n좜AEJ��ۅd����KM�]�-^m�|�$�4
U�ON�;Tֺ����˭���~SΏQ�n�*b�Yim��eiJڃ)D�-�J�K����0KJ!R��(���[a�fZ�j��mV1���KJ���F ��e�Z+Qh�"���!Eb��mj�TE*mK���Q.YQEDb����j�Z�kR�URcX����l��1"[c.�-�klmZ�T2�VR�
��k++Z��Ԡ%�J�����I�e"$���R�Z�QIQ�E���iF��[`�l��[5�R����Z�V��TR��� �,mm�TU�(��-b��(�UQQ��L��meh�XڴF�E����mF%e���<���~.m��>S�q6·e�Ү^�X���u�x�iZ��2I� RH���3yڕq��`����|G$�_uBz*�/p[[a>�Tv��~q�x�HIp{՟I,tnws���r�]��ˡ���Sh�QP�ZBUنw�gQ�撰8ԫ;[b�Tj��ngN��¿}3���3�q�[�1B	�$�W�bu���C#iZ4)ƽyƠ�$����'�(������KV�Џgf�
��n��Q��$�q��p�������:/^�v���4�B��[�P�q���m�͊}��n����^
����{���~�Ԇz5�O��b��",�[��*�S���ͼƹ���3>��PLśw�2��o���@_B���\�<�{��(y���c���{x��i���V�(��ޜ}��eG�[)l��� ~�'��B>D���+׮�Q%V����k{X)�O`ѧ����
Ywo�k�a�����b����ѵ�m�ħ7�̝�!\�-sIb����ᑀ*�o�fms��Г�o4���M��kQ"�twq�U�-���z��ҩQPyFo�ͻ���e��4��� ��x���m������U�+X9�C8ȍ.��
B(竨��Xr����|��=��Ǧ�A�/`�4���V"�>3�B"�73���+�-{i�:⒡�b�v������d�����/Gʔ��s"�ǋ��XUe�\��o��D�1��P"b�Q~���Q�3 P�O@~Y݂�8�gA�q�P�[@8��ig�i ���oV��7�����6���C�a.x?�<�m���g�=@����̷Y�ۆ�;~����+�j7p�U�@�ļw Pn*9�E��G*�{���î2����c#h�;��2��H�޵x@7K�׮�� �Q�m�u�5V/�$R�マ	�Z��������n�2�Ml���ۣ��u�0�&u���W���Q�0w$-5ܥ�85��\�-AR-c��QF�\�j�IY�1	܁z~�m�ε�L���A�Z�g�$��o�s5<�R�������,�4��Tlwr�	A��:��P�Qal]���i�v��x�l��.�E��K{k�n*����Y {�՝���g��]�J�J�c;(	����)�+�N�Y�A�n�f��Ea�Jlb�X�ʬ����}~q�x$�O@��Qr����:o#]s60NŮ���h�c���V������Z�ܩgj�lb憊�Ȇ�ޛ�^GeX���Ã| ����..q���iS/ 7P��h���kN�������T������e�ި��;�x�ڗ:[/!-Њ8��+��7��9�6��K:b	A��>!+z�	�8�t����q�(�C�x�:��m��T4/�� A>��v�E7���X��r����e�E,�9��� օ�ⲢN�6$��aSL*�(��w!�j�m�I��cpn�4�ލD��gv5�uf*�F�4U�9Y�22�i��D�p�r����D��U��'�cqX����%�х	rHI@��Fk)��V��kh�C�(U��^���ڍ#y͸��b�YͮNPڒ�����P�M��֯�U��`;\�X^�;Ҩ�vE�i�;y�gL8m���Q7w;"�[��0iӁ��EA.�69��h�z<��"�U7���"W�" 1���v�u�C�^�z@1B���(e����\{�4��
�:�<�2t-w�:T}�.nga����%�FЭk\���g@{�vkUK���ܲ�a��WJ�h�l��Y|�Go�k:�]�o���\S�a�C�wDcg�����,{�KU[���jH��5譧'"�Oh`�)xWZ��^3�X����úHW�;���+l�>j��f�f�t�K�{q�(3O�>����k����Q�\e���!��]�>}Gn�uxV�z-�Oԥ̚S]��Ư�Jfݩ�~�ў���Jޒ����N 3n�,V �2��fj�#���V�x���(�Q�[�4�smДdw*v<�sT��o'� �.x�+
*N�G ��}�CƊm?ed�؛����M���E���6!+���g��"��Kڝ��/w��W*6K���L�B��WY�f{8�	-	��˯W��˜�麫� ��UU)r�]غ�ˁ-p�8�0�M93�Frb2�������.�ϊ�AQ��,�t˃r/�~�~�:�"_g�d7ۈ1C��Tx�a�A�Ɂ��!èB�ԑP�]��*�m]Y�k��V���ޗJ`9��?sɑ*t�H�U�kg^ٜ��Gf�q�:Pm�8�S�9U�5 �:3�5�56U�\𭛇�[	N�ˎ�3�..4^�\���˾�>ܦkxM�r'؅�����+ԡ��SM+Z6�H��W@��_��z�mӽ2�ǀ���+F��^�cݰ�.J�>.�1a��a�d���r�l@k��&�x��=}�h��N�̸�`PƝ�F<�ne��(��r���%�z#�_kmn_@�P7�Ū"��p냗3}No(OQu�	�{�鈱Jc��ʌJ�4�ڡ@x�S3鹎ՒԚ��Nu*-�E]	�w�;&`I���ba��rgiՒj����i��j�����K}q�[qhژ��JD��k�_wQ��	������߫���Tϖ���be**���d��w��������,���}�(qof�q�<O�Xz�`oew[U���&c)hTa���G��i����a�`�O�����,e~����>t���ȫ��&�삇Z%-�S��9V,ɗ%T�T*���NB�f�ȍ@�t���/N��_]K�Ҧ�Թwk��^���P0����=�K귖8�ϰ��m�ot\���:�߰�oM���=�������܌n'D���F��&0"9�!M��NTT�oS�o��0��G|R��z"Hm�?�QQ�~�����~ 0��m/���}��+w�J��.��M�3�SRv���𾻜�s�;��y������}Qm�����N с�1����ѫ���UC�����h�*�k�K5��̫��tot
X��sl�L�+�7/�\�����Q��ÆQ ����|�{���pG8)�����"Ź��Q�pՉ�3s���-c�Ql�=뙳Y7��6��P:��u�(˛�����<Jj�u'��2����.��~Y��dڗ�!��gF"�������*&a�\���z&��Y�2��"9,�ʙ�.��>�2+�oߎAᕖ8f����Zy7��/��Þ*K\k�
�D����35|���ʍ%�ܱ���u����4o�A~�u�Ȳ��Ӓ(��]�s+��ٻG�a]ؖ�/W�=興mZy���ˌ���vT+�7f��X�}V�;Q��d�6���9�/FKW�]p�� �צT���SΩ���=�w��Ad���;���90u,S�UD��wÉt�b���KQ]1�6�X��� 襂���۾'׌K�5K���Kנ~r��X?>P~����Nh��C:�S��fg��ku�tD���O���GpKV�]�(�x=���� ��v*=�8uuƪ!J�Vܻ�.��v$����q_q*v�Ƨ�1|�3�KEK�yS���>v�ɠ����2���K���uz��*��S��g��ز+z�Q	�ʗ0�_��*�;x��纘w|t����~w���<��g�Β�+\�䩂������J_�l�@����<�A޲n�o����Z���[Kd�r�JLȪ;����#b�t���6��8($�A�oW�yM�!v�+�e.f�2q[��o����&��&!�W;z*����i�t�+�u^wt����%�[q�ۃ���v�$������cB���Tݕp�W#�a��=-����#e�w��D�:MJ�+&��Ȏ���0NC�{T�˫�c>�}��ʷ���|u����qp:�=�t��:yIHff�R�l��r�pX����Q5���z,��ض�lOm�0>��"=n�ڇ5�j]4.��7��X��3'i�6���wFQ"T��B^���OkU��}�������M�	�_i�*����"�-C8me���\�z�f�9Յ����(b(�J��ܑk��Y�`T���S1S�Y�o;�ٿ`�ަ&���N0ޱuS���C���V�I��R�8�FU�%G٧�
$	��^�nw��
��"�4}��ߟ,yº{����	p��ۼ�]�Ү���dđ���^E�dqQ��б�z��}��������Qg�M��kl���3&�"��fD.�2]�4�F��p��l��*rY��͕�R��O,�ܦ�Үu�6l�Pn��*R}�FWL���:q����M�[g�Ղ]ە��aU�ؓ�Qh]\o�.7	�y����.���w���ﺚ��@�lp�|���v�RXUvgM�.llΕt��"�ul�2�:�b���1�Ӡ�
��"�)�Ow'Yn�0�ltۉM����ӓ.r:��;(�7�{ε]j�����[����yS� ��c]k�_�����Pq(V�lJ�Z"��Z�r��D��Ū%���ҪTaZ�h�Km�U+1�+lR�҈R����a��LIU�mU�e�",G-���-(T��)iJ֖X�F+m`��ci*�����-�q�
-s3-�B�R���m�U�Ŷ�U�Rֈ�0-�j�`���%nS1�J�Z�TkR�����Yh�)TQ(�+i[h���-�R�h!R�DZ��[eH���T�U����lq�+UJ�[�*ə��,Z���Ev�aRz\�uq���O�8�\�.T�V�Ry�:s�.�h7:(��W��ץ��T騹�T��J��z+k���}��;�	4�x��w��+�t��*a'�3q71Z/�26����v>,�T�
�ӟ+�la�T'j����.�DR���\���;)�ߣ%NP�4*����)L�C�!�B;Qn:�Ƶ�."�2�f�%H�U"&�Y��Ԯ B��G��E&���ˆ..n��rD�����:�>C;�(Y�x�ճ>��G�v��W˧ho��_��B��\�����}t�6��r�VG��W�ӝN�s�ߑ�>a�H�1IW�I���p6�����J���ט� Y�S��9���,��X�B���Mк����N�~ź�b��Z���;��`\�>�9t��v'p�FW�C��I�c�����$��r�b8�	��gq��>a��E�#���諭��qh����7~^�293r']z����f�Sx�`��$�
�1��ww�����:�J�^sSH@��]XG���>��2�����h�n����kxL��+��c@H��'��d���$3{1sb���̆�:�༨]{Ap�O�i�z�ׄлO�t��Χ;�Z�Odؾ �[:��T1{9�֮���=��XN�ʨk�.��-e�ہ0��M>���S����Nz�I��ˀE��0=�ΪB.7wM�M�mz��}�Q��:ۄiLT�SҤ�kz��o<Eo���K��X�W ��53.�RThb�r4DJ!�K�{:���
����6ϙ�՛6sL�tsh�R��Y�@��8K� ��I�|�]����of���ŅmԎ�%3��v��C��Y��4��&�xƣ���IT(wI��p��Yzer�
�˞�/���ވ�D���7�� �К�n��.��4`�Y#�Y5S<\��g4�D�7��BmLc�\Mʾ�����G���5i5;3{�y�nݥ����g緎M�,�7w:��٨��gF��y4�!��W�<s��?cx�v�H��(0�W{V����� \ɛ��^�S�&v��6���z��<4����y4߈4/��s˧���q���������bE ��זM T�=��
�}��{5���{�ߞ{������%AH���Xi �I4}Mr��1 ��<�Af�i��ANj�$���3���+����C����PY��~��}����{�w����
E����J� T����%a�l��!�t� ��z��i �o\�i&Ь5�$�M}�0;jAACIR7�Ϗ���y�ܜN�q��ܡ�����I��^�z� �P�JÌ*i��vi'�VC��AH)�t�n�
�
��*��*x�YY�ןvv]߶s�sϺ�{ξ!����`V���AaƠk�bAOY6��,8��
�QH):՞�@�TOn$N�S_s �OP�,�+�z�ޘ�y���ʁ�.���Q刉�q��1Ǭ�l��̭؁XLR��Pfnڼ�ήC��=4~��Kf�|+$h�&�GV�q@�z"""#9���y�~'�;f�g?'��
AO��bT
�hT�@�_�6�]�H/��&$�����x� |�!�H���P��Ns�����߹��!�AI�ݜt�3��l��Xm�O{�cmC��H,�FT1%N�I���T��z�!Ӥ����bm�e���y�u�;�~����$��Ol��_Xt�&�j�)�J�]X�0�1�1
�Y3]d�A`zԚB���l*c'�V�	3;}����}��CHx�ԓe�d3�M�v��M���X
��&�Y:�Y<d�2C~���u�o�{��]�q+'űH,�L>�J�R|�N�m��2V��|͸�!ެ�AH?S�J�Y�qN V���'�H)��{��:>u��w��}ri8���'HbM}C�Gw5��U�!R
�q�c>a�8��H,>C�]$��LH���s&=S}�UL:��"���	�r�d���Y��	��AI֨bt�P;J� T��{��Ă��'L5"���V�R��16�!�<���o�~�}o�s��3Ԃ��-I�*C���T��I6�a�
�P:�ba��B���Sû&'���j���*�R�k��+�޾�7�>�>��1�x���q�t��+Ơ(��"�ҡ��&$L��M�T���Z�8�Ι*ty@Ĝg�3���$��sι�>��=�s_N�*T���4��Vt}dĂ톙�Ii_X �}z@״���w�LHwi=B�+XjLB��M�1���s��;��~�o�"��K�Cw�=^]��B��%cJ��Ԧ�j�<��*.,�C���r�"��KO��Y� ��F ��x����W�_}T"�|�����1 ��8�H,����R()d�Ɉq%M���i'hVz��Ă�U6�N$zԊx�R{�� T�g_]$���]n��{���w��o����z�`|�>�P�+'l�6�����M!R
jya�4�Xk�:I����a|>ô$�
ͧbA`�P��������_5��s|:AH�ĕ���
t�YY��B���$<�Yq ���� �i�:I�+'̨
,n�Ơq*x�"�X{�]��_=�9��{��&�*N���L�2��J$�����AH��¦�*T��Rx�O�+������$�
���ή'�t��sv�w���|�w��=U�uG�`z�M}O� �HT�[́��ٶ����4�Xj������AH��b$����)=B��k�H(Z5��^u�~s�öi'�$�ى����LOP*M}��mx���ڝ�T<J�T��a��2t��R�ɦT��;�z�'�T�}��[�~��y���Aa�*)�I�,;a��Y1�|�OP�)6�����+��z�[�*��Nَ$}�i ������޾��$��&��re& (�f���@�>�
E �CL��a_P�O�Y�7�4�Rm����d��<:�bq�C�1'��%���k��]y�=�:H)���礂��t�����/��1q �5i��`z�!�SHVE��OY���C>N0Ă�Xp�x]���������"���)�W[� i'��oܓI&�+4�N0<j
E>@�L
��T<���Y3�1�'��AAC䩝u�{�^=k�3�;P��,�VIY�E����M�yXK�^�_e��-�;��!ʁ��V�n�q���r<E�i���q�R5��CeN��D]梗�{��CK;�O�"!H)�~-<f�T+'̬�����t��+1��ÝXbt�Rm<v¤,C��:d�)=N�PҰ������<��|��y�|�3��6�R�a�$}iƤ��+'�$�;�Xg,1���k�b
E �&���gl�d�+1���׾�������w�T��I�L풠�^r���J�>��J�N!��4�X��H)�h�_X�&%@�Rt��$�s��ƣ����}�wZ�����z�8�a�
����8�I=B������6�N �PS�hbAC�z��@�1
�=dĂ��Ԙͤ�ĝ���N�7�����������x�R�T�B�>���'5�<t�PP�y���S���zΒT+XVO�P;7L`tԞ�^��)���bv�R{���.�����w�q��V��H(t�����P�LV���c1����;ʤ����c��T>t�Y>eO>q&о�b�<�^o�{�>��w�;�M�;k��b
EiY:eOP+���'��欘�Rwݞ�gl����S�
�:�@�O��vH�K՘��������3��y���~�z�h)l
�@���Ü�!�Ad��e �:od�AN����&0=jzξ�C��!P:Jæ ����R,����u��y�A���Z�6aLDTǔ��L��� �Ձ��N�C�"�a��i ��<�hT�� Wl��0�=t�PP׾ᤂ�uM��IP���k�|��ߜ����d�*O�C�'����AH�<��'h���V0�4uC
0��I"��M�Ұ�;I��z�{d�1 �-�_y��w�kZ����;�/:�wwu�,�,\���@�Z)��D�5$��VW����[�{zJ�u��.��,T�1L�ܕƕGB��v���o~�~�$��9y���9κ�jAO�VjAa����'�$�;<��
�kcֳGvM �Rq
��*m%E'�VM��M2bAC���:g��>��~ۭo}��i �;q1��
� ��ی�e���{`h�XAO.���� ����H(�ۦ����!Xjz����<�^y�{��p�&Щ>�0��`h���AH�ݘ�H(k�LO*O_c;d���Af�t�teR)�h>��AM�זi&Щ�z�����~����|!^2i1���Ă����&�
����*�d한d�Z��y���Aa�*bu'v��aP��LH(tϼ��3���y�lZ�PX}��=IU���s �4ϐϬ1�$O�̰+R�x�mH,�%M�x�j���
��)���d�b
E��]{���\����N�>eLC�i'hVO��3L� ���+������&$���f�H&��n'*AN W�8Ì*
E�ܢ�Sh��������w��{��|M!�AgƬ�j�Y���\�a�9�����B���QR�QBs�c*��ȱdGIݾ�M��>�=�N���S��y�pr��k�y�T�~�W��voiegM�.]e���h^�ۺ���Uf�6�Oy���Hl��&_�f�E��d�c׌}�#m#���أ�8%Z̧����r��}�s^��s��zܜ����X�/{͟Q��n�l�<a��b�S�\]�h�jS��Zd8�&b�Bp��=�z(�fLE��!W��(�G@f�Gn�y�hm����ŗ7��2�_�!WJ��& �̈�6��P-�l�;b���c��v���_x�٬������1f�΄Ċݤt��3"�qqu3�s*�j��z�Z�-WI�N�j�o>)���A���B�l�M�C5���e��=Nva���v귒k�}�r�k'?x�S�P��~��00������k�e��a9��Υ&`ٳ&`�7L�L�[��*�Yb��{ro����3�GD�~=t�7g�����G��-��C�+�3������W<�[wP�̥Jz.��bI����8�+0c,�}����mq��@Uv��x�osϥ���ֽf�m�[���KA���x��s�[}��b��H�]���::Fd�X�6C�d��o�	�gF�!X]��G��z#m�[l�ϠZ�50s/�7;��S�S�9>r�%S\ETeR-�0�ÉSj:qѝ���Q�`�	�v�c�PĎ��	�l��9���=/i�֯���m�۾��[h��	ٙ7F[�W��Dú\kdL�G���?`	�����r TMB��g�w�^�}�����@�^׈-�+SA��Ul��E�˘��W�L:�R��\�JO��wV`��o�)Y����]�ɘ�veτ�U��m%�������Y���~6n��T�x�/�:�p-�r-�>A vjJ����M��Rd�F�H��^��rr�OiW��5��{p�(:�0����WR�;1Ҧ��1��:u�?^�k��=��e��dT����������N5K��Z�(��X��
���̮(ǳ�����.���:���l	�����-,¿#��z10Bo$9��C���v��>7^+�I�7�q��uvm7���Y�D;���W�z%����C���;�
�ؤp�K�)��f����2�zn2mP�U;0�*ȵp:��˫P��`���o�Q�
�4��]��coj�.*T�>���˟8U3}]1i؜��W���.�0�5H}��y��g������̣-"?~h���w݊Z�-�7p�ٟl
s6neZ��Fτѩ��qԥ	�S� /r2]���*tu��<h�F�n�GX�����C���ʄ}̗\m��LA��W����3b�٬�9�x�J����UY/v���Y1_i$�����G��K��٨�Z+#�2�5���Iݹ˶����U��~Mķ �j�v��T��FvV���� ��۔#�'<�;�Cv�D��jZ"��oD
�^ed��XW�N�]i|/xd{5ǯNLDhT��L����HHN�9�����h�%�j)ZsDA-rԨ��Emwr����9�O�w��¹�̇�#LD%�ƛ�mή�CA:�gay0���Ў��d톆f����.=����Î�o�øV���D��@�=�!�v)7wS���pٺx{a��@s�x���e=`�7��{.�s�)�S: ��wVe1�JIg3�5+��s2Jξn\̥G���%�ںT&��/�|H����V��i�ϯ�֠3�  ��1��7��q��.��(e�79�4']-a��f��X�qJ���f+4L��w�a�qZ��M��F�5�ɐz_�J�琼�Ⱦ��X��&UuȲ�y��@�����pչ����?�c�N!sVܮ[|f�|��Ҳ��qN��T~�)N�[��;�6ăi�wQ���ˤe+��hրq�}ѳ �l�V��`��M*��zt�L����Y�#��>�E��Ӫ�. C���e.I�Z޼-���Y;[�"<���B/J�u���5����Ѹ�r骘˄0��zp�6�f�1F�ʒS����˭�c��:�]b��[��o#��*�rf�7yÈ�W�ڧc��VP=�"Ji߼�:��6��ן�T��N���L�cf5w8�0��&7���91�-²@U>�(�Q�Rcf��IٺD�ApJ�%���c��@�r�] ��x6V��_=q5�םo�{}3Y�j�������ŋG�f�
[D�V,��U��R�+F-�#��h�J��E*Zت�9C-�LeV
��DcfcY��V72-fZVbL��h�����J�G1��&�X,F�ƔkeKs%p��1�Z�(�bT�[UEa-�̲bc!QLE�������3.J(¥B����J�-�R�6W+h��s0D��X�[JɍE0\�2��`+���IY�����U�H̲T�j`�1�`V�E������NnIE�E���$FD�r90ȏn��[ʶ��(%�{��DCKP<�}�r�{z�T��.��ً�u],W������Yv��{�Ȓ6����f�'	�L\�E���Z��	H�%nFT	��YX+���3GQ�/�TAH�r��a��Bo+���s����,5��mP�B;�v6ssI�>_-�u3U���c�F��?�u�-���1U��{9�y7E	�02�T��V�ϲ�6y�ȝ�F��K�6�Z�N�����&\�<>(;�2��!�<ji�=ϛ['�V'�yu�0���9�������Z�֙e2鬝wt�R�t�����~W3L�Һ���U�0���x�ݾ�WBu�ɋ
mL9���ĩ��*S��(6l�]�=��A-��j���6�kR��w�ՑX��:G��x��gnģ�V�BG%��CS��{!��!$�b��V�6 �5]|Պq�J9������c��~ٞˏ�/�zb�.�Ŋtӛ��u.�iM�Drw\_���z�_�Q�م����{�
0��dH}�G�2��i��T��~r&�\�M����K��9Ok�30w%�θ�[���t��z�����xh����>��y܌kg"�:T�0���^
�,Y��r��<���+����;@0Ғ�f:�g�zo��Ź�N)��(�E�k�W;��ԁ|�Ü���YU	�t��T�t���r!,�m��ť��L��`л��z�![���|tu�h�v҉E��T3XI�b�3R�(��9���Y;0�u�m-:�?:�r��4�wA�{u!�o����� Հ��ۯ�f��Ǐ�����³/ua���4��7,�亳���[˸Rp�|�����C�T�cpw`*:n�����:�o$�`��݈"��z=��վ�鏒�S���X�L)�t�d���@���ȭ���������GV����1b��b�1xne�t����=���V�L9��.��m��*����j��n��Z��P|�N���U�*z�@�g���p��^U
U�����D\�*�z_���ߪnv6�b��*v�!�6�Y[��or/�&ǫI��5�{u�)�^2� :)`�t~�x?Q)�N�]z�P� h���ʬ㨊���+(ȺSs��pri�k��S�37-�@�R��hL[�Zkf�L���f4Y|T�t��	��Khiߨۓ��C�lIʋ�P%S�7k��g��ꍻSswj S�W��&0T�{{2��bm�����*�6�����EE�4"��}�]��^T֩��A���
N�u��8Dfݔy`Er��,��A���H�}\�I�9�U���ǋ�m���S�t�ɺ�ɹ麯�U~׆\�Y]��-H�}�%�''���݃frr`
��ss3.s�P��3��SC4}K��	Nh���nnH��^��Ӓ1N;�-����q�
{j5�)�TJ������ɘ'���]�;msH�^ј{Q�ꌕ7j�Κ��C�y�y��%G�+�=��#���Ȼ |w�j���L���л�ٷƗ�����k]���3Bg������;��'�B�v������VC޸�.*��7���7���ϥ�WAVRj���?>�7iT��3�H���>��ac0��s���͞o��︐%���p�"(��4o��<��{����ݧ߻�=&F� ��M����v��ޞ8�d�7;�:����/_:+ �ڟ�˨Wڳ����m��g��i3�r^�q��p�K�G��%7Crtњ��=�3��˵��]��]�C�z��L�_,�;�_6��9�Qs�Оb��?T��*�5$TmGقMp\
���1���z\�Y/�:��.gE93r&iWk���	��?h�/)O�u�����������'�T�i���R����%�����u����<(|���t�5۪�߸�DO����Y�Y�6���g+�G�����g:rra׍�s�g����u��V�+�6��)�5.��Gh�^���oZ)m{n�T�yFyTF�����=Q��D^�_k�ՒIj��mBꙇ60��5�������Fp�z�M�V���w`U��u�*`/9�5e���w��Q���%�w��S�2�����L�4t(����js^�q�T�U�!��./Z�q{��*�f�*�����#�����΍.+X��Z�i܎b�u�����M'�T�H���)ʛ�Sn��ϳח�''z��eW��܌��F������L�J!��uT���ʑ+j"��^@�����è�q~��>y�Rچ�f���WU*���k��T,��^�Y5�庹�SNa:�j�LJ�R�#�n������'�5����%�=z�[��^>n��.������iugNĉn�a����qP]dI�2�3�M�ֻt ��\�S4���~� �1+�o�|1��nP�Q��o���tn���4`��K�pW�.����u9|o�S\���ܪ�۾�����W���Gj���0�����0a�ӛ��Z=~��k�4���Z�;uQ�U�R��R��e���ѣ�,��to]3AV�>�+>���6��k��o�]�<��m3�X=����SL3c�:���K�h��r���MaG�����G�t>a���nl�D���}[�p���M�E�ʛ�}+*"�������U��iL[�2(
������sq�V5qp+�)L&(ܮ�89D�.^퉅44w�s?q��Ա�s���I����4�t�
2��VU.��3�� X�l;��yH�n���=?]�נ��A]q��S隉����LtӴ�e��7c{z��;z�:��d����6��ܙ�Q��\�Id�dJ�q>�Bc"}`]�Y
���vQ5^𻏽��rxQ¹��~"���?Tf�d�j��j��a�T��<�c�罃�	��K����/�S�s�Y;=1S�P.�3���2��F�%�j�-��QB`�tޫ3���3�c>�B����G�>Ҙ�ӗ�V�V��;�ؔR�k.�t��sN_6���\w�@Mh5f���1W@�^� ����1)?>�G�,��&~Y�qә��)3q��*�1=1���(�ږ&���FdJ�G���3$e��P�O���u�@��B�S7$��}���,���Zk�������r����5Z�!�1vnc\x��m��j�wkQ�4�h���U�����zI�{��pѫ�����ѻ�m���ߜ�:��xfm�U�ҳ�3��;;&|���Ђ�gq��ߴh �#��� �A�>�3s�r����Bo��K�$�J��D�A�F�1���i{���%�w����C������Ȏ���Z��'��2��+�[��ڇu"iTb�4'ǲ�dг+7/�sy������~:`�.�p��A_v��t���BZ�8��G�'�%�Z-p�먳��@��/�l��0�ҥ��:S��H��Դ�.�e��:�
l`�E0n�x��J�#��w�oh���mڐkۚ2"�#hIݛ��"yT\�d܊�����B��q}p�F�qU(ўB����^S�&^V�m�N��y�~�7߈��D����Yb�2ѧ�%jL��T�yڿ�s��ٻ�ę�3�dϜ���B(�DJ��z��G\+Y�|%L��J����t�y��x)ǻ'N˸�MP�N�m`�~�R���9qa
SR�EQ��,���ied���]�[��0,����J�~�	KFVv6�ONNK5��d�
�d�d�\]��
ύ�Ͻ�Zs�G��`�O�W����b���n��KB�hVݘ+��&ڠzD�FW*s�<(Iq�z�g�Ag��s����<R�^�z�n_T;tPP>nT��ٷu�5sX[�J��E�̛~���"�o) O�zbozl���/���2�J�6�͓Z�ѣ�+�DD[h$�t�گ�>ߩ��.�x۸�3H��+�``������Ys7�'$O:��Y&D�ɋj�
�ݽ��n�ŋ�G]�B3s�0v�m_|����9cfi>���$��;7�F�{���P�r�y�6X��e�H}~i\��Zঔ>7�9
�����P�>z�;���wP�<���"�-����EC��J���[w0�L���6��R�E�-WOKݳ=1z��Q�g�!݊ST�3��}5�_+��fN+����ӿ����`V
9qqWF�Y�үw
�NM)�tjrEa��NxO��bT�4~���V�W/.��=g��wQ�`s������n(ɘ�"+ѵ��N�Pf�0�"?N@��/��뻉�ձ�}��9;��0�T�ҫT�b�_�Ƒ�T��ݱ��Nɣ���&ޖ�����3�v�`�1��
u��*hs�G!E;��zsOȥ�1WP�7�1H�d	,�\-앀$���ǆ�� P�E�׸;޷~��>=�i���^�ow�D���_( ��Qc��f��5�+!��-�OM�������g�c%���S��6U43Y��3��g]sG��Ԙ�eثS�Eixh��fS���ܙ�Ջ����V�rt�i���d��탠���s�������k,���K�5̐�d�f������i�b��,��w8�4ZY��l�X�d����.���&��׹��ڻ�N���紕J��<��\5^�:&i�r��]
Y�X��%LIK�N𖷲a��l�,�󴡫�N������������g���nWkHQoi2����MV�.��9ɰ��y{��4fƆiکϔ�b�\�U��v�: ��m[j
�"Y� ��Oi_>������#�Z\�7Fz�o�է���x��]��ͣnI��>�b�0i.�y�{N ���P3��>���F��MK�����]n�g;\9�^�|ଛŪ8I)��j��J�Ms�~���M� �t�"�'�ԃR�b�E���:5g�]җA*g�n��j�H͌������������u�S�n�F�M�e��W����a*������Y�RZ�\�^���_F4n�X	��wѠ�f��w{ß�!���i���,���a��Vog0�N
n��� �!���ڠd91S�[�򌈶ܙ� �X�`%�8b���7XwX���v����t\w~�N�����̰#��0a�>πYm'V��E�q���LrլƤ�a��T+1���f4.\����ۈ-�eF���YP��p2�¤�`���7-��.Rc1l*�����Zf[E��b3b�
��J��
��(8�ۙDV�R,P�[B��h(,��Y�{��)5�0\qe�2�UI�b[aX�i&)��fb嘆 #*J��sZ��J̶T&$R�Qf�,�X*�I
�)*�����E �P����ZgGC�>��p��A����g,+S���L�KUJ�E��r�Q+���ă*�:���pe+��2g/���/n�{��MN���絻�&leN�)���3)T)��Xi:�>d���E�VW����Q�����lݴ����۵�H֘�-f�Gn��nt����$�{Nn6��O�6��]BD�Ź�N(;�pI{ߞ0�uz��0�B�A59��&lV���U�&�C�#<d�	鞠�L�L���5qp+۞���2��It.��Rj��{{ؖ ��"۷w9��m{��Mf=`"vc\e�X�/�SsQTUx�ɜu^�����lE��ieT�n�\=�\U9�����ԩ�0]3Q3�9�Y8���1n�}S^�l;�\i�h���ܻoˮ����3g�6{k8����JsR���	���;�����5�H'���:e�Ws�\ZΛnJ��B&���Óv�FIq]v�]�; �8�S�ﾬe��f���+eL\O�S�������7��F�!<o�Q}]3ʔ�����*	Le���.�B8t�B�iǾ����C^�@U
���^غ��GX�u�;) ����K@'�v�}ɕ|����P۩t��x�wJ�:+�{�3"�p �C�n�ͬ�9��f��jD�rꋬ7[^ʺ��VTȸ$g�v=]���/h�~�Ffle��
�J}F�úT��~��vO)~b�!F�q��Ƽ���z3���{#��v7AMVT=�Sn�a�mP��T9ـ8e�s���&&X��ӕп6r׸�.���ѽ�ʵH9ʯ9�u�+����Zʧ;>S�'gݔmp�7��t��)߭e%�!�D]�c1�Ѿ���څS;0Z��ej4�&��T[5yz�b��t��\��(��ѐ>�nIn�f�<X��5�嗀���sZ�Ջv��hj����Z���Ϡ��r'r���5�n��q���FI�J�&3�j���P��Ox��C�2�:{��`�)xW���G�h�A�%��V��%��ُ����Ʈ�]�]��P�W�L5ג����3��ɫ��"��,ѝ��A���� ��Uq��l��,c)sX��Ҹb��-V��șf܇^��ɭ�'b��U	㵜?Q��k`�ޘ�J����»�V��k����� ,}׫1;D��:�yfc�`Ί-ߜ�,�s&z`���E��G^����=��u����M�ٻ�ɘ�S�dϲ!��D���j�X���S����o1τ��72�\T
J�R�9qUY<�^��{2E{j��k[�2�xW}�?h�]�J�ko����>�G�в�$Tm�.�9�=΋:�-���@�6q�r�أ�$�afD܇�`�hk#:���)4�.�Q��h�K���ef���٩�Eź9^��q3R&+�V����h����
�|�Ow��}z|�ܮ�}I����Ӌ{���xv���<��5���W뎭�9vĻ����K�3�hC�U��zr��U�"D��j2X��B���ç�3KK����쌯�fFT	����>{^�Zv��^��ѫPRO0�����\�ۿ^Rmx��-^�Y�){*N�:�d%��4׃۷@�>��s!�ڈ苡7��U��/�Zy��̟
��)>�R�<*`/<������w�j�Wz�'�	�1R�O:R�%N�S�>�����n[�ƓKj�U�p��Ø�j��7P�����T'�\�Q�����4%�eu�>s7��Y���ŃiJ�{����B���;�ש%�]���%O�Fl�)̮q����6�D����J<�Q����w��or"���m�L^�_��J|UP�.᪙�&c\�l*���z��qW��׫k&�2�V+ɋm�g��w�w'*�g��S]51rM?����F��.]+o�ǯo�c��ŵͲ��a����Έ�7
�f<�ف�[gO
�S��Մ=��"��Uƶ�x]���^iCv��J�?:�J��?+�h3�ʽ�2��
b�Ն��у�/��_h�]�:����s{b��1��M���U�3G�kƑ��Z��Up��ӇI�Su�CiNI��И�>�뗕�v�_ѣT  �iy�g�<:���.`���Ɋ��+=�p���M�9Sg9�i(����%��`�1phL�[��a�����{�?����Bw K ����l�gZO�-���i���Q�8��V�����q^�J�<O �GTEl��� �Ǝ���Θ�+�3�li��_��G������u����ؘ3Srq���2�k&�j�r�myq���
}����-�஍N3�_���.�/�(�M�)ikDۉ�&vc�_�R����W�J�SX���e�YW1���"���{r�9Fp�I�ᇇE
$�O����1w���_o�!���٬�__Aª�J�<^���u\^��{na��r��a��p��
�S}�*h���qhZ)��z��U
��q��TE�_6�� >����眥��;W��]_�&�
ʔ6�];9�����%�:��bN��t��߷e��f�|d�M��.b4�t���v��	1�F�q����ƀ;O��{O��)�H�-�=޻�n��w��Dw07 DJK.9_C �i_0��6����U�ؾ�r_h��au�g!!ʛ՜��-s��Wڊ�"q���D��ޏCǥ��k�[6�f��1vo]o�*3���NNA����K�9�W_�HUc�������N:N��*k}�C�{@hga擼ΘJ�����n��ƚ�^�.g��v؝���M����VdR&:	s�+�v��2��M^3s+t��󅰑��R��6�ݴ'$J�胈�hem�ե��8Lr�ɏ)ט��xu�]l�-�1O�֯n��Ʒ��9]ڲ���S�m̿Hʎ4Fro�ṷXY�)c�0���+���+k�_���FO]��ߎe��P���%�F�䙍�{hc����*����_]�^�����Xcne
�f�E�}<�$۝�Z�F�u/����5ƨ��z}�^�Ami���u���M�N�65�TJ��'�8÷��u_#���x����M:@�מ݉���Ӻ��|N,���F�+��7z�3.,�4uv쓈��(���{[-��yʜ���C4�C�^?z�U�4S��#�:����|�Ӓ�l�ڭ��w�*����nUW�T�yT�)Sl�)"3)��qT���P�U�>�U5]����:���&�LiJk���z��<.��Q�[a
6�K~�R��U;���2x��ݹ�Z���ʕ����f��UX+�G_�:������Y���d�:�{>B^p��U�_�}	'�h�,E�WM�=-���\t�&v`ì�*�b�T��(=���-���{�L8ʁ9TdLL����_�՛dmv�����1���v��D�*C�Ӓ6��߲|�)鎓'�Khϐ�ᤵq<�ٻ��U1n6�S����~ڴ�{�X���9����������N�x��I���1u��TQS�X�b�w���;�Ev�O_��{���ǽSn��S�$���|�*�Q�H[�ޕ˺:;4p1��r9��W�4w�i���\G���f݊lͳs>���<9��Z��m����oX߹��*�����xc�9Y"�́��O���J0m���9��싆�*r)�*o(�r��^���^�H���I���؞eY�S����}�[����0�Nn�ORҢb���Ԛm ל���;�Q���g�;�Kn��w3^i�BI�a,�E}\5^�z��ՓY](T�@�f��}P���M�������32�:S�!%P��t5�k�˭�=3}������&f��j����܇�0j���	| ������������׍_U������Pݻ�����#ݱ�� &���3=3���\���P�,V*�qF���ϱVJS,eí��{Ƕl@k*F�8T6��.WַM
��U*����/��0xAl�b�Jώ�����8�6�z�t���ђ�VT麺w#�興��ۙ����ݣ?{����s6������\=Q+-&��
C�7+&=^F�`x6���b]�����^go����[Yi�眍AU����vVu���.2rb������'pdq�8ܩѬ+Zx���Sÿ�#����x+;� ���Sq[R/$�SM��Ab���ƺ����LW]D��+�"�L���y6�6���N��>O�po��g�Q��y�LYVU.��U}Ji�Z���K"ԛ��.^�\<��ʘ��2��IU
c2�W������=�r�~�����EmR�։v�j�s��wa7���~�s��8eX~.�bm p~5.�3�Ћ�[[U�L�Fe��\*�7�M�,),,pA}�<�^i����s�t�I�Y�Г��a.�	jպΝ���D�|l[7j�uՈ�rL�}[܃fr�v�5��g+�&��!i��5{�ύ�}�\\Z�p�L���-[v���udQ4�<�'����J��BĠEg�2����͢�yle��RʺAVEN��a�[�lw�d��J[ul�s s�zh��Y�	5mYۚ��l�ג�L���ClZ6��l�B	Z��R��,:�cO0��uy����;S)l�Z(��J�*�ܺ��B/������1+�+�붨�$�U�����w���̼�@�=땅꧔V��l)��ⶐ`�Û�+
U;8�.u��ӯ�3N�#Ea��tDp�zYÃ1=I���:�����ڻx�C�*/��6F��p^�����q��G�UcI�k��h�X�xA����f7(=�4e.ʻ�S�_�X�HH��s�ʦ�z�ǜox�C�6��V��NPr6���McI�=z�S�BL��FE�V�x*�M�6�5+h��o�Z	�n�AIݹ�����hY��ԧd�͉2h�E�ӡ�0��w)З�/��	��0��bÏ�Iw���To���.��Z��8.�qN�j*N�\*;ʎKP�)���<��Xt��Mo��P+�� (�\k���"�n!����s�vW������^�@���3"5��t��b+v��\ft�H;T�N�9;s ��Ga��:�E�Ft��O���/q��DQ	�OsO��vY��bN�n��d����U��Д&U��	��%:�����C��ܕ!.�P�WIn�1r��V�p�\�J�{�D��*3nK�a\����/B�3NT�"����]Zj�z��y��h*�ͲfPؕeB.1�9@U��4�1��H�Z��Y��k,�4�%�b�Pe�R[dP��%I��4����Ld�X5*�+Rcc"���V��Xi�YXX�e�(ň�1��dPXTl��LdRVE�����`�V���ER��fP+%eAH,SIS6����i�I*�l�LH�(���t�+1+ߛ���4�yC�M�`�r�1�פ<�E�Hʡ�uY@U�.�̕���"�����L~{E��U3p��!OJT���AM����Y6we9�{\>�}j��꿽b�U��V��F��0S��e�,x�Qr�ٽh������9��S6��Ke��_��թ��L����Y>>q$QFa��W��{2̝�+���~�g<2�ȨR�̑qs��@�=���v��gx�Q�i~32v�~ud��p�<����M�RՓ���eC5mVL#Q3�B{*��.ccX�0{6mQ��7�#͗u�R߰媜v��@kG�f�)Y�bC���H����qјR%�@��9�����4Ex�����Fh��[��׶Q5�����Hm�A�/	gY�~�r ���l��������u	y{(�Kځ�
rD�U�W���Z"�[��Y\�ʺoh��{*����Xw@�TT#v��ʤd�ˆ`6+=���:<��$r�n� o.f�!�V��!Y]�%��{����[o����A�9���&
�l��9!���<%'��i�U���>�[��g��fo����{/�dLde	8�"�nn�i)��t/e��d#Y�W�3�ԇU1��=�95�$�ùsJ�Bx���vZ댜�Re����ƨ��k���L�m0���t�lz��^\���
��C�ƍ�꺸]��AH÷�{zr���)�<~���ڵx� v�n�ػ�r�9UQ
aL۪8��aOq���׀�(U
�g��j?�/_��5�F�X|�kޓ�}/�14R��˻er�Y��Q�k��R�㋤[s@4�D8�6�MU\1nq���p�tI�7P��TL��]l��{|���Sj��ʜ�^�&���W��s-���w���+��k��`�ˮC1[�pC)e�|U�8Px����l��� ��K�W�p�*t�*���;m�Pf�u�ɒ	�7L���\,�E}�{��D6�S�*��dF���rgl�ì�k�+f,���c�C��CCa�W�0�r�\���4"xM��qۑ��l�J$.io6��)b�ߡ�ف�+�>J�f6z\��>;&�8H�7E�
�	��u�t?v���x~Y�s��og��e�@���q�p�D\r�d�@A�(�Ϫc%��c�@�u8W6.���h�(�y�Y}W�>9Y�?2r����F�9>N�\=��.����Jn%J�%S�>��k�.z�"����i�U����x�|�m��/7N��{�ELP�[gO$��p��z�*ccE�ؘ�~��>�t�-�Sg��7H	��3*a��t�P�ߜ����rzW���3naP_GI�h�'6筼��D�1�7�U,P�[aq�7�M�9����+Ym���j�ڲ�r����)��e�Qk�%�ds���-���s�P��.O�Tz"AsI��És2$*s�1Q2��ߠC��dz3�߽V�?����V�JPw5��ʨ`�����Wø�q�UN\�ұ1}Nf�.$љ��j�����6V�b�	�h���Ә�P��S�&fjC��JB��^�v'���M�=��L]�5�1����,�5�]��a�3��;N����}�#��8�C�����;8�q��?3��S�K��7��ˈp����S�s��6bf�2.�n2�5�<�'�r�7�2V �S��ٸuc9{~�3x�q�,hi����(̶���$�fb�F����1r�e�D���D��q�/�@����M�t��OkݕGi�uM�㬘*��^&�pb����VT������[����,����GG@V5�ǻ�x�&����nte����Z�R%�%lܲvp�/|v�d�z�E����5�0�ʜ�E��`�~v�����K�f�+cu�!�d���߽o��3�yek9>#9u�t�Uh���0�Ӷ0�i�-8�#�O����p�B��}�}��8(Úq!��n�2���_I��hǵPTt���Ux�����rK4NϪa��+]��k��Br�ttэ��V��ƊѠ,�+��5tg�ڟL�s
Q���n,�	��Q��b�f�����_�������]���9���ǝy�Wm���y���$�Y����V.���,�g��r,�o��N`])�(VA�.�&A]��.�p��l�v)
7D����O�Z����1;�90�	3rUtÉ;Qj�ʟ-79T&��Lr���Jc�����`Jl�P�[\�T���Vypn^b|�`r�8S}��S!��P�!���v��4dr����ћ�����O@�}˯�	~��,-�K���G!�Sb��(m���S��~*j��?V<;�5xYuJ\�9s���*�"L��ʋu�2��8��A[�J��sS*r��WE���P����U�����J����VgsM�,;��&�:\�Ns�7�W�}/}X��H���l�N�4������13�~?pt���v`��I�r2*���x�,����/-P�[�n`���"�}�1�;�w*��3\��J\���/4g�rhq�&n��A�	9��X��Ǉ\d�L9RUF�yQ�\j��xm��Ñ�'��.����myD��WDy\\���U2d���c'f	�.���b��8{p��rvv�'��?;�u����O�9}���YN�
��`�*��j����3A��T�����31-���\�Ɲ8!�1u�4
�Y"{��d��!�K�݃�;������E7�1�J�7�bꍫ�@�4�풫i�^���WH��NZ�}34��ۤj2'�T�[�=�k*.v`�.fe*c��9V������P��Ql��l��cWW7Z_�FjlEGZ�-�ZX�B�ɐTY�0��p�Nv��5�{��N��)��q�f�J��·�v2g�r�8w�Cm�]�7Q�P��\�9�f�b�u��|-�l�x� W�'y�}���J�7K{sSc�l` �b(޲��.�\�Y�(���K���x}�Oەײ�ׁ`�*��ǡ��2�vP�IJ�g��\5{y�F�b�RV�U��Ch�g%���Jlm�ju��lͭ�wQ[f_M��&�P�̷?<��>ͯ}��5��
�J�p��9��}�{�PǛӂo�p[&��X�޻N��>�<p?*=�y\m;��Gi���fb�X��{y�uBI�2CA>?m �:�ٓ�"����K��.*Va��ʬ�7{����F�(4�Q�Lq{ݘ\�j�Η}L�L�z�ވt��@�b���:����(]���1\X�����|PSPCh�a��u�q6������i��d����;T�`W_�n�{Åk/z�3�۬��T��A�*��"��S��g�����Wz�";�*���.]M����7x��BK���rZwcc���:���yq�JUS�0�&T�ѐ��t]�׼+Te���K7�u9��ڋ��iT>w�4�`�6����:�2Q����k[.���±)v�{�9	B����BZ��W���:�у.ʽ���r�8}S�F��F�a���r2�ƾ$�^�~���FP�Z./�k���N���S�������Eↆ���dۻ#X1����̊-���%Z�[27s���<�ܷ���]�Qg��&��Nfs%���M7����v�$�PqyE
>۴-ڷC���<ZY��w'�V�2|�o
�~���|8+��2��z2YD��iU�2��`D�	�0�#�QQ��=��5�4��.H_�VeU����*o|TIH��t��87\�`ӎ��Dfi�}JQn�޶�/i�)�n��(�+=e�}�M^�U�Ii.2�+��V���
�m�Kb���i��4q�/ĺ���M��gV��s�+4����|����^��A���t9�[�W���x���TFK�Eƌ40�
�f5:kAug7�uZ㐿2H5�v7a��[�D�����㛢<>��u;�Ɩoܼ���L�p:y��D)��^і%��oj+j{UW���~���є���L�"n'}z���������S��Vkn��Z����9�.'�`�Z,���yw-k�2����E�d%hCt��^��J�m<��A9�f���.}�!�љ�e�5#?Kk�^�"s�]jC(�Rō��*>U�ZJ[�Rq�]�c���ը%Y�J�uQ��y�ZU��ڍUi��h�����|�6��g�s��޼��cD����5FƠ�Q��G(���i�^�X���vGV�+�j��� �4����b��1��	,�*�n��Q�W����,�F��Dg�{����@�@3�F\EK�R��Y4d���7�y��1R��AR�D)�Ę:P9����#7��ed��L�[el�������4L��*%�'\�X�r��K�ת��V�8T���*��"�g
��vu){+"���-�Y,�l�:�f�L�9<��q��-��b����Эۤ+�$�HO�����}[��f�����d\�&����J#e]z��F�>�=����Sm����l{u�+�b1St�ݧ��Bn�c�gz�S7+qzow-�su��<���T��G���j�ʓ+��.���n<K��
��B�*t9{\�V�Yj͇=�5y�#�������a���޴����ĳ�{���Z0c�;���ý����!�žO���9(*��6[��计�.0q�^��u��,f��/YZ������/�1eq���Qs.�s��uh����� T��O�(���g^9pn���]����)�k�f������P��F�8���\�iv��u���)W���(�sN*�y:T��FA��e�����du�kG����8�e��Uڃ�F��A���+ׯ[�u��@t�,P#�,��`���DPP
��0@�J��ƶ��cq��"ʐP+1�(����`S��b(.X�c���h��h��+�
Jʋ�I�*�YY(��bf"�J9�B�VV6��[)Z0P�ZZ�5dF �AAq*
Jʖ�J�"�L�R[���*1���(�QT�QAf$���Q���@6A$�ϟ�|��[����2t´z����i����
�= mh�I!�Y7��r��衉,U5||�fv���9�;]�5e�(��
�V�7�����ޱ�ui���ʖ�u�3pD���Z ��D]:��#4:�)�a�`׬��c��,]�ʊ��5W)�Q�D�W����F*����z�B��|�n�K)r)u��[UbG/|c��Ɍ�y���S\T��F��O8��W�R%в�k��ZO4+�cA'���2��������rbt�5�{dm9�k=��ykV�b�Rmx]��|����@[}dez�O�×A`���Vl��ո�n��T8�]E�N�
�/rD�%$�pD��Im�q/^Cx���l�����+��&���Zp�<2�|/)�<Pz���`^�a�L���aj��Y���00}�N�9�|;���4�v�h� �&��W��d�˲��V�X���=yZCXQH�5nz�L��#M�I��:���%���T"�^�p�XG$YN Br�)̩�U쳲��C=p��f	P�R��n�O�9Q����>˚��/>;��C-_��Ҷ]��vVr�A]����at�}r�"���E.��F].�I{j�&�0�#$�'����@��@j�}����������'m�x����0��Sڍ�9��i,��iS7���ےaS%�NVwN7%��&���&n�I8[���L}Py�z%eM�� ��&ዎ3*^ͤ�����~�z��([�^
E$�7a:�5��]s��k�b��{*��>y�޴J���e��f@�n��͡\�GK���+���"�ٽ�S�Te�VѢ�\�R����<�B�O-��w<��  Ě�j�������llp��`���$��:+�Sz�)��Pn*7��V=+�mc.\����ϓu��[�}X4f��Ea����,.D��olߝ��v-�XhaJi���+�q�;㹒t>�aנ跻:u�}ޤjg��Z���b�ׁ������|W3��J��|���{զ2�c1��F�7%F�EM㑲OsJ�1CA���h8/�ċ`>I�����2�YJ���mmB&�Ta�"ޮ���K��7�/RL�F�EA8�
���=�D�V����7K/���A��i�BQ���P�Fez�o)©�
�\�Z�廾�8�^�L���F�y �
�헳�X|M�@��V�+=e�`׊�*V�"�|S��Ҙ;o�F3([J�kD�s&�:|�.�[~��lv㻸8��e����F:��}��� ��w0�{�{�,q���x�b&�a�Hj�I�d�6,؎M&��
�{v�1��v�c�&��7R.:M�3m%Q�rY���D��jH�)<�n��3�^��t�o0�+S��� I�(�W�U���`��|�6�� �c�ܦϦ"0�+���g����[ꖫ[mv�ެ
� �;'!�V�$�]�3�y����~{S��\Pԭ���N=L$�.�wj=��"�7V�v��aws��oMV���3M�tS	QS|����x6hI�l�u�S�ܢ���7}�������@� ������ٹ'�/��B�:	j�G��ёV2���P��=��v��d���U<�Eq�me�้/i7n��q�
K0��ĸ�<�J�Ԝ�z�;#�Gd���,�p��'Q��QX�.Ir�����p	�8�pc�롢+�J��(.9N�q���W[�:�A.�⋻=�x����e>���-9��
�u��`���	�}��1�p��f��C`�/:+C]�1��[�}U����u,^R��ږS}�o��V�����s�z/35&���o�U����|o =��F�ԗ�qZ����-zv��	���a{��Rty��ZD��N	.� %v��	l�4l���*���P�i؞]�u~�XӀ]����|��F�)+���Ks��>;�.��)QF�����۸<�l�mڑ�6�_%��Kq�R���F�x�$o@�Õ<����CB{׹J�~�'�wTJV����-e�]׻2v��}�Y��шŮ��G"TT.V����Y�K=�^�U�u6�3�h�l���ln?R��s6D�g���ю'�����`E4�]ØƮ����j��*�z��|Z헢���B&,]-]��L3"c^�^��p�&�X�rm
��æ8��K�GF��
�)7���/���hH���P浣M��o���W��r� (��BY���H��w��[�F����Ifw����.�R��DB�z�f�E�q��^��;�h�g�.��Xʒ�'��r�Ҧ�_.�et�GNk%��LV��F�
�p޾�h8�N�H�h� %���*ƣco�J0c[�����͗��S<�I�TT�ёj�]2{;�zC'����+��t��+K�z6�Ra����)K\ҳ�w�-�����k9Ȩ����ئ��$��i�{f�!��!=yn/S\˓
4�Ew��p��sw=ۡ�-F�Ʃ�y�]8-���%����^��p�o�x��{���Ƽ�d��^�d]է�4}̷V*x�F�����u3�z�P�7Z;y��oԔ�W8S�9�J:�S఼��\�W�k�9MD9a��x���u��q4T�����G��X+jΓF{ �P�̷�5��"�����F+n2���Z
�5�ol����^wEoi����ϛ\Ӵ��`������p��bS�A�6��lsnk��Rd`nr5n����-�����@D��n+�X�e0m���;��vS{����_@��]�O;zebH,�n�x��M6#φ=�\��[Y,��w²�j� ��tbhl�9��Z����]V����$q{�{��)�Y�9��Ai���Ui��;��z��XykA�)t���,��n@��71N}*��݇�n�];pRj�t!k{�
���	�N��NU�9M�� S~��x��7ohiDs^�>��x!��,���P���]�=u�x�z��o�R�r�r�H\Eɬ�5Z��I=b�nB�������(����H����5��ŃF$q�1�;�Ȯ�аj@�[7V�\�*�x�_z6�[��
8�������"���.:���3cގ�����C��)�b��h��Wly�ud�����s��N�N>�/-[�m����u��`�Q�%o_ÙY�ʮ����E����6E�:70p��
��p���M�Q)�	����k�<�<=�����{n��|��~o�P{�sx��hD�S�o�rR�ۆ�4�!�;o���aەh���p��/��]+8$�,�͊�U��Y�*���o�ĸ��������xu���OJ\�f6p�c7�J�^���͟N�+,�V"�]�'Fz�\����Yv�XS�q��W�KJ�F��+��׸�v�ѝ�y $
n��e�a7\���d
67q'�|2ø���9x�(1��;�����J��Ɓ��mf�eAE�},�󳉈���;�5(���i���g������iܾ�<r�Gpj�PZ�v*4�	�
$H�u��]�G*��;�@T�{�5&����;�ͯB��O�fi:����i.�%��+ή�pD�D��;bVZŒ���sg��o�^��Sv9Zհ���O�Lջ�C\�B��ܣ[ʭ)��%�N�\0mVM�3u��x_r�i·Ɍ�2�7��YO�����n�0	�X�GZyV��>U7t��5x�djP�"�h�ي�PB��K�$�{dp7�::l�_�(�@v'fYi���j�D�5���;�wO��g27h�X����\Eh#�V�* �磬m�}X3	���s�b�{�MM�!V�P���z�F�3�9bG�dB^j��Pv��]�j4�JYDݴ�j��>�ȯ"�Y+�%��z�O�f��� ����Û��7�E]6��c"�/1�W� yW|�x(��w�S�Ys7](&!�J`(�w�|u)[;:T��(I[;e	'���݃:Nc��g��څ;A*�_H����K�C$�\ܳv�r�|��t�
�@��cj��kW�20�`c&$�.3�T2��U2��fJ��
�b
"�)#h���S¤Ĭ�B��B���2��V1ea.Y��f[*0Y������a-�"$Ę�(�
(Ld+r���� ��m���02���Zێ]�TǦ*��3�C	�*.L#��C*/��s�Zؘ�5v���w�O�Z�H-�2[`�j�-�!�R�M�=�w�zA^���}��ܲ�Pib�\�����H"�I�{YQ'o�N�Ij���t��D"����m����[ݲ��^BE�SD�O�8�ԝ��z��s��D�歶ڋ�zY}Jo)SqP����p˻�oW�!	�̰��ZQOD�����r�HM+%[
�q�(��Vw*��&�1A�Lq�͚%���/fh�77"���	��s��p6]s�J:�F!qj�c�<
n:�)a̻�t�㚞��T6�v�<�J��3Lnm���J�o8o��d4a��w�
۾InzSԐ����Y&"�!��\R@�@�7NF�����d��;�[O�M7B�b�6.����gn��2]n����S��ش�D�������q�u����-s�\y���g:��];��/ݧY��)�@��;͝"¼�[!�۸�-�,)�`��z�n�_"q�3��Y����U�13+&���i���m#Ĥ��*��=x'<�o'�y����7DA�q���u�m�Fq��ȼ-,�\jqܕ �J�&����Z���^��E�Ȭ}�ܱ.O{*I[��LJ�gr�<s��':%��������^���kn�K��.�1+��F��2{o��mAJ�J��5;��k���N3�F�
�R���V�z0Eih��~�Q*���a�Ɠ}��:�/*;&�o��2�!�r�	�qֳ1�_rw��̫�{M;nT^�����w� ӷ��]���C4�
k{`��8�}l�$��.��Ћ����\WM_u�*C`k���`��J��xU$67:]ff��t�秶��	�I0쭫�oS��7٘w�BkRЃ���>�;���Z1�{5��b߈ #(�����޹Y6sYa�o��C���!x�ucOC�He]�5���]Nq�ա�:�P����;��Ľp�c��՞��������O�<:(�.I�&N3�3��Θ��Fp=Sܧd[�����>��Fa�$��Qm�X�z�����Y�;h"��=�޺U��w籖�U�J�˥�r��m��y��'WY��Z��\�ŻA�᧠��	���]o#����+M�n.�]�c;�"W�ۊ����t�n��h�M�e'�"����g��\�	��ʫ�G��;��=��&�.�%!% ��K�ʋ��%���aB�u�� �#���5>R&�&Z������}�"�����	��ה�p)�q�d��y��jX��U(��A^�Sn�i�%�?0)^	�e9q"�1�{U�S��v��Q刕�f���,�unZĵ=�	$��E,x���Z�o�LeI׀�������E���mm�5�^oX��çX��J�O2�Z���ve��N ������n�ůy��g-�����أ��	�,<j���;��d�h_�`xE�����~?F��7���c��}��ᬸ���	:��r�Z؛�Om�x.(�%���]�%�8�n�<����і�l���޽ �e�y�г%3�P�g���y�d�N�s�-tu�h)Z�T$��sI��uY���n��3�I��d�
5�L#0��?��K;���=y���ͯ:�2\�0��m�,�2�j��Ų\�
���&�>��,��l�Ƞ��	��/Y)ɰ��xp�Ë��)6��������U�8mk%7�w/+F�a�izaQ�7��K�zQ��-
ٚ�Mƈ�n���*rR�ɮ��\�u�#�-�ƭyƼ ��ރo������1J�dB�ν��9�UBƔ�;Ca�!p�Z�pXӘq�Ш�nL��K�Ls�U�����7�qsx�tPq@2x�U��}� �τ{0Q�=ᾸK΄�Ip����;�tȸ�Xa�M�SW��z���2���qZ����9:h�b.Į��!	�p~V�s"��w�d-ct�����Ko+nb�f��2䚳WV���4�i���� I��ʑ	 ��[w���,đ�.5e�,���܂�k2�A� +�P%�b���ׯ�m{�
 �Xoe�OW��+d&�I^(hl0����
[��Qy�j9����0(�^c�������w�M��n'y�q��ԿyPH0^�8j�u�;��j�*�t����pܧ�4V����z�a��#�Ⳁ2�(�	��1�nc:���̭�[�7)s�I�*
h�b�ƈ�Ög�,>&�8ǣ=�Q�* :�j��^S�Snkw���KX�lYB��'q�L����I��C_#3xP�m9��i�����f��
^d0� ��'��9,�!���n�i5�3�DB�� �)�O�����oV����牧cx�����bɾ�	t����RkU-S�c�zEZ��/E���~f@j�������S�� c���P-�#���p�#M�sC���y�9�~�Lm���k����_GsW���-�f�/7�"֭xFq�$3�(�w���[�`�
#���UG&s�~6���t�I<|x�<��+����ӌQ�Eb{���p��ZU
���W���	��T���t��4�#��U�~t��3������}YO�i�m�˭'�}��C`% <4p�I[����u嚝�՘����W�6�1u��T�!hY,���X�b��2�c�nƳ���kDJB�>*C�{�Z~��=���}ߦ����|��c	��9�zY��`$��YV�����Zw��:�[�008��f	069��n�]�y��:�v�챺���|��z)���FMSך�V\k޶��yXX�w�l(X���7Ǫp:�Ǌ[�U0T�}�Rx�OF� �;2�R���U�2�UgH�0�Ǔ��=�l��*�s�,-R5Y����=�}����� ���atoA��_�� �K)8�LA�����qۇ�|@X�ewc��V7]į^�2�k��D�k;������t'�Y����l�ǲ�MnI�,C��O;�+�S۔�M珠x��� ��%�����1�<��)*��[s��єA~���;��t&�pٽ�����7s�o�P�Ԟ���R�����0��#Y����^���C�Zm0�7���靖��\�w�UR��ۋ�j���jTR�6����)v�r��%ʊ�L�w^+�Aj�1��e4�/�������xވt��R����u�5�LD�@�v���z������r�p�<�..�ojA�fA�b�,�G��M�Si.|����䍇�X�g0�<Q��>��^�e���Ǹ���Qc7|���sv�k,A7����`3*Jx������.�e���H�(.��R��]�P�;aQ��.��s*6Y�ܷ�v
ه(˭É'��q҄�/n0(+�XtAvt��
�������*�u�8|y�e2���M��V�:n]K���$m�����v���!P"���̆6���7�^�����H��*�̕|{� ���@J;�}�vOB��X-4,�eյ��_U�K�����I�p�Pv��ɻ���=N�Y_�e�R��`T]g몢z��v!읠�)|G ����Xj'���s��F�J���*J��Z'8���(z�%����9Tg�+"E<�eI��n�C5ic�&��"�j<_��`�"=���sy�����<�����\��g��i��b�*^���J��R��|�)wk�y�Ì�.K�;�Y�}�y\� n܉�I[}�a�%����9p� ��
m�<�ٸY�~��o�v-]�������ڹ�.��{����.�SVn���%Ի@g����������`����۵�)��P:��¸{7�7cjܢ!|���x:d����-�����i�9�^xydx���y+� >b}��ğ�=u.�UK��ɕm���#�-8/Q�_t��(�MR{-I�`y������T��J�U�'$���C�ˎ� ed�uʯO>���)9��� o=T{C�����T8�)i��`���ob�7�!�R�ko�ȕ�It�Ryx,�R�<C�́���pd�7ǹH��)�]lL���)-͒���h��0��I7�4���]t�W���>1.�;��D45���ܸ_٥���;J�wf$̥f0Y*��d�d�����3fX�+�R+�̷���I1
ţ�P+��m�c ��2� T
�n�cY.X@�Rőcl��1+ �X
�
�A@�E�I���LB�h0@��B�+A`� �s.5Ĭ2�DP�V(�PĬ�`�#l3,*��Vж�d��E%d��,VҊ��" Ԫ�R��Kl
���W��u��<��}�����쭁\�vZ�m9�wT7���|�5�"�)�AƜiL����`��i�{�l"�s#�,�����e�\�[����Q��7���pAͶ�F�?]^d_
����cD�c��m%�zᧄ���k)�=@�ev>�J0�y��cxR:AJ�D��gOi�yk���}䛮��3v/��������s�����ć �J�(h�w���Sm'���B��lj7+��P�ٻt�pNַ��X!�T�UV��2�E֔��2r�8y���*��ܷ�o4������C����H�_rʽ���"����;�-ۥ\��������$c����]�O�����5�N���4p�}k��L&���9�0�$rKI���]�\�E�#��V�.��X�e�;!�����C��%j����\z�7���N8�>�PS^"���1��Է��%�e���ù�P/��P:oS}VO s�o���q�*t�oV��z���[�`�	v8Я�M�
�3�Xܮy�ʫ�Pd3�Yֽ�`� .!������Jw-53���X���1]�dQ�&.���ڴ%LrmTs����u�c=��}���i-���ޠ(A�����M�{��j>�0�=������f�-�ssJ���)t5��e���)}՘r�l��LGr]�r���l�G4tjnۮ2�+7܋4�����3�����k�����n�ܝ��wgJ��lܮ�ɭ�8��u8h_�U���w ��oB�%��(��[��騜\V���hn��`n'Y:Yț��-:����tz�;� C��`��9V�>�|��J�\�c��̃��'*S����R��0�����SO�޽)c��>���1*��pS>-J;%ak��k<1�m?a�}(����ߨ* ��c&���.{����~n���k�NU��H^�J���+�������L *<S:}��#/��W��\��/ׅy��{h<��XϮ�<�Ckz���P�#.�No��h=H��cǗI�Ț]G%�W�Rn���͊t��G���jM��3*�ⶓ�ݩ��ܕC�涺Yi�q�\es��p�\Wwd1fZ�g.�P&K	�r�n�%��ԘVV�ܻ=m̦mv���3Ϥ��[�C��~Z)�>�^K�īUړK���4R ֚{Y�6vs/;C,)�5�V��*�7�W���㌕}o�3�o�;�������;�扝ֻ�!���ȧ�.�=J����������=оvX=U}��D^�k�G%C���HI���S1U�eWF
�цc���>��)RF�_�����OG�x5,�[��M�;�U�ǉ;�p��٫��'��va)ȱ-�ҫa��P�ϔ�>M��eF�`.Hށ�g(	��gnh`3Ѣ7]��T��z9}�Qp�c`�]Ü"�f�sn�p�'�6yK"��7�"�iǈb+��Ɖ�͒���s&ƹ,`�9��n �]*��94a�!8��8�®Ջ���������P�F�4X#"�c,�P�Rr���		��ɻ� �\o���d����y�=��b��q6�F=��9��՜�������2}m,�)%$�*�{�������e�x%�<6�:h�+(us�
ri:�U
�g�/�
T��s#uzԼ�r����qx�]+B>��Z��>0h�v�W0.u�^��T��	��n\���֘�q��7�� �}�/��gD��d+�Q���`ʶZl�oܟiy�V�������w).m��{��V�.r���������3����6>�24LȾV͗�����ª��	e��I�&�c��n�U��2s_�������%��W�u�ʘ���B�#��qO�� *R���E1vE�F�Cp_�&����{������k���=�%n{�������Hi#=�Xk�����2Us���mm��cb�g`��?*k:�x�=Kj�:Y��ƞ��;|ы$|gV�$=�)�RgUΩ����ޝ��L췶�<xv�7��,h����6`�؊�u�q0㝓ĝ���!�S�O��[�2ʼ"Q/k'�jZ>�ZWMA�,�8��QMKs�e&dW+ݶ�9�і�h66@o�Vwm�-Iq.�=�Ro�ƨ���-�2�tK̷���Q���x���;o�=��R�:���<�M.��,:X�uQy�3�@;���,XWǁ��8b��iF��EVƃ;y�&����,���~t����ba����Y�ۄr�C��.Ox�{r*D���;��O6��:�Ug��E��*T�����kY>x�m��9�`lx|3�5�oԂކ֚+�t�W��*V�U��w���G0�v"b�DM�Ֆf�AІ��7���W�	g55B�sd��վl�y:�w3�ԭ��i��=c�[�q6����4N۽���La1���d;�G
�+8�UK^��Wm�X-���6ȱ�*ہ���4 �t��wh)�����^��*�=��7�er�1�Y�%�ipWZ�R}|����t9�V�	��=FT��̩��x�\,+ѓUk�)�$V�|���^5�=CR,C�i0i�>Q?�I;}� O�
��9q�l	�r+�2܊{q��~���V�xb�#�Y�#+3�:h��.P���_gl쀺��u���c�eY��k�"�G���G~�o��]�-��<�����	�M���-,�6D̐I]'�M����J��3ڌ�/&9K�ݍ ^�8E�V(��w	��M�$��'���'ݷ�wu�Q��E閻抸��q�E[��ꇉ\0$ݝ����nч���b��|�)����-����b��`{`��e[݊PjLq7Q��sE*��3�c������C1B݅AM�Y���z���"�rG�^��=��f���n����tW�zS�f[T��,��xw�f�D�'����y=���}�g������Sk�����
/Q���'�Xx��r��L՜sڔ	v9Gzi��u��Y#
��@��Nc�P*���q�,8���/L���s���h�i�%��W�X~4���0�Uas�H��z!�3Vc$�x��u��S"
s5��`Ư`�s�J[��.����E��y�k=J�^Y�@�,9�*��@�ꝫ�~[ JK:CD��|�e�^���Y�hv�请�Lz^��_��	���r�Um`�m�v�Avҭ���½:s��o����H�P�3"Lݕo�>�PomT���Lq�<�f(�!z�:�9 �ò�7aL��T��m��^���~���������R�UU\�@$���<�@
���e�U@���ȽϿx�u,�,���Ο�~��5ў�S֋'�ޓ�E �I ה0;BÀ�{.K�tȵ
������

��bR#8�+ο���}V������NO�s�Z۪E�L�	����;�߽�w���� H��}é�^�$U��VY��� H]y"*� ��U@����������{S�C�?��{����_�@��:w�z�$�� ��c��~�nP�@��"��Y����o�^�l���oHW�V��].��f��m�D1��^�l�'���$U@�k@WN��To¯|` ��T!C&+V(M��!f��p�*���Mh����^���&ǎ�q]O�'��"Ҏ�8v�&F��t+���Y<�u#�h4�eU@�Ì��u�)�����T�)>��h��%�>\zs9;�!�\����A�ӳ5�/����p6 Ta�c��M<�[8ЏD����� c�� ��/c����NȖWu�>�s�y��	�Y|�ꢪ��v��DDƁ�B 6|�GT` Ci�㩸Xk���=uZ�'�=�:�$���[��h�q���ʈ*����~J�N�U�g4>l)ޚת�{�Ov����27�ԛ������k,o��a�w����I��lJ|7fb�̸����+�X�G��g�v�*��P�&0(~�T��k�{\S1�j�C��B�6(A�yT�AD�n�=�>�����eo�o����q�+���� UP7�Muq�۴b��
�L`���5d�C��H!�6�i۴�TY���T����45��#�Q}��DUP7�ӂj .�w~���eq m�%�5�fA�pA��Z�Ys���"�(H��