BZh91AY&SYm����ߔpy����߰����  a~�q@ �    " �@��@ h�(�   �      �    yx (RD��B��(d o� H(P(�;tHWJ�gm�jֆw#��]Rɑ��nt�WXv�#@7�x�z�U,����x��Y�sX$�3bh����g�y˙EQݎ��a��قP�ѐ� +� 7�tH�V��Ή��bCZ�[��
v�����Tk]�r8wwE.̕m�-��.�$�R��� Q�5J�ɠ�
;g#J�i�0hvʦlU6�U���Uv2���ە��7`�ݪU�Pg:p5���O]w��   �4 ��6`��\t�WCF�䝵
��sJ�ã� ���m��
����&`�h6���� �I��
�n�v�Yɂ�䦴ڔ�t쎲S  ��jKs��ۗT�j����W0ɱ�f�x�                   4���  ��x�z�*�e10&#�4����S�BRU(�Q�� � �M#&M'��0# =dd0��H��R  ��` L�C ��BhCBd�dĞ� �4������iDF�*�F�&�dѦ F!� �a��{wH巺�euM�qӣ�r�GO�ӳ�籶l�:XtF(ӝQ�^�ó3l���^�7�7�?��e�8��]��f�n�~�����K����q�n�5���̳u�l٦tC��Vβ��+���[6͛�ټ�ܙ�*���l�wi�-��w��c�~�I�9�}?W���K�?�^��g�_�|Ye}�0�>� �g���H���)��ڑ�Ї�'Î#�E
b���L#l�0��f"Y�WY��ϱ���0�o�,���A��蝔�*!:%0�F[�T��0�B_�fA�������z�`��p1@�xI�:�H��q����}��$��p�j$�#s1'J0291zD$�L%?`�Ǆ��f<'��c�+1<���fc����	��Y�G�b?gfN8�BD|�>���'�0�1e����raD��<p�f>C�@�L';0�(����BX�5�	�"^3	Bvȇ��pL2�c�1 �C0��d�`���0���pO8�aD�P�ߦ9dB`�&,�.�<H�>A8#0�x��$����W0�"{��Ye[1�q���"H�L#��>�zxH�Jf\����~&G�E�a>�",�0��t�a���$o��9�x\����gNJJ3v�$�<$���>���'�~�� y	�j(Kp�0����'Ȗx�zF����v�f�G���xY�L(��f$���c�"<�0���rRS�Ʉ����<%�LtN	�D���Qe�qdȖ\�x�$�g��Ĝ!�LaoI�	�V��՛�s��|O�K=�)��zZ�x<��w:߉* ���@���"�b���D�f0XÙSpb0��&9�G�5�Y��UB&���H�8� GЈ���������D"<��LX���DX����0�'G#�����\�%��T��a=�D���$�c�B"q����"=�ǄFc�D}��1e�1��>$G��xc���:�Q)'
�� ��RJ$�Y��2�s��!=#����:�ȎdL�Y�����<P���0}H D�%�J#��	D���ĢYW ��O�(y	��9�"y�$��j�~A2�|�	�	^���j%,Dɀf'ǹ���%	Lħ9��:dǄ�r�%Ȕ��N����} ��K�'�J��a�"R��"p�X��B9pL'�L�pf���S��BA�Z�OM��8`��O�'��7�lx��~��(g"`�
��DJb!8"y�J"#}��(�Rc����L�(Jy��<�2"#|���(�W�@?u��E	ObS�%�J'a'�x��̧�cO��ۘ�Mc�8����y锡 n8qə8K蔑%b|p���N�ב)buȔN����D��D�O.e:��y�yɄf�0zD�1����bI�H��:>��7s�6̦��E���#��#p�8�ɟIdAјH�ys(����hL�Ie��KS3P����,Af���Љ3Lag=S3Q�)��O!$O9��ߡ0E�N	d]̾���� ~�x����{�4כ1������y����(<�k��kǟ/�_���J=\=nO'���3Ӧ���<�g�E��3%�:�Gn ��bS�	bx`��^����Q*؟=�X����"TB#P�|��GH�%��'!$��a<%>�N�ȎTO9P�aŏ&>��	f'�	�bQ;<?1 �G�$J)�(��8�R�ȉyQ(�o&S�:r"�	�N�1�	B�<��x��&��[pQ�D<Q^ȋ<p����bdDf��fR��=ɉ�y	K"%Lz�%G����ǼH+�	��<3ԯ���¨�ʬ���������,�C�ba�^ve0��ɗ�ӣȈ��?'811?!�N@ ��	�9�"H��x��DI�J"#��`����I ��D�	'�'N�P�J"`��ȝ(o����(�"8�tN��$�߸ �x�,d�QBTG�=�<"�ŘpL���	�U3[p��Y��)GD�<u����q&OH���f8#����̉��J{l��'|�����0�<�zHVy�]8���yz���+��>+�A������W�K��ħ�3<Y�	'�3_E^�ZG��ܓ�:�H0���$�x�}N<Y�; �Ⲽ7C��Ǒ�@ϦR�#�>��/݉�fg�a�d�r/�����C�G�>Q=�	���x}>��s4 �L3*e0Dr0�~�z��ӓ)W3-��/�d����ɔ��'���$}#�D����""�D�D��D�Ƀ0�����М=0��"~~����BsЖ�Bt�G	��J#p�1��D��@��c��~�Kj%:4��'F�0�Q=�Ģ9�p�˨���(�y�%��'9�<<$��I\��'��?7��6����?BtK-�Ja�'�G�9�<_""������'�!�+�NA?X�1#p�P��ɄG����b_!8=�F��8#�BDn�g�&=$|{��ψy~�B�?��I����&3���q�D��)�.�.~����D�bu���(X�ϰ����"?"G�I`����#,�2#�8P�ÐQG/����x�c�A��	^��b�Q��Ό�G�ҊJ&�=c� ��I�A^�j��E��(���������&'Ng�<w!0;gJ��x�Iߓ�\�	h��"P�1��,��&"��Bƣ伉:/&:S>�G��g�xo���0����؏�����dvb�� ��xDN71H	��Q,QG�tF:ON�tG�GD�1"#1�`�U��J$~}1q�87x�fcĔ%�2"'G	����i�M6�4�9l�I��bB�3@��z��t��:X�5d��\�'���Jx�(�I��T|�	Ѻ'�H��4P�y�UH��|=������D�#��N~%Xt ���p�(Q�'��ԃ�@����u������~�l��17.8�ʩ�x�$��G{\r��g܅s�Y6�O���V{v����}/5�Fo?�_�[�`���ֿ"���#9��g<O��n��nҎfr�p]����Ap�:9|Kn��x��$=O+G�J��3�����ݺ����-A|5�3����^b������<��?H�H�m�ofg�(L�3�����E�w���\�?O�/����dq
�tE[�[5�G��V�W���ՙ>^x��?�ׅ?��O�I��T���Ot�@�ݮ;�r��Y��?6b�T��L�y4�m#Vi�����s�~��3�i����{ב�9��ߛ�����aKsnH��c���w�:��:��M9��п,0�睄�5���+����+4��<Y�~U����J�Y^�tEt�8���y���F9��_�#���������'A����vs��6t�L�aY�g�w%j-8I9Z��v����m	�?��8�C��t��l�d-Д��|�ܛ�G�l�~��6��?-��D�����疼��;� �\��`�ȟ�X}����K��2���;7q�����$���g���zx��H|��z��� �/����;���n�������(���!U�>8���y6�8x��Pg�[��eny��Czq�y�y�V�<YXI�v�8N����Na̞X���o�	˯�/p�U�J�"w����Hg��^4K�n��·�%f�x�3^��p����o�.������}�q�����m��:��N=�2Hz��.4�ܕ�Q���?~��WF�_�O͒����O��g�=��I�,�75/X}��r]�)�;og��緄O�s�DD��I3�4f�����/<dnX1|@�?j9q��<���4�W����=��s��g7i��֋ћ��b�~��Q�������[�Xz��Ða�,揕%���\����W������0�����XD*������@�!,5��'¸�9rQ_��$i�g�4��>�r�b>�o���.�a��d#��~�ƫ��#�x���d��!H���޺n��?�7���|��>�fC��.�H߭��J:�,�� ���5����<�C��A��FO:�g�!rʦ��D�-<������W��[��	ξ�n�?O��>�	������.1���OK��s�=}�̩�sY���?�?�Lx�������|���A��m��8~߳�Y�s��uǏ�a�L6�q�g��6#���K����Ѧ$y����7���U��{�l�����|��O����O��.�K���Ø���Ons;�����=�'��T�
�׎�{�w�^xn���l�Ň��ڧ�ȷ�Cs�?�R�o�������D�_�ft�5���<{J'x�_ר@��U�
�V���~��r������{����W��������R��ˤ�p��/�NMh�u6����/{�L�����?O7���u��ó
zT�xԇN��n+4��Qi�gp�W)���V�=���5Ng��^}��Ufg6-�ǵ�s�����!��ok��vG����?s�ޞ���^����)���"{7'������L����g,���4x���'��?����{Z0�\�N��ȶ��t@<��#���O�N����k�qH���q����(����Sx�՚x��)7�}i���j���v2Aq�g���}~�u�i܂w??=��=}�1���p���?9��X�^/ gi�[��	�{8{̖ݰ�iL2<{	�E��;
/��快VS?�>�Z���~������JØ�߳K=�٧���^a�wU��̺p��2�����i��G����}�/ǻ�����f�i���?���N8�?��r��`�x�?�ۺ�����^+�)�1�[��3vU����׏��{ѝn������Gf^o<���?s��2U�o>|n�|=��C�����7����n}�@�?<9�y�YE��r�@��놓��͞�c*��Rs�'�o~�Fb���Ϸg<���gĖ��|������m���[�1����#q�g�ue�_8�P�����ȸ��ui��(�T,�}��P�RzQ�3���#��O7���+�2�{ԦW?��O:$��w:����W�^O�P�0�n7w������|����Y&��	/VHd���q���}�^��C,���Rai���e����2#}�����w����g���S{����ˆ8�{;YqD=�x��l>���~��aP�|�g�g�����{�y
��|��ĿfQ��.��)dڵ	�y!$(+�q�w�s�|Yӛ���ē9�E�N(�M��޷&���D����qk9ێ0�<pP�)�Wv���h���q��(j���]'��X�L���`��?S����x���㝧J��Ô'q�<KH���0�z�'�fC�ò�x��D������L���_��`V߆��>)\;:c�U��_ՏO4��aY�EM:��S�t����z���3B�[w?7������wN2x�<����x��i��ҡ%Wx�9�ֿ:��maRU�)�qX��־كr;��+�akc��=�i�T0���c���\j�d�˝�	�L�U�$�d�ԇ֣��L.��sT����y�{o'}WW��Ō��O�<4��~�)����b�{��g���ᦿ���)w�>?��?���g?~_j�i����1ֆ�3`���o�\;��� �~ل�/������xV�����>qz����g�<g�7�%�N~�>w?^0����h��Sĕ��aXi��
���/6����~=��N�ޤ;���p�Q�s���Xb�&e4�[��W��q��Y�����|8ۧ_2VK��]t6�8}]��|j'��K{�'�|cN,{[�޿�y߰׍�'ο;��7O�s}���:��)��!�i��\��뻷x~;�x�|��-���|��Q&�����^����n���6���A�n�=8�2j*�]�?Jie�rx��m�9؋��s�c?/Ƽ����Ĉ��ڤ�:�=#I�:4������z|y�O�3.	3qT����~#������<wB�H��Y�~�a�ӛ��7Z9�E �Ugy�hÛ��8{��w�hՅ�VW�	(�z7v���������>�윷���_k��GOo������͖����������ݷg���U��$�=�7����b�c?��,��)b-�ȟ���5��q�rir�,�m��i\j��4�]5��v�V�,%�duv�	u���#l#�[�XkvVCjk�ܒ���6�j�*Xhۻ+7wYn�-��[m7c��
��Yv��]M���M�}���l�v�פ����Hr٥+���ds���t�LQr'��l	$u��^�{����I"u�QҺ��]�v��ɬ�<өZ=��=m��:l;d�P��g�z�I�ϟ��P>{f
�$��6en�:n�MZ�Tj�`�6L���|O��b�c\Sxί�H�c��N��1Ϧ�cp��<O�����%ٿ5��gq=��fvI�x�w�Yd-��n���j��4[Y�t,��4�]?<^_wC��p�a㼷<N��>�\�0����Ry�$ڛ&챺�iƜY5_|�L���2����gv��k7m$�<9kq��H�Y�y'D�9۴�%$2a��ԭ��	g�ª��#&#e�H`++,�ԫ�٩��E����	���ɡA����0) �l`DLe6�*��%���jh�~�Q�r�e�~�i�Ge�q�M��wM�&�R$D����^�X��"� �H�����"EE�d�v��Z� ��$�Ы���"���9�$�VTf���ǈ;k%sO&k��XrCY��=c�SƸ7��R������P �Ql��B�e�+U,��b�%��ܖJ�	��hB!%��dxB��+��a�֐�����I�~"A?}eo1�9k��ԡ�҅��s�BP�_C��ç�C�b�V{a\����\�$�k\��(`W�
�{+߱�}��RD����E� 4���)$?J$�#)n	H��n��x?%�+���m�^]r��x��:'~���#m���ɗ1a�t䠲aaFl��Ɠv����4&�wK*;;'9})Մ9�'������
@�5��LAD�/!H���?jDE�=�$ӒқKf��25�ܕS%6�6�HBm��ݙ�I+u���٤c]��H���sj�V��{�T_���w�u{2d|�_ >�3�����d2����D�|�����������ܓ2E0׎Ρ������C�jgω�x�C�g^�k�AjG>CS"Oa�gG=uα�}�N��H3���
G�~�����\bϼ���σ�|��N�|}���l<}�o]Og���=l����✷������~���}������>?��?��_��/]�/�	UW�Ҫ�W��i�yU򲪭�ҭ����^�Ҫ�YUV�UV�[Y^��V�Wʴ��VUU�W����x�I��$��$�ؓhG�D}����D���UUq�U[YUW�Ҫ�W���^*+ջ��y|�*�Ux��U겪����V�W��Ui�<��W�ʪ��|}��DA����|��z���k
�����0��k*�����we�ݪ���k*��ZUx��aUUaUU�UmeU_+J���פD� Ƙ166&�h�www��W���ZU_+*��ª�"��������ݪ�ª�"���*�Ux�J��UUTUUTUUq�U[Yh�>�"t��tm�{==���l٢։%g��_������<^��{����ϋ����3�(I A��P�pJ,�`�&&	����,Kĳ�K<t�O"'DD��$�D"@�B"t�0N	gO@�$� �p88A:@�$�t�$D�(DL�Q"$�g�:"I�0�D�0�O&	�D�,N!bp��D�$���	d�0��<@�$$I9$@��H�8"pN��� ���O<xԔd���B�_����	}���vA3�xJMa��H�^���g%��ݺK$��H]����4��vݺ�H�6��,lN"�l��lH#�K�_�(��].�-�I�k�E6���۩k+�WmRݭ��]��͒+ll�qvRV:ld��Qyt�!���n��c	63Ql��7k���֬K4�Y$���Q�:k���M.�6�]�-�iJ�ٻY4�fUtWa6�7nݩ�Ą�dѦ����[�Mݵ�KX:��i7]��g1��6K0x1���y4E����7mٺYm���Fj�i,�B��v��Ehͤ���.�,]�e��M4�Ͷ�]��I�ɬ6����(�"H˩$�eo�Ӎ��Wh�Se�k6�HG,�6kv�[#-��eFGl�Vm�2�"l����d�B#�$�E�Rʥa��)�n�Ci�Ij#�FQ���0�7f�����w��4�kY-f��$�R��R�TY?m�Åݗwv�Q�.�k.��ٲ\���b����n��/7���d�Sd�Ҏ�.�B��-ذh�l�f�6�_��"�o-u7vf��ݷ���H��S%U�!'�G�(�x�iB*� ����S[�-R)�v��I�m�H��x�9�M�Mde�M�d���vj5�)awr�n�7X��$�vɪ{�iMr4��	\P��B�d�E��+��X����gLK�tX�X����ۑf�]�5�k$�M���k�[�Y�݆�(���6��1�v���J�$7�
�1�A"�C�R�6$2C��T�٭��ԒO�^gYW�0��M�+KsF2~y����l�t��D�l�f����v�+d�v�f�ˤ�,6՛
�7K���]
��k�]K��9[i�$ݻ��Ye7m�6MFAwev�l�ݦ�][r�wvVMZ��t������N	�m9!q����7P!���� m�C"I"�3
l)$&"�[i��X��D�KI|Q0�* ٺM�i٨�l��I�uuȉ�껦�)Z��建.�]Wm�B$É��l��-�ƭJ�6ee����fܺ�ғl�6��.�66�w"@vX��W���8�V6��]�m�I�MZ�ģ�c�����r��B�fIh���D�$��Je�[��])��9m�6d��M��K1�Te�#��eU]���= ;^�罙����� �www{������HI�����ffg��P �����ffg��D�H��x��4L4L,�(J0ç��O��7�I���ܸ�e[I��В	��r&Pd$��jU#k�9��in���-��l�m�PE�n�Y!q�\����n���,��(��H͚j;�b��.-V���ED��$S�Ӓ�a&��5i:>)�Sf�Ă3�H�����]rcwYX[%�Rȭ��YM�6A���Ey��7��e�ɦ���4�I7vV��u�c���a�p�Z ����*{�e*�?g�e����g��5�ٌmwX�v�Hh��k9�4]�ܒ�����VA#
G�H��d�[cg,�{�z|p�Ⱦ�'EQ�/�0=�Ha�&C�x�!�g�Q�馈�h(<�JQ�?(��:Yh/����n�-��4G19��&gR�Xӄ0��U�N���:i�M0�KΉB%	Ft�<!��!�e�j�mup>!��>�1���g ����~8%H��J8R �a�m���o��/�	�.#�壾K���f@y/>�H��m�	Y�w���s��ÂRr}ɇM !d��#�h��'�Դ���IGK,�ĳ�P�BQ�0Oxޔ�����L�+��$i� Up������B�|({�m��}'�")K�1�\;�}�g�Ke��!���Q��^�i���)�,nxq�ъ���уg9��m����:\<pp�<?���'�6���ѷ���XxӦ8x�%��J�0�xC����N2��&�ɻ�gC���0�D#�p�~��Y�rɑ��Ů�'1�1����(�]D�����}R�P89�)�ĉ��L<a��b9�J(��E�w��#��ITR�0��o����q�
��p�����}APa�$ç�0�,K8%�%a����d�(���x��]PD%}�~0��)�,?W��N���mۺ.���vX���l��FS[��ac���ܷy�W#�<c���
�������6F�k�w�z%���Jǅ��z��ݞ�d�9zY=� n��/������88x���D�j,a��أ��8j)I�."Q�.K��%�m�)��uj8ݸ�E�$4��
�9������wq��;�*�g�3�3�y{>m�P�>�(�8T��xY�i*�9B�t�I��}�U�3(���x�`�bYBP�BQ�0Ox����xD�L�L�+�g	�J���޷ �\�鍠����Q�jH,�9y%��=Yphz	��[��xLL�
/�~),I����OmŘ�0�蛇`�����<.�%M+(�J]��i��4�;9sB�l��?x�c (�k�Ρ���ߨ�e��LĲ����:`��QEO�LFz��EH�E#�$��D��b��
�10����R���!��H��y{_ɞ���w��*�nݶCE���m����Ԓe���>�}�:�h��t�aXh�n�:Q�x��Q��Ac	)�?d`�`��R���'i�t��xz�D��?,0�Oi��%�%�%a����N��$�����`R��G�R�u&8cQ��tԄGW l��1��͌&���\�)��9�ǓN�"C�Q%��ِ��.7���G2������5�����ul:O��z,3v���� � M󥃁�Y������!��� Fo�~(��x��,�(D�(�
8x`��&�Ep����6�O�(�I7�B���Gk��l֜0���Tw�[�BMeR�K̲��"�!Vf4 ξ,�cy�%�Q�9��bu�k0��o���N4ؾC�+�Hh�C9-2�t,L�!\��&�Y�|��*; �U+�X��ߪµ������CD�'H$�Qg�$O;�������(�!�cr�Vr�!�U�{f�ldM���t��;��<<7
�O��A�Ɩ`���K$J(J0������^Y6V����t��Ft�nm��h�5HAg�5n�S�llk�Y>�DQ�N#������I�-R*1����4
2<E��D��x�ێ��y�-!Ј�R$�q���z1�n�2
NtC?w	���{$���DB��@�:29N���0E�8���](�E_0��$~�Ԝ#��FGC~*<i�o��Ge�/I&��6�UM�'���I�������$���BF�����N�N�N��t�:iǅ��ziQ�ޏM#N��M&�����h�I4�4���l�#ON���B:hF�2~��X?��)�p
<Fǩ�0�$�$��ŒF���zY=6N�M"�$���������>f��?��zt��:O�#J#G�H�����H�|=�ӄ|=��7�>0�:QD��zp����&��,�4�4Ӳ��0�=�x=o�^�oG�X�zI�Hǣc���(�x;4�,�8i=0�hL)4M9f�iS���18NW�������X=�n���/^]i�q5�s��X�>޹IG4V�.�q�i��{1����IW�"��s���QƌǤB|�a@�B��C涬�G�Q�lW�P+����n0��万�ws*�������YQ����8�̤�hy�x�t��y$9c�?s��a�/#P�iu��v��ﻆm���m�؞�h9���s������߿�7wy��������wwwy�m}����www{������ww{���4�L4�M�4�M(�J4ӂ'��ƅ�t�URI�x��<�y�ܝ����w�uX�XywRv����8i���Ԏ��X��a-1�ߟj)���>�#���F,��,�%���P�y狛�$3���,�c�G��B}P��|I-�H�_~:��T�)v�����Ӡlܣe��A�!M!�4���@-�"z~h�	�_�p� \p�����H�.����&��s;�]���mҤ��� �h�n՘k��R�L%i���@�cA�@�Uw
a2f2����p#�7>��E���X��!��6���	�h�&��G�%0��8x��M �I(ҏ8tӆ���Zm� �ڈ&�G3.��;�-Ӯa�Þ{�瓥��cl�:�gI���sM�������l��6���L�DN�=e�JRWl5��͇m����a�����d�S�'|�z���n�i�11qD$�`{�L=E�pb��n�SSApC886
b}��!E)�2�ǚǂKlpL��: o��뀦{���\�T��xd��F(�c4 T��wq��:�s���k[jg����m�(��d�i4�> _�4�����7-=V���O:_���&�1��� ���s��6��Lr��g�U�L\�"&s噚�9��31�7�e"y5H�4����N|4�4��(�㇍8hT_3�~��LӨ�Br��`��r���11�b��R�&�;\9��ՊR��*�N�"�4D\�:�y���8\%�� ��D	%��$(�XD)i�4�I���3%$�$?튷�����4�j#�i�+7+�z��|:�>Ǟ=ޞ��]��D01�"l��GP��qO��h�8/�V3`�%4��B�8:�bIq͸�u�9���c�e�-��Ɩv���D$�h������y��H�B5PBR0Ϧ�~��0h�$�͈\H"8bL��Ë��Ɉ�a���>Ä:r`Q�""c��Kh�H��n�\v�y�|x������0c<�(i2Q��
HB�P1�P*\%"F��ll�$x�QT�P�bB���;�4�n��gm3��l�����
\���@�D�ǿC��k�
60�M1	�L
�\"h�w�厙nO-9mE�D���S�:8H^�ԌC�!�P���	�
Ɂ��J�,���x�񇎟�b4�M4���<&�4"'��ӕ��R�r�UDD@��ɘ��H��p�0&i
� \&B�
Q3\!r����I]����hi>;���0q#�I�q��S��a57��sq��ɇÁS�8��	�ӿ�Y%�%l81�$�$iS4 Ұ��!�fA}�2��X�BMl�����Y��s�Z���B�p�Xx����@��=ɇ?n8�kB`�D����Q�DO���[��Y�w���w�����[�LMEm�D��{�3S1J!=f8�pp�gOʔ."&���a3(���tn�4�81Cҁ����(E&��zV��B%2��<ʞ���pDLp�209�d�(i�8��a���p���$d3�L��	4�ƚ|t�g��M �I(ҏ8xӆ��q�T����7O<������oUDDL������3�P1Q
H�y�`��
���9��S89�<�qa���:@��a������L̢S��u[I&�-�MͳLv�wuu�M�Nkg2qm�t���p���R1�� 40=!��P�p����s�D�r`&�0ID�����K�[�.���>�!�������y>���9�BX����hiCF1��4����B�A��88
iP��ޒv��Q;9�4�o>�ۮO-,E4���wG	Rq�M��*�
���%���Xз�I9�<�4+L<NRē���x�����s�:c�'E�5+o���u�[q$=Y���5A&����&D�a%Ō�pcb�@BG���:~���a���i&�Q�N�K47[ǲ]H��e�t��#e����y������g�10	�dDM�N�r�K;d��)�[���oNf�p�C�w�����P��Шh[�-��gr��ɑ4R�G(����,-�-w> ����؝r�rP�s���s���8M����ZuM���ۙ	h� $��P�������H����c��a�4��0!���v�W���Oq�Q9�HM�a	.M1��
9�� GBgUg��G#�����pK�pp�`��r��4pB!���\�ʷ�?��L� �z�D�LHg��0�Rb~ÐJ�#���>Zć�a�/�
\�pOM~>yM= �R�Q$1�8:��0�F�|x��<	��i�t���4�N��7��#�*���BH�J,k�)���\C7KL�H;���!nH�W�0E�57�YH�;��j�~�Y�N,���65�lvjWeƝ�UPK�����r}�ç�8~�	*!�a^+8��}zf^�`���0��qSΓ�p�VܞG��jB �0���+Àaj��ԆjA>�(��$?�L>�����l7�)B�fh�.��T(�)Lx�$���Ey�ϲ�Æw�FQ= �����08 8R��A�O�}�tS8&zPr�Q!C�p��M)��� |@IB�u^�KS �}I��tb�f��= "H)� �txQE�)'��&�rx���"��O���d݌�i'����8���EU 5a�x!�D���HD��y��I:~����:'��?x�~4�M(ӧO	�G���&�EHt B����$��&8tH{(�añaDI�3�%=�C�;��[�8�d��A!�C?_�H�!Ǖc�՘x�FI�{��ç�ȐN!�nA\ $���AQ���.�>!D1#�@�0�C<t�� az<e4!Ґ��!{���i��_�����!�&-yi"c*�ћ�I�6�۵����q?���j`��ypj���47��a�1JCp�>4��N��#�_ˡq��	a�XsҐB�ߥ4	� !��I�O���~�m���X��0f��I)6�x���a���<tA4�M4�N�<&�o�<Ѳ��g/.�N_��N*�&	鱑Y�~�����'؄OA�
&�ى�ߩ�h���e�)Ha�|8i�$L�x��P��>*LZyCch�e�<�Y�(a���DD9�đR;��m�ͣ+���_�M��6p �t�TJ�Bt�QH	ܽC$�g���uZaF���a��?�aaD�`�)	�C�l�7�e)F�T�HkI�p/�g!��4�8Id��?I�SI
x@�D���֖ӧ�y��<�|R���sO<��w�H�x�M,D��: ��$�J4��8x�.���,k��� �6�i��1��a�|�66��&p�� |�B8a�ӧ�J&� D\��N�̅���
��@�~��[:ݫ��l&��k6�3�܄w�ދ��R|B�I�S�zL��p�`�D��9�0�"i��d��1Rd2A�R\��(�b�(� :o�Eѝey����*�H��=QӐ��w=6��n�ݝ�a^MR:2Ob�L��2ID$��T|1Gy���jL�ގ���PY�	:> ��z8>#���~,��4��"�#I"��4� �ӄ�i�R4�|i:a:I)�	)BF�aF�NJF�N�N�Nt�N���� ziiiii=�:L�J!�l�M���N�F�G���N���Ѝi�R~)(R~��������ǣc����&M#H"�#G&����zl�#K#M�����zH>>�D|;>._������tz?Ǎ+J'HM'ԉ0�L(�Sf2c���E�H����Q$���$��LG����tviaa���a�����f(ӣ���(����> ��l��p|Y<g�i�I�t�I�i�eᇍ.�#O�=�u;�C㰟ٱϟ�y�՚�W�����=7�`\W�
m�#V�TQۦ�`�2�MEaC��b�����w��w�Vd}�Qy���1S���n��F�V�t��!{��x�+Yq���7��{�K-y�7S�����"�C��<�h�֑ �1�y��KS���85S�k��U�6�̣s�V���t�>�CX�7#9��O���ƋF���F��!T�t�QZ���fA�d'�;��qP�~�]Ώ���A˽8{��g��WJO���M�|pp�H��`ʴ��^�D�ޑV%WO˒4�ṕ&)��	��$Z����r0Ti(	d�� �,([I����P���{Н���oLh�����F0�#Jd^۰��$6�c� �dyT��]��J}wu�wK����KDT��- �7��r����_]����{?i�qTӆ&����!|�Ck,v�`i]ܟk^�z�ѿ���\^�㙙w�
���ffe������j�������oI$O	b"'��&�I��iӂ'���+�c�m�rŻ+6�Y6���EY]MԎ�j;u,I!X�JI4�n��cH�t#v�l���53+���vl4���Y&݄f˹�]�;7h�k5�K͊nIRE�]�ٻ��FI[%�-�b2��&A6�Z96�.�� �XI�l(��#$H��ݻ��H�u7�K��.투���JTS]Օdi����Ů�M��\��l6f���]l[����ث5D&$��c�]����4���Kv�Q�����<c��7�sٶ`�M��JGd�ڶT䈎�"�S����!I�ƴ�)e"h�)��F"��SvJ����ix��tJ���J "���8��=8P|�t_L�����yƜP� ,����rƸP|�D���� <FT��!����L�p?�T�}�'�}$J8�	!�G�����
~|SC]��%AH����O)JT�8Y&8x�������$�J4���if��g�(�gj$������6�i�>Jw����;�Z��3H�U�S���y�<ÇO��d�����$0v2
��w�x�i�.�](R����q|��U� ���kw�uI<4�F��Ǣ�vMI$�lݗ�{մ{�y�.��s=��锤 �d��!�Y�}D�ɍ�#���S6����D���1aG&�K��d��@ $�i�9�4pB] ���f��OOƒi�t���4����s�λ���L� �O��\�m��3�(Q�G���#�,�0h�:8T�p�(脙AG�u����� k�8J��¬iw�,�
h�����$�A���ϰ{��M��x���8����O�</�(^��H�<�<ծ����J�k�8�!p-��8�+㦢ui�w��+��tx��/CN�2"�aVY���Q�7'��(N�<Y�>?	�	��M4�J:"xM,��^Lxy�\,�L��uUq�?��j��1��(�q!y}�fE�xk'ԏ}��y�U0��J��5T�(`Q��8O��!.Q*��8!�. �@�Ԓ��䳰Ak2�鈝�����4a��BTr���J�VM�!d+9Y��h��Bd"S��~,��C%��R#G�_5��°��:E"������wX3	8WF�B���,��|�qEt�a0�n��D�jn�.�
P���x���~�D4�M8iGDO	��������a�[��Sdy7����XH�3fT�b�:�faû_�&��b���tL��[Hb�Zs�����|ƌ�5�Ye+&�$��yb<��˝����!���}�/���"ui���[R�.��zq��0�X{��j�6���e�j6`�9�c���/;�h&0�$�����o�q�&@à������JRt����<S$",&��+�Y)��e����zm�0��n�(s�EG�U�pj
�[֣^D�Wã
J�1#���t�J
%B�;�³���(�B�������~^^Px;RO�/�Ilm�Ѧ������|�>(�x�GPh��<Ȅ�e�?uҙnQ=M� �N||x����'�M4�<&�iU��r(��v���*�������>�O���h�W�D�� �G`pIJ�
56�h�������OK	$�h��1E�����0G��Y�
���28]sE���������|y����x��ts26A$�ll�餰�3�M83ǋvY����|�L-i�O"
 >:II�p�������GRh�>4�K(������D�M4�<&�ie�_O���sr�UTC�����0�����B1`|��&:G����� �-�ڢ��IHw���bӦ�+�Qd��a�����Ζ>?�"�حD}���v�M��Դ��-�V[��>��4�y�Zب��9O�]��f&ר�0�M���,�r��a?8�8�:H�z菭�DA�I��y�yt�D	!���C8"����p�I�8�>�60b">���(�,�O�x�$i�IG�<i���
a��3��4�I��x3t�N�8��!��O��՝�
��Aa=�D���$)}�;�֬�7YFXmݻ���uj�I�UT�#+��M��a�ǅm%w�F*�����T�����]�4�x�d|u3{�q44G�,�6"��i�>!�r�����D?�E�|\�n	�K0�s��A��I����$�x��Ɵ8tA4ӆ�pD�Y���O����	&�A��**����9�h/2:PQV�Rj�Lh��L��B�v¹�Sl��ݒF�a!V*�!�tzy��E٤� �1�$!�P�V
L��Q�5`�&Q2����R$�O!�yk�A�,:+�����Z_P�[��l�u2���A�mA,��J�d��|R�ӥV�cD�r6B��A<UrߏQ�9��4PPk|s�����c}D0:a�Ĵ��iDE.Q'ȴ�:]1��{���m:���ْI;�#�T��m����*�|}�Nړ�IH5��J+�ﾈ��ƣ�QgO<||x�f$i�(���4�F*6��ɔ��j�+�<Xͦ~��H���Ic�k�aE�y�#8��4}�:?#���1�`yB��W�2�5 ���Q� �cF�1E#H*L,��B��n�Lp|��j��D����E%y�_�nnm�Ց3E��wUw,�g["�h���g�~�8�j8`P�*p�t`բ<΍j6N�x����N�I��òQ�G����4}��'%��dQ���ಉ$��4�iA6�d���I��3N���a��HI��4��IM%4�(�,�,�4�Id3a��4�zF�zN�M#N���&�MF��GHҍ'��/H�M'M ���e���4�I���3a�$,�d2���f����pޑ�В4�4z=6'Fi�Y�i$i$@������Q�����_#��>,�:=<E�z^�[��ai&N�0Ү#BtI0�<>�G�H�d<#���i��4�f��/%�H��{��I��:F������Bc����O��a�Y��<>#���i�ON�t�24�=����ɇ�YS'9.i���A^a7|�ט��4�Y�	e�:�I�e9��1v�+���ƺM�,�1,Od-�!��H�}I��q�}�ɴ��@3��TE�0�����w�d
����� ōrm\KZNY���Q;w���9C"H���#���G���ٯ��a��9{���t�d��4�ޛ��M�����w����~���\���.��n���s��?�v���s333
���fff�ª���������^�ffn�x��,�4�<t�D�M4ᤔx��Ƙi���8uM��G�1E"c�|����4���4y'v�I��16Q�Ah��xp����GH~�t%M$����J��8_$��Ƀ��C<�]\EJ-Ap���xx@��}�ik��a�q�ݢ�/����B0�uQE�a�y�ts6���H�h�"[c�^�ܶ�#��g����4��4�$��=��Â~0���0 �M(�J4��Ƙi��k&F�"�� �R���tꪨ�0�~_I�>W9��d*��G��(�)��>�-�:�f�0�Be�(7Є~�#e�9���D���qw�K��I���Z,^��#��0�:BS�������:�_��M��W����PZ��Hpj(��8p�ȳO�Z@�)�?E#��Y��"!�3�"�}ņ(��~0��LH4�NQ�D🆏���j?���f%f�T������C����k��T��x�j�	$O���Yn��d.Ȏk����7f�2��7S]��$�H f��9UE!�b�-ob��
�?m��2�T=�߯�m���x���n �Wv��k�����Ƿ��`����C��<i� ��$��!�D��$�D�$4��D2��EE���g����St�D�.z�8Qg�٘��Yѐ�O"���>�$���t5�<w�8�gJm���e��A!�1����Ӈ�<:���I߽i�
,#II�ݩ���S�$�GO|q}����Y҂�AE#�dIH��Ɲ��ĖY���x选�i�J8h�K4����$�}��~��4l�A|����S���89��xpӁq�����b�'8�KS2�����Mё�NB�0hM�C�����&rb����M|HP@���9�4!�%#�R�\���)$�W���.��b>]�Ӥ,(�A���<��a���s�b�+�^o��枂g�&�)�?h��@���kg��	�ޣ���4������0O0 �M8iF��if��Ɣ��D_�d��g���t�M��������?�Hr�;��JҗԺYA��YF�oܫ��������%5����%����6��h�fđн[ZB�S���ǧ�
}qV�ĸT�	���8
���|�.!���K(�!���O��&	A��:S���F�,$<��ϋ,Ɯ���.�:Rӄ8Y��0��LHM8i�N������<�B���gĄ&$�?*�0�b ��A�눂�X�"����T���~�:IH�H�sY�>�q:�����u���	<W��⡍�T����㈢��G�/���	0�|�:��(iZMK�(�ؗ16��i�=+E���[t�9�f�НXwŵ?�>a���9��!q=��҆�pnQ<��|6Hۯs��Б3�B,�GW�a��O�>>:i��H�8i�<&�iVO'��ilA?�(~6� �D#$ˆSb�����e��5�ReH_an�!I��x�ʐqR�)�P
��1�ĒI�~AD���U�q�'��TD?!A��6=d�:�)=��gG�K��C,��E�Xo����曔p�N��Y��{����!�a��l�V��C�7�Wܸp�MQJy��m!p��F12B82���v�p�������Dp8�?xtN"�D�ӤHb:�E��E#ĺ�%����A!�i2QLk�g��H!ahg��%?�I���ط5F��u�,t���k��q�e��p�a�( �D�|�>p�K�M0���x�?:`"@��8i�N��4���y�"N�#m0�eT�s�S8Ӝo	n�着�y�N����$h��~{s2�Q��Ř�U�@��M6x�+&��gKK�((Pt�*��%[-0���2~mv=�m�ň�8a$( �ߏN��:B��I���c��԰�ȭ>(���=�?�i���S%��;�'
%Q�(�\�cXG�6R�Y�>:tL4���NpӢxM,��|?Xn���ʃ��C�Fw���G����!���k̓�,h�(�y9$0�,�Tq��,f"!�|daP���4t���:���?lԛ�M4��Wa6⋃��&F"ƈ;�c��X��8��y�a�����$�H(h���@ۏ������q�<
�O=�h�'�����C��Ʌ��?Yi'4��OÅ���ҍ(��4�NnNF8��x�*j��׷�.��=UTA�O|=1���@��o)������A�I���¥du�� �Bd� ���]C�7㥒��i	��g�"%�:a���A	�m����>��#(��|C)D>Q-*���G������D��B�E�X�!�}�GٝS2�yBg�EHjP4Lcƪ\�v�Y�I�|��So�|Yt�,dYDI�1�=4� ��J"6]�N�#I4��O-��M�i	���aZ$�3N��N�F�4�����iG��N�M,�4��F�J$�mF=,f����F���N�I4�4�;M%�F�I���ч�'�'�pQ���f@��f������g�#I"=4�#G�����i��3a�!�F�G�_LE���|G�>���4�I�0��t4�Ӱ�M#�������cBtIȍ&̘�*4j�&��$���h��4vi���=4�H#G���=4� �l4�z3I"G#�H� �a�4�m��YF��I�a�+G���~����t��Y>��U�o�\�k��[Cs��0��u�Qץ���*��e�v
|����\��e�z#�֤�}���Y����p<�9!�UfE��	��^�,etTF��͍j��G����}0q�j�ǚ1ׂ�)�⡖t{>dq����2�!-�C�}ݎU�b��q�1���tM��GlTg�_v��0�͙Z��\X�Y~�Dt6T2u�^�惭��`��;��< ����'�0��;��9�dcg����1S�/�SX��s��)D|�]�����?`-ÍI5�[�Z�Mu��L��)��8/q0�VlN&��ʡISz��f�)[���5�h��|$8���TnB�e��CsK�M�e.��*���q)3�m�FTH����Z�ךf�Uf;6�;uݥ���(���3{xse�E��K-F�"�[�6�H��6�,R4�aKR���7�W���%Z�e��_R�����jm'Ժ�R�Jsf��8�e�v��$�򠯼LL���A���������weUs7333wvUW3s337weUs/s33w��i�K0O0 M4��O�Ǉ㶧��� �),��+�I.�$6m�6�MM�5w[���/%���𐤷v��M�`�b��l&��6髆���������n �Y�D!�-֬z��vH�yl��]��lX:�'��U�9hT�a�~U�c(�(�4I˨�͆�mֳVBnͿ�8r�U��jD��,�XZ2�e�~M�!�;CE£,B����]ԲJ���Ld�X�v�lC3�c�H`H1b�L�j1�1���Cyl���Љ7Kl�,�B�tS��C�[m�0�y���^޾e?Ik��C��KQ�|���oCg�}�������4��G
ǽ~d?�(C<R!F�(P�X������o���A�K�I#��1�p|0��=�ӻ�O�O��-�R��D�:�8�a�P4|{��a��������Ym"}?���E�]�Y(�HPb��!�O�5nݫ_O���x<� �e�}�w�[q�:X`�($�Ř|x��:<3ƚQ����G��d6�B��E�aIZ�ߪ�>��!�8>�����u'A�;��U5����c )B+���Pp߯2Y�tb<0�I�N����2F�t�i�:4?j���z������d��X@n�� ��B�R,��5�����s�=9�0d�B����}QoX3Q%�J�	$�0e��_��MUU��xC���x�H�t�Q���t��gC�@�������3���" �k�ϕUs��>�秹Ӹ7#���;�⒏2C����� ��d$$��-��E��pcFA�(�RX`���<�SL�2��j�mP5UstЉ!Z�&�|�?���-a�4��8|IFAm�"QC^^E��M�>X���|4yy���=���@�������?�DU?B�|��ױ�p>�U�j��tᥝ:||i�ㅘ<3Ǎ(ҍ<Y�Ƙi�^���l{By�d����UQ�iҞ�p��0����Xp"��F�_�0���?���l�"��M"I �`��B�	=E�:G�$2Lmg��H�Z��$L-꓄�JcD�Qc%�	���I�}�}ָb>��3���g�1���KE"P�m� �G��H��*��).�w�8?��('�%��9�����Gň��8igO�>8Y���<x��J4�ga�z/�Ӊ���D]]�SX����@���G�!m��3,ύ)E��L$��L�pIU��*���-���6,]d������쳼��-�4����� ���~��`���ڣj��Q+)���d�.�N-�a���W������>�>�yLe{�M��q�A$��=:�A]>
>,��3ȖS��>1TAk	#�$%d
�zo��z
"$��2)��>D"�TR����c����5R,��x�GJ!^�,�k�M�]?e;N4z!��ꨢ�������$gT`H���l�Oӎ)M�M;��dA_4 �x��=���F �!��6�, ���LL�nL\Y'0������KH?4�x�Y���F��xXmz������!��ZA�\��艸9pa�#�!i�cpR���y���N�1w##�2�:�؝�R��73���	���(l��J$��b�A'����󰊦���-�d�2T�$����ʔ��D�#�)�FòN@@sF��7�;8���Dy64��>��DQ&I��x���0O�a����J?p�<'�,Ӗ@D|g��dp#��3*s�UD=���_q��ai�"�(iB�8��� �q�|T"���4�j, >^>,�Qw�����~�\�:n!�ۦ��+��[n�����h�ғ�PiJ�Y�>; Æ�@&���B��S�Hs��_ɢuJ��($�i�'	5 b��$�ã��V���8Y��i��M8Y`�%�8h�Ɩh���Lm��Uܗ�~�=ݷt|����f�,<@�I>m���h�g�VX9��ͺV�[sM�e��5$�n��0g��(��I�R3_�3.E���D[�Fy�p�5!?#��|�!3yS��B�O&̲�;�W�G���BE4��%X��$�<IK����HLr�3�F�q)�O���4��㥂$�i��x����$�������v�����[HN�b$#�3HP�TZjV8���wy�w�ؒB�jm"h�-��ܩ�͗o�o�,^�1�dc�Y��RI�eDO���WG*�~̘U��bq��VMw,���0�P��d�<��Z$��N��&~<4��$-(�x���PB<�0,��cEx�(;�2�ra2B����C�ÂR�&��A�ƴ�|D2d�g<Y���0�Y��a�!�<�p�����R��p�;��� �+�qF��h��}�j	r�k,�%�TE]!� �B�(����oѤD�E����4���ǏŘa����J?p�<'�<?��3�&LEGd�RH� �a� s�UD9�p�0���ä4L���>G�鸂!&�<�2<A�n>��A�IcGXb5IC=7�B�Jd k�t�B�����l���ԍ#fѝ��$��l�XYf��,�0iY�B8<\#�e{�-71���%�;d������������CL���Kcx�-h�Y���$�g�a&��$�AH<%	"pD��ba�D�&	bX�Ǆ�,�<"P��""pD�IH��%	����,�:$	$ �	8IHD�	D�DDO���$ADҍ8i�4�"a���	e�b`�"Yd����ı0�����x�Bx��D��D�H(�HH A,D���xD����D���[f�N�}�mG;=��O�&n��bI鯹���wfF�!|o{F#H�K���Ⱓ�g��;�zz�<߶���Y/|��W�`L�eAk�=Ѹ��s�Xa����֕%j�(�a��{e�Ϊ�M��n�l���Wq��4zDk�Z�f�����D��·���H�^��n(���;�b#޾[�9������:��^�ff��ҫ�������J�fnffn��O4����$�i��x��?`�E��l`���h��<���g0�~gޟÇR��l��!�
cϣ�"l��Hq3����+����憇���	��2�]���}R���oЈ4�0�#��i&���B����;��ц�<��?)	!#�N������Y�_�6C�_ ��p).�Q��QٷG	���5C<�x�G����a��J��D�4�N\{�BG�0���B���IWc�$�0�h�+Qh�\l'�⎇Q���;����!�8s�>��Ȧ��6쵤��u���^���&w�Ӌ�����]�{�񫉖R"Zl�8~i�]�>��hP<4D��0�#oT�����%��� ]xQ����e�"�x-
Ft�M\$�>�A��k]��R��J(��D�L4���$�'ㆈ��G��������I*����4���.`�UK
��]�����ʈ�~A fH,%5[�)�8R��J(��Q�I$<�"�UJ��{!HCF0h��
�N��H��=�<btDrD�˚Q4�]k�p��}���@1���R!�_r�������Z��=,�(a�D ��t�c� ����2=�I�P$J�2L�hÈ���L�ah�Qh�uўC�����y�Ҏע��1cG�@Q�T��b���$�I���HP����8��i�{���d����	>@�I��nC8���(�Ӧ�>0�b$�'ㆉ�:if��33����jy�C����z���p�p��ص�}���<H�8�ᢼo[cR|2�!Cv�#���PA�e�B�a��(����Q�-h�,`�gǛy�B�I	�&�҆5����A��}�SQAPS��D�sD�A	j&9]� Y(w��!���T��#�zE��0>[�B*�p���� �N�>T�|t3��p�f�i��t�! D�4�xN�Y�����J�k,̶ؙ\"K2�����m���Y��ӿ,O͸%�_���~pO��aX�D�Á��q�2!�e�$���k��>!��?����Λ920���.��@�[8ix{�;��Q��}_��;L	,��������Po
����zs���L�>�c���)�O0�|�QEq�v���C
z�t�{p��g��$N�t�i�Y��HĞ4�O0�L4��¢�J�0U�j��#�g�����3�C������"iZ>�Dp�|�GvS�d�ݤ��M�Rl��.7���&h�d�ȃ���i��Y1ԝF`J����P}�H�a!��f#�gȨ����,8@yr����H�e"�F}qe��'F7H�oŶ�(�w�����H8!$/����p�4�&Y�0I(O�,饚a�9��r{.~��oշd��z�F���*/�QeYb)�EJ'���,�/6�ز0��,BGZJM���wc�٭cv�nͳi�L'ĒI��a@�yn�b�f�~U#;��e<�l`%I����+�q�i�r"���6�Q��&�}(,�t�28TD>�G�y�e����Ik<Fxwh��У�@��<� ��q8�f��E-�����Z2QK^=l���]F��^D�(�P�L�ɕ��ֻ;����)C�ɇ!��C�(��4���O�,��$D�4�%�4�I�IuT�3>�?.��NU�(���UD9�>�����O!�B8���G�`|3B�4��A0�,4�D�q�%���߰|E}�{���Pl(�rbI���Ēq^(��wY'��F��%@��p��5[��0|��T0�t�s��#N�.
R�l�KFCy��($�B�o��X`o�J,KO�a���`�"P��||x~:x~~\�O̒X�d�UU�O����W�7sp�?�C���X���""��t�O�����@{�0��$S��D;9?����Vl�E�U��R����$�N���X����){��l��R 5n����cr�(�G�ռ6�����7F��o��V|XŤ�(�DoN<t���ŝ���p�ǌ4ᆒ^ ��8�&[��Z�UU��WM��ۣ�p��	�'��'O��8�)h�iOy'��� ��w��v3�:Q%��p�F<2��'�C����ˡ���lU��dw��D����YOD��$�����ӧ���AH�6'(|;�� a����$џYFi,f��3H,�B%(D�0K0�""p�"��,Ob:`�0�ÂA�,H�J$���"P�,舉�����$� �p88Q$� I L ID��"`� A�"H�pӥ�if�Y�a�@��`�xK��$L�%�%�:P�%�N�'��b`�E�: �"@�Q$� ��B`�"J0���p�"`�&	g*�$�{#�����B���3�@N�g5�	�d����l!�'8dՎaN�9>0E�V�K�r00�p��HF�������\rr�(MrN<s�hZf����d��-����ݝr�jG�Ϊ��|pzd+r�!�Փ���u��i5!D�Ԗ%�2b�P���*�M�`C�ƲH�8�K\�o]��w��_�=����D3y.��(����V5sc�i߫��Ƌ6`��..�}�۔g\�5��h.:E�S������+�+x��o�{{�o�N~�k��^n-Z���#�%���?���2����e��ju��c�y���WwZ�7����6�L�Bm�,Ӟ��G9�!�"����1ωr�4��L:a�J�ٻ�YpE_l���ƾ ͈ZhE�e�e%�md���oe��3r��!��M�+��D�ɰ�����f�5�o:h��1�`�H�m<*3RLEb�,w��L�l�8�lD�Q�沬�"9�%�+�v���c���v�*}�FE]���32�33wwkUs2�33wwkUs2�33www�������㦚Y�L4�,�$��%h�g�ç���W��h�x�m5��Bq7t�8�L��'#i*��YQ��$E'FF�'��@�1)!p)556M�U�c�i]��vB�T�۱�u�6%��d[vYc]ն
��px�#�a		v�k6�[aMٛ�udl�f�M�����e�&GH���c��Flwav��kKb�4�6sv��tԸ�l�ʹԖ;�]f*Aٷmt��Y�擛,�[9#���l����j��HH&�Mlm�U�ی�Z0�Gtuꪢ��y;Oc���źr�G��9pR�Q2C��n��Szc�e�q�5$�yb庫�I�/���ݬ4�2�P@����"H�ֳW��w�8WS����;����A2L��\9h�Z8�(���D3�ӡ(�҂>���J <���2!`�\]�D��T�:�,���!�'���nŖk�k��.<�fI������#�NJЯ��#L><p��0K�0�
?	��ig�;���]���r����q�<UTB!�O��7��f ��QD�AA��H�`�.�re��;��p��FJ�Ӊ�}��5�a!Q�dDA���>�&,_q�����v3y*��ɳ�i�:�!�w�'�{�O�Ȁ屺��';�����>�,�}5yrGH�(/��k�o3K���ab~:%�i����$L(����������T��6o	N"��w�-�UTC�� �ɟaڿ��8q���+%�}h�æ?C8���0����A�K��������;0��*�.��"#���#��H҃Q��I%'��|����|�my��K�}m���@B5J�Çy�M�5�[�s���ʘn�3��Ĝ,��?%��%Q�<t�0���X�K���^�ɫ���6��Cc0�.Js^u��c�
���Dqa�C�Q�c����P���vK ��,]aa��D�>�m�Q�N[tow0�I�2����WXك�D 8�GxPƏp��!�A"<OZo$�$��
c:��2��߇�Ys�sD��C�N�<����%ͻ���,gРħ�T�&
-a����)i��~Vy�}G
?�<`��?%��aF0Ӧ�i����C}�g��fyV;�$�@���j����iN*!Bh]�Hۻ�DR�N����->�JԮ��q�I�M�,(T����UQw�����9��_�ٗN�t+�h�׋!�i����՛X�_b���`��O}���x@чQH�N���>�N|4�M4���/M�� n���O(�Dz����%i��"іPiO��E�����)@I�Lc���Su6Q�-wu7d�*,���O��a�J����B"��:tÇL?	��ı�(Æa��Y���Ǵ��qT��m�����GN"XG%��ӆ�Y�l�F-0�Sh�.� aH��/ۃ�#ø�"@���J<_ò��0�8p���T|!{��=����k�ܳ:�o���t]:Da�c�����}��˧6ʡ�ь6"�)E/��"y#�E�ٙw�x�N�0�N�`�"Q�p�L4�K4���S$��$\�R��8W�2z\R���|�UQO
FBxh��\��DL8u&R(-XAE0�rܭ>Eu�!@y�4��{�Y�	>��Eb]e���?���%�4J@�0��\�h�N�c�pC�t�9*׊ ħ&�5&s1��x���u�m�����t)B.����Y�Y%Ye����bX�Fa�ǧ�������*��R��M)e��l�/���J7$�ËHі��"L<��	�q�p����V�cN��Ny5urt��R�H>������QGK_a�Æ��q���e��:I�]�UJ��(8��1a��%�F#��m�!��<�;��`�W�]��>�1�C�3IA�"��iӦ4ӧŉb%Q�4�K4�J�����""@Dn��bP��҉D�f*-���6i���-�KwlFX�؟,�y<��^�7-c��j.ل(�щ`���$[�Cf�����U�~��w�I6~���z����H�i��1�)���9��e�kg�.���T��Hq�y@a
�8�m�p��������E��(�Ũ����G	�u�9��(N:�(�  ��0�s�� va祅�T]?_�2X�s����Sㅅ��r���"�Ą�e�P`3�	_D�}EQ��ݻQ��v*�Ĳ#"t�{���fD�%��N-�,ўF8x���i�X�"Q�p�L4�M�c���ȑ�I��z��2KȂ���Ͷ���z�֔&o�nI�,��G0��w.�=C����8�,<eK�l6��YR��@t��H�첎Z�!��N�&L�S8h˫qg�2W6b=�0��)�����qH���AA@Y��}<0�y���̸���>E#)�u�e4���x�K$�<2�<�$�xӆ�pӦ�i��`�s�8X�%%�bY�:a�8Q"$�"""`"#Ȅ��A�"�N�x���	d!� I A�p8p�I8"@�@�@�$�""X��p� ��(M;�4�M0�L0D�	Ήb`�`�%�`�Ibt�,�҇�N�'��Yb`�g	��,�I A�$D�
:"%�xD�0L�S;�鍸����{uB���|��Ӳ-��&UV[F�	�k�M�|��bp-3�-���)��*��<�4�?|��r������ޕ{�Á!�xa�����p^�q���C���}-|#[v��8�ZzJ��gDM���n{4�fb�Cq�Uǳ��W�#����
R��0�Ջ������M�u^̆����霹��������\��������fe�fn���U�����ޝ4��<a��ibX�Fa�0��,�@�DDDA�X���SQSn|nJ���db8X��c PA-�(��<�b<:�;�4���@���#��&�ׯK��""fI�ih��&����u:t�B����:D�D�ƩX3�#���oxv81�,�%2�B�||��X�I�3��z�1a��ba�a��,D���(�M0�4�%CW�$O����v���U�J~�0�Z&Q�҂�eHAGQ Yhe��?~?�>�3ku���e��R����4��D?�?���[��xf�E�Lwf5։0.� e�bC�{���`��UD�<I���=�9-��s�x|RI���O��"}��ǖ�Ji�p����߼:@��xI((��M<&a��b%Q�,�K4�I�`��p���DB��Dҝ�2Q ��RŎ]�ؼ�w�9\Rd��J4݆�.��	7n�ϕW&�~��/Hxʫ�&��I�I��Uۅ��1���G�Q��v/�ȵXʙ�ϱ`�C�����yzi���Ww��9��UE�iL�f)82�G-��Y�PiP�ux(��c�n4��z�2w݈�
ĺ��qa��#���Y#j 0�WC���J<=����S��K�A�!D�����ӧ�Hrs�m.����bZ�d������?d/����?t�bh�ibX�Fa�4�x~<?{ x�	^�,�j���-M�m����$���#��FP�kxvȴ2����(�N�!�gFZ)yJ$����/��I�<���[c�ؙ<pd%H�qZ~?����=<�����ce�]�����!�.p�jUy�y����Pzp7�~I�p���8>����JF3�3��[�}�gO�DH�l?<~�����J0�Y��x~<<�R1�[�$f�������i��o����k��<p��a�[�Iu�P�NYӃ �u��i�䁐jsIY��(��ьڪd���IᒋR����a(�)����_3��P�A&i�W����>��3�^i� c�%�%x��\0������#U�"
i���'�ڑ��I��e��3l�E2��0��X�0�D�ı��
:a��i�����m̱�Pʪ�N6�i����^o�����P�q�ʖ�	H��g�x�`�Zv=�eS��mMd���gnv���B�F���b:q�9(f�:�<�*� c:1����{Nj����o��/pcG>�>GƑ|Q0��3 ��E#޼��嬁�a�g�Á�"՚���Y	��GP�,���~K�J�(醚a����Eu�9$vS��T(���mdx+]Db�l	-(���Zl�ȍ�$MȾd�:H3J%�Ll�2ˬbj͵�ыb5��U�O���0󼷗}������Q�IjDF3%�u{�n�na}��two�WS��$�����:��][�rw<;���.I��3���z
�׉,��i�6� ���,��:x}��t��8��)�\8#�)N�h���I����#������K��� �%?�|:w��A�s���n[7X�۲i����f��F�x�g��!S���י�Rf1���O�i��m��QO&�0MK4���0�L4��Lpr��J��m��B<�>���8����d$6��(8"b��ѿ�u9�$����a�˾g"��n��

���3��*F�3+�t"ԏ���>C�����jf
��3$Kq����YCK�<�t�8��G�XΡ��L�2@�1ҥc)6i&Y��0駏�4���Y��i_�ML�Q�p���l�v�m,��?|����b�!��C�E�h�Ξ!x�V`�GQ6,�o�N��WF4Z >�Ŧ��H$��֖�dT���Ŏ�<�k���LGC��D#M�xQc:E�憎���!�eP��:Q	� ���I,���������81�4�%4����x�'�:Q�4�L�=���&)˨)�qN�Kl����"~8zL=V�����QD���ftG"w��ޮ�J�5�c�A$�<>�8�~ tM ����>Q]C`��!���ઔ)D�'��y�\!�p����͂��O�@��AT�>ZKRt�(e���p�(�0���2�kmY�2�@Σ�#��	1ç�Y�i��t��	$		�HN	B#؎�&�h�h�M4ҋ4�0��%�bx�gN	D�������4E �$	b'JO�bt�D� I A�p8p��8"A	d	"%	""`�% �$	�8'�b4�K4�0��	�	b`�`�%��	��'K<'��"@��: ���x�#�$��I$�"%	BH�xD�0L���w��̜�s�}���[�k�>���sA0q��7Zh5�T���~���ՅPq���ހ��~zP�ͷ��&� ��fN�!�!D���0�WY)��g��Q������g�%&��҂y�P�����t.<��$�Q@��ÔH����S�~C��d˫�Iz���̔�2"�4�`�AO�0�\3r�~0n�%�"/���+�/,x�u[o,b1�`Ķy��'rm�q}_{Y��?.�Z�J+��2 ^ٸ�(�i並 a���;7�*����w��a,$��b�����ù��Pwh%�� ������crw���l��DůbP�Gl�2G(�I]@t��C����O���7P�h�HK-��2T-�e��?IoKp��sP�F\�2 q��@`���[
������FCa�K��6G�t�vB��xપ�e�4$�7I} ��$�'�B�Ĉ,$��6�h���M��wd��HK{k-{��U%w��9�o�.�=��gf�������gww|�ww�n����n��n�www_7ww{{��M<if�4MK4���Y��ig�}�+$���F7[�`��[Hn�fh�mt�.�ٴ����n��l�K���l�uJCA�sM��]�������.�k��e����Sdm$5�*h��n]�L����&Gf�stH��Wlml��eY[	b蛶)��R��f�lwv�ݺh�X�kvJ�ۻ6V�]���٩�݊+��Y��J�d�V�m�n�ew��U�I�濧F�?���10_��s�`X�h�z-d#���AяPB����?,����c����b ���=���d���9'�aƪ,e&Q�\�n�ĸ3�a*3�ϋg��C�C,��Ç/��3�M��N��d��� ��ϑc �c�8|3�E�a�1��G�W���R"Q���>�PT�(�/�LI6'�h?N0CMJ�U{����M�AgL>4æ�4�O�%p��4�K;fF����I#���NX�vj��&��Ui��aD�y���,�ll��̮��8xf
����C ����4�!x���OI��C�8�C��KD��;$�0�<��CA�ۻE=Ø8�Cu����g�u<�T}�x����z�E��t�$f��{�X�@�zQ�����'�${��Y�N�if��Y��JN�t�M0�8_��)�DP�MF���Lg�E���k���TX��J�I���.HO���۞8M4�@��?��5�*$�[��XlF��9���8�"�$g�d#���EB��W��
psR	�"������$���C:�!C�K���yf�0�e�1�j"k��8{2N��M0�X�&�i�D�(Æi���xxG�&�^�כ��J�nDN���Lc�Ga�����珖���E�Rh2�	�H�<?�1�EF᳑r�-���S�8|ii������yG�@ϐt���T3��,��a����Ä#���K�6�_%ڮL��:1����n�d�҈f��|��=��g��k|,f�u��AҘ��KD��,�K4�Q�N�,�M0��Z��ey�wW¹��2��Pʡ�AE}IE�pHl$��L�Qh��,��B�F͗{N/9d�)2q��bh�Mص��[��=U\D��}Q����iS�_~��wE���m�l��|9�7�E��&|է�8�A�����pQќ@�sN[c`׌4�y0�x����8�8�~<��ьd#�l|<�1�š�<��ç��33&�\�����������N��}�"�8 f�a3�9-,?�&�D#)��M���!	�&K��u�xw�Ic>>D"lf��`�xOY��?i�D�(��i�a�qn92����\��@��U�HyE��p�����M}�Nl�3�Q!��E���̜��t(�@3Q�)�g�?�Ѯ�D+M2P��[��<0e	��Gh�4O���_�KZ�mR4��c��X�b)�	$e$IU9�Ö=<QC)a�W��'0�A|�;�'N�D��a��DM,�ƉBQ�,�L4�tI�lP���(`�9p�!�U�K�N���\�i��>~��%*82M���9�^%��<3��}!'�s��C'��|�*���L\��^!ľ�,�R:%u���	�3�T�7,�A>�`��">��gY���$g
3��s*�3~Ex��q-(ߛ��}�f|�%c%[(���Ͳ�,���O�i�D�(��i��_�\G�J����\�TrIl�Y\�,�?x�����u����j�.�ݜ���2H�����#2�Ô��Ŗ3��
�+�P����c-2�ގ�/V����a��(D.#��NH�k����)s��*�65xuٺ:r?��8���Jw�E2��˘�l����7�'�kQi�n��L:x�L4�P�a�K4�G᣼%�er���k��x`t����V�f\�\+��$��ر���~���1"a�H-Bۄ��r6Q��5�ѵ]�ݓv.���Uq���k�<�1�`�nF���!I�R<�~���VwU�~h�1�Ө��Q�J\��)PƭCR�#��Ԓ:"a���Ne w	�N��R	�p�K��j%/�,��Xρ5H���0���3=��Β3�,,��83zYC9�Jo���&�����6�p�N��p�ϗ���N��8����Q��4�i��4�N�%	F,�Ƙi�=�Ǌ�S
�&6�i��$=�H'����n���Ӹ�$��$$���!���-�燂n����C3��dѐ/�|ȁ���D��t��*K��t��2b:�]���R���ä!�z��u��9�Q#&'����}O��B��4ϗ�l�~(��w�e}h��#D��N�<pM:t��	$$�xD�$�(Dâx,L0OLBi�4�L4�f�ibY�Μ$A���,BĒD��DL���%��'< ��I'�ÄI�AK I(D��@��"Y�8'N�i��i�a�"%��%��abX�Q�a%���	㤈�"'�<P�tD�Ή� ��I$�"YB'�0�0L�
�n��z��C�'�A�x���ڸ!}��ݪ����B�������W����ແ�%���//���y�x�+_�v'�.zo�%8�w̝]�>>����~�^|��DwJ2j���
/G���6
�`�EW�M���y'0v��\�g���=�'�����ځ�LΐG�.r{ԝ�W�V�n�d`��T�G�Ɠ;�y�6%�As]��n��������7ww{{��������owwww[�����ߺi��i�a�Y��4J�0�if�s��ē��������}4=.�$�<�E��3Rҷ�
"^\6��H#�g�&�h�o�4O߾��ې�vK&�6�v�pr@��Ǉ�a��s��,c@������yAѕc�h�Ff%D�s���qaEQ��8�E�3�|��m��=|^1�<i��0��0�,�N�%	Ft�4�K<���˻%�K�0�~�UqQ������و�1.�3�h��?s���N��?�f��\dfm��<$]�QQ�qQ�� ��Ϗ*!��8H�E(@�B�l+΢I�`��?��'säa��������!��s�'�fB�a��O@a����nzq.��!���}kK0�&i�%��8i�	Ft�4��h�&Bl��>{�?=��d�F�	k�6eO1�ܮl��$2~e��厛�����Ty�K��6YW-��&�RͻCn�Uq�S<���4�I�A�F��Ṃ���ۃ����ݫ��J���8���}T�� d#���p�� `���g�{|:A LEׇ�	�҈�qG�>];ܺ��wG�y��q��Ό�:AE6����GH c_p��(����)-�l��8�5)�aQ��w.~�!D�<0��f�A$|l^���,��DK4ӆ�P�a�LK4��G.;Q����o#�fG����8s�U�K��gҍ<�83:����n�3>a�=9�G$Y����fz!k~1G/^E�(�}C;j_̜"���=�.<&�4�O�=���Yie�O0��p��.1�P�2Đ˞��(������iGap�����nQ�:'�	�0DK4ӆ�P�a�L�����>/���c��0�4�UU1�m�8�;݈�83���ɳK9����
x%�<��z5�ٔ��P3��O[Ѧϔ��<!(YQR"��Ɓ-3U2_��9�)���]���=����hxC�Dq3a���I���&�RgS����D��d�S,�v�D"J �
�~��p���if��i�4�(��'�4�Z�T{�3��N���w�_W���1`y����8[?{v��7x�Zl �q&��ьF�6#���G��-C8`�LC%W7!DM#��� a�Q�AH��9#f�p�- . �n��y0���6B�ݒ��0�R�@�a�}���c! ���#`�iEt�M<t�M8i�	Ft�<i��j�=ʫ�W���b#d��B�ܤ!h(=�Ө�0�����fd\��h�5��r�o �P��H��)
��9�K?�Q3?~$�~ ������ٲ������x<38V/O�I�\�\�][�"\ח=v�.�W�v��3�u��9ؒ!���(��c�nx��P�����t81� �d<����AU�����#����������y��܁�� r揬��r�%�h|�P��p��®�!-��eU��������{p�C���Ƈnf~��|$�ag�"&i�4�(��'�4����9U\�q��'{\�D���F��o�\4��'=��C��o�JG���i���#��mo"(\�e�J	%Z(�656ph�Kc�V�ȓ�r)�PM���*�i�(~���
9���la�m��K-�qH��؇4 &s}�Ah��o����)yte(����K�"[�l��K,�a�&i�4�J0æ	�M,��
�{wk�C"�s28�3-%s#f��!f�Ҏ���}�im&�~�?x�\�%T�s��2O*.�QDVgA�$
/�M�9��⛂q��RO�]J����Wmr�Kh�j��?~�Nς�&Ǉ�8�l�$�g�n"C�a�2mo���&��C�$)3��V�Z8���;�@NL��">0���{�Q_}DHQ'�D��0D��4ᦔiFt�<i���2�x��Q^�t��E��[9���	�?�����O���Y�h�%�iŁW�{2��Ad��TY5#�dg����=�hs�o;����f���R.��E˙V�8J=��:�3|1�y�gOA�p����%a�)�"G���9qsx:�#�<�]3�=>F�n���SJY^�*���F͛5���忹������?�[K~w�����<�8� 	1$
�,N��A�e"S:\o"♮DCӰ�8 �dD[DE�d�"ȑdx�Y5�"�",�B��DE��Dk!dDY
",�"DȈ�M,���E��DYE�dZ$Z"-�mh�DZ!�4YE�H�["�"�4Y"�:A�-�h�$[DE�DX�"��mm�h�5�m"�dM�4i��&�"dYD#X��"d[D"ș�4kh�-�%����-��,�,H��im,Ki&[K%��X�-�%�Ȗ��4�BY-�ɒZD�M,�Y&��M���%�K%�d�ɒ[I,KH�[I-�ZId��K%���,�,�E���"ZD�-$�X��ȴ�b-&�F�D�-"L�L�Y&��im"YL�d���K%�i�dKim$�"[KG&��Im&�K�%��$�BX��H�H�m"X�I�%�K$�m"[I,I-�Kid�i%��[I,��K&D��,�,�KH�L�ZD��%�K$�ɑ,�%�im&�I��"Y-��id�Y&��4�D�H��%�%��ۄ��#H�H��K&D�m&���H�K"Z[%��M-��%�!-��ĚX���M2�Y,��D�-���,K�M-��ı&�d��&��%��Y��ɥ���BX�Kd���i4�&��KibD��	d�X�,�,K$��ۯM��,�-��H�%�$�&��bBY!-��-�4���KĄ�Bd�[HK$%��HK$L��$�I���M,�L��-���Y&�I��Ȗ$i4�M,�Y2Et�̍�ő�n!5�h��g2f���4�I����f�9đ����k%��md4�6���f�Y3��M��4��3H�K!��Z@�a#kM��9�md	0�l�Z�y�� m��b�����Di�"�d,�C�ȑd,�B�ۧL�,��h����h�93�""�"-�m8�2,��b-�"Ȉ�:t��h�m-�h�",��8�!h�[D�mӇHt"Ȉ���b&�",��h�m&D�h鹜-�k.�nt��2",��h�m,�g&sh���D�h��8��"-E�h��8�6�"h�MD"Ț,�4Z",�D�""ۢۆ�,E�H[E�B,��Y,���2-�"ȑ���[E�&�"E�4Z4ȶ��ȑdM�F�D�D�""�"�7T8E��$Z$Y��!m$Z&�h�",D"Ț,DD�6�4Y"Ț&�"D�di�dY�dM��[DDE��$DZ&�dD[DDE�H�H��dDDY,��Ț"5�4[DE�DYDȚ5�4,��Ȉ�&�k2"ȑmDDȑ#Y;�n,��"�h�dH�$Z,�"Ȉ�$H�DDE��-DDE�D,���dZDYE�dDH�"#YD���D�ȑdH�h���8nh��",�h�DY4E�dB��DAh�$Z5� �H���h��!��b"#E�MDE�B-�H�E�[DE�"Ȉ�""ȑmDE�"�i�dDZ"-�E�HЋh��DYE���DE�dH��h�m����m-�h��"�&�m�"h�"�[D�dB-�h�Ѧ�h�-�"�[D�2&�d-"h�$[D�mD�"E�h��#H�$Y,�h�-5�!h�Z$Y�h�,���"E�"��D�dMD�"-�,DE��BȈ�4�"ȑdDB$&�hY"-��$[DѭDE�"�-�Ȳ4�""�4Z&�DE��Z$-&D�D�dDZ$[DE�"ȐZ$YE�E�E�H���"�$Z$Z$YE�D"E�E�h�2"�4[D�DE�H�h�"E��Y-"F�"-�E�"�$Z"5�"dM�E��X��m"�E�&�"h�i�b&��Mȱ"�&F�&�"h�"h�#DH�E��[D�dMѡȶD"�MȄ[D��BȲ$Y,���0�kK��CPy4|��\�Z�7�<���,�i�lmkmJ�R�z���gnz~����|=����؀0�6!�`,�A��Є�a�����y�u�[�nmw�N��yzv�Q�G����g� ���i���i�bLph�,X�h��W/��l����z|�]w�G�ٛ6l���g�z������s?�F��c�f`�ԏ�׬f͛�g&H��[�����-�.��?�{_;�O{,��Ϳ$����&�g���^�mi��=���>�w��l٣ߛ�>�?��$vgq�mѾ�3=��[�n��[�w��)gMg�<Y�?��g3�gw�u�sp���<;�q��~<��=�{��l�;i�KEo��߅��}ng]��m�u�.�gn�07����6��a����Ζ́�`�u��s�������!
B��~�����PY�G�����y���7�0܉
$m�H�D��H6nC6�`��G�~���7��5��<x��������o�w�s{��ޱ��xa�����N�ǿž���]/��d,ٳf�|��N�N�ߋm�<����m۷�����������=��u7���@���6��>�?�<���,��B{����{�{q���y�7�w}�f͛�Ϣ�#^C��D������}/'��ɿa���g6z7��6�m�Nϯ�f����^e������g�qt��t;c�~F�����o?'s�B��;l~Fޜc`ݷl��Ee��ۢ���մ�l��f��h�>��n�7`�<F���Gf��3�g��c���H\xE��(_��K
$�B�H�u1�a��RHHHP�p�_5R�_c����o�3f��:~Glߥ6��g�{sof��>c�߳��/1�-�=��OC�w�:��>��:p�v��������ɾ��7ϑ�>���8��}�������M�6oG0��?"m�߻�m�3f�����||_�f���>-��۞������m��x����Ş��㕴��i'��������"ݒ��c�^��wC��>�uɟK��m���3�l�����GlD�q�E���+J���@���oʽ�����9�,�=����9�@�z�G�F�����y�x��f�yY1ȧ�Mٳ���y����og�=�3��C��~뾡�ugw�{���{�|����3����g]�>�m��xx]�7���������ei�g�#F�o[�����]��BA���4