BZh91AY&SY���p_�rqg����� ����  b(�                                           @U P` �{�%�YSϸ   bP  b  �w   �h  ce
 �   Z   ,`   @  ϾJ���UURB��J���!%R���DBB�
���T��	
��"�(��R��UDD��� iТ������PBAAQ�>@�[�P��B�j���9L�Q*ΊS&@5�wyUz#v���T p����@�8� �   hR��z��Q��O>�!ǒ� �w�EO}`>@2 2� 8g
p 6���@n΀Ocް < P��� �\�"B�)T
�%R�� ��� �9��`���� �z���x $��� =w�}�����` ��}�*� /����|   )��
<��/}�  x���J�� 6��{��{�>>���;�{� ���W����� ��=���z�� � �z�hYB��$��AP���E/�C��w��z�<��}� W���J���}^`��0y 9t{� <��D!���r����@(��  =| �G}�����C���} {�@���w� z��⢏ 0��z��  r    7   ԔQ)$%DP�U���� ��n�F� t� *��� l={�'�`��*\ 2:���   x   ��`#u��xy�)��=�;��n�z<�V�p ��;�9��r��   ��x   P�*B�UR��	< d�709��t8�wPAp!�&�; 9�q�D� ": rU   �� �B�� �v �nE$�k��w�@�!��7H�W ;��u��,� >�        �@
T�L� 0  &��hш��D���0 &      i��I�)L� 4b@� �M��RF���       &���T�       
��ңQ2`MS�j4h��0�<SM��=��a���9/l��@��{j:��]�A�_O:��珠TE�J���p~DAW�?�:E�QO�AE��SO!��W�����?��?�7����C���y�>��v�"���UDp�� �+�d�C�ᠤ����L�U]���~o=k����߿���H'��	�*�ͅC�dP�`P���y0m�C �*�ʡ������ �����1�Eq�S�D�	�\`�@a�N�H��8�	��UaP�@LaA�aT��������ȯ,�2�c
2�c"�L �ʡ� �!�(��8�vl`1��\e�\a�q�`1��t�2�c���c/v\`1�q�zce�Yq�q�q�q�q�la�d1�q�1�q�q�q��8Ì2�	��2�c.0�g2�!���c.0�c���ce�d1�q���c�0p�2�c���vn��i��Ce�{2c	���c�2�!���c.10�.0�c����!�0�cc�8ˌ��ٗq�q�q�q�Ca1��q��`1��\e�C΀�d1��Ld1��Cq�a1��La1��\cL&2��c��2�wa1��Cd1��C���d1��`1��N��&La9e1��Ldq��\d��q�q�`1�q�q��:d�Cq��\e�e�a�aƘq��e�`1�q�Lc���c!���w`1��Cd1��̸�c.2���c��0=0�08�c��c.2ˌfSLd1�X�`q��q���`1���Le1�gLd�e�\e��\e�`1���Ì��p�c&2�ˌ2���w`���.0�0��c=0���2����2�.0�cv1�L��c.2�.2�.2�c	��gq��La1��!�2ˌ7L2���.0��c!�-�2��c!�)��08�pɌ�00��cِ��`1���儘9`D�S�DLe� Le�La�Qa@�G�d@1�GE1�C;0� �0"c<0.2
c
&0*c�2�v�@L�L`�Ld��\`1��EG�T1�L.2��
�2��&2�c �vLa�L`�D1�GAq�WQ1��
&0�� ��*�"��.0�c*�0�r�����)�
�ȃ����/f�Ld�D�㣮^��Z�����َ�;�����,�6�3W���i�wNX��.G��ָqǔ�O�`c���u���xw�e��nw��NC�N�C�y���rG'S��w��38uCcT����n>
��i=�����s�Gw [Ǖ�k�U�Ӌ��k#E�u�Cz�b��n֡�{x���R�k5��s���{�	���Kcmɧ{���K�b��6� S!�;�U��]��н:�֪�4��� �i�F,Cg����m qCP��oVw$�L�����B�����*��m�y$��`]��0�_r�Ni�G^���<�;^Z��ͥK��}�ӯ�d�Ա��'��}�R[��T���}tjio:�YO.�a�^w�{��8GȰ�f�`�l�ƖP�"M:�;U�Q��m[�$�㪜ߦ�#KT�V��f��[��pӠ+Q� ['''F�L�aYvv�ټBG;U�@�n�7F��`bF�ݺ�.�7F�ػ�[sdQ���wy�@��9jg��{�x������H����Y�j�9�q	�3��d�
��܇��ϳ�� 
S��\�&��yΎ]I��`�xw��KS�-Z{��19�V.�P��k\Q�͚��?,2�pooL�:��q��1��88S�	�3��Dfwm��sq+u!d��gl�r N��5�8���V��Mhst!�glYfH	1t�W�0E�-�$��9���j�)�Ѣ�z���U�z�l���.[�a+U0�Gp,�b�Xөq
x2���d�p�>c� ��ɭ�C�h� ��A��WN�I�t�ÆI���W{y|7u��;s]tCH�ٗR*��6\yݗ����9Ӛ5ݏ������ur�����f@^s�d߻T!,s��<�XR���H�a���G�e���&^@�r,Б}.oC:h������4q��yhz��D��3�h�5gQ�8�������Q��}I6]�5(PDl�<��ʩe�RNZagfL�a�S�F�^[ؔt4+\f�ܪ(�wyI��4��_��;`���!O�]M�;�2^;ϧ^�Nod7���3n�����#5cD�K�s�ۋ[�
�Kf����Yԑ���.Sݺ{j�T�5oX��1�u��1'{�@|2Bw�)��Z{�X���D�(K1�-*�܁�І�;��|�ø��#v����]�t����n���m��s�����e�۱P�l/��׻��k�w`&@����g.b�m}3�u�]�CNhƃ;0����GQ�u+Ø�7{��Kfr�f�}�uJd���f�7H��st,�ӫ+��Y���R?�ԠEq{���tY��wm�ٛM���ٻ���b��FC��ۧOqȭ�h��2����D�;h؟�9Ms����J�DH0��8ܽ� �aeXpnU��ܥr[��M?���H��נ&wpE/<Һ������j��J@�Fu�MKf��z�n�8F��3	�swg4]o[6�7*M�y�-��{����ӊ]'�p7NO]�.�ٲ�j�ݑ���s�9F���r�{�w�Q�����y\ѣ�ei��5\�Kxc�Ŝ� �F�
�[Y�=�Z�-�1eWu�اc�;H��=�v�G;��	=v��m��<۲�*��'�O,���f���e����me�fU+Ǹ�!2�)�I
�6N�ě�u�ø��(�
�X��N�ې��=�L
Ϥ�[5�&颵.�t�2���w�(����L���Ɵr圧5�	9�8e��S;�=�i���뗵N�Vd/4Y6�6��٭�q��.�p�����gAz�T�ͥ�:6*h�>�N��Ew��� �E�Ãy�*Zo��e��1���p���u͘��Ǳĕ.���`�lDwu�`=V.�%B�@� �;Vn�|*j
�ΆX���g.�S��v�ݫ�աݮ��C.�-3��B��.�;n�ïqW7��>W��҅�к���3�o*��$���b�F�w9���{�s<�ʎ^�qI Y��Ѧ���A��r �rǃ�*�(N�&�=�f�����է�IE�Ħ,�`�dchb|X�[��RӤ�[C�}�4-�s�.�{���ӹ
C;�m�tR3c ���ŗ\���Q�n࣑՜L��8xO	�bI�k�b+c��g�(�ҮUfT��I���S���`p=�6��k��\/U�f���7n���l�P�,�$��WN"�t���T;�5�Z��-�I痏I��{h�7��]����i�D�q0�Vs��:�;��jN�1�Վ��۸+M��+��Iԗ=��N�܁�ꛪ>S]���eP��5���D������PV���1mVv<�E̕>�]`T�f���۝_iP����sLO܈����6��߫�ƹӘ�
(d<d�m�SY��iC=WN[3�m�\��OJ~=Xu�;(� ޔ�C21pwn�`od���.C4��*m]m#���=Е��퉋�#��\z�|d���$�s[��@ЭTpݒ��f��L����s��z���ں�[y9��n��S*�'C�vm��04L����M܂c� �Rn�%O(9r�ۄ�4��d��\+G(�գs�`����tkA� ;tdQT��=]����{q�l��,k��h2�:;r������ޜ*堷',�:�tjg7���:݋,]��;X���nKV�k{��+����zb1�%���	ײ��O��$��:�F��ۢ {孅�H�+1B�t;*���p�\��>G�ce��K�ԺY#�wt���W%��qS^V��R�ǃ�ew@y���|�[b��%u���3N��c���ד�gfK]ף�Ƕ��d�<&�?�^O�3Td܆��gd����W�|���0p���tí,�~�\�2nS7R{�[^��ާ�:� ]�i���ۼ{��ڰ����!������-�6���bXz@�q��nB�rt�{��m�[�>�Ԩ�p�nY�DY�|C���d�5=[�m#B������U��NX�*x�N��z��m��y��8��(�#�M˰vS��c뜀9gPf���!�i��4�5��&$�{�퓐�H�yf*����;7u�ʄ6��=z9jKGa�ya�rl޴�б����k�0k\!��N�%�4QTy�\���-������!�i�m�	��ᖍ\�	.�B}�-\.0��V���$�)�in����>R�9&�Aq��6óZ����}W�w��5^��'݆�w);M��
��0���@�°��%�u�S����{^�2�T��/p���F�܅Uspv!s��9�Stt��m��t�8�>E��Nr�1e�gv�6�<��\��]f�ݏ�h
�Qِ"����D[R	ٜY�ō�c7�n�.j�]a�n �˔��w��`s�Gc+����>�ȥڨ�E��+�S�ö��t=C��*�9�Gշ�(���M����;��7	��3I�g!�9�q&��;�k��d9݁��66�ĝ��VF���.���gc�(��v8uEHc[p[�%@#Eg-ɒ��h���í�{6�){.ѻ��K��n٥N��#6<T��ֿ���R��Yc�	�+��l��\��{:&�a�����*ܻ�k��7^�\�9t����`�qelY�;����JA�)�=7	4� �3_6'�>�-�]��x7:U�)�ݧ��2�;~��O�W\�<l޼ӛ�~HnpkP�&��'sV��=�^�.��}�"0���Hex�����ֱր�gi�P9u�JEwh;~=�t��PPE�HIA�N_V���T��߻��f����x�~�g@��;�ت�V]o21�rʍ�{
�����K4��y]�M�C��v�ͦe,K�������r!���ݳz$yYi�m9$�+4������jE��$L׵�w�G���nu�����{z��9�sx�3h�v�v�8])i��j��5CQdF��%�״�r鏯Q�hX5�95`�&g�����o۝6�����頉Z�cZ0g���x�����ir��.�����h[�(OC�R\�I|��Q��;����n;�4�*���s1���n-��)��FIP�{1	��LQ�3.t^C �V��׶^.N^ŋr~oðN�Gi��yw�k��w���gur�w�U�sW���e[����)�0�U���Փ��2{�{�l������`�M��vG��UM���w��޸�:�Ўr�3��C��H�|�i���ٷL���v:�Rq�lw����0?�xc�ӉN��Z��Q9�1<�N���U������"I�h�XT�Z�Xv��sל�le�.C~���Մ4E{B6-]�4�۲ L����Ds�A�)۸�u�v�N@��p��x7F��&~<v��9����4�;�Ps�5!��!0읜��]w6�my�#L�ky��m%��a<!��	<�ӽ����m7��sKZswG^����^2�@V�S�kw��B<��!+n�#��������0s�{�ί9��U�I�[�����[ݫN�}\�v��&��<	�Rӣ&WF�Kp�g`��%e@�p+��w�x��0��m�e��n���� b��S}q�	���ݏ-�>ý���A����8�p����a����N��tE����pP�e�Ӟ��{ͧ�Pswqʳr�o��7~��7V��t��m<Μ<�����A\�WL�7,ၐyT���:�Cc��b�7~��+k�#p옟LCX��$��SK�C���=�x�ɫ�����W;;�i���7nX�r�s���N�/�����T�=1�2�����,�3D,��
-ٮ^�u�L�#�NG5>��l�v�f��].��H̀m#^Qx�֖2��� �gq͚�!0A����L�� q�f�bG�����8YΫ�WNY{z�{q%)f)��*�k�\T�g*�7r�V��\lR�����x��;(ㄣ�"�u��]�ks�3��oG^��g`���,��'��3\�	]��W�I��R|3��`h1Ý����oR�ټ�m��r�\v���\;�-�g����62B��f����Ѳ: [9Ek;7��j�#� �YӇ*�e<�7i���l5��+�5���.���:h���9V��Z��Zۓaǌr4��ض�8�u�9p�����\wr[�u�2P�i�wq���*�m�;{�擜o>�e���t[��k�̓+21��3Ov�5�����6���p�\��8U��N���jLY]���&�I��olYɧ�0�nٵ���J�	ݏ^7ypz�̷͖������e�r~� ��ݼ��owD�q	�Ar��=��c;�c�r6Trm�S�9����1��gqbȑ��N������Q
y�غՍvPחw'h�rs����-��"�N�j0K�j@-wG7 �|��4)r�TS�s;�}�FR�����&�M�Ní.Ѐ1�s�+;7f�?2��2&��w�����gk�Q��'Lͬ���&�z�[*rq��lv�X�7;1��q�̙jce����𛼏b�t���FQ�}Tmأ<����g:`-�!!^C���ָ�n�೻��M�4��4g;*Me���L	�f�L�i�d�
���M���O�:����L��s�&����ɓ�<`nɳ�n�R�j�"��t���3r�d�Ln����ZE�#�O-XCY�8]Мy3g���U�;מMy���H%ѳǽ6mBr�`��Mc��)r]�!�φ]Ɏ��Ú�):�	�2�䅑�P�ɮ�V̗��Ǹ{"��b��l�:@$�.1nj��G!�Y��
�9"�lz��[�R�����7qc`Πضjr����dl�S���';��Su��N�r���;.06�G5������!4jX�՚�z�1���r ������Ck緂Tas$��/����Nα�={�(h�6".�xYJ',ϵ����a��1�$)݃3p~Y�%x��%+��R�5����~����J>�n�o!��K�rw�7�5#�wG�����_�.����yo���L��"����貦M�rbk�������r#�x}-��E��L�/��|;�B��>4�>�7��k<s��v�'��.�)������'��8=��`�q��u'DMȄ?]�mP�YT:�P�Fhۄf������k<%�>vD�B�یB3(NA!��#�����l�ޚо�T�qi�i���	�`H�ŨG��-��5�f�ݸ�����_v7���4N&=���E��`ju�ܖ�P1��i�Q�nUZ0 �/�v�����@t>ļ��5�CN�r��
t�?i~H`%+�t6�� ��4���(Ȣ>n�X�F���˔��۶ ��TGĽ�x�Ђ�dqc�(
]�E�bIW�h8��3��b��F��8%�_c5k�&��g"��"*���56~���K~��>W��اk��v�B�6�=�����J�Y4ǹB����Zz	�A�S{�f��ŽF�}&�f�o���,w'y죙&�y#go�}����r��-��Q:aZGm�/��d�Ote���o�M�ĕe��=����}�ާ�Of�Ѕ�.�|��4v-�g�/�g����]86���+x���c����Nؘ[�Z~.����޹���Ncu��&������6�i�=��P}v�����$a��\���T�*�R�hi/����o����6O�`��9��~��y���=�]㏣F�_\(�(J� #B�R�� �#J���R4�R(�Ԣ��� ���MH�@�R�@ 4
�B�P!�@�%"�4�"��P5()@�R#�EJPjJ����*P���	H�SP	@�T@��(*�J�RJ�4ҊP��SP	JЈj��	J P#@-*�@
��"�WP��WP�R��(J	@)J"Ъ� ��"P���P"j
@ �J�SP!H�R 4�� 4 R
� - �SL H��0��?��k?����-���9��.�/�Ą���h����-��Sz��.�x��	�@��0����D'��7RP��S:�n|������_�:V ~m�!���e!{�K��oQ�-��`�h䱖�pP���,Ie�aX���S�|�Э���z4��51��j�6����6L쎪B�2���k�[`���x�RޔsOI��&�5���ǌ�@�<�X�q��pX�ĉ��0�'$�_�_�e��杬�{o�|����/]\Z��by
R�A
V˼�Jo˨f���y��]3�O<GU�9<K���B�i����`p6�
����<@�p
��Y��Ƀ�.LgH{����%�V6��3�G����
�@��|��ao���角�ax J�!%�#�R�Cp�O�h�H����m��L��O q駫�y6mX��O�8���� �
�:�=���}}�@C�o�ˏG�����|_H��O��}"@������������/�'�O0�ŴY�� ��`�F�� վ�#�ӿi��ĶoХ����m�i�K0TM��oj~ﻸn�D�SS����哵m'������:��x\�r����~X)��e>a��QO@�/���,�hI�e�ś��"��8۞~�|��<��xB����O.#Nʖ��y�'|�TB����=���=���$}�=��1�U�j��+��{:%��z��<��>�lޜ��ٻ*��������ؙ7�g�a�=aɢ�w�w_{L:�D�p�Y"�^{ڳ_�73��Fr����s��g�nS�-�wh-G� �b�b��f��5f|�֦��1eM�>]��?]G���]^�~�����(z����ܯ������K"��v��������^h�˗�-��1�u�Fyߋþ=��:<ݕ���-o;�s%�vn��l��n��zO�+�.��{��+mp-���͐��i)��������K�ޒ���x?bC�0���\A�̣����o"m�7T���o*
�G�%�x烼���^qS����KH�}"<ry /||s��gC�S�q�Qw�@Q�I�sA+76�/��3�l�7=��̓=0���W��y�[��-%xMU�����SX�㝎�<�S��r�L�pq۷nݻv�۱۷nݻv�۷nݺv�۷nݽݻgnݻv�۷�ݻt�ӷc�nݽ=���~=޳L�w�~q����=��}����D~�ա����ъD˗:���iފ�ݩ��o�~�L�c��k膮ĸ�{�G���RkL>9[4?_�7�E#�*.�ಙ�_*�G�Fb݋�d�S\\ɻ�+����/��@���i��f��F�
�M�l����^�{��`�ؼ���2*0�|�����%zg���<^�ϻ6˝�zn�A[�9��o�����a��(�خ�����Y����MnM.<�Nｃ�u�>�;之W��֤�h���{��l�:X�Y�{���/iƣmx�'�{*���rAC\}@�y[�Ы�=w�._�)�j���a�e�3�d��-���|���`�7��!k)�-Mo�ݛ3��۴�r�`}w��k�|z+G-�\=�N��w����������i�<��͜ǭ�=6�œ^'�m��{q��ѿ`T���s=�$z�=�OEoI:N�\Nxs��݂����'�# ������`̞�͞�w�Y�n�|׺L̞Y	�G�e��y�n��X���^�~��w�V7^n�m������f�*o����}���ٻ��]�R�����?:]Us���D�=�'���zx1ڮ��}�ٗ�}$x���Q���x��@8��L��y��J�}��ǐ{�;w�ُ��N=�۷nݻv��Nݻt�۷own��ݻv��۷nݽ��v�۷nݻv�v흻xt�۷l�۷:�U2�j���ن{��c~��	�����?�D`n}᝜��1k�ݞ���9�zv\��zك�]��	^{�W�2u�^�s�N�^�陽=#��C���;�/��=���(>�����z���=��^�����Z�{���/W ~gdR�tj���7u�x ��{˺׍5,T�����';-H4M�����S���il�E�LZ@N�ó��3}'�)Lw��_���G��t�̓E$\Z�~�T�[᫖E�7�Oo[��Ň�'��w�3J��ra����f??]��S�H����X�~Z_�O{�����f��C�UO�#ЗY��T��ʯ����4>x�=�p������ùJ�d��n=���ɦ��w��o��P��^f�/>�S���N�s�FJ;�E�EjK�}��a8ě�e ���Zk������j����,w#���G��#:{~�l[*�6��-v�,�
C���w�R��0z�cx���~�;Z�n^�)�l����`�ù�kѽ�.���8q����d��CՄ�)��7n�)\䷻K���~�٫�9��,<�΅��{S�����}� �=6��W�<NA��6�G_{W&��#���达*o��>������/z]h�WJ��;5=���%��g�ٷn��ݻv��۷nݽ��zv��ӷ�nݽ;v��÷nݻv�v�ۧo����y{=�FE��I�:Ɇv�lI��k����F���j:m5/e�Ȯ��e�H�cz���E��"����E�1�/�f�?cN���&q�?f���x��^{ۜ���q :��>����`��Gc�8����<��_np��r�Gw��}�01q�~x=�j������o��No�|W�9I�]+�f�7v�Ԏ_���7-\����=��c�s��A�k��#��w3ٳ�+�x��{��l���1ݳ+��nx�ٯ�d�����~��8B����i}��^L���Ķ �����v]���7Q<�|�O���z���0��bgЮg�ʳ����Yu��x#�}:x�M;<6k��F�ۺ��z9dl��!�5�yz�<yO�|z�c4����|WeM�w���=Z��Bg_�ض��q���$��kc�C��λe�nx�U"H��xuY�Ճ�@�<7>���{��M�G6��?t��u���H_�c�UO_KN�n�Z���Qv�����y�=�ӗ��-@��]��A��ή�3�a���`N���+����$�}�{�6�hY�-R>=��	�Ѹx��^8I}��;Gb��:y)����Şxo�%n��'�G��3&��8{�9�{�>����s������nݻyv�۷oNݻv��۷nݽ;v�۷oNݻv��۷n;zt�۷oNݻv�����۷n���?s}�96��4.n�vL#K�_s�V�i�a.���*���'�2��|���=��Qt0z]Ƹ��YK��0Ay��?x?
4p��<:�ᠴ�z=y0���Y_�phYPX�p�"���������[��ўA{7^d�Ǟ�ߔ�;�p�s�(~�w/p>�cA���%��A����y��(�fH�2�>=j2(0<�O������%�LX!h�<q�	B�kY����w{�`�u�K�dd�����L�t�����C���iɛm��I�Z�'�\��MI���Y�,�2m%ǧ��_,��ů�"�_�X\	%��㾔gE��q�<�@R�I~�p9;������ܩu�v�����n�^'͍\��/J�L��ұ��Qx����N�d؟I�.��^�x��ro�Mw| [�p�TL�l�G\�������ɻ��O^Ր��৒[�Y�x�Ow���e�ȱ�A��F%
����9��'��O�g�����Y���17t�е�����9��o`�g�u��H�.��坓�s\���Wz��}O$�}���r���U��{�!�C~�Bf=�of�8��m��A�,���$]�wF}�9��;Ł	�6c��x<�ݜ.�Ӿy��}�`�7��on����]�nCſ�����۞9�3z��g��˷���۷nޝ�v��۷nݻv�v��÷nݻv���۷Nݻv��ӷnݼ�v�۷�����n{=��A{�+�'ύuh�Z�z���y	䬹�m�@�!��/,�ve�!��Ρ_tg����C�y���9N^ר\X�a�6�M�g���+30��?h����`�'))�7 n�qLwW���)��_Yr��o8��W#���OA���&e�����tK�j��s*�뷴u���lF�����U+5��16�xQ~�f�"=9#�wc8��'�8VƬ��n�ِM��b�M�q&�w.�u��;<'�]���������٫}6�00�]�q��y���^��8����tGZ���
��L��_)�C�𻳽�q��w,��n�>�����:��O�:����޶[�{���f5L��w�9͓1���q�֋� ���{����*�n��4��w�H�n�J�"7�p�r����Z@p>��o�.=�૏�V�>w7Z��k9�{7��>��vxD��Ox�ғ���5�=<����J�#�V�x^:���'8I�zs(�Ⱦۀ���n�l�Ki�;lòjc���1A�G ���Y�q�;/{��P.{j\I!+���g�a�.ٍ?k�x��^3��o��K��.���S�輫��5�);�����nkqE�Y�ܼ�l��ÓѰ��^������|������Ͼ�=�k�L^�U���������y��g����{nݻ{;v��۷nݻv���ۧnݻv�۷n;gnݻv���۷oݻv�����{=��VR��Z1qsFރ�S�����eʖ3.�:<~���^����<�1{'��l^���f��|zV���+�l�w�<9�(�p{PǺ4��碖<>��po�?"�)�케�"�WqM�e�t{<=�Äv��:��;�.���I�R���{����/O��ט��6Il�^]y�T}��fz�;8�.8�O�����hw.��W���ٗƕԏ�5�L��Os}�`�{�Gt����I�[�G7u,�[No��������sL��v�<���'{O�~�p�O�{fy����_'�L��"]���ц_S�E_s�o��"���}�Q<�ӦQ��[�y.��*uLy�Kް�ub'���{��������ơ{���S_vr��~&�~���Dqq[��>/\{��'}:,�
�0k��>���]>츽����e<�ƍ�Ov�6��>�k�J��<>�=ö�K��}F\�M`v�^6��IǛn����ߓǽ�����|��hz�Nq�{���{�(�;_bԩ��C1}���&�{:מFS��e8���=���{qp��G�c�tt������C��3�g_��1�s1����	����V��%.���HXߛ�'�L=�w�����L�{�{Y(Zy���-�����}�O�ϧ��G���z�wף���o���ρ�n-��s��ۭ<�v�{��8�۷nݻv�v�۷nݻv���۷nݻv�۱۷nݻv���ۧnݻxxxv��ݻ��w��Q�,�����7��N���`�Ȼ���S�!R��l���)h}<�S^�����W�|���E�����\'�wr������yg{O'X]���������3�ko�-#G���B���.2����|�a���F�Y�8�Of}��z���u��	�.a����O(��Z�e͂n�(��y�dłk��4:��>Ѻ2!5zOm:���i~\�~��o����y6v.���K�Ȣ���=^rxz��>�0��,y��:�d��w���O�x�������m��3����b��9:}7`g2aP����8n|��I�gSn������_{�Wݞ���溧c��F/b��z�.����>pÖ܉��LÝ���~�(n�:A^�\��e�fK�IA����r���#���`��A�7����^`�^r�V��xb��D�g��g��lŔ��������L+��Z����*��M$�}�G'�̝[�/�;+�=��g�O���,?	����E&���0O�\���f
�����A[%ξ�o��V�G7�ƙ�����Y�!b�J�}���`o!�4m(ꮚ#ܽ�,O0�p��[���Q4��3�Q��]j��qg�t�B����1,j/8��V9� �y[�#ɭ�ȫ����@�v]�Y�N�8Bg��q$�@�n{��q�ws�������q�v�۷nݻv�v�۷nݻv���۷nݻv�۱۷nݻv�۷c�nݼ<<<;�v�����&,(%�Ǻ�޸3��+{}:ĩ�Γ�-�{Ч��u�=&����^+��x\�U�H�cv�Cӏ��~;nt�.�^��ގбO��|\	H���7�e�Wӳ��:�;�޻�3�돻��}���^��j�l��az������o�'�i%�=m9��[|.gԉ��O+��kf[y$�L9�h3O�z����fL�J��%��-V���8�.��k���͇�>���!&Ɲ&OU�{��uxBA�R��/n�p_{<_�𙼞+�?�^����Wq�$lc��vzʛ��_�ٛ.^���
0��x�-{��q Qf/O7Wq=p`>�e��{G�*%��Ȧ��O���ں���"d�x:]~��ʳw�3�ɟ{|Fy������U���k��>\������o�}�d� �`�YG>~�s������<�W�<���Y�ݻ,C�J|�+'Mͼ��Q�Q��_�8q����r���Gb���I�{��M����������vq8����r�]�{f\�G��u����y][�ųFw�8퇱��d"�
/�,��#�ۼ�r���x�;�������E�{P\{��#��}�L�&.^Y̳0�ɒ�靅��a{�}������h}3Ώ���h�2D�����m��c��& �½ßs�_7 ������%7׳��ʆ�py�i�N���������O�#Wq�q��tQ��S�[o܁�Ov{���eUn��͛�k�k�z��5��Gw�/l=�w��<oA��1�Ζ�ɌzM�v�\es-Y|Ώ,o��y���ܞ�����&ն
u"����Xٖ=˗	�qM�q^q�`�xf\&x����7�����Ӌ�k�i�{�W����/�����Gu�K�;;�D���b'׶�{_SI$�����L���gb)o�H��R����{F�4����vY|$��Զ�74(u�t��/vuѾ�8$�_��!2Ӊ���M7��W۶�vU5�I�澾ű�I��{ټ&쾨G���5���}6r���1������x%�����s�3>̒�q=��*�7.�n���2��I�r�SI�<�����.���_z{�Ġ�on[:r�w�c�9�zQ����KsY��9��^o���vi�?C�Ɯ�zW�Ry�ம�I�� ��g��)���k��!/{5g}g|������0x{��"�I7y��7��1��� �A�7�w�(l��$�}��9�yox]QwKq�[���Y7�h:}��n���{<<0�E;��ˇ9畗���N.������}�/Ь�\���Ϗ�a�3�^�y�y�{��g�z��Eƫ��w:��۞�߾��O��}~�TV`��G�{���}+�}�C��w�׾�\��1��GlK��ڛ���|/�@�Ǚ��i��%��u�=z�*������
z��Lˋv�Wl6f*�tb�S2�mK.Ñ!(�
���B�`��]#�e1�@�lݫm�H�afݫ�Z�7l�W4�5�5c�"�ҳF^l�,	��Ѱ��N�Zq�]X���[��a��U��#4�^ЁL�J]E�:��8�1,Zj]��:a��&�l�+uR��33�B��`pY4n�W��Z�f&3!w�F��(ǖib�bE�cf��0��KY������v1FJݬ�Y@�jk̶[Fmx2��F襭���	��F�եXh2a�V:�EJ��e�!2�yJ˝���3n�qRX5ݦ�!Lj:��*�mpu�v&��f[n5ĵm�"�&&�������	B�I�eCg��Rm��s+e���.��;L��A��JV������	�U)�3UL�kS]��rLA5j\�
�8�V�	Hhh, \�N!I�#\]Ila���)aG^R��m��4��j�n-l����$	ZQ�csȩCJ�B�:j-��k �P,qt��nvf��C����+��si#L�6��I��ɂgl�R�GE�X:<43�����xz����dL�LPŵ�%D��ûAF.��xl.���C��z�Fl�s��r�����J*m	�-Ih%����e���m�4�IRb���4��R���m4U,�Af��i�*�c��v��smՔˁɗ�1J�bl �$��J�ud��7VҲ�Z�$$�XMce4�j�C4PR�0�1���+��ڔ��cB^m�5����@���p[�iFT��7*b��*El���Kb�bnk����ʑ���E�0��l�2�A˥l^�-� ��ՔFf���m�fmb���җY�ť��e��V^�� i�]K�%�Aҁ4�6HhF��M��B��Q�9��y�R�tc��67k�SYn��Q�	�5�J�F�U���W�G\5�&�fa�3�e����2�r&��*��;vc��ү
���n"���fKH^F��u�Ke2�F������af���h���c��̓Dbu!�[�X�鉵50G�����ar��7]nIr]��u�C#.9B����N������ƹгZ���^
Z%����$4�u�nmҡٶ�s���5�gG��X]�+��l��p��oh<��[)K&�HB饶j���6��\0Vٜ�IF2�vi 3u�n�\�v�WYqd����K���3�k�JV�+� X�1Q顈���q�,J��nQHi�
�b�s���e�Uñ��2�mt���Y�!sRn%�h䎈�ٙrR	��)P��*c�*'P֛:7!�t���in"m��s&��i[1�5�5ZDy�3��56.�u�sm&K�mn��!��I^6������ ��^Ke���`�s�5�Gcd�;Y�ؔs�hL�-�l"��,,�m�\��<L(.�6�B#��#��]b6��8f��)J��K���V��k�IS�a�j�Ë1��E,�`�u�ZJ0�s���r%e��V[r;ԗ�lvEYq������y�F�uЃ�W�b�e���87h�V3X�e�ct[�V�Tqiٚ�^�.(�I�1�V흲2�eJ��L�P�+J�����M�ܫI����r�x`ʑ�l&��wf�*9f.͚�L9�aq��#�����&��M����+1�e�ps\c� �i�(�b��Gf�V��Ρm���v���56��6�)&^����X�gE��Z&���i�f�ݫ�j�X��X��Єͽ��C665�`�,X�؁�͖5ҭ��Q����]!������m�tI��n	c��pM
m(`�R	w=�h�M4\��&��l#�ɝ6%õ��*��U��#4[�L�ZL������P�[��U�e�J,t�T���-�V�x��
�B�ɹ]��tI������.��4�JЃu�m�G�4��W�R�11�na`��%h]b��.��#�-Ir��ne�5�0(��2�W�G^�%cq�[��rb�j۠���R&Q�&��a�j�fҙ"؎s��iV�JLm�@Ƹ]�)+��5b���2�jHi����m
�mX1Vd��	m���1���u��#�,�j+L��b�1�d�bѱ��MQ�6.\Jiv����GA�)]���-.�-���:����"c���lm5!f��F���4yM5�4��l�	1��l��R�X뚒B1e¤cq%j逩��*6��Sns,۶͚
�h쐘�5�͸.�v����as]�{h[�[2!���j��e�9�\�mi�icT�E��h� �f��Ĥ��e�Fk3������LV]�0gLi���Dʮ�\i��-n[�p�`�i[֑�u�[c�]Q�l��uI����ĹW ��kw�m�Ƕ�Mj&�l@���j��L3,ue�е�,�1��)t���B3lӈ�k5+�X9D;M��s^
�J��a����4�r,ׂ��(gR���y�8�ٍqJC�uGvt�4�#)F�YM��.DJ.��δ�.���.��Fr��i�6�r��Kl�G3��vs��SQ@�su����v�F�$�U�ٛ[D!�Қ<A���M+0�&F����Y6ԥK��P
��TҎ�b��5�.��J�T��lR�b�뭺��hhYq�,����U��q���K@�7-��.�Z����K-�4�&1��l��ٍͥUy�[�%5��a:F�V+�ɦe�!f�(�3n�B#�3Li�4ɋ�����#��t�GC5��퉃KJ�C@3������z.A5�ɍj�*.K��� �S^r�X�P���F�]6\�b.ج\b�󩌌nȎnЄcZ@JVhɇ��MFt`e��*�`�ˎE��<�ɓ!m�F\���q���Y�e\Y���l2l󒩍��%m�I��lKV�n]^��Q�1+M��b�l`�ȅ�����K;;Va�,�B����LG9{d�,k�ю��.E���!���l�Fչ��z�*�i�b�܌�fm�[f(Xsee�ͦâ͙p0����6��՛2�h�#,n�ĕ!h��b\�L������7Q�&�]U1X�e�h�u�:h,v�&i��Z=,a�#���p�,�ڷLR*hLFk[�cK�\=l�vy�M��V�(Y�֢p�[l��A��´�CZg���*iR6qL�u7R��U��dҦX�lI�ks���Ґ�!Ml�%��a�\6�$60��)+���ؐFu��{6`�j4�7@������!��WP��cl�Hh�f�5X�J�J��2�i�j�Ibj;u+tt�U*�J�qeH�/b�Z���{,�%�a�j��0l��-�WF[B��݅W�c��f�.��3�pa{����⑁��v̓�K`CDf�94��W)f����Eש���X�C �je��`ř!�,�l��+�ݎ]6D��v�iEv,�\:%9f�K�Ncs��lhl
hM��ku6]��&������Ͷ]��;L�Wj6��Ҫ	��5�6��6�P)�B*��S*����h8WL�:��Qk�fjS'R� �8qu,֠nuL&�8�ĺj��PɍSL�d�L��i���L�lؕ�5]N��k��9�f&�v%����&nvtYB�6ёu�멭nL����c�/e��˶��A˨�:�X�[�k�L�щf6�q.�@j�jcS�l8��b֛k!`�ci���V1�[��6,!�W$�S�`���4l Qd�� ��3Al����	e��v�9�sT��Y�l��b8�6�dH)�T*i4d����kbu6,���&I��5�-�qtم�	l�ɓn�
����!u.`ф�j3X���+Z%�i
-�D�d5�Ih�ƪ�X'V���Ms���r4�M`$�d��d�n���U�-�[��
���#4�s4Ѳ���L�H���:��� h�#i6�Y�)+R�o9)��kK�a#�@�ZZ�Ʊ�&r������WH��Un�� K���б�eH+�n��k4+�(V�9��i��5�1�h$Y�.ҕ�;�K�"ۑ� ��9�)/&��(�V�:"R�a��7L��/)�E6ɦ+cFV�J\2�뉆�JJF�e���4����](�3Rjڅ�`�e��aV��2���-���&{q��ƛ:�BP�k�V�k�^5��j9��d�h�pi���V�):#س!	����R��Jؠ���i��ʘțq�1�M@�Jb��w-Kt(�ݖ�5�j�qf�����^ GmQn��,����\<�B=�!��0�fEhm��ʹAu�i,כ�j��5�8X�+]-�tp^k)���&���X��̈́ �`��`���͚fRb�IR��n5��Y�wW�A%h�`	YL[��S6u��8�1Sk���f �i��ͮ8څ3��3�Z�bd�$RcX�:��f�.j9Y����.�V:`.���|�p��[����ū{B�`4�	+���he
�5�X]W�ܦbE�P5*B�ZL.t���׉���x�QE5TL�{��Z�4Q��"��j�T���ŋZ�h�s�D�Q=�:zq���t�]i���"�%J(�Ѵ�EJ�Q�Q��V1V���#/%�2rrrkh�Wt���V%�TQ�[*J��UPb[bDEE������̙yf�'''�"�E�J��R̵`�ي�QLJ6�T+Eb!���v�X��ITJ�B�*>�,���rkk�1-j�+V"�a[i*TX/�8ⱏ���*1����;5AQUu����FY�s����K^�kb�n.5`�."�2R�e\��b�+,.+rD)ID\z`��
_�Sb���L�sڞO'�[{j[㘠#h���2�1D�j�.-*#�F�%��p�$ZPc%FIxZ��N�#�n%��JS"c+�F���K,��y<�۶���Lm��3-(�ff�xf(�� ��W!B�J-���y�W�-�1	������N���m�5h[$��me�R�O#,��ry;so2��6���c�A֌�V�Hd�.7l�6P���HF�K�z��r"�W24�X�҉�-q%G �DDJ
��(؍�����5�e ޘ��e�XNҔ0C�H��*�2�!$�������m��m��$t3Yt�U�ˋr;MQQ�nF"�kYv1X�.�ҁ�M�%c���j���F��L�h�k�ӱ����&�E�W7+L�5������ƍ���aw -����ƥ٩�m��&�^�hh�	�6��MZ�ͮ�uK�CUb�Ys*k��ԶVb+)b�,�gq��0�PR��޷�rjCk4c^�]��\+M���
��6^[���
��v���X��L�E�t��+,%�.�L��F�-�	C]��[����b9�"[�K��i�rm�e�;�-��y�����Q��Ak���B�.�F�&���`�s�����Xx�W2]H���	��؈�fv.�p��nK��δҒ�tj�t���	��)C�++e�Lҁ,uf�6�l�e���Kf^��P��۳5uԊs6ғP�m�G6�$5u�ƏW=��D,v�X�Wk`�hu4'6�lT�-��2^��A�����`b��U�U�H��"b�$���-eIc���Dk@#A;Z��&`v�]e�b�(�qn�B��]V�ZMdY�C4�6e,�`�e������jm�d�J-�:���&ԕ������ڕ��4�Ө�.�R�[3ss���S[K-��. -��-�"T���*�;Q�&)�2��f�҅�ձ���<�lݥX6����H�f�&�r9��\���HY�]�uB.�$%�L��5U���7T�\���!��Z��4lMe(W:k���P����]�*�.hQ��	j�BeĻLX��':�6e�����-��F7P�2��K[&�(�R�j4��^�]����ۂ��1�]��Qƅ!cZm������JV�
�5\���خ�m�8Y�P"(1�ٍ�fD����B����eL����3�w>y�%��8�[Q9
uN9�Kh�(^R�K^,��
�����Jui�\*#��2�U���j��Ty��:�`R�V�)-V+x�B��ضX���0y�ԉ-�-���ehȥ����kЍ�d:���^"DF���B�4Ak�A��E=X<������,$������^>�=��'�1%���S�ϒ�ƺq ��p�rΝw�ڦ��ځh�^�賄�;��i��3�8ΛN]�a��	9Q ���9KFD�Q�w�}�q&�h�(������ ���\!~H��v̭��{�M>\Ć�}0c���Lˆ46)�ىF�1�b"� A� ��O���NV��a�Z�`$g�]<@��]���;�jS\6�>"=Y�<�н��b=h'�SQ�zv�$���+�X���Ԝ�Ǽ�;�[%�>T�ѹ���n�@��+y�͸p��+��V$�m��mjnl�����]fw������_���`��o&xz�h���G��L�}�����w�`�� 4Ș���I�6�31ѫTbd�ЌB����E��n2��X܅�7��)i+uy^jdf)YB�FS/q�4cK`֙�*�ٛt��>�$	OUd�@;z�c��^m����N��>���9��$A�o�N5B%���1��	|�	A��q���>i����V�r��\3;'vA�' �M��4��qbY�E�x����� �0��iݽ�����[Ĉ�y0	�w+��� ���n'��R�f��5����nˇIvv_3�?.?,�;���Ԛ�١b��(�#����������v�bRR�߾�}��s���'�_�a��7�y"wv`T��m�q�f؛��{"	ڷ@�4��dS�g�S�. ���Yo��VƘ@��`���|���1ь��l
b˻��dAvt`/6l$�m�|g���;���~�rw��R�j#8_{N�+��GK��ty`���{|l��j���3��e3j��6��b�B���OV��%��5 �����#vb6�@kI�0d�(�wO�fv���v�ނ0&�� Cm>��x��CZ�8'ϹF3������L���>�/Ф+��K���??��؏@$��Lm;�5�&gE3Q6�(�X*@�cl3���1�[J����ᛳ�F,�؍�w��8%f�ˏ8$̘k�'�}0y�b�LG�����B ���?$�e����L�B/Ќ��y���*�����a$N^KǈА����`����=���� u�̤Ax���A�و ��l��o�;>1�#��gjI�. ُ��$ʩ���?�]�:�dFjɂ�W�j"`@-�f��NV���8m���
�0�dE乙~��m�<W�>�9�sX�P޵'L��n�р=��:&/�?�v��o�y;{1�H{��A��@���a�&p�����nm�>;㻬 �����u��QdL6�@$�5[������l3��^f�����/p�˻��5���z��\҃�#{��M,�{�j45���Y��ً&NK��$��m"<r���M��c�������@�̠ A>;��I%�`�d�ùg��yp�$�e��r�^�3K��'ĵ�@o@S�6�0��s�y~�,�ui�+�A��ɲ�)�L�??�G��ߞ_�Q�f���?3f���|ӹ �}�nx��X]3'wL�xGoh+�^yĕ�� �o#�@��'v�K=�P����zӜ�Xe�H�SB���LɃl�?;��o,m�a��ӹl�ݗ�N^���pY��p7��{���YV-���q���l-YF�IK��Y(�bϢ������32�)�fw�m��VY�����<I=K|�}zn��Ҥr�,��`D�'��:&�ԁM1h6Z�]�1��)adك��iN���O<��Ͱ�Z,��p���PsI\��[�C15I�4V�����(�.��L��1d`�����l�V7k�;����k+��Y���sp7f�]лV-%�q�
�@��:�{�)FdMhu�*"H�Hj��u���nk�7teMk7U*Z�j���.p��f��#��饳M����XT4�ִZ�jlv��-nvH�*�`nI�0d�(�׮�"H^^[���7��x�1/I�K6l������ٰ�m�/��]p9O�F����.m�脕�/\@�$����� �dj�u����Q#@e6���$lˇ���0C/6��d6�4�y��n�������s-�9�!<vt�v\A���Ni]^��0q�I� fTD[sa�H�Z��M�>���蠘{��Z-��8��?o��H+�w�%=���e�^7��7�������f'LM�p�cl�! W�0�ᦂ��lɡh��Rذsm�]�)��:�Bm�e+o
r����ت�H$���O�f��T���:T�X��H���@�ʉ@{/��-��Ye	�m��|/��W��?v>IoLWf5F�G���\�:PLG�b��jjU�	����U&v)D�U��Z����@S�q�T�d�*����&�x�M�DA>$6wG��,��Kq,�I��`$g�r�e�N���1d�d��5��l�?���0��׫ixH$�T@�Fy/;n��	�lU��p���-�Z=M��Ĝ׸h�$�y<g�Vۃ�;Q�$��D��7������sc�m���@����z?�C���.�v�c�y؜�؀I-5qP���48�����7���h��R���aD���6F,�K�ai&hk-b氏0&�L_扼�����;�g(3�x�d��k�x� ��/���`��NS���Γ�O����/�F2��������I��r����m'��$�j�9��V�?=�X7��"�$L�sd����M�pH7��I�� ޚ
��^f�Z3b�*��З�����e�X�:�3����4*Ⱥµ��3UZ|ƪ���B�U���yѱ�ʤdPNC�z��\���3����>>
����&,�0�5���N�;m~�!��a����8o?�$�����ښt,H&���
<N{ b�L���	j��D��̈́u�f���D�5bЎV�r|O��ßX1=�1(Ϟ70���\&���eH��7X��&na���vM5ȑ�}����S4�sbi�Y0ĐV�s7����D����*�5`=�ZG��$F�8�G��1���vwd�Pg�7[0���W������4iG�T<�[��+��~�{'ܽ��3h�<��>���F2���r�@F�� R{U�$wn�Hw"�y�ͮ$[['v,S��1�"*vN�&6"�qx���l	&��#���w�MS1�4K̦��`�1Ązp, ND`Ŏ������ꭅ_xl�ps�܃�Yk�{�S��J�mZ�И/\�F=�4���3�y�����k
����� ��ߤg��ʞ���K��v�"�$���S��@�������\%c��L��	M
&�����b��,a��-����Y���|5��h�dÇ+�<r��	>'��u��|��Ř��0Z�k[� ��Fu���iw)��4�9���3�w�q����l���O�3�����	 ��75����I��|��C8�a&'/����n@����/":�ʶ������̦i�D5��|׀	�Q ��iNY�����m���nDn�&w��f �A&����Hݷ1*E�ɧ�x�@#�a¼�+�Ye�D�f1�~?�����j��̟�/�,�~� ���״����n4���_bj�/�y�4dxfm��}�Gѕ�����9���~y�R�v�Oy��W�+�<�sg�"j{:��4���%��|��Y��-r�ǩ+%|�.�	tk4�W+Yk,X�������!YJ�v��95�k\Ct��,ڔ�-٠��n��u�-��U͊�͡f�sb����Xꮠ��h3[�W�!\�F�C�X15�`#M�v�-)v��]p�<0�� t��V�E#S55�Lܘ��aoZB(��Dt�=.�e].�Ƙ��J��tt]QҦ�-� ����Vͧ/6ٴH�R"�gP�#InZ��:{��{��W:\������x@�����%��p�1��z/i�����)�u@6<�`e�EÄΐi�W���Òy#�gKLdMߠH�m�HݷB����w��~�<Os�?��U2^�q�/���bEn��h��6$�檁 �v�PH's�<���	�������6Ȃίa��}��Đ1�5�����g�o�xF�FDNRt
.S;��_�KyU۽m=����ds�U6ڂN�0�_��A �@�0Ld'��	)/9xL����@��l�#qBj�sm��L��K4��5�L��k3��ӧ1��)���o2l`��^rb�a�)ٞbm��m!@�k9靃1,�ط�snKe+ň<K?j��̥�OW��;�� ��Z֪/&We��}@��Ē�_z�����+zR��eחc��Y�9W//��>� �[$�ܘ�Y�?p�π�~���	ŵ5�� �lǠ�H&���t�Գ�m[��$���n�)U�l�N8gr�4�ҟS9l����$�g`�,$H�؈��}{5xl�%R.^�`�w������vr�9``d��H2��stlj���yN'.��#<P$c�����|?~�J[o	���ݢ�ј���K`6��u��V��ue5�3m���_��u-l)vL�v6�9�k�$�}m �Ų�!��2=yn�A��x��^3;1��9�/r������i��;�ǊW�3�|}"�%XzWRq�dI!��nq�;bY�h����~9�d�|<|<<=��0~]��^>��yv���eJR�r��t��6���k��f{�x^����9emg��S��;�XP���y���Ot�gG��n��t�y�H�I����D^�y(��U���޽ {sm���LӼ�	�dg�y �t.�o�
��~����.�@q#5 C˳�g{'�N��f�����ш�sS_y�����4���Խ��8P���2�,N��{4�:���i�@�B�dXlLr�B"�0oK�ML���Hyn�������������N���Kww�r���iBo}����j8���<;��JK�����5��x��v���>������:N�g�p{�\ɛ���:��H�;7;K�����7.ޫ��D��.���_Թ�ׁ;E�oh�捣H��}�������8�x�z�����!�M�=ƁH����C~'�P��N[���x�wc��:w{�<�d�"�O�=���/����Ȥ������zk��i��f�xy�LE�d��}r�����q��iY�k�W���}���Ǽ�Z�n��p|�nv�Jߩ�/|����������f4{}^�{ۆ\�������:��b�վ�\�X��@@��hո<�=��n��"3�O=�gl�7ܼ��� m�`^�̳Ш��3
�.;�Q��;;7�ށ#%<�����|�mּ!���q%z�/G2�6����,]g�*j˫�7&�P!^c�QB����.���h��DƉ���.&̴f,S0��Aqcr��\�ǭ����V�u'T�Q��;v�]�;75��A+F�*(�cU0j5qb��[M6Q�.	�`�bRV�Kc W�e>��۵9<�� p1�8c-m.5�1)�̭T��F����V3\A���[s%L�2��gc,������Ȏ�x���%h���˦�Q*�j#46�
n�"�J[KJ���*�KZ(#�e�5=��ӵP�m�%�R��%j��akc�ph��A�K�[mj���h2ҾFY������*�7�%��QrʉhҢ�IiT��
,ER�҈]�T+S��jvnvf�{aV*�[B�7�1mh�����d���)Yb�����,EP��̞NO&�[���Q9�L��1-�PP(�ed�\n[-*D`��2୺�,���٭����-��;)C-Qb�eє�*����D�/Z[�(�!\pU��ī�EA���5+iSl̲ѵ"��,�Tm+R�R��J�֡P��q�O#�y�R
C��d-���g��Y�Ow�p�bAN��w�z���L4��u:�3O�o��_�V[���}��*s~g�pd�d�������J��+���3��w��=�o���h����o�O8���S_{�06�s��_���ki5��,?gu���n0̲�»]���4��+7ug<����{O���,�9��ND8�c�j����풰5��w����q%a�V=]	t<O(��&f�	K:�>���@֍�L���f����V��Tl&�Q��S���t�����y��3&p��x<H���"+y�0�%g��L*o�~��3%d��{�)�a�a�w�}�y�� �����Ado�{�T�(s�|�~��]-u������}�,��VT
���^�9�Bm>����N!Y+
���������d}���ZS#��;V�~��f?�e���G�g�A��G�xPX���̝����F���5�Ã�c�)����C��5��HVz#I��%O~���ѭ�����0+*a����E2T(�Xư>���a�������5�5�b�I9T�}�����5'���,>�os��A�
C�{�)��Y->��q����~���������/.��9��,�!��B:��L��ݥ�n��֯7s�vK����ɛ$[��3�X��M	��6��;���H��B�������r]z����])����� w��m��$S�ﳌ���������{��N��{�M�Q�Dg���m�(F f�I��=�b��ܜxt�E�zژ'���ʜM)�=e���E[^b^�`5���D���%*_bbYػ��}���ŏ�>�G��Yl��￳Hn$+ �`T����|� �}y�Z��18��� 9��ȡ�lH�Y*I���m�P<�ן�~3.h�i�k��OF?��:��'+'�}�����郎>�y�Ό��2bc�a=���Cq�%�)�����W�	^#���e>¸��@Q��<H��5?��}i��Z�f^��C�٦{�Y�ȧ�߳�:��.��bJå��{��Xg���I��IcL˞<��^��qJQ��;N���R�8_��3Y��<��:8�٬�𭚧iQ���$���������gw��c�!R�
���v��p`VT
�&�����(o�����g�~��q��5$�}Ͱ��0�����ff������N0��o}��É51��o�؏H#��L��r:�jX~��%HS﹭�6ԅk!e��������V�5���l� ���ϻ��.������D�f)���=Z��4n�>����!�=1j>�_rػ�цw����-���Mc���
�}a^]:g"V"O��F�j1��|/�l�Yq݊\����������ew�ک�(�b�&��,]�ZmY1���X�2�-�XĻb�2��e-��X�nYA�l4غ���f���(�tr���b��TE�MA�\�g�\ ���R[3s��kEv\�up���#h�t�Ʈ
G�HCk���tR���� ����$!�8�TK�X�=�]u���2���,�a�WjMZ��u�]{j ))P�V&�ȵ�-�3LeKs�z��=���ZƆ4�@����oK6 VT
�)���l��	*1�׿����0�>��w����p�=���g��zY6�d�$f.�� �zkI&��t�K;r�Q�j�'���*ޔ[��P��B�z����.��%d��=��Ag�����l���;c&!��{���ϓnO��<��Ǎ�+,��M3[:Ox!���?{w��8�P�
!Xk����2��C�AH_��<����1޽�Hm�
5��i��;`rr�,��C^��6E�S��G�;ߪ	�r�N̯�A� ����T�j�+�k���Y�����u��P��<���'E�T�������T�cY23�}�,�����~���}<e`Q�O5y�!�8���/\�Vf�Y�y�Aa����Z�,���}�����
�s�S���w�{;)=M0*P׹���G����{�6E��P�?y����IX]}}�}ﾏ{�<_P% C���6�kpl��[��E���V8��ah�`Q�H�}�g��q�O���>ya��o��ta�Ad������8�
�	D�
~���Hm�������7���{s���CV���{`p�$Z0������E�S��w��s��F���n��@�ޖm��F!�~�M}���].���}�n�z9d���̒f�������p`��'���&��{��>��� �$�#�Oc���R�q�S�h�L��t�d�~�
�V�~�z�+� ��eA��oK&Ш�������x:���vOD�	}����WZ0��ZMv�:�߼�����-20*C���/�IAM��3�\��Y�y�\�bD#��^��MF�5;c���v�h;�0�
��~ޖT55�_+�\�u�C<�Q�#�u�6��%��B7��2~�"Û�����ߌL��̳s� q1�R�{�Ԇ�ԑd)i�oݲĞs������A}�
�&���|!
��ʭH&�A;2��:� y��K6 VAB�T����)�m�!�������Dy�\@�#�Qe�p��!�Jy����B�����?>�l��R%4Dq*ᴺ-�2�D��uE&ơ4�f��12��Beɧ���h�[ó����,�ǐ$$�C�v��%w?R�@+��W3-*ݶ)k�h���3�Q������VK$�3���qNI�r��4��FZ!����	����G�I��P@�c=X��������4��f�	Eâ[��vL�G���Iٺ۪�PW�D�7Hk;/�`N����'�=�/�{6_w���÷�1�+�=�L��n$Y:����)ˏk�e��L��o���|���H�o@�E �	o?R�J[늻պK�`���3D��
{���ESc��t$d8�B@$IW=ҙ0�&�����0R����$�O%14��p��3�a]r�>
I@$ٚ�!*��D%b�̿� �z@I>f�S"ew�2^�˦@iJ0oM�T�x19LB,�	&��ɯ�z�h漲�26�f� 6�iq��"h�,�c4(ՐO�}̂`C��-�S���(	V�D��)$M�� 4���n�Ш֗�r٪<��6C�<Q%[]"@����M�%;�;���%vL�I *��'͸����9��J�W�ϒK�e���~���Xݜ����د�3��霢賉y�O�p�vf$gD�Aw���:�U0Q�8�P�	ԍUl	���E�z@��K��Ʊ��\:,�v�/P�szM�Y��2H ����E��bRI#]�:����HAkTQi��cN�3<J�Λ�S��Ծ
����˷^F}�j��~�������������%8ё���;�x�	 ��L��F.�]�	س���A��@�)$k�8�]�!{�fl�$�;dNz�̂H{ɉ@+�L�@�	�M�mS<�]�Y2�
9tй��nU��j@Z�Ml��e�:-�ҭڮ4��8vA �8�9��D3�wA�	u��e�H6n�����|�����H�L�@cª�	G8��}U"eP-}��{"��"�E,�1��!$��eѫE���������-�291��2��D"�T{-0�|���R���PV˜��vgawix�fD�RH��p���
"��#������}8g��~ȉ		��!!�~�S��tΐtY��H��׼�ʧ�����������I%w� `${�`jwfYƷmK����"RB�φ֝�N �aGL�C�f��D8����jmPIx�wLJG��w@�E ���|&U���a�
���ۿ�lh�6ѻ]6��k~�`�{7x��W]�����$�`��F;2�9�"���в��՞�6I��ѹyc�a "PP������,=
l
���st3�a6!�Be��]���r���
WKi�ݥ���
b�V�Zj���Q��0�r ��
�Q��h�(��cn��e!��.
\��6�x�Wr,�G��.�.��u.����B���٥���.f(j݊�a�hv6���Y�����C�u���{uE63)T[�usCVS�X#����f�LD�Z5�-�f%a3s�4�+�hU��1s�����)e�O��-�fD�~L���}q�f"W���L������3�ys1!$��� C�'���p��3�ZU�� �K�kM�$���I$�
�Dy$�K�z�D�D��Tn䠶�����IlKc � �(��}"D%�A)��!$�em�8-�碌�N��+�e��ɼ ���dO�-�p����x�;'av�����U�E�d��U���. BA%�f֭�L���M�Z����1\���� Dm�IA��b� d`	GEę^�Ğ������;�Ԓ��$�����(��:����VM���k��k��.� Y��yÄ��2]Pp��I�����w+G�s
&ڡ�cT!c�~�=�gЋ�����q��I ��bA��Ȭu�K�����C��U1=�JUur �:q�àS�9����z�C�雟{U2��X,]���*�-�<�����^˕�V]�$*�/DT�u�{��d��N����U�o��)vА�f�K��S�O#��.m�zO�$x���8s�"Vul��� ĵ{a���$g�1���,���6A�'B!�3��$��f�lK��	`L9�[:���e��A$��$A�)�yن	n��B柃 ��������M[+��=AE��d��MWp&<d���E�Cf/I>�R�F��W1by��tC�;#X�IyC�H�%�$*�gogd�&i\�ٗHy"s��eڳ��T��"�B�zD�I$����|�y�̂��G�?�����g����˫�-�F��v����ҕu����M��m �\��ds�����E��F�%pvᄩ�310�v � � �I^����Gs0�;�ж~��}>�E$�u�J���4p���E��v\�>�C
5�{��ò���y�5y��F� �y���-��l�7r4�)���HL��;���1��9�d2A%��@p!
[椵v�6�Ɇ�����_U��ӳ�;����]����儉���5�Xn�������$���{a�3VH�4Sgo��f�π�O{	��k��R�0f [����r��3�PK�z��&��}��&�`	HJ��L$�i�ʲ`ez�|����R�}�q��`�tC��)Ul �37����o)Y�{������>J�Q>EO�_@�7�4��$H�fr��E��.X������X`���C���;Z
[�\��C���A���>�����읅p����W��-�q�I$�t��L��V�g29UWg�$���1���y�#	�O/�K���YE_&^n�z���OI������kƄ�H��!$o����șE//(�jSO�Z虧3:d$_E-l�.0v���f	 K�z$�),�kq&����H+ހ��QI%�;"@��ղ����$�_�j�=�ι�(�ݴ��$�Y�� �H?��v2D�I,~�E`z�,Ի��EU,���멂6E*͎���v{;��xdx�����{�9��{��{|�V�:�}��Y������_v=��Og�����,X�b1 �x%>O,�!s��<�!����W��"L�A,|�Kxյ�M�L�g;S���I�A G�AfLY�E$�7�L�~>{�<>�='�6�>�ff�������PJ<��:�Pe ���QHjM]�Y����sY�F�*���@sIy+期4��A��&<�����iئ��=��L��^M�H.w�S(�$c[�r;��*�����BH(�ʼő��_:]�BH�C���(���)$yzz��\�<Dz���I�I�'<\��,��<��4sEϚRI#�~؉�bI����ͫi�n����`�o\��'�ɒ��x�L�Q�����';EW�L��S��cd�ljI&������k�<&B������L��t�r&d��ͨ2&�(��p�c ��\I8'79��V�]��K��P!g�1&Fy�<�� 7:xD���,��xx��,�3������L�p:���z�@�E�|�����
�4+�\&hK��,�`G�{:��u��s*��л_>߇ްt�u{7_`q*XX��H������\vx���UW{�����Ҝpn�.�N{=��Ra�,���5^e�c�0���85���;f�w;����@���9hRvq�R:��,���>[D�=�[R�}|���}�nߡ��C�wt��v.�x/v�>��o�JG��y�sگ�{�?o@��񋼼���Obw��dˎY�wͯ;dɺL�+�� �;��i�nr|x���pR�v�3�t�V���k۝�p0�q`W,�}}�-[f��iݖ��:���F��3�b(��Y�gy��b���d�Vi̇<;(q`�;�6o�nF����*I�� k�~gW�[��v��4�����]}�Ŭ���c�<2p��Վo��89��׽����|��}\��=�n��(�-���}�N~�����ޞiV�S���H8�A�-y��sKY��Bk���`�D����;�s�Oz{��첖���T*��©�R�E��[�X&�{}�ٳ�����w/c����w|{�U��\���/���}�<s	����S7��;���2<�Ūv�ksʐ9����%,]��y�C�ۖ�*��>�Ե�\�b>���[�ۛ!���
�����6�,�G�s� �f0���!��	 {OeYF+S{1@�PVf��1� �����RQǔ�g�?�I�������O�2d����0<x��/ʟ��g�ו��(޸{{[�����3�������B謥�-�4�>��(�f!2� �6WA��9Rs�4�s��)*T��y�L���O�����*T��DQm�DVE���2�b9E�)�+P�E�¨��Xde�=����m��+��eĨ���TZ�I�L�1*�*6ܲ��Rq&���"�Bp�8���x�����I�*���3��XbUJ5��؇�;�B�Kh1�uKZ.��d�n{3f���r�33
���m��2�e�TX�R�s-%���L��Ј���2�Og�ٳ{��L0d�LpG(z���
�-(�f��*(�eq*��TH��d���&� ��EwlUcW,��r��Ѵ�`�1̥�_D�aR,�ܳ&�'fjowE
YLJ�Um��85��U��+�Vf4�,Re�VV)�e�5;;5�v�(�Ѓf�qE��fdM.�un:`��[6���K2jvvf�F+��)�
��J0VȤnb+Z�.e*�Ce�ec�F�-�1�U�Eb&8�s&
�2�R(�$U-���:�n�[��s.�nk~:1�a�N����U�fPЕ��)fd�e�$y���˦ZD�ƶ�V;.��3��+-�`�rl�gF�Ucu ��XG�q]�\�50��8.!Y�-�rJ�&[�j34�ls.��e0�JX B���kG [�K
�]b���F:���l0�Z֍���,P[F:�uΘ�8�L��W�Ò�FZ�%�m5r�,7<�sKZ�%�YR��l]
2�,�9z�R8f�f�ˠ�ėM0��n��J�3gv���&ua�4��F)c�n�/P�1�BiZ�����	�5-�u�&�I^c)�T��Mִ�ŉ��m�d�iq0LT�S.���G35,��k��jE��ͷ�7bͶ�S �@ڴ�c,�+tI�l��B0s�@fĕ�XQ�aj�T�ű��\�[�ь-&G�컝����XH��!F���m,t�壇Rm`��M5uf1Z\PNՆ�4q�fP�aq֓6�\���j�+Af]]]�L���\��:\XK�V;]E���ō��M(���7�r�ͥt9��%�3���ԡ�Ye��5�����Fa���k�,z�[(L��,�i�ҍ
�؆0[25�2*),��FmMe��
K(��Ul2��-��D䢐�+��jݗA%e�r$�8.���[c�ל�K����q9!�j�K!��ː)Q�Z�K5���ǆ����H�u��.���T� L,!iλ)��XY�4dn!.4��Ý��\¸i�lH�L�f��),�^��a٬�d���Lܭ���`�۲F�������2��V.iM���^�.�7���K�R�r���	R�ZB�+Gk�:����%�3j͆ǌ�6�jF��aM%��s��Y�Dvu�ѱJB2�+2��&\e��tp%V��)�F��*�ZӶ�j��ą�α�P��n��3��I9f`�]��]����e���ĳ2�.(0s�L��uڮ��cQ���k��!M����\0\ۜKVi�����l������-��g<����z���ۦ,����j��&�8Mm�V�¬b6RR��q��d-$3����ĉ@�u	���B��RM3�PVP�m����<l�p!��T���-[��s)3�e彜ʁ��L�43����;b�f &��f��Q��g��J������>s� >Iu��������6��5�ʟ	E�R�݉2�<�A���	���:B$���?[��6m��y$���=�FG�K�6��W��e�7p����_Dz3;�A��Iܠu��yػ��30�}+�������K� �h�(�c����I�o�e%����)`�Q�'<Qww��9-ʹ�J�B�νp��A.���! �I́�H�4�3K�v�<.�/����$�)`fI8`��*�L��K���i�i�o�q��u҆��3^7ʃ"J� ?�� W�;�:�S`��'�2fE�������;�Ԙc�[1�H��癋�\3+)�T�LVz����b"���@�14�o�H��q��	%�ӷ�	I�3nʃ�{ԣ���Iy ���`bkۨ�Cgr�3�W4�T����G�r�)���ܤ��ݯ����)h���Q�ԥ��y`ѽ	]�<;<=x�K���y�_xo2��;�|@�1�|g~�����c��@�	$�]�͠ �D��]��m-=��ę�<�A���:	�T��z@	�]�8�RA(Ǯ���q�_c�y%��ٛ""��y�v�x�2�t���7�˺tª�{�y�6�w.���ٌH$丄���@^<ڙ]�E��z@f�=�^�=��Ѱ B]�O�#|Qgwr�����n�'��n���_)�=�~g�n�%��I f�9L��Z� 4���w�a�ő,h!9��vL�q��S �j��ǩ����i��S9�|���3�'0v�7�ؘ��h���3$�OKJKwj�ϑW:=�b�\H�@^I �1H��''�(�1��WL�@$�MDFw8�HW����e@I2���,I �L��Uҍ�<�Y�>h�Bp��JD0vw!�f�[m;>iI�	��d�؟:A$�{�j��Sl"+�6��ѽ�\u�:��A���iC��V>��a�[����D��w:-��z��xy�;���滼����1�e��F21��Nsݛ�-P�����xq^��不��{'�S �	w,AOF���.�ml6[���@)v��҂I,u�!"K{ $��<�	x�<>O�F �A��cwJ8��ɂ31C���I"@�a����mFݒ�cͩ��`�It6d���Iwd/��ߺO��O@P)eeͮMMtD����4[q,�(#�&e���5#��'���~u+�r�렏w��k��W�n�tI+{ @�P��,m��7=R�E���4� �i �vk0�̒p���f��������.�U;cUpi^H�P�l�iK|�ˁ�"aG�2ֺM&�b�q��!P�����+<��5@ ��ں$:I���W��$&p���c{�	Я���f�i�iI$�[� �Ȃ|`l�Ȇvw!���>F��Э[m��<�ɱvD�@/$�U�!$��=����
�Q�
y۷�K2�DҶ�4'Fj�qfY�?��w�Ι/�.�o��S]����32��N��pm	�k����|=���fd&a�&W�AwMkA��o�i	!�4��f�� ��*~�c���� CСF�	,^�m�<�U�`��"^I�"efX힇��0�&I�����jJ�ef��[��F�s+�	�v�^N���h���?���� ���˺!������	$@(uFșIV��M&Y���M>H^>@_c�1<+�N�ӆl�ۤ���}(��'�o[������~�>rH��q���fd�g��"P%m�z�.ݍi��a��$�h��/�@$�\tH2�@γF&8{�2����&}䏑����]Ѳ&Wz��+|��3J�WH�4�z��{5�Jn�D$I.���(c���ft�@��j�����؈a���.�`��C�U��`	RI,u��WZ�u��0��d�y��@��t��R\�zBMU����G� ��]�F�ݩ��;3��{G�ܾܘr�����*)��,�/`..bG1,>�Y�Z�se��Hv����_Z���|;Y�sP�J��㛍W=s�O6a&RdfP�t8��Gy}_��1Y��UkiQ�%���i�KL����c�ڡc��n-̶�3!rM���+N��mXX0�Aab��e�s��6�
X�Y�+1u2�@�D���Dڕ��-�mV]�U�e{5���5��B5���-5)��.������A#G���٨ZDҝh�����7�(�+(�s�!��Z@R�M)I��G��u���`&��xd���[)���-�hg&��	d�`.�*�{������rA,�~�s`D$�J�2%����f%�zX�J�����[ƍ�ļ��B�&d����	�)���vrP�����d2ISl�&��wF�s==	���ݙ�2y�`����dd$}U&���2T
<�3�O����N��;��J;.JD�g<HIy$�>LiSoD���I ���ky7�(�� ș!�n���0`�atL�P�z���'p�CR�A ���I��	%ݱ���b���<��ݏ	�z�Ry�.�j�m��2&�\@�K*�Xƻ�dßfD�I%��ؒL��[�!T�9j*ֆh�f>Fe��A�Њ�X�-�7j��\p��]F�K`�,BC�顄�s4�D0vw!ߨ�⾹�e��$���>H�{�Á?�W�f�y���{Z�UNH�E$�7"c�G�/X���
�18$3����_t������k;���u4��4�nՕ�M��AC�������1z�v���w�q�k�9�g��#Y�ٮ]E⚍b����k~��޳lS|�Y�0���O��2��(L L��d 7|���.Ks?{�|ym-~��D����clr�ў��ה91��;�tP���+�I��Kw\9��3%%��Gt> 䏕vDI'�3od�	��<S�9p��Ą��ᘴFwV������V���@x)d�H^d��sʃoUH�V���6� HIy�&$�I�z6���0`�"t�K��$I)����^b�;u���zbL�*�3/.Ȁ����IwGH�(��T���J`Y�m�	5�]R�f��C9�&0��up�Xʡ!K�J�1b��F%���Qg1�	�m��H$�8�	y"w��D�1Ū����dݧN�K�yc{!�Ǜ�@��7��"��tCwt���u���	,}�ۭ�˪��	�A^gI݁�|���L�
	���:�Z%ԾIW��D�Y��\�הz{�H,Ky ���|d�� ���p��u혵�a����I�.�*�!����س	�2������D�G7��ӆ�+����a��w]�d!�d��)0)2���ȁ1��w���D��>��	%�}�&S{��&6�p�W�q\�gz�Ph��5��	 ��O8�D�$�;$L�"[7�	����\�yꕩH\�s�b�@���'uQIF]�oD�y ��^%-��jr	ȟZ2/zBD�u9"e{��7�	#!�;��Y\$|W��3x�fg
9mn��R�t��Y��Y\Mp���cś߿�~�r
p����Ңto� IW=e �	 ٽe.z��n�� &2z^I.ɹ�I���!��S'4T��d?��`��*7���~	)��>d��Ća�dY��^�n�$璜՜*:4K4���f�ls��.���w���l��I��I�9�|�H�m�7a�bۉvq�0:R ���mH�IA�z$�>Ez�w<$"Y�C�C?z��W$��-P�e_�%��d�P�30~Ή �I#W�4�o'tT9��KBW=U�E�ꬰ!��枕缷�ۗ^��/�|�D�77�Vؼ�Q����Tsπ͑�Y�Y�Y�����1x�[K�k���P`�Fu�����;��z�dW<���̗��\D-n*��N��l�i���M��&BH$��@�B>1���O�7b(RR�O�I��c�A#��2[��,c�V�T��]Kt(�j�ȩ'����|�c*߾}����r�@($ݺ�>I$�o�<y.�*SEy����Q�[t;A�?�](��(4�U�r$�Y��l+���A��4�V��eQM�f�$��H���2�f�C�wh����J�im�J�o��'d����y��J|�f��K�e#yE6K��ڛI��j�2�	%�� BQ�=��Aû��d�7uE��v��̈́��e��d$��� �	%����#�*N08R��p�z+�$ϒ>O��6( P`K�C�MJw�9��K�%H�{"�W���A��$ϒ%��#Ы��?+��^�E:g5����v	
7�럛�A�w:^Sm�q����l�����+��1�!��?{^t.����C�r{53�q�Za�5ߨ�?.�@m��]aqe�ȨxaD�&QI�R`Pb B��|N7i̺��csm"��U��=u�5Ԁ�Z]-�6d�1	��-�0�dj4-��bb����=�։74�͗JųM��,���E�.]j���bM�.BҩH��,�Ԩ�s��$p�&ۈ�s��w6�Vò����ڽ���&���Ęsv�ZnGj�,�\�k*T�W�5�ff�˨\�bĶ�Եe�.�tˬo]�2ĶCKP�c:���klZ�kB��Ĳ���\] g���f>wt�|_�q |I$�������7�z`̄�f�� ��:Ox�u"W��@�	 ��;ߊvw����]t� )A��أO5��4�^>�Ť������~��̋ �z8̠
J9�Q��,�Ni�[2�~�6Hn��;MXZe�$�W�bR^	5Lw��Ϥ�I$�vB)$�:8̠A��c�̙�`�gɻ���o0�j��H��q @	 �(dlq� $@)��$ة�|;O��=�N-�����Fpt�p��=� �m�=�p��Fu��P�{�W1��X��g��D��w"e?�y�H?wD��j���Q_��Kg�Qi
�5�{MJKM-���=a��j��l5&�0�z���{�0~��1=u��
ٌ�RD���!,;�۬)�����8�K�"�DΠq�3'gA0���q]!$L�v:
��A�R��������^I^ܓ�h�xD��O��N�p>��������j����DUY�C֜.lߍ-SX&����*�2�L"��!0 1	#$���G��b�����/*n���1 �$ޡ��Z7/�"��v�X�K��AI�
�'@)݃β1.ڸ}%o�g|�I�I�ufՕ�S�4	$�����!�z$>In'Q��p�h�]3����2s�H@&{���=@1t�g^	9�fH~��NǶ�x�?�ϝ��D	��2���X�gE� �O<bH$�3^뉅�f��n��($�'�L���� 1 �H-΁��O={�����m�t�V��͸�*vM�n�+�m�f��;v�)mD����}�lb����T�� �$�ؐ�{9ÁI��*f����ꭁ2��K��} 4�m�0H�%�!�L�΁��;�q�v+3"z8w��I$�:zZBH${q�@���xM^����	H*�r���?�0�U'��3��#>H�k�2 �a�<<�3�K�9�u+����aI�wɎw��qyr��ybv����}��7��{�x^�{Uܓ>@�5��쥎{�g��9x��ȼd.wN���O�O{[�Ý�s ����<�ѽ�o.�pv�=����i{^kɎ���:���%��u�H^�����o�F�yf�Y��t�3P�o���'�7/�y�f��v���������4E�U�`��؂м���K��<m��9zt��8T�E��
�{���ሟs���Cw��0��㵗�T�_���j}����gf��c�I��۽�����_?n�ޓ��8g=���'^��-7�=���3�z 0�|�`�q.ߌuN+=lLg}��k��E';����	D��Ѿ򞫶�g�����ב�מ�&R��o�ex�'�yw^����=��T�w��|ݽ�y������q�?uX��y��B����]�,��73��tN��M�L=�wq�����c��A��s�����g��u�wz�k�nS�xz=���ɷ�#O=��K@&.�z/{qo��f��=�l�����êq��,[�;A�@`�k�Z���F��K:%�r��u�{Nx�+���=�qę^𓶠�;�7�-�m����s�|����}p��-�|:�#�f��y��1 v�8� �9�Ƌ�5X*�����NdS����C1<���j ���ў�wq!�/�I�<�L�?��A?�4{ST���EUEkǍ�w��і�7f�T׏sL۫�6�
����`bUE�E�1*q�
�~>y�x�fk[�΂1<�����2�c��f�e/Bn̶�T��,EIV�TƦ0�ԳSS��h�ꬋ��-�B�e�ˋ[,�.�����F&d�ɩ����ބ��n;!�mq�eB�Lb��pĨ��b"�T`��a��y�=�}w�nq��"H^��bXMaZ��[mbV�F�m��1i��SS���jZʊ�6�j��Lq%Ģ�S)C�S-�%+����ZV��ML�����7�+\�Y�k	黖������VZ��̀����'�̚�O'7��@F&R��d`��E��̶,�,�̢ԔG,��f��'&���S1���ִIR��VfS=��iM{��IS�����)�X�e����fh+*�V<J������(R�V�����V�(b�mTvZ��J*���30j�R�V��K���@ܤ�)2(L��%� ��!2�L
�w�Ύ��Z�:߈iH�3|�@G�C�tV�:�9&uqiv��q�x�B�-�]$�]� ��	/$�����$v;c������	��7�-����s��X�E� �څo�3"W��Ή NoEv�&A��>dO�o=ܴ���K˷`D"o�t�G����=~E�S{����$Z��x;0��a��SgB8jny��AJ�k�g��ֲ쇯���9�,�b�Z�d:A*fk�w�I$�譑$���ӹ!<�[��<�l���I%����`]�)r��;�PJ��'�RG�W"�w�0��U1���bk���I%� �a��"e?�y��cN���:�7��Ms_�M�$����^�^�5�H^IbR\��"BH%��^<�y��>��A^��W�=�&P������?�0�-J:&�R��Ѳ�	g[�0�o0â�wƩ"WCGKw��Q����v�]��O� ]� $w�ۅ�G���t��i.���Y�ƀ!�e�����5V�ui�}�{��� $��0�L��(��*I1 H:��/￶jlk<<��:g!΢%/��'�W���������^�}�ͮ8H..B�32J�6E������ 4��P��WG���);�64�܁�`��3L5��7��3̭X��E�K�����R��X/c�p�nn!�I��wt�:b@P@"P�m�i	��ݲ�e��P#Њ	 �Et���2���Y�gfI�ז��t�X�i?��x��q H$�z<����$�K�o@)$�F��kx��2	:Eo�.��{�J�z$�y��@-���y"e���bS��H�U�$J),u�!$�]�N�.��s�\�KhYND�PI%u��I\��(�d s�&����I(���T�ކ>I��U'�jiz]�	ٮ"T�0�"�@r���^��Q*!�nYH$�oQ��S�@.΁��K�{�h��2��SI3'��}�~�Wj|���w�O�7ȫ~C����/~��)���<&v��}鐣�,h�=��a�idX�g�$����/�<�l�l���+���l�3 $0*L0 c$��۾\�G�����԰x����î֢U��V�[��7B��Z�-��6�Y�~x�ȅ�<ұ�aZgn���.�J��%��'^ʋ��G%p�կK%���.fή��ً�%����[��F5�L*�Ս��t�ّ*�,Ёv�8�(M�RWkֳ&8�F�d,�˙�B棊��.��u�Ն��
����jB�
�V�C^�	tn�:f�*�1�5hl\�3c�əؤ��p_ 霄�;}��j�A�A-|m��H$�:B�6;[Y۷��v�ȑ(�
쎎�A �t"�`�"it���Q�&��wb F ��̭����H-΁�I�kgc���n{��*tA]�.5�2��1�X���H$���	$N�0��h��~�"A��eJW��˟�@���Wy�t��w����?s�A�N(=q��I �i�%�H$�IV���	$Gt���cx�-y0e��Ф$��W\$���J��z@	 �	d^@��+\�firUu�� $���b�A~�g�3=-5_{���H 5}�V+�rZ;l����F�*���J��-&�&�rKq�67�S�/��o�3�<��!$A.�p�<|�@$6;�L��3�T�TI�f`�@m�1��V 霄�;L�5-&��x�?�����Z��W��E���Զ҇�L�#Ф�j��r��ƹ15�w����}6�~�/z)��;wM�}2�t��e�g�s��5��4!�f0=gXCi&����&�4���� U�Q��� &	�Y�m�x�$� !��"H$���H�Q�̝�KV!��lϲW_I�ɰǂ,���4�fz)*�����`�,m6NG=�k2H�vE"z+�A�ؒ��r̉wI�Ѷ��޸��_>?<�O��楤�)n��c*KJi_�v� �հ9R�[e=%�LVܕs
߿Z��|ѱyǩQ�2	,�����o^K�h�{*����2�	�g�'N��y�J�:/ԩ$LgKĥY�@�O���p�HI-e�{	��~��2ٚ7����T)���o�ܒ�������W8����)���Ě���J��翟FZ�i��O={c!���̉RD���O�os:���5��P>@�D��t��Ǚ�\hF�1��.�����)>��Hpj�)�H$���K�2M��BH%�u��9K�� ?����� 霂�;LO�ܻ�2���O���y���������G��zO��A�S��n䬎���b�5���u�Gg����:L��E���'����{��v͉�5ٯC[����D<2�L*̀
2�A� �# y��Ŷ�}��D� ����$�S�GC�wdX;P��"z�oK>�0�V���f�h��ܯg��?��� ��! ��;`�z/`�f�1����g4�Y���I��1�K�u��3:]����-�ه�$����RC|���$ϒA%坐l��w�����2��UQ�R����ي�f�D���h��{^Nmq�sl�,�-{���`�:gt��W�Z��+�$�l�x��fd��3�	O=��ݦ�֥�Z��֙E$�x�I�޸��. �����O8�@	�6����4Q�9�n�RI$3�L��X��|���PK*�q�W�ޓ����Jl�ކ!$�vqUK���I$������ӆ��㽕��%䗛�"I$�K�Ü���[ t�AA��+�ʾZϛ�1����o��	�$�C/`D�^I�{����b���wH�CM�81��R�L��z�7��g��J)C_�qż�I�~V��8uǞ�Ԗvkb����&M�vv{�����*�?� ѐ � DBe��U�A&A�&����H7�O�n�wdX;P�Q���I$�������l�S�fz�̖��I��,`�fl��"� ��V�wYƲY>N�w�Mڊ�L�q���.�]++7PΌt{R��j f-i��S�|��R�ߒSׯo���:��9��%A\�<�S��z�3O\���� �C�.�t��w�KoG���v���QD��U�{���{�b#Ē5oI$�hg�!�w=�y(���
 ���@�WK��$x�D �LL�;�R��
�퇺$(r����0+ʱ'b�;�����鷲"�i9���$�p �F{Z^-���L�d�2ڢ<����|;�+ٜ��;HÓ6��3ѹ�#���0�YT��Ze���w�A �odϏF��WA�����d��ձzgzw���ޯD�|��C�"Q�jU�����h¨]�_/�����\��^}q�ƞhC3�*X�~oJ�y����.c�V����en�����$�!2&I�Ra��I�Y=-��zvh�SB�9bIY�[�E"�.�Ɖ0g���Qb)�D���1QM�6�I���ha��
i�0�^�%V��G.����-B�W[Xqm�Z,�cƃhi�X�e4ٔ.�T6f�)�P[��Q/Z�����qa���	���E7��	�T�=o�n���tLf�V�%��T1�R�iBؘ���QN����2����5�
L�k�b����B��3g��x]u� �y��>4gy��y��'=@&�hC�Ύqʞ��	��]X�,Ⱥt��Cy���<}$�*p�;-�ui=M�M7�I Q��oB ��lH$�k*s�!��ȋ����!�:t��;����ݏ9��Ή�@ ���g������>dh�c@'�w_D������
3�r��K�Df\#�d�5�I+�z$�I�~�f9�>c����M��>N�wW=,xj�{� E��f�&�ŷ�W|�H$-��A ����d�9�Ճ��Y�LY�d��PZZa��m%)KV]���E�0ʸ��s3�*Ν�k�.�g �.�9�ɎUC�A][�$;�.؈�yZÍWK�%���@!e�L���fN�;���Y:��y�`A��X��2��5R�z�&J�3Ze�$�x��I��g��o� �{=������~�S6u��р<G�Y���Gt��=��t�yw{�Mw��?�I�#2�L�� �%@$X4��MY~�G<����Q揟� ��E�z��;�m��G�A�c��"�ȳUyeF̒yV�HH�������� ���I��5W�B]�;���~]�G	��s��[��:fbl$I>�y�����]<�8��X���D^�3y�3�7#��NR�<�3�0 �� 8	���]u~5�S9&|� ���	��mv\5���L$-��u{s�aɢ�K���	w.���^kשv�%�J6[Yąg�N�w;����I���E���R떆��gWQ���$�+Y.��R�<��部���r��K��9�\X�S��]@$�]�I��Lb1>L���$?���{�ݘ�zc@�F@�	�/+<�	lf�\����>��� ����&�w�w���%��{�E,���J���8os����GT���?�y��9�n�R�� H�F"��02�L ��QS��~�������@�Gn����E��U7U���fǙ�0A �9n�G��������c��8o�.~�����A.��w�(�݆����PƳ�@]O��O>$7t�Il��Kn��o�{���x`��\��g[th��6
chG�kN��@eX��L�k�|��}a^t������xǈ�W\��Af���6����/4='�g�G^�e�P iݶ�G5�8fI�O��EOm��ѣB;q���PA�6�i��>m�O����5=Cz�
w�@O�[�,��LL�39I��I���Չ��̟/%�J�e���W��Cq$�{�Ӳep����ǫ��0�N�%s`�x�����A Y�;�Q ���X�:�Jm�j����y�(S�dR�1E�Myn���l�������Jr���}|}tNw�5p	���p�0�+��u���{������I@I�BaD�U&PI��	"O��=͊k��p�3f��L��O���TGk\�`v�$☆K�oHo����uǣ[�?&A$�fm�+**S9�j �gfkmq�Yj90�X�-�@��w���A.��w�2wa� ��$���sg�x4�x� �Mv�H+�ʾ�"b,��\�+�� �9��?�vvv�	q�n{|�K�����I����@,�G.ږ�E��a!���B��;d��
��ڙ$�f�z	��=?0��לa��˾�� �:�zd׻��-�w������Y������H���k���H$�t�g�x�J�m魷��t��:���/��x���h�V���؋p �Gg�>sʑ_��_H���g��y 9<�G�x;��9Y^��������A;�����-�(7�F���D�;{7�-ܗ���m�����<�X�c8��a�ǰ�u�1��aB�!���Ūr�2��]��y�%U�B��E�2y��?m��^�ro������ځ��/VjW/������ߌ�+�}�0|guW��}Ft�P���r*g��4�+���=�v��/g�Yڳ�P�O7�rV2$ٞ������W��uvJ�5.ft��s��-��UĜ̪8L�D�6�F=�`��9N��RJ��Υ�{"�-�s�{%�֜ﮆV���o��=5�vgy5���G+�����#����W����|�h�������O7ٳY��˞;�5��j�~�ȗ] h�C;��7�y���v;;O����s݃6sIo8.?����т�U�{�A*;Ԃ����N�$ͺ<*/�]���:KFF�\'�C.#%�YB�$L�����hk;�Z���^>�F�xՌe����k��/��ܭ�o�B�z�7���'���@��w�f>7�}>�&Zq�Ye������CצY�
�.v�|��i6�=�Mm�ԹA]�5���L�}������]9Խ�y����}�܄YW�{8�
r�q���n*6���V-��=++uu�0f�P�g�gQ���=JKsOl�Ͻ��<�<���S}�:�{{��ODv%X,�,\9���q�I9�ÐA )�q$2�gn��6��w�Vqt,��f7�p�C��.<y���hA�%��z4�I���*�!���Z�ī6�ظ�I��0MY�L�s7fҙ��RR����,����	�f�N��$-٤F����w�lM��7��%��Y��h�����(tm���*��#�Ա=J���̜���d�mUQ���`��J�,LJ ����I�X�Uj2�<�5<�Nr�&ҵ%� #��%2��+[L�|�L4jYٓS��p�νq��D�Z��Tm+p��9t�#�ʑF3�&�gf��es*���3
T��E�T�`����<a��V�vd�����C�})�Ι1I���X��36�V�YlBKz	��!C�dL�d�1�+����{.ɦ<�3,%���I�Ay-6����Q\j%Za�+(3�&��f��,C�R�݋BLI[H�&��$%J���K,������Q��4ۊ�-�2�PQ����LALpF���l���eL��H����R��q(����[�'Ru��O��R)Yr�Q̢�S���õ�(�5�Q���)��U�ei�4�kx�u͖.��8ݱ��B�d���d�ж�+x�����:��Zl�M��m�P�m� v��*S=U��ٓd����dSL�(�4��<��a
����������6(�j1��Q�͚ �;AΉ�A���ibv�\�r�Yduc1����K��6���8-eJR3����0�dWmX��n�WX�0�r�F�g��(�2�ۊ4l��������k5. �,�	5e\�L���k�ڢ[+�F[�P	nHɒ)���޶����us�b���ъSB�+.�tнx�K�[e"m��hpu&��a�v��խK���[E�LݮuAp��]G9�$V�g]MiE`6]��ʓ��#6�E��0�am���P��S��GF��N��v3@��Ktp�Ґ��\s0�F�bۙ�ؙ�V[	�Y�a4��j醙(mū�ƎX��"� 2�c),.ɱ�ԥ��i�i�3M�i-���8�׊@��k]
ꔖ��[���Dr��!�a7C-�����%1����%��i��;<ۭ�\dUG��ڶye�j\X<��X��Y-���XTy���%��M{bk21��DEз�Y��� [��3
 +�ͭ�B �������c�.��{�
@(4� ��B�F�4�
�1���f"D@`K�H��f����j�Yf�=F�h�)�����%��J�X�rl�+��.�[sI��56�F3(�R�dR#4�P�.Y�.ܺaH�6�v�lB(��m3Å�cM5�&6oU�.5��`��*��1-0gc�F:���n��L��ZL�Տ`c��.�p��	e�5A�h	-D�v�˶�w1�[�+�-3ټ����6�XYF�bd�c0��A̳0d�FfRkZJ3KBY��Xu�S#^��[(Ӧ������ �(3*� 3Î��ē�y�S�ǥ[���:��:&���0(�͚�l"<X����V�b�1�3��1��]2I��ҁ]
�;3:4nf��M�����RkP�f�8P��K�K�l�iu��v�Ŗ-n�ĉ�(�A�J�&l��ؗ[4+�Mѱ�5ι����X*ۉ��cY�.�j��V�5�e
FkͰ��h؆3jU �Բ5��΢�cK̨��Z�i�6`���"��u4�3E��ܷ�?_�T;9E����*.d�ُA���i��U�^�!G[{�]Q���N^K���� �ܰgN� Ƨ�A���+��*:�	����kO(� ���}5��ݗ�W�"�0.μ�y���3f#��{�H:��7^n:KkXM�=��9�7���<����<H��J��;Ȼ��q�R�u��2�/H��4ǒ Su�/>F��A���K���S�Mh���H,��=���g����f.����m@bI~�؟�8�N=�G��;��>$f4� ����%?8�~�ƙָ�J�@�a.q��&D�.) �D2A]u�0�"�n�\�W%����9 蝴�hsЌ'hQ�b1�^�|O��;`$��_Oz���sC�,�_����;��$w�`�N�$�pV��ܱf�,*��w��+~-r�����
�?� ��2j������a�k�֑���j׷{ۗ���gO��X5��N�5�c�uL�����{g����������ʌʤȌ��ȁ���I�sN���[ҏ��>�.��gT��A�O�$L��d'r��;�Z~Vj�R�� �z�.�a�k��^Hk��^��(Ot�ǌ��L���ט/3����b�J�����N�� g�6g��|w�,�l���#�t98���1��@'O�a�Ln�>���e^^�ׁ6v��~Ჟ�41�Z<H/ۻ�~U��~��Hy����E������Z!�M�f�&�ٺ%�I�5�p8�h��A�F�'!�������-�`A}�؟	's� �F�U��O>��R���̚�2d>atu��P�Я�g�bϵ��8A뼒�- ��W��@$Ψ�F ���=�˾��p8�hL�\:fh�����H>�ܘ@#�ټ���M)�Fݫ�I���MռM�"K{w=>��p�fݞs�y����^r��Fv���wx5���h� 8h�(x`eBa`R`BaY�fA}���x)���Ǘn͞tZ&��^���&N�:w�F�N;�士-@9}<4�vTxg����I�m�LF�Y��� �jf:D�b.%ú��A�ـ ����ޮ�O�s������++�wL����&���}|���h��u�?
�n�]vB�\�IK�	T�[y%�f���R��In0&ƞ�}R�o�jv�c<{�_o\�+�	鷀Y�q�V��8��.#���I|{v�_��f�;���vbꨎ��N,vY8Û�Dc�TFw�D�� ���GN�Ү��
�F�r#�D(/o~W��E��A!Q��a롧�C\m�O����N��A�fr;%2W\�۰6�������u��FG[���ݳ����J�˶8O�l��g���g�v�x�_x��{�~9��Xf��sG �.Mte�R1��l�L��*�5�33�d�>Vae�I�f��1$�u�s�ovk^t�K�Zs.�^"�����ؒב�P3��nz����A��2��A�c�cH�����;[��]�c]��Bie�1�-(ҼgB���.�ĳ�Jd�;�Ucr)����1�0 ��:3#�Hn�ȓ�:l��;�O ^��G� �����/��Q�m�L�3�����$Jp����wZdw�����3q/ �[��D�Y1���"9-����S����m˹��f.��ޚ�>$��݉'���VU�9tY����hC�ۏ7�w�p��$�8 ���zbʍ*��+�g��9� �CmvL�Go@�ץT�09B��x�WO%Y4ahI��?�[�nO���G_t���2ٖo�cN<	W�3�A �tD_�fn�)�x?����Zf�)���"�����d�x~���K��@�ճc�p�[��\�goc��/qݢ��3�|=�"��q����-���G2���H�BdI�&�aI�M^�hW����u#��K�����PYnt&�Sb��:лl*,2�\Sm���56�� �F�ŕc����2���M1s�1J@;#01�f#n�2Y4��j9u�tWS`0!#�R0f��B)�uZ�W"�i)W��Z[S���[����cJ�C,7Mcs�RatM5��%KHʛa��ۊ�u�HX[�����hA�ZKF������8!y%�@u��vK`y��|�����ڮ�߂!��^�O��:$�=���������Z1D�{�3zd�0�[q,��y�c�`A7&�j0ʪ����H$y��I$ވ�K�����ӹ�V��q�'�ȴ��2g5c+�dH�$y�" ߃[����^�ռ H Έ��f+�.�9��M�⊮����+ZkA�����y	^K��{b g�ד�4���U�� �	9�-�E��ք;�`��$��@_�kzuj�ժ�,o��{�D���ސ$����>������~���">M����5�k6�E�M���gh˘Jq]�-]61s4??C�������t������@ �����$����Ǫ8���Z:$�z��j"�,�2w.΃�
�ZV�1 �N�ޞ�d۵���׏�e缆\��&�����hX��H��h���M�_^�Bf�s���#��� ����u�_yo�[�Z�O~��G�P��Ȅ���3L0��2w�<���;6��y�GЈ%���ǉ:�A�n~y��E7��0^g�4gz�	�[`/�U�LZ:�k�|��A �uD	~��&;�J��"�3'HM�OC1����>,��(H@�ca�I�}:,��w�k����Y3{��;�)��gtbM�5B{�_[Y+�ڹ���C�6��"vw�N�Fgn�j �i5˄�1t�Y�����	t�AкX뉫\Dyt��+���lꆆ���v�0
N�"x�N��I|�؟2�M���u�' ;;���q�C'�n2H}$��p������]�����i4y����A|��v�B�"*��gĝU+y��;*�,Aă3�5�fN���w��)�l�|oƲz"H>/9�!��1WY]F�8�̆k���� ������|�ɗʚ)'�)w��X7��>nk�w�=�sip͑z$���}�	�>|2$�3 ̢L�2��(Я�yw��Q�x���Wo.��v�B�8���wt/3�}��F>��������[T ����$��͸��3� ���DzxJT���1d�2+9�?���������,7���-��ZLx�w"�'�ג�����{y�I!$��I��	�^t��R�P6e�h,�b䦪�Kt-Ms�*��[�p;�)��gtz=��Z�H3ћĎ�lA}� Եl�kB-x��`�A oGl��:��h$��@�؁(��O9վfŸ�!H��ɐO�a� (S @@��"�1��x���b���u��!���#=������úQ ����ȸ�19���0A w��֟kop�'�v;c�w;"'��ᡙ1w.і��umxfKu���
oobI���<�F�l\f{���or����9���p�7B~��=E}��.f:;K帻�y�>ΰ����v��q�ݩR��t�n��0�b(a�x�{ő&U�a	�(fP�|���m�ϳ�{�D��E��`��T}r� ?d6B��� R�?�?\L�3��&�d�= L������Yf��_�X���B��Ђ2��FnMΠ���^LXAй̚�Z\͈�1I��{�q�"�F���>&n���`�N�~im`��Q��"n� A��\�r��gw&�U�эG=)�е{�{� P$�}�~K��r_����s���e�r�I�/��p$��9�n��n�W�M[V9'a�)��w�~ͯMod@>$WC��$���úQ>���ݤ��0�5	#*�R^$O���b��-�lh=������2b�]�z���	;obA뻉�.����3��C���D�_L���Z&���UKw���g�7]�L�q��閹P���6m1��ĭ��2�/+k��c>~��h�|7�9��5nT6(5@ �� ����+t��֚9u��� � ��Hă0�d�u�o�٫�陭e��U�Kn��WFQW�(�ڸ�cSH��	�hM(庘v���k�F :]�#.�p0��v��r6� ��%��K�,hlB5��e��#�eV%v��Y�щ�.YX2�K�d#k�C���Y��f��%{^����I�LҠ��m��R�IuZE�km��;\d����)vk*Zܕ�e��\f�VU3iV4�\pY�������μ�*�(����%o���܋���y�~:�=�x��d��AD�_L�k2��+��p5�߈�y/�<J��0�6R�NՓ�1�`���dA9��o$��~""g;�A �{.e�g��w���v0�1����V�U�7D�H'ş1c�N���q�K�ٍ0�".�z_��|��u�����4m��O�>F�4�>1�孽�$�{�/pgYm����:��f�'(�g.҂�;��F|�-����!GCl����}1�LgnĒH=�p+��Dkz���VK*��e�]�6�2��T΀ř��.���JPB��JF��=���=ͮ���7�v嵽�1�{H� ���!��ufW(��Y�� �y� �~z�wp�y����Z0!	v�p�wcw��nL����]��$��x�j�^'u�峓2n5-��G���xV|Ja�Db���A��\a����� &F`��I�e&!���}����
����X�����{/���(g��`��aRoZ>,v��ٌ� �ݸ�Т�����o7�gn̂@ G�]{w���Y�ə<���/��t�)x�
���}V��:�q��{-��10OP����$7�SƳ��3���Ex��@��G؏CD&�Nb�Od�K['��&vs&A���O�a��ne����߸7#���g�f)���j�a]��lv�Li�D���e��J��]5���A�ϟ������2r{�]l�$n�-����|���x�4-~��ٙ7y1�@�}���zѡ�w.΃<�3�9/Bp���SF6/�ݷ �H���	4���݆K;�n��O�D�M���8^g�1�1� �;# @�X-ǀ��Sj��D����^���y����4w {��������|T��?Da����X�/.��u��*�[���t�ʼ|5ɾH��ug��1ym~-����<��M�|��zi7�Z�hn��������px�.h۪�,L��޲��3�a��=��$%�8��{?tR�����49<�w<un�§Օ��~'�i"\� ��[�g`ڸk�i������E���w��K�7�f�n�rm�㜺�ã���;<�]�n7�W;8��y$c�����?zkۡ��8�:.o۾�����a�H�3�h4Ebݘ�c���v^7�"1����zm�|LU!o���-:���K�z�{׷��OM���$(ؽ����Ǵ/oRF����ݽ��ƹ���Gn�7�J���e��}��:��g=w�=8^s;8@��1�� Dw�x;� Gf��5��c�4�[�v���}V����3xw>LF�ǯL���s�o��%	o��K�G"�Z:�������y��"��0R�< c\\�Taɛ�˻&��S�>��8�O�74��O���ݽ;�yH� ��, p[v�z�<�פ<�,!�F�s���c�=�C��$=e��偟5���� ;�n�'�_��,`;�^������^A9+�5�j�w�]�j���0�=��vw���ե��\�N�}�T�ܫ��h��)�~�:м^#����p��9�ӕnrft����[�q3��U�Ǩ���e����������6^��Mda�zzబ!���X3X��7��秝�{�ַ�UQf��G���m��m(����1�qŭQ��-c�Y������X�+5b�`%*��1�s"(�DF�(��6ł1��X���5��,����y6q�--,j��`��ng�֥kXQ�TV-�-�.1�4R�ѩJYe�MNO&�r�ЩQAv�V�+
�Ĵ�b���DV�`��jQX1�vrnvl��ԥC+k��+��n�(�
ְ���l����,-��Y.K,�������=�ZթU[kQ���[E�E��efakb�$�Ӌ��s���9J(���$DDm��l��m[�╭U�iZ�D4G�5J���eʒ�;5;;5�,Yh�F֍�--�*����Z�c-�Y,il��R����X��D���T�����nrrrs��B�h�E��6�lEIc(�e|ʠ�6�X�P�!�ѐ��C��N���*U�JU�F�µ�Ѫʍ��bR�Lk4k-���QF����dŃ 0$�L�!���>�*��ݸ�I폜B�I��G��N�W��6����;�'��I_E�O�w�g�&���ݑ5�j�+R9L����_҆MÆ��/�A�s}m��üDx�d[�=�5wL�#"����������[�(Rmm*�BkzbL����(JJ���u�%s��'vabs9������o����A��wL��m�uG4�؈����H�pP8(;3�g%�+�z,R@�wS�`[���}ݜ�A�$��x'� B:��I�{Jn�q�T�D'�c2�]�z�s��'��;`I �1��ݦ*e���m��[��oLloT���$��!cpgw���~3[[AW�z�s�@o/N[�K��̞��Wmn=�ꈿ�_�s�x�;+��nQ��m\�΀]ֺ�ε���3^V+��T��yj�ل\�l]�.�{�G���+0��L$�̀]4���#�ᢔ�0�	;UUgT�$��j!4���Q93�Ğ���Hי2 �m@�iG�Q~p�1�1��&o��W1,��H���K�ٽHgga��n��˶QSfL��n�_.����ɯ}�	�`A'���bH ��������I�1��x'���Y�'|�������i�w���r��#���|��v���D��]�#�u�����&����=x��䄉�Aݝ����]2H"�j1ڝ4ᝪbz�	&-��A$���@�r�*f�hvA�:w!�0=��72�A	���b_� �
͘�w��<��g��SEz�+:�[Ҏm"�Ub�����/3�~��@$fF>�Ďu��� �ǋ���Wl�x���b����߶��K����8p���P��Ps�pv�K�l�ev�O�:.��-Ҽ�`ٜ�S� �6��O|�n��;�ڣV_��'gu��	�y^^�)a����֋f]Bi��ӿV��/X�)050�	2�nn��ۈ�c[�����kJ�sa��p�5t(є6kn!�P��حcBhk�\� ��Tl S[IZ�a6�k0��0٩[tb�m��P�d҄�mRWC�)�6�Z�a^���uh,�/0
�2�U-�u�A�)a�,�KD�4q�˛&�6��)],f����s�����e��n����+C���s|�4&IK���4P�˛c34C-��f���53D�e��(�.�1w^�g��|������}��x�+�v�����̽�G�ͣ}��*2ffI"�f�F�;9f)ӻ/���M �F��p�-w�-瘿yf�h&�W*g�gb�LTv��$ 3U���0t]ݢA،�$�;A ��.�����$��	�h� �"rD���ٜ���P���dE�gTw6� nc��[�!��j�g���P�;l�3m�u�e�OVdB�A��6�g��w�^x�)�"���A���;Q��&}�	�٭��M<�׊^�[�%0q;}���u��6=߫��Z\�-�J��ڔԘ��C<۶-��(J;ml���ئca}|�e��L�e���7�!x�أ 1��B6��cZ�۠��ʊ��A>�h� �w���p����e��Iv�e�t�pK<��N�=Qsw�l�į�ˎe�|~沍�����1;����ם&wj-�;d�|��2�4d�w�ݒ���>>#�>!&D�a��	�&�|� �֣Tx�6�� �n�E�͗���rvp-�
�;�3坑�̪,o ��s��H5�*i';�y�$L�N�0V^�-l���:,��g�2f�h\���ݫ���o�q��J�C�����k��Uֺ�@z6�dŃ�\�Z�Eۄ�Aó����u@�]�7⊍�*b��/t5b9�� ��6X+2C���C�-?&�	�Z�Zk���Wv�1u������ɚ�K�)M��>???���u���w��=b��1�o����^$o]@�X�W��ol�
<O�ͽ��HV��Å�{�c�c�|aE�?~ �%�L���A޺~�s(��+/>�4Y�"	pS�Ft9�A�ʈ ��Ԇ�X�Φz^�zs���D���N�'nB��eDړ����*߹ܝ��B��澀g?�{��{�G<�8�ֳ:�n����I��&Y���d�N���z���~|�	ﲏ�ntӳr����^�f��eDk���cpH+�����Hv�DGkGO��z��d�8F"s.�y #�-�Y9�:,��G�.A�Q�'����3^;���q�4rû&��4�tI��ϩ��DҸՍ&!����9�����ئph[�mf�Ү���A���Yg��1ͨy>��&�#���ݨ�H�s�yq9X�,�\�����I�Qyy�h�vA�w!ڨ�Cq�o��궭��I�ʈ�1��B$���ds"��m<Ϻ�A/u�؀��;��+��~/�|�6BY]<R��[�)��$��@ ��~Cq�U��v���]+u�;�=��w#Q8Y�p����WCـs�u�G�g�B��ץP`����j�zg�����U�cp����E��I�fQN�z��*��wǱ�]L?1w:��쿺|i����U���Ϯ�'~^v�b��awdh.ƌ�~��^=��']\f@=���=�=O� �M�DUt�a���uAf)�+���L�5tiR��jL��ٚ�1t�-!�F�e�iX�4֓m/�������^`軻GsI=�������Z5�*�J�ٞ*����=�|g��`����tk�]5�!�TD��u����? �սG��.f>�2f�����t�g�;��lj���&�q�hŠ�愷.I$_C�[�+y�6I58,,n��J���҉�k�y1M���	 ��Q�ݽp H=�m�"�0o���?5�A�8�Rv��و�$���"�#7!�_����CD�� ���z|��'�X$B�r��~QZ�q�ü�s�,�X{W^ȓ���Na���5�~����Ľ�ڬD:rr7*�J�����F{\���y�7��a����`�i��d�t��0�� �"2<���3Z5m�sF�ƍ�^�f
�;6X��\��.̠�l��" 8M�жcklA�``I���K��lb�u�붖b��*�eHԻ*��K�	��aee0�l�]b2����]:  ͨk&�r\�:�#���lx�;�
�Uܪi�4#��Wh�v���fc��r[��JF�=u�M��A���f�ڬ�]t�PA#L�n8%�U.!��X�Ř��Y�.�\�6j�=���Q�v�ݑ�4�����A�O�,w��+�1
m��f_�!���n��G��P2s5�Cy����4g�]D��������b}h0	;�� �w��<�u�X��b�A-|F�$��Çg)љ�$�]���.�w����.�	��yr�x0�I�����r�beۚ��4'{���zy���H���$�v��[����ɻ��ȀH��7ww%y�dݕ��>9��+��#b�;���V�I&�j}>�P;��c�b���X(�Z����5�k,�c�:=��\Yki������m\T��j���Q���>��߶�!j��m���>H���zB���_I�c:��W�쩆�)(�ȁ��')��˻#4[���6*;m��J�m2q{����v��wO
g[F<1C*5[�z�Vm�+
��M��6���ǾE�Es,Ol^�5��d8��`
h��W�=i�ቦ$���}���US��~��>�>Q>H��O_?p��a�A"v�E(���Dy���������#�GHb���;gʙ���5�Q �w�Z��@�
-�vr�w�}n�B�!V,����zQ$�4��B�����aT�=�MtǠ���8g�9v�MG@rI��q�Xq��U�;������V�?u�%��0�%����\�Ll�-�KF%)f�An�B�
�Jh����Q��{������;�}�~ױ�������(�v1����������{��@��x��S�~!����e*/��:��A���z�� $��n�=���ل�Pb���wdfA�1 M��䎵���v�SO�Q��a
�NK�[�S{������Dv��9P������x��f_Dxo�ݨ���`��x 94>�X��f)h��K�'ăv��H$eoD�Mf�e�x�E��$��׭�"v�+=: �]����O��'�����Si���\��1y�Mϒ@�;E����]��F?�m� �A����n�M�#u����y��C�� �H=ѐ#�pPg��Ow�^b�`_ϋ5�Z\�\h�V��k1Iwa����*Ѱ��:[�Ҝ�I����_����.��΂	7����#�2 ?�եF�3U���3�ǉ'�2#Ď�h�m�3;8-�|��3s��O�mљZ�랖"��>'*� x�G�Zާv�v��[��L��W��T�1�y$�U5�	;��;0Cy/|�r�r�fΜw�~H�v��^HoLG�҅y�	ư�;p����T��q�W����A�Q�� ������~����m�`�a���832#�6��S3z�:�/�1QE:TJw�F]��nV�T�I���a�.f0w�>��ٚ��}^��}E�A!wh�SA�d};�Xo�Y�OI*��n�b�{c�Jy�����u�t����~�yeK���,�l��[�v�*���Q�3i��\8,�˻2Mt007��0]�3� �A�و>$AΎx�m�P��q3�����@ǖ�T���=L���w]�i��|X5��t͔Y��S��I'��0#��c�A~~�B5��sPnz���$	�A���gg��w��I ����O@��'��Ē{�]�a���sG��p��A�y$�T��[���Tn{���"o"<O�ycT�A�=}��L�6�[C�'�k�
���ni��N��;�3 �ۖ�^Av?<
�nGk��Z[�����O��1�u��<=+�7�G�e�V�����4>ە��;�|pdX��t�|�e��[�v��!}��h�Y�{ge�-�?��4y�{���z���;�=�\R�]���n܎M���}���Ⱦݘ*t�{�a�s��J93f�X����n�t'�г��|9[�ĠM<T]�<;ݧ���x����t�@��}޿E���=�M�q�M��߬×�����g�<%��w��g����\��6�Fo"����]�}��+���������^X���3_L�(�`:B���c���[�'7TT�5skۋ���[>���3P��|��3i�>X
���9:����߽2��xپ��s�c�����f����q���·�����;�D��*�=�S|��y��g�_��ή�kѳ=��ݒnV*Bzjwټ7˦���!y�E5��Wz�{��w��c��#�Ǚ�?Ep8��5��ܸ_fv^*z_L�7c�Z��Xr����9qK c1ƙӂ���Ώ���8a���?ajl	��o1܊�յ��I�����sp4F�N����g�j�.;|<{T�A�l�݈��B�n3�9���F�O�K�q丞�}ݝ����m�à�2��Q����z�������HL��U�f��|����{�{��p��\n�e8�X�8�׃�}-c�e�މ��ۋ�I�zW	�I�r!���XAHh�1eJ9�2�ɟ!�t.�۔g3��g$F!�����iw	O
����+aXo5\� 8� �8	e�^�@��[��_�&e�Ա���B;KH]�e���+�]珏�&x��X�xՎ�]a�a�-m�6�v�`�z+U6I�#��Q-��FʴKh+hQ4�5X�+[VԪ�
6���K�e��O'&É�K�F�մ���5��QPh��ij�Jŕ�� fEM0��5;7;6N+��PkE�U�j�E��2�V�Y[L�#U�(��Q�e�1�d����U8���d��-�ԢU-E��X�іԬ����dEZ���Y���ٽ��)j�-������*�-Jʊ���Tb6�J����S-E�D����Ռ����y7�)DeJ��*UD����G��1(��mF���L�AA�Vk3%�V�%y2Y������tZ�����hKT�*�[A��TA+Q-�X�j��ihWֳJ[�Q��ɒ̞O'�{Qv�kV��Qf�B��`��mJZ��b�mV�V�Z�Ң����ԭ*մl��fL�����TY���+j1��CT��
�[�Ӊ�X(��aiEm�W����#X�h���klD��_Rfo*8�ŭh�DQ�EӘ�-��JVW�Ţ������,�aQz�ߧ��ZW`εU�*��.�L���<���M�8Ù�4��X�J���*ĵp�l�Py�#s � 7h�֓V�	%�lG3]�[%ц&�`��4Y�:%�S�1��l�a�㕆Ŧ�r:��r6��c0[�Y�y�0�\�m���/4�����d��<��enunV�bf��e��Ku0VX�u(������#�����n� ������9n��at��R��̭��*�F-�����*`u���dvr���ؠّ�yb�����6�(�х.`62�\؍��p�!{��T�M��G4�Bţ�6R�f�H	D0n�&MȆ���4�f��EU��^�X��¡�f�k���Ոۅ�	��[��ܘ�n�R	�����u�4n]E���m��]n�E�{W%1ռ��iΩ.]h��63k4�\5�-C$�5	V�Jh�Y�$�̀*��vv43�h�n���4YU�2�9����ڦ��h�u��W��og5��&�	�,�SC*ˁ�+�g0In&r��p]�1V�2���\0�B�W:[��x��"m�ij�#j�]����+ŖL(d�bs�cL�-v�%�F9R@k�%�K�E���il�ÀS;]Up�ٌ�i{�i���⸭J���F�c(��Ĥ��Æ�ZF�j��%�q͎-�#l�-� С��Y��`WD�M�� \��fd��{]4
F4�2��T�;��f��#�Av]0M��k`V�)��5��M�|�yY��i��h�(�-e�3��f�%C�ԉR%{4�ƺ�b�ˑ�܆��l��4P��]`,��e��]��f ���Ƅq��r�B%�:af���l(�p��b�!���h0n��1�"L]����SRQ�ut������Z5�J�L&rE��n�l�B�]��;ͼ�u��m�.Mb�e`���RYL�K_��՚�beLVV1���C�,]�Ԛ��k`�k�#�%M�06/fیC,3� 1�kl26��LWP�Mk�"Rl�4�����R�f��^ͅ"�M�s���#J�G�|�iM<-�^MQԣf�Lʸ;:춦Λ�v&-%�����,Ū�.���m!��+S�Z�H�mun�5hX(@e��%�[��:"�q��
�X���%�/+a%���E�b��a���S�<:Xe�A�����uCvN�>7Q�<���$�vtA9WA��h��M��h5� ����g)��fz �y������X �����	޾�$�~�:�zw �/�J��C�.�wh~:nz<�/o^�D��T����'��g���W���n���ti��p���&;g��a�Į���I��q �ݓ�.��:�^	�Q���c�&�"N;�o2N�>�ٌ�;6`E�X5蓇k�9��|�%vVzg_ze�����L��X������IV�E��+�@#��a��U6�85�\�Ù-U��hE;p���9�A� ��^
�ALN�\@=�p�t"u��v��Z�#���[هQ0hb�OTd�F�qج.�[��Ay�+�C���as��L�ُ�7���{��=nhd����;⺧�7��{�.�zi��E�1,�Q�~|H ov��7������r�r��e>6�:Â��]��e+�\Y�p ��7�"i���3��Om�$��胾A6\A�Dj�� �K��ګ�uGe������o�( ���r ��s�=L��[.�lDv@�!��*�b,]�o;���Iё'�
��SQC1�}/� �܈	 ��<�E��#a���R��C�)�fpJV�J�@mpG��fY IS)	�Jf�땻u�'���[:�$�7��O�^\�D�H�޷�b�'��nJ��#}(�H�́{���v�ݑ�$�LUM���ӹ�q����I5]q$ O�wK�>�L�
�m�FA"�M�-1�w��D��띘�Nt�	%����rR�u8O��c���:R���>�<��Į}�E�3������%��T��ݿ�o�w$��.�y�������烙AMe��O�oK�9@���e�=��c?JY0�1�'kf=��v�^!y!9��'7P�;��� ���]���ahX�E���C��6 H;{��}j�'���n �H�"{e��D�tA,��-�_;�׈8O�Zx��	&Ĕ�-�Ԅݰ���c&%K1�xk��b����ͱ��Y�/Ͼ��ُG��Kx?�	��~����FqWn:7�D[����=$��p��I�k�W0#��^۔�[n|`7����������K��R� �;��6��v�)�s�Jz�Ny,��O�!��V��}l��[ ��A�i�!��EV�G��ӍY�w��D��Fm3�,h:�#۞�As�>��	���I����y_*j�M^=	�g�����b!_\�\<<-ӆXF<뛵S��d[٬�'0$d�I�m����GssRW��Q���{�!��[A^��L�����e��s2O��ۈκ�*hѮ��	�؀I'�� 	�k��!/�#I�%��M,tҎ�,�4h�u,ڭ����4b����}��?P�Y�;9f�Y�������s�~��=1ֹ�q�œ� bA]�A^|�b�Q���4c�^s卧tgZ��m�c�����>�;�Q���Ѵ� ���Z�xA�$6;�o:N��k��O^T�-A͐Z���{�5��H;�OZ	=�V5���gJ�{���o�+�پq�?�ov<�I��x�9G* >Y���a���	��;�l�DC�r좼z�#��AV(��<����񙫲f��<O�yyv�<^K����̤�[z��LR{���Fg��F��e��b�~�l��)���Oe�#U�s'D��R�b���Z*t�|4���7"�Id^��m�#�2	���I��<r�` YH"��q�t`�$�7y�(ܬiY\�sH��J'T&n�,�Jk��ͨd�*VX�ɦ���˖���$.aI��q��ii)-ܑ*�Y��Q�ډt�[��p��4�ʴ�haԋ���(U�h�d�큩���5�e�4�4�Kl��X䶚�a�#L�5�$�@5H�:�:+���X���JWQ��<L�j�v�[Λb6%.���f�j�`�k3��fm�%�(�)��;��F�ĝ��e�o���3�0�z��$g4��7kk91����'s� ��BH�yhZ�����f�y�j�r��H&{����]����phl��~��*��Y�(�\�k)`�v�1�0 ��[���A&V�Yޑ�(���h��g�\A͆����(1�r�Hr�j�u)�k��i64�t@�J��Cz<�m��r�d$9�N�Z�cނ'�|V5���b��i��&�5اn�ìڊz��5ފ��h1�|O�o�y������~}y������i����0��i��A�-ۘ�%�i���MnhY��4�����Y��C�r죎�l@���$@���{5ys�F�x�T?R�r�p;'I�z'Z:=�Q�n�Y�L$a��!2ƫ���2�&�"�Ƽ��a#�1�?>yʚ�{�������*�8���;ҾT�;��{k�|z��|t@w�� ]>��y/�	�$=�� �j��>�4���Z�/̗9D�gw,��P�t�s�\������n?�<S�9��ڼx��C=>G�����nX����t�@�{kn�Z�]O|�8Ym\D_���^/�>'��N�l��e꥾��X�A$5�r����ϧ6b^#�%�nWEܶPc�]R�=א'� �eG�onC�/��NPf
-,�Q��ְ��f��X�ĸ�VR���"h68����Y����ĳ��N�X;]�!��H=���� < cc0�u����[�/��F�A��]����j�Kz�s��)��A /�by/w�b;l�G;�.&�׷"p3'I��LtA �g6`A�2u`,Gks���c����zo`5�p�|te�e��hRX�@�
�}W2��f�ƕ>���)��m���w�͋�xx:�q�&�rxvKǻ���H�gg���Ct�H"�c�^<$��]}Q �O��s��Cii�>��b�
N��b�ToLy E�d~#7U�Ҧ/	��N�K������&���ؙtͿL�3Y�
S�ml[���e�v�Ȳ���\�6�Y�i{;�$�NQNXT�Cc3��]wN��	/&7�>#[y��=�8��;�|���؂I/%�?������bꨇ���[pw�1c��}�Uu�B�@������=��fYZ�D{���tQըT�5I�;X焈p�'؁	�w^f�cC�X0WV�,U6�ؾi��������f<B����r Z�����鄎yc� h�=����Os�{�=�ƙ�hI7]. �}�<H� �8I�̋�i�~o;Ś�F<۽l�Y0���o �O�s���3L�wO=��]k2y����g��k��K��Df�;�,?-Ⱦ�R�4��-�k���:�8��#�=��13�a�뙯/y�y�:׌��'�+&0��E6���c.���:�0z�����jy�w6�o~y�������^���o7^<E<�~�@�t	OdG�z�O��m�Am�ڭ��; E޶/�m�j�]X��mC��Tt���N�e��atL�;�fr0pE����t.��/�H��>'���D ]Z�ǩ���k��u�!��G9�d5���ϧ�o�$����n�Y˚�O��� ��xy5�����{q]�AD����m.��ȸg7~!�&�	������x�����"��7�ך8M=��$��8�޾�	bT4�좁��#�C�9�;��_��-���U�Ȑ	3�5|S�'D�C�'�,�'I6�t�3�I�1u
��٦\hNX�%l��"{� �7�]�P��^,�"g�SŃp�jAלY9�Y^���J2Q��{C�5$RmCI���=���*cxu�$��`V�U����3�SVLY��~XPe�2�1��m������LO����y9b��8�cG��r�q�m7,V�b7�^^t�+CB�^�+1tK��9�̨�32���ͷ]�T+��h���:�F�����2�kf�WD��h�ƹ]��r�l˳]H�A!)u�1�fћ�I[�W�42�(�e�����iV�)-W6iaæ�M �U�ҷe��Pu�e�(!w4�طl�Ymrˮ4��E֌0�1���-�:�m��E�/d�؞���'�+vpͣ�=k�1���ן7�$��m�+:���n���Y]�����pI:�joW��ڏA�$)�oFY��S��6Fn��$��ݳ<����.�Wi���O�tr4�c0.��Y@��Q �L�K��h�)��\G[���Wk��=���Yvwv%�9���7�U�"��ըϊ�u�L��EgLEy/�<�[���"V7(��i��pI��	b=��g�2�y���c��ѧ��D����'}.M[�z��l��O�O6.�'n<���d����4�g�eԗGeI�eѷF]��X]�˴XL���Eئ`�q6N�t3"�w��"�m� Ftsǋ����~�숯$H5o0 ��\����;8fO�?=�Ì2��F�ؼ �ҍ��ۯ�U�|��/�f�@3Ɍ͓Q����ҪN�3w��d\�l��g�d��	V �z"d�ӜȃwP��x�C���r�H$����z2v5�͒��}s��"=7��`I�`�ڨ���G�"�r �A����nTiCaP�$�>K;� OTsť���ԉ.�r����o0�&��F.�b��M�s�H�	�>ѯ$����x��u=�{ �~�j$��CYvwN�sY��`A$�g<�ۚyy1�>�5�� א]s��0	��4�>��H#
�.掘t1C@l\[HC,1�dݘ+�M��%��lίUXK����@�f��
����<A��A�΁яy��@�ӝ����}��d�:I���j�GE�w�8ٽ�F���Nud<���׀O�;�$�˴�_x}����������p���=�!�;�H;���Lx;��+f\�w������w}c���tX��ZP����i}����ow�I:P:
��	���M�z�|�z���m�Hd˚�1�<|G�眱|p:.���˞�=����w{2^�y�=<�x]�]�\oOl٧��/�^{ٻ�tž���)�1w���7�Qǭo�#��b���8����!�����X*t-4�^��^�Y=��gn_��7̧�r{�<��좾���b��<�o��9�������ÌE�ap�r����۴�l�2f�X3���w������>�<�p��o��u�ٯ^��M�t�V�|1��LZ���8�����sz<뫤J]C��;�*���z�	���?{�j~k˷�<_��p�Դc�9�{�����1F���/=�ޓ�	��z�a��T~X<v�zS;K>��P@ܦ�7�<���W��1}��f���0��㋦r��رHt�c���r�Ys�j8{޳�[��~W����3�3��j���=�7Ƭ��fLLgg��^A���;�\K�<��^���f�+���E���+s݋�� �fI�S :�m�u��3���}���G�C�K�'zk�w�b��6w������7�o۷os85�9��X���&������v3D�=�9�3�2�����o:%/���Ζ�@$����`8��k�'�o����˽{��A����ܦ���L&��n�z�Gۅ},���67K���}UZS֩�����z�ܫ:1t�T���%7j�:�핐Y*_y��!�d�P6���Q7/gG�U-��bb1EAm�T�Q�*
,��J4h�#Z_)�5�QE-����w2Y�S��kb�Q�e�w�L(�U�U���[j֊[BѵZ�Z[-�R��*&U�2Y�S��f��ɖ
�0PUQQKJ��䴱�aD+l�*Ă���ҽ�Y�S��PӶTm�
2�*��X���(��6_i�6��E�U��Ah��ҫF��3�R̚���ڪm�(�R�U�el��Q�r-`�g)DT1����G-%�Z:�Y�s��sj���-���cmE�,E�c7aQUW,h���P��$Q�10X���|�Y����ֶX�V�-�UDe�+A�Qh�R(�!ܺS��L,-m��%J"%���mD����j2̞O'�SN���m��R�bW��2��c(�V�Q�ѱ}��j��*"2�E�����2y7<��9h��UV%��ж� ��J�amDm��[ZPF��� �.2�!���%��ш��UQZ�j6�Ub�V-�Z
1�e�Z�����"�i[DD_[��=q�R��=��}�~������T}��@�%^��b�$샰b�T����ڮ�@��k��*�����s��{j�x�p��S��h�)�<N����t]��*�S�yyvm@�����f)�٤��U<	U����+҉ �<�cN���=�����<Q����tU����@Yhi�I�ͬCL	(�u���R�@���C���hm.���p�{͗x�os^$�����̺�|Ss�
���e��3������=4ў=P��(����y��I wvD�T�R���t-vf]ּ	�@Pb\D�f	i��=I� �����x��؃c�vז��^�Έ�Q�y�/[6��8.��4�<j;Z
�5�ț�I��x ���؈$��c�zD�m���s����.�ԉ�r�$ g�b�/��y����o p�/��^�9�6̲�Y����V��� ����~� ��H��߱��]��gk����z|�6vq��Wk�2��ǻ��|Ȃ@'�����G.�h��'�z�����|�4����q/_���f]؏�$�e�0CT�e	M,դ�+ֲ������{�����)wt���:�`@$5ls@���M(S�SÄ?�}2�����Ψ���xH�	���p�`Ux��(���6sp9-V�|O����x��� Hݡ��/v{r�n�<�A1�}�]Qz א�����M5T��3(7�v���	nG���7�l_��o7|ut>��v��Ϻne3l*��[�@���I9�-�u��}�}�rmEO^O�x���F��bft�:g�*������Nn�I��{,��q$�r�ր�H��nt��)߽��?VA}6d�٧����FL�};}�Od�=q9<;Ϯ�O��G@nN{����d�|	CXuٽ�@�T��-������ch� 0&�~N���Ñ�,Qb�Z�#5�m������M)	]c���16ҙ�/aJ�vv���5�[6�\֑�WX�K1oj��R0���B�������E�q�.����(��%e�qtz�j��."h�S7��i���F��
�*�hWL$Yk5XQv���ե�4���	)�ج7 @�J�jg�k�A����MA4���ى 7�ړ�.
�hYc1��ZD1R؍�z�rjni�D؎q��=�����nv�;o��l��K��r� ��}e�t��m�q����#��4x��YN\�!���,�WS�]�4aQ=�� ��L��<A�w�z�²�t%.�����L����I;�� �	�=�ft_��`�=����� ���J6��=3�1�@�E�h�/#�oMW{���O�|<y"7b<H �=����{�%UC�V�LI	�A�
����͘f93[��U������By!wy	=�1!g>�z)��)E
�km�ν����-a� 8�m,SQT��suĿ������Y��'gL�$�jbo�C5����H�dDw��h;�}��
	&=u�2K�K�\�����>�w`��z�%(H��xIQ�SS��vFD��9 �x=�́�}o>�2s�ۇ��� ����9[�}��G��'��=��NeJ�iQ<fQ����7Ċ��g��m�@�N�{�x���H��Xy ���t݁,��YUGl��=�0 ���U�s8Q�+�+��@'�m��ш�Wi�c\39wbɃϳ�x�j��~z�S���3��L�"I�1 �9FcN[��m���웈�^ߺ��w!�	�f�'<E�A$��룘o(ݝ�D�=DH��q ��-��ؘ1s9��G�H�̑�Đ����3A)len�x%��7b�����\[ &�[M�d���`�u�:����J-�ă^5�r����5��_�ˍ�SƝk��3�e�C^ʶfw	;�p��wX+�=-�8�^��$�����I��x�y.�h���fQ-�LZ�r�v�;L����H!�2�9ck��c�Mp��L�
�TBk����vMv�^z�"�ff��i���BSd_���
�	�g�q�9px�nIɌgjɷfT� -����}��<	/�� �~έ�.��d��]U{g��n>@�(��&=���\�O��s��s��|����{��GD�p��ӆLQ�"��x-�CT>�錹�ˤ���@ ��}>� �^nޯL��-�!�&��:�7e�l�Sj��A����WB�vF�sS2�zo��wA���f��ʍ� �c�A�/#9��5v��/8���9��Z�\s����P!'*�E�Dx�ub�`��ݽ�[o�
�Cޡ�[�#=*��rws�:NL�� =�����L�3寮C�C�B �v��H,�ѽ��̶�U]�� ��z ߞ�ٗ弜�v�U��n݆פ�Kc|E�l�vC�$wu���+n!�S�4�4c1��LL&�&S �X�~��;�|/�/Lr���ߟq��,�����їx��WD�Vq+6��^RJj��{�g=��'t�9u���O��.#B�i]|�xH��x$'/�W�|{�"3w��,]�X�/ب���0N�툓 ���8�lk�ū-%�p��9R[h�0Qq���.�˧�?p"�a�x�f�A �ou�`�ئ�-��g�6L�z����f�$JήI�݃�<��WS�����+�8Dyyv�"	$�w<z�E��Y�[��I7�(�bAl�@����I񭻁^E�e4��%���k��@�� ������$�<3�S8N�X�W�Y�T5azY�|��zx /%�;6�3�'M�У7��ӫ��5��FK�6f[%Ĺo'!��Ux�t�@�$��m|ε��惮��7{1 �ݸ��@n�A��lz'�1=+���ҿ�x}Jg9���wj�_s�;583�׆��F"��:�U�6�j��VN�W�+��pQ��lo��?��H�7��3kQ7��|��}yW��t�����`���&ql���䉮�F)eK����3��p��QJ9�Mu��cl��Mnf�plE
�-a�q��c��Q]]��[��Qn�R��h�.�؃K6hJn��҂�邑�c{f�X�8RRŬ�f��s�do&�u^[%J�����Kjk��2�ڪ9���tu&vѹK�K�e!V�ٛB��aˉ��[]u��39b�9u�7j`Ey#��$Y��w��9�>�슇{�$�˸|����w	�;	�=S����T���k�6�@^KŎ�?���r*��Af,e��M.��a�'�h���	��7��{���gi��U��cĒz����4G
s�ȃ.	.���w7��mq�#"�� 2�'��T@����_���rf�$9 ���:΁L�8g�,f�<�;u����nΘi}ٿ_�	U{�e�m �H��-�Z4���w�6���@�,�"���&��j,e��CZ�z�׍��a5����)��<��%޽��K��!�;w���,w2ߗ�'»z5��T4F��Qj� ����Z�lmb	�1E?����OL@t��<!�[tTϞ,�5ܮz�������MT��h�s݇�K���\��m�<����%jZ��T�)k����mEܻ����<�}�A�yG�;Z��"(��oY�������I;gXp��wfL��.����f���3�$)�ӸC r�����Kz�5&kvr���P=Q���H�Á	VUwLB8H,�sn '��e�ld�<aS��b�ư	ћ��$�#3�;�|O��Th����V"E��h�[{�D���>�nt!m��߇��K�X�e`�m)6�uS��ц٦m�0[@��s��;')�X+���pϼ�h �{��I$�^&!�aP<���W����zSRO�|���w��s�`���Fb"�����A{�=ǚ�w��}�̪� _�쨼H����T�P��=yQ.�g�CF�L�%�t��}��~��Cu���"d�罝!�"�r��vb�Hk��%ȍ%��*,4\�����ˡ�Awv�y!��������:.��v%ݙ0zz��֫N��/ă՘�	�[O��~g����$=�Dx�>��ԙ���[�w�R&����b�O�W}x��X=�O{n�
�	���� ���iw�8��1Q��}j�j��W*r��v�a�tr�iz��c�OS���O�g�^�y�p޵�A!���	�Ȍ9�������72��'�тt��fp\3�_�OK�G���EN�K� �EwT@ W�(>��V�!o6ku��>�,V�]�C�v��~ف��~M��anr��1�I��^�	�ʏ@$�����dM�E�0b��]NT��DKWj:�d��{��A�'|�݈G�#Z�Z٦J̃� 5S̡Fy���z�K^����^�└{��W��˥�oi��U�$r,���[���d�z/9�7��	2���b�;�ffޟP��s�� ��ȃ]2j[-��u���v��_�z]�Aշ�8�ۢ�:�]��wN�윰A�Ѝ�f�%�,�"G6��`�l��hgS2�i����/����4C)��7s ��t$�9��rҫ�t�T_�`@$���ѱ����IvcTc��	5��I~9���>z4�I�۽���w� ��7��e�w^�^�DO��E���g�<Im��fv��~C2ð�4𹗓�X��m�;�G����g��X��x�d�Tu͚͗�3|	9��H$M���H��a����dNw<M�t���]E�����B|�^<z9D�a��m�$.���/"{�7�&<�e������B|ux鏳q�U��̾����,b��?L��Ѯ��wkg��8]�0����}b���(r��k�bv>ʰu������f�;ܳ�$��{�Yuўm�}49���wý�6��uD�O}8c��U��z�=�U��]L�=��֞�{.��w�)���;ܒ�:�]>w��v��}��cV[�ܞy�vq>؛�bڎ���ݶ��;��}�������L�{e��lP��)״M����>3����kq���i~��4��ňN�^C��u�|����fzᜎ�k;�������rp|��]����ќ�}F��Oj�����Y4��~�4Oxa�]��������� .�ٽ?v��g����o���}��TX���gܩ4]�#�'����������Gx��06����}{|vLu��t4L�^��Q�槇u��m�M��ͽQl�+��hZ_5�Q/PŏS>�i��\������-����n� gՕ=�e{L3���*ܠ�K��`��#�^�1;��ϰ
��s�h�3���!����=�����q���Σ��3�ݞ�~�
9��Ѵ5���i/��7کx��eL��ǵ��-�Nܷݾ�[<��<&@{�8=px�3�*�|4`U�^���6�\�
�q4��d��c�9��w�l���D���պ�8a0�-�y�
y���� ����_�y��[oǁ<R,NZ-A󻛚.9��2Ƙó8R���p�.o�1�t�^>"L�����k|`k�l�95*s�9����~��}z��Z��F$���v�-s��E�#��狭!��0�~g�о!��ï�>S�!h��6�5��|�s���%5�wK�j��;��Kݥ�{�P3��P��Fܡ��QEQkb�-T�K-%F#R�*UE��ci�̙7;?����崢	X6��c��:Ij��Q�[m���6�H�E���"�-��+�m�&NN�&���Q�,X"~J�4�J�
%����cFQQb��Q�F��X"�1��c,���ٸkb�eA�����D�H�ZYZ"��XZPb0Z״1&U�ɓ&N��͛6�Am��kUV�Zj�ʱ�[m��T��(�V��R�QmmV��UaX�Z��̜������m�DE-��J1|e���(Db���m��"�j�f"�e��S�e����M��h���Fյ(�����U�(�U��R�T�7+B�5%�V��V/��2y<�MmZ#Fq�����m�7��ږ*�1b2��J�\W �(1Y�e�;;;5�j������Фe�����B�-�mQE���mF	Ej#�c��e��ZV�յmmm�dj���oS1��b8�UQR@�^Ϟ&v�-6U`�:��^n& n��Mu����aP*n��L�
��V6X�vt�ջ^"�Z�)�n�y�kK�D�k�L;���=�!��Ԅ�)qΖ]E)�j6��-�RlL��#��XV(P6��Җ�b����EJ��)e/Q���L൶�r�M�"]nڑ�*��jmu��d�J0,ʬ`��d-r��H��RirK)�eݠ�^M;tR�J�6�G+�Z�V�f.���Z�4�[*+�j�\�E�Y�IL�͜�R��Y��S"5�P�e�9H��F�\�L#LԄ*l�.�B�Q�Rܺ%	����WRZ��iR�FQ�P���{8ҖaittE+�Pu5cl�$�1,KKEq4�ʲ�@�!
�-���%���E��г�!i�۱#�d�#����s�A�Gl0IV�<հ��VZZ�pV3Wd��s�m��4`�i���4���B��l.3QvV��]*b��ob�cj4��u�k*�f���[A�Ŭ�M����ɪ�e�7+-).ܔ�EHW�5ڍ���G3��5�vBpAhi+�KB1�*MN���^EW6g-�Pl��J��e��\X�Myu�V�`h�22	�\��3��Wie���\�e&�l3Ra�"`�b��ڕ�"�.%YK{�s��ŧmdѶh+Jnf���jm�2�0�7usd����6�n�5�Ĵ�s+b��K6� ��̀ƫ�,ԩ�Sm(L�I�����.،n���s�l%S�I�"� ���S�XkQ�7Dc�8r�c�IsG�q�E��.XØ	�β��њ7��k۞4!���]������P�b�tZlJ��.eR��K�[[��3�Kz�ȸ��ZK�3hKH��K6��L�U������Tٛ��Vhe�u�"8z��`����tV�vs..Ϋ-3�+�Y�b�ʬs��q&�c5CQh����PUtЛ=����4WM�[���5XLĔ��Q�[T��Ռ���!�X��e��l��α��Ul��tu�+45�M%��;P�L�J��\]T����1�i6��b�:5�pqe�2�Yp�Z�M��4��Xv�2��Ѓ���ɶn�8�Mu.�1!�\8n�Մ�f�)�3	��1�=�~�cGv�?~<wm� os^	���p ]��|��>$G�3fW�kI5:N��4C(^�.�̟O��֭>��fWkh4Iͼx$�\G��Y�i���6=cc�3Q	ؒ��W�k�G���o��\�;��K옏$#�
�ȃ>A��
���&��.�z�Zy��u���N���<��S�$	�#r� y\�zw7p���cYQ��������.�&7��Ė�l1���W��V�i{k̏��D@��>5�� Co=��kX�=� �}�@,/��״݌@�� [R����L���G[�h��:d�F�b!˳�C�]§� u�x��n#iLʺ�<N�e�S�>'ƻn ���6'ٙ�ݜ�h����������غ�8���v�.в�2�K)��e�]���m*�*ֽ<r���8߹kw�cW֧���ז��IM�dU�}�U��r����~$�H�ˈ�x���\�z�w����5��&jEԼ�e��������7�� �g�4ׯ�;։��� ��sq�G{��f���ƪ*z��.�uݠ��6���d)>�W���k� �����S]l���<�yy�E���g�=Qc;����gkǁ����L,\^� H$�v�^^DVwD�=����~a�2��ne�Ҙ�jn�e�8áZ�CP�*���Y��T��|����Wp�����	1���>��H,�_t�x���S��&}AG>��x��8��7ȇ.�C�]L����<���!p�vqC��P�'��Gs�$��}�w��Ѱ��2q��LbHxs�	�1vL��� �;3^�����w�"#"q[Ȟ�cv&&����͔}�Y����~nv&�^��vnu�;ܳ{�,r�^�{x���){�r��x{�N�� ���I��'�ă�:�f����h�[�×9,���a���$�Ȩ�{Ă{����V��9'�wI�Û� �E<���f��;c�'��*�����{4��*�8$�d<sob	�'�* �9�/�Xi�r�"Dײ7Xz�Ako�����@h��&��]aֱM�.Yt�Y����+������r��,g���D
�_lD�	 wmC�L�c��p4L��Oe�A�=e[�v�wA�h똂{k����D����/�6��z<	S2[��Y���d׶r�v!˪�s��X��������Ψw�I��ِH$�\�{�։�b왃̀D��=w�uT�e�� ˒J���	��TA3�t�	�����vj�Y����f﮵�>�o���\Oq�*����V�9ծ�ma-1�.�6W�z�	�v�,(X���y*빒}�I;�I&m	���ez�b	$fFǡ���-��� 5��$nt���Q%��~���q-�\��f0�2�%.l�ٰ	RmgK	�0nb��S,4(�l1CcKg����G�2��3��	3�/ �s����>�]y1QG;� ��Er,�];����O���|���T�O���W4�	9�� ϒ�������d����<���v� �0����>AMMEf2��H3�OFA'�{�Hؐz��Nɐv!˥몙xk\����Hi� ��跂I�ރ��Zs*�=5_ݔ�PtX2.ɘ=7�W�nT��_s�9L���Y��d�w�N<K�'����3����[��-7"ޙ�I%���NI�7��`�!����4�i�躣KKC��݊{Ӥ����<�k��L��@���ϐ�SF.�°F�H�
G+Eaǅ�/��Г>RoY�Cs+2�r�aeJ�F�	�]DΎ���rR��b��f4vl�5�s�4�X�fє%j8T��mT��h���.��q+lY�Q4KR�ň������a���2\h�[)���%60�ڬ��#0��&�Kc�ݷA)wj`���V�cMn�ڔD�L)��8��JX����3ǂyl�d��)V�KA�f��&]`�똘v�1�;F��P��E�ZҫRf�S@o����h����+���_u�HfF��@�OoD=�[&������tc�dփ�`�fC�tG��yN>]}���}�@A$���H'�OoDKy1��lk'���0o�lVr.���A�슧�O���ǉ'Ŕ*�=I��*�A'���x�NwD�XYw�ؐ�����Mn�w`�B�ǀ9�� H�ݹMي6���R�� {bwd�R�wJ�ٵQ����ǟ.=s�8���fk:���y�	9Y� ��wS+T�m���s��&�3;�L��(�B��#Ϋ�u��U���X�^�P)�o�^���0X2.ɘ?p"�bl�x���(��k!��Ng�\sG��<mw<����%1��* �C)�=�~������r��E^D��c\1��O6�d�ӓ���#������g&%I��v�ɲ�>0��b���)C�� zKTs�O�gs�$���t�J`sv�9��������"��f���F��	��wdǊx�m��:r�`!���dA �u��@on��S�wwI{��U��y�NF>uqq��GvD׈� 5ۈ$6��p�F�;bړ]P��/R[�v%��u�ƻi�¼�|]��oO#]��.���]K� �f����mn�aB���+��w��'�4�ƭL��[�eZPL���VWMl���{e ˹`�z���	�c1f����{���3y\ �>H����B3����{ݍ��'ă�w�ۖ�Pt�D4RǺ;OI�|���߇���]�W�'��p��R�??J�_�vVwC�t�~36
Evm���Ln �C(/O�����f�l^D���@n��hsG����з�x�x�U�Iͱ����ѫ#T������$/|f�o�E�k�D�꥘���jW��4�0��j��{��zq�k�tc�,���:f)G ��x��d�|�Y�s ��of<H$uoF��|~�;:/\➮=<�%;�wrQw�'�j��4�A^t��Y����c&�ωW�sV!���Z��V���g��F�6�,#��n���D���A�w[
�kr-r��	sή�.����o����]��l���$v�@��l��`�A�-�Q �[qA6���Y�r���ҷ�#�Аr�i����i��w�?>�9���>�A!jn���d�1tDd��cdAof���E�3�vW�٢|��W��Aё�8�뫟s�^e�@��� �7�"�$��V�E�Dxcj�0;p�6�o���7�"g�^�Fx� �w�Z�-�Ȩ�=q�aL�U��tPpS&�A����oh��j��>�>^WwQ�=�I�*�t^���I��u�|�����vosc���hɈL֯P� Ł!d?&=c�	Mn;�b�P3�<���y�C^u�??dlƾ�1��6�do���1�v*7dSk��F�igEfɋ�%�r�̬]J���eՆ`�K��6��_?'�aTU�N������{��L� H�ꀃ��Su�^��z0O���� �^�T�mbؖ.��
�k���=]j�����@�o/` ���1Q/���g�2u�9�X3���Q>�ځy ���dA��07��$�{�/�[9�@��X�^<I]0 �pA�c`�Ȼ&`�`�sG��n/j����';%���77rۤ��;��[5+�cz�=Y�N0tX�g�1F�-�Ď�t��5�s1zѯ4��=�Jl�{�m�Kko(�"|��5�T�fi��q!P��( n.����c�����4~~&�'l�Ɠ�{�󸈟zy�t���Nm��ޣ��,(�Rw�Z���8j�W@��c�6~I��Տ�1`�#5a�du�E��)#+J9f�JL�,�0��B�l{h̗D�kKX�hf�g:$K]3��iYR�\�E��`k.V�-�����2i�T)�b���̐�����~����r�tX�M���Ř!Hi���eٷ���X4���
	1簧JS6�I]���	�c	 ��Vj���A�ٺGL�ˣGK��&�D�3�kp�%R*879��*6Vl��}�|�}c�tȥ��+��[�I-���l�5�D�L�|38��>�[:� !�$�	�����Q����í��nۧ�|H$�_Tz@im� �	yots���cgq٘'bX�V#jak]��7����v���b2�g ����@ ���4�2�9�p�3��:S";�9����hn4ױ�@>-ʭ@ ��D�kV{�l��z� A�uކ���Ȼ&`�.V�y��Ȝ��w�|8()ϨZn�KS]��@u�D�֤.}���2��٘9k��ʶZ.���m�����b&Ea���B�-nMR����>���z}�ŵ^@bO�����x��{zw�|��8��^M�����t3[�N�J�lM���}<Á�N��jaV�s56��>/"������ǈ�h�n{|��ݟ�/[IƩ%�q�fK�l�B�yO�9��S����o?7�R�PO��Qc��~H�9h�J�神㼀>��'Bg���@��$����6\���հ�#kzS��30Nıv�GtJ�/�&��
����Ȩ��2�/";c�A&��#��s��BQ6�	��X�9H3�3^�ۙ$f�z&�3{rY���#ԧ����	 Uf���'���v����n����%�2�1woC��[I�!���`�+.6��Ip��Y],2�+����?�4�\�0~�������׏A��TAg�tK��h$�W}� V�l�Ø�W�\�ZC�˶OM/��H��x�>'�{�=�:�;�sz��X�<��wv,���A���aZ�� �W�4�����e"�0ӓt��pzE+�g��+|x/���'�:9j�^�o�d`����4b�(��9wf�ed�SxяY&��a�7Z�"�ߖ9�6M�@7�����:>~S��	���fe�bQ6�=O"p�܃-V�Y�G+~^K�)_�pW���4���8y0�wN�����^n��g#��t^U��!o�7�{|h�^�����.Vv�{�k`�����__/u��9��of%��L�'�X��{;�ox��Om`�3��ͅ*u��}����]8�Z���f���M��)/,�/9�f���������`�C䎉��{��{|n6��<N�#�\�"�ȋ��{����nAGi˚*��뻧|y�u`���l��^��KN%�P�FA��\�Mm�h�_���x�����W<���w�ӑHN鮬JSJ\��-;��y�x����;��Z�qoE��)1���j��x�P|�wM�l��^:��R'������{9a��0g���F���5�5}L�tG2�d�py?W����nd���v��"��^��Y����*DgN���ި��މq埨��1��j9�ۧ��3���E㷧Q��I���{��9��Ds\>Ӻv��iy��{,[��{_$�'6�~:�&<G��^��w[�6�P'f�Sk�8{8b����ϭ:�֖Ra]{N�'2�=d�Q{l�e�(4VT�F����%�էZ��\D�Y2�k�m�s��5�P����|0p){˙��+�S�E%�m
�Q�QJ���0F$b�H(*������2̝��M��vQ�m("��-����TU�ZR���)ZT�w�+Ģ,b�b�4ԊG%�d�����vZ��b�F(?�g�f��To��UR1f%R���eʪ�c�S�T�2Y���?M�E�E�
���8�1�"5(�b%kJ�o�(�լ��J����fMM�M�V*���"եUe"�DDԥETCZ�jUU�(bQ�YD����%�d�����Ъ,T"��TPY�Ֆ2��G�QVz�X���"D���bEa��#,���{7��QV�J�QeJ�ŶV��mX��A�J<���*d��b�����2YfNNNMv�Z(��J%9�1����TE�"��Ub�m�aF�
�eOѹkR�j��]<<8�I�D�ui�.ѢV#8R�V���եUTuh�PP�[j�&{���DAWl�`�������ĸQ#r�Lr�-¸�6"0bŭEfb	+V��=Y�]�|�q�>��$��� ����N΄�c�U��ou��~H��<x����y �˫�����ᦞq>ǋ�f`�� �H���A$5}q�ͧ<�������� �˧	�y��1K5L1����GT��ڒ�)�R�mhŴ%��1�xm�)p&U�j䢝�����p\���g1��6��IyQ�˻���P�u;�Y>Q��#���Yi:,Hvdd-=G�����1\���UV�A9WO �G��4.�``��sO��Xɾ�i�pҠ:xs�dA'Ŏ��0�����ۘ��k���E�(:��^0��Tᓺ(~�ٮ�Vz�*�����	e�� �uoF�����3z޳��3��sL�%����`���M�3'h]��Z��o=i���/�yf��:a � 2�f7Ȭi ��5m7��w�!��0W�{�g��g�Ot������^ް:;����#Ė7��O��s��b�.�k��� ؤ�L�,X�!�\���յt�B��Z��Z.�ʬ$�iq��IޫsY��p�����3�0IcW��_���.��� {� G�$2����C=[9���9�w1�y�z��:, �U�@9����d��w.�����^�ٸ1�tX��X�Q�/p�Ofs��g��w&M^��/Y���{<_�kyċ�^�L���Ù~=sّ��6\M��9�[�.G�3��O�wW?|�2i�2`�}
c�<H�ބu�-�@6�_�  ���%�w�t�Wl�[�䛭��x��@$� ��{�ﳥߌNs�ǉ�B���*-�.1d[�Nd&���PR^5��kɹ5��ѥ�t�\5��xޫO�C9&ؑX�Є������ۘ-i���'>>	�7�M+mL�u�[�M��|�x
�9��Q�VYU%��C2��̱�]r�m��4:È�L��i�M��c�0�
Q�d锤l���0�%j�ԨGr6��P�����YH+�+m�A l�F��)����m��*ᄮ�1��) ƚecYs�0��-�48���Ҽj+"��(=�iu���YWD4��D�5]Qn��6:RP$�أu"��CM���֬DL��D'���g��g�w�,o��Ǘ�ͼx �	����[��va�����3��b�oY��p�C�uh�u<E]�����rW�Y�� �C��!�S�ܵf��U��{���FE�D�g�I�����o�G�m�3m�Y�s�O8s)`$��	zy��SH,��%رx�R�33:^[��z�CD��G*��}>I����f�����������>��]:-*�h�2q��I�Z������M���etgN��|J��PmOr��]�{a��ߧ�Sۦ��[`Ʀ�C)�]q��Z�L�&�n�V鵫��|�5��sJ��l�A ?��n�-�y���PU�cmr�֦��/*�@"z{&K�*pR)�;������j����fv�������uLNn��>���f�Q��5=�n��{6א8��Fկ=s۾����n������Rk��O5�C�`p J�q���7�ɕd@ ���_yA ��V:���SxN��s���p�C�uT1WN<��v�,��N����;�O�T�@ �.��nB'ӓ|��r�)3��Et�}�sJT��4W�f���Q�~��%�1�o�}Ϫ<o�Έ�L�=_c���k۠��l�x�A �p�r:!��b��+��H;��_���Y�����i���3��(� :��k�;��R ��%�/�\/h�2�b�����ۊZ������.���ˀ�ؤ�w��vt[T)�G��A �Y�s���M5u!�D!&���fl�X�Ɲ�gI��]7� �s����pӍ�H�$���$��[�#�nY�y,���]��м��&.3�I��;�̞�Q�ēy���OS�s���А����)������w�J�//��
��{ ؉^^����Qz�뼥s̬�2n�Ž�L<M,Q��#��8�+l�����	Q9���;2A�u���B*|l�;])�e�@'ă�=�C5	���tt_��qt�1q��÷��)3��Զ�@ ���@��ҭ���f�P|�� ����Zt)�GF��	/�"� x�u�&�3�
U�
dÊ��e��nʇ�)���M��r:!��g]��l����y�y My/o\��p�^�нR.��@$�^gD'n�PvtZ��wh&�z�"+ŭ����=��l1�ϕ_t�����=R=}�:�K.�hl�ZM�<1RND:��~$�]<�H*�i��mKe\�9��X<k�
�ȏH=��#��f�8��ݙ�2b�`�Qْ_*9���v��x��H�v�	�X�˯%��t��SO�Wd���#'��1GS2���l@��_n������y�����/t�1ݕJ���c3)�%qj*��e��CG������zd���rk���'fH:���[�o$Z�d
���r6R��y6�'��O���v�Csw �y��d�=�xV�#|��\�0����i�	z���umP�vM����~33D�uϙ�����^��A ���<mm6wKwl2����n ����F^��@��X;ujWJ���g̦�]O��{��Ȃ\�j�W�u��xd^�'�î�HvtZ`1wh����/�>�t�	�f�1���r�z�w��^��x���O�a 샲2p�: ���������u�[S�b6F$��	'+�2��C`}�
j��>E�I�˳�v`��wA>�q����Hn|��Cu?G���<{#����^��^&�d[PL��˩�B��{۲���q�wݯ�X#H�o���t�@������K�G,=�AΟ�5>�0lߓ���d�`��1c����떖��f�9�K�D�����R�	��.��ђ��5�g:e�\�e���`1L�P׆�#�(�68�u�ј��۪�]�-mSP�a��[Aoh�f"LFgKf Cg���M3�SvNW`���@����� �.�3��\���l�/��6u�`"\�&)-۵,9ظ�0m��E
An����õ�A��6�1�%�4�"��,��4�b^P:�4Ŭ�f���r�L�WΞ�_??YXe	��?R����@%�[��uoL{M���P*k"<C��`����p�9.JvuO����5����0�<H$�}&A$�Xkw<A�;\�����3���arY�`��uvrn^�9�^ &��=5��{�P��7ʁ��<��	�u�E���u����vu(�V���i�ǫ�5�D�1���A �ݲ ����ΝlЁ9ّ��dܭ38NUUEtA!������w�9�� ��p0�wT���>���Ӹ�RHaG�e�e��G�t]�b�����W��� r�5X��t����ڵȺ��?<^���~��  M먀y���t��6U�ez��L��@%�/��fL��u2z�b�����:Rs?��}��#��Or���wB�˔���c��zl�>�56�lM��}+
��!�b�Y6�P�n��Ukf�a>�{��E�i�byA���e�Ը<�v�xp%��ÿ�����^�� ��˘��sh�7�"tW���x$w��:�E%�&	اP�S�vdh�m�[����Oesŀ$�m��I-�ܓ��|���G^�@Q箱A�س�ΠD�Y����y_)x�����G�_��$:� H����[F�+����]����@֌p��fip<h�j0�mc2�J.�a����4c�_�_��" �ָ�G��ܠ�������zw"���|��|Ҋwgg.���-h�&��I�fI_�w5�w��[~����w� ��qTy��K�T�&%س`�d�G@�W͆�e��瞟fWw��8�{F�Xhxs��007𵩗%75�����t-�_v�އ8�~>kw�Q�dC������7p8yWDVkq��U�M������L�w�Q�{f���� f�/�3�%y@Y�dA��x��UN[#���%�j=nؚ.K8L�N�MN����9���q�OvTG�*���$��D�[�T�����$�DM�	Ņ�3bܭK]�-�+��t�-��[�T������e�~�-�y�A��p�n��@��9�::qݵv[SGM��,��V5�'=�b���v ��?U�y���0�:��f9��҉�[�����v�S�⧢��Nd�k���ȉ{�wwg.���St�ޕ����Hi:u'\[�T�8�I��$w��9�0.�0v��Tv�E�����
� �T�I�;���>K��}���Vg̙¹�,�fBL�݁'���m��QnQ7팾���%�z1�ϗ-+vŷZb�T�8/�f�w��4�`��eܺ&%�;U��Euc�kQgkV0$z����Dy�>k݁��|5s��3�:тy�� F�!��"�g���k/0v�54��J9�p�`qiP3:�Si����>4��S��ju�y"os^�s�w�'��cZ�9]��o&	&�:	�I��6������X/�q��ُF�C�������n��|H켈���{� G��i��;7�xxǩ��T���	�T�~�������*ɩ�ӱY7�E�P,�� ��v���.������C�T����˺Ӭ��M<�H �θ�|	��e<t�3eW\
ͯ$��4�s�`]�w�2g�g� �_�� Q�ٛx��}�R!�f#�<���q �6����<'�>Ϩ��[�����n8�TQ^/��E TK��U���*(��?`SE��  g],a�3M@0�(@2��@0
�@7P()�Nݸd�!l	BB�����@��&@�7�\&��&�&@ 0 �%0 � $
� �(@2*�� � ZӤ��(` ��e$JdD$J` ��U��� Ƞr��`P�&�eE��i�V�V��V��HP10�´��$�������"��"�2�0��B��D���@Ą����!02��"@�+���"�43"��L��+0$��3(,�0�J�!L�! ��C
,�� �(� ���ߏ���:�������^�����*" ıPo��q�����3����:����������/�ޟ����@�O�~�����<�/���G�u����t������'����_Og�_x �+��߿��l?���0EE��$VH�����=g ��?B}���|e�>?�|����� E}��������9��F��k��3�����hq��_�<��x
v:�9�k���G�=A�Z/��a  *=k@ �~�]*,H+	 ?ؕL��J�B+$"� ��Ĩ�+@��")
!J��*�P��� %" 'F� 	B�"!�� �Ш��*- �*,*�(�*pH�TX�HE`�IQfEX%E�QfTY�V%E�X$�AXBTY�YQa�BYQaeE�$U�!E�`�!E��V�XXBQYTYRXIQeIQ`	``�VAYHEbXeE��IQd!E���
�Y	fA^�ph�X��?'��O� ��u�(�� B��g�|�����}�����������a��y��������}޾� ����k���u~S����>�2��w�!�ƽG��?I�����������K��:�|Ԁ"���f:<��?hz�����?c����TE}`(��P|M,w��IߑEE�h<��8�<��R�+!���}��9OW`{���OBr����x�G���N��@p��"��z�����'���Nz=�(���>����h��������<���:�C��?z}G��<�H|O`P~ y'���װ~��_���H(����zR�`��� ��������Ǒ�}��� �|��������=^����>�xyQ,A��g�o`=Op�;O�|{���"��n=�u�3�:G�>��r@�}u����߽>�{�G�o����2{S���ǒz�������w��>��w,TQ~��zN�>�#�ö��v��}������^�������e5��H��B�Ř ?�s2}p"?�n          @                            l+��RE *��H� �-��(RBI

���R�(H(� @�UR�(( (
�U �|                                     x   T        � ���!J͂ �wPDb` a�u��TA����PVw/x 7T��g��j�)I�'x   ��:
��j� tУ�-
��JU�wJ��՚�a��;8 ԅLC9����T�eR�CT�N`�t*�����
�            C*�R��uy`*��2R�ocW��R��qAT.�� �TJ��w�(U)�c��z�J�;�T)y��t
C �A���9���$��   �nc�TY�A, �FB���בO ^)T�p ꃮ't�r5��B��s�PP("�   <         o���
������q��=�.��[i� �ʔ�6Ҵ�ë���㫶��Y
�e� v(����Q˻�**�!x  ���
�7��cp 9�f��k�J.���lX��*�8 :73q`s]�a^�=zm�f��5`@�W�  x         ޽f�\[����0�';r�f73v8 �K;��
�ȹa�M:l�Gap ;@H˩��iW$UP)�=  �����L6���  Dn�M��h;mS��.��h�l�� svNFv�Mr�"��k�f�`�d�J $� �B         =��js�Vڹ2\m!��kq9D�� *1Q�����l^� =�� ��Ҁ3�8�
  ^�G�  ���h�\��� 	��Δ6�H;�Ҫ���t� ����ã�ss����
H��C�O 4��  h?ɦ)*T   4$��4�  Ob�Q���  ��T���*T���C	4�S�M  f�-(�-b|� 	2�t�@��Q��	!I�9�8B�R�HH���$�HB��@�$�@���3�o�G�*?�e"F)3s�.��Eث��H�H튲��zU&Sx�-s:��KO⺄�ğ��`w�q�z�{,�L��ql�a=H?�,M�6��D���\f������OtĻ��"�u
�`����鮌L����lL�_M�~
Nڇn�麰�6n�R{p���^vռՔ���>����F��
Oݗx�,��N몋7'pY6f���E:�q�������v�����5v�9�4`{r���=+�mH���ݙ���\Ԝ�]5�5�4���j��7b�5[zѯup��yۜ�������p��8g�4z�C�}�m�AM��gp�����4c�(~�C�9q�k�i�Rڒ$꽶�M��V୬�'5(KFr�֎��N���繿�
K"���A�YZ�t·��μ�0�N�ou��*@q=�.nTz 9�h�S����{�U��VBs�W��"[�Ք�k���Z����f�n�o��Cܴ�wb[�� ��ŤM��خR�#sZxV!�p�j�*C���8�f^�ګo%y�u����t�뫺��T�qU;�rbb�-�dv�tW�j�Ἂ��uoL�{Yfb<�R��Ҏ���;h��Rf�&.��m�;�Mr��.��	�U֖�8^��4I���N>�lӯVγ-�[��B�<��7f�rŽ�lv���$mx�v�]���8g���C�;�+�\�t���I�QIT��;�w�ހ2S ;p�u����nY1TZ�����+��"��f �~U�2�|��	.
�b'�m�X�-Նs!�˞��۸&�
�uY��nQ+=�<S�Й���Z̓�ON��yC*��������7]�Vn��h��`z1&��",3��H&�������imjc4���'�K�DZ{ە��wh�cE=s!�1�w]B+��<�1��rf��q�Ib�QT+�@<պ�h�^��V&*'"豮���6���N]�{B�J�v;2�up��
�k����f�J\��qk[׌wc�m}��Taka4�0e�wk[)��v�L�r��Ouk����R��3)�;qp�o	�7][J٨s�nNU-�Ԗ6i�ܼ�qݹ2o3�ݻè�֕�5Bٻ�e0�/vj���<�gq��\�.j�{����X0^�hԵN8�`��ŝq��$�m�Q���_��@׽���&؜��>:��
���7�H@N�����tU7����٤lӮ5_wX��x0��M�bK�xS��t��#�8P���Y�V����Q�q��TK��`/P�{wi���,���+�2"�C@��n=�p��i�Ju.�Ӈ�"f��s5=�r�v�|8c=�W^]�o6����p8f�,q|'9�6.!x�%f�u�,ٽtі&Q�qvZ!��6&��W�1%�Ld�ջ0=�UI�.r\9M��Ж�E� �0�OsQ��͏��w7f=v���N�m� ��C�
c����.�����BӺ�:���u�{����N���OM��.iE.nU,�4���Z�A6Hi���p��h��ۼ6��0lҩjNǉ�Fj���M㗈��&[���2����{#���-���t���� hf��k�=�wvL\i燣'�U㵥���Z�{��nN�F��:R嬦?�S�~syw�ݽ-�B���O�7l!�����T�r٢Q��2����{((l��\QՎ��T�,U���;�J4�֭�9V��
�S�Ǣ���9i�[�x L�&]�A�t̙�Er��G&q�1�r���f���q��=�76�8憆�{�qp<�<�U�_j!����?�3(�$ҿ3{6�������c��at3�*%=�u�5�H�ǮܛPO���!d�HMl�T�͌�ha��vF��((���y�{2��zY{|��.8��U8bER�	��j
��������6��3x��!�?Ρ�5���s�tk �&<�3Ayxm�,4-�UۧZ�^�ݛ�gV�Y,�0v��c��3�=�m^
�;���r�n�WG�{G��%N�q℞�n��䐁��� J�7��S^��ݢk�kB+�#O�+l�%;�R���_7p%�<J��l
j-��K�mR�Yӕ��S۠�b�t����eޯ:�� _ҙ�����+��]eB���ͦ<(f�n���D�e���E�r�up����w���u.�=q%9���8����s��(�u 1[q�ل�oz��("�O��K����t]��|{Įa��/���k�H��x� u��qŗo%�#�͗�.nRTV��F�iR��m]q�+X�� ��\y��[��%	��lZ[S��fn�X`�qI=PF��0��;�{wi�ݭ杳�b|��;F,�6;f0�t �L-Vvn�3!�D���7�Թ�#;C#�۳#�L~�_o�G�{b��4-�J���\k^��P��!L��
��9��bZP!H��ٵ�����;��ua����u�oc;۪� �輋P��F�7�79	�$��r��U��r��pm}��2BrwA^��G��T�,�����i��V30�s���F���~��?v-�=�\.�.lH����Yw�&�"p�즣��X���F�Ǡ������X	> 9xbT3�-�&��X��)���yߦ��74;�4Lܐ�r�`�{��lŔc�vo�z��eg�7xbhd6s�M�';7�n��+L#4��ϮZ�� ة�-�z�s�G/y��z�}'M�ٜ���ݭS IwMlܫ��ۜ���s^�àg��`�(4��)N�4X{s�>�/���Ő���B;0����3y.VqX��%�'nHL�s�ݖ�Ûm4+.����L9�U�@��:e-j�����75����R�<�erM�\��]������׹wwD�ʚX]4���v�o��m��B�g$�zΈ�a�?���y�+��-�.Ҟi}��8���Y�-P�;F��rb��KԔT���j���{/w�nͽ�z��o�;��l�!�9� ,��7;R���{�m���z��4��#�T�n��ݺ��7�ó���ZG�c�.��wL7�txr�[��mt�}����Dw,�U+J�)M�%<[qs�N��8K4ܤgl�G[��oQoY�i�N�aC�#m
���s�k��DRn�ӁQ����署8z�c
��6��Ob�b����hM��2l�
�<��/`�FW����,��uԶ��[v���gں���R���sWxv��]�s�ٻv�%�B=Θ���i齑���F�G�&wwqKy2S-@�ٛ�Fp,�`�@Jz���D��F�pW��f���bƊ�9�ch�v:'(�U���C������:�Wf��Ŏ��Vr,>8(o-�y�gd�L�pn[���s���sb��ջ�EC����1�n�aZ�����خ���6Ӳ]�����թ�vuĪ���+�-��w%�+�\-�ы�j� 3��q��8��ƛ���6���n.\�[�jd���L=��lI�K���-��p��l�Q��F���t�Q��C�rX�7�� P��C���3�^VF�ׯFK�����6�C4�pW��]���&��]n!�����%�QYU�`��qf�fjhz�e0��o`a`��,%��D��e�Z�L�.�r���7o�a.�5�9I	�'�z��_c@n�a��̝s��$Bh�L\���u)�����2�%�3�����m��[�u�}Y��j'���k�v��$�s����ǚۆE֬F��������P֒4٫�g.����L�X�&���aI�rֿr��=ji�{g�c��8q�M�W��c\0��"�L`�.k70��Κ7�
��$�b�F�n��YЂ�	�?\f�����������n�&T��n9i�#6*K9�p<n)E�iN8�=�ͱ�Ҏj���f�u����J���;��M��1�����ݜ�0��V�ɀ%���!A��ݜaȍ6�7n#/3t����n����6-d��8i��x�+�#"A��>xSز7>e�ï��4T�]ם�`�h�:GOVv9ʓ�vN��`�#�H5v�_;]}Ѐi# �����
�c�$0�Ysd-wp��.����48���ך Aeh�w��h�ۛS�7�k<���Ѫ:��s{�6�3 8���$mvqG��Mn�wn5��v1�y���a��8ZA�w8g>�ٮ�GWm�Z��.��;�f�����p;�th�0C���=WV�标��X�,XY:S�1{u�n>� m���!�i=*0d�s�6L�k�k	覔���֤���E��{�섹��G\��j�{�܏N�aDb$��=�f�4�;�㔷��m <Ig�ll�7k�ʦ�V+�t+�ga�g-g�ɸ�1�'Ӗ̱C�n��ʼ��Tɪ������U�^�ϳ�V�h�~Y�T3����f�ʯ[�`X�ۈ�^�=��N��ƹֹ�xe�:���+���-��ӂ��(N`xV7�ә�gZ����020�//4��w�=5�tf����Y;��lZY����gϡt�r�ۄ��Q�SS�ǽ�r���ż��'�;�x�]or���[��un%�����K�B�{K<Vud�k����g>3:+8�5��)t�������;��0Gr�  �k]N�G�P�vY;�N��͜���tb�aJ�l��� y��������WE�f�sw5�5����[���!�.&�ܮc&��`W�Z6���*�!*Cj�ӌ	喲�*$����+���XŐ�kܧWwP�z�$��ŴwM�Id�;��6�(�s�W�#�p����)�	�뽋8g9Z�kһ���oT���,�ӭP��f�sf����[�G.�!�W^j�_�qf�w�ٹS��|���jy����ӗ�=L*;$�X���9=�,~0���z4��+��9��I�7�\�l�A�G�Gq�����qԞ��$��nlfo�Ny�In>�� X�C'�ZvE];r���R��a@�����gr5&���o'Dq���"�)A���y�jFk�M�����2M�Л �M�^�]^��HX�Q�.�z%���}�N���w��Iq[�µqz�@z�.?݀,�.6��jt�i]���We�r��&��h
�D�ntڅy6�������όT<1v=�4a��]�]�aH��%T�g%��ۼ"l:m�_N�Z���^�xe���\��u���#���+
��If]F�Y;NR�n.���6�a� �%sb���4������5�׻�C���øP܉�r�t���SC3;{8n��������o=vj��q��v��n^�0X��c��^��R�yw{e�!P�An��M�>�!�ΐ@��r�qɼ�8������{�ۧ�� q�wwr���5f��s����c��)ʞw)�w&�z[��q֡,eL�Xl��h 3{ie�>ޓ-�D	ξ��*�)��vq=Е�;�ۋ�Ð�o����<b���m���P�j���Ļ������u�^/8�������.9��J��$̥W.��F�q���ּ͝8="n��{ǃ܌{�l��T��.���	��|'wr�n@�oA��İ�p�$gXՎn^_+����Ck	&)�{/n���%��jշ*�<�˙p��p`�*���p]=͂3��]�]��+'q�W�i鷸��

$E���Y!H`�WN�3r�L�l�4r��}d��l��C��^vk��T�^�-����� TʠG��9sxM���:`w=:�u��� ��W6�e���`Z�C��ί���Lef�{ab����Q�kG��`��9�j���Pm���gn\$^p�/'�bMųv�Pr�J��ZZ�Ԑi~�"����W��R*`�Ėy�h��F*Ċ�K��p�VvtkEӕi����*!bwqi�Ƙ��k.[�s�^�]�r�ʛ��^�X�u\a,a��	�]�I�����O.o79^�;�;Ǟ�r�Mw^Y-7]��5��s�u~/4=T��Y_&��oq��3��������:�ݱ-��+��lf�.�!4�x0ӊa���]�[�ۤ�ǧo~���l�H�[��BM�6T��t�}dW�%nQ+�j��+�O����v<;WiǺ�M�Jb����x��7���3����w�S�U6��F��R�;�Ѷ~i�A5��V轫xhY�4����O+{1���1`���[	zk:d�g~�I���&u�m�=g:v�*h
�żɐ�1�L+/q��B'�.h�S;����;�:sztt��u
9�&�;zS�L�'�_跳� .�����x�{C�s�ʓ}H:X�ҸF�[w1������U��E�ۍ�u��*曻2���9���Q���g���WV3�^�Sn#�ݯ�g�ܼmX�9Jx���f����7�Z���%��m�p����7�nwS)7FLQT��� G�B$]�}���נ����y��&T�:��ќ��z��|m#q���R���k��v��:v�������gpIv��͖�m�&'���5�l˜X���yw0��叡ւ�f��n���WU8���G�'��?���gH=#k�&wi�{�^w7�}�{�����HE! Y`, �{�!�H(��@R �T�,�A@"�`�H���H)	"� $�d��B VI�� V
���TAd��H� �`BE�Y
�"���E� )E@�E 0$� F�$%d	) "�@$�RH�+B,�a	 V@
��BE�� "���Aa	+	 �I(��,BII+!�%I!R�����IBV IXIX@�dY H�	�,�H(H�B) (@,� I!P��� ���BE �@�*@�@�d�
HH�����@$$?�	!{��t��?�W����;d�Ç�h^ʜ93�x{{۰�93�o����2�'ZX�\K�!ܸ���躬��N9�w&�T㚠����7&���\�h[n�F(�L�~���V�B��vW�dU��5����#4D�-�1�۸	�X��`����.s)Qj�=c�޼�n	���Q���{4�rN�'j������~���uڢ��3����ۣ9���Y�NL�S��[��nf���9=�ҞC^�S��Ʉkr�&�٭`�čmx+�Z�v���=���>WF{�n���ק�>����`L*���6�.�x�0�*n2�I�5�Enպu8.�
��S�C,�S�Tܤ����Nc%D�]kȻ��SxA�
�51tנ^n�݉�/�y�Av���V�q}��'rG�*�uR�C�|�>���<�_uCu2�f���xJ��x�=g{�Κ�4{��9�N=���e00�ܢp��������=>���\5�3ܷ=1_L��V��w��;\�nJ�}�Z�����ޕ�H5P��4x��PS�\r������b*��(N-
D'�P���iƂ}Y�vucT1n����f�v���CgpSOh�u�L���P��)�H؉���cjLR{r�O6e����1b���]����!fpOy������`k_�0N k<&�l�)�9���I�ޞ�Âok�N�^�+|W�?y�m�z���!�/x/.�*�m�X��^��f�e�<�K�D�;�E~��8��'��zq(#px�
�O�{˅�9��|��K�Wl��I>˭��$�K����S�W�n�o-� ����o^��d�J֒cV�7����Y��z�ɶ��i'���+�'�� ���3n�#��Y˩�z�kq�r��}F>ELs�� ��?>��j��ݯݝ욳��Z��(}�ֿeA`����/�������gI�:1N{���F�W�f��P�ÕQn"�:.%C�$1h��x*�m�pK!��+��a1;����X�Џ=�ڢ��1��閎�;n3|̶^�|�R�t��Yub�� �� �9�=��T�ex�O{U�[���ԹޣF#���=��ot/�Ӿ��yA�ݚg�*;��Ւq_�,uS�)H�+.� %�z���<����F��Ӕ8�����OJ/r�7�3�^�=����L�,���i��]�ٍ{�}&�T7�p{{�٤�-b�wr{Ϸm4-�]�&�����`��`��ѳ:��ZAkm谽��1X���ko�yxtźގpC��D>9�xK|��)�X�U��nQ.�N^K��7jv�=6�D���u���������}2�����gsY�jP�O�dy=�(h}�xL�m̈�%4�{Ĺ��Ϟ�˲*/B��u8�A��Z���p�"�.�ne����i_�hij��;���az�6�a�k(�@W�.�t{f�.�sr��������_��vt�=�*E��K�e��r���&�|��Q�+�BIJ�%��:� ��_{<=�&�rxNt��_��~tN;�oA.Ǹ���<��ؕ����{�t6��dG�v%(I/{�T[i��}�v|����6ӛ�C}�O{�ho�ǒ���v%��Q�k;���<��S����l���`�称�c�y�.#{�7�{�J���f�$���pg��#��SM���7=wzk�_���|�y�S7�q��.�E>���V�kG�'a��,N�3�����q{����U�@�
C�������1�a�4�#;��tf�_'}�gG#����^A��THd1�D�TM�>r�J9up��È�dO)e3m�z���/#{ݵ������Ф��uqQ��D�l8�%�+�>����ӭ��i7�~����þ��o<N9�z��x!�	�G���
�F�{��iop�tM�`l>plc�М��R4mm7`"����u�2X�W�X�DU��9l�oĢv�n ���d�%��]㾹�7x�D�C��]�2�ԕ�u�%��'A�1�[��[fq�T\t���+��m]'��*C��;�<����T�q��4n��u��Q�unө�B���@�=�7�����[e�9�&=�q��<Z~��Lu���"��ub������;�׃��c�C������)�}�����| j��F����s0P�Iէ`�-8���E�y����W������G6�/���U;}�ll�vO `�M�׼f���Uç����d>��MC�26ꁽ���-��p^��y��W*A�r��V�uw�W^r�0�bzog�w��v�}���g��vY�n����������N�0�>�o�أ�̚Ӓ��u&�L��r�A�s^�����`[��G=8S���W9�;m,������Ɔ�;[\�r�Zm�M�8�`�j��S��/cuwd*��29�͛w9��a�rj!<���c���E�\�\�n��ݼ��� ������ܰ��o��;&k�g�Hg�<�	8u��6�l���Iٻ��y��~R��p�_��z�r��y>��g-�gCŊ��G��ƽm	��q[��-Xʠh1�#kN��3�����W�g�Vs���4���F���lg�ֻ$N11���c%ַdݭ�n�����Q�c�ER���cbs(D[��V��r��f�d��JI60!����ehG�=;qvE�smr�}��ڷs�}�Vp̞㪞s�N{�z��<ѯ��תuh��o��ݻ�;��[�v3<��n(�L�r�DD�[����S�*�}��hs����7=�y�a}Mƙ>>��:=���cO��޼R�E~v��Rl��=��ܯ���Z}��=��)^y�	�F�,NJ�!��G;e���b{���;��m@b�ߐ�6��#%_�-�jR��f"��p\�\Gۥ�Tc�ã½i�<n\�����P���O^�7yu[m�
VY%�kڳ�i�p�d�0�jk�1���#�Q��W�f�p%e��ҳc;�ݭῚۈ�4sʴ�s3���S��%�þ���"/m��#���c3[�=���e�H~�;Z�c�?7������z�=�=�#C%���&F%���,�3}75o��^@�а��M�<O�rӷ����<��܇�6�>mwxd�lS��lJ=ї �JV���c^����v݉[�
&�V�;����}|9��\�p?=;�|����ss�����<:��A��8lK9y��lD�NUT"^"dE��Q��h����y|����:Yz��;�J��:_n?*P�wWNг���/ ��,�{�M��ù��Cپ�.ѳ����%�EUQ�����h�a�9V	�l�j������-]���Tp���^Lޅ��c�&0%�_bR�^���'c��/&�ȑT��Gvb�h���<��A��Z�\�O�T�i��/q���-�bl�[�!+����] �c��'1�U�ݽ����,���BB"d1R.؊b A�ϧ,a4��T�7�M��f�{���]&>m ��k���>��ع������vzS���-��G�������5q�>���RX(���#ad�-�*v^��A�Q�s],�x?Q��k��J%��}a�����$�Ww#)eL��e��{���/���a�	��>9����϶/"{ü'��u:��8��'so��n�������q5�I��mF�-O^�r(�ddd���\\/==�͋S�P�{U��Djy�=Ӡ�x*� ߻�A�l��I{���fD�Oo/5x�Fɜt O�&��$����y��h��v���{Y��a��5�pN�sǞ��9V>���K�7�8N+dB�x쉭�[J&qm�х$�p�:њtOd<��;�l��P�Bm8e]�%;�f���]�2��H��=_Wg�Ǻ}������<��÷�{+w�����jB�{L�_r���k;֪}�A��۸��'{]��-�9x���W;�w����D���w!X�پ�㻞�7�K��J
�Y����W�0����� �R;��pe�h�p&bv�z9E󳡸9էN�=��nq�r$i�5�ެ�h��ѡ����{f���{x��t�L'�A�^3-
FN�=��	��U�\�q�Z�����c�5�3;A��B;�BĦ�,��U�������2X0����Z���eY��Ӹq������� �ޡi�P�H^�$y�k�7�������f	���㷖�5.��.5��w��sw�4���U�ɗ+.~�ly�=���w��9�&6��܊�{�iU�����g��ɻ�w�Ft����ۀ���ן%�u5�{Ӹ{�1��7��t��l���p{L�yk�+�F;�,JOo��
`�sۚ/�0S�e��7�Ap�%��ݥX[�c�+�ˣ����s�>vI�"w��\�(�J���D��{�'��G,�=�'���N�׾&#�{.�z��޵6_f���Vw_5�Cx���SW�*R/=�{'��l+R�OP'���]2eD@����PFB�-it'��r��i�x���e<Q;1k��zvm�Vg!n���e0����夽�T���XW���}�n��~�g�#N��y@د- {'%����í��sxYϷ��1�@����������<~��mu#2�b�|����|��_׹�~������ԡ�6:p�ns�g�_V�ػ�]|.�?��9���מ��{����t�y��4D;+y���w��V�'���f]����?v��>�>^~�1�Ӳ��Az�][�i�=�˟M�;fU�|NB� /ɿ�\��:���/�,�ޑլ���5��襪�)a�dF�-\�b�FZ�f�;x@�i�q�����DD�4�+�f�f\k
z�Y��#2�p�c+v�o{����B���o3ڹ���{�$/_���l>2K��}p����t���[�����~�jRf��P�@õC7���Vj�{�{�-8�d�BdK4h幂	�1�UNN����=�3��}�r4�f��4�	��� q`��hz�=C-�Z�ڰ��ɯ;/�5����~��h=�����4�!YHi�BDϱ�s�R���zLO�����b?hi�iG)�� 'Y�Y��zC}݉a��D<�-��@�L�1�:.��C��L��y�ʎӲbЪ(��LH�{tWr8�2v�!/{؉V��|��D����t�%�|��G�H���܃R�=׀w��ec��pM\�>���{����;sG�{"���-]ϳ���u<���7�� �gf��~^�!�7OZww;u��{R�/��3�=����h]:$��y/��&���%�}�.���������_�Z��ea7h*����O&��%�Ǟ���{��Z_��R;;j��MOl��vS��}��j�=�H�N����w6A1�C��fs�u���l<�/���٣�|��z�\���>��㮝�����U`
	��;���'��fmN�Q���u�g�׻�';K�oa֟�;��պ��_O��5�����w�O�Y�΃K>6+�ie����n��	�OS>CYy����q�1�^������#2gF�R�Pы�h:ٞC�{�;��ݳ��oI����x�椋�T��Q���Q�)3<�	4?g������������9g~xߞ���M"��D9(�sc��p��bBE��ۀ�;�W�Z�Qg]*�x��w�w[Eu��>n��>sO2��r��O%68����6u����Q���.�樷��ӽ�Ճ����>[���v���\h)�0��X�v�5�(��ҙ�r���Ӊ@O��ɟ�g���ˑTl�j�<�-E/j�S��vNۨ�H>��u{:=�1���'����:�j�v�\�Mb��ҏ����vl}3|tT�	��r�ې�//C����7=�nH�o,�tN/jպ�P�E{�=g�;��}�������3<�w��	��^�L>1{�.{r��&�nbD�;Zt^���u$CB.DcJ:�nq�=�I�'��t��t�����/3Z`�^sU���;��>�{<��]]�u��+�}�,Q; y0`�=潑��҇�x?�s{�Ql���J��/SA�qNN"&�PA��Q`��W-��Wg�u*��#o(��r7+�f����e��p�	U���2.m�30[�6cJ�IE�X#w��Ϣ&���{�C�=��鱂0i7T�6�;�z��B���]�Q��2=o=����n��v�9O-��r�.\کy�:�e���'v���M���1���==_�o�j�$��N����5��%T�f�u��`�e*��O$����ͨ��~���܎��7�x&k���E
Z�Y���@�,�/U�
�ʃ4ќ|�`��b�M�q٧V�0S�	i�]9]>�xe�]���{Y���x�9OmY�cC��N�D��߸�=�n��e�7S��lط��wEIm[�N[����t��]+�7�����!�=�L��3w��r�}[y�#=4����o����{Q�lqcV;H�i�o�������>=�;��P���Åsל�{�m��q�3t���
�C���^�9t�/qH�0�B�|�̢!��y7���1N^ܝ�~*��6b�?vq�;D��F�u
� ^�љ��oP/��}��l�w����$ ?+���y뽁ޞ��h������
��v[�d-n�8TkA�}A�{��{}�3�	���ʹ�&���G*�*�Ra�mM�ͨ~�ݱo��<y�<}��ϝI龅��V�M�"��`����i�3�"�'o�;t5`�W�e��������xx{���������\]����'����谕�sɮ���q�;�:�r^�n�%�¹�O��<͍��ǮH	��@($��n��63v��7f\Gnnt��]��,�/n��7G:W=��^�O6�5�����W���g�îe�Ia�督�Ls�:�K��ٛ���u�k�[OQ�wnX^�h�\���cg\�Қ�u��mێ^���X�ٻoWm�/v�W�sꓭ۫���.R�s�6N�t��quK�mݠ�<:Y�l����n(8��g��� �<��K�F�l��:Ï���{�q��C��t�Z����Ϝ��1��v�\pެl�.��v&���:;S�:ې^���wF�pړ�8D�yB#Ƕ�u�m>�y��ݮgq����m����v&2q{T�xA��<�s�n�Η���i�	���7\�Y�pOB;�eغ�;ug��睋�@�Mn���9��*�I����6	��7��]On�ZwLq��q]ix�ո��=i�ܧDdn��;rc�u�=�51�[�ֹ�<bz��z������I��z�pl����k�&嫭�o"�y��ݶ�[��;����;�n�=���I��3B݌�(o�cymĜ��{[��;bVy,�n$�=r�5�3����+m�����u\;��c*n�c��v�j���dm�u�+�OmW��Mm۱��爼k$^۳��٠�<��N*\����!۵��v�8X^��!�݃F��P�=�����]�9��vL]j'	6�z���GX;ln����f6�T��f�X)��&�A6ܵΞ9�wOOe7�l�!���C��\�3XN@���QaՖr�X��C�]��c��ݚ�@Y#��@��P"���x����;)�t;���wj����:��\�՞��&�n'�xv�
�aǳ��<l�(��7�;�܋�b�0ð���^˃g�s�۱�k�<�r�����w=��-m���ͺM�i��k#]ŵ��G7l��Fę�(;`�+{vU��J=�¡���綺��ڙ���A�c���v�M�l�z���P��,u2v8�.f���l���r���;��7MѶ��[ٍ�$W^�v�yΛ�96�cM$����� p[�Z����k� ��R�g�81mB��+َܘI�4I�q�x%���{5-�K��ZҶ�۞SLr��l�z�{vۯ[�rc�81�u��8k�7j�9җ��:1���γ�S�s�Vz�mB#���n�����b��cGF^�OP/e�r:^��p&�����s��yRn8$d3�N�*�S�[e�����6�w�H��e-;�7[��z���>�ݡw]�vpp{r]ڣ�k]��7Y{9��_m��뎳����;nM�sǵ�Km�c���cg��j�B����9ݺ����Gn݋���ۣ]H�q�k Hs���pv�:+s监���y��;�Ju㰙�����uY��۩<��\�Ԝ��3��N�NnI�ĮNy�{g��p����'��t'd�;��h��s[շ6w4%�`�[����^Giv,����r78��{rn�k�t�vتS]���/0�J���6 h���y�����r�pr��nz�'��Ʀ���w���i�D�t&;lo������ �i���Y�7Pq=�/I�;t�뷕��v�mA��5�(Qc���S�v��tNmqn�7d�<��p�m������ں7lr�Z��p�����κ�3eIC�5�+0��=q��	Dx�6įN#u�Q���L{Zī��W�aԙ;��:���e�l�݆G���N�<����Y.t�\/M�����K�cZ��^p�^
�[צ�:��:K����pBxܚvۮ7]�
I�keuPV��.2Й���+����xN^M@q��6�콣=+θ�2,y��;�Ƹs]���3�h��`]u//�������`��PqI���� =���1���Dg=uq"j��䂚�!�-n�����G
{8����.�؇��+'<��[�]�`7Uڸz�����	����y�לm�s:�l�z�KR��z��l�J�c����c���.ݮz�����/5^F�vhx��md��g*�����:9W��+F��6���.ݱ<FPx64�E<'mnU�{umQ�2l"8��J��#tv��P���4��-�c��u�A�H���v��\�w
���8R2���M�DR��c��Y%NU➻q�M�<t���xŭ�N�ᒮ�]��<Z�ُ%�W��=^�H���AǮ#�÷�g{�tC�emu���z�{WT��e5v�=�\Vl�a���Z�1�؍� F�ݸ�SO(a��f��s`x�v��ƶ5Dlq���[��Xsvu�<)n֮�k��s���S�XЦgβ�v�z��S�Y��q��>����zs�ہ�.��yv��8nҫu����;���z��������z8�r��z�t�d��Xw�*1h�	v��t�8ܯ\a�i��Ňs�m��������Gg8mշ�[g���7��6��8c<q�\��OKf`ʸ�x�^���q�x�9��!�\k�{W ��X��	7I.@�K�m��fnu��d�۫t��uBl;��n�c\�ۻY�l�n�<�s<���k:�$źD��9��=gai�v[U�r=N��e��!{m��vm�!�%�[����b�ʭ�t���m���욫���vf�Xq�]�<�c;������0sA��q�m`Gl�ݼ�-/H����G�m�+�x�[Ok���p�v��l<<�+��%l�׶�{C�q��!n����0����=x�)ɹ�^�)�ks�͓0����7V�@`��	G���I���,S��2�v�m���uP��8^9��I�盞`K������e'H�g���ZׇԝSt��ͺg�n8y��f���>�ؤ.@�͕8��v����vtñ�l���F6oܼ�R�q�܆�e[#Ϟ��ZCv�S�ͅ�\cۮ�Mٶ5l�b�v�ګ��ۙ��)��M�t���۷\E�]�7vK�0�ܝ�\;���A�ͮ�l�Y/n���ũy���9���L4fֹ����qʻ�d�U��Я�6(���x_�08x4\��"�e{[�،�x�u�Ϋ��pt=�#�������Q۝�m]oZzK��d���ܓ�u����ʧr��y�N��2v�7C��M�Uӎ�۱��g��c�s��q�sv���ۛ�pct\vsg��@�ܯ�*m�m�۳pւ�z��8ڝ�;k8�γx)ً����Y�� ��Ѵ��uِ� �x�����<m�����O1�T[��y����C���M��rbwf�=�v�ϰzz�.׎���yx]�^�v%�i�pk�.�������<�â�{u��u#�0�l�M۔�m�m��Z1'�'Z����av�s�1���v�i^ۛ�M^Cf��$��ڽ �//m�m�D�� �h���Ix;�n�����:q�]����nP��ϴ���د[vڭ)m�<1i���Zv;Y��l�)3�nN����v�ɱ�9���v��[�\��Q��9t[�^��,c9�۶��0Zط���s��h������]t���k5�E�;��<�n�j�u�����rleNXϰ�<2P�'mmd�x3{y��Y��y�kns��N��v�PM��Ǟ�u�$���vmq��˞�-��nٽ\�EϷ8�\#Žd-X�n��l�ۖ��V�c�uĴ�κ
+%{x���i�7m�o��l��6`��y����v�Q�gw.����:�G63q>ۧ�.��]N�Z�PXkm�����!��E�����a��c��ݻb���ں�7O�\��pm�m��Cx}��+&��]X���g���x�������.zؕ�n�qցpqA��NC�t6���6��#�-"\v's����q<�vѫs��tv�K�����\�{9�N�0i��ܜ�v@�����V����\:�]�n�fϳ�q�v���;�h籝�:��-�ҝ��]Ѽ��/]K�r��wH��[��OW\ΐ��c�$���َ�i�nj��1�鳺�3Ɏr��8�M�=�`3�,w/��m�h� ��q��WRW&e��a�k�v�鋞-g^�BXM��˴��9���
��ϗ�q�tc=ѻn'�ܖMlQf�����Y��lx�9��s;����&rv��u�{<��&�h�9c�k��nM;�ֲ8��f�b�86�pq3�Ӟp.�=v��/d��dױ�;V̅nH��t���G=rgv�6Ij�����OO>̞�[]���󹝸嶛7K����[�����׶;���*�z�#f��k�6nH�0���%�ɓ�^6����{n�(��/s����
�ap�vՇk��9�tv.g۫�+��ۋ���ZSg��cknݭq��T���>u؍`�lO��X8zr�e6w̻<s��6�>�Ѷ�������y�n��-��we�w=f��j�k]n�U�;O��kۋ�G"1����,��ezs�q];�G���ׁ��m��js<�J����r�/<��KI���f6�Z����ձ�;i�������	�LQaku]3N�����#p����ޭc�y�\Rռ�^Ât;�<��]P��.�'z�\V7	Wn���m����>5��Ռ�m:��zy��tk=Z�v-�i�]M��[qӺ�]�n"HBȅG9p�'WO=v�g��s�'cp�c���Y��*�
�P�u�J�{-y��0��l��=�k�洍Q�N�B7n�rt/0���3и}���ٍ����Y<s�sr��v����FӋq���7VsA`�Z�48�\�ˠ9,9��;7Z
�N�.�;^�&w3�]\�rGV��4�ɦ�Lg���͢��՟����-��؈�V�Ѷ��F
�T[U������X����j?�X�j�ָ�G(����+X+�\h�1�(�ڵ�B�-k-h�X��P��Wb��UJ"UDJ�,�e�VPel�R�UD�R�-+T�娋�--�6���Z�na��KDZR��U���%���k*дQj�h�Z�J�����%m��j�E.8�s����R�V��n5ƥ+k*��kDR��l�
Z,�+�-�
�Jƶ�Eh�Vƴ��h�h���,jƋ��iL�b�V�J��-�E��X�[T��m��E�҉l��Kim�`�R���jT[JQXҸՎ5����Q��+iE�E��j4iemiJ��kh-jTm-�YK�l�e���k֭�j"�j���Q��S-q�6�\ƫ*�+kim�kX�m�IiV�h�n4pe�U��-�B�h�ԣ���Uh�յ��Dj-,m2��H����W
��Ѭ�HE��\�Fa�ǜ�Y�MR�Tȍ2Q��дTˡ�����
'k�{���|�o��Ϭ��pp�8���m�mb^���n�[+[n��YԽ��ŝ�|E�r�W0�m1쯷c;Pg���N3�r�c��Ѧ��t.���Л���i�݋Nj���r��'n;��l7\vϑ.�s��7W<�u:��,�S!�����]�o��s7\��v�8ym�dy�gw[vy��2�m�|Q�Wq�i3�˷Qe-�r ��v���Ў^�[���6�����g�m��G��l�l�>w�v��ְ�v��zv0��[G;B�1�!�#$p�n�K���l�ճ��7gx�n�wm�չ����Ǜ��S��:�y�n#�χֵ�N[��ɼ8�y�fOF���m�k�� ���@z	�����f�ͱu������zt;�9S��g����im!�^�m��غ�[���� !�lۭ\ݵ�K�"ے�7��Kc��;���v�us�89i y2p�<�=f��g�nLn�ػv��m�:���Fw�uu�n��>c����/2�s����]��t%���n%�������b}v�|�E���4l�`�ۖ㝅�{6��M�W�\�ʯ+�莩��9�������L�<�Ay���h�糠:-%7B���ݷF/8Zy�nv�;��˯������6�۲�]�W�qix�*�W�F���!�����6�_+��f{���ڏ8�vQ:�]��ʰn�6���s<Þ��ۻy��ǗN��3��-=���:�@q������\vǁx����Rs�z�A�\'�/�j��sI��L�a����)@��nz;c����(�p��k�Vx�V��A��u�ލ���v�Yy���6<�>;���GM�s �����Eu�m�`E�"I4�2f��-m�G;<7�����c�Ɏ�H��\=zFzI+[q�4/����������yw��l��ɶN��vlC9���<�nq�S��Ϝ�=�d\�g�țv�vr�gnv������S�wr�v}��v3��d;;�s�Lp�s�쁱��9;o)���㳶y�eP���<�m��;�|aϷ>3��n�&��nݻ���J���l!�3����Î{s����s�n]���<@�n!8���vg~��q	�n	_�Uoj�$�{B�ju�DRtn.^�}���U݂;3����d��D�B"|�׌��R[:c�^���g7`�w3��$�����i��@�z܍(q�.#��ۚze)D�&bݨ}�`���$�;���uk$��� ���hI5�ل
�
�dH�_M��_OA8w�m�w�V	�.�(u���Vҋs��n�X��~д����E<�U/� z���cBHПmk��K2�� ��oz��}C�37ܞ/��jT�d����]���չZ�W���4H]v-���x����߼��Ɂ"RH���w���=�$�I�{�)�h:�zY���s�0Y��E�w%I�0%aH� ݷ����Yr���X�{�ʫ�-?�Ҏ
}��1^k�-~�H�=%�M���)�����žIܦ���Npy�2��7a�U�v+D,�s��'���دHm�]��uө�W�`�u�>�nI�`Mxц�O��]�>:�Ȩ�����ur�˿H8gv��s{�~�XQ:�An�`���>�Ê}�"9��̺�I$��w��	 �e[����Te7ă�6�����	R$B�dH��-�0e�~�^��O�s�WP3��go]�Hʷ�`�����C�8PS�l�v�X콵��a��==�p�:�\���&y�k��Hh~��;�iD��E{���  u�]�H$�}vz0>�ir��uS�L vn��&D8�
eH����'�]����$�H�z��9V���36�<��1�RC��J�
`Jbi��C��V	l4�x�����(�uj�o�-�5��?N���@6]�X�k}I��9���zv�͉� �9{w���xӋ{7y-�� wn�� ��}vI�����Q>�3F�s�]Bَ�z�:"�� �c�|	�:g�-���j!_N�54���7��)D�&bݧ=�`|ݡ&���w���>B�u�$��}�/�i��٫�-�8������>�P��D��"${5.��cpV�nn���T�/^n1���l��~���Z�,Y��M��߹�  ?R�����v��yvO���VHw9
:����)���e�?`qw�}>o�(3w���n_u�$�3�R	�eWOGTE���L���
L�	�۷~���$�r\���{3k���K�}v	� ��|.9ؕ%)�(
Eٻo�\���+ne;����$��wb��'y�_\p=�r�� R30W�=Ѩ�b�d<�&!��k;5���Ζ%��J[|}4l��}�{U�}��n�E��{����U7Y[y�(��/����'�!DD� �F9��_=v�2p^�f��x��ܫ'Ğ3�BA$k{�~7��2�@5׿��'m��=H8d���v�qю�qɠ�c�4�͝-�5��./����Ҟ m�/VSˮgv��A>���0f��w9ݓ�|p�lQ���1�0d�dH��wb�5�Z�I������ �=�@���vH:Nv�gb�)�w�v�!C���J)���e�C ���^���&�[F���H:gv���\	��J�Rd M۾�/��q�A���I�$���b�̷�p:�	�n��'N��$�v���� LaH�T�Pe��8q><O
n����!-yI/;]�$3/z��\�m�6jgV����}�z��΅�B�Vg�d�q����{�V�}y�xt=��m�A��fv,��L�$`ٹ��#q�u�׎�o�y�^�;ȍˌmT<g%�7���@�����<g��BV��	�ISE���y�����M��yդ�G��%n�y2���n�v�墔�ݸ.s��,������xm�/:b��t\cqQ6�uJG��x1D��9�qi��b�^�\�$��tvӍ�=�6�<���1���v�F��giF�5��D&�4A�6�T�}�j�E��w3;��_E�u,ݑ�m<�[	Tp��٧؉
lzbL$��i��"I��<���'[�~�H9��V
��z�����2u�
�>��wc�-�D�#%D�&bը}�~��c3)e�
����A�]X$�;���~o��6��U'b�^�)� �#"Ex�����A���	���5���UY��u~$�fm��'�jiߴ 5:����|����Kp�lb�m�� u��$i����=��.hZ�Y[�U�jT̨ȑ�I(�ݫ�|HO^ƪK'�%Eu�N�� �<��(��S��V���.n����W��w<�X'���Ӽrq���n5<N�B��f�{��(B�JR7����ψy���	�ױ^e��1��Bμ�$�ξ�`��6aO�(��D�G���F�`�����agLMQɯ�V��`��}W����, ��U�;n<��t���%���9�\�Y���k�=��!{CCΉ��ψ>��v,N�����}��E��%�<��ԑA[����`�|x��	Iܜ��5,�ା�$�m��'O^�YF�D��T�"E���8y�v�Wn@�v�I>��b�$oc덋n�Ɛ�=�Ŏ��Q�D��&f".�{RA�����s��2O�1��>$v���oc�lWL�����x��{�rj���Mu t'[�/F����L�V�/:����ߟ����������W�,t�ؠI;����;JjH�[��v	���hM�<0�
H(ȫ7m��ɱ]��cFo,{^��o`W���V9Cr�v�0������l(Q")�h��A��5ۊ(;�}��*��nM��Fs"�M3�&��{�U����f;���;u�b�!�Vm���:�k�_>�}�\z}[��w|ò�c�� �t��
�>�{�d����̣%D�Bb$�]�SM�7�t$���$��θ�hc<[p	4i�	#���@Ĵ��g`�˛����C�m幤����'޿7� -�6!T�u����<3@�/�(8󈁰.�I���h�����@x���ֱ�밼t?����O����w�����-��� ~�ϛ���&3(H>���]��&Dh�FFbB$V��X�j��dܚ��lP��_7��l��zC�~�}�d�fi@�L�����}VI}���$�Qݎ�n6���s�a�On��n�]����a���HhҸp�y���_ڶX 3M��$���`�H:{7EGJ�"�:�DGn�����#f`�Y)�$V�O�;1ٓ.�,D���l\�((�OpN�jF���S8+�����խ��U4�)_l'Ѷ����u�q3(�Q![�7���60~/b��ͪ; A{k��$��v}��jC��MU�7nă/��FUHe�ї7u�l=k7�ܜ�On�yi��2)S�����3�K%J���O ��s� G��f0M��Tk�C9w�����<y��4��	�^|;ҡ���:n���ȿ�u���_��`��t�mxH$5����{�Jt����L�3&bB$WN�]�O��͡$h�Xr�&f:�vVh ���I��ٵ'��B�e$�&E�7m��h̉wWR��l��&����H�unlW�#y�\W���qh"8DKv/з�!�}0�%JF�K�$��b���'yS��>$��ŀH,���F��vl_Y�S��4�;���Gl��n�*���v�?���k;��#��؞'��)���'��x�.��=�=(���'Uq@�f���nx�+��=c�HQ"$(��֕Ji5)��w�]���s4�nIL��v�{j�k	<�{�<�qt��>�'�7T�Ѯ�snX�ڎs/b�m�eնڹg��	�8L������݁\�����3@�����q�]��5V{�[�{�3p�[ܻ�݇i���q^1��6{ud�H�n�.뮺�ьq�mr�E`�<�x��WL@n�nکcS�yS���j��cC�+1�H�n���8Ƥ��W�9��sy7$�<W�"�}2��`����yv �^� �/�~l}�������I�<�.�$��hI�.L�HJR�"��s�3H�	�쌛�`5�~쿀�.�k{�d���)79~'*r�L2T]�6�(w^����(/�m[��/j�� �Yw8���`no,���Ӏ-D`�ʫ��c�k%�^�@,�� {���'7w�R�v�IU�T�#oP����I2�L�F���>� ��uՀN���cњ�n+ĂC�޻$��޻u:�͙�-ӨA9q.f�>�P�#�8k�
��'7ɤ�ݨ'�����2q�v�~{���J��0"$I����	/^��O�^�U���'���<q�H ��޻ ���9�F�HbԱ�|�\��_�Is�7�x%���w��#Y�q,e�U���@��g$����o]�(#����p(�f�[�Tle�#��k\j+='�`z�� ̮ߛ��sW"Y������z�G)%�J��>����{{�W�I ��=xວ�	&��]��̮ߛ�䦑�biѩ w����~����=���gt`_���  ��&�g���p,�O�[sw��R�' [(�6gz������#Kc�:W���W�œ�����N�܆����"� i��}K\����N�=kj�Il8)���OlV=;g���B��LI22��G8��Y�yά�O����'8���Dd�*�Z���n�A�ޱ8��'�
dL�Q:�BH)��>�h�㎲���滰I ����R�f���	u���F
�"JIc�oϨ���z��?�3/��>S�3�\�S�ӵ���ۀ�J���$�����!ʁO.�z)'�w[W��˺��+\9U!j�W[E6��a�O{O���^���a{CE�z�^���4g�XrqC�[=/E���͛�bZ�+�*�jX����=�'@�r8=;��a�~��|��zj����5�`:�=p{m�l�}�o2ZQ���f�U��7\4��n9Ǽ���'y��^��<F�x�:w{�0� �_�/���+<�W�Ρ�/�j�.m��i]L*��T%��
�r��]��=�������t�c6?G7�z�D[�1����������z��%Y�֦�%�:ӛ�%�ނ�EZrQ��Or �1rjed#s�X2�+h�7W�{so��!P;s�yO^��{��Ԝ w	�S4�3m�\]�|��+�����q_�����t/�\��'�lV=x�V& Y�r��讍��^|�}�)�]b|�ꉛDŖH���x�2z�zx1:m����^�`��%ub\�疲�[r��I�3-*������:owm���o�;0�y_v>�xQob�Տu�\�ǾWU����8e�K��/����}!�0ɿAfz~��L�U����B��/��0����P<�;6����Ͼ;�8 �_�˵�อ��Ƥ�nn,`1Pؖ���F��=q2��La[W�i\� [�J)3����@.��[�RQr��)�7��n\��7�s~�<6wn����3������êE{%�����P�:(�R�S�g�W�i�L��m��(�J�����ֽi�JTh6�[X��-+e��ケQlq��ՖV�������5)K[P��j��Դb%-ij�J�QƊ�E��)m�.$m¶��e����k�Y���,�KK[R���b�F1U�QJږ1��-�KLZ�[l���s3[��V��A�--��R������k-+Q��R�[Q����)e�����D��c[V�6����KF֕(ѵeQKm\˅+h�V�E�T���S1��e�Z�[R��6��J--�eT��ԭ��R�+Q[F���P����h�kA�am�,�lPXմ�m�QX��TE6��F��D[-m)V�Q��+J�P�m�ce��DVڨ����*��V�-��h��ZU�DkKE-������R���[E�օ�lQ�mh��K�
U�ѬmZ�(�h�[[-�J��J��iT����E�U��Pmz�|ߪ���vH'���د�����)DD�E�V�q�':o8S���U�O� ��lP#7��T���x�� n>۰O\�#~���	 Sc���0޿<}�.��1R���;�]����N�o]���u;�2J�C%�4(p�TKG�wm�����r�e9uӵ���7%�m�\�3���}���F^ eB����݂@#OVׄ�A#w���y�]��8{�T�D�:��2|I�ձJ���A~'���������[��'U$�][����]�^gbŘ町�A#�3&$(�%Ʊ'�=�� ��c��9�y;����p��H$���vNPk�(0T	bfE�Gv\<.��)�	L=�G���`��޲�"T�>�p����_\v>���{������U��.ʉ��7D��Ǎ�qv���3R�W��&�]��J� ���ʓ
�-�	B�5��w�>��ޫ*�gm��*�H'�s[���Iop���mZ�:�`X� st�f@5��.Ml�Yv��>95���vv�9���s���2�6�L�D�*_��jH$o�����`�E<�q�� p�7}R	o[�$y�(B ʅ>"��W�`��zI7)Uќq��Ho�݂A9��� ;�\���Gn����:������2$+�m��|H/;z��|i(�~��/���	-�����/�)�*B��=/a+�3��'>뚬�	'ٝ��H:z�^噂:}V�9k�
T�C�K�ݔ���+"FO7�����ܫ$�����H:z���W��u��N8YrJQ:e�M;�E��)��w�u7�SC�t�#e�P����u�^�0�ُ���`�G� /������Fz6�׎c�Oʼ1n9ܜ�ۑ�Lv0���\v6�	s����1ؖ�M�pv��\�qu�٣���v�;rm�C�m�v� �1E-��k>��6��s����v�v�Ҽ$�����i����.�@��Rڒ�ŭ6pK�<n�(��������+cn4�c�Cu�����[#I=m�����K�溓�{gɃ�L�͸��=��>|�7��oIY,���^cq�Iv�������=��%�����U�|w7z��O�W^�����*1Y��#eW>�$v�6�!��;���"���CA� +�|{̷٢� ����ϙ�ڟ*+k4��m>��&t̋��LyHQ>�]�}vI>:z����Y������;��ZI>�{�d���^Еu��bA		�"B����C��D�s��H�T���$�w�^$�}V�hr�9��(h����,O�T�3 ��h�u� ��9ݡ�v\E3�+*��đ����F�w]�C��9�~=�����8s���{i���K�8;Kag��LQ��g^y�uv������g8z5��Ϸ�v	����'ĝ�}V�i�)Eh��I��k�D*��I��dIJ���{,Y;�Y]E��ν���H��ʩY��jY��z.%�(ȈC��O9/^)j�'8冾�V�)��n�\)�ĞV�#rh:����2i��ĒO'{ ��}v ����D�9�$e�B1�L���eM�,��|I׏�Y$�k+:�<sW�Ig�`Q#w����h�Շ7Ӻ�nu���C6��@2{]I�$-���H���ȷQ[����6g]I�yJ�$&�
�x�����]Ui<�o��T�W� "T
���织Y�J�*��y�� aG�w�f�w1dcD��#a��D��-&�Y}i�
3���8��L;�8�<U��Zp��wY�b}2�I�}�DxKg��6��T�!Xy�{���%�� -�����#�1�1q�D��ót亾�<	��mx��	/|��0����)�$D%&B�f�#�O�m#���O��r쟩}�6߼M,��>�!bJ�XS�>��C�:°�
��[���� "<	��%aߚ��|�,ݯ�g:_*kN�q�.�@��������(ԅ�?y��9�B�B�>���
�.k�qV���&�^E܌�*ޗ4�͜�YLe�*tE[,?�rwNm+�y=XE��B�*��*����S�Κs�K�nifg�c�TK��������4�S������nH,��Ȁ7u��dxჲ����P�	�<�R�ߟ�s�|��7���ĕ
��X}���γ��� �P���>����G� Qk�u�;����7ii�B��~��É���f�f��5R���y�?}��؁YY+,d���t,z����T$D)x=dy��}�u�XVaP>���q'P������ȵ����D*��c�I�PH��=��T��ky��YmS�s�'����V����4�Ns3?D�#`��G�%����s�vz��H(����9�B�B����|��I���B�?E�������{�9���z�R
߿}�Ρ�%aM���MMj�K��6Ã
���v��<��l����BX�4�)�{>�J2�Q*���=�Ԃ��|��^�!�R
{﬉���b�;��y�z�`V�s���Ir�:.�Yy��'u�߶u:�R,d��~y��&б%H,�����{�s���x��
��%O~�ݝI؅d�����]���i���[�MkV��tp�Gç�� ��>pd}���>x�<	 N��8�zR��_�~��N(@�7���,�n�}9�M"7H�}��7]�Or�^�A�7ݚ��{z��oz�%���7�*��WUcPx���I�� �׏��_�n�~�D�mܻ��BI�?�J�C����:�Xw����ύ:�s5�������m%)@������0a����ӽ��~�<
������v%`V�+_���p9�<	�7��^s��#ے`=v����x��B�����͋6��nz݋�ղ���v�`^unmw���߿�q��6x��폒w�~�gS�eJ�_.��g6�IR
y��{�u ���?�>9���!��	�=�ݝH,�ed�+�߾nN&�)��段U��U�xu ���퇾�^(��5Dƨ#*��=�i��
����r���R�#�o������Dx���Ip�c������ 0G��B�O8'�*d���Ci��}�~�6��T�
��>�ݝ�J2�X���w���tw[�Ys��|�蕁Z����~��� ҏ|ﺼ,����ˏ��J�����s=��8�mr����_���t++%ww��q�i
���y��a�|��#ȍ��a�y�q
�Qs^�Y7R�[�rr&�(o;��SZխ�.]6��J��}���`QDx �濨^y�V)�$��X0+u���@�p*Q�����p�:�R
����C�IX~�u�翶_���l;���!K�,^|؟?k�u�������v-�P������i�9I&k�x�Z؉��u*&��j[Z��~��~�ߟ���u�*�lh#	�k!�q�9C�u���/d��qr!�;f|ôa��8�1v��OX�įB���6z�F��;�!Vd�6plv{����zz������=I�����k���g6�O.3��a��j�t4;a�� V�Wc�6v��U^.��C��x���s^�slk��;��n��ɅO��|:��졣qʝ}�bܹ���y>`Cp]�Q�R��ծޥ6#]ʷ-ssq��a8�?��S?�"�ӯ��7��0�������i* ���~�gFu�@��Hno}c�'�Gξ����=}�����n7H6��,?}���p�Tq�Y*B�$��
�"��P�0�������[��w�
�{�����&Щ*$�;��}�8ì*AI`���߶u'D+%Y4}��������]�����6�L׾���iV�Z]�P:��~��ۇ���{��}���x"<	Wsw3�'�F���$` 
����{���R:2T,C�{�Ρ�IXY���Ǧ�:sC��6Ì+˯��gy����.אĞ�RQ
�\矶tgY+*�P/����@�Vk��w�����_�]�9�d�A�HZX{����נ�����gؗ������Rw���gS��d��Mг�Q ����h�y���a�{�70�aXQ�ID������:!Y(ʐ_�y�@����u�߲�������8�7'~�\�Rnd��n:�ܜ�4ˇC�qۊ������n���/����~��6���i�3��a�����y��{��)JB��ٿ��'
��������x�?~���q��J�2T*�����IX_y��_���e�a�u�u���'����Dyc�_��˦!|t���;5�.uC��bMq$R�SL�;ӳ��;n��D+�x�ȧ��������^s�,��<8��k��o�����@?�L9���p�'�*A@�������`V�,k������A�x!rݑ9��T�)�o�]���Ń�Q�Ed��30 +��#Ξ�C� L�d������6r2m
$�X�����ޛ�{|9w�<��?
��%����I؅d�+%e]����m��~����e��V�V��W����?A�Ҫ��N3�,G�	 >�}B��!Z0+Oٿ��$�a��~�p�>���>9���s�8��
}�y�Ρԕ�9��zhӧ4:��Cl9W�^�����T���>�ݝgY3��)�ֵ���T
y�>��P:%`Q��w������B����}��װ$3�;��H���(?M��!Q��etb36��pn2҂e�a�o�ِ�g��q�߿O?g���Z��f}�����:�R:����6q�hQ%B��)��~�����x������7~�B��Y<eH/�~y�8�@ߝ�}+��mˊ�@�t��^|G�o����.; ��t,��P>U�N T����}���td�"�����Dm��\m�d#��!�{���ֲܦ�\�Xu�~�w͇IP�,B���~�gc:�YP(�j4������P���;jD�񽛙y���_����>��璋I9��v������d��U��cLQ����G� $�����<@�+� ��y�� �B��{�u��1��tk&�kX`��,�O~��[����o츚�� �Ag+�����d�IP�+y��g��>�����,�O���ˮ����M2�~����m�5��f��Q��5[xu ����퇣��-@���G���iu�ӝgv4�ޮ��
ӹ߿r��@�beO}��w�����T*�~��H,<���u����7�����eH��Xyr+nحZd���m��ܞ�r��.<�ɞݛ���~��;�����v?���
��l8�i*%�=��}��u���J�O߿{��u+z������.��p=� �H[���w���y�}�q.��m��@� �ﲅ�� |�������cg=�w}�:ɴ*J�IXS��}�!Ԃ��`#w{�G������>�A��o����n���i[�K�]f�n\�tl�蕇���v���?~���*C������|Wջ�N��$x?�'�}���R:�
��߽�gP蒰�뿳�:�[��X���G��@U<��AX[P߂#�@Dya��~�gFu �Q*=��ϸu���'� Q�_:�'���DCkv
?XE��\���C��4E��C�x���{��y/�{���,�}��4�����_�����G\��k�nw�L8�����s���\�?� �?�?�!ia�����Ԃ�1��tk&�kXayN$��~���� VX�Yc%|���p4���s�﻿��IX_��=�:ñ�aXT�=��߶u'P��2����nN	���ϗ���9��?����'�CU�>�{�b���8�e]MnF�km:;9��nv�z������g�gj�~? }��������jB�����}���-�*Ao���r��N]E䞨걩e� I�x�w�>��#�*!���{��tIXY���Ǧ�:sC��6�]ߵ�����T�}��>�����}��Ϲ�Ό�%e@�T
}���p�A`u���s���� �!��_پ�y^G�=<~q���f���s�:������x�YY++%<���DG��dʜ�z���_C�>�+
¤��~���:�Y:2����nN&�)�~��-֖ܹr��%a��v<�g��\�
C�@߿w��v���*A}�����p@�|���^}�Fֻ�uj'}�}��Ȁ�/] aG�t�����Q ̙�H/�~��x0�AID+=��vtgY;���5�{*A@�f��:�Ԭ
5�F�_;��st�il<���:��H l͉�؎ �R���%!_�Y�(�������k��q����O���I�6�<��J�{�������ǚ�yީ�хo{S7FU0�`�+"-��.����!��l]�ԹSe�L�o�S���.	�}����&�o+}���7������V�H;�hyR�u�i�&s�Lb� �}���%�(�㫩=�3����W&>���h~���F�vY1������;���]<ל����`��\y�ջr���9)��Տ<OU:�ڡI�&i���s&֊��rj۝1��}���M�!��grT��F���,NR����|�y�Q�^���=߸~�٪z�խG�o��n۝��|���ø���#᳄}��|�^���KR��sw������y�ۣ�ך��>���a��9�Xy^�Oj��	��}zF����S��k�nO�\�4S���S���b��F���i3�h�t����a�nh�ݱ��-Q5Ox��]c���r�=�jѾ�=`㾋֢Ks����O,����<�.����yw��5p�N|L>�ga�w����o�OZ��f7=�v��I�/���������t�8d��V/xe5/{g�4�~~���!���Ӑ���a�^�����P�y��d�r�2�o'|��5�l��:�*�Vj����S��D
�,SS&�T�̾F�S�U##f�0�������.Lc��ڌ���y� A)x�W�-��eDlE�K[*�jV�ҔF�+ƪ5���6�ʪ5�+lek-�F+-��*X����K�h�EYm-��i[m��B�KZ�TK(�E�5�**��h��Q�X��X�mR�U��J��E�U�(�R�ԪԱAW��YE�e*��F�R���J�-�-��(ԩm�TF�*5KF���6֌kJ��-�j"�E�V�r�6� �V����*0QDZ��Tưpk*X�-�*�+��h�P�F)RZ��Q3+�FE��Z��-*��m�EB��Uj(��5�KJ*��[[Yl�*�AaF%�F)R6�UcV�b�E�����!UY(*�[JKE(�,m-�Bж���e̡��ѭVЭ��UmjXX��mh�h4K*�-J5�Ե�XT����̍-�j��m���)kX�j�le��JĶ���*��E+V�ڡE�Z�*��X[eT�mm���UcR�m*�m��ek@=����~�m�D�����m�W�h����v� �6㱮v��=����\����Anm��9�s�6H�w9^�̨�y:�t{r���uX,c�9N��yLnM����gY��R�����CpS�яK���=J*���qˉm���h�[��n��p7"T1p���s�� ]\��,w9{#&�=�c���m�:��ח�x|x�75�f�V�t�z0��u�����;���ك�Ʈ�	��N�/m�K�;�y�m�7���PvX��ӎojwm,���� �ںN���F^u����Eu!��`瓵eaw�৛l1k�nh���j	�6 -�{JL���δf�q]��8���v�\��]��Nz8�� �+u�H���R=��=���<�MZ�g<�\����Jx�sۭ�:t�s��[<�Ҩ��i���!׶J�[��nCm�[v�n�c�}��=�l�"��E�-�Z��O0��ӝ��v��C7���*nS����\���]0Z^�7\��x˺��vCs��n"�vc���kݻhT�n�Ǉ6���3��cnk�Y��=W`��<����]�[]���q���!�=�/l%G'��
��'w!�����4��5p�ڦ9mY����mk���#�"�Xm���{��6�h,{��ӛ�7[�1'#=>n�g�v�ش���g��7
�T�<�ug��8�����粅�vSyמn]�� n!��ո����<�b77F����^'�l�O]7�sYh�����WOn�����8�91�ǵ��.:�[��6����=�ɲ�ώ����<{>h��/7Zl�3xS�\�=�ع{p��lx{g��]�Ze9�kvz1n����{KGGl�k���¸؁h$�ཹ��N�v���x��u��A�ګ=���z(�Iѻm���/\t�<zwf�u��vz�(�0]��y���R>�.�u#�\ezÞZ�Z�����b�����j�:j��GM.��g-� ��>�U���w����{���q���K��&�C�ۂԱ�W�u�k� A��v��gr:�u�ƽq��V�E.ˤݡ�i��s�o3�tQ�l��PqֻtuP/�[T���v�J�x�^d�Hb����e��ܙ��&9��e�u\�}v�Q�ٽL��Mk�띉�m�-�<�P�0��s��y����y�^9��6��Ú��.G���/��&M2��nKq�˥Èv�79˸@������<�nj�Olrκu�3���?߽�����Mְ���
�������v VR2T��~���Vy���a�°�����|u��Щ4�����ԝ�VJ��Y_���p4���|�3Xj87Z2��#��
�����Dxm���m}A�o �����W��E��߀���@���}��ԂΌ��]��fH�U�gv�в<	�s8A�"H����a��y~߻���B��WÛ���Ͻ�Ȁ�3�����L���}���z����V��_{��p� Ґ���Ͼ�p��i����b`�feD(Q~�G�~�ha�ǯ@3Q���J�{�l�ɴ,IP�J�!���0�a�Dx<��o�G��/�������ʐ_����@�����Z\�r�ѳi���sa�z�RZ �^<}�(?To0n�9���g=��NA�@�����p�;+,d�PC�|��C�J�<�{�4o�{m�D�����Х�j p�����Sl,m6���U�O]nͷ/������Z��{X|0���|�pm ��
��~�ݝgY(ʐP/����:�Ԭ��Y�6V�����u�.��(!������w��
ۇ��ٚ.�.��0���os�G�>�}�}��ъo^*lX�I�шw��)��/�����;ͫU�&��6F��yOyy��'��.��d׳3F8A�v�����w<8�������$��M��~�g�ɴ(��RV}���tV�ID���?�u'D+%Y=�>��'�|�������m�}���a���iռ:�Ԭ=��}�q �;h}�϶s����k�w�a�o��3��i<*T
ʞ���w�����%B��y�Ρԕ�.�<��DDH3 ���g�O�"���"��}��R|�a�߽����H(J�C�X� ���@�<	տ:��>CZ�����=~�> ���kﻸu�`V�e�@�bfTQ^��������O��G��B�}� �8+g{G���+�������,T�O=�϶u �u������ܜM�k�־x��/��o��w��C���U�v�p�Ƹ�v9��:�*���=%�]�j�{vj�����}1����|@�J��{���XjB��y��9�R�![��������O����'~��־��i�9���:�R
@m��a�tVD���DD��#��Yn��|(�"#�ys���'w��x���>��gY+*�P?}�l�bT���_�y�7H4)���ج�O��?�#��x2<	��2 ɫ�ֵ���}�;�Τu�������͜d�$�T������τ}��
]������S:���QGNz�ܫw9�An+�w3�I!՗�\{�{r��潕�%�^����[��u{;���ٮ�o���?�
°�*}��l�N�T��FW���5'�u�艁0BEL�J��߾���G��%���!1��	/OnyU���k�y��7�� T���=��ì@/��������Htd~�{�rr2	���-����7���I���=��X#�~��?C��ٵ�$x ��np�A`u�
���y�9H6������^p�s�S���Q����Za���·�ۢ�{O[m�,v}Eq/A���nw^y�u �����̩0���y=�,���R(�_y�mD�
$�+}�_�>�46�ɇ���#���;gRv!R%_?y��q�5���ѣY�1�6�X{�w��Ԃ����n����-�<C�|?ks�)8�R��'����ì�%eJ���
�+����G��� �*\�L��:ñ�}��t�8��RPB���~�gFu �X�Zw�>�z֨�O�g�����E �?o9��D�e�����ïX�~��tj�ՙPJ� H������7��q(��� c<d��?wG8�P�+���!�x��7�P�<�N�Qʶ��ٛ���8�n����]�I��^on��_a|���/aÉ��񝣯m��ޓ,f����{����O�`�}J���$�$>H,����￷'hofk���5uo�����cԂ�	 ���Y/쏽���9�<8���׿�I�
��������Y�d���
!�y�Ρؒ��y�x}���|�/��,Н�Mh��-;��Y�;��3�<y�p�M�A9�����?z�rݧ���|a�a^_��Ã��!Xy���q��*�_|�ϸu �7��2w��>�����ן}�H<�-���}�p��v{��ؖ�Mk.���N�N��?l�u����k���w>�~�~���M�*J�Ͻ��É�F����8��>�>G�n���ﲲ/�?��?.�R|&�,�k����ѭj�9���8������^�(5!e�{�<�g:R �`W5����v�t����g}����@�������td���
���϶u��)��1���W33F���-�����z��È�@������γ� �~�{���(��(�߶�|��6��#��^��W��`V�4���tj�u�f-��s϶q �����������2m�9���l���_<'R��߿ra��%���:��
�YY(������h�!��|�[ќ ��5M�L/iVv���ע�6��O���
1wxW��!�F�s�9�ʌ>b�'\��Wp�}�5�8�w�ӱ�\<#wA�M���<�@�5�+��8�Z��clֵ���u:뱻�!c�n7n�s/nM#ۣw�wm[9�V�牻Jq��{Z�ض���X◱ǜ���:5u������u�20v�t���S�<( uqbםȏ���]���w=���q��a� ���d��7�n�wS����ɱ���`E nP�ݵq�n헵�)`��<lٻ�vV�u^�nI�-n<��.��n]e��vOF�ѥ-V`��a�Nvu�zȐ��+~��}�5����-�<@��Xs��{��z��H(w�>�Δ���k��~�܁���߷��ٯo�<g�w���p�:�YY*��϶q��,���_ƍ&f��o!�`��_W��<	J��2�>
~��i�$
%@����xu�Vk��������+�x-�wc���TO��σ�p���L[�kYt��@�tI�~��N�VVJ�_o�����B�*IXo�{�3=��������a�°��IS�y��:����+%e_��rpM�S\ׇ�UsF����6�į�}[��җ}���e�?���Q	P7�y��v�����
�w���AK |�F�}���ﱆ����f��Ȉ(�k�l�	+?k�ύ.�31.h�!�a_��?l8�i*%�ﺆ�>�\qUt4ο��� 0B �ﻳ�J��`Q����n���//����Þ>4��fW]�1T�������X��:3�y��iҞ�a�b�17���{]dv�~�w��k����{�n�{��l�t++%e�����8�B�*IXY��~�������[��~��'�{�{ݝI؅H)���|���zo���4ɉ�+i+h~��� p�Dxv����'~3���I��ftK�w����������n��ҧ�v��j�@�P�����s�N��GtP�橸`�s-�tX�������w���l��!m!Z�����wI�
������p�:2VVJ�;�Ѵ&\�ڥ����a�|�=��Ѥ����a���~�8�i* ���}�gY�JʁbT�y��w�{��y�{�� tJ�X����n7H6��������Ԃ����όd�e�
/�aG�����vcbwT��8�J������ɴ*J�V���0�|0�" ���#�;kvk�+�{xi�1����~}�8�@���O��f�kW+�8m ���w��X(�@m�B���W]����$�3��r�
p+*w�~�p�:2VVJ�����Ρ�%a�5ύ7�z{�[w9�3�G҂���OƷ=�-��V�Qٺwl8����[��v����ǟ�m*��F��|¾_<�����T�B���~�p�'FT
��{��8�Ԭsw���eϾ�~`z�w��p4�yHV����� ��=�ȕ"T��*�"�{���ΧD
�2Vl�7�ݯd����l�2m
��RVy��{�u�F ���=��I�B�O<}���7�\M)��G~��KIt���&TH�&& |:�Ԭ9߾�p��R�<��}��B��b$8�k���+��*2��Nڗc�9[{8�O\Zn�9�Q�&jx?}�)��&g��Ţ,O}�ʹ��v���,+�ՕQ�o���{��_�$~(�YS�~��p�:�R
!�=��gP�IX>u�_ƍ&f�\-�6Ì+˯>�o�-��w�6��T�
��+w����:�P(��y��8�Ԭx���:�~���t��o��!�ia߼�ۇ^�+Ny������:s3�:�I�~��N�VVJ��_o?y����@�����T}��@�G���xY ��
���y��:��VJ��FW
���)i"�[������j9 d-G�����8P�3t���+WP��a��	�~�ԅ&T̨
$|(�|/��,���P<�{���!iHV�+g?}��d �ؿ��&������p#z�k�Y�J��P���l�Aa��o�>4���Ĺ�\�Xv0���?l8�i(��|εN�W�I��>�2�a���P*T�>��@�V�H/���W��Hx�����Q����1_W�
��E����5u�io )�'����t@����2W���n�
IXw7���=��א��°�*J������Ad�+%_ן�ܜ��5���ɑ�*bb���#�y�}@L���w�����~���!m����9Ґ��H-�9��@�q�T���{�u���~�;�'��pڲ7�p��c(��wGȥ��ޣ�gfyu�{��ū�rk����U���JX�w=�ŜO;֟�$�O�=g�%B��y��gP蒰����_ƍ%��-�6�]����ID*J!X{����β}緜9y*D����é��Ԃ�����p� Ґ�X~�߽�:��]}毕��xo�G��Y��.�`X�y�q\p�ƺ�`q>̇U=<ϵ���ߟ���yq:���w�ps�9ݜO�
�++%}����2m
��D������y���wO0޵��8}����vq'���������ۓ�m������Zt\��i�}7����"��cqo|��`
ov��������s�܁���R��'�}��ì�%ed�~���y��:�u���x$�,϶�s�K����5�u�F����m%*K�?y����:�YP*T]����㻯|������*A`Q�����)B��=��é�u���N�]�ִ��/�{�w�C���UI��Ϯ~ i�2VVJ�}���IP�+����a��aRQ<�}�gRk���y��|�~���C�J2�Q��u�ہ��=��f�7Y�����+���tz��H	 ��P�x)k�[�Q�����I��i�������i �
�'�����R;*��l�IXyw�{����$���s�b�.n��b����Q!�{7a�O��̇UU���<{�^�������1��"Y�%l�ח)ŲqlSj7e�Pݘ�)�E��=��y�$A�q�����'6;W�]�^|��۾c�n:����m�W�����bh�f5v�kk��&S��k����PA�w	�O]Ee�:6��i�P��۸s�ٻv����&������g���}�]soW�58�c�sH6���<�٭ۈ;�\�=��g3/��ōl�"�շ+� ���9�����q[���cke��B���@u��:9�E��B��Ι��<𻭱ImFH��m�d�/wS�܉TsC�}��}��%��-�����yu��ID*J�a�����N��J�g��p�R�;Ϗsm��~���=��|
:�r����)����W��`VΟ���ᙍn�ә���蓵�m##�#��vg8:ϥ�̥��2m
$�Q%aO���y��¤�O;�~�ԝ+%���;�?{u��~g�u�|� ^��1*��2H�H�V����tz��jB���{��/	<@�c�\�=B�]���o^L�o�Hd ��'���W��a��+�3��+�Ꮔ�1
�W��w5b����Ȓk��T�u�d�v�z��N�Ԍ���g!zE��������8 ��jH��N7��2��v6��օ���j�����$��=���?���/��T���U��v����d�8�Ү�Hsv���= ��;����뿟~��Z�7bh�s��wW����$���#Jt$c���ϛ�$��o�Y�;�"HQ!L��"���7�o�lw�i
�&�\L�	U⹶��焧�/i��������rza}�z�L�[=�y.1���Dӻ�`ݱ��Orh�:��x �߬�I#m��`�I_mP'���Y�U��gn�D4I#�SݕI���ݚ$����"��UY�Ė�:�	#o���UF*�L�
$HO�"�oh�;j���hO�{�C��i탒l�	&b"&��w�D�s^����k�S�L��̻�C���y�볯LtmCȹ6�(K�����X{�7=Y{������,o�u�&b7m�dF�Y�2T����P�]e��$F�mQ�y��UK���'���t�r��Ēv����Zq2"RLL@Wf�Y1I�R���]]i>�H;}�@#�ޱ~:�{_gBݬ̗~$�=�"HS%L�қ�D���gěP.1��56�Vm�ۦ����ɉX��N���{��I={[�V�ئށj��gv���u�p-ޣ]0yF���<Z�x7���d
������Kg��K�xdG�Tv�G%�Z4�0��ϥ3ݍ��J��}���kx�3�ܛ��c�ݒV�Ӌ�oq;��&&��8�[�1GaKS	�ã-Ĉ�FP�^0�&e<B�����ifni���y�:��tS�-�6!�;���b�5Bۅ�2��p�Pa���d[�Rܸ�8T�8&.}�M��V�
���.�<sKμ{X�plS=��2�7���2e��������@{���iӃ�Y���	!.��+C6�[�~�w�eMMo�����~��=�h.f�l�L]�Q��bhb~ȣ��h�;Q����]����C�k���A�j��]s�-�t��x���"^4�g�}��������O�UފW@��%(u-��*i��د:��G�K��پ����m���ah͕���&���^����7�w�	;�7\��e����O�y�Z��N]]>@�u��&�{#jF{��-ǀ�� n��:�n�չ&�э��F��N����v"e�㻕Mn�l�j�v/p�}u"��k%	Ɯ��c{�q�$g�5t���f�y�ǝ3�(��\�ۉ�:wuUs��2I�}a�k={�<�<�o��h\&�v�=���i6u�<�W��y��GHo)�U<�}�}Ѥ\������u`������q�s���&����}��{���ʙ���{��N��a� m7L�[*�ZڢZ(ڢ�m���-�Җ��h��K+[IU�m*�F4�R�TYh�#P�2ڂV�m�����b�[h�J�P�!VZQA+JұJ��[iQ1QQb��R�+V+-�4�J�J��+Tm�-m�R�5�(��V�-Y��E�-��R��4�6UX"*�-Kl��C%V�mR�������6����¥J���[Q����R�m�Z1��"ұ�QQ���-mE�Z֖U�T�����e-��P��*�[J�kj������Ҳʵ*"�e�\�B�R,0TR(�
�b���յm�)mZ6�-(��IER�-�m*1e�F�����
R�j�,���#-�Q�X��EJV�m���--Q�UF1EEJ��(���Q�Z����*�#ьb
���PZU,X��E��h�Kil+-��UE�l����T�eF�lD�F�Q�"ŊV�B����TEQ�&""�`ʈ�b��k�"�2�aZ�X� ���UQVV���ŵ��*�lAL�i�$s�;߅T���ؠ@$s{�ߍ��ʁ�FT�1~�զ�aV���L��_O� ����<α2����uI �/g��F��� �H,:�p��F�`�d����P�Qʊ@��s^'����� ����\��g�a�_�Ҫӹ�0p��:�,�ѕG��=������j��:3mnY����]������3��
<�%��gٯ9��$�w�vP��%�o5�D����P$�=wd�:2fJ�1
3�ZO��R�ZU�f5W��Pe�����?O?�x ���t�r��ڹlɘ �FT�w�v�XA':�j����zTN��1�uK$����:�Ŝ���2$�"fJh*7�ё���3��:�ę�Yb���{vI��p�]�Y���oQ�S�:����6�>�'�6yF��_��&�Epj^���<���y��R�`\RJś�*�^��j0�x+b*)���� <�9����X���#Љ�0b.�����$�՛UuM��wϭ箬z�m��9]S�m-b�_�D{����ķ�դ��$��<�c�a׎�O72�n�7�w�ף�{���~wՎx�	S"{Ǻs+�<�����)Sr��u�݂���ŉrrI�*&M�<sr�E��S�u�T�e;�kڰ	$���*�:ɋW�⮱�O�@YR��R&"bAB�z��HNWT����+��君��2u��  �� ��j�0|D���v������1��U��� �u�dKYN(�Hx�ڛ�A�|��[�'�*��',�\��"d�Jh���I�n���^��=�Sh��w�|	,�:�v>t�QK��Y�l=�'��j��M��~S���;��{=���1��=�c�������g�Z�y��D5���gdmZYw*#o|  ��H������.�Su�l�ʝ�m�;]=�8��<�۠�Y��,��ǫ�� ��ȳ�n�N�����cu��6|��]�l�����s���۲���l�oq8.8{C����l����2��Y��y�� ����u�m�v�z�g�Y l7un�)��m-+ß^���.�l�����e6�ӽ�^P:�n�Z�m��s�ы'E<H����-����e�kkut��ۑ���+�ʒ ̃,=�1#��0�/�}��d��V�	;�u��:ޛ���bUs�$��[TMJ��2���%2&�9��d��7f�\GS�Y5UV	��/:�@+vʬ�w��oq�	rNB����
��vC����o_;�O���ں{t�*�s�s�A#r��@������D�(L�"`�Ȅ)�^��":�J���o]P�	���ud>��s/Q8n��Y����ڣ7Զ`������l7�l`y�y���*�r��[Ӡ{��Y>%��݂v�d�f�?�����-�AY�NCU�#��c�-<�	r�y}��`�e�k�����wﾺ���8.WK�D�m��I}}�1��޻#=]�Hͻ�lgs*G�"aDU���X�tG8ۉA�;x���Z��uZ���Q��y0~�]��>�nv�_zj�8%��_�)���|���}�V֢Fz�9!im)��bV����������H�|��%�}�d���g��a�'��T�$Ɂ2��L���Y��6�đ�Cm�Q�Q;,�{����_v�����b՛��u �`�OG�m�~4�B�3%�Iz�l_�#2�V\?L.�jS�_��_w|���yH�F��Ew^�߉'����;B��m֓y�N���N��v$fgMv�ַ���'
���lg�<v��mݮ�KL�����=s��i" D�a�u�F�O�	�!*3�VfҦI���A9��^&�h�$�#Q���݀H';;n�I�;�B�IR$I�f���^=�hVz<�{�d��пFfu
����Q�k�=3�d���V�*�N9�����,PO9��6��{.a�ꪠ�
�ͩ�m�
� �	�P�}8e`u�{ .F�|���j��i����s|�h�L\i^8ˉ�*��#v�����M�w���|>#/>�D�\eD�&BQ&h�M�\j66e��̠I��ڲ$���G=�}�c�F�|�k`m�� �Gp���/r������.�uS�|���Yo
�{����6:VT�"	:�m�y7O���զͮ��V��8�nXG{]l�21�;҄IR&L�C��e�>$7���A<��َ9=�
�{�!�ʼ���t�mI�u�)�%(�R"�S�vA΋�ѷ���������:�"L%�b�o��A�"�J�"L#4hƺ��A|ۻ��U���6���G�j�	$7��#^�`P�l��
d�������3��׉<]UI���ݒ#^���G�y�;uN�2z��7ե���s�Z��os�)�{;�z ��q�]�t�"8��Zy���h�L��T+!su"d`�+w��<=�$��2�����&TL�d%f�U�X=߶�����M¦ȣ�:�	&޷v	�:��쭊��'�=���8қu�Ym��&����ml��Q��ܻ��Lh1��b8�?�Ͽq�����5��;{^�O���vA$�{�a�V�{���<���>��s#�s�a�ʂ�#kb�>�ƽ9��+�6v�u݃b3�2���n=�v��$k)K�+��S�%�c�#a)f�FDT9��V���@|=��uDU�{z�tgw]�@|3�2� ���!O��$�7W��5V75�;�y����#�������) �-�m������f�A�Ǚ�X��TA��eÈ�REuGU@ �]fz_��o�z���*����P3�v����yz9��(��ѣ�ۥ�F(s��3�»u��|�yL�^���KӴ�~���w���4Ӌ��<���ڋ���5F��:������=��2�#����a��9Kq�3�/�ю�nЭ��cp{]^�ac�vz�^εD��	���ݹ�qԜy.�]��'�m��ٲ�nni��*��H�a�ku�1�r��]�n�����y��zN����[>y�콦i�>�mu��/dQ�y�����ík��gע�Yc��"�Q�b�����e��:n�;w=r	�+�܄sҝ���z�j��xS�{7:�;��!�9�p�V3٬u�s��H҇N7g1cf��'Wg�{R�����P�k��������^]�cb�7v3ä Yו4~�Vo�vg�5}w` ݌���֮�!̒nu 'ý[�<���p���s�oJ�Ϭl-ݜ��6|[�ʯA����� ��"���I	��Vj�R�-��m��@ c�ʯ����'�0vm_��� vle��$c�ʯN:�6a��E
TTQ���+���h;�7Ԕ�-2���@gn�ٰ��]:�@&n6�I����?K%L��G���+�>��gg�C���$�*n���yYUၝ��V�;��65�����r<��P+��`�^�]}5�3z!Pͻ�T��[�A����Ͽ�T�a���>�썪���g���n�]��:�w�����ʨ�G<���"�p����7t�Ǘ�;����?�\��N�l�J"��]�zo�y���B����jg�r�4l������/��~ߖ�FQ uͿ�y=��_-����p5��P�]��{���
�t]}	�I��̈́ �go�@�2�%���)������Q}�f ĩ�D(�&�&i���u��j�������~޺������ �����B�L�9A(�PS�n�]J�G�׺^�)7!�H7.�)W��@+�޻��@#3cj5�+��Mz	o@��"]nUx{b:Ba��E
TTQ�{�gH ��C��y�MŦK<�Ӡ 3�z��3cj��=�B�ߘ�lg��X������ڤ�끅n��\���*H`��M6�S����~�J������J�}��V��͍�A����(���׆ ���Tv�!���%D]������DҾ;�/Qo*X }���m� ��ڥ=�9��x�)����G��ոViғg�YM�͍�@ �ۑx��=��P��zjjd[�+w��)�����B#,^{��yuﾚ��%�]1��u��(e�8�+6�٫��uH��� <</��T�H�~�w` ͍����]�f!���&[�����ߔ>7#�Mm���{�j����) l���:){�ۭ.w�>�����9���29A(�PS}��( ^W��x՝�=� ����Fnm������ڥ��W���_/��w����:dD��Wk[b��O$N���܅�ݶ������zۮ�w��ϫ��3�*n9�@v���6,+���Z�n%g����;cj��N��*P�"}�_��<�Ic���w�@n����@벩xbÜyݕ�r;����pD6�e�&*�]Q�::̥^N&�'z⮪��o����P1 c�ʯUp��10&D(S7i�n�K}3Ë�}To�@���=P evT�6,�޻����#��߇:'?`]A)�{~|%��:��ۛ4��1�����8��\���j��5��IO�Wu�z�T^Yf�]���ؘ'��� I?���
���A2�!D�4O�k�	/%���'�ft,�U��?;���I c�ʖ��o>�Ļcr�*f�j.x��Pȕ���Ǆ�^��n���׭�x��5�ڳ�F����ȍRܠ�L�-�n���؃vUy��޻n���.-n�=���Uxb �]�.�ODl���dj�����뿬>����V�t��������g��@}���w�a�Few�:�\�{f"��	1"'�Q4g���D�ϯ1$>�]�7Jss��^�͎ ~�^b���#w\�(�0�V�tN�/�����K�eW� f��U��;h�����u>��� �~��U���ba9��&j���˵cb��A���U8f��Cܷr���	ko��ė��n�Uz���WU/��ۋl�,�Nl9tҋ�Fu�h�p��ѭ��9��&6sT�5��3�p^�7��=�=;��)� ���wj�`�)�&�yr^;�ގ�J9M��[�_ZK}=��؞|�}j�1`�w�6���ڼ�4Z��q4�FmbQm���FZ��O�Ƿ������wH���}�*�{w=極��lW�����e4�Q�O��)�YÆ5�X��"C��y������]3�ޛ2�	,��u�Lڇj�G4���v�k5����p��F��*�Ȫ�')��hV��l*-=|Ĕ�A�S��{u;ן���dE�!ܙdEX����W}N���H��j]��w��qgv<A��^!�Xvn�P��=195�Tb����hɧ;�<=�S{��)k��o<O@���lPynY*�)������ݜN��A�#v�ⶃ��snX�՜_n3bӷ�!��Y\���2�w�y�a����R���=l�8��bY*���Au�43��F��i$t�C�Ӳn^�$���7'-��n�e�͉�����;�$�А��\�1i
����P�t鸃Q3�L�Ҥ*jSn������Ks��{�E!��Vr�;H%f6�RZ,kr�S�'A�Ue.����{F�=Ù��];Eٸ���<}�UMsz^����uA�<�з�ϐN�:����E`~�B:U�s�#�#�����{��|dh�XO�V왺P+�����K�#�W���{�)GO�qf��`�۠ � eW���D;�obƭ�,NA.v'i]�FJ���|A>R��m�cj��F*�9j�ȉZ�QTD[iH�[R�T�ĵ�Ʋ����A��V��m�eƈŖ�V����Q�cJ5m\�UbnZ*̴E�*QTJ�PU
մ�R�Bƭ��-R�UVR�(1UcZԩK-�jT�E�1b5��V�����"�h(��",`�5(���q(���ъ"$X5-h�[l����B�Bʖ���F,e�Xԋ"Դ-h�R�-mcj�[iJ)U�2�ɔ��-FU���ʴmJ�--��j-���TDU��Q�(��6��J��E�YJQmR�� �A�,�����������X�)Z��-��)�G-ZִU-*�H�)h[Z�`�j�ZRֶ��QKB�TQP����-kj�"�J�D`�k,X�c
�6
�aTV��*�(Z,�Ze�F�R�J��KUhU3��Yh�¥b(�Kh-mj �J"YaT�)E�Q�l��mQEZR��m[T��))Pc���*R�X;�:���k�eQ,��v����M��N~7v�h�m�F��m�gy��-*��{�ݰ�,ga���J@[O`:�n�|k��:���;[��Z��)����u��ڻwlz���V���t�]�mc]�\L[Z�m��+���K�V��WT�j\y�Z�v��!ӌm�/&��n8E;:ՍC<�_A�C��;V�\���`ն�>�E��<!�ȜA=`7��vJ�o磜'g�iT���۪.[9C/[��4��')؝��x޶�=��K\�9��ٍsf��l�t�g��q��{�.ܘ��n��1��u��l9���ρ��q����/I��M�vc�4���۬lSѹ����9��n�0u��6c]�������u���1tnׄ͞v%�l��̌��ۖ6���3��v���3�1p�ݴ5f�ٍ��f~K���=�ˍg��4_>w��|��d٧��cB�Z�m���m���]��G�ϝ�ɺsڋkq��l�t�]�\޺�fZ�!�R�k������|�>��ι��̜��c���/��v��z��.��qn;5�[���ڹ�:��ƕ��=/�lq�z�&\瞌:u��옋.���s��dS�3��gMq׶zq��0��TiN7nɄ�Xa���tsq�����v��[:-�MK�2�u�t8�X���z�5�����i�z���l��W��=l�k��ћ�$y�͍`�n�6��{9���z:e����n@�;F�g�}��s�y�tqV��n����ڝ�PKְ��.M:ܝK;�vN̏ r�r9;;�ʹ��F덛g�u��۵��95�ɶ�ۙ즶Y��4p܅�w�m����5�*���c���j�ڇK��7
Vx��\���V-<^�����.r�vvk�n.�.�R;qm��.^=8�h�^�_�W[�v{d.y��Lcl�m��_<d�d�v˶v��9E������v�u���n->ƪ�ۑ2�N��gCu��l�c�7\�5�ԋtfXqhL�\V��{���|��40xx�����˰"������M۹L��N[�[�ɹ!�v�7GK�����r=;,-��ۃ����r�Ǿ_ ���ó�֌ۑu�Q�o.�$B'n��ub؎5��.���:��ʦ�mn�p�����ѕ;c�۫g�)��.�{g���َ����8�#n�Ƒc�Y=��ڻ=�j�ջ�S�9�l�#M�W.�9^�P�l9'�KN'���x}l쩬l�=�\Lk�H��f#���I����f ��I�d�M���.�H�m�Z�ϲ�v���w��P�v��o��>fv��v��2�KbDʂ��[U��!�ɪ}G��]�i �W��v��KN7wH��dr۫��×Y��WDt���eT��WǺ����w���u����̓��� �gv��m��{����3V�	h_�5�'��$�>�����뺵`��M  B�ˬ[���~@.���wk�!��#�	����Ժ�]y~�{m��)��yT�ͪ� G;ݩn���:�O���!�9�h s��8�)��.zqv��we�c�I3��ѷZ�θ��l�d�~�]�뉘N%�5���5�o�����+�����fo^eݠ>ͪ^�(�rD�2:�]u�T����+L�kx���SD֨q!Q�75
u�7�B���cg��;{Fq�e��ی��U2K�2�K���5������ݳ]u��Āӳjh >��T1��*�kѴ�N��|
$A\��8��Tt�u[T�k/���?(��2��n�ƾͪK����U��荕1*L�FD���*y݃��P���4�A��ޗI {}��@$���'�q�5|��y�t��;1"`I��� EՄ�����I���>�MTu=�qW���Օ4� W}�_PĀJ��o"�W��\y_�"-"a2Ht�i5��I��6���u�3Mvʳ-�`}m��q���3���"	��S���� [w�.�A%��ݙ�#��Oj��2����;��6ą�}U�k!��D��p�L��]����b�\���F+�8Z네��m�{�����]�������&0�o)�-d��2D̎�^�*����괬/X�م�j�w�Y�'I���0G���ی/7��/��	��ݒC�t�{$�幨vv�h�rkb��5EK��M�O��������$�nc�_P������ ���Cs*
u��V�d�f�?;��:��g�k� ������fԬ����N[��{��#���)"�@���{��р!7�u$�����Bwz��%y�ݙ�H�ܛ�0g�����9�p""eA�q#ڬ�[�����]��:n�n��\0��Ͱr�gc��
`��p�g�uu*��v�uZV �wF�E �#z��mS�H^�ʥC��w`/(��}�*#wV�_���$���s]ہ�Ͻ�͒@�w]�	��n�7I��X�'�����J	�LS&}��̻V �i�� x{�z��{z�;��� �������ݪ���WH},�����{��c��{�Cv�K�Me��$�7j( ��)>���sY�nyC;Z�2x�^OAne3w��!٬x`«�m����$M��j�w���2�O3�s<���j}[�\t��3U�N�xB~ s��9�8�G5F��J9��x�?Q�U ��*�T�i*���;�N,�	Gz������T�
ﲩQ��3LvFS���y�@8NA��0���[ٶ٫o6D(���m<v+�s�������Q�K�*T�rG��n��@q���$s;n�'F�N��.'C���� ������&��$R�XV�|��~�>�q���J�wۙY`��w�����`Z$�d�aa�[x@P��!G�8R�""b���z$יJ�ʹ=}������v�F�Y}��#\��X	K7"5.x}�K%Ν��G��M�Fw�A �̯7@,�޻ɚ�0�ɂ��I)�N�J^���9D�A!$CxN{�;�d�{�9�K:����}F��� ]vU*�3�����{�]oNϖ�ݼ<�1��[9��d�*r?7�,p({W�4����>���Q�Hȣ6RK*��.8��CjN�n���{��~�ŏ��c�k�
n�{&r���I�`$�X�L�lōۃkoNvc�������#�0셞#���6�}1�(.�;�;�"�^w`v�]���>�r��M�>IItPC�筱ͅ�9�%�g�:ҷ�\.��qz�wKm�ӻO!���*��<H��%cE�7�Zx�=�t6��8�#����g;��q� �/6��y�M��C������m�`�6Mnxu�<��l��;��Y5�t]�u����������<����[���H Y[��P�@fv��jOX�<�7�r�����;[d�^��:��Pбbz�z{�2���8�P�Ϸ��}��H؀Ok��� 37z�� ��6EWDt,���M����!LL&j���uD�M��I5�뭻��x/�^���+��y���6��	yF^(�i��"DL��[WO�M�7���6�e$���R���w���3�ھ�Eet^Ve�@|.��@�V�Ġ"T�H�f��s$H$�n��P��M4\'ݷ^�Aۻ�V��n������=r�QQ���`�:�	��%�M�9��s����9&�<Wr���n �.1>:~������ʔI�~��-ʺ��� ��V��[����'��C�8D�]Q,��y��v���G|��SS�h۪�@�3U��kk�`���3�yӬ���,��ɻ��OV�lA_g^]Ֆ���oYrm��6�A��/w� aY����Ӄ������B�2�(eA���q_�����@�~��w`�7}����^�^OC0+ެ橻QԀ�B�k��{�iX 8��%#g����V�/�F߰ �o]�	 ��v�H+3�$���Z4���WUVp�L}�W�� �n�R@ �����+ٖ7���IC�wxTkA�D(���|W�JA �=���%�d;���E wm������T����}��y5�����V' 1�5�tbI�KV�4���85ƍU�G=�N37c�:�<�ڐ�?]��L�R8��H�u�ڰ 7M�C��vL�*�I�4�v-�̻� q�U!0�Tp��R�H��U�.�y/x@�weg��u���V��`� �cv����U�E$z�i�p��fWu��eQ�?�J�0��GQ�P۠Y�3�M����}&�kn��sjTЛ�;`����Z�q-��7��d;�w�q2L�I�56�95��c���y�!}i���蛼�u}/��}�� t�}�I#�&��(�|,�����z#	��� s�E������`���$Ki��I$GԓHWݷw.f�V�y��.��O��I`:��>;�$ �Z����&�t�I8���@9���v"	+ם�0��Hw�wrn!X.D($�A,�!�2t��^��t�&�v� 2p\����Gg�;yDC�!J�"fk�+mT����}������x=3��fI�u�H�o3��@ʸ{��r�#��+�[&B�n}
��S���+�E$�Aorc�|���ۻ@ۋ��k��ᶴJ�����D#� ��|9�r$����).��U�;�[��eGx ���^g�{�wh;#�B���4����F7��p(��( 7��l���m���3jVu9���^M����A���KS&o6(��K����M�V�e��uB!�uX��Q��LȑA��ב�N^S�����'Z��j�����#����"\F���R�)Ϣ����X ���Iތm{�vG�H�9���ݷv���W�:�3�kWtx��0PlA8��Y�a��X����<�\f��;�qZ\q���v.�Ͽ߿J�fS"fNs܁U�ρ��ݫ�������W�(eC���έ��T)Wc�NP��A�$�%(���*I�=ʺqlFB�����n��Z@ >3:6��<�WH�EvK~�Cؔ0�$>�wf]���767Ԡ ;��)��u}R�~��ۻ 3�݈J ۃ��$�JTLɻ�A��<�9�w�	 YYWa��ӴRھ���d����}��`H�����d�S

to�6��@����z�j;��[s��ww� �U W��~�`�t�D����&B�eEV:�4͜����]:��1ye̘tj���3T��TT��צ񐮙èf���H���}�u3ty���H�T� K�ˢ�$����s568�(�"b �:N��ծ8����Ϟ�]֙�q۪|/o��9"1�t;[klx�Ű[���*ț'Vۆ|pb���ۜ�<6ѵ����h���*��O1Ơ�p���m��;rZ�܇&�Mcb��%�v�K��/�*]���������7ty��aV3o���m�N�'m̆��&tY;Yޣ���lH����e{s1Y|M��t��d����c����cG��;�y��!��E[ջs�������S-�2S��5Y��%`����@h��U.�u��L���ԉ^N{|��'0[!ԒKԴ��５�E{_z�4a�./6�� �_N�_ �HW��xb�/���%s��H����&�R�"fj��� ���ㄜ&Ύ��la�KT�͹��^^���b
�=��/.�A3 �f�]�k�?l�?w+��3��=���� @'���  ������T�,�z}��ǧmoI�Ap( V�Z��A�Ъ%��;�b<��eҸ�����(���}��;�����Ta��?��~�?��<��[��F�<t4��f&�;��Z�{s�v�=R��2����W�u�=0���}�� �e���gv��Q��Ho�8��_v�@xI9g��2t\28"JsQ_[�wcj�=\r��>��"�+D
��D�٩ˊU`,�&mV�4�U�g�Y玨���d�$�_t����sih<��x	��٢~	$�/M$J�<�sȾ����u��PK�y}	��RI,fb!���^��x@�nի�A�
���o� »�{�lU��wi����($���2�������<���[��߁E_��$�e�mݠ=�����h�4�[Η#����T)/,��# �pa��]�v�>��ݟP5M�[ϛ���O�@f�m݃a��5A�;���s\[O���!9�\�%Bj}sǎ\u㲝<%q��F�gN.�ܶ�}ud�~����{n%��DI/y��/x /3��X�{y˃�m-]�[NG�wI9m�����q�$H�0!Y�.��v�>3议�' )N���6����ۻ@ 6�t�}�[�X�P�}��K�Q�D��!��>���������$ 7_x;W�j:��4�<�n
���c�Ab�]�a�d�b�l�@p1���;�<]���恉����t�ɝ�:IX���(�<�����;�=`1�^��=����8_Q��H{���ވh�)L�{w:�}x�2����A�X)�~>�Xz���MVny�c��t�b�vv R}�]�"o��əב�eK���'wlM��ca
�s�#�dw/��W iq�k�N�B*3m�H��۩$LLS��1�ƋuF�)CG]*6.����wFy����CJ��D2��ez�s��{*�5����\+x��{����Ν.ճ$���smV�V��y.��:�E�I�J��9���w%~%1y���jUx�ֳg�5SP���C��O�H�M�:E� .�\{R�2�����j����@��S��O���z#,�לi��FaY�����t<��1s���0�ΎX"�Dfw,|�7�&d]��Q�P_�Tl�ezc9 ����uyJ!~{��0DN�Z�\�ECتA�լ��diy�s�&�����]bs~ӻ�/�#�W��x��%EO]'�!YPtR��6�YY�rؿ?L�D�E>[頭�{�HӕW7_�frYT�3�nѱcb[ְI���w��E��S�XW�N0���FؗPbJ�4���.�9��f]ɲ�$,�IyQ����;ٶ���g%��n�s�s9F^é����U�I�R��MFxuOޝs�|wQ��권� �;�����n)�̌��0���)��5��9���Q�[iR� �
RQTb�TR�wJ*�UP(���Zն��m��R�-�*�e���EDAV1FE�,UDU�+[Z6��ڒ��Km�J2�h���m�����5,D*TE̹��9k�ZʊU��+b����UDV6�[U�QV�Ŭ(���EQ�m+QR�*֢[[j������"
DR��U�jY-%EG2�6����R�U(�+�TLKEV��iTTX�(���ҙlC-`�Z��B�6��h���)KlTUإA��(�R��i`��X���R����kKTb�R�c�2(�ZUB�*�F
*��-TAQ����Z����)KQV��,+�	����+b��E�*"-�YP�V��jV
�R�G�,I�Tb�[l�q*�Y2ТT�[��0��/�������m�y�ޒp�����3�$����T
��)ޏ�zmq��*�7{uj� �/6|���W}�~�j�E�ߐ.Ǐ3T#�� ��"J���T�� @��{�>�M�Krt�Nw]�"E�˙ �$�����6͊�G��}��������^x���ы���me���i4�uv�Ŏc&یu�����~�����_�~ۺ� A��>����;���]~.^Eɯd�����>�7�8"�3D�4HuS8��.��NF�{;�V���S� 5w�����vz<_�Ց����9�����*%�Hݫ���_y{��2'����{�y| ft�5w���JT��1	H��4�����+4v��(��� mm�Ͼ ����u�kF(���G��L#j"��RH�>n�9�A�%��B5���y÷��H~���ZgA�Nr��sڷ=26�����}��ܛ$t�F&ffAQ*`@��H^�UD�$���1nѴ�r��o�][ާ@؅�����	fom݃D\������翫=�xzR���Ϥ�lv��<Q�q:�n��m��n.#�v�;��������4�>��w&� ���{�x� �K3{n�����[lF�~YX��"JomU%�vYČ�e�	�&�#k��ՂA�����7"��ʺ�&�%�jhy$��m�0����w������&v�r}�a�s0��]Rޯ/x�v�; ڬx��W�w�d_>[�>����Uh	&�P��*%��}S�L�\uT\�9 �o�e��۝�v�@��U��8��� ����x �q�3%D�?mv֫ 3:}@�.=9�yV��9`?wz}� n�mݠ>���p���z���9�҆ȍ���̫�|�bb���Z&�Uû�.��=���&Vs����78��12UC[
�r���7P��~����N�Z��4���8
[n�!ݍ]��v5�맷�;���6(��/D�#ݣq�Vݺ�[�m�mq���<���u��	���Q����k�u�k���7!��s��9�:���:�a�t��\X�V���ܴ��n]�ٱ#��\�ݨ��&I��=���n�[��Н�P�cv�]��Q�׷lc0l��n��Ӆ�Խ7,[W��/e��GY�g�\C�J�֒�Պ!��:9��=�M�}�unl;|����ՙ�L�&)��
�����W`,̞��_�s��X�1��T���Kٹ�3Rl��D	������\uڀ蚧���˯��� lKz�n� ̎��A�7�p}v�TV�<��$r�@.}GW�.���ndo�  =osƿ1�����}�}�v��U�o��08�.�z�x��T�#3=���괬 -̞��������꜇V� �Wf���!��	�"$���y�]l$�	�Us9]�O�����s#hn��{�x�U�J�X��N���J ���D��>]���zv:�\�n��7Kl�{6����ێ�?����V�����H��mڰ@$�w�H|��ښ	8y&�WWN�30$�;�z��w�UL�����
�}��nϻTL^¦�wbVWnX�[
��Q��ૺ.�Qb�@5�b�q�p�c���0锶
[������5.az-2+�Y7��X�b]��Q_���7A1���5�o��,Q������$LE9�{ؤl@�wj��z��gDP��e�� n�R0+�ڪ^q!�J�&\��WUc�}�͇�������ٕ����R@�I����D�W��od�ڽ��o���.!�/ԁGz�U6��n�����yy�=/���**��$��\���۵V�M�{�^{𡵟��</]=���\���
�tv�k8�Ѻ�=�n��<�68d���C�	�#�p�5����m��󪴐I�n�Sv\'��d*�wU# B�ݪ��	u1	�49޽���lc���Zdd�އ� �n�l����I�s�\�����]pp��:��P�d!��5-���U@;wv���dU�Mth#�7UWޥO޲��1O(GGw�˵n�wf)��w���f����o7�v�D�BN	p�kӼ�}�.�m`l]����ws���r�q&�&��Iy���S|�a8'L�f�(3�Q1aT�ַ��Tej~Ixgo�H���� f��������.؁���y�{plI
T�e�Q�Ϥb����!q�VU�@�.ۺ�^I=��3���V�ؕ�P��X�9�	��0�"�&�	Bs�yw^�}����gy��9�l�<@�|t�������7E���?�
7��7H/s��X؀�23�(=tl����RY��tI6;u��	/J�*T�`DY-����FDVR����^z�@ ;s���@�Ct6���ݦ���~�iA��u#��	+Be���{$��u#~H���-��ɇ�檾 �s����FfGU(�{&A� �MM [}����fTZ��$ o�2�� >vd��[���&n�r��FLr�p�dÓP%�Y��f�ʘ��q^����*l��O�Ĕ�q���7�ܰ�{x�L�i/"-`����$gsr�A�����U����}������;�P��$LEQ��� ,������Y��Ӳ�Bso*� ����s��砩��^����}��l.t�hq#vk�^���<��X�Nz�{R����>��V����~�.�� ˍ�}`s��A�vΕ���ڦ� ����P��ɵ�d�@��v��Ywh�r8:�_8�݁�1�U�� ˸� [��_Pۏ���V����󌼬I�!�����(��S���A!��I�%z;z�2��ɺ��WT�`[��J�	u�&BHP����}Uo�| v�/�bIx�󺴗��|��x��
�RIy���	�rt�d@�*j[]]�T >
���$D^�s��b�]�Iz*�m_�I	{v�� �7���'�]�'��}�Λ�&+RN#C�/��u��T͇�NL��4��]"Ω�Z�v�:Ԭ�ЇB�.����ޮ�\ԇA��v��l��ݷ9.Ӳh��;'��r��Ga�ݾ[�����9�lY�y�.�¯=yz�y6ܦ�+��v��vn�S���������u�N���I	�c�A�L]�+���Y�.�)ú��S�x��sh��Y:s͍x"�=�68����X��6�0e���=�;BֻE�3����]W�³\{&�l�=�n���9벐���Me��K2�y.Q�e٠!41�CF��g^ͧmɆ�L��[u:zbB�I2�=Ǻ8��yD�b&"�U��� ,��z�Y��m�]}���]\s;+��{�P1�wj�����ѫ$�<>�YP���^��lg�@�;���$ 
�{n��n�f��][|��d�Tz����CB�%�.aU���� {�W���FDO��e窯oj�@ >�mU�����I>dp�9$q08�tkʺ���t�bT�ؐ6�޺��@�W��w��>(��櫞jE�/p���������L�$(	�>)[�w����;���+��菫�wٵ�@$���w`|L�uإK(�|��R���"*&3s[��Y����]�x�j�����l]����ݹD���
T��@��iU6�v���`����4�5�f��x�;��C ��s��^˨e#�'��.�����;����d���k�N�H�q����ro�s��v)?&����hw�e>k}�����Gb�.{uS���Ϭ��Q�a7B�67��G!���D�Y��`�Wޖ�:����ވݘ�]���{bH!ħ L��F��ݫ��u{�t���<��8��7@{sv�� �w}T�
a�W�S$�%�*�f�T�^^�Z��A[뺻>�.���6
�:��_�f�����	sO�Y
Ba���<���U�� �f�UT���W}��|�^�X ����x`W��TF,n*����vK��r�&$SE�i5��p�s��[ؘkl/�[����w��	-�w4��C�'��! 
$�� 9�O|��2�@#�{�j���a'	Iޯ�	�,T�`@�*j[^��J�s���;�O�׷n�ձI8I�ϚxQ)��`Z$͸�����n*v��c/ьB���� ��<��U��ݪ��Ib�mD��*�,�q1j{j������E�γ�[%0� Z��������+.�a�h��Zi�/fc%ۚ�W�7�����=_x`�Ϊ�2�GD�D�%MR6�.�W���[�R�@$�Լ ���� ={�vz���z���5��R�)��^|1L�.e]������$��;�b�D�-�{��T���SH��uW�1��;n����Ѵ|��w���<�.�tZ��U��J�U���:ڞ|��j���?��߿G��
�B"�|[����@��ΥT�����:'&"}��/a��j�� ���<E�
պ��%j,2��щ�����;�9����ٝ^�ם�l�Y�D�5b���=I \��bR	R���V�R� gn�6�s��Փ㷺\�����^gU*���l�L�����u~Z5ke����v]v��6I!m��^Ix$�Ow�	$�ו4�d.�S�x�䬎��F�r���{��4;���\�o��f�[�>�D���N$�K6In�����:Sbs.*(n��\H�˺�- ���$��c�ĩ�6���X��������jw@>���t��u݀_^z��d��Νȩ]�pv�9�N�Y�F�ݎo���ݯlNˣ�љ��c'��NK��߽����\�&TJ�sw_U6�3��l�f�ߒ��
gn�Do�7n#�on�n��s��9�!LD0���e� e�k]3�>��$��}~�~$���וIx`my'�O��uϫR��_�0LLJ�LIN�=כv�> 1���� =ĵ=k/#�U���3������^�[�N$2�MM/�V�oD�:���&nH/���+����� �Ϊ۷��5�x�W��wh+�L<G�O�&<����I �	z��d�A`���UX]l��` ���x`Y��_QI^�[2-�2OEtvD�z��"gk7&�h5�>�;��	;��� ���S;�_d��=�ӵ9�KOa���9���5���`E���n�S��G�	�i�t���ւ�}�;�O�����tcgҳ>�$+.�;�f猸��^(h�����fL'I�nT��b�MO,�>�^o[�{;�͑���q�ǽ��
x�� �	_���]�o����⇨w���:(߃��yo�w:zOl)F���>tl�l�`#v'̳7Rn���$\�r1���IPq�P*9+�歾9g��|Y�u�'�Oi��i��{x�<2��_c�G;��MN�,�\�H�
CN���ޞ�u�1��S��n�K�^
Y�2(�@�go)�6��(\�_ݓ��uD\�_�r�}f2����=o	 '{���]dSL�)i�@-ufh�nEH�Y8ڻ�ն������n�g#=�uMαh��f�/ny�uθ��b��P����tH����?Mꭷ6�0��̸�g�m���@�.�u<{��}_ٺ�W�d·��%Y�+��x�v�]W7�xn�ѡ�"�cL�귪����׮�[A���t�ӕ�X���k(�ECH�mM� �ه��р{N���x���C~�]�Y�}8������\����u��}��c�R7��T��,�1��L�ɝ��M�Jgbуrs��q0U7���}��K����DwU
��D��[�KZ�Ow����cLb������_�� f�
A�v�5�N-NL�t-���A�cR֕K�b�J��ƈ�h�h��[ibbK����L̹r�aZ�J�R��-jDT��[ErŨ�Uĩr���Pb3ɀ�Qb��c��K���[E�Q1l��fUYs��(��*�,UUDQp���T��mK*�4n	mZ��QEDQDkPXc�e�q�1���.\�+�l��)*Q��E[�\�A��[5�%��VV�e�F2b��ʈ�E�fe��Ҷ�D\j9j��V�Uj�L����UKfabcc�*b� �(̵-��̫Zۈ�6�U"�KK3(�̰�­@��.e1`��e��YS(UE�0������Q��\���PV҃kh��ָ��A�L��iLf��R���C3.2�X4�s��,r�3-�3-¢��T��imbTm�L��D�PU�2�;��=Ǭ���-v8�땣-�"��������wnԻ ��؇��+(m�6�C�\��ƶNU6�3ѷ&�D�k*���r��Nk���	��zۍ�1ɷ��a����-�к�s�����qBN����qճɶ�ݷى콬�un�˰\��,幺�m�kl�l����u��S��8�^Z��ۂ����C�i�\�1[�N��=^�[=n:�.�+�ݺa�^=[����[3���È6%ѵ�]vL֬ر���P���1��n��utKY�w��������q�u�1�
j�n��1c�V���v;��."Kvś���9��W�N*��Z ��1c�|��V�������ld\u�`��PgFyᭉu�2kˡz�^��@�Vw���|z�����.{v���g�bG����l�X:�t6��������,jNυ�7��Z8�E�^�Cڲq͸���簺m��۸���mN7f¦�x�Ûq��I���v�� ��E[��ѺE�=v��n���=ˠn������=�[f�M���N���瞴���vlr�FL���(v�WF��=5�.7.H�oU�u�pf�ڠ䱼����1��kÛV5��/YB��Նۓ�D�[�;sȻ��=2��y$���dw���rc����q�a�<E&}&��4-�![�����n�Mk\Il;��n{{rڳA�lv�Ynxɺ��ND8 y��km�s5X�ؗ&�	`�ی]ɻ/L����[���g��n�^��gW7��7?8`��ۋE�V����1��S�s�B9�3���U���T���{�:�:���3d���=���=��Ʊլ]r�30�����gz���ۗ
N��{u��N9털7���m�*nK��y�q���8�O'�lu�Gn�X:`:�y�j���MZW�͹rn1���2B�瑗�F���$�\�γ�x�g�MEm�ۦ�c�A���ke�;��8�a�Iܘ��2ud�M`��m�^^ɣ#F9+n���O93�i�{s$�᮰v2��;i���6ڭ�9��/����;r��'-�n��4v��;7�n+��ܽv-��bw3����mn�0�<њ�t����x�/Juf.��7O�-ÊN%�fQ�N�mp둸��չ�&��ӭ�ax|ݰ8���8�v43�W�M֬ŝ1r��T䵑��r�z�^u���#�v�8���l�x��ni"�+���w����?�!D��!D���W��,�D����%�ם^nz�ݞYy��>���˻��>�v# ��B(I�fd)`$:s*���|�O_$+�ߡ �r���d�����JtdLt���+^$��L	�RȆ��]eԺ�����X�Su�?۸�c�ڥ�F_}�l�[�����)"����f�����J~�@u���@ ��k� I���q�Y'^����uw;�yAn�	8׶�H1CR���V�{���vwX2̧.)�-������$� �wj�bAu��W�E��7��θ��}���싵R!]�=lk�j��r�3;�m�㮺�r]��+����>�}7<f�f��K�ڤ�6�ݯ���3���7��5���ۿR+�/n��O4GD�V(�X�����2Oc������v� {�k�^�����<<ϴ{�����mQ�z1�����?�/�:���n�S鋘�ɞ��(��վ�  ;���tY�U` ۝�t/k��VR@)Y�^�
fB�v����VgU�cb����O�sP��m�z �{j���yy�m�M�&`I�0��GBf�^WWm�Ǖ�� .�eU  ��ګ@ x�7�W�����!s�!^uU}A�l����,?��}&B'���|y��m���� ����@ �/:��@}���q���9�#� I(����bE��QQE�)��ĝn�nY.ֽ/8��=���ߟ{0cb�E��ު� כV�> �f����5���!]�UPπ]כw =�}���~�s1L}��/��Wo����5ܕQ�	 ��:��@�v�xbuI�ۯ+�뿨�Q�"�%H�\�#��.� A�w}.���XU�v[���>&�Y�\G�Z\��nˡ����޻��F�w8���ib���":��<|�]`j������2����-��c�wx�H�������>�D̎UP.��8�I�Sy��S�@|����� >÷jib1�mE_Dɵ-y��ݻ�'�LKQ!�H�[u.� 1�m*��ab��IӬВ����H�好��PI��݁JDq�x򝚕�8!E��u��I�㵻v��x�[��m�Eu����-�Y���7�PҒX�I>-�zL��&y�I&�Hj|�I�鹳T{k�t���ۻ�nU)��Zq Ј�4���_ 'm�z�㷷*Ս�f��ń�	/�]"��jf�=%���9�|���O~����\�z�WUH qmغI ���;�ہkcw��K��mX�'K�V)��D�*$)R�ɚ�z��E����T� >��R 	4۹�A,��w��)�W�l�N㩦�E�4}V��c[���J�ܯfr��<�I�Ώtd�<s�݂�qLz߲��ޣe��.�K�� \eU}!�	�,ϦQ*eJ�AΪ�W�]gm]�:~�d�\�@%u  ����"�K/y�Us��q��u�'>��3�xc7F���p맷>f]�=��c���Қv�"ጘc�J���q1-D7	����+��>�ǽ��x@ .����B��{���h��݉Ey#ŷW�K�&(���u,AjE�[�z1	.c�<{�}�<��{T�@|ZwmM| ]gmSm�6�Z�U���{dR�m�aDJ�M|����|[�V�����&z+���&�s!��s�گ@^_m݀��=��_��3W.���������~Cp�������j� �3i\O����kλ���`|s�ʯ����LD�����j��컻 t��)3~�ɟ>ݯ�VU�M| ��wh8�Pggm<��	��9&��^V�75ӱ��oݧ��e�N*|�� _�	�-^B|~���歞���OS�|�$����g�Y > �`�đH�V��]���KNV�� ���륞`}��[,�i�)��Q8�dn̮�����.�n=;;P:�d�W��Ӏ��͵��u��Ú�.�[��[��j��m�v�g������ݪ��x��5�M�6f�ͫ	)�t�Q������g&g N�d�Wg YL[k����.�z�c�;�<[\��^n(x�ġ	ی��|vyC|{r�v�ܻ�\>�L�v����S͖����~����S.	�+ߒuWJ�ؐ^�m]����6��h��ԣ/���9�^�v�n��.��H�đL*��S��N�x�}흇��^ 3ov��6#c��I������g�S�����J�fDL��f_��ݻ�����@v���V�/�k���$�H��u&���������QSAO{�x�ˌڗ�{}s�3��W�� ��ښH�F�q���Q���������IS.�'�O�*f*�}�U�H�^����L���'�/�U�]�`|k�گ�0Ia{�t���]-��v�F�qUP�&�),��C��޸7<=g�G�ӱ�1<�j�r�=s�V�KIW��-8�V-[�"�ߌ﬌7���� /z��D<����^t��s3���@�6��NYG�ʈ�.�g3,]����9[EF����s������ZCg$�o���7M�kd�`-��r�DNAsS��A9
y���L8��r��W�w6��� �f����n���� �b�vz�Y5�� ���K��䂝|k�ږ�$�z��6 �ʏ{f֨�̼@ �}�T��$��z\�.-��L�H�<�#�]�DƬ�QZ���.�whe�_��L�:�m%���m!*��3���;~����]ja,b�0�4���T�a.�n�]s�j!��e$9z6��@&	���	'%zHLm��W������{t=���L�]P'5Íus����$���pٮ��h�?7��=��c7������uK���5��*���^Wmݠ	�FPT�7\��Zg��Ԋ$���$�2:a	��11&f��{���O(_[�s���-����@ 0�ښ�>��ۻ�\n7����8w�R��g,�&}șR��s�����w��W`�[�V�G&���U_A�i� f�7���}$'�Yvؙ�7޼�n}�x��Sǻ�ǭ����^ڵw1���OW���DY�qDI�bsH�;9�m�< ǹ�-�+����E�Q$�p�D�S�s�ڪQLU;US�������z�4� f�m݁��͢#��$�l(���:~�����1l��
eC&
u�����I>_s�ǻH,yJ��^7���ۙ�M� �ٵ^=;���}�߿þrv6S�N�U����˪,��wuW97(%D�L��m2S�廩�@)���)�u*��ͫ��0��L���E>�Mto�8I��I	Ty(OTq?L���"u�/ r^��߶��
c�#�6V_UR [�ʱH��Vy�)v��5����0��L��&\�Q�˵`�5���W��@�y0�mW��� ��g]� c�گ1��SlP�&eJ�:��i{����gv�Ս��n���ؓ/��^!�F=|6�̮oVی.ߋO6�nLպ�������\�XB3eWXq,���8w�#���_nX;t��l\�y
����ު�#"�D�."$K5N��	/%��uQOˮ�u���Kuo3 H�姛�&�I&_;�
SP� ���O�
�Y13�2K%�3=<5�sͭ�{�����PpJ�GWI׎v�|�}���F���/���� �_nz] l_i��5�E��^�'�j����ݗv ǻ�^�{m2\!D%T�AO{�,�U{G9R�s]u�"I@jonl�,�u~�IwT�z�dh����%�� �Q��ș��(=�w�D����]��ڈ�N����w\V^�G�n�R+��{j��Y.12�H�s4Ξ���fo4b�nK�_��6.7v������y��e؀)�uW�Ҍ�` ��JKpϔ$�m�96ws���ػ.��$�|��"�[����vd�A�Nnh��y�q����c�J��ѱ	�մ��jb�0Sq`�sV�g��{���	�+[ ��@�����:)�Q}V�O۹V�q`ҷ6��E��{s؃5�nm3��y��:ב��/=rCS�9q�]�s����Z�$�1�ݹ���η<�'� 㷶`�m�v�2\������R�ԋڶ�o7�-��cv[��nz=J��s����u��][)���7Q�p������g[kX٭���rl���0�[nPwNŮ�6�4����)j.��O��7ϟ1�	xG�\�ϝ:�v�Y��f�u�	��Cڞ|�pݞ�^���_v���\8D"H-�E���u�(���&�~l�=B{Q��Οo���Uxg�|s�گ�Lǘ�dp��pɂ��euSԁ_E�hu��=�{�  ��ښϳ3:��A�Q^�b�ȏa��;��+v�d�B�J����wUy��6�����"#:�ٳ@�[�گ��ٙ��vS�|�<���eL�W�>뫪��]Q�R݅>�Ux���I?I&����r/+�Z�ĺ� �t^�|G�.��IZ�H�A.g~ײַ��5�o�x�}�ԧ��j��_UM$ ^fm݃a��j�_E�&V�<"�ِsD�h,�.$��C�2�!147n-W�խ�taHW��i�dg������~��e�*V�N}]^ �Ϊw�	 ��ږ��MFt8��t��X�(7��1%�$�p�$��k����t��g,WE���Ǯfd�3uЦ�9j����z�N��sN6���CR�r%�[����-s�N�iξC�t�sТ5�o�� 7�:��6$c�گ�6�ˮ�U�7�]����1l�AC&
tuVmݍ���}K�g��A���6�ɳ2j�H�y�v� �ٵ.�w���j *��
{�/�w�d�of�h����`>��� #���*��w5
r�6�/�� �>��'�3��^� �w}'�+U�ai�W3����a$��w~�I:_:�R�̂�,b�1��玊lA#���)s	ƶ�.�;v�S���[N�uvwj�V��s��������$��3L���6����}��7��/�,G����v�Wu��'H&[ۗH�E��D50DʕT�W鯀�c�z��knw+,�nT� a|��"�װ�{E5�{L����@̒��QG:��^ ��U��Ig�m����7%M>�TS*�W@�פ�����_�坞���bpu����z�w���ӫ���6{�'�C|���gl�����uֱ�\���#q��Xf�g�=��+���t��^�u�Q��ЧoՆf�({�^�����X��X\��� ^Ei;j��[
򀓫sۓ}��L�%�o���d����/V����C�����M_��N;�w`���
3\�j��.2Fnv.b��i79x�&D��h�7v�ֽ��q�b�3�k��;mW;}<�W�6���������Y��6�Q� �X�R5�퐟[�"�m�����j��N�KH]Ș4s���~�����١�K��7� �0���c|q������ɢ��n<�R3BQ�b����17��vL1�<��]K�u��]��T"V�JMN,�`Y�ZxT&#2-_Ʈq�}g�`FV5qO�J��(�[�}����n++1޶{��@�{�ݗ�N�h��^��w����O_�,wY�n�}|�v�����Ǯ�{Q| 8*{<���{3�C�,M9:1�J��9�-ͽs���e�7-�Ȋ���ڸ0)c�19��2ܧ�zH���m�����NJ���@/5{;����Z����7^�	��O}^�N���4<W������;9�lܺ��"��8r�(�̈�û��`A����=�ˉ�w�9�/6���kI"@�evi؁�64���~ưh���°zN5�>���n�]�ۻ&h>�᭏`��z3�2����T\2��2��sJ�c�E�+F(���("5�Svܦ�.C�N�m�π� ��
��\ql�+2�%�+Z9�[n,2�P���ʔL�T���B��C-��V��+�\��Z���`��գk�m�bfL\���",Q��S31����L�ª�e(�3-�G1p���ZQEj��J���%�ah"&Z����"�U33*�ҹ�`�V�1�Į[��-��KfP���V.R�Z�b�[`��J�b5���E���m�eZ#Ul�%qƵ�R �F-��EI�i��b�h娋)E�-����EZ­(�UEĕV\�.4ƤE��iL�%nfc���e�r.c[�f
ckLf&,V8��%m�Z�k����U�
�QZ
5-S�3�`�2�(���-e�Q��r��I��O�Mp��U� }�R�$F=�����+s0�3*Lu�{�^���k�3���I��WIy%�0�ښ̬λ�l�_�@�����g[LQ	�9U-��v����.�z�b��6�K�%�$�噷$�H&_;�E$���y��5s ;�ɄEW|��~���ʦ�ki����;W�S�j�F(�;f�v훺�]�v�?7߼���3u����{uK��A�wiW��A���W�om`y=����Ub�A%��y݊H&�߰�+V�GV���w�Y'�@�w����LS���� k��Kt��ۻ�`N9V�g;��ČLO��D�"��U�i egmS������]x�����3��y%�n�R$��;�mOFP��." �D����Ք���(���^l	}�_W��,�ݻ��@���u����	��ut�ִ&�Q�4-t�����.�ҷ�����@�SVI��{
/n��i���x<�5�*T����I<=<���#"�Ih͘Vm:�y�H�y�I��TsUsHO���ŕ۷v��ە.#k/Ȯ�u�!��*��"'ҁR&]f�ٚ�{F�e��7-W\�!y��]�￿~�L����U�|�z�U�]�Wc`c��M�]�ﳺ���1����[�wZ���`8�.T��|CA��M��ٻ�r��㕕/���<�	 ^5��W� �¦�<=�D�/�o|�Y�D���a����wa��w=.�	:����}�s� 6�������/�l�?2F�"aJ�~��I�*=�>y� *���X l_i��-��"��Q9F9���y�N�mݠ�B�\����R8������� c����bfBfvK��������y%�ӯ.I&����Jn ���s�;nu�Wy �h��7�&'K[��l]	[�g#���3�������=r��<l���M�I[��wS;>'�#[R��(�:�1ٸ�r�z&�t;zܰ��9�`��W��q�[vy�v�V��Z�Pgb|OgO�z�Wŵvwgyc;���b2�/kR��#g�+�p�<sq]��D��l%�z\v��M<b�6�7a-3�{��M����/�z�8��vVrn�m�\N��w[+vk�8�Z뢰���#��5��ج[���Ï\�]FWu��[vpN�����%��^w���1p�5�ΰ5�{p��^[.~&eC������`�����/  Y��-��=o���z3�T�|�:ꗃ�c-�Bhp�*��
y�U�:|�\�U����;@|[��QHw�T�0&I�ت��}}>�{_yBw�ʙ��4몐��]��x@|�u}yy�z�z�P0ۨn�E�Ϊ�#5dr�d���a��"+:�k�]'��>�	� .�w�H|�q}�4 {on���v��w����6�x2&ي~d�A.URwWJ�|�u�Z��=�$��5��m���-�;����]�v�{/���=m���H������ҍ���q��nd�x�^ןFH�e��bw]������k+��F�E���� �c���W�� nu�݄��*�eO;$���E�UU}��z�����
���ĸq0S����������|����D�-2��=g��8d^�`�$���љ}34.{��yg=�����矍<�]����+�ܱ�/|�WN1M�3��Y ͖���q8@-�w�� nu��m�C'�N=��S����IP�xD"��(ȹ&��b�	�^ի =��97D:jp-��Kt�[�{v�ν��%K�I0G�>�ת�|��Ǐ� �o^f �)3��H�W���2`$C��y�ػd�dĐK&�Q}wv6|��n��ţ�=�Ґ�95wV�(7��1$^L�wt���P-��u[[�;,����s��5�<&�8�[$�m�ϯS���gO�`њ��,��3*#�L��3���$�\�~@��uT|��ٵN�Nݩn2��(���S7�D��Q/�$�k��$��E�Rd����	��o�xm�ĝ��t�����swj��5��R��ڛ��~�8]띵@�a�˟�$�::�r�� �wԼ
�n'�C�lzE-���CoM����F����A�cμ����N�X�O�Y:�=�qk��Hźݳs����j�O"2�Ý�9U^�fn�U����K�f�R2��g 3�~｝���j��u�[ Bh��M  �3��l���G�'�V�nR_��	9�}ٸ.�HԆ,I6t}�o8l�nm*�x^��o�t~�@Mu��v�9��Kt �3������ˎhr<�����j�p�\��s��[��Y���\F�q�9�9�Q���H_߿{��'3�.���E�������/��3�ͬBu��ta܍�ꛛ�o3I%ŷro�l�?2@R�I*�]5^��w��Nм�}PF��� �ݩn� [�����F}3Q�$纑՛�y
ܐ�8 �d'�#_�j���mf�UP D�G^�Ӆ@?�ʺ�[��n���� �3��"Ty���l��"`�H����v�n1DJ��ߩ/���3�����[9/#������s�T�z���h���֦!<FOS�s����/$Ȼ�x�e[���u�(S��rK�"�ԭCڭ�2���G�����1�D����r�i U��T ��Wc�y6�TH/��^�먤|.�ڥCo3;j��LNȽ0�NYȕ!0�qy���:A���7lpݵ=F{�sm�gm��~~sۡ��e�S3\�î�H؁n������=˪����<1�eR^ �{j��cWlL@J��,�s4Κ��Kë�n���l��`�J�Hc�Uh��ګ %���}K��"���D�1O̐�J�@��t���A���j�σ�u1+*��'J��\g� >5߼��&���)�Ѐ��[��o�ڨ�U���38 �Uԕx@�z�f$�^O7`�܊pr��ZIq���:��r ��ԏ~w�&d �wԼ.���Ƽ�m�\�Q=�4�����@#n�}��Ύ��Y]>��6,P��[��d�zĘ�4"^�b��8�r�ޖ����0qR[��d��޼l�n��_��:)Uf
�%;�ܼ��Qr�������e�n%� �I���qwTq�7���9��'j.�@�:箇T�Q�v�RTK��	��qs�n��\�sbf[v6N+\k4(W9e��[ݸ7/z�k�n��+h7�n�r��ت�;+��M�vtG>wsl\�X亥^9z���m�r�m.�Rn��V�m���iM����q��m�q�u�q�O���NͷneI�>�������Peݹ.���u��r
0i��޼�jPCە��O3��|��V�ݩ��4�+�P��h�Vg��"�K���3Q�ЀwA$_�-L�ϯ�$��(:���o�	���m�f>ݪ�xm�Һ)FY�>~��^�9i� J�e��&j��_]�`�A�w}K��3�[p�(�7��ٝ�w� �v���&Ô��Ba7��s�X�\u,���3\��u�ڧ �SH5�mmTw<�ɾ�m5l���ۻn5ے$MD11j��wI$�KK�~Ev8,e_�^�^�� ���P�^v������Kz\�
l�b�Q�H�M�E���kn��Q�	rC�>y�]��o^���7����n}����"�.� ���T ��;ji]eEve/GJ�TZ��ۻ� ��j��q�射�!�*����RU�.��s�68'Y�jV�5�����+u�.�.\�%�)�}����s�(�Ş�V���H����"z5����P�=�u��壧3��V߶�X�O���I�;ή�A)���G}�F;;��Q�|�"�?L��
;��� o���x:��^�Ǿ����@$on��m�׽�.��6`d���� ��#����W����B/n�֒D���si �Y��w=1	�״.���D�b��K%G�Ī���U���^s���s����}�N?��d�ğ��ݵ^��2��1U��#b�k!D8��M]k7n{E�â+U�,p�4u�wh�b�5�y�,�=��I"D�Cd�g|+��W�-/��t�A%��ٙ�ޮ����;1&��U�E$t��_�%����BB�Js߭6��R�Ղo����^խܓ~I;�ٙ�]T:$���-��yEj��>l�ܪ��)�u*��A7��+��K�y`��jN��؟}YS�D��f�ݞ6+�T�[g4>[}UlOw	dH�0sjbjU\H�^����w0�ۊZg�kb
���*�2�4.��ڐ6��o��s3�� >�{�xȈI(�H��!w].N��1PvI�%f��x ��]� !gnQT�2���Z݀�u{R��N��(���	���Ϋ�v -��y�)�~����ꩤg�:�� ,�ʪ9�xE�'�7����|��f��W\�\�u�}L&LOp
bwiƺ5�vF�:��>�~��^ͧ>&V�Oޮ� �fuZ���ܯW�T@��=~F��^��λ��E�D�"j!�f	�B�^W�w��Q���Ny�v�^lA�Y�V� �v�P�����b{F�ҡ�}�J!P4I��!�'�|mVmӴ���: !��ޮ���!����ɒp�����	���U�Eb��>lPܪ�AO��3=W�3yр���� �O�v�@$����ze(*�'��n�6$mY�J�V[{�/EL[�&�L:eM��ӛ3������z75�x6lF,�0�o��8�6�����O��rHI��{�xȈ ��TD�!Gu�*�H8�v�GIɢbU$�^]�H�|�_��I����H<��4O<�U&��R��ۇk\�[uh\=v�ܝ7`���p�nؠs��pWf��]��0șh ��Df�ݫ -��W�XomM��^�����F��λ� ]���H�N&H#�bW�9�����\Ok�լ��j7��X��.��z�#��/HǷj}���̰qgAJ$ML&L�4RB�^�* �ү ۅ������~���� [۵T1�1�mW�R/B�.=1b&b���{�3���3�ܒ�zӘ �W���Y��5��λ�����3�$�ݷ~�й�$�9M|����6����^���S�q;��ύ{�U�� 3/:��1g�����m�W|��۳ӃҼe��.�r�Sl+���me;˘�:�C�
a���,4��++k���N//��+^,���~����Gh�v ���ΰeǖi<zG���a���(,K���.���^�۽��I����5_o�)����yA��&@d��T���h�$:��R�y�\��8��ny&}��X��,`Q��p��z9�퓮���tE�eR ������혳s�<3�{�P��v�?>���0n�&�rH�2'�]1y�S��6���	bY��޼f���j6q(�� ��_.��nVOu�B!������T3Z�Y�ӭ�R�:)��䪷Nqwߵ����;gt��{ժq�GX��5���ۙ�6�TSڜc%�l�z׍W��Q�7n��K�ʅ�vQ4WŤO_�y{�{�Շ������ҔΙ8��@7:]�a��Թ'����`1x��|<օ5u��=�Wt ��Z��1�ؼ��E��p���%����߄7��h+ѥ�)�:k�|�㶷:��ݛ\�~~�h@���F��ݝ��򨙃޻pO(o7`O�{zNy3ook���+Y���zw�.Ig��;���g��^�C�
�M��lC����߳�!jgw���T��I��Ah�.�y��vI�e�w=����!euM������|U�����0h��ꬆ9��Q� �f�v�dZ���MFV3{)U7A"�=��:�^L��JdK�
4,vYW�{�<]D���!�Dd��H~�{�9yE�6/WV;O_t7�,@g�]~�=���*�T�"�S2�ŵ�1q�*bR�m
�KT�QTij�c�1�L�[�e�+-��A�,�-��r��Sʕ.1ZQq�n`V.)s �#m�bԭiZ�.QF�R��[Ln"㖆1T*�j�2�\qf��lC#�e
aA[iiX8\b�ڹm�Ԯ5�.Z�1�Ek���Q���DZ�ImX,�����[K��qY�jf�V���6�Fa�\��1n-\�Q�q�fe�-mQTj� �-e�+\��YmW�1��ŔE�+P���TU��F�ƔZs"���31UmV��DRڕ*UR���bff)TAF��� �#�fEJV��9w>��q�;m�{`ǁ�[h֬�Q�����+R�J�
�a�T-1�U��M��&�۶�; r�	jʙ���S�
�UYK,�Zb���[U-e�qYr��rԪ���JZ֫VZ6���Qe��X����\����`������6�l������f�=,�/[��Y8Mݯ[���V�s��C��7:�<�������۵r��n'�\�8;���F���m�n0��Pŷq=�ϰ�uٲ�/>4Y�a��CE��k���)���y�'6y�S��ct�+9�F�n|�n]n����ӭ�=���2<&S8aݍ�Nr���l��u��e�h���۶;^^��@�\-�-����Z.�������^2!Mն����z��0tm\X�m2��w =�mp�',�y�ٻ6*�m��7m�R���n�	g�a�pl�XL�mm�s��o4�������v9=����mɻ>/E�����/�8;n-�c���l9��ٰ��!�=6���pj���>�ێT�#j�=<4��7k�nn7=��]���k���+L;��b��m�m�$�V�v�έ��o'^��HO/SJ�\u����)����:p��\q�狵۔�dG/��y8��O����nK�n8x]�'�w<�<�Z���y'͝�S�k�����nv��������;Y��{�5�N�ع3ꎖ5��tON��%�;�qp���c�q�Ğ��n$�c�z�����<@�8���d����R���{a��X.����;s̬��⹎ݵ��+v+��\���V}��h��X&r�Au�VϯGZ��awh:�V� �a�H󓚄�����/!z��d29�h��<N�b��ud�ۋ̘Ǔk�D��޽+�����(�L�錙ƚ�8�m휆�]i�����z�����Y�\�b��׎M���۝�[`0����E����f�c�`�c���{':�I�{9�vmӎ�u���d��ح�E[��9�܇4V�'>:�N{�vd�{�p��\�Y�̏���;�#��M��;��E��ɓ��-��8<=Yx���ix]8�e���oEג��u�7b5��n�ܼ�֚�76=%ïU��0V��;T�+u�Wq������\ë���4�Kk���r�v۱И�읙��2�V��<�Ӹ�:�Vm=co$��mo�ɮ��[Q�)՞���5�G	�1:�\��t
���d��#���g�9���s���ɳ��n�A�;�g�U=�N=�,M����v���یx�Wp�+��\��9�/:�w]��[,v��.�L�.�㹻M�un#��EGi�{F���#[fg�WUn��y�rb9j���\m�z�]�v�w��q ?J���C���@޽���6}�{ٙ��Kz�i��sq0��L�eؤP ��^�T�فʂ	���i�ު��\����y�w��� >�s�h6Ͻ$$���9A<>�I�N}��ښq28��Īo\�]x� ̾ڻ�z�Yq6>ͩo�{�^�gm݂�:
Q"r���y�9��k۝1s3�5 �sݺ� ��j� �5����;��u0N����I
�h�L(����FϻnՀ��=^!�vMXyەx����nI&緞fy"P	�ݻ�$�@�u�Y��Α�I�0�
D���f,�n�T�'c�-V9�P����/=�ߟ�����7
��=��^ A7۵X ��S@:Q]�ɳ��y�T�0&����^��x�!�����/�}�U���h��u�V����6��E���m��ݽ�i�����C!`V\l���N������gY�yS�b��Z{�%�ڨ�SuR��B�N?]�Bown��l5�eR����9��t��Y����zHJ���D)���2z�����<{RI$������λʸޖ�$+w���@#]�U%�K��N&G��x&���Λ/C�L$�����H�9�rI6������<9����	!��.����R�.L�QB۬��BIi{��UY��t����K�/f���^n�E�Ωy��j�qV'Z�7�nn�=��kpn}��AQ�wK����n���"a�cr�Vj�Z���
$���"/۷j��m�z�-�w����q��b&;q�bK�/ ����:&
�`A�no�Yo�] ��QDE��$� {}��@�c���Y�
���^ʞ����D0"~�q>�(ު�ZA$����&��נ�W,8"��N��9�$�N ��AOj���mw�����[>��x{��9V�ф�^C<���}�5�����.�~�{��f7�$.���C���W�u���)O� Lݧ5ٕ�M�2r|�HK�����w���m�]�EZ��Xo����_�uTb�A�N&G�M�M�o�y�jƏrׇ,�x�I�^ש �uCu��y�v)�������Y�t�x��C���������b#�B]�,nv)s�F�s�����Ӹ��������Gp28Ӌw[R��uT����6)ҙ�Ƴґn{*[��gUH}*az-�q�"$�_�]v��g-��5�����3}�����3jz�H��#E�9O$��{F`�&Mi�U-�=w�V�> �Q�U�۽Yٓ��gU}# ��uݠ�{1b�O�A>��z����(�[�#�� p���@>z��� �>�og�%|�Է(Ћ�_Bs���N�$ Ћk\ʽ��	�9Y��<r�Z��`�=��j9L��c'"g!"�G�ߢ}���[y��\>�I-��9ox{f���!L�>�vw���q엛������{@y�����'<��g;.���z�<�+OGkO����1s�����|��d.Ηc�[Z=>�0���'l�@�!۫����;�����m�7��	 �<޼��/�g;*I¦"��Rp�5C��ùQ��B($�f7��t�DK��E�{=���#�a�儛1ت  ��y�w��}u`R$���1�A�ّ�D%AI��d�ĸ�&JtN�m݇����}���V�Fmj���O^�ݤ �}uK��Ҭ�%
>n9Mf�;�O4nwfk�I�{�e�$�8�I-�{ΰoa��ٳ�	.��3�\� �C'�0��^��� �cj��]��]�ָ��;w��� s���#/c��*�O"}U�1f-�g�|���9���3[)�����ň�� �Axޡs�8�u����54n*iBT�֓�"�^��q4�4�FM��)׉P1"Z���c19����qk��FCc��lnݔ��v���ҼG]��� ;��Z�M�r���n����݉.+�㪗=uݣ��=61�9��i��u��q�� pX�E����ջO��Yb�<�����"���[��.T���E�mEi�>e�wl�y�k,9�l�d�"�Gn�9Ⱥ����6�|�d\�<N�6w��w���	�'iƔ�Ii�%s�<��=����4uhS�{S
$����t8�`D�D)�{uT���o��^�QAYF�����V�U7� ,��󯍳��	�HD|�%U|�w	*Ge�n��v�H�^=�.���2�:��&rK썸؎������Ȉp�����ey�^�RU��L����x���l^�U�:ѱ!I��dǐ����d�����f�� Y9sM��u�U6�kj�&��8��̰O��}46�v�!�0 �6)��d�����uPrU�d��{�O����>$>�w���ꈱ5iNiǾ��Wk��F���W*��f5���_S�g���c���~�������Ɲ}����7v|O���DbB�`�u.9{#f�白v	qN�0�O�@�.'�I2�',w dufU�7=��7&�ش��#��!��uj�Q��XL��q�˔:�l�_:�8�n*�cv�:�=���vAI�^�p��1�� �O��u� �7ƭ��b2e�v�J�)IbE�yv|Iw���>$�;ow{���Ԏ���d�)�u�$l��-L��!ʊ��*�q���V!��}��A�]w�$��O;��$;��B+"$�s����$Wg]�0�L��
f�z��H$��T�5�;ӭ�s5�oV�2ks��M<�b϶��Q�����}������M���Ƥ�
9�������˝�v���}��9Q��c�s�b��J|�H�os�� �k3z���I����]���av��{b�<}B�鍊��AJ&J*D���!"n�n{�'��,O7��'�s�(e���L�&z�wA>�����幩ss�����"�'���AA�
m�{(��yOLn�b�^P�)2�ʅ�-β��������=���g)���JU�I�/&F]v�F3�����\�"�_(fFmcy����gY�ݏ _ޟ<�cF6D�R�����E!N��G"ꟈ�{�d���$׽R%ٚQ�9�f��2��AL	��#�6�H:�zń�x�S[��,F��P$��Ϊ��[$ψ���G`N�q?)�T;�.�Ӓ�O�n��ݞ!f��4�ֱ��0M;��=uL�S0�P�E�]�>�u^�NooU�C�w��E��e��徭�X��B<`(Rٷ���5l�9`��*q<�MU?�@$��"��{�~"#��fy�gx�^��	(	D�EH�V��D^���%G��ɮ�Y����f��@�c�	�!A��mL�EU�QLޝ���GWmQ �H�s޻��k�����t�I������;��!MW\�LQ�Q1���s�	ӵ5G�D����cowY_����}ݖ���'\�2�Ѕ8�� �E�U
>9jcQE(�H3(������΋�Q�s�5�|w)��^i���jr�} 刍[�\������1p:L��ty�s6�޳���Ѧ��*\�LF��\Ȉ�L(S�W�y2cޱd�	����J�)͞v�ڠ�c}>�x�݂`(3e�F%�(C�v,�v�FH��� ��W���vH3��61����w\�U�R��
�vn���$�gw�_�'�Ъ���]�wKu���/��A"_7b�Ll\� ����^���۱��Bk�ݕM59�ՂI�}i�"�gL=�������b��p& ���0&��u���I{u\�qS;7n�b����>2��X'��}uQ�:��M\�՚&��r�r�ڍ�l���T[�W�u���D\��4�P��x�w����W�#M�Rw�̸45�K�%ϩ����s�=>]o���.��s<�+v��\��y��خ��p���Z�㇮�kv��ٷ(�TmoG'��p����(C]�YQ��� �C,m�'�����9ϴ�u�p�f%����r�[�����qk;n`2���9�;tۡV�nwL�#�˶���sR�n�tv�q���6�������M�#N�]�wes��cg�P�6�@-�S����y��콲n�\S�q����Ӈ�s�p�e0])�T`mL��17Xf�"\
S����z��Ӻ�_�>�N�d�5�6,�m��� �|��sk�����&o�u��vR��6����}w�I� K�v,���=�7��6�{+��&B�1�P�(�$�!P廰A#o��A��8�螜���L=n��A}�+*�t�"#�)
����7v��� I��u`��A��$.���x/���^v�Y�K�%`%e"h��U�(�A��wq-�u���G(L��+*�I ����.���;�ɬ�����O�FA �A  (�;�����c�;�K�\N'��mrv��M�o���>����"��6����}�q �}U���*#`s�� �} �gp����$7D�1"����d���@V*⳻��\F:���7B�I��3��o\f@ȟC{5U����n䈵2��������.�kҫ�%��0r�{jU��:��}Z<H$��ɯ	���,�Gfu�%�z��'bӴff����v^�A���d��Ί#m�����:�Ur��	"$�B|��0�C��Ύ�z\_n1XI5�DH��w`��{�iۼ�/_ H"w]VU٘DG�
B��;�������܎ҥ��Ý�XH3���'/���w��{��MZח7o����u.�����O��j��m�\l���l�^8�%*e�������1�S-�S�{o�(�K�����w��:�x�eq%T)�-�^k�'�OW@�$�I�������$�Foj���3`Q ���v �{�v>;�K�ɸ����|z��2
��$���/�|I���`�}�˧G�gfp��%Q�u
#!��ݴ@��5e���{����n*3w8����w_�T�=�y��b�":���3��X����ֿ`թ��μ�g+��ڐ㊵��͚���Ĳ��-U��q�v�M��Bm���.��π�-���O��'����qcix'����g����\�`C|t�����R枕�}6��}��{�������M=1`��K�y��c��y+0�<����~�
W<BZ7�v)���޹�"S6{4I�n�0xn���} �h*��8:��@f�D8eX��{��z�~����z�G}w$�3�2egZ��^ՓW�+f�9�UӸ�iT����ue˾�!{�W��ۼ�3��.S8���j^�}=�ɞ��Ih�'0��Ӝ2����@����j�,�:xAÆ$�y�W�ڝ�M[-�x餇��S����[�������!�^�^�����3������~z�S��SX����2�|tgm<�y�Ӌ��=�b�8M�,��]��{�ak�.G��{`��ܣ��awޫn��ŊY�(��0��zc˱tS��Q	�P��]��o���g���o����
�x�W������"�^4xO]�A^��+�y�G����!H\$�N����T�2��=|�;�>Z�Ov��)���M��t>��[��ݹ[���Q��ҥ��C#E���ٯ;69�KŸ}:�UD:^���U��o��Of����}�=�D��Z�ُ��=u�n��ЈE׳6�N	��߷ �VQN��UjUլEm*Tq�;���g'lp��y%T)\�b8��Ŷ
�km�-w=�l��n�s��ݷc�ƊV1��2�(�����+V8�
���K���G+lUѣm����Z�qj Ɓ6!�! 6��#�mU(ҋ*Z�(��B��cR�s)*"���h���#E�ˆe�	J!DD�ѥ�J\�ģV��e�ˁ�R�EV���DJ�j�Q�q1+KB�1�iJ�A�R�Ī�9E�e�h�
-��*T-����մ�kc�JUJ�-Fҭ*��ZU�,-��ce��ֵ�jX)�����(���EkQ��j��#[m[m�J�%����KZ����B�ikXѶ�̡��Dj���KmV#bR��i��KnZakU��[m��-�B�UmAUE)KJZ��jUY�V��-�*-lj�$��J
1�e�+k(�.8W��Z�m(օ�e[*V���-Z�E�����jŨ��+j�UPD�9�I>y�v	�U��Z�Jf`)���5��,��1��H��U���z�O������sT�6��w`�P����0%A	��o�>#o��J�+Ϊ)6�O��]��go]��y�;��S>�7HC��@�ZF,�-[<Oiy�b�ݬ�Ukg��X��č���9�F=w�����3��J9��7��H1����C7�DGYٓ��ٖ�������M��d���L�dH��rI�@���SF��{{d�#�]�$��fT��qFz&�wXhU8=�����>�G�A+q7w�wd�@<w2��AՆt�]�]���=�VI>�̠$���� ��f��E]x�XV-��
�}��vU�|I��"�I>�������d-fb`阹g�_	�t�*�=�(�sn)*�4�k�crEAV4 ��˹��Q�]��[3�]�@ws���ʤ��{b`J�@�&n�x�mI$����!p�s��m�^7x���	�̩��`�=o�ϼv~�S�#�l�h!��� z�uK��K۴>�\]2�����+ݝ�;������yX�����vI>:{2��I>���Ҝ��c���\' �C�����!������S�uN�{{�������e6M�A>���uMP�V����I�-�L�L�dME��� ��wd��z![=c2FS]�|I%���>���~$9�:e
Y�D�;�O�q�Q���-�tݸ�A�;��[�S�=kA'�_��e|�R!n,/�%� �o���c^�����H@~��w87=�0�~��K����2DAZ���Y\>��_�ߦ;��g�f�
^$���jA��F�{1i�w"F!�,��˨��f�8p�p�s�8�"q��ϧ�*/%nXܝ���M$���pP�s�:H��y�s96۱lc���\�N�+��v��]��[�f�c��a�(2�B����/��yOlj���!��Yc �Y�	�k:Ը!�k��{q�׍��b47nxNg��cGst�aw4�<�tW���X�]��м�Xg��5�r(���;
�G�X�v۵�@�t�n/d�n8{uӗEa��훞�j�:y�n��\D��\Z�0%D�B/��@H'-�X��@;[�CS[6�V'k�گH$��}l���1�:Pg^W���(�{�lX�=�I>���`�O��z�čx�Ծ��|>A�������hvo{zŐI��udf��Q���s��I�|������)�B0�($�@��B��Xr�i>�IZ�]� u=��{p�}Kn��r��Ӻ��BJ�·y�߹�?|-��koW��Oݕ�o]��2��	 �۔$�Y���N�W�c<�:��LxDL2P�c�w�q��泧AG�n�v�h^������~���O\Z�P��*���U��|Y�ȯ��P�&nc��������}�����1Ajl|:]��ۖ�2h?=�>��M
��0Ȍ�0U��,��7qԘȑ`�4Au/FnM��4e�¤���ື-������A�Śp�P��66)M�y��>���߉$�nP	u� ͤDK&:�I"(�	J@QIDP�;�,��(I���l��I V��H�{2(\�tL�"|bL�vm�㽅wN�IJ���>$�s"����-���WDFC ���m�B0�!( �@�n��Iw��]�{�1�0���A�� Q9{�`�C�j6�5�:� �����W=���gN��)�$�Q���f���GH\�?$@@��[�}��v,Y�ʐ@'/_]���kQ-�F@�f���`�Y7�
�����������˲{�Nv_E�U��i>'����N^�]�I��E�V1X�E�f��؛����7q�5s���͏�`[~���w�1Ko��7tqLJ�/�˰ƋS���z5L/��ҵy�,��oA��T'y��N(��Gz��.\��ˣ5�U�T�o	̩�^�U�E��J�A�Rl�^u�ĶW`�15R|I>w�������A��-O$�tW�k�&e ʐL���_X�Lok���ˌ��8�����(���-8����a���{ǝywC �"����B�v͚�Er�l�z��aM��Tv9�[����i�L��Q �����@:�]���ޫ�;����ۦN^W�Oc�a�����Q·y�_6�}�w��{�4���}���ǉ5��W�@;ՐU��S��it�n�zI�U��*d$��ug`��<`�_��o��6yכ��W1oa�	�]�'ՙ�bä�7������f
����yv4|I{��� �)���� ����Q�>	��W�o}�;}٧O7$�"�j7v�mޜ���LnԸ���ƺ2Mb���Zh�ס��n2�m�"�+�2"�F	*@1�HUvӻ��OVP��j�}�u�v���A�=�	uU�����~�9Z\�Y�*��p15��㭱h�cv�}zE;>ӵ�������X��oϼ�s�>"�9Ւ#T�@�AZ蜌�������O7�Y�ҌX"DD(�L��F9פ���D��xu.wU��Y�݂:g��M��/�����V��H��P��W��vH$3�	'�qT*[����Mf7b�#L�T���	L�Bd(��]VJ +.�À���~$���Nn>�ҵ���v;�]NDjҖ��@56>�X��<i˾6M-��[�`�p��H 3q��7��89�\T�Wx�T1ma��R�W�����׹y��r������ǑWg�N����L�}��m=������~n�o�)�:�J-�� .vxF=����J��gHs�.�Q��C3�6\�v8�z7f)A�s��]�β���;��c���[���N3�]�j�;�f�Y�1���NS��e�����n�'F�髎e.Ƴ�z�qȊ v�u�3a������:�2n��j�ɶ���0 g08k��K��m�������;p|�7<i�R��K�ã�5΁�H�Z�+;�صӓhg���]s��M�i�\��kgmw���|kU�s5V��s���
,:���LP	�nw]��Vs60���\�,X$�/hM�Ӊ�ĉ���`oz��*�j{z$Ef��wL ��wb�'۸���m�=K+���&{�1`��A2&���H%�s�,�
S[�Ӹ�Q̶��;~��Y��J���:$�� D�M�n���4������f  ��M徼|�+؞�H:n�(��	L�d(�]K�I7��VS���dR	�\
��W�I����&^5KB!�P�8��$�@syΓ$KX�.��Zzw�t�:ڱԞ��:_����_��0$�!M��В'-�X�	���]�(!�����Y���	#����"�T�b$�@�J%!C7+��ǁ������n�g
����;�[u�tqou_WmH%���J��9��uF�2�1�t��]v{���x��y��Jo(��Q�Et�^4�	ٺ��O^s� �[��A*��\�eو�\=��Q���T���ꦓ:���6��	1��bN�<̩���ך�����]��gF,"DHF�+�Y哔ef���$���]��Af{,�֨�h���W�v	��N%"&"Q�1n�7��	 �Ȉ�'Q�<��{{�,�Y�ʗ17}W�l8
#л�\����n�=P��>�q�A���ʢ^K���e&���	޳u92ܐI���*i�ʾ�  g��o~m���'�*�z'�c�]��,Sw~Ж��3NiO>J����3���9��Y�/m��$�Y�ʐA�F��C7+u2hEH��eD(��뮻$�� �'V�Qj.���RݹHV��s%�B�P�Fq�Z�X��b�����^e�O7�G���gs8u�,>�Y)�HF�S�rݩ��X�����}}|�X$g���s��B�)#
EX7�z����d]b���g�:�I �R�(I��뙥;wH2N�.���$��LX"`�Q!F�s�y�텗s(�b� m�u߈'������"/c{Tގ;^��{H�Z�+��iƑ걍�^��d�N�|��l���p��μ:$��9�S\F��7�i뜼� W}�cj^H}�r��\s}$����$����㖝�$�%�
E3�b�ͻQ�o#kr-��<=ݷX	$�V�x����~$��Gd��Wp'�s����%0%SvY�دr��� �"�(�34�u�$�;;R;��W�"*������Nve���HϠs����A�Y��$�_f��>$fg;�8�O#t�<&���Oh�޹�ZF�o^��T]�˰����{7��\�a�yG��Ѐ��d����w�ש,���BH��ɕ!H���"��=����oU��D�82R���
�wp(v>�g39ՙ�Eg�N��`�ED�aI�y�&�7#>�U���λvMg�0]�Dm�ٻ�y���g/��0T(�@�2n]	$�����#39ՙ\4evf�s�fmǫw9ݒV��:�An�l�̀%�{{��N�"c�I'���;��fg;�O���:��ST��L�H���2(��N�s��'��"z\-��q뷝���K��jiߴ-$��G\������e���рܼ��$<��,��[G����Ʋt����bĈ����b%��vݻ�I�մ%�,��u];)H$
ʺ��]�;�A �u�5�B��P$�	'� �@�I$��$�	&@�$��	!I��IO���$��	!I��$�	'� IO��$ I?�	!I�	!I`IN IO�H@��$�	'��$ I?�	!I�@�$��H@�t	!I���e5�����>3E�!�?���}����"���( Z(�  Ph  (  �    �  h� �     h  �� ���@P"�R��Ј
"�D��l�@R�Q@ (*�@�AE(�
���	 U�*s�    �        P  ��                     �    (VzA}yr�bT���X���Nէ6�R��jUI�����U�m[��R�l��B�� jB��
N��K�G�� w� ����iDͻcf�}� q���=��ͪ][V�3�!6�j�'N �I&Z�3R�;\�6�͕WK���rEW@ D��{�  �� ��   hz���S�%]i+�hr�ҥ��m{j�� ����B��k
;5.Z��mr�)U ����� ����@��  ���t�޳Ҕ /  :R��X<�: N�<@y�����=� �O^ �  �`�`�`y�^` 9���z $�P�  �      @z �X>����7��0�à�=���4� ;:��!J��z�y�ua�y�sU�n �֜��W3���
��  �z|���ΨRw �������U��6�^�=� �� ��
�j�(reر�9�:�ݪ�%*��-��  �  �  h  ױ������̓�*��g��W�� �uNm���i���F�+�I��ުz7Y�Me������m�C�  :��בs��\p ;�ƛs��SW3N-��Ól���u� �C���ځsh��v���:*�("�D��  x 4       3�+[��-�n�d��tʹ5�1� o����98\�+��ͪ)�3�T�k-� �J%��%V�:�
%@|  {�����MnwT��uЕríU)s w+\�Ru�rҩQ� �Lθ��rԮ�'MJ��]e*�� @   jz%%R��  4   )��J�!�` L� '�R�d�P44  �   ��E4�% #&�d�!��&RT�T�&�2hѦ##@��@*I��`��%=�~�4ho%=���_O����>���or@/�5�����ky�C�����@�@���t��p�~� $����Pb��$}�T������t��@��A�����_����6��0C؀�0$�@$�)4�K��	��J���	[ @���^$���k�}���ВI ����Fƛa_�(2�ţ�
�תG�G�&�����W���r�w��c\���!v�x,�[�a��� &��\���o���#��Y�4j�'�,9��zl���n�+%��q(cx/H�Ա�o&g�UԼF];�kR44SZ۹(GY
�Ͱ�Q�Xv�,Մ`׻:2��I�`̕2r�m����+���+q���e��Vm�S�sb��i�w1�����9������i�[FH.m�Z�~��aЅfc�K[;�^�J� SU w`�b:0eҸ�6<�A�X�Z�e�#�/B�kJ�F�ٙ����j"4C��i!1ط.^�R�t�U�"��i?�g���b(`G0]��$�S+i:�@{�+���f�-��6]�Om3V�:ui/Ɇ��NúJ^�#P٭�i%#��r���6mI�Y,�ikR�\Y-w(�j���-i�M��0��yD�N;6cz��ݙg37NQ5b��qӵ�[x&�e���V'[*kƝ[����B�f!hr�*��T;�]�{2�7�b�R(eH���X^�:i^��R�Z�-�aLrLU�jLj�еY�Wm�1\ ձ��G4�͠��l�y��R�ݻ7J�ӣ	Yo4��i���z��䡶�F�s]��\�J���V���@�t�#M	�X�k"1-���k^�*^QW��B����zr�8n�Ø�!Ȫ�C^شȤkoC��4n�[z�*7��aX%�r)SK�E��)�^�����n]���ӳ�G5Vc�[���Or�k]��ZNn�ȭSw����Aeh��n��`:�X��3v�ӭ+�i(Sb���Nj���xm=�S:f8C;O*B���A���l�۰��%���NR֬�-44�f���6�z�Vi�m�/+,k*�7p,���24!����MH�F��ڎ�^�`�I��7K*�	��hņ�۴"˙L\�;���wpNm�&'1Ǽ�+)e\j ���x#4�2�3f��d�ź�WL;�eRmtr�ɕ���[�b�t�R�sd3���1��j5�7BRB��82�*�9i+V��2�^�!����8��hV5�_<ڵ�<�եz��"U�"��mH4[�~j���L���+���vEur�?��������m܉,�k,��-�Ħ��ôf�aX�#�ͱw4�Äb�����-1��N5��n�I&��>͗��=7$��j��R�����/ :ӗ��Ø6�Ù�j�z6��z5.�B=����VV�I�NU�X���],�*K�T��j�zX��*�f��Z���6Ӛ��6�+�z�L��˭�gv���~zE�v0M�H*ڇj������{.����zN���wM�Ţ��)�j�(+4ާj��Z�����3 �i��x�Xi���cfk�FT�T�
W�'����,ˤ�rƊm�*�����۸�X5XCw6�D��h��36���ٶZ8�B8fT'���vi]���6iuY��0I�%r t���p��El#�*�VD�NV ��'N T�M|E�b�e�x��f�ֽ!C��K7��Ʈ-�otޑy��P䩪������4u����5m%�;�h?�޴��7�Qo���<�w �ni�0Tc8�fͶe��se��3]����2��]&�qd��=�3n�1�X	`Mbفl�".vV�w$��u�#r�%�cgl쀳U�H[���a�-f��̳��'	���g w��s6P�rf�`�ڷ�����m#�B]�ƭM:�h
"���xICw��{fiKP�/(�㺩ac�	D	�4��z(�s-=L����Xp�f�9ɥƹ��#��3J5�L���cr�M�w`-c�%����#[u�[��ƹkV�l��g3HmG�Ե���Pa�E���U�Դb*���摢�QF�۫�Y��[ JT��95����Rʱw�nJ���A���=��RJm��{u8���mn�ƻX�ȓ�kv
d���a��wB�0bғ��(�e)$�g Cc�s1n&d�%�w��p|�e��̟�/��ͺ�/(n:͌n��k�İ��Tz�+!.!�.��dP/U�v�AEaf�Y2�	lI0M2���.�,�	�lЗn��Z���D'���#L	�i�z[�͠r�w�6֜j�[KN�q��f���Ai�F�>hͺ�8Q�tŋՖ��ge���Tz�U@�4t���h2�01��g(l�*:�4��fQE�F_�`�՝�S4+Jo�C$��O�wt�8mJ��X�M��@:9j��E4��iZmio ���{�J�[�(�ƹ-���[���������l֨��<hV�U�s0IsH�Fn�N����Tӽyu�A�B�ݰ��dV�u2f�� у�7M�M�B�^�Z��5zQ�l-Yn���WYW��!Z1�7�w{d+�)�%�2v�UwH�û�"C�O+w'�(�O6)�Rj0&E��)�y�b�{n�K�{�b1o&#�U`�	�M�h�i\��&���qZ]Vm����l�X��*�dy��J�fл�)�3��؈c���f������wSr���������a`)�ѣ�*��$fɻYRN@,�[�f�V�ݒ�R=�%�Q�شE����y3�y�V������r�kZ@�Z΋�2��K�`�m���/,L2�Mߠ!�C��Q��u����u���R��bs�z�݆�������*q��rF�[��o-][Y{z�����f�-������Y4mY��R��9rlH �Ōыٯ^�aa�*�PӴ�j�c啚�,Vh���ɤ2����QUک���;��������J�\�ی A�sX4���
�ەj�ec�$��^薯㛻V�b��c��$e�VF����@�PaJ�G1P����,���f�z轹���)µ�Z���N�'�l`m,OQE󡠝�p���C�Z�.h8]DtZ��N���d�ʟ/yݔ���On����MT�M(]��0eهN�¬��=w�1���^�-��֓�k�WG4�A�4�.�̒�mb��N�j;�-M�÷iA��u�G( �̻�V��׷:�pS�c���Ƣ�>�q�Vi<j*�@��;+�R���$�4nl�m�ڱw�����åN]�T ��S�oj��Ch�ɛ�N"Q��mɸ�wfU꬚�a�Ǚ!d�n�U�F���#v����&I@�/^Vo�[���'*	WCX��3
NngL��9E�Ku��x�L�b�,:�G����P�H�K&���Ӌ0�-��� 7���J������Ii�Ok2K�%��h|���E�U�ݣ��N�L�R������9�HU�
�M"�ң�&�\;�&����ae'���U�Y�z�1���L�aj�f��Z!ٚ��]]	�ӻ�,�ŷk#W3a���n��d4+T��9ih��l����2˦�%��c��'SE���2��OTr�&���f=b5ɢ;1VV�ެ�Eł�[{K�6�
��=��9���M
�V� +S��jE���k5�bG2�&���SJ�4`�;zTyEƈ)��G�����:n�-��(�ܙ.�`2�^^���9o7h;�	ڂfA�[S�(�ܫ-0Nec5��`���Z�Qu-c/Sj�c��)�cX�P�pxlD��&��Hn&�����Ig"e^��^��O,��!X"�t	�zF4��v1c�R� ��S�d"��0�.�R��eY�RĎ�X�Tˢ�8V�@�c%�k�)Y����0���A�]A[�Cڸ\8��:�]�*T��K&��IԤ�l�{�wwe�V�2]�]�a0.�r��&���Z��P�L��&B�D��YB�F�\�d)�R���YaK��+N���/0�آ��L���%�P���x���9[�%�ݙ��0�v�ފ�8ڽC)���`bB!R�a�k�,V�����!����1�QF��;ٷ>m�b���Ѻkn����]��l^KC ����xҁ踂u��nw̇5P�Iܚ�5n�1��hn��J�v�-5�˻�$�Q3-��÷�E��.�>�X����,a`��ҭ��coc{+q2fe�N�_]V��X㸷F4U[j�bݕ��WX��U�f��R���gc��%�V�e�c^�F32�-��r���i�6�0��Pa���Z�c�m���i˔��w��б�n䬹��5�Gbw(��ǂ9���0��١0����z����9�ݡz�fVϙtYջ"���M�2��6�����9M�/t�4e��ee�W�&M��1�W��Z;���Z��cr`U��inŪe:�0���4��8��VV�*f:AT@ Z�9"���].��V��˕b��]vmRhf��+��L��J�4	W
{vE��a�W$x��U�ba���e��5����Y���	�Zx��Z�6͋�Up��!��(��z2����xUv��T��N��S�jL�U��ԕZWӅ�& �uy{ǲ�u���V����t)�If���g6�N�㗂���ּn�Z3볩b�p��r��B�%V�Jà��,��ITѤ�GO-��6�;��Ck6���@�mbZ���	^����*[Y�@�^�`[3I?^�b�٫���z��&�<;Mcv)Cf�:�Uy�H�^=	+��Hցmb�:m�~fĩXc۸�ڠd%�[SL�Ux�ĨEI�F�V��.�U֑1=�/`��cU�,"f��FK.��=�B�!�,�ʎʵ��qfU���$�57\���%�-S"���@r��<�B�ɛf#�w�q�e�j��Kc�U�Jݰtq+��>���v�#�"�@�0��kF��G����kU�j$���5���p�3#�ʽș��Mn�sJ�ݻ���`E���wsiS{Zc9r�j�52�+�k�n\��S�ͦWw���n��B��_ќ�"�)��ƕR����ݴ ���Z͘�B�:2f��F�6�죇K�Z&�vN���j���ꈺ�V�`	�w�����e��kkpi��/.�h7��l3[�ES56��'cyM�u�a0����`�W�h�U�`
[D������̊Y�r]h��7ijc7v��i��i�Xŵ� �˭�ZJ�q޹6����YYB��+KzDI��7`��l���).��ڃ��Q6�T��M��r=G.-z�oFʔ0����9G+�5����2T�WjT�6 �06*0G����Ocݭ�vh"�+�P$�݆�e,�wCVTw����:��
Ĩ�z����i+&�;�K�h;e֕Yn�e���56���۬�{��)�[:n�������ɺ�e�"�ҤI�{��R/�y�V��Ȳ��*^h�1RW++i�.��0T�}�aAee7�ZFe���%�Xmҭ؂�n�C
�^Fi����0�{k��

�%vK���ڟ%�a�E��jн��@bz6��J��)Vص%E��>B0�ڥ&��B%����qvD�{��B�:��5���V�ơ�W& 2k�T]�r˶���$�Y�� �/k>��W�5�s.�'H�wqe�;�*�l-���a6���������H�R����P��-��<�]f�#�V��*yF����t�U�o��5�p-�Y #l&N�q�*�7
2�����a�>-����v��ѲQAH���ƀ6𝔶�b�.�<�����-��i�ަ��BL���8�hpDy���jSol�Y��6�Z�\M�-��R�7yF��)ґ���Afi��+6��j4n<��nܰ�0�^" .��4�c��^���l�g@�k`�� tLN-٪]91[{*K�6�Z޼�L�XU;q�g{z�3ay���a�tB���vn'�ܧ�+E�"��e �s
�Z6��9.�ڊ�V޼���`�Jl����V�f�k4�{RGimOefo,�±J%DQp=u0|ոv�(^��i�4M��1k&�f�uq���slA$��DY�Y!�N�N;ܠ�h�s��6-Ub��J(W�.,������
9V��{�qø���Z�-|-T�9
6��D�D�U��kj$]��I
�8>bܘmj�9�%M�U��gł��R&�&���P�&�!�3t�*լT���e�p;��հ�I
+Ƕ%{`��Ħ��)�.Fѵ� �F��^+��v4�zmf��)E�%N�7n�h�uInaO6�^� m�v�V۱ِT�-&K/�R��W��-Y���-Խ�M%���u�D��M�56����5�En`�X�0��uh��V�M��R��d5�!M7��4�z��/[���B���%.]:U��9H�V��L�l뤯,���l��bB�췑�f�l����x���v��sT��t� ���60Yĵ@ 6�u���U�n�hfn[j�V�^��܃2��m����](��խ���D��U��Gf�yu�i,��^���xe�:���nk¢ҡ�s!���k6��n��ʵ��˭�����iT��t���zi���7^�Ν���ҦE�(�{/2֍�Pì[�r��op<n�n���m+��̴��U�w�`o3\S�XP�붛QN�c(ٓ$A4�Bj(���M"cw;)�̫Օ�7�˷��.�Q9kZ���
ܽ� �va�%��N���B�Q�tM�M6���ա�x[��Vt#�1TB��ȕQ"�A�5�H�J$���/!%j�
�,�X��&��3��K3�ü< ������ȿW���jB��}�>g��U5�韧ә�wn|��I%��I&�$�IP �?��I�6�b@�v�ˌl�0��˱��v]�����pe�ě`�e�2� l��'c����0�˰e6�M�N��Sm� ��4�Sl����C ������m�$�0)�2�I�86�� e��66N���8�'`�m��1�c.��.C)��cBp�0v�C.� ��(�\�.Ć� aq��v��Lm��l)����l�m��M����0�N�8�2�S0`�6�˶ �Ɛ�i�.6P��6�P#@�DbI�����~>>����� 	&��U�@I_Y~3��r3� �@_y�F����{�����6��38c��ɼ��a�[�0�o!���Pw���޾� �SN*��R�m��&��c^�$R�bQiAfG`���MB��K\�����}Kz��j�Iv�j�h�ID���f̘֩Ou�Иt�*�d�N�֪�T�V���u)�Ӆ��$��k.��A�Us�1�ԓy]��C,�����|dT�A�fd}ܜ˃�oK���R��e�;k�_V�
�;o���)�U�v�N��+N3��{%�YH�kCvs� �t�
��@��t��w$S[;�����Sp0`XfZv1ځ'^���UFee��k, �өC��c	%��z�]�Ј�y[4<�̐�O+4�c���4f��-��i˒d%�	�0f��&���f��:��W)�&�����.�{�8S]��lC��dO�c.nf��(ͻ�e�xeK��U^jt��u̧b�n�q���B���=������9&N{N��5Je �jHL֪k����f���o�O�S)]^^��h��wtK�{�1��3/7����̀��X;{2�'s���dRG���n�W-�Fr��f䳘�Z��5�XL�V �G2�@���Sm��+J�ɢ�{yu��vM'XH�zI7��Бk�G��Y�̚�Ƨ&p.���Hˮ!V��Yݷ@t�NCh�
HC���m�M�='I��:��-��u�PfdV�7u3�Q�*���[��ۨD�w�7���NYZݮ�b��aX335���JQ����X��lk(PF�r�8�٫ѣ�k�EM��be�s3F�C;M2�QZ�)��Lwqop��;[|�h�2��P�7t��c6��N��W7�oL�3Fh�xi �C�x�j��F�o,0�ڣ��	l���^hUa�S��ͱ˺��ٵ�ۜ��k�跤��Y�E���k��L�/o���oh�m��bT�N��pʦ�+;8�k=OR�Z��/"��eM�x�(f��-�ܿ<��ۭ�xd(l9��=g%(�-�cu)j�г��f��j9\�Y7b]�y�=T�iC�ɦ�
��Yami�)=6���#e*n��a�wlZ��"f3���Ш�3s3I��J#���k�F����!�6�i4��"
��
`Jv�]i��k:�<��pG*O�kyn*u��'��Iѓ`e�i#���u�����u�n]:���1p�-oChI��n��8Z챳Q&��r���<��Xӧ��;n����5-R�&]����r�M9�(�B�K�laڣ7Nf��@������%򡢡��/s�[�,٥�tgQ�"u[W!�[�%�;*�+qj�vL��o{��� ?;�l���;�Y�,[�"i��;�h������Q���5�or�fm���!��5�YR��S����rQkj�&��^��}Ch���=g%���؋u2���o���j�O���2*+3!y`��T85M�kB���tI��z�K'_��ܨ,��]g90�����9t.Y�F��$q]X�!I��rvw�j�^ا�-�]��&����;(��b�S�38��f��|���:�Fs��T-ʌ�����&��&7+B�ځW�I֧5�y�!f�<0��	�����;I,!]�@����$V��X�qZ:���V��t��CAX�;HV�ս��fùb���T����<I\��<��&]�2���u�N�e�՟M�[b�ff���r�ʎ��uѹJ66f|M�Y}/y����Ӣ�Eͷ�ۄS�h`r^&�aU��8�>'j��b���]glU�ԕ��ײ/^ީ���e���І)c��Qz����h��,�&�X�R�TaE$�L��@/��9��uu��[�6��ּ�f�Tb!]�z7�c6�l?ie�*{�&�l��ԉ�ʁQ�v�b�69�LT�H1��D^a4����UE�2����m�Sn�-�9oWk�!�>�`�A��i[�7�'V��M,��8�;r@B���n�(����>�z��)�Wu�S�@)Ѝ�9p�gh������3�����1�U�)�����V����MK��\4NI���G��Ko3���5$���TVe��4�T�-��(�Z~�ؕ�ɇ[�|f@�$כֿ�9g,R�m3D_[�M=�r�[��oPor�1�����R�}0����pD�[��Em�lfa�Z�FE�,�hB�̽�3�Гp2lh�s�J�j���;;�4��[�k��)oy]N�A�ț����*�u�*�X�*od�.Ef��.�o���0B��&c�AD$R�c^TKs��zP�ۛ�"�ZT��W�R�ܑF�PV�$lL�v&VS��P�fePQ6�i-nU8r���MK�r�WFw���r�u���b%��ݞ�\���_&�wWbм����"�u�u�����V}6�i��.���06�q�u�6:FK�0�Y����rM�5��z��Χ�\���Kz���ʍ�la컆�P�#�o���0�;9[QW"�)��d��A��x ���,ۡ��b��N��g۴ss��3��S�O�:663�-d�:�u>u���ڢo� ���7��Tr[�瑷S/�~��x�|٩�[b��VnublnU�3.��k�A��؂K�*M�����fݽ��M%��m����-E�p�]l��mgv�-�������z�v�.̔vA}��a��3��w�[�륃>�>�r��ꌒf��Ls�.U�5�l[�ΰ`�*�m]-؝�F���Rt[Z�%�b�n;�H����ˊ��$[�S�KWQM|�Ŭ- ���h$��f-��4���IMh�d�ws�&� kr6�6�����usI3�D�N��T�Kɪʰ�S��@�*�M��C�W-�x!j��3q7Y(����xWw6 ����JuޗR�f5N��w]��V��}��V!�.��\��Ux��A�ej��ii�RRZV*��b���q�b�f��R�՗�sx��xs6�Q����nر-��k�E\mj؋i���P���:�n9���\�Q�Oӡ[\
mT��'o<ҼCe��t�����V�2�b Q��;ٳ�l{�Ƴ%}0]�ڲ��1l���LǶ�|6uq�KvQ�s'����	�u��[J.�^����@ ��N�����i��s�)W;Wjʵw����_ވ�*z1�m��eX�3��!N,N�cor��:�`��n>���{0���{�]�.�t]�.׷���1�o��\�Y8,[3�as�1�vZ��>�޾kWv��n�V�`A4V#���;�t�ǜwv�;w|�d��5DOpP�/��֋�4����pVM�+b���oʅ��Tz"��6�j�
a3T�cUn�F����bu�;b���k�����w:[�����!�k�p������D���D%�&˻ύ"�ؤ��L���]@۰9V�E�B�{v]8%��f���F�#x�λq�J7Fⵘ�}��kO�f�2�7JU��![N�昄Æ"v]��q]v>�l����Vq��8�ɖ���&�*�/D�ǎC�0����Q9������.ŧ�w��%㨠�*�dD��؇�⤢(�n�l<�Օ������V�RS�e���q#΂��G\�;�����lg��p��X��twٝX��f=�Y� �6������h�NեnӪ!�1i5�j��+�Doi3�T9�qPbm]h��؎�3�����c'�f"�csxb�R���ɺ&fEa�������u�,�!�Aj�_fIN���9q�r}��7r�e^E�Lǹ����53^�U�hµ}v�BD���ݬ6Q�n�l�|���rf[�X�K�C	A@��	ZN�յ�]������VY��Y�jVm{P��kf�C�n
�We�ˤ����z�;L}���W���XB����m'W	Ro�L�b�4�Ѷی�4���/����`z�����yc)���y-�Ҧ��U�\��5���X��ۗZ����4<�W[{�
�Y�&�)��e�ͼ#��5��h��T{qS�+�@��Y�l7Vm�X�ӛSQ*h���%�v�|���9�%�\��*��F)���pȵ�2��A�!n�����W]ytL�3ow��vv�I�=����z���N^W^aDu�6�(�jؑ�9O�!+.�u�:��M�]/���J��"��e�s�p��,�ȍ�;����e��;�f������p��&�R�-�2�M��b4�*�R�#1D�)m�\Nغ,������'TFKs'D��t]a�ڱGq���́-4��_��;(�Y��C/��ۣ�Yd��)��}/+�swE_+�eX�y���2�\��s�"�:=e}�eL
�r�*�E�WA��ޒ<6/�'u�a�0����b��"Dn��X�&VJ�	`S��o�l��bϛ�EoPA�۩�8s���;,W+W�5]	��*q���������;��iѦ�tK@���y�73jVnQ����Y��ˮ�NE�8^]Ӧ����~��͕�Q1nk�:e����][�rؼYx:?����Ԗ�D��Y��R�V\���(8�lսzE�<Q,���$��ge��D���`e�x�;7wn�u&s���+	�7!��f�m�[}Sb��aܠ��09�Y�wK���l�n^n棻/���К15��M�@�(!
���j����S>�l��ba$�:�t�x9G/;�����˝�q���3�.JAr]g:�CP��֐�yiaC�ǡ��W��Z�Y}�zh[�c�N�Ӱ��?=V�*�Q��a�y�d�-��ccP�6��
0�S���G,��]X�kKDE�ؘV�n���y�O�r*�5ɗ��%'PQlm����y]r�Q�u|H��`G�=��;�ؙL#)d��3g,���by�ir�U��,B��	�W����Ax�u�j�]��0�n��4f��pñ�ŭ�Xv#�n��tZ�h�2���E�b�Bt�eIȣ��P�2o�����[`��{'���Ů���Ы�U���������/ 5sA	��L=�0ԝ�v���f��-k̊ONzF�S��R�Έ�ك�0�73O[�W�˗����J��}�@̾o1�Yp@�i8ۗG,M�l�Ș��j�[X!l�L�t�Nm���!^,!���yn���ՙzz�a���U��}N�������.�+�0�9S;|��VP�A�
�׽?�>m��h�w;U)�>�[#*��[����+}]KD�X9@���EoA��֞d	������.����Κ�8�"���C!�mn=	E�8�$��ul�Y�{3�ʇ�{Hp��T��t!�n���)IHC���oa�J��p!����[���7�q6N�w�-˭{���y�%�f��ZJ��j+t0�Է�EՕ�o6E0�22rNj�P���-p�!4��]N����F��U�:v^a��ɷ�u�զ��Wh��WmSq�=�K;�{�[۽�_Ɋ�����g\�̦M+�G�/��-ԫV�#N-��%���'��9��&tb�n�\U�E>�iuv
��+:�
UR�*�MK�������M;��eTz�Y2ȍ�SS^�m�n�[r1`]CJ����w�uIy��Slڼn-2�ѭ�Y�Gx�u��l���pn���]}wC��u�Б��×�ũΞ�b��k�PP�/��d�"�����y��T��4{7��a�Y���g"�
�yy:˴�ȴ.IH�ʄ�,�"�&m+�f��-����[�����v�V,�AwJ�4���� �]��"cѥ׭�>���L4s�*W>��iK�k5s9��d��#�%���j!�(�{*\�d�6�-ɉ�M[�aF�u���v�"�ݬ�N־�݆���/,D]�v��j�r���ٶ��;�97hg�hד�v�}1]���F C�2��nꆦY��ͼeJ`P�^N����ׯ�����.�uc�Uս�c���֗�4��� �������V6��2R�T4¸�u�奔�̋f�m���u�;B��t��7m0��d��t9�wi�G;�yC;O!����9��\V3�t���ֺ��{��B�:�c.r��vq�5�NKCC���M��v�U����9׉�	����$T�RV�s.V$�j^lFn��nt�qPC� ��s7S�Pb��{�TZ���w^l���ؾx�˷���./4V`�}���]w�7+C��:�(̓)�f�E!�T7h����V\�:!+yWN;)t٦�+7�m�)��sQֶ�͌��������mi�;X�'J����z�*�%pY/%��jO��2N�哪�-���#�Z
�+<�ݖ�]�b{�Ii���c�Nͷ]��7r"
J&��p�RĔqkx���"e7v y��6�N���n,;ee0F]ʛV�DUm,4�HJ��Ҍ�̌;�됽�d��ΛSX}�����Ȓ�V����r܋�+Y�p�����i�lqO2Ş�]�Vd��M,�wS��l7�һ%�W��9��[�����.�'��v̛ڵ�ߍ+z����
�n�x�����*X�\P�s��F��X�l��$�;����.���fu�Yvj��4]�����l��,��T�3�+��¯ȯ#9��TQ�I5f�*L��De�ud�⸴[j�Fn&�=2��T�)�G}%���^�cUx�.[��K�nL�Փ-���1e)&u#)1Vk-0U�3B0^��r����������v�͛�R��9Cuk�Eh�EW��_K;����*��?$$�$��ؿ�2$��'�(hyq*B6RP;�����UUUUUUUUUUUUUU*�UUUUUUUUUUUUUUUUUUUUUUUUUUUUU*�UUUUUUUUUUUUUUUUUUUUUUUUUUUUU*�UUUUUUUUUUUUU\M��A��Z6�i�]���g�v(���5�Tܱʃ�l��p�\/<���Ĝ��;t[<��������t��4��md2�۫u����1�ݗH�g�]��f�f�I�t�bS��;ntbWp�:�;��BSh�`��d��ö�e���Iڶyp�f2��w]8L��D��`�ᣥ�6�1,��;�]z587�l�������/,=���o=E�kj��nx�,�Ż���m�z�l�*]]m�W���cm�z��m6�F[˵s�6�u�.;L�3���9��U�v��$�u��#��wjut6�.9�<�J�&��v�Į��j��K0�f=왅�^Wv��ܥ�ֻ]�pמ�6�v_'\�{u��vƷ��e��7���A���\�R�ٸx�zu�:��ζj�xE{s�U��jֻTg�ܘ؎#q^�kʐ���V�ל2���<����xN1&s�1����r�K�ϝ��]Ѹ��.+vA2]nrt=��"g�b�b�u�9�cRɼU�V2{&=�mn�&�#�.���3��6����\C��1'�p�ww�<��ʄG�%�!����o=�Y��C �n2���v�t�Mk<�C;Gv���8��/n��;<�l:h��o)�����}�n���EK��X�.Մ#�ݮ�2VtX�(���ݺ}Ed=��=�D{8q��c��QwZ|�f�n9�s��Rn�.����ӌeۮ�l<�òN������2��=;8l�zd����0�f���[Te�wAX�ݹ�rrJ�y�>�7:�	6٣u��w#�1�ᢚ�Z�g8��Y��]dLg����)�7��;�ٸ��z�A��e�S��Lu�U�����=�]�s�Y���U��B�]�
�s����+��ơn�<��k���Mq<u����l���qJ�����X����箒^�FkF���c6�mO=n�N:h�b[n�q��rKQ[��ӽ5�^.���7f��ӡ�g��qͺ�P����Hd�����<��4v<o/m��7cIJ����,�N��s�DucI"<Ep[�:���Zժ���;ۡ���-ն�d�F6
@�^����4�=�mK�uyP%�`	�C��˸���Ѯڹ�z�;���w���yt��"�!؜��d뭇����zx�^H��:�svn:�oe�� ���d�wO��ӵb3�7f:܋l�K�<vu�6���k�6�5۶��L���^\��b6�K�)v�01�]!��.�=��]h�$t으vv�(�cq����#�kb9�ls�AZ9��b�*��
�p���B�g������k�� 78{!�G[���.�r�y�o:�����h��ܛdr�gw(�jn�N�w�G�j{uλg�����5�a�&y"�q����Ὠ�O�����4�&���W���ۉ�h�3ɗo:��+�<�q����:�/G�@qz{+�������.N�vP���[��m��\rqc\�i�r�.3*w;���IMŎ-���g<�z�a7n�@�Hz�mr�o9f��o=����Oٺ��ܖ9��v�۳�G�;ZNM<����:��8���[v��,���nل�#����=�ٸ���"k�9W����<\�z�qu�s�3��v�ۍ��P��=��	>9Mpհ�K:���V1�Ӑ���f'`:��c����u�5�n�;6�ޅ�"�ۇ��X{n��i��\�/��&�z�3ۄKPO7-Ōs̛��ݣ��K˹�ճl��������6h�olB�c�o#��+�.b{��N���f�8��V���n��oq�i�{I�#�Op�U��'��0��9���z�	��7��9��z��ݱ�cz���g[�^/Y�|v��q���Чa=����Q�õ�{v}�L׬
����u����@c(��O&�NB�c����M�틢l�:�0v�a��M�\q�ɢ\t�n�A'(��L��yN�����Q��kv-�'2��z�����T�0�.`C�x:{�\D��l]�燹�q��@q�ع�p^�Қ�&9#*ᢶ�͆���m�g��H�7n-Q��:Gq��q�q���Y�mY���m�b0d�n��7�I�s��ٰn��p� #k��;��qq�O'f}��n�kn����m2Z���p�חm�q�l��V��{Wk9k<���Ow�ZN�*���<+�;te���������m�A��x���N2u�d��뗎��v��FBZ��+Q�v��ε��������S��d	�YX��I��̷$u��W���^�¹{c�ر㝋�Ɨd,ѻvle��v�/�ϋc�=�i`{h�b��cn�4	&��r!3�d�:��W&�6/R>ܣ�v�Ѓk�U�j�uxE���'�=`gs��G�����w8j�M�9y����&8SWp� I�0i���@�k����Sh���,r��+.:�[�}2	&_b��7,۳�^am�E\D�Y����ӶpE���V伽�n{Yݞ�=�8wX݇@<T�j��{"�q�r/Lδ��pu{ ��b٤��1�3ěg��O.�v�(�8�8�Wcv��KY��t��u�WI�nlu��v��m�;w��W��w��E��3�du���:'m�l����f��yZ[m��B1�'�Wr��N�,0����cOE�h�r�e�ݹpʚ�;)�\y�E�����q�0k��˫q���oYE��F|����N}`�n����;y�����]]�7i�K1s�/i6z�y���s���ce��^\=t�f�-��B�6]X�Յ�ykG(>�8�6M@�Ȣ�����ut-r{
��U���>�u�q��u���Lm\;��qcq�ڭ<Cq͜vn����b
�v�����
���c��{��=\�n��x.�����zzl�@[���OGŚv˜���Kl>�y��s��h>����U��e!�{Ic��n)��I�N��n�z^�pV���qO.���\�/#�s�onW�nۡs�3r�<d9��+��w�`c9��9\(.랇�ɺ�۩+0�qu���iڈ��>�:�[����
b�U�k��nncq�M>�e.]�"�Ëv|��O�E�8�����64u3�g���AmL�Ǖ�9ȥҽ�r����^���li湷a#����)��ٞs@�8��; �r�ɷkN;G���i:���K������k��5�Nl<Վ3��i�u�g�Ӭ��ӳ8ݭ�-AnYe���8vjy�ĝS>kc�%��p�=��!=�\�;v�K�d8yK�`���kp=�u�� �����5C��<�Grn���[h�W"b��[ڶ�pn��3�*���bՄ����m\q��#�W:�b�G��u۷�(F�b��ҙݱ��/��n�n2{�H)�*��y!l:�鰹hH�2���T%��2��]�s���{�q��l�mz^�8��&0�O[��ۍFq��5`�uOG0%�N�qm���ol�]
�8���d����.�(��d:�1�8�ɬ1npkH�f�^]��mu-cl-Ɠ�����uSj�j�2&]�zϱ��'�<-�N��{O�8�۲y0Qsǅ2�Ɂ��q�*�m켝W5�h��]��lM��9�Fnm��W@�j�q�(k����'nŁ몠�F�E��&z��3�ն�1�f�l^	��p=h��uM�6��ڻ�)��k�s��2�Wb�+ۭ'`�t\�`8��͍@\6u�;�0v�c���Pp�x����õ�˔C t1���BO<m��xWg͋D�	�6<�(�۵B�Z�v�:��Z�9N3�#���.;/�5'n;v�[;��d�';��^^yMz64F�ϲغ���\����"p]M*���<W��׵c����<=v-�riI+Z]��R6�i�lZƹ�sjKc��X�v�w;ѵμ�z ;q�=im�$hݖ�ocm����2l72�<�"Tr^����*ˮ�$Q�6��鋞�h�;a��j�W��΁�� n*z֫�,��m=��;=B����&�"1c�vn�m�M�h^7���@�۶кp�n���am�9���c���%�\���B��"`ŵ�G��\���;E���hw[Xla�`}/s�<V�n@*�7�g��=��cۛh�I܉n������xv۲��&�az�d^f�P�C�î0��Uڂ��x�=�δ�;s�˩��'u�m]����8�FW�ت(�pg�&X��ֻD+������d��l\\�Gcvu�lX�:���J���3g�s�x�.Ȗ�v��b-�=n pd�nG�5GH�V��p�w]F�u���<�p���;X���7	�hq��L]�qg�k��e�z�:ކ�'\]mgh�S�u��;\n֞�5����Wlf���ۘz�l�s���=�W�<� rNe�Y�z��c�q</�ԧ<��m'eW��{r�ƻ+G��k���������;L��ݞn-�rk�[�Zd�}t����y�;�-��P-Δ.y����s����7U�3m�6^VYu�9�l�󕷫�:�M�m�v��̆�s��ڝͩ���v\Rsq%jnJ�����P)�\�A��9v��u2�(]E����rq�2t�n�zq���^#�ݸ[���"��v'o@�j��t�δn�TaNà�[��ce��!9����8�:�!�<Sj�V��`�9��q����\/Q��%�mv6��<9�\�^sb"�ˉsmkf���c7'j��=6꘽u�v�zh�\q n�g�.ۜ㋫=�n��KUT�UUUUUUUUUUUUUU_�߬��ߣ���aL,���r *젢�M:dnW\���3��C��Ap�ͅD���TU0��Y2��N<�:!v��d.�'qu��;H"��/�i9Ur�&�W~)�"�:�BN�8��y$QL��qy��5���Ruѡ����hs�EW9p�#��\*�.�Q�$QEQW�;��ZE9���%˖��'<�:����	�P(�VAqT��N��Q�G�7�$��U�?h| �9�9�ePU�/<���	!��S)Ԧ\��xU%&��v��e���̙AU	�0
�P��;)�Qy�T�I�2������aL�Le �PE˲�r��*�(������ +��Iۨz�P.&wtnEI	�Siˌ�)!:BUvQBeAES.�ga�вﾑL���;z�i4��x=���ww�Ϳ������U*�UUUU*�UUUU*�U3s]���.=���q[�t�sV�uc���{���68�\
�77f��n��ht������%�����ӷ.=�Wdq<�W4v65v�-Ѱۘ�<�)ϥḍǝ���1��L��4�B��Ҷ�GP�Ԝ�s��H�p�F-�N=��{r�ۃ��*W�av�on�n��OJ�;��&u���״w���Z%�8�ںv���t����^j�pn�{"t� '>�&Q�T��Ʈ�{�h���gz�n�<=�<�fv�8lzNmۃ�z7]K����*�9�;�EKp]c��*gms6�C�i�
&�6cn)㎺;n��:��]sM��#��9����{2�i��.^h;FׇW���y��mǶ��2V��'l�1�]s=Q���7chz��cfk�<��síȘ��\���������7�D�,\m���ٔxN9읹��v��.�/;w��4���s���j��\T��%/�o`8�+5Ɯ��������v1�nRn�F�\�ݩ�w\�����n�Y�9�콞p�ɵ�x9ۛ[^�ɔ�,�ܾ$^��y���/�=�}O<���n����pA@�$	mm"'U%�F�@�Jiu؄w	���ob|�Ykms�#6̇�7��Y��n6:iz	��&%s:�b�"O�q�X��{��������q��ۓr1D<5a�mC�-��.S���\���!s`\mۘ�
���OW磜j��;pu��:��D�s=��]���&ܷϙ>w�#�;���t\�m\��L�[<�Z��V�l���XlV�86��ы��ֶˇn�z5�s��Ilus n�����ہ�n��`�j�^��l��c�n�e��s�㝍^m���q�N:Ɍ]bܼ�m9�9�f{Y��o\���f�iI.�+�OR��/Eڔɢ��Z��[�n�\J�U~�����~|UUvw��ø�0�<���;n���
sɎ��{����캦�Ύ{����tWQ��$<[��眹y�x|��6�vx���!�$�s\K�r���rwe��{r\�B����`i��N�w<=�j�b�!�:�jn;��軞뛸��F.8��vrr��<e�Wq�;nJ��C�[�W���{�'���������ʿ�/�DJ��VS>_�}y�f���������zJ�_�t�O���c�F$��{��Qi5N��r�M`>kֶ��;�jk��|�}���m����  ��6ز t�P�~{!4k� ����P`y�.�M��� mv���x����'ā�M�� �~�D�}uf�곙`�[������l����h��k��?Q Gو�D�����r���u��/�s]˘5��HWdV��AŵF�	����[�Wuh�(��w0 {9n�@$w|�w�gT]���{���<�Ӓ�ۢ}���m��ڎ,l����j:	���2�;e��w�K��ۏ�t&I4H���@?Q'�����+Yx�eۀ=s=L���ig��;�_����{�����A�J{��~�]��W��I��ju+QQ-�,�L#�N��&Dj�lh����r+x�g]<��ڸ37�w��,白҂���^���$�=�1I��l h�ȼ��s5�j���]!5$~�'-���;�Z�߽���~�M?_]�bA��� �;�w�ǿ��j(&�U�V�=�Ū~����X��~$��I�$�ӷ� �D���]�[���ٸL�+���\��r(��([/���6:�$�箓5b����%��$�M��� ������ �s�0ŵ�R��8���h��T��J��������vn	���C�{i^�P-�ְ�:j����~�\�]�g_�	�*D�&��ok`H�=��b7U�l���$�#Z��Z�Q�R' D�f0�64��m�@{��DD����	?I�=��oάޫ٧O��t����b%��VP���y��=����ˬH�/���0�g��T]�b_Z��>h�I��nr=Z��M��t9�r��:%�"�L��c*�j�"�ݢ�wj�m����%m]��ܡM�M۴�#=�sx��9��İ>̺BjH��N[i����Uٍ�ڵ�w=���> ��|���s���o�zH�aKD���*X��$��]࠙#�9�I$�7q|���-�{3OR���{�ă��.`�{��H*�N>\��bs��cP%U��jc�W�-i}v��i��A�G�S��UV�)Qk��<�#:�l ���R����M7��d�I>٘�'E'�s�7&.�=;d�@ w=�ɞ��]�@��anL���� �օ�y݁Zu���Bh��#y�'�'�M=3$�I����g=���&�6�eڕ�PKn<@��x����=���۴��"��{�I$��@:�MQ3�.�Z��b$��VP�G����\�$޸s���� ~�{>Z� 󛵽z;y�Z��E���xRl^�R�PG^\/#����H	��J����f��LG�mk��(١&�[��D=��9���CK��8d� ���� #��d����nA�Fܶ�1�rפA�����דI
]�:�4c[��I$�n`
�'���B����^��맸�笓q�qy��Rjŗ��Q�:yy:S��qĚ�/[�R�T��}�~V?��=x}��`I n�$Mh���� ��!��Y�Π���M����[�Xy�(te�����R��%Bh��5n����Z�쏩3D�@�nb$�O����僨g�Ӽ�k���]����anL��^�w��BI4N��]��8<�3�Ě$�ˠlG���x���*�Y���[q�;{0����k5BI rX�5D�N��O�4I�����M{t�x�#>$;1PZ���b$��VP�9�s{�����⏽�g�v�38 .v` "��t��D�w�q�6������u\��RY�6Zb�u�؟!��R�L�9���]we-÷{~˱;+Y�[P������Zќ[Ԛն�m�%u',��	���ͯa&���1�EX�vy�;%��G��޻y���x&y�9��nv;�+nt.�6C8ϛq������񺇹.��n�)[vہ�o�������on^���l��m��l<��B�tcj���3�Fݜk�l\�졨�3ʳmN�n 7l�]y �<nk�V�1������k��N� ns�J�Z��S��.�Z�,��'b�'-�h9���42ml<d�j�=p�u�n��s��??;�F�j[i���ܺ������ ;��;[-Wx��+��j�^��D�Go��c���85�c�J��@����O3���+�;Z{�TI���}�>$��M����|ٿk*���kJ1�P��ke�&#Zｽ� @���5���<P[�'�̘�6��D��'���� ��˟`}�L��B��d�& ofpM�.�O�h�I�|��@9���  ��֮�^��7� �}�f��/o���E+n���m�N��2I�@��H��!7jY'���@ �Ozn:d�4L~�D�K�/q���}}��t���=+�NM!���ok%�=�sɷ=���س�����Yw���;%�2���w��  ���� �0��=�x��,�S�HA$��l�������r����[�F�bD�9�+'gݘ��[D�^�cQ]~	gl�Vjӓ0ڂ��w���m�������Shtʈ�Fi���5F����M�����$�$���n�$���ـ ���Gۚ����tV�9�U��+O0���` �3��Q&�����E�7ݺ �;��l���z� ���!C�-��옍w=��7����_v^���7�]x {;n����2�o"h�O���ɩ�~��S�N�nL��ց o��{�Kg�����y��Ck�} %�.g�؃�ً�I#�}�}

����HDĞZH����ck�\`m�8����@x��pqt947eN�����=dR�����ַ�&j�4H���DI��}�B_�3{q����gw1,�H=��A��g]a̻�x��v�!5D�XI���}�r��f��@ �r�  =�{��[ �����5��0���d�x��u~b|[i��>k�Ih A�绛�a�:�t%.'��F�LD�}5�g�<r6KY���i�A�ԩ��B� +�)�+�h� ��yn_�q��!z���&��������D���.�9�U��+O���e={ܱf�s�ā�" ���!'�G��n�{��~S~��i�7����F؅�S��Ey��BI4N��cK|d���W���U�DA����#����I�J���m����v�s�v���ŝu�Q��l�Z�G4zS���R�,W|�<�u8Q����@�LT��o���O��m?�*�
�����m��@ s����]�*�YV�@7����_KO�i���b��'�`�ϳ��w����ɘ1_t��gn�5��ÙwB�%��$��7���+���Hdִ���q �=�w����;=����f]}S����f��F�g��[�8)�&���됐>�� ����]߹�c���{tR��P�7���8�06��D�#G1��H¡�9`��Ŋ�)�}���zM���U�
�f�2��$-�����w{�`�n���UjJ����m:�I l�T��8UgR-ۮ�ABO�svHH��v� �k�d�b'�3_��U�|���|ܩ��몕���Q�_a༷n�|�|Gp��tNC.������ZZ�y���^|��\��}��ۯ�$���N>�&z�!�|���A���۶��ME~�c��d�& y��}�A�o��񜝞��X��&y��D�O�s��$���D�s6��7֒���y�wB}6�YV��-ǈ0��� 7�r�h A�vے�os�^���l;3���> 7�[��wY��Y]��ڊ��u��R�Π��3� �~�%pH���*$�$��t�e�;~�[��� &����3S_G�O������^���s����L�	��h�^�ݶ� �Lj��#�_-ѱ���j�'�иF҉���)���w{)�Yic鹒��)^��2�mK���n�v�9�GA�ͥ��,�<nk+GQy�*����Fo��UU���kV���9X�즍+�����k��{q���OFݻ:,<^��q���e�OE��F����'�c��t�<�3�w�v�0�����7����.ڸ�f�g{ ��bCs]���t[������O]֘���n�	�Ⳁ3��Z�j6���
p��v�XюG;�����j�Wg��qkX;\�\(�j�#p��7.�Z�@��{�Nў^���屘�.�V��@�6<�o\��]%B�[�EC�%i��L���?!���zw�HL�<���y�\�a٭dİm���@,(�'8�yB��l�~�!$�W���c�>���I?Q#�nZ$G�}�Bj��f�>�z��V�Oy��p��[�Fv�� ߹��7���p�;�r{�xü�@�y�f=�8�'�B��f<A�w�}�e�{{�}�|��k.� o���� ����tc|ݪ�cI2��=�S�Y]���5�{����h ��\�Ԥ�&b�e� {��7���93ܘ�������[}��a,�$48���%��rn����AG�M�v-������/s�Q�:8'm�x<{,zo��`I�~�l�}2�]e�[n��>��Z s��o퀭��}UV��<���@AGm�7�w¹Ŧw��?`��qvSv`�'�q[��Kq�yn��_l���ξͱ���r960F5wx���I�.X�yq�Q �w�d��~;o�n�b
�n���x߬�(�(6yR�/>v�)w�HMQ&���^3D��\X:��ES���D�$���l�BN������N�VKu3�3��~i���"��s6� ��߹3>���tuƄ�E3U�Իw�����2ُ�2�m���'Q��0�ֽ��h����Ӝ�A=������tݖJ�U�TX�B6I��e�I��;T��Ͱf�tB%R� �R*FUK_;����E��������6|��1L��X��RD���S���fOl�5D�w{��54���B�N[f�����h����>�۝�� O�;3��H���r�UD�Z����xk@�'���$q��UZ���>Aܞ�L��]<I$�� �M/c�tVn��5�yֽ��Z��5�G��qknp�֚Օ�R�d��;f�k�Y!^�����ǽ��u��-���ŹY��|�l��8ţ�nsw\�g�N:o+2�웮96�r�*�h����-��bՖ0��b�/�厷&�_wgD7�˧�4;�9��%j�΢x0���[P�}�?�|���Le�y#�s���#Av���u��F[$� 0���V���k�T�����N��{9$s�-�l�7CF���r7��=�2�GW��5�n�
�����P�=�M����а�Y����Ы��sr♪v���f���X��4$�v�pPx��+��I�aeM�F		bv�PӉG ���0��L��qW�����8���,l.��X�	ZB�oX�r�'��#W�KX3�����p.ӻ�^��l�)R)#5џ-!Fk���耱&�����)P�`��.�J��̜!�1�	�+A��T���Zi��Ǆ9
pV�%Ԣ�V^�K�!�=,c5�e�=Znff\��J`�w���#�z����0w%�҆L���O3f�0w��)�#0L��m�8D\m�{�Q޻޽���E9r��\���dR�W|�@"Sg,KT�����"���(fXD1��J�Ko����ļ�|�W^��w��e`x'�}��I♍S��e�B��4����S�k6nmnT�QM��:�A�IH��׈���}u��n6�vnf��d�cGV�O�RJ�v��v���:���WLá']<�[�ìm��n�hm����"�ӏ�N��E?Rc�(�"(����!<�]8;���L�ɔV�WW��US��9��IRAD��Q���C.&I$Qr���WMС �s�}��ۙw�r��!u�e�\ɹ�]�i	B.]̜����5��;��L��RWꬓ��L�F!]�iRE����%Z�'e�b��͑@���w	�N���5A�T��AG9�t"�Q3@ҙMU���ι.��!([y�X_��$�_��ӑ]"Y�XqV�U�0,�j �O��p�^�C�<"�(���W4N�OZO�r'�j_wq:�T贄��'i�S�
�F�˴�n��{܇=o'�����(�dJU$�aD���l��옑�w��k�h���  �ε*� ����$zw�\�*(�n����IQ�9^ȏ~k�P�f(�VKw6�Fz��������뷩����I��޶�$nZ$};�6�����-33��4�K���g����r�Ԑ��n�h�1ݵ�q=�r��5%�����?��h	��~�0����?�H
$�t�l��-���4oܿ�9E��׋���Y��f��Z���?ݻ���$sϼZ��|N�p�(���:o��!< )KI�{:�d�j?U
�9m���ܺ��7�﹛K`�:o��������p�@��f��|�����H�aڝ����{�;v�Ke�ہ� һ,*�@>�v�*�$����+�Xq����ml��={GoR�������Q�D�f5s�aa�޵/�p��oU����f�}���]����az"�������4]�e� ��Q?A����/�3�_�������g9�f�ϛa|���x��@�{u?���:��3�6�k���N����!��-q�����1H7��8�ɐ�NzL�v��m��Ym��{�*�:T*K{/�Fr�'�O��{��>$����1p�\��缂��~�b>�ڛ�>�[����D)X�că2w3�E�9�Ws{M׸����4Is}�BMQ'����d_������sd��谁���z������ 7G�zl`	D���h����J��joj;�"#��>{���?%9�3!���NT��kze:;|�N)��w�������l@~��ɘ�@��r��ћ��\BW��]��{�ޒ�1��u�)+OM�?gf����N](o���S���_UQ�'�$��BM~����o o��Gu�]�Σ��?��m�.�x���u:ڎﭭ�xv[�o.�B'l�򁧵��=�jM�+�A�f�t[��n�cu���_@"������Յ�NR�0&k�1���9xw"��vݒ���;YHҡ��{6e���ɞ�(���r^�Jq�v����zp��la���\qWn+�$�\Pa���ѹ=�潩$�0��V�-�����tpvc��oF�۫\�/��#�U��W>k���]sv���dC"�1�G/.ɖ.�<��ۯgvSS�b�w<48h��k�C���F�4�۩y��#4�>:��g��sݮ����S���g��K*�����w�����1\~���Grx�է�������7���ri�ާ�ʫqҡ;3+�"U�j�o����ݼ�
�&��>F�yM~�my�x|�2�վEg���~�}�Wt0�e��g;�� |�����Fw�ܝ�N�2�~@ �Os�0`�yM|��k�5l,#��C3�׼���[�{����� ��g�gyf� y�w�d��^�����{�̦��u9S��m�<|�}����6"�9��D��>��$�$��r�$����J�imzgw�Y���"t��S��QP���&�l�x�z+��S�]��d�n.j�������n��r�=x;��|Ü���s��f�{|6��!V�h��e �{r�%� ��Kj����罽��ަ=d�E\I�^�R��-װ��9���%��o�c��v����9�wmɮ��2�[���<��!I>�˃�?Fƭ�;P�B�Cڹ��W7�U�I��D���I�c��|�}�b#��L���N�,�L�}Tn�۲�� y��K@��=�����y��Z��=��5��D��sĒI�9��k`����Ԋ"�e� ̝�޽�_n�k� o���� ��{����&�l��a��_~'rf �S�$��S��v�������2`��y��{/�=�I%��D�I��B 4wٺP��W����y��Ɇ�fa6h��G�;-��Z���^x�C���z�e��]�]���MP����]�ʘ�����~�]h7��s�	$��7K���
3n��v����G��w{��2E��褭4��\�V�"�&���V�b�I$�w��f� �8i��	�yz'�Ò巟�k�[T��k��ok`�A޽���HeM��ָ@_��ML�[�o�b!��5
�;N�MŜYڭ#&��-��w��2ٝ��SU` ��i�Ow�j��gfuWވ���������ݼ�`-��\���6��C{���y�H�kĒVwsb~ ��͙�`o۶jks�A�l�4�L��HMj߰߁�uxA2�tJẃ9�Wm]��<��u=�D@�Od�I$��f���I3�1Q;莵�M_��l���(���RJ�N�BX�R�P���x�� �F[�ke����1������і�&��z�d�$&�޽�� &zf*�T�y�>���S��A$��l�L�O�y�5D�3US���J����*
s�l�}�1F�I���n�$�g�`
���d��"��~�IXE;�@���RV�`x��5�o�ݯI �����Nv�����=�>���}���v��8H$x
�̫���+�=n��g�j�=�d��ï� 'vf �'��Їa>9J���fѬ��HݓI�ڬtO63J�P��B/�����t��5�Y��,��,�;��!���Q9{�ȅ������;1`p�9Un7jm�fk�*�q">I��xp�q�\�_� )IK�I�{�` #��t���Z;$���E%��۳�66�7i:;<�qxa���Lm�k	ֲʝ��s����+����u�4g2�$��bD�I5���'��s�՗=�g'�i���۵�}��<�	)b��$7G�:F%Q<���pzjW��� 	}�t�@#��y��m�OY�銼ֳ�9���!��r�'-�0=�Z	&����r� �>��3��!��%�:g ���	 ������5F��d}TRV�bA�M�oz.>��� ��]}�@|��{���@#ݼ�o�/{��\}�� �PL]my[j���{Ӥ�D�^�mv��'�'zat�>�M�I4{�� J��ͅ��vD2�q��ҳ&ev���1;��*��!��n�}�K����О)�ܮ��A�4)x]s��u+.��z��OW����ꪪ�"u/7Tvl�����[���췠�Y�t6���\e1˯����l���=ȸM�8��+p(���n5���}lNj�
�j��ql��܆,�Rs�buf���EZ�뗐�Ȩ��kڨٽ�����e�����lW��OLxe���k�9��U<ۜ�7cZ��r�����.Єѓ�7^r�I,�Ћ�Q�5�,�k��Z,�qY/V�&���:떮э[��Wv�ҝ���]S������u�`�g���_�P��{���� 9�͙����{�^{�ɮó9f� �����5ϩu�XleM���L�]6�:�3V���\�C�s��f�@|sכ1`����y��[Q浺s�^٪RIe������d�	�^�l�I�&!���J���O���j�4wٰ��nh�ݩʘ�m�ϐs�,��ξU}9��g���{��3 �~��׺qy+º5D�+۲J���Qvh����'޹��d�Hӻ���^�r��aK���k|��@|{��3|�F�f�5Ƚ_��^8��ܕ�m��7&�b:-�Nx:�n����|��y{i����1k���ہ~m~V��j�5�o�������L0!�媢@Q�\tg���k�������Xl׻,�cv���`<��q�ҟ�ړ�2Wr"磗[����h�#�t�8'�h� r�{���n�*��"��<�o��VJ!�)^��i�ϑ����#�����L?=�o7����>{����ѭl����a�o�E�;
��xgs.6�|�.I�k{�z.��F���@'��-�L� ~���k��e	)b��0��I�Z�v��/�I>+���'�1h�;�Ϣ��=�_�8Y$�}���x��NT�Kl���ց ���{��fMk|�]��d�W:[d��M~ܒlDDos{���Q=P��d�Uxx{�d���&�K/ZV��uix6������ҡM����1N��+O~�߲��	U�DDDF�7�K��lt���2Wtϰg�$vs�7�+�]��;~��y�� k���ɕ~��\_y�0	&���,�"v��Q9����훷���z�bcr���b3�J����}	��O�3����+��ʼe��M�]��[aD<cOV��!�7v쌰xf�.vQ��fiΥ�n�e�
��_���*��8�[xU^~���'�75�I�B��I$���l,�LH�&�[Y���w!'|�7�ң�m��'�I>�{��I$i�m޻ͼ�I6�A=�t�k\|ʥp�]�Py��l�D�x���	�'�L�4u�S��N��&�7��A��v��m��<���y�<���6�GKA7/q�zݲz׀��;���G/O�����~�}�j٪߉� ?o��	4I�o۶����g.ă��ü�{�{E�y#LS��J���:{}�p� �5��Ve�߽��@$���$���n��-ɛ��1����0~mnRX[����{��cg��ۯ r��,n�f*$�I�7������&%���{��7+N���D��<�eG�vQ&��s��� �Js"#�<�E�lܳ��H�W&tY�����?��+Mh��So�͙�흐�u6��Z"�ͱ����XVm��=��rN�U	���H�>�>$|6��m���6�m�b;�>���r��g>�?�vJ��y�a�̸���ņ�����+@��[�!&�}�o�A���U7nW�P Ύ�u�wf'��nf�K�{v�af{!�ͦ���f�s۵�cf�EH�Yk�y��J��]�P|�9}�%B'��]c �h���{y�gak����b�;{�B8��d��(��2��Kl��{W�g=����w���w�����93>���Xޕ�����5���+�_���A���N�$i�� "|�)umf�����E ǯ۶�2��h�0|�e%��j�5����wS\�r��>��g�M8��@��>�yVݑ������`}�^���i�(ӢY}�	$ow6%cs���n��m��OBU6" DD4�� ~~1d3�w�e1�#&u`/�k#OU�In��(��F����0�Y�|�ދ|�T�t�T���ͣ���i� \�p���$j�n�x����kUA3�j��6Z��\����h�Tn,������v�;��>�����%�E\�U�L�(�޼x��W�X�1#$뉚�.�n����rָJ�D��k���Y��l�G^��H�����þyg[�Q]�Ǚ;&�`�RϞJ�6n�ʧ���xp�J�6��a46h��<����ČM��#��Վ%ۮ�s-��w���a5���,�YHvd%�r13�m%�W��)LmZ-L)�'{���,��9�ݮ����ړYn$7;J¨s1�96�!9YZ��]��5�P1�6Fb׋fi�M���0��t��0u�7���j���M�bo"�k&�x5sL3Sx�}Ip2i2[�#3��jnv�Ehs�<�h�V��4�^u�K�w���/m�{���Elo��� �  ��v��U0��a{�w9;2���3)�;���L���[kL����T�R�n�1I����:FB�!f�*�e4�B���ye'�OYW-G�@j���S�w�4����Y;��,S|�M�ó^��E]�;顷E=)�z��Re�B����y�P��V�Gf*�0�cM,�V��<�o8񷔍,�5-�ю���geӺ��joj�ի���μ�����z+Ž���q���R�g^�׶��C�ɨ�_�V������#R(F�m$��l�!���.z��yQa]*"�G9�qǟ;��QM'7 �[OV�Bd'R�sS �wCԓ�G(1�)�l(�Hѥ+LGw��4��}�;S�Vr�͉"meI	*%J�AK�r�{���N�GK�	Ҥ�2�L�/"�w\�p\6����$J����K�PVJMɻ�'��E���ʧ	��ET$/ҝ��l�.��\�ou�"9fq�Y$�,��%��t�Q](�fp��!BO$<��.����5�����w!#$"�4�($��ri9�fT�L����=O'0�;�24�H�M"�<�Ոa��9��P��H�$��\)$�y�NcC�:�P�>:�#�5wwwwwwwwUUUUUUUUUUUUUu��������]U�ս�ڻ�ו���Y���6ϱtB����7V�v��b�^�[Zx*������v��@<��xcۃ -��e�γ�G846��)w^�0mn1�7G��X��T5)D�ULD�Uj�P�6�r�L�u��u�����ݮ1�=����`�����b�s[[�,�n:�u[b̯c׷C�[������6Fm�N�:�=�������6n����4M� �"}���۫<��j��k��M�<h���n��Q�`�su�j��Hu��S��/�k8n޲b��Ѹwl�\#�^�$�/֝u�׶u��K��;�]t�Y8z�	����;����8�:D	��եD�i�&
볠��R���fM��F�4=�.����wK�֍��=\�a�Ѷ����"[<v�^�]��l�Y��ɠy�l�Xݲ�����n�gq�y����ӛ�K޼���$�}�oE��he�٣�OOQ����q���ET+T�U��iU`��x_tI�"�7yRN��L#޷M������s�N*π����r]���ջ<�i�6���P�u�ʝ�u۝ѷ��v{k%�s\�H��_ivyJ�yӛ���_f{NL�B��\���5Ӹ��y���ⵀq\�z��x�a7O'�����1�g��'�.7u��;��æ�<5�M�m�c�������7m8�������l���l�;�t�������8�6�N�A�S��qڐ�,�&4�����r�k1�.��/ <8��sڶ�y�\jÞw�.���1&����tz��;x�7h���F�%N�{��*5X��N�8��૮�V��Y�k8'oZ^�ѱ�a]��fۊ��Ƕ;U���DI�Xn7<��O%2�o&��p��`�� �%�k	qwlf���f���7D�g�anMa,���]Dk�*�܉tkZ����hk����j�����{��������^���Ex��7k,q��Ʌ{^����@��Wh��a۱=�����絹6�v���\OF5؞{5_�,�b�((��$�j��ZGϜV��ɺ�Q=b7��Ӯ�P�WlY����m={�kՅCC65��{����ce�ǎ�"�ts۱�M�Y�Ǵ��KE�s�>C��]���zh	��%�-m�%����~�?8�k�'*�z-Ћ��V[.n]�j��L�8��{9h�U$��w�ߤ� vJ��̃�g��@�{�J��	�{���͂֎��g�[�ڛh ǯ��$�U�yW��������{�|���]^�saO��h�I;}�`"O�۾�*h�u��.R�\���+..��I��i��p�]}F��������嚱�j�ڜ�$z��k�O�I�ݾ����W�4����<ă�{��w�'}������ ��.� >f���{� |7�M�������I�6�"�#��	Z��u�gv |7�eͭ��y8���$���4�H��w1��97��7F<�/�h�w9n�.���̠2�<����޻uuvz�^����!l����'��UM.�����t�(7+MYgu��ҡ�7�w�������虹������ ;2�߉�s���s9���;%L	f� û̸I�_X����D���:ȷv��ׅf�B�f�ʻ���]z�GV�Z�X�;�WHvҊMv�v�H]^��SW'38���L) ��z�?�	���=���6�2	/z0U�w8vjy��I����X�[m�������� :oܚπ
{cl���7�������@ ��˘
�
vFZ�����e{��dNw�I$����Oğ�4zt��I��˺�����fY$�=���d�1r��+O0s�Ŭ �r����n�!��{��'�@��D�/�c}ݯ/=�Vo7��Ϣ���
'�8�\�<��#sS��X�X��JUkN"�v�]wl�*ő�Y�3�EwOIP�I::L�A��Y��t�{����{������ ����f{�[����5��v������bp61���&�?Q&�Θ�&�4e�r�D�iZ�%����d'�\�����2Y���bZ��>�U�K��^�[�B��a�d�]�x��p*�F�H����d�%�qF �aL�[�zU����ݦ����l%�4⪼����x{ܟ�|��b#��6�n��%�.�*�1�mcy��}'{ZY�����t���I�Mh���7�;�w�]�O����jkI��N�"䆴��2� 3��,=�xb5˥͜���]g� wה� ��{�칝՚��8�6m����V�D^����.����N:��a���ݛɖ.j����vF��]�J�א>绚��|���G>o0�v1�\�'2���tCT�.#8�qr��V�q���a�o�l�˹���^�[�-a� ���@#��l`J'sL�\Y��D_'23��̊�[VY�7u;w��s��ml :�︽ٮ�����@��]�_ >�v�P�[��'	�7��$t���b����π;2�@ �=�fm ���Ʈ�8����)v�x��,�a��NK}p�݊�=6�ī�۸��|g`j��[�L�w�C�������3���"�5�xι7��<Nk<�	�?B{W��s�U�m��7�����-�����:���ٶW�=.�$���M~/�풡�@���|=��t���f�q΢���\���[�x���.��\�t�J}��Y�\f�U�{��>��P'm�|��= �w\�I$�Gg�6O��vO�_:����>F{����խd�2ttRV�b�^DC$OKU=KJ��I=�k��0�N�Lt�4M'��/w�t��\��@.�8ț�����{�������`��j���$+�m��TI�=�����o۹��=�)\�_��	_`�g�����?9P�I:buD�$ї�ˤR����V�$����[�}Iр[d�$;��` >�U�����u�q�d��� �:{q� �!��&���3�²�}S�0 �����q5JJ��T�yȱP�f�jZr4�(B��[5i����lu�ͣ����r��z����G��q;�UU\��^ݚ!�������A�1v{�i��u��MU��n��rnu���gllvt͸�ŷ^%�냲6e��lֺ����Ӵ<��4�-̝�����p�-��3�ǵ�v�kG=����n�c=��d	���:�;qOk�Y��Ÿ�ۭ��g���xmÙ�ηh��9��k��)vcY�#U�%���+je�f`[�ܤmR]�P�,u]�I�����ܜd��G~�V]�s�Δ-��޿���!4H����,[�E����iG����퍱w�\X4jE�;*�f�,�$�=����r�s�ЀI'�ܹ� ��r� ><��4��l\�)����[mh�0��
J��ߵ��k�5� n�*�D�S?u=�/(�n��H ��˘1{�-�c��Q)�HJ֫�׽����綉| ?w{ϖ�� �w��@ ����&߷��x?I�;p��5� ���m 1vJD@߹��1�Ц��k� N�.b�!r����0�21���[;��U��[�klg�ۭ�ݱ��1���C�{h9(�s��,���рZ�g_�<���kI�@�n$I$���7	�S�����eMg��Ā�7�Z޾֗{1�XL9f� ��m�',ozź��im�����&9̬d�mqx��4ugu���f\�W�^'V�W���w�`�t(a�Z/��P�)��W�#�V�`����/�ns����yn� �����00ja]�ۑ��YƉ˨H�F�faX���u� 3��skcg���3�� ���z���x	���"M;���&�cF@	�भ<m�^�����>  �ؑ$�k�{����I;=0��ֆ��> ;��H(�Q�8�	Zˈ]��>�� ����5��m�<w�@�{0 }��}$�vzc�J�ނ��k^���ͩTE��i�F������Ė.���^��Z���4:�V[b���vX�mϯų5�	�$MQ&����@$����n��g�̝��TH�{���߰߈�k2�ɼ�ĳ��қ�̝[�e 7�0*$�D����$v祠!,euE��9�{�u����RI(��|r��BI��u�D��[����2��b��N6�\tm>�QNd���Q��"������*�����a殽2孪�"�"��B�ai���sS  �ovq ��~�w���|7�s�4�A�kh��08{/���z��w���x�I�]�@L�i�I$C�˞��Vq���Η�w���`�kF@$�U�
�O��$�;��
8N�Rקt�~$q����4e�r�����\����Ӫ�+t��q��t��ꇅ��b��?���vD���pQʥ�������H��!+Z��w����� ��k @"_�,#2�e{QrJ���H��I��Γٞ�J�MO��k��d3s�E������{�>�I'�x�KO� F�f�@�}EUo7{��y�{���@�V�O��û�+�� ��t�|���K�ｼ� ����0g��{�i�.�cv��J6�����
���q�z3ٟ\z{�k�$���?Nmj��u�h�\�p�N�ʲ����������v.�)m���z�ẝJ���O�4��ֺj��/{���޸�&Y�T��>$�L6����bX4���[i��~?e��$��}���]R�s;ko�q&���n���Y�@|w��w����x疣\�~}���m�v�Յ�1����S����H�ό%���=G+���
�h�N�5%i��޴���U��I5��t�s�ή�߸kk7��vf@|nw�k��ch]��O�s���OīJj��=��;p� �r� �G{��x��+��|��kۙ��`.��x������4�b~'۽�T'�MuvΝ�K�f����r�$���ͭ��>��;U�l��w{^���u�� �ǋ�$�D�����H�=-��}�����nsz�c�K�4��ɍ�9l���>�풡4I'��u�����S�phK�5�	������ρ�߷4�o��n]u⼌��V���J�)q���ק�\�Y�)�h��׍)���s���je�'��ڊ�i�5�r�U��Uo����{�����UU\��픱ҏ���K�p��(�4Z6�팷]�I�q��tm���v�4	f�#b��M�+�D9����C��;<�5.;p�`�8M��6�:+��2�о�q�ԝ�t�^ޅ�m6]ag���I��{����ndըm�^�cm�s�O[lp�@񶞲E��枥s�ӈ�<�d�m�Ѫv��qsK�r��ֶ�`�͑��z�����Q&��9ۊ7kgl�X2{.B�8��Z�td-����/y���Ŷ�����A��{�Kc`p߷5�#W(@��&n�[媛��o7`Z�� �������׻�q�uuw5�L[��=��l	�$��K2	+�s�;��Y�z� 0u���G��%k+����BI���$�"֛������Xλu�HI5�s���r|��L�r�������3sQ�u�XȬ��c-,�Ht�Y�w���7��X���M+j�%MR��3Z���=�m�t���iF�9[���k,�E5MS
j�����0a�a��;˕~�g���Q��S3���KMF��<X��9�u%�d�Q���wZ�m�4����EEM��`�b�J��������=�^�L��Q������[f�4���MUC�����ҍG�*j�0�߹���k�?�]��I�{\3��-r�kL�$��7bD�����ٹn{v��n�ns��Q�~�ם�n�]:����3��c>�6��m�j��0���gk~�5��T�4Re5M[�s&�,����X���n�3��Ku{]�6��⦔���N�S9{���zf�T�Ƴ$3��v���i��h4W+���e�MQQ*k�ξ�U�8U�|����R$�!ݷn��b�0a=�!�v�q+�1w�9�S�%�Rp��VAG!�Avn�/K���P>d�.k\X6� HIk�,3X���?��mS��MS)4ST����yE��i����0���n�9�[J5e�j�gz�{����oާ7�yF]{ǚ<3mSFql�*:�7j�ق5�-��v���4�֚TTTҪ��'+�����ҧC)�N�SJ���͖vV{�ǫ��Kl�5Q�U���"�Ѩ�5T�4M׹�[J5�T��)��O��Ul�4մ�1�k��^=w�r�;�w��y����0��5L�{���5����iF�EWo�Ɇ��.���j4�T;�w��K:�����?x��Sj*iS�S.����ZQ�������Edwsie��1Y�3�*j�%MR��3��{�=�[j�9R��w�=��mF�j3��w����5C
j����c�0�0��5L)�j�P�1��u��B>�෮A;� �Eɓ)�9{n�����3Ś[���Hy��s��<k�i�����Kl���|?��w{�_��4�4����{��ʊ�T�e4��)�L����v��6�L�3�;�w��|x����Q��g�E��D��銚�L+��0a�fSE5L�d�W%7-˧.��#Zf�)��{�m���T�0���s��=^�w^~Q�g�8�����5M�j�'}|�����Yt�4�������Zj4�Q�̚����Vk��2��s��Ҍ�5�!�8�۴���M-5'=y��q;iSTTJ��Q*f���ii��1ST�h���	�37}�����)��ף�����c�'���� ߰�V�:f:(��k���Z��b4�n��!���ׁ�:��zYǻmRG:�:U�����~N�)E'��
�J���_V</��:��ʌjW��aC2�]�g��4%����&����nk�U�k6ԯ�њt˭�}:%/Q��S��3
�u���Fz�+�:Hl_w#R�j�z%�2�.�Z]Ҡ����fr!+�ɡ���Ά��\�Wi�=3ngC*m�j��b�jP�l����MJ�fsjY_L6^A��±�l�V����u���ܜw38��+����k
2�Hkb`V�B�o���L��oO��RV#��w��
��)�nU.��X��v�e��+:�g�g+��;�N�(�1>�ӌ!i����֦CR�����y�m�t:r�ζ�존0�SR5r��&�����W��Z�a��-��B)4-2:��]��)]G��qweX��F��=qk%����oG�Np��. $x��y�4�#��32�m��a�f�[�J�'E�of�[�\<̚'�P�IKV�7�
:^���?b�Yu.�������hw�a���M�f�K{��G�H�J�ڼ����c0�D��m��NH�MI���/Q��J���ڵ�%�lyP�j�
�������Uڷ���f��7�N���9�wU�4�J�\9��Տ����tj��P3eVA���d쵗���:7H����(�?I�������0��ADd���h�)�Ŵ�F�&�����A'Ú�y��:vD�'n*eiU�\ �vp�C�8U�jy9U8p��y���8jb��ˊ��OtH+ʹ��i��'r�M̜����j�rA4�MI'"T������)�*��	9܂�Na!��
C+�fDI��#̻�;�z"���t⥫(��BPO:N"�4rAwMKJ�.Q眣ZAxBBj�eP�B]Ԉ�VhR�n�'2�KWw�v>�{��^�a�Ћ��&�HgJ��æ����u|1����^�.��jJ�!0��.�ά*�������^둨f�Ei�Һ'�^aB�q����/�N&l�I�	K����]"�S��N:�ȊU�Q9	�UR�.�W#�wC�\(����B�e��y��I �UR��L���5e�3�������λ�:���Jʊ�W1C�#?�6�{��`-�3�4ST�0���W��`�TҍF����ߎ�h�͵Mgd�Q���U[2F�ŧMS;Z�p���қ�gǱ7��Ҫ��Q��/w�ʊ�T�iGL��2�w��v��Q��M*j��=�"���Ƨg0w��m�����t½�{�dh����f:�*U?�U�(�V�&�f{��ki�ڦ�aMS
j��ww�`�յ�=�r�o9����5�������d�Tő�T�N���T=�o��Kf⦔���N|D�����'A}�!̩�����_[Ծ~�Sv��`�og�*�ą����n1��������JB�-��	�ʚ�T;Oy��?�����a����*%MQQ*g���ii�����e�2��ǵ�SZf��j�׬��j�駰�\k��z�pa�a���aMSTT�w��6Ѷm�h��p��Zإ�ًo�����]�Iq:��J���Y�=�&��+���'���Q[J���5Q���i��m:iS)�J��P���aֵ���*j�u��G�6|��g�F	>�&�r���4K��֙����o^���a����)�j��ߵ�M[ZaMST�L���S�g���q��j�Q�ŧMSJ����m���Jn*iS�S9�{XE=�J�X�d�z�E��]�i���D��80��[�����T���T�w>�4�1m�t�MS)4ST�n��"��4�)�iC�>�D���Y����eVsp�~ګ�r�ㆋ�T��JN�©���(�(��V����s��ɚ���V&�n��Y3o-95p�Zy0�sb2Ĝl�kn��u	K�5��j0����w�m�l�T�Fs�MC���̑�1ht�3�W����ZiR���AQSD�/�1�+iS滎[߱R�������2�o��v��6:iS)�J��P���a�ZQ���MS�a^�9�S24ST�W������}�􍽨�pV�(D�Ed^��mۮ�bS��J�7��T�A�����ms�QBG�㒵��ƭ�M����6��m�j��0��j���u�M[ZaCT�4S)�h������}{vR�sjϙ�����ޟ{�⦔���MFsw�a�ZQ��jݺ���dws:ie�4V�}��dvҦ������S��G7�21����G����"���4ST�\�=����4�MSJ5�W��`�TҍFMST±s[��00�ůYV���� �}'�C�8��n��.�&��(�f{z�n��J�*iF�D���0�4�Q�YM*c�y�K����Zg��5Q�*�=�"���J��(�h�����j3+9ڭ�Y,rǔF��4S=���Nnr������g�mm��85MS3��pi5mi�STҍF�+~�2a�b˦���������ƚX�a�Tl¦��TҧC)��=�"��i�L�g.C>t�Yi���Zf�M�^�a�vҦ�J5J�T�w^�4��Q��=��1��7�a���Q�\�;����4�)�j�ST�3~�Y���F��aMSTҌ�u��M-5.�s^��/����~���tu�ݮ3�=��Wa���f\�h����KTnf�M��
]��s���x�����Nb���kU{�,b�y�1wwwwvU���na0�a��ʗ���u۶��]m]�Wd���\v:��;zݫv�r�AU������;w���n�G�9Ӗ����Ϝ��GF#P�u����G�/���-�=���F�]k�:�gUa�Ԧ�����k�=T��2�l/nÁ�)�nލ�,v\ymn]��:�#<Vw��Һ�q�.�b�۞ۮV�\]%��6#3dv�l�U�ɼ!���:�&SI67�R��zqb��j�e�����>�o��t�Z�l���|�MS;��p���4����|�Y���YM*t�iS(=�{��Kl�tҦ3�;�d���֖Z��9��������b�����fZ�e���Q�xoΩʜ�Ӫ�ej٦�f{�skc�MS
j�I�jgҍi���0hj��J5)2���^��Z��j4�Q��������Zj4��*iS�x{�l�tFLo;�)�iS(�j7�U��)Y�ΚYf�M�v̵M(�B�T�TJ��k�ƞض�:��e |$�H�;�n����WxI�τ�IT����,�T�(j��5MS
j������Zj4l�9�f�ۅ]˒]N>�=�2}$oRVbnryvn�>��b���TT�����b��:e4��Ҍ�����[f�4��:iSUP���a׹��45�]���}��2z��L�E5L�N��%Se��,xDk,�E3�޽����ki�5L(j��ww�`��i�W�\{�|τ�'�|'y|����.��*t�4�*���m���M(�iGC)��=�"��i�L����{�k�Ǿ�m
��-q� �Wd�S�X�<�O]��e�x�$���)S��j��`�z
_�����Z��f�5M(ת%MR��3]׻�=�[j�Q��M�3��k��ҍF�ܘ�������3ٿY���F��iF�
j�����6͵M�g�*7]��KfH֘��gu~�N��J5�~���Z��_�K�.�:C�WY�H�G�Ox��Y��k�Eo4$��=�:�rq���Sq�a:�U����\�՜���f��� ���GwY�VҧI�ҧI�ҦQ��{�;im�N�T�tҦ����jѦ�ҍF�j<gG7*��d��s�y���(�܎C�q�Z�2ճ�E3=�y����mST)�aCT�3���ZkL)5MSE2�����z��]V��h<4q�l�9�`jp�#�7�fї��2���߭�-Y��fF,�ݳ,`�������hGZ���CCb=���`i�c;���s/�;D���=���T�iA��k���3L	����tUܹ%�d��3�j�`��@�D	 �y�1�"=�g��3�=������@�40# ��A��3h�YiF!�����Y����~ߵ�r�k/��d�v쒋�znM�r�%��լ���N��77@d�L���>���U�udvK+ȍM��k�0�L#JF��ٳ#Yi@j0 �����c���M]F�=}���q����!�#�9��ї����q���j�����3L^�fX��ZQ�{�����,���}�I�L"b�h�z�p��d#F(�oܳ-,��>������~�����` wDd����Rْ4h�}���!��oܳCb�h#=���]�J��7Ȭ8�[�ۨ3�&̖�5��4h�<nsF��͢Z-����gȾ�:�x�ǖݫ���X�ʻ�c~8��o�����W7߁H[�y�<�6l`F�꽜"��J0�Q�|o�e�m��'�J����[0��q�3=�w��{�<��y۽�0ņ�Q����CV�6L��ܳCh2����� s��u[�̯\���C�Dpkׯa�4������l�dws a�LY�{fY�����g��������T���1�=cb�!�p7��r�h����k��idj4�Q�Q���C[i/Ӟ�9æ]�]W���UȥQ�X���8ܓ�{v��'77c��z��9(��U�?���ڝ�n�ܫ$��bFwZ��؉ ����,��A��d�}��1��f'{�����{�E1��`o��h�h�9ڬӨ�R�ee� ��ƻ���LQ0�,�:�5�f^����m�c86մ��`FF]�y�-P�A�!���;�4jr\�Ӑ���m��_]�I��]�g*�NU�@�4��kVe�`F�ҌCf�����L"b�4F�Lcm�w�S�Nۓ9�)��Db��9�r̴��i@j4�Q���C4��.ٚue�j��$h28��׹��^�k�z5�#�A@5���f�q�������C2��_��SOر���J���dk�\�}P�ɜ�O��n��Q;�U��k3����ΫL*R��ӝ����+���mc�����;/Z�o��B|%�	�0�5��̱�+��'c���tꭙF�4����{ e�m-F�깬���y���f�O|]`D���޳�-G�$5���F��"8�oW�_��>���V[�9d���s�	���3õ�
������[s�z��;h�N����Y�|6�Ϊխ���$������z�fX���j4�=�{�4���Q�4F�n��eё�1{w�g��Z���c7�n̴��iD�iA��{���i�x��Ӻ�$��4�hq�S��)�lEc];Y��NN�s�c0Dq��d9���L�`FFj!��{XE��F(�YU�S�yX�k��oe���9=ʬS��R۲��і��^}��i�#�95�a��Q�Fs�j�^��Os���e�")s�� Ѩ!��0�k��-堌�������ӕw�4�&.{Z�,�sÚu�4؆�Q�߹���1F�4F��׵�[؆Ŗk��i{Wls[�Q�������}ރ�"^|�{H�ū�Q���-�#A�ƏL��E�R����c*����V}��gG��2#��}�4��6�9Zk-(�1F���Y���F��0�ެ��DvE_� I;DU�����V�i%ïs0M�`-Ҩ'F1-ULWMr6�C~n�-yX+�g���y'ݓ�38�����Zث)_��=�uR�����=�y�v_<����{2]�����%�n���ĉ)p�sհ�u��;v���c<9��"D�X�C��7�4R���n�	����v����t�	t�[��9z��K��c�.�p�����9n�9�H�%�%kb�&pE�\�����[�4ln��vpOŎ��Akn��&p���+�wgֵ�hÍ�s�wV�t�*��،͑ڸn2T^qn��rd^����i���qp�G*��5��a���1�Z�>X�ɵ��;���a�(�1��\����������`��	30��7�ΌLkxb.C=���4jqA��{XE���U�ۛ��Wc%ռ��e��l�2��4�]��s�Xᴩ��3�LZa�Dh�u�k(���F!�D��ܳ-,�F!���޽ױ�����,�9�`[��=�:��t�˪��M�h�[� ���y�0�7���Cc���ع�w`e�C20#F湬"��J0�Q�L=�r̴e4F���}��%�ܶ쬢4e�3מ����oo���>���Ұj4z{����4�����0e�ˌCb=�w�����{�Gb����6d�0ު>�*�NU�@�4��kVe�me4�Q�����a�׶9�[��-�4vc��-�lY��}�2�6�Z��$}�s�� � ˳�%��gn\��wj�p���5�YꗲU�h�E���P�/�ok�:�uw$�!y��
���ul�8�ٞ{��"�! ߹f2A�n4���y�4�0#�s����L�s��-������|�,�FSDh�1!�Tw)�Ul�2�6c��pX����H��p�e}��:��v�\�L�b�hp�rV;��fث��-��؊�$un�_LS��r1Y�XּS)R�q��8g�Ƴ*�n������E�|o��4�Q�F�ǹ�-\h"b$����`-AD}�o�窼x�sz���~h#53ro����uo a�b�}�2̌�iF!���y�@Ŧ�4D�1�o\���{�[GF��F(�w��-,�Q��J5�������[ǸG]�쫩eʹ�M�h��`cϢ�Mb��G\���z �΅����F!�s~�2���������k��ea�y��=WĶ���l�FZ#D�v�Vc��n[vVQ24Fs8��a�(���G&}�k'�{����Gz����x2�6!���;�`-A73�a������~�}�[
�7/�c��NX�n1�ܺ����A
��%
��XՖ���q��U�����{�نy��J5Q���LZbDh�u�k(������{q���s
b�{͙bK)��6s��0-�m^J'[��ul���ɏs���Ik\���9����pc:�Cb����@�4�����Fn��a�F�b˺9�b�|��M{�y��Dh�1p��)�Ul�2�6c��pa�(#JF��{c<}dx � �8}�t.y���S�I��A�ATV�����mռ/UB7x`Ś9�oPZCل��+oT��ԫ	���0�X�`���Ū��G�m��5�� Iw��փ�q�lD��}�`�PDh��ư�yh#"�f6Ó�V&�+Ė�ƾ��걧!�OOV���6�4�=�oX4Ŧb�h�u�k(���F(�1A�߹fZ[�q.i�6C���J��҃Q��y�Mm���{�rx*��S��o�?���xb! � �9f2A������8���4�w�w i�`FA���g��-��(�6a���e�)�?�?-j���x�BL�Jݩ�A�݅g/m�����vKh[���)��=n>���?��H�,����6k�`�y�bG&{�k(�`FF�����#�5��n�?zn؎)k�� ֠� ��a��5�[ٓ8�]Wj�%������i��ά�2&bS%��z�g�����Lc9�a��#Dh��u�[FSDb�#��,�K-F��J���3}���f����kX�i�6�%���:�d�Ch��y���؉ ߹f2AƂ8�Fv���x��f:�x�dL��ϵ�[�db�#�ܳ,Chɬb8�%�)ʕl�4Ѧ��w���x�+}9�h��\F�j4zo=���ҍFd`C[�0e���Ab!!�{����Yֳ��u1x֜�'�����5�S�`��ݛ�k�,�@S�����ݩ�DY�\
�k�<��t%\&Q�(��Sk�b��  �~��#���{�"�F�3�b7$��WQ�][�fF,�ݳ,���A��ώs���-0��oW��.sθ.�dh�՜�(���F(0�Pf��Y��SQ��J5�{����0&}y�7������o�*6��1vh=��UV-з��t>�z��CJRYb��x�'�X[$�嶾M���k�"H"�s�c0Db����@�4�������0��z���-��(�Q�L9�r̴e�4c&߫ܢ7,�"4dh����hi�0�-Vf��M�J4r{z�-���20;�r�1�ˌD	s�� ֠��7^�*����o����~Md�o#�!QU���Im���f�Ʊ4��M(�Q���b�� 4F����α�V߫z��QlCb��1Fk��bK#Q��;�w���ū�]�T.ӫfH�6�Og����+�� �����0�7��8d�=�d3L���A��oXE��p�*�s�KlCa߻fZ2�!�bHM�K.S�*ٔi�l��=�u0�a�����Z�Jv�N�=^�(ָ��6��u�-G�$;�w�KPC�7=�a�4�5Y'zN�7�װ�CLEO.JC45:�̐r�\��i�R���lأv���mj��Z�sd�:�w�O/p�*�����Z�1ְ�H��l�s���;b��c��	�˻뙀���Neg\�sm\��o�7wVZq̭s_P��H= ��0�b.�T�G�]#K�H�.�n�ش�l�{�w�3YXE���%�}Ұ�݆k����Jd�ol�/FR�.��Ż��v$6�c�e�H�+��6f�n�z*={y�*�ҋծ\�f(
k�E��E�Ǎ�7e��/L����kt���7n)�L [��d'�����e{N�UCJ�&Xy�o��"��T�T�!�����l�Iu{E�Z�9u&'c�:'G�ig=Z�0]����چf��f(�oٷ�3.�[�T��_7;yWLY�$�]؝#n�f�'�LS]�Z)k8gYc�2c��S�']����]
��*$5ث�j��x��0��-5r��$ڴ+d�eSB��r��#���Ә��쾛�ԩ�j2���445cm��wx	`��r�f85�N�}��&�c}�vGu=�>�Vt��>&�4%�.�Y��s�ʭ�4��\i2�u0E5�݊@��fb�O]����kR�^�eugN��F�r�#��q��ޡ#~����^D�gR��u�0�WL�D<&�6�Yݶ���K��tS��׽Z�"�d*`#(��Լ�xn;�ZM�	��\��d��<���6����n��p�����Vзi�������?PкE�%�%E>���z�Y�E5��"��jK���-6G@�n)Ѝ�)�r�,1!L.�C�]�I��멪a���rI*e?Q9U|�T����L��-4���
�)�w"�)�^m+%f"v�t&�%Q�XPZ�]2�F�r�r��B��+�F��f��D�B�'Ի ����Q�̓�p�eʺ�#I2�)2T��ڥ��FBd\U��EPQEo<(��L9"�\�T-��9T�i�Z���.�HM|A�ĔR7��E�D�AI�Q"�-8��52eį'n��d;���W9?5�Y��QM	�<��bh�sBԣS%K&�ɦWJ+�KC(�V̌�H���l�M,K@�<�΢w��;N��gH�H}�۱�~s����������������������On'�rmӰ�=�uNN�m]FэrJ�N�H�g�%�c����m��onXK�Z�k�zL���pN:g�mS�m�#��+tk{wG�|~p��c/�/>�Y�X�N�����.9}��޳���Oh���V���cr-�tqβe$�[9�T����A˹�pX���p 2��@�܎����l��WOg��my����Y5|��8�V�Kmd�6�w�'c�%���;l�#�(��[7��ܾE�6���b���I�sز�!㣱�L]���L�OU�v�uӚprj������c���< �^71�&�A۳�<n�\A�0tQ��όÀn�H�nD�j%8�m������Ƀ4�׎�F������ɴ�t7e9A��|��؝�γ;X��޳��Nv�=tR�
���g��ny����;�!)�<�\ǈ�;��5v�력��z�����f댠��g����6��Ƭ���{ssg��\i9ڛuՍ��6�q�50v;g�')��FȖI$׌Վz�iݜnݬq�[�y�Ŏ4y����/�k��{7�#�.0�Gzz���5x���)�z/ScFr�az��^�+l6�n9���:�n{��v�e�7We�ƀ�ɺŞD�G��|�n�糖��d}�ۉ<]��l'�'EI��yz:�����Qz�=�l�=��[�x����cu�K����y��#�7d�u���c��8�N��8/VR����X��Ov.{r���,��<n�4�т�i�4o\4�ǃTv}2�t[�hЇ�Az;	���<vy띸ų6�t�q�9�[�2����
5��Y{1v㳭d�:rl�]4S7�Q��EĘ��A'J�)��{k�v�������\�sp�>É��鵛<���˸�Vg��^3�
�u�.�Sm�t��G7*&�6z����냷��\�`��k͑�(��&��G-c�����=�gWS.��d�s�+�\5UU_�{��{�k�ʪ��}�<X1 ��r������]�]�;<�v����t6�\/����&��[]s�v�=]ё�n}r�#��t�	�9�����޹����y���-.Y���^�;RF�m�/.��u5�<��s�5ֹ�I���,�eG�����;z�s���C��⎦�s�[Tq���7hL��ް����!�R�Ҵ�f�fl��f��q˗�͇�v����x���7[���0��X�a6ef�����m�;�����3昳�r̳#5Q�Ҍ�9�`��CDh����Qm#<���񜺞�@2=����a���J&�=�w����=�:��e]J��s&���s�c�$���\g/`M{�c�Dph#�d5�{�L�0#ډ��oXE���F(�V��y����h�Dh�2y�7%�%IE�VQ���=��!��������j1��޵3�g���󕾝h28�A�"�9�s h��L7^ް�yh#!��4�uշe�Ww�4�^�ufX���xCj4�*��`��h��4M׷��؆ő�b�=�r̴�U}ܽ�h��F!��5}���2��U��(�]�V���q����/D�D$[�,�H"<r���s�� ��h#!�sz�b40#Pgk��mdiF�0�oܳ-#Fk�ڻjz5x��>�5�r�li��u�E�;uٮӎk:Wfr&�T�Q�uZ�}�O��U#$�g���4Fc�װX���Q������҃Q�l{~��h,�xjQ�Ưۦ#��k�� ֠�"80�{z�-堍jb7&�t�m�][�`c�f��ҍw�;U9�kҡ�b��x��*�o�Yf�Y\2Ey���$���ֆGmmP�8":��4U��T�M��n�5�X��{��/�_�}_ >�3|�0|&-0�h�Dh��5���2�#F(�o�e��j4�}ޙﴊ��K���X�i @W��Q�, UL[%���ѝ����BA�o���#���g��r��=W|�����^�������浄[YM(�&(�&�9fZ2�/&�qr\�R:,���і��e�3�ɅBz��@ID#�����-a��20 k���h#�D�����u����[�lC�F�����b3��4��n�N�� i�b�=�2�6�ҍF�f�����ø��_w��Y譈mխw(���F(�1F{��ie5Q�҃Q�综�%���T�xX5U(�i�5O�ݒX3��xM�盬�]���v9X��}�{���nwW�[<F!�rw<�y<1�C`k����A=�wyL�3;�zw�XZ��Ɗ�ϰ�b1F��Y���F����?vK.[��l�4ѡ�3����a�!����9�ɵ���cX2�Pj0##���,Ch28�AHw�������6�0�7�o|�=�:�-頌���nM��n����0̱g>�bYQ��Q��;�b�1F!�_}�Ǿ{.�Y����ߴ�>5�@vļ@�Փ��b���s��,=W��ܑ�LOzĮ��/$��;�
F^%[3�]���ѷ�3+��� dm�������07ώY��SQ��J5�ώ� e��x�	S�U�w)�.�i��8щ��s����׌���y��$�s=͘�h#�f��� e�l���Fn��a��7^�M��{~��Za�(��c6a�m�V����J��e��F��Fr���4�i�&�m�ްe�4�{~�ˮ�k#kx����q������!��7^ް�yMgzo~os�}��y��wm�.�/5��gjoB�⁸�X�G��/$+�\2�j���t��|��/5����7VY�j4�PiFk��0hb��#Dh����Qm#�s��o�Ǘ*c5��Q��z̴�5Q�ҍFw��0-�bνe���:�d�Ch��;�#�"���l�/��gg����B�G�8�ɽ���f��`F�f���me�A�0��γV{g�������;v�rK.[��l�2�����]�i���҃Q����m,�d`s��<�]��]�U�4�"H{��0�9Gn��a�4�U�ܛu�ݐ�U���e1g>�f��j��z�5|��iF�Ҍ�g\��-0�h�Dh�[FA�1F�3��,�K��J�_N�e?���s�kTVh3��)�bVZ@��]��	Y��}9'yӰ�R�P�Z���0�I��4���sEL|��?������y��(�f�3�C4������Ӳ���˼�bE��X�D�D$����:�On��~�{A�����5�� i�lCkL�{Z�-�l21F���Y���F��/�4s��ֻ���]�]-������&١E�J�47�!�gzP[��nbv2Q�ee���{BA�����|6s�`<�LQ�iA����k��F�&Fw�Y��#��[�%w7�B��&�?�}�� ��Z�VI�F�7����ɤa[���j�|�Ƨ'D��ٓ~$�e��yh�N��R��2��
B�W�Q�=�葜�Y>$���0�D��紟�$(Y�,=�sK,m�eVW��q={���En�o+�$�}sd�1�vH#��V"��2_s���T7�{��mx�a�:��@��UM��;SX3���ͷ�I�}�`�5v}���Bk��8=��Q9�M�7�����\�]Neූc������=K���隊aujNU{!
j���v��Qg8tL��̤I0�ePa�R6����{��ϫ�UUr=���#�7j���>u�I���������n�v��K�'���=�����xv����b..2ݸ�:|����g;�'sx��qK�ܽ�6����ڭ�V��NK�Gi!C�ݺW���s�݂3�m<��n��u�{tݦ�n���8Y��7�(�^v��u�*.:+h��㞹��$�z�\�B�����6�ַDg�wd�36G2u[�R󎵪�r�v��p��j㱹�m^�RƇhJꖫ,�?y���Z(UT�6�l�y�B�%�j��D�bbz���ZSdjJ���]����dP�F���'M����m� �*�>ͬ�Aj*3P�[�`��$�Pg�&�9����s���H(^Vr���\	����<F��Im-���&�L
��E�.:c���D���/���� �7{�����E�У�R���������
l/y�b�5��@ϱd�t� �%���
�����B��P�w[W��\�5ΞA�x�+d-)*�!�5�5�*v��T�z��U;�x�Jv.qԽ}~~�m�'�TI�3F��]�>$��Y�	�6%��NUuU�|F�5x6���f��@��U��tA�}k�\!tnt�-�S��ˬͥnh	,��? c�`���]]���OX�^��_8A`���+sx{� �R�$�{�����&�Iɜ�4tB��w��_��TL��"�
6�����o��Gěy���K�5��<>���N��ŀ^X�$8��o�y���&ݙ�/Yu�G~�g�t�ĀK�w�I>{����K�P�3W�2I�K���E��Sk�TA�U�(r{ܘ�&���OC�P�Q�(W+�j��s�)m�q���,�x�f���g̸+#mg�`�'�`����bqG;:���P���h]��vX)+Z�����>���]�I��$v�<�
��!�������W�2��~��5w�^���
/�C�8l���k0�AW=p,�����@�Tv��Ȓ�޼.ZfY�4DM
��iF�Ϲ��<H$�{�s�ӫqL5�/gn�-�]���4��x�>�U6j��3s�1Q �RCԎ��|�*�n8�Y)���;wd���9�kK1���I W�o�m��{a{^�2^+��� ]ee`�c�7&M� ��UHo���|g�X������Y�X�$8�險��y��I��x3�2\� f6bI̜q`�[��a �v�j��x���w��܊ѹjvB��8]q���a�a����n�K��-�W:������w�-��������d���xH$��O0�{"N][�� {=�d�9�x3n�0-TLT嚻�M��蘯nZK���h��R�%��=��N�y�M�U�*�*%,46��K�+�����ci�7�w|G��Q1x�|^��>$�N�s�Q��`�jJ��I��.cY���
�:� �n����~�x�Y*^z*�ox;�(lk*���+�uNO�e�=�݆��d��t
d�1�!kv��qz�4g<t�3�˜��]�������s��o9^��$�q�(Q��Y� �U��b\��[R�P&w���I߰m�\X��0�9ޮqc�:�֞(�2�p��g�c��s�/=��l�ۮ9��z$E��B��˨���'�[s��Z�m���lP���Cu��P��B}/7@|	���e]�(LГF�D\r�
l��Oew]��$�m<�A;���A��`�ͦq�g�{�����	,�RV�<o��0�
�WB�㒄[���HK�wK[��5�k�~�R��
������iZUqA\�e[�I��^E� ��:;%�Ð�ʠ(>��u٬��ff�4*�8ݹ$�ɻ�o�w|gL��D���� �nKȰI��wJ`Ҝ�
>t�<�]<�~�U݊��kH͹�	:��:[��x��-��&�&���dJ�2����Vm��+�F��>w�I$����m�ڣ�KS��<����{��sd�mtO+ۀ+��M:�Ƶ e�fd	\�)a�1?���;=���,�Ӹ�n�f��nv�L�x��p�&��i�x��(w;����5��(�͓<t��k<�����IZMr�Y���u��:�Nu��;[�X���م�c]h7<�і���hk�����mŝ�{j�a�&�Q�h�u�n�p�mv�y�d]�͞����2�4��P���\��{ߕF�B��O/�$���$O��<���,�R��=��o	%dY ua�q4b'�5U���� ��&iA��C(�$��I=r��3��`"��u�"�js��֑b*��3����Y��v0IY�Ss�����Is��>��y��"� ұ��3]�����Z���=s��1��$�|���|D�7��\q�+�?���M��|��V��J�f��ʈ��Q��j�Œ)��	'�{��������I,�
f'������[��颠ݲ0%��=�=mƋ�.m��د��5$�r�%V�3=i���u�>"{��a��<�yŀI>�|�	���ʌ"������W��D��>�o�7����=w{f���8����+�fJ[R�T��բ�wH��83jL2�㖻^v�q��ü�^�:��//�x 5�%	>�� H$���f7�%y�m��.�X!��Pk�5Ux��0a �.y�Ė&�<������.��ɼ�H��.w�n�"�H�>��*�p%W0��H=�n��Rn��=���WT'ιva<�M�)�[-��W���ؚ|����h���I�=�������mua.k�57��v��t��������!T�8�zb�|G��}�r�]��6ef��ϼ��[�۴Q��[�	��c���`���z/m_f�$���@��"fY�"h��X%d�I��y2��}��Wr`P2{�?��"�V3"�1ܻ�����9b�A�&`СF�]����lA'�D{���u��?z�xq��Lu8S��#��;��f�⛽k��W����wQ;�9od�[{�gt9��9o�$�[]�scz��P���\͜36�AAVL��"���c��:�/u��Qg:�]��}���4����9c�U�ְ�j�䜱_lۮ��P�v����rDvea�)0��]Lo�"j��$��;B�{�o1�A�n6�V�)K��T�\lm��v�eˏg;�s7���5�,���M����r��4.�^������h:�2b�H���է7V��DLz֖�ډz�UQL1{�	�l���\1��{�ltN����o��>�
֘�WKy�y�ܓe�i�UR�qG�N�ڠ�is{u��Bm�h�Qa�)�)��0�`�y�QMӪM�!h�.芍��m��5j�c�P���c+e�\:([�J��A7��ʔ�����G�W�֒"%��������Z�[���80�0f�ĺ����-�{�;6͑mz�L���6�u,Bb�A
.�Q:xT�)��kF��bi�����Z:��ܡ����.��p��{�j	HҖ;/�N��a���T�٩�;W.b�R;1�!9bvBS����t�0ݯ��x� }�ȥ���1�1�iF�X@�r��fgX�z�z�X<�6�e��:$ޓR[yh[�"���Q��WW7L7����{l��ij]W�^���,v��i��u��w"�f�y��Md��m���%\6�=o��6o���r�l�A��>��wI,��J1,�'�h;PI����IH@����D9Ar�8XI](�ʅi~�ү惝"�EHt���QE	Y�RId�Y�T+*D$�(*� ��鴟]«�I(����U��¬�Z�DYYIi�&�9��XJU�Th��.���:r���BA_��*�w���P�V��fI��D�"K2�%"��EA3�+0�BJ��	Ԕ5Y� ����e!�R�I�bHjr�UYT�&d�NV���+��$%J0�DI$\���KE��L�S�R}��8U�3��.Pf��Ҫ,4S*ٕkVE�,�E��r�W��E���2����J�V�b*k���N�Wg�w.�*Ft��ET\�1@I85#��I ����&�{�w�~��f��3"h���U_9��:��S�Ns������$�y��Wq�ff�O��=�%�j����Ŀ='�dF�����:��W�$��>WN�v�w��^uH�yb=��tƷn|v�sv�Ì�ʽ���q�4�u�'=���5���\H�說�4F���}c
�;`A$����;-�;�9e�	J�� a���:��h)]�Z�}�ϛI����5�MM%�I���`�����ŭ�M�v���c
�12�DLЪ�4�v��6݌�w�#Wb�a�o/4�{:��$��x2�κ�0$I�4(Q�T�ف�/�u�Z'ǚ��G����Mrp!��t��*��!�>����� ��j^_3�8�_k�
{G��pP�Kk*�za�P�e�ᯬ�Z{p����E�.�+a\��[t;��WDP3��x^�}��̏��?Dצj�����A�Y� Jȇw�7[�[��`�ۼ��Nw��g��b��l��U[iڶ��(�e���f4nvv˸�ge-�)ݶ��+[fh����hת`����}.�	5󱄓-r��.{�NI��I�Uf�I:�<`E���;��5��6/sb��A��r���-_MO��M�@$�\�=�՗�-�"0�
ۿV�(�81R^�� �D��a�YMرi��]�$�m�x�L�����&Y�"h��Y��ΙJ��.�$�޼$2�Y��H���%t�O���u�$^�����e�b��Y�2�!/�:`V�\D�k�O7w�Y$u���H$M��A#s�M�s��[��v�=B�<$���Y��+T�.�l��ܶ�;U��tn}�Py�C��������l��F����}Q��(�Ň9�������m��Ts��,NF����\�-�a�i9�K��n�;v��sy��u+��9�h����n�o�o�9�ذ�y�=�7�]�6�<ml���u�r�_n�n�U,�ً��/`{9����F�l[�`�r�ڎ�v	v�e�X�l����ݗkv��df��`�3�pg����m��'Jmq���l���/�T�]�N�A�.��~|��1�|��Ke�E8�#�]��W��ѻU"��r����ƻ�è���\-�~w����k�5T��y�H��\���զɬ�*�<������L|Vu�"�>�E�*�Q�uuS�*.�>��A"�{[*?d
�/�u�s֕JՈ#�T���f'{�w1���6}g���K���:��`>$nOl ��ީ�""��_��v&�*;.GM��0@엱`�H_<ɫ�y#z���v�W^�s�(���qN��BH#�n�n�vF�%��ĳ%�t(
�w���������`�9wf�gV�w�U�κ=M���f��G�����V�%<	�2D�A�G�\��I ��۫ ];�������%�c?/�G{+�hP㕙C>yx߽��@|9C�����U8��Y<Uml���H���t�rk	�y���{��h�}lWk�z�B�*��1�I���'�\(
�{��K{�� ���ŒO����"BZ0��@ξc͹Mz���=p�{7���P<�=.�6Q{� 9�B����N�Y�"@��FbH�6�q���s:Mݬ����I �|���|H4���`�D+���c�ȿ\x��h�ث8pbK�� +7�?��+�x�`��>���A!ro=����u#z�ϻ��9כ��}d(�d�KlUD۴]�<7/=���ua�7�)cC�%���,�6��뮨����$�g
 �ͷy�I$S\�Ж��v�P���2�L[�9����:���Ա�V�v��ƚ�\��-Nf�EL�*آ ��x	�&���Jʧ��	���=�D��AءTx���buy��go�?����>��o*�&dJ���d�I���A8��f�:�W�s+��T���T6]w����b��	�L��=1��ۇ&m:xW�Wm���� ���a�5��a��"���* ����$q�=Vڤ5��O��ח��%���
���C�����uA�MW��6A�P*�bH��|�	 �ko�jR�j���NM� 
�ک�ZW��,���{}Y�K��Q��N4��T�'Σ�H�<ض�6U�]�]\*?�>�4:���Es6|�=X�H��UM��A �6�$��6oTݸM�Np�^�]���7��,��B��VccH��^���5 ��� ����(i~�HZ�VZGq:��ߔ��c��M�F����>Okx�����Ҡ���P�Gf� ���|�;fɚ�9Y�3�w�����p�洪:v�)ov$���dX'���1���mpV!�ܧ��Nҋ$���8ȣweb��Q�{�%dCJ���U��k�V���wuy�uh�6E[�1�7�$�x�;�L�X�x��#%Za�䨒k_^x�%��=yf����]v���ȰOk]�d[ַ��3���;������u���k���`�§��͛�v��p��)j���y�g�*)I#Z���o����-�D{Z��	��FLS�߼�:��Z�Q�T�E���`�Ym�`���w��zI!�,�$��f8W=�\2��uWz��"ѩ&��
��En�N���>!�0�SqN"'2�N�vM�!k]�	,��$@�2jLУ`���M̄�딾�5n�^#9.�>�;l�Gr)�=�z9��O�f$�@ό�MfGvf`'Āq�x2�+�1ِڌ:L�j�$��a �_{�y�:M���Yxj�6�ӓi-��I'aŹ��݆�P5�����x�*s4%�����+�V*���N�([��-�TC�����wZX=Ε(�c�J,_׽����UUQ=q�p#�ݞ�������ף�����ժ1On7N��nb���\p�1����&4b��h���n��kf�|�W]c�n�cm� ݍѬ>.�"^�E<6��vy�crێ׎�g������8j�:�.y�������rm�ĝ�$�,t�+��8,��K���/9�>nA�Ԓ�ڳ�*��)v$n�Yg�j�:�l�%�<��@��QK��i�᪻a�nn7��q��� �v:|婖T�y��Ί
�D�?�f�X@$��^$�7�w]��OZ��xK˔ }�ؗ ����"fH��g`N˽���<����{yu��>������t���u>�p5+�'���%ꈙ�M5}x�0	8�x0�H&`�>�e��R��k�>$�\��U�RM�Y���	\R�dǏO�ZjL�+/6�A9��a>(�l��QܤI����@�r�fx�b˩�(سxl�V6��b����/�qy��~�}X�<H�M�(�l�'wUF9כ��t�8WdU����(�m�3��
;b�D��$�j"*Y�[k-�ί&��Q>rb�:��A �.V0��6��z:hM���3��[���������EA�_�v� �Q�%W_�f�X���@�L䳗w�����oe�LS,K�_Zl��H߉�Q���Yݑ_v�]zrh��n��7�ּ��ĒH��Y�HQ�l� �.M'7y]̞���P&�fH� �_;
8����k'�x���� �k�Y��gl�#"��@�����������݂8�[Jv��| W��A(ų~$�ֻ�9"�������1"jI�STk0�{�Dͧx
����
]�HY�gl� �k�w.fX�Տ62c�Ѫ�`W� �T�2Q����T�����*݂yƊ�nn�&>��5,�f*�&hQ�vz��Ă�=� ����*ݻ��W��v1d�"E�pl�^Q����~�Ķ��aN$~����ڠ>��N����WF1na��c��2�Q׈Fy!@�ֺ�Ć�w|�Ң��:j��^�ܫ�o��Y��D���ʕ��H��8��L�v��o�(��գ�@��Bb�����;�ܤW.uaOٗ�L��"��
~3��_��~�or�"gpR��f'o���f�""��MW�,�;�$��ـ�H�5S��G��g=^�칲z.0!����M5w|�0�I���2��qn	�eL�\��V����'� ��s3H�-���_&���6� ����7lfN��N�{(����#\j�(� �:֞��d@\}5 �UUEg%�ؠOsN���O��|Y�5��V�{6>Z�f0a��M��%U��k��;8��-��l�|���$�i�X0��\��
9�޷4�o�nJ�i�[����m��kk��5sq�pR݉T�#S]�A�5�a �d��0`�x��t���NIqh�L�g^Mwr�������O������ç.�@���L.�'�f��;"�UX��x�����TF7(WL-mggN���f�/-��W2j�<4�]1޼X09���c�F`MD��0���AQ��v!�����I5ϖ
���J;t�B�}��k����z��TݵH����q�f-4��u�n��9�t�q��U�����;~�$DѣUK]�$i&�` ���`��$��fp9���z6�C7�͊��	\�R��m��jw{�Z3ۼ��i�o��n�$Z���ge���;��D�K׾����X�ySD�����/�&���y�vA>)��s�e�\�Ē'�ŉ��3�V��t}��UcNB��֚�<+%��+2���}y�I �vU���o��.�9�Q#[�|��V]u̘�QW�������מ6*)׋d�О�������F6���[�����6I�M��A8��d^'���YH*b*qay��pM��*bLXm�j�L�/f����'��w�3hu�"�x�	��T����{(ɲ��i�d���Qt*E̖A
E�3W�qh�rm��s�^6�̝��[�m����M�9f�C�Gγ	�<4�]�y�t+�i��Hj�d��j��ft9oh��۬��_Vht�6Mɸ�'JD�R�SmSʸʓ*d�t��:F�V�+��[�r���-b�aw{��WZ����8�;����mhm�+�QÕҦݎԕs3w>���Kq����[@���	�z0���Z:��c�͛)�9ݫW�7+�l���HԨ��N��XN�Fް]�*}^��h���JGZ1͉!P�YW-���n��Uf�Q�G]lSy�j��_(�|���.�L�Y{p]¬���zD㭷38ktR���к:jiC����W>��h=��	:�72�&�{�Ўbٚ�m�˖8��������5�NI�r����_k��nؼt��"I.<v>ʺ�	ƺ��T��/s&C�fQ�'f�&�:����H&^NZckjp�J��`�f.�ʛ�2�ׄ�ᷩ�kC3Q��fkn�����4
�n�ؐ.�\i���5�:�,�)Q�)**�������MG�����}i�.Tsl�;d�T�n(�;�͸��r�w�+ͻ�y.���E��h-EU�Lj�ff5�@�ه콤ꂡ�TU���1_��g�$a��ȅ$��02(�V�Es�y	��Q�!��r���Ru3���øF��Z�\Y������E�]i,�,�$j"��U跘��$Ctr����\ΰ��T�%LڕE$Bi%)��U�fME�ԈԬ�YV$-EbE':��eWU5+D̥EԭL䥔y�m+i(�s21K���Z�d��*
�����Q-B6RJ����.���!U9��
��J���"��UIYd!�~�]RKK�Ȯ���d���ҋ�C�Trz �t(!��s�B��E*9s�Qs��hGe��ȎQL�4� �.�
+�QQ�˕Q		QITEQEb�J$�*�Ђ��p1���n;m�=���UUUUUUUUUUUUUUUUUA�����S�%ľ����ۮ��Gn���g9�ȵ�U?�Z�m:-τP*���Mq⩵j6��K�q��6w�|�󥐭���E��,X�p�=���D]=�Y��ny�tu�ƽ�ɩQ��w&y�WS�ۓ����QVɧuڮ�d��Zkr�SM����E$V�����]�P���צ�u�g���-�S�������>Ho���^��,^�d���8ĺ���<e�Ls�m�qsۓ�\쭇��[^[�)��E�δ���{n�Mԝ�pY7�n�-[g�Q+Ԫ(.�6uq����k[����N�\�Z�`�ݜKY��=�L,n4n�ڂ-m�i�0j�j�ڣ���^��av9w/J��=]N��!6�l��Eth��=��n�m�'
8�¯���<GH�5-�!v�o=�8UU���u�ͺ��H�Qx���=��q��A��@�BW��m����77�;��L��v�������7&\h'l,�z���L���TƎ.�r�S�n��\k�7�o7;Z�����g�:wn���̕s(��rXk��9��x��.et��oh�M�-�]���ִ�Lv�.��7�ד�\�`.�V�ƻ7a��m�]\7n�N0�z71z�;��6\u�qC�m�F8m�=m�n�Xݻ�,��q�J�ի��sw��*=�"�;��N��	��j^��V�㡸�
��vpq�:�x5��x���{=Ӟ"�����M��M��]��ךM�k�4�5FܙwZ����F�LF�s��N��]\vΞʈ��gO�n�����(8���F-7zhu1EB��ϵ���t;� ƌ��{]�q�����F�:����n�kp�V�k��Og�	h)vJ�;m�m�9�=��r+�Y�Q)Ϭ=X�½gb']{�ձbl���{7=k[6�{v���:����/L�n�/Xu�%痵�ִNqn�v�]n�z�Z��j���r��UUDu8�۰�狷���z�.5��knN�|#���nm�<-]�I�I��.-vyl���'�qׅ-�}�㰠�Ǎ�3��']�۷�n�.�I�ɳ��òGd�5�V����w����Olq;���ċ�-v�Ʒd�iIv�n�uۄ�A�MPؐ��ַX��r�$���i!�n���ú��U���l۟j�34�{v�4�xݭ�����s�7�k��g��Y��檗�;�W��_�&XԤ'��d�<���d��5ׇ�kj�*�)o��,M���s&�ia�4.V�Z+�]�lXz�k=��{Џ(�0��M��	�v`"�Wo\N�b�~õ� wMH5USY�Jݰ(�A\Ӽ�AY�{�Q>'��M�	�6�0�i��5$,�-�I��s�[�q��o�6����Ĵ�fx�M>m��ELUqsc~=�M6��su���3���ci�|ݼ�U�^�"d��ֻ0���Y|3Y�Nk#�rd:,uP��+v��l�y7\���ێ򋊰Iζ��m�v9Z�mDۀ�;��
�0j�xk�� ��]xI
|�`��'k�Ul!�� �w.��r�"g��HO�>z�ر�M�z�Q�z��=6q ��+�i�w}���h9�������q(���Z�`L@����PF�eֽT"�ܚ�ƛR�c���4����}x	"���H�U�Uܼ���q6��O���-��{�Xɤ��>'���J���ܤY8�y�
��w'�5�Y���^^7��������^,QS|�����lV��<�z���ůs��[[��'jj��k�
���0�K9�b��d\Q���{7��H6�<�J��������G)�����Sۡ�mACry�X�R�T�ժݔ����6v�Z��9]�[^������^��0����H$(�ٰq��2�m�m���>$M��&A��"�L5^6Y�W�$tVCX��2,�w��*޶$�M�o=�Gn͂0��҉���դ����\������f o��=�
+v� �O��֥Ğ��8r��7.Z�]�EUV�y�Q��V3&�i�E�.����O%ǸWl��u��V�6��L�l�xI��'��Aw�st(?��@3�
!Q��*j��v��4ۭNu+bǉ1:�{	$��6	'.�b���l�G�&��`�?Y���^^.E�
�\��.g7{&��3	�#anȰN.�6&��B���PO �Y�˲0�\/N�뫣)���^�9v�Q�Qm��"
�Q�eͮ�����4jU{����I,��$�q5ـ���Й���(S#j�X���6	�C�N�"���r{[�m?"m�;�g�=Գ�@ ��ݛ$�5ׄNu$3�72��o���dE��	�����=j�3Z�V�7�J���o���ȲGk]���תH�����u��p��sK�I�X�	����>$�\�Z<B�)����wC��$�]W&
��k}�N쾦���
+3 vd�I!%�@й{j�Cq���ų��[Ý+w��G����W����Rd;nJv�핁W���H��Mf��u����X�׽V	%�]�J��kTMƓ��z��:Z�ڻge�&�&� \���-�yluj�:��y�{�:JWe���T}%t%�^���ޖ�Ğm;	�4���ow'v2�*��:�I����Q=@��4hEMzʜy�A�u�n�u� �)Y$�w$�a��
w^Ul�&,k�v�kN�Bm8��;��� �O��� ��́�T��;�f6�w��3����B��ߟ���GM,s5��{���$V���
��ZWi�<�`�T� >�ɺ{x��a�Lϳ�k�>�nX���T�$^�v` �I����
��	�t�S��(^Ku�)1g�vhsw9�H#q������7zQǦ�=��;
�L���S�ˬrp�]��������m��i����,�����e�����Fه�:���ϭ������>6�$	��;F��vx7Gd�N˫=;�۞օ��6�ڣ�F�:�Xqټ#��^7=�v�g͞	7p��5������z�+on=y�Y��n-uv�#�n���닖7Y�GN�;ڝ�&��sm�A�t�Zŋ����2f3#ku�뎂;6:���n}Ps:�e����	�v�8�7e�j�C��V���g<ޓ������.�=>�>���"$щ�O��}�0|H4�+�|B�ʿ{g�׊��m��3������h2*�MMMf8�Őz�u��[wQ�z� �}]ܳ$�׵~$�QK��1փD�K�EA�5��eM���>��$�;ݗ�+{o%-�M$���=�����;�@�q�!n{��T'���F���&��f	� ��^����c��=�v���׻�ı�H1��R�8�}�IY�'5�����ͅ�r�n��������=k�r�4���f�c�Ս�Y�-e�mZ��|�[��*�6��	Y93f�ʤ���y��~�$�_����>��	^���}��`�9�eի��Nu�y���j���{/�@���y����eo���F$���L����:"�ރ#/#%�jRe���L�2���-s4�j�Z40��AVr,B�*�	S��R�t�DӬ���?m*���	!=ʰ	'�k��Ai��mE�k�-{�l6d3&��MUf8��d�m;H4Cޜ5�
z�t�#V�Y$���1h����3F�T׬/r�}�U��n��>$@���E%�,�S�3���I%�r�}�;�F������3޺���j��Y��OU���x��YV	���I��`÷wT��[��ҺቡU2&"�Mek!V�-�k�c��3�����'^vW�'�p�n�D�51&MW� CW�dsZ��A&��xr���,U[(�UՓ�|;��1���v�_�	>�O]�wK�=���dA c�ـ�L��=��]�#�&�R'�ό�A�h�z,+���|O���` �Ü��(_j��Rz�CT�D�^��Z�,kN�eY5�E��a���BڹWϸ�#�ظ��"T*�lv+�4�?���V�I7���M��~�.�l�\MIP�ۘ�����9�b�.k� 	Z�<	��(K=��Mk��[�zHV$� �/��*��tw�_)�T���7�@5ϖ��A}�VuA�����Ʉ-$U�
Q�+\�W��g�\�#([�"	΅�ď�%cVEkV��u��b���1�EVB�w���r�#�۵`�٬��nT�Ywٞ$|k�<�LL&���2j�|��#Cg0B����8��O�&�7�I �5�O�v:{e�')�=)D�16�/[��:�c׳��6�\[�,�A&R4;D��>����A �.yT� ;�by_����,����f��2֊�Z%j��g��	)�Ւ	��]K�!G�w4Ѫ��fu���R_p�jb��ٝ�k�7��+� i�32�z4hξ����L�
ZގIf͊�ҁ��k��E���X�}0H��Bb�����~�B��-ʝɨ�2O���Hv-��}�{�﷾M��9���P9��5b����c�׮��鸶M�2{']�LR��Z�Muy�^M���jk��f^,{b��8��`5�n>슸�����$�j�'�F��!�(�H[��%�bǝP��?=�坹ӧ��fH+;(_���4���� ���&v�x,�\Ng3��{9X|I׫�	��:����u����ز��[�c �&����BM��
}� ,����G6��!�I)ky�$�m�c�_G^��B�Ud�nH& ��r��⳹�� w�s|QX+����EU�$�}V>���<I>6���jo�һ�v�W��-*���T��:he��������j{$Ʌo�|�<:��=��F��w�m��ۤƸ�]~�<�*�����y�����n����ؗr�2�\q��u]R��l��]g��=95��^vo4x����=V��W<���m��NV��+xJS��2ru,��9���1u��׶-�ܾ*n&�j�탸�v�e��MT�j�v��uxz�3�����X�nW�	�&]��=�b��z_O=���ר���Q�cL�e��g������^���z��yO4v�����$}+���˧����K-�����i����w�	$[��v�ڨ��J��SY�������&��������sH71�Ļ�$N�;$s���O���߫ۨ�ó�/����xޫ�����I���4�x�o��*�qܬ�{U�Q˷S��Au�`$�o��1	�(�"��|>��{�ޝ����^ 7%�K��	�$�쥻ܜCž&����!eW�D�13��{�Bŗ��n��S���}�<E�n�K�ʰv��MMg�緪K\!SvW��+!ݡF�Rsv�D�۝n<
 ;k�v0C�Ie��}��&�U
�5��k;0E��a$�^vU�����:e�g:��Ni�@�m7��oL35b�ea������m:�s��JÈ�x����z����3v.{���e���1�ϭmOy=y�32�>�����N�Ezߠc�k���V>$���`$��<��ʈ>�Iá\qJU{�eB�T���6��wֽdgF�q#�U�8��@�H��`>$�� �u�1N�J H[��=����[Ǫ߮x`9�z�fa$@=�*�'�.�ȩ�z��Yݺ���(鏰�K�.�ࠅ{=�� I����`����K�t�\�0�|�ʿH�k�<a�)�\��d|Bȣ<���Lu����8�&Z�ļ�/on}sz���_�����^h3��o{=��,�$�3���$�aR��P�����bʲq�H2(4*jDע���DH���v��l�{|	�Ǖdֻ3Ĝ��P����\�͡�c��3&�EMU^ D��A �{ɀ)�R���s��X��L�:$^�rr�Ķ�'m��<.9vnkT�}3��̺�}����ɝ�:��[��G����L��^qOFƓ��wY�j�iw��=���}!�Z+����)Y�XXQ�T�����y�u��9�.��b��ꬮO�A�y/�#�+%˹�D�+�Gj��{#���(��<jƾ����ᕖ� ����}@k�GV���PR@ayۯ�2hKl��7���V�x��_e�`S���o��֜L���ׁEKOl]�h^"�X �)e�̛�K":�rR妢�۪v{�D�G2�W[+%��h�M��w5L.�<�2�%�����vMQ
��|�šd˩u��tZ�[��b����k��u�V����a���(�"�Ju�[3�j�����t�P���0q��o'��v���w���l����Q}KFj��YS������%�����w �T3L��l���z,�{�0#MY����]���ζ`��Z��Ws��j�݁KU��Cm��Q�F�%��G�eTm�.���t�ف�ݼ����)����a����m]B��1V�^HD~��C̞��:w��FR��hz��5�r,�x�b�h3&#�±b�E���z3�Đi��h�z7Z]|N,�Zγ�M=ƁS�-Wdy���q��iж5m-��3��Ei�w 8rЙC�VS���3��F�4�4m�i�$.��T����7u�>��L��k��W��i�Lދ����wC����W;�72�i����ei�A�(Pij�F�&Qr���+�B�D�"�L���e2�A"T�B**"�J-j�h>^�H���u*�"���y�p�.Q2�ue��3**��tVt��J�TNd���GtJ�W�/E�jL�U��J!����l�G5�)b�*��iZ@z���B������Q�'+9V�L"VFefr%��S��Nw"PHL��U�Qt�'�����4�l�O�U�r��(gB��);-�����䨅BfwD����ԩD.Uȫ9GP@�:Ӧ�J!Wrs�Ě��]�P��.�D�*3*4J�7�N�(�i���YY�ʎ\�"j�r���ؖtΐ\����9Q2Ե*�����W*�
�Ts�tD�R�H�܋�t�[.$Y.���B?����||�?H?��X$>־��>z8ԡD�B��׬6�0g���]H��b�>$s���z���;���+:�EѮ1EJ H[���f,M��w���9�vs3�r4�*� ��`�M>kuR~�w�ɚ|���tq�������U/�i6�=lq���)��=��i�9X�6�o���`���n����Y�wDsyu� �|Ո��	�Wl5s`�F�]�	&�Z��	�3���׀a7NV��Ed��%�I[��A&�5���9pŃ����V�?.��d(P��^��}h�I�����4�uP'(���Ox�syu�%&���Yʷ�u���ۤ>�58wk'Fގ�t�p �6�	$�/zZ���YwWVGp��T�tn���zr�|���5������}#��hY�.AE*c���#4WD,͌�u���	Z>��(�B�T���7٘@$s�V\FeNwtvO$�r�'��֧��������r�u|l~0�̺$t-��qq^i�^M�2���c���t{lW:�
v�������箷��m6�y�0J���x��J��$����Kw��3�jc��I(��O����ӹ��2�jqu�I4�+�@'�3�l��z��ԍ�8� %I�q,���3��m�<� qm��+;���ч9ɐA�MXv���FH�$B*��ע��}�twYu��x���� �^=���u�,ݖ�׻������N��a�-�qHB�[�N�*��{��߮>%z��d�Z�fB�ڿH�k�W��7���}���,:��m�Εn��a�c���Z\;!��E���P^�>�f�cʲ�rf�XIme�w͝U�s����ʪ����npn��$�� ۷`^:9�C<u<Z۫v���mڧ4=v9e��-�9�q�Frj���l*��p�P���Gcl��:)�ǫ�\u���c�^ܻg�����j�<�.�)��:��ps�Uʎ6l� s�6�I��\�/]��pmq�&�]�3\s�����j6�����M<Fz�{�Q׿�|/��Mz��M�z�i�k/j6�����y�2ۮ�Y�Z��S>c�G��c-�BDd�V�|]?Oʶ�Q�R�m��a�;n�$���=P��5dhu
�׷�bϚO���6�_4@�UX�G.7U���ߨfa�$ztb��� 	z�f I���S��Sɥ����oj=fjA���b�9�u�$��5�ov�(n�HY�VH$v��3�&���֝R���c�s��ܖۭ��s�kSn�@�����QYw�WM]`�K]�d�'9"`��hME�E�4�fI4�M�'=!��}@�1P��ẃ@��3��D5��zfB�)F�	kA
�R뗞x�;A���<�h,��ֹ|�e{�;1�&~�}���H���ST��Y�,ͧ`K]��N�����d�ݪ�@'��f�uL�ZuKY~�Os���<�k;�ѥ������ﻷ%�j����+��:��D��X�mܭ�2�Z�p����qii�Ŗ����T�_�<û�6��9߄�v�X ��{������3Q��Oo�����z���tY��"�H&&&�۪�^ �k�{� �s�IE�"Gz+�{�СB�g��l�Ԃ�V�6�W}u�����>5ݽ�F�&��*�D�]�f`*M��vQ7'��}��bi��7�|�[��I�Y��7י�>��g��;dM�VDd�-S�!Y�ͨ��U�et���2���=:����`ֱ��U��>��pw�\�5��U��$R����ٰDO@�3�Ӫ�+u��<H���a
��&L�T,�}�mV�D$��W���[�Y����I<�\_l߉���Q}ݞ%��B�2&��T׬�^^Y��`�.��Z����2�>���D�˩E-x�_FuM���NF*I��%�*2ȼ[�R�;�d�{ѹ��ḙRe��"�F&�����$�r�g�t���6��8��T���Ļ/�Kn��֕ �O6>��� M���oI��j�Y�|�-���`�P L�P6f�M�|u��Ѹ�mm�l)�]}�O�.-l��>սن�ʴ=z�7��w��	���Z�${��9�uq���6����9�j�	c�%�Y*���2/5����5mv$��kf�$uk��I5[��U�h�(�ٿ���&�����X��sw�^>}cz�BޱǍ���w��p��d�Ѭ$�Ϋ��фyԭ�]رg+9��c���9��0 �8^Yp��yu@q^��=�7@���h�2jL�Mz�˼֧^�.Oax�KlQ�w<�@'ƚ\X�֌��4i5�{7�Ք�ޫ���j��reJ��6��R��G�X&a�������c~����h�L*�[�V�T�K��QY���]�}���ᤇ�i=_q���F�	n���y�6�N������@�=�L\Rv����{�O�N���G"�w�����m[K�E����qӥyz,�X�tm�%��L9i-��M�^"`��:�@���x�K��|I�k�<I �k�� .=�9�lA���	�7�$#$�Q$L�0���A��o_d1^xfz�G�f&� �k�{"���o���S�=:	��&	
M	4j+�b��`�AT��0�|Dթ��@�)d��D�3�<��At�f+:\̑3PhDUZa�r��:ۇ۟h/�� ����|V��� ��_s����j���I�3TE�י�	 ���Ԧ�+�+��n��:|��$���2aj�����w�w�5��/��CZR��ś�9�{̕,}Ԫɺ����4��4|�,�/M?:Y�ތs.�����f�ffU[���m�ܥ��n\]�����
���k�a�eP�˨��l����.�j��Ѻ�C�)��N��6f{B�ڬںqR������R�gzyD\b�۞H�t��ۖ=��xU�WW+��^����=kWg�`��l� �uq�wO�����ۋ�,�ޅ��<n�x�󸌽���qqs��ls ]��[��Q�ɺ�TFݧU�KgR����7]sە��Y#)Ă�ܜsl��<�m�/7�me����g��F�	n~����6��.Y��[�C���=��P�/:q�_�i���ŊF�c�Z����5��1Ңr.�I����>>T�s�ⷶ��7U70�����&�D��*�&g�:���Z���;��{�	�Իs� ��'�Ӓ&	
M	"�W��J�f���t�d$�ѰCg�  �;�g��Z���gH�*~��U��Ne�B�9���w'T0�D����㼶�Ēf��.�V�>K�{s�kuE�cqd���BI�huz�8q��հaWs��77lݨ-g���[cT������^� ����I��}�<M�0�I5��=���[B��W2�}U��{�I���z0��\�XC*�LB�!���Ph]%Zɋ��[�suˣE5}3�\���y�G��p�+Ǘ��v�+�eEꊦ��A��[V	'ݚ���m5�k۞��v��y��F̊I�Y-d7jş��ׄ�A�9���>�˴�H<�Ր{5�a#f�����	��W�ބ�)Y[αm*��=�I�9��3�ʗj���S��	*[��!E@PHRhI*�2��׉����M	s,��;˪k�;U���}ݘ	'��]�����ڨ��{?�����Z	O�&���p���F`���H:�u������?,㖝����X��z����IT�p0l������M��w�洛ޡ蛃�rF(����Q�:��sY|/��4�q#-���)]����۵��b��'�e\�UT"�&&�3�]�� +�=���`�s�1y=�o.��gE9�S��#e]��E�vr���hΤ�����!J�8:C
��g�.�LYݾ�6����tG���d#AԾ맓�;O�	!J�s	�&2D˩��j��ǭ7��\��vH�wo<A'�v��	�C[7�^�����v����6O�u��,miKe\���"j��0�r�s��:ٰ����s�O~��
���\�R;-��D���ͺ+�� ���=��pH&$�LM����y�ߜԟP����o� P�1��zٳ��t��s��	.y��X�.�`�3Pj�h�o4Q!��ڼڙ�T�1�d��}ѱ^������Ksæ�$�$���-�i3;��M�?sz���{測1���Y�KI$-�$t5�&�M��Xj�6o1OgF����G`Bbm1C��- r���u��S�^�VQpLt��d������[$$���)@��$��h2�G��j�n}�N�XL�Yt
V�5���w���_��c汧#fO��Q;%��?ד�����k��y�J��`��Y�H$8�d���߽��<�i�{���� v&V1�P�W!�n�ѹyt�΢(��
,�O��U/�v9P�3��2ELԂb}��]���HJ[t	 u�v`2�&�DF�܍��8띌$trٿ��&��&k�u�ݘH'����6�C~��{ P�K@\����2�,��mԥ\��e����S4o<l��z�v0�aݧcL\d�*Wgv{��	.���-S=^51��U�;�笶ʞ�{SىU
���C�]�I�"$	>���2�A�Xl
6o1O���;Ѿ�ފ=[q�v*��$���ـ Ʈ۱��髩<�'��%��UKn�kw!���S�]����ڲ1-0M/4�<Sr�V�#Z��9ԶHHC��kh��8�|c��[��$㤻C�kr��eD9��v��ە� s2��l����1e�%1Y���xm��2Jpn���ѥmm�{I7�~I���#׻H`enB.�l�vg`P����(�Q7t�e_8�نI,��W���e��U,o�v]���uݷ0�Xlt��J����J��|ٚT�����m,���,�mP"�qt�iua�Бə�=��(5L��R��-�yV�!�x>�ͺ}*ե��M�3MC-E$E�q�T��͊RNCIn1@M��QxF�ؼ����:����;
!��:�ޠRw-1P��s���N�Z�����{^�W���j�����".iާ5Y#Ca/eu��ӕ;aSw,�x�:;jK��\f��2�E�lL7�kS�k�z�7��4�U��`��.�n۷����}��N�����1'�R.�t��VA4m��	�HnE��DʋZ� f5Y�L�ӗ�����ەw�%k>/3c9%��(�iܕ"b�/Gom�px{+�7gf7����eᐷ�����2EL�9�s���t+���k0٣�����)�.p�Z������(͛N�W�m�x���o��㋓T�pT�X��s�1��E[�Č4Ds��fͦ�!��] \I;ۚ3$���Ѧ)Z㨔�beb��=Ɨ)��}yi���g2_w-�A���	��bt`�� ^9��z������!����[�#���ۜ�9��u�H̳FeQ����e7'!�ubY�y�KNQw0�Ay�L�\�\�AA�*��\9�Z�)hp�1
���=H�P�"�,9"
*���#��z�q(��s�k(9G(�r̃1�\�����PG�UERha��*[8�t�;̮˲��0�**#���<�UD{����4B.�S��a]�z���=@�z���#Q$�S5���r9d�4t[,�2U1w�
5��I
�2"�EȚ�N�*"�QAr�J��&:�s��D
#�\�Qg�Å܇'��EO3�A�r@��(C"�S(�HT*���2�ȹM�D]���r��P�b�G;��(+�${�<B���*2C*�ȔiĒ���U���V��ѯ�	8��I�l�N{|��j����������������-]O'KƦ�Z��rVwX���na���sӦ�e����h`��:,q�ϋ�`^�D=7:n�w<��ŬW:�׃�L/m�rd#Z�]��^��q�I�
����
݋�87��]y�ݳZ!z�#�\�K�;ݓngq���h�ݐc�a���{;Ϟ���ٷ$�vM�JsĜ�6���[sֱn��{S�5:�N:��jz��=��ȗ��{�y��
򥔗c�&�Ĝ��d<k��<���\D�[nx�[�U��a�܄wNu���X]g����a��@��66���l��]�g:;���һh�cV��	OOb��	nݚ�����/qX�;X� 6r�.�<eB�wD��\��ʑưq�񧮍��ǂ;'#���p`�dW�vݱ�k4E�C�d�ݒ���{n��Ŏ�xK��tr�<��6�\�yN���
�wa��y�]=��[��Ѷem�v��$N;r<;:7X}�Z�p���o6���k�R���mن�'*��-c̀؞r��ۻu�"�Ɲ��Ǵc�ys���k����6�֍�������k��Y��n��N�y�t<���<]�8����7d -�.M;�8�	&�Du�f���w���p���v���`�m��9�z���u��&�u�7�n���=6�6�9|wF��Ν�d9v�3�ݱ�g�G��ɼ�Ÿf�.�;j��՞�ۘo]��1�br���2n��m����R�z�q'\�#)g��g6�۷[If}�EZ��q�x��1X����`	�6������m��^�nӘ\F�/7�n��w!79t�nI1Y|�fۑ��NB��n׺:D7���0��v�-����$��˙�����E0vq4�&�H�Q��w��R�m�33ū:{NXڎ'��͕�Kn�;v�q]�x^�ny��'��@p\;����	��`�<Z�.�-c�7nu��Mi�t�0fg�@v�$�����򪪭��;r��OX�^�<�]�8��"H����)j��n�%�Xn�.�Z�VCX�v9�u�Î��NCW����ힽ����͵�.Ⱥ�8}N�b6�lk�w{;��-���^�,��}��%�k׃�=A�;]@<�u��J�:��m�a��X�a��0�u7-��m�i�[���1`ی�;
�'c^�ѝ��N���V�ku���uC��Z7O��R��0�p7�S����Kj�-�����J��;%��'�}�}Syw�ibm�o��gϡD=v���NLM���罘��13��e�] o��.�6>�eY�ٔ]��I�|�	 ��ۘ5|�(�O)-����d��A���m��>���H7cuP���:��|H�m�Lj�N����"�����w��K�b.���8H5���	 �ܳ$u��h3[M�v�y�����N��T-�i�30�ۺ�O���ڤ�Y�	�>0���Р��_�/v23ųˠj9ir^��7]��:����t�Z����<T��\�ͭ�߻"et����.{Z�cm�����AW�V�m��=����y����{	�&Ш���j��땋>3�A�V\ML27�΃�y�t�H�;Ʀͺ�3oW+�7��X��o=���Փ�Y׻�K��o^��c9�k<��[˄�T�[H&y�� �mX"'U�;�O{E�]�r�I�}���}��׽Θ����� ������}�n<Z��>��`�I�Y�VHΘ$��4A��߅R}��j Z$�kO��mz�{��w!�f/.vj�&s��|�e��d�	����ǻb����F�5��mЀ��fH��� ���3�s׏5�|�r�M2�:㢊֫��q�=>����j��\b#U��Hʙh)e�^\'�uQ��U�.Vfa�v߬��|�_7C���`���P��� ׳k�׃�F��7^�`|.,.zg�6⒝ (k������~^6��*�F�s���"��7U!bvKSƽwKM������'Ɲ{g��CH�^�D�3���VlGmEe�"a�e�4�Y(�>��yD�������h��޾��Ɇ*���W���7�/�������_ٞ'j��S騙�$��0��l^Dl��}O�����O��ˣj�-i)U��00H>B��'�2��x�Sk)�R���1����$�=��1�;�s0�tu�5yQu�R����_���!���b]u�Z�w=p8סgg�j]ݩمz����,ԓ&hMT��bݻ>'Ǟ�~�D��0�{w���2�_�)j��	z4T_���*�f
B_6鏆{a�F.��N� ���$�-r���Ԡ�9��Ͻ&�Y�Z�,�� �f�vcZ .Y��A���*͕�^��[�$��r�i��dۤ
ݒ����8���o�E&� ��x	� �6�Y��B���0(�וS+7��C޳ϳ��s��X"ť��כS��R�K���\{�j��Z�ܝ��'�y��莾�j��L�B�&��|O���3���s騙�$�������fİйd6ϲa�z�ʘ�O����gG-����q���>�D��[�@j�����Wk�uF!�n��1��@���g�W@� ��UG�O�e5|H*��I�%omY���{�}S�����I>.��1���,�y�x˛�">���ڳ1�oĂA!�k
�ڰVlL�2�r���M����OV��	i��u{���ݟR9PL�Sn
�}�lL��!gmX3f���Q��D�MM�ˀ���s
%Z��$�������ۯ��B��^骺��%�|fIS8hL�&�j��r�gĜ�}xMj4����1����f	=��`�O�u�aw�X۸w�<3���҂�vu�+5�R�j���S�*%mx��:��Ղ��4�(R�[0��c�!��,��]�Wꪪ���'�a1Hqt������7��cl]ojF�� �&�j6���cm��plr�+�Y�>2�=�L��K�i���;mNu��g���}3�bǞz������v�۷'6�E��=c�&88�,6�wV�b섆�g��J7C/;ִ]������_on��<���Lp�J�e�nч�,�{nn��P�v
>�u�h���Ò�:�� �k���d��'"������|ɾT�E=s�[3!sM�}?����U�׾r�k�HZ�şGn��.�'UwuUv��{��di��uxy!���]�NR�^oy����f;q����	=1@zN�`Uǚq�!gf{[��EI2f��L����o�@#��x	���L��=1Rװ�j� ��}���LԓBfj�Y�y��5�]����b��'�L��$$�I<��cӵ�Ɠ]���ӜQq��[R�X�w7���A$�_��Y�+�1`�� #�ʱUI���BĚ=��/�GeewG�L���kƕ�����%��ЭMJ��B�
��X��v���2��C�-��M�����}��r��}��^\�U"%��9P�~$�g���2ր>|^��h�E��CxU��Q34I���.���z!'P7��������3|�MظJT5�&��[��#dnM�6��Qs.ť���ڕҙ�%�H�kilg����Y�գ�s��u��~Z~���1�����}�VMk��<��הrk<�����V��O�]�ﳫ`���d� ���N��=t��Uz�����-���3��݊��Kd�&;�,s~�Ǻπ���Ǵ ���b ��iSZ�����bk�$ђ?In�f� ��*$���M�̘ ��Z�G���sc��zl��D���v��?F�Ub�e�h���_ST�����dEM�x�@[:�3qd�1��|r�۳��r^�5}��|��E+jBXg�{7���7�=̘$ >{Ub�%����3O�wF�G����"��&�R*ݲV�������o��YM�߹ȹ�}��}	$�&���-�I?v�� "L�mGf����o��Y$U9~��ܞ�)� �ʴ�&���a�ַI��=����SYw9�1,�gq�ն�jT���c���C>^�;P��t�F���ta��m�t?.ֳ��@|~��7�?���=����|������;�o��+�ꭀ~$�&�TI$�I�M/�N~̌@|w�^3���Ecq��S&|i�T�$�'�7��!��%�h����-�I�M���&����.�"��~~��uup����惇�B��)G�i�'�*�Z�жk8�����,����l�o$�[;)"I4OI�7*�M3Oz���]a�ɋ�������E�p�*���s�H@��Un��^3�w� �O;�+�>#��{{�c>�Շ����u��ֵ����&�R*ݲV�>ﴫ�3y�f���9�iuf���o�BOĐ�Ub�MOG�I��i>HՒES��Aܞ��/����-��{���*�_ �s;�� DC���-]��^�X�J�٪2#*�u�N� +yt��������Ƥ�f�RR
q;(:�%̣{;�*�S�����*_�Q'��ث����D��&���e��f����fu����;�iV��=����� >;o�b�{h#kv���ӚldLdj� �ז-�u�#E�	\�*�P��FB:��R�|���EF�;d�O|.�zZ�@����=� �����i������T&yV �������	�����nk]S �iL�����<�ز��OĚ$��z@!'����`��ZL��I6sg����Uv�ܵ�Ԓ�>{Z�s`�{��  y�#����IOs��	���'3��Ȣj�j�L�uZ��cs+$$��=����;KtI�H��Yi
�����C�#�B3
��b���r�k>��qL> \�*��!�oVi���jt���$j���h���qy���3!���U��v�SÕECi:�g6bG{����E�7qW�^n�ނ��
oϯ"YOp��'l���w\ay��������_k��m��v|6�u�p��0��4状��:-��v-�N:�=n�՞���ӂ�9�a�wc��h梶7L�7��z�v�8�m)��A:�]ƵV���,Rrrf/�_o��;�û`�O`ޓxG/����!�qh��,u\��iݙ�֫�t�#v�Ϟ�yx[o&ղ0���R�ץ�׷b����s�㭸l���,ڵ�.&8�7M��':�ʭ�ܚ�c`�{��a7k�i�7��������pO�]������2`�H��J�N���6WM��~��@��iA��o��n9c�Jd�,�����Ǆ>�yl�.�u�Ѐh��=��@#g�b$�~�����}l7��>�n2t�D�VYt��rfd� ����- =�rC�޴��$�I�:���dH��X����6�kv�%�����̫�w�� �{x�������� ����K����P�����U[&ʤ�;I�6k˕*�MQ'�\��!�����@�Y%�&[��TI�j� ����c���s�� ��nD<���ɫ��N��=�.���2�-�m���IQO���Y	P�v��dhѿ��Ӽ��$�MG2�" '$�'֎N���k��5�s-�I4=9V/�g��F�D�d�&#Z�}��_�F�Z��ĜxP�ER�v��٪���1*�I)6;{uՊGy��m�F�.��Xɡ�R�F�����xST����`O��L�ߥc$�MP�9V ��v���A$�y�M��mK�m��^�^���x]�O��H�����D��Z˕{�=}n��\�$�]=��*���ͭ���d�u�,��!��p����K�>��/����;��$����:f{~; OG���Jʽ�-l�����{u��� t�s�=qV��s�ML�X�M{w�� O[�۪�VsG3���d�Z�q�h���U��V���TӻC{M�q�2Ѫ�"[)eή��RV�vX�������y�sٵ��fr�'A��wCN�p��-u
^����wr���Ǫi>��g�_�`t�w�jj�t�6��/{*�� g{�fo���L��{q�ŞrVq'��u`�I\D�#���ul ��Mg�|�������
��^��զ�T�M�+o;6I�8y������A��~�P@�wM%�H�򧊳6NZ���i�H��
5:���M�P��V(�Q�XH�1�Z���ר�j���P+���R��@e��yCG��ITNMޙ�/⥏,�*$��_k7�;ךl#�p�^ S �-���.�'����A�9E�rKz��r���QҎ%�VdXň*��R�hʊ^'Bu(�Ug�]��wj�f%�VE)h�k��h�l��k)ܤ�y+��)vF�45�hD��L[+k`�G����T�0zl�4s;L�:�����K��K9�S�����"lU!�Q��2Bf��M�2��@+W�m�`��!�����uc�Jos�����A۩n�U�%Jg�'RtX���6F��#|^)׀,i�c�wr�]9�u�yJz!FM'��9*�^���r�7eE:�`�`ÏwT���8,ȆA�-�ǜ}��9"����6]�e,��uz'X�W2�l��;]��u�<b��>�]z��y��q����{;�K}{2_�]'U�4���z��1_h��Z���)�+6�nS��Tzjh��w����e/��H�#��A � Vm��5V�ITTU����5������e�η3����,�����duI�ׇ����ٗ�fs���An�$n���MI] �Lˬl���鋣���+x��m�5bSo��=vp�K��2cxu���W�U+{�Q�f�X�m���.�BT?(G0�IC��"s'$�I	J&Teyؐrw\��9LMJ���	"߇�������.pp��
��:�\�n�G!�3#ReD	��J��9��;r5&b%)KP�F��y��!2�����wXNQAy�N��QLN��H�\
�-Ec���
�N��wVS��N	�����.Y˕Owq3 ��ʰ�N�ĽSP��J�EÒID8��*�A:XHr���ЮWTu
�nen��na"
(����E]��.�J���.G-O6GL��a�Z�.Ez rB,�rJ�NS5�Er�L��h���� ���
9��^eˤ��
udW*��ʡZUUD'�Awu���e9�t=�;w8�E\*u�8p�z��gS.��������1�4�>{��I$����-��?rfO8ն����jbB��K�oe�%%�ƨ�KO�؟I?z�m�H��*�{�ZS�[�(���d��9�Y;Tn��.<A�b� mw~�KD�ѣ^��H���gw�����m�A$�<�:�m����_<p�<n�ڻ#z�8�d�,l�����ܼ�Х�m�\͂;]-}���ת�����|s��������ϔ��[ߪ�A_yrj���L���{���0�}�0U]&ʤU���ѭ^U�w{Z�z����^��>Y�[$�IyV/�$�g�\��n�G�Ka�ti7��[O�~1��{�S��D����`D-Г�z�UbO���t�f��J�3�x�nq���}��K������)͢O��ߴ�I�H�ʱ|I�MO{��m���]G�1%��y�2އ6�N���ٜ��j�D:i��Ȟ�eoe�q�ٝH.��,C,IG+�D�f�;�j(��}��8~�$����,��<�ڲ��ۓwzZZ
$��ws����_\�d7�Zߨ�I��U�����2��W�v�a��o0��[�ۙ�+��=q�lӼ�um��O[s����V������іˍ��jk�u��ID�Mw�� �y��:�����b����J���"o�TP�ICNr0E~�Q�����&�46{J� ����kc�ﯞ��s]�K ��ٹT��]�<k��sC`g��r�$�U4�u�K�n�- �C�������w1침�8�K_�_�bA�=յ�R{Y����p�ƪ��U� {�����׷8�Ϊ^e�d��	��Һ��8���	]D�&#]�{r�$�'��h��Oy�⮉#�Ub��	����I�^���i��_�*r�dy�3�e��n� ��wL�;v�H����B�'T���6�^vo��S7�n���0��[��qa/���{�j�;~_{�z��m�ȥ"M�n�� �M
��G��ܱ�r��Y�P�;tpf�⃳�:ad����v��n��[4Sp�WU�R����9;c���2�6&m:�b{�{�ҌG��>Yw��r�m�c;�p�ۃ�����t<����@���uuعpVu�n�C���=���la�󑺽'X�y3��'k�ۍH��tb4f������Wj��DqL�]!����Z������:�@fH�g:�M_����ޕ��X�]���szZZ�=�w���I�9�S�"6����IQy($�Q. 9�����w�u�yEF��eǈ!��V2K~�c��W:ŹZ��I'��{��A }5�L��Ũ{��{&ok��q]���ouTP�IC0﹛��� 5�b� o�֏:��^�!�͙�w� |gy��{b;5�M<*��nTJ&���tkW�zj~���<����>���ЀI5�]��d�'�a�C1�O�zI��F���K~x�M{�W s|�#�|<%ݙW�>�O�=��I4z�l�{ߴ��Ҋ���Z�V!�\��FW�[a�dy.j��S!���u�ܾ.�����\����C�[['۞Hֹ�o���^2I�O�O*�2�Ǔ�=�}�ix�=�{�� 4��l�O�"�����.yR�4H�=e0>6�/�5q���W4��Hn��η�N����}�+Μ$r{Uo�ݳa�S;��]�T�1�ݎ*z�MS!�7��,]������?� ��rf �~U����B��=�e���P��X:��pe��ς�˂ 7괴�:!A�fv��+��D�I���t� ���*޵U�M���I(f#��H�~QXo8�ޕ}D�|b�X�~$���$�_{�d졋|-��GK�L�U<�YDղי�{���?~&O{[ْ����D3�]���uD���*�D�I}�B%{������S����U�
ڡ+��^&��W��{|�:w\Z�9��닚n[����@�;�x�<���$�RnRD�'�Oޞ� n��~I�&ϭ?[�A��$�X�|M?���'3 7�E/{��M���#�"����o��āRnV"M~==�J����9�Ze��ovm�d����dV^Ã1ج� ��ގT$�Kr��ཫ@�n��(4MFc��o��Q���Ω���.�x�>g��^þ�ټ[é�y�V��è�t����G���ښ�x�Z�~i�ϽH{�*�D������.o����V�l��!�Χ�	��]����)�U��@s��f� }
{�X�z��ݦ���t�Q6&�C/eUD�(c�w��ll��b���Ss�O
�~$�<�I'}�B 'oϓO��>s��~֧3+id�N��/�X��v����Ů�a��]&�ۉ-���������ȕKSV�N��ڽ������ͭ��5[k�l~7�H&5X��@4\����kQ4�Z�C�o�X3�Į����]_�R�+iQ%���;k�m�hSZ��.m>L��+�9���P�����K��*D��v�`x{<�U�6�+%I?���W��&S��ʢUt�ܘ-wzB�/_+�7s�a�����l@/Mw�1 �~�4��R��8b�=*���1�z��J��Y&<:��z�H{K/}���eպ[�6�t�R�>>�Y:���U�g�=�߹����K���=b+n�\x��. _�ڴ�{\:ׯwWzD �=��O�4I;k�m�h��sʱQ9��.oڦd
���%�BJO���J9�v�%��n�N0�<�^�'F���Ư�����k��'	C<�{���-�<k�˂@ >{�U��2+8��F�e���Ï���?�&,��)�T�5m���\״����yيLƩ������ zk�m�I�3��������BQ�j|�\e�5-��|3��p@ \��$@4ML�G�^�w�t�I����0m�{����cj(pkd�Sk���+��[��a��+�������I���t��������}qD�1�bXyd�l��ʫ�v��,����}���=�=T����8����$�I��Ub�OĒ��t�h[�>��Y~�K�]����ߟ�J��l�_W3���^ڻ�}�� ��Bz�:�K�{D�N�o
]�Z��/���|_�?�~~__UUU*N<��!������ֻ3q��={+Ƨg�;Kݹ�=�(a�)��M����p#p����t9�2O5t����y�hw\�؎��3�1ό�9��6�N��F���\�F[�6z�\]���No]l:��g��ϮKs�s�˫vx�]lfp��cO�1ی�\�z��,���s��z7xНr;�#u2)q��;����W0,l]�;vŊʼC�@�ۇ�88�N::�0��Wi�O���ߛ��n9�k� �1� ;  _{�$�r���_��^nꢯ_� �d��I���7c0
,^��k�B{�5b��Ң��q\�9�[�������σ��E��^��59���[��y¦���� ��_"h�L��9P�~&���r�ߕY�X��~�I���D�{��Є��*�B��[�� ����ݳ��~� ޳&��I��{���G��ws%K�Ɏ �Z�<mEml�j9}���4I'��x�_�"h7٪��$�)L��'�I�wt�B V��3k��7�v�'ӻ�r�����;���t����	��y!���$�E*��z��uYT�Ut�ܞ�wwZ����ml�f������b#���D@�AIs�旪:b���,��9��ϐsy�y�nAMm��kY{s��r/N<����}Sxa�X{lN�w�v�m˓�v&���ޫ��R�Κ�ⶎ�Qb�y;*ȅ�:���7���@�������{#�\�1`����"kSSy��u�V���BT�v9C1�3{��}5�b� -�tu�V�v� ��E�wI� �I={���5��C��ն�3�|׮�x?\��;(�N��� m���Q$�=��n�Ē��k �$lu�*�B��[���w=ۂ|�.��wq�c�#�¼���k|ߤ���'o_Z�����,������u�S%iҍ�p���R���[�\ ����)�촉<�ms�WE��q�:2��~��E�{�����猒&Of"w^d�+�B{��'ЂHrk����oy�����F޻�z��R�iVO{9� J�kĒM'�$��e;t��N�������*�K.<s7� m�o�KC`x���y;*hgFQ~{��z�3�B܎�@�2��c\V�4qY�ږX.7Y}�rYtxի�^�^*�ζ���s�V}�w��s� ����, o��V���U>v2�b;�{{��ncb1��3D�I���I$ў�t[��wid���pP C/���ƨ�5w�`�3d�/bD�����}������o����d�٘� ��n�gy��ka��f��H��B*���
�X����jpf���h�)���B5��kAe!*矸&�}(IZ{�t����o�� �=��%-�v�ǂ���F�m�I$��] >�̉��і���G=��w��s)u�Xo#�I �N�f*$�'��{��}����5��޽�OУ�2�ª�ܘ;���� �9���� �jz�N��'��I��$���I$�=�l;����r��	mǈ!�������D���	s|��| w��s6  �:��[�+8\pl���Q�'&���4O]x�.��[����Y��wkf���@9H��,�˲'g:ĝ�.��ԟ,�o����j�m�I
���8Kg�F ����%�>>����I&�y�� ���t�4H���v�û�^�=��K(�b�*D�
��pQ7id�Wqm��N�6�n@-jJ�$��/;���U9m��H��T�$�L��9P�j��؟�Ȭ{�<� ;pm��D�j��wI�$׭	���a������=լ>����oۙ�@� ����$����$�I$���l�D�����~�|�M�_|I��jϐ[/�3�Z���{@ }���X ]vMyTJ�&�f*$�L�~ ;���z��Z�
��+u1�����E�V�zh�7'��B�Oǹ�7D�$��'g	]�/��?O ~7�ݛ�a���zX�M@��x/35���3ؾG>��3�B���Q>�#r�4I'�]���)3ګR������}�%���ĒH����I$K�~�\I ^���LLk'�DVB�%e���o��ԧ�iO�C�1�x0` H@!� !UlP��N�X��:���B�ԟ�I ���O�4���?�K����?�2��,�}@3��`i��5���������<�����T�  I��i{���������H @���4	 �%���M�mh�Q�#��������_��on���*��/�_�揸>G�p��I$Ka�����G�z`�{	G�
�}������D���,$�j��'�&���}�A6�����R��"�$�@$����[M�J0�~�ȉ���0g���pl���چ� ���?%��@X�/�]��I$K�}HXd_@��P����|��_Z���K�C�/�-�A�-}a���a#����/��������������5b $��� ��`$R�����H�x�����H�]DtK��J}���?rvR�_�}���~���%��x~��2|�P�I ���/�i3_��C�O�,��64��߭n�A�}B	,Q��$�	/�G��	3��6�����P/���$����Ă�?D=I 	, ��m��.+�L?����$�J!��J� �)`+��\ؚ3Q��`?�@��
�k��\Z�[Y��a��I ��'���p��I N��H�q�&�@>�͇�F����R���Ԃ�����/���ϱC���}��Q�R����O��W���I$�I}��_L��}�$�0o����K�06��ĒH�K��=/���a��a������� T|�����ȘR�t�ޑ_{�|�~��� Z�CC?b��Ϳ��?��~��|`I$�IW���� �_޵�>�|Wݬ�������_[��_����0����~GуH @��L�(?@�>�bA��/��E��|� $��? ��сX?U���e4����:��b_rg��������K+���e5�+?�� ������|���� %]���IJ����3M��Sڇ�a��2f�"F�M0�?H�I�� �$�I��MS&Ѡ��M1S�<��i�d� �� ]H �EQ��������,?M&% ��lJ��,as𝵇$<��)��[|v�ʙNSW����lk�1"Il/��TA��bzaP�S��Z+R�ߣ���W5
?@������O�F�G<Aɖ	��@�B��C(K؍��뭹�g�f�^���Q$�k/Z~GG�x{�M]�lkm���kQ?�9���R�Irg�&#�	��8���>�V��F���i���U�ĺ�%Q:��͵:}1&%2T��/��KbY��U"_5[VbP"<$i7,hy �MjU�*(!���+�����N+��8�
`�dK�L�1f'�b�c�J�Q&���(9��JĽ�g��A'���Z�V�(QA�g �E�

,=��$="��d%T�)a`�i"ڜ[��( qRQ�n�s���ն��A�=�JT����#�pƤDV��Hp��x�$�IHee���U_{����-`�/�	��ܑN$/Hˀ