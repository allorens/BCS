BZh91AY&SY���L�߀py����������`�{׋�  �    (�� ��� 
  ��QI � ����    ۃ�P �=�  V�4}����Gm��v�*"n |�󬔵��[�eB��n�8V��glt�X `������n�ض����u�kH�t
�;�I�{��Dl+Gvu�7n���[[��:�w�  3�W�M��[�����V�]wj3*��7 xa��v���k�iF�q����n�p @&`<�kT�/li�-b��u�`ƇM�K�X��x���k�UB���e:wn�  �c֝N���+v�֜��ٹ�z^����ƂV�a���n�n��� �    (  k�4���k;        WE���U*i��`� 0�HI)U=C#&db ѓ114aH�LA24LО��	�MЍ�Sz�*j�����  `�2 ")QM=5F�h�� �� *��&�R��� �     7A��B�ˉ���.� R9����E4
  �@S��>+UQ9ۀJ����{��^|���)�%0��&�ٶ�2ۨ�u��sns�ʿ���6xѷ���R���ll��^������g��g���ZA̅[���Vga��b���;Tͱ��c�X�S=�p�Y��#��8�gS�\�i���;�R�e1��LO�έ��"0y���{e�kV��9�s�;�\p��mk}6�WP�k/S��Ol��}�n��)���#tb{����V�W'��.O�H���g�6�ۘQ*�
Ŕ'��3D؀ng�-���.��p���\�\����P��\c{hh�n�N-F���V�j�\���Z|(�l���Sk/�V����#e��l3u�-n��,��\��7�RƸCD��ֻX�ǘ��U��K��!��ͽ�l8gy���sS	�0v�y��s���1�j���-���e;(Z7-h�Q8˗Sm���#�Í� ����:q�9�c���z�d�Cs��̈́8���q
��8C�X��kq�۹wm���v8�1��nآ��8ŭ
�nG#�=m�8�s����q�S-�cv8�7����
��>X�7͎`q�5�L8��.�m��8!�v�d8M�B�����_<���7���vk��%���ۅ�F�j-��z6��pC��~�p�h֎plq�Ōq�|���Y�xk�o[��ܦ���5��Ks��8'��	����5��X�G	�o�߱��M�o�e81�;X=-c���)�5�9���b�x�M9�p��W:����W����y���^j�������`�p�o�q��K��8�xC�ޢ�"���P���a7�ƒ��8��e86cf6��Q��!�u���(kF���Z�."�V�ʥl��Mh��C!E��b���W�J�O��S�-j�4�6P�[�wn���YN0�S�p�<soa��PO���G=����`8�}��S�T�[�e�r �*Yn���W[)f�Y�"-�e��x�%�8/� =����n9�kt�E�1��QOľCzC�������d;�+�8و��f��v�[��#7���s��LQ-�bօ����r��q2��-�M�;Y̷�m��"��X�q���V���r���\d�F"Y/P�;�pC����p�h�sV8�i��G�1�>1����山��K��l�[Ѷ��.��ŷR�6&ѭ���x8�o1ŷ�юxk�o[����qNm���ޣ\�r8�pOD
y��#��|<�ŭ�}C�ݶ����mkl�'8|֎:�-��|�#^����~`޲2#�����9�-h\І�o�hM�mknἇ�����qĸ�\���)�����ca�5��-�8�\a.
|�aN).%�cn��N26k�ϑ���p�k�v�k��,[�pH�H�Δ[�v�.G8Ü.bS��qh�p]��E����(�<6�n�!�Cb�qR8�h�b�1�\k�1Ţ� Sm�_��G8p�z��xr�1�(F9F�%ǭ����7��z6��mƣ[e6�����xCB�m8˗��(�*]���ZK����l8�\�qO+�#[y��SP�j\ZۧۉVN8�6��<ϛʯ�|sʹ�^;y���)��V�Hq����8�Z*�n!�W�+'�q�����(��h�+ض�;�q�VtqK���l\6��B�ٍ�Ec��ġG1H�hCX�Μ;���1Ę����p,Z\ELr=��C����TM�B��cx�x���ؤp���-���Z�Inf8�'��ȧ�n}��b�s�s��\b.��ەH�p<q�<�7��k�_}/;�u^:y�۟)��xCz���q�/«b�m
�_��G2G��9J�#i���T�v�|�`�|�m4�؍b9�p�j�)m'
���8]���"U"�#I��h����Nt�Nu�{&ki�j�jӔ&+��&{�	�T�}B+������m&�NP�T��ʅ�MSM���i�h��Z��"SZ�j5�-T*�1ub���(�	��9M�.%��<!��䶚�qjq%��h�-D�kQ����f8��#����l��]8.�J"��o3����V�]��Ǫ���.��y��,D=!��\@c�E[�m�"���G8�Ԇ�O�p�q
q�����r�`�Z�mo��#�O1�(Պe5#lW�ZR|Ct�E�x��groF[��t�^�ޞ��ǭ�KS�J��&+�Zb=�o�'²S��|&.}�;��bt�V��B�P�H��G���
Uj�����'H�oI��z�i��`�+�ԍ?	�%��:OaJ!�z���x�b�,�3�'�)O�11d��lLT.P��1h�Z�H*�J�$L\)���D��.Bt�i�G����w�ٍ7m�Wj)E�NʫZL+C/�א|��MɄ��!����A�]�l�xQ��KZ`���Ub_�_t�1$���ѴeL&���x��ig�M������ߵ�� �'���ؘ9��ޜ��_S��N1q��?���[m���ZcR�Wt��8��hU��8O�����U
�Q��PsD�u��E�������}��ώ���jC������>#�SҊ��#���QHw�M	�Nn���;8�Qg�1s#����H�7E�'����b�5���9�ޮNu�\b����Ӌ;�(�91����GX�L�QG
!y�hj%�8;ǟ�oI��9�[M�5�9����_��s�W������}s���ϋ��}��5��"aq��_ʺ����.���}˾�R�]E��9Ķ�;�,���ҊBr]���>��xｉ�>|:p绛��5�M�nTW��q
��E�/̜ۛs�M�N��;����9�e�a��u�^�������7�=�y��
s�n����m?>�1�:��Ϯ5��/�'�>�ϥ��s�$b[�t��-�>�
'$o�4�{akY�紏��sD�x�Z_�V�h��R�ۧŞC���nz���<�'�;O4U��V�)�G|��(u��q��w��}�{�o9�j|���H��1����ӎ���p����Y֎F{��B�q�#��1���7��7���\(��B��ώf���TFƙ����k��ﻟS��.6\k�}�8i>�M΋vyr�kZ���G�<�9���Y�U�%�d�g�YD�����t�f�	����F�w���T�_�S��t|J��/�p+��ǿm9�'����Ӝ��6o.�{, ���w�����w��#{h��:ZTRO��s$&s砶C�E�C�p���	��^�/_�������Lb��ĸ�5������2#�/���v#\��R��7��)�����7h�͚m6٭ǰ��$9s��gˈ=��HoO�K��o�|o6��4Ν�9�Եě���E�q�n���R�˜#�/����Jo���:v(���oN��7=�K�ѹ���zh��ќ�@��8Y
Qj���{�'Έ�>�+�!��5�&�d��VB��w�F��c��=y�a�wHF�m�߷���$x�D�y(�Ii1� ��N���\��=�>��v��[&-��4�d~���F�!������NR���9�GO�i�8-Ӧ�:Q�.�=4BL�$Bu�w��A����v��Ow9��Vp{S�5b��U���H��t��;g�Q�DWywN����zR}>���!�}�ij����� ��;���[�]о8��r�撈�R�ů�E~W�_ibz�/g{�����CT�e�
�֏z1[�!�}�oWH.Y��MD�}�r��#�}�tur���$�
�hȻh���q��{ƨ;�I{�o�7y�7�Ĺ0L�oh����H?����_!S�����δM���W̵b�w��<n�t��
U��a5�L��c��}.���F��%nb2�WJe���i��6e�9fe��巓�إ���s��U.u���*{[}��4L+DUХ)oc,>{�M�S����/*J�G�W���{[U�3N��s���oi}tЈ��川��F�{*���_g�S�/����f��۰��Zy�}�͝��v�p���v(��y�/w��=��ߕ�w>�_qĻ-����>䨗�����G�'2��5�{�uDGn>��s��/�1x���Kx7D�x���,�ݞ^�?8�mMo��ⵛ��|F���>�996w��-���ˉ��+�⎹k��dm��.�:���v�[�[��D��Iz��b��z*�����N������$^�?y���;~��xC��$��k1��Wusj������{sPB�}=WgD��+ib��nf}8�e�j�%��͏�.M�^KS�Kbݜi�F�b�J��˛�y�j�';�Uw�ONN"<�$�m��|�}�����Է}ש�y:�g��ջ[P�Z۩�#m�4}�s_�;l]k�P�W՜��s�b+wd�m6��֧��r#� �,=��9P���}�����6��I����_Uњ]�q�$NKd��eS��s���u^Ǳ����J��s7Tzm]��9k��������}���Ie4e7��ji�Bx��IA=�3tf���3��"���d��>�M��yܴ����u(�pw�SH>��wy��u�/s5؉߷��*;�4������[���#�z��n�	؉|��>���5����Ӣ����*�!:���i9ӛ�rҒ
���2]8�}j���G��|"f�傔J��%�R��PO\3��!�:��H,H��-m�F�vir����������>�R�j$�붚Х��뻫wK[�rB2A$G��NvC�6>�Yf�V���(Z��?����0���v��wL�ԇ�H��g~�V���S��7��V��D¼{���s�Ss�Su��+鱙91��q����1Ul�\O*�N�9UZj���Ɍ���]�̛jҭ��s�J��<�5�����.��-�-�ʩ�.3QV�H��W��<�/�et�x���Tѧ��>.F��Qy9幷[���p��{���k��o��N��^m�܊]�v�W*�{�v:���I�P]u-5UŎ+gv�����oo{s*��cټ������I�UWW$ۻ[��ys�Uײ����;b�/]����͵�$)�ʮ��D�ڄ�6!t�L;���[=�޽,�C���$;=vj|;�;�zM��.�\��j���=�T�=Ǣ���=�˹�܎��/�����]V��˼����(���H�|i5�u��r��m;�}�Z���(��*�l,[,e���÷�%�����K�<i�#����I7*��$�۩���v��b�����VA>=�, ��8�R�u�k�J*�$��\�o"�6/����bz�?�-��dgS�8�%�S�*��u9�'"n�2�Ӈ�ƞ��[��\hV�X�KR���&ے�VƐ��l��ϥ�I4�!b
.�G����۬sY�"��T���"�;��,����g5��8mݺО���6�p��������V�X�ה�=�ޞWڅ6�+��k�����!�H�����u�jc���!y�B⽜�k�����k��q�{��������)��q�ұe��
ʅfK�/۷9�F�M�[*b��An��o:�8ꚻZ��IF�$%j�Mv������ߊϻ��q��m��ʾN��y#i!���bI��]9~�fq��T�ӎܑ�9"���(��1�������y�Ҵ���N�M��X(77g/�p��q�7�;��������:�&��F�$rI%V��ȅXښ-Z��)ʔL��[Y�����>�;F���N6�G2�F��4�vj"�:�NDҞ�79��cjI�r$��U��Q�"#LU�&��X��ů�}^�i7:��F$(�}h�J��D_w���#�0C���d�']U�/"]k�퐊�؁b�5l���z�w�^�sti4۩��;'kK8Xv�Q; ��^B�:��%�W"��jWeK���M��QkQj�G! �J����W�֔I$6�v�W�ݓ�E�X�}��ѱl��4��26���S���Z�E�To���k��r1�N-i-M�W^�3]����A"�#�5��+��(��J�}���k�d�T��Kb�:�c�V�H�؝�ؕ �U_3��K#Z������l�o� ~�ߑ��*?�U�  �ݜ4�Ki� ̿�/^��y�|�ۏ�����y|�~���P������������~_� �P�  h�  �e  �� 8 �  h@@�  h@@� ����� 4@ `�{��)�+1Y��^���Ͼy�0 ` �� 8@  ��  �   ��HH  0 �
 ���� 0�|�׼m���nY���7&]�3��  p�LL� � �   ��0	  �� � �   �  h� �$C����� �  �=�{�JI����ɥ/ջ���G �  �  h@ X�  � Ѐ   � �
 � �  hB � �  }�=��� H ao��?{���3�� P`@     � �P�8���  � �H X  �
 ,  0�����0�
�^�.�@�( ��� 4@  @�(� h0     �  @ x @� 4@�ܻ�� @`�J�I8�^A9��N�EUH��\?{r���z 5�S�7���s0Pr!A�5]:t��í:�n�뎺�n6�$t�ӧ]G���G[u��z�2㮽u��e:u��GT묺�N��q�:��,X�R�����!r!r,\���u�Tʝ:t��m�[u��u�]e�#�N�:㨧Tˮ�:s�^�c��H]>���+�/8$�l�%v�R�f�a E�6QX8�&Ȋ$C���a�|�͘��"�\c!�4�X�MF�EQ	��kq�R��f�#G�2�F��Rb�f"�ℤU�F�D�(� J� ��@�1�1"2j� ��+;��s�_�#�X���8JA�ecU�+�%!Rb)Q�ǣ��rV!N1��TԠ�O��IYm��M���5dNY$M�7/�9��e\�mej��:�K#�N*Evf���A!ib���2�P�m���4T"ɲ�ˍ	$�m&�,��@�2���i
����y9�����L��_+�����4�UҎ9nXB��t�
X���j�M%L���D��I0i�4F�$LdT�,u�zD��O���(J$�2�)"��]�*�Ӵ���k�m8���x'�����&M��i��X�+ĭU:UnHVʝ��NJ���\��wnG5��OT;��w]�1�ws��_�g�.���kV�ܕc��w{ֵ�r�J��]��Z֭˹*�%ܻ���s���������s��>9�I[UJAE���Z"-W%*������3�v ��S�,�JA)%�$pR�B�*X(�\+��D��+Ȓ��Rq(��i�9�:�p�+�UIB��R+e��ݮ�
,�F���*�ҥ�F�\�'�'�Ǐ���R��TA�&Ƈ�iÀ���kN]�O��6��̚pfp>7'�����˙!A��tI��vb�+MROq�21��$}������"Ե*���J��J���zs&!����X�<9��I�!�p�bvg���厧G���aĮ^	�wy�/1�D�.���q��j��9:h�ƌ�K�YN_t>pْJG�4�?6h�@���G��ŗTK���C�eC%!x�eQ���^�E���V�rm��rO��:�|�=��$�p��*���r�t9�p;��pnB��˺oh4�6���S�rIݼr@�҉Ns����u�tS9n�=M���z�	����>�t�1��p:�s���y�Y�8_���f:BƤŖ��Ta�S#��C8∄�E4ʷ�=����+.Ú̙�$v�"q���8�Qz��XםD�4Q�R���T�7��̑.}.�����򂩂K�y ��kǂ��#4��&.s�I#�+l�cױf��*<���y��GS�lo��h�I "[ecQR�A���6ܵ�X'%�f(e����2i�O3�I"����$h)Ӎ�7��[�ݽk�9Mo��C��[�9ʪ�x��Ұ�pv@���pc�ccBM�昳�s4��?r
>1����dQ8�ҳ�1�S<gL�B���o����#��(���}����Vd�C��^8vJ�Pp��=���4H�����s�wVh4���˞�F0GF&Ē��ܣgi���半��:�,3�p�q$�Ɓ��$>�m�ʺ K��t����1Hta��ld��S�Di�*R�a! v&.��a�a�Ð��1��1���L�W��"�����2C���w�]n�WS��;�nj��|2pt2�J�
��󭁦�qUMU�6*z��܆�$�L=clC�TQM��e�Ywo's=�d0��2�<r���.]�\��Pc�r	���*Q��X%�>}�����i��N=n���s�|�sʾ6��d��K�cq�K,M�:�ý�~!���B�*᝸�f���/< y���A���&yygg���CN��bc�4�鸇�y��斊��4�9FY���ƷaWi�"���\�E�(��E���9ws���g<��'�Np[5�Z�Z,��Z��,�F�-Ƹ�7cR�:�R�pB�OR�eQ�Y����3����&��܄~�̝h	��{a�Bm�a��I,�>*΅��$$�o�����tԪ����8章�a�L��#����$��|=l��ccM�|�eB��I �A%4(�|B�-� ;��5b.-Ϻ,_�����@��7��	�ZR�u�۸�S�:g�e�r��'�W6�xh�Noz�6f0�(��8�C�4=��NI�|d�wGc�7���%�_1���r�w�潏�9RG��ԑ$N�>"�%���Q1�1�D�mJ��Z�--iX�Zm2�-�Z-�KKE���x�iQ)-"Y��-���+ԉ�D����)�>W��>E��"��ZZ:��Q�Zi��E�KR�-��H���Ԫ��h��{S��ҭ:�Z�oڕ\m\O�{S��ҭKN�\uV꯵*�q^"�V�SJ[*���V��K%�rJ�4�Wʕ\z��{J�[*[*�����">'��>S�~H|��KKO�a�y���笼���w��.��罜�4�)��y�vt������|L���Y[�z��͹RLQ9V�;�R-��NΫ�3+�&l�ڎε���Z����<��bܘ+��_/R�?`���z��lh�bI���lCCJ���}�?Q���������>�����`�M���ݒ>^��Կ~���'���w��\߯o�+lK������r���ZĻ����Z��=���K������Z���g)wuw{޵�_�y��]�]���j��Լ�!e���d�-l��,�ߪ�ȑ"D�i�LaC��UUE�i��^���|҆�8 9䏶97��VuNsZ�f����[o�9�[4[�p9�o���=g�ʈ*;aT��n�m�lU˕]�u�����ޏ���χ�Ƴi�!�!�kCS�a
�:@��N?h�bt��.�5|��zon7M3��n����ps�]�F�;��u�m�m|�e���n#��	nV������!�]:t�Ӧ���8��R��6�L����{�I�s���6淍o[M�P|0l{ �@v�:y�bp�F��-qU(�&��i4'3�3���#zh�� t��c�;u��z���zu�5�?�cw7}����ֱ�G�7w�DUn��/��`�f�/���
e�a��8)_8
z�h1Zj���pۿ{�r<����v��m��n��R��.���$����,�D�/?!BY��5�2���2
����C^3�p�f���l�(�ň�hE6B����d�$͓sT�k��8�(�����d��X�CP��Ց�%5'*��R�:���L�%�2d�:T$$$$$�j��$h��}n:�����t��&��Hn�4��L�]̚��n}�.��:\��o��>fGE�;���>�u�{�~�ow_ۛx��4o�m�"Ґ����s��E��Vd���C���R�r���+\�q�O[��[�oK~[�|�&��žﻘ����-i����_����r�M�[�n�֍�No5��}�;6[��7�7�FW�]�Id�髺��Ӳ?!���mX�k��ɹjo?��X(x|JD4<ul ��a��E�C�/���B�����y�w�]����JR����WMֶ�����M�����ۼ|M�o��k�n�T��#���|47֟5%�`�Ɓ����<;sSo�k�Ʒs|��S~�I*�m����[i��!��F������^�\�'�y��������7���w������F�M��[֌�7�o~q�kt�i?�]��{��֛��ܱ����{[�c�o�c���,�8<M9���m�ۈ�Tc���eHʟ��Ye�_<����|��xJR��c�41�EnX?b�C��$��ַ�M�[���m�[�>m�[s����\�ݝY{�N����i�o�������&��������p��컻��By��D(���lul����ַw?n7��sɽ����g����1 e�8�����UT���gq�=�l
��t3�'�T��/��9 ���V���G��������b �<x�!s6���x��+Ȏ����BBBA���~7i����Xъ�W>�YAx]$��J��[m�����%��\y��p�A� ��a���!o�<�|�f�ƥs`�Qv�P�+�4hj��	�]a��
�:8���@<���U-9y�����������szz����1�1�<(˨�*FT��[,����(���m���D���mc)X��6�K+�T��&�V�c�H�B9r�a�K�.����J�V9j$���F�L(������XZ����-q�8K�ែ���_�˟�A����6�S�9�,
i�I8�t@3��H�/��)@�iێ�z@)�N��4�<|J �MFeְ������i�J(��4�4�~,oZ��B�
&�#"5�$�ٹ�����9��]!TJ(�qɏJ-�Q�#*|R��,���*�S>��$��������o#Cƛ2>`��T�k%]Ye�[�xw����{ouUUy69c�<t�u��%1�6���m��s�n��"��E�BLeN���Z�`�1Ǎ����Gf2:^��� D���q��o,۴1A�9��@T౧x���xpˈ�*FT�KuJR��x���,�B�z�"��i�����d�! �`���x~hӬ��w��1U%Q)����c.0]��w��ϸ��#���y���:z�J�qcH�� Gk����6��x������[X�ƴQ��.M��qNr�9�ǡ�7ՎX%��9��z�(ʑ�=)�ԥ2�R���5����������_P�,���rt��㎐�ǎ�.]�`���X�B�q�B����-.Z�1x\ 潋������2��ht6_Z~v=s�@(�,�n�,Fc����=rJ��#���[�t�w2KO�Đ�w"�FXP�x����[����b�Ԑ�FԈ�"'�Ĉ���"Ze)"#�h�n+��8�J�4��m>M'�+�|�x�+E�S�m-�b��2�"�%�E�-�G�z����DqX�RqҖ�Z�q_&>u\G��j�4�O��ǉm)IiɏR%�JZ�i�%�KV�U�U��R�Ե{iV�KZ��J�i�x�Y�je^�U�Qiի�oU�-l��x�ښ]M)l�����K%����&�U�R��U�^Қ]L�l���iȲZZ�ͧ�3��/¢��꺸��8㕓�����sE'�{n��۠��/F\RQ�����gR�i��^��C.��2��SIӄ��1n<�R�;���g3L��7�4�c7��ޱ��b��lb��M�Ag=	�c���p[E���K4�m̡n\Ak�ĪGӝ�NaQ��DcT�8�.#O�ۛ��ү3�����ԂZX"0��HP�(���)�9nL���(��4ݩ2D��k��E�9/��#:�c�;���&ӥzn{	�����v��]�ĕq)>�r�̕¡�N��>���w���5��:�����=�]������"w��RV9�eOe�v�8���5��"�k����_x�	�������#�o�ɭ(��1$%�m��s8,��4�k4��[d�ʔC��R�P��+�?
��*�]W���e�F�k�����:��w'�gד�7l7���v=O�|t]|�Ɉv�GP�mq�%F�٫t[�r84������X���ȔnG2:II9]����Ȑ�VҗY��dUr�XĖ%��n�,J"��MIkRB�̵�능!eU7c�N�)Hc�"+{r��`�U
��l��%JEV,lqR)�p��4���bJ�X��b�Ǔ�l湻���q���+Ğ��w{���_n�^%�n�w���Z�u*���z��ʯ����������3.�_C����O�nfov����Z(ʙE,�֥)�]^tt�
[DG
� B��NT���s��\k�ByW�n��2��d����b�	T�E��%ZQ�Z�\�S.�ն7%�V��H��#@�e$.sٞ��zq�+j�9���O��5����� CQ���!�ϵ��gc�#���j��`��Yt>l��y����{>Y��[��7���q)��9���=��VV��<i�@<�7:���>��C��d�Xah���ؾt��\�87��w����fT��6��ݴS��2ʔٗ�)���J}�{�~��쏎������e�p4hv�eS�F��C�͢|�����wzs��|n���W������@o�3Ɯ��[C�H�p@ûdTj 柇 ��n/�9H�y��&^�,��28��>��䐪�c]0Yd���a����խm�B�sM��ʯ�����7^�P�e�����1��u�!��Fk� �a�*/8�O�t���P�1�I$R��S&��x�{�c���>nۜ�WǾ�29:�pqᶏJ��T�F��1��9%�v���;k�%���������9���:�  �����Çļ����\�0��@��܌�ӯ��8�膀�R�ch���ɠ>7�5�3tw�!f�"��*SF\|�)��_V~��$.���m��6 �޻>�x�J�B��{'�<V!/KK��Ź��F��<g�{�����s�<[N���m������ї>����0�`�h��c�t�m�OڒM8r^�ۇE��-���Z�ÏX���i�E�T��[�)L�$���:z�k!EF�֠�q�MZ�A,9�ɲM�(�3��L�T�pC��V8�CdD��(�-�p��dW \Vrۂ#Ȋ�UA��m�#u��ױ"���T�VHHKs�-֓<JS���^13p��=WSԖ&11��|�EPJ�:��Ç8~��KSM$�0��ړ��//%jdi����
���u���t~�<:lp7��}uUD���}�*�|�[�|���n�u�W����ҕ�BD�m�ln��xu���cB-iJ��ex#��E4cn_~���4N��X�䓃�`�Xߌ���?�`�A��C�!��jGӸ1VtA���5�o0���b�&Yn[��D���	�^o���{���}�������á�͌2L���ٔr�C� 9}�����̉S$�UFi��0;zp����Q�I&��
n�2��;��Hmر��>f��F/9"�^d2�2e�  ��`�A��CD#�>��6�S�eZ�~�������t�>�=틠`�=�r%�#��u��$���pd�4�Ѧ��m�ٗ.��@{'�&pM6�_"�["��g��L��l	�%�~N���n�t�N�lywE��Gϝ�oӓ��U26�9�}`��lb�k�7���j���n"��*R̺B,׉M
��Q�N�j0�L�e����ο9:��[dp�b�"�ʷ]���z�~s�y[x;_�]Bi� ��fئ~ۗm5�?9��3c����Ð(��-�\���c6�BG��@�C���֞>s$8;ݚ�24l�^4PPp���΄<!�W��X��Ar�7t�	FHX2̅�cp���ɒҪ���cf���L��8�7�ծF��E���"YYciS�� Bkj����D�\ѱ�N��d���N�	�����&�xH�$"�D�~����x&4�����;�c��/�HH`1�޹y̥�ݡ$����350ݎ��� P�wxgL��9c�^��f�mp:=�"��������e�`i�~4�dhjڏ�#(��Ӈԫ'�?6��%�삪$�8����c��0��p��S*G�[D|�A�u���j���cf��L�r�{��L�v�������p����N\�t�����ʓ��`xy1��MJ ���|u��f�1�X�������6>Ư!Bu�aFZy@U�������q�U��e_oe�fqۑ�`L��ėkK�I�OJ^$�R-�Rc�h�i�R�Z�h�i<KM��m�ͧ��>x��>U'Q���">H���%�KB��Dz�'����+R�E����iiԷ�e�uV���OV��;~��K�>��)~N���m�6���-�[ړ�n�өn��u<��x�qV���n�өh��Է���yR��im3i���D�YE���U�ۊ���<W���H��^R�Y,�%�KZ�j����Ջe�=s5�U#�Vi�g)��9o9 տԺ.�]o��94��p�w�vi8�P/�{�+�*�Ŏo�|�Wwe#ΦΕ�U��Nif�Knk�(���SKYN�dw��z՗S���-I���rt�y$Tj�6��M��!�~��>k�K-ǋ�yu�|^Nko3�&�'��nf]���>�����O�nf]�����}����f_�ﾈ����}_nfe��ꫲ���|��<ݮ.��W�y盵ܺ������eh��l��7(*��2	�ӷ͏��\��n��X(�<QU	R�o6�7{���w~����{o��ƀ�`<�it�{wn۴ݙ�?�%��.��*��n��&F����6UU� �G-���S�������y��c>��d�O�DR2�#/���~&�J�@�kS�:s?w�)��|\�5.�Cφ�к�|脝ȳq�̹ �w,Hx�<���F�9	HPu�:�ěY���g3䒡��h<f��ϊ�����1�=�u���.�:0��Nw��O��%�m� �@Gu�� \*{&��m�UUttˡ��ӠS1�+�!�DR2��2��	F�?On�3���sq��A� ��7aJ8rnD��sM�#|�)�ú��set���R�ERk"łw�p*Ȳ��h�ˑ��q�Yr�IF���*���_��ʬ6�(�Ti�P)�c�c��������a']�G\`�`L����G�;R5��UJ�|���A��fI*����2ӗ@X��;�q�c �����!.���L(P�<�����y�r5PQ���to|g�\C�~�:�	��O	a�L���e�F^":�0T�"5���@�q�	�ó�������di;⊒5:��=-N6�20�,=J:��.@�Zb�Z~C�������?�.��r�(�$M9	hE}�������9���I�O�E�ԗ|w� �i�M�&��[kݪ���ӥ���Q��#/���e^Y�����c�G�G���l��Y��ƀ����2şm��Q7����g��>^�2I��<�5n�0�+ރg��(,�ƒ�pI�� �L�y�F ͏��0�#@G��]:�v�=L�J���-��,���# �\�C�JV��ۗ�u���G�"���e�"���wK�����Z��g��uۗ5˕�nР1rN v;�m�`QJ`�?�d���J,�n+RI&�}�ϳ��*��r�`Jc�`���K��[t�XS�u>����ލ�Ƴ���y�I:\�Zs�]�4[s}g}��j�ۡɱ��zP�rj�!DR<i�Q��V���m�[������TT��27�4A2�5KM�ڊ�j��G�"�k�Z�o���Ħk��dq$Z�m�D�$J�Θ�i�<��CX�Q���G��� K���3 ��
��m�����E�9�nοj����7����I�.G��d�^����8L?�������l��lx>2��m�0<S\h����y��<o���}�޿|��Rz�m�֯yR㜹�q���t�r��������tޝ=f��B��h�1���skaG�( �R�D8!7��#�����Io/s���^���������և�R��r�u��M7��5U~|W�{�������$�8�q\��7{��~Ǯ�IT8�ǃ� lt���u�����a9q�O�x�6��	��,���坨]SU����i��V��������z�ϻ��+�s�������c�(�)i�<\���@�i��G���E����ϛ��?onϺ�76O���7{�$1�K��FKU���Ik��j����9�u8l��ܹ�>y�@?{���-��:IWWtU���S�4��1K��bI<A���'g��ߞh�ۑ��ɒ���"��������>x�"��L��)���{ZLV�%ݕ��6	����<c��ʦR���`�|$3H5�%����+�I��I���ym�84�` �i�6e
f�[���Qs��-�*��c���m�{c���L�@��0l{J� m��g�Փ̱�e�����.G�쳸.�^8����������%�DZDƟ*%�"Z#�̘�*��i6���Ջr���i�f��GSiKR%�|��|�>N)_!�x��U}�_W9O�9�o˴�-7%�n*�$�-ږ�Qǋ̞"�RD��x�x��-1h���v�'�T��^��|�V�N*өrv���U7R��[�[ږ��Y�:�N�N��S�W�Z�M-ZKJL��*%�ȲY-�8Ҹ�q]z�y&��ij�Ze���K"�d��������V>D�"{RW�Q��{7Y`Q!�5�8���F��ED9Ch�q�hѐv�c�elTR�&�q�y�A�ǐ"(�U���v�z��±S�ϓ���ڷ��*�}q���j���ݳ�o.$qԅ��`��vZ�!��R��Q�^t�j�z�<r���F�lC)���:u��n��H�(�ɴ�H&#j!�������3���z-�2pu���v�ьG�7*���7th��ݍ=�v&DZ-q�r
�T���7��61D����2.{���k�˩�zn�G̢{��mһ�%�|�����,��X�qAEQkv���>�<���q�mS���u6���[��P\��d�!���X��/'�ݧJ�L���+ﴺ��"����q��]��K����������:��s�?.�NU­�}מ'�=q�pg	��3�u=m�;maRh��)�(���*,�B܎F�j��Եb>�4�D=w,MW�,,��]N���MK�l�1�����jb�6��T���D�"��]r)�$DuZ�)b��*71�V#�^[�9�4VԂ�MTzKP�ě��u��c��N�L������?����������}��?�����̿��?���������}��?���{�y����]���|��<�ܺ������Y�V�)mc��Vi�2�m��,��j6 �d��"c�l�HDH��`Q�KF���B+�2�c�Hv�&!�I ��+�Ƙ�m+QYr�"&��`�RѩC�m�0�M�ٸQ��U���-Wǔ��%]�i���bImj�v�|l�W���ʫ��"a���y˓t�>w�9�+.�ƀ�P��5!8���ӆ���C�0sl�*��%X�rP���\�L�`w릟��a�TѭSl�"�0nV�m	x��3��U�X*06l~ry��b�1��f��]�!��R1��������'*ߣ�}3�|no7��l���[t�|;�fs��VU�R����
m�cׯ��N8r��t# )���~]#���1g�fj�<	��I+�P���:Z��L7����ӆP��zn��UK;o;�~|�����};|0c��:1��i��G�����U�lC����z<3-�6�ɦ�lk����|�v9#�烌�j�H�<v��ǚᝦ~�=�эd=I�&Ց�U0#d��,Ŕ�٠��g��#�Нl�֞����W�c���q�1ɑ��Cj[N2466�B��r$ĕ�����H!	Z���zۖ�5��h�
iE)��R�<q�"�:��ǀ�ih����3߳�� �r	GqLD#�V���7����wn�Ҕ��x�[�9r�9Z`e���:�;׸b�%T;5��0���m-�Zr�:�!�c����~�M�t9h0��>|dy���Q�3�����h;�L�"�����\g4��A�1��	�l�r�)�8�ۑ6��<b�J�F�ȄɲY���R��*��J�m0v:����E�ll��*8B��ZM5VHd�d�Ĉ|*|.ƃ�tX�Ӭ���BOS#�ǈLpx:L�^G<�v�_�{4�G�V2�c��B\��썏��3��a}���+Rېi6���K]e!a�?���?x��c0=�8��9-O�\�n�5�����W���ǆθ����)�jR�2�n	�4�ۗ�dp*��L�5Ib�p���C���?7�$&4�.��a�4/.B�q��Ps[
�0�ܣːαTf?���U�׆8�*�c�}���?g�S<c����X�&B�d���-�S��g��5��h�=QJG�!�h�3�������q$ӌDت�68��q�nl��Np|<L?ez�z;�i���G�Kbe(7���*�"���]���R��M�NߴPSC͎��k�j�XϮ����~n���ּ۳�wV������9�c�������f�ž�>��<��TL{z���DS��c>${�\7�ޫ�yy5ˉd��v�4�%�x9l>64d��h�<�1�� S�9�R2
�%�՘�Ky�����G)||3!����Ǳ�w��=$I�n=�dw�=�C��4���2����h��)L[c�yϨ�أ�l��#��|ڔ��kh��Mg=�нS��h��e����4�MHR���.&�&+otee�]����樅����5 �Gɺ�]o�K
s�}�J�B�����a^Y�D�텄�847R� Oh�"q�5,��#[i�?����<a���ch��� H��c��Xxq>��OCC����Q��Sn�j�{��e���\��/��5${���2�;��pdx01�C�QL���%ʹHI8����rH��Ι���~��!S����o�_����3�����Î'i8���O�����r�rۓ�NZ�@��`ɱKp�y���,�x�'�)ϭ�y��c���E-��Cٗ(m��������Ur=8�n1�~��!kQ�Z��Mnp�3�=;=e6^ݹ1(0��4�a!	�	hg:�u��>�H]U�v��z9�N�K�Kx������D���">DE�U%�%��l�h�i6���KG���TZ�Lq-6�Z�-"Z"-"ZD�q'���z���%=S�+�|�'��6�-8ꖘ��Ke�q-<OY[8�i�i�"��M��V�V�]In-�v�Un�i�4��7S�[�%��Od�[���Դ��ԷU�z�q>r���i>L���Ze�1>%�K#��*x�⸵x�yRij�Ze�^��-Q,��,�ZRu----4�)Y�o<�l��u"���<҃�rsdg����BvG��z6Y~R��]:_wO%����{Թi1�b��*Dn�4���w"uɖ�	2`�8S���bm�ҏ����\�LX�ʻ���o�f o"��	�Mp�JZ��.�9U0��������w%�.������<�ܖ任����<��r[�www��y��%�����y疻��.������<�ܗ�!kQJE�)h����x���l%&$S��q�$���3�#o����[��$1���(f��;�1�B`���#1J���zom�����}o��W����EW�	n"u��	��ް�I�����2B�Z�N�����R8��Qx_�I��3�n翜W~�m[.z�����{���@TӇOb�0%Jx>�9>Ĵ�Y	+�U�m[*��X�f.�>n{�����!��h�1��Č%�|��c��,7P!�C����~|� w��p���eK��v|<\�F�T�hpi�kY$���|d������"��W�zԙBiD
,�z�B�LE*n	��o!�J\nڶh����%�s����G�
�C�IqC�����I�U�cw�]�(��<yPԷ����o4`��V�$ʚDbLV˕f�,�|��+�w��[�7�r?�������ˍ𷭔�B������]li�h;
�v��d��n}�b����|#�AƓ�<p�7O_���^�>�::�%UX|4���DS�G�V3���5��c@�!!	�LA�7W{;���&�]�uW�m4P����6�HH^D�4�������J��$�M\�&)��ޘF���m�o�*���C!�w�c%Qp�oX�G^�!a����	����F ���a�C:t�M�LF�d24`�"�C8B4o^7��q
���|Ͷk��I^���	��C���0�!�[$}��~����e�i�f)�*�dn��ǚ,�
������ITa��>��m�/����a
zu$˶8�F�'[����o�2���1�<2�uDS�G�[ٌy6��Xr��wǰ�����9ij�Qj��sR��Sӭ��>|ںQ$B6ܭ�x�!h�E�q��tx�|06�H�y��t�8>>���07�wtgYӠ�P���X�m�n �x�؄3D#���壍u��дN��"!��r!	$/�-����[������b�z���d�-�".˺�Yˢ�,�ga�T�4;=7��F�s%(�me�*XҎ�cK����%���I��9��h��ڊ �b*��γ��k��\:�dv��4����Ga�����<;}�ĜĪ�=��d2�c��`,!�o����<|9���	V[uP�I"#�� �*gs4�u�O�Ϙ��ʪ����|��ȏW��j��Hx{c�-�G�I5*Qf��2!.�㫼�$��08܄��)��cၭ�I6��t��x���������렺�v'i�]�/7����?`�1���졆1�{�N����3t�W�`klL�CF����E=Dw(�������<s	���G����y�p�����syWZ��xr^�����'҂�
���R%���
2�����3�M�n�]�\4��T�靧�|o���2���S߸&G;��4�-��mDS�GR���9\���n��K!�ˌǟ�
t���$�ɉ�~~49�S��ţ�U��BSdH���ZV�b��hA�����2Iʪ��_�S�5l!c�䕑��8|65E�i�,m�h/-?��ᰐ��޷g-�~����zo{Δ�.�q��I�DqH�DO�"�TLY$�Z"Z#�Z-J��m6�KF֥��Z-:Z�Gi��������-$��x�	�z���}Z_WK�?'�������KN:���թ�q8�x���'d�D�"e"ZI-E��+W�xͣ��-�{R��6�ɧ��*ܩ-�[ږ���M:�N�]Ku\OSķ�&��%�R�R���O��N'Wީū��ʓKV��)l�L��K#�ʉ��J�W��>O�n��Tr$S���P�Zį��-i���������?imnA��83wr�e��|0k����Y��=e5������ק��+�-W�H�e�h�VE�f��f�ѱ��G�u���-�a:q�;R+ތ�Q�s8&#D��ӚD!�N���C�:r�m���чz�7�j�)9�F�ϸ_��<5��qeț9�H�*C�_h��w9�;K�1�I��m�k���\zyh-��8T�Ϻjs�%�9��C���=�|���xU(�v���C�����<��tߜ��f��ֽ��9y=Z�.�ёu�95)��+����y}ќs9(�R��Uլ��"pJQ�vD��f��b�rW%J�m�;8��jH�#+����]�o��ϔ���Z��"�׺��ma;ޯO䈓�v��^��q9�mQ5��YT�\��ߵ��NkՑh��Զ%mߝ��{��]o$U�&���5�����b{�{�Zu�k$��X��#cE����C�6����?1۵\��S,PN6�ʙSCd��;iM�S��qS	�;tگ�믶��s|��������s>_|��������s>_|����ﾪ��ݮ�O%���Zכ��%���Zכ�]ɱe��DR���|���tz{�T(����,P ��&Q1�e)JB3%�whY�b#!2Ŗ:� ��m�S�1�dd�l�j�J�B�Aإ#���"�2kn�;���JO�6��H�5�e-2��uV��qp |z�b�eY[�s���K�񪪦���t���u3�%�7E�����2�i�����9;�m���}),�f�$�(�M�d?�D[S���X�$Yޣ�����=�U��s�HI�� �Z�qN�9��j�ܧ�i�V�a�QsYƧ@>7H��Z$㒾(<�TG��g�z���D�������464{cB|�~�du�;2tft��!��YU�Kd�����\����j�}�u��-6�oF4p����0rI!�����(5��T���Q�#��E8��}�QTQ\ �Ɲ�6�衷����d Rp��`���a�����&�}&�l����SG�-M�������&�/��۟����.	�|7�"a�����z4�t�OoN�o��=>��8���r"������Y�`�"9li~f�����8ɽU�E�I%�m���r�����.)���B�J�����=	;!T[���n�iрFVk��]�=��W9\�zߛ�{}�2d��&Gnh�B���>}��xm��QU168��%����Đ�1���i��JS�W�V}�q�j�(�"�F6Z��(\M!�XJ�	Q��h�qFD��R[���%���.�jM�&�:�rB��-Q�X�5s�or,�OK%y"��h�#]�i@�UW�̇��i��e7v�N�fǉAe�og'ꨪ<��_R�rNU�	2h����ڪ�yrĆ�x;��J�k��$v��x5����7G�<=3�t��ml�w}�+b�b*�ĹZIT�ᛁ��T}�<�q��Uz�b����|�)l֔@�Q6�f,Fq�CQ��y*m��t�!����!F�$�Άu|��M�`��b`hqRv����o�e>(�GNG���%������V�j�h��4ɊO�w9�w�̎���y̡��z~tt���K5Ǝr,�x���� CD�h��4Us�#d���O��fz/^4io��W�v�y�o��>?e<q�^�x���4���4Y�d2\��Pc��
c�QE��M�"U�,��j�ec\�Y�<<Ǟ))����q���Iup�n�~��4�h|�1V>l��:�Y���!�>R��\*c1����mX�l[t6��n�Yz)�c.�N��0xh$ b6�ĵ�I9�NL�G�J3GoF�D�Z4��n�0��U���"`,`m���;S�A�����:1�h6�2P��U5E�Z�[�P��#�=S�)N����!>ؔ˴X�շѓ��a���(!���Bq��I�����'ZW���׈�YP��uL�n�+Q�����h�M��-��Pԕ~3��yT���(YmR�r��2��E	��6q�jxt�af�Dz�m���,z>�Q���7q�z�d�����������I1h�ڢ���I1#4�U19��N�~o��;��≡h<@�(�Ep����.� Ǝ�mhhz7O�x�� ⨾`�����c�8��SN�e��rFt~��������7Gԟ�Ⱥ�j��.s�ݴbC^������3UwvJ�f��<~��k�9t1�Ii-)�)te6�:Q�êGŝ:u�
P�4*B	�\'�V�)�!!J:t�Op��m-��������z۬��N�h�N��,B�!j��B�)R�Z�hB.��]z��\z��m��u�T��:t�x񧎸㭽m�YuI�!RhHHBhX�B�D�j��,{7�b����)��s�7�����sQ3S*25f�^�d���*�&�Y�O�w�3�v�Ʒ��iW���ډ���˾�����佥~���a�~4e���W�L�gw����b���%��?)ƕ*/�����ٛ��j�J�[�&����k��Wr_�����k^]��ծ��Zֵ���MZ����k^]��ծ��Zֵ���MZ����k^]�����"е-J(�W�-��C�����pW����COZ�}�C��-.fh� Յ���,,����O��F>�/Cxt,��j��S�.Zxp�C��trw�~ל����{�nw�J�/�[����;�7��ӌl�á٦`lr8hˇ�ؤG�FQ�-JR��Y�a����WUO!E0Ԅ�A��g��!�F$s(L��L���Ϲ��4ۑCP�_8��)�"�`��s��<m�8�!l���,(0p�ގ�5�d=(��l�<9�s��GX�<p��_��a��?���o{��}�{d��N�N�|1���x��9�AI���(wJJ5�!	�$�F�2ݎ������Q�*iJTV��h�9�҅�!H2�(��J����+I"2eyT���Bx2ü!�ɚ�$vǎJ�h�ӫT8�����`�)��U9��� �laʒK�5�P��ӸƸϼ���c�0vfrxm�$$<�8��f����aï,���BFМuc���}����U��ߛ�q'�N�O�c���ϖ)!�U�D�b��1�vT���'����*�0p��R_C�hp�`��c��z�;�X�}�f�_�-�8ѓNov\�ou��]oh�M��3�}��e��i�P�e��ڳN���C$Y$��ێ8�v�}���s�o7j��tg��C���}���Ǭm�m4lmK2:�����H���)�.�6�&�K?c�����T���c��b�̹1�/���(x��m��3Ñ�k��Ud�k��Ƈ$!�4B�4c���E��t�i�ͶscOу��	<4��)������ɑ&�\R4��hH��SF��,�1<x�Ӯ���ӧ.X.�O8z�OG����8�'�Tq�1�e��Dۦ;���L�{		ht;y��h���6:��C�P�h�Bњ1���y��),�aE�ۦ��JԱi ���x�T2icp��H!��Q�g&mm��#�HT��e�5d����ԣ�V�� �6�DBuYRlm�B{-Bq�A
�-�&2��p�憺F��ȫ���*X�b�	dt?m��&�f��|�Y��#�U
�ǻl�A��c�=gM��	ƛ}��ӳ�oĢ���UW��x<�>����r�B�0z�9V�.�ǫ��{w���3�ַUoɈ�V1�>Q�#�|�)뚽K�x�b�89t>�FGC��W9$�M��3���LF�˩!���>�4ۓI�[�?g���ί�sswۏ\������Y#�$��O�����첨~G��w��.���1��	�-��\駉�Oڐ�_1�Ǟ����_���{�w�Q�I�	�B�f�c:u��mV��YP�_�<�MY�zT��ԫ����뢷�ꢥKz���v5��;�
/ti�s��㳖���Dn����+���Mۯ�<��eyfI	'9K��/ [�r�w�2�h8��(��#�uJS��&9�c:�_Ͷ�!��C1��_`�� ptQW`I%QEևf�h~/[��8����=n=-�Z9N�Y�8�s�{���X�S8e2��3�NV�i��&��$�ղ3\xn�����A�����˥�Ykx���Ɏ�뮸뮺�uH�ӧN�����E��N-���u�[u�qӥ:�u�u�]u�[u�)�]z�6�m��:��^��׮�u�\F�m�YuH�ӧN�m�ۯ���[e�]R:BT���	�ԡB���䡪U3Jq%�E�8:鵨�#���4I��IC��J��,:Wl���"�z�^/x�4�Â�Rl�7X�8!����Z�"T��Є����"��m�l8FiNw���΋[��c_kai�J�ɞ\���˷��[E��I�����_6q?<�s��A��\�Sf�b5G�I��r��,�Wh��;����1b��΃���s��GwԈ��d���E�ts~����m9XD�&��i�j(���'��9��Q����q.r���o��I��y�8��]6ZM�+ZH��w�����$��:ڂ�J���o��=�'a�?�w4o>�s�ۿD��������>����DO�������atz�V��
�l��6>I��C�$�+���3%G�����m���Ż�֔v5#�ݨkSܩ���D{�˺����;t^��;���/�s}w��G�U(��)�X�J���$��\\�ݷZ��D��m$1��+Gdb�z�J��J��E�cTm�UU�B��e�H�Sź�"q��ɍ�5%�:���S�d�9UQ�n*�RF�%�����4�D��LT�Q�NJ�F���R�Q��c�V����{�ֵ�>��I�]�޵�k˵ܚ����Zּ�]ɫ]�޵�j�k�3k��ֵ�_-w&mwwzֵ����h��h��?c?����,�e�W����# �B��(�Ѧ��\��y�=+�6,Dcc�&�3^͔E�DћRM%Q.k�lBb��>�1b$Ԙ���*/R��\��X���r~^���ˆ?=)}�=+7�����GF䱏!��pp}�:��O���ٸ��f}��<2�H�T��6I��Yq�}��gLYfL��[�Gb�ڔS(��N�Jxa�]`�UP�i�:����:r���a��u�t�_8��TmԒL�N<p��V�@�WM�v]��O�������UJ����oC�-���,!0PUM6W�p�/d����8���T�8�;UTȵ
��ӌ���$��!�����	���*[�Li����}��{�^�<�%qU�+�G62�&���$���}ܕ*�)��$��$�ϼ��NS��*�*���K�˱���_>�M����pBFxc��")b��Ճ�`�v��tr젬�HInM<%)�+�M��HԊ�JҘ�3�u�?9hp�w&4����e�x�}�7�y2���ǃ�X��^��.Gy�����]8�יc5&$;.v��9�xF�E=DGh�3��?!5[q�QN|(��i�)���E,+#Jd��dY�9a?!��E|j5�v%RF*�Ѝu%M�QA&I�K*���r(,CmQ��J�Z2Ga�n�]�,bb�O��tC�4�X�D���QJ�N&$&�B�р���#� �s�)�c��A�N��n&��)����T���LL�,z<)�Ia�|!*�$��X�g1�љ����R�S�Y��x�E��LwZ�><m�g|9/��2��|��)ꔧ�S���"�J^k�C��3�<���w+�jBy���T�@9Ѯ�^�^=�JeU9��$������>��Ōĵ�"m)1�'�/�s7/|dJ�9*i��I-��c��E��cX��S(��R��ZD�uqj�_�����ZRM���!� e��ՕWsNô��i���u�DXX�-�XHmj+����C��q2>hv����4Ѽ>_����=�z�����ԥ-7۽�11��X*����{�:�,:��6�!�땛��~���ԟ�&Gc��Zp�lS���Bh�~,(���BĔ%�z`t>��2h�$�!D/#~|Sno�Jý�N�k�1�g#���vn���'�r���M鿺n8�����޷�xeE�"=S�)N.k�{�2�,���K�i�E�sH���]�R�b��eKh�MAe��Sr��LUYLR���D���q����\�S$&H(�ur�{��_��u���NoM����q���@�i��*�Up`����|�u�j���S�Jz�h���އ:Ԣ�Cc\HA�
s������Hli	���4?���b�ӭ��hPc��Rԥ<{u��53��J�Y�b�2;L;W�lv���n���'�[���"gǝ1��D:������t�x,g����ԝ��'��{<eo�������r�{o�v�ZJ֤�|rMk)K}��]�|�����dv�9�p p���c��x)�Ν:�:�]F��u�V���-H��,�������ũkj�޷il��^��n����C�u�u�]u�[u�)�]z,V�R��Z���\��\��ۭ��*u�t�ӧQ��m׏��h˪uH�Ӧ�:�:�.�R�/��R�uV�7�f�_]�&�����zޜ��X�^x��|��h�دʻ�_Y�d>̥�T�~~�h�}x��ˋ�X��l��3qYI���]��\}�2�T�T��ݛ}���¾>�ҟT����=Ի,g�>�=�n��{S�ծ��Zֵ|���Z����kW˩kծ��Zֵ|���]˻��Z���Z�w.���kW˩k�e�����Rԥ4�롪�Xr5�2�U'�M0l�I#�$&s��{ٸ�>~��Y%��=���9bdqC��䦪���¸8C�;�H@�$2=7Dm��~~�b@�AAE��8QҊ(铞�j�]I_U���z�Zy)��Y��C�cjox*��뎮��s�.r�������o><=��t������8|;�C��F4d0|93���q��r�F4��U}EV��+��o^N�������BFtc�}K�tp�L@�n���JW�R��Z2i0j6Ь�,��B��.2�亓ت%��|���ճ�%j��e�bIf�i�%G^u�^-4U%D8�Ij�ĕ�r42<IU'���)�k��,�bn� r�#��#�pnu����Y8���� ����c�2X�����ގ���HY�0����,��vU,b�x�KE$D1c��Aы��̓%�(��DF��)Gsf*�{�%�2�r8���q��1�7��� �L��M0|=�M�(���6m�'ǉX�C��W��	_��6��]�ι����c�wo6FB�N�2?8�\����&G���P�>�����s�i�F0FGn�x���d!l��:�a}��D�1:,��0:=��=�y�����V\�L\雟��Y�� �m�edB-i9P�mD��Q$�&c�߄w1�t����{��0��-ہ��Yx��u�o�\
g��FQ.���g	�1L<8��m�jR��u�dֱrL&6�%������z��	P�!>+l�K�[8��`}���o^0~��??4q�����ӏ,�}��~05]��Q�Ӿ@�)%� �Ó�3�2A��Q�a'a0e��A�*(���6�)޼y#��V���7&�VTd*9¾P�����nѤ�Ֆ�t�*ĔtԦ(�I���ŕ��jbN;�e浚#�<!�ESV��Yr]�MC��n� �	�9���a�3n��;s�%�D�sc�ç�g^�����9	8�Ӑ�:UVn=�sK���S:�rₕ�c%HQ�5uC�ec�r����t2P0d�hφ1��j�]!�p�pm铙s$#��Ɏ�W��������}���ДBN�l
0>l��P�11��M��B2"	��~Wq_}�?�����cIۼa��_.��돥�z��vs-ƔQM"#JZ����������+f���m����[��M���Q��x<I&�6=r1x7�s9�D9 �)�۫I5�&ޤ�^�gXSD�Thvu��ۦ��{�n���!�C��_��Lf��F_��t�ǬM6Q�S�Dx��+���T��J��o�Bm�$!���������L�VL��v��﫝rt�r^_[�7������ܲ�����ܓ��!��%���=�M�09l|}ꪢ��0�Zv�C��U��YR��Nuh�_��?})�,��UUJ�Y��f\O�z_J���4	<��[X��DU]��D�
������-�	�d��H|���w�#,4d223FA�,ddb2�h�i�c�ۆi�����mfɵ�#L�[;���fBfC�p΍��жd-�cB�	�u��5����f��!lhY�!lh[l�m��gЙ��B6аB�hL��k��q�Ƈ��hP�&�Bд8��B!4(ZBК��Bд-B�P��uhZ�BhD&��5���B1*�b	�& ��!�su��}�$��g4&��С4-B!4m�B�(Z�	�4m4?���4-�4-	�BhQ��hZ��ZBКF�Bh[Mi��&��4mhF��4-BК�ѵ�2�д&��hM	�hд-�&��4-F�BhZBhMBhZF�!hZBЍ	�hML����д-BhZBд-F��4-BК�дmhL���BК�ѵ�4&�д&��4,BѴ�X�К�д-Fօ�4-B�i��L֚�i��i��kM4֚��4,Bд&��ZBбL�hZ�КBhX���КBhZ�К!�|�BhMBhZBК1hD"BhMBi���f�֚i�4MX���Mi�4�Mi����DM��дZ-E�Z(i��-EEB�dZ$MQ��ȴZ$MQF�D��6��h�Mh�X���MD�dMc�rk��D"h�D�B&����D"h��E�4A#�!#�!4M��,D�"h�M��hhDh�4B&�E�4mD��D�4H�(ډ�4&�D"hi��[D"h���8B#�A�!��!&�D�"hi��D"h�,����c�E��!D��!h�[D"h�MD"hk"h�D�4��IbSe)4�i4�ZD���I�id����&��K%�$�4�l��BM,�K$��l�t��i4��BZY#M��I�$�	4�l�ZBY��S6�2ͣ&4d�h�fі6��m6�4�FX��2m�d�h�m�e�h�m�&dd�hɛFM��L�ƌ�de�6h�lFY��afBE� }����5���攥4�[�;�k�X�6�3mJ�d���p��}n�k�0�a�W�d�g�p�K�����nn��?b��������_q��Zp���iY=�W:_������4.���63�<�A��|/��������3Q�EU�n=�[_�G��A��	�D�H���� �?)�Ec@���h���s���� {V%.1[ ~#_�V���k��~d:J!�ӵ�� �2=�*����~���-�:]B���m;�-b��`�M9��7�II����t���8a�n18)�w�|-�Ǌ�^�F�i# ���nV�8��(R�GPDl
@���|0P["��� D�ء-3� ��5u6���<��^� #�?�r?��E� ��1BF7�6�qL��BM�	0�Fٮ�����j Dz8�kX������C�!��� Dn2z��i4��R�tO����ć� Dg����v�����UQ,����_�N�?����.��}<����b!�Vb<������9?�^�Z��`�>�D�3��umw�ں�q��y��EUr�AH��}�#��Ww#�3����B��`��3��"����+�;K�LO5@u��pCS6�&����7N�������6{���IK���ދ<ׄtRΐAQ� 1,\h�"PǛI����C��M+��˴M��=]<�����L��k����a c
0ً�D�'�~�j3��hqUD������g�1w �j���}W6��4,?e%pX���j��N���<����ҐS�(�#����D�7"��m(C�lT�@���C����ڊ(�����ի+P��M[+VVV���+V��ԭYZ���VV�YZ���VV�SQZ�Z�V�5eej+(����)���+)�����+(��2�+eb��
ee
j(VQB�555e5
j�+jj
e5�ej���jՕ�SVԭ��+P�mMZ����+)�SV�(P�M�(VVV�ڲ��B�l���B�
e++e
mB��
���VV��j�eeaB��B�
V�+
ղ����l�[++jՔ(P�VVVV��VVR�VVVVVP�SjV��e
+)�V���YYB��YB�[je
ښ�SSQ[P��X��MMFSQ�VV�B�5l�YZ�mM[+VV�l������YMB��+ee
��5e
+(Sj+P�[+(VP��+
��(VSj��+څ6��M�Vڅ6�B�P�B�
�B�SP�����B��V����+P�����������VVP���B��Z���
�+++V��
��++)X�Sjj�2��5emY[VVVՕ�emYJښ����+j�ڲ�����+j�ڲ�mY[VVՕ��emY[VVՔ++j�ڲ����++j�ڲ��[VV�(��+j�ڲ�5mYL���+j�څmY[VVՕ�e
�ڲ����)B�����+j�P���+j�ڲ���eemY[R�mY[SSVՕ�emM[VVՕ�emMEmY[VVՕ�emMY[VV�(���VյemYL�mYB�����+j�ڲ�Y[VV�(����Ԧ��+j�+(V��������YE
�j�յe5e
���e552�V���յemYZ����
�j+j�ڲ����+j�ښ��emY[VVՕ�emYMMY[VVՕ�emY[SVՕ�emY[VVՕ�
ڲ��[R�++R�+(���VVQ[VVR����[VSVR�emYZ����������e55b�555mE
+P���յ+V��5�emY�jڶ���aF���3P$�`�NI�����G`#~����`��OZG��]B[`�⻮ �V��7'$�O��m۴�[�*��靖����ڼp{K$���^��b����C��ٔ��ἃ�����DUQ4���ں_$�28��h;G�R�[�����x�g��E=�$ ��5�e�x�@ᩓB��!�So������DA@0�h����?�?ב�~��h��nM�\�;���K�ӎ����8^?�Q��wQ:U^0)������"�(HqK� 