BZh91AY&SY*�L���_�`q���"� ����bD>|    }|j6���$ֈm��M��EKj�����jV̠f�I����"T-���U��2�����-����"Bk3`�I��ӫ3-���M�l�kQ��*�+Uh��,�bf�&�m6m[V6�M�j���b��Ƶ�k*%�%EjЊl�����mH�Z44dy���Z�m��Im��V�)��U���-����Y�m���dԶƕ�fk���ٶlͶ���e+kZ4���1Y�V���l�F�
�.���Q����f؜  Uek[P}����\��U�ǧN'�=&�/nJi'u��=`���jv��kL&e*h������zc�B�غ�5��Z�l�Zƭ�b�   '{䯭.�Jo���ǳ��Q%)����B�]��+t7!UU{j]�S�T�j��¢�R���o=IPW�g<9�F�T���7��]���jw�2��ƪ�T�)�4�i)g�  ��%�*Q�O{һjTy���t�R�+ޯ^xR��Ek���:�J��s�UJ�+��w�UR�-="K^�
���{Y*"������T�jT���l�61ZسYiZ6b��  �R�H�������=:��S�(]>�*{�:v֚x�Zy�T�S���v�i���e]�����
�6���|*Gjom[�/����$}�����ڔQנ��^J��6��lT��k  �m��D��=�>��)T�>������WK���z힫m��S�}R�}ڥ*w���|�*U�����J�}0S�{K�*'��ҩ�^�=�ES��{��Jْ���{�m�R[�خ٥�  ��EJ�k�:��=�-���]5�J���f��ƥ=e�^��G���9�g5��ީ�z�x^Զ���ý*��`�M��g�z��L��֫�U^L�Y�٩�6�CUXH�  �/�O��v����t�zwz����)J�]���4<�)�s�9t�+�vǼ��/m%P󞸽��!*���ރ�N�oC	Pu1] ���'���m�+�6I[cJ���  ���@���h�m�z����E^��{�{�4���S�� ���UR;����zUO=����w��E��YYk6��ږȭ�B|   Y|>�.��q�@Ѥ�yOz
=vqΪI�7W��ATs�� �^8��4uX��Y�[��w��J��'JU�ٵ5�H֕�ڥ^�  ���QVP ;����g =m�x{�H9Z�^ S�zu��E�K��^�瞵Z�=�(Q�_      S eJT�F 4�0&	����%A4рFL�i��d�OɈJR�4b`4`L 	�D�ASU) �    O QS1H4F� � !%*hުidT����D�1���i)�}��_�ԇ�}\�8�����
�!�q�2�)�fW�5�d*��ǜ�� �{ʝ�� �~�(*~�TW�Q @�O��?���*� U���������ك���@*���~������#���+�2�� W�2�ŀ?�� z��3�
z�����FW�W�� ����9_X��@��=`O�@��=e}d�S� ����=e}dX_Y_�+�	2z�����������/���/�z����W���@����>��+� z�2���/����z���!�+�+� }����)���"zʊzz�z�(zȨzʈ}�YQYT�(��"�������
����,"����
��!�"��!�
��"!� !�!������ !�
!�(!�*	�*!���*�� 	���*|���� f@�Q�C�A��C�C� � ��'������ �� )�")��̃���")� ��"����(��(#�aT=`T�I�D��P��������D��D��_� �� ���)�(��(	�
�+�z������z�'���eY&���=aXS�D��>Y�>XC�e>XC�>Y�>XS�A��=aX�S�aY�/��� �Ȟ����e�����zF����M1f��5J�`���FZT]'���W��SL��L��nԙ&,���J�ݒ�l*yYd̊���Z�f�&d���F�Z�3��X�o-���fղ�;K��[iV�3k�4��s<��]��]���M�
�&^�YwVv��F��M��<Ԭ����� �+w�{V��W�ݭ���kb�ݽ�D�m���և��!�a�t�b��W�U�;h��-�r��B�rE�-u���]�Ml7���[	�W��kE���̏�<��Se��aF�a"�%�@���{16�������<�e@�٨Z��o��	<��[N�d8�jV����OJժ\��P*�
���6�� �30���,�,�[���  K"��͋�-N�:C��o&���}��b�^wP�1Ӽҋve-׏��X����91��[I�n���%�ۛ�SM_\�k���O�7�m%aY��)?����[ܷ*�ՐÅ[�Ŏ�K �(���h4��DlQV]�؛W��:����s1�񄄎�I���5�`Ճ5�=c�R�
���r�ҩ&�*�$f��ΰ�DCH�i �<n���ZH�c"q��Jœ���T�^�H-��T����փ�YS*���p���*�EK����B� ����m��EkY���-ܭ�6K�d�Gc��*�Tu�81�J�&�09�	�u���k0�X�cx�������{���xa���]30�#Y�=y�j�Gj����i,ԩP��'����~��Z�&����R�`Ԩ�#[7[��f�X��ue6�_҄+j����L��nє��1�\R�r������Gvetڠ�M��B8j����PسB ��;2Y�ׅH��C�10�h�U�&U�Fբq�vu7��Iӣ�w�qL����)Պ��k�a	�-8i<2��F��b�͆�W/
������'�gͣ�R9VÑӬ��&^�k��@Y]�v�f�trM�OU�̨\�-ˬ�ӺXw#QL���`A
Ӆ3��fn�n�����s1����b36n�+=�t�m����Fm@ ��	�R8+h �S���#X
�X�6iV\�i���"��ѱ�@�a;���:�mY�WO(Ztm��7e�Z���-]i��A�M��+$l��:1]���VՋ��j�P��)�D�V9��2]<��jMGp�J����S!RГQ��卭�J�x���En�[H*�3ZF�E���U�^�T[-I,rW;o�Z�,i�'W
�Vt�\��H�nn��bY!<I[.Sk(�z������4w�7��l7W��Cv]K�1��e�a�aǹ��Ʈ�:�&�U�V7�oU��L���l٪̤��7/1�,GT�Z�(�e+V�r��*��>8�#V�bZ@�|+�{�mA�R46��	P	��<�del��`�I�1���!��vV$k6�*��zsBZ��hE�GHt�[vFw��e<�`�<f�a�7ͫ�M{oҰ,X�'2U�lm�F�PY�V��V� +i���Y�e���kS�y5{�U�PO�7�B�Q�//"�e$7j"�X�Pp�uwj����@�*a�Cu����H��	��o��A�WY�:
����!����f��0�7�%� �dni
��`�Su6��ù{{,�u�ėo)ӗSC[H��u���
�e��4#F<���]�
�xɬMIP�٘�T-l��iRo]����&���*S�li�XOqM�p�x�����Cb�M:"VRM4���m̬��hXa6d�&���J�L��H���ӕ&k5��%i"���[���j��";	B&�Q�`����Su۩���I!n��t&�l&m]�T�A
�u�0(5%����L�U� l�q� ;%'���mb�mVmjV����%(4�=�R�No+���*�3�n�6-�tu�	(��ͼ��j+�̱��5J�;�ef�U|�w��I�=��Ø�J�n	�� ^�Bp��ֵWu�hc0Q��X�[��5��O]'�'�7�xv��B���ۋ^��H�dQ��"U���c��,$�e�X>	ZC��ý�Z����h�b���~��z[�ֶ�����єI��<�5E5S4Sz�X��X3>n7�J�v� �SoCs]�T��$����m���5�+��9����>13*�I�)B���(*�3D�[�����֩*�9���Ou,ǚ��2���E�)�-Z�zV��*��%oq�"���	�֠�H��.Z
e+.�Y��Dއv/*��w{�����ķb� ��mn֓�s1=ݣH"b����E��M��5��-S*�Fޢ�nh2���[�^Q�&� 5M�+7@��C��B�R���J�R��@
#r��mbf�R�Ed�ū��d-ոyU��H���TL��av��`�Zkn�%�u�Y�;

gX��pt��[Zri�&��IҠ-e��5��u�QT�[tu-ُJQv��(�1lՙIU��1�׹GaSp��L��%Sp�n�IK8U��`�����X#JF��Km����4$m���Ͱ��EbH�W����ԁr���1O��Y�QGpQi�b�Voh֣��F�AY��9m�l�
#rA�	���.6B։E����xXF�?CwL�ADú�a�mY��Š���Ĩ/ei�ɂr����9�n�2Rj�I-���R����+{zr���-/��E�[)�#^V�XJ���ej����	�QI����6û4]��ժ8�JV���I�oI�Xq�F�[��.��ֶ`J����d*���`�.U٨��qj�	�� �"�̼wxn#cB���� Q� wu�%fƍJ��I�2i�p*,�1��f�(�K�#��O�Q�\N��΋O0Ш���Ȧ��-���z�+e�l�[1f��T�����fF��4Wol�Q�YI�]X�C4FD�z0
ݤ�<��`��x���Y�V�JJȖ��O� �AP��Qg6l=X����Y�q:z�j���V�W$����I�Ų�*��ͭ�/!Ͳ�Q�t$i����m]�t�V����b�h!ul2OZ�P�YH�[N�Nԍ^�<�ҽ��e� ɊL3I�-�o%KaHk,E������e�dڹ�i���݈�N���H�Z��TcU�aJO�Fv�.�Ֆ��	�N�~@��
�7S6����Mom��6���bc�e�ܬ�{K��%�.�̔�YkcɗJ����^BѨ��]ޘ#DpD��XYm���n=�Y��[Z+IHɶ7DI*�M����X�2�ǋfZ]5�k&\���n�T�L�OkN�9���O�P̻���.z� �%��p"��z�
�6Ӷ��wA1���;]�������N��� �B��c��9j-����Y�uB��J+n��(���cU3�.�TзA�G~&���&�!��9z�r�ܱz�ڲ5�c$Nm���lS����n˳.�^�c$��G{��\�9z%��P5/q-����qY �4k�Ue�Z9��$q��!嫤��h�#�g�X��77�SJ�"��lܡ�wyp��r]�W���2��A�+�Mn|ء��];�Xm��f|U���5]��^F�b�XF�Z�*+p��*趭���!ZqY$Fv�v6azsfDEMW2W��5�4��* �bXp)�LX�Z�Eމ@��$�f�,>�� XU��5后�ϰ�Eif���n3A��5כN�\b��z`0�T��"�`r����2�^Ff�֩���J�ݟg Ao&pU�h���i1Tv�U��9S:�Jƍ�^c0ҋ�/+j�q�K,�"5������tp�n��2鯴b+2�+�yŐoW�xR�V��ض��|]>O'���U�aF/B���k°d�L���^6�j��E�hn�]��LC�r^TU��L�Y˽yD���xR��a
��7#U�E�-)�����t��v얚Ub�e��Ђbi�`� ���!�A3cu�� ��Z�1c.�S@��y#�p5!.�kN���q%[i���R˘&��
��(���3����E��kE�U��t�K�$f��5�a�`d5f�VPR�,-S#����F����\r|Ξs,-t�ȥ��r�Q����'��l�!Uu�Qf��R*[�Z	����޲Ėt�[J��bo�X"��,I� )K*��oYw���An���.���;(ڬX����tbz+Z!�B���GHQ^<�F޽Nn̥V�����A�+z���y��#c%^9{OB!�y��Q��/��W�b7�5��f�d��kpS�)�m��Օ��Z�V�,���ن���p$��D�cUj�+ú���@�ʬ'o
X��F�W�)%ZF:�-q=��Gt�.�&i#�]-Պ����>n�+��--��-fl�;�É��мU����x8v#%)�N�̷�j�a�6�Z�W��G�h�^�μY���Ͳ�.�"��8ayP�yy� ��oӆ��jn�k��-iԕ�H�PG��ݤ@V̍)��q�CqI@jO�cG.m�I��,��:՛1ZԢ�Q���	X��uϘ�[���n��d�ڼ�Z��5"���ɍ豘��\�d�����%�,���t���2�څa��Nk!қDb.�|��2\��2A��.�;z�E*[�ᛴ��^��Ҟ�|Px�U�/$�܆Ҭӻr�	�]��\:���x./[`Xkq���R!@ǹ�����1��i3b9#��T�,����RaVl�o%��VeM9�i�����a�ab�*0a�^��X�X�RW�rLGmc�l�������7P�;o;_é�As�&��6e��8YEdWZ��;M5�}��BS�@6�j(���������Zr ѣW$�&�Ҝ�J�Nի�X�������P�y�gr{�h�Fe%����ݞ$ ��g�kk������nĘۨƺ��V�W(��nA�l4/u�tv7jS4^M�#RP�+(�3�N1�p��L��L ��E��!��*��T/^ ] >#`�{������M�82��H#J�4$��	2�ck`�2�	�,���1�f�w,�ݎlx�[sk5X��t��[�	�J��"��Җ!�N�%q��mcvMwgS/���X���F�U��r�(ꎍ��8Ix�.���(�s�%z�*��)�&n��.)YV�B
[[���%U��Q�aG�%�1��Ui#E%t�p���2�6,��5Y׵l<�PWC.J¶��p���ެ���t�J�0%Lv��ن�I�M-����l�E���(�y��`���#bͬB����ɱ�k&��L<�s*٢�ګ�j��B��
�	܏���q�OM5Qӕ=�3mf�� V�&���F�n	s̚��ʻ�o�ԅ�Яx�y��1��:ܲ� ���Ŷ�EIK6����p��2�KC�F=�;�ml�Q�Y>9�ʃG�C�x)_0��ָ�/Fު���X`�W�&U*�%e^;�&�,�n�&x&Y5=�l]�נ�.+�m�R�(���R�.���-Os1����t]�Rj�m�Thj,ي��wP�오���wJT���=� �E=(��4U�s�[d�R�] 1R��J��P-U�'Vk���U��iH�K�"��x���B��P���6��r��^f����T`c�a�z��&B�g7��������'��.����*(Z.6�$��N��h
)V�n`��J��b�V�;����Q�T ���a�9�gr�F�0eB�8��W7�e�����*�&�{�2�^>����0�4�ݱ4��J���I����b����H�]\-ծ�Q��|)Y�CI�G��2��Uk�7i�|:÷��*F�شު�.�m��P�
8�,�+/�F�<���DS��t �4��:p7n�����Y�Y�1����)Yѣ�>�y,�
u����n��P�)m��	a�M�o7��n��F�j=�n��B(1���)T'B��%cQ�tׯ-��46���p�6	�G����J���De؇,�p+�M��*	rLcY0L��*��"QV�*�z�[&�Zӡy�5��Y&Lx-�0+�ڧ� 1%�md"��L*���И�P�$��Gb�A\
jXM�Ŋ	bnh4�VU���A��4lgBR��V�e�%]�9[+.�Rd���4s]#�Zp�f���X�48;zb(چ�i��k[����Pڧ�tƕd�0��Y��?P�#�
q�
��ݼ8L�Yg!�Z�k)���$3\]�Φ(��}maJ�4��cf�k�J�j4t���L-�r�����uU��d0]L�;��wv�
E��і��Zk�`�A�B���G�*ʭ/7em�owSPRby��=��wZ!�����t��jb8(���^X-n^ٛ���\�.�b���V
շA^ԋb�M�ZG.z�[���R�-u���%��te�D�5��S�� O^�&&$Of�Z���A�,���EY�fe"3z�ַr�8kXړw5a��i�{n����^�`�đ4q�%뀃�K��zP7���2�7�Gb�-s"ʺ�O	Ǚ&�E>b�o�ӷs��-.s��1��b`��x@[W�f�_��ц�������y��_+/�E�̖�o[�C����7Nօ�e�s����n���33,9�!�k*�oz��{Uv�ƊFv*���Nc\��Lꙺ�&��dj56O|2�8x�/cn�i�;e�;$��3v��������bZ-w*�訅�"�)C��&�^��!��2<�-��H��]���#��
��9�$�W�����!.��Z��n�M�oU�.�2Uf�zG��}���Ǥ�Z�g�ے�5�F��C�jv����0~{�ro>o/���X(>^�X�	�����9�pw=虹C&N���&��V�9
�u�d��>6�5+�Z�*4����i�lSm�İ����\�\�B�����v]�K�+[`��\���N���Z��N/k�CGHB�u0�{����.�e�ݶ��P���a�/s��Ԯ�X�Kf�|�AՔ�[u:�p��ԍ�7s�ɴ(�'U�Hdv�iQW^P��K����(Y|l��HeGw�k�H]�}�T X�n���>��^/v5,V�E��Y�e0�Q�t6A��Ɨ�`8�;W5]�oi��W6g����3�QX7I�;�J���C���w��u�Y	��ܬH�Z�h���[W۬͢n����
H:w�Ԏ=��ƍ3�b�	s�ɻ�b�\��*;q�g��)G���D��ټ�۬�����(�r�T�)��:vx�l�7S�AMb.++�L	��'}��K�1���:�)���z�/Uwb����5+��'S����s�����j/��ih���P<k��Um�T�Xu�/4��c69�Qcy�z���n��澁��t���bc��ׁ:%�Ӭ��V���FR�^e&f�v7u�uu��P����7{d�Sz4VA����7��T�v�݁M���J�j�
���4қ7���S�V7��;��c�|D�CT}�x�\y `J�Ĭ���mLbt��w��K�)Gk�[���oY��bm�Ի�M�wp�۪Rh��i#m˗B�-p��U��P����n��&Ñ��1swMwt�q�J�����K�8u�և���"�A>�O �<�j�v.Ȝw�c�;�xf�\䗉R�g��Jg!��j�m�c9m �T�dǡI8���Z��T����Rc�
�*o%3��[)�66�tҲ� 2�W*mD�ŵ.���.k/1�M�U�W�Ր����Â�%%/���2�d�c)�8Hmۈ�F:9�[i��7;�E��%+��AM��:$bW�'YM,NÜ�)f�g7�s��w(��v�͓�a�Q��u��\�{�WR�%׵��f
V+�p���f�D�n��2.RJ�=S��n�w�����7N���H���/fWO��c��AwEݰ�/a_�^���ð,�P��d�F��m3�j>���,..gg=�^���捻�J+��ؤև)�.o��H���v�z�δ�1Н�ҰT�1`��Z��k˽C&�3����V(��A��]�nQ�-���!׆��(���;��=��Gj��֮��gU���q7�"w�ފ����u+X�\}�1.������j���u�>��~�cL���-{ܨqԎ�_=�JG���)tn�\͵p�����[Ks����vJ0�m�|�Nh5��Ұ�[ht�K�����r�TÙ�����М֞�3�ikxM�LN����t���V���V�<r�6q#�Q�BM�����%Ӈ6�]��%X��x!$�f�d�+�\%5�m �oaklN6<�U�_1+^JT�9��ʹ���Wm�mi�DȘ�p��8p;������gǊ5�c�LVc�n�Lb�HA�7%L��*�wS�Z+>,�J�
�*4�Rm?�K�Wb>yG����fH�d�Z3q�'`�4�
�T�1m��o��c�ȱ��g9������d��B�Mt�33��4,�GE�?�7|۰Z�4��]F��q���#.L�Z�TP�ݩ|�6zz`c6����y��M�f�� ���S7���������k���%�[��$D�`�i���=��n�'nl�`#�hA�:�����(�Z]��j�MU�XA��kc�����I��-�|���P�)йbku�0,Q��,�綹�FɎ5��94ư�=`�lr�̦�\Չo(jY��I�NV�p����&��Im[�WP�1Y1�3}���e�:^�%h$�%������V�A�uݗ�,=9�4�4�[�M�K����Ov�I���֒���r�^1o�H-a����<^MaW/,ֲ�U毻8�\̅:�]BL	L�M���c���&[�\�o��~AG��� �/-Q,�H?P���ḱ�ז���RW��[��ܩh���(�w{[3��H��BQ&e��l�6��cq�Ճ���:Jb���:þ��o��:�A�_eX��sN�]���D�Qu�3L��M���e�L:�K+�#7���]⫼��^v�ލ��JA��Q0�,e�5c�oxu��LSA�S��E$��u7���{�1�J�;�R���+��"R�����9�S��
A�_>u39�%zZ�ŨI�i���Ѹ� ����9�S�m;�q�M�j-qW)�5�Lx��<��T������\#�`tҗA
PMw�!k��_X�(P�i��w�����&A,�TU���-갩L�wT^����oF�2�D���+A�@ľaU��-�׋��R��:Ӛ�/w
{bH�ɠ:����z�$�88�|Z���ؤ�Hӷ2����U�_Qk�1�W%��	ҭӫ*;�;��K؈�Cs�^�g�6�0G��2�j��[�.�R��yOmZZ�9ٲ����w�����X��^<��6��o_�-,i�����n�`|p��1Z���&)����zQ�KuR{,�[rx3z[���a��aw
�,/��/Xt4R�
JR��s(�ך��1[T�w,ל��b�8�Fv�!�su�T��a����v��_:L/��1k�*��|��x�읦o9k#��(�d[|mp<��0�%A���&��]���
�;�ѱB�,nV���浦�d�>��ܺ8��ٗ׻ۙ1�8���%'đW��>|-<X���)��>�}�wIW~Y%����o_56ͽSw0�ݫ���bPʘ�EK�2�y`).r��#x1ۧ�r,��n�s8�E�x��'7(D���D�I�%�WN�k-:�`^۸~u�th��0����qś����'2�Z�҇b�Y̎e]�ӊ)�{�m�S��[���
�kw�0Y����6R�'�Ր���2�1���T��,̸���S��*�+PM9{n�!�L@�]p��tїw$�At�#j�����$����t1��u.[����սG�����˧^��{U��9>��{ݼ1C�.���Z���.�i
ѽ-�$l1��5!��XzV��ҡ�5.S�n��f3])�1v����JN�5�ٿ�\�(������Q��h��r`z�4��KU]�&�Tbm0�^Ǐ�#@��+5��\���f3������*�_J֨>��	���]˴�o��f+��5_��M=�v��2���1R[�����i�rJ�\�NmA�1���µdL�|�������X+����^r�g%�h:sX5��]���;���*�)z�q3����2�-�C|�SG3K\s�)�5Z�Q��>N�Wi2��]Q��N�S5yB�:ژ��̉)�@�Cg|��ܽz��ycy�맶(�y�X�_Y��)��s��/l��^��t�d+I��r�),��w���+r�ѐu�0(ꢸ�dȪ��\�gP� �l��|��t(Ha�d[���o�K+"6sz�g*!S�N�kTC�n;�㩼�Ʋs�e���c�̬�Y��ꇎ�Prȑ�7��G�Y�#*1�iY�y���H�0��]m6���䯵[J�pr��y\,U����H�����9��B[Ջh��Tj���I|^n�ZB�Z�tM�ꓭ]��z�K�lf���$T�,�q�Fe[yV��v�ncӄ�j�V�斲�����B��B�1CᚡN�ٛ9�Fd��v\�u���5s/-���[*득�Ik����bAf�g|��L�o��˫S����N\�'V�5,0��s�l<Ä���8�i�����]�I��x��k)g�,�ܩ��A�2���5�u��TՉ�eK.����tT �֞��z����g<��vo9xr�⑃U8��/ ���&ڥu�4,�Х�	����+8Kw++��68xs�w���J���V�6o�m�X����l*����s0պƩWcޅ��^����z���m�z��:�f��t��1rg4���)p�1v9�U�$�-�×�T��{��k$�W���h���7�W�l�/��I�Rq��&��k���j��M�{ő��s͌A�0O�z'z�金�x��Ɩ:�_�j�Z�:��S�OjQ����VvVómGb23
Ć�ķuK.��3
t+C������d��r��ùW�1b�t��PD����P.l	0'\�p8�JN���jjۢ�Qz*w�ECB����^O�-���4cӎ�P�W�:��/�d�j�ɱ���DU��v
J�T�P���{V���E39��Y�]p��]�'dX.��坜Z�����>����!4���:f���]��R;��7����5S��Vw,��u��΅�	�]wY[s��M�]O��=�ꣲ�M08�yV�,�Xp�WN�Q�G}��!5�+y�U��Ѿ�7մA@�qzZHI�'��mA�؄6�>��z�=߱��!w�trq|�)�r�w�������oD�Ż�y�zVb�}Ȩ���B��ԝly��S�\D65=ӻE���w,	?j�yړ�ޗ��t�9�]X��	��Zt�=�֛�]5�|����GѺ6^�>d�#��	�w�C� �޿m=ȧ�D�n�[�����{��K��,Nj��+1snz v��,��W�d*��K�n0���B8G�fv������f�.=�{��;\�gNɊ�-�������/���,�(ɋ�yTA3��kg���E+��Â�{z݋&�U�W���S�����Ҵ������&��y.!"�8�Ae�^�m�޶���hL�C�qk�[u��|P[Ⱦ�O_�;蜎��wwr0.X�M��O�0�u�n	X��o3n�G�!@�MV�B귖��owk�r���GE���l�O:ʥ�� ��q�z�7ʻwC��y%5�}�u��<��Cŏ
���(����AWحt�=�t�5a l�F'�L9��C�Uч �`}�3��Q��{�������s�������&"1gI}��,�;W���t�>v��E[f^��J�s�n����p���uE��~�@���Pk���h�ǆt�'*�!s<%ff�NX�q��w��d�Yl�.�%��R��e	pQ��*�@R칸+b�J[ǫlhJSr���,�`	��˜1ŇV��s~�]#���=��E΀��m;��.�gk�gq8����T��so\��:�qﵧ{k+��ŋ1�Iov����`˶I���Tn���T�x��S2k�v�i��]��0Zph�l�㦔.��k�$U�&HjΤծ9]��UD��"�y8�l7�R�d�ݞ�s�s��@,��Q��pm[�roh��1c\�Fq�n��ޚ��c����:}���Sn�[���j��VE�:�jǬ�Xy��+�ړ;�udqr�ѩG;�K�t�hu�u���ΗWLش^V�$)���K����A<���m��wD���N��e`#zwT�WY�����5;\*hY�xF�l����y8E
�x��.u��sr�=���X�r���̥5�x�Rň�$zVy�B�c����:/T�ԓ�\�tg��-j���pʻ ���c�����{���a�h����p����'������:z���VD�V�{�	b	t`c��d�o���ck���DYb]>��:+8K>�I��+�J�AٺG�v�}IgX]a�;����5!��A�f��d��$�t�څ�v ݁*�Kr��X�C�3z�*u\P��E5'�m�y��Žz�|{���}k�����U��P4���]�Ϧ�];N��q�G�Ek�RZ詩�(� ���/nS���&��,�Y���u.b7��w��f��]�N�XB�k�Uu+���ql:uxU�A��P�8�f����C'(E�o\L]�ޢ�V�G�C�S;��W\PtԵ�|c�q�}��%;��}�)����������f.x���K�0\ ������!��$-�9(_�D>����|�QS/��3x���!BI�{���ݭ�l��.>(K��ˎ��ϭpR���L�]B��t���ٝ:Y��x��8��xj�ff7�^*�Z`�U}��*њ��)�A�8�7
Ӽv��R]N�&==2�F.��۲���n�0�#�U��P�a^Tf�w��}�8Ҷ�����.�W\Uf�W�Ű���s��523��#��Z%f4b���ɾU2d�
���>�J�nj$].TSN��<X��ݥ��j��M(�t�W��R����أ��2�T�X��>��+�c�l9��agd�q�f���6��9�p�I��gx�3\�6z�A���N�Y��82�e�p��Fc�BQ��{���b_;]���&_��L2�9:um��h��&���k:�~��Tۄ�B����}ܭm�ђ���O6	�j�za}���WK��Gƚ�-N��"�-rJ��v9��y�vպl>��7Y��66Z�e����|����A|�g�N�X��E��R�!87$�7yٝ/�U��e��yt#��d�L�SZ�D����9��Q�Q�4���7AΆ�|:8Fl�l�I�x���	٩\� �P	��[��nk�2�[�q:��Cr������J�B]����u*��|��J2c�&�}R�v@z��<w��1yWw�9D܎v�!IbT�t�R-P*1A�A���I�%PdS��T���S��ti5M"ˤ�P�F���H�y���ȋJi��;�v�n�	.Ur�&�H�w�H  0��)��zq�Yb�a�&)T�[pCІʠ�vb�P�`���4B�QB��I��t�M�iU1AҤ�[�o��o��������EE�~��O�� ����߇�S���QE������ _������w��qN���>���F`��B�b�ضգ�ϲ�����Y�T.HM.�0�Tfr�I������+\���U�?v���&��6Yd_^R�p��^̵Ut�M�^	�pS���+g����J�@�gSu��]�=����4�f,CaPzo���#�q)�]��VlL_N;7L���Ԏ�&7.U�>�@f��!y���#b�G���g]��4����c2� ��V�t���I�V|�N�ͩō���Xⅺyl��ܡռ��.V�EMZ�'���6�6�9�j�$Z�M�u�,�DS�9�G��"���^���4�fS9P��º�K�{�"h�d��gz,u��5B_jjӭtM�gpow�N��6M J�N���=����IY3o��l�w�\X�������v�AޛrTB�PG��.�G*y&�`Qa��廃��n:!������כ�1���+g6T-'���J�ō�
�7�qn��WCwd�H����
�ŶTP��������yW�$�y� ��`���U��8��.x�M��y�$�ggE�qE���]��a+�L�t�{�żt��A��2�i�������8:�Vr�ą	]�f�L/��t+.�X�.=����>�gz��q!B���t�뱄p��tл�w]��:3"HZG6�%$���3�i�޺�jih��$�U�<1p��a���据��׮osT��p�eI��Qǜ�9>ͥ�*gn�M�k�F����y5�FIEu�ٝB��h*	G���`�u��
�ѺI�d�5w#�t�dO������cL\���JL�jj�)PEu��m��|�Xsbn�4��M:�1��ڵ�٦u��c��q�]��Q��WI $u���5�
Jm�2��Ifu^�c��pWzNG�j�Шݒy��1Kܩ����W7���b�iN>�J��_
�}J�j9оi����.�J�袦��������n��XI��s��[�E���e˵u�\�vӕ�\�X�{]SDJ�b&�N�L����w�g��9�3�O�3D.v��8�2SyW���s��&����Gm<̽A��LTM.��&}|���o2\y�6�0���RV�P�3�9��P-��k�.�x`}���7�ԖZ�G׽4
/2�DN<���B��C����YL����X �F%�Ӷhm-�HL�[bg��k�.���/�X��Z5�f�L����`_r��8�C��*0��Q֮��M��X�[�JTj��6b�A�"��Ɋt����Vƫ=]kSJ�N��eJ$�n��'q��͋;fuhOf���wK�&ЎF6�ܵ��d� �j
�\;x�L�ܧ)��ލ3�޶utJ8*���I_9i���Ί���V+����Ӹ�7�oi�]K��R<2�O���8���k��==�s���;�w����T��W�����n�I>/^���FE�E�ܭ���JT(ͷ;�[�M=�����4�[3&���X��C�����}5fU¹X�\�;�M�N�5U�.B�%6^����t����#�)��ɝ�z���X������1�(,済*<���x��vQ���T�.RE,�9�b�V%c]��S\D���x33��Tͷ)T�w4�r�2�7��
gJ�T���	���N��ږ�	k�\l`	���q ٘6^'�����&frc�+"JG�.:�/��]�g����R�Ú��f7S�f�	d�����A��>��!T��]���Os��2tR� =cS��Fv���9��ee^��H��9���۫�ٺ��ǁ��41�x����i=�Wv*n��7���2�R��{Cs춒�2��oc��b�����.Y�e�:6Tm�U/��cm7�ي�#k�^\������2�X4���y R�u4B�����p�=�AՏRə(+ݤ�]z�)8��*@D���'��kX�1,R�&]��\����L�Y�q�:�/��&�X�%B�fj�eS�"��<�<�_Z�x��v��
X��(���{+9
���e�48T�,��]'+�߆�����3�}A���R;W��:��-��N�$�&]�1]���1���I�AJPCN��n'T�5f������+Ǉ&Y^|M2��I���q����Z�I<��aùZ�۔q�4���:h���j���@AU,|%@ޞ�����ʛU��.��ѵ-����p_.�NVA�mdp��si_c���Vk�է�u�Pc6jfC�1{�&�.�&8���9 Hvxb[0���;B����KfPz���Qh�>�b�]���4��p��n�y��F����f[W��ft��GWd�.ј
S�j�In#X�3)b@$w]�j���,�Q�����X���
� ���ѕ������%�sw-1�7k��n�O���SV�Y��Jt�p�r݊n�`�@�z�-�1�V̵�Sƹ'��ux�V<en�Ӂ^u�0=N�ޏV>cG]윑m��Wʑ0�k��v�Y�O;.'���y�@�7pUu<��è�ĥu���ձLk��K�H�B���W�f�����V�����+n�[���*]�G�Ѻ��\B@�:�Mxk`�IJ��f1�V�锍�Q��`V�w#��T� ��:)�[��#�i>�Q:�˙���w ���Jr�ڂ=�v�Y[8��)�a�d���#j��{��I�=�/5�Ԏ^�fp�i�|33�zd��x=��u�ض��A0s�Y�fr�Khi;�5W�C��j�#����K8bi�sݗ��*����S�sW��<���SV���ֽ���z��&�f,hJU�j�V�;W�3)c�vNS,1�+VIAb�>�/kv1j[&h���33-F*w]��	�Wqp��=�&.Ýp��>���P4��x�tX:1�B&|0�,�Ձ��@Z�YЍ��u�ޤ�t������Y�S*[] �7�����5��b�D5�Z����XN������ԑ�G$P=�h.�ݲ�2=r��vVȀ
-e�Q��*�ݓ])��eg�{8��K�fY�N�'���Ժ��k�r�=9[��p�.t�VcV7�����C��u�f�p�����Ѐ�|��
x9�7���5��Bʂ�_L��n��N�i��.r�Yh֫�&`�N��V(�%*��@F���̺K.�f���}��@���6$��֪�Isr�k��Zw_T�2��"�Fce#\*,<�g�J�h�be�1��c�HLJ��z����n��Y\��M����WW�T�I������ػ�3g�q���M����ʓ��OV7�މ�[Z^���v5�+zV�2�:�f�F����L+�Z�{b��54��v���e������G��+Y�+���A�|��޳}bh�V܈XoR/T�6���%�/K��v
0;������d�F�X��F�(Y��F�pC���ysxɎ=V��ɘd�tEiާ�i,&V%�o�yZ�.��W2V�nshfևHzȺ���f���헛M��(^_,�\|�B�Z��10�����ϝ�N�MTX�䬀76�ɕ�5��������*����{���ì��	���0S�q[�Sr��]�%ܝ�^�)����D��g7O�.���+�8��Td�{q��=g���}�-��¯e��O:}`k��0�����7�vX���n��v��~rI��}.���O�}��B��:,�7�+��ݚ�&ԓ���WS	r����gko�D�nPoy��먳��]˲l'ܘ��a+���$�;%�.�kp΁g1ǹ�-���TR��0���>�MF�p�n��N�7U,9j��7�e���������������m���t��]�P�:�ՐNU"��g5��чx��n�����G�X
��(�u'��Q��Wu!Pfh�ʠu��4�z)Kt⽝��6�Aef��y_*�v3���5|��TpĊ)T�.��Ba헹Sf}yk�����	�˫��b.�i�,���#�5����:J��ݭY{R��|��֗\�ھ�v)�m�b���s,�5���R�.moL��e�I����rޖ���kq�+�bF��ף�f9 �2��	e1� �`Jc��'0��]�X�ˎ�k����u'Q=��(����ܹ�+{e�����B��=�.������!@ ��ۖ�ڬ����H�m|e-Ĺ��ח�\�lm��r*�$c�o^Ҩ]Xڀ���tlPF�����Ҳm���tb;�ڭa*A*�]J4W**�]��,���i�#i1��O+�V��t.�n�����K
ᬨ�Р�#Eη+���e�g�b[U.�6.�QLܜ�(r����h��cK1j!odT�t�|�����
��ʺ=pc�˴;$�|5s{u�B=a.��D�}�2.4�(L@�yc��.�n�@�j$�7�25Y��at�Դ���:���u�$��V�7	>�!zʋz�\�����{B�@�~[���k����u��
��q��[��rS��))0Min=���x�ګ�Y�[:�JhmqB�v=��'a�ݾ�(�J�&ge��bb�c���[Ƃl:Q7O�z�邢a��qx�1�����Q��Yv�3�g�d��݄!�oXa�n;���{EX�9P�\6+VaC:a��k�� �
2&_nI�v���:�K�&p��P�f �8r;��Z���XA���IZ�����W]����Gj�G7�8)��ҵ"���X�{c�h�M+-�j.�7���a�iK��:��9�{u;]��ݜ��ȫ���R��q^m=%�̪�z�BS{�ʭPx^��1#��w/D�C������x>L�lY��J�רv��|�f��*ʅ*Ӿ�� ���X��;V4�\@vR�n�� ���O9��0��|���1�V^��!��B6�Ʋ"x�Y���esm�|ri�-h������}{.ּ��ʲU�t�fJ�����Jf�Xܭ�b�
��U/�D,��=z1+�=�{b4�m�m��gR�±�Sy\�lta� ���b�$,Q�1�m��uw�V�DT��Q]�|��*��ܢ3gpK�+�S�����.op�+dv��=emp��4�s+�*i�q��`��lH� G;x;����$�e�{�V*��9Z���&�8_`\+e"�u���%]u]$ѵ4/٥��R멐V�<a��\��<�2��WN�d%rҭP筮kJ��0���"����z��J!k����s%�g�ۆ.�wǔ�ӹ/SQ]l�N�YE�5�=��]�]�' 'P�r��ܨ���Z{
�DL4l$r�g_A]���H���v�0Ѓl���c��J܊csW�l�l�Ob�k�-�c�`޵5u�q��ׄ<��f�n�&�u��X�]dJ�m3OtI0C��h���V��#�aPΜ�^c���'��Ծ���+ o�'9�K���͑�s*���ӕe�u���d�%Ns�,�j�]��\zc�VKۺ���tda��r�`}Du�\�\�Y�]9T<��::�q�N�mu+o�kbR\����y��5n��Mn��=�%�r�n���h��3E����o���-��]`�f��<Xɚ������oU��I}�Pr��i�j�׸���Y�5��V�z{R����
C�'�wP_oCN\�,a��(%������5]���M��s7rA7���J�b����W*ei�E����c�8{��v�PTN�Tk����/8�3��I�Ќy�]��
u��֑����r�`��� о\:W��1R��"�[�nG]2���Z�;@���A���x&N��;i4{<4�<4ݢů�
[]��e�_5A���qv"	��9�<�ՙ��m���e_�,�o�y�C&F �\+���'i���.�-�蜼%Qh��+�y\m�N̷ʹ�(6�:�S�6R�q[��d�9��4��T᪹d�kD���/������vo^�"��z�璐�_���k�	+�J���0�/9�ݴM��m@��јn�2t�
n_+�I=MB�F�A�;"0�\�y�0%F@݌�2�*g9�{�	��"�Y5��bЊ�ӹWy��;ئ�j�K��\�c{%Ըb���Ѽf�|���oD��L��_T`]�����}W��܎��N�H���ݩh����Q1�Ӷ��b�纹�ڤ
����n[;�f5̺R=R��u�B�u�{��N\�Ɯ�u�e�[�QA�G�r�k��k�N�]��pμ�9=�24�Hr�`�Õ�/'9_p@U��钑��C	*��8��P����˅�q�Z3QkMYr59'���yݳ%�A�zSi1�U�X����(�[�*���	��Fo�ھ4�i�a"h[�&���x��U2fd�r��x9	�����V9��Hr� �/��9���Y�R͔���D�u_Y�6�#�k�Y�8R�a��x�ִ�B��2J[ �u��ؙ���W���Yf�7YVI��v�BR�VK��!\��?L[��K���5��/v�։K{��}�J����DU�F@ka_
e�4��S���k��KC��"+�6h���_@0��.]%��Q��u抺��5ۖ{"���v���}Q�kS�{��\��Ӥ5$���;h=��º��˾��4��n�&�n��,y�kh<�:fL�/)s2��57�F�x�3=i8ܡ�v�9�vr�0L��Hee�*D�s�B�1s��vit��7��
L��d�.nG5��wm[��X1�wyl*z��A�M�Wt��&���]nN�������r�����&V��|]�A��i��]��Uɰ����ı�ӜV��	���z�hq ���fl�՚���%�?�߇�~_{� ��}I��}�����/��G�����{�?G���������fs������'�T���鏅IN��(Q0�W�kι_�v!  \J���8�̦r�ͮ�L�J���"&��[Vn�ehm`�D�-OE����Ҷ���;nˣ%;5���^�Z�*��Z�������V�nqw�t���;2�-Ц�V�F�����L��u|�J��ge4Z�X���.��&���>��+v���!**��,W{8�j�.�ۆ�������x�˻˙B�Jڗ!E�Q:&β�v�VŦ_0�6�RU�K=�� q�|[�I�v��J�Nf+^h#r'OA�wH��M��Sk0|��]i�rRU,.� ���*�@T�*D��nu��G��v�s$��{t�'f�Q�D�P��$�Ϻ�W��N�mJf���:�f�G�vv��_>�զw�:b�(d5n�]F�#Y�]���]ԌL��.�>ô�����uX��:�g.+�t�HD�]�Gd}�d�{������	3oR�V�*�
]]�E���PH:Y��Yz[�J:py��ٝN�n3Gٴ�߬�R휆�S�] �u��-ݓ����)��$���N�� ��k��6�VE�rjU���f�+�Ƒ�|��/6:
r��4��#�Bk��^���{Z.�W];J.�6�ae崌�2���R�a�^(�؀=�W��6>�+�˧��	�(��A�=}N�ڤ҉%E0��
�4�&�S)�7I�E�
1ƫ��j�{�j��ACcX����m�cAMRP�D����uѻ�TF�4T[`�i�`1�==�Uv�v��@�*b۸^��(�&��I�$I�֫��Y��j���8���s���Em�tk�6�T�3&�(h�`&)h5VãIlhJ��t��MuF�:twdz�j�&�j)*�lR�l�و��4���[b���\]��v���5l�mZ,ƺ:���(:M�*�ѱ���l�GE='mv��K�7c��4v���b�Z
6�h���]�i�cZ�m�H�(����d�ݝ��MvzN�Di�(�Ymeի:*��tI����=Q�. 6�5�Rb4=u�c�DPv�ѱA��;��"]Rv�q5]ت�Dj�1�V�nꢒ��J����.��������՝�Mi��[u���o+[.:��	��nՕ��n�{�[�R���ȫ_�&������
��J�������l�*���V��9+�J��8	0m;3�}	�#��@�T����h�8�� 0Ğ͋�zAs�٤��M,ۼxv��6.�ct��B����=���>����}���6�5{� �[=�u�lߧ�힏�^1��������'���BK��*�xE:���>���E��g��`mm�>���S�zM{�l���"prUB�b/�����5O��ދ��J�G��,�qg,��y�&N��}{B:�:b���l}r�ޜ�|a�c*�ZxEcsI����{��Y�{���a�4�!�����V=�~�+��`Ǎ����9Ŀq����<���&��4.s>�L�ޡ86<K�{cƪk5�Wy��	�6�I�9c�/�`^��+�0lv��y�7l��R�5�@c��3� ���[���y�}^���}�P��8�z�<�0�q���\5i�����U�&�^3]�e�R�i��{}�D�&$K���&�AJ��ue�nS��)���e���"�-ݭ�p�ؕN{v/q�iu���3�jQ����w��Y��Ny@�YVk��<�_HV.�!��w~�xpx�p,�8.���)����W��o��x�W{<F��n��i���:'eS��f@9~���"z/����œy�w=��^�^`�&���-�S�u=:�s�e[�\G���K�h������Q�頪/e'�Gy��{�ߩ��{P�3��V�P�r�_�=�t�O_�.����Z���*K��Y�#k�}r4�4i�`GdO�H%���ʋ���QP֨��I��S���u�J��IJ��܁>��Z�#�3c(�z���t�K���n�P|���Cy�~w��q>so��ğH��U�E|�����ӗc��?,["[�|�9KG�t�C�F����:�^4�y�j�T���އ*8����O+�������{��CۀVt�Lq>}��ۊ9�wQλ���!�m�A���ø1��x��'f��d���W��f�+���y�ze�����ac({^�-bjx��Ԝ8w {u����껿)�<.O.�o�3i�cx>�z=�H(w!�����/��������f��cv`��u�@��ХF7EG]�%�Nn�<m��؜mlPt�FW(*�
�kaI{֬-7����vγ�+m9��Y���Px����kc�����y��߳r���ꧡ�|�u�m�T&L8��\����P;�I�)��}t��t����́���cT�}��v�XCmF���A����j&M�+$�cڢ��t�]��J����}�������0��>/�|HF<�U����uN��������fN�#�]�K\��^�w$ǑO��Q�C+��D;�y���3�6��&�rw,��;#A��h1ʟ2+���\�$�������J�!�\竳��U�򡚝F�:���3%K����(ݟF6�;+�[�U�֨�2PR�_���닙nppNa�Ϋ�{}��1ֵ̗s��:�h����ڮ�ڸ�޿3U������D]�KC�s|����2*5���1���Ѽ����Uj4�9}3���aۓr�#�K�NS���+��$ߢ��q�˼ۤ�[�-R�V4�}��ϒ��=��)i��~<�-��۠��C7A�K:��0��]�6�[3���=���8h�!р�D�+�ah/Te�r�UŒ��b� ����7�s���g��{�Z�%���3G�S�H��2��W����uOL���̽u];@Ѻ��Ιˏf���_�q���9J��W���O�3ˁv<�wT�s΅�G�.��mR�608��{�L�w.�I�9'j���2g�m⭴����]a3wD��"
�p�6�׆�t��=��{7�>i�ZQޮ��}�ْNM�k�����H��>��r�v��{}���Ȟ��<��;�sj�<�����z-��oU7ٔY���ڪ�Λ�k'���GVpf=w�~q!�����=#/���Ϗ�Ab��Y�ϯ�eu�N�Q[Ҽ�)�'	\!��92/T���7]�в +�Ǔ!1����zl䗺Wj�5��^�7|OegXɽ�a��;R�6��^0��[+q�4��%�h/t��U�.���E���my����hn����Ilڸb<Şu�^{}����W��N��Wi!���SrlX1d�8Ζ��Y{/V=u����u�����a>�^tkun��7-w)�q:�����J������uf��K��VJ�f�F2��J����_b�1��
9}X��	��w�M��vj?P'K���'��!��m����-��-��|b�#3�l$���_ެ�Լ������(��"$7k��,#]�np[6�a��G�e�F�V�y���P�!>@:�]:X⏌�f��ӛB�<���V1�zP�JFk���uؽ[W=��c̎�����t����R�5���-��Wb"6���]fTг� �2F���J�s�Ҭz|��]'#}�~�z��6}w�cf&'N�� ��}�x�f���L5=����e�J�y�G8((4�ٵ!��Mt���lo�X�"���!I���d�ow^���)D�a>�"���'*vUO�[{�7�w3�/�oǉ��S�Cn>`zÜ*,4I;ƞ��zH���T�^_~�d�����Y�>�W��N���S����5l�[��ĝw�/N��*4H���պ���Fٔ�����n��t
� JF���"���p�K�{��=��ΏN�EE�X޻�e�ݩS)u�w���i��z+=N@N��N�X�oZ�t�Q7{�R�t�)j���>�"�
�ws�3�Q�h��-S��y�,N�K1!��ך^v˹Y�����\�$��}�{����;z�Q��m��*�_�%����vf�I��x����~��W����*�h���sɗ��@�u�%��bW�dyf�a����I������O����};��d;��U�ķ�k�	+p7�ԍ�U�*9�o��� ��7����e�,���VZ~���<����OdLh�9eS���X(56�z�ț=e���w���<����|3�s=�T̺�hL���^�WL��t�2L����f�ަ�"���ð�1<�	��~\]���CC�s�6� =��Mvd�Ĩ8����+�-@���8h��{��%�2:�,b��4��
IS���=T7������q�q䓂��z���t{34E��/Gx�9�&(�T�n�y��"��;/ܾ��*oo��{���JB�Փ�z_�ܙ
�KV�j%4�:��1���-EX�O%=�ޠ2H��m�����V���z���e�hxhv]0ئv�$�ZP�z�9����U5r���0CP�]J�b�"vC'E��ܸ��:�.��vDfȦN���pm�+=��`;_<0�]7k�Q�}q=!�d�v���&2��TY�m�b�F�y�+�eP;��({l7u�澇Ps�O�+zk�:����Aټ0g�d� ����vN���e�~�&5��A�{�{Of��Stk�P�	!�sKi=��Ǝ����u�ݽyQg_�ޡ���� �������?Q�������Y�z�9�^/=yc�l��M8My#:�̙׹+�"�xk��7lG�[����v�ef�zx�|'�tN�5�����	n�T|N�q��0vu��˿9�n����a��S.W��`MO 0��W�9�P����
��g��c[��d�F�S�O���7}���7�{>���<�pt��Q�!1b{�����[9�%���H��1�d��a�z�s왝�a�z�w����<�-<�z\~�u+if���
�g�CwrRy�O�k(SMh�A}��R����)��;j52�]�59�����S�Y!�K����n�ym���"0�j�a.��x�D��Sհ�A�Z3�����U�����Wf��L�=x���n���"��2\�ِ)R�,�Et��\����7.�˻ʹ��16"ѕ#�6��ˡ+��r�%���pK��/8M�?l5'�WK�j��Oa�$�����ީ��	�y�j�O}��T��!+���ҴӑZ��s��_>��3O�Kp����	KS�M���˦G��X��D�������r�q�@��]���*�%,����T�����Bs!׼��.����� ����O��[5�����j��~~G��,�<�ݭ��z�1�2�N_F����!�4�_@�a8h�9]��W���V�{|H����y̯3F��W��=��lx�K<c��d���2d��'"~���\���l�+�}��=���L5�w5؎d�|f��5���Y���buޜ�OT��'&�z�f���ϣ��x{��i����!}������9��Rd�Յ�7��&�{@)W�T���.��8�`Į��7��PI�Z�*Q��gX]�ߴ�fۤ�HM��3��a��ݛA�cB��ɕ�Pˢ^����_1Z�J�7��p�6��u��JuǛx7%���y1f�-lj��ɋ���c1QV�H��������<��{�׾�_��N�x��Tʲ�U_�x�Q��Os���\y�V3���ݮ�?��zmW������/ԧD*5�����\����ǎ�^]�~�q�z�7�}��{=����^cC?O�뫠�3�a��痢��Gy����:.N�yJ�}��crf/zy=����-��\ӱF4o�!H��`�E�lO<�A��-��R\: -xө^�,ߦg`[Y��AO����(�זek�=h�6�U��j~�J���1ޡ�S�S������
eGCw�y����zd�ovuΞ0�dă�GE�u~�u�M����UK�.��^,ۇ�k"�Ci"'��]Y�w�9�b�#"��|��@=�?�lN�Mx�U�5˞]�0����R�9>��a��^�.o��gm/!�����=&[��V��r�0
*�yM�Z�N���]�+�+�wd���~��&L�!޻Ы���.^e�ǖw%X�L��5����TFm�\���wvWrӬ�v�+�c�m�[,KDQ�Yg��4�T�U�hn�s�t��uf`/��+;�7aC���:���7�>ފ�sV���wA��!������^j�����E��|�����+E�=�s�H�4�]����1��_��`M�n�m�ih�a���h��|��ӄ��7 �p&i��f�5�S]�	پ���KL��Mf�t�u�`C��/�ˉ9�Y��sڹ�ySr�ۡFxea"&�ͽv�bE�K�=|�5�z�}� �'O��W���_�t�ݾ�|F	uյ{��q��������Rg[��7X�K3������|����ʳ5z�_� ���S�M&'ew˽7D^���s/��j��H�Ka�R�%�����t�%������ݯ�Z{�7��*u1�+v{��>��B��<2�Ŕ��!�S��(���O�}�另���\ly��'��r�Y���x8ihu+&eӛB?�J��TU��V_�����^�w�����|G�������y�"8e���cS瑠 R��2,5�yu�Ut챖�c9;�Uj�s@ri�=�A�� ��)�W�
�c��hLç6f��r��.��9�/�S����Ev��6�pZ���9Vwl��9[�<	
ލ_26����@�i%�r�
���Zw�}nYI	�7E���|�t�/v����.�R<�{�rC�FgP\λ;�����;�B�3G@JBCGxϲ���~�7�Y��<����^����ݔ�NU���܇�m�0Ӈ�ڙ6�x#w���RI��y���.� iT!���3�Ht[�2vJ}&�*� �oVp�^��v�ySt�-�E�!Yo[�T���6�x���'F�9�d��vIe'o;*l_^��d����`�J6�c�7ib3�%�)$7!�a�7F���n�3�e��cn�x�&4t͙k-�qr4�e!�⑨�{|03_Q�Z1)��QKT��c�8�	�_j8e�s՘�.�,�Wk9v�s��ǹ�ka��`|A�Y��K=���I4-_xj�
)_Z�*�U�ټR�y1a��, X!�met�,�b��FXP:vS��O����K���6T9��c���%��){��f���⋹Y/C�`��T�i��9F�q����,�$�e�w�v�S�9Q���!A���ًX�)�4TGv�&��ep�Ŋ�u3N�l���Q����L�|h��;��T�Y�nٲ�D�溏;i�Wp�x���eD���{��P�I�Od��WK��my
:HJ�u�W���g�o9k�۞P@"ۆ�u�(׏K�V\��/��O�g,x���ߓu+��w^��9�䌁
7����)f�:i��T]�Zt`�7]t�T.C��n�mc|Xcp��p�o��»A�|�FV���X��ۣ� K�+l��u(���om�G�	�rs8��Is��]��b��U�@��t�S��So1�5}�T��z��e��hͳ��1]x*7t�E�b�	��3�M=u����r�9��j��7[v=�R�\E��J��fYWD�gO+�ƃ�]*�9�wn�+E�IMj㬴q6qn�� ��{r���C7jQÌ2�J��q��aa��mCrM��R����]�;������m��p��5x#�5�5�9�F����!3�l����,ET;D���)]:�T���鯻K�6ئ%\����2��k����z�3&ӝ�U�f����J�U�2�_����c:���$.���)V��Y	Z��5*�eܲ�dj��v�b�{���7u�zV<�U8r��V�N͙�&��`�!��i��cF��S{��r�]����d�\,b},q��}���[����E�r��W�v+�&�v B9˷;X]��S��ƀ��ݗ���^,�V[��	s.�Sb^�ʇ���z*���&��D1Mȷ"��9i�	��(�(7{~@5��\9��RU����qj�y|�
(�Dh��cj�&��lE��[�Z�l�hшkPE���vlն�݊�;w�Ό�b*Ӫ;���U�v;�th5m�������$M&#6���=Rn��y��h�c8�:ӧ�<U�y>G��^A�t9�˫����Y��my����N7]�2j�N����� ���=��c's�w'��Ümև�h��X�ݩ�h�0���Ѯ�1�۪8����4���監�Zw��I<�Ǜ��t����;A�uD]n�N�,^�͊j�1wc��w��vN�i�ƞ�zh1�I�y�::��(��ih��Ƽ��[�ˋ��풃E�M]Pѣwpk�<�8�A�Py�]���Myc���wG��SӢ�pw�w���㸪ݛgwr뮓���y��%u���P룎�'@EAA�iN��#��;n�AI����9�lo1���&�4�@h���t퍌R�j�1�%I���h((:�5JPo1ţ���j���U���[n��Y��ŏ1��(|��X�A�����:�����6-�����>�O��j{/z�%�M�ݶde��3�6�&*�kr�.��;��2��I�[h]KZ6���v��}���Jz��:�h�8�ǐ�5���Ⱦy�iw��
*Sz=���bl�0v���t�<�Z� ���Y��;K瞌:��I��Yr��w�n�1�[hq,O��N��:y�Jbn�9U�yPgGXR�ܰ��� ZeI���MJ��S�zj���l �BR�mR�-��R��l�9{��DS����N�+���8�����S>�~��a�TO����{�\�n�3l�U`�$¹M�)��Jfq��T!��yʑu4�eԂ�FMH,=X:RD�K"�qӷ���3V��p81e�x:r�[���/�:ڒb�B����wS�|�W�񟥓�2Ό�~Ξ<BܨMAP����)�Z��)?b�-w��K=]�IY�^29XM<�4��h�^�2:���9�J��tr��C+_WB�\Y�T���='�+���d�m�ӯ{k��b���*�s�fQ��ʽ�h*��/�긖�lV<���s��j��%�4��43n���&����:�����_{�c��s	���P�+�`u��q)���'Y���c5�Wp����m~���:����^c��L,*P�)!��ݝʫ5����.�]�P.�{�3[Q7�Պ��ɷM�GTx#�"L(-�[Z0�ɮ�b+�v.p]�*��s����o�Y���I>ŦR�ܒ�Y�����V�u�&v`Gm��l���"�rޥ;.~�gzr~ݩ���7z}7�.5���VDa=l5��X��f���Mg?� =MR����els�J;p�-����1���o!�Δǭ�$S*-k!�>��O+H�P_w���r�h�NI,��u���.�TXl�>�:��/���p0#k��D����Y�3��ؓ�?N�C���,���ض�`(G^`�N;Q�l�`A�j�]zҝ�&L��6"㵵�'�E��U�i;�D$]V?1ո��}��4���`cn��3�2�͗�Ÿ��Ipu�"��wV�ǋ�3�@)ZY*��`m0\����N'��%g�=����/a�B|�j3��a�����]��.&Ă���
��}0s�/�9��o碝&�w�ev�bv�5��㰦���]TPۦ�mp��2���L"�v���7��"֢vHy}�u�D�C*_��f��GE�r1�"x]��t/vx1�����KQ{�#Q�I��T�/E�m�=Ŝ���h��uxN�;	uP�eC�$D�?Z�ֶS���B�+�z!��c�Rz��\G�ݫF1�I�;l�@��o4��ܻFB�3743M���b'�&�NJ��X�)A�u��p :�p��ق$�(D�˓�J�6�,C#�t(A;d�����d�G�o�Vp��摮L9j�	�Qf �+CX�����oE���MU
)��\��Ug]�%�{��
�^p���Mx������l��L��"���������4N����ݻ4��6g�z��ܟ��n�(<�z��<븠���󌨳�=�Ӧ�7j��s��+��؃M;����f��B����dc�*ԥg�CL7���A��)Ɔ��C4�yJ/b��4'�ZS�0�%�{[u���L���>�,��S{\��T�	��<{:�sR~[�lzs�gs&��.��tT�*��>(�L�D��o?R�$�WO'�P4sǎ4�N�^�S�f8)���w� ��kS����^��dv����Z�Er�%��T��(�V�T�fJ�Uür��w��Bfsu���pf0U)�]N��Gs���gǬ�'YM���cV��MOpZ�cq��� 5&DÂ�N^�����ޠI]cp� ��Q�q�Ae����׫�B�w��ޅC��d��k+��0I^��� h���;c�s\TOFە�N�VQ�EF_1�luoeRdC酲�	�VȟY=���U�G�����=>�ʥ��#<��o&n�5�E�m3�&TPl���t�{[�,�r�^��������,�yJ��K�V҉���n�<R�z3���RN�0_V��A	yv�H����խQ��ͽZ�Y��j�7��k�kd��>����[��43�]�����ކv\\Nۤ�������z�}🲜H�w����)w�1T�����p����ԥ6���>���4C���+���m��U�A��ć��y ��^
匷͍��9�ݐ-�Sښ�K���hLf��5��pe]lԷ�^�A�w\�s��q�U��G�|<���H'�;u�������{�I�Px��3�����_�#\i1�����Ph�S��P5�K(V;:�D�s�1��M����t_�d�b��JL���5m`C��[D'[���`3aN1�Y9+�XL�����Z�,�8���>}���Jϑ~Pʩ:Pd�e���g�Y�,�j��*>�W<��,5;x �gX�9U2�85M��̬`�ĳ
i�K@J�{.�@v_ݍ��:v��c�nf���/Z]A����%:a`��1n�	U�Ѕ�(��	3������ܳI�-�1F�*��|�NV�9��I�P͐�pԇ��J]���JJ{Q�/��#����~a�V���IGj9���4�n����oZKV�Q��)����P�Oa1B+����A.�
$v��}�&��Y0��t��q��*xA�:Yze�Fg%:����Z/<,�gzY�5���x�͠z��ζ�ձ���yu|x�b��K�̬O>��D�'�hCi���cH:gJu���ƺ�����r�����{3krC�Ǥ�7��ƛ�S�q�k�"�l���}��-s�<͘�|9���V����]hly�a|c�0����n���-��w0J�_��k�9md�Q���w����Wt ��-'Z���	�p�0Py�T:|\X��2-�;�D�O]�rxC3�fU��n���>����.�݈�����#�5�8uن��p���^tqV��p��/r(��k'l���/�V�a�<��{#��ϯ۲�- FmjD�ͤ'��]���U��`��	=���2I�F�ycN%��|d^��%�DL۸�Y�6غ���7�=�b�p�0���������Э֢M>�VPb�6�r��P/D���p�����.���w1�h�:�N��	1��Sɋj������ۡo�,��޻��&]���N����7�Ls��^Ȼ��N�Z>��ã��r�U�����TD��Kg*�ĸ�TS?z��{�h��ü���ӏ9{�n�eZjxIO3Z�ouě����m)��(Ju#T��zE����u0�{q���e<eU���P�ED�|�A��,[l%�M�
ڳ3����`y��
J�,(�7�6ڎ�{����&�ߝ����j<A�ċ�&n�������ˠ�Yܣ6��V��p4���-����E�a��x!S�ͺ��Ȩ�<%^)�9�>r���`�1Wpv9ⷥ��k].�uKFh��gZܔ_R���fU<[��Su��]����F�J�W�T�z����$�s��_l��x6���ߑ�
����M�T�=ߒ�m��w�Y���FF��7�)oA���u���9Ѹ�l�|"=��څ��K�<TZ~8���,�a���_��7t�V������mzc�-Dv�#]��Ts4vuC;N�TZ���N�^�풻���"cs���D!v����j��8�a3�]�b� �A�c��!��6u��'��ӟS#��+9���x�nS@�j5�R6@v�`U�e���lA����v�S�l�r��~�}'���	e�J���\e&���FK-mo_QhJ�cRH����<��nl�{T�\�j�"/(���4��8�]AR*�*����¹@��L{5��RW�6�*'���|mi���7U�RO����W�������u>y�)�l�`F#UZ�	������m�N�[��A`t�KqS���i��[�կW�CuS\���*�}"��q�����~Wo$�Z�4�c�M�ߢ���Q��4%{>L����S�|�qށNMqYq��kJ
���E��k�-օw����M�G_淼���NQ	���J�.����fE����O*�e�tZ46b���i��yhK���Z�@��H}0�\�R���ټ���[�v�J�oc���or����f�'��m��\Vf8�s&�R͈"�K�]���>�l`���{���F�b �f;نj��Z
>��+�	��5����gi9ʠ�>��#&S6)�Y�1�W��)�xWk�'V�i��	p7�]�	uV�73�{N�\L=>��46�i�9Ƴϙ���iS.9��x�e��cIGq������I�k�Lqҥ���x�AM15O��wR������CP���b�m�P��aA֪Z���U�s�KhV߹V���-�x|��8fy�����4��<�#;ŰӀVJ���?-�t�g#���L|�!;��ض��M�ۄ4�ȽG��G�T��bGjM�;wSE���m�:�(<�%��t����MϦ���3ţa��EWb�^={���'+aꕥ:��ʕ:�{"�h-��	�F�A�m�P����yXi���ի1҉�N�ܚ�����؁w퇚f�X@�E*2.=��1-��F�fTnd5d��z�y#�U��0��O0��g����[W�� q�J�4Yu�G��?7�qCq�y�ǔ�}I�_0�ڭaҌ��U����`�1��H�z�花�6�k�7A�J	[5���,�0��_�{����٘]��j���0�5�$[���B#d�7�zq���Od�W\/��V�>�-��W�u<������T��/�8��sW"M۟ @l\5���a��gD���ȋ��5��;`�w2��M93f['�9�đvǻX���>����
�Q��!���/��ζ���8���R��G��ۣ�m}��I`�.����K��e���!��Ñ��
��F���js~�GNu��8�_�5��fH����{1�7{�B�i�9�tD07Z����+^�:Y�(6�C��}^�aLɍu*�w�a��'yT��1�mn8@�ַ�\юf`�6%��0&�?�Lk�p�����ȑ\�q��N�TD��1����8�֣0�����@��Q07�8ǗK��[�f[��z��|'x[,~�g��rV%�_'C<�oZ�ѴMS�{��K��>�s�P~�����X�Z�&ai��j鵍κ��ӡ'D�#�*�`Χa�R�Y�-7�X��PCm�H��5V;���z���Ji��HGjx�GvF�<)�?Wˉ���m���u�} �yߩ���n���R���R��a3�{�~OB�տƇRg�� A ��t����2'ť��V4�Ez���_���'2�����x;��[Fx��T�Wp�I���T�L�4�~a���t�զf�w@R����RD�䚱���e��`���L̮�\�%�x�*�pV�
�v�R�i����O��fR7�*��qK��؞��1��L��_ѪV�l��/��J�;����U.7c�D�S��ɪ�S�˶o��b�״{=���1B�cL�ő�a����%�aUL��iU��/m��(����uqN�X^ˣO�0�&f����75f��N:���:M"�[�Jt���w;�1���;}lD{�P��J�;�zsoX1�1(\��{�v�^�!7P��ok�Pz��\X1J�|��6_[~m����1'�3w��}�Mg^}�WA�<���YnF�Jc�Y},}��h���\����ꎊ��zON�E��3�c���N�T=��"бm�:�鰇�D&ޘ������u*�g�I�m�mR���3t%��
�ým̵ygYwF�7�7�
��p�&��P����{h6[4���a�Me���SI���T�f�E9��X�xuG���{5�i���:�Yo���6�/fZ����O��I��_e�It6T�m�:g����z��"2�Mx��u��#k\3oѽ�Ƴ�g2�/*�l�#�)�`Õb�et��Ӭ,ဵ�螡��36\��ha�M@ ��69Z}�y�vx%�F\me��S�B��=H���j*�q{ ������eu
������B�>s�H��iy�\��z-)	�\]�t��d���G�(�̤���\��L��.�8��Z_+��ę�+1�Zov�%�E�����*��wI}���8{�`l:�e�Ku��j�چZ�H7'Wz1H8Pف�z�߷�xxxNm�7��������Q
��J��ӀT�bڷ����"�=%�cs�FzGw.ǫm��?���i�n��x�.�م�(J�`��L �Kv��O�yMn�c���=IVGMm�:L�Z���� ͘��Ko����^���,�h_\":�&k�(Ju`ev��kAz5�g:�L�~����ն��AH�5���2bķ2�%�M�Vְ}�i6{��h�p�R촢%����5��6	�O���D*wk�2h���oE'I�6���o4��Jo��)��z�Z���-�d֚�s[f��yO4%&�K��G�׆���P���')����k:��T����]����0Ù%s���m�5��_��Ǖ���[�u����2��֦��Td��ݖ�8-�����H�\�,����v���!���I��Z>��}��}��!!=u�����XvyT��m��R�Tqua����x�\p#h;I1RE���X�Ŏ��l)LW�2r4��ˮ*E58h�٨M�{)mo7�QhH
���+�$�[Pః�����}�o_�����}�`����>>>�U����1}��J��
�����BO ]p��%���DaLp��.d��n�{�ZQl�Vi5t�ު��`�����
3����f��w{����s����K�����h�WV�d�/��S�u�4{.D�;��XR��6(��[��ùyφ�z��Ҝ��N���-�M�U�Ees7Q��al�f�bQ����QǇ\E��ѓ�G�[����6��׬<���:u��q���hǭ��93^�J3C����4w]�hHu,��׻W��RZ�YAT��B3y�ŔЪ�f�4\�� �5��hI�<Y�[�x��+��Y3r��w�u�C��Idh�n��-��p�n�m[���:K�g)�����	nR�(���b�[��`�xe)��	ڎ��c����f�8+��Ƥ��L>��cZFR�yh��na�A8�Zݛ۰�0��r���=�z�3uN�Sj��U.�m<�J�Ov�N�ȉ��)��aA����æ���F��6%�n�L{j�d� ��η��z�����̃S\w��.��k�C�,���uf��žg1�qk�H���%�r�f���ٝݙVa�C
sJ�;�2<9x����Jc/BѺ��9�n����i���P�VJ��5�mU�}���>�\̦�8�H�oRº�3��^��7(-6�U����ٌ���l����wD���R^d���<w�QJ�7�c�^Η�غ�Z�B��f�e��96h������ƺ	�M�;�v+˓0ћ)��y��OZHYO��t���Nn12�F���% ��i4��T��3"����噬k�:j�"���<q�aE���C�9hg#׈,{�,F��e�1<��֯6�&L�rn�_ �#ԁ#��·+ �:����V��n�u:d@�llY}V@�:�w�NW�kof�����c��U�U��Ȭ�;����nڅ�m�������M˼�������+��#��sc-F�ڙ�|"�^g|�o90����FrFV$���#O
�&V���Y��8��rq<�AV+�Z��p�/uj�W����a�Tƚ0'u.��$jO݄�U��m��nP{��t��8m�`�Ћ`oR޷���L�$��Ǯ�aR����w��Od�u���N;�v��U��k6�^\z��Q�C�����;��sW��f��������"�PI2idvs+��l����/}O~L�ʾL<M4�y2���[0���74�g����V��^L�خl�u������_6�z��G,��H�X�����
y�H9}0�5�h�J)S��Çw]�N3�q�2�0%m3`ֈ�N�r�=�p�iZ"u��#�uy�5�����b��v�ՂJr�j�SP���oq�mQ� ػjS�6d�&U�J��8`<�&�0^�е)�ŭ.��n�;��ns�b��4A�`��qL{�1�92L�a�R�3zs�JS���Y���y��^�C5��x�v���m��e򘫓�t�!D 	L�d�i��:
� �	$�q$�J.�	�>��|<@ UQ�i���·K��'M!��O#E>G����S�'vth4Pbi*��Z.�����z���H�C��M�tt�&�)���;t��h:B��":M:	�j�ݐ�:��AEy��I����ۻ)�[Z4v���!�T�t�Z�$��۠�$�ĕGy��4u�h�H[k�)��A��MQ��i�lK�	��5N�*�!m��m�m�:Z��A�t�b��u0cl��i�MQ֞�vtww=/N;.�5ѣ���t�&�M5�M:�ib��4j
(z�ә��GvX��\]e�b�uv
��i(�ưTC��bMQD��шthi�����[���"���ZZ�cEQ�F����GGT=$U��b��b�����+HD覨�Ѫ"j��ݹ�km�RUV#M5A].���l.��ƲD5TU|��af�O���*]��IB��T��wC�2'�/5\�o��R���&}�bk������
��)�n���z�#�z��?�c������x�<���*%�����ߩ������*��S������03^0�z�#k%��a�w�M۳��i�'�����զ<�mkQ~U�Ƈ_����p$hc,��Uk�ԽK����h�]�L���R��N���S4y&�u#V�uԶ)�[Y�0޶������&$�����J�~�{�Q?
Z?xS�1��B@Y!�-,�e�06�˘"�q|�����f�1���V�"�+vi��d�Mu��zR����G�\�����ւ�F'J�f�{QLu�84<�B�G��]�s�Vl�>���/jԴm�hB;����]�S���.��|ɀ�}fE��6�&P�Q����ˡ/Eŵ�
E��KP��C�FPn����������t�jzeهX�t2X�͆��X:*�䊨������Q�ɋa'�V���A��,���f�U�)�Ee��R�wdS�k���D�ýx�i2����Aj4କ���t���[������dǷ[b�:�9b���̀��=���9����*k^���b8M2;�I��/E��B�i7<�t��}�>,`��_�Bx9w�����\�Oa����G�)��OFW[:�Ll�������V��
ދ�޹�RZ�o���M|}:���AD�L�F]jɾ`�:o[[2m�^�T���j]�z�m>�Z��ytjE7�D��A{skz�h<�o��������CK�lYn���X�������:��2^�~�~�)��am�Ǡ��s��ԭ!���Ʒ�:�h�l4|�3C甭��4Qh3%��K٘I����m�?aS�f�m�SyC��-�<5���h�;}���;��r��u�]�?a��G��>(�L�:�Q�k����V}���K�<�6͹�k�M��;;�'���ȭ}�*ͪ��Q����0�������y&�MTs[*�&��߬��W��ƛO3�9l�2�ب�@��b��K���G|���}�K�dL�n�D���(DU��ĝ�d?1;�:��7ΘX`VK ��������P��ޟ����T����3����ݏ-:��p؈6c׺�S��A�(P�\'����9,�u�����5L�-��ΊT�W�S�Ρ7�fT��ԠlC�-���coS�6�.��oZ��t�t��3�f��B����qU�8d$:� �7
���IoLq���.���ZԽn�OQO��	��Ds��n��B���Md��;�'2-�v9:�wA��q!���w�Gs�R��z;��?Jmjs���&b�X@{�m�ۛB�AE��J3��;T6�Q�dӳ/r�HP۬n�tzܮ�$���ï�b��+Qj������l�)�����+9<�Ɔ�zLu%�����et��*}հ��f���S�m-r�Sw�������[W
��U��r�Tsz��;�����}_{�G-9HKm9r�_7F�����y�f�j9�w4aM�Ӱ�_��pp��uw]�s���\��u9�.��*�FE.
�g3hb�0?�/кF�5�DIھw4pV��{����t;�	ٸ���&�%n�Q�|�KE�O�U��XX"�07��4��~��?p��5hm�3���%&vɩ=�"�\��c� K9��O�'���feS�W*��Q䪑0dϙf�3f
��˘ d��jʋ�@�0'@^�23*��(tAe�L�k�4'�q�QDB�yT�U5s��&&��U᳉���8�Z�����=t�Eؼ'L
���$ն��u��ͷK��Z��(��8t1�,�\6㣆�m9Ë��@�4���!DQ}k��wE3���ڜ2�n���b���@J��Ϙ�s���ʍ�F�<����c���h�O'S8�࣯!���m���U��p�q֠^��05bI���ֆЈ|!ᛍ���v\ƙ3l��V�����Y�۪��1IG7-��S�-hto&��a`���8\j�[���9�R��̄�t+���L *���aJҧzˢL���C4+�ZΨw1cE@ia�^�M{b[*5�]���3�{�7ҳ�%�h쾩1v��6�m�t����f��w��]�wig0:�o�Vu�9B�rN�B�aq����/t�>���{�x��#jL���ݾ�[V�%E��Ih�Y^�rb5���ǝ�kq�0�sX)�ͽZ��e%s|���p�uΎ-���60��yN���좧q���x��r���zF�L�h�ls4rm,n���,"����,{X@�Z�3c��M�\���bc9���F�34S6�d�-������\�x�(��3#9	��ˋ�m6�V�E[#{p��tn۠����j6ѷ�tD=�  �޸w�u�%F�cO���o&uGf�O�0�UKY�ѥ�LRy�V۹Ԅ��v����{u�_��\'�\�ء+�0y��R�����8�׺k��2���?�������^�U��C'$<̞�ɦ��D8m)��(J�X���_8��_m���+*k{�8g!K�Kȹ�]ЫZ�t ɩdK�Eu�v��U峎��n�D��,�HAk�[�n��1Gi��3�&`k,*�8���J�G.�AtR~��E6PJs��&z�NH���;?N/�������">�T�o(M���������su����J-?�xߞ���;��f���-oZܹ��ؒ����n�tگy��?{d����<�OT�.�R�w挺�J
�	��d�b,�6³*�i  �����ww�ck�z�6U��%6������/�,X��f_�i,�.��ڜ�ɨ�V�R5�g+�5�Θ�(��@A��?{�����D�=1��!��hjp����	����:�����@���^�I��7V�K�<\]gt�"bw�#(I�;F-����C# ��?b�@��Ŕ9MHKʆ�	��f�5��Th8_Ҙ��$��.KS]h�]�he�;;!�*��/e�Wq^ζ�v�Q���bJ�VE��[ �?s���\� ό�5f��	�L�t�����0�ף�)���d��g�QhJ�RH�TQN�6D�e�+5�������S�Q���́3���\�>ʂ͟E��Ӱ���:���Z�"b�Z���,4�~h�[ƛ
s͇L:Z�J9?Og��.;Q�M*�A�v�\f9�%6���\��gww�u��@�Q�D,&��ċ�����-�M�����7f�dJY�*�cN�'I�Po�\@�[n�b�aPٱI��=cBM��i������
��@Aq��&�o�|�=���Dݜk��3��Y^fVTJ\3�����Z�W(��^�`��*���d^����-��]rq��H~s�B������"��A�si4�B�V�Vv�%�[��g�/�l���t��fwi��3u�6p�,�Pɋo�Ixa\�7�z�T���'c���}ɪ�ΙPv���oF�'܆��9�B��c�Q^a���G
UÜ�q�JR�t��N<.��&<������"n�`�����������N�A��	���/_k���x��P�l�wSp6���z��$��&1ݛz.yX'��'�"�9r�=qÍ�"-\?�.����)��uJ׾�A��,�/�䶅o:^&�ķ>f^V�3*�A{����3z�SnK��N�r�T)��F;?9��bUm�����u��V�\.��Ƚ�ku�ޭ�ax�ڷ��|޽�Hz*����sڎ�k�M~D�+��[$��Kh͵��L�~*<���ȚQ�5�v�[*6�s^��qeIΆ[|���CF@�#+�VR��
��!�s���be'X�)���]T0ɛjl8e�y3Q���t�9�)���non��!�:�<���^C��4�W��>yD?�φ�������>�>�Gi�:���j8Mm\����A��!�58���/�H�q@Y�\���/�a�Y��/�Ceﯯo�.U�H�	
,�F�P��~j���߅l��8Ъ�R�oS��ي؄���m�>��S�`�V�RHq�aը�"㦏
��Y.Q��jsb��H��-�&��}ڪ�^��va���U�YҺ]31�.��Go*h�qۗ��>EP���K2vu��h��;h�@�D*����YS�n{v_�a��V�?��;�z��U7{=s�(��G�k��od�$���h�]�*���)l�_^��_W�U_}�W�}�}�  � �
�R)�7q;��Z#�lD07Z�դ��i���Y���w�6k��O�R�9�y(���L�tѵ�j��'�a��K�:�.ML��6%���ާ�W�Z.�7͸^��3���kJbia$):�y`v�;
��V�����㹤��>[NR��V-E��&�����~2ta�^)��DdjqpJ�J��B.�5)��4��Ǝ��R�v�T����{����ˠ���z͊ZD����vZ�Q�w\��m:�A(A��Y���os"�Ӄ	���l����2#�
��g4�<�[�)�C�U}h���	�^��w+��4O���,y	��+�kH�V�9���6,:��;��@nWʿ|���~W�θ����0���3m�a���{$WE�\�=w	��T�b�%T�(2g��eý�������2Q�が�y��oL�[�T˜�M�זgz�U��,Ԫ^�4�W�v�Ϳ������mo!N����	�>1�v��ҩ�1)����{�V7W�Ok�F6�e��/Œv�P��9�F�^�P"��e�ϳ���&R��^�W|o`��'�Zk6 ;�Z�SD1��d����qG#�����SG`:����IH��q�Js+���yP�YO����8�Mj�m�[�k��ٙ�{#ި�IO��n��o3��/���.�6foN/��^�W�I����3{����f�*کhV�.XSO�i.�ѳ L����3�X(�͞t,R[ɭDQ~h�cD�Am���7p���"U�$���-bL!��u6z'�fnXZQ������9��&��[3k3�������S��Z�z�90�NsI����3U�����66��oLCo5��'���ڶ8�g6����$�E(��7�`�[y�kT�o8 ���a`��r�G*:�r�}��D��TyӞ.-�:h�6�r��¥�c�Ā��Z�-��hi��g���&��J[�!�sJ�&f�����"�2�����z���5����{�����@��S^�	��z�>ؿ��|��bu���]��Sius�T�+f���կf<p��3�螡�W\	�����ӆN21��� ��Cͻ��L�qcc���t'y�5���fm�8�3���]�5��z������⃁��(m�\��Vh$Ɯ8������xj;2)����Nn\���ɹ6ݱ���0�P�u;G!�9�w��J�l����*�L�з����8̭��r�g�6d<�]�f�mѯS�{.����u�nT�R΃q��O�d��%4n��k3U]k�'Př�w���@���W���WNmY��&��ј$�N�����{O��K0��c��v�7�LmS��o3�5��ŵ6��x��Rʍu�h6��������@������&���N�1׈+���)����5��K'���c�ɦ��N��e'�0��H�3E�?����ϟ.���5��B`g<�ԃK�V��B�S��s��7#z���5$ǧ��:S^<R�*�P֞�N��u�%F^�A���� �z�H5���s��I��#B�uV���Ѭ��SҢo�̖S�����i�-�3���>�Y>g�b�a#�JN,�4��OLV�!u;UT�`�ղr���f1�y�E���my�j!����ᵏ+�l%���ʡ2Ҵ��\��t\T����7�""������!Y�f�����|���/���^r�q�����;��j��JЄ�mY��Y�Ưo\��x�j���l��vb��/���p�Ó��'D�x��3���񜠼4s��]�"���d˜�M%���8���,h�|��wv�Wf`5�3��0�tČ}�Q(S�D���@�����9Ob�/�����*���þ?f�)�'��w��g��G��˘�2��{A0���D�\T��`:F(c�y��C�P0kS�В���A]�dJ���/�h1�y��7[�����Ȥ�ҬB�TU*�'p��"2f�Ұ���$�z����U�+t�,�%WW��3�}�ܩV�9h�ͫ��uu�,���"�Eo��R��+;e⺗�O��GZ���L÷o�X�4���2������~���A�Qiϯ����}8��+85z6 �f5�@�A�I4�o;���%�Hu�hd{o+���{�M��n�D�
��
�mހ$	�Bޠu�-U�ҽ���e�o5����;���WkeFd��ɭ�!�54��W�r�	�*q+��@��������1:W��kX0[9U��Iot�H��F��ǁ,�uMIos�3�qwO�P�\M��pl'���ה�1�o����L�I�hS��.��uj�4�a��QHA�9�c6b�pc^Jm��E��䍌{;Y[�b)L¶�42���=p��"4���d�oKA���Y�p"��8�~�.���_�
��~�Ľ��{�фA��t��C7�n8�ӂ�W�c:Q��SN�q��\9b��۵G�&�[ܦ�n�-[W:��i�{rEe�����b"������Kр�x�'I�K^T_����\2j�b��9�12���S�����㬫���V�ױ��SO��Fꔱ��Y�,P}�dj��[͏
�|e��I͗�n�9��!Y�o�4�l��V ����y�^�?�����}>�`���}�^>��5o&�ݚ��I��*-˙�l�����o��هoQZԸ���8�G\�*�q���aڢ�z)�U��M/2®�[�3�JΒ���dۙ��@�g��+uK�.�G�x�bӻ�>�Ώy�˲S�S��!�&�Ž�gD�=r�o�8��;����]��6�H�՘]v��[j�u�|�3m���q\*�-;�,��!a'|�g]C���el͙S޶��1\�)�T˸&�I�m�q)1։Be�uƒ튱	�c{u��[��ݩ�	Lʏ�Q�X�ņ ��:�����m�@#˖���r�wOފt��Ɨe���ُ�O��L��D]%|�k��Q]v�Od��*��Z�v=/0μ���n�~���?����=������O5���Ek	��C�E��.8�
�L��)��V](b��;ˈ�;1oC���
�_(c�m��K��(h�Y�e�a�r.��<�]nqw=��7��L4j�j_�f�
cr�y0I��2��+9`��Փ�٫vҾX.a�����Ё�\�H�Xq����]Ǯp��ٷG:�n�=s��=��������Ǥnq���0�:�M��0��6��wS[�ź=��K��3�r�&�����x'%�vt�GkH�r��ʽ�y���^�_*V��{G8�`k1����A��U�j�qh��쎐�{����a8�s��h�;;ʠ7���9Z��4)M�W�<���V�xFZ[�����	���b��J��2�]õ���j�[����Ea�������]�"�m2h��&�!�񴍜�Aie�Ծ4�
,�9����P�����]p�b���d-.}UҴR�\�[�ո��t?���g'dmB��ȱ�c�Ł�+;Q��ii���n;ǘ8[�z��dȱ[Q���9�s��-�\z̈nF-nbb�Y�����n��RQ�}q!�ZL}j�h}o�p#��b�
q�p��\�U�emN�déH��� ����W�S��v�,Q���t��,��=��޻�wW��K,���ws@z�E����f�Η��	��J��1���ɽ0}��fmΨW5{�]��TI���ٔEnV��`��ij�ѠX��V햸�N���Rŗ�i\��Z�j�G��g����eI}�Z���|1t�]�3f��U��R�*�@?�<�bzߝ���@h9��+9SȺ_\n�:	d�q�U�Tf�pZ|xL�K1���Ws�6Vt�rKkl[��-�޺�� �n�T��c��s�A�2�K�q����e�s�V�v�sAM�/�Hi\W�I�t:���N�Ev��(��Y&�v��#+Tꇬ����}}�J�\s�������Z��xB�̔MKˏ�־�]�<�50>.��G���MU=�iN.�]:�nC����v�J�4R�S���ֶ�m�-!�4D��V�m���GHR�t%R�ڪm�k�mX�cC�ֵT�ZM8�#�Q5�=/T���ZwcL�$E1��m�0�A���)�ѥ�:���Dt㍧F�5�����V��)�&5��1N�uF�]����-v���&�f�v�M-%����::H��t�`�b�7kPDh�1&�X�v�Q]h�UkDkC�k`��ɠ�4�bth4�t&�E��k[kb���M�!�]PP6�m�5m�Wgl�K���]h���"�icFqi��1V����4�_*����Wx�� �Fm��N�]�T���
&K�H�r0v�[i�Uv��J��]�́�O\Y5K�R�t����.*���{������|��G�	��U-��B�����={��%��^K��y"��f����<�T+69�S��tv��,1�4��K%ޖǚE"��&� ��y�x�EPn�F\Q�;�t�q��;jG�խͪ'�D�`��+�
�d��ԁ%hk8M�2���]{z�� Y*����N�2MM
	m��i���:�P��}!�Y��c��aa�XA,��v�[0�z��ۻ�����h�ձ�ς��q���wr�/i�����{u��Q�����$��5���q��p�g��er��J�dƧ�sP0f�Ŏ1�oD�4cѪ����Ĺ���ԉ���"M�Sly6��[ړepn(>��?��,!�<Z�G��0��a���O���+u&�����.��UlL#Mu=�b�L=��}��J��z1	�g3s�j�=?�7�Z2��5��y��Q�!!���C�n��/3]6�a�,{�p3���Ғck®����دz��.`M��e��p�6��b���YSJNl�<2<ǳ"�	�f1��6�*ߌ��5�/�L{ƾތ���{�Y�ƛɬmc�q^x+Ö�Y���Q��ܖ7����_!v6=�P�+:�^ΟF��+�ݜ�%������X�[tbQ��v�e;o��?��z���V���P9/~vQ��yٲ������7�:����ּ�2J՛���~;����׾|�}+�UE? �P"@ �{�=�G��t��k�૬�����Z7����*/�����K�F|��.sɆC �����EwZ����H�tP�^M#����q�Oֶi�b�oaWt(���ח�"��w�R9$��W*{=��m��hgb]��C_l��$��oL�]�U4���m��XQy'�j\���l��6o!7�=`h�vO�9�]{6izCϫ��,T�O)�
T��*i�z�E�Sg#��L�fQ��1Mr����n�6a�7�L8��\'Ƒqf)QN�����4
h�{��x�t\�tJ����������b�[�I������me�g:�V_KG����T�8f��+&5q�j�B]ԓߔA.��j/�N���XpWZ�a���(�D��ɧ���mF:;�L���1<��7rÓͣ����0��co0�X,�7�`ɶzj��>AY���O�L��ߔ�c�9xãyg	m9P:�����Y��N�Ƴ��X�*�B��>Ӵ�pO�O�؞m���Z��r�!ŗ����[�%f�8j����9�a&���]+�+��gU���&hy��ԅ6��s^�K�������;iZ�	��,{������[5y�-��A3�����7�Δ�η�ޒ�t��ܱ�(*���ǫ M�����'g�N�[�os��7��b�NY��ls�3sS2]�v��e`Y7�&[��ٌ�ν�{��� ������%G��L�p���G�6��f&�m!�+�a9�UKn�:Fώ���<������{�]��r�驕�stŘV�
!�-��LM0:�X�~���o3R&��2�U�B����&������]�RK\�v)��&� ԋ�Ӈ�����J���at�ӕ6����y3�;.��ۘj
��7/���sY����3d����s0辒�?�f(�	_@LѤ�B�n��jF�w�5̔`3���SOF�oMzӲ|�2Y��%�X��e�H�] �rw�^�����*raW�ʧ�&��_{K��/�:�34��L|c&�3��>k�ɕ��_�ٖ�-�k
1�;K�"�7��i��	�%�4>�ɱn�[������Fe� �eM|���(���H�;wZ�'X��/<֗�Re�-E�
ڎ�[�j����:7�l�|"B�\T�d�Kl�E��s�5��EN�5f�/X��r���L5�������ό%����kW[	`d8ʻ}�7+s\��\چvK���@EE��/��*��R��q�:�B/��qO���.� =Y�L&���x{F9h�i�r���\��\�󜷩�o1Qbv����.`�����u�Y�3e�p��b9���j����������N�\��tzkjnu�6�)��w=��r�Ҭ�Vβ���p�l�їS/�=�{�x{�7��"��wu�МP[��1��훜�Z�~��ɽ��8��r;��k!�**ȳ�����ؘ�3'kv���9���ץ�96H���H���T�,�M%�0Yct{�ю�J ���~I��M��x�_�� �+c�p9��b�@9{R1�`L�T�m��⹡=���XP!������K�V�+r��tn������JI`i�|����b�����ƛ��s���ţ��_��8�\Kcg
=v�K���Q��÷��I4BG=LG>�󮥱�ob\����13�BS���F�6��@d�G9򒑭�S��j��b}N��y06�.`�C�n�F�0�9�4������%���P�{��c���=%s�Z�� �ޗ�kI\�bt�a0{]m�v*z���������L&&-�{���1y��l���ĚV3�I/�0�v�%٣'���J�����u�O	�WN%���QI̔&Xc��L����g���z3�L\��l�_ζ��c���d���h��b8z%�C��P��^E�]�?W���M���|Ͻ�AOo���_�\Y����u�}ί�䜪�z+�ڟ��*�ڃ{�g=3k,���9�T�YRA�Z>3�{.Φ��9�u������r�֩$J�V��j�qW�Փ�;K�B�rI�u)[*\1�e���j��*��6M5�5ڹ.�Z�i�w*k��� �>a�<�� �0 xn�Z�n�e��z�;B���	i.^v���z#���ⱉx�y=�;��3�Ď�3N�,��'��ll/����%�b���m	�/����#����엣��B�.��ޣnX����bd=M����`r����&�X&Q~��O�B�n�M@��V�R��L�K5!�ѹ�L+YFZ��B]�=:�2��m}�4xnr�/}0���,y���l�f�l���U��kw�kXr����`��fJ�2ú�����q���p2�8���w�yEJe�:'�v*��)��eR1����~�C���$�Z��1f��6��a�5@��_(Z�Hg�g�k��Ф.�Σ�q]e����9|9���EʳZ�H�\�Y�vkXc��ن�_��7�LQ��9���F����Ғ��B;ݹ�u�ؐ�ϧ<c݆]b�Db�f� ���Q�v�Z�t���~NU6���Z��g[��$prs�,�k�����TV��9��Lk�擥B�g���ͻ�ѡ����й�,�{vQ���hf�0�n���c�l�G`
��^�㞞9�:�d�S���hy���Xt���U�_�0�U����
��4���s�JE�����u:Ⱥ�i"5rQ��\�5A\��ý]@�J��O�)��ڛR��<�w��(�;����F�ju�[]97��#z0t��}���o��`�7��R�H�B���7����|�����᪴�<]"8�(�������{���|`_yށYV��y��mrM��;R���jb�Wo[x�8f��_0��~�>�m���1k5�6#��h�lG���)<���(Iw�^H/X�V(��L�ӕ4�CR}��<4�4�Tq�n���u�;�g�g4ğ���gN�:�2�Zp���_E$�لC�5��ri�[�J���Ά�r�����}X�ZFb�ӆe��xAhK$����T�;t*y�+���,�UL�E���z�]��<�`��XO	EG#�_<4��z�o(d�r$�,S���,]��I��*��R��x��Q]׵��5rRu�C�v�Rh��{�$���2�λAUL��������V0����d�;���w���ܝv��ү���~�+R��F
,��܆�&��*�{bS�
�-������D���f����j@.�ŭ���)��Eo28oϡ��S3�X)���C����G8��4Wh�|���o]����7�9��JV9�|�C<��#A^�d���md�:G�*~+D.�1X�'/Y�Tb����0M�MeA�{�v�D�LRM�'obn��ξ��b��O��'X*Z���t{.�J���)v�{Yc1Aay�D�v�~m�A��؇�#���.���R�y����Јi�X��7'(x�z�ZoE�����,*��� {�<�P�"4�D�P"�  H��ā�G]Vwq�#	�����(���s�	u��Gc�Om�%�$Ƙ`ֆ��+���@�Ğ�U��U��j��Z�re��55�?�Z���)(-�c S~�%�)j�m��ͽ!�hlY��R)����%���ta�:~\X��6��&s5�P�>}*��Ƚ؋9�Y�|&��)��HT\u_B{�-�/��",�Q�͚�Ύ*���[�'R���AZ6��=�p<�n�k9�,�*��;�A"}�R����D3ly�ۆ!F�v�%r�˜aӻ<���*X���&Kwa�,���t�z��PXѨ
ZDZH�Rbi�6�.�O�
�h�[#s�����m�"X�ʓ��`-�m�#}�Ǎ��q��S�G�	�˃'FQ(c������ˀʢy^@�$�C���x�9:ޣޚ��1w��{���bD�,َ��+�0{].b�3��/o����r�:b=�[ "�MD��n�)�d-U~��o5��vY�3�����iL�=����1���/*�ս�$�In�vQ�aS�����i}Ɯ�NN_P�O�1�m������x����X!�U�;�騥r���>"����غJ�̫���V�� ��]%��<xe��5t���}�8�Y��N��}�\��!ұ��R�;�&3��E�IB>�4.i�pS�������"X�e�ښ���4z��}w������Б
P�B7��` f�m��pt%L¦Ͻ�u݋�P9��)2����f�H�s,*�8�+eU�G.Őn8$��)lvч�=|�@m�"�Q�����=[��ZW;7��hJLy�������Y3&�Anb��zy�m5��p��4��zO�B����E���:���L��[Ž!��+v#/:��x�ͬ�UE�3w�vC0�r���	�K�#��Ŕ:�Ut�$�|�7�0<Li[uF���-<�o�`<dיi����`^s�f��.��gN:ef_�*Fk�I%5+wc�.Y�5����W �!ɔ�B��3ݹYL���O_����^�4��FK-�3����\R���i�qr�����u�H�Uܡ��$B�/^��t^�=s��63�L2�k:x"e[.�M3y������}����O�|�[)+Ձ�Q&��w-1�B�Z>�����t묨���gM'����w�]�-.41�t�5U�@���^�r"i���H��}0�Է�ֳ�݃Ya��j>�Ab���U8ܱ��K����*^uC`:���&���t��~��zK�j�%q�v��
���Z���c��g|�o�q�uΆ��7��߷({��O��
���={��lm}u��d�!�n��D�-Z7�����f����sgz�Y��������qS�z�7)����G�q����@����ҨR*�(��+K�.|�'�����d�c�g���ҧ��&��oKq�;j%�H�)�G�ک-�W/���Ʀ�Z�U8g���3�;��/><�Cm�P���M�ࠚ���8���M���GG�Nf�g;Q�l%��o�{v�N$k	qMܝ�Rc�0:���ཎa�%6��Z,һ3oo�;�
/:Ғ�3Y1|�T����w�D �;,|j}��J�9&���ԍ<M9�XVծ��N��X{��p��Gm����D�dʀ�d{&SϩDmK��.� (��v��қ*�?V��tr�X��%65�Bd^��'�ĺ�v)�qT9q�"�#ݞ-'�/���;�s�d��Z�f��0,P�u�:�p�6�Ω7f�^EfЫuu�7B9[^�]�Ĩ���W]�k�mVqx���R�1�Cga��#yJ/`��N�TM�� G�_b�Ӥ���%��_�=��O�fym�h�K�i�0��E9���1G�?'���&��_T�u0��B�QT�d�j��V�%m$�ۅ����4�)`�T��tj���/���:��L�����y����I�|z�*�Y�v��[3�@6&��O/x�ܼ�l�mR��!���]ooY�'�����t�=U��0�׼c��^��Y2�M�Bh
3
�ן	�'�-D����!8Yx ��E�|�׈�f�[���A�6��8^S˲{�̻���$�x� ��{Ā �D(i��(����~;p�Hm3�ywJdp�a>�L��U���
%�5��;5�,�yk�{:g+K�X�-�|\Gi���^%f�v�OASf!S��C���a �_�
�	o.k���_S���k9X|ʷ�51\������4���N�T�+#�.�D1��V�$җ����l�0Ies�871�и�i3�%���Ν2�Z��eG�cR�v�v#�ާE�;Ri�9�1�@C�;a��*p�	v*�q!IǛ賉
��pjeh�a$�{�Ռ�z���0/[��N����x-kd3z��8g��֡�yH�ehU�sĲ��k���3�Y�A~_�*�����n��=���G��إ�He]��ўw����OD�O~�*b����u_`"���gw�[A�88y�yH.�|d;#[3�r���jm�]
�b �Әj�n�ep�/�ɓF�hn,��q����E)�ˈ��fQ��4��2O�s�ŏ����7Y�m	�Q�Q�C�����7�^-΢��N�#�l�6u��
�b�[��� �G�����z�^�_�����g�������,����\B0�4U5AC�J�ݪ
�fpo��=�a2o��E�A9����;��b��Z�д*'2��S9�ϟ����%;��ח�)`g�XΌ��R�.�f�i:���QR̎�� m�B��K�<��q���ȴD)��_>뼫����"ۛUĎ+�.��*��3�Q!h����>�6dn�\������=�k����Eo�ޡ���P_<�z�ۄY'�U��9O��o�j6�L��{4��W�E�\i�^�5�`3j���M����J�S�baT�|3�@�؈b��xѰ�T��:���k���}�u
-K���Y�:�o,����՜��y�MN��[*�K�
±:����@��vb��Dr����yX;Ky��gt*��"�V;�^�hQ������x����E:u�ێ�ö&�q,͔��D���m4�)O7M���C|c��t�
�
5�y6�:�W��˝M&q�%J�]:8�Gw�LW�"R4�XC1l���(��6��R=����Hy�B�t3b�Xr�ev;ķ)4��؎�J�ʲ�x��un�osTD躥Ɇn��Er{Gh]@�:�i���ҏ;D1����k�;�Y����1Rl��j4��ې����f�0�lޖ��v��-ַ���JNq����i<�#nv"�0]��R�p�5�eʝ�����r�t3�ڷE�7�k��0r�q�ʦlh�����i>Ż�u؍�F���B����sn,�Å�iU����5bOB������ ��[��u�f�ǭ!�{
����
����][��9Zq���8���SԎ�}� y�y�����<W�SQ��¦EO^>�)mg�'Z�ۗ�������y|_̵���\Zz=�[/"JBi�]�ő�"���'A�u�ׄ�L��A7|%�)E]�Ƶ�'C��c��ɤ�b�`]�&4��ݍ1\�����n��tU�K� k�h��=��*$.���V��/6	�2]��Z�D6܀���캺����#�3g�2H�ⴆL}.{7��'k��C�p���fH�����vM$H��mѷt6��=�Smb��y��-�D��i��iT��;�I��m���qtj��fv�ފ"qlɷ�ۆ�oGRgU��[�j\Q��Yf7g�R̹�:89���:J�������V�&�%P�{2��uCe���&^�=��Cu�;���6�M{L�&���&k�d�	��Sm�Q�tqr\Q�UN��Dʛ�\�n��p�l�%ZWJ�;��4���;�(�����^nVր�쩘9+���+�镼N�nO�ڎ
�ަ��P�����y�ۨi����VV,Ǡ��܈ҹ�Kw"�L�.�,�3&��MwM��#l�Ԃ%C-���o�Ǘ�`ñ@�.�.����MM=�V�&T�Ȝ�4A\z��n��+k��|؉�}����bGC��<�EE:I�<�1E)*Ti�B�n�2�1���#�lbv��6��m���UF��m�Jm���lb(���Z�֬clF�5CZ+MPcgF���M���kY��#G�CPDCITD����b�t`�U.$���V�kMkEiӬE��ۭb��;Z�БEj�3I֪��1��Q��n��睝�N�T��;g]�MRv��l�<�k�y���y�ѣl5�cWy��y����m�FֵF"��u����mۊ$���.��GM;N���Ub�mj�m:�����QAbo;��k�yb�t��훶�Ɗb(�N3lFM�&z�#V6��8�J�6#T1���4��]��)"��`6��6�cU���m��Rִmc7Ӹ)/'^w.����=�w ⤕/�߆��lp�(�y�y}�.�,�����(��[��;}�4]��z\�ۜ��#��U֤�:x%t��{�1$�F��� UfX��#u����R#@4@x���Dт���W��F"fW�w��}��t��l��	ޙL�O����y6�lQ�����1��A�@���W��J�	ط��U�l������2�m�6�rB�
~��!&��5�)-��<�4Ԥ[>�p�լl��j�h�~�/&�)�
�%�o:6`=��L8�i`�H�WC����NvQ9�hw�|~��>*5��f��,2��X��>H)���ܬ�;k�m�����s���+$���	ڐaiT7��	�Trr�;�Ih�ڢڽ���ş8A����we?�|��~k�T��vDG1��L���4Z��jU-V�Z���s��s���Y�F�c7�7���և+]\")�?p���!�z�!�"���ib�����$����@gciiި�0�n�Y��|���8��[Y�' �+Q��:��1Ø+�H.�ƭR!GW��F@���ʫ5��U�p�C뭈,�6J�r��B@¾6<���)i�����bf�p���^�aʹ_�\��*�[��SmFj�$��t�ƮKwHZѨ�pQ�fF��jG"�X�-5�Bw��"w���qMQ�4Ts<��yB�1�xV�˒��z��!n�{1
}�=��]h��ґܧ��:+�R�Ԯ���V�����W��g{�9�������DO��U��5��^�	�ӻs�ۤssB�)=T�ev�c�$%�|���9!fcwsř����~� P(R�(QJ� �<<�o0�I���a�͵�����p�7�q(��@�\
�G�'E��1�7�U��~O��Y��f�W��mN��������j����"����x�kI_��\'�l���	_@*�Qj]�Wɯ���, �[m�xotE��mtW�_d�@�E���D�j�v�%�}������_�)}��xg��N��Ly��&<�3�q5.2&�S���u3�7�bM�d��[[��t�����l�w���,P�����a<ɯ;j���t��2��i�+S�퍸+lncͩ�׋u�%��b�M�)�{kml��L�H^�ք���#w�v��e���+�d��u!|M0X�
2�S�T�9OI��/k�*�kP&�%����MD-�ެ�+Z�46�ٛr��*l���4�,��gm⤷���Q_7J�/��w �E���s�낎Ųr�23]��pt�����E3�Ƨj�S��9(�����}1���r�Qر����)��e�R]⨈1��2�S�ǩyN[�\A|�2)�~.SI{(��L=��-��8�^�����,{����޺��t"Ǫ�*��5Aʹ_<�N�ԥ�u|�Zu �t����/>��5���8��x�-9]���s��:�W��s�f��A}|\}GQ�G2=x�w0u�[vX�%�Տ*l� ���Vo`t�;$ꜜy��yV`�������y������*�,��x ���0������A��i�0�|�.�W�#ϐ��A��i�D�0�E��K�:/~����"���L9+����K�~��5fU�4`m���_c��k�l��?�#k��Km�9[�Ly��֊Q�_GBA�adɪ���i���qϏ���&u7�]�FV8j���[�AZ�j �`�4�^$\*��}z*��ဝ)����W���+�m����Ϸx�-nkhp.i�F����UB��G�:W�k)�7N�YK{-�l`ץVH$���e�풣(�ۋ@C��˪Ok&$^8Oz�*[��`-i+����p���EUZ�6��S���&(ݰf�/��'55��E<1��}Ї&���\�
=���U*��'�M|����pzV�������ǏߋE�U�j���z&��2�ûΖCؾ<���wU�B�ұH���nݛ�+��G�h{�L^���;�Y�tZZ�fv��\���K�Ƚ,�/�����gE�X铍�t{d��s�.��b]�Ԕ]W�5�w[��V٣��m���F�Mscg:d^�E���{~J.Йk�"�I�z>�U5s�|vZ��!A>�5]�[p�Z/�Vr�{e�5%��t���o&�Hz�u�N���5��ѣ����:����2��)��\�%Zk�ȱ�ҟ1���Jx_4q�tV_v��ܶ��VIY"�]I�jw<�vO꪿�>���H�	�"L%2��yD,�2a	p�ʚ�q���4{o�Y5��M�)?[��Vױ��6�9F���dd���Ulgq!��o�d��A~�6�d3o(E���N��1�������[Q5�OhQ_�=����Vώ�q�
�{Q=��t�򟖊��P&ƥ1OkSڜ��n���L�j��AD��*V8�Q��b6� ��e�t`����|;�_W�R�Άh����e����n6ᦗ���l�a`�%�
~ϐ�蟎�Q5�/�Z:P#OH�c4�o��W���)�{����R�
z��ar�Y�N{y���Y�V�b �:�U�( `k.do�"��}�~��Q.�c���E2��-�$걸
�1�a>4DA��j+3�>�Aך���DB�ǐ��ef`S��.� l6ᕙع�I�ўi�5�/��lo=�c���Ʃ�����0Jv-��ۯI���0&�8dm2�p������Ț*�]s�|fE\��+J]��F��h�i��m�j]pbxoLY���PYn&+�7��c�nj�(�}�"Ѵ�j�� �����l��ښ2�<h��y�s2��YBD�S(>��T��t�be���)�mԽ�sNX���ANG�����U4�NPY��r�!¿#��1�������y�]kR��[�r��OA��fl��;3��I���F�����pɺ�=�o������"R�D�
=�| >� H�q/-�m�r���A��)�r�9�($%��%)�!�\�����ۚm!�5o0�<4�4���[�t��|t��=m�B�v�ׯ�a�}�88y�_E$��"�쎽��r������6�L��� �8������:�>��e^;�M�y�L��d���pVؽ=������]�Ƀ����w>��	�4ŗd[L8����ݚ�j
m���Y?_��2�k{J��DU��ubk(FܞZ�c�{x����L��
&��:K덁�S�eav|�l>�A��Z�s>n55a�Ř�D�jAvV0�ƕL 	�[	Qk�tj��m���zC��j^+��L�Va�vu��I�za���s�׃P6�)t�דN�R;�R���5���r)��؝%]d_KQ�f�7S�m���s�2K�b��Efo�ǻ��a���X��>H)��ٛ���|e\�ԣpݴsKP)����s�(�oP�v�P⫓ڈ%�'����-��jē m����х�"��o5YX^�H�[%	x�	���[gp�l�>J���ƺ�J5��``��j�ma�1m�E��絵���7��L(�ʎ�pd1�S�4�M����,u�ݱ6��W}L].��%�@+�P�-IygTcTZ��;T�Μl�Cp�Z5�J�ks��;-�W���*X�˾�w]S�tЩ��Il��㫆���y��Ϸϟ_�ǟo��v��(��>> �@ ��A _dc|����Ph|R|�^9�M�����:xյ��J����+��3v��:/7��"e�\�q�G m�@���3,��'۵18�T���03�U��T K�suV�k��{�&���Da���r������&t��m!�+�a�	-Z�R4��wv7������w�h�oCa�>X�iFv@���U� �-$k(&&�-,a��Iv���F2���sC�u��vdg,�	n[��k#xH�)M�	k��C-����wYhS���w)�n[�h0�{e��)�	��Y`d��^eT�n�h����,��u,zj>���"/��E%-F7/��9*zҍ��=����"���Ձ>����^Z��B��'�Ϥڎ�x5�(�T�v��S�)nN;_����e'[jǐ\la9߂�x�~hqy5#��­k΄5�Lf�ud�^t֥Ʈ�s[RյM���V��w��[��!���"'���(	���;a�e�%ص�6�T����"���u�b����0�O�+�A��Q[�f�E[#����Y%'y#Dz&/$�N��]KVMgb�g��}7Rw]QN��8ܓ&�n�E1�b������pr���.l�X�s��L�S��������+&2�)�̮>SM�Ǘ����\�]��>,��II�wJ��'Z�F��M�:]�6)FX��:d�u�e��3�_W�|RLJR� D�������������4�n���$�/
N� �Z~8����E�ݗjQ��?�d��6g:��2��nq?`�s���W	�u����b*,:�/����,YC�@���
!�K�+���#(�)�-�W��n���p��Ǎ�&G'9��l�j���l]2J���#�4��˱����`��X�S!I.=��4�{q�Vb���f�\���Y�.r�4��-8`���Q=]ת멪��A��ym���T[ZH�V-l!ۛ5C��j�Q��>l	�3p�a7j�3oM�7��V��䤳���j���辰+��`�����=�%��a1j��&e�#�B��ڼ
'!h�_R7~n2���7<��[P:FM�ׯn��i ᤉ�^$_fc�ٖ���Sp�p�`8��X���_E��ëb�`�P��u��ZѨPc�֨��^��{��cr�H���p:�)`��z��û��[>���k�Y`�ԝ�P�t�Y)���5T��2[.]�jG�s{2&�AX���W	��*�����Nr���T��.�4�������#*N�3|!��S��^�Mu�n^N��c	�F�㎤�'��^�뜹�)p7��7��|)�C��޹����l�Y�uH��^Z��l��̾Et�N]�i�`�6�$x����wr�� ��L�,8&]+�'^J�ג���46���3/d�z�^%�*6��U�}��UQ ��A �@ �]�ob~��j\s��|��� ��dZ� �\KSo+�Rc�,1MlC����]��քj�!սmn!kd:[��T���7#�ע=`��f�\�S��r[d!*i41yj
��r�rE����[kA�EdQ}���ʵ�5-ɘ���˩��x����Ī0�NhB\�J4�2Sj�u�;�L�03�b��y���W��hF�"i#{f}�=l�=�S�X��e�M:�� �4�W��&ܳF�&�[ �VX12�����q��D���٘�^��X��'������vQ��yjB�`j��*�ȧfӹʔ���T��x�s��.V�An���uo�����������!@L�]���փ��z���a�Xe0��#�)7p�1�sn�mD�֭u�����+w5Ju��d��"����<�y�q�P)>)�ru���j]q�UnD_[�Y���z������D��y�g1�����E2B�c�g+X^8���V�<��W«*��Q����]J�=n�8�k�*Fs�e�Z�� �pEy%���7�L�&��3(��0�B&���ަ�o���W�6wSA�qIr�8��b����U�P�v����X�Ip��E���5���<��yQ��i�^v���$\����77��1��V���źZ4�1|I��$�څӱb��-��6m굇�K ��T�yţi�c�DL̰C�7��d�Φ\��X3|��S0���St���'���EydsEѪ�֠	�g/B�����ԱL�k�u�&yn�N6�{!NO����[��~�k�S�z~�ሕeI|�y����o�K�'v�<Htr��+U�N���ڵ8tyQ�'s��fegE3�Gm9K�B�7w�]�L��u��{���r�G���[޶5�E���z�<[�)�mA2�x��]�iHf�Iun�y8G6�V������0c��^J���tc����5���Yŝ{Y�&���a���Q�����=6�u�w7q�<�<��j�#Y#u!3���hu�'�}��e̩��B.:ހ�,�39��q�D2+4?���M�K��}E��K�"��5j1���Nn�KI+ؠ�Ye��# �~a�����_�������[5�t���z�g�?-b8c��Y���º�2yT�b&��2��t��kd�,(oL�]����H�
L�eC<���L������fcH�Q,¦�G$h��L�۰�ؠ`��\k�E|�D(y���GZ5������^4�΋\�p�G�>���W[V����e=����}�6�ۛ[�)[���XƸ��"sw*��E�����qu��top���vU`��bBMDd��b�XH�!��Ïn0>�<���"�}M
{�顊qS?�U(}��L8t�4^���(��L,aWE����E�v}K���Ơh]�������Bn)���ڥ�35u���S%�����%�yS���"��X��IJ��nAhV��d�������ͼ2�0>�Q=Ö@I�O��ˬ�7����T�s�K�O���8�nk˻������������*5�M�8fl7��ʦ�d�5x��t׎7TRQ��aC��p�T����U�)�Fug
yv8N�j�O��:�B�l��kٜ��;��_Y|]b8��_3y���y�UE��N�F��0��Df�Lm�T:8�TQ��|���څ�����5�����V�Č�c=�"2�jk�M�;��pv�3�׀Aa0��	
0����P!YX�K�/yx�q����.5s�N�įw P�םP��C�fF�bi�6�3Fs��1�m�M�p�vr?#+���S)q��f���������;n݁��e�H"~ٞPY�r��Y��S�w�eY�_l+O�������&p}3�x�w�hϠ��$Iq}%�^[����z=~�W������~C�����0�w$�P�ea�d-����h1e�V^l��C���c�i�.�\b��"��SXT�@���ݫ���\ͥΏ��mC]�@A��fm_XQ�mc�	��ss9�[�]�k�^?�PQ�vfB�Tΰ�8S)gt�sfPo��a.6"H%d�	D)�p�ЭF���)g=��w�M��������=/��a (ւ,��I���.��}�e���C�Xl��ՌL^H���]ռ?n�7U�ݧ�\3E�li)�HF����.����N�ݕwʗ�G��0�;9є\���w�
n�_]�e̥�b�2�v���n",��4�ջ�6�Ҷd���2e`*.�Xs�(˖�6�����'5���]�h����Tͥ4vr�j�saKNqvb�7�k�cwz�\��Σ�)N�U� ��R�y��]�Af���+�Wm�v�Y���O5�j�2�;,rݍ��Ψ�޴���K׍WFs0
���%=����Ib�P�.�S��*6w�б��6�K�]:فŮ�Wk��.֤���=9�w*ݤwN:�����3���V��h�:�S�\�[ʝ^q�V�E�䇰a�������-'s�<*1Օ�yx쬦���t<������d����*0p��k��r��%7���G�\֢����$U'Xgv4��E}x���Z�S9�bwL�2�F��4rh�ǄΔ0N;�2�z�V�\J]d+؞oȣ��*�;�3�m\�\����������A9ۛݡ���`�8C�d��K+��Q�6�1�7tn��k�2�ř���NU����
ɝ̄��741�s��>[��v�ћ��{Gk�8��\݃�m2�^��Te1���Ҷ�\��Kp�E;�n��v�)D��<jjDQ��dm�ɼ�v�I��ۺR��{���lo4�������e5�:���k�����v%�6��K���z��2����GV�K���,���e�^+����`�V�Rfa��$s���ǝ+!�#�Z> �
æ�p͏�b3��Ӷh�V��J�"n�����\�CײS��Gj�3�<j�YE��ƔƓ|N!j�v�D�G�f�sV�M��V[�ڛ�fe���ڸA��Z[4���u���H��ަ�(�й��x�We��6�@�96WN�.�If���oe�tm�i윤{��6����͑n!����r3�:�B'0WAK��*�
�zG#n��6�ƭ���ʋM1s	6�v�yY�F����"���_h�p��K]H��R��.E7{q�rѴ��j�:[`��N�9j�������uϠ�B���L9&�;v42V$��	�*T���iDr��U�� �ܹStvͺŸbk�/]�Y�D���ܾ�W�N���-�� �%R���;14�k��R��E���/d`�c�&o���&�w�tɎk#��f����Rưؘ�el��D���1G�$#Y؊��6��tb61F��sţm���U!��Wk֝F�X�/;����*�b�s�b�D�1G�h���;/�M���Ƌ�SUE͢<�Qu����"*��m�c`�/h:�#O�H�k��
**)��lѪأU[y�*{`�Uj1G�jj6:�x���]�ch�<A��̾G�]���j<��#Z�'n:-��7q�b�ح�8ѻ��"kͼ����󵱨��1�
(�5�1Ky��lF؍�i��"��)���b�)�u�#�z*b"�g5�y�y���^�[��*
�[8���vq�i�ڭ�S���G��d�5��5[�[Y�q�h��E[u��J`�����*_'L�1^F`���j����SA'����m�3TΌ;n�<��b��� ����+��ӯ+\�|�g�FV�͋{5h<�U��u�1���q�\��̘�0MPd5�����{��kפ�Ԟ9r��	n��װ��D\|^���mW6Ýj��{�2x���2}�n���	��^��ĳ��,1[N��ҙ�%<��R;�"@jqj`qy�ʺ�<,}�8V�&�qߑsTf�=��n�͚�sq��3<��d� ";ғ.ˊ�l����S�H�`�S.k����ݤ7v�.�i�ފN��yJ�W8�Q�U�f�<�#��jt���s�Y�\�X�Nؼ��u�a�e�����M'�TY~�-Q�{aU[j�r�\��1N�#�m��͊͐����1����VL����b��/7�Y�"���|W���(u����LA̺l�v��Wc�����t۪h8d��nq:/Y��}�ݫ��z�YՒ;���rT�Dv%��D�iIvX7�!��B:-���~Y���Fs9�̮_-̎�⮃��� ��?}��m����hJ��Fݚ����76j���j�!F%Ơ���d�h�Vs/��z"�l�Ij��lb�gN�c�\�u��RW�k(59%�6����s��L%6]�w�,���A�#��5MY���;yV'��
��L����q*�os1N�^b7]p�KV�I4�FJ۹��)��l�-��{�:�J�F��]4	�R�W��e�gp�oi���%v	m ��N���X���Z�/ �ah�ˮ�����>��g5�{��B6 ���d�C�9�N7
41�,���SZ��cZ�D,&���}A�"�OBsH�D����q�Hu�����)j�5�FW���[���6����O\�-�e��˦oam�sy����"IMi4w�j�^��N�p��E94v��ՙ[��SV%�rh��Z�ǣ���k.߬�撩@��^�Ѯi�w�r����a{MSØm�P/]���xn�t�2�tĉ���ϭ�v�|o}1�)�o��'��N��z~�u�,7_�9*̌�&Fz��^+m�z��e��N�c/|�|�Luҥ��,w�U�73�n���	�U�w����w^[6�uGc�:��dR}��Э�8�[|�E�DG���C����? �����5�B�׋ܹ�(�j�❬��Ϧ�b���lR~�[B��%_s���l�����in���1��j5�i�t��N�K�"E�j�8ū��F�t�O��ț�b��������ފ5��n-�@��e�� ����T�δ�a������ߏ���z�ԥ��������Ѻ�-c{�C�v�c[W�����[[�d�s�t�?��>/�p;i�<Ҏ�>��}���.��W>��Q&��8�x�1����a���L�#}qA�fg�� k//je����L�x��]�{2�Yd��s��0^�����y����y��0������;���Ͽ ��u{�厱1[#����DF4��b��A�P)?'���
�9�i���k��u�ְ91����׍l&���|�"YҦ�R��̯�F��ߎ�M|u�r��d-S�P����H�#qBͪ�⌖��H�L��
�?�%�0�q���f�͎6���37K*e����g�|3�
�*�8�����#���{�xW�0[
����� ��}
�M
x_��OySw(혶a��69oa'U��I�{��֋��mf{#m4ǧ����.b�g�k06��ۈv
��K���ѧ�Z�L!��7���:�v F[dX�AUN3lG��1�-��Lk�p�����dC3�v�it.]H�2�ܫ�w�qW��T�+x帽*}�I-���r�@�3y�ZԽtk�nj�(<S�*��Qd�)u0������L�|I��hT(�D�j:��f�hq���y ���ʀ�ek��͸4�Fɠ��c�TS��8�;us,�#P�ڦֱ��s�Jm�BD�xj�H'�D?�3I��B��Idkg)��s���*��4�<��WG��⼫S��)�;���/~�!#��`j�[�V�nf`F6(��g���/����2����LT�|W��v>q�#���^��sc���3JA{|��W݃V�sNb�z�k��f�:?������N{����>eQ��{,G��{k�ٍ���N9��VP�{խ"�^ۈ��b�n�W1�I�G�&�!K	��<T��V�U��M�3輎�43����x;|��9���*\�舖��p�M��WUH�wP�Q�Z�%RL`�G9)�q�����g��ym���W�0em�G=ޭk��e�u)�z*���Q��.�&��˥�P�8�=c�����:���-�w"Cݠ����"U��o	�[m,�<�&-�$C{ͬ,��i-�Y&�:��uN���-�f�ƴ������.,�*)��"��j~h�%'Y*C<��h�j<E�T����H�N/?c�rR��BL,_����xnC�1��oOa���Y��K��s8�Q|�p�B�2�M�Iͪ5w�j(��-2�#���y C��T]�铚��P5�$��ئ�S�g�⒩��J:1����W*~tUm�{�C��e��J�X���K�-���5g�A��-������i�Vv���D"�G4�#��bp��5�>ua�PlU��(�d{��p&�r8�$04S0�II�¿4�s�a���U@N�k���qk���
;3_U��M@jY�K�SK:z�G��.�Z�����9Y��5yb�YutŤTc3���ՙX/��5b�m�S�Y����ʟnָ�F���'�j��}������1ώ�l~��?,��*w*}��n���Ѝ�H����fV��c-�n�S�hɪL�j���9�������o�:K����]��0U����U\�E-�#y�7�z����Y��C�l�,y瞋[�b�5�Yr�q�v�c ��D���p��5N���9���۟�m3u%���r��~n�Ψ�Ч�Ws.f�\��m�9��U]c%eG1���y=�V*��<�:�����T�4�V��q{�U�b�}�Mz�|e��ԗ�n�����f�^�+��r��]}[�U���qVҙ�%:�2�N.C.6i�T����ʺcK&;U\�vZ�4V��5n9؍̋�&Įe�J�֙��{I��@�3�&F�
K#kf�~�w�sJZ�U�D�>����·�����)?^)O����=�*vMZG�/.���ňvV���`�)��"qߙJR�ջ$4�a7ҩS��J��`����]B��U�֠M�K�k�آ�34��KX�w���C��/�꺖�[s��}�������^�J�K��a�L�A��,���f*���^��_������B^U%��TO�u���#���˼�����Xf���^6��)����]ػ?7h�mAi�ʹ+�����{��FKp(�O���T�l�ܑ"MZḛ\3.���/ L���n��S]w�Nw��}U�/v_z�����o�U�v��@�����/���a�ɧ�y�N��-��nQu"�Tl-����"���+�]�me�{�7jF�v�b��.��lM���,ۇ���8���;�T?�V4r����l�����g��}]ݯ�����x4%X�$n�5���t�_����U��/3�!d5K��-۫��.�����؞�͟\��h�m�������k
s����e�Mj,��ч�^㊊�='��4#A3��ߊ�׊�>PUU�@���Z�����lt�֕M]xҝ�.��N��Z>F�^u�>����}���-�6��`��[N���S��ۯ'���&�������14vc*=�f�'��I���I���}���c����������mIZ�U�2m�n!&�`�?�
t�������q�aM�뵲�}w�$�mu�;I�44���S���.�cx�3�Oiq-M��QHIʀ��V�����ƢĪnSHi�3.�`�0�?��C���I�|�ɋ��ve�%�Wqq$y�������m������ǆ�k���^���Ǡy"�����e�/u�����8�Vd�+�ohzj��U8����F*�fwV)��6%(�Z�Go�,��5v���z���C�1{B͚�\��5��|������>����J*s��n�
)�?���U&d�oL�|v`L���똦4��~�A��dQ}��Э�U�)�-�xy�T>��bsf^1v����W
د3�O�6Y��|���1)��wBd^��7�u���<�P�l[�_��?\�b���E��~�F�Zz>x�Z��(L-'��æ1�cL�L���O�fL�����h���n�g�0���P;6�R2� �԰`+y�(����h�s��[�R{���I�F�2��`�O<��5?yc��>��v.C��;a�0�&jtCsؠ��)-ŷ��ơϓ>?��m��/����Z�&9T�)��*S.�Rm!Bɀ���g�(���+�������ػ�/�{��l���4렌Rz�+�T;q;>��!����pM�4�*�{��!D�^Ȱr�S�WO�1�/Y�_����0��v�6,�*\a����dw8�*K	Z��ʚ1�^7VP��^�o#��K��j���\۪<��\ب�S���-�VȾJz.+�#��gy���ÕtKFU�t����j��p�A�p�L�\!k��
��	x<v:0�֋@�r�ݭvO*�̭�L]�$!�n�{Sk�j[���{������Sw�!� 	S��+�R��Rܨ:�,$�]\�W^��t��)�Q�ٽ�nY�M�]�p��J�N�T٬�����g����]�I�t�@��d�J}�r�L��=�S��x���#xg�q��I6�OG�����c�{�?����0�C���	�N��e��=�jbyY/1���l��0��#0-�:�W�,���iN;Xi/��<d-�)tk9V�7�V�h~z�.v��D�%������k��r8�MS�^qv��b����x�"��)�>Fi�t����"[V:~�)N�چW�0n�F�|I���0+�Qg"���nݴ��0��P�$M��X���v�"	����y�z~�t���)�p�W�L��4a��x9o��Z��K$��YB�ЃK��+�"B����Gg����P�JL���e��g�P
��5��:��߸̲~��B0с�JM�H�NM)t;��s����T��L�ҩ+��R&�S�f�ƃ=ld���2(C���-��%�f�`�L�.�US.s�j�m��+PJ/"z�KBTX^ˣP��Qv�p�p������e ��r��*�iY��^S�UIn��&���H}yeF5	.�J��V�k������p���q�C���댢�b�qy1 Q|d��|���F����+���47�斀���˛Y�	7]7��4+�aɺ3���h�m
�]�d���+|�͕�:�][�c�y\��Yʴ����+6�L�u��ɽ�]�'�������=fF�ms�5U���>�C����[`��ث-H���F��b�i�|�[���}�_�v��%��U�rޠRy#��/~1��Q#��gM�Z�Ŧ�:±�Q�d餗 q�� ��66����D;�]GN�'{��+[Qj&%��pT>b���TX��)�����:9Z���n(f0L6j�:{\c��.-�"L�sV���?u�9y׊�[J��#�ȋ07M:;�:���#�n���Z�xž��mE��Ɯ�݀ѨoC8�q�J��F�|�3�z9�)�l4y�e�Z`V)k�9L86�"q�i{��P��Ƥ��|��#`���v�S�hu25����;"�f�Ә��YN�;���}��|W�=��R��N�4�X�z��Э֢M>�d�Xf�n�6o"��%X�0-Ќ���ϱ�zڟ�.��Q�d�Ȧ:�����=5�����D9�+�oJ->�~�u5�$�uϬ9�qs��՟Xt^��ǃ'~�*������|e8��eA]��~sɌ+SE���}�u׸��&ׅ�����������m)��BS��AwH9���^����8h��j�$���B���%���r]/:��]y|:/.��بEl���Jջ�F���
�N���)�ާ&sZ�F-��`�2`lԜ-9{�)��t�_.�wr4T�v�Hŭ�:z�b�ɜ�R��V���μ�o�Y��*���&*�߯�fv��*,����3'�~�ؕj}��L�Mv���i/�oI1y@���%&\츩�S���gdd�ld�MH(	�_l�����}�I�~F)9^E�}��>9��h�]^#ևN����W=�8\ki��ͣ{�&�j""!yytk�j��m���y�:�\q�T�]�*u9W�q��"�Ȯ�,�b2�����Œ�k���0SQ_����s[Kc4�l��<6�JSPQ �%)�n3d��y�n��+7'coS��2�Ӥ�(�C�����Hl:�?jr��Lx�����t90*Ɇ�{�LC��O��)k3u®�&�n4�v�Q��ڝ�,�$���.[�b�:~Y�T\ŝ2-K��!��gd��:�-�!��Te�*j{(�e���	V*I�k��!��Vt�J�|��f�����|.���u�zO=%P��oGr+�
�V�i��1��J����)��ie���~}���� s���������6玵�;��=!��ξ���b6҈u��H6I%��H�]�����=M���������cN��d�� o�����x��>�O����{�������Kfшַ��;e=Ňܔ`�UfN�)�F�`%�ݮ]xD�N�����l��~�sFݐeI��Q�4jKOp'e�Ǵf��Ŏ�зxP�#2�NM����.�([Y�b�ݓJ�B���T.�|~��Do/���:��q=�4\w�nQ���6]��'T	�kqj��𳂰wd�!����Cef^	��EDNS��D2��ε�:8y!�/����xj:"�`b��-P�P�ܾ*)��e��*��q���X�s�r�:�wpD �
��=�4^rʽ]�aJ�E�� �	J����uݛ��c׏j���p^p3��A-s�g:V����9o�m��E�.��)wV�%؝��<�Rb8��_i�
B��eD�d�u�s�'.x�v7Z�f�*��x̙o���j�/���Yn��Y�┺�h�O�m��]E�zh[g2��uZ\�v�V�����f�L%Q�֫4�H9�u˩��Z���d����4��̦��R5շq�X��<��Ѡ"�i��EYgM���k�[�a���Hg9<�hJv���X5y7�*v��U��I|�ೠ��U	\�JP���^���	�O�q�J�2n�u���p-�A�::\�f�lT'�;���L�K�op<�Ү�e���nā�h�*eBҘX��J�n]�gq�a=�)a�*^u$�h�#D�]��w�{�n�u�����]������\��A�:��[D�ɍ�q3u����Z��jSsU�{LQ���]����0���[Ɯ�dc�e��n��Cy��1V��J��Y�[y�N9pZ��g4���'s�8i�N���Ԇ
0y��f���ɹzv�fԥE��V�T�W��`�y�L����P.���5�������CT��xFX�(qH%nv��c���ʢ�e�v�g7L�qhy��!Ījĥ�[F�W=-�o��J��ɵ�Ӝ6��ϋ��f�V�(Q�ս�u���%�Jj��㴌:�h�{�= P��e�:��|�+i�xMr,=A?`��*�>�
I�!�0w�����	�m*�oP���˚�VM�
[@�j��?���p**��ge�yy�����>�RܗYJ>��EݙYW��۵}$�o4WJ���ʗ�QNY�\�y��57�f;vpK#�C9�<��p�R��IMv0��ӵ��xZ�)ܲ��Ԕ�F�Yx���k$�@� �f%���7��99[;5ՈR��GS��َ��*���k5*V�]E�K;:��������K;U��D���.��4�dGܫ[F�1ܻ�]+ l���O���o�)�+�탊*F�)4l#�V4o^���8U7N�Wvl o����u�ɚ�-���s�W���%1N��a��S3U��˅�R%�Grq�i��\帖�ڳU�K�]H	��@Y�z (iI��"��N9��H�D�@
�k6ݱlڶ���Ѣ�-���`��>OGT���5����b�����H���1G���^F)�"��:����3<mT���N6�W�Mu��h�]�6�w&��֪61�S]�WlE�cXb����ƫc�{Z��t�gi�j*�1!EQu����F��:�;TDZ�u�(��kc]��l��{�Z�n����5QIDGy�1��u]�Z��"���X����(c�Fڊ�,U]b��(�ق`*��E5�Qӂ����]�PUU2w��N��R^I�*
Ѣ&Jk�&���^mUAy��;b���ճ���F��Eb�z������cuݨ۸�:8�*+F$�f��&�:���ͭb.Κ�[b�J�������UA�".Ɉ���qص��q;�5PUQ�h"�ֈ)���t�&*�o-^y� ��)`y�A<@�
5=NJ�u�S$�M��s̚�2 �K\ћ����[>��6�X�R�!��\I�YC��w%�8�0
y�}�f0�d�v�kw=��v�*WǱ:W�jV�E�[N(p銬�v�47g�}Ƶߋ-c��������Gq�/�<���P1:W����V�v�(3���"���	�h�;�:tf;;Pa���(�g�6�r$����ք���o����8S�&�y���S%��g���e'wj�3PS.)�W&/ܾ�a�~W)���2���e�
����~�
�3��/~���)sw��!}p2_i��*m�P��R�r+���p�:(�;�N�.�j�zVP�k����-�����XΔ@��O�ʝn�xMm^��:ה�ض��S�r�VT`��ѯW{��q4��@-'ײZ�[�ȉ:K\tQӖﱦSs��ܺ-(�\z�Y���59��a�V��2��/��t��b ��e+h=�)Ƃ��� (�> ؙ�����A~�&8�P����x�N�'�n�8S�Vj�����mk����<{-4e0:�$4n��~
�x:{t-'��VU�f������9�o7J��̉U��@��=��i����8&,�]�/���82&�R��T��7�:r��J>�S4E*�UJ��:�e���0.�T͘��p~1h=�p�6�9���H.
{o��0��E�F�:	������*�8̕����f[�6r�2�S=�H����rĹ}�-��J�5��ۛ]8��Q-�*�=��x��y�c�y�ZEW�q@Y��"w���ִ������E*p�l��a&�/�Q;N�Y��2ɇNZ�`�6*=���6,�*\e��.��;�e�T�	E�nu[����������i �`G�H'A�P_-t�{�ޠI�cq)1��٬��T��q�ؾD(�]���L{1���G��遲���E�_
j���Un�����c�ɓ٥��ԠL�f��Hp�k2�ݱ��@؆})l�G`coS�6�sp�,5j�S�	�=�H����eV�h
�PX�Z=�´,��+
�f��\oDq���.���Z�f���k���c
���z&j���(,�t8<[߯Z�#�2�Ws!��cV��B�}'ać�$�r�vV�C��:Z;N�n���62�۹�;��Y_Yr]mf�{��Y�؞X��f��2��~5�4P��H)s��ya��ۻ�l��d[2�x�Gk�5Po�X9�M6��)���r�O�l`�}���J�|7��1�f���L�Y(o���ō���vWNL/����5���u��2'ŧzUcM�[5�}�m~m�{��
Z���
R�)��%ImQ��[����-\�!��iʖ�e�Y���E�7�ٲ��	2�Pͬ*�Gm�y�uc�x���XҀ����p�ڮN��f����t�g���������.��#���z��[%k^g�����Z�}V7��5өV)J]��D��!�{�(4��$��N��^��M�˲	��,�ˬ��I�j�mYsl1(��x˥��Q��F�u��<�D�d��z�'A������.]�:a�T�ܡ��G$V>��v���u�����hS�4��m��e::a�ӎ)�����`�(����ሤ�ת9�����Qbؖ�j���z�k�y{� ��C1Z��T��+-���L{r��+u������	}V�w'�"J�ÚcmO"P�X7ZN�'����+m�M�?�����ED�+�Lܾ�T��gA�v�&�6+BP�� 5L	r�)L���]���7��X,�!�5Pt��ç6@��G�v6�9�v�\y����U2ԧ����%TuG���{5��N�Ʊ�0�sX(���rKz����U��h���^��zO>v�n��N޺&�q���KMy���r�����-�br��J���of�q���rzB��ke��)%���{V�>�GּG@��Hl/2/�y=�RTh�"ʓ�cӦ�No:���B�#�v@%ed�sCb����j���A�e�*\��fo@���
��;��T���K������G9�E�rR�dY&A�M����^�]�g��ղ>�l���RT��푎��o9C�u�1�^�E7��^���o�#��l	c/K��`Dx�·��{�ˁE����'k�4��ƅ���:��B̵w2fɱ���K]Ԯ�+$�PT�bﭼ����?pٙ&�����~��P�ӗ�Ɍz��]������%�6�.�8�iI�<>&
�Iv��P��ȉg�7L�X����2F�hi����e�{����k�6�����C���3?�BS��Kyž@�����]x��kn3�P��5��5�dҮ%���ڦ�KkZ}v%d�L`Z��!IJPړz5��e��nv���)z!S�* ��U�q�):.��?F��ڌǪ*`c�:�d�s��кN�Jml�nFw�yzy�)1缗m����{��0��(���j�.~*,��^�m�ly��s�!�����s��-�.B�+8�����	oM�\^wF��QC�ٓ�l�;��{��9gu�4zX��Z���:[�;)�1��x\�.@�8��3����|���^o���n1��K%�<]bx�.��Lke$r������E���l��嚇�rQ7��H�h�$ŹlF�����ٞ�X��k�:3�xӗ��5�-&�à��J�¹�MW����2f~�S��ݖ�����_V'R��'T᪹����w�pY��{���9�.#2^����$�<��������Gx�v��\��ν�a7�Uq4�9�;~ɹ��"h"���ZR(�&L=�M)���u���x4%P1�*J���.l#X-��A��N�T%�θ:|[i��c�v8�L6�)�t�6=�����=��GQy}/jB�~X;�4�;�����3�xt����'���zt��.gS���5���#ƪ����:!�C�(�O�'�+�h�D��R.k�`z�ح�i�j��\���cn���3�AEY�[��Wi��4�rr��__�i���S�|�qށNMzˏ0��CuC-�ײT��[��,�T�7���PW,,�i^Hΰm~{!��Nr�y�k�a�*#7!���8>�j���~!��(,ܠg�\wL1N;^R��k��2-j뉞{g��7tԝ�"դg��G�Ⱦ5���^lԵ{W�<���BڠCVj�I>s�&/�ʖ�$�뺭Ѩ1{���u���o�{~[�)-��/�~��Gb�(Z��2���h%�(��XH��[����@�ld�OD��y�ˆ�#� $�j
�^u��Dm䞚�8�g�'1q�[�����+�t�=S<W��&�Ul���v��G�ײ���ԝE!�޹Y��� x9��[ܹ2T�yӻZ���g>z<��V��q��.��Y�5u����G#�����F=�tX��pg�srͧ
�I�Q�q��D�\i��Ӳ=
��ZnE��Z4{�[��r�I���&xgE�"��p&�����KQ�[��m&y�鱙�� ���~��������R���K�z~��4��\]����Q���R��y�&:9u�!��ޝA<&f����p�T��.R��R�Ӭ	���x�ڬ��3y1@s���#�2�>���j�ZW����o�hPm�A{���a��xԦ��5����+��œ��B�$�[\���x2���Y�g����/�#|;~�RcOX��"�4��;qf��(%��g�W1���7y���V�R�li8{S;0�ao�T�s��0���A:b��ҭ��oF�V��l��=kvD�v��[�S�$��)�FіZ�؈7������.k��|�}�c�N�O���
#�J���]���[���u���b�-1�lǷZ��z�+PT�k��q��}q,��S�΁戳����2b5�FT��ԣbL �C���7��l�k�w��[E�[<=�u>��ey
GRF���<�0�c8�a[�N��$�ވ�l�K�e�e�m�@<�Ni��T��J�V���x�f1�}Z��}p���v7�x:8�/�G�����[��+�=���=�h�dʋ������i��]�w؁�M�;=�(� yu��G�Fl'Is�&*ne�)�F����k]�IN[K�QZ�<f8�����°�|��H3�o+�m��b���uh5�@������Wl{��P��:���V&�j~fs/���������e�89f�a������P�mxr&Ҡ�v�����������HY�R;��+q�f8
s��?2��9��q�SꙦ�\��[8�M��௰�]ՙ����Zе]
׿wkH�71�%E���.��L �>)��7�S?��7dC�Q-�ت[R�mZ�^D�'6�h��tY��ު�=t�ʤ�K52B&Z��ܕ�=}qs|�9òu����
�i�˰��s������"�Q�ԭ��\�a*${���6�꫶;��C�v�
Xe[�ZۋmXF밚������4$Y�]�}15ͅO��˃��%ڴ�:c�BZ��hŤ<�4���TS�Q_[S�c�a�5c�������/̀���8���������}�s�dǃ�c���"��W'QT����P��η7ם׊ie�6W
֓f1jI���z���vhM�b�[gۊ�=��b��t:%��.+�2�:aJ�+��ZMbV�ҭ�����D�W�(s[ ��ua�k��Af	�$�nqF�S�������H-����9J��F�T��-��́��}e�W��^r�r�ZQ�ܶ*mN��yg9�yO�+��|�M�K�T��Lx��;��ks�9dlC�c��-��1CR��th����(lc��,Y��͚�:|\u�g���{����օ�#|��Z�=j������|����qnT�^7أ��]���b�87�iɢ qɹ:��=�ز�=��9�LΓA���Ū�����a�tA�~C�e>#�a����VwG��;�������T|�]�~��{��rr��
�.�^0ג�2N�́
�c����q����Z�ayzg��U�r�ӯ�P°<�a�3�5���SŚ�=sv��Q����y~�0�{{��rs�H�\�>�d����s����ÀӜ�r&u��w�jd���&鍥²��2��O��2BW���G��J�3��2�z�TȦ���.�zs{^c���Jtǫ&��:�p�V��Tv�*��<Rm[Y��R�r�sw0�[�7_KƊ�9�Z��毺R�;'�ʬJ�lx�C���B3(��w���㗎)�_^�f�`"��Nr�����Ru���!b���`4��[Hn���|�p{�b�}�(Ы�p�A'v-��ɵ�^��<��, �;=�B6=�n���o��{e�l��J��ެq�Hsz�g;�6؜C2��D�6.�z�a�%�EL u�Ho�oS\�I��Y��선�GR��WRݝ����Dh�,kk����$LԐz��6�'w*�>1Mr$y�s?��a��^6�y0nZ���2^V�/c�;�{aW\�q�OC�����c��N��:�z.#����O
��e���:w�r��F䄍�A�hm��Z]��������l>[e[>��:&Ș0:䫰�Jq�˜g]�HY�< ���H��U�$�/BX���6���<�}Y�v~�wƶ�T5���Y�u�zV�6ܴpvw܊�m�Ðɗe��6�����t�vV�*:8��c�+�]��V\3�h�j��Y�&b ��9�̀��}ϑ�`)7g�ڸ���ݙS�}��%�NP�Pl��t���1Hx��>q�'����T��ɞ�Ƞ�����zѥ�$�fĩm��z�jʞ�+u=�v%�X1�J�hj�I˩������5eG��
�VF�F�O5M��o^�9y����v�-�{7���)��Ôj-����,\��w�5F�-3;���P���L��=}#�O��l��)P�9v�]bq�Eh3p��U6����_.�k�����noL������%v�S��� ��ӛ�;��$�o�!B�h��:�97&~��7"-��M_d�����J�ټQ��$d�J��X���������^���!7�O�t$�j��ED�Kkݨ(Wxx�k�WA6�*�< �������!.��L������H����t�g4Ĵsu��z��կ
�Gmu�TQ�q�w��*�Ϫ��8�d�C&�}��"��5[�*�J�k�H/v�Ef����G5�Xε��!c-to��M�[��kܒ�)�j$���s��Ⳃ�z�^�j7����]�z���y����ad ��[Bu�h�o%C�"�;�������iB.�v�o(��/�٧H}�7t�c{J���#����= Z��}���j⻊��c-ڛ2��X���jɉ��1��$u	={l���	zg�R��kX�y{G����{<�?����zǷ����v��Zf�ƕIz�o�U�}&ei�=�9YIJ������x�nj���vpT)�N�ۓ�T6)�j�e`ר:	�����:u(8*�M���LV��Zk�(-��c�㧚C,ٛQ� �V$bؔ�9���t�����t��8-Q]���7
I���cN���Td�Ixs,�/�eP��J��2�P�L�k��I��.��U=���˾�#T��F�
6e�qPΥ�f�7D�u��dI<i^�"gR�˼ ��JS8T��M2�Xܝ;�kU/4''�<�ͫ�De�Y8��� �v���j��8�6Ou�]��ioe�S_<]<|en�9.�b���ƛ	=/�VL�R���&ف�'�s�����Z[CF[F��l_��U��7skɧ�f�m�-�G��I��m���=�ܸ�\2��n�8�*���u�bv�N�G�0D=Wr��<k�;��V��9����a�y0��Y�Ԩ�Z����`[X� ���,9
ͧ!ΰ�z(�W��W@^�et�$*��c���vњ~/6�Q,J�Js�QfrB��ҍ����kYx)��k�j*&s�qBt��VVJ{ݓV���H�����~>�Ԟzں�k�_[�G;Ȓ{Y�شл�� �S��LW��rVI��M5 ��{����۝/Fvs�8G{z�_JBu��_ݐ<�|���*�룗q̐��;3�:"Q�[ϣ��U�gۋ����MW
w'Y�؆�od�3���e��w1��c��Vc� $b3���l��:��(��d�P�JD��+)1EP]�)�&�Lm吨Sߝ�r�^Ȟ����kf�,<ϕg]�ѐo/g "�r�{g]fx�d�={��m�����SL�jEnut���b�19]o%r��}șԍ�]�;֭"�$��#F}�Ib�-K\���$;(jՓV���	^�莋��d.	+�ҷ��^R�=��tTfm�jR{6�t�����3"�q>N�i)���됚�H��P�S5� �n<]a�R#�ޮ���I�3�i1&����H��E��2�V��d�<���+����Os�%+xc�l�pv홐H+�����%�+��Uf��'"#�"��mGטq�ҳS��4������z���5��Ժ��꛸�HP��V\s��߮uI�RP�7[u��=6��g�T�WM)XӃ����b#/hӼ��MNզ�2��m��ה��	��e����-��뜞l:M]b��n������z�_l9��8��-�<��ܲ��3~M�N:�&i��75���ն�>��S��<e���1hTt6��r3�7�;��@
怭��E��y1?��E��X�p�R�/%p��l+%Y���s�v\����jT�sy{wD�1^c�j	�h�<�l�}t �qMImدvV��E��7�u66j׭���Fm̦ԩs����ѫ7�-��H�o/�kGW<v�z+�i@vHj��xt�P�)�G��9��t���(yJ�u�RJ���uo����U��M
1U5Q�ƨzsu�h���*�m[cȻV�h��6�kъ��/3�c�RPEd��LZ�N�X4vų�*b+ZM�1u���mc5t�킋F�q�k��y��;mG���G\l�b+��v:5jڶ�Tj��c�EUt`���ڂ�옢#v:Mu]�]���n#%ck�:ծۨ��-��ڻm.���֠��GT�l8���Sb�ֶ�&*(�����)��kPM�k;�������U�m:��ӻ#��v�*�֢��t���TQ���-ݮ�M�Z��Sv4C�6�ݣ��ѧw4wwUэF[-�]�OK��:�]�v�m��(ѭ4���T�UEwv���Q����ѳUl��j��U�3Ѣ1��(��lTv�q6ŃE݃�B+�Q�+��Mژ�nؘ���l�Ƃ ���m����ul1��Սv;�ڍ�уDQ�ZuSU]ڣ���B�D0#ɛ�y�*�kf��9�J�tIO��c�
����rݭ۴QK����lu��6a�F���4<�Q��`PP�����k��u��?~�����f�|��he� Dj4&V�i.;3�S�gb���p�ܛש3���c�q�Ḵė�H�'_\+�̎���^�����gX��rG9�\r[|O\O����A�F��>q����؉�)z4�t�P��t��A{��Es�D��:AR�1��z�l�sf�b^�f�3FtX�F[�YQ6����vw�u �FN�B4��r�������\��rpE7s�Y�D�R�ė�kVY��ʌ䣼�'��X�n�K]�td6���)-�|��T����W6k�T[x����b픡���1~R�*����I�J��a�ϰ�����b�b}���'��͘Q���1#wP{^�	w�I�qm�T��e��]�Wmi�(�q=&���O���Dq5ٴ.#���PqZ�&��%V�;�����w���S\�i��/ur���HUNku�G`^�s^�*}ר�t{��4C�T�J0^ �
{��}A���m]���|q$��?>Hc�������lQ�L�|�n<��'u�R�����	\��YW:����v�tEΧQ��L�|U�L��!��ܠWk�J�Ｔ<��~�ui�KCw⫵X*�U�S��=F-&gMD�OT�\G*�� |M^��fEj��f�mrF�q-H�VN�+ۆ���˰����S�����Q��ְ[���~��P��1�m;H�v�=�cF|�%�e{��U�8�l�b�}�s���ڛ����;��V�s9���2�'�I���u�'喡�k�M�/�t9����[�]���wu�ΚQL�w�u�i�A3�ŭ������^��a�:-X�w+~<��Z�\�e�Fƭ��ذ��7�9,�9w�bH?�Z��_/���>�>^0��;�9D2.��9�[���-ʚ�r(�b	`�z��[�B���6�~��K��G���Y��С�_s�,���Y��V#z�0�����5�n�:g_��r�C�/.�&#�@4��2�"˓��e�z�p.�>���Z�Q��|��� �zCT�˳�YKs�����~˴U7��_C(� �p�uP��]ڑ�V��a6��y������b��\�I�2�qk��;|7���m�%r��!�:ΐ�j�����`RtB	SC�37�>��cN�#k�\����S�/�_��+�}_H��)��c�����BUbUy#Tt���II�2]L祬�z��,��p%��C;�����>zUt�ED�Z�n R��^K'
X}]�ע�I$S��OtMA�&������54�9kzGl������sƬ��)����}��"�-�*��q��m�!��k�AM���p��a@�%�ӵ;�\���BkDOMqʺ�����W��O�f2�2�u��W5��휅o�SU4܂�ٽ��TAu�
�J�
�����ϻ��� :[>�4�]U�KTGk#s�a���xt��$Q.ѷ����<K%��}��F��:��Ń�pd>[�x�������1��W@�S>��^�-n���A��u�8�����,��V�ށoW���DrS�����[Ȭ>��0����m}���=u��;��s�3eZ붭'��@Z:�J�����/<��z�K�)�^-��;�$Ӧq�Ҩ�6ەv�/�!$�t�ь^�O��U2��dL�0_+OA�e����*�:�mf=�O�M��w%�Sؖ5;^�A>[{�)ڼ���5��K��4�Y� �e�K �O?j;��v���u�:���w�z-�*�Q����]�A3=>ݶ3���;j�y�c�®�W##�t��}S�m1D���OU�k�m�ߣ��Ӷ��ca�z���d8Э�ї�Gf,H��빭M�\���lה�9�#��q�ܤ�r�U��d>�e�b�mTT���}0����HD����w�^қ�"��E)\y��^�wMz��S����KUޞx�-5{�"iU�콈�o�ᓥM�߰	�|� ^֕%]�X��'��Ut�`�5Ժ����V�:Zc���B��v{|4E!s�C�M��j��9���+w��L�%w܏1}��k�j��,�x�)��Dٞ-����v�Y[��.���xˤ��Y�
l#,r�i|5P��bF3uݨS��D]_s��	���8��]�ׅ*$�8Ht{Q�:{o��쨙^Z©�/���G:��l]s6yH޼�)�vVf:e
��)������K'=��G�"���׹�r�X��8t��;]ݼTU,8Vͦ��3�s�P�a.�
S]@%��鼩[�LM+THR��r��&{��M����G_|��q/q�{6���f����Z��03!���h�.Z*%���J��N�{l��˴�J�ƑV��[{�M��2��8�c_DT�]sFd�b��c��\�;ǝHa� ogO�u��l�N�-VQ<�t�M���7L������2�I���|}�8�<���g<�Gb5^%+��>?�Ny'��6���@^�(3��OjƆ�8-a���5���ꈄ�)�r�Bo*Lp�-N���KRշ���C��nGr��X0�/��KbR�Vfcg�1q�#�T��#��9��+��g�%�A��z�t�Ki���);kF��ќ'Y�m�I��FK��g�R�z�������4��X�U)/A�5�e%̷������4�L�f9���G�g�d�ݧ�Tʡ�3�+htVBս�4esm�ۭ���R����G�a��5w9+"l�_?��bs4����=*rY�-E]0�:ba(Mx��@	�� s0�a�]��S}�M��Z�4��i�zl,	��S �ړ�WF��j�k׉~��bk�L�Xy������7�2���KDԨ��K�١�JT��n��{#s3VN�]{�eg����f�W��/K�3���l�!u����=�Ǝ�������A��W&�cG��w����v�Kܛ����\�氛�!��c3܊��u��AHWtN-*�qn3��� khj�]
3�l�c������t�����S����ЗQR�z�܁��PJ��A6c�4����)m��9�ƹ�ٕ~�d�8��&%XQ޲�-�V��b�ss+���wW�v%�f�0U7�ie��/�zn�ď2^䊼�Y�$r���{:�s���fZ<s��AIc>n��ȇZ�6���U�O��x�wO��̘�1���K�Ó�Ƌ��s�J��y��}�,�τ>��-�u;o�Om�|;��k�cQ��6s�:��Wu"��!s�����5��Q�1V3�������&J��LFڨȠ9+�Q�2m=J3�Z����xy]E�[V��[x���";�m��F(n�4��/L2�:=�����!���W]'\��x����f�&��>��|������]]hS�ߑ�ԝK�e^�
p[u"1�[�\��v4�uk����}��\��{Woc�nSx�+o{rT��P�i��gn�Q1PH}��
� ݝ":�ܬ��-=ֶ�O^��}1�T���z�ӽS���� }~�yLa�:��3�7\_ٛyg	7!Y�ޛ�ꭳ�
�Bȧ��b��LP�z2U��9�(�{b]5�M&|��޶]�y�y�.�"�%JX�)a�K��J+�F��6b)�p�z�!��ȅ��`��"2@��*١e"�2�2Z�����%��S1���{���UMe�zz��NQ�J*F+e(�<���Y����v�f�9}[�d>J�[������ ʖIĮ/
�ۥU]1Z��#��u����F����)�O���<�4�KoG�!Uv��rN�w��f��Ø��ν���l��aK-{VeW��<
�:�jr���R��G��Is��]�|f3T����ݭ ��^9W �-F���v��!�f�!ll��|�؝lŴ��y���{�zQھ�r�L�/k&��T�C;"�c�Cvc�����͙��z�A*�����#�Wq���3Q��������]>��\R�c{�/T���^ڋ���F����b���iJr�S"�u��v��u>@^�8�R|�1�o��-�tvm�p����������Nm���շPϪ}�8�S��{;��Y���5�ս\'�H.�"��6�oB��L$��_���P��`=EJ�M�'v`�i�3�}�
}x>��s�O��UU�/ �%C_�7ir��ʴ���)���g|���w�@l�0��AF��3Mg"���e l��9�*��03z�ٱ�3`�0y�z��}Do�ز�n��f�d��dΨbx5���{D���#lm�����6�U�
�j�$�2l�hΫ�.*N�#Z��a��ݕ}��׌ٖ4����r��{-�lݖ�I��}y��]U���� ؕ]}2����>�aL/O��������I���16b֜�g��J*�^�cy4ϒ!H�(BU^i���MU�/]��n:x��ħ��6�y�t���w��QXKϑ#$*m�Ɇ�%�˵P�����p�����:��[�#��� �]ut�N=��c���/q���(@��y#��QR���q^ �Q�^��Y̷��rچQ���CF�[�R[Db��Pq����DDK�Dpm��tRO��\�F����|�h����v�̝�W �'�#�{a����=�'�������֦	u��Hh���hȌ�-�UL���]�El�X���9�V��KL�^C�z�sCN/}�"���QF��굙"
qmU�8��o���ɂ��L݌Ź�F��܎cV3�ٞ�=��<���U���m��̆�:����&�8�����t�9���"v�l���#W��� K *��&׶z�me�d�]1���2��˫ި��>�����>�Jx��e��[���!�cTLIa7]�C�鋢���r��u����9	m;_^G��\����~�Եj�Р�y!��/3y�P�o��VG�BVG��%
�.���uz{cq
�)���߄��wnDtv�i�ɞ����\��eAx[ڈ�Ա��WՐK
g/y�gK_d�b@�]��z�����P�Y��1���#�{k~ܟ1�Y���jW[�Y��ebOk�L�5�E���^]�s��+Ďo�9���}����k6��b�T*�6'A��s��Lwu��U�A"d�vt%wV���u�1�t"f��ޯ�� �[���N�Z3S���E5g�����Y�8^h���2P8��ʇ��m�w���Y�3 ��-��ȌȚjRPd�cKq�%��4�^�6�زg�� s���1�i�{J�<s��a[����[��̵��1 �UȸOp�v/���� ��9��Z��f^ً�"B�n���X�P}ʯ��+S���T�Ϛ0�ۉ[�wFԳ<�]a�x�a ����z���4�>�l3猏2�#��[l%�g0�>:~���ξ�+x�(�K'4v\T��j2�q��]-�<�t27'x��n�d�H��8zV�	nG^��$�^�Vz�)�˧�e��"U�q�۫z�_1"����F�q��K�iT��+��m�v�'���F2�a��k�͖�,QY�A��`��)Y�VSJ�f ;Pz�	O��QVM1d��eN���C])�?�Z�����7�0��_�������?����w����M�����Ǣ�DՕSR4�@:��ـ���b�{�!�Tl� <E���7�SdV;��E�]={�k��d�O_>�07ptAD�-f�gxGsW>� �A�쩬�݆��t�ˬ3��o{�TK��rI��u˂�+zr�$��E�Ыl�4��y����y;ؙY�8]�J�"#�wvo�1��}�=�=e</�5�	^����}�DR��ui�`;9Z�DT\u��>�)r�����c�Ρe/��K12�ٷ��GMƘ�);ǖ�d`$#�L	5%\�2i�N�+��	O�}�U.(�*WPI���cɀ�z�y"� ��m���ws6�)�B�M�f�2�-��z��)3B�������u'pc��{W���5X=�/7us����9K�=���ˊ[�,o^��9ՉGc�WZ�Z�#����.�(� R�T,��s��[��m�<��l�Nlj�O,���)RV�`���WMP�Nɷ��.Fw��.��K�x���F�E5��NoY����9����x���ì;v�f��s���w�z�%�/Q�z�ťᏦ�X�Rؤ��n��$9t�b[q.1k*�����⬛G4>��׊Gz�����F��b\ݬ�*>�B���kb�g������+����+n�1��N��ރBTU�ӧ�䦹ua*�9ջתl�c5�i�Ԟ���x��p��-"��9��l�oE{Rb|.�<��$�uh2���h�ekM�O��얤��;2e�"��2��x�t,���fPq�^R�P%�R\���q���̼�Z�� 	k9(N�
�Ѡ㹎��7��gn�X�	�
s\N��f��q�+Z�-Q����zɕ���00�+9i�C��$����	G\�*��v�7����[:��M�Yw�0�Z��Z�j��{��M&�^/hj�i�4�hZݢ8���e���q�O<{�WL	[��ӃUYS��-�;�{X {��j%9A�l!�B%f������BM��>��N��g:Z�LL��G�O�:�kW_�+��ǵE5�w�`���Ph.�9�
��5���R������n:���&w|�	^�⨹خ/{;�sЌ�D�N���=A��6T�z�!��J�ec���`N�+�4��� 8SV��Ӗ̬�������\���5��G'�*κ�:귫��%���N̖�Y�Æ�6)n��J�l�cں
�f��3p=�%.��"́�]N�w3Z�+)�|k�"���G�#j�q[�7TrYg�xjv��v��s7;�����6�`����k�yҸ�+����^s
�[Y�t$�)��k��};#��1g=�)R�ޥ��8��MjW�-8�A7I����Lyͻ���������RG`��=��ĩd�������N'�wR�}]������Z�\�,S�%@S�#��u�m�Ql��hQ�a�R��d�5MĄ� �hFJ�Qo�1 *$��:*�jؠ���]��h��ݻ�m��mv�E�ؼ��<�۶qӈ�N��uUSAlm۫���"*;7U�&�kZ":��ucLTQkV2h�����ٶ������[��lwtV��u��ww1�[[k�����:��5ӶuGl�T�N;Z���v�Mi�bX+m[`�Z(-`��$��V����:�'�uV�&���61�&t��F��J�*���υ5T���(�j+lu�D�n��PT[w:
;k�j�;�롭6�ۮ����4bJC���7[`�"�����4MA�;[2UQGZ�i���h�n���ww\N�V5�UW�WcETDU;*cc0ְ���g����=٨�.֎�'T[c�UlmwgY��d�k���V�vi�:5̝��gQk��q���n�
֊h�������j���ws4^wuX�Ѿ�~��~�fR1�n~�8�ڜ2��"'��+S����n (�f�2U�ȸ���P��[H�|��j����d��T�4_w_wv_!HP��6ZuE�.����{��W�Ӽ��:ي���)�Z�}���\��V%�����&�::2�U�38m���o%8�p�7��u�̫�f,���:f�3��\��+�d�̣�q|j�X�:LA[�Օc������<����uܕ�gcۓ�vs�8�z�Ԃgg�[Z���Nմ��g(<��;
嶚.2#��ʍ�;C����x� W# �������n�13	�7H�k���n��\,5vtb��;����<����0R.�ڨ�X۾#2�z��\`���ƱФx�ю�����>�h&��[5)�yKז3Q�&����j�ݯr�V��e���Η��B�윿ڂ�/�.}rzt��V[�����vr���g�B�*٠#L�p�-��g�#��}�v�`�5~���z����:�����q	紑��`b�R�yޮ����6�u9~+���l�s�<�G��9W�&yc�4���^�0�ɯC�]�$(���s�*6hY�{5^�zLw~�o�.�Ϳ4�:2�$�n�]��N��8�qk��ސ[p�Ӱ��V��,���)�<�����;x���M�w4�w�{2���NsS�J�m�Y��W<m�f�\͵Q:����Igj��)��c�����.�vtO^B]9"1���5c僯��/7���6N��V@&�q�ǜ�u%��k�H@6���ZmF��^b��J�[Ggf3��{M�r��F��6E�)�`��1��vt��/�7rt�nY �"oOwy�J����YZ��{wǯ�ocǜ]�(�͊~���\C��A��O�{�O����ĉt�s���7λKe�	/�Uo���s�������X[�$��L3덁��P�%�����l?.�w]�P��%�j*h�SE�1��$�=���{�G�P�psUV�V��\:hpv����1�5{�*~��a�im��ޏ>�K�����͈%TC�+K�f�2k�����Oa��{p7d���)G�ј<�Z�
�D���L�kh��N��N�͹���TYP�jme�-���X�f�|~�'�f92ڢ�:�fW2��(N�7�v�a��Ao3$�XJ��tι�']��ԥ��u�OhpMDPr�oS�I�u%d��M�cw��'щ�F��*�ֈ\b�hm��1��0���F��]fi�l�Ӕِƃ3X
b	�/uZY��.�o"i��Ǔ:(W@��>�:��6�!ʔ8Ӭ
M0�RE���j��{]�n'�]<�Oݞ��V^�����*Nsт����Di={99m6�Jm�x��Z����&��]^�a�ֹyD���=��n��&�`Ӵ�AC�Mt��&��c5�9a��{51�bubY�%SŬ������=U���B'rO\�8��c�{��<�C�[��HE
sqyx�dS�m�HY8��3���r�%�IV�𫺯Y�Sx�e����V����F&�W�rg����
�� �f�箈S���K��W�뻄k^|���i1�����"�5�o��m�	��6�č{��U�V�����Y��f���K����ˁ��������.��B8�N:˴f�T8�)4��ӝ%oK��N�*i��J���e���.���$3pv�"�MPx,a\�e�遃�T�H3���c����}$r�ǲ\�_%}s_E�qA�\u��ܬǤ��c�h�1�iضf�qf%��Cܫ��������<sN�:]�ȍ[ٰiOz�C�%�������cL��KJF�wO�Si�k� ��7	oce�Sb��k�0	=qm��qN��ӕG	�Q�2N���F�����`��`z�:3���odMgh��{�maS<U��VP	sܛi���r }ŵ�&�rk�Qi��xj`���d�g|by�ç y|7�6�;df�Q��e���87 �O���6\n�c���1�|�k�Y� +���_H�;#��6sA;>#�`��ƑSb��<����Z�	��]Lζw��LEW&�N!wN:��=�Fڑ}i{��u�Dd}J����~c�� F�����ɦ�e�i��*q���Ӫ��F^�Ž��$l�L1S1�ece��x�e0�-�&�YQ9�Yh�P[Lf���UZ$�ג��V٘��ji�մ<��o{=&`�MM�����8>� <�V�U�'?(��w�|�g{�rRW�k饽��/˰��P�[����V�7{��u-�h�y8^���&�l����DtV�t�Hqx�nК��>�bt����,�����V
e�Y�'_'�U���Y��F�pej�d��&�I�6���6s�(h������q�y�� ���]x��ֲϪ��?,�m��,Lٲ���a�O���+�}�H�=gf}�hoJ]`�[B��d[����Oj����E���^<��m���P%�é�us�(�S�槸�F�F\4���{w�����騱�m���f�ul����3gG$"�'���J.�F�ݍO֬���$��),d7WH�f��-�s8qL�eYT����Q���Emt4�D���a��\�l�e�H#���2�Fi��%£�����%�왘�H�=ol̏m�oD���g�R�>�5�KuES���1|3�1Xt+��/���Y��u��UܖW�ƹ��&q�*xL�YW]�q4[�Âȱ��� ����{VI��JC�ds�,�z�p�3�Q0"15.�uݹx腻A�yw��@]�#�ݘ���<z��nI�v����μ�1��A���h��V�vU`��T;�]����;#W;�v�I�&9'ħFjՏ�;\@�@dzJW�8����㔩*�[����Ю��'4����cx�ck�[O�xw���_umNS%ds��m�qï��i�9��~^�����puű�t)��d6v�*�;��>�����WD8� �z�88�Ǵ��,e����!� �r�b��b���7p�_5��<euZo(�1�S#�ΐ�AV���5����2��j��O���/3�|ԩ�����H����PP�*:q[%�ktt@��k{��"U=K9�j�zv�2)�����R�R��Ad�WSz�]�&4\�G6�4Um93��g���Hk�jt4�Y�[�;fVn�t��g&��H�,�͝-�u��_*� �ʠV<xU��_M5τ�p&6�y-ؼ&:���fz���F���(�{��`7KQ�z����5�8��u�z&��2�,��/�:��;Ǥs���2�o�l]Y�)���bѨ|1��ǃfM5�kMY�`AU�e�YS���#���Ѹ��=]��4�C^s��>��+��2A��̳b���/{��c�T'^���պ��¦�U�r�!l[}YY���j�j�o(�kn�Y����)Y}nMK�����=1g�8qF���b8W�k�U�e_�D]e�������5��S9t�qr���̫���%ޝqjS�'nI��nP��?��9L?s�8.66Ҫ�K׮R��I�;���M�h�y�8:;옪o�_
c h�X�ݚ�{G��X��7~�Vy�a�PQ��j�[����?ݳ�g���O�`(l#��+�?�|˂ �%�<ީ�������|-sb��i���Xb��,g���t��M���]�M
�V�LM^uKwi�l�!���1�h�"ڎkQml�&9�ֹ�w�HE�	E
U�绎�Pc|�Ƈr����9v�7�Se7e5;U�A��r4(F�-��{�0Uى�$u$�ʹ9��1#�����/�2��&t5���vY�**�Uuл��ᘚ�^�\��a���vI;�/.$I¦�����k2�1U/rd`f�{_�C�(�15bq���w�z��'��� �qM{;��m�zxE�:Z�y�Qr�CZ��N8E,h�4�:�QV�F'{�9�q�6n!��4^u"��G��O���{Y�5���[4	/��OvpV|�yU��-�&���<���"�oKud8V|�oY�.��o�;�������6�U;��EEs�p�����籔���ڡ��7岺�k�=g���uԋ�FZ��f�P6s�u�~z0K)�o����N�8���V+�Fi�tLΓ�o��i�v�3�KÝrlq��͜w(����4�i�%\��l{�\òO�Φ�-�zWb��m�l�}^�]0h:�4Ok9@��I[�4�g<'܂�y�t�֛y����>&�q�U<������ߠ;���� ��y`���7fG<���,�Y^���l�W����Ś�ق e�>��w+�m��z��ZZ.���%�)c�;������)K*�p~��e�b�֎�6�t�m������ޟDv>j�X��QoI��1���٥ém��ft�іoD��ĒHz���(f|��)+.�n�W���\�B�t)��M�5w#d�c\�@k ٲ�\F<�f`+3b�/V���ܓ��@��ܨ�I���B�ȕqX"��u* ���|�p�U��ݦ��G]A�ӊ���T��D�l�������Ғ�{���C�������:�9]�,Sa��vI&�gt��n�"9���mF&#��Cť�j�RW�)Wl�W����y�����ce>�m]4J���Nʡ�^o8b��ќu���n�v��gM]�>�
����s"��m�-�6���B	��;`���x�c�8n�M;	�1r�
{d��uk�	ξ�#�q�$6}�V)f��R6[Lc���O�u�f9���"U\R<�'u�j��4�埔����n)�j�'�oo��渷]2���\a��Y[�)
㮁8���v]���m�]�-0�,�nU@eV�5_�P/��6:�	JW�f��x&�,�w65s1���'n�o[d�1�8e�Dr[^��:�pK���8��ئ}g��5�j�v��Ĭ��7U@�{�&�Hj�)���d�Հp����G�[��)��}6�����vY���3"�_N�|6�*���d�!x�G5����AØ�ۺo9'���ս c]?��r=zIUf���6��ʐ�B�@�s�ޔ��9�{P!W�r�v�ŚH%�ـe�Ա1^�\��:�'fsv'h�m���)�r�P�yj�=.���{���{�9�1K,5x�,gDn�Χ*^2zIt(̈́\�ݤ���M���<9�������Q��������k3x+�g�MΥ��}L�ģ�鍍�3��]S�n��a[;\���<��7gtg�'4�{<ې��jQ��=��K,c�F�ƞ����آ��I��6�tɚ�ɞ*����dK�k�Ó��!�ROC��.����[�k왝�M�3���aawW���2�C1*śU�����jy�l޷�v�U��.��8�X[�@���S5��T4v�Ǭ�G\�=�=hyb�v�m��z���`�Z� 1�S���<��0�#
�l�uC��え�s�"�=q�j�#3�����V̌��0�k;�NY��M#x�L6V�"�Q���z��	�F�Rz���k���/[0��M��������ByG� �9�-���Z�P�@��%�`�m�ɜ��Pw(�����e5X)�H{�1��"B�����W������z�>�O������{��������.�w@��{�s��s�<�KL�n���8&�����n�U���*�*O�'�o3k�w�m����y�$Lȸ�Nwc�ػ������"j���УB��w��Pʔ���]��&�J�}��(�q���[�log��K"�	iA{v]�4D���S]^��y�|�3c5��apĩ�{ɛ�j��W&��5p_6_Y�Б]�zS�@⭩w�j�,m<N�TH��0Fںq����9���ͦ�3��0�M�aʀU��Ngq�Ym��:���j�j�F���Wi���)p�l	���ɒ�+��z0*������sn����陆�c&'|j���ޗ�0QM���;���iҦ���:J��7�N֗P���d3H�E����#{��Z���,����kk�����v�+���+�@���MVN�Z�8܆�݃�l��3z@�s#��'9vZ�t���	�6 #�if8�wV��$�!eun^ھ3�!�����f'�T�H����<֋��m�{�:�*Iu$�P�.�x����1́���X��kJ�2u���7.��Z�GX�\en�2»�eibXR�9�t!��������m��ܴ�g���s���&�78�F�s�D�G.�Q�'�l'�����96��N�z��*�ɲ�6�6Ō}s�f$��J�qsF���9	�ab�J\�ű�[�0�
Z���^7s>�׷�xğ^�tF��uB*s:��ݷ�v:�R]��q䵜f5a�*��fܰ*,E�%u1�W>�h���"�)Y��w\�4���Z��*���IK���ƍ#]��� �O�U������+��݈�[U.�mr��K�vo��bx�}�G�G^P�
�y��1]y��� bQ�����6�4�~�r.ɺ}�S9�j��Ѳo�G���J�ؙ�n=�NVEe��-y�e2����ۊ�쳖КiI}��X���a����l�3��ao�Ɛ��7��m��wW;zi�뻪%��JJL2���3�x�ġ%G���
�6"�g�&E�T�;N���P�5��tZ�oR�k&��7�b^�L�1���,��,�<� 4�VjGoqb�*χD�b���Mݩg�ʻ�}s�r'���ήu)L�����Åޘer�D�뷴X�(iʛQ	o9=z�X&iyUh�k��������b�aRU�V.�O��� R�Lsfe����fU�ov�`�rEއ��iwn�F3�����t1T� �c���O���C9�Sv$9ԏk���so��Nʜ������k',@ƍ��%�M�!������̮��B)q�s3�،�c:�2^"�̽X�F���ۑs����W��pjqǳ*�Y�٣q4��]0CPL�&!�D��?Z��u�-�)&r��i�Y���'uͦ�9]�-Ԍ�L��ﰗu�^CCs����1Y#�!
�)R�hc� �$�Hm��Ͳ�$�b����A;gA��5��
��8ضtQv�a�ۋ�g��:h�w'ws��{�T�F������h��փC�GN�b)�G�j &��G����j��yjn,i��|٪��q;N4j���|�U��F������QEF؃��n�5�Z�7e��1��]��J
��j*��
"Jmh��T�U��SDA�N���"��$wk�5T��F��5���u;�lh��v���KZ�AX�c�;g��Ɉ)֝j�7c��tj�((h�[���VM&֭6Ǝ��5�UCWgT1v�Q���)�cj���5���Ui(cS����ۣU�+U�g��bj�h�����`�F��l��cf��	��[jF��E��l��L�ݝh��_i��n��O���ۦ��,"�$¡����r_���dA�.L�'(E�-�1��r�Rl[�ʣ��Ū��ʌ�Fbɐ	γ�mof�)�
���˽�M�FJ��U��b���)�t�W,,!W���x8�Qco�$5%�If�9W �-���O���`�_{"��n���.�?u	v�NA���Fj]\�%i���Y
����I�G>_(g��z����M3�3�y�s�Ղ�U���s9s�<�zF5�ke:!/N��c�8��ԋx��Y�9������U|K�J���(��\\�g�:gd[S��r��hQ�(��j��׎6��⛫�0�Z���mƛ&qI<�k2��Z�{ו�Aa�6_l��9͗j�P1�"r7�������ݖ����f6|M�H�ia�y���3���OSӛ���Hnv�4�COA�'o�ZvFl�!��f�4��u�U|+KP��L�x�a��z{����b	�����~��WQI�!��Pv6-�F�t���*e�].��طoxW�:E��Հjm;�WG�:��jE����et᫑����'j�����9g����k�9���:kʽ�Sk�y?wk�y�#�6N	;�-J�ke�c����S�/��Q�ke���=�R؛h6'0޾�|�fVf��[����:�6/�";�����	����n���O�6<�Zʱ]ou����K�2�9�-��~F%���U|�%~=�6�(�T�|��e�_���=ߍ����M�B��s���Q�;v��7�vI
O^jz��PŎ��� 5T7.�����Rc���6Yk5;I�Ί�٭�t5$��$훼�WuOgV�:���O���+#/N�]$gH�FH���d��G4qG��U�걡�����3�2ӳ�+s�����9��U-n3Sc��d8���6�#l�O)��,A����,����Lގ"&Z�Tw\e53�ĸVLp]"Ӏl�G�y-*�\4���h����"�;�v*��/'+�Ǵ�[�\��x7PwY"5oc�s��3�E)����dۜ$�ϴ�TQ+�(��-��8�����ǧ�uO+�ݔ7��ǿ�Ȥ�[�pA�k����U��?<�j{���FP�5�;�[<&>�y���;��8d��+�.���6�A��_~d����09�5�y�ک{;I+d̗����J�Ko��#=uڮ�z��푸�_-�Om������$pgEI:
����\6�|�룂� R-��*��vv�Uf���%\v%T	J$R�1��)p�})0����/��;������T�S4re���å1 dgwqŜ�{q�]�cӋΦ�I�e��m9�,��uuɲ�7���WyYp�f��m�}N-_N��k��g�\z-���+]�}�·O�6�5ؘ}��Y�]X����{E�8�Vv��'x3ʾq3�LJ��&��x �_7e�Ȼ�6"ʟX��$�����wDH�]��Cq��L���2����]�w:+�i{l��>�][����X��F��ކbJC7��\��h���ag��:��-�c]�׳FL�m�"Ԋ����2i	�;^K'+ڱ�K?,ʐ�f-�kr��%�K��ے���/s�H���{гy
��ƼN-�h��&KE�*�����M�9>x���U��k����;Ʒ��vW����}�P�
�]+V3`k䉺}.�� ��<BC�s�m��[���N���:*l�o9Qi�qGu�J8�]2��hH]�MW���y��AP��gW,*r�Qo�&�Rἐ\�j�Ü���b�$��nY�}p�ŒGs�T	��J�{����7jBW�"����;i�D���:�3�לke�Ъ���ATK�|io_�����{��G���6?�.�ڕ��U�k>�-4C�_V�&j��aD�tRh�[�d$��%���g�즔F��i��9x�<w?�`U��+iH��0�W$��z2�U�y�=r��S�c�����8V7ӷ>�*DGoT��ٙ���T*w,���xJ��p{Y��U�N�v9.��AM��W�ty��Ԫg`�޾J�F��*��g-3��x5Wm�����7{zL�5�xw�`��t�2D	��7*��3�SU=���|;�cy�
o����ߠ��z܀r��ց^2��c�����Z]
��[{�5���x�j���rp�=:���G�$�sG�N���l� dy�U|���1��>~\������W�u�j��4�-���c䩬e�Y׼��,���rL�+�K�7�]ʲ�{��Aƞ���>�VVLŔ/<�V2ގ��eU��(޷E���ἂ�&��Y�����]FP�O�	��3�<�w}��Lw�m{�VFۺ�\2��\��5���km't��,��Lv��ف��lg �o{�@_��w�7�BZ��@_��t��,�"��kʻ����ܞ��ς��Z2=tj���ꮼ!l��Eu��\��{�t�.�)/v�+d��)�Ʉ��oA�xkۆv�}�z�����-�ga�+��w����[[k!\��&FC]�cP��@\�!N�,^�gc�E�3�X��&Ws�aƼz�;'��Ue#�T
ǏVc��~��qQ�su}��u˱�+r��g��xKo���®|n��F����\�c���v�UDlWt�� �[)�;d_��Wo:I&�xUꮬ�,N���a�k{{i��V��Dב�p�a����	~a���ޅ�K��x�R���-]>s.��*�=l�E��r[���t�}�����}�~�v��M���d3����+B[:ٰ5��,�����#=#�{�g(�!�"
Y�nK�vj����8�H�<��3����E���.t��g��Lz���wag�Ү���+���U��ۣb�\���^�Q]<���3��S����[�b��&�ifq�3Q���b1]��l�������=�òQWϽ]-ׂ���L�����J�ۮX|[F��YTh:4=��k?򫉭�%v���xԯZ�.��Yc�,��zfvA6� w�Ì�bm����Da�u���N�a������Eh�]%�曖�ݧ*��y:�(7�}�.I��v%\��_ CZwW�}|�װa��v���H�B���0��w��6�Y:޴�*�����x�%ӫ��t
:�w�p�/�$��Nu��=Z��x���v�!����'9ŉ�u1�rnR6ٓZ[]W4x)�F���ƞӺӫ�i뼃�ᑥI���m�����z�T�٥���/�䇱�&�$��s5��&Tg.��(�+�nn�U���_Sl���ti�FN[��7�iB���ظP+6N_���IV��S1;+��2��s2[�7g:�Kv6��-�2�H�qlE��mi�s�Ў�R�nǎۺk��=,�L�j����ll�1�~q`�ZT�����tGuԄޭ�x]�a\$y7�^1�+N-k+r��	����Ǽ�R��We�w���ܛХ6�O��{n
��V�=����ǌu�۱��
�b��uǊ���y%�I��c(����''Y2�^t�z���K[�\�0�͐�yŹ"�(a��Tƥ���Q�qIw�O�=�紿KO�D�T{�.�������Ɠ��f�˶C���F��@.�*����$"mSv"-�<
�K��_^�!�~�g\4�ơRxCIK����z�:�ܒn��*m�F�l����E��u�*�s]�vL�s�����&��*���Ֆ
=e�Ȝ��4�kw�U���7Ÿ�Zوݑ`dVwrL5���V� .��n޳6�]�d��a����b����4y�)���r�m5��48嶸�c�ִ��6NMDɑg*�3+n����y�+��"��̈
̋�z�<Z�i3P���XSv&'�`*�iC��|݁�B�1eD�԰��	>�j�{�3dB�[����#�=��(B4�B4�Ft��$\�����S_�3�}-�e�}(]=�5 n��m��D�mP�o�M���I�o&Xy������p�ռW{�u��������Y���s#�E�Wij�<��YIP��Y��B��V:mK�V���D=�R�>u@����<O+�)K�q�j�Ks�6o:�Z�G�>�>��;.*�c1%�<�b�j���u��!�j_�En��13�&|�	L�R4DV��x��d�X�n��&��p��=�u5T���ԩ���@��	M� �
�*�Z\��q��k*^�������Q+2�w;�`j�cW/��)R�~؎,�Q�cYCB��������2v�fn}��RW�"�Hl��U�Kf�Vڰ�^�s���	"f���ǫ�	W�U�)^׬VG��bG����`TKa�<�9�3%[�RĄC}��szWuƀ�رvG�7�9����N\N���5��sGnW~R�����ۜ��S��r�b�=~|��Z��V������km���-�5z�2�Ko)��f��-v�aP�%���0;>�Z�Dn�¡�&X���u6)�=.���zgccz�{3��z����9s`�5T�f�v{��(N��XjfV�L��F�H��X#뤺� �]�:��).�o1�*P�x6S���n�b �k,^��,���L0�����O˂p��u5W�n<��1�����c�ʽ�79��#�(!�&�'�����J��q8�\�e[CLw��c}��w+�}<8G�ٰ��<���3fs)-l��.K4�Vm��mEnAKp�t�z�|fvI�ǽ����j�G�cD�;?':�-
{�B�z.K�ճ��oXc��O\�5��({��M�Y盀�;��?����HN�C�T�E`Ţ��t�l��$`�� a�R��j��m���w|�`~E�@��%��KC���\�Y��&'t�)���Q�c_�Vq�6!�?d]v����9�0n��<d5*��2=u"��PJ:��L�mc���]q�vZ�r�7Q�M.h��ݶRM���k3���b�|����q/]��t΃����������N%qe\+�|Lu �z����-]���M=<q��̎��W �@ݙ�5.�nxՕY@�ʠ
ǀ*�l���T[D��Y6+A�%ۚ_��A���a�%��
<o&�����u�4z囜垆��q���kq��J�k]u5�%p�J���Y�RL$�d�O/RyfK�T�r�(����\t5�V�
�w.��@�V���c������x�*��Z�7��ď.V��:�0�{l��-ԭ�V�k�O^u��]J�}��5R��!�#��p���mG�iyֵ���\n�O��t���sJ�xϘ�L���oS?Dwi�O#����+f�7
<6硤
�R%�~��˦,65#�{�S|=޷\�����W�,�nFAwh��:θu���lm�Qt��	�1������G���{����o?(�)�{���d[�Q�5����+z��>�z��+\��˭9�X��O��_��9� �w�~��u���9��\Q���G�Zv�Q9V��L��6�#���s���#4f���������-2�6et�IW�7���r�E�ˌ|�噕�X7�#i�^9Ph�L�����N!�cFu�af��;8k+XEO���LK5�e:��I�4f�85ҍt6�vm��)6v�qWf��0q�G�����v��&B>�FO�p����
�Z�c��`"�����}�������� ��x���/��G�� �Tw�pq���|O��� ��U� !�a�a�a�a�a�f��	�fU�@�`!�D!�!��$2�0�2��� � �w�|��9U_��" a��P[r d@�ܠ�` 2��*	� �@ ����� � ���   �� 0�202�2�0
2�2�0 7��P �@ �UV  UXa a eUa�U�� !� !� !�U�UV@UXeF ���a�a�a�a�a�a�f &Q���eXeX`XeX`XdX`XeXeX ���U� !�a�a�a��|g�||A���x�4��((���������������������/���|�����_��?���;��?���}?����YP U���������W�>� *������ j~���?�?����� ��/�?g���$�?����?W���D�x�� ��+~NPaQQ `@ �@
 �X�@" �UY� %� "@ � ! 	 VUVRP �� %eU`a 	X@ � !I @�z@"�H@� !$UiUZUD� Ň�������ZUB��B�o�~@����_��
�����~@����tW����~������|O����o�?������pW�?$?�?�~i��@_� *�Z���TA�p��E ~ ���������_^?���D��I��8 � U�?��_�  �����>0�����ϫ���������W�����W�������_�����}S��a����>}��>�`���>� ��>"����� ~�����}W��O�W�E1���x� ���_�~~�G�� �~����
�2�ȭ,:�'+b� ���9�>�Ϟy) �Wl�Q
)U�)*T(H%%@"*��T�i@�VؐIR�%�J45����)�"
���ږ2�3i�Kk&��alSm�[kbi2�fȄ��6V�l��-kS3&����kj[a_Z]��f���m��jl�@��l2�lUmQ�n_n�*lʭ�kl��Y*��h�YōZ��4�Z�-L��i4�5��ikm���UL��ͭ5V�[[RV�ڥb��FZmE�Z�V��}�vMV�h�X�   �����ۺ���Uq��`���t�s��t{]��ӹ����;[�纼'�-����浶���\y�7�=w�n��޼׽{���w�sݵ�h���v��Ǯ�֝^��U-��&��&���ʶV[k�  ݸz@  ({�����B�����
(P�B�w���СB�Mv�|�����M;��׼�rn���y��m���=^ݵ�Gam^�Z��v�ݒk����^�խ=�ڮ�a+f%.��6UF�j��  ݾi}������^��^��ޱ�^���n�w�s��{���{��ⶱ��P��L������n��m��{�I�����sw=[[�޽燭��{:����^<z�՚�^A�a���nN�Y�Ͷ��  n���n�齷�y^{���^�����ݽg{�D�v��9�u����d���-˷����^�ֽa������ms޼�ڴs=x�Za��uQU�W^���J�y{h�%�EU�M�Ul�  n��m�ڽ�{^z�*�u7�z�e�]���ޭ�5Gwlq��W{;�Ըr����yE9�^�7�zm6��W�{����:��̕��jV[JKbm��eH�  1�綱�����젶R:;��(���W�rՓw5Z��o{�J�z�����B�����pڮ���G�V�������]���,�uQt�jڛX�fо  ����}��i�t�ON����=ڡt�w��j�kU�] 7/o=��޸�^��{����q�]��5�:h�g���[`��Pԑ3j�Z�cjQ|  o � ��W��  �W : ;C �&�@ �N�t�\�  z�^� zuJ �r� ���%d�L�Km5��C[->  s�  ��8@�}4 �{�  �]�  6�n  $�v� ��<�v�  gqp� (�.� 4w,Fک����6��m�4m��  9�@ c�  uۀ( ø` 9�  .�p  .v�Ӡ Sr;�P Vi� V�kJ � E? 2�� Oh�JJ�Pdh��MR��mA `O��%0056�ʔ� �	4�eT� ������_�����_����{F�_�&�]D�A�Fm�FFqm襧����>���U����r���IO$!	$$?��!$��@���@�$��!$��<���������?��h n�v ��g��aCwT��z�D J�t���r��L���K�3����XS���ѬAҬ��a�6�x-�N&��� �丅렀JWQ�"[r�7X�)<���ä��45�a��1���K� č� ë�$3�Q��:�Ǜ��
E%��7�/PØ�N�@Ne1$�5YmZc%ZrF��e�L9n,B��3m1M����5���u�LԾR(�e�J�l�f�u�5[��;�6��H'��������֐>SX�7.�Ō��/��J�-��{��w��C�,HQ7"0��wFi��.�N&-�*gd.ʒ�P��c��K�J=ʷ�^!��"��M2��w��[[f�Ǆ�	�{6YJ�R� 0K�u�ûZ�R���e!�lwBdfj���J�H���δ)a��5r�j(��6�;��n��P����8��tM��T�p�r�ڣoj$m՚�f�k^��Su�ǵ�t��4��Sb7rD�Ĺ��6�K@ܰ�^�eɉnL:+��D��#��[��*�P��x�v)����G�
x�K � n�*Շ��AU
ܰ�R�.�9��Zf��n��d�s��hu+%޲��E6%�r�k),���,�z�!$"J��u`���
]���[46�n8�(7%X�YX�zt@��bR��2����)[%̗X`U��p�@Rj4l���lcW��Ҧ*��c͊�
a1G���?i� �,v��ڌ^:G[�I^|~w��Jn���tJ���F�Su��&CDfeB�3��cc���+"�@J`�^�mF�09�����.��U�n�M�[uz�R�L�PX����ݸ�e�z�/%�����%Tƅ`{�+��m֭��h8M0�_En�\V.���O)c�,ok1����-GIL����ve5O���e*b�<yi��O�m��Q���4���j`s]�'�����\�B͹W�F�]]j�{z�e,��a��(����ּEjN��q�"�&�VpRǗ��B�A=)���xZ�a�(E��Go(n���.Ч*)����aM�pZ�k�ۨ�׉mt�3�nc���m�n�(,����=+qkT�Gi7P:*y��A�!��t2��`7�v8Ӹ/j�R�A=�YD��/k+p$٭PE^ˋ�F�u�	˂�^�;{c7#��&��`���SB�S"Ǭ+�8�%� �	��S
�"vX��B�c����,�p�e��2xi\�S4��+N��Xi5�R^|�]]!�Gs�3�b�XB�N���ie�1l��(���	��ݸ,�(�f�4+iH�m(�7`U��i����\i�#�z"!V�F`�t<-6>NB˻ɻ��2g��
�.�55�v�5��U(0�nPNTM�Qn�
�LU����Zw�j�R��`D7v�ffe,3%�.�f�����eJSf̫2u#j��Vc�� � �S �lj�]Z� �^��+7dڰ1�'2i���a�Y�l��ѫ8t���l���
д4�VV�N����q���B��)��]�R�(/6�U���-Xd���T�L�6�!P��u������<�c7��)XJ^����F�D2��p��)!J�jt��y��KJ�,�[���)Ya�r��HA���4�7Vj&}�ެXt��ВbD�Z���m����-�I*�m��/B�@ea[�K�N�ѣ��3�j����Hr�#�b1���3aXrΔ��7-Z�h	�,�aX#�b,�M���� ��+0L�1i.��� ��9�r�Z��8�V&M��)K���9���Md4Ŷk"i�6�� ���YZ�w��h�5l�h%�m˨8.��+X���d�[�r�;�wmR��*�{y�c����C\t���M���`�jn��s,���?&������uUw�si�GE��� �	�����Y��r�ܛ$)eX� ��.غ��/�/�W�����r���l![��_�ܩa��PP��)$w��:(=Ɔ�[��݌HeZ�,���(ˁ����ye2i�if�L���;u-%N�Y��u��`J��a��p<9`7ù��è\e����7n ��*?c�p4�-�h�z�[�f0�sB��Чn?���xte�n½z�V^�n��,���k����O ��k�SsS��yL��,:݌ċ�NB��#Mݦ�Zx�Ä�J��Hd��bf3m�Y��GX8�ź�.#p�o�Q�.ݣnՇ�퓈#��.�����Fn��ux"o��o$L�e5��:i�1F榶T��e����A�e�L���oi1��L�Rf�j44X4�=}�x�����W��iYOF�]y]��}s�cl��3�㼓fE�k�M�Jxe�E�a�9B�(3�R�灲�r�h,���!)��V"g� �Om�t�L*��c��In��PhD��M9��-jv�e�]©hM��ץٓ���7&#�)j�l׍%��0%���Z\ϖ�7�QN[�6�mD��=�9nժ��x�ݒ6�A�P��f�X٤B[����YݷO(�8�a1왈`�R���#t�^n;�a9d���T�B��zÛ�[X�����O��#,��f�*�����LI8R8��&[�]�
j��V7��$���� f�j�Y.�]eh�W(QC��F1g6hBU�hH�ݔ���R�����:$��&U6�ڸ[�y��T
�Eر�+!��ڥ"�REZ8�l8��|�]��5��!�%f]��5곍B
fm����4ѺM2��ܓv��Ɩ�
h�Х��i��(,U`-[x�ẃ��N��[��iƯ�z��^0!�5ab'v4�B2Aq�p[ҩ�$��ۗ�(��]�`�.���WN($�*Q:8���C�R{I�rl�>;-��n���>Jçk,TNm<��[A�q*�`�W��/E�Yh�A� c���P&��Lf�X��(R�F$�7N�d1fPsA�N��ؕ��́ �hX[ó�`�n�U��]��f�[�&��V�Öp[��2<v�Vmm��d�5�� 6��
.����������eR��yF�L�tٴ�KD8��A9��M*���h7��ڣJ�a�5��7���l���(�t/�l/���+w̳�i`���6u�p���@�X�z`�)�֊��l��0�����V�i�x����H(��C��֯&!yQ�J��Y�����{n�<j�	����֧F��� I@��J�D� �.Q���F�`��5C2��3N^G*=��TL�6,�w�b��F�Ҁ{s
�&��������ܠ��YM��KhQ�,��k:�(R1I�.b���V� �z��-�)�0)`j�en�ڈ�d`ܧkB�V�*G2���
�eK�%�� �/U�e%cs$��&��%J=T&��%�Һ�wr�̰֞W���n����⽤�("���7^]X�*�GM�,�@C���f������n��mւ��Y!��A���K{V�����B�p�ȱV���:�X�M !�އ&Z�MY�bJ���M��S�r�p�vcZ�;����U�2ݴ�ړ*c��mS�t��m6�_%�$o\�h�̊��n�u�5���f��E,�6���e��ԠɻD������ު��W`��keY58�%սy��[C��Q@'[��E�e�,7�1�E�ʑ�p<��8��2^:a�v2�©M��;�R,V*�-�P�72��� @�қ�5��4�K��u���gѶ��w�l;*�l��Ф7�G�w4��7�Ԓ�0�q�M��R�HǄ֤��W2�j)����Vˑ��h��N�P�2f�x�z�pD�:Z���i�[��L!�&���J��:ފ5wMT։�Zh������(�S͵6֜����1`�\�)�t�u���mǓLY��QU���s��w�ș��^0�1E�����@��6SGlh�FU$(�Z� �˘����;�2ȴ��*;2p����Yi���#�9n��GSSR6M�,*�-39lo[�Ev��LZ�p��؆�ֈR���d�Cg�t^�\���Y��EY�Uz$v�j�9B�Q`�&i�
��T�wDf-��X��+�8�C@&"V�$oTasM��̚hM��4c��X�V�2�i��q"r�n�W��tҫ��̗�5v�Yp�-�l�n$�D\����
Ula[��iL��TJP�U�r�k��էR��Wm����íeGW)a�iT��cE��ybF�qH����v����"���wOW�S ׈ƅ8�Ue�/v�Y�`j.;$]e�&��#�B��m��z��hT�6=T���7\0�{K>٨���-Q��f�4���flYa;1�ؙ��St֐�o7.^;�
CjcVY!CcuyV��6�٪���%[�[����,t1��D;�yd;M���(	�n���Z�JfjA���`� AXK��I
��VV�f?�8Y͖u��!	=�8  �#����<�Phj��W���֨7.�&t��Sk��������Uk/U��bm]'�a�n��,k����fabSdj�&�f�m�:�x��F�WWf'�M�[�if�j�wx��l�ڐn]\Z	���v2�L�6�ر����g�,�C��׭V�&bݲ�T��u%j�@Zd�t)A��E,,j��n�S�mU�Wq�h�]5�g*Pg2�� �1R�˺J�(䂮�<�����3!_%�0L߬յ�-��w� �s�(�B�ŵmQ�)�Kfi�n��/'U�Ⱦ�W�PTX^�`Ӷf��a���#�زRGt!(��)ރ�����D�H�lH�f}+,��T�%�HnKN^���M;�pQ&��eelHam*Ѽ�B� ���(4TZ��l��=�\�4n�O��j��C��WW���P\�;5�·���X�:6eViI����(�ބ��t^�w������5�+(�k�v�7O)�]e[c`�N�!O-�wA�i-J��VV�z�!n��,-��n�PO�ᔄ�1ڱCB�w�{{:�8��z@m&���j�{�q"�d\��h��[z��h�Y�l��E[�Xcp�0����ő妉�y�SFЂh܀\�alr�cd
B)�u{6�^L�/9��Ȭ�WH��iP�,0۔j���ʴ4��V��Y�;[�[I)0)��V54�.�5�oZ�X��L\	ύ�b�.���^/�!@�`��x���m�6`sr�Yq�e��<� ����˚�ϥ����d dQ��Vmj���fQdS۹CV�Y��ІL�$���m�q�R����9�t�U���؝;���gi�6�W��c��op<[	hKZ���o��k%*2n)�	7�pHQ�b{����Yl�WWT�`���%z���?c���`E�n��Y��Y2ROO[ R�֍f�	�iN�d��^�����$�	��lia�L�RFҶl�$Z2���
�y(��^�KƝnX5�2['���+��̺�P:��e��ֈ�����/^��(���51r�D�ҊG���M�p� �H���w%���j����czlmul�e&Օ�jW&�9L��4e=�@t4�0��X�%TGj�qJ�ߋ�h�f
��E��j��/&n^�.�[FZ��)
Y�i��Zy�B�rQKvC,c9�ۆ�$B�S�-��o�O�F�&���!mMD�+F��d�,×j�
+Ť=V$���^��w���Ej������>�Ѳ�a��4u��`f������^�GR�1î��T��Fө`y��hK�K�5d������VF��r�Wtж\n���`Z�UȜ	����7V��e�p�O�e�n�85Ӛ,ջf�Z�m�T�{w�n1��[�M�[���vC̡yI*'*�3u����Si޼y�kE+�'�f+� PQM8+&4:ߤ.K-@�t&�ttFHsEd��JbcE�y3MZ����\����p0ފ#U���/KJ�;��G�v8kK\�4U� �ԉ�E�4��a4���A��
W�D;N����-�h�M�p�[������@0v��fш�ml���i�%�
�8��YSe���\��ʹr�ݱoZʃ��5M���bf�X�iHn��ٚ�bT��b�J�Z��	�yNặ�����k�i�oA�Z�`���`�u�S�X�)���T�Z6`t��˫�p�amˌ�sQ�kp�W5�[�*���WJ+�cD������-I��	s$�$�pDkb���Mv��0��8��F�Ywd҂�/�0��ӶhI��T���K��L���t�ć�ٻ��OV7y�*���i�j��T�R�҂4�֦�l��ʮ�,�X��͹CMՂ��4ù���*�
�NY1P��7��*���B�&�uo+�z�:�sV�wVۛ�)!P͈3xT&ȴ��W�3p�x��t��Rf6l�f�@Y.�Σ�weh��.�S�ND�N���C'0?��6�2�f���:��H�W&� vbki���̽�-\؍"��ڍ�Y�j�Jך]"	��Vy����V�ݚ�JE��]v����`�p@)5��?�²��/2��h�nջ��'+ohS���Æ�)JZ���Dؼr�N�:�FYȪ+p
q���#�n�b����n��B'�kbV�j]^�u+�j�4���6�*�acea��^�v҅�6m��Y��ș�0;t�-R����[T�j���ǭ��a�v�\8ڷZ�7��=�4��+�a��nƶ����Z�W���Q{7�Ξ�O��=E	� *Y��\nȺ�
�p5�Q\���b�ocMs+u9��3�tQ���X9&��>���PauH�NQ�^����Qfh�3�z�j���f�kb�٬Z����yZ�]������E,c۷w�P�G�18	�0=ֻ��>��˔�G;m�-ܙ��"�yǸɄ-�W�7T����4S�u�m����W<z��F����j��p7Z��'�q�7Wx�4�.�_1%yf�ooˈ�I]�)�|eya���{�+�Q8~�[��&�t�ܤ��\5�G�3�ef7.u��:�q�jf+ ��f�[���鱅�4CT����=����Y��1I��`�G-jY��UjY��R�]�lr����ARgs�gn�	B�M�6J��nC�į4Rw��
�wah�%�|�֐6��}���5���>Y�Ŭ7��������n�K%=��O{��ػ;�=�6-T�ӨI�X�8������s	��*[��T�M��̶hp��uТ��=3r[J��K�,<g3e� �[j���7�j� N��ɸ�8�Q/FDB��z¾��&ron-6�5B��G�3d�&�6TR��]�'SV�!�����i���g]/e>��Ӫ%��L�Nܫ@>M-����E�������]0Ό�Ƕ3���.�_�+��R�8��9&ErH�c)�:�ҚnYFB�%���ϱP�xi�u�7�g1�G^�{,�ՙY�Q�Xm��5H����M�z��n��]��7�Ѿƚc.�и���B.ʓ��ח���;X�I��ַ�x�
z��,��2��!���ʻ�3E��ӷ4-���ҩ�c�]N�`��;C����e�$�|�ҥF�u`ݯq�~^ͭ;�9�/?XD� &����b�Nإf�Q�.֣l�]�XO:�.�h2"i�}�2�]�ݸ8�q��2JzJ2��:s�k���\��E]m��n�W\	���Z������Z�fwnd�^
���ke��1���qv�S%��3"W�ZK�q��ps9�ux�fk�H@�GO\ô��b���(���ٙ%�����*S�nm\�2����'��ؐX�TH
L�U�� �%_.��}J졶V�zȫ$���P ��X�Pl`ÁQW�n�Z�k*j�o���^.��)䌻�j0+��\td�p�=WM���!��#�,��D';1�ɵ��R�I�����0H�7]R���2wkG�R�yjP�+n9n��eK�����Xµ��%�Mrȶ�OHN�f[��oEJ��!�޻��z�9�Z��9� 3y�ܳsb1�}ad��̷�C�p�e�;�R�|��,3��ue)��E��Cpɤ�����bh��h�U�ʧ���O~K��s�;���*�{VUHF2(A�����|�J��|m<���{`e���ݠi��Iـ�سp��j.{���_,ΙΥna�8̤q��n�3��0n8�Eg
���:�oUC7s���V�M$�7����=�ܧ�eg�\mn�dF�Z�g���Uͮ@©62��ot�Ô�ŵ���OstM}�=
ڦ���RcA�ƃ}��$�K���y�'�{	���YR�H�iWo]��H0Tޙ���Zt��Z�ٓ�E���u�����ٜ�PI6�zA��WwC�{.�iV����{4h��B�CY��o7]�
a���eF,��[�ߺ����$��L�X�[Dm�.�k�HE���;�(���P�b��;���U�w��S#�W��ٳ�]�����PH�z��q^�p�tq�q�7EY�s�p�I@���6�z�]н�vU�ǃ��ؖ��][��e�d�)!\j�ѧ/7C��(��e%KT����,��:\�(�r�m!b�1V�WuiZ���!3mI���]��b4[^�b����A�:�����F{ HI���ۊX�ɚ�ݶ�m
�f��9��x��4p��'C��}R��F��U�6���)��§dcݍ��e�F9`�����U�V��>��)AJ���##%fptNhU3���ͭ���aJ������g�R5�kq��wԪ�ц�9ڜ9�D
�S�V��	��2,[�⩉D<�{WWj�(	o�uC�׬�a��L��B_wY瞁����ώ{5>G�K3�%�m芉��:�n�B�@Q��rgd�'��7&t���W6�P޻�37Y�H�e�:�*tk*;�-6�u�`K�\�q��ʈ��@r��vR���ɖ$Vm����u:�$����H��p���.��q�w���=���r\�m�Ő�-pK��H��̔-6|��91��'+Ě0��D���۽4=Q̀`���A��~[���M�jA�W`�T��C�%}p��cn��Vbl��a��-���~��&oc8>�g�&�3黴��h�GC��,��&*.�����6N�
W!L �9�gU�m�t���V��.R,$����7*����� ���W�������+<�� �RFS߭�Hc{u�|�DtsB[�^�g7���Գ�P�
-�y�%�-�z�p;���C{���zJ.�)��+�t����6��]�3o���鏫n؃��쎖k��14(�e6�u�w |/6�j�+��+��؅,#]����n@�f���.�o{+]�|:�aE��u#: �R��ހ�¾�G;��@�*h��ql��}2��6;�o�F�.ki�|�]z>�)+ղշ �䚵q���jr&���+%����I/�o-m����闪jH�mXLW]�b�=tx.���.���I����=���E�c������Ff�c9�[Q�l ��[�.�r�OM�#{u��]x�4j::��5���usm%α��wKn^�J{�6��լU��s՘;'c�o0�ZbK���y�N)=���+��r��xm0���I��zL�޳��s]��������5E� {W�+ޔm�w+	˙���i:��5r4{NQ
?�+�9m��G��������9�f�i��ro"33UR�$\n���.�D��GZT\�z� ox.Z)�97J��ݣhrx-��cf`��J�rݧ-�{�:�/o$�b�������Za�!��Q�D\��WJ�њ4��5�И�.D��γ�3F�q<�<�<Ģ�)��A�N5f�ħ��&�	K�����-��oI���^���R2��u����](��d49��񧒰���J�q��(�`eY��uB��v�u��l-j������v$ň�V����2�	Ku8��v��i�a���|�Q�G��M�n�;���4/.�6<���ah�A	��d
]�;�{%O#��,3�\�se��u�YLS�&�1��:n�-����ˢ����l:�9^4�Vҕz�T�"Wj���w$lc �4wB{�����>�Gfe�V��jue�]Wp�SU�l�1Ǻ��>���ϔ���`���R=����D`��p�XE�\=�t�6�ɍ��tt�l]����F�f��~�ô(u���IJ^)@��;�X͓��0�J�F Ŋ&�IQW�gs��8˧����NW�wm6��m�wd���:-u�oi�_�T��ն�p�r��K(e��U������}P��7�IF�8]���I���;�X�f�c�a:]ۛR��3�.��Jj��;��g@��]�a<�V��/n+-w���ٚD��"����
�ǛC�#e�&
Ù5�;\6s&�]nAZK��}\��ACwR��&�c'f���f��B+s��ऱ/��k&uV�����MIȚ�F����U�,}��\zb[b�u���t3���S��L9[jUŶk�m�M�y���X7�H�2�1�d<6�[�MMݨ�nuf����r��۸�\-e(FrgV�8��^�Lgs�mֵ�M�hǺr���W�		����m�f*1F�X�l$�P�����n\tI ���뜍R���ޮ`c�d���1j^ i�"�@"r�7��+F�Κ��1i���gsD�\궨bB�.��ȶ��w}%��N���w!׺��ĞSN�m޽~����kh�!�߁WQSrƺ������Q�
��>�Q�m�����p�0^��v���c@u2:�֍i�XN��V��^�8��:�XU;�2�F�fT��k6Kʹ��	w��|F,�㫢���n��x֣FZ�;�u����9ur�w#�;�F�ȕ��ҙ�y�g���M@4g(͒��A��6���dOLI�͈�')�;):Xܺ�If(�+wkۺ��v�%B�7o��dאe^E.p���e�Xݙ�mt׍N�\���N����3.od���& Bv>��ɒ� r�e�p���gHL��y�Bh��5���%�Q�v�kq����6�H��ax�ַ9ځ�1��'l�P��s�M��&j�����:!��&�l���v����1c�B0�ru1�2��x[9m]b͊;yv����X�ԇSD���L啦3.��������D�ܲ�5YO�ĩ��]��}VgM2G��s0�T$|6�%��(��;�.��<`�+wbu�mti��7s����i�8�w��C.�ĩff�B�-{3#�A�w��$�S��ruf.ɉ㏷�Cs�{��J����G�ʻ� ��;b�Xx��M�9��Z�=\��ǝ�v�9
$Y�����%B,�l�1�ozk��o����i��aN)e�ҧ2�U���c��+/��Ł�ڎ���ȷk������Jy%��'�'���v��}X�Dv�CZܫ�pc]��ʛ0RV+����v�	����W�u���@ƥ|;��sSg�Oi�|;OH)��)%�n)���kYʌF١.Z����ڛ�-e��41�FGt��=!�O�S����f^�A/Q��>ų��֍��78d1�q<J�T��7���&��[ٻ���-zL�˨�_bSk{Z|P	u�i�CP�ȍ�z��)��lw`�q��D���9V��i!K�Jt*.i"]�w$�{1�b��Bf��j�n>���l�4r�ũ��ۼ�p�+��f��{�ϭl�Хd��A���QK����}'��O&t�K�aW
�ʍ7��X�Lᚌ� s���:#�� Tw��2��{�������!���.Q3ʳ�X��� wYpМj��V�7`Z�t�iQe��0�Nsl�/CG�ѓr�BUAQ+�>�A�v�^�9�"�L�;�{g��j��{������e��{�	��'W��6S�	����+�=��x&J5qQ��/�K�Ŋ�8k��b����P�ю:W�-�g��U��C�%;t
�7�@z^�6���y�i���"2!`wkn�@r���W�I�^����iɇl0��@���������+��l��ͽlhx�����^t��y�;	g���h���m��.VH�%^�ƕ�Y!%a�B�x�N]cfu�[��sիc�e7��xb��x5r��e�]�6bG9=�y�!Ivw3��K35H��[�,!0p�'���q��g�W����J�0ܦolK�oi^�Zu�J�Z�L��#�X�C����PHMe
tz�T�(���u��ni���X�n�����
l��$F�9�Ԯ�Pp���aulb��&m+�îbx(gj܂P��a׭�s��m�.���;E.�Ɔ,9�������Zz�k��Jn�o>@�t(�=,:�H"�خd��r&�h���fX���D��*n�m�6�?Z�ex��,��'6`뻰�L��pIk-��b P�9N���6�i�Q��T��n&;�f�A�-�d�Kd���Kthb& v�����Av\����q��'r���1�Sbfp4x��m�v�4���Y��@��+ŉ���������h#{��φ,����G�N1�=�<�1:�k�[f�۵ָRn��}xˤ�Lݐm*׭�JY���Y�!��W��#����Kte��f��#���s�1�Z��R]&����5RF"�����2n����T�%֞�L��QYy���e:ɪ�����r��Ԣo�Ԙ����ܖ��"��U��jӜ�W���6�z�ۓ+mr�Wtn�b�-�I�YRk5&rYx�۔����4{k"Zgf�x�X��ǳ �-���mC[nf�z� ��K�Sr����l��#v';Z9�'���n�;�Y����ep<u^8��.]��N��M$4)拹W�#R�rv��U��T�k��,�q�Q�V�m��BR�9q����g�]����a6nv&�Qݹ�q��쥃l�p�����n;K"�١Ô��Ù��^T|�a�+��Fꬍ#{W�/锳�j�5�5���
�����J�̰�uX[Ov��:g�U�k��쬁�{OfP�)Ve��c@�{xH�%��]u֌�¤�O^�������� }joP��	���ܙ�4/��e�Y��-�O0�N���r���qRa��#�%�&�J_-�v���T�޼��`\ӊ�1��NG����r� "�i��R�9�K���2.ъ4�u�=�jWfҴ���Y�]x�'E�N���P���J˿%� �dBuh`�o9��=�FR�$C�2^�8i"���Lvⷷ���Mٳ";Y���Z�;�#(�k�Z�9��a�y\��xy��RAB�1ƳGpqл���֨9f2M �gu���Mv�X:�;�c�C����sp�q)/�V�@��nS��V~}q�!se-2���ά��\�%��͝��βʭN��s���6ء| Wѳ�
�|ʋSѵ�G�m���I5��S�_H3:��ǌ�妵�K�B�['moo١�b��ƣ�|����z�m�p��]{�:n\�z���� �h�YW�6nX�[2,���x�j��}���x���?��BC�I|�^k�Y�ґ:Ĥ����0TN��˫��X�IF��������C�S:��H�|�܏x,6�}u+��|:]�Q⋡�lmm#Z����<#��+���&Քe,0^���7l4�X���٨�5�ue�Ǩ����es��o� � P��V�"��*�������Z�y/lS�2;�Yh~��u;�ܧ��D�k�Wp��k�udѼsw�!+4G2�jٛ|е~��t��[��Y`C0�,���ƫ�و���uૼje$��"��d�U#}Y5U���Ȱ��ɺ���>��-%W�y�- յF��{+2�k�i��B����'1�-��E��
��_�h�.`�s��m��S�^q�ȣt���֬����J��7����&M��>\'^����NMf9��R�������1�:nf�l�A�ٳ�mi�t̛��I��a)=�/�ẗ,�yi%1�4��Y�n��,GA=���e�X���ذ�z���1�s^��Z.S���T�MH�`��z�z�,u�Cw�pKyz ����H|��I���K~s.�F��믔��V���(�]�+�Z2�e��j�i͆��U�V�`�92�D�WL��$D���b�����iZջ+v�WTÒp�T�3F�*�
�7ʎ��0j�3���2�'�ql���]����{�V�7��d��]03o+UL�nOm�*n��/a뺚�Z��� bԏk�{��P}��(v��R�=G]�I��ԡy�jT�b��a����<��V�䅫�i�3&�y�]�e�.������ըv;l}�[4�w\��tP��u�g0�rQ	cFh���E`���z@������SD,Y{u���r:��.�����۬6V���W+*��s�P-@RU�(��,r�]:$S�|���a�����O~�8R{�]7��ځ���*�bj\��v�:���YŢ��:Zfe_v�ڊ��&u��w.f�2;�W�O�haTh��X�᭼N�V��:�&�GG�T���Gh�J�+��ʜ�o/�`V��au�kA74��'B���s��b.D�{�B��0���r��[ś�|
��=c��fwj����VlTPع�̨��zd
�*��a B��ۮ�����6��2�;ڸ���JД�	(��P\���1�f6DAga��ց/�je�c"\}� �F:Ȇ�����W4�`xx�<,tvɄ�q��ɛm?`P��b�M`+^�s�j%��r���6_�pń[�s:��#��4��2N���3�e�ǻ���ۇ;%�yl�q��m*����9��\ ��L4F +�;�寵�:�ɔ�+��� A=��|�n��c���C��Ǵ#���L	�v-yҡ�4�^E��m�T)of��bBǋ�RLn��1�zVm��B�z�_p���#��ػ���b�{�ۙ�q�y���*t��J�n�Rg)��b_V�b�g�;�r��v�6EǍ�쒝%eY"]��!���ݔ4������v��k��Ҩ�gU��ތ: ��[Qћ��� �[��e<ճ�fػ��� 6���]��uIfp[�#�$���ѭQ�K��Z�v���V�Yv^7K
Ts2d:��淓ǝ�l��M�u�X�����]�GCv���1=��r�xu�o^���+%`� ʫ�'x�>s�����)-��m���f����d������L7�T(ucz�+��Ҹ,	�6�`ۭ�$�`�Z����7n�
G�n����N����� ^P�/e#�I���HU��6D��#�J'�P|��,X75���]�i�%W'Eѥ �I�0�O2��[˴`ʆ�WPY7��T��r�):*�T�Z��8�y:#G8�೥99ku��#&m��+��L*v��
l:&��7l�c �R���[%�}�J9��A�� ������@Ծ)�+6QK\��wG��kF[7ֹ��FN��i=κ�mJf�RhXi��SU��\+�2���]q�\My��X�J�̊�>�_�en��%������1�U��� ���s;�\���3¹�D�
��Ț��3��|�*���*�� LLH�t�iF�M���վK-1q�XiL�*�fy��&֠��5�FX޳,�Q1:��v�K)��3�����P˭��Ò������+�������v�LG�2�H��l	K���C3�Z"5�]�ػ��ԫ���h�<��W��[%�y�o.!R��qFep
.W�k���lS�z�ʒa|�&���n��/�����wE���o�gj��>��U��2��5�Ʀ���Ӧ.�&8-u�ⷾ}@�f���n���Q|�]���]w�yO(� 3F�.��mgcZ]<i;��J���gp�#[��	@Vˬ(d�j���z!M����u�Q Ѐ;�i5�o���WQ�VnC{m�r���!|�[��0ҍP�Σm�i�{L{O1.啶�F���9��q|zn�.�k��U]��@��օ���E�.��oM��o���ij�R���8�	�]w3y���[� �mip5ܯ���̾�D�N̙猻֍��-Qg�zb�"��r� �k�sw�Qԫoh!� �����h�rZ�y�"oK��d�g*R��zV�^^7@5�x��u�r\�Yؖ��X�0�����Y��^to7�VemRE#H�@z��i���B��n�4�3g�pb�<x�Rh�C�f��y6=��5Đ���*�r�>ͤ�1-�ܧ��@�mX��Ֆ��Z��pM:[�-�m���4`5XS�˨�.���zJ�3������y���M��8��ۤ�B�����=�Z��c;
y�u��!2�Vt�1Su��d�w�Y3b;6�:���[�4�V�a\�����g��x�_h+ �h2>�WN�p��#�KFB��cTi��|�]��6�U l���j�0�rJ4�̋fPbb��\�ĉ�>+Y�\���MJ���:��ǘJbf�#x�	[Ze��/�8����N���q�J,���W[F�NkۭӋ�q����7�AA�-p�y �����ʱ�oH��g��D+���4�'Bγ����SHQ�}&k��X�5������P����SoV*�gU�(
e�oR�2�.�9d\y�n����[kU�p<��S[��w���D:�T�Mv8g%n�V�� ��ں4�P����V\�g*�ʖ���\�n^7�Ch06�J��#��f6��i[@�L�D^�����2�=EU�������M�s�%��/8}�R�v���4-T���n���ס':���z�I�YGm����.�E*���oPX��Y�Q[�Iܥ�A��[��L�M�d.���+�\/d��x�KUjU����k�m�J�H��m��S̮ȕM��:��O&iR[3x\(��c�s��`��K��4'h�w���۫R�ѷr�!�,ejfT�%��{ۧ�R.���]�ʁ��]���/����2���h�@��7Q՝HءS]�:P��v��*�r�d3�uL���3%��&�]Op�=rY�]����]��D����h���ᶃh�����˕N7��ݤi0ތ�(e
��R�Z��H]YS>�okP��'�Ԭ<�Ű�f���2�r{oUgWu�i���5�2�6ŭ0hv4`t{cat�m�)(ނ6^�n�vi��N���@�fP��o*]8��!&�;2�X�_f٭�i�����gLx� ���9<�����+;qm�2�P�Qk�C��d�NN�؝�A�L�;�-���q;`F������b)޹bƢj�</z�f��Yx����5,K۔����hn�Η٥�M/��*YP�c�Wsh]�ɩe�Ro�-m�0�6Ḉ.n���4�u�%p���]m�uEg�Cp��T�Ӥ� �ߚ�0�o�z��t# �p�* i�o6�YΦ���B�z����k�㎖nH�O�ej���ޣ��ɯ1,�6��e���{BRj�9|MЦ� �hP��6�Y�k��m���N�R�6E��6�s���-�fvN�k��к�Zr8;JW�l�7v�i�2��eZّ�/_J �x����|�\�a���T��Ǫ��7:ژf"�`�p܁*`�5`�.�,�ʴ+HRdX���G*����]��ul-��m�ʧ�rJD)�"@�����s����š�U �'��`��5��,�U�QIQTg.XCn����WΑY�W]6n�)�����O���Zp�}:ny���`Ž�r����$FM{�/ݝ땭��f���+\t�����o;�.�#-�S���s��վk1��5a�B���ƲG8�1�L�FqsB3.aӉg k����K�����e���!�8.x�]�X�tc���K�V %�nP�}X����jMvr$E�)ջ�X).�T`��2�j�tʎrH���yڣ�jmmrpX�Ó{I�r�p��Z��3��Nr�[��S��2�S˽:�ؗQ��P�O-Y�J�l:0�f�):�� �v&R�Ŷs��Mի�;fEԡ�&���O@��Utu]_Պ��E:v�	Z�N�1�9�� RS�V:�u$ݽ��^��r�tf6�F�R�f�ܻ&vh&"֯�֭n����.�U�ȩ���S{h���sE��_�vz��S�U^ᵨ)��83�	��є�,�d�J�J�U�N�-����,^�]x!ܹQ��*��ݻa�TIj�6.��N]�z���z����r�+:�̴���Iq5v5َ�%��#S�]t)!�%�{�j	�jv���FR��ih�.ӀS��k'(�tq�N$�'�N�=ˬg9"e�:Y.Xm���5�ZgQ.�1Ч[4T�ޣ���
EX�`��Ha�R-��Y�l6v��K�:��X�3��~e�x�4	^���wv��_���di��A%���b	Ѹ��F��!�����jJ6�9�ΰ���Li�<Ve!	��޺�7]6\���7r�nr��P@E/[yR��-��/!�i���rfĖ�.���ӟt��w5K�;U�PS�Nt����v�c�z��	&㨸�����`[/��� �O+OmJ��v�)z�1VP{s��Y��s�i�u]m��8��N�92�%^��
QӦ��6�섶�2��;�M��8�C�+�:V��-�ȵ7�[@�;v�t7��)�g\9	P.$䱦ߐ͆�9�e�zڧp�����'��ak����CHO2��}�V�6R�#{{¢ܙعE�vOG&�7�ºYJ�L0�7FN8ڙ0Ќ݇�u�z(��/��$آGF�C�X�*��nhwR����-gk>ZU�9��H6�7J���w� ��ΦX��Ԫr�3��&��}3I޻�]9�\��T;فo_0�	3E��)�
�u��֭�;�:٫ 2�ݬ�y@u�8h �>+��a[wR��]M��ΰ)�^A��M�'H1���uzLҙ��v�׀`�[&s�pl���oq9�j��SC�6��S[��,��3���r�f�W����'�%U��bK<]��]�ԥW��K8����v����X��a=Nxل��������߭'}�݁� e�n��5(S#ܩN]�[�0c�oƱ��t)�1�oa8.��[����0J��o���lC5�f��D���BuZO�o�>D�B���jS�kT�]{T�j<�٣ZB��׋-����u`�/����jX� e*vo]a���YN���,�����K�[��.̷B_u��񧭗-�DfdCA{�v���}�Y�j�NÊ�n�YXH��bX멧n�
�}�yn�F�2�:�f %Q�i��#��ʶo��n_B��u7h�iIu�`�wz�'�٣F�@��c>������������V��xcgd�P�b���\sl^Z׼�#�����S{E�c{C��.�t,^�ܲ+�n�V�=�%I�f���b�w��j6{L�3��0I�_ee�]I�mk�M���Azꛦ�S�ʔ�QqQ�H���X�OXN�H��ެ����u-O�
��5c�ɐ�/�݌2�q�Y��e�%[I\�ʵNe�I�/j��\���d�zw�����`���]-XY�___�4����8�Y���0�-Ӷ�&�Rb	u�{� W�(I��������悤�aB��F�Z�e)�
�Y{�5�V+Wh�X�g��Ը4q�ˊ���Q���q@xr�˳P�9��!|��eB8��Fh�iV�]��^Wc]t+b����I�m�;r�=+X��Z^T�,O��A��|�e�����֭�W�f�������B�V
�	o��ܬ(st%���[sV�sUV��J;qn μ�J�
=X���@���鲍i���olml�Ѥͷ�)�n�[Ưu�񻹯�
�)���Z�f^v7a�ܝ�Z�Q��Z��n��
�.:���@�nh�1�Ү����7����jw�m
:7���O���aúkK�����I�>ԣ
�����¥_Y N�8�@���+��o��z�nw'��PnX�0z5�N��Y��f�i-d��CD��]�P�>�z�P��Wң[�$��R�6���pf����G�R��ս�$�j�.�y4z�ܻ�vX��D�x�h�^��8n��x��f%��Lg����R�ͺ�X;�l@�����V&�儤��(5��k$-òR�g����p\:�%4�q����\�������݉���Y��s��Pץ�\d��(��a84EJ�u��VU��J�gWCۯ]�	ê�Ǣ�yr�Gvj*f�.����"�GW��=���y�-T��v:x�2{E���Ѻ��ݍԟ&����>��7�bw6wXy)�.�!�CΗ��7A��'a����5�.�\�e�\p��
\���r����[w|���a��v��Ʒ�nԷ�na�+L ����:�(v���Z�CF+�<0E;tٙ�K��o^ޗbz�_S\�+]�ۭ���ώ���c�e@�����h�h`Hq�+��P�d���l7@eq]�Go���7E���v՜����xF���7:m�]Mbs��������z�4�m���x��X�Y�ĤԺ'[@v�9X�՝V�C\���L#�� ��`K�6)nA�.��g��s�n����r�T��MD�˧/܎�ͤU���ul�n<�w]@��ia�ыn�1�,bpt�tRc��s�Y��M"T��
iVvc4�n�s��)�vy]��
��H�'�h�ѧ���-�{b��9	@�/<��AVkՓ!J�(mY3�Wǋ��s���։2�Xf�w���#�7*��M�J���Wwm�eY\��moc� ����`�
AÙ�r�V�d�S�q]YM���W V.���BZ[r��9���.����B��Z�����pY{��N�-\����_ �p��g6��/m���H�ↇa;Np��kemƺ�Y��q1��r�����"��@�)�>�n�y�w�-�����7��5s����-��k2*����}���f��T�*PX��P�+(�*)
��֪ ���F(()ic[&Z�
�V�j�U`�X�P�T�
֢�T��@+�J�*IZ���1�"ȹj�ADH-AaPP�X,+m
�
«kE�����S��
��Z2,�lZ�� cd�(TQTr�&*A�dYX-j(,�*E���6X�
IXUd���**�`��!i`�X5i+im,��eIP�lT�Ҥ�B(Q�b"�*
�,1���E%`��%J�**�b�2�
�5�PP��"��
���AYF�XVVm+V��E�-�El�YZ%E��`��ł$���VJ�TZ����Ub�e�Y��V"��Ta��+�!X(
�"F!VТj���H*ł�iX-EQE���V�������T�,�j�Q
ʒ�6Ѣ�(-����"���Q�(����EX���?���Z����n���;�iN��@\JNP�-aݎ�����L^�师O�mv�g�����<�V�W-{"�Y����MY���n��Vg!��cxP��m���*˭{�V}ָ0w�n�{��7|^�)���̗��dC� �j!T�E�a�@���}�����Itî T�c��]L�^���:���2O� ��u�Z8	3K%h,F�T(���8�ײTi��\f���森��kם�E�۹��,��9�k���Õ���Z=����Wg�-�r�kxU,-v�g:4C�9@�D��&;�`q�r���Ԟ5�*�Sʜ#}�'�ߤ���R�}-��B�׺�㲘�a�</�p�c�!�^��
NH��m���7�{��5ZW�ʖ�+ƶg������b{�v}H��b��y�0D�����Ǳ9d�ȶwps����V�s;�۳˒�H`7����<r�\aٺ=��w�F3^��qQqȌIטp_�di[ˬ��0M��<��S��b�K���'��� ;�T���]¿�eb��&F�D����h��s6�SZr���<^NS)��
+���
9�Zik�Ip��W�/K�3�a��4��ȅÝ+��,%IZ}�3�9��3c�@v[�	����`9'��W&T�U�*��9��{�;Z��C2��-�-Y�Ī��[ϮG�y�;V�}��j�r`�n{`O-l��+�(/(��P���{��rWlr��R��V=���r�x4ə���xߺZ9�a�m��ӯo\�l!*����t��7yLhUN�k]��+���20����.�U��C�U�q=�C ^�v�����;K��Ɛ��Ij��%���eI
t��&8;���Tp����G_JT<�bj�zz�S��N�Ql�S6{�Ā��\"����騯���H��5��ұVPL���=�6Z9noJ�q[ӽ=!���S�z ��ٕ!����8E(xp��N�����ȀB �C�pm����%��7���_>j��S6�����:�MܓV� �.6jP��$!��i(V�WH�y-����fT֞��o���%L܋�s��©�vʒk��+N$tm	��噩\��v�{�D��GI�a1=�þUd�a�S��OE�zZ�b��.�!�.�����d�X��lvI��;^��!_�C�Z�`�E�� V����)�JND9�6[��!;o������P^鞹�}�灂�h����>�W�$dPٱ�j"(4� �{�]p`�s-aÞ.���2�x��� P�죂��h�����5�4+A�C�k�l u�o{�q/]���;��T�[��њҥV��}:v���Z�)]��LC;�����@&f��Yt�؉ٙX�����Y3p���(��:�n�Z�̬�`����SB�"����9 4]ݨ�:�MN�V�lbWpΧ]FE�z��-�6���h��¢����2Z���Z\dN�-S��um�6���UO1V�,q���U��l�NW����H�O�GG�V{*�-r���ͪ�Պ#q����#:}lN�r��+�.3Kv��e7�w��6��:$�]��H�[N��̜R�ڞ�bz�B�Φϰs�h� �>4'��XOl���GFW!��Ik���N��:�E��qU�Q�(��K.�<��h�ıc�蕦/B��E1����	f�^�������OՈy�*�O�lD�\Nea�?p_^��x� �K�\�X� ����.s5�1d��cC��Yw ��ϥ��#��\�/qr�x.���.i��L6A&dG�To.2��ǜ}]Ȋ��2ztBWy�B @�ګ�F�^2��HT�N�t��'�P�/v�\ҙ��=�EXu��+G%�ѐWG��3�k��T�|�q-�غ2I���ؖ�<�Rᐡ���E�!FPIڎ�t���n���@�M��� p|���<a+�vJN�#Zé�T{Ý����5�l)ʏ@��V�[B�6�IɆe�:�Q��e0nv�N�8�Y��]5Ї�6eu#%s�<VbۮاG��]�M���\�KʔV�|1&��p��j��޾�~�$MoP��R�w8ҍ�)"�\�ϼ���(V��^���C:]Xd�j�o٩�`��w�(�vU���X���W[�,t#"��T��]���;&gY7[��p`�%p��(�7,��3���|oǤl^�	����H�kt+�ax�B��B�x<;����D���8j=�2�e���L1~4��{:�/(�Gh�z�O\�UC�k�b��{l��jyn!/�Q�W�ڷ��+N��� sf��ޗM���pu�1K���b�b&͢���o.TUP6���������/�&�mJ�������"E��j�ɘc Z��,vj� �^��s�m����nQ�4Vn�]fդ����N�b�eL�F�Qb���/6����Q��]--�n�(nJ�ͷ��z�0���p;��n�[�˞�\r���"u�V�Uym�L��yia��A�"ky����*�:�O��f�����z���_�`��>u�N�ӕ0t�tߝI���S�y�ϭK�e�d��cv\��
��q8 q��{V�(���ݪ��GS5�-�ුݓ�e���4 :-�1�M$�u�N���xJ�{����y��ڃv��|,�# ��
���v߆����H�J���.w��Lη����#��9P�r���䢗��P]`>����
�OvY��;R�g��i�t4xh��N�1�\�h��r�+�9*3��\���"�-��$��[���p.��'��=!��[N���4�j=���/�1�e��T���W�����݄��A�<A��\LO�GC�d�1��4��j� �ȍ���z۽U�r��QA��&`�J�t���ְV
uD�$a��>׌�0���j���h���FYF���n���Ml=kpw� us�d,i
k�m��u-����"���|��U�zn��h�6��PO��͛���q�����L�,��e��B�W��q_�|M����;ח��R�^��'���s��UN��>��p��jJ�
*�gk�չpy��M�"/�\N��=�6�\p�NGɛh׼�1Fz�1���ӯ2bTұ�t��c�I��Y�,X�8j1��e 8JrBY< 6��ϲ��-��t)����7��>f	�ZY4OzQ�u/{ya����y,�':L��T,�=�ER�5nx���]������i\ty�S[�gj�PG-m���g�*�.�Ŭжp%�Epd_u�{K`��[�ژ���F�T�͓iuI�F��6y��@J���.fo\���^W��X9������-���(�����9D�b��{�z�Wx�(q]��P9�U�s�p�7�|��.q!��W�|��J/�h�5s��X����'"���+ڜ�Y��t�Kxw����e=���%#|���ҭ.5ẍ�y\�ر�����hZ_����S/K��҅���l��*����Z],@W�\'�Eg�<35)�V�h尳�K�,1*�6�y�2��q�n_Un�q�B���͇ﲰ���?J���^�� �o�:5�<��]f����E�6����=�p9�3M���#^��\]V�q�V�#|s�G��T%3�Ds�ex���mA�Yq�E*u�[�@��g&���s���p6�dwJ�������2�x�O3�H���^{��ܛ%\krz#赴W{7x�Yf��� �ȉFB��s(!�>��;� &smˆMƱ0Y/>~��|>����˨8d�.O �j#��ي�Dq�!i�T��Ny�n��P������x%�wV{�V��&�]��5��&���mM���2�W�os���V_ne@e�[�k��d�G�u��ܩ��V�9���5-t����3!�"��攕:�
�*N���,"����\om��iݵ�+�8uv��Z�a*�@���תb:�a�}���:�s��Jq�[:��LÍ��(e%L܋�s�����!�9ZM��XlI��H�ԋu{ݣ�����Pw�ሱ��vPw��b�9
b�T	����p�H#��Z�8�����	l��1���z�0¼�zk\�3Qu]��d��� �
�dl�N�p%Vc*������k��y\A�ϡYJ���·�%H�:�ֱ㗑��5cl����x�(=�E�d٫'��+\.U���%���-����N6ٻ��pV �wod{�{�P.?o��:mk�خ��8-Y��X!�#�΢v{B*��-^I�wJL�K��,��Ʃ�"�:��k��7��+����i�W�����zT�;T�������\�v�w~�eK��1{�}��C�=B�X2Z>MK��G"����YgԺ�{TfR���oGr�_@������U\E���U�-̊i�i(XX
��6�����v���w�.�)3�f:vѽ��,I�#k�M@�S�JU�߰�+NǺ8+{a�.���ׯ��j탗ktE�z�JMTC�-�%��Ⱥ=�ة�@�����.B���,k$��n<��Sی����'+0�;;P�I�e�1̥5��k�=�B�=$�[9ފ]�Z⡶�rI�	���Mdk��3t�P^U���4�S��	�ݮ� ��h�{=�qB�:�XJh�,�p<\�/qu���q�<j.��WR�vÕ]�����6s�@���62-�\�n�$+�@Kd���QR���k{�I�k������gs��o[�W靄͗#`t_���=���U*(�GF�G<����
B��y�r��c������xE�!�R��c���T�Xs��f� t�v&��d�a_F�q��C��rv��u�Č�Bb�K��iF�1�	:�p�CJ���V�ܖί,����g �L�;bn���V��s�wJ��eń��b�8�0�v�t�8A�u&�n�a����;yv$\�$�%�n9���
��O����Ee�16\Ie�9]5Q����U�7TQG�{b@n���r���(�e��~�]Dzl:����Q�+y�Ɣ���u2�UL�:�X��y��D��á�u���@�A�)^߮Z�[օm��Q�j~Re�n���°�#������U�O&�v{� >�ƴ��b����q�}���v���'�z�ٚ�FR� "e��HY��q�ŏu -S�E5�X��
ޫF�Й�OFRl_o:�+��tigb�/�`�e�R(Et�D[�:����̈d�ҳO`���b��/����,�}˰�ߕ`�蝔.2f�,��<�����/�j�1"�l4�8=��#j�[����Y{�q���b��L
����z:����E�Iz"��MG�u��T�o1\�z~ȕ�2���������vF��Jvk��u�W�9{T6��ɰr.�jfͧ�]P�7�3�5��������Э�����3�S<|�C�{f���m��	m�,7�aU��E-N�b.�1��<�P�snج���*�+��h���bz�|��f��'O<��5���ꐮ\��c>h*�s��h�y,C�.J⺆U|s��]��I��y��r���!�-�
��_���G��ok���1���6"8D�= ��huK������I���$r��H�Ga�J�2��T;��m�
2>zx���V4�ӛ�zﮪ�1�W���fD��(��͙i�J��=��cv��!Ɋ�ڝ�k�Mn����蔴��tm�B�P�C��B��^l��c������>gȂ�<r�	Y��2]��d�)L��]>fNռU �ʷڻ��M"�D���ޙ�3Q談k紴m��E����&��I=�Е{&.J�d���.�z���.|���7��H<���w�l��[5�5��ϋ��vZ��K�aP�X�\�K*�]�xe��ۅp1.D]�S���`��K�:m��j@hܷw����D�R�[�X�!ϊ߹a�/��_s��S�K�du��XR���t�i�ߴs��UN���<(�� �5%q�s����ɭ^�m����Yg\V�W���J� �c��9����:x;��O�p��`L��+��%tL��\�w#�͗c�b���@�8j*��O
NHK%��`�r��5qT*Q�/�2қ��8Kh^��Ug�ɵY�B�1}��p��u:?v'L��1�.gCo���=��y*;v����F����Ԉ�xC�GC^�w끌蛗���$ ^��,�����WuQ�$��ϴ�.X����ݣ8vӰ,_���wp��U8,��+^v��mɭ\�Ma�;f9��h0�(�2��nGE#|FZ�����Bv@��1�ڨ=��K��+��=��q�����R��>yKg3������9����֊̺c��x���y��.T����WQ�a�&��2�Y0�ֆ&��>�Q�6< ����v�0՚�{Ao�1n<�E*a��k9�k�s
�3�n�|ĥ.��á���[|�1N�S#��f�q`ܳ��+E�Έ4I� nt=2��EZܹq����V��R��j&��v���Rw��H���i�
�ש�.�!��];r���0N��	���ڰu��F�Q�1��,i��j=&��A����/��5�+f�/���:�Y:���55��� +�x�iaS ��;���A�J]�X�s�Ӟ��4%L�lIa^e�SvI��[CW<���7�)3 ��%��Ul�i��Z�;5vu�XKV=:�k|1�D�X[}D$tT&�E�G\wWS౗�NT�$�e��Jዋ]�v2F�2�EL�qu8o50� �dk{t^�'j��g�β#ٽ�IF�^᷵Z�-0O0�2vƔ:�N����v^2^��ݛ��gT;tn[�����v�vr���
�4$�˴�Q����P�L�'Sk[y��R!ld�S2��}3�]��""�8&�r��f:2���vaE��7c��/N�I��V.��A�Q'���'R�sV�����r�d�{�	�d�� .8���36Ю���n�V�Ax�.¹�WP93Νi!�e�ͣ�k��]�v�U�[��\C�����\�0��tLXE�xr�������%HW �/n��)�O*s;�2���m��-�f"0��,7����:9Y��\ވ�Ŧ����70��:�oG#�ֹ7��]r���vˣ��%�Gq����ԝ3Fn��I�ٯlSWY/Jj*
sJ`�kb�7�]��͔qP jjن&ճ�&���6�컻t�	'�MZ�C�.u����\[畮4��(51�a�up��u)��4�ͣ7�|Щ[0ӭp��f�u�cPX�v�������W0�܂�Ғ�۵P�;Pp���s���FG�B�n�^��WOS��:��b�unJ@I*l�Z(��p�{O,����,���՛�#�r�=�������,Y�w&�D��͹Eb���U�XҪoa}���;�%u�;�#U��Q���%�k��p�����v�n�:.7�g'f����O W�z�))�Hˮ�z��Ӛ�����UЛȳ{D0:�0[_T��&���J/��E#y[�F��<Yd�KA��0E�c��Y%���P6[x\���ﳻg&N%�3�:��{�F�Z��W��;��b��S���b��/	j�X+5���s iYҰ��"��]^uո�t]�E%U���dq��$��z�	xh�V��cVr�����v8��`� ��k�5d���/i��B��m�yI U�C"����r�H+'U��-sz����5`Ha�:��^�*��eu#R��٫�r�B��
&�F �z^�Zsr�� �¡\��!ge얅�gY�ۙ����Y����b�갑iT͊�z��黡f$+@�)[�������N�\ͧ���<���U"��UH�P1 �iB
JT����c�ŨʋYY
��AI+PR(�`�QaZ²T�fd#l�V�@��rʘ�Uk
¤R��,�eaY����m"!EjT���P+P�jE[��`
DQX�̸ T�R��%eB����l��
�����(�T�-�-�����
��9�[eeEb��(�QD�ADA@�XAEk�bLUT�T+IX�Jʒ����hЩ*QEAb�-
Q�jEd�+P
2 �%I�0Y����"�U�+
�%J�%��b��VVڲ�J���@�
ʶʨ,��Y�*He*���P�Z��EXİm����Ad�-J�(1+�(�TȠ,U�D�E��*�
�AV)m��[jV[H�B�R�őm��(��*�PQJ�I-�H$=(����+<+N
�'�c�\/To�M�;�>���u(^P'�m���U�k�!M�7��;�6&bB�}�t�7�4�z��0�g�N8ͤM��"N�f$�����q8�����$s)�:�ӈz�!��a4�|§P��������s�g�*��Ϲ授���H��4�z8����/��t�YGϳ�>��8���I��Ȥ�
�Y.�o\`m�d��w��:�� ���Ĩu��?&�QV����h|�0++�?&�u�&$���!�b��=fm �N��}���Z~~�b��DU�f�����Ub��W��UR�=I�����O�T��s��O�VVJ�����M!Xl�kP�5d�4�3�J��Q��LI�/l��|«a�W�k���c�'���������<��y�4�mĜN&=/�j3䟜g��'r��
��i�4��V�szߴ�!�L1���&�++8�^��m��!��eVT�����.���ɟS�i�Qf��}��}�a�r���b�į6=Ç�>����>4}�	��I��Èc�w��4�RW�L�M�bAg�7�a��c�4�^�2$���ϧ7�i�P�r���i�&0=�w4γHbq�b}�����y���+��=z�aS�wT�H/P�<�ͫ=IP8�e����&"��x��|}�!��B�d��sE���K���m�=|H,�,��Y���y������]��}�����w]�����������J��<���SL=g��xj��:�C�y��H*���.��=C��1��Ɉ~�C�������ߛȤ��a~�1�I�*~��6�nr��i|>�_�:�w��f����=�
��'�u��2T�B����LfՀ���e�1񇚡�8��~O~�i�I돬;�$g����z�I����z����8����3����>��9����ck��,G�4}"$D{�c���ϒ_�1�l�Aq?2a���1ĩ���Ԙ�z�Xl>�!��O\VM�LI�+�'S&��C�+�z�_���ϙ��5�N>3L��|{�s?���w���|�ߵ��`"M>3�~�z���~採�:�<�ܕ�3�b~C�=�sĂ�|¦�y��<H.����*��J���1%}O3���iR\�7�&$�
Υ!<� ���]�+�,�NU�25�d�٬�,{Ee�1y? ��=P�	�ָBu6��꾡��+es��"��y,�	=iB�%��*�w5;�/���T�G:<�֚�٦w��n'x�)3�G*J�Ipҡ�	9��j��_G�uhg�v��P����uXo:��ꐡ�C�:~��@��� �k�:ɴ�m�����CI'��4u<a��{t��b|��c���@�~C�b��CĂ���1O��ū�
�ϟ�b$'u�~_w���^gs��{�'�I]'5`x�P��z�|��a�<哌<5�m$�ϐ����O��d�$�O���2|�Y��2C�>d��a��x�i�\���n�^N��O�}#�"$G���ğ!PԴ��O��i6n͠q+%f�����c��'��1$���=�� �N��9�v�Rb��}�2u����s��T4�d�ĞФ���uS���N��G�2� 0�ӿ��=�!P�%]�3��Ag���4��ى6eH"O�Sf��^ -L�8�Cl��&!��&3�u�'���� �����4u�x�^���#�sK�T���wp����} ���>�ʘ���=a��m&!P�%�{��m'P���y�7������Vx�fS�%J���jèi ��Ӊ��0�0ߔ4�0�0}pU�r��M�Y���_� �D3��8��
���8��qd�v�~aPY�ę��t�I�7�|�<I�+*y9܆�*N&�LaXW��z�|ՊL@�W���"�C�o3��;�����z!����`v�'P��z�|�쁤:î!���u:�$mZ��Rs�1��w4��*O����p8��b{�̆�4���=ަ��l8�&!}5�1�Ǐ�m	�G9Ϯi}�{���k��@��>N�Xo��5���,�k=d��Xu'̞��'ْ)8�}a��é��g�=��m�'����f2^Ru�4�Rb�O�s��� �H��\/UD�����Z�l�k��!�(A���&'u@�u�!��<��!����nyf�I�bA��|�j�$���&��J��"�q
��}�`8�v�dߗ�g�w8�l#��b�|�eMI5�����]W�V�|�2T�|΁�ޔ��H/ܰ�bi��+���M!�>La�<5|M�q����?'�1 ����4������
���C����I��u$}���� ���5��3|��N��Yk�2�ulOY�VfΩ6��d(��1}}�Q+߻ BjV��vj�OB�c���]��|#yP�yY6u���j��2+��RB;����gm�G�'2�s� K��:���'A#"�UgW��q�� " ��ͺ�l+
��'�����Cĕ�[�ed�{�aP�Y>f+
�I�/�'�\v��|î'����m ��������1���1Y?%I�}|���Zwp������@>�!#0}@�V�L�?=I�Xbzk�*AV~Itw�l�!�Az���uM��J�Ԩ�|�m��SI8�O�=q�Y��B�3g�:�}`T8�_���qx$Krn=��YޯDH���f(}�d}�K�O�3I��V!�����Az��{����8�3�13�{�f3�b?���$Cӝ�P�iP�����1P�%�R��J������M��ً�)���H��D�:~����R|��.��%�����Ӭ���]!�a4�2T�|�~�x�:�Tw4���c�W{@�������O�Ă͡�~�S���'�-�}k��j�idߣ�9��\=b>#� ��Ά���%Ag�0P>J�i����&$���0ҽ@�߹��V�}凇>��<IP>r��%E��������b��y��O� ����=���v��͡���[���/������s��I��bAOo�+���a�Ն+'�R~vj�$P:�!��Ĭߔ�3$Ǩ}���g�~��hbA}���u��������t�$ ug�x
���|}��Y�:��|�O�<5�mX
OP�;�ISO�C��&�ɯ��Leg/)8�1�AV'�T?=f��<�C���1�a���i�}�=������Y�;�_�עDBC�AT�30��=Cy��~C�1Y���6�Ԩ|������i8�C�9�j�R~�ed�~@��H~IYX~z�<7@�q��M��xD}��S3���ܽś���b>I��0���C�bw�d�>O:�u���b3=�U'YP����C��5�Af���w'�J����L~dĝO%�2�U~@���DP���~L]/zN�=��y����ɤ=IRw)�4�d����<�I����|��I1�e�2��3�S��|�&$�y�Rq�O�C�@���V��H/̝�   ���m[f�{�I�J*7�sp"�TQ.v�M��k�����l��"pK!��8��w��k#�ڱ�P�:kT�V8�c����r^MFa���;7Z��0�C�)���C��9�3�b��Ԥw�����rg]��XJ�Y���]#ɑגy������~{"�Y�I1�:�CIY���k��C7�ǉ�L���1��'H�u�����&�u
�a�����U���;�~d�c�NNө4�ɜ��{�d4�d��q�����o����k������g����;*AVE����A'��\C�ug��Պi ��q7�6�CĂ�o0?0��=C��&<C���<�04�Ĩu��{�x�dĜB�����7��{�3�_�='�W=�"$|��,Gބ���VV>��z�Y��7�kA�b��J�V'����Vi�
����YS=�0>f���C~aU'YP�=O�ن���;����h�FG���YX6��'k� ��DX���jq׬�����1�aU�ɹˤ�!R�W����ɤ�IP�:�q��ʅb��_�O��˥`)8��M�Sԛ�B����I�4ď�I�C%z�ק��6�n��{�1`�OwC;�h����Vns�4�_Xl��:�3���{�d���Ę�|�m�g��r�ĝ�z�ɜ���] u*,����J��V��b����������=��p�� ��~���8�T�����:��2f���3�d���9�����d�~�W�ă���|@_�|�3ӝ��x�$m�w�LC�1d�aU
��B#D��;<��=v�g�ϓ�=���i�+;�a4�Ĩ|�e��;��"��>jp0'����G:ێ�I���Ք��gH�t���N�|��H֋uJ�pp�
�a��@W�X8
��oiyfP7};��0���f]�hN^Be�gr_e����Ex�8<��鿠_KUΧ�C>�һg��8S�cxH����#jvs�T�%��Z�q�[�;-���'�gZ2��҉{��� �*?j��Sx����]KM�-�an
]{�����|y޲ْZn
��qua�j�!�N��=� q���u֍5��(�dh0XSP�Ѵ����-B��9�Ws��p%��yڽm!�N�r�us���]����)˵�y´�.�����SE`��>���gO&�N'wT#��=%Q|S��Y�\D��s�4>�<w�@�1���ʈx�@<:)nH��˹��l>�1���_��L؞up�VNS)dlr7�e���G�d�O��TE>�.�*�YGf�s@��%`*j���kG�>�S�N��q��F>��q�ziRw��&�of܈CX��m[���V��vb7�
wQ@q43'�]�]|�ب��y�Oi՜��=�y@����<ш����C+߬�FA:!+��"�y��~<����Լ����я=�A��N,���j�Qp��_�]H�	˚�_@!���Ȯ�m< $s9t���H�#n�"��0�r�\v��Bf���y:�w�2�a�J#�|x}Z��Q���$�jQ�)���a��W�'��H�<�j#�=�&�ȸ��]�s����k	?c��z�"�l�tB���nq�~�WjR�pg͕&�<�$Ê���o���/�\�˴��]�#X1�n�mTυ��Lv��9U�Ň!LWɪ����}�*L9���8�3��h%�M���8vXAS�o,@��֮���+���H�o[	��i�2_ս����p��R����������P�\1����i3n����k]2nb�]�٭!pmtc����Q�;k5D}�J��5kMp]�x;���d@��<���B�
���ӵ�w��p㦧��9��X/���Cn;�K�t��*B������%%�rR�]fU�_�Z����"Zta��GI->^^�U�U�m��E���_T)��"��lF�:'����V�V�7k��h]��r�y>�Η�@�o�P���π�`�7<�������t�צ���X�ãX{]��2�N��{�|�Phr8N��Dk�^���61�eq�Cx�ϮO8�kmL^C�V3x��p|�@m-�*���%}�o#�ֻ�A7��?4Z6���P�3Sxj�S�
l��������柝]�]�S��;œq�U.�0��ƒ��ٔ�4n�HRz{a����q�<6���0�#Q�3��5��2�q60�+NǺ(�+	a3ې�0�zS����O}�kֆ�1����7�a�<]�Hc%���H�8ұ�z��m�W�ɕ����;�+�}��R��NLF�ȫv�E�U�[70PP~�-�+n��L�J͛痡��kx"=�����#Z��+UFEl{g�7��S�27-��*,��K�cR�,V���aq慛�z��M2�9[6T��՗��L�k��ި�=��޸�`�+����m�Uł�����U�\���̫[����0�w:�y��X���Dd���e��*ޙ�l�-P�Qt|���Deto��Ly�Ou�˹kH���8�/��&Et��Y8���N�qr��@���l	rlP�xng�^�
xHa�q<M�)�����$O�uD��R��q�5A��Rul�4уt75d�9%U�v�Xz�l��pB5=A8��Be������en�W��ɯaP<�l���(�60�Zz��6WG~���sC�dF����d)۰�0@�1�G[V6烪M�q���}�G�I��q:�0X���߻^�8�9��7;AU{�J�����\6�F�LV����p���z�s��e,�<�_�a�0	��6��<J�F����	�NY1�.zV5h�xvI�].g�ދK�x.Zb��~C<���6}�+Omb<��4�+���X �`jՒ��:a����#�f���!�� b��,vj� 
x�������r���ek�AOt7�{���y��H���n����g�������ps5��zc*�`m����=D2�1�^[NX��+��f���HbSR�:ȪS~�-����;���7���Cw,:*�<l�⮕����qe��7�����ň�P��������h��r��������V&	�a��y\0K�bK��;p��{���i��a���?x$�(ܦ���������m� �?��ܢQY�]ws�x|-+#����ׯ�=�v��i��.{<��wN:,*����DV:�@-eX�>g�:ԭÓ�3��ϣ�Q6�=�ߔ���'��.�1��/}6���Ed!�GMJ���R�ҫ�Uށ�9R(@��!i1��z*���D`c��2�
}A駐�Xhػ���l��r��l�ǬH�)��� �g��R]���_����5�ok��c�ro`�!�lՇ��_�V�Up��Gh�_�H���3� ~��,u���0K!zv�l�y�or�x�7�88q
�
���E�0�oĮ:HN�K�h�3'�d|��a����uJ���
�iu[8[�#l�`�O�QH�F��7-h��������Z;�ħu��BO@��vw+�/Z��Ɋ���l�d',���e��y)��ב�Bcb��u�K L]��;��5���5�*����r!�	�;��<��T��5ݼD�U�L�rQ�]��Z�OT�fa���ԭ�]�[v ŗ��2�v17{��(漞�G�]����\��Wy�͹zoo$w��2�.q��u��Iml[ԵdJ�	��p��
C׌��me�q����W�#��ܲl�K�eZQ���\�)�}D-��r�\�Y��v�:�kÅ�=�Xb���)���<��3�r��i�<gimܳ�����M�y�2��Zأ=y?`�kqmu�YzP��p� C��@T���y�����.Cv9��5��07�#m�_��}e؟m��g���u�@�Z�s�!���.3�[y܌�+|�MQ��%<61�3ݾu�$�_C��>�V�ㄨ�3�ί�����5��׳\����ݎ�p�E�.��	;|pk��n>�LmOg[�^�DS��X\��ԥ�Ggy}@�����]� �ÿ�j��3HLק]\,�(�7�Բ�����w���!
�4��3Sp�NH�3�O�:����Bə�_'�q��d#�[/Ou����t+T��UOO>K���Yp�m{��5�rb7��ѢB�&��̭ĖL
�;ͫ�q�gg-bj��"�ܝ�ӄ�[���^����yq��%u]DW�:XpGC��c;�g��܎�V�v���v���Z�B�쑂��ȨN��,3"9�A��� 5 ۦ�7�Þu�(Gwǧ7���/9�`i��f�'C�ܡN���]�r�U+}�i}S3]Iq��}v3+`�	�	sa;��\��K��Ք����~���7ۑ'V�؍5Il��*Α&���%v����܃�<T4Ƶ��T�������K���5:����~C�M��ș���A�N��*B)�$���á����eL��ղ�|sFG��Oã�����$�}P�S�E��U�\'�$�0��o�(��wa���1�x��X�SG��\n2��kr�����3��J�@ul(�
��t�,͙�A�5ዑ>�\��F�cM׶[�����`"c�P|��c�9
c���X�Us���7V1���p�+�c��"�p�n$����Evk���Y倧Q� 1���u���,��r/W�T86�t�����0c���k���L�;s�W�y8!}�8��f'-�EJ�jr���*q"�2ɴ�8���C7�b�܈���5tO	�>V�^���!���uU�v�|3P�*�7�f�K���l�-�n��®����F��FY�{����h����Nq3���.k
�2g\��u��߷S��'�zEB�����}ɁgL?@#��C��?3,Ç�*��j��o�Uxp��yk��u�P�V#%��Ծ9����Y3Pgo��D�L��b�xx=�Z[����r�����i�Nm�K�g ��X���i�
��7A@G�7������v��Ǜ+um*�-�%��[�Q�n���u�irU��9���Z��h_vj�wru����(d��	�*f" f�\��I���
R5�s��[���*tYyJrʍt������[m`��9�h��}۾B�}�*,ymǒ�f۝Vf6>r�L��<���tu���4̺G��^��:��G�Mj���ږ�_6n1{I�u�K%�7[�}��i�ڷ�0;�_@��B������ZO�wn���.`H��fqҞP`�2T�ɼ�[���Om�qZ�-��I�Ε؉ڮ�j�wf6�h	A���3��M��WN��R�g PVo+A����
a!����g���c�}�>�[Q-W5�=���J��{�77e�K���.�ܛ�Pgcޒ+�d��\m�>9�
|z���׸u�b����:�e��`�wƬ�n_�F5J��
��{��d0����q�y��b�W���,֧I{+5��EkI���W��7��^n�œTt/��	��� ,7]��*�u��hY��Q��&�K��Cَ��Y'��ޚ3F�[U���o{��m4��qw��u�����I�js*�mW%A�T7nj�LVS���/z&%�{ǭnӷ7+E��P���u�n�n��%�⠔�|���O_v7T�a���"�# a��͊��ְf������f���%�p_3��4�(#�sV�ߐ8�kY���VK�)�U�jU�G"*��1L���I��V)	�mEi-#{Ob��+�6���٪L^���
�hf��)�r�����e�{�^ճm߈7�݅����:�LP�F�t�:s�Z0���8o'�H@�j"b>7�'�)ڹ]��&�ά�u���9�RԎl����0��s�2�1RԽ��W|�D;uL
����\8d����+)�z��y2��ܦҰz�+���b�P� �n��ne�d�LH�lͭ|�]>��t���+) �m��։6^+s��K��e��^�t��|��y�q�˴!��Kq�Z')f���]}�d�~
'�X\O�P�-�N��Q����Np�h����*��̦���\[x���\���X��R^n&�8s�[}Ę2.ىa��勑��}�u�z��`�]><Df�a ��;���[|�uCY׎	:k�]*��Л�q�{)n��vb
��Eɵ6)���f��gV�.Xc�mn�񣪲��-��e�ּNv�QYAn��ThD��r�0�}���}�P,V�b�4�f�a��1I;�]+
��%��� Q����Ά�n(���d��u�)e<��{��oz.�m��흌��\��B�6��k�t/;5v��)����F�(�Yj����;�Ν3����k����/����(��Ɉ�*&5r�d�A�ejE��c+(�("E���`���Q�P+R*9��6EҐU ��J���U"�H�jT��YF(�-aX��(,b��
�-�Җʨ�,�
��[ER#��[l,X���Z�jX�����Qch�(��UEF1*b0�Ԋ(Q,L�X���X��iQШ,PX�V���A
�Qb��-�PDR(ڥ�Q�+��U��
Q��e[DDE����-�d�����b��QEm+Z"1DX5�T"�b1@U�TUXԤcD������U�1m�PEbƉcIY,R����VA,�a���J�Ю\rDEEb�D���+(�D[Z��X�m�K
�(���U�U~������}}�ڏ壣����h@��KR��u���x����V�"7��GG��Qa��4�F��'B�"�od����~����U|ߑ~I�����̤}̏��R���骤��M�H�˨L)h�F�vZ5ϫi�uQ�prܻ������2��$��P립,L��5O��@�|J�bsLua�F�yi�'q�n�p����Tke�!oD������_7uM�PF D���!���~Q��vw���&3�{J�P�j/�|�t�A�08nlgκ�T7U�-�֕.�^j������X
��DĞ�dX���ݎ�L�������	��h���)�ԍt��Lv���6��.2R���I^�!*a	��a��U�3�����_�J�y�.�X���Ѥ�������b������u'ii��^&��t�]�a�3���+n��;��^��bZ��R�GL��s�Gt���H�3PG�ٞ�a��vʫy��<�+ȥedPX҅m4�*�g<6�&��w
^�	 a1'�Q(nY��nL+z@�
���)a�lS��a���
7�����-�y:��9 dۻ9R����ր��`��)5���Y�J�Rsݰf�=دu��{4u�ؠxtt�1 �V��0>�t��2��YdQ��1�]����wxU�2�i+ޣb-�0��E�w��]sݥ謳9fU'O�Y����HԎ�w0{�6��+"�wk�K�5a���U��UU�9�m^��)���U��c׆���c:@�}N�n�%C�FFvש<��2@2��Ί���*�%r8��Ƌ��o��o��Cu|�yK��l�:W�U��tn��7�����ܑ��r���$a)X9}�Ӗ`��]@�]aC	�67e 5g���b� �8kǞ�v�qn���IЕ�q�.{�z�T�xө�w�AX�J�ōg�&��k$?vkZSu-v�@h
y���w�+}����kul�cyV_��<7�6D��I�ܢQ�Y�]25x�[)���z�1vq�����-X���";ӎz_\֘��\�Z��3ɿyC]\���q����hF��ax��LP<i'�tٍ�a��Nm�9E��ooUsAS�R�g���G����P��Lu)�ؚ��dhZ���# ��v�<�O`�{���!<"���'��-��"���'��8
����i°�_���G�k�p��"Y�����=������ՓPr���q���'�v%q|eC��*/�&�n2���TZ�c0.���="Ă%�c骉���*�=z<k�C3Q�u��d���f�Ӎu:&XV�ͯ:��G����Wf�*Gԅ@i�oZ<@�H)4��&�n�\�m�Y��u!z('=�CsC�@�
�x{���jR�S���ޮ=)�g������B/*�R��Ӓ� ;�
�E.�S�9ʌ<��}�ue�FTP�	�1͊b�>�g �@F�(ڞ"�:�@��ox�Cg���cS���p�M��1��B�	�Rmm��e�-��`���U\Լ�� N�Ok��1j�VE�ë�d<q�P�:�+�W8��Q�g}�ԙ��/ֈ�E=b�M���h@�,�S(�೮��=����t�p�2=����O�]�Ea�_/�+ݞ����Z+����a����GR�^A=U"�z_��*u�r�٘�����c�R:���ΐR�4`����X�WI�B��U�/��sB���$D~���.��Q}o��"�|`S��񖕯Ňy"@Sۑ����o k���u��_?1�i8 FeF����!�v;�X��HN����z����4tq󅗎��p�+�GOf�#;d���=��aN-E;ڭl����f��U�Ƽ;L�<�����a���z3��lW�2�=]pz���mtua�S����k/A�[�v ����B�[�[EǞ܄R���m_7c5jDDsf�m@�Sk5��j\�QNՐM$��`��Kt��^�A�awg�����H^����t�.R��[z�;7�3���(����3{�^��N6AF�l�(� G���䯲x!��C�N���q��;�]{��%.����[sݰ;~��k����V�FY�,�2���ф��,��dR��x&��ɑ���M������/��� �ݼ�0�9��FJgd�y�Þ��i�Uځnx�[U��r�m������:H�r��<�c"���b(6ͅb22 Hச]�2~s����Mɾ��%�Y-��f�ᴨS��r�`N�"<ʘ�"�-F%�E,.���Υ�^q{����>8zͰS;� Vu&+�\��f�h��@k�Ar��>�5�҅�{��K���p2ܘp;�ا��*6�UA��R5����=�{-;ͨ�y�)�AOM�&��T��$���5Au�
�X�:�c~҃��VK+!���y��{A>c�tÌIX&-���|��!{@[d��x���ٮ���_�倭��P�N^��T�<��������s%l�DF �
����rt݉��lN�X
�ߛb�����ۿ���,��>�ܖ㣶8�� �ӊ:mН�p�R��Q�Z���>|�˺-�Y}�/���s\�mhg}k/���A�*Q���5��qM�J��Z^��G�:�I<�_!�" =#����͚ͬ����FM&�������}��l~�������ܐN��͉�h���f���"ԗ\8�NTY�/x�U��Κ�&d�X+Y�ӵ�.���1N5\c�V�xR��eqb39�%�E���ߺ)�늸s�4cPt4Gq�;'��$M*rP���氼'\�uT",�e���r�V��c.��l����N�<���?��u��>n�K���o�QCY8��T�Gf$r�d�~��*��I�c	�jqV�c}���8yI3���}``#�DǦ��E���::�.�-�
k.�H�ˠ���U:z�c����xj!R�daLm�
�@�|�%*�nin��3sw9�m�����;�uy·�]ؗ��Ќ�z:�3Ǯ���:x�/GV�}���an{ջܪ/�V�v~\��F���PR��r`r61���J�ZuQ!:��9��koZy����0PUs�3�v���.f���&h�d�	�Ȫя{X��{��y�Ö %�DV��o�J��TzKD8��=�X�e$�Gd�V�\IN�d�<�^�rj��U��Q�����5����@I)�twvUX5��7��Q!�+�K��9�ץ�L�Zj߼"��=��Ք={į>c��q�{�H��3��C7�7�Qr)�E�E�h��E�c̞���(�f!G9��V@����b�EДg������׽�Y�����_�j����JNr~GI�{��+�e�0R��\n�ҍ�V�p70WIt2�oQ|�(E�n�M�!��"�t�������&�.���}V�dѓFj����܉J���ܔ#���`mY�.�TBj�|�U80@�0zf�3{�.H7��L��l�'iq�#`�6-�q�gY�q�J�.3g�0���P��S~c�|�<�ԍp�k��V��x{R���T��O!��E��F�ޟ�RL�a6�!gZ�c�gO&,88a�b�#&�u�&�T5�wخ��U��=m�����H�u��Ug��zvp��鉨ͣ�*0ԟ}q0�ٜ(dd�1XP��9 b�M��Q9�y#IeЀ-���v6�y}��ܢ2�zH�S!3@g����)yj�~
ʗ������LV�jv���!�N:q��o�%���1=&r�>{m��'6���l\f�v/�k ��-mPL�}^~���=�Ds�q�����B�9 �#�����Œ4o{r�	-:�~2ǻ<'�/=�V��x*fU�� >�7��3v�^��-�i���7]-,��,Zw�fޤNR��;1�i�칆�/���XҦ���#�Ɂ��7JB1慏k3)+��K�,9���K��Qr����^�{�d�bg����1~�pO]p����N	>��e�g�q�pT	��!��`ւ(C�9�I�⍰@�\��{>X0˂�R�>��Gdt<�]>Q�)�c�1"/ ޣ����w��t?Ӑ�t���AH��$zN���*��͖Cο�Q�8)��[u��o<WYo!��XT>]֋�霍x&�J�:� �vĉ�]"D��xbun��J��HPR�QϗH�Ҷ�j�|�{��c˂�f8E|J�2�V��ճ���r�6|��
˰�Ln�\�C&'EB{V�AN����G 
�<�!2D�o*�26�m����]�Ip���~]FU�h/K�~JF�Rf�F�} >.]W��4	5���Ti��%�_A���p��g�h�u��m�35��L��P�-{���DK�(�#y��̍�7�M��� �c�lكE�����x{]�qXb�_/58�o!����%�e-}cH��s� 1�Or�*�{s�s��xkE�V냇�xAaY� W�[���܋�]�n����Sz=hm�B�� ���C�͑�k`�-�(��T֓]�̩�(},�Pj�t��j{gd��Σ���:�72�ƱQ�E��ٽ�`�ua��mC�am�R�S�|��D��Z�t�F�c�)��`�Ӕc75��KWK���܆������?x�{7OO-s/!��D|�k�;�=uj������^��W�����}���n�7ԩ ���J����ޡ �w,���J�iB��E¾�|4g՞��u Z.R\,�QL���OsY*ƿw]�����ܡɅ$^�'o�r-�%�7��TlP{�x��<��x۪+ar�y_ ���rg�ȋ�a߲e��u	f��C���c��e#�[��JI���f\�if*vѺ1A�I��K��
�Ip
���2֎�ۘw���h�]��Bs��Q�U��J�x4�}��My??�b��G�@�ߛ@��3̭��D-�������Wu��J���I߭����0ϛ�a��7��y# ������<�a�]��ܰ͂	ɛ�A�׽`�e������{Hod�ҙ�t��`!��1]�������S�I;���Ϝw�zѱZ�&a��a҈��bј�RC�v)�[��cW�]�0�.x�x�=;�3�S;�D+:q^�����%8��'>��[i*�ŀ���)풏�e9aZ��Нٝs�f(�u�Iy��*�f�7��ڔ!�?+׹�"�h0��y�o�w )�`+g,j��]]Vڮx��z��r�zR��E���&t�G��ю�K��{�x
ތ�N;qK�;�ݑ���ӆ�@�raP#��ok=�Te�TV�$P�S���bq.��W�&������K���I���ZrH��2+�#W�vjv�>�^����.�]��,Մ�8s#��$hk+��
�X���ȁ�@�ϼ�$+��+�&�Yֶ6���-�^�� Tk��3�I���5�y�%z[���%%�r,u�z0pX�SZ�B���c7<��##!3�����!$��J��Y�S6:_C�
��g�����yP�;�O&obh���̝��d�s��������v��C�g��(����QL�h����g|�8��X=|��3��q;=>�:�_�UB"5ϯ@Iۃa�&W��ڒq��Yk&��7`-nu�o���E��/�����U����k�����m�0��A� Dx����P�z��.4���pѩ�,������U &�x�Vc�>��ݰ�UsN�p�{�S�3�\d_�ؕ�_�r�lW}
�D�Fׂ�U4 k>B*�lխLnz��ͽ�((en�'M��i�ǩc���B8�fKb�
�l1n�R]wRoPїYVu���_Qae��x�/fdj�秹��Ð)�U�{��d��%o>�wkk���/T��*J�͈�r�+���-H�Y0�g��H���~���ꪯ����m`uY?��/r%q�
�{P�Q�։zu��������YB�wt���_^ʼ��9?H�(+�Ŵ�>E�q�����q�q�ݫ��u�k���ܧ�;x�+;1K;-�ݛ�W�D���|E�Q�n��ˍnE�e����9-u[{˧y#Hv>���x�w� ���@�q��R��ZM�)2!��4q
2�N�v��L�|�m�S{X뎼9]�7�J ruBP���$�GMO��r��D�R�wDU�ދ��vN�n���fnh}�W*�QR��#�lL��ٮ�_���ֵ�T�ۆ�y���E�[�]kW!�Gu��*2�#"�� �>�;v�E]�u�����<�A��r�t���gLV̐�'��#`�6̷�Qf,�{"CUAtl͙<I�VT�oT�g�dĎ�L��$G�e���;9;eG�3�q ��v%5��['�����y���s��jz�ܷw�Q�}r���5V�
�W��+e���o\�����S���G��wu�<��,���t�Ә�K��1�MՄթ��8�ᕅ����;:Y���;��9��+
&16P4,=�ͷsN�Zt����O
�+a�)b��<%d�ů;�v&�p����n�dN����2%��F�]�B�7Z���u�7M�A.;�w9S��PG�c��,d�8y'Rα��ԡ�L��Y���P)Z>%:����̔Q�TN����'�σ�G���a�p�F��b��A]���[HmiA����rE���T�YX���`�repP����3�gQ6�A�̘�:���(n�&�Mt������z���k� �	�k��ͣ ��*��pKB�M��vt�r
{�5@��'J(`�����^1)*�pU�W���O#-d�kF���Ps��]�A��B�*l�D圴$�{��Z�Vn�u����,地�ڤs�Mf����S��>�a*6�e��2NGEV�+P�b�LzR/@[�]Vﯜ�ЕM^��������k��9N�c�Fb�ņլ\�D�פ�.Ӗ�5J�Ձ�,�M1Pj�W��3r�|1�`��J;[U�*���FY	�j��}�jGKo4Bnd�Iu6\��e;͏x�8i�&,j�i�[���}*�&���C7GM��V>�p6��n�'h�1���+�����ڳ]c�E�*��ǐQ�����7��d�Q��yJ�u|g	�tܫ��s5�o"�A��B�@ꪑ��M�5���]o�qy�2֩|��L[�j1o���x٬
�!O �%�Mx� �tz�t�p[�����C�N�uڠ�4�Z�	����`ʀ�z� T�,ƀ�U����2A��)>{!ݰMe�J�^c9�sgH�ͩ�+8,��⸣y{"��B�TfC�f�����u�ж�tU�jؽ��Z���v\���602���(P�wo����{6��B��M�w���A�&���lD`x�V�B�jIf��-�%�PV{��;�d�j����pe\K���e�~��,�:U�;A�Zt��ΰu*��� ;۴Q����s��˰�X�����\7�(ݷI���p
Kn 4�Qo�D�%�\���73f>J��}r��uEp�-|I���n�=��f��݁j�h�q���c8�rfK"d ����="Ӄ^f����6���oFS���ّրe$C�&+|�*g	&rx��Ty����p����a��z2�t�K�7ڑn�d#lCQ�9z3V.�J]n:x,��ƻ܋�1l
=��,h�6,㫂�Y���
Z+��۾M��Pc���wWX�b����g
��4W3`e|Y��nYع	�(݀1�ʰK�vi@��^]u�5�6>���v�^��CN�iϼ�˭y���ͮ�~�Z�T�Q���T-��"+�
"�c�X,���l
�* 1QT�l��PQQ*��֑b�V�XUP�*ZR*�YZ���J���TD�VJԋ[HR�P��X*F$J�,�QR�aQT�����*[d���"+YV5�Y[l��jʕb̶&5%��*-�Q�EJ��U-��R),Uh)3(b�)�UEJQE���E ��X,D�liTm�����e�
�X��B����-j�+[E���!+YkeV�QcB�1�k`�F(֖��hXѪ���Qq�"���Lj�����h� �#7�ܸ��h`���:�*ڑ����9�zcΠ���h�_sh��E��^�r�:'<�K�:��]0��^o)�7����<=��Vu��k���l}]5�}��Q_i�ڂ�!����*��;<%U�^�� /�4xCv �H3.e�`J��X��1 TZ��\+�a�����nQ��0*��L���g��*��V%
��2����:#oݪ���(���)��� �Etvh��aBR�)��*�-Ho��Cl��Rڠ�^����o9zq��GIpカۖ�n]72ᵹ�ᥧIA齒�؞�(S!*a��<�F$)=�MM�+�0�b�Gy{C^�"�G�E!=�x���Ψ2�!����Т���P��OF�ОO"����A�ڣ�ƲTcǴ�8H�h���Ӓ���|�OQ�O3�p!�ߖﯥ���Vfݦ�z@}�܉_d�����5�ixj �r���.8A�x�������ڷHRb�9������#_۳L<�JJ��W�V
N���wZ���²��yU��o.6�+m��M�CbC�.��zC����A����؄���-�� uBxl�X�Dlc|���B�ӻ)ȥL�+y��~�#�yQ״�IdV�T�&�ԯ*�4e�2�V���;���f!պ�m\N�tJ�{{4�fs����4,�+�*)t7f�A}��W5�=�g$�g|$E���)�9�b�,�O=nC�,�Y�#C&i���^�M��Zr~���yX�pZAӼ"����y&7E��5��to�JF�T�`VN�E�ڀ������-�^�n5��NJ��!�y:N�,F���fk%F����y����D`�;=��G5�~�}��2{���=ѓ^U|��^(G=fq�����kt�tX�ؼ
j�y�:y����m�J�oi��T:�{��js׆)��Ont��8��Eh����>��P��ԸƎ�ٜ��On�2d���PX��oi�`�^۟ ����M��G������� �>��ϴ�ɃΓ�>sY�=wo�n_���_Q�Θ�u}���>��g��n磘s�B/t�������`��,e�W��h���TFXI��\�K�(9��w�`\#u{�w�o����A~�P*'F���}3ҺU�Ƽ%v*L��X��Y_')����՛���j�2�6'ui�~Sײ��+.� ��{"eGy�߲x!��C����p%�+ ��a�g%^���u8�(K��.���|Tӯh��@�;��2b�0��=��lTр�1���v�Y��X2�
ܲD��!��c���Q��<'�[v���d�s:�@�cN�qf��9��;�r�+�A�i.�$��{��j̶ͽ�l��GH��{R�4��j�	7�*B^M�1_����B6o�|�� bJ���L<�"=z��o�y�Gd���,���tw���xzBГk3��B�OR0��VP��7o��#�����,tLP���{H�zH��ҙ�9�Y �ck2���Մ�3jȽxE�騍�vwĤws�לP�b��͎u��V�[ڙ���K�JL�VCg&:nK�q�(x�£��*wa!3�@Vw䘯��/�3h�%§��&�*�{�zv��\Վ��U��9P]^�r�G�#�Q���K�x5u�;lR�:�����V�8�-q���o--��y���k��+N#Z1��[��/E��7�z��`�5��4�r-��%�����#|�W�º0b��"{�I\t���sR�s��-�bJ	��}��j`��K�v�=҃��,��7QBG;3�k����.�*o4t�8���gx�{�#�C����Rۭ�|]�kP�r:�����9�S63������t��ћ��H���&H`���brz2�V�VKW; [:K���l��h�盿t_�sj������^s�/x'i�^���K!x"���k3␓~O*��Th�4t�y�e\܊�T�#5Ȱ�E���fd���9�ט��n�:��u�a3����KGR��2e릁��K������v�� � H�6��g5G��=��7=o����_6+��D]���:<�'g�^6|�8�c�:�쿗s�h���&o���"r��e�
V⭒�qc�|h�z�ܣ��\V�k��.*���W�WT�=���PFhE-].i)T&8i�|�j�:�_"k�e���>�ty���T�'�;� {�,��S:N��|����j��M*���q����w�v#��5F-0��ww=2�]:gxuPĲ#�8�T��j'G���}��B��7p>�ԇ�
�����c��N\���õV��2�QEJ�=.W�����*�Ӕ��4j�
�g��T���G-���m�9��ڂ6�ɿH*�1 �|E�Q�n�m&^�B������td]k=S�ߓX.4B���ۗ!dʢ�6����Qu��0Ō.{_Cr�eI��>#&_P���͙ѬK����9N�m�:}	݉�#.LE"��Q����4�k�!"o����U��X���r�N8�q
b�`I�2H}0ED'�h��f�	/�l��NnH��"�Q��ˢ1�W�R��B В^PL�&t�}��%�yˋt��n̛)�d�YW�}�B���8�ȴ��H:Pݘ�;x���2�b�[c��Н\�ڎ���syyk��T��g��\(� >��Vf���a-�;�uaꏅJȷOb�;�3[�k�����<#�os�t�B�>��zM{vxC���cBVi��2!���V[�ؑc� ~hI�'�a�:���!�j'X3p����6^�������7Wå����Ǵ]}U �z*��ϔ]q��'x~�/�2��D1U��ڵ�x~ԥ[�T��^u��'�x��%���4�f��`��Xt�w�����s��Vmp�V��E���~[W�Ds���	��h3�n��>��q�|W�b��p"D���j�L	fW�6	�EUf��P�=�.��>�����/r������yR�,�)�.צBdlD󂶠���[ϦV�Ӑ��9��2�����F��ZP��N��7_Xϛ�\;H=;3]�T(B�Jo�'���͓>�GDF��m�L��y��7���,p��wZ��=;\1��!��M|1���@.e`�����V1�h$��P�2�Ô���&�h.xw`0���0)�,� �\�j�B�<�Pqp����u�F���[~W�Q�>X�y��޹a�@JZ���G�n;����jdՙ���haB��EKk��:q�V�n�6�n�Dg��39\
HQ���Ye.�EC������]��h;�+ޖ�$6L�����˭�oӱ�������cw�w��!��ݎ�C	�ʪ���淅��Θo���AW3�K��p�-��%DH���`�g��*C�	ֵy���e�Ӕ�pMgu�0ym)�z�����Uǂ�dw�i��SĊ�n��r(���1�E�l�4��\��\q�r���*��xP=iހ��{��Eˑ�,���Ŝs���&��B��/�LM%[F�L1�|j��䙾��7��
 ���U�f�T`�X�2/7FҧƲd@f8f�W$-���44�.���lW)�CS�f�U�"\�_#l�5}N�����v�ѠI��ZN��\+�1�]Ks�o�?�p{�T;�I���C��i���,*��ɨM���6أ�ڪ�(�!Y��i��\=(����Ea�w������i�,B	�ky�X�bY{��ζ�
��W�q^�5l��|/�"�"����v�T+���lg=N�\�� Bq��*:���Wol�k�7�>!���'tؒ���S1��F��n���ӭB��>�P����E�'e�js!0VC���Y�Y������[����8��&�崜���"W �<�|�=�}����n�DYedXø��Ӎ�{z�ֶ��\���wn�8�t;j�l�tMj��u��/OniN���:�y�3��U��:����:̮���8-��jmj��z�i�p~=�W��S}l���ߦ\aSb��C߫�F2l��	�VF�;|sHp����P��}5��lZJv�P�7�8��Jo�S=+�Z\k�Wb��Շ��\�����g9�֞�\w�N����J����Q�=zgw,WN�B��k��F�A�x9�y<�>�ݞo$R�hLu���!�b��aƪ$ʆ{Tl�];���V�hsiX�n��1�o@��*�%"4$(�L��E߱�T��ʛ�U�����Ss*�ɚ��sz�����2��]wS�2nr��mt<�BS]#��zf_���S�u;g4u���7�a������ގ��H)"��C�]��+��[���+9�4���oFe�8���p�G3��zR2}��!���b|Vm�k�����d.�d���T0�M��QT��)��#f'Û=�_lJ���zq�=�٫��a��^6�����ݕ�ò�=�<��^�U	ҤX:�ih��7���=א�pS|޾w�qL�`�w�>ݶ-�҈}-��O��ޅ�y�9��:n<�k/v����Fq��]��r��i������_W�Wݱ����NvA����a�2��W.�k��PV���l�Y�����X��6S���נ�b�����B�φ�wSQ�To���̊箐{�s"��#=Ax��
ū���_V�\;b��9G�x��셱c��*k�o\������^�?���{�K�����Y��"�Q���4x�Թ��g����Ҿ�k'�㋶�^�	G+:�:�=���\$�p���1���H|���r�rm6�:��q���y��4���_���;��m�r�w�/;}Jk�l6P�z|�%z���0l�~��\/C[��yp-�io,=����	U��u��)��!��ӧk�J��p�Q^�e�lt�O��KJÇ�P�d��b��`�F�U����i���gѡ"͈K��k�_��:B��/��\��+|mm��zR��OO�^e�;�,fU���쾦�/+%s���n�ơ&;��a�b��8%.B��"/��l� ��u��Gnj��Y(�nv�x��WH��m���5Rv�Y֦�7%�#0�vuk�ً�(]�@S{D�R��(�m��(-�5�~�����WVz�-m_�uiH�\ %��鐟]��w���gw@�m���K+�630����p��	K�2�H�%�^#�p�Z����R�!�e�s��j��s�]/��f�v:�vD�q��-�lEWqKFlLΝ�AwM-���w1ʂ���q�CA�����_g3��Y�Z��Z�Xn�d��dv��ukL�<s^\������A���v��Jw+&ᚚ�i���-�m:����Uy����հgu:�v��q�q�7����`M�Ͱ�������˽�Zʈ8��|�ū�1�_V���f�P��[�WJ�:������-����趂�qM>��-��z��4!���r��ý�,#���N�E��O>Λn6WFe���*�.���v�P�ޱw��|�"��:9�i��]akqO�U��n-xz�wЪ�E��Y�䘂�q/NÖ���=X��Gnok��7V<WӐcfӻ�еѢ�Yʇ�9gT�-ڝ:��Pu�����Xl�RUŋ^�to��aWԏq��4�Nvb!��t�ǔɣ1W��'�m2�n��0�p�3y�Nz_�o��t���V�&w�磌��]���g�_�5�Y~�!�h)��}̩��7�N�!߽�no�n�1f�\�<�F�ݤ�:�<������`F���K�����c=���I����tѺ�`����85P��⯒�%�)>h/��.t�H3wU�F�7�uݣ)RL�K˰B��	tRjЅ����&��Z�U�n����S�Rk���:J�;r���^]#�V:��qJLVm
Nz����Q�{��z�Y���o�_��*�q>W*z�v׈�N��쩺)Nn�z�+���fXי|[����=N��:��U�J�s�7�4􋰽r�r�>rr�8�>��ۓ^��������T�P����a��w"��L����Tl�b���@��𼎑O�X滖�*Z����;>������!*O	��4^}]޸���oB�:+�)r������}���A[K76u�C`�vj7,�M<�kƹ�9Y�h�/oI�F�IFk�;����T�A�K��!'��k�`Ww�#+t5��N�/��R�&��D�ۥ�.�ƛ8z��I�}YQ;玜��7��!./,��՗eh��Y������>j�[Ww�J���>�6խ+�U�O��xA�aYX��v��fTf�i�H�WY5!�`+�v>�ȯ���{��@�Ir�V+u�Z�x�W՛�]�S���zg�Z��qGm���+�d'r��l���� (n�� tE ����Yn�eE��GQ��9���{2��g!�.�XG^61\T���jX�ċu���F5I!����Z�s1>�p����E�V��B��N����"�W�͡��Ur��$�%M��n�*⒐�����V����b�B���(_b�{��֌�J�Os�9�R��{9���yNp���
0:;{*cBV���e���:�ch�G[V�R�1Cص��ht�z��l�6	�RU���m@��t0����H���B�����f��Kr�e��:{|M2��v:���d:��:��0��4��:�,��
K���G4U�o�:��`����l��37 2c�[i	�������p>����$O5�&����.�cݯ6�h���κQ��qBCƮF�r���:f�`G�|5t�Vd���օ,��Pt��Wβ�lږ���V.PY���TD���ՋSaD�����[$�����}hKpxΖ�҈3X�d�}���@��{.��%֡j�T/6u3;�����d���n�xi�|똶o�X�7̾����rN�SI��M4�GE�{���Q��-i���nWX�*>s�Tub[t*�+�l��5bl��0M��À�2��{u�'0�s�L� 5��{����}��{6��^T��a�dR�׌�#T|�ؖ�-�f��Fu�,�z0T���;`c�� �M�acvʞ5�v��i�8��`����]y�R��ք���n�c��<kt�Ѽ�vL�	���Y�b}�#��ю�<��8�P�W�����Д˛�M�Nl��K��f�_(~�yaoA+�z�*5[%n�A���{��t��V�J<���I��%i(�{��l/�P�^ΐ���Yg+�V�J.��j�4imj�9�pm뷘
�)i}�j834^�M���/��C#c\�!ժ�Z%��ŊG��IZ����P.U��`��7�`�>$,�K+^��Cbij�e��32ؘ�.�6�+	q�KC�U�؊Ru�/���l6�읕Y�.j��[Kk[�L=����#�V��.B�]u��p�W��x�Z��(���E��@��-Ә6�,��J8�M	�ptu�i���s�s�6kJ)k���vԆ�ۮ�˻�cy�q��"�k2@q�hd|-��nd�"�Ns�uJJ�0�3{[�GLU��v�ѶB4�i�C9��qS8� ����m��a'S�Pt�J���H��ڋY*��U��Z(��R�B�ET�eTFҖ֔��5�E��� �(�����`�V�c����"�C,��0���IP+Vi2��PE@�2�V�j(U�Q�ث�V�L�\J։L�\�ˍ.Z
�B��1�"���q��X��1�-bV���k*1�J�L(��]!���%2�q��V"%�X���i��bW+h��*���P-�J��Y�-�S-�c1
�jU��d�QƹW1� ��am��b�˗2�""�2�+E��[J�8Җ�mQ1,X�nZ#TYP�j(#%h+�V)Z5��kc+\IEkj�h���<( {%�Qʗ��넘����Rݲ�<LZ��}���9���&b��0�(S˦��M��%���IV�{�����tQ�8�~�����qH*��E�Uw�jGk�{�r�.�����8�E�+�{np�*VM-�Nc����+��\s�����N>�C��S_'�5��+��+��,G�\��1�pͷ�9C�B��Ԝ_���a�����
�(��񨝽p0�[�F���qW����1B�[�r}�������aɍ�%Y���-,�:���v��KS}J�=6㕝U�oo��Z:c.Rk�:�yک)Δ��Z�z+���L����u
���';i;�5��:X&箻�9��M��g�%Γ����gf�?tC�T%�~_gQ��b���h&'2G,�
uu�,U�i��][�����e��ж���0oTI���쐪B�*��X:C���>���C����ݼ{��B:ܫ��PW��[Uک�W�t��c��w��;}ws�����N�}���OE�S�\a�y�����ɰ�p2������hWj���~\*	�p�Ϫc��ŕh�&�+��z�j����b�,^Qa`�'i,���huOd�|.�+�X�JHJηAmN���ޫ�����\V�PK9J��-�y����ז��yF��wr~��^�YX�!Jxz�w�@}�CU��-v]ﻥ;�֎���^l"��cץyVzm���{gR�*(���!:�J���'�|VW�q������G���Xk�Ej/�9I�Rc��[�im����bǵ�N� ��Ф	�������\jl��u�/uD6���h����y���)�o�7��8�,���U�U��0�4#h5��11�]���}=��W�y��7,�g�wx����b��o�I[	�a���3-b�]J�����Os<,gs*5�?�m�l����].�Rghu81r���vx�m�U���i�W���W7�\t\�W��V��c$_7\�w�vC�ׯI2�I= ��[����i;y%��ƞy�U�8�C����.m��9��%�r����P�'۞��M���쎫C�=F �Q���{��|#��|s��2we�]���W{}�6vΆ'z3s1�������1���Pb��wi�~ȑAԳ�o��kF���r@��V�wn�>ror�ь�R͐ܔ8�H�.�`��t�2cƃ�!ͮk��ȪTd%�x�����9�(WS}�_}�{�p��M7Yy��k�{���YI����M,uoP�zA}űvsc3b�^���8{����>�}]���o��w��[���S\��6�v�)�jz{l�ڵ��9]NT\pޡ<'�EsV�[>V���Ko7���e��u������H�Ǜ��{e�H��Y�r��k�X[��Q{�FPL��k=��FF�����N\��!*�b�]�}��+��-��Ǔ�[9iŜ�q;�L�E¹S˴G9Ჵ�9���f곝��Z�V^�eVs|�0�[�!�v�c>��	f�G�y���7x�ѻG]-�z����c���kݱ�er��IӸh>Jn�1͞�o
f�hTM<x�-lQ���y���x漳�XJ��������NS����c��y�gr-e��^�ˠ^�IP��^�kV��V&�S�s��< R�rge뤆Wui������*U�mM�h���um�CM#�㷵�Cuet��쫈	c���q���U��P���;��b��6�+X���sF
��y�2�%�0��s�j��ʕ���*Ѳ�O�x�"���:�4t�Ϋ]�菾���/(ı���z(�}�%���/��/'+�^�W�Cze�Od\ΓS����n��%ڲ��]��[[C�m�h���-���2�}d����gy\�4��6�&���g�O~�37����[���k8��2�DӉ7xD��箱�繶�̑�����[{��_��̰}MvW��ڻ�����WF��bF��jN���UU�s��vow����8h)�>�}:/o�7���p�qc���㮶{�D��T��q�JN�Vy+��/�5���s����6Pە-ׯe����c_e�\l,���y(I���Id��I�J�A�Y �Xgr�$��b~J;w�i�n�	�.d%��WY)�:�:[��Un_�%�ۜ�I5*�2��-�P9L�úb�X��~P��۰ֈ����?B�kZO�s����=�T��ʞ�v߀=%���KwGYȼL���f_HG���M!1���f��
5��]�u�G�e�8wSi���#)��m����;��4
aG�@��U���;8%����s%q��#Tb��s9�J)}�G:�3;".e�A�=nua���/��&J��!�p����ϼ���/^��D�<�]�П��R���p���.�S��/k�%04��ΜJN�΢ȧҷ&�=�VW�8�o��j\0����ox���iƒ�җ�!y\xK��g<7o��K���9dTb�H�W����ua�b���9��`.adE���Wm]^��W��,���^^��������TD��y�P[U9o���t��~�U������W�f���=��e�5�P�t�C��Q��̞���I��c���!o(w�����7,��fmY�1�t/P���퇲�횝��yn}2xO�-n����.�GTj�#�>�{+fUN��N�
)�c��
{�4��-���Eݰ�ux���=}J��t��Ϊ�	�İO��FLd��}8�������˙�W; pZ3�T֪,�v�� +77 t'��.qZ�稰��=HЗ]��^�s2��{�,�ip"i�a3�hhxu��ˡ��e=�~�0�µ)t��m�0Y=[0V�=;m1v�w�,����`%��x��bVp)j�m��WF�S��4��E�u��GQaV���<=�ZN��l֙�W���Kx��˰�����R���L͔���Ի$��M�ׅ�����>O�Z�{v�{^
i��V�ALƍ��o��������b\	��M���
��si\>�x��r��+��'	=X9��t�9�G�*B}Y��\U{s��O���
ތ�[.���wl��׍�5�	ex���f���,)כJh9��^�Ȑ 6�kw;U��9#籕�|=C��>W*z,�^!}5�D�̿By��dk���,P}72���7�������^\�����g�8��^4���S�f����/o��T��5�������I�6��Sa�F�O6{,�v�oN���k���p�Gܐ�%򰣵=�A�9�7�������
��Cd�k+Z�I�K���8�D^b�^=��`ϫ��M�0��5S1�\PF��Ȓ�Vo�_Ӝ+v�*��x�E{_p���gg�v���A�N5���4u�N2zIt/�K���֕,�(��O��ՙ�(�#<�ܽ��31=)r������$�u]���y#u�d'��0�[�G��Q��n\i��?�꯼�OJ�|�o��O�.��m�O�
��a�=�տGKN�w{�k����%{��O/d��Y.���v�8�}:1t�7F�0��t*�.���7���7+�fmy�{��6��{(��!y�	ǐ���^Gݞ��ڝ�Gc�9��7/���+�y�wЪ4��ݍB$Ҟ��v�l��w����ΪW�&�bv�����X�'���ΰۈ���<�\��}�1�V('_wer�[��[�������U{ؠ�)ټz�t'm�v���cx�Rо�k-h�V��ЋJ��{�`E�KAzv����`��z�F�W���l%_K������y����L�{�n:���W��U�!9��ї���9r�G-�	f�ʾ�5�앱\^�i�E�n�B���F��kyM �S�98�o,�
���������_=���M���yщ4V��u���q���N��J4b�5�2 ̖��ԁ6��oU�s��v�Ł����::ʎ�՗�S���+��R����볼E��5���$6\}�Nk���E��|�3}n �Ec}(	�3+L�c<�>�UU��&�5-ۥؽ��̿��m�k��z�n:^B���A��[���Nx�����H
�F녠��Mb{��eG*Q	:v���P͑�JbK�nDr�/�Z����o��2�"[Cy�K���\��]�jҲ�
S�m�#�WMUt��-�49.a�1/�:�����t/1^<�[k��ڸ�
3��3��N.m�M���Ɇ���u���`㺿c��%j��j���1�^���r�\����b���mi�Õ�7(�(⺹�ˢ�Y�e�{o�|!Qpr���E2:=��=�;קǝ�y=���߹�smC�����)��U����e!uH�<�ڋ8�%�W�κ����y���`;�|z�-Z�t4�yB�\����eJW��S[��c������5���<e��#�u��佼���礯MT%����Yg��[I�|�io���&�.��i���"JY�{��S/�Y�T�Fm���F-���V��sR�ƐP�{�a��Ճ�74��>y�R�������wMty��џs�"��kX���[	�ົ8j�J���ڤ�(t��%eG'2i��U}Pt"]�xS�������*��+l zAѮ�	I�_%Aec��9"�"��M�ȓ��U�\XS��>ʶ���N��
�ꃧ�U]Iß�܉�RK[Һ��t�4��w�5ɥ`k���dӤ�;r�B_%�e�ZL����Y��^�ku�Z�<�O�+g6������+��U��}(�]Mk�8Fvˋ.��N{�>�ז!ve��:�iu��wu��$�1���8]Q��f������Ǣ�v{�LJܜ�O�>
�0�j�������U�gz/w]�:g�����U,j��7���6ǯ����&]�KTĮ����K�h��4��Wmx]^��^�f+I���V+�[������;���=`�۔�����WEvQ�ޠ'ygB�=�K�[m��9����O����9�эGH{u5���k���3������v.H���x��U���\�M��ݯM�J����
��+q��P�km���T���D#���p>�f�vt�_�̙C��-]p�[r�K��f�2�y�;Vlt*z{�l�eΫ(Cr�1b�7��-�P�����h+h�>8�Qy9_/R��}Y�P��}�^�7�OE2[p��O[@���J������N��C!��ą����[2�^�r��e��G픮�Hw|�gPN/7�Fy��&�q_m���g/�,����mڥ�E��J�K�V.�33Z��%�5�P,���#�lg(Z�Y�ոP�=|�I�U��R��u�_&�vz��
o�mt.����R�����W�Q\�v��^�?%ϖ�|�=�׫a��lmzն6�)ʊц��#z�0d'��U����������9[��ͤ�;2ض�-��*B�or1��<Y*6�m�Z4$x�{HB�v�t��U��P��[��ݵG5�5��y��	���ג�+�d�J���ft'��S�$�O��[՗��su���
�z�e\��٤'"����	����RW)z�Sa]�E�v�F	#B��u���G�cu`��F�$+(���ZK)6rރWy� ��C ���ܔ\k[}���VW1�Wp,M�|��OzH;Z�\��G��tM�7*St9�X8�Lm˒��\|f�.lپ�C@�'���Zȝ�Q'mf���ds�&��%^t�:���qպ�sJ���#l���g%�g(Y�r�۔���+_,Li��Ձ���e�q|o0�6�n;�>�� ��ݴ�\��6�"X.����`��@j�G-i�5 ��:H�n�Ό&���R囨�h9:�d�#V��P� K�����s &j�c��2n��:����N�B��]����3B��6zŚ������9D
l5Z^]�fP����lh�2�U�DN��c^�.�]-pI��{ׄL꼽i�j�gv*lґK��Z��B;�2r�=K �N�i#Ybr�N�f�nfM^��D\������Z�b�f�q�ɠp��gt雬�Y,g�J�'(v5
���!�;��aֻx��	�G\EfF̾�Ҵ-��c�ҪL��M�.��������]ef39o.�a��V��u��OO��zEI�+<p�4�V��5�S�|��N��[��"d�h_�V��(*n�[C�Df
�d�wg:;%JWU�Oz��l~�[ٳM����9����$�衤��
�Ͳ���L]w�ɴ;Uo/0:�2��9�2	�>���r˩FT�(R��8��2͝
�,�W}���|�"�7���8vM�s3��݃�9�r#�Uok��'q��r.9���-��������lwܞ��oQS�<�C�S+�=����# ��EY�4
|�)jk����&j�o�9��U=1n$�$�8/M\rC\(��cx)s��.V�0�@��B����-s�<̢��	���(��0��X�i��[/�
���ۢ��<9cq�Tm�#��;[�	R\�
��}X3�:8�4S�2j�mL��G)v�[Գ��b	�wi7}6��<��#0�j�L��3���3)U�Y]�B��b6�:��ݰ�e+s&s��e��*��] r	g!�p���0��^Ad��H5bK.őE���B�ް��wt��5O�P����ςrW��Zf<���0E��/m�n�N��S�#K�.UZI���42�A��
p�fV^��ز�[�1б8��ɶ��ܵn8Fi��v�ԗ�(���*�Y�2���[�dn�!��x]*)��d���Q�f������'��e�W�Kˎ���L[FJ������W�����3o���]��*܃b!]<��� v�|��@u�X��Y��q��,G�T�fJ�Q����8�{�$��]��16|�uu^d�����&n���~�5k�k��,����5>���r��tbvP�ME�z���l�*�H\�X�z�e_`(��,�l;����A����/Qޏ6�fU*���TA��V0W�ŦZ#"��[kmEb��E�X��iPq
*�1X��UU�Kj�+,�eE�L�T1`�X"�kJ���(�DKB�b(T���1EkE���������2�m� �UAb�GeB����[Y`�6-J(��f\E�Ҷ,���S2�
�D,UȍL�*��E�cEQTAQ*cTm���ʨ�jW-
�3�報����s02�ƊDTPL��ն�2�( �媨����T�֘8
0QQ�X�Ș���X1���UE(*�TUŌ@
�+Nmtݙ(�9�wү��}Vb�;���En�x�����n�]�������\��Y|��8;�[���<��ї\i_���Q�;P�'����5�T�
L��ڞD�c�A[�im������;�T��3K[�lqy\�2������)��#f9�נ��;�6���_*��~6}�߾mx�r�y�*�9�Ui�n��<E4�/r��������\���B��װk؁�ݍR�|5�:��.��֑Η�Z�l��h.;T|��R�1�_Q�Ԝ������Rܞ��T�x���UCi_o�ą���}�u�f�����=�cV�M.qB�,�\�t�{���Ҿ�j�'��8��<v��j{�-��[�����]e�$�S��efh��|�i7%�����ʭ{���{�ת74�h����Cu���c���V�C�ɂ�h--�+��v��GM�wV�BH7%	�&���yp-󱥼�=��m���e�e��Z�8a��/�����l
j�h5�OSLM�$Z�D�Ȫ��+�;N��� ��
�ɸ��K�D>�n�$X��k��6�3�X�A�@է�pB1z���"6��P/zo[��N�(/n�ݩ�V8�X2s���虪��F��UQ���Y�ٜ����������0k�%)tVg5�����$�7<�(�ъU�ݦ�����C���R6��2�Qk�_�G+��w,s].�.t���O$�v��dӤh��|BU��	��L�μ��q�Ug��N��=ԝ�j;_=N�7�cut�'�oP#�$��KwNL�G-c��|�2�s̱��Ml=�r,c��ٚR�D�w*�ݨ����'3��ǢV��"{�k��Wڪ1��� ������O��
�w*]�ͦҔ�N �᧵��uD[�8��|��R[����ߜ�e���&�������R�`�~�$%�EnW�s�����{V����Ee'�n�vv�.�֢�Us�v�v��ӌ�{��^:/iX���/�&���*ɤ�9��/y��7a��эGH�zS�x9���C�ۥ�WAdMׄ�z�}f�IW ���u8��kc��<�7s��Wݽ���i8�%�Gf��3^_tB�6�Xa*�q���P7y��H�q�ձ�m��*b4k�J��ڕ%�[��;��]윲Vi�k�tW܅�^m�B���h�a�%L����ٌ<y����ڻܥF(K���S9��k7��B�}M�s/�6�Ӕ#�cX���Z��a�ͱ�Ѭ��-'�Q��7�r!�~=���V#�Q�T,��ŭ�u�n+���{���%��t	����GQ��5T����f��B�q���ܷ���5f���. -{<��{�JEz=Q�LqP�T:A�P3�U�J��qϛ`o*3z��o9����気.�OyMr��+l zN���k;�{���� ��o��n2� �8�Ĺ�M�ow�i��������B\���J_7��\�س�9Tt��Z���:B�ٮM-c�/c"�%b�W��s��#ȗ�=�O6p��#|����I��\�ֵO�s��|�۵�n�HN��>÷�};<?r^�]ٲ󟊼]�ow���;��:��L�]S�VjJ��l%q!\��٤-�)���.�N�峽m�d��Xlh9<R��٨�E�-�
ZY��yN�&����K�Vܰv�i��Q\�V���E��OoO5� ܘ���q��^��r�XX��k���O��G��/�^q���rz뜙,98v�A]s��D�<��[�����"�<�*��P_`������X�Iz�Ⱥ�0^v��+��󋔲�J�hrʦ�}`�u�h�����h]^��br�{�j�V�rʕ�`������O�}=��}Aw�{��ϥ��:,��X�/P��w��۹�y9^���b�'8�`�R��jÓW��*�URe����gA���;�oU^Nb�^�7ԜXo��c��L�.ƧcI�o����ϡ{
�f�߄=g8�h�{���mt�S��Eٞe�{�І�>�3ڻ�Pܞs��*��1n9<=��;OK�c���-�ښ%�q�ة���v��]R��j)��w��#G_nk�w&�7Yx��\�e���^&�Z1��R�[B1 xk�S��y�.���A��]*���ء|��[O���Xanߛ{@)����VԂ��Ju���Hʭ����� xkV,�����f7����y�伀^1Gy�̗�k�yۙ��R������R�۫AVF�N9�B(Pfn�A��l����+fdqa�mn.n�ػ�Rod�����/�9λ�v��2f�5��SpW��__-W[�!��(k�P��[������Y@[q�by'�������彋m� ����*���p���&���2f�zC�--Z�=�~�F�/�L62}N����V�X*f_?}5y�[�z�V{2��`z���Ҫ�eۭO<�VaL;�A*(�!<��+rƣ�v�������^�*s���^��h'��m3aN�'�i8�_�Pink�Vq�5T�r�R�cBp��n���r�TqU�m�� . �g���EsLA�靼a�F�:%k�[�>����ܪs�T����S�����0٫�<�<��!�@ˠ܌Ko1P�{^װf�P�t�^�0���
�a�������xEme�7y���ڡ�o�q>}
Ŵ��mQ}�C�f�y|�t���-��k2���١��,����Ho_���!�Nގ!����w��wD��A�r��]pW��pI2�����3���b1�C�m-3����(��ȧ5���vu>�85���#�����1A;����������g�������� �ZZix�G^���
{
��lq�f�Իkq_K7�W[�L	��3�R�:Ym�/q��j���}��OcGJUՄ�Wf=}6�n��C%�vu��I���>ܥ�ݬѯU�w!и#�-�Lu)���j�U�ͳ�9����r==~�ޙU�"�aՎ,7wՎ-ܶ�8�B�#���	@�;��{�d�[�cGy�o4s�~=�֩��,���0���n�
f4k�(J]|�Z��oYУ6���8n���U}��*8X�i��¸�w]˺�g�t�.JGo]Z���Q�v�����Hv���u�uX{"�"(6�y+������!�.�m��قv���T��e�-n�%4�S�y�֜b��g��H�˷�P��~�I�A�)�>�ܕ�8���#eɵ��E�fA;00X��oDS��h�UU��c4���2�'��+9H����j9����ouT+<-��*�#�߱��O]9�G[]��wí�bó�W��wwI����9}�:���*Q�l`�m����8]��Ǹig�n&uv�^oii�NӒöOEے�sTc4� �Ut�`毊��QJ�ǫi�{��&h�+�z:l�˘
V\�6lme��ǵ<�b��)�;G0�m):�t���E��-�:-�o=)B�ڷ)s�I\�������;�SA����3����K�l�����+r�s�K��=���Y�z٬�����:��o��E�������|���k+�ׯ��:��"�spOC�B�+�r��fˈ	�;�zSk�kQ�����Mx>���3(�p��04�_P�3s9Ȥ:���U��1ooP���v�-���ӡnF�Rf�U���p��4�jxP2.�O\��u�8�d����w٩����oS����n
����'���'���o�G������g��Z�\}͜{�/��kS�zU>�4�U�&��1{�㊄ʢ��B�Z�,�V���g�	��+0��5�SG���]����^��Ё�<5Д��3��uM���s�k��Mk�]O��Ť�gc[Ni�n�C���PB=�^�/����g���GK*�V�ce���
w�Q��9w��W�0>6mk��u��=�;�iXja)-��6X�zu�y��V�+���b}�r��h�dMX"�ᶎ�������C����s�����0���
���F�D&�\�fGٚ��z|��hriX�\�i�e-ܪ
�F=SFu�׌9�xB.wJS	�`\�ֵ_<Jj��ox'�Չ�_N]lB˦2ZE^�h�x�Ѐ�(�U�r������.�;M�5�^QM�]]��)���ИօceY�wa���=���7�'kz�'	���um����൩����l�Qq^s_s7��xW��KN6��i��N��m󡚘������4D�LvY]�it����j8h��׾���+ݼf1�=�{�����*�z��w/`,����ţI�7��j�4��u�J��^NP��ȬBGu7}N�t1��T����Y����F���;f��H��+���y9^�1���}I���]
_&���vW�8GJ������<��ߡ����@�vqg��b�˧2u6֋ᙶ�������H�����4=�*�>K��w�b����D�����2�NfV<��ىqq�<x�Uu'�y6�/l���Xt#�]�cI��r�*��������1��g��0s&^]Z��lTv�[8��G6�K�6��!�l[^r�qh�or{��!x|����]���U1�����6�7�Ӌ�S�����EW/��Y�w.��n�%����z�^�{����t��Z�	�I��}�.�Ъ��̞j��y1�y��-����8�J*��e@4�6:Z�.��q��f*z\��k׹�i����U��5�&;�)�X�;�V�k�J����0O=9�u�|�函��ҬAR���=2#�X\��O��3�����o}FHB\�w�)|z�]#̩}�����]�.̙�%�&V-�߻ӆ������?W�w=
���h�W����T�ssםY�˄��nWbq��w�I�Q	�f�<L�.§��q�E,�f�!u:��_j����hsK�ǷVW*I1U�}jn#d$��F.���@ⳄҌ��Ĩ+a��=�t�� \����s7�7sm��3.�~׎��{M�<=R�5���ևCq/e[��Z9śQ��!o3o��=�RnWX쵶����vm,	Z�q�R������vx��J�2�kȂ�����|{(�/k�:$��v��@+�jH�ά����S�3�(a���ޅg�f,z�;�T|����n�Dv]�n�g��[CsdV�;�ܠs���+�i���]YRo��`����K�g��(.hu��1�6CwS\��k���]��s����o˼����;�wg}R���T��N�z�N��Q~�7p����P��î�{�<����I�;���sq^ykw}����܍ꌼ<m��1���1�g�۫S�:����d:�9Q�X��C�������xv�c�M�S�ɓ�,�~��6��U���B�s��j���M5���]٬���u�CfwgS���K�p􂷉B�xH��*��:���Tш�/��ܻ���\6�n�X���S0�����U�YkGK���Tr4��Δӫ�uӼ�<��y�籒��q�K�lhH�bNz�k�J��֬���S���ٵ�wI0��K̶C�=�欁EP�-�60Q�:��od�Jy]��[���Y+���q����дe3��\K
�F[{g���r��;ٰ�|�ts���m��+��9O+RJ`���h7L*��]B�
L_�V���{Q�k�ʙ(Lm:�M��6!Q_��&��b���Mw��8�=[޶�n�Yq�g���i*AHe��)���T�&�&�z7:�Ҝ�ʍ�py�)e䫽0,ޙL$����0Ԛ)U�ػ��+!l�a�U��G��.�n����a��9'S]�4��B��N1�˭�R� ����� ����o�Y�*��ڋ.�;f�V�@�Ğ�'�J��E�������杁�Q�Q����PV�)Oj%v�.;x���r�e�36������TmR��gi֚o9�ňV���﷑�#�+-�X}Y�9`Kx�U���B�4w�Sy�>��щܓA���M�{P��4{utU����PN�G�Rƕ
��["vP�R](cGi+y����C�AV�,G}�U
��ϝ� �@s����-�5Wl����Рl":V_p;��>���y�'V):�¤Y�+5*��7RصG(�A\P��Htgct.vY�/A�H�cX)�p,��X�q
�Z�����Q�/1NYkr�'2�&j���E�H��k7�`Q<�:9���Zv+��M5�2�)u&^`��ޫ���B��ڳL��ӫ:��L�Vb��`沂���[r����F�X�f�T��%����;�a��4R6�����V$`^]v�f��vފz��]Ȏ�zq]f��P��t�)a*o�wfZ6��S��õ�}y`@�/�jý�E�$�&�u��'��sJ�m��6Pr�A�Z*>\�18��z�/7��2اu�.>PX���Ց:+/�Cvk �=�e����f�ɼ�܎�a}��y�d��:<G]
�n�L�<��yd�	�YMι-��Z��᫮
'��b��^�����]v'����6�Cr�g`l9�����f��X�y��3��ܫ���(�Z�`��!u�W�������R�\�=�4�����K-�=T�a�Mn�w.��!�1�cy�o��0a��Iz�;��	��ȹ��\�T�l�9j>�f����bެp���
��6ep�w&ښ��z9��y�4�K�=[X��W��qE�x��qŁo${x�����
͑��(]�[���^�Ők��o�8ܠ|��F�����	�tu������67n�v#Օ�v���=[@Vz���Ww{�%�y��2"D �	�yM4�k�ѯ��\뒜c6ZWjh�vL�m˺���RtP�r����f)�&���m�=�Y�G%���h`*]/M������n�����s���j9O�3��MlWX��{έXH�ʖ�J������6d��ζ��K�jhm,��=P�@51���EUU���Q"�DF�F8�SR�2�.aJѩ`ڥB��AQb��R�b���E+Y�kE֨�X��"�1Ln&**���U�.4DAEq��0�(�ȵ+�&X��X�S*�c"�1��EQU�"E��(**,be�Q\s�X��,U���$D�+Y
\��m�����QDLIQb�b)��E�2�R�UQVA�AER��ƥB�Q���(���"�Y1mX,�*�`�ܸ���l�Z��",bc1&�YT�PZ�e��ee`��TE����T�h��DV(�X�Pb��DS�U��BcQUUb���QcƱD�[��TYX��PU�E��-��4X��V(���UUR?]�ݾ��;��!�9�m�1��fN�NRW��,[�#̬��|����@;�e��ՠe苌يmf�5�"�ec
�^��˚���9~�]���[i �2E:F��W�� ��G@���D��ܭ��|�F녙w��[C��u>lrqk����\��z�^ͅ�b��Dm^<ȵ5�=����2��e$�CJ�i�|;�oA�;�]ǻ14ҥ$1��E�4����'��+9H���4r*b#��M�F���J��L5�z,�9��	[����ڷ*=�`B��yF����+�c[S^��k�t��>��G5�g��]�y�v!��s<*9W�IhfTi��h�P7��;�j���j�\G7_�Y�c����UJ����6���'�oP��m�ka�j�y���2�����j�s;z�,�2�ͻ8���c����N(]%[^}}9��f����	���'��,o�`�g��^�,Uq�J�V��Z����5̵�,��
��a�u�ؓ�����y]]-��4�^�{�d�q�\�����bȣ߰����o���7i��nR�d/�K�[���D�X���u)�'XOs�����:	��Ue;ȳr?(��{�(�@���U��	�6W�g59����&|���C�%�ڙ�39|B�q��E�Y��5���Q��5s&�SFs���~�zJ�5(	֮9!��+FR�۩���������-�Q�R�e�;O�+-ek}$L&�:���`n����s�|��h>یoh�u��W9M6��yS��qk����Wc��~��i�����ٮM+�j��d��%~�C�u�e.��9��\el���Iq���B�v��g(׫���
Z}t�KCN�Un���ˬPV�u]q��=��Z���	�ݲ�퐊���s���c���[y
�W.z,��-�%nMOv�����.�W<[�xxv�Z�7�ǭ�E��/�`~:�X]������Mdȋ�V�����{\�2�8�m�R�1!��Wm�Ҳ�K���3�BN��,��,t��ۼ�f
|6K}B�w'�B(4,���mqM�Ck�G)͛��6�J���r��N[��K]4o����h���O��polf�]7r�����ёc��\d�#i	.�n�.34p�>����1r����q>��)5W�e������"m %�x�rNͅl�|�J^ұj�X���&7��qphl�f*l_[ف2���\k��xr����(WoWz�pb���Ԝ^T��⡕t!�̕l�|����׼�+��}�T;t�Xԥ��_��3{َ;T�ǫ����7�q�^f�����=5�Qru�ý��h��{k���5�=��r)�x��|����M�R`�na�}��T����I�ӭ��=e����p��Zi��{]7�~�!���a���S ��]���⠫�s�Χ�pYN�O���ov�ck-����5W����I���*�c���9������|����
�׹�����$�Cw[5֍ԮU��M!���:�TჸxT��=<O;�\�V�����EJ3F����Q=Y� gvQ�j�$c�y��Qz5*��J��}����*��:��z�T�2�U�au�i���w9�7V�{��V��{q9+(�1��+E�d2T6���
�*>=4tlA��r�HTǫ5���>jZln�1d+��s�hF���r3��;T�Ջ8�s��x7v���'.U��Gt�����{;u{��9D�^��%��\�'�5�:ۋ���z��eOF��h�e���6#1��m��ohl=Y�9����OS�|���
ò%8ػ&_��螕��լ޷��84�_;fb�{c�V��Q���L=�t�@���P}k��H�oo��x/�%�B�o��K�ޙ��{SԨ��!��s{�C�
�������[����ڡ�\�n�{�A��{���EI"їGz��֫#���n����ָ��Gյ>��oh�*`t���V$����t���>��s/6rjR9���]�$�̥��_:X�L���]�n�X�ܜX���	���ո6��fV�b�	.P2_9ASR��˜�8�Y�C%���jM�{˽r^�%��J�{u}��}�TRI�\̬6]vJ (�yÍ$�0Cj�B��S�8z5/)�6�)���R7b.�Qz��gn�^։�ݱ�2�J�::�;�/��\��H��۶Q�(���5,$���=�c�K{o1\+%��=������$	k���s54?U3o��6���V�v�	;[r�ڥcW�-i�ͻBz�S��V�g$�zV����8���m����?eV�Wer��0b]��u�uG�tk�����Kv�}AMr�GY[ac3�$��3�iF��i�Þ�����ds>�x���3C�*��D`� �.u!��g�,�sT:CK�Z���3	>�N;����)�g��������̕[�,S�se`I�ɑ���SO�}\���[O�ݑ'5ؚ�2Vl������D%>��Z�m��=I������,����m�nK�;��<-� R�z,�^l�S��[�^�O�Q��r�Yn�o�B\6���X��"�6z!��Kh^t�xgֱ���{g�򡵸�[+�Y����*m��;GH�+r�s�y�f�S���eC��C��]�Kkyu,�n��e��"�G��f>��U}���-W�W�!��[l��Wv�K0.!J��k1�GmL�'Y���|y��sv��F���v�v%��k��i�\����2�]8�v��f�5ٙ� �)�VӋ�y���[�F��|���S/���ɋK-g²�ұ�a��1���{~����uNz�2��NP��Eb��n�s��Q�3����'X\]u2مD��{qM���	x}A����}�WR��_V;��`n�)L�7�ug��歾]���`鋨�Y��g.�:��C�κ�Z�Q�z1P�*u��uҶF^���֖�5}����nWe�<��my��m��G��*Y7O���U�4��{���'�s���v7e]G�/�QW�/*����}P&5��G/3_�y׎�XS��n�o��k�B�+T�;�Рn���﮳_�.��#�����vQt��qŪ��f[j6��ut$���wt̓cr4-�W�Bq�zzg�Ϣ����z�z��&�cv��r�-��N�\��S��f����⼇-@��R6=��Bj�x��2�ɛU��G�r�#mĵ�^b�f��n�D�Jπ��r�z��I�C܍��|�S��,�"��`��j�Qm����\����	=(�]][�.�~�����d	��+9N�qĺ��l�n����:B�;�o:�*Ƣ�,ਵL����R�ӓ�����Yټ�K�/�?ѓN�BR�X��`s�WZ����☃1Y!m)�0�������p�+�wy�
�F+��@��9��V�����U��r]7�iy\�jҷй;JV��Y�4eQȾ+oǒ����7c~K�S�}��׶���S���{;�'�d�ԏdh�Fr��f�#�F�f�}W}B�8�v��^�s
����[�TtA�E_���-�A��2�m|^�ķ�̫w�wKoySB~��v����%'�uM��;5&���O9�V-\�J�ďR._YJ����gq�k;��[!�l�,9]q�E[�UO�o��Ѹ+�U�gg<J�s=�X|#[J{�n����t�uyQ�;)Xى�قh��>�;���͊�����Yi7^����{^��~�Es~5'<�}u���쳴l��u��_��<#�҃�nAY��&�F����:����xL��]�oв����[��g�u�gN�J]�a�K+���v�(J���X��gX�l泖��N�N�a�x��ÃV�$��Y��r���
�˺�W��s�[����W�+������F)��:����sίU���j{{.vg&��
���!!*��(��-�`MO#�n0�]���\yב�Ϻ}�ё�������/Ǵ/�]Vq��g��]�.Ϯ7J�D��k��q7�zW���F�{�ǌW��`{�v���Oj�3�lS	o��C����xYYR�@�����G�O �����% r�GB]��.N┺H��A3����~�R׿?��Yj�s[��SV]m�[��}�\�c�l��� ��^���uq��~9��%�Oԇ��Z.˕$\I|T^�B��fM��K��;�Gz�3����.}�r!cm�\u��+��Dzr��s�;[��j�~t��� �T�r�{@@~��7*F���1`�S��ϑ�5'VN�~��:����Gm�|�gĻ��K�5�@w��W$i 9�7P��L+�WIуҶ��mٯ���>��_X�t;��|۠:߶�xc�4E/D�p�;���*�׸���F�����t+��'�����ѻ�Q��Jn]���jY��euJ1Q�{b�^hn�ईڼ뭛xh)6#L]�<k����=o��"�ozAp��$%%Ӕ�/���s��%�G�&.t�F�i��![X�F(�����]�j�;��1}hN��~�ki�B�]�Q��@�>�^�X/���r�e���b�3�ƈ6��������I���T�T���7�(
�o"��x�di�}�qW�{s���gG����`cw���;&�������#s�3�k����x�mc<=���Ψ���g�i��$/{�����O�M�(,��L*����q�;�}���꡶�y�-�#��pf�}5R��t�\����Sz��/�d_�O���2��d�n�M��%ZY��eT&�S�}/�X�ޟ�F��
�+m�唂�n��ͨ� ���X�0����ѹç2k�2�!~������ĩT�������p��Z��+*Y�@:�����i+�;^�;�D{��Z�\��Y�wT��L��9��O�qϽӢ����b�������^*���t|k-n�U{�5����'�d�o�dS^��3���u��b�n���@q��ҭ!��z�����9+��ӣPO�Y���̅�ǯ�트�W3�O*!�H�^޽���}[��:t�6;,ƺ���qa�b�;
U�-ډ�[&V������ /��5��!�nm|�!��X蕘�����N8�.n�
k����{��y�[����6$SVE��nP@p+@�{9,ΕT:x��:3\]G;B��7]M{֡O�D}��+�Z;bD��]"D����ٞ�P�D7^G�"}�y%�{�5]{�)��Jؗ����Հu����� �l��d>4/�#�����/�݈�`�tP�	��O�Ub�����P�������]`���ީD�L�-�8o���v���-��v�h��6Bo��>�t��1�ӌ���
��*�ޏ�&�]A�7��7(z*�X��-�g��s��A��<4�����ww�^�.c�N�˸h\͝��z]~��C���~��9�)c�`�Ճ�O��eZ�?�ְV��s�k��`W˖{c�a�����S�����k)9�yǋ�9]o����8Z�D7��t�﫰,�)��KGQ~��_��޹}y���T�H�����O���`�妴f���������
��TR�9�����Ȋ�Xj>�ڊ��� kj�F5x�O�{ai���}9NT���s÷��hu��.7�k��IF�b���=�U~ɝ��U�Wj����̮���f�J����'��g?S��7��_l_�8T/b��{�W���c�ϦX�2)�y��4�r찲˙|yvt�76Yڎ��/Y��F�@3���n`3/gkvͽD���{����>�&�9Nq�+$}��,�����^��b;��E��A^��v4N0G]�ǈKeeX��7��Tr�f�]��$�^K�mfZ��(��6��
'/"t��+g��,N;,���X��&��걍�m���}��BS,�FVc����<���wm��[:�f�֥�s�Ja���+���^�	�M�ݭ]��ّc�-։�����t�Z]m[�M��%��m<�z�YF�'��+g���R���/L
A9v]�G�,��p���򆌅几�@��G���������w}A��#y+�e3��0����&2��C��#����s��͔4	�=T���9��	W��ņ,��6��q����l�jْ���M�Ŷ���oSu+�����6���x�+3z�o�ɺ���F��b0joH�]|���(�Z벩3b=)gQ:�3���.I;�;��.�<��_[J(����ͬ���ʵ9�i�#�z�kI��P
�ٙuۏ[W8��emb�z�)3O{nwŶ2�n���m���ʝԻ���"��}��#:Ĺ�������H��`��\�+5�u%l���^�2gf�
�a7mM�]�t�C�f��/e-�L��O ���-Cd�A�ƴ�PLU,����
���V;�'���-�t0���p`��Suw��;|R�Vm��S]+P+��V��uq%1�	� ���׸��7��.��1,,��f]%k5$��6���I6��P��>n�q��*5 ^����{o�䴫I���t�-�w;v�2���SC:{���jB�驑�|�Ү��5��ݻb�-s�F����Q�Hh����^]���M����f�ͬ�	 ';��ƀ�ɘ�+�ۋZ�;��q��r�2X�]�=��nf�b��;ْ��Z��隺mokt��z3LC��[��`�B��5ݬ�U,��i���z<�I7{����]GZqw\Z��V۷5D0>L6M0ↁt��X�����;:J�eѝ3u=e������$�E�QM��6:�z��V���VD��[x�j�O�E7�'r��z��#n�0D��y�QR�]ږg��֨�����%��S�{.�4�$�`�֊O��a`�	uyR͜_^�h�6���b��B��6��hѾ�>�r��]�J�,�}��'`ڶUG����}�Emc�����[��]���)U�ΰt[N��T��������1�(tr�Pّ9�yF�n&��t;�R�+*Tv+{+�eL��<
X[���,�V���T�ȋ|����v�!��)�Kn��Y�S,b�L*��(�m�Go%t���VWe����Je��T=t�k�c����|���$�Q<�ޅv�����{N�f���_;�돻���*`�Ur�Ƣ��FT*��Q�(*�\��U!�QDd˘X�#Re��T��F[F++EA"(���UUTD\�V&&3"�H��)-QUhV[J��Er�Pr�AV(����*1-�b0����E��(�*�*���6ᒰPQA�(�ech-h�DEDLB�TED�*��D"8�2V�Q-(��G�,EV1��"*�5q�QU�V2)PDk�,TPPTk
�B�2Т���hUc�J�-"��ePY-)���i*��-eH+�Kr�fU ��LK�J2"�dkb+-�啄�b�A��E�e��k��B�LIX���E��U�"*�ĕ�#�d��pޡZ�E�'�#�	������^���:��e��E���!�}����ǝ{fJ�Xp^_f������Y�7��L�>�˟^��F�SÏҼR>�H��+��Ig��<vi�E�C�w�6��ӝk-���ZԦM\��7�-���oև�>f{C�ӟ{���z����q��Y�݉����|6��r�yA�4z@�W��|Keq��e��#�!b�!c�1����n�>V1��F=Y�ɭ^��{��AX�����Ct�QW԰�-��	�j1�dŰ��*��X�+��=��{����芈�n@!�뉐��O��r	hz���=�G�/D�}ʣ�R��e��#޶ w�g��$�;2�a��
�I�h�^
����;S�W����s�ϴ��1������G"m ���&��>*M�30��Т}�r����=z���J����Fﶼ,gBv.6�n�nb�����c�Is�{$K5�g��z�����õ7�y>�]θ��c��uc��9����vnQ��_�oV����r��&�D> �D�q۝�^���1x}�~�>oi�3�~����F�7�ŗ��x�*[I��L�t����tGp�pm\ڗ@$��:\on�ג�t@��wHe�ԕ���x�ke%ow������׃i�B�P�P��u��;1I}y�#�C�^-�z���R�WlN��s	�1>���9�u�缋E��:�i>�:#����=y87��� 4mV-� �L���a߿��7~ƛ�,d�X���W���w�r�Y�����g]��Z��6e��:X����O���9�}����yo�6tp縡����7��{�=넍�ⸯvQ��,��Af����<Of��[^�
�������b�]����s/��r7��_�G����ym�D]�N-�ת�Tf(g���<}����7<υ��:�9[t�ϧ��y�|Ό~u�z�>�dJ��y�FU�g�ZF��u�YF�L�R_7T����|M��)��U�׸��4��.z:���"f�4u-���a�B�!�J���&C��'��_�P��t������
5�g+�a�f_�H��w[����N�U��	������ޯW��,��CsD���W��An�7�/U'��ϔsո;g�q�~�=ގ�>7ڍG\?RF���G�3��	��Vs.O�sq0Xs��ۢ�{�r�U�����t�@<=�O�_�����u��L��?I��ۗ"��9(�a�'����S�<�WTw.Ʃ�4u0�wu��Y�3���nB^+5���Y�����Kǲ����~�8[c&6:Q=V�#ה��0�uKr�z��9b�D]:�UB�k6 8�J�����jZ���Ş�2LJ�A�}��J�L>X�kk	�	�ԕ��;�RW���n��&iOx��>��r���~�}.�a}R�3~�V��'!�"+#�Ђ�z7s�}����7'�v��=ו�b�����|;�cm:�t[~���n����Ewx�,�݈�a��Ъp\#� ��eO�≺��;�Fz�M}���_�_�=h��*�^53�^H��>��5w(���	W�wC��d��F�cq�f��ݨw�^���ҏE�ё�ў�{�����}ٗ��E�s������=��Vgտ��d�u�X�./�k���m�nf���ў����4��︰&"��#��o�'!\���ڮ*ڣ���;�}�K�ݨ����f��юE�fp�d�V�����Ft�:�����{k�}��=��@�u�]�FmǏ��<JΛf�{�wM�xRʯ������;�{N�׎W��>�"�ث�<�?Ux樓{Mj�o�_��یv�{+����)�/	몇㊥�ɝ~�ژMA�vchm�>U~�&w�f�\#3�⻥#��ex+�Whh�{E �dJ��,%7��0&��
e�y*P|dұ�y��Q��Zkn
у��]<vi�.@QY��l3{Z"�E-k�%����;�3��l�0,/R80\��'�c7��:͝Wg�ޣ�:��-�	�Ƨ0p�Ϝ�pu��s��\�Q���t/t��z����k��NGod�����R\ozD�;���{K��g�=�ǃ�T�t�,��9U�;�qE��/Cp�c/_�gb��!f}����h>r���ՉF�+�dB>�ϸ�ң�/��ެ��g�r�/ :���G62�޻ŝ;أk�^;շB����Ǚ���P�_
�o�ه�/q�7�u#�;4���v*��'�i�l�i�DLL'Q���V�t�wz|�RΫ�P�{�8md˒�YY>�k:0�%}��C�C�ȑnQ�]�>G�baz��11O��p��w>FX��-����k��eg`W���\��7��e ^B����䕁�<���^����?Oڱ����K�5;s�"�n�b�ۧ���>�ؤ.!�׍�~�=�U`_���y�ODς���c�6�[�~�Kht����rCI�=��n��ӱQ��F���q󬻏d3�$��s��r&|z/bV\Qފ��q���sR��̜ѓ��l�&M.�<��dy{�S��:���wb�l׫f�О��T���{��߶�q�%�۝��ٳ��FN��q�7��J�q���׈��g�:�Ѩy/��{�y8����iW��!�d��6��V�]7��"�ʖ2�$ᛸ�F���(�m�\���k��3�f]s:�Z�nA!;҈ ]��}Լj��E��$��m�c跮V����϶�V�-(ۻ��Ҩ��t���k)N��&�`��B�Huy	���:c�=���N�<���3L��r��Y���H���%Ůں�D�[�G݄��:�W��Eh��wMė��ۯYv�ץ_��~`g���n��^Kۀ����_�W�n=��=���������4��IGn&X��tP�}�����2<�F9��s��Pu�Y>�����[�{J��?*�FqQ���ϹIG��'����xq�9CVQ��`V�]��Q��+��W�����D�U�h��*���w���6�3ZۖU����W'�}��ԧ� ��OH�*�S��p��Qn�z����U^gFz�7�uy����@)vg��<�[]j�ʩj�����W��-�M�^/_Q	D<��/y�}>��z�����*W_;~[1�f��Q�~��³�p� ��<���F*
�,8KGِ���5�z�ǍP�1��}3��z˗W��Aeu$}��������{$gޖj=<��L�ٴdd��.sӾ�N+1�U��^Ru{�B�~n��z�ߎmp+#޽ ;�e�O*�)9,.70X򊭤\x�*0Utdf{M�a�*��8sf��:X廷kH���
��C1�<�lm��x@���k�8��dJ�z02�$�n����(V$h.:W>6����M.�AvԤ�wijIW�;.VJ*K���i:�o��"T�����ۍT�L��ܲͣ}�O5�y�Q,��~���F�?��4߅G��]��q�Iq>���tI�|J9˒�`]�:��ǺZ4z�jX�c�=Q+L����b2��Bv*5����)�s��s0����5>�7w���È{� lL�?p�r�sZ�w���j5΃4���c�'�;���m�(��GҖor�����^k=Z��^r�x���Zد�����%��� uw�Y?�1x���&sGy��U�=�TR��TGW��b�����GzO������y�M�'�������߉�+N����9�e�s� ;}~�����PY�Llw{�>�GJK��K�ڿ��ڄu|�0�܋u�Ή{���*�:<zz���W���{g���;���q^�ǡd��I����	�DL��O�{�k�{�
�kK�ɝ���HNW�=걸߯��g���Y�5����_k�b�{%�N]�b���G�i�u�\�=uL=����K��FԠ�y݇�i�x���^G�;'}����T���F��T�[�>��W��>#��2�	?"��D��G�o�Ss~{u�ב�縺���'��1�n���Xq�ԝ����ǅ���Iܜ5���!�Rh��>��yɷxJק�����Z��lQ�uT��%��u�n�W�CMרz�[�wjXQ���	��1U��|f�U�jZ�lҫ�|��7_Y�F[���U��Y��e)��hM����#k�����0y���`d�C�qw�9��	�;�5LSt��¼^�w;�{"%7��uZ��&ϣ��p��"�z'û�D`����VJ�ˀ��'@nn+�@�_����a�Ô��]���Z>����F�x��\:��q�J)��D误��E�Uz��@o����ط�k˸j���ЕP�Ҽs ��]O�����/#ԯ�n<_��I��=�r3�X�yQ�}���øɟ)8IN�鉆�Ց4�tdJӹ�7�adO�_�3�NS���6�u����Y�敎h�JQ<O�O�ۉ���^&&���q�}ǲ�6�s�'��n^GF�Tfg���o���->�����x��"�^������}q��a_���:�W%�kg;0�4e�A���ބ��,c�<=�E���@yd9۱��MP�Q˙q�`�_�A��O���O:vu���i��s~�>.|��ڄ�|�e�g'v|YN�x����%��=�xڙai; kk���:�����ޡ��
�'kf���q�,
�W�d{լ�r!q��g\R�n!�T�Em�AX�&+�k�ꮬ�	���e�������z��EQ����f�i��k{����F�.hN�ͫEUQw#�C�5Y���DS�y�V�$v���س#����i��<[b#��M�U.�Y�m����\�[sm�αǎ͆�1H䫛Ul�j�0�y$�/�&l�ztm��!��Z^	Ì�����bO<��,^������׬��5����~��q�Va�Ix|�����kK�;�{N�אײ��>�#�+����e�Pv=����V/.���ԧF��m�eJ1vqQXQ�ƾ�t���:ϧj�1�\��uK�	���Ą�AV�����R�q��x�������	C�2D���S�5	����/=����f�ܕ�+6�=~�;��q�9/���}^ӑ��[�-իc ��g����<zv��b~����oFn5�� 1*�}��?i����~�z�6����v;��%�|:!NQeַ�ML�]�f�yM*JP`9>���J�QS�M�Kgq��*�]߭�ARg=�F�E�w:�d\I��>�&�GeFw�|k�L4�qdBD��zNA<͋���m.�(gC��xR\͙���~�fO����~������5
�|U����Qt��}>ðKGw!c׌�Gs~[^s5uG�QW��<SL��`���@w��2$U��D�G�&@|o��}O���;����y��	L��E;N�/h&/i4r�����������?<As%�:���oc��lkx���޷�4vb��¹6#���§C��.8��Q�K뱷Ճ�oX�Ӵi|����z�8\��]��T
��楋�U��O�Z&;�K��yMx�9�Q� �?a�)�Q$�,�~��E.�`o����	�F����;'�{O��BS�)И���6}� {���]ǘɒ|ωY�.|������� �xG�OM�6p>����cL�.��i�\yz��/9<j=�w�zg�Da�T`�����/�OG���i�?�۝�����_�:+M���^��J��ᐽZ��+f� ��}WT�E���oc�͜���mΊ3�#���=�"���I��.����C��^=�Zl�**�L�����'��>�X7��HH�|kE��N�/�����׵��&���@��������,�s�׏�ɿ��x�o�ւ�������H\fIGo�0��=���Wy���^Z]���g��nr|�O;�܆�~㑾���b�q�o�^ל7�:�͐%v ��x�Q��R�gNr������&p^���W���J��K~���~���_���U��S�t�{���]$\֋ټھ�6\�z@(�z@�uL
<�'~�A�on�z��hy�p/���q��ۖ�;F,]�,S�L=�s*�iu�+���S���g��oV�H�++��d�p
��8Iݍ��3������%dҳ8؂�9�.�)ϡ�j���k�]�I�@i�Ld��HEp�Ū���ͪT+��3�W)B�gڏ����d�>1�%Ѩ= r��Q�%����+�w>}D*y��,�8�7�k�3d59V��AY]ǵH�W������ �栞�U*1_�Xr	h�8&z}c�6��Tל8K��oйc�H��<
����__�܁q��ðG������SC=�bcۏr&쉽�K����4�w}c�5�%qW�k='"��.=6 }���e�Iؙa��Vo�5�n���Ï��Q�9t�:{x�Q/C~���W�q�I�[@+~ےqx�	�<�=�y�S��i4|f=�nn�:�3�G�.V��wǗcW��\u����y��t��Y�'Ӿ1��wՋԕ�1���&��^�u\en�y>&�΃4����ud�-���#�H}yݑ�nB]��;��m�=/�4=��EG����_���^����k�o���3u�zˢ��=�.�� W���s%�>����ۘ,c�8+���9be��;A�g�A�����e��"v�p[{x���(4vok�ԩ��zu�r<�u�Pߓ�Z��6&X�����3o���C�fRw �j��d9���û����ބj����ÂSy���'\��h�L�o2��OxY�+��|����{S�y[Í�ަ����q9]@��[<�׹�>�) ���X�T�Yl_]$9�fv!��,N�j���Î���Z?]��R�(t�HW:7PoD�S��t�=��1j�[�[hJ��+9�=�MS�vC�-�Aa�����j����u'۠U�������*���?��Z5J�Rڊ��N���2����݃8�u�-���Ke�iWe�9�����)PL(!�,��e[��/�|-�1](ZU<���������@㬖��E a�Ut:+ףc�X��j����aV�+mqX�S��d�΍"g�k�l����/����m�,ZBf��v�/����6��ft�՚["ws�u���C{wz�<1_����v��K��<�}\�7 �,���"T�4�X*#ݛb�.�Z!E��tN�˝�}h��[�}t��V*�<Ȥc���zr�ڀ#��Lpt�]�Z-L|��C*n��.�q6��@�r�d�;z��u�4���yX�۰��nm�o:	F�
ݔ����Z�XG՜��OaV���.k~Z�b�r���Ynܖ��v
��s���n鳝Ԛ灦emur���A��Nt��i�I��s][���em����Σr����ΰ�����iW\t4��������]��;j�X��q��E�.�V�3������X�pޖ��n�ٜ٨{E"��uwan����1�5X�I`�c;{I$�	N�rx��[��V���4c�d�]Չv�W��.pIյy�$�\��^�}�=��#|e�F�lE���/v7��c%^�Z�oQ�C7��JP<��wo
3sH*���jTyu����K�
�ZŬƛU[jPU�KGTd��X���J���[�g�JCDa�Η
Hm�X긩��{{�(����7�<�6�ɑݠ&�KeJ�܅��f���4��+�_X�v���f�`&����ӫk㕊R�܎��
�o�CRRXe%���ι��iB37�"鬎�J���8�cQ����� ۺ�/�ȵ��t��R��/_-����U*���\�-��J�qgh��%�/8n�(�XNQ�W�S�1�.<z��]������.�xk�u����K����o)	A䬙���k�=	��s&ˑ�c6(b��T��V�2�Wʙ��s�m;0�`:�in�^�r�>��;��!����6��q:��S��.�8�A�4xh١�f��)oJ����H���j�����#)E�7�*t���}�I7�1�J�gX=J�)�Z�ZK�si⺜j<vK딠�[��'N(;f��eh��X6��
��Ȣ�E � �Y=CAU��V

�La1�2Q��eH"�Aar�ċUq��i2�KK �E�XV��UE��1��Y���$P���E�X�T,k(²�32"V"J$
 �Ur�a���eJ�b��X�j(�b+Y*
��*Q�LU���k-�k)�1#���ELCB��h�A`ґB��-�[Im�.Y��Z�LVLdb[J�(Ȱ��[DjTb-Lq.fl�amYW(T.R��Q����XV��ƭ�3��LaY�)�+m�X6˙�cV,Tm�m���PR�2�eB�e`���H���&eTe`�"J�ejhʀ*����X�d�iX��E�������T�qaP���,�E���E"��b�$���]*�Φ�5qnE��]b�1�A5�֤�����Ctm��ӵ:�ow�l	\��V�O�$}���id���Aʭy+ҭwE>���p��uƯ_��j�e'ꄏ.�����%c�-���a��U¼D����۪aa�>ܙ�L\렜��=걸߯��z���'x��|n2E*Ks3Ϯ˙���t֡u�G-���H�W�L	��/&u�q_e�yꃽ3�tv��3�Zzr����>^�v��<V�{�yI�Q�3ƢO�SuL	��|M��2���?2)�*�^B���'<PG�`�C�/�g�^�p��3ⰻ��!���w�&�����ײ�p�_��3���e��Q���\���"r��q��>�Y+޿_��,��7 p�u��.�χ���Q�<�#}��A���'�}��
.��)ïZE��y����W�w"ߪ�E��EG�u:�~��3���T�)��*|�`,-9�.��~��+��ߋ���Q��>.cˎ9�L�oq��>�<��<M�h��L'_E�&i�x��>��P,gC~�D���c����-��%�{Y7Q�{�[3�N��{r&���OD����}�^&&)��7�ù	c/w'<�{��gѶt�o#�ҹ�ɜ�®��K���:��f�u�4"EWU����LJw1��gk�'�L�<ByB�.�f�N��]*���q}�-:M#]f�8��F���7�\i��o˵�
RN��s7P��4�k�k���s�V���7r"9ƞ�g�	��j�˫�9Ys�����-^�hz<�_�l�c�vM���W �^������}q��a^z�H��{�>qge���s��=;](`�{�k���T|n!��X�nǆC�4E/D�p�;��g��vL)��W,��?F�w��&oj�|�e�dB�QjNyT5���G�\��IG/�˕U������ ��N�`�>��c/�U���N���c�3yR�Vr�ǳ�N2ɿ��4���늤Xy�o�i<7���g\�cl���ζk6�2�kJ���:��M�`ns��m���VK]�g��8|�����QOr����>��T�Td֖.2g|n6��!�e�����7��ʽӕ>�M/^=䩳�s�{�\G{nQ����/	늨~5��'Y�{�$�ӗF��g��;��s���޷�>�:�=�P�����D��6D����)��`oT�AY7UZ;�8ZEo�}��>��~%���u�>�I}=��/�J�/ⲥ��eh�t�pU�{՝/=�.����n2W���bQ�o��؏���G�O�q�t�>��x/n���u3Q=��&;�6��ҥ��jI��ۜ-�=P�B��O6�`M��(d4L��Q��?f=薅؍/;��Qh�\YW�dE#����\o%hV}6Zbewvr*UއQ22�I���ɷ:Rx��v�S�q����A��q�[�G.�WQ��gf��x/���#���t(�h���<ζ�Cqڭ��ً�>������^�Y+Z;\��=]H׋9Օ�Ҥ�Y��w�LL7Qt��į������]1[5?w���^���<�]�c��3���I��ndLW�S��B�}t�O��9�Z;���>>�^�� �ΌQ�W�[��a}>urn<����X��%�W�[:k2��o���xQ_�׏�jGq:��)��� ��,w����+������@{�� +��6E<�J&�g�m���j�k�Y�.�g�ȴ<B�G�-V���>���.!;q�{'|��Q�n�=p�;tJ��>Ԫ�=Y3�OH}�q�9�(j77>
�ͭ��0̥�Ǯ���/U1~�S���U+��쭑2�P���/B��T��?2�������d�a�8v����L	����{i�Y�{��R}�vN{A�7e�{*�\{�኎��>�}�厽r��>��3�����#!>�Φ�w���k�=�M�u���,�(\k�Z-`��q%��Ȫ�������q'S���'o�v���Gl�%������:�+x.��vM��*>��@-Vꩃ�f�[����ߚ'���W�47�y�3P�i��I{�S�ۧ�nI&���mgm���{����:�MKy�5������[�(J�(cΏ�#���J��al?W���d�����'�1��f	Cne�=*���J�G�g�.�|������;�d��n''�3���5�W�����_W�3O/k�ymVnfɾv�׋�j ������rg��_;�\d�sᏮ��^�_i�[�G��\k��*���]�g1�w<sH�z.��z�*�d	F�v@�U0&����J���R=q��C،����9���9뙮�˻ڊ� ��h�e�G���U���T��=��9\Uz�A-�M�^/_Q
�f�>Q7���n�*�ԝ�ʔ��������xSElt�����Y�y�!���x72���Xi��T�%�C��-�}y��Gz��i�ԑ��P-Ǻ��~�R7ޯ�� �9��d��/�2t<t1>��\���;��5��n��z�ߎmp+!{��mNyT�I�
m��	�q��'+�BQ���V���S�w>����f9{��n�x�N|�hV�3���0�3jI���r�I����w5(o��Q�V��wǳ�e�N�FlCu�sN�
����Fߐ��.� ̊[pUn��W4�f�Rk�w���������3�av���.�v̮s�#k{-�y(Z\�ɯ$������N�c�X�']�$X��+���f0oT����vZo-��m���r[�{�c]x�����/����,�9�'ݶZ��=�%?�T��2N'>���#�u\en�y>'Y�gW[��c:�{�"�y#�K�K	�ꄈ�>^ڱ�h�+�^r�g�~XЯO���h�;j�ޕ7%ތ�^w:���������^�-I�7��˱B�{Mh���8KG6v����ޓ��03y�z]ލ��7����Fu�X�x��\�Rr��xgY'NΏgC������WUH�msU��&Ϣvxe�mü�+��>}7�S�ڽ^%}�g�ި�+��L{c�r�ZO�ˋVE�/�p��#t�6mW��ɭ.�g}1�΅9]顶߯�����y���ޘ�y>���9��W�ϣ�U��%e��s���0&�X�u�g*x7��>��+��Qp�D�w��A�i��JG}��.iTc�T��=��jO�SuL	����8/<�7��2U�z�\=��<���$gW�z3�Z;�uxr�V[F�:�9���PĨ��V��S��^�]��p�{	�C+��!��F�y��3�l�{���g��#E{���
�Yh��=�^�}�Q�Kʧ�`V��=ݴ��J�=8�2��h�&�RT���E�����6�V��Ef�ưr;�Z�/�V� ��Ch�2i�qu켠%��$�X���/��l�΋��CL+X�b
J�򩂩Ruq�Aw�]Pwq~�}��H���h'Q���ko�I>���=ً���2=*`�KGې��O����~�ΟO"�����쑔�m>���*�*��@�I��&b-U
�.|�`,-9�������(����>��Q�˄*a�5xO��v%�J�|Y�|�\��UJJ'>�>G�^ۤLӞ�џl���X���Z|z�~�W�{V$��o�)�}��צw�:�;���7[:ja��x������q�ú3/��A�Of������*�t\su~9�:S��p_�\��e�3�v��^V鄮2o;
���ddŜ���C��WU��cd:�P�TY��PY�5]�<7���!�(������B"��o��w�%�59������Q�ͧ���f���~7�_���g��+��޺��3fb����Ybkn;XU��Uy�f�d�tfD��e�z�z�'kf����&���=�zq�M��3���� M�ua..}��lո�?mΛ�,��*����ʴ���_��>�!�����7;��2~�|O�2�t�)!�Z�;K�t��>���[��-`��C��2Ũɭ,^L��Ӡ5�L��鹎y������	w�x�j�Xt�$����dw�A��JT��u�J�0�V��Jy�j�r�]^���\��H��ҳ�'ue�]�F�9�m볨�i>O��7N�}��Ԡ0Y��n��H��T�	��W+w0^Wt*�į��/��x���}�S��:C{��(��	Hܗ���C��t���wUJ~iU��o���x��B�����z�nC�_��Ѿu�{}��]����(rؙF�����I�6�g��6v�B�-�d����~ꇡ����=����JX�g����X-�3�;]�gOu)��{�(SqE4���L����K2��==��d���}>�NR=K'�ګuߤ+�ͦ���W�Pe\���+�]
.Z&�X�;���Op�o�ً�Ϥ���Oyl�\���4w��?I�_E��p�<r�%��g�H���F�_� .W�0>���;�N�����~���zϟ[��~��7�>�E���'J{u=r棠>:�baz��11O��r�Y������5�Xu��ϕ^��Hz�~���U~8}��Y�^���q#m׍�re������W[��qY>��[Z�}�=�r����&=��?C<�_�G���¤ U�a�ze�����3]ㅰѡ���6H}~��Z}��m)|n>N�F���f�Ǽ���_��Kߟ�Y��D�l�F�1� w�Jź@�8X����o�Q�z��J;�$���O��f tm�&�
ՋVFu}"7rdC^�)��p������2��s�a9B�G2�բ�P-�y�uc�\Њڴ�q{������pn����'���?_@4��'��ަ8��c�	�d{9�����fq�M��)���c���-�TW�*8j?2��D�3�g��FN���N��z��3Q{l�5���|�O�v��9}�^�=��j���E�}�bm�nt��xOi!���2}ŋ�8w7���Awj6P��*���Z��`U��_��u_�$d{e�o��~>�v�y86	�$;>]�T<3ϴ�����T��]�^�o�=����@�t5~�#_���{g=���� �<����4�Y(�L�����E���Ao��c��A��9�7>�::�3���FL���L��wq�?W����v��g�|ߵ��f3����s	��O{q�P�������툪`M���L�>���W����}ON?K�H�\�\u=�s5�mS�����9Y��HO"��|�����ϊȍ�%�z@�]SjyzM��H6vNw��P��g��k����[�������]��S�7/�����N�4��g�@H�/�+��U:C������ȯ.W�B�����AZuo�����Ҽj ��:���ʪX:��~��~�SM�e���m�8��0��Be��Dp�k~��= ��<K���8�9@�Fv��F��0�B�L�t�l���ծ�0����t:��w%���2Ja��Y|:�q�{�;�:�~���m����hM�6�n�,MN�^f*�e�h�Ǯv�P]�����	h�3��D��)#���^��{�H���У�~���w�#�[�~q�#}Ꙛ��_H��g�l����^Ä��|j���qW��~#�<
^��箈���m>���\�����ԗ��o���TD�9�;���8�^�m��,��Ϥ�� k��>��y���o�ےj-�%�1�tԱ��!���"�������\kOvD�í;>ɸꊇ�5�S���9���*d�^�IZr$����j�K����5�A����R�X`��h{��O�_�����e�dy�=4��ǡ�F���$1y�mB��en�s]�������C�����f��� ���߆B�QjNyQ�]P���kGx�7�-J=�`���x�#�U<if�3����f�i���zs��;��9��(�z�D���"�F�8��	� sw����:�9`?�/ԕM/�kC���jY�(o��Y:�q��n���ō~B���\%N�t��.�W�=��쑸O���T��2kK���L_Ӯ�s�ޫ������jx��8��@�Y�c�m��H���:�d�&�����m�w�c�*�7���/�[��N��au1.����)z�y.*�Ŋ�W�*���!@�˪!%�p�:�ھ���K��*k�2�yJ��i�ǚ7�����-Z��p��ݨx���N3��\C��7�����\�+���8_�L	���c	��_V� ��t�B̦��Yq�������)���|�粽��Z�����be��T�U0&���7����ϋ�7]�_��v�F�^G�>���FD{��=��xu��A�����q.��w�I��ͻL�
�3VW(��=bS��0�n|���<�W�s�^��0LC���s(��S[^�����],�T���s>�X��9��e��p���*��u�H���S9��Sw츹�]�lO�T�h�z@��9*�<�n"`��-U
.|�f�aq����ױ+��T�z�7W��ƞ����?����K!�þ�#�����I6w�&�D�S��ч˰����~4�����$Nؘ��＋͟p�O�ߦ3�9O�9Ꝁ���j�x�M�h���C���11MV��K�{�9ꊭ�ˍ�W�'����P�ﻦ����:9�k��R�b�r�@����"��K�}�\�C�>Q�j�}���}>͏u~��I�+O�����������<�ʡ��!/D�sc�x}Y�=&��V
�"�*�go=;&K���K{G ��'Y�c��Q���nu ���DeE�[9C5����[\�NP�3��e��N�Oo��{�I�㑻q᥉�7�+/�%rqT�Fw
wWt@<oM<]R��ʷ�^f��8"xP�
낖���uw`��O@gT��f\��@j��Q���k�Ut��L�Iv�xj��#�7���qm�qQ�;:���c���J�9������:w�(S6��P+�ݚˡ���.�>ƭ��ۼM�S��q(�5x��*;y-
��~����q�]���:˥$,xCBո��եuC f�j�=~ �/n�άa͡��c3(�[Οj�min�ۤ5U�<;����pܭg�`5��������t��~U��C�/Wi��+m�Ң��r�|�'\1���U�=^�s�1]��-�q�p�W)��ZI^�`�dx�Tٽ����z�J�֖� >���/A�Ύ�`5�na쭮��il.QW�k1��2;nX�XF�#rB��nv`�������'R�qv]�ý�S�CXv���t6��@z��6��s�����쬖��g_n��H�6Ѹ�9�슁g��%ҐV��}/U�v4����C0굘�ys�pI����T\:�@���E��S<X�v��.��k�ɂ�=��+��m� 3nHw��:��Nvڜ��.�e'�V�h�)_R:�eZ��8֕�$�^�9VJ7��Z+m6���7V��W���Ք2Ax9kfje�2R^Ұ�J�v�V���H�M����v޲s���(]�����f�)�rW�i�;O.��d�-���P��로5�ˑ'������ɂ���%��)����`WRj�b�?�iȳ���Z����D�|�q}Ǵ��]�ml��L�6���sb�K��ٔ�):&�\�lpcn��Ö���tVMDx鬼���r������X�eP]Sw��bs��Hu��+��W3 i���s��g:;�2�B�L�\��(N�0/�����>jtf�H�t��S(ݡ��psJ�3����!���v�dM���N ��G%��%�+c	�]�#|�b[�[�ov�ogݯ���0���m�(��n�-n�� �)�Z�s��vЂ����h�7Q�2FU���m3D՗n����g�ѹO��LЌ��ʱ���Kc��9�W�2ga���:��bciy�҉k*Z5Nx7X"�ɘ�+���")x�v�[���սr�akVk�]09�^���,PƧdy'-X�Z�p����>
�h԰���K�f�e���[=���;eIW�h4��o��\�� �dȸr{'��z��Z�1Y��pP�t��S�x���7مէS�p��d��:k[�f�otTd�d�h�u3���RyZ�?J�Oz��c&p�C�77�C��$�j�%����6 �g�����pV�w����z�u�ʭΧ�A�:�Z�j_��צ����>�/����*,����i��*\�R��\J�em��`��P�,�m�HQ�b�-�RڱkR� �D�"��(��D�X����Irb��R,�mb��m�X[c�acm�+U���++��UE��U0AJ�"V�h��Ķ,Z�P��ZT�X(TP�1
�dKIF,P��D#h�kR�RUd��(ȥb�`�kX�D[[f2LI��d+RZY��-e��-)Prܵ�h��0�b�"�ŬeB��"�*,T�¢�Qd�%E
�eH�AAk*-�������YYZ��VرF�6�Z2,
2���PR�EX,�jb�
E��k�P[h�b%jԬT�K`TR,Y��\TX�[E�D%�JUZ��j�P�j�Y*h�PYPQ��+
ն�ZȴID�
[DF�,)j1Z�PUR��Ym���+����)
E����h����I��'N�EV��B!�h[�5^E���Vj%u�_u>�3{�1Y�R�%b{Ŵ7�x��&��R,�Y�������ؾ]N����o�Rok�=���3_^�?������������y�s"�S�%�eǩ�t�#�=��:r�x=7;,e�p:����{f{:X������YD��N\��S�}��I�әa��֦���C��3���xLvs�u�U���3�t}��Zn5��Nq`o��bfi�('�弗����������<���϶���	�$;>]T�a�,o�3�<�������{�::79Mg�<���u�.=���k����e���FقR$;'��~9"�_y�����ڷz�̽��h��>U�q^QN�k�Sҷμ�o�������BP��$OJ����_=��f�t�m�OGd�j4	�W�%x��P�K�T?}���9��[����uj�<7}4k>��4\��<S��d����@�QxSqE�1M߁��˿�ՉE��q-z�>�|V��?T�1T@�ι���/�6�+2��f�H�� 2�+�<���!S�|(����3���]�Ω�ʢ�u{Y�D6/q8z"�n���9^�����qt���U�.W�p�W�CK�*g�H!���[�#������WZ0^*݇�rڔ����"�ޠXΎ�	�/��i�>�r���A+��)K��h����v|���a�(�5�'^
��2��������u3&�=S"����ޡ��I9��;8�H����ݠ��t�ձ�0�OM+��m�<�zE���ئ��,?t����$y�n�`lC�j�o��t�����5�{#3�z^X�N������#^���l��z�_�A��d{נ;��D��^6�ɖ�Lf�
	�_�uQy�����>\�hޗ�ݐ�Cҟ��~�Fϝ��l ���#�v��G�
�+b��mu.5�h�L��fl1��C�N���|}e�:	�?Y�{΀�+Vʡ!��$&�*�Z�%��{��ڒj<���.7r¼���6�'KfvK��2=�Bhi�3yO��}#��w��Ǔu<}�۸��\���/
�>gnv�?^N���N��z��3�f��>�2o_��������dxg�q�<���U��{nt��xOi���v�j_�^�Ä'
I���:LpVj���ݼk3�G�ԁ�Τ}���H�{i�|����P_F�5��`��C��۾���ǜd��;k;�=��YQ�ή���5~�5ϯ��{�|Wzt?uք{M!��y�/����d�U�ٓ~�C��aWخ��N�M�e���o��9����o������+���,PQ�:��.��:A'ת���D[��diWI��i�_����@�W��8y�]v���kkD�-�9��ل��9w�=��E�D�F��*�ں�a��(�}��wt�S�̛9;(/4.���rl�}/�d�A�D���f��f���,ͮč׬y-���%W�|=qT���\;ݪN|6#�_��z�=	״�}��j�ݩ��ΉQk�R��Gp�!�R7)Tmǖܲ�6@�jz@�\ESb����A���H�Ꮂ;���ǻ+K�ow���������я���{��6��q�*Y��q.��9\W��A-�L��A��g<���ʚ��˖H��z�C>��1g}�{~~�6�^�`k3bF�%��S��˕%����'�W�~�AU�>�}pUD<��>���{��=�F������>��y��愳���[Q�\<��� 6k�SB���a�Z;��C����qn=J�G��)��;�|�c$�V�z���9�9V��> U�NI���q����"i�i܈��S/M�߅G[��Oi������G�ݱ鬘E���j9'�$��ܓQn|T�a��7Lu稇_\�2+^ׇ X�aa.��:n���z���G���&�"zS,y��Q9������50��m�x|:Ihc����1]�fG���+q��P3��|=p�VO��Pw΁鸅�σ� �� %a!�͝�^�R��D�xF_�li*�.Sz�v�X2S����\�yUڮU���m{Vv8��b�հ�� ���N�-�wu��$ �Q����nq}�4#J�s��6���RvJZ5t���cri������7*[)�9��p� P�&wX�c���uq���zm�-�l�}��|{���� %^�}ꏔ��7r�uB�����Iӏ)�P���N�N����&��>���6�N�x��u�}������YG<��g]	~��q&�y[�Iz=�'N�������V�,>U=X鿝*���z�M{'|�<�R4�U��y�_呖��?V���yQ��o4δp��K���T�έ<>�ig鋉�A9Ȟ�X�̵�7J�FK��>(��f}`��]\��{'x߽���l���H�lUL	��0�~�<}��9��آ�=w�)��y���]��z���9�;������q��P�[(ԟqSuL�9��7
�op�O[��{��ڊ'�R>�{w�ב���V���{�����c �.��!��zF�a�au�YϽ:���[蚍�Y6�ŵ�y��C>��/!^	t��������ݢz��A��l{Z�6},�騂x���B��H�h�vcx��֑�~��e{#0�o��15��ֺ�ǘ][R<�S��鸘,;S#>�����Ӌ���kw��-�7#OI�(����O�+�P��y��)�g�k��"�/ei�D7��J�ƪ	|������mIC�Ϋ���j�=k�U/�\��W,Wo.�t�k������ �@n^�bqn���a���_��GV��μ)eS�>���K)�N�=��ne�D�Ih�����]"f)�x���Zu����;F��Z��<�����ԅnz�1nr���N���r&�׉D��͉���^&&��'�uY�o�W-���;��k�S�'��>t<�>u8�<r�K�4����;��+A��������Gw��tǱOI��>���p��ׂ������@���9v<1N�!>���g`�mf�{�C|d�9�7l͏3���}�q|L�E����/�>^�,��Pt��>�O�T�WL
����9ޅ�r��zJ8K	���ޜ�/*�ޖ=�9Ł٫=��-ߓ��;蜟y��N�'��#�}��y�ΛG����Jq;Le�d֕q��Zn5��KN��ᏽ�5��;�P�k���G���ޝ���l��`��C���Led֖+�78t'�O��֑��@k���C�y�.5�2�-�����TQ��������d�z	�r�b)����0~���Y�fo����/a�vc������3��:�CF{�)O����(�\8�W@��/����h^Ֆ|st�^���0��0E�����w30�6��by�_R�yZ�?L�]�"�iT��?f�G[tbi�ΨSyWԇ-���:�d!o:�y�F���F��3��ڟ+{K��v�Q/���6�n��L��jc�]��w;��΅ү��������@Ms���Je�Ϯ����9^�iϼS/�}~N�u�|��;��T�Y��
��5��
@�Fts!��Sw�o%2��bQ���=���>C�v9^��dW����%�{ŝ����:�_�B���ρ�G�W^��D��,y�}$'GE�yP���TU\Uծ�-�O��{�Zg|Fw��C�r��Y��w�֮�|J�Xk���<��������,�N�G*c��v�_ު�P��Qr��F��ۙ+���`-��&�G}E{����������NF���{~�|=^�$|=*k�t����#ư~wS�@��s���!�\��M���2��bb~�մn>���&O¸[��ȃ�@{�� +��r��A,{nk�Y�d�U�|E�L�>��[flxu�m�/ղkK��+T�)Иڎ~�f�
�GM�^����$w�$}��2=��q6ϋ�'Ñ�af�ѓ�3Q���+��aq��G��"�jr����̪U^��z���s����m�{�8o����G�R����O�!^ �fL^X3,��AI�1i_��`d�2W���F��$�,ދ=X�I�ZDĸs���f꼎��k[Ô)J5T�/����Z/�ɥ�����F�炇k�&��\�x3��o�lt�B���B�Z|�X�x�t˝Qߎ^r.a���K�/��1X�K�i\����v�+�=����N;@�yQf�}�b_��oxOi!�Oח����S���Mø��e����Ǉ�JkM���u�
�Uo�F{�M��Z:��Сk�Z/�wN�C2-�d�w�����'�n�˷��*�=������ag��~'ϧ<{��:���������{}~vkZ�Q�}ì�8N�;>�����Wp�7j��x|'�Tf�^�q����=�ve��vF����R��ў���]��g��Ei���=U0/�P�&S��/�įU�W��qz�A��M��T*�{��ܦR;�PF�*��i\���Q���U0&*yzM���g��P:e�,�J��8K�zFz)z��p\=���}�C��Ǩ),��tF�9L�K���s��=�k�<��'��>��BP���y��w�W����_�<2
�M��Cr�`�{���[�u�4��a�EVъ��^ÐKGُ�
�oq�c>u�l�(~�FU=:!�)�l�C-�r+�.V^�2z}���@l�Z��}^ß���F�����R�W[�ȃ�j��^R/��s%�ls�F�I��f�l��)M�9%c#x,��@%.�dp�v:DP������V�sA��r��n��5����	��ӑ��9��j4���<D0ӽ$���wsf��x�K�2"L������
�F�ۈ��B�v��6�������ol��*�������,zԑ����wN)����Q�I�RAצ�ow*gzogx{c'�K'8ԟBR�����>%���4v�鎸�Q�.V����Y� 9�d�����Y�yX�ۈ�L�Ǽ�{�:�b�Iϗ��V���z�����Kp��uǺ6�q�'���:O�ߩ7H4������#7·)����M�TA�������z*p�=��^�Z�����z/vw?f���<�E�BW���^�-I��:���˱A{���g_+�7އ������G����wzv��oTz�#6�M������=lp�����<u�n�A�������@��j�3=�t�SV��ͭ�d�;s(c7�챙;P�3Ԭ�i`o������Q�|5�]7m��?].k|�����޸H�y⸫�ݶx��$��r��C�gK�s��s��;��N�tG�y�敪��<���Ѿ����f�!{��=���6)�8\U0&�X�?z���_P���6*����ۮȞ��x6|Ό~u�{~�W��V�7>��ύvQ<v��Ǖn�g~K�%�0e����[n�PzMc�[�V7�SN�x_/�>8�}0}@ãRڙ8_j�O
��2T������3nE̓0����O/uw
w����;G�' 8�%-�L�u���G4����:���m#rR�ۃ�~��2p���󜍩��.�Ō�~��%��t��O=aw����9d^׫-q3{⧫B����|K;��&��q�x�������ϩ��G�O�v{����k9d�����w�˯U������J�ʰG��:sq���}���f���^��gE�y�uxf�;{�<Q�}���\.߯G����r`0��P�����ә���(�{'���R(��N�xU\>�~9�q(���.��r*�S���-���^�VD�N{�B�U�m�Ļ�7c�{�6-{��z8φ�o���&Uzb�=O�9���\Nۯ����ۉ���k����ns��o%�!�1��������FX�������y��Ju8��.A�4�����{=
=vk�{�hw'�uw[��z�Mi��U���pn��w���Y��<�uC�b-yʺ�8�vo:K#ќ$�˙���l����ͯq�/���ۇ�7�~/UQ�m���=}954�h��<>�g˲�=�qʜ7�$xܤ�;�����c��ީ�~:����ўl̸�[�:/z�A�oz�%[f�����]d�-�r�FE���Kz�|�w ����+0�e)�~P���Dz��G��Y�����WX�z��1G�;�`WX9��b%��.��C1��㐬G��
9S/�{:�.���Z2ҫ��9��z��j�w�}^tx��bv�Λ�|Oi>(fU,~i`�e��S�/E��o�[p-^���q�Q���m�g��N���\kO�"
5��pyܷ}k2t���o}�饰��)�F����ƽ�}���E�]yߞW����\�0��T�g���ʍ���_�������2��u�q��ۻ��
V�������T��s��xu¬�4.V;ҍ1��)�����/��%�}%�����]뇅��/�T=^G�S)]��W���gNr����C��ʭZ^T��C�%�w�h�)��;��wjģnߖG�ϥG{gn��XNǜ�{Y��M��9�鯽V��#�(���#���#�����c���t-��v����4�;��dW�+��SfyI��I�Q~�p�>�׉b�0[;s�]*.7�H0$͸��[<mF˥����ح
�N�x��{�L�s����1�7 5�ў́},z�G���J';Г\H�[���$sHiOq�n�����s��Ny���$�	'��$��@�$��H�X@����$I?�	 BI�$�  �����$I?��!$��@����IO�H�t��!$�$�	'�	 BI� IO��!$��$�	'��$I?�@����IO`IO�1AY&SY{�B- ">_�RY��=�ݐ?���`o�<**TEU)P$"f��)�B��ɥl�M˝$���mU�TU�*wqL���l�5�ɭ`-�8;��T�� ��l�2Ց���áv�Z�Xm��eH��m��մ�����
r�]�@� h��$@�k���i:�lض�SmJ��Ͳ˚��Q��61hhT�8:Y�e��ѳm��f��;��&�Ъٵ�M�� $�f���k`"Xl�    M�CJR����4 d�db4i�S�0��*�     a�&d`bba0�!�&�O��T&��ɣL#L��0	����L&i��MD��ѦD���G����56ԟ������c?�5�߱	H}�BC��J!1	 �			��ET�$,��?�����?�G�`8���`L�	Hp'�Q	Hza.��0������>�|��rb?��}?g��� BC�N}VU�{��N�Ϲ��!��(�o�;������ز�m�"���}N�1CFJv^f���6�j�:7#�xsj,X؛�)l˻<��S��(��{B��.��m�y�N%��p�հ�e�3F-��Ϣ3-�v�MaYŭ�*(Ņ��-�N�/��M�xb����*w���t�2���X@v��&��EƳH��ǎm�Q7r�,��y���3ͦKf'q� ��w�mU˖<sC�[5�!I�7m���FYi��m�_�.Z�]�)�8�xnF�T��$�m�b� �y`+.��e�&�ۭ�W�j�HF'l�B�J��P�2ӴD�v�z��Fc.t�$;ݙt>4P.-�k�7R���mh͛��9�C�b8���&��a-����,m���!��º����Ҭg5`h��>ttj�X�ך$A�Z=�]Zu�D�8U:��O\#nBt�(����me��݊�*I�3f��YJ��E�¡[���P��mu5Z���A���U�3h�3�$�\`�Z�#LGsb4�m*n�ݖ��a�ϖ�������Zn����nvd!���mCة�`� ��0�kE�P�m�y��2��{sEL5��ۃ&�(C�N-���l���w6���{�Zܒ�#3o(伧u�k�����R�K$�bd�	��&"� �F����EGwYB$�2��pIP�{��0Sp�HY��{�/��{"����t��L7&�{^ٵ32u%n��Pub�^�5���j�U��ӣ�{���a�Ib2B���^��Lf�7{�#h[ӌ�IQ��+�D��CZ4�ѥI��2��eU�t�͆��h�q�����:��5�Xn���֎�p��]ǃHPb�Lo4X/,����ۡ���,��ʴZ��M²���nXl�	���U7�Fcw1�`�6�ЫɕraB��=yY����.�8���Z��� V��P��7En�1-�!���f]��ܫ�j�B��9R�����4�����s:��4���`��<E"p��/]$j�+`�op�t�$�BV1kʧ�JXj�)��jkHk*JZ Ka�i�j1��z��!
�L���N���AT�Z��A�j���S��#�\��ele�qm�^l�h=:2��6�O��J-�U��ziB��kSmI֪�
�m���h��JR۱������5^䗴%�1lY)�n��p֨��ي�Yɔ�8�;�E�k�FQl��4Y��LCZԂ��2�7e(	JDJh4����Z�mi����_�?#�>�?��&��G�{�H���z>����<85�:Wy���{�ۊ��(��6��\�+��z�	ɏO�ƺ3&B�Hͻx�mk�k�Y��P����8��+4>E��9�/K�>ܟP�]����o���Ĥ3��+�Sō_�g>7�/���\7�W��<7��J�{��fu:6�s��$g �$�Ә��Z�Z=�?\BC�H�z[�z'I<��/iR�n����R��I���g�,�D�e�Kt���2��@{�5h���GC/�*u��a]�P�@�ɑe�qѽ�869e��+s0ճ��1�i��h���uh��y.���7F�zc��K�#o��%�֬���s�ԭ�{t�'[Qq���������7�d˄Z�_6����)Qwr��.�pC<4ʖ��+^cp�59c�n�.��s+��RP,�l�@�ݒ{,����n�\���-uL��u_�S*�<�O�9Q�>�r��7�\��ܸ�#��-�����1�"�V�x� �7[��լ3�\��Q�Y��iԧ`�g)��vI� ��UsF���wkA�I�X� ��[�B�F�х6����O`U(iCi)���+�-�^�w�6E4�q�������=6��D�VXWk��õ7�	Q}iݺo/s�s�sq�{ǗУ������ޫ���־��;"Z�aծ��-׊k�ܮ�ؑ\"W�J��`w0,�t�޺t�i=Y��T�g&�܆1F�omq+
Lr��zoo�Ŷ�G��;���?{8���Ԉ��]�c�.{����\��x.�h���"潨j����~�W�M���k��*�����:�9Ε����UgR�[�������Zj���l�Y��K;~�|5=�p`9Q�u�&�"�;�*��C52�`Ǳl�:��,Ϟ�Q-D�{>ذ!��Y7P�##MR�M�J��T�]�4���o�kwX�:�]��O�����������x�kH㼫��N�"��hp�
���T�L3�:�wk���^���[J��[�kf�Z��L�PM�_t�6�h�qNٜ*�*��N�ڷ�i��ջ1��"w��@��L*�N����G+���ѽ.8�m���K�Bg-' �}���xz���|.��[��h>pu��g<"��-"��)�w@ʨ�f�8%gÏ\�x�2��_�2��$$�LSW�S��tI�����e6i���׉�������(t	1gI���ko�	Z0���"��:���������/%��x���ȫ���1"A=����$ِ�ی!���p��q��2�e$�S�Usc���b����>�c��﻿v(���H�y�/ߐ!	!�\�@?D8}�.B'��G��}��?O�w�?Qg�T��7)Kx��O���y�0�Q��@;:�)�����\"V�����W�-kP��5y<M�WSZw}�u� .Gz���K��`* J�qEo|YY�u����I�u�xM�5���T����A;pkOI9�2Us&Q3�:�]�F]��S-��b�u(�f�!0���-�x�3�*·7��J�_��w��{:����C
Uq9":­5�\3$̼����b5r��X%$�����Zv��Y>�@1Xu����]f��e�]��GD���-��.�m3liVI]<<J�66�1Sr��!|B3ge�W�rvy����t��(nB6��Q��X�&��\�0�6Xk9t�^n%|X�m�t3�D
�rD�jjA�4���tn:.���{��u��A�c�Xx����T��}�w�9�ʴ7X@�εP����Z��*����Z�r��z�`4\�
�$�!1�;��F<2#grxzڹN�^��75s��斪kQt&8���%f�Uf��سqHr�J��ݸ�����s&�,m	�UwU*u�2��K-��yT�X�4�gi�hibe)�Kr�Vm�n��ғ���p��Y��Sv�t��cXv�Ij�o�Z�ʇJ%��C
07tթ��S	V�m�ؕ�x
'%>ܛ:��-��x�e*�((2��5�0����,U�[J�KoK6,��d�2?m��[M^��n:���]��(����Z���=��Y2,{�hڵ���Hk�d}hZ�.����)��Ã��ם�)�����nV�ݏ��$�N;5�mp%U�����[�U�B�ك����V~;�.\ ����Y��;9>��Q[�ݥPk�j����<8��in����n�z6�
��
�b�x�+�G�X�/8�5�kYާz(hy�U��z1P����N$�:]i#H���l�y!�\�5]��v];(�it'@�.�Ҭ����j��歶�9JʣZ�*�p��d=k�퐳�R`d����Z�צW9/�7_(��ua�>�;�)��`�}![;RC�T<U�ya��ص�ĺ�!�AΤ�in�ȐEtP�N<ma|���i�B��+oP\3	��4sq�-Шu�=+��ꊗ8JGX�$gnPL�^�w� �Y����:%���� �x���r/��]A��6��P�d�W�*��0-[0��i ucu�YF|_j�}F+�/�-��>�׈��K��*�.�M�9;A}R���Žx ���[�z~q�o���M&�ku������$E�����������b}K�7��� �b��6l��C�R�;����E��e���ġ�S1�o��3X��a��n�4��H��6*�mb�!�!9Yʨ>����&M�-���Ȁ���ҕ���h������^�4;_)^;�S��-��݈=���:Sr�Ħ����w��<Yxp�L��%)���li��.�"�UD�kuX��b�6ղĺh���QTJ���"]5T�ih7JU�H�Wn(.�j���UPJ���TTjU���QB����n���j�ԤZ��ՋUB�u.7TЭ%(���Ș�\~�{ӈ��{K˅-�>W���<E��,��P�}Y��V�t7��i���٬ߖ`
8��+��E�U��z=S3��<��L���gN��N�R#����=�k��5�E��(�K�*a᭩ƣ�m��2��Z�����o�r��ƴ�	���n>��J�/�͝�(��z{��ęබ����
s��1ȡ]�F�}��U�tl��j�7��t�zJ�(��ml+{���]v>{���-/���+�ˢw��B��u-ڬ^�-E����ƈ���q�ة�n�
�G�UR�b�gÙ>�Cz��tWnWzn���ô��뱦�;tB�/}�`ͧEV��m�}L~���9HT�*~�cYLžY�q�@���\���%F-�3�aW�|wY�E�Klo���y��ׯ!�{]L�܈�����,wCu�KZc��<�eby-Jx:�_]�Mc3�ޖ��.������y�U��^\I�S�=��2��u��$t��X��㜶k1%&�̾Dq��̐CƷr�I�՗�~c�S
�L�i^��ת������/��1�j�9W�����՚�J�0�����!�Iw���6�ө\oԳ-n��$�b��Ƽnfʺ�T{�F�aq��'Tk��쮇x���>xUǯB܊��J}w�
Y3 |�z?k�{��-�\#�z ����d��0kS5�����U���\��
em�Q37p���l��4,��ۘ��:��Ty��<��s-�k�]�}�v�؀j%�Zz�C�t�	)dG'�7����(uz��\��Q���!x�Q��o�P�5�[�>&ڹ8���]M9��ji]n!��r�O#�2�:Վ�����Ӱ1�]/<�v*�jϔ�R��.v��Ǒ�7��C�L،�߱����\s<VvN,��&;��J�hzc6����v�td�uү���@ٻV��PD�ft���P��4~O��ߏҩH&��"r��AY���������L���W��qkEe5�Ym���sb�-������\M��n���6�A(�J��m�Fw+�W- n�㽊V@�+Fm�*�)ͪQ�mG2��x������mm��fM�H�m���|3�ߨ;�_P کab�ul�%���(,(��dѸ�C�c8B6b��Ӽ�*�%Jl]��" � [&�P#��5�x�fQ�)<YA�Jth�D���,� [U2��f�b@f)�h�f�n�y$���gO�G�DPF�A  &�����j��r���[���EST� ���E�-R#)�i)EVQV4�1V*���][UbZ]J��TF�KV-4�%�PR[h�[v�Q����z�q�W��&���c��M�W������'�J�M�RϨzm�#g�k�����c>;C�>��?v�N�2��Ԁ�,��d�R�u�#4�w��kF`䡻���(���~��}�^ၛ�u�T�����e�fPfۯ;ca�V9Ft�C��\*�9���8��k���W^&����j���/X�ߪ�i��.==�8��{�wzi�7w�����+=B	,DEʁ�"�����P�����MLQ�2:��bY.,��w�{� yX����nv�F������pX2�(ƅ�F�.^�ɧ$hu������y�n�xyf�4�p-����Y�K�B�#����8߽�T`ְ�_=@2�=0�e,$�I%��ϬBC���Bm�~POL���z`L����޵Y$"�I۠��L2(y� ��c	s>_y��BP6�0�@�!�!ԁ酗����Ǭ�/�M�L׷&�$����ޖ���$�甄��:�����P��5�ַ�Hu�I���IL��I4���!�$�!Ԑ��Ad-���
N g��L�)�!�P��!�Hm������I:�6�m�HCL�m�6��I$�����HW3��$:�@��M06�$�Ix�!�H_=g׬7�!�0��RB��$2��2CĐ�o�/��lL��$��KdRB��$a;���HoX�H_j@�)��a&TL�I�y��Z�F~��W�+�[V	�S�fn��S���2�:���GGoI#����r�X:拏Y�7-
�Cc/e����L���Q�I���]7J Z�ɘ��R��v���C,'�{�tM6�b�t���d���7זw7�<T�ֶp"��>��6��.�=^��M�E���}��u�G_V����:���vi�	 �������`�W�v��f?6\mRي��6��_+��eB����|�u�Yl�9;�4)��;]���w�ج)7;�L-����R˔@����q/�:���-D`��P�=��ӵM���-
� G[�pl�E6ϑ��;i�X�5��JP��ǭ^�O�е�h�ܰ�|#�X$?=��t|�69o��H�>�Ik�3�Ss�㼿�`���\=V�T-��-Ǝ�1���V��
/���;��L\q�l���pb�������O����A�o�U����YTk��{4���s[�{�ơ��*�bfeB�؉�u�2�OµB�t	��TTo�������jǄ�]�
de 1��r�y���˺4C��[�LJ�*�*TXd7$�]���V�Z�t_=��+	̦�*�k;sEn�;j\8��+
������ی^lAI�Y%]8n�,K!�����-M������V�S\��@�n��wX09F��4B�h,ܘi0㬋2�Iq��3-,j,�
d�t�T��8��uXQ2��� h`1�bbX�b����r� �+X	��<�P4�7����u��o������H��j�"�V�%J1�(�-2��#.�,R�H[Eմ��u%]]�j��7e]��)
iU�TJ�����5UL�`�ŊP�;�ﷱ��K�;m��'�'ef���)z�~�#y|�������Hf�����!_�{�>~"V��w�?_�ŧ�2�,����آ��ګ�̯#)h�Z�;�0F /�ˑe�ی�t�F�:4�Ʋ���m��O��� c҅O9S�)��KʵE樌�V$��.��4]�Ye�J�m�nU���_�PM�?|3�i�ܮ�<�rF^.����������$��ոn����H���RgdL~O ��SԺ�0t����/_�{ޓq�RR��U��[�N���}ݡ`U�(�]�BWss�yx��p#g�J�#��ۻxֺ�fd�����Ԝ�-�Q�[�Q>�֝��*�s��q�#��Q�e�L�4�ix ����`��mL��Bj�g��{��)Y��n�E�u�^����=p�|TQ������V��uY��/��s������g���$�=|����e_�5�o���;���T���{(�ؕ��qq9��:�����)�����74R���ys�.�r��m��}Az���{��Fa��0.�/��k����r/��~�~�_�j��B���U�]���x�u��:��eU�C#�����cy��*OxqR��Wc�^!���%Y��ն����	'��6k�ˊ��~�(w�_\a�`����CQ���ƀ�v��������d��8m#gu�3h��sZɴw2~9,1�Ë~��h��̈́�}�;��!]7mvî6g���t�5G�g��v׺5'���a4o�&�vW*4�+�:9�\m�3�L�X*�����G�d��!��dK�N������O�����m��aT�/gc'���`guҩ|n�@�;nj���9�ՅmH�K8�#��2x�Sr�v5�I_���z=���c�ϗ8}���N� ��c?*��8�^�K�7���M��e#��?r�)�c�Ҋ�����Oޝ���/b�{v��<�z���ʜ�3�C�U���}�=���K�&C�M��{ވ�ƿ>�����jw�/N��U��s����Yş��b�c�{��{�eܶ�Eo�ڲ���@��lk���Wh&X���<Y<'�׳�z�4��I����G|r��|��������F8K�u%���")�dE�]Ư��a�'@��foNX�q���/�:`g<��p\s�+�`�7r��]��Q����q����Fr-#�Q�ۯ�6-� UY��h<�l�=�� ���..�J���[����fe�ESD�3+ǐ�"D�edi�v-F���.ѧ����'i���k�Y Qs ,L˫9��.�B-�]`A�a3ȕ�A�Ɏ:��d.�C!l`7�յ�G(��E�lZK�0��6ڵu)��Ŗ��cP�����L�
h�*�(UԔ��UB��P�*�ա��]�8�s�r4��=������[��+�੩S�F��9ux=��j�44�X:V?lՃ�k��lk>�����a�F��Λ��|�*�����O�{���\Zzi���]jS$���j~���D���驇[�{V2��S��ri� xQ?��+�������啳$0
��S=�+J����wD������ց[�@zH����A�u��#�y��=v�E��T���L+M!b���\"���5�Y�嗪=�N��)�|kݽA9��R�N�f�*���x'}}ھ�tZ`���H�W���-LSC��$ѾE���y�fi�ߢ""!����}���L�sz3��<;�}��U�廲n�'(n,ǔ�Y�}���2eo8��=5����0Q%�oZ>bi8�{k-��e�2%~�y���=S�ճ�b�.�����Z��Vѡ�1Oml�����6�c��fwm؁=�U�*#^��߮V�
?�!J�#���^������K�s\�x�Y�[���n֤��Z�<6M����r�����2�AcF�Fw@�WG5����������z�?��U�Q�1��O��~���O��;�dQV,��y:S�Я<�)�������;xn�f��5�����~\�--=ʞ� �LfD'D�J��9�踏Dz65��}��a����us/iٹ��r���u�:��
g����S��9�m��s���RRd�џ/��[������`�M2[5ti����L0��hӗ�,�2s��ި��K�,:�:g��o��'o�%�t�f���%n��y��G��\.J�:0��A�߫�����F���XfRZN��kk��ש�Q�Rc4R38�pk5*���˄0�_]��˓o*�;sښfuE��M!���,p�Tx�~�iu7�/�M	���TC,)8�ǋ�.3��y��r����1�q^b�))�aļ�x>��i��)����Y�>^Z�̫5[:#:���7�ic\���������0x��'�4�b��Z��0z��<�њf��il�o�9�<�
L	�a�g|�G��Rm��m)��k�ֹ�8m���L%�)��;�3gPΩe'��*�m���9al�Sh�/w#�7��6�e	ħOS.�C��d�@�j�ά봼�9Z�9�Z�0��fI�wu$8�@�՗��ׁ�s�g�c��}]�{�=�ӷ�e4����֊JC���ӌDQ.��s�̤ۖy�2�M2^]�)�	�m��0��B��̛��3,�i/<�|�q�ǈq�wP�.��|޵�!�����v�|��(�u��O�ëk�8�j�C��<�^9u5�)6�)���3��!�����4�����ɻ�4\닳�	wRC��yyMָ�\���k��4��:��."�3j�Ù#G�V[��YW�u]{�n�\������i��X;�����sf��!��o�Y]9����*�WJd��!j�͊<�d�����bu���u씲c�ԝ�+Y�2��q.��i�zuT�J`�pƛjhiV�����n;��|O�R����:�����Er�i�:��\�Ž��.5�[��TiU�����z���Ƈ2��[�˼�=���3G:^�8εU�м%RJ���Ha�)))���\%��M6��"�f����Qڊ���]X�w�i���|^���>���NÝ��=�uG��{ֹ�T�-%�;ʵ��y��]�L��8ƨ2���0:O;G%&�/�Y�(o4xͦ�P;�Νy���2��to��M��2�X40]3)�	�Q�������)�Y֒�n�<W�޷�������&겛f�ldO��.`{��F��(u�[7���ڶu�ѬK�o着�Io=��� �`Si���zL�e�f�9qʅ4�u�¬�jzlf���nt�W��4ɬTj��]�5�3:�L�ͼa���k�y��j����T�Y�
a�n��g�L�(Z�-]k a�QX�6n�yՃ�1�4M3,Y�U��i�_��Hm����`'QS0��h�t��]��<���S��5�m�與�cc鈁>����α��<Cn�R�Q�i��4e8�ٶ�]�.�T�1�Ӗ5�/�.h�g9JN��FY��ì��g�z��u�;��ؘd�Jfq�5��þQZ��ZL=f<�a�5P�g���)F*x��{��,2��r%7,s;�f=��JQ�L�����T$���ʾ���g~�M� ZR��h�^c&�+[��)��(��	��V*�))!��.�s���u�u!����9x�3]�nD��G�i��<��9��I�Q<{��&Ĵ%8f9�/Tq6��}�)�L3Nܸ��|���I�Z���x��7�֦Y)j�a�Te��ߝ�t;FǛF��9sR���C���~}�7�3���!�4��Oi�sZ΃w��ƨ�)-��d/>Śt��3���e>7�V�cꂷE�q/��y|�0�)���y^k��/׏Yi�%2y����/������Q\�wQd����:��y�2�&�����C}�����uKq�\�h���,�W^�󜨱�E7����4F>c�܇y'��5���Y�{���b�f��^�����ߙ�<e��{��\ч��Q�
CL6U�l�Қ�x���:��z���7�,�-<�Bӽ�.^2�\Z0�23�p��N3���I�*K��8�w��WSI�ۆx��,�h�b]Q�b��.�!T/�EZ)�^�v�@�S�'�D-�'!Ӡw��U}Q�4�.��=>7�5g���3���Ci)R�]x�v�uS/���m|K��{��;�) �:�]�w�`�208�'OkF�y8��L����V3{��\����Ha�0r�u2��m�L9sʅ'���l�e�L!�(�u2�w�f��6%��-�V�ܺ;��6b�z��V��f��� �7��=m��LFLF2r�n����r�0Rݳ'(��mr����Mf�2�#�e�o�I��͡����w��iahM6�g�5��g�HS)ѧI��w�v�$�l���fǘ����m�u'DQ*��欻�.D�����AMߕי�M'�T�!��V� ��=��܀�*��ҳi��l�ZlB_O�_|�W_�뿺�.\�ya��l��I�m2�5�1�s�+0�L��q��OZ����,���E0�*��c��*��w@x��tk�a��;��2�e'L���Q�S'�W���»����""�&p�W��a{�H������4�p��-d�{'W#\§�	u�&����5�-���]�����%�=���^\��Ii:i)��+�k�״^�|�/!��S2����
*����E���+o�ҭb�0i\�ו��}Ӯw)�z�[���׈q����).EvR]�Y�����K7�ʇ|p_8�Ѯ��<�Y��G�*\��[8w"i�e��E�
Z�[͚X,7�zu�g38�w����n@��Iq.�%e��(�CSB�{/}���r"�%xSf�7]{���8zS-���;;r�1��hn��{�e�R�6두c
,�qJ��%���D����N�C���f�o����˕� Aڔj�ᜄ��Κ���v�T���V�Gq\�w�����V��Zϊ �|�jF���uee�	��i����)D��k{�+��8ߘ��;��.Ѫ
qUiHS�)��%)�� Ĵ�EX,
e2-%@Sl�Mף��u��7��`ׯ��z3[�~������<���������ꃭ�wm �a��#O5�G&_gL�۾ί�͙�b��Q��i=�˲k=u�ǢWӬRW3���,é�Ad󾷮�&���~�{�#rj�߭�i/��.����jUO
����4i8^?o��eJ^�u��A���:K�y�
�A9
�m&�f�k�\�j��D�%>V���8�� n�Ĉ��N���u�zs��}zFm8��eo���ծ�?)z�����j7��
����;
J?���CU�^��WФ���Ƃ�+���Ι;��ތ�E�"=5+�����6�}��//�rԗZ!���D%�w�۲AɎ�{`M��?mn������v��Vq5*W7K��k�5mb����Cp�{���B%�+9�
�T4�.������q1Y	-`��45�F�yA��G����艱w�f}��n���3��Vuq���;�L\��� 'v��L���~�0�[o{6�XV��ww[���uް;í:b��te��y:Ne�67u��n���ߖgۑ��z$��ӻ��w�*0 ;_���_���'�%���o� �����U�������[E_WG`���򊳼�,�]ѵ]8�'֒�q:��ކ �G���hb����_DE.CA���Ϊ���32�$�T�53�q�;1�/;�Մ��׶~-;�3���:�]cI��x�
ȣ�^�T������ȥ�x�LU�9�!�{ދ]�|x@���^W�9�u�f��	�C)Ԃ~Í�A���^�9��ʬEp��&�P��GLц�7l��*�^jim�ڭ���e�,��~���]]�Mw7�k����K���=�����o��"e}.�3v�N�|���kE��3S�k���{r_rQ�3>c�PV����22�����&�Ƙ��\�J��ZD�OB�	N�N-���k�l];�}�W����������K��J���s�@&\��2�9~�ԣ��$�t��ڈ45�]]��f���@U������%��pu�Ez�nt�;+�X���V��'�)��>����k�Ծ}/iNl����Cer��[��[y��%��7o�ܿ
�+ :4O�R�VA��2��ˉ�r����]� B�ΙRYM!�;�7G%^D�YiN)��p]Y�$���U�
(6����i�0�&�+A3n���k,t�W�yF��f�2�eܣ.����8n�����E	cdX�.�7Y++&t~ē������@QW��̧Ec�����U%+:��,���±�0P��d�u`�j r�a$�֎Vfꃋ�˪�)"� �7E6�l,Z����X���Am�TVQUE�P��H��cl**-	ET)�e�gs����s���H�Ѕ���5�74ѯ�ވ��)���?i��͌kc�9�؜q��Ĳ�rG�t��'ٙ���]�φM^3��{��ܢ�����Ôc����y^����.	�΢��-<���U}FY�����6�Ժx�N������/�[��m�p,u·��!/�5Z�{S��p�\�Q})hԫ6>��R���<=]'u�K����^YB?[��M�nf��nOC�{�:=����>�>�	3rЪ�@ϋX�N�S���3��ǲl ���W�io���SM	/���L^"��܁A��U�O^�Yn�0���j�SG�_f��%��. <��u���-ȋ����T��O�.%��5�3��*�IwI��U�}�z�J�a܃�J�s���4�Nd�na���璗��f+�SޝMbdQ'37�-b�V�����R�F^�������]��כ
��Zy�u�Պ$���ދ��s����OѪ~�0~����F�Ŭ�zur=p��<	�1�L���'A��;��%`���y�^v��w|��;�mc�{�RJ~�b�z���]o�{�v��|���%]���=�j][ٍ���{��=
�;}ƥ�/[�V���QW�8f���MW��Q��Z��S��K�]���>�/f�8�xb�h�Us�kKx�o�<��9�`�ڗ)�#������<7���C����� �e����o�=e뵲�<Ͻv��+�����=���n�9"
�Z�n�Y�����b³��.n��.�2ŋ}':�ۼ������U��:9�k��^�97?2�߅�:_I.OՖ�Ū�^G`���m�R�&���b�gOn^���ɕ��1=a� w��O��C��X~�dn[m��j�W3ʒ��z�T5Ֆ���;��3JI�h\�3ۓ�r*�Y�p�j��Ҩ�> ���%�E��z�U���2���&�]�a݇�Q�ɖ�$����S�XN�h�nܮ�KBR�՜2�]r�5�Qr���Q�+ai��uG�U�q������|g��u���vv6Kf��f\L`%�V8�/��xF�7��iސ<I���O�S2��-���\ X�y��륯���K�F]�;+:����nc>�xx<��N:�V�W����To��[��S�\9]�D �'�z����]��ys-�7a�,�q��8��O��`=�V��}�+�p���AunS�E2�eN$V�2����nT�����*Sn�[�Dӻ�q��ee�[�(A�G�,��'���gZaa4(�ڼfŷZ�&�VJ�L���e�H���T�(S#�y���V��R�B�e����J�$W1yAغISwh�O(X�X�ɫ��4UW,P��4�(�QJ5U*�*Ƙ�(�e�t��T�m,F�D[����JAm�m�w(����)UQ�(kR��j���L��6U#(����4�Tj���*-�c`@�R%���y�{���v���ZDj{��By�űJ�ʗ�Ɩ���)�B��|�.M�Z6n8
�川�,N����2�	={�-�Y���ޙzrB{���N��s�uak�}cf�h�������G�eX��D��u`�r"�Z8s7��W	�h,P�螋͝Y���m�Q$�!�p���=���LЪK|���ӟ|��g[Zeu����H%�S�x�}����Wf��{./�yM<�V�p<�pv6{�� ��#���>�X�ڶ9
����O�g�,���tY�SCa�f����TF7��-���(���˯`���*��^F��v���h���5Czw
'�v���tN���t�m�����]W�_��i�{��yqy|����2��pLZ�1r��G#DVv�Ҡ��TC!|�������"���p*�i�ъȞ�t!ݲR�m�GF�X�9d���EY̌����E�SM��eu�.���N��Q����P�Lm�$[�l@]��=����`y�D^�l��Sq��(��fd(��s!�_�JeǺr��Cx�ð}���g�Χ�'�-18s^e �� G)׽3Wr�*�,���){��B��R�}Q�a����f%λs+ˍ���T���Y`W�ɔ��^�E՞��b��L�3΍���G:+��9�@
l�]�Ck ͛Ǚ�j��&�}c%NJ�_���h�Aqk����U[���tf�'�o*쩡���l�m���/A0��Dt畯q�Gzt|9n^�z��1�����H�A��7���Ų���S~��1Z��|r��-g����47��ckc�Ŏ������!>}�.ҿ&��|�v�;h-y�Z�-�x(6�-ݎ�ȬЮ��8�Ͷׯ]�Y,���LR���<��!n�VՑd�����&�W���:9̹1��ބ�wF�3��:dY]�f��-�(1rc�z>]�	[�^F�Ӹ�G�&�ץ+�w��G�AsD���+n�*�^������O��뼌�;�=��:���*Jk���G�l�B�g�jl������g�<�I�t�ȖEz�tB ��U�@�0��F��z�#�����K�cˋ��EGb�G��T�lP��vr5�Z��z�
��R�<QPա�ɼ4�Ό��῀$�9���"_�d͆IO[�]&L�S4�qc���ّ�w04V�kƤ'/m�Q�=�'�=W��o�ar��CxÐw[�We��n%�]^��'X��1u�#+n�A�]�m4v�R�fķҸ��o���rd�G6i�c.c0��t�Y/*�L�B�eIo1��^]ڔ#�@ ��*�Ř��r<,� g2�\�/"b�x��Y���-�F��^;�DZ ��V�n�(�mU]QmZ��TjQCT�JKaUR��MRe��(.�.��eSWT��B-UЭ\��ƑJ�(�ꪭ���H��7T��4U5%�Z�"*��UU\mj����U5B�R�V�
��V��U���T��ӎ@E-�޻��qSs�l��W���r2v/[�D][���-:'(I����u�P4=��[H%�������"�u���v�P� ���:���mv{�=��iՌF[|��f"<���+2w%9_4º���!:�6����"��5�5M�d�
���o]-Ϟ�F��D��+Pf�y���&֦���Ѳ)׽��9�����y�l�t���e�x;��x7\y���٥�Mv#7��n���|^�섍 �YY��M:�-9���8V��
�|c6]�d[�t9���L7�ct<}p���_e��%gH�I�T�&�nʆ�oM瞳�7�	ku��]�,�k�Ǆo��2�Y��r.�Ѱ,h�����n�]�lP?<P��Z�kx7Gō+g�t]�4�&�K�{ۻ�}l��
���/�{��t��F���u��ʞ�q�]����ÍДݹ� �tQ6m`kP��I[��[=e3�4͛���g;�r�9�,�ʅV�j��M��W�{��&�1�Kk�J��Q^g;�6�-�F*���W�p��/�B��7l/})L�!	y��'��򦵬�s/���m�he^��!�V�9y]�����O)!��Z��������*1H����;ܘ��^k�%ֈ�{���Y��E�=z3$�*ò���C)@�F;w4��4���#!����Y^siS@P�Y^�3�s }�ZD�2��S3��wQ�~�*�d2�����q�l^����(w�׭�z�ol���d�ͨ/xҡ�t���?p�g�^��sn� $�x��n�u�Td�k3��)�1Rڎ�b]�,S�Kw�Nu~� _	�f��OH��[����8� YV�,��z+/ U�s���7�`j�q�2��P�[��r"�r�m<������wm��nob�L��=kv��#9���XŅ�j��ڴ8
bEN�Ib�bP5<f;wv���#�	�ћSz˓���	���}�?@g��X=[[^>��o�6�Az�;d?m�.ۨ[R'ں��=�t�q�F2�V�K蛿ą�:R�]YY�g��,:�9c���RTm]ތ�J[`}F�%����t�~�<,����{&��� �U�/<���:��B�"����2�X~��#ܹ^J��C �����ŪO�*���w��7�C��^����u�+oP����u{\V��麊�W���@��t嘈�N��n͙e�אuۨ�r�[���Ɣ2��	�8�'nP�]v�<:Юy�'A��F�f:��#��[��]v��S�[��鷻�sk\��ݜn�����-:=B�R��}Mos-Jkk�U��6y,�`���1�\���a#�ʘ��W����S�����A[�݀p��s���]B��k$��U���4[%4�VꛩE5V�*�WM��-
)m�U�*�����T�@�b*4Ѝ[M�Wm"��lJ�UJ�Ҍ)eZ	R�n�[h��))�QQJd�*�*�)KaH,�e�m(ȈG�"EQ O�(N��βkH��{2o^o3��5��^�Y�#i%��װ�ʽ�S��S%���i���Lu�e�\���3n��;��i�d�Kҟ�]���{�Ke��,��P�t����Y����Aq����.f!\{��؃@����X"��4aQx�6kβ3q��q%r�aح��g�w��^�Geg
"�4��Y�� y3�:��-ۯ2��Cy6�N�睫o;����0��oǤ��^{F:-�^5q��T8��odf^=�P��y5����オ���tJ�m�m{=����,IB��7E�i���Oc~"�¶R	Kgw��s"]&ެӝ�)*_\�hnY��ǙRy��,���v'��N��~��N�J���{�4]�j��5�Hz����v.#��{�_Q�.=� �3{
��\��]�TK�p�Mi��y��s��Η�b�Fx-���]�.�|`���u)��Gl�)�x��ӊ�5����#3@릞*�ȁu-Oso��B�?El��k&{-s�rF��:�:]�m^��9���������.��6�^�](W1�i���2)-��<��
J��;��5a��2�m�o^�g	9F�~#��<���W<�\�l���'���	':�Z�n�����=��Y��ٴ����p��SͲ�G�����	�;C��A=Ӆ�.]����le�F��Ś������t����7M\��ikv��u�=;y����U�2(���9�J�)%���:�x��]ه���R�����ڰ����k����W�:v��V��Vpe�G:��j�9M�/([�x���l�.Av��4�h�'� �C��W�9<Uৃ�����+}=� 4�p�yʋU����W��:�C�0<����Y3o�S�t)�&��Cm��0����T>�I��!�q��aG:_���7�ݟ3a;��=ؚ��ȵ�f���q���F�f���]ha��O-��J �Eֵo���}�!>�݊��c���y�>��~�S�E4����P BB�>��H~�:Hz���E��J���R�^�(Ɵ�߃����$ BC�}f�l��#��@���H{03�T�f3�MeI^P|.��	�$_d6��J�w^�z�p�){��?:�s���󑗊��7��
�rY��^�!R9,=xfo;��@�	��;�������>�H��`I�!!�a�XT�}G��8������I��	����G�{_?����g�f}���>�������s�}LT��K�N��e�j}�����������I+�1����P������>?t^>�}�>�D�_�$����`@��ܾ!��|0~7��Ng�p v8U��IE��um���W�a�3w��x=x!!�4HW����������������*rw�!�:{�2O�xc�q��������_�G���!!��T�r|C�Cݯ��>��=������߯�\�J��~�����5�>��|d��>���~�u�@��~?W�~��}�@���}y��?I?�{f����y�}�>�'���$3�`!!���N8��>�)�>6Lp|����
z2O���{����G��F$�Ĺc���{��$! ��(�6$�#������]4�����B�kT}��aU��Lr���	���}���O�>`@�������q �������?�؟����{�O���O�,!��_ ��G������L����>�K��@�g��~^���������?��`E�!TT����9�'���K?���w�����!�������63D�
?o�FD.K~��}�3����t3������_��?��7;�|L�����!!�}��w���po�_NC�}�
�������	��F��WˆC��2I���A��	��'�D�@�'��=�?��	A>G���c�A�MS9��I�����s�ɨ{�P����I�z�����rE8P��~�