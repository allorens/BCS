BZh91AY&SY��2��fߔpy����߰����  a]�0�_@ 
     ���Z  ���                 � UJRUR���  D�砂*%EU�(*\�uE��j�����:\��&��w��N�u!�
��<�)ZU�x����
����v��uN��9i[-��J���{�H��RU[a)�R�hѡ� %q�i).؈R ֥A�Q0�f$n��+��u[2�`�	tn��P��������ȰI#fBm�C�N�ae Nvá��mD�8����F̭M�7���D� ��:�0n:Uƍ��$6V�+����vHlwp�� �b�Nww@�e��i�]�MeSmA���.̓�#�#m�Ws'�5I�vö���.�ݷT�����8( 
��R;J�)5��ǏݍKM%�9N�%ƻ�l�( Gt�0�]K���&������ڎ��l�w4�-�        h             �   P���T���#	�0	�	� & 5O�	ITTi��	��  �2h0��!�	�4ѣ4ɑ� �S�"U*{TaM1FL F�`M0
���	�5=5���2m@a4xS��@�2��!�Fh4�F4� �����#�8�	l���.��Ʌ{���r������6o��G���fm��6c�m�������	��ٳ|��l㞿���?��p�rv8G�*���c6l�9C�����Up�ѳlٺ��š�ɜ�UUUM��qm�����m�O�����~��ᷫ��~�\����p�~(ÿ�1ꙉ<"X���a��%�"w�%:P�E���`Q�G�xAI��aׄ�BP�ra�&'�
�p�3xNd@�3�%��&
�,?P���
��*>IǄ���1g���aɎ��Lv�&�X��$��m'�&8����nI!�3�2Dh7�xhy��q�r���&�I*S�S1'"��Ӆ��� ��|6�3��� �G�Y�f:IC���xK�;�8a"DD	F\�J��#91?D&�b��^f8"���jc�NTH�y0���1b`�y1�F�"x��a��1dG�L�vIN��Ç����$���ä�1���0�#�1�<Ye�	f5s	�"^$��@�1�%�LǊ$b>A�L`�#�0�'�{	�^L%�0�3YBLBP���%��dG�%�1g�GȐ#0�Q�����᫘N"_Y�YV�|�fbDG�DT�#q��Jx�$�v��Q='�<L�}0�aױKH�a�:a�$��	���'����tb �Q)�K�J`�I$F:Oa�O��_#����"[��Sԟ`���M�J#�������k���8SɊ(N�a�L"5�'i%(N�\G�%8?a����Yr�tD��HD���ag�"t�f0�ԓg�f,N�ax�pL}0�y�>�"<'H���Q�|'�J������!f>A��!�����C1�53"X�1%zb�x�a�|�|�A�D&�0��"yf>�U	>��DG��aĈ�
�"9鄳��	d�S0��pf�0D�BY9	e��$�Ye	Q	b%Yə�K+�K$b�LH�Ӈ�I�8�	c30��ل�T�tFc�D�a�D���,�f/�H�$F;0��c���-D}��:L���T%��B�f�9����<�p�γ2#��>�OLxO'�DE�(O7�%�b#�ID}1�$��D~��ĢYW ��O�Q2G!8"yȔ�;�x��D�"	�!??E��t��	'D�Q)���ı�D���bzx��)���$K}��2#�t�9�K�)g��b!�~�D��ϣ����G�L1�J@��&�$�"#��bdDf���D�I=�:SȔO	}����O�'��Ģ[*��1�8"P��|��`���D�j%0L/�><%�O�I�q��(Jy�X�X�0DZ��(���r'�9��P��%:"^$��$�N�5ٔ�x�i����}����x�f~�U	B<��#p����&d�/bRD���Ç�:'^D���"Q0���	c|��\�u�J�����^T�3S	��D��1E<��8G+�t}�n�'�m�L+,��ل}لn�e(Ϩ� ����Q�3e�ЙȲJ3�,��f���	,Af���Љ3Lag=S3Q�)��O!$O9��ߡ0E�J%�w2�"(�LfC� f,���c����L!u����Ղ||���/�d>U�s�s���? ��S2TP�b���:��D�Y��'&'�5'I�&|%��6x�D1e�8�J%��DHj'�F���q(�8[H����j-�$��Dj,L��P��-D�^BI�E�3��%0r$r�l�B"?1�D��?"B��Nu��D��D`����$DP�SRBP�X�-��{��L��t�D�D�D�#��P�=����\Dx�X�P���)���Җ&���cD��L�=�8<�� G��p,L�'��Q�Y�����D�~<"��xv��D�Ud�������0|��e��"���`���2�x����Q"TY-re$�����
%���b!,K��Ĉ��9Bp����Γ�$��#�&xJ$�X�)(�<��DIӃ}'���E�BtN�1�v'����	��t��
�J��:$�1�Ȅ�2��˔��w�JQӤ'���8wd�O$GD�Y)�c	8�Jbgݹ�1�d��ClO����y3P%�%����q>%Ȗ��g�U�$�����c�{����F�!��H����I}a"q��Vf�%��0���D�-L��>�)������Z>��k���9�L����bdN�g
��I$jfRFre$�2�3!�>���Oz>�����Ip#pG3�2�`�F)�&>fdG&g�@�_��":%���3��Bx��x�y3/~���"r؟?$���?x~f%(ϓ�E�O��Љ�G���D"�O���'�5�b!��$�%�D�b|Q�����$��"[Q3p��'����O7����L'�/bQ<�%0LybX�D�O�I�b~�`�N�@��%$I�'�~��{X��8'~��K�OD�'"(J~��a��&2(��xFa,E�$~N5�c~D��#�N向P�.c�=��Ba�fx@������;Ģ��~}%��8,p��������	y��Нb��r%,N���&}�p�L:�C�$xIN"Ol��"��D������'�'�N�#�GF^����u��)a�82NQ��ba������%|��:��f�_�~4�v)�O^��Q��~��Z'zt�鏼w"�x�#��,ĝ�8u�:��0G2aFp�DLB|�|�Ĉ���Lt�D$�D\$�D#q�O�"��,�Gɇ�(��L&G�,��a��	Bq�d�BQ��$����bNP�p�� G�GD���Ĝf0L9i)҄�$� �>A=u1B=��$�OT�P�ю�H��4�M�(�<A]�4�&<�A-�5?�V�9�q����5߆�|�w��J��b��?��9��3�`���g��9���ο��,�K�	��9<_��x��@������0����ߧ��������p@����������^ӧ�&t�ȦEba����8U� �-F��+p����|z�U~>��t�_�����Ow�~[?k��z	��Mᵿ��S�z5�L/��œ��u`�������g������Qw��t���������2��������\�Q&Q}�?]=�ߎ�]� p�$�r(�o�#4���
��x��#.U��{�eק�낚Ws�}����zc�p�`w&�ۿ�e=W9��W�ke7�fLx7t�M�<90���_o���r�9i�NfF�3O��ܧv޼?vɇ�J^*z�`]y��ݛΟL��H����ẁ�}ⴊ��������k�C�s<�G���JG��V�7�˶ތ�~�~����,��6�b�59���d����I���,��f摉s���tKy�_n����eX���q�c׋$�ޙs�ݝ���>�võ�tݦ_d}�3��XDMl���g^ Z���Qj>|,�٤���9�;�7�=�(B�}�t��˲�G���U}T�9����f̻p�M� 1�]e4*B�sJ5������O�?������R���B���^~y��gӜ�'��3Q���p!����	^%Ĺ'��Y>^����?�\�v{!���7��Χ3�9�k7�w~^�"�������?k�e�5'���6���������<��Sg2u���ѿu�����I�^�b�k��:[�I9��v�1�y�'nk������2���2Vm�2��ZEcϛ(��K(��á���P�������nA�O�Qf������og;���>��qϛ!��7#1_�.�p��)j-YJ�ٷ
!��ĳ��=������I���+���=��8�l�j5��0C���%:i��+��ٹ�OF����k������d'��rB�¶7nc��k�>넒�7@M���<�VsO��L\�7�77w�Mr��՛�љ����{�����{ƣq���n04V�{Y֦�?f�ӑ�Q�1����g4e�^���E�"f=�ZB4Vfx��S��u�)�L�9�XQą�E�o��]�%�m���6,�Ez�nz����ٝ1�LZ*;����sNk�t\)1��6}
o7\�8)3�|���3
��p��_�#<~R��ez@-R������S8/��ɘ�,2���ɘg�3�g���H�s��'�?��ݷO�Z���(�`����&�˂�6@�yٯ��D��g��$,Ml�]2Y�
aǶ��s�l��x�[�M�x�~���^�h��p�"ɛf�q?7�p@4����+P*�a䒿N[���>>�~���ٖ�j�|y���7�zuVot���I������n�\4��m���4��i����T�;�},KR$�{����vޛ3	��gni�$����"2v�%��8w�+;�����=���.��=J�ޜ���O�:m�ͅf������){�~�?a�m�h��%���I�՜�s��*�J[�b�̭J�(�7�3%��`����5�z�c]��T��$~���YY�o�NJ{[�K���Ez1���/�2^���O��I����~X�t"���q��Ke3ν̹@��nzۦHՅ4x������*���O�B��c��~3�Y��,�EӜ�[t��c�{���=��5��ﯧf_7k��H��ó��z�+T5��^ܷek<�f�c�Å�`���,�'7��|9#�+%c�}*�1&��f���ة����{�|]͇�I{�������mDzx�>ޟ�[�1�Nr7�e��:���#Ҧ=٘k����j���4o�=?z�����x~3h��3��Y��h��f�A��Ѩ��CJ�6l��ɔ�ޯ}52_��Ƴ7��`�u]� ׌#�J�\n!��C<�¥l��ݷ�4��_7y���^��h�q�|o��sdh�-�t"��%����kۻ��l�a1�ST�ۛc.8p��ʺT+-l�k�u�����FS�{���V�6�w<��~_����섣St�����YC�}���u�oK�mQ��)^ʟ��~�KL����;��٧??ݼ9PNA�G��VW�Ʈq;����X$2L����;��~�+�F�Tp13���+�1>/�ch��6}n����ޯM?�~3����YѨ��$��6i���q�דC�q�e�Êc��^��(�a����2���=���g�{=0vM�o���b��x��{�µ�G�s
aq��L�������F}���s9s��o�����,aXIf�Y�����}��tڶ�2��=������+a�3߽�Ӟ�OQ�Ef���狌�����}4v��h���iM]qG�=x���EA��>����|x������ߙ̇����yxݗ��I�v���8t��u��N�u�:�%���z��$����p�;V�y��Jh^�w-��}��|ӭoc�aㅟe!�~�0N=�ޘ��ۛ-�95�q<`S_<z����/RI��/�����w����su�����'8���m������q���)��w0F|����>��4s?2x�k�]?���z�g��93�(�^mf�q�v]%s�,<8/����0����a�̾�{#�eu]#N>̮��3و8�]��&q�����5�f�w��Oc��1;�����_����0���	\}���~^��ݘ�x;�-;7|}�ݨ,��RO?Ǭu��������2,]8\��\tُĝn�x�{���~��T���=?D�*?����gu��o��_\��z���L�2���;0\Zm��ea��r6�kh��<�7�s�v�|s�F�p�
q���	|~����I�խ��x�S�{�w@|��K����x������q�#I�K-�߻,g�zv썒[�.&�}߳h��i=���d�����訨��s��1�1۫!*<?C^���,�(��_73��1�pv"��Yi�	}�x���BxI��a'�u����n��~�{+�������*���ֵ+=Ӿ%r��P>�d}��8��?��r�����O_���[ᾈ��oL������z�=Ěg���|7�����?��pi.��$�|\a��h��-�f�i�Z�j�-ݲ�Xۺ��6��!7tݔ�f��[��ZV]����IK,�6Vݷl��]�h�蛤���l,+��u(Ͳ�%���4�-�fGwPJ]�"���f��HݺRo�q�lH���e��$�+$6��9�1��f�&���8jk��n�q֒��5vf�l&���9r7�ݞ%~���es�}������#�����M&�d[��s8��8]�=��s4�H4�I��h��K��X$���O����j�m�mwu!�������=Ӫ���	G�E6�-�c�g�z��Y,>�>��:�9�G��=���ZS�}�h����A��o~��r���Yu�Kj�kW
���ٴQ����\���ʉ��J݃�7&Y�U�L�k�ü�B�]��¬���f�P��Ӽ�&�5�aj8�FX)���"��<��|Of3.��ss�ro�ʸ�1x����EƷ9͠�b�^\���b�~s�Ӝ��.��;�«6�dD�Fg7�F�p��$N�4<���:ҸN�>�-�̈́6A���:!'˲+�-�V���vm�"eQ\�&��3���R'��8�M�Sl1�^�P��qK,�#�"����a�Ұ)R�_�$>��"@Sg���N���m�m�2N٪�J�~�nu����Y�빦������U9��ǮqgЂǘ���|u�C�	)5����>`��>s:�!m5�g��-s��u�H�GՋ�c`H�8��
�$4����>o�l(������^s����Y�^�����q�A��à�+�H��n�ݜ��e��#��g��neb��g
1X�K��g�$���u�kb��y��M
�9׎k����p�}&��>(V(X��<��ᢑf�f�>p���O��tK^���S�`���$�'��%���I+�L{��s6�a���sn�Y�Gi�ǉ^:�~�����Xn ��@���Ll���6�գ]�,Չ�A�o��̆~mQ�i=�{/ށ}rf}���W�9٘��Y�.a����x���}hg�;�L��N!���2������p�@P#���]<�8B�~����
CF��t���_ G��6�~������T���}�������� B �{�.�y�9��g��_-ǵnk���l�m����yW��vه�?=���8�	�\�����~�v����f��=�q��������������x�����k*��ZUxʯ��U_*�V����^�*�ڲ������.0���U�W��Ux��V�a>�������菀>�#�"��#ʯ1W�ʪ��������
��ZUW�Ҫ�������Ҫ�W��^�*��*��ʪ��*���*���U�}�	|}���D@}�ܘW����W��UiU|���k
��
�����v]�ڮ0��k*��ZUx��YUV�UUVUqU\aUU��" 4���wwwWUW���W�W��^�*��ª�,*��wswj�������0����W��U�UmV�W�ʪ����|}�D}��3V6���²��l+Vǣ���ov3f���K~_�������!���{��|�{��ݟW����'
8A'�D�Ĉ�Y��	���&$	bx�,K<t��DD� DD�&	D �(�H(D��"`�g��	�� �D���,f1�X� �
�DĎ�$ ��%'D��'�8"a�'��,L,H,L0L(Lı,� ��'H DN��$	�xB� �D��"�'J:"tNp�LZ����&��[H��s!ʏ�aDS1��SrH"�z|�-�YvHKbB�����RF���g���#I84����"�6�o���:C)� tC�@�9����]M�l�����R@$�����T]�ĘP��o��MZ�B��J0�����mJ!��]���D�	,�>i�X�1b'���#�&��Z�;F�ʖ�Uֳh.͂�-���s.��f�ll�r��h;�6͘O;���F�Y���f�#0����$��d�.�5�*7k�&�e]ջQ��AƠ-~��AH���).W>t"�(�(��J� c-��2؏ŵ'���.[E��R�%5ER+n���Vd�[f߻9��[_�h
iH( �B��1�CA��HV���m�F�.�mr�ewSd�vXSvI��rJ��� ��a�Fc�Pх���5,%���3tDf#�Z*R�I�L��B���v�]lHX�6�$R7N�"�겶Wn�ܻ��Y�j���a�K��rED5���^K1��u��H$���lc��A�k��/l��Hku$#&����i�=z61�Q-n���b�A�ۆ3*"�(�!vYm儲���r�H\f���۳Xv�L��$rHI�����AO���R��V��v�F���ۂF�h&`��b1�N�eVjl%�Z;m)�G�>�}4�rv�R�&!g��v�l��.ݻrU�+��t���Dѻ>Q"�b7Ah�"s�LM��f�1݅�[�[����X�l�esk�[M�J���iyx.���*���N4�
<����W�I��$ф�K���wev�(����]-�%II�#�d)6��ȍim�o�����6�b�$,KZSf��M�QԶ�)�fKe���T�:��l�I�c���ۮ�L�w�Scl�II5#�����M��7/R<��Ͷ�u��}�i�Ɩ�S�kD��.@csX����#%{Bn<��.��6Ĥ�XR[6�IwY5kU�߯n�ⱶ^\��n�`*1ݣ+��nl�n����I�d�+�ֵ�n�|�R�e�$٦�v�26[[���BB���bW�� �ح�Ku$��Sw͜����#�M$gʣi���/�� ;��1�8�U(�`����F�"��If��c���v�k��0�绷����������}��|n������ݻ��|n��������|����ww��t� !i�M<i��a��%�%a���+��u�T��&y6A�vV��Z�e��)i�XQA$�m�����P��o1C0���$�tFmd��ɖ�7v�sI$���mԓ)$I��I��+��4HCj��-m#vY]f껭�Y1���.��pr�c��lK��ɭ%�R;RF,��A����I�aJ|R�n�,�Ko6lѣYf�n[��.si9�3S]�Ũ�I�j��F�d��͡o�����a#��:4����ֹ�/5w��;�n8��r#���"h��(��� ?��BN#��A�������h��uA�����JG�5]��4��<Hp�{��a�1�Q0L��� ��hȎ� �O��@�;٘}�n����l�x�:o�bA���9Ξ��,�p�$�ߠ�0�MD�,�"P�a�L���k����B�q���'@�_Ge�h�C�f�|��m���3>øi�n�>>�a�����LX��B�t�G���@C83���!Oo�����n��GV�Sd��=Gt�T_�(9�0��8�b$�E��e��:&	�%�gD���:`�>�z� �&��a�ɐ������t�e�=9��i*J��>/:�<X6,,i�+E�;��
�$�n�~_�×�#��Hٗn�K�Ȕ��|{����=x!��<E�)��^�3�=���fgs�_�6�/'N��qMn;=؆F����8�;��H4D��ĳ�P�ǃ8Q���6�B��)hi������Y�n�D���w�$@��U+Y�*�GZ��Mٞ`��q�́pI�Ucp��SU�Z|ׇ؟g���۟��&!��D���a�'���rPQ,���#ĢN������"�}�=�@z�ӧQf�A��X���0�,K(J(J0�Gm{l4�ߕB��0��	4�Tr��I9T.�a�jDm��e���n�a""�
6�A��4Yme��l�]Y��4���@%�#���K���jIs��AD�0���k$D-����u�P&$�#�=�N.��IZS����<�!��	�,���o�|IC"<�%�p�0���E���0��8�Bfl�ў+�Ǥ�̜]��74:'0�z�a6t��?{��=m#��p��tpB����}�1�&xD�,K(J(J0ç��O���jԭ@\ʕl� �q��L��1Gv�2'�^u0�i�.�!�5 5�p�_>��C�nm�p�W�?����|��s��L9��>C�����l��-x3a�'o�
ˇM��C���	Ewܙ��d)D�Do�(�`Í��6�H�%If�4����J�0�xB�)1�����M]�`�S��l��`��1s���8�z\9�0����a����ӝ��y��ƴ�Z�7��g$�3�.x�L������Wh1�qO3��\���釬�t��O�a��:Y9-�J %|	*J 񧎞0��0�����:`�}�\��ܞĖ�c�iy]�4��9��^��J���)ID�P�I�U�1Cȃ�9�o��K�#ެw�����'C���D����ЄJ RP���(�8H9��`X���I@2�@���U�t(���p��0��d�B%	Ft�<'o�L��;�j>�"e$b$4�����BIԵ"T�kLK��Y*�6K2�Jb�V.�:㢤�L��,1	8��~������=�`=�Ƀ��X�b���W�NZ���.��g��]����c�� ݢ�#��g��l$���1���nCʰ��B�p�=�87{�d���ϱ�m
�ʏ݇f#�X,�? �~��"�J$�aB�I��@�ӂ�y�8P�8|xy�3��	<ib`�a���J�(��ü�K�	�ߙ�`�9�	CԶmG���Q�2�=@Vq�u�!Q��(�4�tg��Y�c�އ��~b0rJ~�y�:C��KF��@�Cc*�V� (b�@�k�gE��[vۤ�����O������ �����,`j%����Fכ�� l��,�X/� ��a��?D�tz>�NC�4�(�
oBI�J&��6�I'M"
4�ia:F�t�4�� ��8I�$i�i�I���:=4�Ne���iA����重*G���4��Ѝ�i:Q�\�6^�N�i:?��~4= �A��䰋�� z6=M��t�4�#GI9oH��dh��e�=4�I0=>�|��?�#���||��=<N��J&���&��h��L�N���I�zQF|a7�><F������0=��M��Y�i�4�=�d���э�P�CziI�F�B�Hp��z84�F��N�M'�H�����4�{ts{\�0{�ڔ��f9�vn�������zf���`�-�f\��;�V�>O����q�JB�������3���U��K��Dӻ.�Y�1��7t��:�.��0�N �K��&e^z���Ǟ��l��+0�Y�b���������t��c���d뺦D3�[�^I�����λ���������wwwn����t�����˻���7�ݭ���˻��4>���Y�h�%�Y�3M$�J0ÆpӋ���%��i'�p:�en6z�\6�n&�k!���x��';9ɻ����Bp`cB��\! ��	���b��%��2����F�%E�u֡!y;8��A�p��#�� u��1bI"��T�כ��y�I�9����M4��a�;��&	�L�v�j�nf�<�9[o��rY��xy�(:0��A���i���Q*Ha��-��|о/(��M�R�T�i����x�8�0`|E2!2�R44|x�F���� �"�34}�E�jӌ�9&yY�V;�<�w����H��:x�L><pÆi�IF�a�p�7�km�Y�9�Nf�G�ͬ��N��V0�a���1Dʀ�h�b�3M�|<��i*�j��]�eu����b)/���P�Z�P�_"�3Q |����L0�4�7I������.a�����P�1�D-&��8A	�dCsDfa\�Vf�6g�&`��i� i*q�!�08[p�"�!"�#`�P����'舓�G�1 X�X�{�n2�8��c��t4B
h%� Ja��� �C`�17	�tLP\�3��9�v�#%��e�m�N#���&��,�	�!���̘���d�L��
4�ӧ4�����00�H4�J4������/%l����a�:�-��
�AJ�r�&��XB� �
[m{D�&%d�!��q��qE�Fۉ&G%��#n���k6k.�g4����EQBÕ>�f�Q��D����ZX��[�e�P۷7,�F�pW%#��r�M}2��'kYP�v7k��p�G���RT0���BCAD�M�m�S���q��U�r��ͧU�)<�pΑ�,r�L�v�i��|C?�+�L����'���`O4q�R!&4�gĥ R,��v[q9I	�[��˜䙄�0���s9�=��S�W߭e��läd!��4�"��@����nc���n�0�s*��n8Lϰ�\:HLc��sRx�	ă�=!�s�2&���n@\�9��?I����)l\#���a�aḪ�*E&�)�	ń��f���57$
�,7�ǋ��a�%�BSp��2�,�O�4����XޚA��iea�:i��P1�7N��]j�I,��f�N�:B��8͖y��sl�[��n|:����)��s�Ƙp�3I�R8�lI;��2��V�d�nn��8��\bI:M�c��F
FR"�L�H d4C9��A2�"$�[!L�	�z49���'�4����<�AO�8i`8B�D�e{��Δ���鹄	���F�CIS cK�T|�2���n*R0}+����
;��5�ͤ[��J�m.!���ӈ�.1tp��C�<e�Nc�"S�33o�clC�>� �����R1��hD��C=w(!	��PG��D�^nQ�C>"�lq8��+<ƐkS�<�ۯ.2N�"��r��y��?~�DM$�J4���ig�gd�XI)���C�E��'���"y���I��!��@�(�!8Z�).0a,`Y��G*��&\����c�a�#X��4�@���H����apH��r˧�I���"_�窚�\���s&��Pw�9�8�ӇRB�����nD�"�_J>�i����mf��X)BfY�G�?�14]����\�|xN�#�s��C�C,�0��9s)�#���Q�1�DZ��`C�PРi2� L؂�1�0p*h����qInIT�L<4�Vn��c�Nv�m�θ9���ۘ�M�Ntw�si��D���i�Ť0��IP<�ᒕ
j�
�pk��x�<~���00��4�K(�i�G�|�DL-nJ�CH�)i)������`".g�����,�J2�к��>$$C`P�=��ˢ�xg<5����'I������3�w�N�O��(�VHI#,�4�3���úb���\9b��2ɷ���i�D�Q$ i��>D
Z
 "Hy�q�(�12�%�&o��-���J؅>�C ��Zyi���$s���:�q�,��88���X�[wN6��?a
��;��I�78u�s0<��`]:BAL:4��+n��W�F��YF�q��|40��mw�D}��Z0����Bm)��eG7�/��7��᭞)�;ۍ���3����& i,>(��||a��M$�J4���if��V����&��+�����>mf�����T,��wX�P5kQI����t$A�@�ͻ�����m�e�vi���S��-@�$
H�,~�I'��߿�/"t��Y��q���j�r�"���㒐qOs��\`�U��ն�[�&�ǖ�ܜ�u����q4D�\̡hÀ�543��D"ys�2����Ď�P�	���!_�~sa������?���#���wR�P��&�������$9<�d4v[ �c�ѶApA�f"��p�̩Բ|�Ky��E8����5p� d L��X�:L��:Hjb�)8��3��Nl>8C�A7��3�;��
ANu�M!�k�~?^l�m����7gL�w���������Z"��@1�F"P�|?���\%.�ϧ""�X΍1�$��4�~?	�	��i�t���4�Dߜ�ye"��Wp�i����sa��Q)���O��w�jQIOĄ�T��rX��$>�-G�vۉ83+�R:�	(g�Dl�IV@��3!�pp�s��(��13�x��h�*�Dy2�\�P��(ђ��1� �ZL��JQ�Nd�?9�v�����j=��X��gP�<)��s�`��d�/��L��:��e��т"'����n��a��~E	_
�lh�p��b�pd`��!�9K�9$7E8$�d
l<�D���Ėx���M>0�fA��iӂ'���'y5?WꚂ�\� ��/�������&��"��E}e����;#b�󈢋LP3HPZ,���>�����̓H��A:��l�(0ӈ����Hddd��y2җ�G�%+��s�&,��������1�G��e�S��ū�9���ֶ�b�u� \L)Tj3GE8�G�CܼXPI�{����M'<��?bg�&���s`�z�O����($��H,����%�W�q'�P�8�D�(b��c)��krw��(^DQ"��(�è`@���KC$�9CLY��Tu�$K4�?��x�~4�M(ӧO��g�~|��.l�I��J7�U��x?�1O�<
d7�!�<iN@�.��Z(�(LD�0�`8��7	��;|y�>�wJ�]�B��g.���<�wv��0���C����
7��'~�fY8 � <pm��ΐ ��HQO$X��ra��LɈ4�����t���)��e|_�gxe��[q3F.�{Z��h���bW8|0y����đC8,��m��[�OQe�ڈ<�+GȔL�N�H6	 ��K+��Ie" Q��K������(�<GG���8AF��K"�"��$i ���ip�I��dQ��&����h��xY<��t�HH�M)#D�0�,�ZY)���82K"���饒�#M#M Ӥh=(�6A:M���O�#M#FiF�V���Ѝ�������4�XB	8)Ȫ���7���:QiAI94������(�4�zY:I=��ޏ��tGó���|r�ē���tzaM#�I�5"L4�ӄ��Q�N��a�?G���t���C,�X�zl94��A�HӦ�zl<"����S���x�I �HL�4��>��|9>"�G�|Y��t����O�>;�Xg�l�����gu�b&b�2�3[a�* �u6�1X3_�&�Eǽ��U�=���=Gq�{o��Ϭ}�ăҐ����x��`"5�M�رQ����kk��]V�幔��q��}�B�&����g�4�aK9���acX�a%�V̿)��7/r��F�j�ɴN:�uG�}7L|���"2�L���yS��Z$����Q
�ї�9�h\��b,{��H�^�"���{'������W<�z#4,�;�=�{���+{Lm�]�@�ƦT�;��xU��V�g�0��x�L��l��zlXYz�}�w?g6|f��1惽t�-�]'�/��v`��Ǫ�������i%m��":�k]�ݥ6n穣g�\���j%�������϶鰤�y�ַ�DM�kӜ}��Ö�#q�m�K]���f��t�Q��B6����$F~��h�}�����+���fb�QPcm6dn�I�]�X�iNR-r���:؊���Cq�/E�)�<��� o~�����̻�ª��fffn���{�����
���fff�4O	b"'��&�I��iӂ'���0��QQ2O,�H�V[rI1�#m�+7l`آmwmj��%�)fk�l�I�������j�l��t�]��a	�����k�����v���j�w5�]�䲎YY6ɧ�p��t�×wKeIu�֥�l�M��v�l�I)7w+f�,���))ke!���J�]��&˫�Dж�"�%��j3L��F7wlؒ��i��-���]�:���[Gf�6M\�����UD�͜�M~r6��r$�P���;`D)�f	_�ϠQ�ǈ��9�#�tR{_s"z����6i��+�i?㸞�N�즍�&)�pv�ᾏ
8y�ȣ����%gC�-�I%�q���>�c��]5��G��w�1*=��o0�9��'�&�p/F�C�p�)Y�t;���4��I��,����d��iH�Zh~?��Rz�m�	4m�c�d�>g����Y}t�C���ҧNa��pV�zx��p���i��,�M4�M(ӧO	��v}�L����oS������җc�������O�)X�����;}(�Z^eG���^5b+�|$ad�H����lp�ox�"�)��k���ϛb��"ٟ�)AҔ�2�c��{�����{���C������MtvU,�kM�'�l��Aá#q)�$��4��j>rI���ϊ g� c(Γ�Ya�0�$���c�L���gW�u(�@L���?��Å�|i�I��a�4髬�Q.D2�Yq���!�nNύ͊��S�7�����(.�h���2��*�H��@)($X��6-`Qe��b�;��Ja0���7��-4��/��Ox��9o�Sb�t��I��kY�E/����m�@��3e��N��t�e���ȫR���2,]Gz�$�}L(�FQ=�Ŋ�܂�Y�A1>���G�_���7�S8�X���Q���Z�)��#�_��	�ꕤ4�~�DM$�J4��a�:iң��,�G�O�[!�u rL��9e����������a����$��Pu"�tQD�Y�i����՘}�����.�����n�8ɸ���t}9�7aR�)�b$��ܯ"�����
G�����Axs�5��a�-ʟٸ4��Zg���4�B���Q!�	X(4�w��!�CF�*�����A'C�Wăh�Aj�!��>+�-(��$���!�pኖ����<i�p���A��h�<?-�(<����0�Ys^m�F[rY��&��5��r�=t�w����/v~N�O/8n�6��p�AV
(����i��(�V�ald�v���UU��o���T%g��<(���Q���������<ƒf�
�ݔ��^���$v	��uve\n�����B� `�+�����%!=H�ٓ<,7)H���H��rA ��@E(n�Xa<G�qp>��X��� ��AcD0%E�'z�5�Ģϸx,�VB9D�3�<-���D#=��M]^�K)0�׸54�t�V*���d%��r�]����M\��G�ú�j;��.��`�t�$�9'� ��<||a��M$�NQ��ig��&v(��Me�V�������=��������\=��/�vKa�|&����"`qSc��lӾXA�����J�:��D(g�m"*�A'���U�3M�!�#���2C�3���ϧ�K��B�w�k�ͻn�����Օ�d8>O��'�?��~:SjF���	�Y�IH������>E��I
T�>f��(k����>����X�$�k~D�M����Ĝ���O04�M8iGDO�E����L�N?c�ǈ��$�[B �G�u��s5Ӱ@|S
�iH��v3��Z�CN�yP=�} �,\��p.�R���Ѩr[cc�Áÿ��A����4���Mu�����/f���s�F�҇ٔ����g��|�$���h$3�_ �D���+��U�]Xi�6ƨG�e��8(�8@L#N�Ţ���$�I�>><i��,�a�4�J4��0ᆝ9��J\r  b�B	K>r^�ǧdgy���8i�U�����E��ߎj����3��7a�����z'�.yT���7M�[c��?�F�6'��\�ā�r�I�n��
V�(����r8Y\-dP<D���x��uI��m�衲��ng>�l�C�t�ԯ,�>E��BY�~�2"f�:zo�E����h�B�=��@�Ո��IK�pRID<t�>0��4ӆ�pD�X�v#
����-��B���T)�����H��0�(宗�@jFO�%��%⥠j5�M�"��2`E$j�^������矯��g�)Jw9�7������b��g˽s6I�T^�����V��[�@���K!��+����J�0O��7a3��r�nwA���8���6YwѲ3�|��i�����pzC��<'73B������aL���g�t�K<ۇ���{��>))?�y����罖�I�Lm㈥Yjd�SaS���0<a�8�(���ϡ�aat��|AO�<x��x0��i�I���O�Ǉ�������!�o_�ڭUTA����I?���s)��*��"y}>�����k���G
�OP�q�Ձ�9�!�7'�|̠�+�gͮ#��@[`�pԢ�����9��.�ͻ���@m�#Wᢍ /�i�N�BA߈�|>���1Ѫ�,�43�n֣�3��<�����_"P��8�� 䃅���<F��I��>�N����K"�C�H���4��F�E�MΏK4�24zx�8JF�$��:@�OH��g%#���G���ӧI��:=:EC6���zE���tzip����J&���4p�(�zY��4�4�tg�6Zz#H4�C6�X8n�e�1�3F�#H �a�=#4�II=���h��I��Di$@������Q�����_#��><F�'D�4j7鍘I�0�4�'�0�#��i0h�a��i8i)e�ٰԑ���$�<;4�:z_M$��K#{!�C��k�K� f�2ь�0�4�i6i�=4���S�dd~��D1�=u��j�)��`g�"�<�r�[Z��[^<��5�F�{E�5�7�Ϡ0�u�;>��N�H�ez;̨�a}�5{��.vwe��`�|~�rL<��Y�%��O��RWX���p�gĜ=��,���f�z)כּ�U��F��sr�&�J�ɓ��mTl��˒^��{sc�s7��x_����c�K�K!̓F�U���Ϯ�"�ִ� ���?~�������
���fff�ª���������^�ffn�4�K4�M4O0 �M8iGO	�����ڕUQa���$I4�|�	�[�gF�Aa��G}�7�14Y#��~�w��IK�=;G��p����﯀Ї��{p�4�j3H[)G]v���e�����a��1�o=���1��Wͱ�7��vH$4�����%���������8���a�r�#y�ޕ����e�u���*3X�x�!�3x馝><|p�����J4�K0ᆞft����(����q�~����A>�>�:7è�rW�p_8"��u��2����xt����m�5#a+]�����|9����d���xQ�3�������CD�7��\��E9N�'�=���$��i�4��4)����Q�G�Ec����P��$����D=�0�xa �\<{��ˇ1�����#Ŧ~s�~�g�B ��N<x��g���Q��Y��B�|p��wfl��(	��Ú��eB����lH'z��2"���DHqt"N��+�$�&A\��v������eo���M��kRC�z��R,G>%�=��I ���ل�LBI�!8��vf-bؙ�)J�^�mF��K����4���{��9�=Mcn���a�~~�����!����"���;�qޚ��ZIݢ@��tl��8��uyFa����x�h��p���,�f7v�ag�>TX��0�!������Gǉ�'�Z|.���Pd����,�R��	�y�u뮛��V#4���,��$��_�C��W��<`�Q�L?:`"A��Q��Y�4�۶���18�s�UD<��x:%D�Ä)����%�\8B&�8���D��|t��k��X}�Â����x8J��D��=(���4�Y��rwm�KRZ�y��y4��Op������!�\�Zr�������|���7qϰB�Z�W�)�	 �����,�a�4�J4�K0ᆝ��Ա�̷-�,i�i+�*�!��a)#<]ə�1t����B���!�����a�GS8g���C5Ci�R��?��̤�?�|Hm��GiS"Z�%���sh߉Rp1|��H���p��ĘIe�c��E}�}���*�}�]?�w {�t�ÿ�e(���ޯ�t�n{�*���Q�Y��p����M(ҍ,Æt�u�46�c��E9Oު�!��Է��jSL�9�+�}ƶ~���֤�&�nɗ�i[gO}��&|9�تL:O��N~s�:f�'HG�a����1�Iz���8|gQ�H���>6�T���A$����ڠ�p�|x���0a\ ���ӇB#�F� ����Ǐ�x0��|iF�i��B��|.�E�5�YTe���HD�G
u�Yښ2($97���n�/�������I��U&�gvs�y�i,�cɿ*�k�ޓ9������B��ΐ���#э���1�Ҭ�]��V���^��soB�Sꚣ���v'�B��|�ק��z�$}?wpO�9ĳ7v��К-ECᤜHX�qG�-G�����Z;�Ѭ��CK����K%E��)���a���-���ӋT��2a�	\���aI�Z�,�5��T%�@�h,�����38�t<��a�L���L|$����d���s�(�	�wJBZ �~�z�k=�ܖIx񇏎x0��|iF�i�i�]r_�шk�uG*El[���9�����O���Uns���F��8^$����!��P���51� 
��ߌ ���4%I!g	E����Y���$��X|O؏/ߐB������a�QW�mm��vŧ>��"���)���@��{�#8"a�y�O��/sN�/�(<��l�QH��L �0���<`�>4�J4Ç4��6��4+\���!�n)�iM�oʉpӡ�C�$�7�w�D=Ȟ�2�~�I4���2����3�L�B�������lt���4��.*~�6x�OQ���Z�Aध��A�N���D��f|ahgJJf ��A�p�xd��B%��R)Ko���dT�X�Z(�����:����*CH��t�O��||x�8Y��a�iF�i�i�peW�@�H���Vk�;�yzp���9��t_�C�a�P������R�m��P#��X�.����O=�?a
��4..`,0�o��D̮�,�oņ"���Z:$��tcn�ߑl�0ãco>3��璣jk��ܝ4#�U�K�M!s�aC�ђ�~�I?��#���0�9*oB衑c#aD{G��3��xg��=-�t��6�őGH��$p|2 �C4� ��F��'N�i��GM��z#��Bi= �0�t��i8A��H��<t��C#��H4zpѓ�������DI�8&hi4�t�(�8Y����4�I����Y�3�A�����3H,��E�p�vѳH��H�a�	#BH�H���F�M"��e�i�kHf����W�d�p�������4�0�D�4�t���4���R4�4���)�0�|ޑ����2_H��T7c��zG#K#�����|i=�dpz6i�jќ �� f�3a�i� �Ie/H�Hᆝ*�p��.?�_jFѰ��ڢx��n�C�����Y�1��\�X#@8G8�l��JKǦ޿��r]��N�V�KY#��I�˺����X�n�)��pc�7�Nj�˻N���n����D�X�r���쎐�y>fUA���Q*�kYL������+��j{}0��*m�ߗ܏vo�q���V�"���<�0tq���h4m=#sM�vy�U
zeސ����a�3����c}����ϛ�;�X��n�<F�<��6_bIm)���;^�#b�~
X��Rt똷�A[>���g�/^_��ڲ�e{�S~�͌��?�[7��^G�Td��2���}'u�^gq��d�Ŵ|��U��l��,�af]Kv�e�D����ʁc�qVHV�RI?lu�{�Y�'&;6�Z\��)�m��]�k#"&�坰��w�%8����(����[M֑M�j>^%�yY��v�	�!�;T�W��zB6��0�
�����1����"g�p��rr�y��v�F�����33?n쪮f�ffn�ʪ�nfff�쪮f�ffn��M(�"`�:X"@�i�N'�	��棓Pr�jb	8���MH!j&�n6ą����6�Dn�lӼ���/y����<��	�Yʕ5�"k�C
������&��MT䌳M�M$�J7me�Kk6�+&�aUt%aY+md���K;���e��n�u66Y[Q��ݲ���r��Sf��u%��%vXݑ��KJk��YD�i5���ܳt��wK�,wa!#��뭋���ԋv\�لn�GqaG���Շ�niRR�B�o9��E�SvY,^�����?�'�ߟg���;�G�����/�X���8_%����fgr�K�~�%���0����,��%�U�K,�a�p�ţ �t�C�4Aۋ�����p@�����dPP�\n	C(>>���_$�D���'��pAhk�P�;�ǒ^>��L�7�$	��DNJHj}�Ews<���~:��2�����qxçO(��Śa����&�pӆ���idd�w��i�q�fU?a:z���¨%�����3�� ΁^�8P��2�@u��7����Q|�so�FJ3���F�La����,h8�����gX�p�, 3qq�c-��Q2d�Ɇɀ�T���� �:i�H<_��(ґ�up�C'N����"A},Å2���e��F��IGM0���:`�0ҍ(�8a�N���y�`�Q���&���I?|����|73p��D�ۊ?�=��5�}�������Ch�" ũ�A�A�R�6ܘ9(�u4@�������/�xZ�-!�������4�C r�p�������i���h��ޔ���^�:}�����J ��n�,��p{�6�ͳ�l��420qc�Q&�0�L�KH4��Y���\9b�?9�X�uUQ�����a��4r�$���ĩy�9��|�8�IG ٖ���Y��QUd��	9��1kld�Yt|gx�-.A��o�^7�7a m�Dp�cBc��a��DA�0`��շ����2��>��)����>1��dsD�~$Βx��CK�N|Q8�f�a0�~0�Y��M8i�D�ig?'��	��9�2�G�e;H<�CX�f�j"JG_B2�)N�`�a+w[r��t����֓d#�lٓ.���ߕU�=�o����ٸ�-�5�6^�� w��$�s:sZ�:M({��h?%�i����M%r��>J�ƈDcREd���Ȥ�Lk���<�I��:���q�B:�b�f��0���P���e��5!	@�#�#� �

��pR=��n͞}l���m��A,TuM�T��Cu�3b���۝.xC�t�0��-\�M�(���e&%TR��H�Jw�i�gI��e�"f!pGˇ�tӧ
>4�?t�D��Ɯ4O	�K���,��Y�,g5���UDCH�8 Ϳ���(���/I�2�E�&6���l�JáG���Z@�C�p�����+��́�ppI�7~c$���K��13�~⊯�>#<�ޟ�cfx��wU��]��v�B���m��x`�ѵ�Ȑ��3�e�I+N�C���� 1Jl�qd|��Bkd
"J
��m�n��@I'Ɣ|t���㥖�"Q��4O	�K=ꉚ��U.̻8��/���?�UTCÂ��is��L����K���7���N"8ݝD�c>	<����<>M, )">����i�{��a��~��*H�m[���s���`�t4�"M:��,i0�R:PPp9�NUD͎V|O>+�p3��ӂq.�8���(��Ȳ
D0�x�눒N_ƞ�X�<i�a����$�~4�xOY�����U�e�ꪢ����ǳ߻e�Q�VHt>2�� �~!C���"��4���^1!M��U����h��b>>8P5]"5Q����4߆�Cc�W񆢑L�Á0A��D�qCT1�!Z�3���r/�����e���a�#�O�Va��&1�vHc�r�(��@|�%'!�p���&�~,�`�%i�D�4�R֗�����)h���9�
�+'����/&�Xa�l��b0c(����nLY�Uq��đۭ��h͖6q�U�-�Đڋj�����UTCϾ�y!>B� &Ǘ�!���H��/p(����V�#0��v��S	R�g�Bp�oCP%�� �E�Aa�#�E��DDPX�D�����o�����bP�W>G�.�ݲ����t�4�| ��񦞞�{��J��MI�"���w:@Ö�#��D#ݥ}_`�0p���4�{����M���N�����=�͹ͦ�wd�esOj.�;���ἇd�t�O��"�66T��0�E�a���K:`�0��J4Æ4��1��f8&�Ws=�R�?�UTL��p����Q�_1L;��Ueo�\�7
}����	�I������������6�q�C�;�<O�zSR�:�D��ҋ5A!�C�-Ti�4s���jϚW"��tiFe�ȍ]��Z�0���?%k)|��\ �i�G����C����1��i�cm�QA��p����Z�^��>:�ct��>�=W��0�㇏�tg,ᅘY��,���@�hp��I��aG�8�&	�DD�0�0N%�g���K8pO��""x8"Q$�H�tI(N�,DDD��L
0f3


 �P �H�a"I@����H��&�pӦi�M,�0�DD�D�ı0K0K,L8X�,N���8 ����GR�,DK<p��I҄�H D(D��0O'�{�����w�z��r�����&��j��I�bF�
;�u��a��pm�04<�ʐq{�R�(��%��^���@9�$̋qaD_�y�nJh�4ev]{B�j�xox�|p�gv�G/n�v�-����'>�xY�偌x	Ƣh�|�_wx����>�9PDx�xM��шn��N�����I��5^�v��q�s}�ݾ���߿~�Us3s33wwiU������ݥW37337~ᦞ8ib&	gKH(�J4Æi��DJ���m����x��I�AF����"�(�~ö́uG�Ƣ�"�I(��](�#�*�=/�w?I�s�������֗�r}]��i9%��_ڒB	*��t�ݒ�b���Ͳ+��y���j�P��`,�=��2������)����|Kont���oQ��PXoW
�8Q0�0�Y��JN'�饗�8&{�,��bW-�)��UD��K�����]���2�@O0�����9��g�6��4���;�w���n��Z�'�����K��E� ��B_/"��h��Ll�Kђ�*�7%:��,�{����l�9����|yA�Yd)�6i�Z��D��j��k� (0�ՠ�)!�J	a�G�0�, D�4�xN�Y���@��*�����K ���Q�x �ei	B%Fjd�P�$cU7Xt�T��i���M�F7rm�%[K���UQ�����]��]-?��}�5���H��L��*ހcO��y����J%:x:Ϸ���{ʽ�!$�������������� �������B,�40�C�3�3Ea���A�q��p�88w�$��> E����<x:����|��K�A���O[����!`})w�VZ^	��E�x� �8�፨�Y�(������)b0���C���L�pm�H�U�8p�Ο>:Y��a�a�4�/C�6qV�s|���ĝ��ʪ�i2aN#�NI�g����p�uxd�R1I�Kߢ"H�DK����`�����Y���� ���q|��(][8l?{ޞ�	��Ǵ�C�z�Oa��!_����q��L��'�|8?���n���1A���ۃ �E{.@å[ld(G�o�
Q�����~�D|ClgQ�Q�ÇN�p���:[�"P�p�<'M,?����y�e��wc����J��No���wwܥ�	��z8�pPXZ:i�a��Q�2���l�zu^GiD� �<�`pP~���٥�؛V�Ҷ]�.���؏998�SN�O����.9���qCg�:EP��m��*�8�T����b=��8R�H�g��D���ȁ�K>,�<��i�!�w�q�|գǇg0���X�~,�b$�'ㆈ����ˍ��?qUQ����?{m��8o��t/��"l��p�3�����3C�s�o��	M�����%����p��$	�?a�p���%6�SS��<>!��xB⎘Z8���
��$����t<�1�S�̊�k�����[��8�JU�=h��|�{��yx��AF#M�[��x�]����|�p�=8tӇL0�ŝ��ӆ��?�>�>����U�\LH�;0�Jn��%�H:���d;���z�Q�1LDZX"
L�q�Q��U�͵a��$u�i^k�m'��*�!;�{T��lJ$���a�P�FA�R'�ƲJ��j�s��}�^<����E��Q��!�
 ���e��=\�"�|ZD��bL7/��%�z��,�{��+?-3�0�FPz[cm�QF��xw��q8���A��s�H, ,*��V}�Pz�(8�$u�|'��Tl����ͬ]���,1�é|�H�>G�1Hq�2�)A�9E��A�t��:&	"%	�,��/�1�&I�lR	]���UD&���OAh�%�ę؈d��x��`K���G������֫��"��](��d�4�$aF"Cp�!�(�!�H�aRI�@�@��?l?��$A�8�LNĈ0�Ȋflc>Xg��vI)P��g���di6�'�3��S�(:��t�e�('�?���3�3���%p� ���p��t�@�B~8h�f�Yg�5PDGb�&C�p�⪢���\�7v]�4ܙâ��v(��x�D�A�4gS<�t8x�RH�%�N�I�ET.�BQ���3qN����d�vl/���N�{�m�z<�gD�����>Q}�w[b>I���ɶpj(�A��TJ\�JR:2�4E(:%2��"�ZqJ�����nCW���g��3�|p�Ξ>0�ΉbH�BQ���ic�#�u�N�0S�%�M>UTC�?ao�T�O|p�!���y�����8OBy�߳�Z�+0�ͥ弳9Q"?��d�X��VJ�H�@�@�R> r��i�pg���+���Ҁi��DDt�{��[l�0jԜ&���;����$h�HȒ�p��ˇ*���f���\=
!30D�,��<�v,f�t��9���,åYC0��0��i��i%Q��,��@�&	�D�(�"��,�%�H��	�$�(D�IA8'�8'O0OH�$	$PPQD�AA���a�H����:@� ��%i��4�M,�L0D��Ήb`�`�%�pL(�:X�x�B��?Y	�,�"Y�DD�N�$� �DP�Ȅ���������������E�,SN���Ǧ��l��S?r3g;�«Z�$,7ge=9�����q��d��A��L�F`w^a�i\���(����.�.�/F$6��n�i���t�n�����ژ�68�by՗��Q;A<��,���X)�v��~D�-��W���ٮ3�7=�0��C&<�u+<pߩ&r뗨��=�p�F>��r=�l�u���O����.-�����!�1�=�fo��o!�~��{��x���pm+t��5�a�~���=�1����F�r�Q�(⩼��fxཉɁ����
B�WI0j�"��������8M�pȎ%s�>���P�1(�r
Z]Fݺ2M5��n��cN%�/#�ݍj:�S]��#�0`��h)݌�pЕ2B���RY%��f�nݔ�d�e.�]$F���,đ���OP��S���1��Q1�lD���T���p��EQ#�K��0�[��7�d8PP����{��T�H���֋�=�=�><M�/�\��������*�fnff���s3733www���������if�0�L4��X�"P�i�xxh�4^�~���H�!P(\D9�weD�܆�-]�WYn�ݛ3h��SvlX���U��I&��D0XrB2��Q+s��&��#q]弲�Z�N&��F�&���Gw�4��Mb"��`B�l�hY��t��dݴ�����g%Im�
Zݻu��6�-c�B���-)m�@�B�q�#���6X���a]��kc&�]���4�j+��j�RT���l�awM�s��V�#�*"�xs�UD;�z�q�g:�4h��6����+�Cqx��q�=]�\���[d����Q�K|�#,��'B�m�*A��<8V���Iҕ��

^sp�H~|�82���?���8�"H��oQ�qD.�kp��kq`�#�s@Q����A,�4Po1�}@�h���vI�v2�:�y���9���v�곇�%�~. ��0�����,KD(�0��41��%��qk)�b'��dCf	KO;:6��f�CS�9��z�$)������z9$>�b�����0&IM�ԡ��S��qp�O����.��p��D��]\|7���y���=73p�r��}�\���
d��! �	���rr�~���cS�bR�w3DN�=�CC�<6U�_�~��N<��m�\\D
�bΖQ�Na�%�"aFa�Y����MoB������UQd���J����!�����3���b�e4L�L���B0�(�y�L��Q����<\��~v�Y��y�rMn��-Z]�A��lR��\y�(�pC8�AD�ygH��Ӧ�dZ/�zp��}T�0��h��Oӧ>�t�OxMŉb%I�xӦ��[��t�"���VsfT��UTB�s�>�����?��?��p��9��)������V�a6�R2?��@�s.cb�~m��0x=C-�a�\��'��)DƿD2 ��D��R+Gg;\,'iM��yl�OK�}C�{�D�&�f0��6�������}�N����j��QT��&Z�jP}s6vԢ�� �7
�$��Ç��<|tæI�Ox�Ɲ4�P�Ǟ�?@E�H�0�%Ď��W��Ա	��{�ײi�F�0�����1
*2!q�PE
r��T; �B�.�⪢~�g���=X��vs���L�z�C���I�w��%�Z��H7��&�����̎��ߌ�����jZ�>�(U���KMS���pq"d�׮H����Х�3).�:��]<|�������Gy��l��(�p�ǲk8p����%d�M�t}17��Q��$ �z��K~�l�154�vn�K6��we��}��Ӈ�{�B��!/+F�m��:�xx�,��ŉb%Q�4�K4��#�Ic����n'���N���#Q�{���E(L�Y%�8�߸6IAh8��M8�A��RB��D	����?o�O���݀�����e9a�U79�{�KE��:��@2)9��y�"Rܸt��=;����}��f��H!O)������ibX�Fa�0��<.uP���C�5+�Bx����	�2%d�����
!s�\5�0�³��r��<���C<�(�~�C����|��$��n����-�v�2H��i��e��)������CNs.p�1$DR-@^�1��j�b��:ٲ�A�ԍ�6�(�'�p��L?%��aF0�,�ˬ��!=AH�JVo�U�:C�s�:Y��D�P^1����WL���Bǹ��{E���4�k2�����O���������\hM�iK#�ٝ"-�q�|P(��ĔY�wQ���qD���
�:�ڲ"�<$�0�����_��)���$��=i�<a���"Q�p��4�K3�6#���]r���q���;�-$X���,f(�kI����IA?V�-cLF��Sd�#�wv`m����&�=�u�K��
�I��$s��l�÷7r�<y�+1U�%��om�)�0�a�9�[a!I��x?v�M8~0d����8����td���x6�5e����n��F��0f�β"2�g��Le��"�<@�J$���3�c���h�O�4�$���0����Ϲ���4���	����v��[lvR��ӧ���8'~Ʉ<�l�Z7�����,�&8p�<|X�"Q�p��4�K.��S1��"�fS�����DR�x~3s(��џp=s�%p�3s`� �f��M66�Q����u�=l��ꑖB,d��
Q%�<fQ��D|��0Z>��M���:7ic<�Om�����Q��z�ϒ�h���"3��W��Q���Zu�ш��5J�N�,�8ic0�&��8pI A�$D�D����J0�4D��f�Y��bX�X�%�<t�"	$���$�3�Q""@�,N�Qâ"%��BD�$�(((�H ���a0�� IDD��"t��P�t�M,�L4�8`�,��&	�	bY���g��?$"'N��t�0D��:x�H8IBQ ��'8'N����7��"�9�=�S�1�������G��h=:CV�M�v
��<6i	҆��$�]���{~�y�����J��P�I����
C>s��uo�;�]3�?hڽ��?�-�WɐZ1��^��2LG.�:��;1�m�>72�^��O�r��R����]�ܙ��bݪ�$(�������G�_��>��n�A�s]6`����y�TY�AX�'�{1���6���31������fe�fn���U��������깙�����N�if�0�L4�,D�
0ᅚif�I
9l���/"���_'=?�i�1B>C	$�v�i�i�f'�B��A�:N��d��	m٪�|9Y!�K������?u��<^��i9�Ҍ�=�"f	����P��Ğ$� �m�4�4��n��3�F��͈��l��:;�)��a���L?%��aF0�M,��s�vviKE�^�7xi��Uq�=4����H9���ptah��P���2E��%���pI�Q
��p|a����*�=�GVc�'��슃
B��j=�3��V@H|}�Å)�P��zs�c82���)+ÒI���C&f�ɗa����<s�/�R�3�4�g�`���b%Q�,�K4���G�$1f�ar��x�?���bl���08r�dR��2V���N��\�.�Y��M�YOZ><�efT�W/O\�=������y�sL�����\'��w7��|�@�rn�4w�����7���d�����1��b<u�1��pa#7!IZ<5XX�P��;mi�ĸ3�H�*�y��Ff1�r�t��)��euH�Q=�Q'��8Y�cH�*��՝dPX�?���RFefX�RL��y�!�Tpc��D���cz�t�i���a��4M,K(8af�Y��2���0���2ISZ�'�W4�)���4�����	��3Ox},��d|�o�8wܴs���t�K+�:#��7�~����	"�#�ߟ^��c�Yrx>� K��Ҝ���Q/�{�����]ť�p�����E��
t�O����Ӽck�����e�Ȅ�$gW��9PI�}�7t�d�:'�Ɵ��Y���aF0�M,�̾L�S�5�Ɇ����u~U\D�xR��iD�3ن�<�~�KTġ�}ү�����Q�U[v��@�~4������.)��^s��n�6ȳp�E��p�. �;�cȃ�"��D���w�1�ѐ�]]�H�@�e(�K��z�nO�P���Uq�:XX�`�H���J$�G���?ib%	F0�M,О~�%[k�U�DHR4������;��>o�h�lgu���dih�������HI��wv��M����lI$�|$��!||���GL���T{Q�������g�N�OX����1�?T�>�6�X�Aє���$�!<Z7��z]QH3���ITh�a#�2(~9����qAD����Nt�4��~?ib%	F0�M,ӳ�Ȧ�y�μw�d����nG)Y���ț¦ZF�r(I���X*)ܒ�M��v��NNn�-���ū�n�wv[��74[)d��5����O��Z���o�=F�9�?ϓ{������ҙ���el�m]�{udpayƢ9~�5���0`�?h�����uSrv_�>��}��(����z��a�ٔ҈�3��xt�vl�M-���aތuDkl�Z�E^��pgPϏ����Nn7G��J���2��������=R������"M���~ϖ�t�9��?���	_��I:'��b"if�(J8A�G��h�=��
�FA���u��4?W?���5S��"��pNs��6�+>_?�æq��#%�m�Q�w�޸�{�B	�4������CD�<�8��uI���(�pg�x��9���_�?��?�
\��#a��u�tc7�S�w��m�������s���3�9$eB��> � gZ��p涾<�cG�rQ� ���x���O"&�i���Y��ic�$,a2��TDz�����u���83M�������J\Fy��J�Y���zy>�+�$�&	�s��~FF���6O#i8wU���p�=�D#ǈGH;��v;��
'0C������	C���Ӽ#�	$�#��@�I�@�>�eI(����:x����4�O�%p��4�K��(��m�7�6�i��5}���L����{BO�`��ߕ������B�=���|�0�;��:s8j�}1g�K�?g�Os�==O?��17��O����L+�p��MC)p��8��3xI0�����=1? q<0�FR+U%f"U�"'㥞4�tI�	Ҏ8$� �'	0����,�0D�<i���L4�OY��4��x�҉ H�""$F��D�8 ��D�:A���3���2H(0 �$I(H�(� O	�8';��Y��i�����Då	b`�X�%��#,NxO$D�8"tO'���	�#�H(�$� ��'�'D��A�=#Ȩ���d�����y%�/?+播�I�!H:p�k|�0�tÅ��m�����d�b�1�Or���v�)���N
�5�~|�?
�4�,�؇����k�szDp��oM�z�/Ԧ��P����y��<�b�nQs���5X�Ń�-m�����ɸ��kt���챈Q�Ff�y���ޯ�s�!5��Y��- ؞��|�dY��r�k(XA��QW�!�:O,�9��ho�!zk��3����y=�g���
f�\&�^\�tv&XQ2!#�r����n��W��ޜ�&���w���osk�{+lh���w��ɲER�]���fL6�vCX�8�`i�]�&��k�n�wM��\Y-��k�0�&Ä,��K"[��^�`�[�7���k��۩+2�,��D�tn�5�K�����	(�B/ƒ��5A��E����lPtm7{xkrˣ5�f�1'z�a����hk=y�ww���_�www�ww{v����V���������n����w�4�L4��4�O�%p���������{�A��P�$q	!V�u�m�vh�:��tV��vJVl�$�%]]�V�]X�K�&���*X҈�6�S�	ȳw\�l��ܮ��U�f�v�;��M[�nii(���q��Ȣ�Kv��v�Rl۪Ȑ��J�)c�-��6�ݵkm�ɹt&�%��R4�P��b���-jI4M��n2�vl�;4�4�u,��?�*�"~�����z�kM�K?�����1��~�q�X�M�ƗlE�Eri=޹���f:<��<~>�<&�����B���s�H'WeRi�`ޚ��2�?F��L-���~\��C/�h�|'�3���:qi�5FHȋ�L(Tqt��Ӄ-��zӵg c>F�N~��K,��I�f��WH�we��t�,ch�_m�4m����<Q�%����xD�(Æi�M+�曃��k�7�!G�9趝;'(���'ؐ�=.eEOH|w/�s�D���!�Y.~xt�>m�,���)=T݌cՈ��sH��������L�{�q�m�X��u�M�J�tJI:scm�R�#� ��$��y�08q�3� ��5H��U)�ע&��F}��BOǌ8X�:"ab"i�Na&x��M4�;w$����L��U\D���"Y#-4��U���C(��J(�c*�OU^WNa�08w�L�b����g��RD�����6n���A8R:}�7Ӈu&�<\gM��7!ᖠ�n�Fo�}S��с��/*��<pg��c��H�}��滥.+}`Tr9���Q��&�"&�i�D�(Æ~?����E��7yy�74^/�Um�3�h���"����#�3 ��D�߸�����XHM�!�g��J�T�ѧ$�]ckU&�M���?q{CD�|�����S=�*d���ff9�>�q �`j��d���Gs�"�&3�*�6��^ �GK4�M0�N�p�	0c�
4x~?��o�>kU(�	����,���rbA<,9M?0㭮Ƽl�ݱ�����b�F�7v��F�JW\�l��J�Ym�*��z���HeW���H�O�.�ʡ���w�p�M��k���p��#4��{�N�w�A�]︟r�g�3�����(e��eM�
�83�1Qњ��R)����4iF;����5TR��#Ş<3 ���q[��ќ\i��O8td�p;8�Gq���ѣŖh���w�3)˕�%�P_6���!�M�K-r��wƏM9�(��s��/�ӂp���Nz�ē.R���%�:p�:a�tӆ�BQ�,M,�'�5MW&�c�ȱ�u�s����"wC��rvN?��Df��>�#�y��ط	�ߢ\=�D��3p�0��8w�����qut��>�F2C����p�%<�|se�ɲ�[	Թ����Մ�C�pgFR� ��E�gM�l,�Q�3��zo���$(��h�����҇D�zYe���&�i�D�(��&�~ύD��o�ť�9l��*�"y�]�G����w��wզ��8@�YH�b�a�̱����b#���q�!�{���w�1�i����0)m?{9&���[g5pxO�#���D�pd�k��ic,gu�Gi>W����Y3Â���p��t�)Y��Y�`��t�(J0å������~� ���h� �;����N#�蘿�$H�tᙄ�Q&~�<�C��"?��l�$� �a.N�P�pF*(ey������8�V1���Aє2�m2�q�t��
Q'��%l��m$��Hc�8��|<4�%����G��I��6ό(�7g�s��p�	Uf��x�N�0D�:h�%a���4~Ą�D���A��Qke���DrE��@� �p�� �Q%H^�c:\NW`��m��%([F�e\Ҍk)g}U\D����I>H@�Dh�y肓�)0�x�숸��X�ޙ�Fg�h��߆������Zpq�~�RD�>Ds3<�0:R0�$c:4@�A婃�7s�z��pȂ:`�&R$���3��i�����"�I�2�_��dd2hNu�J�F�����(�������8�x��:p�M<`�a�M��:X�4�ݏ�d�f�W}��x!Z�Z��Uq0��|�u6�N���<|-��3Ie��|: ��"���7���YS0~0e�H��R�%�H�t�I�������(�@���'���9V%YŚ�ϳO�?��~������t��t��/�a���H2�s>�ry, f�i�q)ıDp�4��E��I�$Nq��Å	$ ��(A8"x�,�0D�<&}ȋ���'��/H�ǎi�l�h��,N�$% ���"'���'F`a����@�(((����~b<@�"P�""&	�(� D��pN��K4�DMDD�<a�D�0L,Kĳ�%xO$D�8"tO"Y���!b$H�@�$�H����Y�,NA޼�rK���d�/s�껹�a�gy��1�k3��1�#Q{Xe/ 0���u�'ƝJJ���NC�]�NA$���+�{=�б/�
�h�E(��ɂ�Ȉ ����U�`��U���=��g��\3���9�N�gd��W̐p*��|�Ak)���>�H�>�Ƿ:�|�挛��)4���p��'���n�3�+�N=�徕y�#|<�Ι��Y�N4R���sj]a��?�g��H�W���;�䧐�r�*W�O���}�e������������������7ww~�����ۻ�����x�L0�M0D�:h�%a��񦞿�� �������a���ߗ�=�HC;�ykg�'N6�zߎ.'�cj0����Op�o!�9��i'��]�����RX�m��}�����=��N��P�6�
��n0�6":���	��M�?}��5�g�f���ݗ$/�a�����#�Z,�߹3ݍ��N�a�0ᥖ"`�f�t�JO,�4(n��f�m����Γ�1�Q� gŐ���C�/N�H'���g��8kQq$��!&˥�Y�=?�O0q>?��.��~E�'s��4��s�$���%�S�>3���?y䓧�|I��je���#�ID�����1^5qB�x�#J4e��4��$ç��ŉ�"Y��4҄�:`�4�{�~������xܒ�M6ؤ��Ѳ�v�mdVn��۴���8�ݛ����,۴b�����2ºF0\OUW^e�.E�}E�m��C	���p!BC4%r�"
+T�FŚ�A���y|ӑG�O=:|C�zf�G9+���n�Z=��{��'�`����	��xzsQ,���?���9���,G%>��'t�W�?"�|#	�7����1�$cC(�g3>��DJ�����W[vڸC�t?a!�Mb<z"��Œx��<&�"%�i�M(J0æ	�M�{�����*x�N�/p�I�<�ƽ槃y��U�g)R�j4��3<6Z$�27=9^NG��q35�����QWM=<���y�-�<�"��Mù�"C���g�_���Ήy���C�4h��%�_���"G$O��/��ݍԕ������D�d>���t�81���FW�g��$K�_���A�F�A��,M0M�4ᦔ%a�񦗅ɞ� �J*h��M\Qf���Lg&tGU�:2{�Y�|���2Qc�I�738a=���y�O�y熐�&�t��fB\2_Q�8��	X�gW������U�W�D�gI��E��~8H���ω$�Z6N2������l�2�����-����(ҏ��&"%�i�M(J0æ	�M&���G�m��Cd�\��K�h������"x~��;���繧D��R�K�D����G���[9`�<yV%���X%��o�f-6 �M�FB��X0��0�~�
~�8%q=�k���{�p���j4�ao޳�:q��"S_ �$e�S��1�ޙD��G���1I��ȁ�5�D0��,�0�M8i�	Ft�<i��-��O�)�������t\�O��*�1a�A��]R��*GYҬuq�4�8$�[b9n�K��6/$�G/#vK��,)G��U�N������_a�S`zw/{�����1��*�?AL&�Y����~��0����_���� ������p�`SC�i}7��p.�����>\�.���t��@9�c��#:4���*�V�.a��-0K���`h~jҵb��տK�$����9��� ��x���P�if�h���i�M(Ҍ0�������ސ_�P[!��H9$�9��s�y�gY"p�U\~ͻ�ip���!���(L�G�9�|�UG�%��GA���хBH���U��,Q�\�@�~�=s�i�3\�Ib�^��",�Os�aޏs�^?�C(Y(�E	�t�ahd"T1q�#��哑wQ0p�Śt���"af�p�J4�:`�4ӟr��e��9��3���L=����4��u@4R4�H�H���0��A:��m��E���4��d�y�$�"�CL�"��Ȅ� 73K3[�Y�ah�ѢN�yc3{�Ŕ,�(�Hg��"�N;���hˮG�LM|�K�#���:����l���[�Jg�a��8t�0��4�J0æ	�M%�Ap�<��ULSW>�G���QR������?|�yV���ǹ*���3{��"�mk�st�9�pJ�e|F����<�/�Oq9�Hs<�����Oa��yX=�P�O���
.�2�å�D����E1@M|DǙh *��4�/��v���SJY^說�m�f͛��[�[?fx:g�kio�y����L �� $X�@�!4X����M�p��Η�"
b��j@�� �h�mȶE�����dL�h�DȶG���!�!B��d-��-,D�"h�"5�h�2ж�h��$Y,�D�"�QdYDF�(��DAd(��,E��
&�!DBȑ�DBȈ��5�h��E�DY-#[DE�DZ-��4Z$kD�b&�"h�&�h�ֈ�"h�-�dB-Ț,D��2ZD�&�i�2L�K$%�i�H���	d�[I�,���ı,H���ɥ��M,H�I��q6ᥒ�d�Y&�L��M,���%��d��	d�L�Z[F�D�Id�Y&�I2�%�Ĵ�d��&Y&��-��I,�%�I�d��Ki�Y�R%�K&D�--��I,��$���DY$�2�%�	ȴ�e��Y&��H�E�"ZD�!&I,�Y2%�	m"[H�H��"Y&�K�d�-��Ki4�l�,L��Im&�%�%��$�[I$�"[I,��Id�	��"Y"ZM-�KI,LD���D�X�[I2�%��d��im2%��m$�BD�ɑ,�-�I��%���Y"Y"[K$��&BI�4�M"ZD�,�D���H�i4��,����	dȖH���X�I���e�%��[Kd��"Zc���im,K�	m"e��&��%�2Y!-�M-��Ķ����,��m"[%�4���HKd�ii4���i2M,��-!,�Kĉm2im$�[H��%�,Kd�BX��4��&[Kd�[HKi��Be�bB[Kd��ĉ�%���Y&�%�ɥ�im"X���-�M,�,�,�g9�n����7pF֌MY6�m��i3Yf�F֙����	ɵ��ő��&-3Dě,����2f���'6���&�6ք�ȑw7G� ]@b�c�`���ֳ��"Ȉ�$YDE��8�-B�"����9E�-$Y"Y��2(�",��Ȉ��烘r�!dDY�"e�L��D�DE���s��9E�DM-�E�D[Y�ۂ&�F�$[Gp�b"-�E�s��"me��p��"dH�$YF�,��"E�D[D�ȶ���"E����"E�H�",��h��"&��""Ȉ��""�,DDE�DZ4�"E�ˍ�-E�2,�4Y,��h�YF�m�4[DDȑm"�&�h����M,��rE�DY,���"�i�ȑh�"ȑdH�D�"!dH�H�5�Z$-�"�"�h�mE��Y"�����h�D�mD�dMȚ,DD�h�,�E��E�H�h�,��Ȉ�E�H�DH���"F�-��$D[D�m�t���"h����d"E�H�dD[DѬ��""�"D�#Yж��h�m5�"�,��dDY,�DE��$YB�E��!F�h�DB�hYȈY��"!�2&�DBȐ�$k"B�mD�DE��DY��""�"""�m-A�H�$H�i"�-�E�B-��"��"�&E��,DE�"-�#[E�MDE�h�$[F���DDȶ��h�y��E���$[E�i�h���h�-�#Z&�"�$[DE��mE�����"-��["�4E�����",E��-�M�4[E�����h!Ȳ$Y-�#Z&�DE�H�$YF�2$Y���"���D�"G1�4H�-,��,�"E�DB4E�M�"E��dH�E�H��D�"�։!h�DE�k"E��dD[DE�#Y"E�"ȑm5�4Z"-�E�"Ѥu�8$Z-,����h�dHY`�"D"E�E�B�4�D�h�dH�$Z4�!�h�"ȑ�DE�dH�Dk"E�"ȶ�DE�#Y"B�DE�"���-�l��h��4X��m�"h����E��,E�,E�&�b"$[D�b!"h���
g���։��G��V��;o-�n�q����m�l��f�+f��U[:�ό��/_���>�'�g��~�~z��~l�wg�ǽ���߻�����������q�o�n�����6�����坼�S���t�z��3��x9z8p�]������;=G�8o_�Ǧ�x�zf͛7�vz~~n?~>����o����0o�G����3f��s��!,����^o�~G�?�{&?��������6�3?�r�6�=����7�֝�1�O���<f͚=��������$ug����ۆg����m���zۖ���Y��?����q��;�'I��q��ۻ������=��ǧ���\�:�̖����c���q�7g��'79�c:-����e�m�N0t�o&��ĺ,@$*�a�@&JP,> �8ܝ>���]ս^X�o�����<�X��3q6H�(��Q#l�C6�C6�`�㗵�N���y��gf��;z���,�q��|����z��7��8?�x���1o�����{�6lٸϓpi����Ѷ�]�����m���H����^����c�<N��uq��߯��}��>��v?����e��y۽���iǳf���~���o��f�c��׎ߟϴO��q�|_K����oȇ�|{��z��׍�f����lٿ��7�̶���?�L��<��9:���[���6�>�B��X�-�8c`�w\�{QYj^Mʮ7��i����,lm�������ks�u���ݼN��\gg�g���v��g\w��@����put7���g)�:WX�g��lٳq���^���_k�����1�6oq��u��mn{w���s�������>C���{3�=g93������t�f����s|�ž��7͑��s��p��~����z�ygCf͛��V���m�?۶��6n���3������'ŷ�{3���Ǳ���_��w��'�:��SN�e���oo�vvn��GtkѾ����G?n:e����m������.�����_c�v�gF����/����f��׵������gg�=�Y�m��7!��m�[���=��yy!x<� �V�w��� �ħ�����6��g�bf`��kg��H�{Y����q����7�rz�,��{�8<N���x۳��������������������#F�OS����]��BBӼ�0