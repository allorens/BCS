BZh91AY&SY,�a�w_�@qg���#� ����bI�P        �>�-UX�E�٥a#6Ҭ�2j��)+TX�i�ѵ24bM��e*��l��[h�*Q!U�Ѧ��-3��5V�V�����i��(V�l6�Z������c6�*��`) 5�kkSJ�����֍f�lL`жiF��m��i�͙f��V�ڄ  'U�Y��Zh� �]4��fc[{����J��6�����@���VŨզfY�ͦ�6٩D�a@�j�m�i�4fښlf�j�X��l�Gi���0x�P  �<�u�M	��w:�ڦV�`U�j�P7ӱ��܎��l�є6�B�dbhtۺ�]Z�d*�M��]�Y��)*hm���F��  ��� �iZ��@��M� $mh�jƁ@����Ei��oy��W�`� C��� AOm���� (��n��VSU%�����lU�*��}  yw��Uv������:=�=[h -�=὏l���N���{����zW���N�t���(��zv\� n�;��,�Z�j��6i�-����  Ͼiԃ�A�w ��Tk��z M=ήRٮ��n�Ҁ���Qڮ� (�s�������:j�p}=�:{�(�C@ot��V����-�V��i��@  ����*��w@@����(i��pR�;���  �ު��ގ  4wI�j S;�qA���c��;�T�kP�d�Z$
�Ϡ �ހ�Uf�)��]��:�(�ƴ N� (
���S�`vk�t ҭ� :�v�AB� 
��$�R#h,Э��ila��  �^�� 
:����@� iFN1� h-r�  X� Un�p� ��2�*�5@(Gw@Pv �V*�M��c��  �z ݎ K\���� kA�a@�b�T6S� ����(t3���w�:E��[2MkZ�ƀҚ�5�   �x ��` �`� ;tuP�n������ �\ h5;���ܧp�@��wkkV�4Ͷ��T���mx   � j�z� �m�j�Z�� h�.  w P"�F`� �EV��8  ��      � � ʒ�@�  @ OhaJRUM!��&F&M�{&BR��      S�MR��)� ���FhH&i&�=��4��6SM4��G�BzjJEԤ��d�d��h !�3��wN�R;���KS��_;gc4�&[�m�Y��G3L�'4�K����`���؞J*���A U�T8U z�UQ^�PN���}G�y�����9*~�*���J���<UE�BO���'� "����N����<0�F�)�\�e&09��.`s�L��S0L�e3)���2��̓.`s)�a3)�L��S09�̦e3)�L�!�L�f2���a3)��f`̦a3	�L��09�̦e3)�L�)���2��̦e3)�L˙&G2���&`s#���S09�`s��f2���&a3əL�fS2���a3)�ف�L��G09�̦`s��2�S29��e3�C0��`s�L��09��ds��29�3)���2���fd3)�L�f0���&`s�s�f\�0���e3��fG09��&i�̎e3�L��S0���as3���09��ds� �e3)�L�fS2���e�	��fS09��e3!���fC0���&d3)�L�f0���L&a3	�L�f0���&e3&d��f2��̎`s�L�fS10���e3)��f09��&f`s+�L��G09�̎ds#6`��W29���s�\�L�3+�\��́�\�f`��@�.`���0es fW0��̮es&d&W2��3�\���f29�̎`s f0�ds�\��G2���3!���̎ds+��fY��.as�\��30��̮ds#�\����as�`s���� f ́�0�`&0a�9�L�+�Ds(.eE���2��U�� 9� � �eE̪9�0"��As
� & s*�`Q� ��G0��Ef�s(.a2 L�9�2 �0��Q���Ds"`A̪9�I�ȩ�Ps
dA�*��0��ʃ�Ts*�aA�
�"fD\� f2(�@\���Ts".e� �e����0��E��s�3��L��L��09�̎ds���Rc29��.ds+�\��3 fG4��̮d�� ̮`��̮a�L��̮`�� ��\�Les�2`��29�̆`���S29�̎e3#����09�̤����O翟��{��	�����_�6����>d�l��un�7!�]z�1a�����#��M�u��pw!=�f8v��]١�J�(nY%G[6*b�5�q㊯�(^pXś��
��$��B�w�v䐲�Lee�˼����/g.�p"j�z@�5B׶S���u�x+���E�4��UF���éMX"���2����3Y����c�ԕ���&�-⫌�%���K�˚c�2
7����^mL1����]1�G=cei�8���cC���J�FZ�g	J���0�A��3�yˊ�����-ۺܔK[179�K�����s�,�;wE蘯(�f:�w%c�n�kk3쳙"ʖ��Uō��R:�j��ݖhe�����	�K[$��L��e�2��Ԣ恻�X�~�������~��n�r�n��-�2����Vc0F�%L�#f'r�Y57X�Ц��i9�nm��՗8U��}i�\Z��2�,�͏qL�%��.�S%�u�5�@l�KNV�tӎ��<F�N�i��H2��l�Lt֫����e��e��A1�Fj$I� ô�[�"2`vo3�K�Vm��&;�csh�O4sT�0Y	�Z�zx���f����k�C>���wK��}�4[�]\��F%b��]��jؼ!����)(�M��N�W��?��+E��Wt�Nd�f�r(�b�[X��؃�]�Ƣ-����V�Y��)�Btx�ٷ������(vV��j�����W�C)2���ɴR��U�9a�s�UX5��Gvh�V�\���[�Sr�D�ԭ$ؚ��.�uR�\�>.s"_Un�I�^��Y��T�6��f��D� �v��f:�R5{^OG�ɔ�*�Fvf�yc����'6Ys-��UR.m0�˕0*o�M��2�2�{v�.�h#Pnbe��	B*8F�:�"�)��6����ZM�I�KwyOl��i]�̘E�Re���ǖn�������%+�F(�B��,R�<J9v�r�7U����ߔ�a8�w2�tP��w[zγ��V-���g9g8ǃ���hڼ7�5饅E�dn�{sE��wBҮ���+��E��_��U���h�]F��R;�)��M�}o��B圆$�W����[�����pT���x��67��E�9�j��ݨ�ʽ�5̽/]Ԑ6�2�
��t��`�S���.�#M�v�,z�QK�+�s�a:�Y��2l��.75�����"����C]�����:6�n�����L�.XV��%ҹ)fޫa��\������U>6�~!v�R��f-�09&�0�e�/���f�+w�1�EJ�S��uY�:�0�T6�/��4��V��Ʀ�xJz�	b�e]x������7��A��YxR���\�z0�ٗ��]=p�u�Lۡ!2�*6��	7,�,����0Q��fLa=cGsr֛���=iѬ�n�#��'z��j���o���+:�����K�4���]CL�+f�iiݸ
6�y���2G"���he�oQZ˳�l��;׹�#/s��vm�f��[O]�#[�N��Hr�@���e?fl��0Ӹ�X�4.�uP����ۅX��Ҵ�n���$ՠo�i���^�"K�KrJ����)s�9!S�B�:֝v�g��1KM|���'b�D���+V�+6Ƥ���u�q��c��c {�*�������opa1ǃ:ݦms�3}�h˽��so�=J8մw3ke`�4���oX8u��ŗ��L6��,� ���GW�JW�]�o��Q���l�j�P�	�P�Ջ��62��[����
���_�\���j��ҍ�SX��-���e����v���V͚�H����zn�<�V�o
� ��P0��R�d#u��\��@��+=��0����7B��UnZ.�`�E�J��KvV/m����9X���a�3�kk�+��V&i�!t��0R�N��5�"���ވq��]f^T:p&�ӽ
Aq=wk,�-�����Jܒ�c:��V,�n�*��I�g�.���{!ff�ח7X���*�
��$�f�ʹx.�s^�����oJ8yhP�t�d`�b��=5'V���MnmAɊ��V��\.55Y��R�洴�-³������Hj�KE��ޢOظ��KUohb����rVT��R�6Ln�^!IIU�\�A����E�˚��*fT0��������ʷYt�֝iɂf+W�`;	�N3F�)����w��h�N���3m�W��B�kq�r��Z��<�b:E6�Ì��o��K�@��V�N���.V%�k$����JqD�ij��2���zģ�5���"���X�����sb�]���a1iݱ/Z��͒[ɖ�s��J�`ᖚ$���l�Z��ü5�/�	�E[�+�$:��F&�wҺcP���sj�el֔v�Jȥ�4M)Y�,���X�1:8�ix�c`��=� ׺)SQj�m�q]�V)��l:��P֌N�3N(ކ�6�o�5��M�3)���&�PZK-�/K[�Z��)q��S�eI��#N:���c,�VE����Q��ub,� �X�j�R�n
�ʧr@iJU�Ѳ��ݳ�V�=m��>��i<�Ԃ�rR��������3*���Yr���#5��y-)ڼ�`gjz�B��3���SpQҬUa��1�X%�YÓq�S5UӖ�����oL�a�h�]��N�)�2��@�qÏ<o��^2�*n^LY�#ʛu��ZU�fb�*V�2B���v&^7$�n=[pne`׮8[d��ŭ/�V��6%�)�-�G�W�Z5כì���֛,�o_͚�/&�z��81(��M���`H�A����%^�!YF[yc'ׁRu���-Y�0�{�5��D.f�w"͙�Ȧ�n�+fQ��'5���f�8�����Xy�p�����%=KWkٛ*�nnP&TQV�u�-�B�C��l#�iCu�VYTYYnT:Q��,
��Wn��/1��f����e&Ս{��ֶ���rPI�.�e��I��qE�~èڴЭ�����5X�htlꣽ��]r����L�%c�m�<]M[�nB$��(Bmee����շ����?wN���V����eY����qM�$"n�f��D�t���ڣQ�*�t��G#W�*z"�z�����v�N�X�K�S�
�����Pݫ�#[*�l�0�{�+(E���HD�X�`��҉TE�jl�f��3�5�Sj6�FKC0Zk����ӱ��VUk{���W�{o���{��h�X�����z���:�ꕭ�w�c93UY�7A�L�g��H�3*�[�Bh�il�N^�+��dF�Ţ�+��P�غ�W/HN���{WM��/-U�盤�
�#�M##xl[��$���WMn�gZ7��Л6��YǄ\�p�!"Z(Q�d�n���Z�����1X�e��h�Q�wK���$q׍V�)LڳF�	'կ,лW����Լ�IH�֙fa�����5V�B���&���E�UO1C!"S�SD�;��ް�Y�׶��W}t��ԂF�v�>xŏ��-Sӄ�}����
���մ4P4,��e��)�����2�dw���I#L1�i��f�pc=ڵj{���8�;�P7��w�Y�t7���o�mq��N��5��I�Eb�-]�Ř��Ϩcb'y�2�X�Lf�ωU��,����K4r�"�^�X��+[N�l'�l��X�Z"�=U�05)�ct_���5S���2����U|�H�uF�Y�-�-�*D\��d�V��x�*����Y�pFs���,�-�"e[��	�ĞYڢ7QP�V��)m�H��M˫
֧��K�q�$���:�Jm5L(�C�^�,XEr/���˳��mepz8�!ʶfeln��q93e\ER��N��Į�M��;�5���ETn�1M7�Izv	wDV�k yN�l���9��QQʂZ2�Y6qnY��̳iӻ��c����!����ɷ��Ĥ��Z�)�)Z�"�h�S;eL��Gr�[��H�J<u��o�kj���YYR]c���[ ��f�L+6Ț �jکt*K��d�Mi�e�yzwtln�m����d�Hr퍵Z`�"�nW���Q��9��ÐG4ءeT��+e%�eB�L���դTd���Q��ic�;mn�[�J	B�ͬ�q4��Y�D����/%[�ƃ�Fa�,P��ͭ%t��[g6���5d�UL6Y:ijĮ2��S��"�`1��N�ٽ�E�M�al�Z�/O���(�N�i�N������a{-M*"�Pؓ�kIu����ò���23��(ީLR�+e�*\�vTF�4$FsI)��Z��۹�b�+���#y�������t��p��ȉ���Uzݴ��w��R:���,��#07z�G%k�)��e����aTi�1���@�+Ae^c���I�k0�˲�R�Sx1c���\C5���q=yi�XSV��j_A�@؂�3��;I�6r����&�ݘ�P2��J"�Onགྷ��`��3
f�������1�ڣ�osk%e�a�#�'%ث�P���~�B�5����BVN�r/m����O�%��qVa�D�Q��xvnEJ{��㸙��"�Kd��р����R1N��/3n����el��݉�� ���5N��n5Y���6*X��"-j�H0�6�ٍ��:sP�v�D��>.�Y{aVf�a�	�L�p9��V5
Swq��&"ɤo<�ͳ��d�{�TpKX4֍�Ƙ��E`V�n�F��8i����85mӭ�䬈0�����s
V�BMb��/*yɅe�E����,ʼ%���L���fR�5�	T��O�a.��� �6nܪC.����ZC*��Sf�(�G���5�5M]jWR�-b�̒R���9�C�ăک���9�%PFⶮ�.��T12��$LP�%�����ہd�--X�42��S���ǵJ�ՕX�X<����uGf��Bî�>�Y�1�9i���א�n�s'�An�y(6)ՓA՝P��+\Lä�ڽ/mk8�t�Śȅ��&��NS�������Vڶ��b��:.���`��/C6̷�#X���A�1�`����(;��Uh�sn�m�ٶ�c���=�	g(�e:Z]�:��L�i!m'�X�j��e鍕d�yǙ�;J�O�5� X�5Zј�c�;4��>N�E�C!4M���R�ym�p����W�%(TtLySP�aKyY��87cH�S�zT��V��k-ي���"�|^�X��dT��(�)���eb�������!T4�T-y��s+Nehd�a �@��]Wo�.�5cq�W����${��O^j�c*���+vP��#�	Nn��V�M*�"�qk��̨���x��G�B�LaG��Q�ɍy�A�̈U�kv�4��/ElxL����R
E�u�wj�hg����@�ts�
�c�yUs���-l�̩�Wog��Q��;�[ǁ��m���e�4�]�U����u��.�ڢY�/3G�;��-R�]2-h"jV�ӚP7�ZcӤ�5,D#zL������(<Ɇ�sI70���{V�6�q�T�n�
�+uQD�Y(��=T�Ӭ$Ys/MYT�;Q[�l�eu+a��2[ʆ���H��P����b�u��`g&��֖�=����A�.��z%6�����lZ�-��šU�FMN_�L�$Yٓvkn��R�Xza��0�̶���4��[R�Z����y�|S5�q�-ټ�6�1�U�1��3�F0���J�ӧuu�1���=�Y�X�Զ�	�z���ms}%-�����tom^�N�,��"�gv�x��M,�N�y��f�����/t*d�3+*�����1�Y�l̰�${R"��q!Ό,	��Rh�EbpMو�e���	_u;����5�8�4�';W)[lPkE�
.��e�/u�{�x�Y��I���,�hK�ź��l�%��ް�kI�y	��2����v���R���\ �B�樑�]Vj�jΆB��ƚ����L���{e+a���}V��]��:o3N�4V%�T(��C-Q/ODk�Lb��M��/,X-ӛ��ٙK[�4�*n+���e+�B2^e�Um"%gmQҵ�r���Au�s��l,V�c��*Gp�t��W[�L�hnY��*�ηV�Ȕ��EUn;�:�m�Q�S��j��L17nf��r�����d�i��������gI�h�^���>[T��*��*��q��Jd��6L��)Z����8��I�F��u�tF�� A�A�Fh	���`�nY		�҄3ҕ�IRJ��f�l[��,�;����v0JbN�^2u�էw��oAt�XHͬ�T�ͽ�24ia		;OMY#� An��h�D�Oao5a��z�\R&u���}/rr��F���ڮ�Lڧq��d���W&H��g���ǻ�NTW/9S�z]<[[]ֲ�J�')7_:}�\�	���K]�,Q��&�h��wq�(�p���&ؤ�]��9c��ڸ85��uv򻵆�<���|I(�Wv�\s��sxBW�n0铫���1�V�$V�ꐎ�Sծ�1��6ѻ���3�T�Nu]����v-�Kp$����6�O\L��|����h���,�X�˼����l�(����i��^+���=:H,#kn/���O�I�ع�4������i��w����	����j��Z��ܲ��1�Y�V�7
�#(1X�$&^�����i��� ������m��eH��'��w�k�^��c����͜�9%G[fޜ�Qk(1T;�Zt]B��Pa@��&�hWZZC�d���uh�n�#ge&�KL���H�b�f��U�Q
���f�Kt�ܧt.�J,;�2Ϳwe�WGg��7�U��~~�v��l��{���}��������/}�i��ſ���}�����������I$��8�.�-��$�H�I$�I*I33$�d�He����-P�'�L�Y���X18(Vգ��,�X`�;U�Ex�
57�ԜT�n�sL�� �Ob���S34s����wQ�+{0���Um*�[�l�S�1�w��[��#J���os�r�CfL��27u�u�u���s���9�p,V+�탤�+��}V��ӛ��}�ܻ�w;"���CI)ڹΨ�v�R�����M:�	ӗ�����&�S���Ey�[כBm���A|�9��͇l��R�H����IUۙ�F5� ҖUE�P7ѓY�8�q�lC��M�v�쑜���.�lE���� gMWw�!�������Vu�x���*��[*zy��w��:͖� ���Z�]�{ʹ=���9�)d���˂�=�D�C]x�h����z��h��R<.�cvy�n���m�K*>�P���d���|r��H�l�NS6hR��OvT�4js��]v#�(���y:���9Lj�t���f����*ѱ[O&Y}�����FK\@����K�J�o��Bm�L����tg�����zV�`�Q5��^S����lrT6���ח4�c3�M���P�ѽtE̋&�p��ɼ9u��z��e%n��XD��+����Po �,�os�e>�1�-\��������=�X<$}T6nx�f��r��u&��8F�+t����z���%97��v��s�u�Z�w]�ou3�󩩗c�x=� �Œn�Q�����滛�$�h���;Sޥ4T<����ȽA:_!%�ch�����|�]�j�VG��b��Wv�\�}���]�2Q��[sVt�����0�����g{V���j���F����u."���'�
���s�B�W��:PΫ��.�P[Sk��� �h�QgS��uH�����bE�n�ņ�d��Κ��*���{n�b��=/�ky�W_����fιy��i�g:�h��,�خ��ID�1a�ښ��K��]�(m�l�=>Ğ��a�v�n�Xz�C'mm��D�8�Y7���Ҝ�d(ZhmKÇ�|Y�蚚�B���P�O�3��J�w���+�eȼ[bz[�=��i�ZVQ}�e�ytʬ�4j�pl�s�Y1w]M�0�.�3B�-�+e�]Ʌ�9���f榍M���J،�o@�<&��:���jd8��Tz�v�Ob�BB0��Vy=�av�GY�I���봦���D�t[5�ŕ)HCL'��C�w|e A�˥�78���B��iʌ���,i9I�M]�������<2�CN�'/wI|���uz@(t�ќM���E9�8�i=�;a6s0�7;Gh�ҳ��scn�h˄���[���P6�hLX���1Z��m���7x��א�f�_�}(d��s;��h�yӶѢ�wO(_+����p��1:���Q�s���Z�o
'7/	+A׈�2��ò��'�$�o
GN���H�
���W��RQ��7)�wur\&�a
7oz��J�Y�<g)=4M��Y���6A��9Vi{�"�jLA1}�͙]�� "��ت�⦝�w���gn��M����n!��~NQ����O,9�ܧ�ٗ+��Bڍ��ǐd��J�^nj��ESM��\�P���1=ڻ�w���Qo�[:�3�I��ɭ<E5�5���s�ޞSf����كgvܡlek�<�5��h�1��i9A���Ʋ����ŬN8fɺ,�K�_}5d�q==�Y.hM�����u��TE�T��+����bnvVR�4�r�Ǆ��dк���THq�mʐ�wK	z��3��驭�y`Ɠ�|Q��Σ���Z�@�0���T�@-��"��s$XK��9�[ʮ7K�{�sWl��ht��"g�}�Yv�6��L�4�m�7�۬�|�kD�n��+�pT�<�\;{f�u��k�S�}��[�Ҳ�G����6�]&+2�������	{�rRU����Z9Y���׽r��x��q콢���xꇜ�yÎ�Z>#;��e^�q�XFU�\��'sS��Vqv���ht]b�V�t���cK��s��G\�[sw�p��E^�;J��B�xhB�Ƴ�={P�]]7]����SOa�+6�w6#�56F�I�'*ҁ�Y�)��\���vQ�3^c�2��\.�$v����u⽅�4�XS�g��go"�:�Ix�j�s �3,[˺��m�s$�T�8ruV��[�`�=4�I乵�b�W#	�ō�Uܚ�Y��hKz��7�������ܹ��T�3�5�N�؍���O��ˢ�v�UنQ�{ʵ� P�!x�fP�P�]��cׁ#,}��l�#�#���y�U��>�2�ʶ���t���'oG�믥��8�"����:�G#����i�w�������0e�!XF�_
��.;֕rW�t'���D7�g�Q(���@�:�w5vP�1���a�P[�;�i��Z�C[nF_c�)�wgn-1���QG-��7�V����B"|�{���s(޼kv�����}Lu�=/$6]��gK�r���j���#�Wl%�m��������ser5��۠2��r��"0�%���^>=�N>�W��N�/f�^h˿�[N����+^����k���W����ˊNLng�� ����鴷�]:��4f^����-�p݋k�_r��y��K_j��].�r@f��&U
ͮB�
�^����b��7�J:v1kV��D�4�ͺnЕaf�a�165�uq��Kx�oc�c���ΣD:����4�!��)�L�W{�q	טMg�m3iE�A[a�۫k�aM�Cen��v.6Zus~�x5�΢8��؜<�A�ut�pL��!-�U{G!sHѰ���[��[���R¹���;��<W;E��1�;�Xxo,��ݼ:�#+ۊ�����X.�C��*[;�j#������8�S^v1��b=��u�$o�*��TT�kXx�Z��}^��B:��)�Ȭ�Xd���
jr5��s�5��֖��{a}��>yA�oyՍ��Ɏt�o9�'{����C{���u�+'�5.��c��R�Iԯ�,.`�wX��-u3fd����8T�=�2��s����x�Ś���#i���F$��`�O6x򬒌����!��+L�w[5J�qrwf�Z7��t�RI%V֌�ȁO�<�Vع�gV��e+�ʀԜx����ܬ�M#��P�Wp�`}|�L3h^T�P�u�qs��e�;R�J�Ǜ�5�9��r^T�����SK&�ԖVp�{����t�����87b�pe����*�wk��2u����9]��2ݼ�E�10���X����{��b�{ϲm��R�#��3n��V�V��(�hH�`F�*����y�Y��{t���H]0[.�Y4mJ�n�����=�q]��i��fsoᙏ\[[d��o.zfvi+����ȁ�md}�#��5܀դ��9b��ѹN�ɕ�Ӧ˅rQp@��IWh}u&��H-`m����gq�ggen�P�[W��3���h���3 ��J��z�\ފ5��5�6(�j-��ZŽ�nv��+�²���S���.���	��)���+A��N��H�[�i�i�w{����o��1<�f޴���ֺ��D��³[Q=y|r�V~\-"�2й���l�;�D�	a�{n�!�-�2��T��n0e(�){N�&v���D���s7��h��g����}OpLq�;�����7xXq�꛻aoX�4��s)ge��b����K�G&����W�[ss͙er�*�Ӊh�KEzy�;�<)V�xw8,a�9��i-n��٥z��)8�ِ�C�3wf-�k��},VR,�)N�;�n��h+	Rx����r�:���T9)����3�a��5�U�Um��Y.�v�w�Z�ic��e��+9H�b�][Z\;��í�`���{�[qc#��MK�cx��k�],��ڬ�v؍�W�'1��6ܫ�!�ͫ��8&#�ڬ�{J����4����]L�_f�[��%�]��E��2�5�q�H#!��s�4���������f.uf&pl�˝�M�4��S|~�f��0[[h��DRp�f�64��6kDx�2���6:F(���V��!3wv㘥JK����ෙ��+X�_cd:�ɥw�$�yi�ݹ�c&���{�j�sƍ��S��Cp��8u�)����lvx��-�r1�z�OS0h�_jl����j�s&�֑��1b�m�L㛖��IQ���Ӝ�|8��h�њ_G�G����CW1��s`�;���@�{A׳�fh8��U�Θ2s�K�R"�>��"*��z��C�u�5��):��c]����s�ƻ2`
&�^okso���ѫ�=I��*�°���󧒶�i��:�/�����O_m�¬�\3���L]�F���7�V��IW�4�G�v���Y�v���q�F��bU��z�oZ�=���sjE��ˊ��*�I�g5�]�ܤ�>l�T-wd$S�2u�bMPo0+-Tm��u�Z]�kaZ�n��B%���sxsrk6ϥ��.ZhM�E��2��y�٠�Y�����'_v$逕��t��(�VQSZKj'W���16�
�ٳ�t5��s�M�6��Eh�R�θ��p������M�5��(�Pm]�7��V'n.�3Ӄ�Z+oR����J�sf�|���K�#n$a������JR��}(�Ɩ��=�,��6
��фM�K0���;�]�R׎���P)yv�Z�

��:;3�q�n��S�Z�f�*���ڣ3��$�V6Dw��ʔ�b�X�Y/E<Y��m�]��_
�J������7�x,�n[�ò4�Ղv�X\ݗ�mR��h�or\�oO$�&\b�i�ٵ�u}��vZ������,�	��2����>����o�^%��o9UL�n��P�of�|�Gu��2Π�֠�p�X��PTa�/��mi���]me��{q��T��kg'uGiL5��LǑe��ނҶ�{�-��S��o�Lښͼ��&��Pl}�p����g��@�Ŋ�\�k���g����;�厳�Q��:�V��K4fK�wK6�S�u��T��n����g%ҢT��ܥ�Z��N�7-q=���X�(�ZԦ_v�����QE;/[71�m��[��L�`痽؏r����\1�n�2Mt�J��$��f�go�B��ɯb`��	U�A���.R'a
�}6�tV�ܙ6����K�tw;uɕ�]�[�΂��tjD��kSm�3�ql:�����f��{��D��[��/��Z4���.����vQ 1�w�h��a5L⼳C2N���櫨ග������=��S;��9:�5�����;_-sJ��y��7��M>R�ţ5��l�(0��Gj���C}�����W�"	�ַ��i�{P$e��JT�D5�3}T��}�>��н�%��,���|ZT(�DvͶU��T�lp6E�a���X��$=��J�,��d��w��:���+�n�շ��B�];2+VX��:ƅ��\!��_�v���o\K����cs���Ҥ�I�֝����u/r�y��G�+4�{s%�W��!dF���Apì\�U�]Tk��F�2;\�h��܈m��z��qmΫ�:%�c�/m�����E�=�Y<a���P��-٪�o�P&V5GR�9+J�3M�N���+;B�r�V̷���W��
����Ugn3�s��������������8�	J(��ݮ���v�DWV�/�����%df��q��DjZ��rb᠜���c��Uʗj�WD�a����fG|#���9S�)������3����8]A0�m<U;�
<�}tV��rZSyR�Zwb�5�QՍ$�}��N]c�o�=6"q&���W�#q�n��x%q����d\���cm�V�cp�,��mӼ�Y�	�^�I������s�p���y�M��7+qq�f-	F�Z�"h��6��̗9nJ��S*�ŋ�����AjR��c�w\wu����OB��Q��{w-��\��(ܢ��U�]�h�C����_Uc/&qӏ���6k��Xb��Mʇ�\|�!���y��u�v�JLto=�֨�雍+��}u���LW�Gx��0�qD�w������ɗ�mu����Bvl9�d�˽��J���!Iux�G##w�rI$�L�=�i����� ޙK�<��)�N��E� D0���Q!1K��e� KB���?R��(�CNe0*3`9F�bR,��0��.D��ti��++�i��P�U�Iq�0C�B�J�	D�)N��|C\C��u	�HZ0����n�x�2Li�m)�!�O�ہ���R�RFBSr�q��
(���,�)�3�T�j��(*hL�%9
�@�hD}�Q5^L�Y�.�`�al6d�HH�f��l �(��M�T��'k$�
�H%v��?\�����g�ƋR�d�щ���Th4�/���b7I����Yl�T ��mI%P-3��I��T�1(x�44�*1E8R2�.y4)QR\1�CH�l]�&��h� 6W�AI8X	�;cE P.ڞ�T�5T�����&��"J�GI)�Q�$12�ͺ�Yh"���f�������=�(�����y,� �m�#�u�'��u`���PQQ����O�e���������Z_��M!��H�2Lg6V���w�uDFn=�����|a���0K�Cx�\.�6�ŭ��*ͦ�9k�vxu������"Ug��� �d�������Vi%� �,}W�@�R�gJ��^�#+j=�_a�̄:ÃK_T�6r�R�ޭ��|GZk_>TӮ�7)��u4�̼ԙ�m�xJ�ĳ�>������}P*�wW\�*T�BM3r�j��:���~�Rn�MUj&�a��õ��u��&�Ѥ�%$̔�7rƼ�u`	�D,r��U�q+�6	�l�ec�I����;�C����뺼.O�s���m��]��[��2L�'F�Ѽ�ڝ���N�������dp�9���N��R"e=ՂC't� &e���V�e+l�j���.}��Y2P�cO0i��c��^�!eg�L;r�z�,83�`{�W�a{�ZظJ�Қ��*���[�*ܮ� 
�Onw�S&�el7qp*ݞyK"�����h�Yx1�ՠzޓ�1�s�8�{��{���P��U����fXQf]�m�H��W�UJ>��J�3;p�V�.r�g���3��Vm�x&cM�_Ul� N�4��N=�W..��v����-�:��l&���ە�::=��>ӽ�[���q�J���)u�
ܬg�=zÁkU�@y�E���F^��
�$̪D�f�q��=~=z�z=z��^�z����z��ׯ^�z����ׯ^�z����ׯ^�z����=z��ׯ_ǯ^�z��ׯ^��^�x��ׯ^��z��ׯ^�z�=z��ׯ^�z���ׯ�^�z���ׯ^�=z��ׯ�^�z����=z�^�z��z��ׯ^�^�sׯ^�z���ׯ�^�sׯ^�z���z�9�ףׯ^�z��ׯG�^�z��ׯ^�g�^�z������ׯ^�z��ףׯ^�z��ׯG�^�z��ׯ^�^����]+Q�5�W)�)�"P40ڣ3Z��ٓ{k9l����d�]ԷgG3b���Sc��gFn�`c��x��usdԱ�:6��M*�b���s)R �<$�ѝ6��/ �iX �Gù��D���]1R��+(����ñK�V�x�e�nJ���6��C;�_��d^�6�"n��Y�����*^e�m6HZr��{9��;3QljU��=���fr�Q�<Z�iy-��b!��m��w�	\���b�j��][�4���1
\w��L��{1*�,s�V�@�}����T�4�Ndz��qͺW2T��-��ʛ+d�#��[�=r�l�
d�vt�#*Ý-�3`X�휲�7J�gM�'fPV��gEY|��fQ뤠��\:��2�ス?�|���ד�WS���'L:���$�E�E�H3M�)�u^��1ץ];*ҷy�H]<�%�f>U�f��q�1&����A:B�9�H��S7���W��Y<����T8fѻa������UC�:�'���������NbMF���)�^��/Cy*��s�S����V�:�v6��o�J�/7��f����s����=y�f����C,M @���[���1�(����vI������-wv��=�ѷ���U1����b�a�C|��W�k͛2��Æ\�ݖYe�̲�/_^�z���ׯ^�}z��ׯ�^�z���ׯ^�=z���ׯ^�x��ׯ^��^�ׯ^�z������=z���ׯ_�^�sׯ^�z��z=z��ׯ^�z�z��ׯ^�z���z��ׯ^�~=�z��ׯ_ׯ\��ׯ_�z���׬��ׯ^�z��=z��ׯ�^�ׯ�^�ׯ�ǯ^�z���ׯ_^�z���ׯ^�|z��ׯ^��^�x��ׯ^��z��ׯ^�z�=z��ׯ^�|�{���w���Hq�7�N���o����uкܮň=\c�ۮ,��AH��^�g�]q#hV�F��q?7:��c���ы^Tk+����M�y�dx�X��aqÃq�7�;� ut{�6�f^F�}����G.�^[OQvtθr �:O���j2z��w�U���hCoR�Q�-\�M�+��oMnV*=�OR+48��ͽ����1t��Ad���;f/9��ֳ�6��t�N&��Ef	�SG-,t
�KӦ�`��ԕ1�z���j��t��4��G��)����Ul�ڧ�l��X���=�Jv��3ze�F��:bt0�L���B�sJ�2�Y�fc��
rJ�*�`��xk2�x]��\%jߞ/Mo��d�7[��$w������`+H�%í�nvj�.���	�־����i�܇v���.5�(ᣊ�9v(�}��so��T�,V��;����@rqբ,HU>��A�b���!��d\���;E4��4*� ��(*5��E^��d�S0��마���I�]��Ψ(��e��wL�����RɚK�c�݂v�,��9�C�®��^8K����)���5@�b+$X�L�WO�T�(݀�\]����$�=��ns��y�H-ܛ��3�� ���O���Pt��:}V�lIlÙ:fc�\}yH�j�զ�&M3��甚��mdb��m��B�[r�9����r��Ԕ�5S�k�L 63���1u;sAt�aaݖ&�:Y���5.�e�X_'�4�p8R���wܻ�n��Z%���ݘ�N�=�cW[�7W�66������:�r�5��p���K��Kl�Y�G�7Գ6�{o��R��RFT���ٮ(n�3h;U�P��+��vAX�;�I��2�Fy
�hCL�2Wi�eT�9݃����c��ٷ�q���fn�%m�b�د��y���I���n�l��9r��JYǉ�yn����- e�{��!�J��+�ڽ��My�Uu�b�w��V򂄣Sn�'J��v!B��VW;-G��G�@���-��3y���͊�8��>��g:�U{���t \���[5���s�3B�H��y�{%UD�q�}����2l)���;�J6T9��.���aB����n�;w��3�'��"(����Bv3s0��%��� �����ٽ�)�؈l�N܋��)o�t��R�H�fd�	�C�B��I�d�C��^<�Uv�/d䮄�ڸ��\0e-FY��T<k�_;��X��7!Ⴢ籇ZX|����y�	��r������l�I��"���M��ӯ�:��&�=�<�G}2	���2Yd�;��b7R6�6��6���7���4�	��e���G_��g-j�]���WdLBZwG�9�i�7C����*gs�Es�9 �-5{�(a�d���7�6�cj+l���bm�������T��|����Z	��%&�(������y��ٻ�r���I���h��fs�ں���40l�Zn�T��p��|M%�󐃩�n7ײ>�v�P�&��`���-��!� ��m��Т��2�6��v�`�Yڜ��@�P����h�b��ɣ0Q�sD�cR���ox�]���Wu�5�ؕ��p6�Gw�<g�hRG�i)�C�����o_a����v�.�A2t+�yXU�mK�y�;���k[���aHa�gj�(V����dv�V�h���e�acҺ�M�}�r��8S:��G��>8w�tw�w����f)�t{�Nt�ȑ��\��f��hv�ۜ���*�Oj�AM��TQ[�p����{;ʲy#X� ]�M�����*�u��%s{i$�P����4��sm�6����%>��/��J6�(L���w����˖�g���;��6)L�IU��GU��t����	�"�Q��b�mHĒӺ�6�e*M�Zgm�m��q�����;��u��[��pu8����uݕC��M��H��'��"����Wiq+��|n��x�	ݹ�Z9���  [{��N�Eܝ�s��v͚�����7�u�T��bݕ����-�E�öӶ�W#s�\CO`H�T�Q�sn�u �Q6��%:R��ά�����Ie�4
d ����7x{J�UtʅܟT����cYmn䯶�;��8m»p�滐$i��p�o6�g�A<��gsl�wz�b*8�G|�M�MDkS�)*�m`�4�6lŵI��3!�oos�����Yge���bS�vH-�j)˺���"�	y(�ue�m1t���v�>Y��u�,�s���sj�i��:�2�Y�3�Uf%ux�� !&<@��J�vntTZ^��[�K�2eY���Be1�ͽ`%ݬ�%7[ou���ݪq�ks�:�?F<%`�ƹ۽�d@4�P�R��>����l��u���顊jy�f۝�);Q�ɝ�3Ej�k*����s-Ǽ%W�Y�]Mdif���<�p䱺�{�1��XV�|�^���T��!��T�vMCqS�s�.�K	���	�B
M6�*��аN�Փa[J�OdG��)]i�{V��jõ�"S��+.ɗtsp��P��}���HWl�V x��)]t�H2֛��Tl����K
 ����V�cW�,�n�4\r�����L���u��_e`���S;�rb�Kj�S�:_إ�����,��/��SS���ٴ[�囷[�f�YdJ���b�"t�Ӫ�	�sa���e	��`w][�A��
� ��N��k��6����56ﶔG����6+�]P�΃3�]c�@��Ʃ4�Y#�]v�� �R�:��Ohn7�1��u%��[W���k6ω�d2w�g��Tʣ�p�.��-��V�̓��4��nT��s7p'��n�!�M�aT28Y��U�GrƾCkc�Q9��}xn�[�u����L�&R����\�d�v����q=�h]�K�8�����L�`�܋̫�xL�u��;��u��uI)�j^r��sB�%��j��&v�@5b��{���w"�Xt�õGx��į�Tz�GbNܤB�r]�'�HN�;�B�R�v��WB�&-�@��Φ��q�+E��ؐ�c&��󺱝bw2nN��B�\�A�&�!a�����7a��1�V�G��y��{M	����U�=Z��&m�%2�rL"��N�g����\�v��>����F��m5ȋE��r��u�]o��-��/(�Xb�c��j����yX��K��]���}v�E���k]{Ż���E������+@ӊ�c��s���G}��mYQ���I�;*��ǔ�n4���evA���A�n�+wlk}.�=�^wP\l飜e�2��M��Y�9�r�곬L.�;S.Z��e,!�b��D8�}ǰM��l���#ͳֵ�B&�^1 ��4�l��C1]��""���Z/�����ղ	 �J��T�z<�du�4e7��K�.nqefι�����0H����74�C��TA�DՃ�ï-e
�%���Vԙ��z,��(���]y7�M�n+���ۑR̍�wYC�5^��z�� wF|��f۩9#Cx��]e��	�7�ga�fܠ�VZ,Z͕��!g1f���|^!>Z�D9��>|stDt�O��d3������e��[ؒ+lSt0m[�6����]n�'�N�y�{�A��6s90�RQ���Ά�p���ͮۚ��w��X�f+ʰB#峖�Y��s�Y�z��܌;�Y˰��t�IqVrH�s:��.X+����e�Ôa�'M�ĝ����71�;T���o$���R}vd�FXI�z ʘ�Q|-m9��:t�4�u���d.�bp�#A���Bi�Q���ks��x\}����ԉ�X�[�_M�
42š��f��h�蔽��n���C�r:�ҏC���ռ8��G�%�I�ͼ�����3Y�r-9ؑٻ����D�(1��rx$Z	�N�EU]}v�H���w�����,���}$����+��݈�B���|�N��KQ�<L����M%��G�«�o�ϙ�Ô��j!�	���{ɽR���w����	��Jt�y�G@J��b}�����ݘ�(�JUÝ�窍�����@��� �6E� Jn>�2i(3�ڶ;�����M��=꾕��R���]M�Q� M��,@��{�g���&��(m�YΠU��	=q��X*��X/�=�H���8���n����6�Ӿ\x�])�)Dk���gb�wq�/���,��o�`��ŭ����"8�����L��N�s��qA`H��%�^YUu�rsB��Y�w'f�G6�������`�l����Q���7����Q�I�F�Ruؾ��g,�o�/r�1;N�ε��;���`9�B�~�}��ch�}�	ո�u���8�o�>��'z�aJ^)���Ob��%gH�i�����}��݊,f].���3^���B\��}vۮ7Ȕ�:����y|tx�N���ҋ�	ڪ�U'nα��9|���:T6�G��,U�H�ozt:���GA�Z����c��[X�Ao��7N����ʫ]�>��e�Lvz9jJ�;݈�1���Om!4"�jV�A\�ǄV�C�,6��H����yb��޵�W��p����ʵ>����:\��a���5}�ѱr�Ԣ�sY��;H��Ð�Η+��;�j��p��lf�̍����2�m:�Nb^M*�z�b���#4�عl���<�2;�-̮�:v�S{�Z��\�{w��!K�T�|
]�\�״o
i�� kZ |��`똾+)WK�V��^]g�^��a��\�Ι������G5}f\"���E*c�MQMQ�Ѭ\-qs0V��d�p.����k݇�ث�b��x�p���i�T�
:{S��y�v��-��nfq�Ŷ��dh�i*5]$��$=�+��N��à-���-ә\RuA����<���gQ���<9%A�����O����!ұy����}�ۭ��l�7�,�ا�쌴%T�Q��f�jx�#�jDWu=�iG��Р�x��r�����v�-�+#�e���V�ƒ~�p��'�G�	�R}sn�-ײ�y����L�o�,o>o����urS`�i�k����ws�z�Se�"���2�&�]κ`�B���HP�:jv�V�xV����`�u�w_��x�����A�������z��_7�$����������'f(��D^N[	���Qx�)��J�>kѰX)"J,W�	�Mk?�����7/�:p����[;��M�]��-U�?MT�[�d�j��oV����V5Ne<��`持�b@�7k����{��{��_iw֧d5��x��ViK�$�Z��me�ZP{�U!�2/�(��ĊST�-׶7�dh͜�ѝ�T�e�VrM5��NO3kL{�2l+��m��A9���T����r(�8�u�܍X������l��T��ɬóxg>U&�6�(Sn�Nl���.�v�H��Jؾ1�**ʧ��oz�<�V�X+6L
�^_nhh��4����h���Bl��Ëk{��*c�L�9a�9�B�X���oD�������q|Б���m[�tO2j�fld\����q�,m��u8d�eݨ�b�
9z��%N�J��zM�9���\�l�K���WN���d��(��"����)乎��6��rB���q���6�(&6�jhEѐÎ
��j�ӷ��ͮe�5�p���H�ɌfAh�v@£�v��8�T��ɜ��PvEݕ$��h���7�;�x��|�"��w��N�@���q�:��@C���}�K[��^�o���-ykY�y�r�Jl8D:u� �^%���t{p�����{��(e�;Yϵ���2�]�$��4�zG��lA>�ۋГ!&Z
6ʌ�I2A2G#	��m4����b�izF�JH"�%�
m��2da&��0J,���<ܹ��q?�*���"`�����iű�4j6�N��T��9����f88�4lݻ.Ye�FYe�Ynݻv�޽~|����j��-�r��AEQT�k11AU�5EDQ5UU�*���f��,���,��-۷nݻ.��?q����ض�b��5�)���
j��f ��L[&j�6�QLPlk��1��&�-�TV��l��6���U3$�T�cF�j"/@٪[�-f�6w�9�Z
J*-[Nزm��Em����F'cI%^lAMq�9���X�+Z�i"	��m��j��^llj"j-X��+a��"""I����Φ����Dh�ZqLTQ[h�b!��$�W1��mf*-��ULz��sh��9�b���5Q��s�RQ͝�X3��b��kW-r6����.�n9��TK�Y-�P`�����*�w���2փ[����r��B7���ce�ֶ�e�G�	�@ؤ��K���br��ս�*`媡�L槺��gt{���ےg;j��K��f;}�gmcwYl�D1� ��u(Fd�2��x��	Ϯ����eUX_�ܬ}�N߹��>0��t�w�lN�x����ei�/O�@\�������:�w4zMA�>�=��z�t�x�SՂ��̞���˯h��^�#�@�$�����&�O�c�#�`*���=��z�{�����O|�q��yo��o���w���K(-�n��у��C�T��>�ܧ��U�{2!ҽ�p���}��5�La�G)�IN~/=:�g���XR�ٷJ�=^�>�����c=pU�̝�b��u��Mώ��Ӷ��%�L3�6@a�*R��I]�V�2�<������b��.�=3ķ��s{_x�����2y���56�J����f��ﮈ����j���H��s='o}�y��T�u��,�q��=Og�9�0�Y�����.2���m�'(���D喽�����I��Um�;��,>3-½GQ-a�̇�m�bÕ�i��V����l�C��Bc8HkY���M鍪JzD�&f�>��ż�@���h���r�o�m�֩t_ʰ]rSs�N1�;*K�m�ǯ�a����vɝYݼ�F2Ʊ^Z(h��ܾ+'jw0d��=�V��s�%��OT�΅�)+�VCW�F��eL����3{�Vq��l����Vwz7�g���R�N��M��o��h��-�VB���%�������^�������ď�9��+��.��Uq��ܙ��b׋ί�̹癝Gpup�>{��c~����E��FNW�������gW/rVQ>w�HP��tp2� Z���_�D�8z>�>�|_�{l�C|�{�w-�f��O��в�_�x�\�>�wu� H�R9����{3�[X}7�r���|�՚��"��4�1�&��'~���ް2����Tۯ_;�W��͙Y'���n������!�p�c�ג��j���zC�9�o8�bFC����{ڶ�꫾
2�j<��K�;�o�6�w���2vϻ�����{i���B��N2P��iO�r�s].�δ��Ù�7l]v�'Kj�AbL��4h���a�-��hv�E���[`F�V{���3V��5<ڈO˲����[\q�nƾ��>�B�P2�U����u�v�"vt������������F�gK��~�5�%3U�&�3��x�N��I�޷��s���2����z���B�����]zeP�<�q��}7���������G͕Ƣh�ܽ�������{�T@ޣ��r�~ݲ=�a)�Kf��߼��g��]W�E.�.��E����ݗ��ՙ���>�3� C&N�V�6�^��<� �L��IO��6�琍w�=s�>��o�ʝ��!��5(rg�7}����i��S��1T�ԎU1=c�3�vӢ���l����=g��P��Յ�j���4}T6�ٲT�r\U��*�G�~��z�B׾^{��$�~tז|0��%�iP'��㭞��������P��P�S���d��jm��c�"��rk�=�{|xt��캊o���1��{�]^�6oh���_��D�H=�mU��o�Rz��o�jGzmzx��f;�ɜm{�o�~�B�mmr;Yhn=�[D��u�AՅS����z)�B��
�n�}�>_.���8�0�A��f�L�]�ѷ0��r���"��q)��[�������y�{���i��H&�����O����1C�8�5���ީ�^���[�um%��a�sA���[��-f�M���g�����7W����Žtv8�&N�^��vq�YS��Q��w`U>J�O�^^Uz�ﱖ}���vCi&����<�l� =��uY��7U�\�����}*�� ��+4@���oA'Cq�6;�T�k�y]k8�m4��3��e�ͪ� �m���C0�cyz�:f��<M�3��|OK�^�l�ݓ������������n�T�,�os<��ꭋo3�Ё�l�=�k�ӝ���$����h�}����]>˦�y���<��I�s�wJ|_�
�������o�)x�ߟL/g]�Γۤ���˞p^��c'��)�{ϡ�N��>�}=�N�kʨ�Um>�y��X}w��)�5���R�^�W��5�Z��W���%b�}K����{"�d��Bv8`z��]͉�������u��R�Nqˇ�re���]�9�̑����[M�5�T�/y�Oa+����ԽH��)BWW����k��ǦT�eR8;p-�)��3i�e��V�@F�$��:c�-嫛]���d=�̭A��ke�T�� pHa,��A�b�>����J�����vaH�Ci2���S+�4��rm�{�ߒ�����6t�T���;� �י�I���~�峮e,�R�b��M����oO��*'�W���+lP�@�a��{�Gw4�F}�O�07�c�ы�O�՜t`�?z�4u���k݇�jd|��_�%M��}Oҗ.����{`�=�"������pO���|�^yym�ϳ��{8�M�@��ͫ�a5^�KQ�ӓ#Od�&���T�8G3d�֗��l�o�|I=&���m�m�e>�Kpv0�o�����|�v{&�z�]z��*w��׫���zzz�I��d�0.Ϥ���{�����X쇭�(��#��k�������{�����O�fW�a+���t� ?=�H��T�s u�rv}6+`�k
��'�Y�����i��:gI0x��&Ns��OO�g��0��-��M�!�r��!�r�iP9D$��I��z���V�.^w"����|����Eniٕ+��X�W����80�u{���D˩��Y�W��ѡ�(.��P�eH�xo:l=b9�䰖��n�U���G]±%�i͇�
�~��>����1���8����wSR�@룴O?�@�[g��;�6O�v�	�U�+\��ߜ|S)��^��{n�Λ�b���ϥ�����x��ＦWm��Nt��5`���p���$0.vl���������E#�z=�ʹ3��趍��q^̋7kŧ�d����S���*S�)y|F4#��5{�����w�\��?rz���{;��G��k�X~�Z�|�:��{���� ��7L�k�׹?O{�NK_��{�Ql��t?u3W4[��r= h��k�[��i�ꪮ�{+�e,'��8dm!�t˿<����8F���O݃�.�6vu��|�{{�;=��C%=߽�����RE���Y<2��|7��I������w�kF�o��Ϸ�Vs`���P�U�H��7�2O[tO��U_Xx}Q���ge��k�:�|�Pe`��0Z����D��������A��7����*�\$#��FW�;�/l�u�/�5��I��;�fm޹j�4B	fQ)�ё���o�^s��w
�N�����V�^[N9&�-�Rf�A���<�8s/R8mj�jR�>�Y�K��]��Z��e�}]TIH'8ӎ?g���sG���4;���߬U�[�>pD��.�}7���;�g4I�x��I�����1�M3���_y���^���]�kݺ��}�{y��Ǵ<e�	6��$� lx�h
}/l��ӱS��rK�^�cE�1y���LJ;'��2����ޞW7�M���M�l�o����ԛ����s��X9�R���2�lt����ؑ�GM�=�Kn��x�K>O�#��.G��J�}|�{u��yk���>���o�}/l�̧���;K��+y���9��ո��p6*Ry��yB�����}�͑��ڳy9�{�o��:�55E��nr�%�ԧT*�9����R<:J�c��|�.2���R�#ųE)3�ռ_Z����Oq3�F+u���1}��RD�Lb5=*�sIQH���M��U���gw4�}����.���M�lY�	;�����'xmj�/���[�U����2ھ�
�Q~�n|�����6�}g���:�F�4*����q�M��f��x����i]�v�9w�`k��:�Ӆ����stW>�ي�R�7��]��CU�/����g��c4oΟX�{[V���d�IS)�yUo�4gT�񗵻+��aQ��Ժ���ʈ�N��կy��󘾟X����h��V�;�AǗ�M�ݝ�X�3�>ݛz��tD^]��*kVH������w--�2��<1,��?���U̞���-�7L�������>��Բ]]���>���,����E��x����l}�vS�_����xz_�.�"���Cx�{Α�����LB��+��8��hA5꣹�6i�ձ��"�����;�{�$��dGh�Y�=�w<�[�G9�	�.I���o+9ļ��X�Y]g��ty�|����%e	^ϵ:E������z{��Ӻ"�[��E��%���g�v����
�(������3����{�^6��27������>�o*���ƪݼ��+�_U�t/ϫ&7�e��|=7�D^LV�'d �����n�q&�g�C����Q�V^-�&��	���>�wyX�4�A�F�V��En&��X{�m������9�P��F�Ҝ�-D���齢e+�vd�;�\M֍i]���֯��FWr�S��"�P%���Z���ٓ;��� ����Giؐ:虢{��i��-�̪���p�mm52����(�o_b�>0r�}�{��L�5����l�Æl 6���0��/��/J{td��Ft52'�?>������}V��e��9���YW��j��}�a ����|���&w�W�{�Oއ����3��������ܨ��#��,���+j&}��fH�=V�K��3���L���A�6�>�TG��
�OQ�߹����Yݻw�qg��D���V׽��~��(`�b�=`�9x>�E_O{�V*�sok�N۾e��'Olqn��;����"�������}cjɃ����8��?f=�E�����t�ܽ�=����<p�T��?����g*�4Ay��6{�Kͨ��\^�Q�����O�Dm�ߠ]W��NgRu�U'�����w�{P�²�42��_�$��پ�=f���/O�۷J���V'O�\����p��\�n�a�_h��VɯuQ�Y�^0���C���
G ��Zͮ���͜j�%��A���>����q>(�o�1�$_�2T���O5�H����_�W���ι~l�txcC˥���xX�=�:��Ͻ7r��ɳ��0y�'�^��B��3+�G�r�������{9��d˺��e7ޡ7����FW�������-�d�e���Ov�w_�@6�v�Ji{��^11Ꮲ�?L���2��{ƌ�O{��ɑ]!W��W��L��⏚w�{�/"v9%��|�̛�C��̫��G�^�J^����f�ZӍ�ޥr8�6Mq]�~�~��7����_I�]�zf׋׉{���z�yeёھ�\C��M�*����5��PU�Ok0�V��TȤ~^�{���Dʄx���'rs��%��:��?P#F�7��]G<��9�����/y�wp�'���=����9���N5Q�I�p���K
�2�b0����L-���g�E�ř�Pf�~�i�� �o�WA�=-|;��(o�<���*8s�� �4S���0���$��y��6����k��5�)�'y����.@t��t%OWU�̄�G��s뙜)A���ޮ��J%v� 8��
ɗMÔ��Ucnc Eق�Q�f��<�kbޕj�2�7k���%\�]KU�̹;q�^�E�	�h�p�S��S[����w�*P���m�L[�.���%oN0E�'�gt�n�Y�V�ñ���]k(�'j��\�p!��׺KT c8ݩ�=�okN���]�i��w��'P��h6���۽wbWiwl�Ԅ�X��m��Y�d�H5��o16��Zġ+�&�j	�)�4��c3g����p9�R�f��K���"�E��j��ܬ� ͠���'���lA�2l2�;�r�HGb�ڶXw�n�ab!�9���)���lF�),b��^45�u��)��L����Fe��]w����ND�;�1����1j�j�v�ř�d�#�s��LKi�����*��g,d�CuJ���GKu�O��JqwѼ����n��7j-S7B�V��$K5����ЃW�R��h֜��{\��9t�ӹ̼jÔ�mk��A��
��j��k�ٸ��s'c׶`�X��5I9:�W]XҥP'{bOb�P���
@�X��{2>��k1�,� �v}�9P�6S0�rW���Y��p���s�Ԥ�Rp��j�v)��zԏg�t�X�5p�ϪI�t�Bq��j��;�����u�Oeu�4�S�oQ����c��,�Oe��EN�xQ�X�}��!ð�W�Ldn��-a�7tѐ1[�W|q�M�ٲ�3w�a��<xAtl���׫0eߎK�N�j��wk^������|��fd�r�w���D�(�5��"�]� �A.ݕ���]9�<�,��?����'�`]ZCS�]��Y���F"<��GSbY���mM�k͸���`��N�g1�W.�:��[Һ�w��6H�#hQҺ�YLF��u;r�G�����M1R�fN�i��ږu��u�*C2��\�ҭA�le���M
���C��;��bu��˭��[K���xw��i��k[��P;v��ۦ�;�5a��tk%�V*C�s]�vf���W�e΂�0#11��kVn�Y����c5_t޳�-�d�1ܜd��P�$�{�Bʛ��l�kTŊ�u@�l�l�n`ިi����Nb��ɬ��t�2=�[��N�MU���s�#��D�4���n�)��*m�S[�ޙ��١JA�W)�5�o��ru.�v��� b�!oM���7��c�!���w�%�R�r7��lіc���Qf�H�Y��:��QgY�ܻYt곶�����Z�y�V�!�51u~��2���铂�.�|?�)"D,��m��v��s[Q�jmV���m-��VV�X�V���ч;lS�L&5�m�勚��gk���||}_���?��ףׯ^�|||||z������q�1��7�(9͌b�0�sZ���`óV�q�x��Hgy��&���^r&�ƞ7.��Dm�}�+M:h�gg9eӦ]:aӧN��|||z����?�\F�Xض	�9v"֜�S�"��*���<g�0cQ����O��5sp.DIf��6��*��mZ�N,D��;�s���Pk-�j3�,E\6L�kb�k#E�l�#�-DcM��0�Mj+��SVw�3p-Q�6�3�X&(*�cV�KW%�W�\9�(������U�Z͍���lQQj? تH�0j)�(��`1M�y.���ԑ1W6lZj�xl�6(�lQm��[��QF�EEMTUDEQ��U;�-�z���m��4�� ���(���
�a�EU[`�lDd6�TMX؈�Km��W1�k�jj�t�J��-��8������lUD�TQ�&����$m�-5�Ӎbh���Ӝ<أ�9m�:PE�EKED��r��V�5k?�x���X^_]2,��r�|	�G3��.�P���xf�ݎ�Cum�Yo5�@w^94(ʰ}�>o?���Ѻv4�����7�Q~�x`(��㺃t��Y~q��{�D�&�Fw���b������?��´=_��
n��#���@��!�=Kսݡ�>�Ρ~|� �8�B�R]���i�f�Xw/
b��O,�}�\���V�2� !Xk�??�t#f���??˭F�Ȫf�e6���'�F i��7;?�[
�j�W��{�^~{�J{�"�\ ��=a�yp=<�`�	ȡ�f�!5��Y����1%�{���x��Q 3�|�S�4Xml& ��O���gu��=���}>xe��b ��S�Cd�nT�����C�L[ ��T�4�:[��T���#��ړ0i�CU�;�.2�Q%����'6�J�gs��4��}�4J�<�P~�.��s�X]"�P	*Ml�����ȸu]�YM���T�!7Wowv��q�� ��8��кa |VG0G#a�{��|��' �n�J��,9����&��溫`��j޼��=��}A��<���|�o�>�׻>��; �TA1i�g�G�����>?�3�5�6����i>b��L[������}l>��C�����^�@m����ُ�'��i)#�
�Vџ`q�1�[ho�~�cQ�#L	�3�ǜ*��V��*9�H;GS}f=�S"���2p�')��h́�H�/M�d;'r���,��.u�pT��f��5Y7s����"�Tx�k��o[oc�)t�ח���O?����s��F�q���^�^ޅoA�:~q%Z�/��S]�y����&D��
�? 3�Y%<��㢪r ���{�W��p;�F����;�}w�:�b�pZC���h��j�Q��U�;�w;V�n�Hh�<��w|����è�5��=A�����c�F���U
?h~g���f]��n����=��m����^��^���lGf���A	��
��y���� �zT`:j�;��D4*��ps9��F������ glG���>ǘqm�̟<�;pЊ�3E�vb��q���m2���jn�ݫ"���lE'�r������cm��8��/�}S���6<�thCz�a'g��,�B�����]{�X���o��4S�`K���;����p0Mǧ�r�����j�̓D\(��W�܇�c,8� ž��R3���8ʆ@�t��zw,��|�>c���5�������H{����J�-�����5D���8�P�t�@���;��n�; ���K�3%t�����o7�C�qp��m�����O��{�|���Х~�I�5y?���y�_'7b|�T~��j;�mk��U�\J3�S�z��|�r\�&l�6�e�V�;A�Yu�k�X�t4��}±SU�u��[9�d暛;��I�V��ҵZ{Cwjh}j�Jm�wN��e�x���Pln��{����i�˝��lrC����S��"<}�?��{�ޑngh��z�``��<�������^��X�������@7�s���#"���I��HQ�:毲��-�G7�5n=0C_ŭ�WN7�'Ƹr����j5�4�s�{�Rd�0�[]��]�j�i��=�����H+�g�e<7��@� �D9	�ϖ��v�����;y���/�n����=�1��>ZkX��q���\������� |�������)�pB���q݌��W���w���i7��,�\�zJ�i�HN;���><�8|m���rN{��:{q�4<�n)3��xןÚ�Л�R~3�(�ؓ�.�*�xPY�̪º�ݾ�58{���Jr���Zـ'!9��J��ژ>����N[�`k��_�-Y�:㬿J���K�Z���v�[c6M֤yc>V����Cŧ�D�l0G��x��mi��k󧑹E��v�S� ��u䡚v�mS��:�u����N����'����?~�/U��
�{��?p���?�i�>��#'����N�ge�gP}�&F��Xbo	C�^q��p�f]����5�l��s˸'CDay���T[#O"��e�i��ŵ��ڒ�;C�v@z6�?��u�~�Vz>��y�Ȩ�l��9�o�\���ieWU柺�;m��=&*�^��5Ja��2��$ᾭr�(��t��%�f_!O8��>�;8�6X*6g3���������?Ǡ������3��jxF!��4�2� �d��xc���2�Yp��|�4aԍn�=����V��#1�<5s��Ұ����c�Zy���� !���@�П������{C�?'"�k^�;-�
��7����b�1�R%�Pd�_�������u���{0�*�z�r8�Q�)���A���AҞ�����ΐ/�#xRm�2+F|%:8��rXU:v,�����C�OKy����{Z�=[�S[;_��8��������S�A�,f��9�����c�M�=�>7�a0-P��o�v�5����$8���'ʘ'�"���P�1[T�7/x9���;zjo<!�.���^GfV�c(�E�7E2o$�0��qOw0�z�� �Ɉ0\�*iN�;�����=�q��({�C_��[����==�e�xZ5):��g�]~�	�\�+;���Nɦ�������ץ{�{�vhe!6������Ȯ��P⫰�T_�"��XJ kڤ��A8�yxbMP6��1^+�=�����C]�@	���c@LIuC�K���vJ�����]�t<)�d�����J�N{6��3����'�L~�1wD�3$����j+�O&Ɗ�(o��]���s�T�>��ρ�	X��IUǏ��#r�3B���-�w�&�9���Qa.��b�.�h�bX�� �Ep��:�s���ݛ�/�|>?�Ϸ�q�;ϸG��K/SӸ\8��k,:=í~���-l�ɭaD��{��{i�/{�t��u7aC�_A�m����ʈ]��{���?ԣM��=�w�| �&����z����}^�Sv3�$gӮK�r]�k�15��k�tg�c��:Op����4MS�ȳ�x�m�C�G�6��J~�^=%��D�LP���D[��!��ý���;�[K�ۼ�e!oԭm�gC�����+k�|u�n�gs�\����i�A}���=�!��fŹ�\�ٓ܇�S:���'�����y87hmy��xk6�~�5}%�t��H��,b��v�m�C�o%������L�b9��a4�22����s��[Hԕ3e��n����t�������x������c6���_��a�+������ǧ�N0F��W��ݝ�������uV��C۸ 
b�)A�����(�0=�������^-���0<0�p���,k.He�3sU����8��=%���p�	�d����`�R��q��^�t��>������n]���,�Rk�޶7�E��?�.x)�y�az���j�jN��4��av���a�B���K�Ipw}��Og`4-�c�*�T�\��0�����]YF���+	�iR�ݶ��-K���f�n�]���v�>��yy{���|=����Y�R,m��
�äfH#�>��qާN����|��N��7H�I'��#�y�^��U8:���<�.���ԇ���Za)fT&c>���R;$É�i.�h��`��-��˛�A��w���ʛ����ޛ�h;Q�3߇��9�/���л!��?5�0+�-�S�n[���Q{�a��kt� Z~J��]WT�U]�]OY\������*�3L$ў`#��#�#��7磐���S�9��W�yRf�eo��7[S{�H�6���l������!k��i=Xs��C����H쟍L��S[j�H��̸��W������M{��2�z�y2l��X�羨�j��ф$�!��w�'�`w��h����͝(x�sܺ�n}�q/XŁD�>f��9�^ɏsz������aba��v�+� ��̙k�xn�|=��}����?*���ߠ{���~Nf�Q"�g���r˯M�<dm>-�o'�������X4��W�4���0��fHl|��B	���r]���Z
���#D�L���G��wfz�I���D��A��|g�|�KR��A�,�����Q�A	��̫�j(U��P_,�Ջ,���]݊�����=�x��ٗ��v�N��ۙ���8m�1�|�.��'�{\voor�� ެ+
�X��R�I2e�.6�/h�!YblПL���Ԯʋ:�n��x�J�U=�<�l\��/|׾Bu�?+Ǐ>�� z�M�B�T��\"6����t8��o��9����L�N>4��X�p�Xd���]�(#��0Y�W��13�H[E���d��Vj�(zK�!���U�!�QW(5�����8ʆ@�t��N�`���R2R�����f���${�킅 �zn���0B|k`е�N���z��@eE���x3g'w�m���%�^#�����[�DD�J�M��-�E�נ���p�ħGؕ
6%Rf�S.��.�1"�B,��#���b����N����Au�'�=sH ���Ι'�9�N�#B�z��UYj�N��/�����t�z= �4ä�a�e"�Y���s�Gu*Ls�����s��oRC�]��K^���O��/JF��
�����F4�r�L9��C&�f�;̎�=9�ڥq7J�bxR[ɩ(�E�`sN"���f���]�Z�;^}���Vz:^j�}���> �U�n�o�Ə��ˈ[k���ܖ�rW<�*zJ9�r�v��|�|>�ChPV��ZL�/ߠ��+��3�{��"�OR�\��B�x8ⴕE�ΎeO�ư-t�����,���=�C5B�@jQ_�R���>Y�8��@���1L��֥����aL��s�����LƧ�S�!�<�ž9j)`V�8dm�}2<��j��N�f�=���67����fg�V)gg;4�|1�5r�Gc�{e����\�;��U}K�������z��  fֻ��8��[_0tɜ'�905�wxZ�u�_���}��K�0|�,��5,J1U��;�qfTL��;�8aA�3������	�e���-�C�*>��Dy?U���z�4�6��9���.��21�����>x~��W�CxB`�x�6߮a�'T7dm��q�uP+�~𓑕ۻ��{sb�+1ޮ�T3v�x��`$lk�����חt��v���,�3�t���w&k�<uᎠU3�|�E���T}��˱��ɽ����gРN�z�Src;*6j��6��N "�%��q�fBOW�Ar����g�o�鳦.gRl�ZC��f\��������g�<D��<�����$E�ҏE��OT�m*<��cB�ХiQ�>h����ةl�W���$�|=��ކ�}����G�y��P����A>`0��Q�?}�mCƖ~�X�@��7�}]�����3Z[��Zw !�=�	��];�X�o4��xh@�ҜI|�	��ju�����4L�LCݪ´��pjj@c��r���c)*.���W��8J�������d����v���J���(|ꖨ#q�j(cDu�Q_�!&J�'o;y_�L�i٠�	�l�B{TO��L����p���٢���SG�,�*Q��rIld�t,/���L�����(1�'קS�J���΋��Z�'����g�^��ǂ�@� ((���9���4}�05�̤��M��tS$�����=�Ek���b#S�W���j۾��Uyy��,/}�3�!�	��]�a�ݑE�F�C�Y7�tCi0i�Pw����⪛6�iC���p�4��ʦn�;������҇^�4K�o='���7�����2��l���U_�}׏�M�!��]�dx>=�b���"9�	�N��,P:v����VGs�oc���Ц��2�EXgC����o@��2���s �����l:<'�0k�LKZ��-l��t%蝶y�y5�yX�i1T�-Q�+�`}sӍ~���hvB�:xW�ߒ��B
{�L1~gfj�3Z��sS��έ�y�͚ݚ�#�z1���k��OO��gӯD�1�`���GE������Yʖ���E�s�����!��_1�B]����6��3�9��_��g���]a��{��h�X��?J�O��3����vj�����GM*)����X��{��%����2�,��d�d/y���s�;���b=�j衡�~�1�?|�O�w����tn�P��X*�!*����1��f`R37svǡ������$[j�;��q��z���RC"K��G��_Hj�*�,q��
y�<H�HGf-��ջ�����O�%b�Y�T'��q6��:�n�=è��3�K�,����h�z�N\���/�g
��{�ｾ~�x���T) )P��i�)��)ij�)(��y�x"%a6�U!�.[� !�G����]&t�D�����~O��ic^~|ql�RT͓��d���Dv.C�^C_tSd	9A�`O��/�"��hqma�w����	!']m�j���=�鹬��S�l��zǲ�Ak&b�Q��Ҍ��ŉ2��3��0�(#Kʼ!��3�zyY�������LY�j��8�	�d�#�#B���6;�>6�_��	�[�W&r�uP��=˷oyh����\t9a���A�y����>1)Յ�)�JSStvH��/��u�Ȋ��H��r�Q��^�~!���`��#�@�z�}�d����F�v/;�"����Ȥ�=�Z�=��*<ۈ{K�d/c�.2<�aD��	��1���ho 〦X��&���-N=O��
�m~�s�~g�g�lxt5&���`y��4l�Q���AK_��_o�nt���G~����;�ڐ��֌���
]'�rx:�����>ZQ�Ѩw�r֏˿h���|�\Xbf��^�r�O��2�Sm&���
~b�ɷ�+�Aj�#b�ٶF�!���@���N�xB��S�7����8�b+���yl&2,�^V8��#G3}N������w�z��[{���=K���zʭl���]8���4���j]/��>�|��������~����ְ'aO,HK��i��v+�C���h�`���l�����u���7kL�7v/(���s�_[��bW�L;vò���޹s��ڪS͠�@���jdMN��N� ޭo���ci�1�u�\9^7[�m���W�.{2�H�vZg����N<��x�N�,&�ĵ.�;V��z���r	֍.kp��֑�Mަ��nap��}*�9�����R��"QỈJǪ����㻉t��95�oc�]cU^�͛S�;���ú�3hӪH!�%03S�n�\색�{G]�
�	�9��=.��ET)�����7GEVꛦ�N�':�sq�{V���m��E��٨��fr��ܙަՅ�E� dk�m	Ϯ*�%ty���b@5v�]Sü�y�_�]�0���`�����Zͫ<��冠��]��n»��=4f-���ٝs�ш��E�}n�s�ٷ.Bf^�<U3�������t�6W,���}�,�Չ�C�+U�f�@wTZ_K�h�<`�&��y��7�egSb���ӽN�Y��.g:a�շ1�m��WN�d5��뺣����q̦:�0`+YUu�E�)#Q��/1�\�e�Yy?�K3�#1y'��L���$;"�?T6�g�ΰ��.�+{���8j�
5�+�e�HS��(�EV0m��쾾�Ow��]V�&���i�.Ig����Y�[>�k;MDC�о�u[̹���Sw:	3�(��βޓ6�s5�4���x�m�QCK;K�*�4���K�N,Z�MIx*�il����p7C��6��nܧ����%h�����IswV��-��u�����?�gbc��XCu��[q'
V>�x�x��SN_Q�][�ۦ��M�daŴh讼�B`�sJ��9��шˮy;�y0>��Y����S��c���B:ō���D�G�ͫ�n۴M�zb���8VVS�8QG��W_aVi]�F�8��71�r��Tu����h��(lu}2��#a�j^��чZ#���GE����f�X�һ�u�	�o��ko,�د�W)qM�!�*:��&f��=�����m�u����]07��e�#��q��ޙ��\pb����3y����`���8�e���dn�g>0���R�������=�ε��{f�J�(�U6������34>�'�v,����e�+*c@G}@[�Ef����:���:���NQ:!��H/
V^�_��X�j��cj�W���#�> d������c�z��o�'�%}wW0����&���z���*�y��AWۢ�����*$�!�PI D���1�	f�ŕT���&UC%���a�I�%/S'�R���nD�(����"�d�"H�����8R�)<�b��A$�|	 !u��Ѧ��Tb�j��lMUF�-E�Y�"&�����>?�ׯ����ׯ�?_���������~���Q~�QV�8ӂ"��)"j"/�h�����H��V�LTS�j�׏ٗfYe���,�˧f�۷t��]�O�TEQDTST�6�jj*���V�r������j*j�*#F��Q1�����D3QPET�ETD�LL�UTQQD�5EDSDZpSQUUW�AQQQ$DUT���UQS�b���U1sa�رALASDSD�QEM%:ãAT�UQ4�ѳ�����;%sj����1l�����X��$� ��v|C���9�TTL�m�$T)�j��-�QTQ$i���l�5�ֈ�98��*���d����s�j���4UDD7�i9��E�	���[F���*(���lt���B����4��,�i�?�=az�nEk_32��P�t��M�W>)�@����4���P���,��dɂ�:�+�@C�Q���P)�g�xQ��T�F�Av6��kL걫�32�.��G;��]cЗd�ޑ��Z�bK��e�OG�H5@s������J���PWeu���CŘ0��x�	�;&��̜��B6�l��y_����������9�H�&92�w��j�����S�/k�w9�L��0-10�A����wW�k��L�wA�+Y�O;��;�ې�f,���i�����
w�h�29�&
sM��Fl�7o7K�x��r壧��nd�Vg���[Pm�di����oP�x5�RO���'�`+v~��v>o���dm��<y�ux�+	΄C��1b�mH�0Y���"<�О���=`������R��\�lgg����7� �{+/
}.%��)w��s��SU��ю�Ƭ��ܹ,�\�`_�v�R�����6���D㌠&'^S�9g���>�q������(ʤ؝�c{F0��͞�n��9�6���Sֲ����~���|��4��;%73s�I�9�N���j�+��Y݈{�s�6�/
�>�D�v_�0����C�L9��F��'�7��E�g��֦�S9VW2!��Z�v�"7�&ː3Y��H��]�u�0>�&%@��$Ɔn>�Y�xF�{v`J*]�]�;ܐ`�ܭ��9G8bs�֨��bcz֧;�JI�6�L�t*�&6�������5*��4X��x�o��% Çv��V�Z�(���S|ujή�-���4���)=��lA�o�|���, �@�!?7����{;mN쯲oj���$<o�%�F��eU�^���'8�<9�o@ӱZ����]��A���]F�jS���;���x�|�	yO�&D��[¨vI疠r�'�	Ic\����'��|w��3(�����iC��`��" (/^u�uo�$�%I`����i���l������_����[�uV���y��R�b���B�~:������z1���k��x8�1Mў��'I��1g���z�+x�qxoʋo�^ú���8�|�� ?����sS�$nQa�^�J�rn�)R�^^VFw@#ե��3j�����­�!<X�>��d����
��,����N��d���;yzi��8���L��Hz��۽Z�/@�f�z&�ՏhR���B��T�^�'��A��0�U�[=9���y���EAc�7i�G�"���HD?G#.��ʽ�6�ƶ1;ݏ:�R��x�*�����=��͎��%�e.|��zj����a`b@k�#��r�r5��t��ab��;TW��� �
�S�1��qv�uu���b�s�M�)�RXz�wo���ׅv	P��a�X����/3'5/\����Cu�I�f�Pq�I�!�M<�-T��Z˥ά�s��˼g��8^R��uW�u����}�p�j�jը�3��o}�:>�;_*���_h[B
��-���g(�&�[�%!c�>�,��J�0��6Ő�ƭ�[}Ӑ�����䁌'�1P��
�p�Ȝ~6�|����}�
ۇ�."y��ټ�k�n�1��)���H��o��&��=�/�k.y�f
TQ�)^��E��-|<����!5q�w��,Y�i0����p�>�8�0	*ofb�j�O�g�@��������r۞�zY�齾�N C�^q^y�@����L��ĲN�7G�L�R�w����x=�Ͻ*#���"�:2�;����p/����sЗA��H��&GdQt��E�7E2�-5�`Ӗ+��S�ۊ%4�i;xk��0mt�X��ŤB��0u�M$��zNٝ��p)(�I�l�e�������܅h��<�שּׂĻł�O�	�8�������&$��Û@:v��*���W�͚�u׹�{K�R렏�X[ ����������o�M�\]sz:��L&�Aid������5�����q�`���Γ��j� +�cus������ØO�}�3��;��`_�uj0�-ꚟ�ϤO�o�Z�Y1�'J�oDo�^8�G8@Cc��,�k��fBWe�;���G�F� ;ܯj�,�<;G
]�ٲ���&Ί����Y�)ց9�*�W�kF�L"��<�낏;rT8qi?ϩNMP�Z�P)]��c[�|L�%��_�gf�o��M��:�l��נL�'�Z|���g�38�`w�Ld]tYd�l�]��|G�6S�-���۟g�h3m{�Rp�<zK�$@;@����7�@_���~y����<�2t����5�A!R_{��ڄW��}��{�J�u�����	z$@"GN�a�6�6�v���#��%���K�@g��sKHd�ȗ�I�w�����۹���>~���\�ֺ�����|�=߱���/`ʽ�Zfj�0,>id�{{�;0=�������-�.csj�W!��f+��m8�`�R�����[����g��
I�|���g��G�9�{.ze-4�����:},��~�:E	��c<���aVD	Fq��|��>ǘz��x(ݘ�.�C�H��=�����q�v@� E�kA�.(�:F%���5ߢ;��9���C �T1 2�>̕׽�{ ���|�OtJq�0XO�X��p8�uI/O�)�I��bS��S*IRknz:2��ƅ�M��ޜ�=�Q���ê�@�
�fl��R�m��� ���=�a�'��$��)9QWz��ޖ�MY�/���V��PRU���{�T�k��T�U�4&�̵;?Ls��J���3�e�h#;wOb U*�w�C7��$l��(�/��L��|,�S*�}9iJp|W6I+���ML��(܋+)S�g�ׂ���In�	O2Co��W�J���� '<x�������Z��d=\\@i�vV�MA��<�����M����#�K�:�n�d����Y�8��{9��_9�A���RiH�0�z<�����~`��،qa�]k��{����9��$<]ᱼ�wO5��%�Y#YK�J;����I�w5�!����K��U(p&�t���f�<Y���/�ԊnoP��ƻ�ִɷ�Q�5R�lקv`7�%+�.�ݐ73�H{CC����z��E'��0Xu�����N�e݂s�E(����l��v�=�Y�x�w`!f�\6�����C�az�2|�/M���ɁLbXi"�1:r��e��FT?C�^|�4c߹���xg�b ��ߦ�YEn�m~�3��Ch��|�a�fydfg=���ϼ���q������-�h;��4\sO�a'W�-���p�� 	�f��f�^����qCx���s�x��A���`޷���|�<���t�w��B5�2�WmV����N�+3��R�~k�haQ��sl��,�Z����Ƶ����*�@�t����k�u�e��u��]�)�鳎�G\}[؜S�ٿ;U7��6��@�J6����n�)T}�{R�6iHΝ�3c`����K}�׻�|���mԞ}x��R�}��D�r������P���p�wʣ���L���P��}s$U;�����]���Z�j *mi�7����7�u0C?�~B9<�����O���4���$7�k^��^��ʼ5�����vj�laS���!㏭�b�g�,���ʆ״Dۍ�1%����{u��$4��1IՌF�+�j��|�]v>VV"Ө{��,�rq��C���x!7��N�.5�vBnm���2O�&ø��5QX�|��AsO��|+��I8����a#�-�tc{$�v&f,r<�5�5R	�S�C�
���({I�k3�X��-�2+^�&�������摹
 ��r����ɊŸ��u��C�:�1V�7*y8	�d]ctӈ���zi��NⴠM��1��#�YA�#^��_駷��y�q���Կ7O�Ȟ��M�]�y���O`%\�ԩ�HO�"&�GBӛ+7z��;�:T0t�1 ���y.���`h�a'\]�U�����+���ڗŊ���k{W�������0�B���y��C����?!��ƽ1�w�ZI�OH�
/]34Y\�icW�:����/���j9���� hG,K �p~%{ᯠ���8���u�wJ0��{^d�Uc�E����.En�3�O���V����J����5���_�g�D��iz����$m���ّ���Q��js�����E�P�z���޾�z���["Y۩4���Z	�����[B�Շm���m�86�%u��>�γ�����{�G����z=�  ���)vr���~�״`N׉����e���O���みH��a	�1�;^�=p�Qc&𨹋ݣ��x�3롦�є�I�/D�0�L@8�����[As�.�����Ι�"1�_:��W�x���5�LQt�����3�oE��ݐ�?�!���T5�1��^�C�M�W���f�r,�8~�H(?�xGo&e�lf3�Pf3�W�Kߊ��B�O�iv��O�s��9�u�9��>$/���(֙�}5?(S ��Pr�>dJx`�@t-�{yJ�6=��f/�{xr
�/�/�b�P3v6�3��o�L��rtk���~]F���{d�&5`�G'&��������#׸ 
b��BcV�
Or�V���f=[կM0�}gh�Ųi�K[�$d�C�L7.i��V���$��x�C��R��Ij&%:J�T-�ŷ��k�;y4�ۼ��j��۪R��[�x���&ow�����ק�e'@�2N���jJ�+�3ƴ��ݘ//ݏ�SO�xz��e�^֤=�8S�^�Ly401�}!H�>�.�Z5(�o`~�eKMT�~�gY�o�����Q*�T��y�r\��:{��_�qz:�;���/ep$ܻ��\�(�7ri ��$��V��$Z(�3	�9�:�l��O�/�-��N4���Ó�t�J��k�Qͤ�s�e�f�d].;un83���������{ϝ���w�Y���Qn<s���<�q�����m���;�ǀ�.��N-�&m�/�I�;)C��z^��-?3Lʓ��;qȶ����OYG��~Tr��_��!�-��P/��}�uI`Z���j�R�5�_��b�1����;����˷��M�^J�;��Fyy�O�yF;Ǐ@}�����=M Kb�N�[�����F�MY�E9q��l�f{=*R{�݂^��\�|2�s	��:s��.+��zY[cD��=7���f/l�ٻ^M����4:�Ƨ�cя���=P�~����Q��ś�0wV���#�5î���3az��.Y[��nL�G��~�{�?��u�;D[sD���)訝�;�5�G�vküX}a9O�1&l���%^ݠ�#������	z$D��4�w2O/ʠn��]3҇��#@~a���4}�Q�T�"���.��������{���A��x��c�G���r`���0�ꑁx�.���>��(kT+�Y�/!�#�/�#������۫n���ʲwM=e��|����h��	�$r��͜O^Ƕu�$X��J��߃.���ut*���{Tva�ҟ��I�<wVv�V������gh^�n]-U0��v�D���d���%��O�0�5�N��RP�޳�d�:�$daނ]9ss�ԫ����:1ӵ�HL��͓k^ޘF��8T���x��3�\��]#+3�F��,Dl� �Bɂ<�+߽��x =�G�� �X����*�OL�{_��r¶)��HH�۞&Pb��P����a@�f=z���n�o�-�$t\�of֥�ށh@�a� @<}�|���� ��A.&�'�$f�G)�Gc�f�e`���rfvZ�m��\��C���H����.��,�����_�2OnbS�)��xZv���y�Jiھ�,YF�Hɑ~��?!E��{�p?AOH�nNhOu*Iɖ4p�3�q�P�r�G)k��"��&�b^���y�lY�?��M�U;�W�p���n@�SJO/t�N/ܡ�P�K߭)���Y�P9�iG�=��蓲>-(���[c�:�O��ݽ�KZuМ�nXey��d�y#�e��%�5�8��|kgaHd����j��]���y-�}��t!���2$�P�M��Սv;��:9=�}��`tc�/y�븨N"g�}l6��_\�>�	�|C����!�]|�%��}�h_���/��'�ӆgZ�4�vѨ�-k{G^�܁k,?�C�V�^A�幨C���О��Y?_��P��l���O7����{�-~e_z�	[�b���|�6G�I�W�g}Q���9�X�Vm�y�mX���si�r���y���]��ߞ�^�8��F�/��J���PZxs!�<�j������S�g�����ƮY�i���%�6�ۛ��S���?v鮸��=�x�������=�G��=�*�<���@��j��������T^��)}^����jڴ0mN������?LS���R���=�ĸ�b�%	�.I����w���h��q�"&w��\c�۹��]�Z�1�3/�EwI�j*O�c0{��O��Zz/6���i�$(�*t���s�����vv��s�{��zr�}F8fAX�oB�#!�ٲ޷U�-�<΅����3n�*;ܱ��Xc��=��
���Sum��{m���o�F��PȮ�s���a����W.�T?P��9�aϐ�>S�g�}�� {8��t���K�1CIY��|�=��P<��,)�;'��Ӓ��τAoB�"��v�2�66���Xf�`�ǈm0����N.j�A�$������ʤ�e�N0�ȶ�Z]�\�����u'����`//�Q�����po���O�~��	�����&��_C4S�xX�d�����4�Hn�Yw�y�����k�cc��n�iܩ��	�d@t9�n�ZF��v`ug�{
~��Sү|��V��n���$�|V��zz��b��-u���	ڂv���-�{\���w5mr4p���*�JTI`��0֬E$�=�#A�m�D����Ą[8�b��$y��K���3h,����ʨ˹��3N���5��񈪏x�/��gJ9��6J�SFxPaTO;�pPB�����6IeH�aʆ�X�����Q۬�r��:�]�*��TWW)�*����2P��Y�uh;�3sܧ���h�L���h���qcbJ]�m�̰dڀA�Ӭ�,�k��4�Zΰ�H�xlɢe���\�SΗ�L�7�_]^J��V^���cHa;�8f9��傍�G���N��v�Y�4Ϊ��� tB�v�6�R�Vi�N��a�,�;��F�\���˺�`�L��� ���ˇ�R����ogQ��k���"���v��ֱ�o3Ƒ�l��v��oic;���-X"�C�CEWA��r��fW��0�=I��6���6���Ϻ4j*5� �EѣC�w�#��s����LuP�E�v�����'^���EZ���(+�	�Ln���b�}�u���YNf�<�꫚��ܯ�,�o8��p^���������1Kv3I����h�U����ڸ$��AS��/;6�ؔ/��P�5�$4�/"{����wY�kg]�B��ҙ�a-g�u>��$=t2�4�B�4�(u�ovW`U+Is����u\QL*�1*�p�2��-͋�(R۝^�,�K���>��
`��K6��(���[�|�R?w{�?aEP��p�r�*�R�ob�<f,�T�X����ٻ��"BmطǃK�m�ᎎ0N�6b��/Z-���U2�&R�&Ik3�S�ʪ��zg�z�&7Wk�N����O��u����F��R�%f��[t��+`��LRr�9��4[�6���}��.-�m^����'��x���'��|�J]�ohjX[ap��UR!��VƝ�&�d=��ᒍЍ�WP�Z���.���׮���Ϝt	���s���b;�J���+������<V�����h��v���j�P�W{�p,D��s]tp1\�9�y�d���YQ=X^n�9�"9��l�k�0�f5��a��;�X�o�[zG��w+v�k�/1,K�1��)��|W���y\B��8v��&��b�dB�X|�6\�4�J�j%)=|����C�rkGXZ�t絋��i��c������`�6������\J([��fAN3���ۺ���s|i�NS(��k�J�芇�d�m���w���.��iŁJ��DP�73N�}9wlV$-eֆ�9poU����X^����6�����[����i�mVn��z9I] ���E��\�������4ADr�QAA���*�F*"��8�J�A�����?�ǯׯ�ׯ\������>���_���`�j��������RATU5C�梫���=�z��z�랽z��___���񢢖��"�*��f#UKDDRW������
�h�
�� ��(Ӣ�jj")�I�gZbh"���F�cb�h(o�1TUj�4�s&h �X������$��i��*j&*Z|6hhi)����C���DEMhu���&yÉ���CLQ%D6�J)(�*d��f"(�������*��$�l��SM<�� )#�R��v��`����F�M{�@�j�f"#M�3)U�T&�Ɣ�
gcDSh�|A�k�̮�/e��˹V��n���=}̧ys�I�E����i����&��A�!��a4'3�SY,t�� 쐓��@�/&�!V�Z�"����iV�N߁/a�b����t2'=��i���7P���:��	�[�<���M֠��
���_����(Sˡ-�@���=�yN�uGd���0ʢΞe]q���EJ��u\��0C_X��XA�Y��Hh|�=B1����W�����O�W�ڝ�U���ܛ�P�G'�~��q?]�5�V�A���W�}ʠ[�D����z�ﭳ�8w&}���}�3D0np�,��h+	�k\��Mi�Yz/a���>x��h��7|{�c1�PTvj�F�Иf'�+۰ͳ��\¼Lw��f8��d	tE���l����n��8�׋q����!���A��P6eon�1M��3�z�X/���q0��f�&��T�,����]�m3�k�h�'��3����B*�F��<��/���r&vީ&I�GVj��;��c�>2b��k�<��8z���.#��8��@r��d���ZzWv�A�1�C^�H�	��6-�z�*��:)�H��)풞����.凾ԏs0�C5a{q\��en��_��Y��ş��'����.�f��EFM��;;�z�M11��)�s�nCB�����caO+c���(�[%���g��Z�s��u:;���*l�n��j�;ʜ���� 
�������z=�x+/&�,�\��Z� ��ʽhФ���{cv���}O�ǆ�cJq-{ۍ�Yx>k����Z������+3�O�%5 LJu`%%�j�$�]�6s��<�{w/�'�iW�ݻz[�70d/��S�s^��E�;�=�2��c�=�����J�
~��Rqe �~�Ο<������(�.��\�W�	�p�����W��v��]g��������Ά�����'9m(S���H�/�V_�̛�X|B��>=3 �����`Wi���8�(��O^�(�W;[�|f��oBc@YE��;ۻߥ�'����������Ҹ.(���ڟ�����l5Jx|�W+H�)r4e�,�e5��;�{�c���Ag�H�G?4ڹL��b�z�ok;��v����]s"X^e&���O�.|J��ߕ��U#��-�l�����35�9*�n�*�ຝv�M0��o e��s�yH��x��~&}:�LsO�\�O=v��ˎ�R�]��2"�=D�t؞�.��w$3d�J/��g�6�����`e'U�Tδ\S\�Clބ.��궘���De��s���t%(�m�F��H�����z�T!�E/�ҠYzz�k�2J�.Ȣ �&e^MҺ�䨴l��ԭQF�>9e�ݬXjk�Ϟ�%�s�{c��ʾܭ���t���	K�9˜�-�58�����8���=� @f��8����fm������Y��b����p��焾2U�A�Gmeн�=�W7~�W�u�-�������C�nӴ��-�#b*�Ȗv�C!o�p�z��[�ݟE[�/X���d+���חHB�<ë�]9Aw�I�sͼ4�Y�X�f����@{�Nd�;�R%�=Y�53p_o�j��\b�Wo���]5L��z�2]`H{"�����י���[9�gYD���ov��f��w/���M�zF�%6?��A�bxO�$g{��o@[�zW�W��'�^%fT�����Ӣ%��5�d��[�\��?$k�̯ҕ
��-�'��vw,���Y/y�f�r���F���a���q�0�d�O�I�nt�?1)ЉW�ر��]�-9���!��Z���u�C�t��̓�o������9�����I���΋�o�o���3���Ւ��a�E$���<��|�x�Ű���!�l �.�Nz
�W�Ƶ�������'�O՚�L2�Le����R)�1��zi���'�Ql|� ����m1RS�췩:����s4������vo*'λ\�gQ��L���uin��(3�M�*��}@��U��@�bٞ`i�A4_QH��$��V[�;j.)�](�y�"atf���w9���±>ƌ���hp�el��G)�k�U��G������z=�����ݜ��j�|!ᖼs�vΡ]�����\��t�������pT��j\�oo�UCP��152'\׺�Sut��v;�'t�z�s�S3$βӍ&�z�c���D� �,/�x�����}�群�M�B՘�ø���Z�� �z�����?^UD��ѧ�Yaz{��x�/�p�mgh�pZ�E�d��a�a6���zU���3{;�0\����-��������cC������W���^�=ؼ�)���g����Q�0O�l֯3 �Ir]��/��=s��э�o"]�Èh.9��$i��T-S�j�$
����0�,�ٲx�3!PT;��Pm�e�G��Zs�1]퉻"<��y~�/��K;���c����?0k{b�&��2�}]�/��-E\����m��ot=!m-u�SY�1܆���ad��b�����aD=����=���/B�	e1"��\�5��_���}�}�'��g@���`�8~b�?!|��Y��;?k���?jO
�՜����MN�K?ۣ��$����y�����{-J3;�Q��e�B���r�=��J酬��^�"��.�a}����]]F��4	��6q:��3�X"�so.�L���hK�w	ft��d����d��C{����>����7��X�71s�#��^�<�� ���<=�K��J9K_�xЮ�%��إp�6�W�_!����t=��Mc��9,5[���sw5g"���'�D�V4R����nyن��BΜ���)���Bz��6�~�p��O۳w���6��J�B{��n�r�Bd��E'I)���^�o3nV���f�Z嵷���2���` ^|-�1��ۘ����2.��i�H�=5�J�)�}t��09Ҷ�^uu�wA���Y�8I�Cw<1n�fD�d���y���Oa(,`�M"⚐7�+/6�1&���e�#��}][�!����*����#4��.�TXt[񈄃:�f��/ig^x,`:׎Ra>׶֞zp��3��R���y?@��wE�L����q��ub�=���,��{�ٚ~�a�t��?u�5�����x��k���Y'��j����ݝܙ�+�k%�P6����w=~&٥��e���e���h�b����u]s��g��X���� &��s!�$n*L(����&Y�}�}�=�J����]��(�tp&��>�3眷t�N6����'F䬦���hml]��f�.��=)'�v�KQ�i�Wh�ґ��e���n^��&�\rDc�4�#��:��oc���N�l$f<q_Nr.��8t���V��b���$ڜ7˭ڎ�I�������{�G� �G����g{��_Wv�w���b��Tj|���߷v�ٌ+u����<Nz��W���KdVp���2���Q3_s��1'����.}�6��`̃�@_A/�4>:yv婃mɇ;\��峴����/������Ϩ���ƀ� �
~���H��!ܯɐ�=�B����y�z�ƣU�]{J��^ː܅����R�����	���U�L�[P����q��=��I%O��ܱ��*������&BeV�
Or�Ty����[�z�E=�����li�����֛X�:��֔"��#�����_�j;�������RRX&t�����z׶t�|�7eW�1;��]z�S�����y���.`��l-�{ʽ6fu:��%�{]��e~J�0��7TJ��&zR=���9�j��s`L'����������rT<�z):a`#R��)Z���ށ���n�����6ػ6�Nm�hwb<���J�6�̐Շ�Ƈ�k����ъ�ӥ'wygm���n�c;U^���҂ƀ�)߀`('���|�=e���a)��z��!�>�#��iӕh�S���iq%�����!:��g����$.Nq���qq��I-��KL��u�幃2귃'�x�� �0o���'+�1�Nb(�ڐ�W�!�Dj����WC�r�-������Y�
���x^����Ҡ[�Jg矼���b,sr��ɹ@����=�G��������:o����j�^�<D@q��2��a-���j4e��#[���w.c`�$��a1�z{���?��Xx[C���ܙ���y���@�
n���[���+�'%�?�܊��`��6b�����N	��ۇ����C�r���oc-M���W���	�I�N�_�L�P&��c���ey
y[u��o���Qb�A��H'd/�U�SZs��d���#rQ~,�����3��SN밋������� �q���a���*�q����#��EM*����q���O0v=m��v�.��Y�i�� i&^�x����ֽ �tP�T��.��I�^����[j�ț��ٝ����B),xt�r��$^ŧ�sͼ4�
�|a�����_g^`t��BL�U��'��0�xW^�jJ��>;�ǁSl$nC�l�|�=�-"��)�\q��x�������>����ϔG��Q/>���M�L� ��-D����
�1�kx����j�3i�i�x/��v@pQ�sb%�Ȉ�N@SJ� 3^���.(��I�#4Ț~����:�Kv�>Ț��"��Ս��{T�EY��"+����zuWB�nu├��E�e�&���s�ƹ�A�S�6��7]HWE&�����r����G�Y���g:��swL��q 
�NN��1Zr�_�>�|X��u�W�����/��x!G<x D"����?��{��^|��~��^Ol����(��?���nT&"�A;$�ǟ���;�s�~\��:��o�? �>o@�Ԓ����$ȶ����A��0?�@p?N�Eq_�L��?L�]E�f����0�j�����)7H�A*,9�����x������W��Bb���dM�ߝ9��y�uPn^0 ��ٹ�^��O�H�s�"�.�~�D/A��背n^���-�2��׉ƎR�����O�[��	1-�u¡G"�䜐�K�Q�����gw�wGP/"�#��vu����0S�Ls�9n52']t���=X�c�Rq^Y����Ϝ���c�,;uawn��kaPE*�wf�����8>��;E�K�d��Ė@�k-ti�,�⃅��-�i�ý����|�����Dg������G~X;�T2}�ܡ��t�C��S��D�uY��ؖ	 �3;�~�����k�=�?3���ȈV�͔�-��qɹݜ��]�;ma���n*��	�b�L�@��(�{g3��y�B}[!cWS�w���l�g�Z�U�&�jCv~t��\���5Q������&���#�̬̏�df��*r��wŊ���9��y�B?j�z_l�B��"��đ��wmD�uBq�ff�n{�]��d�մ��0Q�%���{oh��lYYē^��0��իV��������GVߢ`ߔX����y��a n�}+���4���j,Z����89�S�´��j�o����e����	�[�a|��zg.m���HqW�C��Pj	F�`�Mu&��_Y�9c1S.��cŒ���+�){�#�]C���[N�I���Tݯg�Z����;/^I���!0Pdy.�g�`��*���J���?!O��[K�
���+�L��}�OVv�olx�P�hl.��P�_�J��d�WT\<��<!�
�����2�pe��L�od��oq�%�y��a2O~u��$h'P�n:5[5�K�,��X2����~���٬��Z���6K�pe�Μ�P�I�	�	{�Z{I*�\�`w�xa3RB��˚��8�E�j�C�>6L��A.a�[�l�3�1����L��m��F"�7���"0���W����{�筝�5����y��Ǟ��n�:��0��y���Ox�3<ny�a^S���Ï�s��D��Cq,V��_���m�/%�xu�q_��m�}1L�S��e:���C�;�%7��%�ϳILsóS��<��ħ�;S�ۻ)�'9�[�J;�c��QТ]ق��f��+���Vx��γc:��=X�k��ڒ�0�޴s�t�3Mu������b�f��ę�cbo����TjիT3{���x0`+
]q�V�*h�|9t��V>�� �gL����:z�B��	��#ޙ�!���]J(�Ǟ�\ݨok�c��{�s�J	^�g��\�q���#G�WᯏT�鵪�}���n�E��p�t!ם�R�����ҨO�Z丌�Mi��\�s�!���e��k:��Ŷ1C�s)~��U[�0����_�x��*>{�0�y������nm��{f�u�v�s{�������r���a���dov��fE�������\�=��-:�_nڙ5���{�b-�<�1���@�}fۤ�%�ޛq�fA/�5i�V=Yz�$v\���-�d	��3
$ךE���]Q��U��|�!�B3*�X"pi��
#�!榨��3�k/ot����c6���u�>���똨s^ئ}�1�`Qm4ϋ��_�E6ZݽըM�1c�	ʖ���,����g�Z4)<.�����zޭᩗ��m�0l��d�������*�y8�و�B��6��S�Z��Oi� �	�E�B�6s�~Ȱ����:\;���v���g+��P���7��ֺ��i�uG�,	v���nt1Q:Q�Fl�w�0��v�g{�@�]>�2�^���Q>��Ity�
�T�����U����ʓEX�l�M^t���gD/�p�#���w���r	t]cN=�co���φ��T�mK�茐8�鹯�l 6������4�v����Z�"IGK�w�Z�u���L�X���E�B�kp�����uH�`ɶ�:Ukt��<��E�=s�l�9���]�{כ���ʿ.;6�z����Rd]�Sp]ĵe����e�-6+�t�djO^�Z��A�e�k=:���I,�!n�|�)�޽�Ѻ��]w8Q�N�Ɐ�pKsQ�{@<�rA-w+v��fХ­���YmN�[lLl���d�R��ڲD< �+3s\�$�٩����q���l�\�-���8�6�m\�4�L�cn�U�ܦ(��7�GBf��XE`@�ɭ�Y%���|�p+������0�6��{*���y�p��3׎����>�++1S�V��X1�o�/��El�kf�c�|�޽�(:Ub%l�;:�@,����3��z�t虹t�?�uoQ�S{6�ִ�'9�˓�yD'�]4��#��b�.��W�쑻�؎%y����@+�	��7aL�ݮ�u;��(>�q��:���ʤ�V��=�=�wW��EjFL���w[;�A3(�޳�ق�kR���X�f�Y�[�UU�՛r\�c��>m?�V4=��V*�*����Zj�g8)��֠�dALf�R��*�4xA���c�=��븰��6"ڃd-FF�\¤�Ut�;S�h:/��c'u�v��i.&��joȳU[�Պ�ۉ�NfsR�0�>���adB����#�r��B���N�8K��n�.l�o�h-/��
XWyt�e�O�KƟGt�W�EعEo�	�h�yN`��)Mlw<�6m���~�(vtC��FuA��PNK�ɛ]�AZ�oV~A-׻�
y���H�^=ǳi�k�ɋ��N�Ӭ�ʲ��������'zF��E+�i���y��>ݼ�"��ӽ܋�˺�ːZ�2���2�Z��*[91T^��r|�s���xA�<���J����zU��=���_5	��]>0��9Y�e	X�R��Y8j�TS�Q��X-Q��H����KٛU��Bcb7�ji�Z�-�&л���Ǥ̩�Wc�١��j����9��/	k0&�T_AvӼ5qM���]���}W؋���t���^�Hۀ�=X����I�xn��L��ܭu2e)]ҥÐ��e����t�Es����F���R4�>ʁV�lw�(F��)=��y��v��2u;��Wn�L��+�V�Z������g(Z�6�[C�d�q:��X��q�n����1�ݮ&u4�|��x�"D���`>FB-����T�`�E�`,��4d$�l(�! ��jAI
�^��L��Fi�� �f9BDQlDЀ�f���H �Ui�MT145Z4�IQ0E-%%-^���j˳�,���,�e�[����n��������?��b(�#�q��tP����N
NlMď_�|}ǯ^�}z��׏^���_������򤠘`���&�J�
"*����(����N� �h���6�$�QE1&0�hb�*�����mD��4UAQ1T�ST��#���"j**h��ckEEUD�D�D��PD�D�If�\�RC�L��lh(��*?WbV$"�
*����4�ELQ%EDM%4EI@V��cEQADA��QT�̘��KcDT��D�����ETPUA3UEQ�AT���K 4D-%&�QA�:$A\�9Ztrv2Q�٘��*��F�1MQI����^y�r��UՁ���I�!�K[�w;xحs&̓���h���9�-��z��oN㭛�z�g+��'n����M0��r4ڄb�nBS&2bĎ�ǜ�d�I��<x<x��ST� � <0�%�'8mGC���y�^���[Bs�T�)��g��2��c�:��+����WZs��6�����)�0d��h@�!-/P��WU���(����.���b�`~w��:���t������:hqsn[]�k�w�A;0��!6И	�}}"O[ճ���0��WB����a�)J�����ZPX֩�/��#^0��}��~��|��l4�Բ�mi�y˭`Z�-�w�UzY�R����9����r�A��g����lu�����n�:9y8}N�LK[T)��OV0��es�PK�\2��ƢX�`�
�]���{P�f�;_r�ް��"~\m29j�_K?/X�u��v%>�z	Aly�����M��ٜs7��s�?Ty��`���(BO C�bz�d�;��w%���k��wwй��y�8�s_	f�KW�܈�b�lC�xw����x`t\H�Se�K�%[�kvB۞�YK�uu���Q�נ��dq4� ��p�iy��&��t-�G��ɣ���?i^���W{�Q��͊�ef��&����\���Hk")1�de��ι��l��؈��_k"�[��ۉp?��%-{���:(-s �Vf�k��:K�9N���덀�"�ې�:	���yn���堩Z��0�2��W�>Ͼ��<j$J@�s������}���vN�6\�^��}B+��XVXB�IwC]���KL�P���3���W������︰��'�2S��#�����R�j�o ���`����C6q=c�:��f�,+r��+��#׸8֌���.=)�;7��D���2�&�j%:F-��o��K!2�g;V�̥6��O�[�!�.���� .y��
b�kS�\��=����5+��=��{Qcg�P
;�=����x��\]L&
odp�vJ穓�q�d�nF,��Zzu����%G��z��3�>�S�#��gG�� �Ƒ
��
�7���R��#�o2_����	��vq��XR��q#ܫ�'�9���))��^�#ϯl)#Ҧ�����9w�y\����0�l�/#�}0ۏ�e�����̤sH�F���Ot�� �����ݸ}ke�Xە��E�/.1���/��'�	m�n]����	��O��c8����wV	��Ki?n����]�ga���ᾐh0u�>�,z�̇��}}t-��z���pBΞOQ=���ŵ��=Y��V���կ���y�f�r�#D$|N6�ņ'�(,�(�#O�Y�֭h��Pǔ�y��nۤh���m3��o���%R��#�76h�W��3��&c�v�G��#sm4�p�On�j��P�o%��G;V��`f�l�er���|x�g��X�������������H�,"�٬c�g��>����!�:/^����phZ���m�����]D��Fi�E��ǧ�1�>�^�h4vk ����?~X ����U�ۑ��������)�P����ӿ�i�x� �3�[i���G�ĳ�~�<6��r-�n7��8cni�@{^���۴^{p������	�mi&z t���xl�w˞�(kt�5�_h�-�0j��q��F��sg��/�E{�O;QS��r0퀾���ܧ��Y�-��߯���
��b���P�P������ϲ��mA!��Ŋ��`�6�m�btX;z[��fSCf������2sm�"�\pqd�? �?��]�o�um���R}nE��`���{ڔ�x��R-״���L� �v8�\�C���3�	�_�D�g砞�6�ym�(������n�sz�C�Gk:�I���B��O��k�d�^�v��+)q��Q�PPdb65�䲱�#���T���mj�̋�xN�#A:��V�6q��ȶ_���}o�/މ%���|�Q��+�2��xa�V������t��m˒�Ƶ�Տ��Ka.��%N{u�iѹSj��5�tq��x�4N{8/�/��tg���rZ�i6����43$�ܻQ;s���WK���>��pr���G����������A�30`��3 �xu9��M�}AĈt��[�H}�B���y:��2��)=��O�|�`pCG_\�-��]�i��F4â�u1�b���4�����v�'Ģ���n��-vw��wƦ�k��;�=݇��t��$���C�P5��=K��"z�e&C�O<ϝ�l�C�`Av<x^�ܮ�4p�B�t7�S7�}H��i�ƱO �2��h�㼨K��M14Tn��Zz������ۊӳ�:y�XWZ����4�������maA��ܖ�U�.a��#�wP���Z^; OJ�I�p)��G0�׾�kÕ��W�K�Bp~'�~Y'�b"��,�2�W�1S(����r�sW�jT��{&�hsH=��,{�]ah4ܷ(��v������<B�0��>�C6H�TXQ1%��{�f&F�F�Ml��J3(k�/l�g�ť_����[S�d(���wh�����vXs�}�S��a�!T�g_F�ݗi:"�F�S�p�`�e�0"������f,�>�~d^�FT���@�}��dk��yF������e��SS�`�U��{ܥ�W^�h����T$��5���}D�W����oL�ѻM#lN���Δ���`�۝���O)�eK�"��R�x(b�":�[1+������[�ӕ`�e�p��w�����S�׏��<"�)e��x����iw0jffgv��̳[��%r�F��.6�5t�Á#^Y��s:N&.��3f썢}�RQ�|�ӫ�9�"����-S����%'=��sƆĳǐ��c]G(�(�WW�Y��b�P�1���tNT��"^��	�Z4)=�G(P�1�3����d��G� �7�sy�Y2�ࣛ�C[����4m�֠�D��bS�JN��hJ�R
��(;=�Y[xn�-M9��흢^��M\���pK��^����.s�a�.Z'�!�{�E���o+No -�wu�\��`�����^�*��I���z-/�k����Z�T��uJe~m�c@�
�'�ٞ��lwow�A;7y���^�	�����c��c��<�F!��J�=/@����9bF�N�ԜKGl�#�67A�t��I�Ք��������3�Н���#S�9"����Y�i*�K sI�EÁ;Pr�@;��P$���0�c�<����ĵ��ƽ�8�s�¥ς��N��x���:���s����f�r��Q٠��-��]IL�؟]>K��R��i��ő4�.�E���8��ۗ�KK�����6�sD�X~�I�w�es���M�	�*�E��ѳ��{Ȣ�JI|�w��Et��AejQ�^�.��i��9���˿����|x��x�9IRE�ϿϽ��U�r�{$0g�;ȇmt`��_K?_O����$%[���ղƢ!�$��j̣4󧷔6]C2��1���>�� ֜����M�	ɹ(�>�^y�ūJ�3�8��C���ohvx��g����D<��'��#�%iz3)�*6�o2�s�������I/`Ѐx�v��-���ב,��\s7S��p�ض��9����u/\����fZ��K�L����R]���Z}�yǆ�yg2�ts�u��GUV�����[$qi��= '�zkҕ3P�1�T���Pz�^�wo�ە#�!�{����e~��q��V��RO���,o��y�_т�^���HJl�eMB�R��ޝ����G����.N�{��j���T-����a�.b$.�E��-W5 �'
pԙ�3C�{��75G"Վ���7)P���ơ�l�����O��t*9��b�)b�|�e���W����ۧPY'�p�M'X��lIJjgہò.P@0-�?��Ԗ��k�}����ٷ���J�e,��6�PY;� /��Gi�(��T�1��>�2��l��B�,�r��(��@��ؚ3�v)I�܁-�͆�MSS�c�Ρ���bq�Z�N��gU���"؛����_���|>C{��ZO\u�Zd7|ct��&<;��O�a1W���*��Ln=a�����0�b��Ȳ׍�U��h�|����^7[�罵0ӹ~�e���`O�n�R6��	��r0���K�Q����7��>&���9�=�]q!�3z��Kmn*]�����_�Q���1�a�5*^��9i}Ŗ�!��r���C�{�	��k�"y�R)�GM�`-����=��Ӛ�7ӳ���ӭ�a���7>�U#+`�"3�����!��a+�%����}l��hZ5JM��v�rmn��ΒÐ��nװ��Q�֞}����ۮ���?M�0�Ⱦ�|K�Y�ـ���E�+��L���[%86��
$@;��nZ�^1���/a�s;<�Y�71��9�0�S=}��OSݴ������ǐ;qP�k�E��Ť�q ��,�z�S06sy��\�#g����:(*ǎW�k������m��̜�#��]�7��=fr�z����/��f+i.���2����:�l#�ql�ߦ�zg.m�PHq|�1cU,����*�w��޷ڻSyvd�M��3��N�7�U���o���Jv�ĞC&qGg�˨������[��-��D�n����{�9���0�TқT���|�3}@�Cξ�m]Yj�.P �оg��p�;��@R��ð�'��?����(�]K)V����7�+��G�Z � ���#!tQ��N��3,~V�;�?d�i�p��P�{N!���c9~�똨sC`3?���t�o�n�?~G3�����-����a�70�-b�+zu2Ǵa2�Z4)_�QaMG�q�^��S�< ��d���u2���V�n�C}s��d#�KkW�`�.��:�@B��]����[B�Q��n���M���p͛��7�62�H8��!�	�h�:D�J��	�M�mi�$r�(bx�^3]�s�S�oNnڬt�m��Q�0�?T�#�E����v]CH�<�Q` ["���d�.Y����yd/��*]5��^ý4�c�peϞ�M�,Ȟ��dS*���"����s�[�.7+�',qv	-�6 x�(��_����e�_m�N�s�������м52u�߸�,s����i���T5�p��ys�Ѷe��Aۃ7��4�c����Afг`��OJ簔��_�h=s��$u&�W�������y.�F,��{�yojy�T7Z�g�ݘ}�]�>�Z�{�4v��$j*#��[�#S�:H����N�,�z����S4i�#���a)%A*��5l�k��J�\fu9y���,�R��ي��Χ���a�e���.3.��;���j*��L�v>�a�B	M��)�4ïO}��� |�����<�83�W;�s�o�9��O�Yy߳vS���@�~�װMzEm�C���ҫS�\�C8i�����+7�@S�l�cXO��AK-u�O��Ә�]��U�1%�f:�IݗmS��c4�Z��3{��M�����yw�`F����yOl+�Ql���7y�v1�=�;������8���q���N�-mÞ)�8f�^�t!\>:O��oM����M7�����iL��X~U}��B��y���㦮��~hg�-�G0A��@�;�Q�]y���i��U:�]	�l�t-��h-}O��i�*�Rp�����h��N��g2��7^��z����a	^v#`��F���ܨNT����,!2�hФ�(�
�1�M�U	�z��b&{z���׆\���8�L!��"B��j5�>�%��XJK�a��N��tۗf���klkBz�K�x�:la(JC���"?~99;��!'�u9!��YSO%G<�~E�q�n�������B.fָp >�M�=O���#�r�`�)��=ۿ�f�]>���7�#�����h��F+q߻&��Ï
y���`U�q���of�]���u���^����>Ba��	�g���9f�\c����[5��v���}bف�ZT�wJ8���Օ�����^^^���b�Fr���a�����U(���KL��`�Ahw��Ђ�a�m��^j4����i܎ȓ^YJv�4�^��$���R���8��p�l#�wP�Y����i��hE���D a�hL��4.�*��,�e4�硉���-N�k�#�\J������U�ݹ�}�C�h�as�
=��	�lT6�S.��aܡk�%����\�s�/e�r�E��ѷw$R��!o0A���?��_�Du|Q'qms�o.�B��^5>���UW*S��QO��Wg}������69P(���Q��?�{!�E4kaz�d�>�͗dCA��a�#����q3����KJB�Ͼ�o��cSuv�w|A��E�/v��I��9�U�Uv�;u}��t�mc�z�&(�D<M;�O�l�P����k(���ô�\q�3��j�v�:�^��./v��fDgt��WA
�$
���Pio��77�+�_�?�/��c: ���`��^��1�睾��{*����x��	�%�ǂ�w쨺�p��M��b�˛R@�Ϣ�ꬂ4fJS}��3�hV�=հ��R$ɓ��m��L�6���;�3���UL�)�+���i9D�b�zŽ�ۃ~���l��BU�Uv,�J�������-�!�����A���}w\.7��c��9���5��!Yj��<Z��C]��*�ޕ�¸���&(��0��̙MG�ku,m�b��ȵ�K�8T�{K�/�k}��`o���eK�)��"�Z���#�,�gBbl��]��S�8yi�(ډ�</���L햐�#����献qq�6�z��k���r�k)�����fќ-f����i�f9\.��f�� �[O�Y���b�r�3O�o� �4RY����UWZ�˄I���i:���y�^Ky��U��T�S���ު�3�<�*c{zL.%��d�����7 �8+W�}���ܱP @�ǹ��q�����jwQ�b����E�Ơm��p�N�g��^ja� �]kV�����hb�{��M�ٓ}�d|[�`�Xք\C��V�I��fՖ��Ӻ���y'-�魝/52�|.�.��W!�ܩH��M�v��8�/!:��0Lc_8F�M��wMwm��V��/O�^4�b�».��"�]���#v�ta��WW[o`+%��y���٘��t�Z���J�0�;��
�Nu�*W=�)I�b����zũ/7{s@o��Q Mبȼ����0c;��r��˴4A*�{2���8���]m~y''������z��p�o6�KxP���Zm��i�p]l���d�씶��fU	��)���RSb�
���g�6pi�]̖�ݫ�{���j��a�s��w�f>��o���9�s}-�G�C5�΍h�ՙ�tS�3�ݜcW��[��FV<�K���+zi[��Ʉʯ����{�J�ؽQ̭����ƕLye��M��ުB��3����B�f�Q�uX���`G����g k���Hv���!k\ӄ���![6�����Ŧ��R��a1�
8v��|�L�f>]�y���X�,־Į�N#z��ebI��%.�a�T{'���ժ����x6%�J��sH'3��#x�D<�-S�Ƿ�Up�dB+h�����ҍ��h-q���W/ٯW_]ź�2Gjt��ӱ������9��e�H힟<�ӑ��5��ބ�rs�X��]�	��$TJ��穫`+2�:R�Sgm�G��	�=�%��=/x��9�C��Ǯ�M�>��9W7�r�b!�p��];{���)�.u"�St8ђ�NӢ��T���FHd��n0��].����i�蠐���%�`���3wF����ǉ�Bww>�av���;X�sht=�?U���b:�)��RӶ��������'~8jճ�ggL�e�,��VYnݻ��߯��|�ݢ
b
��R|l�QT7-AAG�"�i�hi/�׏ǯ�^�z���ׯ�}}}~���_��Ġ�
���)"X�(iJ�>gM��UO&���5J�)��h��I�������()����c��b�`��i��:`*<ڢT�(�(�
�4�C4%UE��)�����֊��)/Ɗ"h����9
)��6)����<�xf�����=����*a����4�Cm�Z���r���إ*+�h�d���s��-ͼ��̴k��J*�� =h��#��A�TMʹ�����pk�G�C��[��a����������"�q�P�Ύvq�bb}+��@hV�ݒ��-֒�|_"Q�ػvKc��'&1�N�n3�������� =I&����3�d�+���(�G�.�@離���n������M�����������T{syt��`y���[�{fkA@����=�d>�U���v����nz������+�%�#9�u�RT+�k{l휼�ۼ	�TIqU0�,����"l�����]Ο��qu�0��1)��)�u~IRkkrD���5�@.-�N);m��V\\ӧ���̽Pᡟ� 3�d:rA`g�L8��T��LU��E*	Qa�K�}|�|��.�f��i�ggӍI~��8����t!�_<��Cl���mL4��̋�����Kߗ�Z����grţ��C��ȟ���U0[�|לY
9��D<6kО�m�R'����){y�B례�RV��Wv�����(0��Oج�8b�����󗩑:�T�n���k�ї�,�<C����}���\o#n�l�Յs��FW��D� ��i~y@�����E� �LWT�[�q/8U_sv���D�a>�m<q�_�s���M0r��h4vg��nm|�V��c՜׸.ju��{�V�=�f�;���[±��\x������m�N��6��%���DU9fsO9�����Mt���fb�yJ�YUz�K�]���f�=��ۜ�v��9�������gm���ʝ�{�q~� ��� |Wf��ur-t�	v����C{`�҇��$#|��*�N?[��^ø���eC1�Ϲ5AYѶ�����h�<B�6&15���#�
ė%ًi0]���.Z��>'dY�Ջ��/�o��K�ִ 2��z]"]�`qE�k0Kȇv����}�w&7���3�OngJlf#��ugw�٣V��O��~>b@>oql��q鑗6�j	��Mnj�V���ӣ"�R�nt1&h��e��T����,��Pߍ�d.��{���˒�j�z�.�3Uygz�����O�b��(�^č�y��Gc�'�r�@lg��Iq#Kl�ļL��i��;�ڪ�L���]��2�\w:cW�$�TXSQ�h���=��=�Y��6c�;��n��M���0y�}p8m�ml}�Ľ�1)Հ��e�2�T�N.�8����Ȗ��/�kT��v�ƊCg[�!�9!���}��$wM&��|�bdU����[H4z��֖�η��c�T�L�3~���_�\�����!���CO�*y>m��j���#3+�_�,u$x��S�R��K��mEՇ7Qj[(�G�rd�r�����ܧil`�
�����̢2��d6� +�$�p�%Nˡo����yŵ޺TGMv�*�V.���I�蔟^��q�5�@;TZݲ8Sk���J;k�],��T7GZHKr)NB�R ��m�@�	�)������^^@7/�<���;��7: 5��y�ܦP}Z��T��-dٯ�Ok���T_���'V.�
n���ӛӕ��"�.�CR˔�҂ƽ�S��'�qr������M\�
��]r-��u�;gWS��V��[+_��E��<ʕN�����9�ñ�y�B��3e�������Gk;�,��� pX��f��bN��ҹ�r^��Ts	 �x��X/n�ej������ӓ=h�5}�0@�;�N��\��vm�����j�^-W�9��7�c�8�P��I�̬SP^��8���k�Ϲ_	kM���-�,&��Y��ʆd3d��E�/�sjQPa��#^
�nw�6��!�d.M��gO:����4,��S�m
t����h���u;�>�,�b��Ŭ��3��x�v:�Y��r3�e��b�'�(1�� C��F�-�P���[�EF6c�xj�<䫐�r5��L�}hg���[Ų�y�O�PqѯyO���{L#5o��vXƞ�!c�A�Z�	(���ӹ�==��������U��u�c����f��غžY/�Z��*�k�P��[	�d���t7vF8M���0�"Ց���"��2}*�0��F��]n�����\�>:�ㅑG��)Ԕ΄�(�Ԧ"b΁qm�cWFZ�jܠ�*>�[���n}��{��G�����������&���8���Z0(��̿��KD�K	��)�ɐ�U�B���Ps�b<����ݝY��Z�UZf
VQv�˼�A�!�m�֧�$��A,CK%	�;,�����.���#�Q		�>Y�8���C��c�v�
f+U�a�1���z_v���V��{^n�d^�E2����[C�MzY����	�ש~�7&Q�r�2�d�Wot�b�(�'L-�]ye�i����y�6�;� ��«^XU�2,��w9Ǹ,n^�	��8eq=�z]�@6��'�$j��͉��l���aK�N\E�����{����{Z�!㟨Lsi�&��%Q��,�e4�祐9�D]v'��{��i��R�[�4Bg�\�=��zb[Uh�)�t�[
�R���A/t뙪�U$Q�y��[�0���ڑ�Y�Wa��o�K�Q|Q&Z�_�:��d�$���y�z��W�q4��5O�^��1�k��� lg:��ƴ����`u�?s��$%#�K[꒤z�B���Z�gn�~��C5�GէN������!�ۻw1E�����*�Z�*�̝��i�ԋ�+�H�S}�n�[ϰκ��c�	�v���xʋw7��}�"�#�3�x�@\�zJ�ꪪ���o���?�<^ZL��LPf����_X�'�`�ó�O`����7���0:.���%KEF>@�J�fl��o+�@K�=�!��m���rH�dq4� ��N�T?c�<��N�e�lh��gq�l�>kd�Ƙ�Bd^��޸n��nd���,x���R]���wyҨ�4�r6����~�ʻ=��΀����:=ŗ71���zkԕ3W�ϥ6T������A/婫/���U�3�s�n�{�t�c�9�dS���jâ�n�mF0F-�ݤBkq
�E<WEu���2�9�gW�Fc׭���3[��D}C(&Fcc�  ����1�T��w5gq�A�8'�N��u&%���R~���t�Os�=�j(����I���9����Xj$h�X��۞���9�x���R)�$�5����ȸu]ޟN��l-o۴"����ӣ����fB�|a���8�wQ���LU�H�B�(��X;Y1��U���]���W��_�Z���|�������a������k��LZ~A@�a�vT���C���.W���h�PE]R=�Q!��$�o��%V�:�3y����M3� �c��ƻ&D(_�Y�
UӊRC��,v3�0�#VWW
W7QU����%�H!n5xJ��j���w��ulg=�nfLtvh�У������{�֑Q�ɷ;m��Ȗ��kH�0a.?j�9õ��
�;'ܦ�����m�54��خ�U���St������ӌ�M'��!���6ܠk�߫�	����m7j(�͇'Z�e�VvV�fj���[3�eک�{��gF�{^�
�Ʀ7ͤ�j�
��[� F�x���a�E��9�其�dWj�;ک��$V��a�Vػ��}�M~Kܶ/^�h��<�cC���YQ(����1�kB֦^���۟$nu턜���P$G��&���n{�Z�#f&y��wwe�)����'��~hq��̀���3��r�F��wXO����˧�-zb]^���(7Aт���wijNw6}2�}bo�Iv�݌�nbcj��������vE���4S�͖�38�`L�"�5��/�z�}[�L�K�݇�ڲ�ڸ�۳�׭�t�Y�̕A�	1l6���������z�`@��;���	r�zM2F��l�RNv���&����Ћ�at/�֠&T�r�n3�1P�u�h���e�[6*_��eϔ�c��4�N���6���O�ա_S�e�����ʴ�v-���nε�k��9Գ��7��XHi�h�b���yo����0����Osx�{[���#=a�J%J�隗']���Iv%n������u��:v��pRP5 y;���y��x�1�Gf�w�����ߛ�%���"���c�d�ehȕ�U�{'����q݂[������g�彎`R��s����nkgG8��^Ø��#!:�\V���cYuj'��ͼ��4��A]1��ᝣ���Ӈc����bGi� ��L�1��-�_���*�lC�Q��7�����v���x��U�Axy�P�i�����Z2-��,�o���%�h�8CP�W�=��S�<��#\CiG����6����O�p��;\�%�s������������F/`��Zٞyn.R{	AcZ�;	O�q�Ç6�X���I��*�l�nj�9�]	yO���:��Q`���Q��	���sӾ0`�m���u3�7�F��Dn頡�y��w��xn����qP�f$�'�s�PK�m~
��I�l�CU�1�R�6�n�Tv�^�u V�+�dY����W�όag�"�^\�݉L��'�{&��w����d�F��U��qX����<�<>AM���~��������׻U[���m���so1E�6�F�oĴ��n��Ì���o�w&�!��
돩���K	+c<E�z��R��V�-�_l��+:�Ϗsҥ;���օ-�yasJ���E�Q�鋭6��i�&�ͳ����P��c��U�[��>�?��?��7}�bo8����3n�2���ȋc^��^sb����{������(�1����;�������*��qC��q�CI�.����x�����0&Be��5�=��h��;;�6���S�s�Z�ۻ��%����{���q��t���C<�VD����M��n����`�����ֽˈR6�[O������b|-]A)8��ٳ��v����6�iT�1�ka��Dh���	f"�=>2Q�/����&BeBѡI�/0�a�ԃ�o^Ww�9;�~�?w �K��Ul�4���V<D���l)�h����D�i�LW�����0�Y3.��3L�8k��8�`Z��~��ǡ�l����8o[Ǔ��^��2O^Ή������ṃ�c�K�����^X�Ju��YZa�-�,T�S�N!�-~/H !�%���������h�]�D�:����2��q�2=0��˦��(���T���9f`���a�!��FN�}ٕ�k�ߴwď�Z�Eċ@-�`A �'���b��ZPX׷��\k��J�}}�R��n!2|��4��Z���t��W�&��O�tp������ƙy�l�Q[[�+9ʜ�*]]]U�o%�^�7c;�1^��]-���3�s}�+]o��cɠ�	�������4���]c!�up��Uˇ� ~~@// =��˼�$�+�d>h�`鹦�gg�P�^q���м*L���c�&E���f�LE�Lۓ�_r�iiw\`<#Xs��-~ن��*T�룦�`�R��m�da���jz���k'ye?S������lgդP@�~��+��h��Ɖ�S/�~�x�Ҫi�'`X����%����x�}�gӮK����f�OA��\6y�p���a��9�Z�#�����}̋����~�f\�=�@�e#�'����?C;�����������NUu�>tNdLa�����D׍({���!��m���r��;I}��6"����Qt��Z���>���4XQ�웋�S�6�z=�}B(wI`J�h�%�9�kՃ��ݱ�Q�JK�E&x������~BՀ������=�����'f�fc����U6GLN�ndWb�o,al���A�f�s�S:��[G�:.���Ql	����.��^��,=��1^�3���TJzH�0<��+�;x�^��P�k ��z焃�/�}{��4���~�i�]x#Kr�j���K�̒����f7ٹ*�i��K{.ޛ�4[�[�vGk���Z�id�+޼��!y�*V��ņ���x�T�l�v�,(Ȧ��V�� ke�lf��ڦLGF�uP���ĩ�K	��=팈��C����?���h���a=d�f.�pK�"�N1�e���PQ����s�:zkw�\f۪�Fnb����ΞY���ۊS�ȵ ��<���L��xN�'�	*M����O"}��[)�x=�mÐ��ئ���V�fwxm`��li����K�e5�nGC��k��k��*��"����xΈ�-�Cэ3W�٪w��c�?��l� ���Bn��������L�H��\��b��ys��0i{���djʨ�ռ����.�a#���[!F������	���mxn*t0���J��"������ �˒���~����eC�l!}�5���$]h5|Ϧ|���fVO^��5�cfڻ��	gO'�
��T��l[�63�Z����� �Y|q9�F��鸓jvo��n{�B_�N)A�,:��2װ	��W�4�r�^�A����7�}��bͪʮb-���``� ���v�C�:�%۟'qP�픜��A>�<���i+�%.��ۙw���u��C�^׆x���.��۝��M��`��#Nm
� D��L3s �l�&�j�����҆[<�V�r�/��f��Ex��Z�ӐB�h��pB�cU�����VM� �ۓr�e��.(�	T��\�.8�z�j����̢wj�=�`���&PT��/GP;կy����z1�j+�Aj%�t�w��3�rn숭:�ì�v�A�;��ĳM���V�e�Cp�,����ʔ8������.qt$AG��Ɛ,V�|�q���i��*�J��촲�,u�}-K��.o]����Q�[�4&$N�+�aT�`��).����3���ٷv2Qڝϴ�,����Q�'=7�s���̸�ޖ!���39�v+VMU�7�w�`�z_Kf�Z�1;O�� �'����I`Zmm1_-�w\�<}e6���Z9%W�Vn�}~Ռ�W��c�2��Zy�'Q'���@r�q��jgn����q<X�}�[�|��pn2��}�����[�dKL��tY3W#z_.a9�h����#H�б/wf�$Fbo���J�3#��jk�IPV�N��15�Kl�*����QuK,=h�1�*2�s��;+�W-�oQ�*^��ݑ-�8,�V�1��^]o���f<����c�RU�7�j��m�{X
���v�YOd/ym��sC��ī<��{Ӷ����;�q�c�
J7*�[�\YqL�����S�Uea0�(1�|v���t:���wv�����<XA����;�v��B@��L9z�>`�m2��1�U�ETȥ�ʔ��"��J����EV�K72E�x1S���1ը�������IbrU̾Ξo\0�>E���U��6��Ly#�m����b
����Frj�*ƹ�40	�!�g�-��7R𸁭�٘��}��V���m�����i1���ܚ�]:pXr�7�K"��1k�X����Ȩ��#��iڱ��՞Wɇ�G���Wn�V3�1�V����v�_Be��os�M�-]�ȇ�TV��I���V}&ȵXt��hc��Ue�,�O�,'ƃ�Žd���jƥU��IgaO}�͹���}�FY�x��{�o�I�n��%�۫f�'+ gF��X|�M�;�OWu���l�{L�VB��[au�ԗ��d�$�����FN�I��E����#�[`�X��*S�eL3u���,d�ޏ0܅���k����.��ꂐ��xF,�defVɝ�M+��WMg�=ke���w2��J�:1U޶�l�Z3��g��C4����7Ҩ5��A��h���]�\�Б�`gJ�y�}��E�FAIW-�u�,��7c�rX�*�PD;m�Ž���;s�#U����]m���9�yӆ0R��ov$+��2�l��z5�+�]���
Q�Q��Y��v�3�l-ӌn����&��:rA� »�=�9c94�p�Ԇ�	H���Zl4c�~H�"ZI�1�1D@6c!`��E�B�A�%($&[�$�XAH��G�l4�Z��哛b�DTQ�TД�\�6�씑4s�ѫv��ܲ�-�e�Yl�v�ۼ��~�>Aٱ��j��u�m�IЌTpƪ+TRo��CIVƟ�������z��ǯ^�z���������~��@P��t򊚣��.��Ēlֵ������-��j��4P風j�t�Ӊb�i&�v-��Z����)4��7�EG1��誨���<�h9�QZy�P�r=	Q-�i�V�Mi"����U�y/'N�֭���(u�A�I��6�@j�[`К���E�a��4me�w"�h�hOV4�yÐ�
+SRi�kHm�J��`ĕF��DPF��ъcU,ly��	ERS͟78h4��UgG$�EV�?9Mo�������o��\o�ݮ�nuk��ユ&��k�����l�=�g��eR:"[͗z3�7�	���F\R�7�DE4F�AF�d&������� ���������_�Sc�+^�$�S�������e} �"O��k���}�������{w&DX[E��L�7c�͜�x��vD���	2���W��g��­��TC���( b���S��퇭���_&j�����ΎN+�`�,UB�{� �Ξy��� ��:��������mn�5�l�_�<ǲ��<��&��$��Z��S+	�z8���s[�y��_m�\����V)
@����@K�<�S�s=�lc�peo~&*�hR�*�
c�ݼn٫���}�s���Ӟ�[���=�zBa��4���6�6����s���a#Ao������R[��u�չ�i��Tl�	9�h�o@���]'�rMF���;�Rd��r�p��ȹ�Yq�7���W���+�>/��0��:|��
�y�/��!�~��B���������*�^;;{�7Sf�,�T�t�YI�i�H��<����l��~��~u���"����~�C��s�����raG"�収\����T@eRÓø�Ƶ@��7Iܯ����q�]��i�/��`��i�4"2�9+���o�"�~���3KsNl�N�{޿J�n�Ҫ���Ŋ?*Sۇ�-Y{D�J�S]t����V����t��{��^롹k���<���n���[���S�}��?G����K��Y�A-���/%���>Lx�qw�U���U�u�$�֟sӽ�`A��k�."b��b���BxF�W��4&(�5遬gۆ���q�����iA/maTsk�D36���5r���]ws�?Z��s!�~'��ƃ>Q�~��\�5ԨO�Z����>�s�����׵���j��;s�O���s=!����o-u�2~�A��Ϧ�ɝg�{�qg1i��L���ϩf4���&�����7�֗|Ci{�����k+�,��5Y3��ݏ��qL�1�v���<i�e�<tD5�^)Ẳ3�`N��ްN
���N����0�3 ̺�=9�oC�<�̌ĩ�WЋ�*�!C��4�m�n��{����9�����l������a������O�mж�.���0�U!hJN8~Բ��2���ݓ�fR�{銇��O"�����s�{`��`޽��	��#\����x�o��{s{H<�Q��9�b��ᩭ������Z�DeO�m�Ϸ6w�J��.�w_,���U9b��7D|�ĩ���lv.
O9Q�Fq�mM��C5�ʱ2�t�\e�+�_sn#nq��

,�qe����y�3+f��2u*��2<�
�Uݴ]�����Ɇ�E[dZ�&d 1��1�����}T��	�ݧg4j׎y�<���3>j����k�:y��x[E&����� !��-q�n!�S�O:�^���N��D��+��RJ�
~���a=k���#s�Q���/O"��ЗA�mKy��I��X1w`���ft��Ɩ��3Q��Z��k���OBK�cr��V����f�AeB`cl��kݔ�Ď�=.K�~n	AcCT�~is�˟!��,�B���םq�)��a�A`^�B��Z[�����si�F��*�����U�nr��;U�P��y
��py�{w�p����Aa$�����z��޺�9���8x��.��Xo'4�t�������DV����9�G���m���O�us\���-�zF�tɇ^���=��"�)aԱ^�ޱݯ�F*�r��d��~ȟ����߂�jzuxM�*-��[˪��j�7.j�}xy��}�-.p���q��Q�|�q2	��%���(�����m/e��gv���B���������E�P����؟��m
{�|�T_a��V��<[;_do޺�����]pN�z549G{���&�їo%,s�l���	�2�mG�4��w�B�<�kk��U���i7�Xs��X_��y�?�{�xN�bD������!��(�H�) �psq��wI4
�#|�C-~��/ٓ��pgu��ز�����X�z�S���bHQ~Y��Ϸ�U�"37��<�,��/�hj8ٴ���M>����㽾YƂ��LV�nwM_vj�H^�7D�i9�OZ�fHX®,*��{��.����3��nv��ؽ�>]�4L"���^�f}�r5[����ֽ
�̈�q=Be���ݽ8$�;P���\;�t��Nၰ���RIP�s�I��]���8v��lS��������囅��%��.6�}�f`��`}�c;q�b��iC�>��Hlǁ���q�!l��^�;t�ܯԠ�S%CE��Ew-1jɮ��!�E�|��S�_�6�� ��1cy�s��ꕊf��3�t������O���._���h.����.�\oc,�l����v�V&{�Xܬ��^G�9���u����,���]�#Nl�v��7��mY}��RB���W�(0Y�.�z]⢎4��G������q��t��+�j��+s��[]U�B��$�{�0.������������8���.K�Z�]]�)H&�������涰�����8;@wnk��:��r��>I�L��'i�x�ޖ�зe\dn,��m��)�1�}]�˸ՠ����gcú�GPm�Y�9U7X�n����W����zA,��m��;���$�z�7���nu�gܨ��?S;8g���g�u[���J���#��d�����^=��͙~�����gc@:)H�e�y��}�)��H��;�HCd5�la�G{�.��k�D��4�r�Y�s:�J`=�"�t!}i�6�wn���uv��@�3�5���HO�����S��,*�!�-6k޶�~���Ã8�=)���E�)]_!�T$�؃�ޛ�s�ȏl[�MT��յ��������W#Y��!I3赲od�Is�v��6l��un�VeE�y��1AR���[�kq����%p9�k�Ъfx�}Sw���v*-^MTa��v�y<4����pʂ��<�{���}�~�'�Jq�t��Pp�hF���݃p��BIsv^�#m;ޒ�Z�q���Ua�����t�E��8gSc�G`̵�>�?�������%��O��A���rߧó"E�������4���.�Կ�j��7�{�gj�jE[t�	-���̌�@��z��"lm3��j�3�*�vw7�r�.x�\zPm;���p�>AN���;Ց��;������ZD�]��w����%�8K)��l�|�y�7��+/��;�7�DH�rpt�W��j��TܥN���ƭ9u�fD�=��ɪ�|�7�����������B;��H��=�h�#)�*�kH�e{wJ�2��igw�;�c/gƛ7�4&#z�b�8U�v�A	�f��Fѫ[W{7��Ygy{��5�a�pa�<^ ��&
��tZ���8���l��	K�SJ�����	��=cM���t�4�.��ynE��'7#�������&e]�$�Gy�L��"x�:&���}|��_��k����~��}CT#�����'�����J
;(��>71c֍�gn΢�'Gp��H��tu����T8X.��Dx��q�e������j
C&��R�x|���EZn[uȺ�T��؝�+i-�1��>ג*��|��y��x~`3k�:Ym��:�:����z@hW����x�ᝩ��m!�3��ʷ�4��n��ӎ�[x��P8���lK���F�+,a@��c$����Vy�_�b���~i���=�S���ҭ)����@Q[Vete��/��-�0�r�^��A7 ���Ӛ�@�{@[Y>sp��q��Q	wV?���:��sy����8�^n�g�ƒy#	*�۹�eL�:�5��)�]����������`��D��a�.��d>�Y[����Վ� H�������ۜ���87h�I'z \�׏Q�t�F�n���bIm�ڭ�6��f^�5ڛSHd3۱�λ�<u����Z�$���ͺj+7;^�u��m��S~)�K�xހ�6ʟA;#q�J06�ГS�th�Ν�3Nɵ�3��7����S�)������.�������Cd�i^�hbE0��E�NA(,N�9��E�{�Jxy���k�Jf�=u|{N� �*��D�e��%�z��ѕy��mu�����lQ�;i��E�<�w����&
U�7���F�?���g��>�ʊ����?��<��r�l�#z��N�������L܌�Z���`D���~�y�H�����UTt-�_���X��s����#��d��ƱOM��ڶܱ�kR7c,�֩�g�:��b<h�!���ˁ��}]�����������}�3ϲ�N�r��"���w_uwl1E(������zҭѱ5��;�{���Q���K��7zwE�q���ا��gAȮ��R�rkr=��y���1�G<%{�������E+�4��k;����(�_��)��<{[��c�T��\X�<s{���G�w�KR6ۛk=>�vS@��F���~c�c-����[�}�
���JE(2J�Ǡz��q.����Ms7"0E��3w��͌Uꎅ���� 0�q�L���ބo�@�d�V��KO��n��j���A��O�WH���pԎ��&�*�y%>Les�4�vq�.x*���0��b��չ��u.U{m���}�c�[�ayX��^��Ӿ�x��=KI���P�s�	ڄt\�T��]�V�9�����T
�АtZ���0Wa�����`��M�
T����r3q����!D���HRU^�}��� �ܭ�ǳzsb�60�Cz��)���!�(��9�RW���v[�KQ��ܮ���;�g�w����3i]�wB��?r��g�;��lO[�j�/��S|�9u��@Ost5�Aly�ޑ�2~#��?tӛ?���{�<�*�{�D��G�}�X���܏>!��;2{�MT��s�Wl���& �Ҩ�Gew%�+�3@Ҁj�D�f�hwQ�Wen�nU�qyǇn�KF�x8G�ѷj�tq�/�h�T�v�>089k��峽Y���>Ѻ�bj����bo�|H;�����\0�΅�P��y�u�>�a��8��gU���
t�tn�>���=�W�AZ�ĵ����AY���W�X�[xo����d3�b0_@xI��/#)>�g_�;iɜ쳜��槐%���D<�9m��S��xB�X��.���wםf-�s��[��dX{��iÝ׏�i�� P�ߠiݓ�j�Z�#�uݖ����#,��c���+HL�3B���w�':��\Q��#3�j�99�4s�x�Z�j>jl}ԁݬx6	��9Ԛ���YLO_��������{�n���yQ���FF�gA���g�)j�X:[7���F\�E.�ƶ�����r��׹���W�t���A#� �Ђ�b���m��VN'��u�����\z�y�t��$�]���끿�}�O�Y���5�5/��#����3�f�nҫx�g���!! �#ml��t�{���ճ�.ǽi�[t�oirMW�4Uێ��@�n�s(�o�xp�Bőyxz���wf8�����*|�3���j�9���t���2��;�;�rh���@�`��h�3Xb
�;i���p��6R�E�OOKo8y9���h�����P�\u��n�������F�Gx�%IwH�YHP���E��9��f���b�7��ω�yt����
��Nu�w.Tp��_s�8{�M�i�7K�h˕R��Ƀ�0�0G�Gb�nT<����;V�1�xq�b�GuM��Ϙ���S�ͪ/3���Ů�h����3uMc��s�:��5d��*�]�$#xS[
c`#��:L�.��m�����yL�:׮sŷj�,8o`��8��>��xU�rB����˚����w�18�fP�5���59sT�̼k��+9�l#e�U�&l\�s�a!FѢ�Kɷ�2�@o^l�f5��vgFU4�h�1���*NV��0��/u��@�B5��7��\�{�;�������Em��eq�W+-[���	WK�M��Sȕ�70E����HVɼv9�BfOmox�)�_�!��p���@��֑�)Lŧ��zy4jf��r���laer;�L�׸�|A���n�u"�MSab���g|K�JWY\�)�G�� �b�;r�h�e����+��*�\t��e��px���m�3�D�/��c�s�m��Z��˰��Xj��r�RɅn����C���2L�U�Wikc�ܷ�NّlL�޹�p��9qj!��^��@<J<�~��)���ں�
���cvi.o^�|oG[Q$є�ƨ�ף��/���d����M&���a��`X����޺�1eZm����{��K	��7��$�`-������]a;��ZPW8:<�T��`s7�T9wVgWI��Q�,�U{ʶ��,ԲU�v�0y�N�慠uuИ��T�4���.*�U`QwPQE`ȩ��~�R���"ȧE�G|���aI޲�U���)���t!��1��ڗ]:nn�(Dyi�e���{ݗl��MMD�׼��q(jx�Cxe3[]�mT�l���R%�D�����𶺞B*�6�(��gtL�3��P� T�;%���WL��Q�b�-,
m_@e���wU�[Q܃:�$�4��Wm7��o�Y�������tFH��9��T��[�{�uN�&���n_T�?o��gI�d\��t�N�н�l�/���үK� �-d������&�*����M߷�7׍�fs���沖Rց��b�\��g��Ѯ�EU�C7�ַ�8�\׻�XQ����$�Z��KHč:��B��y��1���
��n�fqْ��-�I!p̛uE��&c<n�eUSqc=�\y���#a�[�3+�*L�BPW6ە��d���Un�%���c��d����yҠ}�LoL��D��]��u�G�X�.v'9�Nu�"���v���Q�r��0^����٢#�]垐:�-�fp�("�1{�1��qgm��ޤ0\&��Φu���M��	�S��ͺ�R�q�Ј��ue�MOh��ֶ��h�
���6�ި��z�����o�X�wf�Q�Լ��Y(nA�����L�{)�2�ra�ÚR��`-ϰa$ "MSZ��:�yrJ*樝D�k��i(��dҴ�<s������^�z��ׯ�_____�����v��IKA�4i4|���ERxM���PEA��S�IJ🯎||������=z��ׯ����������޺��V��K�6�`��H٠k��6��
+AF��Xھ�(ѣh�i�r��AA�lh"�������N��-h�N��P�t��Q>;���G�� ���4�$�'E�QC�E"7��<�E�Q��7.TSC�ki5Q��ɾ���YtUP:
�8��P�)ӡ=	��Z*�=��\ˠ�e�m�mZ�h�EE�)u�Қ����|��ր�71mZ~�$)�Fv4������4굶����ւ6�h�h
4i�Y�
)Ѡ���m�f��&,l�Ƶ14ME.ؤ���8q�/�����G��VP��X#d"��q�[ٳ���W��'\|�����&G3�g^#�Mu�3&}>������މ�͇z�O�\��vx���?�ޏ8�p� ��Obacu���7Z�vuf��dY==�^�VM��g��P�c�g'�o/��c�9�%Z��SϼaU�dϘ�1��1��}���C8lZ�9�������4�V�Ѱ3#�������+�h��P9���L�O(93QX㮯��g��uû�e�F�0�L���e�a��P�= r�$i��}�LUg��WO�_/�nԟ50���n���
��g��&XI�́�J�(e�2�[c��o��voMfe1��\����r)�B|����Ğߝ[��&�"��3��������o�S��tk�ǤUC��@��w�PL�Spצ�Fgu74�˗9�y�"�@�=׉�UO�s�^�x������Mr�M�T�J*�F���n�uJ�����O��J��U�L��U��r�C[�QL�Y�-��4�BoJ{�h/��"�wo�VaEb���=�\�tmXG;p�.�����a�R�/:U����G��E�>%���%/Wj����7-�� ��%�V1Nj�P�n�S���G�y]�b��Mn�К_kl�B�d�~�����*^nE�i������T'F��u����#H�ҥgm�FE�n�b͓�{�&�&�R�����f����u���Z�y���;,�T��������1*/��WC	���aܩ�v`n%k
�ڌ���S�]Yt�uA�;���i�q�Sv����
��V��/+�Mꍫ�����ׄlm��$Lʒ:f�)>���G �#�;D^��ʆg*��NM��^�q��X��^�;<�����g� ��!�3�n�N�-Ըv��}�m���H���=�u�3���%$��m���늶�f{��//wuj���}��1W�*��ZS�27/��]��8�ci���07��U��Ө�?_�;����P(FA\�r/ on]�>>�MS�;�+���:�z��oD�Z�U�S��g��C���0.�<k����n��?+�w/�����əG��j�%ɾ��: �v�B�;n=��mYL+�U;ܱg-��³�W\���B���1L�P�ˌ2���]6ib��ݲ��cՊGAqζ�Ԩy�eL���eQ��%�D�!�w��|>pѾ(��y�/(]�6
_�^�H����m���6Ӛ޵7,��Z�UxL�m��*������\{TU��B�%4�ϸ���ٓ�s"�Uv�K�n��ƶ��#�)�פ�yi���g$�$�=����F;���#�o[���Ku�<����p�[���T���ڑ�7@ׁ*�8ڊm�zj�*���<ӷ�<C��)�'���
~
'5N�>zM����H5Ĝjs��3�M��ɜ��X�r��8d6c��
��@l�8lS��`�LNFl�^,��;���Ἰ�J=H��-sd�ʑܼ��~��<<�v�Wu�>`�#5C�v�ݾݝ"2;�s�Gu��.�V�k��~Cl�'&(�qy�Ey�frmm�c����o�{ۙ#��L��qJ�L��%�u�7r{��B���*�����#(��8\@�ہ�igC��i�u {��;��ҹ�{(̽��Ռ��#y��e��s1���ZY"Z*Y�˫�_��ƇS �Pd$R��3J�{�|D�eT�-1�L��@ڂ����$���f��N��ά-QH�ڝĪ��}u>�c��Q�Ӱ��5�޳.Jy��n��+� I�n͏���^?�߻�e�Tn]ʙ�� �v#�F���H-����
g�Q{�O������Er���z�7���h�s��ꮽ��Ѣ��1��Rw/77#��n��ʝ{'���%�����C:#����*��L����=V��v��~��Fe���'��!��G�m��q�}���2�3Y����A7��6�����Y���(����J�%.��U���j)F��em-�Z9Ń�窕Qk�.=R4��dT��G��Ffn!����;w'V0�`(���k�'���p,Bf�
���|��Y(�f�vE��8ӎ9�[����'���?�΀�܈HW
K7�j,=���iͻȘ۫=�Ӌ��I�	��K�j����GfD�������8�	m�[���z��zy���$��T�L���U9���>1,� ob�h���ɧ�.lc�K��x૴�	Kz��͸~{� ����q�S��G�;�73���;g�$��l�*r���-��jV�p�$;����rx�Q�[�whޙ�;���Ǵ֘2�tYϮ�-��{�Ez���?�;��,�����~Co�n8�J�a�)���z;c+����j�v�okz؎
�)�I|#m��z�[令a,����5��б�{q��~�I�oޢ,��맟�8D�2�vU{�r���fHx�f�9ahy�Wu\��!��@2��8f�d0K�Gb��J�`��Wcnw{��|r��NwN3hn
���+
��VϺ��ӣ��F���6`�v#�Nu{XyG1�7�D�j�x�Oӕ�FH�} �4l1���~�+��䄖�x����0sOoU��p2��d� �c�Oi����OJ���囂�� <U}պ6e�?q:
HO"���:���L#^���(��d����w&w����5!�h��x�����<�\zyQ�@Ÿ�8"�Nf_Eq�ɲϯKӮ��}D%w&��2�1"��
w+�.���Sy��>u(��ak�L�&hy��C���<>?�7���찥��k]�+O�LӎY��#��f�r�b5s'J܇�k��#�[{�+X�,�o .V��v/�v-Av"�DD�2lxm�v��-�[�egJ�p�DVqMn��v@��>���|>�Q::#p����$wu���S�<��K!T�?GJ�YV)�j{�]�G�7��<F>�u��UhʯB7>/��7V΁9�i�~@EQ����p��M�a������� m�)�+ #�ڊ��S���+�d��4��EY��*7��v��Zp��!fD�=В�0�-�$�����%
�=9���gj�5��|5��?.��
r�/{��#(��^�.hܾ�������ۙדu�6��C��#V�3=����������t�l�fk���ԛ��O;l�� ?�i�4�vw����x^�w�{��#�c�Rn�݂��;��2����Bo0[����,s?ST=wn^�-��.g$j��;��^J��S����O��#�w3݁�HuI��cW�6@.0ߕ	��ռ�x�׻������m�3��Y��-/��\��>n��CmR��8��
R3|��R�4��lٛ4��|r���}�u^3P◹��:]6x�R�W7o���I�r�����"��9;��#n�qA�H����<�Ŝ���|��d�����V�Z{�㌵_Rb�(�BJDdM���{�///]ʴ��^v���Ȏ��c�^�,�3`:��\�{Ѹ�Qv�L��� wi��d��;�F*;����̡r�?�؂���"VUE��3���=��L��J�����7��,ߪp50[���t+���%QW'r!hS7U��q{�W�ػ�.�w�.(�ȴV��YA�;!;Uw�CD�P����דO\c���q7~\���U%Il�X.�@��p�\`:��5��"�^t�_`�NT� Yي�(*�e@Z�I��vd�Ӗ�\���L��U�F����tJ��oXW�Mf��H�B̥A#*�#<ͱ�q!ʳ�/�F��H��=����h{�sR!{�;HmH�tbd��m��T�F���<s�@����:��
����HW��P�s��<3��k�W^�������٢O�l��H'�Q8Fc��p�z� y�#q�x{'.���t�u�]_���N��v�/�A��X��㎙����7Y�V�9{�H��֯ha�X.�0�#wN�������sU��%M`��2�lK�.<e>����r�fHk`��EѶ�dO8�V�l�닂�.�O!��������6�Y���~��o�gL�5�9eƾJ�=��[���9{ө���k�{jkz���J/�^ccdm�����R�K�ucl��ȾX�:3Z�/_U�U�s�1Ӳ��tvUw%!^�%���htx� ���ގ����`o�(�T?�E��,�������T���D�d̼u1����2�����<�����Y�l��%4TjS�2���|�z)���~������]h�e��ߞ��gWu�rK6^�h���̓�o��7��G8l#7?^��rr[<tQ�·�dl3�Q�}�Cͪ�[v(���3����Fm��̲�4�]����e
ߖ9�,� �@���7<� 2+N�n�푃����hע�de�(���U!>K�
�Y�jD�����e������=x���ꧪ,􈺁�+�}>C���%ʶߛ�Ay����~*��;�i�}�3�7���o��{��ڃ����}����^yPW���۫L����8��$�E
J�^wX��
��zom�r��
Ј���g�ۨ�i��C��b<��»)���"����.�Os��٢���ܞ�������i��|g"�������>��> Y��y�t�FA�p�z��E\��Y|-���W���P=�#��&���:C��9���,��]u=���NwQb�+�%^��cFp>Z��uٙ"��'��*Y�9�8��;`a���<7c��7$��7�$N�V�U9��S�iia�3F�j�.>᫳�����;�C�!��m�t�'o���J�#&I�)Z_d���X{�H;�FY���ή�cH6����тE�h�v�r�[�&���S�ь�-��l�C�L�$>���AS�L���܊C)\?5'h�3�<���u��EH���<Z��ka��`�Lv)��' ��BG�&��p����ޓ�~��}S���G3�`��/|��D�O���9�G������vz�ҍ'��=#�tw���8p�uzv��W��^�Al�+&1;�C]�F�:t�ozRJ�)\W;���D���JΎ��n�K�;����;�S;��+,6�(%r]��.��&,4���ݡ˔���������#X�[t��{�P�=1����9SEw������)�1��|��
2���]���|��d�� ��U�~������n�c#W��Q�[���3��a��O@�<U�&���_�_���H�X�,l2k��/�m��]��]�
!�Texjg@�x�0���&��33>WvaQޑ70� �U�\��3�����5�rej��_���/ƺcd�k�+
���0��w^ңd�B�$��=yjni��Y�
qA��uW�m�}�	����}�A����䶭N�>�����C��".��̋g
����6�S��u�����i��T$�����%A��frۇ�Ϋ�7�%����dǼ	�\Dm�P�K�ɒIR��VI�&�}��x�3�9������b��Gg�����6V�{����ESVja���e
�������U��7�7��	��jt4?��&5m��:��7X:����~�;i��Cv��Eb�N�����sE�'uc���i�n�5+�������x0T&�"I�n�zg)�ݥu)�ݱ�%���L[�3�X�>q�Qؓ;����6�s�ˮ�2�e>�\D�r��N�qntՔ��C���{.1��Ҷ�!A�� ��]��G���jẵ+�մ^ոJ�e�b���.�v�T�J��4��yc^�&FE�ް (��ծ}P��O۝����o�4gn]$D�%~ݹWJr��x/�.N��h��"�p��jue����\7K5��L�p���/0L��dM�ȁ�)�[bI �i����?>�B��{��+2e������2�����Uxh�E���1V(���泴h���(���7��W�\���|Wt�r���YG$ti+��E1>iwطsV�g+r:s��s1�D����Ž\bS	Ɏ��-Sǂd:e�4EXkCʇw`4ղ�h:_7iYo��L���)�x��o1�Y��-�|���n��8�I�/4,������51�bT�[Kj:1��p���U���.7Y�޶�jڌ���۔��77�������fkoZu��T�$o'7R�pmѢV�t���wr�{�/g	vA�[C���5�﮵��*���p>�֡���'�}���o1׹���aT�j��k��NZ�C=�]|ꞿN��:N�2�,Ԡ!_!)���	;�k.`�C���ijzN[�b�+������F���SL�a7Zٗ�T��zz�犏/2�jm�c	<t���i�y]�Gb���Efs�;��Ť��U�͵u��gl]�7ڗ]J/��\É̔B9�����5e��t�ѧKZ���87S&p��**�T�y���� �Aې��8�^s�����X�ҏy-�T�"������ST`�p^=E���-tkoL��6+��$MY]�0�ͫ5���Y��M��76�K�M�qP����V޳V��HYծ�K���@���Եu���Ft
���˨<x)��l�P��]޴�M�ݴK����\ז�9�o��u3)�����\5��v�>,᫠���tŐ���^�D�zV��+rͦN�b��i^�Q�z�u,v�-�峘��oMbܫ�Φ�F̈́���<���z��/r�M��&'�n�ܵ�5�����Z���iՎ{i��,B���c�`]\�����<��9�i��	�� �G�ߢ�{A�/����dܚ��Ƨ}�IG[X���9�:u�n� ;BX��<��k����q�ެ�[�7ݝ����_x=��\;�M7��i�,��U�ėVv���.vKn1��˛�$q[[Tj���8���z�u�KG>8l�}���M��Km�s([�<F�5�q��[&®�q��Z����% ��z�QJjm���`ˑ��E�Φ�b�/p��҉N���7j�"�WB�j۠m��E�l0S24�;(���h��J���N��(�1A�(ª�������D2Q����, ��?���$��A%#TU4�SEQMi�tj���ZMV���hb/Y���ǯ_���=z��ׯ������_��~=�(�����٬MӤ)~\�4�UkKU��x�}~�_�_�Y�ׯ^�}}}}}}z�~��RQ]�$T��\��RP���.��9q��F�B��E''�r(1�m���M�4h6ƊO����3�Mj
j�����m��j("��)�Y(����)""'lQ'��#A��HkcA��ɍlUCN�h��0m���J�������m���֍���3T5T5b̚k��"��3�Z<KkY4�PZƱm�62�#F�mhjѝ�V��d�bm4ל�LQ��[9�Nմƈ�r�6��Q�cb�A��G�޾;��h"�5�**���*M�I�o �U��y�lhu��<�U��/=�|���P��Zγ\k�i]�/)L���sݵ�ظ���4�^_Y�
j�d��ʘ�U6��%Ea�U9��T��Q�hQ�$Y���//?�k{o#��<ls�c�7[��(��t�=��殀�d?��U4\(��L�Wq;�{�G:դ��(°0����k�.N��4y�q���~�

;3*�wq���æ{h�t�����"fT����I�@�j�&��s�������w#Txg�;��nF⭡�6��l��D��J^��g��8�����Ëf��h�{���Y���]3��p&<�fDqX_7��g�v^qLؠh�u�����{pV������;��b�³X~J�h�[�b�/n�H��e���X�iΉ�#x��pR���d�rЮnI`��LK�d��Q�3$�����/ �#@�B}ȴ
�S�Ng%�s�!�eUglȭq3Y��V�7g�sO�A�u�w�>�()*}��:ӽj��!�Cf��ת��kk(��d+�"*�Ϥ�5�P2)A�֨�c��U�J8~]���!����(���aP�+��/3��1f�e\<�úodr�Z+Y5�i��\�M��)d�ž	��5�H;�k��|o75d������M�|�d޸m'hg<���frN���Rq�>���|>�w|��p��6�@G�B����:���|�^#�0��2�v�H���x;wu�Zw���ח|X+����8@9���^��K�Ct#-wt��հ�{j͘�����;ʺ�ISuuK�< ��x@�a�MJ�1���c�j$�V+޾箌���6ɒyq6w͘��lBҔGLK�FD�i�Y�#O?.����hK��ص͒;eOsp��2����}���c��Gk���S;kbGYJi.�Ս1Έ'o%񢡣`��7��P�3�C���^�"��L�t\�tvU{�)W�c�^6��Z�5ʧ*����ۺ�"����pހ�"���YU�=��տr�7Sڧ�k�ӭ�zѸ�ɴ6�l�m�pG]��:��YQ	?Xǜ�Ǥo7�:�cO��U �;>'���`l6�i���W6�inM��\(�t�H1p}�ta�o$XX/�2cZ>�ٷY
B՜6V�n�����W�U���)_A'}����������&����mW[��U��V�*��T������-SP���:�v~�y5��C]�+���K������˒1��b�O��GE�G��wb������9��c�:��6� ��	����Ix�!淨f(�_���h(�y�r�U�r"ƺ\�j s�U��ww4tG��{�/7�q|OW���T��E��W�N��VA%��f$r{���m{l���U="�}��ѕ�WW��9���*�`8�hY
?x�آ�*�ɂ�l����&�]ak+�b~�HϢ֯R�%�µ��c���n���<@�M���ʨ�d����dR�r!!l%�4�zeQ[a����1ٚ{�xϛ�$W��L�P�MS���{2$Zh��U͕Aag��W���ԗ�����y�۝����S䉖��T䛨�xޱ�ior�5����`R���/nyQ�\l	}p�)/�[XT�zK������=�]ݓe��p����zD.�>������ݞ��-��'#\Qy.N6Z�gN�>R��m����O�n�Mʨ�竸K$$T�c�q�7�ݸp��²v�4�pr�omI-�#�V�����	��bӠ���2��Lt�%�EF^7���&kKn��r}��|�ZtU�j`A�U_�����~~����6��2.�7 @v�9O���^�+��}z�rO-���c��;�%JG&��?O��U� ��g�L�1���5����cI���������ܫ64�}2-�y�hx��V���\��X�6�go��fa�O�4���*,����,�{J$'��<};B�q��{,�c����3���7g+<�vڰ�ö1�bg5��7��\xe�h�2 ���]{��6�[A�����:j��� 6����t��Ψ؅��;���2��>�^&�I"��q��5'���]}3՝�EШ����q�
6Bc�j�[�o0����j�n��V����d����
>�ܛE�yz���  �����
�eU�;Vsw����K/	^�*Ԝj��q.o� 3�^�c^e��U��w���ئ�G�޷8+�)R�.z��>�ɧ�l�gT�<�"��قP�^�����Ђ�ϻ�x����b
�gh���]P�"˷�ȋ��K���Kꥬ�tԤ��B$�����Ås��Z�n T����1�+0��am���7���c.�0�<�J�-��s��nP҅ڑ�eL����h�H�	���Ęr�AD����|}#�kO�����[��x	8�!�������kd6�g��o����\�UO�t��<\0�X;l`�F߻u��3���O���/��o�o�RVtr��^NY�h�{��"Ei�=�[͵}p��/��x�kLJ�y�y@�/��vL�;v����ڋ��w���7!����*@A�c�ܾ��E��\:�wc���}��$���H�Ԛ��5Z�'��7�J^*��Ou/����;��ш�Ĩ�c�W>�4M�j}ƛ���0��Grw
vͨ�n�:9/8Ԧ ��u�co������S~雜���!�h-�5k�u_w��n(�� @ˌ��C�l��ygr�'�ͻu;�8�,��X�tn@�p���P53����홀�+��q����Ǧ��usZ�����z�Pg�g��0"άߢґ�퇬�>��cc������s�fc�a'Z�䂬.����V���ȃ�O�e��veE�:t��wo!�U#�u�,�9�<�n厛�YԹ2{�Ƿ�)KZ�R�h�4���h3"�ʃ�
��Pݝ�*]�y;��-����/�<�����{��7�wO^auGvQ=��;�ا����;�]�)���eF�^�V.���C���qm��~G�V��3�
�Z���W�����Pd�3!4@�{T�uZ�ٸt^@9(�_zz�2�@�C��)M�4��Q��u1Y9�S��Z�ͼ�5���;��t�u�}q,:џE\{Q
�P2(2OZ~,��yS==��ݻ=Y���O��F�W`B剥^�8�2�j�3���44B�y�����0vd��@�����y�9��T��b�G m��tV
��i��=W�{��8`�3����^�U䒪�t�K�X��8���#'"f�anV�t-CxFRW��ƛd�<��Nl�dO��-�,��]�y=��Wy[����/b��={[xΓK��[k�3�T�w7GH�0"�S�֦ܮ�Tǅ\x9��_�wl���޲��K�ucsvu8������E�i;Z&_`]լ���Q+j��%�U�LT۾�e����FҒ�v�Z/F�V@�=IӎX���������Lz�q�	��ޮMդ�V\�yJwnE��q&N	�Q�����>o7�/����ם�ԙ|0|c�ˤ=x��O�M�����,�3F�֗cs��Nk�y!�Z��oh͏pއ	�m�Y�ǅvl�.I��ĳ�d��UQ���ɍo
�L3Ͼn
X�8 ,���SQ��Z:N��[�NooQ}�D���'��_�u�<�#�6�5co5g��U<Q���9�n��;���"�@n�����`�<4�%�zX�4 �wb�xֈ0z���p�S��C1��������Ey�r���C��Yu[���}9����}ɝ��`ȁ��=�5s�V-�|A*P���7���8�vLzM�uԌ�n��T�K=���)��߫�N{�䍵U�\CT�_dnt<v.�="��'O\z�]x^��!\`;�W�{��A3�?	z��ڋi�J��t�~�M�Vz~�BW�xd�:��(6;v�[�Қ�e*�{�X[WeoH�X�Ӿ��'��ZS�Az^��Y�ҕ����:�޼i��}Z�
��������A\�f��٣��-#zŶ��g��8�Z]�;�ȶ�P���k�Z�oj�ي}��&� �-��"�e���W�������k��pv��7�����bL��yG�r�Ohqp��h�`==Y�[���:��C���m��G$J�RD�ml�e<�COt�w{�~��뜉X������x�=PF��7L�����x��#Py�:T����kSng[ᬞ�Piq���!��cd]�]�=��2ى�}�=�*�tN��z}��N�7!��d��o;���&�n��k҃�+�m0`�b��;��t�Ӽ�k���*ݓ{��2���uyu+.�O?ev��v���9]AF��	���aWG�VϺ=O���h�`�=��s��#5l���4���Ư�d�XmU֮�ԍB������ov�&�ɔN�Z$����ή��b K>�*C��P�ؼ�N�d� �b��_����^����,/�#�C_E�uF�U��7c�̶��&hB��e����@�UHʈr��+/�>���ŵj�
#x'KI�v�4"���a�uc k����ߴA�佮��wޣ�uM�+��wzd��|�mh��V�\�ƅ�]j�{v��O�dh�T�����n����P���!�t$��ή���u�	��"�bQ�A_����쑍�8̝W������p�f�A�Q��4+�� !}�S�O�j��ɘ����^�9|��L��i�״����Q��j�;\)R��@���3uWћ�gN��������k�X�9��t)��K�Hc!�,Tb��6lf�Q�'�_k�ج �z�IsՁm��Ӛ��n��2�yj�f����J��?t ���[-�=Ւ㒸��1��۹��e?ӹ�ՙqDe1��q\90�q�2;�%`1��th��t�cG6O'8��?p�m��>^7��j���G����׺�q������GʀӔV�R������S�� �n'ѫtf�*.ĺ��������!z��׀��=Xh��%�A3���Ԇ�m]cGN.ާ���$��}]��g�ˣ|sTu��+�ƙ���:����wE�s�gV����i-?i7���ov�}\CN�"+��u�Z�G�pa�N��N�*f�[�SP۴X�5w��Z̙!ޙ�517�e��.�V�Ă>f�ܮ���ē��U��?��׫n�<_a*���3���ER���ϯ��2h��7�πa����z#5���r]^H��
�n��:�����\sy�p�3��Լϸ���`��|����4��l�s���S��yE�x±E�WMD�;�u �8������>ِ +���|�G���;�4O\Z��+�Oڥ��_G]&��!n�uzFE���j'eD���sL��N�?7��Q$�sAox���ǣ������9U�tEdM#;����#����R�wI�Q�
�$r-Y*�)��*;:�� ۆ{n��a����KU�P�m�jHMr<i*H�fҋ��f�-�3�6F��1ݭ�l+�`�]���W��X	@ȥ �}/���1�;g��	��ŗv�i��2�@���X��Kw��D���f}RdF^D�tk�hY�;�}g�x�.f��N���'1�U� |������$�`�֞�&f�"v���ّSma�����5k�&m�Dʺ���|��i%0��c�g@�VK���_a�$���^Sa<���ԁi�zr���*Q��e���~1�6���Q�4��=h���Lu,�T�D:�ҥ%���[y�ii��Q6�������%�-������m��>�6�[&����ܠY&��Y���2iF��}�r�I��ē�L��}y�G�쐼�!�����SsMT���a��\��
&�m�mY�[cq���-�q�n�H�̿�L�:L4��xėD�[�ٝ��k���#9ƵF�Ad���Q5K6d�b	F��6iT�eĮ��U1wU�.Q��ԒsӗGF�!N�3�N<��qFl[B4YF�er��ʬ멦��-b8\A��b�n�j�=�m���#:z����MfajW:����E��W��c&oN=Ł����fKܾ�"��M��i.��Ռs�Hes&�S�s���<����A�7w3�Hv͘�s���/�i͟��֚��s�KM��m2�z�2�jh��}W�����E�*�4�:�u.홊t�1;7_b�](��x��t[��gcZ�(p_sI�x�Wa��ce��z�G�3����ݏYӁ�Ch�l���9��M�:)�B�y^3'���Ӳ	D�����'[�q*Q;���oWg�5w�ҹ9bA!�"�P�%��:�z�m�@���BW7�ǔ7Xn�eR8V)�j":uJ�&��T��tk��D���8�{�ʗQXNZT��gI'g3\��qň�%����U���{��L��|%�-՚{g��݆OI����֑k�īn��Y�S�$>�؞Ɲ�� ��;o0,�h4�#X��m���Q"f��,���xv��ť����X۹��0d���s����ޖ�.:!&��3�jY%����iO{����E����8�Ab-�m�}�V4WR"�t3���8��r.T		�m���f�Y'�]�[L��N�n���إ[�Zڴ-�h?�Ӻ�osc{ZN�&��.�T�#�n���=@M�\[7�Uӵ;���n�}f73QU,KZ�{z�^ѲM��;�F��9�j�}��2[�f����X�J1E��5j[�@z��'6���E:����U�:��Mx:����iMn:��֜�%oq9Yު�er�针.�F@��]�&W�q�J��g�G�]�+�w#�v�R�8��^�Czw[�B���Nخ%����o�v�u��Jv��Pڡأw��;�Wv� V>���a$�R���^$�f�vɖ`{���i�vܽ�ӹ�3T�W��QoS��r�[�u����8[����g�ՃV�M{O�/���C�_w�:�E�NÕ�0.kQ�k&(���)�i�����4O� �J@��ڊ�h��-�
�5��&(jj��$G\珯���������z��������ׯ���>Gg
�֦m�kI��Tm�*(o��5T[ѭ#Z�*}~�x���������ׯ^�}}}}}}z�����%m�h��|yϖ𱍜i�E����v1�Ӌl��V�I�Ӊ���k�<�C��sf�����Tlk[m['bؾmr�T��cXkM�C����kF��QA5���\���8DM�TPQDQ^mZ�j����Th�*b�ŭ�\ɽؓ�k{f(����.`��X��gUTSF���v
�UU:��.�Ѷ��k���*�/`��-�5<�6�gP�ܓQ��E����Ѩ�.&�"��6SZ�*��QO,F�M��1EL�E�.]��TME�-yi�*������^Z��4�V��MI���b6vƢ��H����F\9�8<�9��o@��cXɹ��ԊSbp��s~������+Q��L�sG���˹Y��\=�uNVVfyy���3{���oW��>��2O;�%T�qQ��X1x�u)�e�֫��w����Ű4����t���ƃl���l�_���N6*f!��Xf�H>�t
~�gm�2��'f��\��Zݝ���h��D+��Y�����l����҄tl�6������]Հ�k�e,��vl����y�(P����kbe��W�ڋm!���<n#/ʀ�7t:;*����E���w�0�t���9�['iG�VN���q�`�7��FDi�G�ߞr[�?I��3�>�c���!ͯ{���md������~�uce��+o��`Y��mov/G�9*׾���q}� �|d>ё�붎d�ú٢j�%klʵ��gK�҆��������4�%�g���5e�\���Z���0ff��6z����)��������p�ܲ�'�O3[ﳧ�&���5�v/
�B���i߷o�ǯ�W���e+�t{]�^�0D�C�$dLc]�Q�KE���Q��a8�*}��Ɉ�}�|�H��Ő	��rК��67!b��n�ft��oPh�y�od�Lj�^j���:��'�UIͥ��y�7�\E�&3�ץDz�Dx�0� >b5s;wk�h� �z����qj��5��n{D�۩���.��`���w<��3�~�!�N��Ƀ�=���%[���m�N�u*�G3�^=�q.gu�v<w����4������|��LP7�Ux��l���ʫ�Xv<��xi��K@h�;L�μ��˕�n�Z$enD�c	RE1&s����[�Q	�=%�u�y�[z�Typ��o��,�A[���a���ܒV��
�rQn�b5^Va�3�CZl�S��p����mW�� m�*=+�U��4F��4i�(���َ��t�'�C,�3�ຄ.�F2F�5Ӕ�%\���mŽ��Ž��z���~�%�v�k�0�DF���AM	��d<-g��s=�k9����Wq�Vwk��Gu�w�Yn0C{@a�����nm*z��|l��$E�W�"Nbuv�)gZ���1�Y$CY�{��=1.Ԍ(1ۂ�T���b�CP���֝��|��	5D7D�B��N�p��Fޚ���w�ۨ��油���-��{U��-�U&lVs��Y"���<�f^L���7�[�SZ�����@�R/7��SLw�L�i������,�'L=�4�J�tճ�ݾ�UfD��6��^�`L��v�Î��P+�IsO�l����f�aR��ҝ��v���x`aB�F30n@_�w-�Yv�n2�4I���A ���
�S��_����;b�y[�v �,ꍈ�GtkH�b�N~>�+�����S6|��_�$����痟U�pA�//`3��o<ǹ�B�`��?~���S#�N��"��G;�c؞��<��zЂMX�q��jfwj�Y���z�k��5Yܕ��@�� �%��yj�\߶["\ZS��Rv��ѝ�kk:��;�0�����v�"gu��Z2�B6ņ�C�]��b�ʶft϶��D�(44�6���ܘ�r��t��kp6�g�=�'���哳��Qs�z̛=A��f�����G$BQ��#o�t$�Hm�����Ș���ߞ��Y�
u#���Ye�Hp��E��1�e0���q��͸9 K%o�=��"H�{��yX�퉬u��/_J_�/��Uh&��E2ҳ��뜲9زR��-�Im��p�o��l��Jk�T&깉g߾���o��9�����z_� �Sep�u���:+jx(�E�F1ž���Y�9GM�:��\�RqH��@Y��;��1m���,v��ͬ��:�b��Ӫ� v�O�;;�j���Y��J��~��R<f��L���̠�~���c����-��j�(Ā�O�ݓk��,'*c�;�I>��ڴp�������ޟDb؅��}�)��	Q��
���Ǯ�5e����wS3)��8�4b.2�/�η��L�Zʣ��)����mN�~B�������X��;}A�3��s:��p�lϢ�N��f�ۨ���|��t���8�n�#��s�G��u�q�·l{0�þ�s�e8��z���><�(a/��Wv��sO4�G^_���P�s<dbn�UlMs>�����.�盃�����y��T���h�cS#f\��CҀ������-j��
;X�q�ܘ��F�qj�Zڑu����U�ƍ:��W Fp=읚��E\9s��̗kB?Y魢�Y<ڝ	�9!��v�H^�H�nu��k���Oݼ]tj6��p73+���O�87x�S�+�^�x���g7v��w[|4t���� ��n�2C�4������3;��(�]f�L�\v�n�
�rj�TO��j!Y(����ɢky�N��$�=�^�un��P}�=��?��;ѧ�������n�Ʉ��Vn��蔬�4��^�%�V�Ϋu"����5"U�Ӝje�ʝle�W99�f<����Ӡ��-đ�N��RIU��zu�K�6�#���*�)f��n�����3���	-ˍ6ɒyux�-��ƻ>j�n�֬mPv�Dp���O/�MK��[�6V����|"�;VM�|:o{�Pۭ��?�̆�";dA���;j=���)H46&eܶ�]oY\��Մy����� ��.�<d�S�k���2:��6��&�}��[y9�Û����eg�VN�x?�3�$o0(؍�Y5���py}��q*vg^�c��)8{����!���ٳoR���ki�t�X��יZ�{����Ey����Ҋ�=����up�ZV������H���rv�]���z[{�SB+�LMG1F�g!��yQ���{c�̚�j���n����h���������Rڴ��7��F�}[@�T׷���m����.��N�H`��5�5��{���]@�F�H9�����*�g�����ca���w���W�-}�6�}!��P��ku�\_Y���;����a��F]߳ �u��7w�-�l3�QZ���^i�����$w��m�Cli��ܱ�xٙ��� Z��1ngCXP������]�'�m��s�s��2'W���X%��p��Fu[���d%�T�a�k�:�b�����E�ߏQ��S��*��q�����20��`�&pg���͆��ؒ���#�S�-��;�j礹�5㹝���4����g�37gwo{�.�<!�p�L�xs�A"�9&�)gSm�8�m��ǥ�t�Gl^0��M�T2Ӳ � V�����vL��$�7/S/L����kQngs"��=��ޔ-���/��o6�,j��}��a�	8M|����	<�>�F�y+(t�7�� �I b�����1�����1"\�w�r�Y]�;ڸ_I�y��\�L<n��,��7���u1%���"�R�N+d��dN���9�дIA��"�}���i+�����_���`��`�:iڱR��9A�tɧ�}���1���G��F���ď�d��!�t�t��==즗S���i
�wQ�Ÿ���od�Ge��T�^)Y)%�}̒�q����d>���M����k����;���9��r 3���o�ҥ��h�o����]���ͻ��.���5"�î�V�qa��'�@��=�h��J{OV��S��h�l�.��p���ʂLӃP.�9v�St_ѝ���Qm˷+k���q}�Shu���0#|�r�3F�H
FNj!1nU�O��w�����pQ�V�z�:,�xT^n|���L�Ǫ����sߒm��˱y�m�Vodo"'�h:*��O����'�d=��p��۪gF+��n��~Kܰ��k�O*�`4�i��#��=��C��L�)��_�H,��2nav�qY2��{qr��'gK����D�W���&��t���{Յ�r��̺Wv��N����� �yr�E�@P��$w���m�nP�ڼs�d�t�M�Ӌ�Nl7�0��:T�٥V�N�/�Ҕ� ;X��*'��lR�O�}_��+�&)�F�zz��SC8���Jm0K��ז�\ӑ�P�]�r�+��#F=���=�yj���+�ܒ�F�J�u�,�Z���nɬʊ#&�M[!�@�ܺ1�dF�����1�rQz ��\5�w0�Ӝ^����Z���fʤ6��ҽoBÓ	@�q��6y���M��G-���][=T����I%s���N�`��"�8%2�s^�LM�윮����� �� �%H��t�Y�#��}N[�5�v�s�,F�=�{�wR9�s�p`�p�0�f��/�;ҵpK�>/CRn[������l��`Yճ�G�/ :�A4 ��Ĩ�aU�N���13f�r7f���^wC/]��;�T<��O�1N̩����x�DԽJ�7ǯr�ʾ�˨&�x��wz�-��P*���)FO��^�������K�ߛڜ-f��Q�M8���%ފ���i�s��8R�T}��-l�=�����:�;#8�>��lL��yX�,cM�b]��-č�;6�L"�;�w�ݢ��'���}G��e�V �5a�yX6m��9�1��dvlD�O�"���^o7���^�̒hguR·�����ƃt,��Y�"��b�.��v�mu:��_��������{�*)�:鳪�+�RU*��<�u\�8��^���ު1۹�6�?wW��H0)}��G�4D.�ObV�'Q��(cU��6�%�Uɡ{w\���z�U�#��w���#[� (R�]ٞݿt<쟅<K5Z�5�!�b4j�%�����ؐ�C��%l��/�̔t^]��vVwk�ٺm���(+�{M�vL�^�s�q�YT��扈��c�Yѝ�G������:�a��QB5�s�o yµy�j��]<`k�λś��D6�*���0fJ�W*����܍V�}W.H)��NXA�ew����̾�;z�����n�IR�$�_�0˅C���9H�;���ݽZ;Hw�>r6'H���Cl�'�P'
�>�W��3gE�^7T��2Mެ��;�u0O+mV,�B�PA}��BY��so[���7{ݯ�V#]�I��[��1H0�O�����lxtL9����V�l�s3�2�k��B�ԕ��:�xGs��@}D�ENO\�hg�úk�����z�����lC���t;g���37���=F�xl�`���+�ڳ��F8��'�l��o�:���m����>)����������tl��^�i��^�,�;��\�n~��_R�ky��;>[\ �lx0O�s�;��#�ь�$L�f�6�.�����@���x�d�0��3H���ѓ$���c��bӝ���'l�.�մOu�ɽ��m�a��jsL�wթLL=��ھђC�Xa���vN#��l�A�'�j`g� ]�����5�;���fjO�G��s!���4�~�tR�n���3���Y�;��w5\�A4�d[���p_f�̡�Mg���4a����撬��#w���Ÿ������V��ov���7.���nv�����(Ǟ�W22�m�߃�b�Y�Gk&�>E�=è��n{��!��@��T){�>�����R��QUEi�T}����?� {��p�@���~o � 3 �
�*� �2�2�2�2�2�+ʰ�2� C
� �0!�*�(ʰ�0�0!�+ C0�C �2�0� C
�(ʰ2�0��(C*�*�
��0�� Cʰ�2�0� C*��0�2�+ C(�0�0 �2! C*�*�*��0�
� ʰ�0�+�C °0� Cʰ�0�0! C*�(��>�� Cʰ�2�0� C °� Cʰ�2�2�0�+�C*���
��0�2�2�0� C�*����0�2,2�0,0���+ �2�2�0�2����°�0�C*� ���0
�� �2�0,2�2���M! Ȱ�0,0�+������fUq(��@ � (�� �4� � ��ʠL�32�0���3�L L̪� ��鐙Qd�Tx�"a�&	�P&&@�I�&	�&�Bi�P78<Q`&@�e&�D�fE!�Hei�` � C"� ʰʰ°Ȱ�0�0/9�x Cy*�a�a�a�`XaV�� C*�ʰ�2�0�0���~G��{�?/��ނ �
*��"�,��ρ��=��z��g���>�����I���
>��*~^T�_���yN<�TW����<AT_� 
���=	����=h}H*��çxk��7*���6�����&l:w�@��*��0B��"�H
  B �  K" J�������H@VT �� %	 � %PP� $HD�  Y@� %@� !D �@� !HP �P��	YVF  eX%Y%%Y�iTB�T�E���Sȟ1AEF!(
�����_������|݁`d�;�(����ou�{?�\	�A�} ���.u�����+��!ޝ95�L���+�EU�C�����W��U�A�BUQ\� Q��J��q�C��@�}�M],p6)� *����+s�pv!Ӳ�UEy�i)�V�g���y���ِ�9'��=�����TVL� �����@Z�c��"�nԡ��a<h?|�l���BWUEn�DD0�pv�<�`:�P�newh���DE�6`(��E�}��<����D;S�����)��uaa�qhl�8(���1"_>y��cmE
RkM�P�!����D�iKM�l���!T ��J�YPf�U*P(J����*��f�R�m�����aJҙ�X�U`٭Z�6-���M_mC�f�*�����Id��e5���e��l�������B��ֺ6��ڴ�Ui�*�mkiT�*���LjSU���%�6��U�kf����ʶ�٭j���5�[[+M�4%�lU)��d�if���k�2�-�bh�%�V��m�@�%Vɭ�gP���6��   M^��:�IVn�J4ݭ�wYU)�]�i�
�k�t�������(n;Ng]	�;n([w]�OWAa�Ol4���ln�
�.kkR*��ْڬ�Y���   8��C�P�v:�S現���2(hQ��y���
;bB���T�Ҹt|��[��9Δ2�nշS��������M4(m�7x�^�V��9UZ�ˎ�u��m͌ƥd�ղ�UV�-m�  k��j��F:��A�o.��wv�ڻW\]�ZU��v�ջ7f�w�45�-�mr���U[N�P�)T�v黺u��\�]��ݩt%�f�M6U3UTkT��  q�GF��{�}���ڻWA�{�S�Uy���X�Qj��Ӫq�p�`Vee��۶� �E����=��QE6�ն�J)�XE����Mm�o� �������t��u�vu.���wU�R�0��MI@܇q�EUa���uT��Xu_Z�=�7�5����P�tڦ�X��-�c*�D�  z���EW1UJ}���pR�R�����Es�9]u�+���	Pwpn���ja]=������TKZ�Ҧ:��Z�M�ZZ�Ydņ�-��  ����A�U�Ѫ�z��z�^��]{��y��)J�)����$�J���z�m����=(P���x��ƒ��M�u�*P�<իMhئѫ4Ԫe�ʯ�  .����%&}���$Pn�[ޕ+�R�t��TUM�n�IRU=�ު�M����۽T�Jνyꐪv���)J [��z T���3]��F�2M��BՆ-P�   m^��	7Qw ��!Y�k�R�JJ��N�JT{�.�j�)R�w���A��{�ÕI@����萒����z��[<o)BJ���/X��hUZV�Rm�   M}�]j�)]���֕��5S�۽W���J{��ޕA[eU���R�*���F�D��S�.�AkK�3q*z�{��D��l��O��)P  "��b��@  S�b� ���%)P   �� �U<�  I�"&ʪ  ��`�7�������%ꮾ���v�Q�f4��,1���yO飌1�5LD� �������S?�?�1��m�����1����`�6��1�vm�6<��?����I���4��#�d��.�j�n`����ջM��<W�&�X�;9Ne,�.�$���u�X�c/ Y[�с]��+(hJV�nc����[��}�u�ky��y�|NR`��۔UM�w�Z��l`��K���Z"o�	N��k7����i�\�Ǧ��x��E�L�zYܐ��f �D�A�+�G6!ً�����������j�o�_K�Wq"t"M�YkH��(�I<��Sl`52f���S3`o ��䳈d�x�Z�mB�ZL/N� az�l���؊4ME��Fk;�p@�*���\
�Z/I;J��;��������d�j�	*�Tpm���l�R���Л& q���
��n�Շ(̠���n���o,QB����	�5E)�.�c�@���u��]�e��e��(JMЏ*^6'��1h�-]��1���ï^�olJ�R�B�-ۃ/Ȫd���v�eVF�"��o	��*�يܺ��d���d�ѫ6��ut*4�{��s�f��z�d�%��DӘ�7�NiOKˉ: ��}�v��0���[����"B�n+����a-�
ӭ���ie�yD��й�e;�\�jH����j
aC���kC�S"f�ArP��2^��Ӑ6�b��D,Qn�hXf�{�I���_����:��:��iɋ�*�ogb�oհ��]�Ž��]�®��YL]佨��@F�P�v� ��g�D��a���7EA�R���UM9Xo���h*���a����[�	J��%�u;�P�(���R/�j�O;׏.�WH6V����-/��մ�o7m%�-�8X%��&�PE�m�y��Sݷ���'2Խq��b��L�B�xEciXd<���R��O��9%���]E���a4t�ѭZ)�m�$C�{W=�ĘZ�cIm=7o-��<j���1=�3�*��;Jlu�3��ڏnM��,�m=v�Z�m���7�n!��:� �h��1w�Ihu�t>]#E%][���u$�!X��tɪ@�W��@���u����4@{��z�ou�P]e�)�"�+3i�K�M�7��GF�.��j�*@� *�mK��'o]/�J�]���rS�p�q�'V@wi-�������F���C7��e�+O�MeŢ]�g&�َ�u����fMo��e�є����-�f��qZ
�엓ie�P��p�32QY�Z5ޚi�v^=.���-4��P�F�B���L��Nj������Lj���[o^x��ãq�l�������`
B�Y+o\���i��`�5I(`�����e-#l�	�Y�vEf7��=PZliʺ7vPm�Z�[��I�t&Q�;���j��LZb�tv�̼�c��
�������[�&,Զ �	(�[�s7[�^�W�[�AQe�ըYC�p�Tp	a�WGM��x�S\�-GW�3\���q��J�4�@%%�=���M`s$��d��R!+�4XkK�Ys��r�V�����ծK®�ڠe�I��xv|ov�V�tݑ+kr8j )\�@��q��N��[b�X��36ƥn�����	1��ʽ��j��6��P�VJ:4ҽtsSTn�H͚��$ɁDҕB��J�R���4�A��1�-�ø�`�"�f�ޓJD�����6���\��Ԩ����B��)��Q׮����+/#Wԕ]<�4Z9*�(L��e�0^��b��hτ�׏M����,�
DK�M�.�w�l�Wu��6�X2|�d�H]:č$�R�[�t�-Ж[#1�a	����i혵�{�������ꗕF�����ԓfk׿J�Ɋ�Gp�0t��4"Tʺ�xPw*�6�V���2 3%M� R�$"R4D�˻�L����wh+�����C�֊pA��[>�1T��Ms)\ѐ�Օ`�����H�[un����OF���/l�Ac�ܙ�I*�ݶҭ�;,I�h�0n�X�&`�w�
b����T[:�S��4�1E�����3�!�u������KY����"x�lK��g6�M!
8�h�3@'$ݼ��Mᒘ�t�Q�Rr�^�N��9,�)Nԫ���9+��֯d���h0��=	ˊ���]&1*��,ǫq�a�5�XC	ʺ�`���ո�ʊ�um,��sh4���ؤ抓�/�K�Y�Șueab)̤�Z��A6�,u�2bm��Z�����i�r��`w[��^�]�xF�"��P8��ʴ�Ջ'l�] �x�*4j�5�9jνTkF�f뭸���0 -7�fC���&c�f9xn�'��/P��ֶ��N�AX%�4��Hh��3��C��an�M32�Rgb֓�ˢv���cU��X���U���U)��dS7d-���5=ܻ�w��X\�ًbN��*Y{ӱ�֝i4Ӭ�����1�5�`�L�g��kmq���m����)��ۧtݽz�'�Q_J��~
Lh�[�BT�qd��Y�`�-'w�[ژ��VW�jQ@F�Xt��[ݒ�)I7=�r�Ԧr	WJX���h@S�Zȏ@̚�{�e�vܢ�ܱM[vkr[�X7CM"N�B�8��&��r(������޵�k��9�X�7��.:"��Y���p6&�JM���.�ҵ{qTc%����]-x�A��v�c`�F^�{��J���t>�3�-�귂�0�����-ik���.��P[b����pD��u�e,��
��I+9j]��j���mȖLHc7��˷!t�u�W�{y�mU���[�*±]�Q�N���<����b���L�����ө��)��Y{�.juɹ�7Q����f�6m�Y-X Ti���ӢG�H�s$64��(�q�.�"�����wh-�n�V뫖�9�Me�c~Z�-m�5���0�7��,�7c^Q�UŤ�m�a�I=��Y$�ۥ\X$m*�z���.��7�+!���ӊ˫I1b�qJ(�{5Ʒ���k���TH��5���$�����׮��\�Ti(,�"���L�Џ�T��ә�w�F�Q��E��V'��]�6�"�2���y�V�P��D��Yn��Ӆ����f�d9�̵��a��B$:����kHZ{�-���oO�-%�x�h0U(��$G7F�bh����"3&�
��<�wSkI�-��j���!.M�P㼩���5x7�S�������[�$�nZ��R��%��F�#���殕4��2��l�M��wm^��yj������r2���V�U#z�h�9l�*	N�Nܭ�\J���=g�Y�P�5���d�D૷�:��"ح��ӧ�kdŬF�4�D���P,w.�=d�屍�ՉG �v4�R��8��>h��*��"����4�a�"�[�a���I���M7����K*�%��h:�I��`���h&b���#[l��iY�[������:{�噛[Kh��� Tm\�6���%���6���&Ve e�H-�W B��sm@�L���h*������E֚zCu#�DA�V�T�C0�Xl�
��Gv�6��U���Y��q5�ӱ�7H�xu|\۱.���j���"��d�afk�n��m�����n�i��Ou^<t�)�A�&яUG�r��v�eU�(K�SN�?�h�kl�j��Sst�c�h	ԛmP�LYF�됱�m��0
P����l�4��\�e暒�Y[�*)(��Y���4�����e5�X׸�^�%��@�FcSiV�$^X�r� B�����܌�X�i@C��S:�*on�ZK�Ui�m��ef��(:4W�QP��d�#k#Vӻ��G^C*\�gR�IܕuSF)	x!0ݸ�6���*���d��!0r��!Ef����Ѝ�e�5����#�B�*8��"�4��vV�߮�:5,��F�R'F��०�^X���,�x �t,��rb+T��	M;%�w)��v���q�č�.͂�&��mee�K^<�P=YJ�4����ϐ�^������̪�uR��C�m�zGh�qIy07u�Z��*�"�K'm�1W3l_!W�>�N�oR6)�:��~�F�P��Jjn^�v!��'��S�����;�yVZ�_���,�V�� ���C+eɥ��3!ǂ�1���<���Z��v4E��u�]��&oN���hQR�nr�U-��d*@�0EԴ4{�q���.7iO$�f�qf��HAL�y���Y���	�Q�Vh�by���Wr�ؔ��NB20F8�&b���6��<׋0T�H�y�뙰����o6�S�67J��u6�Bm9{��Vֵ�����Y2�f�6f��h�tԦrF�Z�5e7x�ho^&iu6mc��/4wa�C����`1�kו�)ج֜ySh�͌�b�ԍ�^�6*٭,ăy.�Љe�̅�&�;��S$UջP�Y{>�*nUe3PѸ��u�.��x��tcr���bU���)�-�A'Sv���"$�*�rIM�Q���fVm�j��!�H�܁k[���-����QX+�(U%��2�*�0�vi�(��Wm|3b ��J�4��D�2�[���w	,h�$J�u	�a�϶����lBZ�)N�����Z�-�T.�t-ږ�Kۤ,:CB*���u��������i�BdW�g�a�V�I��Ɛ"G.�#�h��z��ս88hm�夛�;Qe���mJ�.��Z������Ss[D�1XN&T��V�����ۤem4�VUجU(Z6Xu��X��Mn,�0��"�q��ǭ�ᨲݛO��ee)��{��ҝŦ}q��kE8��Dlz�R�B��]L��91:Oۊ��!]h�VM�����y��D��&q��÷L1Xnka��cF����ݥ��k2�*dj��Ӳ��U�;,bR�B�9�XX�XT4� x�X��q
Gb`3]����ܡ`�:2^2��h�u�B��S�֛�6�CR٢���
�i��[-�b��d�����&ߙ���B&l�x�B[�7uYN�)�oNL���'j"�{x��o�-�r�2*�r��!˦C���;0�6��t1L�;�w�f�6E���Z���k4k;b7�QT+�g/4�l�^�Q]�KC]��f��7���ߦ��0��<NƗ@�ƩP#jS�7f��k���C �H��R�kj����XY��m`�t��j(�1^L�e%.��V�*�^<آ1Yn�w�r<߬V�c�F�4+mi���eV���6�&���C6ژ��Y���˖�kbǫe�VEe�(,�h�i6����w�m=i�xa�(m�Z�aך�Ϡq��2�`ֲ������+q������RfB[ͥ*R
��$��v=�{��\I�7@H�]k��PfXs�74��"�-!(�M(���e�XB:���.9�4�EvTpm�0=ĩڦ���87�K1")Kr���X1!J�t�^�)��q�2R ��*w��ͧ��ڃ�#Ӏ:u�n҅�E��K&(l�-�������9�(�УO,�ԋ�/N���K��ŹQ�ᴲ�@F]K�.m*�Yو$00,Қ�n�w{��J;��fJM���.Ѹ%O�ï1�]�"u��2o�w��oY1]ۡQ�S��P&���]���a��M�+�A��/v,�@A�o^�f�Tei��ʽqE�5j��t�[�/h��XkpB��+j�����Zn�F�6fˠ�����l���ige�7SZ��5K��jIz�R���ݫP$�7Y��m�f�{�iZZl����h
_Xi�F�wt.�H�{��[�E����Rnml�l�R�>̒n�)���@t�H͓pG����tӗ6�D��X��d�0o2��H���h�d]��I����2:����N�)%��/mL���4�i�C����qѢ�HG.m�W���N�롻BmR�F�!m&.��usq���*�ԑ�U���iۛ�,���vїg �K�n� ����Ǌ}�Q���Y�J�̈́��m�!b�Ц��?Gj�,hY@2t0*�U�B��{Up
��ߙ�����6
 T�h�su�����<����Q9y���v��zf<���bx6��hz����ރ�������x!r��ɶnY��dw�l�XO�m�K��u)��m'�Uj
yr��h*;=YbPMUj���fB��&�4 fސ���u6+�Ն ���պ�Q�̦�+3R��
��A���:[��Y����.�"�JY7Jњ^�	���goij�.m��wD�ph�i��6��sl�Vj���M�Y�����A�cZW�V��u�WS+N�n��S��Ɋ�М�n]�U(V�K�xw��!�5t�cںa ��S�L�
 J��͈�&�H�0K8��[du�!�N��7��%'v�Z��/Q����1FC#T,�n�;�eXxjZN��`��f���1Qe�MP�d���f�L��&�/"*=Q�+7f"�Z�Wt�=n4�m����jgj�z��o���$�B�Q�2s"�-s"�������o5)�X��q���v��M&���
���<hЭ:���)|2Q�S�K�$51y��Ɇ�

V�B���Z�i�w�U����.�L���LV�fXi0ö����C[�xMi�6��AS\˚ޙ$oR	F�h�+nA�5W.=ѱ��v�է�Ӯ�v��r�a����Չ��ܣ(�ak�e��Wo�\Ԅ�O���}�n7X#��h���f�i��WX�5�����oXV�eQٸ郴Q�	c��Rp��R失��\ȪK���h+e��j����k2n�%�f�E�YG��&�70	���{���9'N�8���͵֣�)��ZyX�N���4�{U�=�ǡQ�����k�����0i�]��5&����ɮ�U��Hű7k�P�������Hr��@�ݡKDKx.�޹cq����R�;/![�Z�K��*sɜ�F��A�yc���,�+�k����	���'K�֜wwց\�(73��+�e�����=�c�r�=,��<�2�H�m�]�k�x��M0�H:��{��ۈ%�W7{:;L���*��jn�� y\���f�=2�����2-�n�x�:�l!"��RT�ҏ�!���R����l[���[��=Rt�a;�x�+��A~�1�Z6;����3#����k8��V2qO���L���:�����d��w;�`��4��n[.��'c�K��j2MFv�AZ�-lS�C\1��L�3�����ÝF�-N�_����A_su��X_JN�ض�XA��=�X�c��˾ܽ$'�WZ�Į��q�d�.>����s�R4�+���*G�3Rn]�S��)t����{�ݚj{��87rV�ؠ��Yu�nc��� ��N�3w�-8���I�ŭh�3m�P�d�Ka���M �����=�-��c=��4�D|�	՗ö!�/��� ���ԛ}BO���:ߍ�ʞ�ʻP��N4TR��L��j����+$�=uۀ���yHV���D��R���A��K\�B�p)�t{��|KzqD�PsD��K�3���'^��C[6v���l�/�����==y���-\��*���5-�A�Nm[�eG�Z��kH�yv�b��q��*��tN����WU5�O�Yg9�n:���u7;(^e��T��Ӑ��Ks*�6ye�e�'n�T렲?��4���A|Ĭ��Yy̦�mK�e��oAA۽N����8��k�Uk��-���=��H���N�׷�G ����O��WCd�	��RfD�KoUu�7�7Y���$�,<9��G�T1d 3���Z�/�0�3��F4�Yi�$伬�Ծ!y��D0t<�V[9w1m2鋥v�8
�W"�Ř�Q㻄�S��k�|�� ��A\�
��:+"����K��2N�q�ʟ5{�z��u-r�$�-}ٍ:��y�A�hwd��2����$⢹}.�^Q�s��,G!�󝕫�+wo�D6I2Zz5W,�\���)[B�Nѯi�=�FH�v�;}i�J�]�4��N�V;ޙ
�j)���#ӏ�a�;e�7Qn]=t7��9[�sI�bp�EK o�}u���D
-�����!�7&]���]K7��_p r��Kd�<�f�J�3��Aۤ�#=,[F�^�9�
�X�8/?f!�i�o(��r��!��Y��)�N��R�yZ|�tt�\ZT������a0�3i�s��Uw�e����� �N���ͩ]��D��t����5�7���|�f�gWkh�f��]������<Lܑ�
w���Rx�;u�gN���;�E'"s,�(r��N���d��t���gl�UI�$"f�ʲ9�=���ηG���Ad̛ۏ>e�V33mT����ޘY�v���
���'�8�\��l� Z�۽\C��x�d->T_m���aci�-��j��s,nыQ���j��P��p��_�[joV�g��վ�ד����\�&���֨vu�QV>-%Ӵ��(hy�s��d��e�tJ����FjB�;+>���խ�x4ueGj����BtʡĨҼ;O�W/Q�PR9,�V�����BZ3�s:�T� �)��p�Kt�����/6/��ù)�-*٥V�F�c�sB#v����萚�dk�N\Y�9u�Շrk�|o��=�Z��͇O�O��HRǮ�sM��9&;��L�лi��u�w(cf�*�w�GX�H����i�f�ܙݦ��V�w��FGٙ6��f���N\��m�SWY[An;���Г�=J_ ;�A)�BD�H��uPM��e8��&+�a�kj�I�;�[-��� �Oh69q~˗b�,O��Fvu�A��}��mo�^󬴘O��#�vw�` ��[�a䄮�bݎ���`��oX�uݩ�7B�{)P��Q3u�{��J8u��ֹ3�*��z����sG�{D;Jܽ`vSޏ�)���✺*��:�Իeb�e����׃q����I�zi���fJ uC��k��GR�p>��|.�c�Tpp�L��)�@+<�h�R껴��K�)����PB���GS�o]��C&��h6��UN�7��hԝI��/V!V��
)���ԔOj�N�j��/4��Ƹ��:��2;�\��a<6��ϯ*t&�d����F����V�Q�����r�6۫����j��M�i�=�m2F��nX�Y-�Y)�|;�N�I�݉CwB�m=�M�H1���͑�j�='�lҴ��!����_tJ��f��R61f�9�\����Bs����B,��u��nJ�2ri�|�=�I��x�a��s�B����p�^�����\CLር��}�9m"m؃nVkׄ��Y�V5�5Е$T�2�;�)�����2���tvV�V7[��͏q���a��0N���b;�����W��*_W1s�V�Ȇ��;h\nwAa[�#�$�j�4c*�7>�����Q�������V6N�S,I2��𕢕#���wf�`+ c�����]qs�#�x����6:GoEǝ[��ݢ��ĩ�3��ڕmǂ�Tpݚmǔ�G��u���:H�B�k������0F"�[�6 �z^B�Ԋͽ�����Wj���v1h�zuS|�:�>��r��|��f�PI�����b�m���]���\��:���J���N�:�b�)wf,xj�"�c�9[r]�)�P�I��9]5�PU�	�ܵ��+u�
�9I�ץ��������B:��\&}��_\1-[R�@�'v�
�`U펺��>�v���U�QZ�]��L�8�.3r"��=����d�͈}R{��u��n
�@b�w���'ٵ;�YewJY����+�'G(� �GC�g��q_Uq�1�oZq��ob�*�6G*���".�uIfR;��i4�hd�h�c�(�\�m=��V��W�lV͖(�ӠsHӉ��^��H2���DJ 
��r�D]�����2 �P����a�ݤ^r���ΜY4w`n:
��kL���B�̧��niD%l)���0�̽�3��`��B��2��ۮkx���u��A�U��L{�24r�0�W,�.�ʊ*W���9łt����}�s����R�e�����\�Ƶ.e�5^$ݷ��Q�o�t���߱��(n�����i�M���X�W*���R�׼dԕ���,A���a���B.2����|�*�vm&�����v6��t&���t��7�,Dt�7T����]�����a*N�{Z2���W�Ε �w��k~f�e�r���w8�l*��֯esǖ���R�Z���c��*�IU��*��mӓ�]����ne�U�$��W�>�� -Thq�p��A�H��5#�|���FmyjI�����p��[�y�_'�17F�S.�1�r��ܐB&Nj�[�zn(0-�S���;(�w����8�k���/�:`PuHYtv��f�5�"��2���Xz�Tx�&� �r�GQ�T�v�@FQ�k����ͫ�a�YW����fNap��~�X��x����0;!ץ���O�P�ym�M����ZF�����$��P�B��������.x��^�}umj�f���ejC.��C5d��4�������dC5*��Y�&�{���Id���y�SJ��P��ܝ
���+�w���*Ȯ�6l��t�d���PST��ғ�On�w]A���e�ݠ�VgK��i��Lj˩��gt��c���tX�\ܝ��Y2XnB3�MnZ����k�ٔ�̼�I׬�u_���3"�\���_��hݙel�t]�� Y8�5�����#�#��� N;����˺wHi�Ien'4�;[yk5l�S���\�F���<�A��(C5�qzq���o��:N�j-����*`2�A���k^B�ӶU�o�p��]Y9���Dt�5d�f��5��|�̀�1�v���,Y��E��;駁6R��Mn��׏�N{uz���ѩ��lZ�Z�`���ň�[4�U��46���eг�k�WX� ��[����{Hk��LQ>OVd8�U�)b�o����{[��o^��N��;���4k]M��F؉6��mrn��8z�nb��Z%a��N��Z%�ո+5�Z��;	|�Ҿ�f\9ژE�dC����̝�]ՠ�˫�m������&9��w{Ne�2��<#�ٳ!z��5����ǉ_k�8�׊�gh]��ͦt�]8�qm�u�oj����͚:�59+������u%��W�+t)��w݌�J��Je_W�S���ݧ��i�0*��u��D���� �O2V�-����B�W6��tqw	���9��Y0E�[t;��^��h�{�,�6R!Ǵ7E��[neZ���T������{n��e�wF�������.���&�c?XW�6Hn�����=pm+�XQ}a)f��%ChRõoL"��+����E6��Ю刨���P�}YuԎP�Թ��e��U�Z*��l_?�u��;��*�ͥ�e�ހ��`�����Q$�1N�M��M��K�j������/v@]��e=�h�
��2��Z�1��Q*-\ֺ�r�vޥ�^�c��fˏn��)��,R���&CKT�5fmZ���ۮu�X��y.�S�"8�V)�� m^�[��K��7���'x/��˸+)�z�Z��0fQC]��w��zn���ysdx�ʢ��'�k��S^XøK�����+8�2X�:��b��S����o�=�_d*�Jt-��|���g����]�]R-,��*��,��9٢_V��ڕ����K�*J��엓�f�q�Yz�E[��Zi���S>���MM�z�Ɛ�xyU��j+v�R���*�6���9a�<��)P8c���\���&�1z�[�F�0D�܇;�/e(����R�Z{��
��E���{xW���P=��J`��»�.��4	F@�[J��ʾ�2�f�goQe�����YU�����i��[�e���7R�46<��ǰS��m�@�v��ϥvЋ���&���K�F�a�S�F<�qK����*����*����.a�of^!����[���#+��F��.��D[���=�����ejZ�ۊ@��\��k@+M� �,дvJ��ŚJ��u��Eה͓ݭ5{pN��"B�����b���UcX媈�rr�k��([�(*��h`}��CM�A��o��vq긢��&���8�Y�к��ۜ�ݘ�9vd�Y�t69��NX��躚�D��8��R�K%oJ�]���J��Pޑ�SU���;I�J=n�,Pd���0��c���f�b�N[r�d}
ս�:B�*�l������>U�V�=��͐Q5�t�^	��Ytۅ���;n�Dn�L,�x��a]�*�Չo8N"����T�BGR���q�6���m3�]��lՕ���N�V�*� �]�;ǻ;+�L���e�!pO�b7�&F����v���1�����j��FI��dW�Ɨ��"7�6:zۡ.kq�B��uk0���}����[�����2݋�z�hV�]Q�S*���m5a��6���u��9Hd�ج���C�i�Pju�ѐ�V9m8��B�ے�B)�
`=����9v]J
���T��X�s6{f{�i2�������)�$w�p}dUm% ���ě(+a�L�T��FI�.��I��`���Ż�/j�oNM��g��d���Sg:��p�a�4�U��@�[0�%v$j�n�]3��S3Uik�����k�ٚG$$���Q��b�����̐0�F��-���c�]_����((5�;{^Ln�4#ʓn9�1Y%>齭�WFg=��mV�G���@bU̠V�ג����4��&�ϻE]�/�β���Y�o���� �"{h��q6���q�z��D� �Xp4��݂�ᯖ�5��R�J�4�̢y&�\��|K蹨�t��wR���>�/^����)�녕�sm^�dWYzm��][V�rXQd�%�#�/8,�*m��m��u.���Z�@j7��4Z��4fk��<U��!�F)}ikX����z�?�u_]M��;/.�;їPca�t�S]�r�zV�XG�����RJ\gI�D7b[��N�N�uJ�FHs��Vf��yh�����mwj���}�F��Q�d����=Ϋ$ͦ�QgX;��UCr׆}nA�X��jZW@�;o�����p��K.AFk��i�m�@�4�$�6��{�/��shs�e�k��b��J���*�#�"��`۾)wo�0m��u!�tv��t��;��]��B@�i�G3�Op_�����,bb����r�i����1�GdT���u�U��ՋA^�fY�܂�{&�]CQ�"�Y�����IJ����a���NrSL�PG����ʃkZ77`���K�S�]M�o��P?�H1ǂ��J���gc��l!eN�Ëy�i�|�w�@�M�ل��)�:q*�#�,�&jQ��i^3$8�>�M�A��*\r���y�`���MD>�,�p��d<3R�{wл�=]�\�2_P���p��i!]�LW'qx�s�4>��l`��V��n��P>���ӮkX苀gT��Œ����:�̮�.u� ��=щ�XΤԭpoIo��i���*��H
ܕ>�9�K����]6�V�fM�9no92'I*���N������������1���ￎ�����O��VE2��'G8f~�o�uG��HT�³�ɶ���k�R�� �"'Pgh��]N��U-5�bug{FԆ���4
�m)�]�#��u�1*�^ծ���+��|��S�����җkY0��8讬[i,=T������,�e&�\��:����=��mđ��ˬ�-���4�T��K�8��t񒲲,X;ˎ�ܳy:u18��:�y)*�~2v���{�A��4 ��kh����2�D��"����J��wMn.:�}�]t�r��ݛ����L��1�� ޟ�:+�i��5t5�̷��3w
U�y�ܧ���GJ��5Aq��c�jz�e�2�$S-Qpʜ�єR:�l�����PK�!�Ct������\��ۺ�����H��W0c�u%���9$��0��D�+��Nú������ll�9����5N���_V�ƋddS#G&Y�֭�^�u��s�K�ٳ`4� ��ճ�{�9������U�����A� �O.�f1q���Rg
݄��%�S�̸�x-*Z��B�O����:U��fP���p`��R�X}4$��ց����aƻjˎ�M,:5�����!bRpIo�o��"ѦH�����-o6���]����^p�՗�j��Zz�
��CԈV�"�ha�Wt/��:㒊b�} uڊ�v9��ƁR#��ڴE�ח˵ �Tw��+�Q\��tƏ]�ԉ�\��ĆqJ��2����j�mt�kᶌ3��������hYJ�i�j���VX��a���fM�ʷ�:�a�oN�-I6G�1eբ�.�\����r�T�K�pnu�N_n�ي�
x���Ȁ�����KѾ�tj]t�ݩ`�w	׊��/�eNȁBl�hCKj���k�m���G���nm���u̻��c� �*�Z�GE�|{Vʵ$E-��F	nj=�Q�A�y�D��̺��>�r5�����6����^��{�l��Z���*��� v]���Ջ�:����R���9�V��m΀Ic�VՍ=p��n�\�c�˳�!��
5X�_-�*kx0����]���{PX�c�R��P��YU���\W�-�i��Jw�*a�D��n+�v�X�s&�G-V �㦠<�u˧M����q�թ\��N�%Q�Ek�X(��l7n���ƺ��2<9|�S��j�B|�w[��vel;�o.���{�P�ԑ��S�
-�I� 3���)��ʘ�\)�����>AD�EDn��@AgA�%�Jdy��66�@^Cج�$�W�-��S>�g9zt7��K��[T\�	���7\��[[A�G�23H�&�go��6;�:e�j
|���u�6(LkqX���۪ b��kr���V��V��6Mӷ��o$K{}��3EoQ��/3��e��a�z�����#)wKзaN۲���d6�H�oh9l�����@�ۻ��U�1�l�+�����
�Fi]��ӕu׺B,��w��r{�&Q^1���I)%
,v�ԧe�ڛ�Ҧ��(YV���B3Y�jhԏR�Ee� x�@sνE��*Z�pEW)\]�f�{4h2�EX��u�B��F���w9=���V� U����N/_�M����\	������@V���Y�v���1��t9�c��f�&M�Q���5��GU��Q���k4M;�	?�S0�foL����:[ݬ�{�jIu��T��ķ)�W�C�fƟT�ǘ'Z��=D=�up����t�r��<AQ��Y1�4JxM[��R��,��2d�d��ݴ�VKA�nsڲ9�r��*�h���M�4 ��\�}Nv�����Ĭ�h(܀�ڽ2�-���ӹ�*B3\Q7�*I"k�X�E�Jp��21{���[�H�镂�|D*N�6��0���o�j�.K�V1����o���ĺu�3>�g�m��e*��IP�ڵ��n�ld��KlǤ���(*F���'�mm��"6���<�0U��j��h�[s�x�k�']�t����3-��e$k2�<�<��R����Ոt�-Q��/k�O��d�-��h�u��U<�e�S��Q��,��ۚ֙�ˣ �y:�b�����@��N6���+��p��ں9�W
�2�lH�Mj�S��a�[��
��s��;.�4g�^:��:`�7���D����r]{\�O�)@ۺk���-���UǮ�-Y��eD[�Nv�֝Tn�K�z�[J��Rk�����w��8q��t���K����b�r��n�HtL����-�MЅ�	�ǀ<5<}q[��QX���Z޽T/��I˘붺*��w��ҒjB�}y�\ԁF��₁^%N�Go��'mwd]q��g��Go%�X�]
�kyP�.rJ�F�Kr�j��.i�+_]��VmBVV���O�������>t6k��de���ؠdts���y���&k���,9}�,bf��o��Z�\�n3R�ԯ�1����%�Gx7�%e����ݪ��'/.�t�ow �mp#6�T�&ʄ���m�� .[�\���݇������;]@;R����-P���0�I,�j���VgI�?�����Y�m���h���A��m�h����ؙ��,I&��9>hQ��/E�qS�������-�gM@�[+hD�>�!�=��]l:r�Q �iGf�1^��-��J+:.����Z�P]:*͔�w�1TB�W
�&F���ź�,s�픮��6P{.�R�}N�-6�*�q^&Q�]��n>����Gz*�d�07`d�*�Ǆ���8���g�T-��5˭�2ľ�]����줺K�ɥ:��V��tZ;C^�%�n����L֊��S�|pI��ughM�����)A�[D��Z��P3��9nj�ֱ˔jK�,w�
li�՘�pdx� ��>�]C�C�V3�~����걈3��j�jJ�۶m��6��ݰ�BT�ՠXc�ڂ�"�E�V{�)�N�JĒ�����ݴ����f�K�j�0��)}�t*5����;�&[�LѰ��wo�ʃ(�A�3�jgKI=g�i��X�0k.��;��ߊ�Z���R��.H]d/�lm��'��:�֖�F��Ytw��yh�G.��i*��8'���G���1E݆'G�g���)�y�*V��K���m�j��u��C*�hrt��z��;���lp�R���L�7����,ߢQ����(吖S�Y�M��v�]x�9gj�4�X���H��M17cu!�'R�t�r|sfX��nAB?���oQ&�sųs+���iA2<ױۻ��m�y��9�����1¦�s(].��\��9b#�Y����F��u��D�/n����r$o!����i-행��(��O�v ӣ@ˑ��"6��k� �]��C��#u�v��0�RW-�c%vJU{B{حQ�Q]���|*&�{[G��.6-l���1z�{`�]�v����/��K�)X�Jl���b���+�j&
W\�3���7 �
����1Q	)ө�d�X��Ɂ�\Ӝ�@���gnJ.5*nņ0�pκhlGA;k���v�:���=�%����|j���<ʺ�F�l��3�����]}3k&T�(u%�PDnҖ�9Nd���SMY�kn��n�ک�P�ph���!�ፊ�����k�Ŏ��pmmEK/h�K:2�֣0Ǌ&�9���U�S5�ŕ�wp�d�G+g7s�+:Gg��Z����TG�J�ZhF;(��vR
��hgf�/E��;���/��EKz��,�;.Qj�7���͞�M.�{�⩶C.h�}D��HY�D��&��)�����DZ�Y|+"�T��V �ӎf�/���Y��8�j92��ְR��t(��U�ur
�.Z�6�r�R�m�b�%jA����wܬ� ���\]�y�gv;�R`(���մ�i�YҀ����|oP�{�_(j��R�u�_-α5�ju��.��v�5�+hf�C^<L��&����q����{f��\ؖ�g�y#��K�{�@�lr�녨�+suJ��<�",˦�����UY(L�qQҝ��A�-�d�����@uJ��fک�wR0����]��`|��� V ��p�u/�����b�W��@�U�ذ�'��'d|f�C�������`�n�o$	�TRG���O�=���)wHj�RY�;�;\)�k�ݢ.\�\�@�N�gj��5+
�K�f���_Wu�ؑj���m��^mû.���jƺg�8C�wG�9����(u�&˽�F#U�c��&��Y.���ޤ���;3vZ�Jl���;G�D�rX�b���ay+E�TDrw!�.��b郳�(U�ݽ�|��[��8�!]c���vQ�8�vK�m�wr5�-�Yk8.jKX�agY�n�����ͨawtS�����f��y�*��S�f�5��:n�W(xf��M���� �C�>H�}�J�̗����Ce��ضЋx�.P��meǔ$�Y��s.�+�v�һ+z�SO�%���&}!�����t��}q�I�9�t-:I��}ݗ|���i4��8B`]of�-uN��Iq<]��^���C��o�,8K�8�.��yl ӯhn$�ͮQ��%�๏�7���#Ǖ�ʖo�ά5��n-ҮLWZ����&}��V��Ȳ�/��� ��s��Su�':Y�jaCv�V�U��]uES�����o^�o���#�GyZ�ݍ�Ze�jK�̪=�U�e����j53�����e@�^B�喴���r�T&�Mf�P��62����d���m/�2{���� �(�6'+���C2 C��-����ʾN�����ٹ4,Ư������:a�܏b�M�z�_*؊d��R�k��]O��#��*\�ôt%�34u���A��
珰�]nѼ��o�vJͬ�<	\g���tm#�YNB�<�ƒ�c�gE-g!�����.,�
�|�Cn�1t�+��v����S��"����8����=j>�+��v�U��+�G.�]���u�w��+jҸ	$�$6�s�ux��q�ﺞ��5��X:'�f��	�P�ra��f��9+Y�2��6�2u���]�#kv�8V�YL��DŲNm�岈T#I�5��)��Z47:_hZ^�������E]B�:V��5zʚO���:+;T�⾽�9̻(�<�M�GX��Z�O��Y��[�Q,��pQ'׽��g�ْ>�4ޫ�0�U�l�Q���j��)&����9]���ɫ��z;"LU;�\���J��.K*p=��X�����j
sk¶u�0ۮ�pw
y�7k�J��M�ƹ�]�{�VG����^(z:��5���z1إ���H����p؍Pu�m�O�{B���V�W�;eo�[r�!:+�����Z�s�T[��c=D���4��t�&�ػMx�s�/��m��DM�Qq��d7m,�=�2Ӗ�w`X@V(r��{����e�+���aR�r��b��i>wF��� t��[$!��ﻓ��sK+:��S'/�v����x�\�CA����MOr}"u/��ܦw��w%�̮�5�J�ԤW���� ���¥\�n�7���m �U�wGQi�_,�s��Pc �÷;#yg�b�5�u�I\��Nj��]�P�
h ^�������XZf4:.�#�aj7gju��w�(f�1�|����_E>���b޳���8��$
�E����Έ]ZB����-�N���(R
��I�9ѽ;��1-�md��qb��A�QfI@U�2V�6l'˜ڸ)(�;7[����*r�1��N�Q��gb�9EV�N�x���<��gEB�n���>O��wO>U�4�V��
l<HZ8 �nИq�� ��]gud�7GS���"���3�ojk�9x�\��ɝ}Y�/��o�KE��P;t���)'[�%������wR��Һ��p���r�7[���l���*aXM6v�4r;hgu�q�t�-m�gT+��4HB�אc�9΂��N\Gk熵-T�3��}E|F����j�X�ms5ˢ�eK�e�g���+[B�8��c�@h�8R����Ư�ՙ���'z5I�����/i��̏(��Z�N�Ch�U��9���p�d���	��b����6HJ���G���vթ����[\��Z���l"�Fl��K���4�W���O0�&����N�S�wE��.i�3�4�X[�/����r�}�o�L�-&�jf4�o+p䢂�j�:B# V9��ٗk�

p�5�̀�L�Ѯ�Z-�n��2�:0�a�cy,ʎ��
��%��q�)N�Sݹ�����J��M���V�-=������*��qC ��T[�.F���z���[����K�6��L���jsw}R�(�J-�[v�Nt*�<|��\2b4u�+�T�=VfV����Z�R�����tlm�z���Q������5н�.D���N��v�52�ɚ��K�C�����:�i�u��E\E����25W�h&��D���"�x��ѲS���S�ܯ�������\m*ݚ�مh����Y�=�譁5"��u�-\�0���l��Oj�p���n��Κ�p���n�}DjL�N����ff�f;b��Aj�_5W#��{�%Tv��%`בk���*��[�+r�Z}tpRY��wSOɹu*�y2�a�p'L(%�Ժ��F���ʃ;.��к-ȱ�hLA���h>�U�t��i�ݗE�Do;�I{��f�_���I�J�<������t-n�Mݸ�2��6:Pg���BXհ̄u˦�Q��ݻ�ie���s�5�څW���Q����^Ƴf��7ls�x{� ���\�Ny�������4嗐p�jgsUl)j޳g:[q>�du�����f���G{j�[E�l����ݎ%6��ޞ�c�X˹����P+3i��8�Pq���SD��'Qu�[%A���XbU��r���^�t�mJ��Nq7��i�e.�[��7y�N�kU�������k�:M����1wV-�r��u�ػ��ɨ�Vou����)\P��7i��Z���yw6��p�ƫ�WGV4�t9����z�12�r��c�������SŧF�1Wk�Hn��|�ސ�����*8��Ʃ���ƻ�س'�b
tR�9����c��y/��o�	t�R�xͪ�����>?Z����N��ka�O)0s�B��:�[����b\)�N�1t�Z�h7����R��
���J2�r���C5!��oc� q�{��k6�=#H�c)
�@e)\ѫ�I�}K�.�Z�n0�7n�v��T+N_8l���U�����:��	[�1���%�7R��w�6㮮v\ԛ{ػ��TL���&P�j��mF6�ZB��]�:�S�V/i�v+ �O+hM	q�c�o�F��ʽ����%GY��n5L1K�]���rT��0�:6uÔ_���_\��j�����'qS���Ob�;��o��^]ࢮ��� _8v-EB�Qh3!ۻtr�C�21j_b�@a_Ԣ�DG.
!ʈ�"��s�E�#�EQI$�D�� TDEAU¤R��M)�!r-D���"�D"8L����9G(�DDDTE�\9Lʱ#�)R�F���UQ\��*���EfTɑL�9��" ��h�vG*�M�UvEQkH�r�P�!$�̄��DAU�*��b!DAQʊ9�T�XY!E'H��DZ��:U(�ȮW4XAZ�A�8�d�Ed���I9�Yȕ�DQ\����
#�$�Zˇ*�HJ�*ˑ�d�$�G.Ur(��%B��+������s��\�EʙDP\�$�*r!!#�UE�HJ�NT\��i"��(:c#�����.T�1�UE\��%)QEEI".G*�(�����*"8F�]ReUAȨ� �	P�( ̈́U�T(P}�[�.���>�3ob����w3&Ĺ�F�)�=̝B�n#�*�d@Z�H�s��̡y�q;�viPZ��I�Og�d��9l꿽e�9@������	i�Z)}�����B�( �����$@��>n�R�3�)�gՇ�W����tqX�~r�{���P])lWv�Q��n�s}�R���7Z_˝ ��a��ks#y�ɕf�E߆�/�Vׄ+�'��{�ew�έy��^����fq8'LJȍ��4�����c* �p$	
��-���U�w�)����d�{L
�K!��t�"�X�l7V9ds�F4U�ӱ���on\�y�\�X=B�:&��ȥ p��Z:���ˤ�ȯ/�z^�g��U�)�k���}s��g	h�\A:!Qbx�)u�ڠ�؈gKqn��V��g���;<�6��/G��n��~�=�
$��$� �����B��Y�<?NL��x�λI�� ���p��Ա��,bh(��P$�`C�*me�?��V��F��+D[SW�������}Ie��!���p�Ù�^D`�J� ��=OA���w�v��7\����-�<�!XN�{x�!�r�a� ���[��m�k�4e���9�ƒ�C�k5永��"`N/O�y�$�ř]r\8%v��R��\ow���t�<�O�dŝ���Y�&+2m�3]v`fs��!��m��n�J��'s�a��&�<�}��ot�z��O��F���E�p�8��Q.�W�
��GAy�`kr�Z{��j��@����N�ϸ�_-uÆ:j����,nCu�M�w��(�?�[xy���g'��5R�o)��d@�B@�0[��"4;�0���	&���D��1���q0{7��Y��V�v��7�~����yp`��x� ��،�6�����Z�W�ύ�{V��V��I��L����i�8\3�v��6�~�>5�邶�U�S<V��2��i-S��}�s��ri��]���PEZ�ɓp۠9�3T6�~�'��P��ŇU=��oؕ6^v�����n�pXZj!��������k��5W��{���!VtP�퀵�ZNV��usU�"�n�S��E��Wv��/��FDjt8��`�:�C[嶈G���z���ĒAvJ�7�CX��aC�*�| y�
��`�J�1���:���s�b;%��mH_{9Ƅ�	��¾>��u��x�ڡu ���ex
��TǑ`����^�C����s'�ke��9��g��Qj�����]}�S�lw%.�k.�ȴ�L���*TporcSȇf���r2N�K�s��G��5r���(z��e�(��ޣ�ͮ�#�8E���q̕��QݗH�2���[��푸�冺��)rDG/��b���SܱuH�tBy�F�V����ꑪ�9G����7�y 5$zN�?9  ״�uN�c�|c6��Tܞ��$�'��0vSKھ�J���r����r�y��ڦ4;��n`2��7)�՞�����T,Q�1YeQ��%Y�b���ƛ���=l{2���5bV:c��:C��sj��)�g�!�����z�N����i�� $H�=0�mUD����(),X߾ki���8z�������먼�Tb�.��ʷ��2J�eR`ԡ�d�0�~3 ��,{QMӸ�����L�-Тj�@�K����K�SmAtX��2T� #>�&L@Ј�]YȘψo��V7��+���������3�,��-����>�d��,�`P<X�Vb<8���5�����ۄ�^�Dt�p6���&�nc�1p�q����d�w0D��0��<�&\l^ӎ�X�w���y��ct�{/M�:!�A|jLT$��6��k�j2+�t0�Q�*OfXxUm�����XQns�kx�x��΢�]t6*k�4��txC��8c���6�7�9y����ބ��Y����K�e9�tR���jw=�^_>/��}B}����[[cD�q[�OG+���o��;q�Z��v�JIۮ�� ��Q�w���~�B޸�f����3MeU���m߸��L!��_!��H�s4ܰ	�~�!�&�zf=���OL�w`���d�(u�z/0���rH�c��`p�x?������7��v��s��h��(\ܺݺC�M!R����=��ss���j
�n_x��=~U��ar��+�����|Kj�C��ߞ煿eD��8���Nu�Zn�x�Z�f7&�<����>w��dJ��@!�gz���#|�K����Y�;���h֯-��υ�}۴շ�L.�:ǽzU�	�DLw:�X;�2�����8����<lF�oo��gb�nX�m�����:.*g�B=�&����+��7)�ϩ��dg7y����)���ܵ,�SE�f �>\n �SOqت�!\B��c�2	�1��,eN�t��X�q��y��-�S�f��J��*�)'�3��O�
U<1�FS��yϱl`���"G��SXDGk�䍸N��d�R ޚ�(	�)���	��4Fj	9�������涟�==��
���*m�J�qZ���[]O��.��A,ef
�߯��=�9�oӭ�hi�t��l���Y[�.�9�yQL�k�t�4�n�t�8%w;�4E��u*�Nl��f��cZ�����qř׳+:^4dOX��Gypq�b���Y�6�gj�w^�yZ꽞�2ߝ�W\�"��DC� <�����ǧ��^:w�K��?\H�#��{�ò!S��`9��ȇ3!�19�m����\��٩A�ӭz/Aq�G���@����и��c#�	Z���C>rՖs�F2U�_D�v�$PM��~�3�#[};�v���"u��i����\bs��A�˕���=G�IS%�X�;V<����mOw[�H����U\�FX(l6}��˵�P�R�.�Ew<�15W'�8��*^�F��٪˕���� `k���c3CC�?�d�|�K8�u�9
�ߦ�����zV���6�9K{R"��o�ޜ�S���#m��Q�FL����M�p2~Ut�.��92�f{a�k���(�+��3�_��S\$ⵜ�Tĭ��-��l���5¼�+�u�cFZO�b|7�j��.Q9}����k!���Ҹ���X�o����p��;��p�	���8����n2��IP��=T)Cᙷ�e��W����|��*u�it+�xP�{�yͽ��mGb��kx�¤��ʶ�:g1�N�`}� ���/9�:���ƒ}�c��X,P���=c��Y3;n�J��`/v-z�8�pɍ[����l1!�\S��j��A�t�=�Tu�������R�>
脴�t�V�$+�	>�g",�)\����+��Z_ϐ�#c®�qn)�������w\t�RX7s��o�?�4�mZ��]#�,�^Ӕ+�8r,�!��r׉�(��-v�)��n1q-S���,�p��tv�e0T+��Q�X���eA͸���q[�|��e$Kz��Ϛ���4C�d�)�`���>% �|���ޜ�䫦�pf���T��n��X�a,u�W���~ʗP�+%�by�U��b�w��ˤw����i�,��s�f���k��_&sK��wp��O8
��޾Ѽ:z.p\������A�� h������%p���V�C�H��ml�<FlO�I�y�ٯ��K�J��x�$@f8@O|vH�[O���o~�ϣ�)8'V�\��C7��:[��j$���\
�i�8_�� �S!M���=?I[X*Jg(��Z������Y'yؾ��jF����j`��)�%� kbdc�� ��zh�<,{5�j�
��&o,��Y�:����� �sms��S��c�z+�)f�'P���=u�2��U�+G��oņd9��C,qb.�zsJ(m���1�a��ښŤy�9 ��=T�X�nW3ڱ��B�e�z��w�3r7+x�;H��{u�9�+���,@t�ܗ:�����6������\,�����̕��;q��t4͛� ry]| E�V��=j�Ⓛ0��
�S�����Ѱ�R��:c��;�b&�AYʆ=΅5x�W�������m���Һ��r� �(b�)s��T��l:I��ά�M���JҊ�
ퟞ;ˡ��9�²O�&�0TD���0������֗]��Z��1�Ŋ�+���1^�l>�ņ�,���B�7������W���kSqZ�����]�����>U̺؋w�
������nO
�I�%��Pu��WI+�p����Z�/���-�u�8�Cن�5��s��۔���ߘ�YP�F�d]�z�jo��t�H���gi����rLP�Z폭�t�d9���6�d)�g鸞�'{R��^�SbqY'A�.�$a�ڪ�w�؅�R��ki��N�h�Rn��6?iΊC�g��jp�>5�}F�P���Uo�gC�1�y�f���ZG�2��,��%?P��e��m����u�Z!�XL���zR3I���{��[we��Tר��Tff���]��'�{�M@;����+����WjpaKb ��.�Q��_x�t�6tn�q&�����辚E!�|D4yGŅ���]|�@Z׺�V�q^���;�tB��0\$��@������6
��"H�����kyW.�:qs��&��֪H�9��ȇ;X�6�X �ЦIB�����`<(��<�r���a��k�SϜ��(OW��7x�K�ɶ�8C�9�d���*!��H�sq0�K�\{��<o����r���b�s$T@Aa�Ұ�s��|jL$�=�s�����t0�i�,yV�ܕ�ίGq��I����L�f�m����S��\1V�p{�n��s4ܰ	BA��R�Osq��p{Ս���u�U�
C�^Y��Y/�/
L�
���;��X���(@�,]Ɛ�o�-��������7��U�E�/�j
�n_x�gm�o��k�L���%d��I��M�LC����ܥô޽1�!�K�����ei�;{�1�Q����4�/�*b%�녟J��@�,c=����|�x�b�ƋY'm]��s�}и�l����ߺG2_��E���l��ڈ��ṵw�t�y�[�k��o�v�e{��U�m��+v�s�,��������,7P��Pgn��O^�	m[�y	��[�oNa�م!�x+��a�]�_JZF��c�-�(r��b�ec�3�gT�Mh�ޥbC�֩��
r��ތ�8饪�-��£N���uR��S��XO^F�xv�p�*/Q��o����*B=c&�쁪���LE�ܦz\�|-e���V�EeW$B��Z�&���B �6A�AT�q���!_��tcT���c/T2>��um��]�yp$w?��Y��Q��	�~ӄ���7ae#T�f)\�'��Uyܫ%i\ے _iH�k�Y��v9�ϧ�I�,�5�I@B1H�ś�ݵ�V�He�K��"�էqVe��p�a�Ӑ���~�Zt�HKh�u��Y��Y	�Ë��q�=@�P�
�..���f9���s1�+��D�f����I��ql�����"#  �k��Ҙc. t����).�ȇ-Yg"�W�5�H�P D�q<z{�[ORAn�/}�r/��GY��`�(v�YU������a��������ۂ�u�WSn1�uڐ9�^��"0	LTD�T�; ��|}���r+�Լ��O��e�hsՄ@�.q[=�'.�S۫�.��e��Od��Q&¸�[�Ga�`y�]AY�Lbe8j���6�j��n���"�O��������ߺ8I'��z��V*-�W�_J(^��d(7�R޻����	w6=p�e�ɝĠ$�N)�&��k�Ydt;[6d6��4�u2n	�T���f��/f���fԞ]k+D���d`p�lB�i���N�rn0�b6۪�FL�0�p�r�_�'尭L(�uX��m�p��iM���ZN�͞f�_�T��	8�ek�b�}��^����R���눪��=��Ns-�fjS����NQ��d�}�H
�k!��]+���c=�7V9g;�k`s:�y���r綋����#@tTn�.�W��_Rv�R��P����A�;�8�I���Q#=���ۂ~V|�����(�% ~�d�_'��폆�"�b �;.,�P[����=8H��;�����x>�b߲=���$���tW?��״��]Cx�yfJI�pt����o�g��@5���N9D0���&b�Z�;%m�Y �10��J˸��ʋ��Ș�h3"�����V~rpv��;��o�CRY|r�c^uB�q���(� p�D6{s���U��Ir�c�_�O�S-�v��,p�ik���ԝ*�8��_K�B���p2't�鱟?sr��2���4�O=��eZ熎�M_�^�3���$}�}~[��g�����S2�o{C��i�e4j�*Y�\�P����i�o�S���X�����0a����YH��H�ꮒ�禴�۲��tګ��4k�I�ٶ�[Q)\8ֶ�[`��Րg�M��+�*c��eE>����*ٛWFu+�K/��2���k;�Ub��T�����<�u*n��Q�okVEۆ.T�F���(�#c�ǚ� �\�F]�P
��L�#�f0�Y*J��O^xw���gɿZk4��XT��t*�O.�Tw��\�Mắ��9��c���)�9�V8�Q����뛼sE����%�j���w���I�LEԼ���-��t�(+'� ��-d��ft��n��2B��D^V3�H�!�8��0f&���>��f�-˷��b�n�Yfn$7:E��bH�r�X����n�Z�f�8cWwą��w��f˺j���0Er���j̝�(4��=�R�W_,B�Z�J mT!���].<�vs�F�SX)�n�H���t.��;-Q|U̾��d��S������j�QP��ab��Ѹ��Iq�]���]�vu*9-�	�t
f����]���s�$��}���_�ݞׂt"��.�k���J��[��]ؗLub\��U���ܿ��f�)]-.M�nذ�CChDV1�\�8I���[�����m��Rtk����!�7J���өȼ�B���w;�fn����7��ym�U��٧KG�A%�gm-�{�9��n�!���b�s�]h��}\H��9��\4p_b��ކm*ȝ�<�R���P�NP��V`Nػ��.�qL��u��g=�q�&䦖�wVS�Cj
甡�)�]w�;���Ć<�I�[�5(o@���+�:)��.��"c��8�kݾ�`�绰⼲��7.Jp�.���\"�Wʌ}KsFL[O�j��/��2�K{ݦ,�y�������]ja������U���ui�W�N07d5
pcF������"@t�#� F�i��%
�®��9Z3��ӭm��b;L	��k;��nf=�@�e:O�8o��ʺ���Őm ��+d��3
�����.QSk��ҡ�� :r쒑}K	ہ��dj�R쩂:�Δ�7O��"���ܪۗ>z�1l`�E�ZMt���7�#�K�E��ѽ�'s�D��{2Kɪ�p�����&W
J�,�������;�%�ؗ*�SCW_-������u���`p�����q��wKw<�[+�MU�J���Ҩ��GL�l�U����l,�e�EY�m2)2�P���=��)�Wl���M<��Q��+K����#o�+-�הEN��xN�M�&m�m|��8[u�aN�(��c�v:�aṇY� �OR,��;�}4�%��Ϝ�vCJدi �F�1��y�� ;:�/��](�C�䲗VuIWO���3Ѣ"g��gV�Sc��f�kX9�x��X�:��:j�}}[y|�(����ʊ1S.D�YU��QEE�9ȹ�#-k9�"�W5*.T\5*(+�(�APp����5:HvAsD*$���Z�p�9Ȋ��TE���Td�\�3eQEQTE̐T��T\*����숪*�Es�҉R�����Er�"���+0�����.U�dp�D��Ar"�9s��)��Ȩ�B����*��dQU";(��(��r��D͜9r�
9tȢ"(�QL�(�9(��*�J�""*�("��EEL��*9Q\��.�*�`]ZEAT�Da$s�Ef��.2,�"N�p���L�TRaV�"�*��
��"9�e�D����Ed��I""��ȊL�E�֑�Q�̂��p�*�QF�".TUW"
.r"�QVATr"�Q��$��A�EʹG#��s�QE/����/�����3�"t�YO�\;�jC�rR���x�T�ڧ�1oɀ���8��k:�ɶ_E�#	�i��xv��E�>����ߛ������~N�w1��L*��X�(I�M�
�];��u I;:z9����n��;��O�k��0t�|��o?|�t� $�~��b��}���3T��g��|�+_z������������ۉ�O}����ڭ�u���}L.�'׎P?$�&��?�G�\�N����;OSv�M�;���?8�!۾%8#� �#�0ճN��U�����o#w�$>&�=?wї������S�~v�oS}���7�N�����M�	'u���c����t�z���p�6㴛���w{���J�\tp�a,�� �sȻ��ɘǫ���x��C븇�;N>���:w�?;����[���\|��:�q	���9ב�C�ǧn?}�ާn'~}~���7hH;��`�N���a����;�oz�ozXuL���Xjtٝ����ν>:w��o��ۯ-���p=�o��7�]����m;���w��η���]㏧�=�����&���u������6��eӸ�'������������<�`�|�X�f��^}����*N��=��:L>G�>Qһ봁������^;봝!�~�q8�}7ϼ�I�!>�|��}��㱯wL�ɵ���f�����=���a���8��Ň�H�s�E'���w����4�q�R��|x��Df�RV��_!V�#qާq?���s��aW~q�q���L>G����;q�<I�]�[����o�;]����
oP�e�}��i����D͏h�U�b+�~�g��߿}}ǉ�7���ywN�o�����ޱ��j�]���o��>!�k�o��t��8�!�����&x��q��z��0����&�����9�oP�q����q8��������g�5��tɻ˵�ε��a�` �^���y`�M��������:޻v��!>��;�~v�|��<C��n��v��q7�q�o�_o�V��o�������okz�$&���;x	�p�sjᯛ/��f&X���0fS �t���3zw��?tiIۣ��zݻ����7n�
OL<��ox�����x5�����R��i۳��x���n�;��o�q������'�c|O>��ߟ~���o.,��yA����W�^��eO46�k�quи�ҍk}��9�Q�j5��6�B٩���Z\���l̚��[���QS�1q��-+א��⾫�>�]u�њB^k�{2�q��g%���v;63�OЫ����V�e-6z��Q��ԥ��<1��G��um��:L/ø���׎]����o��:w��,��qt���z��q���ӼO\q<O��xz���|�����8��A&^'��Gc~�V�ζZ�����Yz�z���[ݧ�,]�ܭ��}C���o����=��=�m8���6�=�` ���$�7���<�(x��:<��m��e
lY�z�]���k����os{�L(��o�$=�7?�q'��ԜN:����ۉ���z���	����v�i���o�����@�/�wζ�Ӿ�N�{�7��m㸛���}�/p����X�}�>��#�u���N�o�����ާ���_��}C���PP�O����a��t�r��7hHN�w��ny[G;�Xx3{[�=����$I�5xt�M�؅yS/Y��]�{��ަ��x%�7��?;z���?���i�B;q9��q7����y�ӞF't�� �n>'H�����7���pz�p9yn�v���8�z����ߖK$�W�t�fOU��<�L%���� ����	�I@��7�0�����e�=v��޺�;w�k���y��ߐ�'ν�;��q;�:N������~�ݺN&����'�i7�z�۟�(�>5C�d+*�;K�l�5�x"�o���C�k����:w�z�!�_ߺ	8�]��<����]�p|}�I�!&�	>oz�}��N>����>��O��ݧ��n&��xt��?3.���I�Y��ԥ��E��(A�oS�}v�9�pv���;O�X����qݟ���I�w���?~��ަ�����t�L/~y����zC�|���?���s�����Oޞ��ذ�tݜ���K�-��B>�zX����n{a{C����}չ�o�q0�׽��W}v��'I�׎�>��'����:>&�!?��0�#����y���Ca�]YO�&�+"�z����s7Y�ަ��#��ǧ���0�>������ӵ�;�Ѻw��O�;���aw���ˮ�!��G��~���t��	2��\o��> x�����\ݻq7�N�&%������
*�ˍ̈�Ok��:����-^���Ӓ�B!���]�u*�yT
N�����Oى��[�6^�����I�q��8qS�+Z�N}i��ݹ����s�,�Q��ގ�)�ވB9n�k��ܲ�Ko��0���J�p��fM�NM�E���N$}T|��%�oy3� S��-�	�������t�!����|qۉ\!&�8�Cㅻ�N��q$����0���ݾ��z��N���$����w9��������xD��`�>u��q�uκĞ�]�����8v�����|?��ݡ�a���<��>;�i7x��S�ۧN�����7�.[}w�I�wo������������|J4,
�zs�]z�������C����q�'����vQC���:?!�0�m�9�ӿ>����W6�Ӿ�m���}C�©���{�w��@������� �G��*����>�>�;�wV�a�',��u�]{������@�:W�����v�9�1?;����?��>np�;�j����ﬦ@���z�7�`�v��~���z��� ��f�0����c���g�I���]�q��ܥ�ԭ��<Y���o O�� �/��vr�H$�;(�V�v�oP���N�{Nݝ[�:I�ǟ�|��v�'��?o�:��p�v����$�;q�]��xn�x������5��=�e�r35������Q!���aN��!�ݻ�x�v�Wo���)��ޡη8t�v�ĝ��:q�~;q�û�:C���m�q�n����_}�o�v���>O���k�IV���ު�e�X8oz[Žm���q�o�����7��x�Տ�u�1;��X����8����w�N8�㧉�]�S������;;�;�x���;�Nߝ;�������)��3�[�|���"����V
��O��ͺ���&��8r=v����X�X ���3�,q��KC [�98|O��S{��n'<�w�ӧj��'I���A�G�NS
����n4��
�L�M�O5x�b��pq��|뾌N�O�Ow�=��'������^��'�?!���p�]�i���{�s�I��?{�޶���N������v�n����r����$�c>�/��۞1�L>WYQך�x��{�?�S��Ӆ��2ɿ��qǎ%�w 3&��	���#�����ң|C�=N&�9�����C�� 8�>!8���z�i�����{������ K�h���:!��Α��.5w?j�!/���&���wB[���*{�_�IOq���s�B���U�iovP�:X3m%ȱ�R�\��S�'�Ҍ������%Gx��T�M�h�A�P���]����X���}6���Rl���^P�`�����܍�&o�����q����G����i|��HH���o]�'N��zv�8;z���n&�����~�J�S}w~y����B�1'�{�=M����q�X���L����L�i�Ӂ��-*���%z�®�>�y�|OP��z���wN����;�n��n:w�X�G_�|C���p�v���wNב�ۊ�����|ϱ�dxxt��7�}��c��UGsEu�Y:��<���a�QR��:}��R�r+�ӷ\({:�u�Wl'Y�yj�8|����X��健�3Cl�����������aK��W���\p��)==��{����g��*����9� ����f�T&�P�#GG��=6�t٬R)���g�q=Z2J�p�l�9ԫ�*aወI�k9ꘕ������p�L�ٍk*��Q�$2I���b\�\G�W�������t��U�G\7V9Bר�l�t��zR�f�vT:(�QU�
��
�Ô���b�l�O> �G<ڼ�}K��xv��p���Z����'������S>��l�d�#г�]Dy�N�m�>H@q���NX�R���o�!�NH�<����i���N"Jw}�ӕ�RY��s�#�4n����r��{�!W*�@<z�u�sa*p�ɇ&XEf��QÜ�Jr����̐YH!3�����������ޛ�`��b�ԧ�wqXP�:�h-�sPKWH1Y�gD5Ͷ��]�+Qp��.�@I"#�N�u�M!$�UV��9SÑD0���&b�c������������	1xu�Ca����f�:��'��:9��B��-V��5%�� h�6��\!9�e�`�����[�0�]۝�9&�&^0S��:�.��=X��K]�v��Y�~�uӝ��'�r�=�
�M����F@p! +�y��(E-uÆC���/KcD�jU-s;ѥ�ۉu�D����lظ~�hB��|,.��<6)jg*M�h���E+T�ߞ�V�󹩼��a��`d�n��x�&�4|j٠#9EYW{ጬT+D��nk^�m�{�~����j��۞�i�8_��?7v��6�~�>5����]�r�z���͡��r^�A�ˈ�>e��{Zj��R�2[r����� U���ίb|����w'u�B���Ǭ�?O�����«u�]>��7�25�̚�ܸm���e��TCU�srgw'�f
�A�v�u#^����b��c$�A%O�3�N���z�7bt�X�|�w�U�q�ҍCt��r�.�T���`���)���Β;������z���&*�-��w�������Z��/M�oK�{���"4۫��1ʚ���RX�fj�J����}�R<�km�δ�K�Xi��xb�v�#f��^���>�a6���J�/�n�?���i�9��m	u��9C�*�| O<������a�viV�j���/櫹�s23OF���3�4$��'1���{��_[���:km�^����[�	�`�(�(ր&t�
wPQ��+�օ:�X��zb�[Xt�8�����}f�����^>���38�1	����u��ʹ�[����e�|��r�tG�I�f4>쾗nH�Ԉ���C$�s�9�Bن�5���^nS+)���
�'��VS�\���+mjY� �t䂨΁b�z�\UK�9�ɊK]���>��`3��m�+y�ܘaq����y2��|�U�=P�Kύ�.�l��}uIR�}�����0u��\ˤ�y���mn�������85ݻ�����j*���=�b�|�5�f���~�s��93Ӹ��}��d�ޤ8���mE	�S%Mq #>`�R�ݴx��������o��==VEFi�
��'I�Έl�9��o���.�Q|�<5ڞ�mW�d̉�7�޵���A�
���N�9a���?h��ȏ?:wנ�$��t��s�[���a�Q�0k� 5ܺ�6�*���6qA�9�\2�֣�u��2�3�WE���PY��*�%t-fX�ip�"�'��ͧϩ N	�����#���*���6 ���zJӃ3����c+�ܖ�pa9�d���)��H�׾é���\���sV����n��y(�6bG@c��Gl�7��e�1I'fM�1�]�o\h��ηswd�Ҝ��:�7��6ݗ���a���+�ʗ��&�ꯐ�N�Eb������u��q�d�2�t�	����Tk�����롊�l)�yf8W�}��@2�MHf��N9}Z�rT%U!�'A�Hs���P���]�ɽ��څVSF���p+3��	���F�9��o��2q	S��k���-���B��X��3����M{��.��z�S��F�J6vb'����S\�%�g������^Тj�0޶b�՞P��C8��p[�3�GҐ�n�\���<�S��ȩ��ı^�:n-�=eMu�'��<
>����-���t��;cܡ:��-��pKJ�>\�۔�fi�J��g��O��k�٠"?w������R,BJ�s�u^����7������s82;j���7��z�����+*#&���i� �A*��8ʺ��5k�iQ�<��W�Vܿάs������eue������MntV�q�5�-Y�6��[��䕔4�n����dxTJg!�\n���}��C;K��h =���&�:�u���!��5�@��_<=
��(�Q�x�����¨�)�j�Kl�v,|���Yb�'�r���jK1���zm�T����v�����k�<2��� (
�Ľ;��ܩ(��C4��+j��=���1�q�":�x�FK�Fv�"��NTL�&�k;3x��@ḿ�;��_����0��-���]6a� ��G!��
�u��7¯GM���m�n�N.[����C�8\:�#��@:y�Дa��,$x}{	u��C������Ã�nw�W=}����s��'j�n�&���<"`�=g0�j��=�Q�"��}�'�Y��,�ɥOw��I��UĬfX�c�uJ�.FX(t6}��.��^���@z�����ɾ���W���U{ܝ�0�7,/�~�t��݆����Wr�w���C޾iM�"�,^l�ژI:�.5:ɼ0�m7T+��roExV���i���Ƅ��3u;}��?:�Hd���߳g�Ω�R�xb�p�O7�*:�{,���\�U� :5�ƭӄ�蚲�&D�H�8N��:7�j_+ ���#�C��1����}�t=��Λ4T�v��]�I��r�|�a���]�<��a��
�\����U5t
�	��=�Ƅ�8���E�[��:*��	B�'����}UU-�l)��ڼQ�������t��&���'������Z�c%�D$����WRgQ�:��s���Ҋ�7|�_�\6W�n�]
�
���
���9� o��T��[p�j���z{�b�s�穎�����O�ˮQ�d��~Bꌺ��pϖ�ݔ� ��|<��׎'[]�
���_N�/b�1
��׾���j�7xI�F��w�v�������o:2w/���-.d�P����4C���0Z�7�%m�G	�GA'N+��,;���ֶ\�]��ԭ�g�p3�6�d}?��<(M}ڭ��jK,Fb���B���-Rɞ=�,il6�d�J�F 8x������[m�]*U�Ҕ��:\W�ԝ+R9F��_*tX���,}���
�AYⶈ��z�@	�y쬎2�T-u�-������W@=���-��:8��:����/m-(!�顥}P������F������fu��>�-��D����+C�3�1��_6�@�x�&��� �7	o���M ��ԯE/G��۽�u����,�[d�u���mr�v-fR��wS�<��Y[�@���%f�Ԝ�^k�;/�ZQ-Jx[B�����{ qͼݼlE��S]�̣ș�^Z�0�$g�A$�4�ntƬM�0�#v�4*Ve;G����<�Wsyv:�Y
�K���Gѹ/T�]�ԌÞ�_p{�c7�5��^C5pB,�)M���4tgtze����>�s;y�ͯ�Ū�W�JGh�wJ�i:���"��ɓm��<]G���|��M�䞜���5Mŕ.�"�p�F��������i�Y�'v"��̚n\��m���z�rD�	�ܨi������L<8R/Ɯ:=�c��^�N����3�9��7��KE`��:�`��������'@�^G(1��Y^X{��e7βk�����0��-*|�3�����/�}�q�'^��7]
�������5�����z����x���&ؘ���u���P��(E��I����\��5��ʻ�v7ӠT��%��{"�&me���5^G۠� �nc��u�
�����Ud�
+g@��U�����Ij@�0�'��e����J@��c�b�
0v[<�J���B-ӽ�qyk�Z6��iB��H:+�!zxeT�S��b�-t���5�=_�/q6-��V⓫[ݜ.���.���:�c���n����.M�*��Sl>�"�eq��.���:	�Ŧt�#%I���L��]��ڮ0Nv��s�z�� �w�v�M�퍤T��#�h+cy���HOϷ/�Vj�:�֪�xn�,	�佻L.Ŵ���Q��z�go+5��m�� �ި,z��`�\�HR�@�叺�Hm�E����v�0V�tp^J[���4묰	�w�� �M-[Iǎ��ᱱ�ұ�8s֥�&W_6[9X��*��OdF��Vv�.7{��˝��jdP��khoB�����1�m�c�f�3��Y�n���\Ե%t�Wa�ƞ%<� ��&�A�n��ܜ��&)[R�ةSj��9ǺB��i��[�Z��-������{Ҋ��=�ۇEco:&93VD��D�\�$:��\�`�l�Z��Dz�����"{E!�c�m��erǲ����zS�w[	�+ �n0�D.����^Qw��'�V�)�!;�,����u�kX�gn�T���*�%�6�@j9��\�t�f�P�fAP���"��ucְ�l5�5�ŝ�5�akܗ�Qĺ�od�a}N��и�&8ˁ��i=��z�{Z,D/�.��&I�_Ln-���t��\X�x���ֹWA�5iL��_���\�DY&�5F��n�Hgβw�!�ٍuԡ�l��R�R�o:����w}�"�֥����[v�o �����n�s�88�I�]��ەp.w�/���˹�\���k�w$O��Bmb-��Ҭ��i@��mk��� Q�nCM8�/�,$�/�S���,�p\�壙��U9���I!���י.�m��g�5��P����r����w.�[���*�5��3N7umf;�@�[[�Ve@�-+�vMȠ�.�໢@�yc�"�w���|3.�uy��l}7r��28�mØ�xx��J�0j��c[�;nʭ����1g2�,S��� f�8j�1R�G-�u�ͥbJM���鵒�]���鍌�ﻢ{Ez�FvA@���u-�3�	��mګ�UG�lVe��#ي��K��f�l�]Z{���ԩ�]d�n=��Q��z���\yx��͵%+�ܫ��5V��1n� C���q�"�]>�j�(gs����Em�2��m�ǆ�:�|lQt*��K�̆��&m`������\8ϝ ��Kl�K�AU\��o��/nWC���D&�]�q_ht]h�ݚv��m���Ū �`�ݕ�B�ն�p����:��m��2Ɠ�`��U�=�.K{8����]�uw�n�˥[C�����N
(�gJ;{���fX��+��N����;m�+v�!�'�h�:��=���^t�0�5����.W{WL��U����� ��o�mA�(T�e_` � �>��#��%��-t�b�[�wM�i��a�(v��2�yx�y�=_>���JU���{W4�)���p�.G+�r֗p�T�(��N\�+��+D��p����ʲNQDQ�ʉP��2�s�T�"9W�qe���8ft��A�vQ��r�Z�&�"�T2��.�(��A\�\�
9\�%B�Թʊ(��� ��"�1�,��r����\��PEQ�r�r��#��"��E�ra��fQEQp�e\�.\��"�-@��QQDDr���r��W*(�E�E�J�Q��p��p�erN�*Aʦ��@��G*"��*.d%A�9AL��r"���\�˔EW"*�Tp(��*�.AZ�D��TUs�.UD�E�9vȒ$ �-��~�(
�*��B�B��Nrd�i��cX.��7�-�ؤ����c�o�j1J�!�D	ϰ>f �e�RcS� .���O�F���>�������C�9둚��kkϽx��,Sq'r���C6��]�_b!�w����K�M$�C0�od��c��_7n��"`}�c�OǺ���O��yE=�S��z)��,g�9'���R�S���s�Cق6��(M)������M�Illc�Y��nu$�m�����Rt��s:!��v�m�qsb�}��kqvX>'��lX�bY�{ˡ��M h0�]Y|`�
��L���vŷ1��3����h�1Σ�'��oRBs��Q�1�6��$T�11�<��:!�Ƥ�$���TM��W*'�F�7[�q�&.t0�Qr����T���:�t�{�_b�=pt��;�bn&�Vc���5�eHp7H隆��}��V4��u��]�AA�>Wf�ez�"��sD��\��U*��-H������1�'A���;-����Px������2:�Z^oq�t"w��}|қ�LX�'Y��o���C�IK�����~{��Q#/�0,¼���:�*p+Z�k��ƌ�x�fI��K�ek�a��,�+��t��wkp��P���֒�\�� ��I�+p�Rt�Nhm�̙�8Ř^�W�9�hN)�G���B�[����]__f`�����6���ћD�6�w:j۫�[�S�������DG�ec<��֦�����#Q#�f"{\<�S\�X�{"���]f�V�*�bjm��O9�C��ULGZUj�/��^g�Cڄ([Q�s�e���2�Ɨ�mI���s�8	7�zj�tUP��Q�6�F
,F�������������3e�՗��ش����t�VS�g�#4��ƃf��o���O�ʦ|+��L
[�no���Ԁ���r�1�c-�C�n�|n!VW�.J5�<I��!��#�7¹����e���}�¡��p�kg酪��f1}h�����Q�	����fK 'wC�J�p!B���������^�� ���nU��B��(xjSv�nH��x�FK�E�9�ʩ��S5q��E���=��P8���:`7_
�Zc�����m��se����R�Y`K��:�^M��=Q:�ݳB���q�U�}��^cUk�T^7�����p�k<��oue�~~ȳ�.����n�D�2��t�	\	��0yL�4�H�{>�����@X�{��L4v�={sS�OQ]N����{�ܴ<ѷx�������k/Ih�f¢�m>��	���LJ����,9P��ղ���F���JL��ڢ�-�+,y��u�ܡ�A��-2�rs��ը�/����;<�z��������w�Gmc{̛�#�q��4���,j"��[����T��d-!��DJꁑx�#-��<���ݼȌ/�ƈ��-�MUɼ0�ܰ4��f��q��������}z�/�螅N>za͙<���Tp�wV#��s0.s �~��K���zA6�R��6׼;�CDR�^���e��$�'�l�7�u�|������s�uL\�yѫ�f"��Ԕ�4Ǿ��;\|MEF�mC�����o�Ǹ�O=Ҽ3������Hk-Ků�>�=��Z�y�uc�Ds�F4U��F ��0��O��P�|<8Ⱦb�@�-�Y�vgu�H�����\���}�m���Ԣ��*�(����m#�E�1��U7�j1�Q���}�:���LB�u�7�Wҫ����$�F���~������%;�ݾjL��X�
�ū����!�w�w	��j�앷��G	�2�����5�)����t�������`�7��ǅ	��o�5%���X�.�-�����ץ�άm�w�oب+��Kz��6���nq�b�	�w�}����O+&��w�˙{�cm�"��S]AJ�	M��}6+��z��q��7�;���K2��*Z}���b�ymD������r�L�},J�sh`ATĎ�D}Gc��E�}șH�x�2	�X:x�?\G]S
�}4�0\%��0G1�����.�<q�>����
��@{LÐa &	粸#���:�����[y�H�Ϝ3�X�n���z�'�ѡ�����"��A����F���C0�ܗ��-�JE��u@6ա�g��"�'~mր]���F����#T��W&nsǼѬ΢��������F�0���p-��4!n킍9�����?��R��w'-<}]��˞*���+���������JS&Kn@֡����qk&s����e���+�}xz�<���?*��������\uҷ�ا��P[�ڴt��쮋��{�n���C{�a���ڳ]0]A�ס�������6Ǘ��BQ9)��R�,�]��TW��;mދ�mΜ�,��~��¿�a����n�xSgN�uw%�Cy�XR������sC�����8Г�	���} ���OoY�`׶|�f�օ�"�4������g�Nގ<w�<{��F���}�E6��SY�����r�$Y}�4�����i���Ӎ�2�\�=M������E�{EAV$�qJ����Q��Q]qн����R�^h���ꪪ�׺�2��Jsb�d�	� �]Q��C !�u'\"᭮�ɍF��$5A�v�j\ፕ�K].�z��*�=�P6���s�e�S��V^�͸N����y�pns�-�Pɞ��#�g���K�xk	A�i{U]>@R�qW��r�v�e�nS+{�Sڌ�����Of�)��v������S(Q�+�VQ��|+���躦׷�v*a�����S�6�<�r��v���������������
��&2�T��^U��y�~�s���J�#���E��6��(5S��-��Y�sn���rD�>�@ӡ���� K��P��ׯ���3yJ�Ï��
��늸t�8\)�|v}�:�o�Q�3�:�H�i 
k.�yD�-��<'iv�%����Qx�.�����͟��:H��gD4q��m��.lAت�j�\��mku.֥CIA���n	��GaB�Jf3A���a�1�d�%p�)h�rM��wo��$I�U�Ż�"zf_�kF����\_�^�<"7f�S���w+�
�첡�l���M��oD�z�U9��-���]�m��ʙM�}C=�Z��l���\�i��WS$s�����R���N��ŭ��al6f+��LK�P�gp�LBggk�z�N�2+�bI[H����;�zA9����t���0�SP���긃�]��&�K/n�����)��cmr;u�?ET��K�W������еa�NR���O����|��_�2�Cr����*A���:���/�}m����.���%�^��b��0��Ӷ4`�1��x�f�A�ͷ1B��H��K'�X|Z�<�Q���i?I�w�&1�f�V�ţ��ֆJX�.#T���</�쨑�\n�x�X�����I�I!�4�'8�8��	Bو�}P�T�2[:�W�MB¥_<�n���6�|<5�̖\��+����F���g/�[<>�ι�
cp�saA��J�v��]�+zL�k��h~�M�pm����\��׃�����mI� -�� &�qu!)�eK����1P�*t��`��3�B�e��N��P�]u�m֤��':dB��H8|&ˇ���V{~�;S;���$�~�.�AdK{�;�ɗ�?Lzi��;Yv���*~����}%�ۇ�C���/+���k �{
{x/d|��<Mhn��V=�5��1�oh~$�9c(<��3�
�§�-����ZR�|6�N����
.����2����_ �)F�g8�NM�n�`�|Y�#��@�Mj9R�8:�b�e�Y�M¸�C��9:��k����ʯ������]��7< ��I�'�t}?	��ʰ��m\U�g��a��|�H�x�E������L惡��y����:�P�@�&|*�xG\z���]6a�9����D�N���]�[}��]��������.�2��ԋ�xm3���6o�8�����n�s[CC��e�������]���F\�$���1?I��[="�)tQ�ڞ��r�Oq	Y�F��?T6�x̰9��L}P�\��C㧲�@.�#YOָ�����T]�������yld&���"��`ix���.0�8�y�d�R݉~+ϥ���S��>9ly�Y���y�͘�]�b�wzr5:ɼ,M�닥����A����.O�w��Q�+���ݟ_��a0���S\:�0���bqZ�au��6ޭ]�V�/.��*��ꍣP���C&/~0�H�5s��}p��qp
�{�x��d�o����+|>muk+yՎY�;�i�p�.��\½��N�.�_�c\)\P���t�@�ҍ�� S&��G7���3���#h��E͵/n	��vfju�c��b���3�5~{�<5+lnN�V�q�A0��jM۱V�f�]e�gku1Nl5sA�0*��95��j=�镦��W�M{t�v[���-��>�ƚ�x�wq��˷�N���_}�4��N��� {�{lq�<�dK�g����3�?,ck�=�z��1i�� �=a����D�(G�b�\�\��6X4b Ot�R��1��c7�_��2��D�p-�z9�K��HN��s>"5��E-�adtɍþ��0Z�7����&��P�Qb������J���qE�J��`.�rH�%�F�(MB�o�5%���cu�����޷��Z=�E��ßGdtJ8�7J~�몖mZ���R�34�tΆ�zׁY�OD��ȶO�����uC��If�Az��'�a  粷���#,�sc7/��2jhP*�g��;���q<beO��Fx��XFLdǑ���=[x^�ϓ|����5���*>I�C!��3ƌ&�mցq/Dق�0�#�I���y��}���R�=W睇j��Rb����%Pɦ�p/�h� �S��u����~K�oٱI�u��s8U��+*_�}Ҹ�$�}I�A��L��M�믭��}�-n �$Dڸ���1�Y#6+$�9[WiLԥ?�g.�w5�)�0=ck�uAY}��|�;SC�T!O���먣{��G-U�0v�D�:��4�� ݷ9h�pĺ������KT��*�i���c��0k�(s9A*��.�;�D�[�IW�}_}�DG��r}��$Mp�~�%Li�xD�x0x�?O���N���wSU�[�n�	��%����x��]�
��z����NC
&
xZ��`��a�����`�[K��]��e�[���I��8E=�S��a���w����mΜ�,��~���Һ������^�k�䧞�����4����:����iS�1��:m��ή�[���wn��ַ0�0�@��񹗼�R���=0�D�������UP����Zٴ�p�����\T�GdqhɑO����ﰂ�}N�L���NJ�� �s�e�N�a\�3r�㬭����y':�.L�!&�F}x�����(9�U)��AɆ:�*@ژ�-�������[w�˓��g�$ߞ���r(�h�VA�2!zxeT�R�Ąn-�R����V�ݽ�)l|�tu!��;M�����?Xb�/��N����iW�oٖە�m�":�i�^�-Ա��hKF/�Y���p8i�w�F>��3
��z���]-�^
��5�wR�w��,J���TL	Q$O=T��i�\�TY~����,�@h����r�:�#wٮ��W��6���AkT��	N>k{^�;��y�P�ҜZY�87���p5�p�2����k�\�S:�ͷ�r�V��5ЯUW�UW�ŝ$���ιp���<��
�\U�w.�>;�7Dj7�ق2����J��\���JL� ���������S�|�����.�9gD4s�;X��Gr�zSR�����'!�����(e{,�zL G3�*J��`�h��2�.��D9��^�,s[T6�g��w��	�W�\���	䨅��]�B<�*�B�m�|g��a[��ve�ս�{\I\��(�l̘=C��ք��|� W\�=p&~ڀ]����.%K�X&�g�4���̦-�g5"(Z���6�܋��f�� h�g��*A��d�@Ʌ�	�?��\��QoO\\-W�)���B8����YB�IՈ�N�3(9ٶ�(=�cB�C�u
̘"�}���u�S��u��^j.����N^����Ѐ���c����瀛ك��f� �.���ә��;j��^�"}�|d�w�Zn(�'M�鈬}P�3��䱌��P/I;z+t���iv�QR���8�����>�a���ET=r����X����dX��_s�q�A���WSl�"b8�RS0��D�Ԅ��}��-:\1h���S�jM;l&dv��A��'sY��ԉ�������rMX8�\f�Ӯ�j�)�oA�!¯ulr����fm>�f��n��̡SaI�{ݪ���(��W�N���MG$�G��r�l�:�����ܵګu��L����W��3[���D[���[Y&�ظPrSD�O<>6�����3�l��*�Uxƪ��sx�t�,����]tB���D���7-2=՛9�8	���|�����#��jϥ{_����O7]*���4�4�f�Bh^��H
^����;�Y��Lܺ�IC-��7Zq���ަ@4�s�%��$����C����O0�A��U���!*e�&�4���ϡs8�gZBІ�u<���.�\ޒ���ٕ�Κ\L��m�FeN���6Q�)��퓨����u�&�Z�� �Kd�TG5{}����<��.��QH�ɛ{����VH��`-m�#��8�VQuA�%tj����.���]���3�ܖ-w1�9�zk.��%��j\AL���z��Wt)��{&]�2��Ӽ��̟qQH�e=]�N?��]y*��a���
�\ŋuyu3hĪQBV�Y=X�9�K�B��Ӈ ,���X��7�^�a�#�7&�4:}��2
U����[v��}\��][gO9hV�;D�Wt� 4���s
\�vkӻX�]�/�9��t5v�cf�v>�-\ll�:r�wa�v�+8~Ȃ�n�c���y���2j앷B��x�7s��<L�J�ӘiaS����`�X0�d�]��P늖�IY+@�#̃�Tp�)��_�����O���B&S�F�&)�gn���1$HϷ�.����U�[Vc�ۥ����:䥝Ie� :�d�jv�\Ww0Y�x�=X[rV:+P����m\�뢀������L����`��e�ƽ�]����>�����,:�7�P��Z[}��Z٬�z.�1�7"���G�xX7~��^#��Jwly.�(�ݖ��]����:���z�g�(w��Iզ�Γ�=ђ�>N��s#����v��9���n-��]���˽d�+l({�cjuvv���/-K{-A���"�_;n��>���w�+������U�w3����R�	p[V�\K�1u�ʌf�<����֫����B`;�VI�J�Ղ��#)^EyC���	�I�����y"B�;y�pTfk�!�F2�ƞ�\��[K��c�!R�k��Z��\���b�t��j�?�l�%,���؝��n�aM2�G)�N�ݞ}�d6���SP��%n����}�]�S�s�㾫sQ"<�P�ѯr��b���+�m��p�]���yʗ]���S���S/��6S����r�mebAW1�ys�9�گ��
�q ���*�i��N\��E�W*�UEVE�E�AW�3
�v\��3��*���Tr��S�.29vP��+�\"


*��"���˂I�"�B�S�PQQÜ�l����A*���P\�

��

�WdUr�\�f�Yra��.S*�r��Q¢�AL(� �����*8QU2"�Uf�G.��2��*.P9N Q��������G"��<l��,Nd#.]<x���6���PUP$��DTG��P��Q-���=t��}%�o.��V�'w����nH1�!z�s��K��'Ԩ�"��vEz�ͩg[#��|�����}�|�f�VմՋ�Ӏ����ϪxFm�{�/�Ӡ�b;� �P�B�)��R�o�v	�iA��H�1\��Ps(ݯ�oy��S���u�Ӫ�s5ݢ��@R�??]�ܩ��
(��D���N��j֙�c{T#���0�_�i�����epY�P�x���ѕqhw"��v���/y��X�[��\7��uӟ�����[oh���J^W����P����z�J��Is��5dˎ�験�H<>��G���	���WfY�7	L0��C�":��UL演{�'����V,�g���Di��d0��g�o�aq�������Ƣ���w^���AV����q+w|���"�㨝uT��L�T #� 4?+��.�;C�%\t��u�c�K��MC�kU��-Qe�1�M���Q(Y;�$�ɫ�����~��m=�dBԶS��jk0���+#��<����^3,yDF1�R�rz����v��=|��]�6��J��C'�����|���xP`��nX^#46⏪���\���8w��;�l�v�\�����Y�ӻ����"�{	��\R;b��[���M�Ьo�y��f�ڝ��e��l�P[���5��nP��n��)���v(u'�3�j�4=�����f�����[}��.7j���jmw^ �y����v:�5�I��ۥ��cV��S>���EP:�V+���������E�t�������=���r@��reY�#���d@��TK��Yq����7>U%ב�8>�+��l���<@����t��5.}F}�LfQ|k�n�K��Ԯx�x�\k <����j�q��9��Hz�fp�'8�.uc�s�F/M�6��Fa	�<�ڇ�c����`/ה�O��	xa^u�"�y'��u��7_o�z�?ok�2���31;���r�h|��j��{3}ϬR�ി�@{o� )�1&;�Z��n��K�7��ݝu#T�g�eL��+5���$��FB���F�GamS s�M����0_\��a}ó�WeטS�^�f��č�ɔ�T)�e�T�V7���.��+�{s����T���կn�q!b�:`�#�Hiu��jV˞�3���e̹�͝ir �5��>�8�7Mؠ���T	D�窏&���j����s�L���}�}Ɛh����te*/��7F�򉝯�����doL�7��V�t�^�k���+�<(��Evj��I�6�o!ڶ�(�ވ��(^[�jsH����Fn\u/
��z����^R�c�Pأ�p�&Xm�C�����:)�vz��E׷�M9}�[���ED<gi�)�B�^4u9��b�|�Y��m�y��Z�-�awB�I4��s[ϙ��ob��P
�����5v�me*��ԥ���R�2�4���l%��;���C՝�����C;ڪ����¶S�{��=s�/�k�mw0��;	&�wd��bN��5 n+��O����sbv*c�9�����r�V�eE�,�.�Me�Kl�ov���k��Dk�"u������b/,�yѹ��z��x¾V���x��__�K��ᚷL�_CW�/�c$[��@4c�u�j��_4���ض��E�s�*^�>\�uF<��ە�I	�=�OwS�]��v�3�w�:?��+��:�(���ʞp,Ԟ�����6.��zQɛ=�u�VA"<�oo"T>��:��c��c%��>�!��L{1tYP�yz�z��r��6L���C������k�힢!�J��
�b��V�V9�p2l��9id�)xe��ǜU���n9t�uwK*MJ���p�%<�]�����!/�)�,���6 �B�a�Bn�`=*� ^���f�� {ӯ�;;i���K��M-�f���
mY�2��>U����I3��&�N��k ���Z�_>�+5�v��T��y�����ÂW�Zؼ�\q�݋i�HI�����o-���zyl�sF	�3�8k�Ы�'��s�K7���Y8���*1��\�w*L�~%��9���{RI���6_d{�l?�lH��}t�K��r����ؽoʗH�e���4��ƹf�	��j�:��ڡ<�~f<�,�~nRO�W�{��rMd��K�I�*��C���	��V���|��T%�8q�.�t:���+b���)[yB�q��9�9�4�x��b��\}yT���.ͷ�md�7�γ^�&Ƶ�F�L6c�G"a8���v�[Aܕ��=�����e�m9]�����9�v�!5F���mƴ��q���{��Y��_s廥�٧^��(2+�J+������%�x����ȗE�ܿ�O$J������3�e�S�\E��z���P��D�U�,�����J��Y'��
�V�p�Z�=S���sxtA�s�I/�����,�s�_UW�Ux���y�X����Y��{W�j�u���5n�����qf���'L&i*��S��I F�^�b��}}T��<[Ï�w�s�&�CA�R�SNT��R�*�����}#1TD��Oxev��|����v4��d7]��I�秱5�o�����;��,�np�}���Z�lwWI�󨳜�$�f�&2%���}�p��=Zz�����ym��1Rb��׷e�}�l]�Qz�����SM\�}p�:�m��p������o*G��Y$K�MR�H�s��B���z�S�i���9D�``���,�����S�3�`kډ-�I|�Z����m�����-�z)u_Z϶v.��o��1a?�ap`w	�4���;�>�r�ƶbLdT;|p�V5�8��<��<}~���LS��(��.寺0\��mmK��ڙ�W(]��e��zޖg��4��Smb\��֩JV���Kд�]:�g���ɛν�3���1;#��v�uw3���v��b�X,��YvX[�wc����Y��;�xc�"�R��ڏ ���X]6��OZ�m���q���*]���}��u�v���B�g���<g\˜���]"o=��ۮ��9ʜ7Ԙ�I�ݽ���	!��I�����y�5�,������U�K�|�w����~�]ו�=��k��2�]�#�0ݱJ�������+�qr�x�mя�.{���;MQ���4ۍv��dmtvAM\���os��=4z��U>_^ȯ��9طS�[�X�z�C�7�I�q�����3�M��-@������LѪ�9��Z��"�g:V�e�Ŝң|��׌���j�n����fQ}#1W�oj"V����eMv:�����޵pT�	=k>�[ׯz��y8�]�s�|���Oe�밫NI	��%�cJ�m���c��\+�ϛ�K���޸�{�V花�(�й��^˹��WI/g����"\.��(���i�4��/�o�z������W���qX��8�=��@��]3���jG9PP�Z���]�N��el.J�?b��]z���Qj^2���m��T;���o\U�]����;L��h��F^I���i�#ʔ����K}tU;�����r�@nG��|�e����=L%)�u����[-X��=��i�
�}c�K��>Nx��G�րB}�%U����T�v���˄5���lw}� k7c����N7p()Z;�4��K�����rw4��aN�H
�jw��k��zm7Mؠ�}�PJ:�u�X2Iƚۻy�u�Nf�M�ꇯ����Gk{��8�R��B���vM,���w��:8)xjџPk۬���0�&��9��;��m�Tl��޻�PMƹǗ7�LB{�;�A 㽸���oK���l��"^q��=]ʹ��H���V�|�T�:��sQ/�{{6x{�]�e�� �1�Oɗ��6��j����}�5_��N���Cc�rWf\Jy7�8,���U8���-�jֈ���ʍ���c��渲5���]�{E��n��*i-m���:��qK�Yi�H�U�����^�rP�=R25o��Kj�7{lk�g�-� J~�.����z�۵��������[�K���1z}7��$-�7���/��z�Q�7-�ж"���x�M��`Ot5կve�60Cgh��խN�
��!*O��}E�ێKV�03%��ڷp�����j-�;m�SW�5���U�� g6�GL�w�w�U�n'�Լ]��׵�ʗ��I�Y�:X�i;��ĺ���'8ֹL%�!�5�z�n:���Htb����#�:
��	=�D�T{ݱ����n���fO+a���\�J��uQ1ϛ۹���윸�{i�V/y�=ܧ�:�]�m�@��|��G\|��\܌�}T�+Ԑa��Yp�}K��_-��ՠhN-�=նN^����ϱ�i�vV�J�O-�o-�z�yЧ9\

V��B���<Kɋ7�7\��5]zEc��yJ)�h5�C�y�*!�n�9OV�K(�yU݆��)��;��TO�#��Z��Q_u�8�s��uC�r&w%bZ����	'{���2_ڧ��KE@O���ov������E]֔z3a>�].�m-���}��J�+��e�'�u�n�;��msT�[s`��v׹۵[�ǟ��7f�䵢�~:��7��d������+���{�l�͎�Ne�����ʓm��\�&��uc}4a�e����}HǸ�r͖L��	�}}�9[�^�5wz=�.Q�B�`�9����_%�1����9�3J֓ڧKu+��p�ଡ଼a[9ݳH�1�u����J��GF�r�6�B�Z/m�h�o�}%.a6\k�r&���Gj[Aۡ����2����z��}�M�Ee�Z����&��p�j1?��UY�o��呄��f��MvoDS�m��̯�b��[_^իI��'պg[�5�;���&��M҂�3ZUqƜg"�Fbٷ�`���u��r�*^ZN5���wv�=\��ҹEP������݁�����[/P���/C��ΡA��w}��{T�N�|Z�>��5�o������rP�����W��Ց�j\͞�;�|%�j�a��*.l�)}��w=Zz��pUp�1��O��˄y�>U�M�:/�bB��{->/V�9λl��WE�W����Y���׽�<^�0h����n���b��B�7K�g=Z-+���Ǻ9*n�Ɋ͌���S�Z������mX����>�w`���vm�ܕ�Ơ�O�V���p\��H�%�eJ�P܋k9 �2n.tZ���ٷ�E�9+ﾯ����w��^r��Qʖ�PƝ����D����!��H����Fz�8����:��;.uR�/��3�B���k����s����)f�2�����aL/���#�HiwT���MC��{VǙ8c{7��b��.���c���9R�+���%��>��+���R�߮�͂�u��'12��x�{����溧(��.�"7�ʺ��:���O���f&�{�)&��Q��آ�E��v��KUn���x���p!�緕q��$�Tp,��}M�����-M��O%uY���Ւ�Zԫ����+rj[��Y����j�E�����k5��$Qw�KiӐ�~�n����eo���e���oE�4�����]��6�ڭ5����Q���j�dk1�P�U�
�yy�������%P�e��@�p�.R3fS����P�g���M�0��F^$�q�Z)�;�ӮU�=�ᑲ��i岍��M����G�n_X�mP�Uvwa�&���ȈMaf�,����4�U3n5��}�����	�ף/��@�K����|��.��)j|$+eD2B.���OD�A����"̑�6o��Σ��kf
��1���"Y"�yVn}��V�̏'NM�4���c�3����ѣ��poC�¢^���%�)�)���Mm����wK��<T��	Un�4�2A��E��5B����ts��w'ž�ao�S�f�o��:�Z�XR�)S�Z�o	�K8"�,{{*���6�P�8�q�$�"wz�ҩ2{8���W�i�l���+�%0lY�Ł��'ـt�A�7%�m�-k}k�;ݹ��[��Y][�Z�z��j2�Kˇ+��v�r�Ѻ:b<ċ���Ƹ����G������ͫ���Vk�F�U�.���m�ڧ�u���kO���D��(C+KXZ�D��p�/;�"@�[�of��춞��d�4t�ۀU�s'X�PM�|�㐡�5��C+4EЂ�3x��u�eF��4$9"օ����#ҥ}� sM�nV^O�R��Q sr�|�{���;o���B������*�݌n^I���c25����wJ�2�-���������δ����gwj�m�u8��0"E]Zn��v�Ss'}J��.^��u�j�Ӗ���PñM]N�qܬvÊJ+��&����;�f��KS����$9.�Ҭc��,�u:��t�+���J�)H57���B�4j޺7;1�o-;��g~����n�ܫVʀ.)�j��I-P8(�Z*�(�9��s�JW�&I���kI��6̡`U��1���	�Zԭ�qU�fP]�H������h��謱2��@�b�	D�n�O�)�$9aZ3~Wg��e�{��
�Ωe�h{P�]9�ڮ���w�'ښ�����h98f��z�]�lҭ�"D�N�l��@�T�ݳY� �L��-�j
W���8݅G�6uj)���Ԣ�Y�"Cv�mf�wj�}5L#�w�w^���egg}`���Y�@˂єf���Kb�S��8+��h�Zj���7Y�n�����H(�2�Ek�	�T�U��q b�J������;k��:��f-���`�56��Yg�]�)wY������ʶ�=��W"�nto�LỤ�^�G��W� Ա�oJm�֭�/��w7jռuצ�g�\(�+���͗�Z|�K_U𧕎�*-H�ʜrK���&��U����4�e�٩�K�7I�ja}����]��}���6��VXcpD�[�>�K [|'���܃�X�2���r�I�yЧ�NT-R�Սn��m�.͌)u;\������u�}�P(����UQ�M�["�	aDW
**+R��DQ�K�2�(�T]�ʹUE\��C�g�ʥYJ��#��,�W�8CL�S
�e˅��:d��0�:r�8��Ъ�DUQWYT�A�&\��U.'NU�m9ht���\��2��N�vEQUSr��E��G(�9r�e1�Er*�9Eܴ�D��
���\*�w)�\�� 5��r��
e�q$�g"*(��tȺ@# ��ex�*�#ı�" ��EQC�e��D�J�v�W&QI	���9E�:�\�1*9v\��
����.x�(��&E4�B�lJ[\:�[�W}O+�N�o�7v�3I���t�F���n��N�;�9��)acӝ��9-�v^\]�ȑ�S`�2���}E����iX+?|�V�q�F9g��Cw�/X̨/�b���6ڹ(�Nl����;��	�ؚ��ʗ�'�����5�{5O9q�/�2�O�)�u3��#o��w�2��:�\�1���2^>mf��y�wmS�ʥs7Z�*�)^��8t�$0�U���ާ�:U��yM5K�؝c9'{�RIܧ�k��Z�S���yU9�>�K�y�E��z�ՊV)[�B�k�����Okz}�*>31 ��(�<�Yo.���ٗ�U����4�A��c��n�}�9e�i����v()��t�P`wip���Wc|��Zu��8B7�x��޹���^����y���n�Pk��*(���Y&s\��)�w:��y��ܵ��9}�[���C�q̩P�Xo�Θ3SWY]��w{�^���}B��F���3Lr�O%l淌��B����;} �MgT㨫l�6\�"��u�z©J����G��#��V�^ty���n닼�ն�k�[<��m���-�n�ec��Kz�.w+:7�>��I$�����ۯ��u��D�4F�.�S����/���T�����մ�HA�ﾏ��͑ͽ䌮>�Fˑ�QA��I[w�iMoԹ�m�pa�9B�dg&���5�\qȔ�
�T�T@+�u�ǧ�^�N�tn�x.Y��A�{qr���rVn����r5�E�#ë��#���J�֫e�:Ʀ����u�=_{*մ�է��f�q�N��-m@�T�Pq*݅{�<��lcW�)�EZ��om^մ�ΌN��L�_5xr�Xɨ�qٱ�œ�w�Z�Jj��ɛ\U��������K�i=k>�C�#nhL�:QGc��7i�Y���vʂ�`<u{}�[�uҺ�����~�3b�ecaf&u�Q��f�Q%_,��<�ۅ�2�*��>0�{4N�_	Ւ�g�.<���򶺯[V/��M\D��O=Xz�wT�@��Y�˕��b�ױ2y�,�Ȥ\�\�w�}Cym��/�\�P�
��EG��ޥngA��ج��Q�N�ѵv�����Cź�of��Ҋ�9B�e�8oa8���t��W�ˇ.����m���l����-���He_����X��%X��ղ�uKx��۸f��N%��b��Ճ ����n�kv��y�;�J����6_Ľ�������1�-����/�]�[N�+�\=�[O;�9�����Y<�Xc1wye�k]3�B�Þ��|�Ot�R�4��=��r��ov�ٽW�f�\�z9���}S� ��c�7�|������q��/f�&6U$���3���e�Y�!����e	�<�Y�>���/�][Uik�Ȩ���X�Ю��o�隄B���4}=+^\h\�q�]��N:���[̚ٽ͗��3�+�r&�if8��rV����֣5Cˠ�d�}��s2\s��4�J\�l��h�L'H�D���M��u�r�Wl34��L��r�M}x���x����������@��c]���r�3�l���n�jD��D���fTKǹ�:��ZN���m�9�o1�9b���MF��VuB�xm>��	9[�U}T����o�y{��9�7�!�h���KV�JK5q�ᛚu���39��{X��\�h���Ž4������R��T�{j��oR��l�� �rj�k���%\���n�G�H;2=�j�#��G
��3fΫK�E�_,��2�I6� =Ku�r��������k�8�������3�Ǟ~�7��3(��ᘪ��*���Ԣ�����|<�#�ds|���Ocu�q�z��N�,�U�}3���p٠:e��Ow���R�|'T��Q�͂��/�nިz��Վ��_�.�4ܞ}��<Wf���{��])O� d���
[���D�}js���t���%�����)~)X>yVcϮS�Oo�v�7�����Z}]1}��7͹^���I�/����uQ�G�ʳ&Y|�)������X�*�V�������������k��aL/�����0�i�Oo���!��9]I�=^՗�e�D�i��O���:�3��+���|;�*�o�Ǝ�;A&$���z��u��q��o�S�u̹�B�`���:A+�h����+;.IoԚL>C8�Co`:ekﵸV��LE�p�J��t��*G�̛:��Q����erq����뷙t�aų
��۫�=8�58jLN��J��-��0j<���꧛D�Sb�u9��}wOkE�*.�V�w�"�Vڹ]���mM��(F�q[:���y�o�g]l����G���׊��<����0`��_D�ɭ��!�˙��Ì|�EX�`�� W�5���$n@[
ٞ�c��GۓR�Mv��v�Tj�`�.��:ƛ��M��Q��Vr@�V?��n,�k���������s�n�����7�Q��U�k/�[fy��jہ����g�5���W�$�~����ty�6�+�זb=�t�=�=u�q=��_s�.L�̯��}7�Q�u%���rFT65�4�������&�s��ഞ��η��٪yˏ�N�/�^�}F-�ft��2��ʉ�:��~�\(���}/6�{����*������wcK�㊰���;��%C��b������M5�����_���}[���=��:��V������K�Qʡ�42�8P��m��QO� ���>���Y��>2�����m����s����b��4պ��^xݾ�	NY=��۵N�l�,��{oy@�iIk����ǩw�6Z"���fk�.{K]mK7�er���nVf�Ui>�]E�Wjȕ�X��
�,U'�vo9tC�]�P���#ì�3�u;����:�r�}6r1"�b����U��u���� j}�����z�i�n$,ZIPGp�N-�NyY}xS���*���tv�=��)��Z�gφu<��t�����y�U��RD��ffO'�Uuu��|������\B8�r��uJrf5�;9�sd֦�y�r�	��ȍ1�����r���q淐��5�#�l�}�kWi������i}�@ўw�v�3�Q0�G�MM�U�y��	\�9[yB�Z�Æ튈T�T��\�V���_d��h+�ֱ�Mr�J���M���/��q���qq<����#���P�C��m�m��Q�٤�:5i�5�_s��q�k�7Kk3�y0���J����zWo��[�*�ڵiKیN�,�y/�͠���E:�ȴtO�y����Bs�܎Ʈp�z�E�s���I��r7���7s>EZ!2���꿳��V�f�oWs�qx���{�Τ��د'��z�lQlX6������B2AV����{d�I���2�4�a��n#Y�Ӝ+�ʶ�NA�RW��K�e�6C�{���wx؁���q2zu�zٴ�8�к��};�T�ƤW�U�㮂DuקJ�w:�{}�z�ե�1l[�3�b���t��.N-泯���E��`���}^��[�!��z����ws\�u�LdKMכ	�?�;����֨Ωo���c��Ԝʘu�s����N;�W�Cyp�}�~~bk�L��B{��/�o[���P���r��Iި��NժW5������x�ޞP�`��T������w�ԛ��9�=����KήSJSƃX��{��{^�������,�Z�v�p��`O�Y�	|��Z�S�/��}���>��.�;^���;F�r�]3��o��{(H�U	��1�D�b�ѣq6aw>�ۮ����N!x����m�.Y��t�G�E��\^�ex]�����r3�֠�$�S\����ض3�?6�Uq��������|�`ڱ<����{l9:Hv�޺��N$n+��/+�j+/13Q�y:Ȯ�=���*&�B�H:f�et"�[��$�g\؃Jn�nr˥�S�A�&em���+��-���9��u�Ow��%n�)�{�5v�WH_������55�'.�g/}�t�Q��L;�������	>:n5�+�uU��)�s���)��^-��x�5F����c�g7c��"	O	�X0ξ���Z��Hz;�A�/�z��"��ɝ6�'Ϲ��؜2d#�F��+r3{�Ԑ�����W�P�Y�A�P���E}s|��\Sa����9�R٭��+�|��׌�_�Ԡr�z��6
�U�痣��X�7F2�Ϭ:�2�rPr;֮
�q����nzn�9x렑|y����N��Mz���ؒ��5	8�{
<���KM]������(�������z��n_���H�pmN˨���/�bB��{�M5q���;�kڹ�&$����@V�Y|q�IJ;���Tr�[=���o.�ܐ\�ķ��ޮ�7�+��Ʈ0�
(>UR�/��3���L�ыr55n�<YYu�K��\z]�G1ɞ̨�{�Y-�z�h]���_���cpFu��4{#��5��vZ�hh�W�=+�y�Oz�~|s[�\�+D�*oonV��nfb��Q%l��9�K]��h>8�s(ΓX��8b#�mSɩ7 �]�_��z@r���������Z��
W��E�!���]'��o ��ƅ��Yj�$ET�Sݖֵ��u<g*]%p(.�xC�8o��{�R��tW�ܜ�ܐ%＼�Ö����>o�T<gjS��B��s&Ӷ{K��Y���>[ym{���ȸe$ҿ�|�3�Sob��h��3"�jY�Ѯ�N�,���bGg�]1:���rQ˙��|1����DNR1"&]�Z�_$OCJد�q�u���$����YM����@ȵ�>ɭ��}�'���k�,�͙��\a�!�-m_��ƻ<�^tڟh%��ܓ��{�jDR��V�bpͷ)���E-�r��I��ꎚ���ԛ���1��K���$^Zq��G^=�n����fT��4*�X�֒��q=�����qX��R�$��u��;��N6��H�!��N0zrE;ǧ�}x�p�~�t,գ@TEf�����a�,F3+kSʱ|�f�:ft�{�I��IQT*>2s�/��A�ZZM�2�D��v����6�Q@GeM�ye�y��k\J7���j�
�/-G�2�Uf�oJ����z��BE$9�5:���luQ1ظWǟ6����]���"cv�N�}!]oR�WV;*��w��s���@�COv�﹊7h���N�t���q=ٶ��z���Lf:
m�3)�U��-��#��X�]6N�]�67��m>�i��Yˬ�X�WTes,��}�t���}�����;��^��C����k-�{M����AO�@���$���[s���u�:�n:�T�j��cZ�^��n���]�YKe��d���?g~��'��⺖��r���Gn7�)�:�D��O^1�>Ks����??��t�Ak�⺖��I�p�kq��7p�<���R*�{�D�v#�7�3��[�H�g�0��B��:���F=�XҞ��-���q�h�7Ld*g�.χ\��j/ϯ� �k.�j��q��L�*|y�J��F�ؔWf ��5{-'�F��iIʋW\T�kF����0u��\�V�BK��4r�t>�a��j�)�fS���u�tԣ1�zΆ�pq�2"��D�YYc��g��9�qU�So�6*-���=�yf��;&F]��|�K�cS��WfQ�y����5��@uCάq�ݱ���]��k�Rp��b�5�훤1�'K�sb)d�v*�߷|qTC���9U�Jf+��+@4(��iPdk�{�E�8�k)C��:+�c�%{�=La�w�]�>��U/���q/kb�e�O[��y(SY�^]���cuo���G��Њs���;]�a.���n�L� WTG�a���݉�%SB�<�ޣ$��K^�8���?�����I�u<��w}9���$qW�k.���w��z홿w׀K��kq�]�P���:�wU��i��&����?n������d�H���I�e	D�3��ۜ���F�O���iD��N�^��+�p�&M��ӂh���I⥮���#5��Ov��@�ZL�=ʜvzV��T�\n�|<U�{pT#��z�v�}@I|�!N�e�[a�ݪl�]@���/���M=�*w���bP=v�eq��ﰨ�6h�@��n�-��y�"�C�5��v3�ǑH\̜�8*�T	^�=�3��	KU��n��
˕�Y�	�w��(`��Ogyv�s�l�K$mKHogD�^@�wnSǗ3ǔ���@yX�3@u�U�ly�ڍ�EZnJ��5М��ˮ7Ѝ�Tz��'۬�1�uܦ��z�=�mB�B��Ut��3p�ۧl�rX更ﻅ=Q\�Q����ob�{O{*�e�Ѣbw���آ�U��M���]�U���e;6����:���0әx�"�QK��t������p`�d`�N�c�������x�Ȍ�]�T�,5�)�,�jo��)a�S�ɮ�[�P|��Չ�Z��<o4��(&.QD��{��o#�ؗrR�����X�8:As�1+V��ϋخ�f�_R�*��Z ���OP��췀����,���}�J���K��׹�٦�u��!&�fةʜ�����c�o�]�a&�N7[�)`S4��Ì��-U�LJ�Y\�����v�������U�Z�� �1�ۮ䯗��M���l��b�m�]����+�c���Q,��Sx_Q����ds���m�r\!�z@�\iwE��C,�;�'b`_ua�����Բ&�MD8��k�P�[��ih��+M�	%}Cyl� Wsr�6�^7]"W+dW��al�׻�N���V획W%E�=�)u_nK�wbf�։�4h2��T,쾻P�ܻ�A�w#1ݡ{B��Y}������*�N�j�TK�g\b�|n����/;B�v�VR��ݸy�і)g���땬�u�}�gs���s�޹��"��"��$x��v\��p9D�Nd2��M@��vG
��NҸ��"!$��]P*�����ȇ�9IvY!JШI(�"�Je�`��\���'-;�C�!�"#��.E&HsVUT�5aQRIET�ULN�-Qd���ˑ		�%J��g��a&��j�vh���Vl):UMT�L��4�2.P\��*��N%���@��q&��\�d��\�T'��0�2�U�����T��¨���9GQ ����#���
�%�W.<g�D�E�쫑Q�J���]Q�IJT�Nd�X���'9�+����PU�r�ɡ�epI8Y�p�T�g��`r���Up�á��9 
�֔����|���䭎�ͱj�	@$	5�6�J�ל��ļ��n�t�[�.��d����*��C@�&L����!rJ��Z��"�!�M�I0jq��G"b5����lb��_�+/�'�ڮ7}�M�O�{�_^-�����N���o\Y�37�8gS�!�a�u�ju)�S+/"^=��[_^իJ^�pʷL��l�Q8�����o*Zy��s��g	t�	9]��X2��:��vT�	=h#��0L��rM�QR)�gSw���0*�B��o��ԫ��o�1]my[UƲ��<�RT+��z���Ǚ;keA�t
gǺ�W���A��C�+�>�V�}�	�p�.ld�����OU=Xzhwls�:�we�����e��|��ƺ�/�bB�Z�m>���낳�aU���X���׎3�u�Hrz�]�Y�K�+T����7�C�m=�9� a��%��7Ic�R_���TC~"L�:�:�MB���m�al؇�w,fsɲyhV��/�r��i�n�znkt�ms���Hd99Һ��6��6�=-N�Tkwz�R�֊ u�N�jy0��@�R��
\OBvMHk�jX����֯�7Y'o�snL�D2H!������q�bc=E����3���j3��Y�Hr���h����>����{�܎_���~n���A�M�0w��=7�!pί�3�.��B����0��W��+�&�,��.�r�Jx��5[ǻ�9�c;���v��L�B!LGH]�A ���y�w[��9/���O=�2�歗��8¸g"[�Pg��O�{���ϒ33y�i�������jy��!>��a��q��Ȕ��meP�C����[��I�L��-v�{m��7�i�=�2یs��]Q��df���8��}фL&:E���Z//"V=�ز�f͓؋��e���]�����ᕅ�u3���G8�u�t[쁘��ȕ�*�]��2+��Ѻ���)֥�����T�����k�.����4͕�WL��7_��y"�[;���rgU�\8��Od7[����us��fL�]p�Ow�����=�q^��\��X�ۥZ���ZM��V.�A
�|���"��*�%�X̵}��}�ezO���r}t_n�j���˩8����QՖ�.5+{�"���uow�G��:Mm,�TD6����;6�"�&]���]�1��f�(m�d��Z�_OC��~�\*>lg��W�6�oz�z��NXkae�k��Ά��2�ӀR��=_J��2_\HTB�or)��%���l���.)���F�S��Y��+@�-�ʤ�*9j�ꁍ;����{�\z���u�i?[�cetP�~�$@,��0*�)W�%�j�g*�q]�cM$�q�9m��=��rۂ��XS��z�3��P�!mt�'�=K��(��}��"6��r�r�.ֻ�x�TU�$т[�;�׹>^�jk����躍>�S˃���p�寷����{��h�x��C�r�W5N�&-1)�Ȝ���{�Og�}�N5ymN�d��RzO��q�m�J����n�tOo-Il��/	�����䧲�88�}�1�~�k(�w���I9�8�/S=W=hT*g�}C�Jܚ��k�ս��.on�6]D%'-C�tҬs9P���B�CD+�w��`�Yb�C�ʛ��o�]��[򖥖8�սC��l�D���������Z�]-��;�JZ�yz��E��	N�3C8���ۻTY�Ъ��_ʸv^��U�֫-�Q�YwۙN����ỦY{�8�,���Pۍw��F��&9��ka�ϧ�*V9[��٫v�y��w��H�o*��N���jہ��s0�Y�c�����em����	[y�[��z�S|�X�y��i�^8��]�z��TCw�.5���O^#/��7�{�:}�K�JO^�_�^w������ӟ�=^L�)��s���E5Ew��v�ih�*'꽾˞_|1D�.�62^>��7��W�.ܺi��.�U���u�
���KeG�˃�Q犇�1�TQ8�P6��͌���Ӷ���{;˜�͸窾z����S���Y�ʫ��"s7z��	}�#~N@�Q������}r�낳�vQ�l�>F�wC��n\�3���;7���9�;u5[���OC����N7q���n��I�;�үcס����U�	�ܯ���Kf���k]��gT<��?���|�S>�N��˄����U�7^�]���V|Rm����efn3^���^�\�t��[9��mK�.R��{>Y�;3�	{��O{%:D��??���q��9�o1%kU���5g]�ѭ빹��n�V�ikwec#J�Gc��yL�5�Yy���пT?�I�!���Wܵ����!}��	E`��B�z�)�i	��3s�v���G�	��Y�"ad��V�Į��vUM�\�munp���E�5�=!u�{m}W�#�=�-��-�1�w���D����А����,���u�=<���7�+Re:r);sw�e�}\�k��:���BI�Q	��p�F���1���9����y��kݐqש�{=[�-\�^=��|�������9�,�tN�����_ut�ԉ�$�f�Of�75mE�Z�J^�p�9G��J�}s�o�6�\�q���^��E�����|Vϣ�;���K��C�uX��t�w4����N�Տ5:�����ۡ�_^�e�]*Ն�SyN7��z�H=��<}�7��oV<��]����5U_����+�҉�_K�5[����A;ډ���Ũ�쿎l�	>�{E�B�u���Іr�*��t��E(�8ݪ���&0��׮�郄N��ٍ�u���r6���IS(Mj���m��U��S�w<����L�(��@](����-Gz!\�J�[��'C��;��-�^ʡή��l�)}�'�����V;��� �T��l�/�|��jL����U烮=��
Z����h����ش��Z���(JE�`�,�H+k�=ľ[�JƷ�CyoCچ���̥�ۙ��OKS��ʝ
1@�*ʢ$�Q'��W:�<��[��kP�VAvrm�kH�q�NW��w�_od %�K�#��\*���i��~�^�u�v�57b�'��j���\�p5�!S�h`q�u�@3k9m���kR.����i1z�gpT6��_��!�؎��羐����.����;�.{;!��xeB\������4�0(CƯ�]��ʢn��e^�<0�J]%u�bj ��;	&�.5�qyE*B�ÝwܷZRc�'J��
�˷���_^-�v�Tk�N��Ml��~9p�����]n8�jݙtw@�p2��\�)��R����<����tw6��{6y�����f.�d�5���k�'�AF�l0�u�}S��ʧ)��&�Q�-�jKsy�^��?y�Vdo.�jޥLS>�;F�]su��/��m�H�-H/k;�C}��q�b�􊯧����O�R���F����=&�Kp�8k��r�7��9�-g��~�BNUo�_A=!���{��M(��p⭤�]��Y�{r���mOû(�wT;�{���u�NR�����ү�Syg�[��'���#�v�)�F��us�����t�����b:��4��7���+�Q�Cv.y�`��}/�n�2k�1�y�(�w��sĐ����s ꨗ=Q*W�%�bAf��)��7)�ܺ�z���L��n�'_��{Qˀf��0*���G*[)_�[�*�@qIM���wܭ`��k|Z{�s����!h0T��RR�/��o	���zsT;K���kw���kn����[p^7'}>LJ��N��Vy�4���^�jUe�Nꕲܾı�P�gW���-��_���I;&�����4Ӛ�40mM�qJ��'N�s�:��O�ݝ=iAN&��Z��% �����6��b(��Ri��=�{��9�����q���۲��a����X��Ebp�"��Anb�m*���I3#��S.�4�&��ؘ��$31���FU�w��_u�i[9�r�͇T�f氨9�e���jz��	��������/�)R��I��6q��ʅ7�k�Kʥ����D��*ٯ��?G�����j��Jy�Tp,�����qT�Y�y�W^P����g"~���S=��zbk�����N�"����ʞy��Tj"�`�6�]��V��'��kj ;u��cC�������w�u���]��녑*@�Qs[ÌOpk�稯1�3�����/5��k���k<�z�|�l�ܳ�.�y�ի����q�gm䨆�* �}ʴ���8�1���Θ���6��V��X��R�_�=k9��3����#�������z�����A"��0*�����TQ1ظQ�͎d��wG�)�n����2I�9�&���c[=qV;�z��T�}P1�N֗N��ځ,ٍ����C�Q;�Q�m��;�y�	[����)%�l�2i2�qf�N�k��r����E�D=5w]3���F���Ǻ���uS��_1u��x���2[:�r�_ή��y)�-���j�X�\u�+P7���S��-"3;��㕒.Cnv�܀�,U�ʥH���� a��Nr�h���窞�/~���*eY��m)� �y�mrԣc)�v51P�7��}r�낱���tef��W�Xב�ɹ�Y�gS�V�j���Y=jOn�����vH��ƇB�w��d��>|#S�/��T)O-�k��zm�N�oof�'ǥ>�J\�P�oI_%7�Oܵ�ӗ�#��憹k�u�[o��P��S��c���g�!��Я"�3}b��4釮�aۥu��Z����kY�;��{�(��;U�{m}}�/?B���Ӧ�V�D�ю�j|�8�B�>n�ɞ.�}A�)Fͧ�|�C�[r^t��e���}��O��$�)��ЎDƸ��F̈́D�I=NOdiܝ�'�6�3���ŵ�V�9:5���n���qH����-� �O�Eݳ�j*��v^����o��{ou�gA�^��IN�}�pL�YA�J3J�]��~�,p�����{PL���i�._D��{��r�f��KI516\�����RA6���GT�#)� �Y�+�)xv���[���W�ʦ�5	�����I3i���=t6,��ϻz�yo(�f�E���EV�����o*.GW(��o�j�n�r���}��m�ĬڟE�s��v�}��MmosV&�8k���C��zb���ǰH�<�zqfK�p�xQ�h�j`�r��7z�G�w�<}��o]{�UOIx렐rtn�k�ލ3���X���ĕr�p�Dq�Os��KM_��6��_=Zzhw=��9�s���*)��*��_�<~z:An�O�"_>���Ÿ��gp�\]M������\E0]`�=�2�\+T�kyoCyqCی޾�(Z�X���o"Vss�_�����_>D%�'��+Y5
S�b�5$E�)t�&�H5o��i�N[�����!(����].��K���,��Z"�\)����}��އ��K�P#�ޓџ}�q<�e��Yy[��4��۳3D�������#C�r��O�А�x3SoP��EM��.s�3)��⳥�Nb�f�p�����$V��H���)d��e�U7�% U�nV-��e},դ�[�
Z���d&	@�w�����J�v.�V)����
@z��{R|���WVO7n+(+�;�Z��d�)ڂ�[�M�d�Ot9O��'�cnL�W���(Q׶xɜӤM$s��?��r����ͼ��N�櫨&GM���IBd��TW*�j�j�۸i�8EwJ��ϡR�o='�P7���]�M:�8zl2�K�9��r��7�^��čD^n}�C�)NȮ6�;dW0i`0�-�� ��kuԲyب��V�w#�;��5^��Ӝ�>�W	�r)q�K�aP�5�PtԴ:昝9u�����a�[��J[�7���Sˬ�l�T�&�n��l�1�e�|�ˋ��4�'ʶ�c�8KgV&uY}B�t<���_ã�7��y�7l���9�W�e`�2���N�@��� ܻ�).Nu9sX��V�
��nm��/.��f�U�q�\���`������I �N�WLP됭*2#�FZ�˽�z:����UҮ�N�=��n7M�W̞��#���R��wH<�K>c~���o�_f
�*TS���Ȯ.̧
�vCɻ�NnW;�	Y�rև���������K�h��V��u��L�m����I�*���� ���#;M_p������_V�J��8��
ܖ�P���p򣭄β��3���{�"N����qmJ޸��S5陹W�.3�-�X��\�<^�z\��5�c(V�֯��N�$s+s����ޗ��ZvX��9�v�b�E-����ÂZ��b Xթ�B�w1t�a�w�DeJ[�=
���þ	���ے���c��)����K��W+���#1�iW��ӶB�\�t�Xv�v�7��$��ͥ���Yiw��d.��X�9��e1T�_6��lp�޲C�G�T�8�ZI�p������;�m��Et�R��MH.�Qս��y6*',A.Z;��jFD7�(��j�o�E�
������ԮW��V����2Mf���_�ݤE�.8Q�YN��t��1a�Q�QP�*�^�h�G�V�E�l|l�%��{�� ��`�P+�U'NP8�nu9I��E�4�=oWi��龔���jͻ�U��Q�.�@�3z���7a����ݳT��]��,vN�<�r]��s�A�ECCwB4xf7�e�R�s �&�ڼ����s�"�k�y���ꂐP�{���ԾN$*nqW�. �.�����2N+�HVte<J����CI�Inc�u���(�����I�k%5��dX��uh���w�t����oT� �,�&.M[����W>�\a��T��o'1��x�[��id޸�r�k�w� 5�=���Cv
啻[;��![D��Q�E�'k�!f���>V��*�����9T,��avE���d�HB!S;I*�E
�t�:.Ax��ٜ��*�9�<˄��J�˜�!Q"����Qq����g"�51R���"��q"��YhER��\��&Ej$�	�I�F�!f'*�FJ'�Z��p�c�'��*9gK�GUPL�P�"��XV!ÐG
i\E����*��#��X�i��X��E$�p�"�'9a	Qt��(�N$ɔp��(��C����4�L�M2�#1)+�Ι�)�����
�u5D�C���j®�'(ԪեfIFT�I!"����G;H�*�2.]T����Aɦ���np�-(���H3g�t�����ޯ�N\���zj]<�9�mf��K����_h��{��}�QK���.ǭCVGuX��K�m�l�kL8lcyZZ�o�w�7�fR����Х�p�kX�ਆ�ډt�qfW;�0y��,ݼ�꭮CC��sS���%Kxe%�0�4�0���혦�x���[��V�f���J��db����vM}ښ�B}F�I0���4����ً�ɞH���q0�N�����)��^-��x���U�+ک��}�^m3z�9���.8�39Q��c�Z��Y/0�y�f���ĔTQ�3�6y�sT%k�|�o�k�t��z���y�A�P��U�HrןVP}�}�:\�6��#�gZ~�/ݲz�������S�Z�f���\����Fo�6ͽ�n�ۧ=*�Z]�+0��pS���okηW9�7�4��S;��Cz�3\���&�+�P��b��� ���}-4_^<��|o'%eMu$���f���P3������c��gp��<��F8W��ٸ^엤we9ƌk;�ա��k6l�3U�t9�
v\�fd[^�>��S2'�B�#�
yg;kG�{�̌2�jfXȺ��eiZ���'��l�-˦��gc�5Ǥ����(͐{*|9�昁 ʵ��7b��u��岺�_).N���=�_<�J����`��Y�ʹNDdV�N�����w֔�t�G,�z�\���Nr�AO�@�*ʤ�Z�Ȱ���ym�쮬�=On���{O9hv��f�=W�*5nE�{�2or�+�����/�,kS�O��-�A5��ns����=%ݹ3�_[=��
�{n��+���r�b��7�3�T�%[�6�m�2H��3��B:��7t)������.8���o�4����w|�(wgB�^rxږ�|]�H�<B�	Z�nMF�t�JiħJ��[�k+wZ��-��q����nبT�T��\��%;�LNټ����^_g%"���W�j�ZL����Fr��<�L[��Y/11��O.����8��j/�uZ��;�N��n���Wφ��:�Tw���di
\��q�xv{xV�I/4�X�0�uW�ܕ�{�F�5�gM��<��Oh�򮧽�웁Q{��S#�d<��o8���Xn<H�6�S뮨�E�K�n�^��ڻ�1���P�u}bQ��n�ͳ�+�k�ݩ���J��;��E}T��<�I��k��,��c�h�f��-,�)��s����� �τ�_�*���꿩c�pT��֯.��C9�1�v�(�O�o����	�t=����W��N�ظ':�<s61֜M3���j�v�;k\6����j禆�T�ީs���H���#/v��K仔	�ȟ�.ns�i���>[�?)��8��`;��
�}F�*�!��쎝�Z�����v�-p��C��})'�v�t��z/L���~2'��֞{�^���W�^�|��;�D�����r�3�JljZ�9��AG$%�W<Z!T4�i]�)�P�̱Y���^Qr��Iȃ<�}-��Yu�N�Pr�X=���VǕ+i)A�~X��9ڑ�ĳ����'ơ���`�@Q�^*��h��+���Z;���bb����v�λ|QG�l&B�آ#�/��< ����?끸��dB5�ߔh?b'� ����Vj��'o4:�TM�%%����i�V���{q"l,T�a���u�]������6������}�q��צ��l�Ɂ+�J�� �V�8o����T)M9٠)�u9w�^���m;]�g)4��x;��z;9�J�Q8N��W����N��#i�-�����R/#����%���A~�*�f�9�ڵ=�����fې��2�h=�)�Ei(�w�J�q�fI��:]>��q�9G�"3�_'KK���*�7���O��B✽5.�ú����f\���%�"�Z����E����%�aTO��~Q�y����3�@��[X6�>�W�Lu�w����r�"�C'y	:f9���ke��\�Z�f�(V��.�N�jp�Y����(�2 ���y<��+&���;��tB��v���KE1�}�Uc�Ӟ�U��ʆ��D�je���zu�=��3����T��E��4����OU-%���)~�0ȵu�<�.�׶6n]��x���K�&���c�d�<����z{x~�&Ki��_l���5c��Е�ͭsK�/ѭ�2����^��D�M)�*^�^��E��#�n�F���z�)�G�B��S�D����W$��"��7v���H{I���xd�S-��!�p6hy`�l�z|1G�O�O��5�I|�8:<�==�T�4e�#�0=�&�ƨ�x��݂�0����� Ӕ:�q�r���9�m�A� �)e��[Cw���x�r����e�c���A4t.𹉵��Fyk6��u4����i�g;m�R�\���A���ݡ�$��Z�%���ˢ�l*�J5#mQ�G=�F��z��{�,eK�r�{WT��lJm���7���2s��7큕��yp�	{����V��f��x���8��we�qS(/x��v �v�1<�mU��u������9��Q��S#;��@�^� r��Kbu<[(���Eė}�a-���CƩ9�!
wMs���m'6vU�v��U�6�Ae@Q y5��{�b&o��kw[�^@�H�Dx�F�*Ac�[dP	�%q��L�%!�B��a�������j~��3�������'�M�s�7@6�n��-Yݲ���u�Q�'{D�g�-konh=%׻���:���0�m��>Id(3��'ۑ̧�����Cn|O�6S�N7�f|�<�:�HLӋ�d[4�Hh0�����a��?d]�y�r;Ґ�>Y�[��1���[rT9^Y�ͮ�&k+x�5���*����6�^��Qz}�m��٧�cr��K+����Ar��@_(fNdR�L���6jv�z����N�g�(=�Я������V
����Q�U(�f��2��u�ofW��U�������$�e����9�j�mV��Eʐ�'>��u=��o�ȴ�y:
r��Q�q��"��{tx�ٴ�)���|ƚb�r�e�Ūp����oV	W4�nWf����H�Ŕ���$��nP�dّV���Y;!.����s��W�����MǿNx֜����9FEx��:�8Y����O�\T�]>'W?3E,����U<����Q-�^�4��}`�{�OP9Yu�jwTaXl����{ �6�kM��+������@���~ש��8���Wg�yZf��$�E�N�E�9�,��BM�%�Qc�+�H� 5�� kvFc�&����$�ٽ���b����힮��z��Y�п���q<I�B�L>�3�n(�	�#̋W��K/kR�A��6� ��*�,��^�.��C��[�����'�e�0<�c�c�,�gj����?�9:��?}S���{=V*��q�)>/�yc�r|�dvP*-Li��Y�^+{*��&��y��Ir�=��@��O�,�H�R�Z%B�kj��=�ֹ����=v�5Ɂ���#T����w�՝�m�}��L�t�d�)��a\>������{�M�>Y9̗3�	��]�+��i {�(�߮)�|uʾ �=G(�>܄j���m���
�@�뜑�6���'��(f��# o3	�P��tfP��ܻcQ)ŝOkL9(�ܜ�+]nD��q�[t�F��om�Q���/�v��S���(3��k��o�����P�鵣�Өv_l6s͉�ޖ�w�n��}��h	�О��V1y�C��7��9J�^f��R�i/m��J1�C�TG;�xFIh��&%�z��|v�;��Y�*qbu[�#v�o4�n�f�9I>�]�a36*b٠�S0�����Aצ���m,6s]�]̽*Yy�����>a��ӽ�.dV�D����lU�!�F(kw1�8�X��Nv{W�=�Y�k�u~cd�4�:�4H���@ݚ����(_!	����9 %0ֵ��/�9�i��)�-�v�_M�H�I^������ꕧE�9�nj�YMd�75wB������<"�s1G��u�s�}<�j@��*p���`��쎿EB� G=����f�6�SS�)�'��.u�wD�a8�ә��r�^�3K�^�S�4�a23uЯ��U+�ʭ2�( �yC�e��5��n����/=dw'.�R�Ժ1��d�Z�;�8Jq2���z�O�Q���,j��4��be�����O���S�*!@�:���{!{���E�$�_L��FFC��*�+��e���-��\H�v���Ǆz�b��VAEY���:�,��zy���{uש*��
��Gep��)��Pވ^.�Kýܓ�%6���S{?���.��Xu��:r��df����*kF��uI}�ٙ����c�Y|���z+NrDwq�2�)+�:om���b����k�8�ꭶ�;p��)J���]f�s���A��@�����֑���WD�H�ScW��Q�k�z�HY3ԟ���\�U���+"�5�6aE��<Iug�L�"�>���ˠ�GOV44��SmK���SS���(�����[���C:1�́�T� �n9Q�p$�@Q�^*��h�}�qKװ�yjz�.�K�ugk����O�m�[	�+P���D���<���^<	d\��3�=�Py�)w��ѡVe��!2P�ց���≬)	�-����f��3�Y$����6zHW��,Wl8��X��-hP�f��ȿ##�Zwl':��%	��*�ų@J)�:]>�R��flЭg^�EcO]U潡ڃ(�(��k�lč��3����[2�O��Is>��7{!����-�a�'wV�u�"Z�Ԕ��Y��}r���d��Q�nm�9՘��c�+�b~��x�C�3�؆�����]�w�fhuL�s$=��v8x�������_�at���ٚ�4:���:m��Ƨ��X4\��S�i���G�j���b�d���D��Usu���i��7p:|"�i�A�&ˎ���Z�c9��86�$`�s��p���C8I�}�a1S�V��{	�Ea�f�M�+b�����Hc��ⱳ���.^*�ԏU���&84I��u.Tf`독�RQ&��͈�-�;[�MwÑ��ૂe��Ƥ����pw+���W����nv�P�yN���꽤�>�-z�
��ۜ/�~����K�Y���ۊ����!r�u�ڜ�ו�Pz�FM���/���8���ͭ���up��:�ٷ�Se
���m��j&��uۮ��wC����r������_%�^>c�Q��["��'�;FC��t[���U��4J�����!�i�#�����C�"�`�|=^��?c
�5��]K�~��܁􇞂�xŵ�,��Ol㑀_c���6C������)��5�X�\toTk�]��v��`�;��Gd���a���nOp����l�A~�0ﭨ�U� Gjơ�g�9x�u���2v��W>W�Ae�^��`�7��	u��j$�$7P7:�~�'�J���^s�5��م)["��<M#�['z=��>�fY ���^����x����UG���-�<z�`6
��U�.��k�f��=�W��J�i�,�IH�����И-D�]0�D/\��%N�jU��J���AgR׆���כ]7O�6K\�l���d�I��=u�cS֐�їV>���I�1�=}RL83ig3��Ρ:��\�!�J��l?�"�޻��wrY����T� �E�WϕҺ�%:�o2�KrcjÑ4H6�U���r��;���CK�j4�0���꺹:���@�t}��
�u�x�!����˼`���gu�����������2�ҙ!�=F2_W���j�u1�i�ɴd�N{a��'�ѓ;��m��&~�3�9�T`�p+�t�����z���9���*�vx���6Fl��R'b���6��JjM� 9n�_��}�ېk��M�loMΞ�L_-��&J�;t�3Y7�ru�k&�uw)�4/�3'3�S	�(%�-:��ް�:pӦ޸m���u��=Ӻ�U����U�n*^����x�d쎧�dW���F�D&}��Ꜳ��9
������+7��ĒN��:@���9'FӖN�.�^�dxdK�솯?)�v��Kf�WcS�gi� �=+Os���������m�9��٘yQ"��Y5���W��`W�]�E���xF�e�W����v�w��֖�W�R�=�/����������y^�FY��mP�^���s�)�^��H~#˧����c�+և��[h5s#��<H^8eT;����l�t*u�h�ڰ�t�$=��gDc*�gB���U+����.��^��A���-��%���V�u���V+ml�Ry+����ASg!FJ{��(V�Z�[ӕ�Kq���3[҆<�
n�;�Ӽ�,�ə6 1���J�4��=#�]˳�����)t���1��e�U�M;A΃'01:ER�AO Yk� �:],�/eCs���u���U���Xjn� �<���'����eޫ=�Ξ��v��tC���]��U��.q����]�7�Vm���|��o6x��#$�W�SS�Ɩն1��a�DJX�Z�X�c(��Yd�����!��`ɂA{��l;����L�ԯ�S#��e�`A�:�(S�X���r�Q�cNZ9n�Y��]rl�-��C��B�Qh�҇M�z�i���]�+�p�L�	TX�m,��ݣ������g��k�U��я�˝|��@�=�v���dK���Ÿ;��	�R6�t˱C%�>��r6���tv�F��+���R���H�,���\��AQ�U�d	D�YYs��k;�cW����7uB��ʮ�	����qL����oL�M�n���Cm�De�8j�U�a<�±Q\�}.�}t\���ϕ(A�âe��Jo"�ް�=.����F������F��bPJܾ�.�qSP�V�*��Zf<]�m�o 2�����A�KC�مv��M4�A�p�:��|j�C��!RY�
��%�Lܜ�GSV(��޺��:a5.��ʘl�-f��l&�8�-�����#Hdǵ.��S�vɣ�ܬ�206� ���Km� ��S7�p�c�⏆��F�U't�u�c����]��P�=I{iT��GJ�F�dHr{4G��=�ue(��
��㆖�Un�Pj�*Rf�J�7q�k1�B�);�`���vȰ�Ӈ3�Rc:2Q�"U�Go�"�v`1�۲�B5�J��n�f2��s�䨙���Ҽ��Y����+@�w*���;�6�j���\[�=4t�pФ�*ܕ׷��.�꜑���e�q<G~�\7-�&��.�.hp���_`B&fu�&�����'0�i9.4oEg+t·c(؝�/VE�8������``̝�WIɜ�}ךʅ;7�+��)�r\��toXj�ـ  �_l�k����Y�R�Qk�S<Kׂ#bP�|y>�`U̫��c�/�z�R[���l��]��ܳ\&P/�7U�j#�Z�ei5z㼮��uP��xv!�8����)\\�2&�I���܏�9�� LB�4qT����G�����Y�v��Ѧ��5u)�kBCK��Nimm�l�iE��
���=�S��9/z=�9Q!Qpn4S�\.���Cwv�r�sއ$ڮ�k�����LCL9��Ѐ@��&-N|E	��n]Akv�nB�k)}|��Lp�K�([}�>�M�� ��#V��u��egYWW����p<����q#��u�<,^�$���\y1����5?�Or�@�M6�*��sD$��i�ڊ�$����Ci�*΄fp�m$�%��fD���4�Bt�,�����I6�E��j��B�i�)RP�Q �֗!M9�4�jQdt�8���i%�Z�V��O"8Rᖄf�L��UnT�R�ХQLꢉ�m�-l��D+�H*h��$���@��s��Uf�r�4���T�-5L�(ȺX����X�k3BʔC�"�h�)BZ$�S8"��Y�DZ�O9<���LL���EMJ��ER�!��d�D�*�XXUB[ER��D�b�C˜^:8J̢IH1D��D�J�쭮r.8�J�H���t�F��TӦEkD�NRI�+Q.i���.Uk���)�Lt�qQX�]�]�����v*;:�ibMbp�![u0\K�݉j�mV�r[Ʒ]8��5��gA�6���i�&�=��w���W�Z���g��=�+
�Q�<�(䀯dv"���X�/2q�@����n��^�<�'�0�'֯mLr4�։
�[P��m�{}Q8��z\x��kA�ǵS�@����騏A�� ��E��Z�Z_�{kchP�y�=��J�cF�j�Ms%E�;��]�*��/�Cᐦz��d�H�A����7E���0�|��<���\�����V�����w5>�^N�I��/l����f*T��S��.Oi��X�:�^��n�J[�O���Y]{���R�h�a9В�b�L͋��ҩLg����u�@:���_�s��r�}{��׻9��4��C���+a�Ur؇3�x�(y%ع�ڱ;S������ڳ;��c�m_�UM楇��
pz�*V��S�b���|R��i��HW�Bs"���%)���,�=����[y���f�%�L5p6�;��i�qNt�͔<���d7^������j���(��w[�h�4^��gZ}ʮ^�(��.�g�#�*��{cr7'��o�?�?~��ؽ��%�`qE�F�fM���1�lյ�g��o٫ܽ�F�8u	Z�(}��wQ�\���s;�Yhu<�n/k��wlL͔�v�����I՚�pu)o7��fUn��e0���{���u��Hڊ:��Ol��nKy(�C�)�×�U�7�Ɋ95�V�^]����%�MY�j�a��=�w F[���r'3��E����Z��{���K3%X����jN]8���^u�y�!�S�y������Pg����d��wQB��R͌]e�Cg���5�3G�z5�R9�!l��Օ�+:-ζZ�J�� &�/�n�'����jE�pN�(w��}	�y�ñ��ء1X�Ex�{��q�֣WGq�ȇZ��V1י>թW���I��x	��%J�o?utKD��)��k(�YŖ���qc�!U[۔��y����������g�(�)+��mNB˨�_��p�:~�,l�;�|=���|���V^݃gd+�g��(|��X6l�9�hQء�i��+֠j��uW0x��^q1B���:�z�ka2��ު�+a̗5��$x��yjb�c�J���)�ͅvo��n��2{��N��#i�-����4��E��捇=��)�Gr]U����z�DNn�Y �b�$~�mx�x��ց�;�S���Q��h�\b٣�E"YDew'�/msjh�=�ΤiQ�2���c55�φ_(0�����'�7�����]��L������,��Q��K���ga]��F�H�*a�w�<idz�3�뎖l�vSލK�*;�����R�$N��|��G��wz6t��HK����U�lb&8��mn�շӹ��^_�U=t:�TJ��>+-��%�#����Ŷ�%��t"so73&ާ=��7ICGl� y����s���d���Y���5BWxO�R7:�1A�� {f����tvmMn��1Ĥ=B���D�����};�h�>�޶8z�q�sO^���S�v�AlGa����(�O�IdKj��j�cL��7p:DT-=���_�.�_������c�ĳ��h�u�c>~�VMwBl\�5L�j�G*��zi�'�aU�]DP/˻��N9���$G
�t��id���,��Б�J�f׼�sL�{�|bRz3e)�j�y�c:{�:2�L��>��b)��;,��u��G#�d^G�;���j�b*}�'U�!^Tc�mOY�R��,I>��e_�f��@�l�z|3�H	#A��I�i�a��k�E��ݩf��'��0�j�b�e#UO�n�ЇWn�I�1k���e�ͽiH7���)��I��{�Ǹ��A���f��J��0�I�rgsP	r�:����*��:u��d<5��ҮAk�J��Uu��˷�Dp>9P�{�]��f`�\|t<������Ws��).+�u����Sw�Hr(�u��Uo ��1X��V'@LZ1�Zf��MLSk'%��(X��^gnj�Z�rZ7B�v��o4b֙+�nDHQҬ��+�(,���~�R6߮�=���@�d�7�Ygʯo���U���;ǝ�"��H��;�����7���
Ի\���,��������=��efL�-J��9�:BU���C1h�>T��^��W��J�i�,�IH|���;�Fh�6����s��3禂$��ީ!+��DĝZ��#���7h�%�}ݲ��������!�m>�ɚ٫'3X��ui�a�U�GN`w-�A�n�z��ǭ�dxVfL����ӳ{sYKw�^; ��I��.��s@�k�!R�s��d>6}�/�t��ڥ���Bz}果��vBh�eF��]�Er�d��ͅW��5��.]��N���9�oM��i-W	�Moλ.������ו�P���5���5�0;r��B�C2sJ3����jv�z����2�3e>ZhU��;Z�Ӱ�K��3j^���͕�J���5�0ߢw�����V~�}�L�l�w��G$"��͎���g�5������_5���z�m1������&��MA�5Pj~Sh�[HaPZ�s�Z�Ӷ5���z�h/�=Q�Ps7��o���}V{�����ɴ���m����Sq*��!�ų9�=�@݄;��"�l��9@M[r%��wKW&��N���Jy�����®�>���Z�W88`km��(T��}�k��x�-TNH�tB�����W1��&�K���:����ɭ2�]�D-v�<O���)1Qn�"�;e�/���lr=^�׆�Y_���4,���<4g��W����������d��-j��]���hnA�6KJ�ԟ,J�e�
u�m{��Z{j�e� s���������U+i�OT9�/6qv�n"uy�B�K��dC�K�:�X�m��.��O^��ˬE ��wF�Q��R����5Tm�L�1qOѼk��薉��Xk�\��ic�rB���I��U7�C[fEu���	f*��T��P@�T�$)@����C]?�_�
�P�Zڻ�Oi��͝w={r�U�/K�����o���J�EmޘqD���A�=0}$Y+�s!a[�Zdz��;Y�9�\���y�o��ٸ�d�jC�B�!�Ë�0�����>A�=�]#P�W�"p�"�-��/u�2k�c!��<���RcL�I=�/:�A����	-�=$��9wQt�'������2�k��p���o3��ol�2Q�U �&f�\b١*��G<�}f%i5-ƪ��c�KL;Y��7�4�^�zY �Z���/�8/���O{���r(��rث�)��DOݙ�Z�j����)~���^2
c����*X���ͳ/��̳0w��T�PU�Ej�}Q.�5�m@8�����,�U�6��^jS~`�<+�-��p�_�P�]2��%��%ث�C\�P�Zx�����z^j�Ow��,����WR��L+��5q�g۳R:���^�B����{�����޼a�"_s�H`^J���#�'E���ۦY��#�ɹ�\!��7>ۇֻ��];��Bwz�T;Y���Лq��xE���8������q�;�cʾ�a�e{�ӝmu�.�����(�f����ڶA�6m�wB��z�[4���j�a���n�x��,���VUi�}���	�����{x��8 ���"�:^#%�c�oӣ��}h^��ѝ��������?d��pi&����d�!�`�e�M��}ۼ������P��/5\�hY�nu�\���Mp(����R�Mz&tt�ȩ��.���v<#�ء1��QVR<�p���j���v�rd]��d+�H�t}��k���A�,]J�/��s�X�ޯ
#�z�׾R��6B�^UT�-��%��N�3�B�O�U�<`8I��~fv)*��quQ>�k�Y�����E���y���3�v_nuH�L����z��ד�|.�p�>FR��O\Vފ��q�ns��P�&#��o�^�R�}[�ӴY�ԥ�����Ob�[Ґ���c�Q�kj�3\�p;Y��޷�n��;;�*(r�Tan��^�I ����3��ʎ�~�Btߔ�A(����c��s��>��7�z�O���j����FY�$�*���c���,%�L�Z�l�S<�>�s�K3v��9��z����f�w�uy����Gi��h#�OqD��6����1O(��<�6�޸���o��e���z��&[�*�_��_���*:�~��i(�k���-��!+����ԇIn���K-��1��7d6�4:|Fa>ى܎�;�)�.D�r�䮝Nf�����;��V�^�A���PA(j,��Nz(��>��V��j�i�����0a�e�܌�C#����wm�t�̆�y	:f9:�E��.����jq�!�쎚�n�O���57�</ՀϒԈx4x+��j�腆��2/"�K'Ǡ�D�꫘k����cL�ɻ�ֶs��%!�&��l���yYEA�&̅��Ȭ������Л�Q �uJl�.ֽ��w�[�ޫVC����5��W��8�q�d�DY�8���x6����Y��z:�@��.����*��])^d�����_��A:OwI���԰�fF%Z�Ӡ��8a��
͕]���7�6�bkV��=�v��˟Sͷ�g�i�^���֫��fJ��s�X��s��ghlO�	x�6�.�$�#Ð�]K�}s�uj{����㫧XXG�.���%�Q|�H����퓧ne��3�_�>��✏)�;,p5��K����S�x�S�*�U2zխ���%��ӚD���^�D�pe��g�3�n)�eX١�]�,�p�� �TL���ݦiTַc�Y^�<���Q��������f�*X�R=�UO�~�T�����E��^�=H2�2�1���t�זAe���,5�q��\��	; ���V��9.��5��}���ޜ*�yR�>��Vis�ϔ�,2�;\��e2�4O@�fl׽�0�{���g�ݤ�!����P��>϶�Yiu��S�hs���l$��ϕ�vۯU�1һc|��+=ӡ%mO7��Ae#��ͯ��F1��Nxi~�>����u�r{�\m;�5���E�)8�V^ffKɺL�J>��b���H��a a�dTJ�f�
�oYi+a�b�?GDĳ@I:���{w��sP�5���L�ZT�<�.�ƻ��|�c�.ݴ�̖�E��i�V'b�^q2�c/vl˴���H�f����	�۳�%��a����_V��Bݱ~3D�̨���s #\�]\�i.���o�^𗧨��MR�����dv�w;��.���du2�96�T4�ŕ��G6�n�K9���=ך�g�b=d�WA����8�zF�͘��Z��n>��i�gu�5�1J&�w.u�j5}2f�����4�p�5H�+UBm��.f�C2y	J���}�ېk�>%T���S�TH}Ħ�Tq�]y��+�Ў��"YXj��Ș��g_(fNd
S	�(%0Ѿ��.����u豂i�l�!��>�x��Ьl�눬�6�^��4�֮K�VEw!�Q	�T��Y"*#d��ӬQ�~��3|k�����T6t;��:.��'WK���#�%��@�c����&#�S�}�;v�V���Q-�C�jj#3������"��Mi�r���`n�,���N��2�՚�� ޥlr��(ּ4�֟]�jM� ��,za�W��^�߳�tn��e�r�uM��3<P������W���9NW�26��t�̿�8�X�}��=ۼ�eP^�Ϡ�nFGdG7Sb�F�9E]yd�Z��6�EηPc$��̞�Kq���Mw7i?;d�f@6("�q"F��熌�+-r�a��Q���xtF.��\v#��3I]�CC( Y����k�b��[f��)Q�)ֱ�7޶���}�Ygm��|��&�/h�7��ڗ��QG�Ns<���&E��^��k�aV��L[y�6��z��3�j���;�L����l��Ï�%���n�6�v���nc��P���9zb�n��KDXur�-�2N]Ob��cd۽�FPj��ͭ�GM�3�Cۨ�Gg�\�@�F@��-�+�W�^#,+�z�@�j9��h,�9/����]��'���iF�2�H|2!J����K�ٱ�ꌃ>��U�'���������]��BewmƔ�O5y:�%W�{dL�%�.�Py���\��>8�<
x/q��W��u+����ѨV�r3������ $�X��flU�-��Lds�w֮�.Υ9�T.�毶+�
�OM��瑨67���W!W.�s\y�.vk�8�5���@F�B�W9y�/ͥ�Ǆ}#K�NqR�迩�xU�m>)U���g��!9�ڧ�|h��3cE<��H�$'� ߢ�p�GL���\2a�Z��N�gI�ͤ=y�x&s#����\a�w;jL��]�؞�<"�V�Y)�z60�n؅��vGO��a��7ʣ����嗠�%�Az ���ldD���=έ>�xk±dkO�U�5�j���,��j1��+Y�ӳ��<��m�2qn�,���'�6� �ZՑq+ԼF}.�NC~�>��B�ζ�Ϯp�6���p��ڡWn#J9�ؠ�5)_DN7���J/S	�no�G�[?.�"0t��$^J�Y3����XRQ�����v�aL9Zh��d�T���WQ�n�t�R��j�vd�h��7����v�$�:j�7ݝ֙�Ey��hl��x���q�*�9XE<vގ��d��y��,����;�(dJ����$��P��.n���hsB�N)��+n�eJ]	����9甋�*k��[ڠ�y��ǂ�C��;w��}\�.-H�%�.����5V�V��u�����޼��3V6V}�v�rUɾx�f�&�Lv��ض���јsN��[2b��
��f� ��Ҋ���P�YN�� ��4�|�w[[�0�ʰ1�5F����xT�-�^mLˇ.��� ��ߥeخ��ۇ�)�'{FX+����gێ��m�8�\��5f'RpC8�#u�e�z��؃���:m>0�eܝ��n�H��7Yr�#2�ķ�4{�7���S�,�W�q�L��q�JD��_v�[R�\K�u�������ksu���|�&�L����X�\�ڶ�&��.e�"�ts���:��[lt�6`�|ކw�J�p��4�j��>��=Le��؞t�~�r�0�VNŎX���n�t ��i���^e3p���� �Opn�J։j���P�;`7�n
.�����]Y��|�dݷ���%L-}\4�)rqVe�KXL	�k~�e��;�u*T+k�P�Sw����e�tc�؊t�DT�Q�����P;AM�B�j�^�b_
\@WV����\v�}z��p�˫̢���aM�Q�f��s]_A���͗����T����v���M���Ǐ���o�h����q-���У����&T;S�����.�Q.��O��ڦ�hW�����ŚnM����9���Bn`��H ��p		�B�o�+�nBb1 �ͅ�z��'C��Е��ʺ&�HE�/c�]+�Ȩ#(3�e��Q;�46̩-i��^:{��-����[��S#���7��h�;���ZEfc�n�z�65�يXmv4$u��*�U����������lu���-����M��t���ث�9�#���o#� �]К�4�:u)�ow����+���F̵[Lnk�P�p��GH�Y�R��n>o1�#x�6��)7ٻpLF�'��<Y��%�ڸ6�d�O	����**�ȴv}���8JQm�8`w�����f�r�`�<�9jm��X���R�-���.�I�ݔr.�t�6��R�V�H#z[B��9�d�-&�
���N_��.8��M'�N��U�ՋW8��B�/J:#����t2��!�8��D�v�ͻ>�wY�jv������bU����+��#I߱i!\#Yb]���V�,3�����4�R���q��[�{mr@�KH�Fa�L���k[,2��z9v��M<x���s��Ԋ��ie�.I�2�6>p�^R�K+gj!V�����J���	B̚f(D�Z�"�%�$D���-$��-%"�$4i��ʒ,3U�)��jhq-�9R��fH��D�T\.�\���CH�h��H�������D��(�UT�b+JQIjE&�
�NlA!��Բ33"LZR*�I&�H�s�`��CMT��"�$:&�V�dQ�Q����Bl�DY����VR������"�E��A#VB%�j�)VʴLj���R+"�QD��Q#(K,��4��!T��)Q�J�r%LC.$R���aX�Yi��,��4�,Vf��aȑC	Yj�'N��S(�(���EBF�D�E�͐d��EM1*:T�ra$����P"��.�Xi-R,�2!Z�(�4��h�"��>�(i�jX�9��͗���=7L���b5��)��꾣�dL��A�e�R����oZ��\�Χm�n�v��z����v��������7���^7G�7g��tBN�*.T�G�B���+�_�ڜ5��Y3��!�ԝ���]DL���3��S>N'����=��6(Ld,���A'�w;o�r}�p���vOr8]�>�F�ei����Q���>E��T��O�����S�W��Lss>m��v��`�7�J;�K�,�x�B���q�N�/����⟸�Ɉ�����%���nt��n�+wY�KC/tf͵.�\v��6vB��{2�!W�\����`�������*���^�b��s�^k�5�3
X�DJ���\�NZQ��ʵ�"�3Ϲ���Y�S�ɸ�7o���>�>��>CÏ�u`2�p����#�ZH�{�'{���RS��E"�Y�w�ޣsUy��v̂�6�A�,w�Z*��]a~FGf��ݲ�ϒu��A;�%XfՀ�i7���Z���/��u�$_�T�S1�aV
�=�B�Ҵծ���/Q�~Wr`(�X�U�j[J��f^�܊�\�n��A#ء��@/�rZ\vO��{n)�����:��6jj��z1�z�E?yu���:T��'���jL|�E�Q=�1�k�om�2g ��ִ�vg�v�&��up�qa�5l*��A.!�����и��3c��@U��A�!ϵER�;�w�{r�0��fV�N��n����7��-M�*�]�t���w��jD_�C�N�E��KςN��N�g�v6:'a��d�{�:aEٞh&�c�g%��^V�f�6o��)��VMJn�uf�;quJ%���	dKN�����:&�1�Zk�J����E'��݋��lb3Y6gq��d즧�d��؍Q �]t���A��n������'�����T�Χ}� {e"*"̀���j<it���Qf�?(�u*���/u����t�L%G�Ϣ9��J^��.��1�KG_�~f��?r��Q��o�z׏�����&#��f����ic*ê7d^W���$,��$��/�Q�3ŉ'��E9���C�ͅt����s5��kR@O��:P�}�S�Y�C�9�a�L���<I�0�k�*������LIt{V��׺�_���!���B=!��������,�%<���n��<c�u��ҡAK�l����w����  �arq���GJ�@.r��,2�;\�S)�1�x̆ޕ�L'����)�n}'��s8��U��t��	�n��h�I͝�j]�r_,E����[arZ��V&Vb���L(��m�Qۇ�v�5S#ێ�0�'I:�?��"48a�۸�2
����D�+orm�>SV�A�e>�ggNͨIYʳx�o���{��ȩX�|U���TJ��y����pX�pyk����{ivuj�T�.�s�p�dN��߾s �AU}2�7\��P��h�>T��^��dzw����@�R ��x�F��w[�*��}�$)��#��Y� p^SAE9��
|�VF��Z���*�c#.�e㡭�N�ON�����Е)#��:In�r�?d(3�޶���"z����"=#��}U!wt"U]3b�2-�9
��6c��v�2U@���1�e�Thm���ך]�a����9tK��r�d�l*����>�.]�����&&�1���U�>y�ϏN]*�7^��x������g���(t�xSEJ越{[9}'U��fkJ��L��e���������鿳ex�u���K�VE܄b3�h9
������Vf,��*�	�D~W�~7�����go��T��r���S���������#��~���/��ou�6�e���h�ٴ1Ni-U�a��ɻ�\uC:��")���a��~��]��j��Bw��Q.�w��	��Rcp���׆�Y��]�a����eA��j��]��&j�G\�d��Tϥ���!C/
���0�fT�:��ۻ1�zUI8JL� J���Z��Pq����[���z��(u��CC�צ���/q*�ҧa�*��I]������$"�H��sn-�����&sC�;{�)Z�����e��H/kcf%�L��9����Vu�?m�?	�C]Kg����c��^�<:�B�ʑ�o��73mJ"p��f��t����/���dvDsu ءQXJ*��9k��m��n|��"�պ�۫r�]i.�:bOC�38�L;�8��x��薉��Xik�{yc�p�]�꘧�����׏����Mo���8 r���& )@�7(\,�~9��!W����U[6lw=��*"��n�:�+u͝V�=`�]�>%��A��d �_B2��ﮒ���^;;ط�4�p�Λ�2=7��|�uZ��dB�!狞1��v�g��W����C�����i��;��t����h�4����I�i*�{dL�%�!�*>�t�\����5,]eHmn�.�i����kE��lT��q7�7���@���NRO�Rg�f�\b٠�S�mfV��=�I�v�am;� ��>8����h�C�n�n?a��rr�2+��.RN�iӽ�Ŕv#��n��'��t�#�a5e������i�t��*����#vjGV��3jB�X�������	�툲|V�x尯%�g%!�%L�d�t�V��ΪS#k�5�Yw��շV�����nm�W��>=�8ƺJ�v�Ah�&����J� =���1Pxv��|�s�J����:�fd���L����p,�G;�l�:F�����`+r�]9!)��[���D��Upz���t��2�>�ymx�^�Tr���(�}i�@����}���6'�O�ڋhl	U�٬(���p�<Ӻa�e{�,_B��Y�S}�;��p<���f�&��1�QL{�_>��%�N+��6�k8N`0����O=��|�O��ꙿ���� -j��^����Wc�r�m�.�֑k���k9+���q3������&ۓ�р�0�4���6�6��f��Ѩ���ޅ�/#=S3�n}v���{��J��Ԫy��N�J����P&x9'�bY	��>+ý	��dU���E�+�Ż�b}�e��E.�����nZe��A�2��|�*��>Nz:�W��� 4�P�j9�����b���cls] �
9!.����|c�.K4�U`O�
D�>�ȕ�p&��,�����y=ךZ�xCg+�B�Sl��qŎh�W�fBR�*.Q�Šr�0�>���ހ���UN/b襹ܫ�f^)�EyL�-�	�ζ�s�-9az��}��>�b[�.w�Ǖ����\�ٰ��
xlp��G�)���<%[7w�Bs�SC43�R��7w35�͒�;���<ZΤ�W#�)m�v_%���u�|lS_<]#Y�\��m���\�iJJ�v��]֝4�9:�XOp����qmb�˶�+��!FK[��W����b"ծ��P�+]�����	��B2Z��\^d#P�|���~��z^�l'ȶ)(�hԮa������S�Hϟ�'����OI�P��~�mu���g��e9H�%Ē��.^U�<K�}�^����)���.�s����M��gGh��Ga�7TAtn�UFL�M/o�I���i��K7d����بq�b �E��_�䆗���nm�9՘���=�'��&Z�.�em}Q��˔˴�(d�>I�1�����Q�]j�O:��aHkڻx(J9zUS�Q�{�5d�n���ee��ƑY5)��!a����xd��Ȗ�j��k�tM�E!c���o�5�NU�u-<W������l���5����PЛ�Q ���:-��ͩy���{j�l^Ƕ6nC�� ��ON�m����jk�*~x�Y���E��;.�yU;��ǲԻm(�������N�O���yA-t��`���?r���p+n�]5 g{���+j��X�.:�SG�ȼJ/��vK�4N�i�1|<$�#,�{ޮ��j	��� K`�ΗM�N���-��������7�*�Ϩ�m����t�%_U�f����7��eMc��NE�X�&�`�Й]�:Ф��Jx�S[�m\�X�����民]��=Y:cۧ��k8:p�9�B�$uE�����{����[E^m�T��͙:Ť,e	�'�s�
5��=i;n��8I��#�9�l[���Uj���^l��(D=��S6C_t����#k��Jy����.x�<IO�e9�8��flw��H�P<uTeє��S,&]���.���Z�����W��r9L�Z-cL:f�ao@�d��	{�o)�>� tԞbu�z[+�Kv��["$(S�x�Gl�I͝-]�a����y�ms�/�!z+���$v�T���`�1�P�R:���]�2����js��]�:�+��ɔ���S2�4����-�4��4.)�x�#���;��S��)���D�����̊�(�w�OR0,4%JC����k�n��$���Ό���5s��ecݬ��uwoTkl��%�O-�v��D��f�\d[4$�!�l�9�]��U��L��0'x��׍�{^�=��E\��;��5{�D��+�3'J5������F܂z�Ͻx�u��&�=�Ku)��������[���O��������;���P̜ϩL&|\��^[l��#���C��Ś��U�ɇd�:����=�f�С3��L���,b�E�I�Qc.�;D�	���Cy�y���q}..K�Ӽ����:Ҏ�"J�/F��Z��qL��OV�����l�(��"�v�z���w&�v2N�G��N��?�~�R2e��Q�9,+�l�s	�a�ɳ>�}F}Y;#�TC�ɢ�:�NV[���$�\yq�2������7�NxΜ���go��P���*r���S�������;�&��eF�xx�mr�yd�����:��^h�9�M���5�ɻ�@�<��g��϶�4]�M�CX~�:�*=�� ��~ש����Ho�����>�G,�)\��|Z��R����֩W��ꑿ��+��A��[=�>�KN�hx,��m�meH�Y|a�]Q99\+!�^�)$�NsP5���x6�Ȏn��
�,r������+μ�̘�5|��OF���K�W+�7��<�O��tÒR�u>��D:薎΅g|��=�Ga=yB�EOW)%k���j�8��`�N��,	��P��3�O���B��k��қ�Oz�5��id�:V���6vB�!�Dz�x.K5�*� zd �Y�_b�1��k�x��#�/����G��ؤ���-(�&|��aJ��8��K �8d}oP�x����4H���ZD/ڣU㦽f��+��-�<k�ӴN����B�2K����VGs��6�&�jL��X�r�l�rg92�<�w��aN�����tS!�9�#:��6��vЀ5�D��o����o��y9#�:�$M�V�jp�;�X���������<j|���~v��J�^�)(�i�Py�t��w$��od�:ɜ����%��rAnU��<]��dos@���Ne%�R0��q��9���{�Y7�)�ܐ=�S-���i�zh�-�D?#pgq�����r�L��>��f�	����M�s�i��k��������o͒����i��Mo�svjGS���*a)s8�nJ�! �D'2):rR�k��l�7U��<�*�_�8=5�/��	�F�u�Ć�w���J��g^�eMk�\�6�yt,�W�д���jq���U���MU��[ 3Ց�S/�rhf�r�EƼ��ו�W�^�܅���=7�)���б?^���4,�i�W0�^�nڥ-�\g5�N暬Z�Gl�EDY�8�� ���d\�R��1�����[X�xpB�]|y�*̒���f�ƗTb�?7���z�����g0o*L�S�L�w�+h��3UE(��{[��y�s���Z�J��aT	�I�Br�ϊ�r��o����\e�蕛���k��-kZw(��H�����]F����\����]X�S�p�b`���)�C-��u�'Jy���5�bMj�����Gk3��'R��ڻ�a{ؔ�[[\^,,N�6IǸԷ6�{��kK���sf��Lrp�xޟ|���W�ǖAu��+L�\H=�e�Zy�C�kLC��e��y,sE]��շ��T�!ۓ��Ak(� ���H]�9��E��<ITe�1 �H=5�Y�z��q�y��}Se{f =�R����Sb��V����5�̄�HTK�c���p3�1n�U3�x��w���tx�C4O�TV�L�-�-�j�NXJ5��
�;d�
g���z�����e�Rհ��y���Y���%��(�2ǰ��q�wݚ�2{��N��#a>E����q޴z]o�ʿܑ=�����d�᪤�SpzH���B���ѹ�~6�
�������Sjv+pC���}�W$�C]��ų$�k.���q�5�?Oxи�J�V����
�z��lg���i2�b�f\�]�K�E����zE�2˓�.a�������Մ��#Om�����fWf����fi�P�e�k�2w���c��T"�!N�p�sCS�ʚkס%u���'ݬ�pE!
�M�Z_g����:���n��u�G�ߞ��%�-#U\�^{�]qw�ب��g��h|�j'�9�K��N5�)uI�3f�΋J�{�<��I�x�V�T���R����F�=���	X�5�g$��n9[XԖ�&��iFf������b4�G�_�@p:xE3�r�.��:N��f[���Bs��p$�;TT���7Kn��z�]	3VǼ�@(u��q�΁��.k*�$����Z�7���ެ� �,3fr�_��$켈�ū 
�����O5�	��:�u�Q��e����7���rWA�ʽ�F#���fr�יr�jIe&���)d��&s��I}װ�4��AX���q8ְ֩`SOm�2)PH��wtу�P�is5�,)Jnɓ�e���:���[�f��fJ�S_��L雑�ݎ��ܮ���;�u3���Rñ�O���	�n���f��8�5"{ul���3+�JH��-.;C66P��e�Ze�]���AtcO:�����\�Jn7��Woh��r#��ٹ�z%�9Z �t����FÆ�4�����1.���XN6S�l]�(�E����Y|���	��������;���j���-�$�++���}*���%��:T�o��PP7P�I3F���~{����;�s�����]m�3E3Ң��p�g����̫L5�`�\�\*�<���[{��X]��YVs6��]�֨�	f�Y;�^˥����ՌV49.�X�`[/_l�jcemϝe��*�*�
��"�d0ԋ��B��Y:W���(2.۬���C,�DL��>�|S6Mh����l�ubr�g�LlZ����;��J%5{}���ŷP�Y��m.e𲔗�aA3�d���+�4궰�1@mǇ8����2oM|7�7f�����j�'��+J���sWٶ��w���x��X�{O#�-eo@�/)���o)!�Rʇp��6�KR��}�7@T���Pǻ���α�f�V.�0EٌY	LU�W�j�v`EPK�{,ᙵ'eK�ڼ���/z��T��$�u�܏~3�_C�u�{y�q�ee �EE!īYjۣ�5��g��D��=t�����X�U��.L��PoZO:ێ2+6�خb�ஏ��4��V�ȃ���s}��fb���`�Àb��k���!�wW��R��Q�Ro�o3
�[�P�d��C�am�1�Η�UG�!�#h�	3i�H� ���4'��Cj��Ʊ��
��\��:��ŐZj�nA�/�QeIt��d/�,f[o��bZ|0�Q���uU�6�zz+Y�̢�։G��H�ű���YJ`qs��Wt��P�ya���E���f�.��(i�OW<p��
���׿dX��aݪ�sm^I�@j��r����S�pKK+��L qQ���oV�{n�d��Nk�\���P�cJ�uq���L̻cV�_r�ky�wd-Lؔ�ٴ��}0�)k���$P�E P��(��BCDM�,�"�P��5$*H�-BҢ�3-*�hGZ�hW1LXuJ���B�H�UA�YF�!Q0���)X������UZJ�sRT�!!]ZFHR��D�.i�.fI��dZU�"i��9I"�dV)!iT�T����VeUG6�K$���9Y��DF�
,��X\�%�Iji�R$����(�4�E�Pr$�ZtȪ�QZȥ�(*�Qʄ�0��EJXl��d�9R�
�(:�R(�C��R��Z
��QsVQA�r�(��FHr������MHMR$�(�(�T\#��� �UQ�W"��QUb!��岨�*.W(�DDJ4&*�T%r��"��	j\�"��5�J�ʕd�#Vs0�*9&\"�(�Q(�$b\�(��R��Y�@
&��ğ�P�y�c�a&�Gq�(��{M^�#�Ftn㠆�l�Ms���{�9�ݸⶮ�r-t�d'���*;U5����w6�c��~�{�,j7v����7E�:mt�εi�?D+&�t&�hQ ��Y:���<L�{;:�j@��{�V�܇:�����Om�"�0�D�o��ml�@?<j,/�pz��rm9ܜ��W�/��q�Χ��H֌�FO��:;i���t����Z6���n�K��u�gv4��@ɸ�<�B�G�ȼJ/��vK�I�R�2�T@3ŋ��#�jn���M����k_4�^nxkT�S��P��~G:h�q涥��<I�a��������A躴_��9�V��{�"!�tð�k�5,gH�ydY!)�Xk��[������n;��4��/�n�]9&��(0_���ڍ��#��Y��W>,r�ΫU#L���4>�y�ҟry��p�_z@��	��
�z[+U��D;��N������	�m@k���[���7r6��~3ndiAQ z���o�e�o� �����/�5��g�_lQdq�������ҙ�a�s��T�Չ ��yM�����W}u}�1>�$��%j�w���#���`l��E�B&�y������ؿs��J�4����=�k�x�$�{/��Ū-����M�s#�ɅA��aH�$$j��vD�Y�J�[�Х;o�u�Z��p��qNT�l����g	&�&���F�պ�H����W�Ǌ�(�N����0,4y*Rx�s�r�4[�H�~F���_���so��L+�r��B��R;zK&�[2�#����|����P2>WNOs�$[��A���]6/�&�6U��@P!�b�r5*�v�W)��D��\��<��3aT8�5���:�/ӕ����m]GzA��'��8݆M�6ȅfD��ׯ��D���S<s_�I����n�ͨ�]㼐�x';�Cd\����,�ށ���O�mK�t�l��Uf�;�M]����&�&iW=J����'Y�o��%~�[���ߧ<gN3������·'$����X�.���s��Z
�e�jѪ�S�Go�J%�qE�-U�a�6MܗPδ�E�7A���u���]��bJ��3d���ͷѬX��<�B�G�B�k�^K#Z|���9g	KBq����7xw��ԏ��U=3�^��T<|5�OyϜE���Ȋ����������t��x���j�ջ�8��	tI��qc��Zr�3�Ȏn��
��QWAd�Z�m^D�7�G�{Q���(�F�|�J��0:�(�%�S:k�&,��9�Nʲ�i��W���N4�S��+z<�����r�OH�ER��&%Z��r���^>�d���f���'7k���Q��Ґ��j�M��
��=��W���;�Y��M��o���|΂N���tR�u>��C�V*�;���{nF���
��%�2o�t�z�����珐65�*2��
P4��2]?�^��Q{�u�H�v!��kj]�{M��͝V�=`�3�u4�f�A�A�= �@~�5B�A�R��ת�N���y��X�[Z����A=��J7	��H|3�R�<�s�=��v�uŶL����E��؉��d͌�o0W��u����-�#�t�PN�IT��"d$��:�A�>�܊��2����v�aeL�I�}��&%uz��|v�����LTd�l�2��b�#	��SBO�ٌ�b �F����K��'�Cy~��ڙ@Ѱ�4�h�~F���~�;��*��.h���|�wl��7�hv�+�\����lK���!�r�N�^c����k��ߣ�E�f>>���n��R�#�ޛ��xj[�8E_!	̊N�J�����g
'`58햸��*�7��d�,ƹ-��^�g4�'�(M��ɳ�P�|��=ZxE���Ɩ����XQ7r���/�P^�C<Ga���p��*j�JS��]C�ҍ*�"dak��WV4rU���㧔�X�Z��u���t53*�a�G�n5��t�Ϯ����a+/1mr��0�F�"��!�����̛B:-�],�}һi�s���!�}�ՅC����NI�|k�VH�gО���Jfh�[)����V�{��1�f���������׵F��ZՆb�kb��ed�1%�=;ٸ)�����"�W�x��u�r!�W�\���F���:]���z#����.p�k���/�5Ӿ���ɷA�C_C
I���]J����w���ʵ�_+JÌ����C�c�u�P�RIU2¨<�L�L\S���>��s�?\�f�;�Q:OR���gT�nA��k�?#���-ϋ�FᕦY�������>E���R�bB�L.����D�Nh�[��Gyl���D�H�Δ��Y?5+s���Z�h�A���$� _��f�ń���+&�]9��SXH�9��WU�V���G)�]n���l��z8��
�K�\;b�Bm�.�5�:`�(����3@8���0;L�-�	�ζ�{��-(��}��c�ᬉ�+tk�w��^�>�̝�� %5���p7��Ȅj=��/;���w�)Zb��W�F�s�/�ժ����U�6��̒�*����"b%�����_�e��BcV��`������E�^���csR�����TW��[:v��������3��B�������38:Zj���[XQлjk�]�`��g�6�R��z�Rm��Z�[)�����G�%p���c��Q�;�<�z^��5�ڃw�ӯ�e��R��v��ˤo�I�i�h��֓Ɠ��U1l��D���s�\X=�C~�J�Y/��!�}�eo�"Zvso��z(,�-�lC��ܤ��Pk[�����F��G`*Hǫ�x��f���nvr���Wڔ�/1,��f��"[�yD;N�;��3�T"���v1��V�U�,�B�ZUWK|���'��1�vf
���'�k&���tB�B�C"�J%���K"Z��U������+&���j^��ne�A���T-2 ��f}����N�j��B�k�Л[����2�E�b͌����u�)T\�LhՃ�d�t;���tW�F�����ܔ��e��~��k��{�������8�����{��呭�2�/t��M~����򛞩��H���lN/.�����ޝE1�
9�["�(�#B��}5�4N����͗���<��%<����|�����B>��C� k��|&�����Yms��;j�6s<5���U�~��"��g��{��y���a��]	���6��+J5��4�\y�Vn���sT�p�3�{�.$ j�]�xS\�IF5M��w�{'J¸R�v����6_k+S��4'2���;��X�9N�mcj�C c�=��2���G]�;Z8@��+w�����7���\����魵V�n�q=��7soU+R5%���著Ğ�1�S�2ٿ�e�<{qN]{�W>R�,��䍢���K���m�i}R�}w��8Kd�H`t�|=-���N���"T)�*�k��C6q�ܱ���v�`Օ��6uZ�jt������qU2�u��@/��FZ"��h���,�t-�)^i0��tl�I�%q��L����S2�4�w<`l9n����M��ou�u�k����9������!ݲ���N�J4��z�F���z�m����2CYʨ�*fpH�>��zz����c�>u�dy�֮�=CN���2��Ή\��lT8ȶhI�C����n쮫Z�s�/��3p{**"_V�)�r;��r��<9�\��<��0��1Gw�V���\��(���J6�{����6��"]���V��g��ˇ�߮���d�l/m���j�9�Q����Й��va3�P�S�;��Q��O���·VW���/I�q�+ű+��g����k�#�h+�"��1���9���~�}��~��9�;;s?��:��'�LxE�b����];ܞ��Oe�PvP��yY\�*�(�r�	�N�o����u�N�N���]<��ot��k��H��l݊���"E�U|���{&�9%�X�V��Au��yFS�����;�,u,���ٽ�D�-3���]k�jpcmX��U>K�GUx�5BSk*7soY�%�}\E�CΩ�~Sh��(�͡�sH�5�8�7rfP��n���z�{ �ή�2�˕yѡ�sL�)�����@�����;�(�y��U�	dkHY�/�cZP��l����G��C�N���.��S�F��Xڡ�\��g����c�+և�>�&O�{Fm&BV�R��CU̍��<I�Y"�\v.�ȃ����vDsu6(Th,r��:��2+�&���a|��Ͷ�[��]^Ӕ�@�.��$�D�<�EL�1'ҙv�^Fߖ'|eb�:�I T�c�=��9G%^��'�EScƜ9W�e�1J�7('�'��_l�mY��ż�ז}
�1W����"�_i�-sgeZ��>�x�O��͛ �2{���l���WY��f@��~�]6ϻ�kR��̍d&��Q�L�Z��dB�!�qs�e�F�5�u�̗N�]|���}@BKU�n���	��ϖ�}ܺy�O���E�2Q��6#&c�;N%o-I	�q>�L���%#g��u��ȃ�n3 r:o4���BJ5��Q�Q�����aq��T�&�aL���ޛ�Ƒ�^�S��S�SR�
� �Z9��U΄&�Ep+/��GN^q+Zn.7l|�q����5�l뙕w+�Rv<�S�b��r`=�S	���lY�z�Du4t�O��Ә�̻Rsq������u� ^�3�N�6��2���#g^� ~ȶ�������27U�SC9��]��ۙOt��k�\ʇ)c��BJw���w�i�eH��h������Ok~ݷDt��|�K�Ĕ�n��u	����B��9>Ja�k�/�J��\�Ӽ�U��\�GFo_�E�<�9웑W�Ed�2j�P�N֟�i�ڵ8�ҕ\��
&�+�afz����j����B8�9����k���<��6�SS�)�5��X��TKf��,�l�{�{w7-Aܾ�嘓���:N홏a�>U�*���_�V6���d_ҽK�d��}4㏖���{}����I��~~�b��:�*���o�L� ����R2#�v}\t>y]�.����j����mq�^����W��Y^�9�S�I����G����[�啣�����7��&����pyy�#XϖAEY�$�������ei�k���`"ǫٱS��S�kF;��:zʼ��V�!�q�*Q-�إ62�O�\�
9>K�,��Z\��J�ɉW	�ˍ�W�OY:MM^��`��~���i�8��_{�'�;�>�c�Y�K�N��P����+R��C�t�ǣ�^����!���F-#��ٲ�մ�:�6k��\��M���u�u$��gZz�f��3���m��Չc�H�܎�
	�?Q����R�lP�Oף<�����\{i	�!)Ry{������-3�73:�5�+�[Ɔr�3G�>��^���b� ([Z�i֛I�5oŏ[H�\Nk�,5��ސ��z&�S%� �b	2[����j/�����[g��cWK=D��U����m\-��t�����>���̒�*����"c�~�*�ᶺ_��Q�ʎ[z����ךL2���PI֒�'{D���h	E"[��g%^��:�忋ߖJqk�O6/.���etaj��!j��G-�r$wr��@��6.g1;Ifݗ�8 ��J�n�X|�f�ST0�]�k��K&ڡ?Y�p�'vf��yD;mr�N�t�ruP�21�c2(���m����{�9:�nq�,�dd�ػ2 �+*�y��²jy��՝�Pȼ҉d��Z(1�5�UZ8��/u�+k٨��Ή�i�L��>���D�t�/�Fu���u^�_gHS�yO&�fKVV��*mÚ��]t�G*��zi��z�����*#��N�����u�c�_�c��N{͕�g���kI�֬�yᢣ���7�?!�ԝ{*rU��H�>q��OMa7v�J�������n塐�P��̩bѹ�[�d�l�,���
W�U�=��IN��GJrł�ۼc7�5.Jɏ����P��tqW1>ɡz��K���nj~Qh�r3kT�����ٹ�c �*}GC�S�eO{ڄ�;�,��N�y�K^�h�S��7
9�B����+;%��I;�y���x�Qu�����U��e���:���Zf1������.W��O�ez��ȇ5��W2��ʜ��3�rG�I���FTkO�ߴ��m��T��+b����,�R�e���|�{���
��m�vT��Ŏ$��0�O�ʡ�b���uȉ*��W>_
��n�.��X���k��ݝ�E�J�vC��S)� Ɖ�� r���-��,�^UP슶�r#�FIX�w\���w�+����[둷^�fn�,�(#�$Xn��_���3�*/rC{?[�^�?t�3v9�:��9=�(��p$�>HS3�B��f�IX�+ݷ�B�V�C��sG��hz��;���������x0���eM"y3��R����?�SKS�H�O5w�`�/<��-b]�������R٫���r��N���%L����T`�>�1����`�6��`�6����[1������l���;m������?�l�����co���m��1��P�1����ckc1����m��6cm�`�6��1��P�1������6cm�6cm���e5�fx�`1� ?�s2}p#ݷ���*UR��J( JBD@HJ��UU*�BETQ*��P�$��R�� �T�T�RQETT�D%TJ��BT! �B�T]�Zյ5QT�U(�޺�B���UT $"U��͈P�i����cTR�W҆���$W�����H�ʉ�P
��!"�M�J�fKLH#LQU���H�H�IP�M �UA
�E����j��H5`
��飙�(�]�� �_{�n��]� �h�Қ�+Pu����͕l�+���A���p�u�u@黮�\v�4T	�vUQ}��5E(IQ6�O� k�}c]Ws�����]'O��ҕS�Nݯ� ��E�'Q@���;��R��E�ǼEh�E���|Q��EQ�R�:4h��:4n��Ѣ�(��Ѹ�@�*A�c��\  6���ֵ:�]r�P��fw��{T�cMl[.��H�ج����7\MJ���L橕��r��n��3�-��'I�D��J�JP���|  ��l�n��(��]r�uN�-�M�ts�S��ۚ&��kv\�ܖ��M[3�k���uL˪�R�wI��m�:�:�j	o��b�UP���( �� �>���f5t�w8]6�-�[b�֫}t�{n�4:Uʭֺ"�]۶Crt�N��)l��5�7��obU�ݮpsk��XU-������-kt��%"���� ������.8� 톕�f�Wu���p�������5΂�7I��S�'Z[�΅+m���7��{�Mwu{o
i�F]p*�6�aK�B�J��{�tԵ�� �}�
�d���������ή�R�Ε��kYN�fK��Hk��շ��s��N��.앪u�ڱ��ۭպ�kZ���U��WB���wD$(�$�T�[����v��L��s���mu�r���L����;����s���]ݼ���뽯n�t��[v�wmF��s�ݯ{P����KL�܊��u�P%(����FR��� �My�m���:����vW]q�]��M�2۰�tl+*��s[v�h�rV��݃��à��M;v�ozz[�n���7�[.]��=���tݲir��)R�J��
�k*G� 6{_Z�wn�5��u�B�wm�ai�حe6���N�.�6�Wk�v����M�:WF�v�[���h�*�Q6Q�H�:֭�ln�';wv��N��~BfU)H  )�IJ�4 4 j���������  ���R��  "��S��UM d��
HLʨP������g��[�طO��@���9�]{)ūK���cB�Ėh�|͵�����W�_}������Ȃ�S�Q�ED��* ���QE9�_��g��w�uw࿱���,�դc�n�IJ�ʱB�-�w�����lV��1x6a�nт��u{Q坑�P*j�V,�*[�[�9qԫ?R�E��Tk~�iec��,b�AR�Yz�;G2�<Ͷ��ɸ��#�a�.ƍ��T)Q�ifJ`��M���Eb�JIf+��RH?�R�Z�mn�����Z�ú#s#��v���Bm���&l2�X�
�ʚ*!�� #��h�Y�1(F[�b���gs�ln��fn���GEc�X��YGh��0]!K$�r�hj�"�'��y�r���������m�4M�ȑ�%i�`]d=
)4��jl����=�nYY+r�i�H!���Rm�V[��n�J�w`S�j�;�5��!�����+r�����Tȱ����.1z[cI�}x�`�fʗ�W��T/�i2�����1�ܬ�LĀo�z��0���dZ�J�ST��7n�j͊�Tv�����qj�fi�K�)r	XK�eJG/hb�{�J�x.臭*+Y���NૠEJ��Sܭ�H[�	�2���bY�����
�L3���t���K[-��.�Ѓ[V6E���@]�z��͡�i���]d�1��%R���U����լ�-��.eN�bX+ �L�S)�q�ʺ�B34H.������À4�fS�ܖ�-.� ni��'1ӣ
��{����lƖ��b 7��cV���&\�f���P�9�w@X���nٴF�Q��*�i��z4�1�a�JZ4ĲE��j߶!i��7�:y �(bP���m_���)�����S��h�gY.�f�8��Q��4�n�*lã6�E!V�i��Z��Ua�tk�͘�,c d�n�/��ds7S�,���I��{f�:$�̭
m��a5fZL�&8Ք�V��2�v�f�kShh"��R��]��ĭe�N"V��v �ZfI�0*���!OZoy�(E��%do-:�R�uh��HL��]�])b3C�b���
�ˢDER��@ѱ6��B�ѽ�.4�[d!y*�:��
��@�­�[BԿ�ooX.����E�Ɩb�AN� �z0k�����
ܚ�u(Kc�X�T�ES3H9:`ð�	�7D�[�☲�7��kHMR�h��e<Na��Ce\L��H�M4oJI�d+��ɪ�h�j�ݺR�4�֊`��4����W,Jm�W�����.��3����Lb�6*
��g%�+*�^ 4�o[�	�ěHػ��{V(��Ŏކ)k���̖�Z�Z�H�yIv�麚tf/�IU��HZ���x���*^�Z�w��ٺ*b���s�L;kZ�l���h�4X*3W6�Ջ�c#�ijz��MAsnX�f�z��褲,��9��&k�m�L�ff��mLT���f�tj7f�F7l[Kk^�v4�wJjf�F�ʻ�'2bqc�!�yY�I*�ق�ޔL����H3X�ҳF�N<p�L�b!k�m�Xj`Q��(�oX�t ��zijqK��I�5n�5mJ-j�v���x�@bsU��XQk��zo��Uf�茖+1��.[v�"��g~	$Ņ��*�"޼4���!�%��!�A��Ȋ;q��[B���H�,_�4a-�v�DL��@�{sC��B]$̢2�6�A`=����[ �
��Kh�m�0�0�#1]$�J��2o>��x�`t&�Ӄ�(�Pm�Y<f6p�D����&AtXe�vM��C*�ʕ�QT1�ZO�*��٧S�t�ɹ42��N��U��v�<	�����;�-�k)Z,�I��a�]�^��2n�7xAuxޏ�7�dnV����7,��g��(e����kՠx��F[��B��&э��
��6�/�L��ݓZ��6��p�J�e����nd�)��d�@囥�s y�hM��┅!#���84�m3��Z�yk�=[DŲas���w]%p�8�ˠ�Y�S6��t�1���Z ��K����CHZ
���<�4��y ����`J慱�h7�13��z�h��!b�3Ӳ�a�L
ko�V
;y��]^�I�m�ӷ��ݓ�5�fn��f�h�.��0����3�Vk�C	�DnZ[E4��{�Bh����x+p$�Vŗ"�7��Tp�����M�WHā2n�5���w��nΒV����%V���wZ ��NC���ùQ�q|3n&jM;Sl�<�I2�M�AЋF(�V��i�&䎐�L�D_�6fZ�j�zp��v�g[������^�Ȭ�L����ϷlcH����Z���eLr�����R{�,u��fn�su�����wi�oZ�6:E�Տ]�+UǊ�W�n�&Dl�%�y�aUg*nV���.杖ĚX�Et/���7/4l��2ջ/5]�ӖK�f��2lze��X��s^B�A�����(�z����kY"�h����� � ��Tq��ǚ,�䣎��Vv�J��,�ב�OB��SF���1���x�lf�sNAIЦ\�w��N����J�U��V=n���&��S��`
,.��P2�(eZ ��Y�-^�	�M�9�V��{��T^L�N�Уy4�ra�eާ�mږ��q�Q���N�Nn�`�+Q�ͼF���CElݺ��;�A����!��j��� ٺv)'��Z�e��SRJH��ϖk�%�A�]Ч�Y���4H���=��u6�Y�2��Lא�.�� (e�����r��;�i7D�*e��Q���R�c*�m4�f�zP�.����T7f�u���U�kr��ژ��Z�u�ƒ[B�1�����q��n��6��ÖC�^<��-�5�Z��/f/jd��3m��]Y-�V<�l���U��hM]����0���x�3][e+6�ⷰkAjB�,[N�Ԛ���aHۆ�T֋oM5�{D���dԩ`낢md�[��1sf�Y[�ةp���g`�ۢ���Pa�슰��tq�EGd���n��:���Xd���Q|u�A`�������kop9&'�������1�@�ƛ�ۣ�Zá���
��H��
�P���x5$J��EFÛ���~���8j �v�h#�
��Sp�ܕ�м�c�	Xu��CD��<5gҙ��N$F̭zF��CK1§�5���K���� :�t�a��ԋBÙ�\sqR��y���YlK����xv�
��ie��.bm�����w�\J�dH�eF�YV9+�oD�e^i�	H���Y�m��r�[��M�H�3p���MH�yfL��`B%�-C1{%;��V@���sQ�2Lo5�`V�<�d����R�+l5x�[t�(B�7�+X"��y ���#,`���)2��YF2�y�E��gC�{���ZԤ��`�/T��j�RSn3�����Ҥ�����;��_�>	��X��ԍe^�mR	'�*����DT�;�IGQ[�L���x���^�X̶^g
��[�m��4 �F��U�oh��%�r=�)�h�(	���ѵ�TX����D�b���Vs�V2P���ֻ���y�ڱDMa�̍�`�
�q�n�Z7�Ծ��{/P��֊�J����.bO
�-����x>�tA�r�\�L�F�������GqX�2�a!Pd=Uùe�Wd�5�\�	��v��`cL��	�
W=�͡�����B�lLHTEB-��H�n�KӽV걲mb�n��	�,����kL�݌���Q؈��A�"ɨ C[*��p�l���-ɧS��Nh�Gf���n1`=�6cӔu���8h:��A�m���P���%ђ�.Q�Z@�U�7�t͚x�u5,�1PyA�Cwl&7nS���n-f% ��Hp��;�[����4�uWx�F�9wK^k�RU��e[�,8�.�� �,Tmb[�X� $��s&i��0٪��U�:��ne6�n�m�SX��S��<�M8��7���;+0�����1�[)��˽Gh렖\�W���5(�`�o\��Z6,�{a$��5��CV �]�������b�ذ�^n,�Qդ�a�Uַ!�֋���B�����L�*��B��M��V��:iP��H��Z5�-Bc�j�˳��B�in,ՑrZ�^��Aa(N��e���Ղ����|ɫצ�]*@�q����Y�&FٲFd��2|�Ƶ�D��*�:��L��Y+;7A1xB��R�_<�e�K4��e��#I*B�4�����u�2�,��`��e�[[���%�y*3V`w���6�%�r�In�"1
���s%X5� Df< Ahl�W3��=��\H�.��E��%۬:�4@��Zf )D�E�5n�	�R7��WhRQ�F݊�/��'yz�@L�A��m�76���YK�QF6�oUf��Z7i'e멸��z�]����H�wr��+�5a�wi;.��Rvh$�e!)�osT)�2��V��V���b����s1S�E�P�xbSbe9pł�]�?D�5VT�2]JX���ۡj��x�Hd���ڛ����,1Lm�e<,�T����ƶ�%BZ���ɡ�A�%�n��Ow04*3�vM3]ӧ/%:�)\��07�f��;�ʡ�GQ���"|v�m�q1�v��5b6�i�vSu;Xժ�ڕu��_K-��n���N��Ł4�ܥN]��������ް�;.�f�r�j]+v�ʚ��<ۨ ɢ�fY,GJ�ҩ��p`Oo��/j��d�٭u���lޅ���ԭρ�QIq�Ժ[e���mU���,]!��JD�Gt<���)XAQ�ܡ{�]��g)����
��M�5'�$h�336Y�0�N���o.�k*L@aڂ(5��Cc?G�������d&Ri�ǎ�
Y	�
�t�-ѕ:ט�5z��\@��f�z���U����c#��s�T�mIAJ���J��)��n���A�-����l2�e�1j�:����#Rd֤l�Of"�뛗��ݐ��5 ZՐ��NnS�z+(�ź���-1l��oj�`F��������`�yV�K��v3,$t�Af���d���+F��!�Y�<�V�X͹��7one�2��z�%��`ݷi����m@H/)�,�y�]��ZE�qىc���� pK�u+���0��;P֊�opnn����"�˧�N�:yd��f�t�d��5�bj����	[km�pc&R��h�Z�Vo)��P��&���WV�S�Vd��Ԓڽ�e� �EZ��h�қT�X���	�O4d�LjdN1�/PT�pV��(��`���w>#FݻZ�H�4�%����ɳ[�K�ӿ�7w�hP�� ֬q�
�ܰ�$kz񫐑$3[
D�b�D�S���b�����Y�ȳ���&1l�uf��n�@��HJA���m0��Tc�
45h��2�f� �MX ]:����[����Ƒ4Od�CJ)��l�	�7\8���5*Jà5� ���H��vnLs:u�)��mh6*[��$�t�  �b��Z�5 �	��(ύ����!�@ue�f�����SsP�`Vn$hVڹ4óqKJ�6h݅�m8c�25�):��%���pL�Qd�����x����lTj�cm���-����ˉ�ɳI\���Q�cm�ZȨ�л;z�QuX-��,�E�Q�
�6s[P����*6���d�R�"h�*HtnX�C^�u��졒⳹tn��M����ͷ�a{@kna.Ԩ62�U�(�L�#x^���d=�J�Fh �F��WCV�+���V��-W�lzJꈉ�^�uyw�Y���@���#��:^+��ک����5�c�����D]>C�N)MYC�f���N 	=ɚ�l�fS!]չe��w^���	&Э�����k>%�}���+L爵l��v(Q�`]4iXN��Ӏd2��8hF6�weV8��Bnj�2\�r2�ߤ[m�ئZǲ��x�^R�f��1�!���H,��B-�)dݪ�z�@��ݢ��#V�,�K&��R����D���k��sg"��YYT/jW
)�Ym"R��m��N�Aeټ��b��Ln��JPhCR�'b��Lj�R31U��&��F�Z����B�ҫj�Ϊ+n�K�"���-�ae֭[��&��&�T�M�Y�	�o�C��ka���w(�X��Z�.If�ul����	.���e��}�;�DL���Iu�[����x�f>]�W#��"�{R^��}��*�"�e^R��ӗ.�T��į�����r�tJHLjLX�]=Xm��H$�vJy!*�M��#�6«��!x�I���"R�RV�j���	�[X�magHu2`��]	N�7Z�ٸ���a��M��)n)�=	^��58�b(�H�(Y��^7���W�����q�����nm9I���̵���ۀPX�H�.����Fn+ɴ2]ԌC��I��i'X��Tb����̙U���,қID��`%l��7L���K��,fѷ��h��f8�Թr��c�����:kV��;zi�*����Q�5��t��� ��T�E2�;y�:Gef�	�L�e�n��(]y[4���a��� �EKkQ�Z(�X��0a�����('��gKU�Uv��6��IaTq�*H/"ܢL9W��XbM�p��trf����%ƛ��a��
W��Ɠ&^�Pf<��q�bͭ����JR�ѩ"��6�OJ��94	{�E�-n0�ޢ�����/P�6%�i��ʖm%��VȒ(P���7�`�i����fE�]�p>T�s������VW*��O�`�9}M�\�,�7��[��v��f4����H�pb�ʡ�wu9��s�z�3L��yt՗�,�CW�۷s-H[��W*���2�U���O�Y!AV�GO[H�o*��j�r��rVqgt���sõf�:��酁��I��l��ٚ�kk��;�f�˹����3z�Į�/�A�T�h���\�okp���n�-Q������N�.`ͫS�WGWf�AՊrtnu��Nî�Lm��4�ev�D�r��_u�����+̋��wsę��W�"A�S�	̱�@�A݉�U�ba�
�=b�2�и��1i�Y��B���t�6>����0V+���O�ʀ ��,λ�2�U8M_9�O1 �p��KH��ݓ�u�vK�4�Âr]Y3�U>�j�No��%d1r����ԥ�w��լ���缺�E|�x)pX�/08`YL0�C�9�%O�����KN�!��M��:��V��Uh7�5w���鄭� �Vd;ː�	��9zU��wMp'f�gHa�̛���1��%k�ً���x���b��͔���d��T���35؈6���Ì-�Z��h�L��B���_.��z�VT$(�讔.r�a�"�ǵ%'kmuh�2�Np��*�T��z���9L��φ,B ��.�Y�T�IJs�8���h�����V���ސ���,�<�;�<�]�� �qoZ qopl�.3+����&N�.6���̭X�r���f	�s�X��;N��x:���맱%r��c�=�4n>��7gb9�"zՋ����:�M]]���٩z�����bX�ZMq�	��a�*��5c�ٜٗ��`czR&�����n^�Tz�BV�):���Д��'[y�)]�|󦱵��q��V
YU�Y���������k5ҳkL\e�!��]��s�VNoaí�e	�¾�
��z������+�:�-�[KXi�﹁Pk "1���\\F�s'z���i:�[��a�З6�o�}�<83�����"M`��Thhj�v�P��o%��Z���n�e��@���)B����IC��a!�0t�Y:uMu�ed����O�珄��!��v;)ut�']P��n�swU#C���OEc0Z�a:�7E���w� f�Gg�N�79�K��V��}�*[���j.����f��&�N�����Kl���Ĵ ܱo��iG|���t!9�D@��8��Ո:�;�[BC���*�C*c�o7�Y���N�Q�,"��GJ@�il������}׻1���,!���X�;tD��s���F�j�:p�iֺ�a�N=�O&; &��,��i���(#ċ��J즻�t��9ϣ�k.��S�uɪ��єy��9V\cn�b�{�TmVd;V,8���k�ޕ3*�gW��i�sAc�}.л�9���X�u�jHsu�tc���:0S���B&Du�,�7�(q����M�-�����o5�Si�Z��n�����Pb�a_��
%��#����[]��ǭ�J��`qw�Ѻ�v��dY�-������v���]��/��3#�rN���-�:���q�C�f.�ڴҚ�r,�,cGf�j��m��
�1o���)c��R���!X�8��߆�l޳+�k3�#B�j\���}��d{b.�͹��3c�"
ى�#t�<�h ��U���l�=cT�0v��Wd�iga��ؼ�D�;���ˤ��G�/q��b[!qӟ�\sT2M�X���
��:�f�%�\����X�&����L6�x�X;�d�KB%���l䡌�hQz~�F��[�&��]�ty�V�m�p��˙u>`��<�҆[O�������J��&Y��Ic�b�%�@��1�����4��l���(�xD�&���]r��}ʥ��b�gJ�-��`6f�����^)����\�>Ԑ�q���!��i�8e��,�䌇�ko/]G���y�A�o�����C5�h�V�/7�t��Y�z,
��,e��Vu�j؏e˫�}�-�.:2J�k%:ۍ��(u��B��W��*^-CȇD�ml͚n_"���s���u&Pep�w.U�h�wƟ�\;J�D�s��
]ۙP�r��3&"�W��$�O��w:Nh�̆D0�k
ͼ����v���e@0J�2����*v�.,��$:��¬v�Ь�%�Sonf"���� 9P�R��=�4�],w�:��1��[�w�q	w��{��J�8^_ew*7�|O��C�rǠ��:NeY|�w�]�p�E�Ka-�Y
�~�f�LR�d_ql��8�\�X7b�����D��wI��<F���mo
�b��r{Fqziǟs��_9�:�`u�1�)d$�(�uU���;Rh}9�y�ԭ:�����<z�͉W�w��Z+'G5c� ���c�S6�ZFP��+�lrWQ+���ts8=�P�U|��!JA۴���W���,�ҺJ�5�-1���lv4�1
�Y�ڽj���a�6b��"���������?�����])�5h��o�d��$
��7.曣��A>�b.�!��`��Mz��O�>E�z����_5²-��[�r3Z�ى�WM����h�Y�9�7�ќ�Q+!��R͚"D�M�Kg^�Ja��M�����+����0��()�/m_W]�c�o�tݣ@˾�M�[�0I!���V�{7rwp��4.�����M����ӥ��o"꺉�Ȇ`�]�v��y�[J���˵�;�eT[ט;C�Q��W]W��5)C�v�5m��}e��׽Z� �ݘ���e�{��r�)����$X7}�I}�<���I��c������6	I���,X�)��q�����Ed�^}~�N���x�+�.�����k]z��72�^���Gk���.����xii@+��K����eԏ �+6�Yv�6I��7vUuc�qW͘�������:�6��h�w�X��lh!�컽q���jW2塕&�1��(&���̅p�{O�T�Q�.�� 
�,fv�g\
�ݾ���r���Ǣ���m�g�0 �;,�����72�;-���OX�J���r����Um��{֩9�t�i�֖Υ����V������X��y��kb5�'g�R'�C�lp>�������W�����u��娲�+�s{���s�5��[��.h�*郋�Լ��N��7Gh[Nb=�dY�2�^F���G�\��"Ķ��yw���Uu̸�=�&bRW���wgkr����<S��e���:Z��'����PvӔ7��m���>fR��݁��l�JW������:�D\�m��2k��5t�mB�n�m����.H9z����jvU�lӏ��^���St�*9-��Gʔ�ˈ<	*��B��:L�jʨ�����c�}��#j��.v�nL��&o�>Vƚ�go*��v�D��.�q��#�vVu��I�7K�]��j�i���R3eEܘ�21�h�����O;;���B9ۛmR�@�x��Y%�d�z�F<���wwf����mh�oL}J�y�P�u 7��0ڭ�v��["�ҍ\h�tV,�@Ȥڊ��:IwEK�s��9�k��z=��;��[������
4$��V���PQ�u��C�2�ZR��W|��j�ꓢ�e1:Trf=��=`����z�ՠh��]Ҷ���6�حX�*�y�����)�s�y����#Z�� n��qj�������'4w���������[��n�f�����Ҧ���4t{@�Z�m�V�D��YC�Q�e�H��5�׋q�k��Tx�j��\P˫�q�4����
5�Xw)�)ބ�5�S�{��af���pT-�`��x��w�h�i��8a]{��Q�V�ϳq���*	��4ր.�8��-ޚ�
��[k�v̬���
v��lt�/��W�]m��&|E�`���D"++�#�c�ulO;��-AG7�m*�)���&+wS�i���n��up�}���5����I��y`�V�\�OJ�C��g��E���'��Hu�.��*7A�F�]�zyO����Q��f����{�c�+^��v���K�9���E<]��Prݠ�x��m���L ���&�<���9r�%`�ioBt[@�f�*�#�A�3��T��)�P�M5�O��s���l�T\����Ů����G�ջN��{z���8�b��c��P���c8���S�Q���-�љ6S��`��aɢ�Ee��`�e�[͂,[��Ň�_!�P���r�b7S� 9��#C�;��pf8�ZH�.X��o7�*��> �`�Γ�:�S�U Xs�Z����dq�&L
k���+\����뤲���NP��(x{ ��0W>h��J��S���æg���ހ�0h���n���Y���^n�"�{ �Լ��0	��n���u�﨎-N�wN������1,��_Usg���P\zf>s��3Wڋ�1��k|���W�����`'�]Cr�.��*Ę�Ň�&�4��vk���Wn���o�֫F_`Q�#YMa�ؙ2����F�}Lo��úkh.��k��ƌ[Д\�z������qg}�\���@P��^��U�W}��\�𾦜�y�pc'un]<9�xpK*M��`5��_\�}�z�|��\�3n]���+��C�_o@;��;��Z��f�Χ�H�]�����u{��Y6�?������4�þc����I�]S5�H)w��bSq#[���Z�5b��f�#�K%Ճ
YJ�|W��8.$�����%7)^}jmnN�!Z73�e^�o#H�g��_, �[���=ݲ{\Jf%�C��,��|�4�a9j������j�,gŇ��n�NVG=5�171`؇cW�-�P&15֖���	)Q�1�^�e���s�Q�J��r��f��YS�D�y��ũ�s��Ӧ7�a�YsIڜ`յ�m5M�����7�aGP�$a�y�+�0�h��r���!nD
�P^�d;ފ���p��Yi�a"�o��s��;���ڧ7\-gt���I�N�k��ӝ����{pP�Z��Y����[��&4M��]Q�'l�OJҷ��;J�-Ѵ΅�#$�]ϕ S��'��m��H����`7�X��Wq{�M�{˩ʘ�^��^􂥘��$�n�����T�ky�bj3�[W�*�������b�[��z��u��|�oT�iU��O[3�hd�y|(b��"�:�mе�ڳ�w�����A�u��U4�/,���W��8���Cp�A�a�����+��<�k%Ŷ�D��-�t�&��]+qIG�[\�WO;2�s�oa<5+d�u`�AL��V�d�f�ʙ;+��$ֆ��.u3�"�hi�ҕ����[��lI'�
��$�5��7f�L�B��B��"�$�v-���+���u�Fs�t�Z��=[�$�0��гz�2K��x��i�t��V1�.�ɬ�J�̝��T��!��f,ceXz���dB�a���(9h�� ��&�(n�ۼj� A���k9p�S:�K��)���;�~��V&��E��4�=q���s%�Y+DS���i�"���#��fP�r��x)]��7�*^q�E�Wj��[2l���n<�S�hf��u��9��b<n�1�]�:�,��Z]�����;�E��*�NW2�����W�-H LuAP��b��;�D���y�m )�tͦ�Jݧ�ݷ���ϲiIX��A�*㎮�����s�2��%p�oAe�7R�jm�]X_^ܧ0T�o0�ty*!	��̼2�Y>ތ�S�B_k�s.���ا�����5*r��pG%ձv�;ώ=�LCp�"�����U�uyH'�/��6�Β�)<�Jb��h��ٲ�]���X�θ�Wt����s��V��2;a3�k@��P '\�d6��Ͳ�\��omY���q�v�c�WaF,y��dU���mr��p�P�e	+�s������eb8��}ؕqB��ܲ�[m��B��Ȋ�"�mޢ�,1�^ͳ�j[�}7B�Vm�k��w>k&=�r�叝�E�VK�0�qE��F��0Ԍ����H�!03y��)���,�����h�-�-��x�"�4^q���˞{B�%vzzG���x*Q�}/{i��O�������wA��M�.��7�lG��9S�|o{�d[�ͧg�ފҬ�/:�[X�M൵�]'���j[��]�F>䔙��w�22�\��4�T�^j
i1��ŗ{p΃F�x�����9��ޗƑX�^�ʿ���٢���x�)��[����4+)���r���<\�G/j���*��zd��Ӂ)1��{jIس�u����Ϩ^��OQ�u� ;ˣ��Ul#a�B�w��U�͡ϕ��V��o�*�U�pw%���hsv�8��<(`h_[���.�f��s0�S3�*6�PLou�2B���� ���_Q���g`�3n�#��uF�RZf���!`���^rATSe��u���y�7C�=�C��%��Ҷ��N�$ε8Ӓa}Y8t/�f��Ϥ�m;�����!�W�i呵A�<\���u9D�a�_pV�z��0���M�����z��!�2t��L�pe�\�+_]`�#1�ޤ K}(�Z+�����Y���'�+J��W�һ72��gl��tOw�Zc��r�xo���H4���,+��z=*u��2�ם��i���ass9ՠ�2�L��[լ�C��_ei��J{��f��إ��ܐf�[�4�{�^>���Ot�ĵ�j�'@f�u2��bʆ�9:�}w��������@QO�D��s�}�����Jp�s7�p	ID��Eܠ�7��ֻ���J��w@�"+U������SM���V�WV`�@��,�Yt���ژ���Y,�	ǃ�6f�Av��eӡVebv��/Lf�+��`�s8��g�9biC�]6_p�3#]j�l�x�۹�RA[vF�	W���5nԾ�N���՜��w�c���So��T�cr�F��du���l��5�F�(����SRpi��ʶ��f˘GV���F���n�m�����%]0vd���G���}�ƫ�Y�t7��Cʹ��v*Xk���-�{�tv-Q�izs`�Xv.S��z�'�P�=�쳈�ْ�n�o�Sw�T����5V�m���H��JU���`�q][��̝.Ro�S� W>�U�����n�j�Θ�#�..2:"r�_2�����T����3C��c_=�n�=A��@�Q]� C�]_JZ�����]��K�cvމ}.[��O';��ɠYu�e��s7�[�:W�%0� n�Gu�g9	�7�ƒ�w�Ef�UgsR[jf�)TIw,Y�#x�|�*}�N�e�v0#M��p�]�zgǦ��������p��t�]s��t�VlgS�<�T�2/!&T]XB����Ey��|Q�@b����g5;J�:K�`o_v7��>6�#ZT�0��;��*b��*�{ϓ��G0����a.ru��2��:�F�C�df[��J4)J#���.��x��[�VJ�ۂ>��1U��~�����ݚ+�H���#g���X��	����2�d����Bv�����]�]�xs��[�ۙtZv�oW[ge	R�b�ӣ�Sk�9�[l1Y7�҆r�0�/m����Xa�٢5��핊�8ͭ�wJb('i�ƃ�uM�e>�$f=*��]�+N�N����6��w.���zHٰ�b�W�[G���������*�[Be)����q�,l�A�������3N���.]��ҞV�)�0Y�rL���=k���YN&�,�6��^T�Uk=F�k�ss]�W��{7f>�
�8F�pAe��=	�Z�.���=�K�A�Q�֏�l����s��b������PL+&� X��QU�v�L4��Z������Th�L1|��������� *�P_Z�d��"^uu�y76򍨝�k�޺V+�n�vk�1�*Nbp�yʯ7-A�7�M��hF�����q�&kbȤ)-�{C��g�S�� ��*Z��`-_&j��X%`��������ᄙq�u3����֝�?a�5q�Z��5�+vf��Z�#��̥v��},����H������!��C��h�L�S��yiV�:e����ծs��XJ*�Q��j�Hag���u:��2�8�E�c�d�i���vR\��4���(0K�2� wЅH7E����$aN�5ն4pۆؔݫ�GP��[ΐV7�P�m-!e�Pm�Hꙙ��M��z�8�R��le��i��}���mR�@�2�Nf��<���&E��
�U����$�P!��r�]dd�]��j�"�$x��3���&�W���Н]��W6O	�]gd)Ө�i����V���eݮ[ثM�e��1��jZ�W�n��ӧpT&/>�
3�5�TYA���z��U�p�b	�4�7�a�|i�ހ-�utќ����r��Қ7f�e<�qSY��br�kź����
;��X�!]���ٕq��g'jj�\w1�j�^n���}�Rч&Tt����z�2�%�:��Е��}|�[uˠ�ڦ[:�;l���3��p*[}���XڱJ+�.��j�d.o������U���0���D�F>ܖ���6�gL�SAB����%��	F�G����>K��Gk��V�� ��f_J(�����/Ox4T�t@'�ef�S,��|��$�5;<�`�F�ɧz��gJ#��+8.�(.<�b�N��D��},���s׹i�5_��6��,��j���܀��["�*`$���W�/��)(Ea�o)�ݗ��),�ƻ��h��гb��uՔE����h	�x�����F�D�pc�`ٌ�8��wE�ld]�<�z��g��s|So���
���\�z�<���:��q�N�3z�i�P�Ь���h&�.��:N�����w����
�T�����L�P�Zz^�|���Tm�g+UY#J�a�4.;��4��ڄ��
�r��Vmw=
�+]�Ԭ�Y� *��_�z����K�p�� W�g���A��&$��.B�vĩ����mUP2�h��xfǑo�m\������Bmq�MŇ��lf^u=<�m�i����ÂZm�N>v���m��\h�q�i����w#�\e�4EnM�)'0��P�{�Iݽ1+�^�Э�<��������ƲA���ٸ�|O*R�8S7fjGo(��wܫ���:_��S�E�Lɇ�NX��u�����OWt��jБEgĻ2��6��x���ҫ|����W_��Vm�2ZUvzv���4��J���h����x���s�4}$�m7�k2*&���Ǚ� 39���7��N���u]��$oE�29זu"s�2��=�⮱���w�͹j��4I��)�U}Z��#x��3h��L<a�f��)��n樂���vH���V�L6��ˤ��+��t�_�Ɛ����뺻�8e�̊Ֆ%��E:-�Ċ�R���­Xv�i��TG�t�\��2'�P�b�䬙cI�+/��� ���t���pR���WCb�L�gr�C�kT�׹�[i�;���2�t@�h��Ԧ��}v��'n�����jI�_h���<���;!s^�V7����9e�B����N�8�V�jLwcWV��n�Ӳ�j��������\�[��l���K���]jf�Om���7�2n��ݘ�kw
�=�!����]݄��}c���ՊR��v���N`��C**?]����"mf��rח��r^�S�6	ǠA1p-��!�n���H
��3�ǉ�W�H�콰.�Fylt44]�3K�.���2����)�Iӭ�����Ke�����^�)�10���7�#wh6�a��� n�P�K�Oc�A��wx�i��GT�Y�l@���н�9ϸf*Gu7�g���Uu6�:�7���u��ZtT�jO,�OSa!ʺ���_\�IE�.���f�̮��Qs�$�"(.yD���-;�h{�	�oY��� �|��`����5[�����!��>��>�,��8T���}��r�m�2�~�B��w�}k�t�$�n��p�=Db�[[��C�Զ��x�G�䓾#8YۋB�����d+ \�eY܋f�ȉ'u��JUë[bE^8\i�˽oV���lO�`�30kdZ�'.�aܻc{O�#���P��.��Z+Dė��M^+�cz�@!�*CR�p����mL�D�Ű�%q�K�q,竭���d�E�M����+,�B���X6��飋��&��S��Ww9��r޲�ᷴ�;.N-P�P@=�e�Y���O.��\;��\�.�~�{�'n��|`v��6�b�R�I�l�U&d�|�[��K��2�Yώ�\��.%��Ʈ�md���wohD��
4��,����d�(�-B�s��2dU�X�u�o���My��8ٴ���\����VG��k
]2�]��=u�t��ۆlKXi��`d2RYHr\������|�^A�d�v� �\/s��$͗xSCV���6b�����ͻO��۠�@T�����9�7a<��طJɁh<�FU�*CPU݊�����yok�����ԇt��i�ɩt{]0.��ZL�(pyv��U*�o5dL��^���ep*J��@�5�-���+@���������]G��w�\Z�W, �����V���'��YW-T�W;w�V侦�Gm� ��N�r�<r�O*}��9Ν,y���ʙ*Q�xz�]iY��㘂��K�u����7�7��+d���>�x��Ӑ�+��x�=��lvo�]m���d�	���7r��/�J���X]j��<��[ouh���ʨ��U�vi��`��ףu��(y��|��Kƭ2��mQ�g�y��p4o��y�M���Ԏ>�ۜ�1�-�vkD�������r���`����Q5)U�,}�(u�u�I���}�]9˴yFd�5�XL/e���Ӑ��Xy9�Ȧ�n�gY�wKX���b}F��԰_�M�k`tЭ��\�$f�]k6�@0�Š�Gl�ɪ�֟�0\t���s���n=C#3F1���MqOnc�Ƶ��iX�[r�	�W��jX�L�7{)en�T���x��7�)�(����M�F�&��֌Ǌ�
�j�����Y9��aܗ�^N��Lד�N�R�o@{����3I�����[JQٻ��n��y��|cS��	�,#cO�8L��1�-�Ӻf:�\[geN���Z�8 "�BCz�B���x�EZ�J[q�V\I�œAr�Нf�bo�)�t�m�=�[�GU.�B�u�b݈����QoTc�Ҵ�#j����,u�n���c�[X'gbt�ZX�Υq[����T�R��K}a�a޺�5hIeݏ6����a�F"�����xl��A��X[�+�5%�*��v���oR�'v��s2ڱ�3�6�;���c@�LÏQ�6��Ƴ:e�T�u��P�o��p��+-Lå�WG�ܧ�o*o���[r2@��'K�sZ@!�/E���}� �9��B������}A�Qޑp�Ҩ���G-@�e�V5zYN�Ƽ�kvT���OY{� w�Z�<mɃ���:#��b��w8"2�]ܗ*�|uSJ�e��軩��[�:����C�ӝ��):O�f�fKl��b#.�ꖶ�m�h弅�X��1f��3��؎Ij��2m��q�7ʡ�@>�
뽸��P�5٨)��87rG�`r[@+�c7E5�!�M�6�L\��	܎�gm*Ik& +�f��6m�-�&��{�:�|L�u�4n�c�dlw>����z��o=޸��$�k����@S�f�ɽS6�,��s���Ǫ������}o������cm�y)�njCc��R�A�
�c�|��s5�9r���uw�Yj�$H��ɋ�T<�65cϻS�p`\חۮ=y>�Y=X�Xs�ٟH��g@���:^E6+X�g$��r���1�:^�QJmp� \4>1B��c�t��͖�fb�}��N�Y[�닝�n�`<���=W��P���K9eV����w܁��yCVj���9-a�ݒ���d�p��
���g��]̱���M{�������{]4%_v�1�����k*��Cq�.�K̈� `Wi5�`e2���@��)26�K��u�o>Dl]��Zx�][�ֻJ�\�yNSYY��=A��er��(�nq����
�CL��}�v�kHm9��wY�7/
�����4�>�U*��@}�&.�]���֮��Q4�L�s\��GZ�Ch����H�;��Q��F=义W�ܩ���T:�x�ueL�H�0u4wxG+`�X�m��7�M��쒻�X���Ig.��U�أ�r��w�n]�6���>�/�_ B�Z��͡�u+y'ݴ�Z2�$��\6�ݱ�E`�gl;}S�ϴ*I�\��j޻�r"�	�F�Y���.����L'��i�gA��m�6���n���eX��@k��a�+&�Ԑ��������Whu>Ձ7ǁ��@��nd�AR��=�ӫ�;����1��x@#GudF��c.l6��[�@|�%�yǓ��Wܓ��J�G�šr�6�뷹I9�P��79oTNb��F}�s��Ԭ�Q�q��Z�jv�p�>,�����5�&�YYjN(�< d��n���5�YVy�گ�!<����@9�e��L�╃�:Wm��4�W;ᯔ]M ue����b�wS�j�J̒���wwlů�A�j��H����;��ӻ�aU�Tzm��#ŗ{g81Z�4���(Np�,����{ˆlB5�Ey�Q�(&+YZ�uc#�V���f��9NBX�x7:��r���n��+J�wc&v+�R��w@�f漫a}3�RA��brhNqh��H��;}Ĥi���VI��Ya8��8b��	�R.-�¨ܝ�*aYO%��[(��u�ˢ�VǛAk�2MF+�j y<�ʇ��P��ݦʪ��극v�uy��pWӆ�+FH�>�Ζ�s�O���`ņ������l�;�d�5l���ݛ�������E�����Gg�DhE��dv�c�]r�ъs�C���&�j��e�v�+�v��g^j#n�R���Kw���r��ړ��[��b�RK2Y*E�����[��;���503��v��H'���"�}E��w�{l����]9$ͻ�ﭳt�7LqL�=�Jn��]�X���z�u�ĬP�{�$}c]�t�
]�+p�I|��S7yl���hl��jc�Yo�81f�(������j!�+��y�2�����ۘ��'�1N!@P�7�6+��֞{����0M:�+�ܳM�1c��9��-��w���k�����7^@B�߶�m+�g���#�Y�H'YA&CX��9�/���9_mlp)�$5:��jv�k+k#�a��
R�����e���2T;i�"�y2�sA��"ɼ�V~��R<�E���GvP��D�z�� tƁ�!ި�/A^a5�3{��Ҳw����u�\AS��7�����ݮ:�d�0^j�I3�}�R�Qum<@!DU��]��x@�����nN6,c�.�ȡ�ӫ��ux���s*kVa���<y��#�������|�}uU3�:h��"���YI�<4:������竻Q=������Ѯ��Y�:���z�pn��e��34+�S�Ai3c�ɚ�r'����F&�>Ş��k�f+�k[Kԍ�}�����r��s���AeT�JU;WRa��'k���.�jV��D�Y�j�#����I[W�Jm�7���cJV5��.L�%��S�$���^`��}�(ᶌX5͖��]��ۻ�x�u����^q�2,㔦궆��K/��&1�	Z����Υ�S+���P�9o.�%�Z��u�Zq���.LNv7Zk����qn �Sa7���a�j�Q��\�f��!��\ЫNw�z��MB�qZ49��=�Y��1SE]�)f���$�R��Z@�bF^2����%Z;��vA���D�Q�Zr��F�x8�Yb]-�<g�z�>�3�І��lh�������,#���}B�O��%�5�O��bU�w�>��L\����#U�o����GA0�(�ȅXы
�^��"G�:���Q�u�w�{���+M �h���)p�s�rƳJ"�C�7�bi��J��.9��9�uꮶ�G�U�7�ͼw�`ܣ�oZ������Fr�m�yS�z��d���Κ}�:��}k���/�[�]��wy,�
��nE��CŁ�{c�Y.ZUw(���
��6�C/�0v��{��A�}wpUdNa��d%NM4����YfJ�!F@���4	Ja9@UP	�M	A@Rd�D-BPP�bTE�a��d�AC�R�M�4�QQRR�d�VHd�M�f�fffbc����d%deYCY&DE�EENM��PUfTC��d�f`DE(VAf9��X.Y�4IFE.IfE)IJSP��!f&F@�Y���E8A��XFTى��@�.B�F&YfaU%PY�fb�儙�de�`Pd�4�V`�f9EE��T�9��T���1��AQEYQATD5BU @QT�����I�YS�}#5�>��&3�ij�}����w���02�ցQ(��f�v�5tn��t��ۺ�¨N�q�n�y_��Xzs����4��D�:5�[��M���3�㧨���9={��Ԍ�B�1�'M>Õ��|R���2�X�=�~�����%��j8=�-��*�a�7c]Z�tM�Cb��Dr���EV�.�P�o�wdB����l;;®�����y2x rm7@-~�'���L�wfg�̚��bKbÕ�Zy,7����^�nK��[����N�P��Pߦ��3=�jG�?9�}=KЮr{�x̩�q7�ؓ�t�g�&�'��;i����|���ݾ����=���K��$���m�sf糴�sv�׶���ymy�y�_7/�C+���c�*��zlnK�����wܞW�њe���������׷�B�}_��c�����N^g���G7�V�њ�Ky]bɏV�>�7�������qtN4.
��Ų��NtƤ�zsކy�xa�H��VS,QLݱRJ��c 'Ҳ��쬥����E��u�K�.���!A^�,0UXP'~b� J�B�qd׈JsR	�`���m�75<���])}V;�T=�a%���5}R�֘8�˻��mL}�v�Q9u�������fI����C�e��"�˯�_�yo��*.�V�ˠ���f�~.�nt�c*no+�Z���I�cc��5��E���@���u+���;�M�Wuw��Z��_T��E�#H��oJ�9��X���Q�,�u�C�_W��Ɋ6�응�+l���/��w���Ղ漧M�$��tWǟZ��&�!ʶ�Ʈa���c.[��y�w�~���g�����:��6a����3�Ws:l����ھ.�g��5�J�v5/pI/�}.l�C���˦��7f�7vK�:�����Ru_���ǨnC��o5,t��EO�y�z�^��&�HT�Ұ�	��ݰ:���P�{-=�b�P��=u�7�u>orW�"��b�͸�{HK���՛Z�Iu<�:��g���ꛓ]��m�ܺ�D�g��ӑ{�89<�����ܺ�6������=�N��h�T�]�Tu*ՊE%������ve���)�=��b� �)Hnݼj��y�N�5��r }u�i�=�W��˧�
�֝�ci�=�4B��)9�7��+�d��v�{(<<j�v9���y������\�ކ��Evr����{s�/|gl:��s'�*�`I�N}�v����5yZH�РС'�l]xQ7*�����;s/�lg�o�����{�}�+���ϖ���K=�I���,밧������`�[�y�s�Y�|���}��c�ˮ��&���ٜ޷x���`'�_[V�/�\6�<ݨ�Nf���^�y�t��$sz��ua��4�/S'g�0��p���A�y~'unS��i=�cC��5��?n|����82<����̼���z6�'c�:��|`�-��V�'?xl۝���G�Όz��og{�u�gv'�n��/C�:3}[�=�D�3I��e�ݬ����A��fꬫ;�MmnID������B����7��'��<�dyn����
�i�^^K�����{~�����a*���������uѝ���oh��v��{i-1J��^��\m�M_K��].�m���z4�hn&957�����PJ��Gx�y���������qR�ު��O���[�G]��y�o���{�Iem�:�&�+Z,bY\5�a���(7�u��$L빉��������9�Ϧ�=��V<%k:h.�WOhd+קϺ���r�:5ʜ�{��S�V�vk��dg�+C�6V�g��WO|�P>��Gc���`lm����>���h�$��<&p�ܮŹ���K&?zV�x/(�]�<n�f�=��cC����=BL��Vt�yYӝ��i�h��f�������t�����3c�(�9����[p�|�ti@�q���X>�I�s)�?���|��r�Օ{<�{��-�[1/�r���x������g��D�i;j���ݨu/��u�������z�t�it��m�$��)��m-C}i�^}�q�A��
�<K�3�z�����'.���q�˓�&P^��LEl��.Kw��>p*q�x�o�X	Θ�ޏ=�w����'PƼ��,������5�T2s]�-�ޓHrI��P*�ut�-��X�@3ұҫ��jlQCz�ݣ>iY�kkR����En�+��3뭤�� |�q��x�iL5����h���EY��������7�$^�.X�1��h����2bfN�y��:�^���g�����nl���Nz��*��8��]̝{����*�f��/���1��-Mr��/�W>��8��Qr�{Љ�fu��yP��[�_�`�t�ή������^܉������X��[�w�R�����<���l���*ٍ�8ׇ+s}W�����;�w�K�ɕN`v����NR�==X���݅�:�}���}h�*T�{�5ދk��/�j ���z�"ѼL�u+��F|��3�q���2G������$��D�\��
#=E7$W+{�&V!�W���~�VdK��zK���C-�>����|o�!�mn)G���;74p�;Y���w-�n�����`�-��Jn�/<���/�=9�7�nƌ�����2�<�Ͱ�՜X�6>�ʜ����5*�r�;:�A·~�M��%��m��e-[޻h��^=�֝���V�;��c�*��\Mv�ͧ\^�f*�d.s�ֱ�������ր59�&�AN���{�%�|�S+��ȹ�/���jt�ν'���V9���;N7nw���]}���.^���*{�Nd܏]'�ugdՅOԶ�h����=��G�`�d���75\�lVG��p�z#��^e(��n�1����:Zޚ��s����]���G�ӏW׭�#�=5���
aW���6��	�|��3{t�>���]r����硹�}��O������w��Ⱦ���1ѺĔ����z� ��b{~��^0��'��e��N�;��E�	��2nOx%����	����}�	��ɵ|�?xlSmkG|vK\��1VV,
�5�+����}p�'�:\�u�5�c��w��[����q"��۰��:K.�z����r��r{26���tu-����@�r *e0OH+��]o�f�|���ŒK���!(ֆ���k�ߊ�6��]��F`�Z���Vx W��Y�9u�z���ދ�yf������h�J�.��V,~�����_z�:X����p��t{�>D��%i����_k��yw1�G���>��Mg��Fۋ^Z������۴07�'q��9�v�k�{�y�BP�t�SUWz���w7�}.3�F�6�?�m���61����f�_�͊��V��'����G�tKw	�W��Q�[ݛ�|���0�3�׶�1n�xK�ޏ��ʶ���v�l������Y+���c�|�oDh=�P����r��.�vv4z-�%����˿ٲq�d������0oz>�n9��ǧ>�,�̼]�nq�;��u9O;�ީFm��_/؞-�b�U�1����o�)�w�^u� ��u2wS9�Sij�:�0��z���uz�7�\^���+'�\�l�}��ҏ3�I��	�y��u��Z���^dw\�Oэ7�M�:���ߜsX&�+P�5��x-��{d�����y�S���/q�>�I��G���?n|砣�||�-�UF[C%s��u�w��;]�v�ahxX�;)t�lrU��T����w~�v�%�����I�V!�y��8�h��A��Y��Y2�iv(�.�3��gzsk/OZ�]\�|+x�`+Rf�4fv�ᗹ!}jNl˶������o�aﻛy���V�cz�N�������s���xl�v.�G���f{^ܾOt���~\�?���q.z�u�:�s����&y��k�u�N���{1�ݾ�+��6�����
L���k�]7����%��}W��=�Ĕ��v��F��4��i��79�C^w*F�fW��|b���׻�m�u%`w�ì��Ӫ��Cg��$�L�N����o��%����y*��"�ܒ�93D���·���9Ǜ#>�T�A��`O��(G#1�����������=Eft
H3͟w|����Wy�7vf}�ѧ�W����o��3�Cx���U�3��Y�n�nP\�����Zڞ͘v�7��؊��p�=�љۤ��JYQ��P�ϝi��>q�v����w���=]��ŧ�U��b��(j��g�R�%��籎+u�yY^�t���8Zˬ��x���Vb��<ۧ�{�v��e�t�8�70u�T�p��2�K0>�0e��Ry��5�9���e�jl��t���c5���.e��of��i�v�]�s����3�y=��O6�C���G����;��X�hŏ�v�2zv��{h�ʭ载8uzI�}�#j�eO�a������8�w��S�����z�V�i˽q�s���������Y��ˏ4\Ra�i����W�l�~����gDzl��d~s�{����Џ���.Y�b�VS�����w�%�lm_CC�c��]76g�No-�v���o�Ƿ�{]�uc����ߵ�$��+l.ӛ�{��d%l�xp��<��
�y��3y���;\���u�9�l̿=�6������h:��G�h��^�Tչ�9�"#���|GL��<G��K)z�F�ђ0J�d�	׻��s����,6��t�s6����oc[Ȯ}���>�\U��~-��{�K���am
�y�45���1^����L2�Zro	o����h�g|g�b��OQ��1���[�:hg���L���tʚΞ�M�����6����V�
+����8sY[����3Gn�zH���]*J��`�GFoUۙ��:���2�(gB�x��]��7O������u�w;Y�G�����X��Z-{��?w_;)z�oem�r���ɭ�V��3�3�ʮrUae ��"��WI��=e;�1��.`xr_�[yTuw-��ے����f�l��<�[�0�o�(|.Lx%{�����-P�<���эT��ͥܶ���>M�^���u^�E���1;�W����ya�	���ި��m�O+�9�>���۬�A���r��c+ӛ�Ӟ*��O]�zݿN�������)T��^��l�Z���8�9�s�J��]�ųB��l[}>��T�׬/T�
��F<7ǡz�'!*{.����s�A��ΓޟF��I������v{�L/��[��շ�ط[��<�*�����=k�����'����N��c�����t�<����omQ ��G��n4J��T���5ydT��	��@t�V�;�-ެ$h��5�]�3UKF�'.���:
Ҍ�e�A�u�/\��4��/�D*�m�<C�dH��)�C�t����k7�y�C��y������c�����չx�ʸ�[h�F�	���*�p�_TV�gvVm�HS_	�K�Θ���]���v�����l�A^�^d����;{��}�>���rS�wg3�n����c�y"V�dث�M���7��s�v�r�ɞ�7�5��`�O�/]�\+��Z�%ݝ���O8�ֺ튝A���W��wZ׻���}��b�������j>�{Xd�H��^����M-f�eҸdt�T񽵛�m֠i�+�2C}���A�k9��h�hjИ��6w�CNs�T4xx潗\J��zvִ�P$6����veA#�.���?�jw�ڒ�7�,���S/���Ng���l�������zZ|�aT�ќ	�թP����T4���w����b@���YdE3�R^��(�lOu��26��+�No%�.�
v~��7��O�u�V�>v�C�l�{��5Y�l�ȷ�蹴As�[�d�6������).�%�h���pc�Ƨf�,�L�7�5�0����PkLT�W�
�cN$0�|ԭ���8�uT����r���k5<-vu5Ֆz���8nӧQ�l�=M�t�f�׊�D�jKh}[0K��m'[�G�Azs���A�����$wn��I�;�$��xE����Cv�7���h�T����1�p_Z˸f�N^͑-���y���ԓ��E�S�ir�­����-��u���z�	cs�8/��u�o��K)��������e�S��X�J����z��Wx�n  �_#9eu�����E�sO]�4�O��lakyF���xz�Y:�ov���
S)s+-��*W�YC���U`Uv0*Y��YD��1m����5apt���g�D!5hʼ�j���a�X�ߢ�7���}6����JN�O�%C���GS����'ب�"&�;+�ŧH�ͩ�fM�40e�"��E��{[�,G���_V�=��T6%ݙ 4>
B�c�J��b��ǜ�>��
�{��]��ɇ.|>6�	��f�!�%ú���+��f�t|��+G+Wnh�������y.���Vo%>������c_Ҝ���4�{�8����Թb�m�����q
�)j�j+�j6�_J�)پ#�h+�]�e���I�,&qWwY�֛I�t�]�[��Kxr݀�5��*yvٜ���9i��Ʋ�BXU���Rj.纱h��J�L]No;Y���<w�$Qf�XpY����Ǹ���o2 ���춗�����D*u��Zkt#�0MC�&�Ծ�fN���H�+����@%,�E�MEE)LE%5HSB�4P�De�U5MS��@RD�YS�-��EPEKA1���AED9d�@�UUR��Y�LU��%�AUQ3E3I1YQ1UBDQIM,���$I�T�PD�TSKTU1�P1	UDVc�D�M�SIM%	QIKAEd��S@�ҵU4UURSAT��Q4�EC@EIAQ@RPTT4QMDd�D�f9U	TD��%SDUIDITSA�I�8MSD�1IKFa�UT�DdeH��MVY%DL�1ME-��������z��~���8�A�j�4�pu�&��`��8�]g��}n۳���e���:T��Q�ߟ7J
�º(V��}��g���L��mX�?xl@M����:(왻�n�V�f��9��kw��ƽy`�sӣ7�`��)�Sq6�={y��v���[�.^��m�8!��I�;_�_q}C�Np������hMfJ<X�]����>�S*{�n��`>wS���!�\�._{
��{^2��op�f:�n�%1fiUx�0]����ܦ}l�;��a]�z��}����Ld�f�[�nVKxJ�w�[[k#��C�T)��/��D=��I�$�&48����˘_p��<��t=N��y���{r�:��\K���6}���\��3r]WÌR9�{�Н�z:�����cZV)����O�o���QC�rcӟt�NI_u����8fǾ���r���ߚ�N/tw�jV9��^[���[|%��	���gn��sw=t��J�t�y�C��Y}���f�=I�[�ۻ��cR˺^�s~�`��ړ�9x����9�����L�b���;&�u��k����`��;x�m�������Ȯ��Ow�9n���gG�������9�]�,A�}@��OƮ:���+y���+a����V84�zh�uI�f�sk�؛5�bF��3�5�y�������E�`�F5��=��9o9G���;>�7��9[��Qw�&t���<�>�V���֎>��3c6'�f��Ι�Q�=��՗Z��nkCѮ�g�P�	�[��E��4^�9��Z�d�ג�*��0�j�!�A�2��'a��	k�N�Y��N1����Onsa����3�����U>����|4(!�W��}��ov����Ԅ��{|��E=�׷��y���<�=,L!gI��CUx6��d��p5���7���c�IY�9��%z�L�r�;xPΚ�ͬ��wf\P}`�n��Ou]�֤�dقU�
�o�V�O_ҰKxJ�w�'�5�v��\�9@˕����47&��h�G��sz��g� F� �ö{-���X�M؛O�ڗx��5�ók~�rLZ�, ���)��MQ�:�Z-Y��#S6ʡ���b����%��&���;�Vp|is��J���]�%���B�-#K���J�%��jS��=�Y�2����m��܏���L`Iw1�IT���Z4T��p�W�_�)*�1���Ϸ�4�C�bÁ��|�MhxWZO������N�=���p����J_*��͌mv�7���\
ǡ��t)��t��=_Mͫ�9Z/!w�Zw:��[�ف��F��,���[�X��(��G�k�T��*�4�>�.>F�F{�N;�3З|�� �M�lޖ���;�����i�<^"�q��.��W��M}���'��m*�y�x
�-9w�?c�v����~>.��I�?���\�N��;�\���-u΋Yl�z�:g�I�������;����c�d���b�](�:ё�2��e�.���;~.���BfgaX����~�����'��7��{��{���@�d�R��`_L�{{
1}#}rW�51ԫ�̓N�7���9ܩ���a(��N��],��(t6i3X�gUX����O҅f4���ǩ�\�d�G]�s:�kJ�e I�������JS�,]���u�M"m��i��)���.�ݺ�}ƕ�.���3��O`P�Va7f�X]���<�����p�.	;{9�݉غĢ����,9о�3m��/2n_9yv�GS۔;w���zo:��9�nyK���>dB?}��<��w/Ѿo�#��߼�.���k����ߞ+�j|��%w{�ܼ��_b�C�잟u������z>�����iy��Ǉ<�P��t���ߚ\�H~�ӿ�?c�D���}z�w3����s��P�/��b;�����%w}��r�S߱�/��|����}�w/�{�b�:��)��z�{G^�w�1����V}z?K��������r2G��9��rK�yu~z�w�y�_���C����{�r9��oG��w3K�:��u��7Ͻ����Y��7�\J��
}������>뾎�y'��ir2^����!ְ~�����z�~��ty���%ܞ��9/pw�ܮFI�k���o��k�y���:�g��#�y�K��9�%��^Ϲ�(K��y�ܯ$�ߚ\���ii~���#�=�GgX��s���aB>�=���,Z��[�c����7/�s�k�B��~������G%�
C���y��roBd?���]K���r�W}��h|�HhW]}�Y�VOEX�sŀt�z~���C����]��>w�H~���
�ߴ/�9a��r
@�<ގK�d|�!�g �1���ӟ~��^�;��">��?n�f��+�����y�}�R��'�?�s��p�����w)�1A�w}׺�7g����W�����q�=�sHn_߰|NJ�?}���0zg����kW�S>և����'���po�O�z������(P��qf�o5�:�0,��8m��xq�mm��Qdu,�v\��C2��ʨ��t'2Z��
+	E�Tq�[jq��P�v�^Q���n����G�6�p����T�J2.�)�B׽�j��1����9�$9�4?Z��w�~���X�W�����������
^߿i}���O:�@�A�Ǒԯs�r������}�3�h�q͚j�W�y����/`���_o�.K��x>�P��������B�z������仂��hr���vo��>�~�A�L��x���t}���^~U�'u�r�y#���}.���^���_/�ޗ }��r_�n������5+��ΰ7+�����N��g׻mgp����2>g�C���%�N}����֞C�^�8i���_s�K�ǆ���;���g%�C�1`从���}�q��s���|7ƽ��~$�F���!��!�~�;��<ߺS%ܛ�^���ǐ�}��� �^�{�I�_c����}���2_`��[��׿����������:����>����G5������'�ԯ.���~���ϴ�r���hC�w���]�Կ�@{n!��0��E��c���Q ����W�7E������A@��{�%�
N� �<��٣�GOx�J�{��yw)��h7.��}�oB{#������B�o(}����������_��o=��;���Ͻ�7y�{������+�;����ش��%ְa�g	��u',����'�������>_A������,�����W{3���S�s�����w��{��|7ށ���:�wf���d���rd��Kְ^K��G�GA�',����I�>G����_�~�����J������p���8�ގ��W�7�:��@s����>�����:�C��r2��ܙ/����ܾ�ΰ�W�/���?���,ۉ�K�2���)�/�I�-7)U�FM�O��ȃ�E����-��a�2n��K'C]�x�iV� �����,S$��.t"c�V��}����==J��\�/��_<*�����
e�F�w���^�{���;/�
��������� ��i����?�sJV��O���u'�ގI�^�sOP�
��IA�}��s�|��9�Op���~irW�G�4�f�+G���7�e���I
����_��_��~��`>�h��%�S��4���^A�k����~��)]_�����
�sHn_ђv�z!��sΞ�z�:߼����Z?o�k���~���_�}�C�CNb}!�{��:��^Jt�������w�H~���{���$��r
WQ���~����y&���9ym���n������ǿ �����z������Gb��~���9 r?w�ԛ��<���;�ÿ�_`�_������I���r@��sһ;���=��Z�6D�~��#�������}�����������S���Z��y�|����ܯ���NI���5�:��/�9.ེ�ߎ�\���+�ʽ�*|>�>dî�?a}�v�n]�������~��w�!�_a����}����%�C�1N��������1|! �����ݹo����in����z�g;��w�>Ҟ˸���p�����w'ه%������r��iy!�?�:�K��!������ޱO�Լ�ַ�u�s���u�9��k{����AB�:�`仌�����$ܻ���7�A����د$�a�wy#�����?�a��?t�����9���������q�I?�&�ؙ�v�Q��s�`���_��a�_`��u����7/ђߴ9'%����2]��1�	��4r�˻��Y��;�_^Z�.j�[�l��¨����~prW��irOe:s���3���;������OP�]���)����ܼ�A��iL��w�/���.�΋�z'���+�_�O��w&u��}vVd�,�g�Z�����d�Oc��&�=��:��︓�P�\vXڜ\�v��a��R���z�/�N�^��T��8�R��rXon"�n<s�-�\��4��0!��!�u�r��\5��-�SX�M�5�uf?���/��s}s<�w�� yy/r�'�i�����t���;�Z\���wC�>��^F���y��ԏ�۬K��N���7�s��s:Ѭ�8k�W�|���}��k�{!��~����/P��.�r�v��}������A��4���wK�d��>�r���G�*�Ò������"�C����;o�����w	�z������h�_a~���?@zs�^Gr�w��@����^t.��~ir ��9/���H �����l��ٓ)��_㕜7��ع/qԛ���×��=�N�}���Gp�W~s4u/�{!�9�:��)�0A侜�΂��=��N_��e��}��4~�%�W3��|��u!C�K��jGr���ߡyg��%{/rv��J����<����接�'{撃�AO9�J�mA�ߧz�/�����j�O���_~w�'$w��Z_� :5��a�=��O�9w���K�<}�H{��=�7��>w�B��ގK�(F��{xA=�U���ص�����2oJR~��߼��D���.w���Z_n�2O�9w��:�r�;��I�{~��?Gr�O~�$}� �Ly��V�������n�i���i ���G��K�/o���;���>�	I侜�ν��^��K�`^���y/#�X����vy��;����Լ�p��}���`9���3A혼��}�H���P_ �N�ގAH�?��!��ǜ��?K��俥��~��^����֡w�`>_��;5�O#����ח������g�s�&�܏0�u.��4�>��+���rO��#�^������Jv�����{������~�_���C�Խ�����z��u����%W��~~�VS6=��R
fz��u���Ahf�c��խ׸��,kU\ph�{��7�XSi\�s�a�.�HxZ��<��1��`����ot.���\�G���L�ѹ�W��f�Z�W��Ń�hY�@{=�]�Ż��|��7�/�����﬏�)�_g#��NB��r^AK��������q��>5����w����#�a�y/��vw�/$>��\��W^��J����+w����>G�~����;���O#�~��c�`��O��|:�A�y���&C�w��H�NI٭����$�a�y�#���8a�,ix��|揄�߬�����rW�;��~��f'���'�n�]C���jW��w�&�}���y9!���&C�wf�iL�ru��7����W�+�.�%���~���?}������#�s!{�����@�����B~3��}����ù�%Ǯ�9J�d�C�����u�:���y�5�y�}����������|��/��ßiL���Gк��Ð�}/��o�������t:��y�\�<����'N`���y��W�7=��g�{��9���߾�xw����|�k���S�9�众��?�H{!�<�[��z��hm��Ǜ��w/g>���G�wδ����/�Rw��o\ϼ�<��k����������?P_}��'��9d��ܞ˿1O���r���~7֎K�{揭��?@~�^Gr�'q��4���;�
W�s}�~��{�?`Y��֊�mٟ|����ˈ������<���F#�}���9d���1>�/e=��;��}'��Gr�#�٧r�'�旑ܿAO��ֿZ��>��z{_�s{�{���>����_�~����~ir2O��rg%����]]�b;��:���?I�{惐��A���w#��;oG��w���o������kSqu�m���/�������i(:��)�x �/�뾎�y'�����]{��%��C�X;��yuvu��C������.����/QY��k/n�-�¿�C�Zd��^�M��:т��@�)e�*=�Y��"�@��zXqV��}��ㇷ7�3����q���6J���ea�k)>�-1R�ٮ5dw*Z��Ծ.�)�7Ҳ�f�X��I*��"�$3h� b�VZ5�Y�5�3B�u��ԣ�j������3�=����er2O�����Gg��ܻ����4����������O7�/%y��Z_��2��=ߣ��'%��[�˿��f��5�y���{��oϵ����;��x�H{��<=�\���o����u��仂��9���g ���&C�^{ގ�z����.^J��Z������E�9�����������:~��@a��*tw��ܽɸ|;��?Gr�
����A����)]GG���~�����;���<>��_e��ߺ����: zܯ�"������𼿫�];���e�9�Od}��o�ø���=K�9_�}��w|u��������W��~ގK����!ܾ��ۂ�Ij��%�_�Wp���c�|��Y����u�����=˸�X����;��=A�w�y�K�){>���K�+ǯt���zy��>��F3�?�c��v����z҂�����ѹw/���{��/��x��z\���p}���=��GR�2w+�r?w��)]u�
^����d}����^����+s��r%�����-���G�=�>���s�7/!��_��4���w���/rA�r]I�?k�K�w�5+�������_��Ϊ���~�~����4��!���C���#�~ҙ/$����^I������#��!�|�K��~�y#�αr�~�g%�NAޱ��]��}?���VW/ڙ]���V����T��'#�_��`r^FHu��C�w��~�L�ru�4r�G�~�<��p�.�xi_ײ�ϼ�5+�v�.C�&��	[���*?g�|����@GﬀO���{�~����w#��>��~��%��S�>�n]����}�2^I�w�{}.��_;���!��7����~�"B��:����jc�X)鬷&]k���$��8��	�j?D;�]��f�t��e~�I���[+-LV%�7�ZJ�h���w�M]�g�E��J=�eظ�9J%Ms�D}�X�e�[f�:�30�t3�%s�Q��˼�5�]��Ͼ�}����S\�w��J�?�{և �u�<�%�
N��>�p�{т�����Gs�{/.�>�˸|��n��=���z����_�m�������_��b�uvg����^���h]�r�~h)^A���A@�����/F���?Of�Gr�;��!w?��I�>��xg�6~�i��?o+);�~����~U���߬=��@p��<���N�9����:�wf���d���2_c%���u��X���:��_�<?r��ԫ-�y����>G��>���J�nO\�ܜ�߇3GR��9�&AԾ�Oa�iNA콜�΂��;�#!|}�ɒ�yޱw,������'�W��G~�����_�+����/�s�R���>��+��7�9'%w�3OP�
�|�Pn_`���Й�z�<�����K��<���82���C���ݻOa�>'�� ~���_��n5즧Wr�/�z��!��_ �ߵ�]FIѿtr
WWO���w	�bd���=y�	����:���z0Σ��'��T������������y���Zאk����<:��]�w���������=��<=�\�������R��7�%�2S^O��ecx&���rsG���;��_ԯﻌ��}�(K���ҽK���.^H�>����=O�X���y'RnG��5/!�?���r�����94'�~g�(�����Ż�\]��9��U ��p�����N�7��O������_�����z���hZ��y#�����ܯ�����nG��:�p Hz{b7��g��+������ϾdW�/:�?C��Z9=������仌���9/%����y/�^���~��d�K��X����z�r��_��+�*��3��߄����_;����B��oJd��r�tt5�^ֽA�U��n�	7êv$�����}Q-���b�"�d� �箲@��2���&R�oIΈ9yD!�G75*�:����V7���ḍ�V�;�N��Іu�(g7)��Cw��ɺ�ou"%GNj�[S�^8����@����� �����eG�֓���
�L�q�Q�l��F��>�G�Q��)��W�^��,KR���M�B���__�j��]��V�U�>y;���u3�sS�(Ӗ7�]Y�-V��Rر*nWw.찮�T�]�E�j��eIJ�2��5�[�m&�ol�[=�"���K�m��:�V.��@0I�x7��▥e)R�߱j�1R���*ҥ�vf��}ģ�CS���ɧ���8�v��[��U\I�8:�V.�3n����@�}�r'#~��҆L:���*I���=ԫdf�2�=bBb���n���QrX��*�e+���$�I�4t�{6$q��2e�%��I͚c�㇯"���U��`t���nM�mѤLwN�*K0-ݝ�����ϩ�r�R�onNV���T��́�K��7V�N����"�u���턒�V_��$k�y�Ƿp^P�.���M��]���̫��ۙ����i[՘ڮG:c[ȂX�sH�2�+�(_,k*���!�]&nPˮ;(D�[����Ӻ��t����9��Y���A)*�CA�ۺ6�!�����/�EMJ54�v[�E�sϑ��E���A��l,���&6���g�t
���K	�˧�.d�U�]1�{Wz�D����]�]E�;U�Ӿ&��]�9Hh5�U�<"�~�E��E����r��W�9�����FN��Qw��Mg�g��Y6��4w�S�e����������sv��zg%@�n8�=A��)���}X3A�*�a��V���&����RB
U�Î�+�Y��kz�Ȳ�����&��*�J�b����y��^�ƙG�%��eMgWu��g*�5{��_�!��M�����M��E�n��/���xE��$��n�4H�)HwcUƸE�vN�{Kj�C�y$Ţ�+����.ql<.ǈ��=7`�Y2�9n����)��s�,\��+4g.�b�4=����&�/�����R�ĕ�<.����ĺ�t��̹/]�s�d��w�N|l;�7�m���F��R�]��Œ��˓/�e��m��Z�4V�x���5ݥqV]�Z��5��ﻲ�S�AK&�1��Jk$�hf���u�<t�rM�zR�v\�����L�u}��_lqgt���Dun�]�����`�ئXNGY�uޠW�e-�|���ÌV�ҙ���o�ʹ&�H�[�ѕ�y������u�,�-�ԔM'�v�L�݂@;=��]�����*N�(�l��$9��>��
=X�l=�hf�@+��n����o��y�_i+o���W}р �5e�Bfd�!ERMDUAM5M6f)MAEFa�9	XDTAT�A$U1CLEL�QD�LS5PU4!0US@S5PDUEDD�QDS$M�1I1QTD��STUEUD�M-1Q�TT�S55SUT��MU4TEDP�T�SA��D34DDTQMPERQE$SEEQUIRP�EM��QEUMQTE%TEIPQ�1QTS13EC$41A,M54QEIMR�KIy�]Ư|��9#�����u��Y��ӛ/4��g����|��˱ƺ�+��GTL�4����ꃫ�&;��������~��k�����AB�>g�9�;y���@����꟰)��5�{'�;}rv��fKG����e�e���ww�%ҽt^/����x�o�n:3;'�~�q��|�>U���{�Y^u�r2P�"�XKe�Pu[�C�c�=-���Nl�=��Xź�����eXu>ׅ�{�:(n���'ƾ�76q���pޔ�ڍ�>r�9Gs�����.h�Ί���B���wN����Hc����M�S����v�9��d�y3��Se�3��>�:BF���(���m���%Aޏs����7�:\��%ؕ����pe7Sٰ�ܕ߯ܥ��RiyN�:�qל漕q���pI/�	s�+tsM��� �usrx3'[��[��:ĳܝ�&G�S��S��t���}~oӲ{���c{>�*�ؾ=����_���̗ٝ���W�t/+qP�����>�˾'�	��*�B�ޛ�N����Z-�i��k���(���� ���W�M��Ŵ�_>�<��֤_��=�V���BP��M�yݜ�cf�Z��w�V�`

�K%�ki�@j��5Nn���[��B�bL�?W��nan��r{v?���69�W�e��{k]�{e�O�~}>��~~��\HNc4>����q����X�Lzs��	��_V�{�לTg��.��5)��V��ہ[�̦&�G�{G�g%�����~P-C�B��E@�l>;y��?�Cڷ{�oG��|�gڱ��S�k�����rI�w���g{_`�cc��]�^������a�����k΀�M��^�t��ގv�#V�{��#�0�OAi�9]v������w���גR�c�.Ί����dP�����Z���R{��vk�G0!���]�'"���]��U�i���֌�*�6{�W��=yϣS�	�=os���t�u��-v*WZ�º���A�U>��p�Y���g���W��|'�N��(�Ί:���{�6m��+��Eb�}w�ɍ���c'?T�w|wN�(��۽�x��8L)�A�lk,�J����&�%s�>]|\"�{����1:�V���@*Ō��Uj<$����vp��i�+W�S��_�AzE�1M�]M�׫Cn�V2�Mk���ٽ6#���2�f_$�P{�3�eM�h:�y��)�f�<���� > w3��e����ΰ�����9���m��:\�_}�7����֕�ȇܵ�Oq�In�颹���*o~�^��(����|�e^,f1��[��Ӻ«��T�f=׎�O8���F��-�b�/󤼩{��n���b�XM��y���p���y:]�;����U�����R�oK��x�ͮu�8������qٹ�[�=�wt�����ֆ�[�\�oPs-��ݾ��{�q�c�͛�W�q�&\�GI�mP8�����[���OT�&�Vo�d�+�4*�݃cqiHO[��ӾYS:ӷ^�ۀ��%VW�Grz��w%�����ܾމ��Ӄ࡯؁|Ϻ�v"u����Z���C��{dZ��˗wԫ�e�P2[����'Dzs^�&畦��г�;ƅ��la=�x%Ve�醥�"�����x���y[Y:�v�Er�xwU�S��� ��eI���,�r�e�Ʀ�\�+8�,"�s�� 2�n�ދ��d��������Ncv�>�M:�+SA__é�̳�Km�
��]i�u��9�X�u�4pUcvvgꪯ�}pH��ֲ2_����ӗ0r��#��Hŋ��''w
�ή2�^�[v�\_�����e}�G���s�=!���ӱ�b2�t��%��s��SF�O��b���������&�I����b�$W���!I�iu�DNO��>�7�^ު3|��G4K�6�0ٛ�c���\3����hM���gE y�9���ge�ro������}�r���T�g6���f�[��xIdg�Κ�ZP�.�;vAo�|rŹA��M��+�!�=$Z�=��v��=:��Oq�J�n������y�}CكdفK�"��HkE�&�{~�v[)ߧ�����kk4�d3ܫު��_e�{ �w��r<�EL[��_H��=d�y
����\�)�� ���s��?g�هa~~'�</+��g�N�W�|oEG�d׭Ӣ��)���;����7�-���E���^��=h�X���IPnez(/@��_�efmf7W��_���[[^�VMtcz1o�l��%�T]�)%ê��3F��ۉ�d�7r�L$�܏kt)p�SE�-}�V�{֜���q�7���O�#O��&�����S˺�ݿL�`uO�K}a�a���䶧B��'f���Z�d��	ζ��G������Gx�������3��@s�s`{�62gn���S�ڪ~g'��_aNuۏ�cQbHb��b}^�
�vK��62I��<�l�ز<���{�!��^��G�`�l{���)����;jM�V�y�\�+,�����=���m�������/�M�����9\��WI�>��3M{@|�X/^Ŷ�Q�wCFr;r��To��x��z]|�l�옒{Y����Γ���cۮ�4w��v;�.j.�O�w��v���m��h��G���=)���ɞ�:h��.��>���[3��굻&g�9��l��ݽ�N�y9��L�/>��nyK�C��y�,�4�ǻ��c��+ٸ�Pa��-$R��u˖�����B�.��f�{`Q8�;��V����L:�C���[��Q59*�q:�٩J�eWm��Ⱦ�E�/vv�oU�.&��;M@��Cn\QP��ef<\k��5�9ܫ�b�Os���}��}��?f~��~��癕�&�jO?	Y��L�L�ןL��싵�Q��=�]Iu	:���i�9�����;8s��J��E]����`�=Z���w�9j����O4`�3%��~��۰3ܝ�2<�*bie@��o���yzh=�ĩ]cnJz��M�^����W�{��٘;�0�3��osٷu7];���yR�W0�S�>c�kP�^߭r�}�kw�gi#g� =��������OP=8l������ׇa�c�z~��݋��z�`���y�Y6��l���=I���z{pz���Y�T��q��#���v�k]|^���;]O�/�Qd��~������<�஬�A۩��4;$�=�XoeԌb�Iko�^t쇽���<���ZRS�ǡ�l��� zk��{����l��ųa�\%�ޟvSh=�>�����~�I���O�+MZ&��o1���К�p��L�Az�s�$��|#��ȷ�J�+}�t�'wz�].���-�8���	���)*f��-���^�2�oru�d��P�5yJ+�L���*v���7�w�|_gԻ�������Lˉ)�+��j�LtF�t��y�ne�}�C����1��vM�r���>�j�����Y>��vs�3�Nz���ϖ���Yo�@} �I=�yV�Σ�z��P�f�I7�N2�v�s�18�bv.�G���H�{U��ɷ[�<��;՞�iʾ�g_�7=�fNy\��;�;�nX�tō��g�\�VA][�tH�u��.K��|]��o���m�9�zd��Ϝ�*g���3؞ml-\���S¶g�:]s[���od�vju���	�˰�cͺX��Wm�}|0snV�	Y�=�O�إ�Y<2;�~������}�&�<}0���7���8+D�������5���V�O��.�4VhG���עW������d�"��a��,l�u'�����E��<�[IM���C=�*m}w���T��|�M�.Lz%{��di.'8=]�ҥ�ߕ�e���$��&�/��\�}�F^�^X�cȮ�l�6R��Cu��j�־�6�tߴݢſ$'�Ե�Zz����S��l^C`;|i��:����65��xZ�.wӱ�1\�=��>�ە��� �*ӣ��;�B������|n�[W>�%w��6�^\�W�o>�z����1�7&=87>϶���վ~T_L9/�Վ�om?M��љ�_�ܞ�<]^���-�7
�w�}�o���oԸ��O9��Q�X�f�WuJu����$�!����:�����2z��K��i{��&畦��в*��].�����Y�c�8o%�e'԰=�Ǣ��3��t�t�j�
��Az���ax�ISf��Պ�zu>��Hlw�f��s�5��@��$����+�y�&��>6fܷ���E�]�����/����O&������;��9� ܗ-�3��=�-WZ�U���������Μe�Υ�	���`͞^޳����u �v�4F���9!΂��ryi�z��b^ d��%�{���{��u;'e�y��	�C��_.|C�ý�`z�Ͷ�����7@g��)�b���S��-�ca��;�:��ۨ���c��Qv�Hg,W��Y�ɽ"�۟^�ϓ�oF�cKD�pJ� ,t�@ǚN�}y'���n�^uo�]��]K��du�p:%_�g.��D��pv�Z�nھ�=���_}��W�V���<�j���}
���{��y�)\��0J;�YmL���.�+�\��/��C���f)q»4	h�&ܬ�xO��{��H=�5��æ>��a�E��`T�~sh�kF���TŇ�!�ʡO'�C L��}R�%}�e)��UY}�lٛ�`\�P2]���uM���󓦇��-fƞ�=���<Q���W��j[�Nyږ�ڵM��.�-����P{{��ǧ �=5⿶	�N���u*�kܕ
�u�,��y�<dnw��{*j���X�N�����7ܦmR(?^�C��Lͼ�U�jΐ�+e-��C�	^�¤�X緳�L��zI��<�T��0\׉"c���x�������ԣy%*�y�z���r��㝵&����T��k�m��I��԰�N�
q�l!Z���|��:3&�گߢ}�3���Y�����^�u�gR
���)�ۭ�);�2����[���q��cU��-�v֔��"p��>�2�.�ε-1��e�[JKa��4�tt*�fчGr���2�9V���k��]Ҕ�j;�f��[ú"&�5eg�g#�߾������l��=��{w�������g�'g
��|{�<�������]<Z5�z5�%a���Sœ�W�cn��'2w�J���;0S;�=�Q!�W�I�O��N2�o+w���u��XtBΊ���������k�s�9Fu�?�>����d��ɒe�λ��)r�\Λ4{|~W*I�_����5��wd�o��	=�_��b͞�TR�U�XX��z�c�\�G�l�䫩�����k�*��23^��P�z��<�֤j.��ㆵ�l ��y:]�;��e�7��<�������2�[�g��\q�'�R�Ve/��*1)�	��Oc�W���<̞#v�7���g���rQ�`�{W�;b��c}V��G�]by���{e��s��f�ૢ�`����A�}�z�ޚl>�V9�Ę����nmX�8�p�L�����x>{p]�lWWW)H)8�����>�}f�/���;��s\9��|��˨��ʸ^Vu�5Q�غŹD��J*���LY���v���ئJ�e���yagt�4��T��^^nqɻ:,��tg<��2=�Wϫ+N��=�b뫵:��(���0N\�r�,>��̓{��5�6���ކ�NP���2�qaA[��b������m*����3o�;%�\{%�����3��A��#�:�|�]�vs�AI��ż��s�b�S0e���H��W��ò֎��n�Ӗi�b�P8�W��0Mk�tY�X;�7t���ug�F{rGn�<�/hvz�U4:2���?��NLo`}Pr*Ss:�1r���A�8�����z��R��5����ܩ���є���V�h�;�Y�h�N�^рzs���9��M��G\Ӑ�{�t.��v����Dl�͑�e���P�]6�f�s��2�"і�����r��TGA�CK\�ZŬE-�xi�e��v�!V��-��*W��M�֭e�b��r��op���rˠx:�To�z��\'T�JHGc�������рb9}۰^GN�`�o�KU�DAV�j�}%�곲XsC�|zR�����N������|����Ew@_VwB��l*i����!9Qv��o<�o�&��SAn>���8x��]8�qɗKB4Z&������^��W���=Ԇ����UD�:�5�TF!��KƜ(��YDl��AX2f�ϱM޵��˘N�2�&�U�Xܸ�dů0�Uk��	�E�cY�3ۭJ!IjZ�|�GH�ͫIp=˸��u�M��O��������8)�,�*�¤Y2���ʇ[/$��آ_f-(�{}w\ژ��h�/�2c WTGn��,=��+;R*1�x��-k:*N���k���a�]��gf��p�5���h�1�'[ݔs�}���Ԧ�[\��x�;�D�=t,�Y�ԇp��G�EJ�L�	�}4����s�9}XWUٷC����[Z�8'�g�1u�d8^�z��G^tڋ��.�j(/\\(d�u������TM�8kx_;�zԬ��D���$+ �w0���9%+���D)9��]�wz�oP|n��/2��y�����4P�)'��ל��}P١���=�8*��}���=��v��4Mp�\��/~1֍�h���M��:��d��Ի���S�T�'#�<+�&h�f
�-��,!ruf�v7�®�#�n�>�O�q-�x�z�n��d�][�����(:[�A]ghTv6k=�fK�2���ۍs��_nS��oA�w�m�r���-kxiYt���Dn���2-�R�rSd����tV��&�g�]�t��oe��v���j�d[[�4{-�Ӈ{��(�R՛�ls�����Z���.�6��u�P����~ �A�5SQAL�RUQM1�%4�DREE%,E5TAđQA�ED�EUCDC@QM4	T��UP�P�IL�5AMQD��4�4��MPUMMPMT4EE5!TRRU14��LLE)LKTL�AM%ESMUL�MTU14EQD�����ULCTUD1TM�RSEPLPQESE-SCE1�L�KR�UAATTCDKI�T��L�HTEKPLSCDCE2ԕRT�PSETTPđP���?_�ֻ����u�#Qe)cp�2�4����\��9�74��<!	f��w��o*܆E�p��G�{����Ik�wU}�}�W����颹�µu�����6�{5��l�]�|c��O~~PO`�n�&SXg��{ai�ɣOJ�D�:�:N������;�����w��̏ct������-�����7�sv�+��{`�Q>����Tz/x-F�Z�~�w�-|�}����7ΰ�zk��_��aV�/�[8=꺇��5�3DV�T�Z�fOk�ٮ�s�`�T]�'"���]\���y+7����gf猦�LNr��[��&�cl`ϳ���wC��5]m�y�OT�����.��&:�%�nZ�7���ބM�e�b���׺�gt���)�6'�s��������{f̜���g����g�2�	{K���Wk�o��BO���w��!҅�t/g�o��^�{��K#��f�L��b{e�^$���H7�,L!}��Ϭ ��@vq���\�%ާ�q�(V�r�F�-sدj�_K�N��GX�LNH�`�HT��U��;�n�p7L�9Y��*w��6��	'�m=���x�o���oSS�i��)u��r��W���e���3�=��&�4����%���؇u��{1�g�������{�qX���ž������=��KΚNu'����\������o��KK���]��8S�x1$���|�N�ׁ=�W]xVi�2׸��1�w�	��v�ȭ�bÁ�X�=BL��K���$ڜ�O�����2+�nc[�U�3f�����q����Kt�]�K9:3(��x�WYZ�zP��\�Ӌ�I����ݲ��hE�#G��T�ژ�%_O^e�n�w�������{<����O���,�S���F�mj��.ʛ|�<��9-���ƣ4����7ݰu���*e���k����+Ϭ'/0s�pz9����au�V�n�C=vў��0���ϑ��ۨ��҅uO��u���~��B��̇ê[�#P�X2��7���k��o6� �NO>^�nm/#*�؞�ɾL�ؑl�Ҋ✄Ϛ��{�|3K�\5-�Cr�&O�G�j�=�����&d!I�OUeNso�1�rUh�w���]���F���C=�y�5�OPy2t�����Ckk7�.�]�7���3����1А{k;r�Ρ��vK��o�A�AjV��Տ��׽���{��}_}�}W�uc~qu~�(�ŕ�f"�͹v^}UE�A�״��s�+ P�u��k�'UK\>k'w�p{���k�QbQ-�ئR�/.��s���9p�zu�*|�M�/wg��_{�������U߃�֟eQ��ݠE��I槀�C�Ǭ��W��vjh�	�XT���,������_I������סIlA��h�/��(8��"�~;��o��tQ�]�w��<�qP�Y%L;����N��Y	�Q�fQFy�x�f��ySb�>�T��Z�-��w��2,����+��JV�`r���.p�'��]Iz��Sz��J�H�WTd���A�UX����y��UBC{�[���
�C��bF6O+w=�q�3���~�s�h���<ʫ����.�~����>�ج�<�V�zc	��/���2���=ih�:
�M��#��[���6k��C��x^_��u1S⼲���Kݣ���R1�1pِ\T��Fǹ�GX^��,�SspY��>��L����|�i���va��4��k���[ ��1�z�nR���{�Ud`����ٸ�_u.�n;Rg6�\�|p��x\�M1aM����Wys�J�z��s��o�m��ƩqR��Wo���+��*;K�l2_8C�ᬾ�oc�V��.� ^�V郬fv:Ӭ������q�Mu���?��S��*p��J8Ϣ�}N5�w*���T��a|�Չ��ǡ�m���}F�*l�o6���iem�iԻ��Ҽ�A�r�شl,0�Z�zܹ|�����͞^�W�ŕ+J�vM_T��{|a'+i����~��sW�A�ڏ�u��񢄱N	���_,M��l��X)qh�=),
��
��m��L�-�u˥��2;���t����-�;��gg*�-O����Yk����f��M6U@x��4�0���P��Z���{Y̒������S�����^R=��l.�:+�"��Q*�\�Z���e�exj=�A<Ҁ�-/|'b0�9��[ޯ8i����Y�Q>r�#eq�eM��\�)>b���S��ך��2��i��ڡ��s͵1B.�L�ذ9���Ѡ8o��� j���y�x��'Ԕ�}J��'�W:�[�S��7�.�%���=s��f?X�7�5�s��@�n��
u�p��P%����P�7�s���K�9����a��-���G:��r��6�KT���XK�Yc���˲Mܾ9�t�&���0�Ay�)Xs�<%g�Pq��Z��d��X��H]��>G�H*i�;4�K&�GW�����ªJUh����a���72K2;+��Y]Y_��w��ڵ����]����}���4�gҰn+�ܭ#�����CY\�k��w�S	���*�>�G�o�g��V�y����WȖ�z�}(C�*����ζ��h��ip����*y��R�i�Ou�O��-��N�	_�rEg���৩g�,��1Y��hNGr��=����27�O=l8�%o��W�'����v!�oK��X���cKL�oL'M�(v�n������F�V�=jC�]J��|�ܮ7�v��ͽ��:�,>�������^k��^:K��TN���JcVr������Q�[O��ǧ�9��5��",__�r��~��e��#���=��0l	�_)���c�|]Y�IQ�L���m��<���.��������v��e�,=C��ݧ��}�&o�ӂq�ՀR�Bӡ��0B�\F� ���$����=��Ǥ�<�;;��jP��zu�]�%ù�e�״� �s�T�~��N���Ge���.�<� �J&�=�Y��T9�|ׄ�Cۂw��+
gB�\�Rwټ:��=����W<�I�)��fr�|�%]�;�����T���K����쇺�hG�z��{��R�|�'@T�r�%��eK{z^,ǽ���wI�,7��'pI��[��o@�5�{�X׺(�b��s�,U���\I���}��UT���x�C�T]��-��ب�您h�fSl¾���{�P�^��q�ȱ;��o޵<W��iM�tZ�m#�>+L�(&e��켪��Q�]2�A�/M�8��~"�y��v]]ֺ�k|GaK��kx�vS$WJ� x��|��x(S2�R����uޗɭ����?�2��-_���8短�D�A��J�.k�P���	�W��(LO���^-������/��4�*Z��C|�	��` �
9��/�{�ZU�z�>�llt�п/0J񏥮^��9���5]���<2P�e]ه��hGb4����X�Z�u�Wa��O��;��V�t���*�9���(���tٙuܽy�?������ƕ.�D�������1�|1�	��v��&$�����kR����x��Y�Wuc�8�뻑�������,�T��v����!��LE�<�ss<i�5t��7��2��Dr�J��]�z�^��(q��Y�,q�VՂ=JE�g�����mЫ�o���t��J3#���>��@�#R�3�t੯*8IV�ے�"�S�^u̗���޲ٳ+:|�]��[9�cHc�.���QZ��ϝ.�q�$k��⻻n��vQ��Vع�� n�k�6�F��-n]4�3��{߇�|��C�bc�ߏj�G�;�����ݎ�q�r(4߀<5�j���鷾�����&���!4����{��<X|`�>�9AYr�;2�v�3�Wm�vu����/���)��N���>�Rj,�q'.���-��5��ɐ��Xo	WR����g���ۘ�3�'��X������_S��M�ޤ[+Ҋ�Few�3�����Ŝ��Ht�z�Gٕhe p��\^ܻ-(�:���E���xT��'���zIRv*��t��Vح���<�*#�--ئJ����g �O�r�]����՝j��|�޺���SE����{׆�:i�U�v�Y%�L�C����otx�9d͞�W�X��QӾ:�)|E�9��|'��,����E��va�k�"M8��Tic=zU�/6�z�1���9GeïD����"�z�ISg��2�T;Q�#�U����!�b�e����6�������:��ﳍ�o��W�}����a�*^9brV�*TZ��g}6�^��Z_�J-�5Z�]�r���p}��dy�Ms>�()�]f��Eq�y���i�����r]��T2F9����t-�ܬ���}�9
��7o|8�su�-ok�R;��^�+k�	AZ�+�}U��w�b����؅F6O﷑fR��I�\5�,s�-�0g���(_Ev���]��X����]����:����f����P�	�(�Lϛ੗qp�8=��4����B���`��|���u�@U:��
�YH�;��l�J�Ye�^���1S�ڒR���+L��з�J3N�T�a>���a2�|���)��-�MB�I��1U�e�9�
���s}����G�N��i�8k�=���q��Wܴ �[C�]�����Xc���D�Ϫ�ԯ%Cc6��_�Hc+lsY�=��id���{|z]�{�iZ+۸1���Cㅭ����|�`3�5�DX{|a'+i����~j\��;W��Pfcc�ջ"�z2\����A��Q~�G�����K�AuPOWx�+�\��b����6�zZn������=\6r�����Sz�����\�҃>#�4P���<o�tҙ'�Ï�b��x��xN���v#.zƘq��gӍ{V��{��,��p6��"9��mz�����c�}B�Fﳗp7��c1n���4�abØ�.��՜��a�]���Z�v�Zik[P1�Z/
��/.�,��Ɩ����_e���`����Ҹ�y�Н�C�Ktj��#�{�7�����\�彻�Yʟ���������q��9���~��ĬE�N�a���}2��^�L��(��Y�h9K��c������}�8���<e�ԇ_��|��OP�(_�9�u�^���ϻ�_���+�2�[��wo+z�QO}@��Z���dHG��c�t�iC<�L�0ҳW��bz�ᑫ���ӔQuOo���P�،��J����di*���Y�;�lh�7�W8�n@P��s�{�{r,�9�?i�Cih1�B/�X,L~���ai-r����_Z�xO�بcGb�ޗ%WX4���ge=k�g�U�N8)�8%v�Q�xM	c�w��O���a.�Y�;���X���{��I+�����$VpEe�a�OR��K'l)��9�G��{�����t�Ln\˾��9e�T���̗�{��؆����*ǜ���Y�	�N�e��T�V?�D�������}��(����Йs��}�J��<e�x)Wl�Y��X�y�J�~�%�@�������w1�쵈����yX����0�#)��!jb{�B�uk�_�#����5_�7��z�$�S�D��tUy*��X6�9R%�㙈]��b�]n�����a�>�!�[�v+�;[�vo.���EάV�kc�M�f�8��A�6wlk�d�0�\��W����j�77y�4����������d�禗ް�X�$���^3�k�K�����Yʋg��w=e�맸�Q��v��m)�\�^����>�_K�#�q�Ԏ��:��t�^'K0�B���r��΂���k�YZY�)���u,x�u?-y.�Yh�aiX=),g�"�2��1����xM�0�n�ȟT:�1*�R���"͂�T-J��Cۓ��YXS9S^�{%��F�K��u[(�<$�)]��w�U���5NJ)��f55�	��#:)�gq���c�՗��6�>�bG�Omj��xY\\He��ت�t�_�߶��'z�3��~wa���N��^�Y��ڷԈ���@�&��k����8��8�U���Y�5�/9E�}o��RK��/�ZO�Qx�e}�x��R A�CZ��K��L�(�48��>]Ufɒ&�����6�*��*�a�F]C�/�K8p��KJ�I��Z.�����}���6�W1�^��'��^nXE����ާ���vUݘ}�zi�}�9:IA��� ��v-��o�Yŷ��X0�X��:��mtD�Gh�Wt0
<V���8v?�i�VU�*�rn��*(�ޝ��:�ލ2aW�v][�q�UgrS�]�L�t�1����[[�7�(�V�j�ؾ���m�tWb�!�f��Eh߄�-Q���&����|8X�1��\rԓFv�T$l���R(�u�M 8��n��^����{���^�
����ni�|W�ptk:���w���TydQpE��7�i��.Hf�1����晪;���!S%�N���dx�pͼk�$�ٲ�7Q�/�a��[�:,��"��u}�K�yCy	YO �j��HMA|2%KY�7v#�������W���k�z�Y���To�1yZˮ����wT�R�Cpk�a��CCn�lբ�[n�*쇛�<�Oh��D�{��W[ϳz����˃2�a+��8n#����Cpuϫ�"v�ujǤ�A�J��BtaS����
<y��RV$�N{E
O]7���Q����[��R�Z��CW+�ȵ���!����T�y\���{gNp��^�e�#�Y1U��%�Soq�wFl���"�t:m+�"���Fc+�xR�VHK�HAE�nf�VB�+e��R��{�+�<S�:wd�jo
��f]%5
 .�v�2L%�:����9m"#/^f��9��Zٌŭ�}�*ˮF-X5~�ia�u����L��a0d�T�r받V�S8��٠�F�[�[og!K�wUz�Lb	�q`�,[��1�nT��@	�:�.���"wn���W�3�X][�H�(�}�Ud��\xӶ�H���:���sz��5�(�G砝x�=5���'��CA�%���tY�λC�@g<��q�ۤ{�[��Y��ݠ���;��O��3�[����[�j}�ϴm�uS�ǒ��d/1l�{E�����\ejSghw;zu���K�,"��Z��T�����. �'X�.���}���"F����e>��d���B�u�ڭ%Y1�	BN����k�_Sx.���A�Y��1Ǟ�\W�͇��{��,����yzl��V�J��DS��jJ�(`�3F��Z��$�� �Q��"'yݤ��d��B�ͫ�����a������xj��}���Fd�P����ܠ�O��y�)8ky>)!��1&����7�Yee���!�MN�� eAN}�vV\�mJw>E��}��Z�]!Z��M�cHܧǸdv���+3NV��M��IK�Smuq�&�5�4�;�cK�j;ox]K�CWE������=;�w;6�y��'Pǆ��}�ӻ�y�Z��T�̘�$=a{��̵�>7��8��`a)I�<֮�!Xov]>����O+�Otx��"xr�Elۢrŧ�
��e��D\I�iv�P�Y;�Z\����K��n���-��'���|�UD��E-QAM%)IERU$�Q@RQQ4�ERPUU3QTST�ER�TD�1%ADI�5JDEIUB��IMQAMETTCT-ECRR��D@�4RR�C�SER��$E%1R4L�UTA4�%E%U-,I@̴���UP5AT1QEB1	@PRDPUATE4�USKHT�PDAT%�5RQT��JTIL�USIM$IMQIAMPUR�AU-%P�$AMQKAEKJ�UT�IITP�T��
(���)p�{�����:���J��l4�gws�-p��9aem(��ػ�����On�a�e7�k'�����]�k}��o��� 9�{�e۸�Z��RӮ�����}�b��0$�J�'.�],q��`1���
�Y����R��ѳҫP��۷�f��+��*Ö:�>����Zק�8�Z�K[>&T�p��$;,� {h^w¬�B�S>��Ə����\�I�E��w˱t^h�SŠ
د�9��V���Z�^ՙR���#Ԥ_^���}녭��c_�KS��A�Wϧx�=tٜX��vs���^���P�\��&Wv_��t2'ٷ|#Za��3>�s����χ��FԬ>A���e�/6�m�� n�^�m`s���υT-+
���;Ԛ���W�9����B5���!�[�ջ�4&����I�3LZm�U�T�}}P�}�E�����V"���Է�������u{�����✽��J��8Nx�Z���ҟ�)/q&�zh?,�"♰A��-Wo�
��E�X(��Նl��G�a�8�I���Kb�)W�N�9R����⠾�#���z��Z]1[�Y�kl�>�#S��W�q�;�Y��>Z�)S�{Xt��7�����}OM;�S H���� �}��;d���Y�6kl���A]]]��ϭZ��bP�[��U8j�M�(�ey�إ@���գ�Tӳ?}���Uk����߾�h̛|h𹽞�V���Ϲ�B��YA|N��T�z��g����׆>�+3��Y��Tb�K�͡=/�}=z��D8:D���Z��_���ߣ���D(dY
�g-Ջ�ïD����"�z�K�;��~����x�ר����S�Ѿ����얌Լ��U���w!��+��j�(*d�����)Z���X��^ɟ�R=��>����[�y`'�#l�墓K��,u屆	y�^����k[��N��}�r֨g)ПoYfO%S9�L��<ʫ����E?_2�e�s�ok�cVpnWm ���6��2M��I�b�)b�V�X�P�}w���<�f}t��
b�N)�o�F�q�0�~KGK$T��R�Xj�ն_�;����u݄���K��g�4���ږ~Ռ�R�v���Ҏ���q�����B�z,K�{��즦�S3Ԕ�ɣn�O��>&'=�mT�x�:��4�]����c$�r 2�sH�y�Z�N2k�L��g�����M���z����j��-Ս�əl_����Q%to&cV��W�2uF������N����wu��,wuL�͘���� 3/�U�yoKxUկ��Ҋ�����W ��L�-��P��9��L僿��W����ns�۸;������8��^��񄕩����d_3�AO�EYw����{���]�p��F��E�+E_�j`/�����N$w禤I��p�<�)��=~��]ds����Bl7��/w>���XM~䟩P��JP��6Iy�B�����J��Ͻ����˞��u;�Vyy�#�;�8h���o�#d�[��6b�Vz����	�o���yXߧ�5ߜ4ˏ.�2�%��2�^�����~��j�a\|m!���vK�,���i�P�9�ژ�}3b����x�'6c�V��hO�Y�U�	�>��|h;C��|ꡚ�L�<_J�]�9�=�J�������i�dY��0�@��H�V)�.�]����̀;w8(9yl�{>��9�������;+�{΄���P��P���B��\�\�y�o�l�<(X^��yb{�je�
Z^��wE��b��h�
z�Jc^lW���:�[e��q�yb�N�|�׸�u|����sF�b���y. ח[����5ƙ��h���&�s��8���A\ϋ�b]�M[T�&��\pD�;2�k�!=�[Kw����5l��uH�kYƘ�{����終:��X���u-ɏ����Ч�yc\��Z����d�&O�ܑY��\�.�O��1Y�8��޽����~��AZ�:.�]8���y�}]�g��Ƥ�
�_��ñ �^��%����`ݱ�׳c`�1�A�Ct4;7�E�b^ُ!��ZE�����ih���몋�ߞJ��$� K6��(r�J�|V��b���a�#X$!�����ܶ�V���܏g����3���/{�@����3�}[K"G������E���]K�{�v����鮶3˵(/��`�`ob��^s�ݵ�?�`6��O��ȫ�>낖�F��J�R�g9�L�l�i��V�eӹ��<=:ޮ�P�]#ŭ5�S|pL�I[oz���|b�J��Z�PĻ�4�������5�o�hUy>����_A�4��eu�y���)j6
�"�U\f]QuO�����Ԣ�'�e�C�{Əf*4����������+�fB�y#�"6�:\Y�̿�ݗ�C�Μ�q�L�>��N\e�R�%d	���3/}����ج>g;u��x����v�m���%?�t��{�^�Oe;C8�iꣾ��I6T́�5�p�]�č�`�V�s�P�t�)p��u�e^hP�y�������cD�ۭ�H�!����!JrG��;������G���7ґ������O&^Цe�����`R�?Y��l�=��`���g�ˋB����������	�DwCZ���?eg\5���m�Y-ݪG�D$���Y���Vf�eKZa����'�w � Q�X������H���S7iy�껪�{M3�t�g70#c�dA�+����Vx`�!�Wva�>���
4s�^��
��N"0�/���X���Ir��V�gJ$����V��y7[]4��ݽǼ	�6ѳ��PWf�Zco���O�|�=�P�����n�k=��I�&�^���\�!��˴Ǝ�(��pNס�s1�"%R���Ԧo���<di�;�W���$\�~kåw)�Ν�a�ﺍ�yև�/�X�k�<�{���Bgu�y^���,Z'.Ϳ�{�����l*�c��\iܪ�7��W�v�:�����3��cݾ����B���r���N��<Y�)����ڭ��zl���5x�U���y�7S�G��mDX�m-V^a�9�{g�o+�M[�4z@d;l�͉t�Y���:���.(���q�"z��\�^h}�(��H�	;6,��2�8���[�K����w���q�Py�k�׷%��6������K�`nN�z��]T:�@�rĚ�;��b�́���jq�����)���=�d�O�t��^
�l�=��	'D���ZE�����W�S��o��C��k��۵��G���i�\}��^�L@�Ij[V�8�����)/q!�]f��T�X�de�oE�ܯ	Y"I7�<+fs��{WG�a�G$��m-�e*��:\"�S�ؐ�Y��έ�h>����}��|*����ɡ��,;�U���hl��Y��z�={�.�ۂ�0͏�yN�0S��9p���"��m\Ϝk��������^�= I���T�n�'�7�!�P�A�Y�ub�p늳�7�T/V	*b���p�L�����wޚ���x�����.${�%�µB�b���:��W�K�}��w��Z�LL�d5��V5���w,w�p�I/}ґ�,�q��.�c�[`���<�<������ry�N����葠ؒ���#��>h��<ʪ�z4�]R)��{��!�6d�z�+��W��s���+�<�)��T��7���+�Rt����j�M��n,;^��m1���,��v+*y�W�U n��~���U�V_,JZ��l�7�N�d9�0���u�w6aXqj�k�j���[�z�m��c����AӮ���	��h�d��8Ğ���^A�
�+�Υ�"A�w���=�Z�ׯ�=1ڸ��^+�\��ǈ�az�t�EM��g���o�:^�C���:�O^���Z/��Ʀ%^N�CՍT�߇z��.'�5�w*� �c�����Q��]e�z�4dκ-��z*�Ԭd�lf��k�Hc�lsX���|�M*�˪t񙝛���_�Ĭ��<�\�[a��)+\�9���x�]�G�`�˸vܺ�+���Ml���l��N��w�F��eP�|UYh�/Bє��}N$M)�������]���m�Q�����5Rm���z/w+-q�p*����H���?	{w�}$oP������SJ�{���˞�������h���g4F��"8/���͗�Cb�(��_?vS�ZED��W}v&}R�!晞�،99�+{���^G��N��I���n!��Y���,�@��C����jWb�˩��h�Cy9�ژ�cpZUPn��Sk�#u�h��h�^5R������'.�%d�=#k�BW�e�0m4�WV`=^������<��h<�z�=k���o��}�u�ߗ�������9[����+9�N��^G�0�@��n]��W���_i��ÜI����u~�W���+�f5�PL����C��J�LT���i�&���j��J�r7��]�;�؅�jZ߄���hw"4�K��8߆�TdZN ��D��i`�Bgd��᜼�k��\5�K��Ж��&|�i!Z�rV)�y��<k9{ك)�h����Ϥ��X=���
b���ma�OQ�%v�]��P��z�;��]y/f.�9�J$�O؞�[����ʉ�'�B�P]*��҉��XlÑ��G�0�W�����v0	��V�n՝�����o|k�zX԰>��_��13����������f��N ����1��G��s�>�L�ͻ�{6���A��}��t���&��\�;�~���c���Be�G��ҵ�ǥ���1>#Ԛ�!x1'��(j�S��l��t�{�b���lq�8�Lvi�x�����L�JC����hP(4�[�XX0�]��g
s0�å��`��unJ�����GL��E-�8q���`IQM��.�t����u���b�{�����pU-��v5�Þp�Ubѫ�>����ٙ w��m��X�Û�$���3w�b�Λ���YVDiemc|�;�]���c�5hq�{ۇ\ cA�0���ن�%e�M�͙��Ї�u3�jN�#���vN�u���)���L����t�r��Ա�/�����ȣ#�җ�'[h�-�1��Ƒ�8���P� �(u�bUޤ�OQ7��nW\[�䫧�}�jh̏���5���gX��a`tu!���U��H�uW}�����au6�*>� ����W7��':L�A�؄X�X�k�iqqg�3Q{T;<��V��-��n8��?p�����μ�-��bET�"��������}t�z'�'�2뵜/d����H{�N�ɩZx�������Ǖ֘3�	r�!�֥b�5���u�V��[{�v?��M(l?K\�7,k𕙧�R֞�(o��&\;�K������Ź;�r%AK�KV�K,#�u�^ӟ^��o�r����:VD��z�g�	BRg�-U�'+�=)����b�X$xi��(v]e�{׷��u���XIw�T!_�f0w���3B��.�ǞuŞm]^�,z�Ƽ'Z6}>�@T
��~�|/���`�`͗d�O݅=��h�����c|9z�t��&)��%���i���Mj���ȴ[g	��Ǒ��5��!oT�����3؅��`jq�m�t����έ���'����A���[o_�E�kҷ ���R3�w[Y5��\�ͥ<<��L�>;�,t}��Ӭ�Q�J��v.M��퍱}h���P���R�&8+�LL��yǼ�~߷�n��N�5��>FCǬ�	�w	"��zW��]�#ׂ�)b�X^՘*X�|�׌^����N,�u}�~����r=�T�p~�z�~���ώ8������u��G�Ïg*�<9�}Ur�#;6��u�w-\,j��/��<F���N��:����>Q1�q��T���θ=[͈�n�Ԟ�Vw*�iઇR��P���u��}\��U���{qv�qF���5�^O{�N�L=Sg
Ƞpn�bX_$�yyt�x ��Dw+��6����R�`!�٧0��,b��^�/D&}TTԶ,���V��v;��q!�{�;S�7M�Q���#�N��E�9��C9׏��[�#��*#�$��l%�L�\Y��m��������(pO�_3�"������2hBS�l��֣�����6hR�²��r���v�{��צen����E^QW)�Br�ת^��<�<>������Ͻ-� ��g5�ԗ�R��׻s���H���L(���Ν�;tJ�ci�&�C�y���!��O,�Y�vÆQ}S�}~KM�|s��|*i��f���+6��1�f⩺-�ۖ�m�9`�r�5Y�("nF�p6�F�\x^�͝��%٬�8X�*ţ��y��j;
]ݵjX�M��>#+*��+�������vó��$��I6E�܋R���vWM<�S"X�F��;-`=υe��L6yN����{+Wfȃ�jnw.*���:C���l;��R�3M*���=Ӏ�c.�T~3%�9X}�/Kμ�vL���5����l�f6.����j(����A	����=�igL-͝��c����`��3��ks�Y����k]�uz���k�F����ܾJ
�v��l�EM��qܮ o�����It&��o�u�ٹ���Ҿ�/sS��ۤ����+�)M��u��=x�,�㙣BZ3ԗk0rX,����������܊Wӣi���bF����>�u �r��ߟ1j%���+�u�Ze�'������S�%�E�A�ŋ�wR�Q�S]DQ��ꩍ��Va��ɹ�:��4�!�B�+��̼�d�������ޖ3��4`v�lJ�r��4�v@� /��H�.����Z��:�Ǚ�k'A����{�@R;uJ�JMK�WgWq�4��ɼ�rL�'[+�u����%��)�+Tg�'9�P��f��������Z=��&&8Å��{�a�=e�J�Cݐ��\���s��2� Z9J�W���e���$�f���]�yw��x��A�u�Y|����'�oSSIǖ;��>N��{�G��Q�˽޾��5�u�()�)lǺW���KV�ݑ�g�j���:͠�V-'{��k�:_.��r*�vyiD`={̆��w�y9]�i�����!\��ҷ#�9p`�:�}Y�N���_�|�+S��-�/�Я��z�j�uT�d�Qs��9ekV�M2�+��.��#����:�(�}�﫶��G)O�0$8{5^>20�R1�]E^��T�	��v[��m��wKC�#[2=̦5A]׷B=����1���&�T��J�c��#��p�.��Z�bY�p�ӱ�
���	\+f�����IS:P�oo���7,���ۮ�ھ�n�%kt�В{��v��[&���f���w���<��L�2< ���yӅ�O^Є��*¬K<֜�BL�.�U��N��gs��;;���;�rX��<F���[��U��ڕ�N��ms�W�.կǅ�T�Z���%�(�O%\�G��\`�#�CY[4#�iܺuu����u��0Y}]��Ʉ+s�cR�	d8r>�.�j.�"��ѣ:xMQ���hg���I>��tDV�hWRv⼈�V��Y�m�5�ΖJҥR�RE4�% D�MD��PR����RRRQ0�4UU@QT!CSKU%QT�#ACTPACAE+B�!E	SR�!M-P��HPUCABҕLKAT�4��QE%5AC@R4�	LILER�T)@R�%�A@L4ҥ �4� PPJ�E,M"PP�-%4%40�QB�D�	UCDMPTBR� Д-�U%R%-%R)@P�-(TE1*}�.HdQ@����}�%q�a���\6���'3^�ܽ�2��M�����ޜm����VI���e8�Z���uX��Jv"m��/�@���dD �p��ƕw����s��h\�{�~���z�J��n%�qѼ^����k�J\=�җ%b��Ԭ�v�Ca𧻓VpA��*d�������쮩<�uOE�t�h��NY����$�y`�\i4�k�,X�Yla�wkfz��˻��vkc7i!�^;ƫ���$h7%/+�قx?ZJ����Tȳ�K�9a�u-B��-M���\`�LŀoK����j��6�6#�}&U���Z�>��
ވצ���{e��K�r��n�*�h[Y����x�iV�ѿ8��,/R�D�����Bǋ�2g7:v]1"�Wa�z�-v�d��KO��]n�c��y�N�p'�q>q��f�Μ�=�҄�6�:�xX��E���쭻�"\0�U<���BS�����[�}��U�: .�3���rٛ��f���}=�Fߖ0���+\�9���Fv-D�	��J�y�nBy��^̩��j��/�y��Հȯ$}Jz��V2�%@���䯛bƞ+=;4���SE�3���Xh�|�moR��93�Iv��o�n��Sdո�k8T�ݥo{�*Ek��\�m[y�ݘ9��7:���9A}��ovg=�Y\�c�s�*�.%ge]�g�q��Bq�r�v����l��NW"ֶ�g0�ܑ�+y(&�"�s�O�M��)��;�VZ�,-4�:��:pR�����X��A�u�w�D��\�#���D���x}U�Ս���dw�
^ǓAOJ��-��{�v	>#I#��T6
w�Y�L͝h��NyG&V����L��7�iacIC��T�eM�s��p�:��.G��!���u Ԯ�ປOV�ڡ��sʹ��^��}�+ξ^l��"��|�p�H)rWT�k>����t�ϓ�f�ku��.]�{wެ~NquX�{ᙪa���i����>R�vu�Ao"4�W�+�7)��!�vk�o�+۞�̏)-I�^�r�yl��j히JZ2�%`�1��B��k��N��$����Q���lI\Ǒ�2��8"���k�3�Ȫ�'��#�J�Ի"U�^~dA���jO6g�
^���{���>�����}{Y��\Fgs����"��Ee�n
z�J'�!�C����&+�x�ٞ^�`�s�Cm�f,r���y���C���gϠ�W�����ޮ�.c�k�z��H�3X��x+i֭�)=�79��7Q���/juK.�TϜ������Cf6^�*�=ݍs4��S�K�M�3r�t1p��B�E%�Y8�c�r�ֱs�g�f����2��Ê��):.���EéOg"&�����\fv�03�����b*z�6����pLo������T�x�ଓ�g��]�mt�zz�-��]B���J������V�X���������(Ox������Tc4w>X��tHS����&w-�[���Ӏo�idH����	ю:��tGe-~ꃇ�;�6��m3�g5��!���մ�l��GN}�	��17݉��yn���p�{��^V(0B�����L����,
w9Bԡ�&�yk�p類ރ�po��m�92s'���2�mDP�<1C�&b]�k~{��`��R��:ux���*�-v��nd�J�J�n��l��tHI:&|��i=�����\�0��׃��(���4z��ݙ{x��<'�\��c�R�:G��
��Ϩ&f:���ʄSX`ؽ�F]ve��2�ҟ�SY��D4�9�M�d�kք.�}:�U s�M-�e��)��������e1,���y%S��S���;�`�����������,3�	bP ��jT$�7�V}J��ôtG)�6��ogV���Y�K^��M`�\���4�ts.�=�mC���u��p M�N%�\q�骖ms�xf�oF]�t㘷]��]�'G������D2W�=��~$����Q�E%��4�kd��9���ܪݗ�R���^'���gLnX��Y�{�T���C|�}2�ܗ�%��츰P�}^�j�u�3r  �Y�X*��<��U�S�|����z�[/��8R�/�ZC}[���H��.x�ů���9 �u�
�xV���i�ٹ����gt���%B޴�aU�?We���R���$��Q�$�tّ�	֍�M@Tp�mMۃn��3ޙGMU�~o��2���uRS��*�yWPU%�8K��0���C��=����s���{��qS�yZ��1��3v�#��<c�d�:����zWE��G���}k�a{V��OM]���s�䜃��j�V�-�=����x�:pyǈ�ޞ���#�=�����W��Ja�OE���.Uz,R������!�A��٘)����/�������+�r���F/^�ݓU��M�j�Bc'�[>�xa.z�*z��:�G�������w��|
�u�#U��x��s7y���N��UOO
��(qz|�ē�e(���� -vGp5�ԃ#ԩW��b:�+�D}�))m�yl���8�!YJշ+zm��w-�xQ}���р"��n�'%��sE=���Ĕ�0�l�,g�.J��[��9F�����P��o�y�Q�����*�hjN�"����]J�{5ջ�Kba�����z�S��ib�<�B3)�v�L�/}� Z��j[
��\^���J�Ebs����[Yoy��R�$G�A�MH���
ϔ3�x�l��?+ƒih6إ�ܘ8��Eu|�ַv�R��O,�9p�zu�/�s��׆���V��G�RK����}��]�la	f.�$��L讨ϏEp��t��������k��ks56RGn���=N�}w��հ V�M�u����-�<�t�ڇ@j٧R��ՏGh�h�1�p��=�4A�R��XD*�|���.���.��X֝���B���s��"��ޗk7tn���t�h�����z�%o�fR��I�\4!c�]��ou:���tq�)�VJ:���,
��,�'����`]G�W/C�.̬�B��;�eF3abx��a���9���}0��B4M�)�lGH���ׂ�
��szt�N�&�q���ud�k��4,fи�_�ء�W>�q�9�gK$X�G�t�c�?{p�#Wy�c�5��N�²������f�<y�K��'GN�kҦ�k}d��jF�;���e6����
���%m��W&o�	�Pmf��㛍ގ��	Դ��cq墙�:���� 1R&q�s�uA5��9��k���mb�3��z,����ͫI��W��a��V�c�nX�X\O����r�VVfg��W:��.4:�Z\���j�Y���J�J�5@tW�Haui�czʳX���_��ۯSڒ�^����T;�jv=y`���k��d2�,�`P��/�`�{��q��3���ę�z������5.j��j�I|{�7������ц^�Z8iWwѾ#~2�dlb}��9��R%�n';�j��`��^�/w2��:Pf��3�|]�1ik|^�����@\�Q�Gc���}��~�̵ٜ�P(mF�-�[fK�G²hy �2��<����\D����a�|�3};��Nx��Y���#yVtz���שz���\��Qg�D��#�Wm8����4&wa�c�;
�# ����X�#�ogZ�?W��<�ذ9���t��)rV*��g�"����:mP����ύ�}�Ux��l�=xw:���Ӆ���離bs�1`��a��ց��N�9ϛ����DA���k��9�2D���6F኉�`�N���T�}����w�5�uӕ���l,F���f����n���(^�C涴Q�g��W�*ն�ƻ��ċ,Fzk��ՖDy��*�����W*���X��P�Tr��}c8��:E�c�%Nۉq��,w��x5v�xJ��*r�X�)$5��::�r�ui���V��Krw�Ga�7c]Z�tO�oeg���LP�U4N�>G%v�]��$��q�����$��b�����a�fߢ��#0w<	XrEg>���������{�<�9ޮ�=�[��^�4J�!�z��#᷊�q3fKȟ-�8oK��X�����=Zn��/6�w2��a�Zug<'M�;��*u�Cl̯E��o��U1�(oeqBF�jr�:VpsӍ��q�Gմ�)ǀ+ظ@=fկ�q�x8�~�ӥ�ǥ��X�8_Y����r���4`��z#�/��c�d{>{q�/{�@����쵏�X%��PSB{w���s�Q�O�����S�`��f
s0��t���w;�⇵�3|���k��[� �X3&�|3wgG���R�B9]U��8;M2�|+K2��s�-J{ӭ��+'�TyBd�:�z�����R���X=>K��P�w�f%C�I���"͗:�W�o���ڊ{.ڤ���-v�@��G�u��ݗm�ul[]J�2`^>t=Nf�#έy/�$�J�X`us˶d�wۙD�Gs����51m���q"8�\�k��Zuz�tW[���wH�Y��J�s��3{K�A*a�nk}M�gg��^����`�L~�>��g¼i��r �1U\e$Gz��5����=T߽�W��zt�BQ�眬Ϛ����A���V;%��ZG�����(&e�.w��G��{��uU^��٨{V�^UCX"��y�O�o�r*��D�NP��<ȴ&����*��ܟj5��s*�}Nߗh�|l�X||��8���Xg��lҖ����F���S���()g��^SJ~v�`nX�ߏsU1q���reý���E3-r/��ܽZOB�������=Y�c�-r���D*���k�Х�b����B{A��� t,X�M��l=C�l-�<&�ʾRm�'� ,��0K� ��S�˼�"�÷3���c�N�.�����A\5��k�����Z��o�[�Y	�]s�Q[�	�Νt���Ab��5䷥W;ٖs��^S�9���*pwf��9���Jl�'����u<\|3v��0����j��D�O�l9��gz��,�y�i� ��u���Y�v#ˢ�iZQ�o�9�d�W�egeIn�C�c˾u�y�I��a98j���/�nu1EX����s8Gc�l%���F��v��8-�u�ԂC*�GR�-�_?v^3�F����iܖ�9���E��RU�LNcs�9�[�ܙ���}�vӽ���j�`qg�=����~-�h��q�9���n�i�˦��^V2���Y~s�;`��xZX���,j��ȡ}v���lPV�3�;��Y��m��C%��|���Ԙ��ȸ���z��[aN�,�y��X&�C�X�(_ ��z�Qg��qa;uެ�ԧ]8_����c�oW�j����cp�x��$�yyoW��|{�m�Qv_]�z�G����W�S����l	�jb/D&U�%�lY]V^R�u�ۻ+����=��-K�ą4�~OR/�9�a��o,���ϊ�U��r �[s9ny�ק�-�p
U�3뮵
����Νh�&�57��t:վ����~Abّ�N�#����>I�2���_Zer�r��Pga�.�͠�8��g��B��ѵ���'����l���$�������A��9n�s�u�i��G�T==���3<{��G�d"��_�Âx�4:R�du/�О�-i�y�׷0H����tA�	�T�f�6&�|5�<+�
�d/Z��=u��2���:���wK�6�6/="�������g=�H��Y{%]r.T9��i>�F�ꖓ]de6e,܆X�"Q����[D������8�8�`����3�؈p������O����5v<rJV�`r��D�A��7��#Y0�'���噡M~ۨ�YԻ�)�2w!���5Y+�!��T�q<J^W'�yI(X=�
oa��E{S~��c�v���Z)�������tU��	��h��K���Hשmj������u���kݻF����[�3��y���ye�z/���:��B'����.�S�Ů���:7XشH���,��X��m^��}=W�Uz�[����Ze^���o��j����!<�39��p`Ч^��hz}���_%�	O/	�z�;X+����K7�D�ᵑWiΉ!\��f�q�W�Pn��v-����p�1�r�\��e8��\222n{�m�9Ϡ��G:��L��f}N^�Թ���&2K��y��`!�^W�/Z�6��*L�^�n��@s�����D�|�ԉM�Asl8�6���Sz�����/�;b���v�߱���{|TǨU���*3��oMC7ӱs�4���e�8׵P�1H�G��GEVh&����t���d�f��q7�tsq�������x��:���#���{�Z35czy5�k,���#<:xx�d��fh}��q	]�#��A0�Z�*l��[�մ�{�ƽ�+�}��B>��w!��=��kD���9��C��*u�_i�)AB���R��-��|C���m��.��ِn�н T�n�-qp�����7n���H
ޓ��$l�E��(�t'z_Q���rۜ�T�ձU�b�Ю�/vt�n�=s��Hug0��%l���Z��xXa�2m��u�F+���1�R+�#g`F����q�y�̮Y��]WNޝ:�q�������>:��V�n༝���!�h��%:7��K�YXP}��8�[n,�o��ײLբ^�<j���c�,`Κ�:1�ӆ�@@&Rp�GIV�9GyN�tޡ[����x
�`�ᏄokY[�FfV�.�R�QSu�6o{��:�ͺ։��:�w ��N�y�H�j�沁��l�䑽������Q��O:���r>;Z��`�/�'��F�6����po^������������[5u;X�Y���:{:��ʬ���3��eu����`1m�VIǦ[��7��I�Z�co\y�����F��V�O����v���{P��m�G"��j�7�X�؁���Z7�Lܼ�+����j�����)5��CK)bi�ޱ����]Ns]G�b�%L'H�u�[�y+�l��%���YO��}}2�V�<�,��O���4jcKF���o.��A/UK|&�7O�Z�32Y���-������#k�:<5�;
�ӽq�f��}|9CM_;Cn�=�1�Ys�}�z*��v^[�S	�h��t����j5�{Y��`���>ql�C�i>�M9�U�XN�Nӽ�vis[s6��V�R5F�-�֋����)C�����S�˦\�wV��-��1[�2NH��Q֯��#��>Ki~ ��c�k՜���ӛYF���l>��^#j17��Nܰ��wO�Gr��B��&�w}���2)�����-[t�a
�
�n�7��;�YR�5��LD���³chr���ذ�]kWoI��$�t�B� �y-4��x��4�Q�q[63е�[�w7V!\nZ�WԦ�P��Іn�U�yw�XӼ<'��W�B�����q�maV���%����/x=Ε΄�i�m0����K�8՚ �G�˵XVa���ئk�)v���q{sw���WT����>m}�^ԭ��v�-�Zk{;owt���Z��\����6%ۮ�(t�����������=�	��n��
U�_D�^�Z v+��Z��2��z���u��$�ʈ�Uq�� �v[|�;��4����o��릤��������*�>]ɹ�'w2�Bﻠ��O������|�%)��+E#e�UP�RRP�@Y�@��P�9.E4@U	CSI�#K&@���d�S��E�@ҁFAHR�@�d�CL��9 d
�@�NK��E%R�-CMPP�d�"�DC�����1R�,JPP6bE
dلKCH�HQBRd �J�4��f`#CU	T�CBR��R4�������y��5��7j�r�ݜ�Ǟ�bR9�B����WJ�W��bVz]��c�j����͖T���f���I×\��{x����FGB���\�[ſ7[=&��^�a����ޚ�db�����'l��7������8{腁9K����	q~�b�����z�Թ�z)����G��Қ�z�T#.]���C>�Hr�%b���PN�e��XՋ���T�B�7�N�)�ˁ�Ry^0����'�bpL����,7����H�V)�.��l�w�K��'U���0��@�O.%�tY˝�����z!)h<ʄ\�&?ZHW)���mt������T�;�����P��{+���)��EV�.��>��k�vCn{/���K�y�LJ�� xMߥdCk�zwz�k^��.���������Hp�.�=��]X̴���ڠc�qםji���V������!\�� �)�l��'ճ<�K�
=�� f&u`��;ݖp*u�Cl���p����7�28��O`8�/t�^kA�+H��X�9m,�i�}�����-b=(�-�K��s�z��pTk2�1-�(��w�	��w�xFb1�5�:�77�:���DV�VU��Vj�)!�� k����=����*
C���k�m�����6���d�fH2��!7 ^PFu�o��-ʶ�[�4�5h��׷�YM�N�S�uSݴ=�G���#ɬ�5���萧��8rE��J�X�V���Y��2
�=�q��5�T
��܊�Ϋ0>��U���s0��t��GSv��P��,N�@�3���U�|�/#��YKm���A�l�}�i���gS��|�XV%J�mw�o�����x-�ֿ|�#���`��z"�E:]J����Uj�Á�E���A8���պn�H\�S+�m;�{`�흘�,W�2y.G�q�JIh��i
֗h7�^S>���D�ms#~c��ORi�mف�y�x	��"��V;%��'H�W
	��g�{��;d��֭���xu!ք
K�k~��E^��~�x�]9Sl��$h^�'(_Cf�;�>q��ݾt��4X��-a���Y�\�:���}}&������:5�b=�N�Y�9;tT},��n�Ԭ
N)��CآP����5�J��̩kOE�,o����9�u�3<��~P��VK8
��u��|�{M3c�-r����Ҳ ���=�b��[K9���S��gl�w^���\�� Tz�.�r�ߪ�,���Ք�	˟�����v2�k�up�*�i�1]06ph�� u�ֹ."UJ�z�S��j�=��}o;+��M��цR-��緸b�j�;��Ɩ�ul]����GF�,��&4�-S�{�Γ��AVxa�va�)ƞ�r׷2�R,��&߁��Ƈw��Z��w�J}������0q�-hr���=�u�g�P6�p�5y����{��Y1Jk8l���`͗d�v�b�9a�bJ�Z��J:�w�,�~��0u�^ˆW�;��^�/�=����Y�������b�!��1ݳ�Z�� E�2ޕ�һ�}���]��������Ǖ&`ay���o�`�R�_����X[u�8<��pzz����:��٘��6�c���k���ʬ�*��)CV��}v��Cb�/m��KXT����K��Γ[�k�zϵA��#](��;2�fa�]�g���	��W����I��k�	+�t�=�С^�"��}\��1�u;z�cP�{&B7+��(�8/�}wz'�@n\V���w{�����.�LΤu��m(���fWyy��ڠz!2��-Kb�]VZ�Ew�&-�Bҹ�v���Z=Ho��BG`4�k�E㝂�C9׏��[�#��#��o�n�j�6�
�ꕀ�s�'���{���L�*��h�-�RS����j��78\���괢��f�ll���NV�6`�"qaV闠5���g{���/h?��.�r��W>P)��3�:��N�Ke�y�f�]f���<���9���>�U���.�T���Ӵ�T��\�Fwӭy78��s{<o���T�gGnɽe=�}����^�;��R����}KW���Ev�R���hff��H�3|�[�W��!���V �u�y�;�W�h;Y�u`\�k���!^x�V��S�V{��9P�M�ks��C���'�#C�.J�S#�_��v�O0=s���\���=q���5��TɁ��ǎ	)Z��	�V
�ORJ��"6̥増;giv_h��~�K�s��8h����:��eR\��]�q����,�'��޲LN�㦽������FN�yx4�Z)��:ӂyf��*��ՇB4M�)�o���eh�кĿ1�Ƀ�*4Y��s����CS�t��;~1�vv�B��ȃ�OWt_[>^,����6t��_FrSU��P�R%��-�s���z��
�(��Z@�]�#���*�_��ZO�5�t���z,4����V���g��}1�P�?��a�nV��[vW=/8(�m�)Va�I�J_�w��Jԫ"�%b��&KU������;�����ᶨ�}#"<����O˒=Z73��d)Jb����g�c��y��|����0�l(��h���5���y��dov��I����9]�;���	���*�������:oV��)+������zI^H�Cv��Q3=Q��m�d����r�?5.j�A�ڮJӼ�qjψdW�~uB{Eyѿ97�{�6�x��ŀ�_P��!#�=5"X&�"�s�O�M��
���a�[�»����=*����� PІ�#�;�Cf]�x���oMC7ӱbzƘp:������Ϡ�b�f>�v��H_#+���DpTt^�Ep��҉V��夯���c�� �a���^e�8.��+s��yQ��!�^G��},�4�.F�\a�C��ԃ���ZX��_�����c{��P����m�OT#.]���j�e$�j]T�k)Q�WcWu玶[[9S7����m�~��zp����'�breLX%�X�8*�� ��{j{���Xr��),��K o���@nE���z���m��{҄����P������32���x�N��O$�����~JN�����^�TcS/"�h�
|�]�7�N�"z޳t���nGm�cĚ�*�<����6�w���q������X5'����8�5ܜ�f�8��YM�����<h���Vkso���]����˄�`�� r�NLS��X�Jj�فl�)0<��_8�>����n=�i�lV�[ U�j��g���\ _?bp���^��D�S�1ݽ�?Z�k�ޥ�ڞ���`pVa;��(��C^u�m�8lş8�:��x�j�~=��1�l2�y+�⵮�<�I�*zL`�3:�t�t��le*V�����ދ���� Ϝ��"�`ߙ�3oq@z/�>�����9{�ڵ��.5���njV�ߥ�L��ڥ�?WCk��z���,�X:֦'�萧��8�{t�^Lw��f��ي	p/+��@ߥ��p�T�B<���c:��p�S�V�3����t���w;�{��o�M�Y$gc�����A;�ze��{Bxb8�3ʴ�A����)��if];������UYlz�-
R2N�Υ��{�ֽ�E��+Lߪ��E#�����P�Ri��P������3���a�7��R<`>r���qo�k�jk|8;b�#�t��K����W����ڸ=zX:ʟ7au6�*>�!���[�p���:U.Z�#��\\V>�(yu��������x�;���Uv8�^>��Y�b�4��J��nqZo���Vr�.3ݒzf�-���i���66�}x���Y6����e�3��;Y��u�$u9)�ݕ�ΜΙ�*�d�7��C��qf�KZ��l5�f�h�s��jz�vM�Z�c3��a�$3�%]/��闟CX"��1~Qf��"*m�$�@�o�Ǟ&��~��s*��=�x��R���:*��a�Z�?�f�,]u��'E���A�R����w������u:u]Ƶ+R��nTJ���偹c_�fi�|�L\H�uҲr�^��薏nod[V/�k�8p�5��`���˰�{Jg{��/7��ŔƼ��ݺkeV���Q��C��30���H�,��t��u�H�֭0��w\�~��S��������B)˶�(���N��̺��yL�u0�zט�74��������f�+Z����7�Օ8T�]ؠix4|�����"U8{�0��y�s}ó��� 
>:�qCEӵ��\�s�������a5�P�4	2ޕ�Wr�W���j��)�����+=���:̠�'9և��Z>����{�������<GMלvw?^�W���f�u�ewg]h����)�*ӑ�
O[�F����^[&�+s�kC�˳�8�̬���O�.`;ucD@K�5�l�e��y�[wKI�ˢ8e��ڃ:�o!���� �csCy�M�P�$��I�P�"���n��=s!3�y:ڕ5�-��U����r	wgvmH{ۃ/��3��{1�M���yǄ�a��r��҉�ó/`6ݻS*�ԯ �W�<z�#B\)��0��Z��Myu}ڠ�3!�T��F���S�²}���qz|��RKG�V��&,j�o'h�{�`��d��}��>NBcRޯ}�S;��z!2�����wۊ���<9yr�3'Α7���x��4UF�zPx�=�]�s�+3z��E�ڜʮ�^Hm����+lj��
��Y7A�7ǧȭ�xO�yu�z()�����=�ǩL�0���wfj�1T����ݾK`�7IVe�6W6hR�@%�L�v_Zg+�yg�9p�c���,;�tRY��g�q����f?u�,�L�+Ęl	���Α&�#���
+ƃ����Fg�g�B}$U|ot���j��t����*b���p���p�)��+���Ԭ�ת���r]��E�1y$��������YS&8��hr���_�Ñ`>��q=�9.�Eۨ}�f3:U���Pk�ōyla����;�åB�P�@�C>��*�~�O���j��53��}�/��<49�%楮����̽wt>�;�u#8�i�����B�p�=9C����bގ��d�V�ma�W���}���h�����3H\�&�ǫ�B��������F�]����uzgi������E�����+ n��ɝi����]3��LŀoK��>�MXt#D�U�����58<U#O�^Y�#ҧR�
H�?Ue�f�m,�ꗗ��<ja��o��S�.�J��\�����o��{=|��N����X;$P����a�kP�RR\/���1��>v��	�O$�Y�R��9Ü���:�Oyq>q��0mN�wbi�+n�a*�.�{n��1��g�e�}�`ϯ��mk����'K$�wW}�o�zV�7��WS ���]����vLJgY�q���N�M�":�IZ���9x��5B[���/�x<�Z����=����cz��򂗭j��Z`�8�ԉM�G�`�T�C�l7�Ÿ�w�*	��I_��z��Q�4��U�Vل��)CB�_��DI�0���*��ku�wU����{VN���T�:��O�#��T9u�5�:#�SMG/7�&W��h���<��S�3Ӳ���_9K�����F�p�k�6��?E�y�|�;R5�-���"a��Wۺ�ix\ţ�uu�-3�(��=��j��M���i}��+]�W�����TՑ�	O
�gcS�u(�Xwu.�3�&fIh�li�� P�����/D�5��-i�I3Iu�������@�W-�0Q�/�F�bʶ�n�
Sjj�ڡ���m�}=P�����`sU�) \KR�cN���^�63&~?�^u>���<�	{A͢�3Ο�v�O�o��~��i���uӭ�\�K�����r0���#�AY^.��uj��I��7����\[�^BZ�reBc�Ӽ��xh�e^_��r�Z$�h:K�tG��N����v�����1LP����e�ϕ�S%����p�݌�F��lW]�|��WyX��m�fٷ軖�|s�����.����u����n�0j���b�	�`<���53lk�Vxk�k��}�/"t��Ӝ��w��R����Ѓ�X԰>��_��13�:a:nw�,AA�P���Y4�ʸ�y$�,��k�N
l�g�ٷ��>�H��X��xKظ@���񛖈X;A�u����Ǘ=}�M%�Z�u��&'�F�	-LOWD�?}ا^��=�s��w`>��L�h�/[�N��=]K�."�(G�]ȯ�����N%�^�3>�3��KP0.z����XU��Y�4�d���D��/�wfn�!s�>߱m\{o��%�:��Ҭ����&�\}�^㡑ol雗�#5����}v�����t8]�1�9:Nz�!(N�8�vwtc�u�3��{W`���?7�֚��Q1�_ P��ö%'g-�ASÉ�F����0,ɰ��j��1�w�+�2�=�+��x̛Ègs��pr��*�XZ3&�/�����s��u�o<�þ$�ָ��d��g*f�G:N�h����K��ޤ����ۮ���Vī
�l2��v5Z%ג���,䵺�N�� �*&J@��ɋ�vq�<�3�:���$�	�-�Η]����H@C������ded;�e��Ȥ��icr�m_>ݲ�mSقǅ���w�ڨ��OoU�W�[�~%�[��d��E{$t�����VܷA�[F�Eo�H{�:�\����yK�����Ond�ěxrN���Ƒ��[��fD�����ͨ(���~�Ƈc�bͣ�Y|����c��B�X������c5ĳ5��b�J��N�l7jv�����M˷�N��nT)cr9�^�\�T��9A�-v+~�Z�
Uz]��U12Vmޖ�6[[Ѧ|��m��j�<��GY�>�:��ZU��� 2��4Fbƨ�}���N>[W}�t5,a��I�,�����mM��m��21B��#�6�XU��;3l7KfTÈ=ݓh��0$c��뵦hӫw�9�*�pQ��c�F�`�ff��ځ�a���Ȟo@�yd�+�D:�p�ٺ�mJz�%�9�Ki���H�"�_�K�C=��k��psbg*�}�1���ѲW�:cz���M�Y/hT?�1s7z��EȔT���n��r%�0��	����k}�����ٗ��I����M�uܱ:���,�54w'�,����2�U83]�>�����YEu%n
Bs�@W9t�br��Nhj�����ܵ���o���Y�;�i���]�M����k,K�5�n�x\��ٴ�4��j�n�XZ�Ξ�KuEIZ�ofN,k-�8B��� �j*���-�Jf������KJ��4���Zj׸fh,�;^�j�J�F��q�]������#����ouAՇa���)���KWi���`��ܡsr�Y�5:1��؃����)-#"ʊ�Γ�a�w�Mbl��D���
�6�ǧ8^X�J���Y�[�Ba��V�N��'�L ��w��br��, *ɴ������+���]���xR���m�6�H녹��bU9-eq�$�C3���ݍ�k
����7�nІ�=�l��3�eɝ����hK,6����}w��4j�Ή�*-dF�ͽ�O�Lu�Rl>���f݈`W�����T��g��p"������8%�Qo�@� 羲[P/�V��w^^�s�~w���i)ZB��R��ZJZ� ��r(��1���)�R�J

�ZR����hZh��hiT����J���)����
P(J�\�)Z ���W �J ���� ����� i(���
i���r0�����iB*\�r �Z,���hJhS$Ȥ�)JF$�L�)2U�D O��GĀ	�U�~ykPV�Z��خ�`E��Q &I����qY�Tg�sR^�k�ݼ9�md;��Q3a±�6��{x��ѱώR��5l�7�~%B��f�9�Ӎ^�������0B����L��V�fҭ����k�ͯ9�"�;u�)��ù���=�^Z,�+Lڭ��
T8���Ř���D��Oҗ�^<����A﹑r�����-��U��T��pv��_��Q�"ڪ�Y~{l>2ٖ�ͱ��VG��Q�`�"����QXϲ������"��V;%��ZG���x��V6�yM��4e��=�be�o�#��e�CL����߀�|׭x��X�H���!(�}�b���Ѥ�-�N��(W?��|�-a��}gO+;5Ab믽�ڄV�Hu�Y��'4oi�RA
�H�Z��*%�;\��nQ*㡏;�iv�ot[��ӎ9�T�:?�y��0g`�=�7]���{җ,�a��w��+D�sú�γP��ޯ8*�(a�Wva�zi��[	3�!�<#���h+lz�uj�A�y�-\�V�EXs1��QkF,�"]T>~��9,��������&Aˌ\/ ����r���tp�$M�b�^��B����)1�0�~�!�mR�bg> ����?%�_��;�^����a�y���k)K�~9%,9qj<��Hy��bKd���2�Xv�
���['�2�m�n�)Z[�;{Vs[��vu׃§ԭ��I�ta�P���I�)��J�Z��J:�eݙ��Sν������'�E�m�hAi����ً�Cۦ'l@^|�@)<�|	��ק��+�7v�:��3���Je�gèL/)yև��Z>�K�U��c��!c����O,j���_ptY�)!��w=ˍ;�A���,ʖ5X�����p[Z��"YR�)v�zBq˽G�}��a�AX����7�ע}�>J����0��OR�:{�N觚�F���w�-��]B{l�jW�.�3!�T���5��d#pV��J<M�ů�j�m��1GW�����G��l�|Qt��V�#�}O�B�)�Lj[��
gyxE�Ϫ�k��r�����*��y_�\>������3�e�G^���E���xQ�s�}OՎ
{W
:���[��\�/O����h6֦}J��N�9R����L�"�X���w�L�ZY�,��s�;Vz��v�Y%�H�V���O���~ɏ'��٫K�1�'U��Rv�E7��Y�3�oz���ud�{RT8{O=@����-�ܙO�A��u� �i�J��F��ut�S�mϐ�h;K�/��L�[���Z}�*���fې<��C.u�TD�`BM���kz����{s�r��R�3�A��p���醉���$�#��qxg\����Xrc�Q�.>��è�شgeKOs�*��1vL�l��p��4�}җ$�.�����CpX�Ӟ�s�|�͏X~�����ز�L��d�kF,NR�T:�$��>�e���wЊ�^�r��[�a���^�<�-�Xpo]%fEȮ�8�F�rR���ݶ>c��nmJx����i&m�����x��t�~����>͊��κ�@�Hy�z�|f�ٹ�|Ƿ'�e�(��N��U�+�Jƀ��-�
�;Bگ,�4.�J�k}Yo��۸[��x�>��F|��gå�(M��bVط]5�%R\/֟�eLn�r_��K.Bc�^�sZ6�f��/�*�o��/{��\�����	ᄋ���w -�7/�u5�(��%�0_�H�V�����N&���\=�q���+N�ժ�w�tKO��C�Q�o�Б�/A^��m�G��h�^_���R�D]�����-Һ��m���k N��l�R�����P�,]������b�-�f�������[�T�6��˫	�ky��A�x;�t>�sc�7�z�Gt)����Pvgi�U�u��Oٚ��[ݓ��bsU(t�<\�@���kN��{��/3�,[���f
���VZ<e�V�=��8�zT�9���`��=Chcڝ�ѡ�#�Kρ�x�+���:i�
�1Z�:EVz|ߨhN\K��pLT�7�U�����d�mXbUm9��+<��QުG��p6��#��������`m���j�<����a�{h�NyG �[ޯ|�^G��},�.%����A\/C����"�ױ5��{�!�����G���Y�=�1�Q��什[�ћ�b�B�Y�Z��"p���̗��\���e	u�����=��:�k�Y^!��'�bpL��>��a�����V���ޭX�Y�ݢ*���Ԕ�دIc~��^�r�᮸��]K�����/#ӽ�-�<���(P�4��$���W�}z"�Pk+��6+�Hxy���=��5/����^��m,~D��Wr8v��vD8;�]E�zʳ�qz�����8wN
I��]SkΥ|=:Y�	Ov>Vs欰m�OR����J�fB_Q�R,�b�qp��5�R}�kb���iR���PuB���{�Y�����^�=f��~8�ZtX-vl-�oc�;�&���^#iyҞq�T�>���0�,!)ϫ��ĭo=j{c�{���6,�V�ڷN��f��x�v�2��E��7��y�l>b�n)���Q����ړ���zX԰>��_�s"Zg�{��{�
���l�w���x�mR�rR������[�ཉh�є7���K�R�}�[㤺���|�Wi�۲(��<ޱz�r},�l��LB{���e�"��������
~�S���ܻ�-A��J�����[6����V���X�<EF*��e�=�ī��Js0�v�jfnÎ�Ę�� ���V���	��t��q�Ք�д�r�(0B��\ �4�H�%�[������*�H�����:�%�_a��y�d�FG���z%��EV�t��o.�P�ϧ�LX�m�X�^g��n#s��o)�P��ӽ�Y�x�'��|
�"�Y�:�����z�ֶǛ9 ��:�T�q)��N��>�,��d�C��v+*� m�og��l��-��{�N>/�Q��9���a�w��[�,d��7r�����ھ���:�E;���cn��2v=dVϫR4.��r����(S2��iK\G���ߗm;��vj��2kW7Ԗ-z�eMF��8�v�n��,��x�dz��qP��`i,���r]O1Q6�[��W:�{˗�yR���{B�ۖ��ȋC7�r=��{���t��s��_�4s��!X�[�mdfp��4�r�:��-V'�/�����^�8�Z�vcׇ'z�,�!,	@��kRG��)�qx����[�gI1��خ����e��gs�����a������"�	~�Y�p��ZU�qu��a����d�Îk=��~�yE�#��WN4/d��?�ޯ8*��C���0�A|8V���i��Un/X,z��=��} ܙ㾝e���0$��*V�`��^Q>0̺�>~��9�aoD��֌���<�ʥx-&� �ك~ޗI[�,U�,0lI^kR�J:��׏g�ow��"B����`�c�֍����#���LpNס�u3�.�UX����ꯟ�;C�םv�T��[ܞ��ўFǫ�$�>5��!�5��g��U^+��Ṅ�x�:����7Q����~�z�E�8p�ӼG�q��3��G�Ïg*��^k2��V2�"���h�;�X;��u�2�n��>���VW��%<Xu\`�>���
�J&3٫nKi�b���g��&������u�,4k'0C�A�sԚi��.�3!����q�Ϳ����)@��%I_�Y��~�:"'�Z9H����7���֚7�a�ʴ�k'�{��Ojzkbo�mH=%J�N������ֱfmf�st8��ңOQ����e�kY����wI6���̘��Mճ�����61����w��������R�$�3��k��w�;i،����-@[����"�Y�F+NB`j[հ&}������Do��`����Ѣ��Kb�]Vf
U�`�vZQ�u����_c�ᆇ�ӱ^��;�qS��C1��Oۣ��ߕ����@%�l%�DW����r���
n��'q�.��d:W�.#���1hCϽ�þU����F��,��K��!�r��8+�yq��|�Y|Nh{}7���,/��mQ��Y吝��%x�����Α&�#��B�C&b�z�eZ����l�*��{��}����������<=���Y�Γ��h��[oN��M��*lRG �4:�YoN��U�3�zWAwLg�YG+��ñ:P8C�]��q�-�ʕy�<0�>ݲ1�^�j��j
ϋ���Xpo]$$P��탎Q#E��X�/v.b�q���0z��D�:�0/��2�^��.h��ᡈ���.���a57��[��N��v���Li&��>�'��zא|�MC��M�LT��j�����2.�E�����QKb<�k�����ӯdo���YO���;+]f�]24X�ytg�':ez_f�x+$w(�<-�}�/���9R�$4��kcO��C�9d줅�Y6�ھ=�&l�q];<�;�H�zN"m��}�Q|��J�9������ui[��h�F�az�t�B�d�LlWi��K��U��J�z5������W-��f�u�=t1��p,
�E���k��}p`Ъu谪���45(�n _v"��z�����9~�"�9��`��q4�d�rg�˞
գ�r�E���x��#q�K���^3�Jюɡ}R#������)ՎϹ;qB[���z|_��J�y��k���^apL�Z�ȯ+�j)\V�0h_S��ɷ���=Լ>�yֳ#�K�H)�T8a�VZ�-i�͑Ԛ(l����tҿ���k.�ÇF��ώdt���bp:�8_�+�;m���l�A�D�tH��J��Uw�`>�s�].{Mi2������8?�k�F�o�gm�4O�����A���b��c�s T��~�
�gw��,�$t��ϗSi��{T99߭p��F^	�;5\9.�%�-zn�l㳽���1�F+V�*��������:mbu�[���J�]��LB�L���wK�r���۵A���#b��j������4�-��iu�ܣ�j.��4ɥ����Y"��}����%�9�� �1�S���c];�]�X��2*f=��w�G�Y��.o�^��.j��|�sp���i��y������F�.�o,��nrו����<�Ө]໇��/�����oL��|6���cz{]�{P���Q�A�=����U�.�l�D������-ixnU�����Cb�䇶��B"6%B��c�ms�pg���	�u.�$��TD>	�/��H�[uL×�ȳ�y������z���-���a(��}��)�](�h���8��%��ާ_#�o:^Jr��3���m��P6='^j�}]�f���`}�����ά����13Vv|����s�^х*�qƶ��S1����^#�Acs�cK�y�J>&���וy�5��v�=��j<*��k��[\2e�#Ԛ�!��'�$)���i�s��Q"?&y�N�{�}$���P�Ղe�Fx�:)�<*�^񹩎�(^�U��Ϯ�i��V(�-���9y�˂KP���wV���}/؏��5z������0B���[�3�C�{�,�5�_�VN'Y� �z�;���u,x���z��C�+-l-5�eV�x*Du��su��{P��#�~���{w�x�Ԥi�n������j�x��)6���N�|
"���.�Y�m�\�[��R�:�jݥ��E�CEM�K���ct4�����?N�z�x�m�Շ��ɒ.����!�)�weAZ��|�7�tI���N����Bҩ�M5��"͗:���_5킾����pv��UGl�
��:�ݝv1�t��W{��v����V��fSiEby�Yơ�8�dM�Cs<)������.�n�\��|'�i�`���1ݗ�U�:s��!�^N~�~�|׭x{�*]�I�����X�1�R]���h7�]L��L�M)eq7��o˴.x��;��[W������y�E��ޜ쮵�K�P ��CZ����o���#��쵛�T�`Yl_�	��M��eK����7<t?��i�Pd� 8R VVu�Y�uy*�,���-x3z���%x��Z���oz�
��>uwe���4#�X7���sd��|�fr����Z��YW�u��;���*R]�u�-pr���2�]�d�jJ�q[��o�OT��jCCq�Mۃl�c>��4Oo�U�E]A}%�8Imˀ侖6��T��g)��]܌d&�@^|��P�n��φn�4}�P�L&��sz��B�ιu�A�]X��ʹg�p0�5@�K�������V\�%�^�Pu��^�E#�xo��1ZU
���wW@ͮ�Nҽ5Di���4w6�TGRZ���j������j��Z�U\�N�*�Qu�U�힓5��t(M�{T��d4L�XGi:������K]��9��?�ƒ!
ȏn=j��; ɫщD���뎟<Õkh�	F�V���:[@0Q�k���/7+'Y��z\�[����1*᳍��,Y�ث�4�%��p.\u�k��CH.v̫V�m�i����U2�S[:jT�xD��҂��e�Z�u1�pX�Щ$C���j����/`�Ύ5���V��L6�ŬǏ�>ӊ.퀑\�n�w���YS��y���e���0j/(���8e�j�e����gEZ��I	�ɵb9� w9%��$E@Y�^<���-� ���"H$˽��9���u��k�]u��M�+TB��Ӱ4$��K0��f�#�k�R����XlT/��W=�W$���t4�;�\uU���!SN�������{Aı�ѽK������_CC�� ��uV2%�B岯;W)�p�0	��{�����n`=��ZK��ǂ4��|/V]]�a��έD]����[+(w7�[��n�+-��5�����

|��8����w
Xݨ�����s;����=��D�K����n�0P�\�Dt�X�*�`T�������u�붋o������rW[��BrioNp���=�k��Kf���{H ������a��]�e����C�8�����ː�A��)r�ǑN �%uw>��a���1������ܦ���JIge8���rvg5����ڬtG��֋�QR�䲜��u0�2��;�;9X\�CfA%�a� ͭ���W�ƕqx�����9�W�"�(�P+��k��b�v�J�e�Mqx�}-���C!؜�;�2�K�;N�h�zl�G/�v7�/Zj�[�%9���DJ}CtWH���{}ԑ�G����)�]�\x�u+hV�=<Zޤ���ET%Z �ή��]��]@��V/�Orȳ�]���5�ӒŢ�i	t��u�����3��ݱ��s.��V��y�#r��{k]�jZ��K�\�yWw�xD���K׈a�laU5��Q���:Qf�������k��w�o"�!nU�z�}J�"��2�.3��4��k��\��y?�y6�Τ��<J��R��f�R�M�G���ݏg��;v���g/�u�v6�dߙ)��>@�:]����}�m�Q�0]�*1�L�B[�y���Ui��Z�s��:���,K�I�H
tm)ǃ�v{�45����1��d�j@ �,�iT#Znd�7�Q4�C�.�c5�b��}�)*�+�ŒU�����赈���r���SRT7����;W�1��J�/��+ބ"�e�jf'Iݵ�A+��t��mZ]}�^�R%�&I�e���e�@�
P�Hd%�!B�	�d9 P#@K@��NNB�Rd�J��)A�d��Bd4���JR!KCNBa#�+@䔴U!��
U U*d.BdM ��U.KJd&K�&KI@����@�d�.I@*䩒 fcI�R�-6��&TfFH44.H䁐�R`�f!�dA�Q��}�}D}�Kv��Z��P�U��DZK��,0R��un�e�O^ �+�yq�r��l��d��1Lefifh���v*�d=�uLF�h�;'Xλ��^g[�<y�4ք=}VX��{j^�/��V��eT�pu#�����3�x5:�z�M�L��v~S��4����v;��>�����
�5�Rƫ��ר8��yUY�_�o��}_�8C��z��SŇ���r(+._�g6j��E����)yo��R�{bS�4�z��+`�V�0o��&�����s2R��p���>>���zlԭ)�2{�{�s:iÅ���]މ���Y#�.��9	��oW�
gyM��'Ws��
9�(��}�V����f��R�.�Q{UE�A����w�9�놰��s/�K�?cJ��Ȏ���uV�o�*#�$��IئҮ.��Ί���9p�Ip��f�^�pU�E�����V�NGٲÿ�V��m���4>�YV@�<k+*qɃ��G_F��X͜:��2�rѝ�b��͠��.g���g3�^$�,�ps�I�8����7v��xK�{����)𺊨���C�*� ��P�X$������.��=G;�:|�Ã��B����Z�Q��i�̌��+]��)}N�M�����sX����K��p���� �Yسm9��훵����h���)9�b��4����m�x���8d��N�j��Y� ��սAfӹ=�(ZV�k9d��X��PO��W㴷xDY?�J
�_¸b�hu쵧Tߺ�;KɁ�+����hr�յ���!@S.�\���Y����%V�#l���Uw�E�;=a�2�y��U���%��m�B���?�G��m�J� ��&�.Z �{�9��KM}��YU�QεP;��=�`�p֯-��ޞ�{2\^�̺� N���e�ԍz��ּ���I�sw뼈X�-�4!4�h��S���o���[������gK$M��gü}a�Q��`���R?<��5=��<^ﺚ�R��V�'y��ʜ5ҋ�.'��\7r������\���=�P��06)�9Z�̼�i3��P�m�/դ1���5��`����c$�{������n��Ȼ�;���qg�}��4U���X�b倹̚�_T���o�$�m32���K���{������!�ul<���vˈ<�Z�ȯ+�jg¥�W���N$v��O�(*�}C�!s��2��'���ʣ��ڇ>���Zh3���Y�ߨhuS��o�yԕ�̍@��2�
�],���\y^���Z�B�m��6�g��2���J��DT�j�����7���V���\R��:o�_�k۞ɴ�h�)�+k�$���7K���j����\yzr�>`�ʄR"�T1Y͒�ʂ�P���_^ѷ7���J���+���B/νn�xJ��/�᝶��͑��ж�+�+x�֦^ZiU�A�l\��+���J(a�ﾝ��y9��C{��L��<g��NR�qm�x�S9���Rq����z�	F�1�5��[�y6��=���6ק���0v,j~赎NK�҆��ir�� �}�I&dHG}|h;��t�ϓ�f��/׃�P��.;�4���۰�-��'����F4�T�Y��e���냗��S�%�W%�A���Խ�T�R���|�_tO�n:k�v���&�I
�i/��G�o�l�<3qPؼ�IB�s[���К�2H3r�ϝa���[D��
|�J�Ի"�4%��>[uLÕWu!W#c=���=�|��W��0%a�H������,�d���fW�Qm�v��.���s!m���9g��^V��2^5�����cR��9� �L���3��ϯ�����o���<HG�QŶW��3n�ͽ����H}h�Қ��HdH[n�$���k��L�:w/������ts�3'=2��b2Хf�*�j���'k/��Q�:M&�5FLm��������s�Ы��Um���פIx���WH�Yd����۬�|ci��k����J����gK�a��.Ƣ�Z8Ρ�+�Ǻ���SJ��<"��Y���˂�e�#Ԛ�!��7�
e��8��ܷ���S��@_0jgw{`t}�~S���>��:t���e��ڜJ�G6�1�;y~��s��̈́�6U^o���]��Nr����r'�,z��<2��i��Z]*���,Jw������K�����3��������0zu�]�.ϫ-N��%�NZ{��G�2�*o����AC�(bT;Ԣk�,�ΨqԾk�`���=�|8Z��DǺ��9<3W����6Y�;�>��3���S�A�5x	Ԣ���e�y�`N6\`����5�+��d��*ݭV�#�.$1���C�Μ�tCL��<n;�kW�W�g$/Z^�,�i�DM�h�Z���ϨS2�SJb�0�s��ػΪ)kx�s��R�V��j�E�e��x�0!4J�CZ��K��=j%Otu<+�ݾ��ߥַ��(<�����������s��a,��H�'��x�ѯw��!�oA������7j��y ��{{#����\Ӂ֛�*30xK܀-�*x0��W��!�ԮO)Vy=�q�l�:��S 4�7/4hM�J�����M� ��Si̶�E��
�V�j�\˱M��J���i����r����õ_dcz����ZnzZ���z+�8j�ɸ*�Pö��0��F���V}��D�u�C���5�\�E�|���Y��`IX��
��`�r�\2KEܾ�x�WM���g7%���8�0�����z�5YV{T;j��'�P��������}h����5���K[>'��0��ۑ�֍�M@^�����c�v����j��^p�nS�<����N^h��h�+�}��N�ʯk,�����\U�}⸡N̄��f�8�*yvכ��g�y~/CgN}��x����_{���.4�}o�����e1O|#��%�6j�H��+��f:�t�ڔ�p�䧋���9�D�al�,�%��o�nm�)1yU�d�	��خ
�ZY�@{�I����+�́���]	����>��wG��$wU�9wȧR_����c�o�g�,���2��ꄛ�R-��ΌV"��Ʀ��]W��̈́&���a(�f��g�i� ���euYx)W���x*�H��A�g�i>�y+F�sÚsW��- +�,��HS���=.N�����CxhN�}v�I����T5�6��^v��ɏvN��f��=�{*Q��nv]�z�uaWb�=!]��3�=�*��[�0�������iޱA����mv��-wF8�����X*..:���[� ����Dq��Z���0R�/.��r�?.������N9U��Mc}�#��h�&�9s{<o�C�X}����?24y��
9���V��J�M�:A���J�#%���Ń��y�G3�Q��� �}S������$��o��F��z߱�E�D!mL��_�9n�ҡ�bU�Pp�^[��1vL�l���?-+w�����X�b���e���g���
�cZv�ﺃ;	y08j���%+Z5ͮ��i1�m{������R���u�J�ȍ��j(1ʱ�����U��8�bmˮ9%�j�T��q'X��4�|_�?z���0/��2��z]��G:��F(�Bރԥ�z�ud�*kxM[��&�pS$�J'�'��y�5��O	���w7��#����J}�t��n���v�c2v�B�q�=�`�d�����}�>��umd�]����%��9{%g���Agr�hf�;~����8�r�X==l�h�t��^���d����R#Am�v��p�w*�fmv�-��)�wY�k��*}��/�nںe M�f�맩�p�:0ȼ�<���,�fz��e��D���Ώx7��4��Ŷ�*�7���y��v�aU�QP^�K�B��o1L,�o,	�R���̃��{���U>u�T:�5��w�~�!���5��`��q4�J�uz�Q����
C7�	�_k=����񚆫��Ux�,��iV1�4/�D^�I`V�0�{Mrj�kг��l�Y?��;��$�=盋W̅���+��4/�Ď|�ԉWKWs�<5��W�.���q��hxl7��xùYk����6IإCf]�x�ޓ=����t}z�g[�S8֗��=CL<�v38�����H�A�N�緾��q򧍥��j}r�n}N�^,�=�v#���QϦP��8S<���E��C1=�.^Y�ˈ�m�԰���5���jWb<�]�7�2s͵離�|MB=;�Z���И�l�]9�F���t��_�LƲ�dP�4��:m`N���e���}+9{;zC����чg'�}�9Y�i�FV�J�z��diV)�.�]�����+��9��Q��s��뾼���*�����3����1xS�)N�>�d�Y�i-r��>o�]���֐�J��:un��s,w>�j�c�>��+ʺi���N�)#�{y�`�Su���Q1نʮt�S��m��B�j�mk��8ŵ4�X$���ʃ;`G�d�Q��Ӧ��� ���hb�vy��%����Tm�J���{��j4q^���A�v����7�w����KA{Py����Xay[Dゟ#�]A���@��u6����Z�����Չ����{%�W���3�XK���H��VX6৩g�,��+�q��GO��^�le&s���
ת��w����63�^}]�g��ƥ���V<�0p��Y#��v9uV���gz������c�
��C7`�gE�b^ُ!�o^
_v�U���_D�Z�^�����f�-I����H��5Mc��U�����>b|D�v�{�_�]���4\��_Wz��m�y��wC����8+�b��X�X%��]!��	FbCG�F���a�����ד��bv�`�a��KP�Gs����~�|tN5z������:x��2���s����8�L���:��P�:�<sӯ��z(3��G��x&t�Y�7�o�i=������W>�C�.CK�z�M`{��eΨs�R���}��;�e��{�����/>���%i�JZ���Ȓ\e$Gw�O��A�5NJ&'�e�jk���ҥ��5�1]�55-]��a�.f�t��<��S-�V�3�T.���ns�/%Hỽ��קO�n�+��2�B P��6�d��	x [)�fL`�N-��;�N=��^>£�7fXjTu�6�e~��ff��m:����$����p�v�{���ǚ>��c�ݮV�#��\\YA31��U�-s�6�0���������
�ݽy��%��|�����EIT��ɥ��L�2�%'�\G�$�4��EC����z��D��|�W�n���o�%�(BjW�.k�L���z^�
������pbJ�햚��/��}/�c_�nx�uH��y�O�p� �Y��7�=@?L�8ԗ-[��U�e(�>)��|����[/��8Rz�g�|0�y�a��^Y�*Uɓ�2%�W�pNWW����u��;���%B�&c��
իۧ�����{����D!�#Z&�6{H���|]�&�5�1=���.��^|�"��!r���'�P����n�y.��#�ѳ�Z��#���oVx���p��Ry��,?x����^�WJ�7�)�J��b��6:)���Zlӭ�,��*���G��ܿ=b��f:�[>6���K��/�c�l��8�8�f������δ=zW�'�UO&��K�?H�-i�}�,G���enMqVR��LՑ|�X�e^�Ɍ�ex\�,��m�c}5�A%�#Gƭ]ZL��@������c�t��?F,	�2rŻP޸6u�}��a�"_@�c��Մ�4��q��b�������Pn�������mT��T�A�{�h���³������%<Xu\`�>r(+��a}=6X��ݤ1��@y�Os���N
�u+
�=䚋���W�9�@���,N0f�U�����m�����zX���pf������bKG�����V�#�>�
�i������.�V���S�i���Rw�~�gyx�JP-PKRؗ*-űr�Q�l=4��z��3({�c�Ov /���4����l��G�a�TG&��N�\[���f�%֪�q���f���y�ufr0�-��F�X�)�����Y����
T8VPD�E��cF�b�ye�X���j�y`	ˇ^��|�o6����|��p��[ @�����&��N�e��|fֵ����h� �q�����A��[�;�^ʿj�*�$����Od8j��=��W#���gKx��z��"w#���V�������\����;}/&���,�#��vc4��k���r�~ORJ�)��E"xm�b�e����։}�PȆC��B��b~R-9NT��/ki�����.�F���1��ˈ]�^�)���i`1�jp���SX�k���Gr<ufp�ʋh���^��-ۡ8�V`B�Qk"����
h��"��B[�@�s��F�n�����`�hPLPW����Qoܯk/u�7-���Z�׽F�R7G\"�ºi�uЌБ^P�{��sO��[ܔv�g[��y�v�%\$�9.{5s���ݺ��y�'$�8۱�m���>]���e,�
燲Y��Q�1�[��$�t63M��5��Z��R������)e��Aa`���"$���>"�Sy����27ieq�Tz���U���$��Ij"�9�6w{+��u�Ն/;���nggSfBX��m�L"n�=J�zmm�������m�w$�:.��v7�2'�<I�����jEM�"7{�W$�AN��.���3Y����#w��[w�N|���.5gV!�Y���z�ܒm)2&������H��E4�OD��R���3st�sf�s5��:.fm����\"釢D˜��GOPB��_�1�7aKq&գ�(FQ"Le�}��z�\�Gj�3v��O�1X�}j��m��9q��M�������A%�K��Ŝ�}x���M��	@@�����
S��e8Ku��{KX"l؇;������k� ��]D1\YML�ïZ�[ �yP�9�3X��ݲ�+F�U�7wyX|��$�-<���8[�[�t8�����[\A��e����)��G�,S���Y���v+����W���:�K1�o1w��� �Eerx���c;&�}�s��Hn.Z�;�JB�9�Վ��o��Y�����`Sa&�ۓ����q1��m<��2�bͮ�b��Vy�X�ñ�m�:Z����S>�m�ڴ>J�#���������/��^<��2�ԝ]o��ҁ#��[�n�;��M)peE�ֺ|�s����m���1Y�b�i��U!��E��5pQ�]�KBe���<5{F�� �Q�G���l��b���xe<X��CI�"T�e�f��.Z�o��s1��1fQ�H"��|�jϷ_6�Q��}w�*⒝��SLhR���w@ �ޘ����L�:RK^uՆ<���+��� �m�wy��IO���}]I_y�F��O����9@nŧܰ�T��R��Yjo�K�9��k�Zl���f�r���) S��=��^XF�|��*�5�+|����j���wu���uG�^�o�іN忴�ʇ>ٗ����7�&���wl[ATV����s���̮�z�.-g:�a�;�6W%��6�Jj�Y��)���q]�֧]Iq��&o;l�ƅ<�!��#Z�r���1��nCږ	���u�]T(�am�y�O,�)7WZp]Y*�D;X������{*4.�3��gk���Tf�ިFƜ�^�S�
�sZ붷��_v
Z�u��Wҙ+�FIIHe�de#J�+EVX+�f(�JDHіAJ�R-NHa PdIMd�J4�J�f4�+�d@D4PR9	��M	@Дd99S��Ed�4���R�T��9-A�K��%dQ���e����PTeE��-d�CV�@AJQE%9!��d�Ye��YS���d�Y99d�KTNfP�&I�SA�P�Jd�
PR�@�d&A�-U1�ًK��cI�W�����GZ��{��W`�-oR���!:��k��W���v��ˌ/p�{��B��&E�am��ZĎ�]Lf�w؏8Cgegb�/7���Zw��w��tH�o�)y_�{0O?Z'èt7K�E�2�.
Ec�����תz�Ӧ;]�/�:�}0��B2��| _l����R��Y��յx���C��"�7�ٍ�-�i���V����|�\;tw�}��_{��;
���77�Ô�u�d� �l�^;yVOԖ��ni��Ln�%;YU�u���Zly�ize3�¡��<��k��s��2d�xX�ceW[��]�������p_�HamiԻ��؅�ja�*�y�3�'�K�=�%f|y�u��/e%c!��`.sU=^���o�$�L̤P�:�w�f��>:�^��9Zb�/�k��.��-ɢ�P����m�-*.�������՚n��iV�,}�&�OR�=�"�s�FT����Sz������\����?rO���"�u�۾��A��)�sMC7�N�e�X�:���+<����`wh�aq�,�1��]RQ�{s��O��Uωύ��-%3Ä�7�A鼬�C۔�p�/>��E��t�����Zp�n�j������YXF�'.�ˍ ���+�-\�$�����kv)��d�eУ}6ٔ� A��S)+�i���N�g��l����E�æ�n�����p
��:,ЏWT�:jNh*�aw��ab��t�Cΐe����V�[�Ή�3���`�,�G�ԃ���XSi���'<�^��FZ)�sv�G;g-���xl/)#�Pz�+4)�\��3@�+�P��i�3]l�[�1W��>
�xg/`̆{�9�E��g�*b�/��yHiK�:���5ڠ95�غ���8�y�_'���X��j��^��Wl���Z�s�2�+����B���S�2���v���t�sea��q���%���Fd�0�U4N�>G �!��ȇ>~W��Kl��`��_��of'�td.�~<}{Y˵i��W�ܑYȬ�_z�a2���a�Yr��~�NW���Hv��PR����ʆ�d��ϫ��ƥ��*����>N��\���%�WyOs�=Uwy�
�_ڄ-}@��>��ؔe�e޼�e*�Ď����y���:=�zb� �1��oc��#��U-��X���*b|G�5�B:��w.���t�)�zq����K��x�Q�8�Lv�x7�V���RF�aY���Q9��}����m~���d@�x`J�9}��A	��	�q����_��Σs.����ʜ΀�Ð�nl��ug.x�z���Uӏ=��Xs��2��S�N����H�ނ�O	�]Q�S{���W9:ۚ;
|�5Ϩ>�c�=D��٘)������S������籑��4Z��8�9�f�~�^�Kd7�}��`�θi�Z�ZY�N�(|K9��[���K�r������)M�ݷ�zgx��O|�3ġ�(�Lī��&���f�.uC�:��l��i�G1>�%M.�_rh��7���`6=��t���$�zSHV�W�
�]��m�c�H'�2J���gPy��N�*�|�3�Y�h2'ӱX��r-#��qq`�����C����s���$������vL�&'�COO�w���x�j��l���F���r�;l�)�yM(��j9���ݸ��,w���=�ؼ�:���}}&�u��C�H�`�kR�K��Z�c9��\�4Z��$�x)��`\�:}[�}����k�s�D^���D�
@
�do)Mi��w����J�s�ʂ���˱8���UZ�:[��z�U��s�R�.�U�� ��'�o���xp뫘�R�LX��D!��H�g���w2X��c�;���IP�I���f`���{}�l��PN��G�^����;��Vd~�I�V�b�����u�,Y����Vf����ĵ��}���e
�O���5m��ϡ?4R���tAY���;�����֫M���������;*8X|�t<�#�Ƴow�2��#�w��z�kz������m]{��F
֗����g���
ᨶ����^���=��������m�ű�G��.�cYN��`@>���Dퟹ`C��o
�������sǅz�j�˕�ڡ�|7&���']1��x_S� ������>5��!�?}����t�}�uy�{3ݽK�����@Jzo�(u�~6t�q�9����:��#��Ǧ�Ǘ]���k���~��5���ʖ5^XdP��`���f:�k��z�zK�o��~;�U��W!�ɃU��:��'������P�V2
����5;��t�d<�?$r�S&%�MTlw���r���g�Vj��V�Z���/ -���;��W�xƜ��/�lvf�v��'�ӕXyn�uS;�L�#���-Kb����U��ltK�H��Yj_Zʿp~�E�xt�j~H��� P�u�킷���2���M-�Kb�J������6nZ��j�f�
��5آ���h�ɹƎ|�o�N��Q]�X�rF�X�YC$��'YV<�kh�^d�v���&�����(�Z��Y��,V���2���(\�
����pe��p]Ƈv�����833jP���JT*�}{� ��Y����]Y\�N��0�ݹ.���c���u�WD�r'[�\
�݇���VVV�˖�\�-	ˇ^�z~���Y�)��|$�+ x>�#�sݔ	s��۸�'֑'�-����A��[�;�;*Zxk���,2�y`k���D���׺����i҃�sF�t�w¶ʡ\3�]s�Ӷ���ʶ�3��vVͺ�1�t�z,�J��n��Gt�'�W��Fٔ��Rt�tX���[l�S��D��=V3Ө��R�^����H�2%��=�'��%����Zk�޺�5�S�F%J������y�����*�L&�:�o�2F��.��r��f�v��z��JGv�MGނ�K�ۥ�ڢ�Ո�\�V#�ѿ8��԰t�EM��g,!U�Le�-�0sΞ%h|�u\\}0z�!�T�~��Ƿ,z,�����Ͻ-���d5��
w�f����mhAܷFr�V�>K�T9�P��ZChs\�H���
Y�m^������t�rG�e��v�i�cs�1[ �c�`/��x�]�G��`�U:p���^���p�Nj�3`��dަ	�4�֚�\�ʽ1���ڻ�]�����;LK+�6'��8v�os[f�MZ��!G��\�Ǚ�E̋{��\6��"INŴ�WN{X���p�_0t������M-��ŵ�7\9fy�u�ءO�Z��v\���y�sW����p�Oy���ႸR�Ѷ}����lmX���~{��3�5@,�&�"�s�FT����Sz��;���!kM~䟥���C�+Rɋv�5�w�y*$��g�v#,OX�:�����v�c}��ʠm�E���;����`KH�"$V.]��w�X�e���rs�<&P��x8i�����S������׶�j��:BD�8��u/��&���9�ڪ�8�.鶔%�����V
o�g��r] i�\�LƴPL�ƃ���k�f���׋+��7+!�|b��0ެ��ꘅ�jZ�~ �h�H�'����S���{�-Jԋ��fcxN���{�K�g��gx(e�&T"����yI!�5��\e�<�Y��-��#������ �@�Vn�Fd�0����s�>G%v��vD8�M��n�+��=P���Y}q���T����=�~��wW���\����WJ��}[L"���Ϭ'�̧��a�b_���W4�t��b�lU/v�&`�����R�/�~�c��i� 9V��w`f�3b�������{���E��__sa�c�8'w���<n^D�b�����Nr娕�bާ���]uf�t�j]:�Vrd퀆4z��k�ji�H���t����^}]�f���`}���1��X���}��o��f7{��ؗ��3��#�����APs�B�Y����߇��<��7���j�zƧι�p��f?y�R����x�@���z(v�5�U-��X����\C�a����l+i�[�����E����!O݊p5�$��ђ��|g���-�q#�Qdb)\��'{k������R���f��v�ϩ���}���=M�c%B��L�#�h6Ͻ�綠��W��#Q�F]5`P���Lv�e���t�r�Υ��oWnK�N���v������s���t�V�>��S)P�.��֙�Wz�Mc�E�.uBԮkA�Z�3����f�ǻ+��k����Vf�R�A�"�U\f]Qb��W� ⚽:�Y�ٞ^���>
�F������k�C�v+��r���xX+��(&e�we�:�����{6]]ʪ��_1��}L�N~�~�%�^�!t�u"%�v��ɥ��â���aI����]�#���Ԩ�uƖ���EPM䘓���ǖ BM��vv�K8�la�����v�e+6�-����,��.�+:�A�q�©�a���H��}�(�}Cd�)m�hDԾ�QӍn���1�2K���W�y3�]�cz�wi����[Y\�W�z�&�;��FD��E;�`�������Ǖ֘3�	bP(���*�e�)l��־�M2�][z�<9��9��{>�~���s�C���G&\;+,�Kv��Vf7����5�@S2ρ_Y�yz��ҩ�\���n`G����"�z���+��[�Od��Yx�qk��.y{�5�@dm���u�������1f�%bJ�!�����ZY)�=SYO��r�.�t�3.�σ�/)�u0�zן��]$׆�#���3��Ώ��e^ݓ�*����/���	�C;5��w�#�e�chv|Q���`ٝ�� 0:�[6��3v�#��-��kΡ$l�oJ��+�`�^ܥ�y]}�W���g,rq��붍���j�`p��x`�ݗ�چ���ǈ�eyh֞��*a�{=���	���8�.}U�:�,B/��>�6(3��f:�k������
�@�mp�MG8(��:��)_�5gr�֦UC�dW ��ޤ�>���
��{�YSuk�<l�^�����Sy�����S+�5��*��;}�{\k]BB9����jV�.��o���ڲ�|&߮�c�K�9���Rs5�zv����q�%J4��G!��֍C���idAm��M�e�$��Ss3vF%y�x�8��Y���yޚ�:/=����%(qz|��$�yyt�x�H�!i�y���7jm�5kx�XyO��q	�5-��>����2���-�>��/*��U�+��
{�LשJYĉX��3�ic��X����`^���Xx��5�<NPtNx�z���ꍏ/"$ʍ5���r�k�T��'.�N�e���G.f����Q]�X�}�~���^��)[���$c�I�[(P�+�3�WT�ς���1`�Ut�mU\ϧ��1TfS�q����N�z�XG��|��3��qA��9n�\�qVy�z�i�O1h��\�g3.��f@;��4�A�ő{,�*�m��c�@��V5�m���BQɅ�(AIZw�/c[*+���r�s�+Z1��	~ORJ��Dm���R%�_ŋ�q0�����O�x�>��tq��˲`��ިR��`VPU%�d�U3�h����+뗡�&�o�e��c�Qb�x��a�=�>ޗE[�ՇB4K�2N��}bE��š
�����%��^W�B��7H	n��X��D.��[�w�����|Q�M�����B[��������)��ƵWr(rWdCu.�{����gr���.j��f����23z떈����u��i<z��F�v�V�J@���L�tEL����)oK��pκ�C�1Z���L���)���À��R���w��d�l@RS;�&��2�>�d���$a��#�[�L�ͼ�Xͻ�V�c�rǢ��N�w��v�=��E9i�v��������ܴ �[C��W�JK�꧗�����N�WW��U�J%`K����f,V붤�סϓ��c$�{����ޕ�M�5��JJ�C)r�]T�������vzS<�Mmv��<�d��[9ǉ3��3�9x�R�C�|��/�;��/�9J)ZT�_?	�׹�:Œ1��|��i��%B)9���M����B!�T�^4���7l��rL~���z�O�Pɟ]�0�Ji[�P���F(�`��s}���o��֬lݿZ4���ƪBͯV��:�hP�N���:+�v;;�ɖf�v#��e��˻-Y��A�b�y\�7�{����f������\a��Y�R�|��OP�(s�5"���2V�����F�gj�ǌ�m��u�������UsF��9k3��s�F{����p��5�W��TA_��* ������"�
��W�����Q�D����+�b* ������ED؊�+�* ����+��TA_�"�
�aW������ED��TA_�* ���PVI��r5�>Z�` �������f����$��UB�%T"�DQ}��R�P�D"B��dU)HR��@T�ATR�D$�$UUIBJR��J6a%"*��R*PU�*���R�I(��P(��R�T�*��*�R$�	@I*QDE*��^�Jv�ID��$*EID!)_lT]aT���ԥI(�QR�Z�PAV�J*Q���T Wl�J�IJ����)�   ��ln�t)��ni�u���w:ӮBv;��mwY��V]����]4�e�a��(wb��S��P��v�B�Sr;mM[gw]kC��]'RU�aPR�� aH��  �}SA[WvՕ���m����뭲��=�yi��c�
5Cvl��;�6��r��;b:f��Vë��8��7q��PP�n�d%UJAF�k_  s�(P
(]�n(�(P�A���@ (t�0`���
(Pܯ��(P�
B��.�B�
(P�43�.(P��@њ�um.Z��Le@�vÚ�Ψ(��!	%T�$
)$�*�   ����n���8�k� i\�]�
�n�ԫ�t��9�JkJӻ��5�t��W��J���B�mFT�N黁����A���%T�
�EP���  g�+�{�\0ѧA]��ik�E6u�΃������u)Z��Ғ��SN�.vB�4�l��-5V�э�t�v��2�A��v�R�֩%P�!_f��U;�  ����î�䲀�Zj��飛(S��[�wX$v�8�[��P�w+J��kuSwl֝C��h:kKb��MC�T�è۷]��6Ʃ��v��)"]5[j%   Cx=SN�v�"�'B���5�Y��Tv�-��n�[��W��k]n�nT�:�w� ֻ:]`;�i�ZT���Ua[k��mCPv���E�S�H��_   ���
t91������  m��F��v�j ƀQLcP
���)F�:C��RR*J�(�TB"��   ���Ti`��U�
4j(�qV)A4`��v8( s+ &��sVT�Vt��J�UT�P��HH/�  �z� �e��0AF��� *%]'U�@Ь�`Q�E`ڀH jcA�%P��S�0���2��4"����bm4  O��S�   j��1�U@ 	4�&eT�@ O/O����u���̫ؼ�w�?es�N�O'�|��<O|���?e_�����$�����IMHB!!��IO�$ I?�	!H�B!!���~��k3��_��4!
�c7&���qД�J�B[����\4Dh&���*���r��/\�T�7�5X^�W��:h6���J�� ��xn�x������]h%��u��c8)i���ջ�Ԓ�#�q�jx37tKn���r��O)[y����M� ��Xӕ�چ"D��"eAJ�l1T�ۧ���1��r�nJ���?lL �F��������Z��Bzk*��)*�us^�)�wӧ���kA��z��1�e�T�ix��J�o`,��"��4�*H*m�L��U#'�z�f�̼ѫ(M��Q�)L[I��v2�ˁJ�8`�w54[6�m]�$rܼ�G]3��@������Z��^$���қ��6��]�4��B�'��+#���Lڊ,�3J
���'��+F�9Z���+Y��
�:���|𪚵�@* 1�Vhj���Lf��f��M�u+-|�gnR��XV��<j䁪��4��jN�!MYH�������Դ�����H��H��/0����SL�:S�b��m�����EN�^��X&P9RP�������(��Ř��Yo)Ccd�{%��Sa����G��=Y�Y�;	��DJ�Č{��4nJP1�
�b�6���%Z[I�+/5۱X �YI���nYyn�ȩ��0�N,�,�;P1�큕4�EŘ��f���*�u�?E����vr�`m�Y�j��5S�J��oD�a�ߦ2ެV�S'&��E���oZ���E[d��t1�����4��c��,)[8�l� H�qZ7��Y)�_ګ�����J��%XO���ciԄ��LZ(�VKԫ/%�ںp��=n�)����]yFV�6��ˆ=A�45���*���8�]l��(��a��0����\{���Ty��7Y���YZ!�uY�6n:%�,9J�U-`�M����Ln�D��e]��V��b<w���
ؗY�{-��Cn�f��WKr�Ŵ��k��XJ��x�]�)�Y�(r]��YV���7R�h�vؽ[����ɡ�u��4i�a�Jx,��IG-!��vݭ2����36凲K
���d�̉��[Cnne�脰[WL�@m��;Xuӻ:��+�WSQY�f��5��V�Vc��p�����1%��`��[ZT'@Vm�Ww�� ��u��I�W�IO5���)or,[n1��q���`]��20�2.�n��".JKv���I���u`���]ӫ`iJ� ��=*e6�-a��2艑��n�نg�1B.<	6��^��w�aF��[uvLv5��[E8KY2�KC�=�J�ڣ��qaXLD�m��h�/oZ�w�0EbXS�!
x-S42��y��ZR�܁�lZˤ��٥1YT-azkS�kq8n�R��*A�̲�q�;��cݼ�j4�&�R�xeZP����ҋ��x�m#�qd�Xo7U����h(���op�j̨�jKT��v�aUb0����h6��l�6��l�;�/e�^�\I
B�MGv�ԑw���^H�*����qs�(6�z��f��DOq��bxE��)Z�-[Xtm�v�GVK-��U�c8);`�9C���oa��N�̔�l[5��^P8�Ӻ �.�Ѧ7i�Y��=z�)E�v�l�������f��/3dKmQ���-Ʒ$��h]*asAV"F�م!��ī�*��q�7Z��u�����`�X��ۥ����U��̗��xEWoY�j�˙� ׭ڣ�
m@�:��V���2�7$��6�[S-�Y7^���Q�u���4Sװm����	��LS��Sy�����1;�Zy��l�yt������]�M:v��q����Tl�����v���˱�q��ym\����{�}��������)T�n��9.<V5ֿ�70���^I����5�qR�顛�� U�$�2�Թr�\��qk%�oS�Op�U�*ǉK�m=��D%b�"��	,Ŗ�X�i/st�mQ��M�[�ٕ��f�Sf@e�cTD��ZA��v޷�*mS1cr�h��ؕPe�iǮ�T֤7[{de�h0c��Xe:Uq�Xr�f�\b��ba�n�r�G!ih
��^���%��	M8��)��է[�\x�d�Wy�$b��@�ک�f͍:�K2�,��ͳ0āD�" 5	���uy�i�!��%j��ܚb�77h�bD��e���D�Q-mcݔ�];�n���xXf��6�.����ݣWsyMS��U���
71�C
�&Q�kAr���*��?#��XLa�:*��fL��L�j�D��Yv�;�Qr�Ƙő 0(#�ɻ�ɗFآi*:n9LB����)���j=PJx��D]PݥN�;��J�[ h�x��][Ԍ{%v��ʂ���d5��b�\IAu.���n��
�[Ee��,F�؛��
!�l��f7Y�fI�p-��*�2-���ڽ(����-"�+(�:^� �paw�Ie	R]Z`��[7C�vl8�H.�[N�\5��d��L55Q�q#1���S&+����e�Z�Ji�3S����:͌�w*���kr}�_����L*6+.)jM�]Z��ۈцk�L#�t�2�T(^JF��S;_��,�03��!f'V756����h�m6֕ݻ���!�Cn-5�255l���!2)�����e -Veh�%Ʒ����E��	���Чj���l[d%0��%�*n�YBjʮYc��)��K?6m��d�V�9J�-ܫ (�ύ��*�����z�Պ���{B��ۺJ(����[�S�ǻ�n��R�[;��և�8��U �/�Q�#�ܬ���n�`Km�)b�U�g�jB�H�t#sVn��л��j4�ԩ[�(�B�^�N1�]�9)���� ��+A:I�Vka���l=m-��kw���3�^�1� ٧��ಲ�@��PJ�b�n��D ���K�I��>ө(n�:3��*\ux0a��m�M��e}Z�Xl�ˀn*A�'YUe�ʵV�N#RI�\�%кF�D�dpʖ	��Tke�̥*�\j,����r����&!���.�9B���`���h��X�{v����Yw[MaiP�	aRQ�.đ�$/[N�kwkj�=5�k]�m���z�+,j0���b��Y&ef�Ȥ˽�u�;C�H����Ï�d�i�/E�4�ۧ,j��h#m��o�U50�����d�����	�#3+p3��ڗm�Źl;���]7B��hy	blA��'ٚS�'I`�WB�"�Vj�$k
��A�ר��pՋw{�Y�)���5dmm�Kn:��:޷N�nG{a`N��[���Vk
Dӭ��ʵ4
��f����#a]:w&�*�eM��Ҙ2�t�@;v&hĴ"��jT�,�����E���J�J3"�T@�*�A�kpn#Sd�%�B�d.�V��P�kQ1��i�Vآ�<��^"޳4a#Y�@�ŗH۱�#CoFn��ޔ=F�F��ܨ�j(�x��S	����]n=�[h��'�3&��J\�/��|3C{ٱx���E��5Y��B��4����v*���ZՑcC<�0��=�"�]�-��k0��.{���K �����{�Mw��#�)a���Ã&EH*i�2���{�јf�f�24���8�uxҭXǕ������&^Y��a�mA�Z���,��b��Œl��Қ�7&�˷�,8Ӵ�rY�=wV�;T4�8u���eH\Ҏ\%5���6��i��,ܦf�ԕ���K#b�I+.�i!���b��;�vK$�sF������.|d�ՌU�
���
D�I�]���
ՙ�)�wO.
���0�,�m��y2]ᣵ�E���NZ�ȃB���QRź�h���K�ʼ,��qb��]-;X�Q1��A*J��j���u��,v90���B�R���v�+)�
���f֙g^J�16Y�6f�ؽ1C*�b��ɤ����DȖ��o "�J�dCn��W�խ*q����A]�T��)�n��[v�Q�d��YBiP�#��kkpD.ɡ/lcoM� �ĵ)F���L]VC����X�W"�N���az������!w�xo�b�c%��ʰ[ٺ���Jօ�ǘ4!
�����s�)P�s	b(�Tk�=�XՓf�V��+ Ut7^n�k �l@���r�|��b����h&xr�hȂ��YW@�V�fO0Sł��&��AӖAʸ$2b��F:<ډ���Po.�n�ص���ۖ��h�WJ�2�%撃���#���u!k6�X��'���[�c�cQ�YwK&�Β�v�72��L�F�Ke,d�YŶ!X��%<�Zb��H[�j�����nK���N�����h�4�悡y�]��������-�W�J-���1N	�N�]ئ��Z�w
�w�c͂�+N@<�(-c;��dU軚i�uc��F�� .�U�Z#5��CXH��j��p;RF�Y�J����Ǝ��ڷ�t`
�u&�9u#:��RA�Q�q��R%F|����2��IZƧn�� �ǩZJ����ylYn^]'�
f����6��̃*-��ȭ�K,�FM�ٮ��E��\dØ��B�t�M��Sb�,��֢�n��:��������U��n���ѷ�+f�_0�
�D�<�� �Zv:�[��Km`AR˻x�S/`$7����ã/m]�+ḃ(�+y��D
zEJwC
�=��r�䢩|,Ճ�M���h�b�7p��ZD�)�fRƷ�nڧQbz9�N����J%x�իk6��v+��7f�էQ@�*M�b�,��Hm�M�f�Jkv&ҡ[$��Y��ۡJ��-������C`���i҈��LchjͽɈ_�JTj6/lh�޲��Dk��lFؚj�j%lA��w�
u�Eم-.��-�UĪ`v%ɐ̼��2����o �����{�QV�-�p0�ʼ�{�cX�[�J�Q:�7m��	&�f�d�R��[y	"19��M[GTf�ha�v�6�+�[t�	�U����Ɏ3/x��-дb����SU��ұHh�v�a���v�4Z���D��$)Ve��+Ya壥1��7�Z/;�t#6���72��T�h�\{wXkVS��T���*��
Z��
��Ʀ�݅R8�E�q )��^H�z���Jٰ�ʐ<ݥj�u���5�Ȧ�AS
�[2�Ǚyr�AK̄e��M���X�n)Pwe��w�UK��U2eǱT[��ik�[�[`+H��� n��L�=�ƥf^3��
�L&�NңlЬ$iҐ��?X$#�pۺyf��6#�F��ӎiW,E�j,�d,޺2��)+b����Zv@�@�7����24e]��r��/oF.�t���j�-m�B{�-�k\s[�;�H��:iѦ���H��U��9���J�Z�2:���NV('J����ډ�
�5�X�JΊzv����`M�)ѭ�+��V^)��r[;p�c4���GDǁ55�s>��.΍��AX��w#~K��ܖ�n�,'`e�d�U�����k4���1��1T�v��Q�V�9ec���"
���-ꕠ���wl�*J�,�N!�v ��!Zu�m�+TM�j��H�ݧS+V��Z^K�����=!�M���RB�Ȕ��tն��ֵ̈@7��l�p�a)J�>ۢ�����̷��RٳFJ�1�Wu)m���K@�7����8�fh�ӻF;��:^e��� bZԽ@mf]�sK�u��+YW�R�D�/RЁ߶�H��(�t��GVlz�+m�@j�$F�)�,��M�$h��Q��[��Z�Zt�4���D�2U�[�(쉻�ر�
�t���x�9��2���Dvٕ��GFX�l�eٺ��v�Y��X*��w#�ʹ[���B���WQ#E=J��U�j�Q���z�;.�l���!���ս� r��A��ӎV�7C� ��lf�}�ƙI�&%#3%#Q}�^7��B�U悬�ܙ�Co{O*\nf��S����-E�� �jUiV�z�X�̡v�Pڳ[5)�0^JBB�*n��5��"��b��U�'&�\	e%�7!���Ġ�!��M�L�>��3h<l���0���<5��ض��XJl���'�<�Ec�k�v��JQ����4�/B�XI ��V�5`�Ŋ��q������hf�Ѐ7�pAdV�.kĎ�Y�L<�t��*�v:!0�$$��3{M��ɩ�áu����
����o[�vZ�R���rK�aX$5��jn'�!sdVb�eXiU��Y���5i�2�8���I���@� ��2��ŃVՂ���e��ө��	�v��ȦT�-&L29f���c0,I0�f��%ݻ�HD��r��[A������b��޻���f�Dc$DZw��	r��MfP�+fơBiE��
4ܗ2��_[N�k.�������D��g��~.]�-q���d�+�M`wO^�����JN�L�ua�x�fcv�ʏs0��N�c�#v�:���NZĀT��dk���nm�AJ
=X����tD�mR��1��n�����̀�dJ̼�Ъ�%�md4��R���Wm�c@7�����Ӆ��t�eM��2��wI�����YNܫ˅J��W��soV��gN�XCͪ[XBe"-^PN�� 7Ң�8�=����q��J���P�.����o9�r����C���|*�k�/q��8�[8��˚;InP9Y���6��v@�ͳ����w5G�'q.-r�g(q$��^̫ƅ��T�4iO4��r���m�E��֮4� �6�R뫨}�5�xe�W�3;xp����3�2����}ԅ��.����#�u x�+"�]��`�T��ݑt=c�T�;Vl��Â;��(}�h^��z�`�p"n�uv�$56��t<qE��=�ޕ��،��Ɛ��ݮ�n[X�%3\���]����!��Ŕ�ǇN��Kt,�{VIø�4VwDή�D	A׉��:@�����/8��]n8v�U�Mrc\����̻u�m�-���׫e���C{�s���]�n�O��_U�y9i�Z�S� Pf�+T����� �s�(��"��ⴻ�vb�n�Z���s\�2�Q��C\e�=�.� ��aV)؆U�$� �d���'u�z��U���	�F����ژ^W��|Gqq����8���7���>��ok@��ʼ6;U���S,r���.�%���������O�+��F�;�� i-�Bp����9b���R�Po�[�z+�z�I3��.OY-wh���[�øx<���]HE���%���&��s�Ǘ�|L1��/�6m pWsfj5d�
iT�AT�v����� �bW��ܥ�t�dY�3怗� ��u*p�f��l�?�R��]:F�G}w0��g���/*JU����P�!��e�&�����˸��{!D�i��P��н�Lx���Z����ގ�[�,4>WO��E>���j�s��O2���+OL�k�g,�c��]�]3�D��sWd\
7y��`���B����M���B����CiErv�n	�0<�ػ�7l3G�<̈v�9ժY�Tu�4�f˗`��H�V��c1�,.b�<t��)b���,�5��'^PYV��8��C�e�0β���bXn?�v�V���z�q36V�t��}��[�����r��v�,������&;ir��^f�yX؂�;CI*]��g��9�y�όo,�}w3+�*t�H��W���M|�4��ڽ��r츑�p�I�����kR�BҎ!���cr��Y{[���ҦN7�|%@Ӭ3��g9�6*��jX��1\��,�m��]�W��qٴH��̓����sW��.v��t9gb"kEwմvHSwt9�s�LW���AsT�ʠ{���u�m� i�����N�k���̕�؜&u�]��WۡE���k�ru<�F�id�*g_LG���31_�謠�=�4��} 1���9
�I������W�V-*������I�:��w��݀Wj�i��^p ���v�cgN꘨ŘFVr���ʵ�4v��=l�\	��(-�qݬ�ŏZ�z����s�/2�mp�7�:��b�P�]Mfjу{�j��6��Z�S:a��xv,x�y*f����,оMU�ә�$�Go&���wK�?���8�E�V�����x�8֫]qwut� ݭ��s�0�_F�ô���v*�e��EJ[�xԜ�/n��0�n*Rv���}y�O
NgTC2o<�ҳ.�/���z�Dw	�=�z�q�*����,9��TYLsZ@�XR5������jW}]�����������\�m����zŮx5r�]�I�\s�U�d�s�n�2rѕ�9�}Z�R5Ks�]��+�z$��6�Yh/s�[���{��1��Q�թ!�3�;śn��5���:�{{������t�V�Le>ݚݭ��>�9�9Ѽ��A����	=��������08�u��q��o��V#�gt�I��4"�C�����V���0Y(m�^���P�;�\v��K6E��|���S��]E���B�����Zg�;�^-
��)�DwP�T�`�"$pӵ����v�]0��gF�n�[��[���س��4��Ǵ�tGx���V�W�ts���l���)�E)�Y�.�#V^c��43#d�s��'$���
�a�ofwe�A�b��a�[C�R-��H�8V����c�X�q�Du"ܰ��o<PA�r�����mu�q}ܺ�͸r��˔W��O4�T*��֎r��'��;��հ�=�M��ܻ/C'8��i2J�>atF���s�0����#30�U�lM��1���K';�x�����]w�-r�,�-����i�G,��+�9��SRk(�+c�0Y�yfv� j�r�*��X���2���/{��`��{���퇾A��E�FZ��+EF��Y����S/wl��ybl�,�sV"Y��m���p���
��;���ᗨ��j�q��K�v�W�[�[��9�]�^���ܝ6��p��`Ya�j��y�+� �[z1e�z!L)�5+@=Yx
�t���8�����ˈ����Z[8G�˙bh퍻�|8��Ӥ�fz2PI�ܥ[	���0`��	Yc8���s.��!gJ\���u��`�e`|�o~2�Ń7Z��ŠbٔM.|:����WQ�Xm�9(5IY�7�(R֥	��qN��C�E�p�v��5U��3k�3y��,
V5�����α��@Xt�)��q��}�O˩����������h����;���1��Il��Ž�L��F�[kC�ΐ�6�X}�]3���t����5:/�E5c���<�r���ė~8�.���zԅB�^��^m8ZG�]N���2�4:Λ�����=����N˓�����+�:5oVǝ�bض���5m)A��o	o�Xz�q�􌊳y>ޭ���dY��T�7w)k�t�@�x�4;��QT+{[Ymm]������Nf�fQ�H�]2��Cp��:�>�p֩;�����q�#�K�ֵ��mc�qZ��|�z��5�
�"8��χ4(u�ewAɍ�-R�-����n�r�f�=J��́De��T�^��hg_I�bG�n*�)vi/-t"�ӊ�Үېi]���� έ�hNO��¸i#ⷳ$���ow��Kb�y�i�(u-]�Hs˳X�C/!�2�{`L&������e�;\�]5U�:�t�W��-��X�^+��%sVL����6��R�=�S	v�l��\D���k��)�>�����-�����wr�uK�	�Sd�]�]�fʏ�3
���=�"M����U�k�6����tg�uվt���Na���G�/b��V�v>Q)��g%`�ս�h+�T�<��ٺH�7���#�{u�Y,�3����ス�n�����X�X���!�鴡3sq(��\���}S�bֳ8���Lw*�m��>o�^�mg[.�)&F��x���<��l3p����z��(%���b��G3p�ap���mVN�f��B�jM+a�´��Ş�蝬j�����E����"�vJ[0�R��$����:����-gA�3-�����\x��0]�Q� ٛ,ݓe��ZEͥ�c�t\��m��%(.�d�fQ�V�Y�d[3r�J�溋6�v��	��9W��p]uu�˱�VP�ɮ�K���+���[y��{�V�f=�B���j�fp.�)w�0��-�r��",�]��Ω�EF;��9p.L�O�Oĥ����Z�ua����r�+�����:*m9��,J�-�gi{��c9��Z뻐 <Tެ�ii��z��·#nݩѾS�
Vxs���a��0듻]@�+AaE�q͗}�])=EVG�K��������¶��jr  �\�qZ���Z:ri�Jv��D1Ӝ�8��L���ٮ�cu�Λ�m�.�q�5:th^�����56#��)B�[�M�:d�hMA3��Hlp)k�u���2�[�;�H���;{���� ��*��N� mT�Ge0�x��Kޮ����Vc�9C*�Vn��ǎ��Z�ƒ�����PN�t��drr�bWR�p�m���0ͳ�uM��]�AO��k��(����5��m�ƴ���ɺ
F#��=� �!�9M]
o�vjh�;�$��~��N� ��
�8�p����.���_#��=���(�g6v�J�^�3.+2�.+3����E��4��w�����ҍ��bƐ �{���)٣���a��}¯+txL�o\4?��6ŴK�cꛛu���)y۶�fwcm��Q�3�� ��L|�\��n�]��qf�Z<��|��ŭWTN����݆����9g)��MH��$�V�mS�E%�u���n�D�S{ܰ�Y�A���TWM�f\��Kk���8��̡�鮝�VT��qZOe�qO8ɕ�50Fy�4ŵ���v�7j,,ǣl�if�0Q���ײ��L|9}(}r]�,���\����e	+fe��l�F	ܫ���֝�ȁ���5P�l[�]���m�ғa�-:&����]&��[�;/��MGrݏ�k��%����I���U�8B����<	��s>�)��1;9���纺���{�NO ��wGm���J�f!@�9M�B�:���l���-�Ƞ�@�&5w�#:����;qlA>��B��e�2�jvP��"�O��m`��>X֞	�/]8|�������ݗ<�p��=`�;eLޥ�x���C�%�6b��<ݮ�����/����MM.	�lWh������]��r\����)�hx���u�X�N�q{��#�!���c'l�!�զ��`gAn�+k6d��U]���x�#zc�=�ξٔ�I��5�J��qF�ɇ�<�kQ���4M5)�U��GTR��K�X��.U��H�}OM_wh	f���b��@�ۭG���;�ۼCqkf��l���3n�gL��o,�!n_�E���ŞW5�h��J��Q���R"��xT�j���l�a�j�tO5��w�#�yد�EF�"SA�5Zt�Ve�yY�'c+n�Kˤ������]�k�h6a�ZhV�W!cS�]������b��.Ȯ�ΗJ�cW��G��q��h��n�s��Z���1���6X��!J�|�����(c_=�m̷ܻ�����]!G)C)�-�սO3Q���n
=Zn�;���nr���?m�J�+���z'�F/g&K�= ������� 3���r���V���%r���әl��):ً���Σ��t�|���!�s�XW#�̝t髨��W�o&r���P�7��3�r"�����We����y��N��:mt���F���B�n�$<�r���y'v�s78�C]It���FJ��[j��L�k��{��;�]B�S��/�
�b[]/���lei��@=3^
E�NЇw�dR\��V�����f�'kq%�/h��w�ꮰ�(��ĥ����F�_M��fbp)�.�u]�g�Wj���:���fR$�P��mF�w=9/E�h�O #@�%F1�<��%�Ƕ�,WG�#�Y��[(s�8�[��%@�-#v�:�3�qb�z��E1��%m,��/�۔���t��v�ͨf[�A�_7��tΩDk�/��gu�Y���9F����jΚ�̹���V9���\���8Π�Q�w��<�f��/�S�ə��9\��]�Ym^Y�+W[����J+9r�tAh���r_4R�4�F�N�Ve��\7�0�t�Y��}/	VUaX��W"� �����JW\0��i3�W*A��.���,�\�q�¹�a֩)n�c�a�$��=D��/[ֹ��2��y�J�7�X��5�e��"�I]sg�GKV;��B��LOY
��净�"���8E�GN*E�]������.bE*��-�O�ޅE�;��salZ�>�|$�Vm��[w��RuJ�m^�x�������u1s��Ǵ�e5E�Sd����$x��y�1kr��@Y��T�õ�U���L�ǌ6�xؒ�"�tx+ゅ�a�u	ޝ
��t� �wQYuyձ�J�LĀ;N�Z��Zn�J;S��**E-I��V��ʳin�_o9oN]��WZ=Z�:���^�fŧpN�`��YU�U�͛���Z�4]p=�o	@�f��V��1�A@�v��ٮ��Q��s'����8'W0�1��s.�Y�:���@ͼtF�ҟkmn��jK;�u�6j�� Y��A\��1���{�܆���k ̨��y�����v��]�0�F���`7�)d�֪D�ZJ�g����
�.&��]w������*ڻ�:�6��}������+�V����4�CNu�uCڌz1Tb�r���{D$E-�̌�Ŋ��nU�Lhe���*hTV�&��v�
u7�K���[DII*�5���U�l�oZ�KD���]���)BBe�oM�\���@�tԸ�wI)n�F�d��&)Hnp��)R,����=�Xg۔��4�֐0�1.�R��n-� ���)�͑Z�e���1m�t�E6h��/pT��(�m�!L1�֩��sk�4o��iu7�����:��]-y�Z/�^����y����yK`�)�(#EEY��ָ�o�^+�`�������%K�q�ד�λ�������3ւI�׵��5��#��}����C�*�h}��r����u2;�4os]�N^u$I���(A���ۯ�4y��R�g,U23-Ӿ5gx�4EX:�R�j4;���|,�S�:r��)�d��t��T�GWOb��q�RBͶ����Y�;Cr��d�=��t��jQ|2Q�����Hi�ڔ���RP�R5T0T �bEQ(�R�b��$�yX��ݫ�*H*�ܴ�W��6��9|.����M�S��j�����BC�!$ I=��s��;�<���������� )���s00���=�//sz|��S6v�8!���#+b��a�YH�n�2c��S�9@�f�q8*sd����}�豎«U.������	ɸ�i� 췋�+�F���às,�HΆ)%��ˆK�g�o�*@��-֥]�
T�N�Ɏ|H�ƟҒt0<Ҙ8����-��_U�yؐ�ǫ�ɷG�ȫ�z��Rؚ�M�#����%`꙱#hT�#�ʘn�O3�7���3����s��4wqd,�mY
�_;�eᲝ59^Z�/t���	j��9�D"��`�<�ia����V�;/Wr}l�%eA�!l���G��N�d˧/{(� wwCWwGz���]b��*�h3`�`�68�
�yQ��XSr`hOZ9ϻ�_1Y��S�/'w�Ġ�v� 1<�ͦ�0���9�^Ш3X����� ��3�<F��m�j��v]b�7]��y������/r1�J��t��l	,��[j��dȫ&#��2J,7V�,��D,��`�)ƙ�����7�B�Q���}�ծ}
�x����^*���Ʒu��fj�K�ѡ�t��^*��ڏ��]N��2�6uKtoCSh�U��R	�R^���"�U�˴���|�����q隰�6�s�pe����AV��1�pӅY�ʋg�s��v��L'VX�f��RqnM����s�-倻y!:����Y]��};B�IB���J2�v��1��u�т,V���w7Ia8���$��$I��=Ԁ�Y���p���2K=��V^Gjp������s��� �d��p��+�۶�s�z$
,�gQf�}��;Z�4�^7O��V 2�*���Vr��QGV�T<w/k\����d���Hl-PP���X�.�ػ9�eZD��]�n��6�1�에d��׎vch=ŭ�Y���A�����́7F-ˡT#;q�q���V��=�Z���F�б�n숶u�5udŅ�p�I������mi��'J�t���7�{��5e�_r���F:�bP˳G�N��Ε��T)٭l�ڸ@���yu}:q�f�����;m�4�B��si�*V�H��\t�T2P��I��mou��K{8b	U�<�;3Gr���]�oH12,�yc��g�f��B��c5�2�"�x�J�v�Čor���WY�(e��+uY���N�PލV$+x�x��ó��S4�$�<�����u�tN�Tu:��^L�q�@X�V<�u�Y�(��`���kV�ܫ����C.4 ��i�W:+3o�}��y[=لm%ȻT�N�����v�]�>�� 2S�fgdoM��.���J��Nb�i�!$�mB� -w�`Y��	P��q��Y���lڑc�G��2�:���X2��ZV;1-����Q���u%'3��Lcc4��j�Ǯ�K7����׽���w���'Kap�5Ϝ.�nX�~��'hz3R��L/W���4��đ}��}�)��{�=k&��9�3�;�X���I���;j�S�F팙�V#��c��̷�Ԕ(��v�wN��.�V�k��t����=E:�`���TR���3n��/2о7
{؂�8h͑�)�ɕ��տ	L�ٶ��&"�J��S�Ӗ-�.�/���9F��Q��Xn�v���ӠJG�q�!��V~��9�ՙ�ݴ��3RwE��Fk�u`�C:c�2�2n�X�u^\��ʍ�t݉��zž�Pf�[�%^*��@�헽ʸ@��I��e��Nvt�����
���k�����xqj)��c���;S�\u��r�}u�/H���<�g��I
LC��*:3m�e�0��N�\�
z�.��2�j���]��"�y=�8^k
��Ml�}�5e���DX�;&��I>Ce�c떫w�&h�B�uB`[��՟ࣚ�x3���0/ah�ZOyr�j��#�_�/.79V�VN�q,�ڸ�w�aH�!���7hP�&߻���`���5�<�5�u�����0J��|h�Y�̵˦F�׬�|����%�v�o7��o"�pY�����;t(������ݬX>_l;� Yox[���u�e
t�Z���j���,���M�E�Ho6J�y�����vYS���ΠC�++��W�,�!����s:K�֗;e`�ʠ.�M�i��&��x����=����Oi�L��
��[u�K��]8����.71SWY���EEt�-Q�ˡq4�b�|9_v����yNͫ�pͨ��}g�8�����F�&�_*��bkj��̧oy�d�شpA��-�dZ�ξ�$ޣc�e��5��e��qʏf����n75>�%�眤#;j��[�-˻���z]���ģ\�rJ�L#���Χ��!�ٙ�w0ņ6ӯ,ABi�AjQ�n������(Y[�&yz;	pɮ�J!_C��Ł���+���.+`t��s��R1���,��Yxu:�\i{-�N�b\mvԶ^��o�XGԨ�#u5m7���G��w�n��E�br8�I���;U���d(s��.�Eܝ��Uu���9�:˛s��o��t�C ����Y굔�C�`yʮoa8�T	HB�ݕ��i�V*��	H�o�4���eG���&�7J�=�D�9`��V��w�[�r��P=��j�AЩ��8�쏴��R�w ��\�QQ�-���I�f�Oq7k��߹���A�mθ�^St:ΊRa� w[�cB$�����˚h��b�4�Z�V�b��Y�@'\hfR�Һ< L����T��+N����nУSq�����eΠ�\��7�՛3v�����3�:�9�ui�u
*pO*�cT��G�jgV�۔�S�;ܝ����bJ��mκ�K9�e�_^l�tJ���n�m�p{Yt� v����H�7}�*�*���2i����U�f7������Z�1eU��-� QS{DY-::��sC?KF(�8:Spc�)�r�wa�Knص�Z�GxG�[=C�jPrQ�;�p�)Yo���R�f2�,ׯv���hp���G��m0�ջ��d�y�-�!X���]�ӹy�F��]J��]hۗ�����s�����T����҇�&,�9��(Z�.�T�/���ظ}G��_i����޷���T:=�n��ƅ���� ����̆�":��+��j���vV��_N�+��:롬�Y���f��S�(
[�ڴ�F�FL��E)Q7�fi�0c'%·.b�i�/W�����π֪M�l<��kwJh\�9���r��)W�\Aĉ���� ��NQdiP��]o�U��.3&���$P`�W�ۥL�\Lx����^H�'����=���t;]�m�]���W}�C4M]�)nދ��Ǉ�q��,����l�w�h�m�!���>��Y��Qw	�Y*���Q����9���Y Y޲��`Fd��X�2��ي���qйVŕ�t�7fZLT���T�Lw�hكG͸��)��NXn��h��-�?VݥY�pa�m�*z��X�V��s�ʱ^�թ�\��_�p�!�6�:��<�N�䚕�h�`M�΅mcmѣ�s�%56ŹY��=��v�O~7:7W��Ԧ��V���r��q���px~Jrt;ص?Bh��7kGmn�
�ޝ���4� ��"��K�|�͹o�B:��s�dmE	*e5+Y琑�u�۫����G�E�N\٪I��,�O;;"8̚�|F�i����5�+���ٵBXI����(�u�RSN.�.�L��捙�_]��VqĭV\=�D\6�r�-"�ӆ��$8U�t���CI�uo3R�E����.��Y�
���Ȑ⬾κe�:�.�>y���DRVa��If�˻����Q�h[?j��n_f���vt�}����t3K��޴m����"� �#Qh�[s!�5:�J�9*��Y���>�w��R�^"�Z� ���yO&�J�6��,�ldA-��:x�q'#�s�V���1J��vj>�oE���E�z�u��n�/,�f�街���k,�rTt+.��ӗ�ZAUu�׊Q��Q ���2����eYz�'gP5�U�mw;��"�k�u�4Cɂ���-+�M2�����ʳʦ���қ��꒶�qn;�S%���(W�w�EN6������u�����[��U#����i_s�>�i��U�R�%�����ƪ �&J�Z';��g�o��*(��ò����Ƨ�B���;��B��2�"4ZsH�J&�Q���^�.Cz�He��Ʀ]� #p�}������3x���4�Q0���u�T��z�I]@�+0���:��چV�,:��-X��*=�Jx�=�Y��}�)*K�p(`p̦r��)�-`�մ��R�E�������ֵՁz�r5��Y�� :���-9�E����nm
�Z5�[�;�lat"���u2�!�*:Fqtb�\ݫ
��'^v��K�����	�c�����w�[`�KPҊ9KɀY����pv�(mi�\�q�:��<u�]�|�%;
%hu�k�'��嶀�_n	��<�`�ٜt �|�L����7��inT!m݄���FڸXd�wi�����8y����ؕtfJ������=��-�*�A�����]wwwo+���:�M�gr+C��YK�+���;�\K���pr�o\�sXmR;��=yWQ�:`vͳǅ�F&N��b��Xr�Ʋ�Tj�ɏm��OGW�+�f�/2tx��V&�c!yʦ�a�K9���p�K�A�K���2�-��2>��c]��p�ws*��;N��ޮAw
��k*jm,��,���J-妄������ȃf���p �<ճ�ǶHT+u�i� ��=d�d�WS�Ƙ-�c9R}�b�O�e�Gkg�uN��gP���܂v�R�/k�:����ͫ��E���V�P�X`��vj�F.���o.۷�=y�k�+v�3 GKzp�]7�t�#�x��Ζ͇pй5^c�u���y�:ݧ[�3S�8���ZK�W#ݥ�=���,P�YuPd�S0��F�{��Tz�b��;w���}�_|q�B[-ےWt<�&lu��SR�
E��_N�:��p�*X����po=�wfV�碹mkΝN"e7PP�����@��n�6&^��}����sqKU��ce�h�ۭ<�-eeL�Eu��vT|��5yt]��P���Sߤ]���U��u�Q@� ٘m�ڵ[ƃ���E8mL��V�db�:;��g��^EC��\�VWM���uʰ�}��Q:�D᫦��硑׆�z��=�š�]�p +�7vF����%c�i�q�%���k5tI��<��3�1O�m�,8��Wt�{�:V�#�p΂}�Һ�k�u����E��0�kT9�^tK�^p#���,7w���aO�5��2����U��Z�UL����jv?����A����u|��+R9�7��[8*ScU_is���no���jޛ�[���r模��#���*�k��[�|��.���)N��n��.�XhwAۣk�Pǌ�o::�K�Slrk�{����q�N��ۇxǅ�7ǖ��Zv��
���|���]L}83�W��0�����{#U;-sV&�]ms�u��5|�Eǎ�X�4;��*��{���k*�b�m���=��]"��i�r��5Y�����!K7I���:����e�K�Z��Nj���L��H1�8J�dˎ�7�-m�/(�l�0�w��l���Ҭ7R��)E<v����}*+s+{%{���C�\B�Z�����4SO2�S6�*<��v�ɧ��D��a�I]>�M&R��+I�(��ۏ�=q�zev�6M��
���' W�X���<�t(S@���f�rz,G�QV'S����N��g~�kMIW+*(_2��)�B���'ۚ�4lG%XF�*|����	��:�+2���ؑW���-Ou���X��D]�&_iv�0]��V�M�2t�F�N��b���}���X:��)�v�UӕĦOI[�6�v�F�+8��Illġ �q�5R-4VR�S�b�+����'9B�.nc�:�3�k6� �y�,J]A���c�۝wjtJk��}���)�4��Ltkpr+o+��,f�/��١��(�Y�C��sJNG�j�\6Cc�ћ+(\1yN�:��4��;	��q��:�������H<]x�-ޛz�t�Y�eہr����ᴥ>{�a�#A!���5�+�Z��R˶�����h��&����V�}�ݽ�v]��c�j�s�Tpl��j����\�>�Ūq�4���Z���y+ik"]�m_�F{3w:�-��q}\,S�a��W��O3 u�u�Pw�|����MP���'�q�����ҝ��6L�cT:�M���3�\�.��w�=qc����+v��P���d�``��w.�:�Ƈ��K����q�L��m�N�ogn,����xa�D���S�-w�X�zgp����:�j�d�����g1ۓ��� �ث�yXn&�ve�*�Տ��D���[K�����i郅<�tv�W_}����K��1$^���d�O�a�$=��joV��4b�N�R�q�
l^��m^Ϋkz\���	��a�֬�]F�0�5��D��N�EʋL���g�+F,���r(s��a@��ڛ�L�IIH�e��Nh��#�M��a)wn9|�v.�]A\��#Z՞���j���/+Y��.��Mڨ1�]��w�d�&+^��8�[Vz�Vh�#�޾��#�6H����S��iу�~��������Mc=k��[��
��.rm�i���f	j�PR��1��/-S5k�����.�_t*�[nn���h�Y@��ƝL�ӮڇH����,�J��7���=���٦� T���.퓪Gu������$^�yt��!8Jܬ}�,��Ȝ9��r�@3�1�i#(��K����w��,'�Q�9�j��/�G����Q�[��-ڷ�Pu�%v�_HꝎs���>�|���3l,`�,{k�R����J2:��s�P���)�ݤ;�%W��s�Q�����ufo`��1q�v�4[�N�Z�:Xs8��Қ���n�V!�&	n��Ё1byj��{�]����hpW��������=�a��:�Q���;f����,`�ohn�O1�[TcF�5�.�-r���*��H權]����Ft����'B��Y�nw_Dq�������3��]���ơ������>ť�[y��oR[�3Kض��ȯ�K{:a�׃IGd!s�*%S^�ja�%\Mv̂G�&�+tE쩶���-����J��2�Xl:��S"n�����Хk��OnF.!ְ{R�Yo^��GĜE을Kޣ���[4[�WŷKEcGQ���sɢW1���wo�&@Č���d|6h(NP�����\7�p���3�`�m�#�8AZ��+��b�p���Ͳ�E��"�b�[hV("�(��QT��+(�(����X"�Z�
&*V#Z�R,P�dDF)S�dP�(�"��W)(�+���QJ�������m��� �
�R�ʬ�Z��b"DB�QQF-�E%���DU�(�,RҹJ��Qq*��X�bµ
�Lj�ET@PE�Z"AEQEb1@�+����V�UVTm���EEUD*J*� �R%,�DQ�b#��9ebɍ"��#бH�QcDPm�Lk�Eb(���F
(��l
1A(1b2�H���*,bF"���Dcm"������,�
��k���H�DH�
DLnY1� �b`�*�U[Z[k,k ���"��X� ���V��0F�b,V0+Dj��V"�(�(�`�,���"*��*��*"�@h/�����R��t{)�����S��7�Wi���_#��t�S�S�3�jK�/M���ky�*u+�L���e.�w�÷�,G0:'��?�U*<�ʔ��uW���.tr�>ױkjD|!�W��1�8��{�Գ~}�����{���JCY�{��˓E�D��� �b�њ���7��t���RGէ_�=G:5�t�s�L�������aU��8F�^Gg�7�E��� G	1����3�G��U�>��q�?-���QMWi�\*���P\a�yPK�w{M���Jb��M�C��(g����x�ޝb؆eg�(U�d�Y���E�"	L�����j4@�T]O��+E��:���}��R5�]R,G9�A�^,Xr6�s�1͕>Lߜ���<�^�6�w`U�]˕�z6b�S(8�FFCu^��wW-�pln�Bo�l BH��E�Ыq��2�nj�[�O`��3\Ҝ��Y/h�j�ߋF
}>Uc�T�|o�q����\�����'^�Z�I�k��/�,��ڼ��a��%��&�{���Hw,&�'�x�@��f�^Mޝv婝ך��c����
.�=�5yn�>XR1o]�=.(@<�(v��IZ�`�-��nIW���c�wg9T	�qE}��}+�]5�V�YaN���M7�o����J�ut�賈~�˷rK��4H1f��WTw��YW�#��[)�W(����+��g]o����Oj���*F�k5��Ӑ�;F�lt�ٺf8�Η���B�D�!t��/<��>t�]f��iV�r}^}�v���j=~��+�9��R��Mv����ةp(�p+ˋ�}3�ްE�N�y�AS�*��:f�#�FNb�aZ�-e�xh���y��J7�bj��unVK�����#���f��ҰE]�sO�dp�<F�&1*1�@�<l48�T'/���-�:*���|�ءo��f�9B�٘LG���pjG��9ER��)�~.����8�9+����t�-��{ �Z��/����gaX��PmJ�
p��$yi�
ui䴷��u�s�Dk����v��@�~.�������P`�4��\
�@V�'%O�C���NA~���� iP��9w�J�7�S�֙
�����C����F⊶�v�/:j�A$�;sW!�R%� ѡ��@rt��6���Uk� ��'B��I�_��b�Vj�f��' ���oH� A{�c-�{��r"��h^���݈<�Gn�S�];L.�uzz�ShçF�
�V����f��G5���c���n�R��틞dר�vwU�'c�>�ã��Q¨a�{��������3hf�]ܯeZｦ�5_h_!�^��5\��~6hܾ�w��٥�x�b[�{kX��N����5ǦezལsV�Rx:	�VL��K�9ر���xɼ� ��N2�ػ���CC�l�jU����|0.5Zr������:��uF��G��#]���o.��F��,C�v�"�{7� �Q��Bb�4}4P��]v�{O]���}����3``}�f�Uţ��175!��]�sG���xn�jY���[�r��bS�#�ԥ�z���� Y�=���*˭�����T��Ar���:�N[k^O.X��Y�]��,�M����(A��4IrjEC5[�����p��5�v-I���YQY�%R��}�.�ˇ5^��[�
���s�Jx���6���?.�*�N��u�5-�J���+��tԴ�xv��m�꘺�:m�Ҡ��!�#HE�P�kh���	5;J������ml*��X�Zb�+�T�8���l�K�:�*T��+�h�Ѝ����"�L[�Y��Pz�-�U�e�띗����f [,Ihi[%�"���-�����LzH6�=˯��RN��l#�AƝˉ]�sc��Z�u�K��l͎�t9�����=+mY'5z3���{��o7�}��=,Q��>�<�\e��
��W��t';'�ߵ�3��L�pd�^��j���}SQ�3xaa�\E�o�aq�CV7��s��%7]R��������V��nGC`���]����j�����L@�r�x��PGh�r�ɗm�Q�x�%c�W�s��W����6�X1�@��s
�x$q\lTaG �}��K�
�e�	��_y�b���� 3�tE4������\����`X1�^-�Z���44��\���W�b|7kM�g�g���E��]e ���ipoiX������YL��c��ͭ����ρ/k���Ox.|n� ��F������ ��8��zZ�et�n���0��^]��F�4��cb�m����|���}"��=��N��K�&2l�K��od�ǳ�n��|Ҽ庯ږ�ݕQ��M��Y�wd��N�
�v��ݶ
�����k��CL��j��R��:���wV�+pE�#4Z╭|�]��Ta�>��pb��w�;�$��7��0z�A�6�Lz1��G �H$�57��d�x1׌��b?_t&�����f��C3}�Vf�rB_|{���,�e��������rmpc]=�8����+7�L(^��.Αg	q2Iωߧ����N2��{�rq:��A}���!`�k�z�іW��9��U�N{E��O�`�,l�uVN�9�ǒ�g7^5��J�	Ch6q|¶ 'Aԧ������ե���͍Un\�H�*��jӰ�[%F9�4������80Uڈ^��_�vC�fs�2YN&:(�}jٜ�X��T�1�L�����3�M=<��r�֮�W��y���Zy���S��~�o���ճ�J8���ڝ�t�Th���*�:�:[�,��d��X�π�BV	�҃&v�A���Tts���3�˒��RssU�k�x�eF��p,�Z=!B�"yCm��".�:
"pxN��o0�Z{�3%����\t>�������y. �%D�AX֐��1���du��Ni�ы�n���ůb�H��P�l���yq�\�$��w�
|~�ZF
R��lX����ø�ڙ�9w:��9�P慦E��#�;�!Ł����;�$&X��bX��>��xpE��uڮļ���(��y�����//��!��4)�V�ϝ�y�.�=e
�˸h9\8�^��$y��I��x/p����`S���5,M�1*n��@8�t��5�*�4�.���s��][�a�i�g'N��
�rb�z�J{�.��{�a��p�"J�1�1��j��E��3�QPS@鑾�5���kMܛQy��DښbTz��0�

(FFCw�}�^�G c4���M�7ʶ �����Y�N��#��VZ;5Y��o��� 6P�2�b�"�.�Uc�N_\���`|�=�b�7]���P�k0�n��!��o�Nl�~�	�ڊ�(�R���\%#l�y��!A>�ѓ�7���x�<NQ�k��>��y�fņ�����l�<��ЩA�|�|1e�x�rւW����8�*r��Q�"B��ڢ��g��!9:α����K���1�������%�,��SX�GG�'�e#���֌:.�!T��j�N�x�ΜSy1m�J�ķ�	w���X��0E��P�8�B�h�Lt}A9y+%�ASʖ��aAs��u)bk��pܞ�=�m�=��σ�M�ݴ���kj^��E�Ey��W��c��r}[�R��J�S1�뮫Ct��@����HBV	���W�K�;H��l4s��f��Nu$�i�e���EB�e�Vb�=�IڡMA� ��k��İ7ٗ������(�s�7CmϼV/�+��-Ƹ#]��'x��[�r�V�����`�K��u�b�~���5��M�Mn�R���l(�.z�Ɯԯ��_*ΐb�|z,��3��>
�5G>��P���!�Îf�-�oGrS�����_�8��T�v��NS�P,�.��gr}~l���	Ȑ��w ���s����h�{����2�,)�#��q�W9!\ئ��`�N�.oZރ�SY�	�I��~��� ��u�4,�U�5�����G᪦�N��g9.w���cq��Ro�v�
����t4)��|VqPj�b�� �n}w�T����d�}'(����� n���"�}J��¥v�;\i_R�@}�u';��(lm��ʧ/-VcJ{�=��\C���<�����e��S�W{�k�S�7Q|�����������K��o.Ӟ��2�;�>@��ٰ��1=�����
���	��B�
F-����6r�J���6��z��Wqb�9ۻ��l�͝r/dVVE��i]��Ƹ�ЊM���"Xڋ�P&��Y]r��+"�F���F_���X���"��%1�޲r9Ow[��j�Lu�
�m��+��_D�4�ݨ�V�4-�٠H�vXs(qV��a�����GG�PdSv��W�u��8qWS�y(�W��圫P�N�5�2�7ܳ���He��p��2'7H�W���'��.6�sśQ����͎���2*��,S�~�%I�T7U���}D�=�^LTU��ڕ�\V���qdj�z���w���d{��}�bܵ�`+�Ӽ3�^%{IA~��������s��/D�D>��B�}��SXH�KJ�����@rKAJ�֚�6��nH��+�dw��[K"�!����!��M��:gj^D�M�ms��/�T�j��;{��/�%jｵ9~�H�*�e��vζeF>��ኁ�Q�{A;�|/���b��B<�.	P��Е
	�����v��	MŗCT�N�Cv�ɔ�M��$�8�K��P��?!>Y4w�h��*�?P=����$ˇ���a�].Ck2��n�w-�ьV��m�0D�h�� �My
�����ǔ(ծ�m��o|���rR�;v���ona\�ˋ�T�a���Mh0��h{|�E�{捭9���S��ܛ��[�VM�y�Z��N-�d#.JG�8-u��>"�i'��U�مިl�OնH��;޼Me={���?Q��v/<P�X�r'2��jY��7�*1�R�~)����g�����l�Q�D}2��6�N��+���
�-�y�_u� �`q�jc�m$Z�����Z�~������j�ײ��-a��t��.X+��)�
g^���G:�-d�g�3+�v�P+F��s���2���/b����ħ�Wt�E�cFPS7��9���;�:��[�ޥ�N��w�Az�!�����U�tpƗ]�/$>�[�PIt��7ˍ >��N��5# ��3�\lXօ��w�9�S�dЫ�ĵ�8�������p��j�N|4L(?Z�Kꊬ|x�V�']7�	�z#%:�q�ST4��{����Ѽ�{ �}��Xe^ŷ����)�8#c�H�]𠢀��-͞�i�=X��r�M��g+`>����u���*q�������X}a��Q��46��̫�y�`�0��F�p��\KS��V��ΑNU�`�I��:��R�P�roN���v"��7��z�p���	�u�&T(Po�[3��c��Pj�T>�����ט����/>�ߋ-��2pY�/�>�;>i�4��t�@���E�W������\>�5�����n��c��X�L��b\Lj�i.OT+h.�||�k��;S:ѷ�s&x���b',����R�A���\���:�����Y�d^p��LM^�VS���ʗ��b���p�_n\£���GA�RU�1�#3�B�'s�ֽ8�q )�?���r���0c���/vߐtC�!�]��v�Qt��4��c��z��u�FlW6sۗ�o�;�e����֩@�!*�T�C�R+d��E���"r3`������݊�Js�W�q��<�����y. ����VG��jz�uӻC�F;F������kĈ�����E8��'~$.3ˏ�;	WN���~��e&BtbS8�̋O�P���eC�jоdQYב����ƺ�/���� &X��p��I�J!;ϸ�82���ءT������`,����e�A��XF܋����/e��n�������������^<>G�+iW
�c�K�2Nv �E���>4 7˓�3/�ڢ^���^�ŵGf�d\Έ������@�(߭�Oo�
��%Ծ�r�R��gz�Xu��ن�`L��PY&ޜ٨6�ɒ8]>�Fzf܅��7��v^b<���{y���]�4����dc��Nw�}�����l���IU����o3�̻� m��,OMAS���b$!	M�j���L����9�##Ch�R�z9qqy�S�bj��"�v ��$��i؛����"8.Cؓ7/�k�b�ŋo)�wjI-��aHk�d�v�;��y�kU��*�L.���2y�Ӟ�Fk3v�}Ǥ���5r�g{zLD�\Wj=����e�N���^�V��r�Ծ��Ӧo�ӔB.`VK�z���WD�V6�Ny幼�k�j����
u3�lZ_t[uq���#��Vry^9O���r��1�*�x�"z�/��݀��r�z�^(Sk9b�f��O���IɨeZJ�8M%A�eM�F����|֞�9>o�AjN�r��eX[��v啌M -���v�:��{`�J�@e�v��N�ދD�le��B�:��Oݩ��h���"bh���3��)�Ӥ�4w��M	�,�
����C��+�������9�%�A1lo�V2G%�\�.�!��t6S�<gNa���V��M��s>XwQSn�i����U�k�W��mވ.��p�����K��� �T���n��U�V`�J}�eIV�������p�_KG���p�T3t��e��dDam�fbA-#5\��\/DgN�ε�C.$���t�y�\$+�i�+1G�,�إ���FӘ_5��v˝q(!��E#����ӗ�i �<���jJٛh��8�ɜ�"����х��k!�W@�J��9�hj�v��u�X�A@ٕ0%�gT9#���K�ePCvP���_>��a�Ȥ�9o�^���S4�9�Ő�c�t�1PpїNG��.c��]�k��Vs>m
�Iq櫝���{u;R����+��]>�̺� ��U��z<�t��/j��U�t��*��vi�(�b!�\��s��6˙82�emqj��>[hZ2©��I��4��*$A�˾	�Pt�B�T�V�#��o� �V�Y{��$ػ�O���a�}�:�rͨ�<�MZ�Ma�}9�Nw�Wu�6���o��k��nwnZ���n^r��r����H΢��Y�msq����qhd\ >��2P�z����u�3����5yJX�x	w��$zv5Po�:���:�>]avV�iG�)�&�U�W^�z`�����.��p���� �kam0nS�&�U�� �͛崶��ΓXn��_+�QƞcE������&��Jt�
�o��us���Y����ۣ���&-��!�Sw7�R�K �
�v;J�&��%�P5:��h.f���ʚEn���e�C~毵�v5�EkQ�Z����ʊ��=�(����� �ʔ�૵b�9�v!6nS��ϱJ�hoTL����G;��̼��C1x�����_�1uM�\��kKzY�q׳iq��49��-�˶=��C���`��%IN��k5&��<�|lbuM#]Eu�9���p��*�����b�K::��w��s�J�;���+Y3�rp�)����\f�P��ޭ��ݓ�Nc���*� ULmP�)l�0Q�1��UZʂ�b�EE���Eb���((����b�TU(����2��1EF,PPQE�
�**1",UR
�UDE"�cZ"��EU�1Q��"+�V(1c���"�Pd�UU�(�PE�"�b1`��DT`��aZ�PQV�(c
��QX�*�ʋDQ`��E�`�R
,Z�EAQB*��Qa,�"���"�EV �����1#DEAUTTX�b,Uq���Z1V1E�����"LIPQF ����V(��`�EUQPU��"�U�Q�b���(EQT�QX"�QT�T�J�G,)��ьS�H�y,�TVR0�׺�p�ӲU�5�=�b�Y�����Mj�%%�s��:+����?eOU����Dp����U�v9ֹӖ���-VՏ7���dtlEڅ�$R��P+�� Pon��&��7;�5���K���NX���=RB��6�(>�����.Wv�_,�5�reU��vdD����m�Y���1�TᯘX�DI�ڋw�cL�=����4�0Y��j�3ˢGo����||��a~[2�%��\�ûuP2�B����ct�́�X����3��~�;2��㬠�s����B�ﺲ��wa]M|�EJ�f��]�]®�}�W�ܻ� ���`S;��ꮧ}	ȟ=����%d�(�z��D�u6 {/GMz�]îr-p�p/˫����̵e�Z��:�v]��%�������C)F�X�F��$�?6��R���j={��efI"�dN�t�f�у 0&�><5x�����U�U�O�l?��~URc�_�����SSG�ے{fX���^�C�����,���M�Z.��S}K/�P��ٱ]���)�ҵy>�۩[��/�X#�C�h���~ʌdn˅�gz/0C�ܹƵ�2ç&M�:̌Hm�:�d�S,�m���v�֫��6�)�g�v�k!�f�û\��P����O1��"͘x2P�9��V���W٬�Dt=�;l����A�\���<��^�nZ�'N&+�,�a��-E]I%��:���'fkڟ����Z��ˈK�����KJ'����	{p���V����e�1K�ѥR�E]z�oj=:ѝ���8,Y<�;�g�o�Bwu1�� �w}>���a������\;�����Z�g��|�!�Y\Z��}m`}*˭���΢�/>*-�J!��[�9q9A���ܖa4[װ1�������(:���*ECw�z#%�D�	�ͨ�ػ�9v�����t_�?vڌS��qb'9�Q-���X�|F���|����W/��:���.�l<���Y�n)���U�Qz�yc� �[/&c�)R��'�����tD�쬝0�[�?Z�&�������9��ȱ�R�zʙt
�)���%�)�C'��aU�U+{��~t��;7N�I�-ȿFZ��JN�;ޕ���_��(m_�0o�d �v=K�t��aY�����0��M��.*	�ul(��v��BSqe��4����X����n�-�u��c�f��u�9'�3���Zѫb���+����������l�u��s�����a��S�E�]�X���כ�4���a���T&�Rۙ��Vj,y����B�DE]&,V�xEJw������eo+��2�wVa���3#��{�KN�M���p*����|s�|�)�(�\>t=����^�ջ�9��4�&Nα���T^m
)���[d`��N$BD��l
���羪���gRɝ}��q�Z��&�V�_�}�z��s�2��U!�G0	}:�׆�
z�MTXDӔ.���y�\a\�#e��Dv}5~�*3��x�{}��g(<�A�_v��z��a�[��{Wj������io?GA�(��8���̯M�a@�޻nps�p�8p8=��[��X6�]r���4���?N*��:�u�-^�,^U����dhͷ~7���|����,��<�[F^f�֊��xS�{�Y/�0,��3"� NC#0�ؼ�B�`� *�JE��߱hoP��,�9�,��I���>.&�T'�����a�}�����=�P��a�n�r��^&��y���(�;e^ŷ����)�9���#�|*�!V��je�hJ��uF9�{���9���%{$�7WQqn�vN�H�J����
�T��1���x�����X�{��S�J����\A��9����7rb�(�J�l�����5Ҷc�΢��l'"�S*V�"��k{�(yrt�%ٻԐre,q|gA2���ѻ*��L��!�1ܺ)�v���ڋ�x�({;7'ݵ�l�6:��@E�;EtW��B0��r!G0�Q�q�����؋�;e��h�� �o<�ȝ��#�~�)蛗
_Y�V9y�@#���n�d�`�ʳ9�,�6�,nK�G"�y��W���Pjp)�4a̅�t��߱ڋ���ү��־��K�������-���r��(��r�W���!w�E/����=t|�A(�9�f�c�u��͚w�E�3OӐ�)7l�u�ہ�-R����O�EMP�-fV|=U8B��ƕ�	��C\m��+a9�t]X�����lމK�(!*&�cW�I!N
tNk'�_�y��a�#����1���L��=�)�����\+�.�L����St)l�.��N�{�`3��Po���o:O�e���y׆x�K�N�		�#cʎ;#n��Y���p�~=>�z{#�`;�Ʈ0������VF܎s0��=c�QWT����v��VϽ�aR���XǍ7����X��O��©9؟�^�X����r�-�P*Z=WήR:�5^\��FM�+zk�a���%��" :P�zP@��Q�Ϻ�+Jd�f�߉�h̏YVz�Ĺ��)�y:���]ٙw֒��_-܎�XS|��yu/X��z��u
�V�c6{�ѓkr*S|pp:Ξ��ǋ��	�?�b�T����x�L	�`7c&O�O��
�$T���C�7�d��FHL3�m���s�:���;0�,L��������A��ɒ8[_`tBո���f^x����+f!
;R��tK�=����.�^F��u�E�Ua)�����WF�X���E��ˢۨ.��G�Ldb\oD�!)��.^ϋ�Br��6T��cz:72��{w���Ί���P��A8"��b��W����j��J]�`�E���?�������(>�xfy-y��c�c��$N9�4�G�`�t�	�Z�*DD&�pa7��e1;��}u�� [��!_��钇R�BtC���X�(*{�rWj��i[�޻|�u~ń(4�ϧ�b�+��v:�o�q��|F��ô�ɪ�Ы޷`�Ҕ�n�oe�/����Q��oö�H1~+�C8=n��&veX�sQiQ�:�����6��U,ʖ/9��Q�UC�S]9�h�
zd��弥͂��3�~��v�k[a���G~�8��]��sYӶ�:�ie$�K���&�!�n��R���!�9T���cK�Û�"�]wVV����XC\����\�0�+]�q��0��k�o���q� ����@�fD�2=�緌���k��N���\�Ü�W�}_�P�7}��pQ��R�*��|>�<�e�!�9�q����E��p�2d����<g8E]�o�7��8"���
aȔ<�M�B��f�����u�_��&z{�@ƼP��'&K�8��>=g���t4)��|W��@5\���a�����{Rm�$�[]כ�7{�w>���@/Q���_A�rp��BG6�+z��@a��j�f�>������7]�W'bԋݣ	�5�1~t�b��= �h�fKQWS�RE�b��S�{�E���O��{�Ѭ�~�(�{�[���ݧ��{6�{(���1Pb�+��F6{5�Ii.\wтr1��*mm���-�e�!��qb�9ۻ�
��R&�v!����A7�/ä^ȧ���!�]ū^��M`},��!�D�SOi�&��3N^��b��p����P.��``n�f�>�5��+��H{қ�]c��ٵ�%j�Ea����ul}5�Zˋr��"s��T�S#��R�F��+�3��ca�~Q{�^� r�y$�m*c/A�'�7(;��<X�&M�E|9�����#��=CuֱJ��K�F>䜖�Ǫ]��n@��E�����̩G�����*�e�Dœ/��E��q�w��Au��#`fv���Ϻ���3Ϊ�c�[=^φ�gM�Um�Q&��W��֡g�+e��te*�*��(W�t'�"뚹�dƣ��: �^�DM�(��*xΩ�!{��])���Թu�-�&����INW��c*%�}AP@lq�sCԩD��܋���_���g NζeD:�6y�.�o�s�^��)B�=��"�ؾ>�j��fߧx�]ŉ��"��%ݜ�r���\�@n�������J������v4k��{���N�m�w�h��Ƹ�x�}r>�u��0D�EĈ(:����l���NX(���lR�	��۵�l9�Aw���be��RrE���߸J���y�g.�n�0'{V�O�>i�VJ��L}4yD�/����9C��E��]`�ψ���KQ�Ý�ySWe��m������tlp�~y�t��w��v�(~�m�|n�p�=�fie�p�s�5\���Բ7S1!.t�J�YX�ᬍ�Ddo�mߍ��|�{�%�\h<��>dJ6�2mf��)\�Sdj�%"&v>�罙;b畑`s}0�$�j�y=���'{g"|�Y�9�!E�Lσs8J�=�k(e���>]B�Ӗ$*�ժ��ջ�f�;�1ݹ1Z����B�+� �)i�i�>�����*����6Ռ�+�64F�ʑ�U�J�%��foV�CfL�g�
���a����(�.��Wtz{jU��ؙ�B���[���Z��K��d������spÞ�
{3p�Xz���U�[|��`�W��I�_{B�~{��,=�H��\<�h%mff��i��ce��O�C��
N�&�@t��:��;�mO'��d�Զ����-美���`�:ĥ;��ˁ��S��P+���{w�x�\��
���{��wMU,?^��Z4:�VR�iUr�Y���ٜ͊j��Rt���ӕO�����{W�.=�#{h�*�)1�'�^
��A8��FAG�ǙQ߭�95�0�����eaW�7�=�e[���d{K�&O��⋟-!��l��a<;����Ri.w�:�������$�Ӻ'nX��*��P�}�ϖD����������(=7\��z�������3�v�:
.��t2<�����Cָ��P��s`�Yr�+3���غZǿZ�{!w-�J�[����΃�b�����v�C~2�37��Ա�vl���ibHE&e��LT[���'1k��u;����"�$s-d�x��'R����/�f�s�����|{v�)#�,�*����)wu~���}]�q����63�UC���:NϫDe'7�S ���)��'~0�qlL�D� �z����߷��%��G�~�0�i��Y�P毙Vu�z��5�Խ��`ڸ��KA��¤�$�$���A,5<
��Q�!䪓�qPs;��mϝ1��Q�*�6�ݷ�3jz@�w?b~Z~i���V�!��������9B.��8cD��]�����Fzo���[ ��>Y{{�H�Mȹ�'�Cc�꜀P�b���8���t{�s�p���> v�������7<#���I�=9�Pm��'�����V��E��īyYM8��R2&2�5;j��U!�Nv_f���]h�~�XJ*y��'� �-��D��{���9E����k񨍊�
��@���ڢ�^��r�"0P�̺��$��#
������oV�s��F��A�i����洊#N�]�f\o�NBT������P�=�q���^
�}ْ�����_#F�vU5]Js�C��\0��L�#N�&�<�	���Zmj{�LQ��G�t(*X)7s�����qaj��(�P����)e���X}���mm�\�բ��;��}�3�Qt���ӏubr�{]���=��yH��A��9m+:�C�����8F�l�[� �=F�*��Oc����WҰK�����#��yÑ�!XRƥ_A���hp!^e˭���{Q�8759ℿom���GA�
>}7��#<D���m�������0�7�l(��5,��f�3���";X�����V��r"��2Y�pL�ʹq�5�7B}QY!��ylfd��^�
���P��;���)�9
�l�����_���b�ܟ8]t��3ְ�(�sy�,�z�B-+�d�X?g)_S:���|�ˇ�cUs��pkz��%������u�-�K'Su�C�4¢jFB� 9�Ң���\U�T�v�qo*�I��Wv��6�L�l�7A@2�6z�;P�hSU��⦫��Q�����wev�֜�Tejj�g�^i�'�u��%�U��o?�`��sZ-�VwV;�N#�\�Nڼ��9���A��w�"�TZ�{�a�Ƹ�-Ӊ����S��a/�G�_9!���y��0e�r{���:m��U��i�[TQ>����(C��|�L���{(���\Z��V�<ǉN���v[�c��������k�c(��3n�Y\��޺�J�JU�ֻ���D��6����#f���Nm\G+6!���T�����;8����Z�Y�M�$�V��ģ ������9ve��oq�v�lH6�k��
�C��z^K��ZĂ�.�n�=Xi���S��9�׬S��c7�"�Ja��+7��<��مʶ��1$��=`��Jh�þ`m�����yӷ
fil���7�n�AB��\4�4_H*;�~�U����h��w�m�˧��&F�H>�tƍ�pU�ҟrWt� �[��e�r�Pw�'�j�7[�Bs6��M�g�r/��!ڂ��8���	-�!]B���F��б:ҫ&���nd�������+9���/yj���w�d�ݗ�,u��a�)�5�y�����ڰ�d�9�x_n�3����.�ۜ!V�Z�O4ګͽ4��ecR�������ݦ��i���b8���ř��B�+�������ޡFeLu|�ql����ھ��E"��:&�D%�Q��ʼ�7N��9�\r��r����j3���u��H�(�w�)�����S�&��V 9��u��-XE�	Ҳ��h�Ѧ�"�B�1M�{Cy�λ������M�m��tЧԃ-��n�U|���[��\�oke�����9megf�W*b6�^7�n���[��&H�����b�d����9��]\�Nt�:�!�>�s30�r;�1�[9�s�����V��H����k:�>�\�A:�ZX[� ���ެ�K#�"o�����E.��J�h���z��nl�H��R��8�ѩi탪�X��]�X�N�9�W"W:.���"&z\���8N�s{�'g�k	��MX�4�W}��y������S�/y\\�3���t`�c���DrB��Iv�ۊʕ�h���a�۠�opV:�X°	moW/��\+��ձ�ܺ��H�:Wpr�t��Q#꬜v��)q�}�4c磍�M�UԎK7a�[���+���f8l�OWJ�Y���f[��,L�r� m�[p�y�eM�젹��'z����M�ʥnQ���s��0��Y�Y2+�qu*]r�R}���R���f�WY����>i r��8)����w�cÉV�AlɓWiܚkS��h���fJޘ�$�Hi��;�$�D�l-�R`"X�Za�}zpa�s&E�7�u/�z���<�m�!O	:���C��}�U*�m:�j�_;�� �x��>2���]�ڥk�n����8[���;[G�����n̕��GI�!$�*���k�o����hAݪɸ�ޫ�,J\�u\K�z��ʨ�-r��d�p�����
�
L)uƉ�|(f���e��K`�w����!��Z��5�+�2�n���w��9�[<����P�0��?5��("���b�+H#H��Tb�QE&6EDqa�m*1PQ�E��",PPlF+
EX�������JV�*�L�YXr�&8�D�(,-(���
�EUĨ,���Ub�ZTE�cTf[Ib((��A�H�[X(#PQE��[@V1E1	QcDf&0Ʋ�lR6�� �-�(1�$DU�PF��JP�*,"����(G)V"*ֈ�d4UPPb���K,� �Q �,U�"�H����DfR�E1�U"�F6��"�7�?��w�����+��|��K�V���ܤ��
�}�c�\o���@�'Z{,�pٚ�}k��@ԙ����]�VR�˺_�� ��x��cO&�b�z��W
q�����)��Vz�O��r�a�v�Y+�M�;�
AO���'���Y�}�I�T+:���S6Χ=:k�y��tN�i9qZ�r�`Ǯ<&@���v�<�����{;�G�Xb,Ӿ����P�9t��SS����!��gY7��=7f�z³l8��z ��J��0�UI�?3�~��x�{�c+
�������Ǯ*<{�_ԅa�:��;�q�M$l���>O�
�Oӽ��x��bO����~�V/���i�T6}Ef�dě�1aS��xn�'�T��~����˹�Rw���Ͻ� |��m�%E�C��2iE�'S�{掠T���S��2f�HV���T�'9��z��i*<��i>d��E�
�}�Ѫ)��a�?q���*�b��@�h���|��&<� J�,��AOSv�0�d��k�:��Xuy���9i��qd��q�����'��'?9�C�c���2k��<��I�|�\C�c�����~�]׷������AM$��"N+*I}�7`i���f�;��m ����m�aQ`oϳI�q�'�mOy�5�ì1����HJ��ɷ��������$��1=�~���C�u�wg�Ug>M]��Q��!�a�>aY�|�� ���sX���T���Lg\a湐�)
��ϰ������H|�E�o�&����o���<H<�T׾}�NЎ������ЋŻˣ�d
�
����{��g�Y1���,6¦r��٤�B�5˖�'�0��M�Lz�Qgb��'�w
�@�6����'���+<�������{*��\����G�{2�r�d7�O�Dy��q'�zo�H)�'�>���T������XbO�é��J��]5���SRc�!�oT�l�����y�4�R�0��jq���"�j����~9w �[��_{�*P+��4��q�P9�i�XW��r�����d��f����)>C���'�ʆ!��}�+T+��,:�H,�S�P�=aQI��1,{� l ��_�;�q�F	��e�n�<����&V.Rkmz�O��L���s����ķ�򑜵� �#w���z�ua.��<�/���cfC��[8�L�}Ի{�:�m��ÏY��V�͆�2;��S�w�VPٯv&6�oA8���]\c�Kq=����mL�Y}_{��I���%�?(3���P?�fOXTJ���	�����E�WO?sxLB����p�;�m�XVx��N#i�`������_!�h��x�8����R�>s���\}���Ç2/��������4�m��
�����C[�CiVMϿoQg����Ͼͤ���d���J�0�߬�l6����w&�E��:���`J��R#�4���7$a�86����W��� �Hw��q��o�Y?2���!��'���{7d�~I�7?~�H��O<�m��
�u}=�$�<a��bv����gU�3�+�J��ޟ~뛺���翻��&�I_�mN�� זzɭXy;�B�m+&���:�P��aY?8�@��5g�4��:�l?���+�&�~�=d���|ԝ�AM��dГ�ʇS�������x��bߚU����Q�ǜxt�^��g�i��TP�;�I�z�Hm�w�<H?�1ꨳ�*�S�RW��&0�j�E�+��<7f�~B�����}�
����?�v�m������o�;��;�>G� ��w�������a���RxϜs�7�B��]�����bO���0�1!]�f�
x���QO�A�Cp�,�q�2c�1'P��,�2�������L�F�f��� �<&{��N!Xy���N���~��mįY*>w�N2mE�wVM��
�����=e����0��9��N&?�� V|�CF�"�S�;���8���s�.�!5z!G�G@���&0��O�u4������0�z�Qdߙ�N���a�<�7���'uOӝ��@����w����%@�f
|������q�̚s��+�|�~������V���X~��<xLS����H,��k'�E ���4$겠���HV}<�3�8�����ugXTS�@S��3�����O9ܞ"ΰ�E,Ɂt�wQs�������7�.�?'�LgOu��(~I\}g�y��'��'�u��>a]����uH,�z�4����(b|�Rc<3�Xq��!]����xì�b�y��?0�be��oI�i|o�=[���|~�ݳ[n�� ���*Y��=4^u2��b�4���=������;�]X�f+����Px�W�Ú�~)�c���G%�+�5��t�Y�fαŃ`�s�7�&N����ϧ��2�b�x&��h�uZ��\�Ե�;uݕ�x{����$��ٟ�<"Ǉ��s���ă�w�bͧXc��'Si?!Y����ɴ�°�5����8�f�d��Y8��7��ҽd޵��2T��d�M�+>����<�"J�/w�~0���������{��'���sĂΤ돜̇�T��'��|�����;@�cr�Kt�Ԩ�5ʪL~`V�N���a�L�A՟2d$�y��|/��h׮h�?k�{���a��&���{��'���=I�'?�z��n}�Y'�d�!�d�$��A��$�UY?0���}�/���~�o�]fw~����Y�1�2vkXAM3��{��H>X?Xb,�
��☇��u�;>�i$���w$�>B���k����+���p�<a�9H/�N�V�>��u�����^���]�߹â���I�ظ������Vu1���bx�c+&!紘�SL<��i�Pć�䕋4�a����T�N�Y���l6�Xi������{�i_�.�=R�nd։ӵ&���}����Ɏ3�}�XmĮ�y�Qg*S��bu��H}�'�^P�t�aXw)5��u6�Y��~�^$��H)���I�l�T<��CƤp*<>R7W�8���'��\�/�����%@�;���uRW�g���T���9�P�A՚a���q�@�We�?[8�Y�Y1:����n��x�O̟�u�B��
���ړ�)������^�}l~�g�l����OS:�&�(��M��m$��*l�rqP�=a���3l��3H{>�I4�a�w�C�bAݛ��"�0�4[?%C�J�:��n�H(~I]]������NӺ_u�y�{�@�N!Y���I湄+����xè��}��=d�]��C�m4�P�?a�=|a�哜�L6�Si�~�<H,��g�RbAM3G�,0�� ���i��&���Q������JŜOt�@�*N�Y��;�6�Xo���6��|�����,�q�߰?0��^��w!�Y�%I��`i�'���'��6���L����@��
� ��0xӉ�H��#�#��ay]��56rzM ��5���O4k���c7n��t�!PX�N�H1-7w�\�������᳽N�`��j�޵�F�Jgu�����ڛZ��4o�!��$@:�Z�gWX�����70D��ٻ��ur��}�%�����������9��S��Af��9E�M�E!��<d��T�j���L`��@�*��ލ����d���kD�)+��,� �γ��}�����$=�z�W�?k������Ӄ��]_{� t{� ��k���1Ϭ]yHV��n�ɾ�I7��&��w(��*~@�N>��4�R_�.*�a���{�L�:�3���rm��gY����߾�7�1��NO��껣uF��귏~��h��
Ν�C��>I]'��`x���CF馻@ğ��Ϩ�o]����L�#�������.��)>B��6wXg_q��5�gsZnr;�/?�zE���c'g��H,�����������ڇ��?'��k!����1>g�{��J���~�iE��,1?v��>�xH<�ɠ�0��L}��Ue۳�
;�T���=���C4�P��������ϳ&�x�r�����i
�l9���%M$|�w�|I�*,�N�E>d���s5��Lg��8����S�=1�{�㾪��&��m�����N"���}����Y�>�9�T��ɴ��ͤ�.�S��8�s��i'�Ľ��HV'߻�o̟�M0<�sL�%|d�QO%�)�#�-IZUv�onL��_!�DG� p%�d�4ê�g|�oxAf��͚�CH����OP������a��l+�d�&��%z��<��E�|��\@Ĝg�w+>d�	��ú�hf�^՛��3��Wl�g�4�P�%g̕����=B�P4kXJθÌ/)��m��0޻�����y/0�!QH}�a���ug!��&�d�Y�m��� P&���*��Vz^M:X ���>��d�������P1��P�(��X�a�r鬕q���"��'S������Y<��Mr��<a�։�u1 ����;G�����݉�_��r�^����� 6O`��w�H=�x�滨}����g��Ci�~T��'{��H)QC��a�1 ��,�jÌ*��I��3̠�(�Y7��q�۪B��~���&>�h�gJ�f�=��ү*��+f��`�[��Oo��Z\���J��$��p⬌^H+.i�*���|�˫�u��f�L���Ok�cJg!�cx���p�^���W��D���'j)���c�9��o�Q ���یj�9;��SO4�m���=�sڪI�杯��R<& �*�<W�M�d���4�d��;���u�
q����qY�<I{a��!��
�a��p�Af٤3g2,1���h��~C�bM�nì1q϶z��I���w�?( d	�LG�|Ɉ
(vy�&��1&��߲m�d�����XV�a�r��p3+}ܚUI�8��y�I6�a�s���6�&3�Y�Ă�&���Jjf	6��:�����}�P�&@2��a�1��c�v~�V,��z�H%I��sAY�,���{�i��T�h�;̇�m ��y;��Z�VM��&ߙ*,�O�6����P*\!N��d�n��:rZ߹f���?!����Y�R��~����bCsY�Ԟ��Ĩ��Y1<d�7�g��~~�G�;�@�*�d�c8�+������S���woXz�07�q;�{�Xszw�.���y��6���6½��I�6��f���M�(�a��.��'�n{�+'�ܐ��Y�>�y�i��v�Y+�M�wz���7��4N+*I~�﬚a�B���>̶g����]�z���d
���$��a�>aQH.�y�gx���C������4����z�a���S�L@QM���O1O�c:ɼ�I�4���a��~��ϣޘ��U�Ǔ�ʖ�^4��{"" x�T�:�!��3�u����!Xm�L뼇��Af�;�P�<C�*)?���3�|��w��~�V.�M0��P�����ɉ6j��0���=�Q�۬������{ߵͤ� �������s(i4�ϐ�{�4�����|��
���~�3}�+.~�>�'��b�k3�8�IQ��'̘�7h�!S�:G�wr��z;���N�_\n�D9�� ~t��������$�)>O-&<a�1�Ϭ���N�È}n m*C�N�{�&�S��~�ω�
���ɴ�'�v����>a_̅�1P�h&qU|7�y�}��ǽ.!��QH)�MQ~VT>I~��a�B��Xq4�Y��wl�
�~}�M��1>Chc��d~��E<������x{ܛx�Ɉ��^�[:w���ֶ���6��.^�c-%,��]���{��t��PɗyTd�)��0���B��ޫB��	��m%�-;��6����cgh�R�'�{Ժ+�g���:;cGQ+u�޼��d�W
�e1݂�3�nc�nX.���ս��������������roS}��=0�P?���6�Y5��~-�0��f!�UR8ɣ��T�B��dRc:�5̆�HV�>��u�LH/��0�i�����$�x��bM���.j����o�������ts�L���c@�W���|���VLC����,6¦r���i'��h�z��T٪E1�%E�M�XiE��S;�N T�Ce�Z��^R�w��W�v�)��Y�_��|6<��@��4q'�$�^��$���>���T��{���a�<�é��J��˦�TR
d�E&>����Re��N�É�7f�*T����M�?�>`�}pӞϼ�ޘ B(��x�~@�:s�P�z��;@�s�m�XW���Mzyp��2Wi�]�}���!�w�~VT1�s���1P�a�Ă�NQCL���괹Ea�^��L������|�Y��C�i�A�0���d��@Ĩk��x�d�O/�QC���y扈Vu������aY�y5��F�:�w�iUIP��4up=��齹u[_U�	�1n�|>��R�=h��zΦ l�1�a��=B���a�����!���&ϿoQg����Ͼͤ���d��{����
���;܇�1
ɮw&���{b����9�>=�º���E<�X>����:�̕vy�$���h�i8�Rm6}GVO̼�+�P����c?�c?$�ğ�SH)���sl�T�����'��������p ��"=D����r3vn�=o^�~ϼ�߽�%|d��;���q���hbx� זzɭXxs�@�VOX�:�P��0���N Vl՟��~d띰��0�¾�o��h� ��Aiſ}�
�����Vn,��� >�5������ɱ'�ʇ�Ӿ�o�B��Y��sl��
�M3�4�TP��M&��M!���'���!�Uu�@�*h��L}N�c��C�J��3I?!Y�N��<��~�}����آ0�i��xLx8������FI�3��`mUI����O�'����}�0�)
�yvΦ�~g��>�`Vx���4�vw�i ��1��E6�$�?L�b�'c#���~~�
(�c+d�^]��N��<�(IF�$՛M���b��}��4>`9��I�ޙw�7zV�U ~��ku;�Qd��7ǻ.��*3��P�Z{X�2�fԌ�f�_c�x��I_6I�F��[���Mz��-���T���[�o+���{�y�;34��L����B�ײַ���
,4¦��4�|�a�~�k�Y8�����mįY*>w�N2mE�y;�������A�,�2���0��9��N&:==^c��* �
Y��2{j��غϻ��OQH)�:r�����^P4����bi'ɈJξ��	���M�fE:�J���7���'uO�;��6��+�!���J��đ{��5�^_�n������{������'4�t��&�u�q���H,�������QH- `��ʇ���HV|�1�a����4��1�aQO�ـ)�u�'��Dp<#'��v���=�^
;�k����_�����x�6 z��oz$������E�+�����q
�a��:�V0��TXz���oY&�T��`i>@�1����	r<&;��#�����h��f�����y�����}�4�Xm13��(����n��b�~��{��x�a�<�u6�����3&�XVk�q
�d���q�{���6��&�Z�g*���{�k�{���6�Ճ�|�=���t�Ǿ��@s�q�t�N����;��'��w<H,�N����z���&�w!���+&��&�@�1��C��@�TJ��U&?2TXV:�J�x�/�_�/sʶ�ձ���@���(��xdx�J���Y�J�{�H�>q6���'�T���n��r�|¿3����x�Y�{�L�e'��'(��6r�L�!P�_������{��������~~�U3��;Y���ΰ���S�O&�`|���^�4�8 l��!�J�:ɟw �P�J���]�*O���3�?o�!X|���f�~G)�ϝ�8��4W��=��k��W����y��2TU��C�&j{�t�����0��1����tea��4y��H)����Hu:�$<�����Y���P3�L�N-_�6�e��N���*��Dfɇ���2Zf�|�O�ceA��!`5o�
���#���q��D���w�+�.ry{|Cqb�k���c9�We�dr�������w��a�]SV�oĳӈ��$G.�����AWiU��&�*�^�e˩IV�j�=QK��ƞZ�/x���:�z��o��;�8^r�y����[v�H�5F��jV)��wu~����7��'�ݙ��σ�$��,C�5栃G�A�,p"�g�b]_����t�kw�F��M��(��ԋ�S��EF�4+){���O�<��V�!�f�v�_�ѥ)�T��^E��r|���3M(9�P�ʶ IUF�e��^ ���7��dɩC���5w�X�{�ί-���&ǫ�t26*�vU';���H��pӡ��zerk�Sz}�̧���+�U�=$��R�c(`tCKڇ|���M&ЇU!�S�]�ٱ�Y\Ŋ/8]�.�u;7��i��#��xV�V3Q�x��VD����$�p�gK��#��g^s�w���!�qڰ-�l�*h3ci�b}F#��5���5�RD��\�5%��g��r�UҬkZ����s����ݨ�65��A_-hAx�>��ᶟ6��N�u6�A�����!."
�1�����#܆�5,pڷ���{�,�M306�W��CG��	�:.�oE�A���JbT$%����g���t�#O=��F,ĺ��}��U{V	}+����u~4-�V^�J.�R�1&ô�=�vemLe��¤�vm6���خ����p �U��D3�u<��zJ��;�Vɍ��5d]�r�������X���2�ISz^B��3�a6��mn��(+?{��� ��θvn7��zn����9�J�x��mc�b����z���	��D��Op��\�Oӓ/���Bf&�����
��!�å4��:�r�O��0��=k�Ffɫ5�fK)jW��m�F:��>��9Fq�K����p_�ǝ44���H!�9
+mKR�e٧o0�Lh�pi�d+���n0K'Su�C�4 �5����MY��'2b����z���(�`wiqb8GW���	�P���u�$��#�z+�Q�]5�1�L�l7Εd�uW
)�;E��^_*z���D-���98Wj!#�f��#��m�ɗ��>�+�J��V*r]��c%ũ7h�s��!���#��^��^2�Ř��֒~�g���k�\kB�X�^!�F����w.��2�;��e�V+{�_=�,��7��\�9������1D|������>ڍ����`v	ϰ��8�C�^js0J�є#��R
���<�#y:�^ȧ^����*�.��C�k�k����W�웑fۃ{�A���)��G�[ۘ��K�{�˝O���t�i]]Ǫ���쭋[�j'��ywu�YRR���V���l�e����ΐ��}9v�3t��'���Ee��=�/�h�&5u�;V���
G_RS��7{�xvT��s�6r�G�v��1�R��� ��/:�7W�]���:��.#�0^7����U��79�;�%��]�\�lד�v��ޕ����q_ѽ���Z��/��S�W%�}�4��d�'�LP��lэE:�74��uZt�M\(��W��֡c%l�����+ݮ�d�Ԓ����cj�$��>�8�B(H�"�P�<gTې��P��qX�ܭb��w.�ɐ�ۇگ�V5��Y>bD;a�E
��nE�2�t}s�==�e]�mU�X�(>�[2����T�*%\R��=���U�.(C��c)����դ���g[s��%7]Sa:�
���*o7,*����$T�:Y��	���*��v�1�î� ��+T�	�h!A"�_��d`��N$F��M��ss��3W�'W/^�bf��7CJ�t���Eh}+:�v��uH@g�����;飒��ƮeS]'��M`:WySU�Ѵ뺃��E���.1�z
�͙��x7�B/�V^��V���04���X1%�l�2�Q����;RwΑ>ݶꯌ���q�K�:�[���[ᑝ�|������Wr�P�����g�$�94:��ɵ�B�v��}��Tk*�2�9�^�Пq��JSj$���2�0s���}D��+{���.��>�2��s��r�.qaW�9ۂ2\�,裇Sa�@�TZ|Q� Ԩ�"靮���:BoB�\�bq�Y�\��3����j�7-ڽ�t���\�2�w�H��$��ʺ
B�>�ܖ!�\ʙ�e�O7�k	g�q�A�ۓ8�c9�X�eJd��ї�'�C]��u�)A@��x��]Z�ۋ3��p't;�ms�dU�Q�R�؛�ٔ��ĸ�6�4���K.�YI%JJ�t,P�
)x�����.�z�Bw�9芠Z3z ��o:}��3�z`۸�En]V5R��(��8����ub�7�s��[l�H�Pb�	�m�]�]c.�ǻ��*�:�9�ّ"{w�84�z�	�Qg#j�DIS3���]��B�Wz�	֯m�s���l���,��(��,ܲ�	G�Uӫ�J�%����\�ő��&������K��;��U�	�O%��+ECժ�m�X�FxF�����
�ٽe�+�=vReH��/ht9�2��t�XB��Ӿvr�Y�l�r"�|��B�W�����҇+{}6���!b��Y}��Z������LV����WDh�YV.��Tl"�s4��[�69R� �S���&K�`��C�0;�cx֒��LԍBfLu=L��*�ʼ����onޕ�>�\�7�i��`�5�]�ަ})���Ut\��A:U�#l�A)\ܡ.�D�yZ�!X�Wl���h�u�ͳP[ ��q���	�{�L��gK|�W�b����ԫ�,X9�o_t�Z��0��ƻ��w
TUI[�)��.l��y�t^)��!����ؠ�o�X���Z�]�����>b���<��C���5���k��Xܴ�_\��v�sK�5I;�
�t�μ��7qe���%��.v�g܂�s�nw�v��
��nl{O1��NRP�ҋ��NW���[j��gb�YF�U��X�c)�l�x�N�\��Mn�ur��mR���V�R�ϋ96�l��и��k�_	�9��Y�b��)�	F�X4쮹�U��M$f��ڴZ�a�� ���x/�Ӄ�7�r.�\#��/yX��3_�!:�Fn GK;��P�m���,�"��i�z`������n��6��&�s�{ƺ�hf�Ax�`���a֡C��f�h����-K2Θ��	b��s}�f��.�f�J��Y�ke�y�<�!,<�V�F�E�Z����9e�N�����gZ{u��֪8B�F���������k߷u���R�F*(�Dr�`ۘX0PPDEE�"�Q���B��E��"�$T��QUQ�D���#UQ�����0��TU�(�ZTX(���ődTTrыE��1�������1q�`����X���*",QUTFF(��dTlUTF*��,��V*1`1����X��T`�,QU�m�2�"��"
[kUC-#"�b��Db*�`��*E��ʨ��TX�"�UT��h
�#EF�A�(���E�UEX���(�1E`ʅb�"�8��TTX�"����*(�1Ī�e�b!����EYF*��Am�QF""ZQD()iV���1b���V/��ͣ��W\W�Z�c��2l��wsu.S�>�tOe��י�H�3������<�E���9\hvj�º�+����x��\��o��t��*.Ezk�('�d("�:���#2�5�|k���O��!�e�O��ϞdӃ��C�z�����Y�Q��^�mJK�;w�۳�����Ig5ӈ���p�|����i��<�<)��J��}�e�hՇޢej�m3��Z��p�|V+V^��~��j�i�V`S�z�����w,���+@]G)A��j�iV<�ŝ�_�V<�R��,�]� ��F������e^ņ�^��*�q ����ˮ�"�I$�m+�ࡱ�jp�W�N��b��
t����e�M��wKo��B=���s���=R��Q&�#�Tl��'(!�B�\�S�K�t�r�ǔ:F�"�m�ۂ�wi��Q�q����j$���hh�ƨ	��%G2����i��@�S�w's*�٫ǀ�~l�s~t�E5��QҠ��OD��)�Ah^qƣ���]���H�}����+�s�W��a�Q�L&�����b��E0���˳;!ڇ�Q� v�Է�����7+�;��z��sQ�}B7Nb�ӥ�¨j��ؿ�w��n/hl��=��-vsǇ�����^�\{9o.:1�V�!I7!.
g9Z���t:�c�e'�e�No7�f�6f3.�bڑ��WpY��u� {�ދa�b�'$���O;$=��*:9ɻg���p<@�-R�"$J�<������k�������T1i��y3�������[�t]_�N:�*痔�2rI���Ă�{��(W��
bgk��.��b����r�)��x>���}5���1���=���w>�|pt>R���w�
�(���O]���[�8%ﬁ�1!T���I{�L��ƃ�ad�N�n�	L��,D�*�p*{!F
��U���w��g��>*H�3��Zj*�탪����S��QPS@�����G�kL9�im^��ʠ�b,�yWGG['�.�\f��Л�[ �5e��^y#}4l7c&]JWn)"��ѹX�?_���v��@��2]���[��:�����p�&GA��$��0��D��:vn�����.���yI�TL�Z6���(C��A�w���$M��<f��t���GGF>��4|��IU��*����F�s�����p�I��F�����B�umĝ.{$�G'vR!�(`ɹǣh�	).6z75���c���}ƛ�u�C����of{+h�Gta��W�JIJV���խܝp01��oG3ڍ0��*�d��bWHGbC3�Gήw�(��Z������y�\�=(rjw��\|U�Br�gX������*b��Nm&���٣�7�F��%�{���Z��$S�cX"�eǹ�t�V#zB�wzk�_� ���=�U��N�qf&�[��������r�r�.$�T/�������o����\9���n�0�ck��1BP��h��	�_;P��t>�	�P��'��g!o��o��m����J��qF|p�P�q�]md[�܅��/ڏ��,�|+��Q���5g�s�HOx��P�ɪ9\x*�U�U$<xt�ɦȻ�] �:�e�ɨ��/	��螄d�Cc��mºgr}a�q*��\
�p������K\'y�F	Td�F_Q�	���V�C�n�]s�������d���ϠR�r&����YF'�v��;�z�m��ְ�T�z�u�UL)�P!�ì$5�#��t+q�nJҮд���>E魟%�C��&'��5�Ϯ�PĖ�b�:�¿B�sHxm,�TN�����Ma6�x��/x�{��]���=��[�b�t�9�݀Օ����k[kM>wR�c�HΖ�{ڻ����%�]^�mc�t;}cߔiq}\��7q�6�=K����	�^�sX�/���2;r�j��;�f���HJ�7���xxz�j{Ԛ�x�O��N����>"��Vl��g�p���:q1v�&`l����o�'��_l�����U5x�9Pf/�׹W�"��_�ܴ�j�bf�#��r�����ީ��Y-�=�a�И��І�q�C��b��	�}}R7���5]s��,�r���%���P)+���7g�AG+��_ڄ?]�+])�B�N�@�^��e]����}�׃���$���|\[�
t��^���_Mv}�(j���Dq���g�¦�"��QP��A�%�Y��w��c�v��aL\fH2輺:�;�	�3��%k��oڗ,��aޭi��?����x_U�OB��
/X�#��B+j������=���7��x��֩^KAuԾ�~��R�X���-� �QS�pj�r)�%
�+*v.�������l���z
�<���*|���t����
���,��6R2���Bq�_O$6��r�����!��C��k��T
���l��j¬�����nu��Ok!�Me�L��Od���chg9P`!�Ӌ��b��X2���t���v��ur���K�|�M�wuN&�B�2�s����MO�ei�̃���G*��_m]`���Y��Q균��:L�N�����a��:㛞���F�F��c��E�Jn)��<���]�T����	\����������A��g2T��ܶ)V0j O��Ǐ��T�+\��õFE1O���;h���v�5��cb���u���/7�8h~!��W�@�~�%�b�q�fu�2���p'^�s��M�^f���"+���´-��U捧�wP{lTO�q�����O""��o1�Ve���˺ᒄ	�������Qg\�L9Wk�OJ�KEo��g���^N����{z[�7d�p)�p�3m��U��$?�.!�6�����x�״|tX6ڌ�*R�hfûλ�(ko����C����/�X�=Y��٣~j�I�{�0,�0��+�l�NO/=Em���N6P�V�N�̧ł5w�9��-�(h�Pu�U	z/���*��H���o�*�Z��.}W5[J-�'�����PS���8��|�̫�o���զJw�}�zl�ܕ>��3X�=���P_y�c�֗r��FY\F}�80�����VQA�2�kyQ�
m]�����hm�_R��J��D�l�%�S���� X��9!�ܫz]e�ܠ���u�9wtN7���-�S��j�G��mG������ҧ*	m��ba���.+O�G`8"��5���V.HɎ[����X�to<���<<���lA����w{j�d�4�jy�D��"���j��:�s��<|+6,�B�3�{B���p�}"�W`�u�a�uJ-�$<U��Ъ����A�j@P���X�=�ۈ�Z�L��=�v̜��{�9x x�2:����t�E<R}
b��p��W��^�R-��� Y�zғ	��q�=�E��c���ϥ^?�7*6=�>�0|�;�y�
���]�-��c3�j����O��3�����ؕ�ضz:�����rB����W��Wbv঒�́"%��3R&(w��@;�<9sp<=��������]|�1�sU�1�KI�z��`Cָ���B��;;A�����^���ܽz��K��Exl�Q\���ʎ1����GP�%����L�U��x�<'��]4<W�|�U��'���0Nݦ��j�=��(�5ԙ}���N����X����Dp*@�QB�<�����v㹚א&�+wu�W���3��<9r,s���l��>M�o��aCG��4�{��+�����H�`�2����[��Rf��#�Mky}�3����Z�Cm8)滬<�\�tE_-���F+BY�b�79���UҖ/LSٴ(���Ҵ(����Hu�Q:����-=�;���t�|��\��l�Rψ)�u�!}�ښ��x{�%�׹��7�C�	�'�
Mv%�^1>��o,O����Lwi�5��{��x[=:s{L:U�MN@*�d8��|{	n{�T0�s(�~L��{�z"TB���3q���A�,f�٨6G&O���(���!F
�2D7=]�8�!�y"��9B5(V�񒛜���Vȝ���j\�^�XJ~����Pc�A�K�Hخu
��Uł���po�*,�:����y���ϋ��NC��25�z)c��P5r�N�m&Y�խ��m�a�z����q��P�$R�z���ۏ9ӊT�@��ݨ�"�W��l�
$�Td,��1�׏l��4aZ\LZ���PN^��+=."
�};�w�,#�B��"���!,�ʎ]�\;�y�H3/�2�(N��>�E��/����GA�
>}6�X��v�Q�:����wg5.�ު~ޥR,{ӱƩ�J�ɪ\�Vqϫq_�1k���~��.�Z]��n�k��Uʎ��>��ЛR����UT+���6EߡW@N�������o�����xN̾�d�<T�jےz�$5iWN�8쎝�ʂ��C{���95r��Ƨ�hB��`�r��6�m՞�
��S5�.�q��@�A�ڔs����I�r��ugU�M�ڒ�h�6�ґ�.MR73�E��#�6�޾��_W�W�_@�.=�j@��W��]S=
]eϐl���.P!
Q5� (�G�� �tػu�8����E����(����"����^��!g�!\ߩ�[���~l�yT9A*�S#��B�je�\�Ԑ�\��x�証T�p�*�UL6��%�nC�'�A�F�Zq-[=K��ɽ�����_�tJ{���1�.�_��� �E׼�[��S�;�y��Tߵ,��`�{�aM+�|�h��*o�����G#!�R;v�78�p�V�1��֝8i����ba��P��L��4��Y���JFx�£����;���q�R+p�s�K`ִ͈�����W]������V�q�j6\+kmV g`��8Zk���k�)�bu���XF�q�;��q�-����e^l�$/E`�r�tel������N0���ɂz�r^�yR����ѪSO�*�*-�AN��`cu}5��@�]���Ӑ4�=Ǎaj.q���y	*fƼ�=B���%�X6k��.-�v���8˝�᧥��5�xT�ި�A�NѺ]-:��k6�R4]��EL&��gi�yCI�r�찄4���W�Omf��Ǳ�X(m���T�pÊ��A�|7R8����y�.M�ӊt�iW�����J�\�l�o���k;w�u�=�����x�ɮ3}5��S'�:СX�0�S�2�%63�ӧ�j�(�'�!gG\��Os+x}��]��`"^��3J�*��B}��>�8�i�H��J�QS�w"�V��0.60�ٜ�J�!��
����q�>��>�k��?��G�&j&��Z��+����״�Yuz��w�;��o���q�*x�S��]
�,���,��tu=�Hg��M��1�����+NL���t5M�'Y^�V��o+���-��Ƚ��	It�T!�S�T�+��ʂ=�+\��õO�!A"�_���"J��p�azDI��������@���&4<!��+����ʉ����t��ڮa�� �qi!p�4I�2P���ˣ
q�C�F�8Jm-���DE���I�۩�M��~�ܹ�j�ށ�e�с�������]�j�z�����/��ipo�c�O�<m�����99#�5?sCό�������uN��0%À�xE���^�[�h��qM�l;w˜���Wb�_����<�Oq5�r=��q��
�L��L�P:ġL�g�4������+�jݼ(�ٮ\Ǹ�:�6�ݙ��ú�\��flMN���Q�R�mǨ�SWP�}��i�2`�Сў�O����8.Z Ͱ����Sj8�Z?{���:�n��s��wm���Ϗn��>u�� �}"��=Y��٣`>4����G樽qn�}яV
��`��>�.6/:б���@Gۇ"�y*�A�w�:#��j����b&޵�#XO���t~\U+Z'���A?y���S�9��Q�U�^�j��<�Ӱ���Yǩ���qM)3����

+�2����
��N�BW�
t�i�x�s�s��1�{�ٲ��̨��%kR�mB�#���l@h��<T�
�<�9�t�b3;��n�+�ii�Y�E�	�p�R�r�E����,WGA6�kJ�u�1��q+���g�l`���m[�gU�^x* ��;S#�6E��霊x��(*��81�ƽ�[�A�P�%�#���1Tx����m�ϥ^����q��&��sO�f�oz�����f�C�L1ޝ�Be�`�x�*,�,0��v��
;ʽ�;;oÐ���ڼ��n�w.��!�:��(J�ӪML9PEH����E؇AA�h���U�1��1��A�Ʋ�mmؓ���P�|MĭE<�u6�2�����bÎ�bܬ�:u�*�h�{�zg0fj��Zew9�c܀���U��j�W,jJp3�'"U�P�d$�>�݈Mt�H�Ј����y�5�k��i1M���K�2֍6н�˫��*ﶺ�&�'m�<sU]t�c��t�0�OQ��.^�ox������0.\i��\h7���5M{�NnPT-*1U!մ9�_�3'kW�{����`΁g3��N0��o7�*;{;yϜ�ަU#�r���P>�9ػ8�qj�3��b�$�V:�R�;Y]�����Ŋ�]d[�>E��ʌ���v5'�Kv��#�KE����۴h!��`YV��� f�̻^2��.�cWq�1r��\��q��+�e1ڰ�OKUi�w�_bҪя������l\)�w��(N��{d���8���<�Q��mvѣ��TT��ק�Z��	Fs��
�"ZƓ�/\����H���}uЅc�5�a2��KY֨.�lp뮙��	��;'&3:�l������]����f��)WW 0`���-.�r���i�څ8�q�Y�6Vf�V�Sf��#�&ބv�>� m�m�������,��{2U�S;�=���ن��n fAu����+���x�a$����q��銶�4���9͢�����02��v����LZ��}�z���Er�< ���WbF���4�Gm�i,�\����V�u����Z��{S�F�'	���KU%�uj�;<��
�sS?]�G�3�7��Ч���w}JL��,�<�oX�Fg=Q.��ө5 �Ĺ4��{�[�_K"��9��2�rS'�Uƛ�v��X��H�>�hR�b/�T-][�qwn]�\���+J��w}�wFQUq2����z^*q�.�뼬鋪�>�� �kD��Z���I���}�#wb��G�K�;�k�vM��peU�jֳ	jht���{�l�n�g*��<�����p8_*ԙ�,Z=�;}��+�1��l:�eM�tQ��]�e��c�(9��d��3�\C/w�dWw+5j���v���b�ה*fs'��%��-�U|�H���@������Snonm=�ò��XL��e�r�0x�u�����ڲg��Y(N9V��;X.���fQAR.��l� �|�ՏרW�{�-C8I9�,�Aè3�+��%=ʵ�:�[VB�8��bHӺԻw��@���Bh<y�å֭.0-�j�V��ѵ���b�%��E/m�N�t[wJ�c�S{k`Uˡڰwv���ZF4�6G=OTb�_s�
S�(<��}���hv�����^Q��z�논,� ��Ÿ��r뼙��/Hc9��L�!�姹EB���+Uu�<�]�
�N!���]d;�^�*޶��%��u-[߇F����Ɨ���9�}��g�k������޼��E��E+�����F*�Q�eF(�#0A�,X3�b����DQEQb1Da�T`�j�V"�(*1�B�"
EUAV
�F1[J�b�U�,E�ł��(���b
"(��1Q1����QQUA��*����ԫE"��DFEEQTU-�"���""
!�*��cE�0elEEUQEAQA�AA�**�����*+%��������Z,b��T**�*��0E`�X ����*�Lq��#T�1"�EX� ��F�(���"���
(��U��`���D"ŭB,X��DQ�DQ����w?f���g����W���f-���.\����+K�ό{r���a�	{u��l�<��-��Xl��j�.���x-�);��ڎ��+z�77�E������$a��G1|�^�ː�t���n�{,��s�_��(�����p�\\�pT�L�Ty�Q*8Q㐰P�]�S�a��-W79:)�X|,k�2�<���b6�,D�*�R�2�X�u=��t���㸉]���#QN�W:�Tngb�pr6�X�`0|�Y�:
�]ʭ<Z~i_�����}݇e:���o����X(8��dP��bP�E��c�Gxت�ԇUu̘"��D�2�!�gw\G�os���ܯ��'c&K��8� ��X�����%���P0Û�n���]E�p����9h��6��Y̡�&ޜ٨6�ɒ8]:��g�p�������o�xzb�8WtԺ\(T��9���
ϩ@=`��>�wm:lv��:�*��1��"c .�om��/&V)�l�lDr��.^ϋ��NAu�ca�[�O��Ơ�A8�sEq�/DW��E0�3!FÚeB�J]�ZL��9�W���wzAfp(�+�>̖7��kD���l�ǡn=�c�k&��{����<��F�s�u��4��l�m�F��
�W��|0e��r�֎�([����;�������l�|������$��7P������Y�G-B�z�(%p�-Vr�v_Y��Ꭷ.��&�~�����MF�u�1֨("��r��5nVK����A�7�D��9ok4z�����C,��w�5�x�"�DI��Z�#�ߊ>}6b�.�6��ܤeU�ow�A��`v�V�8��p6��;2�%���U�x����[a	������H_ ޞ��ݐ�����ql�ʱ.:��F�M�J����r�Y��-�.�]ҕ5�M���^��]���覗<Y��J#�|�P�AT@QQ�r���36�.J��ō���R���JE�p�p/Us���̾��U����
T9>���Ƿ]��˖�{{�Ѡ�\��t�T�\\p�*�UL6� �-p�`��\����v���&;���wt������]�T�!�U�@n}��ڛ��^K��DSC������g��ޢ�}��_�k���S��h�xҿ��
_���UԜ�2#2j�.ژ&�v�ѕ-.�v�OU���(���ʀ[�dΆ������X�7��tp}tw�z�7p ���]>+s�j��9r�L�٨��h�J���[��%�%Y5n�*(���V��`��i�H*����z@��.���\��ޣ� �X�:����wV�ء�حe,���O~����C/����aٹ)��)�U�M�}�}iKo�%;���%�\��~1��Z�{7� �Q�{�LQh�(�N�l��8�k�Wذ7���*<����[�!q��X�s�Av��<Ce^l�r=�:u�Wџ ���6�]�o�W�f�W�z�6=�<�5[���R���Z��nV�E��)�>��{��bo_S�pL�z5���y�����҂4I�"�T7`��
�Q豔K��lד�v�������{�A���s�����%�R����@ܡX�0�u�q)N�:�:z��P%������/5�]���.��X+e�����VWD�+�^�`�A�"ҡ8-�&lF�v��B^�����wM�~�R9�P���2�]��v����^��ʀQ�%�U�m��Ow���Z����\md�>*�e�	�Py�̨��u<=���BTNP6z*{x�#TA;!q��i��1U�S���U�����s�!)��CTߓ�uƟ�X{6��x��bw."ʂ��kaDyߦ�ML-�f������Gh�rӧ��O����s����9��'THIX�9=��Ѽ��C�v�u��dxCŚ�3s���a�
. �����:�Mw��C�d�gɽ��to[�� ��+��>����f�pc� 降�-��Δ�`�z���y8�������l��.��4UfלX��I,\������-{�V�U��7����'�iW��(Q�]�c�t`j��s�RC�|�
E�>]��7@� �'W��)�{��
��)�Ζڧ�Lr��fy	��z�蟙&u>7 �t-����R�Yw ������,�3�,B9@�Ƹ�&�t�j�Lk�np5����h�t�;���D��چ+i`�,��u�e���N�� �C9����6����C�ga�l��`F���~{Gf���d�WxT��.��vU����	�R2
�NC>�*6/:б���>�9Ӄ�*,5n������jCn��z��ɻ���=9T%�EV�?-4+)Ŭ'����8J
{�pj>i�6�^��L�k;��a뇛���qMEg������C�iw+�tg�����%�j�]pɣVT������r�Qp�G\�o�$z�g�l"8�FϫӔ�!�B���������(�<h�FZڵ.@�)xkZ��8V*1�y�,���B�x=:i�h{�nb���N��o���ÙԷw&Z7O�#��J���kbOE'�̻k�z�*�j��(Jөͩw���V]rc9c�x�r�)_$$Wǘ�=���{��F=��La��N��
f_\��Ѧ�N�z��_>8�&���whvwb������A�ﾛ���T�ޮ��:�
��fq��/<��c�2:�"�ۦr)�G�c�NT�õ�L���
v	aʳF8�����̨����^�>�x����S��>��&6���U$�6���٫�\���5�)����
e�J� �>| ����{K�7�ʞz7Hl�8\�5צ��{�Z�!1�H"��5�ϖEA�����W��x�{�u���|s~ॾ�d��8�y��RA�=K�X���̣R��kh�*��� ;K��ӵ�킳��ͮ�����T���S �ߵ�8��'~0�q������y���(��a���c��WC(�:3��I۸������Eμ�X���j^�f)��b6�qb%��U|
�8z��Y��e����C��:�x�������Φ͕&��6�ٮ��[]���:ۭ[���>�b�7t��,w�7��9@��x=�P��`F�V�r�K��o:�7#�w��S�`�?{Ɛ���b�^ՊYC!�گg��-�oP0Ø;�nr'#օ��`{ww	���ڀd��m�X���[�ti�����q����:a^��ޕ(EBR�)��M��8�B�����@�r�[�|`7�Q=w�:	�ۄ����]���KG��G�!�C��1�x{J-���y���<����xZ��OUM�߼�>��M�9�Q^*ҡ��f�&�p5t��ܴ�n��56�8xe�$�;D\0����Nw��6,7�ttg�Pٚ!�ؒ��;F��/��ǚس�{(��R��3��D�!���.^ ��n�r;��u����K_��T�t.*��SS����</g�����y�!�p�����\V�����U�q�!j�>j�u�3���p�Z�N�L1�k�="s��F>r��^�!��9t��K�5_i��3�Ĵ�������
m����W����Cx��A�XG�ag�����Gϧ	�\2{��w�,���v�`�	�]3�=�V�R/�6��c_�u�M��k��SלC�{��഍�+R�7�3��G���ٕr�aA�;�Teq�U`��CǇF�Ժ�e;ۘ�֮��λ���#X��*���PS;�3�>��ʛR��*���
uO��Ͳ����K<n�3�S��)��ذ���\8��\�,��e��%��*�l�%̪}ڮ䩢��41f�R���=2R�~�Y����΁�3vY�R�����
�{�mW&�s��5=h��}Vi�:x�Lŉ{|��,.�s�L��es�P|ނq�X�^y�����n�{��$�{κԥ��'5.��i��[puq�꯬��g���,
Җ�&��ʣU��	R�� ��O����!��+ǹr<�������e,��f���B���|P��U5\���0����Sy��[
�E1<�V�ʅ�d�H�;��k�=v��҆'
����׍.�b���P��Nv%�	Ƽ�q=s4sn�Y��R���f�-�t�b��ʀm��!���:%�<+\�S�7�SnR�٧{&f"L�isU�0��\�lq�!����{.uч�Bb���e/u�a��3����}�o��__N�+5*`PmW��!ơ�X�bq�.û���e^l�r/dQ�ؖD�kl`�L�˙J^w�?z���],]%�5�]�$����E�q�+<���8 �Bq�F]���Hu�wZ]��W_M[��(T�X�%�"���Y
�;�D�6k�޻q�nq<��2���]+��ԙ�6�~<
�w���L��R��6�
�=SP�`����Sc:�:q��M����[\�]3�0�W���P�̕����mrZ�������]Bw*.�_��f�Sv��HSγ9vE�j�r�����,[ᅶҢk,.&��*\D�53/��q�%a�c����e�61:V1��8�#=,�8]rME��n��ev.w�fs��,$��׼��_C�.je�ηw5gn���-"$����C���g����y�v���/|�(V5�2�]�3�/"z%zB�r�Ḡ�!֎���#�ٳ}��Q�X�<�X��]�U^�8���fTv>6׾��<p�tt$��j̜0���a����45a�>�ޜ��E9��u��wyS�&�F9)���'�=�w\��W�����#yt���eG���T�+\��õO�!A�r.����Qh}\���5ћ�yB�K�\H��a8�G���c�_�o�x#M-֢��V4�RP����+fN��>J;�/�W���
z�A�� _�c&�l��/9����A4�S|&'ٵ���3��H��]`�ψ���x)[J�I�狯D�/5%��d6��k_�c��>K5�Xi�{����
\8���3~n�j��A�Z%�w�i�cŌ�Ռܻn��Hi@��<�'��mߍ;�vn���F���a��"�]��ڦ�+ꉒ�|�,l�^�ح�H# ��<�q��δ,vw;i�V`��.�<�[�z���ܶ3pv�rgYͰ����W]p�= R^L��{��'F�e޽��<�\��E�M��l�<���ΤJ|�N�_���K"aeu��(qWWF3eGW��.�T�������U���G$���fȖ�p��Y�"�2�Eǆ�vk�����ig?�U7�M���	=�6MG�<�s(�}JkՔ�����T�����8�p]1�]+��媬����j�;�8�����/�Ɔ!`�k�xV�3֟���Yy��y9�-^j]�Q{$U���*qΨvN�{�=R�>*$��"�6}!���(Y9a�uVa<��EF��Y�cU[�:E9W�`�I��:��R�U`�ޜ��h����6�u���qڗ�h���q$OB�_Z�gU�^yP��jdu�E��L�S��DL��|��􋞌���+G�O�[�N�S���y���Qn��������ɻ���<�Xz�N�wKr�����C�[��:)�Ѻz�������U�.9�1OO�N�KYj��ڱnʍ��ὬU�^����ϖEA��"�H�D]�tbyFeI�v�$�۶q�!�lfK�Aś㡚yy�lމ�g«�p3�c]$0��dq��{�Z{��E	�TRr���8�U�D>Z2�|��p�
�ŉd੶����S*��X�8�9�_�7�����t+i���䑋�*�3��t73+�4��gT�������k�>ה���²'^2�z.��q)�����=���7�3՚Y�R�l�����d�֭��_<���m�8ė���2f�2�o3T$cs����}_xx1�s�<���ͧB�g^G�wC��L�L�W&X��p��M5��.w��(՘Q�ә֮��0a��qU!��0����#3�`<���` ��QPk�������&^jcW�]���4�Q��<��)�Ү�bǽ����ӃۦЛ�[ 5E��U��g���;��:Y~��eU{���~�� 7�C�^�X䊜�U��C��G�����ê.b:ra��.�kt�v��/�u�>�;��d���2��D`���3w����cg�j���
0k��;�p�_f���#��Pٚ/Đ��;PU
��,=K/j��s3��u}!�����uĄ!)��.Zu�n�)
oH�K�b����p�m`���s�i�6�w�TxAN8�B�kH�4ῃ��B�)K�`�W��ǈ���5��ʭUt��wM���k�\ǀ�T�_ o������ҍ�s׵�˯�Oܥ���=�^�5fN�]��S�G�X�!���K �|��x�8
�����e��3�W8<�g�	�#!l]Fm�!|�B���ն�-�Wd�Z&���	�/v� ���g]��7�����.���k��}B�_c}�,��
��9Yǒ<�>�&�M��8jh�|�����j���n1M��h�5�c�S[DM��`s�yÖ�*̥b�;�I6_CQy8��C�G���^7�Q�;��I5p�����&�wbc���F�fWA��q0����w���(j�*7;*��8]Ջ	��P��[������ؕN��ۊ۱F��:���-�e�n�����\� E0�����8�՗n�A\D��_��cq��]���yud-ۢ���#�-�V5H�{&��P0���Dw�8��J��I
S�]G���WpҌ��;G���-�r��
�ȝ�����.�E,�Qгy��7)-F���z�����+K,��Dm�CB�+���Q\$�]��P�*)�L�����.�z�צ�\:�H�#��`�tϳ�嗱U>�_�]dR�O�-O�Ѻb47�y�>�ɯ��2�R5�)��VG-�dvrcn�4��Xb�:�����o�������ܭ+�x�ND�e��7�2���<�١�xU
Lб;�ٶ7)�:����{����Ǉ�s����_8��S�W�C��#��3v���8+��,(������sQـcμJZ����NS3�崪�GVh�Ytk�l�E��3�S�s�j�5��}Jr�{�@U�6J��z��y��i�����<ݬ��YL@m����(iQٔ���s�s�[�VO�Qݾ܋Ww`���_TSlB�YntƩЭ�NK����f�*2;��m�e+Co{(ի�74&����7A	l�On)�N�2�a1t�����f�TG�#t���]�a{x�5�Xn�7GU��k�R6���\�+�)��-"��x�1W�YՔ��|��*ҡ��9�ݎV���'�\r��v��,ozh�A�yr�*bO�>@��I��i8I���:r��DpϜ;���ʹ�J��C�d{R�h�'�Vl33������;*��h&�r��Li�"B���=��;�K��;�f#�ub��^�;Ԓ��`��]<4PzfY�ɂ��l��Ӆ.�v���2�*X��,>Cb��m;�z�����E�F�Hłe�)�ݵ�_>Ogt�8}9�ㆷ�����}{�m�/�Wׯʇg�ֹ���f�Į��Ԝ]P��˼��\��l],�#����hd�dp�U���U�b��2q��cY��_êg��}n�tc�����,ұ�l6�k������ԯ&T��M�*��Dڃ,C9��+Rr�ǘ���۬v���q^ՕX�ZVsP����k~��Ej���MA�[�f�e���{9n�i��K��J�aڔ����=�Nt�5��FJQU0�U�V͹S��O��I��� �X(��E�
ڰP��\�U��X���1EV#l�A��(

Ab�EH�R"
����PFE��Tb��DU��F
V��X�T"�T`�X)b�Z����AEP6,�iPIe*��`���R��f2UDQU��(*����["
�*&5��ıF*�"#
�d���������Q��`�"""�1PUt�DQQ`���b�(��,Q�2���1b"����DEDEE*�F1b1TQm�V�U�E��*��(�"*0TR�fIAUFQEU�"���rʫAQH��"�Ub� �U�畴�Z	�IO]�t������z�\�u��^V�ܽ��0�����'"z+9n�o��:�.ཙk����6{���1תʨ��wԧ���P�Z��8�eU��qu"�l	�N�T�%`�\ʟ_�x��A�[�9���{k}ӌ�b�R��E�w�N�ep�sPE�n�ڕ�p�e�u���U�"ԇ5F��W>��.�R��'e9B�(V��b�ܟ6ߚȸ�b�8P�"�F.������uK�7����h��M�O
=*m��U�B�B��S�,�Xb��`AR�y��)sK.��j��h��E
�'J���xˋ��U�U0\ߓ��Uj]=Ten͡Ro}E��,44z��VR�-�]����9�q���XeUa��cs7������fU�"t�ͤi��1'�ܮ��Ǽ�C2���6eu��js��욍R�\n����=����3����>�.	�V?��7^���I�����a��NE���˴�Dq�!�i�&^͇ �Q�p��!���kCpl��"��gWn��6r:W���� [>�|B��ňw8�n��6U�ˀrEI ��#�\��E]gA�T<k��ir���ն#gV|[�X#����-H􃳁9{����cw����]9쮷)�n���:��hL�{Km'�!v^�k�y���p7%7��X�Au݃�cH�	F�wF�N	��K����V�w|�Y���}Ul����N���C�+���l>G�`��m�+�=:��Q.lo=Y������q큛'f���D�#��%C�KB,i�
�¾�S�ȇ
+;�U�u�s��n,�Rݢ��"s��Wt��u�$@�T+��ф �N���%(�h��r r2�T^��/��5p_���8��,���	���T�z'P�mO�C��B�[��J�ڪ�	o*�_���>�E��U�E��_��2��E���L�KȞ���!�	ƅ۵��#Y�6��]V��.)Z�f��t
RvYL��ζeE�|r��*%DT.����sy�oe�W�Q,e@�qL(G%���45a�m��,�H�}N����d拨������P�]�4�9�>��T� >5����])�(��t �Toh�r�2��fl��_>5��^��:1���m�0Dڧ#Pt&����G�Uɏ(Qb��!��]��ڵ�݅]�� ���1�u�ˋ�� 3�tӫ�{B�1��T�E�x��{�i�kT��۱j@b=���^]Z��(��[����6���Ez[����K�؆���M���d�h};���%B�u���6�'�|�ֶ�Eof�:��ޮ�R���v�M���n���BzԷ`�W��fu�9�,X7��*wS�߽�:�P�r������"�Շ��9B=�ԋ��Z��A�Я��p�hvT*�3��D��K�M��`�9̟N]�
^��s�q�c=.��Y�n�iJ���B�A�vs�Ś.��w�+զ:\NNt��4�;3mߎ�!�ga�l��~�� V{;[w'���Y�Y��3<�Κ/����xT����o�o��P��M��Y� ���{�k�!�o<䞇xߛ<\�Yc-��U	uEV����V�'%���Z\�i��B1�hK��<�*ֺ; ����?2�b��+�Z��4�=2Dz��J�/�Z>�S}I8Zk���U6&��7�9���4G&6H-�&�@t��T;'c9#�+ |TI@���o�
��pQ��3HjԄ���i��Un\�S�z��y;�Tc��U`��zp>z�	~��@2E��,�o����$[@Ju�$J�
��[3�j��Rwa�#�&E�Q��̕7�{�S�ol���^p����l+kL��Q�T_~�j/�U��nEl�3�4fe��y�-WϣVu5b�*�@�`[���]KD$�[<��&�\y]3���˷�w��f���T]��� �gW|��]%�is�)f;�SM�� q�� ��2���_
�(��t�$�ݻ�A]ur�Sg��Y+��X����䎉Y�u>���X�L5?���__��0�'�P��T>>K4m�r�=�-Sxoю��.��w�v������(_��W�R��k�]�,m�ƚs��<ڴ���h����
	�	��^Gg�7�E�υWP�gR���}Ǜ��j��:��ҩ�l{�}�o$L[�������O�>����8�?x}� š,�g2/�0�OCYP�P��|Ȣu�{�:�ԙ}�'s���.X������Y���Gb�S�T>���`,���0�.*3:ՃÑ�"�:��QP؜�#:�l����17ݭ�PH��S
�"����pBŏzSXU';��/*��=��[���׮z_g%Օ 0���NE�Gf��v2d�Ux`�rjrR2hh��!�J�&���/�>}Uη@�lv�X�{P�U��x��t�J��1�0:!���p�h�9�>�xZ~�������Ws�f�P�Pb�8۾͋������xQc*V���lvM�"2�5�K���ܻ�!�X�B�F哴ML��c	A�`�p킌Ivr�Գ�4{�dr.��LVJ��`���z�zw���M����@��Nu��"��lǋ5�|�ɸ��Gir����ˡ�8��w��q�.��������{���´�|F����� P�Ƚ��/>.�!9:α�ڭ��NMU��{�f<���iq�֛p^kH`��v�o�3�ߵ�-&\zn��LA �g�H9ٽ�Y�>��.v{ӁV����P��\��yW5Wx��M[��mͬp6!�-��fDA���c{��d{��BxDƥPk��Xhu^ov�ߌ��컅M��@�(CN����~^-�i�5#���m�ܸ�@Y���HBW�Ar�k��i�}˽��i�IOC��͛�rX+�C%�w&vg��S��G��Ƌ�>���Z��8f)M*QR�X4\�Wq�Ϋ�nt[�����b�ܟX��6�����v�V�2�+���O�+��"��ύGM^S��!�9�q����E��l
}����x�6g�Ҟ4��/��djB)�>�A�9^C
�(��På%�xm�����C��S��ٿoD%�r;[ۚ�E���6��c��N��#�(�9H��P���b|g�)8V���}��#3� 0#]��T�.9�䄬tM�+�;�����h�Qw�o�ZB)�Ǘa�њf��c�Z�����YsU	Kx��V�_r_q�`ʾ�+k��QGa��{�:
	���o��~]����p�S�g:�1~���I�I�;���� ����|�����R�Y�ʛ<!����V)Y����z��,$e�C�ƹWM�~�QjE��F���0�8���T~l�fO����4K�G
�1��L:�3������nNjb�#QQ�y�]�=��(C���L��A���{��]׹��ʹ��}�{�����uQ�Eׯ��Bv��8�"�y��x�ʼ��T���u'&Œ�v�vE+Z=�3���-Z�>��>�]hf/�\�6�c�����W#\ˈ7���k^��ڡ-A]ڦ9}���(-$Q�Q�C���
����MB���r�g+=�}�u�ڻ�+��W��n&F��P#H�w�Zf�}̟Gr�_*�U%�3��w$�R~
j��c�6��J�x&c�)U���(W���8�Y�\,�0���
ʼ��=Cӭ�u1�q֮/r7��{:�B�i���V5�
Ҽ��i19ϳ%E��gFg$�`:G@X�.+=�ܾ��Hڏغ�	���x�	��]�ͬ�e__��f�*���=?)����#��!\,tk���1�-�m-H2�n���4r�9ŌS��Gk�����C����vT;Y������F�wk���@���8��*l�]����v�����b"��s��-6$톉����a<��5m��kԳ$��+;��Lc#aq/��qPGN��9ې��Yt5H�q�X�Qj7���Wz�$�e��
�r�'�"���<*� v(p��I�8ZQN��B�.��[����b�8$S��X�d`�6��B��;"6mi x�x%�.�{}^��ڗ�ϟi�l�׮��g�..��B0��3潡B���$\XG'�M���|q{z�m�a�#e�DQ�"�j�qQ�C�0��1\��J&�W��
Pm��^���p�Ks��^߳f��	���Q<B�V��s�q�c%ÁOi�6�^�P�$�*���(:N�_+ȋ��2Ɍ�Օ�^x�F���lXͷ~;�����G��A^o���
6[��@�s��r]+&��$
��:���d`��@ž�f�C�j/�ڮ�/r��"��L��窲����*/�[����PC�2P�@�R����}Q@�z2�>[5�J8xe�s7E�6�Á}���*�-�Wд4qM)3�"}u�P�h���_J�����|W�J:zo<ׯ8�M@�q��l�����2�y:K1,�����p�:�:r�n�ʬ���ko��.p}˻fƏs<��m��Q]�e�<K���zRn%����g3�κV����A�es�Y�^�Qwwh1��ַ;#Ts��lr��l�S��\EźU�p^�=G����ζ���H�T�:�VE_���O�� �2q4�ު�.t�r��w���:��Pȝ�ʉ���i�ke˼�a�ֲ{"_
�P@����$%]e��ճ8�r�ʀ<Fr9-f ȫj.M�2�E]���v�[������ѝP�lE�3�G�Q}���xs�WO�m��n{+;s���,.��y��&�f��q1K��>����˃����Փ�(�k��fb����X�%��p���z:���ڃ�=!���,��h���{{/ͩ�ز��yO*�m���Npy�
,�㡟S���lމ�� P���}c�+���]㹻(�]�̎*j��k�e^�)��xM����#.6Y8*o��n+ru���^��X��7��0�\�(�*�s�Ȋ6��=`wC�s5+y;�$&X��xbS��F�zԃ�~�6���C�����cB��U�WF2��3�`9�F܋��S�1y�/�[���(>y�blE��{�]�z��ܭS܊g/�tq� ��̵�q��sr��1������Qi
Ø��mmԸw��=��,�Rjh]b@���m����zn��.�!����8�ͻ��,�N�<�!�׽�mN��#�(�Z�=�]���ЦR�{����{J��{����<imm*અ��_X����/�x>���.-B���ҟTu�Ҫأ�[�� ��A
�L��sJ~�NV��/����lS�Hd8�ȭ���3���´q�IWr�	�=��a���I���>��M��6jUs;��n��Y��T*�g���v�S<�B�S�G9��tK��C�p)�~����M�;Xğ[¯׼O�O;Bo/.�~u�"��u9��q�����E��&|[���7�dnǬ^q�]�Q�wL)�S���n^�r�8�V�Bn��W��Ѱ]j��)z��vrM��^w��C���0�P/fK���v�`��W��D㞰h���>�AE��TG{G��Q�X0o.��)��Mj��47û�d{��Bz&5*k��3�!��R"DkSv�13�Uy��{h�ń(6Y��LJ����c��{*�7N.����N�T�%���T����Os3���M>��S׾3q_bS�z<�z}���	����PN�Ǆ���p4pZ3��Y�\�-�uwTd7/9�Ǹ�)B�����Eƥ��Q0[������<�U��S{����w	n���s����,�o�*����'d�����Y�7��q��)*ͦ�΃zZ��0����@bg˒�v���[q�rro%�E�/�U\m�G��h��U�u^�s�˅E������ҽ���Qu��z���5�3��䞻>,XP�D�<ܥT�M�R�y��7ƪ�!`,�"5��fi�z�	�:Zpߪ��Ux~l�yT9A*
����QPEߟ�C_ ��ٕz.�^{�Ր��õ�"��+Ǭv
�Xm\�;�b����� �nG�eEA��'\�$�����r�+%�T")�-��{�z�X�F�.3��T	V��3W-�8ih���ׂ��nͫ�Nũ�F�k�����=��l�fKQWRtK�b������Ê;��8��v˩nn���7.˴�uJ�i�&^���=i��D"WRJ��m?[�f�m̰K�ONe�~�X�lu�ǌ��{�}�-�Bv��;��]���[y['���<&S3�=���զ�O���C��<e+^���XXU�(����O�r�Ah��e:�b��^S��+0V7��]{���3�@�Yp��Ԋ��u�Z���U�3z�f謼�!4[ל@v��*�	�B�*��\�{�gK¬��Y��ڭ�RL�f><˰�!��]e������������B��:mu+�����o+e��J�\�vo0O�s�����E8	�cZ	���\<en���#���&y�*p��C ��֓g�������R�j�[sbhi�b��$}���S81f:4���/�LC�;�>���U+E�P���0�k0��a]f�ғ�d�=�V�$�R�����.|VZU�:��7�ٕ.?�ܴ�v�eB&7N仓��]8.D�·�Q4��+rЮKz������:�5x�B���E��R�K��D�3Ktx#�{r��)R�.c
��;] �|�o�s(�[y7v�"ԘW�6ũ��'p8Θ��\�#gh�������Y'MK{2�)o�R�=�FҼ���c]g����:M��U��]i�ȅ�{���=���B魀��e7x�Jw�/�?Z���Wږ�Z���`$&�+P>aQ�}��J��^f��;J�nK�rU���rm1]��	�h0��o���챏d�2i`�KysS�w��$t��R��2	��\��U������};��a�;S��:��\rE6s]�a���L�E���d���4�R��t�ĚcE�(�X�d����S6O=�o�U����yy\�X3S�wҁ�6K�Q�t9�YYk/8;�^A-����V7R^s\8�&�4U��oh;�{�޻�~S�B�!#��`�k���ȞK,��x;1-^Г�5��m�D��j��ӈm��VG�'jEº���wwV2�1#!wTs�";!L����5&Vu^�Kn��]ms\&�n�9�9`\>A��*�}%X�j�ޓ�3%����T�r�9�l ��W+Z�j�Ou�bm��:$4Z5�%�ǵ�lS���F��i�a�l���Ջp�N�m�����4�
�s��i�@����-)�ܨ�޺��*�):T:T&i]k��{N��ʕ�e��A���8��~��D^��ܽq�ތ��|��.�ƥ�j�}l�]f 5$�����$T�R�uz��V5�%�Sf�"8�:�S=h{K�����J��m6-oj���Y/�X6�X�Z��M,�A 6$�ij�z/J�ڌ�Xh���Y
�ieV�\녵9q�}���-J�\b��m�P5�"([`z��X��'1
�g9>���;�s�Wt��/r*r=�l��Tr�]���D�9� ;�jT��]͡JKC�r����3�Ѕ�Mm-*���뻶��{����;(c�������`V��쾺ׁ�V^���fay:���y�W=�7jAB�Sz�̡2��>�����c[yV�E*�5�Lv�֬.:��[/���5�D����:`<�N�:�����S��%��m�|�R����N�[H���gԅ�KE�P�G����9vv�:~7wLERcEb0SƢ*�"�Qb�1TETEW-T�� ����1��F,���0TTAP@U��T��Ub(����
�*�*�����TDR*�X�VUf4Vڊ12"��
����EP`�5*�TE��Ҋ�
,R"��E#V"��Z�E�"���`�D1X����Db�",��QQQ�iF��V"�b*���
+AjҊ����U+c[TQ`���V.YrՌe��[%q�(��q+ɍEAdTQj-T�-(�*+�VZ��XʩQX�b�R�J��X��"
�U�J�Q`ƫQF��(��R�E��(���kR��iK�ڬLkE�E����+UJ���j�F��ZU֖V��1(��%�5bԪ��"6���??���_o^�}Z$x:uƺ3�%��ϻ�Ehz�Ұ>�o�����w�FqU�#����^G�o��u�E_gIM+2���Kx��>�i��ׂ��Y��.�7J=夿�h�T�_�Ƙ���	����vb�c&��c��c٬�Um��5p_�����BA��\Dt]*�U�$!^�q�v�u�r������Y�"��"H�@"���3�Uc��J���2��E��L�KC�����ٚ�]��Co2p�U����p>J(Uk�_z�����p'aA�fT�nP�Q��+xׇ�꽝�/Z�A��i]�dbҁ�%��u.ul(޶S��Lt�4+F%�9�R�ڱn�[,5Y^����L��W >?w�8�Do�Jh
.����xj7��M��5�8o��Ƌ̜k����/O�y�0D�h���:A
�3l.?n�� �>t{n�;����Ť/eÁ�^�0��&\]�� 0���L���J��<��bB�̥�[�ٕ��L9�DQ�"���w�!��}+ބ>��������A�R�Y����qR�'oww�,�
�<�93�X.ߦ�݅���\n�y�!d3���%ٛ�tP��R�iSL}�z�2���y�y�O��2Zy]`]t1�#hf��1u�G�yE�"��:Oâ��U{����1�9,�nL�˓E�w��v��aB���%��Σ�ı?����\�p����ޤ�;�hkOnb�Ք��[]��.إ�Q�Y�ի��0f]���z|�7��~?Ok�U-<���k�����qu�܆#
���k&�D\�+�6(h�r}R2
��wt�"��F�I�4��'�V���7�Ъ�b���գ��>��aA��B]uEV�ˊV�'[ j����p�2f����s��S���8;Q�U�'��r��4�=2Dz�
�>ś����I�\��SWW:;eq���d��g�g :T��T;'c$z�>�����0e3�2m���fc��	T4A㡐.i)���ˁ�"��b�\��[%F9B�9ܳ,�e�ls��V4��V�N�`ck��贯 ��Qt����c���<�e��Ngv�����&G=D_M�gb�'�^U*	���цj��Q�TX�ڋ�"�6����H��'=�e[��ͩ��}b`�N���E�>ZA<����4o�
W��7�0�@1��<c�~�2�#�.zM�=i��}"�F�T�H�����:��TÕ��v�ogl�Vvr���������l$:���hD��n�
�%�>�ܴgp�0��j��҂�PPYf����A��u�7浯)̊��Xݏ���y����[Z����\�ܗ�I��+te@񙥷\:*�ڰj}[ڦ�+m�\��̐����=-���P���u�V�s�PQf��C"�^G`lۡF���g�C�&�Y�F�ղ�ݯ#����|4ORCǸ�di�~R���^�Sz��_&}P㌸~�N
��		%ԸU�*hʥ&�/޺/���ZS�ei�s^�dQ������T�K�N�	�i�dP���5��"���At4}a�=�RYKBA���w�An���W{}t�l�rs��=�#mn_+��L)a����!�����j��z���r	�\�,X����aI����"F�EGì��9��w*0[�|&�*�%U嗷�x7�F�v2d�p�V	�9꜀V��*쪅D��h�-9
�_U';�@�lv�X���o�Nl��ᢛ{�P�2/S��-f.��.���R���$nz�(C���C���a�'f���Z�L����y�-��hZ�J�bX�W}���.E�T�q.;bB�߶��iש��c��+l�}ۡX��ˣ�����E,��^5r�O�<u��iF�<�T;..��G}w��)S�w�jsZL>���/*�u'f��}������1Gsw����,&ސ��i�9���뼋�����gfc5�֮=�@-m����@Fn������Ů6���s�u�Ҋ��g3�dy�����f1����aV���91��]����q���ڤS�5B��Oi���z�(���Gw�F����7�n����"x�����%b�Bgo`��^����MEW�ho���Y��4�����9C���z�=+9dg��V`������=��Q��LJ�����}[m�w>>hx�-�a�k���xa�B����:ѫ��V�o�w���v�9)ut2�߹:ٕޗsQiQ�<�PPZ�f��3������8�;'ԙbt3��[��@4���u�և�Z����\9q�i��+�0p�Ƌ�
FH����L���j�d�]*i�/�xWU���G�| *b����=���r�q�Y8"�͟@�*�4WU���F������~~�K����DEl�<ͻ���9������(Ъ=���U�CB�� _��H�B%G�.�!�r�N��<�:ٟ1���޺w-�ķ3������q�5$pT	VǏ>�'"�*Nf��(n�H쬖�
��c%E��F�k����� �>���]{����8'Yy�6i�j U���R���P��Y�\���:�[��بb4gC`E��,��~x(��:��/���KJ�/"V��|��{��j�x�c�	���Eӷ'A		1x��xk��4�m�+5;*U�F.]Lx{#�}��'"#�{��[�9Vn:�r3)j��ȷ�)t�S�7�M�7.^]�=#���O�N�K�[tc��[˜��w�QS�����!z�?���xc�0�kNWT�����C����8�"����n���O\V�'C�z��S���g�;���>T3�V����X4����}��'�N��3��fU�����S��s�S�8����c>��dT�	���aΞ�lg)U%ԛ{��o\0���k�߆�q�p;E���<Wt��z�]<��^G�VkX��ޭ�Q���S�uĵ:3�ۧ�M\5��#Zu����-r�rZ՜@H����rsZ��1>Bi5�-��ʀ}}EORȽ�A�3�gTH_-5݊H�����.驳��m���,�J�Q�	�.\���S�s�������u�Se1��c��ŝ�����@�ja�`��<�0##���Jo�aq���>��9�S���/�Sȼ�[�N�\��a��Y7S����aTG�/N�"�糏ۗt5g_Һ�#K���d�ai�⽖7+O�T2�j�sA7S呦�����Z��շO���k�{��w��,��˻�%���+�X5�!�co�D�\�ѯ#�C��ͅ�d��5�W8�w�n񔶸��u6�Ɲ��K�����EL�DkB(ٷj^�>��S��Ej���m�PH���бc���.���W�F�߶�û���G����t��`쮝�:�W1��`L���B"A�n��(�27Vh�M{o���3w�MgȾ:*R"ʪ}Α�"�Վ�������s�2��Ȑ����0n<+���W�ޘ�(�^�Y�������ezk�n[ķ(s��xx}����6��72�=���^�V�$�;��mCA۾]S����N�&|~���U����^g�s��u�Dڼy�u*���E�4�dh�Ѷ�d�����&�dd�3���c*�1�5Z5�s�z��m��0kh���v&����{��i����=]QU��ˊV�'yr�YҒ�5�{�O��`s���Q�s����{�}Z9�\��m_ėfx�Bm��w����]J�~6�d�ta�M8�1	^�:���(���d�g$z�S��:T��g�+7�^����KѤ"*�g�'(1��\JS�U[� ��^�E��vu|��%^0��u�M�{�y@�w:��ԝ�"��\��w��/'d�h�;��3*����������r��c������s�0�|�AeJ�����b3V�O��@��bw70�֌����:%���<���vk����5����������R���D��WGA4P�PODÅ
;�Ql/�ؼ<r���.�U�A��9<z%U���RӨ{�.v_h��1P�
��mC�
=~<ʌtT��y�bw�c�޸��t�ܰ�c�}��L�;�y�U����M�ܚ��0��ٚ�'�,ql^�=w���6%GG9%�Gw����u��R�"
��^�S2#���OR��v�a�B����OC��wh�����[�R.6�<����葐�
c���WJm%n��Q/Y���2b�_< ��^�^�EEᐾ��N�H�
���:s����]�G�k�������!F֚��U��L��H�UJ��ږiL:u90���ҌS}�{3{TG8e��x>@��*4�Q0J��Ì����V��P�5�S3OBؙ��m�kc/d7�08�QP|�Lߛ�٫z=SCL9�����n�O�3e!Q�px8���3b�]4��5](67M�7ʶ >I����/7�E�.g@�>��X�"9Ul_;&%���-X�N%�+r,��&�N�cs(�3�Mr�|M>��:��ق�z�V%Qc���uv�����u�17�AZ ��x�;�uq�1�;���nEX�`sڴ�GM����jQo7���K�ծ��h������>�R�jR��6WF�8�+c�6]����W����n���2:�$��ɨ-U��X"�*�1�Ǐw�)ݽ�*^�LR���LeNz��tJ��C�p)���lXo����V"5�bI����$��ğ�
��1�,O�֬�������/<��h[ �.��Sۮq7�e�d06��lcH�R���P͇[Mx:X�Q���L֌��p�W|+��8QՌ:����Ƨ�R��_[~��W��ސ��ޅ��_� �����z&Z�^��F��C.n�u�i��P���/�K���ARF>�:�n��6О��Ԡ�Ƅׄ�~5Us������C��I��-��Gݫ�pp�.����o�q���F�Q�"5��7mBx���ۥbﷀ�m(�P��)נ�j���A��\z�w�)�'����A�^.��c>��#>���ǌ.T?<��i�]�W c�Z�=���:���|ʫm�.Nay�A�Z�Bޟ03IʛR���(�UT>�m*�Z� ���vָ)�Y�/��^��Ǵ��x�ԅ�%�Rݫ�>��Kh�����t4����ʫC�en �Ц!҈�1 4n.yQs�u�X/M�0Z�Im��ҋf�h��Y��ɕ)*�:��\�ש����w3M;�A��n�ַ���ǫs�)v��fn�Q.��]1uI&)��9�;��r5��;��-�zY8"�6}��r&�T(��PåEC��U�}���`���&���#��p�*���`��'A@��{�u�$���R}�'�t�|+����;RU�܇�e[���b5O��M���d�
�E1'�ԅ��}A�¥v�/k�=�����c3ͥ��{�.�@d��
�>%�HtZ��5�q�c8�zi@9�϶gGIult�]�M�u�}���,�%��"G1Q�,��u�����i@{�n |�{/��ݛ��Js�EՉ�Z��'�����&(�4}4S�ٍ�+kmVx3�������xm�P�<�HA-Ȩ�v�j֧��A��<Z*�g\��I��됇�WEqjס�����.�@��sff����q�����	���[�P\�)�2�`cu}5�Ϻ9�J��0�:��i*�;stL2�*5
7#+���\�5�����9�h����X��=�sj>V::���Y�m�}�g
���R#8��z�D|�����a�t�~���R�0j-\��! z�f��^����;[H ~[����U�];�[�d�rR\N���4�GQ5�W\���gd�2�V�d�:6V�)i1�+�q�{�^�߻$�0��;�����%p��u��B�u�;ToAw3���%�c�y�VmQ�`�4���P-+�]]���CZ�n���q���2��Ε���J��[�U����*�zR�����z�k��7�{�lfѽ�ϱn.~iB8��H�
���F��Z&;TdFb�c#5��ss	,�K#4�b�L��ⱬ��u#PKڮG4}CL�Ն�+��n�s.5)�ѹ��F�`sJ��2���8$�pqhb�[���u3�9.T
�()=�@�doG�o�2�dC"u8[���<�\Y�$h��\�1��O�%�����z�8���[�t�+ٸ�"�#R�]�{i���������Ez��.�лv���v9�c/"=���]ɤUV���]��C(��$��44:�.��W�뵄�ْ4!3��0��چ��ow��!��6���F0h{CF������}I�P�-�I���q���[����N�@k��	R�彭Q��ۃ��.� ��y[9Q� �4�voF����v:�3l��RM���ZjW�\����d�|"{w����cS�l�78$⾡|�]uN��uܪ+���TA3��VXz��Y�h}]����;���U�}!%ģ)Q�{��K���ǖ;$&�;X�ʒM����:	�,m;���"hŵ��2;W��W�V-���Kl��h�O����F,.����7GKX��Ѵ.a���m���t��R�ek��'Q��7���H�*Q��8�a.���L���]e�5�	������7ǁ�L�����՞F��R�oC�f�[�
X���5�ʵ�k���(Z��1��d��������z+�/oJ�����Y�7W*�he:�m��4����k��l�#�J���CM6ߋ��\�Ϻ��K�!��V�	}r����%L��3�HϗI^���mwF��l�<U�t�rkn	.K�i`{>MK�)ASu��[3�i⬂�����]�����D�9(̌;&����t���E�}��)�@ނ�һ���T�o,�o�P�w�@�òH���M�[w�ܣ]�O�_"��D��S�E��7q��c�6�]�볰䡘��ۄ\R[Y�6a�w� ��<Z9����I�{҇G���"{+#���o]ᎈ+8fՈ�I�՚Ǒe�b!�8����.�X��l̮����"[��I7��������NY��hR��]S.�S+,�]-Zjd҈�آ&��f�;v%�\ܻ��P�M*�M�(�ϳ��9|�i|Յ�%R�gM�[��cy*�hÜ�v�j�����A��E�;f�Ŗ�ZA���U'�R�pd;�N<�(��F�#�Z+�ԃaL���u
��VO�T��0�ef�f@���3ֱU"���𬜴Mo+��"@n��$��Q�'(K�F�R��,8�͔�\*�wMH^�T���[���묫<�9�h8v������X��Ɩ�!��7Y�q}��>b�>o���t3[�p�ˮ;��C62c'S:�SN���+�gJ�x��27W���Q���ެ ���C�!�#I��_UɨRU��`���QF��t'G�^���TO�������g�Z{��O]k��t����蓋77oV�q��-�r|*����`Wh�]�%�ѧ��!�lШ��q�\h*�b��kJ���upP�uu\��>�2=LC0FI�;��1������i�k�u�[U�C�}�����R��d����Ff�a�Q˘x	�,�0����շ&n�O]���O*Z��E����X΍�GI{3d)Os/FW�F�w`�=����f+�!a�����Q��X�n���[+��F��_3|�w�|�`�W�2m� �i��p�x�U���m�t-=/o�>}��|� P�P�`�;h�kml�V�D_���U������)mQ��`5lV1Qm`�6�-���B���-�Vв���1D�X��J��kj0�
������J�[lEejҕ�DT�*��S--KRԩb�m��bԨ�T�Am(T�lZ*�9�����)�[cF�Z���VQ����m���Q+E--V��Q��hQ�b�*�[VŶ�µTV8�D1Q2��f8��dQ-F�(*�F	X���V�m�`+j4V
�m����RĨ����cU*�"�#j�U�*�X%[Y��f%V�TJ�[e�h�%�eUY�R���K�Fb�kF�Jʨ��*�"�
 �X�QRҖ�R��ikchU
[liDJ4U���
��jU�
V�E[h�A� �K)P(V�f��5��!�=�ٖ�m8�¶k�'s9j�p^�PJs���,ؾӈG�E����U����vB:�Bn����C�]����������K����}{4Cˊ@�	Gk˅�'w.(J����3VkFt��(,�M�v��,O;5׳���y�x$�1YP�eپ���u�?ia
P�^
�g����N���a�˜��U#n�����$��IcؔQ�1�J/��K6�M5cX)���	l�r��=�V5�t'_��r��� �rQDv���<��>�)�ޡ8����5�G5���x�Q�ջ^K�:X�cB���7�)
�V��ZK�
�{=��׬�K��4�}�����R�C���ۂD�t]�7Y��v1�ě'���m�6
�ue��ⱬ�ZFA!1z`�纪x^j��$7�UuNq"�;F�a���|������3�:��ͫ�5'�2�='tO(q�W�΍*�C=i�U{���P5C(/p��x���!���՜[I�� �}C0�IW-+.yу㫩.���2���7{�W��|c�+�{�jͫ�WLZ�s��6%Z�\���Rkk(����l���v4.���78c�b�sD\ ԝ�oNb��]�ܞ�w�.��2H�fPq�Q=�(9:��,�����m�l�d2����"�}����Ey���E��iz�/����x�@���6ɉ�����g��S����-���*k�WQ���A4��;�����䥛oٛj�n��b%5�p�	�h����.���.#b�V�5����]�ͻvz���X}�I5�k����htDB�����֟$v0U������}q(<�ja�v2�3ۺ�%X���x �n��ǹ�j��/6��`�-���r�Š���yN�g�'B���	���7�Dכ]*����9\)�� D��&���Ȭ;���qV��Gi��\���GɦC
.U�1{�y�|)zngQ�a>M����w������T�]%��
8�8׽���!Ǆ���6���1�XoG���w��\`9o0'���ql ˥���̼��:��8m�A0�O+�[w�Q�-{��%�b=�u�B����������q�YR���*I�T_B�+���Z��pkf(m͋/�}��/�'v��}�+�>���N��qm�кw�8�HI�$Ge�6
��	�Gc�f\l��Q�uՃsq!0�֨ODU8J+�we�6Ws�}��T�U�`l����c)_�����)4V�O���CH��[��]������U2(>vi�]��nvFi�9'��PQ>CTjGU��\����g�NY��������`-%���Ĵ�j'�b���t�Z���=ЫbP'��)�/w���^��ɪ���!؊j*k�Hъb�)�4J���3��r��}&O+���`��}υ��*�!tT��=Q�/˭C��j�!�]��O�:W�������j�n���ib�sA�XA�=��)&sr�ѽ���-K�Ps|1��b�׮���gqA�n�=;V$������{��e�7�`}��G�+�>���s
�VU������F�&`"�f�.��-�ᇷ�ah������L>����i��
�;`�[��zb��I����ϛ�ΤIP��(`���[yl��U�`�_m[5|ҒT�88;z�(c����R��n�:-ʑ�,�T_cR�J��%utAݣ�:�3����K�I،�ߙN'J�-��S}�5����E[=����׳D<ؠ���J�s��Q�@�1q5/L{���#t,�I'���a�f�vu���)9�<(_r5v�f�KS�=�S�"��4�͚N��vL��v%���v�s�.[$��B���2m��!-#�Z*_".R g�{��cX+$�,sҶ�Jb�<��yӬl�P��BFƐ���H�⺵�����Z*��6�9V`��O�U�m���/%��>�w �S���6}�k�a����kD��w�.��M�D{�}r@�������F��Z7#+4T��MDՃ����כz�4� �B{�]\�d�j�#�����ǌ܂'����s���� Gs#�j|�=O��/��6pI���q�Z��´�����\��wH�t���ގ+T:�	�e��2!��.�ջ�#8)ɞ��ǳ(��]u�:��4��[t�ʍ8�is:�n:B�� �S�#hK��ql��ԫW5Zxs��TW{r���
f�
��-$$*��g
(��v}��7ǝw��ܲ�-�d��O��̊�5�9�hӬu��3d;���┎������N�q=��s]{j�ù۾qO���$���Yq�
�m
�X��#��2�QSC���i㓙v��Z7�v{xe�X�:�0�e��U���M�2��8]{C+�%�|.��R�I��� �x��I'/VNg'Ө���9��ק��ӳD�(h{�\]�&��K��؇�D��M)�����(n�	�=|���+�P��o+�V:�ީm�	%�P7��ʠR�H-�5�l�!=[�^�d�A�vn��cT��J��
ڜ��
�F��l%`l�i��{{�DGsa�J߮���y��ӌN͆큎�� D�G�)b-�4�徵ʺ�\��J���)#s����\!o%Gl`O	k��iZɃ4���y�ƅW�����Lf�+��j;�j݇/%ߔ�R�`]�O�V�nq�edU�7�4�E1p�����]ʛ�>�����b�l��z�ᏕǙ�������XP���$�{��t��:#MwD)���Kn5V�|�޼m\��L��)7����ޖ�0�,m����:3�D��
���*oK�z���6_|��k�Z�����M�����7�w�M#�lq��ٗ~�@^��&?]H+�lJ)����g[�Z�m�6Ws� ����:�B�2uV�59sj��&z�k�
��8��h��4��/������؉TKDBކnoq����L(�!�Z�'"1�Ѵ�j�{���@�j��o�E��{��P�"ZL�Aġ��������p����塶��T�׻w|����1]��M{�SQS^hłi�W�������,e�mV̱y�ծ�^��jt&�Ql��*t9��\1|�!z/%&IĠ��wu�U�k��^�@��IJ��)VMsW̱7�z6�8��ಷW?Y~;js
�+]�7ž��ҭ7�>+j��s)l��Ȳ��Y5�O���h9�z��S���>���0��e�0�R�̀����2�Yy��hTli��
-��:�
��|Mj� ��ׄ F��fl>X|�Χц5!� ϼ[�kSO+vY��{�.����Q'���F�K�H�u�32[_^����u,�&�J(i@������z~|yw�R�]�v�w_Z��S]˹m��7��>��!�� ��)FKyYH���Y[<Zi��e��M�1ڊ�Sq�y������A��N�� gy�$�Q���"���.�O}Pd�*c<�`��n3�(ܝM��;hH��ݚ�nȫ7�j����%�<֋��視�Q���ͫn:�r�����1�_^��ê޳�F&���."�H-�k��=����H�Z���FS��ث�£j��M]�N����R�DU:�P=��[�K���7�=�t�F�*�z�S�0��7��)H^ީ#ꭡ��n�}��xE���V�,��\��[U�����us��2Q�CUxH�:N#��j���3�:��I��\�h��5󵅢D���8Ӂ^Aġ��5��ً<�J��Ǘ��H=��&2�I�.ƨ��D�h[�v!���}���]�"g�fܾw�BV�B�o��ke1 5��i�ɪ,q��.��	�hf��S�a�v��5�t�kYS�"��T`�;4>DE8��8��Oc7�n���(�;��D����8�Kc�3���ZcS��ؚ��%�܎G�o Ξ(Ӿ�饽'0ZSW{n��z�Pa�����W+׮4�혴+]�OI�^Jy��z&�ʼ�.���V�6�֖,6�j9�&�ݝ�K�=�x�VO�A���U��ӘU��Wk�-�u �)��W�"{2�3��*��Hz{���-\V���\fR�+*�oU
t-�ps;���� �b.�g��W�NMpy�A�0R��X�*o��
q�Y)њm�Ec���x3�V�l�u�吝�ErrN��#�PN�e	�]G�3�����=���Ħ��m�|�;������������{(�Q��:S) �δI��wczս�ȓ�ם�G5^���ˠݿd�OXsЇl���R���⺵�[;����7j�.`.�Dc�V�䱱����.�v%(�y����R2;a<�#U�n�!�D[�u��,54˜Ehӧ1nu�;�'5���wԊ�O/q�!�����{s8qyJ���7���c.���\/h[�wu:8l+r��� ���U�y���50{�l�n;o��|��:�m�E���g/�)QPF��S׻�9}�a4�=�q����e\(�/o@ig��w@N�]
�gP����������H�/Q	�-us�ZfB	{�"�v���'MX���J��
A�$Gk>�ݎiZ�Z&__X�i��8LM�؃ݚߢ�!gN9�����T=���n�uz6�fw�Ł�-Or�Pγ((ዽ5جP���ҫ}��߹�>g2e��$��O�Te��ɖu��]�R�X��҉���\�>r�:a��������{����4�M��y����p�S�݁W�:��1&�]��4��w#՝Ln���oK����N��,�b�+<���jњ6E��r9ѩ��حwn�S��#���������j>�7�ش5���-���W��{�]N���.�[�Qn�j.�Ok�����-K�b���5��i�2�.�7�>��U����d/E��k�J���y�!}���2��hi#�n�y����]�'8��u[�9S�h�k�=��Aъ�]qjÑ��[:�M k��p��4�Jktܴ�p3�T�/dx�Fh�;��m���+�Z3.�%�vK�%��s������l%cf�Mp/(�F��=��U�!��ӹ��0�~�bw���Х�������#���/xf�S�ee!�S�Mh<|�jå���w��#���S�C]z0B�ݥ�僲���X��㪟���Gڷn^K�=�*5u��e 93�b����w�z�z����������l&��;��2������禎��d����XZj���O���|l��V_q	�+�rJҵ���cV
�F\m,��p{��BH���Up�ѭ�i+4���Ņ�J��W��ֺ3U�X<�p�hg@ֲ�Uq���4��P�F��:��.3k{�*���0�z!Չ>i�A�!���b��\�C��&�R���%Z\��^��o�>��U&�;�b(55�
��1D�R>=)#)|�s��?Y��v#�H]p��x+)���IR�Kϻv�C��S�A8�)�,T���V���L�*�(;첝`�E��A]�|c�tT�H
v�8rsǢ����׳d��_R��z��u���r�c�7��z��"����Iv`|�^m+M���f��l힥�JwC��3��ݗf�����6��%�B��7V��#/]$U��qۻQ����O ha<�-;� ;~��d���J��ˠy�;�9��-\�Ӕ���2���Zo���#d^��MN��6��^<D�L	�xT+���>Ӎ���Y3�Vg\ռ_cqX��G�ޮ@U�F���u��jԳJ�#{���@_*WֶP�tp�ƀz���M�5�Y��$��9k��C籙�V�!���v*�vS䦪��Ȁ���حx�Vڬ��*Wi�8!Tz��*�iڀZ�A�q$����D�i�Y�nI72��3E�r��z�+�-�Ɜ*��PԆ.쑜�f/t2H��`㊂�ԱՃ���;�~��Ϭ�aEZ�kh�w`S��$�!���G�%vSK���5���v�³Z��)��ڇf�BV9��	ˍլσ�w-�Ic}�+d�ei�)��c� ����9ӻ�xRg�g7%{DU�}M�"��Ɣ����بx��Ow�8�G�X)���uJ?4o%,��I�*Z]J��M*qn\���;]l������o�78�#���R��Nﺷ�i�{v�Sٺ��c6զ-<�z�������SN�݁j��^ٗwi,F5O�K�n���!FJQd5!Q�W�	Z���y�m��2�>��ȭ3��Yҍ���W�AC)�T8w�Y���#]uպc�E,�<f��
��d�����i4�YXփ�لa�V�5�>g%MVl�moG��r�0p�b=>'�hM�ן��i�Ra�2 W��wS��~1��(fuԻ��v����]����E��i}��dB��%�sw��0s,��3N�����%�al%�1J�Ru'b%�Xlp��5a-��`�V������+6ѷ%e�VՒ� ���VYt�-�"Ym���Ʃl��]�syڣX��a=�eud���*6U;�T+SU3,��e��P�j�y�+�(m�J^����5RnL��5N���+^.��ڃ���d���귐)Mipܐ�i�V�x8;�I��X'_wH�EC���m=�umn��D�� ܻS�/��
�TG�5�֌��һ*$kL�-��=���*Ȕ�m�GP;�(h �4�ڼ�.��F��ڧ+_mx��-��z��.�L�Z8^$-���$�ʮ�X���Yt$�2�`�t�`����e��,��X����2_c�\臬�b��np���iV75�,-5;��(;�MZڈQ��],ȦShh�C8'1-m��z(�\���BCW6�_C�x�7Q��s���5'b�RD�Z�f�D�P'}�**�6\�,-�s�������w�+Pm*�!UB����-Z�Z1m)Ph�mF��B�kU����EZ"Җږ�V�"�`�j4��li[lc�1�U���T�X�P�6ƥZ���Z��S(6�P��¥AF6իlP�֫ZJ0mh�ETb�T,��,F�D���ڂ5�ƬV�kEX�+R�,E�l(�-�Z"�ʌh��J�)h4̕��T�R�Q`�b�)V�Z�����UR��-Z-aZ�
2ZY؊�TX�T
�`�[F,mJ��1&e*�ikڥeH�R�b�*ԪŌJ�EX�R�l�Z�V����Zȗ2���U$�4J��b��Km@YYDR��"�TYU%�A�TX���+X���QV*$UTPT��PZ�lP�E�,X5��Cr�X�m"�UV�
��� �֍���R(VfTY�-��J(��V�-��0m%����6����[d�V�@PQ9�8�����ɸ���i�ujICe9���E�ф�0f�!���\���v��C���b�'T�s�ڑ��6�n��־�(?Q,�
v9�0[SI��[9'Ϣ����1��������'5?u?KIߪ��c�[��{V RR��� �٩�K��:�ML���^J!�G�ɛ�J�g�-��/`kž��ñۥZo�dZ���3s}��~�Ʌ?��,�k�ʌ��"��A�L>3�7|�]J���Vy�z��mn.��Zri�����J�)����x���+�1�&a����Ƴ}�I�W��v�e�vn6�U��A��N�+����gܷ���&ߏ{݁z�3�-.4���!�v,S�=a�Gj7�Jr�KdJS��y��تB���o��o:KW�F>� 6�ߜ�J�f`гU���� �ю�`�4Ă�Q�
��[�0���ܳ�w���[o�𻳯�F����P����,$}T�(�ڈ����t�e�c�<]��g�\xJ���}{^��kv�#R����𩦦k�u]�tgi�2V-=Q����V�[s�.<g;���c�'dF�;uyy�6"������*B�1}[_Lwd(	�7���Mh�k',�zh�Kz�o��,�][�˗b�Z�J��$ZFBX��Hi��	l�ս�ˬ��RyK̵�#��n��_(xy��@ZfB
0!�5��\UU.�����	�Z�Z�nqF�z���Z&_[H�8��.K��Pd���`�O��o?ep�n&{�~��_�D�h[��56�.xEӣL�̒����-9��Ne�7zUn�|�n3�W��r��X�R�f�y���gK�4���M[v^P�Y�ʮ�-���<��eE��Q�e�Yܺ�^YXoώ�QS�C�Ꭷ0��[�v����×j�Ã��3���S�65�=��ק��{{4|��{C�Ѯ��u�<�L<��Â�+uZuܛá�w ϻv�!��q���6��`�n�q��c�$���w0�}K?��A���սE�)��y��OX{�(���:4H�.eSv�ԭ�E��w����w,�[ �xL�V�-�Y�I������Y*��"�+#�P�>l-�	���hd��\���s�:�.�H��P��M�Y��_8�讎�ST=Հ�%o�q��.pEaS���C�s�eYT��.q%�(S�zY��%�?l�w�۰�e�v,�����y�O���x���7�_����w���/��H�����kj��s�ήeWW�z)����P�D8�	}Q�J�Q��֑�[U7����]��1�r��L=	j8���[���6'���`�p�m�{��� ��H�cרߋ�t�H{)T��^��$4�o���0���L��T�nu)�;Ry�zyV����z�	�-us���PA=&��j��윞�s�Z�t��Cվ�ݎiZ��>���8'7b�b��#3��e$�˸63�F�"��qI�����j�[�4s1b�=1z ����Wz���N0�|�s��5T�b�>-���W��n����6��X�$�Ǳz��*�����䆢��*���uyWjb���G�V*m;d��ׅf���[�o4���yV�f1.:��dSR����XN2�]�����oXM�v��k�[כ��X{}رI���$�0�Wroegb�o���ms�Ὕl5��1�+9��f�b����!�Vy��6�oc���.S��nV��K����Sur��G^̪��(%�R����]9���/B��M�Mna�a�W�Pw�X-�{]g^��h�^�}Ϣ2uJ��wpդ��Ĵ]�͡v��6����=|�Ǔ^��<��<�a��Ճ=;��ߩ��	W9�ج��l] �5�ݨ�em��9)�j&��ij]{�޽���7\)T�7`WR"��l%~٤�m��Y�]��w��Eqs����Sގ��$c�NR�h�H.\6*x�[��N�*�O���5�ưQM5n�;s�;�G;hzF�</��75ru4����o*�����E������5Cj݀��	ib�hzF�lJژ9��F3.N���*�b�<�ﭣn��6H���㏮O�f[ٹ�n��ҳ�wS7
3֜���UuJDv����]ά��������b��b��CN�#Z�SȌ5�ڶ�X�~��e����Ak�����@#GA��P�7 ��HFd��@��kh���n�Ij�y�f���{7.��C7�l��7�%��ܰ�E�hX�up��RY�v����X��io���H.+3z�R���M�Ԏ׵P�� Um	�H����n�IY���0"vs����{�v���8�8��R
$!�R5��'"1�
�]����G7,�4]�{���>��؇V%�S�8CU���t�FEEuϫB����\����<C��\%��5K��j�׃%v:\#}FޟL�r`�%ΦֱV��Mޕ[��݁�)�S@&�Q�g$����	(͆�T�V��wqN��y�S��5�g��ߒ������IM�p�i�zЧS�M��ĖE��j�uC8̥���^_���z�A��
<rH��F�{��;���-?=��-\P�r�R�&�S�M�\�i�ۗޭ�l'S��}9��U��Cz���w��(`�Br��VR��E¾��S��X�3�O�;�w�MߓE�e7ךk�=�W�)�*[}J)��0��`���=�ù�Zoi��	����Z���c���:�m���z�|�U4��J/Wo��BhYG��dÛqN׽���ɡ���c��q�-��a�U%��%Z��8��]׌B�_E����ү�w\d�q��vLx���'� ��O�^2��9���N���O��;=��ڈͪ�MS�
u��d�k�LHKMV�_E��7���z�GGոd�R5�^��,����:w#a��R0>�,�Q����*�_�	8І��*��wQʶ.^j��q�|e���q�=��A,N�)Ex��;-��]7#2�q�f�IWV�^k�,|d�R����RF�hKf*�Y�F�Z�umR݈��'K\�v��z���>\%���rH��i����ug/�o���n��kV��ǭ��٧i����4�\�S�r��ë|Ӂ^A�N`�UU�{6Ms9-s��Ow1C��M���8�Q/{ɣ�"5�H�;u��Q�Z��;�+șcB��t&�;yV�׮��^�c�Sx'&R�{��`μ�`u��1B��hpuC�*����y^�XFc�W�[���!غ�=�}�j-µjf�*J�	d�u�! �*@�8�]p�V*���^Pa}R�\v��)��g@X�q�b;���VP*�Z6�/MP��,YL����:6P�>ӯyݥ�!8J�]���'D<��f�GOґǜ9�iF1���p2���|�w2����T�\�������!�3CC��q�JK�v�j���jm���������qa�A�n�|z^��oof�j�C�Ѯ3)�qUt`��Ӛ��y�������R���ef�}{4^l!X J+tc�;3����o�tר9�!̇[*���a��<��n�z`"��뽹6��U>M.��4Z+�	�n�����N��۶SǪ]ـ�Sq�'��E浱��#�u��@���*��|��G8�󤵉�ݠvc�v�E�oWn�˻�����W=�l~�J+ť�w�JaŷDJJb�Z��4��|�s	�Gc��^K����TԻ���t���8�˼�'Tf�<a���;-�]XM"9�,|d�Sá���=��g�b2E���Z�]��F��B�Fu�xZWT�r{�Ƴ�iԌ���w�82��JW��"��I��˛|����iu�8��6�كZu����$v�ʁ���\e�����[�ˉH�7��ldo7/0eLo�l������ʜ���N��)��Sĳ���\,a����Ӊ�B�gK.I�ʡ�]6oKkot����{�
��^O����~0����sJ�����Ƞg
+g���-�k#�PP��uH��(98��z7���P�c��yJ�o�|V����s�2#���O�TOb�C$�=zU���a�S�v��ۻhi�Y���U��p�娙��WQ.�
�tr����햡X�a>j�e��걬�c��,6�{�)����f��\1\:c�BU��"�aju��%1v�2����@��I>y��2{�����%:�;��Xd���T��%�q{(�Zf�3M�v������}y�v�J���Go����kJv�+A��]S���e�|"��5�9��9���ң�	�]�l�y�����̈́A��Ӕ��R7/�[	`g.��<�\Y�H���sSgd�x(���t�vi��h_?��)f���n�V�Dt��ea��}�3Y(�>�я�O���4)M|�pJ2v8�`�S1c��,��^_t�ǹ�m� ������LA\V�핁-��I�1�y x]�z�S֖)�WK��כK��U�C
R�\��h���[�qt����d�S9LE6l�/4��j��w��~�4ӕo����䢼Gm	5�k&�o��3\3��A�N(�F��N�p�����E�r�]�O@��;���m+ZL�����;O���(�y�;�hۻ������ܔ�������}��0�t�'6u�t���CT;���+�����ᛆS�yBl{#���VW���unU˾FBX���4�V�*Wv�nP��v���j���;��飑����i�� ��F�E8�7�u���.���K^h�׭���'���ëZqA�(�ĚW�sv�q���1}V�^\e�~ֲ*���Eߗ
}i�&���b+�������W��q6�U�-^{�Ot����;�X�u]�'J;ݗ1�����ɿ�X���+ȩ`pڬ��m�F��a�v��K#V |����uW(g�ʁ�����lx:�ﺇ\��L`�[��i^hQ�/�VV�r�A;2�7� �YԨ�\̈;|���Gz!X����o��7\�-t3+BҭV=:m���u6+����:��Ÿ7�����h��	��k/�Y��6
���vo��7ݶ���^ϧ0��ī�����z�s�l޹�=���n�\�u���u����F3�3+��*�*�oa�'o�0O<��^&�f�ϐg��l���m���>y�\P�H��\(�h企�K�IvIL�PS/�+m`2�s�����!��Yu9]�|]=�{y;�k��@��=�)��l�w�e�e�v%��"M+��9��S����e��"�fX�\Z[���/��q~���7������5x^$�[;���R"���=�M����:��@��UYuV�J�{<��狳��	��>��60�O �e�t_��R����/c/��zK9�%>��8���FH	/o\���ޝ�#$��;�cN����6ﭧ��uMjy}a��m3 ��{Tb(MgT���R�嵋v\���Wtھ6ս��#���n��c+�n�]Y�&4aJ�v�/�����֥�Z�xY�+�ۆ�^Н%�̹l��[_@Jj��P{&q���Kk�Ỵ� �]c��k�|렝�ݭM␡�t�P�Lt`c�CS�&WaIZ6i��77����1㬇�ӂK��쫴�oh��٬�y�.I6�'0si2�o+ǘ�mͫ{�i����|r�v�ǩQ�!9���+�Vj6���צnmHm���";7z��C[���H+�2�!��۩��ָ'��pS��zsU	�&�4^$%2�fٱ:�����%xU��XA��D�
N���M�S�3����J�����EAq�؜���-�u�:�����{&M�G1^�As��:�u3r{�sd��:��_9b���JV���%�����R��h�ҕ����f�qkX�m�Ks���.�oR�;s��4��>ݝ5��Z�I���awn�WrE��ӹJ� �Z�u���w&�9B���]�g,ME*I����r�}k@�y�Y���=e���	�8�/��$�;�E�=�VP����6��cFE�O;c7/�������b��h%gL���mԧ��X�]��Ee�2�6�����ۢ`,��G�@Q��+ ��Xx�;4�Z�ia��\"a����n�)k�t�]�m0��>�ohaZ}���y���Z�E]L�{�W���"O*�Fʼ�#���:�}��옥�u{��Km��� t�5v�Ed�n"�#�u��p���+.�e%�������z�����F��u.�n9�r����O {�U���Ȟ�=� ��܆�jw@�@/'F0c�h��n�LA.B�+�K�ѧMg9�vq���v8�%#q��H�Wf���w酻{�3OS`��2������HhX<]��ź��c9Փ#�'՜���:��f���k&�����/%]龩�maO��u�[`g-���M�'0�NY}�W�λ0�����!��"꼑�������S��}��|*�uHa�sqE.��)�&�g(��낰se�-���z�a;�4�M �ՋS ������J�n�9(h�5�����|����(�Ͱ��nV����eAғ������ �~��Ş��jJ��B�)�l�ۨ�
ܼ��U�u8@���ᔫ��VԚ���m.��8���`yB1��w
\{CЗN��T�WfH)
c�4����{�K��
*՝H[;�E�K2�_R��bX%f��t\n�_���ɻW���|#5.��a��M��G3YC�hd�,�(���:���f\w|��+6��=ܝs�N�i�=V�Jŉ��lvB��r�ںN�۶.f�#����Y�_^
D/U����*NҚ�z��n]f��$��w�D��������}��w�BO�/2_f��T)�G��աn����:q��>�ETEP>-��J��Ƞ��0L(�!Q�*J�R(�Z�Db�"��k
��
(�F)�Q�U��b�¥UE!YV�R"��Q�aZ�J���TQ�Q����m��ʒ�ŀ�J"�1U����@*,�[h��#(���(��b�@��
L�B�����Q�T1��VehV"VE
�2���(�)Td*AQ�ҩ*���Z5X�*6˔�X����q�YYYX��H4�����dQe)dX)PXR�cF�T�# �V(�`Uj@P[md�(���ijFT��*(��V,
���Z1AdQkm���AE�Q���2�E��PR�B�*��Uk�V�QUUA`ċej�E�("��؊Ŕ� �b�-����T�1W-�TTr��Uk�S0�X�
(�.%bŊ���DTm�RUR�DUED26�UVE",J� �E
A�A�Q�!�2jPL8��h׷�E���]��ĵ�����-Ӯ'��H�$�i޾�Ϣˊq2��	�b�h;AΝ��>�΋@�Ds�������B���p���5P��7V$��
�Z������a�Hf�������Ό��Hv9�o�uo�t7���>���F��p3�q���+�~��yR��t�P�.	o�2{�x���籌�|�ش��g��~�B݈ڹ]9�dh��mɲVݲ��� �s�j�녝5���k��ܽWX9/���T8`�k*��k��֡�@Z/FƝw&��n���&􇧰�Ȗ�,kF�����9A��.%�]�\��Y�y�������\G.��Y��٢��Q{z��(noJ�B�k^�hU��.�YU��wԒQvT�vn	��o^�F�Yv����o� �	u7M��h/�]�M6^�:�혛��;�s[�����ힰ�A�#zez���[|��M=hM�:��lekstwh0Y�(]f)in�ԣ��둃���u���3�r���,�6J�+)�<�t��]-��ƅ��II��l�N=Nv@oSOS����rv��^�M�.S1^-#'E�9���_�WU�8i��;۽c������R��z���Jå���O.�C��`��|��I}p�Fۚ��x��-q�W�ڰ9���-���<~��5nĨ'WMM\0Ѧ�N^-��-?Iȣݷ]�|z۫	��cE�2CH�
4]�s*��~�ػ7����f��-����Lv�3����.~�}��(tw�-T��G.Q��%��9��G$El�D=Z3�[��+���eV��ij���5.����pN/p�"F>���l�F�v�V3���_Oh��ܨ�����-0�E�̑�D���N�_�)�X�C�s��\Ͷ��-{�U�|�J|-�w^	\����.�0�"d'��'^ow�.0���gK{j�o�0ڝ�|2��9$�4:鼽��J��S��0�����?U���vӫ��@��	%��Wv�����bSil�4鉴4��ٶ{�[�yaDw�_η ��x�kv�N���l_5��t$l`��T�
�ص�X��3�]��B��6hr��o;�u���ĥ,��T����,�Z��nd1T���r]2�F�ʺer�19�ԉ�E��:sn��K����/eQ<��&�WmSKa��Z�[b����!a��&�u-�y朚-\!Y�V�K�76z}\��ݑ�#!X�]kI묻O[�Vy��>�o`}}%��|%l�7u*���N�&�X��r���i��G"s�M7)�s����Ҭ=���NR����
�q�;wT�;|�N;�JZ\6i=b�&�s֭N����'��k���^���.P����|S�e�b�}|ڷnn{+fm��1b�ʮsydcF:������揻�h�w�XM-�G���k�5S"z�;Ϻ[���j�|��=R�C݀�{m���WX/�mks5��[�_�$qvI�����o�u���h�z�E^�������Qɾʹ����ݛ/������i����C:�k�H՛Y�}����&�)=�4�O����b¶j+�fv�µP�K[Ͷu�`~*��
����-x�RiuM�	+�E�õݜU]�;Q��zdRs�r�/$A�C�nt|�0+O�h��rvV��{8�8 �啋��ˆg.U��h!>�v{�[ohv��*E�Ξ�֦z�F��V$��q(b�Ƭ>�
�9ݩ�c��RV�AO�EZ{��^\)��:M��j&fʢ@�錩Q�],1ݺ�z_�c�	�j�W�mMw�$��8��9�5u����Ɲ�L��^g7�}'�e��b�M�5d���j�t�����W�ԜXp�S[ˬ��YXoώ��F(�p�Bs
�r*��~�m�9wR���qyT}�=���Ӊ6z@z{ӓZ��h�1T�*�en8;N���K��p�<x�wi����dv2�3�Ck6���h����	gIƗ# �q�n{�{���9Oknj�@�.�)�9ٹ��8�ؖ���
�;Wug�\�7�(S�:��{HsM,٤�YD&���S��x���=7�t��.7�X�(nT�{3�S\�qM�S]���Z
����>s�Z+/U���ӝwEnE�R$"i��}�̬��.��.CYˢ�s�t����+�z�=ێ}�Wǲ�3s�jw�ARΩ]�Eu*��]��u5��xъu�j:��v�롕�I��ۨPk��X��jT��˷n�V�wB_�����:}�];��{��h��Ӗ�b3J�����U^ٞ	�����$u��1���K��:�(e	->��׈��ăö��Wۏz��z��|��8��ҩԗ��Hi!��97M�ǻ�g9���g׶����T�_[g$�fB	��UQ�K�k���9�]t�܌K���%��:A�&��Ưڹڦ�����X�1 ���zC�+[K.�1��tgP��!�8��7�:����_�F���.�� �e�2�ᵭ�X�t!����:��X�VInk�{j��dEٮB���r�)c؊��\

L����8L��4����gWT�;�,���';���<��ia�<��g$��44:�.ڷ**
�7�t���䤦7s�xS�n���PM懧��{�-���z��mVЛˈ��Q��7�`����s�w����J��3N�=/)t��j}�1�f�ݴ�]֔�����t}�f(Rug{��J�
]�'A���������؛�:�a�%�,�T�3z����RJ�6��,غ���K0ծ^�~��^ao/�ѻ���M�׽���B�L��繞�X��MbO���0U׬R��.�YTV�î��OQn�����{�%�����C��f��oz(dp�St���r�ܴ�Fw���C5�7�fkQ���*{�M�Qщ�K�Q�/��o�D��=�a[�G>�WwS}�twcg��I�KιxׄBt���P�O>�`���`�f-��p�:Ţ�^�k��{�o�8w=��Z5v��$?R�q���45����ʽ�{M����i{-�FV�t�1.�W�U���z�P���	Z�z�";V��}+��/QOq	s7�`O �)y��i)t�r�׾�|�|+���v?C�Ftkw�+�+�m�6�x�ZKk��;׶8����$c���q�9�n��@��uҷ|\�q��q���h�⣯vXlv=m8���q�;���p���ԳhN��7��b!�(^�����������\,(��2��l�ޕm��L�ܹ� 9�Wmi���ͧm(󷂬쭁��/���N �;�]��M��RC��]��m��b.퇰�[h�-2!��2x(�LXf��A�p��y,�:�;� ���.��)���&�;�)���
�e_h�������*�������|_'�7h�Φ�:`�����\�}Vr�lLB���l<����O�8��U���m�҆�A.Aem�{���S��\j�fg%�}4�\P9��������/���]ֽp�&DA�G�+Z�}d���ʹ��� r�
U.��]QoHrW�g�q���v`���bz.���S5y���Ё��
U9M߅J�V0:˼�����i��٦�&��t��nny�ҭ�Ex��6�.;ws��L��hA��mO���l�w��|��R�~��G{s�`S�w}3�+�|'��@���>��Ձ�F>�-�o�-������Ĩ��N�3�z��gٹW Y93-ҭ��o�vt�[��ղ&��^%�|��(<�HU�*6:h���>��|�(Zv�]K�|�GZe�s����j���'M�eea��v����T�F�I*j�b�Y��gt�	���G�ѣN�[�"sVZ؅Y;����v(�H���e(��wţ�������C�7u���<<%g۩t����~��ڔ;��u-P=���7u�M���/f;������`�>���%*��K�`>�*��F^�OniLd�ۂQ�ե�f�M$M=P���6�
AD��^��i��o&�N�f�f�?k
���GhҬL������A�(�w���
�Ȱn�Go�W\N+"����&�)�bEZdn�R�/y:�&���Fq������YbՖ�W�2ƅ��+w꼶��ܟ���`�]&qb�늝Rx��Z��b��KQSC��ኦ� Q��XFc�V7O����M7X�\��G��Z��� 4b�:�p����*�3e�UU�J)K��B��itb:�⃱ۨ�ސ����٢W�0b�M���xAo��6�!���f/�n��cl�X�Y ����:j%c�m�$���,���Ϻ��팛��8��=S!Xq�$|q�^��ڜ��FeH�2�xO�����2��Xn���C�q<C骷9�����Y��wr���=2�y%|Fԩ�9;����?���eߙ�m^k�ɢ͊��m��%���w��b3{'%m�Ѓï����'��vny����C�b�	$a��ɥհƂ�Eu	�fw��{K�if�'cYGɦ��2����ȼ��}�lq�{+g��Cr�[�*�T���#8��W7'q(�J:2Q-kz�0k�X���d�S�^C���R{��mV"_fG�{��=��c2��	-j8�}d6�]�n��juv��J��"���t�S��7sO�-�xy>��8����#j��w�'9=��u�����쬉��^����E��i�'����"�25�����޲�����k~O�/(HZȡ�㌑hnj����-�����Z�0��8f�)N�(x�]ez�hb������׎7�:�gC}�ұVL�^eƻ��hQ��Nŕݘ�q9Lz�Z�J˫��(��P�
B:j����Ɋ�=���y�#4�F���ʴ�oZ˕}\��glh����X�+K��b|��|��*-�{K���,A��������R8ut��eBY�+����܃�1DPJ����FҘ3ˎ!��ʅ����˶� ~>l��wXb���@����\��*xF���n��*N_�ֈ�;��t�q�e�yLp�{�X9$>�5��pɪ*]7���6�E2��T����Wo�j�i��&����6�M5qՊ�	!��*��r�w/\��mzs	�۠Z��C4AV]n�f�Vl�׹�f$�<��^Eݤ���Lb���b��W��/pA�S{��=�V9��|��5��qt���}���W��W����C���x1�ܴ��nbK�17hj:�S���Lv�V)�9���g��(�R1��/T:P�ݗv�B�"�����m��~�kX��>J�,v�O.�vБ�l{/���vg�'y�pV�֮"��V5_j��Ɵ�ՈW(�2>�������>��$��H@��	!I`IO�H@�HB��`IO�BC��IO��$ I?���$�xB��@�$��$ I,	!I��$ I?�	!I�`IO�H@�HB����$����$�H@���
�2�ʲ�b@3��������>������*��HH�@@*Y�v�2��T��6�[���(*(H�������嫜-�fZl�ѭf�l��uWaf �V�m�L���U���]S�e���k2�  �;\F$+\7t�2�Fm�j�d(�m� �	݆�3-c-��k+m��U(�av����խH�6Y�R*�8���F�4b�l���n��Vg�ۡl�5l@m��;�����Vp�v�N���s&l����l�U!k��VڑhPS33cF�[�    D�mJR�6�	�FF�2ba �JU*0       sFLL LFi�#ɀFO��R!L��   sFLL LFi�#ɀF	5H!��j1S�"dɠ�=I��_/��e����[��x��@J?�D��� �Q���`$�$���K�� � �$k�������h2�ͤ��bI D�?Б�@!8�T�2E	Ē Bi��׾�����}����l�I Dce^jW�{���?������XPQT(�:��c1h_ƍ/��k�e=��:i�v�&�[Z��f�/��WV��U��
���wc��ڬ�M��B�5�ޅ���ەuc���X��D]�Ū��\��TCm4��S;�,Y1��3 �z�cD�gi%�`E�ύ��7o3�Ԓ�c��1ۛ�$s.��oV�T�u�i,���EHI҄�;��Q�B�F�Rf��н/tw�&���#xs>�4�I�7n�Ĩ�M[��-]�b��H�5{X/Lxۼ	I��c�I�Y45�`�7v�#%Ă�栣[v�'5,YZ����;w�"��Fw>{�eA��k�����+�L�-|i�HB�>Q�\[L�'&7��MJ�%���
�P�r�)��U�dp쫹���Wzh���+N4��F���b�Z���(�d�	iՉ,���+AcVCD�s#z;��VvM��Tq��.��&(�����;�2y�a�� �U�SJbEh���W���9����
�����*h��l*�-9����wy6�f�#`��X�7B�y�*�S
��m%R���4��n
x���P�
3���k/u����!��hFK���>%��[hɶ�^ҽrQ 0�[�����- ؖ1HKnкx[X�H�fhCo6�VEPNPL.�� U�om�,�s��6`�8X�`[B����"��.�PI�� 5&�k��
R�;v�u���o d�f�cٚ)丮̎�T� ��a_*b���n�S�u�锝��W��g"9��s 
aZ���q���#^J�t�c �ɺ���n��D�䗻l��벵b��ƝT���k�{��b�e�.³�������Z
jj�X4�XTѢ9��U۳��"�D	*}�P0�&��si9��R�lV��	��{VV�!��R�aK�@�b��޽��0//B��S6��k"���0]�Xh���J�M̡�j�<0SF�V��V\S`9r�0�Ʊ�X�f�:+S�U0�7-ꔔ��v-E�.�m�۽t4�tf$��0�/�NdN������͛��*���]7��_�xR�j�b�s3 �&�w�AAV[����W�!5�ZQ�&fݝ����Y��֭]����jĥ��`����}3.eޓE l�ٳkB&R�,ԭ����:(jH1p�o[;��`���Xv���ˢi't�ܽ�&q����Dͨ�S��"�V����T�CL�w+�ӕ��g�[��^�3�[�Y��N����1nn��z�A�:��*"�f��aj�Ҩ�(�īiC��*l7�Ѣ�i����R�0S���R�0�NՁ���-���֩I+�	��.�ᵫ�EE(�9��+ʗd��H�G���x�
$��
Wvw�tw'3K6��c�Q8�Jˍ���U0�K�lS ��ݬ��K�U�>�^P��[E��e	�sTsu˺�M�pof���x�1��S~O��g���L{ߕ�hH�Q�]�Q�g��=挕��oD<�H cD,�z|U*���me�İD�9"v����%�f�U)�cX��Jp����H���V��_]�dEº�,�Ca|f�/�����Jmn����aQ�c��n�V$C�f��E^:�Z/�m=������0��Lɜ�VT�lRm&��oQ��S�;��-��|I��b���ږ��b{)�^���Z����[0B5\�x뼓��+�B�f�Y��ZK:�m�%�58�J�ثy��u��ɢ�R��w`��r*w<+z��{r�d���ܑc�y[��*k�_��h��'��;{uH٩I4����I�]��f� �E"s��>�!�<�)r��֮��mm#��꜕r��rC����N�dh����:�c�uz�I�)�J�� �@IF�5�����*��-�h��[D��G�+V�t���v�tݷ0p갷�^.
ƚ�;9T݊��`�����}g��ujح��;v�p���2S.g��k��1q&�uXN�S1q�1�r�T��>�U��~��:�O���˝z3 �.S���Ec��{Mm�f��G1�`+-���ox�#�݋�)g*'�ܚ�u4��ٷ�Ǔdu��.�@c��k�\�&��K�c��;�M��=o:�e��S��)r&�{rn���;�ze��&��GW�3/ze�}���
q�m[k g.>o�g,�-	W�7򕤈�VՎ�TבLT�=�<���L9\T���'���y��'�n�t9���o,��Nn���	#t�A}����x=ս�urU�����'��7ۚ��
��Pل92oqr	��0��{����6��˷��D[�e9x��"�V���J�$+�;v�����:ÖޗIY�{o�v���� /^wq )qn�U�e{
Yܷow
�)�щ՚� P4Ty��Waz��M⸌=/v��r�MT��zy�w�ޔ����*���9-�	��S��芽�Z��F�X � �62�1.h\�ѐfX�MThD�-�-�mt΋3��9��7�b3���� e2��,�@,���(+����."}�N���,�Xٴ���ͽ�l���e,㘀L>�9�4�)�+dC��,��b��r�n��Dh�3s %�Y���L�%�Te�v�%�z��R���櫎���uM<t�-�omJ;E��΀�J���Q*ݐ��v�t�y�Ih�ҌF%�N��؇h�ѐ���I�e@��
�YJ-!�KȜX��z UJ���D���}8��lPV�mgc�u��8��qN��m�e����B����=�[ۗc�����l��� 6���P�2Z/ �7k{�,mE,�2���ӸK W$׌T�pW��B���Ӟ�����Y]��lWC
�8w	�vV�{�9�t�T�_Y����×��Ǘ?�gE��i��z�E��ז�b�P��o;�'9�x�G�';�����������vOw� '��'��fI!Omv�@����� 	��f{�׶kߍ{����h�$,��%���"e�2��]
�����չqPt��/&e%gBk@CB�Z��rjӔp�-�V��=v�
'J���j�����S~U�mEY[�a���X�^oj{�!���(fL�!)SPcUeњC��ҳ~NWg���[��/>�c!+E��8f���Ӡ��.�z���K�oS��{��z(M�dlV�w_We1U���'w�5q�O�J�p�t~ޔ����MoU[k.��K8��Ry ��K-|w>�k�(�r�3khhb��f�&0��B�s���B_��9e��z�o*Kb[��Pb��ޭ�w���\��sf��7XB�FX4C�qm�2ܗ%�/����Jx�A�w�U�U����U�$DQ���X�3S���HS����7@چ��t"S���q]�C�p�Wy�P��pu���=���u{ƲΙH�T،�6�i��J�U�ʺ ʛ@P��L�,W�Cn�[g��=�ʛƞ��m����n�F�����Ct�SU�A�l"lVJŮ�s:fs#�:OGS^��u�v��۽��0b��l�2�bCd�A�Blq`g��)�c�h+�,�x�r��<����F;�����;HV�6A��k��q��x�I��99�y���f$@��Q�F&lSwW\��,�ǐf��-X���,���n�*:�,U�O
�+���v�Ŭ��Ӷ-�+!�{�53�����T�Z�����-O�X�e�E�33RM�Z��cq]�u��OJ�wcg,���������?d�y6O���f˗M
a=���R���L��M�K��
0�r�N�'h��-��j���5P���Vlap��n �Y��+�u᳒��A����nu��h`h)��$h9�ض)�z�xX{D�'%��d\�c�ҭ���6��U d����6���Vn��݂� 35�{kt�ߴ�5�! �KY��Ms�βu��skV9b�ƥm�-펱��skZ�k�Sc����r��ڽWʐ3��-i�u�����g0�d������v�v�LZ N1֞V���%.��ʬv��"q\U��:�uk�K���P}7���i���ޛ$t����W�9n,˵C<��p9sK;��r����5��Wb�̸�\m]s�j���\]�����AA*?��q�NLD�nX�Ѕ!��)l���!]G���N�Uv�ΥЕ��4xcq�	k)Md�A���Q�bVYǂ��יr���iQ�'�K_?��x̒��W=�y�Cws��p炎\6�a��mc���.�t��D���j�7�sV���7Dfu^wZŧZ���8s��y�wģ�z�oyTcء�Q*L�t��l<+��[���tf襟9o��:�%-{4[�2�;JL%>��;�w�� 6�RpTw�5Ѿ<�DÄ�{����X�M���;�_5�cΗ�=�$�AY�@�.C�Wd���eY��{g<絸ǵ��.ڜ{��i#����Ѯ�ˮ��W5���mX۔�-��%jƗ�Y�L=1�<I^T���D8qQ�� zg��H0�B��]c�b���w~��-�5��B+P�j��iv���y�������xՃ@e4�9x�c��{���:T�RRR!Id�ՋB�I)�H�R�@S0)��@�E�H�,�����#Dg��ݽk/u�U�����o��AhH�3��e�����h���u����V��Ju�\1�^�f����GX�a2P�����w��f'�`aL��qiV.��>�9�Ec4����Fﺹ�r�o�Y�l-���_n�vd��>U53�i�l���r�a""�4b�Io���;:��gCƑ«�)��K�%��9;b�ž�ѹ�=�5'�l�p_\|`u�c�2�y�2:�e��3չ,3�֯��$=t|��|�po�@�e��JZvK�isX�J�jw^=���p�)��zwc[�u�kD�:D0��({���Ȏ��70t�<�������Ѻ]O֠C吭���7]3��w����.��h�%].~���-����!���	o�Ա�^����9:�z�4%XYF�`~�-��5Oe�=�Q�����vݕ܋v�)�s�*/c�F���Յ���W�s�n�m!��]������)e�̪�Z�!SP��B�l�"�2Y��V�Y�c!��V�Y1����Nɶ2��5��+�_c���~��w���k������ܲ ���c���o��fԐ*{����_�>J�;w������ߑ��*��?/L@vk�^�n��=����9ǡ��0W+�r��`�?v*�=�6wZ���}��{ɿFU�#)�z��㢐�
K(@ny���� �]�^�C����y?o�iP�ü/�Cמ�8]�n�"�_��Ӗ=f���Hb���:M�r��/u^$���n�������%ű�E�V�1%$s�[*��k3�ͻ�}4Sף��ų�^P5|1���Bl �{6�oRJyZȧY/XNUm�ڋm���V�X�Y��Q�f�	,�OmT�	�h����IsR��%I:#Ӱ2�_=]�vhWhH#�[���6���:gkb��Y~nc^�Cr��z)�H:�ڸ��&�x���ݜ����%m\+Wxo��-��fK{�6�/:�g������F�Z�eMAK�W�<�3�gS������E��uiq!T^�Mx���y�Ŷ��x�L$.��#���̏s��,w�hVח7�{4��)PK������P��_]��fa��Z(d8����k_И�`�6L���諣�(eG<\]*��7O,r7y�/.x�Q%$���5X���m��Yp�Erk������%�*�<~k:��O8���;pD�z�1aѲ���gfS�M&�Rd�����i�; EX̕���뵤Zǥ߇��7PY���������������~VQ�t�����5u�^'�P�紩�*foU�7(A�j5aT���\�n�&�C8w"�w�:�0����<�|p`���zw&Wq��V^S�(��W�m�۟<+���aN��m���O�2S�����ϐ�.�҉��;�J6��g�,��4=nS:!KҌI0F,���L������#���ļ�i�f�W�j�Բcp�+z�Jφk��� ��8I��"ö�9�ݗ��p����3�����
�Fs�I�q��)�2^��@��{��L8>{��M�S��ɉΓ%!���VL����B�Ɗ�K6#k�LQ+,��,��>���4���(
,E`,X* "�٥A@U"�`��V*���Q@�"�VH,XEREj�H
DUb$D��F,DVH�-0������_=v��(��"�w�s����!c�T���"ʰ�T_�	�^��Gt�sn���U����\s����z��bu-����d�]����J�^}9���� Ev��ץ�=k��+�8T�6A �lTb.,��pY�|��t�K��e]~�����[
J
HQ��?S˴1ޛu	l7��ڂ�!Η��~gs߭0�:�]��EDTօ�T����F�R>k�-��0g�w�ɵ�1~�����Ӵ�yI\e��8��{48NL�%�#�zJ�v��]�]��^H�(�]������$+\/��8x)=�5���pfa��Rv�w8���qSGa�9�^*2y �9��Z;���[B4��j_�g��( ,��k:��� �ν�e�"�/�Q���RqyL..1���q����V�!�~�C<r��)-��82���'I��ùAO[V3|0{�g�,L�����;���x��߭pڕ�wGC��Te s�q@�<'y����+���<�-����&�]-��v���<��3ި'�D�Ϻ��wo�<g�ⴽX�+�8gn`���%�c�Y@�[�ݚ��X0"6��tGX�R��b�=�z]�>���O.-�4s�g���H�Z��񋯌t���Poh�"[d��Ϲ�1<?��|�[�O���]���5�m�I�qή$����Qʋ��n�:�^t�˂�o$b�td�%�>�B�/5Hg7E�c�U.4�V|O_���M��>2���:k{��EY��X��Zkc�؞e%��y���uj�u��H8=\��n���kq��͹�J7��RҊ��J�s.d�i/(G�j�9�}�$YJχӭ�}i.J�UX#1�s�֭�y���U��v'zE6Y0?f�nK��SD��=f���_�#o����4����јJs�#+"�渢�����͑�Ob'�uw~-�ʹ�s�����-�/^�U|�)�ë��W�6��O?g�0܇g̷}�k�2%Wv��)P�)���ٕ7Y���5�wc�Fg�f�v=w��-N���n���.
��U��Ӷ2������^n�ѷPZ�y��5S�![�#�}-<�C�kdӠEn���Þ�m�e��o!mfd(�����=�}~����[~ۊo��`�^Ώ�Z�kt�
����YTt\��Z�<���|�� 䮭$�0b��Sհ�i���C�_��V�_�Wj����0���yf��;�t���D!���!R��������ػ�(��娞ݤpV4�8���Vu50��)�:�[r�S�y� ��\]��� Sտ����̔������w�.Yȳ��U�i���b�����70��Z]1v��h��V��+9�#�p���9i�;{����S�.2� ī���}�2J���JUyR2X!1��&��aKY�����?9D����&a~7�*`�bpZT�1Ah�'���(��s���D�.hac�T��c�M��c��{[�oRs�= �F�Ԧ$��"�� Yj�KJ����;d�B�uE�ɣY(^�� m�վ�K��q[��H;��t΋ݢ��N��V���/wR&I�DT��f�!���U�z���S���,�!ޠ��}��M��p�"%-QU�K�P��.����(��,DV�P��]Jb1YUQ-�J��DDVR��
V-�"���[C-DK�WE!L��V"ƒ�,��Ң2�DD`��auH�aB��X����U�׷�=���k���_�Lг1>w�͙k�5�>Un��}3A����0O��~Nw�yT�����˧��d6dzs�7�F����2we��2HtT��n����;�i(�G���N��K6T4�4�m�f;o+�%��&�������)�x־�j뜲] �VQ����w'��!�����!)֌�u��)XR��خ��в>��r��d,l ���:���.1^�ԟ,�`:�1]���K�>2퇓��A^Xte���s[c��.��u������z+#em���d)�m��Fo3�r�i�������x�N�K�0fh����\
J�C@�;�א�u�������V=�����&�H֕�9�S���e��ȵ�kW��z:�tD����G��Ks���e3�:������UW�w��2S���
c8�~��-��Ӻ2��^�5����Y�p��XzE���%����;\���{W�2��DmN��xfY�hh��W�z���y�#�m꾞M���඄�@;^�U&�|]��2(h�hĔ�/���GODN}�Cĩx4_�rћx8+��H��-�y��̠��js�*s��]L����/B;<b��zL��{���^h�/��׊׊ZV��݊��o�J���b�z�o4B���]���vc��Ͻ�{��S�}so�������v\��_�}�f��,�i{�����WE��2=�`�f��K���%��ے�'��K�X��M#��q����\�{�[�nzN:Z���׽�J!�g���k'a��g����}j��E��C��{���d��5G2ǪQ��ߔ������c�8����P6Ūn%�U� IE��Jc�L��|�5�d�9w�v-Θ�l�����EK_�{���b�/:�@��А�	��r��RB`�IԒil!��o�C�����3[��F^fn�6�[Y�%)Q$$��tj��f	^y�C��fI=�a�_(��@�fH{$�`q����u�S	4��!0$��A�Ha��$;�4xy��䆱DRI�N���H)���L2JHB�w=z��9 �OL	;U$4ɶ���� S$�a�J���I+t�M+o�x��M2������@)�l6�x�ÔHo�IH	ā�Hf���l�2��a�H��@<d�Q!�T���Y�����[$:��'�C��0%$��'P4��L�A��a��T���m%0��
d=$��-���!n�8�g%��d��P�Hm$1����H�fR�Bc�w����㗬���+Ĭ�@ND���}���ήZ_#Ͻ�� |�ضN���Hm����!^�@�d���$-"��ε���0�0��N08�Be���I�&C(置�2�L��=� �Hd3L�� �OM�;�;�C�Ԗ�I�zd2������;�ٯf���m+�Q���E��]��:��4��hב��Q�G��g�m�O3���g���^V���r�2-�8E�^�1%j��{�n��_k�-_E�fk��ʢ1VȾ\��.�ͱӻ�Ud�E��ԙ���ܜM�Y^�kIr�:�<"���)�=b�O���pwq��k34-�!i�"�r���*����G���	��Mp3@ի��8\�K,E��Z舵o��k�T�v�W�� j��r3���Yc��J���;(WM��Vh\]�M�r�.|i�"��B.�1�r/Y5��w.ݷ��+5�9۝*��0"u��k�mv�Y5���SM2�s$L\{��x��۩��?*��op�}��ߧ�-�k��*U��Cg8��A�$&�yyHI���ٲ琢���N��ӷ>rph��uueY�q�i =a�K4F-�1��	vG!"�7}�(��!���;�y��Cl��&��A�jD�����I�ӫ��e1�>�6n3|;>oF�����B�X7RSIJ1T[IKwv��J����ж�i-��I*�����)�6�!I)X,7��>v��g\�c��,Wh_��o7���_*o�r��-|{Mf]y�r��g�[���dB�T�* �y��Q�4���H�6>{����3�{$��X�_	ܲ�x*s�I1���)_�𚽾�Uzl��v���}w[ƣ[gw3n��$fIax�>����g�x�����ߚ�7���ӧ_�]�'3��f�t)x/oX3=:άV�����Kl<���u땇1rC���5ynzP{�s�a}���n����u#~�U���w1�}iN�4���ǃ��^�ᱵ�YEfK�b�iн��4�7��7����x�X~N���,���ժh�p���.�� ��Z>�܏����X�5���'����M�G��v�d�=&����Ǣ��@�^5�xz������(c]I�%v�2gUⱹ�\�i���7��c������QT��ߡ��6�0rW՗��)/t$����+yɗ��y��{R��0K˗HgJ�^9숣=v�_ud�ipOG$�M�f�Z���bF�Zu���!��Gr�o�� h�,=�"�'�ftk��`}������|�R���0���^����r�*}sSj�[R���{w�mj���WlWYγ�q�%�G�:�m;�as��r#��5r\��a{��B�ھG��a�����!�n<ha�Q�%�F�{#��v�33{�ݟc�"v�?�9P��G��?�vns�	ދ�+ڶd�/B/j�֥t��V5��F���k�
�v���;D1��Ti7L%2�t��Ҧ];9Pc�ha)�[{�ޢE�՘�:
c�b!�~����|�5ikt?<��o?s�/Z�'�$�*���2���}��~�ϫw��i��]sr���x��R��B*����e_�C�U������p�1㰝W\�z�/�?�[ܙǥK�a�M�ܽhr�bB�u͗��j�,G�o7��'֪雦:*��������-,�˕�鈍�s�>,�<�V�uL�4�mbW�C#{I��wy�λ�I�۵��b���u�)�����B���Pϕ�����_�
�i�񪐮m��Ć&i����c��_]��v窋?rC��H�P�
�7_W��7rO/hy��w���u��peסy����9�c(�z�������yN��#�M=\={�cN��:�׮�+��L�� �Ko#f�B����A�y���I����fr�u,_��3p��@�ߥV�C&^?(>�b���e����(�øg�fC��ݢVK�O�
sb*k��]��n|�^����1(��ď^����1Uu۬�kG2m+J�n!ŧ\4nl0mE���6�֢!��S�c��IT
Q�5Ճ��+�5�±�$_76���i�[Wuӂw����wa�ܴ��+@��H�u@Ù[�igh4B���2k��>΍��\��'0��'S�4d{U�33�W���(��=���qKj�.˷�sc����璭�/���q<�62�h�DnxCO7wUŎ�:GN��[�{i���jH;��>�r�*ŤU`蜋���&klYZ��M�ɤOxh�(zZT��|���UBh�* ��P��!HTn�~m""q0]�����UVUF���YwV�]J[�ij�Sl��2�����EmJ*�j"�IM4�2�b����5��ghv�v��ճ&��m��Ŷ�7���ByȾ���ϵR����4��X�k��@K�C i�H:rܨN Mn���.׷���q�yA�6���p��Q��]/kJK��/Ԙm�q�ϑ�Ei7sm�2��ؙg�R��;̭�F}�{���_}�y��ݛy����}ĩ�w�+�{�h��a�����#T>��o�Y���N����H�Z�kz�WC�ǝX7�mj��h
Oj����͠گY�D��nj��/.�lm�T�Oh����AI#�y����ϟyՓ����t���3�p;b���4j����� ��u�|��`�-��!y��in����K+����2�q�����؂��-�Hl<;I��u����/q��l?w��`jEN��V0���f���������۳U,}8��Ws�\����Nf��P���$}~�4���(��ܕ��N�ϕ����zV�h�;�M�+y��]5�iy����в���Z.x��Y����y�KuJ/���I�z��B���ա�������Z�O+���?1U?l_�_f�����e�k����pw�`\�u���
뀒!k�w�n_�&5n��I���=��T슰�댊�M��V"��X�J��)�ڭ��1N�VZ�ت��G���ߨ
�<��/ן��s�W1��	�^�yz8Us��6Y�u��[l���)���ɜ��Ϩ��;VRZ#.�gs�<>2���p����z`~N�(H�����ohK���9�41��kWC١�{���Rw��]w�|���e��䷴�����;���}~G�/n��$^އS���}�^,ʚc�sPp��S�2@9-FѨ�X��/55���km�^�GS؁qzhĔ�}�����1u���"��Q6$�Ή9·��Wfη��g��3���N6��ػ���1�}��m���|w�[:y�M-K\+�+���35;�6�i =W�L�x�=d��X-v�[/lu���B����ݟ4|ۊ̫��G�&s딣g���K�گ}zݦ�e���V{.@���7��yM#I�FQ	��}� �k�+�)�"���x[���w��iԔ
f̽N�j�l4��s�]�]"�/V��3{���s��j#���M��m������i5C)W~\�]k�Lk$�XK�:�g%�.�w�Pc�s�Uu�'����W����8'��6��c�]�*� ����Ӫw�)ez�ڨ�Ht��F��[�0�n�����و�R���ݸr-P��tN�ؕ�թIK�gw0D��N_N=��_u���`�̩oL��|�k�����EM[.�!�i�S��|8��/���d�q��ZNe1�OwVۍ���yq���٩@K�kJB��K�ۘ���z�I�ɹ�]wsU���}ڎ�6���	3ld�ʶ�M���@EՇ��qg`��X�*�{���^�ЛZH�����w���A�����\��1�k[C��u���zK�F�*�!�*j��E��.��(�|�C/��Z��Uj%5Q��E]��7U�R]J�"�%4�l-n���SH��)��m5��J�BRRQuH��iD����R��QEB����4P����Tn�WB�E����i(V�R�@UR�.�#MD���H�Z�X�UE]�Wd���*5G�k��O�O�ZCVe�G�ff�����u\t��1��#Y�o�0�Eo�fҶ�]�ġ�cA7dA�C���<r��ܥ�K��ܫO��'�l�5��J���L���a�M�D��´���S�kݢ#[�l����T֙x3wu���,�+N��O);�o�y+w��Wq��f&3��7-H��Y疭�E�����-�V�.~߶���əh$W<�0-u2�+B��8�z�vJg��)nM�V4ƽ����B�(�+A�3W�����(���V����i����Se
��iY����y`L�/0�E�T�+ƻ=ޝ��J�V31��j@���q�_S>}���)�� p!�i��{��!nA��\�����ޮR,W`��y���|Ȩ���ؤ���k$���#u���u�Y=��ڥ�Q9$J+-n~M]�,�s<xvve�D��-���,�ػ�ŧ�D�޹��.����z)v��X��;�!n�\��ĥ�Qz���{��y��OC�+�b���}�j{�3���b�E籝h��������N�x���'X���=F�Y�ޔ�{�=2%��v$��<Z�:�~�puGH÷��U���G)���n�@1H���4�_37�� /�h|����'��Y!��Y�X[�2�Ǽ��tUw\�
����媚�>#&G=)@2��¬��6�Ey����F1��ʷ�7������nW���F�#�sq�h'����Ⱥ�ԝ]�'$��W�W�{�>�3����~g��*�[��?3��u�.��YB��0~v]�[��o�Lآ^7���g�\�N�}~�'��j��Q�OAJb/��d�,�ټ�/��5�8�R�S{�oJ-�y�����~wn��~{�|v3��'a��m����� _�M�� ��6aU7�E�ݨ<7���y��M�9�?Ed�vo���˺k�+�3'����_x�� _�u�qI����)�Ob�����>j]�y�gC�v��e�7&�<�Vюӫ�w ����O�{�p����t睓���xzd�[�f�(��8w���6���	Oe��+�]Xj[��y��P��i^a�f=d��jU�,Af�����5�}���9�f���.�r��*�*���#�$nhouxT��k9e�0{���dC���k��ةg��w4�w�D_Gs+���,t�������Oj�Mx(xa�n�����md�6e����#�m���d�\���<��G�X�����р�S��y���ώQ�G���6�Zx� �V@&z�eB{q/S�+X�#�CK��2�]�#�ٷ�ǯ���Vl$�:-��L����#��\k8c��C�l賜6�|1Qgˡ����x�.P��gN�t��ݹi��&u��DsS��ܔo��ˇ�@��F{v�sf��P��oGa�ժR%d�!%��W b���6���3��xqm�I�ΧE�"�V��M2XJ$��,@�x��J�UmN�4��K6�K,oSo
hE����EP�5B�TԪ�j���SB�[.ҩ�-��hJ�
���)YUB7Wr��5Wt�e4�[j��J��P��R�D���U4���iUP�����0R�)����%QEU��we�TAj�4�H�ݍ��m˻�%�����ե�We�R��.�JjX�St�0��312�0�%�0�L�!�Tm-G������ئ�ѻ���J�c�*�4���6��Ϩ64w ����Vn>�B�q��z,Q�t[�Vk׉��,H'�+(A��"7+dԝ_�M`f��V�ؖi$�`��nԝSttJ>��\O�+���{��W��3�1sN��lOt�bOݜ��ݺ�Z$W��1���~|�7u���$����7��doW���L�~(|m���;C�;&(�z��ת@�VQ�`0<+xf}ZS���_���Y�y�G��ݣ�}�Z��(�<X�UgRf�q���������&���2�2�iS;����n)���os�+�v+��Q.0�������͵"����4%b�� �Yw�,���N�.���9�s������j��K����}�ek�ڼ���f7I��� ����:�o$��z)l|f�k���G^=�im!����ɖ"������S1M�Եt<󺻹��}^k5(��}�SDm��g��8���4,�n�{��t1NE�70�w�y��$Y��N��3�O/Gw�f�����s+���[�ć뽧�ޗǼk��W���_F��F�IAI;�j:/kT��d�A%���x����5�].��S�v\����;�8��Ȟ!r�k��j.�.��]
��L��r��x�{.> c�m��h����ڲ�]<�I!��3�9%���Ak�8�m������������K{b��\~��k�e�v�{�,iJ��o%[��ޤCWWQS}i7Ndr���-��zw֧��r�Q�G3e���J�K�7 E����e��^���!z��We�ظ(�/V��Ŷ��c_v���T6;8�C�}��C��C؅�D�,���	�z1?�"�7M�f��v*َ��U��+�L�<"��S�^�^�
~��R�Z���9����f�'����潺�V!��"W�/,؋�m�֍m�#2�&�ػ�89��<��W3ʳq�=��ɲ��Tkh6��>���&Q�O�]h�BXg u�k�}D}���8`�~wx�j�AvnFX���:a�L%��.oL��+�5�a����rv饇�?1c��M4l��=��ܪc�FaII��3���c0�i�1�a<JMb�znx闪�0��j�I�STwS�a3��v���/P�)���48ꦙ�K�z�4�&���iiH_h���9�j]�����j���]��|_/��k�~5�i�Vv��|�������z�p7�N0t7ݴXU�5���x��ɚR)��J�ţ�,�`�-�)%�^gj��y��ܩC�V����oot&�ŷO;�\��bᔟcl�Xz�+jL{6��ݖ��P��Z-��&U��a�/[��M,M���]�d�����+R���Z�];/4ۡ�H[�#0�f�G��W��P�eݘ�h�ś�OY�O&�2x^SU�����u9��F_W������E70kZ��rǌkn.�۠��1�k*�3P���� ��T��D�5j� w����p��ġ`�wY/ye��g���	�Q RDR �E"h�Q
�$�4M$B� ,j�J.���K�ij�m�QE�)T�UʻA��RYT�wM]�T[uUt�WJ��%[t�E˺)Q���lh�1�1�����Ф�P�*��U�ST�
T�T�3�	u�n�%$�濓�;8�
IM3�c��0��ja�!L�q[0��<�����Py7O��2��YG(�L�N��u�oS�lۧ,8g<�i:i8�j�j��Y�Vh��)�'ySHWk/tw�ʙf�Y�x�ө�U��u6�:�2�i�>U���g�'��*���;��f��5��6Щ���m�x���c�+z�L=	R�f�fwi}5����Pl��^I���c�Mr�[�)ȅ�RUT�Z*�#v:�Δ���2j�#�2B2xd�w4k�-���"��9����e+�|�ǌ2¹��!�Զ�G���]&�S����כ2Él�4��w�i��na�f���j���͡��,�V�b�b�ί7=���H^�S�t��+��v�5�Š����N�����O�γ�;W�Q�e&R���Sħ�w%��7���c��a�ƹ�޼��lyʖÉ�����<�o&�L3�ʃ��K����T�t�p�e�Q˘Ǎ�g|���ΧS	L���&{ZK�S���c*�Ŕn}���������z_]�T���2�v}/�-ZyR&��5e^���\@7�l���=��'��_q}�
=�����2Rx%��Q��]q2�H,6�1^9�:�ٜ���L0��=�n����r��Ԝm�`w�w:���f������y׺�83IǯY�ѝ�Z�^u�g:P�i�1�,b]�m��vٟA@}�
���A�tמs�K�ri���b��a��{|��3Yt�N,|�}��>R�{��w���:nfw����B[/�=W���K�w_xgް�9Kf5G��偦��2��h�I��
�12"�)&R�֨�멌j���2��LuYz��uV�m�fܥ R�^|k�I�����!m��|NyX���ю��;G�
�u�/��x�qGS)�2�y���Xͦ7]e��:f���s�<�x%��ӌ���ff�m��<�U<ݠj��UQ��@�ʹ�-X޺�i�N3�*���n��x�AgY���}�;͇�����
z&x��q���oQ�i/tb�p�<���8g3GP�Il�u0�ߕ�էl4�	�_�lߗ�;�<g�u�%"����k��L𣎙�0��͵��Խys�T��6���j�%'u�R��:�亥y����h�9�2���Z=@-x��k��+�R���N��Ӷ8�Mγ��8�aL8�*X�|p���V��)���+�*�d�\�gSI����:���_s׬�u�e��T�I玻���L$�c����c�K'�#�_.a���y����:�ul�LyF<��yW�(�z�f�[���<p�v�̰�22Ps<���8���U�!�ǯo�{4D�=-���{�N���W*ku2�g��[�3�D�a�,����	��7�u�f
eQ�s��v̳��+=�xRe��k4q�c{�����b��2�%0��3���̛p�Rj�Ǎ��5]�%�NRS*cc���o���0�g�k1�L�3~T�m2�^ܗ����ŏ�5�������	���*���7,�V°��A�����û��*�0Q|��DSF�/[Yzɷ��q��No���GY��l�`���5aõ�L�ۇ)���)�y�o���Q<�[�>!�S/��cX�8aԳ4u�ѧ��ޱ�a�6 �B�����k:�e8�UH��L���;pmS���љB�S|���so���������jC?N.���Q��P"�*�r�g_���� os��C/*s�m8��^�!�I�q�є��c����a�ƦS.������^+p�a�4����Nnܙf�V��I�q7~Y�I�ԬP,�[�;��y���+�0�<L�������7���0ɿ(�c�v�8��(�>f�^QT�Y�A����
�¼)ez��K��1f�M�Gn�y,�a�>\Z�K��7�n�*9�p�)9Q[�z��Ħ���JR�ss�8��b�-�Kٺ^��J�[z���c#x��q�ެŖ�	l��U������On�lC=���&U��y[#9��Qt:����ys��E��y��$���c��r�9t1s�ܺs�9��pufrUս����Q��n�M y ��8d�[yʏ�I'WGA�h�k3:�A$\%q�Q�5}�K��k�]�[}mim�]δa4��/5�7��Q A�/@�R�����jmh �3sq��Ӻ �Q��(��s��3�wٺ�U��Qb2�����R�AR4�X�MUR�m�KT�5H�Ed�U
E)��� �X�tz����v�Y�|�)XYF�`t��vo�]���ݐ��̹6f�f��Tˤ�)�Hs\��f����NyF�{��1���r��a;t��嗺�7Um�șJv�:�3�L�yre��,O�J�{|ɴXqS)6̦��s�ώ���m�C,|7��6�!�����q�Jv��x;�{�`V(��կ��o+ԇ��/��uT�c�W�+m����Ŷ ��s>'L����*NV�g0�|f3Xa�������p�2�[8���o.Oǩ�,� kW[�k���se�Y�T��fп3ya�n�9ZE���nZjC�cF���4(P�X>SU�O��'�՜NU���=N�G+5���:βR��,x�8����Ѿ׈u�e0߻�Ǒ^�ؤǑ[lL�k��z��[�&bR���Vh�l>??�z}[���hp����Gn��Q5���c�ͳ��򥦘e�o���2"���Y��S9���o|���i�P��n�I��g\��B���4�a��\KL&��l�m��7ƶ�N^2��f�i�5���Q+U6��r��꯶k�M��Q��W[����Q�d;c ��mm��M�R����kC��3;��v��7��������a{���u�2���a&D����f\7�5ڛ�x� [�Vy���Sz�y;s�Q�q�_J�����B�f�F��4݆�9�A{̴��1�9��mgz��9KF�=���p�_�ofos��-hos��TM�ͫ�l�����:a�V貫�;Vþ�s~�uU��Q�Ů{t��<�Deo���hfՅ<�y�-EW������������PS�+����{ۋ�`j��)���ՠ��f��Ɲ�m*!V YA���;��'�R��S�����Z�wҮ�B�vYp��\��a�q!��o��<@��Mw��%X'�i<�yEa�5�t;)ƻ ؊�؄�0Nѫd��"�HIj��b�Yl�s�����-���1��z�q�W�*I�s�#~���F��zz��I�ڿ?u�]�)�Ѯ�4�̱+y��0������9s����'��
����Ў�ۃ:{Vl�R�2pXf�sT�Q8�GU�#T@���͜��]��xq��w"(T�LC'w����-~�ƺ��.M���巰��ۀ[�D[���f�A���Ŝ�$�4�G���N^�1%j9�"�W~_�|.}،s�n��w����1LP�"'s*z��:��;��M-xM1�ӦU�ٵr�\�gj�-�/x_SE.�%ئ�Ҽ��#�|zYz=�K�q���E��¬�������e��ۻ�u�_�<��%+�(�K�v|v�ewb���Ul˯eƲ����-Q�Y�����^|��A4�Վ�;+��\UF�Q1�R�}�Um)������M@���x.Yk��{�lQs���Ay)ꏶ�1ޮ##������ǀh>��5�ʸA.�bT5��d��őA�{5k�]̻�o��{f�ZU�P`�qK؊�*��L?c�]ԓr<7����cE��Hdl@o���K�
��ؔ����u�s�k] Z�a�T K�N��Sם��N����·	9��|�"�^�"��X���ک�L�Q/:4�A�fZ4le=�i��>���Uĸf
<���O8�f[���Z}��'9�T#�՗�`)��fP E� 4�sj(D!U�m� a�V�
�Twcj�9K�M��?V��r,&j��HR��ALX*�QAUQ"*�5�	M#���*�eR����AIL����l��u�j��s�c]�KŠ���Y1U��-Q��Ɨtί��]&���uw��k�X=_��V�`�p��nJ҆�����7�Kr��+����5A�M4���+W&��H
��t��ez�Ȓx��3C1|J��LQ���r�!ϏN��~k6��ve�Bh]9�ӕ����4}�U�ڼ�]�\e�m���n��޽w\�'����J�0w���{!����kG��9�33E�9���)a��l|��C�k�X�֞��up��%��g�fk�c�H�u�9�S�­A�Zo_��y�u��XmAd{*aԪq8�������oCמrA��hw�ݧ;�_��ݟ��u�Z��~�A0/,�R��ޣg��}�괗x� 2JL�.P��yZ��QBV���)��l���稳�G�{s��B�M~X��굜��k�
W[2�G��/7»�����1��ՊI��<8fwA3�Ө�^U��g��W��R���^r��~kw��;2�������t�k��+�@Gh��Gԧ���E$3���1��L0�y)}e{��9���D�f�S6T�j�����/'p�&��t����E1��HV{��o�=���r�ծAe�z�'�B�u�����CK�����V�A��N���s�˭��}�ճ�w1���W��Q��@����Y"s���fT�!W�Y����j�,<�ʲi�}�ʇ9�\���|p��=�C��gk�ak�<���E�u��N4;ћ����8��K�k�f�!�M=�5;Ouo0Lv���V��6��Q�(!v�政�x���X��xxl�;5�=7{�"���T�yd^������Z{1K�b���
�����Z@p�#aם�6��Y�as���"g>숭�j��k_��f` ӵe]]���s���?xl.��KGc��2ã�ޯ�'�*�.��] @�\���4g�l�f�K��o�+�*0G�im^Q�,nZ�v.9���S�c{I�}���L�9��9v���8tfwu�/pN�R�uz�z1��ݾ�Ou.U�5&�^�x��R�x���@�)֓f��'UG�����IQ�K�ET��M6ђ�#�h�ވ��=3��Q#�ʧ^wjM樗����Z:�e@e�0m���'�]��)��u�,��凶��nB7n���ܒ��f�w��'}���N\O4vl↭h�n��^��	]��{uw�'�|Z�'�`���V>���1�1��t/vw���}������'�E4��+p���H�?�I$�'���S��Iz�h��V�(.ʔ�nQy�`�/�(�B��7l��I KE4�C� ?sA�9ꤘI]����� !?f��;I�����{�v�T���߮��5�����@Cr���p�ٽc��w��>0H��z���vc}�I$	��y��.�|�s��(5�@ �� �� '�!��"¤������a��}a����Ib�����}��}�C��t�G��$�H��ƿ�����TY%��,	���hh�F���&dy'�
ՠ�
���"�}D����}�}����?��*I G�z���`�nk��$�@���t*�w$��ϵm�WM��~I���G�$�H�h�HW���O�������$�~Y�=�4>�:{��'��������~���2��h2�$���9Q�O��a�������2]C��S��(4I�}�O��ϲ}��Rt���>a�}|=���>���H���<��"(~��z����,��jDDb��C�I$�'�~��	�s��}
��1��+���N���0?3^넀��>�1��(|?��{��#3Rd؀}G�4:t���IQ?Ru.Mj����T?=�3�T?���L�$�������x��섒H�>��#�OxbO�_�?�����:}P��t>�,��?w�z�G����>p>�_�}=?�? ��>�����C�?��$�@�a�1���E�HO�����I$	��0������d�g}���8Oi<=�/�~�ɜ�̑�?d�с���ߪ�ߢ��������~��������|�c홄�H�>%�|����`ߵ|����I��|G�����k��2�P~�d��d '�ē��?_� }O�~~�_��@ ��I�i=�=h>_*&�9I�&wu>��I�"�~�'���$;�4�]��BB��>�