BZh91AY&SY�)��_�`q���#� ����b2��                 �                              �+@>�,�@7�
RF@��
     � ��  �` L  (  *��
 �  }    �
 ]��BR*�D�J��R �J���"PR�RTE
��J"�
��D��T�B �E%!$��H��|�I( �)G0*��R")���LW�e�����'�� ���yJ����vv[<ځu��9ޢ���
r3�i�   	Ϥ��>�uB��k�>�@<n�z��<���=�9S� L� %������O�:�v 8�@�   q�RJ}E�	H��H��ݎ���>{� }�όk����� �}��U}@� ����=����=�=������R�C�}�=��:�   �}I ���`	�o� G}�� w؎��{�� �>� �>����{���|@����}�  �P>��>�Q/��"�"�(�A+,
Ux m����	w�G����v 	���/o`wq>��y�*���{��;�+�ly ���  �{����۟))!��� ����w�P�x:P�bv�X m�'1�ö�w�UC��� ����w`	���P�  ٣|����A�!R���%U$���| >��w�T7g�<�e� �����=�y�{��/`y�:31�` ��EQ�NF��w`@   �� 0w�;� 'w�[�������
�9� ���"]���<{ �gG�����9   T�䔔= |�T�EII"(Q�mI(x ���{ {�+�w`�� 9�R�c��v	t� ���� ������W���(  _[ovH��� ��@sި�W���b��g�{� :=� ={ޥJ�@��9��vs���%UE )$� ������4�&�ɤ���	��H`E?�RT� �    OѪD�RP&  F  � 4�*$ԅ  4     �I���@     ޥG���UJ���h���I�ڦ����������w�Ib�-�D��?/�~z��|?>}>o��IH�z���@�BH�$H��d��<�D����>�K?��g�O���?��~O�O������?���$�$�d���Ud� $������@��ĒH�C��?��_��?��ȏ-����*C�u��9Dz�Pr�:�Ql�9al�9b`HiF@D�Q �Q�&�!'��ʜ�ʜ�ʜ���%T�NX�X�NX�NX哖9g��O9c�9d�9NX�X咬哖9d�X�NT�S�9S�NYV9c�9c�9c�9c�9c���T�OV9NT��NT���$�z�S�9NX�X�NX�NX�)�r�)�r�)ʓ�9NY=^SŎY',��9NY'*r��ʖ�yd����',NY',���br�9d��NY'*NS��<*��NS��r��NS�',�\�NY'*NS�I�r�)�s�,��r�9Rz�,���9NS��OVr�)ʓ�9d��NRr�9g����r�9Rr�9d��)�G)ꜧ)��*r��NX�U��I��,r�,r��*U�r���$�r��)�*�)��)�r��)�r�,���<Y',r��,r�)ʜ��*�)��*r��*r��ʞ[+����'*r�,r�,�d�9cՓ�U9c�9S��9S��S��c��c�9c��X�NX�Z��',r�,r�,r�*r�*r�/,�c�9c�9S�9d�Y9S��NY9SՎX�S�9c��r�R����r�,r�)ʜ�*r�Y9O9c��9NT�9S�u��V9NY',r���$�X劳�'*r�,r�������ʜ�,咪r�,r�,r�,r�*r�/���,z�ʜ���ʜ�NS���V9S��NX�NS�NX�Nx�9S�=T�T�NX�Y9c�N�,r�*r�,r�)��,r���,z�ʜ���ʜ����%W,r�,r�,r�)���<������,����9Rr���NY'�r�,r�,r�,r�,咬r�,��9NT�9c�9j��)ʜ�)��9\����,r�)��,�������)ʓ�9br���xU�r��9d���r�9d�g,��9NS�I�r�9Rr�U9d�*NT���$�9NS��r�Y�$�9NX�r�9c�I�$�9c�I�r��r�媜�NY',r�9br�����<X�Y',r�)�r�,r����,r��*r��ʫ')ʜ�)�r��r��%W)��,r�,��9d���X�r��)�r���[)�r��,r�,r���V9NS��9c��r�,r��r��ꜱ��NY9Nx�9NT�c�9NT�X�X�NUY9c�9c�9S�9NX�NX�z���c�9S�9S�9c�9NY9|T�NSՎX�NS�9c�O-��9SՎX�T�S�9g���X�NS�9S�I��,�S�9���c�=T�9S��X圪�*r��������\�ʜ��')ʜ�)��O-���V9S�9S�9d�r�)�U9c�I��NX�S�NT�,����r�9d��NT�W��9d����*r�9c�9c�9Nw�T����ʜ����ʕc�9c�9c�9NX厊r�)��,r��)�*���*r��9c�9S��yNX�X�X�Y',�')ʜ���,r�)���NX�VI���r���'��r�=Y')9Rr�,tS�9c��9c�9c�9j�,r����,r�,r�����r��,��=�^SŎS��X�r��rǫ���)�r�Y��ꜩ�r�,r�,x���r�,r�/���ʞ+�9OT�NX�NX媜�ʜ�*r����NT��r�)ꜩ�r�,r�*x���z����r�,���r�*z��',r�*r�,sגr�*r�*r�*r�*r�,�e�c�NT�9NX�r��S��I�$�NT�9d�����r�,r�����S��S�9NUW)��,r�,r�)ʕyc�'*r�,r�l�rǋ'*�ʜ�ʜ���ʜ��V9c�9c�9c�9c��*�,r�*r�*r�,���<X�NX�NX�N_9S�=Y9c�9S�9R�/,r�,��ʜ�ʜ�r��sבʞ,r�,r�9NX�O�9SՎY9c�9S�9g���r����NT�X�U����ʜ���r��r��Փ��d���$�NS��Y���)ʜ�ʜ�*r��NYʫ$��d�9OV9d��9d�g,x�,r��,r�,r���NX�T��9NS�'*r�VIʓ����$�r����x�,���9NY',r��:Ke9d��)�$�Iʓ�9NX�O-��I�z�NY')�r���$�W��NY',r��)�r��OI�r��9c���y$�9d��9d����,�\�NX�9c�er�*OU')�T�9d��)�$�9c��x�,���r�9Rr���$�z�ʓ��I�$�Kl��,r�,��9c��9d�9c�I�$�r���$�r�X�r��r��NY'=y$�x�NS��r��NSŜ�NY'�$�r��9Rrʱ�r��9c�',��I�',�d��NS�'*NX�`U5,D��b�DFI�ybr�9br��9d��*u��I�NQ�G��#�eI$�d�:�A��$I�I�ʒI�C�=XG,NPr�'[*I',����!�Rl��Q��9Hx�9bI9dl�Y!���#��d��W����#��_W������������_�~�%�y�LoN����E����%ܜ|��s�]��Y��P���n��Ew�z��C ��%M�x��{�"��4FňА�١nqˋV[�]����U�%oݤA���U�#�vsWj0�L���}���M`�@�n6Ƥ�8e͈�J��-�j�f��5����n&��KP�ʦk�S1>�:��,}ӵ&��}�`
����/8r�PΝ8����r�ս�����-�������>��R"�0�Ѱp�!�Z��#�Я�+K��$�[��遮ё9�{�S6�*N#:gi҈�ک�[Np�6g1q����gdZ��n��^��sL����j+�oF!�w"#q.�[��sN�����y '5F��]��Ϧk�v C���ܠ�V6��v+1v�5���P] >ܗrk���)wY\f�u��*3�r�!}��oz.�w��{Q�{���Y̷{�9ٓ���u�ˆv���- %]�57�^{�,ټ �~�ُ��t/s�[	rDJ�����M�[�+��2�'mܝp��U{�5f��������L̬�C���	� ���\���Gx��9N�o6e�;���Αs�V��v�L��q,�5r��4��n�����1\\@�1�G%�ظkDmMQ�cǼ�`����=����|6� �Nꛮ���۷i�;&dW����;Omթ���94^5)��e�w!vGm���7J}����d��V�o�pE-���zʻ�g;�`�����L�. �7��t<nIv耵Ű�/s�W���q�c�h��{nr�nu�2�k��&Z�p��`7����r�:���� 뜱Y4��]�9<�C������T��Yf��Z����Q��ٚ.>|��=Eِ��&���w�ŗ��I�]��5d����(�L�ȨcŽt���d��+9v��\��t�n����)�i٠X��Nb���L���-J�c�L���٤toH✝���
��帄�V�󎜂?���yaٷ��wdن3ݬ��f�9��/VK;�vzLz�x��r� �Y�%2�O�ZA3sqB7��5����0r��h�VE���:}n�u M��e���{��&=*Z2����ט��h�2�e��<�B���b�ɑ����?=͆7����7��UP�s�*4��Ձ�hXN0O�.�cmp��;���l�J���cw{HA��������HS�2Ԇ��������}�c�qQ� N����ۼ�S2��.Aa�u�#xۡL�_�^N����XHD��{k#��������y���	����Q��5oi�ض��\,��,�1T;*�����N���]�9j�*vlB� %�m:6����r˩�X�{粃il��G�� ��I#�׵%�:��Cץ�iY$�Ė9nι�"3r�8>�j������]q���v����m�#�m%����[>���	�@!j�k�wRpB�U�8np�E�� ��Is7�=�ˬ[ϋ�Im9�g��nq�xaks�^җl�x��;����
�)w�E]צ�#�0c��g$��sI�<Ի�1���p��(����vK���sv'��˂5�ݳ\4䃴t�G�.ӏN[���-=���z��������ѕ��G�Md��w�g �G/���6�bN^$m�n��H��zv*���{Z;�m[��ػ�i�5L嚳q�G��U_shW�ǤCjz@h��J�E�\�l:_l`j�ŉ�Y}�=� Rٗ��&�/���Mdn���[�^��pZ�Y��0ONj���ۆ�������W#��!����A3S�	�T��9�`�՗Y��)�5#�;I7fn> �&1gF��շ���=U
�Z�3�?t��ﻚ�V��弁vޏGB9�9̸t�#�2M5,e����GN�}7f��@n<8��/����!�܀r3���$7-!gH��g
�v�X6�A���\�������`�B������ot�N�o��J���4�M�%�휶M�kH�9;�.��n��F�T�d��G~Sf���
EL��-'^vn��W�=hYzU�^q�q�f���N�7�w��k��#�ߏeX���$�q��sBպ�ܴǹFx�9�|r��:��AӅ7�^��ȹ��\�N�냧r�^�:�¤��΍os��2���r�=:��Ô&q�
���4�r���`+s��n3���nu��`�|����1vƸ�2uwq��wz��w��}u::T������3�wژ�sD�#����$G�h��^�"�wqy��[���^\��"��Wã]:V���7x�p-�Y�J��ħ�[�<�rLp�O��9j��盵a�4Gt��/ �M���U189��tB6�gv�H�& "�9�����TwwYr�z	'1y�ު�oy!��r�E�n�0���a��4h�r�Y1�2��F���{����ܸk.=i|�۳Ä�b���N�ċ�Oal�#�^�I��Np`!�vI�f�Ewr�1�ە)Y��l�rr��	�
yɘ�gU��k�W�#e�wn)μ�bP�B�6y_,-�ӔD���y��y�_q̳�Ly��NF�Nx��ֲC�E# g�x̎e:��r��M���ޤ`�!��w���t^{��V妲�r[�v@���*X�㈔sR:;���kX[�0C�4Dr�z�����h�2w&±)�S�$�p�p�uo��w��F;e;�i'�	s�����Ƿ;�c�����4C�d|�d%�L9A]�ۡ�x�0>�q��^�Y�(7�}#�+':�\0���re`C6q'gS�;K�@��m��n��]l)iS�^�������o#4�ovq��¦a��T>35c�N�JWC��H�n��{���B<��Ȯot<�N�:��ᮼy�2�~��ٗ.��wE����hc��p��S8����p����9v�QvHl7�|r���ģ2��}��v'B��˱�&i�M6��ˬ��n��'	�ܭ ����O�Q{�娎Ӊ$3i{��C�М���-%Z�U]��f$r k;�]a��F�n�n=�$��8��ӻ�f�t�R^K��L����]ظ҅������5�;9"�f��Kq"�A˼Oۺ�����d���v�7uw3��c�h=��Ô`�hx���U�V�Ul�y���8*Y��.W^�ob�{!��y��95�Ι�v˻��vI5Ю'���h�ܔ��QN�\��/�Ӆ%�aMN�l�}�pR����껤:���h���֕���ҭ�R�|j���T�+`"�mɃa������v��F��=t�S��I��ͩ,��)O�n;��Cɻ�bټs�v�9���KK<��[ۨr<�����7_ڪ�яov�r.�d�3r����gK����#��}���ṩi=Z���[��z:�e_0�R�ސ��	ǌ<�67�Kj��4�uݏz�p�Ĳs�9#���F�|�;L9�v˱,�i)�+�f	��f��G����^+��;�\�2|�7sv�3{;P惻Pp}8kw[w{�v]���4k�޺r)���bZ�A�{�m� ���\�/��wv��ҙ����U���wG����I�z��9�� Z׎�}��K�����:����t�|Dɼ���k�,aGmӏ`���S��³o=�7�*��N��W��	\����7���0I���^�Ύ7�vT;�L4$�vtTu�ܶ�p��ݳ]�Uz	.�L�w`Ҟ]bq���
ѬԷn�@=�'e�k滐��Ⱥ��-374lܫr5��xٻ�ֆu#e�����ev�2l��찬�*ǗD���n�rz����n�Qn�U�"��eB��sb��ۉh��m��6��+�F�v�#V�y�Ӹ�[�ZT�{��t�M7t\��v���c�r7Q�������ԯu��3n􉑚P�F�nMɬ�u�':���\)�^�#����v��cX�|ծ��v��/.�0����5㻦��q�X,���8�]};A�;C��i�9{-��d���gM�[M�u�N ��Xov�p)�����2��`b��Cb-�2��������y���V-6^�����y�$��5��
�z�5eYX�^��ܔIH<�ٛA����5D�tt�	�Z���*����i�d��.�ݍr2t9��q�Nj4�u��re�v��0���`�3�����7�]=�˱�W��{����lE<GB:�bvMd���t���n7��V�9�8��#˦�V���^\K�ˡ��肽���A���ANO;#�2�Y�Ld���v�c�{ܜ�Hk��W�<��`�S��]��׀t�\�<m9n����p�]x!��C�j�2�3.����rכ4wc]����n���]�9>�7 ���wl����qH�;�񥇯�W�e�,ٹ�7n�/eof�G|����z�6�w~�\��Z�@{s��x�n��\�LԴh'�ƯN�%���aNtI�ڒ9ۤ`d�8��|���>�Eg;��Wt��ohth�r>���L���*���[:�D��.i���͖ertfJ�#�N4�E\O��qsl2jY5`�6eW�{�����8�y�nv�O�w����h�pk�|��ʄ07&��u�W��P�����7�b��t�7�F�g@�\z�m7J=�ɩs����!8:�4},�F��g$$7LS�!�uY��♤�[fW��4��Y�܃7��C�#/&	a�U�K�:[`���7͆�/\���60�2Ǔ�������n#�%�=�ü?1�JtL���Q>��кP�J�� �FB�$T$����K' ��t�|��I����WN�wvĒ|I%���N��c�ȥ"i�5�
��4�ϊ��$�Ie��
L%����f�_H4�'Lls�X�R��O�ɻ&�{Dih�0�it����Y4�G?Y�OC���g<���8�������)C�g{�'<h]����u����`m.I%���C��,�)���a<I&�D�a��f��&���D;Gz�ݤ���Y)���x��y"��Z���Q#}�敞�}�K=�v�o��M����QԼ�D �kQK&�����d�N��E/��aݍ��}���M1�ˤ��`�Q:J%�	f`��&�t�M%�Q$��)���V��_i8�n�gP�z{I|��}����d�,�'K���a�wOL��'��Q>%�e�(�V	GQ�� ���l�Mga,�%Di<K'I$��PeK��\���7����f�WBU/
l���f�I�I(����$�K'}��ԙ�������\v͐�'���%����x�rWQ:W�?t�<����}���~+N���N�Ϗ� $�(�M"d�8�O�/�������C��Vˁ  ~+I�0??��0��BI(�
��(`4�gKd�|wzK'IFf�T��8:�	�Q>%�I��Z�;��|M'��N�I�<I'I4�^���O��I$�K%	���%�%[��<��Q$�OH�a���xYL d�� �����O��$`�0�W{>.�}�0�t���N%�0z��xIR�U��:����&ޏI�I?�>�'J����G�/�=Eq|_����������m��&����OB�G�o��0N��3�^ӥ�:+�iW�K7�
윙���0"t�O����a�B��4|N����I��Lwޔ���XL'�qxF�I�}��Je�V�4��p(���:��P��a61��+M������է�0<�5��=�t��y�I�y�N�JD���{�y���<wǭ�:O��.���|L���u$
n.��.�����'T76�����N���x�l�t�%I���n�3����D�<WO���+H�������^/s�{�^���8?����u������3=�
��|���} >��6 >�����ҡ<J$��|fHt��x�_���i�L� �Ҕ�n���I%�	d�I�.~���x�.���O���nK�:H���V�O���#Q,���,)t�N�%��+��J!��=�ݨ�u]Lc}���+J�R�X�[��[	%	$�'J�ꓭK�أ��T(���'�]J|��eRpa+D����I�Q,��x	���y/�EC��}����}/��J� `p|��ނ}��pt�K���3��E:��O��}݃�_�
�1�V�|WȂO�'�Փ�=� ��Y:M'Ǵ�ޅzq��I�`p�S��f)8=�q��Μ��q�&���'��������K���On�/HFHN�3A佛�X�I>%�v`o�w�Xl`y��tu�>�~��0�}�s���(iX=��v%��z�`7����������Y$�W�V��9�۽'�u�t���I
�Ě��yjm���Q�3c��BI�����]�?Id�����w���$'�D�L!Dv�7�%>��?��t�I�!-�y/���|��>�%p�Q'Kd�4�L%E���dD�� ����Mc~%S�f��8%�h�(�I$����s���1`y���~MRi�I!X'��,�I'���*��t��2I:H�3iN�#$f�N����2t�J%��x���]�Μ\��=�B��L'O"<v?H�>+�ذj+ĲY$�*�'4�w��Q�������޼-ߐ���~�h���~;��!lB�'���KIT�d�l%���I%�BԄ�H��!* $R!%d$
�!��
+ �AH+H��� �@�����$�Y )!�� �D�,�ؑ$��'� J� HH,$�T! �
E��P � R �B�$�-���[ZDIl!T VBH	 �P	 "� � �R��	h��H�<�HKb%��$<�G�X�Ih�lI"�B(@� ��8�`)�L��:�^zo_ΰ�!�.��zȤ<=�XY�hd&j�᫶��Bx欹[�,���X 	�&2VJf��Ň[�5���!:�Ր���j#�l��E�@�3��BNygI�\)�!]��n&Y�)ۉm:�����dM�����s@}k.��Hzç�o�$��u�zv��H�ӏ݄�m;���=ІuK�n��ͷlR>ۭ�>zsD�u5j`�N�ޙq��*.C4��p��o5�'Fw�s(O��;�#�y�a'<�m�Rm�Rx����@5�y�`I�I{����7O'wi q�����H�<t��$�����@@�@ Ϩ*���A�Y���HtrX0ѱE�
A� a�dzT�`��k��H�Hf�q�f�Y`́&�r(�D�E���+�bQ�"�r��ڍ��c�J`��/N�	���]�{;�=@�5C���xj��^�a�9��P��v����	P�L�7��YM�v��vI�:�0�YB�ڲO7N�Ӓj����A&#�	3��W@���8�4������z�oW�n�岰R��b��x�������5��_����D��������$!???W�/���?������"!?����������G�?(?��~�~b=^�UM+�d81����X@�U�@����}����{�*�K7�y�E7 9t	��s��0��6�#u}�F{y%��}^-�,����u�y�S�³>�G�o��{�}����On'�}r/L�r���i'=/&9�>��<�x�kѳ��g�#3VaX�^�UUt��G�/�p�r��ޝ�OJ=�.�����W��m@^����8�Q#��d���,W�s@EfJ8R,w����������G} >5}���L�@ܼi�g#0�͸̘�Mc/���~���7�^���Q�z��x��qpb{�!ڗV��\�7������On�{�����LJ��}�w�'�����s��,7}܇k����WF+բ��`�4�����ߪp/1嚗�ȖvP�e��gλU��=��'o��r��:fl�F�:���ܤqg��{Wd�9K���"�ch��x�5}|�3�������7(W��y�sG�b�WV�]ܟ�[\��ۑ�x0z�.�dyWֻ��O������3?_o���������񕙙���Y����홞�>ٙ����fg���϶ffs33>�������ffg333陙���Ϧfg���϶effff|fg�����}4fg333�+3333>2�333?�3333?�333>������ffg�3<fffg�Ffffg�3�ffg�33����ffg�Fffff|efffg�3=ffg333陙�333�3333>2�33>���̬�_l���y�����dЉ�z]~�>��;������{(ԳN,��G��qݨ��,�>��gu�{���Տ>��v�>��^��=_a�I��7{�~n.ON,ϳ�{����E���=7v����V��w����Wz��� N܄�����o\N.*,���'��L�mOP�ո�t� �
ݨB0y������^�����4/q+�����ø_�OC����ᶠ�X,@�\�?e0�^��!�ft�����}�b9��GR�C�V;�}�;�[Ở��v��t~�{�������U}7JX�h�Y��{�g��k��u����E���6�s�o'��� �<^�"�Wܹ����S�~�yi�����;��Y(zg�v�f�����x�8������a�O4�4��v��;�)�*����}��%M79�@�8,�oh{x��ާ�;�"�;��ϳ�6
�޲x-�	�6��4�[��B�9�/� ��0�݀�P��C<�܁�<ׯjd��)=#tu7��7}�'7d:�l�2[y�Oh���zb��Y�~�o��3�3Ffffff����������񕙙����񙙙�lό���϶fz���϶fz���϶fz�����fx����ffs33�ffg�33�ffg�3<fffg�Ffffff����ffh�fffff����������϶fz�������̬���ύ������������fg�����h����ό�������Y���L��fg�����h���϶fz��<ff��];���|�>�����w��H��S��j,L=�4=x�����?e���gM�v�f�S&	�}�(���@��B��f����I3��;���[��G�xO3�.@=����y��vٽ���y�����G��dъ�{=f���F�]�Z�����w��xA�,�q��Q�v�c�^��zDG�,�}�����|E����t���&�a�Þ�}�>4k�s���I�7����4�q�\��ݏ��QI
z��a���T��1 ���H�g��߈c%KV��_t�·�}455�4{ܽ��.kރހ7�Vm�+��WAkܲ�w�^�A�0%���c�3(a*�0z+E`�G{̓�S޹4��|��X����[�w�η�y;,W[�u(g�׾\�^>���w�>���\'���$�����ٸӛ!�S�N\O��<�aWr>5ia�з��~���흖���"y���}��|��� �Q��D�8y/yv�&�ȉ��eYk���\�}�|���<��~�=�3���s��ɒEE|z�|~>3���333홙�333�Y����333334ffffg�Vfffff�������333?�33333Ffffg�3�ffg�33�������Y������ffz����fg�����fg�����fVfffgƊ�����|g���Ϧfg33�fff~3+3333�Ffff}�3�ffs33>���333?333334ffff~3<Vffs3>3�Y�������<x���7�|��6��������3�uX�f�V^��	oo���3�䏦랼0�e�܍���}�6�Խ3��C�y��rv���<��7Fx�q�Y:{�u�p����8�Գ<�h�wr��R�s8G-���]�/{]�pc�/T}�l�^6sޛ��<����{z)#��:�pe���2J���n|��?�&Ѿ����|e�XP�F�0�=�#|���^��$l�Y����#$�|��I�_3�
"7����]qG�^����i�~�������D���{�G�QI�sA#~�c��W��ݹ�D�cA� +7o����9�<�ܻ��������6�7{s�c����zQ<��w�S���>ٞ���Qe�.�1�=��r$��%ϓV��Sox���x���d�YG�S�V����`�4ُ���,�b��2��P�Ԍ���=��e�HQ�+0�+��i� j/зq���zP�<�[]�5f}����0gvm����0���$�� ��>o&�Ψ�A�컾��л�5J�0��u��ǯ���>9��c'2���'�*�:��ŭ�����lhlllfg�33����L��ffg333陞3333�Y����������Y����������Y�������������fg�Vffff|efff}339�������ffg�33����L��ffz����fg�����h�����fx�ffg�활�������̬��������϶fz���ffg�33�ffg�2�333>4fffg�3=ffz����zљ�<&�Ʀ��=bT��>��\�YJ"كNd�K�|�P���ˏE�POc$B�i���:uv��8��l��l�o�&�=F���ۛ�O/��sxU������?Y�W�"{��s��z<�d��vy�9;�=ގY���i.�����`�z�-�v�v/���]��_{��-�[�Y�T�^=���{M[�����\[��=�+��_;3��+
1�>��:J��g�������@S����@��Ov�~�wǆ������B��m�>�#�\0�)���c���o�F�3�m9�T��.�.{��k�8fh��Ug��d��'=�ȃb)��>7�e��{c�O2ڼO}\=���5�S����߾��߼��ݹ��6{����q5�����R�~u�w�OӅ���qW�'��ػ"�Z�{ᏂH.��-�vF�t�=�ֻø�҄ a�^
{�]\��gq!׫�xi��	�̞�=��~۾�k���r;�.�	<�G`�U�Y9M�w�k)\�'$�T ��\W�%�3wO���Iz�.G��T��'�xn蛶c�s�s]I�
��ٟz��*M(��3z��+�����?^�H�@�
��.�g�v��
�Y���o{�C^����+�}08��i�q^���>H��y�j��<C|I&u��L/.^�#�s�{�kq����(b���V7�w�ۻýO�0�_�8]��j��v�.(�p�O��
g�]0j>�1ދ�4{�|O���7F{z��_)��^W�/�vxT@&��&���3�®K���C^V���oMK/�]Ԩ�[,]QZ=��l��'�1{�v(�u�^�-
<S�i	���7"�|���y���O��-���1%²�-�Z1��TVd����7s}m��g�Fd�d��Զ�+w��x'�N�}��_<�t>���ۋ#��.Ӥv�M�{՝�<�71m	�=��3J�?x�1��e�v�I��=a;�Ro��E\�x�k��*H.yÝ٥e���Z;Z�q�����}�c+�b����s�i����L���������#}EH���f��Ke���T3މB$ �5�5n΃�=�G�}�p���]�L>�ɾ�n:Nx<W�w�	����w�%,�ɸpY�`-.AYhJV��Ⲙ�nag�/����\��� ��Z��D��]�ףL�4e�Z�O��դsaV >�^7p��Uu�����4fÂ�zmٚ�ado�@���
��5۵?x��ޙ������<"�k\Ͻ�p��y����s=�?��^�|��O�x/lW���8_h���Ԑ��O��|�p��T�tM�d�H9��Ӫ��&u������Y$����Ȏ�P��`�Wa�g�`@�Ԥ/���A�e�)<�ر�PZ�>�����S�E�C���w�Y_Vl�������ũcx2�Y�{��y�����[9��o��+(���/xE�� 2n���',���({t^d]۹:|��C�֍���F<ݜ��!Fhc31�xA��pot؍�X��ۺ�d'������c�~M칼r�n��^{=4n�6Zxa#>Zo���>X!�8�w�͞C��tM�F��⶝��2Ob��=�%����3Ϩ���߾���I�����;��d+�34}�nɣJ��V���ok6;<�h�����Q�=33:2f����������Ǟmʂ�Zo���t���F��������F"��}� \��/:8{����R�}�&�y}ػ�v`�N�#�i��y z�j�]09B�q�^�p�Oo�s~[�����"c�;���=�=-��b�Y���'�b�9S�����ff!��7���3��(R�\��NMa�T�f���y`���j#4�����#x�X����F�(�W��S{\�W	�iN�r���9�}�6�P�������j�W�C��y>��r/�������k���x�Z���6��`�>]D���ٞCˌ�6D�)�og��s��=�{�m�-�ϣ�<������蝞�g�{�'�>�vG�gi���m|/��;��?f����=�t�>��w����e�޾��oO{'&��wv�E6	�e�"��jeE=�1!n�߉�/\�\m�˷9���ۏ=h�α�����E�<�=��&Lqc[�BUi�f���*KV�W5f����e=�z�=���@����� ����s�����V�9��@�R�����Go�g�#���6G������Xu�i�ť�ײ*�j��1��Fnn�5�y�M�d����}gd�7N�;ғ���+���R�v1�dk����U�M��������������ԥ�;���ĀϾ��@�<��f�]wF��׏{=��w<g�w_xy���U�7���sw�ޔ��x���?Zq`ضd;�N�������j�Wkb;g}����iž�)�0��^L�V�a�n�b����b���&m�X�������rs:����*^*9Ͻ'm��X�;f�do_�/����4��ß��<�Z7�.����n.!c�}ԗ�i������[���}7.u���\�~z%����G��zwh�7Ǐr��g��ם��[�F;���O	�{ۡ/+�����v��'�sY!1���w�VM��=u�F���;_�W�ߥ�Ua�o E�ƵzlG�lY9DOv�`}��__pξ� ���G��H�5�J�==����x������+/�?o�j=�'=�ָG���AΞ�OR6��ϸ��ΏP���L�ﹿ{��S�BSӃ��_��}����V�nv9X��o>�{���{�w��g6J_�[Fw��%��0��\鹹���;�I�̭�M�2|��]z�Z,�yl��²o���j��}�<z6l�����k�9f�O_nv�N':zi4�	���9O{=������JQ�.f�!O�+2�����s}����s��g�:7b����EqO��I�ON���׭��_�����N�~0�P�f|wU�*u�ݹ�v���y�8��Tv^G@���p��c��8�[�Ǽ�>�3)�1�������\�|��v��"���4-��~��>,�*������/_Tǵf���݁��#���ǁ��%p>�ܒ�<�%�䧽�����|jr�n�@������0`�@!���U�����Xc�<O���sp�G'��n��5���_pG	خ���T��mz�ə A�Hym��F=��њ��{�����f���N���8��t�#@����:��~�G��fD�Ί������{]�ǡ�۠çC���gd���+BtQ���V�t�OM�7�ɼ6�V+^��2�1��]��ed�Y���h��e��������ݹ��{��8g��x*mCe\���I��b���usQb3����u�
 �P�I7�Yի��f�T�!��y�doF����{H�����C�wޢZ��E]'_k�ww��-h���v ۬h�f���滞w��6�cS������`�Z�_x��mm-�b����s�'�Vɏ}�C��3�O�*�z���_x�G����ܨ���},<��N�lɂ�+�פ�����d����-��ښ����'����7}��w��x9|V{����%S��x�&ѸFhjU����3LZ��{&�����NT��"��HC�p���ff  �E�������_�����1!�O�?�_�׼���{��7���W ^�f��f�Ч�J��i���H�]���/��}�[u���61���`p��%������3׵M[�.�.�$��yY��ީ�Z�5�"DœU�v��PlT��J�Y��A�6��쳦���[@!���8Ԭ���ءyôE�o��� ��e�Zc�(fj�rEomÙCCm��a������f����}�H�ԥkh�']�٦�1�샪�ڌbVhjn|:�u��ZٖĩZԕ��4_�~ǳҝ�i��ؖQ)2����!���em����9j��m^�!D��͵.9�Ż_��q灨Z��H�enҁ��	�D�@�O7R��K�[��kU&l���K��1��S2��M�������̣�5rQve�3.�1�hZʸ*ٔ8<yu\��c2�@kl�w�w�a��2ܛJ�e��M���a)Ff��2�L�2��lg��#��AE)
nl�Ky�M��t/`��s�&�Q��	Y��WcSsM���1i�{m-� �R�f%�]�u!�V��Mt��8@UMSn7\L�kZ72�
�Qb�\�.�����(�]4$[+r-����	M��n�앩��Z�@��;<��<i&���)��MCQΆ�P��c�n�)��T�"�c0.^T�<��%�`�n2�\:&MBÔ�n\V��`��kj�K�����Ԥ��K6���ȭ�:5�2;rf\ʤeXB��Q���/4٭�a�,a6�fH�JK��ʝ�#��[V%c�7Rj°�D���SM)�k��H��,�WI�t,��3��^��Ð��%��ҽ��lҐ�L9.ZA���n���^$ 6�[J��u��b�lnt�F��öR���TB�B��-q�-�[k�s�r�D�[#�Y��] �m�Mm�f02�lI�Hk�nx0kD/5��2F�f�R� ���bXk[iu�kX��M���ٲ��B���H�+u1�U65���m��b�jV1�-��,\�X��T�5�dѺQ�@�Q�k�@M.��!�7R�lہ
1� ـ��9����P��;R��VFdMf� 2�ۘ�h�/&���!�]eB9���`t��IbIT�֛[6n3LiR�#GIW!k��v&n%L1r鱪8�R�mo2�N2���
.���#A����FcS#�hfؖ�;5IR�9����!�bB�B3`�L�Ċ�X��	e+2�ib�]	D�e�)��Eu��	�k�����eE(V$hƴ��X�KM��42]
4R�`�Kk��v�l0F��m�L��-3���T(˛xf�6��+��@f�͉]��5�F���SY���62V�F6���u��%�*��x�E�,���aD�����c�6�H�m:f�����j����:&�$�(Z2���x�,�<a�iV$i��f�6����\��ж�^TM�ҫjĲ��b΢*H���I��� ���f�\Pj��#56��[��׵�h�D�!�ىLu�q.�f�C��e��Q��
���hʩ*b�c9n�f��\K��L3L�V�e��X�v��,t�d��)��gjL"��Δx5���u�Z�a��m���Fg)m쵕d������,oJ,q)И�4R�S��q1x����Z깭q��Kr��ҚV	e+�u�\��䍋����aF�hbl:e�"�L\pZ�l!l+2��%ɋc6�q�,f,/R<*m0�X�q�R8ⵔ5˙��V":$e+�Vf�XŶ� ���Fl:f�b�.D�vbH�x���SF6�S)KK&ۙZ�\�k�1��A��GU[��QqVY�E9yD�B����[�vv�A]u��0���ii,Lch����1����a��a�qLM��Ԗa�մ��c@��F�3�Ψ�	Pv�nA��8f[7M�p�<�q����UtK��ɗJ֑�c�!�*�����Ƣ$��-t2�8�Ц�3����i���%���9�b�5��oV�f��զq��TLl��Z˭o@����{5��ۀ��mA�����������(R�(a닳Z\�h��A֘6n�vګ+�,Ѕ����4�S �,�*����6����պU���-�K3[2����P`�ĂXQ5�Yi���Ë%T�R��l��Ʋ�LK��V9qieB��X��[v@d��c(��䈑�[Aŏ��lY�������6�[a���Zb��6�tsr��ˠQ� hq��&��XTᆻcK�h�-m��ΤJ,0^l�]q�Y�8�,��ëͦ&.( ���1t�HM�ˬkhP�q��Х���v͢$-��3KH�.�X7B��6,�aH�9�Hؐ-�u4�P�W�#lQ�3fM�Y�[v�a2��d�ق0�5�ػ0��E����К�F�3Y��%�m{8R�%0Z�u�%e�GK]3v�H����س\1�E,�K�pL�Cd��5�6f��U�2S�a��f�b�;GCU�/2��)�X�،��[��Ӵ��E�֢ �69��ͦ�& d��l�K
ь����۪%n��sf����{UꙨ`���չ�%��˖f�f 53�[��k�i[b8AK��Ԕ�a�!U���I��um����\��l�2b���
�GV��F�A�]���+.s��F&p,��)q�u
].l�e����Yi�Y�ƍ�:k2ήpI�bW��A�W��Ҵ[`�����h[��3 ���*��-����ᵠ��V �GG�tv�1�]3�k�Ŷ�+Cu�n�42�m�m��q���G�Mí+S^kS��3�ef�5�MbV�4&([(I�\��pq%G[r#�������	�*GRl[��4�`ěXJ#�1����J5ͨ]j���S)a��$��@c���\�pYT�	�B�H��#Si��(�����G,n�,M+s��uli�++=���)��hM5��&���
gb�vɔ�`�LDک��7h�&�1�kcvf��Ԇ����`ضʔ40��]�0J�I��hj<�^�x��ԑ�̴���Wn6��,+�A�P���!h  WJid٨�c$f��°c0j[[tTGL���3n��+�@;,�������Kn�Il1�Et)f�����eo���+�Z�p�ƄU	�&�n�;eB[��hD�K.;\��MuT�(Q�vn� �m�)
�4ͼ�aqʄ�3ͅGC4���f�4 �3uj���R+�[�f���:WM�L��L��q��F��+��FܹÂ\�,؂��y(���Qm��jاn��)�f�[öRl��Dkk��f�"%FѲ�+K�Q�r⹱���	��2��R!,Lk�1vƫXˇ�J����嚺��.�X�ku�`�[sND��h��Kt7dkuK��`�W1�*i̻0s�lq����"���L�`�:�R]�6H��o"B��G5�G��K��؅)�aI�1,aiS��a�.%�і��(E�Q��]
g�n�[`�b�j�:CK	v�[.��R�иZ�YNj`"�ۙ1-��sA��͏a��JM`�F�j�Ԇ��5E6�ƺ�j�)5�%L!�FL��%�c�Mh�E�v&m�	�L�6.�iZ��L�Miq�4�V���j畎�����&t��ٶ�tV�^1nq^D�Z�:��x��\ͳq��T�0�B�X5-�;Jk](::����Bd�,F��˭*�feu�N6&����)�(�ٍ���l�0�ȖY�1�m5�I��� b���楙v���q�L:7Úg0����bhYI�.�I�mŅe���ˈ���U��e[f�U�͌�� ��ʮqj2MC����,pi�-�qV����%���6bn2�Uu���$�V$Cڼ��p���ë�Lѣ	��U�&8i`���bŅw$֬�t&ՈmW6�]E��-�+a�mK���ڈ�Q)Rʒ��e۶a6�-"�6m�u�0���X͜�kX��q�2�]n.�pf��٭�aa�W"���)�d�V-٢�j#3fu�j��+�0����Mj����,^me�t,�{ސ'��:sb>�[k,YN{CX�J��8�k]��ݥ�l%�@�dkV�φ�zn6�"VB� �k�эҳv5NYD�j��mBkK�H��6����K����r]�����m�ecv�4.������zc��o;�+4���ca/3m�(�]�p���~��j�u�̻K�2�R�͹�[��iII����D0�b��VYxR:}���w6L�� 2[��έ���&k����͋z�eZ
h�Ζ�PNJ�7B̺�]Y`ʅ�t�1���,E-��jK�<�+�tУJ�	ʋ-Z��R����kܥ��GZCFZ�a^*�+U�,�5o�]lf��K@F���e-뜻l��Mb�bQ�]]DXyLx�9��&�\�@����//�"P�^�m*�`��L �1�z�eYA�E/��&��6���Iu,�P�v�.��mM[��PÜj�"/��^����Ś;G|��;��n��X;Z�ۻ�lv��1(�]�p��a�l}��m��Y��#JY���w�������4*�X�lϝ���]��R#M�41�6����L�GPۃ-�RؘK1�1e��a�x�c�\��iB%d-^��6���&�i����Ɇ%,�Q�3���ﯞ���y�Ӷ�D����e@�(L���u��ӭ�j%��*�a�D��]�G����t�j�] ڋl'6���"�e]��ͥ(�@�1�pW[�22�%7)��lŴ�G[B�	v�jj�����R��-Jm��6,]��mƌլq`h��bee%�,P��o��3�^�(�֊�V�s���ر�R��j�Y]�-ɩ��u;'s���w;��ٚ33333�+339�I奢�V����S��W-yo��DU����qpGY*��u;��?>ߏ������������y��y<�MN<F��5DE��ʂ6Š�mm���r�7�%�g۟o�|���������3Fffff|effg>�s���O'�y+-�ڂ��ݔӦ�ţ�SV}kR����y;��gQ�O������񕙙����Q�({�P�������Jl�&-��
�t\�#�j��  ࣤ�
�Tr�+1�V��˙d��T�4IXJ��i�i�I�^��Z:H���P��IRW�� E_P�bI
�0Y$��U*)$
�*��+6�"����Z�9`A�F����nP�p�V�f�I!YB\�PSi	��ˌ�d�eVT��wX�Z��㻹%��^1$0@���b�T-���paT���L2�fS2Q�)��"�O�1)�2Ʃ[J�!�9m�����YIdkI+��1.
VB�iZ�̤�G9��SM��2U�\���`JZKm茘&�a{=�e�6����ԹDʖ�s	rѱ+E�iҤ�ރƢ�e�%C�JBPB�*���jnK+�G+��fn�Tb�!�+��*+^e�K���e%m�P�D��Z�j� I��̻.���ߪ��,:�	��j^�t�ݢ` h�7l�G�82䕛u�@��J������F�;�.�S�g9�yv�j�t�M��1ԥ�v�Kwz�5*K�'{�
ԍ�r�c��%�i��i�2�0[)�9��(�J��ae �6��al�hԦ��\��*�E�S��]H\@%+[u��W�:�[��X�@p�V����.��%
�u*&a�ѭ5�,hK5��"彴�Wj�B�؛�sHE��(DΞ>ym,��1"�luٱ��i-%��\(�H��nl�fTs�v�m��p�0���ԍ��cFe�Un�hU˹a,R�kv�< ��X���],o-Ek[tt�H�:]s	h��#�v��4���*�(��l͚e���ƶ����3��i���hUҼ7&���j6��S
��L�;f&�U�<��W;Ź*�ҀWSp�� ��v�-KYHVd#hk35�5F���UP+��a�a�)h����V���`�y[].��%�cX�M�fe�V7��u5�m�X�\��\hTwh���@�IM.w�.�t�V4v��r ��2ŷJ-(-+%�v�B�.�BlcSmQc2�-F[��q��*�ì��f�֖ip�BX,�F�1�Yb���ݫf�q��� ��ئ�(Y��[4
��b��f��j��8HM�dَ�!Mn���Sk*B�Z�36�`s4�X��E�ڴ`�k�fva^��l�J��n`����cf�Wv��M�2g ���t%��W�îЉ�X�k\�4D��{e�ȶY�x]���]��K\��$ٙ���m�uH�j�K1"EM�[HA%����׽e�GJ�h*)n"�b1m��[Yk��7�if�Y�ЋƎ���f���%
`�����i��j�5(YaSvV�ņ!��:���"��y,aeR]Z�;�5l�t-�u-�0ꨣ�������a��f��3٨��bC]�7q�-R�s,���#A��,a
�¶�U�(D�y�#TbT#m�F�������[F)V��P(���+kQ�PIW����[)*ө^�:����(���)"5+��,�2ե��H���ae�6V<KlB�	-� ?^6��m��%b���l���U�[F�&��
�K�K�(��FL�>b��e,��8�Nv\��Տ��v" �N��[��B@N�M�.��z�bvE7��[R$�@�Y�#-q�UV�yܓ1���j���Pt!��[Rآ� ��;0ɼ��V>8�O�^�q�I,s6<�,ہ%�`�^u�!I&�]�U�gs%�0��{fL�d�ocL�IY���3T�׌Ѩ�)��KF$�\�|�o7�r៾$��~~o�[��	&6�;PD^�"|��$	c������������In�F��ƚ6�Ҁ]�m��Z4s�|���'���w'���?����ol��:�e�X�q��j�\l@LQ���Ӵg�B�`����n���?^aI{3^K��&?q�yB	��nw�Z���>���!�D~�؄��O~�z�/���J�;��u�r3'_!��U
�����~��>�;�=�m��}H#����t@-���[߱��9����P�L=���0�7�_����(k-c����[��=�N�:��RN���9�U�%�܅P�(�p���Ԭ
|p��%��4�2۱��<C��37�{��~��y�͔h_O���3 ;���[+�3,��8p�b��W>��;�C�=?����۵�]Āꒂ�ٌ�	��!�W3�O�ęO*1���D���I����?���qDHf�5�wd��֑ ���`�������A�|1�xv��c�	p	� ��n̒]��Z�C���C��F	i��0�Åv>�gB�z�Z�u)ټ�x��w���]���oe��%{n����I�a����Qe..;��.��u��z�~%����1!��oMl<d��-݆��{&@AM�Q��g�_�/��v|K�,`c4�E�!��w_K���kM�$ϵl��k��sCC��VOy��������ζ<w�:ڀ15�$3[,"
;�N����vW��1�w��TBx[x���.&ku����6�we{!9��w�{}��w{]�Ԍ����R�y���40�eȂ��Y"*�^��=Z�fCkS{D�D1�<,��I�H-�p/̿���y">��}��	2�j1�NX�H�'ĵ��8B|�3^�Y�9��J)zX��ՇZU�5v�$�);۰� ��Ċݍ����b�K�dl\no��Eg���v�>�޶da�E2j[�-Bq�_~����<�q�6q篪���˧{=-���x|�Jb�|=�3 i������d
�n�^�a���cX3��������2`�u�Rx�)0	�N�،c���_���$��d�d�4I
֘�{��*'x��S��������]��/1�4n��6�cn�^l��K��M2���M�D���u����F(�И���'b�� �f��F#���Q;rC8���^2Kh��B�0""U��$������7 �3Z�t�'S>-� *h�� ���N%:EDCH*��D�6�,�u�12�&�zh؆�����53��݈`_A��bBNBi��l��վ�آK�lIb���y�|H$ͣ�^6�4�� /X� ��qA�2# H;�(J�Q.b	'K�i�nL1$�9�#*d䒴P��,R�e�=v,�/7nM�����yzt��^�U�ۊB5�P�Y~�گ>x�j���9~ۡu{��<��kʧZ��,`�10=���)5��2����ʰŗG��n��n[F���m���Q�n���6�A�M�c�ŋ�&(]���?[�N��֓2�83��k&ҥ��aE�3(���knvаB`L�h�+�)�Mh�D3gh�(%.�-d6.m��Z�l�雫f�1��Bk�fR�Xh��Ua�]r�,k�vi��n����v�8M�;m`ww�
%�� bL�0::o�� �m�'�%q��\��t��Y���vr��g�`NmU=�7����h�C�p6�!����@�Y�6 �"gDAP)k�g�F��w[k�'wyඈDa��w�3=u��������>�R�ݖ�X���X���	��j���N��̜ȡD`�<('��`��Y;t}�)�~S�>��Lps���0]�^TxOy�a���$�͈���� ���]%+���5��)�0[�C�w_"�I�3t�~�����z��	�Dz �m�C�I�*� jd�\>]իo&ýR����?���M�&��>jӭ��!
��ࢃ�p͗���W6˲M-�r�M�̡2���4��Ji���^��A�Ê���i��$z�-��}0	z�F��ǴS�l"��I��X`ø�C�:�Rs49��ciz��(ޫ�q��;ZN��sZܘ&_=�ۓ�o|�/'}'
Ǹ��N�9X�w���-��).*PJ �,X�@c�γZ�-Y����1Ѓ=���*u�6VQ�����&�d;��b-�Й�I/j�D�s�{Y����Uvm@7�ĂA��@&�i�@1[c������!Yg ߲['a��rIw|���k:$nDlaȺ�J�oK`Kղ ��I)�'D����@�yz�$��>��8�J��0��:�1��#6`�^�i-�{bZ�(�<�㣭�l���cE�Ǎ�D4��v�H�3�b�m%�hxM~gs/2����|6�	=�����@{b�dl���$����8���Mq��	)�z��<5�Ưc� �J��`b�l�x �I����NhE<�ߏX���`�z�b�}QL�i�۰|���r�R;��눹U��Ȯ��{�g�� ��F
�Q$˅�֜�ly眺󙝝�����b�ř�X���=��d	��̒"���̃�[��'ڤ����DԲ�w�ނ�����=��{:��Yѳ���FyY��~j�0f[�"q�M���-���y*]UO��be��_�uKjLKO�dI �l;�Z�Y���N�?o��/���
�
:�:Ѝ^ke �k�җn�,Ҽar���=�_)U�b��Y�s@���$_<dk���渁���1[<�ʙ#�Ԛ1�A9pi��pߓ���!�ߊ j̙3�<��[��	�S�)Z�fA��%���2B��g"�F2��i$*)c��LY�44ٳ�*� 퇘>�PD(B�w&����z�a�A15��6�v�D����|��6�O�i�+'TŊ�5l�cw�N�TY̬��Q4��!��[�ݝ;�.׋��7�~v	:�c����w���]��J�-����K�p�m<���~YJ�#cq�lnxk��b[���	�[���K��N���zI���p�Ӌ��j��5��D�SAa8�!<�[��pG���,H-�l�Bv^�q���ЄK��:�2� ���`�s(�*!i�0��LaK�E5g���w�X�'ȒO��Ŧ	��1�,&`$�lۻ�1^E�xwy�d�� ���@����鬲�vJI���L2
&�ǚ]�e����pۢ世TU}�>o�6Pa��[�� ��3$k_Ll�{ac���1�H$��w� D�m���!0�<�k���B�&���VQܬ�S��`Fh$n�L{k�{hg}d��jɗ������i��,j����}�B�!yЭ���u쌄}<}��b���Mߊ�F�6��`f[-��ԝR�<xe�f������ �c1'��~K6�ñSa���ݡrKie�8�:�1�XL]4I�6�� ��T��mt-�d����1p�Te�t��4v.��Á�%#�8��m��mk�4m�][+
�)V�j��r�U��GL�ac"�^clƉ�-$ٖ	�Qf�	��nVf�Z�#�T,jK���]sT���X��V��7��-R��A�m��g虤ϭ0��ID��0�V-��fU�@�a�Xō��uP�h�=�NH9/`.æ� �@�[�c�ׇ�a�4��� yqq	����d����OB�o�,]�Nkߦ����;��v^��x*�	$�ǉjd�_ծ"�$U�HIJY>��z��F�Iw4��$HV��b�3�x$1�Zc<�Ɉ���0BYo� ����^�J䢞ܙ%c{*�Dk���2P�вBS7	[ll�'�?���(�ʡ��|s'�a�ED FFZ�����(��y�r���1����N��.� G�f�U�y�(��OF���~�grM.�a%�n]����!�D&5�߇���l�n_T���!�RO��
�{� �q�om��U*��E2,��l;{rDʱ�]ׁQaԐm�s�(F2�ጦ��;�!GS̑��Ɏ�i�o�X�N'�}����~��~�a�!��v�8�
�a�c�Bry�o҈�O7'�E5�=�2�"�T2�a�#�6!���� ͭ�0�2Ef��/6G�l�ғ�%2U[�bLo���h'	D&hƭu7����M�����#n5���g�9Ј/	�^N�ϓ f?ngb)��孼�#\L��A�9ۏ'��D���,d5�	#&i�H��7|�����=��f�{>:�[c�����f"�iV�)le�],�5B�5�LC��:e�r\k*e�?�d�9�x�C0�AI�#rtQ��2j���>�g�ua��r�ҝD2%����2���:LSm~Q �ב�ޏ]�_h[kD6���R
�s�m5ϡ�}���3`�}g�i�x$�u85So����y���3G���B�z�^�Y<�\w�w��OX9�'��z�y<�>�ۏ�~��샨��s}���[���܈��75�}�$�Y���ln5�.Ys��A�p	K�\��z4���4<�/l�7�
�J.y������3�h/���z��ݛ��Z
�g��k
v3'�{z�f��;q�aG�֎h�"s��;���\D��&�/x�Ge��a�hŒUm��o��z%��w���iv�WwG��}�$�m�ůuO-�ޒj�*g�Z����e���3YG{���>��1\�^ѝ�e���V�G�gJhݨ䟏�����Z�!�u�&i&n6�;���:����'�z��iU3��*��<^�D��%;��~����7X�W�9=7n����qu�\6��,~�D������Sc��^��9�9�\UW<��yU�N���A�:^���g��v.O���=��'������"6�P[�Z�y����v�N���.�!�G���dvz��3VF�����Y$�˼�rh�{ˤ�����l�����//<_����n�8|j�	dI���H��3�~�c8���q8��L��{�t���z��ׁ:
O:n@<i�ٗ�����X�6���n#����a����Ĺ��cZ�Lq����y?.���?�A�FL��P��*G�N'�mҲc	�5���9�F�{�{k�z���ub"f��\������if��8�H$ɈZ[EiYm�32TTQS��FԵ�.�X�S���};'ӨΧs�������3333>2�3=y8T�{� �������)D�Im*���Ej6�Uy��332�?��̬���ύ������"��,����"!�G�m^�F��A-TG�̭b�=��s�������>>>>3����~�333��O'�Ɂ�ݴ-�*>��A�����\�e��A/�/o}��}�������~<||||~>3����W����ff|h���N�R�V%h �T��|B�"��h���Ŭ�+*��e�k�0qb�*,��I���Z0`���-mV�J�Em(��%-�J1j���=���U1�Kj�EVҍ(�Q�8�B��@�C�lвT#���Cv�e-������j�iiF�m��l��*Qlh)m��b��cˉ���*�V�TQJ5+iF#DR���qQ�l[h�4����ܣm�Ь���*�z���y�m��FYIe��YIe�
@��Y:�n3�d��J��{q��7M�L����`Q�㢞�C��@j,0���qמ@����4��dy��	�I�,fb[��GOg*Q'b�3LXY�`=�x��E��kgAc'I/���la;HSr�u���!���k���S#�j�6!�S߽�M� {�LaFg�M�\������:��: n��Gy�}Aі�$��\'Pa�>+aw2�VA&�qn����69�r��]�g�XK_�	L�3��^�!��	RE����&�$��z$��sN��溾���x�F0����C^Y%d�'�f� k��\��\S$%�Y ts�71��)/�o�!u�'p�X�ְ�=��
ø�2���sa6�,�'#&�]䆐��=[��`͏4�,�hDD9a:�ѪO7���2V"R�CϷ�Ā}�f��ap�u�I4����!�A��a4��fF{=^e�*!�:�śz}u޵���0�C1`g~�ShD`$|��Hi�D�~��4+w�8z.o���zG�Ñ��}1s^��wd�g�{��+>�;��������8�CN�f�f�*W�
�:~��O"�y<Y�W���~=x����7Q�M�[g^���T���mLe����f!�1�$��c���� �6��k5U2����0`8�rc����n���X!t�MP�\�Z�E�p��]i�����f�0��fo�r]΄�<"�נu2`w�)��cq�@ʺ�jl���g̡����A�����wj��~���}�?|�w	k��]��'_}��Q�i��J���Q�����X��	�q�R���Ɣ�׀X승}׹����qD�7��n��2@+���hD<:
G�ߦ�	�F;,̀��b���$&Lgt��$�C��NgMn��c�<p��V,rTC�u">.��,�����}�v��9�j`��n�D�����i��[˥�y�}>��>��*�F�Y��Y�	�^~��/��y�W.����-{�=�*�g	�z�59UN~�pa�+�0BBg�a�}�K����Ԥ��K,B��$��
O�|��֏h:np�[)�`�An-��n�u�Kunv
��eژ5kTn -nC���&��2��j��$�1\��d\�vpCGM�4�A�G5�[�ۦ�Yz�e�TcS-f��GT���t5�bҪ�Afɴ��&�Q���ZL�;q3��p�E�э[R]���H�r�sZ�Z˵��Yn`�*ᶺE�a	J�D�gP��J�W������sTj-��Rj���8�lZE� �E�]o}|{�^�˯��r�!h����̀�� �eLy6.��x�p��p��g�2 `@9����j�5w���
�S��;V����,å\0�O�L�Z�5�2@'ٻPo��|�m���'�L���	?�����O��[=1%��^m�ɨmgpH/}�T6�Ű�y�:t�@:�}�!�et�� �O@���0ۇt�[.poO��}�\;:8�/IN8;��`xƥ�4��{�EC�s�_����{ۇ�J�X0*�'��1Һߌ���XD"d�|�Wu@�I7`G���/�bo�4�72$��2gp6��r�D��z��(�I�cWP���[��vk��J���.���dt���=��*��F��5e�$Le������%p=~�~���ގ����9w�$U晧X��TD/P<ր�������gȣ���<��w����wV�������3�w|��Y��wf�f�����u����`�N瑤e��X������~�@c� �H���ѧܶ�� ���X�0��%8�Nx�<:=�^�%BC{֢��E�ii끌i)����)�!�H�t �VhK���ꉱ��]�|� ��H t�D���I8vgYm,�\�Lw�,,��f�.	w��+��;��̤W���׈d=��tY���]��]�0ֶ���=���Hu��P�G{����6p�>��<�Ͼ˪䅆����n`ٗ�-!	�$s��n"^��Ԝ���̪)����xt��{��$�]��X�A�d��^Y��M�Y7Mdq8�~��A�^r�B0��4�I��2�$CM,��Y��c騀<�$�M�P�<�s -~#�WO���y�g���@��?�<�@����``'ܺkk'9�7m�l��PՒ#��>%��9�{ҽ�^yzN����W;�y���=��V����n�zr�2�0b�[֌�0��N�%� JFX�2�𨊫�iW}���9)~�Zп~�'�u��
Oy��y�WN@�{���6J���@'yA�ѻ�VPgi�� k�FdD��V`K� $��Zo$^�@&�odH7.cy�X�2-���Ik(
�P�����q,Kv��h^z������A�!�������s!m��� :����zJUS�:���;�S�e�5�}/,x��blX+��>���V�� 	��mj�Y8�@�u~BZlo�xt7��2րL�Y���;����M�d�j�P	�w�(�M�oe���4����a�<:�)<%�&X>)vWhS_.�e�����Ms۲�@$�wkU Kg��xNTD*v6���h�f{��Ղ�>Z ��`� �H=�-�M�ە/�(�����������M��j��qg��"�M<���T\�d�[�Uo�p�������N�Ay�0��k|����ĳ��̘a2ds	fL
Ŋ�Q$�h��=}Mw���[�E���س滭ə$�O�ou��\_%Ļ!���f��@C=3����R ����$���d����!���~��ت�,�4U���F%.y��ڶ�1@!���=��$!��2d�Rl"S-,�e�+z�� 또I ����)�����.�����bG�]�r�q�Ulu����
���lcԗA�vH9�]늢H��h� ���jsf�x��{p���q殎�h�#; F��{b��`�F�c$�c�X2�ɮ�xC+g��v�vN�-Y��,r��u#�M=���x1�x
m��M�ܱ���5ߍ�R�C��?w;L�	{�*�P���Td}�h0�{�J�6 �)�j�h�l q�52 �s�=�����1ݖ'��2��M<��l���յ��w}�탰��/�ĥ��8p���B��c����Mt��Z�0]�>�GL�Pbɜ"�Y�&&L�PU���G��:��vsԃ2�2h�Y��I[F��X)�B��$�9X�p'�y�X[)���
H�F���9���s`�(�j�����KTTtQ�F&���D���s)�hZ�60���G�Smؙ���f�^(7*A�m4[B���m6�+1w.-�m,(] ��Ap[ˀ][X��W�M�.(�cu�CiF�WEe0��c2�~�����IA/���t�B�s�IH1�Lۆ��3�x� ������x�V�mBP
˅�O�~	���lh.� �	�v�vCbwvP,쳮a�2�ý�	��
�T"^<�yKF�N3�L��(�L2.0�Kz �-S���Q�y}��<pU=|��w(�e$��Ɔx�v���>�pA�~�Λ�7Q ¾�,z�����PH^�^���)���P��>��kc�#��A �.�ۀ�H%2C�:okJ��WlA�K&�"���P�;�P] e��8c}��"�/M��G��:��2 �F���.�ь��L
��o��3�}�*׈���Dx�,o�m	��v8���-��R����D�*�������0�qXs��o�0r���Tr���H�`��%�5Z�0JqA8I�L��Eut��wb�D�o �7��y�j��T��w�X�����w������
�i�'�{�\����o��rl��q:�7�c�WG�:Oĳ��\#2`L&L�
�%�0!U�	�T�X�d&�o�w�~�FlFz~��6	���m��
�T"^<�{q�2�[�4'����$x����no2wW��^�wH��Y���Z.�03#�֡�>�L�̐+�||�����C��ʀLW��p���B��l��ȶA���/�8@� �0�i�&tF��$��vv|�/������/�y����x`��ulX�iƦ�V�C�,��Ι�^0��,Ť���R�9%E�t�6濰��|��!A[�Ƣ������q���Jz��N��`�!O(,��e���>/ʈ�!�Z��" !2��^.�v���@���ݻ,!�"wݍE�3Gv/����ܩ�.8Rq�$�@-��� O��p��S 
��{��텪Q'����������&���[uO0��-���Y��^�EM[Q��H�>l�<�Si W�&���L%�0��̘Ha2d¤�I"��d�$��B`M��?ݓɘS�t
� ~�x��%��/
{(����z��F�=]�)�*R׻ĂE-��{~����@�Jn���{�3�N�N-�j�p�i��w!A]��i��%�"������|c�<W+�������3��W�e ]�B0��k0��Y�a���4q6� �He�Ц�$:�8�ۍ,O��qd@�A���<��[�S]]��&��^�|+A�X�;�PT��}(A&�U�8�ke 
��[��]���0�Sk�)�Z����W8b��h���,#�NTʈ�(;-;>x�g-,�����"�K����T6 Ϟ�� ��w-,e$9wP!��ԓ�p��y����9/�-�,��'���WL� ���+�`�	�N�^_|�	�+	ӗA�=1OO~��|Ut�c�a��LQ�oP��/۳"	fQO0�E����<����g:�33��MOfa&̘@�a,ɒV��&B$P�"$d&B~N��g~���!��5	g�������?C
ӏ�*�=��h&$�fv�1-+<�8�uٽ!����0u��7�g`�7��wP��dX��F0F�Yt3��f����{�d���~��K�i��Jx��A �̇$؀R���P]�0y��)�]� K�i�����S��xt�5{������X�q]x u�	�$�|�!�7wL� �{��Y�6<q�c�A|5q�)�B�O�K:��pMw\H�Xe�/g�g�X���H帠Ogt�$���P\�xT+���\±�Kv�t�E7�Ú�zb�0��mUX�&׸��}f�N���稩��{Y-O�k$<^��xC��$&�g��,:����y�N;�0g34
% ��C-]A̳z���� �ޢ�6���E�Ư�,c�5�����}�wN�<X��G;Î�z��4Ud`�X�Λ�)��;[�`�`z��b�ۣ�d�� ���]�|!��K�ON��j�3:b���a���WTfw:u?̬�ᅾ��'.�#�z����64���>�M�|��Ӫ�#/�fo���p1�n�d��;���~�ޔ��f�&�4Z�u�^;z�gb��<뭼r�}��I�S�R���7G����->�9����X�k}�i�x���(4q�(�,{8�οjx{}����������ho�l�p�3|rb��y��F.]�콍�l���ؗ��W:���Y�T�^z�<�=�����]g{�|����P��g�y��n��?_b�����*V���ń�|��;�쁿U����p��@OG���r�sc�rK��)�\�m�ډ�ƫ�N/,��Ɛ���,�tm��������%0C�rY�_|�X�5�5�kLvp����.�5���*�5煨�ˢ^�wv������͚X��ƍY�?���kw9g�e8�p0d���g,���"� #�>��U|�ӏF��{�wvw��ӤCB����%�3@<���<�H�!0�~�~�I�3�e��~�4|�IK9�Fr/5�^ت��{)O2JS�uP�R-����	�"3�um�r��Cw�*�������`� ����s�o����o����� 1og|�߸Ѭ닗ɮ�%ERھ5\�UD���2�[��k*U���]R�"�F�m�S���w;����|~�U��~�_��gƌ���ɹ���R�
"�҂��ZTmG�U_)`�4�1EEm+T�f*8�Z��s���{9;�������~�^?_������~�4fy<�7��PZ�QX�DR�j1[���lh�4�R�K�6y�{��}���oǏ��������3���~�_����~�Y����y��}��VJ���J�[�pZ�yL-�]5E�KE�Z��gs���{:�N�o_���3<fg����~�?c���{2mf�1�ҕmKEkx��A�(�Z�I��eB�� !�Rdou��B��kUQEz�N�嗽�GI�UAsW�V*��)���Ȋ��Z��Y(橊��&��:L�B�9qUJ�Z��֣-�ݴrZ��fE�c#�*�)^��-�̔�2�KmEE-�UQx」,/^��V'^�>^y(K
[q*,br�r�]Ķ�*Te�]h1ETrъ�kE���PJѴ����m��3%���d�ql����o}�3:/e�.c�&1+F�f6�,B��#�f�%�.
T�i�Ļ�5��ͼ��,Zq�Һ���(���a�{�;�;4D�n�G�w(��L���6�U��7f�v�as�f,du&h�i.�LpfȗTLLLT��5��e�#]�҈�RXИԌ�t�u��&���ŋ#MX�e��q��LFkG�f`L1��.cb��i�,nG�p`�Ƅ�mm��K��\;�ufXcV����͖c^Yls("��Q�ōi�p[�2Q\g��I��i	�V.d8Ђ�͑	��Q� y��ˬk��K�Z<�����&2��Ų�@�`+Z�]D�]��.�M���J*�sԈ��ٮY��r�-5�y�p����J2�GB.���ƍ"��D���ŗ�����+[�n-�Z�,��9�Fł8A�������: ]�5�Œ�2�d4Aظ]�!b�����j6WX�h�L�%�h�2��t�3�ی͝������[J��6��V�Ks�
M
]�man�j�@v�J1���g9�i���4��EZ����.*��H���d�l���)�T�%&6][,[D�[h�6�+R�1�A�Y�+���v��y�XVdȃ2�Eˌ�C�&��ذ����ʷLP6phE�F:�l�h���[MS��W �v3M.FY�F&��-,,���e-{b�� V�M�:�]14I��-
cm"qef�&�V�"�.����s�/n16�2D1pͪ�2��-#4�T�J7��YK`��f�@�y�HBcU,ݱ�6�Z,���-Bۣ�M�`hF�ࡻ.fu�f����P&�f���8ю�5Ōl&aI��U�vZZ�e%qcv�TJ�ɄaOA������W5��h�
�k�����d�`�Mݘ]�hv�:�M�$���)n:�[\R�J94^&��qfs.b��B���`b�ڿ1f����&���$i,�S^7mkvX���̮�:u�'�8�ΐ���W�d�i=x�^�{Q��z�H�ڄP Y"�����cә��S`!�Ʒ4*	�3W8�5�Dt��yqhB\k,�%�ť���\@Уjb��c�Ka�M�L��d�H[acp\&d�\ٍ �-!qi�va]a��G`5F����8MeW���'�v����s�r!KJ�GB1�sa�X���eろ��q& �R�3�˳i�� 킬x��b;[P�RRk,#�a͆?$�?z��������.[�&��`�ʑ)r�`ۦ�+�t���������k��<�'��&	��� �"7�$W�)��>����3���nuj	'��fY �o�^p��[*�@��%�k�?X�����bFx�{s}�I �޴Ϙ�O�"Y���g�rϷ<3à���A�Z�6ZǄ���F�%�;b��<1f�]��虆^c�w��	}����DR<X٨�-��N{c"�5�"�2��a��	��c�}Қ�6�5��U�x��o�
���Q#��cR��\�^�VLzl�� %��w������ ����@br`z�tw�D��=o�2��>�ww��$�A�mt+��d�r��%��Ys6·��O>wt^�~���J�;lm\qJb���H�ܠ��@�e�o3�ǩԀ&�^.��|����C̖>ְ��!,Yh�^��@�z��C�	:2������޽6��h�q�O%ի&e���;V��es�7П�{s��f�����s��3�HN�`�J���$��d��{=��O^+ע<z�^�=�$["Ij$�����#�X�� 0 kd��0�'s���t�뚌���HK>f��Çql�]��x#�l6�f�٦�f�:v5���IFB�]��KWy^>�p� øR%��l����:���$�l$�9 �ݔ�.���s"��`2b��zf#<5Y�ww�Ëσ���3�7]'�B������L����m�	5V�@R@ ���+xb�}�k�,ɗ��C����։]������(h,5ΩU�چ]=ﯦ�be�}�C�F�E��7專>�ͧ�l'����OC�H�T�I�p�Er���c�rg�C�nb�@�w����gjg �*��y˘����{��`_
|��%�C���o2l�!��K��,��������?�Zǿ�,��E=�g�#=S��M=�_8>w���Я{��ۮc�Y�����B���a!,�̘c!��d�a �c2dA@Y
$��)�A=��čd���K&P[+���XK�;�2�+�,�=�lO2�9���-�J��=����oYM�1�C�f�=*ȑ�m($���~�/ÅK��@e�nfd0��{:m�Ջa�7���o3��矿~�>�~�K��F62m�Қk2J�T���S6¦`����?,^[��x�z�X�f���DZ))-lG�ؑ̂����2%k흎�fmt��`�)8	 ]�Ē�zO���t��z��L�.`�e�v�,كc�L�O�>S��e�Y����E����S��1�N�����N�8J"�V��HL��s�J,M߽��+ ���އp�H.�/$I,쫺`��O���%.O��So�㽜�wX16�o��d���P�v$��?ε[���m�O���֭#a�n���"w�^lle����8y��U�����Kk����p��y������z���Y�W�X����R'��^+װ�h��{� P�3&@�2 
�`�,!��j����%n'6�����m�@�����U�-���k�Q���B���$5��I�n��(���3�]���|a����/��f���l3a��%+u�o*-�٥��;�/$=�ǹ:�QB�p�m��B�@Y#cL	ο eME�z+K��f"�nb���֙L��:��ww�JKx��Z�w������D�	�H<6^cy����M5��c&p��6ol[X4�HwJ h�y��&v*[���e��n8{1�ҥ�6 ���%3����h�B����u���8xx��Mؼ���X�Cr� 5�ߣ[�N"�gT�g� �z����z_#���H`~���B������z������2ݛ�I�V�F��^���Y ���$�Ɵm�쉁#��{���%��BsWQW�Z3���tg]�P��ܳ4��/|�;�L�3���ۺbC{�s��}w�[IL�a�XϦ̕��=W�`{a��z�#ڐ��I9'}Of�
pպ	�[v.����c��)lɎ0�`��F�lE��`fd��c�2Tq�hhͨ�0�)��f�v���(k�:�ZұXj���I��kV4HP%u��1u.���3Ƴf����f�q1,�ܩP����R�Jk�6�e�6���!`��hp��X�5�]�i�h*A#qPj�<�9.rl+\)Gd�].��WV�c�wi�Ӈ�x�w�cT1!0��-(�e��4v"�\�&����>��*�x�()A�e�|�["	 ͬ�gƆ��b�ē��> .�N��I��}K����r�*C�"��i��$��*5�@5�2{w�2`m���
�s�� �@�I�50n~�ͻ�ӺwԹ P�T@�Z�10�cT�sf�w:m��$
���ld�Ϥceݎ�Thl�wćt��_�a'�L�"��UvQt0�(��.2y��f�kx 1�'�]�8,B�Y�l���]��B�"	�tņ$r�=�Yپ�`Y�: �/ �fĐ5��~s\w})�
�Vz/l(���ϱ�W.m���:�*�d-�嶕�aukT	PVXy�YCQ���g������>����<gt�vNĒ7��{}'�P����� �{�dT�aJ�t]C")�?tOUDDs;�J�B�=�{.�����?L.[c���r�|l9{�_;wt�����tG8{�t�5�j�u�����Y̹\ފbGg;p��A��*�"������a=� 8�jΘ4����w�ݑ���f��|B��V+3K��Ѝ�鉬h׃!��q/����;0b�����v{�cK���h��S%�C$��}�g���_oR=W�d�<z�^��,fL���a	!�>���~@�H>Y�*D���K[N1�_�������/\C��]� �
!�o{�=2X�؀5�?���V�c���|}x�ey
��An�馤��ށ�<���'/�&�I��&�:z�^]�0�dI8�
o<N�\� X�^b�.�1�Z8d���� @����K����C¡Eg��r�^i�^�⳽���/��҅�̑!�s�3D��[��X������]DR�b�Dr.�-����,�jK%`i|�oD<L�Sd1�o_o���onxw��֒`60��a�zA�  ̐\�p�c}u�XLn=�р�d(g^�1��}P��P���뱓I�K����c��D� %��h|�{��/?�V�-C�e�I��6k_g"��t]c(�c�gI��-��� �m歧:b%M#g'�*�r-�$@��K��wrD	�	p,8����z'��0"�n�2�x��Z����R�im����,g�	$�#2`ā��d��%�ɀ@�$a$��I�����;�NA�����.0Ku��uD�{�?L��T�����1 ���~3�*<�7r�\��*8������vW����9�����ʧ|Ibv�I;%o,���Hk��>�LZG�Y�*$� ��;�.�;ׇ�oi���ϯ��䯍n�Z�J9*��ml�&�R�f�3&��7��Ѣw���~���7�����%�7����}�j�j�ہK��g|��{�@:�0=_��T��˙r�L̍d��)��E�A�X )�AbI ��M��������s�< 
w��)���
h�YF�dO2E����MY����*�-�ָ�aS��n~��������*���Ug�H��yLF2`��{�� ��|r;6z��"�R[��R�\S�;��J���3�h�,���'y�0��j�RuR�N	��DD�ݘ2�ʼ�D8�� W�H�Ǫ��'�B؞�W�C!2X̘����H
8f�9�L�I�Q��?�˶D0�H�,�_������CX� )��A�I���@�F2ޗ�=�[�cS@��9�yj�ж�W3�2�ցJ�GD��a���]v"�=�XM
�ѿ>���uɮ��?.$�����d�2@��A�o8����p?�y�C?��A ���%��ASćt��S�*��~�qy��N� g��d$o�&I$�s�i�>�3�x�X�I"2+��N�;���o�"I$�� �*_��@6�M
��6luI�y �.�Е�B&!B��vC�;?����k�۶�%����L*	w��s�ݏP#gb�ib��*w�;H����):�ATWs�_g�Ո��>1�X��o�Z�vvZ���a��<�ex�p}��;�N��*݇������<Bgφ{;^��_5�Ǩy<0�pJ:/r��|<�l�Trշ�	>���!�H��{#�bG���I<z�^��1 �@��
ߟ:ݶ��XL���f��aa��&�ܧ�"��вț���`P�m`;D�u�p�G�.�]�(�c�..e�����`#[��aI����VQ��H�m�bc]e�����SQ�2�]�]��a���i546���ĵ�g5�&�1X5��T���b��5٭��X[�׺u��@ʷb7l�S��t���j.f��<~I�>�N��l75=TΤ�--��a�э,\�61L]pVlX����߯���4�]z�"��4��C̑.�&D0%����J���h����t����'��F(�Y��F���N�	ԏx>� I�=��;��<�w"�$c��x��D�8~���^��{_f�|=���AvM��I�C��{��L�@'t��,e�x��t�'��
�����8��0[U1rLw8KK�zP�'���#za��DϠ@.��x-B}������0� �h�y��!K%�URv�P+,B%�B�4J{����gՕ[��l�{����*�,�$G>��&@[\k��i�ӄ�]�^�]�Ӥ�X�؃.v��#n��]��l[�}�Z��KCK�y~��ߨ!9�ڐ�2v��)�����"��i�;۴I�ڄf�]��\:��T����p�ɞ0P>�+����F����h�=�������ng�H|�"ohײ�$��F5^����
��*Knzu�P�W^i9����@'�c72�L�3�$�=W�Dx�^����Z`sGe8��cS��<�|���D�a7�{�C{e��H�7/eܧw0�7����Ƙ�̲��� �q>��E2@����X��udB s`7��A!�(x^���s�[=6ׄ�{�J�f�5"X{�D�)Y�$��� �F�ӥP��O*�z'`P�x�<c&�
|�1�yO�1�4Ş��dR@�!�ɀ.����o����}��ٽ�4�&���F]�b�mkJL0�24�\�9��F��4������f�I����ba�c8C7��A%��B[o����N�8ƽh��-5}@T2��p���]��%{�J�s��$�@r��i5os�ib�� �q�}����oj�2���?W�y��bC����` �06�s�hty�)�����Y�#vdQr�����T��4)��.zB�y<}^=r����^�o��gu�o�+�1a�{��c�ڋL��CC��:<?9�;�����5��1����{''���x'��.�l���U%��ns.hG�[��e�������Ysz�G����A�uξ��&uS�:ϩ��4��T��[ձ�je�#���\չ��K�{WA���{^:��f�Ɠr���^����{���X��;xf��$]�0�5����cF,pS����j�np v�=��?#�}yx�g<�m>��pK��^���#�8ɾ��� ��9�/@���\�A_^��,x{�7��7���)s�m�7��:������x���3� �� ���v�0)Щ��
o-nr�=���d��&2����]]�p���q�J���F ���od���yv^'�gs��.�:�.�F>=�*,���77�1-�q�����wh��A�6�;�#7Q��~����7��/}܅<t;svl웞��˞\󻰬����_M���_}�و��	�ӶY���vb�3&wOr�1$��w�O>�I=6br!���lA8�>����_r=�_!��r� mh�d8��:.Cu21ye>x�F~9���ۃ'6r�"�������.ĵ����̀9�������^��M�^�3��8�񼌜���[���	b	%v��)ĕb������b�*�`EZ��~�?_o�ǯ�����}�3�fg����w='����d��[K
�`�(Ɣm�
��QV#Q���񪈢��vՔi�H�/��������_���3<fffg���������,�[|�[�^e�*(���pTU�Z���U��RڢZTTT[ibY���e�=�}?���}��>>>3��������љ��~��>�/�|�ڶ��ҥ�U=��B���Y�&�b5��bՕ���{������f}��Ϗ���}33=fff}�+3?_O�ܞy��UEUU��X�"-��")�SV�K��f�,�V"�>�&W.'-ujW��V9lX�b�4�7T
*,J٫bE��t�TN�1Q�m��wf8�E������Ub��o	�-��4�(1D4�A-�bZ��+1[ab6����Q�+iQ(�JъիDUGMj����$��e,8 
VS�D��(�PX�Wn9,g$��bU[�j����kZ1*)JԜ��PQJЬ�تXT���}����BOg��L�%��^�#Ǫ��=���{!� � v#�3��S��w���P��"!���<��;��4!��">j�~��(Ee1g;�ĒKݽ�	'r�=1;�ك�-o�2d/}��	�Cª���V8�%��#ND �{71pf(!�l� ��ԝ ��@ �˹��X��O{�+��:��
w�lB�j���Cg%5��H)�I�V�7���f�-~'�A�����s�.]�AS#�� r!����u��z���@�C�1Ŕ�_���%�B�	�θ�`�S�� SA�~O�7��i�MJ�9�2�b'[|@��:��tS�2i�u��4Cw��*G�AHg�� 9k���|�n�f(� �D)a������}�v�Dע ,I'޷̥�.މ�Y	�L���3�:~����ʛj>4�"pc�[�X��8�/{f���3(���p��[������ߧ�v0)���/�1ǌ0���T�/����R=x�^�#ڏ^+ײD��{�Ԅ{'��}���Z�)û��.���� �]�U������s-�'{!�M_;D��@��_�}&왅w��fۆg�\�&�m�YX�L6:��CiI�v5�xq��ǉ�;/n�3��l�݃���1��� �N8�b;*c���౓ 9��*��>�k��J��`Ic7���N�<9�"ďz:�
$�a��+��	 �$u� H�n��G';��~�溚�fzұ��,o��a `"3;��쇘׳�'vy���0'�-�����#�l\b^r৴Q�&��v��*9
�rń�ti�H�#�H�T�CJ�Lۮ!Cy�	O�b�0�B�{���k���L@Y�"�uX��O5��0�g޹�X� wt
"��t��V��l	o�lb�c�[�ϸ���}3�������N��:��8��-{�w��ѿ7�mʧ�������_�^%|��|��b�����$����{<{2Y� ̙,��>c���ՙPr!��.�z��v�2��偶x�7f�j���Ը�6(mm��i+^ �hcg+���&�e6&Ա�-N,p�:e�d�_�ƽ��Rf�l�ƵVؔ��(Ma�� %��]i�ٹ�i��ܦ�X]N&��b�˖,^Q���L�R]A{D�V$hv���i�Y���"Sl�Iv��a��0���7C��ჸ�/)ri�ىt\��޿���K����Ǌ��)�mۮ�T�,]buTc��ԡ��<��{���_h�c���_������y�E�߰ٷ�Z�Q��|��]�3�w�\2t���@��b���}������m�"�̹�@,FwDc%۬l~>��2��"��0��zxx�B��ճ4��O=ô!�=����R�w�5N\X"���gi���<�Nb����w*R���I���T�w 
��$��k�%r�=R�A��
����HL�ىC��=��H>�����x	N��q���/��>�)$k(���<�5��>1�j�#�p���f�1k�,���\:w��"�'��n�v�dHZ�tEnaJ�F0�׼5��ü��X[m���^,��1��P��Kf���@�|܅g͒#��	$X�,�F��Ӆ��� �H�k����1pk�3����C���xl��x힞��e\�v�����'/��k��sw�<����p�9�U�\%7;n?{^v6X�"O�j���� ~�MK2H2d�$�z���$�)<z��H�Y���J�8v툁���x��[��Z���>��9|�ӣd����>-�O��	�Adw���?�{ �@��@ �z�Ǜ+�%������<Ar�⨟X��v��([�Vd*:[�]�̓6�aa$���l�M�$�nM����vH�O
d{�;�r���0ٌ׀�6g\H�V����9WK;wg�Ɛ(;$K{&��dnGٹ�ٷ[ۚn��tz/�όF�x�0�@D"\�s[^�%���V8!�#�Vfe��vij�����#��F�~����s�,'1����ݛ�1�]]�w{���ϻ|�]�� 9!��28׽�Ǣ���7� �;��ȃ���=<��^��FX�F��d��=+4�@o��wN�D�Cx��[�i@Q�͊G�}ezm��*w�@�9���s�ZI���m�~y�U)bK���}AFd�ߌ̔�f9��ɜ0 ���zI+ׯ�+ׯ���D��lگ�}l�9/�[J,�gv����p7p�ӣfAa��Ѧ�t:��;�˘���d��@!~ٟ50Dr9qrop��c�` ��@,@��}z�x��CĢi�H躜8a��T[�	@��S�l2ɣē+��n�gXдú^ڶf6`��&����4O��nx��H-<M�(Bh�&�K��K@�pZ:��`6�`��x�$�xKܻ����)9�(w�� �@�^g�ځN�����I'�)�مV��@�HO]̃�r2��w�Q���b���r#�w{Q�$vKI��[*��ֿ����q�:��0DBj ��m�c�D�� _=�n�� �Mwl�6�{z�=�eӧADa�ۊw53>���H�:=� �q��2�7r��A_<=��mJFH3]O�zD��E	�*�U��]=%S��|z
�,�"�=����P0��Q�Ğ��Y�Y�TH0���9��w�o��fk_�C��rY��2Y��׏`�^�zD��$�I��a�z�>o|Ά�9��ӣhP _�n&H$�(7�^ˇ���N �g\K���tWc�1	�~0b��p�U�~�t|� :wmT��n��k`Į�e^e�@<a�SevR�ټo���e��Z�cCJc�-,\w==������v��(j1��$Lnbw���� ��@���f�+��Utxy�,T��L� vK9��b��v����}��j��t]˒�d�
RI��fv @ �ۮ �<��9����N�N� �XN�g��7�9�	~Xj �1
�g�Ӝ*�={��ivB'� �<ֈ͈Gw���Bӕ9��� +���]:tA�8��@2ɑ�G�"Au�ٖ���!��sw�޹��MZs�.�'��(Y�yU�yo�*�A"ͯTҥ�3*�f{ׅa���!�!�r���%o�"��T�X���@� ��3��v�f1,�f@d�f�d''�����ݟ���$gk@��f�rr�(%���,�k#�s+sTa��CsjC0vk������r��nnST�u���J27P2��aW��i�,�kc
f!K-�Yv[q��.*2�m�����E���TW\m46���,2��F�mf�m���д�R�hl	��(۱͎�,�G6�j��Ґ^�c-�4�����|��DH�&�h�6��%�ګ�I�I6�+��$v�po��r�u��e<;�0?�Ժ�+γ��bY�$$�C��Z�<f��x~5xm���	9�ؾz������Z�xu��	�U;_��~�2%���[��D53�/��"ALZ�Mr�{���/m�>��.���sdV5� :�TZ��&Y"O�`ו�+hx�}|�A̐ݛ�ox��}�
� ]��j���y�}��v�����'�!̣yĶ2Ce��I,z���de,u6Ǳ�1���Ϣ�{�Ӳ�d;!۾h3���]�(	[� ��x[��dHI�ƟU~�	�]�Ϻy��;���#s[@��)��d-4X��5Vk�u���y5��?�|���ؙ���e�)�>̉ �<��WL��n9�R��\˴չ"������ш5@��C���\J�C�s���m�݅y�Y^�fO~_���`�ƒ/��ϛn��ҳ�^]�;�^���[�ie��sW��Ry|��������+ׯ�%z���{e�d�	&$! K�����Y�_}�|�
آ��M�My���WUdO}��kۭ�R�'fTDC�t���Sz�_o]�椘��Oo Aʑ�h��[z�I%ƹ0yy,$�M��������'J��{���mZ�>[�h9�,��d%7j� �I]�*�|_K����F4geQ �^�N�.�J2=����	}o ��ƞ�^�Ӝ��{d�k�뿶w���A�o@�f��.N����"�)K��~��Pj���6�q,���"��0&ֳ`���{����|�c��V��g������<9�	9y~A$^�5��3��OVY�֤Ib_<u�݀�ܹ1E�Z�S� �_�n��G�� ���6�&�c�U\0�K�(gB͈�� �k �Œ]Ɉ4'���p2'7��cl@q;�����G�M$�<:�7W_з��%ƌ��%�^9������%�)��C9{ݵO{�w
�q�y���N[@���Ŕ�%� ̙,�̙,� ������r�g&���b�}0ĳ��ù�
!�n{��&u�q ݏf�h�"��|��#��H~����үS9���LH^�r��%	@�}�-h�d����1s��]�`x�� �>���e��߷zgnu�f7k���c��٢y�$YI�>����6�#uʶ�32�*Ͱ5�j��QyA�sPR]����Ѹ�X�;=�I$���$�U��U�y��� {;�5�/,=���],Q우�O{���p�D$4�,fa�>��-!��]��DzL]����GU���\Nш2+�R�Ku�/f�$6���)�݀x�d��M 7� 
���s̀��o�%X=�W�w�7j����'�� ��͛o"u�3�˷�=���v�}�{"�R�/aϪ�3��m���>��è0������]����w:.��S/��m��P��������I���Ǐa+ׯ�^�x�
��&v�d���L ����;�Q>ox}q2� �_&�g&M����b��#�}X=���b�Zr6(�=��_<ʺ���2Xg,0\��y��-�3Uѭ��{��	�&#�Ӑ(x�y4����iD:;:�yq�<�ϞX{|����X�L���	��S���d{ŝ��w=1��i�Oma�qe�S8{�3,H8ǹ�h@��uC��(dhw����C'ލ�L��]��P�jw �o+yϺ�I��,�a �m�o?H�	���g��:p��A��<ꗍ&,�׷>�	>�z%�"X�TOv&MT�X�������t=*�AD
�&�=,:�y;P)Ɉ3 �؇ow?�>�~��\��5ݼ��g���p1A�0`���hܩ"Z6���/�/z�~@�r5J�w�[���rվ��������y{��{U}L5��'y�K��ūN�oOy��D��H���;iĽ�>����}�j�f�r(b���a��x���O��Ŗ�Psȇ;���7ES���V��Z|:{�n�FN�󦩉ފ��u'�������n{�s������6I�d��]{ ����X��ra���g���[��X�kv��Wxq�:+�icN��G_-n���}�8w&.�R�I:5��n��^�zOwx������Ѓ�R�Ҍ�<w�Y�n���*��,�μܣ�2�cv�Ll���*>���gб���K�4j�u5����N�U�<� ��w;�(��r�'����y �Nae͒p������g�w
�v�s�������������|�"�g7æ�X��w���F�*������pK|���r<׷������c��b�$e�K�ˋ�8'!`�uH+]Ĺ% ��k���繵���w�8��e�6<�ɞ��g>"��n�hø8{|Z��>���<@�ē&��~ưg_^
ܻ��KW�|ϟ����!�״�f������۪J�x{�j��P?�a�FӉ��Q;x���ۆ���TX��m5����f�+(a*/�ɥ����N<� a\ī3�!:qR�N�Ne;Idż���W��(#���ٝR�ok������,�dT�/VL�;|��/ˎ�������f��d-��|�%�E� ��T2�QcS��IA�v�强����Q�҂57;�����������ffz����f��y<���
xd���i��*3�1Ī"�4m-���(�_%KV[��f~3���g�>>>?_��fg���϶efg���/���3EQE��PA���*�� �&I�P�m��x��~>>>9��񟯦fg���<��O#<�O&�ͣ7J���E��ZLV�UXRʥKR��\V��V�Zuxɂ�˶�2|}�\��~>>>>���333����̬��Ԗ�Զ��e��c��ADb�Jw����`p�O��5�@7ᦶP���0f4Q1�(�DX�&�0�i`�I\-+e�Q%]7E+�p�̢�	ӁF���S^���u���Ūin&�i����f5�TU-l�ӫf*�N��3������JJ�3"#hQ(�^��bs.���x-���J���lM5��SL��x��i6�TճK��R�:s
��A��(X�Q'��i��TZּYl}>�?-����s��Z�̆��%Y`�D�vRA|k���+I�u�t�l��,�ڒ�B��� -rA�j��hk(:jڭ6њf/��vGJ�ƣ�$Zh��\ J�/��!K3x'�\M��u���;05v�˴#kCc5��ìHa@��KQn����M+���Q%p�L\[[%�cCY�[��v;)�-�^KLG)��V˩h�� GQ�ݤ���P��Uܬ�GL¶��P����a�����I��m���2)n�[ ݘ�4�H�b:��[�����&��`vٷJ� ��[��Q�R.q-�i1vk���3V7	S5�TceX��"�T�r��ю����4���V�l4�чdsh`A�jb̻#Ԛ�`f� �f��sfcv��-���v�E�쫮rd!��[(�0F��b5�����]l�.JQT���Ȭml�(\�2�x�`X�"�:б¸"�-�7m�A�kM�©J��s\U"�k�� �͗,�H#�5�Z�b$B��T�m4t�-Cj���)]�"�%�-�H�ً�j00+�Ci��e����f��g����IZ�,9�톏�	&`�����lT\ĽW�%�ː�����bfSNa��ei�"+��B6a�clsط����YV��7]Dƺ�NT�;b�8R5C4��Rb�YG]�2�je+�,��J\��4�^�+3L��2F����7�c`�p������k˱��v�#[v�J6�N�7,�,j���i6�BlAc�P��*��K3j�+e��3e���f� v�spF+t�Ks��F
��PƱF� ��2%ټ��d�vˆeu�ھn���^�,�
�,n7hh�bY��\W0΄"�(Y�4j;:[(%.�����9+�ilX�,�5B�kJiqetE�+̡�cC��,%�	���6�i����!Π��˗Wl�5�-nj�0��ch��jL�ֱ�n.eѧ��?O�R̐�K,�f@�%�!��Y�̒��=��oZSq�pJ�85t5e*�u�d�H��Xr�֩�1EԍZ�l��bkm@HT�ѕ�6<�fV`Mcm-�ڑ�ږ�9�hݢoԚ�6����f���ـ)������ũ�ME�������cV��2��%�k�+���6�mp�\L�&Ыq�m��T����"���XKm�EN�Q�B����.���P�����΢`p,�Df^).����u�T�զ��|S�J�O3Q����D-ߋse�S2������.��i�|�.����ɐi�D����)��
�ű�"v�os/{"Z"'���$�$=�� �.��}�{d��YU�'s�'z%�;�}na��z}����V�c^�aY 3�1������ !���ȧ���gxJ`�L���虂#����8�%�Jd˻z+wq�r���n��z� ����9qds]�R�H =yj���l�-xKv�O�H�ܖ��1̚�z)����u��?<�/���l�����Ԃ�W�-�ڬ�F�̻���T��W`uM�&��8�N��i���8�Cn�;x�ua�^"��Ўb�ѯk(�;�Q*��dk��·O�=�X���v��c�z_zxŝ���ن9���݀�t�{]��=�M�&rz6/#/=�QE�+� ���2gfr�Y�̙̀,�1%�d�B!ε�	${���w��U1 �G��#Sm��m Vήr���t`@�/����:W�����z�E�oGeAj�q�,��;�&���'z%�~��祏��M��bN2@d���%T������v����Ӹ$�����D]�/���Cª&�֊Q[� ��>���
�A�0�IbGW�@�r�HkDn�Ϭ`�6�O�g���(�\�, $�$�0i(��YYF��6�������H��8�b0D���"X��p��N��;��6� � �f�1$(c?t�e�I�\���=j��ی�}��f�ykQIч4(;C[$i���̺��Ǟ� �{�	$�	o&p8����W������zqp�0��P$^��U	�AodAHc =s�7�\#�S���mn�J����.�jz����qH�Z��r����6�q�d,�Dc���>g�`In#Ņ�<C)I���Ys(hCN����?Of�� f=x��z��I^�x�X�_�*���1��|��H ����W�S�%���}��}�w5
��m���}H��7�	$���r��yeE�ݰ��hA;'�	����)��t���%�d���`�\1�\��M��3�2C���R��9~<t��d��?�1!CC9��Y����n�8���*ͣ��%���[�	:y.�A�q��xN;��oUKY X�����W�I�\��R��c��"��.K�T��d{��6�l@t���w���#�� �mz�o��c	#�^%�;�☵�3Q{�zU��z;��Fq�X<BN�9��u�A n�����z��gC&����΅X����J���q'['�G�ã!WO�"�oCEX��X��/I$&��Dnw@�Ӧ3߱b�]d3������Љȑ�y)黊a���ꔡm�
qh�sX����u���ap��W���|��h�㱺����,�fB3&K0�̙,�2d� �y�������cq��0P_~q�׾�E��Ǥlk$%��MTİ27� &@S�ޙcͱ�V�z��K�@�!9�� AA<��G�E�e�^)���aA���ӛ�.#��;�1���3��.e�D�-�.�������K�guP����='���$���NNZ���(�ozf�d�\uJ/WX��ҭ��zP"A-]}!1rzOv����1Y��ܹq\M�x>bɈ�{�kTxBʛ�����x	;�@ 	ӹ2H�Avd�-l��#ˇ�N�C� �]�LS�3�(쀅}����5�d}�^C蝻��nd$V�y��	Ճ�aш�ڀ�뗙%������7�ث\�N���]�F_l� y���8������0�+}�o��"�U�YE�2`��,�� ^�ȇ��~�%wxK���	��xrGw]&��u>���%��~���]f�3_���� ̙,�Fd�f3&K2O����s���ִ曓T��)\V:�6��(م1�o9�k.\���L��*�F��M�3I��W�����1�ō�jD�"��n���MNݻ&30ڸ3@iu�ZR�z8��J��VRneѭ�[l\�l�sV��6)��m�V�)�͑��@�65���9��0��BQmJ;`aZ�53��R[Tu���ܥ��c&,[��C2X�����DC����(x9D��4�.`j��M�r�\�CXyOTFrD��X�aɩdٚp��9����q��_�ıi$��In��;@[酾��v:ȁ �� ���{�L��c��t�L���oCQ ���艽��0���,@9��,��{��g{��	�X�2z���"!�LO>��2Dc.ǈ> ���<7XA��Z�zߚB`I݇��. ;�r� �Tv%��%+|(�	]�3�rż�w�C���ۖ 7*D�p��E'FԃG��7������qx��b	�l`A2ٽ"M��6#��Z�OH��|��9Cm���)k��cM1�i���b����[�<��_<�z���1n�/���A�����&d����Z$$p c,���;hS=��w6@,	3 A
=x�9����"����	.���Rw�r�ɢb^��-�jr�����o{fz�j����%ㇷ���^��=�\����G��埵x%�}[�O�����^�x�J��Ǳ^�y2Ld��������{޴(�߿jH�}�����L������4���5D�L�H2ݗ�L�>��ln�:�~�������4K۽1�Y~��� ���#�(}�AFy(�����ti`��2 i ����+�$,��n�!��o������wr��A�j[���& s�Ę�L�{@Q$�  _� ,�	���A/�U�ߴ<w�=Y��{�k� M�ї:]6ؘf2�+�\���ZG�QQp���4�H�.fÈ�����9�D�񇸂��y��d�n� �`5Y{��K�����d�����yp�*�����T���=��2o3/ �$���h�oK�-D��g��)���c�?s@�)e��Cy.׈L��K;:$�,�Bǻ��M���]��Q�V��C�޷&�mE)��{9��U�X+!�*��w~�؊�)�\��U
�8&b�|��pᝲ`a2d�	�& �r����ji����A ��XD�wN< �U�]]�U�-�5� ��N5�:���)鄒k�7I:3f6�̗�_K��kj�K��>��$���}򊞟I�	�&Wuαa@�G�Nl�{��O^��e2� ��[��3��-͌��*�,��2k�j$����_�~~�ͱ���[R�@,Je=}�'	� &��6/6|���z�H$��$�����I�ß@#����*�؇d�Gs�R��p�bɎ��)T�"w8d����ص^��q�s�J
��cX:�X��c<}$H1s->8{kz{��>@nnE6HK���G�]''���Y�>������	�����1�H�Hcwl�s-UѬgj+z`<�Y)ר�T���TY3���F�����ht�����B����+�4OB�zk�xZ�q���Q1��=���Y�RYfL�),���Mt������	:�1��q�=����%���Ա��YNt��Af Ws�cbq+3�6ݞ~i�]��cj��u�X-V�\;�l��]O5�2�>w��� ����q$��@a[ݍ3�@�-"UgE>h�\��H����m�A��>?�1����9���t8q>��h���w��D�H�mw��D�Yw@��:{��ny�j,�9g+�M��>#�E"��A����	�s�*^�߱�R�����{�����@�gd�ݽ��h���WTl�Y�Qv�����ҁ$<�s"L1S�Ӿ����\E��'g`���$���:NO�'0=���)�:�c"e���Tl{&��q$g����m�ظ	vH6Wt�'ц��w�?�-���4��:2���g��^�������b�SǼE<A��3�����3\�ƴ�f�4
,U�Z��1Y��N��0�2RYfa2d�L�:O�xh�e�����^D3P���-{\&������#��WC*�f<H�@�0��&�X�+��7�j���B�6,jˆ�an�M]ZQW8�`��R��
�]��V�k��3��%ʠ��m�Љ�66�()�u�{]؄��%fY��J�r�*�
m
�^���$[�Y�jۇ$Mxb�#���5��u#��4������=��F�ש��f���Ӯ��EΨ�j٘fm��}���鷝����x�.��̧v$�7�<ҩ+��h�͸M{��1˨�A%�9�2C����x$<<$�E�t���O�����fHK�zg�z�aK"�s^{�￉�߿'�Y���A7�m'�kr{k�AX��݌�e%��:�˟�1�P�H�GD�/�yȤT9�(� �{u��5�;�w$�:����g�H� ?���E��X0^�Y���P^ B��6�.u�;:vL@~=��^^�>w�@-�q �@ 3_�fE�nޘ�ݬ�U�1n?-���ې��6��;̔0�a`��h�nT�͍���4��^G��H6������0|��I�[w��� ���tH轟@&�L��@2ɇ�׷�d��,a2��d{���hIॣ��=����>���y�f{�4��>$n�n���mC�{R�o�*�Z�,���=b�<N�M㗽h%�c�V`����o�ȫ�*NS���SK;8ggg����;;;0�O�d�	�I�����,�?}󆎯8[�jļ{�`�[o���	�P��`%�Y��Xf�S��y���ñ�K�ٞkg��A��ā w��;�.� ��c�/�˽��٫u'���@ gmD�	�g.ia$�?G��^z�+ܾ�@���}SP(`$ۑ�8u�6
�=@��H�b|��y=��0�X`�X����T2L]�%�[7�X�@���	jd���{�J�:����]ޙ,`�G3`Wl�-�[4pj�W"��q����/l;��ϟ���Pb C��Q��	;}$�M���q2z���&��ƱL�2@nD"'��riBs���x j�#m��h�J(�����()Ͼѡ�������Wq���&�M�A˸���@P;==~w��vAcJ#����R�r�(?��xu��7��sбt!i�$�s|?�P�q�q�K��6#�8ih�| ۤ���x��/�$�s�b[�s�M��*��So���0^�:=����z�Ş���a[� ����;^k"U�y?��N��y>G1��6T�T	��x�vp��(�M����:���.��iT�p�t#�B.������'�3����3�PÚ�����7#�{�f�����B)�o�>��z�+v;֜O҇:?<3���X�˾ɾ�y�k�і��rc7r�n�ʘ3٬�Y�l��ZD�ħ=�"�|�s�n7ƱΡ�7�a����q���C>8���Ⳃ��F�E��hsw��s�������z0�Ş��c�ۛ��T�!]�#`{؆�#������n����{�)�D�ށ����ɷri�����u�ҷz?f��y g;��ZC�{<[�"�uqo>8�V�pΚ�4W�z6.��7���L�|<�m�������?��8gg�b����>��^ɽ�z�C;w;���X4�
��..X�V�,���iea�r�eT�����Ȉ&��"��+/)�T�@�9�%�
7�JQ
���4�O<�oOH7U�Z�X#��X<�#�_(��_3�`�D��{���|������_W�:����7��Du�q�弡�c���g
>_A�v0�T@��8:�?�3���*��%�b$�WI���39A�78�C�K�v`�j��a,
* O?L�Oo���ʮDm�a�yƅ�����<`��@Ӈyd�;y�&��Ql���=;���
�.o+9q��0X9ӆ�%{�Ǻ*��[ѕwL�Wz���ӆ�h�Q���k �P{Z2�R�B&�� �D`=����|�"X�x	�	I{S���y��;�y?/���MLA�YI�U�f8Eɔ�%�{ս�I?�8]��f�v�I�0�U��-��7�[󩷦������E�f
��&
,�
�b(��5K,�L�fs���|||}>>?_�ffg333陞39���2z�S)%���I֍�D��ε�A�Z�y����z��~>>>>���333���������m�l�X"E+); qZ�|�Y$�S�C�/NaI������y2y9<�Ϗ����������ff}33�y57��U�H�b��A���B��SI����hUEm�������ׯ���������Y������fg��{>�Y&��⢋չi�.5�2X��[LfC
ƵRڻ"WH�-�I����b�F���%X�*�j�e���E�:����H�x��S��#����3)e�*�X�\�Z9�(c[l�)�E1�fQv�ǪTv�$�Z*Ŋ��P�f$PP��;�7��X���ݫ���Yr�l�-�*1X��TM�k��5?C�Y�&&JK,�������\? ��������;�̀��ע�!�D����͹����{x;LP ':E�I8�k\t�L�t�;�L�J�0o�w�!×qh
`�za�Ǚ�ݻ�� W��G]��M4�̂I��k%�bs��{[��GMc�5�",^'���	P�]���������0VX�Q����{�s.�/�w�c/�!�#}�HS+�؁H� ���$�vs'c���Q��A�@y���K�u���<xCc�2X�r�:�#;F��h��I��a,I-=�,%��,��;�߳D>{Γ�B�j�,�d@-�h�m�/2Ki��/��ND�s�i �(��-"ZS�!���Y�t�]ň2_-T*a��^	nI�Y�2ı%�'��Ʋ�씕]X������5�[�3�-�#�L�G�����{����b�aև�od��u�~��	�����,K�s� i�k�,�RYe%�RYc��{��Қ����c��]�3��#������I��",8Z���e�����Ye�T�H�>LN�>��nzG��̟yr�ws�D�ƍF6�s-�4��42�E'Ll�7�$:2o�?���8r�"}��e]�	�H�F} L1D�߮��cu2oKd�KKN3��t�͕�/\���"���� �o��s-p�� �d��� � �<:����z��; �B�-׋�*!C����ڠ@$;^������������0�I�]�����_O�9OE�;�@��r�_���C`Uި�"������A3����{u���ދ�G��N�a˸�h��ȆN�"z� � ����PD�42=d��[��� �@\wt�c/5��/};�SF&��ҡy��{����{�\�w7��Oo�����;y�h�\�z�5<�cͽwwy��|oc(��w�p��L��YN8�q�=����nh1.h�`��-�&�b��@ͻ�m-��5�T�(�bR���LB�2j�F�X1.c��d\�
�Hj�Au�V��.L2�h�6	�;k4�j���-�h�J�����9pk3�A����Mmq�dV-)�l�q-]d%U�܌�Vx�Բ�J�IFX�P\�H6$�6R#V�[��3bH��l՚R\��{<ߧ���O�ى-���,�c(���6D�R���nѢ����=���õ5��'w�� 9Q�*���9� @&;������#8�)õ��O�uXFw8�$z��� <.� �'��&�O���˅�Ǯ���@x�M n�0���
{��ąh��M㶢X��U�Fs��}�5���ÿ��D�{o��Ч�x���>숶(ow@�@"����
!Cշ�=ռ�R=u��LPb2{kX\<��������:��'�r�8�z������T��!3܊�`z��x.�&H}�2ǢM^ۧ�9�̗N��H�I�s8��H'Ew8���YUW���׬vL���S� ��.hG��@��� ��(���Yk������X�K�q�d�&C�qbv%m;� �L���I���bXzҶ!�k&]�2���ݸ�,I��~.��@��1dmE�8�;�
�@��}|���5�`��ں�?"�ǈ��S�ϻ�%<w/+��=6{���맥�29��),��&JK,�@��_@$Ϳl���/�� P�<��
��mݛ���.���x�(6- a*A �L�z�D��aV�;ކ����2��"��K0`Otd�R"��rE�\C�KY.�;{۷�/��'�"2G� m�Ic,H��A�F��X�g����8�ދÅ��U"S��@Ēs�;�u��1�g����]�D�-0����!2��d�H�q���|�%���I�l"
<�	�c �)`\��W\,-��o�4���Ɛx��K��y�f�A4H��w[{&AǹIM���S��X���e��#ݜO!˸�&�^��*�
+�su���}�Spk�y�@"Ab
�q q��쫍=>�Z,�r�n2CB�3D��=r)��4כ i&}Y�dr�7�c;�}��G�Y��/�����>��ݸ�S���g��������B��N��!Bg@����`��1���q"LH"��J}�%��I�(�.K��F��9�����ɾ��L��p��������1�I �����@5��#��.Y:Nb��J)�Go�>xO��R�,|�zj�H�{w�Ӓ��&iF1@���ty�);��_Iig�\�@��5D���]d��Q	�z$M��Nzh�h�r�jP$s${%����%ݐճ���wW�ϨO������l�:JW2����`� N��C��$���nU$s�
kB�q�s�:d�W��L�$��q�����^˳#�̽lP���ݞ�E>��U� �D)���P��j�O�W���F���1��C����a �0��QIOwvϙ&�I��X�E�Qt �{-�@!ʮ�]�Q0��P�!q���ML1�t�b[�{ouǡ�* ח�O��Zez@���ޕ�x�F��YQ�$@�� ���<� ���Y�\����-��N��]Rkz�w`{�帒�~ g�[�9B��'!��f�EUb�E"�F�qF`��*|N�s�&JK,��dɐ��$�<�g'.sj�ǗXP��u�$^u�:@�H�Boy�C[/1pY�z5������h�1��-J�P�}�y��3)4Q���v��� � �Mma��!t�O6fC����H6�s�7(��#Q2Y��	�[;�\L+��<u@�A�Q ����H��uP� (���Qgn�ɠ9.ewq�{\�Q��֔�$s�v_e(!�������<�!>f0���w�N��ziS0�=��C�� �}��$��}�T52Lk�ۚm��tɖC3��t����5TQG,���VPA'0� �l�5�A:�ٵLe�Q��N�k���w��IEG��c {i���0S��Em��$	 vc�|w��*SCe�М���"��{�Z)��N`�w3�J|��{�nܪJ�<1/w��<�瞝w;��YKc�!|*Q.<n�^TN0��{ǉ��
"#��7Ss0�2d�dɐ�dɄ"w�K��=���?s�=�n[��vG�d�M�Rd:�F4���1+6nb	Lˮ&n�l�S��fl�1jQ�͈���ia`���[����kwGAr�kl�7�@��
eXj�K5��.��Ҫ�2R�q]RbX,tY��!���\����M�j�aq,��2�F��AtH����3��8k��wJ�۪(12f� -׉'z��^�4#W�'�>ߗ睻��vY� �p����j�2����3�5�}�����3���˯��ZaF}��u��KZ[�3%�$��ɞ5�usn&�KÝ�˻z�jQ�&�|��z{�
����]To��m�%��(�!�,�n�d3"I�s�H�˜R 8>Q�� �"�/ܮ������d���oJ�S�ߞOp
��*�'�0Q ��~薶Hc%����7W�S�p��
�|�5#��SA�rT8��eG�u޶
 ��}��u*���N�i�=vA�駁5��>��a
��CE11�-�2/�b�����]���桮BDr9>ha"Y!�p �n�:ح��4�V㨕�Әx���D�kR�Uͪi��vs,�+.����l�m&Oϟ�,1rv~��*8�A�:D4�YF�Pr����:���2@$]�>��p (E�A��]ش1%d^g�^�"�LL��x"iH�*O{5��zx>�A�"L"�73mY�=���Vd�"c)yZ��`����z�-^g7���x�]5/�~'&�L&L�0�2d�dɓ}��u��;��������<�/x��M�&��f����D��U0���,w�PY��	c����1BJ�xo�1�7�v�|T�OB��YO��zC��>��C:,d�CA-lQ�̘�<Ԉ�)gn����ω\r�vI��-Sn�z.�,��%2nȗ,�Z���&n9����mYhr&�ǃ� ���5���o�R���\;c�*��L���iv�je�`��bcUsp�W�<K2����bjb{�78��I-���y�?� @g��X��H	�=gO���3RS�o��}44�ކ� 'ޯ[�؀\��#�{c�mE�̱��{�EF�d�l������&������1qG0Ar1g;G�/W�p����'Q�7氫����7Y�$�A/�3:���A.U�7}��튉�(^�6f3u�&\;�6f���y�ؘ������i�z���*~1��Q&O��ܤ���L�0�dɓ���d��~��C���$��í���P=@������[G>�59y������kj�=}��ȸͨ�p��a�yy�P� (���m�f�K[���9��/Ʃ,�۞� ���:B��gmT�)�����d^�e�j�u�w���
r�K�lն� �6U��;�mK����?��/5�"�ign�ȠKs$?<=/�WS�f%��d<�k$%+��S
��!����'5D�fG@�d��n�E�e���p&�a�{*��@�d�� ;^�ۥ���y�ng�q#Y .���D�D
�srA%����0�������X�b�wK�e)0��v0b���:�2=��.�9��� ��0��ȐI:�+�i�"��y븘꙾��٫7�^9[sc��3O�|�pt>I+�������M�1���7�w�7}���-a��ɫ�cB�Չ��8�vs��8�q����fz�S�6�l:*��EX�	��$G4�S�
#�xWT	8ǹݠ�!��!��o�F[����RT��Ò��3�f��p6�CA��.Sx�Xh4�<�Z�5nI�@��q
 '�Z�Y8/z�A��,-�'��w�Y�뺙��t@c-PO���GtT��GW��R���wp�n@��=�:A$vO.�w��(���H|κ�lCwup\ȶ�>� ���^A#�3�xi8�=b����X��H����<�K�Aar���丼`�o&m��{g�Z�À1Ă��w���{���_�htS�p���� ���x-=yy��Իc�����h���B}n2����c��h�t&����Ըɺ7ӕ3��{QT�Ow�=��x�}RZ�F6{9.�r�(>O��65�M,���A�'����s���
��:3z=��f�����~�zq��)ָ���&��5�����ny�ܼ�d��q{+��O�O2B�����i~�#�٫�t�[��S�	��Sw#�'���fG�vX4p�	!�c������A�QOVj���7C�{;^�^�zܝ2�����9�3��ҷ[��j��7�}=��/z�w���5<��`_{�z^<�~�+6�kڛٷw��.��s��6�ƫ�5��Ć�{�9�>><�N�:��#ۡ���{��Ƅ'�W(]���X��j{ t2p�J�ö��:�z�����i���3�a�wfu�ɜ���/���x�<)��1{}�47��[ѾΆ�<�y��1D��=��.������z2e"/cZז��b9|��m���^��b�O�k��= �룴��{��'&�.�Ǫ�q]���r՚g�U%�K�ؖnvc�9a>�gt�}��u{��{�������{6*+3Q��p���Q5*!��y�ٷ�Z�׌�C�D���N�`�z�D�wB⩋�yq4�g3�����{��wn�U�a���No���&vڽ?_~QI��
Ȁ��й�bя+O��.��"�C�Uo��y�_դ
h>:y�ڮ���3���z���������>������׏�K��u=a�v��x�Sw	Ń��ώ �0�S�ۑA��e��ڊ,u�[d���~�������������z���ffg�3<fy��ߞ<�U��{�1�=�TX�*�҈��b��Z��e6x����u;�{:|||||}�?_�Y���L��fig�ɰ���X.Z�Yc"���Q�LPiV�;`k.��S������������|~�^�33>����O'�ɓ��'�=�QUb*ő���c�3bhb��t� �ϯ<���Y��g��|||||}�3��333陙���Y�'�ߒN�KJ�8ȳ�J���ҩ���QU�UU6֡X+ժ�b"�G��&R���"�!bx�:hŊ�Z�M�"7������ƥMڊ�jk.�� ]�N�� I�I��x�����ck��b-�o7a��X�h�[��r�U��m ڸ�Y�h��X�ի�Q�J�e�̘�&fgq1Z"RV!-aպG�b�j�&��q7�ki�5cg�5��ZnU�)��PH҄[�ys^K��ĤƆ�;2�ضk)5�4)��4���̀KUo�Ҥڒ��pň�����iv9j�,4����z؆�Qݜs4Θ�/M5���3�of�.K��](S,��GI��:]T�@ܺ���j�3e�K1��qXGY	B�Lܐ�:��qC#�������f�0�n�ec��kPL�.GJ��^b�h��Ft;N���č��؆��du������Jf.����+�)��1�Q�a[L�3�IK0L�Z+J���a��[8����MT��n3[U�����R�L��Y���F�V���f��d4�E5eD
Y�5$ۛV�n�j��[� ����	pP�uN��3�ma�kYZf�6��R��a��-4�<$*c)�q������a+17k#��4�E�Jն��-�\�4	��u�,2��5+����m���l�hmJ&�`�B�V9j��;L--h`���WKV�1&�U�XL���Z���m�m�Sn@t�k��L)`R[���vEv!,�;J�j"�4c�� ��,�m�f́��b)�����,��$q�p8�q���0k�Tmд��u�]e��a�SL-+�d���b���r���K;�B�쒋[L1�����K ��-���%w\���µf�ޱT�]���ƹk d��L�0���1�1I^c�W�	tf�s� L�g��a5�s,HE�W�6�v]���[��CF�[3˵�t�ar�mNlf͌<B��Qk��j�t]X�-Bh��nq�P6c�����]�l
�����6,<�ٖ#��WCnWLR��͊��r�u�萵��+����2���%�H�2��L���Ų��&��.F�rgr�蹲�p��j^U.m�Qe�l%�k���e���t��j���:�B[�]f�IUaVِ���~�nw),�0�2RYfN���o���
��Ii�H��Z.s���tæn�h�f�V�1�4���	��&��ɰX����.,NkH��͗H�0��(���+mY+�&h�cK�\,�4E%�GF���c��Ij+e�[4��(c��0�@�)t�Z	.��]+���!�L����m��5L.u]
�5#V�q��R�;
�vr�V�R��Q�rm)�U�bM+��ߗ�>��g���U���t�rCE.��݃9�0�Yb�F+�|���jiG�"�|�x��ɿ&Y,��2	2vp�Z�ӱ��>����؀�cW(k�P�
!B�%��>���HK�ٛYތ
Q`Ggt��T	kI������&�h|�^ڳ.+)z�QO��x���_uĂ&���r	:�V���2׀�Z���Ad�;z8�����-wW�I>�>~�[��wc L��W��L��wb��bA]�퇝]xKs&!���� �w���AHD	�YgT��8C�dWnv������m�XC$���3L�@c��9��"7�'}[\�j��:l��J)c�,�@m�whi�Ω&�p��[�7�C&��{�^T�!y�
a�@ٗ��0Ds�+� �1�~�i���5��Iy �ȩ�a���ug�DE@�
�P �����N�;��QEd���Li�������I�u��|�z���y��i{�z��?z���Ͷg!�����+)�@K�ck �YIe��Y�3�3�r�KK���9FX�`@,w�������LDd���-0��P���KU��(5^�A"/b2Tn�
�n��&�L���N1�C��b��K���x�C�'���Y$i��X�F{.� e����]TG]��H�d�(2[��]�\3E���  ��<��c��UzZHj:XS>fK%b��^�u߸�rg�cƐ��Ro�U�z#�ty��A	���-�9m�P��ݱmFZҮX�L$��~\;-�~��wT�"�<�z8���;���Ļ�h\qJ���U��F�Ā�@�v��=��r� ��x��@����D���#*=>�$�����gz12Ka{9o
����������P([-�\eq��I���P|\觏E�%����u�*Q��lK�J��]$����,�v[�)7�-�BW<�qS8���6C�}�T�r����C:8�l���A�&A�&A�&Bz.���X�i�?���_�������x[,���vI����{�l(��@�-o��������6.b�^''�K�;Pv�"��%����|a{�������K� Gu���Z�9�@�s����}�'� e���ivX�c����R�����6���)�p&3��@</J����s�Mu�&L��f���$�F�IWL�e�)^I����g�Xbv�:�r�0��Fi�]kM5�c�# A,�9n�K�HD	v�`�O2g_7dAٵr�G2P�@���*�"G�zd�����o$���rl�=� 'r� ПLD	oge��XJd���a	Z�q-^����3����"������SyO��r3� ��n����dM5�����v�۪��hp7��؊ǆL�m�����`���~����!7f`�t��A���+sɔP�^�"3�U��M)1 d� a�Xs.Ax�cy�k�&JK,��q8�m'�oϿw}>�<6��&@�ɭ�&�wL o�7�T^�.X���{[����	5����3�<���x{�n��d���+t���m�+��suդ^U֞�L�'�Z)���e�E�Ǚ��hZئv!n�M2�l^���¶c&�]�{m��A��m�fH	��n˻��9C5���I1��z5�r6^`A:ٻ����p� s+�fr�;\�!�z8qF��p���S�z@��N�@�I�O���cw[ı�C p/��ۈ	�Ј0�G�_�z=g�!C	a=̓Fl@Ĵ��u��<�;s֢�`��̛e���|ʁ��
>��i1��c_vxMUw��X-��ֶvrV�"C<Hށ@�g��g��^��w�x�۟'|�qZ�ݼ�n>�=������T�s��#H����>a֓4�%�0�Ye4��toĳ�Ie��YIe�r�fx��wtL��**��]W
j�5h'+�WB�5�ɣL]�ZHJѥ����.x�\��KZ��mD�q��V�Bݡ4�`K����f��CX/kD�+��ܮ��f��j��4D�m�[jǅv��.���Z���Rj�h�sA��P�U�����73�,r`)5����.˯'Y�ӥH��كөݻQ�)�K[_h������|��/4�{g2LK
LdjYu%�ՙ��6\��&r��qU1[F�qJ�(��"%��O�d�L�@��8�$�$ǻ�ȋ~�꺦e���2�"4{˱�K�\�����>[C�v��$#��3zL��*�з�=s9�[�}��n]���(<u��<�1f^ǃ�lve��~E��2��LI׎!���^�K��tC�kF�rs�o�������:�JȜ����4��` ��
�v� H���vr N�L����.����F'v�|���o3��Ή����y���ᙴ�-�=V՞G�3��[}�Tod�ا,�ϟS�N�Sd[YnѶ��b���m�ss��\�8�W5)����Q4ʁ� ��~"���|�Sfwz���E����?� �?\�4�<��$����a(��$$����vZ	��4j��C��
�������<4W5����n==��*�ޑ�:g{a���f�h!�|d�0fLk�q�8m�#�x�ngĳ���),���(o�١=�G0�]���b��wNV1�5�Ӕ��s��׾E?�pa�H���<��d��!�ګ�� �R�Ơ w�	d� @���%�t�C�|xPf��>�#}�ݼV�# ��
�d@$so�(jZ�{��������٤�Q��ɮ^�z�C�r�\C���>�ĒG^@k7�`�>�%�֞=W���$����پ�]��s�珷�χOx�Xhͬf�4�;W���s�㫠.�f��+T����P�L�L3���u�/��n�����ȓݑ@QeV@��3�	Ԛ��XH��8Nprl;�ꁆ{��� -��������-�Ṁ d��vmQbN����h�����{�Ô
��X�oo�D%�����꺙b������ ���cO��:5y6�Y�{�( ���״V��*�T�uu'W��X�w��Z�e�B�[*�? 8e`�����	�U���{2Y,��L�L�߭k`D��@	$�t4 �Lv"�Ipa�RXRIxD�u��ן�> �!��xC ��vd�%������#�mD����H�V�CȺ<(>�]�4Zڂ%q �p'���>�>��x%�张;&\���jE���}�����_�UHV�5�`d�n��Q,&v0��ͥ�Si(�A19��A&5�?��� �x�,H�=�(k\酴��¾�]5��P�5�2ǚ�#��K�����w��4���;]������� �-y� �%���@;c$js�+�e/B A��m-���{���>���w*0��P5���KN���]n��[��vm��≮y� A�ȀX�qw !�n�{��p�B/	�ގ����{Sz%� '��3�F5�:a�:/���K}��&�Q�T��]ߡ�>���?}D!��O=���枝<}����}uto8A�����{H{���՝����J���T�i;�z�.o{��:��%�P,���(ϓdD��S�F�[;Ʌ�]q���s�{�k�{�g�$ҹ�$ֽ�$3;�C�[����x.�Y������^`�G%�r�U�Sfks��"��ƍ�<�x]y���"���u7[��$��7���rA'{<���|��N� �xB Y�.�}�l���8t(�L9�r�^tu�_W��F� ���A��ΐ<	�N���		 ��Hn���.�c�.�����E�L	�ĵ���6��&��K �4M��"S9�Á̑�މ�$��hC����b����|���h��q4ɑ��hO��5<]-��ϣ�׳�Mmyt$����`[l�L�%���� ��������O��:@�\��I�doKG�D�X���do�.c��މ����]o9��=�Zb9u�1ڽ��O��q�&TV	�ES��������2d��:C��>~�WJD�D6M��Y��5��+��e����њ�\Xf����\�F�َ1RY�j�8�I��K��-f�tp�i[	b0��P�M��P�R��m�&-�=e�0�v,t&�L�$�(�5���5�����X$\�`�kD�&�q,�Ɍ�a*�:nڑE��e�D9	r؂�;ea�0q1�)6ю���eHh=����|4�?�fc�LhR*�-6�*�8�,(Yab(������{�1v�{��E=�\DA�n5=�`I]� �=���^�Ja�B�jAwC�!�.d�_�<Ƈ�KȺ<C�&��@V��[#���)�צ,4�l�w�{�1 �N�DK�|���m �=���@+7��]9��2��6�& k٘�N����*�T؂@ ��"��8[ga��t�"&�藗�s�*=��^�r�v�%��@d8H�$0wC�Y}F��5�;�� ��/.���W�w�|���c�FA���|bw���$��� C%��@�e���~[U�b�˨>�m�̅����6�f!6��f�(չ�M
�sg��������0�ed$����pOY2	 �>͖s�P � �  ^�a��Ô��d�d���X�z����Ew<H
��������v���x��Wc>\Om����"�:�ߏ�-VNk꛽˅1N)�wo}�������W��
��Qg�to�g%%�RYe%�P�=�^��P{�!�z��@,}~������p<����Es��	 ��țH�z	��c���{,@�H3SDy�B��@ ���~p��wΪ�{��g� �d����-��I �޸�l4�M=���'��#��/qŐ�ܨ�
Ex��2d��$��g��/xGK�z�F2	��fX�����u�ښ^����Ø�"�:��MaKv��P�]�0V�C'6����\[�c3 ��r�!�>�v��I��g���lS�MQ��hb�Kw�C�vw����O��5D݂�7ь�SkC<�1K���V+�����>�@�%�}�`d(�g�"�����e=j)鋈�5N������Ļ�j��z^�"+�Sz���n)�ft{|[{�Cz��~"`h,[�Ͷ�о3&�@k��N�����s�����?"�̫6�ѫY`oz:=lH{�>�8��������ɮx��s���\��C�A������#kf���M|3xA���Wf����ɸ�]ܮo��kУ�kz��;� {��v������5��3$����c4��Gʌ�l:����׳�Lٓ��#y�}���}ѝjj�'Y_�_k=�Ӎ�n�7]�vyr~X��ZUٮ����,vJ�@=ꦞgW�z����O����r�G^��(�➁N=�U�T�����<����oOW��6f�^0枞�!�)񣯍X�^�`�Jv��;���a�ݽ�;�w�M=��@�Of�y�T0d�lg������c쓽���{YŮw��-I&���j>��Q��I�÷���b��*3�
h���Ud��~�}{Oi���:Ħ���W���;��W�=�_�~ǖU��z����� ��bCO��7�|� K�b�={G|��%�񽐜ٕ�ݛα�4U�'��g*�����a�_��������/ft@͗d:	J0�ӏ�b��q��Rd-�u (q��Ϸ|�(�V���!�h��|��Lx%���/�^2R��\��=��Fs�[b d5?yb}׶��}1�||�'�;�{���$K�OP����S*͍ut�O����s�r���l`�eC�gW���@R�[5�H���[�2���m��?L��x��||||||~?_����L��ffzϿ��R�e�m����2c��F�X��Z�y��e�[g��Ϸ���������������x����ffs33�}y�V�&:5�
�j���[=�y*Oo���W���o��>>>>>>>?�׌����fg���Zl�q��c1�j�+�I�V�G�Kz�)l��Y�����z��e|~>>>>>>?�׌����fg���56�򖖻j�PR[X�ҥT�3"8�qr�UQ	S��P�(��1���b[*(�Qy�֪BVH�PX�Pmbőeh하�b�n�)���ID�FQ��eTZ�i�9L���-T��t�DC�qՕ���O2�l�b"%K[[�,1Y��b(԰b
DV,iKor�j)Q�[Vw��!�יW,�iF�`q��A�QJ������K,���K,���㤂X�[n @0�s��H�'�.�Q(
3�}���� i��w�}jDk����;�����}���]���6��g^&�.ِ$�{2"�'<�'�kg����n�wve��s��t����7,�r���N��V(�̬G,X8m���0���5�3�i�9�c͓v{�4ƂA���I����=���4l�]ݑ$�ǳ5�#�����L�F�D��P��o�H4yp$�w*:��<˙�$hE�y�X$muα�@&z9�|�S�#�:{׃�[FOD;�$� �&��2CI��A&����N�����髕CY���$g<�,-�#j{QO�t^H�2o<?:�����	6$����E�4�����Pu�,;/	��\��6��Rm���Rm�n*c{����ON�U��h��Ocw��Nb	w�q\_���fgĲ�K,���K,��=�|���:|�w�p↯&�%���ǂ�(��7���I0��fK'gd�:Cyןt���K���c�xS<0Pw%�d �Kmj�G6Sah[x�,��<�U��V+ө�/�,��Ӣ��-���Hf�" �Yڰw���$�R|y�J�M��<ԩ�D�v=~�c7��(�:�w�b�D������{��	�s�fA҃�C%����b�gQ5�ND���`�I��T	�]�$%���נ�x�pH�s��Ņ�� �F�@����z�:ud{^�����WyU� >P�'=1�1 �g�����p3�k���kf��@�y�E?��xu#�ϝ �u�r/π��6!\��.O@�'. �@%��;�
��V�*6��!���>�=?eU�N�(Z�}"[V���o��������O~�7�H	�oBn�3⦤s��bә�͵��ϧ��K,���K,��K�-5���V�q�6+˿��v�N����V�r1l+i���*2:�a������2d� \UuP�yL���v�К�l3Uѯ[�] ��]m���#0j�:L�u���y�Z�\�,xۣo�Ё�xG:�cK�6]4U�ʐ��fm�2��-�f���3�%(�
�i���:;�)�K�r��3�o�/:_} v�nN�ʈ�2�Һ���fЬ���y=%�l�o����g.�����u�?L��y�>���s��Ta�_��x���}�ݰ!�w�Y×�Eҷ�,����g��??�%��'ה(�@���q�>��㔲�`��:�@w0�!�
;0��JYveT�$Y��WP��.Iө�P4ɏd&0q��p5tĘ��$�r�U���jsn�T�d�ZS�<���v���� �ƻ���
�)�����L�W�
a��x�T���W�D�ƻ�t��혔��`����!{��Q�=����Q{�~��=�E�3��4��([�QXn��smѤY�w�	P�tb)�'����e� ���8l�	L�=� KO`$žw�*�L{�r���Ò<��p$e��ȗ(�=�tEk�q�=<fѺ�7Y-5���]��-�n���->Zn��M���09¨O���G�j�$����4$�x3�2�2�2&^�q� Bm���;��ɔ�FWy��!�-��fAg^�%����ڎ�������,i��ܼ5��d��׭$��H�0o!�V������)�L?��W�芏)�9�$S�vH; s^��$}\�ﴟmo@�R�K�T�/��O��P)1MK�P �}��x���R%wT�����<�ށ���sϳn=�pE�T(j�Up��-�G]�A)Rb�nL�SK��x{٣;��m��v��)��C�y_~v|璅��۸��ށ�_�����O@���� �7��;ȧ�p��Ao?6"�U���@ ��+��c5����K}�@��DwƟ�+����{$�H8��4X��ƻa�B0�w���H�@z�r���������K�V%2��=������;7����nr�s��������c
�Ax��x�ǙIY^��ډ�ijd2d2d̙2m���I&��)��r���M"}��_��~ڙ΍�{�����d�n|����5��O�+��� S%��q"@1�;(�D�cXd��a�*<��$�g���l��U�%�l;��y2
���z���E�����x�	r�1c@�(������sU+��U]H��r&��⬽Q�4�#\�h:*.�$�}��ZS���W����˒�xw^�)����a���w1� �s�L�@��_��˟X��$g8�H��� ن����q�}oF�)�9)�*Z��<���otx�d�5�
�=����fAئ��%��	�a9y�PD����f:��Uʽ؉�xbA ���Wf�ڐ���o<�O@�������w�(���P���c�G�yr��<����{#���>��^�3��ǨC���z��WW/l�h矣���At$��$��L؟�g]�_�ދ���i ���de�l8�T�\a㿸��wz�'v�*��ї�o��к�{o$8��2a����'5��q���ɀJ*ixU�>A���Z"��5[�?�ԲYe��),����<��&���w!��B�lE��}�0���b.gl�.��b:�rڨ�'o�CnOV(x�w�υ��흉��*��nk�v���#�1�l��$��sdZt���~/e<ng����V�7l�жA {��xS�d�rA�oE��Z�8���E����rA�� ���q I2�Ӻ����"c���,O�.q��� bq�~}|3W~d�\��;������\�!�� �$��]��$9q���W^H�C �y�;O!�w���w:�'}`c溾��;�,���8�FlD�F��dPS�xn��#)�_R3��]<�(225�&=�p�]fʏ0H�y)���MM@Pv9ܜ� p�j:��ς�]����ZO��w��w@�)��o3�����*dnZ=�x�)�1���C.����Y>������z��*PR��]&��eQJ�Ϲם�N粁e��YIe�3�q�k5�*Rэ�(�*�¶����f1��F�Ű�����ۊ鶚[�!�Y�ѕ��j�a��f4PȒ�!��K��sqcB�ts����t,��a4�ɥ�Y]lH���N�*�u��b�,�ؓj�A��0f�˶��T�XW�ap�������3e�4��s[cdn��Eia�tY�[�2�-��SWBd�p������ѥ�Xx����.���S��ҋeH%a���% ^�n��7��̉-G��3�T� ��,�b��P�Iު�hǼ#O%��=Y|���E��9w��"+��yv�dX�OU7��8��2y�"!������W����'қ��n�S�_�ܑ-o��bgE�nH4�T���
�widA�K/W�;�s�[lD�6��2Y� &�qz�Ax�!���R�~��=�Y��	=��E�8L�ݛ�/����o�Ts�l9)K�����x1Ti�bI+��):�ME�FV�gk�l���A3�c$������U�^:^0R��sd�xxxIJ�k����R����E�Dc���;��|ԥ�1�~�m��`�)|�[����\fC��Sr7D��z�ʌ�o{�@53��6�=���,t�MUL�;�Y1�2�P��~G_מ�nS`���@��y����D�����D9DX*���1�o.�D�������JP���%��}�v�}�R�K,�Ye%�P;�}�Y��Ȗ <ɹu��F<6}}9��B 7�;M×xObG���5	)�V\P�1���*������#��o�Snt��#6�e����9E@�L���t%��&t"u���O�L���zם�+3��u��k?]GB�D ��+��Q${����[s��VG���6,� G���̀�B �ށ�&,�Σ4_?/|�~�Ͻ�~f��Φ�]���
����5ұ��s����x�x3'kQw�\'�\���x�$�tL7A ��_ē�<�u��k�4�)�]kB����F��eև��(_�K�Ģ�=�/C��A8� �I�A.�i1]oì�L`�o^��B�I�~��'̑��AY���Ɏ��w��j��;��M�M���j\b�2�����>��,ZjD��f���?/=�2�ʽf�R�3oy�O��줲�K,�Ye���뽝ǹs���kA�|�����������'�0Ew}��iw�/5������n%$w��l�q6+��OЉ�Fp T�=��cQP*��6)� ��s��2uӋF���b���L�_t1h����e����i��3�פ=	���ޚ!$��(�Q�ڹ"Ls5����4e�B��L�W,���(��=�c�(Sx�* �Y �-��e� ��2H^gC̼�ƹ���5k���&bo`P�� ����e�o��I�E�&�5��w�clϧ���+Y2��wUT[;� Wt0�&󁹠G��k�@���pS�������� 2it7�|�I�fA�jX�A�l���	��
��r:H�.���C��~K3A^e�u 3'ݲ(,���٩Q��}�{�h����9O0=�c�������p��n�O?��i]f�Oz�~��>�`�z瓶��I9mǏ����4ω�줲��),���H<��oy��	��j�O��w�s�K�οwSDn�d��c$�e��<k�&@��"w���OB�<G���L���l1��m�Qс���0�4q�g.�\��4W�Y�"bZB��x:J�o]��!{�L@�I"���������O2J��o2��i�,_D%�yw��D����e
[��8��h�z�Q; ��4]�"�s�Ɓ�dXs����37���A�C���4b�gGY-���>3�ލ��7�1��Yǉl���"k�djX�N�Z໧��Q��O|C�����X�/B �I���+���G_H��6�U��qx��
b��X�a�>fp��:H�&ݼ��t���sf}���b��2��q���L{6 C9�ť�!AƧ�naS���DD{��\N�f��;��ܠ//x�	�k�a�}�����Y�ꚪםn�HN�T���k��y����Ba]��J���sW� 5 '[sҢ��[�����'��T)���
4.��o�����u�j��l��V�S|t�U��S�i�&��zI���|�[}VV+| �3�����q�u
ҕx�*��<��MD�W���`P[���7�hF[��^�[lƛ��ۻ���'x�@�u��ݥ��*�y*��Bx-����h�����~�MB�,��t�@�Z׾j YG�p�d<��9��X6]��^:�Q���uW���#�7��=��\�)k�گk}�zZ����o�L��J[f��8p5���8f����7RH3w7�yK�:N>��j�{r����ϟ�섞���J��<}�k�j�_{F�R]��������]�ㅔ�����d�8�K��'d��`ڀ�9=�$�L��f������Pn/4n�ԝަ�.�0B��|�Y��{�������p�p�����S/���-���.l�㣊��74�y!����	��ˈ��z�h�ڑ���P�Ő����Y�҆�ʆ:�)���N� =/lEM8%� 7��Q�)? M�A�JC��{�O�
ۮA�t�3_	�d�LU����^���5���/�h���e�	AC�M�S(��72�X�����qJ������<�J��~�_����~>>>>>>3��+333>ٙ�33:O�m���E�.e5n
�X^��.�1�Qu�E�6n|||~��?���fffg�3=ffg>����O�/�y^Y疒�R�l�R(�]�Z1��o����~?�������fg������ߞ��=�_��I�6��l��E(�mm�-hU�R���j�oXUʴX����ɟ���������Ϗ�ffff~3K<�O'�ɩǈ��CJ�oL��9#���(��2�vO2�c��`ԪV(V��(�z�V4��֣3
"��,.�0�1ۀlLp���C�s���ZV'30��D�,F��dU�S��N!S�۔������0m�kJ��FV���T���J�Z�ڭaU�$�2P����b'-�f[nL�)mJ�jt�&T�C�Q+KK+c�c1-���r�+Kz�nJˈ���*Q[J«ֳ,��ۉ�-+���%Y)+�ol���-������XX�Y|��qv�Q�	�֮��Yu�?X�,:�&��ˈu>���q�n���h��X�LAF��=�y�(/�5&�� �VA�A��KvB[5MV.� %@phƍ�H�4f��2��v ���[C`ҳi����t��A�"s��gj���L���J�tѴ���+��SR�̈�mT�d(].&�F�^�2��=H5hT�F���4&�"[*��s�[�\�`���
ֺ�i�XCK%��Q���](�j`��E�l���Ȇ��W�
1]���\�q4nݭ�.4j��\�Xu����lW��D%�8�)��t2�q���W+]Yh�͂�u�S E���X6�L�[y�M��)�Ü�#E����aF-����qZ��6����v����ل���Z;kF�e؛��֭�!c�n��	G�L.�I��V���,��rٛhFfkmҺ6N5u�г
��-�X]Ƅf&Mf�p%�p1&��-�a3s���%��j�G��ΰ-����d�2&��qa�#�q�2�Ҙ�ˠG�6�-�j2ǋ�yX҃0L;D���6������H�7
b�ΗT��.��X��eH2�n:䦸5��k�Z"�).���3f���q���bh+\��,���v�݋AiA��5Zm+EF�vs�j�tH���թvj2�upgF�8�o\*R�YYf���i�-ãIXͺ���SZ#5����.6�Zܮvh��Xl-nG�i	��3.�l�`k0�\����&Aq��U�Ѻ<�qF�ȕ�ـK�ڙ��YZ�FlnkqPF5m���fa�U��A-i�\�F��׺�4ҩc���v'_���n������$�%Z�l�f�2�lMU�,���Sν,	���f.vu�KX�e����Ќm�JGXژI��Z;��a:&�K�`���̻�M\F"�~%���nIA�gj&7�b+j�K�VjҖ�_zÜN��ܲYe%�XY`k��[��7�"A�"��3:�ZYv	kbg)��	t�&r���-&��K.�� �4\��ù��hE�е4R-Y�kc��m�Ǔ2�v�(i����L��&Ֆ�̼茺f�AK
����ɜZ� �!����.�a���V�&��B��ᖙ4�M���`��$M�������-X��6�]Vd�ڑ�P����w��ybZk�d@�x0���Ij�b.���ٮ�X�:�|��o�\~߮3�y��cg�n�$�a� ot@3q��k{ت+�16y�u�	����2�C;�p�9 �t�
�#���h�����8H�'�Ltm�I�����۴�Vzod�����vH_4�*!%b?�"�������8�=���̢����'X�RvL��M�����(:����u���JQ�A ���A!�0M�g�dy�&{c�(z��FR��SC�wP�ө�.��Cà�X��^��p6��N�l�đ�Κc�E�CkKKW<�^�dm�|�8V�Ɉ?�' ���^1M�@cjWh�R-e4�Ρ�p�������p����~�G�{��S!�c�����fH�)ҵ^����-޽h�Sc+�>[
 �s,=
a����C�?�@�Q���S1������:k���g�ʱ��%F�o�=A�_f�r�����њ��y�i�z[�h��׫O�����F,ŋ	�Dc�;r!��J���$�Zu�z\�a������1�l:J��^;2�-"�y�9��m�A�ʭ�Mv�����ԁ7���ظԇ ��n�w��15��:/=�8�d�9�Ib�"�W �1�� ; �7��低��GMf��Ǧ�9�U��?�A�(�@k�n�����!\vG�-V�©�m�L�(b�"�j� @��Z�؝�ƻ��A�t�\]��L*��Ԅ�+�"ẀY%���M5���n QqO�AN���<��)�ż��HגA�@n��V���yb��YS�0��@ 'k��4�q�D̤�{ޚ��C� ^���̫Ȅ�1 �mt�$���P�uV�u/oK�״��x��a�Hv��y��A�ȐZX�J���PuR�����/��v���$/�Kx��|�{U+�|%��Gf��FN6�F0��'$�����f�4�xX|N�#1#Nf�:Yس��[� L�\�=�/�l:J5)�h��V�Gu� H0�2���(s�%Jy��׆y��bpk�~cd����q脔A��|���X�I��8�i˚w��c��km�O��4�ȂNoy�������#���b������ٛ׊�Z\�ܙc��o	��"�ɲ��%��[�5k��H���P����̂6�$�#��N���[�X
6��A2ݻ H+$��)��:�i�e�ɤC�������`Kb�	�$��ZY	5��{)?P�[��v2�"%��Dl�v=y�����q-p�����ky=2<�1�k(� �a�p��Ø��{�W�4ڳ,��ȓ�G��47w@�]�S�Ҹ��*8�*z-M�z����;]�1����6���^J��6&7��o{Ko^c�3+ח}�e�����h�MD�db �c����[��pW�-�:�|qlN���n�O��P�c5UDS ����4�;d�[q�=���̑�LU�R�Gqu�Im��3�f5t�GF�V������嶯k/7s��IDB#���m���q�=mْ9�&��<g����0��ՠL��*3�{�%��]��)ʇ�@ki�Gr�}�]��+U��K ,%�k�A������ LR����	h��'h�S��uX�
69�I ����$e���ft�{|	&/�c;?�,n6(�m~��y i�뤌	玌��������Z���4�	��ꩭ�Vz��tlw���8� s='�^�#�ד�L�G_S�NS`���5�UK{}� �	�zg��=
���N���[�ϕ����E��ɃX ��!Oӻp����P��^w�}�)�wԁ�z�9>-�0�@���~'Q��^�~������X�����DX].�!�������8�̦�Y��+�6((�T��W���ÃK�u��n�3é��	bò�sC`��m�ㅚ�kju����K�ml	tr�ȱ�l�f�.� ���^gJm���y�L�Є�\�1�Sv6L� �¬6�h �6�i-�+13B��q��W"YH���ǡ(�ۂ͛j�[�J�hh%Z�;ejQ��u�Co'�?��MmGP�n=	�ׇd�%�Y�����8�JՑD�l�u��G�>�)�\:J"�����v���c���|���"<��BΊI[P�z�-V�ڞl�;�Qٮ���C��>��9. ���\1�.��_��qM/0�3ݒ	^�LYX$���ކ�Awy�	D�]���n'U�eO�o /���{P�� ����K��0�&\A#w�n�$dkS]��L�E�@̈O�X;�Nz @2�S��� �kz1�A۬e���VLr�a��ʺ�0f��8�l��è�u��Gf���
$=ߍ��� ��y��W�MnĽ3�%���dۉ��RbC�n��hD����f�������c��]q�Q7R��W�?��_��[rr��c=��׽2��0��qR�����
�Ć=ј9OWP�4��&�)��%;��I	�V�f��,a�Ča����eQ�^����&7ٵS|�=���R���(�Tk����D�`$���F�H���+��w�2�ە���vH�$��D��X��Jr�᪁]ϝ��y��2��\DI	�v�"dy�%���5��XǢ��A�Q�$��A��EC~{nd��<����*�� h@P<ɻX�� �g�;l?��\��}}���r�VjP��;���r�.���UK[��X[+2�'hI�lݨڔ�&�eO6�c�Iϓ�$�hg��bG�;�������5�Kn^Ц�C5�%�/M�'�	�D
�z%���WذL���Y�[/���-�kiQ>4�p
6�_�w�NR�S$�je�3~j��� �p���B{��#�z�'���|H�ӻ.��|��d�:g���`��r�p^������zE���P崆,H/�����db@�������L���g��6�����YJ���{���/�\��v�~L�Aw�{vA��Q���C�-<����C��w<��I��	�=��;�	L��X��1��}2�����%����;��]�B3\h���PMGj�鮬��ʠcJ�/�Ӗ�~���^���	A�K[o�I�G��wa��Q$[ws������H}��x4&J�fZ��|�	�GZ�ߞ8BeM�ޠA���O��)n�ʀm��������g�=N�����g;M�Xo�O���燃���%M��4!&�I���'�cT;�!"sw�*�Z��	�P*����◻7�KF�l���	�I۸@����K�j3u�H:z���c)�}��+�=�r��0��
]��º��w��w��7�:�p+<2�Sdc$�3�j21#a;�������;�����P��P7�`�R�w5	�-dٻ���˓����#�22D��ԟ�s�}wx��w���۴k���1k\-3v�f�5��,161��$�E�֣q�I��A0
�����]c�e;�!����NV���s �A{��T�b���4�q��S�bٜ��(��ȐI��mi�����w��68F�4s��D�����,�n؜�f��i���ʘ��%�X��e
���!���N���Nꮝ��;ތ�-��m:��'"��"G��(S���T�V��!�$�K;2Fs�Ɓؑ���ڿ\C������	�P(6)�\e#(I�6wUP�A��M"A�G?4�"�̄j�u�Iy
k�S7��&L䇤�^����Ɂ��y���^��������fު����f�{n\�����O��@c#1 �w��(�Ҵڊ�s4?<<�
�f`�F\3�4j�&RR�60�)6`K�Z!`�q��p^�c�WD�g���k��5��HbWu�f�b+���1�Vm���p6܋1!����D"J�8�,��$f�(���|B_�q2��lՋ]r�!��A��q�͍�v��R���:�hAc7SZSj��0�z9����w���b���v�WX�K"��k1sM.�Xf��y��QĬz�\D:��t\ύl��zDS.gD�{0���h�!��{2ı�J�����)�;Ďo+���e��J$��آG2E|�Ǚ#�t(%���7 �`�������J'76$A$�o4�,Z��q,�{��52�A>��&%��]�xa�ܜ�f�홁��³�l?���0j�*H��ؘ�I�l�	��$,��I����$�D k=���� 
'
uM 'o�]w�{�^��X��yTH$r�(`Y sc�ck0��z��rRN��w�g�u���5,ta.�j� ��6�<?�m!�k)]ӡsc�
�NJ���5��&i]�r	4��	�`wwS��an��1ַ�Bs<R���C�7��}2H>{:q����@�eMF^��v-�m������yt`��0�fz��L���2l��Z�lDXR��p�0�z��λ������@c�I�u��}73�����H���1Z��mvI��ǢլsP
s�T��i�2C:r&��^���u���ݨ�18��$��x=��9��H>ݵ��U|	�VUN2G��2RPY��A�q8����%քN �ۓ��RΙ�	$��ַ���P��MS8�ݙ"UwH�~��,Y`9[�����N�Y���w5ip�)5���4m�-�e���'��;z����A�CW��'x)9��6^8 ��I_lI#Y&'���z�r�z`�׽�F���72fu!�/�a9*7��ZE[����n<9�)�mf���#�@3��<q_9�(V[�8�䔽8."N,�"�;:ke}�!�hh���s�x���Ҹ󏺣;�^�N��<.�==���>{���]�Q�w��A<}i7u�^�4��Y���UZ��V�`���V���%��-F�J��.�=y�(��{+	�^�A�<2�RF�<�PŖ^=��(��w`��/��P�wt�Q3����Z��ـ�ǽuq7�OH�חg��N�]���{Okk�,��ӽ����=q��MHx��z��5��ݩ�ﶾ{�4^�jﲞ·{G��緢�K���`�����zn��x���gX=�}�<��7���d<y��{�)��]W��0x�������Gw���3}5u������G�6X} �Vn�[��K�����[<�W����
o[!k����}����u>믆p\��F��I �=猄�K��Z;�$8�no!�Y$/����y��W�7w^o���U��
�{�G�c��x�37f����A����a��yzo@���o��=�N_f���Mس���d7{�x�Y;�G�改�ޝi\���׉S�l87!���z=.�\W�y�̎��!]�������r�����}�g['�p��L�Ss�ꠛ�CW4s�fIpfj���w8��0�-�n����&�س�r������ً�� ��$�c�o�H|s��3���,ONߘ�!�B��cL��.%%����~s���F5�i�4�ë�{�5���S=F�Zҷ�U*b ��ح��b⭾R�DB�1\b[��7�X��j*�h�w;�O�����������|~�3333�Y��y<�MM�)l�����\�������D>��k8e2Z�Z�ҍkSS����zN�S���w;��'�Ffffg�3�ffs���,z��F�h��m��!�o�����kqʺˋ
�JZ#RK @����);cc[cho7������߯֌�����g�����ߞKK�LjgY�
h�HU-��*��M[+K��Q)噊����������������h�����fx���}}��ye�[e�>��&�LWL.R)Z�T��W�*���.��hڶ�+ۚ։��nV�0�R҈��Tj�,����S؉n�KY�2�ANwf����5Z��m�g�D��d��mne��"+i�P�]j�Qn��4�؝S\N4`9J���q�+e��%m*�˔kjx�j6ʫ�I�Tt1���(���P&f66����YJ�-�-2�n����JH�3��`��S^\��ڥd��)j�挸e�d�@bF 1��u�����ϵ�!�%�w?�����w�$�'�ـ���G�����c:m}�)�7��n&i�iMݒ[��	8��zs	B_:��خ�;��Tn��$��
�y��>2Q0��IZ�`�zy_�G��G��8�dt�R��cB�t��i��e�B�4���\���b���2�����M�Y�E�����i@�eܴ�>���K���站�g�p��)ڈ�)d=zb!;��8� �t���`MÓ9�f�(z�^��-�lg� w?��{A>.h.���b9���@�cנ���HE����T-����$w��c5��2��ē���y��[�]{/���fh�!�3�>�Y�d���R�h��Z���<�
����r1&n^��/n<h3��t!w}-ٓmqg��&��[��^(t�3]��`c&=7��y10c#4ɒ�x#1:q9�xB��.�I0���G�'}��k$�7�9��D>;�idz:d�;1Pt��*1�$��#	�0eQ��Hp��)^t������^4R[å�;ØJ��b�� �A�Y��ݱ�f��F
�?8,u�φ�����|��Eڨ8��$�v'���݈�\i���7{��� �Լ��j��*#��7�ɀ�$rNy������KQ�W�9�����Z�̷7��'/��Z�<8P*�6v=>��m(��A�]�Neܲ����|⚣3�X�/�fm�*����R+��%��iW��<� �{ʛ�����`��^|ީi��t���l���4z�c�<�&��a�;?���:{}���i%��#��S�N�/4���N�Ǐ��X�z���.�鸃�B�����u����KB]R5��3LL�sn������3&�h���[�V[��h;8�#\1[�t��u��h�u�tŤ����Rhqڱ�+����L�f��- c$v#5ėb�6��Hk0R=�hU�U��ˊdڽNt��L�6�X%��M�9.\j1�Q�ԥ����J�2�!7b�k��M��lՖa�2]t�(����II׫]v�<���	׭6���i�X�XŖ�f��S��6����ۮ����q�=���@e{b��OK��e�m��y�Lb���e���'�0����S=��>�ݓ�.�i��,F7�7�0�1 �M�����8��)����6��e�
)�dtbA���	c_���Խ��"��Y�'����7�F:�u�R���{�I�0u�u�-LQ ��O�2C���D+��;b���
���)��
�Q�$ϭ�B�1�Pd핎��h�@�>�\1��b�t�O{���⻼%ɬ���d��X���ajmZe������fck.S�ɲ#"x�N�y�m�ʿI�H�$
��Y)d�g?jUw��(�.�d�P7�Z{*�:qa9P�TH`���T1�}(�<-�O�mß"qF�Iw}�ދ/��{�o��qW�����la���"*��H>e���{aD�bN���7����Kf�鯶(��VDc���w�|��k	�F�aӁ[:N�BN�Q}�A�^�%�gMgQ��tR�W���&2�dF� �	��ڠ�Q�A3m����7��z�{�g���l��H�tX�$_d
c,k7�������MnS&]sE;E�9���8��.!�={q ��W�[v=S6���}�i��h$_oL�U/���c��H��VX��u��V��k1�X�6r�vu��{�g3O��v���<5�eNf�cl��e�J�E&��}=���:�)�*�`s<���<?a�e�[e�/��'�j����+yVج��H��IvC;��Ys8\�Ț�.6=9w��m��:q�](x�I���-Q�B�tP%�/^��8�N���{=7��yhծ�{}J�����J�nX�*j���>�x��C�[�����wZ�kc�w�U�O�ȁ���Z�a�z�lb�w�)2QC,�I�I�]�n��Geߦ�c�y�hvrv^UIo�u:���A�� �&w��m;pQ�I+�x�]�A������~�׶��<@�.H���D�+gz`��򗭾hp;gj�)�޿+$DA�l4,�n�2�h��-(+�W�K�J�����vc��h8b!'��%>DH;{�$�&$s�A��<dM�r$H��$OG�B��S;������W�H=>:&p�\�	�,���(�Eo8��Go:�]{Ѹ��M�{��*"��{��ȊH��$׽�����Aq��l��nS�]�=�1��8�](x���p�׼����A���$��Pވv>ez��GG{r��<�W��&Ľc@�{2b�en�^F��
��u\�S�������4"��� ���cA������8#��������M��8q�;�h_<נU H�[��y�C(�;u;��D�,;�r�T%�]�,v��3�۬V8��Ζ5���sn�������w���L��yeL�A-�="X�I;q��1�Ӓ��^�q3�O���p`9�����>]�T�'ŀ��G6+�@�Ip޻�dȲDgt�g�p��y�d�v&4+��4"�� �;�����A��+��پ~9<���U����������t'�py�TD*��sWb^U+э�Ft��ă����y��R�}��9\lTp14��ͲK��$z{�E҇�j��]��H$���N�^S����6��츒D2[�����&�W��y��b�ߺ�yRR��ȨN��H3>���:ѝ�k��ˇ���@�1WyY)�0x_�{�dDa��8 �Ց���y1�`F$�}����[i�bh�.����d6���-�0�۹�aJ��؛T`9�4%�F�3	3BWcG�4.[T*��m"��e�`�eīn!1���&��ė�pMͽ5$�栰�×q�Ԉ��"�Q�KY��6f0a�pl2A�k5�����5��t:+/-��3�2��#��c��vI�6%�/h�v�.�V������=�6u�[Jh�a�k�"��o*�q]m+�|�� ������]h��a�O��b��+����b2�$�tb�(��������DCċ́����v8�@r~����[����@ʘop?�Lsǝ�LW����H�Hg�����d�_�^ɝ
�΂d^��'�0p9�� _vĀI�ɏZ�nn�[�`�ޙ�H{�T�"��0(P<��]<vT5��ئ �ȷu�	j���ޮ}��'�A>��TD)͎��s�˘��t��X�n;�:S`���I gn̙(���[�>�]^�Qs�1B�;��L��q��Ķb�̴�04���a<6k��x�UM;��kIӃ�Q8g���|�,�tI$�#��s@!N�i�ŵ���1$��ɐH�uBz�+{ �y����S/�O�P����n���<�.r>��U�oo?
�sS�)Y���O��O�[��o׻��s�U{hF.�\�bŋ ��\h$��hƁ��q(�{���V�7�=q����n����(�v-�6�L�,=y�N��76�a/z���$W{�{��d���͔�x��ho���o�г���O�Ab5�/���J��`�8��ݩ�"5�����9�qǑHC�;�'�A'{)i�x�8ȁ���rI1uլS["}��[���	����K9�>0���/��C��N�S���:�Z�fj˦���G����zy�)e���3}\�V���6�E2kޑ��� ��嫌�����$�'�"9��.�r���Ý�["�<�35	Y/'��x�{�kjg��A ��C��D[���v<�XD^܂퀺���G�]�0I�˘�da�ዜ��M�{��<W�z.��"�cz�J:��˅�^.��3��7Kّxg�+���Ksf/m;o����ߩ[eF�����],�.�eK�9���fhT��-�e��41�s�bss4S�~%D���:O�������O9�$�g�w-隈�Uw�Z@�����|r�s!W����>0A��4�����s;��[-���'!��p� �"/-o�C�I�c��Ա��.Z��-�k1�-�M��,m��-�ZV�ӆ��h�!� ��l{fH�I�os��eD��L���9_�u�k��5�q�N�����R޸�I~�5����9�Y28��"A&��Ay���{Us�ӃQQR���@'���m��>y�-��Ln�{�ı)!5��IuBy�����,�ŭ���׃�"#:�&s��c5lQt�Gm����s���+�+��3�n�/�k�/���e��M����n����؁��D��20bF �:��i�u�O^�;n1}%i�n��j���)��޼&d�1��D�M]� }`���wO4�1���Ѻ��y=��K4ߕ����X0��EY�cCR03De��������x���b٩Ru�d4���0���E��� u�v1��3,g�fƁ-�SM,��D42�8���9�<Ǜx�x���P4_��52!I ��Q �{�	�#�!��]tƉ�=��a�����k. A���O��p�3��g�h���zd�����h�L������(���Q�|irl{��pm�O\�c�^  $M���b\��m�d�DD,�K�I�{��b�˷ �gʨs^�Q�*I0�Od��p�������;7��� 0�������s�/$D��I ���0�I
f�]JE�JI�  $HD� X�X�1	 A��c  �ȒŐ*��VB%Ij�bI�� D�!	Ȑ��"1 	�H�A�@�eR,Y"�X��-XjةlZ�
��*Ֆ,@�,X�bB1��-YV$U�jʲ%Ij�($"E�H�X�X� ŀ� �$�1H�X��H� �d#$RXJ��ȱ%�E"ت�R,I��`D��I# B0��! !"�B0��!" !" !�!�
,�"ĖE��bK"�ȱ%�E�%I,�,�"YD��`FH�HFH�A,�(�(�*IdX�Ȱ�� !�!Ȱ�,�dQdT�ȢȰD��D�9�h$� !,�,��Yȱ%�E�d# B0 $# B$"H�HF �a#$B0#$B B!#$B0$�(�,IdT�Ȩ�E 0"@B0"B2D"@B$# B$# B@B$# B$#!��! !!" ! !!�! !� !� !�!A��	���� �`D��d�F �H@Bd$�$2�%�	d�$��H��@�@�HA$!�$ F!��	����P�d��K$RBY"�K$XBY"�K${�A<�)	�	H�H F@�@�� �	��# H!�H�!,�a	��#�BY"�,�bBY"Ą�E�H D	 �H	 �H�FKU��K$RBy�ybK���H��,Id�H� )��E"�d��DHA��@D�BA���30	��B1#	!�F �HBA�H$a%�@��D�HHR2$P��E"���$P�H��$D�! H�D�H� Z��Bň� �"1 �ŋ2 a) ��� �$�*KVA%�VUI"U�Uj������Y>�,�O��?�$�D�@D��@ 0��a}���o�������O�'�O�#���?��F����?�����X$߷��v?
�#���H�@�	�r������BH�C��Y!$�������O�g�H�'��j�?�?�O��i?�$�$����'������I�_?���O�?������������-�j�$H��KX�T���%H,�XIb�E�,"�X$@$H$�A�# H! H	$@BA�!��$		� ¥I,��X��$�bK$	�!H	"@bdH��" ��PHB Ad� E	 B%���H�Yd����KR	d�A*������ �$!A��	,Y�%$�RT"X�%I,��D�aD�Q@��E�$�I)�*AbIR$��
!KR,AbIb
E�,�O�$D���R"�w������_�����y�	hI-�D�[$�$�B"_����O��_��_�Kd����t�$�	��_����"I�?����s��?����S��"��,��O����'O���?�IHO�I��������"$�?�I$�?ړ���?��_�'Od�H})?�=���$�O @��?�
�ԟ�8M���P����ǐ��pa��tp��0 I#�g�O�����?�O���]$�$��~��O|�|���a៊��~�#4�� ? ����_� I i���Y������$I �I��'O��;��XY=7���� hw�P������&��w�0��� �I�pa����,���'���{'��|?��ߧ�	"I��C��H ����??n��B��H��d�Mea �<
[f�A@��̟\���0 4�  

@
  �@�P��E�  ) >�[ d@�@ � 
��\  &��J�کJ$�T�c
�Q���5"m�VU*UQ[[a*P��J���(�BR�l�ET��+f�JҖ�JZҢm�`|           @  
            �             P    ��=� v^��@ � k j�f� o`{ښy��r � ��3` dc�TT)T֪�   ���p\Ɣ�(ׯ �@��@.`.� �)J^��`
J�' �4���
q ��� r� n`iJR��QTC�B�    �       � GN�
P]��p
<@B��AJ^�@ �R Ҕ�����.a�y�`x����y y� p҃#�@�U�5��*/    8@=D2 s� �C��\�
����P����4:�� �,�JDf<��V��J�G�  �  � P    �ʥ\�ݔ�q5I���s4({� ����XP��f���	zqB�� �J��������AD��S� � ��y�
g �B��:�B�+z�����nc!N[��&u�B��� 4퓐 ��RQ(�5[� �    (   ��de�#�-'@���� �d:�v(��� k��C{ ���ƪ�i5�R�   �@L@o[. t(͎��G 9 �,�V ��dk�������uF�RJ��          �xJz�4:F��rt'3s �i���@2=.��GL���Vl�  k=�^B��:J�"�O  ��G!�=i�v8 ��= r��5@� � z�G� ��e�:����b	J*��)�0R�)�@d��	�&i���UP5)( ��CS)P  ��
b����hh6S���g�������`���79���'�<��^3_�f��]=��3��a��f�3��x�`fg� ��3�0�;�����'��\���n�{���Nβ�Y':"4�n���Z�i�Ż2:�w��\��A"��{k���y�҈�\{��M)`�=^\f�4��pZrf�u��vq�n��w��X���@Gٽ	Tn!wͺI�0c6;xs�,�ڻ�35|�8��gK�m����W�/�<��Xp�����B�D��:8�ݫ�(Bvo.
[�Xf����]3G}�����آcz,���A@�G�LՁ-m��/ֽ�˥���Se;V��5�s�b=����d}�d���a!�O,��u�d��n���7�}.�;683w�� g?���2�.�{\����P5��F��:���,�1#�d��������A؉�F���i4N�,�H�}̔A�E?�mdMB�_�k
�z�"CYWp�mH4PJ�]3@��2ُ��UW��:���X�v5k�4'�.����)0���(%n�E1�%n�C�5K���8�e�����0n�� ޥl\'-,��?��9�J>���w������.U�Ct��PYf]�FQ�s��(�4K�]ˇg%�_w�};P�#��S�79q�3v�Ӥ������d��C^���,��ƃ�>0/5���k�{�M3q�z8����A]�nG�}�T	n�W^��ܥ��sK�����]Rv����D ��ƞBX֛�v���#ؐ�.*5�IJ����'x��C�g+�Lh��5|G�@;D�P�T6�EfҁZ���?t����7Ob9�h�Y%i�9]E�,��xw��R	&Z�aU�?9�I��<v�M�F��Ӡ1f�ˑ������XƸ�i��j�LcrOh7;IL�AbOg���1�m�$����5��%���޸�΍�㑢ŬvÉ�k���;nme�M��� �ɶaK���Uf�8i�sD�9��nA��7zgvq���סZ�hK�L $ek�Ɛ:]8<u�1�`
Cu��A�����K�M}��i���i쓈N0�pgl�CK�X�>8x�ʤ��y���}@$��h;rp���3��5���&lܥ��"��/(1�w&U*!�t�ܤ��u+V�ʔ�C@$.����͆b˷���ł��q��8gN������y�QU�LRΠ!�F�n�䀬��3��˽2<A晼_M0d�y(å�2�A>�jt�.����vn�m����Ղu �{�6K2�s{&l��o$�(��ZI^ˑ��	�:q/�l�}0��r��Ž�HT4��j�^Z.�V��_V��ɹ��=uV�̰����͸]`�$�I�E�R���t������d�7ͯ뫞r��%��,X&�I���ȅ�:�'z;f��*���w4P8Y]]{�8b9l͏!�����2E`T*�z��*c5�r��;�$�C,G��pP�A��W�#�۱m݂BnK�́��a����e�p!���U�����^c�1��+��i9��Vu8@�Ӻ�ٯ`$��#�AJeޗ"�!Y�Ӎ�*-˨��P0t;5U~I����5U���n��ؠ;-�nk+i�e�	g^�� h�HXYp��D�9N�׶u`y7���9g{D4�F:��V��x��d`��,�d΋��Q�snAt4�p��Wn�z΍Y�J�����8j���X�Xo�"d.8^�j@D'e����#��4��EY��خr�w8����$�G�Uni3�;]�y��Ki=�t��*���x�l-+�E9wa�%$)���v�{�L��U�'����j��6D���(&��Z;c�I��>_4���N�#���'ܶ�l����3�7�[��
W2��gzc��7Ʒɔ1;Eh��d2T�x�A�M��#��{V�=��@�:V���գ-i���ArI�!3� ���ol/M,���_boOn� J֓]7�����9#�%w]G�gJ��g�6*�S�c>�<��V�5�8/v�k��&��k���L�{P�-O�:m�ދ,���/�V�<��k3��#��$}3s�8kݳ9$cĺ��-ޢS�<~�Y¯��氄�tݰ��#/�#D2d5����N�gqR��H=����\�֍�~,8�!��ndd�󏊕=�S�v&z�=��qh%�Łڡ����YI��^�g5�5���,kήv���Lb|�[`�wr)ֶz�t�ۻ\�[�>{К2'x+GFWG��.���L��P�%6c���0��K��p�x��{����dWrmԣ����6�`����\ �׺���Bǀ����Y�G2�/T����*+z������m�8�e+"g���[˭��]�x��(�I��U��kjj�� S�!����ǅܜ�K6!x.��Bf�kA�8ɣ>��vP���#M9�'o��}�`c��>��*�
�6V�-
m�PĶ;�E ����]�
Q3��N�wM������]��uqLb-G��^n����GDw{���B;F#D�
�2l��K��K|%o%l�Ue֬�1B��x�*n�VSM�oj}�<i���f��@��Ef>b��҄�N�v3�#�X7�2�N��Ǖ^殹.m%I�7+ɘ��N�
pP�1�����{�����Θ[��n�xA쥌u�9iH77�#����e;n�޽�(�;�UN�hu�>8:��z�w{f\`L�ZgNb7�g�Ҋǻ�v��)��5��կf�"���C��SƓR,�aޒ2�sF�e��W�e����wQ���E-�i�7�u�4�p�}7/��j��XpW�v1�N&YdV������מ��F�M$�D���l�2�]��i��+�\�ud�:�ݲK�M++e�}��ye�` -�v�)���$�Ƴ�(
��w'%��8�L]���8~�_\׃5'�(ŤZeP�&�.��y�+&U3�m�#|N<�(�05�ˮ��^t.i͜�Q��4 �%�ؙO���b�D;��Ç�'�:-�[�:h!�vU��wZ�r���`V
mH�]�����a5T�K�qoQ���V��9q]vÀZ����F����L�&m4)��.۲�w&�F��w�˴E��1�4,�:��b�`�z���T��9p4�u��3��#�����m ���F����s�F1��j�.����YhV���ʫ�\�ql��]�7n�`��soQ�d����j�Wa��n�j�X��"[q	Ru�Ԓ�p�$Y�E��Ƽ2��N��>S���b�&ǹx�`��U�jiӼ�ٳaL�n�Ӧ�R��"}5�v>޼��6"�6
_1u�7 ��7��U��C�S9��Qjq.��kp�|
"Cg�w�:E0�0��B�R�r�	��7�]×H'e�sj]S��C�7����%��P.�ѣ7��7�n���[��nu���޼�n�"=7`f��
[�*���Љ��m(ów훩b���������8�$�V��۷4�AVɐ.ɰU��q�aqM��v�-��uuMon��2�W]���|�F�M��9���J��p^�^�t�m����l������F1�0�-����-X.�٥��P��Bak1�q�pd�����q,�S�A�����Y�/G��E�]вwT��2�v�r�5�;�Ʊ%�
B��wq��㩖S˷��iW{��s�W5�#�pz�������T�u���x�R@�q�M �Z�n���ⲝ�E�@�ٿ�@X�E+���eҋoXU�F�ճ,ݕq��#+f.��iu��ja=Ul�����Uo{9ǻ�����o�ނ���Zlb��&��Jד�CIs����ct�:̄V��*�2B���)F�űuI��X��e�zi��m��z��9�nFl�3����9�&a{o��w���ڦt�Y	Hz��+Y��7R=�U)'
��n­���Ԃ��j�c9���Qn��y��[�&�#Y�'lp7gԺ>�O��\��Ff�Z�8�ݢ]l�:��6�*�����T9*Ǌ�pod�Zl=~sN�4�غ�N�Ў��2i�����wy�s�&�<��>��ܪ��b"F��wH��J�n���*i�UO��IE���1˲���i9t�������	�>�N,ewv�=���� ,y����]�����VQ�����!)Q���#:�z%�,��^���۪�����:3���>��^�Y�F��x++	�\�I�hHE7T�F��-�6yU�fO[�+�.� ��㋙��㚴L�c��3��q�h�6^ү`�(f�EI|{��_:2cgP���Ps�^�j欱���2�Ӈ�l��ȕ�	��Ź��F��d����c�C.�}���E�T��x��l\u���� �{��wv�K��嫥�oH�]xI��u�K���4�$�S=.���r�lf��7�N=�L�9�j�l��ƠX����d-�"T2B��Z���3l�QB��b^�v�%]��7��	��Y�{
���6�~�=�����n*9���ly�wv8d۫h��	rC�Vv��p��o�j{�-���谱������y�V��5��-xΉ&ޅҖ�1Gvu����;�$5�wX҈Єu���*z͹ld� e��^��޴k��Mh�Y%�*	�_+����,#z�/o@��	
�MH�pS����ќU��LZ�-�JU-JYI*�v�P:�8s��G;Ƭ�����:-��@IZ�M8�觛��i�ظ��V���.���m���<H���:�3�K8��`�r�w��.����u�LC�b�r�� ���'>uۙAb����K�!��)�B�J|w��"/��PE�ͭ}V1���(������i����x���h��{y[�{�N°�\Jz"ov�e�kSQ
nR'NU��0�ea���V�n���{ bEή؍�0��E/��"��GvF#��FD0�l΋xH�~��+����_��궒�z(װ)Kkb=K�,�M����TRku叀P���y�N!4���ī�c�)1we��k��I	ZS;�7{v���߶�W�5�+�(V��mY�,9h$b�Gl<-��y$����iSW�JVv��Z*i۬�n4f�<�;�p=e��z����/Tv�.L��r>������DG��w6t���"@A�n�e�l�R��lQnUH�y�
Ȕ-�b�R��l$1�)Σ�s��,Q�D}��)mdB�E�v$�p���nU�e�:�fqKv�/���p&vѴ愲	L��J�V,�~�J��G6l�0�9f�Z�nր6Q��J?Q*���v�*�i圴�qLnT��l�Q]�
j����Z�C��ҭe��N�D+sb��K����d?[���G���J��׽�Hʤ!i/ R�Ǔ8r�޿+��6�R�q�9�{��� �u=�}�[a�↖&_��vn�d��Y�C�c����w'8��q��d�������{�j��4Gk;ԛ��,㢣Eu��A�^�����hk8���A>Ʃ�i��nA�(!,�x2Ы���ؙ���o�nE�ה�oG3����c	�X�'Y��*@�\��q�桻�1�R��9_�ړ{@���[��N<��:� o]����J�kW&.�Zp!���A�FS�iQ���()@�7*�j�w�Zǿ�"v��)�ҭ�a�oRKD�r�o�u�PY6�Jm���J��,�6�i��s&Aۊ�׿m�^I'pHe]FȲ��f'�V�9>��f��,���CY�d	�����;�M$۳S$���`�dt�KG*���s�N��	kզ�=47%P�j��bz��.��#�r�y����>";����~���:�.�Mvws=�%ٻ�w�cm[)�Fk;�*;m�q��v8�ʒ3�B��D��J=ڂ�E���6�B��A�B�%��vY9\���;���������Q5�"�F��C8a���c]�)V�N�O�wos�
d�Ӏ=qCYɳ� !4v�8�n��~_*q#��v�9 �bp��ww���M��Ckb��t�5RS-j}:Nk���+xr�w�M/�4�{�]�ô��c{��&�5���ݺiT}�S�N��٩�ގ,W;����Q�f��k� ��kG��ovjNV��,�.�9��".%�vd��NPra��OPv,��uf���J͒�TKtj�Kq¸��Tx\}�7K��
4���r�;Ҏa �B�C�Qp�d��Ĺ��L'%�^�ostΓ�c�Z㯙�W��ۋ�� ө��j+����ۢ��e=�ChF�ޙ�g�j=��H)ÉkCS����nhK�Lo\E�Q��0by��Ҫ��}��b�T���ˆ��&#�&n8jpk��C�t\x�rǽ����x��Ip�&�-���Zp��+x*xVx8qNa�>6p�K�B�7;�nO�]e�����D�h�ɥ`��_W�abZцG��h[`��7���ߣ�+�L.�)!��Ź7� ���d�;H�9`s�#�t�9�����O��t�r��)j�����?����sM����K���a����
�a���Na\��@����P0\������`D�0�s33"G0� 0��30\3 3�E����0\��P�30�C�0 S30\30\�\�3\�@�S3#�dL��0  G3s0\��0\1@p���p\\�� (a��0��G30�@��1p\����L�\0��fL������0���.fD0��fD��P����\��� ��s0��\0S ���C��1�0�29�fb� ����(f. (�� �s3 �a `��(`�)�`(`��`����အ�f�a��f�g��>������k�_�h)R���
���Ǖ�Vi�!ews�a޼7i.��Mh��މ4Ԃot�^߂�wڏ?z*�t6������<�Vwh�QWT���.	DI�;�:8�Hq���WzZH��Ϧf#f5��MFCN#7�p�#ۡ^�Ru!��-��(�'�����g'�;�y�NVK}��4[X�r�nc��_37B[�xp�Z�p����h�[\���8��Z,Lh\���j�gMx�ƷH���+Y�t��ʨi�W�D�U�S
Cw�S)��mQr�ׄ�#y��;wR��*�k��+��P��$��n9��mvd#��k%�$�!wwC3WgJ~��E�4�9M��F=�tSFH⇷o�r�f@�**_o���ۀ�c�g,��J�����T��Pv�Xg����%�I�wPNG��ZN�6��*H����F��4�Ю.�5�}j(�7å�.�Jƞ2h3�okP���u�砾'y�r��t^�D��\����a�E�ϫn�Qݣ��WU�����Je�ޝz�|K]rC3 ���Q����K3�֡��g+��*��c��j}�H�œ�N7'V�>�H8}"V=�{��BWh����t�s����[t��w�OOUa�\nX��ۑ��U];/m���.�8�|94N�5qnqwǴЏ�L�k�j>|�lڡ8QK7[�w��*�h��]�6f���y� v��Cg7<V�vw��pu������ύ��j��i���{�W�k���U�2�6��!Y�����5������W5:���4���=U��уo�=g���E.��M}��Mz����݇�cތ���DI��X=���ty�+���Y7&ұw��'>��v�[��1'��S�M�rG3E6�nA���d�9�n���x���j�ݥÝ���d��];�,y�}7/���G|s���b��R�bA�x^<���Y(��n�l%���z�쩏diu�}ov%�;r�G������<q/���w�'�l�+�z�٣P�x�V���~��g� V��o���AY��jmݛȑC�x�媽��Z�ם��wUw�=�H�O	��^]-�ʉ�\w�Wc:צ��dr]+p �a�)�Pv���ŷ9Ҿڝ9�T���/��0�u��ddX���'�vel+o��̍|�_�7���z74�l=}�tj�I��9�+'a�k�ȟ���@@��OmNiHӏ��ɀ�����^s̡Z�.�Y�륧���Y�U��&���wnY�u�oI7k��N���K�/��Y�J'�&��RY/ya�PH�c+��x�Wh��8�U�vu��ۏq�m����{���	cZ����S*�,nuH���S"]��4+F`�Z&�G� ��l�ݢ=����H����ƱE4ѫ�o$��3ط��4�	Ӫ�il;�F�b��釻��Up���G�]��^����G.���1�t(о�����.U����q*8�gjm&\����Xf���ƕn��,U�w�U�˜��v4����_jv�iz��Ó
`Ӭ,���q����[����*�Fm�lUS�Fc�Sz,b�IF���8�����2��X��vU!��z�f)���Ua�U]�m>�Q��!h_m�+U(2��D7���yu|C���}�N_l�12>�.�����wJ�=��ӱG��yqMQ��O������v�r&5��[k��լ��tw	����Ƽm�9��u;>Y���,���.��w�L^ـaiڋs�ƠkO��ȿw�C^?=u���Ӿ�H� �T����f/����^�����wep|P뮋j*E+�~��$�Nu�]T��nL�_��[/;5P��<c-�r/z+�Cw�E
cWf`5|*ꕰ[�����=�����$��Z�Pԟf�}����;yZ��$�^4�@��9;���.����p�����5��XwO\G�lo���d;���_��ڱ��6��Wixj����l!:?H�ҋ����z��ϲ
ͼ�ǧX*�}Z0�SJ��#,�]A�K����!ӗ�������oM=�\j	��V����W.収l��]���b��UM!e�4����9�o^�M�#�dǷ�pu1e>U�C�	��/��7|Q��Q�{�ؽ���T\�W�ٚ�qO�n`��[�m�wr�V�T=�ɍ&�9ɝwP\�)ʊY�}hW������wm�Y�
���:�{=�V:ܰ��ݯ.��ڀ��|(lg�]A#�ȼ^"wv6l��7�S�|�\-~�f��w��;�U��ES��� j�����pBi֘x���uI'pc&gϝ����ǈ�n�=�Ozf5vc��Lc�}�W�"¤�l̮!7�Ue+H#����{Fy{9b�Eq�}�ț�s�	<-!�zW�4e��X���]!kK|[���Uת]4����V����	d
�RX�i@����<�w�/���{��{{/(+�a��Xȭ��r���ەu��O_Q%�v�fL�{��Ju�����xb�t�������8�`V?TX�0��nVT�{����RIچ���,�������1xI��V���X��Y1�۪�����4w�K+��sU�X�y�_ؼ���s���!��XbM�3��D���0R(n��p,�R��0h.~J5oN3�����漰_k���iN��}���JM��U{q`N��O�2@���pFaa��0�MN�:j��^��)���\
?d�G=]�'G��'�2Evi�6l?5��F`����$L�CS-ٹ�h(�p��*��<�#��3��X�;o�OE����E��w�V+�n�D�oPZFf�R��;����_��CN�H�r;�ygb�OM2�E�v�ݯ�C�M�*|/� �˅��/=}O*	[7�k˷AѤ�p�9���ju-=��'H�xwz���]����ۂ�pB�
[P,��X�EK��*�ګ&܈t�q��������#�]�`�0��^ȸ���u�eCkCU�ecQ<�kl�]�*���р�fA�ҭ)a�c_YJ']��j��`��l"҉�q�\��D�il+�o6�s5c{�R��Lc��D�(�X�O:HP���->��[�t�g��g�8��Cn�~�X���1�Uh���aA"Dv�#�^0�b�"Az�s���o^��ҋz7Sr�5��eua��Uu��к�����ot��]΍b�RJK�_\}�ş=�{�Pa.�N�����{�Q8'��ʇj�Z�N[a.�o+;v��v�k��+�u22����g6j�tW�+;����bޒ�;]-}��g�'X0P#q$V��dW"�&�A�U���%���Y�l��8L�[*���n����!�*��ܲ�c=�5,�Q�v��<���~i�$�����յ�������0mglG���%���w�^D�^�/��^�m�S �f�.�9n�U�o9�Χ���_�������z�8�&�7���_{}��+��9)s��دq���؀E�V�nw��{����#�}�,�5x�w^���N�h�<��砬{����G�W����>��N7������j�UQY"�V��6��k��j�}
V���@s�!q�6���؎�W{�|�¯�Ӽ.�`���L3�VG{��|����]ae❃�Kk+w�:I�����P8	��g&k>Fy�{��v���;!xL�p  A����.�p5����E6��ھ��jM��S�k��ˈ��
�|{f*2�
�J�ԁf+�h���3y��w"d.���a����N��T���Ţ��f����,�/��ǷL�(�Y3u���B��B�;Z)��p1<R+;�
��貝w(�6���r]�==�t�{XN�lx}��J��zf���#��ލ����}繽T��bAUB8m�U��N�k�^h_wG��Y�+��7�.��U_s�/�wrBd�9��4uZz�/�i�̳+3�j�-�ة�8�Ţް���N��׍¾���������:A��{�����f�=q�nV�9x`L�Uݵ�>�I�u����׃��Q�Eo>���x��;�,�!�+^Z�_3z#C�9t����ǗǦ*�`��7n�O���y���w�=��Z��J��O)i��u�f�:��T���8͝�3wWb�O:�U�c�����F��.�4�zD���z+�,l�e��z|���Og�F��IK�`Ƚp����}��m��s^��.x����Q=�Bض�u;,�L�����ɵg�V����-#+/&�� ��Cu\9Wf�6�uG����Ic��9"�G�޴�����Q�ys��%Ӹfm�#�y1�w�`��/ih�ӽ|�˱U#��G�[q��^m���;(�����S�<^�{�w�Hhƫ}gr^��{�r#� ���m��J@��4A㣢o4|�ݵo�Q_���.�7X�]4e�ԗ<�m���� ����ؚ�����K,7�<֥4G�2��3�'����ח�{q0��̛ۗ�r��M�y�P�[���k�H��g����םHTǝ����E/y-�|�[�7�Y!J���(Uos;1h��y�@���އwx(o�B��]f\L��#'l�p��Nw:�\�wEaW���D�Ԗ㌑9�w���&h��å7!�y�Qi��i���E��v�u�bBt��|�h�:z��p6���6<~���z�����[�9�����x#U�k�/���̫��<۝r����7���[W��B"p�B��A�`��gDx.�����V��s������xe�l;��eE�-��ֵ��Bu��Ek]lk�;�r�Hyy�����g\pYP�ͬ��X�_*9� �vhP��p���j�2X���Ð(�K�^�s}0��Uk'=X#[��1V�`��f�L�yT��-�&�����3|I�{���`zx;3�R��*4f�p��fiAʶ}��,����}�,��N]�v�|O�
���r�ܝ�2A`ʶ���]Q�0{�\W���������E��,PF������W��ce�lVЉ����F�ޜ`��I���f���f�X\�ဿ6��*�NΦ��8��������`���C�U�k�N�w�lqZV�mЧ�k�>��r��B���`��m�� �:�i̕�Nw��Xl�<�,��gu���V��m��y9w��_�s*�Db�S�><"o��}�E�[[f�������7���Ƴ�h��ӗ�m)ng ȸ�S|�5�5�Ӓ�D�z�lObB�9���:��=Bͦ��<�f��ǣ��^�K�o���%�:y�o��]�`�Ǝ�NlY�3s&ͅ��Uk�������H2`�K#0�=���	�͝��}[����GkFL*DV�=�x�(لk�U��J�*9��Vy"MfU������������Чס�=�_W������aeR�O%���N�j,o]���؝�Gq�ְY��s9 k��%ow�5�24@;�g�z@�Ǜ��q�3|��E��Q�����/!�75{9��wx/)fK<�����p�r�I���H���A֖ j�bg�����z�'���s�L?��
<>m�4�n���jZ��X���I�V�"ǐ�1�}��t��b���/��-��`�-S�.NK���g��q^
��%�����Iq�z⽷�ڲDl�h4�|�,�h�����Z� 삑�/|�gwlhn����Q}���ϱΞ�*5:Ү���Э�l��FS�H���Q_wR�a��(xU�<́��٩᳀ɵ�ͻ�#/Qn�g��=~��>i�g�Yw�f��Jͷ{�.��샭j'�.U�:e��nd �w�oͷ�Mu+�犼F�:뺫J�6�Nk{-��S�irݜ��X��Z0�9W'H�KGs���M%j촕 ���ܷ{)���t�I*��;��)�菒���@�J;�uȽ��<9�RC��V32�e�h�wU�te�Z�i��Τ��ĵ��R��M��qv�( ��n[��`9�6�[�Sic\��jT^3r��:�E��w/:��6�G�Ϊ�`��کd��3p�a���K��:ү'հ*�yn�j�6��'��N�Q���E��=����40����� UM�N�裺�,mt:�XUk;9��GzN^Vt���y��=��Q��{T���x]��ޜ����֠���Εv9��|AUp��N�+oU��t���՚ց����͵��G@Ƅ��t�����>4��JT\�WV����X�:�R��;Yw�V���;�j�va2ƌ�`���z�TZ�5#x�BW���Y�y��x�r���l��)�E=._'����j�����lЮ�fT����Z�j.�O���7;#wE��Ԏ�g=�t�pn\.���׈�!3�o^'CkV�Bd��l�M���Y7ӷ�:�����hN�rOU�������;Ƣ5g��h�["��(0v��<%�
�Dϋ��t�z�H[��B�7��n�mN�j�X��"ۃ�=�]�Ңj�T�{U��iڕ� D0\;�=��c_Z��%��Si�o�B��xn�#ekٜk!�
Kz��P�TM���M��&��q*��!� Wңz&ԡ�kT�%�,�צ&M]��#Z�\!�B\VVt�>��\�rW�������߃��]��o>�{���A��=���K�N�]뜙V�u��!����,�P�H��
��.-�M�;I��>�,���&|����>^�q͡zb�x]�@�E��9��}�	"P�!Z����֫'���2{Í��0���O���ܛ�lov���<L�w��^W�Z���X�H|%�^S<O����37�feã`�օ��%�50T�]'wkr[pv�H�v�z�wa����`;=h��q":^e���c�q؝�J�]��#�n,ʓ��A��z�X�	��ݹ��m�q ;��m��<G���ˮֱn�����v�V�W�{<��e��n��4��=����1&�-mL��5�g9�؍ngF��X�gJ�[�B�m�l[�!ͣgn:��q�i�[G;�����i�j74.{:Þ�9��p�p�hK2��M�rN�svM��+��W�9��΅ɒ����]��X��"���ͺ�H�&�ض��͍v�5��"wc��{� ;��]�t�8,f<�t׳���9�,�8Cc��Ս��ݱs�����D^9��it��W�v����+�=�Q61���OW]�]���"�1W&sû"/�ؼ���)acwBn�U�n�v�x�yL#�q�78���x3����nMzzz��F����k�;Y�l/g�]�0t�97\7��z�Nۭ�5=���$ӱ��Ygmm��,j�ս���$n+��8��ׇ���5�E�����c��^�&��l6�Xܛ��Se�@M[�����vM�ڇ����s7&��M�nv���C���3�ܱt��r�1�8�;CKx��Yw�!���܌��T͇�8z��&V�gc'/9��P��]y���f���]�k���6��ۣOm�ݮ��W&���u�>:��z����ؘ�Y��ݹV��]�>p��i7��N��[]	w0h��y^x�n;�n�W��+�;nA��r��H�km�
kv���A�o���dƬppw`8 �.�:���P��kb�ɛ;c�s������X�Wu�<V��9��#ۺ�CK�.��5ڞj��p���y8�;���幪^��[��f�,��j뗶}���n��x���t>�ۆX8N��c�q ��E����]
��0���[�Y./ZW�9�C�,��v�W`�nݱ�����u&��K=X܎�L��=WUÎ���G���^����g m8���X�k"�=��e8��[�f-�m'�u�8��v���$��Tu�[ku�v�+�pv��7�[q�u�9I��Ϋ����۱.�'v{��mZ9z�gZ��3s{/K˨�]����g��ޞ��m��ո�ݘӓϵ5�OvW�"O\od*y�7/nK��(q��K˯e�;t�`�9�D��u�s��"k��e��PӔƣp�A��nQs�6���6-�9���h��<����v�V�cnrO3�,6�Ÿ�B�����p]��{Tvvۯ l��wm�	u��tnz�%S�r�"F���CK�x�W��^E��7<ե;����q����hi����y0��&5��)��Yx��x��p��6� j6]��vŲ��n�z���F1�L�X��\v79�\s��rZ8�1ع��\kr��rH���r���&��{a3���#ƭ�jj��������^�j;t{+��<�2v�щK[k��y�z�V�u�G]m�D�k��L�Å�p�	�\��vs6����P�[��ut���Gqi�M���pqY��=u���6����n9��R+��^ �+�% ]����t"�Z�.��Ş��z�8�wpyt�����n��%뫌l�9��mv�|��9{rHqn�n$l��Jy'��iDc�)������$#�֓l瞢�ȳ����r�����9���v��]m����!X�ݶ��(�7�pd����7e�;<st��q�S�;`�����waɽ�����s��x����)vO����y��,v/g�d�/s��`�(�ݚ����{H��i��;Am�^��WXu��Og���ι��y=l�2M%��os��MnC���FP]�z���ERgel���BQ��ۣ���ۑ���7h�O'e�Nl����80k�����ܽ�����.�&��`�Tev��u��S�������N����F�r�%9m���h��2���nn�]���6!ۭ쵌(uf� ��%�6�֊l����aӡ&�V�MU��eպjXk���ox�x8�l���9��k��l�8�]�u춸�r䵡<]�"�I��Pns4���6�:�����5��yƻ$-�݋��3�NT|���]ի��h��&ӓ&xLχ�.�V�G�nC�8�zvmN�d��̈nm5�+���y,��;.G��nbwj�3���Y��v��6���xGGA��c��x�ɺL��}�܎�*�YxúMWc���Xy�Y-���
\X�5�j�F���Bۛ��>�
BL[����z킖�u[e�@��=�n��u�2�Z�Ee�$Mv9���t=ŷ89�t�FH���'Oc����[�x����[�2�A��m�\Н��P�+ٮ�L�ۗ����mF6�Ұ��Zqex���I�5�n�͐�;@sv�.^=y��-�Q�Aħ;��H��Mŷq�x�y�k���ܺ��x5��Փcn1���G;��/gH�|�\��b�<���4�65�'\�S�Gcϱ�3@��Ƹ��kr�46�r�{)��hz�׍�� ;^��%ܹ����c�yU�G�ܩ=�ɞ���m��{n���wm���$�l�X;��s-��'������އst��z([=�v�B]�r5X|"ڹ$\nI�a�]u퍸ݥݻ:�E^�<vlr��;;v�Y��w�"�XM�����ٶu۵�;r�s���r�yW��p
�˹��7�68M���Q�ծN�}:ʝ�:�v�sn����Y��ǭZ�M��]���qs�f.d��q5v�v�]n��hj�ݔ��N;��G=�q.�ی��� �xP5�2��{)��wn
�6�:�nS�zh�m�N�o;v�ڝ�qg]u�g��O'��ڹŻp봜8Q���Ǝ��rml���W���$q�nj�k����Q���7
� cj,z�q��)ۛ���8�^Ϟ^��ٝ�s�]�F듙͑�{[A��ܸѹ�y9 ͮg�v�7����ݍlpݯ"n���ۓi��u�Gb��&^�k���猵�=�^�\�,���tKa�9�.�v��u�^�&�^�ݺ�|�ŭp�V�YA�^:XS	��n�܌]΁8C��q��b�8�a���g��6�t"o)uϞ�5�zx���W3��g�b�[�Ă�6W�q�c==����g�ɮ���郲j6*��� �M�>�ٍ�=+r�N�^����v{.W����OUu��6���w<]g<n�	X��7j���j3�Jh+{p�^ܻ�����#Gi�
ll� �7`�k�]v��6�n����Gn9˂��N�sI�{��V;thSq�r=��g���/5vZ��	v�V9�x;���d���i�v8�'�#�vc��Н���m��v��ˑ�;��Ѫ|��c���:㶆��w5''��I����W<u�ۗ���zI�S'
rc pTt�K���l�g[����ފ�=V@���B�g��jz�e(�yX|p�����yC۝ָ��M�殶�c�,�ܮNjݼ�G7�%�r�ǔg��-���zѻjt4�4t�m������JA���B��d��]J�[��·nܪ;�&�Gn��	�68�8�5�ێ�0^nl�g����,���v�!rB��j�'c[�Iѝn�"�t��X�����CCq+�jT�ݳc�$p<�8�އ��m��V��O�]���k{&�ƌ�`ՠ�e�\7)��m��k.�E :裭Ak�x�;�wU���}�z�E�ڑ1lx�i��u�T8�tk=�2�n��}p㶹�3��磃v�ޭ[��ᶻvPf�.��ɔ�x�����iΨ^csO��D�ꍐ�62�gv(�q۳���=�ݳ������e�ytz�vV녺.;]'G�v���خu���l�^؇sۖ.�]���c���*w�q���U�q�s��6#�,�n5Z��<���nڮ:#tu���jxXf� �TO�9���	�FE�i�E�0WX��F���[KD�OG��)$]�C;]�۰��ך��y�s�ض�-mv��s���]s��j���i�l�X����VI�{Z���۞��\��vM��`���R]sjp���3��q�\=��D�x�q�H���ˁ�m�r Ru緱ո�޺w<<z�,q���d�k���Ƴm��6�0m�g6��ֶ����M�k��XG��5�֋�P-�n�9�n�q�	�������Ƹ6�l)ۮ��l����8�Ә�H�n�D+��;��Mc<:7=�����kv��^&�ٺ�b�os��x���[��˛��g�{x]��6��Ǯ�p��b]��ܲ��n��X.P-@�"�s�y��G)g-��8Nuݮ�k����V��C�+�v�v���qt����0�s܇b틔SCgY����;=�������l7/=z<�vȗ����]z02`��3$��s���p�䰷)�:[�:�416���f�;vڞc��K�=�b�Tݛ����k�����m����;���n-���k4��x����uv۵���Gt;v0J�%���ٛn7S)�^*�\Vɂڣ��� �����ю�bzS�q�C���帀���]�Q#o$lzH�����V��]����k`��fٹ�Wu���Fv\�Y���[l=g�+#��rKsq��0���iu{h��5ӄ���6\˝ؠ��v����#<�JM΅�.�뵽����C��wj!��l�չ�=%��+%��8���]3�ܞx����Q�sA�ٺ�j��s 㭧Ɵd���Tw�Z���֣pM�Ȯ�K���m�s�yMv�Y�v;<�l�c�v�,�l�p�lHM2�0E�Zk:{[6�cV�箟U�-�ƭ����<g�<�cn��cE`9�`�-�m`Ă�eq$%�i$��
��i2-��$�V�8��(��I��V,�(0AF@�A"+!"��V
L�AfD�)F$$�#�֫B1H�EdX�Y"�"2�G$X���+d���HFV��\����$$(D#�cX����R$\��	�A���qY1$Dqc$���"đr(��E�+�!V��X*�U�I��d���q����ċBF��c�R2F1��U�&�XDd�222AcrEI�## �D��c!dGd$RFH�VFI0�9�(���-A"8��Qb$bLE��$fH$b��"E��,�QQDTUVL�#�����dr,b���Q�eVI���BI!aF0d&#$�����(�9fL�$d�bL��Y�,I!$�Q�X��H̀��QI&""�@�d`��$HFb.2Dq�E�dŭ�&$HL��$V1�$p���+$\TH26�Z�����s53�MM���K��j޳�iL�ݫHZ���uM�-��n�d9���v��۱�x4�G�Z�V�tWH�m����9wn���m�ɠC��-�W+�ق狷)�n�^C�qj��0�u9m��5�@n뷎�ټ�w@����pzn�su��9�%�ϲ���[��'�kҷ0�����k"t�>��=��C�k+���X6܆�m���B͹<d���8�=r�μ������6ڮ�W��<N3ь5ly�0G��u�[usk��lv�d՜�{<JK�F�f��m���"������
�����kӞS�eGOj2�m�����w>7�;kq�؞�:�Un�[=�O��m�l\�N���t�Wl;� �v	�<�nB��cfK���eQ�b�4.�=���m�hN����zݫK����n.۠6�I�c��;�4l�n�t�y�[uu���<��ZɭBL�k,-���7�Ɩ��>�su��7v޴�`$�mL�!���]v�\9�n0׍� #=;��t=��y^�Ib��\�X����W�M�[t��:��d�㝽y��C����i��������%���]��E`���;GY�緦�+u�r4)[0����oJ
����yۓ��r�zl���;��l\5T�+�z�갏J��N6�]���t)���cv
9���sq�m�-��=Scۓ��٨��6rH�r'6����LNp��v��b�4oo}k�|�n~��Nw������!����NҜY�S��c�:�덍l�@뉶��v��g�v{I�Ϥ� ��Ϙ�����ۦS�Nj���7���,����Mx|6��!�=���9\v{1ƹ{r�Q�s�b1�ɱ[�>u&l{v:�n1�5cG�Q�Hs�z���]�#��v��98�;��bօ�l[�Wm��A��P�]�0"vi�p\�������":�Թ=u�q�[]g�Q6�.����N�� �Q�<O�������X1T���ձhZ�r1�,�\KZ�I����(��$ �Z�Z�E+�F9I	+&R�b4Q����QkX�h��X[LZE�k\�*�d�%���V4�dY*9�6�Y2�k	cF�l�e�u��XK1��XRʕe��@�R�RR�-�ib�XH��D��JZ�lZZ�����b�V��Z��Ȓ��J�"��پ��AL�����˹!�c��I7��haw�V}~;޽��I3}��/E�e��E%>���$m7Ԟ�-7��� �f{X����8�
�4	�s���]E�I�A#N��z8	�{�O��)1i�t��v�H3�����'�)���Q�Ӥ*��g�>��:�M��I� �e�2�>w��緭q}�f>����$��j/���ʘA�J�����I��t��n�'s�p���bo�d�A"�=����=G�����v��� �ח�ݢ&{n� �:�f&�x��t�JX]UI�=<��u�V��=��	{�d�O���zX'���A��A���$w<�
?]��B�d4����]�S��V�M�Gwc'Y�՛�_���8m��48.��3��O��Ou����~@S`�L��:+ܚ[}wl�ھj��G���?|I ��a��O׹ޱe�K_R�ywp��~'�1�t]|�TZTR��.�� �f���~1��^K�xy��4{w��@��z�˩��)2�T僸��bݐ��l�W�8$�=����fg�q:�>3/���|N�^�XD�I�LU�g�Y$'f�x<-��=�w�����H��u���Uz�V�D�>1�ܡ�8^�띡�k;���C��=�Џv���q��8�%։m5K������$i����&c��A����$�����:u���}/����u��W��L:m$�d�u�$�����7�ݼ�[������H��� &���[�{����o���!S_4傶�� ���s�I3W�ݍ�'��y^)2Ba%�W�r��p�ŗ� �Wl� �<�'��,il^s��Ғ���ᚊU��>�I��d�'�����_�iX�H$gg�b�33�R�E�ͅE�����ױ,W�Ʈ'��*�پm$���	��c��/x�ɬ���X'f�|���)��������~}�+����s�.Œf瘄��c��+d�j���k�SJ
�l�Ai�T	�T��ͺ��Z�4 ��s�b�����ʹ�?��]lr��5G�}�v~$'�\$�N�� ���w���w՛���?fg9�87�+@U!)`��9�%�c}��o���޲H$��\ ����?]{�-JB+����Z
a�i$%���H=�� $$�������s;����X$�� �I�{X�ߨ�MPH�vW]�nJ���c�ֻ�@H$_�`�����_yз;n��c���;��ܸ����/f_��}%!�%d'j�K��U�}tׂ{��b����_7�Am�P��T� �g8	��<.���
�J�C��zA=��F��wfm��|	;��>$ۚ� ��n{�`����3I���/�F���[�K��v�p0&����@0�n�us���a뗣���|��͵_=������I �3s�w�=

�����?�=�����2i��5UFϽ�g�OA<X���瀐	=�� $����$����;�Cv��n|HѾX��R�٩~p�I����|��.מ;���b���83s�v>8�
a�i$%} =;�<����P�(��)�| 3s}w� �v���ʼc*�3	��m�u���A�e�r��X�	����wOz��'���	y��@$��4�)ú��k���<�����t��ɱ��\��mfAXZ���m�c���أ��'�W9w�ڥ�ز�-1�7>^�B�Tj��YM�7{��nzw��("�{;Jr�i�i�t�0;�-Z���rx�O���n���s�׎�]��W��lW�v�c�}x�G����n؞�f��;Q�a�n����3m��ma��<�gn]h����Ձ�1;c���A�g��mp�����-�§��Y�v�W]��'F�c=Dն0��^�v��V%�����i�m�Pq���]`���3�XpImu��n������*�����s3\$f{���r��A�f���-嘽� A�3y����䯁)���
n�긅�t4Ǖ���H#ݛ�d�F^y�A�<��ܚi��^���@⢡�&���۳�$N�pO�'�}*���=�WC_��3��|� `R~+�2Q��O�	��-���W��d��IN���$gg8A;�ƽ�I��v<�O,�]�	���S�I �+��~�b;ۍ`���C�-�w55.	T��t���Û�>����-�UTȪi����Z(�#����9��n4�Փ�l]���X�������Bi��D>�d"fs�	��A�t�O]�5�� �e�0�/���¢Ң���p���[)���@_���qg���R�����̦.�]�"�];�T�ڻ��$�,�G���ޤ��i�4�}��U��7�3��rw�/��$��w�ρ��;7Ư���5����oQ����n�S�:��BA���	 �{�;�f�{�������e��$���;�Ѱ��4��4 <��'�o��c@"�5�@ �~�@n{�1��F�C�'��p~3B�K�5H4BWf�x�$��۳������	x� ��0`��ٸ��-��I����C��MR��j�SF\x�^rF�QC ѺƖ�m��)�f�6�y燞�i�J�%}���p	���$��n{��s�~}�3���8	'�{��?b��E"L�Eخ��J逊6�oQ�<&_�I����A�7=�fb�k~��_��vg5������5TR3��~��ٞ�`��C����Ntߞ�.�ռ��i䫟��}�\��Dx���یoZ���U`y�~z���^G��N��	G1zi5�G�n��F1Y����e�` W���ߓ�d{x�j�d�J��Vy���3W��k�z���A��s�I�s�vH${�Y,Xa��%S!$���p�zC�QP�U)DX>}��"_������^�=$)����Ad�{�
���^v�T�"Ȩ�;����r=��������Cl���=��1��z2_�Mw��K�h1��[�����<����Y����〿/仇:�>���'��{������L6�I&�@^�{6�B��ŖހH��oK�/|�'�߰�p����۟n��T��݂�w�d�/<���M[�^M��A�o]�H��p�m��4�L�MU�=y�G`f/jݿej��A�7��&_s��N����y1O^B�2��V���E/<�qn�x}6H^~7���#��xs�ʑRj�w'�:g�(Z�uUOLo;�mjj���5�+�SY�(���fX��u�j�`��S�:�� �>7��!��=p�z�ݒ	2��|I��*˹�5J$�
)6
?&�i�Z;]-ţ�v��6擘��]:�-�-=���cI��ߜk��*��-�hx}�b��}�O���� >��8�]��D��O H'�/�����U�D%4׳!m��SW�o2���A���$���s��Y���`9+݈:��/�<�<�l:T�%���'��{g����:>�;��� ���� ����Q	��/���n��H�
#{#��A=��'Ĝ�����v��+t��'�<Ğo(ӤBe�j�$=3�@$��z�ߎ�f�n�s~#�	 ���$�����љ7�����^/�V�}:M������
�V�2�:����Mo��Og\���cX饜[z����|�Wݺt�>{����߫�>���;��ֺ܃��an �^���'K�m�l�T@��4Rq��Q�Y���g!��3]N�#�u�Gmvz���9[sɻ\V�k��siQ�q�"�s�r����rۡNݙ:����8Wmul*�R�"�w�`����G#��q���vm�n��v�Gs�+`8��s<�&���O9�nx�M�c���#\j�v��M���}W�=���ջ ��Q��W �O<%w��0�lc�;k<�8'Ԕ6�Kn����ϛ�9�[%����:�\��~��'�A����p�'�^:�B�k��6k����a�h�h@y��Y�d�Ok쁦��A��������;����:��v��G��+�ƪ�4Ph���{1�	7پ�H9�@����t��|�'�������ͥ�/�M�a'D��ﱍnG�c%;��I�;��I��c����{p3.�<�z�IPM��|����߬Y�/<Ǽ��t',������s�O��ޱdK�9��=p�N�����O6Qd}Ll�k�N;f�0\���/k��M��J�;P~wo�%M*���g�cܫ���w���'�A��bϭ^�9�,�?@$v�z��,�E��-�i�ڿ=�OU�	����-��Kb�+�s��ʪ]�����&vb����븻���aчs�k��)!�]��t��.�I�T軼�7S�Q�zl;�:zݿA's;�Y?{�	���~�*�;n�li�c�Z1h�A��>�ز �~� ���sl���`߁ �g�_ĂA��s�q�p�j��EJ��cNϋ���oĜs���I2��A 利/e{Y���ޗv-0�§D��}��$����ꛭ)���j� >~��$�g�\$7��P����k�k@��M��l[�ѐsW.2+��b���u�%.�x:�u�K�t���D$�&�b�O|˾�d��3�	${��C�gmN�tg>���޻��f瘂[~�N�I�)*����15�����W\d$������z��plt�%�*���̉R�UB�%U&�9�Ȑ ;7��$�>iF��Q���~`�/v�)�nc����x8G���xg��ۮ_y�i�M{J9fyg*c�銔���{	�.ɼ������y<�U��ɘ^zg�7�鴒�h�I�X�Y�{���v2�\��}��B���.��%u�G�Sn�Mp�f�]�c�/�����b�{�J6*J�G9,������Jrlsl����*#[ Q+ѳ�5}&�9qn�g���ޙ�wW͞`�'��F�fc�@X�K/��_,4��[�6�o���[N��Wq/.r�33r�?��Q˧��g
b!��R��^�G6�k����ʥU��m����ED�R����'�,���s:S<��-U����vn�ݒ��A���p��ܮ�gh�8**1��ݲ�-Ժf"/nZ�B��/�j;q'䷰��N��:3E�́J���i�Z�;H��Ѳ3M��}{���u_TZ7�)���{+%���Ŝ���kǃ8�I�{����C�����.�r��L��{��t�RM���SЯsy���+7б�.>����.��.�����0�u��Zy�Yi�SRf���/k���#�ԏyXׯӕ�>+�f`z��״��J�}ʞ Mi�v�D�����U;�-xuߵb�,�C�Ә�*�=7x��լ�|�#%ݷ[�1�m�ґ�����$,U�w����ej���<|�eXϺS�ޭ�]�%}鼽7�v���L�����tx`u�ˬ	\���\�����L�]��sA�7���X�ĸ��!�Z�Jſ/���~y6�ñI���!2HHȋ�D����&*���D��H(1��b�rH"I$���X�ઉ�.Da��!`(D�F*,����&H�����"�2H(��d\��"�Ed$!��"��b�d�$#���I2b�`�IPqd�HF$�(�H�DD���LQ�@��d �����k#$�#��Fb� ��+(�F1 9����X�"䒶�U��$I�QlH)1�Ebc"�HBD�`�r!
�E��"I&Bb�2d�F
�A�1T`Ԯ"W"�+$�$��h�
Ȍ#R.Fe��ř�$��G�� �bI��#H$R	��`���D��2Lca�0�bB0��	�REb� �I$qFGY"3$R
,��Œ,a�G�I�H�W�H9�TJ�F�9T#�$H�(,�"ਂ ����.2
�1���$$!$,RĈD��d�EE*E�R���b)EE� �)$��Y���j�ݫK���� ��n 7'ceTTTL��E�;ޥ����Na]� �� G��m$��4�.[�Ԧz��@���\���52|�1Q*e7�m?Sa� ��U�\����\k���
ʺI{�դ����7J>]Px��4FE'�e�T�a�/vmAb63\=�T�ckc�}2u���ۏ��ϛ|.[IBU\��
� �;7�ؑ ��i(����)N{8=r�J�vw��.�Q$�71P�����w��0��{U1�y�3kK��7NB ���������4�J��!u�j�Y�9Wn�`Q���d�]8�mZI����Ӏ>�#ܣrn&��0  �w���D�wU�.k2%HT)�URl3��\�}����뼦��7��������A��૿��f�趬��b�OF	�����wj6Ȯ�N��nkM>���^�$j���^�	�X�Iv}˕Zy)�=�:NS��;���~I��r�V����7�:�J�R�y�O+�Z[D�4�
gS�W����ǩ��L�Dȓ��͛��j{���K��צjI�>�9��1$��|�Xq�`�G �D"��A�!Q�V��F������Y��.d*T���gl�d&�i���2�;�ǵɼxx	�GO2�����jٌi������]~���:=B�R�����~��q�L��*eB&D�����i�8%L�w�v?L�u��.d}y�I���� R�*��}^�T+Ow���V�j�n�h�B'D*^{��6�CHW)����;�~���4���A��@DJ�B�B�_߽�}C�jP�������m3��27������v+�򂷾�_�I����w�D����\:��#�����L�x�ʅ�ʓ������-�eB�~����ݭ/��w�-��,���d
#�
�B�\�{�ϵ�:�\�TȄB�K���f��i
�C��ܒj
)�)*��0�>�ސ����jk\�!S"3��s~w\z�S+G*eK�S*[�7��T�%L�Q����߷�8��/ߟ5�/�xg�DȄ�����z�P��k��+d��%k�s�S�/���ͧ��9P�\r�_�{�{:�P�k~��>���������T+��~�P�Z�p��*e,/kݛL�D��r�V���~�>F";���3{-p��Q�j���Y�u�ٴ��OQ��.rbΔ.�N�{ݻ��s��X�$�n�e�x�_�א����
�WL{��%{�+u^M��9��? M4�H*!��-=U�ڌ���sqjCLL�FH���7���Ml���r�@��T��;񱖷b��<������7l����skq�ۄ5�7nscG�m��z���f��[kq�qk{qcX��:�u�E��of� u��'T�9:��r��C�N�}:��k̆N��N�ݮ$Lbz��mm['K�Z7<�v�z��lp:�n�N��L뎌.蚷.���W�i��}����%Ѧ|)�O��~����^�W+S*,2����f���*2!y�߹�:�N�
����v����Ǳ9�?!�	￾�����B�G*2$��f��i
�s�>;5l�4�[y�q�W_w�������s��~�_&���CN�����ΦV�s*2$��f�*q*er�2�>���C�P�P����7���|w���aorH@ӧ����~�m�I��&b��2$��ͧ�!S"��B��߷�8�C�P�T�W	�O��y~��߹���?8~jB�[ߵ�ͦsP*dB&F�W�{���S�S*S}��,����e��i;�\/����糛�ߵd>�/u�I�����a�'>��L�Nd2�Z�P�<�s�u�**
�K��~��������]�3�VG����@�>�����pHW���rI�F���^u�u�W��}��^�S-�S-�\'��}���eo�>�|��߾gS=N	S*Oߵ�ͦT"ds�L�\k�{���P�a�	HeBم���ohu2!�{���ϴo̧2�ī�j�kN�F6�+�	��f�����,�L6���>�\���?���Wk���S�B����ٴʄs��
�*��}�ι�*�P�P��~��m�u�W	�ߟ���o���!;�W�vm3HD���*eh9_|��N�Tʔ���x]��ti�Χq+�߿y���ȄL�r��~�o�y�N��Ny�Ya�zY��[�\�}�}�e�g+�.o"��1K��oRw7Г�9�a�v�xcO<�@������&��f��P�Q�nǴ_��V�
�����B&D"w�W.%���ohuΎT+�ʅC�\��M�I���6��#����~;m��Em�C��u�oxq�а*e��Oy���ΦT"dJ�2��|u��Nwϵ�zm3I��2�A��ˍ|����C��T%!�ra|����L�G�}�w�m�֙tCF��2$���5�&�l�p@��Ȁ���W���{:9�*�S"�߿{�6�\:5
�A�T�X^��l�g���߿{�L��T��+��oxu:%L�C]�[R��\:���W�������er�2�K�;}�|fп��������_k�w񟐯
�w�8�N�P�P�W*_߾�{C�uʅr�P�PJ����6��#������o�o��ɵ�W
�R &�4L��n��m��FѸ�<�Շ�;����������P���-��x��>ơ_?y��ǨT˖L��\'��}��s����2�J�R���p�fӉS+�^{��e��߿}v��:y�oxu��T"dB8O߼�{C�\*��<�Z1���q
�y��L��9P�>��y{��י��~���u
��T�W
_?y�6�\:B�V�S"I�>ٴ��S#\���>�����[�3�������)��hL3P)�OR�]���۝z�P����T��y�i�B&D"dB,޼�����},�'�Ҋ^�'R
�gO^�BQ�����'��ڒ���F՝��h4Nd����tec9:�;a���a��B�R�T+���Ϸ�:�\�W(�B�D��}�hpN!\/�zv�*1���ȇ\:�+��~��kI�|�篵&w,
�l
�<ߟoo\�eh�L�R�T�o}��6�L�pjeB>}߷�8���������^P��ʅp�����{�
�����j�u���Js�"I�{�i�!S"2!|����:�C�kS|�����~CH~J�p���y͡��
�������f�8rL��*en9_>���B&D}��~����5�,��3Z#�m��V�[�=�#�����YK�`5d �����/��̺��3I�W������z�\��ʅ,2�������-eB�p�V�}���:�N�
�������W���<s�_���huιP�W*
�,��l�fЎ9��9H�WD��mãP������CI���d��Υ�>�~�=!����2�J�R���xm3i�*eB&G(�ϻ���P	HeB�����E�H�{����@���_[��EUP�ht�5�*N�,���6����B�D#��kݝs�i2!�T~����F=�~[�<����?!\+P��,,���g@���T����ϵ���2'}מ���ZVH�.�#�#�����O���}�3Nz�ʅ�ʒw���g���p�W��^o!S�T*Q
�~���,�W�:X~��_��KW���P�g�'}�h��Ź�X�y�Lz ���U|��O���/&�4u�z)�/_5i��&��\��޸��� mϱʅB�K<�vm3hG�~��TcM���tj�}��G�i2!)`W	��>�ރ�L����{�ó�>���<NbTʖ���6����2�A���5������:jP�PG�Y߿H@��� #_�y~��9�x�{�_W�]q���n9���.<u�;b�Mu�MFc	�Z�]Lg؂پ�??��!�7<��w��L�'{ݛO�!\��
�r�_;����:�B�P�Q*������L�G�����^����~C���<�6��@���T��+�|�{èDȝ9��Ȳ��4H���T����������pjeC�y�ޟ��g䓻�f�6��!�
������9�P���B�\�{�ohu��
��o��:/ݗ�_���pB�,���I�x��.��l%�PۇZ�~��w���
���,
�;�ﷷ�u2�r�T"dG���o*��~����L�{��2�F�W+_�������DȄ��}�{C������J�!��i�j���}DU_~�ފ������4��r�\��
����g\�2!�T+�/����C�jµ
�l,����!�sڻJ�%�B>��?">E������0�Gȍ^��L6UT[!�S8�J�~��ontz�\�L�\��U��	t>�~��⽤Ǹ���e�D6��
���~�0�:!P�q
�r�}����s��
��T����@�,�����uL1Ig�w���Q��S@
rO�����o�����?{�6��!=.f��������i�Ǉ���	���J��&�A�?��<{Xo�8�?���ng�;����8��C�IA؜��v�8��ۙ4�^�b��������̰��<j��cj��v�\��+7F��nn�;��u�y�\m\nq7=�$+bz�q�ݷgn��x�аfݸ�Z�'�=�<s�D�Iظ1j5��)ٱq�ٟmv�����6Ů(��Ü���������g�-9%nȕ�/<u��#G49�\���\S���>�+����*\cՆ��y895�ƴ�Zɢ���5����ֶ�B�ko����j�~���3�L�p��{���:�Z9S*T��-���L�29gu���i�;���^{���C��T%�eBم��ﷴ:�p�V��;9&��ZkE)�:�N�,���NbB�G*��	���}|��P���<��qΡP��
��\-���shuø�+�j2�{϶m3� Tȣ�#�o��K9n{_����=��|<@�>���s�VR���:��ʝ�}���νL�\�P�RO��f��2!8T+��ݓ�Ϯy�g��p�2!"Ή}����s�T+��T*T��}�hq8�p����é��%B���@G��Hw:��U9>��P��L�`W	�?w{zc�L�DȔĩ�-���L�pJ�\�S+����oxu�����<�>�_���?!7�[0����z�P����ZFkC�Y�aP�dI9�6�q
�r�\�T+��{���s޿��������
%B�[�>�C�j��P��$���g9�F�Tʅ�ߤ�YB#�C����?��:��pot<�c���h�s[��R�O��3^�b�Sϳ���}�����Z6.���S?!'���{C��Ϛ�P��$��l�g��������!�T*w���^�듞{���z���;���:9P���J�y϶m3hG�����+Y����uíB��߷���
�l
G҇�R���~�j��^L4�-����L�ODZ��9���&����D��1�������P���������Z��u]6���}��!�V{�!����*eK�S*I��vm3iĩ������߿��:�r�*2!;��{妚�+>�~�4�?@E}�yWT�z[�)�:�N�,���N!�+�ʅr�P������9�*�P�P�GK���?x�o��{�8���P�����<ٴ�g T��ʙ[�W�����S�Tʗ��FR���N���|�ψG���C�o����������{��\��ʅ,2���͛�C8��2�[�
����9�P��B�R�P�\K�}�{C�:�{���o~����s�9P�T�g��͡���{�é��M+n���;�B����tz�L�D�X�w�>�����%_���R��{�#� QQ~�6���%L�\jer�������P�T%�T+������Ǹ�P����Ϟ�����¶���`���BQ�7=�ǞwO�hʽZUqt�ӳx������d�7h�aP�dI9��ͧ�q
�r�\�T+��{���:�B�T**������p�P������g�������兝��6��"dy�T��+�{����Tʔ�^z~&�i]Uu��3��+������ש��L�k�|<���?K���!�B�D#\*��>���2!�T+�/}�����ʅ~@����E��?\��mg�AY�S���I��Yh����w�u�oaרTȄL�p������ΦV�Tʕ*eG�߻������u�A^�D����������]����6�OV[�(\�B�ɭM���	�]iKR�4�u���"�bz7��U�!���|�;o��3��|�6���J�\����k������;a���&�{���׮
�����e��u�E9�P�a�������߬�������@����|�ι�**
�
�K߾��C�jP�������i�s��>����u2>�S+G+�|���S�Tʔ����)�MC\:�S�%p����ntz�\�S*�ʒ~��6��!��6��pȄ8T+w߻�a�"tB�R�P�\�Ͼ���r�\��
�ĩg��f��q
�?~�;�~�ý���
]Vj�X�7�"��P�tjL�8[��5�Х{�?߿>:i�un��߽CnB����u�2�2��w��oo\�ek�2�J�R��~�͡#�O�{�k]9�͹�^�߷�:�r�*�2�nL/~����*����bK�ԗW�T:�B����Nq
��{���5y�:y�~C�����!"R�\-�����Z�p�P��$��l�g@QG�G��{�Y���+�h���}'��"dOu�I�ZGU]T�3�G	����������P�a�$��l�0�qp�T+\*���;a��ל���j��;�0��L�DȄs�{��ohuΎT*dB!D�g��f��q
�~�N���kE���uø5
��{	�>:M�&xL�p�}����:�Z9S*Q*eKo���6����52�F�w﷼:��o��{te�6Fx	�CS9���	��\��Y8ݱ����K�s�`K�u���=�T�lּnE��o�˞�}!b��O/oyɗ��[�[����s�0��;�Bʅ���y����^�
߽���4�uk5�iy�P��*Y���ͧ1!\��B�\�W��{��s�T&�\޼����>�==B!�J�p�����L�DȄL�XY�|ٴ͡#�*ek��?~��
#�!����WЯ!�� �[��v�S�i�A�F�fY�ټ���N]���V��][�N�#)_)�j�_&T��^����ΏS+��P��$�߶o��!i�V�B�<�s�u��T�<�y�z4����	w�����:�B�G*
%K=��6��#�����4³WQko:��:�+�}��C�G�P���^;����p~��$8�S+\��*Tʗ-��p�fӂT���W+_;���C�P�!���~�?�/w�
�d������=��bK�ԗW�T:�Ny�ͦm烕
��W������P�PJ���@G�u�F���o���?��@���j���*e,,��vm3hD��r�V�W�����S�S*{|��M-T�p>�3��/_��*e�W�׷�&W:�ʄL�'~پ�!i�V�
�;���B&D"u
�?"w��0���o���u��x����B�D�^y�hq8�p������&�XYȇ\:�+���{�B�R����N�����ΦW����}7y�����g�"dOK|�8m3i�J�\�L�\k�~�{èDȄ��ZL/|��G�@�@�P�m�Gi�b�Ľ��s��^������x��Ȯ:�H>O=o�)-�M�P���VM5w����c8�<�:^��Jb��7W1���бǫ�+[:�Ũ�V
D�Tg4:u�;��
��Ր�Ѕ��,�9r5�{Ww�$�ѫ���xc&��v����A��W��J˺lf� A'�E�tj-�'��t�nQbG�D�粰muH�Ӗn!�%k�uR,����ս�^�oW�!�$�q�VA�q�ْh|�,u�kzFV�p46�Ř|��7R�s������:=���BP>i+N�Y�m��%fiMkg���Ł�+8g�dy]*�Vu���;�v�(�59�u(oXxsvQ�k�U#}�����x�j��Vx��x��ص��<�]\x�[-^�0=�$�c�C��݆�piɾ�
�e��,��lG�Y�>J�ג�ޏ��WN{�8�ge�tr�Q�f25+j���*��������W}3;{���Z�P�U��n{�KOe�
e�WS�+��t���;�P=5�p�Mr��l�Ag;�k�s��,E5v�Gu�Np��	�FV�Q���F��T�!V\-�!*CQ�H�^�z�`2������Zsc����`w8������q�2��V5�`����YS�7�x�\���ܻ͒�y麮�u�p�A�]���uS�����j�Ï"�+��2��a�7n���*h��:�{`�W�&���`���)U��5�2&�ޫ�y*T��{��،wvG(�1;�5��c�+�������J�Q�G� �9��$�E	�"�#$�1�r6B��������&"GEȌ�$I$���H�8"�ȊCEL#Q��"�#dG�"Ed�bW#a�$#2pd�DdV2
�I��F1��IqR	����)��"�c$����
�*�&"2!�!*6ڑ#qFI	����D"�EE���aBa2L��AV3"�!l*�,�2Ec��d��U\UW$�B؃��Tq$�1��$V!1ŌA�1�V����I��Y� A��QaX+�Dc����229�&XU�b�E�FHI&1�$I�����$rD���FI�! �*1�"D�a���F�a1G �(�$�&"&*�"�$� ��1EH�HH"�$c0qda�++EK�ĉ!$�������#��d�I���8�F,X���$��0E$��!I2*�1��㍘HBV
��d�#*EK	2AX�Ud��Dd\U�da1��"�"F#�Ib@�����&GI1r9$"�`�	����$GG&H��E��!A�R0�"��*P��D�y?yE���m�Q˷g8m�tmظ��o='�n5�&۰G��r�έv�.k��=�H�9;aN^�Ѩ���o3�n�<�\�Z��`�m�@�=���R�溮�[���ลz�GM�����x�Ѯ��k���8�8�9:�X�z�{�\�.�n�<Oa�A�u�����űm�]X��:��v��A���ɰWF�A@����8n$d���'�vr�0�v�xg{vc���v�N�=��|Smۮ��ݱ���py9l��m89�ۗ@۶��Z���K!�$��+\�nk��_=qq\���t���q��͎4�<a����OFk�����g�#@��2Y�eq�y�<-ӹ籃3��8'ds���0n�����������''[����)aݺ{	�&N�<'Z]�p�9w,.�<Wn�ύl� \l\<��;26�b�r������`.���k������ui�c'NW���q�eix�=9գ�x5��
փu��c���R;ZޫoX�k�:M]v���N��n�;:8���u�r�VP�Źzwc���e��p]R!�)�k��m��s�֒�r�s��ɅN㛒��<����9Hy�[�����^y����z
���֞�r�����c�ݞ�p���,�{��zy� l�/<؇D�Q��z�^�;$�C�x��ݸ$w�Nz�.j��a�+6Y���������D�s��=n�x��up�7��#���GU��l��/u�z�$�\sS�H�I9�T퇳��TnR=.独Z
�3�e��6:#���f���� :�z�狳b��n܋��q�n�m]��a���Z%�k��$�c:�<���)�fݹ�Q�:��v�<�'�Y�mK�u[�];�<W@�&�Y�]��V8�J[qr�u�&������pmskYĝ����Fټ{��9�<q�e��:�!���B�ַk���@r-�X��6�n�W/u�!p��g�ֶ��.�M �����8��֥+��[�\��U��A���dZ)���s��'mm��]G���c���j�u�>�=4M]<��6�g��΍�TQi狳����H]�Z� CΫ�Ό�Ѻ�7[�n]��k%��;]��q���#v��Ŏ�=�]eĤ��x��e�����p�'s���q��umn�0�aIo����]�M�OR���7\�����Ʈd�P��G7�zt�K!���eM�&��n�cь�N�D�^|�ۏ������ԬճZ�I�a���,���ͧ1!\��
�r�_����s�T(�
�J�p��}�6�\:5
�߻�����m��{���AW^���D}�L�G�}����S*\����2��4j���T�%p����۝�T
#��O��ݵۏoϣ�P:�􏚂�D#\*�s�y�:�N�T*T*�wϾ���dB&D"�w����~�z��#�@��+�iM:Z�Ρ��P��y��z�L�L�p������s����S*rY��1��|����6���*er�2�F�����C�a����{����T+{����u%���PD*��"����n���a���2!{����:�B�B�D�W{�Ϲ�:����а����i��|m��{������ȏ�@��}���S�Tʗ�}���4if�Ii�i�N�\/����&D"dB&D�y�~C8��<����_]o�=C��
�o�{�9�P��
�L�G.b^������ʅr�P�T�g=�f��q
��T���3�U[)RT(�
!�M���
�y�8Ź���`��p,���V�D�f�h����x�u	��}���]w���:�
������y����enTʔJ�P�J���#�E�B#�~��w��M�}Dʄu�����P�P���}��ǣ�B�ϼ�冥um��)9�P��
�w��6��2!{��i�H]�ߦ`��#��P��slw�S�rpE9����]��%��^��Ŷ4�}��+�Ȯo����m���z��73�=������x�����B!��P�Q*�߿}�͡�Ȅp�5
�l,��6���
��L�~���١|�����y�w���|%L��㟈�ST֛];8��������hq2!",2�������q
��*�}�\�z����~ÈD�B�R�
���ﷴ:�\�W(9P�Q*Y�~ٴ8�B�S�����*)�D����|Qw~������{��;���t�����D#�ߜ�{{�u2�ʙR�Tʗ-��xm3i�J�\������~����w�{��8}��<3�&�eBم�~{��׸�P��7�k]���0�L�'��f��!S"ˎT+�}��ts�T7�g�~_V1�Ѥ@��_�z�ãP��T�XY߽ٴ��S#\����|�oxu;�S*v���/���������~sุ�r^��`���0;�W]v{[�Bv��萋�z{N���������b�->6���J�w�ohq29֦T"dI;��7��-�T+\*�s߹�:�L�D�xo������u��P��ؗ�w����r�\��
��g~�f��q
�{��e����r!��P��߷���*e�*e���:��~�~p�o����L�DȔ�T�����m��S+��Ͼ���,2�"�!��NݿA�����_q¡Z{睇,Ԯ��kUo0�;�T���ٴ�B�G*�T+�>�{:�P�Q*2!���/o�x-���q~M^�f��}f����n���ݙe���k�r�B��u�I�\��+U���F�f'՗ڞ�Y_ϳ05|����\?��p�B�D��}�i��
��L�+����C��;7���e��t�:xu2'R�_{����}��蟷�̧�B>���#�@AP�'�{�|!�B�eB�¡Z}߷�P�dB&D#��~�����o��}�2�����ϴf�\�^���mT�|p8p��<�px�BCI��{��(�v����{��>��D|�E����m8�2�F�T#���Xq�a�	HeB�O?}����
�y�y���!x�~l�L�SZ�4�lr�C۞k���t5˶�l�k����Q�����~��s�q��&����,���6����B�D#�;�:��P��
�o���6�\;�B�y�y~������"g����͛L� T��ʙZ�}�u�S��ʔ�^zt�4if�2ӆ�:��]���,����� u��fv̚>�*����-!�
�p�W�w�a�8���
�r���>���dB9�ʅC����[8�y��6�A8�p�����:m53��w�u����=C��������<�{z9���*e QQ�J��8��Ƕ�g��GЌ���52�F���5�P�dBw!�I���>����p�V��ǯ,Ԯ�*n�w�����U��!��&�;�}��~�W+�
�����C�T�T(�
�<��w�8��
 ">�*��A��uJ�����?������z%��n��A� ����3q3ۢg2��^���׽;e<c�����g�~Z	��]o:��T�euN�s]���30��u2?�T��r����{éԩ�,ߧ���hXi��ȝĮ�߿��:=L�V�T"dI;��f�C8�ן7|�p���C�
�i���èD�
��W	��{���:9P�������L��o�Sf��zO=����$����5q��M4��\�k��<qt�%2��s.��/kg��:����>qaݫ�����m��_<���:=B�[�[�O�y���#�*eK�S*\��}�i�N	S+�G6Nb���g\��_w�����DȄ����Ϸ�:��w�{�l!�����C��
�y��Nq
��s��޻;��xk̈G�~���9�**
%B�\�{��p��+�j2�Y�>ٴ͡#�*ew����io���]�������y��hѥ�4�NL�tJ�w�߷�8��S*2$��͛�3�[�TȄo�=7��]ԯ�����2!"�{����L�DȄCԩg|�f��q
������:m52"������_���~9K�:��{�?&D"g�p��߷���S+\��*Tʒw��6��"ds�L�V�����A��Ϗ=����Md2�i0�s�ohu��P�����R���Z��a�"tB����ͧ8�L�G.T)����������_�a�<D+���y���Ȅp��*e,,��vm3� T��*eB?����B&D���
��?W�"���t�����6�d6�WgF
N:���,�}�R�'iܕ�cY�l1���:�U��j㵔���:U���]q`>� � +l~kb� �FcD8�<��G�Z�uky۟Z�&����S�/8�3�9�'nqŞ+7G4l`M��8�.�7B荻0ݓ6����Sٱ��]�tF��]� �ø�;�nۮ���!���)�����^�v-;r�8�{=C�p�H�[����Ìf��z1�m=i��؛ض�`���$+1	��	��=���g�7N�=��nD�P�y����W�+��m�\ط����ݳݭ�����dݞ�`5k#���O}#)GZа���dO��߽����2�Z�P�RN��f���ʅk�B�����èD�
�u���g�ep�g�!w��~�� �\r�P�T��y�hs�W
s}���eGWQe��Cn�|��w�����D|t'��{���3���9���*eK�S*[{�6����2�A�������{èv�*2!<��_����!���i���Q�)�����4�"I��l�fЎ{��
��W�w���B�D�TȄp���O����s�u�����P�j2�ag}�i��
�������~���tJ�S��I�F��鶛6���W�������<�����y=s֦T.XeI>��6��'eB�p�V���s��T*Q
�r���>�����������'꼞�����@D}DUM�"N!\/�9���t�j$g*p�5
��{�P���*dB8O|���&GR����������ɤ��([��xm3iĩ�ˍL�Pk���{èt�ʄ�ʅ���~����¡Z.���ߛ�Z�?�ׄK�KUH�XL�F.8��r����ѹ�3��64�;=��~w���b���Z���=B'��K;��6�C�W+�
�r�_7����:�B�B�pJ�p�|����p�P��_��G<w}�ן��3�XY��6m3��S#\�����~}����Tʏ>;���]kB»8�������onw�W.5>D	���6��S�*-�v�T%�X����֮+NL�ض΍r��9������]7��k��:d�^�b�p��S�1ͧ+9��R����|>w�}dU<��C8��ʅh�P����{ÈDȄN�P������s��
��T+��ｅ�B�y a@G��W�L�.���KΡ��
���aרTȄL��\'��{���en9S*Q��&��|-}�T���D|��jer����{èw,2�)�W	������¡[����VFF�u5uy�d#> "w���c�w~�<@niʅr�T+����!�%B�q*��}���Z�L�D�ag~�f�;����jh����s�u2?T�P?"��'�G�Fy��&�a�6Yi<6���%p�����L�u��
XeI;�������^ޙ�:�p�W�}��ÈT�
��W*_�y���S"ιP�Q*Y߾ٴ9�d~~��6�OX��"�A�]Pb�[����=�m(�.���rprk�ƻ��,;�����a��P�#>�x���5݇�P�e�*e,
�>����s���TʄL�K{��6��"dq�F�y7�~��:��W=ƿ~�^���C*�*�ozB?@Eo��.�(��&X.�:�N�R���Nq
��W=�����[���;��� 2>�*�����shuø�*dB&\���}�i�B&G��L��~��y�܎������N��=��*�J���ߩ� ��\ �}��t�f�e�6]2��Y��۫���!��2�h�]/��������R��m�}�c��e����Y1軱�;U�����̿Y� "�~�� ��Yv�e�R��(���nt��&�W�}���ާ  uRV��̥~��q���.�ڶ�^�U 552�,쫋  d�s�)��ߧmT�%���� ���� ��X�>2�y���=Eo�߿��7�!��mᮅ��i|AR�%���.�^�V+�wE���2c�������KZ�*��W�ZK��mR������ ;_������3�hU�pJ�}�+T��"�7-�8r|�kѭ��y�Ā�� 2�y�8������XF'����-�
���0ى�%�H74���X��N!����G�.���o@ |fԥ`A��M�+�~�$IURPD��^�����Q��QV --��| ���� 7��w��(R���%����mf.[m�A�+ԁ����Og�ΕIlw��Wm�y����䳙Ŵ.�3�ޅ%߰��=��BMN���R����M�j��tó����$��m8e�eS��Wt��������H2���@��o�����ϣo��;(������Pl-i�r��z,/l��к�8ru�.y��M����3�P��$�*Z^=���:� oSa��:W4�����u_� �W��O�/aRU*�)��α�\��F%1+��ʔ����L��u7 �3>��t����Q����)L��yO}M�	�u6�z�:�ܬqP�zr5������ <Ώ(w4��I����p}S�˒n� U�8` ;��#�J�ꝸ��ߩl�̫`)ȿ@�dJj�%)��^լ� ��t>V�8o�y�� {�M� ���t7�b�������x�y[`�E���"M�e$z��X�'q�J ����.="$�(ul�U@�}��~��+7:��eB�^n�V�Ҫ�h�W�>|>�>���>m"v$�@��J:�����[��8���vj��Ľ\z�<o��汅��>��]v�՜v6��{������ܻ��t��/X�96�sɻ&�W�nu4�k�c�.7
o>�i�)��ʩ6�nL�㐬ct�������-qY�<���PWVx�m�uB�����	o{'c8�}�nI���|/�kg�7g��W,�\Ѱ�b4*A���8� ��d�5��H簮x�m�q����J�:,ϟ?��qeۦ&���ngS���|	�m8`]�Id�L��ݩ>=��G��oU�����UP�j	*J����dX@{q)~�A��+�:�*�^�:�$�*�I.��1��������n�p4�j�4�i9���M� 	W��ď����,��,���������l >]�v>�D�A��hTj�
�/��Y�I��d� Oݴ�@VmRI\������[k�k���J@�����;!�uU)����*��Uؑ�{M����sy�yeM�I��  
��IXu�7�u7�/wz+�3u���aQ4TҥR�\����mQ�^�ڽ�:t�F^M1��]2�|����dJj�%+|�i���J�*�� ���^{O�B�^o�i{�>Y�v]�eM)�����J���Zp	��WV=�?|����n�����ǜÔ���Ӌ3��q��N��z����Ǿ�]�eW`F����s����/@{�3�m]�h?�����}�p��UUO�7`�g��M�"s%�Ob�w��.��r���MB���o�Y�T� �_U� @�?l �[���o� U����q�W���J��UISM���X��Җ��<Xx��\X@ Do^�L��{�Mb�����$
{j�'�BS"�1U0�!��}V�~ަ��ͼΩ��^����ih7�V ��l @�z�����;}�q�?~�o��;��lT��:�}�+Y���sG<<R��vlG=��ŴX`��0H���6(�� ا��7��{V���>ަ���u�x+� ̀]WWb �:n �N��fD�h�4���Z`���̞W�e:�}έ?�����@P��@�ه��U+��I��e5N�6�nm8a�	�mZ`��y7����~s�}� �9���jn��F讽�LX��hz�#S���n�!���D�/X��z���^^�Mrת\L��:y?XQz�jX{�s���{YN����ynyrc�/������@�e=���@1P������0��'(Iw�a�B�ʬ��K+���0�񧏽�bk�U��^�|Q������:�����>�0��n��PზD���E�+=iCƟ6�e������j=�9|H����taB�xz�MNѳvfX�[��+�:"z@,���^�w\�X�hu����za�.sY����]���e�m\.�+IǛHپz�=�㗊ףx��:r�EP�{>Ӽc�����wW��QR�WQ]Wc"���].����/s��H'��5�]�<f���J���/��X�/5�{��I��}nt؋0ϯ�~�P���.v�ol��b�����U�>�}/2�&�U@AK�Ӯy��ƽ͙��dN��:����[Q���wz(�q!��{u��n���J�-�zރ{$y2��t��!�+�uU�|*mׇ:
W{&ٯ{�W�UN8���~Kh�w�5��A�&���\l
����Ԡ�}�靼X��W��X���Rzs��҃'�y{���M�0�.�1F]��X/0�2�1�J�n��_eȇJ몺�}r����0���-���Sma囏�R�9��0��1J�WTK�3��1m����F�Y�:q��E��:�<��'���w��c<|�*ʸ* �mX�f$�(�2b,v���F$�$`���X��1r��XD��HEd�ɐK#B8��Hȑ��*UH�ETU��F�G$�H�@d�d�VU!$W ��X�U1�I1���"F(�	�&*���Q"3 @f �DcҪ��
*."(�0���&
�H0`LG�"EqE�d�#Q&1I��!$��+\�bF(���aX�b�H����"�Kc1��Bdb*H"����\qbEŒ�+�ȱ+Z8�E"�DZȒ�Gɘ�	 �Ir,����0Yd�$�QI���RB
�*����� EE��D�"ȵ��H��eH�\dEŒ*��"D��0�D�BB`��QqLE221F�\l���#`�$�#	 �0fED�&,�"��dQE�bEbAG$�ĲRLŌc���V�	U0�[q��$I$����LE-�DT�#d�%��`����H�"����B�,Ȭf,��$�V���R0qȐ��ȹ$�3,���$�	�~��$���[�#�������T�!"j�%M�������!�WVD�U=�> �m4� 
�*����6�n'+����n �:��5H��UI�����#�J��qd�^4��_����N � y�M��$��������K͎�r�*�G���� �b�jμ�O3�n����ǃn3Й�6�Q{V�<�Q1U0�#x*��p�� �m6 | WeRK�G{�%����`��:����;��)�f*�����ڸ����PS����즽��Y�=�I�
�*�D|�?�^d.���} B�C�fD�hD)M8{��` %]�J�	�ֺTꚷ�}>��׾�n�p	 ���Wq3RH�&��LYU��}[�uS_v;b���y�H�>
ͪ��o:���
����2�I����`�y-n���dy�A��f��������<��^1��=^>���=e^�w�f#��퇴��}�������n �����MB���i,�>��>~�S�{��n��4�n��/~ �}M�D�ڤ�� ��Saeϛ�B�}t�����"eP�"J����GG���լ��i8�,v�6�쳺.K]+��w??�>|��7J*�URig�����U�W ��i�s�Wv�����g���� |�기���Hu��b�a Cs�6~J�_Q2_l�}u��J�*���7� =N2���/�Rq��T�R�&b�
i�{ꤕ��z��Ǘ�6�R���sܧ��@*� ��l=��̊I�BR4�{՗������� ��R� ���� ��fq����]N=��� c�����㉚�J"jjIIˀ�nէ @'ٵk�����> 72���w=M� ���L_�{n�O$i�k\n���{�s��+kz�^Br�)�|�Ӻ9Z��v7�x��co�u�uqP8�yiX�ϯ��H��|>�h��IJ6�k��q�J�1�;r��[�]:ys8�s�I���v��uɧ��*f�X4'(`6��Z���;��la�c�6Z{n;]V�]7n�m���a�ڦ���=�F�h�M�!�睑ᔁ��OL��\�6����0��L�c���j�9�����������]��<G=I�����-�ǥ5m�h���˫�7m���z��:n�iw:�8竮���v��[n�p[�^��s��n9z??�ٶ n�R���7���,  ~�U��'��nJ�&{q�����A����ܧ��
��T��M�o{�ؑX�Pzn���W�e/_�, ٞ�� ��U����u?uk���p��4yy��m#H6� �¯}V� �����u
qm���^�V� 3=V�`�oU�{�.��� اf��=�{yt�������M�@$۴�p�ud���;uX��^' ��o��Z��2)&�	H�Uϫ �����[X�\��D�[N ����D�%g��dY�w/5�ux~��k�
z �����۝�3�2��V���Rs��s���\g����.��?��d������%,��m6I��� .}�6�k3S�^Ej;6��$�i�"���H� �*[���W@��x�ד}�|�ځf{�wE25g7��t�B,�/�z�V��v#ݭ��}��Ob��}U�e�|���a��bљ��O����^^?�]UQ5O����T{�g� =��xa�FGv�� ����&
��5*��p��ؒJ�ʿ��  ];�u+~pz��׀�>����� ,�U�EnB��!U0�!�����"v��R� ��qbD��JI\�m{4�q�kْZ���V��߼�]D�L��TӀf��\ �굻���y�_���>~ʻQ�{$�'����D6�}@�T�(�ckm���&點���7��;t�n��zx͸0�qo߿���yt�3B����維?����W$�޶����_�T�;j� AFo��VXJ�I��j�1]Wf��D�T�y���Y^� %]�W� �_U�I{���>&��s�D��NB
�����RȀK�������.�V7�����򠬔�L�oS�Io[H��G*_�[�(��qp��Rx�V��G���?gy��υ�yט��O���6�_ﾈ�>���^K� f�ň�??��nz�	��j��T�l7�ꚪ���}��6$�����3�V� w����z�cO�I>ڻ
�B���S*�a Cs�8bI'��3�p�-vS� ��J��>����� }�M�E�*9i�+���_x�䈩y��'F=	py��޵�7g��/Yq�CE����}�g�D��LUA:�} ��W��v��8����B��M��5ӻ�#lX��z�N�5�&R��RR4���8b^���吥߄��^�" �w��	��n ������b����vY��SRMLMUJ����w6�0� O�i� >��)�rȿ^���U%��z��@w��E�T�B"f������{�%����/��۽V� �m4��D�uuG���T�T����)��%���3|,�Q9��P�c����}�6�T��u����Y��K'b��D�=�y=�����f�7E� ��!� ��}M����*�����������*ܫ�������HY[�����N{�� ^�'�{#o;=����w��vu����m�<qGB`݋�=k�����hۆ�9?��n�>v��ל��������>�~�l> �+:��'*������ٸ+/��@'��l=�YJ�(R4�b�6Q������|
�8U��T��� | �6��  U�L�U����S.fL+-抠�,��$JLU
U���k@ �{���:�^T^lp���#��m4�q �:�,"��SI4)��&��w�r�f{xb��n�N>�~�>  �ʫ�H�5�8���-Ұ^���/�LT"d��QU-���`y�8s�K��fb^�;=�� )��ŉ#�8|��L��q�V�f�婙�Ԋ��_���QnRZQ�w�K ۤ�d�ݵ��S�p�ِ��P��g��w|�M",�T"����7c���a�[��4�U.�F�";�n���	�[qx�d�œ>��<t��4�n5��k�D��/��7W-h]��d��:�ݾ�5���gA�y1�
��=Y�u����N��\e�v;>��Ŷ����;]�M��۶��oby�;vi�t1��۷=ɷ��%+�٬���������Y��Í��n��٥�q��i����.6�=��RK�W4n�O\wz]�Ln�SЖ�\�d�o\�;{OSʾ�D�^��������q��aTJ���^�@n?U� �S�W`@������\�©���7ަ� �>;�vWd-WQ*&UTO��aV>p��.=��㦧W�y� �Up ,���G�P���Z�z��7>�R��(���Z`���� >��D w�q��ٹޙU����INeR�d��߼�^�;��m�t5��M��ȼۖ)x�����X�l�9`} ���j���3՞�>���{ށML�LU(I�ݝnO���ڵ9ٯ��J�2�U� A�s�Ȁ��ҹW]*hȣ��=�D�4�*�9x���ܮoh�e�ʻ�k�פz��3��I�T�w�yM$3R���Z��z{�� ���$  ���R\�{[p�1����$��oW��P퓅@��e�n���~�ĺI���W�n2��$�K��)����k]�-^��pi6*�[�/E�w��]iNŦ�ۋ��BM�=�Ǫ�w�]Mg�]�w��bkַ�qi�� ���}�nBI�L�_��'	$�s���	�#^U�uAVDn������\�D�RUD�o��|��O���a ;ۨJx�?e��k>�]8��" �}�M���S.�LL�1U�p@�OvyZ	S�v��!����@��n  �{��ޘ���.�1�ʸ�η$^5�eH��*�IW=�� S�p��><$��k����4��)ޫ�����-P�|�!/̙5YwXY[�-���S�8�9Y�7bj��I5_�����%U*�	��%�����$���>� 	ުH����oz����Pf��p�?oSpTﴚ@I5��5R�^}Y _��HsW~�ޜ�$@$wi� S�Wb��*�ۥ^O5Uf�{�@��a�n�WOc�bI%=�J��$�핳��6���ڢ	���ތ��@��!Lҁ{�+�61�{,Ҷ�*in�h�+��weh��ec�������w�O�����X�#�"N���
�B��TJ��'�CaM�Y��xO��}Z�K&�����ꫀ ^�_>3ro!�N, ~�SK��)�P�&`���md}기�o�l��_�����u7 ��)�U$�����`*�N��v�pCu=���N�S�M�e�#�uv�X}�s����{Om:�8G�uؽ>�e����]�ʒ�JJLIV<�� @%>기����0K��J�.&��u4��u]��	UJ��j�	\����R[6�M��/=1"�i�� ��ʢI��yz�*$�rc/*���~'��j)D��jje��mR�/��� ]�F�K�̩��]�� �U�J$�~^�}���,"�i��Ut�?;3;���/3��>������Ռp�	�u\�ת|�)��k#
�)��Z�4ɫ���GekY��6
$��7K_�z��V�/`5�	���V�/c�ڸq�No
�&�yC�����7�UU'�T��݅�Ԩ�%TO���p�?����q8{0�03������I=��t/NL�+۳��!e�r������{g��=rc6�C�#.�]'n�۵:���0H��=�4)��ا��F^6`�+�g[� {�M�ѵ��U�^� ^�nA^�^�RI553IH��m6�IН�:Z^��V ^�c�> }�M� e�)pAs�3��O
wτ�/݂�M�L�Dڿ��yu�h���p���:�w�{��Kۺ�F�� ����D >��
ͬ
@Q5򚚙��)��"�1W�չ���ܐ@��:� �uus�:w���2�����H}�"XF�i��U�ޫL�]Wz}��]��u���X� {�M� .������}���L�~�����y&��7xG�[gv���v,X��y���px�k+8T��ܥ0�nLX�*,�L7��7�l��Vذ�P�{Fu��-rd��N�w���w.���_^��TaW��U6�MF�QtvA}�4�%�[��nǊ��w��=�z Ǿ�M�^yzm<7��ޮL�Vn�gULtL�z;�M�f�ug�}K.��N���L�l�HK,y`;�vM�u����znM��g�=t�圭-Ӆ������N�Î�J�{C�\^��Os��0+���Tk&�Z�lb����W������h�o\7hr"��]a�N�(���W��O����)s�;�:��a����\6������Nd��3�}��e;���%ҧl�֬I@���9�E�C^v}6`9�U6EP���[��S��$��;��4w��G��ū5��E�G�����A>�k�շyRh��XTr��O�q�렐�u��)q���L����o�|�,nF	��mc�v8ߧfݥ����kI�:�z�2[K}悦v�~�d��+�V��'�����2�5��L�Lqg���%{_M�;}b�����a���̉���dWY���(�^�����Li����Rn�΅�|Ҫ���{:�\W������:�
�w>���5L��RDs�腪3�-�vpާU�_���eמOngܨ_�$�v0��V���[����b�V�[��,�[_:Oa�6�w��
���oocmu9+�
2i=��ݠ�"m��E��+Eb�*���#U��J�S#�XB.9\������I��G*Ak�W$�(�#�"LU#�8!�H��� IPUc#H�Y!DZ«!##��(���V̩rL`��H�G2+��U�X�V3"8�#��FA�$$b�9r+A�QrcTd̂�.*
8�c�Ȱ�1�I�\���Q8,pd��I1$-�J�d�)2c��,qH���d0"�!\��1�U����ȦH��X3�pX�q�G1�r$c��1a�SL�! �21EDc�"�8�(���GH�A�#��"ȸ�2dpR1QQTED�(����r"��� ���I�dp����b����cEcUI$����"IE1d��
��1I �$X�QpQ0��Ɍ�Xa�+�
������I"E�U"LP���U����7��vGN�֣�̛qɞt�7#��*��eX4��h�5v�|�q�3�q�ݤ��gb��3�+�"=�b��w"����a��`��Is8�\�y�mW;+���%#�'��h�������I�f=�:݊�u�ɷ�:]�!p�)�������qǎ�T���Kn:N�c2�;��X=n{���ͻ,��]��}w�&�U�m�ధ:��*ݶfL���L�`s�V���b�p6�s��O�����ъ�R/kX�sPb��z(����j�ڛ^�F�9�ʔk������OӺ��:�u�D�;��B�n�N��e��r�sͬ�=�=��:|p�e�nhݲ�c����7m�:�'z�{Y���ʣ��%���񅾱��&�+DklR7W�ĨKu���������]g[��!�l���L�V�ܓ�����.��0�^\6ϊ�'�8� {z�ڶw��'�[c5��-<�7m7#�ك:��G����g��6ع���\pR�˱%��q���x{�;za���.��q�,#�]�nò��4j��-�;n��/v��0�1���n�vX8U�m�M��Ÿ���-+�(�Y��Ů֪-�g���o}o����F:�V1�d�A�"	[[x���Mk!+HĔ��GJ˪U�i�<c��X�u�s���1
��h���r�m�����q����'���u�3h���j���[Ѷ���۞y�vr�׃�����\�g�(#"v�ɭ�����k�2�,b%ͧY�[��v^�K�X�Y���2OR>�,��E�v׮��wn��kP�:{�6�Qz�sT�Y]$��码%Yƺ�N�EQ�re�>�=NOc\5��v�˃�����C}uu۔Uڡ�y�X���TvwK�:�=N�ǣ��	�[��p�҆!����wH<�����u�"�ֺ��6�Y$vKs�DMƞ#�c��.z9��G�`��3�ոЪm�9N���P�lkێ�x�4���ŜmtK�]��w��>�y���s	��te{0%�6�x�Em����㎸s钇�l竉э��:rc;�Z�u+gM 9o&lWn�D�uwG=�J���-Gy6K�6��W:C��]nm�ڸ��u��.�Ӳ��z�u:/h��v�{��rll���tVӌ�Q�*<v�Cf�%��n͎������vl�M��t!o<RZ�U�x��+U�&�A�Zڨ-�����1m9x��%�Zƍ�FFz�:cB�����ɣ<�q�:t�Ͽ���E��Z.H��w��r���y�UU^~l��H��P�ȶ��W4F�Q��r�Vx��H%HSa8n�[�L�\�Qe(u�8���>��� �]]W#���#���nbي��J�M ¨I}~p�H]>��� <�c�r3-�n�؀ n�����B�蠕@��Jh��e�&�Μ�2�3}�\�2k�	/ou8a  �˚� 2�y�Uffe��� }�vJŸi��t�4҄^&z�������ކ�|�q���InwU��H�[�ID��^��^X<.WYMv��ݎνZ�ph�`�HX;a�=L�	-�K�\�t/D"��݋~����$*(��6���|	B칸��s����P�������� �ܺ�v�cS��"J����1�t|l���͕}��9U�Rtw��]�5�ʸ���dCÏ�)���=�-���Q����Q_ǜD�646�t�҇�P�S�p����DG��7����@%�uV ,g���@1���������w��;hR	R�N�'��	D@��� #gD��q��y&��.�+� ������%��T�
�7U/��S�[�~�bӤ�J�l��>�=�\ @���w�E�00
���dU�Jh��e�&"}�싪�}�O�eY0�W������\ �f�P����@Z�)�|�:-������۷���קiεrn�fz��jވ��v�m��WGns��n9z>��?~i�En�ML��竬,g�à������{���C[)*{W����^N�nMF���S��U޼p�Gĕ�7箒2��Iz�zĴ����%�˘pp.��z���K�U������I�Pn��n@ �u6 ��;=q��[�D�o��C����H����3�ЭW����Ө�o��p�;n�N����A<1p�'�MU�!�Sm��\����kd����}��{�~� 9��q">ߺ����N�	��`����\�{*�_�)�����H�����I-���ny�+Ik����W�?J�ST*��C[ޫI$���"Ȩ���3o�Z��LC��c�">�I�$������ml0ʝ�K=�nqZ��&�#����i�ٽ���7p�U�S�|k����
���SB��4��x3vqÔ�O;jӈ  �ꫀΜꕝǻ#��7=<�� �괙���PU(SSI]�To<�&[������^[��-D���M��ꤒ�]�b���O�ઇ���aæn�{����ʥp	oG�s.��;�Y��� {�M�$@-����F�Q2D�R(7M��&r1]�T �������J�c��6��}7��f��X��S�In�*���e@q�Ѭm]̥�0����wF�w�i~�9{���{��s�7�菢#���M�ߢ.�S��0UD�O�]�Uŉ���9��f�� ^�o�  ^���$�z��E�����g��}�L�(&z�Ooj[V���q�[��I��A�O��`5d�߿߾���"j�3Ӌ��ˆ ^���H��1�o*�W���7�-� k���m�:-��b������۴K�MJ	�HOV`K�0����c��r#�*���x�Ӟ�5���π�՘�PTRSSS-�~꿬H����� =�9�{h��˟]K؀ �ڸ�hU�/J6=��a!L:f�K��Ni�f��[� �z��, #�+�����s�9x~N�YުW�G2�BI��P�SW=�$ �ݖ�z�Jȥ�O��[�T�� �_���$C�Ζ¾�*�����I��ݹZMK��rf�͏z]�D7��O�������o����3���]��Y����HOb~�l}���x�z�K�������[�謦� X:�j�����Z��8���sr�dG&�-�[b��e
q�l�-W+۳5�R;��cnN������:�'Ti�"��t���4�/���lYIL4�9����;,�e^����vw�N#��ݐ���1�]:v�\��T�{�\�^:z֭Ӊ�0V8�q�؛�v�m��X�H�:���"d�MZ���Y��	���������qyƺ�1i`�b�v�=.���m��xu�c�����������WL�PN����\X���[� �t��+*.ݎ\�n�+��$���u�W�?J!R)��Csے�D@<�u�V'.����|{'s�������� �w:[� �)��7ʸq"����Jt[E�&�;����h3:\0�J�[�a+�%>�*�z ����$���iw �h��U%552�{=^/|y�� ���� #'����KyҎ��7|�]H�� |^l��C�v�銉H�*���_K� @%����:r7�v^4�d�'α� '۲� @-�Wf_���ڹ�?�7���qu�s�5���v�Rc�غ�K�:vڧ��(&�!��S�ѼTH3SJ~
�>p� 0��L 7�U�g8����^�\b���mȏ��wM�>�}e�b�J�lR�U^6eT��]�}��_��5�Ӽ]i��u�t�>Sn���cW��A�I�̛��2+`߻y)v��Ru)vb}}��+��|>����� ?��i8��uv .r/����:���w9z&��ץL�"UB��}�ؒI{�\X|����PFf�W��g�=>��� [Ω\)��B��lm]Wo���y��������Q4e�$@�T��/>���F�s�蔐:�� ��"�U*Jjje�Or�"� ���'�1�N�-���ή����q%�ͺ��߇�������߮7Ǯ;���-��Y)��묝�x.��A�Oe}�I:�=I���χ��gb��Ϟ)ג� ���, ���iUS�zlۢ�f� ���D6�1�"eS��
�<���O�HU�y�O�����0.�U` y��Kjŗ�^PB�{Wo��u�MPj�i��-�������r@n�'���-�ydȪ��Xޮ������n��K5���Z��eɋE\B�{aY.�w�>�lta�����].I��j�#�'.���I�����Gї����@$��]� ��?���W�ץL�"S������Z|�Y+p������W1� t�:Z���.Ձ��������L �$�'����"gM�ߖl'q��s=w��R�˪J��N7" �gKae�y�~|�o��-�P�2m��z��kC�<g��k�u�-:;�-�[uP6������݁�ٙ~����� 2�<��I>Ζ�g�~��0�=9�����"Đz�q����;��S�����5������L��'.�ŉ����=�6�)D���c�黇��J�<:S
� ��
�����.=�6�a�_�Nfu]U�	^�7#�:}�-�{�^LT���*��)�	���Tye��C� @N9m� }���n �>�겶��Q>q��ǖo�;�oo�h�'8��-a��ι��ed���ٻ{��~���.�j��z`�슔\b�%Ԕ��	uO_�����HOw��9d�{�;ZIu#+�����i�	~˫��;=	��w��a`��$d��[�>w]R��S[���O���7�~�e�&��BҚ�W�b�s��y���dkX�5<݂F��??�?�g����+岖nO��$ {�[.몿�ܽ>��w�d�*$�s���>��n�����"`����e\X�����mr�!�@t��[�H�uv"c���{�N}f����HGUuw��4C*�wb��b�����s�� ��O���oЄM`����l�K����tc*$DĕU�����9�T��M#e(�� �(o%�,˪J�׳��\�Mh3���~�SPh&RA��;6*��0UP�����v��n�s�su�9o%��K�U�b �盓����s��f��
c�*wwJ]5v��U�[[N��x��3�S܏o�nv����0�����F:�㌓��ő3�F2�z�˄�v�T�T
�r�����LS[TƁP��	ѷ�m�:h�]U����\ W�=i����Ž�TGC{s��q&x{j�ɍ�O`����/����Kq��c������]�x�T�-��)��RОZ�z*]n:\Z�Zy��S�Z�d�Ӎm����P{6�b��\u3�w%�XG�Mݑ9�3��W.Ŷ�r]}v�[g��[t4�t���dИa�l��-�p'[*Z�k���a�x6}.4����n�y�=2�~��L�&�����{f�.˫�랱�e�ɸ��>�K` 6��>]OT*�_',3�q���x�c�:V9ߘD�%�uI%p{\��6*����v���'i��6I��
�����R�1�X��={O�X�<eNd  .뫋���uV��!�eSn�
k��8U��R5�a6@UyW  �ֱ�Dt��_M~
��{u¨�=�J�<:SRF���An��p� 8�l�d�-}.�`��3  �ʫ�7\�r#�>��l��Y����P5c:��A�%6���(ݗv痖7O\�;��[��4T�d ��5�.7B��{��QJfb�j
��{ޫ�����r����n�n�	�=�32�m�؏�=ޝb���̈&�&�"�A����`aZ�Ի-�~{x,��M�(��לt{����]���t�׋+�v�m<3�`�C>�b��E���$4�5geߩ�������[�π M+VDX|�����}�}�e���x��p-�W���U�SB���������� ��Lq�"��xy���@�y��D@>���פ�H��&
����)y�K}u�y�L�%���H �f�p $���f��U�
UW�Wv��D4A�SUVʝ�H�캸���Z�ɾ����?�#�ٲ��D WU�[��A4W��
��4�:.�M�i0���N��F�ƛ��x��{X1�#=@�kc��������@bSW/�����e� 6k�o�ޗ7Na�}郯��$���l� Dv)�1DM"f�UA-?���ݙ�f\x����9#'���$@i]R��w�k7���U����9����$D� ��!�K}9�x������Q�R�NGm�}YI��j�M�%&d�Fy�~�������g�,0��0�&[s������no���$Ӽ�/��S����L��y��r�j��G�h9X��ȩHO9��:"�5��#"��aI
��վ�X�فop��u_s�����N�j�27������7y39��7�d�޸��璎wn��-�j�����v:�WZ�$*���ɜ
N�v�}W�jE������l��j��^Н*i�=)Y�!jrˈ쥤W8`Y�Ŝ���M�#�g���ư���]�~��{x����˕LY�:�Z�����f���N�E.��}��ȧ}v{���~��z��/L�z�S�n4}��mZ�k��D�v̺3E}��b�܈�D��׆j�&{̥�?�5w�%��Ζ��J��t� ��kmU�0�M��DL�'O%��+s��ιxf�!�o�7��x�U�2�<,�3a�\��)���w̻!�2i���Y���s5]�Uk3����9o*�Դ�_,�隋���0�,u�[��b�V�İ���6^�z�W��EzЄ����D�04M���������˔V=أ�V�� �]��7�?e������������L�ǒ��u��P��7���P�%�җ��Q���XH����{�ZO��ن<;=!��O��_�{\����ݜ�1�õ!|�ɥ�8w����9�	wD����Z�\����׷�N���;�M3˾J��g0��/d&`�w�H�H�䙑�qEQ�A��$a�s9#I"*�"
�".F
�d�LQH2�H�#�E�8��E�q$D&$`�L��Gq�����$H�,H""��$�(� ��1�
()����WB,�WB#�b�X"�
�QdQH��LU\QTb
VBD��.(��$��ER1#1r*��#�8�c��c���D@\PG�����EE21�d1U�"�⪨�8��Ċ���� ���`+$��F"A�$b�bAqE#��AI20�EULU��dqI����$�������� � ���n � [_��]��n����wU��
�.b� g:���+�� >��g�zi�n��U����o�>����(*h�������$��Ǔ��ǳ��ߚ��q A5�M� @)ܫ��|/g�^��}�_ϑ6�.m���]k^ٰvnt�&�a3��{lj���ME�%b:;����ߜ��=*))�����$�Gee���F_W1)����OUi�p{��o� �S�T�Kcl��&PU*�>
�<�r�y�9]%+�]k�"w*� ��o� ��G����Rqڝ9�"�5ETL��^���� 6�u�  ��Y7�I*w\�r��Z�@���� c;��W�x�L�H)�HbU}�c�w�-�̯�+�Φ�h�) �9�r����΂������r��y�U�-��n�*[�\y��J&��"�Θ���o�ɞ�U��ڠҳ�>�"f�Ut8�7è��^�������+�w�~�>�� @,����7�E*��A_'N�����i�ٲun���E9���j�>1�������G�擟���M��$Ѩ:]-MCDĞ�����]�(\j�޻a�Y�vw]�'V�p������7n&"`(��@'�W`	c3n_�{�V�.���/��w�W Y��V_[$�UKm݊��k��b�\��{�\�, ���㔘{��I7��B��/ъv�"���Ʋ�"
���U����?wS�a� �o��^{Ҫ��U$�}3���@=�;�U^�n�t4�e���G׍����>&���v���}�V� �S�ez�9�MêԪf���Q}��̕UH�*/zq�	z��,Y���<�W�U>�[6zo���y�M� -���9��fC+����3��d��5|\~��[U��}K]�f�F>ʭe��J����޿v�W?/j�}�m���R~*S����W�����{�scW���ݟ�A�ms��/h��e�E7[=�Ǭ��ӫ�ǭG�7n�������58�Kc�-U��mМ�']v7]r=wK���&�<X5tnMz,gd�[{]5M�=F�������H��lt����.-n�O!�ݱ\m�n�(z�WV��^ƭn��rq��j�n.ms��]�8��`���;m�qquCѴ<��i݂��2=;y�{�Q��e�r=��S�'���\�4�����RV�{~�����n8t@$�nӆ  muU���ο-&y֩�.܈�n�I�{^�j����
(l�U�a�J˄��~w�F���� <ͦ� Imu\X��7>��S������Fן��)��%�瀣_e8a ]YW$@GE+Q��}�]N8�x�$3i�����J���"
����V�޺����p +�t� D�U\@ �yաU��5�$��s������TXt�a��i�-~�� _N�=�G�ӑL >���� Y]Wb 1��q&�NI|��돳����M:���K��h]*A��v��G��tm��^��=f���n�������eK�J�: /}�� ��j�#�1�Gy�ɫU��y;>�i?���vWM�U2T�D��t�Μn@�ʞs��շ��/s�쁰wsףF�<n�w��6�ͩ� ��u%I�v�\up��c=��y���2���?�3q��܅�[�����}�����%� �꤮ 2�7 FR��];��+�u{	�"�jb`(�����`%�������9�5��=��u{���ʻTl��c�g�S%Km��u�_s�˿���\X|��c�H�S�k�.}K`^̪Y|.��PIL
�*��r�'����M`�� 9���  �zq� ���궹������T��j���*1ֶ��xb6��ӹ�;bcpl@��Ohmq�����`UUEN���T�|�����" wSp��(���݄�긡$D��bqe��*d�j�TJ�-�U���^��=YBD�oz�����߿�p��4'~W��=JIB����nH�O�i�� [ǖ�/UYQ01���"����೜��؂�U&W��4��7�����\-.B��Cv��kVɯ���d2t�y'�ﾧ��O�������D|�u7^W���*f�&�vWnO.�y,����o�)$|<ަ�  0뭆��s���� ��g��G�oiR�RP�ER���{2� i�W�Պw���Ϸt��1�D@�6�� ��Y1r�WZ��2�Ȫ�_2�LҤSOvA��뛌v���6�kE�
���#���}V�������<,�� Y�)��r|����8` d�ԤN2<��S;�:��q" ���l����TUEKO��ޫ��	�������ِ��i�>�î�(Io��L�~�w�>��KW�x�S*j�J�,aoz��^:������O��%��z�x O;��@%�G u_7�)�Ҧ��4�6˃;�M�'RI,�u8`	,6�n �>3�<���f.�Ǉ3�X�G�u�|��+�Ձ�s��د>�� V�]�.��(.�`�O��0��"��;�{���
����KV��u�M���{I�"��E*vU��fzy�C�O����������w�괒�uP��Yؽ,*�|_���"O*��l��o�(6��k%7e�jlݲ�u�a�@
��N��6�ܶ�OϿ�>JUL�J�J��|��i�KL��@ޞ��yM��nG��u_@ i�R�<�Z�*d�TT&�
�<ܟJ#�yu�dT��nn;D�B�lh�N�צ�5T��w�+6��U^�a��uJ�(���nj"��2��> )��ՑQ[�����	uqB 3�<�HE��x*&�B����mONZ��p��i� /�P@ F竘���ɢ��3Ն����T�ϝ7�)�Ҧ����WIgl�Ð O;i�s)=�^�g�����Sp v�y�� �i���Xw��\Pa[�VG5���]�{��r��O�(>]��.�i�<=��a�������#���c�n���H���Ut����uce7�hcO�;>ׅ�8�w<�Ɋ��=�h������/k޶�g���ԛ��rw6�R�n5���ִ�ӶI�mVl�qc�,���]D
X�s%��М]�3�H^gC�J�G�t��&$B8pu��r���ͶC6ˆ�����ݭ��ݘ�G�vl��g�h�o-��x���9�e9N�n8{��o���}]o���ڻdyR㖶��=�m��n�Ѧs��'�Ӷ�C�g&�����{���ET��C�{*�H����) >���ϧw��h��Y�7W�P� y��'�w��532*TUSK_z�%��|��<�1�P oz�� ����o���/����R����bu(&aMEAn�ο���}�N]X?]���.�@� �zq��D��:���^�ETT��U*"��Z7I��~8=��~�����ܐ	'��i8u�;�ٹ�vb� �s�ĄE��x*&Q5�9a}�M� ����X_�ى0���SbN ��6�@,�U�VL�<>��ˏ����jf�j��D�2�_�g����gF$���,�	c�����s+${W�N�r|	'��p� �K;�Vջ���ݦﲛ@>ͦ���MA�`��u6��s�J'MyY���b�/��ɺ�;z�r�W�fv^�b�v�A�o���٥���)�}���q�D�"�G`��vYF:E�6���bӧn[������I8��es�NY�v��E��xM�k�i��]6窹����>�=T����+sd�::yB�V�  =Φ��Yή��������Q��r��י���Ϫ�u�O�Iv:��  ǽL}eױ�����5���5�UD�(�UAZp}� 5��dc�K;{׉oǼ�H�[���@,{�n>��'�~�y#�[̤�"�4����JY���|u�]i����u��(u�]x�j�����w�NI�"��JU��w�  K��� F=�i)��63n�׆�E���� Y����k
��f�QE|�0����;}�o.q�e-�mg�  K5�X$����Q��U|��dZ�ӷ�	�[�ZL(SJ��Z�X^uZW�{ҽ���>��5��E~�����!kƃ�u2��4�*�S�s&�j��7\G>n��/�z�<��~�ʃEz�搸��.��ܧ]�@ .�Wb 2���#�*pE4�J�M�'����G{�.U��H�>�z�,H�/:� ��U�Q��)����| /<���ʉ$�U*���S{M�	��8dk��'1�2��~�J�2��������(M�R�oH\�*bJ"���	������Ů�	9�M�1��Gcvn�ѻVۏ�����W3
*UPE\	��J� �ݧ ��i.=�M�\�g�x{�v ���M��sQ�RTML�(r��1-��j[�`����u�[O�?wU��~Z��̋�l4g�"�.�x��&hW����l ��V��G��'���z �N�*�#�>/=�wUK�qLSt�˫$�����m(�s�M�8`y�V� wz�3!�ۓg��d����Jdd�.�������yg�Ο��R���!ݷ�J\(K9�sF��j��͠��^�u=�U�z>�oݻi���C�/ܒ�;/��޳mJ����(�*���u8a�^�8&z��kȔ}.l�H'�o���~6}��%��i���HS�T��aR�u�k��F��c��V��b��pE�ݫ[����0R*�:l�>I}b�đ{����u�b�vf{s�ۗW��w]�&��b{N�2 CE����3ן2	Ex���W);�|m�煒A?�s��E�{��:u���7/4s��2�����L���/{$�t�rI�Q͵+��5Պ�I�߷����d����N�uEӧ� ����p2��	���b�}������.���+%�O�5�)�H?�e����tg�@:��_�uY�σ�o;�@$���'�����:Aj��`��xU�WLo2S��n�����j�nEZ:����=�ܝ�2ޭkpY;�F��6q�r�އ@*���Onm:��=O���{�;�8P"^�4yq����e�8��>�S��7�.�mꇨ�X����H��[�T����'�~�[����cr��t���V0����(�:�qж��I���{/�vΊF��5Ȕ�G[�^=��%���� =����x�D2�p�92�&�t�CZ;��c����ު���t�'r&E����jc0��l�Q�Ovާ��#���c���o�w�y�uS�n��Y��c��7���x�}��U��[��P�:�#�쵳-�:�nZt\9s���-b���_o���S�.���11*�TX�_#�̖{�5t��UK�#q�ʻ.�/*�GF�̽��w_U]��\�Z�y�����j�N����%��*��K������?h���"�Pwn&��=]�~*�t�Ֆ��8t��a{����M�G�q�;9S�/ת���>}�a�yeQ��cN�ͫ|�E�b[1�3J��(O� �ֻd���_4�OV3"�׏GZ��E��K���{���M�d��:���4��ؾ��-����.��3��ҏyq<����������ۋKk���+?)p�{M�\|���.��Vن�ŀ�^�7��h�p+ڋ�ns�։嚎�*�k��}����<�.N�]���f�G�%i��u��W��~���Z德9��j>��������|a��ξ85Ջ��Frb�dͰz���.�˥������xJ~z��'W�����*�E�I"�*�& ����\EE�F9�E�$!!!"Fb,pd\]�Q�T�&!&DZ� �"����1����\AY �9$�\H�P���$`�"�86�.L��`�H�PK2؎,r+��Ȋ(��$��\G������"LTl̒LDpl��A��̶.
88�8"��2�EJ�JČDE����3�J�q�X�DE�qh�qA��$DpH�AqGȨ�E�FىdQEU�APU�$B"�a��#�1\J�Z�Ue��رr9,"Ș�E�QbI"⣉`��-��2�ܭQcnL$%$X������=#��������k���+��v=���v��v�ڬv���]v�j������|�\tY�`�'C��u��;D[t�Y.�y��rp���.��_��~��/�v�r��NxK׫<�aC�:�W:붞�cM^:� X��ܠZɮ�p��-�Ss��H�Tm��ݷ�����*�ۣ8I�8�;�kp6�r�3Uqȧg7g�S�]������s��;sv���j7�=�>^wmpe�cq�Ϸ{]��iR��K�x���Q��]�)�5�]u���k+�t۴s�:��j{L�x,��YS��o��:���[zL{���L=���<�1]��o-ۇuϔnx}�y)콰^v�Z��%���p�]��K�Ίp�ݰlq�;��x���L�z��n����V#���*��I�=j�G;T����)Ml;T�pL�=V�9��g��Rm�B�i��wK%�ݞ����v'����vwvH�Z�:Kz<u��J�tK�֜�wa��k��y���{u��9�v\v�v�Xms�5v+�v�J�y�W��g��v�̜����ɯ�?[v_��Q��v��}�����\���>��6��`������I���v�;q�%�n��l�����a �mv#lvǵ]����[mʧ93�q�'����"p����Nͻ'`8�еq�ݧ��[ۂ8��Ό�g�޾���cv̊j(僪")5Y��-Ӓ���N��,�gbv�:�n��Z۩� ΃T����rr&��������4r�Pu؟F�\[m�����e:tLp=�Tz(��ڍ�W��[���=��s��ɻ��vÝl���Gn��mێ������ط<ή0{n�v��+��b��\�H@Wln�y�s���k]Z1m�����SРΞ�i0��ӵ�N�u]���w��s��:��<h�O���ރ�f���V�Z�YSζ�gn]�(���8��|�2���v�.l�e0x��!R6�0��ے7c��q���������p��j7Qsڅ0]І:9m�c�[����\���z�R�m��;;��+���َ.����c�<\�Vr��8��$縜�[)g<X�<bxK����kX�n��M���!��4)5\nN��cx���7<��Ž��K��FB��勵ٷ�ʞ:ӷ��n�d��<	ۆ��-�-��ٍ��8��\��n��)Ijځy���.@llu�^��]68��/���θ{�&�Bj0���t?��~�ߊ)��T�:n���뀒N��(O������/�g�p�Gٺ_[����ݑ�d5Ҙ($]6�0'�엛�Zޡ�պ��Wn(	����x�;#mR�W���O��XTh�P�{�p�o�Q�u7��o��ƀH>9�����}de4�S	��uA=�t����s�BI36�� �o����%j,ϲF��S�MQmS��������"���Ʒp{����e��	S�@"����}�p$�]t%g���4�@���:�J�Y��*xA`��S�ϲ��cnu�"sn8t}����.ȿ�e׎�P6nt�A �o�.��C�u�<�7��l�d��H���H�u�QM4��L�w�뀌�D����oF�̰��א�]��̺�w=�]�:�V��x��G���^=�����O^+ʱ�+!��	�פ��0�PZ0gjͻ${�a��I[�0y�8	7i
�~>�̆N��l򅂂E��f���7������	$��#.�U�"�v�vT��A?��v �y�p���f2 C	�A�٣���g�;j��c��Iy��I �s��N�^���| ω{nŀ�l���*a�*����ǎ_��Ul����#�@�N������$a���f��]�]����?|ԝ�YÛ<nz�.�V�`�Ƈ���{[�.f�4UM���󺘦�j�e?�Fn��'��s�N�(�L}�U]D����e�$�y��Ƙ���-�P-O:�(Y�~�}�����$�y�__��__�P�׍�:�3���y�	}�s(��IS�i����� �>�P]x�V��?/O5�y���t�m�ݣy��z�����P���i�!�����x���	�ˇP�]�mB;���X���{�}	'ٵ������.Ǣ��§H��DR{露A�Ot`�Kp'+/�|A=���!�?�'}-����XTa6�:����O���u��K{:+��U�DVe� $3:�_g�������r���th�\Pmn���Eu�;z�Ǯ�-��/b�J9�;pum��?w�u:T���U^�。G�t�A���eW��p��^Z��zg��L��=�{4���lz��o��Wo��8	 ���!����E�S�����S��1I�T�-�P=��BF��X�	=]���.���%��I ����_���#�묢�t�j�M��~|:�1�H"l�BH'�g��׽�^�{=v1&�|}�}K[�i�ҩV�X$Et���$:�^�ͅ��y���&M6.�����PoJ{���j�SCŲ�����_^ۺ��Kݒ�m6,*t�6�0�7�����#su�g1�M��_�BQ����$�<ޫ�w��jOb��n���.��Gl�a�ljK�M��ۊ��t�.�����L�B�=]������;u�'G~"�dH:�:�~$���5WM�_��#�.	8��a�]:T���UX_{��W��Y�Z� �3a$��ٷdo}�!7���ra���Oݎ�5I��V7z���� ����LH��`��jh[�p�q�u�ĂM��9�h�b�?�e��7�2���ޑkˢ$�zm����9� �3��̾��ǵ��36zŎ^���4���A7w��p�A�����1'���vd$��ݒ	���?Hο:�m�/]��>��m��⬸X{��=Ys4�Q�6��|]ǝ��.w���gf��,H��x$j��2z��/Ws��8���+���o��r�qn,=��k,����僝u���J���7=ub��O�k�VL`q���`�̘��Zx�t Us�!�Wk�������n�7�9�.��rk 7d����E�q�V��g6n�a��v��iS�llZ�;u���؞�g]�l�:v5�Q�np�Nw�_����	�&��Z��n�g���N�ѧ�{;����r��]n��2�exc�._�x^2Q�&9��7�]��%k��@Z1=�}U�����|�uِSm��|S����H���|I?�~b�I �k佾�o�����b�0�T]�^�p0�����'uN��y��$�3��|x���z�����:��Qh��h&UT�cx�2H1���,��^��~$�o;�A����K;e'A&"����n��bv��W@�F;��~�f℀O�=�ۼeJ�d�]XÜ�����Ѥ��iө���f�%���b�ŚW�,�ʴ�(>=�������{�AT/�x^l��2�}|
�ި��t]U:��H8��`z�\�q�.wmyo�e�aW{���M*h��M��x�H$��#$�{�w�^��^�o-�����I6}�3�e�G�N�m�`9�񗣽����W�Q��>]o9���W�͌�ݞ|oY'6G�}�mPY|e��ݮ�s���%�@�8��f�{�}5�Qq�8�r�O�> ��	���ݓ���nٙ�(��^�)Y)�AԳGّ�OvݐH6P��"	�q�g}o '�O����[��0SF���UP���3^J���_)�$��l�I9����'�:�����@�W��S4��h��>��g�A��>"��-&+)��=�P���'3��6`�e�GG�Ӡi4Ixbc�w`nU�X�c�CK���Y��l�^�I"�W��-O�O��:�8o6|�ă�}��~$�{��n����	#g{lX��i$ۦ�6��}�ph{��eb���4�g=��A雷`�	3������Ӭ���WV́�_S0�T��f�u��7=�	8=sǇ�=�}�H�@�u���{ރ7 ����z��L][����V��AL���tqT^ỗ����Uv:�Im��I=3�vH'��c�vcb��M�u4>�O�c������H<��X+�]�꿒K���{��I�|*��qa�F� �*���� �}��۷b��A���d�Ngy�A{���H{�1���5B�h"���i2U3���U��ۂ�6�:��8��3���`��;	c�������'L�"�on羲I�� ��?]w�@O�곯����`���y��|��i�)�t�i������=���a'=$��! ����5]a�P�Az,O/	�ڞ��m�t�w`���A:}�$]|i�������Ēw;�|Oăg��m�G��]�l�OܸU,�=�`�xG�1�GĂr�ڡg{o���OT�����T�H�ppEf��g�h>E��3� Qr�/z�ٜ�Lm�sec�#jj���U
.����=���G(���$ӑ�~=5�H�@����fO�d�z{��g��{�R���{mρ ������~�����ovNYI@P��Wɖ��t����䫇�����(��V"���}�m"��L|��! ��l�H��m�s���;>33'�M�n�~J����SeЫ���$GU��ڔF�c�~ �g�O�;;�/�~�~;��{�)��M�L2ۧS���A ��l�H4j��6I���~$�n����ݓϪpM�I�M�� ������������D�1�	�۷`A�����V�ު�
1�@�_T0�D�[m�
s�ş�ۛ�	�����d �Y1O�7�,�����]��Rꧩ�>���M��I��K}:n��q�������<�.,\�|�=��t��uQ�4R�f"��ej�Ʋs�nx��Z4Ok �q�9�i��t�nLG�׊Z]�u�s��h���:;�.��Y��m�Z�絋����s�q��v��W�u�sd��YV�+�&�K�mŮ���,,�SS.��w���C ��ӧ�����ɉ��:��wZ�޽{���KǶ����a^"�u�O��5ۑvn��'g�vP�s���;���rT'V�A�JX�Nź��Ɛ�p��J`8DҲ�kAkv.��cn�L2��$,��y�*��[iY����� ���vݐH$�{��m�hi��W�� `�齶,>WCH�٤)��;/�
h���Y^�@���d����9�%�Ј����`��Ŝռ�*��[��t*�ܝ�?��p��'oqaT��o��~'�ݶ,����'�|�4S����M���*���vM�����,O��p�l��v^O?V��C{�w�?y�O"�RM���j���� �Q�Յcv~��EǢ� ���`�	9�� �p��|��<���H>����HC�����:6���#���{f��=��R�ª0ɫ�r���J$0�l��;.�$���$�FW{T7W������t��� ���a����i�]�Gא3��X��S;��p��҆�fP�\�[ܠ�Qsӯu{1j�ۻ����ssP(���h�B��H��|��Нs,;!�9�ў�YB�A�ד��$}��@I������<����e�{WCH��R��ӱ����I��j�&w�/���|Ggs��A����X��
�n�eЫ�{}��c���$���H�gj����wm3o�1�t�Aվs�~�ly��e��n�O��}�3� ������^�I��m����H��˨P�_{�������2��|��)�O���C�G���gs��g��.x�j�Ps�(�"������"�RM�M�J��7��O�`�	�����\/x�j���:מ�I�۪_��0�D�m�c��M��d�9r��y�$�OV��>%�g��#�.��Vy�W�o�9��[�QtM ��>���K�g]���}�7���`���L�	-K�=e:9�æ�_Ar��������ܗ���"ɞ�Y����ᬛ4��M�f�����t	U�cFtj�9}l����û׷�WYԻ��I[u]^�-�� ��j�����I鏳��z��݂�]�U�����h��o(-H3���a]Чm��\�\U#�h��f�C�a�%���z��dW�'�ݓ�U�x����i��7^�aq�A!:����X�&w	y��
KoL՚b �y
�pѕ��6�겡�X�Û���=�ğ���K/��X�ON�Tc��	���A��<���%�uq��ry�ON3�Ƹԙ��R
	�lvS�Ď]�^�ӕ[��%�[e�E}���9�q���>᧗G�Q�R���ɓ��싥(O�o���l�6����vD4�;V���h�قU��m�n��[������k~��>5��.������֫_M�QB��<��f�M��|e��W.ヹ�ߵl���pJl��8�;�۵:,�yI&�S�ã�ά�C�Rǣ����xK�V���,�2��]4Cnf9/�ؿnFEod=�h15���J/4�3�;���rr�$сδ�t�Y�+�~�Q��´{f,{�1f��f��#ݣi����*[�b�L�w�֕���
J��b|:7�]���Wx`}����}��E��㞱i��� ��)�Ub�M�Қ�c���ݾ�)���U�-m����ga-r���vS�v&ńJyҭ0���P3^T�{y{B�^�||8ׇeL�2H,��a�Gl�ₑ��RV��PPm�VBb[k�cEE��8�����A
��q\�X�r�F
HDFI%�*�-��\µ29�!%�
��\sZQWk��EQr�DPdȑ$$ĉ�rH*�AUU�H�c��REQPPTU$ �(�LY-2V%`�.�G$Ȋ
�`��fF$�ETsEsŲIs1F@�D��B��$��,dU�"�2@��b�@�D\,���"�L[m\X#$�"8��eI���,�2ER8�U#�&W8�Lqr"�ȮH�Q�Z�#eTV@#�D��I� ��QQU\D� �0lm�D"�D�pbET�L$�UDY,`�8�b���TE*)"��R1�1�aU��I&��2%������4PIe�|�$ �W/��ɋJ+;���Vψ�i�t�`���s�w�W"{����2F~�K�g�� _�ʷW��9~��|F22��*�J���t*����@$��p�U�O>":�h��	7=w� ��y��|������*���:&:7i I��k�� im%��e�{z=%ܼ%q4)]�Út���:��y���?��v@$r��>"�����6}$��C�g]�@��g�L�n�Wf�<� ��s�J�R����~$��ͻ �2��K�bi��_��YYq�_&�a��&�3�޿��A~�>$o¦�:�d����0��g]�~#/��&�6ֲHL��H:�4}y�x�M��V�8�K�~�'o��O��p��c=����G�*�>�ڨ�;*�4Ҵ�Q�����t��n��I�WnN�,䛢�7�U�-��磇��Ԩn�x��Y�e��s���#���U���T�%U$�==�A'��`w[��Vk��i>�˻���s�I{'��{Ѕv�ޯߟ}��ƹ�][�2J$<���=�l�c Tz��h��G[7[(�%d/����egG���vu��3|� ��� �y�;MN�3M�Yv��X���	��kM�lSi�M@xߺ0}83o˪��W{n�$��o(	�����@s�{�y=�㙛���_�A��)K���H:s؄{�W����i�]<�}����]�P�I��d������2C���d5�����|�͐{�S�(P��x�����':�yZ�o����b�}	�mT�Ch��Y���˸��ٳB^6�}�ՄO��}뿌U �8I��ֻ6�vnrG�r�/�D��͙W����ئ��k�]O��+�=��Ѿ���
��e�'��S��"�z�RX�,g�^��9ݓX�Z-c���nG���cA����m�]�z��7[Ł����ܧi��$.�۶����v�z��>��y�^u̦@z�r(\���}�ۂ8���l�XL�G�]�O vy�u�����k�L���h�%��'O#�3��ۧ��;N����Ξw���6R�w<�v���=�^��k8#��N�.�4dyjƔ�ݍu���ٝ;�v�u�h�Z��]�F\]�F.7��[lR`���u#H�B4<f��}ܲ
?N��]�;�g"�/*��B I�r�����RI��t*���~���Z�<o����R��%	B]��"��v�-�ք79Ox�s�,�S�y��6)�Ӧ����@:�}`Y�o�}c���s��OD,���>']��d�s5|�4���%w՞վ�n�=\E�_��GgJ�(K��	BL���Ÿ��7�qVt����a��&�3��]��w|��=�c�w��p�zOĈ�u@�~��A��y|�z`����%A�>.m�֑�91A��X�h��נ8�+��m؆�6՘�ޤ�T����6��}_e=�BP	��=�a����=k{�s��ϟ@�:�vX$/+�����A���ߔ$~�у��c[Ż^�;lY��������f'������i�?�f$���[5����z<���C}g�7]U�8R��q�.�:��r*#n��~$[}���C=�7�P��R�U+L�ۜ�c@��m$�U��߶�I�{��",^������)��|N��]�A"�=�'�s�e�M�����wc�~�"�ٶRP��m��M��!	:}�v��o�3MZ�����]�Gy��2�4�d7I_�-��H:s���g��L���"�w�$�>�F��+ֽ1�c������!�O��=�sv1ڡy����e��i�p��Q�g��0��m��N����M���B���B���{���&R�!�s����k���RJ��
�"KhWށ��Y<��2zo�A$�o���O���T���8�Ǟ̲BŔ04�(#��`$���d=7�>��7�ҭŴ"%xrC�3�n�a��$$�Ӛ�cs�)����u��@|
.<؆1��LZ�&2�+�Ay�$���C�����!��`�I"�I:vu�r�����s�։�v�?O��݈@Ho�d%��k���7��&���>R�^M�L�M���>Ό�����f�D���j@$>܀0~+oޖ>'�8���9]�M�6�H5T���#���t5qtS�޸��=��uur~~o���"/��J�:�uB	ӝ��I!m��f�.8n���^9z��	$����ѿ��2C	��1���G�8��z]wSُ�'�O�P��[~���^W7����o?h�3%�Sj���Z�B��_�A?Ѝ���wz��-�&�[�$��{#�����
�h��3���b�7}%����E㝰0I]~�H>�U�����{��z��::tx��mp��R�Aٗ����}�n��a���㮸��r0�g]�nY�W|��3g+��Cǎw��<��T�Rt*����'�p߹@s��9W�I�HSڠ'�B���� �_yH��um����1T�%!}5I �;�������3�ܒt�Nv���6��W?�߿��k	i�m�~8s6|�ĕ����?e_y�����[I�G׫��ݱc�;檋I�m%p�i	��o�L+���+/v_�a�����4�R���Ú��H������ꎃ��a6�l���ă���|I ]'���"n�BI]~۲A9W�!>��3Y%�M:iWf��k��Wb IoӬY$6��P��k�JV�}��ć�04
)�(6�Ω|��8�u
�O�/c6/�L��v	$m_����Ԉ>x���wN�|��}���nw"��������.i�e�|!��y%R���?d�e]E�ߔ�ɗT�`��-�)��<RU<z���W?\kn]e%z;r�9�,��+qۦζ9�t�T�n�z;wm�]��m�[��	��nb���̓�7;v�)��q�d3m��kUۍ���|a���%Ԩ񤺷n����ݻkb�m�8��[p]�r�wuEv����Pq�㫜Ӹ�Dq�m�0��;cU������-aY�u��l�܃ڊB|�h�۩��p�r�]��U�b��Kn^�f�����5�p��{rv7]̓h�lç��?~�����TJ
8��wo��	/'�6��BQ�����)^�nl��� ����+��.�i�mӫ[Ǵ�������\����I%��ڡ?s�����B�d�w��Qi �M���ڧ��ܯl�#�'=�K��y�]�{��A��s��z����Q�6A&�0����7��$�S�I&���>'�~[�����ي�9�y�؟h�3Y%��4���jWdD�������,i��ٔH��8~�W���g��*W�����IS��&�T�i�ű����y��y3u��3��y{2z�lh�K���þt��h��>���~=�݁������#�:Q�S�W�� ~ͯl�o��E%I�i�vs��,ﾝ�����8�̞6
���n��X�H,�^z�ݨ�c��A����,�է��:��q��	�t81�]G�<�y�_zA�qf󙠃xҺ}�/:��Y��	�y]�!?-�z��
��vp^���~+�͒�m�m�s��Y�	n� ���nX�yMv	��w+�>@���K��9�T�A��IK;�׾ɇջ����}R���I+7=v	'�3�y��$*�#%{k��'A��0�l�o��?7|��zL7�Y턑\�(B~Y���Ǿ#ׅ��;�����`�ū�b�h���.��d�wHí�z{q�T�][声�%��4���ߑ$�λ�3�p���x�:�.�U�+��,�WaQ&��$��^rd�on]s�c�*R� Vvz���p��v�E=��~~{�)*M3M�=����BP�϶���S`wxqϽ�[�#Վ͊�j�X���-�ʬ�:B���YC�d�f,��BU�<���=��k;}{��-�Y�۰	$�y��0��ZM�-�n�z��)]��G�c���{ޏ�0`���H9���\Y\��z0�n�,X�.s*��A�M���7��	��^ؼf���Lm�kٹ,	��s�	}^���|�ߛ����wا�jB\jf�֊��n���f��{J{7Y���e{\���f�c�����z�{u�L��_��H#o��A'�^����f�����I~��c%� Ӫh%4ԯdD�w�J��On��_s��w��}y�����.��o|HX�-RtE���>${ջ @�P�y!��w��|}{�'}岈x�4R)6�7B��u�r�������������|�����/��,/���imUM�S�fU�xE�y|�U����#�Y�,^�S�l����t���	e�3o.��^LU�����Noy�@^�-a�J���Ǻ�h�� �����������O�����;�H�m�����ߗ׏��o�ߧFH^X�g�.�㫰���wnM��*��v��XlUg=��������cAU3/�����{�.��}��M=)�46{�~;����=(����0�l�c���9hOQ	�]J�l��S�~$�޻���E�_vy�Ď�5�J~���	nf����u���%������U���{� ��݈
����^̠Z$���0������Љ
@���B�y�d���������-Bϲ��x��U�m���W`��ݐI�>ڿ������$k|��S;KJ�[�n�%�W�.���O��d�IE��_fL	+k7��0���Q[�d��MB�-�ث�yi4�,޼���el�ʉ��2w���+�}w[���f�T�@xt^*�0m��"P��vr7|��ݮ0�!�(���T
(!��wBdݷ)�T/n����Pwg:���Dvc�vyV*���g���Sm�Lqne���0�;��c�=6��e�M�d�EV�d�թO�2��zčU�>��]��)�^�v����w����J�3a=�ꊨ�V�6D̂��OMv;4���AI����r�%u��8��+Bȍ��l�Qтb�ʖ�EA{�e�#�\��I0���1jU��u�E.��+�Ic������{���NˈK3dh�\뙑�3�5i�T�s�hnG��WBv�tv����T�V����=W�=D:W��w�m~�Γ� ``�^9��GrGv��5�����@㌻�>��
�x���`ޕ��_�Δ�����"/b��of�'=�)�j��9�H�n�vh�o�]�\ױ�1�V4SM���}C�D���Z;�-ۡ|�K��w��,�WA,�Sz�Z��x��֡�!��kj3����Wd����r睶�j��;���}����6vn��x�v�ct�Yg����My�����l� ����vX��*Ȯ�CxM���K�Q#�g���[�7�n�i?m�`�Aاy���Y�V�Y��r'+}S�=��όf�6�є�b�ll��I����R�5�^�� Gg��W��,ވ�Q:H�\Dc2clU�UK��V´R���$�B
�k��Q��B�PqAE�"L�"V����R.b�EpcAU���\l�fHA��b#�BԥVH� ��b�#) ����e����b�#,�U�Ɉ���V���I$�TLE	d\ĲY�22�+�[db*FBȞR¹TX��"T��H)U&*.+b##@I�# A-�2AH�\Q��U��̊�#[ir#!1�1�	R��"9\���*X��K	d�J�Iq�kq�2HF���$L�b�FȬd���$KB�Z�B�fA\j@r�ʖH�"�D�`�2
HIe+W$X#r�pb�@d�ʕ��0Tb)$�X�$qr[!e	�Bb�eIH1��H���H#��YJ�'��k��j���۹ǝ�1��ܷm�k�;��5���v�ε�n�7�^�n�k��<�S���чm%�ڶ��%�WV�DC��ݍ�.�mvN�4�v�S�;3���onk�<s�;�y�GV���d�w�0p��r; N�#�o��޼�	>AdÚ�趭�n�h�)uBd c#�ݻV������:��ۊ\۷=�뒹��.{������z�����5�]�ݤA�ۃ.B0�r=q�ع�e�����F*�X͠����`��,�2��l�r�Q|�;s�8x����=`w	�[r�dEuI�}G��g��!v�ׄݱ�����F��ݶ�l�>���^����v�.o;�$ދ�%1�GH�9�����E�u�(4\�ۊW����v�on6�}�y�� S��t���v�յ��;�ۍ��re�1���厭؆��ӷ9��<\�u�j�88mۓ��6�r�I%g�삞�����ݮj��wc�l5���͵�k�N�ۻ:��������3��c��%���`�� J�K��O[]�9�,r^��f�	�WazWdѸ�#�N�P���Fǅ�{Q<��2��0/G=�E�n��l�#C����F�;U���'F�n���.�dU=n�lv�q��.+8�.���֖������DR���y�,S�ݔ[=w���󞳤kfqӝc�\.a:��M�n�M�Q�N����c���h�Gn����m͞&��!�^{tі:���c.s̘*�l��\v<�y��{%�t��Nm��ɼ�ga�p��<� HYA��q�v-m�3��뭲N'r��[\=�z�1�� .�;�)x�-q�U��z!�+vxv�ۨl���]�'s������\��8ջ޻����Ju�Gbf�s�7����^�vQ��ٮ�<gm�=��<��Zy��'Q���a�4sNdS'9*�)	����N�G��6���ݷBm�\/eե�3ڞ6i��쳎��!:qH���qЁ�RöqllX;r���vn1�`y�&�7ݜ���Ghnj��;��[s�se�#pg��^����kŐ��HRQѡXU���htWF�<����q� :]2�O\Y�m������Z������qq�Aی�k��녹��8��69u*�s��ݺ�����ޮLvĬ�U�Fͳ�v۷.�p9S1�j���1e瀋��A�βvD��
q����v��'m�t�r��Qu׺ �h�)7M��Vu
�ݷ���M�
}&�A�=��hc���	O>�Ҍ��i)��U3-�;&҅�#���>0�%fw��J��m(��<>�����=~�a�~�u�T
~!��d5��~:o|�?~+�
��}�W`�n�V�+���	W�PG�q�J���
TA-�����X��>:�v��f�ş�$ef�A�W��8��"��=�����HUהD�١A�F�� ��j��h]-
K�l���7��$�%�k�=�N�(���޽N'S�8Jێ�=(�OFK��h�n:�]v�Ezs�y�o��	�A�Eo�����I#3��?	��k����*�����'3����-A��h�n���3޽�ʗ���Z�}j��Ok���QC����u!�=�|ݒw���;=�#;���nj�!��������hH��@{7�k�g=�u�k)�_}d�?g������3���E�Y|�����\*�A1F�I]���N�{b ��eմ}�od�y���%��Jg�)������m�
�~h��iX�C~�$��ݡ	�~��C�շ�'�#1�>87��-%�	�B��jW�~$�u��v}�>�����r��N�n���w�]���zNG���&s��j�n���t�.��h1�{�o]���mֲ$��&���ŷc7n������v�U6X�ڣ�M���v �$�����r�^ܬ� �m�H�}��x�4RUM��"��=����h6�����W%	%��9��IFS�n!(KL�;�sFi���xi��2Z-M�c}W�������v�t!�5��Ǐhe��Ȩ�Ί�N����$_wWt��6��n��/�_y�\f��G��Ygj��zc�đ��?5�z��U2�b�6��o��罘�fɗt��'ޫ�� �	��I���%��=p��:�7�U��W�M�aSo�,���8|a>W���4��* I>w�b�$�w�<�7B5���3Б(���gŻ,ns�i�qsK�b�7	����dwd���9��Ə�����ˡK�R� _k���� �o;�eB���%�ǽO�O��ؿ���*�AT���'9ג�Qc�N[��[����}�Y&��p�|Ȗu���W1�q�J��m��v{o�,�E���3��W�z�З���#���d���8	��-A�Ѧ)6Ӈx�0���k~ė˷�8p�f�M��K8�3�^hU�N0&���vaz-�R4[w�W/��y~�<~p�-�0�,�9�=�mK�L仉���宩�d@�6��{�P��lg��4O��S��<���F�z�Y��oJ�f�	k���?v��IB�9ܝrk���dS�vP�K{/��!�5S�q�GV����	����_��w�J�n��T�˲O�^�� $7��S�6��9���X$�{���I"
eХu��I�@�J���zY?=YܧĒw��Eڷ��fJ*���
�.ٶH
��Ӫb�$�UPuN�	��m�$ߊ.�ya��+w�~'ᵝ���\D���J��m0�
�=�x�toB
��O�{�$��Gt�.!B�;�is6���`Ga�jO\�a��
i�=�� ��3��K��֫�P*�?r� �&�k��_/S�ُM�:=�d����̋^��/݇��X��n<�����KQb����7~�6��<��>2�5F0�|~��c�/|I�]����h�5��H���+m���r�'o;���v3N�7����CCɆ8�m�k�[;%\vck��Q�x�7`ˋs�u͔�gpx�vn��q�r�vkB��<�):�g<7\L��[p���i�R��h�IX��6��Qħ=�ݷs[��\��t��n�<�n��Y������P���,v��]���n|��04m�]�����Xy.݅�͗�Ŋ���\2��t�r��]k��L�pl�/$��������λ���A��n��v�~$�]s�A w�K�wEN��@��8	#ޮʂ�Y�JD�ED��M���P��&���o�Y���H$_/eBA#��dN�F�f�K)�=�՚�J�2�R�]u�D����/�w�d�����~$��d@�wނ®����M�]*���^=^]�^͞XH5*� � ������;��˽Q�ѸH3k=/`,*T�I��W`��l7<��Y���6ME�PA#��������ܡ-5�Z�x���o�C����8�9�b#i�3��۔���y�k�t��t/ �h��i��ͯ�L��,�I �yõx�D_n+רE��Xޔ��H ��M�PM�?tUS߅����ю�u�xo`���-eb3`:�l��.L[�陸��m:�3�5�<)�\3�ϖ[��̶=�i�� �3<]��2O~+�!dW���t(�=9�ܻ�Ε�j�,��a7Hϊ�~���Hn{�$qA랏K'���'3�b{V�i"T)�D�Ћ;�DݯA^�<%�{�,�7;��{+�3�K����f��'�^����M�]*������n��j��a�lM�]���9� w���>b�C��U�U
�I�l�àyqn�=�cu����<��u������#�	c������&S4�h���}�d�Ff��I$�Ӟ:���uT�6��-��\$T�%��h��Vt�o�I���|���P�{��$�q�}�o
��S[̿3T�	�M2����� �s+�B|l8F���n��5B�Z�Û-�-f>�Н��cc%N���7��-=�bC��p�<��7*N�Ò-ڻ��y8�����7����p����_�KJ%*4i��F�߁���/x�U|�}]ޫ�B�(�Na$���=�S�s�3^=���4��\fUL����%�E��O;�]ɢ�n��� �ߜ$�s+� A�~����P��T�	�N�y$�aSqíqt�f��������m��e���:�m�d6���ǉmӣM�YUBl��A���v"	$c��ٙՆ����fm7���'�[��N%�E&Ra�
��g/I���Я,z ���j|I#]��_�*�)����W���A�4�m�ެ�	�y��L�w���Ö=h��~s��H�}뿉�o��3T�	�.iL��'���8W�#��	B[O���'�s=�q�[�:Eҭ� �|���야viߩ����sh�9@���]��O�t3��s���7�����j��kWo1���l�|�W]��30<�7��A���P{�|�4���l�h�����F{���Ftd�7�t��iu>ۿ�'3�s����z�a��&�I���ͷ7lLOŶ�U���L���]�{q�D]h�.>���ک�"T�Q����I.���h'3���w��;=s7{�3: �����n�!WY�SeѦ�,����p�U����{��~ۿ����g�����������Zv\��7n�I2�f�(;g���AÛ�>$�M;C�����	6�v}c+=�>�..���U0�E�g|��(p��^$�{},Ij��~#O��o���t:�Ͼ'귘�,�^�	�M
*b�m�1���$��؏�p����^~�ND�2�,Y>��P@$��� ���v-���+��FȽ��g�Ƌȫ{D�O�n脳2l}sb�)'=��p�X��#.����ܛ�R���׾W��];��V�[T��o��h��r��kr���F�r����.���.+��x�&�vx��q��g:�S�7�Ȉ�[:ޟv���[[�<L0Ku)��9�vC���s ��r�������s��7�zwHs�ہ^����[\���K������b�����ۗv�܆{`���#�ָHMŃ�k@���ۃ�q]�sTea���t��Ye��V�=;fě%ۚ�)�Sp�c�8�9��՝�ߝ���s���������?��P�$���jl۫N��ϖ���Aʾ��'��ES�B��4g�2]�h��Ż��l�	ʾ�����l����fԞ�[�����[�	M�*�����S�Oǽ[�@7{�iu+3C����&�(	$��ys�4L�٪
�����}��<A'o��?{˶�$���X'�����������>&�<.���SE�����JIK~�~��8���BVvt�'2�hB���gG���;_�غx�(C�>���4[\���q��n�����)V;�Zm���M�$YbB�����n�x�0� ����?i�L�E>?o��^��0��
�&;�o�,�����`����[��~�T{���t;���g�7ף�ܛ��辞��ň�9�������g��2����h���?�niN>��PבG����wLsK��I�d�U(&�=.�k��_+����^W�x�|	�������]�
=�	L6'�EUO���%k����Z�Y�i�`�g��I���� ��}��7c��~5�{S�w<)���h�c6w����y<�&�b�{�����/䒟>۰Aʿy@q��N�xq�#B@�b�)i�O- ��B�8#�'�Ƿ������N���_پ.�e�iSmS^;�� D�Wy�d��>�Y�>�IW7yy��O�|�Y̜�U�D$R����d�5���]f�?[~�O��_yB@5�({��[�J��{�~aU$$۪�3��߮�o܄$��:tᇵ�T\�����:�MP'2W���b��+�U��9Ž}POݍ麺�Cݺo:1c��}�`�vWO�������]�K�۰qCs�#�|�lm�g����=$D��^��Êw��o�ވ�1+���+.�u	��.�A�9޷�z��޺ے����������~y��AB�=Zc���z����P�;2J�%C�~��ۣ�L��O�<#;pJ��@��,�����<����zՉ�hHi��M��j��11G�˻��a�f[�'��V5�T�&�U��֟5V�-yP��w���ʾYu�O-���D���ݦ2��ۚ��B��XX�O�m*p1�}�ǗD"p����7�'Y[ed-�k��.���C=yZ�v�G^���!���0���p�>ѳ׵C&V�9ML�=7:�S�{�w��*f���O_1D^�a��5���r�K��"����@�wy�+�����{,}�_�/>��^���5�?u���kS~}=�Qc/�=L�!��6w;��u4J43D�k4�j�gJ&�����!؄i�1f7��EZ.����6e�#%9����_�E˪��7-Z���?r������?MP\jg)�_\մ*��[�;/YUr�Y����Qt"w7�)L�nu��1%�\�c�����3K����E��P��Z��N�Wt���'�����	V$ǎ{N����1��[��s���ifX��;喆gR�Z:b�i+�(Va�����A'�9��V�L�3�3ɪX�[,���dE��ȹ\E$��$Ye-%U!"(��,TQ�c �"��"�A�FRb0aj�+1D� �,f*����Ĉ��B�Dq��2��e���d���
XDQ��U$l) ɋE�YZ��!"�cY ��`�H*H��IJ���,"YUi,�D�"���,U�E Ȫ9���!&$ �&$�!l�Ȱ�J�Kd"L��HH��&8đ`1�!��"�YV�f��FBI&[����IX�F1`H�$r#���5%+F�����[H⥖��+j��&e��"I ��rȕ%,+1b�F֪�"�	�QG$c+�c6���"�-˖6�;�pl�ʮ9�<�ۃpe㤂�5\�"�HIb��0G$��0��a%��\ra$FLG![�d� ��A����J!)m\��#lilJั$�3$�d�cbZ#�?Z����w���r�����	�Ʃ|�*-�J����4���3*2Oo�����(��V�$���Qy����|�??Oz��B�Ä�'�"����8	'�ޭ���p��`�A/޾� �H;~�	��w����y-�]<d����H\ɳ��n˴�&�T/F��b����lʒ!��{;�0�T�MUP{�{��Y ��p o���%"��cb7=v	$�y�OՑ�t��J�j���Y�"�1�rm�����I$�s��?���˚p���]��BQ��v�4
M�������s+��F���H�WV-3$���P��k��g����"�RA$�:5D%��k��ڲ�Jo�\� ��[�	o�|��ut<нs~u1�1Ǟ�r�S{���gm�u��s���5����e���nz�-xs�]v�N�߸ۇ�����߽������դ�0�ҧ�IR�[�Y޸�����ee��R���9�$�z��/��zC��;ݎ4��o�E�-&�)4[��<�a�6����<�9�v�8��x���m��?�~o�7P)?�*��M���݁������g\��:�4���o��ys�4JT�MUPr���9�:����� �ޯmB@$m��$�w��K":��5�q�t��E6�5��$��В|��Za�oω'��[�|�o��'��Ŭ�@��	��7��;������D~$z����s:��އpe�C��Nʾ��
s�PI"�F��qk�Q����Y�݊�������Mʐ��o����b3�v��;W���~�)f�G��D�����Sq�<vϟ�Y�7[��]:>�g���,�����*�Ulq�rg�o#PJ��IP�5����V��ׇ�v�=�=?�}l�}b�Zn��G/�n;�n3wp;iAޜ6��p�z�۴�/Oj�M� p�K�m��C;���y�ܴ]b�3Nu��l��u;v�\p� j�G"�:8�=l��oc�8��r�^5�f��i�N7:�ڑ��t����ܾ-���d7��/oD�q�= n�Ҕ���8�m=��[i�N��:^������a|�hqQ��%��',y�Џvw[q�;vO<��=�=ë��W�R���ԬȏĀv���I��8P�۹��Zں���r��oނ*�ܢ�l��Q�����-�;V8SϦQ�v����\%��2����,VWG�T�I6UT6�B��<�$��ftn/e����_�!$���d|]��M�M@{ظy�����{��쐂	��p������=��HQ#Wd�����̣D��	
j�����?s<�P7P�g��o�~�G�<�����yl���S�+I�߾;���mڭ��`Aױ���j(�7f�#�a�]Fhi~w�%�����am.�$���!�G��p�?7�zBh{��L���kϷ'�����'��յh���d%vjyd��]���n�����q�:u�\t�&��F�]j��p��bRm���<7Z&zer�}�"���hj+;{�ă��p��'{�`��ړ�s%�����`%W�e�`��$�����j�D�,]��>li ��8H$��\�T�QM
j���=~����NTǏ]�M�m�z������	o��Tz�}F�:�lJ�}N�e��M�MO��.�Q�w���gT���X$�� �ya��@���j��}D�1��4��|���T&;t��;1�hMuK�V;��j�A�ׇv�=ut|�����4JM�P�v6�?	��Q$��zB5���*�ff�qe�?�c����D*�L �¶��o��I�x�?
��A����|O�~�u�,���T�7_��c8�eV��l���N� $|H=~�!�e�Nk=e~w�۝�ä�=���ߪ|��(��uIO.{m������mu�9�T�VD'��B���T��Xpw�@$���6��xn
LS%�A$h�^��eo���W�C	���y�I_�����W�k�ȥ����
���hSUT�=}�B	��y���CF����p�_c��_�|��U�	�9�
_\�=�ȟj�EP	��TAm��4V4�v\�pI㭝jÃ�[�vn4�����ϟ�:�B�t׎f-�I���$L�yύ/�*�%^�}q��_���޸��E�(�M]��� ����l���C��|?��L�󄃋r�:�����?{��T) �AQ�����@"o�����f�r	�*�:���$6�d �oz�/��<��D�T�e��u�����z���=/��	?��;�c{�
{sr&��7��de�k*�P�Oاα��,����͹�Q*]�v��4kn���2��(־�BP���^)�v﮻��2A��4�Z<S~p���I�b�,��~�b��9�<��*��{�쏺I����}�p2��LJ��j񍊣T��N�td��Qn�7���]����b{XJ㭍���K���dٞ�U��qω��%�8I'}�b|f[;����꒰@|D��H��1>����[m$�t�=~����n�߻V��В��H��8~>knDq)�מ���.eA&�(SWgrs�~�p�J�������γ���	�ｌO`S����h��ϊ��{�U�c�jq�	lq�I$���|Oč�z,���c���O������r���	K5=����U�F�ܗ_V�$��?{���N�z@r�rkK�3+�MY�]�ɺZz+��r�|�2%I�=��;��&���e�J���f�N�<��d8�&g]	+ ~����+��*�ѕ��ɕ\>�^�`��-��vC���ᰁ3L�7�/ri㇗{q�/m�<r��RLj�0s�ǣ�����c��w�m��F��^6��tӁ�QlǱ��y�������r���]�����\ۈ�"<��;]P�1O�^0�]�ۗ�J�������6�jD�[&�5�9�7&�8[%���-�6��׋�Ѫ�e��:]�%���*��cWA$FOf8�j�qͩm�LV������Cj�n��(&m�-#G�w�� ��{q�#�v��C"a����	�}q�$vn9�?d��h�:#T�ǯ�qioui���x�QW�����TZK/�� قV�vu۵���M���e$�t�;��BM�y�~7W�Y^���?�z�{}�A;~�}qk(�	6�!MK;��-��`�,�i�$�{���	�퐟�_��3:���=U�I���'<�tQ�R
��	�o�ό���mL�@�n������	$��9�{������j��t�B��II���d��[%��{T�Ob�z5[�f����ߝ�?��CD%��c��~>�� �/��|�y�)��R�wzٗ�� ��󀐼��Ӫm�-#F��	0n��ꮝ[�n�	��"�����,���Q`H賎�w~�ă�t��[��&&]��S��3����p����ѵoKv�p՘���w����1����+U��VF=�xH�s�h�
�#T���8	e�������޺�i���N�t��G^y��<|]3E�鴛����Ļ�r�wp��$��8~�z�T9��s6���A>ݺ��A&�)���<�$��[�x��ܵ�l,�^ߜ �H���ŏ�ݞM�0�k|�.b�^&�qP�<[���v�.룚�������[b'f,{0�[�w�aA&U �����B	#���A���޹��db�Fw�ߐ�쐒A��1��uZA�J�~���y�0.��	$���p�@;޷�%级�z������-�۠ڣF��>$;�n|H$�7�~W�TE{7�f��JQ�R�^����¯���1�y�hyfg,���}��ϊ�w8�����!���<��{%�3�����w	o|� ��[eΣEPT�i��t��֭T���q�� ����'�zm�� �� G�m�O��TӪj���f�A��砆��'6[$��S�ujм��֐dh������AS.e�}Q]��Ѻo#��s�hҪPt�N0�N��^���v���j�&
�Ч=�%	B~�B|I����Ʈ�������  ����#�)���IҤ�[~����,�Y)�=��A�����I�_����5�.y�?x{��h@U!+�j{$o��b�?Uq�r�b~��z��{�� �F�{�d����[)�A������D]_���8�1>$�������y��/e!'Y������jUޏK��*g���)��p޽��v��=3��8�)i�kmH�~]}�>����*��O��|�=+s��}��[�D ��CAQY[~�d�w�p�S�nZO���H�:	�g���?y��0��բ�@��R`R	�D:e&�c��s!�ۚ��q��a���Q�[���c����ߚ4u�Xi$2�_� �fo��D��ʼ���U�P�y__�%���ҍ�/)
&�"EJ��w'�$��^��jt�B���Oā���I��p��o*D�΢=ޓg7�<�4�T�Q���zş�"vk	����/�����`$^g�쟉33�Kᕈ�*���5=������'�/ă/ݶ,I���$�����o���a�=o�쐳��H�tڠ�TD/��|H$����㥺����~$�w��W�������f�3��� ��3?큙�fL�033��30����3���f��X�`fg��fa�����fa�������f�f��f�030���`�`fg����3?�3���f�� fa����f���30����fa��������)���x�����0(���1M�� �      �      @ U   � � � 
     @x  {u�
�J"()AT�ۮDQ	u�S6�UF����J�*��R�T@�M�li��*�QJ��X�2Z�mL)���                                        @       Py�UFl���C��u��4==��R��� \�R�w{�U^m��r�����ͨ"�\ �L�@W.�UDP���   �� �2=���  Hre��{���A�� ����` : � ���*�ko�            �A�XCT\�j����^ ��O{ y˾�@^cD�}��4�R�]8  h-I�@q)x�J�BJ�    �_-BD�=Η��T��` f��R14��
�r�A	B�f�u�r�IT��}���Qf��(��R�ۨ���EPv����J�B���b��  �        �AUI��ї�0=�-YA�]� ������ٽ��>�q � �Aۜ3� qʶ�H�_  !�>� �p h� CU�9z�rҀ�� 	�G��z@�oC��a�Jg�%(�H|  �         y�J{\�qiU�Ώ�����]=�^�Z^Ӽ <�+3�yʥ垵���6"�L��:7 ΩGns]�wmG�ӽ�T(22�  ���
9���R�>��������ԩ���c+�JS��-*J�n �
�5*UYa<mR��U�5���
6�4�j�J��@          |>�F,��wmR�Ƚ�K�v1��� � f����Cy�=���:��A���w��@]����t�+������W|>�  7�sj�צ��p ;"]�͗U�����\�P_m{���� ݱJ�d*T2�B�Y�$��'EC�Sɠ))P4�S�i�R�   =4ѕ*Pz@ ت�%%005Oz��*�   	4��e*$� ��?�ɿ�O�G�{�U����f�~�ꛎY����$$ I<�>��I	O!!!��	O�$$ I?�B��BC��y�����N��
~\?��|�[�s����_Sf������Juj�H�:�t��?D8'���OSY�f���دM�a_���XY*�x:'՝�B��O��2hc@i!��,d˗ޏGd�(>TQ}�>tz`Y���u�Vm��9U�F�ʴh�B�a�;J��r����'[ݽȹ)��_b,�yۛ�p��˭ך`ƌ�NƳV�k2�m$�xي)4���<��Εk|��턾���tWr�bdۿ�W�����a����a}4C��T��SKU�磶���{�bJw)��7OcC-��Jr�٦���S�\�ʃ8�n&���p�F�zl��!��3����L�����֞�s�w&��h�>#:�ukE㤎�Wa�|RT݆su�����X
h�v�W!�[S�l�;��8vw8�7X�<m���ծ�,��KI�Zu�Yz.Z�hij�!s{�b�t�Y�i.s�r���t�Q�z�7��go,H:�-5洔�Gc��X��YD�!��'"N�8���C1�����Kwpn42wP�(�(캩tGJO�,�JbG����r�S	e;�C�0'!��K��� d�w8on�q�@�UvZ�eϸP��+�N�,#�����ԧ;Z�Yh`S�p�8��@��S]h�9��AIns�x����s��Z�V�D�,�{k�#���e9��.�ޗs�b��1�ݏT@�W[��.!���f�Uw+қ}�	�(�wQ�W}ֻ؟QfA>&'v�7↨p�Eʭ�.����8�9����Z;P�u�tt8S�hp��mR/]�Ϫq��kN�X�]���$�F9�gn�6m2�-��M����Q�uݒ�� :9���vpn�7����d�����N�f�&�{Gn%�aȎ�{5\wVC����b���Ȍ�<���3`Vh�&�Zۛ
�d�7�^W&w�n;�[���8Zѻ��WDJ���;F��InVn���m�������ޑIT�����f���Tr������T�u�7g�tm�(L�ˈ���i��ຂ�7_n��ө���<��>a9��cx#�Ӳ�d�[+���ړ��х��|R�eB�J���:�l�2���ƩFڮ��J�<U$b�h��
�l���\��kŒ��9��t�f�""]�ŀ�N��[�	h�`Oq�sp�(���Ať��h�TҸm;wm,���O�W�<���Q��h�g�e���dsu���[уw��(��*i���R�Qڴ4=$�;;^v�흩��22n��c sT���Y��<�f�{8�7�#�Sb׊k����FN�],��Հ�Q�י]��i�7' �Zw�q�&�[�q[cJ�^�͛������Zv�� �JZ̷O�����ɽ�i%t6֢�_�f�Mb3rtIw	��]�;5[C�V˦�wJ��V|�������^�m�5���-ֳE��|�l-L���X���'x1���7�'����\�f�rj��8�Xv�c�ؖ�>M��򰀻X���(CU.BŇR<ͿMT�ݖ��M�>���+����Ȼlp�:tn���M���,��Ook��AvU��r�r�]ц1�v��ܑqU'�����;����۸C��L5��Xv����K��ps'�lw}|F=Հ��zĢ�x�ʌ�����%��ܝ�+���n�&n��F�by+��Y�sA'>O�.\n��PxN��Ȏ�pG��{d|���y߬�,��Y����s��T��2#�����V����d��-�Gtsv�^�$���J{B��z���3��0j�򕧱���Ł�$���ᷚ0M[����T;Vr��e�;��W7.q�f�i6����z,�(Ӛ�7zQrQ�[p�ζ;w��vg@{n�(�S"� �&���{�m0���'wq��{�qe+K+��n�`����X��.-|�"ۢ�tDI�]ٻn��\W/�<���⣭S\�h�Q�N�yQ�����呋ǁYD�����s�7�V1Kv#�A$��Yy��yӨMEs
��-�Y�d�՛�
�¦� �L[���C��:xe�w��%�a� v�������j�=��D{J�B�ºs5���[-�1n)���932�r.r�qc鹇�#^ܯm&�O̉e�_�=A���xvO�oC7ko�����.Q�{a=6��J�T�k ��J��d.�{{dd纳`�4�׎��) \7Cc���n
{>��y��i�$�u���ϻ�\Y�t�qӁ�gw0:��|�|�X��J:7�1�AF's�%�M�5�u��p��:)����Fn�g`�jB�ع�w����`�]�Gd.n�Nw."۷9,�q[��q����u�ٍ�v��o7n��ŕ�F� ��Ϋ�K��R��q�k@������c��x�F����ΫDF���"; ����Ѻ�l��Z���A�d��xx�k����� @/��t��[�a���j���y�D��;ja}���׺h�� (��k��Kq�NJ������k���z����X�ǱG��mܹ ՛N�^�h��x�%�ͽ��ǀ�D"�F�)�Q{��u�G��{�6Kٺ���AI�.��A�k�1D������-������iǄ���9��0+Q�@�A�"5�ޮh&�]��(�]�f��W6��� S��g�כ{U�-� S�r�f2���e�`۴�c�y���b	÷�s8Y�Zt`,Z�@��.�7R�eԱ\�b��)+f��V�+P�5��w���;Vs��3�q-F���O��K���*%�m\�i
|M�5F'�P�=�6k'ݎkŹg�yݵ3�.D��'l�l�g����e/9a)�yp�d��b�ue�|�v�w�d�NIǖ��w	��q�`���U���g��=�ڻwV��`��qj�N,��k��a@]�-�s9�6wo+yʐ�۳�,�:�T�t��]3u���8vMjC�_M��tC��B-���y�Z����B�u,�3/NW�w�<�Ǜٸn�+8�;٣Ff�P
9x$�rgE�^�]��2򛷎�ٚ�J�{N.���Oi�{�s�H�T]-Z�4V���лS��omhl��L�r�'��I�{�U9�t�VQ:���˸�WwN�����)���B6D��ol�Y�6��Yo�*�r��a�-�n���	1W	Ԭ氵�t��j����wf��eUi=0�b�M�Ak���Co̪ WITޘ�Ts8����\aS���@�ڳoonn�nV��Xq�4'�:��uL�Z�Z�!ɷx9�;�G�Y�����D��x�9Q�r̓��#4�L���f���x���g<K(�&n$��۪yra����^�5rȲ8.q�f�[0�{��2�ݻ�c�� (*z�2�u���ѫ�s����n��x,���Rš.6t4m�Z���5��9¤�#��u+&�z������t�ޟ�q����:;����Һ�빓�S��ѕ	��$[�t�pո/řsm<�<ou�Ν;�諱�IJ�1�hm3�V��\p��f��B��ka�1�yt=�P�\r����mz*�Ge8a%�C�1���$�޳��m`w�TR�ף�m��yf��=�FnTf��|kЕ�]R�c(�@�!�7Lt�N�4���k�M�\cJh�����8ܗ�m?5E�Ը�Y�y�
d�4�x��DA���2��WFH�[+�o��ˋ�ְs���]V��4cgic]�㨣�߮_��x�6�àn�!�'Y��;5��M���=� �3GsJ�7v��b��-7%�B���n�A���5gZ�V�ܑUbːA&����r�:�[��"�!��vC�~Ek�e�M��SY��@�vᇦ�O�e	��N�>�;^���4�y�����+��2��5�X�)�.�n#�>ٻݹ��U�v�@C�]8z#�)���R�ooO;��Ջ��KU�'j�n`�rX@Ϋ �7E�K���������g+`?iK�A�y���Ү}�j�'syu���jٽK�;�S0m2УM��؊�	g`��3%&��{��-�{f��w;t\�2��Y���!
�A�"�H<(!\Z��Ϲ�v`��BZ��0�"�p�� ��x%�����l�%y��jU9�m��^�#���5n�+�&�o;�Ѻ햢=wh%i�t^��;4�X�՛_���cyW9��`Ǧ)zS����؛`�]��N�95�WC�e��U�R�C���j���@��k��i�j���rf�d�u�Ztlȫ��Tm�%p,k'bb�I�vhve����5��f��B �y�K���s���MN�ߴf��\� �u��ؾ��G:��*CWV7pL,����Ǘ%�&3P�Ņ�6���AA���\�w�}Y׼����t���8,�w�=�e�#pN/���ݫ�n:A�Ѻ]Vm�,�ĆN�}ːo�+;�������j�E>[X����=�<�]�;�^�ݭ�D�[��`����T!;^3D�	f�[E�.�	0lP�N%P˽t��wtc�4��Z0F��oKh��nl�c����v�vn��X�ɪ���X�|ϓy}�XJ��=ٱ��bǞ̻۝�1kcbV����Ѐsgv�;3[�_W/&^�= ��콩���o����v�[�Pؤ���B�n�˜��G��&2^�3S�1�n=��}A�j��cWgb�դ�jYp����q���à����1`���:ީ�N}�]T�	��xnm7q��vu�h�u��ˏ�8��d�`r;��/,ɱ��8f�>�ssnǥ$4Y��@��ДZ�ooM@a�lI{�߮���ѫ�`�u���ܲ�c��	�Os��յS�U�[u��t�Sph��ZU4���نҰ�����n]�2�|& �L5\Z<���F.E���7�V֋��\.�JZ��0����}ͼ`�[g~���F���A�r5�[�l�	�K�-ws�es�)���4�5P�����tI�E��6�z��G��D=��k/���1��¬�M��[;Zv���a��gQc��ZK�ǩ��wQ�J�f�xGr�4��F�Э���vPr���M͏RDW�7�[��!'x=⾉H4 ��8���7�Gs0�$2���sT����
4��٠��H��zA���IL�y?ۥ����'TI���T�ڮAƴ:�ɯ���˗H��]O�����r|:�!�]����p8ob�d��s[HQ�ͺ4�fq�=��1�v�=�^X;��:bŶ�m��qñ��0L]չ`��A�h�o8�w>����V0�*��@�#���a)�ݛpK��M�GS�7������U� x ߵ��<Y;O��X1vҥB� �k�v[�'e� -�>�5�u�*�
֬<���&�k����3������{R�h<�&�-�=���u]�7�3��u�1��I�I9��!%Cwնi/`q�{#Gl�8niD[�s޲c�g*����^�Ҟwf���l�H<#hݶ�+x�&6��s���w*��VE3��ӄ`�c%�cЎv�z"L�s���0J�94�����2Yh�,"�h%̪���˕�i��(�M_�:��0�8:��7oR�6�	���3�'�>��{�=��w�f���d����zK�lC�5��EU��ԭ�.̅�\�׋��!�ז4��B�8�����s�ӻ�Kk��:`x;�Z�ѽ�gJ�؟v�tIj	�;6�ѽ	�v:�S5j���!;E2�:�m�zW9�m�wIü���2�'#��N�roT�q�Yk(��̕�{S�z#��&����|�o;��g#K�rTpgI��kD}��6]]N�&ӗ@����\�8�\{��Djo��c��.|�6;�뱝$˸Ĩo%��)�9��S��ԯq�J�r/va8��o3�-+��C�鹢����l��@�(윙A�b�2���Êuc}����������n�/;f���m�[�_{�C�����/���&��_�y{Y���rM����<5�&�3z�S����9tB��z��$t �K����ؓѱ��b�-cA���Ի]w ���|���7yM�nܳ�2�)^�Pf���3OIpN4X^�*�Uk��V82��v
���װ�oo#�'	��=��{�:v��>y��7P��Q����s���%�y�}� �x#��9���F����e��GZ�X�J�8F6��:���.�P��9�B 	�~����/bWxq��NjԹ��z�R�wYE�'�)Je[�j�D�1a��-=I8�D�r<`��3��o�J�c9p��\�ڥ�N,[��>�B<Q��d1 �fl0�59�q6:T�V�K�;TT�T�6����ܐ�\�`I���/(6�m�V�jVJFWB�KDt����R���7\���7�1����z�RAN�QT4%��pіdG����\F��X&��c�n[����\}�La��w�;5^m���2�fmc�8I��n���3�������;�8N�wj}:5ז�Ŝ�Q���>�$N-/8Y�B�:���w8�e�˯q�r���1�@� �Y'�$ *"���@�IR	RVH ���	Y	$�	 �$�$$�� �I����H��* 
�R�$RH�HII	%`(B!$�H�$�"�E����!*$
�(B@��!XJ��a��a I (B)  � d$�H
I$�����H�BAd �E�@%I
�H� �HT$!R���)$�B
��HAa%H�H
I P���IXHIRJ�X��H( (��@��I@�(E ���!!
�@RXY �Aa A`+ �$�		������W��-��Կ��(����̓{��
�%��r5V�Y��\��������˽����&(Ҭt�9��)����PpW�ŅH�t�������y����W�2�����Nt��!���
�U �E����{�ۥG�fe���d��� h��p�ڍ��E�,e��%�ݓ&i��S��Դ	i�kmT�4��V�,�ײ�����pݭ�÷ �����v�,��4=/3���-�v��o&�E�۳�	�+Z�ڥ�H*�;j'�j��;!�{���{�jK�mm�v��YZ��ƪY�.�v�cX���G���u�;'l���p�0�L�z�46�]ù\����]�{�]a�9� #Y����ۜ��K[fD��̸������|O���݌�jcHp!���瞋��e6�m� ��h����V\��3�p�]��{V��1,jݞ�"g6����8�nH�dµg�59"�J�	���?D�5.�!�a�{%����ݧ;��f�2ڒ<���P�0��3%f���*�,n�8�f�xxF�a��Zt�Q9pA�-��c<��\�(X�IZ�,�e˸h���nn����G����p�i>]��Az�ˊq$j��N���r2��v����#ð���0�V��'[�u��փ�9]�-S�3�9x-r�2�i�2�Nf�	P�Vs~5{�j�`�sV�n^ZZ�ގc(�&OE�L�N����m�/{z:�������f�	^d�&p�r�V��,�|唩e\#U�UK�{Q�׷1k;u��*�R�g��o��2�d�-�6G���sIg��ұ ��a��{���O���
U�+������qv�ʌ$��/=���fb1a�y��p����M�y
s@���S� �-OG?mxtN&J���7&T�7F��aɯ��+��!7�f�|������=���Ǳ���t���u����b2�6�v^�b:�w�s�8��e}�9�)ɡ�s�pE||*�r�&��E��H�3Gy�ʡ����WT5W5*��ON��ͼ�^{B݆�i� ���Y�_R՗��ǌ���J��2���Q�؟����;��MYӏp��@c��w`�Uy{�3"L����Te�hi�9�F��q����]4R@����ZP�����M7Bj
E]3PrI�f.ʽ��w�Wd�i�%�|�L�O�,+ۏuU*��1��=��-BwT��Or_FO%{��<�IA��~�Ү_#�X�a<K�f-���)c<Xo��3�{}�&�Sj�.[E��n�u��2rS^^�;;Ên��i^+�N�.Ey2<&���%�|7���v�LPs@�+ŵ���ߨcG�L0��W:x&z�I78�Z!�B>C�ݫͣ�)ٳat���;�ʁ��,���"v�YsqT� j�U�Xa/.�M�X�w��1f��	4Y{؞oq��q�@qL֑���aL7�}Y�7���*k|�=�Y�^>�����+��O��ݶ�[k�h�"�!�c�[ʮ��O2��nբ�̴��4�x|��_��Z�$����#FC�o��|*󩗤{�,i����s��<q���ބ�1n��77��gjr���3y��Ax�a;[`�nn���R��w�O3��bOV���c�V���PdY���{���8w6��^�}��c:-�tŅ!�BU�;I�;t�ACyq���{���nh��Pw�kw�9u�ك����av���N$vi/�M�h���1'����A5#Zkm�Jy��L�Hk=�,A��.G�+�u��T��ͅ���sA��0M��9�ޗ^�My�6��V߼.%9Ⰵ�|��짛��͗%m�}�e<�NcP>W��ǀ�I	2�,������$��o�W%���g��/�tw(�G�c�N���9q��Rx��x�#�b�o�y���V9(t�����;�l~�%�0@��^�RZn��Љ/�Dr�;{/�Vf���*j���7ub�f����f���Ӥ�y{n�������x���h�JJoFh��Ԯ�0�m��1Āt窨�����2ph݁���!�sB�N��n�d������÷z��H`�
��cQj�����
��6�(`���T�sI��oS�0�����X�8�$o+7@����ж܇~�ز�nBu�5�c���j����3�9Xvh��"/H6��O]u�̜�\�@���/��LJK��
��zx\t<\�,Z�8��ۅ���ڕA3Ќ���T����@�B�&:;���'��׎�x���đ�}� 5�,�VS��'j�\��TJ��V0y�XN���;�El<��w�e	���F�U�[�V���f�X���Ξ�;'���;W��ON��x�U�h�<�5�XCR��{,f���h�P�!�o{S���k�xN�>孃;;6��@؛~�*%&�%���3+N��Y�WL��^�U#O���w��Y��ے��
$x�����OW��2q(��J^��{ Ů��T��j\�mi�gf�/�����l�;��8zJR��:Ƽ$k�+!��Y��!�V{�P���k��h9���z[�}��� ��-'��C��o�J@]x��dN�aΒ�^*�pu��	�	��3���¦k���s�wĦ2�Ċ}�U�vWv�"Ge"2	%���{�'l5����Z�.�T�x�FB�Lc�W��vv	ݞ#=8�%�uu�[FP��u����
�!̜�','}�B�k���F��k*�<A����/&�^�x�� A?!�4r@�U�݋��������:��T.)�/�(aA��t������G8����9(��R��ǎ��o���Z}��HEm�����@�%^ޖ^���B��㝝��$m��=�wi�=V�2�X&��&�ۗ����q��(�"�sa��8�F`����Ö���-f
;R�W�Pǿuq�:�5�����5C.B	��٤�z{����U�����{e��U��Q��s֬Q���C�gR��Z����<Ӿ�痀�|t��̞G����J�٩�1ʃ�ö���"��cY2��[�l詭-UT��j��:г`f�*o�J�xz�Q�II�x���r� �پ4�-9���vWm�m�0�Fc����$ו��2 �*3��/y����#9�.��ky�0B<(A�L�ޗ7N�4�oaׯF��9O+ޜ#I{7�щªGe�V���i�̱\��]J�;�I�ٛ��w%��JL��9��	��cwx�7�g.gׄ�8Pz�k����R�	v@�n�S�m���:/��2/j�A ڑ�{a܅�{��ieE5��6�d(����)�7M������)<wqA�յ���/�s����[��&H#�\ܠ�V�_�����x���]��AL�GS��g(�m��)o��V�|��qw�����𩉥Y������rI�4o\��್%i����U��ŝؑ�Ǣqx����n(q<�{�� ���xN�{��@���D��O��s��=���<��1� }��6��x�~�x[В �	Γz,�\�{��7���5P�P�L���Z5{��w�XA�I����k:��s8M�F(ލb�{�Ƕ��M�m&�$9L����_o�dAKʼSinr�y{��hf��J�z�5*��3��f��"����d4�:D؛[rv�e��a��7{%�}q��d�JI=s}D`�������'�Uiƶ�.�����%>8�=;B���'�&��T
�z�ਰ�ča�HG��\8������,!��b!�Jp����50Յ��aVk�ԯh�k[ˣ�н�� �ߧ��[�:��,��{"��q��3ޡ�Qx<��k�ʎp�l��VE(U�����E	�^G���'�6~=�I�x]|}�4�-x����y�\1�m��_���I����o=�vx��<�f�@����b��+}6����8�5��֢^h޹�	�Iv���V�����Se���q0����|/{�ʆ���w=�ɚu�Uzң��;�quc�Y�/�N8�a����m��st:GD����Ι-�΋��J��ɓ-�ޘ�G�R��{q�W^]9��i�r�A�mA�>��m^�n����٩��8��
�9��uEx^��Wӫ�EVQǗ)���1�S���wH<)FcM���^��,]n���҂ p8*�C�^�
��Xٺ;��E�V����$����|}s@[*�s��K��f��d�/�]�F��s�j���9�]y��m	cd�:�u^�HwƹGv�)�n"[=��uV�U�̜�\�on�^�f ��O��%n�f,��]����:��e��1� �F����!��^������Ps+z`y�x�ݸ��2�>y"�y���L�=.�I�;"�{yu�v��u~1fن0��ͮ�P�䷓�r���qy��e�5YϤ��-E���ٕD���@�O�[�m����4���m���Gm����t��-{���؜����|��{�WpQ�>VV�1�J���c��p���6�=i�ghw-���~:��:����᳑�sn����&g��ݬi��3p�/�r[���Q�Red��ҫ �`,z���J��Oy<tT��5�/t��4�ٻziY��Ca0�V��TF���rd�0TѾ�jԌN�<&�=�.4D�Xd�m&��}��=8���d��8f΃�O��Ǆr�+c�;пz�����$͑<h��ƷZ��O�5�o�n�,wXsVn�����Ŋ�a�|��p��P)���q�X�C�qG�OZ�41PJ�ZjE\�r CrMFrI"� ��8��\* E���T0�S�Լ3�zH�k��h�I�M��bB��*�����JC}��@�;R�L����ݗ�$��G�$���ܨ��n-��L�R��^f��Z��i��T��4�*�崤�@�KFZ�� ���i�F��ǪѾ^�D$W]���h�����vn��`f��ۓ���.d��*��ۋ�t�ˉ�jy Q��'���4��v-��|�����sG�"E�������C@�gn�[*�l�q=��7�G������7�<�w3X�:K�g5O��l��G1���l^z��O�=/G���b7JT�=Y,93õc���яC�7�8B�Z�0a��m�܇�SP�R���hC�W�&����F�<�	�cH�h^�\�>�_v7� ���<-�����"��!�v�����G�g�4�H�)�[5d�y�N���66�f�\���+%�޷�m/�\��^�Ëӵo�i)"�L>���s�yM�3�3q`ǎk�j����d��V
W�W�\�{�0GS7KדK���@>����7�.�sU������:�Gj���n-n��Q�9L��0�ŝ��z���������=��>��1���X'x�u��N������Vf@�Ⱥ8OL��K��9�\�Y@è�wv���.@(X�rT��tt�r�������Ҽ�W��l�G}�Ty־�sȞ��r��H��	f�����Q�`"2��e���-��6ۆ�!ӫ$>{ܖ���(�>���:���Xy�{J�?p�O_N�<�:%��LË�������V]�5ǸbXY}�)��{������0�|�[3H���oOP�1zg%6��{�r�}���z!��:b<hB�ُ����P�[��-RU��܄r��q�4�q��d����,��+=r���tS��t�*��]-���^�p`J+˚i�;!�â�x���/��*�
�`u���dM�)�.A�q���k�/����P���B���5����V�%l��N�����9���5z�^aつ@[f#/:��ܼ��γ��ެ&����ۡ�j����:�hu�6�x=�beL�
r2[��z�sx���a���E�va4�$մr����w\Q�DS���9��^�{B��Tw�;�o�4t�pO��>ht7�2��3n��έ��f@�<W�Sg�c�??�2����/nρ}�N�����bD-,�p�?g^9g���y������0A"�8vF	
]ڷ�$:�t\"i�P
����<����/#�K���(��
����>g: |z����uu`���B&��)��fТ�{0�=�0�3N�^T���ׅ��v�f+�lQd�A���p��"�ni~[�I6{��c;�{ּ���{w-�DىCw��.���3�Nr�ÌQ<�&���#6'c��]������P M� 
`���z=�iԮ�y�ڇq%�`d	F΢R�30�n��U/���7od��>ܑ�^�|�L�YR���㦬f,{a�Q��O8	8�84s2Աi�a���ƛ�Qn���&��LyOb�*s��9P��Db��^Ð�pR���*������Y�s�#��$�X�9b��Slʬv��A;�^Y��G@m�L���I]ph�k�^�)�HG`��TN�a�)J�@�}�a�6bf&t?\ط�ȗ-ηyA��*��N����xso�P�B��6%�����wr�c�>*mW���.����s��~(�"�Y��)�ހ�ds!�d���&�)zv�\{����e�Nxs9"V�����������AZd�����՜�+^X�������US
Ї�ȅ15�X�o65'��}&�M6RNm�v,)9� ��B��_��4���F]�{{J�#�BEs1=���tr&�8\�'�q�+�z!��`��s鍂�u�	!!I�$�K����c�<q�𥝝G����̹��Z��J�I�t8���]���d�\�幛vk/Κ��;Lj�	���{g[L��:Ŕ{f�P2h�ǈҙ.��Q�X���q�����gs�Dc��vz2�Q��ۀ�<��k�)�����Ƿ��s�.��H��5��Y���֝�����ap,�:��-��{v��[��np=����Ca�V�a{�T�6��e���׵�ۭn��=E�x�،=n�%	g��<8է�-#�حc���	�9�p�ɷ�Ms\��-@M��B����ظ:�9���9�l9;Z�i-�m��(wl���Mep���|#��۶�R#G�>���#K��P^����V�!:��9�x�f�8��\��_P�@�i�p�6ݘ�9�XBx�0/k;:<-Ӷ:�f��M�Ԝ��X��玒n����=�3��Ok;lKd��nܜ\��D�l�V�s��l�6�q�IGGg��&&o8��!K/.�=�f�{1̛q�9�ÃRIɵ���q��	�cg�q�� �[����<�n����=�9�u��n6�m�n5Κ%��s��v�8�Gk<�]��A��.�ḃ�G+��Nb�e�Ӂ�^�8�l��z�u��G��5�¶�O6녰�
���7cV=��N���>_l�uה�w)�w��l���5�;f{[�ɮ1����xL���tV7��WM�.`���!wg\�ێ.,�L]��M�q=,a8j��U"J�֝����gq����hnv�wu�����n��rsȧ�9�g��N�m�v��
�; ���;=�� �a�N1��2c*�7
���pezls�jz1���m�3rv��i�'��]n�ne��-�d�l���C�p�Ɍ=���j��1r97��P�uB�h�]������u�4k�l�v�F�sj���7/�񹛳���e���{;.���wb���pmwb���VϓX΂y�݃��[��F���r�l��u�ȑ��v9�5�q/n5�wl8v���ܞ����\/OXN��u���^u��r��p+ն��y�N|�\=i���0v�S�Y}x�y�':E뱏I+���	=��s���8���'��mq�m��ۋ���N]ϳ�*f�X[&���<Y��6)�V��tór���{v��E����w\�� �*��qq3�^N��6��p��X֎����3ɬqG���J[4��ec]��j��u�[sہ�kۏn���tq�7\�v����.��5s���G��ڻ-�sp���+��Խ�5s�K���C=�ț�!n�7n�2u�u�U�kl��֡�,k�ř����P���m���"v6�t���=ۉ���<�������9ݚi�-ĉ��#)�� �����e\ƹ�Xgp��x�mV���^j�m��=
��v�P�ώNG]��i�z����
�u�ros�z�7k�ݪ��2��u�X�|]���N��{qy�:zw<s��x��A��;qͱ��[5ێ=�p��sۖ��L+�����c�ܖӸ��:Χ��c�ѽ��8�c.�F�Y�r	����Z�:x��֨t���2۩�9���[�We�we�����I��X�snۋqѳ����Ͷ����;�k�Nw%K����5����ۺ|W�\=z.���[u�ByM�N�k�(��t�M�v�ǒ�@�$+��#d��:v�a����Й�ڤ̖��ŭ��=>K\n6v�j|��@�v��q]�\]ѹy6�ۣ�.v�\�vzϧP���=����㞶�
9�yi�JX��㜽M՞�΂0�q�}�n{pni8-�[&�	�4����1�m��a�6��nL���6�g�$�8v �t�;�KK�Yݍ�ٍ���e����U��iN�Yr������mv:�%vzV��d�i��{��ؓn�Í��wn�n�n�)<�u�n���5s������9A��r�d�ݹ�M���v�cZw{���nx�r�X���=�ͺ�.�����#���y��nG��׵�Y�X��%Ѡz�������9�%�\���Ɏ�7&�9��L\�f�Z�Wh*rX���
^/A���X�}n�Z��ּc��0�z';�M
��7Db���1�%qڭɵ�C���t]<��v=X�][��8�v7z�\�#��vc��ݺċ<v���rsw.�q��w5K$���\t�Ծ���2�$�:\�{�T��Ι�<�&�v�5ˮt(냭����z�:���)�\��c=�nw�6=��i��p����<�r��q�g�V�ܔ���U��ۗ�8����7�g\vz睰u���5�ٲu��v;r�ޝ��n3����c6���.�tv�9-�/sXzÍ��tN��nq�x�(l��v�d�>�N=�ێ��&�	x����]�I���l5g`��C\񺥱t9�&Ş�N��]��%خ��w���I�;��������2�[=��	��P�ӷ����ׯW���{n�[Nz�{
n�Y�xpr�q�b�xqoAk`�9ֈ2��x��O ni.<�ez���<���k�k�l�s��\����X�r�O�wS�8q�[���z��݉�z��j9z$z���!�'�>��y/ ���]i�:}I咹N�`�<j�v;��3�ԁ�]�vL��sO;M�u�5���!|��6�E�թ�W���[o��K���(���)��2�1�7Q��& �ur�6�v�ѷ��8����;n܇hx�ؗ7B�����5C�fPT����w.N*s�H�Ƹ���;{�ka7g�:�ڀ��,b������Eۍ���t�m�,َ%���\$������^\����R�#ۯ`�&h��x��y�v݋���+[v5���$�3t��J�T^�j����NG���=�f���R�۬�2K��;m[5���_m��k�hJ3v�@-�9��8m��i��F2�Dcq�K��k�l�󜶳"훛�+m�[�$f�n
Ɪ3X�u�Y1�7`��])q��u�^�;r�[e�%���v��MM��sֈ�.�v��Kn{E�7Kœ	��J�M�Kgg]y� ��c�cIvĚ�����;�ZKr��k]n4F���lZ�ܠ��H���'s��^n5�Gj�9�,�T��vwk\9�����tm=�����[[�fwd$k�A�:�ڨ��4Qvծ"S�󥓝�u��|O]���S�9�ֶ8wZ��%^��Oj���=m��i��\��F;�v���ʍ�vG%�m�Zc���:����3Ż%�n�l<j���lv�SWɮ��m�u`Gֶ�bbޭq.ݎ;lE���Ɍ�6mt��n�cP^�&�݌�u�Ün.+���
:�f�AV��OSt�ֱ`�ݺ�/d�[��^�BTc,�[K��
l\[9ʪ[���Ⱦ=�S���vJ8S#�{Kv,nc�ۥ�9Jz��]vvs�kgk�\v�*K��X����ٸ�6r�;�uå��gn���!.�S��8��c��q�tv�c�v��9��-���n�9`�6��&ٗ���o�9���ʭ'o6�q��G���U��؃���у���˱�q��|=��X��۳!�oM9�Ɲ�t�o�{���glv��d�dmڋ'-/m�/r��rk�;�iذrɹ�m��7:E�{nn�j}�
B����,a0���n׌�Ѳ R�r�9�3+Rs����X�1�Nٰ��$l�2[���s�u��Ν���%+�0lbs$�զ�B�v@%�LQ�3fV9�G�z�"��9ի�"����⽇�i���C�9Z���62q�Z��nr�i.��x�+�[��κ8����u��1B��u��j*l�Sgő���`�%��l���t�C�m�v6D��ͤ뭛�vՀ�nzƳc�c:G�Nݞ�@���6�����p�w8^tqТ���`b�ܭ84:�׵q�����\lhr�;jڹvٷ
��4��\]\�:���n���չ��gcx��k��Fp��o/9�=�z�ee�r��d�2�-�@����:	��6�qٹ+Ɨ��I5�k��;�plර�grf�Xݹ�᧋���۷�u�����.=g�oY�m�x�\�:�����#�v�L�WY��-�3��>yǎ�m�ls��pD m�\�kv5�j�ng�z�k#��g���;q�V�΄��\�g7f�6�rgn�yc��5λ�)ρt�����t�<U/s�kűT�Y��u��n��v7t�k���؉I�p�sl��=h��Vڭ��nL���`�q��\��Ǌ�ǳt����3�:�#�������۫F$���mH�b�v��°����(�v���ݶ��[�����v�<��v9��ܢ9e���'I�ka����b���miwg�m�bVs��a���[�u�ho]o �Kw�[q�r�i�N�;s�
����/P��Lf�Řb���,g=��v�@�f���r���z���ٮ���A7Gn�@.�N�aC7/��S��[u��}�q��<榭�^+���n��,�k�\�x�s��<Sy7n��.�c�Dviљp�bH�eI����p��t�c���ey.0n�ӄ�������q����^K����K��1lŮ:�b��r]��<�F�Y���ێd��F��d�8�]Ɔ�='cF9��=� ����"4[n4۱&k�õn;r	]�������2y"�.�D�z�;<lk�g���9#n.�g-�
�)ɍQ�Gb�ݤ�h�}����і^'����f��t��I���=���^}n�͹�䖍���خ��r۩u51�۬�M�����n���+m��x�dn��s��Ꜣ�=�	���p-�#�f.*��H��Ѯ���Yݮ]7�z�B��5��y.�McODLBS�_���m�m��8�p�-��5���0���mJ��E���Q1Q��إj���AaiKQ,�J�UT��Q-m�j(�lQ�¸AF��8��Ŗ�ZU���KaV�Jօ���8�ڠ�1�+TkclR������80�D���+iZ�FՊZ4���Kmh�T��h6�aKR��[R���m�jEZ�B���JҪ�����+KQm��(����Y[[TZ�ڔ�V��J-�I[J����Rԥ���6Z)m�����1��R�Qj�R��
V�h���ZQ�X"�*�Z�kJ�EF�l6�qK���Qʭ��J�ղ�a&1EҩJX��0�\(UjV5J�pb֔eIF���e���h�,�R�TYm�B�e[V5h�-�A+J�Z�Dk
6���"�V�m��5
��B�[U+B�Q*��Tm��jT)kk�R�m�Q���KmJT�p4DT��ʶ�J��S	\�)AjT(Җ##)j%km�-ZZ�[T���V!V�j��E`�J�*°��(�a�(��ҥ��UE*(Ĺ$�:|�xy��<��=�Cݬ7�ζ�gyF���jp/�3;��Յ��]��h�m��[�'"��Ύ��Lln{I��,��E�s����{Uݷ�x9����������E�Q����m�;�$^v6wf��n�G6d{O�W�a7=[�M1�2��ᧃ��N���Wd�v�r[������=.�c��ksC\�����ܾMچ�8�Q�I�F�m�c��Gg۸ힸ�����i�j�E�v��q�pk�Όpۮm���m�GR�f�J��w\Z3i�s��n���@= �v伸&ֲ�]f��.8�[f��W3���j{)��g�8����ۉ�ݶ���K�ݑnͰ3�zd�N݉���U��<�3���<C"����Η�ޮ9�u�$�':�L�s3�/+ۗd��>|��C��:8�g#wat����/�l�v�]p���X�0vx�U퇰n�t7k$���.*��۝>0��FH�N;�㑵:��t:K��<̶\!�Z��w�n3����:�ՐzZ�ȇy빺��'����	���vΤ���*�P�q�6Cv��Ӓ��bxݫ�Ɨ�۞�G��L�j]��	��q���o<�"�:��a�q	�\��	��7o�ۯ��6�wGC�PXNYWn�����ώ�f��[�7g��xy��q�Y�n^�ݪ�|2i�ɻql�m�U�N^�]���Nˑ����k��탸�<<{m�r��'6�q4�:-۪�G�s�:[�����*�&K�Hv�����밠�.�x�y�	�=���93�t��ղqs���d���]�m=�v�'���S��5�s�]<=Y:��m�sBt8�睁٘ �v�\؋iQ�ۓ�[l�5�Lgv�=�)�y�����ە���n��gN8�ٵ�\��q�Ҝ��]�|c�=�'7�Z��g��3�m��q,�7̥ָ��n#�;lk-ݰE��ˮ�uN��w��y�2v2v�x+����ʪv6O��{���aS��Svwq�M�y���c����s�;yx{9��ێ\(r'���*�n=�{a�QDxܛ�L���DK���%��Zc	mZ�8�8�q��{8��r�{n�¹y�Gy�=��;c����|�����ʩ�ە�W�66y�a�q��Ap��mɄܣ�{�96Np��Eg����Q��0p����	s*|�$�Gn��@�s�sh:E�yN�eݐ �t�L&u�PE
>�UR�Cb�z� ݭ���s2�2ݫ" �l"�����;gǘ��}�;&�괆g�9�ʄ�0*�E�mM����|�Ӣ=tv⬵U�Oݹ����ܓI#�ySI ��d(-��1
]?��w}�=�F\��>���[�>$e�M�Aowm�ۙgop�D��s�+�(��UE@��)ݶ�`��w���i����- <�M��x��wwk��T����\ͩ��k����;j��C���-�ͻU��l�kZ/IW�sn��i���tG�	2����{�y� ]���4�#{�[�)�j�O{�B��l������������ઠ�g��˪���i�n)Ǉ*R�Fż�L��Q�w�jA�KN��\�F�7V�m�K:���Y7�b��}0��E�Ȧ�.d!��&��,x��y��� ����!���ݶ�/��]�l�6�2.�ܔ�F�@��m�i�i0 /��ڰ 6�Uy[y�W�(�~h �ݷXu��_�uf7�����4���H�g4�����ۻ  �ˠ�k1��۝���ԀJ%�~`U�ߦ�T��J��\�����/�"7r���e�E��������CA���E��f�עk��I�߯�ߘ��n8���a��[q]�.f�x��8�N�/����kY�p���_���ѫ��Z�t�?z;�v�k� ��ܺ��gR���^(�m���>3;��XN���
�Pe��N��	��.�Ӌ�ܛ��gX�fwsv 3r�7�+V�ю4b��&�S�u(�2�4\T��$�eКI/$^ƈέ�RH����F��PfL$��GZ����L����;���]�`A�)���phW��})�,��6:Z$�*�Vv�]r�L��;7�ݑ �˦�)����(Q�J�B��&9�dm5V�]�ѝa�@|w��X |we�E�fz���s�lܢ{׬��˵a�oџUAEI6�Gy��>���^9C�����n7�I�#�2��D��nےI�k�)�	�0��tlSUג��m��	P�}��ӹ�f��ۧ]ks%��tEl� b;cU�߿����T��J��ny�wn/�>A�o� gf:i�����7~�}��`H��B��Z�E�A��iTPZgm��#oi�������7^�n/�Gn�z!���0����4�M]�����D�qB�T�����D��K� 3��L0t�q�nK��Wd�興����L���d��.<�ԉZ�����	�Fs��5�^�`+��r� ���S~WW�o�e��o���md�����4�F�AtJ���瞹���P."�l0�l��g?n9�y�x��w~X6y����r��I3g�I'U�MDe�%��a�5H�筯������³sb�P���� ��r�Dww]�[�W��/�󔷷����<}q��n�x�C�c�M��C�3L:#Xs��{#m����߾lD7w���>~`�fy�gwu����"7���>yM�|d�9��|g��M!@pTTR�껱h�A[͢���7Y˹Լ� 
�s�� ���q&E�r��9���,�K�h�0[-)��]+n�4�D�ou_� �%�2*�T���e�lF ��1� ����)K-2S�S-TV�E��Yaf��������A-� �7v�Y
k�}u�4�o\��G�𪦪&��;�� >��y��^�m��5���YW�� F�w;�" �ۦ���J-�i��7��B�	T��*�v&�N�,3DO�gUuQ�mE�H�B�EӬr�G��0h�C�QD�=ו ƽ��ju�������i4������{s�,����p{\���E��w5۳z���g"��"��.���B��p�ힽ���vS����n������;[k�y����bM���2�?׭�GͶ��7��xٹx �y{.)�*G1-���^D��:��:�q�<�b�A�nƭ���=c��G���֮ݨ��{�ܚ��L'R��{KJ][n.']lm�5���\��=<�7��Y��N8�4��$"�M���~ ��>L6��Q����@�s��� >�t�'BӅ7I�n{^_�~�����j�vPoџU!���D�s�&�Id�CQ8�.���]8�{��v��n���2�0��lqt�"�Oud�Bl%�QH�{͸���~b��y�U�V7<s��"��dF�]4ý,\�-��J���ۧ" U�P�6M�{��Հ #;.�H�g����M�����D�fݫ'Y�QQIE���v]M��Y�Mvz�	��U�y%3>�O� ���d$�?m�@�lc�IG�پ}﷿L|��Җ76�f�G�d�֪N�v�JVr��)�+]�]�u���~��㩭50{��ͻ�@|ۖל@�Ә�׵��?l�Mj�����q oeס�3���(Q�J�B��D����B�(��ep6b�Z�4��w�Y�(�9�~��#����_�y���r*ހ���MIݗ����؝:�!X>h���+���N�� 	��_~� x��y�#I������3�QD�M��m�� �??�ge�vy������@ -�z"!����w�(�m0TEE����cٚ�����@/�35� 3���vwu�م;Uڍ�H���^��협b��B����r��6��� ������IS٦2����78�H$��cs�����g�*�7I;�n�Ģf;�����]�����:N��뵽&+�<h�+v��De�+�&�)�)��	J�y�! �1��D@��w������ef����ݵ�d$�=��֏�$��s��h���g0��vå� f�71#����p�6cި�z�g/:��B��UB6�<<o��A{���E�"�ȹ9�
q�Yϯ|��LY>]���8���]�A�Է�P�h��$��'�vI�����ݰ�<���̮!$��g(W�w~�͜nb���wgF��*�QD�^a���Bݯz���6� ;�w��7;���H$uM�D���
��&�}���ȃ>���TP	�U�I��c�쮷>����q�nZ �� �lM�P�WBo���@��m��G�^�Ŭ^M#ƕ��-�ݳ�p��;]���=3\p՚p�i�0[--���]u�	v�u]����g�d�_�h�
�]�O ��w`�cN
��*%9a'�Z�|�T�a4���j�{���@�{��"gײ�d�j�Z�mu�ThK������6ۇ&�Z��Z%z�� ���66Hw~Ɉ߀;;���IS{ji�@%2E��@�yGYm��Y.o��Ș�?O9	�	$�����y���k{j�� ��7��0`��_NZ�7V�5RR5��xfd@��X�v�l����(Q<zȺST`�\����0���'�U����,�"*�EQ��q�ڦ t˚kr7�v��܌ހ��۲m#�w#� ����-k�2���:\L(�#��=�ˏ�p������ֆ�(�*m��S�u�<:A�(p�^�A��ۂQ�����U�����3�+��r�[�κD��y}�~�I8��+Ԑ�u�a!�@��o��� v���ūeiW��n�� ��nK�a|e�_� ��r��X��o���_%a=�pT�AQ(����$��_S�e�� q>s3��N����;y� ��nKd _N[���U}�!�89��3���0�j��RW�.b��'���E%e��N<�>Iѽ�&��v0!�!T�U�P`�{���U��Z�Y6�����%�̨&�K˳�����3�1#��2F,�<�E6��5�����|��X�>�J�s})�br�nE��8��C��nQWY��rgE�n�!�wo�ȣ�=��I�+��	"b:�Xq2��neh�ۜ��-��g������͵���=p��igp�uݤ앻cZ�a�í�s���q׵�nEag�;,=z�W;�o[�n���W8�I���<�n�6�.=�o�zή�n��N��pT����q�u�h}��m�����Нdj�SS�q�Z�8L�4�7��>�nΊ۩�g	Oa�ZYԯ'S4m���ò��Ϟg�k��qSv�C��:d�0�h��s	�Ql&�l�;�r����g����vK�<:��+��Ӿ��ԅ� mc���s0�5墷���`{�7=UVs�T���倀���� ���ճ��NOF۪�����a��R5��Q��u
$���ă��'��NL�'Ď�̡@���!
�v��C0-U B���$^ł7�rk���ݽ�@�3&�G ꈪ��2�nsċ�M��Ai�N�zu
'ۓs��݈���qLT׉�j����{7��I̛bk�C��_?7Ǉ�̻\��]vz�r㵛7g�<o'-�mvz�r6�̹����~~���[q`�����	 �wuQ ��M��̓
"�T�s#	7��^��°�$&�4�iP��s̊��*ČԺ��I�J���;w�Eũ��)��6���B%w��#�d���j]�M��G��ܫ�osUs��Z���>���A>9�nI���+g��<�v�E�!�����wM�͛�>$��W�r+��L珯{��^'2m�=�$�& ,6R���դ��v;�H1��TI$�>$+{2�w���}��>.窅!ZL�q�fe��B��$��m��>�ueY�φ�:��ė��2ފ|H$V�eW9.�^F�=;�8f,��m\��]�sֻ��pN�^�pf�9qӴ8��լq7�P:_��e�|vu
�ɹPCgͭ��$h%���}� �>V�"p��2Bi�BK��W��ܹ��])���T(�n͹$��̪j�7��{��nM�'h�&�	�6!�'�ʟ}�|s;2E�sP+#aQ\+��TwܸA���l�W�&hwu^C5!M�go#�H�vR��֛kH$�����t�4�/���?KwZ=�ڈP��z�%��:B�[�����"^ш	�e�, ��o�p�����Nk{��[M����K��|��ɚ�*$=��)#�;�Ӌ=F����N;z������1�FOd�3]MGR�ݔl�*n]�t�F�kq����BU#�b|C�>��qIL^��1/L�4�۾{�5����,f5!��N���yq��#�+T��/7�����ɨn�Yvb��cjk+�������F��l���%���_�o�~�\��e��{]*4�}�茈@�]Za��r�[�2�Z���yY�F��R��M��a�g7U�g(=�mܾ�V{�2����8/�L����lW�n���N���.���Y��Ʈ���uZU���Rs=��Y������r�e��F��M}[�n�����9�;�J�f+�ȬIoiꭦ������Nw{�<��g��s�ӓ
sVrڒ���s��SlҜ��޽ۗ��8����dt*�	U�b�ͼW���L�����1>���4��5v�h[11[��Hp�*n�J����=g�1�R�n�w"vNl����w��m�X"�a5����[�,�(T"�;U�ǇtT�$"��S|��k�l�� �]�����"��f��	��W}�8���qY��ȴ�5��Պ|�4�l+ؽ��l�X���݃�7|`��|�K���8}�X�,2�Õ�I����_�}����lm���V�(
)D�kcj���L5ҍIR�TD���T�-���
ڔkJYb��+QZ���,0�%�BѩKF���i`�"�+Qilim��J4,���QE�d��)ҕ��Q�c�F11cm�#D�%�DQm(����F�J!Z��E��Ш����0!�����(�DX�5��1jX���B�VQEeJ[U���m\cJ*�[eb���j��B�0�)i,bֵ�hŭA��X��Lb�%j+\`�Աm�*������1lQ��eb���U���Ʋ���aX\R��eb�-�iڕ��(�-�R)D���R�U�)�b[+R�-�m�!m�P��TPU+�AER[b"�ԅE�ѴX����X��хcZ�
�+j�X6�`�*���Z�J�0�X���H��cmE�0b��"��Z�Klm��ŕ��`�[�6���kb։m�
���1������PQ+Bڈ�T��Uil
6��\*�څh��[jJ$KkiH�Ҋo�}�S��w �vd�>��im�!C$���x��7�g5�3(ׁz�$�O�;2��A���y�Mf�z`� 5\�H$tA�I�L@0Xl� kݺ�	���+�k��o�Z�1$�yٔ(㹽�	ʜ��/�yvG�naqZ���;=h�qnή�Oi�*p��Z��n�͹���(�߿{t�b��kxr�C$gnd�'Ăw7���;�����nbH#/s*����:�
I��=�z�-����O\�Y=�'/s*��n�W�:��.�\NĂbx�ġ�K��2�R�{B�O���Mx����Q͒{�z(�o;2��㻽�(��ND�CP�4�O0'������$�;7��	9�o���K�X����5-�A�4�)7���d{f�S�.;��ܴ�ٝ��rc��S^8�c\�Uyd��j]�N��%Y�O�T<��&;r�!� �����޺�H#6�g�u���J�&�ω��ݑD�˷&�ml+jk��z��+ؑ۷T��I��N��s�6����YM���#��e(���Ӻ�&���\9��P$����>'�2�ψ�Т��ۓl=TI �wuQP�z@b��j�vu�l|�olݚ�:�0( ���}��7g�9���>�K�Ԉ�!BM�˓�禉#r�d����:��rc�5�I7{�Q'2��19hjP�%�pB�El�p�Y���b/�&2f�$�ݹ �[ٓ��M��	bZA
/:�D��@�!�[e4'��yR�I��ɯ݇N&���[�THvչ�H��ʠB�PT���8�c�ٌ��s��\➕;�>3��~Ҥ��?1C#��?��
��?]�޽�ޓ��H���(V�]f*�Un�c�+u���/���?��z ٱ�o;6������������9�x���է;û[96���ލ�򽍺ꎌ�]��͓�z�n�g�,��z`��s`�z��B)��tw;�t=urG�c�N�X�9�s�70u:�{o���w�~`��wγqØ�qѱ�<9'�|i[k4옭��z�l�P$�ˊ�&12�ZDT\�6�y��ݦw�������F'g�t���(���s�1�q��G=�6�c��z������\�����8姶[l}���޺|�j܂IݙTJ�#=/K�~�]R(A�rN�9IÈb�e)�>ܯi':ˌ�Tn�pQٵlI5��TI;��+9J}���B�����"�U�[X$�|s��hIۢP�|%�ʾ���A̫rH$WveP'*&�h���m���{��2�߹F�$�d�A>ٙB�'�{���N��#A&�m��}�rP�%�q�R�ܪ �M��N����h�b�`�N����*�'�{��&x�sax��F%m��1�r�·���-�C���I��س�h!{m��|PZ	m�-��Dd��gfM	��{�c�0��t�P�� �j�2��2.�&!�UQ�޺��AP �Ij�Dk���B�eM�:&D^�H�6�����W<ױ���Kw@���h�h����l�Y���V��[�;���{{2��|w7�E�7���m.wy1;��S�	�L@"a����0�{�����˪��u��{�����w7�h*&��N8%�U@��t�8\�W#��~���O{��� 	\W"�1����4H�}�+n&Bh���M9��s�(�W>��5�z3	̚٢|I����H7�l`�����(�����]m�)��ԃlV윳��q�-ʷ��lq^�3Ą4�i6��YéC$�4+�'r�T �>�� *�=�B=�v��ڤ[@����/�"��f!����Ē�F�IE������ �y��@�M�[��ՈRJ��5 ��7tN^ 	�ln��y� ��;��2�Y�n9�VF��)- ��V]�������gEl������sw��A�ٜ�����K�,y���"��3�d��C��rDw�a��m����^'ֲ�$�b2�C��!�3�ν��؄��2$�x�_e
���$�v����+�V�:	3y�T��8&a�Mx��r'�����T�}7�3}TI8���F�^U3��(��ł
q�ˈd"�AgJy�ʘ#����:ఴ(\�
�.�.��%�������~.p��1�����N�^Pj`��zc�eP �1m�O�M<a�A���ns�����$o�;�M�m���>$��ו@�r,Ө)aun���n�}�%@��*�I��2H7�y4@6@aG���a�u�@z\�>U��s�q��D�1��%�M2��,B$�۩d�{:�H=���m�fԸq���g'��#����� L�5��=cT����<�ƈ�8z���f��:ى ƺ��]���)�]��9�na?���p�ʶ�I��
4`0ё״(���g�ꈞwK5�<A��ʢI=��=bdh�2i�B��@a��V��dݭ�vSF�/�kcs�n���;\��v3z%�.
���.
"�,�Q���|{s2Eww���0���t:cTnǦ��*�$]Å��!��p[�'��M���Ӑ��Q�d�ٹ�@�۽�(Tvy8�ΗH��61�p+S��g���ڢ�+�bJ�:b\I$��̡^$��mQ�}�%@��*�O�t���˶V5
߁&�&�$�Ov�������Ŭj��r)�7�(�;���(�U�![D�
���`�	8kn|���D���}3��Ngv�	e����xKS&�M�g[�BŪ�-`�BoA8���5�b���1.,L_b09-�R��3�L�ӧ]fJ%;��NTj2X�� <ݘ+�
�	�D����v�nnx�����w9�6�az�P���7=��=�5�*v�."�v�n�#7r�
z���rm+pݶ�Gn�n{y���|]g��p�=�<���ջ��/�y���N�;$u�;+���նwd9aZT�`���vg�Mu�����W����r��;��=E<�e�C�[��d�v^��*ڮ�&�,�I�s墭ۜ��3�]rv��E#t���7+�v�pk�/IW<7��wС�F��/�*�$���G���eFZ�t����.�>��A3�j�����
n�*V��lK!)�=�r8H��T')e�'*�b��1EoY	��&\�V��� зW�=TI;Kn} R1��ȰI���	>Q��"�-M��`6&�D��"n\�[�Nf�UA3�֤����tt�__�����p���@EPMT�	7�jDo:�h���6�FM�z���I$���Q����;�s��ib����~K57���y9kG�Wk1ce3�nW���>8�{(P�?^-���0�1���b7���H3��H$���6"G��3��T	>���$��#&8h�"l�������H��G����n�)��:CY�g���su��#Y�J�����M�9���,]���3~W-ҽ�̝�F�6U�����Ӫ��������w}G��L�m�$�����R�훞;Ҍ��ٚ�E
���hZj��.�#���P�rJ��s�{��k��eo\O��뮹�8[	�d��1���koe
U8�eUd�T��A�I=�ۮ%�v�#�Z �>US	�ȭKS`���W�.������bC5&ۍq�V�"���/+n�x�{w�k$:;�?�#~����j������9�������6�u�v�_+Ї�\��{���� ZD�gM?^OT��|{w�k�;3	�4Ị]��N�e�ҭ	�#*��o]Q4R���[����/3:H��yu^${w�}F-��^�$�׾$t�0�)O��r�|{���|}8���gjn�"g�s�y�;
5͚w�M��(�W���x^����".�M�4���q���������ݙK/-��z�v���Y���ָ���_������e�H$f_e
� ���@QB���4��MW���ꔯ�X�� ]�r(�3{��Ă7.�"&'I���(V�8]	�d��9=�z�DGm��tt��Z�JQ���N^oUH;��T�ܻrw�\�I�Q�F�A�����a%�A�b%�{(�h-�k�֤V�&���������s*	��3���A��ڣ�Ir����ё&$t�^��'ă}��_���QA��DB�>��#)���0���}s�H$gwmQ�r��'b0vs���-�מ/*��B �H�
��u`�H#6�}$�gk��R�.�x�ow��Iܻr	2�Æ�!��R#3��N��A��FvuP Ֆ䃷}u�0D��љ[eһ#�h�����o�q�f%��{#�N/62�=��^�ocN�<螺�%NǙ���c!ѷ�uo~� O�n��>B����BQ�j�
~���{r$�$H'#f�*�$����]�ȵZ���L�Ҥ�뮋���ٹ���zϜ�6�w-\u�8�����OfW �Ye5Uz��h���q��>$��� �F��׺&K�P����'/{=�J5���'�ME#�&�%7�޶�1�����pj�fh�FVےN���x�q:��=*�c&��|_���QA��DBGd��� �_\׈ ���]��Sˌ�o"b�Y'��ω�=w�TK��,!a�"PKz�H펈����gB��I�'ۗ�T	 ���y#����o����� ���a��C��F�eP$wv�q�]��]�\��$9�A����4�w{Zm%x��xL�R*�\O[R`����!mm��{4	��&��!壻hѩ�̦�X��~���	�Ax��C�)�%'46����{ �L���1�v�xYkXH޻}L�Ǜ�7xy� �=�g�*W7��e�t���ʁq�7���n���t䙬Wv@��?<�Yc_��/Qx��&��h��C�=�DO�:�{Ƭ�ZF�C6�G77S��*g7)
q䐀f29Y��Ұ-ͽ�n�k�uk��Z="�)���l�k�d=Qx�e+��p����T]��RtEmA�G��%�34i��=�A��������hWI����G_�-�=�UvB�7�Y~쾐�:x������I�+:�D�h�NΣlɽ���GegsL�ͩ�keoz]�_*��8��>7޽���Ê��8[�l�>��	թ,~�gC"�O4���T�������QYڨZ�_.�_mi�h����Z��+���<���릯2�⏪;o�1wc���q�sط��bim��ɶp��cG;��%�S��-�n���=LS��˻� �~��B�F�v�"Ff�`�շ}ٌǄ(/b�js�5�[�z�_T�pp��8 �r��(�;���������P[��n4G!��k;��9�v�Y�Y���*�R�l۸��T�S�-]�+	��`�=ΈӸ���Z���^'�+7Z�˴��J�M��
��^�ȫ�Rh w~Ma��ה�'q��ee*¡p��L"ρ�
/�ҪEcYU�EZ�"���PEDh�7h"

��b�lQFb�qK�T*�ڔB�B���b%F�YEH�
����U���[p�Q��)�Ra��mB���&-E1B��	�",���TAkEeb���*
EEaTb�L2���� [b�Qb" �5h�DaR��*�F �D��%A�T�Ej-��E���E���imÁd�1-U(�J�0�V�TŔ(�j��
[(�T��*�����*�TXUaR6�XE)[QJ6Ջ*

�m(ʌ*�VҲ-��f�+EU����%�U(ƶ�JՈ��J����#k�*%�(6��*Ԩ� �E���Q�*��*L5U3���F�qj��-H�b"�)Z�k)J���-�E��PD��V�5�Fж�ЩU+*��ej(**V�T+*T*VT���b"�*�2�EAe-�*�b,����Z%T+-e�dF��ԂZ���h���UUX��E���b�.!TUb����hұQ�Y�ZZ�-�E��Җ,8�8L3��CL��O���p�q���[���+n��4gq�wGd��I��l=Vy�kv��s�猇j⵶�\��tr�U�y�u��8��h��nx.Ō�n�4�u���î��k1#:��:����؛���=X�5n� �3��'k��ηgˋ����.�k���.�����W���PdI�����9�zxc{oY�v�򝺼�;��x� ��mvs�v�9̤n\]��c�b^ü�^��贕#^�Ȫ]>���X0���n�ˋRu�wZ!�N��6գx��r�0w���y��u�;i��{v�V��3�2Q���GV݀�86G�uX��/#ϳ'�eι�\r����y&Ӹ�`��J����OH[���I����mn�c��@6+nչ7qڒ�m���<.i��=	s��S����;�C�qGLk��]�ʜ�8m���2��U�K]�Z�:�^�<t-���,/j�nb]��ճ<&�ܜ����w�M�ĉO@ܻ�湃ל]�t���W�.s�\n=�z��:�����ݨ�;=-���br$��wc�k��g������r�!�MN�Vq�'E�݃9nи\f�#��c���B���pc�s���̸��V6���-�g۴�۰��q�x��Wk��z�ݻv���]��/'H{^�M����g{7%s�5�=��Z{Q7n������bK�ڜ���O#�`ƎϦ�h;�1��X#y5c�U���G�X�[��դ���cv\�ޮ�u6��&�^�m�7i�b�Y����z��˱Wkx��v��Ɏ�kF�9�������eU�۳;�.\;���ꇕ��.�<\�Z֍g��㮮�7S�l�}C�HK�jX�t��]�ε�g�6��W.�v�/n&����c��k�vC]��7��=sv�r��-��Ƚ���b����n�{n����c�z�,ks�4Ls���j�bP�t'W<�$|7��={3<��b�v��z ��ԗ�����{��㟋��I�a�n��َ8LZ�:8��Y7&f�\/!ur��\tz�S��·�ѓ<6.k�� ����G|�g� ]pn���]�C�)�7>�ZK��n��4�-�⒨wv]�lq�y���@'�B{;nGv�n�#���5���>ʘ�1�wX�m4>�klj�e�c�DC��]. 亱�v��]��#�lnc\�\�S��,�I�FقL��ZHr�D89�jvk[���n��-�5nk��J~��{���ҥKgx�9�$��{sD�ww���H�(��Ù���k)�����[h�&�l0S!�=�z����_fi�Țt>&���$��@����W�KM��zK���az0
�3�0�y��D�7)��i˯H쾺�H��ڣ��|M��q
���,H����r(�;;��|v��ٚ��Vq�_EP���� �&���	��[C�g)ʧds��};T	'�3{hW�9YlWe��~|���~c(tli�d*�g�.x�:&v3�v�c�q{b8������I��?>��������͔�Gv�W� �wl������������]T	�>9��^�+7�q	@�ٟ��J�yY|g8N�����"uw%;/�5�-�A��v б9�ۺ٬�j�%=d"��
8�����9$�&��^��k^���^!��ȸ'�o�����o=��S�s�h�{�w�A+�>���Y��<��� Ҵf���Ð{��xQ�>mmȓ�T��Ӹҭ��X	���P$ee� �za�С��MtMm=��T*Z��d�����|H$ն����F��7��:8�zuz�DfD��1"!	#q��}y�s^<)TOE\�Wh�Χ �u�H�캠ofų��9Ӣ ��Ky
7l\7]cs�]n^�u��9����C�{y������x�%@�Z�*���Q�[nA>$u�]P!nI<�z�j0o/�$�m��d8m�fe��V#;r�ė��p����D�I��s�|H�캠IZ�&�};�Q�9� �Ht�š��wdI'Ƿr�H$ F�l���E>P�KTf�ӣ��V3w�s�׎�HIV�8����9���*C��F����v7Qw����v�ެ�1��{���~�5�r�ߤu��Tj.	Z�����;�{6U�t�t�#&`�7w��>����@#7{`�����`�A��r	r3��|� ��o$X"�rf9�mz�& ؞*�}�N� '�v7%���&R��DA���h�
����79+��%s<��س�#*��������v��Ug:�H&���W�$gom��O�U��L����]W��魳�	.`���z�P�d��wD]=�>'č�˪��s���ݗ��f��L�'�\L6���h�vnUx�A���I��ሻ2&bdJٗ�e�\�>$��E�.5�
���!N�nw�)����k�l׉�;���ĂA��qhk˛�ܺ����ڋ���t)i����ΚN���ʻJ�����r�囿jv	��r��}z�JC���	�w�ު�y�H�����d�8"a8-C��9���۟M�+1N����券��O���Р@$�e��YQf��{�|�����o�H|���M�9���8n�#ێX�qɥ�*U3V�5qP#�&�%>[-�i 2�~�< x[7��O�2~�|�^ol�h��H"R���^�m���ޒ1�3�S���3w��F���^1�q�z�q#��m�H�ApY%U��'�櫹�O�Aʖ�
�ا��`�/;��M�]��
��
��i������nV2�&{��W�#z.АHۮ���e��oC�@����D!tA��LD�C���A#��$(]R�n9Ȍ�@��T�$�,�$�]�@�#�g___���G�.v'��js�;�&�mB��U�f�ܼlEܩ�۱��l#�bp��(ސz���ћm5t�^<������F���z��%�/� ϟA?'I��{A��qڸ덺^5u���^+ag�ӵB�ɍϴ�6c�*��a4���f���Yvv��/�p=^�]�u���'���r�c�W`+�O[�(�cl�0��lx�%]�6��{��<���vg�m���Og{l��1ۘ��R�ƛ/.�z�]$y��tzҚ�����u���Q��+][Vm=8�E$v���u9�z�
�غ5��\ݹk�s`AdP.�[���h+ی�����!��P���Т �,� �F�vP%�,�		oOz�wc-J�S�V����I�]-�DD��_N_�Y�+2��$�z2П6벅�F�6"�sMsw�Z#v�����"�V���I��ɢI7/*b�po�u\K��$���R$��eW�Mj��P ��J��Q�����,55"$��̪� 㝽�i)�ot��	qܤ�TYV��؀�i���geW�#{�k�x���� �YW�D����U���ͦ9�Ω�@��<�M�[Q��b�v��ۢ����yM������t����7n�D�A�0���m^�I���b�����ɾ�lIGM�T��ι�(
v�Z�(-0�P��=TM��4����4��uUa/��3��[5(F�M���v�\6��!F:�r�y��K�
^~�>�~����1<f�D\	�I�r~���x���|O�W�^$�o�T4E]٭Y�b�h1���P�P*�+n�ĂA���� ���ط�ҫ��N]^UI9��T�8��Jn"!	 �[AIʮ�B'u�K�ښ�A��٠I f�Z�TS���)B�͡�8e�ApY%H+z���'ue��8�F�m]�7~�8HQY�Do7���62�ɼ�8(��#󨽀�x�a��������-jЍ�n&sݍ�	N���:S�^�W\���:y�؀�i��z/o��$�����R:˺Y9�Ϊ�ݽ�D!�A��LD���aVȂS.���p�SE�9��H�w�j�>'62АM\.�ʱ5�����>�; �n��1|��2�C
��u܆�H,��������<d�ʁR�gF�{�����,�d����.jb�l�;8�&Ro�I��;�lQ����>��e�C���,βn)��4�[ؿTS4�`sc�|q�ā �����R
B��?w�2�H6��C�y���FK�40���&
 ,�{�}�,���h��q�돠x̌� ���}�4��V0�)�����
MT�N��{�l�㫮�\}�=�~�d���YS����7h�_���xy�.0�X�a�c\�0�R-߷�ri �z/����<�����}�{�6��*eO����0�2T*J��w�ri ��Wt;��s�&N�G?�(*e2i����¦���Z+��x���s�y��x<&m��?�����O./�����*c�w��H,�2��1��hg����@������m`kӫ����� ��{�@�� �	@��;���@�B�i4�l@h4�tI<��{�i�
�Y��y�����1�i�s�d��y�2z�hT��aX^s���a��T���=߽ɴ�ɱ����D^���8��k�A���=�Y !l��Ș�0"F��`�����ZAH[@�7�2i �c���~��;���� �AM��=��0�4�P�J����6�q�a����y�./��q��,4§;�w!�{߶�$�B�VV�>�a�MFT
%@���捰7��H[O{�� v��}��9�_8�hBݧ	���L�i���8�Ty�)��Ͳja��������r�a=��3����bVl�M�Ν����?�?�!Z��y�s:,�4pq����4�;�sy4� VVJ��S���Hs��=��c=�}�����<�u$��*{���M�led�������y�n&�=�߾���p������m��0�L�a}^	8'��=lٵ�5�{jcggD�����ߛ��gv��1q����5�;�s0�CAih��{�[
B�`V�
����4�` ��nk�}�	>dT�����ިT�~������)���u-�R���1�m��
��� i&��\����{[C�f���LmH����>D ���~�&��R����2����S�}���A:�g�� �C�20�i��A�ʠ@���ܛM�
�YY*s��2lI�*J�|Q�ܦJ����4vr���
��I%O~߿d�&�Y(2�Xʟs��I�6�q�to�+q��`m���@T֙�]A��䇁 �{����`T��w��4�h*|��{��ʧ36>c[�q�� ��G��|�B�d��3�$AN���!�H)������g��ֺ�����1��e �jck�6���jB�{�{́��)
�=�{�a��Ed#Q�Br�g��O�M��G�x5��jj���+����L�w�z�p�mAq4�أ����l]8��>}K�ݘ[���U�Ʉ�i���J�t�Mï=U���Ѯ�����g74ܘ�쾧�7]�a�Qe6�u�����k�����8��uŷn:�ּ4���6S��1n9��]������0Ý�\�ӸE{��${S&D����\k��uv�uӰ�0��6����F:۵��f����W����t�`�A��P����ݘ�"����Ŋ)#c.�;��5v��u��r��
�<�Aш����nW��z���^������i?$���6�Y�J��S��d�$�AaF�=�{�a��T�ƾ����(&9���l��� ��s��6�@�8Oz�E��y���Q�1�sy>$�����ut5�y�[)
���/;��@m6�R�V�{�a ��%C��m�׻߻��H,7�ﯵ-����1�m ��{�C��%ea�c�ri�2Q� �s�9�c�y��|��X�;���f���h����s:Bi���M��J�Ex�=߶F�]�~��~�������<�}� i��,V}���0�C
��T�N����l���s�掗���㝜d���YS�{�lM�S;�}��1��Ѵ�Øƹ��|H)h���Mn���\�����}��сR�ֻ���K
ʝ�{�a�*%B�w���|,|&����W��ZTd4R���T	�x��)��]��M��Y.��b��wPG�g��P�a��xI���">�k� QhVJ2����ܚg���Ĩv_�Bπ�Q�eG�%T��~H]�y 6n�m!Z!�<����<�L^����c@�m'|���i��}���R~F��\�*S�
��aW:��nR�ZD۾9Ҡшغ�A�e�hg�k0r�.�X^ z���mOո��^�?*������4<=��{�����Ns��'�B�J���9�>�P�*J!P?{��d�Ad�+&ﹸzy�w��اq�w$�@���;��-����.0�X�a�c��0�Դ������5����`T������k��c��=�c\��@�P+����0�PВ�s���a��aMw|_e�/�X"+�υ��"!�� ?��؝�:��e&`�d�+w�a����J�~�}�F�`Ԃ�s��@�y�}|����_�)�{��t0*o��\�_<<<��c�rPI�~��6�Y�����9�w�Hw�k=ǿo�c�V0�,�~sZ�haRX�ID����6�Y6��YS�w��@�ǚ������w��>�mZy��Y쮗Ǉ6�����{qn�q�MX��z�ԠW���v??{a�����0:���!�ą�����{ϲi ������4�
]y��۞\�|���1�<f��o��
ACBw��|/��-삹��e0نb�$��§;�w!���Q
�����/�|�}�0ޱ���g��2�Q*>��}�l��Z�����@�7H6���;Gc�ﾌ�_Vτ���X��J���S�i���[�M���YFJ��S��d�M�aX$;�{|�ls��������76�'�����3Ac�Օ{�8�����ݹ|��%���q��y���x}uK	o��_{�1�lː��c�4�璼�o���s;��P�[������*P���=��X�e���$�ތk7�\�fp���0^;5�^ٓ]�yJg��pir�1ua�Z��-}�=�&�e3rY�����ڱm>�f�y��<'��)�{^'���*������5q���Y���sb}���9��-�<���>^��B���25�H�<��#&OCA��:B�܅X	�o���=����ɤ����v�LG���sң͎����B:�cZ
ݲ��׳����a��H��y,��"���c^$��_xHJ����]OF���^�fEk��b��g����ޫ�3����c�b�aʹ7,ض�-̘�X��F�N�4OR�B����w{#8��V�Y�6��i���K�����s��+=g���̏z�l"pz:���$���}݌�D�{�gP���ڧ�� ��t�cu-Դ��3C�1�R���Z�؁K�w�W�Y{B���"������gK�>���o��f�N��
����T~wVfwXTH����3��4��]��v��m�[|����<�R��+��,��ɏb������&A�WK��a�qY�]f`u%d#ԻO>�Kیr���2%Q�w0^�6h���Z�\9�5���&=���q����d��iIB���gE��0o��EO�:Mӝ'5��E^��PKQ��li��U��~]�gY���i�Wm�Q`�kT�j(��*�E+ҢŃhQ�1Dm���)Uim��,UX#Z�VT�"���թ*U0�W��R���b�T�h�ʕE�֠��QF���E��(�Q�aU�.`��T��TU*��H��QV��������",PV,b�**(-�\W�F�ؠ�QTUPR)��QC�֩(�J�TA�UQF���m+�
�1��R�FT*�5���	Z���(�	l�5��0�(�	m��.UX0X"��Uh���A��TF)mQDAU���XXRQT�J$TZ6"(����j8��`�Y�c����QF�ŶSQŕ�Kj��QUTQ*��5���b�UUkQb[J�ڂ���j�DQ��aƲ��Q&-ŵ�QX�hԔ�#bT�����1+U�Z��X�W��P��PdDAT�L5�+���HI?}��0�¤�'����d�ʐR
{���I�6���=��p�y��0�R��C� �IN�f��y;�x ��$�Mo&�HV�
�Kϻ�h��
�Xs�k���]��<����C�IP�}�7̛a��}�/��
��>	�Cl6¦<�~�lCi(�H,>�5�M�~b�{�y�/_b��T{��&���R
w��2����v����@�D��U:8^�~��H7N勚�p��Th��;����1��� �Y��c�>t4�l��i| �>#Ϸ�dY T��S��y�bM�D� ��>�_W�
>�eT��/����t���ȚNw�}�i�q���T���2M�6�q�to>R�qG�F�ks{���B�H^�]�\=�1�t����ܚH)�`T�����n*e�u��x�@���b�?P��4��#�<	��\��qˆ��b�%��T�u��6��Q
�YXw���5�%eH(kG��9����X�i�w��H;)
�9�k���L��`��$%�
 Y }�"���}�5��gvp������DM��i�+
+�wj$��I�^}"Ͻ¬��C��#"��}T$]eU]�3�������������7��-�i�C��À���ܽ#hd�ݹ1f)��S�/\G�.��5���I$���������w��&�m�3�se����b����ǜ�z� ��H6��<��R���M�o����L���@m6 T�a��f3C%H(�~�&�n0�.�{�s�T3FWMO� -�&�l$S8=zN�=n^�u���d� 8椏Go%=�������߾����a���Ly���؆�X�d��>���43,���@���4��O�3��FF7vG��}5� �<������G�"��B��e��m* A F��"�� G���G���Ȝ�N3�)�{�rlm
$��>�7���0�(�Ibw��ܛH,�Y<�3�^Ou�k3��;5#�� Q�Ѩ���`lk^s܆������u�H�C��E |!�ZY� ��ow�=N�( VX���0�d�T�
!�w�rm ����ͼ��c>CE�*�$�Q�Dw�_H��E�20
I�
�YXv�߲j3,�� �}���M$��
Z{�w��zg]���6o���%!Z!�s|�<t��H�ZA2Ye���G]Ȣ4ed�>���@�<�{��LzJ���n����%�(�w~��l�R%eOy��$�&�>2g�F�J�"%}5����mڋk�X�3��&�n
��T̷�cD��M)	١;���dF��ol־];�,�b�K����x z4 y0�q�L�u�l(Q4��ˊ��4pwX�(hIn�OnS��3�^N7ֻl���n�5��	y�;=��E�dE,�m�W��Nĵ����\����y��P�Ս�]ҕ�[�p���ۊ^8�\/l�vv�6Q����c���v4{P�Z�:]c=7�<�+��g�A�m����϶�vܸ��Y�jn�W(��=k�D�qu��x�xM����%�#۵��y[i���p����w���>1����ۏ>�<H�P=���Ml�+X ����4�h���c+�m«��Quσ>��$(��D9��ܛa���5��[�K�ơ�Tǜ�����B�y�������a��w'Y�JʁR�{��ܚH,� ���y�77H4���7[I?}�ϲ|��ۂ��6�)��T �(�?�zE��O�����9���6�hQ%aF���y�D�21�Uw�>�#Ȁ��#6��&�&�+%T���2�6��CcQ	��phY�
>��@�ς���Il73��	 D�l����60+X9���I��+*}�>��{�u�Cu��� AD@���G�>/�R���e�	�*�����λ��Ci(!R�}�a�%�����A@��ލ�65 �,���w�{�)
��Ͻ�<t�����kۏߣ�^9����7��A�Y�i����n7��oe�v�8�Y�'b�m���>�;������j0t�Rs�{��M�
�*AO��y�4��V�a����0�¤��ף�=3�e^��/5��"Ͻg��Q����;��$�M�y�'0�7<0c�.E���;|�
A!�g���4Lo�Ūܱ@�n�o.�܍ߞ�uj{z����2���4{Kb�oI�&\��ok�2'��Y:�<ySybZ���$�����k��k�/�����؁R�Vs�|�Y�J�G� ��'단[�4{[#H�'� ����R���1�m��T��w��6�Y++��f�,e@��˟~��9�Yu|�uÉ�֤)i߻�d��
B�C�{��AO{����6�i�m) A��ߤYx]�_<o�Tq�1���{�rL�$�'��������H{(W&��H,�S���M��.8�[�}S6⧘tm����w�!���Դ�~�&�Rɇ=����SG{�}�M�K+~��!�i��A%B�w/>�dx�#>q��<(p�C�q
\�Wl��ۗ+��uW2��H�G��m��5�6!x�>�Ծn"p�p������#vk��6��VJ2��=��e�L���ϨY�Q�*j�dA�p�^��H)���d��a���˦ �O�d�
ji��@"��ϲ�ZAf�+)�}�}����I����y8�hQ%aXV��C)&�*K�����&�T��r��\_�M�����z�@�8O���a���`h�a�>߁�t���)h��{�[��l`T���������c��6��t�(*2Q��y�l�W3
�2��k
4���P]X&�Y��_Dn`=��2B��'���j�&]uw]ʥ;u.h[$���/��I�s<��K+)�w�s�J�P?{�d�Aa�w�]��R���^|/���}����uc��i�������f2i�Ĩ�7�tm��k�!e�9�� j��{���{�.7�H>R�g�ه�5ϲ;�<�y�y|ǘ�	��w_w&�h���G�Dw�}�/�z��b_^Dƻ���A�a���s
M%�w���M�led���eO���$�m�u���~���YB��*!2��I�h���Uv�mlg�v���^0�[�-r�������@.�0���Ѭ1{�d49H)h���Mn���
��9�h����~��u�s�w���>�GC����PިPIP����M��aXY�w�y��<|�����x�L*w��r�Ad�t̝34�W�{�c2�YR
;�����65�F�-�y�� i �}�f��@+���g�����[�MBx�c�]���M$|�YY*{�;̛I�,IXX°ל���<[�ǜ��o��!��
��RQ7��̛d�ʐR
w��2�7<���=�1�ˋ|��H,;q�������y�5!�i
Z9���[��H-Jw��4���`����>��֥��a�SY���n±^�fLg�="���6}]r� ����/B�(>��{�-Fk<o9m*�L�C�/�����{��J�C]�����
�����r��a�Lja�<��l�Ad��|5vd����{���~� �B �U�`m�
ԅ��y�d�iHV�lvd�3^ �A�+����ɀ��S7�p�K]����J����n,��0��y���/Z�0���>K�Q�8p��|���Zm��T���{̛�6�IXQ��ٕ�υx�"=�>Ї��N�RpM�Z�M�n2�Q� ���y�m6@ѧ
�qID�г�,|!u�CNRKH>=�y���y�k�w�[�+FH)Ϲ�d&�*Q������g���<�C��W�>@��H��}�����v�6���i�Uxx�C
��u܆��JVKVy�"�>�<	 /�v����
],ƨǼ�N0:5�Z��Z{�w�f���� -���G�"�p��Bf6�d�uԊ#&�����0pI���%L��@���V����,40�(�Ibw��ܛd���7�u~�c���o��ed���=�2M��<ɇ�yc��\�A`�k0�C���~߽ɭ��z}��c�`i�����\�M�( VT���s�Q��RT(�}߽ɶV]�^�Ϲ�]_�������|Ф��m˄q��9N)���9�3�A����[nf�Y�f�̻M;*%¦OP�d{1��U�wh^�=@����x{��w �I0�N���79|�n���@%�#cF�Sl�!��g��c���ݍ��.\��Q9���"M��۟k�>�ӫ���;ngmk0���L��vݷ�{g�͆�^R;!�WO(�z���
�]�0u���x�<g�TV9$5u����v�vӝ�S�����n8�qY�A6,�Z���|V�N��c��;c�KIv��nΙ]Qd���=�]�"-�.�.^"�]�S�����ɷh{/=�hlq\x���a��������§�s�d$�B�X������Q�d��Ĩ;�������3��=�C����]�7H4�+�{�a�@�B�-*D0�i6M  �#�k~�i�+1]��8�}��I��sܛI�,IR}��a��IA
�����6ɰeH,�ߦ�3������]�@��;�ی`��n0�aɦF�q��!��B�B���o�d�AH.��.��;�w�|�K���6�*T
�%��}�2�P�J�C������#�y�s0�L��*|��#���o�����s�i���RT+%e`��~ɦi���
{��捰6�jANs�w s���^u|��} ������M �wc�+��pڐ1��&����VQ���s���I�;���[���5w�0�����w�e��T�
�߷�ri�l����9ϻ�o�Y }|�M����\���m�CM�x�;ۋv	�/GY^Ǯzz�\'ڝvv�"'�b����߸~�\`����;���a���HR�=�~�&�R�
�S����M�T��~�����|ͥ�3�a����%B�����a��a~�7�r�#_ơ����7܁��!Y1y�>�޵\�]c��aF�Z��#!����Rr���s�۞�y �.9�r��R�n�u��Ε31e��S�hį�$��������JʁR�S����6��Ԃ�S����@ٺA�<�ۍ�{���7a��I�|!w�-*D0�i6M  �#�kzE�d ��>� �{߻�`�hQ%H,>�}��:`���7���C,40�*���d�&�Y(��FT����&�m�|��|� 6��!��g�X(���'��q��m�<������1�uܚ�HV�
�R��}��l@��/�߹�Y���kw���OP�%B�=�{�l60��z��1��a�px3�@�";���6!��!R���5�K���c���|<��������&�mHR���r��B��7�a�L
Fq���]\L�6f�V�:��JF��R���G����<�t��S��:Y�n֔7a����c��Ӏ�k��ޜ�E� ��%e*}�}�M�6���V_�����
�<=��}��)=���ɴ�ɱ���T����&�m�fs8��\`���а4�|�3�<wR}.���;���dQ�~
�����i��R��/��ل�Q��<�m}ز }g���.rq�XV�w�;+q>	�Cl6¦<��m�KX?sd�f�
 @�@'�?,��M�?-]+J���u1���h�9÷%���qOc<N>	Ox�i\��k�G�Q�Y��RؑFf7��Y������������-�;�d��R��{>G�"��B�Pi6Y��d��I�~�2m>Ͼo���׹�3�>H,�%M��}�i6�IXV�9���C�aRQ
���}߲m�י�ٕ �|�D}�\�X"� ���6!�Q6hZAao9��Ô���-��>ɭ�@����b���,��` �@d�w@��J VQ9���a�42T*J@[�Ȣ<	�kߌ�<�!��cE֡%�ͭ���M�������אѱ�ڑ�y�����fC�_x3����#���7�J�d��;y��i�d��%@���4���|r\���pL��C�i��~��iHV��}���"u�P�6�M�T �,�Vd�l*Ag>�sq���{&��޻��&ТJ°�,�>�ڇ�40�(!RX��}�&�7Y++'����l����>����Wr=�@D�3���%�L�B��k�5̆��AH[@����hx"���|"'��v�z�L��� � ��
ʞ��0�d�Q%B�w���a�����a�[����Lja��Ly�{��=�[��LzH,���/��a�&���@������6��HR�����u��}u��q��c�y�Ǧ�p5qv3瞘=�?C'h�b���]Շ/?f����j{JSφl���v���m�D���v��:�_jߟ}�������)
��;�|��D/�B�Pi6Y��d��y�_��i�
��R
s�~�M��w���W�۲VaXv���0�
��%O��~ɶM��VVJʞ�w$�"�D)ϟ�IC(l�h�`'��;aۆ��V�#�m�N2PRvb�ԠW��v���1��+q��ǧk_��CC��-!K@�7�2kt�H-=�>�@�/� �=�/ald�QY�_?�|}�x�P�IP�s\��6�l+7�A�Saa�
��|��r���@G�j�ȉ�"�Fܝ�[�>�2|���%@��}�tm�������Ϥv��Hx#~�A8��\σ4�D'ק��e��2�5@ ��H�| VVJ�*}�=�MěB��(>�s���}�n}��������H��%�w߲m�l�����T����H�N9�||n*��<���÷�C޽J���Aפ��C��o�EZ	��[#�>��M�T�e�lv��3��D�d��w�#Ȁ�\ɦaX^�{ò�����6�q�Ls>�!�6�R�>�0��k�ǹ��56�D������m`XԂ�s�� i �}�}�a�AN���	�踹'�M�W����K���q�Өҝ��m;y�nX��~F���3����gp�_M�g�:y`�=8o�������tiQ��;���29�S�A�F�KVņv%7�>�7ʸZ��+/ӹҸ��QfQ�Uܒ���ݞ�
gZ�1cZ�0_%�9P�"_p�r��`�������R��Ox�������/�4o�C��䙹�7\�����n3���<�|�S��0����ɫ|�9�3��o3U��(����Sc�EV쳆g37��p�#jS�m����^�h������/kg$�Y|��R��Qf��Ub����;��.�t��hL�}�dv�-`(r�6�{r�X�
���WI°`��'sib�$o4-�D�u�g{Ӷ��!���M{�j�E������A��a��H�����3k�o��a�A�ڑ�{6�)�F���Q[[�tv=A��(͆��x��^�����F�����}�5����)�~����{�%]�D��2�X�W�/	�s0T��n*~��佤@��A��vd�i����=B�z!e�7��G�l6�#1�4�n���9��:tp�j[SZc��+Ź�S6��������-���c��6���L(��C��*�N��g������z����V��fO_8[({Vхw��}=��O:��]��ң*��{�䗰�_�gl�u�5i'��]:7T���hX���Gc��6��c��$�����M9$�`�2��
�ޛw��\\5E �Ëb,DU[h֑Tň���DW��Ķ�*1V,*UUL0��b#5�(�Z���Q�#`��-QD&�
�Q�D`�iH��D�)�
#+UH�`���d�h1@ee*�"�dm�h*((�m��T��qK�Q�X8�[�b0QF��H��K�L$�`5�8�aSX
,U�-(��DA*���TTTEV�l�*�QQE�%X����Q� ���UU�
�KJEFaU��EP(��b�)U��U�j�m�B�RV%JJ�YmJ�m�b(a�pʡZ�EU
�.10b�J�h���j��n1����$��m��Km���b�����id�*ň��1���U�mTX,T�[��;�߻�΁b9��ny�v�v6�<f�����A<���y�8�Q�:�K��A���/m���, v�b(�����F�^G�;vtwZ�9�]�<#���+��8���vy�u���Ϝꍞ(2=��>^ܜ�=������3�v/n
S��t�6��J�nu�f���Q<�Et�n�l�=��cW5�v�[��v�n��$ q�^kg���g����t$�M�_�f6��W��������6�y��h�ql9�A���G�:Nt����s���)Y|��ܽn�r�(ga6�YA��>��@�sͼ�x�c�q���>_7\����s0��nl����uƹ��Ʈ{;Qc�8��Ν���{Ii�5��7��۵�:°���4�'@���n�n.بr�!vw�Wl��=�K]��F{nE�ˍ�l��|Ͼtm϶}�|�6,r��w]Ƿc�m��ͻ.�ڴ���nz�n벖�W�B��.ݷ':������d��ŷ1��lE�ax�b�&ڶ�p;[^Y�u�^^�I���q=y�s�p���D�Զ�hx�R;a�P�n']�[�.⃉=�'٘�$v�x����"�t";n9zV�62��G�s�Zݷn�Kgo�g�8Nw �ݰ�.���e�Nyۘ�
��N�S�<��?+���t�gtn�;<m�=u뇱��7��wn��{ksڡ�I�#��G��1���F�t��9:Q�����<�p�_�v��ݺ�v�]��g\��ax㬇��q7Ct��v�mÎ՝�^y��[$���l:6Q�6H6��+u)@gz���+�%Ź���rF�G��cx��`��He�J�N�{m��m\�R��&���W`�2{و��8^1P��5�
���h8.ܶ��^���ma7nvv�k�k���\�ex��8�/\��ڋG��>�:�`d]��'cO=�vݧ�{r�3�:��pT��M�q�Ǎ��Nc	[vÅ��^헷[(��P�n�Jr�������Ag;���(����p7.j��^�w{��~v�6�6�j��_\3�Od�Y;]ر�6�v+��q���^����\/lf���K�^���ѐ�q��e7��z��tr�m՝�=+�#`5���d�ѳع	�[q�u��y�9�ܩH���&����;�1���5���n��kx���べ�ӣ���nyNv�Iʞ^B#Ihy��m�u�ql\������p1�n�0�d�����!�v�{�l�ڠ����4Qv[�m�����뮺�NK�Ha�_o��_�e��l��� G���"ɱ����2T�;�rlI��°#ཱ۵���${c�yV�u�d�+%ed�*w���H����0y�n*y�L��������!m!˥ϯ�~�q�������5�`V�
�>�=��l@�ba���f3C%B�*�}��;t���c�}���TȢ<	��t7W�#�����|!��!R�}�a�A@�B ��tlN�׳�,� ��DxS�����HV����.�K�]���fb�(dY��\�#c��s�-���J�*}�wy6�hQ%H,-�>�P�AH)4��~�&��VB����G=�x�A�"�~��,�H�1��� �8�'�W�>�\���B�A@���ܚܤ+��u�;�t���9��&�*T
ʗ߾�0�5*%B�߷�rm����ֱ�Z�?�����^����3m��un��n^�ѧμ���6[M�����7lTb���]��g]e�a����;�r�J	h'��܉ ���ɠ��+#l����z�g]�#m�1!�l��-��FOm
v��]'Q�e���h�IDG�f༭��">������%��w�[��_N.D��4��O�q앆��b���N[��|��A�������=0���$�۸� ��_� uξL�:I�f�BT�Ca(�h��$�ܑ@�"��^�e�@��Ab���oQv�$IܮʢE+�b����Os�Y�wVM������  ���h <>���Q�/�"������8;����/7:qTMÓ�����܁>$wV�p������3Y���}��A�@L�.:'^���*qjBzԗl�n�ZY\�j<��D�l��ƆҀ�p�81�����I$��ΠOod��P��rw�>'��ʾ�'ٳp�"��,�^1}B�&�kn��ً8/���W�������+ݺ֣D��j�7Ċ�(ć	��h�J�F�m
'ǻ�hQ'�.�َ}JU>������k�H�>��s�痴!��8��T!��^>�*Rf�9��o`v���L��:�L�%CJp+ˁ�N^1�3~ϻ6>$3n��D��~�:id[i��Pl�v����WOx�f��h�A���	շp�fFv�/*��)=
1�p��pO�� �;w]p�Xbw�0�r��|s��E�n�AO.n���ɨc��Ƅ0[!&�X�'RƘ�۝F�zݨ�k�Y�<r�u�ؽ��h��p�N1�e�q\6+j�A��ڣ@.>(p��O�*b��Z���*�7��^�>q�0nx��l�u]�uע�vӫٝ������r�I8�3���g{�d����w
�
<a��1@���D�p�\H$�ED�Am�1��G���B�'V�ĂE�T�	��D$2��wSd÷���}?x��r�I�]�^n���}]&��9�B=SLh�����G����P8�%�u�g&E�,<�����u}Qٚ��wi�C�S��{����H;��P��%�L��&�׊?N��շ�G1R�E����wC}���yTH'�eĐ@���y��í:��5��eFv�d�dZ+%m/.�������ܷ�\��>�~�p�����Q�7�j�A�r� �����Dj��*rz�	�2�W��pb�p���^��[���5�8H'ܳ2$�N�_Ux�DJ�J�3D�Λ�ys�]yƈh�B5�gǌmr�;?s gR����1�+�_{ ���I#�/��λ�H�0�d�� ���֗�����H'���ĒHU�T ������fۿ`�E�Ĝ�(���,6J�E�m
� �uu
/"7�EV_b��6�LO�ڮɠI'7k�
�y���q��������5�7��v����D��U�x{x��6��J�b�7ybkb�A��-dPnT�ZZ�Aȉ����1>^*��i �0�B��.��&m�5�VE3�y��m�&�A��W��sm����cn�3�0��r��g�3\�]#�.���ا��ǮMżz&87n#g����89SI���L[�c�_h1�)Ơ��=����F@�bެu�n=��Ҍ����s�> �<��{s��sZ�]�؏n�u�_��9���1;ZI�4���ú^m��u�b��$��pN��tBm/mm��m��i<۲F�p��I��������e��y�X	ן���[�@�	����]}�~4*��� ��� ʘ���,C`ĝ�^����&iSc��ɖ�̒	WyT	�';o�P1�q�poo��� ���Eh��5Qo?%�D����^�݌"�(������'ăy��m�#`�`!�8t뢄����;�=�4	�$����W��s��2���`���NzEY��� �}?60ONM�_�>�;6�	!FoUE�_W�uN�H-�S�OT�AL�("l8-��)����Y�:n:e^�|�k�Ru��R������u��uՊ轮�����$��� O�e�C�'U��ʪ�>#wo�5����[	G�58G6�3�;V	��Fz.0�Y��vr6rנ-�=2�E�� �����9�r=q+�Uoy�1��p6H��E��!�͒4ɽ��Wo��yEf��������Q$�Ȑ	�XC�����i;G[m�!�b@;�TA �ȟ6�����з��T9��khP�c"FE{4Â��Zn*�ӓT�qӓ!p���ʈ�#b���]n9'���s��QV���QC׽B���ɀ�8k��#�vduY�G�V(�{����E۾�@�w��U�TI�n�Wd��ܩ����]��c�o�7A�	�n˶���z+��O�d�]ۥ�y�6��$���|~](��IU�+]�Q$�x�O������Vv��*�F�+]z�$��$�ȣ�4pJ�E�u
�ت�Y���WΜ�I7׎H#k/��)�V�2�������2�J<ᩯwj$V��{�㦺*�;}g	�/�z�N��gMu��{�1�6`�/�F�����!����!%���N<=~���!%޽�:(�_��2���JM_O��ႌAl>;:�V��o�uL�ξ�A ����� �o7�:��j���2�f���_ҍZ7u�)k�&������e-�SL��<,�RH��ʠI��T��f5'�HXw/8���P��>}ra�Ŷ�Z�����j����.���8P����}{��	�M�4��&�/�Q �wd��M`��[8�ȸ<�$�>nJ���ч~�Clw��'^��Z3��zi�A���E��P���ڧ�������)�D8)�ÂT�/���n�cN!mot�����!D$��`�yݴ(������I��T	ݞKN�U��ŕ}9��z�6h�	�wmW�:��)�T6��t�C�S<�`,��!eը�DH��ܣ9�uˈ�qx]���%�
-�n�n���*��×YsJ��x�}�o�TwKi��F �
/�g���o%�$%��1���s�B�s�j�${V�D�4o]���~k��~���J:'$f�c�÷K��C�۷SX�	�M�/]�a������ٜ�&�{��U�|O�v��Iշ� ��Ǝ�����/g��77��Q���	�M�8���IW�nĝ�ē���[�H=!�.�ݬ��'����"	%��*�Ǣ{(P'�K>�Ę�'�D�u���s�s;`ov�P ��s"|m�!�XL"3+�7o��$�c:��k�"I'�w}K{�ν�����;��B���Yq�	?8j���R�۽�d�+/&u�"��t�NcΡ@�[�;�}T^�Q�%�r�Ͷ$��2S�1�m�ܙ��w5��Z\�L�V��>���N[���L�ky�.�Cn�y�C���?���o��F�]Q^�S����ꔱ�[s�lnڹ�碎�o<Q���������]a6QG���3�7�A�l�[s7Xӎ�dI��-��ћ�G �ׯ]H���,����6���-�+�3�u��7kN�q����w\�x�t�z�s��[i����N�7�ƶ�Cn��օ�]��Msy�G�>ۋ�Ӂ}=�mQ�S]�Z���N�^�\21�u�VN�̖V���l��mp�Y�]8ڶ��ݎ�D�K���߿���Mۅ�������D�;�!���M�9 m_��kzn��̉���i�D8M4�UtN�{h��zm2����O�,́�z������o��+j#���?��V�L!6|L��'g��	7�}5�A�N5��;�YIǳ�	'VfD��{.����F�!�Il�J��؛���3��,>$v�$�{.�h�Ff�T�}��MF��'ܳ.$���"`�p����Femm )ϟ��{5��3hVM-�U
I%o �3����qn����n�㇕��穵�$�r��3�E=L��.�\6))6f�p�M���i@I��[���Rω��f�O��3s�����4S*\��w�@�A�h��2��.Sⷺ��A�4��g�syK&��w��8��<������s�{v�_l@E�&�v]�=�qs���B��r?g���J[��pݺ�=�E5���m-(e�� �y� �~˿��g��P>5���+�R�f������d'"&�n*�'j�Ēww:��]%4�0Ema}�q>�]�P$f�P�_�&�(!	��d�'b�E\mkXQ í��|H$^vuW�$j��w�}n�ѫċ���C6��B#Ų*����D|p�d�Sp�G�nY]:$�������s D>�:՛p��#aPr�%�K$L0pN�v{�fv*�\7&ݎb����ы�a�}}~~!�^l
���@�7��P �5nd�.UYCz�'U]*�$a'{s�����i@I��U@��R�69����2p�Iwo��>'V�D�A���j{&��SuS:�&���Ap
{g=GĞ;�,�k��X֓�&���Ũ��f�6͞,�Q��-9�)�׼-�*�'����쯢���4������Ƨp��&�R���b�j`��0񱗙/��̑*��<���C�*=ܮ�p�,��n����}�qc���1,u���/|�_.�D�ҋGڜ�ѱb�Md2��X`]ck�|0K���څ�KZqU����w��0]�z)��8(�B��[ۧV��\��C"2lm�Z�ΗbS�Z�Z��¶0�|����/h��Z��Jҳ��m��X��}��F��Dp��^�]�����m�����9ɕ��A�s4��2��ĵN�j�Ϭđ��u�/%ۢ�˺�ΏO.�,���ŉ�a��o�٤��ؚ��'�$Tn�d�����$>��3�nњ�tҦs��IM{�-eE��LQ�LDz�JS��S������d�}x�Z��7w��:_,Px�:0>�3�s�Z����?I�7�0��L�7�ݾ=���2u�r ��J�������V��s��]�h�KC�nl����r����Cx[џo()z
��5^Rc�>;�qF�g��uDk��cT��\�⪾��.)r��h ���T+E� ��;�T�7�?s�#S<���㺹z{3@�s
��V�y㑨.�?8B���[�������S}:�+/C �*vI�������j���Dߐ1}�f)`��ZVX�JT3f�#]݃n��w|�WҴ��w�2��o��'�w�-��}�y�_����Q��*(�QkEUT�-e"(��+b��H��l�Qm�UUTT-�b�J�QA��Y�`�"�EATEP�Ġ��5��b��YZ�1l�V��`���E�EZ�1V����65�Xa���"��Ţ�F(&�p՗��Z�1d-�+
�Z\2�F*��Tb�lqJ��\ba*��#0�pث*
�T�b�11+Q"ĩF"%�P[h�j(*�V�TXyl<e�0�P�*
�*$O-#Ap�mZ��IU�TŅQ�,|�S�A�T��Z���Pce�(������Ua�U1lOt�yٖ>����Ex��Ȓ}�^͇���M�WN�S謪Ȝ��M�'����Qqܸ��j������I���+�d��0��2�y,��uY�;��'���=�B���q ��Y��q��5�.zk4�&	����0�61�?3r��v�F��8�\-��ʵѻa����7��ڷ[}�'{�I��$�OUgU�C�C�ت��-�m
����A.�H��!�^l
��Ϊ��RL��1V�gU
��4(�H#6��$��Ϊ#F�qU�}����ϓk�L�J
����������B���;#�c��tI ˷$��Κ �Q��
 �]�
�o�d>�	U�L�A=U�U�	���YxƵ����,����E��1A�K�mm��	�ޛ}��"�:�w�����s9P�fg�x|s��$�V���(���qT>���$�y���F�
��v���}�[�+��w6��(׿~����ߛ&y[A��u���ϋ�izRwn^:-B:�\DU<���E�Wo���lq٭�j3��A���A$�mu/����d&G2e�9 �Wm�Rf�i��S�.6�h���{�.��v/7X�H�ڢI7�}^�|U��T�ӬH�s�H��"\!�d���E�uPw���D�n���U��1��$�n�k�o�:��:.���'�W��ı�[�(�d�I���O��ggUA ��37�T��;2��ɢi���p�\�x�>��	#��g-����H�;�+����u@�wk�{�$��1�+0ysR����o�&+�|M����vq�4�Pn(��K�w(y�O���
JjY �9ҩ���y?�q����k�-�YYӨ�q�8�m��ֱ\q�.��*�l���3m����F�����V����7;v��6�sض�뇎�6���N�� �8��5Ɣب�OH�3u�Y��mNTݸ����u�[۴�p��n5���sn�0��-6v6��K��+��{P��D��6��8Npvw���\ǃ�m��ɱ�!������ڎufxL���ع��Ξ���[�o;�;���rt'k���_ߟ����b�i����B�3s����9��wv���(n��Q �ٹ�(��t���0��2�z����r��Z������@PG��	5��&O�["9�}m���n
�PD@%��%P1�ӄ�3k$I�>+�����Q���|{{:�Aݬs�jg�-!�d�����J�l�yD�I����N�c�I�}QU�w8�mL�^'�*���غ�T��5^;��I��f�3��T����ʿssU@�/+�}�w�F�Nn�h#��^�L�sø�f�Il����{
��Ν7�����&	1���لb`�W=D� ��w�^828s��Q��N,,�=��M�c�FEa[J!�e���D�P�oo5�u�i���n��M��'s{s���ho�P��疸��M����¤��*�y�&b!,%�C�q�Vт�ĜTV�i�9[�t��I��H'��� \8�÷Gb�>�y������}���I�>&Ag�A�}4H$�[�H�;���� �yX���w�;ј" �A��<S޶rf��n�� ��� z��k�����x���K�c	=�.|Hٟl��3͘E)�fWU A�;��=ؔ�{j��d�����yTI��B��t]�Q�@��b��G�A$Bp^�n�.�=������XG�6,�S��=�����������?8k;�.ڙ�������C�E�Y�[CtI�n|H�]�W�^�D�h��0�S���|g���>u34k�$�H�ʠA7��B�<{�:�_�����k�'�E�箃JZ�V�	��oy�	$�� �o�Q:t��ͣ��M��--�V*P�|a���|���{s�W#"�o��P�s��U�n3��+
V��k�	ڲq[�ݮ�WZy~=�WI��� ��w�@�I�߶V?qm��@�ω�:���޾6�
�A��٠I ۽�@�v��ȋ#�EGPD���	�f���ZU�z�Q�3k'�7����4.I�ut(Nwvר	;��L���œH����[h���2\0݊7��=4�hn�6,q�'[��ӳԝj�+}��{���ay����g�H#{�j�n�1��������w���֜,��iǵ_�"�2�$�᪯�j}$�;�XB�]�O�hM�vȯ�X�i��mGd�V� ���&�����R�s�D�;k$Ie���k�9�$�ݵ���ݬbFEYZ�n!�%��W'�9=|"h���d��3�D�Oec�A���V��ߐ��}��4o�O�W�!iB��X0��zl�3���7�Y9������TO�}��u�� zD��N�o�ن�Le�Ţeյ���3>�p��W[��i��E$�>&Ad	 �Yw�J�u�à�<���|O��c�	w}U�N[��7W��d�D/�#�2Pnq7�/����y���&����&���˞{=]r�����;��"�A���:�>#:�|$�@'�O���ď��'�ss>�� ]]�}s>|��/6a�3+������u�c+���$�c�I��|uL{'�';�%;W+���p���[m}�`=�{4H"-n]�$�wٓ��Ouc���U)�B��f(N
��0�5۷(�UH�O����	"�{\���S4�y�G8G����5O��Æ�-��bv���3{hS�府N��|\L��Ge�U	�{hU<8���� �W��P�1��N�.�T�t����\!��m����ԇ$1oQzf;��6?����Oz�L���[0x�6�H��g6��������EXa�if��k��X��8�b�k�]OujO.^L��n�pc�䋭�ֶ�gO��Y�h�ۓ\\�Ď��	�E��Ë��ݩiCv�u�b�׳���pz]+.�]���<㺰/ciz��<i��x �;q�+�Ou������v0�â��˳g��M]���g�;pͦy�u����=y��{X���8��Θ�ݙ�Nv�s�ۋ�v�Ꝏ_i��L��@̗gi���-[��<��D&��?:Ϥ�k.�h�I7��T_8���YdAH=�.I�zJ���#Ѡh#�l���~�V��B��$�M��Mx���ȯ�-^�;"t�#�O��>|��/0���F�uP�vУ�|�ּ�W1�E�<�յ�D�A���}:.F�� �(�0�3���n�@Ͻ���{��ĀO�׸��o1��P�-��H�T$�0!BpT��L��>�>�yyblg-�PQ�S@�G�ovW��qȈ#͕p��Κ��׳)�D�P
J��jZ���<'u������S.��Ӧl��z���<����pe���Kڪ'Ĝ��Q׸䮍YB�<'n���"���ow�c��o��g���Ϥ��}�eF������1SK"�#z���r�2E�H|�T҂���6���i�[x0��=�ׯon[<s�*\�GLm#��ʌ�a�?GN�I=�}�^$�{�A�ٙj�I�w���ۂ��$�A���ϵS�<T �d
�0����<��w7�}^;��A73�̡��	I^ON������Đ���u=T|H#:qω;w}7D)�D��Ƒ�"��UNgPʀS�MO�d�����׌��4�XȜ`����$��� H����ۼ�����;�?;i���ѩ��!����n�	�Y�.�wZ�pmtK�7�S��o���X�]�N;u���v�O���}�w�-�B'����c�(VD�P �w'��ɽn8nl�^蝪��ٖr*�R�{2���rH���Q$i�]�s�c���ϲT7�P��2�z�˾�@��vS��$aoE@y-�Y�gh�����6���fhN
��)
�v!Y�o)�p�#.��y���`�z�<����O+`���]�g?u��~���S}��c� �V9� 6���eu@I5B�pN���qw���gn�6�t,��x��n���A����rI#2x�DϘ/���ze����ay��1�[B�;��^��*ek��h���$�w�^${���[]o"g{j�E@��.PD1��\���GTA������3ZB�9+�h1_����z!� ���!gT�I�{4H�{���jp�l�O�����A�S)��Q�Cz`%�Ye��	�y�@$^��W��&�{d
�����w���L���M2[-�V��UA'3{h
$���Y��Q���Fe_P�/��V�s�o�P��8�z�.�׻5u�Wy���s��$�����ǎӥr;�з�	���zk�?�'���=��aA %�zi�}��[����FP���]ޝ�ze盅x��&�����G��QE x��9��w����j��I';��w` ���D4���茖���_Ϗ}~����]�b�5F;��pf��Lgm�Q�;b�4,�!��ECEV����Z�	��{��]��;�� Fm��Eyle{Ss�~���m��Ȉӽ�رU�*&��}U'��N�m�G^����u5[9pz�ϝ� t�l���ݼ~d��ng��S��^�����RĈ�Q�䃊�O�m����w����6{�+���� �FOv�L��禒AS�\6�&Ke���ζ�ob�Y��?H�<j�@��x��Hs3��Q��3$����� ��KL���׈eCg��!�v��H��Ϋ���x�V��W�m��r�@�o^?4����+1,sQR�m����k6�A5��yxFpE�C�`2�:��4��!�|1g��o.�+�،k��ra݃r�i����4�v��j��2��i�f���zs�9��Wr�^��R��i����7'���zrㆴK��
�=��[M@)g�f����h�h,��vު鸕���*���L�0>�-�6G�NFv	�<eXIK�y����чmm,�j��]�,'�fL�7]����R�	V5�YL�W��c77<�-��fK��xr�f�<T�l��S�|R�V!+_W-*�l�n��ӛ�z�1��TMl�5yW,�H4?A�z�O�u�Z+;9?XIk����w��И���3x��T*��X��G���r5s���>�͌��=��t^B{	<x��M�y�b9U����1�����E	��8��#X2s�:/vNû^�����{[��*�{�gD̋7oybq��Yx=�|s7J�x�y��R$�C.��է�9d��8/��`Xr���eT�wƑ�]�p��Xx��,���K놽&%�۴l�釪�չ����>KS�b:�Q4{����4��(/1	��d��}�k�����\徸��캓�Wq�+_'r�t��WZ;�5J�5�Z���v�״zW�;#8���sy��{�N�q>mr������$�쳡�̡�[��5���P���8ݱ��;.�q-�Dr��¦S�˺K�����Z�Ӕ�?"Gx�u	�H�H;�O��V��U��OuN��C�Qs4�W�iؾ���t�}������ذ�������d��y]0�x�)�X�a�F�c-
�X�"ʠ�b���խť[kUb�)jP`�5��y���<�Y�x����ʸ(�*����F"��ep�#0��Qb�m
��V*��A�qd*��
[DY��-b"�kE�QX���*&-�("%J���%�+
*#m�lYV�����jւDQEX�cj�J�AX�UX�Ŧ-Y�Q�P�>aTATUm��U�ATE�l��TbƲ�hQU�R��UB�DQTej�*��1��i|p�`�[ePX��a��� �E�*¥�"����O�"&,B�E�bDb�<�6�yǽ����cH��e�����������w��gK�©�tnAj�/O=v�� =��n�cq����q]gZp��O��Uۖ2�����mZ{B[�n`%�7]�9|��>WWFH]�1v�3������� ӵr\�׳�&�c�:�m���6�=]@�;v�;b���yӻ�����mp��^7<o��;�絗6z�B�`���=�ĝ6M�Oj��\۵��x�w��A	='�۶����qŸf���ɽ���qt��=���t9Ň[n�)g�d��NT���`rrg�󬳄G3ו���ĜL�/���8㗝�n͋��F���83\��OS����t�H�Su�\7h9L�ƍrn�u��o����O�y<��Ѯ����n�ӱ2�s۲�s#����5�Y�g^�����[�vĭ��Rv�g��ܙ:y�4<�㰈H�ݷ\�$�]Y7cb�=��#����a����^��<�]o\5�k9�m�0O��!ô����rv�qb��<��\�ns�,��Nl�/�k|���nǰ;�m�]�N��D�n�n.���%���Z�)�x�u�򝗝��Ý�r���٤�RV�ԵB$'�kt���ے!vn"�nwg8n-�lv�W!��ب�m׳m�1���>ܒ��W�6��l�3ŧY�n;1B�n����	�^=nL���M^"�^Dޛ��C��/L��Ζ��]s�Vunsh�rc�7'k��-��m�;+����n�n�Knz҈m����P�I�ݨ9��	<j�[��S�ۑ�ۧ���{ns�!��c�>GØ��k���;xӧmö|,��ܛ��G���z�n8��t�Y��3q�;;���۳ڍ�[	{.�v���Un�֍�8�8ڇAǣ&�r2���9�N���d������ �<�]����(�Z�ݭ�Z3�{YF���󛎌kÕ�� (��.{s�MVXݧ+em=W�)��ρ�#s,�<݃۵[u�3>q�&��Ti,`nء��5kM�烪:�+���Bq����:wo����m�D��˰�&G�5��'�K��F.�}����F-��n$4<��� e�C��u]��u�v���������:�n����g�<�z�j�w;�z/mƗ���'m��Y�2!�;+��z�sn���Y���v�s���x��f��{,����3պ:���8:�q�<Qpܨ=���і��K�����S�Hq��=�rZh�R���&+��������n7���	;��` �o<��vfuݠ̇�ɺ���6�L��t�@��/��
�P46!��%0T�����I.��.��n�t��Tπ@}����73:�֊H�*ھ��W���E�^8��J��M}U#�Go�� �������td�����B������v��D��l6�Al��ewi��0�ݸٟ 
��͑@+�ͻ�F�/.A�s��qkɉ�`	F[��p;wRGJ ��g��F'Ēi���M�:G�Ob�6��I��k� �3v��w����z#��ϭ���f�眦�Q�f�.��n3t<4/�ttۖ��33\��~�Y�[��s��ʆω�C�P�H ���v M�K�gnb0ݨ����5��4 Gfv��1�]�%HQE(D6{y�`k�M;�E�i�J泫{����²�y�����opyMW��{�޷
ɹyE��Sٷ�\[Ȭp�� Ě��^�w��{{��ɀ n�mݠ 2oz[ �����&�:�6jI�<�����)�-��wa���:b'֊��~��y��^�m��7�-�S���d7
b��U��ku����wk� i{���F�����/϶��$��̻��,8�M�ш-��yu{0�v��b1n_9v��~��7�l	�'����d ~��xJ�.�ů�~�����1Μ�L�I��f�qm��ܖ�)u;��J�8ҝ�%�������!l�K���k�ۻm�T� Q�x��z�q%.���]��=}/�
m�:��2�k�����	Dѥ���7���v�X| go��D-�~�|���W]u�V\Yjff��b����L@|6�ކ�#x(��	�*}P�m"��{Bg6�v��@�as+^\��W/]:E/����y2o�q��j2�}�W�G�-��:z�Zh��r�v��a��L���oe�^w:��>˟0 Q�x��H������b����g�K��bMx�q�Ai��¨��v�U$�={�NQ�yr��>� �mܶ �x��D^�ۉ~ɫ�Ʋ� �2I��P��Yvq�4�Fà[���H�e|�7&n�A�튇4po�l6�Al�w����:^I�m�ׅ"I[{�w~INL�n����.J]Q����_^??�	<�:��A�7T�����KNJ7��:���v�?4�{�wd+'�"O���I��eG C)��MR�j� ���Y$V�L/\��X G�+�'�o�2l���"��D6o\*&�'�=��o����۷v� ��ɣ���3s��e��}�3C�J�igvn��[ٝ�B:fFY.4�ܨ۞���X�������4ǒ�O�]�<�q-|r��T�Q:ޠ��H�WT�OU@��m� �`���.ŤD����S����U�$��]I$���ۢl$�F�D���
ΒN-��M�����)�v.Yy�t�+h����a��c��'#���B���!�RZ������ ���v7��}Y��0�d�� �)m�mѨ(h��6#[3�{U�9���0*n�� ��^����;�/�DBy������:���j�%���|��O�9�0��LH")<��U�o�Uy��rI���݋E ����ȓ^sdQ�⦪~�o�u{]ߺJ��Ȯu� �n�V�iݓ���r��|�u��z5��IS���Z=f���E��B2J]������f5�Cen������˻ >F�vKL����ݭ�7�����8�%c��Qs�ѪE�^��Q��:c�XF��m��2I�������<4�<XX+ խx�>ՎZ���z��.gFΜ��۳�e�^�zytN��^}"��m���*����I��ˌ;#y����Z=9ݹ��y� ��G����v�<�O7;��]�,N5�/<���B�j�6��ֈ�/+�bۤʻl����6��1���u��Y}s����˻-՟5����]���!���綍��jy)�p/k��l�=��G���ڜjZ�=+u�0�f�c�����+}~�J�T���SJ&�&�m��8��L�7/�ϫ ~V�ݜ����ӻ'��mD\�&��*��N�~�+��<���l�^Uu�I�ݑ5�Gr�H%�lLM��on�����y�UH����r�+��8�m�a�Dfድ{]2m��^$�AdodI5�����Ur�p�
h��Q�s���:��+�i����F���� ���u��S�]���+�Q;Iy͐eFx�ˆ���9��RIw��~�}�e�����휾��׏� �]y�wk�b��ڬ~1H"a71��|.N�xg��@`���<�S=����m���o��S$ET�"@^��b u�`��;n��R߼Qy�.�i5{-&A$��_<$�*�����:t,)�*���2OA>�_M�~LN�)$�~�*�"�>��s �zn�� �6��Ub�N�~u�E�T�˺���r�@l�jD�TF�NtE^)ۉ$�[W3�$�^v��(%�K5sE�9wq&�<ɸࢂ�*��cu�� A׻��#�S^���v�����//� |u�mݤ"�i<�&�i@��:K���[�.��{�� ������>��ۻ��2w�"cp����z!g"NwU$�UҡsS0QU#���� a���wE����{}��  .��� �;�IК��N��ѻL4ÁCp�d��u���b�=��-��dN�^��bū��~m�;�K.�]��9ړA$��ڻK�!�N�Kh;6-\d�g�R�o��	 >:��Y��%ET�"�$ޛ�	:���#�t{;"s�̀�=��@ ����2�k;��qw�r.��zm꬞�I;�K��"�a:��uG@A�vO� ^��l���u�~�������;J�fqE�^�m�?{?ܭszE�ao�U�ɭ�"�D�Pi�W.v�+(Tai��F��c5�Fĕ��r ��ݻ� �7�[�J�Q4��ML9b����1t���c�w`7{)� �x��X<^Μ}s~@�6�X}6�"6�J�PJ���u{k� �v�y���ƺ\�o����� �7{)�� Q�x��®��H�ō�@p	e�iBL6K��s��]m �㶦`ӹ�a����oa�����7M��U'���v�Fwey� -��y��2aΤ=�b�I/%���ל�2�2H0\4�&��{8)/% L�U�A��Z���I9��	#�r�$�KQ8��ՙ=�l���1(�*�#��G{��� 73ކ�A�;�L���� w��d�^�??�
��z"�7&�a:��ub�"��)y���@^�k�@|���膂5�k���ނNʩ-;���<�2�<UZf��!�8ܯ�7������._�)��B��f��K��Φ�UDЉ<�39NMTp�e0�!E!�[i�=�v��&���k:�W�@��E�c�@$�{n�����v*ca �� D�Qm&���I��͞N�9��`�h�d�n�n��c\�p�a���������%L���'��� gfy�@ ׽����a5��Q�C��t� 辵��Oǯ�@n�+F���?�?I���'>���	S]�� Y����{�v��|����l)������SJ+�%k$��L�j�Pzv�ҒK�[��v |S~�=Y���ٺ� ���� ם��̸�-L�*� ��F�]�Y>������x�{[�#w�����~�����0>U�S�� �h�QA<�ˣa$;ݎR�'�?�ՠc��v@��7{R����Ol�P���D��e$t���c��J9�\V��o���f�5��$�.n�h��r0|���:����熻z�7�Z^��Ԇ{#GMI�mgLÉG����0[�u�m�۟R�kI����j�:�T�1��Ν��.���N;�p���]�S�rX��;�*{7���n�i�CXg�K��b�H�wf6��;�A�1�{R�=���]�z\�k ��x�������1t��6㎓b�����C���X���K�N[	��R���S��/Yɻۢ����Nʅ�֜�����kL��c�V���}}��~���.ӹ����Q� ���V  n�Sh&*�^�a�����L�7n�ڝ��-�ʁ�2J�&�	^���w�dt�E�z�"��v�� 7{)�A�a��hb����w��$�𕩓b"iL��s�������� }QW7�7غ{+> k��q�Df�SL*}�W2H!�j&�<�N���4����#�v��a��>h���tw�Q� ���݁�
ƈULA	�o[J�y��x��ML����}�$�@&�]y��I�_J���&A���4(N��i8D��.z�'k�e��.����P��뭻<�/d2�>}���ݧ��*"�*犽��V  �0 >����<�:O:��Z��" :w�Zi\`�e0S�85����R'v'J���t�x����f��b�!�vG#U#jy�)˰]8���x/g�{ e��MiOR��E[r��!!�{s�]h�����vEI#�yRM���]���`����؎'��m�T�C��q^�L@ Yמ�0>
�����h� 7����=�{�fA�S& 4�(b�]S�ca����`s���� ��7/� y�q�mj�X���d�#&	3�\��z��p���(USDmk��`�Aw����w�{���3^g��l Yמ�H����q��͌zD���LT�=\��W�:s�Wms�ohy�<:�[gc�7��������A�QU1,���y�FF�y�י�v0���!�9�g��i����������TA.bs_=����5��7�k��	S/k�������d �4?���g{i��j�s�f��}50哦�興���+�+�]1Y��"n�a�`U�%�V����.����43��G��b�,b�^a�1��s{hy	�꽰����������Wn%L��YW�
 ǣ��tUɁ��F��{�0�X�\]�8��ʸ��4�_nJ�'��N�r��Y|n���س�������5wi��﬎9m$ew�*:*��oAr�Z��ׇ���EvW��y���\��Fǡe-f���Z9)���+1YYJ��Ai�)r�U�Fv�������+�I�����Z�]�\���;ނO������	�5��鳚P���ٽ69���	P2����F�c�"s�i��G�c��j��9���FbUo[dvfܩ��:�$6}�Gֱk�h+����0�x��d�1gU;��X.�'��|��I�e�]S��ݪ`J�<Ef��wy��p��7Y.� x�d�D�.�x�s�,��6�x��_&/��H�{�.$���@��,�{�����K5�gz��J�+M�X�;�nl�v�s�:	�uˣv��uS�L��r��uZo���jaWo3\���X��\-XV̤�B��j\^�QQ��N�1ڮ�0�_:��^eBFHYaGD8�60��<<UW��0��rz����1-9�$�;D7PC�gmdgn�fc�}�zu>�F����z ��VU��i	`�N��%�b�.��qL�4	m����f��G�x����v�Q{7�>�Or[Yq1I{�kٳPv��+a�cm
ږ�Z��X�,EcK�U#��(���DUa��E�J�DV��"�+X�mQKe1ep�#Tbƒֶʖ�Lb�VکZ%l��-j����!J��mJ����U���E��8�kF��J%�UѵZ�ʵ�RR�J6�UmkkJUZ�Ue��KV��qmC1� �Q)l�[kqq0U*��J�TX�Z��k-m�"���`��
�D�l�Z�����n+[-�07���L8¢��-�S��5W�jUV�+УR5�UE������m���
�Em��,ALZ"�K,J��-p����mF�1�8+�Up�Ubƶ�R�F�#Z,APR�m����p�U��pU0���4�����*�qj�J��-�
���0�qCp�{�v�7���cxی�(�D33$�G��)����ez�	�����3|�Y��CtjA�S��7�z��;�PAٙ�v�����-v+��m��$fo:`q�jTL�)I4�F�ۻ�Ȁ3g����Ή���X
��t�@#�3n����g��ڨ��d���
�R�m�:7��\�&q�G�.v᥊�aOɘ0`�{F.`���@����1�g;� f�h�W�o�!�E7����bqcDSBl'g�ˈ�v����x���|D gfm�E��]�d���=���dmo�� ��ePJ��
QQ���|�X| wOi$�K��\M�ʫMv�I��g]�+���?�F�W8�j
PW�SY1�ܯWz�"�'$����� �v�F�@i���}.�Az�c;�)�Q:��Dg���?f�y��#�w�H�;�7�zTx�#��.����o�:���b��1Y19Rm��5��u��=f8`�D��n�2�h�՚��7F�T���|���@8�3W��[������-n�h�dDM�t���>ǈ��P�8��0�Z��l�ف�雉�]��`��j��s��b9IN�x֒�������h)Ґ}����E�l�����co=L	�t?e�z�����#v{F�W��+� �؇	�\\�P�J�W&:��su9��� �3k�qi�����G
�zJ�w3#k*�%��*PE����	��=����^"�[��Vo_z����v��h��:`V:��Ah0�,���hksU<.S��@ �=�X����� ������C���D�� ��z�q:�2�)��
mUzQ(%ۛ�v�"z׷� >ޭca,:��@|���v��S�3�E
����W1nQ��q��uPֆv2y���K1B�J5]\�Z���Vhh:Ŵ"���vT�K��vd>ۇlx�;76� ��V���N\��α�ݦ[q�s����:�ڣkSh7����GqƎ�y��1����$x���Л0��8/;jCHԻz��;�����{F}�vm��^y�X��W"�K=��@�U(*Z�H\�n»L���9�.�m�]	�^��i�.ݰ��oBa8��{w<X��\���4��|�|�Q�]���4��@S����9hy��&�[�qѱ�Fn�������}5M���@-D0IP�p�=CL3[j��%�'\������5��s;n�'�H$Q>̵z`���4�>q���q�zQ3PR	� �:�ۿ�l7������ԥ� ��x����v��O��zµ'd�s�t�Ԑs���	-�q*!�D��< �v�� �/b��^���9v�p� a׎� ��n/���AA�����J6:���]k�4ٍ�.)ߟ��
�;n��]��5��f��W�;@�d�2J���-��R)ED�'w���t��q�W
������π�I�n� >:���Ȃ�k�UK����E�0b�r��bܝoc[Q�2�ӊ^5�06���0g�:��\�if��O"h))����c���{��'�@9|�R�ĝ�pM{g{����@|כ�v
ncHꨚ)TL�M2-~y����W:O*n`A�i�b&���7����z��/�n�y�e�����{b��ꇳ8ͫ��ja��6F2ח q{�Aq�ޔ<k,�j�i�����_n��� ���""L�Q��k�^Yfb6D��BM�_��� �6{0ީ��s���S$�
�;n�h���k�UI9��\���8�M0�cBr#s�VXI ��_;��7��m �x�y�[��FA6�w��Z<.ұKm�4S���Hy旉w��r
�י������"�Y��� �x頗�?>�������o���^<5[ [3]�ʹ���Yn�ls�:�-�\����	\��������uĢ�	��V�e��A�9�K>�J�$ʺ?Og�ٵ�~��0��Y��0J5z�uAH)LTæ�1�����goj/~�W�u��;� @%�Y�h >�/0w�+��eT�;[S�3֢��y�f �j]y.q֤�	q�ɯJA%��⅞��UF:GD��R^�����������6��W���P�:���S���c�f�*<|6��v�F�W��o�"/[3��g�D�Y�d���M�2����2��4�q��k�Ǳ�&F�ӈ�.s� �/?�@#�;m黁p��0I۾T)!풱�	0�5�����	K�{��v��Ψ�;�d�HYu�6�%g^:` >7s��Y���@��	$}b��2�"ÀBL���P:W<�3l�]vg��ny�r<����o�����q��?���� ���?A}۝�v6�s6��e8�[�E$�u�:���T�Щ��	s����;��T^c��֥��/D4���v�#�fXW\R�=3*�#�l�*MAJb�A��x ;su�� vZ���n�2��Q�����4���b��RQ�Æ�.�A.q�F�b���W���1� ���gfu݀�Y�UD�ﮥB�]���k�=�KI�8�+e���(�EЫ � �u֧J�`�i�x�rV���oQ�net��|kO:��j��SLd6cf"�m�4{� Ӝ�I�)���"!����cz�� ͞�-�M���yٱW�I��M ;o9ݐ ���=���{Q����+A<�ʱ�6�t1m�'�B���S�W:��<�>1j+�������s�|������ ���H ͞���=�3����[�N�^I+�ͺ7��j`!EU8�g�K."t�5���}��}��@����n�A�]�h��V��K"w��Nk'<�*2�h4R�PK��׽v� A�=�K ���&�4�T^2u$�/:��I/,�ڪ����*L�̺�U[=Բ�y�;%�r�m�7ݮѿ� �oU��1��8�� �v^;���Q�Æ�.�^K�WP�%���Е�:j�x���fv��� oWh�dACV�S':+#���	��.��Qoܩ�	�l�����=���Mn�������p�׏����8�y�7���e�e��1�.;��>\��q�r�|���'Q9{��c4� �5 ���"BU!�w4bV��`s�����l�s�nz��)���]���{f,t#�3n�v��
��۬�%�Wz�@�nM�ݳ`�5=���.7W��;�.�=�E�4��ˠ��hx<�������z�&��3w\'>��ý�[�5�u��G=�=�6:���o[���tN�瓱�]vu��{&9��Nky�����!�4�7�O]�����r�筐P6x��X<�lTZ�s���	e�Ͽ�~;�+�r��e7�j�"3���H�/4/�<�a쾻� @��z{��ĂL1�ˋ���aΉ���x뛻 >6�F�A�����~���P��\ac�B��A{vz���#o<ׁ�+�� �w���u �F�v�� ���MY.zjfjU"�TA.Z+{��c�}��h��*�m ���X� ï?��nv�����Jb;:.2ˎ yY�a��	��)�b�G�g=)$On��d%.�e�B�f`v����x須�ݷ�F�	���
G��i� �h��m1�n�6�E������v5�'no0������NWT�rς#�o<��| ��wh)z�=3��-��d�^:`��=
 �"IQ�s����� ��������~�v޿0��.
�����QH=��.TɆ#[���B�������T�L�rc�������,�.pE(ꉮ�K> 2��@ �۶�- qXո��Sq�]OR�Ix9���>,(A�ض���H���+" �q�Lu��Јw^?0	��n0�c�B-����Q���rx�]{��L�2{%� �{v��D;�>�Twy�W&��ۚ����n"���e݂��7u;%�w��	�o��	 v�݁h�$��7�$��B�D��?#,����ۡ��t":r[{Nu�0�M�Ά[P�	��'t8����Lk�#:�" �����@|N�ˈ�����v��idڊ��x}��`��l�*`�&}^A�=�4���V@��o��Fon�` d�l��_vD�Ndx�^��>ٯ$k�:b ���Jk˜���@$�Ž�4&����q�^����v,TB����{oD����$ߛ;;����I���|�H��X�Պ�=:.���Y	{�=AfY�p�����Aˎ���p $fn�@|d�l��W��D����T�;I�CLFj���>��� �{�[@}��x�ލ;��WLOu����ۣ`d7fKŶ��A��>� dm矂L�Y�m���W��wh ���̀�^:��R����rnL���R����^M4�6tth��r�U�vU+�������ض�l_�}��R�F��&�����݂@|��y�a���%y;�<�<�됢r���^	 ��j�R�����v�]wٕ�hő�שX ����D5�^:a�2W��N�w~�Ss�N���C�qPODOg��Ii�ɩH$�#��^o�y�#z�F� e㦄��
`鈂�a6RUAs��}��N%F��w��� ��t� ��ۍ~���*�,�Ӵ�g5{��n�_2��Ǣ�pY�{Ist���	qiM��/���4���vN���8'|��=p2DјYG�K��Rh9�1Ē1�{9�I$��ڢ�]Eɋs����t�m �u����DQCz��NZ*XZ�K�Ah�����s����+[�u؞���5��a�&�Y�������pz*�}��zzܰ ���? ݻ���Ջ�Od]��v���%�@��/)גG$V���E���)�컴H��T�u�w��0��o0����v-�h�}0��+�޼ي�$�o�9�%(����1�n�!�����"ä��dzy�G*�ʖ� q׎�D��۴����5D��LԹh8���5�k�$�v�Y�$J�����Iy%񓽒�}=�g��QH���@!�<�I��E(��;޽���饱m>�13䗄��I4��ۢm$�7�(R��vN�J��	�w�U��j�ގ��s8�7��:�D�NNB2�4WE���AޡBL�|4T����y ���k_f�&U�͛W[Hh�d����΄R-F��OE�E�T"��P->ͽ���q�%�L�JNgK3AV��FM�f:��a��ۑu�ej�Vt�+2��/'=�s���}��q�${�VJ9������nH�w��������؍�E� �%�1���Zr�DO�z����L�s���.����J�jμ��o6j&e!��s��M.��Gs��%PC��k���F;�@�s�j���t��� �6�Lgv썷�
w6�t�^+��]Powf������ �H�"@y;�{ ���f+p�X�b�@�n�b1i�J��S�5����̇=��~�(Гy�e��ݡ�%'{�M'G��36�����c���8-:�F��0&Ц2������
�{e��Ɉ]�0��+%Z�ڨ�v6�v�:6�i)c�C��]b�\�-�"��M����L�7%�/ݰ��$O�z�ך�1���0rS"u�u�z��[�#��O'�}��:�܋k�PI3��t�Εo0�kh�B�J�6��� ��_%�666*�Sw*	S� pl�W׋Q1ٺFH��nj �[J��ǂ�q��5�a��	N��*\�����5�Q�0p�y��}'7�r�Nt��zT]��6�Y�mv�wd*����5�3��pk��.d��i���1B�V����6Gc]Z�{s�g�X61��&ˣp��i�²��Ip��t(U�ER�D�++-Z2��^��9�ی�+��ȡ����\�.0�1F������Km�dE�����%�m�n�m�9�{8��vو�ƥ��*��Uţ)J���*���WT+.-E�6�[G%�F�*
4��k,�(�2���l�\b�YEU+[me�[m��Z+�G�(,���
�Rڠ�J%B���aVڱ\b�����0+U8k�U�+�శ����R*¶�T��kbm*���1�UlX�m�h������l!R�kYqf%��Q�j�p�Z�X���[D�Z�Uj�k(�-J%*�ËD+ch�km�[J��R�YJ�RYJ��Q�EK�
�pƅЫm���.%(�Ů-kcFQ�F"�j[J[R��F���QA.1L-�mW��~c���vx�u��]n#��6[Y�/=��Տn�s�U%�]iɶ�y� ��s��gs��i��m��7�97\ۃ�Ϊ(���]�z��L�9��3�t=�{q.@�9V��\�t�EN�S���xzR��7H��u��t��F�G[�[\>ԣi�s�0���:�(ƀ�lk��'T��ɇ�˼���;�)���g���F�2��NӚ^��������{e�-ݧ�ܠ��gڼ��uð���x���;ۜyD�Iݽ��7]��\�J���ᘨ�C����7���ў���)f���������=�j
s��M��ԡ��<N_�n����Q�)���<�0�j'G1�{!ɣy6��&�i�lRΔ\=<�n�Yȼ�8�ˊ�t���wg=��[]��<Z�l�O�g<�٘�;aNTv\�����kgA�F|�N�m�t�A�:�ui�9ֲ��9C,�֍�c��V�d�Ps�m�O<�U��i�Ѫ�=� �(�֠ݛ�nqU�p��:�$�����f;>5����i��7��m���la�����F5v�Y��q+�r�z�ܭ�8�e{{��ග�m���]\[6�+���;]�vݸ����;n(���=x"xd/&��]�ٚ�<�zХǐJ��sֲ�^ݨ�n�gԙ�%ݖ�Ȯ�|nvo]����܄{v��VM��!�W"��K�ʬ3���ʛn7������s�
-ӣZ�u�����]�)�l��0��<tVݧ'['n�v��:�5��k(��0s���6��>�k�7���en	{f�\�������x�c��������l��yz��x��n�}�,��F=�uŃ�ng�ͦ��1j�
�x�Ȋ�4lo]̻���6�vU{����&��y��{Y�ݞܽVn�-�y�cc��n��xp<޻=�l`݀ڷڳl����z�:��va4�q�ͭ�5k���6Pq��vҫ��ti���3��s*WnNդ�ˇ��-�\NC62l�襓���T��[�o���- �k�#���x^7��um�FLv *wkli!\��]��Fnuu����c�N|v��;v����V6G�[�a@wmqѲ����n 9��w1r٥9��&���v�O;s���7�9���=��:�w��ut�9��M]%�I��n�:��0,�̉�k���ט]�n:u��ntkA��Evy�GtV��C��< Wo����ݟ��Y�{{��b��� �/{uڰ@����N���㊟�t���ݻ�᫘@�*�}�oc� �ښ���FV�E�{�����n� �FN��T�	@��$�YsY�7/H��!�DQ,���z���|wk�S�>[���p˓�x�"W�wn���@$���تH��	��	2`�QJ�ԛޝ��Ev_T��� <ͷj� ��ت$×��{<�s�/Y<l�]�79=�Q13S5.Z)�J����^����[��|Gx^v]�� l�l�@x�Y1]2����Г�����z�%���׺�X��U0W5[�3̒�qs�5��}~�����v����^�����a����/?�מG�.]��iiu�e�$�Y��H9�1ĒfR��j���)�`�Ww7�MhᲵ��UOJM�p�>��,Αh$�v�՝O.称WKwYj�%yi��WKg�L�*q��ׅz�y���=�-��\e��tf\����$%��T�h������RXH��t��&I8M�� B��;['����|�;�/�@�x�R+�Ca��e(�AN�u���1�A%=t� m�#��m]ouFlP�;��ř�&�9 �M�@H51I�&7m�m��ʇ=~~��퀗���h 4��Q�;o��d]Sq�'�F��@7��p�0�$�N�X�b;A]ss�KÒ�}75莪ݔ�lW������MA�N��=��hy.;y5(�P��wa��~t�"jDd���D@�x��\S��ª�����^]� �Tq1�1.�\Nݨ��'<ӷ���Kv�n�h���q�Y�"�&c(���	 �a� � ��ڡ)$�J��j�Dn���_HN�NθF����[Q�%�5���Ys;'��▯�ǂE�mC�N8�u7Zb�z�K���V��ܐ���Qv�n�)�-?�QT�>l$��;S����WH�^�4���۸��FN�H���辛܋uC0ߒ�{��%�Ejnd��	c��>�dA�q���z�=�q.+
'}�� �;�:�Ȉ�7:[*�����
�����jp�$A�ό�>k��N�8ѭH��͵��y(ֹ5�D���~~�����jA�1K'������ ;o5���@,�Ζ�
�<�����w�� ��봬={H%q$��$���H8���A�������/��x �yy�v ���l���]����]{[�:�n)�eLULEL �6�.��ns� �^s:�+�&}�� w^uݐ ��Ή5��y�H0�4 ���ڽ��\du_",���}��� Kg���>��s��LV��-�Z"^]]�e횊,(l0��&1�fZ�ê��ԃԸ�Tx��nb�s/8�euOh"-��0�Ĕ�a�m�	��}��I��n���,�MD��A8��ة� y�v��T�C��]���v;�/�@�lm�#.w>�Y����vߝvD��س�:���[���t�rΰ8�]E��7O3a+����7��N���`~Ȭ��d@�M�j�DA�^: ��#}%g������m2�_;}-���Vj�jAA��r���ݶ�6r2<��h�=���FC�{ژ �Y9{-�����SA�\����S��)yH%q%Tʘ���V�T��tm��|󽽮���Gfi��&�8��$�.9y.���*}"�द�=�=�Չ3X�hDaݎ�A�	q������f'YjciY�Kbg��ID�,`�1���k~ >}�l�U�����D<�c��|y�` �|��u�_��|6��ڊ�	�{�4�<my�\S~7~�1>�9Դ�� о���K�����������&`�܎�ּd��~�D��W�V�-���ɦ6�q(�:���&�|p�|��6�K�'mu�-�s�������s�������[�l\m�u�ё��<�IԷe��y��qu�������\�p]vp��k�wd��.�n���|m6:wE{pq�v��8��՞vM/�\�z4�u��:�4w;��e,��M��1��0��Ÿ�muˡv���oo�|v��uP�q�9{ixu�T�捒�-Uq��U���P���q$�E�>��P��&��K^K$�C����슭��zf���6+ԊJ��K&�®M�a�\E@K=ϛ�0Av�?V=�e�מּ�� }��:h �������}�����ɴ�E�Y�I��D9d�m���#�s͂�SNh�x����� �/DD?����}9uJ⊩��h��A�fE~��=Q�������@��m�@8�aA�G����7��頌�=�􈊩���<����DDE������麳��S����D��m&@���/,��O��vR>��g����=�˰&�;Xc�vOYٍ;vT��s�,�6E��s�F�L"A�!� �yi~�P�D_vy��x��woK�����t��6�i�I8m�o�d�3��I��l$}T1��4��H�L��j6��0�;�Qt�ˌ&!�t���ÇB������'�⬾~��el�"lCݕ���i�ܽ�""���  �}^�{���>��uJ��ބ�%\���d�J%�S��JH���K� ��`�ƾwo A۞�C�"//��.򽘒J" �����v���e�ձ,V��ɇ� ���m e��+���G�7�s�#{y��I���
����h��A[�/8�F�y�ό<޻��ة��F ���@ :��" �/)�b#2e�ЬԸ0R��(e�v�{r���kQ�ϝ�.�nNm��i�7��������DULQ ���s /������t�
9���n�M2���E��Ez��K"Ʀ �Ѐh񇳒�H��C���V���޴� >���q�Ո�)Q��N������]�@AT�>m�|�$y��@p�h�/ZL,a�m������-�z����:�HNR{1����.�^��:q{�%��\4�YO����s8[����98 1��?�Yy?����Q��a�S��;�Q�dU��"���?Z���`�^:h����C�D�1�������򼘒JR(�,�ݶ�D۹�9��Aݷ+cm�<�����^z�D����ź�^n�4��P#
@���z��F�2*�to\m�Q�kr��9���Y;sna�ߜDjN��CMd�2�:%%�o&� ��w����;�a�^_�~2^ܴ� ��D3.}�0����@����� ��y����<��˚d�>���"�����a�*��:�'�Y�H� �f�Z\�P��I+��4ȁ�FxfS�w��^:`$����kj�nb���h"��'ѝZ�ٶ��>���|� [����$�W�̳��g���Ʃ��^U���T�㱵�Tt���9��B�Z,���#�F���2A�������-�8�*��f�;��y�����y�I�B��`6Ja��Q}�2p$�;��Ҷ0ުs<���C~�� ��i� ����V���}����^��D�ELv�w-덤�壋�]�g۔��-	�V;r�,�����$�P���Dl�:ߡ�����`��"������];��yw2�۶�� ��m��h��T���3EZ��y�,\j�i�k=~����l ��m�>��z"#��;�a�-��{6��*}�E�-EM�v����� �Y���P������@|��� ���i2}1�DT� #��ˊ�\.=��$Ky�T�D���$�Hr��q��̨ݮ�#����I'ϣl�rqذ:�#��$.��?������G_�ް�[m�	m�4�te�#>�R6�<�4��w 7��BV�Yܥg�(T��	�5�yM"f"qf�	�Q2n�����\�(�o�N����RK����R��-�gqvv��d�ږx��/o<;nt��c�u�c�x���Z.��˳wCc�ۿ�����ۍ�v���v.�X�E���qK������$`����R��v��w��mjr�I[��{&��["rb������VzG!��0�g8̶�xp��]l�ͺ�݋[rzb{��٢�-���<mk�'c�J�������͡ 5��>Nu��n],��i�G�����N
�k��܉�m�3P�.�%M �Q$��{z�������� y� *�)�'������$�Kr�Ф��p�C �L&�AQ���xgK^���� �>3����2���F#-?^���;L>R]�r�SS3��9h#�q�0y���ɣ�v^�am�4� ���t�F+=���"�b)IgW���]E�,�x�"5�?0��/0 ��w���W���D"=���'�s	$�	� �..v�ҐI%{�4Vv��6nt�$+?.xH��Ҵ�$��7{g�ժڟb�!���S>����kkj�6D�Qq�9���/J'kƢ�����>��L6-ލ+A$��$�d=H�9W�2I'ޝ�w��g��}�L�l���4\��Q��R��X������U���y�hS�N0��<�.͎���]�_A3��r�[ع�S_�E���Wx������\�u�pu]�d^ES��u���cl�Wd�3��J[��uI�����h��cv����#�s͂ 3'�Y^��uz�q��� v�6�I��拆�x�-TW�:�6��쾤�Xg�� �gv{� �ՑsV����{��d�=92I�}wF���H-�����",���?q��D�٭���I�n����2.r�[;t�������'?=e�t����.w\F���
+��;[�u1˺���IA`D-6"�hA� ��d g������}�� �>���q7^~��Փǅs�r��d�^]ݕB�X$�\AA5G͠�o���D+�S�������/ݛ���/����ZSRf7�Ok���с$�&%���u�� M�S A���O�iS��B��I��Wf��w�,y���	�L���U$��d�ܻ�>�&o�*w�S:[��7�nN��	�O�?E�!)��r��>�I@]^I}e_�N�|]p�/g���f���8n�&C;�꠼vJC2Ft�}Y�+�����M=mz�\��l�{��G*�J�K�o�ԍ�"��Sj�,N[�)v���o�q����Ax�;{s)���NtV�Cm��o��R�:rM�voX��{^jX/�"3��t��>^]�"׵K1����#sz�قi�7M��`�0��A��J�KO��q�x�ž����{��ʓɓ&�,��y(	�����ʺ�`{jmJ�A#ut��bj�=��p;� A�O�N�ܯG0<IeȥoU�����\��^����n-qK����G���#����5Mp���H_�6k� �LOL;�v�4�{�!K3x���yq���=᝹���ܮֺ�Փ����O�To�-�#w��I�l��L,�{�L�}��r	�e��"n�ƃ1�m�y
$��<�qJ�r�ܗ*'շ���u#V�*hlձz:+��#h���W��̈!�b�Ӌ6F�f\B�-�)�®�4���U]"t��7f�۠�m�\(�c�Z�W9E=�)L�޷��@��'C{s�;&,�����PY�zchk���p��/W<�5;.���	Jl�Z��9�V�rk�(��۫���y(�s���q{.9��e�sR]�Y����2i J>D+�)�ոn(�UkR���*[kU��[-�Rƃk[�UX�0�5�m)iQ��c�c�DIh����R�m�1�r�<;cnW�&�������*ڍF"�T�KU�+T�V����YD�+KX��0�Ҩ�����T�KUJ�--����[0�F��0*�LR�(�����&..*�me��0��qL[lZ���m�-TmD�e�5(�kKQKLZ���Z�Z�qqŴEQ�Q�[R�
V[��Km�e����,QQ-RV��T(��F����Ÿ+E�DT��Z[A�����0�kJ1A���J�#P���Tb�)`���K[[Kk�a��R��Z����j5,m
Z�m�E�aFPcl,cm*�ij��DT[FRűl�F�Acim�j�Z���b�W���A�TeQ*jЭ�����-*��T)��4U���V%�[KbZ���P�Z5�-�UU����DjTQU��-Uh�)mR�R�kZ֥-�kh��F��J�R�J�����л��j�"JW}) _�bHI�h�RD�����'=���sކ�l���q���֓UH�����lQvɎ,8i22�E%��Pt�K�q��T	�ӴR��g>��K-�l�����l����t�qO��V'rF�d���s���,]Q՗��F5�A^ɫ��q��L[�Ze(��yG�1An	bU�\�Pd@�;�0���?��ꨟF���}�$�I �:�(
J%���`�i�(l�kk�Bh�E�����0 s���:2���G���|c�+z���c�虸� 	����
:��b@ ���?�5��Q����|���^�IC�^S��v`�6�a&1o[����μ&���(�Ʃ�|�o)�H$�f�ۮ�w�oF���i����f&���m^D�-�n2!F��5�V5������,=:Ad��2�H���݃sjr���+xP<#�*�@����{e�QW�1*�R�!�D��D;������)䖀[9��x逾��wf.YO5�Џ���|��s��c��a�6p�A�� �՞:��u��k�[��f�lW���ݟ�t�n����
ܟD4y�����asK=�ND���g��e�L��,��M��6�i�"pKT��uѰ��������5L@��:` ���I� �
o��S �
�Sx{7�7��QEB6����� ���VA�O3������ ��x須���wi��",�IJ,����ػ�n�~��'���={�/@|��۸�H����[d�� h�򙄜��?]Tĩ��"e�F�uݫ i����Љ��1 I��D0��V@���&gut�n�������T�΂f��:�g�0�@�OA�ky���/x��V!�+sc�k
Κ�[�^\L���y0� ��	��aA1�Rz�K�h׃�k�˷6kz��6=*a�ĎWrdux'x�iKm�[{'m�[r[*Nu��w:[�R襎:�]q�wkͻu�/8ڌ2c��c�\�O#upqky�!ql�G�����"X�Ʊ��"��u�<� 8�\���G��x�[I�B��@��-خr+��]g�ܓ��˴6����燩���А��:u��i�-䶥���h�fx��;6��=�=��aܬ�����LĪ�AJ�2x��� ov�ldn�Q+bs09���w&�e�I ��Y��tS�F�a�h2S-L`KSܧBA�:{�S'��7�Q� ����@d�쿙����/_�s��@j��.��SELE* l���X|;v|�#�bü�ʚΈS\ɴ�Y��w�E$qn�U$"^�&!��(�..v����sDR{�;V ����������7�~�c�I����;Â"}T�]}^t�D���fkkHʾ=���>@%.�.�,t���>q��ɧ٭k��e8$�M�RNG���}��{Z"^�WQ�]E��K1�5\��߻����SH)TD��O���"4�����^S'%9Z��R(�
7���h�KcwbM��0!&J����uK��i�{��Q��ε���1tIޟG��u���}3������r��:���Ʃ���CyC���~Z���}��a��L7���>[�6�P�F���o�� ���>i���t�a�\��5��pKєɋ,&,��U�=�4^K��MJ@$Nd�_n����]x����i2�q���	b��l)�UE�����}~VMGu4 GVuy���x�3;����e��>}������M��ֵB*"!R(��\\�T�R[��V-[6:�z�x�-@#��� Xm�3;��X#�S�z�����$}�Iĵ��c�CíVNk�9fh�]u��F�)�#m����n��٪�����
2��>G^y�� �3�����{����6�2k�ZdDm�$���na&**)mW]ݤ�1랼ٕҽ�{r��Du㦀@|���V@����3=r�`�_�L��(AJ��cv��|��ݮ����lC)v�̬��
Ns!�ը�y��o5�����ޑy���%m"&/��;
����P"�P�6���e�L�fE�S�@�zbV̬thR�i~��q׎��7{m���DM�(UD9h4��.�}I�'w�l wwm�E������E��@��$��d�"̌16�%���[\��X �3��q�۶�.�n�%|�u����7{n�� 72�̅|�'d���Z�B��.h8$��7���\��=�c�s����M�^�� ��h��??�{��DB�QP(|-�k0|���ȁf�W��C�zos��8ح�~i �G�{j� :��A� [��2*�/�k����x���{�� >oom�� f�9&��WV�sV�۩�$����J�A*��{�]�� |�7s�`EgGoS2|��oڀ�_wm�V@��3s)��Gyi3B�����۬�*W�2`��w`�ٔ� �/=�~2em�Mzy���y��뎭l���q�2Dۣ��jT��bX�̲(�μ� �ol�6+wwSٻ/2�~������3�GEY:��r���f2b�I�\"�j��<����:6������y�u�m�A �}j� y��Zd���@�M��ߣ�#:���n�5��eH݂�N��uKrs�A�m$ ��G�MÂ��<{w��ٕ��Ge��H5�:��s>��-h�����@��l'i�C$��i�R��i�J��͡0�|���"w2��"�~�c��A(�Z��u�"$��SD���Es��|6��0��z�5j�w�dǭ����|ve4�.��y�*�a�R���	T��L����N:'5�~�������Q�x�� ;w��nZF�ԷF�AG;�T���@��"
���7_��Dv�k�'�0\�f�g�	 ��������ۻ&�u��$sU<���$��%���(�S�W-��l��fdS0\��F��l�eV�����c�@��׏����sN��Yyc����J�����..o��Oj2��Sb��W���r�i�j�u�7����.��8�aܦs���nZ�.�b\x��ƚ"�V^�����Pl��]�Y��5�&q�Jp�i9�f��x��r�\��&'���x�䆎#�\vn���pݎݓ	��g�;*m�w'm�1�hڶ�K��D��͎.�M���\���]�<�Z2��̜�Z窮��N�u��ڶ��g�����d�^#��]v��k3�����dCP���1Rd��Z���8ܠ��"m�a�Dnom݇z��,�"=�3�ds�^�Iˑgg��ĈD��=�z��5�k/�n�c��RI$��=�@|vomݐ �E�f��^��`��P��"*��T6���m�/7���7�~���[7 �6�$�om_�.��A7�8i�ꤟK�ƽ�7oI������/����f��ӊ�<��V���o���zb���P*)�{�X=h�wf���S�U~��:f+4��u�� F�v�a$k�RJ��9X���{DP��6�9��zV5���A�svܛ�	q-���p�AC���To�Bl��W�<�owk�`6�F�z����U[~h�E��ݫ;uND��-TRZ�r�R	7�F�@\�d��H����w �I��}*:����̻ZuHp�計���yr��B��O 9}��o��I�b:���&��٫!�ɦ��5��j'/�ȁ�ݷv m^����<�U)5��ߒ^�lHң̈́ȥSf�>���9�K#�2&#�=S���@��w���ͬѦ���Ha�f�C��<�Ĝ�r 	�|���6�F�Ge��鱗8;�s�TK�7.ť�^���N�P	>��$��y5K�F��[��fO�9��$�f��^�PI�ʒ]�u�N��uH�"��
B��-��wR����N��e5�q�n[���\�&���,���݇��JE>	�u݋H$Olfס� ����/_�'��q���n[$���5��7!@M��M�UEyݺ�^JsC�3^=�}���6�ܾʻ ��8���x��ŉ��<�=R�ߺ�l'�D��"�QC��mF���Hv�MR$���"N�OI�2�T�MM퉕���U'^[��묒j9<7����Z��Jz��o���7���9ؚ�Qny��72��Go8t���<�o  άѲ"����n<���apUPZ������̩�������,AFe��C����3S.�aĒ�}ʅ%��C���$0��k��������Yn�6���n�F� e��Dgvݫ)ld?
p�*�ʀ����I�0�0�B�>\Zv���94m�F[9m=�ۦٮ�_�[��ݿ�X�d��A]/��"m�` ��wm�p��^�_>���W��?� ��z�^vi�8��P1�mO]ش��Z�������y���-��y� Fv����5w��1�}3�ra�]�J*�DIU��;�� ����j��&�w[�dL�H�ܷ�D��yRM���ۻQ�Y�I��jb���(v�5�lG����d@�7���� H��ɔ���h��n;d�l�u/`m���X$C�w���a�&N���Dz�ۻ*���5<�Ll.o�0���%�9�X��u]��zw�̟Ft�l"�
������"qv�:"cgt�{5
�Jԑ��RM$��w]�$��7r$�z�7�j�Z!��b^.Ό��gq�<ܘsǜtqn��<�H�6̼���}��AE�HaÁ �
�L�I �f�U�%y$27r*�JvE3�8rM�[���@"�{n�9eF����	(�I��}[SH$j䷂���$!�<)�W��wiNn�E%�{�H�q⤻�.+�I�3m�[)@bK�.���  �ݺ�DFOG��l罿 }ݷD�I,ݷT���.la6YS��ی����Y�U���> �׮� �n��h���p��}��vN|�&��ڰ�z�$�*AP
i��mn5�|�y�D��!��o��p|`����ղ߽�2���o~y���	O�H@����$�I!!I@�$��	!I���$����$��IO�H@��B����$��HH@�p	!I@�$� �$���d��	'��$��HH@�`$�	'�H@�@$�	'�IO�1AY&SY��i ��Y�`P��3'� b&   �� �hh օh�� 4 ��� @      4  4)@��� E�:���()C�ƨ�����J��Q!A�b�(��
 $  �"��� 1P�R� �(���w|                   P        P       �  �       ���[s��[[j�]X׷^f�R���ꭱ� 	ӭ[s�ơ�6��Mn�
;m�� �� l���(.���C��@�   #*v2���8 J$�k���7\�eg3\�ٖtԩ�b� ]H)��m
ۜ}�W-��ҕS��A� �   <  �    r�i�}��=4/1G# �j�t�{��M6�F�U(�ق�i֬��N��m9���H�h�@D��  	��T��J�� ҩU��_s�X�:���^Z�6]:uJF� wv �ڝ���1��盥��J�6�V�U��[�   �  P    ��>�������yg@ ��֍ k�;� ��(� �`\�4(]`
{� ;� �G=��` 4�o �@ �� :o,��*��@(�  �@6  ���`  9� � 
 ͝#�
���wcB� �:<Zl( �=o :U��b�9���l��i�j麛�
 �  �        '��)˨�}g�Αj����^���8 ��v�Zӛ�Uh]s�Cm��d�8 ܵk;e�4��b�PQ @�   �;��+��Z�W u9�n]\�C�	�Knv.�-]c���� �Gmm���}�wG�:�wm�����+a��J��H   �        ި�����l��KR[��օ��ֶ�8 �9�ʕ��6����-���Sp \�Sk�x�=6טnB��ٟ   	��v�J��mu�F� ��4欫�)�U����Wz��ۀ�u���Z������kbۛ�Tx�~��R�  �)��J����d�b'�J�5S@  ���R�  �)���B   "ji��TSH���?���@��5�U�5������m�uO�$ Iq����	!K`! �����$��BB��$ I1 @$${����ڟ�?���[����k�����[�uo�,&���>{�#h�o�j����
YS&N��闏7�\
��{�V�un�E;nLI�b�v��Xl�	&�ŌH����sr�U����Kiމ���:�{�T�{�=;�i��:�ܰ��C�����n���*��x��NHfm���e�6KV��ڴ�P��J�����sw|�wZ2<hJ���,Me��ys�SM����jɷv�>G&�f�m��{"A#��Рf�ot+[�˦%MV���U�#r��z��
GF��3��yq)^T���`u��;:�V2�fb/�F-�����Cn��sp����iӦ� �L��`����	��ܷhy���R�[��#f-�k2V�$�L���sIӸka4����כ�5H�����^�n�P�f�آ��CkA�c]��l���U�{���L��D��`�I��7!��$̓+�eb���j�^E�-�M���v���V�V0K��m��6�i�9xM�)�w�4*l��nl�䬺"�� ���qTy�^�H+l��{��4��c�fKi�N�.]-7��A.��!X�,���c7���
�0ɩ��E��bJ�wA9���d#�ї��(�JjyS7U��H<��R�&nl�'�]�a��6�n�LH/EԻL��-n����Xʼ;���rc����n�ņ�"��(�2��eA�+]�Z�1���ʭ��K)ǫ9��wy�١��9{a���7.�efЕ{g4CI��cE�Yn�/ ��O^#8��mлj�_�X0����`u6���c+J"♣ۊ�,Y�
1������\���=���
�=��]�����\MZ-�#٦X�y`J�?m5j�9�"y<�ż
���(�r1�Jփ��4"h�`ۗB���!��Pf����.Aj�P!�$�j ����V�Z�a�L6i����b�H�#��lE�͛z��\:��2��:M��0$Mw!���ae�BJu.�=׈�@R�aO���n�8�l�)�a�6fM�!M��k�Hlڢ�DK�֫o����e˿�-�ҧyJ�`�x����5%����D����2��qZN�TX�c�fc�]ϝ]e��ې͗I�o�n]�{k'�xu�+,^��l�;q�M��3p�wn�2Z� i�^��l=�z̛�ji��S�(k�ݶn��vE�x��މ��öBOi��8�]�2�	��bIm���x�{OatV��hZ�]�j�����_m��j��A�<7��ycVD��(HHV�ޭ�����'ɋkB��֠����9�(��A���Ec-����^�6L5e�9*�^���$+n�b`֩F\6�Q��f�7 �ִ��Jk,� ;����TC��V��Zɔ>��n���dR�yW�h�Pg�M�\9�c������1M.�bBl�Z��Mѣ"�`�jb�m飄iM偬b���6L��ԩ�u#Xi�‍ē:���f�Lf=�v^L;e��t��*�%0�2����D̻��E�
�y�l�-�H�	�"�4܈�f�۠��5�X��)�ǖv�le�{�u���/cp��ٻ5�H[j6,X���A�E3��UI.-��z�l区i�Ӱ���ȡ����~�6�u[�����Q�vBC{�$��b�+A����&g�8qd�M�2�[$�U� ��H�ڙjfI��MՑH-�<
��֯^��ԣ3�tl��4̸j	6åC��Ƒ���Zŧ/or�� =*
K0U�x�X�3oI�KiI�v3qX�^<$��n�T�sI2�M!��`�2�agwI6�f]n��Y~�r�c��b8�?f�z�$
AQ]C[u���Y_��R��GJл�����s���ͺ�5��9R��m�]e�uB��V���6��-^To2P�$��in/��L �u鬕��!Uso,�*���*�n�m�e`:h�x5ܩ���v&��X��V��X����x� p.���2�,�[Ķ�n��M2���ږ�d�j�&�=>󄪤�u�[3&\�Z�-)� �m�[�(��ͭz3&�s)e4/S�	2,e��Q�-Kٖi���a�43B��r��j#�	��Ĵ�4��X���j�lϷ�X�7NHql����M�/f�f�1tk"۫�����Z�ؤi�rV��t���7m�Q�]��Z�=�-X�"#��5��4X�&��1ۍ��=/p�5��KљJ���[�s0++��ѥͻu{G�f�ӬO3#�i���T`۔>��@Q���U�^��Twl�iٛ�%؉��/a�+,KV�-!��Ю�o�+7d<j����a�j�moA�H�mZ�n�����`�C�z+�^i՝�
��f�?[�X����j�	'�� ��Ltf���e"�s͎�k+w	��c�d.�e5%*pV%im̧AK�[c�t��p�ѕ6�NT��@�[&��e�p捚2��V!���k��d/%j�mH�E�	�I��!��s�3z��r�P�BY&*�^U���5�mLūK*�iT�@h��f�7���1MiC8`�78
Ti��D�U�ə�{�dɖ"��r��L+Y��*�Ș� vXjY&޻Y+I��~�Sn��Ѕ��/$Ol��DƷVl�X����C�ulY+Ub�sn�a�j:VQ��nS:����a9�VV�o[���n�	��ʺ�C�8�r�Fk�˷.K���򛶲�&��5+�ѫjf����Swk)#��%
���ձA��M���E;e��b8FR:y�f�t�"�	��'�M
��^?�nI�%�l�k#f<����P���=�Kf�h��ݩ��%66�\Cr�$!j�!��NY7y�#f\�ѵS1N�E�جJ�"tmG���$����+��F������:�X[G�vv��#�*���u���X7)���6�M�:�0u����s4�3R�w�a�Up�cF�2(�Uh�J�;UD޻�`0��m�C���v-ǔP��R����˻�m�i�f6�HF�+r�51��V03�j�ˏI�e��֤����JKr�b�ߦ!X����甯�t.�ʕ�"�m:�Pu�&�ŏ4JMݤm�ڼQ���K4V�he˂k��
[)�j�3N��2�f�'@(c�ZOt�WV�j��E���T���'����� �ݝ�KA�R����ZVN�XZ2���8]by�J�ʸ6�SZ�f�ȥ�G�xY�ю��cb/�V��R�w�>i\;w4�lR[� �~���4�N���XrƺV�'�ԽH�`��Jˆ���b�&5��a�m$���aHܙ�+�0�ͻy ��L���'j��ɖ����D�!�X��h��ab��Ś��m�ĩ�)Մ�rƙN�
=�IH��h�sv%�Y9f�Ѫ���V�C�w�n<�-�Y�se��.�L7W��3Umc]ϓ�uJ�:`�b�2�����v6�Z�IЩށF���3>L
�X��ee�;�^*n)�x��YM	4� Ėm%Y5��tgۻ�ީ��{Sq�丑��ѭz��j��*CvK�T�Yv4d�5%yt�\3,��&[9�ڄ�6�������W�#�(#>���d���b7N=�ɪDfH��.�J]�Y�(�a5�\:�4Mf��ު�7���Vc��5�1o[ǎhʔj����Z	�6Eп��,y6��e�ǔ+mJP���`������K3SbfV����3֍b�!q{,ʵ��0(���m�p��"�`�vr.Vm��g$��\SV�a�t>{�]f�$t���d=�L �uV�OmnTYl����8"�	��K��Ձz��vH��,�p���r�6.&�x�V��(c_�e**�E<WM�fKaR�3n���oA����Q;�Й���.��
��=MM`�h=�˒-�T˧�Ub��Q�W�m�5��cҝ	�����70\��C6VA3Tyf��dMV���K[�d�ҍF�O,"��m�]5P4f�����=�6�t�a둛([]�{2	f�6� A�5���X�;a.bz�M����,_-��ʅ+�^^h�]Jy""�Y��e���SS�z�]e�oj�zԶ�Xbʪ�Sݘvj#4��u�BˋT�#��i�����m�u�����1����,�2M�+�w>uj�,L�,�GK�PUu�#?^�Rh֛�#�^P����T��/�\���v��&�B�-UU�.��e�hT��ۢ��NGiZ��4�0&��*�vE�n���yu�$Q���sh]f�[{�T��%�Z���.T��Vi��n�SAә��y�E�&
��˔è6��F�T3(�e	!k�+t�C�/>z�[72��� �x�:����:p��Od��1���z�R�3��C��f�+6�\��ӆ(M�7)����ɛr��h�{cߦ��Xk ��,fȖ��pѴ��X�K`"�u짋4K���֬zh����a]��*�6�ą��挚(-t��l
���R����+b�����܄��ф�&�і���iYV�S:��b!�ՂUZ���`��Q.Z7M��zԷ5���N��PM1��`���ku�oc:&P��`;�F㫫Ѷ�����r� Q�j�E��3AM�jS~���l*��n3*d��\�6���ɯv������a�$sNŻ3���EC6�9�y31je�+#	X1���(ެ���*�;�N�i۲���YRi�m��<&��%�n����Ż5���6�Ckh
�D�{s%G���mU��ˀI�����yeᕁϛ۔n�lX?�* ��7�'2iǨ�V�e�ǭP�M��d\�s�S�咥����4��u�.m�����-��̡�r��Ktƪ�[��5-*�/.���w�L_7"T,�N��T�̓)j@��ï2JW��W�84��r�i�4PLW�)	٢J X�"�o>vj��ٯv�Qnf�
'7^m��VՐf��V��6:���Uf�5́���d**ۓ0�-i&���lF�XB�c�ݢrn��l¢�N�T*nܕ+*(M�f*ׅI�e���5����#ن��{��W%=�uyv���6��
�P�ᨮ<j��j:��ܨQ�n�Ѕm������xq
�ٌQ�Y
ͳv������(Lե��
՘f3�w�`�N�VC"|FZ:N3ZD�a�љ�v�9{@��Щf��^�6��C�>q��Tgi�v&i͐�j��$%K�8jr޲��5�nKS[�c�F!R��m�!�DA��hD�f�i%����N���r�V��Z�ѵ�f��[A=�TE�6�;���\U���:6��u
ٛ4�qn=�j�j�$���el��s(5NڀX�TP̽���;}�k��Nܛq!;Is^e7�Bo)�a�Е�;�%f
�*�]]ڕW��+�`*��P5��w�(��h��#����p:��"���R	�v��"#5,ߔ�I��Ц�;���Ykv�����/͵�0�;�\8Ӳ�h�w@��4�i�5n��3*i���יv�Z�����^�3u�WkJ:^R��Җ�Y��2��=9�;�uw���u��*�A馨˥���=Ȧ�PIO	ُ1�ϲ�ì���Y,^J�� �kv�^9�.���W%�����
a���R����b��	Fh��%�-Y���wtnL�ndoC�D�ݫ9�E^뵙Zۧ���6�V��ժw��ćjksV��X�@e�,a˺���4c���v��,}q�m�J� V�B�u������iB#/�[Z�Wo/~N �l�v�͍ ^�B"@�F��E=�o�"��*jк;�θ��0BD)V�=���x�m�I���Sr���p%�偔KE�D�X@����b�u�hI��V���F�����i�4:�u]�d���ءm(�i��$ׇs�r����+q���.����m�w�bܣ��2���t���&��*H�~$�6~�[��zm*՜�_t�	���c.j2�0�ˡG`NJ�I7��۽ �����уD�(��ë~�51Pfa��t��1T[�8v;v�ͻ���3�k�S[sXgC��j�q�c�-�]�ᠶ�(k3���t���xtݶ��D�����u���ij�/�Z@�m��o��$ڬF�i^�ɚ鴅k����[�0-�܋2�s�ZE�R=�g,��͙�����/ۗvm,�h���;�"L�ТY�nJP�N��lǸ��A��RA�WY ����lń��p�Nr���ЌP�p=
�ꩫ4ɡ(;�U빵74�ǒ���6�o*��8��F��yq�h�R�+]�e��`�-(Z��C�t�ma�H$��Q^:��ʨ��To�fP�c��f\H�(�w��f���+-DyY-�դ�W�\ab���zR���)���f�6�5h��g5.=�Y1C�5��frcR��%Ҵ��]�M�4�f�j��X4�oL̵t�2�Im���n�s$��{�)�v6����c��+�w�V�ZV�y����5f�e;���b�G	u�E�ٿ���1��f�'��B(/[~��@��Y!���j�L��.��G�,���R M���[.�6�����ެT�Á�x,�SX�g׳Nf�ZLc����JZ�ZW�"���T��b�$�[���V��Uc>C"� ʊ�r�m�6-�4fF%�Z6S��"#�j`�A���˽[/F�NH#w�&�K9�=v��b:�'YH�=[�El�3��'>ۓsFd9��*��#�������$шE4�;����;�:�:�請�����˺�������ˮ�:�����룮�����������.��묺�λ���:.ꣻ���*�����:��㫣�Ϋ�Ϋ��.�����:�*��讋�;��*�ӻ�����:��������:��;�����븺���;����������ʪ�:���軺㨮�;������⻺:��.��.���캻��$ )� T�
bI	�@S%���]�wwguwu�E]Q��U�e�u���wvw]�w]ewwg]]�wE��ǹ!#�$ Iw?�9���3Y�x�Gf��gC��1�,�RԮ)Ͳ/t�Jvm2{k`���=�RB^ǹ�3:�B�q-���P�s��X����v�f�.��if��M��Ǘ��m�M�<U�W˂��`"�er��8��p9**�1��}�h&p+���Sb��׭����ʑZ�E��pZ��x#n��J lme�X�F�Z����:���uC[rV@R��#!�ƃ�-�	�+�*��[�B���f�W%W]܎n1^L�P^>o���
�e�eڃ^=�
�n����&�!`]t��\�ԫV��.�^ɬ�R0L�OT�ҽ��n�>���Ek�'-˵���]jˇ�������O0�X,K�R�/�cͨ�Q�8�y�r��6�r`({*��1��RԂ�����v��å;��;gsQ���w��g�N����cv�MW�U7<`�G��7���*ն+ѬW{[�Q��H�ޘa'4'�Ϙ�һ�Y3(��2�MX���n�|��f-X�ilJ��;�f�ۜ,��̶š��%+�|E�~y�"[м�e;�����,�Uu��S(�����eJ[}��U��zk/&�{1Q�j�e����u�����<�y��Dr��;H/���qVA��˒��T]Um�	f�3yL�8�.;k�|���=O&� �).Z�i�����e�;EJ��e;M�vt�ڏPO��r�\0�ie������
sĀ���Rm�j���,,JI���p��/8r��Inʫ�Wu��{�� S3/+���Ҙ�ʞ�C�T6�S�^�hլ�z`�X\T0:ȥ̷��d��Bzѿ��x&��@K���'pC����݋.���J�̮< �fҽ�X�MgV�Щ��9/x�n'��Z��a�J��T�T�,�q�t�G=��
i	��Rյ��"�V:V�á������њ�[8j�gb���GaQٗЋF���4�bB|*��E�3tK��J6�����>ݫ�:ض��"��G������h�fl}��7��j�=���	�
ԫ%�}J_n�nf0n����*�;�ĚZ�6����@��Vx9 Uv>:��ӛֲ�I��˓7l�c�M�Usu���JT��1/"	�=�����kE� 1�m�9#��=�9{x����F�n���J��-��m��&�U�o�c�3s��$g�#�s������w��.b�����&XHnu��ġ��#B\�FcTJSV^ߍܪҍ8Ǌ�\OV�A{g8
�x6�^U���L���1i�}��j���8Pɝ��x7�s
�ɖ��4���t�6��)a=E�A�/rtt�(5�B������f�m���1M�p�dx������U�)�O(G��tam=�3��(O}x��js���c�9�.e�'�hj�����a2���z�{�\v乔T���y�mNc0S㭭����M�˽؋����XEĒY������h�%��a
+��ژ�ܛ�k�Y��[��H�v�J�V6�&Ң=b�h{�M�
�X���~��
��N�nt���A\�����ܡ�u��C�w�3F-X�#�@�P�;]�Q�]�n�*�Pŋ�ԨΛv���&���15G�6�8��65��ɢ�V�����r�R�l4� e=�,;���I�Un�E1�Dj�+��s�e��91@�a��,}�{�`V�՗b&EL���n�t���m��ǈ��2�\�i{�x���2�P����|;k�I=}pnL'^�ܖv��v��U�p��̹n�ˋ6�
�V���Qm	�yj��Z���ۍ��J�9C��f�If���Ysk�I�ԵX�7w3�'y�9�Yf�LnoL[-F����<r��q2q� ݣ�8];��{]�;wY�C��6VE
㇭m�oF��c�� v��N	�4���8A��\(b��~�tQ[t�y˯��{���2ӻ�F�g&t�Ɖi�6�fK�7niu�v���%��)����+*�Ƒɺ5�wǫk%�Q⩡���*�إ��C��o);�Mg\ګ�^�^�{��q
ڗ �H�-�RU����7h6<=P����v�ݜ�=�Y�w.��h�vޤ�;U��#l^��@�b�.S>ƷEmůDC�0T	G�(�z�㲚���ؤd�۔(�D+��W-���9Ajy���/�2��nvo�*Os����5u.\�8%>�Y|�R��u�t-���L��	�,��0V��e�M2�LR;�(��7/yF-]�\b`�F��xؽ��b��[�YE�Tj��:�\�u-��n�(9��q�Tc~��qJΧu*�d��E,�]��¬Y�އ=�?��Ui���&�4d�[mC��-��c7����ƚJ��ge"*>�2�$�r�{~��)�W`�2gҶ��YoVRE�&��b�J���iZ�Q��v���^Կ,27�#N�����ځKܒe����,�*�������� ����I�H���.��Ѹ�����v.e����IK���P���k��<��Sl+�uY�כ#}�r67�uzl"�`����Ukn�ֿS��v�d��(�Q�#��r;�k2�X��vB��e�U��s�Qr�YԾ�t;��E�\L�ב���hڱC_%���ɍ�+�3�CeAYv��}�S[���3Pm�3K�,z�;���a�Q�Z�O�.�cOPHV����F5�]Z2���^v������G�F�j'����������'�چ��7]cga�.��b�X4*􇺨au��V�鋨;[ջN�?�#�v]=wy�T�%Jj�����k �����vr�'`�|sx����X9�P�M��D�T�e])AY�خ�Sd5���%��XsYXpoi2SX�Q����{0� ��+4�+߱�*(;�5��h��Qj�9�գyd�$���&��EWF�ƴ�*����CG���Kx2��ǽ�ey%`�1��H���",/,^�XL0B��ה`̔0�#�涒Y(�y��p�m�
��"���H�Tٗ�-Y󱹙x=x\�*
��
�D{3w�M��y���Ϝ��j�Ө�-�]f�G���6\�Γ�Y�0�	b�U�s�e�.�j�q�4�^�)�u��CK���f���JU(vZ����Yy�*.��X�u��)܌?�n?d��
��0i��˿nT�R�s��+s:�m�2�Da�5�>�휤;T��f]gm�	%��{6�-T��uI��jo���L�/4܏uY�.�c���}1�%hSo�ة�#Խ�37��,�s'INH��F,�p�[�_�J��b7�)ꩴ���mE�2�kbv���Xիu��%N�t���ql�ӗ�嗏N���,pk��cǫ�m�w)|7J�>]��w�0���׆}��֙ZY��)x�K�4F�iXG�-�V�z��{��(��q�9F�-�X��T��+��S3���͋��V	�G�|���T���ܹ�����'�/P�N�P�T�M�* �N6Xޙ��5�������E:,Tz�@!��=N;���x��Cj�"q��0j��2��E�ɻ�J��j}��f��Y�}5fBs� �E��\�-ࡉ�<���^�������}+�����V���7e:d���$n,b�9�9���9Ls/{�jX��G6�M���Tk*�#KMg4S����bC�F�n�5�Ǭ���1)j�����[J>C7t�j�k��w怽��{�1�A�����Bq!��g֓[3K�\���4�[$���G�T�ڻʔq�[�|�􇅉���*`�)���/sP�)�R�׵FL�����U��������#A�eKZ��i�(���-V��uc�k�K,��ᴅ�2�ݕRw+;5��\Z��O��B�`�G!XNɫ	�j_�+f�{b��&R5gv�s�׋ᕫFWb̰2A����p�lp��m�vMז�H�Lrӭ�{���D]���GNZ��'%ۨ�R��-[뒖f���K��B�i�thMc�5	�w�!��>��gҥƕN���Z�w�_l�U]�Gi53Wa���0��($e
����!�Z8�����W*�af��y3�ю�9�Fi��q]�'UL�y�$�z����M/[v���<.���U@��<�XD�so�t/����5g�8�f�ق`o��vn��tV�q����M���g��,:�_
��T���4��m��z��;�bt^�������I�8�鲬�+w30%x{lTy���˰���ѝ�u ,�}�j����|5cs�]�5-��x���$RK�߷�+;Y!>q�vOW�n<�]Fl��gq�[tPy(lc �[��o��=�Ǧ�]7�<��n�\:�v[�긞�1�~�M̫:�Q_z�Cl���4&��%�!���P�e�v΋��mք���_�us&t�4��w�Y[�ש	r6�HLD��#H闩$iva�V�%M{;x�kR�uY(��v���iq4v�/z�W+f�d��;����{]��q��\���yL������ǹys+53/�,%�7��[7X��YJ߲�T��z'۳^Р��1��&��)K�������|PW��ȼ֋�m�u2��hj�]�Q���Yx�*a����Zz�[N�.ֻ�j�)��K;;�#���"���G���[�ȋ��3y\,+z{����cm�Ue5l����G��ݬ�w=
3p4�]��������<�î��-�zu�T�7��]�����(�M����4��X��ڃ���ʝ쁲���c��7y�z�����xl�Z!�G;o:�n5��Ζ��1fm[���&���R�\��� �n5�l����|�Bh���v��\�]�9;��5;��!�X�u������Թm(r����d��Q���w}֜�:�'��2��lZڅ��͉:+':�MR�l�Y�g\���c�t7}l���7�j*K,�9CY���� z���J�����%�3Vi'op�t�8_1�C�d��P�,��v��������sB�N1�,n��nѕ�h���k��N�R��q�I�y�G�I�|�gj��m 4��k�y+]\�OU�T(`�Qz��@��k����O!W:�=Gp⻰Э�]�v��ewZܛ��p��>�����u�[}Xl����ܱ\��Ev.�Ԭ̉*��ؗ�w���p�>�7=��8pkL4��||���vEh�����R�bBp�5����*nn�
�|��10ȝ��e8V�qz���ʲ2��/賰��q��n(��(i�/�/�ta^��S���n���BM�dͻ΂.���_@��W�^-�W�{"�4�bQ���'F`HU��MR��*��M�.A��V1}�#��"�Qn�<���Y{0�)]w�k���nm�|a�uow�e<�m��̑���2��x����M�S�>�(��H&��8�Uء����D@k�ۻ���=k�3&ʲ��V�^��Bf���%�:s�MR�/��n�=.�f��jj�9
ʌǒ�{�V��I�5���7�8�.��B�$�]}qpV��b[�����I�ˤ��v%�T�3���*�;V
D�4-�z�e�#�L���ˡ]���.�ӈ�T�&�`��Uk0Cvp��N��N���m�=t�j�5T�l� �=� 	ax�h�Ɨ�FT������z�r./ �sr�&�$�����'���I��.ٽԺf��)��g��DR|:�h�_g�4���i���+��J 0Z�WM���[�5Y�ǈ�{s�RVS��E���;f�>L�]f3���o(P�z�F���͒G:�Jh�:j;;^��{[�a�\��cnf��5�
�/�-�}|�#��]0i�q��<{�:��}�o�.u6fW���AB��0���KX3+*)��N(gV��m
ȑ����"��Wa�I���YY���D7��Zlt���54m����"�ԧ,�s�k{�]�zf��L���B]-�[|L�٦47��J�o�m2i�盄�
ї��*���o���fd-8�r��Ӳt��v-���LH���tGg,�Hʖ�c����@�rNM�t�N��I�b��MNN�8v�%�Juȷ�1αj���Ү�g��ݔ��N�<�.��Mq֬tG�1�mf��ٍ��+�ض�9�hޤ��1�з5����9eC%�}z�Q������*�7]㔝��I���lQ��	N��;�k7���;�J�/6��+.���r^h��]���D���e�Y�����.�ʴ0���]�A�9�w]#�{]�r�u1-���>�;�n�,g�9!�s����{��2n�̐�#ۼ69���/x�NG.��pf]I�YS/��^"m�y-h4j�ն�ҧ����/]7iS/T�5T�Ns<Wp�l\X���j��Z�{�/�-j��N*�lms'E:И�g,�yJ\j����os���=5�h�*�٦6�GfC�9�8���n��yj�h����%� �0�ze����V�+�[����M^�9|����K���k ��ز� �M��5(���/#�9�����Z��)���}�$bq�vv�6'm3Lw]��W2�
�uĵ�� :��l�:ӓq�+�u�Rm�{]��'�ݚ;!�KMy���F�žN�ʙK`��ugP��Yg��i�YÝ��;o&&*Х¥�%���)nY�`�&>��f�w����6���h�ݻW�oM���%՞��d��P�p��(^�P��K�J+�=��of����g!�c2��;����
�0f�����o��3���̗]���_c;��k[��L�۸e��U�e&�m��b�lcnI�����Y�b�iE�?l�̲4�	�@?d���5��z���`�c���)�y2����U�l�+]&��<�ύQyxh�i�O�� �$�$�3s�E�2�,w�-l%	��ʥ��ۓi�]xK�۟)pu�n:0[s�}���+c�7�8�s:���6�X-�%�*�]ۡ�;�U:N�<�vPG%֠{;
�����G# ��B��B���:�Mr��B7<����A� ��y-���x�\mAm�6|�d�[b\v��N�M�ݲv�u	��W\km���q��*���Zq�i��g!α�C���9�8�M�m�+������8��S�:�XŰt�Pq�j�]��Usm>:��v9J��{�θ����+�wN{��\���2!���.'e7�;�N=cc�����۞ws�Lb;<u�e���l��&B�m���I�çs��xջtět�,���'
b�vq�����\-��n"��s�۷\�ݮ5m".�F{E0X��xc��hUثo����wc{�k�u��z�W\Za������.�I�\�7U��g��,��۪�곜�賚[r5�ק��-���C��n�q���붞,��:��t���s۰vy�`͝�N�ub�!��ՏkG�mvz9+��̎�N�k��u��GS��Z�<��ny6.s�ۗK�qˎP��z�j6��ր�Gm;���U��.{D��v�������n��g�rܓ�]�9�y�:����&�������v67���-v⃘Z��Q�{/$��e3��i�h���7!�\�5��]���N{m�]o���&����cs��6�b������Y���)k�m]��D����+A��7<�`b��z���t�;#��8�Z�qz�.�U;*�9��ӣu��<l��1��tf����xD�]ù6��ݣN�Ʒ;�n�7�89kn1��������[��؋�Gn�M�u�k�z��d��%�ݡ�B�0�Ɲn.�E��m��宖ˋ�f�^w�0���|�vqΞ��.nĚ��M�Sv��=�)lkv1��0`�ׅ���^�aj\X����sպsm���P���{Gb�;)���P{ul��������1˒G�	�!۳�z�1ҝF�tz�����N�g���;��봖`,������-0-������$�;)/A���G��]�#(�8�.Y��56^ў^.M�ڊ���
���6���u��ݗλE��#q hA��]De�S�o�:QW���s�(�v��ݫv���N-١�P��x�3�vx�A�vz�5�<�p�mp���W����lp	�����V�T��GC��lN���u�@J`彖헃d@�ٍזZ��]�r���v�"'$����/e�u<m�����85)C(A����qb��mi�y��gg�ݲ��'F�|���tY��:2G�&[�U�y��Rd�yw<A����η[l��su��{m�F;�kv��i$�w�v�X؞k���n�A�����x��663ۭ��	��6^]֐�s؜�s�<��s�!��N�C����食:-�g��C5d1�Q�^(e�)�{k]93�AW��vnIK'r-\�6��[Dv�g���
;a���;��^�v� �ױ˻p<�w=Z�\����8z�{��ݭj��cuƝ��7��c��<P�Z��s��zwd�[�se������'nؠy���:��u�v�uG6�z뛈ܭ	WC�Y��nx����>֎4rR�|t���ͧP��1F���k��8wzw$����zyUx�q��cVp�&�=���vn`��v,�;qڻP���4G�^�]<ɲ���C���a���^8���u��[�kn7(�B��Z7�Av��sr�l��޼m�R�v{Y��;!��K9��a.ׂ�y�s�����qz7��m횹�^ȝn��x䬇�絣k5��&;� -�{O��ۑ�m6]�ݮGnm���8w�]^s,�<u��2��m�۶gm:�zۣsP=��q�k�j]�ݵ��Q����}ɶ\I�dͭ���wVzα�F�rVN�Xm�m�g��������Ӷ��3�v{h-�˫u�^�p����%�v�<�Z�4��[nnti脼{n�'a]���e��`�5j��tF���am��lt㠶#�X:�8�1[��=o#6�l�%��n|����Q��&��R���.\����79��aqX�3��:�-�Ů����we+$�+3u��-yT
�M�\�1�v��z�'m&����3��ݺ�^͹�'0��<�E��ꣷ��.{�N�m��.A�j�(qI�vx�ns���n���ƥ�:�l��Ois�k����Y
Tz�v3Hm����;��	�5�k��L�n|����D�A���
g��t���DFv�yb���T���[ےx�Kϊ����`�X�q�X5K�U����v=X�xռ��W��𼎧�M�(b�S�Z�\mB�}�\�+�v^�G'D�l�Q<X�Xn�3�ؼ��[Mqu������\&z��2�O6�fS>U`:,��3��&��k�;]���s-���/b�)c���tk�B:^�4��s�'#n�ݧ+��v�)&��v圾ke�^��	�5�n���1�+/�e�ۇ���v���\��k�S���=���|���0c�iqծ�N��M�mm����t戽�.�:�{��v�a�u�5	�>9��m����ɳlc�Ɉ��gY�LT�-t�Kmj��#v��z==��ݸ�N�S;���/Q�������>ᜫ�^Z�l[]�+�8��shg�]{6Y^�60U��&�XfE�u��n�p[G]{;����uI^�:��ˊyvz	�N�'r�;��tƎݤlnNۇ�p$�q���nCm��"�ǰ�����x��S�ȼ묳�u.�� ���O=�p��f�vsȑ{)[JgD������ 9݋��ښ¸�����	��&,`�\+e7�ɺ�zB<�ݶ��+l�W�4���)+sQ͔�u��$��*�v{'D]�7���H��rB���!�En9���8�&�Y�oX����u��4w�s��.�7mg�5ϰ��+f�v5ڐ���p��0����u�ͮ�&콷�pnݠ�y����;�L���Gm�=pV��:��:�7##\�wr�$1���om��;�c����ݳb�T�]a�!.�l�qD���77�9��kbM�����K<��e�B:�]zU|���7j�/e��p�Ɯ4E�[V�7'^Lq;����1�p͹u���N�Җ��m$kv#yاv�;v0�cX�,�v�[<[��6��-�kyl��WL�2���q�7<m��PW�\3s��6|4m��'��R��o�m]���;�E���[Y�㶞u���Q��g�Rh�[�q>}�[��\�v���&F��x���޻%���/���n��6�Ísn�s�*�sZ��&�gvۉ��n� kN�g�";��G�o6S���S��p��;A�9װl�m�tMi��w6�z���Q��nq�i۬�wZ��uf���2����c����Z�ng.f�gI�sc�z��]��D��<G�lt; غ1۷��7oi�X�jլ��C�cl>�����kq�w��ӵu6���լC��# 郝�&�����ø�\W��Q��ظ����2��]Y�V�nL�m����{r�ѓ\�`8Od��z�wjq�J�0�q�n8�ݔx�����Ѯ�v:��+wJsB��,ZZܚ*�J��x�6��5n���W<�v�[��GW@���6�[����7:����'���� �H��k>��f����s��Y��>͹klu�*u�&-�8�M�LŁ�m���f۶������N�.����:���`�D㮸�֛�y+��u۳k�U|zE]�ٹ��{v8\�vo7�b�vx���dtQ��nm��!(���v�Ɍ�m����۝qQk�n���Jz�^xz7s
����cs�f������;���{g2	����7�b�
s�^w�C�+�n�����q��4J9z'���V�v�;���'���w(xN�+��\����l�:�s�]$�3��� ���݄mh��N93or���r�k�%�+m�s�'Gn�7sv��V���r"&�`,�Ɍ8��Ƣ9/<���g��Uu��"���;q��)�=!a��p78�����L�ʷ6��8�{�]aU6�wg\��ֱ��u��)79�KuO'i:]q�ݶ��9��ͦ�+;v�5q�Z�.�Z9���e�a���W�q>1�0k8�иRC��q������G\��E�Uu��b�s�v�Wrrݺ�Z�v#��v��G3b1׷0�AS�p��O>=z{s��u�#�����R9dsv��n ��M1Ϲ췃yJ4���{m�۬�`�y#���wm�gs/�=]O$��q�N�"b���q��N9�[]V���$*���F�qۃ�w8��\�<ۧV�+���q�x�c���V�s���ҽ9��Wl�s�mUѷ&|��lq���Ѯ�q�^<�#�n���,&�;d�uԧg�p����v�]��]���w:7ZM������kj.|^(ۗ�b]��&���A�\�n����A8�l����s��� 'n8^!�39��:�@6-;]=38�vqzsp�cvZ�9��]7F2�a��MLmҺIɋ��r���y�{��V�&��@G+"��ٞ�p����\[a�^�U��m�:���Sk��7u�phwau�W��5Ӹ'^�������q��u����md3�v5���ru��v�U�ݷ��R�p��i�N�'Y1�a]�n�&xՒ�JÓv�,�W`lyz�T�[����]�2�\g���<5��#�O.�ݎ
�a#m����;t�m���Ď�O=�v��[���)��Q��-���n�:zk�����M���k���c��[�Z�.z����WZ5	.�\f	����8�;��(��(��BI��9N �r��dGGt褜9s�DR��Pڤ��:����D��8�+��1��*!s�#�;��	Ӥm�n�"H��Q�9 ��qܒS�%�i��'r�	HV8$�Ӊ��SkN3��$8�,�C�����;�gh�q:�q8:p�$���ӗ N	��p���@�I�N �D�\䓤G9�9��%N�ȉH��8��$N�:��8�	8D��I�.	Ί�#��$PH8R����HN���Jr#��;kX�KWr\c֜T����
GN�����v�]���N73�NW����m.�>��y�۴�z%5��#��k��5����w.;v�g��'�Z(s�gJUÇ�[\�)�k\]R�"������	m�ƻ5h�=���>z��"��miDY���#��Z�wq.7q<�Þ�]�mI�i3�:玍�x�N��wȰq���m�9:��ۅ'���c\�5��ی�{��sύ77n�U/n
0ܼ{e�n-�ǵ�������G��u�=��'\m����]��K&{��J{�B�J<�n�x��b:�f�x��:�8Ą�=p��5�tq�"���:��v�f��I��ƞ��n�kH��g��mCmq ��\�i'͸����H��+{gv�$3ob���Ʋ�Wg#���%���@�Lmh=�;��`����' X���uS�2[��،b�6��קm�K��<�լ9�Ԃ�Y�4�m�덅��$]�qst�wu���u�r���C�t�}ax�`����tv�W�5ثa</v�g���)�f�is���i��&�z����z�vݶݥ;9&��6ѷ�U�\�η\EQ�0��l�&2s�Wج/.��{d�έ�m�&��r�+�+:	�6ػ��*�<��g�� �л�'q�yh��uݻ(6������u�LÖ�;�Ɯi��tM�Q�v����0F9[����Q�chzyѽY�Y ������7]�t�/����+�:�xɡ7c� :��/LpS�����`����:ч�7���T���z�����.iݻ��8�������{>;|����	i�v�|v�~O<�yL��ڹ�M�<jx����#�vܝ�m���"�/]@��õ�����U����t�x��!��y�3l+�;�iڭ:���N�oAڱS���\\ձ��E����m�!ص8���NMͺ�A��wk�����olki�U��'e�\k�n�����y��}�g�cgd�".l��
����g��;<�D��˞w��;{˼6~Xۡ�ۓ.���m��w8�vO&O8��g��ϕ���<&�xy�l�p�o/*��v컑���n�s�
��#ۓ�=��s� <�r�ȼ��w����N�xs܇���s�;cc����c��ga���L�9y�E0J'�^�����%�+m]�Y����e[XI%�v3�f-n���bS��?>��>*���D#tJvM6=��CknV_4׼�lP��u��u��	���Tb�t��KX�yb�U	+��o\7�M&���n����y��[X��&�G� ���|�|�n�.���vZUGjfc������|Bm�sV@$[���9��'�+��y�I������Q��s��Z����͏O}i�y�Ϩ
�we��(:����9�F��v�b�OP��g��T����ֻx�ۮo�+���]���vŅC�Z�D@k9��Ij֭R>�h�d�d񞾼�Oܹ��
^�6�:�^��{^����$�O���mg��+$���9����͏��X>n=WYH*��eb��E���M����<.��p.���T�����n����K^�	UX9����Vt�՘ֱl��G�WV������H'�� �˜߮�Uޥ��wa��o�E���GJʜ�����4�{��`
�03��~��Ӗ��T�s_	�צ��Q��P�)j��7��o"X��q��� I�Z�H$r󛤂<o]��Ů�kޔ��K�+:d����jfg���3>϶�74��U�X=���y�K��g����Z����j����B�+h����4D:U^�ìx#\s���y�u{G9m��Ԁ�ﯞQZ�t���%���w:`W��A|������3�hM7�9{�ϛ�;�G" �j�#�Z3M`$��R��mt'�.M�~���o�|��2�[���Y�v
�(���U�4��~$�S�	$�rἹ(���r�3�P݋r�k�k��WPCA�f�nx��g��lבc��`���[3k x:n����U��j�X1���������9����Z[��tN�:�}b-I��-���z�y�0�UmNd����97����%�sM�P�me�����:f�@��Il��z-&�;֡�Y���t>�sۺA�-�	M��Y��SZ�������إ6,f�F�q׹L'�5�=s�z��F�ls.�����0Q�wWtj�8q��?�a��jٴ1����g�n�	�[�Z/�7]����wI9�����\]ɜ#�'o{�I�o,��j`���yٖ��{59�����e���Ҩ=f��M|������EP����7�.G�����Z�i��wC���)$���-eL���kz<f���Ř����@ ����
}���&���A׹ObA� ���?����)�c<��N�Gb�s�)j]�W�4�֏ ;S��D�]�u+�vV���ʴ�V���pK���sI�ť͍F�v���>O�s�o���d3�]��@P󝊀�>�|���e����T�r� ��*TPF�5�k�r�cm��񹺳v�e�A�;,%b"pAcMQO��}�I]*��߰�4�M��w_1��f�]?AK��w��W֕��H����!��'�촴e��]�w���j�tD�"����{�|� ���`P �k^��#��.���F����u���D $�s� �s1�4�Ft��y��sb�=��i	����bo��e���Ӗ	o��U�k�3۵@}C���(��۠�O��ι�%y�Ȫ���Wh'��zf�r͂�J�]��]2k�����{ ��4M�V�pU@|�7�� }sJ�n�$�\/-֜��p�R.G��VY�S�$����gIT�O�#$�͉�)��׎����pH�7�U���
c��I����y��Q#{�/�t�8|�<]������\v�\�\�Z�<z�J����L�t�q�uv�cn{`;pe��8R'��6� �x�p�H�ی���,lZ:����՞mT�6�=�n<����[�����r/B��=q�鳸�מͳmG����t�\P��6 �r�6K�;��`�=�<�9��k��n�6^x�}t���{�v�*9��ݍFO�:.8����X�vzڝ�Q���X�TAx0���lX�(0֯����F�A��:�r}w1�y\Ϧ�}$ބ���w3��u��BJU$��e��'�oe���b��%ɛ�$�y��w�������i�=����t��X��C���,�(
�>�WW��gյ���H��������`�X|���v:�]Ӟ��}��f���m'�w�~�	�%�XH$ε5�݁�@�}��z�׻�dV�0���M��o�/�wi�o{.�!x�:���F��"�A�ε2�{0wM��wx
�U��u�7k�{[��㵮����%�0��k��g���wX��7�AI%D���/�5���o��7��I3��ό���ۘ|G�+웣O�&�iz--�E[���f?]��l]����:^�
��{.�� m�W`ؑ}f��y%�������d��5��E�wJDJ!i�;���ٵ��^�j�6ѕ�/�4���I :S�	���y_
@�U�@��-�Zy�'�*�$,3������`��'�_V�+��WB�7!?%)�0��v(p_��һ��Uv����o��C}� �G6,'�H=ء��_M�{�b�8��h�}�o��E�/N�:��-w�9���}�7ryq��"K7Yʧ�U�?|�,�u��|g�&�#;b£f���
�v�Y��s¡�i��'�a1yh�P��N[����[��1�g�:d+v�0�h�rk��̙�S(�I�ɺnZ��#��V�u^E��I�59�����ऒ�WIk��<49v��R�h��B�Y��'�A#����O��ɻ�:�lpN����?!`شn��ߔϨ�Os���o薽�9��0��9�~^�2�+�00��P�w��m{���:�5Q����Z�ң�v�B�;����g�cS�i{,c�ذ��w��C��(~�웠�pw[�drҨAU�����o�7�龋���*&|	��f�I#�ߕl��ˌa���M���υ/q�һ�n��o��Nn��(A�-�lBu�����|O��p�9�h�~Xjr��}����o�\�E

� M�:�j֛��:0s�d�vci@�)v��%�Ѿ�W'm(�Z��-�@����$��ߖb�nƳ=!f?fNi	���s��d+r�a��U�C��yt+"X|ϳ�~$�w�0��)��dov'��^TJ�+Յw��ٺA'��,'�~5m�틽�m�=� ��vv�'�ߖ H�0?Q�&�"�~��xz^3{*�?ɵ�/���H�W_�|H��N'�a5O�Λ�}<m�v;j��$o<�Uv�Wo��rp�]F����0����u���+,�q�R�v�'��*�x.�V,b��n��c=/kn���G*��Os&�$��2�pgT�I�G�n{4�Ex�%�> w������"��^`�`�Bv蘱��{vֻm���r��<��6���h�����ΩIm���.,�sZ�m���$v�!MV�Q�.�pp^뛤�����&���S��;h��������F�s��=���fd�	�N�� D�O(�J�К��/��Ѥh+���Uѕz�I��0Qpt&0=W�c`�}R��;S�#��U��Wdڰ���k���=���L��  ��m� ��&�҃��ߙ?*�ŀ��D"l��t�h)�LH�yۣ�}jWK�,�W��A%�T�+�=�7O'�W�	+M�{z2�e�#J�oN���ϕM2��˂��+/;xz�P��̖r��H�wQt�n,j�{�P��+�,�y[X�t�}��۵�����Dwv��K�v¯���7�kX�/k)�ݠ���,&�l���qΔ�����F�U|>7��۶�2�c���q�=��lv73����c����wO	e������v;6 �G+s�9;v�;p$y�]ogb�����n�܇%hm��a|�3S��ցs����+c�o2;a�u����n�"9mo\���%��Z����'�ѫs��g�g��*��ב�g�nۛI���ˁ����B�`��=��������X�U�_��v�����_@�˛���d{h��Ù��\o��t��!vlU���zn�B����� ����˛�(lt�E���vf�;�L�C��쌴^\A�roC�o��-< -���7u�e�ѽ|���d����b���L���$��w03S���Vm/k�$o\t�h�;���@����⟽�N1~�4���D�-u��n�[��Z�Z�����,�� ~���9U�6��5��� ^�/0π{��Y� rn��y���7��]�荰�l�l��"c�]�A��{;��9sfu<WE�#�2_�?ߗ������~��?��$��R :${na_�T�5k�U��i�Y���۫ �o7M�h*�\��F����f]@��֟:�v��q��=��w�C}�L�{����UrT���*2�gp�Y/��ٱUǳ�+�nYOJ�� w�f֖7wa�4�l�a�Y�@?w��6I�G�ܵd&?��=�״�-7�����d�G<�-�Ek������O A��sAQ$�N��X�+;yj��ׅU
��t�Y� zrn_,*ຫ�!h���6�u8n\�ݧ�	$��5H:$��,�@5G��^i��\�����dg��w�Z��s^�#��+��FMNZ�$�D�;�u7#Iޒ��9u}������&���k� �;��;3�=�**��'��~����;+ub�w>�,����m�tƭ'%��7=8���"
:�|-��:(K]���Y�F�s` ;74�|�/{/p�[\�:aa��.�I"\�d�r�p�D텀XL���n}��d��9�57~�T��I'��,��4H��b �ST��wN|ﺺ|I
��2�^f]�0�_[���	>��D�g�u�{š�Y���ܩm)�[��Y�Oa�q�� ��];I�Tʁ��f��r�:ڽGGW "�k��śy�&��/IC����W�R�{�,��w��N!Bj�X�R�,W�Kn�Uig��5�Ir���-=p�*�n��Ԣ��تkg�r�M�V�C97���m��{�*r��4�YWY�rD��]Jo}o�9Z��9�L�X��ͺٴ��sm�ij���P�o���LF�X|���e�Q��S5�S��ڇw�v���.���+�����Y��oփ�IVL��N%locۻՏv�_*;��`ε	��o��k���能&I�t��YyϺ��v]m=��'�#\�Y�ܵ*]�h�r�;���d�l�E"͍`��8��ܩӕL��r�n��P[N�ۇ��n�Ł��a�:-5�-c����фɏ6��}��哨o;��T�2�^?��h%妻�Y�2U�)��+�f�$��Wk�n(ÂC;n�V�ު�����ɽ�z*�
�Ņ�����S�!�z�o�����Ϗ	F�mMRվ�3f�5�a/)�@
����-��,���P�\�&����Ƀ�v���-�'�m�n颙�(�%�T��܅R��(���S�]R�o	qҠI�Q
S%e�.�d��N�=�V;�*��Q�{[y�T��i^f,U�t���0��j�4ɭq\�̾bw![���}���Q�O@�˭#�m�<gsY��G��u�#4���e&��DK������7��K�c�ޮ�O+O;e!'H\w��e�������=�se3rJy�*� $��(H�q	��HQs�����(�A�u�(�D�C�s�[i%B�"Q�(� �K�r�IJ8K�RB�
R\�������!�9B)����9gX��"�8r�
)B:,Μf��ܔ,�⸄:IK�%.$�vVƹ�
me�PH
rpe�v�QA���D�$��ݸ�NE'' ���&�J�I)�D�� 6�e�8\AI��㶭$�t��q8�9�ĜD�v��քwD��Yn(1�u�#���6��I�H�A)9NN'
R�IȎmhtHS�Q6�	D�2Ê�;������e��������hhm��Z^� |vrniA��v���
��VPV,U���D���.1�v�P���M} l��ǀ ;�y���<����{�*$�ǯmڲ�W�w�:B�-z��7t� �|״��&�}���{"��J��eIϱ?� �^Ř�&�=��>�f��{��������i�$X���k�\m/���,gx��vG�sv�n[ߧcB�ZZ�;�d���3�마 ��b��&��zu��O�n�#~���>�捊�U�ڋ1�*�2I�`�t��7��ەVMQ ��� v�*N�4Nf�r;F���{~���L�7�a5�}��dO��Sd�I���q���� "O�7������ױf|K�����D�t���&��擫V.n��˟` ���L��UUɯ#��5�xdӧP,�T3	�Ī��ϓy44��Ŵ���3f4��N��c���J��v��3��<5���&Q�ۃV:M��]!c9��u����z��qJ�.�#��qg� �ɸ3�T�׻�Βc�0�4I�ڕ  Tz�%�i�g���yVO�,U����Gb�����=�(�`mM�j0ι����@g{��w�U(�Z��f:dD�橲����rYTO,��:u��a�X� �k����5�|Ձ]�����&�&� �s��^{�sR_j��>罘� �sJAV��xX�����	i�N��F��7b�h��U)�D���,�D�L����Ǧ���<@ =�ō�?��Pt�p�,d�߮v���^�%7�s�|��K0 �ɸ7�>;���ek|˓�{5�Y�'��m����7q�;=95 �gn���3^���G���{`s�s_A� �{9sK1N9V6����]���e���Vf��m*�o�I[G]\��C�ˮ������%Hy�j[6��iV�{�����Y�H"�����-����x��򏜮��f��-��-���m�!ѫK��tZ��l�չ^E6Tǎ�\�y�8ywm�n�mp�磜�cm�O���v#�lO73�mɹ.×,��
ݲ��s8��|��&`�8:���b���z��v36#-�y�QmǡG�re�.r��\�ǰI�C����,����
8�.�����9�`��n|�u9��zuۊu!��[��`��'���rv��k�ul��*g;�ݮ�Gk����s}ŧ�Ijɪ$�'�z�d��k�b���ֻ��b�NM�%up^��T��^�$��ϖ {��J��y�uu�.��x��*�$���L�I^���2�w�-t�=��b��k���ɩɯ���o;s� T������H�� =���J ﳗ0����;S��[ec�ޙ{%n�TH}j�Y �k��0�$�O�yRFvw��1hTI��oר�slPT��$�A�o�>�@ ���,Xy��s��yb�*�w�� �d{� �j��NJj�
�^�#�s��v썰v9�=Z�G��[#�N��3�I��^j�}ͯw�߭������rj��Q=cd�j�������W���������Ā=����`��M���
�I���}T���K��p�����L�Y���i[��t�3Fײ�<Z���g���)��wK��ٔq˽G��,�����;���DLw� �|��@~���$/����u>�|'kn����^�w0l�W�0> p�5�=���L�d� #;�ىA�.�Z��z�]j�\�B��L�d/!�g1�<s� �kS��_ �5�<�>Y�kP�>
X+y{�{�k��G�����4q�B���rj��倀�����H��^�'�3̲@3�x0&�����Bǆ�&�j���⺘<��]��q�G<qڮ��&����$����#f4���u��K	,��A�ns2_Uw,�����I�,[�� �ۺ�k� �>�.�cj���[*������;���^zxwny�������=�\S$�&���XA�%��~�ͮrIs������nWhE*����ݝ�@ �;-}��~%�ͧ/ws2�L{OE�]=˙˸�k�V,'{n�fe\EP���mڅ�i�N*�fq��T��뺞���#^��D��s\b~��S�+�$�n��|�ssT>�S���v���VV�3N�{�]x�l�5�O ��D��U]ڦ�r�1�Q�%��J���/���XT"fɥF��;�vJ��ñ���m6�)�I$іvZ� �I=�|ݟ���m���u��ћ��筹�*Nl`wO�3n�ۯ!�R�%F���"9HR����nk�� �{s_P@ }��`o�Y��̱� u5&��H����c�Օ�K&bA���,�O�	o9������}xp��hD��Ϫ����7B�N�	m�!�a�>8�����HW��w&� g�w>���r�s�]�\��5O�D�~;ge� �;�C�Q�	
��RF�+Ӣ��!Sv!ٴ�Z��A��� s�=��@/s�ǓS�Iؽ^�PeI�������Lr\�l�ܛ��#�^XD;��6��;e�n/D�!�[�x�����cgu�!Y��~��z��q���� v����*�H������ �S�O���o�a��ۙ&�Z��N�F��=�S�� y�c�@�����ǬQiu�*�$�,ݬx��k�t@��7J�9�%��o� ��s�Z�%p��<��55F���wF �c	�0וnz[���I4g��j�换9d�U+��ċ}��X!�@��С�)�V}�9��~$׷Ɇ��8c_L��=˰����RVU,dt���Oh�=��y� ��}�fݯ;� Tf��Y��o�y�=+͎�m�DN��]6��ۚ�h������~��=`�x;(`啾%�P����V;��f웲r��\d�Ľ�/W>�y��=PY��0��m�=��ԝ]�MO{*mSn��$��օtB�z��m�Y��ez�ə����Bج�۴�GN,I�z���!_H���V�Vz���|�Z:^�"b�pj�����+5&�WU8ݭ3�\�;wTՊ�U8G����(M&ݱr��%��8G��9��v�{p��8�x��뤸�����nn4�뉓���FZ'�o����[��xݍrv6Z.<�qŽ[n�m{s�6ɝ�����;�6s�X�q�t�6m��#Ձ��O�[��8��o��g&�����ڳ͹��۷E�;�B`��8��kwt���m�kQgH��P٣v꧐�`�?�?����t�����^�ކ��5�0 zL۵�'�
�/��n�G~o� �&j^� ����k���UQ0�sS_P�1�� ����;?�g�Q ��I��u�����b��Gj�$,�W����������}F�Z=�7��oO��}���ǡ��S�S�-ER�r��A��h�t�?g���os�3 ���� ��;pw����ݝ�{f����6;���;8ã�y��%��?�9������	sW�3 ����;���A��p"��0pl�6_�Hꑢ�	6��s%Mk[�ܐ=�OCO��4W��K;�&�v�T�ۛ�{�I$�;r�Y �I��&Ğ���s����P6I��?��jɇ(o
�n�J�7�s/ l��qy�.ײ�fvՌ��F����N�gJ]Z:Rw;��LCj�.��G�ٛ�x�4M����z(�X��g-:���k\���%��x�e��� >���|}��0�}/)�oo�^�	>$��x]�VZ�����D������ 9�S/�����NM���>���P`���Ͻy����,�W�����fGǥfX�_��P ��� �>Լx��gjai��F 2���+�br�8�rRf �o�0ݗ����:͋am���k1TMS��� >�^�L�(���3�RȜت��ut#²����o��u?cR;�<��
&�G%��+��w���`��.�㳓&����3�ۧ� �y�<ϐ����ߟ�;�d��҃7�����v�k���q�s�pm�k\�����g ����<@ ��� @��k�׳m�o|޽75�<�~�ЩF섫Q�=x��I����2h�D���KA(p���QX.�Ũ�mH�R<,T�ehL�;�����}s���`��z*���̟J֡u��[����?!K���? ؑ��ۘ��=�_�X^�������uT\oS��뷽��s�<���Om%��l�M�k��h�l��xƛ^���"k���}��VWFYl�+3>-��0��[s=���s\��-A� � ׻�$�j����D�9
��^�g2/U���

I,�J�U���%l	n2��\e3����H�F�z��?}�?�e�,�����s�o���i�߹7M$a�Q��Q����G�� ]���D�K��������oݚ��|O^���o�k}�{��  \��Lo rn�A�;�պЈ�Ʋ�����k���q��w>�����z�7|u�]���}��l�w�^39��ʟ:4+`;!*ɉ��ս�=�a��\�9�1`�a��٤�}�����U��Z�V��VZ���B��vJR]��J��O^����r9�K^�s2H2���gq�� >k1Js5��sZᷙ��_��H3��U/�������z)����U��q��tlH3�v�^��r���ռɴK��)�I$�<vb� �H�>���gCw��0�������9��+uvyy��a�(7���Z��lV�m����9�GB>s�'�����\Vg�m�� ӻ�� ��wX���������vr�7� 3�T=UŰr�"��o�J��l�wt#4z��Aܮ��� ng,� {���@σ�ث�w�\>���;��sh�Kh"',��ٸMh�E؀��:������fu� ��r����k�0{��]t�X�<=��4����ü�w==�I2�$�I�ڼ�d��O��^.�\.����/6�B��	a���1[�9VFO��2I4L�^.��̋-�>��m�vi 7�r� bw�^3n��z-T�,��3�ۗ�Xu�k�M����f��5,T��d[�q;o��t����fS�Sۭ[��^�`�0:�=E#s�7*M�+Y�Gw/�*��)�4���'�:�{��t3fL��ں��J�~�����N]�тW�*��X���ޔk��w�Ԝ�!�k%�����f"7�[�鋶
�!s��Zf<���ͣ3��kѡ;�������ô,�u��̛dfl�a��|jS:��vD{��g&<n!�����0`���(>W��4�iE�5�NY9� W\f��}��ci�蹻"v5R�����V�|�7�W-'�)��h=�2Kxs���Z7�y3T!2=��/�&+�*ɵbCp�N�'�5���� ƜL�FغYE�Ǚ0��'V���¢^f����棻��}�QS�Z2�+K	��U���Ҋ̣�%�\�/4C[��uc��-m��z�s��|y"����)b�ܸ��܃O�L ���vc��!NP�)e#��e`$,/�w-�΋�H�#�Y��K&�x+��Uӻ޹�S)7�&'�l{u�B��V�>r	V�5v��5jWZ2=�9)d�:�g
�f���9��4wI�t���'L���*�E�B*�޺MIgY�6���-�q�N�X?i�vV�:��(`���V�k��� �g[f%ͼ�����	�	�ٺ強�Y����ãz�(�����ړ��o�[.W �Q���n�g��Zn��iΔn�u,`Wt����&���p�5b�� ��?��縀 �/�ؒP�
����ͻN$:H 8�q��P�:�8�9Y��:H)�ӑf�%N2�%��@��Î��;�M�BPrGNBaӊt�GS�'$�gi6,�98 �$ℓ�'(�N � �9�8�좈��GgZ�96���I�#���8�C��96�!�Pq�NQ�HE !!ӎGN�(RC�S��҇JH��r��9�Q$�
[hGH
Gr����Iߍؓ�Hmh$��%�"����8r r�$�G$� ���R䣁N)(��BS5.!$%^�Om��$qB:��:��u�Y9�Aq�s��9˒�������|��������.I��WOhG�\��o"P�����$Ѹ�;V��K�;^��ɲ��������qpa�[̹m&���NM��'�g�c�NՕ�xLn���Ϟ�=��݋�N���h)�������z��9q������z��u�l�;v�]���Slx6�>���^�h:�<�2�[�b�����k��P�F�㝵�97r�8��m�\ul���vxa�|����s�g�RA�w�Bm��M��.�S���8-�ٶH<H��z}V��U%���ݹ�f�΋���=��ݰ��(z�<;&"�t'�vܝz����gm���v�-�u׳�۷Gg��rk��룭]����k���8�n&�t�k�ykl��F��Mp��d3��;xd"����r�!<�� bos\k�6�k�94���(���Q�O��$�������Ƌ.[��>c��!�N^,u�Ŝ<ٺTѦz�&�S��@�vV�z��J6�L{p��";�E��@6I��\K�����s�,اl�6��j���d^ؔ�s��ZznLmݜ3��X,�]q.�;�&�&o��x��0�g�\��dm�of�=kSZ.;%�NݷK���z�X��:l{3 ��n�ͽ�1em��*�<�����r�^��u�[�]n�h�n
�p�t�;#����
X�����*DLeA�>�"!F)$�ƫn6{[;q�Q�;y���dtO<�gf����̸���u�U�!ͺ�/#��m��H��r�{n��������lVf���X�q��y�mE�xՎ��^��Z��ۭ�GYOZ&ū%�X�η�{GN�k�����Ƿ������.��1H];��M�0��[IS��nU��mxl�2kk�qi g�ݞ.۱;h�U��<=���g�q���ۑ�5+X��7g<p��Ƹ� �9�%��V{n�9�
=�;Һ�!��2�;�8C7=s��l�'tݗ�]v{q��<�wU�f��ai��^;n(�������/on�8q����ٹ���F��t���c��r��!۝���bp�l��F�K�cwCn�➯<q�10wm��a�>�\m�O<��7nH�r+=���975�g����w��������v��ҵ=�k���J[]������E(1��.��=��k��݉��v�ri�,q[d'�/<�u�&w�u����d�ܧcn�k��ݙ{[���n�%�OPݞ	��"��s��z�r��s�۪�6���ҹ*uZ���ă���_/c�I$�U������Z��r��+�4t�%��}��%��l���nT����\Vc�kƛ{�k�Ǚ�z=�+�SW&Q �^-�h�5����g4s�=/Uql$��[i3_o�O=鮙��6��{�M��5f�@�z�o�צb�fq��mE0σ�v�mV�v�6|�n��@ �;��Ā�3�p���{洧@${\��A��v�] WO���ϰ �9t�<���k=��%��<@$9�M7�ߌ���ɼ����eDV/��ʻ��u�Ө��<��m�׻���� ��j-=��"��B	�;���1K
9V��dو:$���$�}or��|�=Xp�9�]u ��3z^��%EV����r���ٮ4���zǷ���Q�꽢�Z�ٰ2�l�4�U�/�R����R�ªef��Ø]n�,VȜ��,��95��ܾ�>�V�U���fo�W�	w�����TUR���oj� ?����5�Ywy���s�}u�{�y�o4M�]%��٘Ys�O �gn��[�ʹ;�g<��� p�5��r�P^�4�����6�9�ؠ��w-�,2� x���d� ��Y�> ��ۖj<��n��|9�i�O{�[����
���*��7�^��~$�>���2ǎ�΍e_p[i��@|7�ң>��su�����/'�s~���"�}mN�Ȃ�j<�v�i��w*S�h�P��n�7���d �����i��\�T H;�v������=g�s%�v�2��U�©��b�4r���7s��Y�oU��S�LX6|ޓ;&� |{����3�٭o4r�v���@z^��J�]�)s2���>���۟`��T�{���-��i>Û��y<��F��RaU�FF�~C՛�ˏ/B]��V�F1�~n��2�R�!��T�C|���^-��_/��)�w7� ������k�1 >������X;3>,�z5�ź�E_[��� �k�  9��$����[�Ź��ۙt����`��5pE��M7�ɽ��L��;7x�mG� $�����]�����A��ʮ�O���֑�n0kg=��ۖwy�WCʏa��g Q�8�e�J�������⡖�*��<n����n` ����1�����q��#m��=�\�4ty�J�W��,;U�xt����Wp]M�&i'EUEo�������ǵ2�꽈�uQ��Fr���=��X ����곝��w5���f��s0�/=3�����U��ܹ���sӻ�ms��o+����w.`|�n^�f ��\��s��/�Y����z�u}�Y�v��'v�v��+!&�$M匉dq*X���n-�{�Nټ[���3�����}_}�W�l~$�ŷ��~��N(�NB�P�1f�1`|#�]��t;\gE���۞d�'���0 ƹu�.�J�C���^���`���\�u��=��oh�n86�r�R����*/8Ud��	�ͭ���k��RVs��ns2  �}٘ �Y���;�{�����9�{�ZϠπ[������.ʆZ�hoƻx�ܜ{y[/ܾ����kG>@|ܗ��� ��<tַ�����rf��Y8IT�W$z���&��HҷH��(M�5�N�������~�����Q��V5mV�^OTT3��{q�*�ꮧ�  ��@��jw>�^y�٬m�S\�Fv���ln]=��T E|�v��q���{�_f.�$іV��?;��;5��K���w�W�H��V��ma��S�:3�����}N�w�YO(z�?����+h��<��w��ڭ��p�em��PV�#F�>�� U���nR�)��Ӑp�kZ�j	�	�g�<���N�V��=����l��e넻v��8[ѣ���£��ks�I4��ȤG�1��˼��FM�l��I�=��g�w8�s������n���9�+��i�<�#�����z�Y28zK���鹠^s����x��y�������t��f:Ź��ێ�FuA���8��1T��s�猒����;��i����<�vn�ۈ�5�(X�cl���WߺO(�REk��s�fk�0> �k�= ��pxl[�<��Y�W^l��I�������Y��K\���C���>�|~юj��Z��Oj�U}UA��"p
�݊k�`׻�]�ӝ@|�.ʆZ����5��6|�N�� ��߼2-�ڝ�}�� J�XA�$���J�c��J�T$u\x���d�os�\�:�zY� >���vW�wX�L��U���ՠӣEXD�򕿉}��H���뭻مF���5�ԛԚ��j{2H�y阃�/�m����~Ec�B�R�ػ!�0z6^�u� ʏh(HĽ��z�v������҅���ܸ���P@$ާqd @z^zf�횪��!�#z��=�Nf(z�+c��-r�afk�O(��z;#�q�.���Zܨ3�uo�Q�;u9u>5���rvj���Swd��y���ب�I��ŵ�>��EWZƷ�������=A ��u}��?�o�L�:��t��d�XMz���%��P�k'�#`x����^~�J�9��|I�M�n��ޗ��� ����F�*L1�v{�ˋo�����;=�l����@ ���4(�7ܣ qQ\o�&�����@��uLxzs�3|riRw�z�nf������8^zi�@$z䏝�7ۭ�W��:�q�%F�|7aS��:Ȇ��;uZP�bvQ��lQ2X7�w�Όr��[*������ 6^zi� ����_%IF��K���Y�'כ����xH���[�1�G�[�&�s����i�gg��@/�5��k�_Q��^R�t�Z�Og���*U%P��33^�� ��f�N���)�ŷ��w�o���ݻ�}"ϏW�es��RW�G|��t��Q��[�x�6e��f+���7���'l�I����|�_g67�K����k�J�j�=�+[�R�3���w�W�k�㘀�<w{��@.ɮɤ ?{S�\��/>mԀ��ɘ�wO��#��2�a�g�� =���������?kM��I$BW��D��N�ܯ���f׫g�;X⬪;�Sc��1�'Y���z��jF�cVF�O���������cxs���H �k�J�� ��^���=n���c��-J$�$�+�V{�[��Q;*Ɂ���d�O��C���j�b�@��5�4 ��ThU{�w�0p����S����I���]-�˘d7����ާt`�t����T}}��D�$�Y[j�`���σ׎�QYc��;a�E��fb$�`��h�O�^� *$�\��*�+|���������z�l�=�
>A�J(��^.�	�Uъ�'{�r�0��*p�������1�j;Y�?}��}��?|9�G�곸V�+�:I��\�� >��f,yvs��;5���pI��H >7�v�o>��ă����ɷ�n���Dm��Sm����������}��q8���eBW[)$mZ|�Q���}G�h��X�l���9#� 3�������@vZ�˷�ܡ��'�� �h��c �Ք�8�S$zs�3���wOpz8KW`$�輘d��O^o��$�Kʷ~�$�(����YJ�y��B�"
�b�9q`|��, m)�5��`����M�禱 ��ds�+k���s>2s��osW��{}�_ā�l�h����� �:���v����1��	��� �5筪+-���l33]�� <ɥM{�<��������X� 95��� =d�6_�M�g��A�Q�
e���,Û��[�!]H��8�{7�=�B���݌��{tT������3֨׶����5d� I3�u�BW�L�=�fMXy��q�l/c��r�p!`�z˸�Y�s���b%q`����x8�88@��5۵ƍ�c�w]��]�`h�v<lr5�`V��p\rw-�w8�N��'oc��e��W3�ѶM�Ou|���=��Ů�j�>8�v^+���N�@*�W��ޝ�����hY��r�h<�Ć,��q��I��9�<����^�3���;J�j��!.;�s[��n{��v�K����;�5��c���w���kr�T�Noۺx�~�eP�&�'����s��G�]�Jk�x�y�0�#��J6X�a��;��� �u����罻��賸�I���uڬ ����44��=�~�Ӟ���T��{��g� Bu݅�&��}S��Ą��2I&�^x� zɤ�.�i9��P�K���m,ˡ~����wS�UD��V�&� Ի�D�I��c޴�k;�һ�~_]��zU�3�Wk�X�s>2[��ɢOĿt�L��g{�7�5&z�$Gomڲ	#�����;��*�Џ�8[�Yn#-����\j�����b.ݘ��cD���x�T���c��?uQYmv*:Sj�y` o�fM@@$��w�zl����i	Ds=i�I$�}n՞T���r�I5�'�7�d����[ߗ�*甼@�,%26ly�%�7
��X�"��������K.��S�+O��
��{�]\O��t���$"T�NVk}�g&{������s����==r ~�ټϠ�;�G�{��K{�M��WO��%,e4g�gf���o�y�h�D��=�qW�sj+�$�$��_X��vo1@Y{���L�*1�=7��v{V��j�_*$2��Y �I�{�2�8����zd�S�$�^_^�%�M':���IVL�'3 ��zb�]��O/y�&���@�� �g3�01f��T��AH)�NSZ�c��X�s����v:	����@��6�Ho{|#<�r�%���D��o�w�x���ә鍯s�U�>�69�jnv���L�>��q���b���7x�h2`��v��X��R���uV ߦ�b�s=5�wg�;��3/g5��57�Y�e��厒f���dl��X �.�zZ�uU|����YFt㇨�!oI3��h��C�۹��ut.��xJ���=:PX�*�J���iE����:�^�f�+f%�Z	���k9��[������/��ͳ���6w4�q�g�;W��^�s]���F��vЫ�>�\x�z�%���V��4�"O;��;�\q�=}1'�dcx톓��s���u��6y�g`�w�����ѡvբV�B g,x�����q:O]���bjc�gD;��Vig"�q�d�l�؛�d�?g9��e�:�÷�u�n�=�w�\\s]I���T�]�h;�V���k�V����g7Bf��Y�w�!�*r=���ޞbvi�Y���:]��w��I2���|z�շ�	�2�<���^���nhW�_M��vh�۰�Θ���[�sp�̓�hڌ ��߶�6&���c.�aFPp��ݧ�m�w[Id�����(�4ӷJ�r�)��ۓjJ͒�hɳ�@ML��e��r�W�p�]�Źp��qK��W��2o��E���@���r��z�bEc�7t+	�~�R9z��X�}v��z��P�]�>�)�6UNZV���_n@��ս��-���۩E�NGѪ�W z��"����J�nV,1��=�u�y��ꥬ1^²*%���)�{���ܫ����.�f����moe�a^��̮7Paxo��L@���qZ����#i���w���]��Svt�.�縸"p�4�A�Nk����vx�L��"e�o̻}㙗"4qP���U�V�*�F�ҐB�����}�_fs�'E��'h�(��'I8t%�m�!#�#��nIĎ9^�K4q"A.)�!ĉ˔�E�۱��Tr$�;�@�8�Nt&��q�qK��'�@����∐�D�]��D�@�wH\�S۲$��!�'JQ&ڊ)�J!9���I'#��3�#������H�D�N�ٜ�'	NA���Bs��%m��G9�XN�w ps��kr�
N(���Y�
!�X:;��ؒ�� ��S�]�nA��H�҉%:�
!=�"���]u}����1 ��o2A��k OZx�V�h2�;�����e��W�O��$��E�D�>�� x�˴Ǟ�1�k�32�w�����!J�7�ܯ��5D�ܵVI�Ѿ��\&8�< N�f` $zrn����,֯5�������=�Cp�F�fg��nf.	ݎ�ti��d'HI[��gs|D��V⒭O ��0lH6s;4��>���5�`��h�W,5��Mnf��N�fg�}�_R�U��˘��ri@�ō�oa��̇����� ӓsJ�����K�t��y����ˬ��z�$�٘6���% �ַ��ή��ȯ�,��z�m�I?_&��,��"�G%�f ��͜��Vz��:�/�a���~$�L;r� /����.'�l���������Qc�^�e[\�9 �Է����vB/9�L��,�|܎��A�{J�v��7S�j��}_U}���D���m�h$z���\Ǉ��dҁ��o���ywd����կn�m�3��s_A� �{���Ǯ���W��26�W@��˅��q�&���E�k؇���"�[�Tu�;���t��R���{��i�7��sP�h�]�".�o|��ٸ�`2C��s_@��"um�8��#~�r�*�s\~])���;�Μ���NEaI��O�A$�7����9�-o3���C��G	ce�FK�4�����7�G���u4��  �����/^=�d��Xܯ1�����&����4�@�����<@߹����S����稑�nZ��>T�4j�Y	kvLςs^�� �5�0�ML,	��Hv kmj�� {�q ~��^-�H���'�v.�ʺ���q��X�]�2��W>D*	X�l�z�a��<-�S���c��R���t��ge-[����݋���}�}�}�}��Ɖg�0r�cW���5��l]�ywl�q�F�&v�Y�b;��m����ۛt�U�������ܼ�"�qm�x�!����q>{n]ͦz�z�OM;l��y�#toE��l��hCq��Hr���*\�ʯj{l
w��q�c��K3���;g�#q��&���B�9Ц�U,@=��f���<���r���8���s�h'���a�q�x�Nn���ز��`ݝ�1��:/OYv�c�.S��n��ekn(9�z���ѫ`�PWo�F�r� �ϱ�h�v��l��oo�k��:���٠m��3�1��יִ$d�*x߽ۧ߰�z޵oe�2�  @{�� 2O�/�5Dͬ1}����ݙm�t�V���%Y1w���� &��uL�$�ӽ��oKQb'<�� {�v��sZ��ַ�;,��	ce���yfײ��w}���ֲ���y�:�@/r��ty� 	��u/io�R2R�D�0��u����j����ȻámZ�L?� ��o>��@����Xt[���U"��#��!M�|sm���/$��␔�!$�-A�	��.w�,h[Gd烷�s�ׯ^S$�I��V�Ԑ�m^��c��b�5ט�X�:5l�
�ĎY-���4J�4K��Ϫ�
��1p�x��s������z���O��^����myW�-��件��&<����fc;�YSn����;�K�������� ����0>?Mr� `^=��O��)��9�� ���N�R@^PA�{|�t� B�,I�}�}O}Y�n= �^^^�I$x���4�UT��A]�D�g�����av��a$��Щ 5-E`�&��Z1u����}j_mÓ�h�:��ZD�Fˬ2oVh {}˘{�o��=�����������;����;��Jf������dV1�dE��ҙ����^�rv4$�N��dPn�)�`�|^�JFKe"���ș�u��7�^�� }��6��ԛ~$��5�� ��l����EP��vMg��ܹ��;�Z-�ǇT�}��������D���a~${��4����w�ֵ�x
�b����ؠ���{,TI%��:d���(�D{�����9L(C��^��&�0��ܛ�b5LѴ��kr_^K�$�����^NT��U�QV���탏y����kF^7�$��fW}UUT���f�� ~�ܹ�j�����H�Z�<��/�-��sS��z� ��p�OZ}Y�3��g��mު���m�f��WB�b-y1w'3 �A�M�l����2!�B��I�� �ӓ0o ��=1�^S��斖��Sr��2E�۟.�����8��^�]�u�t�o<�39���%R�ܔl��'5f� ��[t� z���'I9}�]s��;�:���vf�(�[��`Kc�TU��In�߶����'lk���(�r�� 7ۘ` }�zf ��Z.�|צwvkVt�s������3z�f,�<kݘ� @��Z.�v�A�G�> ��31A��\�� �Z��ѫb,@�<=5�9̗�{仙���ޝŐ ��vf l=5�#��4��j��o��&�-�Հ�$I�F��	��p*���[ciߦ0��Oez��TJ��fG�RSܚ�����J����Nf(j��N�E���7����m�	0��TO���cF�E03�����?K]�`:$����_���{��Zb��m�ڬeI� �%>mE���r[�+�<�Í�j�r�\NK���?WB�b-}��Oh�l�;3  �����C���I��;��-�'j�����UW]���*�F�eǣv͠��w�E���$�������b�zs,�@�Q(�=3ղv�ޫO����ʧG�c���f|I��ϰ A�f�6�1n+&H@}k��$�~>�y`*]ҹ�a$��Z;&`z�f�}�����խ�<sޘ�> ��h {�y�ў}�췼X�I�-��O��:�8v+bb�����= �ŗ{�����;�v���,�nf  ������bG�z7Xk�xyz��f6bxf���j��dgV������g*�HNӘ�7p���7Lx�.������ssG^�a�y]Q�ӵ�{N-��/���� >������g���SK��1��m�ŝvH��wl]����v��������O3�F�/Iٓ��p��]��4�lF��m��c���.��;�$��^'���{vrv	9�)��ǎ�s�	O��-�5�	�h�&�ō�������5���uE0VI��۳��pq������\�v�2�I��'�;���$1yS���]���S��7k�v��T�{#��I����0�#�k��sp���
����{���$a�����]o�@4L;jՒI�MW�}�マ�S;�h�}�tU}Mb�T:��-в؁�^L�̢A7ɯ=sz���i��x��4�����3�1{�M�;u{�z���[��B���e�2Y������S �p|��7�۩� l==55��;�b��-�btv+,��Vb$׷5������R !�ٯ�| ���b��׻3.�n��[�����P9�s���;h왈9Of� ƹ�J]ﯼ����g��� ��m� �&�k�m�ײwn���cpX �m� ˣ)��W%��w�_��=���&��·�����i�k��]+�ڜW���ɐz@�x�V�$����ɾ�{y�,���Y ���e5{�N�Fkzx�N{&��;{��>�:����pj�4۳���]���;��ǹN?8��������Lm�A��bO�iU�nG���{m��oNu�>���z��Y��-�~�L|��?LĀ�����ޟ{8��2>�vp6���t,� v�S<g3)�M
�[d 4��U�z�z��v���Oo3�6Ͻ5�L�>���vJ�\RQ���7b�b���nk���f,��\��| ��Y��k�ٝ��_�?l�k�-�bt�T-�س&��M��wVp.���zo8�&���A�^��|��4�;�z�4���qw���۝�n)��sb=�`R���gN��9���k�*՟Ʀ�/��YhZ哟�Sى��+�Z�?~��V���5�՚�ѯ�ϨĀ[��f`+���+7`�xOT�D���Y��M���T���w�@>���� >=9�h��g-淹���Z��5u�j���P�E),zy���d������$6�ɮ�
C<�}�,p[�W˛%���4���k32�0��Ga��1����(���d#�x�׌a��HJ��j���k�B���rz��\����f�y����Yl@�{'5*}��|����
o�4� 7;��@ '�돆�����O��m�'o(z�%P�)(�s�������o>�s�9��}^����z��@؃��t@�f� k%�f���;���K̹����W�v�Y�9Z!�Xr�!gdE�v��0�@UX@�+D�ԖkXv��&ݒI3�ܧU��z��`��v�'"� �}����\۰�Yim%�����H������+���K�o)q��$��u�W� #���Ϡ����K{�tN�ӭ�wN��Z�nW�s��$�u��~%Τ,����� o�����>��5������ ��Z����NCE�r�n�s������t���0� �\��qv�,�췖<�7��«�DW2�wN���u���2kE�$^+�m���̬�D��\{�T��(�(cohb��}�s߀ٻ[�[�?�в؂�̙�g�z�$�L+[�z߯<�Ǿ���LȰ"I#g[D <s}h� ��;+j�����<F���Yͻc���[��1�y5�-�1�s�(�a��?/Ic�
J6^�3��A$����d�kַ��S���5�u=x�;�p��ff@]����Q7mb�$�zb�A����y��䶋��;sĀI�눿� ������";��W��\�t�\ҹ�a,���e�1��OU�Sh�]{!�=�J�hpֹ[xǻ��ٮzcx�<�En�j��^������p�ٿL|�{�1d>��zf  s-���Ŏ|ǽ���W��%u�^<G�=�>��|�[�5W��9s���g=1 e��n�4I�}�1>����)}y[�>�jMZ��4^9xs4i��U%Em���u��/#;S���du;E��"�����5-�k-*�������:�^�wwQ\AW�fǆ�aݷf��E_����H����6����k��e�ļ#K���[��QR�[��#k�*�b���-��Q}W���/4߱�k'�A~�t�$"�֜���nM�|w��Б5{P�S1[�k5�tr�T����|X����gy���-X�)F���9J�X��J�q���T]G3���R�U,2dsD\y!Ji0��b��و[��j"�r3�QK0L�R���xv�
�Nbp�S�	&���0G[\��ƭ(é�!7 �`�vOmf;t��5a^-5�ޙd����W��`���9�b=`꓆#�ٛ
P�T����~�V{���+mC��;5��E�x1D��:�u5^��"�D��[WPpkMg={y
tҮ�mWb�m�j\Xŝm�A�Î� ϮR�M��5��6�P/3��v�hc=x&��b�YXB����^��

9*��Fc��Y�]HI��b��7���F���'�i�)��fn�u��M��Ð���1�\�r�u!u�Z��uւ�iٻ�f�|�-6�K��+1d׆�ww5��5�p�}0<}2����M��)��]�@ɋ�X7'����9wũt�6(g�ڛ��>�%����~2:G�S�����rb��t05���fV`fHNc�T��Q��vR�U�oS�]���*���<�3n��^�hd�A�P~m��-[��yI����V�l��ޗt�G���;�rs�C�n$���
r��q9΂�E	��n��e�s�P���^Pp�Ķ�rslG{V@K�GHS�'D9'�GqG��ks� �;�
8���rI"H� (Gu怈8���K�8����7������q�#�����)-���S�)%�dD��"
r�ryjI��"/2���N���;"8�Aei�Ӥ)����܉�i's�Ap���(�A#�299fH�n�����,�rQI�p��e�B��m�^�<����M�y����6��qʒY��㎬�N&Y�i�@'It�����??{|�q��m�l��Y�J�]׭v�כo<�Wg�z-��I�%��<)O�:�X�9�Yg<�5q��֞�/[`�I�Ǫ��d�k>�����
�L&ﮃt]��}�|l����3��X2�۷����z���/%�v�[�����2m���X���v4^�1�=s�P�}���I�7Wa��m(��s�Ƕz��B`����]��$�e5��q�垆���s���<h�0��*��j����Z t��M�E�^��n����e�)�^y�C�u��as���ilZr�(i9�ay��/E�r��q�N�9� ����QX��[�e�ۧ�-<�����^���"�z6٧�kO3�q���tV穸6L����HK旱^��ǌ�rrey��[�M�7^�z�s�);6���^��O=���ݻs���%�>� 7�/����]������'�]�l��G���;��l]gt�q��=�����D=���+�ͽ���@<Ik{=�m�us�as���w�ݶ�|��}=�7l�a�� [��y샭v ]�u��8;r�n$�\�����{Hn#�&��.x��;1���ٚ�+�wk@k���x��:�f�V"�t�n;;c��z�cs�"���pt���;��.|n�Mknj��{x���T��C�Z�BB����:����n�n��Z�W�r�����۫�8�̹�g���u]������<F�.�K��l![����9�V�w@�c�\ܽ���U�ݳ�	�3��s�z��Q���7;�>�Md���-`���\]ö6�dѣ��:6� ��9��^�.�\)s�!��q���˷ko5)��-�kx�9�p��\�k�#r�����rW;<vC�2m�3;�\�y���-�tm�^x�ʹ�j{�k\��DE�vi�]�󝝌����/��]&N;R��v,�۶��	n;`���R�.�]�r�YYw=�6)�Nw8�I�+x�"�9�qӎ�z��g)9��;��۟tǮr1�ۅ(���Ǿ���������J(��䬽���k���컝�����gs�4y7\�ږ�qҚ���p�oEs��vx�����;���{qܺ����<8��l��Fwn��z� F�N����v8�.D�jy6V����r���\�ݱ�)勈�n�-T�qx�.x��:�����n��kV��k���Wf�Kb��3��\vl�7Zۅ�7U.�����T��:�A��9㭛wk��ve�� Z�T�C=�{��WB�bev�O�A��\� ����  G��W��=�}�c)}������zf|ޕ>u��j�l�ާ-�֧���k���32 ���zcxA�n�|@��Z��Eyu�WN�[��=���8	�h;b$��ϰ�f���7x�_�]�n^{�5��� %����H >rn��ҹ�a,�ҫang��vf�����Q��`:f�3 z�5� {ݛ�E�޼�7��o����<�En�j��^�{�tzH ��7�&`��ɽ�陹��߻2�(0�ٽg���\�ឋ��J�U$"����V����[Y�sO:6�;tg�V��J��j�n������#sN9�>>��;��o�L2P�+��e�[	(Q�ph�#ﻯ�a��3���sZ��{0��=��^�cX�a��aD22}9�[�SGJ�z�R�Wl�4��w�Q���t�i��1k��^�q��8z̯�<�t*�4خ�\ѻ`�sv=�c����1י�=�f�̏]m��Ύ�d̹�AC;e���b����t�|
��>��^�2g�z�X�j1F�L��f�b�6��Q�(�q��u��at>D
#� S0w?�����z�r�X�G��κ�F�Q&���-�3ɒ��ٱ���F��j0�=�}h��#��#G�s��n{.r�/}��S
h�#�{S�f��t��j1G��c0f��=�k]��v�vi6�ƶ�+s�_ޟ�=>�Ϻ�S0��Fd����
�H�Q�q�0�}���F0�T��a;7�^�m��z�U�9�����#23��n�0��a%��u�ɪ�֫F�+[�у�#�{Ya��b��1E(#G����Ʊ�={�{��W.��\b�:��/Z��i�L�����Q�8���֌a��F�F�̟��|���]Xd��t���T)���W�ۏ"l��_>�,� BDuW�+D"[�5�w�:�N�b��_�Q��(�,��i�al#Pj0�D�a{�}h��F�L�#Gfsצh�F�׷[�v�yl6�%��l���F*pj1G��澴c�L̿.ӛni�5�����=��/Mc�(�q�0����?W��p�z(˓�]T+a%
0�4F���֍����b���g=za�`�a�F�sF�F�kW��#�W�,�@G����-�R�2�&m�_�n4������Q�����SG�9����b�)��!"*a��]�?��^Õ�M	*h����g�R	���;+��2���5kE�7Y]��뇳�r}3�K�9���=gّl����t��#�#�#aLT�q���f�Q�B�IH����L1�Da����4kE����l6�L#3R��Lٿk�w�{����6��j0�F��ϵ�15�4��#0�������у�#Dq�b�zNe�b��/*z��������SQ�822��}h�����0�#�7Cz֪���Ō�F�ky���SX�a%
3�w,�l%]���W���4���9����1�f0�##�5����0Ʊ��5�#��gw�Z������)����[˙���'�u,�!1<zp�.'��\�GUd�(�3�G�m��i���=����ҩc�����y����Xc�b��1BPF�L�oL6�O�Q�db����4Ŧm����Ӣ;���G��`��_g����
�(�4}3��0���0�U���=h�!�i��3F{S�Y�m���D�ay����f�]�~��>k5�:�0���0���h����za���a��ڜ�4Ŧ�L)��w�=-[����њb�����9���rV��c3F�k���X�5�
b�}'2�l(V�Jah�#�������^g�)�C�20�#Q3��=za�`�a�F���9�i��[�=-�ލ�Z���0�F0�=��	�����2�[�b����߯L6�O�Q�21FOk\͚b�6���q�0��w�1T�?{����!��Mn���=M�*ڳa����a���|{��/��e;2c����\��vx��e��s%���7�\�_e>�|���g߄�~���(�B����^�c��0�{V?z�����MSu�[f0��K��1i�5��a�F���]�5�#ǿ�\�w9�{uÌ:�20��w�ޘcF'F�8�1S='r�1i�1S��b�5�߮ь�F(ǣ]$�f��pz�;��i{LK{[��L���GV��cC�a��y�=�L%F�����+cj��ɵ�Z����Z�v��<b�G�Jgd�Y��+a��84F����aL��`�q\��w~�ky�d~�?_����*0�A��1S;'��0�-�h��{�JYiT���Ko��J?���Im�b�PF/s�woϯ��m���=q�X�j1F�L�u���1i��Q�(�}�~�F0�P�
�
0�{6/o��}�u��{^"/��Dr����V�j�4�a����f�����F��j0�=߮�kF��aF�ͽn|�Ǿ�W���L)��S	G�;�i�e�F*pj1F���v���&﫴���M9+Z{1��SG��n�\����ϻ���鞌[aLT��
2�����V�Q�b������1�3F�aF�����1�h�_]٭<��gWXq��F����ig�i��zi���uUj�t��h���˰�x�1IA���k���O��W�/u��)������<������3$�Y�-3l�Q��aO�{�m�JaQP�	
G�|���L)��=(�w�x����<j���E_�B�хm�}�ˣ�e�UӮ�S41���[�XX�R����*�(��uF+����f�g��k|�-�Gxo�{�������*v���ݧ1�$�:C�x��p��]�]���� �p{;u��]��XD�<g��1�^6���s�r7��.��w���h����i�=<j���v-���s�d!|���Ǡ^�N�D�6�v�B-s�cA�@7S�=�[��;�Y!�u��Γ��{V�����͠�Wd�kGm�n�<�iˍp�q��N{V��U�7\��v:2.�%fM���4Qc�#�p�XfO+s�TB�*�ʣq���ʅ&����a�?0��K�f�[��#Pj0��w���da��4C��cF8�4kO�Կ_ݢ�/�s�8�L�5��b�
b��Q�8�{��ь#3�a�ʭ�ֵT�,l[g#F���5��(�N1Fz��k�_Ϛ�͜٩;�k�
�H(�8�G��m�3F�aF�o���m�MF��aW{��'���=ew�5�~ޕibkM(�S�~z�Iim�[+[�р����-a�PF)(#G���o��85�"db�hZ�}��޿aʿ��1�릂�O���n$ؚ�>^�=~X���C.��k��-,+;�F�>�=a?M��&C�w���B�q��S0���볩�aFF�F��;x���4c�#%��Y�-T;�^J��*q��j?gr��db��w��=�NMMV�b�`���{5�`<b�)��E(Q�I̳[�[	[�Myʕ�S�Za���0����ь)��F�aF�o���m�j0�TD��js,�i�y�������#N$Q�$x7n��\{	�!q��:�ȝu�h�,"�JEU���=�o�Ƈ�7���S�a��0��g��0�QJ�%h�|��lT��S2ֹ�4Ŧm21F�}߃�Ϙ��e�6Ä�F�L)���u�x�Gkg���N�Q&�+h��Lܚ��3�0��5F��f�O^h��H���V��#ڭo|w���|{��:��K��w�t��Qx����(_-x桵kװ䷓kp����}l��~_0�{�nѶ����0�#�'����a�T1��J?jsvi�at��CQ�<��O�ԛT�{�h�:��͘snV��ӧ�cb�
h�}˶�x��1FP�='wf��V�Ja#�~�e}��u���qaLTфa��o��a�cQ�j5F��������F���[�)--��\�����n4���޴�����T��~���b�J������l6�OQ�221FNk]��1i�db�)�������h��}}��z�g��
0�(Q�h�w��a���p�W���Z�QX�-��[M(׬�4�͌-�j5F�Q�~��]��0�7��<��J�+>4ÌT+�~�a��	���S	G5=�4Ų�#85��Q������>�w�}�Vg�?;wk��i�B��( ���8�b��t��]���矚��"nn�����{x}���D��x�*g���}���1F�q�0����ݚ�
�HP��Da����aL��a��s�j^�YY^�a��2g���k��j0�"dg�;�4�l��/B��h����U�oi�Gﳗh�
b�A�]|��/ۜu����4V��]�5�Qƣd�'u�of��ͦF(�q�5�߮ь2P�
�B�'y����|�f.r�� 罭4���Q�_�/r�J�&�+h��a����b�
kcQ�j!��?}߮���aF*`G�,~�3���~w�^v��3��)־�j��Y����ճB0�*��Q��������"Ol�/L�Bѧ�VE���ܫ�{�I�_����a���� c��ڞݚbں�NF(���w�c0db�����r�7Ѫ�M����w��~ϩ���mi�(��rw,�����GDa����aL��aF����������/�zqm����aFFsS�Y�l#DW�iֵ4���Zݰƌa��v�0�T���~��5�Qｷ��9�_*��Ze��Q���f��Ͳ1F�MA�ﳗh�(Q�Ja"�M{ݻa���<�o=�����yL�okQ��T�ڪq�ݑ���bg��Ρ�ۅ���eW�(�H5i��}<�N��!��^GFy�gu9��f�[�MF��a{;vcX�0�#�L)�����h�F��W=�M�Ԭ�r�q��ro,�]b��q���r���!��v���kEI4l�*f24{�����
b�;�;«0Q��;f��V�B�G#��v�aL��daF�=w��a�cQ�j5F�=����O��g53�V���J?���?*�P�B:McJ���G���a���J�	A>�{�&��8�b��������N�M�տ}��b�:����Q���3�h��S0����n0ǉ�0�~��y�:U�ϖ�[km(���,�9񜓜����jƣ�j0�~�.�kFdaFF������`��a��{S��L];��9��g~^��2�2]Zr��T�����{o�Vx;��|hmaC4�����B>�P�hN���Y}l�mi���>}���o����S�5�
��]�l�db����sE8��UjllX�dh���\k�(��Jg�;�5�B��[���i�=�豇\h�#�{���aL��b����}q�����5��L��ݚa�[�F���y��+�_���?���
���7U�k����V�ө&�T%�\��GO�������;U��V��Dֿ[4~as~�x�1BPF)(#Go\�q�k�����!�k�٦-3c#i��W1���V��[���v�a��T
a%#�}���h�#����p��j���Fc�jw�4Ͱ��5F�y��J����v���G;�ݘ�0�"daA��h���wcF'F�8�1E(��7f����5���;���i���g�h�>db��7�Τ�D5���6c3#G�y�6�Mc�Q�R���ݚڡ[�L)��0���J�9��G}/��y�1S
b��Fzｸ�ƣ�j0� ��jsvi��[�a͝4M��Tz��b�|4��}޴���Z�C���}i|0�,��_k�\x�1F�L)������Ŧm��5�Pq��۴c�33��੅t�FR5��\a�#����^u�޴B��+h��FL���͌-�j5F�j0�=��1�ao��+�����20�}��n0ƌa#�#�ONn�b��F*aLT��}�v��F(�<��w�?qC��\��}���9nP��N�
?V�dY��ܜT�قum�w�W�
��ҝ�4�i��X~��n�S�Nϸ�[Ds�d#n1X4J����ܜvzl�n��\��+{=m���q�!Sț���`v�1���{u�/t'�{������sR���|�����\W'U�1�9�P1ʓ���u�l��Q��;q���5܆��]�l���X�u��f��MҁӲ`�]3!�f�Bb�1�&�s�9��v�u�p�=�h�W([�z�bm�]�n��-�K�#.��5��٥����5�����F�Ui��I
1�\^�r�O��z��Ō��ѭ�>��<b�G��]�ݗ���T#��w����2���[^���o���0�*aM`�aA����e��ZiG��Kk��ZKUE�����n4G��]�����O�j�m������Y��G�]��b�֣d�"���e�i��Q8��>��v�a��F�L*�|��o�EN߻�G����6��#���?�A�F�)���1�f0����-�L)��F*aO�w.Ѷ�#�L)�ڳ=S��o��料ף�<��L)�)D���l[��T��b�)��˴m���2��NoN�N�M1�������Y�}�*�]��l\kI�(����Y{�[	(Q�q�0�9�F�S1�aF����ی1�`l�o^�{Y��ך�#�ɓ�Yl62�F��=��D�h��oi�Gﳗh�
b�A�(#G�׻q���(�]���;�q[Yё�2I�}�ح��Pq�5~�2���aB�#E�\��x���>��>��\׸E�ZO$vr�+�G�R�
�\F�v�O	�ƽ������ϛs|g�cv�9TG^g�FJ���f�m�jF�5G��]�5�#��1S
h�����щ���������t��a�*eW��[#t��j1G����h��L���|���T��U66,aM�o�G�~e� Z'A��о���]l�7zc�w}�:����ˈ>\u��Fg��V���?�x�xY����V[��-D��V�e��h׷Z-_ob���UK���H(�84F��e�6��20�#Pgw|���L)�j0�2��t��#��U�춗ZƔ)x����e��T[�im������aLT��h�kݸ�k�
b�A��3{������sb�bdb�)���?{�v�a��T�FR/��\a�T�|+Zu�Q�5�F�F|#%{;e�|�����M���m��F��a_�]��0�TFF���{q��1���SR�^�,�/C={��{�z��1S��b�5�̻F0�*fe���ޝ&���=��L)��׹q�ة���IB�U=�G�@�������w��k�����#��w�c
f#�#�g7~���5F��aA��~��i��5�(�\�}D?8s̹`)�t]s�vlj+=Ϟu�����C�W�:�SHt��wZA���*�P�B:OcJ���Q����`�b���RPF���v�Ʊ�0�*ddb��{|�lV͌�Q�����\+�e�ڧsH��}y3>@aP�
b�
Gۿv�b��ڿ:�F��S�%=��c1�d��,�+aLT��1＾�o8������ϓX�0�#�20�޹�6у�#0�(���Yl[�b��Q�%f>��.?}�ݣё�2{x�sUZ�H��5Scb�`��{��Ʊ�j1F�L���e�([a%
0�T���8ػ���#�ST��I��*n�}
|��Љ�6�rsS�(6�Pᗗ�	Z�4v�<�Y�zX��{hv����n�Մ>ͭ�K�V��or�P�B++�����1n��#
��α:t�A�6��v(��8�ZY��Mulwȥ��nѫ\��XL/�7hk�e�l\������}O묬��?e�Z*͹t���m;�C� ���
�wr���v��>�q֙��E&rCZ�o��*��_�cY������Y��6�qV6���.}�qtZ�[�;����l��Q7�(`�҇X�9Fl
�9y�hV�p�͢���=K�e�Mtq����М�Ov������w��%��&VNB�R��ڻ��ow�3E2ⷓ�<� M�	�sK�ڬ��p�l�Ʈ���]��x��T���ɑ�g��,�Zpe�*�1EC/r�׬���}Zwv֌�3#�8d�/\aS�M�@z�ݾf�k�ã�&-��Z>~Z&l�*�J��ܸ�ս�Lg2��-o<��5 � �"�i��P��-6#��ݳw��^��-^ZlL�Л)��3L6�ؓ1��k�|����]�ø%c�(.ɱ�!u�g����w��f&�n��h�ʕ��;�7�Nld�BE�`�>���fn2�}9���`���a"��x.Z1�8ࡻ�X32o����^#|��?jC%���/yԬ�l���;9Á�U̎���3{m��������s-�P��kb򜖶4�p-�����w�f@3b�]����}___))[YEó$��﷕�7�.�:(�s�tBNA	��).r��t�$	��
6��M��d�q�;"@��۱#ls�p�cE�IeiHHt�m�-t�,$��.�݉�;4Z��΂�΅��t��C��)f��Jmڌ��mn�(q"Y�O2���7�̈k����w��ݝV�7k3gvYM���vۛua�[jA��a`��;lY�sZCk'L�v���jf;�Y�����RպkqVa�K76�:�Z�H�$��$-�K3�N+9)�,v�m����'���͹�ݶ���[V[(��J��m�e"ve'����M&n�$����E�~o��������aF�3��v�k�#Q��1S*��Yl6Ͱ�Z�����%%����Ko�Q￷�%<��n���9��b��Jѿk;q�X��Q�1S+��lZf��Pq�5}���p�sӸ=���\�aYB�$T�]�.0ǀ�G��x�֪��=5��F*evo�[80���SQ��?w�vcX�0��w�W�?w����[&F�����у�#DN0�P�O��e�l��L)��S�=�h�1��2�}߫/�+S9��e�˟j�v���k����L��ɶ8�㴥��%X�Y�9�?WX��2X�/5��;�s�m���Q��(��o�^�V�Jah�#�y��ь)���d��{z�h�y���2����5�#���Yl6��zæ��5�G���h�q�~�ܻ0�RPF)㝯�p�>�xgC2��t�k��F(����͖Ŧm��5�
~��aLT°(Q�λ�vf�*�F�컦&��8���=HV�QSES�-�3FL�e�Ŧ��Q�jF�=�fc��#�F��k{ϱfNkݦh�#0�)(����Ų�#85�
}��f&F(�������*��G��LX�L��߮���\�p靲�����q�0��]�z��
�HP��h�#���h�
f#�L��~��"*��&z��67uP����-瓣[w�'�ŷ�f����s,Z�n�9���g\T�k:��omhҍ�a^ݮ!+�o�h������� �ɹ��l62�F����_��M9�h�kv�1��;�a���"PF)(#G��ۦb��q��7�+u�,ddb��z��[������Q����˴c�(��JGw���<Da-�|�{=5}�{����5�� '-�T�B����ٵ=��۲�;��ֶ�ζ[H�Tv��U��(����l�al#Q��5�#��˳��aF��SGy��h�F����٭�
bܢz{�[��#0�*q���e�1�1S3/ݪ7��F��N��ٌT=��.���(�q�0�ǾW>�vk��T��-�L)��S��G3�����2&�j3����5�Q�b��Wod���ٞ���Ã-�h�!�?�DִT����b�����px�1S
b�PF����Ǎcq��S1ɮ�{����o�ΖŦu��5�Q��|��v�a��T�F���z��S
~��HV�U9�)�-����'>���>o{�u��r}����#Q��?�~�15�#&F��SD�o;����4c�#R�露ئ�>=��{�w�t-��Z�Q������1���o�j�P��u�Odb�c#E����aLT��靲��V�fs�w�(ԝ��?
�i��S��>�ь)��F��SQ���0Ʊ��5Q�aFOL��c-�h�G��3ῦ��Sݖz��{��d�7j��č\��E�Ϣ�J���S<wK�x�~�2�ON;��(`�~�}C� �߭��϶wn��������F��m+�o7v�c��v[�r�x���W7T��b��6�kO%�s�l8���']������s�<��=�ݶ�g��!]v���˵�\����;u۝gk��pN����q�v�A̯5��7��s���:�m�]�3���Z�>'�qu��.�u�ݴm��6�ݜ7Q���Y���^��s��ݻt�{gv�Ϋ����e��m�\����6�7L�w�:Wj�Ӡ���zx�)I\��[��K�����y�a�F*aLQJ��k;q�k��F(���^��-�L��������s�b�Q����h��
0�P�	)��n0Ǎ�w�a�SZ�z5&�գl6�L�M��g[��#U���~���}��
~�}vu5�#20� ��4E�_��a��F*aLT���YlZaLT���w4������c<��2�ꭽS�I�Q��{1�������m����
b�W�;e�l$�F��S�4�n����.^�Z�����taFA�a>���k��j0�T���Yl6֚Q����O+)Kj��fm��n0����a���=sStݹ�0����RPF��_v��S���S2N�=�ش���1F�8��e�1���v��ש��+�(�4_5�\a��Da]���^�+Z%CR�[f&�'>�ٴ��F*aMF����aL'7�l͑����4}����a�8�1S
b��vgl�-�A����j>��v�aLTǫ��ܺ��z��~;��&�W��1�eM��a_k��y�7n��;��]\�C�֕ͷ�� �k_�k�W���^1F��Q�1S+�=e�[	(Q�b����ь)�0��Ng�]�7=���q���;�"���a��a��ٞ��m��4CZ��}��Z&���[�щ��=˴m�1`Jź�;>��J����ލp�[��I�!�܊��w�5����f�����xX����h�����bG�7f�q�|���ɋ̻�ܔ�\x�mί����g���~��85�##d'5��lZf��Q�(�}���	B�*P�	[���w�+��k�������J=b�\V["uк�cK�ezo�[8�[�j0�A��?w�v���20�##���w�n�OΪ{��1��0�q�b�W�r�bں�N5��G�{.ь���2k;�[z��&��Zӛ1�3=��n59Ϸ�};�gXS0��Z���Ŧ��G#�g}��1�3�2&�j3���q�5�jۿG����L#Z�#�ɓ~��le��)ɏ��e,��:�ʹ��m8ҏ�s�������QJ��5��<�(��o=Y\���5Ŧ(φF(��gl�-3c#aLT�~����aB�$)���1�h�#����_��.h�UmdcJ�H�Q�Z�d�:M��=`��
��TeP-��n6�}��謈�B-HW�l>g�ɓ�Yl�a��1S
s�v`�0�##�20�ܿ���1���w��u�g]}��l�}���L[.�1S�Q�0��{.Ѷ`������:���+#ٌ���5��5�g�OwR���9��I|�YB���S�Da}��ь)��0���a��/�\a�T���0�MS��oT��=ŏ�!@G�kߒvE�VU�%+� m�as��F�S0�*aM�_n�Z�(����2��쮎���X�X˷�s�(�\�3c�}ۣ��b�-���֎M}K�s+vYT;?N��z���e��^:��h^���LY��I���i�L����1F�q绗h�JaLT¡H�>߮�c0��+��m�7Qm�-�����k�^�G�e�3�ߛ�������G�g�Ѷ�F��SG�����1���SR�jg,�/U#Ϧ�]�ς1S�j1G����h�`�k���}:7d����,k���߽|�k��Q�(�����5���ޫ�]|m�ްX���?kyv���paFF�j�~߮�cX��#Q��0�����Y�e��{����׿u�Y�|�P�&}c%��xp]�x<1���t&�l�P��P������o�M+=b��aMq�~��v�0�QJ�%h�>��<�(�Q�2�Q�=�g6i�L)���W��}xl�Ok>��Mm8���v�a��T(Q�h�>��0�0���흆�:�r��
�-�3Ff����6�i�j&��٣�k�=���<���1�aA��aF��Ϸ��h����S%�k�i�m�����#�n��A�uo�q7���21F{1�oN�A�=+#ى��{���x���(�)B���v�l(Za��8�G�u�׹>+��ֻvk=�#S8�0��#�g���t�ƣ��#��k5�4�i�a���'+UIYep�Zic_!뿹��W̦v���s���%b��4]���x�1G�Q�21F}3]�LQ�db�G�
}��a@�{�v6wX ��v#�Q��&ͧ��Ĝ��'T̷�̓9��Fc�_�Y[��?C�j;���Z"��\��c�7�7��||�ҧR�.0��Q��#/��t�oo�Q�b��ݶ8�E�.|��ƾ�z�3���F*aMF���f��÷߽(��M�0��F�{/.�m��#Dq�b�����b٪�NF(�5y��1��b��y���>jj�����\(�2�1����Un��ǳ��؉����:
�_����S�w��� YF�kZ��L�#G���t�<b�)��BP�>��٭�-0��Fƈ�>�٤m�ى�a[�E��d�}���6�m��]0�X�a�Q�aFsY�ڭ,MV�(�L����W6��8�?_��6�lXJř�i��}��s�=��>&��8��ddb���_6i�3c#aLT���6�2�T�F
��ͪ����}r�t�6��O��5Q�Ӓ=HV�l[S7���#J���5M�w�i��)���SA��_��;�����Z�0�GD��a��M��i�z��T�Q�85���1��(ɿe>f�h�r�l�X/z߮5��j�����}���c��8�E(Q������(�4UJ�z6�$�k�?x�&�^��\g��6���M}	����J�,	f��׻��1�O��g<�R�A]ؘU����D�=��A$מ{�&�/�Z��8Z�Y~�7r�:Qn����c�.:�L�~=6��W��3��Wa��fZ��wTo�'L��9�F�(��!vs �;
-�1���8��T^�����Ն�q�l�۶㈵u��3kvlZ���rz�s��{oK�F3���鮸󎣡f�,�x���얂.��fJ���g�����#�@$��s����:����n�ڸ1��,�b��wm�7RuH�;[ֺ�r����ƭ���8v��۶�*�1*�Л�k���:Ƴ���*�qkv�/|}���M�u��<q!�`���8�x9���v��N�]'5�����P�k�0�����}.��ݺ��D�75�o��n���{PaJ7n�֝��V�����ᓰ���Qu]��PH 9�{X�w}�0��^�vj��6�L�y5C��_�e WGUǁ;�\�H ��f�=���O�; V��M���׮b|]��Lπ^���R2W$vD\�!�ν,S��3�#��I1{��I���d��~[ǧ�7�k%r�`[�c����农����}�0lH<�J�����ZO7�@I�L��d�O��Z�=��ߞ�N>��rh��J&-c-vbv��瘧d�۷Vy��� ������w��9+,��ͷ˜��@ �zi��ད��W6�Vl�k�y��������r���V�L��gg��v.�r�"�RooP�w���ΩKt}�ʅ!؂�u�!�޴뺕��r�gBX��˼e��a�����t3�r�sX�N������ٜ�� н��>A�;7�2굘��^Η�����5A�(�-�#ӻ�� l/-Ua �#=�gѣ�S*W}�'�!���H�^�S�k�����Q��>�ܬ���u�}�D��=�ɢ@=%���k�:[�kl{�����Rfnf�\����#�"��o%��'�f�cg���
�&�j���n�4E��Ut+�;s�����$1�y���tc/]���##ݶ�l�l�r��6�8N����pܠ���o}���	ț�g�ќɤ�:��|y�{t���o������}�6����(̋ۮ����d)�9��}���B�!���Մ�A�W՟Dw��m��^o.��ϝ��ۅ�hUUc��z��� �z[���ֺQ"ƕtt��mo�su����~�2��;=V�c�P�*�죘��ܝ/���� �c4Q�d �w�f3���̃o$���<�=w�A ��� I�}��m�X�$�yyt�y�ӛ<�͑�ë�����Ut(	�����_��l���&߶f���uT)J8���y��"~,�E��E�̞��J���~�Y+>$w$uoE���
�`��B�M�q�nx��F�ѵ�������Q�Ǵsnwk0s�X?f��2��;b/��ޔi��_k�B���<�^>u������EEWD��ǻ�ɔZ�iQ%"E����^$��p�^��UD	�.�H'鋥On<�m�|Y3��|r-�v��r�t)wG��O�$���n�����.�o�p�~����t�6��ʪ�P"�����8�>/wLN���lA3u`�=�q�V��і��5ӻ�T��M�C����'ͱW�l��>�u��Ң'�Nf�+t5�V�����v���I���!���L�xp$9�o1���betA]�k�vkƓ5��Zԫ���Zk�Ky��!�IXI'�/u�/;�M�猺�(�Z5��V�z^�ڷa�.�S���D咸�"����AXD4o�~:��ԥDW^{��X�ގ��M��^�zm����r�k���'�>�'�/�8E囱����2+�m�xw5����z.�A�	��I ����6/�SL^O`V{>u����ϛ��̡���V ��	K�>So=�lb�;��~/u��EJ9c����f�i�׶�ϑ& $:��g��"~�z��c�n̰H
�:ω��𫿪�UaX[����@$�y��g�C�_]fm6�swV���ֹd���;���w:����s
�?m�箑�}������}�3����'�YY;�e�3v��i�R`�ν�nXL���4����왁�
f%��9�����<}g�a$�����5��؜b̆�=�wjxpH�ѽQu+���BEXɲ@��7�aW�.9]ݽZ6a��n���:�t���c�tI�
�G^����Þl�����5~�I^�n�ħ�B��$u���N�H�k�z�O�5]����������9[PԦ�࢟E��9���lS�Y`ܗ1l"+����Uy.wxt��F�<���Y�룭ڏ7A�N^�Ʒa�[�1Y�����-��m�a�U]j�T��Xj�M�w@J[��OfI�o9H�9V̶)��wc��sB��i��%:|��?vc�bn�=$[,�/�(NfX9��u�3��z7����{��v+R{8[]�y�&ۧ9�y^d|�雼Q��(	�������7G�t�tL�g^�*�j�GQBq�U;JP:�.�l�2�ǔ6-�z�<st����[�#�o�s�ӭoF'Xa�v�d�i�Qn �t3xl�}�fݸbV�RP�e����:�֨Օ����6�s��e� ���N2�gsU���X�0��o�����w6y\b���h
c]6w�nd[����)op�l��Ge�7���A�^`Q����q�j�>��:�Ӳ�;��޻��G�7U�>������KDԱ�˲�n����6��:o%\�!��i��{k��I�de�&HPu�Q�����눲ȷ,�+)Ȭ�N�6�H��쬈�͍�l����N���m�Gi����.k[me��Q۶��;:�5��c�,��6��+"ʎn�,��g`6� �f6��mKl���-��M��Ф�l�4 +�r���#�;��m�Y��tq�ҷme�������(I��GNm�m�V�ݶ�K:��E$�,[t���Y�h�ΏmI�r�:2N�2s)��ȍ�z��9ֲk�gw��۝�m�����4�JE��]���ڙ�0G7�uA���WkL��*[U��s=c�lY㝋��͎�R�:�n�Hی���I.+�`:�6���';����y;a���R`�`Ҙ��q�����s�q�8�	<����G�Ocv^��u���=�$���I�Z�Mϝ�6D�6���p&������|��)c���vY.ȃo<mP�a�i������RI��B�au�����vY��d�nK<k��^&*����[��O��c�<vٽ�l�۪sɻ�l��S�竧���]���\���n��=q��xǎN7]m�u��f��ͤ��`w��vB��nwf�^���:�뇷���n�ۥ<u����{\˓K�4�޵�F�79�C��y��s #�+mH�:6;���w8���%���i���v˻�`�VՃ����J��/nû��o	��-���Q=nN�$�y�uʍcn��{R��S�<x*����p�\��ܖ��;�I7Wm��ύ�j�6�9�x����x�Ӟw�	xn�Mjt���mk�<bL.���=�{�������0��,�H/O%�7d����ηI�n{z�5+�y=&�Is�Ǎ��OU�=�7N�`쳗�v�Dg�frGJ7<�5]��<�Sl��SQ�n8�&<�;I�eB��x��O9��'�d���&�:�+( i�,�H4*�B�;�A��1��v��t�mf88��G�۶ȇ�^��#�ӸQ�p��n@�Y'��]m΋V�[A�5��>�r��N��\>�6|ttd���+��	vxn�֨{�4@�[��v����0=�z�p/��l��qư��B����>����lZ�赱�kv{<ӝ۲���e�n��Bv7�d÷ogN{x�q9���ٝs���s�F�`���q�n�<�ptv�<B�;�-a�̔a���\k*��� Ӈq�Я����6�-,tN���c!nlx�=��r����F�E��Z�s��8�����mݦn�:��1���r=�ݛT�����
g^�m���6����n�E��2n��9�S=���M�瓃�;z;<�c���2��YR�C'g���Y��۵6n�޴�k���2��e�Z6:ȵ�ێx:�����C�1�ڣ����Hʵ�Z8yV�M9�:���A��-���hƱ�pf�m�j���n��Uz��G9獅�90�M���z�=��\t��/<n4u;��a�YĢ�v�pk��"�j��%:v�ۄ���Sp��w5�CG>+,r�"�X�Y����F&WA���w�\�o�헇�]�߳>����'U����P P�9�V+��è-MJU#�����3�23Sw�P��j<t
)�� ׳́B�խ�y�B�{���j��(儍�ˤ��
 ;�����d���������|�}�>~�߳W�g1Q��S��U�Q?�He���񊟱I�~{�����ח&=���m O�ʜ�FE��"��SN_s�X����S���u��Yl����$��ޛ����f���矇]���{�`�4�@�āǱø8T�㬏aܒ6�y�9���N�~���4i�
��ͭ|")��V{��H�%_��U��%��gO7Alj�
��P�-!�S9`$����s2YZ��b^m-�WJVwW3�ꬸ�3/;�-��>�j������ݭ����^���u�y#J T��9;g����Oĉoݺ	���谐C{���:�������xr��&;R���P�{�|  �[���)d��z�P�d���k��ٯ����0�,r"�]'�3kY��Nަc �rw��m1�W�B���ֹ�sh�k��|پ�x�_Q��Gr6�źE�Z� ��Uyح�Ӑ᣹�@�%#b��Р=�9^b眬��-Eo�[�+��m��y�l��vY�8��玧]Y*'&�U�di� ��<���	��UN*�MA'�tXIsY(\KkR��1��wn���?]��5j�"jº���r�.�%r����;"�H#�l��;�Ӿ=Zyl�	��� ���Bд�	]ڰ��^"	�͌BHӖ2���j�t�����e�w�F���z�񗆵�����:�So,T�b�+*���݌X2�i���dΧ�_j\����ă{����S0�����U#����s�G&���S^��l��g��H����I�{QJ��z���4߲k�׻}�7b�P�ZʯNf�`����6���|�2/]�Y���η�Lw��g�T�#��(�7hZ�`�Յ�\���;r%�)��k�nq�{^���~ܣ]��TB��O���Y��z��G;��Oou�e]�Ҵ��fP�~ζg�4������*��i�k�ı��o��_p�i� ]��U j~n���L>��������B��O��5jɤ�^��=L�5�O���Uŝ齽=|�`�;�̲����h�9�ޘʚ��B��v�J5�����W�`�q?&+�wƇww�]�`��ɠ0�̝����b���S(ήU� �99���I9.͎��R��ɳ�:m*M�;�אָBǺ�(�p�<pS��Er��V��r2Z�J�w19�k����Þt��\��4=�U@P����C�{�]�c���L[]\�iV�
_�SL��/k�8�����kf��D��0���A07�{�:E%E*Wf��9�׈�H�6n�A�O�~ћJOy&&�@v���}�tr�ػ��k
�(N7��n��0���MO�������B�QV�u�C�P���*J�	X�Ϗ^>ߴ�x� a�f�{-�g�� ��`�wրV<N�Z�wvU%ah��ѽ]�3����'��n�H'���C	�OR,t��'��=�߉��#�_Ԯ������Cާ�S����{��!'���H�ϖ|I�{�[;~1��݊����÷�(�ܳ����_#R=����^���%��� �W�u����k����X��z�Sf�W�%���KT�
���E�#�ݯ^�M��i5��/7�Ǻ��pG	�*��0aOk
�w[�f=���9X0�s�u�L7/M����Mx4�f�\{�=��s���S�أ�J������wny:�S�狒�Z�v���9ϭv䝍u8ng�yYnº�Έ��z8�Oh�//<�w8T���K�xvu�{�s�mk�!�Z�:�Fs�7,���b�v�嗗{�wnѐ:�.{v½���6v*��z�z��E/T�n�bi�I<���(��f����f�'��qgǗu�n�Wd�IX�ÝZ�u�X���^Μ��B���� ���bZ��ͱ�W[��m&��3����;��)��C��V>�>xc�w����谂y��$F����Vغ>��	�şm��F�?V�?s���aUK7y��g�F�~V4�*����t����{Q�D�zf��s�*]����]G�#��!��c��}������=�m�$�:%�	�*�Y$�h��=��C�京Ý�p"V6�4ӂ 7E>�w����(�.��5`�I�O��$��y��r��������
�t���b��W,z��E.b~�5��ۢ��z�kN�`�Ϝfj#6��^r}0��8�Jx�m�=�{	�� 7צ˱/H�;Y��K�'W5�W� 
��� �y��	;b{z��m�Mhh�����[����=t�iF�O9��,i���z�s�;L��2T�~���9�F����5c>-���=^���uX�����7 D��=����<�����gvjٲ���]�Y�;��6�<{�`go��{o�F\��~$>���H'��Y�SKڃ�^A�!�km�{qN����v��Z��n�ێ:m�� �;Ym	����7�~([	T��ts����r�����8��Ք%�bo��'�>9�%�~�����_Ԯ��B�]ڰ�Ǣ`��^�qs�s�&L~�$�)�Z� �1��'Ɔ�����'b����M�d�����߷A���~$%VV���y�V�&fo����2�f��4Oe��:#I���_�5�aM�1��7��<�ta��3+��x�t���� ~׷��I��~�I�N�FD�[����5�ｍe�Q��|�`P�;=hP������8�#k�����/"/l�Y��m������=�w}x1x+r�)Oqs`�_�| =EW˧o9�ro��9�'�)P�BT9*�VP�a;���N�knzp�vu���H��������Pr��wa!Jz~�O���	�)��|eӵ��D:vn�$����~V4����G	����=��S����t׾ŋ�>Mha �T� �$ʃ�z�`���Č��Q�#`�!t�	]چ|F�~�I �s������[@P�օ�z/�r��Fҫ$�an�x��a���ޫP��Z ��~����z;��q���p���������Wv��b��?yK�g��\a���f�VwB�^,wWoNe�P쮗o����6[R�{�D�u��������=���Dꨄ��O^3��@:�j�Z�VѳB��#XOW�־ 
Ǣ��=��:U�k2�ؽ �|J�"�0�F$���
�U�c�n�!�r�m��� ���|��\�b����M@����
�^��x�&q���}�5�����x���PX����U��5�O:n��Ԃ��X�9�X	�Ci����>�^��𛸝�{<�4x�+-�ʟ.X,���[���U��({�F���鹼&<�'�H>�Og�{��������
7�#`�F�]��3�{vP#�� �}�( 7WF��;�W�hӑB9ռFe�rFҫ$�an�=��Ӡ �m�Z�S#��'��� ��Ѥ=]����ۯa� W������\��B��[Q/�3��˸�YN��3^G�u}�>&V� �ۤ���f���3uVjGo���wU��9���[�7o�z�c`�ϴ���Kƚh��n�M�든�nQ�Ȋx6"Q�&������籷
�X�c͇�j�М��]tGn�w��ذ`�1�^��,��:�+r<[	���=���@�땰��K�D;�W�	�/�D�i0���nt\��4�ꃪ�s���i�:4Xڰ2���ct�{�u��MXG�{n8ݺѸ'��۷O���&մ v���7��t�7Ζ����?o��t%�	c/���F�w�� ��������[���V������wg�ar ҭ�uwB�a��>r���bc��-�<��` >~[ q��|I�L�Y���P3�T��?*7�2�Em�I�=�w6���4�M�֙p�sR�d����XM!��&�eI\���Gy�кZo#i���?� h�m�� zylN^� �7g��9*(�LVV-}���_7�o:sjlY��$�ӡC�������H&T�`${�7O>�~|W�Ѡ�PF�[0[1�ay �mv:C�$�F�-�	�J���������J���]�������	����|H'�ީ���|PU�i�={�Ov����ri;�zUBP*��2�>��oZ�^5�=�����N$��`/5{��0++9f+��ft��ݦ/�i������b,��qB6������y���w7�;}��L��g��ꛈ^���e>n�gwx2eU��n������~$�Sp A}�^U2<��n�woŷ�Nw�M��y㹥P[Z� �H��A,���!~�W�㝫� �|wya���m`'���y�WR���j~$
k2-q�d�Laic����5�6�˵����7�=Z��
Û�H�>t0��碢�rUr�W��R
�]�DC'I6r�nQ�b.yz�Έ;��Ȗ�GI��~^��Q�����^].�4�?l�iO���֪�a�?��@?T��3l�$n�Y&�]��[~�4����E�ZC'�ZOĖ��a?�s� �����u%�"���|�T%AP�U���m�y�~�O|7ږ��e���C!�����5�VQ��Y���AZ̖��3�m�QJđj�BƾMl;�f�\�0
����q+&�Znfu-�h.�{�s�H[�fr��[�)L�42��[ťETXQB���ۨ�+-�=�_�$��Lx{��eN�Ү��R�խV�,�ox'}���%�(��6�Gy�3K��c�[v���%��"�Y��]�,V��V ��5��^�aj�3�Iԩ"I:wUm*z:�f3'k>@nX�F���%΂i��{.����gP��&�j�?mA��L�x�v���Ĝ�[���7���������;�j�,[v���D�٢�9�"Z�¥m]ɗgsX�$S�uᱷ@�t=�۩�ǟ��ܞu{y[��N�WW����9g�`�&o���t�yk�[���^�M���z�dݷI=�u�n��q"�V�f���9;
ut��B>�v��sS�Æ��[�ƹ�㹗�b��J����;�t�S�Z��j<�b�.�:�䮮�oU��cx<�,1�5-�^Ě��U�Q�Q�1�9�ȩҲ���N�U�*�!�}��Ks5,�G+�<$z;��jJt�s�C�z�����^V��v�5W=�Y�Y���.݈w"�z���5��6L�2n_^�)p����K�D!�խ�ì���4�M�T]�TzUE��%=7�&�1ui�e����c@Ym���Q�9X��T��� hA3c*g,'���5>��]��)�ԣ
��J�^]nb�h@�s�X��f���1_��1b{:�.�/kz�A�2��Q�uӗ��{c|�i���m&���,������Y�L�:	��a�۳�mqf�ųm�m��ڶLVۣ��Ֆ�F֙[�3�[m,�L�[dv��kBi�g%bQZYi�6����E'$��a��&ݧ$ln���dv��H���s6w-c[m�ܺ�nٳ0��[,��De�hز�;�c�-��n݋vV�m�l��q�e�ͳ��β��ȭ���mmm8�6��5���lu�e�e�q�d�.�lGi��m�f�m���'92��$s[����٣1�aܗͻ��6e�4�%�5�6kSkN�81�i���� ��),��VM�;,�+L�3��[sj��N��m��6NSk�9vW5�ΰӨ�'m�L�Zvv�@V�~�}<u��@}轭�/ IU�n��X0�m�9|���m_pU��� Ǎ�OWF�{=د�n�c��Ĉђ�QV
��%�3�����X>7���;�6�(�v�|I��<�	$J��
}������z�n�Q7cnq��ָ1�<���%z��U��i�a���8���a��T�cWiQ�p7���d��A?+�X	��{UKּG*pU��	=����;�E+��Z����m?M���L\�)k�7mTꄂF��I2�5��y����W�޼]q)�_9+�J�Z�,���ѧ�~>=�I&�Ϋ�֨lxo{z��A?7��I�����/���	PT��O�g\�/��4�N>�y��H ��=�7�g:�� �������^(�r��UL��==�ؖ�[����(j4�,
y&d�Acu�ye>Zf�N.�A�s]6��LV�
N��/�^����
���{.�����Ij� ?G/����#u��$�)�,$�S+3�����R�U#���QJ�]�mjI^Bo9C�1�4�m�//v�r���O9�}�i����#yL�:w�t�8��z�M/ߦ����v��V�'|G� �p3���ٳ$��E���ީ��ܯxs��eN�I7�C�瀣Eu�KZ^/}4�m>��&�x�GMj�~|߁uw5��'z��g�Y���Uvh,�z�fFZ�럽4��$��ha��X	&{9�7�vwĪW�k��ҡkeL-�t��sQ���k�����޻��c�7N�`'�K�Z��^�����\/7�&7�J䘤���n�[Y�9̂��vs��1_O���jn��5����r���Nf՛������w��8:�zY�F�kZt
v>�����9��N��q��q�jz�G���X��bv'�{<�ô=kk'Al����0;v�GC{8v�E���kft�Mq�a��57f�3�:���v�����)ؠ�ka���9f��2I�:':l�l�N��5��v��f�s��8��kn�psΪr��f��g��]Ŷ�,�6����Vs���#�V��[��I�����m�V)��V�E�:�i�le�a��wIU�u��*�8�:�th7ΰ��`}h#�^j�Iev���y�kg����~Ň��I4�{���jo]��E,���<�EՕ�����^��	��X	'���I�]ᓱ��s���OԆ�.`�5�/'�����ˢ`�7 sa��׹h ��}t(E���]擣Et��=鼹k㐉���� A#^w�i2�4��u-.5ח�Y�,g�:�ŹfEf�VEU٠�D�����UB��}�P������٤�U���q��>���>��������I��j��B �-���>�ƹ�-�cm���������p��O[3��?�O��w�'�H����С�.��@�H~���ن�'!F���f�-��|��Z���R��m!5wm�\d,~�aE<�y]�'fE��k'���{������u�M�<hB��^�V�\�R�c2>�ZmwS�/���{����, �}���;4���6�r�B�)e4�u�~$�}	�,�.Bʳ���ߛO7�sX���{4�DX�M�lV�Xt�TmU�Ŋ�^<������������6����:\��]}7I��]U
�n�*�G܃"z��B�g�O'�/�ݺ	��$_g�z��I
�@����ك�����Rl=�y����c��cƶwݎ,v�$v���m#�vA���<WU����w�]����$XI?���ڳ��&��f<�ɺ"S���b���	�Ul����;�'�[O3���A?ꛟ A�Y�K_e{yZoDׇ��'ִ�Gu���<���M�;�K�J���&Y��>N+w�ozb�I��L}��i��^f@��{s�s����t!�	��kp���А߷b�;���L��}��M��x��ޏWU*�A��]��G^�|H<벰�~$��$��s�5��i�P7_7���Eǹ�c��s�=�(�|�����)G|���z�L;Ɛ6f���L��3��xs�ݱ�����Q_R �S�.8�۔wl�n�rA�. �UQ��� ��\������**u��쳝4�I��vs4�'fs�;��w��,��VA�]��v���]�,��4�soF��/�,}����Vu	�?;��N�s�p[��j6���O�Μ���Ȥv��s/UX���lPT[���-�(_����6g=�F�I3vH������d<���:=����V �����	�������,;�ou��P����lo=;�(��rڲw�X�f�k3���)L�NW1^M_]�CT�D/Ff�w}=���y*�_������34��^�WUZ���׻�oީ+>>����kI˥g�y�y��H滦�׍(��~���=�ֵvT�)�;��[���un:u��n��L-r��mς�4&�ߗ= ��U��UV�u�W� ���AF�P�hV>�J�{::J�g�;#�'�<F�X6M*�F|;�u`"��rǗ��0�z�|(W��!]�@|=�'��D7�[�';�~��*��O���k6{ՀIc(y�=ӰE���=���M���l�qs��)mdR;`U|k������O��y��`�� �G�k�$��S����s����{c>���*�R5kA���^�7�i�gvs^+�E5����璠��üz+O.�n?d��b�B}ڋW�H�O�dY�;7g"��y�kՂ���'e6��5^�Ss=�`�4��n�-�s!E%��������ѣ�<��n��j�rێWz#�����jz6w�*-���ͬٷj.��8���v��x72�r<�tq��WZ�\�d�lm,[Ou»[�J�㶛n����6�݄�&@����e��ny3�Q�;�0��zy=k�� ��et�r�t�$�]����gu uϷ{75r]A�}x��N�ላ�p=��M�:��pv�Om��ۈK�t�mz����]�]8�x'=�w6.w.vܹ*�G�f���t�PnZ�~I�g40�O��ڙ�A �?)���F��˥����9����������6�U�	�{*<���]K���V!���A<��`$gT� Nș</�.��/��f�� l����z��Iz��"	1̺n�k&��� $���x�V3����h�PS1'��?]f��N����O��yoP�	ﱌ��iA�ʾ�&з����)�.�׎oQ��r��qvZ^+O7|��ĭ| |_+�����M]O��{����:6�g����n�xoBy�;iuų�>_8Xܒkq���3�T5`���2�Z�H$�V��"O��� �n��Nh쪂������[o�3�J6om)J�#��i9������~�]�ܺ�~��ѭt�H'>Y���υ�Q^]gi�C�����n]�b܃rDc�s0��v&b��6�p�y
�
^�f]z�K���L�B�Pt����gg���ݙB��b������#����?����y/syv�� ���<�vtW��&!U![Z����Әus6���<�&���*� >�� �w�ԩT�yX�:j)�WUeZ���A��������v���ý�g	$w�f|Oĉ^�,���9�U_y��\�e�Ҋ�OQ����ºϏ0Z���q�F���rY�N����Bʈ��iU���D��޾�$�O�^�,>v_.�;����7�u��gצ��QJvTŠ�^�S��Ʋ��b�$췘H0����,��W@Qָ�O%]����T�ŕY�]��@#�?P�~<�KHB3[�m����n��و�?���F��7�!�.�o�������೐J�Jy����������YS���}���3�O\���5ެ����W�D�b����*����P����u�^ O��OՀ���"8L����H�����z��D*�Vֹ鮚I����[��Ƴ��c�����繘H$>w�0{9M!�UW��ޓ~�HPP,!+N½��m4�q��a��X�
���࠙\�>����%es/	�^�L�_*θ�P���UM��/H��.�s�9c��~8S�-l��J:�̙���ygn��u'�շ��>�M� /_#�_t�N���n�2giF��M}vE��\���H;��Q�����v�K�~8	'��]5�i��-������#���'{��ՠ�ذ�$t�g����h���ko�\ʈ��jN]�������BF}��BM�Y�S�Fמd�G��6�gV:�n�ϳR�U�݂v�n�ۦKLwH���P��/��u��fF��b���q�H�r�c�)�OHߺe�0�����`�=}�7�P:7���Gݣ���d��A�$Ӻ-]+��{LW(1�V�;d17HQ�g�2��v��I!Q�[^��������V L�*�%麲�����r��Mɂ��<j�����ж�{7U ێr�/�Ǩ (1�m H���$�9%���*��q����j� ��J�>0��Y���>ϥ��H�+*�-\a��=}�}� ق��5�����!gĩ��}��']�	��t��L��Ϳ8��𭜻-��UU\4����M���m�g+�ct;!�7�B���隗o�:��|뮱�D�\*�ʕ:��\�4d�{[Ȟd�ܰr�j�(�s��M����2w(��WzSu�:�R�^*����{�DJ��,�5K�q����X����Y�M�٘��#F�ԽQ���;�[2���H;��	����֫dʲ�y���?T1�V[Ik~���u�|s��9�s��ۼ:�T��=���P�ٖ�9���̣�x�v腕��k�Xv��.��eI�z��27(�d+ԑT��q6[���Nl�n��vj���.뤊�R�>4��k.��#GUG$�K>jMߙ��FO`�~�vK��T��Sny}����`�7�|eotn����_��f�֥^�X�V��/�k��oE|��Kj�3:�������n\�ݩ�������T,��A�z�)V�D=o%]Ҡ�y����=&��uQԭ;aoƩ9QZ�f-��o-��.�5m�*?���gqW���yŋ6����eO&��5��sQպ0`y�op�%��&ˤ������6f5ټzo΅-�)ʽ�8e��}�P��1ʊu�6p��Qs��VJ,��]�s�uIx��/a�=a[6pF�j��~&&0��@��Y����I�y��y��VILU����.c��k��m�)$��0�Uk��z;�\k����RT�Spp���;p�
�Yu�|����&���k(�������X�#`_+s!�gy���!���Wӝ�I���f�t���� �o���qm�T 
���ZI�p�٘�aյ�%;��5�"̶�͂˰rF�'l�d�\Y�ۊ6�m��f������gdd���̶��59��,�Ee����h�%�����d�١�%glյ�D��;e�δ�r�4���6Ͷ�q�'Z�:2ƛ��5���R �Y���8����m�-�w��LЎ��,��8��4���f����L��ӎ�
*��f�t��a� �+fkq%���v$N5��"����&匷e���8�Ӝ v$M��(���v؃��8�0mYY��[�9�am5�����l]%n%�S�흶�c+GA�n���;,�f�;:���ʹvY�&i̛-���E�n$�l̶�v(���m����ݭ�s5[i�tK|�⮕?���
&UD*�)j�$s�N�v\Q�9�G�^�M�kmvO6{�1q@WT��n�n˩7Cq=^
��b�]P���tE��Ϸ�Nv�rD\�g����(Ŏ'up�ǎ�6��YSx�g��v�=B>sc�p��Z6ۇ� ��{v�F㝺��2�����Ô��.q��N8@S˫���!kkiu6�`��wS��'	�k+�̅���s������xu��;�q����f�b.vJ��������V[6���nx�t�����M�W������Ɋ�0���ݱ�,�l5���=��7]tmӭq���<�n�%�����lظ{��@��N�r=f���m[���N\Փ�։��{h�)S)�nwMۭi���շSn����Cktv��=�v��m����euV���s���l	kEa�*�2�b0uB-�@��;��ת��շ����ѭ�����3Sv;z.��۫�]:벧n�k�O�y�=�&���ݜ�5�l�R�k\�tqٹ�zOn�X�7cv��ǂ��`N�Z{z�k<s��E��>k�c����kY����'B+c��\��e`���=��n�������������rb7Zs��k��e����=������NtI�^Jn3�g�ewh�\xӻk���tmV�sۙwMnZ���I&pvٰط��ã�,&{@���6��Yy컵=���و�t�b˸��۪裒^�Y9�eX���Bv6]�vܜ�9���v+OT�ŭ�*O%�y��szQj�o=���	#�{����a�3�*9��uH����p�����cu���Ӯ]o�s&Q5m���[Y�Fs�k�v
ԬV �V8Ub��{l���۰;�Y����sp+B�:����=r:���8�M�۰��r�#�:N.��sz�f�ɧQ8��|���o%��BE`��競��78�&��G�9��c��R%/d� ��S���m��W�j�tm���s��r�ܾ��	ڵ�[�����y� .{v'�ˣ��T�e��TN�wXz�V�n�\�<���:���⺃�3�۫<era��=��`]�jy��v��]��b�`]�ƭ��^�ODۓs�pV{[��j���bOkV�n���/�]e�\m�Į֬n�n,�9���Gi�%�I�m���� <�f�r{\�;�v]۫v�lZ��l�����x��y.��O�kt��Y������@��&��]:N�Ъ%�T����L~$.^A1���~�}:mho�υn���vU�# �����o�������A�bE����On��!�Kވ�iYVU]�tm�A�^8	�<��>G����me|�;���G>���r�"��H+7j�:�	~���&�O���4��� �AJ����e{�Eǵ`?.H�����f
ʶ��x� ��S>��~��EN����fA l��ω$�S2:u���ymǕW��;5kQN�GUp��\����l�f���DvÌ��l}��Ymb�������I�z5�0	�ۇ���͇�F��֛M���۷��V�bh���Y��Dk1Q�1}W�[&ge�p땻M+S�@�Z��]���J�b� yYus]�%Q��ЃO$�Uv��g*H���)c�����OZX~$�#w��j�a�:��&�'�o������,� �Ms�u����NvS{Mq�{�I�z��I=ڦ
ǑU3Jʲ���Y���c�
����}���pT�<���1HK�iM�l�nw�uvTJ�K��y7�@���>�з�z��G��]����S(H���O��x��D@�YW��iZ���:���waٛvL�u[j�P*�D�n�����u��dU;��U;Cxy4�t�iG�m?n���)�,V/<�k~��VA?u�>E2ﰲ��Q-u�Ns=�7z����;.�̸v��P����^��@P�+�9�v�7ڰ����o�]��֊�$�Bb�3�Q��~������Ԡ�m]G��vc�A<)���No�9�[��Vݬ]�����ud;��e�����ǂ����C��AW(L�λ������\�~1ּ�H�_f�����V�)Yq�;ݡ<w�j5/�Ee_`D�H�z��+�z]fLtsy�jP8r*���s�u׳P 1=-P�^�/�D=�Y'�r�V|A����A���ρ�[����{�����m�REji�7l��n+�g\A�s�;sB�V�aT��i0f�;쩑^8r�1��A�r� �zZ�{;�ɂ�rnn���	�����'��!f���]倓'��$}vGJ�aH-N���~����$���w�1M�)&��֪�)]�*��}�A'�z���>�:���v��iΡ�yN���^�XO��d�u���	���}�8�G��<iF	6�����&��~=ղ�r��#H;L՛^#.E}t��[�a�W�4e�;���Y�S���4|�G��#��Q�s5Q���;ۆ��|(�=~��<r��t�4�u�s��ʔ�����;��o�Ǭ���$,�Ǯ&?�}duG����{�|�$T����M4��ҞΝ'zf��s�N�`ꬨnx�:�>���1rvƲV[��nOZ{v��4�#}�?|L4��*��8������H$��=J�2 �ѫ�y�R�Q�(
�����f�;*r9[��x�7�Q	�;�ŉBg� ��V��x�WC�w�O��jz��K�ߡ#�euPT��M�	�F�Z�*�z��P0^�Sٜ�i����]�݈�=alb�����t�
İO�N�,��~'��V(v��Sji��Q�� ����]��,PIXJ�����I=�{~�s��5o�jO�|x�ń��}O�?�}�t�Y~�{��V��'����(�T������]o5��}�'|2����]�#��1D"Ȼ°�ɴxF8�'�{���?*�~���`Z�BU9���Iuǎ�6�4��\0r�y�;b��u���]��9�K5�ۑ�莽s��|跓,[����k�'<w�|�:��h.͜�m�S..ˤ7vg/���os�gr!dla�]�%�m/W��ŬvY3�װq.���\ۍt�m�ۆm��s�v�_�����-��|=��l㮸�lًb�ل۰ps���ϗ���8�8j;n�q�`��5�\��J�k�/=2�ۢ�w�]^�I%R*���5?'e?g��'�f�5֢<4wfت��`$���m��a�eYUvh-ߏs٣G#���Q��q�`	${����Og�O����V�=f�8�����[���זH�t���@7]KH�8{�ѯA'ſe�{�=�KǼ	
��hҲ��5�^'�+�vX����|�A!�Ѻ���o*��	L����B֟e��Ud�b�`)N�ify`<���O;�[������A�~�j��2,�����sk�GZ�������GA0ֹ�ks����iX&V m4��3�~�T+%R��� {��lP x�G/�s����L�<��t��Ʀ�<-*J� ��FuL�	g�ȫT�>�Zq���5{v��s�l���fN�4W%L�D�'t�qQ+م{�yh�A�{5kǌ�x������7G|֡)� ە���>}�F��<vK����xO���X���o��F*V��n���� ��� !�X8����������i���V�r2�R����;2���~�9����>���{}v���s����	 ?vM߉f�H�N"�W�Z'74������ҕ���g��>��y� �}%�>��;����q�ߡ��m�r^Z����74�f@g�@���������/ӽ��KT�9k���'��b��������ߎ¨Wz���G�F����̻f9��U!5��Gx-�'�J�󎻽Y4o̿y`�OǺ�� NH�k�oD��ǅ���	��˭}@ �-ڌ�Y6�+�w����� �坶��OX̊��8��n��A��q��Ê��(E�+c˽���g�;�X�Ubd�ԬB��Ш<5+�2��ā)�V	�Χ�ϭ�J-U�B�ݚt�"�j�������	��]��A����J���v_gJ�氕�n�Q��)�Uj��.��?w�=�l[�3xK��o�J+T �����tOᴙ]#�֔�+S1mp}�:�r��*i���V��=��b�pR�>Rܛ�5�'���o���N"�W���^��>=�(��o�7@��輛ݩ	<}��M��|wzJ-�9��R�쥥4
]=��5nW@��\�14��K�=XO���ۤ����ˮ�t��s��W����ajp���sJ6�����������H�%�-�(P�:����I��O�J�XHX'>W=�����0IJ�� �;�{tOV=P��;��mn\�Z�gI���5r;KR�sX�WTir�0L��yTUm�,��R�U��)������1<Wu����_��������>7�,�`����ϟ·���9�c��:�+�(�M~l���P[=���']�Yph]�T:��;*�2��*�nܛ�V��Kn�h�QƢ�����A�Ge���ί�P��6
�Z���ݔq|=��� K�t�����P����FS�,?z���g���v�I��ɺ	'�,��;����V�@Z¥���j�]Z�/���� <+@C{���o��	�[�� �H�ǋ4�kOV�
9�,�t3�s�G�n/Vb�3�k�@q�ŀ�OucrV��u����\'����S�c��I]	�ê���{Տ>Y���z='�z~�NG �j��H=Տ����/s��T;u�~�c�wA�>�/B��+%��r֍��_l8������[�j���%<3�A���;�uZgK���h��T���RomC�gV�s�jwI*Ck\��b펺�p5�����W=zS��'���S��೟1WX��sbn�]����W��4uO6d�6:k;a�狷-g<vǺ��Þn�㧡=Z�t���Cuh�ݳ�Ϧ6m����/���
���+҆w-�6��7vxηC+Z9I%�9K���\���/�h�\��"��j�mø���۶�B�H:�ݟF����HE�0T�u��*)��g��P�7f�ѻ�4��ǈ`$άu�+|=�݁�f��?d�0^�\(Q��tv]$�NoQ���>��ٳ��ͮ�I�+;V A3�|��3����g`�.�]��t`����j�B�R����#�-�A��4�	o�V�M:�:�0H�X�`$�X�R�]e�V^]�@�:k
aK�c��@;��� ҼP�]�������zڞV`��z����f?"R8;S��<g�����38�Ƿ2���T�4gb	/���s��������k���^0��*UP�-�:�wZL���Q�-Fx\
�r�׵��Y�㤎H�T\������Q���Mi���GV6����R����Z�|t�&�`5i�E�N��u	Il@�rr����&�#I�:��F�^�t���-K��/|)C��NmG�i&�M������;���y[�^�_c�/��Gd�[Yo$���G$C��[+> ��7F��݄�&Fm�{b�	Q5C��A�T�O�9�(�m<�{��6���w�U���u�� �s���'���j�Bѥe�R~X����ܰ#�X�
�;�b���ss�������kz=�|���䥪�;-��?N�ƒ8�՟�>�]��쟫e`�[y���ix�ji�z�=q��G[#�pn���N�:��O�/[v��5�;5z]���8q���q��f�7d�~���0 A����~�{�E��i��^X+�O�*�>@�	�v��!��J��uLk	�\�GyuL�A#޷7I����'y��vu簽.��B����4��?S�T ԭ|B ��bR�W����Z=W%�=M�oJ圭�����$Wczf&�W��įRʎ�ʵ��	���fY�)roAYi�n�r�����q	*c�,���"�6��؄���Z��5��#�W!X��׼��V<�U��8�D�X6�\ŏ);zp����/7M�$��%�ʷ�y'x�r�n>�qŶ����H*�"��VM�r;�:��gN�}��lO3�&ۜ, %���'�a�H������[J�p}ڙ�nsɶ�6���b{��D��f�̻�a+-�S(3���Y�Ѵ���Ԅ�Շ2�s,�EHNV�oo����ݚ�쩡qKLq�v[�ܺ�Ո���9��p{f��+znA�����^nl�ԥԐ�2��5"�_���Y�W����f&�˵���R{���]����P�b;�M���PӥVk�%���:����S�X�����v�ε���wJ�n�I����i
��q� )X{�o(�
��y�hU����q�s
��*E���v�&U���אY/YR�,�=�}w� �{oV+�t��r�z���oc���J�̚$V~�f]�cip@��G�9���8�5lM5��
��kO*Ykma�O�͜��S�4=-e:.,��!o�ۺ�M�o�,�9�w�y��a�/��T��'+LɰR���Z5KʯZ�7�U�@j�"�a`�rK¼�ݲs7ֵ8s�0��o����&}��իŃ�V;tBy�mO�6�ھ�}�9Ҽ�;2Ê��嘊}z�)����f�f��;1��H
��������A#~U��@��D�	I��n��B�����%kRڶ2e�k"�!�V�&۶����Y��fՃ��e���.��δ���e�ks��L�b2��$C�-�L�p��q�F�lԅf�f��(�	�2ַbm��,�3��h�m�ȗm�)�N,�mh�8d۹m�gm�嵌�g6ZQB�dfֺH$��;m�i�*PCj�A �mR�vݦX�1Ȉ� ���:��.Ⓤ�ʹg[4�9	va#��ū8[2J8J$���.�I;�ZGGGE���D�8%2ܹq\I(p�RY��E.I\���vYD�NGrNHI
w'��w$�9�� e�C���(��'C�f9�)AQNB~?	 +wuĂ~�\���y�^|	SP!F�褊�
��~������~�C�q� 
�K ��q��6m6�ğ��wX���40N�W#�'������_	��ȏfVsπ�Ny�K����I�Z�$(ך�;)u�W��J�#uY�{0q�7Pv6��Q��.�n���#�ۣT&����R�J[-'�g3\ń�D���� �宰��^6����ibm?{Z�_2��FP��ܦ�;�9U�/��Ԏl�S 'b�B�կ$�÷�ά��� \���J��Q̠�O���^�����DA>��q4��^;��P����V*��:͛F�ٻ4�����t���g8�bj�/]*�(
�o� {7���t��n�f�-�ذ������5	�I�U��+��+xva�x�����O�mOm_�Đ�-���zn�qtR���BwS�Ÿ��3��mp޲-)��Ia$p�U짾D�ɠh��e�OVT��	�����^ I�sɺμ�b3p{���:��r]���v����+MR��s�Cg5`��l{��@�������'�N�ެ$�4~�Y�*�o���O�3��ɧ�KU���M&{��`*�/r�/eӠ(z�H
���l
�ޑ�p{7ٿ�WoΖ�[��N����v����bl�{{�q��OyoĂ��09��$'c����v	9�1��]c��|:c@�2�Մ�H�웠��S�[�yWv�H)T�Y��F�F�ٻ4�h=�}�H�z���N=
��@&�l
�q�j��O;�*��^�Za;c&�v�׊�:lz��?=��5�~�̽���;����v6IT��S��e��\Y#e�|�����n�u̹��G�Id�ПK[�-���W.�֤���v��v�>݋�6��<+c�՘��vM�jb��X�	�ͱ�n��=�����ƨ0u�AD7����o����#rV��g���y�FVNy����9���@t\=��m����z�m��#�{p
�l��E�7q�cW.z���e�[���9��3U��[��N���;�����u�n8�)�89P���[Ф]���jۮ�W-%�����1�S�ک~�{�g�E%��IT��>�~��&L�H'�ެ75l�.<�#�~4�$k�4o�pd�Jѣv;e{P�Į��_�[��[W)�H���$��!����ʼ���:W��"%-�!U��i3��ō5�۩��w|��pZ�������#��Y� U���]
F�nS���x�����i���W��A2�����{H��<˯�w��	����J���c���Z�%ۄuV��g �m�n�I.�bD�ׁrt����A��xƘ6��'�.�Q�z�g�P�y��r��t �ZB��]ŷ���DE�U���H� ��&oğ���I'�宅U��KV�͠����c$*f-7�pꈥ�22U*�9�J6�G�>y_wz��w�1�PY�<�!�ōfR��P���B���ŵ�����S��6�p�_��*ez�{ܯ5��,\�!Sܴ�,��l�K)�U�+�R��;��G�����7����
�#̤q�T(B�U��="ܿz�.�T(C���m���}<K,���m���&�g�*�]�ρ ���0_�e`'�{�;��^����t�|O�ǌ|
Dꈦb��F��O۾�����D���>&�s�H=ս��=�������R�Ǭ潯i3��\Q�4Y"�]ۖ �y{cQ�<]�wJl��*�(�&X�TS����NB��w��桄��׈�I�nn��Orw#jF>T�,$d�x����F�V;���ߴJ�J��^����A?t[Հ	��߉%B�*�-�{.�6�\��TE-���\�N�����=nh�~,u�\�wa�^���/����Ϝ�\��0�n
@͔��Zک��'�P�����_����%���fGg��<ݍ���W��^����|�>�olb�.$�l��u���?y�H5%�V�W5���}�e�w{n!=�t�&K����H�w�`�F����߶]�]�7%rW$U[m&��ױ,`�x�����"��$ID嫕��	�����<w���{!s)x�
=ߪ�]sn/���n>p8��T..�=��iz�v���1���M?u>~<*��N~O�7�F	=��Ѡ�z���i�?I1�K ����mw��7��˳,r95�4V��a�滤�N��^~��1 s|ء�^�d�7aC��fy�׽�+�j���o(e�]��M�lPJ�� ���mۛ�4�.v�$�5�Y�$m�\���"�Z�+��2�h��s ��v��I�����ρ?����[�L[���Nr=Ү��d�b�%��٥l.�sxR{�\��3弝�`��X����˳_���R̗K/�%A��W]:33b{V8g�f�C}��T�+�B�$wie�UT �wʎ�/݅�(}�ɾ��������a$��O ���U���{�:�>�F���	/�ʈ�"�����Fn7&�;�[O&�*ڄ�jZ	X���s���+�*����4�;F�@/�^V|���m� �;�nAբ�rV���ءS׈�����f�+(
��z��}DY~�潽+,^V�����H�^VI3�<�+��_Y�m�9`�R��b��B:�T��O��ޢ>�lBU������>��v�DN��oW
6��Մ�������hv�~+��ω$�j��y1��%k�I��N��}�gV�#�Yt�5�(�~��o��q�	/q�ڽ���O�{S�9��"�㧆����tu�o�q�BH���#�ZW��=x�}{���ݜ�Ql�y	�45{w��{vȎE���I(��?�Ќ]E�fv:3ӓ�s���C[5Cj���f��z_]���ӱ{K�L��7Gn{N�p{8�GYֿ���͞���'�Wm�ݜV����݄�LM+k�:��م�04�	�Zv�U`�c�E���vvռvqz�n��q�`�V�[r�ZλlR\�h�b-�Y�q����#�7����vt���q;˷�{D95���t>�X���66�@���lz�$6�[�Z�8rO�j�u��c��&8)H+c�~KVg|�}�N���;ڹ�T�̋k��9�E 	���5�g�VJ��ZI�\�,i���f��O�� ��W ���&�!����X�p�v���5]�'T�Zc�/ȏ��zyy��C��Iv��P�Ajy@�'<��s+�
E+�-_ƽ�Q
H��)��\D ��o�>�+�qڙ�s&\��>��e�D}���d�Ala���w1cm=�\�O$ץ7�J�W��4"�ߎv�ē��V�ߣ8���=�^����Jڱ��6/Q�]�=<	�	���+����6�,�A�9�Ѻ���XV�Tk8Q��v<��~'�z��%��fi���#><�L�|��R6n��*�FU�XI�&{��H�vg4������a]𫥧v\�23lE�d�%����Vi���}w"��;����rїQ���6�[\q�e؀#���C���a)��	;�;t#�ެm��}۽j��Njnoh�9���Em.��{�$q��$��^�uQ�P�I�L������ņ�"��@�V�h�]�Cw*��v�I�rh��]z�	=ڙv�ڿQ�h`�_s��|ѽ(BKEU����y�I���9�]�ž���ז� T���P��P���d�ړ��^����[B>����Ƌ�ܲt���J{�5A���8�o�(�­O���y�a��A/�M�ءP^�@ =�K��V<�p�b��� �OV~ԝ@��j�%V�»�x	��;y�;��p� �)MXI �c�)�y��So�rg���I�蔨�f�]��ten5��w�^'���S>ܭ�2��]!x�c0n�>��$�[YV��j�u�Do�Sf�	��]qk��]wVI��=�H���D}���(7���7�k�I��z�-�Em-�z�nnθ*���i��t��`'�F� �;W3� W<3r�>�C�g]+��+ڢl+T4WoXd��ghܜ*ܼ��\���鹋> ��K��sɚ�o)|_���_���2p�'�O�{p%�uk�y��9umq�gnq�U�*���DQ�9�Ii[��%��_p=�w��H3�L�y�=�㒵��5ݵ��r줷]��9�yB�e�OsuLs��B.��C�L��$���0�O��&�?��[:3���f7�<uEc��K�������f��2xT��L3:��� ��B�mwם�mo���8뢶8fh�n��5��@H:�/$�F�ɣII��5Ҷ�12��㷖�*
�.�c���M�^���<���];iۜ�}4��^O*�
�N�3c<=W�3֛{��x˛�r�FYd��	������B�[���S�w�&�~s��OZ��x���@t_*ۛ̀���'�U)�O�����p���Qrv ���ƃnV��,��\n��`�����}^�����~s{���O�z��� �~�V�ʮ�����5t��6����|��Nj͐����h7��'�����|��^�L{}��I ��;��H�ԭ�$%���߹u���̝C�ҧU���>��X�kn^M&�&���p��ھ	������ma+,|��m	(�wI�ou]g7�f��E�^,AZ���	��Ԯ,�~3�ٻ֛��������@$w=�I"���v;g=��Gz�2o��Ӂ����|���������B�����	/� I_�H@�����%��I_���%�	!!K���$����%�i!!K��I_���%Ԑ��%I!!K`	!K���$��	!K���$��	!K���$��B� �$���d�Mf��phf�A@��̟\���0 �                                    X  ` � *� J  
 (   @(�@ �
P     
B�( 
�                                     �   @      J��Az�!ݴ4��Wf6s�ћ�t%� ����u��7;�&`r;�!�&  2 �
<    Q� f C#T 4@� �  $� ��C!�R PPW             Ht �:�CBF&�  H 	� ���@�� ���``P�z�W�   `� �,� �=C� L�����=� �C�@z@ M���
�
$x  �        �f<�2(  �� ���C d�5F@����5@N�
 )^  i���0˸  H�d@dTd�.8 �R����T�(Qي�iI
]b�M)BJR�  ��  < @      #Х$���� S�)J]e ���\�,�R��.\ ������)JH\� \Ƃ�Y@
]�3JHR�����AJR�#HJ*���W�@U&  �3J^�{g�2� �4ɺ�R�7q�j�ݣ��F�ݴ��� �л9:�Rr�:j�']�P@ t( �  �        �Jj��;�\�nfٹ���W�h,p 9Ҩ��;�*�3���N@1ͮN��g ��P��f�8�W)��� *�  ��]�Cj��k��p ,V�X��M�C�@�n�b�.u�A� ˪R�3��K���̗6�N,�uB� jy4)Q�  "���R��   �LM0�b`&���T�)S@  ��MJ�  �H$ʢi@#�=����������� A��/��}��r��v�0$�	&�O��xB�R�HHhB���$ I?�	!H��BCgݧ�������o0�ޜ޸���w&�񣽕�K"��iWNtE�N�&��p5x^����"�s�0��7��w
{�s��{��������0vn�Y�3�pr���z��tt�p�\v�n�m.���Ƨ)sqU���Ό#vl+��2��M(�l�5���{~��� �� �r�8��ڏ`(����y�e��@�������X�dãh
={ronoL�΃�Gr�=�v�|_uƎk����zW=��Q�p�{�ݘ2E٣�ni\�݀�����)���I �?�zA���ı�&��)��5I��WFτڸ�)�� -3S���e�E�6�����U��H�Kd<�3��ҽ�whʹ��%�na)ڞ�<�
���0,v�:cN�-PU��t��=����H��C�(�oeZ����ުN�Fےi�
�`�1�N��	�Q�7��r�nnfao������x%FǽZ����"����Z��X1c�p�Y��w�#);) mt�o����%ҽ���L����uzT�tŇ}�N�{�X�̦rv�ܽ˂� ������9v�A����<���]�Xƞ$��X�i[>��0U�48��
���,B)o�쐳�2e�0aYxѰ�>oB�Q������еo$�{�Z�vm���j�Չ��M��{$80������O>�F7�j�V�O]U��m �m�=��"Z�m�q�C\�4-�q�pC�^��ʮ�����qa��õ�'N��#���Qw��f�����1�"C��t�v)���Ƽ���*{��(M]绺`�`cn�>8��5��Xi\�s��U�m��ީ�s�u�����!����ے����=��q������UL��_=ݗ+�uXX���"�y�'`Ե����#\���ū��u�=:^r�Fj�򅑽�w��`����NW��C����y�g&껋�<[ܬ��8�Qf��Sf5���f�>�F�=�ƞ�p�k���X�s[͇��;��:wp��2�\�s��ѝ��z�q�������J����j.t$��U 	�Y���v@OnG�p��Ss�1d�C�׵j6=B%9v��`�l��f��u�z��LsCV�\�n�� x\�j�$	�2�x�� �@O�x�N����s�x-�08*(M�����w2F�.�z8]�*�`{�JP�:cwXt���"�Ξw9�����ǷF�u-�я��k+㶥�d�z	�z��xR����nn�=�W�jJ�ˤO�R]yn�3�o��u�V�Ļs���p�E]���=<�Z�І	~ױ�qAyǛ���)��`�W`(Q���Q����ՏI*rOBg�Ӫ��-�h@�.��朆��Y*,�)��y�����a��@*��svth&��0v���`Ō	��<#5sj
����k!�=�vb��jۊoĘx��9���2cX`$t��xh�݇8����Uu˄�DN�lh$�,��������l��ok�/qP���	x�v�tq�PC��7�����6�P��+�9����N���P�V�0uc�����q�V���ahh�r�L]4cM��2Z3EI��u�H$��ك����n��wMu\a�s�M�6���&.�kt�9N�q�ue�:�ت���0s9�X�'��kjVm���gn�(6���1�Gv���������D!��+��5����Y��̳CC�WF��F�)t�]�v<�:�Dwp94M� *.<�\���>��WOnB��/��#���P��'�u��b���ͳ�Q�;�m�vsʖ�*K&ю�M�7��q�*�w6�	���w��wɶd1�m5Ȼ�M$��;����&��&�,ҷq��|��y��y��vcqh1=�E��i�ov꘳^�.&
~{��§`<�W����p��Wm3y�9�ӧWL`%ۄ</y0B��=e�]9��.鳻H�Jy�ם�l.w���A��|D�{��O���.�"�^�{�i�k�k7YΌ�}�����;��}���7�=:����Pf���7����ucsY��Qr�n�#� ��y��wl���A�~'�[�މ��H.��cI�ij�Ul6Q�<���n��Z�Ŏ�)����o-Ho02w5�r�\ڑ�� �Y���� �����4�ݝ�p��� �*;�Ń8r����֎�X7a�lX��7s��~~���ܞ��B� 8��m��l��ÐtFR�*�Wu=�ڗŉ���B[fN�fn<�d��U�7*��ƍ�ز��mp-m�|���o|�B���L<,9y���Π�.9t�£����'�G�����|�v�_\��{�s�pX8����yx�~��z0RY+��Q,E����P�/�jo%e�üZ�lԴ�b��[F��v�˥�2�І��������ҥD��V�;��Yo�ݒ{�f���{�o�6~ٰ�^i��|m�6
Y���QVt*��m�]���)�*��N鮽⥥����;�xS�H�|0�r�Szx f�p��ݪv��K���'Ქ��:�Mᄂ-�c���vh/�S�����1��۵ˈ�9�^�3r��eŠ���5��a�#k�[�)�b1�¾�om����n�1u��;x/]͞���7��I�*؎.p������vjtf� ���ÃQ�Sn�u��A|L�ٱ��z�x��	sk�Am��D�x��Y���A^��ol{0��Цps�C��@��*D����v�����.�=�wq^��^,*��ŽX�ռwpq�CM�P����h=g,�}!f=�9H���b�{qE(nQbкn^��4�c�gE��4Ύ8�6�N�f�c��/�+���A⑼!Н-X#yt����+F�;���4h���U���M�.�6�}Y;�6jfA��w��x)u���;�E���Дy�pd*^�(ˇ�Zo_�\���]�8�\�N��Y��ۼ�͸la`��M��mU
���.8�M�yavL ��n�mZw� ��V�Y2�іK>ݙ��j�e�rAM`�h|���yze/C�;tƨ����|�5�������j}�2�s��
{����	��A���DϸݏcOq�޽�eX�׿�p����c@�Ƌ�bحS���n(�)l<�n�5�۴�|��js#D;�HU���=�o֏�W��]�x����ti<;WW&���:�1���MK����):�k4�ݦ��y�"n�m��؎ܧt�8�<@Ď��_>�q	W�H�syn�8�ă��kXv2���1F�k�2(|��[1aރLou�Ę�[��͠�y�v�Z81�]+�����Þ�S��ԆU<�ε�KwW^B���b���ԗ�>oڦt����؟�����"�l;s{f���-U���m�θ�bL�������� �3N@��m�Y1�z{�����;_6���8wF�XA�����B	�n����i�7���{�	neF�Y���D��d/���󒦌s/h��o���v�޸�.t��=���L����J;tc���9���ُG-|Bn�����T£��f�KqD3����ϐ�~���;�f��u�w\7����x��],�Uݯ�Uכp��Q�IW�Ej�ϟW�2s�j;�F�]���SX�����2��o�@ɇ8=h��zA���̬�����|�n0�Q2�a�0� 9�"�`�^�O٣v��썩��2���"�۫`[Ͷ����3�d�,5�h���uur�ʷu����[�s���
�K��qY�yb읍��NDA�����A(����Y�i��5�'7��р�]�)7lZކ�釟hCd���`W&�"y��Dv�v�k����X���h��RZT�"�f�-Z��	L�ܵ��	epD�L��4:(��ã����3;�/�q���l�@�r�l����po�y/C����R�r�;�wo6"���ڪ��J�i��p-��ι���l@#�+�{pt�OW�`���t��>ú6j��'G ��R�l� 7������8^ypXu�U�X+q@ٸC�aܛwTV}_8�<�ە�ۅã''�}��h�jK��+&�&� ��孙��.$�f"�1H��ߌ�GGe+q�PRz!������<TSv����\��RE�ի��*YI�ۣI�s��y��)��%ZA���ۻ���J���$�6�u�ܺ�W����kr.ڬ��:�'j:�)с�6��S��<并��)�{ȋ��}�s��vW�S�{���F��8-V�9��`���<'L����g r-�N ��{&nAZ7m��
����^�����y }��\�6�,K�&"�ޯ�9��Ʌ@�1�-��	c��K�=ؓ5�wN2^v;�2�������Cw/�ͳ���۔�<���s��;82�m��<GC:;�s���%��M��H� ���uZ� �(�w��
�\����,���eK	;ƭW�:����^6�޷��!�`��}wm�r�3��{�;���nL���ilue�L�k����wyț��n�`����t)�T.�B�e�݇'GטE��<஠�uժc��V����yL�6_�9I��N��Ճ�}:�;QΝ2�>��s`ْ�T���񅜎=��{��Cw�N��ږ����T��
�Ь�6"��r@�}���H�㗍���xO�ꪳ՜m%�V�ɍL�B���֮y��n����Z�F-D3�i��b=�����;�^�ӓ�ۗ4�"���4ri-p��8���%&��ߚ��w��h�s�I����:.2YoA��vJ93x�����ûVՎa㛝>]���pi��]��9����v�.^%����60W�*2�lD��׮��wY�Z����N\J�c�¶�+�K#�rn��n���4��� Y_=�d髂Jn��y��v<L\,�.���R#琲��G��#��oa%��'FheCgH� #:b��)�H�a؂( L�N�F;n���f��_�f�Fv	)�c��ෑ��Xaf��HvҦ��f������nƎ+��nnL�>��&!������(�Ŋ��
J�q�@+�����zt�&�cg#;ݛ���O-�eCkrb��4���/�����o#���145����݋uSF�9����;�3v��R�Jw���*�9�Ȇ��i��(�˥�XyG5ޅ��vY�B<3B<$ ���eO���k�v�Uh,�˞m[��M��K����z¬3��4�U�9��a�f��M��5�ϴ߻{�R����r���h���ػ���oS���4]	�����!��ŀ;��ڲE�m�c�P5b��p�q�*���WH���B%ݮ�t�6;#�
׸���׆��v��zY��g`ٸ]!Z1-�؜���.4�g�;%�'�/@N4�es ^#��� �Ns�ٺ7��e�ڰ�<p���e��� ،�v��BH������]X���ע!8g^	o:!�ٰ(�h[o.{K�x,Ltҕ�m)�N���Ϊ��C)�s�7x���M|��7h��wv��u��b�H�8��yr�,���
�%�-��s�yrwg3�H#�0�4�a��x��=�*�,N�WpӨ���]H�����C�Ӹ�U��,92���J�n����1�1��ԯp[����᳨���偬r!�w@�mv̆eKq;�.��JϬ��܅=D��dv����fE�i�pwn�j˚A���k&�W�b�E��0��qR>���u���;�Z�m �Z1ʵ��#I�rd��4�1�O��S����xqi�zKˍp��6������}�7�+�vη�i��3��}�C��4)�vb�f���AyWuē�f��_�
�7s]�Zxl�R��D;�.��K2Z��{'k�oT&��9>�x���NN��<=�4�R��ocG,������
ݑb��2}M㺒�˹7�c4^�ܯ\��(ݽ��yH4ps�]�k1�tOk�,u<Ќ�̜��l@�
�:̼���3�����=��.�YIV\��l�դe�ӆ���)'�h��\Si��m�qu�:>SF��7���r��S�³���4�=!-n�)w[�V,gp\�Ç����wy]s�=��e�"}ǜM�v�׶��$9���#uv5�z��WA>�!,L�D`O�wFUg�-3r̫7��v�����j��c]�t��E8e�@3�s��\�!=��֠+mh��a�+��e�x�<�=�S�n��� ��W���](.�&���"�e�+8�A�*�#�v�=�i{�pۖ�Zt�ӳ��ۛ� /-�m������n�����;#�܊,S�zlV�Ѽ6�^���g�ZX��O6�h9j'�����{�Ë�Չ��wa�1���>M��²�}a��❢�-Q�n�H� ���d��lX�k�E\��fS��OۻJl��p��v�δ����Gv�H�������Sn�RD�+f*����<8�xxxt�T P� �@��dAd�Y +! ���	�"� +I $ ���� �$X�I*H� HB,�EE�$"���	$� V
�a! ,� 
B@XH$��$P Y	 � ��B,a�(@
�I$��J�
�Y	"�H,����X� "�B)!$"���@�B��� �BH�I"��$�I!
� Y ���`�X@� �d�T��B,$�P��(� 	 �� �	+!	RB�a R�� V�!Y	"�Y T� ��
H�@�T���(I+B�� �B��5��}�Ë��Y�������ޚ}F���}�a�C�mg�{��<!��l�ISn|�Ȳ�Jf��ޟѽ����tW�z|���}C��sE��b�����o���iQD$�8=.�\ �B�б�ѓFl1���P�G헇�9�r���8�H���ׄ��Q����w��ň���z�i���ݝy�Z �o�1�w_��D�iF"��gnj�}��Y�W�W���	u��v��l �&>������d^`��9]0�#���ۛV��z{�'�x�=���V��h������/�|��Gyo�œ��_j��T%��7V��A�ϵo�z�E ѝ�n��t�ȵ�,J�a���׾�{Q���ٜ�DwvV{���Z�y���V,�5]�kހG�O��X���2{���^��&<�ֈ�*{L�4/KŬ��"Aú�f�o��g��e���H��.Z��-~+65����{#��+��`�:gMã��\VC�W��gL����p`��{���s�/��� ��gOhK�Bva��Ͷ���l�V=��B��Z�}�|��D�/K��2r����8���^�״y�7W����E���P��+���0���Mh��[;�&	i�oIzN~����4��1?x_d\d��U��py�i&Κ���|�v�O��֭����5������y[zvA(��D��o�Ź3y�pM�חg��^�g������*������Om��ͻ�3���R�bѻṄ�P����8e���f�i��m1��e�"���P�,$�={5����j#��m��0���V�R�x˛ U3�#hei��.w.M�Cݩ��,���y��wN���N�F.���mY�'7f�lnnU�˙0�Έ.��V]ޥ�)Az�v���m����豫u9��yK÷w�|1S����7�>�2,���pL��O��֖3Ȍ�SB��h��̟h�s�.�5_gN$���ף��}���
�^>ܞ^��]�%�*�*�%>����p��m��ˮpՠ�����k<����vz���fs5��p��|��#�V"yyZxz�<!�&s�fM�_]�Wr?t��/C��z.�WW��^�I��h���W�fK;8
�a��ǗN�D�$���}� ��3���U�?@��������� �� W*������.�o���xol�@L^�K/����җR���a��s�]�lq�!�w��H��S������{�q��a�,Ԇ9�(0`�{�#��gW���2���e��>�r�����5׺��罺7��.��"�:�\�v!����7�b{�޾�އ�u���Ɇ���L��������ܻtv7����Ô�w�L�rx����/^,ܛ�h����v�e���wME^d�l�ɣ�Fn��:w	o�zr���(��s�LO������|jK[��:�2�a,|1����Л�{c�djbh�+�okt�s���_{��M�8��Nt���ni]��������_'J��)���/g���`=���g���k}���m+ڎ���]⏱n0������'
|J��q�V���w9�<�=��0��;�/s�q%z�I�Fp��]�M����X�F�-F.�ϋyM�A�;�� Ӫ�v��7�ۧ�<�]Tm�؈��Į˜{�KhFs�M�]��0�{:>WW��X4��e��u�7��ݔ�e:���S��+s��f�=��.��q2M�q�n�K��pm�vogE��wы�=�/���������D-ǫ����:Bt��K҅n/F:�9�S�@��2�@�ٻ��ㅭ�w���v�=��!w�݌����p7B\�Y�04]��r/t�59;��{��mҏlHvE�M�oo��;��Fjl��،Œ��4d�/ɞ\Ҩ.�^��ۻ��Go����Æ�r0ط�=�b��2��l�ۉ��wT�z��\g�m�d��2^఺��������I`B�A%5��Vz�ECEj�L�W��q4�3l��8&��o���"�]���͹8�s�QI��g���Ň��yn��W��oMo��o�F��� <�&nu޹7�Q�Ŧ��R۵�B	�Éyi�{φrGc�FI��j�i~�p��Ia�	��f�􇣳r�^�`��d���$mم�Dya%��H��j�����.���@{���4��l琗&�W�U4�__r��/���_�����} w�u��oۓ<�&�w����n�;Ϭ�D{�X!���ܺ�����r7ņ�{�����n�vz����|�>�	7r^R}ڷK� me��[��ѓ}�}7&']�]���7s��9&<����{����w�<�9�_�k��	QH���xwm7����"p�BN̼�Y�j|�=ݬhԳ���+Z�wf�;��>�G7;i�=�;�����7����]����x��>�k:� h��<1��q��n3�z?Gi�9z^-YHo����.��v}�(�.$5Y�դcM��t�B�H��ֽ��F�2��!W�y�M=����њOye�AP�s)���Lv[�}���6����DޝS�O=�f��y�3�)�/{�9	h!�*K��$���o�G�[���g����A� c��)9�,[��x���R�{N���}�e���Ty�E��^C�`׆N:u�9����8�"9�{�qnmW!���og��{�S^8W��W�Z˷�Ljs��=�1N;�:���f��ϪSpn��3G������Foa�5�g1JD��6p���w���Q��r�.���G	S���Aa^�Z:�����+���.��9{�����N�{���zn`|'��ji�oxA�i�����C��O��5�\�n%x��.ʳ�%i�{:u�tn>�q5��^�;��^Ä>ݽFbhԃ�e� Z\dޯx�T��,����ъOo�G(�Hz����gxG��ho�uQ�Q}|h�4��Tٺw^�9���ϒ��߼ˠ�����|���}X'�X�����]�����������]��ډ�s4��gu��L��9bQz���kl[ۅL�{s���|׹�oo��J�u,^�Vp�����b�Z7�+Ľ��w.��w?�pg\IQ���ޔ��O�����y�]�7��D�覬�/�^�=ݛIU!�J�=��T�o/G�N[�O��H��2�MSt3��_r󤉝��Ǝ7����FEn����s����|.tt��^ߜE�x.�۞�*]��������L֔ի8t��p, X7 C����2����jnki�j�	7h��U_��'��FB�s���S����Ь��s���w�9b��b��ｾ�ȅ�~�rV�ݽ�t�|�����n/y]�njxP�y�ڏ��9 |�F�ԉv�C��'.�볌�,���&f�9̗ȃ�پ��"�"Ӧt[�y{�6q�}�}�[�j����!y���܁�!o��؎�) ��QdH3{��dMQ(<��{�SP����ʻ��r5;=��vy��>�g���3��`�O�����{��2uk�q�4oD	J�̃S��o��C��o]�>��-[K���O�����r��}=��Ac�� �m�.�m`�[��2z'�	��������5���ƽ���%]�]5O��{�&���4KB��s^O��^z�۶3&�=A�؍Zvע�ب�;7]���)�Ow
 ���|�~�懟v����a?u��ټѮv�Γ=,u)���.�7O�'KM4�����ۻ�^T��%%��w�n��l�Н�yW54f�B��&N�nopU�7VC�I>��q��5i^�sZϕ���!��kub8ox��c��0N";."{7�*�F 1R��ܺ2W�}+)]Z��CDZ�uɼ��]�����7���x�h;D�	���m-»����6܂���q�𽌣��7q�N��}�v�ڗ�{�� �亥s�j9u���bvwvr˺�9�rO�}�b�;��:H	�0c�j/7`9�[x����.�W�~�i�7�W*	�n���m���(���l�	������LE��m�sU�1q�/_ v;Q:˷'2���z#/N;���Nr7׮_{�|F�+�D��������go��|��zA��W	��^H�"��I���{�Ďz����_+>�:�����@z��^�����B����2�y�ob$yǻ��X��fμM#ؐ���)�.άW�)��$��=�Ki�Ȼ��7���NU�8�2;��^�{��g63�y�%��@����^>8���2�糼�LY���32�>txވ=:��^y1�=���	�>�v�^˨�^Y�mOq���|���<���֑u�q�.��k��$���=4TX��O�珗�#�A�[b^��j�N����Rś�y�bk�#x%�E'x�Z-�PKڦ�\V:Ak��v��'x����M>���P�����a�Ʉb���]��q��aܹ��x����{���#+�?$@q��g,��p������;FV�y�'��b�8v��w&�KJ�#mNg�{w*睝�C���l�tr"/y�Ԥ�3�<`�؏l�K�̝�{����Ih�N�^e��ӯϳ��`�~4���H�A#B!C{j��w:7;I�En���b3�@�(�3��'ޏފw�o��j��W�׹��,���T{�����Pzw�	ї��>B��JgQ(n��'��CE����n��������#�8�^�zI�۠�x�%ZD�G��@�a<�M�١��u� c�A���oT���׻��l^�=�_{��㔍/�w�G�ۿ{:���\b?F���|p_	��d%�p�Q���SñL��=ݷ�"=Cu���������*^u���2ۍ��Z� �uV��t�pTP=sN4o����X�Os�����eT�ó˂��>������w
��N"�����2>Ỉ�U�U�ּz7,�|,�,U,���Y��,~×7��ƅ�kE\1��ΜF�� W3;�v<[��y�"+��$b?xGr/ �4�f����h�n%�k�n�<Q!�#��n�����B'V����=o=��>��鯮�}_Ol˥�zs3ܐ|۽�^�����<���]�µB۾�p�-�@��ӧ��¾]���ڜ����^{�.�mGٽ�a�i�܁���v7���{�X׹���;b#vPpF���r�w4��gP;�<���{�yվs�yɥ���t=0���^����dV�ڹ�x"�E9;[������P���+@�%GD��G�u�9s���r����ڇ%��nG�������^G���ۖ��b�NtQ��W�>L�,D�8j7w�=���y�~-e�6Fyog)�*�Ǖ]�׉�3����b7+K�=���wg<g��-�x��7M��=��>;��z�w�����S�k(�X�O�<��tE�t��C�I���z��"n��޾lN�����<o_5����Lrr�N6՝��>���ڪy�ny`y=�p3��^R^�1�ջ��=�<�����g��K�����������J�{��`����[7�7{�Ğ�/�kr�P�{���2�
�S��g�^���۶��>Dl-0{�~�f-Օ����{�nm'XQ4i=s}�jg��;���_j�OW�k�'k����|�]��+�����X����a��VC���8ߓ3�r^�p"��[�˓�Yϭ���#�Ail�{ԟt:arZ}�O�g;�l9W�Ļ���eK
\w��3��[� {�h��K(�Ù�xx6�6��x���d�?
G�'����3��>�t��noS�s�@V�"��`�ܞ��Uo��,���^��17��T�|J݄.��3xn���ǈ��S�
Ag���٣�Џ{!(I���ί�ɶ�I�j�Z��ȕ9g��𭃰$0F�pod�l�4L͛��8��kɚ��C����f�F9v���gs�%��Y�{۾�\n�z�w�/L��{o�Dk���es]�� �STg���ۮN��޽�/s���p��2�鳯��Ǡ���{��f�y��N������g˯1�xt�����q=#�$�}�eg�c4��K�-��x<�;~���o|�Z/���"��'+n�խ}1��rd�
tH����s�(>߅��ڞ��샼�yf�ձ>Ma���?#��E
������E��Ws�ӓ�ItV�o��fȼ�덾�(>�/%�y���)�B/s6�]�A�`H�
ڹ,`b{![£�i�$ÏJ��Z������a���n{��'Lx�m7Ӽq��\���\���0Rzn]`��v�ʾ@N�=!�����7F����C�a�����9
���7Ӟz�.�0��n��>���{ݽ����=��47���ծ�5���o���}��C����Qoc�;7o-]�̾{���w�ڪ�}��R���c�>�t�jf���9�^��@�ê�v�ّ�ql��7H�s��y�n��Ӏ¸� 'I[8�w�w�A�w�zL��p��b��H���'����w�`>�ǀ��q��{��=^�-)<:y�i�̜V�Ǜ������7iԜ��z���$�z�~���^!s�|�����v@��E<�=^��e�:����7���y���~J9��פ�/v��ۅ\�wۇ�X�퉽�툿#�qrH��%��������zy(	�O�r�Vѹ9烜r$��'cT���rm��C�sG���w?p�yNd�;1��b�
F7�H�A}�Eq
��P�)0ʼ�ў[���tp���4Q���r9X2�D"ƈ������%VFf���|�����w�=u��\9�*��v��m��SS9�-j	����������}'��b.gr�v��]Wk3�;��z�#�V�h���!E^�^���N:w7I���W;Bs汽j����nn�L�#ۇ��K�7vsG��45��;Q8�s��۹�����Χ\3�ӭs���v������ ۸�;P�;[<�;�OG�cvd�=t�R�.�Yj6Z�8�vB�`�v#��}ab��:{S��|�B=ta�4�g�xd���#h-�NX�*����^I]\f1`s��������=h��wW�v��l�,���훝�9'&���4=;2�AGs7��^9nǷ$lr���u<���{���8'n�x0�����x�j�������n��B��i��Zv���Y�rx-�q��j|�i��<U��"�/N��v7.-�k:<n��=5��d��t�vy�#�a���h��ڞ#��g�1�R��v��ey�p��m����&����w��;[`���pv����pu�ݞţ>��s\;q�ٸ�]v�V��T�+��`�6����'kv��=��*��J^;�E��ˣu����%	��G �;�n|�v�Ƌ��1mqiғ<�p�ˋ�H��d8�y(c�^�]���۱�q��) 9�[{v��"Z��M�x�����n�W]�L]����t���ָ�80�O*��j�RCwU�ќj	����5����m����붒۶��X�*��;m���ny�`�n��'f����'X��G`��[JQ�WCu�]�\�۱��Z����k|[���Wb@�cUm�][�<�ȶr�m����ƫV�:{Tp�=:����.�.���w�kt�C��<�v�q�q�.�r^q�cq��9:"��Iz �v�ӹ�k6,񷞍oM������GZ�̯�rf;t�҇��̭޸�f�`�v�ռ#���g7m&KK�:��l<������]�rO]Q8{�p��D-��T������&�>���::,F@�vGf�� d��G��;;�}c/�i�E�n�s�Sv�,J�S�]��{%N��΍��`^e��px��1�}�`Q��N�k�Qi���d�!{�Uyy}�K�9��oj�e8ƪ=6N�Բ��r^z���G8�v{;���l@kv�G�s�:�t��\�dn �1^yn�cJx�7)��G4q�m�s�1g)f����m7Ks�nӆ��q��=��v�.����[��81���r<�����η��n#����[	��)vю��ؒ��۴�8�7C5x��fĺ���v���ܽ���v��q��\�a���v{kv�;�M�vn��c>�^�-cZ\��z����)m���n9j�^Kls�#�.gk0��㤸qu�ְ�c�ŞA=��:|7-�g&MѷG�8�Ӻ��d��A�/\�Eۍ���#���vLj��\�^���"�'�xݘ���_���5ԝ�"U�qd�n���v�t�v��k�!�p�p�۞�"�73˺:�ç��P���\�X������u���se�F�Z����D�N��m�+gʦ�.�N.q͇nH��6�;\���g.͓����[ �[����Ǭ����֝��v�=l��ѷb�=�GyTponn�z�=�\ǜm٦HǄ�Y�OV��z��v�I��vN���ɬx�R󞸚,@Xpn��m*�s��vt���s��h�l�C�k�m�����q\��}���Nl':K��3�t�9MI�����2�\ۉi�uO=6�<�����O��Pv��%}t�[Z���ú�H�"ݸ��λfDgc�����ͱ'v�R9��m9z�f���d�u�J�=�ǂ�Onn����gpv�wN�;8�8wm�&{V"�u�R뵸�](s�K�F.�h�����ݮv�m�i��^�`:��J<Ce7 ���(�q�ݍ[Rٮ,����3^���ݚN���J����ז���"\���Ǎ��Z��Wa��[��ػG�4v�^^�n����ol.!�cz���sA�b�t�Z��\��sΌ�c�u������۸9�Ŷ�#�G�)��\v}�نǵl��nwn;J�hE�tf���ٙ���ٱ��XՆ�Suu;I͒�d�����;z�du�s��t�s��P�g���r��kN�gL���k98���s{0p8ݸ�]��[K�yx��4�h]�Mۭ���xˋ�'u;;���g���w#��n�\���jvz����<k�{9�O;Ov���vR��y65e۶�/j�;tci����+���9��t[�kv�+��X�i�c��P�N.u�!���-.��V6�{2���Z̧]�덃�&��d֕3��K��ۍ]�[�O�ra�v6���bvx�s��n^2��[p�κX�ch^�ۈ�� �/^��6N8Y�ݎ���w�m{�lk7.'Y]R�Y19^@s��fÝu��۷n]�I��L�۴�c��<k;�m���9'X;��7X��j6���ps=��A�O��ݺǙ}�2����&���z�ݺL\i7���o�;�/k���;�ق;4��4U��ݡчt/��;��e����OZν�b�8Й�vw���q�����6���k����y9|��C�^�K��#И�4*v0�
�1me)���s��oCn���O:
n:3r��u�vw6���飞Gm����=��D;vnsk��@�/=j��ͭ�zܛp�{<<>VUxR������!mu�5/F׉�\b��.�H�Otn�e��⮑���;)���8�]>�I���8�놦(��jv�%��g&8��sy�h巆�6(�C�f�{gh��,�<I���Fۋx೻.�ۗ���Y��L-=�^sm��X��0����p�n:y%a�^���u�C��Z��^1�UM��-�Qhܙ�.��]�lRx#M�R.)�뎁Ŋc	�K��G���k�y4V�s����t\��g]�;��y�e��p�#��cu�n:����[���h9�fF�d��ѹ U-�'�;i^.`�9v��w(�nӂ�ò��Wb ���t�ɧ�q�8�uX�m��ݹ����psa˻In2�"r�]����(�5���nx���<G`�Om�Y�6z�X�.2�4�����`{�9�.L�ݓc�c]���.��lc{�O=�O㜞�rob	�m�,�L$�d넱ۛ�d�i6I�{i�*Lv=y6�]=Uτ���\���e.��=k�n�,jr�W0ju��:BÖ5�=�cFrxܡ�7OhDW=�q&��;׳�Oc�GQ�l�)��#���.�n����l��^.�n�n���[{a���/b<ج]��p{;x\�7n�q��b^���z}�6Ƕ�����@��-�a챳��c6����)\T]j���$��qˬ�ݶ7<A�{���Xް*\ю�k,F%��z�u��3�nh�.Mk�Y��ͱ��F���Xn�u\�ػ*Z��{{j�X6��\��|�cph�G2�V�8��#�����pQ)�d��v�Y��9�޵��F;t���n����X�u�T�1����#�B٘<�Dlr������s�s����c����r���^��=G<uB7M��7T�,C;���-�; ���6��f�;�q��u�����k��*^(.8�rF���3���u>��zݺ>����Lf5�N�j��O.ϵ5j75��nq���m���ѷW39�耙@Λ���㍈�&���m��gs�vݸ'��굺�v)�1D�����j�؎*�m��c���a��t��q��.��{[�#�i�z���wo9�Uz�������+�Ep��xJO[H<݈�N��Iʯ.�
�^Ѡ�9���N�l1�m��svX=��T��y-nS��7�y�/vN����ǏImmi��xS��wY��t=�������q7Fz��mi�խ'i�nʵj�mݹZ�ux��S�f���v9pl�3�k)��u��{;��E%�ɐ�N�v��j�u��^q��n-�ݷ��ݺ^|�lH^ ��v�s.�ҧ��q�j�=x�zW�4]v%�Qz����m��<�j�.�\�2&�랟V䱒�n��\�[��F:;����snp���1�ݹ4�C���ݣ[c��;�ۍ��v�vhy�<T��x��2�.x����N5��٧vs�7� �I�uǄnp!P��n����$�&m�7��S%�j#��m�ps�7�GU�퇳ٌ���mhۋqi�s�s�����]���'u�v�m��`^¸v컫��}jxG��׋p�܌\�x��2q�m�4ݷ^Ķ5�/g�����ù��Y���-rXփb�0&u�S���ϟm��F���٪��L
u�r���jZ�^x ��6�<Ɠ��#�Z���M]���p���j�s�vgs:��HY�۞K�Ge�}��s��44m@�1��Vծz��[Ac�v�j�ۯ\�v�t�\趥oY$8��ˈ:mն��s���z=m���;n2c������=��oL���p������7�ٚ��q��R��n�tk�����9�M�;;��.��Brq���u�r�3�ֵ\��L���N0�#u�Yd�O!��n��]]b��Otg3�^�ֶ^^���^i�v{so�s�&eܓ��ܼđAt\�k�΃�Ọm�ț�s����vv�_Cq@���Q�<݁W�]❎�N�lWm�VNl^A�H���㧶zM�A�r�Wa��۝۪�����(GI�m��g����ܜԽo��\J�cOO�"{]��p<�݁m�>��ܘ�v��0n�N�n����.�=�\ǎ4n�ד����+�y{�l�[��n؄�$��M���R��G�]z��v9-���b�������[���kV�an��좈��m��� ���cUVұV$[j�*UE���Ҷ�R�H�@Z�b�5�Q �(�IYeJ1��c���F,Deh�1+eeD��E1QAձUT�,U�iE�U�UTeF�`����TF(��A�6����b��Ȉ#�-���(����b���*��#mQb�UF0�+T�D[j)l��+
�Bԣ-
"ʅҨ�`����ac*����mV#hڋUAV#lZ��E�Z*Ԡ�)P�dV$UPV6�X���V�"*� �Q����( �"*�R�J�Q�,Y
�e�("��"*�
(����-(�m�mm���U����YhV�#hU�1m�E#Z�U���KJ��V ���X�j�����E�j�+lQU�#X��ET�*��%��TTADEEXԪ�U�E��D+dF"����F�҈�S�ݶ��{־[��`m�:�m�	��"��#���A�n:l�	����p��n�ܶ��X�F}��g3�8v��r���f�le���z��Q��й��8M�lG\���v.2��q�� �[���n:wv�[�vֺ$����`5��ynwk6WX�2:���:(��%����kNsm�T{��n������v����P���n��!���;��;=M8xM��������cG����0�����&��:��/���L������6�ŀtA���wbsd��V��U)u�]���|�[�����۴p�B(� 'c<m���nӮ�vR�'N�I�|����ӝP�o�o��C�l*p�2�w�î6�|=��ܽ�62��n���[�78�n��>�zy��ϝ�6����H$m����ӱ��7o+�2�֜;�c��]�Y�`����Zn�ۦ܅�9�����aϲ��7lv���f��#�90ܜ'n���V�ں�'��b6x5�og�a�����^�g7XkOlz��x,-��ۘ����\û]s�4��ᵺܮ�ɾ@�)s�s������}o=��Pe�Ƀ;���\�cv���vvy� s�(kP!�i��1�R�����[��6ѳۊn˭�\vu����ۮ����ۗ���z9�k��k��0���nW���Z�z���s�`Ɲ�:㗶OKۮx8{m�9�V���k'��":��w�(v�	��sruv�K1�n��=�����E�p���p�2�ƼJ�n�S����zW!	Ԛ�';O�vŵ�b�5��5����;+��rp�dKuc�2��C�\ഽ�����DWNEy��Ox��:�����>x䞫���w\W��;Qu�M����F��=��:�T��H�ܘ�gwc��n����f�R$M3gpvy��-��{�n.;,c��u��y����{b���|�O����q��ƒ�7�U)�{���>�-��y6y�_��x{m��������N�}����
��»�^x]���gWn-�c.\
�pP�6��˕�s����Twlw�����]�<���`J�0���"��q�Ts1y81�}�v;xNC<+�m��L��+���*�Vb2�2.&�< ��۔݇�ܟ�_l�rv�.x9N�_"�\c����x�ߧ������>�*�����K�@"7*i<��m�9����Ʉ����\��Q�"��1���8r贎�W����}���o�ΰ""��P�}�� ���r��:u�W�}�/lE�r1L���s6�˝����N,8��Ḙ߉�܍@ �l���>�v���L�)l&�,ɇ_�8�H�����W��M1L�����e�H�v�5�`Q�`�b��#};4�Sl5�r}&i%%��W1�� �M����$���)�N�;�/!�G��u
�����-�oh�՛M�h�q[��*�[G�wNnƼx�M��{���58�}����6e8�w��".'3�{R�h�;�I2 ,{�� �'gfĿ�%�K��w����ǘ�p�K�V�w�v����<��wƍ��.�i"��������ͲU��(��5yyckaLy0qn)��w_�'ܛ��,{�� ����K����tq^?�\dƅ+�4SLp��gG��j����w:��Ve_h�3�f�� 	G<˫@ ;��#�!�9�L��jsా����:�7�߁c�����Ow:�� 2vš7��k%��l$����J_8������%�ZD��@|�!�3v�s�1aY��
'����}��� ��;b|�h�sd��L�`È�Ey�D,kM�ڲQ�]�.�ק7�pGN���Fy��W}��o���$r����[�v���V�@ ����؉Jfs���7�PU�����@;]�Z��A!�D��A�뙠�n23�t�g����	��Qh��$�u�d�Y��/��.���M$�#�`���C�J�m۪	$��=�L@.��ޜ�8�%���4l������b���o_1���|�s��"�]��B�QTH�H���;O-��v�*�4mkۻqr�y$�W9��6�"N�I���#'S�d�#���]wT#�/���� �����>���|�@}���,�A�/خ% �w���Nu\h�B�J)�!���`$SΚ�M�Gk�]�y�$-�MI�P��L�y�5���wA4���\S�d��I���*'�7F�Ѷz��7;����B'��3+�s#L��T溈�D�ɖI+ǞuM%�8��a��[U��$I&c�4�]fU�aBM�ߓ��N���.�˾���P�$���>9�]X�zX5w=Y�T�����$ `ԎTL݄x�L ?eZ� A�j����鱓��0�A'��ɐ N�]Xdf�8�R�je��g{��x�#�����*b�>��ʚ	/$^�9�aܭf��+έd��>�B$R�1�-K{����/y�31z%X�Y�t�{+d�j�����G3v�bBl�NOM��;;352�+u�z"��$�9�K����j,���*��H ~�u`g�V��[8C�"�f$ ;�u` ����=�@����@��^X�M|�X�,4�m�G]���cn���64��m�k�Vxg{�������63xjf�E��"+�Sy�Q` �oUŠ�qP`W����5�A�>dE N�]Z�s2�6D��5i���Z	ێwex�sh"�w]X �;���@���X�K���W�)\��~����]�`	��V:}ѓMπ�κ���N�;��V�H@�����Au��v��Bʻ�� Of�ń@�����������6z�k�/r�p��Cdt�_U��%�W�D�T�Qf/-e�#{�h$|;��� 't�\Y5*=�OQ�`#a>���?m�o���o}��H������_�.��M��\�!�� ����隃�D3�s������Dn6�ݞ'�����-g<�[�*p�$�N�GG0n�sS�	���XF(���r� v��Gm]c��O��p|�ݨ�s��\v��#]w����r�ha$�g�l�)v�t�h��NAz-�v7��2�vx�؛4�l�ѻ�厭���n�3� 3���F�ŉ�m���v^�re��;��i��{'..���-��������6�zt�p]�;n��'B�izwU��mX�d��0�!�ج688I�`��=���뿬>��g:� '3�3��L숫*_L�H���tO%�eBD��jq��6�ױ�L#<Ok^�UQi �S��qh 	��k�@7"��ߧ]���RY8���j���DDD�{[>@�����ܑ��U� ���ݠ������"f%66�ؽ}�1-Nd�\,7�_�Մ@�g�f� (�2��o�\�݈h��;��7�eC��f��ꈐ�";2j��Z�^�i]ˉ/ٻ�qh97f� @�{��1�W�����>����m9U��v��9��]��g�������-�������z��f��S�I�W��I%{e�*�1��y�t_Ǫ��"-��Κ`��Fjd�6!�R��u^������"��g��9(H���9��Ng�G
���f�j�5�O�#=8�^X��T�a�=ç�̸KY����32�eܬ���g�r��4�|���v ��ɖ߷�\��=�#�&
/��iE	����A�	�Ϋ�|׫�K�	���,�{n- nM2������+���VR���N*���uj�:���䃏@Xg�&�N޷ �ռ��Ì� �v�����I�Hi
�R�*D�-�;��ޭV":�]XR�u�<��@}s5�4�@(�ܺ�� H��ra;������M��x�h�H,/�'s��Uu�a�lu�(�8���p�v�����}��
d�'	2E�l�d�#�&Mx$�K�w���Vm,؁\D�zF��4� +�l$�4������'��{p�)z��NNz��+�� X��;����/�s�Ly�mM���J��Ԏ�6���߽w�@ ~�uh �V{�j�Z�]�8�������������ƌ�q�g	�~<2o��y�K��s!J-�����f��2�Q�ݭ���*b�ʺS�d<-q1�Hj}�� �y�G.��p�L?�[s59�X_R*������� ��u8������DNٹ�%�z�����v?T�� Nm��7���� �e&�꯲�Uu[�^��wn���v����N٤�S2�ria�P���e<�-���!�́ZJ<p�w�9��#�>��:ȡ��N���I&�o���w@y��� I����y��b͕����w� y��-R��&Hs1e�)0�O�ߛ?�y˯�X%	&ߴ��(z��Ѡ�%��L���poTV��F��]����s/͆Ke���vꇒ$���A&���c=�.v����|A�;bA l��d�j}�Uu9+�NON�{*�^U�9O�,��6_mK���ڕ֠\̶+y+�����K�������J���O*�'"V�*&D(ۓӖcw�D�ۺ��ôɺv1d-���ɑ�1�.I�2��m(/�N*�4]t�|O�K�"��]��њ���=R'�����H=/����03(a����ڹ�\���k��V��uEэ��p{����)����$�4��6"4��aC~�q���~���$��ڠp���
o^ g�� �
��I�Y�6�#6��*����H���4.�Qkk�@'Ы:���T
��{��z��w�)��� �|l�ܲ	=/2h�A���,,���a^����=#��Ur�f���e��0��[�=�;g �j�Y� Լ���=ʛ��[��"	�����>�:41	��-���U]
�����MR�g!C�����H5/r�ĒWw9(���%A��5�r�R�EbkpK� �^�p�2%�[��z�$7�}�w��:���/}�B����>bM켹Glo��߻ߡ��aQ+c�5wK']��볲��](&@Zz��q��5�K�Z��-�=w<\az8��/<FI��d��y|�Z3ś�{���bc�5Ճz��l$Kٺ��`����L��<�m���k���a��I��g�n�F�7���`נ#��V�<��m8��;�K�{�녵�-�a�7]��[q��8�`�L�y6�.����^֝���q�Ɔ��JOF���,K�aqk��7<��MB&pwM��,�i�q�],�I�}�^$�GGt��X���cQV�u@���5�Hq�"$��aCb5&_s�|R�q���y�A>$t��|H;�O��[af��\F�q��p˳h4ay�q�T�uP ���$�(D�Ec���ǝ��'��%�U|F�s��%��b�7���H���I9����*���z��ą.����6�g2��e��0�vM< �O�7},�e�հb��� ��r�� ����A)glI��ל{����\Dy��$((7���l惖�-�>�qIy�c$]��c�����]�ߏ�\�L��Mw]UР	7�A$��vĘ�w\^��ں�I9�I�TK�7��륐h��E��3�Mks�g�]���L��Ƿ7��������`��&�<�?� �Y�f�����[vw��,˅�:�;�R�귒s�Nù�A�fϤs�$v�fLݜ��ol��DI4�&�0ԙ{�I%����"3������A�#u� ��vă��ɲх曏D�s}�l����P	1N\��HJ�"@$���YAU��j��|?z�����I�)4{n|� ��ɣ��u��On���ޙ	'�n�	'�/��X+��.귤��D���H���RA�AA����;u����c�,������;&ʍ����uz��f߁ޫbI(��I ��j��ҹ=�#��u��Y�$�b40�)�[	���ꏎ�_teL�M���$		flH$��TI��ٗX�dY��>跄���a�L��u^2]t�	�}�@�hU���+�/��*��a�n`�Q�����y��:�Mi���������D�1���I��n�r�.z�xY�M$j����������'=�ӽ����ꏼtN�S��y��C>��7���<�8q^��y�:������}�{�K�ݨn�ɫ�1X�`^C����oo��}��kC��9���@�!}�P��O|�^=�j�M�{ٱ�5���q���^[�A��]k��.OB;=�	仹H��s��nëh��a�o^���s�HI�;N�XB�������t���]�8��FjZ����74�KR_QW�Э�XbFDSt�6 (8,�պ���s�z�ܝ7�b�G��<��cy�у�oK���������Rr�>a��q=�w�9|��o�хںŵBx�{�ڳj)ȝ&����F�v�����q���x���٭`��=f-�|=�ޙ�A�����ߦ.Tf��"��[���Z��촵���[*�pl�����젢��f3=�g�7sw�ցwm��>���&��zPW���1�ˀ����qay�(�o?=�ķWc���E��V>%�N{s��ve�`\<\K�y��������_�ѷ���?j��x�ޒ=��wiZ� �(�rѩx�L�;c�wP��[P�|X����}����?,�5��dh�c�ܞ�j<�'U K��{¢ov�S�?@dMn�C K4ӆс��JLنl:6��w{������C��]������������ʑ4�o]�^��g�z{]K;i�|c^�-u���gw���h�PH��b"�"�i*�#lQ�j���Q�mb �*"���J�mj1E�*�X�b��hX�Kh��5��RŴ�-��@���m�ȶ�`�R����2ڋ�P��+Uh�ѩ[�ږ�ȰEBҫ-�i*�P�V�*��Eb��F �(�ciF�R* �1����ĩFժ��Z(�mұ��؅���H����DQX��)R�mA[lQlDamR�J�*�Qem-[BҠ��VҪ(1���Ɣ���-j"$KF�R�QJ�*�TE1��ImU[lUX�A��b��֫X���hUEDAAb��6�UAU�"*���T�E�"�(�"�F�h�kX�%cb�UX��1(��DD���R���F5��Qb+AQF�+Z���"�����UX���b�",E�X�"����j�ƭ�حeKe+*�,���*֭��%)eEkX"���֫U�elg9��		m�O�$>}�.P��a&�0Հg��s028�\ނ �̳�A!�ͪ�s�vݦ�i8� �*;b|xV�6Z0�[k�-���A�z�ƽKk�Өf��Ē	��
������2����O(3���q
 `��`���G8�ض
���8�-�[�9�6��~��~��]���� �ι�=y�^$�7�H��nֻ�zQF _9tAv�j����o͈-4��T{*ܒpegB̴B�9 �珶���rA ����T�l8w�g�D�S�:8� 4�d�jE�U�x��s�H��;�C�ڈő\���MA��b|�o�Ɇ�2�mלO��z�L�D
�b�vEx�H�Α$�
���
ۻ�OVZ�A��݈ ��m�9sq{&�w[Fm9���1�kk�{��
���KO�[���b���ݵ�`��q���O0��\�2��M�a�2�\�I-���C"<֐8$���"A �^� �
�� �!�w���}}K���}��^�֮�9�9����vqu��.�:v��C`�P�!�&��ф	m�9�3��^$A��r	$����+v�/T#��@��ڢA&�9ω�
�\�A.!�""@"��@�����S�=;�I;�I ����E�r69���}�֋�.<؆��L:�{.܂|	�
�I$�×x'u�p�w<A���s�	 ��bv0� 4�d�jo���D�zv��VH3N܂�� �Hz�h:�S��o��� �oK��b�i4�DU.��$O�k����S�sUU���O���$����	S˙���O�\�B�Cy[�f�'K�7b����u?`�z�&��G0�]�_{�]��=����y�� ���-��l�qq��}�ۄ^,�	��nS��Uy�1"��wd݆�91����`K�nP�ȶ]��n�q1��}�=y�
���sT��y�6ʺŇ��h,���z���ƣ[z�gnN\���K�a�2GgX��sy�:�D��rY�G����MX$��m�$���X|�y����qT��a���7]p݋�w�?�|��|,ɝ�	�xθ�
��N����)�y���ӌm]� �0nQ ��AGv�K�.	��_x��s�I!wd� �}�@�TR9y��$���A
���F��
�F%���&o����c*�0��n<$�
��>'ć�������´���]���r�X]����4H��Eg\�A�̚�H�+M�ڲj�OU:	���rA���T�s�����d�������Ư���ԖT	$���I)�ȠGGs��x�����$��9;l@�e2`�5�WTH���$�Q���{���� [��$�����\Ks��o��$�2�kq�q]��Z���m���bɺ�ؼ[H���k����-Â�q<D��� �b�l� OGt��b�n0�x�k�}�Ē"��Q	�JHjE�����rI��%a����[T���X�^���x`P��#0�W(;�*�Ӭ>��tjLO�R���>b��Z�M9�}fR�T\�vu��I�1���67���r�8Tz9ߍ
�
�F%���3}�D�����>$��w�ۦ�Ă���I�|�Ĉ
���N$Dz��MĊ����w ��̚� ���@�^��c�7��>�yuD�V�.<�m�t:2���[)L�'n��@$\��
$�>s���k�=�"�c����r�(��.%7n!8מ�'JJ뭵ָJ�p=�K��(�Bh6!���V��@-w�*���H9���$����P0���~6DwN	��xV��ӂ[j"��u��n�e���N�N�|O��}"I'�w��/3��7:�I�]����BRYPZ1ړι�$D�d�$�ܲ���D���ږ�)��R"N����,́w}
E�:�?=�kK��Kkd�7r�r�z;�9Ǉ'11\��.Nfތy~����O�#���k�OQ�n�MǝP7�N�,�l�t�	'�ψ>${�I����c��v��$����X1T�E8h�$^m̒|_<ɯ
oi�T�ٍS�A"y��A%��	���C���W;k�������%08�n'��㍱ѻ6��n'׷��ŵ�'4�y��K���]�o��$�ޱ>�}�^555Ք3�ˠT�?H'������A�YPS}ut(�Mw
��f��K�I$��� �Ϻ�Xxν�Cj3ky��1A��pKmDM.�d��]>�A%:g$�dk����đ��ĂC��^<�L���b%�f'y�/*.n�=1�H�{>@'���ܡ@��y�邲�n6=
�ʈ?��=|�aw��(�tz6���x�"V�".cV3uz��l�p=I�����N��������U�{f����'��|�G�kLE�P�i�󪙽�I_f�2��ȃ�Z��NۢLgc�|K�yTI �o0Ѝ�CQ��;O?1,���&���;5�NOm�v;V�|�1��[��	&��n�i�A2�pX"#���I$�y�@�A�ꕊŲ/*���[�H'���P&�_ipa��e��6�Ān�5X�q]�|O����z7���O'7�lgF4Ve���jjlA&�y���f�F�̪�vv���|K��TAcy���b�-2�ۈ�7<hL�.-���$�w�D�A=��H$[��P�T���=�9��B�WHJK(C&!�[Rgg\�K;�>s:���0���H{yTH#y�$������U�V�!�۸v�wOvzg%�rw��<��V��R�sE�̫�rN5��y�&i��w�r�M��*Mf��]ɭx�����������V^�ǯ���{<X�vd����t���B^m�[6����,�����V��m�n��᭯c0J�ۂ|���j.�u�����l��plދ"]�Qٽ���;��x���b��1Ӯ�#˸y�v����Sf��q��6�u��{2�-t�Xx����96��.\�/��s[;�E]�.��<zK:yC����wj:�Dp��v��ɖ#�gXӐ�x�9��A�g��u�s�%֐%�?�pa�1AP�ny��� �ǮA �O��ؐk�,�;VS.�����L�ТM��$��j- ���l�\�1�0"gVOk}7�I$gNȒA>k;bA%]uټrս���X��=����!�Ty� �Y��d�T�a��˪�$�o'\�Ik3�H�����T̎˻�%�L��&�y�� �!vlI$���Y�S��K2� g���0�Z�.��L�����
W]u#�LU�S�ĂI�,��>$>��'��ѵpi�H�9�,�@�7�{V��K���6�c/���=ób]�������c���2b%��1=�O�0r�C>$ӽ"�3k�ݬ��7)���|J]�=�(�e��Ϧ��H`���i_����֞N�~��Z�(K%#�i t[�|/��{��vM��oI뾗}�sE.X��>�좏�Q.�EꚘ'RXo�{����$|�gD�	�ߪ��ى9U�g1Tn��̌)BE���h�t��ә4A �!n#���#6�� �������k/�b�"�7].s$w9��d�1=,�Iw9�D�
��6,J�SBH�.�$�cQ�"�T��MM�IW��ǳ��ױ'J����Ă�NuP$����:a�b�$)��K��H�HN&�нD�R���	�)��pĮ�vŭ"��w�}�����AM��L��g����٠I$�wH�cB������J++�I.�v���z$%�!��-�2���p�1�3��F���گA'��ψ'bnn3���t]�x6�q��(�-�u^���H#�uω$����rp�o��<L�*���s{��8�L�����j�n{�ܜG'�߬��.g\`�/=�ut��Y�~��޹�Ѿ����^�z>�>,XWq�.DI��|!~�i��KH��ɠH'āq�"I������㌍�3�SJ��3R*�3�Xl%C@˗$��Q���2�M��m*$N��I��s��	ol{,�|rU,vc��J
,6A*6������뭝E�tνu݊Y����m�N�����#�E�m(%��u��I�u�$|	K{bM��nb�==޿�Ϊ'�dw9'�j�A�L��j*����%td,�`sG'^��ǣ5����s�A#�f
��t�F�'9��z$%���-�㵋���� ��k#'oq�v�/��H7��B�� ��V�.
0iǝW�M��w.��,@}�t �lI$���s�I_mv�Z�]���R��	x�ĕ��o�<#vH8�ޞM��f�w0q�}�w}c�;����h�7=�qm���A����65�}��{���=y�ŏ��	d�, �޹|I<ɠE����r��Q3Ւ$A[x�K��^��sĮ<����"N�v���F����{uZ��E���������}��-�
������U{>�	�z�f�ǻz"jݱ��`IW��P5�.iA,Ⱦ���Iq"�F��=��c�I �ݮA �=}�DI�9g=_��U���|��Y��i��6�W��vH.�l���b��ݙwy#	$y�|A�mP#�ARYB�;�oJ��j�ڬ��������Q�حE�)Ǟ��i���[�04םP��ڠO�'�u�������݂#�\�K�}B� �w92 �<�W����Ѽ�{
E�z�ܛ[�o\L��3�gd!6I�n6j��m{nw%�`g7uj1BL\����O�!�����cx}�c����w2v�ɞh`c# k8x�2������c��߇���ܻ�O0��a3w� k�+ʹa���]�%��8�A�o�{K߃��������>���<�/�@`����g�@�Ҏ��J��y����;�{V��	�o����3|T�ȷ�N����ǻ�y��`]��sf�tv���Kw ]�G��Ƙ���4o���E���g��D���Q��Sa^�)L�
k.J�(��,mݷ=�Ѧ��{<��<,�ԝ�d"x����5�{%���Gi#�{~�c}���uӻ��y���8�8{̮�ո�g,~��� {|��oax<��y"�с�㫞DM_>ް�0�j��N���a'm]躑n�`��=�`�9t��`�oS���=�̓�n,շ|�	����7;$�
��n��0a��ֱ�7�{���˓����-��F�w��7�eؤ�Kn|o�z��^�1Ҳw�f���������`�؆o�ݭ������;<]s��Lv���E��uJ1g�(��b�ƶ8������Z�|�^���{��[AӾb�}}׽C�1m�Ȅg���3�|�S��7ٴz�g�D�,:��C�rX�P�I #�:�����}=d'h1C�Ǯ|���;u7������oe����Nt�&#2-C(��������DQcTm�J،b�-�Q��i-�j���U���U�e�UDc
�)U�EQ��ȋR�)V("�+**���b �ŕ����Qb��EY[[�֊("�,�DVV���VkX�(ʍ��mlX"��kV(���mEQDkU��X��`�hш֪EEDQb5��V"EZ5m�Z11KakAlh�m��h�*��cmҪ�*Eb#KT��VT[J[QTm�Z%�TPEEQbE*QQm�P�-(�Ŷ�T�(�#FQb��R�-B�QTb �B�V* ���j��EJ�VұEPP����Y-��"**"T���,EA��Q���V�eUQ`�"�EVT-(�"�1��1b��Kb�TT+R*�"AH�h��VE5�إ�DaU�Z�*�c-*ETe�PU��F(�-
 ��V�YUPccK��J����c"��[X����������U�$�$��,L��ĳ���q�^/=�N��F+^�;�=n۝kni�[PlM�v8��mp�0���FY飱n��
ή:��gq�v;v�Gt�1�
Q�����7OY.v�Y�^K�6qۮݵۑ� p�'wm�Byh���Ѻ9\��ݽ������^�֬����uNss��EkٍE�ON7:����-u�z����5���s����ci�a���vs�Y}�N��ꖰ����F�����x�g����ui��y�Jꫛ�6�mj'S��W�
mEyݰv8�%�x;m��u-Sn�>�M�l�ݍe���^!��V��5�V'q{��`����e^S,��n"��!:�P��Z@��:W�nܝ�ܝ�L�݄�cu�t�c��7n;��؈B�c���Z	��Ok�%*P#��m[sٰ�Y�tg�Ϝ.x�1u����a�m��E�n��-�= ��ǒ�=��9��j��rQ�+X^�E��n������Ak�s����������ìKǎW���qY'��ݚx{m����Ʈoa�r���\Nx����9��Z���GW`�N'�����p���[N�G����u���r�lu�c��y�[��<��-́y�Jb��[s=wn�t�N��b�Yl��<��d�ف�ӻol ��x#��6�܏=������/cԶ�'iJ˜��<�:!m��f�J�'*��M��cr�ݱ���j��\�]�x��0�Q���v3�����vF�'�-L��s�gf�s���{c
�C�ma���zOoo\�vb���nۜ��L�+���᫷N���p%����hM��1À/NЩ�zm�v�L.7�s����Wv2�h���;��3�e��/=��c1�[�tj������J� �΢�O`x�h���^Cį�E�ح�Ra���3�-]�%�gh���;Go�����6�w*����l��;59*��Ѯ��;4q!��]��������]�n��(.;��<|7͂a�>�;ۺ���m�۶���ޏn�ܱƄ�飕�;�ѵX�]�۳��e�7gѷo�=��:�=��V��=)�.��<[d{,�<����;�����v48��l���+��c����u=>{#�w#�ڗ�g�����;;n�Y��\�z�i���_8���B3=3���׷�vkY({[t.kq�ӭ �LS���a�X�s�{u���p�pZLf�����O�p��@�Â����'��y��$lwH�o���Ӯ�%�Ϊ�"���l��Uʗ$��ʚ��2��ݐIv謁H$�w9 ��s��;��k�O@�<D���Y�뫪�M�sO��co��e���s��v�W��>=�A<1��Æ`Cm�U3]��蕵���q5S^$�GF�'Ă���RlRFk��oo��r(%� 80�.�{�|H$�L��YY[4����@q��I+{���tf$��w�������얮�9�#s��[�\����[V�u�`[ ��j�.��Ek�z����>$Ѻ�H$��rE����&����������U�$G�a�`��"��D���F`#���{U]M\�Ui1ɾ.hy���;��=ͽst+�պ5E�nt��.]��SӐ��qm�éj�8����L;�t{��u�>��� �s�|Wr�����Y�ܻ�*�_7 ��	AP�W�NK�A���LE�ԍ�9sfWL��s��$��� �:#Ch��3u=u�i��u/N;$D�9$�@Ks�I�!�vT�\�/��W�U��w�}�����8f&�UFMWK �b:�h�Kk��[�$��w:D���ؐA��ڠ{:��U���|N�|<��̀�me�v[��Vi����t�\��;���˧�����߯X�7l�w�����%���A$�Bg!O?w@�;ź�� A!+܉$mJ؈�Q�a���o��A ˣ�2tnI'�v�H$�wl׉-֐��<N\v�X���2.����}�x���|�c�G.j!���w�D�v�%�-����9���o��{_��T|�s��Wj��-7��&�WD��G2#T�bޮ��;�  =�ع<	�}A����5�G[d��	AP�Qv�v��pުF��>d�DF��O�>�Ml�X6�e]�	KW���3@�N��X�D�eŵ8H8^\H�b+v����zn��a��:�>�t�Pӈ����]��Y�n��tu�۶�t�F1n�}�?}��~?�hp��MO5=>d�������;�A[�d��Z��ŋ]7�@$���$����%�bz�<�^�:���]��U�A�̪$��x�:��Z����f٦���?9�og@$�$����'�:f�LF�UH��$1��I	a�a���b;�u�%X.jt	$��>${�"��y���G�f�
׵s�ܛ��|wD���<g/�|�@��wg\��f�.�~�zM�(|��j��{�HB�2L�W�LiN��?���=_~ݿ��$Wu�d��	AP�Q���J7}!�>AP&��]4A##:g��tI[�o������}C��n��;�s��cA؉�ΉѺ�-ѻ�[c�#ֺ�뾾���?���x�êv�$�GFl���w@�wZ����1�}{TH$.3��@�mt`f!��mLѯ�08��,��(շ|�{�g	�>!nk�|Q���cr�j����P4�
	pa�\)"2�D�Q��dc�
���	+����$�KY!0���
�����99��󺹒H$��r"#��lm�;\�Qئ��32*y2Dx�����En���}�Ff�Y���˙u�z�� V�?%��#N*����R���ܹv��d3�Yݧ�Z,d(�QV���.+)n٩��ر.$%�c&�he�3���܇:�[�[׻&��{8i[������w���㿮��	�tmj�Jv��n#�w<`�}'Eq��`�o`X���g�h��;a�W���u�oJ-�B<t[���݌n���Վ]�\z�S �h^���:s�x���n{e�Qz��8q���\�78Q�0\ʋ��k�n;v�������{�{.�ܼi�9������u�]��'c9n�.���[��p[���]�f�hT�Z�z���-�|\���ݵ��7j쮃�.���.{�v/:���������V�]p8���E�L�]��I�$�#���c7����$�y2$��9ωH���6�fET��Aw�:�λ�N�"L=�$��y�1�4|��zvB��:�"�+À��ïL�� ��}5�I ��w�jNb+u_\g���9�$���TtăM���%`�q�t*^38	�]�H"7�*�$����,�>���.d�y�I�R�HL(0�uU��TI>(�l���zV���ܐ�&���D]��x���*F�C��\�0]�.�� �c/ˆ�8g31���6�FC%��vLg$b 2&�^b�L0a�b8��2A&;'&��>$.��&�&�z�8�� H$Gd�Q��:�$6Q6f��}0|vCӂ�̉툫����/��%J���EyxD�'�"kd���]�}V."��[�C�RvrEЌ��p��V�,�Y�u5�{��N�������	$�cvz�|W�~BA�)�˧W�<wa���!�V�h������$�˵	)w���%�ڜ�,ד��o.�
�-��`���&�g8���K��v�vh@$�� ��ϝV�c���,�'��(Zl�l��0�.���@$GvH��r��T[�@��WU@��oH�c����ZF,բ�E�y��H�tK�uع�NNh:������ D�@�dO����q=���i<ﯯz���gLI:��FF;<���=�U�+t�2+%IHL0a�b'�WWO���j�GC��5��w���,� �I��b|psY�F�ܥ4���;���H�Q��t�)�{��>'��&�8��H��s�gz�%5!�Z��,�Ϟ���V�l���}w����Nȭ�ȹf�Ǩ�1�C��\zFz�_G����7��4�A\��<|c��&8Ƙ��C0�eWMM�D-�3O�MF�h$P��$���z;����� v^h'��� �}Ь2��Km��D�T� ��}S@�AJת�]]�i���u�I��pV�0ttP�%�^����ف��a���ۋI!y5���;���H�[�M�M�Jm���lW Aײ$�I;�T
��zo��d$�o9�b��HL(0�u^��ڠH"][���ѝ4�8����$�|cw� .H>��u�e�,:�&����(���0��|���I�%_eM�O]�ꪨ̩s��f��ۮI%ouU+��`bx��jL5��x{���4��w5>�	�veUx�#�8\,*|zL�6{���k}�}���{:hh{�2�;^��W�XQ~�}�y��h�v�诿WQ^�xEˇ.������-��d�K����si�'��i��E�8H&j:jl	1�F�q:$1e�Z��=R�U��׉��{���������n�?��&�����ћ�.�������R9�ut�p펢E�������h���y�"k�dW\��$�V��$��èN�O���U��P'Sf�dD���p��2
��D��ݼ7�P#+����;4O�v�>4�$B�
��^�R:��	��VVuQ �#�Jv��F�}-���g�� �
ݎ3"�B�	�	4J�WO���Ȫ�'Ă�#����x6hB�6�v��������"h�8q@ܸ�@��3�gF��2�'�A��r��E�t�A&:��7�_9�Y��P�'�m�\���Ҟ�[�M��y���`��쀷n��\���T�G:�s=KT
��{݂)1�nb��{�p��X���5���-�kRԦ��Wpc�0���EB�8�c�������S1���9;��;s�[=��gi-]6�=��i����.���ml%���I�#��u�X����c���C�y��]Gkd�<���-�������h��0�ͷ=��<��`zu�a����j�n0awtL\�Mu��'co�g\u�mɄ�]�	�m�2뵫mx��]��ׅn����]m�67=<�GF���y�瑷.��ߝ����nL�����n��$�c���Ji�\��gFDeH�|Vdt�9��pYi�l��&���V��ʃ��a^�T��$����$�ză��*���|P����`'�f�f"�H�Rv�� �Du�g���L
F����ⳣeI��s�F�#��1!���+�:�Ss�!���Tt�I>1��|A�ޞ��:ka@m�z��Lu�du�B|�0�, �H���򾜑s:���ނw�dO�$�����=TB[ǟg&��a�DA��>�3fڽ��6L"�*�c����@���������6��F��Ƹ����ɐA!wOUA�BkP]q��j��59NA���� �b4�a$��HPf�]�A�0���
�%����tVy��lZ0;̍S�unު0�ECֽuf�J�p�A�k��	韟j�(�;h>;�un�T~{� {�v��>$�}�I�+離����l%��\���7��ӄ�.u�;7�>$�=4����&���I&:�� �����N��&�EDp��;��n�r
�\W�Hku>�	�+rz��
��!e�k�q=�}��U9$dR<��	����V�uP$
��(;�ۤ�Y��A �e9�@WӵD�V�?O?ȋk�!3�5�$�����܅ɜc��v��y�ncE��_<=���������Xa��rB���$|Wo1':w6�V�7 �O9� �����>�����
mEP���q���te��I$��W�$��rAN�ՇS�}/M�uG�I1�A�ꩳ�ݮH'��n�y����WC����LR;$�jh wv�[������ǂ�������&ݞF�r��Ւ��/�݃)�^�BO`i��$�'�0��vQ[0.I�G���ryG��`^�7b&.��!Ė�C.���Y5f��x�Z�/k}�Q�=�M\�R7qVn�Y���K�l�GbԨ�*���dĢt#���T�v�w��9�w��W�& }̆���=��a�v��D��	��f��]���n2M��L�G��{�*����,�F�`�w���ٮ.�I�J�wL�\��� �X1E�^!���O���8�����wZ��E�'����'�M{�^[�{H�X���^��`�����;9O ��o�.2��qSڱi>�=��M�!�������:�mB'9�3�)��cLk�;����o/wr��������1Id�{s���h�u��Cz��&#�����z�3뗆�w_���?g	�;�z���]�V<x��coOm����Yh8��r����׌B7hE[�TC����B��6 �����;�I˗����̮����:oϮ���7q����O6����)^轺��\���x�Kr�3��$�9�f)�!d�b�ݜ�������_p`r�˵�Xm�G�|����0�W�I�v�ӽv��p�=��OD1t������J$�|TP{|73f��|'��{.�ճ)��[`�w�Q�}���'�e�`]�sR�aVY�;���ri�2���K-�{�0�9��/A����u�2-�ӗ~S���s����b���E�*��Z���V���X�R���EDb"�TX�-�����TQUA�b֊T���F%��Qc""�EX�UKJ�b"�1�ETA-*
��ւ�A����TQb�b�+`�Z��E��*��1�(�Ŋ�����*���[YDPVDX�(��e�eb(2,X�%J0m�"�JZR��ш�*0U�QV"��*��jX��#Q�2(�X*"�1U�ADDE�UUQ6ʈ��QDX��H�(�*�FEQʉ	[X�E�*�A���PU�F*�B������ ��E�PQEDV*����Ŵ�`��TDX�Z"Ȓ�,DETEPUb*�`�b�V*�dDUmUb����(V�*�Q���E�D+"-h��QAA�`"1(�Ԉ�*��AQF�%j�� �� ���QX��I!�g;��$��O�^$�����9��[�a����m�7�/E�ʚ$�٬H ���v�{*��|+���y�J����N��m� �#��Һ�Bn�/DG]���ݪ$�y�O�1��L�N+�������ﯣ�=��>����;D��e�1�=��T�}M��i��8�(()D�؎�`��D�fv�g�%^s	��� څ��Ļ]<���U@�|U�9De����
=]=��
jn3���v�i��$Wo1$���ω3P�_�81E���5�z��aCm��7=.A$��[�$�i���O��u�4�
���$��by��h���E>����CX�|FFS	 �V^�� �-��ܦ��M;7FjzH���Q�a��0��D�m�?]���o�x�骾�����zn%D�l��&�\ÁRÍ�rg&��r+�=�xO�#��rH�?�q0�ê"��D�H+랚�2�Ef�u(br�N��	� ��rH���`���2�Q�J���c&E���m�����=j��0�]�}N�G�̼���~���BID�iq��bA$-��$�	�ޞ���.yS�;+�^E� �Vg9�R8����?A�םT	�ܡ����@$��$.��I�������1)�LT����0�a�{nw$U����H-�$�*3��O�F�H]��@�u��
a�ۈ���M�o�R�"ϲo��V��
$��{Xr#En�3�n�(9�16��!�����>���J��$J����	3�nI%]���|Wv�4h�����+4S��BXMRO5Q���0X��U���O�Xre�����-�*�Z����i�0ȝ���v'�������{��%���q٭�m�n�:89��s��g���-��G\���f�s�7�k�����n8�n{�$H�����k�a��a��;�r9�۵�v.M��x��1o㤵�\�À�P��ܨk�;n�{/<={b�LS���Kk����Wkm���t����9����q���|=�E�9��`r�q8�=���v��p<M�h��B��v����g���`wg����mP�=���sԤ���F���K���CE�� &���MuL�W\��$��$��]�"v��[�y�$�vɀ6!L$I)`x:����p���I'��V�P�I[��$>"6{3,�m���Ȩ��$��W^uQ$+�s�|H:h8Y!V"ftN�$��]w�G�
�t�)<g�M�u�^9��S�	�
�͚��Wvϧ��W_:Χ���v�$]wm0�
!�"�7ă�[�%9$���2��U
�_��W_9���N&���������G�v���1e�ōn�Zr�l��#[����A3�nv1G!��HPxsۺ�@'�vk	����	�"Y˷}]"�	_k:�����T�ڟI,��,T��s{.�:ؼ�p�����k� ��r{Ɓ��9�IS�.���>}Q���-�Ë���_U�ĮLJ�p:YS��=���}��#�I��d�W��Ij*�i���X�zx��I���2���l�|��@�M�Y#{.�	+28�$��r;�Db�	��P����}C�.:`` �n.Q �J��H%v��F�{�u]��5,D�|z�2@G����Q�� �|F]t�I%_NM����\`^��3/��	7�I$-�� �ۈ����a�����.�6��NM����&��lݔ�;�n۸�ۺ���yk�������E��ZO���=(�EGc�I!wOUxȸ�X�6�̣l�c:*|�'�"��끪0!��EA�}wT	���|9����ƣ1���=TIv[���s0�:��# ���n0m�x�[r�A]s�@�B�3;[�%�����ͪ˗S���:t�����ыBA޸��s����wv�U�n�N\ĒƳ��%��D[����� {�^o� �o�A$�w��D�T1I��$�e��=&X�$��ͷ$�9TI ��ؠS���0yQr����@Ȇ�K�	�V?���gN�%_Fϗh��gm㬇!�y�$��ڢI+{X�3�o6p͞�?�:�p��Ns���V��jӣ��rݗ�\jM
��@D�3.>r7��EȈ"@i�л�g�A%_NM%wl�8xtS�&�7V
N���B���[x7h8l���Tnz\�2'o�E9c+]H]��D�A]��&�w�NyZYs׉��hBN���Q�S`�I]��I���T�'Į��	[��:���P!�ڍ	�<E�Τ�ʚ��y�I$��_7qnz%���K��!;ޤy�엶����x^�-^���~�sH���8������#�U���5�M����YC��Y��� � _�7s�9C����"<�*L}_?IE���\�fb+Q3w9U�A>+�\�	'��ɋ�}W����8��w�?��X�{PzH��5��sA�Ӆv5��#���+�ZAc�2�X��r��h��;�d���D�����$��|���ʍ�&wVueP$�}�I��a�$�a��f���9A��u��w�>�H[�"A$t_9���8�{��:�������SP�UF�dA ��ɒ	;��y�μr���Vdt��'Ǣ����"M�ACc��<m���f��`*-���$���=W��TC��������8r�4[��"uD>�� ��릁�g�<K�zgĒ�x�ĂWuuW�F�f�%+S�>�T.��eFC��;ˣX��1��-��c���)mj(5G'2W��s�1��-	�3���� �a�'�p�i+�34*���Wc�;�hyG �b��F�xp�-��Y����Ʀ��X��q.��u�V]��j��v2a7^�����3���p����eY�Y��#I�Oc�m��x�'fN�n�s=�4�g�2V����L�"�Ɯs�tl�u�L��K�.���-�p��kщ3n5���ø;gf��gf�}V�q��Vݣ4�u�U��f*�t���'N�o!��W/]v��Jn�g����qw������
+��_�]0|Hu��I �oWUY����ܮ��sp$���$��DdA�C$A��Ν��N��ڽ�=7l�H�x�Ē�uW� ��5�ƴ�ʽȃ�4Ϥ;kI@�	&�AD�:o�H ��ɠH$�Qbt�J����׮I%wWP����m�C
�ٞ���������$��Bݞ��$�
;��IDx��|I��rN�mF!�jPf�n��{6CT�X`��&�!�� ��'j�$w�\���� �ߧ�9��==	��B����g���+��ܲ#����0�9��p��M�+ͼ�u�!WN��;�O8.Q�1:��� ��ɠO�0�Ã��T�#�fH;�䪄�t�L�i���s!4ɏ�봬������0��W���}w��.��$�޽� ���o�J�TTh���w*v�^�Vn/��_	 ��g�O�!w�"|�p2sb'i�FƸ���H�37{=�A$+��+��v�鞦�A+r���A{dI��E�$�%GM��ݒ�#_j{��kĂ|W��	=o�	���+W3хx�N����� ��4�P�U�},g��y3k{�Vȳ�Koל�Fx�gL�	=o��k�Yχ�5$��\<ڜ��^��9���<A՞j�]n
�^w;K:q���F4 �M�F�ºn�	>[�ĂO[� ��iq���f�NU	 �ٲ'����I�%y�5��̓t�4v����ۑ����:�@*튵
=���:Xba1�dW�O\�G[�$�TL23�uf�«��O
D��;3A>�-h�j`ˀ�mP��1yiΗA1���ǊwT���^�N�N�+�u�k�{��<<�w��ĂA��D���o��z��.!(d�5U]�[6��8N��>��H$���V��_>+�v�cx�h�d��!�H��$�((�m��뫝73H��9P�Jg I �>rO�[��F
����1��'ɵ����[�?��-q�Ƅ�pn�ĝ]`i��+�ɠ���00Q�1�l��7�7$�m+��d�:�H�	$-�꣰\�M�����0$��H嶌`A��p�#k��enԎ�t]4E��Ⱥ�I5���Wu�׉9m_tƇ�"&��E��6�4�n	^���W$⫯��I'D��9)e�Q�H���|H$.��`@p����2
�ukۧ�\�rl�j��$��
$ݯ_L�G���Q��76ŋ�țy}C�sH[�$�,ʁ�eR��
�����H�s���b���]z�J��e��:�)gr? ޑ� �u9;���6��4*�>� ���r�J���>�$��� �J���D�ݮN�@�[�S�i��.->t<n�f2=��%Ѹ� �M�6W���طC�[p ���D�'��_D(7=���wl�Wq�wH���������5�7|�m����SF��%ElVٻj�p��r�+�� B뼯W���VS��(�J�v滈Xw��B`60�&*�n�Q ��r	$���Uq1z��V��Q��s�GkC�.8Ez�#]�3�������'f�f�|���$�\��yk����X$MuUP�Ɇ&QBA���ֹ�$�\���8d���<b�t�$�}�|A$��r�E�D��8���X�A��l���L)�4�uO�T<}�{yG�"&^��fѡ�̿!����������Ry��|��]��w�	��	�Y^���&q���������X3�S��Ez�|+�=�m�+�um�O݄�ݺ����wpĶ8�o w�*��*�j:j�+z���]�\��A�vz�}�8�hYI�����r�,�DM��پ�7�N�v˹�S�S�٣s�������@X^=y�CvS�rVh�F摚����yl��l���)��S�W�D�g�)�M�"x{���VL�1[�ѽ�`�9�f�P�My�,���b=�!��b�t��Ϳ-eˊ!�Ibꦴ�����x��������r`}��}8`��zaqX��۸+�(M;]3�\��nڙ��[�S��Ftm�w�&И�E�C���=������\�R�����Z�)��k���� u��=*���*�XU{;9J�uwU�gk6j.���bøx��bf�%�_l��v�g*��|��|-�p��Z�rV��$�:>�ܛuep/)���>��M���Y����7wu>�Ӛ9�c����F$��n�pN��r��M�U��GN@؍؃���;k���ۂ7��.�璨�����}Bk��t§=�x�XJG�m�nsQ���	t�a�ۚx~�m��ZT�`���]_3���55l�7kP��)ԙ�;��2��ܜj5l6�24�C��ͧ����:xb\^��c��I��S��|n�nl-�,N�XwzD���w?��9�!�C��u���݅ȋߨ`"+DEbr�TUUQ�TUTV#H�*�ұEV
(�X"(��PTEX�mR�-V1��V���QA ��UEE���"���-,Tb�-�TX�*�ADH�,EQ-�Ŋ
��((��,bł��PA,b��EQPUDU��)��
�+PX��KF,���*���,bUPQV*(�)UPEF"�������(�Z�b����A���,TX�X�DX�"�*���b�1V",QTV�X�� �""��QEE�`�E��R*��V
,QTX���QX�Q�(��EDUDE�X�#��QDE����b���*�QQQb��U`�b((�Q���"��EDEb�UX�b�??:�+��<f�f���ל��/�͋�<sɲkLF]ۮ^�Gv��hs�on��6N
���V��y {(�6��p����QŘ�\pK��.�v}�®��<�A����m�0r���q�<8���U{Aצ��GG<��@h1�Ϗf�[������l6�\u�d��C�d�vm��l�x��g/P�s�8��N�u�V d0��냓���c=u�������]`����|�3�7�8E9*5�7�Z�L������w�k 4k���5�I�6���uF��;����y��#Y��l�qq��o"��la�z���:g6\��]o)�� ۘR�ۍYv���q�]�5۷i�t�ۓ�hq �$mֳ�k����i�J���2�xƻVEٗ�۶�ܯ�l�l����]�.�>ŋu/]��d�1͍��n�v�a��B&�F@�q.��5����GM��;��ˣ�ڵ�����;SFpsǣn��/}���Z���;i��tX�mնS�����۳��]<� �|;[GW�%�k�b�����Q���t�W�9r���cj%���4�sxLv۷6�K;љ���ݻm�llu��{-�^�yξ?�+�l���u��v�O�л��*�"�X;b���ǣ�e��kZ�$�-�s�J3���P��V��:ܱDm��6���gW�/<���[G��v:�מ8��*��Pm�O���&ȳ>��ӟ`cٜ�<=Y�>{]��<�8��#Gd�8�p��z�0�qN.}Z�W�]Ҝ�*���g��Ϸ1�m�����t9ݺGW2C�u���Wfdd7F��˖��qΝ���p��11ʝ�v�냗I�:�m�͸�3�@�RZ�n��L�٥��ewn8���y���D����R�պ���uncb���u���.uԔvۓ���=nKh�����v�0�{\V4����c-xpo���=���vѸ�-�����^3Ѫ9�:G#�����:s���G�-+�Eg�w{���@<�ۘ��m�/�Xѹ�usȕ�.�M̭���`�I���#�8%�mѴtl��nqĻZ�l�7U[����k&��ݟ���('�y,c�u��h��n�z��0��I�Y�Ŧ���v��M���v{X��s��I$�6;uø ��u�#�uđ/@�����u�s����=;7m�)3�]���iq�"kqp�U�up�f9Z8w�:.4g[�v.D�5OZ��ڽh{s778f���;dw�?������q	�W�WoU	+;\�I#��{�$Lc]Ndd��Q ���Lِ줊L���}2A�b*#b��8�����$���I ����$��f�6���/q��V�Ef��n �ᶕP穉�Z�gݳlܞ����Ios��[�$�V�1��l&b�wV����pV��,��q�ĂA'��Az��E��+6��OVD�F��+yH��C�W���"��AWOM���_wN��>�Α$�F�H$-������_���3$Qh%�4C���	�qׯO -W8}]ς�]��j�q�z�/���������eN�$�F���$t�W��o�JL�q�NA�Ѻ䕢Ed&
p[z*_gH�>�g#����*�w�����{#�=2��J���
���6�c����~k��l\w˜�#2څ"\�K-[�<����� Kyo� �ߜ�W�OU�p\�Z����FC�)2�2P.@#��D��'&�$�,UV˩�8,��~��=TM_��ۈ)8�ʪ穮6�B�������I*�z�����"�1>ʡ����>$R�F0 �p�f ��]7u@�A]����vEb�U9(`���$���Q%ok�lKں��}+�^�!�m�/g�Jɀ���2n��):��u��c�R��]y���!��n|�i�$[;4�������(�Zn[�I!oN�x�pXR�!4�Luk�@;���+����S��gf�$���� +9�GSTy��M��77'�^�o�lɽ�T	'�gk	J���C�8F]M���L�J�강闷�2|�&,���nan�	NaT�l�W6&��Ώ^k��|��7�zN�o��8�����uh�� =��$��ڠH!}��&l�&�E&R�Jψ��3�DinW����A>���@�z/�:wCQDe���� ��9�ͷ �q�Tnz��EF�Q����R����>������x�,+D�%��ٴ�h6�-oV�qs(s���p��.��� �]�:�sn~m��e�:�8�.Λ��I ��rI W^��:U>�s3UD�A]��@�!�C��P��P"�Ӑ^�m��<����H$�vD�I+�\���b�髁�'1ݝh���&S0���$��׮I �r�,�'�Ϸ�$��~�H+�\���k!0S�k�i�gU����MILc�I��r	� �1�$�5��dʉ��v�
u�SW����j�zU��Ž�IpeFmX��ȩ]bo��y���T���;�5�V�2f�u�����I�r���(�� s�V����,��I �l�+���|H?<��--��%h�aaX���bI$��bA>�������g��:�ruv�Eu۞�g��t8��M���r��;����u�:�AP�ACa7������"U����*��$���Mx��Q.��o��>+3\�5k�ӈd��Ϻ�;�p���ulI Vw9���u
<iz�����QR���,���"ABuDS��I�M�H�F���P)�F	+/����M�XR��J)�A��w(=y(�!��r��H���Io��x�Ww7�������IyT䘚�1���_mP��
�� ��b��4H5�NI �9��H[���Ϧ\_�Y$�tͻ6@�	�vq�9�}<�#����w�w�6VP�F5S̩�:��r���ɳB�j.�s\����R�Dc���aX�D��W��������'%n������=b'D���i=���q�t��s�N�4l�V׶<<�ɔ��\���sh�	�[��sH��S���¬��k���+�nn��s�{wa3��s�<��Z_\��q����Uڋ�=�k��|�dS����M�ֵ���I��^���\4��H�����;pb۴�O�e���6�k�sV�`�c�R����jr��<�;��ѥ9y��.�:���zÝ
%�ltF����)$�p���omȒ	�̚�H]������q�21H;YLH'��z��NYݏ8n��j��G`D����7xH��K1�$l\�Q$��c��V:��ĩ����^��Y�SP"}�7u^˺6|�7kw�����!���|	�H$� -�'L_�D8��4����3����'\�ȠHwG$���1DV�)�����n	?$�2��d�2��g�J���H�NT��x�5�T �Ѳ��&:�� ��1�r���qH�5��Z=��	������0��;[�K��Y�ɦ�i�5`��a&!�+���]�T<H$̎�H>1׬kB�Vfh�)�;s�D�#:6B�.��(�	�@�WN�|C�;j&��4S���l�1�̬2'������rhp3Ң�t�"��aڧ��A�;|�`��x���/QC�x�2�DT��<<%�uO�Hy���A&>�s�@=�$Irb������!����!A[�A>.�*f���c��^mI�F� �c��5k
��,�H$7?t�$�y��spb���@Fv9$�kު������
��DN�J;�NB�5�e�S<ăM�M,��n5ʅ��%L�3���� �G7�TK�W݁�2
�B!���8�\e�z9�nݞ���q���ݷ�^��X�������/)C���x��\�H"3�d�����Օ5J�{�ɋ��^&;��:l&b2����U\{g!�SZ#��.�ω�>�}�^ �m��l����z\Z)`�%��~���$�z^d�'�Hz"x)s�"ȱ��0��p���h�\닓�Ж�;�Gk�l�o� �z�o�����׌����j��j���+�\Bx�ڳ�F�^R#4Ip���B���$��� ��٠g,�ǜ7�jfhŧ�%�ӲK�`��y�>'�/��Ēv���q=�x%t�n�a��8N�9�˫�Q�]�"(���U��zH{��$���T	$��>���yp�aB//z7�>c�����k���izٵ�L[)=�D��n0���b"=�6(�B�B�e���@5/�h�I؍�$������O�=�NA ���U�C\����$�%�&O5� G��Tr�[�I$���U�	�[���ᩝ�O�9������LCl/:��ު�����r8�y�0��2y�$�r�j�� �-�騱���Y�{�MDưO�ڞ��	��Ă|gk77�j�63��k��12�܏F7��:_��h^�9�I��F����RG�TmF���wyuܨ��ywм�������R⯉�ܪ�H�ᱤ8n"��j;= �"�k,Z�B먏H��z��@;�D�gk�l��edD���Mp�±.���׬�Y�tm<�lNk�z(�S�c�E�1!���J�a��
 �]��-[�#��v�/�oz��s [��J��p����]Q眂�T���ҭS�� HY�@'�Fv�� �<�W�`�����o�[a&�. ��]r ����u��7��*��k(�FB�G���rfx*�L$�6�󚚾�Mވ��wv�A�rD�A��r���]����JʀH=U>Nڎ	Q�Xh�ͧ����4�襼���U'`�� �vk�I�}�&#vd�Sͅyea�7[;4K�0�C�5D*��D$m��b�3�{��d�X��E�W��t�9��l�{С�y��w�~�����/~��s<u�e6M�m�u��Xh� v�ݗ]�v����<P��[�[;�밦�ͺ��B��=mֱ�,Z]�V��;K�v:���mͶ�U�t���<�н�;�v������e;��9�{Xg�'�n`���cIq�:���M"�Sg��Z��\X��V��ܽ�E^��<��m�5�`�3�0(��6�5uJh�cM����C�3�룳��|���mj�G����:]�����5ʝ��t�C��e��������� 6l-����}2	#e�����fv�3�1��b���!��b
Nj"�˻�$��u���'R6Kw` |I��s�I�گ�����bz�E���3Ŵم˪K�$S=�D�j6 �N/s�b�[{���>1��A ��ТƱ%��	�`�ρ��e\����;2	"r�}$�ng����c�-�gd$:��ws�Mr`����ο� a���j��|���2�ޯI'��Я�oH��n�4�L͉<�wJr�5����sV^-�mf�5#Ԩu�&E'�kr��0J���@�M�p�A�y�@�W-�'�Fɺ�uc"�����'ՖV�fM����>�EҲ���M��'��������h��:�z���<��U���x%�qӂ�:cdP徠���2��篧��S�wB�Xf�ü�D5������	�{�D��oO�:��t�{\�3n]"0�*
q�gr��P'�r�S�A(5�SD����Y/��}��*�>��[�#��z/ŴمښLO=�Y�!�$�GFI �w�@�A*�I$��ֺ�M�����Ӹʍ�!�bK���n	�c�܈ �#;$Noj��U�D$L�Úɠ|�f��|c;Xy=�LUd���B��g`�\��nɑ�=���wV�;��!*��nW��B���ɃC�������Ă|V,�A$Fv�j%���3���gLM5�`��.A�r$��n�]L,u��;����N�O�Z�RA3����X}��&e*�|J�O��.��tq-��h\(���"�I� ߃[�\LSd�u��-���J�*{S6$�ځ��R�F0ry���G��<��͸	]�����ܕF����
/i�N'��l���wjG�G��ݾ��˘��dܥ	��%!���L4�*��;�'�<�W����c�<y�#,΢���q2w=��,��|�j��ʏ����2��<���+�iʖ�o�mcodN�B=���cO���
w�0���eIޏW��.�S<�AVсM�`K�\B�6t+�N`�"�\�����1+sӻ��.84Os:�F��=E_z�+!����;S&�;h�n�"1e�ˆK@�a���v�^f�2�{������a�=Q�15�z#ge�z���8[���,�R��������/,�;��� +[��{�l�v�̵=p��ú��vhҽ����t{܀O�;!���A�ྸ��!λ���m:agV��"]{NH�����������z�Ξ�F��>�鮸����w7��n ����{�8�]>�y���D�\B��=�xgwqOv{�J.�n��)����N�d�^���@���*X���-af�ƛ3�5^����?`���C�4Ƿ�~���_\Y��9��tq�@�i���OL�ͫ�����2����X6f󈊾�k:��=���ڡ՗u�ٹ�z�}��/f[vQ�Jקm_Uo1=��7�'��o�f�W�$�Rz�z��TJ�Ia�o�����r̮^��ﻲ�?ew5�����Ac1X��`�#)����$E
Db���dEb+TE�X�R �AcF �T�E`�����(*�`��*�1�AQ��*"�V�TA�(��Q���DTE�*�*��X+	`�E�* ��PF1b(�����AAb���A��F �([Qb��%B�������*"��AV(�m�ۈb����UTQF
e�"�EUTL�dF.4ETC-U`�bi�1Ġ�h�EX2,AfP�!Ecl��T�kj�E��Eb�����F5�V"����"�8���b�(�TUDD���q��A-(**�^s}����RA��iN2���0�v]�n4:�Y=�.�
n}	1���힞����g�q�@���ߗ�.
� M<h&ؚLN�T�Tы���������� H;y�$l�UW��,���}:v��ɴ�:���k���u<e��[i8vc��7�t��w����Hˮ����Ӯ`��Dwd����S@�r�⸸ ����|c�X�灥��'/:sݳ�����SUz�n$c;�OuU|@ޝH�z�ftꜱ	������,4��� ��ʑD�X��t*��[ʁ$���I��-v�a��q�j�4�.;O��2�R�IuR$�G>ڪ�Lr�X,B�7)TwF�L�L\���Ê��
-t���D樎ى�,��vV���en���"Ɯ�"�k�֯NP��)�Dnm8�9zF���Gx�=�qF�()�l�#�n��$��.�==wC��6|��r$�O�jޑ�fS���u>���Bہ�3(jp50$+gc\�[�v�N�\�{K��n�9��J�ms����?��,8-�g�s�2A>5�4$���Vz��r]�)K�./*hP�2Pp��4��/�\�)N<}rd�Y"TՉ�
�ʡ@�弄���ꬣnls�HS�ʴɆ��9���	�Y� �A�X�4	޷��)ω'��T}��AL��J`��.|��4����P$�ܹ�|H�F�H1]�p��چ�* �O���Eص�ن�i�Kf��O� �y3�u���izł{f�H1��`���bIƎF��Ni�~I��[���EGO��o},�ד���}�N�0�[��~]�⧨.�%�nl�}��U]x�k"0��^��D?�k٣��X��\�p���3�����MeN5��a�r�;<WW�up�V���1i�f'�2L�{k�k�z��F=�j�A
�j�m���=vx9����
�����=e#����q���cv�n�ɸ;C�� pM��J��Z{����V�x�;y{n�6�qqŝƹ�<I��/f���a��W^�#���W!�]���-��V������n�Ғ�&����7���
�F�m�Ѯ��ئ�esι�������_����R���?gU]W�$�-�|	"+����"�݈u�II	��� bޑ�΃�`�pÂ�f��=��&H=c�Ī�9�"�$���R	�b���T�b��Wfa #I2�P�pL��m�A �����	*j0y��*�|DjޘWs�|�����/EUWv�mEe�rn�,㘟LA��rO���먇�+on�MwHJ�5#�GS/� ����=�$�Wf\�*9�tEL�T��^�|�ĂB�� ���*�lDJG�	CN`�pAp��ɻ=��m�ܻ�l�n֎:K@;Gf���_�����i�Kf��O��Du�ϊ�� ��[}���3vD�L^�7��[�!C�uU���Ά��k0�c�qtG��w|�!ˋ9��{�U��wՋ�M���v:���<uD���=مB�C��.$�R�D�i�-a ���>!ou�A)�u��t��l�W��L�;	�8-�j�{S2|IU�s@���˼~ݽ�D���rA{���P�$�-CL0ӂd�]b�r���[��B��	�>{r��#V���7�©c \�Y�����r	O����<?)$��I� 7����_���m��`���>%ofUDrޟ��_��_S�.	��9�p�ubA���Ҟ)�z�Ӣ����Dli���4BE.a�_x���I]��@|r�B2�u:L���� �geP$NYCu�6�L�[42v ��}���A�瀟[�5�|O�jޑ�P n��N)�c�l���!�"}[Uu@���dA�yf�ynyM�w��BsmzB�S���OS���O_Cl>fj^~'��!먏>U�}�}*�K������m�׵fiN��ć�7�ge
$ƭ�G3���8a�m�Tک\e��f�N�譽���L\f���t�1�Xu�VA*�:��h"Qi����j��|Et����;�F�˪ �@1k:@�H��r
�2�rjL;��޴�p�!@0K#u�sl�d��8�<	qǋq��c�V���_����؆Jh���w�+{��A1g!$��� ����=�FDd��cVt� ]2�BE.a�\���ϊ,�W(o��u�xO�".3T��Et�I�B�M�uT	vP�q��(���A$m�1>�V7 .����H1��@�A&�y�$j�Xe�B�2D�U]���ZeNv��m�7ӌO�{�������&v��kl�{�����9z���w�v$�s�HEhڊ����̝;}����Q���O��n{E�F�d��js>���=�8a�n� ���$*�ɢ��gc��j� e�J�o��%wvM�������U}��%Dc�\����P�x�vM�Î�@�P��؞��h�y�&�`#�-�a�j��u�$S�$�H]ݕ@Ը��_��0��$y�@%t�؆��I���z+�j���l�)���]����< �	]�J�ܚ'Ǽ"#7cELa�� t�r`�(q2Z.Huz�|V�d�Śȉ�ѧ�ӓ~覧đ�1�-�ʠL�:6!�2�l�x�'�FKVc0(�����~�ؿ�.~���`u�!mG} 	_^Q7�s��E�����C��r|$���Gr��-����@G"N����������d����v!�~���q����,;V��rH)�y�8��2�Q������~��!����A��{��)bQ�S����_0=<m�ҷQ<y���K�\7<pi$<�9�i�L~�c� �p6w��]��\ო���n��@�F!���Zq�.1�ij���4�+�'P�^��=������|��\����gi�d+�E$`tmG��o=ӵ��KAX׵��s�{%�8������n��;g:��]�X�Q��#���q��b〇ٱ۫n�lcmiK�؛#�7[���v�m˟Enl=<�^3��C{=�U�O5���j�b���wn�p�67����Ƽ�bdl��{��۴��P.T�8g&3�	pptt[�3N�x�a�eևF��|z��5���͇#ą��-����9Ґ��|!y��x:j�U��� S�>��pd�X��P�^��gXtaXeu�)��х�˸bAM}��a�G�z��C��G���$_���YP*T��߶q�������}�)��H�$���7��۹��"]�!�1&��: Y��wH�: VQ����5�>�g&��*Aa������9{���q~�|�a�
��*J'����H,�����5�}��Ț@�w��q�����������3��w��$5-!m�o�vs�![����^��18�R(���>}��G��LN�罤�<�;�E�>�nbA���A��3��T����i%B�VV����Q��}�Su:�a�#�����Y�u�
5!m5�~�`p� Ф+P+t�I�|"���	_\�1u<����S'<�ۈzs']|6��,v9�jvNq�z�S0���n-��!� >{��|���@��%ed��s������+����l8¤���￟=0�@�����2z2�Ped���3�vN	���[��eևC�h��cX>�߄��A!��˽V��G2'�P[�Rb�����a���\�Ǆs�����Nm��.��T�F�^ì�LHͬ��e��b6��E�_ 'z�E}HV�H)���'*R VX�����l�%B�*�y�����G��s{8����u�x��5���ya��M����1'+%X=����}Dx ^!��p��`�t��U���X���H[L�=�`p� �B�B�_{�m��3�?���\�.ifk�E�=s��"Ȝ՚�`�l��yH�S����+/���!��$z���#�ϤY�����R��mﵓ�VJʛ�>�����x�������xm��k}��Ãą������6EZ�6�������i��m=��bp+&�Y�{��l�8Έc ���y�o�,�`#��v���Ԫc��^g�X��AR�((E����-َ�L�Nޞ��k�]0�BPD&j�	��h41�G���Lf'ٟsp�4���c&e���~~���:Ɍ���1�׿~����2�R>�X�d�Fa>�>�A�����3�#�K����8�=I������٦�f�5���YS�1��?~��x0��C��|�����=�������׻:ͳl���&3`_߹�����'\f$�����>�^��#�}���ǫ��iq�7<��Lp<��_s��ht9�:��V��6q<zɌ̲c3,��Ͽ}��Y<f8��$�b}��e���[���k�7v�;9-���UH�-vg�e_;��f*��z*	]F�h9v���v�n��¬��̛��}Sѻ3�0�p���P������i>�d��ľ�϶u�gb�Cc1�����<a�'��7��^��]hjkf�tLf'3/�G,���3_}v��|O��`��,��y��vY�L��d��Lrk��{��OY*x�&2��>�p�=�<}����x˖Lf9�����8�&3xs���r�5���1�N�1�~�ݞ2u����VT�g���fٴ/}��ϟ��x�0�Lf0�|���q�S�0q��}������1���\�zϽ�4h'ނwC��⯫ 6 �M��5�^\G<v���/f�:��@��YK�=t箹�pi�_?�>=r��`��?d�>�0y��l�v=d�VJ��&;��}��,�3c1�GȈ��^��G���F�~=�Z'|,��^�϶u�d��u��d����vu���1���)_xj�T�.h�Y�DA�Hd�H�>��OϮ�����u��~�g=�����Ɍ���߽�gY:��S�1�M�>�p�8�c.�A�u�}ӷ]j�y#�߈�A3���*"�*��E��Aϳ7g����f3�bo3��83l�3�2&3}O߷O�����ߎ��=Lf$��bLqמ���:��|�3,�޳�w<M�c�m}/���Z.�,��|��ꪑDt�nM<G��~�&32ɏ<���;�d����	1��oZ��!�i8����3=��lQ�j�ϯ-|�홒�����7��ߪ�#��#CT�Ϛf�����u�ǳf��@�)��%ځ�W�:��)�����cz�|uw�Ӯ���i�c1��o�}��<�c��/Kq.�55��L;�������I��1���{���G�}��I:��Mܜ�z����_�xx��x8ɉ��LeM�{��r�c.Lf8!{����q�I����{���ߟ������ 1���6��4�I��n;{���xݦ�i��<u�	��ߝ��������'ц;��{���x�fc1��3y�{���6�YXbc1����}G�ȃ�#�wV����G����~��'YY/�c&2��>�p�4�^O9���b�Y]��l�N�<�߶u:=}�>G�G׹�~yq����ud���a�c1Ę�Lֵ�܆��Jʜ�`�~����%eC��b��s��g��{L}]�>��>���H����4ΰ�c1<���ٴ��1�&Y��s��t����c&8&2cϟ5߮�]�y{ǽ�ߏ̟�󌘙d�a�ֳ�3��c+%epB��>��q�H>�9q��*F�p����wda��l�6�p��'�|�}��bw3�l�6ͲVV�2�����8é�Ę3`��|��2s�u��3k*�+��}'�\���zn3��g͒�;��{s��h�\֎d�t`���gS��&32Ɍ̲c�<�����1�sYE����{��G��ȉ��g̎0�c%ef	~�ݝg؆3�c1f<�Ͼ��'YX �����>�8���$��]��B��]@S3dZvogPN!S��~z�ɩ�r;�O/g�47xp�>���y��_l\y��\}���<����#������>��j�`*��I��w5�g��z�����ZQΣ<�9D����*^�*�*�6�/y�}	�b�c�x��.SKA�~��ڸ�#�9yt=M�o���*v^���ev0G��9c�A�V��I���[��k�q�x�;�h�L<HY���ќ�\t/x5��m��Y��R�d��PW�{G�Ao���'�Ʈ�N�s���J��[Nb���m�*t󴕓VǦ;�o����q�\�>�-}��]����Q��9�Z�e��d�3����y��I�A�<������h���ŉ����h����F|M���M>]}g}ۧ��-z:>��NkJ�׹�v��ws��l��>�f�W{��5����`bQ�,N��/���1��V((�1�؏W9{�=��,2H�L���@�z|��ݺ2s7ݼek�}/E�;�Q��*B�S���� z�U��|AĴ�ξ��>O�
:��'�X���n;l����O��'%Ō��Sʮ�Jsz{�3mB>Lnv�&���䉫��pmp+���7&Ȉj�ym�^)'o��7���/����z²�!��v��P7;Cl��{8�l��7���,%ｷ�Rj�Nq��ٗ�xd��+;<����^[�-ʵ@������uwvU!���O;oO�<��y��v�:�QF

�D�1U"��+
"���c,DF�"�+K`�"1TF(�*���[j�b�v�D�*�#*"�",F �V
�*X��b�Kj�*bUE�,X�1ELE(��F��
�(

V�r±iV
�Z�Rѵ�b
�[iD����UX�+F#�QX�m��,�+���-X���UX�#
�Q��+j��R��2�3)�����b����D��\DV5�R�T�
[EU�
�+F�j�X�TV�JT�kE��,�F�TV$U�1�آ���Qb[b��A�4j�U�F�m��V��6��RVҊ#U�R��V��

��Zڨ�J
�R��[m�<�ӎ�f��jd\��܉�\�۵�9�f��ff��7�m<=�m��^yy�����&ۭ¼W=���I��+���.+��r��teۀ֨q�\Y���:8^�t��k��/tKlZf��s�&�չ��4��O%��%�nI����nx�U�Zw���qveڑ�;�:���0�Сwv���eۄ��)�� y�͸9�Ҙ�
�-x㭗����U���&9�)ʋ��Ӱ��.�m�'�z�wO �,Yz�pN���o\�Iw�"c'j��!�|0��WIs��gK$��g��2esZ4X�p���f����qJ: 8��bM���Gv;�
k�;�s�7Hc-@`<{3�}s���fM��m��ݝm���:x��a�J<��A셶��:��ng��y.yKc�Y1^��oݗ�������3v�/\�;o&"v���焳ۣ�\�k���s��(��.$y3�v׉�c�׫�]A�]�ѷ&5ry,>
lt��+mĹ6�q������A65��وwE�a�=ku�y�ےyz0���i��s���}�G�ڷ=87P�:��1�m��ta��6ܐLC�kT��m�7j+M�C����\\ف-)��@=�=`X�/�d4t8��g1u�g�������R{u��Ҡ�;���*�n�(|X;���v��Ň���ǶF�W[w˸;����=��sv^[\�\�s��e]Ʋ��.y��A�=�������Bz{	��b�N��q�����=��7����r�sڵ'niX�oWc��ㆊ�p+��P���q=�{d׮�Z�&�{��l���&���ݧ>�l��x�͌n�t�ݑ����c
9�B�&^�����]ɋ��<t�
�f��������&�g]�:��2�QĽtg6��p<[l�N��/���N���v��>?М�Rs�y��u�:�n�<�kn�i3;��;b���qո���-d�Q�{qv�"h���5�j�u]r�\�����r�i6�:����雀��^�l����sJ��0�@�d�ۢ\be�G��su����d��+x���ܼ����y��ݍ�m��[Ds�	ra���ne����}n��Mێ��6z.���>N�.�푾C<����9b��7c���vaƱ��qG9�7a���������ٹ5kp:��f�VM���������2���cqX�x	8�Y�v��\�m�Aqc���^�k�a-Z�Nt��*M&8k<=��[q.z�5��~f�	���g~�q�6�����߾��t����f2c�c&8s�>����'�2b|l��TVY����C\o��ϪW���ɕ�/�}ݝg+*}�{��`�pֵe���x��Ͼ��x0��C���7���o���Cl�}��v~fٴ1��d��2�߻ì�%eI��bLw��}����1z��z���_����No�����}�&=���1u����ٶN'`����gS�Y1����c���ݝ��a�#�}��":�Hۭ�מּ}��o~}3I��d�����8�3��Cc1��y��<a�'���h�*\�A��Bb�>��dA��T���ot*����0`����>�g;gY3,�Lq1�ߞ}�<O#���8Ɍ̦��{�i�7���N��?I�]�Lf8���߶u�z$�bg����M�Jf����u�;�����<O3��d�������ͳhw�n�7��+D�c�߻��Y�Lf$��1&;���l񓬬����Y��g��y'ރ	��~ˑ[Qn��H��
!����>�F�s�nѴ���4��m��r8;���%{n�����c��M�d�|���:�2Vvd�fY1ߞ{���d��Y\OA��>��g̊>}V�o7�.�~�Y��%�{�gY�uf!��b��y�<a�x�a���{[�.*kf�u1����;f�`8�d�{N[���>И���B_�R�YP�{�-�W֠�BuḰ� /{���w�YћoK���e%�T(,�*,F�3:�f
&lf��ѵ���5�R(��++%|1�~���2x�����&3&SZϽ�4�M�1�,��w�x}�Bΐ~�l�Qw�>>�dz���
������Z�.�gY+�y��:��VJ��YS3>���ͳhc1���=�{�o��s7��{~�����Ę�1&8��>�g���c%�Y���bkY�����J�w�4]��l�e`�߽���s�3��q�{�Led��,���~�g|�x�q&3I��ɭk߹3I�0�bda��`��~�γ��������g���l��Ǽ���<a��3a��y~���.�6ΰ�c1<���ٴ��1�2�`�����Bβg���}���W�\3>��y�A����}"Ͻd`0ɉ���ʚ����pݓp�c1�B���l�8�YS>�����U���x;?���V5�n��i��x�!���<=6��\�5��̡�4g~9��P��0�q���">>1��߿l�<x�f!��dC���}���f����a���/�����/�A��o��N��7�}�{������Y�����Z���x	�Lr}����&\ц�֎d�v0~�{���>�#�#�G���K����0���x,�3��pI��ɭk�3I��3++1/���γ�����b:�q�&4���{�w�Ϥa����| Q����K�
�ǇY����|�q�6��c&e���y���%�ɇ����k��0O˕1x�Y��1[��M������jR�G�:D3k�{����y�No,ro���P�7*U�ȤF��>8��VJ�2c0�kY���L��˖Lf8��߼��q�Lf&��Zi�@n��>�,�o>�F'�~=���}��{G~³�tC��1���߻8ͳhc1������8�0�Lf$��1&8��>�g����}׿Q5�/K1�0��g�nx&�1��s�^�	�.���N�c�}�:�2VVJ�̲cϼ�ݝ�x�\u�}��*���,���?f}��L�%eN��f	}���:�3�c1f3����>�Fzϑ�0�0�S�!
%fF��-ۋ%p����Ɲ�lg��N��&v��l&�j�s]���/٫MR�e��u��1��fo�l�Lf2a�c�߼����L��1�Ld�~���:����LO׾�s�˯<��d�5��Y�w3L�����B���6u�z$�bd>�_}�nh��4�Y�u�:1���߶x��Vy�a�ݝƯ�
R��>�""fGI��yY++/�}�Y�Jʓ��bL��{>�F{1z��z�jގ������)�s��<�&9;����&\ц�֎d�u���vu;�c02Ɍ̲c�<�����1���VT�|��/���}���{��i�N��La���{��3��3���C���>�g��ea���m̗8�5��L;�bs3�6������M��������н��o�)�d�,�Lq1���}�<Odăރ���|��3;�����d�����Dp��GQ�>}V�����Ezo��|��v<+o���s���TK����W_N�+"��臆�n��2��M2�VW�B��;���ؓ���UZi�Fn��>��#S��,�0��C��!���g�pfٴ<�9�������xé��/����Y�Lf$��bLq��{��:��|,�L��!�O�4��b��r��՟]'�ǯ��H�A8n��Nzr5�����a�î�� �l-��������I���0y��vu�d��Lfe�����c�1��YSZ���3+*]�
���|���'�}����E�Q�� ��c1����vx��<f0�w��rCH4p��'�|,�>�K�@�G����z��,�1M~��~��k�}��1�Ld�>����O��LLq��B��|�y*^�A���9v�X���l��d������٧3B���j�ed����:��3�c1��3�>�@�O����>DA�ןEF���7���{��q���Ę�1&����x��c%ed������<L���>�*+�C��>��`��?]܋#bd�z�n�笘ϲɌ̲c��~�g|'����r$�b`k_��!�bpa�����|}}"���:��wգ����}gҲ�W]矶u��<f0�����K���W�Y�Jʛϵ݇��i���VS�o��azϽ^��(������{�#1ß{�<d�<q��Lfe5�u��sVLe�d�c�_>�:�=���2��q�M�^����wz��GF�۳�ʾ�o�׊������Gw��l){�Im���L��Լw�[}���R��S{��;�_��a(a�)���r�d�N�G8�ħ�RU6{t�\�d�<�GNcQƳs�YwkjG���=r���q�`�_A)��v���B�$nN�6�뷶e�ק��-�gѷm�]{+�u��u�����[�^5�]�=.�K��B�����i��vz��͹��C���7N��ƞ�YnPό�ݽ���	8�՞K]���w�jB�vlȁt����vn�vm�^k3�;v!���f{?]������K�[.��3���=��~��yx�fc1��3Y�_l�6�!��c�>�8�0�&3^p���֙����:�c�����<d�+%�1�5���ᧉ�Lry�<�j�Ɨ��:�q�Ͽ{��׬�̙d�_5��y�����w�|�g}�x�d��D��L������180�bcf3�}�vu�d��,A�R�lN���Y�ɩ|8�f0þ��2����-�]6ΰ�c1?f���bN8�d�,�߻�g;,�&2�W1ϟG������|oW������q�d�a�޾�ۆ��ՓrɌ��wݜgĘ�L�篾�9���گ>D_�����l�#:OǄ=�\�a�|ϐ�c1f's�y���f�++%e`��l�8é�Ę8�OA���}#��s��|�돴?���Z���|��1��3D3�A���@1^J��68u�i����vu:Y1��LfY1�~{�βu���j�����8�I���޵�93L��8���w��3���C��1���=�g�<O�3��9&�}}Ig��&�ɂ!l���<fˬ�^7aTJD�79���ո�%��������?[f���4���bs3�6�i0q�Ɂ�c�wݜ�gY3,�Lr&2a�����{�ނ}ʬ�}ێ��]�2c72�����vLe�&3�����8�$�bg�9��c��֭�\�3�ц=�}����`�3�ts���Yb#���.�N�m���)7���� �'���S�w���g#�<��,���qx���E��+r{W�ȁ�8����g��6�YXbc1�_w�gtLf2VVJ��>�gY<<�.c&}���H��)}�o��讟	4��A���昮j�E.Ͳq:��~�gS��Lfe��d��9�;�Y<f9c1�=�G��u��|z�N}XNg>�$��a�3#f3��=��q��c1��1���>�g�<��1���9���A�I�}g�Gȅ���;7f#��{�?x�Rq�c&e����g;,�&e�Ɍ����9��2x�8ɉ�2c3)�;���[���nK�&�ޓ�ރ�>��EQ�=�Dt|w�Ȉ`���^ed����:����f31��Y��8�3h}ͻ�-��ߺ�1�a�c1�����Y��bLq���s��<d�yf2\�313Y�ۆ�&�zY3�A�����uhQ�t#	��thEvۛ��m����Ѳ��wM��{O`}6�`�c|�f��q�����w"�����Y1�2ɏ�s�vu�������>���|$��G����<��)n�o��Y��K���g؆3+*3<�����1�O�x�d��l�vq�a��b^g�l8<f�++'�}gO���s�}���L`��l�gY1���&2c�y�~��'�㌘��&32��~�p�8nɌ�Y1��ٳ��~y��o��]�{8�>�1��<9�^��72�j�u�c:�c�>�ݞ2u��D1��C����l�6͡��f0Ș�`�o=��/~3���k9gdNZl������˙���0J�:�G�Qv���t��:�����6�?�*�I��.^y�O��s{��?_�3�>Lf$��bLq����g��Y����嘚�~�p���&8y��b�LW5[����:�aϷ��%��,��v�X�>��l/z�,����l�c�Lf8$�bk3������f&1�̉�����u���>~�w�U���q���W;���:�Ȟ3d9��9��զ�][����Lf'���a��I��1�2�a���������.�i���3Ks}g�f�Dz�w�2x�8Ɍ���7�ﻆ��J�ȏ��@�/X��6G������K�}|~��y��\�l��F6ԃ�[�xWu=[�9�͇d76�d�˂�~9Ő�" �_xa�'�1�������0�̈c1����=�p�4�c1�&3d�����u�R��/���B~70���}��F�dY���c%ed�f&����i��d�'����y2�N3Z8u�i�s��GS��Lfd�P��������O>ןn�%B�+����m�aA�IS���I�+%ed�s_���r�'_���l���3h�y�3%�u���3L:��Nf}�Ã�m&32e���y�3������Lz��ٮ���G��_|q���q�1�7�ﻆ��J��Y^}�=��u���y��g��e���b����"τ���Cc1.��[��g�c0C��g����f����a�c1�w�{�����Ę�1& ��~�$a��7�謏�`�(Z�wIt輪���6{Y�=���w��_=}�6��59m=_\��p��rj�H]"�KZ!\c�gL��+63�������>�@^����f�}�9;�M2	�I�]�d�+���g�zɌ�����OvH�^�A�?�������i�� �c13z���4�'c1�����}���%eC��b3w��l�x�abf�?3.L����p!�a@.�Wk�����H�Ź�U��V��.󝚏�����͌�][��l�Ɍ��3l8ٴ��1���|�l�K:əf2c�c&97�}�0��|�����ZQw���S��}�>yO��~�4��˖Lf9�s��:�=I���}��]&f���5�^C���| �ٛ#���}>���׹�W�7ܸk��g�����Y�mf3bc1�_��:�0�c1&G�0q��}��{ ��>��>�w	����E՚�a�|�'ރk�R�D6`1�d�+{��8�2VVJ�&Y1ߟ}���Y<f8	1��YS��G���W��4�2VT�f3��߶u�d��u��C#1��}���ea����E̔�i|υ� ����Γ1/�_h�f~I��c&L�>w�6s�βfY���c&:���d�u�LLq��Sz��O�>������u�b߾���y#D?W�:�=c19��熴e��ie�������:�a�c1f3�bs3>�|���Pd}���>�|]l�gv&3c�Ę����GY8��zY����N�?}�i��d��9��}��"f����ls���k������"?z���4�}�?��x	����&�O .��X�y���ݮ�Μ�QB�6j=���>P{��K!K�X�`� ��k�nE�{5��O7�vs9�]�t�];vL)����Zů5�����M�(�۷�v;^����6a����ݦ9�,;���َ����v[��݈R�y��m�[��kQt[k.��{<m��')��+u�h;n�q�)�vo]�������o%�����s�ړ�β����i�vy�[35��NIX㋶�b��X�<Z�c����^���K��u�pY���n^��Kŵ�`	�_���߶�5�_��z�0~�϶u:Y1�2Ɍ�,�������:�r$�c�H>�#���^��^>}pu26o{2��g��=f���l�8Έc1f3��������Y�09��s=��ƗV��u�S��3l8�I���G�;�<���+�~�g<�����\�����}���N�ɉ�2c3)�g�}R��>G�G����*�2�푧�}I���}�ߝ&kBj�֯!�T�w��h�'Y�1�̈c1;����� @�}�}������K����0�c1&8�I�������t��r�d̳���nx�d�>篸�bfkF�ءg�dY��j��Dqί��b8�~���fY1��L~�h�K'Y�$�c�Lf's<�p�4�YY++����2��|����ɽ���� a�A��^��'Xt=?�.d�43U��i�S���|�q�6�f2fY����9�Y�L��s���}L��g̟2�W{����'S�2b`�&3�u���4�2V^Y1���}�γ�D��Gf�?��;�߷�Y�;v�k;��E]�m�[���O.�=Z�e��:嚵�~<�>5�.9����C��0��y���Ff31���bw3϶p�m����1���>��Y�DA�̨���2�0����9|şz�f2\�c&d���߷3L����^�f:�3��:��0~���:�zɇ�ރ�kO��:��b$"wv[t"�G�\n1�����r�c�q[�bGU�F��^�Qp�S�3DlEn½Y��^�;:`�A�Gv���7���d�1Ę�r$�bgu�=�4�'�d�����8�3��C��=��j>�w�̬����8�h"Ϡ�E|,�i�q�պ8m�a��b~���;f�`�1��>s��9�:Ɍ����L~?r���������ޛd�=q�1������L�&2�c1�/���}F�G����ŎhCd���^|��3�cG۔��sU�]�O��Օ���b}��8ͳhc1���2��}ì����Jʓoߴu����9��&�/��d̳����x&� Ǿ�=	T���lP��2,��5_\�N��LfL�c0�&>���8��W9�ݝ�j��b��>fH�A��k��3�&T����/�~�gY�uf!���C����h��Y�<߾\��y�x>~���~�	i�7m�7���O�6��9`�l]v̢	M@b!`8�C8�9���O��c19�������q�ɆY�y��9�gY3,�Led�k��l�'S��=����˷᰻��Gޓ��8̟3��˖Lf9���u�{c10�y��.9�����3�ц;�ϴu:0�1��3�������xg����s>�g�mc1���}�߶q�d��:�1&G~��d�l�K��d��n�ge`�56rF���������"O�=s��"eAl�$��E�>w>�i��&3�c+%u��ts�N�c�0G�����"�x�DƩr��Õ��x��	��I��7��Mh9�\��������*[Y�w-�3�,��yU�w�(DG3{Sp_	���Y��q����L��%�vţ�G q�Kv���;.���٘׍�顮#�c$Mռ	�����&k�rbV<������-_p�R�R��s�Ky�iӪ������W�`犬��p^�x�m�w3�`ܞ����5��N������:�~����o��+�8�ȣ��"^�|�Ƀ��G}f�JfC�|��3�~ͼw(�}��.ꏀ�z����N����F���R�836��c/a�bJs�'����� O�����:B��&����>]f�n�馤��d�C�b��7p��G4}������H-a��ڹ]׺ޜ�^5���9'��4�y�i0��/�Z�����f���u���U�*���}����eL�\"������k�1�"����.ةv���"��9�����?��	�><�	
Ϻm{�D��v!܊k�"��8�W�M�T��W �sBJ�9꽾�%�{�g��{{��]����7�����^��s���g1fo���$ yq����.����
�6Lu@9�A��{�?g�{��>V9»�C�o�-�]�Wl�%(���v/g�9�}Ewr����<����ᩢ78��x�u޵3�:��/)F�@�2IH��kMe���7ˏ���:c4R��j�M�|g�K޾�2��S�=��Z���h@{�gn],,uŽۮ��� �������QYT[eKlQU�c�P`�ڢ�*��b#"*
(��X����R,��������cmm��Y+P�TKh�V��iTm�ʖ�DbZ�����("Um���-����B�Ե�c�UTX��F���[[F�-��*�ր����Qk*T�+[(1e@�lUU*"����eB��QJ֢�QZآZ�bZ[b�c��E����Ym�*m�JJ2�kcXբ(�Um�ګe����e�j��cZ6�[h�R��"�%���*�"���[-�*�[j�[X�6Q����[mB�e�)��[mU��am(�JV���j}��{������3��Ľ����8Ρ��1��d����a��1������JA4��'�}�|�؇��_Eg����ʓ�33,���vs�βfY����\����:��VJ��Yܦ����3���O�-Y����|�����@Y}�,����>� w�I���Zh6�xY�:�>�:�u��C��1������i޿�p�gݞ3�6&3d�~��gu1���1�_}t��p�317���ᧉ�Ly���g�4dm��)��"e0�!	�[�t���^��:�� `���#����u�������-�ӗZ>8ɤ����vu:���d�d�&:���8��W�1��Lf&oZ��@ϙ| �����ÿY�>��U�ru�gP�b�f!�����u���;�?u�L�MiSU��i����=���'�G���{�OV�"2����ܫ�;4w}~�`���l��gY1����Ɏ��vu����LL�2c0�oY��p�m�3����gf�&I׎TPP�@J>�Whw��j�"{����c-M��ɺ�H��{j�PN�HiwpLP��*d�uHOgQ<7`��	$��&�@9�t�$7����Z��U(�ҽ��Q�������q�D��u�aHy�B�7^IQ6F�*qT�B�8��t��]j�����+��[�rލ�>Xz��_鿥���H��l���cF��
P��Q�ؐ	켫VDE�!v09&�V�Q4�inD�I@�WTג����B�Ⱦ�xc`��8���]zG�m�=7g��n�T�T1t���sv��������&ّ�u��XC���ѽ}u`����W�{�7~�� ��_0][Ԅ�-�ڹ�u����"�^lDY����V �ޙ��F��ՠ>S,ߜ[�λ��:�Ц|�d�Ѩ%��~l��ulɤ��գN��Ն��W^ �('
�%�J�ޭ��}4M�H�A.#钭[�쎫�ݹs�D("v"@A��Rl@ ]׵V� �a��EWRʁ T��I��鈚R	���)ub�ͻ�<ڵe�s��}s+ҡ�>���� o�n���׽RnWk���lUfADR����*��t�ۖf�I^�\w�2��N�]��.݀��t���4zh칠�s�(
|X��#%�vY�)����>���/9�⽛g���`6Cqn"<����{���;��"�Ku<�4bի�vS��N5R��o9퍶'@�z둒��ǂ��Xf,�ۮ]�4�^x�'m�8Ů<��˹��u=���ON՞.�\S��d��+�u��G������իE���{������.��.�s�痑l�g�M�vl3c�&؀�u�㞚}h��2M�x7��z��p� v���H�G��Q����ۿ��t[� i�E�;���k2�X k޻���m`��A�1���R@ѵ�u`n�(�*[��nl����wa�q$�G���2$��9 GVm�� =� �b���6\��iexH�1���U�ڰ@��Z�AT��v�Gyɀ ^�ʫ��w���G\Z��n""��]�3W�X���{U�w �C���l-fU�� _vMmzT°����5��bV������=���}�����d rzjE�r�`Pv.�(q�!ˎ�ue����Ʌ�����H��on^��n����Ip���o�H�R	���)u¬ݺ��";+j� T��(+��޾��ۇ��h�o��d%�5q�1a��Dt,	OYbߢ#��dlи��H�4���]��3���zz�r@O{xyP�eK���`�j<0�(ꫜqX�z^#na^�w�q�J�ܪ�@ =��vB^S�K�7f��q�w6�X8�"��*,��]�| Q��W� �Wr6�G��,��ԓ~I-��H�Q��!����$	����͡u�٩�.����n ��Q`S�d�wV���x�⫗�l�ɠ��AA��D&E��t�J@ W׵j�N���c������W�%)����"J;յ4����Q*�8��"�%PRpY2�r����a�0���כΞ�򛵗H��b�{?�_�����L�.#�'�����@��1���OE�����z_I �UU��W�A��6H�D<Ι:���t,f�6j�H��1��L���RM%{5*R�v�
���n�wd���d �s�0s�P	�o�� �r}�kuz	
*J����"��:p�!<��?V��{F{:l����8�ou#4�����\÷�{q�`�z1��(�)�c�ͷѮ�v#� �S��DPF����[����D��m�4N�q2�rV ����@ w�n�7k�}�U���;�
j��D��x����QM2&\[�m���| {k�����Ӡ��=�7e��� ���ՠ>��Q��;uY�(�P�0��� L��j#��b����+�h�@�>L��	��Db�w
x��!2.x(��|�@���V˶z���bd���>B�)LLT"J������Q!��jL���$��e��4�]�l���M�K�z��!���{��j�ӱ��b'�� �C%�)whUٷ+�A�[V�>�ɷ1��y\��{�| /e�U��;k�}	�}�⩖� ��r|M%����m�^ǽ� +�꨿�@/uu�E�	�}7�H�Ο&ʛ�]B���=<Y�we�kЏ~H�0�<��r��/L�_Cƍр��`p#�p)7�1=}-{�D�3�QwF!��D�	 �eI5�O4h��٢y�NRI ���!�_�r�e*�	�' =��4���ڴ���*Ot�n�	���Mj6�03���m�є+�z�z�4�r&�,<&-5!?6�]�d�DI$�șq��e��X쮫��AS>�A.n�b5S�{"�S�����H�໧j�%レ�I��@�DS	�}�i/�D^b�ss*�+]��q R{�b(*�MX|�8��ݎٚ$�ʋ
(����켾wh PvRM�"/B���ƞ�vV�3+]�A�����۾H#>!��`bra����E�׶e��^��_�| T��� �#z��N.��s���u���}�@OKr� ���`k���YՕjʇ�R�v��DZ&l�́�wV�Xz�ݢ.ܪ�7!��S������hژ�*!�� ��{�=��G�Ů��������9�u��!HFK	bP�F$^l:�׷6L�<tdz�z�G�=��oj�ڵ�X�4�WY�c��Vû�=��;΍v]��m-�٫<��Zl[�`8m�C��O�i϶;�����縨�)磍s�x�zR��D��覊��A���E=��k��:YशWnB�(W[��;�x����q�'Wn���v��d�a���uě���L�T@@.of�|6��[1�{8��i:�Kc<s�d6N��a6-:�����X�D7?���@ ���I���۫A�o˜�߰�e����*Nɦ	s���D�KL����W]ݥa�r���ڕ52��	��Ј> LGlA3�zv��A/9b�.���m�G��Z5g��2B�2.l(/i6 �w�j�1�z!L�:��� >*Od�̃�#����	>�'��I*e�|�v^�;�M���j�AaYM�$�Gzr��	 ��5Q�I.n ��{1����aa����/�! ��Q���{���M����d�$�YU`#��݁:_5Yڡ�����G?5��._&n���Pyһt��v��3�t�Üs���K�{�<咘�M�;��lά�V �]W�����:��|L.��4PHU�L�ڨ�nL� Õ���;�����<z&�Q���a���m]�c94��_d��餝��ʌبmݣ۔��qcU�p�8z=:�m޲��Y۰���Չ�Ɣ�6�A-�l�Oē�O� !#�p\P�]�YvuM|�k���D�7��n�]Wwd@�{k�Z@ ��p(����]s�I�ښ	�]�Ή�pp�!X��"�!�nE.���˚�Ӧ z�kԗ�%nN�H�)vA�Q�A6,�H�}RLcq1 �mz�;<����sw�9�G%F�4U�]Z�>�qa;&�b.�ᾔ�~��չ�ud^�Zk�v�]]�>��]j��;n(�q�!�p�ݓ1'|C&�){�]{�v �k�	�A�vD`
\�)�����L�#{��5 ��
Dv���-����]VM�!ww7I$�K^�^	9;&�A}�� ���_���nE���i��D2b��v�h$ҽ��'�Z�h(��Z�x
��n�7�d���AQ�z����{�x�����j���:�":n�c�H�aa��+��7v��Bv
�N������I-{��$I'd�a�<�DI#pșqnЫ��9[5ûI%T˒m"P"�"RA!Gum���V*ܛݴ���w`|�
�b%��5��o͒H띚��[�q�V��t�a��{��"���I2oV�D2��']=[�Jݶ�6��7	�⻅�z�Ʊ[t�]�U��wm�v����v�rg�"&TKl�������0���շW�r��s5EόE����I�mZ���rA�����Wf�� g�.�~v|��H >��ȉ	/$�&�ےu�y+�i��"5�cLP8s�09�` �+*���z�z�_D�7����|�*L�@��;�n��ݕ��D���M�Ֆ�y�����V` ho�7|��윩��=��M��geGuԅL���YV�F�x���O+}�y��H�f�\*��Aw�R�UuU8.Y������7��s�=��a�}.�s��3�]3&J�|9Z��F�2�݋n��� =�V��y�j]VWU{3U3@Gemՠ>׼���&`v��:8��9Nz�.Onݤ����ls��:����Oӯ"�i�N9�O��w���m��Ѳy�|�A�{]Wd@���\_�>���σg�X̓�k�@gV]Z>���)��>l�-�;�>[s/faU!�3 �GeuՁ�׼��	�z��'����%H)��R�Ы����	<�W�GNW�`�����F���e�E�9�;�>*�E�^3���ra4��y{X���t�v�]�@ ���"- ����{��Tx}]uh�tv���Y#�,��;=�v��M�oi]vKπ�2���- c�w �9;&�+�;��lo�������r�x�Bv���]��ӻ�>9l��ڰ��{�'TKQ���L��xD.�ꇣ���%���LR���u<������5j�nx�cpLK&���[iUMJ��7��k��-ޜw,�(:f]� u����bb���{����~z�ק�Ě\��N�;w���vNG��*��#�d�����E�c�&2[�Jx���fr�;�}���k�<5�=�=�f���I�����W��O�貵������b�Y��K}_���I�N_A�"��ʮ�N�	�6��طa�O�g���D��=s^Y��=�\����=�O��l�<��zW�!N�f�,MkO�\��z.�AW%~��s�����	�6p�:$�R����FP�;�T���ʵ,,�3ѧ��s_gmc�������/��j���\[�}7;�Pl����'����j)U�->����y��o	��Uy�V,|�gH���yl�c��i�jn`r2UrI5o@<��P e��x�8�5'�B��,�:o>����C��l�-�܂�*�)g�I �{���"�[ń^�h��Noo�a�g��|n��NO^�q�'V�ѵѯr�صs�1J��0:��r�7����q�!;�Ǝ���)��%�6ڌ��m]����tQ|;ӽ�v���h���}x�ro�����<����N�սz��n ���V�����#�u|�}�m�������k�q{۫^�O��t�%eV�64b�Э���Kb�
Ѩ��ƶѪ
�)Ym-mH�JV�(�F��F��J#hQkaR�J�V(��P�ZՈ��,Z��2��+ETR�Qb"ʔVUj�m�XҶ�QVҵ�R�JV�+P�R�ƨUDEmPQA�KX�Zʂ�m��D���V��-�[k(�������QZ։E���YTE��QV��Q���+j�U�j�V6���b�إbZKmJ�6��Tb!T��[F�%�V�"�+kh��j�jѭA-( ��ET��im��mV�-�j#V��m��aF,���[mTUUm"��E��YX���Y*Q�,aF�eD������(��J�H��JKmZ�T�h�(�J%Q���TUH��(��J�U�,Aeb[T�[`T���#���v[�Fj��r�睋�y�{a�\W)�Kp'C�:g���:4&�:�!�����v�qۗnr����8��ڵ�#:�{<h�m��[���X�vE�h�k����ny����d��9n���[lms�Q�����ݽg�NS�Wu���ֵ���C�q��`��X݃��&�/���EKYy����v<�0��6����Z�WۗK��d�Ž�-�=U왌�=i���v�8�5ɕ�v��xz�p3wg�M ��C� �c=��t�vwg�;m�5����������{�ԎnP���w;:�Y�ݹ蹵��s���kd݊{
��ϡ�1�o���Vr=����rN�r[>�VZ!��m�s�non��[�!O\�|v�Z��e�ό�{q[��{W*Q�����a�m������y��wq���6L�e�n^�걠q����ex��v,�q�fb�Pt݇�U��)��s�ٽ!����8�n��1���dA��Ʊ\a.s�����o1�q�{t����&�g�`t@��Y6֊���.^�C��'	�}�c�kv6�"�T�S�V/TV�;����[�ۋ=���7!��c�[&u���0�l�d�H��g�Uq�G���1���3�@�n��+8g\�ڭ�fޞy�����rk��N����۠R^.���x��I���GnA�=������1ݸ�kxNݝ�6�'<'K�M�e���2U�u�G��I.�b���]R������onɫfE�z67:�����qv�m��5�r�E˭�p+bѸ��dp۝v��'h�M�X6�b�k�8������p����;%̻n^i ��ꮻ�&^.���ʐ�]�s��ѭ�`�<vFE�Q���7�m���Ĭ��\7��N���.��y���ΒtB�Yι�ӵc�xs=sw����l�GZrgv�{����;`�Nl�c;����R�ӓ��F�R�8��8x�yں0UnoX�0�̉l=n�c�>��-���қ�k��y�NNFxՃq�6�W�=7n�W��6�:5[X=�ݘ{p�=�M.�6:��]�a�q-1�t�W\u�q2���2v���۾|M��3vy=x0cV���P���1Ѓ��st-v:ϐ���wF1�s�����z���n;=K�1��-�LF�.���j�Ov��ت\OX�f�mvq۞y����u�cl�+�ʇ��:���)����\O��1�7Suز<�ۣ8&TC}�q��(p�`�R��SUT�z�]Z �	��L�4�#_Od ��h�0.�f�I'0���O�?.T�L�Ə�7�P^�l�E�=O��ʵ`���y�DX��i�G�߰!��m�|IWu(�8P	�|�v[�waò�g�aUJ�V�ȉ�˨�� z�]����`���3	!� ���?Vc��"�,+}��� @|�s&i oV�eY����L���:��փ��i��L��V�j�>쬫VD^w	���*z��$�/6h�D��^�L��ښ���Կ� G4�)�h�g�`�9W[�f��B����S9sv���?��b��0�A�#{�wh a홠�[uao�e��w���ٶ��>A;fb��8�D�匁��.n����0E���꫍�Ӿ�oo*�pH*��c��a��Lhb+��۾Kۘb�������ޞfوu�p$�e��N���<Uy��+պ�����Uk�@ 	��&h�7��-9L�����T�L�>dT�
ٚ�W�uXA�DMCs=��G�9;&�d Gv�Հ���m����},�E��Wż�[0���6I2�ֆ�H��Y�RM$�N�5�
"B�v$�!d)؟4���A���	���$�K�5͠��u�pz\mdS�^��s9�5��S4�'�y�y-|�)*p����S����u���Ҝ����FMی�[��&z��LP����:Gi�?rU6 }�U���기�LTV�M^J6Jɤ�;n��7M�ء�)r��v�� 2��z�ͫ�	�I�"�]U�@���v� 1��#Y�t�ys�q��%�͸Z�W��� �o:�^�˭�>7�
t�{3}�㜌7�v�-��=KTCq��oH�U���C�\�I��9�����f�C=:]o$#_p�,l��S�O��=� !m�Ur�:�����+D�Lh��Sh(/kޅ��t�tc�]� _���!���rk�Z]�q�*_P�WJ���$�97gĜ_�RY0�H���3N�@ ��K��U�q�Y�w� Wk��� ��L�7W�ʲfl�v�y�GE4Qn0A0f�7qtS���2xލ8�s�/i�"��A�r�}~���9L�R�[�v���5�� 3�3I cS�'ʻ�/�.� Wk�@"��2G�1@��v�0ꯩ�s]��x{�z�Z� ��Q`$�t�>��8������r@(�7Sb�Х� �;}n�""!�ڦ|�H-Y�޸����wa  ��F��ƄaC��I��^t�R=Ӕa���e_O�
���E���s@|=�U<(n���n��F����"�-Z�:�r�c���Ȟ�x��|��((;$nkJK
c=Mm��ne��dڝ�X� 黋�j�C���%��U�1�< -��G�"��D8��7���D�$WN�R�w�u�*Ӝ�J�ꛋ�" g��́ �z���7:�<�=|�?>~Oc���;�G�'��a�a�<���G��u�Cu��0kb���~�~+ߦ�,K��O��4��H���BD�{�jI���I��,�;s�"�%��>i�W� \�꼄�mI�%&�U<�]�}sn�b  �u� ѽ[u|�a���O�=+������0��h���#�J��ެ�J� �]]\+e���I'BM^8&BH�;SI/�t�M�%��� ��������^x�	3r�� ���mՀ�y޺�vO�F ��[��sZ9�D��l���h]WwQh"<��Z�J開�s��V�Z ��y�A���#.z;f�5�d����EVf�=�Z���_H7��N�a�碭�J�P�ݐ������]�lb�1掞Ć!Վ^2�ZOR(�Cm�,$z�	gW�=E��<)��j�u�2�zM<���ͱ%�1�<G��m�2�Y ��қtX��m���t��Z�O�_� �y�S���rݐ�gc`;9p,�%�!�=�c�T��J�[ n�ыr8��.'��py�v��&�����i�F�iܼA)�
q�mj�U��n�s�ގ�{�sRWɐ�������w����B�m�Gi��u����W)�	�2.>���� +�ڿ��y�XWG���{x��;Bmw<h�������阈�*!��e�-�;��5Z�v�z�u�Y�������@���D@Ftw�y�dF��y��+��D�.D�uA	�ۿ� 9溿�AN�Q�ܘ=��pO�읩��H��rM	���-�2!��N�#��dmɔN�DG~��� 5���@|v����W��L���+H�ww����n�b%�%��T������I��^8ѹ����duf�Z N�;���;\�0�2�������_��Z8Z%|q���ֶ�]pN���p�*u��et�r������?�dn�����˻���9Հ��!��i�,�{WU���ug�����w`iȥjb`�4|ȹ��/��`-��]k�f�j���mΓ�t����n�t�����9���wCq��f�:��蔠'�F��١SOB�)���`��������0���qa gk�@��-�Z�e:��6o7Հ}YU3*��$���h��w` �Tπ@�����E�Nw:�|������Z�	%�h��	����ET�������@w��W�F�몍��6�b<�:��$�*6θ��\�!݄a�� ?eT>-��>�DT�r{�/$L��ϼ����SA(�K�w���0}?�lĦ�=v'��/'Oc�Ӗ�0��1ϟ����bӯϯ�������z��� >����k�����L�Y�k�;����h׈�S��E�ß��d p�&y��^�V� 
��1�s�ADxvV��Wզ���$�hR.�&�^h�XE��N"![�V ���l�N�d���.��򅥘���eK����U�;�^K� Vr��jLՈ��}�2��|����4�avu4��./v�]T]�I�w9�E$5�L�^����h$�
=U(��Wf3]�fc����hVW͈ ^~ʫ���w�1��*���k�El���Œ�9L�!��gi$�J/��y''7�<s	ճ9�4�@E�˫�	��w�^�3}���S�����@��
[�,�ݽ�O;��,!��N�ԅ��ϝ癏�����Zy���;�A��M��.~ʵ��9�W�7ޟ^��={FI�4�sު���:��n&SlAe���@K&ǹ:�0-�M�|�2���ί����nѕv���sX=`�nd�͸[UU�>�ui �"�{�#�]{��F�[�]X ���z`��>���>s7�X_g5F�8]�F�D��ْMy$-��I$�����v��C!���V��.n{8ʓ��_(�-�s�Y4��`�:���3�[:+|�8���Sf�p����F�}l{h7wf�h��;�7�w������E�Z�dQhs-B'�e�Ouݤ D4�$7�)L@�z�!zɐj{�i"M����H C��i���s����TT	�����������G)F[vvw����˲tC�7l 8c�Y���)NS"��Y�v�>�瓵rDD9�ٚ@s��ݫ*}�xw~��I�G�W�|��W��k�0�ݠ�����=z�Uwꨴ ���� 9;fb)Ḽ��=59�{[����r8Cq2��e�vz}dZ {�iG_#�sx{�~��πG�O]� @!��5�k��c�L�6�!u�ߩַ��^�s� >���)$FlD�J�mNI�v� ۓ�jC6b��>�f��b�����b �ڨ��nw��m.��W(2�n�|��4�s�Ͼ�St�|�\D�U��UZk^8%]MZ��Z�����M�{ۥU�պ����xq	ܽ�VU>&��}�@��8��s�6H8������3ڮ �dI�:�g�5�\nM۵�c�Z�Iu���ͻX��`gvt����Ǟ{3�=nBp�ݩ�lr���O���R+�k�[���7�F�Ey:^�oeLt�Þ��� ��n����5���{Pt��,i��P����m��0,���qs�V�N���.9����˓���c/\gú[��)g;v�Z�;f� �7o��)ڹ�ur�9�aS^�v;����E�2�"~�W�E>��,"vRl�\�j�5s��Ͻ�z�) ivD��Y��	%�)Hw�;H�?-�M��ߌ���w��"I$�iuHE|s�e���6c(��{=�z�}��9Rᄌ���0:������XEb�U��nb{ӹ�� ��1�϶�����#�4�\H�,�˛��]��G=��H�~��$����� #��^dT�屓�&N��c^'��[c�L�4�[wwv ���ԗ�>̇L{1����}%  �-�]Z v��i2����"�;q$B�l�ݹu<�v����!m�)=`��u�㗵�F��WWiq�l�~}��97�}����Hp*{�v	�=��	��K럳|Z�-DH�M�s|�#�cI<_ɗh�+�b��,\y^�?H{�k���3]7�*��*�������/��*���������r�ۓ�\���P��PP�盞Y�<.˷~~ȴ�Q�I����uh7J똋���!��*�:����!D�L19>9���Bp ���qa�]�}��ܞ�`�-� ]v�fzL��fa�	���A�M���J��A���z+2���k�� ����ަ���"�#W�η�;��%̹RQ�����==N}l�������3bGmۿ��lemڢ���ٯ��l��={G<s�{}{�Oh�Y�1N2cNt��wl�⹝*x�;On&n��������U3���躻� ѕ�P �O=���[���;-� ѕ�tyMy�T�	�85�*���!j��a�Wf/�h��4��v�H��f��|���ΝF����sԧ�b4�`�~�������"(��+�O�uet�ָ�nq���;{��oM�����Y�b�_����+�:;���Gݑs#�ه/�f�^�/6��Eԙ�i��h���`f��Aq��=�ϗ��|�e/n?S���n����텕n���m�"�eԬ�H[3��a�otD�rcH���!�m%��]��-�/&Fk�wYr�-ʫ���q:^�\c��EC�/�܇�>��;pɋײ7`ab�VA^�x&�VD\�+�PŷT{i��=��Â���W2H�R�d/���w�c�sٺ�48ˆv>��0;��������kGm����z�i/[�9��n��lФb�Om�b�U�ӧ�f�j�b+כ�d΋���^����v�]�v��KՏ��s#N�"��y,	��4�g�OM�Зq�� ��K6x��&,�}�$#vyEQ��<�������"l�D�x(�Z6����U&��a�~�/Q�k��K��vL�"�
��#w�x��=��ڐ���h`Rx����f�$VC���)��9m^�B^"�{�{=��L���c*��z]�A��ݐ�z�j��Ǽ��3�M|�vqȥ����aX�Ǎ�]����g`4a���Ѿ�8�tT�g��Z_x{���KJb�4D<�|����97��<{���������1!+�~N��&nՀ��M[Q0B!�����S���)���ԃ��-�l@�FRŖ#�}$��q����ܽQ`�N\�<��$��iF����my�X�ŧs#okc6	٨���6�h?�q����aF�J�X(�kh1-,`�kQ�#RՑdB�(T���F�R�%B����)imҥU�����b����m�UEcZ����T����VmbR�mHګ �X��b�X�h��6�J��X�ZX-[E����1DEF�Z"����1b*
Uj����,EQX�h�Ԉ�b(�"*�ETX�-�E�AUU-�U���B���mEV5,b���mR֢�*�j������Q���$-*1DPD���*�U����[K�֋F�YEF�b,(�*���ڠ�TV�U�U"�6�X��H��DEE���jҫm���"+mQk,TA#b�*�(��1)E)� �F�F$UQ�DJ�TZ�+b�B�%eZ1J�V6(�V�"���Q�X~����� ��� @=;5'z=�B&�R"ғ}���L�h��\gzhJI ͞��������×^ty��#��&�=�Ռ$�,$�+fO�5��\]��f�b/��s�%��-��a$9��"(m�A�6���G��m��;qVu�m�ru�8��"��]2sY�N�ңE���7o߯���-�Г����w\��3Ӵ�� 4}��=ī�{��[L�&�p�Z��Q9犣�1��p��u����J�x{�%��*�6g�\���>s�d���݀��nW��x���/�����c-bBЊ|K.zJ@|:�*" ��gaqY邯+�ݠ C���� 4y���+�̊-0������w�u��[�U����0��NO�H�̷h6+z�1WC���2�	׺��n��mm��/��C���
V��B���Y%{}��]�F,Ӭ��Y��Ы���8�����U���$l�M{wo��(~�N�~F)vG�D�$�!K�*=�w@ tVm8�]0v���l�:uԔ p��$�\gz�V��g	�{Cޑ�����u�olk՛M�t瑽��Kv6�K�x��#����V��}�9S2���}�㦩���̫T��n��Ӻ��/�W�3ӒDR@+e���݆8R�$r�%�ڪ�<�#{QY��*��p�D�O�n����z�&@-{�ы�/UW%��'�x��cM��m8��t�BA�7��a��2V��۞���@ #��ua|u�1kyS��D0����*��]�-\�TMQ$��ɒc�,�޹��@!�N�G�:z�#R���@*�*�	h�K.�-��ڐ@:r�s�̪�Snv�^�դ�v�I����N���]C򕱖���o.�J/w4=⍋��N�ι
n]�NH]��j�����H��ج����يY!r��1	�K��4c�h�^K[s�ݞ=��{��p[r\3=��G1��۳�j��ϝ��=�.ɮ�G<��Î�$���]���3�2õ���g����ӳ=���n�����܆L�:�^���3nyv���q�T<.���6̈́�C��7�[��MI����5š-s�R�m�<�W��N|��� ����`�5���\ks�2tp[�b�$������K�6��X����ێ���v^��@�ȈM��ct�
 �2Q䇛�A�'h�@ ��{$Gv�?[U8��+3�V�D��E����,D�1L�&� æ����f����UQh"Ϟ� Ν��"�:�۽p�Y�s�Q۰�
Zd��)�#��� ��9r��g����u^umZ ��" �sӳR���2[s#m8�~�v~��|�r��$��DZ=9%  �}�Y�ڣ�DߠD�ö�!?�lm7�^�CT��b��I�f�Is+�G�!5>IUz�- ���"(�n�����魗����v��;�Pm���;����cl=X���۞�<�-�0u�\���~'=���^Y�E��v�_ ;)�� Q϶�Į���\Ò�gr�S�H��J�%��b�
 �2Q�}�B�I��GcJ3Nt�|�f��;f���N�m�>�\�cY��T3�L�j�}�j�)RlQ�I�h�NcE��q[Y��D�/ad��u� �grf��@}�4��O��/H���������O�8K-��e�7�&���Ф�D�yq2��=v���$�I��L� \�j� [��)i���P]�n���V��#&x$M)��8I��yS^I���X0�gQ�$�M5�~D�hy*�2�i�qL9��I��yՠ}^�'�>*�w�@�&��_�
1��DX���M:���X]�������Ym�;(]t�G��L.v6����E:��v�T<S�ػ������\gN��˞��@ �y�t �[�q��rv���â��IA�}�� +��R�C%���Yv[�wh"'�=W�Ǿ��=59> c�[���wh!�_E�@P�m�Ttp�zl\�!@��C��ʏn��@�#�5Ձ�+8p�$�`c������.�����Шd��ub�\��Q��R:�ùPK���z����1l-��E,��r!�y��n1a�r;�r��I3I�Ӥ�Al�:���1K-��. ���a�}}�1y�l >�]|ޮڸ�����gծܺ9ػ.�f5 ��z���;[&��	d)vZ;}�v ����>ҋڽ1C�P�xλv ��w��ґ35w&���cc�I���'\��;�Z{]�Y�l�>M�Ku�]u.��k/cfu�d�r�{1�U� ��u �9�D��cvsc#{��<�<�]�����S��H�*l,��rA�t�=7Y��s�ꮠ@$��٢I4���L�,�7�"u��:T���	;wQœ)�a���U��
��NDW[�uι��=� �}�i"��k�bau� �P"!��ܖ}�R�f�X�=����"�� ���) ��G�o�e�nL���Y+����ۼ۽0n��zx��D�-�+�W�kG�8yRxԖ��d6�5x�-��4��%�f�i&�0��>�ω��wh
��X�m�q�F5�$�۳K��͵��' ���|I�E��I25>�d�;\�ڌ�m\Jxc��Q���KWus��hّMv]�rc�l�x�m�^���@�e7���2T4D;\�.�P@|�M���݇��`���=�u��@Ó:i0�1�:�2e�Ke�a�;d���y��vO[���� |�}�4�6m;��W���1r��Kـ�IpP�
�PL�[� H.m_��W�_y^B;�� "��3@%��j��I�@�&��R��um���z:/,��w��n�g�|�n"�Gms�;b�w@߻������bZW���&�e/7T��'�u�y*��ҡ�Òi.��	$��禍I�|�BG�׹�[/��R�5�IY��qoK���F�!\F޴��_��-5��g�3��{���<3K�86�=�}��ݖn�?߯~<a����iӳc���Μ��cz��ۚ�j���m[�-l8yWp;���B�vw�T��O]�ûb#˻�-��Bޛ9�*e�5�unȝ	�������ݑ��(p�.6�㌦}Eu�{+�
�#6у�2�un�%�7A��wq��>�Y����[�L����n�g�<*�^{�op�����{Bsq۞s�fN��u��w�ѻ����.N�(a�j�����w�2��1	J�,��yK�L$Mq_�� 2�XD��qa:�d��]���KW-��/���a&�����S#�a�/9	?��9N�&ӓ��"�η`|;k��DB�̬�;z�����Hs�q�j!�I��.�z�+" ��:� 7޷&L��|%{�$גAv�:'x�f�Y��T�.z�?c��ު@ Y��iX ��qh 
���2��v��kY���3��rv��Bzf@�-Kh�e�yZ�� (��Nnk�{���D�{b*=^��|Ǻ�݄��baOt���0�ˀG��Ų`������F �˻�77\���g��h���߽���"�e�|��*3��* ��ՠ T��+���Zr��^�� �\�"L3�X�-�H�&�7%$ȕ���b�κ��z�է�h�Fw��zkiF���NFWS�5=�+`=�ϻŅgt~�qέZN����G@]�g~����TDDfW:� ��f�� ���za�εݻ�U���Ѱ`�a�K!K�μ�� Q��Nb"*]Tu���=���sF��\�"-QӲF�9�����m�����u���gy�E�ܾuh""SϤ�����DX�91�$;�U���&�3$s7�Ys�W�����'׮��{]�0��u�Q��R@����%�F:�M\�"i|[,(\j�&7c��n7s���v�%ѝ��a2Ns/v;�����(NZ��%�qo�ݠ>�t䔀��N��]��΍�o�َ����9=�o I�?'!�߽&�M{;�N/n�������_O[� �3'$� >�q�6�L���c����S��!�a8�n�a�t��2�X&���yy��Y4��6��y��$�]//����ZĪ�6�V]�j#��8�o��׭4��7<�x��}�˚{�{��k�C���1!�{u�w�!��MI >�w�2vvaLK��Z"]�v{���.��S��YQ�����˯$�G��1��(�IylTtO�!��s!���8�U�c�� y�:������}L�'s�H8ɹ) �K� 5�;����gK}N.殺��T@��($������9�v �#l;t:�7Fu\Bl�O��������.c'�˞�����W��\���%\ox��&��>��2*$I�vݠ>���b�	�R�Ĺ�������#kco#��D��2f�'  h�m� ���@h�����nk�igL\g�!�d͒aB���u^Ro��� ��� #�v�t{��b@ ��݄@����!���0�#"$q��tQ�wa��Tp�I&s6jQ$���$�I8��#�$p��Η�v󢦅W�tG�k�8�Β�˻��3��(yE�}��=��C!�a�{��_OW�ѯol�w��<9>�]}�$Q�HŒxb��t����"?0��C�{f����9��-��L����Q��
�[���z���Cٯ��������~�b[g��6:�0�W�N�u��.�1L�n�ݘ�w�:����������V�zo�l]�8�Vk� "3�3����k���&{����՜�ú"�ܐ�S���0��[��n�����8/Um ջW�|�'l�̃���Wu�R�1~�I�ME@A��m���k�� �;I� zV�f��)׮n�� GWk� HsӳR
�B�Imß��8�m)���K��g Mu��@ �y%���M7���l�{�;�,��|I�P�\,�$<qݤt�9��)�]�{�1�����W�����Kʘ��B���IO�@$�	'�`IKH@��$�	'��$ I?���$�@IO�@�$��H@����$�0$�	'�$�	%�$ I9 �$����$�P$�	'��$ I?�	!I��IO���$�B���(+$�k)�d�HHK�B,�������>{������4)�D��� @ H���h � � PP IJ�*��A!�ց� �N� `� ( �U �P�P$zi @(I@� *TQ@  � Ъ 5�)  (  ��                                 >  �      #|U}9jN���貹�G;�Ф� .����m�����97kF�ͩUG\ 9��Yjt�.��󂃣T�� ���2ӰҔv� ,�UMa�TN�.��4T�*:ٸ GRE���KZ�"fԩͥѐ���  � �       ޯmɹ}u)�Ϊ=��ԩ�{�C�'��t$Y�9�U��Js[NmJmr�u�M���NmU٫mu�h� U� �O���v:}z�-\ ԉV����֥u����R�g1�T� Z�J��]�]D�j��ۻ<�*����2��E ��  w�(       �J�Za�iGLK�#���Cu��L� &�����5u�����Tq� .�+�����t�J���  ��8��'E\{�����`.m8�WX���W@� �UѺ�-V�1ԝX���`z! �@��  |        >�����+���S��G � 0��u�U��P�[�����;j4� ڨ`�;�S�� �{�  x>����;� By� �@ 4���=���@t6�� y� � {�;� ��B� <��(U����^ � �  =�       }��9|� � <��=� <�=�  w��x�[ֹ�Ѻ�r�uQ���� �s���� QM4�  e{�끛.�T�n ���;B�f���
� ���*��yGgmC�waN�| 
  ����Q��	�   &  �~F"R�Q�      '�U(d��Ѡɣ&&�#bh�`j��SAJR��hM �14�b��*�3T2=F�&���L�z#F�@��F#I触���F����<���~��}�ZBG܊��������"8�SO�HBHT$[���`��B��?��T�֫j��ֶ�����)������w���|���o����+mZ�Yr�e��mm��-�J��b�ȀB�����c�?���}��鴒$����c4����0�ی��~�>��@�'���+�n����ש�
�E�U�nm�r��l��i�/QLS�r�ܧDL�{2��k3�m�6/v�����SPh�qS�ldQ�Y��fO�5L�˨��Tf}�0BXX�1��Y��4����e�u�W0��L�2�õ�{*Z�֝b��\�!Cb����
�J����90��V��٩�*\�6��w&��kv�e���ԅ^��:1�Ұ^�E���%K��O��f����bi)���EԻCp�յ�t N�fF��_m���5�9x��|f�E.Kɉ�n�^Ue� ���+)��fSYE��j��5.��rr�=�s�oV��RI�iӶ��ݨ��dVf�{xHWZ�*^�Z�n�wA�NU��e��iiM9nc�f\��$)���*�UgFefH��e@��[����47��n�Cvm��@#�7�å�MOgŵt]��5%�H�,�
��ڻ�~Y���eM���L����3�R�����r�Ꮫ|��[qܳwx�8��K*��rI�iRw{l�`Rsq�Ԛ��Z ��Y'%[f�&��Z���əQb
n�J!{y%*a$n���&�ywq��][k&*�(�	�s3d;t����d��l��NZK/ �3vY��N�H���W�{�����AՠĖU	Y7"���.�:�f��
�Y�Y��ۺߵn��ɖ�@�I�&�Y�ȧ+�׵�.��'l����0+�k	����ǉ5F�]��ѕ�3Y�r]��D*�U�Xp3��l˘(��T�qfL"5�%=f¥6�tI�<8r�9aM��G`SƥPz>o&��dޭ98,6��E�&
��v6�ћ��]�-�,�7"���0�%
17j�a�c	/o"e��j鶋�<���*{m��.Z�Z�p�sr�@Vݍ�^틦�Z��`'7����{�@D�q
{;{2Y�f�%p�ލ�4U���y���ܹy�^aL�B�Kj\����d�Y��N	�8���RN�$�j(K
T���UEZ�	D��[��on��w[�M�ep@��B4��b�b�ջY��	,�Y����Cw�(���6ۘ�"��PV�2��H�.����"�Z�ՙ��TL�r��0۬�I��R0԰*w)ko4�������x��Ndq��S��yr�
�8s#Yp I84.�ߑ�N����.��K����l��2KB,�����o�O��f�f���1�����cš��O��e*V�{r��I,<�Y�(��\��sd�n�s�i���s��MBEEǝ�fU��5r(K�d&��&�c�·��$ǻ	�Rr�g����5��^ڙ)%��Z��R֕���3)��5�6�ե���I�d�3&��3M:IK9T�U�^^ &ל0mÓ���́ ȅA�E�K*�VJp)lJx�:��s!��;�E��a�R3[��Q66�kem
�PK�l��{Z�6�T���J��ɸ�v��1����6iQSYvZ���-(��7�4��U�����0�,m�&�*)]�l�bbxcCQԴ3�O3�I
.�:b�Rl^:%�r��U3^�`�v�w�p��2�%5Md"�:�����EY���zէS4�7�E��{WkA9���#
zt�5ҌV7{wn�%[��5��A,�vrA)`8I�b�Y�kom"����&���B%��)y*��Py���]z���!��J���T.�nH]MGv�E�����U��0u�+�Õ��sW�����{X��-1P���ON˘�6�;i����a�jq�U!��W�jC�!@�,'4�N�������UY��Y�Y��B�5�r�i)����%�H0�B��<{���e2���A	vE�G��i��b��L@�zMХrE���t�,��^�n��Nn@� ���e�ۡ3I�HԷtQ�պ��3;Ё�t�]�[�Y�?���n2�W@]j!�/"v�,nؙ�� G2qk͆��un����]�"�h�c0�]ؔRǙu��^�7��N�B��˘V��`dݲ�]�XՕoV*�]��E	(�MV�o.��%GV+.�=e�jy��բ�X��+UDwg��Jp,ݥs�����lɒ�`ԥXL�u=�붥iy�C ���83/ĤNCaC7U�ʫ��h����d�&��n�.;H�~��^'c��p�h���be�/>4mI�����:v�e�(��XI.�Y��w����o\�yI.��U�$"�I�rU�m��\���XrFFe���-�d����`G&��:錤�A�z��J���L�]�X���n�����]�Xj�{Y�X�[����8��2����ڴ�Sv�&�6�O.`�r���@١��F�XN�V}�e�_0�|Q�mh�KG]!AY�ۭ�V/,����Eown�f^Hj�.�=�D8a��c2�~������
KL�i��L�P����#!��jg($�)X2��ƃ4��%In����ʏ5	A�L%g/_�e����뭣rc��k֭����	,JR*����`���)n"D�d�4��KH�F�J�nJB�y��{	��q�LW�А�7X[��*�H�R�]��3k�Ŏ����2�N�%�HY�DkA��ߴ�����
�X'5����+�v��5��F�K��*a�l���]��(;4�wm[Xj���B7���y����#(Q.hz2��yQ��ѥ%��{9���S�U�qCOZ������fF���ڙ�7m�̣0�B��t��D��e]�B5����L�`�,ۚ�{���4Y�>ly�(���pQR00�f�A�k
d�b&*h��dX�s쉓�2aAfEv^^㽽��i'^����yt(P����;��6f�cb�H�l� ���Ѻ�d��^�,]7usR�l�ۺ1ev@�a��m�[Cjm��Y�صv��Q�oK����5f��$�F�������,T�6��V�-�A�e�X�]9���GN0-�0%�:j�,�!�f�]^�a�z�X�!����Ö9[7^bc3B�ɣj�^�,8o�n]^Vb���"Y�*�oa'�YJ�[���n�l�(r�'F�#f�ϙN���a�5tI�$3�[)J�.G���t�\�Z5D7wa���乴�T+Sea�bR��@
ج`8�2��P��F���1ʸ�.Kr*��ݜ��D��N�U�u7/j�����h�y���C�U�0&��.�7��,�ȝ9�#e��vb�7%���o�k�-��;;�%A��\O�[r7��&n kn��h&��%����[tm�ӯ)���XX�tId��h"it� L���ǵ2�ly�n])"�)\Y4��Wt)j63U-�
�`'���Gx#ڊ�f���L��;����F٬{��P�!��3�3-�w�����]v���ڪbuǖ%ɢ�`4ᡖ�,&b��A/r�����h�ua
܅�.�[�bm���m���;������̥��&� �B%1�Z!e֬��I�a˪zL*E��y6���qs�թ-���M��Ҭ�ڋ6�N̽�C2P�Q��w�b
�w���V�ӶJq���j^��T��M��V�7��`��of��l�	��#�u�M��$+v��2��b�^�v�)+!@h��2��,�r�ywm��v�81�� ݆���M�P���黽���l(�X�n�R�����`,�k������+w-�����n�n[`n�S"*j�g`N�s
����/Na	�!ւl�.Rh��g�嬥-5VpdZݻ%���^���F�Y�V�y��4� ��.���{M�K'2՝nJ�Z^�;�,�T��R�f�ͦ��(C�JA��ٰ;�a��,8���N��b͵,C�c�cS����Q��x�p��ݍlCq�
=����X�gd`e�B�"F�MZA���9����QG	B�K0ӧ����}up+�N��7.���XE�5�ؔ!��N�B���Nc���P���qHe�)`L�VCd����͐�Q��2���]�C>��c�ji�2�=�6�X��*�1����ڛHۺ�ג�"�LO�Y�Y�d�c�k׵n���e[V�,�k���efX�IV�-�A^��#���2�L���`�4ٺ��)��+$��	�N����=cj"���`۷O�c%5bˬ��Z�s.�1,���K4��2-7Ga�l�y����2C�t����z!��,��@(�
�-�W/F�d�[�dn�Dсe���1c{Vs0ͻ����N:4��e����RVҽ��:ܷ��j�휢�X.��t��d�{�K�Ϭ����;YN廡�ԹVN��TKE�O��ˎ�v`���
v�CF���`�z�X{���{�\�3D��V0�:M�/%LԳ-�\@��xJ²�H#:�V��9��+��(Y���q�
�m���F����J
�i�]��ءEB��h4��V�ø�ƊA�ɃU��3^|+iЖ`ͣ��v�F���vR�ҩ��j�t`�~{����+�����uI��CIz����L�E)KʺR�i��CYn�� �K&ñn;V��4��������h�XP�/�`LA�क़P�SWb}5n��pNV�r`R��0kV]2�E��,.h�u�hxA�sK�wrqe�jE�Y2Q��"���:�u!�����(o�jQ�3%�T����Uk%�Nc�ƨ�f�������x�0��'$c����f���M�-�ګ{ub�#5�oEj�r� �Uɖ���@(ӵB���r�S�P�:�/$ɵ$�P��5طN�UfC ���Bطxi�d��p��6�fL�ssn�0%�L���j� �n�7�*vn�����j�I����4f�aC�iK��M�,��˲7�n�B�]�ӓ2�Ki��t����^��\�x�+A�.��T �V�1�S*�=$m�H�Y B-���#�Ӻ7�Y���V�� �YM�j��5uǒ��D�82�6��)�y/S,��9zq�n�Z�:�]�-'���4�ř�F<�����֥e�13ynb��úҸr�CC")�	ef+w-��\��Q-����benѹwI�edT�Y���(�G,`{`� �I��ըҺbX��:��G��!����{d��s3o+%���~(��wu���+N1��J[����Zw�aiU������Y���"&��m� n;2�9S*l�T/�ŃP��`���m,:�U4gK��G+,9��CA���c�E�;Z�+
�ʷ��Ʋ�+�YY�h{���ʷ�3a�f�TkUkc45��lJ�$��X�b�<�2)��jZ�Ez.�+�s6���JQ��O�j��#�	ųv^�)<�R����um��m�0�MqT%��6�v��j݉Sw�V^���R�7u��$�̎���3�f��JŗQ�t A���T��FAb�˵I�Z]:�浇M�J�7�ݡ=a�pT�ye=M0�j�1b�1��������Ǘ�����U&�D<WW@���U�؂���oB,-��T�,ˀ˅��e���`c��с5E;��C�,�wi k�C@��B�w��;�Cj0	Uf�X�XJ�u5hձ=�n3Mi�O%�kL ����J��-Ѽ>%܌�2L��W��
!��Ш��3(U޵����y�-�$�8�C���ZE�PBdlZ�[t3cяE��˳�5����b���A�x�7@ǈ��,�4ݼWzKl�����l��ݔ��9��~ƪ���	2�4�z�h�/���O��Tܐ�V�3��S*-ōS� �7"1[@��e�E\�SA�Iۡ�4��ժ���TL]�ְX�PI�1jYr��{���&+y�����%jB�\��NL�v��,�p;2��X�-�Yxt,����r-��ƩK��ȗd�e��5��6<�M���[��s7u����@Yj�ceđ�sE�+0�b4E��0���E-<����k�/1,H+��55dn�^���M���{��Ԡ�j�סP���7s%��t�f̧��2T��Ŷ30}��b���hm��n��`���)�yJiD��N$^I�Q�c�J�=��Y{YV%�������Yf��ղ��pC�@��c~I��f�[�ْ�����!�x�GKAۅآ'$]8��vC�1���#-	(b�w֞Ţ*!���Hb�
�fe���p�bGrc+wf���~ƾ���+O��e�L���� �C�#Ψ�_V��mW�-F��Q�b��5[�Z��m��V�-j�mW-h���5�ܶحnkUE�m��ۚ���V��F�Tm���sZ�wV�UV������Uckj5�k[�j�+b���h����Z�lmZѵ��kmW-T[U�V��6��\մmEU�Ulkm��Z�Ʊj���Z��j��V��6��mh�E�cUmrչ����j�75��j-UՍ�5[F�5�h��m��樵Qj�Z�r���Ur�+m\�lkX���V6��� F� 6�6�����O����>����D!I	��cY HI!z��H?B[?���5�~�*��WϿ7���m�{���v��y�����痂�]u#wa���5�����0k��#���d��(�LY������O!�٤�=�����=yov#�b�޽�F���.�$����h�v���4w,yO��(fȆ�pNP�z�[p`8$�r�3x���$ᛉ���l�t̥���!�g�7�2��\
��T�\0�j�e� ��8���/,U��@���͉h�E��?[�d��m<��3:Aڕ�+M���̋^d���d
l$��fg'�KB�^ˢ�#�v��R3�to���칙,�fe����N��Ń��ó�mO��c��b��%�� K\��B�/��9\o)/6�5X�t�*��'�X���؉�hMN�����xv܇$��s;����u��ld��3V�L#�hbw����eq۫1�u)>Hỻ���w���{�uq�Qnd��k�㔗�Fof7��E(-D�u�q��gB��"N����+�ǫ7f���x�
Cɣk��*#a���>��k���9.[Y��M�,��K��74#{�����H�r�ktL�k�8�ǝ��nvgVk�bgfo��S�sJ����w:���n�s��ە�붷D̝�}��D4�M��ʼ�Hn�ڔYԝ㈈�.�S��Ev�'j�T|��lׇo��5��q�&70�[��1�r�5����K��t9z9e��tG�^��� ��Ne�}y��kaw'l �'�9I���\�6�8E���pۛ�0�5i���Aa,�J{8���J��֥Պ	ɓ�'ќ�on�F�d�i6��V��z3�#
��ƾed�v%)�HY|�u��f���㫞��w]Υ�u�+cĭs��ImUS�5�}7�y�ԏ.�>ᔹ�w�3sFRt�N��F�)wS-���D8N�tV��s�qX���ԛaٷˋ�tiR��!�N��g$��	��݉���b.+�2�uc�,�z���d8���Dm�Ƀ�����cVn��������3Ԥ�8��EF�I\�v�2�4`�u�P�ge��׸֒�_v��`o�AYvi������b-�|2�WNxG<U2�يý�r�m��'v���kAO�wZ�ov�S�y���ܮ1>��0��cA�з$����U�kMA/��>����k�2�G�:�X�V��6��N7Y���V�OA�M*�����{2�d��gQ!k�`tWS[�6�ɘ� ���73��`3MU9�q+&��FK�ܻ��ON]�p����v��^�މ�m3��X�pj.v��=rk^m���u�|[�:���4n��e�o-��f�`7����f��v�+�k���y(�ѩ����Y�^ћ�-#I2��:��v���'Cqsx��8X7O9��·o�%Ϣ0��6�g����\���y�ןj�����.
3@�k�g6���H�n|���;pT��YV_/6�D��1�	w���x�n,�`�����yԌ&��TrZ���)���]�/���6sN�|:�D�;�D�"k���7�4�/c-��5�q�bR�ϱ�Q�˵B�֥���Qt��o"a����l+"��-�4UJ����x��zG�⮨�;��43�f������e۬�Y�,�_<.�Vpl]�t�%���E4l��_��o:Z��q�v:�W��P��7���u����+��V�e>�`�K���-y�s��i����fMR�Z(��ؗEf�̗��;n��ۤF�-؉��֣l�c�y$[f�'0�Ф[��I��)ͩe�b���ۀ��#=�x�/l�s3�u�k���[�&D�H� ;o�L�+�+o���Z/Ґ��a���ȵ;5w��G圗[��Q�2���@��ʳ�/�%m��w�l�f'�9nQ�8-QP���B��W�8'\��hN�*K*�L;r�C8m��^oso�%XoU���3E�������ʺO�8e�'��(aP�:A���v��RlֽR��+S%Ը�-̝RΘj-Q�-ǵɣVW+�ݪV>|Pc:�ÚG�\���}���`�v��=oWajc�&�s/5ew�/E��2G!�Xrm���� ��c�3Y�.�����N�A6�і�*X�6�����S����5�t�����#*T6p3c#�[�gS۳re�ҕГ��^��\�LL|2�m�s�]u�.��oI:�Ģ�O��5�W\��RyY�z����!�!C�n��`�M���wqU�u��ѽ��A����B!�M
���!�r�y�k�7��5%%b���_<�1�)虦*#BP�*C��[5z�xҞ�'rW� �j�6MpS������L��1wB�N!ݖ5�橹�*�� ���ywp��cŎ�/Ws�ݰ0�;\�t��9+�����c<m6�yR:Du�-Ǚ��qYZ�����b�=������7��uYi���Li��b�g_نr�#Ik:v�:5j�t��Of}�:�m64|����f�r�(�ὪSs��Yl�geT(25Z��>6v,��K����ⷭ���h��B���Ã��r��f[�5��xX�n|Z*�༗.1���K���E�a�*����ޝ���'��������\�]i[�b�����bBthYVZ+Zh��"�t�Q5����?dt�GJфns�ӣy�����P3/Lw$��]kw����Z�%2VRݝ��ɕ2Ӂ�N��Ip�&^:t˗u��-멙��-�9�8�����(֞�5`�medf����NΦ�e�o�0αФ�	Y�����=�z���/�u��p:O[�ׅ1����e杒��'Ϯ�,Wt���0�;g�;�`��kXj�g�z:��7�a��ႁ̙�}�d'�	ph�A����td��Dr�ܫ��G������@t�!���q��3oK��W���w �[����u6�a"���6�R�|�2=G9�)EYO� �"q�wg���/��S��n�^G�vn�2��2�"C:��J�r�;�][c���yu+6a�-
ܼh�:�IC��	��:)Ƈ��3���*��9��t��;2ò�5)i�S���vFq�b���{:l��+SL-ۤ�b�� �D^c<"��b��rU�͵/6+*�y��N�(��/�su�]Aܺ9�5�e�*�k���̰å��k�sĘݥ4�^���Pzݒ� �����-WKM�q�|�C3eN�67d⫳��=�<C�t	��ȀoH�%YХ$�̎غw�5ye"C绒�['�i���Bh�E��t�
�����a�ժb���sC��Q.h�v��c�K�̫<M�S�o���Y}}��t�FJٹ��p5���/�x�����2�m_f>6�C�2��^!8dj�;|�r�Dnqyb��"՝R������{�4N|�v���oJ
e��͖axY�ܷ���V�bN6:E��lN(.��# �^��Tw�.9Ym�x܆��ۛ��Rۛ�	��NL��Ӈ�y�o:)���n���N���.��O��"�8*U]f8$�%7����fk/.��"4l��S:hv�W��vG�3&�qfn���tAǊs$(fE�-)2êڱ(��:��̕���r�������}Ef��6���Ӕ��y�ø�?�{1�R������t����^��4t��.Rƪ��
(���dL9�p�����S֫��$�S.v��]yDn�j;����b��b�V�k�كk�ZpFѲ��EN���4�wh4+wF������[5"D�
��\PGp��΀eZ\0[abV���{DU����P��T�@Fv��w'7�f����-s�	�ٜ+T��Wm���lGZ��D���p v�[��E�\15��B�oEE�3;�&�a�o���6L���c���N���'��Y�n���3���(�6����̪��s]��Z'V�n��̗�����Q[�_IPT��T����yŚ�E�uҼd�Q���$
���6�e@��Wݝ���K�'���MT;�3j���Z���<��<�́�^<������vd�}�\����}�2��(E���ªn��ŵ �~�!����5�(w�_^^뙱�\q��p�|:�ÛL��*���+V�wQ˕�K�T�u,ۡң��U7m,�x�.�#M���c%9��v�O'Xtj&�YP���dOu��7�'jY+h�tM�5�H���M\�YZ�Y�ݲE����Ze�u�6��7�����E���Y�0��;���m����Q7�<�9�Kr�^��:Ԫ�̓A<5��'(,8�H�NT��y��5\�_*���K%yQ�5Nf���,���lKܣ�N�a�ζ�'Ru:ڝ�jA��&�s�t��dRL?X/Pt��j�k�S���*E���PNnX�;�u`��*��Y[�bsl���=�y*��W!���x�#̗�Fv�b����ݚĝ� a�}ϯ3���:�*]��"6��W����ZC�D�v�����������<�'�U	y&e9G���:�b����ͻd��m!Թ��ɐ�X�����W��KA��nvu�Ӊd M����3/!^L�L���G�3W7X���h������v�M�u�z��%n�;�]ܻ=��سrz,��3WO6��8GI���s�p���-˰3*ycT��"]N��k�%T�fs+����j�2�V�W,S6�n)Փ%�']-�{�t��;M!V��Z�qX�Q�s�Kͮt��&�|�Ω� �)�m��,���)g]wC{�����E��� '���F�5{W1'!z�W*�n��)�H�pˣ��o飃�F=��5�5a�RIa~,�VJ�6�wue,vxᙃk����I�}�[�d�Lr�DA�8������oWf'���sZ�26$V� :s���,Z(��R|�O$;Z]ư�klvŋ]������Q
e\\�~�s�Ý۷��N2�Xa3�v-[3Fq��M�޻"���ۭ�����+�nMT����ܗ5�#s�l��1�`�XgT��^�v�]]m*'��3����pS޺��d�AkE۽�.����9Z7��� �j���v���ܗ�����$����OO��0�i��w%]��@̷g���C{�o�hr˩*u�bn����
h��H��u�*N�e��@x-�f�۰Fآٮ��W����M\E���<C���������S�gqb��n]!�И5!3sR��^���nG>n4on6��3N��Ư[������oJ̴R��{fm>ں���t�Ϊ�Ɂ%�̑�v�V�B�Q%Z�ǒ�uUw8i��:`Y;�w�`>��q�*�Qw�ɫ��
mc	�KE�Eeo(�(V��k�d�K��a����oP��S��uZ��Z�g-�>����U+.��r�k�=CRvcXzP��]q�OY���R �PYj�㽫�p�Q��#e��T��Lik��w�[��V�Ce9�{�:�q{`lK����@�)�����q����*VZ��kuEW),u��`��x��ƸޖOA��)T��@M�evM�p�Ĥml:�7T�>��C�י33�V/�����=���Ͷe���sf�a��0fg0�&�-�53;SM�V��4�gy�1<X�.����s�)0;�k��a�Y�U�����F\��6�f��J�O�n9R�S��q�$+�Y�#�)�$s]g0�*�`w���T�׺�Sn��O���Y�/���(.�ƌ�ͣ'C�Z�603αQ즎���A�nul�.��ap*�6���7Ow��s���k=Ƅ���Eچ�ZW״��
i�n�%�wWo�@v3}#诺�uj}��F��'}�Z��1��bݟS��Y0����$"�����b��D�h,��_ouo!DmY(<�sL
�{�S}6$��g�E|��2SY׌�A��0:�83��YJ�u�/ssNd�+�.�,�j��4��p_tW"M�׀Nĸq�A��un���`�~�2.kY
�U�v�3/��ݞn�}$	��]��<�n�Qn���X�Tk�k!�`[f���H_M�Vu���+�� ���_EԐ���9 ����{i f�(�mC��cy�D0s�zs��}��_�D�����'-e�̭�]�fp{{�a���y���v�_-���6s���2�ÀL��{��e�+�Q�	Rއ7��s��a�p��^��9��X�ue�I�V��)��N�Om_مRP��s.1ݘ�v�[�؉�Yz8�IYp�_>�g^�Q��P�T��o9=�fJ�:��)�_i�𓍎w��e��֌gU[�䛌ԩ��H��M�R		m�h�/�"-��~z��Zzr�@�q��^�����s�Z�1F�ٽY2kv1����<qqk�йz�۷\��C�	��vp���mⴜn΀��T��P�g=m����6F�c�t�\�MLm�f�Xy��zNm%Ʋ�a:��϶zP�&
v�j���E�Vo=���B�Q�������/V��.r���㣱*���w8.u���ʠWr���f5�Ͱ&����<�v�+��Z��Bջn1��:ur���cu��M1�=d�'K���%)�Ϯn�v��l��n��F���-��:xɆ�'��s3��b��ܺݤ�E�i8��q�Am�������W㸢�fa*c-����^h��v�ghX}��=�_7s.�v�u�8��NAk��շ����G�7[g%V�c���n.��Y�Oah��g#%�������>{$��l�z��R�Lq/.6[��-Ƽ�8x�m����
�=��s�$a���'=��{$֦���	�8�M���y��V�
&z�d8�r�m�ۯ[�מqs㸷-2pl{^���v�noF�O�c*��=����9��ۤS����y�[��c=�qi�_y84n޹�[��k�Z{�n�T����>lp����8�3g��v�9������]�ڞ`9�+<���!pv:�{�pU��U��.��e�ú3؃s϶����O�y.����8�m�J�У��eǃ��ۮ\��(m�cy��VE5�xqΧ��q�ݮ]:ۂ8
�e�ӫ�v^y��^.�\�c`�y6��hs�mV�8+q��=I�n�	m��Ӯ:�gr�*]s%�a��-�c�ܞ�I�!p0nWf�m���t�$�=��͂�]��8.��:`��y7<ػs�K������nw=�-��M���R�K]����6�Ol=�s[�^��.Ɏ��P��j�{k(3��7lv�-��b�]�tt6x�7I�p�p��
�a�B.��vC�*�2sE��z�6\���x�%�ٝ�Y��Ͷ�S V��:p�pn5���g;�<��������-��ƞN�s� ��k�m{s�����P�m��sX�N�Ƴ�>݋�^�v�֮9/lύ������ڹ����2u�ޮ�(�/yg�b��ѤAx��N�`�>���TfE�2�җ���1(.����]�O[v�BN6x'nLϡ4�t��\�<��i�s���lf���V�_\��T�-�q�@cOi���p �c���<sC��A�ۡ�u�qfk�î��ۜ�(=:K�%O�:x�r��'>���E���i�}n�%�tk�]X5���P�Mӱc�]��v,�=�7�<@f�g���n�;X¥:k]������8_FC]=@�ng��<ge=�N�/>��c%��l�@����k�5�˳%�qф{��Z��N+�w�Ds���%،���2��Ba��lv��ɭK�֑�{1��ƘL<�"���Uu��q����f�q��������h�����'=�ƺ˶�6.��;s��lG��0lTm��w���X�A���gS<�rsk��z�ǛȀG5g�����Ɯ�[qv,������f�f˂|	\�f[\=5�=��2f�M�k�۴f9�3��K׭��z8�9y.�f{^صv^�f�����mm�&�\��v�tk7At0p�;�K�c����W'�����m��#�z#>�{m��73�8^x�)�� ˙��n�0R��ۦ��ؗY�q;Ƚ��j�Wm���͐{FeH�2M��s�6��|v���q�q��$��r�� �-ֻ�[���v���7��0�Q�un.��%���v�&�I���YΰR&���89nP]ݐ�2�+u��3��y��G��<�=�Q'%�{]�Oq������g[���a����D����g�7o�G�۴�ify�[������+X^�����N�5�ϷH'S�#�W\lێ7<�� 眽�͕Q�k�՞�����Wo�6[%���*Ӯ�`�����И�q���^퍆�kn��<W$n�Of��Y�vJX݌��HA�@��z�r\u�tֳ�ce��n����=�hM����\z�W<���Nle�z��lur�!� �,���\B�ă�\�nHMq�&�	vw='��m�n��Ƀ���!��=��s��4V��qkJ7X�臭�]��ׂ�\>�kFP|r�u�(G�)��� acb�Ul"�7nn;<b�����'��/Lc�0!瀲-��J]�kub�	���z�'�Ԧ�:�������Y�ڀά�5�vu�T�K	ƍl���
v{'[��;s��S&�n���s�u*��b���Y܈�j���|�i��h�����V��z�CE`8��j�������9n����=֬��3������q�ʆ��\����s�m���9x�}�/F�&����g����/;	�N.�V�'�5���qԼnB�.ٳ�S��uΎW:m��l�-\���k�Sr�ݸ, ��M`ޞz��-d�\��m1GD���2A\W�dNq���l�#p�]���;n��r��n��k��&A����n��Q��=q��������_<�n��v�]�s�'mћ	����ɞx�읲f{z���v�q�xh���9"�uc9�y�$�˵��r(���/n�of���c8�,���n�n)�[�v[h��3۳ۅ�ne�K�D8�O;��ùv�tz�nu�mu���1�F|�]�v�A�k��<�q�v�]�-�h���MWO5�3���5�7gj�nƇ'7NK-��4���+�0�ۊN�]n�h�ɜ����k�������T|p���%큎�'Y�ovpi7�m�8��#�8�.۝��ظ]Ⱦ�`�<�y��%a��.Ќ<��I�9i�=8�sX\���j���k�v������&2q��OEcm��VW�`�λ��8���\��p�����1�ǶuF��vY��Ş�m�s��n3�v�/9��!�����ג��8��7g�x�-�䗁*Þn�q�8�>ۉ�d��k��9�ɰ��gH	<{v�s�e�n�v�y�v������1y-�q�-��ob�]����厜�VK����N]�tr� qn#���OU����Wnw�s��3�<׬�۪j֣�:�Bz���`py����6�LF�a��ݸEڹ+��7�޷�c����٧��3(�1�gv;16�d�w&�py��pR���k����q�]/M�=���$6�V���s��n+kl�h͟�u��N6O���nvT#>�˞#M������S�tg�g���K1{3���u{m�q�q�������=���	���D��l����	탨x73�D��_'nc�����g��^��B�9CnZ
��LCD��v�u�9u��W3���gFP��`��ջ}"�ka�n��1n�c!���6��;���=��Ceb筞CHj��8a��iC��y�v��%8uȼ��r�}=���=!�g;��nÞ[�1��� �m���&��m'g��W�v�s�[�p�`��ۭ������(ƺ�jS�ۢ��[�
�r�����.��Mq�ݛ��q�l�S�cm�p�3\�t�vs˹lz[�a3��G>ݻ<�:y{\{gS�$��7�e�L<v-�K��@���y�9�k�Zmoe{Oh����=�[��=�c; �����v�x�8�a�k�n8K����o*;U��D�Lu؞�86�%z�e���hl�q���rH��p�]����4�е@V����le�7�C8Y�³��P=��z��U�v��b\�̏Eۥ'r�RV;n��ڴM����Y�W\���p�6v�K�ݒ�9/]!m�<uzrIY+s�mb��t9�`a$r^i��!�������:�7nMZuv���8��%�m;�&2�d��nW�����k����^-�v�/������]���;,���y�֤�q�f��9�CH�{{3�#���c�;.74���G�j���1/Y�����	������/m���Ж�î��f7��w\�M��M��h�NU�`�U(m�۳wN^�ڱ�b�ng�nq<�g���+�V�����oK���m=|�]X���v�0���m��[����3m��w\��u�d�z�mtc�x�+��5���s���q鋎�z�ڍn��ԫ\j{q�Z�l��eݱ�����ϮEv�t���Ny�����9Î��׮my3���鮊'��zt�u�v�%��d�nm"�-�9yn��OO=�v�gt �������ٖj́�8�A���8u�E��p�&¤=u�[pq����n�^M��n$�#�� �ۄ�.=�f�[v.�pwn80��w+Gc9���u��8%�G]RR��K�gi,��ݗ/����ߍ�K���k�a�Q&�
a���ƘI&� �B�H��u�2��G7���'.	�2���!�ɰE���C �!��1�%�L���FdX�n�,�&���Y�s�A�a��W*0#�tl�(1�A!������vΆ"ŉ�@��0$��%+��&R��2�3CF��ܷRM��!d�H�d#ݸ�4�$Q�(�C��)6�)�Y#&���*I)J,`��i(��&�h�X����b�*1�$��/����s��lpTu��%��"����9��E�'x��>�v]�n��|98v�`�-o=i��<V�؄�-�;6Z�Ǘ��s�=��ڮ	H��n�kv<s�����	�hۯ@ݹ���̋m3ǛvyE�"�Ƹ�j�즞;V�x-�x��&Ӵ�竴�nل v1�m���2�B=��h�ݍ`뫘xK<c�����gEȽ�'�`�w3�wk��nt�+����f��V��e퉳Ǳ�Af�o^.�a�D���:���U�o ���'݃lKk��E�E��u��<5�,N�!����t��u�"�8ym�c��ܼ�x=�&�.��^��&�F�^�q��|{�p���{cN狭�N5{pF��o�p�`8>mѳ�t�m�@��wM�϶zC���2C�5�-��au��6���7��=�L��:�}b\f����4@v5��M�Ѯ�m�l��-C��n.>|l�q��K�,�C;Z:��۠���.�hq��wV-ۀ�)q�1�u5c�/uZݶ�rvN8rm�2��˸c�WY������a���%�Pp�2�����z�$];tx��.M����!�MM��j'	���Z�r\��E�N���g��xp�,��4���箬�q�2���jK{p�:u�z{i�T���0�t��8<�=�x�ˍ0vq�e�7' 3�t��sڎ|�O��5�q�=�ˎ��ۣlea���w��o;��9�ֽ�+k������s8�ݸ�36y9�gm�M���*���vö�g��y޹6q
�g�q���Z�-ڀ�ػ�]a���ɭ��M�]6��%+���]�\z��s��Ō$�y�uDf�6뮙˱u��ݚ�+r�	�y�����e��o`�!�y�Kn���9���x���)�r�r��g�������9x;��=�.�n;���y�{l��w��n�s�r7{�ˎ^S�l�s��d��N�����o"�]ts�=޽z�=ޜ�Ou�:�n���=�����{'.{=��p���9]�92.Ll� /c;۶�1ț<�\���09@	?��O�?�E%�HZ�����oKI��ܔ��/�~�!�.�ެ$���/�@�W�J=5�!<��&�2���O�(OW4���������6�� ���H�g�8�u�yO�t��j.z=�����\g�5�m��sKMD,�H*���|��qq�"ň�cVx�/zQ���"N�v�3{���}��b}�,U�
��׮���H��z�]�����R���onQ$�]�Nf�ݛyN1���G3��9yN{]`�OD�G�|�_���v���]YJ�n��)��O	�5�F�di�s�$��^#3�i�̝b[2g�$r8��O�U
�rD&�G������6'g����dL�����~�81�k<��i�ʜ�ҝ��+9��^<7�-�u����b��֥nZ_X�[���/�MS����]&�O�V�@Nguݒ�����f�]��zu6�:�h~�X�\� ���mݐH7��*�&�t�}�i4���}��޽�,A-�!�=�4�R1A��������|���%��}��>��L����߲8떠V�wRwd�7%\LU9���\!��H%��b�=�(s>�$�U�Y#��m�v�ٮaӱ�\����V��b����96J����TA��^�1��"�u� �f܊�r �~�=��"�z��>��תE���U�/St��MMb> �{v�
�s�@5�� �cJ�OJ>"��BU��s��o~ȴ���4I�ֹӽ�׫�5�Y��5�I��ko�Ő���Kx*6྄�Sw�H�=ۃ++u�1��A��̕��F�	�t|s|�O�o��X�^7ܚmlu�gP�dT�����A��98^#'/l��r�Ak��pסl��ՂS9�1"[C1B{�I��w�h���{3��	Ӎ�V	%�u�$����X;����͘i����x�7ml"l�����Y����p�*u��n.����RʅBy箻��'ǎm��GVrG&U�힓��+˻$��ۑU���&��5����|X2V�P�6js*h+���	 ���:s�@�әdI���p�D�hQ��T�����|z�R$�´չ��쥚	$dc�@��՜�D&�_*��fbh]����6��>Y �9�!x�:�R$�ۖ�:���*f�j�hIs��C��w�ol��=��,p�XW��
��ɋ5�K�X¹�PvJ�!upF�P9v��ۡ>���^����WJ%���&0DA�T����H���]�Q�.���(���Ax�f��٬�91F��~I�ֽ�qwB\�v.����37hۣ1X�H��z.�"rX�yBs�i5˾��UN�F��~��M�{-P gr�	��M���	��]sX��MrhF�=�*$��ܐ$��ܻ�\gC�ܺ��#�U$��5�(#>n���P�� �e�h��J�PYW���I�m	9ݹv4X��Bj(Q���f�S���{r�O�f�{^�߉ ��ێ���tj�}S� l�� ��H����Vfe�ټ��_� 	��J�x�Q��hgwԉ��˲|H인^9q���v��D���,�!SLhu%�kI��e�MYQa�;3;����|��yv?SyO&0ie^E�f�'��k��A\�����O���v
q7#r�(�T#�S�v<���k��f�0m��{q�g���Q��;q��C�#������m��6��%1ˣ6^�W�{8u�t�A��g��+��R�"��!Vq�:�^S�n�t=�S��7!N2�;��n1Ջ�;;���n��<�f���/��C�����ݎ�[=c%�����]�S�Z�NUp0���m�c���`k��p�[&�;[<�cVI!.-��l�߬Vy'��k�4���A ��ۄv��vú�	?{���f���eda&d��4�}�d�����^>��˲;#�&��u��=�"y �U@���{�5`��ۄ �3�kagM+'��>˰H=���d�H� ���]��\;)�QrO���`YnF�/A�Π��n8>�у�^����sy���T-!h�Z^ټ�	�۩ksdh�L�]]�d���ʡ����Vx��|��/,6j�ϰ�9�ݺ�u2W�� ����<�<i��������G��
�̻�7����� f��}<�,|9����f�6�����`�э߬V#�ADop��\cm�mTڐ�@ڕ�el!
�Y��t����i�vr�7Y&���؉�5��^��#��l��Nؚ�)�K�y�!�j���}����^�����e$&�M�%�R� ���{�.�ZA̝�@�Hw:�� �U@���_Rz�sf��ˍ4GLn@D�9ܗ��7�/s��&\���^9��$LI���r�"C}غn��[�x�t��9�A��VH��Nw���m�x&�W)����;4X��p�1Ҧ+ ��Z$%��_�=HZ;
׾��٦�������6,?2��<����
���s;˯���j[a#�f;=��vD_2��A�.���L��^$�v����g�j�F��í���#g�7~�X���Kė�r�d��S�w5s�F��H�^l�C��]|d\��2EqE����iW�훔2<�77��n�=3/Gh���m+/f�� �ﴴ�߽��(%�l�Sd$$���ROv���rq� y��}���{:����Ê��0��E�D� �P"")�M_��ٲ�f!���'*�/_>˲|H�겍Nd=z4EB�L��mчI7[X�;N��]�K��vk'N3_?;�1���1^���\��#vX�I=}VAv�h�۴e�`��Ax�we��E�5l-�kK�˷����$Jr9.'=�Zoz7� z{ �C՗���� 6�F�ؾ$MULL��w�Sݖ,�A�f��/�$��g
n�yq_�d�$��ޖ� ��m�Ú�nu ��+��=쏯���my�D�K��h�N���F{|��}�	�߻03}�3�y�F�z�{��������}{�	ϲʎ�-�UG�m:*vi��=���^��Ӽ-����@#�=#��J8I�O^>` �ϖg������>=���@ ���2	&�{|�3k�*���H������X��mͮ�%��cC=YƸ��uͱ;.���Eޮ�{�Nښ����ӲTɢ@?g�ͺ%zf{����I�/7˘�@��]���� :���;��@{3Ɇ=�d��� �v��A'oS�t��/{ӣ��$��=�c��u�}�]�,n��Ř ��0������D�� #=�Hf�/V�	�O�/}���us:�w��$�Os` ���c�g����~�]n� z�q�n�Cs�~�\���M�M;�cg==C�ņ"Oؚ�� ���2ē��R��F���^�f��5�pu#��r��p���FQv-ʱUW�blM�r�D��
��Q�8:nPk�;R�����V.�`��@]�3i�k��9k��텧��7ۧ���]Rom)Ny�y���s�þ{-���\��pQ;��rRr��\C������z��c6�G���w]�rp�盷F�0W��2qs�9_r��;�	È�Z�5	(ţ�3ɳ�m�e�\�n][�5�z��v����.�vz�B)��R͞)���NK6
���m���H������j�]!4���A���$n[�x��p	G	;��]y����{Z�	�s	[�7���&̃D���ٲ��4(fe
$��7�%�5wf5���w��0�$�'��� ����t�!W�Q�8L����g��9"/�M�k�Y�F��?� �BWv�껜R�����]���؎s۸�^��a��#�ã�E.7�D4I�s��6j�?N��0#�٣^��px���M�Q鹡�m	�$��� o~�zw�������O�{�tI$ѝ� o���/���BjV���v�[E�'��dsp�;��ݺ��n:�ilɺ�+M��?_�ݟ�^����'9�� ����ŀ� /o���Le��+�J��=�mw6�$��� l��pBf�]zx�U�͐�uz��O-��}EK۬<s�ea�0D��	���O�y�哚�ζmTN�A5b^Q�)H��,�)�N9z��d��6$w���O����|�}e�h����d��n�-�mM3{Z�Ńg��������z�v��֟]<�$����$�������0�f�^}m��P&0�a�Ld�9y���	'Ӗ��H�o����b�^T[�wďw�'D���X%e��c�jЀ���m�;Cޖ��Q$����N�� 9��l�{�7��ֲGt�0�J��#����n��nܷEOpں�`��F���_s�'���$r���s� o}�x�l@]�٘�H9��v��_n� ��\y�\��i� ��r�N�سػ}3َ��oo0 ����Cd�h�����h�z_�75g�s|���#kЄ�����ŀ�%k��w	$����5�-{�6�_���c8*~����b��kSb�u:�ܙmf�4�甛v�Kp�K�sD��~5[��v��Ԧ\�Zl�Ŷ��+��hX�rVbC%���j`�=�e���F([���ɢ5��y/0��-·�*�[S2���:
��M�z๥���<�I��vwj2W7�=�Ko���i.n��퇮�/|���j������	5W,�N�#�dS�9b=O&�cy`>7WL�w�T��>=����,�B�	V�8e$d<+C��J�Н��0h���N����%�mpd�O�3�u��;*q�!�h ��a�$���N���s�i��]w_�z�_�B�W� �[u�<��/�-��׆�̻��5�q��g�饣;�Zki�yyۺ�G�9�5��2n�`��|�je0ϲ&�n�p�3e�b�ݭ$f�a�kl\[�j�Cuvz�hNJ̫<1��J��X��bN�V*`�,N�����s�X���c�7&��>ܣ}3[�F�5�W�d�wn�b=J���h�P��(a7�[���n��l,�c4�Pz9r]G�oy�[Ap��o��Nf�u��tg�}�38t|30m٘����-���8��(:{������t�ּ������F���ݹv�������Vݞ�C�ƚ��K�)���c�a哞�!��7�6���3j(��~���̒�Ԏ�÷{�2� L �0�[s�w�F�`X�.V��yB;ɒ��柾a��a���hLi�m��6+�F�F��A��CDAwtcb����(�Q�S�r�6(���nF�hɀ2e���%�ו��d��-˦-�͌hܢ�X�Y��r�w6L��w�����5y^jJ�b(�����)s�K	\� �r�1r�ws�m��y�y\�����1�p�%�a���W�J���:HѴ��0ȣ������;ޫ��9�u�JcJL�<ݔ���OB�I�^��uh���A"i��7�F&�HcLA�G��s/��@؎o�����Mg�7�pq4쭌s1 ����Y�K�]��;=.�o.<�� .���_�m���u�;c���42��E{��5�w]�P��f��ϮBy����D�F���d�&�,��W�9�u� lE�}�� ����������a�"�,�H��b�Etr�C|�z>es\u��rKT����e��?F��G^��fA��4H��O�M�}��)^N���+�v����]2	#'��̝�TE�`7b�tr���́,Ò��{N���i�d��'y� Ӿ���H���~�>�CKq�7�J�2�D�H���D�rW����i����1��y�y��u� y��`�99��Ā��������o㗞���z�0;J��h�{˒��}-2Mh������X:���1��A{Jߦ�����y�G9���M�(�s�d�b�Q���joYźa�/%6/�����s^׌!�����Ĉ����-D�����Z1�f��f%����gm�e}gw��z�{�	Ku&I���w�*$���"�� ��8+�D��uv�^L�j����ኹ*�N���6�6낃p�3ݎy �K����g�0@ ��nbX =7�L�{�>��Y�;�4�ΤOo٦����&b^���r��)����l�|���75s��=������0 M���9��L��=�m,w1��Y#�c��{s0 �6oܚxI�m�qتg`��ػ�@>�s�� x�ܘ��Ճny8�ˈ%��w�s����É�h�w4��=7�L� ��wE�'^�{��I��˭����7Uo��p��� /���3�����w����g;�0 >=7�L� _{��a���?ߋ��;�?څ�7
>4�&���t���|�WvJ]&�U*Y�N�nfjv2�ߩū[�9^n���ܓod��.j�o��ͽw�Lw�AV6���!�y����v��&8��s]V[���v��Q,΂��u����u�Ź7�j�kc=-��ޕ.��j���\&�s��82rv�ݬ$��pۍ%���J�&��4��^��N)�l���6��8�m�e���`q��v�m�:'Vhl��ѷoV%��qv��5D�#VLWQa�Cn�ܛY8��U��!��&zold����V�Q�9S�F�skg;*�h ��Q��Z�<gm�I&�5���&�;�9��m�TI�I���A��#g��H�;��wY��R�_1�����8�u�m�I$�/sl�J؞g�7�\����}Pz�XA�c|zK�d�I��6�Ēg%D�4�ϽkH���I�=s�n�� ��M����C��H�X����gu�u97�ηL��$���tI'v��x�ud�W'w;��e�L�^��&���Q\��s��͒I=�̺�NyB�N��Q$�.�f  G���� >�/���NN���s���o���q��ƥ��-R
R�m�{t�
j�-�=s,��cqۮ{Ѝ�;�v����o::d�I���ͲI$���e�'�D�3ڢ�73Yl�D���N�L�h����-��,Z[&���@z��~
O ��sMW�m���m6�Gw֦hj�쟡����ʼ���)�6��禎��9�[5�M��w?Pm_���I&�5��I;����&Tʳ�r��zl�C���)"��^^�,�σ���0l�w��'�3�I��G��� �j�s�f�>�;]���4߻7�Wf�29���$������ w_2�&�4}3t��w���$&��&W��De�vS����$�L��P��sc&��oW�33 ���#ۼ᧽ۇ��f�k��6e��I,���S��k��P=\��؍��0{]��cd���O�S��Q]����f6�{;�,�n�bto���7�e옷���m�~'����5Gg��o-��� �N��}rz��w�Q�9��|���ɦ� {w�1`���v���yņgM�-�c�~-���}��&��O���͵���e���\����B+�M��xI�^
�t�ǲ!�1;�<iL����J�c#���M��y��;�����I�O_�;`2I�5hl�� �"�����=|�NfҾ{^{��e�� tI���CQ �>p�K[Y3i>���EzZ��cj�X3���ãݪ������P�^Fd����ӭ�$�'�'��� �=����s�_7�ݍByVW+�J$��<�EL�yw"��wA���e����Kj��|��et�������Ł�7��<X	 �^�w3�����0Ě2j��:����-��+����f엫�ɽ5��g.`���1 ������$F�-9�[���v��{:�k-��˃�@���d�6�#��C���d� ;�����;���l��mc"�'9n2�;��u�uI�3��ɢI&���d�I�����H'P�2��LJ�on,y�+�=������w�+�ҧ���'sy�O)p�����Z7W`��gz{��*x<�̗_��M��ϭ�}���;�<@�W"�:I��\$�O��l��<N�A<��kY���<��*�6�+cp
�C4n��sKɢ T�Z$$�;�?Z+��~��y��K	�@�?$� ��x�Ļ˔��[���j�q@�h���{\�"+/#,0����@���up�,a	D�wލ�$7����7,6�WA����J�O�[�~�����٭6��{��6�v��e6 I3z7L�	���#_�5��am�A�(��3����f ��{���ǲ�`����>#]�f�d�8eA󶱎f�s"<" ������cF�Z{�ͥ` 󼹀��NpŁ�)v�O?gk��ْ�����V�:ϭ�w��z8a�ühk4��k�c�scL�2u�$t�,X:V�!mE�	�7�X�:���3�G)����bM����^�<۵b�i�%�~5�'�����e����=���M�Q�n��F����M�`<ObN��Nn���j9��c�;v�Z�5ۘ�+y�nءe籵���V��j�kcr���j7c�p\rcrC ��������:��zYr�gF�v�[5+a���TM�-`�tu�9������� �#C����	��K�=�ՙ�v��+志�y��
F�/��ֿ� �>�ܸ� �y�3���/o��[����s���;˘���բ��0����at��^&�����l�% �wܹ���Np�x��2-�CFܯk�IL���)��aÆ����:$�1�il�MQ'�.��z�z/{��@'}�.7��y�O9�QO���~�yp;}�2�}��o���, �^p� }�����,ѡQ'�9��l��`اTs	����⃢MQ3�f��4^Md���7�&�����it�$�މ�'!ܩ����os�Ek���7J��lg�A�c��7ۗ+vz&��u8�JAB���:O64�Z������$�w�P�I�w�l����M�	�E/{$�I1��tˮ��BJF�/�M�^�M�1���%��l�s�����v�|)gl��,R�"����i��j:�]x=L���3E@:���pҩ+���	��~�8��v��$�~7���������{q��{N)kV9-(i�f��?w�N�4I]�������t�.��r{�,��﷙���ͭR�R�ǈ;�n�y���l1�[��dO��@2M��j��x�֦M�@���3�H�ӭ��Q]V�|���'�F�v:g��:֬���73x�D�$wz$�M��n��eV������EY*,m�Ղc��ʭphٻXM�ףY;���E$n[�o���|�n�g������4f��� T{ܤaK\g�0o��i����7vT1�����h�^�8G��.m�S$�;މ0����r\R_y��o=�`b��E	)��Lς�]��ρ������s:J��M��z�sd�O7y7igr�����$uvݶ8R���U�V�y��|]��8nMMT�WQ���ޝe��{�Oē�Ѡ }���5��#���-��f�q�8r�|� ���0 ���` ����޶k�����F߾ ��s��6��QX�H`��d�&;�(
>��;���$�����?h���l�[��ޮR�������ʹ�w+��N�5f5�����cm�18�u�,-f��E~���o\�i�A��t�$;�(F�q�+�%���s�߻ۘ�G3����fwL�'��2`�����h�����?<�(O�1��//W\��X�c�T�t�@W1�q` |ﴠ�.�vJ��{ݰ :���`��^p������)��M7=y�D�w����r�w  }��� ���5$`�M7sf��+&L؇��L��[�B�=z�"��ӽiL�U.nl�ĄA�w�m��o-�|��'��C�#ڋ�m���s]��9%Q�Kc@x�V��&���7��R���$�E'1�MO��m� �'������{=������a��*hjگ�mIJ�����F�e�*�1��C�p;J�jH)%��=�c���os�,��;ɘ >߽�����ţ���/�s  ���b��R(���s�5�=��6h�ʮ��;����2I4O�ݴ�H��2	4�(������~=��	�����1"�������`
���Qb��ѯ[�|��s��������I�?eN7ITq����t�=���U}�0�dŀ�6o>m�I&o��g�Aܵ���=��1v�!~��-�0 {��¶��:>�]���#���D��|� ����1����G���Z��51��B|e }�N[ �;��0J�se�Z��S,T��U�X�)��Tۺ����n.��.�+�s��J�5*6�ճru+�Q,�s&�ct`�`�ƙvcBj�V[;G�ɭy�7�l�2;�ճ����&z���[o��Й����>��]6�x�p=*�;��r$�>�	^;����[[�v䕊خ�΍���U��])Y�5o\��=p�+.��寴V�(v�Zn4��yH��s����XՖG3{2�C�+�4�Gos�Q��t�ץ�~rN�u��r���u(�����kf�WW��*$��Ԗv��}:�S���b��.@�s\�K�%��P<{)�Vu�6͐��<�=� �]��uf�cJ���(>z�q.}󗛶�X�,�lc�ǽ2��u�.���x��r�9GRvg3n=����nGq�C}��	|���7{�ʋR2���ת��s����G�U������XYyp�]p� pGWQ��Y]�02�Q�Ѵ�j�ؖ�����p�g Z.�dՙ��p���6~_vcǄ�[/�NX���8�>���nS�w�EI�oKx|p���[q���oq��I:�z��e�C��d��[��e�@/�v]s�Ԧ��x��l�h��U,U�d:��R�]��&�'`Wj�3xt��u������;�t����w��\r�9�v�F�V���7i5,�	�8p�JE��9z2���@��4F��w'aχ��\8O.����^���Nxvc��!\ݮ��wq��������G����Ww���=۔[H�q^U�^nk��#E�mٽ�Q�+�Iy�z�r�;�޽�����b�,�Msg9�^W�F{�9o7JM\���q�]9��\�CsWwN�p�=�������yq6�A��\�v���6#yW��j�;;���$W�4I������Z�v��]۫�����{��yp�ך�ݸlh5�n�j������sW6��<�u�F�;���[׸�\w\�����J�s���o.nW��p�>��~L9����Ư��C7���^m�˱�]�Vܞ|���x�3{V��s����6:^� k�K\���L�:��1��v��sp=���&�V[:�v����C�n2�m����kj��-��k�f�1���ج���6�r�� �ع�j���d��6�y�b8z9�v�c�͓Cv���ٽu���pv����a�t�<[hL�Ӻq��g;�v��nѶ9 ���.v��u�-��뱋�T���;��1��l[K���gu��;u�y\�v{�{u%țɦŷaI��ƭq�:Aa�-�t�c:�X�\s�i��1��3Xt��S�&n�4e�v�9�����s�\k�y�u�n���8�>5˵8��s��ɽ�88֮&�u5�X��\��6ݮ��=q�u����n�7��;]`�v��5;�Qn����rKG-���g�(+wN�Y�!�8uvv��:=<[���nɒ�a��{a.9�a{��6��v� ��[�a�;��9�*:�[���=��݃���S�;��b��lscn�;� �k̦�(CN7cn�םXQ'�ƶ�#�ŝ�	����6F�R��m���9Q���y�]��8�8 �ɫm��3�;Z{{f�����Bk�L�żf�������t=�0���<����ۜ�!ʘ�,[���a�q�`��n/nL\��8+�0[׶�n$��m�"�)�&#�P9�u�Ln07�Q����-{qRݤ�]��*��'��/N������N��n��<�
���A���
:��b��6��砬��kv�4���Y�qn��9�ӥ�F��]�T+�b4�1�]p�p��7���qq�<t��E���m�'��n]7�ژ�����X�n�)Q��e�a=w�^0b�� ܷ�d|.��:{m�{A�ٴ��; \ݯ n�s������>]<۝��eF��^��]ҏv۰�\��J�7B�l�zN�ɥ]��	m�wgd�u�ՅJ���Ͳ|���d�lq0osZ9[�-gKL�x_i����:�lq�)�`�llqv�Z{X+Jv.�	��������ƺ�r@u:T�Fƞ�`^۴8��8�,>|���>p�{�9�J2-Ɲ����������;%�{��e� {���?�����o�%�	����^���+��ďk��a����v:I6�=���|�v���,@ $���&�}؟ğ�l	��6$r]�/r��3�2$Ib$�z�]V�ۯ|��@����X �|���(�=�	D����h��cd��x��jZ4�o�o44���[��0 ��n` �w���}���]�� ���f�C�j"uʠ+����&� y��QN��>�v3@��<������l�=��Ł�Yʯfq��mݓ��(9u�\Gb��;�%��ݬ્��k'&B�^���,�B�8ܝ߾� H{������\ϐq��*�G}��K ���n���лX/	��!�=�b ;|]�#r�<�4�,�"�,��zgyt��{hb���[�37��'E��/�
��^�a�b�n=�gM��-���導x�D��N}*��<��R6��r�r7$��t��ko�Y�}&tH߭-�N״��P�t��|�����., P5������O��@?�v0'��w�0/5b�>�2�J��wٝ��ׅ�٬����{��������G�-|B�M�x�$+�SVV�i�;˦�C|�b�=�A��k��7Q}��� g9s o��Ň��U�>���c �$* �UM�RE�v9-���l���ݧT#�v�(GP���w�#�����PW�Aw���H ~���  -�=����I�{X�o�h��+���4�g\��(I~����f7�y{�'}w�$Eon6I$���l�>}�zx��j��'v����Y,���f\X��d�}�s�}�y���q��k.p/]�����3s+�9�ǰ��)[.���ri�qƕ���qn�ݷ�Zx�����1��$^�y���BL�۫.6��~�}�߻�|�#����f�vc��g	���t��]�{1���y�_z.nOS��W���OIOF��'>��o��� �'M�8����`=���$�G�|��5Fv�$�ս��9ݎY���ϧ�$��ؐ�h筻ts�1W�ޝ2zvk�3�YSVV�k���ϰ>����I�ؙ,�}%�~cS'sۈH{��ŀ�jz=T�%T���ŁD��rg���/��L��$�~��m�I$���`?���c:�c s�*��$VE	/�X��{Z�>����$��T��f����}D�~=���7�z� ���sV�V<H9���'���gR��{٘ �=�z� @��Nbg�ˡ"�I�v��-�h��k��$��9�区���Y~�w<�����a�JbݒRv.;[F橝��zo3��$�Q��*�����׶g7�2�Lx��� ��\�as!8�f�]��0;�z� �g9s�/�^���U��IWQ!$���� c^��#�͸^���K�+��#��=��~���{33>w��� ��\�Ww��z�.`M�3�s�M��q��p�
��ς�����f�ע��>蹗��D�;��2Oā绍�.W������9��U��VQ�
cs������w�0 �|���^�3=�lF��\Ā�������\���K��}�7��|�$߷�u�=�߲�@ s=˘�@#������<��5�[�m���`
so��XAتy�>��I�{ގ�X�a{|;'׽��I5D����~;ލ��Bfn��ީ(od<����p��ڹܜF۝�9��{��ԫbti�zꨍ�1���Yf�f�s�ݡ��z���7de�O��|�F9�����E|T�{�ƻm�c;���I�`���.pG>Δl�uocvn2g��p��q�On'bW� ڜO�&��^08s�^R�0+�bQ6%�[9��/���\]�N�$���\v�%����Z����e�9���F�G�cF��6.c�֝��Ų`Xճ��nzc��k�W$�\��8H�&�w#u��\�ݴv�.&��wa��׭ΰ�t�+�d�:�%Ϸ�/@n@(��K��� @������{��σk�o�*�b��[ju�ğ��ۈ:̘.�����ˁ�{1f;�ޭ���.���ru`a��.`�{��Kߤ~�F{霻�jz�Z�w��縡j+�������b��Ř 8�<sU��<|���wg�I'��:d$���t�WH���F򰚴�,��^}5�ۈ�wt�� ����0�F��\��{^���e���z��9%��rw�K0 {�]9ؠ��^c�n�&��� M�H ��l�^%.,���Xq�7c�#��0�*���n���N v��@RK���~��uCo�{���	$��g�OĚ�;}��&B\��A���m�G}��`%շ�-Q
@(�7D�?cd�)z߬�h�"ĩǓ�U�/�}����ˎ����履�g�����8Bbf�ʳ�ss�+Ω�U�'R*" ��u-8@�����0SܤI�{��f|�?\�����0���f�������G��Q]\H;��kI��A�'�oi�|<�Ļ��@�0m��=s>�縥�:�mC0%�m����u����9���6|{��o�MQ$������Xr_0 O�u2d��']��UAL���]<�o^�.,8��sT�'<�` �3w��d�����B{�e;5ay�xC2$H�d�EQ�@c�]�;k����.�)=r3���Μf�?�����=�rK�� ��ֱ �箞a�s�1 ��*w���Ȗ�y�h�Gޝ��&on�v�)Pǈ9�eŀ�������{��5�� �'�ޝ��&�?����h����u�		�x�S'�Ƕ�5n+��;s� ��]<@|	���t+ό����,K֫�c{%v�7�.d�jW:�
7w3b;���m[�9cU̍f�V��۪pt%
o5T�=��(�m���� �+߄A!���q����]<����A�Q[�z�7��M�w>%�]wH�b"<Wn�d�$���{޾Ƒ-�Q$��g�#���)eN�[P����ŀ;�U��	�j�'�x�I$�{q��$�>�F���#KiA��o���<�GR�xz�%����j��,ayMp�s�:��ND����:�j��
i���倀���L��$��^���XlE���\�> 5�r��מ�Ʃ�rK��A~\�$��rv�b�w�L�$�J��n�$��{�t�$���]>��M{.m����
R:���=uy���>�G�`k���[�/Ky��?~%on O�ѶMu!9lXt-�Og�.��A��)��$�3��&��I��n�4H��Ŵ��>���faJ4+�C��Y�Ф�@�˭;������{���d��Y�R!Ђ���/��mȈ�X\d��=�~�'�Ζ�s�q9���ˈ?k�gق �t�TΓ�y^�3�����$��g� w���Hbǭ�y�d:K�lN��;���,:�\Rb��:'��`�6���vk����Z�%�|�Vސo��Y���}ޘ���͖��ݼ�� s|�ŀ�3B"��R�L���.`1��{�pIׁ�'�O�ͶI$��L��kM�h9wsڜZ���Z�7]3^�����$���H�$��"徟Eϵ�C\���{���`�}���d0�`��c*��w�����ǳZ�w٭` ���� H׹U[媣մ�M�����'#X�.������� �k�s�Ćv���$���}�� /�5�{}yù����um�����Q�y �$��2��`�nn��y�,��2��zY�E�Ni��ڔe�Y�>�����q��X�+�I�q�c�*�k5n1�+gn��W�`M��䢈��\q�H�{\��=�-FyP����ava��N:�L�L���OY����u��.�GFV��Ku��p+�]�e���+!AO��C	u�Wu��q��.�l��L{q�����◌�����<����3��4�����$][��w6��L�%sv���3X
��Wn���m�f;\vx*�s�<ID��������䲊����0@|���d��4�7��;F �1;n�pc�s�������I%�`K�^�����9�aj�M�$�zb N{o	&�jV\Q�����q'�ꈨ�F9���^`؁�vih A���5�9y��� �s  /�+�u�6)b)Q%�� �����/�~� |�� �[hD�{Z�U�{�����r�7|a��et��i�=�Mh '}�5�h��e.;mZ�mL��l�I&.�H��'��khf/}E"oq���v�,�y�i=�#]�]s��6�u�����\����\ƹ��YaG:��n_,���"I$�{[l�Pb�������{�h���Z98�s��eˁ��t٢}�o���/��+)�Wp�]r���8�42��l���u�ըۻԖ2��Q����O:��ί^���u{R],;��Y"!f��~ {�	���/���������fAos�ʋrܻ��?<��IF���i��u�� �s7ڨh���:�4�Mh`>���X�z�j���1���/�_z���I"ӵH���uD��}�{ث����MvJ
!�G`LV;S��s�\ϳ �=��,��}�Bm��H^w� Ԑ o�{�m�9/�:���{9�r��n��'*i2?��5�����˂��u�-���B�XՍ^oߟ��etR�6����D�w���Ğ����%�޿{o}F�!����"%9AA&^����1�F�A��Od� %��ohkoWR�TH�i2@5��Kl�%�D���+|�������nu9l�Q\����f` p�w1`|����Ox=�z�Bװ�Qw/{��^�Ј�X��/��������q��2���Sr�H���E�k�g\���*>O1���k���y"�s�r��f�{$�ˋ2�b��S�0��d����2�n:�x�P�\�-<�(�)�o&��n��Ad�&��Y����1
o�î$�ڻd�2�T`p��Λ���˞G��ݻ��Y�m���sz�NP����k�m����x';��ެ�:>=�m�� ��t���.�|id��u�	GW���/�&�Ʋr	�:;(��$��
���2�ʂHȫ;am=V�l�,�nU2J�RuE���z☋�p��2�˔�������\��(Զ��ѵ���ê�kΑ� {h����j�&`U�6�rw���3��ZU��nmϮ�+ȭF-";H:�7ϠI"����m����B��3(�llp��}l`d�Y�5�Im棋n��@A�68�^��ja�T2�;�k�nC��P��j�j����|ؽ��h����n����f�A���hx��wNl����2m=�,�X4s�7a�S�k����.��\"�Ď�;M>vU3���(��M�H�⫻��O"̬9`�^(�r]o;@�Z�-�Du�ZJ�93�Kԟgtt��T�$x��̓�2*.γw���Q6�f&��9�ֹ�w�ٙ���/��#gr1�K�jo��꽍��(3	Pccu�o7wn^5��wr ����ݽ��^Q�[��湓�J�4�7��snU�'wy�����r��;�k����r=�ws��؇��Sr�wtn�Ӻ��zw���r�y�GK�Ho.[�u�$����I��!��n�'u�<���6�v��{�y��nsE�&Ě<痛�'��Θ��˚y��.���F(i�7+��1�ˇ%����t�{�wr]ݨ��is\��yo{��nlo9�b�:k��{�����\����l#S�[�F.w.����r��<�+��W7�s���0$p��4� ��j0��	!o;���������oӟ����k��v�IF���z�ݻ�f�\z� 9�t���L;�Ӫ$�&���ξS��ӵ/4�~ߵ���ɚ-j���3<��tI�G�ZDj�&���(�$�g�� �;@q&�'�mU"�6:���������v�q�!#�vIN���G;vu���&*����8@v��蠨Z����|z�,�ϐt�1` G��ZA�\���{��1���F�y� ����$�XdX80��&6��8�	����#k{����I��Kn� �>{j� $�S�{�2wMw�N��vǇ���` �;5�h�J�� �.|��|w��I�rVp�Φ[,TWW�=�e���wz�k }�r�?���K�@'��̷܄ҫ�|uՙ�a����w�>4��m�0M����:�p#n�Kxw�����w�X�d��^/�C�5ی�TPWvK�׽Ƶy	����s���$'m��Ej$�j��-�4�6�s33��x]Y�sA��٬��vkC =�fbX�Xf�k�<�rЍ�m�~��t[�g�C�0v��6��5U#�RF����dj���;�z�� >���� /{����h���ʍ3Z��U�DK��@�X�(*�%�� ��1f {Z9g|�7DKq�$�"=�D�O��������ź�(G7����
���v2�)T��W�}D���H 6֛8N��vFI@��Zb=�fbXx�6��'hLm�{(�d�=�[�=��w^������&��{}��&g{��/~�Y����J������m��+�w^�� @�����0箸q�p���Mh y<ӦA�����ctOW�-
�{=�<���`�Ʒ�
�JvM�]�T�E�v�{�S�O�2Dj����I�;�e%]��anrξ"F:26s����W�w<j"���\;<v�y�7c͚����؇a��,��:�@�t���mg3���N������|�a��<:=GS����%13۷��m�����]�[k��7�$m���ڥ�t>jF��h�`'�]�V��ی]t�p6��6�t�!�4Q�I�sr�Gj;��7�cͻu�:������]�;�j�mu����Y���q��m�c�����s�Շ�]����^�"��J5M~Aof��؃9�ֲ�?h�����A{2���%r�� �H�����4��>�Us0-�n���9N[mb���\D� ����'�ݍ�&��8��;���w�n�+���(*�S%��0@��ۋ���\jhve:��&��H��f}�l;��� 4oo�$+uʤǁ��oOrc]n��� l�m�$�~3��l�D�|���[�M�"{u:fA[u�M�z���@ {�Mh޸C�go�y�]~����$�>��n�� �2ih3o|ֻ����#��PB��Ƚ��@f��f��٢`��H�5H)%�;��N�mTW����ـ �����/�s&���{;�_��=-�#m�3{��F�`�ВQ�k�SK@�����{��kwSDT�. r���fH�����b�>��g{U�24���G�:�U�'i(-U7�.�r>�� �t��Ɉ����1 ���+z_{�u��{��Mr�mL##�}U4$ɛ&'v��z ���ց V����X���b o���� �2k@�n-�
������3��JM�?Oo��� >w�K@�TI�$w<�{��m{H xĻ�A���Pǁ�٭ ;�oZ׽�o�9��6�{w\ �M}���o4�m���ӱ������A��P������ۃ�z��e�rM���:�%�?>���������[���9�DI~�m�N�p�g9����I���s ���h����m�����'��l��Ǫ�H���l�M7v�I��z6�?��/��n�^�M��-��c���T��J�o=��X�Ě'9���,�Y�Ϸfw{��4��8�Qq:Mw;q�ua���1��6�g�M��]�1�8��L��Y�YY���j��B �y]�����wx��$%��h2�.�o��ʱbۢ{c������:h�j�ȒOĞލ�${�j����]��s=+�-�~�U�S%�����0H ��vg�zw��" �v�_N����A�L��[d��� 6$i7��kն ��
�*��	\��㣉v^K��lq)o�'%�}�<5%�¨q��f��"I=���f��I��u�D�O��.n���ֆ �w��{|{ZuX���1�wޖ�}��_p�e�Q ��� ���3�o�������:�}��e���o���`��{4�σ53I?m�y��Ā'����?jv{�d����rB�S3�֦���}�G�o���� ;� ��r_Of��1��:4��˽ؒ~3s��x�1������3A�U�իEM��7S�r�s1T�/�]=��Urԅ|����9���<F�1t�[*�9�z�t�I$����#G��X[�x��6�$�ݝź$ '��ȅ����C�~�,�۷ j�'���]
��w�+vH�ц����ӌ������B5e���s�{�b�l�{�}�@#~�֐UL�Q5W6�34{���x�[�������ԕK%P�ς{�Z ���kׯ��#�6��׽��$�D�lֆ|}S������O�رW*��[-�����d�'m���{�ng����߁�zwܙ�o��ց]�(߫v�j��q�ߎ�S��7�?R3�@N�h?��H�׀*�Oǧ���pMZ���I�����޸���!F����r�$�}5��7�n���Vw(���~�$�=6� �OO6�{ZEݰtMoO%P����J�éoY�5uCI4۬G*���348�D�غVj�:���Dvn������ݟ�|��$���ŕ����JZ�$>��Tz-DS�uvv��=�T�n����g���>��6rc]��v�����[\u�x9q��\�o �/]{g�B3�n7����ܝ��)3��w�#N�ͷ-�p�m`K?��|�ϝ�����vv��Еq�]�wWj���q���]�g$ۅ��l�U�7<�	���'F�O�F#\ݭ���vΌܽ�IHۛq��n��H'�z��gzs��xxN�Ų�P�-���_�����o���>d N���@?t�m�<h8�n���.w.7����.�ۄj�P[��D�-t�%/�d��j�k��ӻ��I �� �=�ffH=|��	��{9�Ս��*���>�k�Oā���l�7Z+�o��>$T^WĚ�M���1 ��ٙ���9TE��1�G��^;m�r�C��@+_"h�I�w�`:$�_�m���,�WQq&���ZF����imTSW_{3� 9�L�3�~
�O# _�δ��$�'�@2`t������'�-�9�gjk�$E	����g�=�7g�,�+�nY
���;+cErF����S�� Q�w�-ܯ_ ���b�6/Owm��뫮l�ޞ�|ιH�D�>�y�/g�>�Us1^�b��ktQ�F{u�-���hU
�Up�U��{��n�7r1�	���������D]�9A�{%�����NK�e�ܵn�*�i�Y��,���������,W�H@��g̈������Hz{���K���c�����=�}�&,��eJ[PK��A�k��` x�y1` V�w����y����m� ��m�D�2m�YT��x�{��sKC|��q��/;� >����f  _r>�֏[�+ĀE�fg�
�mi���-�ϯ�[d�I:�#>�o//�o�W��d�e�Kn�$�s�k�^C*�N� }~0��Е��D�3XM�]]r9�ѐQ�yr��XZYg3�Q�*���;[�޵���iޖ�$�D�����i�~�0�������3> ��ד'Ō�T�	{j�$�oW���u�d��$[{��@ ܕ� ����ݓ��~������O��G�,���� ;��hl��]A�Tm�P�ƒ+�5.�	N��+M1["z��6ĝО���F��\S��ddƮ��P��0�)Ir{B��S0���g�QB�14�o�yr����I=��X�RBI%{xə��IVk0��M�ؙ>ż�'v���=��h�l����lH��֒ ����;�`=�6�LD�K����TК��1f�'yZ�D�$�������{O��x�[|��� ����R ��kh/�v��a9��!�>Wj��p�y�l��[u��[��"�T�K�u�Z�,��9=��< �f�� {[`J�<��k'}w��o�$�f��rqF����\�������繧�gS{̘� #[�ր�w�[��h���@^����|�v�\#V9F���i- =�s>� �1�9�u���^�~$6� �H���X����RUs0���{O�˭�zK�?h@�{4� ��u���w�j���,!1<�ơy�B�j�>�P�t_-�=�wh���f0�!�+N��.����f��q*�M����s���I�I$�u��M��ħLfo>��f�M�h��;3�����".�h�.m�I={�m�{���˭�f���+\N�,u -෣����v��Hz]Ռ0��S2�w~?���M�P���'�V�$�w��tH���ۢ{=�=��.�%Dߕ�@���l��
Wf��.�-�z���2~&	V�씊��D��o��f 	zs�3>��P��ݚ�)ɵ�epS. �׳0H ��v�D���4��>P�=>�	4I���f`�9��9=/"F�v��`fu��g���j�x��1V�^��`��ri�@ �r�{���-���HsY����3�d���a��m�$y��L�/K׏!&����D�_��@�m#�c����G���?�r��d�b�3͂t֌����X�i�9���w :��m�U*�3%g���w}(j�q�YK��on��Y�J�N��ф)�Mʊpbu��L{��	�o{*)ՔQy���w-�gi��zbʐj$�� �ª�-�za��d�ۥ	����+�FJ"��N�L͙�� ���c��ZL���h�ݹ�w�C b��S20]nWs�ҋ�x\�+��UM�B�j���B�ٙ���O)��b��a�39.�wrTٴ�uQ��O4�K0���\���G.it�v�'r�n�n���\��S&��/^s*9��V�K�*�j���ldPT�cwgN�4�HJ��;t�E	��ZB�skfoU�kΏ��҃���Y�~�-N�&i���S{�V��f���x;�����or�u� ͌��jU��nP��S�'���_g���C2/ua����j�n�Խxo{ DB�5�.�`������ڷ3/7���Uf�,[ijt��ѩѠ5��M��YYC��m^���q*���W���A��#l^�{ܳ�w���r���i�6�x.��`>�ga�ճ����P�J��9�tfky�׈be�8	�7��]�����#ʕm�8�ip�'TNjo9�N�b;�Y�qvQ�;{���^a��*:���v�̹Cb��v+{�}ʖl�jz��f�=�k�i�&� ��`a�m��W�O5����yzW6��M����o*��5��y��幮U��t����.�o:�=u�{�U��K��E���v��r���b��̽���c\���.�E�����s�ݺy�Z�s�ח+w;F��墽ݮm�o+w�^[�k��Rn���{���ywb��Q�9��^h�����^myk���X�<�k�6�{ڼ<�.oJ���J�%�-��/7��u^���tG�����F��p��sos���^���y�\���ƹQo6��G��y^^.y���<�]��H�B0�&�	F�8gy����-�̚�u"hx�jnۮ.y_Ig����x-���;��z��/]V�<���X�d�Y��tw]�k��8r��!�u���1Ɠ�vwWcC��k�ݲ/̏����p�z�i9�:�Sj��ŷd�^}	�SW\�^�i�D��� �F���ޜ�c��tkK��|��n:R��K�qs��N0f���[+�Q��c�툺���u�9�v���m��nxLu-�Q�xֱ�=�����v1��PT�-t�k2�����֬|l�5ۅg��Q�Ǜ�7���3Ό�8La�o:����N�[�W[���{n���3sv.6Jqɶ��Gf9�]��ש�;tgy�V����Zy�����HvĴ�O�9ujs���^�&�G�v_US�����^=��]�d�rc���x)�6^�n��ƽVvϙ�e���q�8=Dn�q��� �\E��
>ݹ3�˧�I������Ez������:�t0�bu��6M�g���{nh�7)	�i�*���<oA�6#��]������v8���D<6w��N�͹A;]��v�� ��i��v��㍹��b�=�z��1�8�;sį=5��u����|�/�k�,�vpc�Nꎫ[!(v�\�e����\��/]��\��֡�b�xF�x}c�m�o�2<Iq��-3����b�؝]-69ө��Ȥu����-d1���X��ݸ���]c�x��N9��M��ss����ݯh�K�9��Y��m\w�.�񉱶Zɺ�W&��qåv�3�2��gv�͸ݹֹ�\��K��T���+3α��;G�gq��c6�j�q�-u��v�{N�%�����5r]&�o#ej��[j�x��qm���e��K69^l{u�Y�R����9��x�=]8y�D�؇3��m��p�GHJ�q.�9,�b�5�3��{����/|~=�Gb"�ۇ���7lƵ��hnÞn:3`%JN'��wY���_A�LmY�����X�ͷUt����1�^�N��'d�W�����f�[o]zU�xz4��� 6�Br�3v�F�j�q���͓T��e���ua��9K���OǷ8��5q�p��j��<Ur����g��=sv�Pz���H�+G]�wd�����&x��l�t�6Sq݋��!��~�/��啻@�����n�1f�|�I�Ml���}u�ۡ�i�|;ܚ��F����-���~���Ŷ'��=���=�vwSf�4I���MI��T�$�\�;��`W��:��Ǩ�V�,ǈ���ϰ ��k��'�}�R�6Z�+:-$�v��� bA�nW����b���_k���w^���o�0������_ Ǽ�������@�ǻ�I�o���U�HՎ�T��Mh>���f{����޿[tI$�3�� ���$���y�O4�.��Y ��%u��B����c��Ȼm[Sr8���o��q��U����,��İl�䭽 }����zٿK���J����O��v�?{2�J��������f���"��~g��=V����J�J�E�7��x��n˻�����Z�Y
ni����x+��n���G�䩭JY�ʬs�������� �~��Z� ߳��`���ky�ռ�'�:߳���ڥ������hl�;����]{�~��c��{	$���v�6�{�����m�ӂ�XK1�==��{U�y�7�^�� ^�w3:{�������}f.�Mׯ�}V���+�p/u��0H ����SO�����/�5� >s9���w׸f��u��g������9+��Tu2���ɮ#n7>�n�����Xƈ뵑VTԷ�|~]D�U-����^�kC`s��k ���3]'���v��� �/ TI�>��E׋x�`9��űw}�'�MV�D<�s�Oğ�2?6�$�Oz���$�xM�N�{��K@���%���\o���`�A�N�` 9_��CE�7�l����Cs�m��]2�-Y��4�Sa���B�*n��꽥�sB�$AY��٬S�sf��x  ֮{�{���y�{����q��ZKm ���9�r�=�I�.I�I5^��-�I$�]��� %ɲo�|JpR�	f<H﮶b��{�M-��,5U �s���~��0��k��׾s����9���B1uʂ(9Ki���v<���TD��"�"�*�� ��;ިߕU������\�$��['�I$�m�D�'$�1[�Y̚� :�g2�Q&��
�FF���S0-�ր:�����m[˙g^�� �̰Ě'�o @��[v_a7��1=�?�J�2I�M4��j^S�ʪ��h����s�$���Evŵ��Br�W��>�;''���݊P$�-�ާU���DOz*T+���r�p��w��>9����Aw|�3�k�bYۈ�J����Ω�X"��o �R�S�*Ȥ+��=�|��x��|Gz*�f��b���}=�O���jm�Ύ1�/ĂAֺ�'���3u�9s�:��OѠݥ�!�X�,�ળny��ڌnbqg������]d����:AJ�%��9rk��d�Z��M �y��cl�	1jF�$�F��Iw�g��Cf�&9���Y�r4�ص"N�:D<��\rJ���:��$j�l��I���i���x�P�������]����$�  ~M ���M��ƫ�4hɻ��rb/}θg�f`u��^%�j@�O�=�L��E���i��ik��o#��P�z�;8�� �<ԯ	
��v�oR@�o��N�jE�䎛���n�!����CW���ʍe0':͍ޗ.��+����e�:�r��)K2���:�[ǜ�g	��M��{�L����c[�rv��-��)x�9�����qc��z���6Ƹp��<ݰ�ъ��-�9.D!��l��uL����Wm><q�x��� Χn\n6��.���-η��1�2�ՓLY�7��X��v]�WH�
ݩL���!�wc���=>GNǳŖ�cR����k���M�=sh���m&廃X۵=;��8�����
��q�ę��3%Fއ#}~{���U35U3�0�/"	�/��$�F�5(����3��{�HܭH�,�6j������;@|�=��p=�.@�	�M>��#$I�y�݊�X$�F��L�W$I,�D�₺��gbsW,zA�֑$nT�L��&�$TX;T�4O-�f��HvAܫ@"I;T�}ܶ�+H�TC �J�^�5�ύ��a��}���
˲zMm�2�0ORix�:ԠH$�S�G�7��<���`����8�[Q�Qh啻v�(z,ol9�ˠц�����c����}P���_��}�־���y�	�Z��{-K���IA>��RC��*�f�*Mَ�^D��a|�w��;�Y����"�n*���q�9�9<����,�3��N�W=�/�=(h��g�aē�_{��y�DYߔ�|H��b2�X�=�-y�5$���E�٩��I��9�B��(�|:w�H�� 3��x�A�v��lH<+�$UI�t�z6r�����2�x�5�B$�$�&�\���<Sy�������#EV�S<{�A7���1�i���ݔI6֓m/{���O9��T82���7n|�vkS�qY�1�FӺ�GK�%mR��jE��ÑOR�1QFJ�ޔ	�'�Gă����wV�w�����I%�ّ��1&�jW��ĉ�7"j�aq�s�ͻ�H'��$��C���<[;�Uz�����7`�ԉ�) H6���YN���b�|�^z�{�7���#����3F��MA�{w���8��C�~�ǉ5t����y�w.�^���/��{?x�H��	|�"gx�$��:'�oo�t�q��KȒ_vR'��g\�K"dN\�����S���^��"��H�uܠk^��[byVy���M犀�y�	�J>��Vl�Q��r=Y�v��⣎��vq�h�ln,��kp<&LQB�l�r ���I#�:�LGug$]�A-�	��H]��z��R��;y5�mq��g��y���$A�m"I�ι�+*Ť-�v�W04�j���z�sX��'�u�@����vY����^�;H��	U��着f�T��cb��L���$tg\�H$瘦`�w-\"��� �3s&�{B�
�!�1I$с��al�
S�����s�L�����IQ��:vw�=�`���D�M|	�2(I��bz�	 ���)X��k'A"o�"A7rB'ǹ�Jx��4�*�A��b�7B>�$i��mm��@���8���rEM�Ih�MU�9'`׫�UF�3� $��%	�<Hˮ��1[��� ��۔���2`Ъ��jAyY�~[��D�z܅�N��>;y�e�޷��&��?�r��R��=y4�I�v�D��n5�N���\wd�H$�szZ��	�-�v�W��Sh�ۻ�n��+��{�)A#s��Z.����U2p8"��h�L+:�I�{ւٹD)�*��J��JW� ��؂����T)�1��{	z�H����|v�%��9}�fR�T�j�t,L3�5�;���O�ESz�gˤT �y^�+�St��o/�Im^�L[������;_�7Z����k@�ٷ6�l%�����W��;�3/C]G''���w͵P>��l͔� N7v�Χ��\�re8�uy��7R�;v��4r���!�����;���j�E{bʆ����:�Ce�cp��6`2fq�*�MFD��v���n�K=j]�=sճ{���d\�b�d��q]u[�cY�;���t^ݼ���l*���߿���n?b�y%0�|�k����׷쪨���`��L+��Gݏ).ܓ�hQ"j���1��,;�u�a�F�|T&���δ�W,�{g���R��O��P�33�TP�z�"I�v�>$���"U�� �o� �u��.�D#3�^���&�vkb�M
鎭�O4��1�^ ���F��k�S��ukȹ����Øgب{2*@�zZh�N��( O>��'��(���^U�7lJ�b��7m��qoS߶��{��t�����̄��4�I��U4b�0��A}ւ$���QH�@�i	�7ix�U�
32+�P��J�'O4{��8��v&�o�o2>���>*�ʼ=gqѴ|�n9����y��[/w*�$ܪ�ӫ/TX3-��Ε�Dgi������+��> ���Oџd��y�ҲtZf���<|@���^a7@��T���Pڴ��=���"���O<�	9ꡢ&fE
��P����r�����
�ԁ��J��j�V��j"�R���]7��>���/�J��P���m����崑���eܕ�I��
�G{��F�K[M�㴪"DԲ�e�Q��F��҇/=��T����gW:���������6u�@'ǹ� \J�p{�١�r&��NwsM��c~]����13׷_5�ҳ�uܢ��>'��c�D��7�m�I��z������ύ�
��� $�y�+���r&@�Rc4��]NF��M�e��T��F�ߦ1M�ڮ�֎��A�.��.���c��y˫OT<�/�G����
��tUְ���b��*��r�W�
77*6��f�2��]�����.V�߮g^��q1m�T�0�o��K��ZU���t��W�u�\��s�2���W
[��h��5��ņ\�Xq��	��{wlJ�#5�r��"��̊��0r��{Q�^l:��O ʅG	K�7zD���3q�&
b�x���7 ��)ʰ�A:�����sLJP���x�-��V$C��N����'o��f�*rø#7U�8)�uQ(��t�{��H�ؾ2�Y��i�2�U���4�fV�{�hwWc��{W�J�������M�*�t�J�`��;�c�q �t�&�׌[����y�O.��sn�w6]���'��ՓW[�%��΅�Z|����!�L���K�Qu-u��y�9��!q�3�W9�S*��3�)�A�WE�njs&ZEs�{�q������O#��\��x�3,�.)9MΧ\��+�)X:�sk�l��Vs[vٽ���^����Tl�<:�/{�:��̭[F
�ރ�+]/�4	�}j��d�5U�B{y��x�oQ9�j�"�,���r[=·%�rV�Ջ(�6.�,^��f��2��T=�.�j1	�<4��0LL^m�.n[�w��+�ܝs�t.b�{ڏ+�\�����{����׺�ڞ����Lh��Tq�E�ܹN�*9n���׽�����**\��U捝�ݹ�o5y���\�/���\���v�{��n)y˔\��ׯv�h��ƹp��^��͝���9W6���\��{��4��l�;]��&�mz��{����{�G�������\�ۻ���Ѣ9��Ky{ݯ.s��[���w���E\���{�w�7�gs��Koww��-y^��9ȯ9�I���+�<�=ݷ-{�^^�ђ�k����1�v�s�&�w+�W�^zkys]-���8�Z�u��{����;݋���
��<��;������
��|X���n���7��I���f7��<��(·"�v���gZX�_T���0�(��l��B�(T ]rH�{��+֬��e|s{��i���5��M]*�+�j�AQw��tr��g��Spe͵�{v�=��ٯ��}��/�|N;�nu�(
�� P<����Y��g_
��/Y������Ez�=U�v�Vl�A����y�� �u��bg��2v�5�:HK	a�*���T��1���I{֑��M��}Rz۾ �־T ��Y�B�^�cg�Y9�.��y��@ ��  �����,Q/����]�k�t�b�3Ѹ�!hޝ�^e��E��ȵ��1
n'�n����KpC������QYbU����A�M/�ၳg>���L~J���t�=z
`0��$	&� =�A�C�Unu�z��.^�Dn�B6%n�7>���K6�&9���X�T�3�də*b�@N��$��'c�J�S5��:X����o)g�jO�W\z���ަ�)ǭ���D�wy�H$�y(��b#���:�+���2*����#�N�OnO�%:���-]5� '�[iI��Vߗ~-��S1;=�kgw�c�L���I�ݒ��}��l�55Q��'׼֝���Y"�2Qi/�4�Ms�����G���I|��.���'�d�yp���Ŝw��N=].
WJ_QU�G5u;�b�o3��Wà���r�Uҩy��g���l��\�ލks�T]9G\5���wk��|_���DO0�;il�ݭ�+��o\�狆�G���]ɟ[���m��&K[=;��$��nxep=n���3����D;g
b�v��jw;u�)�ok;e�,�v�t��q�u�c�x�|y�m�u�M^�6�H&��ԝ��@�,��VаC�4�n]+=lX
D��Iõ�Wj��/k��rY��8�Q��kvŗ�ݺ���[�u�=Jnu�V��\�B
Iw����H_���>�9�k�6�|��� >��̌�WN���3�@�hpQ��d̊QB��$A�C��*7%N�GĖy�I&��ybz�ov�9g")s ��F���ݐ�-��"	&��!T�Њ�8��H�(�A��H��$LȪ�'ԏU9ԖAr��F�J�om�I��[�U{ٰ�N�$(]�K	l�Fj�"��Ƨu �/y�@�ٚ7W5�j�	#_Z����i&f�u���U�y�-�G/�Zլ�t�b�#�������)^�=�PZ�~>�?f7��p�g%O|I��A|g:
��8�ݹݽ�-T����C��#bb�B�����y*T���5���<O^dz	B��, �<�M�Ҏon38�'e�V��f����m�JPow}�z��p���M���S۹N����_$����� ��i���H3c�F����Uw:�F�L��"��B Ǜk���`[��M�ZhՉ����M�]	��!��
zdhѸ1�<8P�G{�]�iIx�/I��s�*/��d�� Tז�H�DL���b}H�ӤI��r�;p�%���`���"@'c��O7������>���?��*"VΡ��'aE�d��pih�������o�_����qt�������	�Qx�-u�3��3��i��y�M�c�GUd�0tu\��ױKCt��M3B����Z^$��w(x��2�S���ڮ�}��'��}�����IP';_
D�+7yΣ�jZ��w����v�ܕmȐ�+�i��`�k��M,����0��AQ�ɺ�ʉ�?x&����ix�G�ɦ��u�H�)U4��ky���*M�U��I"����f�����B<g=������lM��^d'y4�\粓�j�QTN�Z^$z;�Q$�����������Y�Uq�G������ݮ@�X��t���2a�'9kq��[���͢�,����}���_qݹ@�H��H�VFowN�";� E�w(�eƈB����+��Aq5i����^e����ւm�oE{���۾�7GU��Oݹt�o�� ��hx}l�P P~׋� =��湶zI-i�[F#޷<�t��PjMp$j� 	m�@�{�,P
3�/7��MQշ^nR�)�=/��U����+)i�Fv&�n���`*�����;En?^����� 7��؝"|X�Q�0"E��P�w� ��<Aa����`.��łA����[�A{�RYޟt�����[@Q:�G�Z�����z6�.x���U��<�-��B�||�t���W���HǶ��y�@��۬�v�]wH	��A=T0"j�L���A�5�h)��H7�t�$�����e7��{w��[{8��[(��Ȫ�G�p=�F�.�	=�H��_y%�Ac>�xi{&0��[�C�yH���ă��l14C�H=״���33TA��D]��H Hy�H��7Zj�����"I�ؗ���P��n���YpVxˣ�K��� L�MjƆ�Vꬊ��\�+b���[����H�����a�N n�6�����o���n��Y;Vc�TxͶv��vbNN�v�"�tmVL�n���m�c��ׅĆ��ƣ�d�uh�4xgZj���+��UDns=u���۰(U �v�WklW��aM�`�X�����mـ�l�;v.�F��Z��9�,���Mb�����2	�L	;���qۮzX��v�n+��4�V�u��kgp�:zt��*��=�m�`ykg�ge�3��v�2+�7-ߗ[���T�T�?oZ�Zi���"|Gs�^"�ma�.�z֠��?{��i�c��*�-y�N��&߳�b����}��F�Z@�A�yHn���,��Zw֯&G%��]'�w��I#{r��C9�)�諚р�δ>>�̤�}G��yF�t�=��ә�j&��[AAor��'��.��Id�(��iD�FA�&�Q5}7C ��)�th*�0��>$�(�Lig^�^o43�-RV�cDP�:Bx9�1c�=��^vmi�T�l+�[���$��-m��3r��'s���o^1{ ���V�$���(���"�TP�^�$�i:9�;�v��7�X�w��G��^��G�L��k�Ō��tem5�B���XR5��[��Q ���{Y��e%�{��3��	?���$�}k�M���y̾������Jۖ���'{t�Z��L
���+GAz����5�;j�b,am���n޶�s�=!����H�i	��SA�v�{_{��b-��fe�v��$���))I�ܤO�/:����oK��kw\���,�T(�r7]�íѧ�L���tg���9�MNLȧ"rW���}���yok("A��H�H$vv ���ҳ����@�I�֑1��35&b*�w�;�#�bkx�y��Eu'��u����t� zz%�c��}B��<Ԭ�Y�@���2(EE
��ܒ@���D�a��s�����Ek2h��pxr��:���<�����yݽg���d�͚��gȐh�ܜ�̫4ƍ����q*fsR�?{���� ��֐$�}��D^�N;b�Y󓽠�ފ����t��WiA#u���L�N�4��v���� ԓ"��}H�V � ���@��bi˚D��)I��yH͈���=[��U:�uG���|ՌT����]�Y������d�cV1�}޿�S��Q�;;믛��漉 ���5�o���f[��O�v����>(I���wM�]̈�Mcntՠ|O��KĒ{�R�$廆*&w�V�=�n���K ;[W�^-4H#3r�$����QQ�r�'���-����q�ҡ8�)U6�=���:D	=�t� �qݒ�$b��qB{^���6�[@�sj鄷xޑmH���ؑדzG�7{v�w
�4��E�AMP�b]ꚛ6t�Y�	N&�\������j���3��L�V)�V+;�{��c ��ד��)]+��p:�R �ǒ�m罖a�u^34�����%,��.c��n�{v8�GH�R�4�R��q��{�O�,N+eO���rD�Y���$]!���I�V���Ԉ!�<�HJˎB`UU�w�Sڑ<n�m�&��\m/"H$8��ozח��9b�2CS��'Ҳ:�h3T�6�Q$>ۥ�|b&���_BS5xI t>r�>$�u��32jI�����&R6���CC�T><� �}�v�]z�����f��tA�B�&*(T�D����z¿��Q$^u�	 _sK�к�¶ꣷSFb��P�l7�+R���X{L�N�1	�	���}��jp��ԩ\�\��,�����l�z�T���w�}f����5�E[;u_u���(��[����"3���%��oab*��c�kU��*�(��f"Lm�U0ܔ���,c���@�ځ��lnˈ��ҧ9
�G� �T�� خ�u��J\9�/�#w&��#%�#�3F�xڅ���Q�����#�IW�]�6�t��3{NXi��M���fH��b�;(�;y�S����^�L���a�Z:���؆��a�9}����p֎���Pנ�/�g�;�'�Z�ΠfEw}S#v^M�ѵ�Y0�|���r�8Vh�p�IZ6so]�뛙:�6V�i�k\��o0���v�C�0U�� �U�e�n�iV�@i��x�H%��配����{_a�o2�h�� �[�� M@g&�׍�Bt۹�v=-�:�SR�Q�16�]t��է�b]�6t��]�v
}'R��d��ڔ5�\8p"~y�b�*BP;�f���@N5c2���ɏ�Z�wJ�̰�T�8	����ɤC9�tIM����0�R�y5��,p˫[�͗���s��.�9��V1�Չs�^!�+.Ԧ��%��`eF�f����.ٯN��uZ�B�����OHhpriw�57IS��Ǭ�;]t� k�/w6*}��8��1���i�O��3u|�j��i�m�$���l�4G���*�s���w��^W�U��k�y�����\��h���y�w7u�+͹�snr+�".['wnk��r����\��n&���$��Of��7v�ew�{s/t^F�6��׻��A��{��R`$���9h�DX^�F+t�M�F�t���(�<װ�wE�B�v1�]�{�����U�$����t�E�tQy���������'87]u=tmvy���yt^���\����G^mû���dۅ�ۑ�N�5�ݝ����zyn^r�:�����t1�{�wtk=Ǜܸ��v��˞���u�;������]�s�z�3���n�n\Ѕ^ss���������y�su��ۧ5ӗ�=ׯv���r������r���]ߓ?��$�]������$oJ�6���K�&6�
���n��S��CvOGV�s��Dn��=�'\�b+�mp[b{k��Ҷ؝�E�;v�v:i5�q�tol2]�@:݂��q����#sN��[�u�m���Ĩ[�ڸ�v-�U<��meޡ����m8�:5�%v���=3Y�..���������]y��&��gNW��v�9�`c��<WX�sz���5�3%�pPh�OMt���v�$bq���Ӟ���^��`�t��v��rޛ�>�̯3�ӯnu�g���c*ώ���{kq��C���F�Vm�g\�Ƚ�^ܼd-]��wFh=/MQ�i7�Ǆ�O&"d#�hx' lY�&�o/�2��dNٌ�!�k����nٸ�
k	��;�cr�����nSx���ɑ����h�7:��7<r谛��Ϝ���=��i��{�׬rMu��|/��Sk�j�\:���U��\r�r�ey�vv��e��o�s|�~h.�$�p�.�T�����k̱cn�Hnў��:��+A;��a�ac���>�sW�m_6|c[��^^;]�Q\b;lq�n��p����B&볣��sR�m�4aݖ��u�g�����՘x���i-�p3ζ���Ǜv��r�[[b��ķ[cu[O&b��uvl��6yq���v���8}�Y�d��=f۫&ݟJ�㵝��W�gHv����[z���u�������(Ba�^mج�v�ۮō՝����5��G=u]trb9<u�V�nY�w[�<��-nz���Ξ���7��ac
�{�.��Z<�L���Bݸգs�c�Ѵ��.ڹ�6��cyhp�pɫzm�]����Xqͅ��kmϚ���:�p���/bVN�Û1�&ìa��� ��p�|�|����A�V�w�V�N�;���0�0����gV��e�狇����,�z&ز��N(�G0ֹ�uؘ8�=�$j�J���[Uk=��n�u��z�;mdpd����O0��=s�[r��Ax0�G�K����&�d,���<s��gq�cu�sϤ��f��B���u�vbmm\�l�΂9:*�λ>�v3#\s6,�p���3����7a༂��x8��r
Hݷߗ���ڝ����!7ɤ�M�q��� �sC�Yɢo�����A�h@���*���:g3Ȕ�E��U$g��)�A ���$x��ؐ$��:쮵1<��ZM��O���(L
��n���^D����&�Fȉu<a9�I'���'��#5�pBMfj���]B�l׹��\B��>7۔�y䢘'�v����P"S}�����T�W~3ܐ�0��x.N�՜�MRw��C��.�T|n�b�l���s�-��Ҁٔ=�>��uS��d뛖�۪�g��h��P��|I��"H'c�J1���]�6�g��j@��A&�����(����\w�ԕ]˫��c�^ƽ�yW����r�J+��o/.	.t�z�=�M��QK~zݏu���Rj&\�:y0�
�DI;$���%��i�랽Џ��P��3F���6g0"�ے�H$^n+yf�֍���F�bD��y!%e��&�3(�l�5;Hٴ ���B�>ܔ>���U%�NZ�G�v�L�A�
�(3T4�܌�'Ƿm!��ڬ��x�J|�$���A �u�����`�i@�2W�DM,�������G�e�6^�+cxt�T�&P��_s��I#-m����u�oo}�^ �κ��E�N��Y}�|O�3rW��;�f������'�t����-���mZU��������u�A���Ns{�%��ųR9�S��W��=��H'��Z@��z�g;���bT��8���"m��ځ(�u����N���-7��o�OqGf�K�Fb�]ʸ��N7_d�Ր�y��2qے��gf���UmP�߮����B6�95WYM`$ǹH@�3��$�vTK��;;��L��_P�pWu��F�tv�罔N)�3�u{z�@�H6�א ��ārXM��VBR9��SB*��c�o
�V�n<��	���WKgU�mb�-���7�v7�H��\��$���H�;;)�����j�~�1�_�sHV��|E�D��*��w�������'�4�T� ���֐ ��� H����v�����	"*hT"�$�$�y^��<Ȼ��s��N������S$�P���X�ބ��Lɑ��T9tHD�}�z9��b�`(��ޒ�3''Y����8r��5����E�K�c�8�<xlps�zB�N�R��X7hh�\��&�2��n�����%���V$�ܔx���;|cj�S� ��I��A:9䣇r�8t]�pf�v��g�Z�aI���G;w\��$�g�*��pr5���"�hĜ��#�G�����y(�Q���𮾎~5<���n$Lރi���-Z^=w�|�UY�����m�b^$��y!p���z��-˰�1��"A�$�HF�48srP���d^>YC�l�	�q/F�l�@	�h�dY�'/+
�ں�"mz| 眐� ����P��x:��,�2=ىU���1.*���7fgv�$��h�H�cԛ3P�W$�$���x�O�gZ	�OG�j]���4^Qj���ӹ�HY:p��Ҫ戸Y3�>9�W�|�k�JAʝb�N�[9�W��v�Ԅ»M�(�A���ȟ�ѭ���<Ⱥzق�9��?��v��+�1�S��9wh-綌��#�K���ͣ��;�z��.�n��8]�p�7.#����*v�V\h��֭�Cn�!�us�v�j��(Ӹ���c��`�c��n��Qc����=���]-n|r<������t���uutP��L74aܝvNm�Y�;��s&x}x�F���m-�m�=6�z9����\.�d�+����c���Q&&�����$A ��t���֑��Li"&��9�"Of�D���ЩQl�h�T&î��ެH�c@fs��A�k�O��.��a�:�kNsiU�����e�i�w����~�լ�M I&��D�A��Ldp��jI5DU�;\�:��n�6X�|� B��D�E�ZD^� ض��|9� �Ŋ�vi���y`��Yhw%��Ol�y��A��$�}i	��K�3#�ƻս{5��z9j�QR�"p�;K`��#/>8��F+^E-���Ơ�����A�m�X�z��Nv�m�"�젰߱�R�m���K��������8f	�&&��@��$N;3�]�L��h�(���'����e�Vv4�u��J���r��D�,��gX������̰��B+�NuK����+p$�}t�$�v$O��U8�
�d�w��0�;��ˬ9��o�sݔ�w��2'n����kI��t�݉��V�rկ��r���z[�����'����^ ��訋���/��O,�1"dTj���z�$���BNCD�>ǚ� ���"N�t�b���ug�H�*uD���&ܶmq��뀭�mG�����ErF��x#���b�[�6��|H#��XYb�d车|{1//����iU��[l������m&���Kc���r��y��x���fVˡXf	�&&��^3ՉF��D���5�y��hL�cA�X#`QI��ˈ�]�:!9�t�<2��������5}͜�t\hu[����g.𭶹gv���>$[�A I�n�J�|(EUU���;�K�	�D���/�a�&��UG��ix�7qBA���>���$���yV�(���@'�� ���!]<�rs��4���J��������Ӟ]�O��s�=��v�݇l+�۽�sȉ�Fݭ^���kO�����֑�C%���9!v4�$��u�[��"�aj�_?wZ֗��_���雥�v�$δ�"�j�vt���ݷW�t �Ґj<��4�|߲�;��&��MJ�H܄H;�ii�;Uۂ�ߡ,j�9뻯a����@�`;@P7�� �j�0j
�}{�E5�f%c��iN����:�5��D��ۼ�]<m��.T�!YB�b��ދ6d�~z����r�I��j"*TTIB���w��}xrN3�Q$��֗���B���u�=��TR
D픪I]Q��<�˟0��bPP�����C�uV����a۩���y�D�/���rd�i�{"��A��Aؼ���MQw��"w�N(:��N�2�B���� �� 
�������M&����YX�j*�e�D��j�1�����--��$k�A���������'ʋC��������(IU֑$}��>����g��#{�3�E��U鉊�3��$9�P;8d�)k�}�lF�W��b�GnЫ��Y|��8k�;f�9~��vF�Ћ��l�p���,kɌqXdU��n���j�ʳ�R���A3foX{x�xA��KpB�l�[F���㋷]n��:-�{h���:�q/!d�K`銽u�;t��ӡ�F�ܛcO<���I�5�l1@���=�E�[�%v��G�;�:��Px"C�i=uq�9�\�+��)���=+�,�N�wu:�QlOvz���q�Y���d��dz��(�e�.�X����C[��7���-˓tvIn&�	��Ư'u��N�p؟�]�� P~���@э� �ƻ��	Z�ჯ�֟�Vk�g����W�^\� �R{%�ȗ1�LM�k�'��cr�3�Gf
��v�=���Q�0�3c�6�d�35�����������ݍ�E�����Q�b�E#ڗu�;�͠�>=I��㙮�$���hN)�Btp ���`��B*A0n������δ��lC���5�x��q�^$�w:�	�+`��D0�c2����5�R����ܮ'�+����»1���e�f��|vf(�DLW���}vINk�/�֕�b���A2G�(�f�	:�	�2��L�HP^�"�#:��a|͒7��3B�Do.�?u<e�R�0�\�s�rWo.v��]ɋ�@�;�ڌ�7��:�cs�tMgoj�1� i�$"7:� I#al ���ׄ��*�=1T��R�#��G�������Of��8gd�GgZ��成d��3:�ߣ�ۼ�x�zJ�(`��A}�Kăϵ�����rMX<k�F�����
�4#ܒ�}�V1}������a#c�e H$�m�����k>s'�����m��Y\VW��D�f���y�N'pl�N��K�1I��s���?TX�}���|�$�n������rj��r�A��My42f��O�$ר�n��S��x��h�)�	�k�'��w�ŉ���O��w�U�Z�{�c-����|����ز ���̎���TM������>@�e�Ik53L�ֻ�a�Ȉ{z���3��H'
����!�%�q5{��l|0�.���ЎL�K(�Wua�V6E�b-�y̒��6�_LW�m�r��!1p��U[�����U�G*v�QҾ�����5�t
�ٍRB�@T��!���!�x�Vt*N߰1�'&��#��c�6�3jO��ᓍa��U��/^^�/�����|��t[��c�#C�'(l�Z̺"-�'�VD�|�oY쓝����c����^՜BY��Q�;���L\��-S�qo��8b��c.�o'r�|��2��I[�>ᒏ_3Gc<ne䷃��_e�c���ٷ�L��FN���#��;���o��.u��d{��m�r��/^��ɭt�"�0�T,�94ٙ�b�HWZ��ֳ.���n�]�]AZ}c�����ԕӗ
R�wNںY�ƨ��c�r����77��E����|L'1j�)fv�r���08����+�S��k,�sT\���`��n���e���sӹ3�}>���P�r蠺v����+�@�U-^�fՑ�O�w.'�ɵ{}�fQǙ��3�-�2.�<	�
�|��̍�ȼ
�;uV�a�Y�AL�-9T��ͧe*9��E��X���TP�g,Q.(�dR* ��[]ۆn�˭�5}6��3�Dt��1P�;أ"�Q��5�<l�f�ĘbM������4{�Oc��o/=�v��L*���{�YݮX��b�\��^=q���y�Nmwu�y�m��+����K��.Ou�˗�К/4`�(5��ەr��s��sy^�H"��s����������;�o<����/w7:XK\������'9��+�^*�ƺn1h���v�B1˶�9�\6����h�3n����ݹ��<�5���HkÚJ�r2X���۹uy�uwv���D�h�*(̹�ѣ�Gb��]J
�{�F��l��*+�Т��^s$����ny�&�{��7���S5幋��y]�wwvܢ��:�����8RoCt̓9�k�Fd��{��wU� ��&���'�z����c�e33T�)�ŗ�'�H ���@�}�yݑƶ�b�!�s�� �o_$C���2Mj�����d�5�(F^�=]j𒧱 	$fv�O�+nP+�-㶛��|��V�ꖦ��X28S�v��m�-j�έѻ:·,*jۮ��eb�T�v� E��vA��";+��mto������yݒ��@�&�EH&��r��s��ȣM��[D���Ղ|z�n>���iF�_��˻�[��oY�l��\��5&�H��^H�0|'�ڀ�p��BD�;��n��6nk�/�w�?l��@�؆�A��̣L4�D�F�c=�i��#Eލ�{�<UMD��d{D��@e8R὘-u��
im�҃Q���y�CZ`A��L�Y���1CۿP��H�!�w6�n�>�.��ףA��������cU�p�؇n��ug�e�I�r�r��:u��g��o7���0�]�(�٭^���,��U��i��s7�jƔj4����(����^s��b��&�~�-�I�b��h73�f�V�iF�����+m/3�:��δ~�V�G8�+n�T�b�#/s`��ϛ����I$���?&'��Z���~c�~���4=1H"H�s=�i�lCe�Ȼ��@�Z`F����L���R�[L����bQ�'��g-�Ng�K�8c�P�b=����6�c~��w�]Yh�V���i�F!�&��^X��[�D����X��7�\����/��4�0#!g��dz�:��v�����3��iF�J0�Q������,h����N�ź˻�ib��F�=�k9i[Q��Cgw~�[-�Ǳ�s�U�I�K9h,hǳ�d;��ʫ���6"Ԉ7�g,Cb-���(��iF�o���d����م9���@�=>�b�E�Dh���'��<Ub��Ѧ-#1|��-�m(�h���d�֘�]c8e�5�������I���-�4�"How��n&�80���eF^���}��SM����\Z�ٔ���f3� L�j��e`f�"��Yt������J�ô�J1A��U�I�Z�G��@����Н����+���;7N�8��Y�!�/��I���a��Ӱ͎���XG�	�W��s�0LnLs�����۳Y
�v�|I��ŵ���ã�����<-����m�7��ԯ9��r$�9h*�%��W68u�9�<��^�5���SX���j75��:i��65��cs�z(���̛q�r���W�:�@nW�F�x��Wa��t��������f%Ux�)���-XҍA�A�3��QlV�1F�4F����QlZ`�<��]�HNV�ʖ�z���>���J5dg9~�2�_5�}���^�8��f��[؇�9�x���ΐI��i�A��/��l�6��o��Q���T[�7^��1W��4lh�o;�^)�%b�h��#=������Q�m߻̚�21��1+�ѿa�X�SA��A�����pCq��߻̢٤���;덑�P�q�f��b���U�뙣�1����Nu-��f�w@e�m4F�w��-b��1A�iF{��M,��W��缾�Q�cQ�^�Ьe�����:�2L:W���1]�2zb$�$�=3�杍z�5�=<��6�,�2gZ��6�(�����-��(�1F4{��LCh��jV����:���a�3�Ex[�F��=�y��ٴY1��%�R=�}~~�s���*������3��y���Q��G���&�������dh=3ݪ#�� U��3x�K���� 9pCq��߻̢٦dַǈ�K�IUVe���˼�V�Q�Ҍ5��=<b�_6UE5e}��%N��N���4qd>뙩wk7@�3Sh�_f�eԄj抛�LMџ��ж��=�|�w����Q��-w��LCbA�]�i�m.5�9�Q^;jh�Lw�.���M�pt�6ꙛh4�Gk��QlCbA����AMdC3�硯��b�����2͌�iF����~�4�Ca(�4{γLCh|�cЦ�	�4
�Dy��+�9E�S����J55��yE�4�������3������BC�ר��T�X���~��6!�����4�0#!gy�(�(u���4��f���6�9�z�b������i��y�p譣��+���F���F!��;�gY���F����o^�[-���ܭ�ӭ��ǣ�qH��c���7~-��i��9�ٵ����f��������lh#�{O�&?��w솇�!�D��f���l�2{z�@�X��{����=��w�6�f��o(�1Fb�#Gq��i��@�Fk|p�B�,�>[k��w�Ii�m&s�����
�4o����֘���#A;�^��h#�D����,Cv4��1��@���2j��`�L����zW3�ki��(�1F{���+a�Dh����<ޛ�ޝ3���S3�j>Q��sz朆��o�=79/+Ԗ^s�1�$����	⋷U�!�M}��"n�>�Z���"؆����r��i[Q��23�רV2�	|ᾎ�uL�4N4z��d1�������L��Cb4�A���i�n����׵�,Cj�Q���ea�7���4g�b��Ѽ{:�4X�!;o���p�	X��2�l#9�����j4�Q���y�[�ǰ_51'�Q�L24�9��1�lE�k��`\�Mq�}��(�4������y�'˘�њM���N�Qu�nR�}������xB��#y{:�f��(�(u�����*�3��ڱ�F(�o]�2��(�#D�=�Z4š�b�1o��9Zi`g���4Ұj4��b=�v�l��c՝��V*��0�^Zh�s|�i=1���wrkx��8�3��i�h#���@e���4�Q��̣L4�F(�c{՛��v���g)>| �Z�'��h�V*��ش�Fb��L-���9�{�E�4�����}5��pt����(�����	s]�.����G���Q�i��17.�%UX���k��5��u7U��iq�l-1F{w�-1[�#Dh��eŦ�0�(�v��᥽�˯L5��6�ҝ��^m$���:z��-'H���\ ��W],��w5�c��3%�x���.�f��}�>���@� ��.��Aj��~n�8:�^�8�U�s!��")6�~�5�;h#�_�7���S3�͠�ٿn��-�lCh�}��é�0�h=;�f�-�4w7�?��jkJ��B4����4e۷e+k���F�p;i=�������#r]~�]g�DH����b;����^j4s��2hkLC`FF��y����h.�L�e�\���!��\�h#����Q�i0#",﬊>J*`�;L�Ҭ{<�5cJ5Q�5�M��uf�l�k4[��h�Dh�}�eŦ�0�(3��5�iX5Pj0|с����a��]�-��;S=x�UVs��Ac��o�=1AD��NƂ8�F@`FK��g}f3U�k�u�L�iF�{��QlCa��0����/4�cDh��\~���V*�F���3�P<�Y�w�<��b�%�w�i�1�F������b!!���N�u��9����!��=�{(��+|$0��2J���^�{y��iF!�����X�l,�w��y�<�B�G#D�oܴi�I�b��4�;�r�M+j4��b;�z�c-��d�tǔ��?~�b�Zt�!F�L�b�Dӡ�oY�N+�uc�� ���)�[$dK;s7v�nH�<A������k`�r��#�EMń���$k`lI�p1�n9�s��S��to`Z�4��'��Wc2�g<�at86�����.� ��V\͞q[�"#��)N{UَH�)ۮ�krl�h��o)��0n�=���8y�#��ݎ�[�;�����J���������i1��S�i5ր|VT:������Ű*��`�p[s���1v5%���6o��U��v�6�c��C���"��y�Ӵ4�l�����؆�O&o1�K-�yE��b�#a�c��i�ƈ��l󗊄�0��QLV�F{�t��Q5W�wXr�=kM�}�Mi�l�oޮ�����^�,�!����vo3���o(�8����Q�QSq�f�U�g���iF�J0�Q�޽E�V�Q�&���ֵ7��yԓ��'��ϑ�!�xaPf��k4Ҷ�J&�23�רV�h!����%UUHL:WM���f������c�{�Rm'���cAh##2滐-�lCjپ���4�f)��ﷱ6!�{��4q�4Ey��N��Ub��i�l��h80��j4�Q�\���I�0)��x��UZ Y|F_e�<	�Zq�l�5��n4���̣Mm���g5�ʗ�����"t���Ӈ���{Q�^�|�nZ��`��9k����v���^��Қ�o9jƔb1F{�����CbF��s(�-#q�n�P�����=��9iX�iA��������[A|ᾷ	THV*��IƊ���LDD�z�u���`�^�t�$�����Ԑ��#��yD�S���j���H	����a	ۀ���UŚ���G�2ɽ��l�M(Ѿ���-��a(���<L�|4�{VѶ��'-�K�	�a�)�E1[����[J5���s��-����F��rk��}\���ƃ��N1$;���Ao��2�3I�}~�
q�+G@�hiWsʶ�ww�nvw88�Z�Ҍ"b�ﹺ-��A�4D�&��rѦ-0�PF���-,f���%l�{o�,C`q��u���
�&�Ī��	�K4�X�G��k(�#R��=�]e�oW��u���m�1��^���ҍ@g���(��hb�"h�9ulCiI���ԪM����EF���P���b0���a�<��;)c9�ߟB���`���_~M(�_}@e�m+j4k�߲hkL���#A�r�,ChK��ي���������a�{\�V1�v�0ǌ73C�{�Uyx��5��0��n���9���b��1��w�F���6��{�����Q��y毺f(�.k�\0���@e��6k��U:�C6�6�c��C��$���Yv���F<	����������(zv�e=��e)��m<��i�#�ru��ߕ�/���]GvћJ����F}"V���f�.�5r����2�r���iF�w��QlCa��0�D�9y�E�F�M�]�*b��S�#=���{ݿ{����c���5Q��[�y�[I��m�9y�An48�6w~�;�������Â�q�}�o(�40#"�>�r��q�`i�M)^�3����J0�g7��c���pP��Dh�Ϲ�F���1D�4�&���ZV�i@j0##=�n��A���7�u������]����IÄA��,��V0��`�HC�uusr8_���ʖ�A߿V�M�����<����6�����lCe�#'��G�>���������}^#�}��41F1F�w����#E�~q�`�UUV!�[�3��pam(��.o�;��c8��F��w(�����s���Ac�Cb!!�{tX��.�-9����K��@GԴ�L��%Ud�iN緜�m(�Q�LQ��7@e��F!�s5O>�y߽�g��#�Cb�Ҍ��/9bJڌCg��Э��_8o��ꇇX�f�'*�������]��ȏG�> �z�`�G�1������mX3}�����Js�LP�S7��PV�omL$_���[������9�ф��L�.kh���[ܟ���$U�ԓl���U�W�U~�_�>�3��#D�����&&
�7h�+L#9������(�h�����;�}���&�0"dh L]�報Ƃ1��7@YpCph#�7�s�Kmo�����������'���]%gq�=��/�{���u��c�1�b�7-�����b*��}��JV���mXҌ"b����-��@b�Ch����Ѧ-0�U��k�$�Í-�y�rҶ�JFdf���h,+���*��&+���h篚�i鈒~�1�/Z� s�r�6!�C2-s���`F�ҍ�7��hb�C`���4�g�y�G���}u�P����BѦ-0������Q�҈j4k�߲�`i20##A�>{�����߽��{-�h �$7��!���0߹�ef����c�T$����m)����W�<W7��X�lCaLQ���E�[� �&���Ѧ-0�Q�iFOsZGާ�)�*Lg���}A6�z�m�ooĕ%ìT/LCh�;�d8��BA��y���Ak]|Ǽ�m��9w�l���DҍF{��r�0�b� �A�{��r�cDh����Q����M�Ȼ9u�j.��ƃ���՛f;���tE�f�1�e�=yc�E�Ѕ�u���%g
�tU�8�$� wҋ��˻�ޝ5�!�,t��\��u�;k0���W�{�`]\�"�����Y��;�;�[�8u��uq����}-\ �1N����b���d�|_rEw^�+��S̽���c�cM婖e�Rأx	+���*p���s�o!�u��Յ�!�3��'j�P4�9���&:n���BV�x�B�v�f����\4���롙Yζ�����AOL=6ec��U�2����yB�t׷�e^Z���AU��"m5K�-���6�ü	7XF���U����:���F�;�J��g=�V���]L��E����ΣQ��*�,kop=M �%�ٙ�R�XF�p���R88������y�y�ܰ�xqU�-�;0�J�]@����ąۂ�D����%tl����յ���:jۂ���vkU�&����e#P���B;}�w��1b<�U�k39e7���&* ���L�+7�D�ƥپ�F�U���G25:�{5��]��00�(+����)OT��x�c��Ĺ��Mn�C�v�*�fSt앙1w]�/*I�ӵ\ؙ�i���Kt���Џׄp�'�1r�wڪ!t�j �WO�etj9�aI�%�/�bY�A��B����P=���^1���:�7w\��J�����s�ۣ���WwQnw�Ey��\���wwk�<��r���v��C��fD˸thǗIB�ǻs,i���/uyW�����"#�2E�7OwE&Rb,�A��"���y��	b5]9�u�"��^������I4�w�Ή��B�(ɯ.E��E�w�r�w�v�۠)��^t�.s��Np��$��4<�B"�nk���ģws����^p���둌�s(Wwr�w����Y���C�8Q�`��fQ�\GͿ�4��7���l��-j�I���˭�-�����.�6IH�V�wa�3ۮ�x�y^;�^�]��U"���g���;O��ny�e�l�Rpm��%l9��{s���X��r��\J�g�}�=��Mƺ��>)�B��'=�e��qr��{������/�v|ۍ�m�c-˞���o6�M�ۧ=8�A�)����ݳ۶��c�Wpu��e��Gf�x���v{lg�֤�n�9oT=s�M��ɺe�Y4�K�$�F;G��[�{3���N���؝��õ̓v븋��8ԝe�"z��!`�xk�N�+�s�DbTs�:��*z������h��C��ټ%{�k�N���\r�Î�+�qi�by�a��/�M��@��&����dqO��q���z��.�1���<�����q�nH�keP���zN���'��]�g�4*���d�'&�N����bb�,�Vyk����x�9���4:;v�c�pO��c�ƹ���<�]u�j����kY��u:�U�9���K�������j7K�������]�ɘJx�b��������5��C�����mr4wA�t��`���Zwj��۞
�fu��wa�Ի��g��<��c[{k�1���e���j뚅b�8���y��	�����O6ٶΏkk�5�����Z�;O�1n%룂��ƻjضHMB��K��\�P����#�c�ԅ�OgT�n.���V^ܧR,�[e:w�;.�N��\Jn��ȝH�m�K[s�.�E��k�3
	`��W"n���:�օ���3��h�=W,Omy:�mV+�t����!��1�{QȩX�s`�v���U�)yn^��7ecz}�V4Ev�R�t�l�ص˶.zkV��8��띣mѴ��X��ƚ���q�SmQ$(�s�ġ+�����kq<�pi$O;���gv���ƽ�x�z㷞6t׫��v���'k��<�v�܀b��8�8�N�p��s�9]���x���۵��l�7f�g9��ss�;nb��:M��t�����R����۟f��q��=�<[Gj�z�����V�Xh�g��]�+�{ik�Đ&z���5�C�Vs��-یBsNoF@J�(��N�y�?���Eeo��Ce�@e��j4�Q�����CZb @"���u�>� ����:����"HV�t��CA5�o�E�I�/��0s�1U#���@�U��(�6���oesX��ʯ]b��4A�4w�߲�b�Ҍ��7����ҍF��k[�I�d�{B��h%a��T�UT��R�h-Əz�������BD���mq���ɏ�X�rW�f���m���g{��(�Q�l �&���-�#DY�z�;
+-��ϖ��m!���R�����bK-F������6dh���-�Ƃ1C��(�v�����h#���Q�i�]�cǊ��U`6Xҕ��rմ�Q�F(�o���+a�ngz��pQ�m[��F��0�PaQ�~�󖕦���s�+e�<�Tf�!'����<)�m�n�m�lu��u�un����]v�t�nT��w���+ь:��z�yƌ�=̆����BD���mb"`FC��2��5��y��sFd�V�x���[1Fb�"h��7��[Dh�oM>�t񉂪��S�������F���z������������N[�rnim�ryf/%X�_�0\��v�P��yS��|�B���Tj�N9[��Z���jz�����T��G�ܼ�Mi�dh���,Ch,q�l����n=�|�����5fb��8� �����
ê�q�f�Jz���Q�Ҍ#g=�QlV�6!�k^����⯪vz�>GX��1A�h��g,Cb����+m�>�ʕU�Du)]1����!��^���X��jD7�g.Ƃ8�F!�[�(��j4�Q��̣L�}��j�6&�ca�}��h��m��%B�UN�̢؆ɟv�����Q��F��s&��07�np�n�m�����{�o-���6{��e���Gw��Q���CW?!x7�_�{H��*���4G&tj�nս�ۇ�����6"�+�;��������T�� ���s���Q�l#g;��acbD9�w��1ha���^c5����Z��`�iA��������[A/|��<a�u�UP�4h�{��hzb$�%�ԙ�����zgY�;h#���Cd׵́l���Dҍ�̢�hb�#a�Wk��ww8�w���GF���m>[t񉂪��)���3��������iF�G}��&����#��g�7�Z���oO������@g��]��Zi���w�?����+nb���)���}����XP&�ѼٸJ꽳H�jL�u�q�l�5�,Cv�G{��P�<	��HsԚ�� ,�>���U5�]��۪���Kma4���5���lCh�DhﹿeŦ�0�(3X�4���ou��j4�5���~�X�h$��YR��P�Vt�[��y������$A��^i�A���x߲B��f��}���iF����Ql4Q�LQ�M�=y��h��ٯ�}�i���ʻJH9�7KL��<�s��.�ZN0�9l��֨�Ӗ�{���(����˭|�&y�0�!��Q�|���Mi�l�Nz�M��f�ٌ�߮oLG$3��j���h#�s��Q�i0#9W�I�&7*� 6X��3��5cJ5Q�;���f��y{3����Q�4F��w}�i�lZF�k��V�iD�`x��g��[�J�����e���t�GXuU�A�ƌ׷솞��H" ��/4�h#�d�;������ �t`F�ҍA��7�L4���jsךbC�_�"həR
�<	u* �}���&<=oS��Ҷ�En�ܢ�d`FF�ǻwM��D������{����q�룵�K.s��2S�p��#�ێR��Us`Ck�Y�(�ɨ�����IN��neNl�z��|<	���0�w�ef��ϟ�`�#u��c��44���3LCj�Q��9�j������r�5���E��h�5�vѦ-0�CiD�c���JڌC`A��ߵ@e��z���sϽ�ω�)@"4k��s<v�ʻ���du�h�tr��UE#n�s�*V)��?SA�5]���� �H�SݼӶ�1����TYl׽o��gU����Y�o��4�@�F(�ǹy�!�^o{�+�X�*R�i�l���q���j4�h��p�9��,4gٿd�֘d`FF�S���An1��ߵ@]���G��ᚶq�;�{9Fٰ`FC�������U`6[K���i�mXҌ#g��Qi��F(�6��r�>Y��c]G��1F���4Ҷ�J&�23��P�2��7���u�UPͱ��Z�C�{�돼�d��5��b.A�e߳LCv�����/�Yc5Q��{��Q���U�S̙�8-���D��w��1�����*�V�S���4am(5Q5;�o�E�(��1��]h�̍G�\�ᠷ8�6sw������{��|0� !]�iF]|9ܔ����h��Xq��`L�*:qL�V�k�T$��k��]��H��&��X��z�<�j��I����$C��t���G>̇F��v-�;ݴ��.=sa�+�d�'lpl�۰����s�ۋ��zv�Nj��v�?�����\����2��8�9[n�h��n6�n���fw����f�]S�MEqG�V�q����[���Ÿ���]�Ĩ��ö�h�t`z�1�l��R�	��:��]��ӭ�Z���q$��v��sK��y���	~#���~��L� ��$����7�ᯃJ5�a�9�����lCh罾�Ŧ��ў���SE��o�ᥦ�؆�v�B��h!0{vT��l�wM����5���؇;ޱh+��3����d`FNr��-�mZiFs��oI���}�ɮ2w��&��
�U/ٌ���i��ߕ��td��֣�ݰ.�:,�;�Ax�����gH6��s2���7��eh��o�s!@�ONl �yY�#sd4 J%�F��h�c37C=�ʝ(DTp�2H�"|H}��d}-@=�5{��hvH�2R���i�Fʚq]���h��`�i|�n4VHB\ο�:µln.��Z`��z��E��Y͌�Sy ���Y��e��(��R<�8�;g9�?/�U��6eV�9y]��Kw�S��ެ�4/8Վ<��Ӻ�Z���Ǌ��j��8D�~Us�B�e�ל��=���KPc۴F�ݤ�U�Vi՝�K]�����31��Ѧ�@�t�ʈ�Y}�I�k��vKP�>JO�8k/2��̓�~����mu� �{'T O�>�<�]�ft�7��w~.n�hI"��픡 I'�ja���"�<�� ��-B>�My{5�u���=�9�=��Q�{�(E,U���]^�$8\w&�1�Og(�J'u1�
�-�����F�v����H9��#y:G{��t�u�u� �<����u�"`UI2��H.S$��3ienߺ�T#����7��-���qz��[q���� �&�$�M@$��,UЗG��[����n�g�}���H�����Y�j�`7i��k� ���i��{��<b�3@sZ�����Ȉ:���Ir� �&��A��b��@��@�(��s:%��'�9B'��Ŵ�A�m���	����tQ�QFf��z��m�$z�m���I��ި�sYNb�$�ϖ�;��\��3�rs�~`�@��cuң.n9����r����P�0Yʜ���}�F���tUP�^�P���H>��n�=h�3�Ƿ:�����\���I5&��!�7�Y5JZw�3N�ƨ���֯gur���^{}d����r���e�!���-� �_ruf`��|���'�jT+�'ysc8y�,��a{M�!FS�����_/ A<�m�$�)<�R�F��.�1o/^x����oVm��b�Q���x%W���6��E��;�s��������Uj��r���C˼�;����&�����B�J��b���n� zF�ɀ_��>>M/s��`�{!�@�Э1�^��3뵱�w �c�#���w���95�������ӍW�{~��R&EI�g�����9ں��	��f�x.<g�א �frۿ2n��(EU��J�&VQ��&���u~D��F�-�X��/TV%܋���mc��x@�&��T%�w$���|r�(�'�C�|�=$��vm�s�>�i�:������/��ע�`�Ի,X ��uB��w�A����K�yb�iy$�$A�3Mؙ�p%�u�{�m� �l�f�wd����>#yrHz{o �5P(\2/#�6,���J�W�ٽc5dҰ�\�m˺�r�
� ˬt�	b��m��1c�lǝֲ����+r���j��mv�e7@�#۞���f��8�U[�Q�Sɗq+۰�C��\�4z��l�8�%�j�Xƈ��#���=r�wn��#n��ɼ�u���dz��c��^7^�p���f3���D���r�]ku�mbs�x3nM�bݎ;=���W6��H8mB�T�Ok�sk��3�n�G>��*�=u����Li���XQ�ڑ�r닜갬R��x�Uݒ|w#T"A �.���/���G�$��K�4�N�,�fQ��3���i�c����$սJŐI܎P����6����Y	u�'&�D@�MB��!�6�O�b䏉0����O,-b��$��P�	����M�� ��Y����=���Gi ">F� }9jČ��������� H;DkAbԓ(�Z�$���}᫖��yp�'yuNmv������g�4�᰺l]�n�d�F�͹�1p�`"��]�ct\��v��g�|�RL������y��U�tZ9
�|�!O˗�PT��,�4A1!�GU�x����*����=W��F�=p:�����P�.N�N�핖t:@J}��j��s��.
�I�q�El�wTf�E���]�`�\f������6�]����d��&�׮���K��u�&)Y[Y���?�-�gOj�NMF���"�UP^픣7dɬ�s�C�z�	<��$�-�m��>얡��Vn����F�F�H*��fI��L-�25B�NO\� x���O#6�P�Gd���t�ӄ��7�����~�<��΋�^,��2[�e��u�=�D��,*v���M>�5X)cs�3.�����I�K�@�O,�p�5Au�N������`���"�ww�P����Y���|	�d��O��Tf���qy��ѓF�Tģ����'ǲ6��������"�����9�d�Wљ����S���b��4�;'P��OM��ok%:�GpJ�ɱ敎�vf)jl��om�x.��켴4�ϴt`�9u�{4�-\3�f�+��xh�y6�Ndt�.ϟU�Y���ŉ�f���{]!�(AB�;Ed[}k@�Q��k��5�d[�%3L5���{�직>/-�p^�=VR��3�v���rM-V��}�p�0X�]����޷�vi�p9SM���\������m=W�F��p?fB33쭗�(%��V657���[5��n���ՠ4V�+����~��+,e�'Zo�G4ND��8M],G5S�O+rsS6�%N�p�^ۦ2�ō5r:V&�,7H�i�)�@�O����O�QR�!��:�[ŋ�#�ص��.K��Z�v9�v��Vc�9C&�j��+���Č���9��R��ae����"9#��F+��;�qzfl�G��i�j�/%��󶂠�0���8�����.��=�d��VH�֣�[Z��|��۝;ʶhG����
Z�wJ0����ɘr�͗b�Y;IXs�+]�q��b	����N�*!�9j�m�%x�cq�L�>۰���Ҿcv��f��Ӕ�a嗘��p��Q��>z2�2��G��a_v�s�e��d֛ψS��P�+&f֧�.q֩��GL>��KPb@���.Y���aY�&l��]��m��a��k@Ң�3�9SsJn�������R	'��@�||tW��фш��������S0��M*{���DLds��!0$�$N�.�,��2w;u�{��L��0�$������9�㻩Rc�����"9ӻ�7��H�D�9�ܻ���"B�Y��Nq�Ƌ��H�㹄��1H�wr�)a�0����2L$�:H�&Y˄�3΅$Iuك(`���BR�$)��M��w��)�	#Q������� L����2R
����3��		J��F���6i�F݅3  J��)L��� 1$Ќ����jcw[�c;�s�m��cw2�-z&=UBԚ�����wPz�	��DUf+�>9��;�vV�QQ�o��{wi�UN���(�Td�1�̦���{U�}W[X1�k�;'nw� ����F.ݬ�f�X�UDH۶�P�V۷n1eJ�E�t�w��d6Gj�RAI/V�����]�����+�(����1G���i�C�i�����j�R����i����U�9 d�__��I/'n�$��/i�k`����>Zv0d�	�0d����"H�MI�VN��޼�`�	̞�@N�Ԉ(^�4`MELJ/��%�0U-�1� �E� I �i��ͧ�Ų&�T�Sض���af�g9�w{�7�[:Î�4�����u�ql[׷Y�M�mmj�B޲�1��̖�fL�דh�4)w�8}k��A�&��"@-�����osgk���D��B�7�	9�uߎ{��_�yisr��T�$w�b���-��u��Lm�S����Udh���<�z�]l��{�Z4��[H�H�}w�y'7�U��΄%���h����������Y6e�w�e�R�	$��}j�% ���Í���N�?�ձ��OU����1,Li�rq%�S���j�$�s٘��_�'�)Ty�N��3����/y�ȏw݋$vK�L=�A��	�O>�F��ܟT		��^/Rwd=CSI��8\u�r�g�� 	�>t�����IqS���E�K*�E'wYv�Y�|�6�r7Ժ;&!}��:=���ː������qeݝ�Gڸ�6̸���ܩ��	�jN�;���#v0�u����{�X�Z��/3v���wf'�/|��2����`�x��S{;f�L�<q�w��#X�ib��=��^�Y��cg��UcO��ۻR\Z��^1βS��u��P���s�!i�(�Wl�Ҙݷd��n$�˖��Ur��&r�6m� �D��ٷ�/C�M��m������7m�H���ݶ���������X�j
��{��q�Z�Q߻�1��>���ŐGd<�h��$�^�o<�ኡ��hE*�.�J%Q�|�5V�;�"I>m��$Gd���!���.8���z����yd�fvj{��|dnB'��G��wS<��ۺ���/!x��H5�����&C�]3�:l�"���,����yE��vv�fd��ޫ+OB�1hL�*�gv>��*���՛9�T�wd<��D��oW$�̻��7#�f4P�wL<�n8�7jf�\/8wt��t2n�3\F���[c\�T		����]vH��D�|H˒�;����v�زw'��-�&=B���5�`Ծ��R��s�+:ۥ��dܿ����Üz�DM���K*�zdV���Jy4Wf�t8/a˞ˌ6�"F�.�ĭ�rT��`�H����o� �9Yu|�]b�]V�h�F�
�U!{�R�#ښ�$t��e��N��C�n�I�\����<A7�����vz5��_J���B�{H'Z���&�cP$�Nd"|v� ��&�L��$�#kQ6�^���齅�� �o���7��X2F��������M[�ֽ�r���z��v��S���U1�Vkj*�Goq��}q�uH�פ�餟��^o;�����l�+Cff^B�bt��R}P$P&f$C�n����5(�:utF\"'y4�>��w`��T=69�U��
Y��z�R&�Ϯ�S���~�F��k�WH�1��"�5��\���3m�
�ϳ����ʵE�#����N5��K��:�n9��k&G����6��I��w�u
���z� �&�{.���D#BP�����a��W[��o;�񝴑� �o��Ăy�i�TΉ
\9�N`��yt�Õv+$������+�ɞ'bD�obt����J3]y�.)Q���뻲K�G-,n�a�텠�slU=1�	�^0b�.�q�Q�� �$�B�L����@��w/��'��θ
n����ځ'����֞��D�v,'����� =�f�j<}��|	;ݸ�������1���@�I�T�@���3ܚ���5��Ǵ��̸1�e��(��F���M^{���H��>O��* t-�`�ܞX�	8�\/	;Y�{f-�jt�Q]�m�%� �d�Q����7��z�[����fc,����>�=V1m�ݮR�]�[[e��P�m��=D��p`yA{���$�ծ�lʅ��c�. ��H#�9�j�3*�pud��	��Qa����=4D�\e��-ú�FM˹��:�),�G����˼��Ѻ"=�  ��a��r���0廬۰O�(��r�"�� �S&P�U @uڢٺ��H!�n� �g �raGa��+OB&��3&J��݄	$��H�����(�m�|";�B��بg��MH��Ġ��t�����+c2����}z�.�|�j�5�M� ��n��4G�Q�5�va�A|u�e��`�����ٻ�alj����� ~��ѱV��wJ�؇^���9Z8����]Y�%D�Z�=w��K�{�I�w���Y���v���Jt0C��2+�%?�yo��8ݩ��8
Kb�y�s�;*�#��nU�d�/�s��6��ܞ֞�����z'�GE��Ǔ��4hN�ru�笾�&ո�7��q���=�2:-ŗ��8X��;����Ÿ"E�u�:���iǭֻt�4�뙳�b�ӧl�
 Z�8��>;�(���QZ�mQi���۞��KTjyy�v&�V%{��16�6�.6,vz���9�K��*�Yʜ����>�>�ň�H��k!GW4�"��+N��=����I95�O��z�\�F�e��]/��/*ud�՚�Ҏ O��f�	��/^	��U3�ꛢ�6#�$(,f�R&P;<�s�ܱg���~�]���E�	+Z@�|�����3 �Й��g�K�T/DV�3I+V$I�}�d��r�g
��$Nu�66��"h�3����� [,�PY�{$f���D���r�	�-�P;�+�/w�ҽ������ls<�X#��~O|7=�|��v���x����uU~������-xs��r�|�;�V�e�	���u�� թo�[k�g4�+(�^�4��ǝvs����p*ʐ���{f�D�mGgV��׭wy�{����d��kx�uR>�I�YJR�e���fJ���MB��y8�i�E��Ds�b���\"���ռ��M�k^هFYKe%z^���`���8Q�l�[.\a�U�W���c~��Oj�Xu5���lx��eG�*�v�A=r� I �gt��4�;_Swy�����Ŋ	�T��2I��� �Y��5OJ�=��Ƭ��H;Y�)�ctH}F�a�T�hЈ��N�ںےwe���fw�d+6�&�ѣ�#9������&MD������'n5�D�՜�J� �WIs�&�l1�FD����@�s��Y��Қyd��-�՜�>3/_K�v�c��=�D�0h�ˮ�� {;U*�Ɗz���S[zé�p�f5�v�=�u�mdװL�15/���\�w3mt��F�Nkn�k��[o�^�Wx;0Le���!�>���g�r�fe��	�Y�v��f��$��e"����R�o��~
sžI��L�lZO��@�q��+����H9۹~���*�����	�4�����ܻ�sw��*,���1"j�Gvۭ�:[lz�3����5C�6}J�"$n[�|�^PB&L��p8��9/{ۖk}���\�xi��/}��Ňr8�ѫ	�g�]��E���{S9��a ���_v��'x�u��{�M�@���1�$MA�-0�/#�I���d�Le
q�Y�Sj>$��@����OhQ�D�]{N22v3�#v� �R�Ww��^��e\����M�5�u8��<&|ߴ7�.���Ц�k�s�P�m��:�d���������[��gV�{���R)ŝ��w���`lu���
����sT�J��]M�>s���� �������)��A�;L��4H(��z9�6���N��R�)H��XӢj��
�]�^O��`�z�T�78��ۊ� ���P%�R��%nb@���V	M�bhDɃpc�_��X�aR�*�ޢI>�޻�}е�F�C3}n뵝��{�H*��Ӟ�~y�E��L�NT�������Y ���(]�"�ј�k�ʹ�4�Q� �z��/��| �{}GE�9-b9����lxX�F�R(���VJ$����5�ew�)�$Z�H���$"Nֺ�a��������q�� i�ڵ���}ϣm�	!~��(��@����ln��X�?��1�������M�cjA��BH���"��h�ZߢJ��%9��!	!~�q����_�_/�~�Z^G�1�p?��h�~��
a�%��lޚ�׶/�n��'G�2��� !	!r]�����_��}��kmo��|�V������5�v޿�����?D��A��ZX�=�������̇���I>��$�	!o�����?��ldX��00�S0��(g��.�e'���K� ��`$�X��_����O�i��
>�C.}��$�!$'�|h��ʟ,����ؒ$��hG�m�o"�	���A1��Y4��|:����@���
�lD���澇���,#��1��a|?{��8|O����0���??��f�g���IB�I���/�������'���1?��r�ؠ,K�}���>�����.�h}���{��K�/���������� BH_$}�0{��`�����oa���Hg봜��mm��}j����m�����������D��\?q>�8l� ��2�����I!	!Z���}a��#b�� ����if%�C ��Ь2l��39�2&~N�Zia+�~�kD���(�n#�`?�dI��������G�$�	!W��ԑ�`�?��>@}l_��ς?��O��p�����>��!~?��Q?��F��>�_�J�<�r?p#��4c�~�����E� BH_Y���$&�1���~"H�ؗ�(3�у���_�����[�.�X�~:K4�)'���}С�0�����������9�0�������-o��3�dIB�ϡ�_b>O�>켍g���|�O[0��ٙ��
I@��d��i�$����~�~�0~Ϛ ���~�����|ABH_b_Q���4XW�>ϲ
�9�Kcu��T���1�/؆q 9Ԏ|�?�.�p�!�ļ�