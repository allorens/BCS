BZh91AY&SYl��p��_�`q����� ����b-��           �                                    h�� �^�QE�ް  ( �   �           
          *� ��x�J�W��J�UR���PIU(�D$�P
 
	�Ih�J�@�@@�%AER���.4��h =�1�(�I"���
U���}P7YĪ�l
w7J���ꀆz3�@�F��uU�������<6d��{�׌��P  y���罝 =P��%���U�������I$+���<�mJ%�2���:�@{� ��:�R��6 vtPrh
��� 8  �_<����U!U)T�)�(�}�����]�w�� �V��R�[/@N����Ó�����%<��r�4�@ !{�[  x��>��{�'�>�݇;�x>� |{�A��� ���|�
�}ϰ4�]��ЯG�   =�|R  zEB
RR$v���>��^��]���� ��O =�ï �z+�T���;��-��H ���<���   W��  ,��>=�����^�R� $x���=����� ���U/��2j_@<��7�t$7`:   t_>I  u i��J���R�"�鑠vtD�:�{� y]��� X��^��� ��}�s� �Ϊ)\�v8���@  �n�� �}� }v n��� 2: 2B��5C���"�1��av �    �|�H��m��B���R�H#�}F*vH eN� qܩ@��8�70r݀�� 8n�Rpl: �Έ  (ϔ� }�@����R� a���rM*�`��W �@��r �d |          �$hԚa240�C �O�4��J z��    ��U(�h�i�#&��6J�TH      )䤤�2``�  �RI��D����bi22i��46D�O��~����??��O�B��fZ"���+���~��(�bz��QE}� �����������
(��?��?�p������O�=��~��?��T����+�eU_�QEc�'��'�E{����?���eQ�*¸ʩ��8c �2 � �0���2 �
2���0��"00�c(�0��"0������8£�(8�#� ��+�(��3(�0"�28�c)��2����c c+��28���.2���+��	��0���+��2����(c!���8�����0�������28��#��4���.28��#�L28�����228��#�4��+�.2���#�.02��L�0����.28�� c�.8�#��08��#��28��c)08��)�.2��� c�0L2�����0��c)��2��c)�&4�c)�&2��c!��0���)�.4�c)��2��c��08�c��0�8�c)�28�c	�&08�c!�2��c3�&2��c	��2����&2��c8�0��c	��0��c)�&0��c�L�08��	��2���+��2��c#��2��c+��.0���!0�#��0���+�002L�0���+�.0�����c!0�0�28���#���2���#�.028������2�28���.08��#�28����0���#�����#�08��)��08�L�L�08���08��#�0�28���08����2808��#�08�c�2��c��)��2��c��08���62���08��)��08��������0�����2��c	�0���#�28����08������08�c�2��0���2���+�2��c)���0��c)�2��c)��0��c8�L�2c,��)��2��c c&0�08���08�c�&4��)��28���.0&1�����08��)�038�c#��28��)�1�$����0�����008�c)��28��#�.02���#�28��)�28��)��2��c)�&2��L�	��2��c!��08�c	�4�c#�2�08���$��c#�28���2��M��08��)�&08�c)�.0��c)�&60�	��0��c8�L2��c)��0��c)��0L8�c	��2����.2���c�&08��+��08�2��0���+��0�03��+�08��#��0��Ɍ��+�.28��+�!��#����#����0�!0����+�.0����������.0���#�.0��2+��2���(c#�02��� c#�28��!�+��0���#�#��08�c��#��0����0�ˌ���.2����.03��#��28���.0��L0&22���+�)��0�L�+��ʣ���+���� c
�0�2"c��8�#�
8�#�8���8���8���A�4�����c1?������_��#�b/}*�T��
�2d<e,L���:*�6��u�A�����7�
��R�%QtcѺ��$�K�"' ��=��ecɆt5�'�I�v��֋	�OFT�f�;��*|��sR;]�0b�:!�[2S��9����1���6��F,@��ܹgf�^q3� �A�
�e`#vN-qj�����XomPrO	Fw�;�O��7N͚*��Q�s�eg�3Ge�x˛�Ի�Ѧ-�V��\P�X,N.�į��ɼ*��B��ۗ`��En���U��/^O*C���n�������Q�)sYʃ��I�����A���d�y�j��v<x?v3�c�>��>G�o����S����WwU��C�e��7j=:�w���:\ci�ζ'n�6Q�9��u�Yu:�u�����w�;{�A۬]���y�Ia`��pmӈ�u��]���,���q0k0�O&�L�`�&�fk{e����vi:.1��l`ӏ7����,PӉ��b��Yݭ�m��\���*���~AÌvm��{��[)YE��-EqM/s��T62��⛝E�J�ה�f�b��-h���]XIP9�U��#xr��,C8tokF��w�%�4�,8�fq⏗zل�t��5��A�s�/����d�v�_t�^���_�vMk�v�Q(��6��Go`��)*e��h�"�0�ע�WH�W#jR�M�p��߸�����'^��* ��I�gBylp�]+"��Z5��y#k�z�[��#�(L���3N|�o��9� B�k/�j���;.�x.�od�c)�gM=�����S"���[��N}�ִ;�� u�fo5���}۝��H�9�G�����@ 9��	k�J��k&��9�Γ�[�tvK�=�J�8嫶^�#kHza�oj�F���ь�Q.�`�:��S&oOj����gp���lM��.�^���_?��;��S�m���[v�8[��65Z�.\"��i �7��߶��s{7��`PY��8�Gr(qԔ<�g��v@QţxM�SQ���ۺ�c��q}$2iy6�e(ɻ2���7 ��̍�H�Ε�d+bC	U������<�-� ">W�`�9�V����yu��T-!���-����2Pҋ	>���vwv�xW��l1Ÿ�.����-�b��0�ײ,]���%�F��"��f�kp��`��Pf���|��iy`�t��0�k��ٚ�]=�*	В�ڇp�K	3AYQה����t��敜l�*� Z{nŨ����+�96����{h$1m��ʥ7Ztv�oQ������1�����Ǐ�y` q��F5=vM��
����.��k��]nak�%n�"p;��ـ������s�qc7�E���P�Yq
�����T%!KS0�<*X5�7K���e�2������78�e��׵�i5���ۂ�'�wل��i��,�P-�U�-ݮ����G_�V�Y��B��S�ґ��^���Lv�h���(]�N.vo`Q�Cޫ�����������@}���g!j�dZ_�G�˔���p���K.��c����=� !E����nG�)�	;�c[��J!�MV��6�y�u��l�h'���'Q�L��I�%[FI�]�W��6�tO �`����y.}��x�*!�w�O%�w�;�[����Wn�Ie��WE��u��[�6�3�� xf��(V�2>���GqAEZ���qX��O-�B_n͉,#s���
ξP�`�#��t��Nΰm]�p����B2�;��Id��_�θ�������k�!�9���lx5�.#�oMN=B�Bi��f�PFE���ip-��wa�ky��V
�{�f�Z�
����i5��hv��S�w9�i\s�e�c����u׽�\��#n��Hy9������Ν���2�۳i�xs��JD1Y��9�9)���W&Ø��X�Ï%Џع�)μ�V����$�#";~8�����ԯq�7!�-�\�e������]���]��dv�L�'~�*ڶ���6-{2l(Y�ȁ#�A�/wq,-M�������AЮc�^����w+�G������q5w�uY�4\aw�y���7AZ��Scvx��={�;���vu���tQ��q9G��	�zU��^^a�Ц2��`»�&s�L{�p����	z�,��6ZɓO)xp�i�T�1����#����d�	�Lۓ]e��BӓQO�k�Y����v��/�Q�䚓�9��8�����j�X�;��<;5ou��>�jͤ�VM��@�3u�;O�WwL�E�`셐]'�Βuܵ\v ��ʚY8��xW�7;9-b�rۛx����3mH�"�E��(�	R�7��Z8;�扮�ꐈ�܎�E���ٗ'-�t�x7.��]�-ЦLD��v*�P7�ïh���h]��ԇn��k��(	2ask��������2}�-��D]�6��̩6'C�G-��G6N�1��	k��Aw<��L]�GN�n�OT6��%?<���0�e`�kn�j��M�]K ���I���������9�	=W�2�,����66����uok��n�UIVY�j�D��F錊��yR�wJwyL�҆�-�-;@>�n��dp�9^�>�X/��#��pH6���G<�g���g6���5'��ֽ7�,��|��A�8�D��w6Mp���� j}̇��(>OL��Pzo�)�q��-O	͹c�$�s��4��i��,�Gc5�;v�wr8�T����ܧ+�pxw0���U�'�s�b��=Yn�ɗ��_L���6�{�H�VHb���m��J�H��D�Eɻ�]����p��-��-�Ժ����	Ihb�X���;ӂ킢"�����r�.�$���h�4^&/nl�b�����ݽv���d��E�<������q�:f����v��n����m&����n��ݣA�Y\��Pd=Z�܈9l=�T��ɩ���4|�n�C�Xu��2;Ȼ��@�3��ټw�.�Ky`�A���2��Bp.�v�F��g1*1�����;_w�Y�Iܠ�i�ʱa��J��s����Z������S�+�3��q��io-ۃ�l]��:Ez�Ҟ�����ٚ.�J��q�9o'�����%�#��GP6��y�r��ǣ��]�w��q���&�{��w�c�hb�֋Μ��T��U�ʽ��r�e*oVǮq�oi��uΫ��3��b�����`��kk��O�D"���#���<���o;��(��2��ƯU�6�F��|�����&
�;�S�ᱣ�~���<(kS�w`�n�6d1J��ѩG�jA���ҎN�ܸ�hd���&2��YFe顲��(���RY��'0�����m��r<�$�s�n�4M�s/J�WcL��0��q��8_b�cz7b�4�^����W��S�^s�����lp��V���m�l�O���_g������/h�jq�ͽ��/�z��N��A�~���h���`�'q�bX�ݻ�������An�]�&Q�/78>��tt՜6�I	RO����ؙ'm�я�s��G^;�fYٲϹ�0��D�
x9����L��,@=�w��0��p޻y��hy^�>�^`�̄4ہ�;19��ƞv��x�gbƞ��wGsF�w#�vk�Q&��`��[�
d���m��OC����n�83��$�\H̋Z�gն����"9Ȅ����`���$2��f�w(�D���f�KKeT��s5*�-��Sй��pи^Ū�@Yѝ�^������R5r�`wk=�;h��6s+l�g8,�s7(��I�TȘ��nw��삨�_�ݥ�=������`gN�nY���� ���.�!��1a4��oo<�5�s:l;:�ml�{&���g��{��K�#y����^��׉μH���QF |;t2��Mv`�{wm�;y������'nN�nV�=��pg��H�ۇ��/oH�Ӽ�������b�$խ��������5;~�{�R�Luǆ���}��ô�/G<��d�jw��������k�oe����N;/r��4P@�@2�<��wc�`�i�̋��Pj���bH2�f�[�v�l����!� �W4����RU	�w-�w{,u��,]�x�N/�{�z����s|I.�����&�
t7~��ś6n�sv.O�'Hz�hI�7�����&/��pj,OV��um����G�R�S�ڍ�U��]Q誑L�C&��n�(�1��.��{%�xM�u˨���_�e�H�dЉX�� �n�������<���z��מ�ӌ�ΈC_L�fT11���v?��z��71�WO+t2x8�|a�}�\ygk��qD��s�|ix�̡��mb*���4�^:&����n����om��f��B�Ȟv���S$�W�m�6���ɶ�	�������w�o��v�;�Kw�l|J5=�A(��vuxe&ܺ��B6<�����ù�~TĤa���r�\(ud��1,ɗ���d�捽A�d\^II� �ƥ%7�x�F"��mŰw�.Z���ѡ^쏨{�����צb�O5���X-Gp�GD�-d]��+8�t-7Nnm)�2�˻��xך�)wQ��.�1�-��qU}׊��n+ם*�.:[ӎ7�˹�첬6��a�Nп�y���Pü�s�<c�Ziɤk�^ם��s��s����׼�X���A���zf��*�4MUol�~Jص"(`�a�Qe�1���"�܅�!�;��/,It�)99�U꣸H�oq���,g���u_X��g+wO:�¯oj���weӱ�
��5-&������Jn�����QWH�op��+����v�ł"e=�Z*����)�s{��K�S2��g�xR9N����8�&\����B� �·P��T�ƃ�Z 7 ��D���g8�g��J���k�T=�}T�'6�ݚ�w��,�>�۫(M���q��[��K����$[}�n���ǴiZ��ze�.WUa���GȎ�5sq����+J0�v�s!�-���a�Y����=۳;)ͪ��d��hً�U;J�p�+7��鯠\WxVz<-���Z��kA�`�+�0�k8���iŁX�UݏO-&�Dkf-���8�\r	�q�滖iJEܷv֌眻��4w<�ɛ���<6�sd����N!3x��ۢ)����p�]�>�������(��R���zh����V��m���y��R�kp^����ۑ�A��m��o�p�Ǝ�X��S�κ򸰜gTͼ��� <|	¸^�� �ɼؒ[5vTWF-�X�qH^M�y(�븪�B���<@������I=���v}��s���e�S`�u�n]�>��dٰ,Tv���޳�x������8;�0{lt���V5�s�j�b�h�*�VOr�G.��U;sÐ�bG<��n�܁�i�=5H��E����ߕ����ז��C�aĈ��"8�ٛ���i;nJ�L@ۗz<���gz	{zk�;�`妃J������;i�k���q8;n���������7J�`YO��Z�x��պU�v%�q�+c\h�k�Gd�FƜ�wGmg*p��+W�xr��=����5
#��ソ��V�\�hv|�wt�	Xu�[JA�t�`Ph����Vo9����J�����{^�_����w<�\s��z��Av��|�{h��lar8�]�A��/Ia3Mw��g\Է���ӧ\\/^���lY���{8;�ڏ��OJ~�%G��W��������w��Ӣ8�#"����~���I~�&��l���">�al�d�ٸ��w&�Y5��a��	#\kw�R�y�e�a��O�lDM��&l���T�f��t����I��i��9}���ǣ��qCs@`}p(^{fq���HP�����wB��>����܂���7n�M9��D�F��rm�gv�w|?��_���P�O�݆�Q��J{��Ϸ4'8��{wd������I�����w�HZ�������;�6sBi	��^ӊq�Y�q4���׀q���}o<3Ϧ1�q�E͓�B�K�յ��P��Ƿ���):��Of�\L:���Ӻ&��Sܼi/�.h%�N��\S2��逍���;ݎ�4{��n1o~�u�Rq�]�}0�*;N"n�E�\X������/ �o4��� �0n��"��{�x�
��w�$���mg^��JC{'x2S9�D"�zh�q���R1�<�����r��涍����r�JU���a�{T��"|�z�(`�<�xn�P�Q�_{iqz��.�0е�w��<Z�|��һ�͐z�gS1`�q�};p�|dY5�8�����Ś�	޼V�L����|^I����#�5C㑬D�Hh������M�M�ϼ���L�k����`�ag�G�3�x�֒�g{=�Q�qn{�ӬZrV���ⱦM{�	�-�{��؞ �C4�tZJމ%?�?~��F]���:!���Yf�]�{���-��2o?�޷{�z\����=�a��3?^��F}���Z�.*^A�V��P.�-����L�
�f�yq����5�<��oMo����}zj�q�Ǹ���O�n���\O�E5�cB�Χ�"M��D)X�{HW�㼖��:F��y��U;6W�`�s+��G�����|[ߨ���?51��gy����R�
~�A&�R����E�%2�TT�A� �D\�(�)iU�D2T�T��JP�A�G S$����V��iE2�D�U2D�$��EZ �R�� iB�V�JUh
!C ���D2E�\�DC!A�P�R��Aihh�)2E�AhD$2�2C$V�PJU�F�D��@�rD )R�D�B�F�EiA
@()A
Q�A�����o�~f?,T2W�\8���O�	@@pbX��BDN�Ǜ��v0 �CՌ�è��t@��a��m��s�g�Y�v#��6��sAbqopf��?-xn��L:�+G~��9�O��VU�[�����j�'���<�Ii�Y�}��4�#�٩��K����K( �a�A�x����ݓ5n� c5f,<�+{���_i�81�f)�n�d�[�O%��2�.�߇��e��>��H��`�`����1J�������v3���0����/�/�0k�Uf�[�"��t|��70�/X�jf�y�p2D'��U��{��' G#�'#xq�BP��O����6^.�A���σ�I��'�Le��D��M:x�x��l�1MctI��	ώ�BL��In�<w�i�����[���fE��04P��?� ��c��7��f 79�� &%�,ўuܬZ �#x�6JNs`("xAx���0LƸ��n�B�-o��		��Oc�"��$^|��b���8b�(�!R:*g���  ��\K�k���������ު���Ԋ�`,d�@�Z�%V8I�%xA��r������S�O�Ҡ�(~�?H�O��`�����G�P7�?����>o��K��~�R��9��z����z�z���QO7�6�^v�ny�s������UA		���g?���A�f��^���>�����t�	g�^o��ٚ��5WN���=�}yL)|N�S>P�dG��S�T8n����G�><ǂ���s��6y�(�i�s�P�~���D:�}��c�=�ڴt��)(R�~���bZ�t�E����LRr�۬��Ƿ}�hbz8�M����E'��~Ϟ������E�11� �Lw���Ya ����y��8�'��}Ծ�{$�zzyhq%��{�+��v����{ז�y��g���Y:��s=s�sk�@�do;�h<}��z���Ǌ�5����Qo؜	��vi�"߃Mn]��h��9��\���;����%��_�ޙ[�y�Vj��|R�O��h>�:��~��o�c���c+�G���;ۗ�փ�!�>X2N���Y\�hr���'&�|���)ܞ��H�'�����n�s����Tx��
���Hx9̺�6}��e58�]�
���Q�kO!�3+��&q���k���N�=&�ڲOb��(Y�1גp�6&�oU
�b;�K�����·����}��;�@�I!��� �}č� �����y=��:�n�����^���\ eP��� Wc����|�$U�y^p��"�_�glmjjlll���뮺뮎�뮺뮺�뮺�:뮺:���]u�_g]u�]u��]x뮺뮽��u�]u�_n�㮺뮺믎���뮺믎���뮺���\u�]x뮺�n�뮺�ۮ���뮺��뮺���]u㮺뮽�뮼u�]u׷]u�]u�]u��뮺뮺뮎�뮺믷]q�]uק]u�_N�뎺뮺����]u�]u��Y�]u�]{u�ӯN����_N��N�뎺뮺����]u�]{u�^:뮺���]u��]q�]u�]}�:뮺뮺��:�8㯷664��'�E�Mר�G�A�N���3����r]�`Z`��=��Q��d���^{�h'�>�������Ѿ&�}�qh�����&c����<��V�)��n��^����;�����ŝ��p�ϳ�\Ӛ�۞��F�*Y�q��c��sfndqץ��R7�{ �EzF�Gq��f�՜9w�]�.d�tv{~��ï,�f�&+��G����.�k��D^�.�œ�V��}�:�~�����e<4β����vBk�O�۱{��6�{g�)�s�Mf��̾Z|�E靳f9�ϔQe�;�Y6�9V1T���\ce�N��������̂{�ٚ0����p���Vom��	;ڇ����&��e�ݷ�l��{���p�F��>׽3�S�ݜ*��_�bw�?�H�ѹ7ݡ����$���:��o�?��ׂ�E��K�v��/�f�k>ea����ȱ3�SY��]��w���f|� ����������o��C��}h�ql�2��۱EY���������x��
vy�v��v?���3}����������5��{��ycV�^ͻ<�%���TS�'�8�홤W.*�n�1�h�Em���=�-���t�=�>�v�t�S7T�x.�TE�ە����ڢ&U/U�Lҟ��--MmM�Ʀ���]u�뮺�뮺믧]uק]u�^�u�]}:뮼u�]u׷]u�]u�]u��뮺뮺�뮸뮺뮾�u�]zu�]u���]uק]u�_N��u�]u���]u�]u��Y�]u�]u�]u�]u�]u��]u�]u��Y�]u�]u��:뮺�n���]u�]}:κ��]u׎�뮺��뮺뮺�뮺뮽��u�]u�뮺�뮸뮺뮾�u�]u�]u��]u�]{u�^:뮺�뮺���Y�]u�]u���]u�_n��x��]u�^�u�]}:�:��u������A^/0�ϙb(߃�Q)݀9C�bo;��4wgG6xr�T��D���*~ʻ��\%�z�wJ�G84H�M+0o���5�\#ĮRGC�-X}ͪ5{��92�w۞���1p�����ϳ)�X������i66.�;�Vf�� I�s�?n=省���Dբq&/���u6^�m:��wA��=��J�̚���0���� �L3�+�ӕ��߻�������>y������g�ɒV��������{w�g�HB�M������e�Lln!�G"��΃��_r�:��몞�|gOo�&ęH�A�l�֌���7�}ؙ��\���\���b������`"웳=��8��\���A�O/<{��N䜰�q�ȰAy�nc=)ý�㽹W���}�2��;�_=�f�ӻ�s�+;�@���Z��������ӧ���/u�s�x%cG)�ǃ3A�<�1�ć%�h;�z1��7O��n��m�$򽝪�F�Oo����~���p�߯���.�CŇ�2g3����W���9t�͟��{S�ό�:���M��wkݓ$�O����=�2��Bl�W��5�w<������M�܌,(����A��Y��ѷ���c3��.Wa��M��9��A��<������o+͙B������L�����9yh��{[�����E漽A�n������x�.k��;��w����H�7tYV�|75��f��ݣ=<��y��܎Fx�2&[��W���=��]�1gd<6-k7�6ٗ#,.r8.j�������U���Y��r�S���̙#��<��;�{�{� �)L���w��k���){�]�k͎v5����y��L�¥u����n��Y�݊��C�E�jY����9ge�2�D�� �︽�I���K���K�qe����8���!����>K���>̝��������o�P�^����%H9�B�AE������}�I�g�}�U�ɣQ|zK��ӻ����+��z�����������z8M�E���ތnp�</S<N-�V��X�(D�g�k8s�!�� ������B�}���!h8ڙ�r�}��FDs`������x�}%�hڽ}��;s�Y�Əҝ�{T���Jk7�{xxr�5�<��4{��<;�c������v��p�� �Nq�-�w"�h�����{�Nν쌓��{������|�s�M�]�pt����?p/|��o-aw��hJ�8� ��8%��+=��w��ƨ��sY�!���D�Ѹ����hw�9z�3�t����n��z=��n�R��֧���Ҭ<@g:Y�8�<x��;'0�$���	���"��w]���o0���|ݺ��C���y�Ө�E��k=��d���$#}���b��ytA�{������cm�f�X�Y�3�ѷ}��Yu�Q�����9�g�iz��k�5a���y���z�,ى�=캵{w�;��e'����'��OL�������l�3ޜbm�A�x������"
�dx���D��(S8!]GͶ��OYk������V�ڼũo����̈́@�H�p'�<�r����6z�קJ�a�z�8n^���Zo|�b/6>˳^�^OP�W$���9�Ou�-Zk$��n����]_����)|�0�����I1�V�x�*9��7��ׅnN�����؉Ť`�7�1w�=;�./ݥ�xߌ�+�7�A�,�K�0��)<��4=T�ݓ�xv���f{Ϗ���d���o9{�:���^�'wuk����O��+�M�JH�Ec鮢��J�������;wf��}V6w��� �//]����'vQ��������������z��y�8��27��6���˴��3w��k��c��=�z����r�am��/$��������S�7��{ޫ��z9�b�z�t�{yo��H;�l̄�ʳ�
� �z_2�=v�OKg�"o�GMw�׸��X���.UyeO%>y�z�9���Ƚ�c�z���웆�����񫯀p5�ü�j�qM�A���_f]��s�>[��������	�����pP�xs�{<��\5=u���3�=ۻNn���T�@?LWx0t�FOy��5л��M�GӺ�u,�^ɛ�{̢J9�3ˢďVlˌ����	��b�m��̝ݕ�.��X
���x.P�U=��ޞ��7ӊ�7M���ǻ=�������[rf����YwG�746�x!�8v���\~��+D8�YVTج�||0�'�njY�ުyc"M�～h�iEջ�#�֙L3|7~F^E��K3�U�u޳\��F���q�}w���o/nM��j�HU�|�(�W�Yu�<c���ϣ���|����lC3�z�^GsҿoJ��f�o��S�����癐t܌��h껷F��o]�k��DlA�A�9c���h�w���a㽬o5�m^[�q%�xx[)�'=IG6���1k�w��[=�j�E뾸�2��NOn{zyK�@���x�����I|,�����j���փ��^�{h������:��*�{��G���*�+��9y�kWHV��^R2r�A/I�S�CֆA�ar�m���޽7sn�[�n���<�*~y]ܘ7���}�ˏ�ݡo�0�ަ�Zmޚ'50��{'!����}��R	��;ޞu�<{4��"�yJ�:��g �K�k� �xI�a4���f񳜈l#�}�����[{�R���o�=�C9��QC%w=?_a�!:=v�tS	��w�=g���5O��LJ)��s����O���v,S���w������r͠ŷ��Ԑ����z䶠&�&y.阏���9����}�=��z�㋥[Fw�%�-�?n����8�T=U�L9�7��&�GUk��}>�����c���邽�/�f	F�\�1~�h��K�����]�{��7�oM�^��K��%r݇�0�Z��j��,,yz�9m����s>��g��:�F�~¶�g��_PB�6��%B/�s�7��r��Ft��A��k~i6��J�7��H2{xL��d��a�P(�#I0zz���;�V�O�^�K�;7��p�����>�Ye�<>�r	%=�	3�Ў��g�l��=�D1�~Ӷ��[���5��C͜���h^֨/)x��J 1SwCz�+w�;�O|״q�>xaz'��wǕ����9����cE�O����" ����(� ����t��*~�v��򝽔�,{w����=�|nJO��䪹���='�Gx��^=��#�?	�mC�So��?7��|x̉���@@�Xq�����3sF�͘��n;�xM�zW�����Oչ��?"w!<��MO�����^x�Ǧ�����W/n�[��$�}�0��ڱΥdy�G�W����z��6��!�}�|�'^����Ꮷ��7���Ĳwy���]�?z{ܺ��n��[�q��gv�Gn����]��{�Ǥ��|���Q{��!��Fc�J7���ޯ4�x�v(n�wfԖ��������o��b\ʻϸ����[�^Mx��Bj��|���}=�ױV～���3_Xsrz���=r`짲��|�j�hy|�����/Owjݭ���X�!��� ̄&g��^�o��.��١�:�j*�-�;]Έ�v�}�e��W���zw�=J9�zo}���L�>ٔL\�o��s��<^[b�&r,#���(�����dͧ�Z�k�/�˛��<�]�Ξ
��fr�;�W�����4<�rŤ�b�Fb�Ի{F�]-��I/��ZI�w�#�}�d�r�i���v����F�{���	gP���x<	�=�=��>U�&�o���=�}zG�E�<���ӥ�Z@�{�����C̟>�.�ůy���3���<e�,�����޽V�����ޱi�%W�]�A�.ޏ*�;�Xf����wN�.w���p��F^�[޽��6tZ�?<��wӜ�MxC�f����0$�L�k���.U�qގ,h^��!{ǀ���%g���Q�\n}�w-]�g�zy��{%�o��7���_y�ȜD�g��G[��������s��w:�q�v��gO�_���X}���4������a��J�X~��ɗ��Avo���} ��d�:�S�GJ^=xg����h���gz�Rgq܊i����$Q����A�#�����=:��Iǟ�o:JV��ޞ���yL�ז{�u�۾�oI�N�?Kf�������� ����>�q#y|5*_S�)k�@��Vj����]#C<t�/(���lrEFa�E� ��ˤ�� ��`�{}�Ʒsqj�n�ud���es+�R;��s�L^��J#�������g3|石�A�KÇ.��Argol]�� {=㋰����z�³L\�4x.����{����}׺X�Ϸ<w�G��������',%��_����i�X�"�ì$�q�R�E][��Q`
O����1lӆ�G���Ov{|��v�2���O�fX���x�?�rD��`���OY���e7=�e�ܼ[ӹ�hA�e���OL�ǯ��+���[�;��|+��pɳ�����1�nｶq:���Œv���xb)�n3�#/&��㧬�6�3�q-�s��g+Kgd���������.?`�dU�u�B���~لl�2=Nu+FoLT���^_f��+��6H}!Oz_}��Y_�C6����C�v��ׂ[�gz{\�.��3ҧ�����U���/s�ҋ_o����/Z�-�D����$���:�C޻6�>͓�v��ZױOyܵT��p�w�q��Z|�^���9ލ�qU����o]��{�3�Y�N,\�;\�t�;�FK�����N��k��ff���^{�{;ٯ1yo��hKs}�=m������v]+��N- ����}��Zq��:{f��a���˙��y�����e������`���8d�:ݰ�9D+;,�?O{�.��5���|,�E�w��^��=�w�_S!�P�f��.�^�̺�DW��\?�d<��ٚ���Ck͛3�w���'%�&��G�>�z�������� ��3�Z?��?���w�w�����>�?��vu���9����?�p��~#D����2���;'njyC,ak�3���G,qa�<�(��K?F�4���M:��d�V#u�Ms+XY��l�V�M���-�P̭�� �n�ƫ��m�kV��J�%v`؎�����4��N�����.e].��ڸB4/2�Y��Ll�k�W\bDK2.H�T�e�&�\Ԛ��KwU&Y�2���͘�Q��2:�7�ڷ� @�7ikL!	�U�v,�f���"kF���Zq&l�q-�`d���L���3F90[q������.�D�G^u�@��F�<�n+r[���)�I�*�GKX�Q0a�krl)ai(j[�V�z��v�CG$t�nQ��MC��iW,л[�Y�b�J�Rl2���.�����ر����Zj�������b�ɋ�Ni���C)luȅ�%(�^ÍB�[��ǽ"F*J�������P)e���,[�sWX��Qk3�� �h�M[��+az�3�#t3[	��jX�X�瘗[`�5�P�P�Jf����U�:�4i.J��4�PK[�+�4.(a�����(��LdJl��a���F���Ձ��C�4��x�Ŋ8�\F3]�cV`3a�&���Sq�q��R��"C
;f�
±�����GQ��[�UC%�$f�;	��M����c`њD��ŀ
��i�����ָC.�@�/\D*�ePݨ�]D���qIjԙ%�+Ms �vqR�p��^�bcT!����q��`�Z9U��%����I��J�ӰhR�X-�۴+��rS$M,��n�m^�r���ct�FkGY��f[�fu�[X�f&�j�U�CnB�hf�D�q���a[�M�ih^Y�Cg&��ƭ&jK��6�XToJ#�HYB�MMF%Mu�D	���3j�SGV�	�qYZPr��q3u��TZ��&�I]��.8(��E���K-��8��A�",(٦v֠ePlK���T�[Yt�D5����mH�� �9�BW�G7Ul�]G ^� M��5d��[.[��p@ع36��)Ś4���\Ri�my���&0�p
�.���%��@vZ�X�K�
�q-�ׂXe����AF����ٚf�-P��h2��AH��e��n����Uf �"k0�\#��3��	����+ah�LcVd�(��2Xbk�� hWGi0X�1&�eXe4��!6���5[e�H[���s]+�-`Al�[[���mW(q�ð���.4ڣ���f��7ZS�DZZZet��Wh��j�4���.����v�U�d��!�X�A4�U�9v
�@࡭��V5�aL	�MZ9�p�ұ���6Y\� ��c��5��-p�54]ZK�+s��*�����B˷l�J6;kJ	f�!�#c2k����Ez�4���Δ:�CXh��t��85ʥ̮ъ�e�����M^a�t��R"f �q`�m�[2hYRLSVZl6�����(v���\��j��i`��&�q�b\`�6�i^���k�4�&�-t�[�g&-[��Qe�-�-Ȣb�
k��v�6:��Cs\�ꗝ��m��uK��i	�YK�-,۪�K0"�T��t�,+Zhۆ�D��Kvm��D�E�e+�8��m�YF�
:[5Cb�`a��f���c[�����e��#1j�v�%����v$�fm���Zkk%-�bhd��̄fq�S�Mv��V�m���5�Kr�T���st��і��A����snu����z��Փ8[f`� 
�m�	��E1⮫��K���I�vrbV�3hAsKl�AƖU0�rS�"��S0u�2��K�m �q�α�d�]�j7���3H 7XeA1��M��l��z�LKP�@&{Ki�p+��su����[n��&hu6ʄ�׫-X��6�N؍��^&���4�2T]����жݺ�*$�8��.��v���c)-(u����h3��]�D���`�d�1�ZRKVf!�]4���0�]��"hhf�R4q�`��"�f��p�]�R�YQd\A��I�q�l��.��XKU�GSn�9�K���.�^BR�3t˻m����2�����c. �XGYY����'��F���Kr�� �X�)�*-�!���njpն�X�R��Z�B�R�B��e�eP�&����K�R3[.V�9�j�Ŏ�v(�M���Ye�����tW-�
E1�͚�`����5��[��bB�L���Ŷ]�MH�6�#�ػ��XK�IGMf�ub`��V�fq�.��l%QA�]]u��^�J�\�І�4xV�-T�E�v[�]R<�C�pZe�kv�Z2��+�.,�<�.��4ģ��ٶ��d�n���,u6K��]Y�;,rQ`��0�bRK\f˘��ňJ4�C([^Z[*�XiX��b�M	Lk�"��B�0p]0�sL�8и���H�)�X�i���֔F岶۠��ʎ]��a`�hs,�G%�ض��s�	�-t4Ʒp0v�hp$�����[� ��[QJLüb/o�f���)�ʴp	��Z��6\�	����*��k���իhҩ^v-�M1`�Ń[���0����q�!ͦŋ�U%L�m�k,k6b:���2bEt�iI�ȥk�GJ;���R����7[�����W$�X�^V�Y�����Ej���Yl��t��9�,m�5eHH�m�ncL�fb\�3@R\�)���R��i�m��G�ٺ�U����2a�Gf,*�#�؎��5�u��D�Z1�fYs̺��ɞ�@��&���D���K�Eٙ��葉��Q���a,XU&ō^��!h�⥮�vˆ��B,�d�P]!�Z�[�`kT��1�n�֬4��BX��`iS�\�V�X��m�JLƎ�uu�f�2��X�XUı!�䛭m[ʎ�5������h�&�X�ĳ*JH�[e�(�YLM�Ks��U�-Ԯ21��1K�h��E%�28�rT6�[�=s(�8-����Kif&��nu�KmF<��n]�5׍���Q*��;&2#��F���@��bV�*B�1�\\���M�x`VU��@���ȃQ�R���HbhJ�n�[K;G��Fc:�n���`�0Q����&Z�Qv(������9-ͰT��M�@ 3r4:�M�Ԏ1���1l�IY�p���fى��9{FVՃ�����l%׬V�͚R���b�do6ص�](�d��;m��3^�궗YkH��0��F�V��m�匼4f�7�����%e��o[ڱ�Z K�+̶�Lֆ��&j��K�ͭ�U�9��^N!��	t�:l8�l[�WS:ۤ �"5���)t��`� ��l3[	h�@�n�fm,���,+([&ر��1,J��E]n\��]���IGU���F�X�d��E�զ���9q�G��l�f+۶˩[UlM-�(�@�Wt��锻i�T�f�nř��S9���+��,m\�ԃ�L:i���\t�5΍�bJ[�Q��v�+K]aa���^%@eT�il����Z���!e؊�L��-�"An�2��-i)�T�Y�3D5ܗK�tE&U&k5�Ž�� �c��1��L�`�Z�Fm��� �M���H�n�[4YCV�$LL�ۦ�o6S38ZfRTZ�Y��X<Rf�^6֥D`��0KYV�`gWm@�����H�!4X��X�&��s����X�&B�-��](�a�:��+����]&�6f�i4��vҏ6��#��dF�Ԭ��ekZ,*h�7��,�y�\�.U�;DŮ�ݒ[lѕŌf%��S0Ö��7X.����Q�&[�)k`R�״�mf�/�u5��n��G \襘�:�#5���������l`DwնU�7\F�Dx�\��k�����	uH��M�ݶ2������MS3h�n�\�.	�o)41n��,�1�i6FT�8ы�&���B�2�m�F�nY4.�\J�02�T[-����`����ͻ�Z�iLgMteɬѪ��r��eݣ��h\A�P���ֈ�c�K(���2��H)ڹ�V8�Ǎ�D]��p+��&sv��7�6������9nb�f���;�3XTnڴ�M4�b%y�V�cSq�R^��U�Ѓ���m�a��i�P�
�͐a��4�������R���L<;2��u$ŋΎl�*M�
����ε�{3WY�Ѻ٣�#�2�P��r��&\�\D�Z�h3iz��e���8vj��\)��mҐX�5�:������lѺ�)e�fl������٭6c��2�U�k6�6@�m���7e1��i]�L��<M��)�8�n�����d�;S����U׽։�R�`.k��F��ہ�FɄÄ����"b!0]�����'�/�۠a�a)��D�O��ہ�)A &�TgL�#jx|s�:PŁ!2bވ�'���L~�>L��t��W��jDR�G��dV��p��c�N��:=��u��]u�]u��Y�]uק�q��Ȅ������8
*��bP�c��JÞ&�w�~w�߷{g������㯎��뮺뮾:κ뮽}�fEa��d��ʎ�2�~m��j}gvM�oV�\�x��JV�L�kf$~ou�.Z5:"�䈇!P蝠�IEH���f��TQZ�X��ԙ�[I�Z�B��a\����T���v�Z%�=��Ð�r�i��N�mJ�bҵ&N��"�W�cID�%d"�km�ۋ%�"���/sh2mJ��C<J��"��P�+���!�mD#R��IP�nf�uNZ$����j]�m�n^��H|�std���O�R1�B���/J�j�F�Ф�d������Yr�N.�{'���S1�&�C���O .����q���z({&�Y�L��'��N�L�Xʐ�.�����`�b`ܝ;������K�1{�;n��++oTq����(�����=q��n�K5�SVa��ec#�����
i���d�P��Xq6�s[�[e\�S,�&�����70��뀴��ek���G�%�еq�D�����$�,�� l�����gj���F�\����xփ�+MK4x��J�lئ�m�la��#�A�*YIu�6#�-�b-֚als�ta�fjT��Fٝv!�����k�XF����� ���Ϟ>W�J��e�-�F��nLKD��h�W,Av`���0K�c1�+X)keSC�i1-���f�\m�fZִ`���+2B�[����ˌ[�@�����j�[#f�٢,�4F�[(۠`!eY��p���Y�sf�\�9m��"Q�rɈu����&����J�4�a��-��m�u-]{Z�2�B�n�f�"�	��We�@��j����Z3L%%�R]LF멡����,3����u�Bء1p�&�M������ІSF4sV٢Me`L��Y+jB��1n��ltD#f1H5��]��m*�P�ۭ,6][c�"6MF�-MSf3WVY�C��H���e%��,f%�]l�`�j��`L�6��mf#6E*�XiWc]��W�WFǮU�<�<��#�F�"��Ў�-M�L/b��ŋ�
�8��fj��d[lL�ˮ�f4*D�F��\���*���իj�K�ؔ�e��:���l�ݚ�u*Ĥqe����,e3�R)�⹣�K�)�!H���%Ɩ�颷��.-6�T[l��x����5�a������1�r3&m3Fi��r�`�*Ѯ�e��4f�A �
R7:�6��V��ՙ��k3oņ�yf:&�1��:W��{��s�����f���tC��H�6ɚJ�Q��mmjGY�3CLƤ\:�ñ+���(#-KU��Tlx=z�)�2��f+3TA=C�6j�	L[/"�%�F��������S������v^U�����.�2�S*�U�l\��ʤD�tD8��0E��*�l��.�|�����`���߬����2X�^;{j2�Ǟ �H�<�6v��r�y�B�n�~\'þ� �Jpf����	�d���K0�{E52�Y����C��J8�ō������K��A[o�|�SI����������i�
d�5xn=�\�B����;>�M܁q�L��MH}��&[Z�/�C�+<殤X�s��l���P"%�H�6�d"ĀE�]1؄}��B}w9�j�\	*���	;������@�-���k5����Ћ�ƺf�Uv�
fQ֎�E����׻�ƳV���_^��,
�{2Ř�,n�hT��_��l;^KѶ4�r$S��&Iy�K`:��`��&1�{Nt���jf�5����XgW�|������հ���Öx.
�=y�x:n=�<5�t�Ǔ=e��ż@wH�LX�7�H S$"0�$�su��e�]��FW�d�ԑ�i������W�߆�2��ǘv��ۋ��m�g/u�� �-$n��$:�U�,m<L����c�g�z�~�g9>�q��� �a��$�2텲'&�ر�Ϳ���,���~�>��H��*���������}��Wv4�q�K۷��H�@wݙ��`O���� ����&[lY��SW��t���e��.�	�6bE�o��/�<l2Y���9����	���y�I�W�xw|==T� �%��<��3����wx�ݑ$�����_6�K�x,�v���`y���^�d�`a!g�A)�b;P�0���1�}:����Āv�֖Z;{r>K.i��o��||1`�3�`?
N�r^���x�;�կ{��;~��7�gT߻�v"s�$���D�>j��b�8��!��x�,X���Ā@'2ݠd�vd��
IT׆�r×@�D�Ñ���R���e�Ͷ�hzd�_��W��md�F��s!�j��hUK� \>vm<L���Sِ` ���aE��|�$���,H*�r%1@��A������6R�Sg2�l �i��(�$9Q���D�t���δ�i\,q�KMA�kqS5��� ұHB~�ϗ�Ȧ֭n���x��fK�����%�/Z�������ҧ�Zx�d�W���ڸO��W����8���A,��$k �i�$4���z��&���F_^�K/�X�/E~���>�2  >���Cj�<�Vo}��$���m����;0�'�$�������,4�
?NC��A2�Ք$�A5������A��/���˓no�۞�����/=��=po�׃&�����������{8�BswR��M��í��^��;PO-���.�I�,촐�T��3c��C�r�����x�X����jd(|���W@�盙$�z�DN���.�K��D�|�u.�((k�H�`qIH�3!.%�۪�,��9�k`����}C���@>��	;�� Jc��mAK9�ȯk�|�)8@��KH'�>��n6%���?��&��D���ǲv@�d��g�L1��x8ɔ�{�,n�/<O~Nd��"�ƃ%�����$�؁��$�2Gn�F�����A"��a������<�-'% ��O���o�0f�O; ��J�H�L��x$��7Mcϖ��HEĳ����A)��_\�LB��`�ygi3�-9Z}>Єb誊��@�{�RHm������O�bi���1�v$��O��"5v5���˪�)�e�W\X5\�h�r���^�sE�>����������x��9�1��Xav��2��)J� �LL&,�8N*�-�g������/�k�51X���R�*˲h�pqy\]r�{˥�#K`����+�q���lh�e�4M2ac��������͋���h[�`��Lː���ۗ^-�\�R�YP	hWf�H�������<�ij�<��2��:����݋�n(SQ4�L�1i��5�ӯXuD���Q�1��TV�%��h��ڙ����[� .&�br��)�ݮc�ĊN�+,is����3���C+1��Y[2rEɸ���}0�D�Ç��<��cI�e�0����?�˳���>c��� ����I�ݙil�p��uV|t͜bX�Pմ"�Q
�2��H6��Jc��b.�p�_�lM��A,u�a4�S�9������s��]�#¤�,F�<C`� ��ɒ"�������֢����	
+q'% ��h�З�O�Θ K�y�p�W/��'��gl�"�݄d�q4��Ny�=n��<���>2�詈PAr3i���)6x#,b6��+�W4�-f��r�����op�CB���H�q�	�����8�	d�ݘ�d2�o�6�xxR���@�q�2]@164�{u]�Ӌ9b��¼�K�Gح��w|�W�d��5���������9�Z7(�-�Y���"N�X��0i���,B�� ���H�����xyc�}��{�tڑ����xb���D�X��� �;[w��rP��P�	��fئ$-�,D\�ǡ!�D(OT_i�Aq�Vn���~md�eT��Jc�W� @$�לFϔ<�z��5F�L6D�)�0��^�:�I�d�Ǧ&�N�U`%=l�$n�0ı�ǂ�9p6nO�I�B��� ��%~��o�gʵ8�A�U�k�`��C�j�iF1��j�:ɮ��\���
<�w݉bM�A,sq�	/>�"=�z�N�D��ke$i��/���&B�%�Ƹe�Z�U�� �$m��K�� �K��-�[�	���%ė��M��_�$H���d���^��١����x
�`���k�YQ��.#���5=�bT�`��yv�^�,�-9<P�~��!({Y#��/�_`�^A��3���%�ر�����I ��\�C��K�1��Әi�����}��ď�<C�	��\�bA3_rE�뫡^1~�$���� z�ߗc��-�U߂1v� ��d	/b���^�Km\c$��q �~�̐ۣ7?5}�f���-�PK��	-�t�^���S%��S��ګ�X���H�񁍧�����a��Mf�/�`������� �s/QǼ�/�H$���I�9��� J�h��~����B#��"�0 ku��,�@>8�Ha��K3	!�r�7��Lc��e�'�鰰%	,Z���� -���/d��&B��W:�@$��ZI �£�}7���ŵ�?� ����G��X��$�	�>�W5ۏB�
t��p{�:E�	%V�y��4�����A��6�$���>�^�1հ�6p�G��>��;<�&8�x�4�{������QT�c��!��kbš��ꗀ]���"�9�x>�=2�P;z����b��:%�")%��<0$W��H$�l�g(ίFeW���L�b�:N�l��:;2T����
��h��%�\�ˡv���E'χ�O�C��P��}�I �^�I�ظ���m񨧉�Zh�y�Y � ��dIA�x/a'E����{b7;����� ��.dy� �݁�_\����ND� '���p��x�*Зy��w�La�LkrD!43f^v�Կ��B���쥉mہ���}$<A0�	f/��5��f_�%�����$�d��|1�A��ߣ׃��{8��������@D�$��[9Q̲K<�fA$�����~�{���wc�~�<�l.���gC���:)�D����E��/,��kd��s�y�9���(	������L%��)l���G<U?��B����n��x���_� Ke��8�?[�H?��mF�a�6Z�c�7X�`\�q(��љ����G%�ٕ��a%�����\SvиɆ
��Z@��.�)-��͖ɵ�X��1����c"�%�6�iM���f��0;M)�cxH�����MC��>.oOZ*K^�5j��!��,�r�%sLฃ5�p�B� XY�����+q�2hW^46)�FV�E_;J��[��$�X�5�����-����5�Uv�3L�������#�0�>���O���ȱ� �͇�F�{={j�ۏ�`q��=�ߨ.��|��oR{�D�Ꜷ;��}Spߗ� ���O0����9[�����O�ucI�%��`��da G�$k����S���h�{�%2M^V`�I��l�^7,:	'/��י��:N�r��=�Yc��-��� ��-J�4A1�hy�\�~��8�>v�l�g;��S�eV��s�x�,6.�$ܛ���S���f���q �m�fV���S�VM�K
,'�Tߏ�}�ۨ��z��y�V��J�b��%YVb���d~�ݻ�5��!~_Ɛ$m[�o�5d����+6(���F 3�P��s8 �_�٘\�q���|�|G_������.	�]kn�gWĒ�qy����_s�:���������8������>c���ږ�q�55lX��(�@6����\F�L����4�A��5m;zG�H�Z3��Xm��S>w� ���݆�/i#k�,e�#vd�{.!<t�<���O~1�a�iu�c�L���	�פj��iz���8���D3��A$��<:&)nd�A�W
��U��`7�I �͙[1��U'uD�XK|ߵ�k�4R�:��Nu���^�WQ`��;.h�W�����ك�Y�׼��,Y=��8�k$��a�[�N��oN��@W����d��"�}.�:%�*��9U	��f�o��z�|42
j�`���a��!������י �F�"!����&�=2Xi��H���0f ���^�)���F�݊^�.|��y��ʽ��{���y�kO�\����Y�©��}瑌'�|J�>�{ֵ�W��x&��'����Y�����f�m;�%qO��U��������fř�d���^����;���z���"��#<s��xeݥ,�#��ď>q����b�����e�4��ާ{�<��9��p9����L���G���f�~lg�\$Q{u>l���A�o @�p����V�Ǧ���{�s�m�f�W�B����P�/��85�Wg��vo�у�!7^�\�<z^��!�g��&a'qu��:�����x3���ӴA]����Ü�F�a/���J����Ǵ+^���S$s����/�J����+�ɢrO?+3���~+�����~5�������ܝ�G�醅n<��_���G..��F����A�ʳ�3}�񮹩�{�|��~{�ٖZ��ٯpg�W�Ǐ��a�qr@`�^M~���X���ݜ}�/s�<9g�)���T��h�댵6q�r�n�7�K#Ha��*<�i�M���w�d�USN��X���×p����/]��:ǻ<9N���Hn�+�Zw��̮�����3�Kv��|x��{oM���r�;��}�F����N�4��7�@��g{t�{�!њ{�ױ�{�Y'�����\����<��r�P|~�<��xvNu%����x泆��4����'�fn+��Cٓ�*ƕ���f����b-܆��{#Q���g�|ٟ=�`��v��}@�Β>���'uSV�f�'�h�%�ĥ`-z�&�ӹ:����N�%�vq�[�����eH���w��v��׶}�>>>>?���κ뮺믎���{>s�,�wκ��Z�݇��(��ā�R��n��;���$�NK�y(�^��A9e{�����:I�Q�,�l���TR�VvN�)�᥼�o5�7�5�5���������mllu�]u���]u�νEg�u���'�<`�[�p^yye�Dfu�����V:�VϽ���.�c
��3hj����w����;�ww���{�2s���d�����|��V��>A8{�׶tTD+ڏ'����&�,_{fz}��Ђ��9����vqU�����oKue6m�{��U�$2e�_�ol�ʌ}d�@��bax���y�58vU�Y��J�������ϴ5D3�,�޶�:"7�n�PpTԥ԰������lD
������J��xn&)9,D��S}�ו2y�Ъ���25s�}H�a�)U<��ϢBa����T�jD�!���{q�*�$��*���.*6.��J�*�dy{6�tl�/Bүǽ�Ȫ=�QR����BsK9�I�\�/(�5y��rȈ�6��fG�[v��\痵r��N�]�O��;��tuӋ��맩J��J9�|�OR��	N�~��w@����~ �T]|�<�!TF� �P{�[W��kC7�R@T�ߟw��^�8K���2���Ȇ�,�d*�,�6��q/3haC"�y�D_O@a$0����pb �N�Ǡ�(��{�Ȇi��	�D!�9>�nÓ|o��y�����Fu�z��.�O 2p#�ξt���;�%(2��z�R�Ҽ0���)�5D$����r`�b�D��R�D��Z�aTpj-&p�}��5���3��xɑ�n��I;�'���D�~��O���FH�}�箣�=�$��u�}y���\�^�%=����Bw�)JV}��C��z7r��VN��èQ#F`�� �� E���;�[�n����G0i"&:��w9R�&{��9)C�`2\eotAf�$�!���u�׍��x�z3�i
!���(�P��x�&y����2SӘ�Lf���>u�D0E��JW�톗��6< =�'�9|뾇 �	���;�%���R^;�N�K|���-#�9`H�G��.��Ĺ��>�f/Pd�'~��O���Q�K��0�q�
,�$#z�0�L��P�l�7����Y�7�P�p��Ȍ����a���p��M,K�]�i$� �>�7�9ۦb��I��U�a��)��}u�8�=��q��J�Ra/^��2"A`	4��z!�u!׃
#���|�>�2p�(2\�y��Or� ��k���fV �ŀ��=� �Pv�a?}��:���(��Ε,|�q���1K�	`d��\`��E�I�gۓU�v�Y�E\�"0��YT�>}�>�v
5�5�>������?:��z�� ��-��&�`�-Y��,"+����zJ�s3��j �DLD	ؼ�c�yC���z����]��XY�us�g;q�C$�>��6M}┾���Έ�ٿs�aE�;�7r�"� HL>��שJ�!6B�s�Ͻ	��H#ޯ,�pTm5M@dG�"�c��w�a�(� �D��%��&JQϾy�ܽ���&}��ￗ��>��w�C��A����}�R�@�p ��X �D�dC
�yqE�藈���X���r��_p���5}Jtf)������������C#w��;����0�O�y�Oql`�Ӆ�փ�"u�qā4z�K	!�a,�p�hODC�D7�`����ɇ�3�a�C"ù��9`)���?J��� ��Q�
s"Ha%��$#0��~t�ݽ�L4�d�o�=�f��{
�tw�i��*��у�p����u�����*���/f���M#����U��8V�7��p��ǈE$4��BG��[�D�ƍi��,�V���9��'s�D�֦/i��v�0K k�	t6��ewf�U*�*Č�ᵹԉ-�	[Bl��ʩ�:�n�Bm�]�x�"	.�\��kUB#Ζ\AM�LVՋ@r���m��[�HV�kPq���v��u��c�-l]"�l̳j9k�R�diU�r�e���R�ړ� %�m�J&��.1Dn�ЈT�3Y�A���[�(�
�]����vj;d�-(�3Q�+�͖0�k���������>z$6>���:�}8'�G[��Od���.I�9&|���I6JP���DtU^;��0��E��Di
g@ɜ�9�r*3� �E�n�H�^�� �BN���cX]>C	.Y��dϒpi�1!���,XCY(Z9׿���{d2p������]��2  ř&��%�O'Ӄ>�y���f-s�{�6En�}�C�d��>���ܹK�'��ΚK9`��,�C���q��b�WuDB| �L�R�y�z��J�,
b���,XB�Ԑ(б�pr�B�1�Da +��,�w�>��q���>@dGL�����Or�2�,tl�E��X"�,�6�xr�۝�`�Z��k����
"!�yqE�藈���X??�=%31J���ԥ^{��<ߎG{���������d����x|٨�Y�dC�q��d���u����=N>y��Vf�k+�an{�Kb	��;�&�Teu�P�j;�W�ّ*�.~G!���{��Γ�;���������k��$:c!/�{�OVI2r"�q��5a!!5} k��)�,���P�"(��j���"Pa�Ͻ�����{a��>��|��Ʋa���������g�����O�s�$˫|�m���w����&(�S'$g�Ν��p,�P�nҁ�O�ǎ8�9ׯ:~��C��%<Dl�d$�.��e�>V��[*ǎ��e��#�SE��^!'N����]��vt�3��x�TΉw�_�M��� C;s�H�d������I.�x�TԵ
�o�;������x혉�}���y	,�-�ٌ�J)LCa`X�K�5"l$��<�K̑�����|�3�5	D*�@3� ��5˗�
(�e��5�JR����d����v��PJL1�()g�^�M$�%�o"@E'gqm���6���}�egs���6�$!�7�R\�PVW��p���'/!3aL��S32���6R{�k
/��D�Fog�WH�HH��ȘgpY�	F�H�
�ȝ4=�§+���L���א��qĒ�~[�aAQ�Cċ{K:�y�x%׶l)3�T�f����$�&Uv���p��:z��Hܝ�����ެ�'���ư�mm��z{iI�$����4�$E����sչ_���ʮ���#�u�u�/�w�j,e���S��6��o���Յ=9*l#^Qg&�������Ukr�oލ�n���������pq�׾��>%�wr{��J)"��"���ӣ�P!@�r�x֏Z�.�܌�?^����O���D4�`�$�V쉦I$��tu!7�Ũ;c1�4:M,���ƕ��;�����.
w����Ԣ{e��N���u��j̠�0��y��d'��EE�@�l��D������P�@>r�q��!
�m���va��i�1���hWUE��l])�>O�������I��;��Ԥ1�ɎݟAS:/9�=��q�Ιf�	_��L����5��yl�R�?P�M�g�^�I�6G�L�ס��?4��w�3����!s?����6�L�\U�|o���]��fiE��$��[�aAQ�Cċ{	gVM1��	n��I�3�f�����x�P�����K
�,�ַs�)	&���໨��"� �� �ѻ�|O3/����F���4�H��� )H������<��Q��$��W�q]��.��➚�:3���Gz͞�� �Q�qg�=̱�}��$X��4���Ӏ��>c��A�&Lȓ��B�!VH"t{�(
��"�J���9���_��n�c2&��y�b%��ePK���W�ҹ�[^�Utx�_�9'Z���M��[ȚTYF���԰θ��y�4�7V1����l���q�໸x�F�13��dV����Y�I�x��:�eZ����Q��k��P�h$���Y�(0s�/Q&�Q��)%.n��Uej�f�3��y¶wt�zbL��A1+��"QA.��Q6�'�g��|7	������D��{u��I$�#^Ǒ)$��|�����t6���C(����K�2&QI$N���[�aAQ�Cī	u���Ϫ�n�!+���@'��d�H"�7z�)���C{8
�f(�]��$�4���w�.b!xx�����Ƨ%���c]�����[5�H{�$�H�K6�SK� �ޢ�NUc����JE���]I��麄��[�@y�'��z慑㦐ؗ����9Y����Z��~5�����Mjs��4��9��1�`g�	<~y�e�(��k�s�iAZb7�y���޸�q���<�_R���g6�U��ʻ(W:��v�L�]#�u�"
F�.�F��v�R]���9%������*̱Ђ� n��[.�Åj6���U��:h#�O)-%��\̨],��LG�9h���D�����`��.�U�6���Ãm��M�-Dm�3�*n�����ر��h� �k����Y=N0��	pxF�e�.�śLEIB�[�Qt��hՔU�&�_'����"��w����}�>z�QhP�ߎ��%��"h�	1Oq�]���:�SDtHBI 	��M
A� �՜N�/��߬$�;��U �|�;�xp�޳o���L��y��"��7�I ���w´7z�������.^D(0������)�wt�n恤�	S��Fgq��x�\������Y*	$��MKd�)"*��'���x��O�y#ǃ�٠�&"g5�R	 �a辬c���w}�2�^^������H@"o����-ȇP^"�NO\zl% �g<��N�_g7�ͨ�Q��L��Ut)�c'�gމ2�<��̗)�$>�[�Q<��4Ҙ��i��M��˥�c�b���S�5�.��������V����o��y�"ɁW�L$���gtI���޴zfͦ�i����)%Q�BMSE�����Ӽ?��l�[M:A-l�� F)^�����j���E��>�i_nD���G�����+��͝�Z1p]Ŏ���/�Տ���eU��`�`	hP��Ml���٘8g'�_�jw���mnȚ	&I}�D�kw�H��$��{��6���}���XO8N���OwiD^Țd��ǉd�$��zG���.����F � ����z�Im�����$�ps�(O����nC�U)�����f\�I��hx$I���K�bL��L�v���6���[�^\��$�6��.:PA�.�=��2R���^D�ۈq�ˢ���h�I��L�(n�I��I.�y��+|���GB��{�����L�s)�-D�.�n�4p��b���Sd�&7Ze�����u�]cW��o��z�'�^$ ��m��tw�����}~1��y&����eL��c�J���YgNwx�"P��>9K�^XJ@%�lٌ��ǹU�3g��t@$���[/���I%��-(���fk�	����y��y��vEEϯ]x���~w�! pH_��R	 ����j���Sꂸ��������"��`�;����|O�ٜ���.LR��ƾy����Q��V��z׫�X��|�7��;8g���p���ʙ�����$�I���x ���*�� ���W���
N��7WM_�R�;�L��m�HZ΋�z��RL�U�7�W���f�j r��I3NwS
�ý"_9�JR����ύ{�V����6F��a�ä����2�	$���m�4�'��
O[��u�Pdut5^˥(;�����q֋Nv2h�D�,�&�V�.�`�a�Y�{����֨�"����I$̂G=�"RI$�Gu
&iOz��,��ӹ�2��wp���D&�0+��a��Go�����:h�.��8�'�*ُ=����� l��M*�����
������4������C�B�x��g4I&s�Ud��)��p�m��dV�� |�	$���J�N��w�U%m*�l<;�wN�����݆��������G�יI$����B��:[L����?�{N*���6��<w4Ӟf] ���f�����0P��똉&=��?�K���^+lJ�}���GJ^�:�us�g'�j�}�:�7�^uU���:�x���ǂ��y�������}X~N	r�C���	D_M0��Iϵ�[���=�i�mn�e� �q�RAk8gzXI>I�{"M�!���}��*S����)b�:��Tx�p�0v@�jE���ͭ��L��Z���_�r�O�>l���@�s%[O2�A-�ɡ����(��D�d�{��G/3E�>�E�/Gu
���ݗ�(D��������&J�/|q�ug��:I����$��M�PEgA����L�g.
zJx��h���)1���A�B������ ���x��	Ϭ����tS� `I.��(P�wv��L���p���<D/x%�o{:�'�$�6�I-�ɶ��d��t�GD�*��ևt�/7{ދK����RH(ܪ�4Rт��èr����O<�$��{���F���w�̈́�tȦ����Y�'��2� Q�k��vg��0 ��I�\h����ׁ��yW �W�BvŞ�ڧ��)�=ς=���O}�2��1؈ɧ���=��ڐIc���5��m0��j-���Ԣ�{��HRd��x��F+�s�_���X]�� ��%{輡X���:�We�{}L\�|o�<�g#CĬ�\%�=�>^ӤJ}2��S�V{/������Ϻ<< ��{<���;�/�N�v_��x��K����N��c9��6i�N�3����]���X��PB��ўQp����q����^������_������/>��>�'��st03��t�kj̘����Kr�����5s��Gڮ�Y�%s�<}����8��iÕ���t��o�����c����,9�f����'����y6���-Q���2+ӻ狤�y��$��>�����w��#��ЃgcC���N=�U|�u޷����-ўyr���E�����&��<�꺭��bQ����څ���+N���b�� �)����ux.6�r���M�y��x�����A.	6��P��c/s�e�ƩY.��ۇ�y�����/��8/Q:n*{w���|8� ��;����ڙ{�}��&6�7��y}}��^��O�
C'��;�{�w�&�DOމ��p�$Lد}P<2���x��pԶ(_���q�x �P��r5W���xzU!(�'bZS@�D���;+[�\��K��.�;t�j�����@cmk������!#�Bz8b^{�ga����Q%X�Ȩ�bŠ@�(Q&ME�3��M[�e@p=O٨���~���z���l���ōP�P�����WO<�cRv��Ғ�Tࢄ*#L9�B(��� ���0kΟG�qdh,P�Z�` �� Xrw=� 1�h��q}4�&$A�b
�+ZŐ�Jb䂀E*u3�dEP�WffL�Ng!r��I�����H�:��\(�d�Q�������������㮿��������u�ۣ���~���>Y��$��V��̊�$*E]F��W����"U�xV2�"�wݍ�mMml�mmmm��M����[[[[[[[���~:��Dz�]u�0��b�YyD=@秙�URas�ʃ"�Р�$.�"��G�SpȪ�ڞUS��QEQ���t�*��ͱ$�O��vT{�^�B(T����#¬��H��R?P�z���W�Z�.DM(�Q�{��^�#��=���<,<�ʪ̑���$�����؂^!��"rtoq�H�,�@/mI�IEԊ��v{a�v!xtMqp-K<Nz�*#=(�h숵.(���$�T*���W���J�g���yzys�E�yVeEE��g�6�]��C2(3"/v�*�}��1R(kc��G��h�!��S�Z�x]l8B�d�'�U�I�m�:B����~��r�m5�b.qv��7:Rm �R�HEd�͢����lj��8�KF�Sj�^aclK�i���V���m�C6�P�TmК\��i��^�`JʴZU�֣�%.�����.�q�0v2�DѐJ5(A��zYKkl[+��B���CB�:=�L��cf.jĆ�"���.�i�rl �j�͚�R&.�m�+�%*\]�I�JƄU��6T�t٘���
Q4x�3JKM�!,�Y�n.�䆻9����K�2\�lj2�5�B�Wl��͙�d�v̯%f ,�`ښ�%�ֱnK�+Mv	�j[i�T�h�dl�`d���]�!�R�-�8kĤ�D�{Kz�u�/YW��6��F�� 7�ҖjQ�G-(R%��*�n�ڰ���̡�J��:���q b����(�m�jku7e3hR�f�1i5�6��W@�4Y�;m%wi�5v�6�h���[jjD!�v�4�
������m��+�L���r[[�2�g[Cc�`��3�Tдtm\�
�Y�e\��e�%�{��l6i��d��TmDX�ʺ�Ba��٠a�k
�e2�c*4Fh��Q4�f�.�B4p��nfƺK��
A�����T�m0�i^�)ăP������Y	���Y��WKh�#�[1nH���f�ZJA&���F�-��SWj�ʷYA���Zm�e�]Va�\qfZ�U����ec٪a�,D�b�ƍ���t�9\���`d˵�(鐷E�� h��5�+���M+�l�RQ�=�"��YU������(*�E&��W�D�ݙW8�#	I��K	]�%��3BT�.Q���J,�;�Ve�e��G8[a.2J�l��Z���i �2�-ԭ�du]a�Km�����M�������0�.)]�$:��fhJkGCh��,���{�^���={v8��|~����9�+���Ep������*[��f34�:Ұl��k V�PY�&�"�.�����6֭� ��jg3&�5t@K�n۲q�X�ъ@Z3W%�\左 ������t�Ĥ3�̙��hj�Qb�6s�uх.U�&�M��˜ѱɝ�q��Ri��-,�:X�fM�����C�S�k
HKǩ�x��i�|qlp,�]ift2�m��ٖe�˵5�8ZB}�����Y��F���ԁL+gwK;^'Y��$=|�!)W�}�vkga���B�A ���)*�+�]�D'x.�OIGkȔ�ݐ��]���\��c1����T��$�3�<I$�����N������ѽM��MzF�\6�Z�B%���O�y��(;��c��@;;�{��F�c�h��6Hu�I���t��M-.YU��cM#���f�;�F�L���͒Y.�x��2!;;�\�ke$L�7�r��Z��n9��nڙ�"�ud$��z�\<;�A
��K��e���cO�K����kk�Hz6$�	
	]�ȔRGczER~�ڸ}J�n�Ι����lo�#4�Te��]��0�L��*ĳlK���ej�љv'��}uqv6s�/���� 5���@H$�����B�(�)]��l�>��2A$�u��Xѕg���;�P���S=�D
A'��k�$l�=ǰp�@��riw}ٺ�{�Qĺ����ڷ�����^w8c���eC���s"0��[>�&r�ks ��~ ���{x���x�������,e���_| �� O�B����G��ח�TB瓁��`� �u%xk�������%�"R"z.�4�L��{�(�3�x2�\q��mD�,��[]�E��e��H�(<G������>�v�F�K`bq���|�yyyd�����PȢ]�Q�6ܶ��{c|���'��HH��͌m4�2ީ�7�	��I�A.�x �z��>g]R��hg����!k���U
jE$��D�P�A�ٱ��^p�4�����sa���B!i�D�iWSmn�.fՉE���tX��u�4ѻ��<C��<<-�l[�H)C;�J�D�I%��Y"�Ue�d�}�i&�� J�N��7B�$��b��C��x9�J�(N��je��I.��@$��߷�L��@/Z*�ok&ُz�e&��s�仸x�M�J|��4J	gcĪlh{e.��ν�x�sf��6�F�_�4\��U��r�3���f�y�yVƟ4�vh�NS��O����-�#��f)Sİ�MF��f��`&�ǀ�B�x�����s���3 AdvP��i$7�I2� �꒬s�������Q��>ધ����M���MH�dW�bL��I.�r�QS���IC��ID�	�����N"����y�@$�F��Pۤ�A�kI��P��o4BJ��P��-톂fp�z�?z�g1U��uW��B�!4^)e��6�R�,���B�.�"����C׿�w�"�k�7յ�;}�`�H��x��I ��v�u#c�j׉�Cl67��M�}�ӥ��@I��B"���x{̗E��I*j�YZe
�c�ޞ4�$[3�M2H$�0w�kД��y�Z����Ͷ�;��K�"�h�E�[������ÿ$��y��Yܚ*Nqۘ�ljD�>�MM2I���Al -�+;�����uvJ��"l��ڪq�:w3Q�\msĤ�%�י��xޖA����O����G�S$f�=���E�J�|�瑽NpK�p��ǳ���W�g�q���޸z2��O��|�ŵ���ǌ��	�#/��a���]��3Os���nk��߯�<�@��恪�_�ٶk-�W����A.�y�RIdwT���=��޹��bT����߿&����r�&��cIZ2]*1"=w=�&��Eՙ
A'��'F��uܣ���ռ�{�d$	$�^����$��u
�!��x�gC��e���2�L��c��<��w�xxN�(�zJ�nhL����#p*۬�ݯ�) �$�A>�P�E$�g�"��A�u�ēEWs��N���n�-�y�($��o�,�ֶwO>���E��قM��Y��(�O���|�Hs]h�=ДN��H��3�&���NC�k8A#�� J%�}Π��IotI^���f;��3>S`��K��C>{�� X�6��}ؒߤM�A,�Ћ�C�8�`$���2�w��B�@ ��J�VP�� ���5ҽK�h����G�f��L�F=��)�ޒ(�K)d��{��v�ӄ���g�6`ڽ4<uy'{���c�a�E���s��b@;��zb�&����H�����p�Er��>�����O3ǂ*�*+��]���9�:0���.=��h�s�]�3Xhk�K�bR
��]�Y`Q�b\G�j滃ij��bVR�;R�D��f�W^5I+��t�L�;m���j[*M��B�BY��h�d�5�˦���$� ��A,�Gj�����ٖ���h6��kr�.���A����!��мT�-Փh,	u��\�j	,,�~N�,|.��P�뱈��Vd�5.�s��ak6�G*WϿ}�1�ggp�䬷�J<��D]�I"Ȥ;��J['j�P�������Sr�(�d��U�}�5�;��9�Px{�YK�c:It���ܢ��	ٗ��~͑4I!��&X *�!�J�7�<�l[,�:���I����{�����~���8 ���#����<!-gBI��wD�du�%�/��xg���u �-��:|�٫���k7��A)�T�$��e�%%��no3�P^Uo��τ^B�u��#¹��4p�+a(�x��XI2H$o��T:�=GR�>�[[/P@%UB�$�N�}4i��$~igw�{j�c�kR}ڋu�-�B�g
$`b����F�(��ޣt 	��R\�b�(�̻�4mpER�����|��wqbޛ��	L�ȚT΀;��A$%.�y�J���Gʺj�H�gw�~����9�<����Aj ��1�Oo�7���[i��J��������������������r�kֳ��-`�h5{���ӯئtI�s�'KQk"��=DH?� a�C��Lx���c����~��y�Y�?J���[���p&QA /��5�|7ݚ7#j�K*��?C��('��y�֏?U3��d�5�x2� ���T�V;�v��}���hHc��	$�w[��S��c�^"�
"�����e���1�a�x[����$
�vI$_��$�}ޡ�1cT�ް�I<��/) �Y����<</��h�gw�w&r�D��Es#�O[5�I7-�yK�"v��Y9vHǺ��yd{NU�������-N�y�N	�P���q�m�ɋ�l��4L��t��!4b�~�V}����.�"4��S�BIS;�[��M(����_g���T,,�s5���R�e�$yL����H����i+oķ��7���s�!���5��ar@8H��Ĥ��O��l|<�I�m[�~~�����1@��o֟��澤}@~�|��T���gU��� �[[pxN�g��}���3�7��ុb�>^��xd9{�Go���^�|��������7I���3��C��?
�<g�E�A�3����9t]�����I���P��� س|_a��«��:2�U!i�v�5�*� 	cܠ	M���B�$�aއɫ��Ƭ0�I2UT�Fͺq��!:�%�����h�2M�a�nQ1 �d����Y���OhlgV�my�yM.��~��T��%�����+�Q�S�#���:��!��j	u�#PnGFL��\���n66�WcR�Mj��Ϟ���Sg���~���o�BI'�٠Y���.M��|�Y�=l�%ݏ2�$��:�
@m`#��)çE��ˌ��"s��{R&oMC`g&�e �I3�u
��Z�8�����9>	Lg���3
s�Ȳ	�<Qt�$�C&3��HM�߭k�]�@��ﭻ�L�H%�tp�D�Ib��{&<����I �}ˡT���!,�y��snU<'�.a���'�}��htI���2 �ד@�������v��P��]v��fR��yC�<^��4%aF�^�͒=�L����?r���}*��b�<���h�֮�];�����������>�3��@ǌ�� ` 	�ϒ�O����C��f����

!]�No� B%}h_l�	]������5���Y[�*�$���@y����Ews���u5	�y_��H%��������H���,b�]P��aCM��2m���� 8x���t��
��#c���M1�A �sba&I$��<��|ރQ�^d}��?��I�����I�����l��g�1l,�@������v�:�ح��l�\Ȓu��q��O,�d� ����%k;�Q;�y=�|�)��&�`"z���xz����s! 9�;�R��	W�lp}ǰ�]p/BD�[���E!/�ܨJL6��
�ڋ�w�b!;��J#:j��ڍ�'�-��K��1!���PI+khy���I�x�ٰ�O$�wO�ޢ{�_�>����䏡~~OA?z恧�Hh�����|�!j�^Y$�@��)�"��"�d�W��D;�ɷw���n�-ɀmЃO���T`N_�hY��u�:����й
�ǣ�7��#�#��X2~A�%���24	$f����t�,kc�/	���E�uκ�=~*��L�x��x�U������h�J�t!�����p�Q��ٖ	���ۮ�G]%.�@J�3YG&���Όc@��rͶ)�1�-ff�K�`�33rX�q6l]�](`j��m00eSV�hmioW���h@y�9	u2��&p�
i��Z9�ʥ�͙MU��Զ��&���4��ea�ݖ����@����,�l���G]P�͒�j"+B�	��[6�a�\g�|�?����
!{~d]o�:��	��A�H�ϛ�*���y{R�
�ze�:��7��C����]�E}���Xq�>멣D�޽��G�%�`d�N�ʀ�Z��Q�)S'�z�rf� �p����4k:Q�x1	���x{˞m@cĂZ ���D��%�A�^�P���M��y��X�
Hwu�B���w�3����BNc_va�.OG��K��;�VϚr�$�+��	3����^�I �Z���=>6]�SLBe�\�H�Z;=��wq�Bw�����7���RXw"Z;�kގ������^(��L�O{�(
E�-�y	>Wm�KFxq�	�¶�M��b�Q"����`�R̙)������ÚL���Xп}�>k~a�fR��n�>�:R�p�ȹ�5�gwd���.M���z��*�yH�II�z�U$:����� ��v���f`�+]�*0�������z�*8�Q��Ͽ��c��^�-]��6�y���gs �mڗuL0����Y>��A�
*�Mr���KZ�� o�u੏��UOO]^��ί�33W�S
��dY�/��&@HO��͹��.�sܤ캱ӎ1�Dz<�u4ƒ@�՝5	$m���]\,�8����ta�������՝8�A� 7���i'�h;�'Ӓ���z�f��
L�S��B��	&Ib�2���ws�~~%���z�I �l�����G]�w�xp.³7.d$�F��d�:���>�SZp�GT�&�Kd96��ϒ[�k(��*O��Ä�Aw&!���u�<V�a4P%qX$%�f�]M�Wg���߰��k�z�(���h���ؑ	�I��2��\���G�%��T���H/�����TO�q6�J��RfL�~4��O����M�-�yI�[���QIGR�}���1֝vMp���{��;� ��RZ�m+�}�*�$=��	�e]��A�'�Mп�-��F�M`�<��R֜~G�'�/�#�/�ʚ��v_c�A��(�{�����}Y�|�zv`<o�n�9DR��q���r�2�9�0qsR!Y��!3N�j�F�yU��w�=�ro��/�$<(]��T�{e'{<�����=(��`��R�x=^��{�qzɾ�?Z�{�`�{�C��v,�c��a��Ҵ|�=����}X���zh�������{'����f�8��/_{W?#}�,�xL�{÷��t�r����<��u^	�0P�B=�bb֡Ws�f�٩W�/a-(>T�{�ǡ˂G���4����7�!���c��y�OnC7wFq9%��q/m��ľ��q��g4gqgn6���w��vr/\r�j�v��zX��'v�}��6��Ľ�^-m! ���.�l1's�ۛ��d:��9���������M���ϸ����z�1xd�t�ҽ{<Mך��}O�<vf���p������!3g��4s2U�^���+۔jg���N�����������2k���0�5�v��׺��V��^�ޓ�3����ϯ���z[ZRS���ny�l�T}�齜���{�Ş�DL���j�䵆��������0�1sc��pgU����Vq���wU��m�3�#f��t2�ב��,�|E$�l,��$C��vj��D��%�"�Ũ���FOqUi�"�4�5A!���ѣn�a�i 5B�h�<�=��M��0���	R��W���:-��d��<��ϗ�ou� ��=ĥ��R�Ir�����J��ޗww��XA��&FW1�1��O����������������]q�]u�_�����~w���k���y
@�����/X���Afg�����`s���-�E�;��ߝ�޻�~>=>>>?��]u׎�뮺�����;��?=�XV�U�[g��r=�R�QQ�g�/�&���gE�*��Z�T{��I�����ֲ(���ɞ�n���דxJ�|ɯiUY]S�/z�W=꤮���N�I)����2G��U�QE<�Q��経�"k�Kk/���MTC���Kk\n93�tm˒TTyV�_7�}���$Y^a�B�g��u&�Oj��"l� �H���.��{�z�A.Η�^W�T32L�O�
 �*��D
g�D]I�y'���}B��!$��M�����mV�Su�,��K��QOQʏ(��Z��=�@����M�}Z��j���%®�p�қ��^T�B��PdY�]�G�/�<�h	�}<Pq�<x��'��}����ǉ_}.� ;�CDAd
�y�JO�A{]8�����Eť}7%`�]t��GjBI+5�0Xk:g@$�]��)$�}�3<=eyTԦC)����A �p$�w��"���e�X���ek;�c<���ޓ�Gs��Z��@�1y��h�L�U�Td��[��h �'N�|�IZi��v�u�9�v�\�FQMr�K���Z�j�7eE�� ��N��w]NϚ� �L��,H��H�>��{��lt�,D_\ �	9�&��1���{�K7F�||�w��4�@ l��Rd��h�	g�w�S��dѷK��x""���$�|Ϙ�%��_q�x��w>jعvQ��$�b��?;��(�G������vT��!�In����LE���J�nu�ڵ���>R6d[WN�������G=1~{�Ms�H��ד�b�fg�gZw����Kof��~�b����� gY�� cĳ����X30���'o�$����K�û�=��I }��H�V�ӾL{���g�/ٲ%���ɓm�.*�R��Ķ��K-�[L��L#3�+���Ȑ�7D#���8e%ux�3/�^��������>�޾���8����L���77��{+`��KO�̘<F����kڄ�:.��n�zdoz�qn�ɮʒZ�C��)�
�j�&%�7a
�z�n%޹ �Gd���1����ޢ�_p�=�|��L��>��#�.�?e�;��ƛ�F�.s���J���;����������4ĀH]�2@�KY���O�1!S���X�
�w|t� �R��-�3}2$�]=ˌ]��FeԷ����D�d�,c��O���ĥ��$�C짾11�w6%�����o��N��/pκ[K$C~|�ݻ_Bgo	�����4v�=�g�2�ڵIM�  ��ӌ3�H��c�5���u�AL�@`�$�+�������q�@�ǎ<zt��>�m-�V" ��\i���&�Kf��Ib���[�L ��bWl��v���&��7�h���ت�`�k�345�6l��:=l0�K�E ev�44&c���fn`�cik;l��v��ԖQ+(r��]Kb+Fڷd��g�l����7���� _֬����f9,&u��,lMmP}3Mm)	�y�<N�%�C�4R���bf�[�EYSqIBe-�SQ���O�M?���U|���������+;`H�H'��[̷ljoT*̷�BnTĶ^�W�jj˭q���xy���$ύF������Y��!�w_��y���f{��(�����N�Ӣ���{�2H";z �*��ܔwJ��;YC:�̉bI;�Z@����%��З��%�֏{�;�=�o��4�D�d�$��D�*V��y�9+�}2#^|�뺇$DD%Tc#fK[$_��A��HK��a�X�?f�1��J�[]�te�phy�(: ��L1
����˫x4h�28�ۙv�h���e
0v�=���"!���fAjb��gٓ$UoG1LsM�\m��2��@�d�,�l�G��D��"Exg�ɠH  �ʰ��.j��d>d[׳:��]��VI|z��H���tQ���k�A~�os�\xN�����_�n�����tܣ�߭}z�O&�!f&������|e|#f�Γ^�CX\Y�6��G��ZOt�t�gC�f��z���2��e�����Ǌ$�� ��w��')}�
���Ŕ������p"ctP{��"��xs�\��M�t��:"H �͑��ګ#d� �w@��%��%���	mۄ��'x�k�_���ln��L���p,X�! J%1_�p�J���k���������HR��$��@�.�)d2�j��[��8�1���F�=��4w���"E�tcA�L��"XȘ��GT\n;2�dH �r$���_t�P�CD��.�-I�����_���\E(gj<�c�Sk�2:��r��5A�<D��w���
x��L�X�ˉbA �[��d�v=���6�m�e�U]�c 3ă��ܞ"!<+��s �d�|�Ӫ5�˳D�J�\�$�F��j^��}�r&�`�nT�` Ⱥ���D]����ڗ?lIv(�6���������z?�s�8'l�y��j�&��d���Z���Yn�]�pwz����4[�Q���=���/@���׿]����/������I��"��S?��ْ$}�}��%����CØ��#�ן;F�m}mk�T��	��,e�,g{�t`^v�7sr$(;wT'p��;�P-��I,c��O���]�^�i�u��4	�J�%t��@CSC�]~-"U�1�fi簏����5�Ф���qo�>_!��ӊˣ�Wj�4��+��\0�̷$�����g6����|	��'�D���H~��$��;�����H�֑W�4�㓨rC�C�7�e�A�� ���0�"뾉iA&`�����n�VG�f*tIx�Nػn��B'�4�G�f��d�2�x��|��3L�p�I;�$�H1���0n[����������t7��v8}6ӽqC� H%��A ���#}<F���皜���y��2�� �O��N=GT��2�k=z�]ڑ��W[ys~�u;>
dN���ˑ/��"^S�ڼ�ew�yV����	~3�ӏI��
�P��~W������������r��H�q�2@$}�I�d��e^��3�$�&Le�H ���$����I�~�*C��am��V�˙�;��lui(��&���-c�*�F)��~�߻��m�w�������X�]�"L��]	��צ��d��- �Msxlx��Q�h��5�y������}�ѫc�p$��ĂX���<�o�ƶM\�g��R��$��;ȯ���.܉%�1d��;��+X���"#]��!u�ͱ@���"��_��S�		�[K{�6�v�ut�(����A~���I�L��M ��oI����+�Tn�Cc9>�Ͻ W��x<9���l*�ьKd�����^W��L]�*p1�C�L�b���P W�{:4Q��M8�~ן`w���(>8׬��r&i�4�}+�r-��9��bӟ��8��O�x��o��Db��M.�T1�ØAl��:�,��3��x�q�<x��Z @�Qx��������{k�a����CV�uM���X԰��:Q��s��	*k�c#�І�#�5�D�e�X�0��f�1
R:�h�j ���"��Q��L��+Zۡ��6c
4����`͒^J��h����0x�(�jkm�覹�kE�L�ל�ZBZD6�@��.��&�Ҫ�Fƥ�Ҵ���6�b@�4l]���a�[����u�BZ0������u����������~���ߗ-%�2��(��蒢=獄=bZ݊��	+�e��D7����A��w�l�FX�{��(�'sn��L2H~��1�̑ݎ�bCFA�x׍���i�t���i��m�2���  w��?�?�ܗ�����@o*M�M�gd�1$�FL�"jiy��*.���1��=���u���|���Ǌ�,Ƙ�͙Ơ��'����k�"��mn�i��6
0HO
E�{�H�d�VN���⎅��h�F��J+*D�z� 	$]�Ou	�a[E����1>���	�u�y��\�aI�i�i���ѳ.��*�i��N���1p��R�_�=d�1��<Dh�?���v�G��	 ��L�;Jܧ�v�f;2�dH$��ޙ�Jh�f��^"!���g�nd���=�������F��ݟbq!a��H�Z<�����h�7;�3���Sw��go��|�T;�z�;�=�+�y�^�(������Vx�ǂ�30f ���>$� �̎��O�2��F�����{�5�^����;��.�n�LL43�d��t�$�:���So5����L���i7�=AC�<:��z�]��=\/���oo@�o�8��� 	j� �d~�ck��JjlG��̜� q��In���2������e����n!Y�������2`���5_;�H�U��V���z�}�Bc3������% ��,�Y*ۓF"e�K)a���iu�6��(�������i.oߧ_��[PE2��@>wH�v�fH|م�@�Ƞ�u䴑#/��1� �DUjD��<�g������0�*��@ K-�H�����)�s�撷O��D$��F(V2ά�����E��$O��~<"��Ͱ�۾òA��;���w���o�P���oi���:w}��=�_y�w��HӸ�f���\b�3���1q�x���x�:|������n �8���~��G�7?7}1�1r�}�CbY�-��"'x����@��Nr�Xv>��IU�"Ib[7zW���;�T��x��؜�;AC�<:��z��X���r;�+ёF�T����ĂF7rɓ�[o9��ag�&�%I��RZ�;<�bK(���0\4v�
��i�[����~�x���ϣ�|wy�d�ScQɚ � ��L�o]\�w�N���5�$�zZm��>�a�D"v�\����@)��ob���$�d�%��<Ɔ���I�=�)�:�u^���FϺ?��3��`�e��	�����	�:$�
pi�Z��2�.�$^�� �s��A�{zTD$�#(y���n�f�$�TH ��fL�~����m�>������и��!�1{���M���v�o?��7�����ϗ���Ǽo�mG���r�!>�DT����?�f�-�`ߣ������*���8����M� �$�҇��]<�Đ	{Ι���8V�-vUt	)�W��D�{��{��Г�53C�	��P�hpRp��2WUB]WP����
�sU��j�i��������ɕr�.��~�g�z�R}���!	���I����
�i6���������:�%�����H���]�=ꌫy��m	������5)t�	�N��7)�����o~>���D"��ۉ%� ��R	5�?!���QuZ�ċ�ِ@L�,_{�����T(w���#�7ӑq*��ͷ�����`]�.�ؖ!�׀C�֯��J:�1ػ��d�I��D$�#<,���d� ��ĀU��x��ȟ� ���-(=vI�b�g��la����0��&;�:�2g����!����[L�Բ�0y�����p�˾><{��W��Y`zqX���V<�=MkF��Ͻy�O��7V�=���5A_���~<79������mGؗ�<���F�x qw��qK�\ְ���f����t���9���#f�y��f���g/&���?(|���T�����������)��p�zN�	��>k��ׇ{ݾS�^�z����_��[���5�f��B��spu���r�dW�!��?��l���'��_Z�b�n���z���峔�e �������{��	�<���V��7�7�BE�Ƌ����f���;�n���'��]7��#9�^��u�OQ����>xt�G�p$H}�J�^�O?v�����\��c���x��t��W�Z���s�$YM[�8q�ݼ���+�g�k�{������tgU������'��'�z�;˹͞����e´𻻎����{� w���l�a��y{;��Gnl|�|��ey�ZΔD�c��k�Od�nR�<4��Ox�z����q�K�O����IG�=���}�ִrHgY�	r��o���UX�<3%c:��P{��}���\�"m愺�^^	�xo��Dv�{�������cC.���xƯ7����Me��"��r�36�3���2l��E�=�s�����2E���Ń�\�$H�&�9	����u��܅��~�7�D�ѨOB��Û����A0p��q#�`0a`d/3R
+[g���h;>~>Di'M5��wd+J7�c�	�<�M(��KFT).Uı�0���|<�\b�ݺ���P���V��V�<M���ꒌ�5O-�5��$Y�m��Â�~��?3��6<��tE^I�23��z�G{y��4q2e�e�D=NN&H\38���������������}:뮼u�]u׷]g]u��{��#.⹘nX<t�/3�|��t�'H���˓��loO��������|||}>>?�N�뮽:뮺�u�u�_w������EZ���@QL����$<�z%�{y�4'�t��Q5"�L��c�a��h�Y9�Sؗ����^\���B<��������-J�3ޮt���2���QА��0�ȫ¨Br��{q�$�^�z��i�Rb�����9t#s����T�=�H�S���#�
t�\,���@dW��=-"�!���I�S-�v}c<�HTI<�z���&xʋ��F�&J"zT&N!�2��'���L��%]�$�΁j�z��]e�eg�Tz�N$�v�4P��'�^QsE�ϡa���--�Xy<����uH4r�<C�xU�DL�g��*	�����d\T|�n�+6����"ٜe�XD-ٹ�U�yՆc�Xͥ��μ�i�HIEm35[)R�KAs(tb9�(Mʗh�K��7l�]]�Z�Dsy�:�dl�`��`[���Z��3�|:�H-l2cc�8����N�G�\�b�4X6�b*��De
2����^ҽS.�;�8k+(4.��)C%����ZFd�B��3�5�͵̴ 1��ƴ9J\4�嶒͛��h��L�3X�H<bر�rfhbƵ�R�(h9b�B��Jbk��aƎfh4���<�.���A.%�2��&Ǝ��gT@�\�J�<ܰ M��M�2�� �Sh�T ���2�a� �v�T�f*�a��CsiMvq�r��۴�+X�eٰh��-y�6��`��e�M]A�;c*fd�rS;g%f�����ke���j��U%�L�J�_&i+Ĵ�Y���6����,v,\�2��K4e��-���F��M�њl]�t�.lH�EM�6Xb:=�S�եۚ(G73.X��D����فsͭ)�ȸ���,��(�b)fUt+6�X��W<l��(q0k�4�����[`��R��
H.�Kņ�)����b�4(5���(9rf�y�,7��GX���T�ZV���j6�R۲�%�GD�m�(����M��F��&{!1�i[�+I�K,��U]�)`�,6�I��a���4p�c������˃)Y�J)�5Ѧ6f�C]T�CWs*Z�1���������t���f������g,��,���%�ђ���H�[=�����m��=B�i,4x�0�՗#� ���Z�)���d�R
Q��/�u�-k��;k�Y�u��)`�c �ʭpf.�QY��P&1[]���Y]~�����q�$��㗻���~�~����W5f�n�ۇ�L�W��`3�H��6�Tյ�ѥ�,X���Xp���N�S,!�+گR����1٩fm�(�Ƅz�Lr��5.�r6�@�A�Xh1�ڌ�@��M��(�^*����t��6;Y���eZ8�b�q�k�X�Ms*�e�kr]%�i`��J6l¨@�L���-�X�7�s�(�h�`F	rӌQ��7g����E�D$�;���̒C��� �B����8s�wq��{ٖ$ߺD��	��`��������D�2q��٭��=�@ ���3���dH��Q#]�U&:�rX��2�[�K�'�a<wH�
bk.%�<�+y�}�����Ez�[�#�%���H$~2QI+�c���!��c?�L���w�� �_T�a,�|���[;�]�;�:�����/�?�p,��a6��ϞL��b�ݥ�:3�;C66�Y"X�[�!����2aE��R�ǖxࠓ�pOhL۩�h��3�)u��ʶ��]�c1��M�3F ��7t(�IFu�^nD�H6��2ɂ{�<ԠN��s��/X����GlEȒF6��׃��I�<?�zU��1(�c����p����z#nj���|���i���dҰ� ��,f6Nx�qJ*͸zc�C��8Gᙾ�-̙³ǎ<E�D)�ӗ_=~z���ܑ��"O2dy��E�Li� f���O���&g듍��m��S-���� �L�v�� 	.�ڽ�j�I�o��1,7�H)��9m��@�����O�i�^�ݙ���LB�7��K�tM �,���L�,<�t��ir��05�9��O��")�H�kgX�2:vdL���̡�	���,N2�݊`I&��Zs9���P��wp)%�YD9�LҖ1n&����\�7�&P��]R\v�Pp{�0��"�G0�GIo�'���Y#=[�Mc������0ϙ�
Q=��mAi���DBHB0#��ά�%����{hE�>�,I�����XK�o�rY�]|�z��3���O��Շ1��]���$��dfw�V`.��_��6Yl
gn�yb=4,^�RnrՉvE��:�ĖR}��>�ϤI�P�5>��x3$�e�'��K��*x�ǉI@4�@В�1 �9��>$f��AL����}��k���x�0��Wz�]�A��8�.�� I ���(	��;�}�\^�w\�d�UL��°������
.��� ������"�=$�C��%��CI�(�:;�H';e��2�4�<b��A+�f&�	`M*i���`l����6�Ҋf\�C,A�:�D!O�md�2ė�Ȓ��1#b:X��W[��z�[;2d��y N�C��х��"$Cx Oed�$��)Oe���?Li���ܼ�2D�����A��z�Wz�o7�밢!$!M�X�X��D�����z!B�%�|z2@$^��SC ��ӽMW���i�t�	<D�:=����J�V�Az��%� j=p$�ݽ )�+��s�>M����N��fz���+a�
����=�����$|���p���yǅP�,/R�����5>�p��`>u��ĥ'�x��% Ń��o���#��oB""<C�+�d�v�	�����׹Ͷ5{�N�!Q�"A$�n��2 ����ML�����̆�b���9��[k��Kі\0�bZJ�b�D�Qfv�߾yz���~�}R��+��w���FLM2D�۽a+S�N}ٰ�i�%��D�[¨/tD!O
�uD5�N��[�Qƺ/fc�$�>g�N���#_ e\b���ٍ�y�Nr6aC��'���n��	`X=y� H*�j�)�Uwe K3�<	n��:z]��
�A��
"F�@ᾬڱ��f��y y��;�5��� c?.�L�/]� <y�k�|��kC{ղ&YP����I���"|��d�6μƧ���3J������$��栀$�����{�s�
�i�}E�Ow�uD>y����A3��#����9���H�{<7�Yi/���Y����w���N0�y�A����Ә)62ѣq�j]2�N��y�Î{���q��P�R4 z����ݬb�����%�]0�t7e�XW C8z�b-�la�#ͪ��`���Y &�e&ޣ�T[�8�s���+`��I��E�K��X���0�-�Yu�Hd�VZ�Wh2K0�
�i]MLB��4��8KXٸ��a�s/2��1�` ƒ����u�D�逘X͋�t�tl��Z�4���f5CbPb�x���ڨ6&���`�&]���*ƷY�����3��~[�ʎ]����{|~u����y��H�ޙ�c�^�A܏H���'̙�ٓm�aƻ�!�C��b�t`(lb2|w����$cu�ͷ�$�} O��P}���UU���?�i#8t]��<���\�,H2�Z@,I����sSc�H0�w\��$�n��"w����"=�|׳�G�5V�5WzhH����dԆ�K�#�Θ����~��@��>�"F�<}�r$��^�H1��^��H���"P���˷�a���]j��/��d�w����L)<9G���G���l��䗚̄.�p�ق�u6c`*�F1����Q�#���v2K��d]�%���Tt�����kk���c�w�F��x�0�"��C�����*0��\d�{������~�]k=����r��pZ�Nd�<���;n�)�Y�s�s����4��Py��(����O���Bx�ǀ�	$�J����v�[�_�E���G�,A+��ă�����&�ݐ���bE@�NM-��ȇu���ȐH��$���x��y�և�=��>��H��̍ '����]���a����R)mty��^��L11�fE��M{,$��� Y�����PD��"kQ�b<C�<U�C	`m���o��
��#��2%���$I �)��L����=7�冦��9.�'p��!�p��$u]f����2�F��tk�l��7M����|�"
	�@�9Ւ�
͸�%���_z �	n*Μ��L`���%wt	><a�)�[���w��l�����J�I�H%��H�$�o@q���5q�bN7��?�<<Dx����t	8�.nn]SA��������,���p�i����r��Vn�VN}}�w��W�e��z��u�NF>U-��V��*(_��a��s�s���]��!:���H
��x�#,�P-B@$3�L|�&%vl����� �F��ؿ�HcH�U�/_�@�ߵ�%��zgG��6Ɓ �3���#1A��L�����>��>���eH-��ճ0��"{�����kI�x�x��7��2	�5�ٖL���d���V%Ƈ}��?ԖW����G�]���,�+�QŻ]�����j�%����׺}ݕ�{�͟M5 �d�3`H"���@��[�s��+k�vZA�w@�!�u����s6�q'�>t��y^�����1 ���2]�nvy��md�#wO`SU��A`K8藪�����6����0�D�{�2��;C;�U�H�@�yꪽ��h]��߮�5����4y�T��#�:^��x�
"Qw�ˬ�o�QĀ@w��ԁ ���)�}�]ٞ��۾��W��;x�0��yGh�+�)���	���;y��!�{� �s���}��-o}"_��./��k|0��D�Y��9[�y� ZC���nkg  ;;���@%R-D4	b4���@�|Ms����
ç�����J��{'dT�4���4�{�D�J��Lm�Hؽ�&��E�D:�B�spTHb$���&�tҳb.�
D��,cM*����.�?/����7R>�~��&[Y�^T���hel��$|���6����A�˖��x{a0��m=������������o��? A1�� k ��t�P���gu�y��eJ�&	Ɂ��I���I�,��Uڌ襾�O�4���Ī� �d7���^a:x�t�J�w�jc��I͎�D���Y4�g��k#-�:f�-���zD��B�D@Q�%�� �LY�;�D�H�x�J3�� �w2ĀK*͖��ޙb���I�d��a�f�q�����F�{ػ������G�ܘ7���'�z�Rw=���T��,�/|� (z�G�ޘ�M�n�u�K�"^���C˧D�<<WB��F]�>k-���[[m�ьO+ZK����I	�'}�;D8<x��5CD��"@Em�}������c�!ep����L��´Lҥv��E�,�̭#�jj�]u�	# �%�2�\�]�6��16����\�]��aγba��Ўap`�5ɰ��r�%	����,�۶����L�:(=N
,�	�Ks��5L� ��JM2atqƠ`Z^���uά!��Bh��Fqj�q3��_<<�[��ZT��اR�H���Ԕ�eseY���Dj�T�Q��\�wHC���7�S;R�(�X�nD�"�ze��WQ�hԝ74���H,Vn�*�t<'0�Q
m����[Y#(Ϧ9b���l���$1e��$	n�����;�gl�d6	��px�"".��}Ēs3�H�H�Uc/�+��7�g��$ą{r$�L�gt	����0�xD'&X�7sw��nn\Vb}��C�@ 	���� ��[Qۧ����en���������̈́S���`�K��]ֶ�'^vL��\���%��$L�w5
=�s%ܾG��q?�h���-�Lj���a[K�6"�[�eЅSX��[M�F�z����vYU�O�LF�5���K4wt�;/tN��n�k���� ���H�m�r�]�!b�1+�I��x�3�ߩ'=:G�r�tؖ��ݽq��gl6�8�yo��x�3���G��O3�}�*�=s�����<x�!� �����H�Y(K=z�Ƃ#�ߟ�i=�kH�O7�aOM�+�x2	w��xw�Q
Z�tù6��FKy�S$8ā���Oo�ɻ���sۑ&X�;�2i�V�aBO�D�{U�ך�$}�N�"1�w�25���Ynd�x�w���LOai�H�Z�����aG�ne5��%ߺ�����9�̗vL�r�dH,9��zD�*��iY��p��I�Y��Bd�ls��k��;k�!u���
O��ߘ�9G<��ɹ���+}�)��<F�7�#5�7F�Ƥ	�oH�xli��DB��l;X
3��Po��]�M�AY�$�%wt���^�}�OE�{y�Ek����s�h���$�\I'X�����,����kz� ���&Y��D�����^��Fy{t�{Bâ�{c��}�yzU���^��~xU�7'�7Y�/�<f��OU�xx�n6p��o^��pv%���`�}���y�B�~�y�/j;��`���?_?kl��n{.O{�bG�ӽ/��g�R�}���\@Ӫ��9�j�ic7��{�(zf8�_G^�5��U��������[�o���|��ym#��Q�b~7��ޢ��_-����})��MK�o^�Oh|>�zFp���y���>��;7p��甼��yd�7�r�IiO�/����<ޮgdj}��+���|d��r��g}�����ض�øc���;{V4���OjD��w=�x��Ϧ����wG����q�y��n���=O�[�gx#���MB�s�#���7;��P��'���R�s���I�s�	~�b�*�����7�eŞ��p�ǜB�|�z��w���;7�vwq�d{W}Wnb�7�������nG9!�o��{ݷ}��X{�0M��Z�f��ٯ�}��o����\z{l�p7���ej�uHI��:!��.�z?��ۃ��݌c����iz������=[p��0�����s�#,��3���y6��j_�w��<�����_���x��{���)�ʜɓ��M�$�j��{=��,黅�t�6�6�1gy�����G�W�
L���?<�=�����Nv��r�J�ڥ׋��xiJ�*��ߨ˜{{�t=/b�9\K��π��T��~�S��H*����I2Z%Wϱs�T�-1EB:P��������kkkikklnhmu�]zu�]u�뮸�O����x'�%ẍ.K�ܸ�mD��,��G�g=��91��]fc����x��}�>>>=�?�u�]zu�]u�뮸�O=QL���%�!P)R�
��
�C<��$}��~Hx��$���H�"\�̂�����9EG	6�"(�&zTRi��ܙ�Fn������A)��C��F�Վ��2�#��\'�=H��z���TE(Fy-�3!$���l5��J�3�M�^}J=��	Qjy��^_m��x�y���Ȋ�=��"="��/Ip�"��l0D�<��U0�WB��ʣ�(���ȧ.E^TY�9�������{m���/a%%�Td�<�&yy[�\5��/!�4�<z��L����/dʺ�S�R^���Ji3�G�L��=1^ЮnU]\�g��<��?��[����y;�����ĠJJRZ��Zj�ݹǫ�2�1!���Lx���!"�Z���|����Y$��L�d�/��$� �8��Չ)��ѼF�c"w.�D	�������C�3Ē��'o�H�Y�7>�I]� ;/wtX�b�����g� ���	[���^`�V(��ۦȒ�����u��^�ux�3-�}�}�4����מ�H%���}��,v��Q$ȩ�~Ȇ��s�?�J ����Ĳ�_��ͦ���E�X�@ ]�#X��5�!�/3l�&W���=�����H@�4uq��D
G���e����� v<y׶kMD!�5�1��i�wt�#�^r�]ˡ�'���}w�b�/@�";b4L�;���A֖\�5�wPv�i�G��E�����+){�߰v8ZCۊ�e�0�|}�	�o�&����+��?W��3������X�؎�Rc?�0�>�����M4�HI��X�,G�odL�i}��!"�x~��&�7�'i�w][Y`�bذ�w{fu�>d����E=����ߣ� �����׫���r���IP[�ٶ`WG%�K��[�m�[�Q�����>��ʎM�[2},)���~����5�Glhv�����Xd�͔ҡ�|�ɇ�Bp`E7d{�#��8�`z�٨� m�N������� ��'Izt�u�`����J �Ȟ�b|��$
bMt?�jȽ����Tp�	'׻%�"�-��I��֛
 �@x�R.�����F�ϋc皉bH#��"A-��,
�N�|n��{�[���/�ܺ�C��x��i$�)��LcϫS�;C�]D��7Y&��̂H����@8��$7A���b�Ta	�z���*(�{����ɸ}��\F�/�=9g�����5UKɦe}�6�����-u�nz|r��,�^��8�m��Z�ߢ#*��͚�����:K:?�%�$d(��~�{�lل�e���	��m;FZ�f֊7�'��y��,�.�n·]H�A�$�c�S)��m�H�1�i��[�fkb�쑺�l\��+8ݜB#�ݙ�`RV���J�L�G��,l�˶��iBQn�x.���p����H�[�i��ʹ5����&���%�l��p�Y�c��Q���1]F�[fv�h�ш�[a�-M4��]J8�9�شqDáQ8/�>��NbBED/��~�bI"�dN>���^ƾ�=�9�;dv�L�$c��2Z������@1]��n���U05� ��z��S$��a,I�72^.7$t�y��-����L<"��<=��+)��H6��$<�_#u�ܩm���Ir�	�zD�Q �Vp/m�]�螙�e�����N$�}�$@#{:K@;�.�����̟E�F �������&R��ؠ���t���:�߽BA]�M(�vt�,rnŮ��:�@�(:���r� e�m� ��4�4˞Єj�2�����1�Q]��qw.�#�\�d�%���2i�$��Ι>�V����ٴ��}-T����	&�w;���Q
���ne�iJ�������Ap)G��d�,�1�5z���y��� .��F��S��\�_Zg��Y_���/x���>��}{��w1[�t~���� px���j�bXĄ�cb�����g��m��<�;�ӹ=@����~d�Sm2�9�PɎ�la �Y�}�
O�if�	 ���M�-�a�\(M��Iy9���B$[��p/� O�
��,䑛�2�ئ>��*"�j�fc޷cD�j��Ʌ��%���7�'`fI�Ot��b���s�\��� �[�2	����᤾� �@���K����136!��D���Wm5\Z�a�j�f�aТ�����݉c�p�/z�I$�u�����io�w{{����Bl��j'�uùxp�C����x[��u睋$���5	p���,�eM4�	l�ݎ�A(�#�,��L�D�*/$4����ʤ�9|$_���:����g�ܭ�N�ϯ���[D�=�j��J���Ի�FD��s�M�Q�i����C\p��w�����|��?�	����<9S*TH ���� �f̚b���-�$�F�J�""��6*.�]-�5a�[;�q��� ?gC`[�#(eʄ��xݙ2	}�Y`��H@P#��]77Z�LtH6�1�^˻��]X���2�H>�K	5~��Z7ޯG �	%@�E��mZG:����[�CgeA�]6���!4b��~z��B%D�tN�v!�,�B��a ���5X��,��2�d#3�I�NC�
 DD/&%WE�H��zښ5~����$��h�|j��;�P'��SS$s3�=F�����L�'\�.���Q�<6�]����<Nl�EC��ؐ~�:������s
 �B�-w\���Ndc$��2�$���������I��;D�'Z�(ɫ�4�pz�ɔI��VJq8���{����!U{��=�^{:n}&��c�J��D]��y�8r??׷����8DRQ� ���br�M�
�BI��"!G��	�l�����q�r��%�?EL�J��v2#;zA����2Bn'���~��ĵ&H�U��%��QŌ��J-���;����(D��8�gn������Gc �d��A݉ ����J�ޯ	����.�&pj�^��ЉQ ċΚ�1���3ނ7ؚ���8Y{"I��������~�$e�>K`���:P� �B���lC�ٻa���u|��N�O�� ,��$��ޒ�S�Wr��(�z����Nf�;�>G�� ��,K���[1�ٳ�p15�gk��5swx�w0��	D)a�@�5��a7�-7q�����]^�Z��"I'6�SmA?wCI˽��/�V��$���q�(Y�v�MG�_��^�5�S�|qu��>�3����y띊v�;F��X�7�b��0T�}�1S������"���n}ۈ��r����Mz������C����G�Ĩ���(����7�V���U��6���ЉK%�r��t&�R�Q�2����T�a��k���fmE��Y`�9u�r5����h��VM��a.pи
�]�v��K�:� �K�^rqf:*6�\:4�g]� �`b拂�%�ť���13�j�(�cˣh�)��A�ak��6�̒�Ҩ�ahk�ˋ��Sj�R���Z���AtՁ�.�NcqZ��&!�l��˒�U2��R��Y�/��?�g��s�|s&�H$��ĒH%����{������D�d)�9��s�P�R�^Pv���r$�)��w�ۗ�	b{ݲ��t���b�naW[��|3<����y�D����
���2	U�n���l7z8��v�Ud�,czdN7�O´K-�[[��V���N#������	{�1�1`D>d�%gt�X:VL�����.%`����Q�=�/�� 
�Ȑ|�K���M?��Y=9���b;>�Рgo��*a9꣖�~|�鱼�@�3�z�,eU�-�HҒ��l�i�+r��=ድ91
J!H��ə$_�fq����D��Q%�g�V&�rf�>K�;�����̔�M����[	;ǭb}�u��: ����:y�.��ē�������q�a�&�=˱���b�Jv>Y.�K*�0�#�b-c�@�H�|�9��� ����|��Z�|���Rf��b�{»�1�7��>~簔BJ	xX�����HW�oq�8G�jɊ�MH�J�ٖ,�zZG��$�ЁQ �Tt��|KRY�ϟ �M�����$��d��Gn���FM{��XG��������DB�z���t�g	tlI�;�s�p^��A]�,X�n��s&�}pH\�[=�}�1 �] �@)��F[/7jR��ʛ��"l�
kV��m����|�G06_�S�t�Ib��$O6�<I|�@�߄Ǉ��m���wl�d����q
I���s,��V(�
g}�Q`H,@+2�I�)�w�[#y�Et��5�txI�b�'w�w���<�T4���K7��߼���Ȑ$w;�{K�nA������)J_=��.h���F���ϫ!�c*=e
�q��ɓ2d��/�>j�_���idIM-���y�(�:��IA/|���v�	��2��������ޙ$���o��9���ʢ`Y0�;�'�B	D��la$�(Έ�uݴ���J�t�5���H$����~y}����k�-�#lI���A��Wss4�p�ܤ3v̸
���M�A�a�{���n���Q��;�q ���%��Z���������I泛zexl9uਇzvؘd�}����Q��v7�����N5�dsPG�e1q2�Ɍ���ަ��S��h/� =����c)3�<,>�@�7&�h&dڵ�����D��̉0����!�	;�;����5 O�Ҕ{joA�]��QS�,H�A4z2e��!��"�yQ�HgUBؼ���>-l�.2���A�b�e�S}���v�p��u�靁槻{�hݝ�B�D̓���ə2d �	�����H�o�/!%��^ �x�Eĭgsq�D��ը�M�k�� ��Ȗ$��	-���"A�o���}�C���K�g�&��%a\jL���M�8��	�Y���X)�F��ަ{�}hA'�P�Ȝ�bKs�"H ��H�z_�xgc��bfChD�nL���[j�x���.�/1 1]dN_D�Nƾ��I�g�l�vHk$:zdH%�Ƚ���z��@4�N
���Ä���i��@)�D��"IY/0�ݙ�㬷�^�<�C�L�"� ��z�0$k]/������/�t��DO�Α =�� 홐�H�&}$Β�4Gt�o��P/^� �>�l�څ�����w���l�T�y6�����)�p1V>�]��iaL�\#�zdxo#���"�`�U�<erR�f�$M\9��j5c��]{6az�8�p��,�~M����\�yn{=Ӈk��[�PKǌ{͜�}{G�г�7M�\(_p �G.{ �km����$1@��L�J���uBWi��}t�ܜ�q���������Y���ѳ��ćom�S>�MΣ�I�>����	���=���C�ZI��\ܾR<&�مA���6B�So�=���L�x(p]������=i>�o��u��ұ����-�Vk�<I����K��a��֝������kY����7o=95
��$5q>���t��p=��*H����ؘ��떎���g���&*���Y��6썮�t�"9�g���vaQ��{�Ȋ�e�bq_��U����B��D^ b��|����y�;�C����2m�2�V��U=���:�4����:��y���>��^c�/nxo� '�/����z痳{�	��S^Y����=0/p}���k�K�ݝ�_�0�/,�%9�T�d~�e��q�<�5d��ٕ��Xq
�K�3l%�k�gx�{�'����OK�gU�'�]�aK7,��R�#s���i�p��bW��|�=����S��ǩ��I͇�TW�-�p
�E��'}�����+�E�B[8#���|Q�ˋH�=�Biز���e����̩��f�m�BȊ֧�Vj�J�X�Y��X ��Ww|��������ô��0�k�ץ��{��Oԫ_LWuN�=�|����O��,��<�s\q	V�f����m7� �),Y�N�>�N�ځ�%pD��%�8`)`-h@��M���cA�-&�	�� ��&�o�<�r����+i-�Kʂ�+�F&�f��W"���H&�@A��f=1�8��{~8�����������㮺뮾�u�^�u�^:��9�X�e=���RZ�夤n��W��VE/�ٺ��fq�N`�����0�����q����������~<u�]u�Ӯ��Ӯ���^�G3"���$�NQd&{�9��ocqk�Us��C�gnA(�'�D��P<��x�AyD��^QA�	^'�h��Mqb*Ua�e�e��Dk��\;XNQ�\$J�ʠ�2s<��/L�"C�>��L�*���!Q�xPQQ*�ji�`��$6�]wTy��.Y �)I&L�<:��FSc.g�a���5L>��O(�S!�e��Vi�^��B9.D&ff�Ρ^��Oef|wo;^�$�s2-*�Nq��xz(A�z)͔�oF�\���ߌ�����$5��.5�n�W�3=��Q�&GA�v������շ@ 2�aZ���0ё�Yo��^�Kc���] !4�j]��@�3tM����+�t,e�s3a.��J;X���i����`nt 2fL݌�*^H�%��V7aۮ!�#m�2E��[���!J`�u9��e2Cu��\���2�XM{.� �s�
BSXB�H�1���+i��	���˰;;Vli��f����'�Xh*@ķ�4"6�Xt��=ZL�z��>��rZ�ι!�kiu�L�nЦ1�14rRb�&��6LJ���h�t]I�Tխ�����*�l��c4͵��j"l��Hi�a��uښ�e��K��8a�����&�5ֺ�X˳��8��$�{[�I���[Q��Sm�а�YO�-�l/���Q�Zjh�d&�ء�i��nˑ�v�G��,�If��شX��4-V�9�a` �@΋��Vۜ�GE7X���۱��
-����tN��vx��,���b��f��˶%Rۣ� �f-!nT"BFV/9�a�Ü�T�Ka	Yq���)��:�n�k�ֆ��1�J���#uWB��4Z��c8ζ�M�K0bll��fk�kp)��C%���eb`�� m�X	b�;�\mi�m�`�U�f%�5]�Yc7bZ�0r��,������a�٠K�3��ˬ��faF��K�F<�J����w�-2l���n�J���&�M,^s�a�u=j:�V��庮�J�-,�ѣSv�%��3R٢��)��3��j��wWavB�GV$HEE�f.�GGv���D���6hJ�����vʔ�(��#!����6MD�.�,E@��Vr�����a����5�]pA��L�M�)e����k�`�bM6�ӕu�SB�dQ��2i��hLB�>�y޺�^�{�;�O?	��K��4����j��B���	���A&ir�����E����B��U� �(�͵�m�T�hשI��[a���̐@�4��4eZl�4��b��ݒ�6kH&���&��JQ��:WX��9ٛl��^_<� ,"�tΙ�k(r�R-�[lc,յَnaM�r*WS!q� �-'a.�q�w[��+b�[Tk�l[ڰ3��[j�=C����"�P�kǡ!�?��H �_D��"�*o�x
~�4�,S�䉖K[�{hA'�U��t�L��Ϊ���kw��u�>d��ВI�oL�@����|GM��zxI���P�C�D'������H����"�"���h|��1[`�Y���H��L�%��|: �xA(�z�~����a�^ډ�@�c�L� �_{���"�v�$
�I�Ι��X�L�)�������ޒl����_w\gT	Mm�PS޺]�����"4���a�@w�`�X�ғb�4@���\3KSL+B��/(XR�A�� �:<=��'wP���T�SPYy��1!2B=�2fg�~�S���s0,	�͐$q�}ED$�x<}��A��>
A'���w}6e���\�o�W�s�yz��Td^+���!Y5��A��V�<����媷�[K/���ɜ�`H[;� X�w��5k)$��@"Ư� �uQ�8(�SC�������Ђw���x�5Ū�#��Q���4�5���B�Oz�dI�;�d�P��(N��"���c�{:M��lSc
g@W�"Y$�t$G��A7�w�ʨ���v4���0$k��K���C���� �n�dӲ���bܿ��ے:w&X�I �m�����Vg���K��/�l��r�k�ÚFh] B�sz�J�d�Ѓ�3gH��;��㹇w�<>�ι�K���2Y�&�[V\�x{���D`�~��ɟ�?�)"�a;>���\ u�v���\z��蠙&%�������G>�c@�Y���땩����Gy�%�p]�z�񽛐$�-��IbA�d���]�0�
z������=�ρ�	����E���N%=�3�����g]�Z�Hu?�L��_eg���"q�	O��kld2o�1$���ă�BY羪�4�}B�m�{E?�N����eR�:��$�&H$����7v�Q���b�X9=Q8.:�"���	��Q�I>�ؑ�@sU��~��Hܾ�$�O{"A$����3=���a�aX��J^ai>��.�r9��[v��+Mkw1�cf��c�]c�5����=��4��w�8��"��ȐH'K8�ޠ�S�
r��얐I�ܑ�i����Z�	�C���[2".f�bbF{b�/���7�6�u�F�o)��
�އ聍s�A�1����% �h'2�Q��� �^t
$�Ѝ�X{|��d��tv�H�{r|	��{`���t�=@�Ȭ�f�L��Ͷa��P$�5���$�z;x�Ll���I]�hB�W[=��2��xp;���O�t��M��{��T��0o;��.���{2*�����;N�ѝ�����Vo�?W�Ӄ�8'�1L�椄2mY�2N|I>���S�B	�R3�n4�doG��q���� A�2����d�{����3��@!�BQ��~�z��5�[��Բ���L���1���[���0�?�߯���9�s�������=q�Θ�D�]=�L�%��n���ˡ@� ��[Z|*�D��#��l�o2|٨�/Lʕ�I����cH$w�fKGl�F���������B��z�=��k�:q
xy����$	載�Bgb�(�|�F�yS�,hu�̃���ȟ8$ȡ�6w/^=l{"�����ܥ{��
&j��:d�'_z]���މ�K���%��L�����
Q	;�O�<s"�Iid��wBb��_��^vmz"d��-D�ӽ2
��n��ݎ�����J��N�܊c1�'�8z��K?�����|цD�ix�~T_{כC�"��B2�Igg�,�䅗�5�$�V}��G�	�7\ߖd�0(`��<���y�o�^/^<�����߃�����ǀr!��=v���κ��
%��nfbD�ƄIv��L�� �[`���"�6(�F���/q@Ý+��b�j�鄰Z�óWYV�.&��j�9�$6��v��RRR+r����&B^m��+.�9ͼ
����͙��R�UE�ڙ-�W,[r���[V���ˎ��9�u.565)�(�K�A%5��@�����Mpaꩠ�N܁%n�Z��ɐ�ͳ5��HM�����e����~5�mH�7�$�d����#Z�ףo
1�
{�흔Ҁ.�9�$�I��x
!C�'���/���&X��m�.�;3�y�l@�M��N$K���i`��좺9Ҿ�S[��j��@p��#�4N��M)��1�Đ*65�׎������8	8��jݩ�!׺�n	&G�{]�ӈpS�ݱe�qw��|z;��\�J�%��rA�ފڞ��d�� k)��q(t$��9x�>Ȩ�,� A�Ή`�#���S�0`���%�Y�"A �F�t�%������%�;��=�tAK�C��k3�:�M���T#\4�X˨gB(�B
i�v@L5���z��}}
�ط3��>������n$�ogL��{&}y2�>���ĭΒ�G2���zhA'�T����%��3�����Q
+�3������W��x���%}��
>�����ꯔ��h�-���v�����M����U�"r7-QH�E�PY��}�!���ǏR�Swׯ_��#;�Y3�7�gӬG]۸~뮞l���$�A��ݑ<(x���3�L	`Hf�H&�#٪E�֪�Ͳ+��& Nnt��='���vx&!ި~�
�xWJ��K�6%0KY �$_n̒EGs����6囓V�C�����u���y7)�L�!�O"�mƒ	˧6��)Q���{`@ӬG�����d�d{�d��]�}���f,��I���l��2 ېy�	m���Cv4v�mu#M�Q�Q�X��<�����p�
�H�y��v�E1��2c�*�湫{�+3 Ky�m��w.�����u�u댸�=z!�d��,X_{�A=^��5�X��^�!�	^�螙$	{Α#��=��O��*?���oH�[��4L�?k���띖/pd�͞=����*p,4г�jk^@py���su��}F����2}wY��!�ǜ�$�>�ߧ�,�f@�I/�t�ގ�� �<Bxx���{F�/A�F�:$�X���2���2iT��W8�� ~��-�����p��LC��	��Yn�H9F�[�FY�3�hA%�6ZA ���'�Gu߼��|#����E���r�N�s��E�8 K���G��k9&3R�Ilv6\i�k]X��|��B�)A.��˺�X�d���$�$��$�15��nI%��2]�H�	8O�xc�I�|T��^|��Op ��$��3$M�h���a���O�Z��HK P�n�%� �P		�%�B^a$�����$s\^a1Ò��<!����b*�bI>e���Syԫ�S�{� �{ޑ,�H�d��cvʸ"J �v��n{*�nr}�M̑��H������G������4�����齋qK�B�@>�=�lWo�M��A��7q(�6m�g覵�ۋ����~儡��;C�އF[��]1߳p<@�<���9��-�G-�g�~���#�FZRS�S]��yd��!F���u���]���g��~�#�d��-d��M�����bIc�IwlI��ʎ���,dǣ�Y �32D�]�˻�(;K�z��c�Y���Vj��L�f\T�\P��+q	���d0 2��3�kf`4uv)��׻�?��0LC�����2A'.$�@n�@�YV���zvd6��$�^:@J	w�M�?uȒ<���y��y6;��Kč|�	�ݽ2B���z�w�����<;C�.��/���
d�͉ y"(Q��ǾQ��DOk
�~�i����i7Aӂ�|w���a�wx4lMw��#Mzf/q��Ln��$��r$�K�j��H��[bWuC�}N:�|�TA*G�6kdI �wC����ϵ���uȒ�p3�ܑ ���5Ww��}�R�\xzz��e��j*K�*h޹��tv����`��S�Q��q �������s��{멺9AD<Fh��%�~�x�6��c�H���M
3���������y_7M^%��s���qć����>�V�Z�GM�z�,n��Ĳ���X+�&�۱�\Me.FbQ��^�Yl�Lƥ�YK��D.\1Ȩݦ�İipjZ,rT��c�#HkYl.�1��du�tQ����t3��!d�a��(��%��ap霴4N��3i�����Z�]7S	���� �17aVk)\�m� �Ĕ��	`Ɩ+�1�v�@��tЏb� �f7 �5D6�QZA���n��E�!����p3=�,I�I{�1LhDv̞�h��/G����$�����X�L��~��s�NUq{�mE1�!vfL�@ ��̂l�����F��X�M"t�
xE��:�[&.�;v��]�����*LE�Х[�[:�D� �v�Jd�dH�t8O�]������w���r}�H��-�; 1��	a�}!eDӜ�2��@�z$�l��0<K���񻉙YrH0%��G�����붠��:d�d��7�O1@���$Q�[q��w��}\p|��5ǜZ�sJ2�i�,�tsct����3JWw����g1�ܠTA+�"rZX��D�d� toH�PG�.�����U��݊W7�p���Q�H�3=�4�O_�1���ѫ���c9Z���7���Ӟ/�_��ő�]�ù�E�j��;����\�w��X<B��V����UWY��%&�Z��2d�2dɎ�JTL$�ݹ�F���{����6�=qz�%�3��p��LC���^7��J>�ȐK�x�sDO�����)���1�0�I�����(xv�(�'x���k�uz���`��O�`"A �u�$H'R��k������ݕ��cݵ�B�v�C��p�9x���TH	o:$�LX��6X'{6d&H���$�;��'�;~�ǝb�D�O����DZh�F%����!t��`.^��U��h̿~�ϓ �wx��8|���X���I�{�S����v�,	 z3$H�� ��x�xI�	I���4}1��דM��M!@�ޖēݽ-���Wo���>EU5,��|��DD<#�f:$�	>��Av)����|�'��H�t��rn+(��w���dX��>�I�v{c=^��NO�ui� �Z��q츾���m��@U�IAҷm�M�z���@#������狍���-���X|}ܰ_1;ܫ�Ł�=��W�n�Z�m^��"_2�ڰc�p��o&���V�}<�@�5,I���s�����r��<��b.:b�4�����œ/=�������T�Vgq�����-O�oA��x�3��tw{��e�=�|E=�ޘn�w�>��	k*��ݓ�g}.�-�r0<�&^�n�rr�׻G�y�n�:�_!Y�9��	_��}�ؒ4�<�����	�Fo]�Ӿ9��������9�O&��?�_ڂ�w�*/�9|�#�O>����q�KЫc�m|��Ow� ����;�y�����x/"�<c`H���z��]Ýw�C����Ҭ{�Nl�7�/MÜ6�+�M�;w�(�޸�׌�FOS�=��"��i#�)u��ݿ�l<�o��!�4H4U� �;.���Oo��$�V���ʧ�<k��� ��X������'��1YKA�ږ;���]�X��/��@h1�ߐ+pM�f�ƕ�����S������gf�%�p Q8;W�s&��.Y��}@x����<���<׾���Bd���������.�v�%�_q�����F�q:���ܹKc(  �����$�����W�h.R���������aE��G�{B@I��>z@��NO�6���%>�����m�_������e|���������9��������c:?��g�g����|_)��o�����\��� �H(?0��{5nG��y�L�����J噆Vd�����������������q�]u�]{u�^:뮼u���=���0̤���\����&h�E�4T��,x���~3�����������κ뮺�ۮ���]uק׫=ggrr�������	$�=�Qs��� ��:b�.6���}��tHE
��sʧ8��I�_����<>�;���L�����,�	GQMί\^���	�l�P]M<5Wy��*Ԣ$���OO4����5�=i�B�&z�Z(W�8yyI��+���²SK0H�"�ȧ�;�E$#m�eVF��W��q�#>M�ԩψ)�H|�)��g=���R�����t�"�z)��PO4�����x��aa_�c���92����lbZ���r*�2r�0]{������?ze���dI)���2KcO��}.䇀b��tt���7Y�0�(�1�u�'�:$�_�M�w�����b{��i�E
7^��EP9�SӕD�JFu�uS�>�����y_L�b@ �^M�"�閔�vʟIFwr]ˎї`�B���Ұ&R8av�K�l���ݸ`�3��({��DO��EF� �%ٽX�wL�QQ�[9���|�1R�Ķ{̱#�Ò��(P�㪤���k&y%�;b���d �E{6dL AGv�	c��@Y1j|,�<�&���	 ��.Z�y�I%�:$���]�g����?��b��]2	ۙJ���M�k�""!���[�te	��2m�F�`H$�e�� -��!��N;Џ{�-�=��J�=JD	�-�g]R9ǡe���} ��(��?�[����EQ}Q>p�_���7�����nFY��f��l�&M,�Hus$�h��@!���zfؒI�ˉ1X(�v���,P���%���̩�� ��Y�7�����g�f�!��Zmkcƒ�C��-�C�$s-�F�c�*�=�S���M��<����<@�d��lI �t�b�î����ݹ��^m�?g�A$���j�R�!΂�"'�x��Cmog��f���x�gg��i�@)���&Y�_�4�T3���Z��;��a�wxL|d��'��	,�k�������;[/2dOWL���F�t�%�I Ջ�k�BO��Κ�ѫ7".��@�ۖ�̑,�H� ;&�{:\zw��Y�bR�"m�D�UF�Km���HL��5d�=A�2A#����v7`N2@��J��D2�`�y�P"�|Oi��F\�B���G���+���δg/������{���w!Jc�.iZ�y#��<�n^s;�Cs���An,@���O�?<���g����Q 4��r�.�]>���q8�d����:.�m��j\�! �H�v��HU�5ٚ`
Ub�P�Ɉ�LR��,���@�%�b��#��/ ��+V�-�й���b9]16�"��hL��SE�b,��l5�f\1��u�ڶ�Ι��nc�R��9--�↰�cD��vQ�2ۡ���Zwk,Q5��I�ut̴�H84m�v-�x��m!��K�L�D8ɭJ��m.�h�4��nc@�2�5b����џ��<��b�y2I2�sD�E�]���,�\ǵY��60�톚~�]�kP�������ཷ0d�g����A�=�t@��\{(I,N����$�K��Y{�;2U�ylؘ;C��DOGn*$��Ή�I�\��{�����&4��$�$Bn�ya#�Ò��+�ț���I޽�J��H'=y-'������wDR:�4h7ޏ1�K+�	�$�;��s��@}݉ɒ�эv5��s�wM�Ǚ^g���20�Vόz��&r��/��j}xRI�@�+!��1���(y5�,�j��34�ݘ�X�p�mi4.���`�?}���w���b>πR�$���$m���̵#��ȗ�r�}>���,�ِLxM�Ԡ �Bz��l�3�9��<�������=���8	(���[��YNí{ԁ�d���6���t��f��w3��FD^�� &�A�&P����3�� �I�톐SYu��܊��ܚD�a�0\<w���3���HtfK$���=���>~�M�� �ِTv��M�ϡ8��	���*T՝�w��︁ ���b7	cs��2Ac;�":<�P��o�y�I�Ɵ`=w�?�X�%@.����x���$�*�4{�ZzB�0��}y� ��p��\�b���$"*ܩ��ξ��V�ޥ��m�`�L�R�4)`gBWV6ۣE����qeh�"���;���lN��$	�jbd��3�<������M�� �d2{�H�72%2���͈!<D<�k
f.%��=�q��&�޷��&�d�d�#���#)FI���{���x9���1	�%� sg��11 X����0�c�.�F���>̋���>�{'�����ǒ۞4ٜF? �{*P�zs�b�J�9$E�=�O �jhd2j׹��S{���7�I)�@�\u���$]��ɬ���T�&� �TOH��,܁ �@$��2}n#S߳4�������V6�)�_(�  y�%^x�""�z�칖!z��_Fj�wV;�y�9;��w9� �+WM�̱6i�In����H�ںd����g�>{�>H�T��86��I ��	��}#�d�5{wW�]��f�P �C�l��6��^N�9J��蛙.���/qw��������I�d���$�l�v���D��e^˗��>�=@�7�;�<DD"����l�ɕ�LK@!��h��l��1�}:MB��	c̘odHƟ	��9uD'�/�t�F�{}�Lu�O�0I��X�{��rhq���3��1f�4���>�|�tO���W���5s�W�sU]���T��&uS�?l��{&NzX�������.0K����2d�o�!�&D� H�������*���Kk�C��S1��.;��z�e�7��؊jhg�ʊH w��g�5��-�3�%�:I=�	�ɇ%v�h�sey9��iR��l�2�l������~���Es	�h�>�$�A�ކ�{������X�a�J���P:R'�rdǉ����xY퉖�7���k��vA�^t�G��e��ڼU\)&:���l����r��x� )�˘�ly�1F�������i&��d�6��CC���b.���=�:i U�X�TMy�OWL���H�NVp�Wg�IM3��9�]@Q	�\����jB� St�MM��e�m�,LZ�鍙�"}9���%�:�I|�=��{j�A�%+�~�OK��m\o�^�}�yQ�<�Dyֱ;�>�f��3ӡgt��^������c'J.Q�|��B������J�@��s�'�ď�k����1& �f��Poe���;����������Xf�t�֘�΃j�*a6�J奔[�m�AunE��F�W�aR�7X���MF2%�ݬc5T�،X:��j���fX��фh�W�b��� �Wve�l�A�4!���j��)bnm.ΉX*��a��e�����\5�4��� �YEu4�s��ء��lԪ�PI�6�$Ki�+��L�K\Q �sM���.�� �B�b��%��e�f{���ߵu[��#y���u��zwu�P%?�[������^��$K/Ne	��i�D�����H!6@ǋs�z�Z��I$�#c:@�,�'czD�dz�cq��\V쵲M��{N��T��<ݯ�ڐ	� \�ı,y�S����;h��̖����#u�0 ����5ԯ'�������k2�geg͐�%���÷:2*2<��S���'��v���cE�z��Dc����+�ܧ�{
�d�i��$�%��5��
��,_=�~� ��=�R�UZ�?�iHD���hD��U�]���ԅ3�冷0L7-*�~O��>���O�p.��$�|��,F�t�̐^zwOWy�@ν�$�?t�ȑ�a�����)�o��$-��ه�\�R����Ջ!µ���7�^���ǗuY�I}�9�X��)_#K���WS��SO�կPv�H:̙L�C�:X�d	${s�L�,���Y�z\��giL� ���<	DH�O1d�e���)�1�XF�r '3o��-,�l�H�X�wo�I	�8"	P���`����BP���̑�tď �s��3��
;_E��E'����ikԼ�Rq��oJ��H'�f�T�wj���g����|�2׽ S��X1C|o"_e����>�A' ��rD�Yl�L��"ZnG\�4nX��ZA�����E����7������H1� ���C��O�2�l����nym�U"X�j��$E6:)8NT�wܛj^d����:_��]{r$�L��ι��H�Kg�X	m��wL-�y׽@/}�PJ���]�S~���$@ ����� ������[w�?��{B��slY�{��\*�50�׹A��:�����{��_�S�-����=!�<}u\����n*�o?�����6�Kv_D�$tv��UG�Bp�`%^���bҴ扟mm1'��<h��L�ٱ�d<�s�C'���ܜwª�S=ϦK� Нb ��xn��N������D��<�d��')��ckt��IToC��r;�I�,��Gy���}f�m�t����SL ��*���YY��+L�JU�En�!Ŋ�<�@r����=�L�1A#�zD��*Ew)�":�E2��;HS<�i~�1H�v-�y����3����!�%�wd	�g��O"A�^���]QO���sO���9�]@Q	��39�${�bH�ePyi��2��Q�o9@� �O�3lP%���H&`����<ER�l����O��	>~���d�웖�{�!p�8�B����
s�\;X괾�N(3��gU���0g�m�>���PG��?�)�F/�~ [��7w� �r���l��L�>�Ődɐ	`b6fy�-T99	�@��G�+��t����>Y�67�}�q�}� H$�-Lk{�]�'�2�z��W�d��@����CY�p۪�MS�L29�`l�k��-\ݒ�X�Fe�={���K��g�����d��6$�ov��{�����5�v�p=Gl����6n-cr��P�s��GT�,�=h�뇜T�׿`�#� �i.�#{�dc  ��������zw�O	 �=[�/���"B����D��fĒX)��S��i�0��7"I';�d�&ÞP��#��`S��s�_*�<b�A���;;c�A��ZN̂mxC�ɐ����xp�@t�z�5�bO>d�6�{+��1���Ȑ@�&D,���,v;&]���3������wS���Q*�.��y�o�Ŕ���/�����,�k���{O7� Ŭ/'�w���<w��S�'�gq7�������c!o�x<���26؞1��9x�/q�z��Y�Fi����)����YK��Wf���}	5�38�f���Ͱ�>Y���D�۹����=���M��s�h������ճo���of�@�;�j8V��i��*>� ��yW��9 �v�:o*����w�yx��}5� �5�.�]����)�rv�{�����Ѽ��7���E��M�9<3�./ol�7�^E�u�Ի�<�e��] ���Ԅ���R�c]���G\���+��O':o�ʹ�M�7��ǝ�i���?{5�N 4ݚ��n��{����tn���g�x6�����9�ٞz�&�;4b3���JxTNs�g�5s|�O|�o� 4c��}�G��0�f`;�u_yfYȇ˽���Z�^�}��m�;ޞ���(���G��2(��1]���{��L�����ެ�p{z���zp\C�W�ɷ��U�o6dwuY�t���'K�P���SV&����hw@k��o��SKۜG]��/<�t�g���WB΃ϻ�٩�hZC�@�E��p�
��sHz<=�i|o�5��JЧ�L�`��x�w��Y�{�{Q��ana:�m�K��?��[Pi�ɛ���"0﵌y(�%h���sv8'�<�p��B�,J�eK�o�~�$|bǈxϝ�"~�#XJ�ޔ�{����'P��>/�5D� z/�q}�<Vi�u֦��8�8pFYB_hŚ�#���,���j��e�``���`�l	|2���	)V1)"x̥�z$���#�����J�H�Y���H��h�Is'ͅ\D�Qd��[�W��ߵ�lIQst��E��5���-B:���]���~���������������κ뮺�ۮ���]uק�܎��3
�'#,�c���Y��$�!&rNU#G8f==���o���������:뮺뮾�u�]u�^�OvEe�U�̊�j%��+�!Q=.�/H�i��{U��I⅔u*�ml(*��]B��6�!L��6����,�����덮3�w9�v�2Bj\ۨY	V��3�5
��σ������g(���9��l�Tؙ3���������۫&�ܲ�N��ԙ��l��n�==Q�g2lO�]��I���E�RU�3�&�L�L��Ԑ�z�mUG��T���x,a�*��Q�Eکk��dK�����c�M�{m���j��vB^"\�[`46u�@lF���9��s8XiMk-&1B��%�YM��J���ˍ5^�{�U�����,�c��L��.�����B�T�c`�M�YA�\n:0H+E�LE�������[,2z<#ɪǌ�����[XFք6�Q�]2�2�GDk[�R�Y-�5���:�4!���Yv\�HB���8�k�b��a\few]n`�,aF9֐�ƶj���F��Q̹�+��K�����M�7!t�XRĬ�*3kl&���9�W[6�V�1�k�������驕3��n5j�c�����옶+q�R(�kŢ�ҷ�K��\Z�M��mtA�6�V.�,^��!6t�Ѣ�+�L�3S��Q*�7�^X�qj֥ly��Y
�;F�m�GdN���B�Ii��$��*)� ����Z`r�a��T0��M]s���-�M��AE�*�S#)kSbjX�tًE�kvřfq1�bʔo�:Ơל�
Fb��9��ଦ�\u�����s*V�jj���lҘVL��f9#4Ke�ΣYZc�D 0�fͻ13��CW&�e�V��B[��J�jf1����#uk(K��<�K]r�$���Rذ��:Tv��B]���Lbl�kfҔ��t�4v���s	�������e����X�H#�k�V��U�j�)e��lC1��[H�78��2�1��:�6v��2���d{1!�U�(�k�m��!����`QBtji���BfʆՄA�4v,׬��Ns��b$1Fٺ��k[h���j�:u��c����3��5W5�sV�ښ:h〖�M��M>N�޸�q��= �R��G2��JXJ�M��$�oh
�i��tf6&�l����z��F3����L����8à8�ݕ�;�=r[�cj�n�R����]�X�ԌhQ�����+`�3�d��4�/2�)vѶ˚��)K f���)c����m�%D�غ��q��kb�e��72�M��Չ�[��`c
�RTh`M���s2R��[`m����a�W0���>���Q(��yQ$��݉��n������=쩊�܍Kv�OH�=��4.�0�p]<
a@��L�e�6�7MB�����H$��D�$?d	7}�W~�x�D��n�i��"���<66�m�'�v�#�~.z^��1�s1���5��pe�~�A�g���ks-�cݿ�;�+�y<��KoyAގ��p�f�x���by��V8�˨F!<��@x�'�P9�1 �|(�q���@DWt�$���̂!�힚b^�(c����~|����~�_%Yh�eR=��ɒ�D����)-% �%�M\�.����
��������8���;�{fIc�L�H$n�H�����?lk�/��!$'�zdϨuРD	DUg�<I'd�[�&.�����*���s�vj�wF=�H7rB��������"7ʗ103�1l�[D����R�m7a{�����"�����>_C Ɏ��q$�o�,$��ޑ$�s{9%�����B��"����Od ���Ic-���#<��#�#�Ł<��e��%���6���`<�G<Oq]�Z9��eN )���H�6���L��Z7��V� H��B�~��	�(�&v�"vl��3j]_��zn�ؑL��f�K6�ٓ�^��I$���W�75SC�$�)te�z�2�l,4�3.������.������$�~����eG>^3���i�(���̢I��฀��'�{�2ă�"�`��1��vP�A���/s��G� i
&�5m��yK�?�o��x� ��p�s wݱ,H$��pY��SS"h��W�����79�!��g{�h�����ߞ=����v��p������f�Ń�g�83�Y�4�v; I��]�1@���s8.��[�5x�.���N� <�jbG2L	��Ϛ� ���<���8���d�}�i.2�'�Jw0����~�i�Y- �wH�y�.:%�$����οq���9%(��ҧf���3o*��!uu)��m d�j4��� �}v3b"�Q� vg"X�I�gD���N	
:fA�WW���1�OC;��ْc�09�K���O�mB��~�|�e�tI$�e^́M�c-��Ƶ��u�s� �׸h'�RN����#�^�̒!�=��I����vj�s=�Z%��jJ~ٔ���<�%(�Ƶў�w�ب��j�� �$��D�H$n�H~y{��5�<����g���6/�A����(~������;�s�;��_�'x���Խ<��v睴���ov���gRN,CM���t�&�>��H<+i�����0`��@^���A���x�����K%�Y`M�="X�ǥ�!B��O��ܺr⪖'��#Wh@�U��BR�؆�G�b��D�u���+����z����{���� M�l��(����G_0֦n0�A�͙�P�^�4<D'0���OD�VFaP�*^�@�UMN1k蹙b��GH�� ��G�#��z+m��i�<�%��<�X�싁6�1GL<Þ��d[�ȐX���H'�<U�N�x$��H�����fn�>�l�Lm� �%���9��q�j��*��wH��[�x�C�x�R������o�/Wf ��7��ȶ5읖��[[�l��\���a�9U�U._��`�.��{�^�c���/Kg��{�W��xWv�4��T�pǑ�p��� ���*����bӄ,|���͏<et��0q{�|��Y�O� �%�0��h�r���E.4�k4�v���Ʒ�3�\ Jk��%���%�2�tR�1XF�V��<��J���;�Ytv+��V�z�;�vJ���&Z�����l�)B˫x[b��F�Ҝ��;knCL�H�]�ܷS%%�P@��ZʛMC8��3�n�5�Խ�J�a�e����u5�jg�Y�tè�M�#M�B��0� �c�4�ZL�M8��8s�"�����=qP$0�I�v̗��+j浏�-<�d�s+`I/�n��<S���-����H0ﾋ��|����A�R����y�AG��"#�v}�sL�ޭ�x""�Q"���I۱!2LO�U�j�Vg"}���s�$�,�-��	�DXs���
՗~݌]:���4Aa�#o�`I,Kgf̒]ٴ��n�x	��	+� �]�*�V̶�H�vD���6�UO���T���Ku�� I������Oϟ�-������VVl���)�RSR��X�M ���0�u�4%Ɗ+�6�jB��/�^����J#�/Lq�gN�}�D2^��M,�Č��W�F\��a�6��R�i��<)z��(�k�{�)�Q4<7i�wQ���U�U(�p�>��)��&O��ߑ���w~~��~;�v��^��}�}x�ԫn���OTp��<NM���Kō�}H$�nd����- �)�"���ޠ����d���X�<S���=��	8��i$�7j�����| M�t� ��Gm	<�r-i�	�(�����z&'/_��y�K�5�0�NDtJd#�zC�{ ��3���$q�[�Dt��7ă\+��P�N^�~�i'�=ę���u�=�M�l�l�W:Ԉ$��̂q��KO7r�c��>rFU���S�R[y��ĨS9V%��,��
7L�,Ҍ�]+�h|��Y�_|:������<��H$�!ѽBOz�tw�s"�U\̒�˙)����x�Q�������y�o���������)�����vHdwH�m�NƔ�E�9dԻ٬w	�����$�</P6{g�"i��ı�;��Hf8���>��~���ow�{�g;�w����l85��p�Z�g->�>�Sww�!Z��{��oV��=Iח�*�X�NQ��'�y�b�K����1��Kd�9$�3�w�K��#0\�Ll�S��sև${���X�r/ cd���7������2�}3'�X���������zg���{b��e����+Q�edP#Y 	�fH�I-ݹ2������0b8ߺb%Iww�Bڰ�\�!6-���a��.\�6\�����f�b���Ψp^'/m��Ol� �&Y�$�X�;��mK�����d�,�޸Hj}�ċ�A�҆�a�.�}���\)�Fh��˟I���%�,�K&;:��%���a;���$�A:r�F���y[��'�X�~w���vVM�I�gD�M���cË�e^X$�~�jd�t�[R _���O	(!��9�ב~D���/�G���KooH�N�u�z����9脖�!��c]�ۙV�n�����b_�kZ�"�����������g�	�2�UG�9KZ����<o�l��˙���b�X$go�I!�F][�x����{ѤL�=�8���S�w<ۥ��c����/ݲ�=1�>����,���_r��O&�)(ٳ��k1[�&�Wa(�<0b��>|���x�t�H�b6�݁.�˻dUd'�����	hd��ɐ	�\���w^o&%�c	ǻҟL<��tE�I$W�$H%��Gv̂a�bt@v%��Q� �ț(`\	�����w�2u��}�&CN��1�X��'F]�$�2ݱ^i�rE���"�G��^�y�<|�0v�d��ĂAC��H<���^F�b�E��;71$�bI�{K��B����<�O42��S��*�/y���[r5��햐A,��-L�o���.%_�Y��<j�����[��	�c�3'{���B&��q�$�r{fk���������Z�ف�y��A�;������\S������a���5�����u�?,��?�d.1�uH��p�����A��U����[e.�������4���Ҹ�ͫ�Y�
�7=n"k�P����b��5MbͰ�%t�����9\�M.�6�ĺ�R^ R[�)e�)����\C%c�n�F��%�bꬦΰ�3�6r ��D�v�:����7�<��Ś��^T���1���
�)4"�b�-�[n�ډ��)��h�$�>z���6F�7}�{�מI$��:D�A,��D�~��[�Y˼6v�I �̙>oI���"�]G��t=�(����`I�q$��$����'��!�5c,�%�	�H�b� IL�.Ȓ	}�0{I�� ��ۄ�	�$m�\u�\	����r��%�m��(ݙa%���ȐH v�G�'Σ�{9�o�-��wh��x�P��G�q�IbA�vĂ�7��.����$�3�,}���{�����@�.ˎ�}~����e?|���Y�ɤc�I�G0�T��Z��[yQ�8��3�-;��O�A͗�� Iv(�ِUz��Y��t�t����b)�ψ( ������	�kn�m�T@"o���,�H����9��~�F�	�z�9�O"fQ������G���L��9�ؽ�3�m��2���j�2�41X���ī�ȒOot)�)�>���&��}Ws�H5~>�""!'&"E��ȒX�o����`�y�#{ z�4p&�2D�,	��&`f��?%�	�]��ӽ��-�5zv�v��w�$�$��2I%oj�w���Sg1��񧃅���Jx�5=<�l����X2�a0=�<3���BX�}}�$���D�/�������N�O{�:2���.����-C;B;aFkY��pY@�՘��h�0�Jz�����"^"Gqw�D�H;���2B:6d�ܒ��$���f*��F5�m
n�$�7��	�%<,�ﺩ�0/��dǶ_�K@�^H֤X�F�=���wEJ�݃A#��۞.� x0�Z��dA)��tKth�p�ͻ�����-��y��(��/G������/���~�>��6�m�ӎ��@V�j����v.�7�s۞I��ğ{��W¡=��Nw{����;��G����˙/��.I���JP�1d��]�%�u��;Ѿ������0LK7t��G���-���3{�y8py������+�t��;�_��<�:��J�<�Al\tb�3�{�yz���xs�����X����MXg	T���/�b����<����h�mXq�j�hp���{���zy��y829\= �3�x����Oq�|x�x���/{K>#���C�K	*s�s��w�7o��
gw<a�g��wP�&�{���/{�y�w�4�=��ܽ��� g�ո'����>սm'^؍v�^E�w��i���|=�O}29��i�u��;�K�c�^�[��O����P��?>�<�pn/kL���;G4wv<�͐�^��m�P�9��Y&���
jP7LFZ�f<(e�d
׆�*��]cp ��yz]�a�C�b���[�
��ɓu/c�/tV�o��׻��*M�:RѤ��蓘'x��`��CH�K�n����|�9��Em�x�{�C�2R��Z���{z����J�qְ\$�SYH�e�6:u�2���t=���@�L+x~�Q����{�i�::�������S67��7�y�0�J��cn��5g(�]�ֱ3�S��h��7}߮�w�߹ݾ�~::뮺뮾�u�]u�^�T^�3�Ts �1�Ç
���p�3G#Ь��0�����q�����}�>>>>>?���뮺뮾:κ뮽>��33���Ŝ䧜�+��ن-B%5�T%+�RGn�5�$6H�Օ����H�fy�G��y�&��c
jYɑKZv�}X_��RL9�X�&�U�6O��{I�,��%F#R�G�&����|�S﷞�<�C4MR�=�ל=J�\�mi�k����t]�[;X���\��م͘�D!憋P�5Uq�ZͶ��"6�+��+����Y�
�[a�n��N�yWj��{�{�2�����*��*��PW��޹"_O/BE]B�Vp��'�U��[VnV*�Z�j�!5��"�w�9��{�vH��wd;b��"}0����IɈ�=�s���� �����D�	*��H8��&tp39��i/Ue����{��-!���{J/����햒�����;-��,�}�(���$�&Oyr$8��$�v��#�{z� ��r�`&.��gK*[�F��B��Z�kZ�Z�Q���K�����4�	���v�-�8�G��ZK	�ޑ�u���H�;>�}2K�.D�� u��(����^v	���I�,�w������q���Gṉ!�`���H�# ֯N<��mjt��k��wx
E
7qS$� ��r��2���w��AW�2b�ony��@*!Bs�Aou��;r���!�W5"Ik��H5��{��=9;v��rs��'+�Q���AҼ�ic+�ك|Ǽb��\��A�:V�b��}� ��ɳ���;����;]��"��%ͬX��Z�?UT�\��q
!(&"�<t&�����_g���NPL���e���H�!����|"i���W���չf­Hݪ�#S5��"̶��sw"��:F\���g���ϧ˾Z��'u�b��	6�q d���v&6��.���CG��2>�CLD��N4#HO#�g�t�k$��֋����H�����$d�(x��;�tԒz\z�w�=5rm�2���	�/v�eq�KN7f<I�!�R�V�ׄ�[��D�)gY�� �K����x
G����Ig>��k	d��VD�  @':�$�A]�({�
��ݒAX	���I8�=��w� ��	����0���3w\%�C�5�'v:ZAL���V�$���_��9���9���]�{jt<��+��w�����xr��Kg��^��;�;��=tĎ��5�w��s~	���������S��W�XX|���2�k|q7�����֫��Ӛ-.�j2����+v�X�Iu�K�Kz�Y�$�6,�:�-�.).�u)��&��E[�/\�S[ce�$i��vN��]��GR`��k�t�46tf��FVˬ�F�lR���YR@���RV�q2�]�M�&���1LFɤ"g�m:�#r8��nK�F屍���v�K�
jcK[E�!K�K�4�mf��	����[��b�6Q?��K�5�0�F+���V41�j4Ќ��6���_O���mh�g�}�� ,�6%�9�l�2�u:�o�����;ݲ&�NX�����'u�k'�Ȧ4K@�=���bؐe�[ٱ,a�3�1�2$��V���`��G`N8#HO#�ϵ��8��יA�����i �Y�.ƴ� �c�d��_Z<#�x�xo�O�u��6��[`�9�A"�&L���xx�������5��gT��7Ƃ�0"�T�ڌ
��I����G����$�I4��]H,HY�"qWEnD�UA<�`{�^]ӱ*�t�R���A�u�֓P���	چG6�f�T��i�]@ұ������?v��D�H+�e��	e������K��?T̂IU��j�[�	B11���a/�j��{�sR��;�b��xDBʊ,�͜�+$d�9��f_�l;:o���V�����˴g�r6b��ӛ^��sc,gވ�`1D��q���D�D�������l�s	��i�Љ��'u���$�U�ĐA���zS��K��Q!3��v>cL�h{�q��Bx���ˏe�MWg���D��I��Kc0���oH�@$w���Wvp��H��L��&�w�����G��\	b;۱�8��|�p����1�I+�r%�2DoGH�Go�go�~���Sm���XX�]�ܻ��L���7@ZM�)Yc���3���߳�=���(�a��EL��A�:+�"X���Z�w�F��^k���U�"kVǷx
�P���~�bX؟?^ԕU�9�a�-�y�.��%�CowL�Tf��4������d��x�P�#4٘�D�ă~΁ �2R�;��sA�������S��/r^��3h��쟞�k�^�ڦ�} �ۍ˸};}I�u��ѩ/�gy��<}�%��V,@���̐%���I�L�{�N� �a��D�uû�ا�V\Z�nY���$��D���ɶ�E�c����j�)���̉N�O��1��O��$y��N6�U�'��H�UH����ݑmL�GtF�e��^��ԡ9NS����@BP�YA��yebr��X�Af�l�������g�N��.�x�9ؓ,�'��h��ڻ*X�_�������� �$1<��%����O��X�xYo��x/K&S�����=4�7��i�Y �ye�ޮjCF�����U�����V��嘓�����n��={��2�o�"K�sF��f�����à� ��� ��_�'�nin�<(P�#a{�6;k����SC,cy��H_�%��w����3�A��Λn���k�(>����FN�����Ⱦc����UAt(�=/�1�%|�Gݢxs91z�y�g�o5�9�ŋ;!��T�ї)t ]:�ZK�	>����o�wuԇ��7y�"�1�5
�)��.�'���9�N�l���+x�oY�ϊ
�X���ƗLR���̀0b%��[r����6.���hO߿���	b#�+���>\�� ��B@;�ԏ���Z�]���A�3}�	�x	Ò�&��{�A� ��곹�/\wNǁ$Č~��,�%��q�ew��ݓ��{�8��s��qp��(�6��$WnD��ۚ؞]� �{�C��D�%����x�(O�~�P�.�w�Yf纄��~ݡD�F���v��UY�6A&�$Kl�P�BP�G�ޘ�H{��X���Z��Z[5����!25�I�s�͜P/��B�����מ��)1^ۇ�ӆ����D�^ĹUN\=n;�ǎ{i���1�?%�(�����旁Ş:\���X�"L2E���{�������m�'6X�T4��6m�J�0L@��)���U��b"i�(2� m�ʆM5��f���E�$�\�1ͥ����5�1�����l��ոB�t�
E��YkJ��$1�s��2\�U3�)/��XK!c�lf,� �R)��x�e��eWl�ju�� - �(q��*Y��X��RP6� F�|�d��	�ZA�A���:�\�� �*��]�RڗM3����ߟ���b�|�%_�	"� ]��,	$��ٜb�i�-}�le��Mr�}p$��W@0A""�t�:���矆J��l���J��I-��#��/N
�謋�{�g�p�p��%<MG�$��u��b�N���{���}��2�v�t'#$Ke��ݲ&�E��<<
#�ǲ+�c�+OA3������[��F�L�#_�Q�����W�;$U\��i ��w>���B��3Fzd�A�Ι�~�#��ӄ�>h��%�vtI�(�GL����o�3�@�-���[��kk4�69�M�����2��Gi�E1l������(��~K��g�?}vĒM���.����w��'l��ܑ(�-�Ϊ$=�R�@�uû�~ْ-�����r�6|�<�x����r�|A�K�
�紘�n=��/r[�*�4����s��;�]���Y����fv���5�b��20�b�od� �&`G\�b:+w�êh�}�SEiu�H����$�*I�r*q�"N��֨�v�k&й���bI<��i6��UX�B�\9.�W,�zz�!��X1�16�$�q�2��	d���<vP�B�୼��D�d�!5�i+p8xx
E�6U�Hyr୾�%�t1�ϭ�#�&I���3,B~�'���^�G�s��"�$�CK�����gG��3B;#k��aYit��Q������}�~�����n���%2F�:g��%�:D��{%k�E$�3,e�cQ�2@�(����P"%�S]����,q��@��SΫ�=�z0�� i��Z�.H@�- ����}��0h��]K�P�;�x���yM,���$Cx����LE�������<#��(�a�@��Hz|�C���"�1�:��o/{??�{�߷��||yr�B�N
�@ �y��˷� �u��X�rA��%�H���e�ӓ~���̓�d��A c'��i%��f�*�x���^g�I�V,���K�{���L��K:fdp� ���K���W� ���2P�0B\��q�{��4J�۶U�d�2G5[c�R�ʚ�:Y���6-�D�������(Q8ة�2Dr� 2D�;��"����R*�bb��Ze�$={$H$y�ñ����
���	�J��οO�<�6�^\�$YWt�	�$p��d�AD���{���2��;:T�	B1�ӱ��S���-l�3���{��/ݲ$F���5Sa��.�wy�x�5n��^XL��uD�$�׻�1������J�N=pFy��h��7��ROg;�I^Ô��O�ވ��o��}V�,�7��Q�H�b�!���A��,G13��	;�l@�""*�N̂A �˙;�����;0$b��K	$��W_nI�)& �`2
�RR�YKj�d�K��h���l-��ѥ��*`X,��z��~�p�Ď㓙A;}�<���"��M��`�Д,^���\�c6����Vpp��(���YK7��G��w)���n���%� ���$�
��,PpAT^�d�^�tv�8f='�$�B��[�I*��A>d��Vzv�.��c$�K_��N� ��2Z���P"%�WGBg��ɳXI�� �J��J����FK��y���3�JY�m���wz����;����"��u��rL�t�$/_L�A+:<�O�����͉0o�W?�@�S�����@F�����A�}�J��ʀC
+B+��ʋ(�ʋ��ʋ(�ʋ������+(�"���ʋ��J����(�ʋ��ʋ���C�2���+�0����0��+,2���)�2������+,2����2������+�0�2���)�2��,00���0���+�2!+0��� C�00��J� C�0���+,2��w���d�1Xaa��Bea��XBXea��VHaea��FXea��Xea���V�RXaa��VXea���VXaa��VX`a��VXBXea��VXaa��VXBVXdHaa��VXea����Xaea��VXaa�����PE� a `!�a ` `D eP e aD ` d=s�!�P��P��EB@HTHPHe��AR� ��G!��D�HhdE aE!���THhaE!����PENs��DHd!�D��P������D�d dT dT� ���1@��@��@��P aP ` `D d eP d:�<\apQ`d$T�eE��X`d��0Qa�Qa�Qa�VQa���?�^�û�?���R���*��2o��������C��G������Q������8c���8�`�3������w�c�� �(��?�?����?�TE��J*(�����?@����4���?W�!��
(���0|����K>�ܞ�����D�3�0 �K
�� "��@*�¨!B�R� B� ��D �
�(�
�@K !�$���!+"!ȈH ��@�H��H�H2����"!"�*�(�"�!�� ��@�B
�!	"! �(@B(H��2"2BL �@4���IE�?�E������?j��#H �@ B������������?P����:@�'����i((�����ǳ��?_�?�8u����#����Ln�G��~�
(���C���y��QE�DQ_���?��O�������(����<�
�+�@c��ژ���a���3OA`A���״��xI���}�� �@qAE�S�O�?����C����Q_�ω��0?���Cٿ��~���[�?pp�I�������J
(��G�#�p�����PQE`���'�v��O_�8~�,��?�����^�<�$��}((���������	���=��������o��AD_�=0`~z�TE�����O��bʟ�����)�˜ݴBϬ�0(���1��UJ�)$UB�I*����RR��H��	T* ���B!UR��)$�H�H�TQUBH�*
�� �9(� *�V�5�f��(��JJ	�ҫI,�E(T�[1+F٨*�Y}���]h�T�����wi*��J:�YT�{�                                     
��       H��1 �n��Q���  l� ��2 �d4����w��<�V�M4-���
 	����<�  �ܼ��4%;4�r�)T�7E�i��P��� \J�(Y�w�uJ$���]�ʑy�
�^L\�R�S��7jš�h��  }         ҤP��J�(Y���nP<�R�����|�R�=p .�
�M.��T�yaT���W-J�R�q��P�O.  "��} u�6iEP�*_z  �y�M7�t68 ]��R���J��+04v�sgZ��8 Ӡ7{�ƚ��My�R��˙Ӥ�E��   �      � >�U>���t퇗GSMK�ܳ����x I�u�ۊ��p�j۶��ۛ��՜ ����m.X��m�����    ���[��͞�6=� δ=<\u�E��z�q7�������ђ�� wN����A�-ڬ�\θ�fk��v��ѥh�   > 
       ���s����v��]o6톧�����k�wA�nv'kjӍ��F張�N9����� �T�M�9�ƃ�ܫ�J��ͷ�  ��M�n�S\�:�Ep t�i����^�;P�T�%^#s:.6k� �*����=²�6�^��=��3��P�YKf�
e� �        �]�r٪��Os:�N@ � �-]��!��@��C��� Ϻ���8��P�5��� @r� �� ������ n����(2U� p����@r��5_ 5<����4  EO���T4 5O`�J��� D�*��I@ h5Oz��*R�  $�ALR�� ������ID��?�>����K������
8lRO;u�$��	'�&w�rBB�P� ���I!!I��!!I��BB�������������E3�N��v�j�7r���o,�9���L��x����7���Q�Ö�"��8u.-٣ �`zI4W�p-[���l����m��ݜ6�����w�AoG.0r2�4ۮ��א����d��0o>Տ�u�$�dn?�sS6����l���༴9k���=��9�,��K��h����л��LS5�ۋ�n�*�]X7��R�qq�f�Kq��-�9��7\0^z�v,F��j�����+�X���y�c���E���	�n���3��"����Y����&j�-	'u�eh��x7��ٛ�y��t�ٖ�0:��kӒ�u��6
872ը�*�@���pOXN[G{_v*+��� ��%%��;��&A�K�fV�	��3{�$�IB[Cm0 @���N9��X����e���v[�����/n����Ƚ{h2����$��gw's����2�ç:u�y�9��{��3d���.��8rm�]�Q��8��y�'%�a�Aٝ+ތf^]ϓ	��*k���31������b�o>8@��YE0��{A�-�Ѓr�5c�%TZ�,��t�:�#{���SUӱ}�w�iWN=�%�oL*Ή\�^iA�(ǥ�7�w��"�d��v��əs8;ٽ]��K�X��K;��M��8�]\�n¯a!����b^fj�&�e�2�ێB�=ꁼ�,��}��x��n��fn� �q$2��=l�Pl�7r<+�Gw\Uj��oHm��f���Ԅ�o]4%�q���T�6��hޘ�m;�n��>Y(Q�6��	�c�����[A��;��o��:m�ߍ1K
[�;2�s��{ܻsAG�0���5��_l�
f�0/,[�Wg��|/�c�-�=S9f��2�}�*8F�(#�@��,N�8+ɍ���1v���v��h�%ƛ,Q��a�o1�YJ�3;���5rP<���
��j���\�+�6@ �T����g&eך���P� ��Ί�қ�wNq��F+�f�a$ژ�����Ժ�N�AǗR�(�b�tY�t�M��ܷ��*�T3vˏhI��U����':$��Z�4��x��t�L3�Nc��I�VݨbGR��v��kD[��3,��n�T�Z�4\x��1�[�Jƍ)<����wi���x�D
������l�Z�qVw�] %��CS70�d�j�B��]�x$:�8�]t�7��9ʞz�x��r�2bz�Y�PB��:��|�N5]��xҶ�n��[vj&ɔL�j=�m[�rNgtA�p@��kk�E1%��{�VͶrX���=�){o9"��hP]D�kW�)���C+�;]j�r:�!�WAg1vs���PͶ欋�Ƚ���&(�Cp4$���>qi�.=�ݶ5��!FF�;�l[�[Zc��jܤ�^ [��4�g4�BU��5�=LPi�j7��sݮq�)w�@�Փ�����P��θ��I�1��oE�=���k��qNŶ>�^�M��l��zT�ub�.֘�z)�#�c#��Æ��+p�<�L���٤9�\��)�5�׬�2-��FH�?���\�7u�cS6�*w��&�'I	]P׬f��i��gGIȟ�+x)Vr�2�o'��7:�,��86�r ����f��Hn"��e�l��j����M���M0үw�9ӨYK�3��ʮ��ҷ���hf�ym��=`#㻱���U���v^v��D�_�8���G�<��$�dy.4�<X
�i]���QdDzRh��5�'p�j���XlÕm��0ܫ&�:�t��y��w�3�V:��8��=�%�;7��;(�ꡓPf��Kn���>��p�y4	�f܌����5bUA`���A������_�E�U(���9;�{�=r�V�U3���\�m�X�-���خ�p�F5;5(����¶S;U��S<�N�ǈ)�޳�[����îm۷�n��2^U�5p�)T��Y�b%���i0�F�f�Fۉ��#44Q���Ev�H'��1��A�ךp6�0�ΦV@��`���X$�yG��;��ոy�v��?�Gbg`١̝�����q�pʏD�.�A9awHs��L<橅�&\�$Nk����1�o�������pj1����8�5�QIj��a��]Z�>�c�ig�o[Yi�ƮC0���ɪr����0
y��苮��9�:�<�\J��B3��AS[���T���gp\�_����~�K��{����b38E��!W���u�+
�	�X�v�v#��ե>�75��RhW䨛yn�{����,�ɫ�����"<}I�:3q�M�>��k�0b@�����ҋ�+XBT��t�&گf�ː����BiB:�[+�û�F�G�N�.	�N�$`��Gv��̒�ٵ�<�w�z�܏�!G�3y��D�z�&��r!ْ.�`��l�ػp�1�)�jod�y�С��e�4m��H��;�̐+8H����n��M�[��gQ����ڮ /.��ig^k����7�����h����Ak\�F1qS��-�^ˋv��X�s�&vk'��cyd#��8&SWDl�=����D��=��=!�3fT��p���2��=H���Z�0L��de$bw
o�0\��5�y�17p���M�{!�3��sRCb��P;���U��`�-wGN�i�%�,F�Qx��������0���Z!E	H�P�Wc1�J�!��{�T��0,�*���5Ռ��L�|�.=��:,�Q��5��u#�{�F+}�93����4�h��7��f�Q��q=�(=�
y��Y_���D6�x҉��`�#�]y%&��(�����#���n�����?����Kk9�a(�6F�@�;t��pŕ�,,(z8q�*2�i���E�)!��%:���""��sи������ךa8ע/�k�y��ȳ!�#�,�#@�ͻ�܏-��'ΐ����8���\/'l��os�%R&;)�It��uT���2�Yhb��<Lk=]mdt�E��Ef��xۚ�I���'$9=xs���:�.�n�4����F2�
�ŨLw���)9�v���MҩH'�wl��A�0��-���J^h#��Yi���{�pM�C)&��#�q��1��R��ڸw� ��F����Õ�.��B����q�e�1ؑ<ݦ���9��L�_dZ^q�N���mM��1��2�f�㗮����۫ Dк*8q����갾w�n�Tz����s�s�5d;ϟ<�|�6�̔F2�!.ι����W'1m$s�%u���d���o>[��y��f�q
�e����oW4,���{r���
A� ����rF��e��ՄWm[���s�'fK�N��$*�Mq���^�V��a�e��86t��������]�8�T�M�wR���p�oi;��T����$�r���G�o�\Azs���7\yw3i���D�q,��B�f��t��l�z� >������5��a����q�]�=�?Y��#S�ԡn�1i�3y��9	bjx0�d�:Z(�f,�ϳx_��Ia�,-� ����wRc�3���Jܰv��ͬA�s;��ģ.eG�>l�ر�h�U�t�Lv��>���T�n$6+ӎ��u�n�W8��{��Ӓb�ۡh;0I�i�́=�gM�%,�c�ʔ��lɛX���N\ ��Y6���פd�1ud���I�i��s��í��]�:k��V���Vwfr�hz��zrQ�3�[�xW���խ�a��软��գ_mV �ĽyGoe���t��&����#p�諃�tv�Ƽ���c�h+�ԉ�Sg����97`�֏>�s�.����q�Ӽ;p*�D]�/8����N�e�呙�k%��ڱ�Otz�6E^ft!��#V��O����d�->�Z�gU���1�40g�d{�FظB�ƫa4�D��J.p��N�k��Y�&�iႾ��0�5�햠��{cf��h�2#gN�!��A��;�4lFѝ���H恥J�V�����[ѳ2��ZxA��|դ��!+4ݶr���0��e��*�Y��6r�ڵ�a�Sʦ<��jή�%���:���@�tF�ܕY���97���ח��ۦ�N#a,״���v<��sZ`�ŒM�6WuȰ�Vq[&��:rb�P2�����%5W��9+��͑��1Υtdw6-7MZ၊��U ����&�!�B�b�VM��"ݚ�;Ԯ��L6.%��,32����S/l�ˍd�8�@TO{�l�^���C�����Bd�8oI��2�fvn��':�:Xg�6c�5��f�{�#��W���bj
��{@^G&�Qv��!� ��Ҵ��Q2uԛ��e��v�E��G#ٙUek;�9��bݎVGI�XN���f�d��G}�+�oL#�9��Lno^�3��&+%�)�w33��˅ΰ�<�ǰf���7K��0mƞ( n-UfA�����ΥqI�� }�h�B���!D�� a�����8t�%����ՒS�v�ߩZ�	0J���������0^�I,����NV�s:�}�Q�����C���{������P�0�7%$���9닱;3����PA���|E��W��{Ge���w����r�� ���c��[M9�K�Q���iwA�ܲ��R{�d���7(�'�(���b�n@�ox9�ۥb<�;���|��1��Ww�n�\c\:q��Ѧ���Eа)�媱��Q���ìh\�3rr�S�;76�9ҎX1r$�G�杓C(Z�e�B;�Ⱥ��}%C4g �8�=���ϕw낌�a��{;��:�坏��%����� ���}�019�����0$~���:[�*O��+��qj���3э�i�V���Hٖ�{�fFd��Gp��N�ƙ��&ٕ�G�Xݛ��V8r�����M�qb.R�5�ф��B��C+��7Kn��鱭���}�/��k׺��ugty�9��n�'z;#�����jĳ,�;]5-ֶV��!.�i-XѯW^qтosB���v,=���IUB�[�3�X%}zO���n鹰?K���^�n��_�{lZ�Bz#'#w6Fo۝DP�����v�΃��ga�/����+�;j�����[��j�!k�S�z�7*pE�Sa�Xu��=��'�t:I�5��"�����@�E&�F�\�9j��4�H}ܢI�Xd���!�@f��%]�2��d����xq���Q��8�y�Ƹ��`�'�IIEõN�"K��Q��`ޢ��"B,<��{
��#"���!��1�;�rY�Z �	���*�[4����N��܏�����P���3r���?(�b��3���$��݃��͒&�И�n�pq\`ס�xBE��'T�b��$=�N`�ݜ��	!ۣD_Q�uu��d�%�j��U�lM�}��=͑�B���ó�b��V���y������\Z{������)b�Q^�߄�gu�^2��T;���WZ��U24�8��3���"K4�2J~̰`���F防�h�w{��.��D��Du�ol\
R��ݚ��%�9�� v��t���b�XS����y��N�o�� O�[a
A��i/S\���m7wG�j��_����Ro�VE��c�����n�%�d9����O\�ko�;���W���aȸ�'�	H������J���B(ٶ�udR�����voI�+�ڏU�0����5.3�qr<�M���Lh`�0�p��Y�睖�VT��6-�.,��l���x�+��I7��K��6��4�Pfܔ��*Kq^��`�n����ʎ=�{��,|��o��.��������f.��B	s#KZ{�G��+ǲ�v��Y��R����ul��dc&��~���.�62�z9���nx�gMN��n��u��Oa��X�ø�$f������y�PEw>��=}�񱕳�[�#]���	Ӓ��䒳�9�X�J��{C�p<叱�w��дt�KF]���^5������w.j~��4@�T�j�p�9��MUh�wfreu~${�Sݞ#��l�9�[��k��hF!�C�.�a^�ç�p��0�9��C�^wiuZ���F�ŧ��n�2�	X1���^pQ��!m|��|$�Վ�v��k/`5��݊�E�f$�Gl��t&�'�.*�:�<R!�w\�Pi�&�����{\!��g��gV�v�7#I�����A�����-t�ܕ-ge����Էb��X۩�U��;9g_Z�'�+	���ɶv�$u�#�o�įKv��c�Ć���\�V+d76����(�h�I��Y��sU;��;��4�����q��6�6e�
����{�>R;�0,7q��g~}��.�=U�[Q1Es��r�Ԛ�}�ˁ=O���>-�u� �ޮ��iߤk���?��	����@!���,�� ��`E�$"�BA@P$�I!Y �a	R
�P� �a!RBJ�I�)��T�P ,���dP,�,@��E�� �dI!R�VT$+ XB@� a`�B)Ad��$��$��	@�BH� ��B�d�I"�
 `Ad%d
�
H��"��@*H@*E� E HH,���IE�$Y E�A@
���!
���!Y$�d�H���H! 
��	� AI �*T! ,!� *@
���$�Y�!�􄄄	"�	O�HH@�o���J�C��,����"�+�?��̢�_Η׳^�_{� ��i@V�7&����״nS��k��Ѷr'�S��uqZ��y/��tr�K�}�5L�{[
u���uj��J5��a ��s�˝2�9�5�ˏ{q됿rs��	y�T��ny�Oo.�Y��Y���gEHg���}ta�|c�.O���^����f��<v3�)w�1���{/��ʗ��Ǜ��.w0�7&B�� ���u�'�p�����.����i�%�8���<�z�Ё���s�S�a���y�ջ�*H0V=��{g����KJ!����}��Lp�5Nr�{/+�l��	Z�8�!
�>�B��C�����#���F��{�>��ދ��4x�)����,���5�-yz���v�ql�C7��M\B��!��'���S��@!ُ1w��&t����������/`�}��{����ܩG�I�{T�G�0]<��ܟI�K(W�v�7MEX�|�xύX�稼��-�����e���kGÚ�}����Oa[8���yd���0��o0��:�3�]�W��g2F��-�g����]ӽ�u�}�s��{Gb\��"�1��#���1�C͙��W�w�x�;=� 1Xܑy�7yo��2N����J㉱'�o�ڌ�L^�^��rޘP���!2<���o���d��r���]|\�|�0��d�� e �<��{4]�i�C��N�
fsawn�,�l���u��	�Wn�f���c8vx{_A<D�sB�zn��> Q}ϛ�;I���^v�*`��x���0b����=z&�ء��nfN�f���ʜKt$5qO�o���c�:r����r�{R��J\����óާ�q٣RPW[��4��1��{�wOp��[�}��?,����=�e����! �3ã�M�9�}��=��.V����"��*[�4t�:�"�I�#�Ǟ��9��O;0�	-��Uc���g���F�^����x[A��S���uk���ysʊ��E�!ENydf첼�f7���ݞ�~hV�+����_<y^�f�K���_|�����<og��ϼ�rgu�xp{H�j�{�d���4k�;�Ҧv" C��X-Ͻ�	(Uͩ��f�cK�4ǻ;K�[���<�{�bd9;W�H���a�(y{ %� ��Fǆ�0�rm��m�H����7�#�[��j��,�~<�P[:�φ�M�X�����N�Sy�geaU����z`�ˡלD���'no}!�����9� +#�令Dm`���)�L��G:O�w���xx+��9�Nw�?���w�e�L#O��C��x���;�8�Yv�N���)�$������!�,R��4F3}�e<�fŻfF�D�9���{��/xQf>N�74lg��g=�O���1���{Lͅ�� a�{wۊrt�ճ���ޯo�m�Aâ�.��E�ܾ^D�&�d�S#���5�����������P"�#��_,�4
���,<�{�sƢ���]���z�F�����V��KU�������A�g�.-׷��Om;k�U����gL���Nx]�o1w�ZZҷ"҄�35E�AĲM��k����|���L~	��_��O^=[��[�kf�	��ٌ��,wx{���b�>ɮ���ă�n�<_B.)ﯱ��>�&��#_�Ђ�匣���}�qzy{O-����5��R���nW����'_0�aC�!9�I�{�/6jʻ<ncG�ߊ��;�<�<k�ؗ:�>���U�F��W�`9<���=�5����Ÿ�so��{��憭�_Y��G�;��r\�D�g�5�MOݺ��lძ�_=*]u�����}3zgxp)ψ�^�Cк��,l��Bn��Nä��hkCͥ�Y�7�3�@��T-�z^+һtC5xxe��_]��۞�/;.�5D䍻팤����R߀��{�� �پ�5�(�F)�<�"�����k+W�%�}�/�A4I�����zJ<�E�����z룰��{F�C�=X�Q�}Ҩ��_����$z�\��}}�Ż�
�p�2��[PhY�GۻPŐTnS3�[r'��7�{�\j������k:�=�G�A���r�S�rz��7�2�ΣÀ�+��#�n�^SQ�N�sVJ2A�3(I�u^����ߗ��e��yVZ}8���3u*1 E[L؜hz��鵎�/^����A��5f�X�.XKcC�xb��4�r/�]l�/e��מW*# ����Uf�h�ٍEhXSw���=�������i��wQo=�8xY,���x�\0��3'.�,��;y���-�������|G�������;��w��Y�(]sk����^�66��X*J߈��my����=�����S�w�z�����É紭�[��^>��p�a����0��lɺ���
+���^/Y�\�*I�}yťq�<��!�
,e2�n���7�J�lh�t.,��H�#ouCOѻ	�a�7l�ne�����3Zwx�yN���Z�ܻVe�33��u��%�X_7�tX���U��bјϊ>�C��F�+��+æ1�Fr[�k���+�&�!�B�����H�T�� ��n�6��N�Z�*\�&��=���=��oo;e�̝����6�͋s���^�/ވT������B=��F�����ty�z�f�,����P򡜱�\�V
q�R�¯'���~^���D������s]���l�E';�e;<Oz�۾h��]U{�h��^��nY9�pm2��5��N�||�}h�W��L������s��p%J�+�JN�G�>C�~G'>-Go�?�7�:�כau4�}�����|aD�b�h\����PS�"^����֣O�Pw�Z�^S�^�4�؝�f7q��"3�a�.��{�2�`�$�?oq�� �[/��\8�����X�ڿ��/��o>ԩwYs��П�h�ǅ�����N�ݏ������<�q6v��O�i�h��Nעzoe���/y5�;��Y}�g��v���y@��ս�u>̆{Ȭ�(����Z ���V��ኛ�L^��ޔ 'FpL}�WA�r긌�̵�|��Y-�=+�yE9M����k ��g���	��M[��jb|�=�cK�&|��6���{�8њgK����8fɉ�zImT/R������q�r�˶�,C��D}b�a���ɘ���OC�p�_���q�_ww���K/�3;�݅�ݔ�%8��d��X��%%������z	�ޣog%CxP��<,�N@��䂸
���:mDm��
��/w�)ޒ���>���w�:
T���@������_%�o��\���U���LN�蕅\K��u���0���n�͗.�kN����/)�����F����W�{�j�^��+��%�욗T`�}�p�_	���#�,�����;Y�,i9�~a/zyy�G�c�Ԧ�t.sؠ���z�В:�H�5���yj�٬��J k�Ej϶���*`>�;W�o��'�px ��=��On>T��k��=�b��w�5�աW������c�h�0l+�tX#0�n],�hd1��RA�5.>܃��/r��n�J��7��z6L-)�eC�n9�Tg��{����m�p��I'g�1�cڍ�^M�p�=V>�vo�908�n�������"g�3�kD-ѳqۺ��у�����F|�M��]�^ۥ_|��\��ꗣ�&�L��&�3��X�g�	�,�z�:{�${��if�ٗ7���y�rE�����1Q�G;����p����8?nl� �k��<OK6\Zb�`�#�Ts���X�n.B��囷���7�=�x�Q�)M��;GjH�;�&���8́�޻��N�=�i�ᾒw�:/{��2�f<���r9n�L���u���gc��hQ��ސE�G|V�f��l��S��߆���ފN֮�f�ा��sc6�N��YҊ���{Wy	�ߝ>$�7����(�H* �wg���P\~�O��)�e�^�Lx2}|�{t�v������t��m�bj'����b�8`3;Z]NLk4I1V6k�v��z�����@�_W���0۴��[r���Q��9�G;��,dB)&^:G:{5�[Cw��]�X�)|ǻ�Z�U�ٰ����b{޷۩Sg�MvZ����6�=�u�c��LN4�M!��ٌ���4�Ԩ�<�{s�\���_-~�=[[��_��$ɧ���oo�)�!	�o2����g����X��xq�}���1;�78���E��ou*q��v�zH�x��o�fu�,�]�#�¢}H򫻽I�o���S|#ԭd"l�;	�a��zsZ�1$��'�G/v�w�m��p��e�~��M睵lO��Z�<{ǚ��<Ƴ��n%J׷��9�h3�������I�<z��_^ �?oj�5G�{�[�|��k�jݖ�.��cZ�M�A�O5�<Rܓ���hξmZ���{w�P��/XݜfZJ��k!k�=�!�b�����Q��/."�cg=���3T��f���3YQUzF����CJ�8ߜ�NGF��^þaQ��vS��g�w�q����&搄�t5�l�*!�y��5�ב��#mں:4y�2v������v3@8��x�4���J�o
=�}ůsb1^OtW��k8���̈́�#,�j	���~�3(�O{'/e���Y~zyBK�վ���k�<�V�/������.Y�ސ��~��������ٱDG�<Z��θ �zz����[7����s����!��Ǭtc�D.�������l���oE�9���;d�)Ԝ7�Yr���%YQ!q��x�0�x5���5�R�E��b�^��ܸ��誈㔍�us�=BJx��Ѐl-�Qg��U[��}=�y������py���oL7��ѭ�=��0�'�ݗ�T������@���.U�C>Pj������=n�ͣ٭�T�9�,l������+}e�3ѯtP�ޮ���R-��W�ٹѿ$|�<#S�it~�;����)v=�䜀P�/oS����|n�x�}�=���nN�=�_5���z��&������/��DFXV�TZww�V[��<��a��f�*M�7M�{�tģ��W��ӣp�����/�ޡ4�����ӥ�g���`ʉb�>�FErg�c�C;��[��1n_^�*yÐ�p��yc��l7*��=]{7�%Rz7ҽ��|%�-yg#|V#c:󇕬L��V)�Ёm�y�����]�"�%Ƹw;wד�*��^���� a�n������Z��L�w���M=�1�^��C�^�#J��_���+yp�Ӌ��4�!}z�f�_�罼�%�����F#���}��!e�u����Vcz�^���\�Wx\Xw���Oj}�7;WRo�x����	#�u:k��Ǌ�st{no�yW3L��N���������zY��]��ξyog�բ�Pt����.�O`X���[�����#�n#.��.:�h�,>�Ä3�\�<�m��q7���5�4����6��ղ�����@-����)��<���)E �xU=�\�p�~�g��y�D�aߒ<�B�:pt��2@�s�橚L��X}�P��3������؛\�A`�L�A�sٞثC�&��0�,�E����,~bt�	{p{%��{�aթ���;��h6��g����������9�;ݙJ��S�H��-c�c�M���V����n��Ш�����3g�|��'`��򝁮ε��B�����F�YHKK��ն1��w����@�C������dn����>jZ���/v�*m�[]Gro4���{/E�zxw�얫��=}��O�B�/���}�藊�1��\��>�=\���2͍b��ιBu-��n3�]Ћ�F��w��gf���&���}����E��>df���2A����U����k���?58E�;cg�z�} d,�|k��{x$�xg��8A��+s���Ws��*���{��$^/.�����>k���C2t������_�ٮ���EC����_{٩"U�k�T�����r�}�2̓<j^ #r(��`�����Gj��l-�	�h1x�Z�涛�����]N\�m�{6�j-�GLg4q7��13�l�������ro6��}���s�4�Tz���]3�8 ݡ�l�q#�a����{��/���鮧�E�o��7���<1����x�!dr>g�_O�ZkS}��; a�b>��B���ެ�ة����/�y��<V<��Eɳ���gٓd�gy����d{a�q�9�~�zn���w��q�S��zTY� ��7A>��h^e��Ř$g<p�(�S��ݹE�3��WĖ�ƺQ�'
�u=����c��m�dð�tn�*�:�GwDU�n��\!���u�IcݐF�ˈ�&:/���;\���7$�t-fz�p�Nb�ӸQ�����UZ�3�=��>�f��Ƽv�~ym��枏p����5)P��[��){cOl�	,��L�ݔN��.#��p�l�n֥�����jg�$"{��C�c��9LU���>�w��u�ww����/A��&t�3�����MA��Nh�:b���Kܙ��Q9yGD�JN��̓�˩;"���5NN����T�t5��B���oX��=��2(Ɖ��{
ٻ�o�P�W#P �*���O_�Z�(�س���������M���֝j9�����4&4�x��[;i�۠.xlcf�g�trt�1յ�5����P�@t�N�iC���B��5�Ųhk���6M��駭��]Gvy��ڭ���z��d�M��{:�Mr#�ٺ{k��z�z�h͛�]����v�=:��U��ã�lGd�6.w[����=��ls\���]ys�k$n�GmuCu�݌�rTtn����N��7��*v=�t�QRS,��4Uɹ6��b��[���=�&�ɷ\ۭ�og�ӻvz\������㋃�γ�����6S�l�h���y�uf.��땖6:�M�;�4��3�)��������v����Y�V����lrs�`��-���'�ٻj����i���^z�=�o�y��h�{�y�Z�;�2�*ڎ8�gY�+�x�[�g�n`��"W���<�ӃR�v�+w;��;�K�Wbwl��=�g�7-�st\��*ݺ���`og�ݰK��ynq�Nf.d���{t���ׇ�l��c����Y�����).�Ҷ�6Epp�.��@e�f�8�v6�^]Ompn���q�z:9�5��\�K�׶x��ڶ���vT�K���ק�9y��g�/:��멶8��sld�b�ژ��
�^�θ}���=�`B�
��Il��*��q=<OC���[�L�:�c�l�$��lr�N=�2�m�',\��l��l��l�OV�!�+�Gcp��i�'�:�����tۦηN�k��M.�^�ۯa��v#�9*�ڋ&չ���m����׳��p�Ft)�اu�ֺu��<r]r��Y�mf��a1�oL]�S[�n������K�l�r&����{Rō�`⻮9���v=�A�x���{q&c���+V���s[��<���Q��9�$N^�O\��'��ff��M�v��l�+��������@xn�r�rTxgt9�����u=�S��`��/j��K�0lE���OaN�p��|�J\�x�ۂ�=�a3�(�ّ�����f9��Q�9�o,X�\rIm;<�Xuvs�n�8qV�嫰��g����gX���-���{���XeY�=��{���:�n泀7h�Y��kv��]̼�lf���k��۬����7P��z�':԰��Qry�
���n;m��>s�V�9�e����r���h6��ME.�H�Z�mi��
���W!ڙ#r=;@�unwtۮ��jcO8����Ş9���;��L��ܱ�m��]��g�0gv�Kcbŷ �t�gH:wgӈy���z�GW����q+a���^�c��%�v��Nr �<X0]=�E܌su����g�m�%���vn�yw]���.��u��W���n7ru��3vyn`���pc�G��^s�Rea�l�qX��q�%���C#�6�n��6�S���#&{{����9�4��6g�Ŷ��oy7�4��U��}s��&��k�ݖ��T�<v��0���Vz4�q�ӛ�=��h�tu�馈�q�Sfs�mu�ո�q&��t\��v�=q����zI�In���s���[�t"zB�uF�*�A�N+��&���96�P>a7({l8�����a�8t[���ӣ��mF��r�B����V�n7Lt��E�
�Űq���v�wX�,=�l2Z@"����-��zۦ6p�$�h�q�[e2��ܚ3�$[Omp nj6g��yG[��V�9���ۍ����tq���c<�=�sѻF��u>�q�<���[tn�B9/c�Kp=�u�&:Čmc��z��.�⼲����z�*�Nx�h{h[�`;��k��バ�lk��g�lc=<M��va{���n�g�c��8�u���n�w��ۅ�͸��Jێ.{[]�n v�v��v�5���ǵ�Q q�������9vvD���9��n�&�݀;"�Vӗ�������)���{Yug�v8��v싷�Ӆq�����ڻ�ɋ��.s2o��۴���u�G]��nm�oC�h�r��m�m�����ۮ���V��]�\�>�ꮂ����U׷���9�]Z3�j:�0t�M��̛���]��.�q۪�86�"�v��7=��˰���%�ͪ����:��r��z�J�j�ҺPö�Ć��i���)���sՂ��a��=��{c���O�ў|�1ݡL�0�q�#�7k�u8�՚��9�^�^���ͫvAy�ui���F�RuN}�������s�8p;&����u�=�����ۯ=ۥ7.j����Y��g�u!�su�x�kK���.5�ۧ<��3ۮ� �N;q��.x���nV䓭uƎ �e��I�D�b^�P��Tp�^�V�\��4eD�
��\m����G���v�;q���u�:�^g�s�ܣWi�fڵ�r\n|\N�pb�˺}+�Y�L����;j�cq�;�4D���=�9�����>�^U���w= v�۴f�Wgjb�y�ƶ3��v�[��qN�max��ҵΌ�ɮG�K�7��=dq�n,H���q1�687e����[c����ck�N�����n��)s���<O<�e�y۞z^�������m��:]�4��^|�X���s�5xNg�^����ruj����a�D�:�#��죳��v���[���.��[���m���q�;7��^�����\���b�li*�p:�.�m�sLk�ݸuTc;��]�\f۰QQ{g��p���<���0{,E�2e�66h؊m�x��u���[�l�mӭ'`m4�6�`�Mrq�y�嶠�[l��c�ny�g���۝֝vQ�����l�;
V�c�ggg�����5��dm�3�������I�!�ٞ�����/s�N˸ptmۈ�={s`�<���͓�����:7X�`��0��<b�[Yn�m��n���p�8��7[wZ=�n��4�W����h�a������݌0U�¾;h'<��2���r��c$Zyv��A緵z���"��&�Q0��zS�b�8Ѻ{gWM��:�]��^���yn)@,$��GrX{%eW[�������E�W#�6�m�7t�Il8�1őxpva�s�ø[�vwPs�M��=dJ����pj�X[F�q^I�r�lCn۟J���:F��;�,ɜ\��3zw	�N�u��uۦ{�C�CqV7��;r,�\Y��xɝټo%�먝�Ÿ��q���t��^���Mc[��#�+ܝ)˽X�9�m�>7�9�e�n��7rc;��	�9&ܥ"Y���/c��vι�c�q�kHɬvxM�����m��V�ۡ;r�+l��c/ʠ�̝x�Z't�r�M�p�z�v�m�6M���&ګWg��Q;ft'yۧkn��x�ƕ�^C��2<;�@i��sƥ���s���z��i��X����tgV`�ۊ���#�fg��;j�q瓜8�G	kq�:��9�I+k�����z���ٳ�py�ӓw�+�����&%x�:x�m� x�&��.���za�<[t=�p`�N��[�㭼pY�sGc�y[��B�<f��V��.��qs��׳��:;f�{��c7n[�e��VcV�\����׃�&��T��;,�7�̅윦�����[�N����n��U]�;#����u� �!z�u�(l#�l/���9�vĻ������9-��x�&��ۮr�\����m��c2�ڷf��I6۞{�/Am���܊��ڻ{C��A��v���/9�;n�"�v�Sv����vA
�[��սs�e���/n�V\B�6��=���</mn�;r&��WS�p7$�o8�6�9�N부�nx+=�:}R�����ϸ��E��fמ�ێ��ք-��9v&X�^�;A��q���a�5�7�-!��n.w������s�FκݻJb��[�.&�qc�s���[�b���n��ݦ؋�����l�k�a�#�@Ep;>��GN�p�ێɶʽx������H���ݖǵջ�o7X�Y�1�:[N�x�vI�zf�˘7N8�7;�y����1c6B.�0����^��m]����:ħ/�f<���P�5f��c���l�8�;-�,��q�/&���e��h��
�y�sT�YN��U�m(���%�;��nwp2�9ę�آ����l�R�ۮ�k���C�=��D1�=�6G̽s�8�ݲ�<m����\����'k�sګ����z۵n;q�	���㜂�=c[p'a�A8y�n���73�9�g&� �a�۷o@�pˮc%�f��������z"+�%���ny�v+�����v{����)�<�<V�m�,�=\�#gv�����eֵ׃��A����Ɍ��/9��s���x[���w5U\��%��n�R��7O���I�T����p�W9r�w=��v^MÂy��d�����t0����-ֹ��>�vg�9�C��>�=�.8�f�\�]q���{F�Ӽ���Ӷ\z�CY	q��Ŗ.�i�G���.5�����Y�x�ڽ%�nc���D�%�	v�qNX�,���%���wd�щ�,���Z�#�ډ�v�w���&��mqu�\�����ǲq�}C�n�l�Y�|�[p��f󷞖�0��4GR��̻��n�]#����;�S�p�EJ8b9�뺻ls�]���g�]W�֭^��P�ᗣ+[E��e3���]���u�ۮ��������G��[z^���]�7�z<�5�k�ی�V1 ��;v�Ɲ\pOco^�������	Zp�-+�g�S7	�f:Ę9��͋Es�z�ɺ��6��=�e\y[mpP���m������@�b
�uۗ�b�<Y�g���N���w���3o��/]cOK����u�Z�㛩�&�;{]��3�j��(��T�j�(���!jn�j�w����PL�ejE�Ts.,\�TfZbPr�-TUr�%l��Z6�2�k�ƱDƔ��q1��2��)Q2ٌq̭���14�-����ܸ&[�1Ko��!����ܢx��YUh��+��Z�W.c%V�Lf9kW-
�qB�ff(�-��X�ҥG2b[�q31���K��b`�enB���f���h"�j�(��mP��r�."�TX�´j(6ʫ�
��\�\LVئ9��J4F�����9�F*�G,��cr�jF+�[�jW�����n��ZX�5q�DŹ�̢�c�*�V���][��)��r�UQVZV�1+R�V�f"�PEb�-h��[Dh\�7m���n;�<&�;��9�B��E\,�V��AL��ۜLv�ۣgd�;�=���{5Ӌ�j�ʸ+U30�fcQ��Ki�fZ��J�̢����ܷcDW-*ڣR�:�t"�W0�1�(���ժ�Tr���G|��\ֵ\nc����Lq��`�T�6�ny��6�����gF���̾���x�//Y��@8j�9�.�p�֤�,ζ���x�2�b��5�>��
�[���f�۞vz!�(VU:;*��7g�p3��k���m�1��B��<0��Gt��n���5�q���[E�a�c�'m�;`Wa��nN��v�;s�W8.x��t�b���d�`ָ�>+nNa��Ƽwb{C�-k.֐�kkA�n� �:;���]�t�z\v�wC���X#�cn�.㇍��=n��dچ�[1��#�l�ڻ��v��%�(3e��`��X���X١3�cu�j��;�w��ƺ��m�zEp;j�M�>z�b�z�tv�����j���Ë\''^vm�]'46�x�F{Sˉ���{M��9�<��&ؾ/|���n�X��뱹x�K���n���v�ǉ\/�xx�Bv��e���5��^|;�ܽ�8^�v���c�q�|����/��s�ݎ�mu�O��
:wm�Y�^ݔ.�W\�-�ۈ��s�=9����-a�{��qWctW�ssbk�L{��Mɻ`�f4�{����'/������֗�l��Nɺ�8z�[�k�=�� z��u�q����1m��,	8�{ey���0�.����k� ����۲s����69���&M���!�ݠ�Y��`�θ��ٵʎ�_Ym��xN_Z�0��NWtrKt��i�n0*�m�j�nkەǰ�θ���7���\F��餫��XOc�qa�[e�:�v\��z3\�V[b���6�ӝ�a��Y�+�\fݮ��ñ��{���}s9s�Z�o�$��Á��0�ukrmg��=qŎN��ذ<e�����ם��̽tq��.���z��ky���*��T�8瓊��j�۟=gu̺���w&��s	�x��G��v����7m��-��W�A|��n��q���3��b��]�a��֧�7M���찆x{/�x�9�e��m�(��Nnx_� �g��9^��y۞�}�s�	��P��cl���ܘ�<ny�x�8ǃ��n{(�;p����y3�7d�m�e=ȧs�����ʻ��3���c#�2ʷ��ۉ��rar��es0\��.Up�rR��%�Ld;m�݌���]�|�����w�/��6ۃ�ۜ.T�q��a���������b���U��A��"�'ٲ�*
��7��I�z���[Xa��hę�	��ج�.��F����j���a�y����j��/��O�B~[�wNL�xeM�
v�y��Y���C�H�u�B�;�ĉ���Q�Aa��)2�ߔ����
`����	�`�ޫ�5wY�,i�Hʙ�}�z͢�"��Ku@�L0H'�'s��EkĨ�� �k��A��� ���#i�WME?��7��z�[ru��m�܆�69���kϬ�7=���]w/^¼0�???v??lfl�������Dw&�������7շ9U@�A��f��፷5�,M�Κ�p�ƍ����Q�b��}�9yϺ�>��Α�~�M6�xv��i�֯ײ
y5CwcN괣W��Մ�3]M�kӾ��^�L� �@̗��b�z��\д��a"�kJn!0BL���>��٠Iꂳ�����̿A���� E�uP&�ͥ�ڂ�h�������h����X�b* �����'Ĺ�꼼�8�ș��G��@�7�3ID5��	I���I.{vh�q�2ћ�	��":�f� �;�U�q���3��P�k��k3d.�V��t-��mi�x��Я1��n*WZ��Bx/�����b6�j�5��bw:�O��Κ2�!q�@����~Q�[� Z�+RѺ���/Ӱ�rw��\ٵG�mĂI�ʼ�����P��$e����`bk`�6ᦠ�E���͠(�K�ޑDv�;o��M�|.�(y������C�5r��NW�O^�ʴb��+.O�s�ۑ�D���f�h�C7v��O����i�B��$�۵D���Q��7�!&R�=Ya^̟:u�� �K�ͪ'���T`mq����A�$/jz�f���`��$&j���*� ��^S���;އ�o��E Hs��@wT0m�5��͎��H�,!�(��&�D\ݻf��g��`��[mRg��ܬ��������?C,)��P�[7\(��3��D�I��ʊݪ���W#&6zA̽�L��
��1H�qB%�	ѕ<.�0�g �O�=�B�O�wC��]Q�À���ڲUD�!��Cn���DvC$�t�;�}իCUu���3��(�c�>ɕ�.8i�,��P7{}V`5�-��ʢK����F<�I -���E^T�EӫG$0^��,C������p[��<��ه�9���:�0�^Rf�qk&���k���'f��t��{���x��j�Gn���Z�jBe(�{;�	]w�Y����m��ޭ�$>��+v�h9#��A�A�S'�M�����93.Z��=v��[K�G�1=���=[�gy-m�)�d��p��ʠA�u�$��o��s�ة4E��W짷U�@$�� ��H�5e�	O�um���Ϻ��w6I$���!n�UヹKQP��LE����1H�m�Ks^3S�I��o���n.b�[��I&�u��}TO+%TH��4وn-�t�y�G7d�5��Ă[w�^'ĉ�΢���v� ��'��P����-1U�w��� ��ޚ#��ŝ��/N�j:�I#�^��L��UY�%�Ⱥ�����7�C�i�s3�(���|C�Z��|u)��v�@���=��g]�>Q{�?U+c.�^�����~c����%��k�'�c+Ӷ�u;vPzUX��a9�<Q��2jn��%e.�c��Pr�k:0\��IN��q�e�v�\��틳�g��sc�r��9�yt�=&p`�ssC�C����0{��n�{B͎�y������m�Vz:�}\[I���۳cn�&��{I4���h���
`�[s۝Z�-�]�������ڧooZy�E�'P�V�{X�-�y�ͳ]��v�6��]�������B�֝�J-a����c7�J��q�$��{TI&gs����*��r �{4	��ekl�N$&ig]�sa��"uWE��x	!V��3��^"�VN
[q��wR{���p�0ڂ�e�	o�mm�fo:k�f�5���z��U��׉�g{��v�U0�m��4��V �s|z�c`�o�D���f�3=�4	�r;��1�ɽ�Á�&�r����U!�0�E�����rR�}�a.�'��Gd�UA36��*����?��N���/I�V��˭5�m�[:�)ݮgs6muЮ�6�;��(�c���ᶜAe�+�v������FGt�gNב��4�� ��ު��&1�4a�!2TI��rO�UV��Xet�6^�-3��;x�]m�T�f~��|���~~���S��iB�$�>�UZ��{�z���m�w��d��N�lr����g6"�x�fw��A'#��{p�<����q�ڼ$s�f5�`��5@FWe
$q����f�z�'������g�j�$���',�J
A�ل�) �����l�5\,]���s}"��9�$�����J�v�L1���Q5u�T�e�	n�u�I�����Q��XY�@��t�$��� �	[[�@�X�2B.���hA	�7h����t�Ȩ�����k��8�n��[rv[��I؎	�Ya�q=�וD�:;\��A+kz��xofU�V殨�	c9�;&hF���-1B�w�3��»=��d`$27d	[Y�^$���I¦2z��]�&16�CBd�����|T�l��g1yY>�ܽ�C��[��+�������؁p����|w�B�&��Zz�CS�j�	��B�s����y!�*q��%���q�o9 ��uP'Әl�8b
p(�U��3�֧ݢ�`���'��s��K��yyPWU���9� �u��-6`���K�Κ1d��㛔���@S��D=��j�K�E����Q��Ӻ��'�'$��3[�S�n�|�����PC�]�|>�I�چ%��u�@ �5�4I!��U��U�z��{/��'b�� ���;*��d�D��!�Ċ꾪� ����o35�N��I �9�TH$>��A��w�q94���cI��M��Zb��ޡD�^�t�$o�-j�:�"��N�MI|���>{��ۄ�B%D���Q���s%^O�vv�$>گ	9κsX.�}y���F�t�
��N?E~.�d;���zMK�g܄�����<���f���f�v��0�M����&�GN��)�d��P��ʠA�9�-��\�kMD�H�zP��{T ����dw9%��onh���F�QO�8L���A��=]u��{xm�kS�g��}�Xq`��߻���rӚM�P��+6��D��6hI�� �.Zތ���g�ͪ�Kכ4"�p�LCjl�ꌺ�$a�Y{P֎�T(_=��|r;��|o������/��J\�� �f��8�J�u�[#	���r	$�ДV�z�/���ڢI9�|vN�V
L���F糶bVԥK,t�o:Bn��I;��Ov�E�:���i:]C�fr��z&16��HBd�����ĒVWl���bQ�͆�^U��rA+��h�n�#a��ie�=�3�VN�0_6ӻ���D8�\}�Ɲ��o��׫�+����y�*P�;�F��0���W;��|�GE���?%�=z���@�Y9u�7�N���/k���r��\91����ݬb���[�ao3����e�:�<�;Q��@n׷��U֖�`�|a��qg�����@%�vͰ�C��g��ۊ�e��@%���V����O[���uڝۅ\�3\�xκ�@쯟on�����M���ѫ��z�܌����;�V��P�Ru�^θ�;1��wͺE��d���c��Ѱoc�LFn����ߟ��nq=�S�M�UH��r	$��{Cz�;��ؕ��X��f���r	g��0�!���S�@;lm��~���� _k�􂻯f� �W1B�UQ=c+7A��l���Q��bH]w�Dx�M��D����	$��H ��٠Hma�m��þ�ٵ��7�� �r�>$,�ʢA|�f5.*�U�ťb�z�ωǨ*�Re�E���}u�D��M{�빤N�1���Ϥ�}"�O�>���}O�	}��j��!��e�e��8�>9���F�Gם�8��͋�t�gu�p�����trmÆ���Qǻ���U���!��&��<�.�	�ǄJ뽪,e(�AN%��M�Ux�M� �sg��U(�]��je��{:��L[������e���%����+�'�4�{F�X����7�x���2�vgV(��T;�i���կ"�v��$�]�P�϶h�1-	��ù�]N��\���"f
H)����l�$���c.&:�O'��+:������+�A��a��n��O8OVٵ۴l�9T(�K�T	"����!��VoX>&b���$�\E��qC�7�}TI ���#0���Yg:�h�������2 ��Y}�_�8M���ݮ�u�;�rk�rm�jd=6�E"6���l<D1^�wAI��Lgx�e�׉��@���㺶#�W�2
�+�ʠ	�/mQ!�cSn2�&
�;َI�Y�D�W��
$�@|��o�?I�3�1n�lnT�x���i�)�d���M�Ux����|s�ME`�{+t0�S���)g��#d�Ԉ�z�3Z@h#�R/`j����D��l��˘~��/%�/I�3��]�[�aC��޷ݴ��)p���~`��^�����'���v��ޖ�w�-}�l�ib�6���O�9�1���g
��5�����¤�䋛�AO\�G�|
y�v-{D�[�{<V��Z�A��m��[���D��S�����sM�K�p�KMy_\��Lv������8��&�i!m�b�ThE�͸#4�uW��ٌ�;���}N�2`y������-��c9'�׵�s�ޝ�,_z�{���l�:n�u2T��ˀ��Y}�iW@�P@�����#�7ۍm(,�1�(i�Z��(i�N��Ǌ�y݋�X��o����Q2�{/�b�b
x�p_!ѯj�� �RI��w��[���F�'݀�=^�%�l��*�=MK9q��P+����t"6�{��<p�:��O�]�JbVU��<F�q�|o변��V{'��l���p��λ��g�	�p�;A����G�+���bh!�e�Wt��h�j��h�����7gLѸ6Qt�����p�y�_g��@e��|����6�2V|�`˃j:of��ష�_��=^K�~ث�����JM�E�pA���{��AJ��:�[����x�y=���.���O/[��.���Z�$��V��f� �^�7����bpj>xx2��Ξ��d2^��� 4�^��@s)�./�V���V9mj%Tx7��vwc��/Gom��`��Ǝ4-�"UJ�k��Ԩխ�ӈ�L����1W3�(�8cV�PkQ��V�ګTS-�p��֨�R�ƋKoo+��p�N3�;�l��ƪ�%���LV�T��i���V�kV�mbZ4̵1J4�
��jՍ��E\�U*�e�Z�U�eE���V��Qkm+iD��,f9(�m,h�Q����l��UAV��1qK*�h�2�1�%h���T���V[r�+cJ�f�ѺLq�U�V+�B��r�e�E����pTjTAAT�\�!m�J���f�X���Q&���TlJ��.lKh�+���DZ���,�n�� �^L����wl�����#���}�/w�R�88�%*Y�r�Ս�҂V"TQ�E�h����i�MҦ��
º�V�m���1�Ҕ�Q�iZ��L%�fEʢ��f8VQkEmDZ��1 ���I�̇#�C�UI7��n�D�n!D5��m��q�N�	=��z7nh	�u�{�f�Vi�LBִ�ܚ5{��Â�a�[� �N�$
뾪�R�nj�m	�Qd�l���A>zy�I����v�������{�ܶ���t���rwmF���q����CQ���6ݕlض����_ުi��}��� ��:���J4���W�V�
��N�#vP5`����F�3�Pر�yt�uF�0��u7�A'�y�$�.���1^F����O�=57�Z`��{��I*���x�#U���j�.���mk��u�P$E���i�)2�E�No���Y��p���^$��bI�>Y��@Cܞ�9�����T���iɫ��������.��ǿ>�I=�ע��}I۝\�'z��{�-ʞ��{�� �+���QAĂ�m�_l�ё�O��'ݝr$�U��Q�ofI���/�r���ȉ#O��3��H�pIP�b�on;s̈́z� ��T<^�^'���߿O�gL�f��5<�|WU�
$��F��+$�;Ss���y�[�I��ĝ��E�m�
�k���SУ*U���ocr	�U�m
���P ��WB+"Z��x�s:�,:���'��� ���`��딍�6E�m_���٢A1}=B�}5C�m�[�TI��f��M��N�;kr�I�oNТM��.uN�*s���	�@����^x�l(�m�Qj�*���&���7��ݾ!�!V�Р	3'�����|z���5UG!�.��)�aPe8}��vI8����}|w]D�.�Є9��k��sRקbu��G/u�l��1��qS�������6�v���Y��<.�����nb����g7Ǿ|�?8��qm�+v<bìms��7�[<��Ǥ��ct;8��y����x��f�v�<=�7l6}*��Q��Dn�s������9B��n�Z�<�+\^丽�XG7Wv}�x�8��涳�	������:��guUus�^n�\I�6}�y�ՈŸ��8�N�`�J�4�"�r�:
���<�L�]n:�jK��ۘ�Lmv�q@=�4����~��,t ��ﮨ���@��o��ݶ��Y,͙�� �}��^���Â�0�C�3S�O���d	�C9��v�H�O���s�.���1B����FZj![-�Ӈ5�yTI'z��6rF���>{�<��$��;U�	��bwL�vL$� �Bb��fu�؝���w2kĂe�$��i�1����r��	�y[U�c}��YnP;��IYהu��"B�"�@�-��O���A�+����/
t1+D��5�I��=ls�;F�/dѶ]ױ�^��u�.H�d!���5(�"����z��A��bI�+��k���HZ]i�mUF��n��)���ЄO�}�4
�����Ά��Y��:�����������j�����7�a���KuUOLo[��y�%4x�A���{�,4e��C^S8^�|��w�3��+���op�*Q��}��w����2T;���b��|�\��A`���j0�L0���υ���M��¤�
��Xg߿}���%eH(�|���S�z�Q _�G� 
>{����R��3�{�q�`V�]؅�Ã��$�#��fȲ>C:7���7���,�%ed��}���%H(Q%as�~���AaхIbo�y�Τ����pU�����G�6��}�!���0�nN!1B��G�>��@�g�"��$;��!�ڬ����<���|B�����y�
q���L���ngFJ�2T*��}��tO#�W:~��=#�$���n�����\�a�=�U�i��֋%�u�/��w���ۿ߿k��kZt�Y[�4��{��oa� ���{��72u��@��{ϸu _�G�=�Ǻ#���|�n�π�*A����=��ۇ^�+u����r9�H�� u;g;��N��d���߻�~����ߤ������R
V>��܇Xu�aXT���϶u'P��@�z6'�Q;�g���f}�!�u0�M�:�(�|#��@�g�&�}�=�ăҐ�`W϶��ӯ�D!?'j>v�f�j���9r5�p�Ž�m�i۸2ڹa���y����1�6�p�~��g%/�;���s��)�J�YS=�ngY++%B�{�>��:$�/|���u��bxY�|���@��X�j�Y��&��(�a�~����u��T
���yϸu�+�X|��L�	��� ʎ�;4xx%������g�"s��LÃ�.'�IG�~��ΧP+(�YY+�>�{82T3[�q��~矽��D��'=��rH,:0�(���=�ԝ��2��}�ϽD" ]�����V��
(&��T��r\� �+:%�������J��q2s�N��a�~�	�"�&>@��fw�0;�)h��}��)JB�0+�>�{��
����sߓZ�����|��é�d�Q}���Ԃ��q�iÆ�	S�φ�{>ِ(G��H��������3�u�ߛ�g�:�P*T9��é��k�|��o~�!�;����v^T�q� ������u�2�� u:$�}�͝N�VX�YA�������J�T(��}����z��熟��H�W��"�:!Y++%e|��orq*��9ni0�M��t P!��$�A�{�~�����R
���6s���!R~���� T��&s߼�:�\�s����0��6�����
�8u�u��ì�pGs}�\�r5M��f�xz,����;>�����v�r/����������:ײm�2Tyϼ��;#�����p\&%�u�g�ς5W�0�B��V���Ό�&������g~�������T9��vq�X5 �o߷���B����{���^�+�:���pX�";�d7@MC%.�k�&l���;%���k�e9mۛ�׷\+�����G?�u��h�g�6�O���6u:�YY++%~���g*AH,3�����a_�u[���+���M��(�}�#��VW����'"T=�����Lֆ��tp�bV���w0:ԇ�ֻϽ��ny��'$�7�i�_ ȁG�z�� )ȁR��3�}��ԂΌ����HN����F�0x�#�e��WY�ֱ5��y0�a_}��I�G�>Y�υ�H�DuGْ�k�w�����ȕ�F�,k���{���)B�9��nz��9����i�$�dY��6E�=W5���>�2VQ������(q%B�+
g<��!�VaRT׿}ݝI�<�y�|g���d�ʐ\��opN����济�u��� pJ�<�߷0:ԅ <��V����~�ڕI����|<+Fu�<��)�
� V�>�p�:�YY*�����Aa�;������?�Z�a?���r�^�^~�.U�[ۗR�鍺8�,T��[�(�kI�}r��ƌv�7N�]%��4C����;o ����[�Tn�2z�f8x�t�h硺y�U�0w!��K%��v�Վ�;go[>���]�cI<�2�n=3[pn{q�pt��UwV��[��[ʰKh��f�.�c��4��w�k&�9�W�� �dר���9�v�kx��	��w�����8n�\�i����e�{Tm�`{�5��ؐ�]u����`�YН{��S=G\G%����.x�a������,|���'|y��E��.F�࿼,�~��F����*J�IP�3�~�gFu���Q*�����A+΋Ͻ����`x5��9���i����>�p��i}�*[N(p��E믾�E� G���G��S�;W^��;�A��ɑ��DT*J�9��70�aXQ�@}��"��'ް|���u�ވL9_��\��(|��\����Yn�@�J��}��^���}����� ����s����~�� ��eL�~�p�:� �k߾��!ԕ��q�CpC��S�υ{>ِ����s�{~�
O��a���͝gY(2�T�^��xu���Z��_7�۟ ԉ�C��&�<<�t�Q��s���rj�Lqu�N��}�:�++%e����>���k;����[������"Jÿ����u�ac
�����:��T��FW�}��'" Q-^����h�QO�3Dz!��v|l�ݭp�wMR�j��;<<Sぐ�5˸����߰��u[�&S>4��y�l:��cR����9Ґ����_}�@	~��+���QyW>}`�YY*���l��+�?}{\�5�X�Ys5�u ��>���¤�T����y�{gnNBpʣ��0���\�9=M��sY���T}�=�)��~�}�z�Bd�4�^���(+�yU�>���ǻ��އ�9��͟�%e@�Ty�=�Ă��R��{���� �ldC��_9�
#����R�Ŵ��˧Z�@�q'|��ݝN�VQ����2(y�D�<����ݮ�nj߾ּ���a�0�_o�vq �u����kﷹ8D��^�o��kZkb����|2�ߤL���"ֽ�� jB���~���H[HV�+O����8 T��&s��:�k���m���߉��Ɍ�d�Q���Ԃó�,�2��pC��U���'��O�#Ȁ�����dX>��!���ә*������\�{�@蕁Z��_w���KH)���{�u����?��{��.D�́,��A���E�0�ݞ��Z�=k-=ȴ�E�����{�nh.^o�ݿ���>�i�.����$�w��:�@������������,IXXg>��C�:0�<�^��C���;'Ss���N�Y(��FW�y��'�P��_sW.�WF�Wg@�V�>�����R�54���nOO�@�9�d�Ї�AS�s�w�
q�Ͼ�p�:2W��ȁ�_H��Ӏv�}#��>_�wI�Ä���υ�n��@�����T��9��2u��P0��ߦ:`@'��-���e�8���V��1�ڰ��/&��9<���������c����0�	�r{��O&p.�{"����.��*�� x]n��� ���Q�������l)
�9����
�۫�g.���N�7i�w��E�yȅ��ZcT� Q��y }�\���q��*J�~����+
|@��W�,�|�w�N<������y#7�L��� !ykD$[d��L�Ԃ��>����� �)h��}���y���c����>� )��+��}�8�Y�J�����8�R#�o��-�cv'��"���dǔ'ِ��n�Qά.=z�m��ʰ]ӥ��@l��|�����Ӭֱ5��~��|¿{���q�H)(�a���:3����T}�>�����S�Vۢ�~���8~��� �Xg;��ïFy�����j�i��7��I���u ������~��s~���'_�������RT(���s�y�u�F�T�M{�>�ԝ�T���M���>�J��^orx���i�M�Xm�0"�x��mvH=H)
Z�����ii
�����'T38�.���0���G>��ì��YY*���l��+
�~�`��i��!ׅ����d
��o�����r�È��?��a�N��J�f����bVi�}�π�����x�Gݛ����aM���T��q�S�G��A�������nXǏ�e��m�wq݈�ϫ^wM��s�;���o���C�����<	��&"F4��Ex�'}��6u:�R+%}����p?x�����$�)��{�!��+
0�,M~��l�N�VJ��Y_���z�Dי��zsԾ����[^�;m��-�6v/dW�V�t�9�F�]�F�׬l�[�0歈A&�BL|4�>!�7��XjB����l�e!iHV�^�謁"� ";켰v��X ����{�é�*��{��u%a��L��!�D��dx�L����!R_������l.���?3��eH(����@�T���_����"C��<�����\��)��<ϧ���7����j�i��9�ԙ���gS�eJ���{��*ABĕ�v��0�_�=���a� ��T�L��{������A���~��(�D��&�0�N��#���]o��������R
5�{�����!Z���}�@S��@��k�����k��;�v���gY*>u�G��9��a4�MDC�>�F����q�ID*Aa����:β~�|���R���L=�Y h!���@B`V��{��H)��_wϷ�|$x7�-�q�.�S���	��ە*n���vv�[.���gn2���}�A���|�9Yy>�]�K�2�Z.:ɹ�9���
��bxP�6��׻��ƣ[{������ፗ^zow.j��s��L�2� ��m�k�\�&��N`�>9�ܺ�����ʳ��N7�tf�ð��.�1BH�}������6�{Ur��;7�q�{f�~垂�,�[œ.Wl`�*;�� Eu�/�zs��;t�u���;j��sZ��4,�"1�YO�
���y���SO�ӫ�H��~$t����OC79Y�A�q;ݴh�V��Ң88�'���΋�Ays;	������C;�o��
�>s|/�͂��p�k��XY�ҰƧ��I���^�c�%��Ui�Roq-B[1��Ǉ��{�/9#�rw��:n����6��R\��V �z[�����4��a{�vl#�S�]�n����n��c؆L� ���o�xo�x��|#��K�v��oq���<�<�9��N�#n�-Jăn��ɺ57��v:�.���Uq����t٨�Q�q�?BVy��3|�@w��!])����_w�юס�
��Tɯ{�7�;;���р��p�Nq�:P*�f�=[A^o�����j'=����^I�2i�M��;WY���#(�+̥�+�}Z5����~�)*uG�k�k�3��JwiO�8��pOb��� �{��Ŏ�/��Z{�l2���Ƀa���7-Qp�������s����a�F�[1�Z5F«j[h�TZ2���h�[DZ5)m����j��5sʖ�b�J"6��ˊ#�UYB��*6յ���
�B�H�-l�n%B�u����Zж�h�m�ٙb���G2�b�PH����i�)R�%e����-LF��V�KQ�­ZQƦ4QV�5j*84h��.�b��ZS-U�TT��ڋ�Fۘ���X�%B�TU�c5luu�hڵ+s*�+B����h��S-�J�P�Z��J�[n8��c��%r�0K*�kk��ֵ��F64��Q��iX�%�f4�Q���-AR�Z�V�WZe2�����m��i\��.a���V�Y�" ��m�LZ�e�(�,������T�QF�s�쉻`��x�#��6����6�DG��m�%�[[J�Z�c[Z9�\�Q��S��bTUT.���(��]"�D����b��Lb	��R&YQb��9Kj�[nZ�2�W-4�SH�kU��]�{o;v���؞u���x?8K�����wN��ȭɬ:{W�ph<5n�۳��r˰;P팼o[4O)O���63��2��[���smt��+���\{;qk:�v:1��e�p����̓�ۆBr뎅V�c���\��j��Pm�!X5r��CMʪnLfxr=��oLnT<�ɱ��:ژ�p�U��.�8�I�qی��ݏV���1��'��z�`�ؖ�J�;LQ[�_G6�{���}1�[jr�-�N۶wiF��b4f;�xz�6P��wHr=nMB6�qX-���<��m�/B\�8�o>{[�c��Y����6џ]�:�k
v��
��y�Gn�"ƍ��QvkF˞s��܉Y�pю}
�Z���n{��s�F�du[X��{s,6�/[���1t+���5�a̻r��8,���H\u���By�93v�n���:����J	�d;!:{{��c��cn�Z4�zr<v�	��V�K�W;���S���뵹��ŶNlM��mv���[�\[n��	�D����ț�9G���z��o`�z�\�<�n����:��p�u��<nk%4��p6.��F(�t�܁<�[x�����V�i�ӆxz�Rn�q�����3қ�Kɍ�3p=���-�Z��'M�5N.��qc���ǝ��d�-ח���;c�r�#��<n��gP�:�w]1Sn�a����k��]L�̈́G�ۍ�׸ePB�N�v��WK�i�8�n����g��guIn�Q��=�8�֟(�������ۈ�k<˅��d�Z^Nm��qEm`�*�ۊv�x穤w>]��u�ݮ5n��;km�ҌU;gŎ���6x[&ܹ	:�g��;D��'��SNV�nm����^�qr�q�+��#=�n�.ø�D�x<u���-�`��u�y���壎�qf[���j�s�H��^5�t1�Nm���qm����F2�H�n#�ʭ�=�
p�^01���;�=���-$p�Sw����{�[��j���r�4�1��4��k]'5ś�s�o;2�ٞ2܋z�t���T� �뎱�=��eW,��/a��6&�֋��^�[u94�����ƍur�94K"Ii�uÓ���;9����b�أl�y��p�2t��.�Q�)X-��8ݻA���E�z6��%���n�9�r��9���&�zՀx����|M�p��t:��.nۚ�[��8zv���ӳl&dy�a��jgum�\�ˢ�����/'�������	=��<���@��%ed������d�X��RV_wϹ����5�����G���ܑdz���2��=�{�������r��h��G����l=z��R�u��]<��7�NȬ�	yQ����U�� T�a�wϷ3�%ed�-��ϧ�Ӹ����2> `#��pq�L���D��g¼|��f@�D��ID+���nH(J�˾o<�e�_wÈJ��`X��>�{��H6���>�����_9~ˆ��>a�d ���Gd�3 ��`|��YY+��{9*%H,(g���C�:0�,aRQ3�~�Τ�����������R}���'"T��o<��UsN�n9�8%a��l;��� #��U��������>��Zw�󜀧*Aa���73����Ȁ���Ȳ�<��y5�շ��Q������{���������Jcv;y����&69wU�Ft����������ѭ*��w���0�y߷��
��*J�a�w�72te@�P,�}��:��+�yt�m���vb�c>
55�π$xx%��{��Y� �줠�ƒ�᨟)ȓ�}�͝H,�%g6g~��s=�o��>n�&��sdv�خ����Y��8"��5��P��}Wݎ�-hi��Z��E�X���#rR���pw���x�Lu߼�βT,IP�%aa���y��aXQ�IS>���:�������~��_��.���D�"�@�ێ[tp�bV����`Xԅ� w}r*�	yQ�󍿡譇�]}��s~@�=��}�|�8��J��P��wgP�IXzk=�iֵ�Ђ�T�3�@�#����Z�w>UXn��Ow�R
MVw�|��Τ
%@���ݜ@蕁cXk��k��Og�~������_���	/��υ����|��.�ZM-3p8�wϼ���@� �s�}��d�<?w���Ni�^=&!�IX^o��raхaF%?{�vu'P��ed�es�}�9@��ѯDMLyD(I��$0�b�On�u��u���6᛹-�Lv���իk�&������ë\֨�-�Ă���a�z��R�3�}��t�-�![��}�����߿~�y���m�'�w�ۇY��YY*�g�{ݝC�%aC��~�qti�u����:ã
�����$�&w�]����9͝gY,e@�P3�y�� u+��F�����L��#�����RdIg��2{~�
#����4���%!����@�_vl�"�FJ��_y������%Bĕ�<\�}���&v�;�3ZmVD��</=���p�o��Ֆ��y@��V肩G"º��T�sֿ=��ok�<W�18���l�7y� �  �����?���*J�����ԝ�VKR���jND���;�h�F���F�  �|3���g>�<)|Ql���II-����s�����`V������q�@��3�����$xr���Fw�?~ܜ���s.\�V����I?$�;��	�<��sӚM�ó���y�:�X�+_���@�� Ґ�3����Ă���g�����Wo���C�9�i�61��M�vk��;f���� ��m�!��Q;��PM��B>�G�z+�}���++%|ߞ����*J��+�w�y�������{���'�g�~�ΤN�����}�@����_����h��/@�J�7�߶z��#�8]j%�?
� cʹ���Zy���'*Q��s��:βVVJ��ߍ�}�����߶uVw�y%�Z-�P����&�s�G�B��B��}���JʐP>�����!=-�Ѥ~! �>z~�P9�A����s��:�`V�;��P���_�\$����NM����,s�5�~�׀Vt*A{�<����*J�IXg=��Ì:0�_o߶q%�=4��/�,�U��y&�H��˥ؽ{E��o�oo;w�5A����1��]��y^��_T|!�{�E������������I$��6��R��s�rr&�)��s���i�2�����a�����v=`Q�h�~�l�Aϩ*Y�%�D���x}�~�P 
������7������D7���E��O���G�-�ۄ�8&��n��^��*��\�Ƌ�.�2q���[��xҫX��������Z�a���U�CL>W�g�l9i%�T��9�nH(�P,����@B>��w{s�|��8�g�Ph�e!hXg=��ïX����f:�ZM-3p8�g?~�gR:2Vg��~}]~�k�]g�:�3߶q�HQ%B��.s���a�°��ISz�߶u'D*Ad����_��瓮��~ܞ	�����Ai('�A P#���a�AHR�7���g:R��
�yw�9���ª��^O��@�!3��{�u�d���
!�}��:�`���<���:4�5��5�q�XW����s�Sw3���x=�������,�ϼ�*�o_��g:��F�+_7�}�޷���y)l9��wp�сW����a���7iĝ������
��YA���>�gM!�k���Y����%ag����aхH),M��}�ԝB�Q�����y�ۓ��.��O��m;�W�/謗�թ����,f��#b(ōL�'Pε�4�[����򛾻FxnT�ͼD��)·�H����h>���_�<<=�#�ۆ'��gn�ܻٞ���%ظ��m�k�8��n���n���Ϟ�����0�ܷ��㵢�.P��q��,y컙s�<Ʈ�y�t({d.Lv5�#Ҩ�:.���uv��2��z�ۭqMۃ#Z*����W]�.�;�u"#�ݞ���5��%�\���v�=w���f73G`��@�dI��6x]�ޱ���K�ҍ�[i5e��r]��a�΅ŷ]i�v�#�nJyN���h���((e�)$��d��|:�
$�mz�߶s�H[HT�������E#+4�F�:m�<���O����7������bמ{��tIXp�؊���8h�>�Q�G�>��|^ "=57Y�[�6t>�����}+*�]�����X���ہɪA���a�=�/|�|����8���z�~��c���44�@�v$�߻�ΧD
���d���>���HyG�3�+���r�������aXQ�ID޽�ݝI�
�A� N�}�� 
�s࠴���T �(�|#~��;wA��:ޝ��0�<	 t��l�A�HT���kϹ
q��}>}�9�vx_{���� <���Ăýם|�GF�Zu�s\�Xu�{��4��T�B��w�2g3��s������8��%`X5 ��=�p9�A����~�p��0+��~��������M��b���I�{R���s՗m���eW��Ӕ��j۵�<�_����r\��f����w}�8�Y�%H/�Ͼ��M!D�
���{�ۇv0G�kwl���*Ϣ���<���r,�Y�VVJ���>ܜM Y������uq��:��+�����X5!2><B����TG��m�J�nD&)�i���p��"���ˋ�d����(������1jk���f>�bcm^&�x\���_.e�k������ �ۗ"�)JB��Z{�}� br T��&s����%ed�{����v~�߶q������Κ�f��j��4Ì+���0�J!R��y���%" D" y���D�I�돴q |B>k�s=�p1 �-��~�p�g�"���]�2J^Ȳ=�d�N�w[��\�����d���>��M!A%B��3���p��+
0�y%��H�<���ΏR��������FW�s߷'Hw�o/��V�]\�1�V������Z���o^���t���{ζ�}������s���9*Q�����ngFJ�2T�	{�H���|&ɓs���]1��;񴈺��z�f��g:S���0n��u�OPi��@�|�[��D�%��>�<	�Z�p*AI��s�{��:�YR
�Ͼ���+�[��w���bAs����y���Xg;�ۇ���t¹�335�� m9�翾���YFD}�W[�>���C���G�r,�A*IXY�����Xu�aXT�7�>�E���y#�]>�L��}P��N�>�ۓ�1�r���sN�-��@蕇����G�!K@޼��臂#�����A�,2��.�\p��R��[�
�y�.�xD{���J�y��}yEw-L?:6z�+����7�gڡ#�9#E��ָ�c��ïr�x*AO�YD�{���Ԃ�P5�}�E8�#�[�.i�*�g�G��YԽ�%O�G�#��
�͞Fu��T
	P.����D�
Ԃ�ϵ��_���u��;��A���fo��͟ ��X?b�"Nd�#�:�������؁R
A|��gz//
�pt$�����3�y���raхaF%M�߽�Ԃ�Y���;??��" �\l[���(�~pX[�m�m���Mr�{Q�;��ܜg��Nȑ��96�չB�PP�| �>!�̟`tjA@���ݜ�H[HV�|������}�� Q������Y��%eJ����8�D���|��ѥ֝f\�!��+��_nI�*O~��ոW��p|��}g�@��P)����@蕁F�(5�k���x����[���G��]O�>~����i�A�P�(�$W�����,��2VQ����}��ɈQ%B�y��c�x>��w���O�|�I(���~�ԝB�VVJ��������@�����X�dx�}�|�~���>��H(��y��)
�Z0+O��rH)�L���u��
64�BGꢑ����q��&eN�[u�=��:_�'�D������>���I�w��1^��c��xJ'y�px�����2�B�4��J��}���:�RV�;��5[���tR�H/߿��a��Q
��Xg>��Ό�<i��}���� B �ꮅ���
Ԃ�����p�AH,3����Ǳ������X���q��q�P�	Ɨ�f�뫬u�4w*��uq�����v�q7U���������1�:�Z�L��?s��:�� ����w��%H,3�����aX~����Wp���~�ĞT��`���5���b��y~)�-�5r�ى|�w a��Dxs��D}� t���!iHT�����y��T�{�ۇY�J�2T5���y��[�߿�pכ#H�>�U���ˈY�C�:0�w�{�'"%B��w߶u�H)�g��ݼ��>�^����Vk��~k���e �B����u�`V�<�T�c�r��@.~�$Q�TU�_Tt������;���8���s߽�:�Xu�@=�H�=�����	u?���O��>G�G������D�<�a6�Rh��D�?w��n`t�P7�}�g;�J-����U9�È�''���F�!>B+s�[��h��.�C�W[>���R�8�޿q�����(�L~�9w��#0�m�<Έ#M����F�z"��C5nS#�܋��WR݇3s����w�����n�K3g&�<�D�9��\��Wi��{��r��:�g{mp����q�-:�ô�͏]o'L���1u��j���W\�Ӱ3�Y~��g�om�mcq�$��>n3u�[�X���3=a�vӽ��U�#�{�xg�:��<��{0�� w=�r���:����\9u�y�dM�+���꣰���3m�.w��x��"�i/%� =���㧜��;���;�N���ۈ��],�g���w���?�i�(�oFO�� ��ʢ$��ޡe���9z�ތ�%M�M2�ˍPa���U�o�P*g��7�ٵN�(���%N�U��w��7Vd�I�Y�h��ei&J5
�Vm�
>'���٢H|���WUYTϨ)��I!��U}U9�"b	p�DC��4�:L��8�̷��3U�(��ݪ$����DRX���ٺ�(����'Ǭ���
!BhÚ���N��8q)سT��	.�輮�����j9����?�����S��`�d0sg�;=�.��s��������;.���߿Oϻ]���#~���Q$ݮ�^ ��|E���1�!G���
����w��Fg�Y�<$�e��
'�o�$"}��lM��A��pp����:��~k5�~�n���i�[8K�g[;�'<��
ξ-������̘�-񈡱�Z�M*]~ {�xT�ӳ���� �������w�ܪ�㮴��z���L��U']�D�2r:@@��4�du�3��Q ����L�$� �4I!j>�su��V��gz�`�[U�@�#�=2H$)�ꚭ��T��$__u
Sz�D.��u@Ө�@�9}1e+�֘��3t(m�l�|T���*ר+�a�Bd(����g�n:zعwfK�n��[Z��[Wv�7���(�	��ܾʢA �����G���W�*�8��dV\���]РO����Dj�%��NI�6n�:�D���
[7����m�q�O�
kz��zb���V�#�AئJI�bA@��D�5�^�I�3���V�u�3]lmE����K��Y� О�X{)�d9�^	+kT� �j��؍YXq�$�Q)���#;�EʇYn-~��ڔ@�\�����aǅA�j��m��Y��I��_Y��w��i�璘?�lHs|����xP�Q��^���(]it��d�m�rɧ���:�a�w�.�N$㷪Ƚ�!{��jX:�"��^��Nx{Y�彞M�{�&\�t��}�3�vg�����t{�y�Q�۩�7˓�H~��bk�gS-���n�~�l�&4v,/���y�=��`ζ=\<!<V�04���j�<��>�0�^ԫ>|����dS�'z�z�3c5��ͷ�-�Z��������%� �k����;�v�|���(H�ש�_v�TLvw�y������oA��癅-|��>�O7x��su�A�k��'~$?Ű������Lx9q;܏�{�\��������8��x�,C>���T�|6��:?=R�����t,'��`Y�Qp�>�g��K|�Sv��I��;�z�2�W��P�.���8�0r`����c�ޙ����
zE;4/4�\ø�Lx������e�A�v�ݴ%��b�~��᧰��I��<ٹfƴ?o�X�<)8e��,�]�&A���C`~ޝ��w0�^�w��7/��^���"�v��Py���O���E��t�{�>a�Ung{���7�����N�QR�����~8EA���'�qt���W����;�7�,.��O3^y��~�cM3����Z` �o�Ǉ(|]g���ɴ�=���iIQ��8�2���J���X�#1Pm�m�i�W-*���UlA�5����D��Z�(,Z��U��
\�2Q*��J��FUAb2,��G,�-��UQA5prж�EM0�d����-�LX�"e���1̭[�\�dE��ZQ��Z�E��&R��b�E���SKn��h�.��j�em�,�\T���R�DmlmX6R�l�l�
�
[[M[��iF�,�U�T]5ŴTUh�e���k�[L���eB��bbE��iAm�¤Z���R���[K��Z�E�j#m���0�R�q�KE4�-F �Z���-
Zֶ�jR�U�mQ�q��G-��#W2\aEiEQR��`���0��6�Emm"�V�)Q��nZ�X
��[b**�e��kU�����(|F����T��A��1ɘ�I�DN��ڪ0��Ӷ�����@"	%O_P�O>�}8y5�5'����t�4 ���PH�{�5�<x0}�춘���r�L�'=9c ��3!Wv[gR.�vr��K��TƎ��u��P»l��W��b�����"�x,�]���4�"����7�۞nD K�sŀ��ݎ�`{ՙ��;�tt4ud�I 
^�f`.��B�HI�.��:��/	��xx����y��9 @�7�πUݖ����7��w�&Y,4�q&�Aw�գ �*��i����o-�Q��5 �u���3�
��o�TI��H
������ج��Ӿ�}�+�u��Q��L��O?\-��X���'vn	����e���\��f9��ۻɸQ��87���}3UѮ�J9�Nv+�H�ƹׯ����u�LS���߼<�O�u�wi+���pl�����l���K'#��V���a��ݾ��πA
�r�d���dgyT'���}���"�9v뒹/ms���J�zD֊a�����a�ь���?>��ٌ=9FK�/q� {r�dA�m���4{^��qW[�~�̈��V�7�7�J1n 5iI--�������?X�ώ�_�Z���� �W�.��#o��� �Ⱦ�N�/yO��I���Y�`��
(�vг;���$ m��r ����V��zA���"�>�m� >F�GUKD�ń�E�Jd�R���-�
yk<�#�@|
���a�DokX�� �;�#2XM�Ӻ_ �|��4��$�R����4�:��t�S����e4�r���l �O2!��;�L's�#Ђ<��ks�I�<� ���*���^d�U2�,�Za��H�"�O�2vݍWK7��Y<�.���1�d�9b�ș�՟��
̜�m��C���==�������9�)v2c�(�p��cj�)����qmrz�;�5����)�q��[�S�A>®NcU�[�����'�ۻv���;���v�M���0(e+3��集8A7==�'Z���V���{SƻA�۩�ŭ�z�:��E�(x��������r�*�;^��stdOn6ݘ3X�jP�=����t�v`wB�q�iƞݭ��^�3�̡���9�˄��y��I| z��p� 'Yݙ� *�{j�ˤЇt�P�W�At�:&�c��!��H�[���!�{K�bb}9�[��I7{o��e��ကN��2#>��P�S�nd����ڦ���I�346���& �����>����}wן �={�q���3 H���`1
!�5�.�*�1h��]�Y��3w�p�/;�3� �!�W�EQܲN���TZ%]��h�1Q-��1` 
{��,/�z��ɀ.���`��7� ��eB�crwj��%��דM@���
�nxc���9{�ƭH�=W)j^m��EJů���O�y�	)T���f��`	y�x��
'���-�^u�<��dDCR�{3Th�)�J�*D)�S٭����|*�������{:���B-c�q���i��n�|�gI�!m��=�fT�r4VlYG;x^MGms^d/\��0rR�gfM��I%�ݾ��b�߿f`)���d鮬�T<�q�-�^���r�"0�(����n�3�"�O�-��������ݍw�`�۹� ��w9�t�*Q2[�Q2�9��Ҙw�}���Q3sp��D���"��;"�#�T\x���a'�8��h��'�I�m0@�O?�ߥ1�f�Ty�>��{3 B��o�@G���R8���~�L]�����qBƀ��N��C�n���7e�Һ��O,�^�z7��}���ѭ.[o����ݹ�  Sݖ� >�\�9�.{s��z7u��Ă"��Q{��&)T���|v�@?GV�#0���ǟa�}v����C�x�"�c��oy��]�&�L�T��P�m!Oo�`�=G��G� E��3�V,35U`��N��T���9�7ή�LGY��A�q����EK�Q��K��x&''crc�p�4�PDDj7�~���{��r�0��HG��B�^H�_t��ɕ�"!��D�T�n��Np�q{����{�m&D %�k���S�ݙ1�Fs;�ñ{��nj��w�!ɂ��Q2��d�}�v��q,vaА�un;h�=G��C}�ّj`sWWn��k#YpB�} YL�^�k��.�;xaS=ub�^^�R�7n���u~}�������S��^y�p���;�� �gvfW��%׷%͚���;�`g��@�\�T�$�D9fnv�,�E�1�'ʻ��*���>�, '�ݙ� ���/mF-��u�"MjT��H��F��jN��	��<� �7�gin�K'^W+����HF_u�$�h��2�R��"$pG�^�|�r]޵4�'7� ����@ ����� �{Ͻs��^ܘ��W��Hs˿9������g���=�������1.>����e�0�}�P��Pʇ�}/v^0���{��K|sٳ�b��z�!Y��? =�����$���mPkﮎ҉�&f	-�^��� L>ۨqs�wsQ+����H��u�� '3ݙ� 	f��/`̚�}R羈_�'�s*�ܘ���Ԝ5���<k`�۳����3�<�C�_ٛ��d���چ���J�iЀ	��x���s"'��w�5Um��
��|{�J� S����#��iV��Cq>f?�d2NT۠�˹Ok;��8���7�{�l As��u�]�L���4���\I��f���v�, ��ޫ` ��ۍ�V^tGv�)�_dZI%��$��y�;:,�PXM�ג�]����� ������#k�����C�]o	9[��	8����%����m���Dz�sN����z^y:�P_�3"0MwSa ���c����ܔb����+t��#�>��ɉ�"��D��t,Q�	�9<] /�D]���X&ľ�Xa�7p/AqQ�QqdnD-��{��{�&��)A-���c�qv��h�/.��]��W#�c��3�:u��8�YA�On�$v�G�>�Pr0�s�l�սy�eÁ���v�c����D��x�\��l���em�H�q�v�c<\g�3��6t�R�h���qqY�7d���Z��%��mh��c���k����Osn�h��;���u`M��;'1��v�c���\E�Z'4)�C�V⣥��L�ޏW�p�q�<�������J
�f`�����X �ݫ`  K�=�Z7�}�����tmU�u�mݤ�E��5��W@(�LB�p�4���}s��v�ǽ���g+�ϰ @*�u�h"z�y���'�=F��: ��=�I�D4�+@E!��3��[ "+zy��� վ�֢�f����> "��V�{���^Ns(�T������,���=��/ݲ�;� ��m � S��c���fOB�N��M��)��H�&b�b�BO��:Ӑ"&�y��Ț^��W;����c�"Nt�"o{�"*���2:fzfDn����m@�ʈ��H�Z7����v�w(������`A��a<l$�G{A�D�%�ަ�@D�Ӷ0 �����Kq��w�kb5�鿂 	ݝd5�Vt�J
@����gf}��w�{�྽8���{}��2|gO@|>�]�I��?��.X��\������ċ#�������������W���'� �	�팟�"RJ7�R�$J�ߺ� �.uv�t��Э��� �v�b�)�f���������{��� *.S���������|Nt�"M�t�	#�CH´R��="�����������=��>i�� ���3 �<��Na��(�H��7 ����i�ɨ���v�֐	=s����s��q�8��Ir띱����&�3�5�F���}�����t�puй���/A��3�>�x��ی��qG:�gunI����0XM���Y�Uy�����9ix��{FN�ٶ�}b��ȂI�]}��	/���R�46�q~mPlG��Ά'%��jrD߽����/�� ��F����3z.����.P��;������/����A��ޥ$C�-�����)����{"㘴%"���36L��Xx�2��{^�5rq�˕,�9���x�YV�	$�����0��/�TT��b�)�f������k�HWuT>�z�ɻ��B| ^��,"}��	���=ٱ���	��bF�Hn'��3��$�%{��kI�U�^�50=g���0�H�^�_Q ����E���c�Ys��㾚��{x�C���dӝ�#<W��t�9{s���o;.���v�jh?&YQ��o3����\��0� =]\Ƃ=Y��S��N{��w�^YJ������"54�i�G.��j=�c�o>� �릀 �t�rA�v�{ݵ��<���pcEy�ʥS
��F΍�7�� =^�i�����W�H�~u7�s^���� �z�y���s1��(� �$m"w;�!2���~���U��Ln��4/kX�/=͍�Գ��9��6��c�k�O3a'�J�r�;Ǣ�o"*\��~��w�4ނ9^���c=Q11{Ul'4����\�?{������$�����Lul�(RT�46��i�	~�������{1t�F��逐���jH M�u݄���3=ފ�>Ma�Bed8��6q�1vx#�(=�0��tcە.��u�N�2t����qB&�I3��\{r�� ����D@$�=ٙ�gzU�r��.�^��S�6� �{��O�D"���	-�^{9� oU�������[ܝ�^�Hջ\�� ��ݙ� �|~p�n����IF
��h��BT��z5�'� ���a/�5B�2�}�9t�.oz��� V��jH ��vf +N�7��~jA�C��f.WDl�7�Dǒ���D��v�o�D�:z�& CSe�z�S.�y���4�T��$l�g{1` �z�-��w��B�N#WnV��	����������G�p��;��m���k2rgM�7=�L|_H\����V�yԜe����W��rW��H���S��D/}��W;j�?\��<����4|:+��<��]�=���{<�l�&V�H���H�}�n��^���`ޠ�g�i�0�t�4��A�sB���>���� @oӚ����O�}q��/�b���W�6a^J�����ڧ��2!�O^�HF�7�E�A#v� �����Xs�2�~���{l^9�\�K}=&������}��o(�G�`���bt<�]�
���[��7�h�Gm�fw���Cۃ�s�Kf�xy��-��"�Á9��GX��O"��s�U-��ܪ0�m�������8�p�E���у����p�UTn���RVQֿRϱR7:Լ=�=�y�o��B�	y�b}�,�-o����o��2�'L���1���0`��n��\����G�����K��)s�����=w�+ڝ�b�݌&2�Ľ�]��ٞ���d�v�y%�Гh�DA`}{�e	x���^6�c�*����xH����|5qt��1j]|^��w�)(�5�9O����} ���L{4{��]+�=�MD��ӗZ8����_Ւ�w��x�ף�oia6o���Vs�N9����1�3=�M�=������p��x��+��d�M��2�P.)��eN�� �U�|�8|	>���E�%W�$z��u���cΏ^>:/�{��&��g+���w�`���L��&���1�$�ԥ��&Z�mQ��Ւ��Yr��	fe�b����H��T1�1�h�X�Ķ�R�h�1LjAV+�ci�CTR��TATU�*�T���آ�U
�d,T�b���Lʦ5Q��E�(��,�\m����QX�.R�-YBڵ��F�P��V��1�(�T�-�mml�*��ckJ����-ul�b�Q��YQV6�H�����ʍ��U*��ImDD���b�t� 	j�r�qR�㌖�D*Z���iKFڕ����#DU�E��m�u��E%��F�
�MZ��X�*V(,�m��Ԫ���ZZ-�������VՊE�l�+�m��e��-�E*,�U�b��+*�*b�m"ږVڊ"�)�Tl�*iDX�(�KeF%�R��\eb���(���-,*-J��E�����DQ�KQ��e��9�V����dm��J���V��TU����/߆=�v#��%�aw����9��y-�+X��֜P��d�㵼��r�s�Ľ�x{��n*��<���3���V�H���Y�˹���ᛛs��z��Mq�w[{.�Ù���m�{po��m�«��hN�N�I�q�Ll�ڭk��d�=<�%�*o!���粗לn;l����q��;�1�Ur�sZ���xֵ�;L	٬�]��+�u�4�wM�˴v�4�G7H�j;nf��m��ܑ��)���a;k�n�:�6����&���vY�l��B�ٻ�e ����W��#m��H���q����v騎m	WD�����uc��vW!F�=N;q�w3t��g�ctk�\�!y�`��T���"��=�n��ێ��������ӛH][e���1�:$w���s���F�ۋ�͎W�����Q�/CZ.1s�NK��Y��[���ac=r��!�+ŭ�m��a��2�zǙ�=v�s�ێa���[�{'ps����ے�<�������7�Ļ���	q�Kݞ���gmJ���t�>�f�4�/'�[���\�(�ӱ<x;<�ۤv\�llv��l=��W<�a;�=۶ݞ�^�1���5��}���6{W���\�vx���6�>$��<���x9(��N�d,�=�`�������7H{v�]���t@�>6K��ݺ�.nj��g�]�Ǝy2 �'g[�n}GJ�.����k���}�^�pM�yQ�:.:=���+�0Y�b596W��\��}�ɮe�v��9���IO)��p��8�C�\r��!��5Z#ـ�RaMP;�{k���cTb.�v^�.͗c��Dv�#�*���vy��7bܝz��Oa��M�h�ԥ�ò7h�hj%\�J��8�3���5�k�Ѵ����6��4�M���٭��<����qLG6)�Y�I,v�{�c��[>r�������.�u����qɭ�*l�H�tѱ=x]K���Ԛ۴S��m��m7@{��L�JhF�c|	�Ó8}e��t��.�G�1�^�p�d�vi����u��ჷgH9�CC�l����clۮx���b�3�s/�NN���ǫg{��콅��vT5O	�.��N��W]r�r��0=��ͮ:�z�:尵�n��%��pvc�Z��m���<U��^¾������9��v�k.1�tP�;x��3�Ŵ��[���cy�ph��ض�ғ��:."9��0���ؘn�{Zy�߿��J������w;�r >	��7 ==u4��鳝�g�\�I�D�������"��"I��.���lr�'�^^�t�9>@ %�vf ����d	���Z��sl��I�
�*L���f{ێ0"_e� 3�����{u��`}/�٘�*���d�)Vm!��*]%�ѥ�	e���U�|��x�� ���m ���w�m$�c��&RS��vL�:\� 0��LL�觳]�@���;���͸�&�s�=��� ��
}�� �����3�E�# z*��
Iu��^���:<��%�g�ڑ�9��a�uբ��������iB�Q I|����K 
}�m���+�'�h�U��ˉ���$Wm� >�On6�ϰET�SD��_?��I�^�3� c��;R����F�JbvZ���ާ{�&R���<����h���.<%��s~/|��g�����#k�&�/t��� ���q������@D��v���Sa ��n8�GU3�97z����"iL�)v�w��d@���� ����kո�n+79� 
w��@5���y�
3��:3RՁ��^�I���=�
�ĉ��B�(%ռ�a�yݘ�ؙ�[t9�@!Of��N(��&�QQt�w�j�����z��;�,R��k|���M�/;�0!;�m�J��O�B��HSP�A\]x8�wJ�+'�i1�l-���\M>6��3DZk���ʤW�L�{���7�" �����$�~�I������r��l㖶��|sݦ�g����P���	����DM�io�x���V�+)T��`�v�0_����QeO��P��Df�]z���Y���j��}W����@|]��cm����{RJ��x�l���l�<���]�gntZ���Z��i���}�`��v��;��'�tJq{͕0���nxt�_{�xfef��$^[[Ω"J�Ϻ�/�X,��
 �4���1�e
1���)�A�M�S��	����)��|�ܚő��'f�=�NI�J�*�}S�LԨ��f{�1` �)��i3]EMGW���v��4 K��� �"w��:SX廈8�r� ��$��xP���:�l����õv��u���c��Zz�j4�D�
"j"��A��M0 %���7�v�_plת!盘�˫���
_v�DbMjط�ʤW�3-�O��`����7f+��]��&���)��i�6:�ؙz�)�7�p����� �pk|���|
o���ܲj^�]���h��������L��=�UTTJ
��-�v���Ԫ�>��x�@(��;����?�����T��׹{˝���;����}�!�R�Y��+M�����1��OƲ�i_����Jۅ2�ܵC(Q�>��<��&OJ��,�81niI!��3��[L#o�SL�O�[���\F��v�` |)�s2�=}��0�4"i��������<����B���Z�N�m ��X^�.ݹ�n��sS�=���Ѿ�N?;��:Y�u�gv�}������ ����0�W�Sj�8����� �/y��$�D�
"j(!��m4ȁ�"(�E��{3y�� �^�@#��M� �闱8\7��K��{*�;�-j��*E}P)�lS�����|�nag��y�� !K�m&@�=}����"f� �
Q0�%�vQ8y���͛S5�H� +��� |�[=�F��IF_u�x��oL2ц�	�;��2�}�wĦ���%�I��̿	���K+�H��ɽ���� �^�6O�ݙ����Yɨ�:��{O��ӏ�o�͕N�qJ�������tY��듍��C*��6��m`~������__�w$hd^�$����;������{�w:%7	Â�Kl�4�u�Su�I���`uE��<Z��n%M$������s�8�uy�v=]�[�Y⓶sw@U�je�M�d�'�۴M���=��mX{`�$\s���K�[ۮ�`ؠr�"��{��xi\a�ղ����Kq��Kkf�W=[�n,��M��M0v�t���x۪IϷ=��u��t�i;ui�Z�o`�v�Oc�1"q�۔��z��^Mv�xn�^Gb�������P��LR��Yy��� _u6���wa&^M��^�XfvUR)#��W�4��H*&�E������,˃��͊�Y�����.�m�&�����I��m6�\�%6)��L2�!S's�� �	E�u]�@M�Q/�ɣ���s��F^��"@%;�����H��
Im
^�tzg�����f��w� �Φ� ���� 
^��ۘdu���_J:% nv�`}��r����*"%�[�����m2.=^�����p� 'w�� � R�������ϵǻ��ٌ(�iM���xz��:�y&�\��6�]�'���>g�0�$A.{�j��Ce�%�J|�Msi0��[�@$�/y�
,u��=g�K��� ���70��;�-@�(
��.�B��m��ⱊ2j��[2r�N�Pߍˈwc�����y��?}�a��K��M�ʲ>�ll/h��ڜք��ȯ�p������Ʀ�ȅ��ۮoԉ%z;s��$JB�m�|�VZ�D�md]uv|��#}H�TUJ3;�s0�K޶� n�/ݱ3�Y�9�nf  B��RkӠ0��-":Ks�󺌎YZ��U���|�{�����B/OH�5z�	=N�n�$���!�J�$�)�s0@ ��S������6����}���K���`$e�URP+6��ۚ�g��Ca�L�i��awb�G'V�kTb����n��w-�r�8���}ߟ��-  ,({���BI���  gw[�����x��8߻2# ���`�q��T�PERH�;}M0@��7n�j|�[��~}�@�Q/��F_O[� �mw}�'�M��rnL��$uB�	��Aԑ�O�����d�O����B	#7b��(�H���th�t·4��VB��f� �zJ��[�2XM���n�c�ݘԅN��5u�m�s�Խ{��r�K�A`��< ��{Y�DS��C����&�#}H�"�8.��������ܦ��HCܙ����?�A/��)�dM-�L������5��D�PB?��ӭ� K����}�魚��i�F�s���ӭ����>��ٙ�N��V���~�ω��B5�L��=;�jۡ�խ�r�cQ�)����$��h�B�`��"a0M�۸�A���""��٘�����_����c oU��9/Ù#х*W�m_]��#"�̋�-�';e��| z�v���ٙ� ���^��Tu�%�t��&��p�D*&\�J�D��y��=:�x^�^䄬-�ׁ|z�y�$���3 ��a�@Q5ARIJ]�,}�T�϶%�oKi� 	K���� >����s�����/����<J`=�V/,�Rm#�
"�"���	�e0?9���"O�M[�w4O:طW!�a�W����D?�8}��m@3p�F�Ջ�����ϰ ���l>�QQ骚���VW�� '=�o> �/y���A�Z�Zq�ȎPf�bBMf
�lS�E����u�;R۞�wV��]��������A�Q�s� >	�{�%�D�|��+��t�gEc{tz��TA%I�7�Z��R)*��g;��*��F�gjd{=Ӣ��7	8I�'�$$
^�i���WI���d�N?)݋a
f�@���� �R�m���B�W�*��S���@��ۙ� /y�x�w�T��T�LŰv綬p���i	��۱���ǟ` >%�;h >=}<�s�æ�bb"}���zc= (����)��Ǿm0%��Ғ��|(�y��0��I';�vN ����  ���#���.�Xl杊s^�ձd$�垸��jn��уr�{��a���ua=��[z�oMj���B��=��1�/l�����3?~�Ө��\���#<Z9d�f}��n��ql����Zڍ���}m�y��;t"������un�Mf�z\k�]��e۠'��rg�c95�m�1�li��Qguci�c��_�Y���ok�J�F�bǫ�����]��������q��ö��Gj�Z������gq�v��\������v��j�[v��;�����7�{;�A)�H2ux��O��mK�חfS�d�M�����95��[�LAQD�܉��BMÁ�]�W� @��]����4���5O��<+��̈������檨�&�"v�o�u�"�q����5�_�^���D/�� z�y� N�t�8�c���Zܓ�4�
IlS�����O4� H2r��F-�^��'�� R�[d#���C�=�8!L����;'���_con��B}�m&F��X� }>��Ʒ"o޵���V8����۪�����AN �pa&\�RI$�o��ָ��|b#ӓX����� �ݧ �_u݄�zfik���]�	n
-CVǵϣkq�.W3<��ny��`�eK���N��A���G�@Q5AS2R��6� :��� '��� �_�ŗ���dF!���!�u�����y
)B�*��.�3}ۙ�U�>���s�Q���qd˚W͟I6`���[=3s�Y���9��n_AF��q�*'�͇�n%ț������P=h�}�7�$kZ+�����{�ǟ)���RY=�M$Le��X�H�{���=��u�֪��&�v�}�M0@��n3�9�KD�^޾��J�5�$IQY�w~D��z4P9��3AēeX�b�eI��(*�Dwo�� ���f W��~�'���2�6J���$��UD@q� �m���X	 };dnyF����qW�q�׽�� E^�[��<��=�S�O�Ql�i��E��@���ca����τ�l����7m;D�}���}��0��.u�H�{�V�"W��`�f�غ�q�4�״��:�vf|�<��S3%"��|�h7*�|�2���;�O���]�w~I$^�tЄPH���$�Y�2w��4e4Z$AM��U{�v�ROj:kЉ^JBgO!�T�I�T\qu�%�y�s�'�������m�ǜ�����C��9oAդwٳ��}ކ�U��Q�J�����ǒ:0�@�sb��?��7��|������CV|��=f�������Apz=<��1���w��a�!l�N�͐qi���&��퓖��k?3:;s��}��zM�y���)��f������3�;�fN�I�ӎr�n2�[8�Ћ�{pqݼĿ�6���uAv+TՕ���y�8�!3;��W{�?f׳�љ;5ɏib�.�r�ʟ�č���:��55�k�]Or{�89�|�9������f2[���ʋ:nck6<o��ٟm���i	��w�/���g�)')e���#�69�޶kgY�6݃r��j�E���r��;G-���[��Ī2^8v��;�L���Nz�T�[n���D	�cӜz�I��v���̝�g�`��d�AW���L
r�u� @����Uw��8q�s�T=�k^�q��(e-�f��`n{�nAsY��5x�φBjΨ��	���ߗ<R^}�}�����V�"�^�B��x�_{&����"g˽�~���~�}�[��l���&	}�xLKyQ�y=K4�NiH2�(�����ٻ.iR,�v�pBh�U�I=��h�J�8�׻3��=�L�r���7�P�Jsٝ�A��'��R�����z��t�:7jvn��7�Q�t����'�>�uY�;��H]���{}���xY����=�<�����̥�C���]jp�ޚ�o���4��w�f�q,V#yk��Eq�1��ֶ��%r�b��Դ�Ԭ�c-T�EZ��JQ`�P(��*QTb��"�$DKEb9B�Z%�b�F֢�V�EUTEP�m�I[-+Z �J�J�Pm)eEKh�Q
4��h���څ,�ff�Q���Z���J�b"0�9�-�*���m*VR�Ҫ��
�,X�Ŗ�)U-��ҩR���Q��Z�VAZ[lJ(�,aZ�eKE�TƋl��k)mQJ�-��ԪD�mEjR�ZѶT��6��+UeJ�D+R��F�YZZ#
�"��֨ ���VŊ[X-E����T�emK��T��f��mb�,�VV�""5�iTV-,*��
����m+m��V�Q�T`�(�5)mc[�FcmU�b��k(�T��m*���Zʈ��UmKkiKj�l���Vҋh�DkDQV(����X�*X����2�TEZ�UKE�����X1R�S�"0�Z��*�AA+YR�Q��$�����Z�HSϾ�$�	�G�P�$�Pl�!0�������l�dC��3P'u�� >W:�D4�H��N��]7������`T�TT
f[H���� ~�2��sP�E�@}Y���^s�Ԑ }��=ԫ��f�k��ƹ+�k��=�^p�0��J�۶ခ ��"���o}��D¤* 	��eg{Dg�+\�� �_u�h^���{:&mJp߻7�""���l�;���Ӹ�l���l�m�x��_�n7���X�@|���^���[�ur�a'�8�(�5$w�nO����_u?� >�����w�ڽ�ݨZ笈񯺛FD<,/Bp����U��q<����rW�1���r =�p�D����޼�8�:B��(l�#)SC���Y�㙾ͯɖΛ~�p���
��<�b�٧��g	J���u�o�S&d����;�� x�$��Q�W� �
�R�������#��տ0@ u��0Ɖ�s|���ec c���z��uF11�c�Ĭ��(�&#�(zwN`÷�����Ӏ5�]\]��]c�#�˽�2
�*��LϹ�y��y��$%Ef��9�2*8`���e�FOD�啺꼕�:��PCD�Pf�+��&B��3{�}q�$�{�D4�of` u̬�j���٫H}��o�%Jj�$�u}Y��/}���d�U����4"#��V�".��&W�:�(�H��|��b�v}���^`|�w2�/{�1 �s̾�;Y�<�H�q�D���lD����Z%��tב>;�-3o(��s����}$�I$���G<~���Y��=�D��R|����e���au��ɴz���d*#�+�=�g�������w�հ�{�*6\�唓Ul����{��;ru�]��ۆ���N��ɤ��S��
���{�"�=��z�6	���//��=���7X͹#����E��� G0�9x�Iy��{Cq"%ƞٺ�On9��[;��;U��7V0󶛌�T���lrz��M	��� �OM�X6F6�MGT�e�3�1v������
�OGG5ǎ�w[�'ǆ�wm��;�ݘ�	Z�i���8�=�������H���oG<[A\��r����D�"�-�Y�j�ك8i�~�W��p�	y��D`V��?���2��@y並� ��ۙ��n8��)Rx�AW��r�	�'7���ٻ_}H�� ���٘��"��[RDD��N��W:{�,͚��PCD�Pj����q� �s�Ԁ��g��n�f�5  �����@"��2ޜþ"
J�U2h��zwt[���}�׋ ����X�}��d�3I�����Ϥ��UQ�BI����<�ʀ���j7̬����G�����$����>�m�����N�~��{��}��c�l��n��8�c�[O/�ֺ<�=���(��˷�z7��}���m�34U)u�5� DV��� ����F�nv*�$���}{wdߒ/�t�i=��P\���F��[����Ou��CyFmt훘{���Q���gz.ip��׺?�����ʽsN�Ie�.�����r�fH�	n�=Ӫj��n�!q&��0�o�wO=�}���M����t��_� �?�V�@��<��ρ�[�0�T��I�K=ͪ c�U���E���ױ׽	����v��Exz� �>���(�L*""�����Wv�! w�Nz@$�����)~��U6z���������4�7� ��S [ojဂ^��K����8�Χ8��}7�Z�;����'}�i���:j.�v �ͻ��Kx�6��rps��7e]���96n xn�?B�S���1�	���1^UP >}��`�)�ofbA�;b�(�3T@�1�S�؋VH���%�b%����K�3�S��y����=�p�O�{3 G_^N�o2+һw�Hz�ʦQ(�i�I��}ݴ���;^` �N5y��N�͕b�E@9!��=������o��i�����v%.X�1�6��t�v����w��o���N+r�4�������/��s��� s���!�>�����[V AL0Ȅ!D�+:sL���nݢh%�m�&�H�ͻ��H�W��\�]��K��W�J/��$���P����%��^��>�@q�n���ǵ�*��^u��;�ّ�Ei����T�B�f��;H��4#��7
OT"����vM�o?������6�5���}>��w�)RTL����']�����D���Q^HU尯7P�wSh ���� ��;�±6�I��w���Ϥ�DE�μ�x�ԒH$���n�&�՝T�$ގ��l@����}�%hХ
�ۆ����=�{s�����[��Mǫ���P��{� �����>+Osj���*{�"�Ť�������s��V�I�H����\�[���M�� �}���WvUl�3��Beu����a�B竒�q5r�gǘ4ý�b�����n��7�4n�c�2�=���ƖV����������FBK��n�ߒ�é�S*U
E$���~�0� 1����%k��\^L��z����fb��;f�D����RP�B���������u��ֻ5PN��Qm�1�����-��ط76��F�I8&m��݂|��,$��*{}v��N��� >금���(�����un�ݤJ
9n�5��a�p|�n!"�.�� �//OM�FE�6�� >��1y�U� ���l�9��ΐe���������+L$��l��^� A�ٵ`O_�����}}��1��숁����i�LUEM*t�{�r�޿�z���m+�B^�Κ5�B�_]��9�3�$M	�R�ӓSR����S."�4�����s �{9��3U��O>@x��O���8�`|��;3�	W�7�C�s�[�CdM� ]r��uF�s�Q�f����}��{ϥ�C� A3�o�w[x9m�⯎�MC�٫�Θ,���������;�ٷ���^�d�r.,���)0���<����a�=�����*vw7Rꖶ��Uk��Փf������8Ӻ��H;v�5Zwd}����]����wl/2Bu)����ۮ^:ؠ��$n޶�t &ݰ��b�	�7q�k��k����>n�y�Ky�F�[sqok8�M��m�lU���gϖ�n��m�8۳�8�zk:H�k��x��f���k�s�(%�''m��oYcSrs~w�~����.�܊I�"�/����m6)�����dE6Y���K��J(��s�{���|)TA��m߻3F�+:�f��q}vՇ� �w��HS��M=���+�r�O���=Q�"�>�ML�6���i �}ٯ� 	#�:��*�須>/;�� >���HIPZ�@��Z��VT�UL ��� �s"1|1��!�Mc�%�$�gs�	.F¨6m8F4�+�ݺ$�JvM	G+R�T�[�ϳ-�_A;�ّ�'N�t��8��^=�8���A�,G�	��tc��[uYx��q���iwV���]���~?m,Jh�w�������n"1���xLk��Mɷ���>ߓdJ�|�I1�f�zd��(��v�4K�p�h�Q�W��X8v����=%5,��/��oA�u���y����=�O��Q,���G5��+=��:��fI�W����	���3"'O޶������;9����F�f`�!��	(3�EVu���}n��-n����t�x ��f`N���ý�RD�ԉ��h)��GEl��D�7���;�@ �N��@ �Ξy��3�j�٤R@+������zH&J�U30;fq��� �ͯK��{�P�='�� >7ͪ �^t�jL�U^�q7��7����G��j�k�铪���i�EŻ�.��+�ӝ4��p�/_7���}�Q&k~_|~��s	�޹�Ξ��K�ر��e%��7a �����!��i)6�U4�����-ǫwx+˿s��A<w�Z ^t�rA�)�P�_u�����u�4#Л&� ����@��O4�ƞa^[��
��W�Җ�#d�{��f�8ch]B��o/�S��K7�Nw��:��(<d��N\S9�lOk�{�u��������3��1��h����:���ԤMŴ�~��3����U�S  ��tD +�V���Jq�f:�X�`#8��A���ʩ"g�D�̃7;cA>}��竳Ϫu��%�nX �o� @}8��1��Z���Ħ��7�T!�)�ڀ���[��p"GF�;�<���NL�]#v6�3������S53J�b�|o�t����r�N>���US;�|<�gktDD^y{�'<a�4hѡb�Y���2��
����Ν�j����ZȈ�/��:���}�B��iz6E2ʂ 1�jI���[䉍��M�*z�Q:L��pI8��UzA%��&č4�w7�q���s�y�r�d^$��s�0|�����;�w]ڌv��$�"}s�lMh��^8��UƟ5�C:W�l��r�J��g�	�`f��od7��$�Oȋ�i���T�Np~�͓�.,[�������!�o�ԤM@��a��~��� 	�}0ro7q�N�юw�n_�ݼ�M|�{���@�y�];���N����xߛ��j:�Y�t���m�&�Ӫ��۷ ��mL�t&���}����&_\2���&��DA:�[� �g����i[�����|��"a'~�Lߐ���[�P��g���7)�<X�q�:Ӑ��q�f`�Ӽ��}Mk�s����ѣF��t=fz�� �s �ޙ�*7��6y��7�	��n# 'N�t
vc��*	�*��"����;w��_=���w������i� �/�������o���.���)T��)%�gm���秛�sr�29R��fb@ ��mQ E����?}�E*��A��cɾջ�-X��.MD��HkI������JG��n�$�P�α��� P�a�#n��kvR{F���]ιV5��<6�C[(?wf�Ӌ��{�G*�;&�#��)�%��7����^�z��?���(ԛ��]"�ꐖ�������e��A�����Gv%�DN6���a���=\ʜڋs���rK�m�s����|��<��C���"]���x�o�Ou����q0�_d�#�=�ٛ�,��<����ojOߢ��?yw" y\'b�k�q��%���ז$�:���I��pFIs�a����]|V޳���|� �e�w�Bi� �Լ�d3=�>�<߶ᝃ�6uRV���#�k���gGQ�KY6�K��ܐ痔�������=õ�`.���ƍE�8i�����E����Dو|�|���,.���,q�����B��$�#��Xl\����r�1�) �
~�|�������˱��ʸ�>� ��6";����b�0�*���lK���3b�UO[}�}��k{5D���ފz{���c�,�����9�g}|�z��_z��aQ5y��ͫs����.�r~Bq�;��=t��5=�qv����ik�/W�x��<���h/������g�;m��ܘ��Lx�pW_���zLK}�4��=�����Z2�����}�k�(y���\|�׳Q"j�М�探���y&;�c�c���,�Й���2}�3(����M�U[`�1�Db,�(�DF�ѤmTm�J�QT-�b����֬VյZ�F�TT���r�-%b��-J��*5)V����$m�V"�jX���Im��U����Z��4j-��J�E+F�jR��Z��,H)U-���S-�F���jV�DX�����,Z5Z*�KX-A��b�EbV��Z�ciX��*���(�eJ��Z��Ĺ��V�EJ����TVЪ*�[F���b�j1Z1E�iKR�Z�EJ�Fڠ�iR��Т��6�EZյKYZʢ�j�-��f���J�"[b���V�YZ�FZUm�j��5�Qk**�1UZ�b�1m�5h�"��X�`�T�jQUb�5���J�eQX*��#B��QcahX0PV�X��+,B���h�b��`���E�DU�)Z� �F��YD�h�Q
4E���jPYJ�1�QJԋEU��Bł1--j�����r�5e�����n��4;�Mx�2����|w�gy�fW]��s�ݐ�s�sWv��;[ֶ{X����^-��nfn�ug7��mŷ����Y�.1i�WH�c�s0r�vÍ�@�d3Ӥ�ݍ����ٶ���U�O�Y����c�s��.^�0=�<f�]{a��p��Fp�W\�j4��]�v�83��vݛ3[=Ag�b����zChuۢT�E�ܦ�ZV��t�&�*Z�۶v�[���\nʵ���=�ոͱp����1��cp���������Ý�W&�ϗ�_	�1���\/B�mmX����秉���ݻXr{]�y1���Ֆ{vz����m�<�[��S9itgu�]�L�.Sn��]��Tg���q\=vr���w�vM���k�2�Ք�C�����<)G�gG
 b�e9ܕ�9����f�<s�Fq��_#4*�ojM�K�wl,ΰn}���%�]�[����eg�g*��/\�����{;1ѮӢ�c��.�]�|;���v�/|�ݶ3t'm�q�auv�a�ƣX�;[õc�iн�ݚ��$}�s�#�фhk��sغ6����]�l�����Wc)�v���Fmu��g��㫯=mϋX��Lĕ1���l�L�4=��8�K趇9v��\n�u#2'k��<t�'wҚ�ݹ���L�v��c�ڗ)������sdg]�=�\��m�"��b���RY�}[u�ϫp�8���������k���XS6p��W�[r��Q�����n[c��BN�lq��.���A��M���O���e�zH��[k�|���I�mI\u��k��r��78�S�.���y㧅������5�{Y呸�ca������Q�϶�=vzݮ��ps�s
��a�����ޣi�.�γ��e�8��a�\vs�p�q��V���m��ⱎ�!/M�d��<�<�l�����X1�oF7�]�\��b-*zm#���j�X�5V����>V��͓�oj���]�{$r�����7=OmO]���aQ^}�W��q<<�=�O��w�^�麡�n�;1n�-n-�^�[�:�f��X�ɺ��q͔��f]�<�|��W�n�	$ck�n�kk�$�_N��Bq�s�3��'(E\n��Ju�����@��\�ʬ��q�.ܩ���wۜv�d������\��y�"&�؀��Rv��Jan)�n���L\�!2Ew?��?5��b���^gf`$ N��* _���R����L-��e�	���|}Z�"Y���n�"z����@zTt�[� ;���w�$�I[=�, �O7$D϶+ǫ�c-Y�y�'��B1�bL�W�2�4J�/zy� 	^G)�;�~� ����~���>���Q1Q*j��3=ە�bv;+6���� +ݮdC@+���i��ѝ�.��$_��tz�L���aJ�*����f��r �}�0��A���=�/�>@��mJ($���;�j�/]�F

غ��n.��n5�<�v�+nv.G���΂��m*�&b����?IJ�>�I>�Y��@�[�����3\׫ӉQ�����'v�N���|~��r�[����AD0�=Y��0�
Y�^��Uy��&&����!1�yԢ���aX�$5[�{�svӡ�3�lmu��K�MU9ޱk���>2�I3��LM�|��_��������U�nr�)�@+���4@]g��Ā�dwL��kɿx"G/w�XVa2�6��^�T~$���kŀ�H:��x^��___�F��Z�)OdmP�(	w�vM��j���n-CP/��U_��9��Ψ>Zf�9> &����=Ӎ�9|�0�N�o>0��)�б-Ǣ;�z��{g-Ȑ�uZ�"ꀺ�v0o;���	�mHNN)�a��:����c,:wdI@��m��!�����{rJ�-�י��B 4NO%�ѭ9 	��<K ��{��UC��a\���[8ܐ ��f`	�[lG�0���WTl���+��_Q�5酏�v
�I^����D�(�	��m\�d�%�����o�!�jK�L6O�;1` �� uB�N�{ӄ�c�����׻[��X�,�6w��Dt���m8}�ܸQ~��b��}4�OH����S���v��x�Y&�c]�;�~��O>��I$�O}�d�aG�U�K#�ЇTXmBJ�M��MofW����� �ǘ |�*�I�2p�WU���d���o�ĝ���@�fO�d2I/z:�D�}�x�r�	1�����D��m� �nH{W��9͙�Ț����=[AQ��N<,m��E����l幹D�K=�q)��m��Dhf0"��u�mش�����j@�����`�ģ7.�ׇ���OO��~$ ��9��5)��,bD̓{ћ�P����g*���'.��`|��2!�W�y�" ����]�L�&�o� k˭�B��)�"�\�o�	Eg��� �Gt�FÂ��+wP"w�-� ��^��Ԟ��3R�i� �9�*��E�����S$���Ґ@[��0��������:~��-wW�;���.xhK!��R��{��7�^!����>Kw�:���d�"s�=�\�
z�<���)��8(c��iE�:����*����%��.q�R�$�Ss�' &��[�Ȩ�{����=ܐ^d���"�����7}�V�:\ʭ�#�6��a�|By��tعל�m�P6���&��ḁ���8.z~�o��b�p[-���/#)	$�tu
�PA7�٘�^��*���Y��y�)�D?�+:z܂�4N*���S4�33ݹ� ��Y��s�>�R |��ZƀA7����$���2�k/���=��؋f"!��dԓ}њ*Iy(�ޫ��%�^�x��������K��F�$ M�vf ն�!IJ�I-�_E�P���Zk���oU^4)D�u�$�
;���E DK7䒪��h�]��1-If��	A��X���Ӗғ=�c�����V��� ����� �$՝Q��^��g���`gR�{�a_8�q��q1�[U����lq]��?�m��Ѿ�i~СDEc�u�ɽ�4�<��`����n8��r��K�٫C���m0�s�8�1�7s���S���[u��e�8�v��u���p�\n�\DD�gn]��]v.�g���N���;;n����ʩ�ضz܏<���q,�v�W�3��h��F➶eڹ�:�� g�v�/���q�../n��5Dw8�:{n^^\Wjz񞱳�9:�+۶��r�4���{�&�*�N�1�mac��\v�R`�F౦���]����<`p������A��ڂ�~J*��P	${��g�|��XƐj݌��<}>u^x�8I�޾�w�D$�-Ѻ*�v�3:|ڐ�v��E���OY����vf| �N7$Ds��Ȝ�@����7x���r��T�'O�3ݸ�=��ԇ�|��S��dZw5�g����w3 @|��d=���TH��D�jh%{ѭCV:\\��d�m]� �O���^��w>�Ȃ�6�4�~��˻�T0k�$Ba�"�AG�y�@e_<hT����I�{��Da;���`"����%�q;���Wv����9�5d��آ�ٸ��L@3���Ef��Up�(��&K+w��p���)A�Q�]����l�@W���')�o}���ge��3�D��[�^��J�%J��*��l%���#�ɹ��s��]DQn�g�υ�듙�(�I��3u���L�jeNWE�����Ș#��Ǎ��k=G�)���Y�ێ�s~�n?@��W�� E{��r@�y��ޥx�`�D"�ѻ�I��Ȼ*�%$�����������{�v���F O��j��
�O7����-�Ap!1.��v���꽷iJ�s��{�a�A]�̈h8��%��o'-��I�s�y5y)�!-��>�������"'^��"e����i ���r��g�RDD��oy�UV=�������A�+�sV�
ݝ�t���v�s�O��mO�۷���no��߿~�r]s�1�>��d���q�%G���F�(dMVD+�fGv��� ��N�!�W9�fj��)���3 ����P�c�����تw�X �g�����u�$��ܱ#�j\	ү������CP�1DU �Ks�� O�k� g��U��޼Ư�dNoB�5����^��
`�;���yY�����"WW���P3.����Ȗ��X۸ն4!�
��n��{����v�('�U��]w]�a�Z�&�m3S^
��Қ�����W�= ���� �'�y�I#G�^�P8�p���x�  -��؉�^4~@�Gq��-�I��$z۳2̘��M�:��W1�>���wi$�=�,���Ӻ{F��l�D��M��m���'�ܶ8[sX]]��d�q��6��;c(꾍fF!��d��	gtl��F'_sq� ޺����{��v3ϣ*�"�Hz6��ɹ6n	�&0d��1٭��ٗ��]��+��,��_��� ���[��K�]M��^s={��s���AJ`&D�vfaG��Շ��:�[�*Oc����@����b 
��7���W�T�(SEQ0��=�}��u�����C�v�X  ��t�@"���9�]��0vo�0|�x���zD�%f�<9���3K6/b���:���]���h�����37"ʖf4�t��LR�6h����d�EU�a!+qn�%���*� �/z:�D��F�sef���&d�]�~I&{r�J)"󣦽
&6K�G����Rq��q7\c=F�a��ٟVy�u�lݙj7��n^����x~��,�~_x���ٟ`|�Q��`�v�1�˚��y	�U�my�� ���[��j}38�bH�MM%}Ѳ�v��8�΢k�������:�`�<�R@k+�|r�[�����$�hٱ��^�UyDvkvD^���DI�D�u���|Q�ʡ(��펤hf>��m6�R�L������sk2{����E�[�ȁ	>Ǵ�"W��z�$Cs���v=VM�.;�U){����������ʰ�
��̆i�Ey}�.�?��޲@�=m) @N^�f����ϯ9N���u��}�[,�N�Gs~����E_���>Y�yNS˗y��g�3�f͛�'��{}|VX����=��t[�v�:�?!���R� ��fa!��ȗ�&wacS�O=yx�c�{gm����|��s�1�8�Uۜ���sr/�V�Z�Ջh�m,sj�m�]d��:�^,�ldM��9]�91�m�;.�uW(\�y]�ӷk&����NuS�nu��Y�^B��Ok�R=(��cWt���N��EѮ|y�[�n��z�8����n1�K�V�&�Wk=x��[�\�����n2�۶W���u��v�����߿W�$74@�������<�s|���|�/5��[
̪��I}��^���aE��)�S7�]Z- �F��xv��R�bo"�_X  U�c '/z���I���۝�
����c����Qh�"f�"*!�FoO�Ȑ��<�����+���'v��b W�y���\�]�bF���m��aEPPz��MΗ�n��� ��r�� };}��BN}Xr%���u_�~uVC��s�3TU}$L6�/;3�|�[V{��{7sc
vM?����D4ӷ�vM��g�)����]9�ʑc�T���g`���Ӆ9�:��ٷM+�U�V�;.�趦n��8���� ���mG;�D�u
� N߹�� (���T���������mI N_kx���L�SH�(/���8�}\�|;���"ծ\wM��[�#�V�����ǃ���G
����Z�W��i���u)Ց[�Xvo�Y�js�:s˫;̨���D~%u���*;�o� A�Uc��dM��-ɀ�NT%D�4g���0���>@�U�<Uѕ�ޜ 9~�$^	�쪔��
�PQ�e"Y�mq۾z�8����������Q���@ \o6���7۱`|�{3�-�S��*>�D��1ٮ��Ex�7ZW�[�։@}����_ �����v@�+��tV9��
���[5�O��=�t�9.�[�fwi#A��fq�oC��A&�JG���I��/�qd�/��0����j� t�9a��399~�ouff��6I����ś�>�KhB5^J%WW���i�N�9n�k�"��iD_��:��yܰ�3�;�M���a6�U&�f_�� A|w7@5|�t�Ωսɔ_<k7��- ���YMꗁ��Z��6���ǖ�}<>Y�գ<�w˧q��{ݣȞFk��;��o��B��y+5ȵ�?\����{���@xs�{�<�v� ^ޫ��_I^�w���i�ry��˺N�K��/�b�9� D��[$�zVȇ���*��f��]�W�mTc�����}%L�t��/�d�AmՅ,�9�d!r��ۆ3ߤ׫��&?a7�ٵ��슒�{�v��۲��zr�gvhH,�Z-�2��;5�b��;L�R[���#�'w\Jy��fj{��(���3�z�2�*�c�g����I�
�s�;GA�^���F܇��羪?������=^���p-�ξ�&�"����0�'��$pOp5��Z'<B�S�o�ȴU�{ں�%<��yz��%K}F�~k��f�^���5\�n�r{@��ܨo�3�z�*��6^�ֽ�_M�����E�͎����M"✇'3����������W��f�7>�Ɣhxy��Ze�o���l��������[
㽒��ӅV�[�{���t�6��E������Y}�*X��s�ؙ�:�pH��T7�)�cfu�Q�=�����}���*��=�?+T�n179�_g��8lnA��yoٷ���v��{<`�u�.����a2���)/�cV��ƣ9�4+w�Gc'0O�$/t�����s�nI��a�d��_��F[��s��s�߉�ea���Z�����J�*���%��b*e�T���5
ƵJ�TH��"ڲV�V���Db�m�ؒ�BƸ�r�B�+KE-�5�m�[aX��*�ZXZR�H--Ue��1b[DAD����kE+R�DeZX� �+Q��ȵ��+b(�lP��@�X�h�X�m(�*��`�QI[J���T�%j1��"���V1��R��UZ�R�"�`Җ�ڥ�-��+P���m[iI`�,U�mk,AEQe�U �ej�����%l*Q*�ZPX�2�kb-kee-��YQ[K@JU-�K����
�k���V��5�m�JP��ʖV��cJ�ʖ��D�T�m�Z��J��DIj�R�U�DQUX+m��"6O=|�@"���� ��y�A���\7&�:
�/���N�#�g>��S�iX ��}�Z 	��̣>t����,$A����j�/A@�*����mi�� ���7�],�W���L�/st@�����灞c\�lh�
	6bQ	���1�;qF�Vۜ:�뇪�ŝU������������3J��$���a�~=�:"�z��Ss���nǗ[L��IO.�A�[�5���wI�Ȅ)Ϥba/��]9����� >���, ����D�v�p"�Oe�zR�j�2�*Hl&-�I؀	���|��sS���� ��mY����H��x�"TT�*������y�rOd^�,�6�Hpm��݈"'o��~$�'��]�#W��AJpBP�G^T���J�N����3�F�Z��;���z�J��ʆ6�	�.���Z;����+4�^i�e�$��=t��)X�n<L8)�t�_]�D����n��6~��x�g:h����f$ I�u�43�$͜��.�n0�F��a�b5�rvr�
&�{\����2Ӷ0��΅��(��,��p�d�{�C�� [=�_����.'��\?jC9=L�	/C�ۻIz����l�DaKh�v��C*zc��ӕ���N� S^��ĀH��mQ <�j殻�&I��O��~)n��o�B�'�L�J�rڠAMI�ۊ�푽��@)�w]�K�"�u�4��,0�"D2�"�	�|�9B7٪+u ���� >��t�%䌞ޚ7�F�Լx��I��>�����P�QSH�*Go��O�P�D����M�\�X�O.���M�]ߒ$�蹡�����^�w�w�����.|��i�A�{��V���3O0�_��oَ!]�'��v����i�)�l�C��a�
�Sb�Q7�ɝ�Ҍ��Ѯ>���ro=�ݰKvg��7Z��e�����0f�6��+���y�p���6ݐ;;�5��]v�v�'%�c��3�m���*��v ڷn�o�[ԡ�pu�9��d�d#���M��üC�g���/�7;c�	�j1�v����lձ#g�v�]�v:4����rC��U]���lFs؊4�����!u˳��瘌i�A��m��ȍŎ�P��۶^w�-��xnMc��n�߿���i��L�w�ggf`  @}goS&7`vҨg�872�뼻��I�d?j��� ��`��<��^���&F��k#�*�$�o<�A$2{zh	D�g2�2��-{wR���S��(��I6�/�[�A ������ ��I�J��8;)Q|﻾���ɨD��ު�#�4_�3^R��x��S7�~k*:� ���rV{y�@ >���Üf_WuNչ���t^d9v��@ţu~D7��9��?� �_kqx&tϞ��@}���4 ���Ր ��fbAN�|�W����n��Gp@�9-�;Hs������+`�.8k;.a�D@I�.;�90��S`����3������n�)���ρ{Z�"��f΅oO2!�q������M�AN
b�y��F�yHjkg�*ۏWvˉnr
�͈b��q�T�iv��Fj�8c�kN�@U꥘)Ǳ�z7���M���85�����G]��am�u7fEƽș������$�Qs�� 	�\I\x��l�T�\�2��TDED;F��� A;}�>����8��]~p^�]�"�|\{��d ��z�4=�$&�P��
(��ٱl.|����Z 6+|��;}�� ��eI����a̜I(5]L��ꀉZ�Ӥ`X�e9��! �;~W�"�~�^3�x}������t�;}�� ����!X�^3�����r�b"�Ӻ鹞ݮ���v��l.g4Wl��ͩ����.�qMB$C-ǡ�%k�¥{�;~׋��*�1�H+gٯu��V�'�@FNu��!��A@)�[L��3:|ڐqQW1���v �S��fbWt��R@G���p�s1F�o����j��
��N�=�^� �>� ����g�(��ͪD_�{��^͢:6����t=��H�R1���}�5�(���. �ɾ1rC�o��~zEy������}_�9~�� ��6�6�ӓD�SD�M��m�#)㮉�(^��$b��<K "]��0�7�U)�c���D�-$2n����JQKh����> +Ǻ��7�)�j��5��f �]�����+�zܛ~�[�������=���B���:�=�\DD�*κۮkrcsR':��k8ظ٠����׌3�Ds�m�݁h��l\�%�O���:"";�5�
}w������9U�Hgd�)�D�e��#D�1��U}���{��}sݯ� >��� �<ܐ ����^E��'�6�#"}��B ��-�1S^W�T!�J{�hT���{Dc��PrX�˭�I/'�8Ȇ�/�y����x�������u^Wy}}��hJ*F�)W�,�r&:kА@ �z���&�{3b6����En�I�\S��u�2'�5�ڣ}�^�C�k�X1T�-�����^��?_uU�}1��}�,;�JXoP���&�.�3�B�5ڼ[5� ��v�k�;.h�@ID(���7�Zr k{��_S��nV�[�w���/�y�" �k7�-,ñڶ&�в- [P @��0Ù�z!Փ<�.��2���f��;u��J�s}�����]�5A0��&����C���[�SY���7��t��m�D�{�גA��͢r��� �Ii�0,A�*O����[�:�W1eud��R	 ��Ӷ?�k7�1 ����ʔ���ʣ�~r������������M��� V�� .j�>�E��7	?�8z��oЊJ�U`�e��%6Kp�TҾ�ʧS1�%�Jr�%���*K�C�ګ�D�����<���V	΍����U�LUC�ǯ^�
�)��bKб�r��K��̼$�����N��6��n�{�Qp�W�>�ʫ��Z]f�tm��e�z�9�$ķ`�`��������yz�ic6�zuTd��V���S���F#�7�1�J�۶�q��������9�=X���M�nt�	�A�kѽ�gȖ��\yR�V��ֹ��Ig����;l�==AA�x�^9�Cofힶf)N26�N���B�"n�4��=�kz��1�\���\�q���\����n���8�]6(6��E�6��=pq�bޞ����,u��s��u�Ka0n��n�ƹ�X'&Qoc�r�[lv�wakaػ���]����'�+��ewN�Dz����ښ&P4B�!���[��	��y�� ���4��r�-�T�3���<DJ�~�	�{y!�����Sd��nA�]�&�۞Ϝ�"	�����>+zq�$/�w�W��|�7�氂�-�H�X�eI��!$��yN!� �u�������8 �{�1I'}򌇙g�(�J -Z���xJ�=s۱�rȂ�=��<�@ ����i#=����v0��!$2���D/Ta��ա>fz��b$����:Ә�����\]ǀ[ۻ�� 
��2!��mI�T���_D��H�URn�W���u�'0��'��f��Ⳛ��x[���V�ߋM�>m��ݥ�	<�F��(Ok�D��~�9�]�\�@Wt�jM�Φ������h3�vU�x'�����"�Kcw^��q��I_���=��^������G-+f���Öo�=Mb�����g|�_�45Ki�`/gyxG�6{;�l��,�Xn�f�3[� V�c"E��[��eUס7~޷�5ʸ�USH�DĒ�ľ�mHE���9 ܹ�մ�������+zr��@}�̏y~��Si�����V���R�yb���"�ݓ�C ~��0k7�<��L��l$�6|���'�Q�� Z�,�\�ͣ��ĭ��!���ފ��o�n�64� H���D?��k7�1�]�gw��VP�#�!�$[P_���=
�N���6��N۲��0�v�<�D:M|���O���V����]���r�:Ә�&�y�`x-δ�&����V�A#8�&��~�	��i�6��;�G��)y7.�������)��̈�nm	�ϛ�5����5W�I@����L;a�v��""k{�, F��jC��0�q<Ӛ�*l���(�5cM��f�O�Ί`]>8��v�Ƥ6�蹘�����ċe���=N�5�wђ���j�Ͷp �y�� ��ofb�qzLTT�*1$�K�ֽ���r��>�i �k���Da[ӎ�/V�U��Oa���%��H����M��Db-���ۺ4��A]���W�s�O ���׻s!'	8w�(�>B��B ���V����tG8ըn׳kEӰtV9�GL2��)	�Oo��(��p�0���5������!8H}��^7d���X�Fl��Ԣ�K��z��F;!XF ن��z�Ϫ��I�ƅ��}j��������{s3� EoN6����"/Z����:m��R���Xm�ӈp�:37;3���t忤9%#�)C��M �SYۙ�oN2����H3D(���+�v���� )�s�"��uc	 \v��D8����m�ا�/A���<��z���	�������'e}�G����N��&�˫\�e�y��&'5`�{/M�9�Y��/\����$(u��!A��}:ڐH�4���[��"+��z�H��nH ��݋���������]���8n��ގ����)����cm����`��r+������v�W��_|Ngf8� V�� ��t�]�Mw5Wx��=�� �ޜnOgTO��0��aM%k�� �	׽]&��[n4 {k�@$\v�j�Rsw-���5��H�̅~Qe5:�o�.Q<�ڢA9�3��b#P����A�ȩ_v��#U�0�Ch��p�HY]S}�B�]��zI1 "I!�gU|
�ޖf�u^q$�$�8�G�#��h�H�4Ah���(���B6NX����ό����$T^�Q�^v헷s�囯t6�yQ5VF=�T����ӄ��
�j���vo��5��˾�����7��׻ ��O�E��O+��|�����#�U������z��D�e��=�j�EK����/l� |ǁ�w}��喎b���q({Y���|8��W{�yd�X����W�Ȩ��Ύ�z��:�����F�N+��e�=��I��ġo��v{/��x1��{�=���􁛮b�{)�s�Q^<=]����R���L'bz�!yшi�N�Wگ�ϴN�˝���T�.N	�̈8�S$��a}�z)��O��O!B�n��f�Ą�&of��wxH���w��&�-T:�#U��1�o�"�ן{�%�c��=�����t�x�����sd��h~7;Y~���в�/�>i���a��r��=�ݓ�) ��u�t��.��wK��r��x��PyxE�l@kHS���M���_j��&�G��wn_aTo��۰[㻢��n��	nw�X(����q<�:m����.yX��ּ��F�i��������,%���|D�և|���:���{ҕ6{ŬYHe��k�xOt��1嚼9��_=���!�r�W���a�QZ"�i�4_j]�L��w{�������ga�	�ۿ{kp#z�{땺��ج�^a4l[ �~�5���k��V��E0�C�����i|���̊���:��]���m�Q��^�X}%�e]�3��0�am�
p�����4/�-�PQjX5,�km����7i+�
V�V�F5kkib-�Fе��"UD�[B��-m�R�J�*�"��cm-,A����Q����[J�Q��؉�!r�G�r�����EY��Z�
k0�B��b��MֳEWe��X֍j��Z�(�j�Q�)�fq

�fd�ֲ��ܗTl�e�PX�k�mL-�q*8ႣR�aW*�G1ʊi���(�K�2��nfeB��8�.X�
[�90�b��b�Q������VQ�fc(��e��SJ�+�`e,F*8!��wn�;�}�Snɷ��9����Z�k4�������D)B��LIR`���"��F�EE�����Qm*9s%�U���3*�*Q-�X�
�� ۋ�*bVڪ�-k��q�+�V���J��ln5���4fa�2���G5��t�v7�ʺ�6��zÐ���&M�NW�x���w��mv�{ ��"	�W)�w�q���د/7M�p��{vN"����l\s\^�nܹ�%���h�;0�2��L�۷ko-ն�v��t5mx��F4a7\݈[��=olk��ݷI�&�n7#���TG��nÌ�A����r搉ۊM��<WV��;�����s�ݞ�x�F�����	�tRu��۶�vx����Md��7 �@��&}�c��l��37uuQ�C�{u��E��燩V(�vq���[��szx��s��O[;;�����q�u=��s�h� ���l�m{3���m��cv�\\�r��N��e�P�.P��6ݵ�Nst�e�m��w�nL݂�z9E����;����<�nӎux+��l��m���.���E�^�(��6�y[ú㣲V$�u�hx��pGv�Ԛ��g��v��hM.�ѳ�/I���v�q��i�ld����'Gm�|/nE��7Z�����K�azۓ���<��Op�'a������\O=�n��h�T�����u���1[����69M��tw��Tq�n�W%l[��I¦��Wr��v7m��m����`�']��	��]����h����8e�l��4�d1X�xG��t��4�2�y�aM�7�-��=�Y�LsN#���Nݏs� x�<��(Օ�˞2�\z6`A�yBu[Or\��ס\����q�ɣ�g�c��9�F9;����N�|�6���ŮvѸ�LZB6wP�Lफ़N�q���;��q����^\�nDn�F�8{R����m���A�۞�:kn��8�z�+�����gzq���㞋s�n���=�����L���v��2�N���jM��a{g�DǬ[�$\����E�i�XҺ�]��7i��\�#/���;�+�%���Q�*�&�_Y��ns=
U�U3�q�۷*3+@E��7;I;q��y<���=7q{��/�P�wn���M���>˷�lu�ϛ]���4ᗝ�r�����R�pk��ڇv�>t�:\:�+b���1�Q�)��v6�H�l�ye���nݏ�g����W�t�u�ˮ�l%�5s�<��n*�O�d�9z]���nq$���(��mq�W�|n��n�ƹ�tk�vc�ӝ��3ю��綕����s����:MMW;h�3�|��~~~�a��a@/#9_fl���ު�]-�{�{"��x��v�3/�T6�p����}��'S4,���ܺ��ڠA�ޯeM3Le�"����f-F\���f�q�o��ⱹ����Qbn� �
���m�k��c=�b��7���4��E�c�P��,�뉣 �yY@Q'�F��Az(&��j���&몁6��BD��C��U�uD�J����lwF�SաeeOH
7��I[�RDU��vl#bD/h<vu�:�������g����\8ͽ ܊]�)(b >��m�	#����n�J�ޚ'ĀJ�tduY�l\we�x�T_t׉�����l��2�=���4����b4���sWl�س�R����8�V�X������ܛè�zE���y�[�E6y����ys�5b�ec�*�uߋ˾�|T^t�>!oEH@��tKd�b��'2�R�D&���l������ʲ#{k�tTMd�$(�ڢI+z(��B���iҀ��w��������$��� ����4\��H�1�B�D@�l�P�Ux�dY�wmz�.�{����s�5�O�]�R����$�p�������[$�M��1�`w ��
](Y���Z�P�Վ݌�f����{}O�b-C��:���A%^�J�}����3k��^��U�튟#��M���b �j�7}�T��7/ED��N�I�*�ѐA��ު ��QRw'ۃh��3:	4C�F�!A�T�a�O�}��D�v�%��I�e���g֕��G�/s���\'���O�.�>�����a�ѱ�Naqɖ6�U�¢�-���dM3���I ��$���Ne��6�C���+�ꎥ�:�&1sd��f�*/��n�s�f��|;&��~#�ڌ	p-:P0��ʭ�Q��v� Nn��"�TP��I�!�f���M��2��
.���oSIsIU�j�9i�J�F�S�m�v���pc��X�s��x'b����O�W��/��"�ȓ��j��}�@�3q/��ۂ�c/�C���VU@�S-=K��F����n-���`�˾�3 ���}�T	�ﺅވ8j�[Wh�wSmI��,��w��@���MA �T)�3��+���]�mP'��}�(	�J�����2�8́���#��ר�IO��P!oE=��s�j�&]��G��97�\t�=�}����nB���~��|�D]QS̟7���t�d�n��� ��i��H�����O5�n�Kt�D&����+�*T{czqd�T}w4H$'}�@�oE-�U�9�r�A��"XA�k���\�:2^�ӐL��Rr�nkg)��v��<>�M��~��(�`�`�K�U�y=ݚ�$�V�'�H�ӗ�T窉)���&3�+�!Bq:�o�,�&`!U�c�4��H)�l�'�oE �p%M����Q�/�ĎVSd�S-7"�:�$}(���Q�0p�بu���T�uW�$��DdvSmBE��,��{���̮���W\���[4B�tg�{�S&v�����oz��l��%!�CL��T�d�C�ίV]�<��A��;o2�ĂAY�R �}�Tw'!�ZX';׶J�F�o�k_B *�\@{=%I<�˚�3�æ�N��I�M�rt�b���e�Bv�>��8��+�PEc3(0�i��gq�Q�mVv��օ9���;�6�nf���ɲ�p��7\vv�p���=���1
M�g�<��x����\�7eۈ��'Q6�<��C�y6n�᱘Xf��b�öƘzuҊ{���nM��:��s��o�|����too=��{��˸M��n�+v�Lj ٷ�����;v1yJ�4������v�ۙ�;;�FϳeW�;D�;K�-,��uV�'\�����r�t������~��L�*����m�UIn�H@��{���۽��fi��>��� �>��0(P����	'���>錇�����td	��:��+9�}t�����įЂ��MCNE��b>$���Ii��ʘ;*��]gmx�AW�R����uX!H�8���D�g]	Up�r�w�#r�%I/����|"o���c!��I�1҈Ⱦ�ڂ�1 Y5@��uP ���2�*�յv#"^� ��;hP���&�T`�{U�8?�6��S�/��C��FrKٰ>�sqV���;=�ݍ��N1����O��0�����]f�
 �bo����\C�����Q��g���}R����T]uQ ����Vj�g��ؚ.��'�ب�K��%Y��_��n��3�{��o��r�l�i�^�YA�A��8͕�r7n���R���2�o�뻪�	���'���Î(.��ˠn�A��!52N�Т9�5�1E�v�.��mP$��&3�+� �0�PӪ7�o:!mD�����|O�s���I[��tRQ��b#��+kx3�f��F��sw��� ���c//X��Pb�$�̪ �D�mP ���s�;9�*d�9�v"!�Ƹ�dcll�턵e[i�l�.g<s�X��nYӲ<b!���m�(#��B��dp1;�4H$��R$����V7
�@���$���$mp1(j$5(�;'ǻ(rY{����$�DNwW��O��*���@�����+BԎ��a!6r몉$��r	$��_'QQ:C��9"Ι#��5-��c�;�\n�p~�*�ީ�{G���{4dv�"h�N{ޞ��}��^�/x ��\)�&���$���
 �����1�ʈ��8j$d��]>K�sm�O�/I�=��4	!nSO�w��z!9�M��Av̒e�Ux�ؕ��5
uF�-�'�����Z�{�ĕ�=�W5�+2��.�zh�6�F
Ӻ��.��
�Rq;���U����D�r�&a�W�5<��Fu�F���3���e�q5�<H!^ӟ	���6��%T�̳{�7���NNGe6��aɑ{w��Dxʜ3�7�d�[S�$!vԉ�]���ޘ)���̊�
��OPI��p�AJ}��%�v�A��D䒢2�_<��@$��r>'��z���Q�DÃ,"�e�Uat�oN'Q&^��㧀�wٵD��D�u�;�g�E;=���RC��f�J�����h�PST[� �v��׊���w;ێ/�tp��d����	�Ӂ+���-���� �e�eDBE�q2Nu�A���uj��^�5�Ī��$�^^mW�$7�Twe��Ur��'��3T����8����XL���#�n+a8܎1ۄ�����A�/�u-�8�u�{-ω �x���@$�7�B�HZ��������BvIq�
D�ge
WGc1����C���$���q�m�:���7z�נ�d_SmAA�,��}y�D�;�4A���];~�K�ͪ�>$7�TO��&N(i�D����iqL<��k������: �V�3|�nԕ�j����O�rr��vф��
U�]U�H]����0��m��R(�j��>+zX@��=�Qj�,��%��5���"�����{77��ٸzL�H=��H{�@��Yov���۲bl"{��ǣ��u&7o�T7�^��M0�-�\��ts�	�y@��E����yw�'����<���y�q�[����� ���Ĥ�Io�����=�;s���pWY���i{[����J!�����෧=�#HFs��n�n�sɶ4��y����rh��E����ۋGm�����hsŘ7f�`�-�RX��7�y/QÒ8�eO4�=*����Ƿ�n�	۝<�y���L�p^vZsqEn���1]U����"]t��)�����jQ	"�8�	 ��m
�ݑ@�O�ޙ���Ue�U�U��f�%�aW�Ԃ�5�[�7� _�'�=�ns��=�h�C�ݪ��oK�A ���wܮ'o5>����`�6Ip 3
D��ܡ@�}.A$�����
���V���C�ު� ��.A9��PW�0�d���[wU��[}>�V�ȟ�Hw����i�6���oX.&�k��L�Pӆ.Q%O[�I �����d��p�"'��Q ��rA$;���\�bݘ;_�|�K�V���n��ˍ;���ۜ�5����m�/ko�S4�bI%Eo����O����<�� ��c����<�ޖN?ww�(Pf�\c�V�U%I!�o_4�w��|�^��!]\8��e����C�Z���I�6�Q�C}ic��V�ÖMX�Uյ�N��l3._E��8ܑC�I=h�ƌ/u�kg�$�,ɟO�w��D�ST��c"��z)�aV �.���c�@$��B�#;�Iz�ƺ�<H$��r%�wM O�X!M�\��n�r�K�b����@//zh��u]�9�ЫnN�$�_E7PF(M���$9��oTm�j���"u�� �Y�^��uQ��E��e�pMCh �!;�̀�>���p맣gtmoT]�v�5�i��Fɞ���դ�0AMT� �]fu
>$���n�uV�x���C)y�� ���j�>�g��pa4�`�q�N]@tٽ��Vˎ�|>'ϻv� K�Ϊ��'��}�s�A=F,YJ ��M(Hɉ��9�٢I<Lي�b�4��6��m��S�}���{�����w+O�h�q.~�U8.Ń:�wq��g���������-+�I0�'M��+�[1YONnkgm�*��R��,ގ���Fk`�(e��5܊���j^(n������m���`&飯�f��w_9p����Æ���XA:�aѸ[Z8.V�Gt�W���3RcjP3��Ú����}��rޜ�t� ��L��b��|O-��pO��9�OS�����N#�C���@��^?�<Q�/fZ�z��Z�g;�5���䅫P;>�b��!Ѵ4�d�`��Z��_�8��(Ӫ��M�O
�"͞�vQ��}{;��zvEN��@��=˷#�o��2�����?y(ϚX�|�Svv����fB����m�az1�p�F��;����js��z&���^s�6��`�֕����Ϛ����6"��&��{��4w��xYl�Ģ��|f˒{�W��Ul�sy�u�6��T�1T�ذ�T�.�#����sV*da ��P�1:�ǟ�yoe�V�fu�5��)�Ϻ�L����F5Lk�+^��$�t�z�K�uͬ����Q���s6cC�qv��CӦ�Np���<�a�S���`{Ɋ|O��DnR��������܊�ط��7����u�١ }Y��ǚ�a+wYk��H*���|�o�L>:]�;��^�ɴYl���9Qs��i>~�k�=��=:�{y��>��`��-Ղ�����)=�|��嗣os�`K���W\��h�m���v�_���\��<lV���̲�B��X҆��"օq�e��r�Z�̡�a��c"�A�q��e�3&F*�j�2�֕��Q�j62�7Vb��-�Ue���F�Ur�P���TD\�b����cis3�֦����[+j�D�mY�3*�!Z[)m��Ɇ�X�S��iV"���nRٙ�����X�"12�nP�2�m��s�#j1\�1���DE�V*�J�n�ӬQS�QC0U�-�����2��-��32��+E �U�%f8S���U0��QEKK��YF1�պi��'`�8�	��=����^��ȥTZ��媊�����カm��1���(֡�J�#\J�kj�V��cF�1������Z� �F�F"�m���\r8�Fe�e̢�Ĩ���j1EcZ֕(��-�����ADQUF0cZPAV%�V��0Xc4��DPĪ�Q��3���gl���Ϊ$ׁX���N�7َ"4\��a �>�A�sv��V����7�O�e���b	�L�jn�G}[  gݽ�/�Gc�#����mQ �V�� �]>�u��8˿��;3G;[�fqֶ��}��lpn\�]e��xJ	n٬	(�EC�gG7PF(Nqܾگ9��	���ȓC*=ҧ�"���V��@'�sv���:��SID���w���e�:�]稒Hs��@�I[��K�M�3�ـ�����a�����sĐ�e�$�}u���ƌ���$��ڣ�.@'�F8YJ ����$d��r���ӭ�A��ɢH>]�>�]��f�0��C�FH9.s���Db2��J�D��[9�HԵ㞢w�&����?l�.A�q�����/U�z�������[`�[��(t���-Bp�뷄�^�uz����y�,����+z_��;��Z�
�6,���>�dB�j0�J��)��qչn�\��nǞ�vV�.�'��Y�?6����jCo�ӽ�^$��e��|�ޑm���s���ra�ښ�J�>'�#�S�	�Z5@��mz�:s�4E�˜j<�����'Ă@Y�"I�oH�����=[����u��9A&y&�&I��@1;nI:��i�K��fU^���� �.H>$;��O�И,4�`�Ad�Vf�@ꑷ9׸ �\�A}}�^$�=�P��[�s��H��x�\�'(�IB)�������>'��n��4��e�^�H�;k�糪����3y>�FT��R���6K`V#{K��a��AάB�/�ij�A�m��N孳׻m�Fd��D�=���X���<����D���q�\k	v�E�8��a�������:9I㨦�1��A���v�/�<)Ka�9K��84f�e�U�q���uО$EM�s㎶�c�v�5�u��u� ssn���6�$Kټ�Aݸ�od�����r�8;�b�� u&��t��M�v��9ؑ�FwH�k&J9�|�=$�m����b6tiy�^��:<�c�ܗn�Ft�����F��v��O�L�(���oj��Ȁ�j���o3�H}}�O��uW��,0w�s�uR�Ho:����(͂�\����+���9�����{���{:�x�[�����v&&�]�O�u6�!�KF��vH��7���Z`�g���U��C��^$9����:�j$�Q �����꤫"=����$�;�TO�[��w��F1p�󘙝�;���L4Zh0P�8�g�v˓z���ku�-�41u7u@�C�Ϊ�[��ak���ӡ��ۡ)q# ���m�q�W.��q�'.̧)v�i۳�w��پX�ݎ4������SI�f!���(\��� ���;�CoV���b_MU|Hs��}bQ�ӥ�^O�� ���l�*L+(�).jՇ��Z1F_NO�=�w�E~^�o9�;F���ǸYqJ:�;��Y�/�� `��:�r���A.oz��I]��⯤*a�.�v�F��y�G\��!�%1۽���|H+�\��e��G	ī����u�T$���rr��!�KFh��nP���MZ*�v�6h	�!nL�"+7�i�QP�FO^Ux�ěP�!&R��r	$�omT�8�Lt���J����IW��	�VwU,����������;n��t:;`©Oa�`\U����|�n�Ų��IpQ0�]��t&�E�X(FpOo���l� �A>���[=���.;2GAY��Ċ�)%'	�f!�1=�^�f`�Uc��Q=Y<I$��2$�"�z�Ĝ�
�}��d+���ji���> ���u
懵�.m&��Law� ���{3�S?8���2*���FR7�i��1�����z��N����8��Й��y7e��ɝ�	Y��H���}������mȮ�����̶,GE1}7D��=r	�c�6kĂDugW5D�q&�T����>5��p�i�%�4���A��� ���s4���	�ѽ�U��ugSJ9gj�u�ۮ�etE����&:�F�í��{6v�Lv2]����ؓΜ���Ͻ�\u&\I�����s��Vn�H1՝B�%T�$d1�f�\˟y�D��Fzi8���]8	���[�X �����lf�Y���TJ����;�Pp���bz��WV����Ź
#y�H�I1��T	�՛T	/��f
p�BM:�k��9��{��'��*�$���T���Eo�?��,�G_ô-p���3f�#�I��B�9��[ z�a��͉ܳ�.B�E5y�"��Ω����ͩ�v�WP�n	pbs�� ��0�0Fc���UDdu�� ξڢI��~5��9\�LƋđqi����Ϸ�Y䭻������	�q�L��������p�@m8d�+�w���I�{�(	�t��K�k)2J����w6��;TH$O=�|6�8�.$�Q'��N��W��Ge��N��I�&pѨ��B.d<�Sդ��F�i�
��.��xt�$
�����m���'ā79�s��"pk4���AhiH�;���S���m���o00g�r�H�����΀��&���˅pЄ�Z�:u��`��g�`�VL�
�Bھ�P9�A�����A����ۡ�fy]�o�����@L]5l���;#�f󹷺�)�=��s�;L��9$�������|@w�77b�u/�,E��k�2�E���T䣮��M�V3+mЧqs6�q�]��|;uڳ��3�f�x�k����u�ȘrZF��[v�F�[�-�6�q��s�G�F͸x@�"��N���v�Ui�u{Z9�ik���w���ȹ��Ȗ�\�ɝn݁�8���ݶG��f�S��@�o @�W�Ş�f�x|6�z������i8Hѱ���\�h�����=E�E7n=T�XoNh��v���r{�����c���T�D6��2����ɆA3���9�n��H9)�Ɉ�گI���n���Ibl��uxQ�P.��Z�@Ֆ�7'����1��T	���vZ��1Y��ޓ����pX!&R��qd�On�{{&� ̇<���':a�	>����etCh8�����wԪ0��)���d����H���	����gNf�[;0�8`�v�f�P�.Q��j�g�vh��}$d��$]fP�L��U,�Ѥ]������������z��Û&uۙ�#3�5�f��r�v�u����6�5�����]d%���N�p�Ln^Т	��u{i�GV����q�?A1y�B����H7�Q���ܪ����9�}���O)twxQj����N1��csp���5�˧�����}�> c��Ν��@��,���j��B�Ӛ��rtչۻ8/S�13�lp$	�n^U	��gP��%��wCp��$\��p�7
��}��@�;[�@�O'g:��;�H.��hI��TvÈ	��e(�g�1E��9�x�;u2P$�eexQ$�&�v�w�6&ﴋ���`B#{����3KbA�L�Ps�Ӟ �ه�	3wR�A>�ު�L�gMx�w�]0q�ݲ��w��G�x�4�o�ݞ�']�u]���
f�;&c��#g�����m�d'\���sD�=[�(�F���wPT�;�(�3���V�P$�7[�^$z��
�L�$QM�c����f��Z�鮢	.�E�1�t����3:	�UL$��(����nP�H�a��3��)w�|	$�s|�{˞��^���se7c��6�:������{�l�ܶ���p�&�����/Ub�2-Nn��v�Iޘ`�щ��6bċ���6��̾$��d�$��,2Au��c�Q���V]Ux�6�LᆜI��>��	$��Uc0_<|�;�Z�V8�WuQ$�ɆA'γz��٥��C�b�`[��u��ݷN�l��Mp��@�٧	L�8�z��4�ف���؆�*!��x�}U�A�O��z������3��}O&� ��0�3��6���҄��W]Q1N�T"�ʞ���|A���|�7��$��w��y�w�s�բ�$��Zs^=u�|\�t�$ݘ�Xq�:�} �L?I��'n	U0Q�DCn_f�wt�َAU[���D����$o_V� |��~��֟��
��EC��CV{��[�j��[c~ݹ�Q��p ���9y�ogH0�P��z ��tՌ"�nH��r/�'����P�Qb���mz�'��oM����Y5X� �^�uW��/�:��Or����~[��u�7
��8�&��ۣ��Wi�[s�e,)�J��SZ�Ggg�>����~�$�BM�5�� ���T|H'ϫz��q[�"=bX1U�^_u��tCi����w)�U(9���\���U��	!��U A{[�^$��"#g�I�ɵ�X�T% ��܊�v���u�#�,��	��S��T	'��,�:�� �l}9ު�@�����,��	97B��$	�ݪ'ĝ�+�m��qd����x@�-Z�In�m�V�>7���(ʈ����t/.}�'
	����!!I��!!I��HH@��HH@�Y!!I�I	O��$���$�䐐�$�����$�䐐�$�����$�i!!I쐐�$�BB�����$�Y!!I�d��	'��	O��$��HH@��!!I�BB���(+$�k.no< $;�0
 ��d��D;|v�QU)A�UR�(���*H��J�%EH	J�B�J���%*���� �)PE(H	) ���(�  7h(VR���Qf-kMKF�h�IHSZ��`jl���ݜkMkl�j����mi�5fڥk3Dm���[j���Z4kM��i��                                             (飼��s�p����v������빾Z][m��>�)��;u��H񷶱q쉹a]+j� n���n{t����oP�M�i[�   ���p�ۛ�P�p .�nm9m��*���]ڌ�9�[�4�8 �
��1��hY�����G{��-:��I�jkZf��   �        >�6����ͪ��B�ojTع�]�6}� {��Qnn>�+��M&�^����������� <��QVa��(�U/zT�6	p   ��� M�� 4*EӀ ������l|�	O��U���f6�T#�� �
G��W��@q�/�P���.`��
}v�d�"�M.   <       ( T_g癡B�F�}�t�{��f�/� C �Ǡ����}� �>�{�
� F��f������  .�|�:S � u�g;z�a��5U���N �-D�z!��В�Vl֥l[f�          ��Y���@bh ϳ�p 8 ��$��L�N���t�  ��
��'�r�eJ�  ޟ ��4\ `&@M�� 2 7g �n��������_#|���l�e�V�           >�������֯3B;�4=���f�-�׀}�y`73rґsd��gSy�A�c��Nƭ� �����0-�1��B64���  |������WD�� Zu�S��6�\��5���U]��E�=� ��K-zjh�[�z���	͹�Ҿ 5<�Ғ� 2 T��JUM4�&COa2�*����COb��������=�'��U4��$ҁJ�  b~������o؎��o��?|ϳ>���L��>����@�$�{���	!I�@$$?�B���IO�H@�!$�	!��@$?�ฟ���?ݾD��7�|�e-'���Z�6�%6c�5*��W����|�I'�y�ϳ�]�6��b�c�)�׋�n�J��JҕW��k�n7�Z\j=�1��J���FMۯt_Z�H�p4m�m"�њ�7���E���~b���ʃ\�l�.��l-Ҝ$Q��b��ڨO��Ɍ�� .�)!�y,;���ҶR�i{f���Nt�E�,ཐI�!ܡ��h�^��x�K{ly�r��k8,��k�2U*���dO�ɻ0e�H���B7�uͳ���Ku��U�0����9����+KZ$כ�,;Ϛz��@7��J�|���:W�- ��Ix����p�̭��z0�Ь���K��8J�URۗ��xY�c��J{���\�䨹��/���KqI�ֱ����T��"��0��3�lU��s~�&�Y�nj�7�F/�=�M�
�N�(�8��qL0n)�Ѫ�u�3x��c���mf��8]�:3Tz�8wmYj��eu_��5�����8Nw�ܤ*�4\x�%W���"�:��s�+.t=:�v���3vz�����1��v�m�s�S���WoL����i�Mc��㭐n��{ݦ�Հ2R k�~��\���N2����{SI^8=�%�0��da7�������G�v�;_G6�����4P�n�ȼ�f�8ctov;j��-�`�L0�msv'%��ȶ�Z���J?6�✔� LW1���� ��np;[���}��z��sg,k�vr�Bi�ƾx�}&��&��y6��'�E�!]GU�ƬX����X:�cA��@�.����mN,�����1�r���Ĳ�3�jx=ǯևN����i[)e�OYq���o`�.�b�ow���j^��W*���J(�G�k�Yy8Xy���� eUW1��3C<v�s�����(���L��H�㧰�ƘyH}�����gx�{=�믐��c�XS�$V*��p$��:
�Q�[��H�E�DA뗦�
�� sbZg�grZ{���hb���j��j;�¶��&��r o �D��HE7��ɥu�q�X
Z2��GWg>,��1d�^,�����C�h����v3�1.<&�X�Yх%R��m�5j�����̬e4�{�ؔ$Vl��^{9s��E��7C(N2�}ؤR��kz��{�
�7�e�8������:�E�w�F��8%����X�ń�~�ƞ�(؟�q+1(��V遖�<���2sQ���ga�׳������=jwPœ��ZjB#(koR����9���I3��F(�(����W������f;h�����UA6�6��-X2�Nv��j���@c��7�e�{vc�62L�>\s{���R?ۈY2�
�����m�czLl��Ӵ�KI���p���}����p��m�7�ný��2DBb�V���8i�Re5Z��M����j#m��#��Ip��"4gQ�l�0�\ѽ�%�*%f�@���i��Ȇ��SC����)�������-3Pz�ja�� PT�7��k���8���m�-c�ƹ�wA�T{�ۊ�x��ŻW�[ɚ2ol-'�Ǣ�ը�"��@�w�c)l�Ե%�@�$��
�44��%�e�ki#5��Ņ����A6��z���^��vU��<֞���Je��a&��3O�r�c�[�ƅ�����`$�*�=���y��z�"J�rz����s�CM1؃�i���Osb�\�1$	�T0�xl��>�����*���2�dF�a�_t��9�q���]�� �nqֹ$�����c�h�c	u�Mjg��q�Ѻ���U�!��a�[��''a��ܶhm*��b4h՜A�G8:;ا3�kw�����H�:3u�obg�y�X���h�I�nmus�3��Nli鐵7";8,hT�^�n�6bǂ�]�(��u+D�G��ZӀ�Q��E�,<�OƄ�3Μ8��vܷfL�,9��&GW����rC�|I�/3�̊���ڙ���pc�l�w�����<K��*�����L�dٚ�/�c�����Xk��`<[�NƿX��HZ��b���gd�CS. ��2�%���y���ӻ"X�9N��:��]L����u1��^�nw]	�q�P��<�����n���sS�C���q�٣t�4�ݵV���IP0;�8u&.lG�[F�F�����E������~�^n��e��a�U�*�6;x��&w<� �3�T�4�Rj�EK�9��`���%�_rO&3��[�J��{�����Ϋ6�K��c�^VR�ֿ���Z��	�Z��V��^�H��j��q|2U���6�:��z��M�^��!�/��V��o�I���7v�'K�ۺ���H��1y�h��p��[�[��ZGf�MJ�s�j�X��˸�Y�c,geM�3�.�3�*���+e30^#�m�>���)���V�&!i��t�^�q;�b���t���򣡜KzP�h-Ә_�~�&lǥ�%F�B�C��
�v��"��%$ܫ8���j�8�a�����'y��L��I�9b{�0̂�4��^�ŗ���I �R	P�t�x�n�����ѩE�V�Xw�5��uT���srcX��' �4].�MmRybF1���V�'y��ŝ����?B`��Y�#X��7������	/	��O�窦!`;�v�
�Iҵ��Tk԰b[���
#�;���z��Ǳ�<gv���v��{tC��\�y�l�qu��b��=�����֬ޘ��K_�d{�`g�y绷h��3�Θ ��w;h/kM�6@�¨
�ۣN�8�7���B�Ooq��r�M�۠�(�7cw�sN�w�*Ҷ��E�!�YÜt�Ѩ�f�b��v�Ӗ��zw(�`�"gWˇ	R�����|0�1���#ÇF��T��&��K�h�ǚ�Xy1�Y�_-C�@w�G���s�`��X:�`^f�%	�P�����A�S���R�ݥ��Uе�ye�zU��T�z���u���78�6k-Qy����;Bk�]}0��vj�y*d���r��\i������ⵕ��}�d��A�лϴ�bo�-���9��-��W�v� ���-m��#���qL���M|��"rՑ7�ͦ�M}Yu�1����Θ����n��>��l$ɻ�_��z�� ѱ���+�:�����E�Ό���_����mW.-�(���;�Y���{�]_/'�Ϙ�Y�(8VV�{�P&�h�/��$z
��r��{ax�c��	`#Z�6�)\������(��h9b^�#K���lO7��-�Y�b���5j�P�&<���)�};
V����`�8�P�����P�яI����:���P\e�������cxLG^��WQ�u	@�K��Gv��Z�5��������c����(p.
u���j���-����X�b, ��id�ݡsF�K�	.�#8N��;'!9m�Cxy�`�p�9��^˃ef�w�8$7F�8��B����5wUʙkLr�V���M��hS�d%��4��i˝�.����I�m׬��@�sonM\��)G'+z����m\�W��G=
����u�滤2;:�)� ͝ \�����D���+j��Mn8�ٜ3��
tӸ�}eY�;��1��
K$?����c�c�hU��j�<R��	4�ޛ�vPF��XZY5��}�v�wF�jxn)�Z|!�6�b�	�Z{4<xnv�>���ں��*����wi��f�
O���1���x�7���( ��n��r�܎֫���	]�׀O�S�2���٬�k6�2�$νd��Y������x4�|��qp�	�ӝ�xi���<w`w�y��c{�'��7)�@ ���a.=ǩy���yþ}�rc�����-�r<��5����f!»�i�ӍE�*׌ު��~J�0[zH��3U�`�S+"#7:d����u������e���b�X���Ғ��v�k�k��P�mn�:E�*m0�v2���dYS����\���9�u��=���uZuh��&�.��0Z�%�Os�蝌�ۯ��r��`�h��Q��j�����EM��6���3��nW�F�)��\�2N����
�F�&V���q���s�T�ˇثSeD�HŽ�ս������]�yz�3xγxdy�� YxC��{��Nw�%�l�.�k�rv��O��xrOj��i$�8fۍ����N���4J����PIA��%X�1�nF�%l!��Q��1�^�N2O.��-u�WƆ���f��+N�Ha]ٴm� ���v
:��ޮNh��%ܴE�s��\����gD76BŅ��Ua��"aS�0u�k;��!�y����lF-��;��9�Zw: Kogj8�[x��0bY�n赍��X5#p����fn>ŪT�z�����8%q 7:�x�v:�:���P�<��D����5p�;��vuZ(X��em#Q7��.xsFkN��Z��+��k��i����;Ju���d��>2f�[ژ8~U�q\j|�;��r�f�F#�!�D��z�*?4���Qޚ;rf�Y�q%9���Av�@{9����I<�n@����>ް��4���A,���Ԙ�r�G��]�!�vFA�,j&7�ͳNr��2�-�k5ŷ�by�S����ӵb;�cd�V<���)�%�ZZ*�	�A�UH�v�.!9t�
7������դ~���j���Z;��2�fo ;�j[�v	��4몍h�s������*y�e�8�	���z�VG���җ��1��5�4��eE&1���7��7�.5y/�gzi|n'�ʥ�\��8����N6`�\�-��6�i�x�Bs��n�\xD�#3}�1����C�q�s^o�|��Ʌ�S��5��EL�gtS��ُD�����^l'��{Df��R �X��v �6��l+�������e�� �6n�̓�4!cN�Y��c�_�9������tՄ���ؕQ4�]�݊s&lsM?c��aC��V��e^
ڡ������j�7���ԂT\�i��o&�����^��cB=-�VƉ�������
)����~x}Q:�&7j7��@�j����-,&wt� NC$�w�g��-�� �&�iIAϬcA&��V�=�Cw��MX|N\��ks Z+�<�1?]}��34�4�˱I��3�I܀r��!�^t��)R>�kOkhW���jDB���e崊�ë�os��n��=@;&$��U�Ìi���U����X��ڮ�ز�ccLM�����Tb��"a�f@5Q4�־|�&�*f�(���G���t��8c���9z �ȫ4��4b�s�N���%��\�<ᯑ����t>�S�O��ӗn�h:^v7�:%^�(�dx�SG;��������c��v�r�]nv��*K\WnR�e�:iʹJє���D����2�srcr��k��A�7�`w��'��<s4DL�>�y."V��7^Y�uf�&����1�Z�f��]c���y�~3���`��w�U�'؍�bܷ${u	Rս�l�<�H�y,+��ĝ���yߒ51��nƒG�L]Ɉb����7���܈.y*�M്�`�u����#�鸍�8���pZ��כ��{���(��:N��h��>��Kڱ�TZ�k����Lex;9h�����v����n���Z���֬E��Ok�xU�Oi�ta�-����L�[d���RXm"J�m�6<]�e�eh���A\5��YRiO.:�;�#R�E��������ZTE�n��@�l���rF�Y8�u�8����z�<g�B�[lø�9V�����q��9�f��f�e�nJ��F��g���%�y� L"�t��K�1�*�E[%3�S6wN:�.kR��V �qc�m�Mp�ѥޣ,��+p�����f6�	HR�{9YJr͚D�`t8��gq�i��z��+�����,nvL(���C��N�w	�(� �VD�3��R��/��Z�n��w`�0�6�낧���X�@;gU�})�s�o��m�>я&+��ȑ�m,�??�O����Q/��K+�w�;�}:'���q���� �Gƶ�#hC�uŰ�1h";��P�oJd��B����>%��J���j��S�����LxWB�4k���Qd�����~Y���oq�3�1��ޘ�joU���z7ЎYE%6@ٜaы�n9 [�O������{�[Wv,�����Ҵ�k,�F��Uk�Bi�w8UHٜ&^���ȹ�sYRd_���|��9�g�+�ĳL�?˖���Gт4���:c
\�1�H�F�jsR�qV��,Gt�v��DaY�%�Xu���lti��\��>BP$�� ,��IT$����� � ,�(E!��A@�BH "�H@�P � $!�T��Id�I!�+	��!X"�H���BX�IA`��"�a
�d$HY!����$��)I
I ,��P R �(Y"�H��IRE 
� T�VB��Y %H,�H�Yd$�� P��*��@��H@P Y	
�H�	*��$RAHI"�"��! E�B,����@�a J�d��B��HV@�!�	 � ,$��	�HER ,�R�P�!XIP�,�H�!���HH'�<����ߨE\����e�S��:6[8�,ֻ���/n"��Z�x�eMX�{<��ŝ����ݠF�)T���Ou�xyB�=�ȸh�!�~��`[���'A@�B\É�8�̱�H3�_�,�q�,��ͅ��	�:?y\5JSS��ϰ\봣�8��v"��\gT�g_/
��J|h�����5��/K��}�����xr��ShR\�m�=Ȟgרƺ�?���=M�F[�,ݥ����0�cUa[����Z�����ʓ�6�~�����jv�t�x[s@z���[��z`));%ț�x�~�౗�s��༈��>��]oS1���<u�}p���ᓵ��sc6�-��uꂙX0e�'Q.�3'ڽ^��t��ǔn%�d�2�t@ޚw��Q�z��&v��A�Q����-�g����hֳ٠�z�ld�w
o�A�^�C79f�}���&D���,)�t���e�䰏b���j�����n��7{s��0͏�%����J�mx^��8�� S�/���r�}���W;������s�c����YZ�i���@�6��8��u��'ьk������A������x���E�o��s�Y�y��<�/�*��Spb�Aw:�.�E�۸�P7_����,;�&�~��dh��O�a[BU�rፌ�/$	���2=
��� /┧ e��n�a!����Ҙm@�}X��)�Bv����g?_lY�Dg��i�������|V_t�O4S����HV�m�/,�K����{�˅���H����V�����C7A�B xg��6h�Í[;���A��d�/|`^����í���-�`��&#�/n�#��r?ó��=v�\���m�_�� �F�#Yy���|��u#	Gk��ث<;ܳͬIP�]�t.��6��u�[Ү:u�pyL�\�-�����M�y��3��W�y����Y�pW�9�3 ���/���=�������ώ��q�.�f�8L~9ꗶ#n������7\cR̓�pδwu��B�G���`s�F�Z+qb%;$Э���pm뫐��
�+���e�m�i�y�����S'��m������`���8��=�Bz�yx�7��V�E$�6}��h��[|O,�}�`��G�zv����BX��X����wH�6�P/S1;4%�a��v��b��g�.1OB=�b��Hz���qh��7�C0ܓ%m][��5j.�8���\����k�n�q��F��ƿw+�s�]�7ok���e��� �q����Zr@�uz�0�䅢��yw{e��21,ݣ��i8�k���h�곁��jD�fw��h4�m�q<����su"�9M��<S����.��.&�p&{Oy�=�}��k���u����������5��3Vu7�Gy6�kʽ��y����/Bt��,�c�6����X�^�|�$=;�r����[kA��u&!#@�b��1ec���m]�گ9�ͩ�����]˱�_��燪���A5b�G�eƖ-�+;�7D��P���ϯ���y��0���:m�� ��6Z)�|-��#�P�/=��u?n$__yί��0���r>���I�;�ޤ�׋�V/{׃��`�p��q�8j.H�G�����-/UW'o/E<*4=t}���Su����;��Jؘ��!��v�/
�,����	��ͳ��oF�%9Ȋ�c�.�ō�]�.�
N�^�j{}� �ww�X\S���K���if��	g��1��o�zL)g���ҥ�{����M����.�_���!6��������gM�{RE�ۯ���u���"|���d%��
:;)=�~���54���i𰙂�n�P]�������Ð�D��]�?�S��h�ϐ���|��� {�!'��gC��W��a%���ᄦ�y2�n��Kp,<�.x[:�݉g��=��΅�0��{(#;;ئ�&2�5�s�-�Χ�ͯuft���h���4�nH�I��5����nNW��]<�4����{� ��&<��)~�����G��&%7������%���Z�I�����3��8���{d�"���]��%�eh��0~o��=8^��Aa�]F���	$2���M�{�C�T�$�]qd���i�W�q8'�c�v��o�JC�w�iQ&.m�hx��wFf��MM8r��r"5��N�����!�b���\5��\�Ҽ�w;���с?x�N;�|B�n{gF�<Nm���U�]��z,�����,�ٴn7�y�ܯ%�������
�(ʑ3�`GM�	s����,�F�{�z�}x�m��x�>�*1Q2��6e-�v�z��gr^ަ��?M�O{�ATM�*�Ϯ_�"�w8T��^�r�":��͞V�{��c��'LG}���X���S�z����;G���u5���D�f-~B�<�"�}o�o��&�!y�-���j�����W���U|<Z~/#��Q�u�:[}xƷŝ�Ϻ��I��"b�b�����+�-#��j�)W��9�8}
�6^*b穮#���B��^o�"�f�y�h���a��DG�K�-��ILn�hAw;. "s1���>G��}�L��֮o�h�P���+aƋ��֜6.Z��,)��	a40^\^ja�8��p��p.�nd�:-[���AN�J�����MC<!���ֺ�ugZ�S�o��Ǹ`k�'���)U�M鷇g�}�>����V�&Fx��_p�Ҽ��p��$]y�㢅�nчk-5,ct�j���'[:���b�l�8���O�¼�{�jz}�&^�ת��M�~!l�֎�h����	���Bg���lT�/l�b�,B~��2Ê�]�ȓ�^�#~`h�H��v=��EL<�q]���,4K��v/湉��������E_1��s� �-�5y���9�x��e�uv�P�+����LXi��u�S!�Y(�4��q=�J�ё��Z�w϶ѣ9��Y�rs3�{�pA�G�N�5��8�P�}���\zfDvs|�+���� ���~\Ԟ���)�'9���,��'��x���yK�񘲟qX�B~�p�f�M4.;_�����l�SPʀ�n�Yt˼�jq��9�3Z��a>G�ۍ�E��N���JƲy��d_BJ�ȑ�	 }w� �ǇbD(׫K��q���w;|CzgP�Cj�� �����=�;&fʡ��f·/`�ː˘��"m� vUb�aǝ{���e}���z�����-{o{)����	¶��G�g�L�2�Ța��D�Kx��w��|�ME�0�!��*qb!�PY4��1�*sy>���}����3�X[����cU1[k�M�
޽���!�ɯp�On�"�5
z��O9&qA��Z�����O�\ۅ�N��o�۔�'	�,A���D�5d|� 5~��L�>K"�U���y�������z�LEۢ��煂d����?o��.д��=�F�b��\�zj�t����F����8��D��ݎ�Uyʼ��A��¡5{)�K�R1J�9n���7�{v��q��_u-͑��M�P�LBu����MG��L�/�#q��>��=|�J`�����yH��>CE���*��Og���@�����ouC����6zc���a�eM���P#�*���䟑7-��sn��N�M�ۙ�P�hZڈw4-�݊����tn��l�3��[�Ǽ��xxU��������^h���%Љj�Ӏ�31�[E��rL��c�Ⲙ�5q�7�|mNG�6Lȥ�����<cE<���"3{풥�fq�D)K �yNUdS.��7sѿ-�*���.k�o?x>O�W{|g��_��-o_?Gv��u����B����dd̡�i���e�4ͤƞ�q��Ϟ�Y�&�Y� �]�>m��U<�R�r(��X�>�W��cT�T
×EJSD�bL�!�0����zY�<�BzZ�A��ݞ�_�{g7�
��W�m[f>��xd���n.C	{˧]�l
K�+ɞq��Y��2/�C�M,�~�++�g���#��G�Q�Պ�w�7`����:��j�T3]K�x�ÐFg/g":�.���$����}��o�"Θ[��L^ãҼ���u��1�o��½�c�;��$<��s=}��Tu���� ���hs�a	�6�Ǎ��ᘕn�F;�ԗ��ܜ�q]7
�߽󆬾9>1��m{�7h
�솄��V	sU�cV`��̚�n���,���ok>=6��ǖ�n�"d�d)��
�XG����wGb��� ����G1�u�<#�X���6p�<2��,�a��.lI�`��
�X����U3�n���)�K�˶/=��e�����h�/r�4r�~�vk�u=Ic���e�8�*���3��rFw9�0���+�v�G�v�_��4N�}�k
ǜc<�K��p!k%w'�)�Ǽ� �/����~�������{���A��57WE��jL�1����:uv��X��_>$y�}X���{�
~�W���lAi��{=2�L˾8=��7V{�`�w*�󮇪>�LXt�^l3�K3�vG��=��#i~�������{.�.��;���~�Km��-�}���'l��$.�Ѐ�[�,^�\���q��G�H�U{�tk���!^�H�Os5�ܦ4xo�u���a[�3��V�a��騸D�U��4�І�}�t�7Dy��(`/�v��s�{������[+�{p����~~��w�M�~��$�Srk�2� P���	���4!��0ȧ
yu�A1�;�aN˫t+_�3X��[��/9���>�#](7�ֈ��C�f@�Z~�$It�b*�QP�0¬��QI���.�%��5��Cvv�TDǂ�G$R2�ǲJ�7�s�^�WC�8{����c˚61���s����T�:C��嬪���{*����vѾ}{:�F�y"�`�ʩX;�����?h8�3�J��w��*�2�����u���ӽy� 3d�^�%�p/0��>��5.��p!�6��ur0S�o��,ް;��T���d�6�}�O�y���I���������97���sR��]�p+��{�W����\�l�3S�a#[���N��}�8c{�-��s�N��`O��yJ��S�	���j�7n���'rՀ�R��������OJ]��-���M��\�����^�_�� �9(-�s����]�^��_L���G·�׆'�,�2�pP�PY�;�i��DMãX�� ��6捴Z��P<9��\^(�=�:c�-�wh�R�@�n82 �:�+��]���Ѵ����'��s�x�.�v�����E�$y$�}�����뭥���΋�bGǜ�	�Jʂҳ6H:�ת�9�N��AN��k��x.x��nx !%���`���<2��O��4�m�XA���e�1u�Ų��x��g��,�=�0E鞢�.��9�E����� v��p�{;��0q���M�"�Sye��zhiQ������v�)+~��B)��(�No��#�<[A�vў�R�L]k�}��7&��KVzK�[7��^�\�o{qs9����*�h?{��/ͫ�I��zt;>xz\])��B�y[�^�M8��'56�n��a�nn�Ý�b$[����e����G�|&&�
���!�{�y�F���OOƩ�tG��Y�DX�6��zL]y��E�ظ&���X�s�kgv���;�\DwS�2)L����sV�s�0��?|�����wU�r�8�>(�'�3��
%��u[4t���{��f''�z:=���i%�04`c�d��{�����+�]I<�xx����E�X��k��q.轑(q8�^����mJ�7�>}�74OU�B@vV=�e6�i�&��
����E'�\��U7�pE��C[
C+.&��Jt�Ǽ�A�7��ePG�/x��/��Ǿn�@{FV=6F���)ȾT�rx	F.[��=�������X���3�3~y�X;j�����uMh��g��2�w��ϋXW��=�L��$ksg	gi�e˩���&�kS
��+�R^f�*^kr3��ѹ'�p���&�PûݞHi<��U�9�o��}�ɢ�>P��?n���C�����!A ��{��Z���u��]r�B����<�,���)-�VѼ��z��h�Z��q�W�~� �
f9���x|lj�;<����n׺�C��o}��P���=<=zf�2�x<^:������Ҩwh	Ŭ@�`�E���\a߫d���@�~Xy���4� �=tz��:��3PoF�Y=��i��g�82�$o����t��;�\O:�F����l��u��H�{�� ���\M���E�8�P�koH#M���5�8n���Y�i��v�^�2E��f@H!��8d��#ӛ�z]�s�����#���S;a铷�-��ߧz���X���w���m�_�º��}��F/��8l��d2��7%S>~��9v�<�=��o�����/t�����?l�����<\��{��`��-{p�}q�ho�x{O1���7���6,;���n����ǘ���07u����Fm�b,ڵ>,�/��2!��huG$&Y�B�g�@ÉNm�
��C��x,Ҽ���z�j�xN(grY$͉����8����<�%z����m����Mw��>����I)�q��d�%�\�3������v3[g""V��`�1�ʹc��;�=	�s�9�-�q�Gi�Clΰ�j4��z1�ɹ��vݶ^��^[�6�vTw����-�B��ێw���^�6� ����Z�ݞ-y���d�&�\�)��F3����=���ƻ��d#�t��^�5�J;1�cO�᭳��V�6��#$J\6�`�瞶ݻ����M��V�$�u��T����m��m{�:�Y��t0�ۜاcy�#��l��F�D�l�{���p��ɀ3,��g����3�_.l�u���Qz���2p�"���k����9�=�7e\\�:�x-x�:R��sڴJ�w8�x�y�C�e��v�)�b��k��ଜ�޷Wgc�mɣ�8�utr����^�ʷ`�oO\q۱�v��b�����ɛ�uP��$�ٻm�%����b"�s�E���\�n���quG<O\mJ�gc`˹�ԜW[f�pfݸN�9��v�r�,f�`m��ڪ�N��sg�V��`�Hp�.4$A��T�Ηs��%�q��\��>�8u[n���^y����N��P�1�(Y-o	Vݙ�/]���7���^�O/lΦ�1�˷c�k��\v9zw��Ŗ��nN�6�+��/\�^�;m8�늃��!۰����[(r'��{���ݫq�9�m�l;q�]{Y.���]C�l�m�F����;�pfN��)��=Ǯ+mx}vG��[w���S�����n�L��n�vܸ����X��Ü�HGuv^0܀��]��z�=h@�5oV�Q5�)�����Ƹ���[a�A�ݶ3u��F�ۓ�&����-�x�6{v5Z{y��f�7[;ٍ�4�;�x��f��ۜ�����W��G�[��M�7,�69�O���[E�{q�L���"d�9�k@�̓��S�Pt�2��J���/D[v��l�G9�*vQ�n���m̮=\�,�\үX+�u�vk-���x�u�vݷt��D�����7`�-V.��Sn6��/�Z�.���<ǰ���v��t����:�7�ݮ��V6����d���r<l��u���=��ـ��cuc���/Hp9T�yx�[tlu=\��-�G��������Iż��Ɍ�5 ��9�v8�z����d�gaZ�a��=�'lku��Y�1�[=�y_*[�b3�c�1H�c�c��m�cn��n-;.�(����C���m���ϲ7j�e�dyv�<��d��;d�Q�-�pWѷn�n����Ϋy��=6�m�講�w���Wc�n�#m�p�����6�,S�ִ���.a��{p�s��T�9.�������7o��`G���o#�:�S^n�I�.ۖ5�=g�H7lj�`7l���;<nX�fw){^�����u���:y�nQ��K�%��y�-��n��u�; ��惰��Zz��Oc	
v蓶�ƹS��{���6��b7��݂���v�����6ۂ��������ݺ����k=iw/u:l��d^�c�xA��<[�CxE�gp��!n�96�I�a�i7v�y7$r���m/q��V���vlp�ʹ�l䘂O�������Nn�0H�2�^'\S�.'{u�y^ܘ!�oe����܀xt��F붩�|����6gum���h�Ґ��v��!�=J�&�@�40��g��&�q�n�8v���[�'�VNxK����3�ъ�a�f|=�r����ԝ�p�]�v�ѽ�^�0c`���]�Y"�v�R:F�����m֒9붜��[��8ǰf.�n8v������WtZ;Z�4�����t��v��v�Fs��͹�&w<��K"u��'�Z�V�g��B�g��
"�1�iR�0d:}l��:�g���v^�^#�A�g�Ʒnz��$�u�X��H{%.6�:�<`�-%�;��\�vuu׆���м�=W�s��'<�N��ӻ>wc��"��M�^-��Ɗ잶:w[z��[��.M�9�m�u�Y�H��=n�Ɲ�:j{/+{v'��=��9\����n�$X�֡�m۲�1��ہg�k����ڮ����仛�M�#�;��������z�H�{s���r��q�$r��zW���ܳ�n�	���-q����cv�1Y���[��k�g��v���{m��nM�fw��t�=g�]�"�n���g��:�K�[�Ƨ�$ܖPn�+���/�c���������gY�ô�뚠Z,�Wls��pvm⛱^�}<xYm�s3�G��:N8���n7�Ԏ7m����%��l���З=���[��cCד���(򱱢�u�%ծu�N6����+��/7oat��ہ�⠺<�"z2��<�k�;���8�&��v�=m�ʛ�9�F�	�G��緲.�q���'�N��$�)�n͸���dr\���+���b�t��Tb���q� ��ܕ�wX<[]4�	�c0��p{[ݖ����v8����>5̼&qq��sĸW�qc/V��Lp�&��N���z7�qa��vݧ]������m��U`�ֶ��r��󛣳:�T�y�7ch�F<���yM�Y�|�+�p�,�+�-��ܵs�^:��cof�;�5��g:��[l�؅m!ˇwn�A���\�[c���:S����ۇ6,��a\͇��4�� Ka�@������y{�O$nG�:Kx�;�y�Ro8�9�])�qѱ�J�b�׀_7;:�7Z�����q��m���mk]>h�,�&&��r+OG����<tq���!ȉ�wF���k���v�SF�vͥ7�Q���s�����^(�=�z�3�v����v�`�xSY��3��t�]����d��QD�N֮+w;Y�g[����:p<v�G�[��isy�����œ�8=�p,�t��+�0����u1ؑ,gt��!�8���֍�=��S��c�����$�]�n�3��[������j�Y��Xd��Omۍ����Y�f�2�͵�C��i�sޞN�[�N��i��뺚���z\�����v鮔�8O+���O�5G^�MlF��y<Td3u��Ζ��^�,�ٳp�&��<�i!��u�lbp�j�.np֗�5i\V�od���Ӳ�u�Ӟ:������n��9�ѷl���
sg9���gd�U�!`�s�q]�l��B�l��N�;�Z[������-�c��7$��M���T����{v�&݋Z�v�90�<�.�=�]������8�=��nX�n�Ԗ2=����g�f�8�]N*T.M"�la�qtb/3���k�ѹ��kl�;�x8�{��|U8c��xL$j��=��("�/�x���U�{���ց7Ys�lc8	n4�7vtwl̓i:�l�c����@g����� ks�2�Ol��knK�g�Z훛�<`��Z�Fȝ6���f�l틶c�٢��^:�C��������s�EfM��gs���ܫ��cn�x��gq��<�=;{j����{Y��m�L���>yU��M��7�k����v�.�ݝ��t\vG���"V�H�HS���[lv�����%�w���5��G���SgtrՀ�s�g�w�%m�F���Mʇ�'K�llu����7on���c��Y���>K#v�!�Z�'l�*��.�X��wC�c�SB���9�q�c���&�ކ6���r��d��2:�����냒���O+a#�L=��³���gN�wm�����cD�Y4i�nv�t�=�l(��ەy9��[�G��9s˳�P]�h���۵�M�%Os�ͫ��ι�"Zi��t��q�������֯d��ccm�n�.�vv�^��X��hS7En��n�hm�v\�Z�糭�1�y+��֏.8٦T9���n*C��k�a���l
�<n:ˬK	ge��3��F�];6��x��e��׮*y�gcvr����o�&�<�4��˹�DHn�B4
���=��p���,�ɍ�N:�ږv��`Y7gd�ź&�t)�\�ά���ȸ��LD�zýC����sɍ%�
)����v99C��|W[���.;t�]���Y瞈1�;\plK�\��!�����=���ɍ��2we�<{<��vx��DVg��^��x:�9�cr���]j�S����ι���8bYݛs�D��mQȓ��k,�F����>�kh���Cf9^� ��k�q���ݪ���!���}�mM�N[������]3��/������x��{t9���۝ݭ���Su�����kS�>�u%�:ֳ.�7c�"�:��9�<;i�W<���g��u��˂��"U��/�Y�e��W.:��Z��&�u�W]�E�k ��7�d+��\gv�nN����p�I�F��Y酃��Pyc�Mm�7q��uXxz�ͭ�j71�����y��P���۶�9w%7\���8����t�M�uȧ�n���A@�'C�8x;�&��K�՛nd��ƽI�l�k:N����v����k�i�28��a���r�f�!�{�A\�ε�9����'@O���1���G�9\�[��2]�ܘ��k5�]�M���6zά��7=������^ppVz��h�TX���I�5��l��٬��3�699nc����n���9�p��`��+q�11����qoe6�n������;D3m:Q�s���a:�g=��[���zy;'h:{U��%��G>�:����2�g�q��ru>�٥m\D����s�b6h8���6y��s�<'�i����5P�c���]���.׫�)�V�:��Vh����u�6��\�"ʗ\�E��F��U�kk��K�
ݚ����E
��n,;u�]v����-R^z��	3�!th��R�Y��p ݨ��[r\X0�7l1���,Cq<M�u%�X���g�oc���Qm������1J�++Eb�hUk1�0 �Q�iJ�j�1c0���UD��0�FҢʔaZ4[`�V�QT.,��ep%��n[���*,����XT�n0��d���P[K
TQ(#-�YPP���ش�8�)mDp��Q�Ԣ%ekD���ËAVա�Ä���h�1b��,��.,FV�Vj[@�*�%J�m���a�c5����-��ʵ�Dm*��."�\)ZX����*
��T���(�bֈ�։P��1HaG�1dp�F�QD*1��(.)Ja�
ZT
��Ԭ��-�r�����Z�V�+hʸ�0R�JJ�i+m�fJ�J0Xֶ��R�QV���V[Lۋb�h(���hڱ�P��Z��DcJ��u$�ofva�,.��k���X�ݸ����gB#b9��c���t�����
�b.�8�&^�n��5�<�`m�A��u���/�c���%�p�l�x�l�:�[YՂ��mѓ��e�ۭ�\ݹ���F́�{q�6s�u�ó����&�cp����wn�N�>釳׈{�\y�$��ڱ�7:�լ�i�t����kc��a8��;R8ɍǮ��aun��Y�k�3۝��n�ô>���f�6v���ߛwc�p&������42u��n�T��׷+�~w����E���ϥ^8��Fl7N�<�xx�tp����G^�n��7Z眘F�sXkF�1�H��=�:�Jb��h�m�T�5�i��g��M�eo��+�9ީ�xd�Ǻ�m�@B�F�n.��u�[v��v9�ݬ6Dx=G=lm;�U��|v���-�]��6�덓��>+�j&�3w;i��d��8�u�}Ppv6�-��6'�WN�n7k8:5Ӕ�ۢ�N��qm�+�����:�W�.�Y�9���=#�W��=��y��d�g�M�,�M�n͌<N�:��K�l�^� ��f�Ke�*�8��9�+ly�*����O1��G^�؊_	��L����y\�wjv�ہ�2� ���ۅ�n��6��[`n�v���nգ��i���nɭ�lP�㬗N=H�`{r��1��t�[��ݗ�82G��;!e�ؼi�sٳ���f�s��*nb�k8�n}����u\s� ���v����z�������|�2'�-�Y�����g�q����Olļ[pq ���x��bn;q���C+(��:���������d�ޔ��Ӡ��	�D��@�v{���LY�Z������~=�_kHu>����5�c�v7%�5����c�P���oS۵m!�G��a@띳���F�9��x��5�ez�С]�Okf�qmqB�9V)��6������Gm�oo(�{r�q��N�{r��m���.Z��0�M���S�����Us�wgd6Ǘ����� �1ˌgwx����p�yq�݅�l�Ɏ;l<�q��@w#��x ��c��yܜ�cv��
�}�{<�vq����gq���Ǐ<�S��g��9U9�����=��xπ�܀��r��xO��?���m''(7����+��"M=��I!���a��9���wd��e�ܞMM4��1*�'W�d�	'!�b|l73s;��� ���h �ίC��\iJ,7.�v�?��̑T��D�����tĀ�3�k�" h��͏u�t$E�I/s��Iel�(�0eX�1�m�1'��6f/�>	1�T� oz��H$��<���m�};gx��1YSd�;��ՠ��N��_}7� �{��ՙ3�� *k�[ ;��က�mݝUԪ�S���"L���Q�KԞ
�8��n�[�{ۇ�g[��\�$����[�Ĩ��H��a�&[j����"�{n�,�z5E��ǌ�%۝� ��K�&&	�	��fӽ�B�D[�z�!�3'
��tC�A�\���_B�ڙZ�>���f\�*4��=1�����{eY�dzk;��C�lY�Xж��V.�NK~�� �{��Y0i�=�N0�����U(�*hl�=��;��j�'�(����`��ʜ�j ��8`$�mݕeϦH��k�"J�t	:�pt)ʉƏ'X�"PJ�w[�5�U�SY���*��p�S;#	%$�&�V���`�H$]��̽���R��N)'0�C��s� �}��׷垒$�7��P��h"R�cFX��7X��ۋ3��=s�gp��v�q����㈃"bJ11*"r��7a"PJ��y�" ���M��(��1�}O��g�0 �mڰ��Dq**`�J�Lh"s�^�%���H��;�
ڶ��h�%^�<�� ]�4�>�,�K��o�r0�:�`�`�k�y��{v� �#]��	8O�/D�~D��1T7oڏ%}g�h]R'V[�y��i�os��0��o�\���s7���2w�4'��I�EóQG���x��s��4������  v�� �}M�Zi��AT�d����|��u��U�k�U������  1���s;�*.�~n"oμ� ������U�Ÿ���k�"Jms�~`3�k� ��n�N��^s�n�.��y�膐��qo�2�l��a�պAѺ�8������n:;p�Ă2g�U,��s��F�3L�ܹϞ�z��G,*����|{���+�y��1  �߹�N؈�B�ɦ{��d �p�y��`�t��*�!MMI2���m|��b�WH:�'w���I"�\ՠ@ngy�� �뜹�!���7���]�K�QJd���&DA��� A��^�0��GT�z��7+נ|y���y�p��Μ�I�$ ��N:k������ܑ���@$=n��׻VI��^��=aK�;ܰ�g���g��X����|[�q�&Odb�/mW���0%�n���tV��Q�ecC�wxssa߈�>ݮi }�ξ��si���AT�����G7����;ؼ�o{�����|]fSh�[���7�׽�dr��V����h����1okBb2v��c�ܸE�On�*=M�lPA&B$�o�6a#���
Y%־g���^` �Y��wa�u�Dc�u���xZ($�f�Y&���p�"}$��h�}��/%8�D�l�4�ע3�.���@���V@�����/Uf9�8�����I��#�E.֏oe6Aۛ�Ұ�:���u��Q����! /��a'�����;L�P$BP"d�-ZF[�N�Ƴ9���^� ��7.� y�q[�p��A�I~��q�~z��@1>B���^�b$��z�^ֻ̼U�A%�$���I#�~�B 8O��[7��Q���͂}�w>��;Yx$�)�����1|������{�6<����޲�j��l���DR�E�,	tp����зv��!�' ��I	6t痎۞3���u0��۰�wI����k�Y%��v���v�b�����ka8��c���!]5�.��;zG�8��q8��w��7���v�a�5:����tq�m;P�62�Xیvz��5��A^	�.s��r�/8˳��9듃x���⣖��[���kJ�Q5\�ɇ��4�[@e������G��&�]���QH����ձ׸tu�c��i�Sv�v�젓�g��p�]��L�b��hJ&J(���ӈh �����$�.���R����Ŏ�ܚ�, ���V	K�Z���k�"Jo��{�y�%�g�=�cw^������� 5�SdDt�yefdY5�{��X�`q�BO��2�םlH$Iw����wg��{� G^>wd�kΦ�o�fb�TW�RQ'���}Mn"z�x������Y�!$�O�����O;��j������l�%��3=�zF���b�(�W�m]դ�y�j��-�n�_�Z@$��]� �E�y�Vm+-���]�F�F��"�<e��&��՞o4�V��9�wm=�J�M�ɳ����u,) �r�[�!$�G����H$�y�VI�ͼ�b:L��(|�-Y 1�W�����EM"d��Y��l�Jn���G+���{@���i�q�<�q�%sWoh^Ĳ���5 �}M�׮\�qˡ���{��FG���,�^�tXr��p[6.�˾�� y�� ���က���c����n��r������Q�7a"��Ձ�e�ט ��l�w�l�=��ĐKozh�]��$��GN"}$���{7:�y>��r�z|��4o v��� ,��8h�����2͝���a$���i��A2"L�&�76��͒M��v<w�����r"Id�M�D��ά�iǝy�����& o|����\"L��y.��4�=c�����s�u�:�0iْi�}��O��z헵co�Ny����u�ך@������Aqq�Jʠ��tشIC��Y��_�u,) �s�۵��O0qe����0 �w�D0>2����}�-ڂ�T����-r�vLJ@��S$UG�9�����;� =W�0g��v��g@��p����G;�����w��k��ǍM(U־�&�L%��ɝb8;��s��ӯ��Dp}�p��{}w`����B�������Do��^��2�my������� 	���f���k͎f�<���"��W�1C=��v��K�w깹�˙3��;��1$9�V�_]� kίA�T����_��1ئL3�Z�.lq]��k�c�yO٧u�p��Ý��g�s���߻�Ԍ��g�~�Oϟ_�DC��w�� n_Sa�/Y�fv�o��j���۴�>��)q*�Dʊ�"�&�ך�_wK;�}�Y�~�	$J�y٘A"^�M�$�d�됶�扤u��@QS$!M:���I$/s�U���:�ٍ�{Z:6��$�g��@	��k���T������P٭�>&�Mw�gUf��>	��w`� 7/i�w+��D�e��@���:Ly��s���:�/c􊚒Uv�@������׹l�C�h�.qd!x��Z�rG� [+�����TED��E��k� ������VEuM�U��U��[ۻF��?����Z%uf��	��jMH�@�j��N�^�zX����֗x��.%��ϸy#�y� �q�����L�2�3{����/qثH>n�y�E��Q��_��O4o�]ݐ �r���:b����j%Tæ{�)�0��M��/}�u:��Ϭ ��o��ngy�@|ӵ�wo��׊Ҏ1��@�J�fJ&�%F�VJ�Ow�� ���;�׽WJk�� ܟk�@���<$�/�u,)b�wFl�y���ݼ�"��5m� E{�^`��o�4 ���#[�@�>���豾$�'���y��I&O}�?X�ѱ��Ā+�Sa-��8h"��1[��ƞwt�C�d;��5� �3��
�}����3�I7�ӇA��ƛ#DۥڶVL�J���НFg�-��j6��}�A@��з���󈑙t	l;^\އMҚ���4���,]	D[<��=<��(��܆�����om����v�Z�=���9xx��Ņ��,��`q�G"co��åy����ϊ�ڀ�c���/^�|��7����u����{m��+�jw���Ob��g��ⵖ�;X՜x:�fq\��7]��/���#ȱmI�1�6���#��*F�[2��{�~�8�ސ��[��V�I-�sV�$�|��%�z���u{ւ��?����?���KH� D��&ժ��3H�}}�c&��m5�#��h�^c�=��)<|�"�4h.�FZ)���sS]SG����e����UL:g���@ ��w[�A������8�#'	����Vl$��x��'Lt��	QSC�X��j��xld��y]�y�  u�m݁�7s���_(��!�=ėO]Y&��� �R���/b;�{w`�A����$ܮ��
}u�h#/�]�d ��6ON��l�T�F�!I��#2beJ*)�v����i�nޔ��1��gL<�+d	�5���πQ�LɈ�fN�ٮIy"s;�� �('��d�Vc�R{i���uY&�I����B��Ԋ��;y��碝?���o���ft�S�q@Nl
/qլ��l��`hA��ݻ�}�n��!gOKx�7ⷪ����b�xz���J�Z�׮�� m�cv ^�UNrѢӪ�Sq�v��$)4���E%
j�gvݫ���~g��>=w���v� �>3s��Y �u6��=Q�3�aT��ɩ������.�2�"%��n- y�M��׽Vdk �Z�R��y�Z���%$�H��=V�%����#.�t���KϺ�0��H%��7�D��{�f�X�|���꟭R�1B���5RI��Ӻ�q�)�6�7ۡ,j.�E%�[p�O�����*TTЅ|���j� }�^` 5�y�D��c�Sr��ͻ� >��x�20uh�sJ n���x
K@X,�7��2��>� _^�`|��ဃ�7�VT�f���)���""�5�"��A��y� ��^h�DX
l2��1��SS��7�✐a�ҚZǸwh���=��{B��ع���c��Bǧ�w�����_�L��Dڙ骸}Ǘ�c_�@@�tc�"�����q���'֬Aa�����Bs�}#F_g�,��Ҙ���
�esOA��(��l���k[�v����5�GenѾ��d��o��]��;9�ڑ��1n=���S�^[xg��{`�!3��S>�j]��U�&3��.�z>����;��ˢ��h_ST�8�}��mg_�9M���� w&�/�la/A��zF$[ԜX�{}�����]��<�}����e��^KG'��7p2��uR��4��0��v�RM�NҸ�!ˬN<���zt#^����'ģt�1�sy��,߲-�1gC�9��]����7ߡ���m���mC�~/�/iM&7�·׽�� `��*�u�2l� �fU�t/c�S̽������*��8-<`��������xolz����~��#�+�<V)�L�chb���B����ۈװt�J�ɮ�L`��q,q�fR��o��S�!�������c��x�܀co9�sq�6���2ș�[p���SSO ��/�B}\�ӛ�s� /ַ9��ۍ�Wu8���<�� F�D��k_�%*���W�	�Q�w0	;#o!�I�Rop����p�5֜R�[�p�5�B���*�C�:�6�5�e�Q
(w�c�s~	�&?��;C>�����氋u��U�m�-�J�8hVa�D�h����[lE�Z�m�c�iB�*2���#j�j\چ--����3(��%�a�8�Qѥ
��Bŭ��e�-��T�T�iPU�T,�[�U�D�-JᩋEDaR��Xʪ�\�`KeU�KkQVXR�"�K�V)*W0ڂZ�[mj���6ъ*Z+h����pP�PL�*��Z�KFQř�\��$�J�)\[
����QQ+.i�.aQIKF�Q�+�X5��E���#1�*TB��-�F�!�B�R�
�T��J%e�jŮ1���V���"*�L�(�eJ��j�[X�qV�-.s��čj(��P���R�m�0�-)�e��eb
""D��f-p�J�1EJ4�EZ%�(��X�UeaU���`V*�Z�X)KIR"���ъTiCG\�	1sL)�+TX(�X�,Z�(ʔQ�\��,���bU,�*��ѕ�cZ�ib�0��X����*TKe��J�PL5QQb���)*QjQ�EJ1j�BҴYb�KDZV�p8�J�pю�hƴ�j�Q�8�Y�L1"���Z�<޽���h[Ϲ�w��oz��%��_�0d"M-U��]�[�qF��D���L ��� m�nl�^F�$��:�,H�o(�S��&$¹�*�ٻI$Oc{vj�e
w����\�9m ם� >���Y!9N�� ]�O@k�| ʗ��ׁ<��gxk��\��Q�od�s�[;���r��y;�v�i��O��T��*S�sd������> �컰�꙾U*���2��̃��^���U��**hB�uW����~�]秷�� ��y��6����" ��&M�]_s�F������*)Q$ET7�η� .��ڰ@c}��7�uY鸆�̈�i{�v�)�����B���QM�|�/'b| {:o�H }��E�.v�^�_z]Cs~�pћs
\f݌�e�.v�;(ʦ���{��F/+cM�JE��1~��' W5��h�;��n�79nr��7&��s��$(4��!(HD�V���f$�6�;�`4��W��� �s~<�@#7m��>ry6dΝ��/�����/��t��f�qֱ��;�g#�t��=�u�\��b�N�7[ߟ~�2t�_MID�\z�q�  >��iX�&�Ί���" =��vDC=�z_����ܷ$u��J��b
�PȊ'=>�{����܋xnuO{�> >{ۗv�}��o��@���܎��{�����TJ&T���	���.Ղ�m� LP���Eᵎ}vj ;�˿���!��K�����UJ)H&d�uQ����S�%d��ĉ���vD ̽�0 �^W1����S�W�EO�@"�w��*��Ȳ
�"��:��>���K��3.�xQ��	w�wi@\�����|��s^n'�B�x���dk�Z79h0t[�h<
#X�R��gi�DL�E!{K��e�o.��!��o�\�����_�nc�*1�nhP�u�L^27�� �}����g��,Mc�6�m�	��@-v�[�����a�u��..i��Ən��@H	�'�l��i�on8,��Ov^;���J��F����=)��������u��!��㫬��.ML�s�PY�$�.۳�ז:��u��{v�x٣���|�u�8�=����7U���#���86���g��-��v�\��kn����5tdݛ���n�n�;rǋ =�U�&�n�E����.����2�5��
J�K�ws��JE��>h��c���oO��ӑ�t�HA$Co�d��}�-GP���N�^�ތ��Lt]��b�ms������d���͖��+��3Ҫ��u��Yv��=|�RH6�%J]��I|�{�C�oh劷_M�tDG�mz!��{�@'8{�IDʕ4!8���[��3�!HI�F���3��
�kX���ƻ���~�����Π$�'�����}����H�^��G|�K=��Ň�N�	1Y>$��ɫA���"�n]�d�z���O���7۬v��$=e��]y{)�4<v[a�I���L"��3]�L"�(L�!I��#�:��2�w�?� [��w���C�n�N]��),��"Az��e! @�4�ʟs�8��`�"*Jq]S�}uYX��w �Y�y�r(q��G�=�y�e���	�1�Wr�:M����d��%l2��k�M�׹Q�]�w�πA��� ��wd%s�,Su����6N`߯�hZ���iԋ������"I���b@$�N�ХA�vrz;�/7� >7{r�XI�1ҫ�
�A�a(T��{k�`�z����4 �ܻ�9�%�&����έfx�aC�ڒQ2�EMM�M�݀4���9�����i����lR���8 �3wr�E�>N7z,Z-� �D��rfd�fD�����qͺ�1������[9sTvy��C�]��/�1�32!2f!���l�<�9��� �3��"%����^��z"��˵g�������R*+��}>a���Q�̤{�2�� �}�ۗq�'�h���i,��GX<MLM� �FiqP*JT�1��ݷj� �i��mx$L��@��r��zcq�S�5��x��N��y�x�9ˏ?R(D��{�V�X���r����V>S&Ei͍įh�܀Ɋs�x$�^\��2��o��$m��5-Cw�Y��z�=������޷��@ ���j�A�Nf� �/:�틸��)��9��_��ڰQ+2EҩJ��D1���ֳ��l�o2pI>߯ѩ��_�`/����� ��Ζ�/;��l}w�oͯ�|���v�5`=.]�N��S���7i핛��A�v�>u�8⎓���g�����#��MW�ׯnՂ��> �o:���W�c��.���N$�F��ȗ [���)!��|���������������Y{�Ұ�휽���~� xK��7�/ww_zn|�-��a��z`����"��H4���0"2�k� �H/�}t"Z�z�c�+�q�N=��>m�s"�����T���j��{�eq����F�%�Nu���O��m$�wnn�bb��n7s ��{�"F;b?��>��cP���/���湂\�yv>����{���Mů�'��l/��ͫ~$�i���[�1S51U�*�A�����!���7�f�[}t�����r� ^˴I7�m��b�]�t�蘺�\��#���Sd���tn-G#ч<U�������e3^�&b%D��G�fAQ!� �*۟D?��'|�� ��wh3�{�:͛����� Oo�d�wO|�XR���+�ywa�Fml�zg�U];�S��'ڀ.{��C��v������͙���M��&-p�%�wJHn���_ͪ�@�{��d=�ϣ}��9c�=Sl"��r� =��qug����L	
Lݤ���׶�k�d3�I �������� >6n�W\ҙ�p���4��v{�����U51�MC��s�ĒA&���18WM�!�&I���r�!��7`$l�����-��t#�5���~�YU;�cg5�B��Qf �\�e��߇�b��9RܴU�:	���Epb'e�����1nѽ����nV�5n��\�/#�Y�ܛ��<�Z:���6�Ǭlaz�F�;s���Ի<���qێ������.��#�C�~��ګ�k����]�1�ntn��=Q���/l0:�>�-���Y��R�/8�yN�����O&�E�;��>�a5���#C�rj<�莥����d����+��Y�ۇ�qug�y�l�(ٵcW|u\ԕ�������ζ�r������m�۝��5��{<���>}���ί.�?o�����bRI����b$���idl�����U��r��>we݂Q+���� ��� 2�G�z�${�ȹ~�����*{�ݠٻ�l�b���{)����uɒQ2�(��&��f]�` iwΘ�H3gs�U'�N��~�� w��j���Kfjp��wRHj=Ǿ��--����\�#��� M�K�a�ozf��}�$� |{�$̀Ϫ:6|Q��`Z��q���b 2��L;Ȭ貱EB�g� '�na9�,��E$��}pK=gmN��; �k>*=��� TD��X�^�=<d�̮���V�>�B{&l�2�~o�ͿƳp�J��?�:�� iw�*` m���x��f4vk۵dD7{/�[�1S54W�ET��{N����]ܾO���ԧ+��j�����T����lp�B�z�kܮve��7'�/$Z�\��"����X�.̵��S��/��������H۝�倂��N�4���ǰn|D�R[�^�V��A�gy� �W�i�������O�m��^�PLLQ5(^���d�wY�k�v��#��� �]s���o��z���\�D���'א��V�I!�6~e����u�(���x�S5D�uQD�Kِ���D�o:�b7/�e��I�AG�&I�Η��&#q�Z��Ѩ��q�=z�<s����[4Ϸ��!�MJ*�*+܃��tπ����@��|��ǻ�W��k�'�F���d .��r�ƆDYHP�MC�=λJ��];���c��.�@m�k��#oo��)�mU*�;���;.2З������B30�I��+h> :���� |�ދO�\�g���Wv�����٬�=Oob�e<v��f�E��׹�gh��}qM��%M?jŹ[�}[�gW�I���+�H+��uX�Z�d�����ē��}qi$��O�!87>"���(��/	G�=Q��o��5����ny� 
�{.L$�O��%�F���T��i�$���L��L�MJg{חX|e���eV\��p�\g\ZK�$�nY$����O��ќl$�"�-�ڄ�[��x��ܑ�s׳Dm�v�#Zc�����<&R&fb ���[�$�K1��@ l������Ϲ�gc��Z ��嘯F�
���EI�%���6�W��/!z�߭P ��˻��g/���kOԞ�m��ʾo#<��KI�`Ą�m���Z�w6�K�,��q=�WCMS������j� H���i�V�r�������QZu�Ƕ"p}��^�ӟ���;�� �Z��7��}������8L�~g`�د���9��JR*����{��uܳF #l:�n��Ȭ�n��{Zu����t���*�Ik��x _�#_d�Bsψ�|4�+p��%�z��ٟ���T�`��]{KN����Afl�� ns���T����E*���v���yz���z7Z��+�Aظ�!��ڛ �ۅ"~���y9͙㿿x���ݑ39�g��v�X]�a���"d#�w}cMV��2R���A�UUS30�5�m� ���u�}�ޫ  ���l ���` xtDe��J�̫��d���QRf�M<�d��gza�A�B���s}�>�{)k��%��]�(�I<��lz�[�0bB��6�S|�Y��=b�a(U|��d^�L���z�[�N���D���ޖ�*�5QTW�ET����;� ;sqڳ�������&zܶ�ok��@��we��O��b��[=+.n$ۼظǳ"ܓ���V)޸|z���:��W�t�*t������{�������^V�N~�����o�{���e�ԣ(�G�pW�7<c�q����:MZc��i��N��6C�֛O�莸�7^I���>�����$p�Я��)v�F�V>���y��l����=�`���"Q�&�ݳ*���zH�w�2��Շ$�Av<8�:�����/B���S��=���.���
���|�\]�)�J.ٺ���DC�t*4��+�2�i��M"w]�0hX}7�ՏT��q��O~�9"�{�ҝ��Ө����6�W!Y�l�jhW��n�^\x��㳘��d?ޞ\�X�/m<ר^�=��}b;�蚮o�����f�ӱ��ԙ�ǰ/0�u6���Bه�*Z�I�����������>�۾I���k+u�������̟�w���b^P��n��z��H煮\1�O}V�O�����Y���%$�Rf�u�!�/\}��"��ohx�^|�T�իO�w��k)�Z��ToxOnk�q;=���͋��y�������j��gn�ǒ4r��6����{ib��_����=<,)h<}���;9��:̆��B��*K�[S5LS<k����/S���iR�;꠹#���L~�� �V�;��C��=���+0 ����B!��;N���f�N�0K��Y���m��[��>Ntm�
B+D��b���Q��<�by��������.ݖ�)�C#���¼�AX9L27Q���z׉�����~s � ��X
E�a
���Q-������Qel�i-lE���b	�A�m��Z�W7��J�(Ԭh�5�Ʋ��B�)Z�����V�f#m����iR�V�Z�%c����meQZ�(����"�kQ��ը�#e*�-J��X�,E�R�X��QED�������!���m�*�(�F���-�EX�,qX�.��J�
�Z��ZX�ʥ���KZ�B�TiV�JE--)Qm[DmUq�Z\B�JV+*���)iV�j[Z�%��,j�(������P�cV��V%�EUm��ZT�D�U�R��X��,��A*W�*�QXѱQm+jԴ�`�Z
�����Z+m-R�
���TR�Em�ѶV�\�f)J�)me��Ki
���+50���[j[b���e�b�TDb5��3JdKhX�aZ����c)j����ŭ�bT��Y��a��Z�ъ���AQ�[Vkm���b
����QTA�$EA�(��UR6��m���*(Z���kbV�eE�DPH����������n������N�<��<�������n+ۖq�����hm\<�gn�J<c(��{yoƞ������֎�e�6w��� <OWg��2Iv������/�1�5m9]�%��ֶ{Lp\q�{�z���N|6�v���m���M{c�g�C��t�:n�ܐ�����;���m�5�n��=z��^����@�=s�s3��6�����W;��׎�p�,����;v�Wf˷6��v���I�m�l��kF�F{�{h��НvS���'N뱨�M�����j:9j6s�^'qOF�Õ�K��P֌=���hG]��[�6�V1Þk�&��
��Y�8�k�.�1Qrq���n�/A�NN�L�#�+@��:�J]�\ݤ��Q'#`4q{7r,뎳��i�
�db��������r+&�=z'���X\/8�ǧ��'f�<��=`m���w�k���nۧ�ۢ;\�y�"�#i��;-��u�*�Î�g�F�A���+ۢWB�糱)���)��Y}T̏j��J��2r^���Xc���(����k���xn+p8:�W����o]�ݢ��> c,���;6�]�3q�4g]��#�!��t��n΋<�F��V�b.cQ�״�y\�s��d{H n������v���z��z��7g2 ��pU��n���nխ��H�i=�qۛpf�r�*=�n�3{n��]mie�9xwc�M[�Rsk<���{m���Ua�}�JdN��֝YG�]�m؞ �5um�FƎ���;v/4�����Az����Vԡ�*�[�i���}�݂��x�ާ��.ˎ��Z�ͮ�̾![�z��e�)�Ǆ�:|��v��c������$]s��f8y�1�;��:�"�i������s�ܽ�!���Mu��%�(�r�N�kq��W48Gٸ�è*�[b�Wb��Du��lN�]u�d�&�:"85 �FR�%g���i���mZ������\��<�������d޿2q�v؋��硳�M�T6gq��ғ��]Y'_��A��� G-�]�F<�v19����M��e'� ���۳Sq[=�p[u�\���!�ۜ��՟V2qո�tHÝ��4��B�瓧�{a��5؋H:$��c�a���!�p�Ϸ�-���n;unl)��v����auˎ*w+�Rbڼ�p�:��5n؟<�ׁ<Wr�2�3tvA�;:���\��]U��"��+��}7ݿ���En)��(�޲HU�4I z�d��}�����/���M�p�J�Œr����qn��p����ɐ�ї齝�)Q�6���N ���c��=��rp��8>o�����J�ч77wRCPo���DL��͉�����n���7}�H����I���y����3�d)�T��&�uP�`�=�����I ��v�� ��Η���3��nm�xI�@@[�$Q5����3Z��FD�I�3�;��o�C@��wd l�t�6�����P5�F9�T���!	�$C����b�Ȧt��˱�g�V����El~�~oߝ���DMHmrG�'R |�������m���y����i��ձ� �v�y��09$t�
 ĄM�R�X� ���|���"��ǚ��E��X���?)I��S{G���f���U��~'��b�dH�+�{t>�"?e�,j�n&I��-L�hƋ�� �GW�@���w@�����"!�S�/w�>�O�D�e�s<�XA,'�w6mz��Y|fs�S ��+�s*��wt� ��۵dg/���f�	O�77wRCPl����O�ӣNΜ��O�1��e������f
��=+3�K���f{~�A��"f
�7a.O:Ǧ�D�l:�!f�o����o�o�n� ���� o{�"O��:����>�WI}L�ԅ*��fz��n�9:�n����Xn$*�p��':=��������P�`Ĉ���4���}���[���H����ᇬ͞�o[��d d�8�~20dDJ�J10���S�$�w(��+o)�D���}��0���H�>�7�H��a�\Tn��}��H߁����And��z�'�>����#~J�;�Jɗ��^��]��8�\M��=��Q��D���)��.��jL�V�]��a�s
���C}���h��G[_FW�F�`}.5���_/��Ϲ�� 	9}-�|���`�W�q"�H�Z��n�9M�/�*�M��!���L ���က6�:��R�{����Nx�@}���&\�R�d"W���e7����2���u��l`�_O� +��8��h���?C7����v��������~ҔaX��.0���璲M�fvb�bL���߿wg�m��j�Uo}>i�_fטDD{�$�^�Pk�4�Y�5Ʀ�O���U�IzS�00�0�@!D�Fu�[Đ]\�o��]\]������ ����K��oIݳZ��v�Ec�{l�/�R����&�4{�q��A׹�Ł�T��%�!b�����>���0���z�b�-'�(1$"iZP�l�yqާ�;�ǯ΀ >���Ay8�膣��vTH���ဥ��f�X��j�:!_��1S��$��*gu���W�����_[�nw�M��!f�2�V�򈟜/xU�?�%��$���g��K��O�d�Ĩ�Dԡ6w��v�>�e�t�z\z"�7f�� ��ϣO��&̅9vg�wִ^-��Q��z�.�ֶ��t��,��0���5v�봑2����"g�*������;��0���n/�9}-��]�-��n���- >}�v����!YHQ5UU7�i�Θ��q7���@�+�j��os[��l�����ݑ�?1�sM���X0��=}~�� 4��L@��N(ޘ���=�$�׸�D���E�H�<��fL�D-D�g�?V���w�q*�@��XO���jȀ�r�[@ 7g9��ڈ��p,	%������sm) =�PH-����z�� �w�=��T�s�=�Ɉrݷ� �8��i� �3�/����d���:ܾ�YQ4���ojm���Dc��K��W��B&���wI}�~��[>��:�O&����=�o:<9�Ƕ�]�$����f�\Z`��/h�C��n\�[JsڷiB�9tƹ�8�78�%��\N7:��㭻T�u�^�o]�qq wIu��.w=��\X5��lp�Ƙ�vv�y����ո�u�v�j46bݺݗ��v��w�b�<a�f�K��(+�g��v:vX��n17o9	�[/g�� �����Yd�i���pvN���=����A��Eضm�'N�㪒����8������b��v�m�v��r�cn�Bu�Gn(�;=���{�t)�*hB���ۗvD4���0K�&�z�҉�	ؒS���fD�|��y��YIO�7������§�49��o� ��0��3�,�uC�t��Uy�{r�_�Ь�bd�3d�w�l��rn��a)X���Q��� l��� ݞ�,	O`��`�m_��{���eخ�3�� ��>S @wOk�� m�u�q�N���c����%��Gyn���+�"jA�G��n��:�5��-�l�ȳ��<�BX��(��Hs�w^$z{�9s���rd�,n��Y(�+��Le�\��l$��m��NiA�a�~�{�"P�-rP�n��H���\�@ ��:�"U��jՇYE��KL��;�_�d�u�!
e4!6w��w`�UK��o��5�m?Ud�����,�*�Ė��ܘ��K~3(щ�	:Sb"b�2�Y��*2d�iЦ�W��V<�ᐻb;�
J���� <KT���d����"Kǿ^{^	����w�~a3̙��U*��f*a�ѯب> .�9ڰ@��۽�L�۽�l"/M�K@ ����v)j�!�!bd�vi�)V8�{���Q}�D@����@ d����?��W�J� ��&�d��� � ��S
&j��Ł�i��S�gT��*�=㧽Ys��,w��Y�g��<�?x%@� $ŋPH�h�\Ά�����Əau�a�;^w�c�؉s�������(��aIQ\{��0���n- ����o�
��]6��^9�a{�����&IДJ�DC	6�4�z#���o%�Ћn�Ud��x󛈴�_KL�/ǲ"X���ޙ�8�[7rBMEM�o��v� 2��g�3�-��c�[�+&�:��yB*YFק�T��_?��a��riO�#w�9�7��qxN]����S�tad��<�pr�Grب����:Z����|�]�@ ���n"� ���-�c	��T���d��4����3b3�e�S��I)o2�N{�q��D�v�OD��
��ٻ�E�ڐμ��Z��.i
%T�A^h4�機 ��������֌��{�L��G+ܽ����qD�K��;�X�,�g�Q�G��1�?�]��W�ힸ�]v�t���f�Ǆ�:��������D�H\����0�L�-|��f"RMn;��H��:�	a�S1T��]�ۙ��|�N^ϡN��UML �(�TW�����܋�g2y��cI$��/��n�k��.�#'����]�����Y�$�J%M"#�	6��"7�L0��{��������Ƚ�-M�;�m��HJ$�]��y���UC��y:�Ibז&�$ܞ�,�F^�\����M��T]>g�d�X�uS��n��5�Ρ��&5�j�-�7��L�5'v�'/M�X���ޞ�6ɛ�+]!|�'���E��b�W�!$&��m�x��cN�1�[�rS&q����F��o� ]�~wd�m�C�������l��1�/s���T��2���	F)$�S& 	$��p�v��[��7C�\f��ҥ��Ѱ̿�{���碕MT5�H8}��A��w��@^�]�W�G��3��������l� 9�/y�6����-���d !uR:��n.��ڦ ��-��Y8��;o�;og"���k��QUEL ���t�q|� :�5�� �ᐊ�X��Ny%���7���v�Wb���P��D1�������z�zHQ�2X�<� �3��I5;�o��Y�p���(�d�/������	�o��wdA����t��׷Ue�/k�Y���Z #����{���a���2a�	�y�u�N2a���iO��"j�_X{J�#v[�Dɩ�g�����7���̜{�{V=e�����;X'͋�ƽ}3_�}��������n�����v	(�D2wd:{"�%,�7<uA���Ak1X1���>��v���m������pgd����Sv�Y��m/^
��vwa[q�^_fNHϱ�Au̓s��KkW/�em��r�`ձsyw����vz+[�ru�sѸ�r�3��`z�H�������Gs��)���ۮm���=���s� ��&��d�=���ڠx9�9:]�N�٧2˨:�W-��,q�ۮا<j�Z!#��юk����_�:�\��O�����h�r:d�0bɆVJ�y����3�����'���2�#<| ����,����|+�{Bϥ���VT83	��w�񓌬1��M�����3��Ѧm'�����:g)�>��U�������~��_�/B��0��YY*`��;��d�<pɄ�8d�*_w�u3�,�ed��{��s�}�Ƞ�5�p��I���DLk��q���e�8�'a7��g�x�3a�C0�%��}��6�!�a�a�0�0�O��}Lc�w�fR|8f++%N����<��2VVJ�0���wP�6�Q�^�����j�+��i>p�}�}��V����ƭ<>�>G�G�ނ>�w��ȓ�a�I�a1a�L��wp�8�>}��A���>��-�ע>_<׳l�hf�03	�����x�0��ޗ�72��Wg��3	s�y���d�,�&Y�{�{�|�i�o� gѻ�F�zLxނ#������F��Le�_��u3q��RT����0�a�G�F3��m��f,?H+��]ӝ<���D{I��)��n{Ga��ZL͒���K�\������F�sK�aS��~h9�J!Y++�o�m���Q*���ݜH,��~^��$5i���h�!Z���wPӸ��!�(����A�`#�]��0� ��'�[�w|��YH�n����F��[1&+kS��t��8�|���2��4��=Xb#�H�������&|��:Nl�@<��֯e^c��� ����vf�h~IXV��y��H)&���������}����8Oss��M]����s���l���k�g-q�L�����!m�wߴo��h0*����_[���?=�G9�� �> (�Y`��<�P�62T������a�°�:��8�p����]Ï�E�?���o#��o�!�A�H,��63l�P(����ݜ`r5�Z����{�t����{�z� �HV�\��jv0*Y~��m�9sR��W`a6$�{�tq8�YY+,d�߽���<2��s�q�#
���z�ᤂ�`�ID�����$N2�VT��}���c��s]s��u��ϝq�Wp���Uպ02sm�=q�ָ��)=�at�K���<.1�ne���W��������ii
Z��ߴo�!Z�E �C����a "2.{��LD�hg�/��u3q��RT}��m�#
�����im�˚]�a�;��00�}�Nx���:s�|u�CY���D��߾Ѵ���R
}�P!�PC�����S�z�����i��R����c�L�9�.݁��$�{�8�++%H)�{��N!Q�|>�[��nn����X����i�2�[�����1��\Y�{8=Io_0J~�ѐ&�_x����r���{ݔ2  �*[y�ŗ}�]��.���ت��7^yE��<��;�x�O�nd��!��d�˾/��X��t�=Q|g��YV�<�Ok�+��3zݕݜq�/���N�帕��{nR�����^z����&�"s�m:�lQ.ՋȢM�s��\�'^�Y�a��3��V���6�w�D�l.�BEݙ�˕3&,x���ܲ&a��=kH��gm��{��:q��t)�gu�Kў=�c=xA����yh�ag�������k��+Y�{=G&�3҈��:��8�ҙ�,^%5ޘo&�T�Aw���e�=#�;ʌ9����㶉��×b檪;��\�|E�'����Z})Mn]�����B��8����p)ҍ1Yi<�b6�l��ʱχ��x�E���ח<������Z�S��b�$�O6^�y<�|ƒZ��<U���v��r!�S�za����>(P���ʇ�?V�?��n�����q��F���jǖfя=�c�{���r�4��m�N�ʫ w�� �0��奨<��8�u&;�s��ƁC�~\t�N����Wn7�ڮ��#ݗ���'�|��?>m6����eƴ��N�>��Ť7:h��F�=|V4���@�4�T���={z�t{&�ذQ7���	����ɻ�x�Vf�x<�>�P�R��� h��<Gř�����^�z�c��C�ۮa18מ���9������{����8��Í��(�J�,�q��� �,aYQb(��[* �hҵ}�X���Q��-���"�6�L0ˆ*36�hV �p�1fAaZ�21b��8�ص��*,QQ#D���QDam�J��U�bŭJZ*���e�EX�Pk(���)E��*�#dQKJ�"1�m�W�V�W)��J��5(�"Um��E����g	JQ�j�3�.T�h�ʱ-�0g9S)U�EFe�0���`�im1�adT�p�c�,��J1jc�0-,QR�8�Qc0�D"�Q+p��*,TQEaPF�DAF*E��b�8K�Q���IR���X"#�E���m�Z��PX.��bԔKh�����ȵ(�kU����8��	�L�c�����&..&S8�0Զ�hcŪ��+R�m2�F
VK�B��Ŧ-��6څ�QR��lq�`RT�*��" ���
��R[k�R���HT���,EkRұ�E��X-b�QQF�j�e�m�m�UDU�*V�$ '�}�9��AI�
���߾Ѵ���VJ2��}���q=��*IQ�Dx�[�������s}�Ć-!K@���7�R�
�N��{�6�
�����wP�=��=އ���<�Hf$�X���<��|�Q\�ƃ(��o��$S����O������6Ͳ]{���3L�_w��@�%@����l���
5!B��>���R�+P�y��#��>�5I�"���wJ[0�LD̡�)�{]���ba�W0�Wh %\�4pt���%�ݬ��H��@ē���}���YY*AN���h�q
���
����ᤂ�E�����~w�9��L�߽��N2�Q�����{�tND�>��c��ˌ[rQ������q�AHh���;ߞ�\�7�sF��*Ah��g�{����
�YR��;�i�d�T�S��<��y����хaO~Ϸ�Z[n2�pXn0�����!ĔB�Q����%P(�[\�w�|���<�1ޞ�;��jB���>���R�+P����v0,!O�$υH��%P�W	.�?�N��/~1��}��@� ��T�w�IĂ�XR^���H)&����2V��D�A�S:jJ��Ŗi
���V-�w��Ӊ� �&(�e�G�E-����.y��p�W��Q�w\��9�ݏ��NͲ~eH)�w�������&L�*"`�(�|;��fȂ���s�}�F�R�~��Ƶ�}�w�H)����' �R��/�s������D����$�w���w����o������C�]U���r��l�p/n��p2<�*�on3�W�WXW�������<�q���AL���h:�X�H,�纆�6ʁA*����08�n��z���C�No���� �HV�_|�u;`T}ם[\d�[G]��I�����q��Vj�������<�I��h�𒰣
����>�4�l*J!RQ>��{���T�ɝs^>��0��wC�������T�"
RQѶ����`� �}�ѾR�
сS���a�߻�@�>@�D
�%��P�6�P�J�C�{�tq ���s��Vַͣ�,6�V:�z�bf�d{���#�f���ͲVT
����ݜ`r5 �Hvw΀;���k��(��U�<	��u�GO�DG�qB�!!LL�h�[�F����%H)�>�hg��7\{��8���a�aX[����L7T������d�ed�+%eO��:�0�v`"�*�w�.vws!)�9sd���	�����z�hϓ�W'����s��}�[�k2�2-���FQ[X���\�^&�r��L;O���w��;c~���z^��ݗ�xݑ3�m��n;\�q=�p�3�����u��m<���������֞NAX�s����M\��޻e5��^�Ny��}N��n����&�Nݱ[���]���X��Nm�1��`ތ��y�L��^����4��d��-�g�ע��O+��s�Nݝ�įh���=>ɏn9�c�Z`�Į��v��Gn��v�nɻ^K���8�pm�z�� \�:"�W\�If�������~�����쬇?�ߛ��������� �-�w������
�0*_��}�NO�v������~�hK���CL�%Bĕ�����0�,�>�=W�G)���
%�΀���>�O��mlS�����{���ͲQ��P/<�߶q���
5!KO��}�H)���s�Uz�_��G�D/,�$bD�J.2�	�'{������X�S�s�tr	8�VaXyq���t���3�9ߡ���%�{�tq �q�����s���s����;���a�%�`r5�������[�8�>Hf��;�{��R �`T������� ��	��^|�z�J��8�_R�M!蒡bξ�Gq�ag��9���n3�GpXlaS���8!ĔB�Q���wFٶJco�}��s���{0�Ԩ�߾���`XԂ��Ͻ�R��j�<c������;����鏝��[K˽��:y�8:��xN�����;�H=r�X��n�7�����|玸��ށ�tI�w�4q8 T��S������T��aXR���4�R\�����w}�|�CI=�{�4q���������g: Y d��
������k�y�㴅- �y��}�O��.�qݾ~!R]����W#U=��&��x��{��1�w�U�.~U���Ll{^��Z��х\vk���Oq��~y�4o��+c�`T��~�@m9*T
�'�y�0�6�P�*c[���o����tu����0�DI2Dɯ>|�}��q �VVy繆�62�Q*��{����;��ְ+R��}���� ���w0۱�R�u��k��*��G`a6������0��{���F�ïI&��;���"y�}�A�"��׀u|��^����@�yx�_=��F����"(	H@���0��S믗�|�@�B�n��'b����^�����
�����AN��<�0�ACq%B�=��Gq�a��)׾��Z香�[[���.lۋ��6�v�݇��[��Es>l������������\g6��Xu�O��{���Q
�YX{�;�`ͤ
	P=��Fπ�N*��u��tT�$xHHU�eÔ�i
���s�`T�|yq|��s���[�6��u�h�AH,�u��3������.�ȧ��y��'�*AaO|纆�
M�T�=������Y��>��o��I��;��zH�����a !/rD��%$"��O�;��HP��-�w�o��k���:L;4��Ϣ��37����Q+k���OU�g#�[Rb=l�{����c�3U�i���\�Ə����N�Wo �W��cN~��l�W��
~�e��>�4�P�J�C�?~�Gr0�1�>�ǃ���%�3�P�E>���%�V<���ad}�}X?g^h�ͲVT
����}��|(���� *X��{p����i
؅���P�AM��^umq��Z��� g]�tm=@��� �|��{���#�c�|8|�exS��*%�����8��2�VT����m`#�Tf�̚�{.Ӻ�0[0Z�+c�xS��ݣ		�lx��<͌f�+w����������cX9ߜ�4��i
Z~��o�!Z��,�ϻ���AK�kN6��?s����%�u桦m��RT*�����8+�s�h�h�9�w���N�\t0�}��Ԓ�uN{O���T.3l�2�X��{ߴm �8ԅHv��@�$x嵿*巌	Q\�4���f<����S&q��܎��r$���8�Y�J�2T�ϻ�$�%aXV���1�s��.���~��q�I`�Ib}����2ped����>�g��
�$WZ�
�(&h-z>I�|y��n���go}����) ^?|Ѿ!Z��=�y�6�*T
�%��wP�5���kxz�l���%P+[�vvw�1�"}�f�=3=YI�5�#^P˕	[B��n�;�r���M�i��"�E���x{������
�=���Ă���ػ��qs�8�r�a�aS^��$�
�X?y�tm�d�^�g��]<�٤���]�<�Ă��ԅ-=���� ��s���
g�^�[���춷��Ɋ5�u���L�68��� ��i�G[9�����D�3/;Y((����@��B�� T��2T�Ͼ�G�B�+
0G�����G��|}�����\�{Dϝ�8��VJ2�Xʞ���h��wݮ1�s1�L��l5�����#����p{SG]�`��#���k�<����8�
��ľy��f�*ACSX�q��y�u�k}�tm ����u���1����§��=�H,�e`��;�c6�P*T�����~��=��>�0>�`PjB�y�{��A�+D/�s�����"}�"������l�a��6����������Wp�>�>G�D=מ��IĂ���/�s���laS�D>���y_��
����Y�DAd�ʘϿ}�6��>sVә�08�3m3�L�����A�ii-���h�Axk��w�3�s�Q�R�����8�S�eK�n2T(���@?���t4�Q��Q&�wٛ��WfA�0�v.ZN��וjS{cU2�hњ(��:�;Dm�t<����1zQZ����R�ew���s��[��!eW��r�0b�#q\��2�wC��z�c=]C�"��']�[o���xGUK�/`n�{<�v�
��;i�h�9�v�=� 2ˋn��&ӛc$�jn��nu�gi�{��"��Dm����ݷa�ۣ��s�㷶b۳̃�sώ�7�7m�S���\q�-"�r!��1q�yMۭ���1�%9�@2�sڜ!J�ƞ�pu��{s��]V1pg]�k`Wl�8�:�ƌ�⧚=���s�����gg4�~����c\�7	����?0��>�!ĕ
�A�����F�m������~���aG�}<3/��bm�<����)��j�s����
����q��W�ؓ]����e+3�Ow����{�wG�N$0�-��p���*%O~��h�'Y��������s����� �vN1��c�gk;���H)
Z�{ߴo�HV�+X7�����1�w�@�p@�P+,K���P�6�P�J���{��0�°���s�c%]�H)��~�;�[��\��ׇ1�q�}���� �s߻�q�d���ߴm�ư(ԅO�����[�=P�E���(�>��n!o�H�����F=�}�0� H)<�����N �����]�q�qͽ&x°��Z��aR
J	����8��VJʐS�>�'��n��Ξ����ԦD�*��UQ3� S3Rnz��a��Sd�m�u�kF����/�����#/e`;=4��k����HR�
>��h�)
�`V�
��>��ȁS�o��Z���~~��s���i���
$����|0������$L
d�!9w0�
�������T+&y��a��J�έ�7o���ޘ�����^]w���C~�x���⃋��IN�Fҥ��DGo��LOa�VR�?  ��<ַ���d�*J�~�������Ԃ����t��i����*zeO�4	Q�ׅ�D ��4n24j�#�0�k���N�����;��{��N!RVaXpζk�iq��0�aRPB���w�}������eO|����}�4����P $Bπ⏁��@dI�;�b��~�C��)h��;�|�+Fk�;�{�8�*T
�%�~wP�/��٦��rT������0�aXS���a�j�3����s�t!ĕ
�YX>���d�����������]o�sg�`PjB�O|��t��e!Z!|ߝ�4�SF7��b�P��~�{��ݍ.��h�)Yk��T�.�<��o]�q對ҤX�N���7�|��h!�'A'�o�4q8 VQ����<��@m	*Aao�󻆘m�I�9�}�|�o�������Ad�+%eO|�o���+��� ���Q34��$�>����dx/$<*��ϣms`ϩ��Az��/�{�v
Ag�k��H(n$�}�Z����y���|0�(c~߼�L�qs�8�r�H)�{�4�'̬��63l�e@�R ���z����VZ��
�Mabd՝������g�澰�c�9�N(E{�}��mA|�q��$辇k3��~�#i��2�e*Ү/�����:���!�Ӿ}��Ô�JB����i�����h�dh��G@a6$�{�ta�ϖ����yW� ��'��������8�VaX[���p���%�����d�~�1�/����O�Y,eN�}�pN ^����̸04Ȼ8��X9��m�B��P>����|
A�}Ū�����DKm���%+(%�^{�i ��%B��}��0�a�G�Ff�]"'h���)
�	�����8u��T�m\��M���c ��1�t+v!DJ�߱��^"&J'�G�#��hi:�H,�ϴlf�+*A@����`pkx���\�|Hbӽ��� �HV���CN�.>����S38˛��@���6���2Vs�����W���q<��y�6��+
°�}ןna��IP�,O~��h�Ad�)��᧹�����!�ߨd �vRK�c��٦ư{�~�n;HR��9�����+X��S{�>��]���w�s~��@�D
ʗ�y��ĕ߽��6Ã
��~s�8�,)1`߆>�|����iL�q�):�d��=�7�JʁD������08�jB������1���P�Z��UY3�iNd�=Qf��v�U�3�}���+�}�cU}�Onl7�E����S_q��Y�9M�x�	 ���B�!{�jv��o�����2Z5q��@�s�6���d����|��t���J���H,5w�}�i��%*K�{ߴq����ed����h�j~�v��鯨R�G��^D��9�d(f��e�V�3Lgos��.���M;��+�����ˌ+L��Ԃ�ǚރ�v���������!Z��`T��w��$3����3W?��|�SY��G��R
~��q��a���j�8��嫨,60����t�q%B�}�־��O�E��w�=f�,e@�P)�=��8�R
C�i��i�!^��嚎��L�ӟW����'4څ���.n`q8��>�8�*Ae*y�{�$�AaXV��:��ޜ�����CL>�*AIbs߻��2pR%S�;�4N'.��+x�1���I	�G�_�>��@8�:�g�G�����o=�to���`V�*_<��l'*X�YR����i�{�n~��`>�M�,C�<�ĂÆ7���s�����q�8w0�
������!Ĕ�������F�m�����������P)�7��8��XjB��y߼���R��c�g�տy��ċ��9?��w
��8��RÕ�KD+�D�qx�O��#��u����cō����9�vo�~��	հ�t4�qH��2uL	s5�彃;�W����wOٱT؇�ԗ���}}��$5|YyuL�Ɣs��3}���|���־~�{rqQ���>>A�==�;jyx[�e_Us�����@0�|�5�W{ܢ(����!���W;���ߖ*^�#�ض�k�����4�NLJ�7U%�����o̱���=9[ ���d+Ѵ��4�̘cl��9f�1�*�UZ�
�\%(73����y���yۿ���jjX��S��yEJR��䡻�(��;�r޾���JNK'��y���rP$�𩂳������!�I�5C�N�2��S�p3{�)�ߔ�����Q�iڅ����9���R�f_{�v4��_?_ w\���x���彾B�����n�|�M���=�����x����2���Nq��YQPBwjG����N��07���aCL��!����|�],�Fa��o^���]L�v��u\V�����%lX�2�t���3n�4�͛��R�Pɺ0}���<[b�q�8L�g�Ω�9��i����]��]�:�yk7�Gn�!:C	�_-w~OW���Y�:�U�h-��n� �ʍ��ǌ(y2yU=���v�3W�;�[ZUL=��m�;��냅$���٪�R=���ê�����u,���v�yT�Iv��b��;f� "A/#����eQ�m�R���X#V��+.�P��PY�L!��Q`�p�P�E"�U�1QJ����V"Ԭ�Q �c�آ"��PQf�L�QX���)���5��
�(*�ʔJ�R�Qʕ��"�����F�[�)����j�Z
,r�U�J�`�.[dŤfnU����
�+�mEV�1l(�[Rڬ�B�+XR�)AeDDQKh5+DUr�.���.�D�5l��m*�#-�#j)mDV1UDr�b��
C�+J��0�0���A��V��j��5(�mm��V�V,H�UPT1Z�DU�D���#K��F*f�PV
�`���E���*��0Ţ�E*�X�eJT��-��Ts��*�\b�Y���,�A�QKkm���*T��0
.AUQF(�D2{��W=;�;r;����&٤�B�k�+��R�OW���ޖ85���o;��֎xz{Cے�g����i8g���soc��nd�v���.�͇��6-��B���g]�e�Y_�����VO)��-����*n?n:�3n�0]Ѷ{<���v���R�J��";q'�ݐ��ہ��x�6ηq[/<b�;�$z���B�=�����p���#0]�9���W�q2����c�Ul����p�h��kW��]O/>�:���ݹ�`�kq紏[����`���y����<��-�w�~C����g6&� ����.�ֱuq����A�]��v;�X���O�M91az�W�a��I��Y��&w%8��yGu�F;��筻7z%鱶{:ݺ�ol��wW�8����Q�m�0���r�r�p�Ϩ�^��W�\�Ày]�]#Cl�9<��oQ��y�:�pcnrK��8u����}n;P!؞9���e�5]
TN�;�]Q5�m�|Kggef{��l7�#ez:km�ڻ5�5�;i�:�uɽ�v�Ra�zۇ�kx�>ϗ\OY��tч�3��t�E�6^�d��v7==nsrjg�ɑx-��C�|��3��: "�r� ;�u�����k���a���l�l>�'��O�L)�e�v��1M��l�=��j��\9��0b��uvmI�`����9��jx,靽�u�x��M�|a�=f��������r��T9�9}]�s���rs��s�7<�\%�(P�e�Ɏ�ݹ�iz��p5��v�KRc�r�F�a7n��G�7]��k�3Ȥ�9#ƴcs�xl���9��Yz��֭��чc8:�M��������q�g;5n9L���݁�˱�z�}\L�.I�sƧH�g[a*5����u>�\.�M��f��Y]�8�w��:z������9y�3�7b�d�>Y�=+N��6Z�L���/Y�����d���m�L���/��MS#�h�\�?� �Q֦&.6��q�g�s'W'W[+�^n�����nt�Ӣ�u�l�t�\׆a�b�[-4�աܘM�${OZ1����c���C��֤[f��h�v^��	;�f���;�%�m����y���'��vOY�tG.nWZ�m�OZs��bw����;��3�f���7Lێ;X��ʻ����}5�����P��s�᧮��;�v��n�uX��m��fS��s�-�3.r�;�n���\�d-ջ%j.�������1�)W�'�_s�tq9+(�YA��|��4r$�AaXV/�ﻆ�m�I�5���qw��=Mo}�G82���y�|�8�@���m��8�V�g�ϛ�n�
B��y|����9�o�H/���)��́���R��K�m��D����fޗE�[��Gz0�)�s���q�WpXm�N�\�A�$�VJ��۾��l�%e@�PG�Z\E�gכ���8�<	$>߻��� �B�y���C.�.{�j��fD��F=��:G���q��,����J����@mD��aXP����)&�*K���q�>p޷ߓɖO�VJʞy���q8�����b"QFlQ�Q��}��+��W�w��/��*����3�{�����^��S�|�N ��~߾�H(m%@��������~��������ܙ���@�sN�g����Squ��t9Nv��n�g�������_���g�va�5�{Ib�����6ͤ
�߻��6��Xw���u��;���y�=�H<��h!{���i�����z4��D�W�,�W���0�G�>���f���}�E�*�
n>���j�&g*�:����h���}}ɯ,���'�>�cQq|i�}~�窻y��kY��~�gٟa�O����?D�Bĕ��+/����%B�{�}�l�ed������1���z�n�h{|F�6m�#�V�g�`��sP�Cr�����h�)
�`T����������7���>O��+���CI��PC��ߴq���s�3���&3)~�_��#�t��m���0��*A`�߻�`ͲPe@����{��$�,-=����/1���>co�`�_R�/������Ly��G39ɛ��ND��{���
����>�#w�t3�{v���A�aX[�9��%�T���h�'VJ�=����pN o}�t_�:�O�q�e�W�\
��0��{qn�b�l�!ΈJ����,�H]B�Y�t_?�>�뗳�9+��H,u��ii
����o�R�
�J{���`q ��u󯵝]`���:����3c%B����P���{b�bDD���a��M{�}�pC��������}��;�KP*T
{�~�g�H)�w��R�+�Z=��-����Y�xQ�����BH"\dvq&��;���
�����|��tpI�*J°�;�w{��i��{�w������ti\v& y9,G�Z/���)��5#������� V�ky{Ѿ�6�Ϭ����7!�[�Đ߾s���
�P<���h�'Y+*AO|���h��u���Q�$c��Q�2�(�݈K�w}R-!m~s�Ѿ�H),���݁��@�D
�%�~wP������:�l�Ʒ�C ��b���GpaX^��ysqͣ�,60��k��8!ĔB��󺆙9�[�3>cXR�����Ĩc~w͜`q����y�}�H<��lB��;�i $��d_օ���2e@
L(��/��v����ۺ����z� �z�p�S�����q1��8/@�;w���'
��YY*y�{�D�H,)V��;�i��T�����]�>у��'��w�h�'Y(2�Xʟ}���N \��ט�b�����065�����5����Vu- d_�B��%� ��$/��`q8 T��/�󺆙���bJ���p:ǽ������ޏq�af7����%q���p�0����tC�* �~���ͲVT
��^�w�w�����+Rӽ��t9H6��/�󺆝�h��~�Ȉ��UO�g�Ɩ��S����d�]�'���y۹�.zn訌���J�;x�{V���{S',��A�k����C�\N�D��7�H����r��	�^9&�n(�t�s�=����w�����F>��$� ��!�ТI�ߝY�y'&�LM�5����I��4AǼ�����m�|��Y��#4�[��F%�6�5ʝWC��r�OITj1��l�B��g�����Lz�������lX��@�Fv�1C4LsCFI��#��O�X��-V�ϝo N	*Og%�w�O�@ ��c�^$gsw~$�\,Q���i��ו�VQ7B�J"�fh���M�� �����)A��wd����>9��Y!T�9��(Ĉ��(ݙ}�˻��������M�B��o�%�Nbt[ޑG�4�""A�3$��}�`��ͼ�먍Җ����彚'ć���>!�yv�*tc�w[W8��aq�sjb�#GQ^��}C�g-KcQQq�_Z�/�W�e��.��VB	���gfP:ʻ�WJ�^U��'?|��#!~w��۷e�ۃ�E������K��uc�:̛�\�7��mk��=n�-n'i�(N��������6��J�tt�d�ͭ=��L^kF8�#On��k�I��n�n�����Q�w&�1X�-�G�:G�=��O=v�WMY�u��n^ۋ���݇�����pe7^r�����뱶�ۛ��N����<{v��`���1��9Ͷݹۯ]V��Ki��/HQ��OZW��˹���:��I�y�=�zXa�~�����|/n:�_�DV]z�������[�gB1,=��1��7�ƺ�'ķ�ݒ9��S��&d�E z.��[Z�s��/E�o��߉�>�wb���lU�/7�<J�&}
JRU���ܱ`�|��_�&��K�D��S�5��mP$�۱r' ֌)��n����<p��ʅ��E�yVA%�wvA;���9�|�b�V@��_X���TLbDD��kL�vز	�3k�*�{��ھ����n�@$�n�� ���C�rn�s�����w�%��6M�y��7r�Λ{ht���3���(��"�+��α~$�����|H;��@��,�!�׺�]� �����p�c�<�H&��E;�D�i=S����A�F���ζs�d��	�(��f�-n�Իk�L+�ۤ�{�Q��C����M:WB�)�ޓ��ǝ�K�Ǜ�E#��x	�Yu�'ă��	;���$n���AANG]M����z����\]e�>>�Ϊ$��qJ�v��0	Q���P�,��QּHТ~����Zy��e|u�3��4����,$��H'�s��QSQ۝ʨ����˲��n$��D��m�I�7���T6�;��c��$�c��ۜ�Ȝ����s?��	��3�d%*L"!�/X�=�L�j�}i��+���6��9_�~~�8�!D��_�_7b�'�<͡D��;�ļ�g��I��b2��_�/3f�I��)��D"�*�Sλ�%>qXǲԅsQ��,�I���4I#�9ݒ͔�ëK��^	F:#� ��k�v�Q�>7�άAysGi�9۴E��`WF3=;>����9}2�; �@�υ�ƴ���A1"�b'�ʈٴ��M	�b��I2�o7P!6�����*�������t*��y��S�q��6b��r��*�,�(�|s1S����	#����I�z��I%��f������׳����o ]�Иp,D�GBo1�����}�b���3�^Dm�x�ۻ�d���f{'���9Ş�W*�J�(��T�"��A�����v�nA�MXs�s�j:���=�ؗ��Ͻ�2B�J"�fx�n�(^v�O��ݻ�&��*Vh#:h	o�����X�D�F$(Re�/�ݓ�b0on�=E�N��V>-��*WWVLF�=;�|vq��L�"d��+A�7�V	�j#m@�;�,��Nx�����}�b�8R1��bRDՀDS�o�du�}�T��{{v�I�Ε��Gxw�DW��O:ƫ=���k�3B��r3tˬ�I�V=���l�Wf�%�,��Ѫ��Ɂqhua�W���v��|���f<��#�F(^��&$ Ex�[`X$ng�!uGwk=�&UFt����� ��v��73��ah�54��|�xn�;~Xu�@�BY�Z`�L�ԏ\�mx޼h�a�%�V��6��~m��8�"��&3���vHc����|F�t�.!{مb:�D�U݂=��bϥU�sP���U|Uzg��/G�9Nb�er���z�w� /ֶ�,�o��ț�����r��2b�=���$(Re���vI!�mQ#��A�ɁV*q���I9��v���㓥��f`�3$��쨎��{ZG)� ��U�� �<^f�A8�z��2j�X$�c������0JF숧u����U�؄�:ܞps+F�^S>y�49۽w�)>ԧ����x�6F��w�$�?l�^�5o]c&�Yn=c�;uP&t�n�G�x��B6��;��7ز8x=��ul�B����3����$��P����Ĥu���:��k��Wnz��Fc6�7L&׮4��EV�
��B�c���$;k�'%���������Ȁ������1��E�<�ϱ��N7]����:��nyr�ס"���wm6ل�ޕ�F��ή��ms�*�Qs״�׵�0m�R�5��m����Λ]0����$Hx��;x�sv��9��n6�ժ#�m�;u���<K�m������6kcZ�jecMͲ¢���(!y	���u��H#���n�߁и��1�&�вK��
��` �f!I���Y�~$L�鞚���mm�},����`�w��غx���1��>�:-D��
�|�h����7ݮ�`����
٪=
f��3�]��~�b�3�-A�BӤX�ݸ�eL]-���W� c�wd�絜q��Im�����6E�3(�%T��$�ͽ�k]��������$�N�I��w`O�|���M��W�5����jXJ+�	�ѷy�5ύ6f��u����ݱ�:6���0<V˷$LNwE�@�&`�Gx"�����I!�{aJu3
C��d�E�ޱ{� �Ay	�G��n�1ε��o��)&��/3�}m���y����0[Y-)jF�)�Jw�X�s��B�IF�O%j��/g-s�<s�s|kكT��
���	'~{�߉!��ذs���v��=`~. �L5&!I��畎������Ւt���U���$/w��>��=�fT�J�*	�7k����n�w�ht^��3;LH/��X ���4
���3�k�}�}�`�5�Т`���F��w;�|C�ڮN��UtfR���A�z�݂I�}�!�E�����'ĐV���Ոbҏ=��-Cn�T��p��ͷ^0A�\��p�]s�����:aL�3$�ݼ�$y��~ �s3��i����&�tK۰H#{�س�����&d��N恞��v�7q�`	'ϵ�ߏ�3����5�-m:��wY���
>BbBQq7�d����N f�8�Ѻg6B�����@�	{���x�)�]��+	��{D����9�3&�
;�Ǹs[�TWsfh��[K�%�9��Y��^&vk�]'�"����t/Ht��XŇ�2��E�I�~�-�{��p�۝��a�#���~:8�քR�W�������5�z�	�l�Ç�7K�F/{]ѯ_�p�H�.�"���C�4p��kk����<����j���Ï�pt�ח]���� aTy~<��9����q<��� w|o���x���~%��ч�f�H�R�ܱ"
zC�0�w�9��q��V:��-���Fp�ܩ�I@��{p~�������歆g���O{C=���=DrEWE�ֵ�=2'��jve������*�<ͽ��䝸iB�Vv;��m��~}[��LbC|��,f�G���i�"�x�c�D�nh�<	Ӿ��K>��l��ԮVOz��p!p�^&:,�S<1y*O���v�9�� ��wo��c����-jŀ���]�bvm�嵚a�����y����j�Bsa�.5�
iZtFz�Uey�-���27��S�$'�܄N�y1AL�����f��\=��q�F,9Q-ƙ�7�V��&bt9e��)\�|[��a�~8���ӯ�B;랈��of���#L�`ǲ�JU#[WX�v�y[��%���"�:B��J������$�;<�ъ��|K�#k������z�o�@=�I�ܽ('��ikE�J~��&���yZ�>��L�����";�0�ͨf�ËAY"��b�*1b�V��R��T���A$��EV"
�1����(�T0�TQ�R�Y�UUX���(�4���KDf-���V,��$Rb�"ł1TQ��E��*�f�PD�h���"ZUs�0��("1�*�"�E��UQ��ZTshȊ
� ��(*��Ub�DUE�Z�R��║H���c��b�b�Lڊ�AED��,���+`�Q�b�F*�TE��Q�TT�F"+���IX**"��#�b��VT\!TQp�A�E��m*""��T��Db��FDE�ZȨ���W	b)� ����V�V"�^����>�Y�|��6
��� ��<S@�H�M�δ]�9�2�`΍a�]�$��� �k����N��:��{}��%s�UAS�������	�y��}j�7p����A �gMN�7VxI�Բ��^ޣ\)S"��n��,�M��8��5�n�X\�8lv۷{��d��fv����(��hCok�<͡D�N�n�{�YPw��%ٶ��\mu��vc��>9��30x̒�O_u� �wRJ�j��t��|C�٠	����H ���Ɨ��}��Rs"̃!@�)u8O�y�՟N�-�8���][��@'�s� �}����\��BH��BW�F�W㣣�Pr���`$�n�P$��[�>n��-,v�WP��3v:��+��|�w�wL��M�s���K�i���F��ʹ�&��r=]]8i����
�!�N5����;��N���P#R:y�?�l`���d�r�QKwAkf�H$���$�|�
���:v�@�)	$��"`JR�Jݹ^��^^���.h9z�i�qu���z/��߿A��
�L�,�:I���d�����]� �n�w`�)��L1>Q1(؇}�Y��U���T�/q�$�����H-�; �lT����/"�8�82bfd�%P���`�H��~��NVe���	��I!�7b�n�س���S��12%"�4�)Y�������U�	#]�v	'س:.����铳��`�'B"�D��z7.�x��Ω��[l��ǅ{k+lY �����:(��;v7�w��lڹO�7�OipD���%��� \:��;9������y��N,�HN?bY�^�R�4U��+��Z�_��~)���f?��������E��q���69���i��3�r���M��+��g�A��N��lҨ.jdv�mRu�-�k��;
���G^1!��I]Ոϳ��s��`�.�r8P�����qɮ=�sُ%��ڵ㬇<*��qn���.t�f��y��fL�<OTg���tU]�]m�4v���	��`ݸۯV�V��.��{[k	���/����]���뭡ѭ]ś�!D3��xG���SLo��{v	��_;��3��Η�­V�Kt#m��$�mسD�(��	�v{d���l�};�Z$�����3��<�C��/�5��)�'�&%�=��dg3jA9�W�0!�$g-�1s5�8����O�ftP#'�&&fA��UOvu�zs4ͩo��$����>'���آ��� Α0H5���Ϧn�-Ӻ�'q�w�~� ����=s�|L�Vݒ	f8�A�}�DV��VE����ࠊ%ET= �;m��ù�#���QfN�iz�������tLU��L�D8�~�	:s:�o�;��r�ղxM��f��߬U���
`�Qu	׿N���#�'�}#��a���}�v{�w0��c���[��x����cr/U�W�V��@�e��3�r��RSf�Щ���)d�������Jp��mu�7y�Jo7�`�ĵ���7��ݓ㻑���t^���f+f�BQR ��L�;=���� �i�P���W`�9�	7ϝ_�SOf
�0b|�bQ�2�p�ɚ8R�$3�RA>'���$n��[�B���(�r˃&&fA��Uz_g]��O;n�إ���v�/K]�x�����In��tc���/y�0�)\Ҵt����V�i{�'7s��\�0��<��b�?�;���ʹ�$H>�ԒA��u`I!��v[}�9��'	az��E����;�$�F	����z7.���X0^zq�4	9�ĒN=�V	$����
����tq��L7+h
#��:���@��uhsīn�D��w|����|���U�'���Ըv�O�w�-��,��@~���}���}!3_=cv������92�J�o�=s{�� �s�$|[���V�"���D(S虯;]��:6�Q>�oU��	���I>řйѨ=u���8��U��X�v�0`̐�bQ� ���Ig3j{�*�M��w_͌]����>\�_�>�Ͻ�v�<�7�Z�<�����e�npkiS���=f���{���s�Aε?�~o��5�x̒�6�q�-߬�|Hՙ�@�e���Pݮ�q]�`�H-�;���XLȉ��eDH�0e�	�'Y"������$�<��A��Ί�R�1��t���}�� 4 �� )'?�(��� ����9z3i���I ��׃ �O�`��	�`(�:��ݓ�����ɵ������H'c�$��;���xb'��Lf�m��o'�n{Ȏʛ�Z���p���esrn�ʨ�s2�#�C΋�甆Fy8=f��G�b��㹨��W��|�~��|�|{�� P�>�� ���z���~(]f\�S}�Ov��$�b��A9����9��#p���M��G��J��D�mk��ǚ-�'��ы�'W6Q����Ͽѕ�).����g;� s6��	�>��,�v`���Q��N�'ڳP$��pd���3�2J�}���Κ�jEVS[\�,_��ftQ ���~$�Nf"u�3[DU갮��ըi(�<!^��?��~���<�c�� 9�	�6���ޙ'B0L�0�A$��3�re	��T�I���H$�\�L��if.��)���Q%Df���f_]�I�\��]���@�`�j/���7��u�����{\:'r��$ެw�]H%����j���0��^ݙ<�^&OPk*J5$3��e{n�[�-ѻ476�s{t�N��Nh��{�,�%�A�"G[#�F�g\읳a�mX:���g�kJ�a�ԩ��!�n��e#q�S�In��r���OZ��⹝���7����sv����rh��CZ�F)�=�ۇ�`9sB��ђE�S��+�g����$r�yx�e�'�������u\r]��+v�x�$��g��$A����]�8 n�C�ި7n6�������x|����8U�^ݱخ�3�����6�=V�<<aLE�܊����O�c�ǩВ	6�_�$��s�2$`02��-�Y���@�H���e�좢!I��)`�����A;���U��O���|Cu΅�%�V�f�{V�i>.p�31&D�L��y�݂I<黲EA͋G�mܐyA���ۚ��7\�]�,�dD����H�0e�KO`*;��:����7�V	 ���vA�:&_XA�]�$��b�P@h(�� <���`�&uH�2�)>��w��u�v	>�:+�y�{�X�*�UޑT�
`��-���]GM��s���sE�W1�g�3���>o��*!!0d�m�mq>$u�b� �Y����N�1�	�qB�z�� '�|��Ria"!�D�x�����C=�}_n��1��{z�>�^#n��l!�ˍ��[�c��tEcv� �d/�S�(��������֔�-߳��<��In���>$Y�Ex�sҠ^l���Ү��D�^�12Q30�]��}b��͊� ��rP9TЎpT�;n�#�o]��VgE�yA��*eH�)�UO>�'����	56��gē�3������*o�R�C	'��l]�XLȉ�DJ�"����^/3z�i��ljx�!^��w`��Y��A>���;b����������6kI�+PgN�v�֤�*Й��mƪz(Tf4���g
B�{|�=�;D�I�F�U��1ВA����s�Q����X�$�]��>'�c�$���0Pa	FLݼ��Ү��Ư2���'�łN�Ί ��U�wU���7~�Ӻc���!7!o嫅�٣	��ud�i�3�Q�U��A���V}�|��z&}:!�ӣ��槴XP5Ϣcn:�щ \+`D�2���b�x牾~���Br2�vj�Y�}���x��gEx�F�}�d˛�F""$JFf��-�,]�5���|H,�mI�q�v/�����e�-X�r
1��;�82eL��2J��I'ǞӱsX�ܹѨ�	��$��;���u�J�i����6$"�F�$�Q�3;k6:z���f��u�;�lO=q��f�M�����}j�$J�#x2�>���H�-���ں�GvI�=�H���~$oD��J�bA$��3,Y�Uﺡ�I7�b��I<�z�Ē[����T딫:�����0�w&j���h����o�$�u�W�A�WP%�w=*�+Ē�}b�-�;���EDȈF'�1GuWz�&Z�3��|	��ʲ	#���� �������?kz&��b��K�G����~�����j��`���.��֚M� �}�</�9җ:��h��ƭvʬ�;sO~�>9n�ā=WҌDDH��LD���;>$���'�B�pd��TŗՎ��F�s�,Hՙ�)��?/�N�� ����.�N{zz9fR��s��Z�q����:��Ԙ�y��������E^+c��ۿ	��v@'�NgEx�
c0���+�6�Ēu�bȾ僦fBQ �Pd]�2���\�oOtu9�wՠI�y� �d�v 7~Cl
��lO�� �J�bA$�.+r��wuz#�쬜�'D4�f|Io�ذA>�����x`�!D�Bn��g\�Ux�4/��l$��fFr	���j��s��A2.�l��x�q"�Z���܆����0���B��F}{A�Ͷ���B�O��޻87�C�Ľ3x)S�zcZ��'ɺmeL͑U..��ơI���w l^<�Ӻ�����Ͷ�i:\P����8�����3�1��c���b=�Rg{���Yw�w�����3�l>ԉ�~�'�t^�1��a�l{�g\�n�>S����/���whS4{��`����I��Ws"I�i�Y�,-R�����NBt`�!�,%"S���H��7���j@e��D�R:�nw���x����~��a#�w�Ƃ����w��`C'6fl���*�ٷ�w��'�'o���J6��DIl'uB�5�8���敺��iR��/}����P�ξRm�����t�2o`�%�N�9�M�:^��n�J�<�����Lvn�&T�T�������7j��=���Ӭ�|}��	����/N���R<��	�X�����B*^��,���|$��jm�B�K�s
Ÿ,�8�[�5�*i��x�!��J�i�ȇ4�����|�����=�O�]؋�>ٖ�P�[���\�$9��8"�y��l�id{V�R��. v����tU嬙:d��x7ئYB�U�9�Hp�`��/*3��7sO{��Qp�^��}���7���6��<Жl�`�cwNe
����^��H3E-��5ʨ7�G��g��^M'�~�����+1�cR"�ߍͷ��k������]sj�;�z�=���pY�k�����rF����sY#���l�=)}�R<�����bg@r83H���:��q��������Wz7�G��z�������"*��QUb�*"*[
��b"�Y�Q�*�Q�
��LZ�X֋"�1��c�����8JEX�*+F+U���1p��(�����	���\%AAm��H�ʌ`*�`�U�U+Ab#"�E`�"�qJ8`)E��TQ�X�qj��EELXQD"�UDH���EV+QDPQEkb��n."��1kmUUAb)mDQDQ��X�"�#m�"��1AE�(�`�EEf"²��ȬUb��b���X�[(�E��"1�֣+QPc�QY�Db�c���A�TEX*�(��-**�������VDQE0ŕb�G�v����~^v�mC�b��yd���/I�zةg�m��H�t�jm���ゖ�zT�9;�b���k�l�%pO9 g�]��r���ݺ���[�v���ښ�-[��q��.��%{�"�[Gn:3����T�m��+���ߛ����#�Ca#��n����y����f��;q�5���1/\.�{Dnj�۰��H��cє�rfE�f\rK�����x8Y�7 7md��.ц������+'4��pp>9�:|��uڭW:_n�FK��]���g�`N2�bs�������$�=��x�E�c�=c����^w��S�����z��8�oY7�-b����ݶ�v�V���F!�m��gc����Nxܽ�ly5�[،;l+�nv8�'a�\?��o�H�Ѯ�d�N��ô*��C0��ΐ;a�s6�IF�8/Ê7�����*�ܼ`{'l���#�F�@�cg�r5������O�����:�y|��n�On�<pf�F'��3*d]ї�s=�a��ۅ������:���&��G���q���ٛu�x�6��N'G\���s�:fnfC�N@�l�Z}��۝n��۷f�қq���[�c��{`d;X;��n5��}b��`3�M��D�ug��L5��,�\��Z�c���㜓�n,�y��퓨���&[`�d�!LvQ����>+��/8���������xǞ���u9,8����&���e�]���y�3�;7F������qn=���LY���5�X�5�l��p��h���oC+�⺭�/4/=m���L�ݎ�r'��v�p[��1�ϰ�2f�FE��
���Ð�#�vȣe�����:`�	޷/.�a�m�c�u�^W��������+��ѳ=f��[tr��!onX]���l�iͩR�:|���s!��{a�s���z��N:�8�Y-�6з`��r���ݜ'�X/=�����;Fu=��5#��Ok�BV��n�\f���a&�J���w���jۜ���u�ȷ�S ���㮭�I�v�&�k���յ�v|�U������a�T<]���>m���]���15r�/-r�FS�F���Vv:�29x�JI�룱��lk5�'��Vz��7�Kd7�ӫu��;m�q��c�tq]N�8A��ّ��9�q�v���tI��Ƀv����;��O���t9Su��m�PPS�M����H�8���]<�����Tݻp�݄�FBRf9�����H�P�"E�޿$��f����!����P��S��~/#5Q �PpdʙR'�d�ݕ��g���P˩�ڊoE�>̌�@��P�	��̜9N�_*��>�j����AP�l->���-���3��>�T?I{J�t��� ���	�yؽ表�PPH$�=����6��2|I�N������`7׵��wq���FFڠO�Yc�!�%Jv;)���>�~��;�C���;U I��u`��wguΜ\J#ş�N�0�"t,D��l�d��r��땼��2���o%����_��>�:��O����>$�sud�A�;�h��<�bF�9��@s���Ju{(�
$I�*bEߍ>޿Y ���jqmP��R�0J=�N�TZ�YP�i��eXx>��<�����q�����"<�9\n)�ѱP\��3�/N��ک��W�W1���w:�I>-��ŁJb�b�x;���M�O����Q*D�D���ݝv	���g�����g^�IN��K&	;��X ��پ놦fQ �Pd]��eF�ML�&B��VH$=ϱذ	̌�1�5�#��Z��"��.��T5$ J
��G�^X�'qg%�3;/+h�����H<޻���	����'W�����/#��Vʎ��\:=L�y�6���;ջk6ր	�dm��
f;�I�2B �R��t�۰H#;�ݒG�23��o.�k%֎��+��%����U�I#I*
��wUu$l��gr�3)��|	����dg!^:-��4:�Q�5d��r���D���$]��ޡ`�Y�P2�Wwn.�6�'����w>�C���}<O����������5|�JQ���G��O�:���O���V����ujgv�dl�6~��o��_�k�d�23�(��hɕ�O�I*��u��jpʽΪw�Y>�:��H'23� H�"��*��ޚ"'1�'3v����NbR	L�& H��;Y�|ww�YΈ�Q=�޽�;�<���,j�H&�݃��e,�d�u��qa����{m����f�r-so�$@qp�붇��v�~~���s��ٻm����ʿ��T&�ՙ�V(���"��j�����Yʁ!V2pL��2N��S�u�`����ƫr>s�<d�Fdg*/;��'�A���1�ݥog��v}]uP����L��(����m�u`�]������ �O��f��/;���b"�f
��B_c���%킜�{xO�Z��F7��`���트�j7}|�,3b�	�˝�OD<��&�a����hFm�ܑtK�O>��S�2��왝���.�0�T����@�##1
��4`ʃ2'�J������o]��D6H4K���ۇ�Q#��w�I ����"�]N���~��<#n��jc�^R�;�Z�e0��㕈�xqUH�� }�l�@��B��KQ#|����B�$�w~:\Bm�y}�v�GRHǭ݃��D@�	�H�9C��?���"�� �hޫ ����0���Y}[��S묎��Е�M��BJ�Ogݐ|q����t[͑f\n���ud���]��U	B*IPT�
b��U��@���A�}V	��ݒO�#9Z�5.ȶ9���y)A�$�1"��ޱd��fסX�S$J���Ao�݂Ndg*�ܬfr5��j6�a3�<�H\�mFkhm�雖{�2�Q�M��*�
��-qJ�TlE�+�Չ��7��	��R�C�^�����+�"�(��Dn��r��=�S[f�3��N���۞��X|���y���\uz�m���y7n�n�g	���*�Y�۬â�f�q�9��c���덜�K�EMr��}�r{B�����	�c�nz�3�nӰ�N9컷p��c�]���T�;��qŠ�ic��i8��B��p>�C�}����	x�ڽ��t��'�;��]AF��F�og���tZ�J��Nk]D[��{���朎�+�����h2�̉�D���y�/Ė޻��|Ndg*9���bWs�r�X�k�}\��0��D@�vbS�2#���¥ˇf��Wx�=�]��9Q>,(>����Č�u&PP&L$M�yb�'�qgW����p�Q�����z���̌�D�g�$�Ġ����m���ƥpf��D;�I�ud����T	$^w;6,��L��IO��4�����
 =S�m�u`�E�4yޱt�����H$<�j�$޾w~3�&b��u�ǿ��߼ex�v:����`��.:{hu��i��ʱ:ڍF\:_������y��w������_ O�śB�@�|�@���G	��#_P�C��TH��P���A�����t�*$k[�T�.x�Qrtc}5�3�K�ҨS*�M���Ǎ���+�c)����I}�z�x&ي��WяN�ރ�9g	F����m��o�?���y��Y �F|�	��~� �}=��+6��yG=e_j�[�Cs�Z};����<  <���~A0�_w`#�f��$�׽v�u&P�2&
&�zefd=�5u}:�b�;]�s��Ao9�o��6*���}����BfP3n��w`�1�;��:]�ؓ�W)j� �y��Ao9��ep|���H� I���0���:����c�sNo-�ƣ�Uð>��_������	@�2B����I��u`�-�;潃:�)��GfwU�%��
 ȓ2�ċ���'#y�@odv*�A�1��	-�;�@,s0y=XVtV+��P����2��<�n� ���X<�ځ:�1T�$7#�����"��i]�6/�X=>����=c��u�����K�%�伽J~O\w�r5�o5�	.�Pn��I-�;�&�8��HBf%<�TC:� ��{*�'��$�Y˰��>Q�q��o<��v
BN$75`��N�^,ꆲ�+��	;�����g*9U�f�"��d��T�(���#���f�kc����y��R�Fܹm�7g�3�󹤢AL�`Npson� �}��`��<��@��2u�Y�Sӎ��H9���f��(���S$(��Oh�‬i+s���I��������|^,2	/�o(@��o��d�w����FN�:������ zy�7�����MtZƂ|��v���@khpP��2#�%�W}�B1�AS/�X �;&��(w}��B�4���
��
N�sݨ���.k����(f������ZR�Okp]�9��-�m`z5]��]���e��sw�{��{�v|"�l5"S �PdXP��n�:��c��0��@O�ݓ�Gdg!@���9�HV�T�4�?�����Zt�HR�m����Њюy����N&�&��G�ߟ��	������D�]�{u�y��_7��609O��܌j�5��D���������Y�58, �[���� ��3�A>���`��L�s��������MA12���L�F��<������N޳$�޽���$fF5@�y��ɗ��TDD�&e)�f�o���jHZ��w3����kg�r�V��V�V�d�����D�*�D�}ZI�]ت��RaNE���A9���$����^Sbq��!d�^���.����.�q�w��Ä!�ۊ܈�w[��N�9u>�4�j�d�U�.������"�$�.�Z��G�?��lN������mķd[�O!ub�e&ۮ�<vd��8��ڵq�:��"�m���y:����N�I��e��OM%����;�w7^��W)��6�N5䒤�'&[׵ٝ��:�^x�̻+����Zɻp�E�sm�n9��-Y�ֹ;F���&�����Y-�^��l�E�4�����6r�'&���'F֜�q��V+��	��:OМ�;GG[T�;Q��Y���;\pq��
�;���~g�rb�r:�ߺ��� ���B�|�ߎI�$L�ү%�r�O��]��TNʈ*D�D�].���\��nM�v�r	�/z�N�n�`��4����I�虭��\L�������3�	����d���$L���T���+zР[��d�A��ػ��IL�A�2B��j�X.�(�;���}W�I$�n�i��TW[��Qk����pA>��wd���"%3)LH������ͨ�n��0�8��i>�H� 	�������%�{��ߟ��ճ�΅����zyj3E���d�+��)���r��EL�R����D���D��n�I�mݟi��@�9�9�(���ݓ�N�7V"��tH���!(2,D'k9���X���g�
I{!Ա�'/��%Ľ����
`R��j�v/���Sx�3f�s;3���m��ٛ:M����6+���K|݋񦳕�d�z����������v,�A����evC�H=�V&�rg���|{�v,	�ʼH�6�DHB`L�n�nvخo�#�����˛�Eb�TH'2���ENNU^}��g�[T��A�.�i��G~�	#�W>t�����wd�G\cTO����!��/��������2�V�&�đ��6�v��<u���,��9xu[����Z~|���Ыԥ1"�Ǳ�U�K��PH fgu��y��t�9}���mg!V�Oy@&bJ�E9wդ�gD��J�ki����ՙ��d��I�t�sܼ̳�C���%EىOss�"<c�S*︥�ad/�t��^.�+��o6ye~�sע���i���r�@�4�8��p8����d$Z�>�g��=����m�=��Z�\�V3'��Ճ=)����&�{/�u�lN�ܛ�P/�{B,��Ƣ��[����]�p�m�U� 'a���J�y�A����k����E��#~x;�� AȊ�0^{/��4�����/�*��{q夛s��O�5�wS�:>�j�E�- �-���&�Ǆ�!����%��d���&7��7x'�ۛ�Y�}����o�y����_B�󩫾vf��ݦ��y'h����*.e�$-s�k!�b�ڲ2��4(�ڷ<��:��;|���vr�}�y�+��Lb<,�4eo#	Y¥�;x���P�@B�x�֧��<��P�b~�P �si����u���k�����Ƴt�>V˶%.�*����B(�9���}f��������2�����<ҟ�����W�A�N_r������9��2:��'P�rK��׾���в�!o�Eh��r�{��!��{ș����Wk�gyzĩ�]nִ��֦���s��A�1n{g�7�Q��X$[ZKL��jx����3���<��}3$c٬sw��sV��W�+�tU�4����I�� �Ǜ�`��{U���<V^s�P��c�������)���cVz
}{�5>��b����Vx��
2����3N]\H �G� I�����EU#*>2�UcKj�D`�@EEb"���Tm��QE��EV
��Q
���R�EX��EqJ1bek`��Q�1Ac�S��" �P������(�*�b��,Š"�UR"�Pyh*(�PU�9���Ȉ1��E`���E��"�mG.1�Q��rʕ���ؠ�(��DJʊ�1U2Ԉ�""�[�DE�1Ab�AUAe�m���b�*�PX��C�Yb*�ͅQ�jEDŕG���1@QH�������X�Z�)m"�"��1���@Qb"�h�5F(*��h*�VV1V
a,bD�c*�,m V(,X��*EX)���|��s�����6/ǰBQGsP p�o�ߨ�	�vn^�|jʨ��}v	7��Y�J�3%TF���G���iP�UJUJ���A$����ײ����e�o��W� gg;�	o���2�<Q4Mٕ��*S<n���	{ �q�0��ٖ{F������$��Ht%M>�JbA��%Dw��N�K�ޫ�$���Va@�g1Bn�k�f�r�O���vH���TDD�Be)�`}�v@7�DA�x��];��|�O>ޱ`���9�MY"w#X�X���@&bJ�E9���I�nłFÁ"Q�ª	����N7��H-�wfp�2!)�bEٙO1�j����	��*�A���	$nFruQ������/��L�
�s�o���� �����sw����;s��T�p_��'����&�l��}�r"*䲬u�ɍ��Ml��V�]������~�A�`�& Ȉ(��.%�X�ŝQ�ʄ	�ѐ��0N���_6��F�g* �6�nC�ޢ�L���j:4��Y�HG�r'\ϨL�網��]�G@A�Z��O��������&DI�:���x�O�w7`Y�r3�q޵��r�/��$�݁f�*��H(�0�ҡPuWT�ꁓ׻*������$�w�wd�7#9
*����ζ��k��%����un7�����`�eU�KհʨtE]���I �6���Fr�}jt�(�I^Q(�=�Z�88�ʯ{�.��cT ����ˮT����	9�άGg�	LH@�.�JyB	>9��V
�]#�\�]t	.��=�9P$������ي�5��MhUYӝ(�!��ۊ���М9NvL�g�Za �pտ2I���{�X�j�T���Q*��4�.CT�Q�՟�����w��/ʃ�6���[�.v�K��g�vY�<� �;2�ۛ�ݷ\��>ş3�����3�lu=��]����޺�ݻ+cgn�=n��p�nK�#������.���i������W�l�fۙ�p�.�\��r��W�	c�����+*A�wb�Ǝ�6��+�]/F���S�N�d�ܙUǔ���|oE��Ʃ5[����������;Y�k{;K�Lm�=����Cc� ���M[l��r9���߽��v;R�$��嵼x�}�` I����b��r��݂O�#5W��&�D�BP�"���u߉vum_C���&��Y�'�g!D�3��Y
� �0C|���*�"$��S�P��ꮨ>'��k�� �%��֣�e�����X�A>���a��
`L�1"����wgb�H��,�A�Y�w7z�<H-��S�/01C����fGr�	��LĤB�E9���A<޺;Y���V�l�	�ʼO��z�Y%��w�a	����z\Pvg�2u��VB����us��u*�F9[�vy
����������M�n�}5+2�Fv�U�A>%��a�l]l��T�O, ��k� ��qB	�3�|���IH^о���7�_�ld�K�Dk;��B��+:pet[/�R����j���5
�g%�c3;�0qEq�dwUi��*6����m��8��	$���vI%��B�Yj�P��]MtDL�ފ�R!IBT�&�Uu���ز	����Q5}%�oe0	��n�Io�ز*��b"BHʅ ��@�W�+61��ۧ3��������/#9S��.��.��7�ݶ���=�D�L	��$U���~�<Y�"�ّ�Y�B��vH#��߬^Fr�b���O-g������Uă�6�l��n������{���s�S�s���9�W����}���Ⴘuwm� �޻�H%�g*h��˱܁1c��]�H;�]����D1!��67O� ��>�c��Mﺀ0e}�Œ�3��O=�;l�Θ���0R�LH���iՓ��g*�'���@ڮ�� ���v}Q�I��d�C6�M�9WsH��uʍuroiv��;�}X�'f^M����Տ�$kz�������x�B��� M�ٻ��ˍ��$V� ��u�$��TI9���u j�rN��� O��U��u��D��� ��@���@m���I�y?��}� ƾu� �J{$^c�S�r��m�o��ѲB�J;G����7f�3����ns�S��V$�
ukj2���|eB���)LH o�]�d�^,ڂH&�;������d.��&�v�����dcT���P	���Q(�n����Ѻ���c/�ge��X�{ĂE�>�$�4��ː�W_p��atȂ�%Q�`̧� �|ws���]�r��ao)��$����H��>��#WPZ"BT	�	9C���8�Ǔ`�x�ՕB�-滲|o��ʲ �<��	9�PR1��2�.%�lq�qwÑ.��272�+���5~������[uF�!=�{�qR׾���0��Llt�Ǩ�08�qmQ"�M�
JdHBn�m�߈ ��v,s�3G�yH����n����`\���+���S��='�H�J����ixx�n�U/:���ַ.x�\�����ɉ���`0x�+u��}��dK}��櫌���ټ$vF�A>}���2����0&R��vm�����I�R���D@$>��,�}���rN�#2K���-P$jt�f%"J*�'�u߈'��vH9mE��6!�����V	����ܮ�Q
bQ%�V���ݺ\�%T�=��V	$�o]�$󶃮���$b�4�#�]�G-��A�D����wv	y�5�i�99rH���I���|�o7�u��U��;�GiF|rQ�_M�g&�S8<�^���n�����^!b��WC@䘺0��74�!M�����<�:/c��^�(@n��f�����(��(JF��b��I�s�r�B��9��6(x��u�c��!�juC�/n�ò[�䴝��.����ݢ�>u�K�w;#;�[�d��Wh��<�Qf�t���.=��5�(�Oe��4�l��wd4fO[n����zzwlD�m�.D;)9컊�x'q�'�q���'�����A>������%�+s��V���vn;:{g�tW�]�ms[����m �f�d9gnyv�������RP3"B���]��H8�]� �睴+�h>�ΑT{��|A �z�Ȫک��!)1 ��@��'��)�Ù[Eg82��ւA$���ݒHy�@9�����2ϳ ���$��7N����}��`���D
Q'�F��ٱ&��� �u��	w�B����Dx�JD)�U	o:��1q��eR��[�Nջ�Y$���	�7��d%cg�a� �]��9�b%3�E�36�	$��CbKZٜ�H�|	��s��A���x7���{��0��9�hň-`H��6�K%���� ����!I��]��k�YY�����PFT	�A�+�nŐI�q��$y���&Y��u�ʬ��_��t׉´䂤�fD�&�l�e�" yṪ�9���!IC�X}9��|�<">�ep�j�Y7%�����X�5{����M�
��n�6=��Ӄ�l3��nM�(�3)����]�i�I��b�H��^V?�~z���;~�[D���RL��g|E�ޫ �H)=J�fc�N�X'�}:k�y��`Sl���̩��V��`uS�(���G�_C�"	�;�������6�ؒ}���x�s'}�2d�2���λ�|w�������`�=7f��8�,׉$;z�� ���ݝ�&�q愮���IL13 �Gq�y�v+{n�ֵmS�sրi���tĨ�;��f�b%11($�F�37�� ��:�	=�: ݫ�����8��Ȣ@�ݪ�$�X0P1dYv|r��p�(��Ɓ7}�VH$���	�VyO�eZ�ʮ6O�hv#	RP3"B{RIǹ�,n_WK2H3�P��o������Ĵ�f�m���%�(n��z������`�e:��ߖoXlj��*�]DQ�N�4.ed�� �u��d���s��6�b&H3
�2aQ{ђ,���-��ݺ�Y��$t�!ԑ!�$�}�`��^"T)2faH�6�uY%���Lf�"����� �]m#7qؿ<��G��,��8��uu���:�^��R�[&�7g�]W��y��g�ҙQE5%"�s�S?EM"��������'Ǟ�>�Ν4`�{W!it}��{�O}�iG����v%ʴ|rru��(pR���|H;������5���fNI�`�ʁ��-�D���p�+�>ǚ
�.a�[�c�h�I׸�X'�:t��=7PQ3"Bv�e�׵g1sg.>3��d	3�H�N��Ysl���Nd;�7l!3�;o�ĩ��,h�d�����R�N��=�8�i{�- ��@�.͊��Y&���b4��Oq��e�cc9|�R���p�G�}|�� 7��<�4|��d�?�2uu�?�}�p ��}vY�O�+���*(�H<��k��{q]<	mՈ���9�9�z�4��L=���J1*L�)��������>'���u�vf{�wvX�|K͝4	ܙ�B�ĤB�!W�^u�$·�K��B�#}.��0W}�xB��U��N����S5))T�h�s�G��;[�@ 4j��Os��霻��@ �r�O �;�ұg9�Q �R����'<O4���k�d��H ��:�� "3/��'��ﲎ̘`R���$��&$�H7sp�����I2 #r��U#����[�fN� *jn$�U��3؉(�3�� B�Xv�Q1��VK�����3bZ�U`�T͍���<}�n�M+�sD^�z]Ս�vZ��8͍�Z! A�%�%�i
�j`q��c��ui �}�A�j�$���rdί
��:�߽�{*R���J�c�WF���6�	W4���n{_,�{�v��5�5{;��xt�&�=�{C��|���*���.�����:�OV��65϶�ک��ش�Z\��*��D𭊬3��B`����w���R~9\|�i�[����N';����}|��==p�o5���;1oE�q���:v	�C�Ʉ�w��O����uy��3"-�.�������e��r���GG�BW����E{��s\o�����`��}�46�������b���q�����3��qw#;٣�k����\�t��K^��֏5���=�9�̆f��"���@��U��o�>1K��ӽ�ti��=-���o�	|��!�ר�u���ggMCv�5�1O&���I���>� �.˶��Q��[�+G��2���d�{�W��&���~�WdM��6��b�3�p=e��
.��e{�)Ɔ)\�===���y=����3w9��:��x=�ݹg��ޚ�<�	����
?��JlC�р�2.$aӷn�$�4-\�Q�)���Ow2i�T�e���5�$d�聢�f��=����7}��uF����A9`��Fl�h��)��^/��}�?Bڝ�KN���(�����7�����Bẟ$��zF0U(�-M�,AV�6�"-h��b�Y��R���mXTPX���j�-m��`BV�AX*%ePcZ*�0AX��,�(Q��V,e�&X��F,b�!c3B�KB��DQb��PDX*�(�
,Z�p�0�DKj#���*��QEŢ�VAb�QE��nma*(��b*5+�`���j����%TX��\!�)�YL!�Q�"�+��͒���U*VE�*��cZ�ڙ��iF*1A�F*#�A�ŕ�UVشC-A0e�-�\`8[e�B�T*�-0�-���-Y���b���qh�*8�b�D�R��*�R�-0��J
a��ű��UE�~�?6n�욋v;"��z�<�)��m���ĭ��;��1�w-�)�q/e��s6뱱ls�*Md��-v�v-��I�2��r<�L7k"Ʊnj�.�+�q��+�v�u麽�z�x��m���܆ֲ�=$�r�K��\�|]lvدvx��l.�Yݬ�;�p�� \�݃�3�;p�Vr��93�ѳ�&��.�Wm���C�cM�;o��$�p��#ʒTaiN��]c,v�����lG3�z�ö�E��o2����m��綩�0��n�Y*�#:�r�\6ŷW*�Z�Ll�!�[b���γm1<+���;= �Pv).:�v�u�53�Վ���9�	c���(�u��ͬg������Xȷ.ڛ=;#���ɵ.؜���o7�W�6ҹ��gzL�ls��8�{Ŵ7	v��!���#���cթ��k�F�8�v�Vy^�5F�ya�\87KX�V�.r��v�����^���8C��箹��a�V�Vѹ��y�T�f盻rDnޠ.ڸn���Mn�mwbM;`�k�F���7`���]�u�{e����q����o-��klclf��z. �md�+�ݱ��ɸ^�nz�u�l�mLGd퍞�0��v�)���ȽVǓZ.{T�f��ux�۷q����e�5�9���;4���)������;i��\��x��[qrl��ػw�����]%���ᳵ�N�c��\x��䭽��C��]W%��k��9����n�xz3ۣ�J����ӛY��5�]��O\+�ے��ki���ú30v	�<�����6tX.���f;A��	mjѪ����W"��u���;�w@m����k�:FwЩ��3�a��»m`���N���O4�G5�;���ۓ�l��Rv���1�k�v,y������c������ų�����·�=���z�l���<v����Lp��v��z<qb������栴�bb�i�R��z8.�Mtv��g�f
�����[�Ybc��IK&3��7]���@�ݧ��-�3��x���X��G�w9�v��i��)�l���F��]���W89�;m������9���A˜ɘ�[��@p@�v:9�Oc)rVSaf��rn�z�_9�;\X��nb�ݶɣ�C���ݿ<�۲ur�ȏ8�6�͡�f}�lN�Gu�n�l�v9��g����M<�v)=���z��M��iK��n�.�n\��0��<鍮Ӗ�¬�ڕo$�ke������t�"�G��ٹ�� y�s�`�]�7�NZ����Q1��ӕ�{� �n�߱%�$b$(��3
D�-;��$>mO����OM� �ٷv@�[��E$AYC�(�=l���"s�ެ!
TP�&)9�:�X4w�� R}���}�8 ^n��I��S�H��bY�b�4��Y�s�{�S�="u�`� l�lY$ێ���:�V��PZ�{3؃wa*��/$�6�� �N��)	��4�`m����'o%�� [=Y'�9�Ƿ�Ւw����$*"�L�m��Нr/=k�Χv�D���:0f��ѻ/�ީ�D�)UJ��g#��� �8�Ʃ� 6z�H���1��g���}�C�˷ �:�_�y�TUM@���F�N:2'��RB��}��H�ΐ���A�����5E~8�Vt�{����MBk<�[�r�����P�t.2l_���G�\�k�����Mmu�>$��{6[��VI�"�����ة������f�%QU%*o�ӻ�� ��R ����[���_L$�Q�ٳ膀Kf{&}�
���!J��T�����I9�a섒\��U� ���L� û޺�Y�}6_��4pD��ȸ?�'��G5Z��R��:��� >��wg����E�E%�W���^��Hr}��4�茶c��n�仳���Ǟmņ�n�:�G��<ɗ�ђLZ�&BR*���A ����Xr	��b���A���v��{��{3�Z|�m?̃�����s����,�TDJm����,�ג��q�m��̦ �ٞɟ  C�޻V@�7�&��NϹZ}{����7wA5T�E��6N��� w��DXy��^�_{���H�J!�2˞y�vU�½˔'�)�� �u�N�7�A�Dx-S�n�a19}û��'�p?➚ ��Y8�3�Ib[��J�f{O�1�"J��J��7�W��~��Dh{��DA�	f��݀ gf�� t��ϐ��!
TP�&(\Zv���y%�z��uFb��EX��Pq�)$;��x1I��6-t�"���_������XyM�=k<���띳����l�c��=5��*�+c��ߟrqy�l,|"B������"��M��p+����S6 ܼۻ�s �
���LK���ϐFu�G�dQ�nw����kq���l�)DumN5�Z}IWvQ*D" D�D�� �{v���#{5�8�=q�ֲ�g
��ks1�Fu�ۈ� gf����r�Ț�B��ED��'\�ty]�)*}� ���j� >�ݯ4 hvL����G7�{ptK乼��4�.F��X��qCM�mD^���O<L��M�����\��=�}V�w��Zzw��h���s΅��M��q������ɐ���J���I�&dM�{�X�%%�n�	6r��*�����˻ ��v��y/�]���.���X�<żPa��BD!�=�z���8���ɻ[u3b�`��^��wU[���AU�b��+wq�� |�����dϐ#}{��&3�|� Bo���N�G�Z��R��éS�R	O]!�wLĚ�ȼ����H ۻM�@�g�g�K�1O����F��h
Q��1�K�������>T�ۗ>�M�r������"�sv�d�=�>Ͻq �*d�&�Nn���r�2���b��WDZ� �9Ȋ�yV8{0�K��[,��UMR�%��=�>� ��kp�{��1z#w}M��3�3�����b��1RD����Y�9k^,��bC�:�JL[�2�&kAt�i�O��3ofK3w� ��	�i:�,MMdY/�߇�n��=���q�t�n�q��U��d苶�8n���-:wq���z�c��逯i8�8�8���Y}�..5�+�7%sp�z@���7ez�ע{t�BY�4!T<gI�N��v^�ƗL,Ƿgn72�<oj�ܗ�׏I�dsh��ˌ�s5��p.��˖q0���n�ps���Q�s��Ɨ��LnyՍ�q�m�ɝ��whj��ώ�2w�ߗ�#�{?�h;q�=9;l�/7'�v�:�dݲʽ��'Vvt<���ߟM����"�V�F���� �̟P���waJ�n��	�q.zkd s�}R��݋�� 2B*��-��ļ��]h�ڡ�i�1V�H�q��H��u��IM�(�;����̜�TN���&hdD��P n^sq` ͹��!����@d�T��E��;V���TI��'}zY]
3c�/}�"$�W�T �/����F_mO�~W
]�$:oj|�u�RR�����ז |�����7�OG����>=;�> �w�n"�3�i���y0݌�<�H2#�|Q�����9`�펗<1jz�O���gqtB���/�����ER�E��3�����}}�Ցٴ���+���W�zg�g�|y|��4��HFL̓0&�$_o]ZJ�����3�����S�<?�d��;g�W>I�iQ��=+Yn0 ����l�n3UBB�$��)�HވRE�~S2?���=�  }�}�q gc�&ұ�ȩv�",$��Q@*d�Ty���A"��ZI%�L�Μ�:ͪ�π ݾ뿕��e��`���&}&JQ�Z�V���g&TS��E1Ÿ�w�$�׷��A#��ՠ�-�왋k�u��"��}v���#H���
�Lh"v���H���C��-�Q>�$��w� ��\شIiv�W��;�(RV�����#6Nܜ[g�6m΋����➊�t�anNW��nx���7�f
B"T�%_#|�ݫ�A"�ՒJ�v�W��;Dը3;{�7Yك%%��ݤ᫒�bI��*j$m'\��+������W}{��X  G^�6�H�=�>��� ��:�ͩ����)���>�S0L§��y� �̟* >A^�F@U0)�`C��l��QL��I@4< �e�"�|>\G_`����^����hCY����E�w������OF\J7��33g'���Б(-�n,Z$��I(�N�"S$"�Q�2�m��K����y�Ae=tπ@.�ܘ��J�f��qh�6��d'�,Z��+骊������Ͼ���9ڳ�^Z>e�R+�>`$�3�3����Iw����D��@!Ė�#�=��\ہz�-����d��^��Wb�pFue��G�q�����I��8���ܟ|��7���� �q�Dgǧ��@��L�Nm��D�� R�����vD&����|;�L_A���DI/+����I�.{����*#9�e����PUM(�
�"e�9�@ 7���j}Nթ�]뭞� 	l��ϐ 7��j��� ���j���N#G�ѵ�=�Y����!��*s��@ d���WS���^!oO�n}��P�C��֓>#��<����� ��W�^���o����V��8֖G�a�a�X��L���^� zo�>�;�yDD���A4C��gv��`�A��j�d����\�� ��۩��k� ���`���W�9���v�D�(1!���
2 �g�z�c�u���s��Ú��p4��u_�?~�����P4a'����1�sq ��}���hm�ްf����$y����?`:I�� ��fk$�h�h+,*ދ�'�c��7��2_l�@
Ǖ�����feLE�`�|J��P(�Mu�$�T���	T��GmS��R:H�y����fB	$�����9�+V�g���F�G��KY����9��$�O�&�<>����c�2�m�����n����X�b��� %���}�g� Qn��v�`�h-Z�H�om�E�l��2 ��� +$���۴z����T>ʳw7��K��,KS:�,���E�U����oS�h���Gy�Q�w���|�'��G,�ɭ�ܶ��B�K�b�F�"@�ش�ͨ���_\q�k��-�^��N�l�M�Q���ҼAWkV{���=v$�ݯO 썸Z<��(#&\c�[�nۤŝ�R����Ń����\]��׺�ɣ�8��M�6�N�-�7�:�\�Yvi;w��;��G[�A�퍻��M(���(z�޺�.��#��[�΄s��=���]����p=��s�����/6��]M�7]u�]*u�k:��^-Ʈ2U����ٛ���a޹�в\}��}��҂��?����q �h�g� 4���:k��l���~�6N��ڲ�:^��tqj+�)T�7�Ｈq^똟	���L���`�e�ˈh;=>@�QQ���E���[�Q8�i
E*�I�mS6;f�]2���M���d��8�qD߀�N�O��됥��)�U{����x�qQu� ��� %w��AM*���Q��g�D���	��IZw5,;�BLQ�ۚ@$����z����W�q�yt� ���@7���W�AN�E�z�W"��QEMr�1�5��cU�;K̸�m�ΰ��,��i\�'�/�A)I0�Mj�ٯ$����� y����h��WH.���Ȉ8��&�7�׈�T����,*��38�7��Fn�Y7�O��+��
ӛ+y��]*$�U�Mc9M���p�E���p����m��ZsA��	n���ey׸"/=>H���j�m_�q=x;*k�}u�0�ȍϊ�������~� 1�s���_�t#r��@���{���z�+��4� ��}	�N]֙����A��F�&��l��� >o���/�m󓴔gS��+	5I�Q{p���i�����!$�G��|���w���C�MG�@"������l���ޗFtROd,޲�.b"A�(�jvr�`6��<�{i�n�����8o�e迟~�M�e4.3�5��D7��� #_m6�]:����׻k��os�Ղ�VD�%ST(�T�F����5Ǟ�Չ�q9�A.���D�%��n�I����5ZP�9��>J%*�[ݶ����v�����0�N�f��o~f��j����yv�c�m�C���!	�6�@x%�z��l\�r�sVv{:{\g���v�:�@��@�L���7���z[��gcH�j���|WH���5���,�!�>��h�ވ{D
-��#��'y�q|�8r8��dZ���e�վ ������	��\���&��Ŕ_1���Ѿ�xc������,<���B�~�"{�˩��z|��b^1y�r��q��z1g;���p�>��v1��6��ͬz�W*g-fP)�2���'�V4$L��>��A�^�����*M0�p�7�W�	�������7��\i��� ���D����8�g?a�sբ�y�=�|�k��8�S-[.<��f|�֗��ܽ�1e���?s�c��r��g$Ր���L�;��LPU�k<l/@�]�Tg�I�¤Ȋr3�W�m^�w}9�������LY������|����m\�ݵ��f�R���jX�*mԟ93Lּﯥ�:c�V;� �i�c���b����i51�*$��&�������ӷ���l��� #���	qʅ�gzy��O���}�w�u~�W�D,f5�{�ݞP{f��ugK��Xk1���̝�٧���4=^�*K̡���~�;Vn�k�qyrY[�X�x����Ǡ#�=p<ъW`�_�ty{������}�GD���h�R�')}w�nvTӷnx��n�FMVM�sN:�N���g3�2��O��U�Qb�QEpʊ �b�YiX(�m�Z���H��AV�.-A­��ZPV
"!�ciUF3�Tb�J��j��TQcT��."�r�0��,TR8p�TE.i��DX���-��j��Ve0�TQE��P���T��+[Z-F��eAf-�XV��0�Q��E-��+2�c�UC-UE��
Z��W,���67�ڥJ%d���sI�\"�V(U�Ѫح��0�DqiE���
�[V�q��
	l-���U�Z�+b-K���QVQ�ZQ�մ�Z�J��U�K-��q�3Ym�R�%eE-*���km�lX*�r����Q�-]���m���s�숁>�i����>��������>٬$~�^q��3��d@�����W�S�[�]�o�?͠�ywiX)47�HP
)WЙ7k�@ �ؒWl���ůuy%��٘$�|���G�xl��~S����&
�"�HMJW��u�sڍ�s `�tn5���!l�VݪUMOf��Sĩ"%_#��v #����I �f�<�P�J���t��e܄�I5�u�K��ҵ u�I����ϼ����Ջ�<�����X�+��G��������z�~�/��dLRU5B��^s�y���^@ >7F���:��E��_e4��^��K�}�(�UG�4Z2���k���W�׳"Ȏ������ɨ� w�Eޙ2gg�Y���}O���J*]�cK����%��r���ߎ�[��x�]$�5�q;�h�}�{��}�_-�nOzn�_e:�[{��^u6
9���}JQ2�S�$�J�yݚ�û3���w�^i ����{� <��YI� ?Z�fG�~�}Q|D��N��g��l����=�$'[��9Wq_�߁����+�Xw��o�����@���HON]�jyF �ٷp����p��̯G����)I�J�R"Seg���G]�k �����+�����p�OޫG �< &�K��R�.�5}����z�GHҵL}����y�����DY�W�sYN#����y$�F�_^b7$<&�12��V�w�9�.���=8{5�@|��7h c�;��O��э�G�	߫��>��=�(�UG�4X�� Amث���ދä�����)e�y��PH��sb�W�r�T��O��<�:F����;ƿ�-��"�[��F��o��J�-ނJ[Rgf�a�/f�9�"�<�z*�R�� ����/�I�
cv�ێ�+��q��)tj���:j-��O+X�@��8��[7��oSڞ#����x��7%��İ���$�%��v^:Ƿ`�]��dJ�t��=Ylݛ��!��n�O5��wx��W9�m<����أ�us�2�[{	��TSЧ�^�������\���.Y��9�ݣ;ӌ��S$p�<��b0mV�+93��9��s�ny��u��wi�]�x�;���-A��9	�����7,c��ث�cU�TA�[������&���w>�  ���9��o�ݥza�m��Ǿ���H�{�waDa�hB�"���1��˺�E�>~��d[�	������ 9�ss� S��� ��_gw��X���K� ��wsDI�L��LJq�\�X 5��m�	*��־f_o�N��a ���n"�FM��I��p�uR�csJ�u1�Ի�%��|�~~n�"����e��zs��VL.[��;���i�F�~r��� Cs5n�o�8}��La��;�2�0�+�a�շ�v� GM��L����|s�;���s����=Pp�������W�Y��-�S=O�q�ܽ̀�ùW�����n���=�z�X|�4�֩�-��Ax����Fm�e�eݐ|�M��LS�����V���g�ȒYb�J���t�ű�^M��Y�Pf{qᮈ_-5�����!�ګ4���׏�A�S�'���n�@;8�a\6�������A�?{ ���Wr�E�}���|�W��dz�z�o�1޾�����@�e��%	�X�&#{&�=�*�^�۹�U����@|�M��L�����ӛt���	��E߂ڮ�.��7�(4�4�v(�Ivez<� o7�_=ˮnlmLr@>Ζ��<�ET�U*����4f��#�|�s�{8��W�����.����,�$גA]�vYɥ��U�?tg�����=���nK������ƶ��+"�=�ss��P)��]�~QQIT�
	���8}�S#/&�� ���쨧��1��z$���i� :��@}N��P�QU�9hy��j�7���V+��>π@u�z< y�w��������=v���O�X�@�5 7���;�x�A�;[�����Yn��s;.�"�j�Xف�J�4:K�M��n��"�+t��٪}OS�R�u�5�j#}��/��\��~&�-��.���)	��@�e��(�̜���db�� �MDx �븈���}��瀽5Y�O� %�uz=�x�t������+��=�` h�]8����&�
���� c�۵dD�����Ƽ���n��9�!pn�u�â��.{�m�n���u����k����2�|�}ﶩD�U3S59�=�x �o���|�l_8�	do;{.l�ۉ-$Am�쳖�)⊉J��D����?���X^��٫� �D���� l���C�L�8�k#f2���%9�
d�(��,y��j�����e���X	$��z�=������H��	4��SQR9h���_��?Gmt���o�o1$��^qmŒM�<�vs�\K��U�������QȻɿ{�O=4b�������K���M�dg<���n�ߞR��ȈD:F`N�����̴O&����)GqAP�/��.ڦ �s:��w�̟�C~�on�,��RI��iZ
MvP���w.ICez��/<y�	���)5��s[��hs�E��PO�c/�H3�%0D��S����4}�S n�y�@N�vnA^�j/�ܲI-Sآ�q��ə��H�������7� ��^\����K��X ��a"[ޚ7�K�i���nK���4 �`3�fD���o�j���"w��h�^�ܮ�UDGW?n��@ l��i�|۹�p�Uq��!@���&(d{6��Fr��>��v*��qwk�7䗂If=�vwa�\Gt��w���!�l�c� �ұh�������@ {��Ykfi��2n�#+�^�&[�0�$�=~lo뽳b��2^�����'.a���goI���#��$�y�Kf%pj��f�o�֣�m�S��(i�-����x�f�s���x�/YD" Q>0I�
bA
dA+�nm»6Kw �]�x��c�iZ\�y�����8�ķ9�wP�cr]n��]6"^m� ;'nG��nI�6}�=c�e����8��&�������V�������z-���0�=����C�\�Yŵ���T8�Kٴ;wj�����n<��zC�^5��D��/�OP��<g�h�A\��ݺ�b�p�ba�Y�fc!����\�������2��N�b�K.O����>m��}N��k�@|������n�Nb��T��	��i� /s|�B���3bS�~N��g��$���k�g�b�Wy����� �{٘�K���:��*�3a��놨X��bJU2T�پ}M�.�9��DD=&=�gs��;=^�����8�E��;�MT?b*H���@IM����:�<���˺� {�wh$��7���RW��6'ʸ�*�������g]��A�_��Ǡ�Q5�^� ��λ� >�sE{��G�f�`�݊9Ģ\)�"F���@�fػ;uΣ/c�:eշ<�Y�6��.�&f��$ȉ�1$���৻f�$�I��V����M�s����sPwwU�m#��ݜ���d�F"S�-Z!Y�d����ZK�����ū���o �8���EgF��^C/��7&�ra��5�&�-�H�w�Á��aQu{^�  }w��v���&�I��3N�,�	 .7nA�)%L�ҜmV���k� ��Z��|�H~޼��#os�� �e����=�7u$��:��}��fU��WN�}�v����  �e�ˈh7s��ߙ���@N��X&�8*H���@IM�>橀$ٵ�f6g�}7��&���os0$J	ŷM��ޫ6�ێ2��YSzg�(fB�
g��xm-�۵n�zx�Wi���5ӷ���l��A����PS'�A��+ǽ�1��V��L�uzT�G�g{�#��wY$���l������Z�-<;��[�";����G�af�����h�g��oz��a(�G�u�67�9�R�2P��T��D��X&�A'��V�	 �M����+F��{x��Ī3�h��z����u��c��	�z����ݞ����N�Շ{KSml	�4Z�j𸽌W7u�ugN��i���:��X�)��Y���}r�AQ>�e�Ӻ�y2	��	���_�%{�Y&�{�~;itq�5�ǐD�}-��<�n�H-��uil�kxH	��y����E������#o:��>��{.�7ݤ���۞=J�2�ASEV����r������{m�W����˙q�f_���~�L�}UJ�$�w�8y�*b@|}���+�컰���c"��0����⥷-w7��3�c�	@Ϥ�U-���qiY�Y:���`D/;�H�c��'F�VL����w��<�)T�LMDUH啽��  ���j��\��λ���z�'�9` �o�0����*:0��M}�	2��Gb�+0��/��y���� �}�_q��M��s�yLf]�E*�<��0���Ѿ9=NW+i�0ٗ�7-g��'�Ue����&� ����Lѱ�m+����טxIƯ��ԱH��7�����H��SV�oީ��6�A�ez����=���N/�X�Q�{��Q�Q5��x�LN�T��-��mؽWN�)[j�H�r��\�Q$����V���&�T�4>��=�� |{��X l��l�l�ɟGB�^���> ��۵e?��T�G�U�%y���5L�޻n�;Vs����o;n� >6_l�!��7����9���m}j Q_E1C=��v��G���/�ΟD�s������H�y�I��Q���DĘ1$��s�u�s��N�k�nj� �}��� ��e�	ngy�nڞܔu�\���{s$ 8ҙ�*
�g�-XA&[t��s:�¾��l�"��}w�m-]y�2�-�s��ս�$ I?���$���$�XB���$�؄��$��$�	'���$�؄��$��B�� IO��$ I?�	!I�	!I`IM�B��@�$����$��$�	'��$ I?�	!I���$�!$ I?��d�MfD;#8��f�A@��̟\��o�  ��    �       �   �          h       ��*�� �    4 � Z *�� �h��QAl �� 	  
5� @  �  P  ($  
   P      (    � ( 
 @     (  (��7��*�ӓ���s�%��^�V� 7���<Z�hr��������*�9��m�A�   �-A�Ǽޞ�����^��g���� ���x���R=�@8z%�Ǽ�.`9�M��^�ۧ�����mi �   x   �@���g����w�0��u��Uf9��Ex� �a������ݫ s��ڭ�o;�E׼ 9(�������t 5�^   �y {�R�����{h�@d]��@W8z �� �2��Yv�4F�)�
�  <     � ����݁޷F���s�F��y���(0;�s� �� �
\�Ҁs���`t���xЁ� �o�N&��i�5�[�  �S�ҝ ����)@��� nzR����G��R�r���()�gE �����J^�������s٥ U�j��0@!���)M-�x  x   P    �a�d 2�w���� vJ�j��D�9��Y h�  ݮa�AY��d4 և�  �yt(�e�"�p 8:#�*Y����҂�� c�  �u@na��ruG����
i@�  �B�    
 �C����sjN�9ځ��`Q�p=��1�:�!�Nl���� q���n�W�4
 p   �y�;9� �p 9�C�{��'�̀v��Y���Op�y�E��@�:
=��y�!��mR�� )��R��� 5R&�j�2 Љ�UJ`�H  )�SD�JR   Jz%��H@ 16���q��;�M�V��M3�\��e�V��g��cv1�����`fg�����fa���f`�a�X�`fg��fa����f��a�f��������Fu�7�h����0w�����3aX�R͡�Q��T�b'��A����q����"�7^<x%A5��b���̫BwI�$M���vg*�o�f�/�A���`f�gU�����J��&���0����G���1�,Cf;w��؀�R�fk��Ʋ�A��p�%�1I]�'�Oݗ�v�3X��,�ͷ���w8:b^i���M<��tLy;t�k��r>���^m�7��R���)ȇ��=}T�/ �o;���(t�^�S�)Yά����/-��k�;����xݒ���-u������tG��qae�ݶ�5�4[uG�N�c��Ν@q�oiP%��:�N�c�B��s��P�Y�t�f�u[�(DҶ� �J0�x��![ڠ�`6͐��Ʊ�v���]���a�n,�Hj[Ib�0	՞��'�ᥐN�E�{/��z]�^�s_Y�+���lCw�D�WdXz�.�r���%�^�k]�N���"*�]��Q4�2Q�w�(��U�c��*��VG�.��z�v���{n˨X��xnq�X�\��7��<Jp�z�Y��v�s�g#u]��Y.K�:��j� ��[8.W�a\#�����p��&�ߚjok�3��\��)�ƅ^?�����{vh	�#�&7����:CH�N������W��53�N�9A��/Fq\*����!�Ǽ��lŃ��Ν16��z��k��9-pѨ�C�y>L7������C,�N�4 pD,�����0�I�Υ=\�5�yd0�ݲ�.Ҧ��5n &�4.����2h,Xk�ιFm��ce� ��i����Ow����C�æqJ�v٨v��-��!�E�{������m�_��R:ZK	۳�(�]�����qtP
ޭ��l;��^�����8�lFq��e}�h�fwG� 
�8�ͽ���ݢ��3N�gw�Á���э��3�q���L%�u��&��yVfZs��EӰ��t�7V(, Ō]��p��������ĝq�x���o��o6����8m��F����wc���� �5�z���n��I�<�ި7 '5�'�^%�Z�sm��9Ntu+%�t��C��Ej?��)�����>g�w&���
����tM)��;���k�p���P<��!o7r��9��a�eP�j�r���">X����!٩�\8�:���x,�v(�*���u�MH� ;7�j�R�5�ݦ�ƾͨf�L݅�͗-�[գPp�8(�	ObȞ;���P��_T/̓F�0�`��r�D�����%���t�Z+tՎpZ�B0U�ǋPwYg��sF�Y� Ԗ��y����#7h�I'ZD
i������\Nv�ۛ��
�-cHYus�u���8&3OsF�p�<_!���X��$��SӋr��J�lU�iwg=�VlM<�T��敕M)M[X��ry�9C󨖊����]�ã���w�	|]��mx���s�G7Ѕ�LQ�R��h��U���ö2�1��-h	۷�mE�n�y���ΒW0qb:�]'r��ڻ�Eۉ���{rI�]�ž{�c{d�&l�I�u���sӨ�7�B��{���z����ۛ�2��Y�`qRv�[��-�=f�>��28'��sN�I���V+��@Eƌ�puk��S��ԇ8�0F�N�>�6ȭn������eh��>�@=.�����#���{qÝٽ���شX .�q�N�/@�"v�7t�]���:f����_Q1i���d�"���j�E�M�v�q։ÃU�F��s�.���F��C�����&u��j�Yw,٢njNk���!�T��-��a���T���Ĵ��i�.������&q	uQY����B{�rj�ԡ3(s#Xum:uoj"��ߡ�U7� [;��i���tAh#�y�\��0m@�6˹��%��-�	f��y,����4���'�k��3-.��V���3^m�7 ���G(F2��©��B��ܚ����s�c�^�&aF�(��nq޼`ǈ��݉2$��0Q�pC�{;; Q�4�.�{��px�wWg+�K#��\.=[�(Z�d9��o;�}{z��������z�^��ef�5 p�0���2GI˻����V��Ut]�^����t:7s��B��uQ4�p��v� hY�)g�éq�@�rM�x�l�{�{�U�,�dw �(Fu�4n��Q�%���
���561輜�!z-q��z�;y����fw5]�[F�)�3a���6�k�Bn�܅v��s�|9N�re��ĭC.��PE�`0/�=f�5�kE��� raf�[���Z`᦭Hk7�5���D<��Ν*���R��h����Q�6������w�7@���	����2��Es�6A{���z���4^K:������{ٳm[�ۛ���ደ9��é=��N�%�+@G0ւ7OR���gt�$v��N�ᶓq�v�AT�ئq=��_I�����$��wB}�{�-���o8��X�����_ݔ'�`ͻR �ӏ\m�b�_;wY��z��.y�j�T&�U�څ�g|�to�}��i�Mof��%o��w#�p ���7��������J�Gu!�q�3��������>`�:b����г��ba"��VX�+��=e&E������������Ώ���9�0�n�)���W�s�tyb��˷+�Eɺ8=ɦ��w��ÇnQM�q�>�0�-%F������J]#ꌼ6XW]͹���s~.�w��F��N���v�>���x$Ge����Q6i��� �i�\$V�a\r*�ie�����n�2.�1I��3vb'u&�I�����s��t�����&�teC2͇� M��Pcv�X��p����d�;�n�*� \�n���,�6<�!v�,c���"���ݓ9r�v�;�}8������q,*�N�o͗I�bq*0�֞�����!�9)��GP�x-��j������r��u�a�U�lpН;��!��{�Ȼ���y��G��M{ԇ�9��±u��`��C_�ȃGV��q��s �E/�TX-�<�;�z>��;4𫸥�1.��Pa]�Ch���檄�#�ƤNOh����d�8��&E^P..]X ����.������xw97�'ô5�V�����s���]Z�oU��3]�xl�9�{.�=��X�z#��������"�D=�m�ت�0�n4w���}�4��$��`5��y��Ǘq��<�{�׃"�6���A���n��#JA�q �guO����9�F��ozW@��*�o	v�]qմ �m�U6x�F;�Y"k��ǣ�o5�hr��M���p9���{;V.���y�=gI�ӜE�45� �m�î8��G�t�F�eH���J�am�ۣ�ow�F��O�R��=�M����;瀜Fao��Sq�W.��$��V���\u�$0��
�vv9��Fv�+i'j��!;/MXz|�f���Jh`��ňm� ����߯5;���mk����c�9f��f��47�d�Kl^K�j�vgZ;��;6�Mܣ48ylp��v(����U$t֤9@�θ\�u3k�ҏW�u��?�u��l��9HU�Tj�nA�r��=��-E�M�/�ĶlUʕǢ��9(7�E\�Ǖս�n���w!5�ʧ�)��{%o/%�`�;�_�5�r�	�Z�jV5�ˤ/9��d�j��M��ZUsV�v9����T[�x=���u�{�];��K�f2��B=6j\�kE��+q�k��(Ïǡכ[�O;�k�F.|r����va�=����
^#(邇p��ap ���8Ӏ�1�����v<�R�CL��RV�u�B��H\=w���/�M�2<{!JE��l������N�¦:���N�^�\3#(�v�4�^��4��yGV��A�ee�H�DF!Kǡ��>cU\��ϧ>��j�5A���vr�H �0DF��R�0�ڻ&ɩ�3n�ᛁa�U�qփōy���|�`4wu�J-L�A�8�X�|��\�vn[��=�U�`�"���y.]d�iÇ/6������˛/c���a��~��8�j*��G ��Y˖�gA�cRs�;4|�J^��Цo�3a��"�_v�	�鸓�� #��םC��.���0\ ,�7W�;y�Q�o��ø�����^�O�GݜF�h�-	c��H�Ĺ`�G��:9��gGn�kn��<�FՆw����K[��2�E|OW؎��,�'oM;Im��[�{���z�8Nl:��ۃ^�["�on��}��|��� .o��"OC��ݠUaS{u�]��9��Y���W���3�9�ŸV�Yݗpaە��.9Ѯ$jȒ�ct^㛒L= �6s�P�;6���Qwi��A^�� AA��v�Jn���qd`�	�̀&s[�~�{��B38툼g 2�S���T2;*��q@2*��oݖ�Q	=y����(�!�cD��'95+���A���r`���ݪ�z�ˇ�(��׬�sB�������m�:�\F�9nnL����#��DK�сb<Mɽ���-�T��\;�wH�WՆӇ�4H��ou�ۦ2t�ބ��,j]��%'�u�oL�����%B���m�����w�y�Bl:~��/p��,�A��<vE���ndM�/t�ҵc�d�w�.�i[4+�������wC�.t�pn�qpIH�)�U���{"٧{ULa�(wG�h�#�d��(�&\z�\�9s��Ⱥ���S��q�O�o�{�Y�G���Hc��Ŏ&�]���m������5���m��I��+�Gk�c�#��tG�k��R
j[8�܏r,}�^�,1�� t�����{MZiw������64MWLp�١��w�>�^n3�xV��P�X5�y����Y����H�ۼ4�ڲ�w��O-�.�����L�b�W8q�<�;��m��UXF�-ۺ\��B˸fQ����"�j!���FO�Jk�afBӱ�t�{Yڎ���
[��.�;����(ޯ�C�@� �+��b�ݒ�껢���qݨPZԷ�#r�vZA<��ܰ��-[�\�ͻN�����r�D��we�L�D�d�WRG7a�6tb&���珜�z�����������^�[�(QeA�8dm�6�wە���5�\���hBo46n��=�[gN,��y@a�~l�v��*T�m'S~��q7Nv��Vmu܋W���FO�u�-�:LYڬ��oG��m�P�]bX��)鼁��<��:�#|��a�#��9�l^�M��h���s��]��w��S�2E� �
����83�ݙ��i��׶ͻ�á�9�� �?ZmB�l��=��K�v��on=.��p�q��J�G)�M�D�A�.�o+��v��rl�$ixvf�<@m޽b�Ŀi��t�F����P���|��x�Z9����\S���8�; ���N�ޫLjNQ&�k��d	�L�0i���)^�i�K�){f�
����#]��hg�`�1UE�ߔm,��51��
d^۷A����y̗�]VL��N�s�ȷ���q��5v�زۼq>��V�񕽸ې�����e�79�;zF	���No���z���4+
��r\�iJo`$�S��Jq���Ƹ��������Sd��e�N2(����{z����wfi��\
ꝣ����0�`u��x�6;��N\�caq�����-���`�Xf��F �[��]�T4^u�?�8��9����]���;-�'COKᗊ��I֦�Z6�*��V]Ŏe*F<ޓR��.;�Mxf(�S�J���3��ϯq*���i�>�N. ��7.Tȶ&��0ۇv��-��&N�f!�ܗU�#OD�4����y��S���dݸ�����}��Աfӣa��p�F�ޮ�n=\pv՚�Q{7�����s'Y�^ �:�|��t��gc�XB/5f�qֻ�lpؾ8"�d���8���/j��\�6��3]m=Ț�2tq|>����[�aGt������|���w�E���㝔��ȸD��Y�d]����G:�.ǧ`S"}$��s�tr�Ïh��%T���wd���ib�yKt>u�\W^\E�k�[ �G+Wv/���f�8��ӫ�5.���}U@e-��Օ,Dz�fX�jH�E���.0Rl&�U�JG���Sd���U��txY�n�>ŗ&�8w�:WY^R�ק=����K<��8�k�992�iW*�V-��c�!:�,�_l�i9f;u;�h'Gm��cYiq� ��#Kcm�6\x�3�A�9�֣"��b��azsG�`�LMv[�n���:tbիK޿qyj�^	1��)�PXtw
�r�}�HoQ�y��ϵu�{��|(4��f�9$��6�y��k7��pޢd�3&��g:����74�X��R���f�n��NHx{N����0NL�����h����cA;�`f����f���P0�00�QL�331p�&`�31s 0� a0�P��p#�f
`.fa���fDL3�3 1@��30\�  �@��p�1p���1p30��A@�1s3�30\��L0̉�D���3 �p�2$L\0��28�L���@0����f`G0�f�30���� \��31p���9�`D#�f`�`d@��#� 0�#����dC0p ��s#�����L�S3s�����33p�S3 S 1C1C3300S P���0�s�S0\33�s31C0�f$���`�a�030���<���~�q���?Χ��ݧ \x�s�Ӻx���A�2��[����o.E��'/a�y�����"˽���o�G�m���'}��zW�t@H4UFj��|yO{�������+)���:��`mb塍b)�A�������nn.��Y+<�:C��8�m��ޣsQ�Η�n���6���w�����a�ϸ��b<�*��F<�+	g=�R�6���I���U1��@�͈��Xr{�tE�/cVl�%׈.��R�kbZ�V���x����[nQ��SU#]<�UP�i����������# 8��=YN�V��x H=��,��L�}ޱ�#���-�O�y��y��ׇ|�{��L�	����Af1۳�z6g�@ew��=+�d�>������-wI�䪂���{ٯ��3�j��X�ǜ>|���"�.C����ӒG��9��X^�h8X�qSJ��z�����ӷܝx�3�TA�8�d����)���3��3�������p`�=����/�D&-p�}��#ۛ�/1����H�ţ�Z�{�I�����5���s<c�=Ǥ���EyLGk��6X�'7ݖ��+�!�4��W��P͗r�΄��y�y�=�1q���W`���>�%!u=׌������VA��/R�b�;�\l��m�/SMas8�d�jo�!l�{��rYM���'1�w�vqZ�][����:,������j����O.ya��@��լ)�4,��"ixo��b��c�����b�~�^WE�%b�랊�.�w������W6}�׏����=�=V��n�Y����sx�!L���-���	U�Y�������֛$	빚Q�.�;��ܾ���y�2�Y��2�9�>͘{W��{c��v��Q@�Ӕ�q"� G����o�ޚ�E��Sj]�ĝ���2�T��G�{d����b�/��~�V���w��!9�7�@���]�Lc �̡�{WV�v����(?)���=����L�}��h�!|#���Ƿ�����$���b���xKT����\���>��O�V<jŔ,�-���w��� 5�z�=�B�7
\=�q
lo��h
/M�:�-�oh�S�A��W��m\��]}���Qa{�G�6R#^3��.vx���MPd�^��Ã\�g��< 9ȕ=֨�fO{�{����Q�&\ ��D��q�� ;�v0�t����fj���t����f����9���͠<�s�+P��u�ǩ�_{�g�?`��<��i��۹ϺE�������
=�/���3;�m\�W����=��@a`y�^>���X���"��0���uo.��a�#]��1not��f�c{y>^�&M��,��<f�y#��;��=,����V���=�6e�*��xG��|��>��8\}�)*��<QU�3��3��`.�V�޾\���޽�t�BOC�<LC����)��S����vI��ݞ;L��.Y0x4W����N�2�E�,N����|������9�[oi��'��=�	����>�yc �:d��b�>��>�6F��q8_�7�� �0o:��{�$bkܰxL�d^>������۾�[�e�K��մy�T�=�=f,�={�?��D�:�d�a�'�m~@1�֤���y�ɮ8P��䦣w�����Kx{��m������(�0�Nh3�[�w��~��������^�^{�ޙY�v�56x���ʏQ�͛��#��y�7 ����_��FlJ��������X'y�<�����uf�g�ɯg3ӽ���;/��� #�!豝"���8矺��8�{�lb��>�))�C��j2��/7	�w�z��z����`��Wi�VǺ�v{��v�̠9w�1
�\1{��p��{����7�I�6����o�\f��g>M^ŧ��n�;��p3��[{�wx5q��צ�v)}����J񾫏/	ǎ�3���7�$y2n����=��Tj���g!�6���K�I����0h�GpV�f��O%B^㐛��w~�Ȝ�D(��8~>��=�Dї&O{�d �33�<�h���o��)8���;�`N��3����]|f�;�{'p�T%Q���r�����kk�ɐ������YqW���t�����h�7��׏5XN���M6ԫog���1�/��O\E�}<8}��}u^�07Wr&v_�?��&�>�����saЭ�=�o� �t�w��XE�αů��u��Y��ˏ���^�[�=�V�����_)kf�/
�*n�����C	�Y�v��|w��QV{�9�߼�/N��o"��¼T�)����ޘ��+Y�}�p̖��ʚ�Z|Ojx\�G6N�i��<9�s����1�)r��z���=}$p3�}�g�./|��{J�q��z���_�f�z����p|��R��E����M�O��=�3b>w-�n��Q��^T7&����W�b�8�;�5����i�嵶���{��i��2�t6G����̝�r�u��n��)g�JnjO�!�ç[r����+g�mμ�,�����[ȿV�w��}r�
8Ư;��Ny���KM�ίRem�{8��d��7OjHd��^����s�cN{GA��y��ŪHl�q�||�̵<���C��vÞ���n��2�ٷ��R׸!��E�0;y�<Ҳ����S����a�0�X�v�sڷr8����w���{8��˦M��~���"l޸�'�5�	�}���4!j�^9�DP?cu{;��x�g��J9���=����:�]e����,"Q�#��>X=�C���G���S��jǽ��ՔT�(�w�|��8�í�e�q��쫐��f�s�tb�*�HX)G8t�� ��d��p�)�� ����z�O�����C>��^y����;�
\զv�Łg�r�0#O=����߆�ז��{N=�J��K�n��|7����u�����Nў>B�������&�-�]�׮<xG�Qsg���|�gyd���s���f��F�������l�d��6h�d��Y��r�sǅ��r��O�9/z�OLOT���#���O�O/�$Yɷ}��VH	�����7��v�������T�{:��2m��Ȁg�|��&q��bY[�f*�ܞ��-��x{���w��B��v��8��șs{�R4؛�g���t�O]��vT��M$UG{���n�89�W�y=�^���ˌ#H��zQ��F������ǘm�ӡx3Q:y��;Y��n��y��Qo{W��J��φy��Q�.n�d�z�fC
��5ܬ��f%o�&0��@8y���@~N��S������3�z��=��c��bQ��� ǬU����}tv����;�ln�0S�'=�Wqt5yz:����柷�����i|�����t�3���#���y����=�z3GpG��#�V�Jt���7��,G���ؾ�H�{��OƁ�z�y�������g��n�ZɄxi� 5F]�'�$6�>+{��ӾNӷu]���bK�7;����@��9�F��[a�F��z��mJ�n^w!�o����󏷽��r�VE���?<U>3Ʀ���)�r��A�0z(d���s:n�1f�5yu�� ����� �+�zc6M�5F�5�hܲwx�*[���-��=��ɞ v�*���v�=���Pױ�og��D{st����ͽ^��Ap-�f]��O�*��{�g[4����{z̫��{���'^��I�Ցs�|�{<��l� >��图��\Ҁ˧~،'N���@k��qUÖI�`F�S����ve����^�z'w�q��������g���=��j�b�^#���><��{�1��������8��x��Jp���>=���T��Wmٻأ'��o��7%3��+d��:��&7	��������^n*X�&*�m];%�F��ٗ6Z߭xS��߶��Y�{�0\wT����XGN���,�-�Xq�7z��+�a<k�e���8�M�=� �G������s^?c����Tf��j�7�-�>���
���i�U�W�q�Y�;�fUi��oN���r���>�=S
 [C��JV]�ح�S���L{�A=�[Gq�i:�< b�3��О��:7�e�@lSX�?Ģ�� �|�zl�����֑G���퉀�N+�l�l~X|$����eo���Ż�ԉ7tiZUN���=�l�(�����uqG�v�ݐ{_b����{�7���j~���C;�b��JY;�}��V�{a¢�V�w�جcQ�9���\�H{��Ĥ�.vy^��4w��y���JR�\��iF�֬��ne�J��S ��m�)F=�����%F�$�W�j��c����F�bx&��ܔmK�����=���.���v=�҃�/��w�������:'�yc��.GW��0�'#�tR�H����^IW���dY�ǝ�k�����"Y$`|�;�����n�b\A�ϗ��n��'L��1��7���=L���ܸ=����ϩ�Ƽu�SW�jM��#ω/wnm��]�Êq�[8�.�Y��,�-ҹ�C��[}��q!ȱ�^¨�1�Y��p��׳pz]�o��}�(�������Ʉ�wc2g��C���X��7�K��vK5��-L�M):,ޫ��"�'�捋��:�C�6�c{;ni�5j�0�)��۽Sr��d�R�ŁG�&����>�n�soϗ��嗍C"�v�T�p{�OJn�}��,0G׵a�A;/��{�䖜�y�s�a)�ڕSy%_�#��gw��r͖a�>:��͚�1,Z����sѕ����3
���G}������ݞ9�
�	Ex6�?a�W�W+��־Y3�^o���hX����f'�/@�Knjɻ�t��*ߙ�U���Kr�Pl��&��Wy!Cx��Z�L�ұN�4MyM�De'�n����P�x��T�gCws���ӆRgC���4�~>�4vvN�O#8�U�~��aK=;�D����w���F�G��l�J8�F�#{/G�;������OԽ�__�1���a�P�ݞ���$��Af��U��������\w�_e�G��.��A3���z�=>�,9J$8�K���{7J[��BI�Q�)4�c��xœ	�}֢M�7���<��^��Uc��ZRه2m��}�J�ZAC5�e��곘��yc�0׃��֮(\��/����Z ���ן�����tP����q��ʼPwk?1��S{��Ð���伻��^�7�����	b��ҋ����\穫pZ������f�����Ɍ�v�y������)a��Z�f$;/��EWn���T�T��p��ʽ�چݚN�����f���`�s���C<�JER�%=���<IR&l����w�
��G<b p�>�����K��T�V�}C����3���ܽ��S�I��Ýv�t�<[0�Vw��6+r���9����1z�ys׸��ܬs'u{�n���`�A{����5��'��X�.T�%���{3���s���������7qvwk8��Ub��{=[[m����t�$~�+o�Ks���}޾�]�ao`O%�O��+I�����s�� o��T>�pL�І//z��>��G޼��g��/�XG�'Э�nȣ��y��Sh|=�����}�bc9�����§OǷsg��W��ӽ���Spb��Dز�[��q�zz��{���5��USr,QiN���K{q'g^�x=���8��8�qt G4œ���I�^e��;/���EyJ;��0��\g�Y� ��e�q�ټ`ͭ�Ō܈���1)�ze>�}o2Y�=x3[�Ft�Ч{���|�f� xysjg�w�j��ӽG��ﰡ���T������Я\);_{s�>OS����:�92x�$�{|���W���#��S����,�nT(��յ�H��$!�s��$��C�ܻ�[,n&1�wZh�t5�Vo�b=;�?h|n/���X�=�L�JCK������~)��;�����Ň�q��ּ�w/8����ҟ] �TO�T�=3v6�&�8�Լ��(;5r��}�K�����q���<���'�q��H�^!��|��޺�Z&]Zc���{<��b3�d�]�u����'��Ѽ��3	]Яb����ه7p仓nO�4R�ǖ^��X����^���K�uRA�׎��fg`<��q(4J�%��n��h��w{=������]<[
�c/gc22�Б�����'a�S�B�<<����1�u��j����O�^�1�����w���r��B�{%M@<O��n����uJj��ϒ����	��w���6�W�`�^#l�E����]���YKv���$���;-�:[��|4�U��i�g�k���!�|�U�y���}�7��;gS��ӏZ��ۧMZ�o��(�gD���{8��V���аLZ�ׇ2v��P���Q	��%�מ>\�?s�_z�;u��/�Z%ب�t0�:��}to`!Iǈ�ǳ{�y����R�2z�W�u��S��ӄ!���%SJٞ������ʢ��|�q�x���?_�.�nrTzo�DSn�Y���cR=��;�P��ʼ�+�I�"��T+>�t�\�9���F{n��Y�w�>����FF���������2�fM��N���{޸7r/v{�L^����o��ucYq���VIa�t����񇔥��yz�9��O��a�_!���f�ұ�ߐTn��>vy�*Q�-����ǧQu�uT��{fP���^�qC�ո��__ �b,s�)GD���՝W��g7�:nǳ��030���ffg�߿���tFkn�unܠ�Rgk��lnz�\7o=]\�e{[�v�6s۳���]��R0n�;�=vpN0j�7'=�98��v���3��g[���Zh7piq���\�ݶL��y�q�KGc��p�f�)y���p]��[E@�nƇhAxz�]�m��x�FێT�T۴�d��[�ݴsն��{;nm�ɍ���[m�Vպ��S��-l'�%ag��]�h�L�]��s�ˋ���w9��X���v�Т��j1͖�����i���,r;���7^���wMm]�g�N� Ӵ�gq�<����{�� ّ�N={&ܜ�,�<��G���{���΅3ۮ�c�qІ�y؃s��[s%l;����j�z���7h�hsd���wtŻN��pt���P�;s����M����\nų���3�{�[S��؀0�#��6����m�n�v׵�Y���K��r���g��l�[��㫃��SϮL��>.�/����c�B��l��rҾ;Cj���r�j7=���X�v%̹�l,S���]����k,#�r�h�H��K�q������;�8�F��v�W��n�j�ۨ�r�gl�l�Lݹ���U���
z�Oj��� ٣���r���v��wAuX���Sm��<���nL����oOpks�w=�k�؇k.�bhڊ儻GM�A#�𹓬�]��ی�EƶmŊ6��/�a�s�B�V�9�h-s���:ф݄�@I�Nx�Gn݅캓�x��'INy�s�!��H-:�<�����aLpX���c�3���v�������v�l���[;K�w�l���V݃��bXB��i��u�[��H�FF�c��ܼ�*K;1&4�;�'U�Kg��.@Y���Q�=�m9����R����9c��úu��8�nќ��v��{�{F��ݓ�\z�]"�ۮ���9U��]�l�u�z����)q�-U���h�d�M�#[z��r��ɹ�+�
q��d9H2�OgO6��0���::��v�ϵ��3uӺ5ɐ���ywX�dC�U��z�x:y�U nm�*�����5�66ֶ�v�n"L��+�qth�L8C����cW���CG7^����3�Y���/&y���MX{	;ѨCF$���-���g��ݥޱ�x8����Ug�ڷ��κ�eKR������nCXN܄<���b�V�[����tSuEatRE��\��}�m�����'��Q�ƍv����z�[�tN��3����ó��΁|Bk]l��b���g�s�ַ��ٹ�܆��62�;�@T��Gnѓf�6���1���7�3�秴��=�˲�]lPK�t�.���0����<�����oW�iEvۉG�N�c�N����+�=V�4v�p�v�����7]ڃ�YGYǵ����ݼ�8��8�t�:8��=���Tsًr���x;Wm��y��8s]�Gs��;{�;/Zz��b���o`��j�ny�zΙ�v]��3Т�m���r�ڨ�=b�i]۴�]��q;��ɹ#t������K.�n�s�n�ֈk<����8p��Fݷ	�`춲�I�Z���踈ˌ+��V��q�Z4���l��ݫ�����LX�Z6u�[,�%�.���j<b͕�c�nz��䎳slı���ֶ�]8]�%�[�I�:�"��+b�۴����r��.ڒ�
��rB	z�.;[��r��ʝ��3�2�@�nw���K8=n.^եʛ�g��{d�{���C�k�٤�s��yl9G�\[	]2�},��zn.�&+[��PY�I�=�k��k���:�q�
m��ֳx�o3��nش�Wm,=ǂ�����+���˹�.cÍ�:��bw�y��n���ư�m�qƀ��
n��ك�r�����Sra���p��7Iɞ�2�w���t�>�;f�v��=���u++�i7Q��2�]����ql�p��<��ݹ��!�T��\�R.���v�5u��#\�R-cڪ��1�e�^{j�����:\�<u[�Tn����ǣme��1݇�1��0,)7Otءv���l4H],�A�[�<ꢓ1���t�5c�{<�݃���=BqF;��T�q�6�ɲ�=��Fp�l����W�;\V��}�������[����w+�t@/�Ƿ
l��8�ݟk��;;�n˶���m��庣R������r=v7/9�}��i�"d�F\��U����kW`$���V��i���*9ݕ��{v�n��)���[N$�q��F{��,�8�]��6z�5c��U���N��m���Hzh-6�xθ^{p��X���s�]6���p�"��n'�V�3ۗ���:.� �ɲ�p�7mֺ� ����\t���˗��i3��;o=�}6��q�=�n�m�v�kZN��"qs�\��>�ۓ�m����7f�˸zQm�<t�Փ�s=O4ny�˄iypm��wm��d��}�힊�x����U��,�ȢQ�]R�dr7EMɵH�;�,N�v��㗄i�W]ex�e�����pc�˶�9v�][�y���q��'������O�9	�V1)/Ic�ڞǎ�cC%��ᵹM���[Ǣ�bP���r۝8��и�u�8�����v���T
��[��ۢ�˼�JKf*��c�ܧ.�[���6:맪��s�������8�v��ٶ�'-�f��zlnK���(`�y�''G<g���6�'Dϊ�OVK�;��b��8���������Ѭ{Y�p[n����RJ>�G�=�*:����.�mnɺXN[�s�sfY���.^��|�v9��nݶ�5��=�A^[�y}�nx��vۑ���]v��9N���̅��ck'Ì][5�vNY:+�6�x�v���My^��^V��9ϖ��Nۜr�z�L9�<��wN|��n���Cvx�����5 mp��mwTq�W�C	n����ރ]��:��t�b���c��p�{[ɮ�|笘Ī\������@��]To�'[]A�����v��59��4�;�W<v::ч��\�re�OrԽWC����3��	�k�\����r:�l$��z���,aN��T�u���]���>�u���\�wF��u�-����5ۣj��Cm@th���0np��O"�t]b	��������u�I`�sQ�[��q�[�ob�t�s�Oo�	��&�Au��OIຝ���k'\��6#7�V��'<r�S��kEXi�qvz���]m�D�r�u�i�c�]q��8�ے�ۜWX��B��Y�'^�C�n;f��ݷf�Ӄs�80F�i��H��-k��n:�Pw�^;�n���a&n�d�^x�K`^���㜱V�'$�Eny�]O/<�s	n8x�����l[���׭����]�x��r�,�$��X�f���ԭ�L��W�R�&��]��vr]b��>�Ű���(�6�e���R��l�5�g.�=��v�E��Ŏ�tЯlv֚;vΆ��6d��X�㣝�Og���DWtvHl�����ȋ��K�mnH�G��im�� ���s���ۇ�vL�<E�
��%��lC�$���y6������ƼWn��N���i�gr��p��vK!S�!u��/V/6�$�����y�|���k�������s�� D�95��m���#��A\M�nps�&N��n#\[���7<Zq��s��O#�7�==a:�.7e����n֠$�s�k8-0�b�����;�:�r�={�SOJ� ����5!num��E,s��N�j�`xn��aSdǢ��k-��ے#m��>�=����ݸ�ۭ�Zq�Z�WVݓd��Af{\cs�v9�|�#ֳ6#��v7J���磉C<{2m�5ط��!ӹݱ������]�@�d9\
�<�:����4�k:�NcVn5!��$��g�\Glݺ,yk�^��=���s�-�����Ts`kA��ۍ\�m�5��s��W=�q	���U;�9^��=u��kC��C�����Fw]��]���<��Ŕ4���|س:�%l�-�ݮ۱!Ǯ���uOA��ۚt�7i7n攫��;v�\l�mt&J�1�\tR�i���k�k
[l�+6ҫ��79y/l�+!�7[�s��l�:�@l
����`��j,t� ��5�vN�r/�%�re�MlMu�S�.�u���J �N�u���u��4׵N���ǲO�]�瓱�1k�������i6�V� �&��1ȇ���ty]<�[��ڭG&m���}�۵�jA7Kdf2֚��G.�,#��6ݷnѭ�^�^*@.]ٹ	�;���V:\V�g������Vns��7�죷`�u5	��Gb"��f,�׬W>`��|�K�'��PQ��[5Z��f�8ӭv��66ۄ���r�B��>,1�<ؼ�VW/I��'gpbc6؎W�C�[�z��$���sv���h�:kݺ�tdJSY*�E	�n0��x�X_O9�jɞ��o;z��F�k'�ZFr�g뮸�wc'<yGP@�v�{�hΣ=�G��VL�Z���zv�ۛu�rs�n6-�m��Iv:�9s�ϣ���=�g�c���V�5�'n}v��5,��Bm�;vb+��c���������L���k'I
g̸�.;f��d8�<r㜸Ͳg78�s�/nު�������=uS��:y:x�g�3�Nΰ��!�qά'Z�M�iÓ�w��m�u���swsX�5Z:3i&jX$��g��j�C�#�V;]����-�M ��q깱���綳¼vU�!W�<C��w:麸�Rz펖�mZݎ���m�G����`�=Xn�n�RL�Y��N0\qN�`rn��LLm)��n^͓�\�]���[�ڎ&��Mx�=[ͱ��zu9�ansv崽����������D�UX�1pW�2$TU#�\qTF! �B3#X�A�	#"�"+��\�FEb�!� �RHE\��"I�1q�E\\H����QD�G"
�DaE��q���q!"c$�q�H�⊐qp����I�L���qc\Y(��*� ���&9$�!!	rc���"��!�q�d28(�����($$UZ�Ak�&8"(�`�ɐY&I	"�b�+i##
�	2���."��I&"
���")��c�
dEqQ�H��10TQQU� ��&D�2J�U(�����#�I$�$dpQU��$QGGRI�HH�3q\�I$UQqD�H�.Fb��I"���AD"A#"��đ��,��A$��
"$�Q"F@�b*��BIbF �EV8�`�Y�A�DGDE�GdȪ��*2AT\ddSd&	�(����A!2�dH�fDqB*
FHGTX�1AH��*��+�
�����#1�1Bc#��q�Y �3��������*��8�U����5���k�a�m�=�
G�3��G��u�XM��L��ۋ��E��Q�\���n6˭�f��A�����ؘY8_]b-&[�
����9�.;uzxK:��iTK���=Bn<���X��։���t;��u:���c���v�Fݔ+;�����(=�8��ɻ9����>�l9�]Au�Ns�0��=�OW���ku����rnv�=�8^�twWgZ!�"�WL� pyS�'���<<�j�<��n{R6��L�|�8$��Lw��=���;Z��g8�%2.㱷cۙ�G=������6X��`踟J���y�!�*E�m����㛂�x��<ulk�t��R����r���#�,Kk)wi4�Tm��"�R%}W.�t�b��k�֞x3�9������`�̺�vN�c^�6����Lvwm���=4�X"��k@޺������8#�,m�<gF���u��9��a��	�Ȕimlj�j�,�b�5$��jzI�q����//Wa,n�tnu���vé�V��]�����6��I{x�g�+�=�N�9��ɷg�q�λ�=�����j���P=uاpA�������s���Eخ*�9;��Wl�bM�/n�Kx�.�]nm��z�;v�y.e����s`,;�ۢ�T�� l����-�w���@�=�ezvۈ��2nQn��i�z�y�]������u\�[�������m�)-�� �<�GGX�p��$�o5/\�R��8q��]��g���K��]�qx[S��r�u���-���t�q\�[��F{���vsnz��v��-��@�.$�y��E�W��JM�5�%�Y1!77j�@�eE�[�[p���o����9�\$�n.d��ݦ�l=j���3��m���'C�Q������\�;<�^��纺�_>�K��=�n�ح�������c��7D�-�ɞ=�9n��&ffRYd����-n[(U�e�[nBIJ[J����U�(��YQ����h���l��J%���b�F��FLX��2$H��6��+l�M�i%�X��F�l���Y
�N8ݝ��8�`x2dG�a(�[Y��2��c�K�V1��V�)2���"�U�� �D��b(�IRH���,��V�#
�6J-F���jX;�$&��n\�Y9nP +�zJ#��o_�Sf����ߛ�0��������)M5�J6c��WM�z�-y�TuR� g��% |ftp�؈�ү}Gy��2�j��=M���#���V�]D���Ѳ���;밮���J�y�_(K3g�_E=��Nd_Ď�սn.��νw|�)2j$}{ωe�M�U�uKo)įt�� �MdH$jɉn�8P��ҍ���� ���J��'<��7}]T�g��� ���|pg���͹�V0Z~�/���F���y:<!�v��Л�W�+���v�׬�l>��fe�aM�q�H�,�n S��Wt����J@�/��^ʳk<��m��gtH!V�l�U(�����!���{/��g�xRw�]��+��<���=ʕ�2`G}���~�������}a�z�o�5A��)͡��"��O{�	���B+%���!�y �|I��טxO�O+/����7�|��i��{q��|n^�%B9č�w���'�L`����v~������S�r���w;�|�&���z��$}�y�_ -�vDfN�:]�O�{�Qݮ���Jߊ;�����c�>WdHn'�wYޛ�u�L$o\i) }�ٕHG�����&��q�3�R�+���8�fB�sɝݸ�6�2s�mu��W����I��j��n�8��q�qR��E��J���;�ə�ǵ>B2�2j����$J�L� )�
��(�^�4�k��yï
�̪�}ޮȐE�B��z���t(ʉ�	��)��R=��J��"@٨p��U*�߷8��<�ݲ�b�!��,6�����Ó�Nk'�+�;����~��W�������_�ں���;.n�����{���s��s��7��W��J�k���C��6Y2�8.�=����=�wG�\�f�ܐ�]IP����gG:��ݴ��s�0��گ�*�;�؛M2>�$�t��>ݮ�J:��˚�$��1�G�B���7vMY:#�[��9#A�<�'d�v{����w� �t��)b���G���qjG�y�Dy�8��ɯ�
�q� Ef�/"q���UuYJ�"���r��n?48�x~��މ����Hg=�ܼͪ �ƥ�gGO�񱖝s�F�Gw|	L���~��=�*���r	F��J�d'���O<����)@�͎�J<�^�����H̾[n��߷&c�{�VM9@,����VU�YQ�h�&���?�ҫ��ĥql�~o����^%�gD�L����)�R=��^F����p�p;��7����������t?D4��C�������nU�*�5�D���"]��})����a��Oɺ?6���A����c�Gǯ��V��VU�X]ܬŖ@ѹ��g���h��8�v�r]ѳ���={t�|�$js�9�@�܎��7��#�<�Ď�o�~<���zŕ����| ���������A�wi�~y�m��wQ8�d>��C'3L�Y�U���;+�$NM^����~ۋ� GwF��B
�����~��x"i/z{b��kGnl�����^ ��ʤ���%Ы,�KВ+�� ^�C�R3��+�{;���r�ɨ\��U>����0��$�>��ʯ�z{"Q]~��~����~s��8N�l^�i�8�~}����L�Z*7r�Mp����zygL�vh�of��w�+~�
�"܋�6I�R&lMB�ĹE/c'n�y#��[#[�nۚ��K<p��r�\�p%s�9�ItV{Y�G���'^�/�j��*�8�n�m�öC;�v�l��<˭R�v�JB�"���Q+vAM�]���������r!���ݣsq7sՁ�k&�6�{���0���a6�vL�X;:\q����v�,A2Wb��U�s)�ۭ�ظ�����Ύf���[�틑�8Y����뺳�Sqv��s�d{Y�������8.�m\�A��n\Z�J��]��Ys�B��ؼ�t���}[z�pᩉN[�1��_"�r��ˍ¦�I ��ڤ�{"~u;�*��̪S�c�xO'�!���6(!���on�>Ȕ ��ǟdu�^����]�@�h�&�l<��D���&Cޖze+��E	�Υ@ ���"P /::<�7��_��]mR�����0�E�@�+�1o̀X��r� ���>ȿ=���j����&��b8�����aW��O]�;V�csr�YB���JD����`��H΄eo\Z�=Ƥ>�9�%ZfC�?E��Rs�r�9�Y�q5��Q�Q��5?����'N�W��t��Vģ�=���k����5��wv*�r��S�Yr �S+����n�PQ*Dd�������鋽��G<�"y���"^��#f�t��^�6���S��K�۔6�6W���ʻƺ�đ�r�*��<�)ftp���7���8m�ߵ���~^�=�-1p�Y.P/���Ă
�ή�'k�]���|.˷ Z{-ǏC�!��õ�>.�:�[�ɏ<��Z�$�Ee��>Vll��n��7��G�e���l��;�$�@���F{���Ǥk��6��!n���n�1�9@K�߿�:�7�/(�G�5����O�
�����ˈ�u�w텑h�r�6�8����QԀ�X��u��L���f�x���m��P|U�J�-�gD��d�c��s���� p5��n��:R������v6SZ=Q瑔9��?OL��¸�C3������aTKO�Ԯ*]y]­ǳY�[W��n�6�5�yz�N�wV�P�Iu;����ve��!wti���Ϊ@�ګ�ؼ�
����Z���<�^�|]tT��%�Y�_�ǚzUe������^>��X����N<��G^����5�f=��oI�u9>�u[�A��9�Ș��u��Q����M��L�$��v��6��y笕���Y���ؽ16�������L#��B<?rFWDϐ�uY��@����ELEr�[bwE���J�mVm*��l��߅�H����.��gr��w�U��^u;�@>�(;ݘ�߈�wtU���מ�� �~E�����㟀>1��X�Z�-l�l����Ҥ.}�A�r�C���ח��P�:����ov�m����o1��n�RȆ�vO�M=�+K��ƭmM��t�a>���
�b��xs�!m �}���L2$�5vM(s/&J�L��@�nQ5$7�z\��G����f��b��qq�B��kr%�A񽑳��lFgA�(�� 1�?��7c�/2�_V����7��^O�58�v��ΐ�̘���q�׍J��jv.�m��mn-D5CN<��G^��·�Ԁf��P�c����U�z���BK��7"$`9�L�[ޚ��Rz2/}��O] �o����펕�
TTM����߻o�J)�.�2K"e�AT�Ok�@�͎�}���2��"�7�jo�=�!�|f�q*��;p8�Ny�R=s�*ʋ����/`9b�HY}nP vc�DUNuw=� E�M
�u��yw��A���74��c�/ mM�V)��'0��Χ? �>@%U7�x#������B����������'݅.��x(e�@����7����{��}1~�n�S�K���j6��2�9�����J�3��8�f�A��}���	%�u�E���@페���F㲋뺎��r����&��6����<��?�����+dc��`�6���<�\���md*����]��q-�vy�.6�۠�!	a�$ʌ5�W)6�L�lڷ7Z���{ma����v��[u؟V�v^t���=k'e�ɉ�'�s���ѹ=���۫��v�l�l�.w<��v�g�Ǣ�gn�o����m�۫�H -��<&�.�ۤp�@1�p�xr�3~���W��B@n�l��*�:i���-aWo�[��;.P$,̎��jyr!�^M�CUH�ۺ��qv�_^�{Km�ρ -�|O��UYҩ""k(���~w���A�Ss2��]}4�%��J6�^9=��➙��n�J�����)}KeL�șlBSv��|�yC^��.���� WU}T s�rgV������r`婎��3uH:��νJ�.{�I��qw�UO��ϧ&8� ��oj����XFP��{�K���`�in�����M��jm)�b�<�<0��|���b�=��8�3 ����w�e�*J_���l�96b�v&wf�/�Ltl�!Y�WP`6��Զ澅���B;��z�%����_ΫF�}�=烯��t��x����=.^j�����ݳ�t9hu�wp�9�+r�t��"�匬�PNW�}�Qs���r�ue�W����T{.j�v�Iz�oc7�T��CP�����j��n��*+�� 1�M]��ދ0>�w�_ =�@��[�	���2�m�םMVu+~�����]}BޜȔ!�[�[���+n�����z"!�!��x���+޸��#۽؁}�UUHB�V�J^lt��Sg�����,��n~�r"��c�����;+`6A�<�0m:�ڷ�.!�A�`����%���Ne(����˵	|i[���>%��:��zv=KӞ�yW�<]������I���{7ܿR>7U3M�|yc�o����Y�?�͎���9�yr�ܻ���;ӈ�2q+���Ao�ey���/r/[���N�=wfU�	�X�3��G�y`��i�3�J�'!�4Wզ*�l��m��O7���~��{������l34�追��(���9ky�ا�4��j���bŇ�"�}�����S�v���&]�;d��;�o}�o�J�;����\��r�|�;���W7�nK�}B;5�%�ćf����y���r�;Z��n�^�W�*����]z]d���T��A೽������{��P������7g��f�<��ry|{d�������B
�<�p�}tyW���T���{%-�ݞ(7Q�z�2�Xwz`���7��r?w��7e�c{�f�<~ƌJz��w��Fkɏ�"u7�2�Z���[�];�d�Y[*V@��������{vs�!ǳ�Oo"uEÇ%���2MH�����	c8C�]:��á����q�I�6��#�Z��rk�o�h�����k�t%.2��ܷ���7PQ���x�e��I�uNm���#i�7�/�Fn�z�^Ÿiک��F9݋O_i������[B������7������_bpQ���䛕m�}���sʙ�_�Cz�}������7����N��!���ox(�1��������,�Į!��e*ݯ���{�so(BH�㶝���! ]P>�ç��F��=P��Q튅N��QH�-+"{ǮO�g�����E�s�&�E6��k�e�v���ʖ}R;�N�����U����=�����P�K�)�����؆o�zM�qn�>���#z�!;��}�^�a�󤯴�߻���-N�iFI*�r��1{���=�!q*�EpE�I���HG�"#�EB(�Ec�EQ�+\d����*��$��H��D\EqUL�"�" �8�+&)&Gp\RH�����8����"8����!c��Q\DY"�� ��ȰTUQ�EDU�1c��QE��GDP�(��"ɐq��8(Fc�8(���"��Y(�D" ��DQA�QWULU#AT�F"�
������⸤$�EUEQX�qTQ1U�p�	����T�IL\#qRL��$q"@DQ1A�
9�,H��**������ 䄃�"$b�*��)� AQ1U�\d$��EQDX��$I �pLU��$Ȋc� ��X�$Y&*㈸�ET\*��8**��#����
0b(�(
�����ⱎIb̒aEW1UQY�1TQ$��(G&$�RHET1U�sQEd �& ����{���k{� �ӹ�������&C>��F�m�ܫB�Ⱥ��R��R	U��R	UVuzwQ�m�ގ�٫�W�Q὚�Id7��	���2:��@]VuT���2�UQ>Aގ��;PB����ױ���١=�NCg��c&�N���[�7��;'<֎���n}g�轝�ff��I3-�2���4�%
�c�������W��+�+�gLO�}=BWI?(c�2��#*���y��.l�'f) ��z)AU]�H/F/r�b�<ݠNz�zDy��x�n��H|mV�P��r���c���[��H�::R��Uv���<�8�!��%�,���t6M�T��+��U�U� �����J;�w&Ɵ�q�{�
Vd�������;��@c��&j��B�:#]xc��[���{+�"���^��j�M�R�ҔXe*\�u���Np�x~O�G����R�
��#���&^`�T��K*��Rb�+6y�/=��o]��ݑ���56���T��W(5� SO�Z�llAwϾ��?mȭ��h�Hڸ�O��gR���?�ϳ�ܧ�y>���w����QIj�-�>^��c�����ҪG��>��11��
��j�|/oc��
�2�%l=�EJS�p9�#7�z���ID��P��l��J�:٩�U7�B��?
"�:0�3#��&[�U[=ѝ}�/lδі�)*>���!v�w�۹�ڈ!r��v�aO��i�y�I|����F��Bw;s<�e���ҩ%;����=D�&��V�#�m�C��Kq:?L7�H
��c7Ց�N�td���o�0��o��tv9^�=8G���S[&��~�I�����w���1.r{�������w�ﭪ~$�HJ�u�G6V�Y��k7d$	��-�3����z�۪���n9\Wl�t�ܦ�ĳ�d��o]s`xC��ls��]��F����
��ڤ-���{q���q��*'��m��:vN��Þ���x��n��CKh�;Y��T于0'�n�ڭn^wGF��c��k*lu�g��X��EN�xX�Ѯ��;{\,^�ˮ��S˲y&�u��\�9M����톢M�߿_�߻f䃯G�kU�~J�}oq� �|J&-V�w����뜪���joщDG�q
<?JF����[x�T���*��c� ���^A�S�zr�}/r��ݹn�!/}���4�Q���נV�[����=�� F<� ��;c�/4��1��Bd���[;���|�!����y� ����9!�M�=��A�8�~�։!�̷X��z�!Bۯm}Y�WN:�/�H��rȫ��^G�7�l��헗9gr��T
fR:W�G����vs��p>[F�(����;�ό|����46�G���~�ӟ�ݑ��$!UNuR/���P�j�1W�R ������}�)q#���]���Tg*KŞ�/=3p�5����Y� �Z����:�B���~ZϹ�K)�^���I�"�8��G�/v�����h��X���۵���&�h��%�6y�@ �?>$����:�d.��=ߪ�� ��U�Iy�������g� ]Nu*���~����R�]�!�>B
�Ϊ��/T,�e���>Ev���)��>��;���U7�H ��� �Wq�yG�S���#�'�09#+�z��"�$���9Ez��:��Nה��:���9�i}
9�:�q99�����}F�p !Ca*8��n��fC���h6w]͗p���$��l��75��hR��L�~��}�(Im׶���铓���>;��y�7�I������n=(�t��>�tpOD琂�s*���9@��vLW�q�%����jy	��T�v�o��@����O�*�.vxN=�F��{�����Q�����m���0(&^��^��gc�s���]�|���D�?w��8��հ�����M�����k��坓���S�f����s��P��^��ڈ��z�I{쎹��/+��	[�jP#;c�����CW
=��[��D�5R"�Ƽ�4z{\��+�N���U�z/zi ��9�>�힨%���u�yQ�$�Dı���W�5��#j�Ѻδd���&�WM��F�kMnز���T1��d��eoU���:K�;_*QE�v��	f�uP9�9�9{��
?!�M�q����܋�}ӛ�R[�r3�:|���EW�ɋHs��
�q�`�n<	���n:r���~�3��^��6n�9�9A�v:W�����y�M�^b�F��Ԓ����z2nN�9@�����1����!�����W۩Ѡ�<eo��z��ݗ�1'��v�}������ϵ�Q=�_�'5�w�_�yoDMR�?\�M�{�amB?/�_(��|m�9�g���Pڈ�_�ey���T]��^���!��@�)�>m���&�f��k7x��n�5DG-[:��m�<ES��4k��g�V�[�flr�an��_[W"!�Ak�{���Wlt�@UVt������n:-��E9�? �#�}�0>`�;�Q'4����?��E:z�j��l�C�ԂA�v�% UVuP|m�tΛ�b����|�^�xM����D�G�^�}��x|��u�=#�#��HUgU��M6��m������TU�=���GE�AmWeR���$��]\�� y~]�?KGp��ıR�ٹ�W�Pc=��,�n������r����D_f���kU՗�ӿRRv�z_��޻s�gI�rd�����k�%����x?���eu��l�~�/�x�{�jᏡ��g�]�yz��3�̧��֍�7]���9<"8Ӈ�<kn4P3�7M�l!�� ݢ��:G-ʻ<��z�ܼ���	�I����y�8s��zyL�t+z����W=-ǪI$�lغ�-G��#a)�bŭ{i���yG��6{I[�ĕ�����cAx�&�F��u�d�t���f
�0�6-�n	nH�/[���=���-�SўS����/�������ɺ!�V[�i{krm�z�v�����V�3�ã�lQ�3�X۵\�}�n����ͦڈ���ؒP"�k� �|���=�˕��2��uV�P)�9R=	�C�!�<A�tt�y>�>�.c�3j���� ��ꯀ>F��K�^�x����z��K+�8!�e��\���B�jA�̜������eel� ��s�'8r���n��n�=�4��O>�v����r���]9�Oį$P��ϳn�(��8Ci̎[�;�Oо��u=�Ϯ:&�Z���#�1� Fns�q\n�O�M���W�k�+sc7jM�KG&�6Ʃ��vN;�����������v�>����0�^�vkx���Rq��nt�H��O|��s�;�wTW�P��k��m��@�&�˔�
��Y�^��-�u}�.]�����j��ז�k�.��E��\�n��[�w[=KJ�n�z��ս!^��r��^��uW��yj���K�nnz |~���� �����g���ǧ7rV)�5R=	�C�:�z{\�@���( ���¬�d�MP��q�n�H�??5�?dD8E��������f�	�1�@�3:T�*�zr}��mWK}=�HoZ��]�26�~m҇���>6�v�����ʛ��`�������U��Q��y;佋�E���08Q2򢓢DEOe���u;J�'��m���>[�`"������Dy�	�q��FS���π�]�U|j��[ʓ��FWS������_a���7����R٬�O.\��.UT��] H�|JWs�_ B�}趗fFdֺ�=�"qy�d5���.~��/�˞�i9�Y��H����c:�vۯhg�Q
F�_D�Ͷ�wq_�Y���{�[��.f�94��i����d�-~��sNnt������>�3�3[�~���=Q%~�~�Jb�	�-�I�|{�\F�ޝ~�ֶ*{Դ��:T��ռ��{��l���Ϥ����N��Ys��^�י%�����X��&����Dq꼀]Q����.��Jn<�z���D�������aBm�;���G	�6�kS�tF�������Y��Q�d��~�}֣i��J�?@�w��|k�rrٌi�{�wfh�\�U?/���ں��D�3#�Cm��˱ۨJ!v帣/E&*ս��z�HB�y�H����_�!�~�,����߁ӚCx?KcT ��9˺��5��1 m>ꯄ�������C^��i�L��{�^׻��ځN�}�P 0��w��}J��+�mQr;�ջ8nk�L˽P7H��יK5޸"�uo@|�����|R��羃�5��"��莌;����>_/�I5��S�]�b��?�Sd-61��~�
���=�Y�~�W��|
�v��5�9@�w�jTe�ws�U�`�C�p�ɸ�7�c�0Ȼ��mc��:��[��1ʨ>�5��>���8k��"!�#�7Ԩ���ԡ�މ�*���Tr��Wy�uU_Gc����3��"1�n�Չ��S�F�/eN��G��w�r% @�7z~hD'fL��ae~ɳ�������3V$���q���%i������d=��� �<Ȑ@�3�S�a^�~�4-��vKTx���%����P�(�gl)����]J�u~�/|�Q(=�#d��6�k�?JG�~`��:���;k)�f�؟�"�$ ��t��UgU���?V.���u�^i��/�g����͉If%�㚼�|�43_���6���:�W��;�[Po�w2�cOC���q�N ���/�YH��ח�ΛxM���F��K���w��������ѣ�����9�@L��xU.F�������z��qKb�z��R�T��2�J�u�/�d��B�Ġ�u������zw���z�5U���̎�m��kت�R�{��3��+ӷ|�t�:h���m��u���_Y��z�=�v��`跴z��CHa3~��v�{&RpQ{<e���~���͸��k̕Y������������z-�N��ݾMH��jץe����;�fz���gn�>�2�݂�V��E�h�<w��~��|���!�&Z��~8n3����#s��m��\^3f�TPz�2k�Ą����T.)=��Tcn�/p���ܚ�؉���z����˧��U��n�[��Ė�ji�m,�:�n.C�y�+��MZ�W���bRYF�:Q&����/C�p�Iݕ��W/}�� Z GC^ٗ�ѽ�ݎ�����D坻�5��{��?!?x�;/T�߶�۝ݱ�u���87�֭����5{�Jh;�Ga��ڪܶ o���������(â���ӻ�v#,a{2g/:9`��y���D[�p,�{�^K 7ׯ�!p����A~O:�I;�w5c��3�	Uy���o��.���|9d&�y/8����2N��΃M�G��ɱe��.����K��]!��]�'��\���Sw}���ߜDd��I�*."�X�2H"�8����\I2b���"
�DpWbF3q����$b�☡"�Tq")�L�&b�����&HEDē"�*� ��a\QDQUBL�8��"`�.#$Q��$��Qqc1��"�q#$�$\EV+�*�b8"��ɑ�`�"�⊉��	�Y ,�H#�r	c̐D�H�Y�F*�0��Q$�d�&BEa
��c1F1QT\�\Rb#&U�U�S�"�
,b*�8��L\qVL������b�&�W#RI�#�b��@Q�H8��AQ\DXL��+
�a�8����"���FDH�EA�H�8⃎"�I"FI��d ��2d�qqUDQ�B8"(�dDUU�9�TQ�FL����pE�GqTE@DX�$�f
(�"	��"*����������FDEV$Y&=u�����$�@��8/[�ռ �t��7��]�.��gƞ��h��G0�kP�q�n:�L�\ˬZ����`n��u��W0;&�l+=��m�]ٰ
:,,�6g�F��t<�F{1�v�P�8XY�̰vמ�D���wco�3UAs�s�v{��Zܘ|ܵ�cF��e��ayt�ױ��3c�L&9	7[�(sz���ݻ:p��k�v�����O��8��s�'�.�n������盍�}#f�����)���F�ZSN�v̐Wt�OV\(�*e����.�w�;�ַ0˖9n��b]ht��C��.�t�\�g=��5�ۃ=3=ۓk�S�7k��=m ��e$h�]7^�O���G#q�N�*�|I��G����z�ݎ�ޤ^\v���i����u��g�8_5'\ݒ�n�۬�)�5��T=S�ώ�qʚв�������إR�����T��s$C�롹��{���-�v����L�&1"q��ڛu�ƭ�]Q�d�����p<��ݞy���E�v�8�b{�<�.���'^�8���]�7.Ի��M&��˰����f�͊�K�@�Wp�B��ۮ."N�2�z���\g�ڶ z
�cn������;x�������B��ڞ�Ǖ7i�;�yy�,��8Up�|�0�f˥�nui㴺��kÎ[�v����l:h6�8��c%��ȉ�{t��!+^C��vK�Cy�wF������m;���)��1d@�-�Yۭ�.ᵋEm�e4�̫\���k7[�8ˋ���ݎ5�ZY:���t�Q��n�Yǯ@��:6k� �z��ycsV��7����K<s1.��nʽ��V^׌��f�taw'A���m�A�q���l���]痵�cm�f9,��^���޲U<���\[&ɺ��8�׮Wn9�W�^W�e����mɷ(�=��3{n\q7��IM��C��1͕k�nǇ�V�J�h�utݣj�a��^���x���k��;��w#���GED�n�T��m�6��ţz��nuJ�v�,�q�)����9+�GcuX�v�mvֹ-v��=�i�ț�s����p3lG3��y�n��Z�'��X����ܝ\���n�ص����K����[���K\S�����:w���m\Ç�f���ۑmwd�Ӳq��kb#���O����<=rkN1ʳ�����x�:�7�ԡ��J��2��nMn��^��%�	�Sۼ/�"f���WtH�^���AUVuW�/U�Psw/���(����AQ陸�ۤ��[nކs��绶������f8���J
������W]u}�����X�W+��B�8m�|>�\������H��Sz=�"�+::W�T���Yz��=�Cm��2�ǭc�R�)$��j��%�}���Y!U�׾��f�O�{>ݷ+	iw�t�%���lx��W
|<��'L���ݐS���#�u�T�&�O=#�0�ʉ����M�0��n��nݱ����vҗq�!�*	NC9`����T,�l���#b���u�T$>�t՜�;Q�[����[_�p���x7g�-��B~������FT�U�Q��>!,b��5/tAg��)��_��o��sNc�YʺG��OM��˺{�wiݩd۝��fJ9�_e˓{���s��rӷ�0�0�����U=����=�u�IB����ŸG?t�G�O�K��ă^dD8�y�uP�㍬�����w���(�GO�V�i o��%�T�S�
ۥ��6��7����?T|�'�Ww��o&)%}�ӗ�]3M�ft`P֠yyԪ��Y����4	�qލ���΍<�U�M�Z��O]P�udJ>���-�d}:�I����-��8���q�^�[c���px^����=5�i$ݱ�����̰??���{���Y_P�"ͬ� 
��R�.��q��]�Eo+��T��K=9�(>���S� �!�@�(��r}��Ʈ���^�U�Ѐ;���!V�9{k�T�e��gz�
��L�3;��>ؐ��Q�ݪ9c��jy��X{�[G#�-�Ú��N�C:ٽ#)�{��k�80��{��i�n��/;�3��^yυP�w��u�w���B���pԸ�12e��oeC*-�I	 �ؐH��Rc����Wx���r�ۅV��=Ǜ¯lo��W��^�C�W��>����X�*�&�.�WsP��.����a�a0���m�Snpu�X�]�j�x��k�����Q�x��?7��9�B�֥ AX�*�4EiOv�\�]�ۉG�{�M�N�ZF��-���-�yO=��0�aH|U�(V>ʠ2|���=�^�����P�(r�m6�L�6��^��v|.�qY7�sb��vs�#�}�A]���F3�:�}�{~�ۏw������s� *��T��WdG��B���]�����%�q�$��)��۷'���w5Z{��vo�%��0>�Q�:�7����g,��S��ѷq\���/�J�5�9@{�������/k��HG�"~�o�]̕�5h��(��4�Wd'��z����Q����;z��G.̼l^��pD�YՎ�t<�Auۍ���d�����xm�R�l��7��p#q�U7���^�\�5Y�=�5����יw	_��R�H�P����Y��r1O{���Oki��*��*�}]� �X��}ўЈ~�ânZ��V���%�Eb�����_/+오�OZ�*QWu�e�� J�)P.�vD�{|#��M���?J3���g[��O<������"A[��!��S��j���ۗ�G�ID��P�)ݘġ{���U뵒���=�T ���U߽��Z+��Zy�&~g'�M���Vw��^�&��4��I�M��I�*p��k�7�c��Z�S�h�?4.���u�ڝ"V�N��_%�F�H���/&nv�p/���T��Sv��f��b��׮�#ݖ���94v]'5�ۍ��붷g{��.�d{<�&s�{Y9ϲ��L<Y �5닗�'r�Rkd�֕S����.Ck	����yv��;F;��u53"sy�&8t�:�v�z���;y�t{�kq=�޺N��ng�,z=�3���"]�b�GR��:���V"i)4&�[�ۏ�ѻ�c���.x-�c������)�h͢V��� h!�e�������G�����#���@���D��$	V�ʐ�{2�XGoW7��o�r'�Np�ɸ2�H��>���0�)՝}�B	�oF�O^Nz�7Q٪��,���0h�G­Y3 �l�s=�YSY�]n/-��D� �[ѳ�w�Y�?�Ch�R5�d��V�e
���Ws�H*휮����wo�s>�/b�䃞M$t��P�&����?x��O�}~��rv�辛�K~[�y̎��Q۔������������6�e+r�������UT�k��|��mrS���[����������:���� ���PGnW�&�Y���z�������A��;ԛXM6ۻI{w"���{I��<{c	�:;fH����.i����,����TK�TN���Gޯ�P�����j'�ӥOV.�{����f��}��/�Q������|J@	T~ܪ@��κ�+��&������'5�17!8�C�s��������7���q��7cg�@�;r�2��D�$M��M�Qc����j�S{;��EO�ѻ��]��~Fe��u�C����_b�"����"�c��@>ȟ��-�Ǖ,.��KݏI ��ʤ	}��Us��:o����2f$C<��<ݶ��GZCa�,�tY�����α�j�������jll��dl\�� .7rU|�dp�֎�]�\���p ��[�>+�ĊZ	Bq)��>يD��s��5M�gN���*32��	��)��M�zff�r�2�P9D̷5
_n��=� �!�t{�l��I�C���Ѵ�잸.���+NI����xnOA2���^��>B��~�ϫ3�{j����j*���|��%{_����?nM ���9����<2<�>��s�Opۍ��u�uB����>+��jqU:|�$n�٠��dG���	��.�n������z�Z�e��w�S���V��c������w�ݏ���YW7i�7�p4�m��`�d���:�B�eB��V�w���n�c�n����l�RT[�r 	V�w��x��E�nѝ�]	%�c�H65&i�$i���x?�Rn�v��Z�w�0����򟇓su��-�5'ڋ���)N�!��P���wT�uޓ:fk��/y �o1�V��)��Q�3-�)}��}q�o�Yݗ�B��jAtn�J*;rW������3�L����YT���>j6�b�������SD�Z�kx��{坓P9�
g4Y~T���-�������+�
n����{�H�H��R;�3�TH��cw*��J��α� Fw�e,_�y}��?��[��,D8
��F�5���|����h��v�P�I�o<���v�䵺\0h=���"�k���<�������E�U"�Q��^GD�S�#;ݳ��dC����h��k+*�>��G���*�S��
�f�P|o���@�9�g��3,N�<vx��^jli�C%#{Φ���4*�5q�Jz��j:��_�eB>
��T��ԣ�3ġ�S�C�oZ�dz��Q�vT��5��Wc�{Ϯ!�4�Tz�T�6Y� ��D7GOm*���W���+	�f��{�3�V�*�.��(ʽ�7TEYّ����OJ�p����Œ-��5v��gC5eC���w��c��s4�X�ws�^���B��T�d�?����w߂��v�M���ٻ��Ƚ��j(��vٯke�T���=�91�Ϋ���tw�s���{���v��ױ�lpc�۲θj��cVcq���.��ѭ�ʴs�7ϖ絜<u���q��^`PA7gna.˱�tg=�gx�^%�c��񱔺{b�4�ʧ��y.t�6+��w7����`t�n�pW�c+�Ny4�U�gr�q�v��9���۪a�G�l�ݴ�/<�`����	͎7̽�������n���_ď?v���f�U�@��ƹĿV^�os�{�R���R��&#�G�τ�]��%��)����v_�A���ǻ+.�IF�c�P�8.�_��_v�5�'�,�~#��k�4��9��@�u�Ԁ�oEp���E�={Q���ӕ�|u�:�-�C���pȖ�b�~�ګ���34��|���J��>.���@Qݵ]��D+�u�i{[sI���=�g���R<�\�"��;���_z��/�>=ξbH��v��D����=��9J��$Gv]-ݱ�`�)�r<�k^��v0۶��W��ɟg���ߟ��}�X˞.���>��� >�Z{]0 ���v}YS��f�E�v��� {]0����0,�N��C�~y�����D_������]���tCZ�`U���)��|{���叏�{M��'m�������d�6�og��}ڗ�\^ozj��� fo������Y�?r���HI	���w������٫-�Mzu-�c^�ț_(m�7�4�@�۷��	9�U5d{����7;� |��_D����i�׮���k�^/tNdc3z����A�8*vj$>Wv�J�ʿuO��\>+����||�k��Ni���)��D�/����H�:�im� _?b�+n���:|�J� �׳n�@d�d����d���F�n �r��<�one�=��	���Yؔ�s��u�@Ԉ%)��GJD�$H�Jft;=5 @ygu�$��Փv���ݳE+K�95 -n��A1���&T�Ù����f�Kn�VG$�fL(��lH�7z�� FK�J�[ܚ�ʹ٪�Һi��9�"e����@��&���ܛ� +���V.����̂��UrC�&2��n���A(o�vl;�NJ����~�^��=�8�8�7�UpAJ��^E��Tas�1f�S��mےac�k��/=���_�}��d=;��TZ��j���q<\����#}��e�s�xx��74��^���wt��l�z��w���y1��+�����[���0�L�(�?,����tP�Tbi��;=����ԥ���!�0}��xz�Ry�۾�y&��N����2y�ƌ����4��c��%y:�r�J򯍷{�|j��˪|�i���.�
���w�~�I.c7u�-�H.6_*���MA��~P�^G��������=�����_D83� )�P3�/x^��b�[鳯�x=�Вʣ^�xvņ/p�컌Q�PD�����<�U����D-gЦ�xͺG�r�����R1�w86�ͼΩ�ghH���������}��^��m��.����ު�Ʈ!�d2c�ρ�`�9}���g�=6�����.��s"�zM�*� ����۽w�@n�:ny����ژ�sŖ՘p��fI���%�8\�0�'�r��:��s��O�-��R����v�|p[N�LX=wv���p�������3ܸ���j�80��q{�E�d�Ә����h�[[Ŋ��\�ӎ��F��ۦ{���Uǲ�I�7ޞ�s�ܡ{�{��-d�[���sw�^��^'
����<zX�7os�|��S����<��q�g�H>>U���Os�y�;�-�Μ��y��J��k2�� �1�����*��*�dQp��0X�DR�E�*�8
���8�Q���ԃ�"�Ԙ���DS⸊#��b�*�ciPQpEG,����*�A#����(���DQQQX�$.I"�1ȢF`���!�#&\UX9L#�*F�dŎ@I (�FL���\d�� �d�#8(�"�,[p���WDQ"Er�q�D �5���dŊ�$	���B"�qd�A��UĐ�H2̉$r1"ɑH
���\d��
4Q��Us�$ad�I"��b"�$"
(�ɐAEU�B"������,�������0�m ���+�$�ȋ�""��EV*2b�
�"IUH0QT2FLU$�#�FL��$P\UF�h��H�!>�� ;�so�����pđ�d��7`{��#��sa�S�)0��[����e��$}��&ҿ�=ν����.�m-I?���w>�!dd��C���f�^Mń ǹ�1�^mz������>��M�`|v:�C��Ulf3��M�G�Ͳ�m�M]��8n<��,����qgX6���rY\Jc41v�(��MD�: ;
�ų� 0{�qa  t�9K�1�\��磌~+�u�C }��&��"&wQr�-I8�vv�bR��sMB�Q�&�L��-���2i+ 4�r�@+�sE�]����Dv�rDʑ8s2ۭ��n��|@.7|� 	�/j�[5�ʼ�� ���7q @�c�a��݂%�_LL4n�����ܾÊ
=�ou� q{�qa |A��� /�z�:.�|y���{�m�c���l������F�9/��|=n�9s����p���}���7qh���9�?"���vڬܢ*ﴺʄ��$��}��۳ie��06�P�8:t� ��;qs�TK���g>~�&o=7`|��1�T�=w)���w�T8t�翽������Kl�u���kX�+������Ҁx�����κM�����;����2>=9y7a ��T ^��. Zэ*��s(���V��$���}'j���2Y	��bY�n�
��"�s��w|��O�H6g2f������	�ֺh��Q�f%��1 wq#���d��4�gO\\� D�nl~�)%���~�'���vi /����F^��b#sR[�����E=�a��׭-SP� �;5��X~꟔˿��=���R6.�'�~�JՃ��N��]�~m p�uO�\��Lw�y�@�9s5 ���;bW�zz�n�0B/;f���:�II����z7.��y����S�{�蕛�"^��n��[U5�O-���cd�J�g�����Q.�}��/��_��!��dG��)W<�^��{U�hα��e����۩|��S8�p����hX���X��#��n�6�9͎��H�]��=[��c�8�sf�Ǣ붎�;]tvm����[J�u�Î��"X��{tc+Qú��[�A�]p�m�pv�`v�عF�9�ִ���q���z9��ݞ��#�N�Wch�\���_n-ܖ��2u�/f���t�W�7k����z�͛'v�#ݵ�����12�r˕�.0��v�@>>��d���F{:�S��}wI��4��'n�>ӡd�?��;w�mf;� �޳%{��Ꚇ @��ˀ =Վ����:��t����,s�Bj%ؗk�˓�>�YՎ��]2��[�º޽��vN�ĉ#��X��N�zR%�"\���pL��5D����� 5���� mc�����}~���޸ԓ[ ��r���ܕm�L�mL���u��, ɯ�x)��Ҡ"{��p����@'d�2���=s�������y�r7k��-[&�Y���O ]�'��87Bc�]�a��5���߿�vܻX'�5�� ^㸰� �ٞɔ���ruR�Rn�7�n�$D�c��=�id�f&\AYsaçL ."�Gv)����};���o،N�whɼ�+k;�W�)vwi��Y�JG���.y�^�)}�oɲ��5��;��q<�`2J�g#9�Fӿf�����}��侾wQ��A� A���v	����#�Q��/{.���Eo�ϫ�����X� 2�l;/ŀ �v:a |T$�꫗}}f�oV;���N�_0�Oo���!5ڿ�:��Eծ��j� ����PD 
�y�U ��\��	��]�#��* ���N�zT��H�3,��$�u �=�=w1}����n?�e�J���t�@�N�Ď�=�7�{|w�v6���n�e�^���n����=m]z�s�\�H�y~�~������}��k� ���DE�=����Re��9���*���Zn:���=���Q2�19�	����>!��q�~7���I- ��s@�Nؕ�ݨ�Z�{��|{Z�!3. r˛�8t�$�v��� @wfd�T�c�u�wb�P�����Mi�y����R{:)<&)�"S0{���r!n��[�|���y�����O���~�W�M�=����5��~��>��,�Ǽ v9J� ��;w!��ѐ��9�;��皹���~%č孀i������� =Վ�Dl-�ꇙ� ��2U�,i�����%�����uc�9�U6�����g�����5���z�$I���]6�bO��!d9�a��ZAc��v�;���k7m��wg��mr���f\:�r:dĸs2���5��f�\\�D {�������f漗��pĒ�����ț�C�\L��Jz��KO��r^ʏN�{�Ƹz����X ��v�S���N���Ϥ~x��N�B$%2�19����닒 �X����J����%ϳ�� >3�vĬ=Վ���K�$�-�Y�O'��;����/D�vLr�����ۈ�  �w`�v>���VM��Q�1�rژ���g%ׁ<�)���x�����a�=��<4�=X��6=64�=Yv������mh��;��;��R�K/6�����}|�V�ux�j�y�@����p?Vc��� ���P/�l��ǣ��O�}BZ��� � 4�uWwr�^���S���<��+��8��q˫n��jU�N�v4�Z}r%CԗD���܄����	�n�mO��f�;�Ĉ㧱�@uw�zb}Z�P��J������;���Cl��ZA��q�'y�?7�_���2 �X������G�2��1��������W,�e��wz�n��q��W�D��]v��o�Uf��Y5  i��s̅2?������C��옑Lb����8~鸰�  ��sP	�Nدn�����u�v��𤙘�0�7�C��/6�sYg�4��X�y7� '��t��N؊�}^DWg3|=ɖ��uMz�(���<�r��Db.�G'M�'fӯ,��)��׾���y~���o��4���Y��#��/��%U�w���'cS�?�_�q�Kg�:��3ڛ��P����u;�Ǆ �<��( pm��/.�!˒�K�x��bEI9�u�d5SJ@���ej�"FK!�L�M�ݞ�.��3���BvE{d�#�����-�l�r�#���5ɍ�a���s�#G�C1�m���4s΍��TՎ��7c3��N�;'o,u�#Z㖭)�g��WkOco/�u<qnk�k��	��M]�6�n��c�{[s�rl�:�۪�j좶~�||?n�ɹuپ_�޷&��"x�r�����%D_��\J�n�&Vd�V a��Ӹ��VܝӁ�a�7�(񣄎�~+��]�ӡy�qa @l�9��ޝ����ș���u;�Ժ&w鐆�%�,�	;]1 =�=w$ x�S�����>�� ���LD@�N�Ć7��d(��n�sײ��8�9;5�����)C� �Ϭ��" ��d��9򮥻W�T 2�0�=�S.T%3	���Oe��Y7X{cƫ���gs��7�=w OVM�^����.�v�GGJ��?������:Itmţ�h3��N��x� ngR�ơ�7��)$�3�,���}I-ݝ�� ==Y7S;z\Ue��܀�y� |wd�܆�ѐ���i7e��Y�J�Qw�2z������(�
�q��{�y�>2e}]J��;!@�9@�W"�	_��]rz�v���}=���^�~ʗ���">���渿?� ���=E���Y7q �{/�/%{EQ����"[r6B�ڰ��Y7�}��ӵ�E��c��a /��D��<$�����@�d8�$��$�j��#Om������ӷ����r� ��5]�H�r=��O�|e������"fB[�M���;��������5O0ĽԶߔ���݉X�nҸ� ��ɩ.��sdw@��d�I�i%�z�yրS<^�0ر������Ԓ' �?�fD�����r�)�L>�5ӷrK�-݀$l����suk�WR�a�l�����ͬwq~�^$ls�ÖT�#��A9�>��SUY��T%�uc��	��U٤ �=�r�ߪ�0�˂&@C�ZM�a�����vMCL��~���W��q����{Au;,��O&3a�n�-^�W���{k������Y_����Cz�Կ���Ͼ������O��X�� ��&P�aTܐإCt��|㟪u��vh �{� �w&k� ���n<�.�Zp^�w L�#���d8�$���&Nٯ�@��닐��R����=鴒��ܙJ��/zv�$��~��2j�/)�h!H��6��$��6�����N�n�e�h��.Dϱ��f����7��3�M��ϯ��H��ܚa ���%����_��o��6I�E'�!�Z�KP�%�I)7�J�����l�.��� �=�4	+�� ����稽��ޕ��ng��S#��bIft�ܤ@u�j*�����I�4�@+�Ttd#����n�6k2s����%(��4�4MC ���� �OVM�S*Z�J+�HH�أ=���K՗�ng�<Mhޭ͝��I�O^w@���wŚ��0��.�#z0���ϕ;���|���O����aw��Vܑ,%Cv����	S��<�@g�Ֆ��@?���Ns�=w ��d��)�u��ݖso1׶�!�9�ݎ��=c�cnvyo]�gu`Y��M��	�g<��}���&ꎹ�����풽�޹ ==�7`v�ʍ����M'��9@,ޞ�����Ey2`�8!�jNۜ�������
��$�ۏ���/뚸 .�E=�/3J�����o������0D����_� ��f��O�ճ���e+ ����	1N��%�!5�����<��:��˷��J쿀	w>��#gՓw @��>�ϲ�}����.���B!�4��Οg����욆,��������_��w�����	>��� :Nɔ����y�e�w�����7��G��:�~�8f�-s������T�.�`��Ê�`��{�m�/a*���P�r�r{;����s�S��&Llk����z��x�3�7L��tc׺c�4n�R{�u����Z���u5��<x��7+ꦪ�4�ܼ�g�g��{��Z��M.XF�OA��v���[��==��_�����x�����{�\կw7�^dQ轇���y��۷0I��O��G��ޜ�N>�h�s��{Vm>^��뾞@�=���P���^I�P������Ƣߡ��K�NE�z��ɒ�L����o�D��a��T��{�l=��۰���o��~���M���;2�y! ����m�N�c��=��^��+ֱ�1C��^�c���|����9S��/�M[�K��फ�7{��ۖ���}��d`�'�fַc��Z{��Nz~�l)yWk���|��j���>Ү$��=��_?k�;���N�@�Zu"����^F���ZI�܏K=V�m��T0i}�,��?>��� �{Ì]�������]��6�ʴ��;�\<��U^"u^�Q��To����$]⍻ެM�/x�S�=�̥�'��K�_��s�	�7�p��+�{׿-���dOl������{��ܫU�,�R��Q`�=o������Nv�Z���U�+2��3��'�Լ��6��U�Vo�vFp��V��9�"C&�8�r����w	���m�[y����;����qA���Eb���B#�� �Ec\D���"*�9���8���1V1�,��S&"8�$�IWT��0Tq�`Aq���UkK"�q�HL��"Lc1�$�`�F.*�(�*��ĎW ��T`�8���rH,W�6��$��%f*���*(�b(*1dŎEQpQDH�q,��r#�B2
��8�2L�Ej�q�Vq#�I�e��8�AbFb�
��&
�!��QE���1�F���
�8��k��e��X�\�,�qqpU�,a$B�EX�!"�$J�Aq�Eb���D�"听qTU$$jd"(�㊸�j��2dQLR�
����z�����a�n�]M�-�Ǎ16+���k���0j��5�;����g�'�;rn���h�v�!�aɹ��*�Fwu��	�]8���mcF�b�E��86�}���֖��.z춑����>�k���8-�sz�8��vH����6�`�֛��Ź�9. ��8l=��u��^{o!�9�cfɗY��Gg�v����;���ڣ�=v��)����m�2/���k�]���)�Rj��O?���dy�7G7j�'8��B�Zi��ng�㗲��n\�-d��:ܝ5v��z�ې��ì����9-�1ņy�W)��aX+W<�2�V���9�G��0noY$6�ʯ��a�{Y��^'�e�)q�n�8ܹ�,.���=�'��Q[��/��۱>H��/"��M�M��Ch�!㎎pB��kgpYŭ�1�]#�,%t����n���a�P�tv� u<v��F�jv�<�D�u��[gaݵj�����E;����z�5�����/[s{�z��n2���ypog��Ӎ�ϭ��v|��Mϛ����:����m=��抷i@6F��X7'��9VMn ƷZ�븋OR�L�e�^�۶ӣv�m�Ox./��������֧�����V<�/�����]Pқ=�)�8ۥ�U�Tno����vU-
���d�ڲ��M�\<��bfz���2��:���nk��蠭y�h3Z�{y�N@+�z���1 ��<KS+�d;�����XѺ�e��[H ��=<V�;pm�1\.x.��A�]��s���
�z�:M۵<v��Q,h�k�-�5�2R��;�{q��דs㱦�\�|&���In8�X|�]v�{��Ev��G��$b
'��qĺ$=��l�'d�����A��}\��d�n#,(��������`��x�S�M�V��I�{\�;�ϱg��n,\[��	�~�ym��^�@mWn���Bm/V^�GF^pf��q�K�y��Gm�ԷHl,�3-�:fC���4j���N5s����ڛc�����m�V$��l�l6��$�A$�D�ij�6��`���r�q�Pup��v��ptm�O9	��fS۪�nmA�<�D�����㧘�r�s�0,�2�s���l����]0u�^�i>�xxV]أ�t���H��
ۅ��������8�[���<y���F{kN�:y�i;rw��n���ڌ���R�yF�<���]i{mf���������Hу�s0~��q_���oW�9����KV�ń�t�d��!�����;����+�>��l��Q��6�pܩeY2v�C�׳7�u����;qr }��ɻ d��<��}s]T��0�q�^L��%�m���/��� �ܚ��:�ttҨ�S�@$G���v	.ɯ�E�+��J�Zi7p��IY��*�&M��JM�N}���|�{&j �o[p����U�t�zn����yȦ[s?L6˛�du5 Ν��u�^���!_�n�ݤ�kzn���4�D��~m�w�s}}�>�O	�=�a	-���E�3�N���v8�;O`<;��T��#��8��:2;!��&��O�&����� ;�Yp�7]�]��gz�� �$̚ar���!�J��Xk����Y�>9Ѱ��G{*{Ϯ�}w��Uz�������yr�_8��!����W�O�ґ�vB{~o4�都�5��F�ߩN���Cr����}�o����L�ɔ� �����q" *hi�w��SNf�u+�}�l�P�!��G7dɻ5�0 =�=E� W�ײ���,��sw��fMC ��=Wc����	�X�i������"�۷���� �{�L �Ϭ� K웮��Mv�\�{��������45
:t!ͤmOe�	h�&�;"�ߥS����K�$�H���4A$���l�p���W���QJ��A�&4�RĦ\�tcp�����f�z�����+����:y�<o�m��r��;�H�eP�ӷ) G��&��?my�&N�� A��ۿ�4�B	�J!��&�ZVzs� ��I<�^rw�^�� D��l� �OVM�p����L��na��٦'-!
ۑ���n��k��ܤ@aՓqa��yZ�k?
�/��7��	�V	���E����ov͝�Ŏ��A�ޫ��������=:K�w[�@]���ok�Fk�W���u7o���7?G�D<{S?��3g��X��_��{쑼���a�at�ͽvd햯;���߃���,=9Y7 �vL�=����<�W�<�z�$<�"��0Kۻ����ń\�٦,Y�]�p_��%�����Na'��U�KC�esF�K���i��|X���D��%\���]� .�aDr�k_?>�lKhD�i}�9s�r@��Mؑ��L�)ؾ���OX���Y5qy�'�`������pK�D0�8��:7�x.�;G|�l�d݀�I�5�][kJ���>��=��}�8�n�6o2o��/d�J�:�L6��G�����9Y7q I�3�P/�ɿO"�˵�Һ�|B&D#�_o:���{�է7�ʄL�,
�K�{|���#�*eJbTʗ��|���NҦT"dr��o�a�>�����O����������U7�~����g�	[^��_�������}�w�� ��:O{���!ћ����Y�2��}��fo���eBه���jx�P�������ͅ��7�*Nb7o��jv!�2!�T+�����;B�緞��:9�y��(��P|��~�bV|p�p�B�D��|���ΠT��ʙP�=�}�Щ�����N���/���qpv.�U�t�W�� �olyn{=e�Mn��\F�ۭ-���޻	,n�!���g�G���Z��*2!"{o�toa�BP�p�V�=��{ÈT�%�~^wke��1w�KD���-{y,G�
��T(�>���i�}���wd%�5n��qÃP����R�X���uӛ���@�3Rgſw�Z��+qʙR�L�O۾�٩���S+�jer�^{��u��������w^�7�(��g��X�|�J
���R]ݷ)���8��D���S�t�L�G+�
������s�T.%B�D#���;��s�o�w�}�v��5
�q�T����F�j2=��2����>�8�J�R�������қ��L�Go~~�\�}����W�ަq�52�l2����F�C:B�P��
�i�{�xq��*(�P}���X��N��t��%�}�(�J�m��F�؝!\,���9w]M+���#��~���q�2�S-�\<�sε�L�u�<�������gi��2���w٩��L�v52�Z��ߺ�!"2!?_��֡��B������w���z~;�Ϳ��r��}���o�3��뚞�ތcF��bԛ�#��LCu\��z
j"a#�3�F�|W/l*�K����?���}�D�:�1iCV˸��Sn
0�g����T�;x�H9�s�qf��ua�x-�M��	�7[csvM�Hͬp�t�w\�J���P`�p:�:n7iy��ǂ'"/e�v���R��a9��=�k����ǻ+�f���6�����;v۔4�=�lJ�D܅SM��uĎ��Q7|��mZ�v�V .�gZ��nSƓ��d��j6��;�cN4���n�����t'�0I���[;g�[f6�ܭ	n�߾���ؓt�o�"[yѩ��HW.9P�W*���u��s�T.%B�R�\/��\C�jï����o��t��a��{���B&G�ʙZ�|���!"y׋����n����3��J����x�&T"dBn������Y��t��>���B~�eB�*���z�Љ�*.!P�T��y�C�s�W(�B�g�w��q1MùL_1/-_�?"˻$nɫw�C���~�]����*e,
����{x�*2%J�Q�=��燐޼��zT�p;c���y�Xɀ�����n=���������nR��T�L��֕9�K�Y���rR%��}P/�%��dʳ�B�D�TȄp��<���À�+�j2���}ѩ��Oo�u�>��y�x��ʙZ9_~����q*eK>���xY�)���ʜ�{�<�!�ds�L�R�*~����3�/��wݎ�Ͽ��p�V�\�;�!"8T+��s����
��T*T��~�ĨR%����*���9��6a8�Np ��F٨@��&�)�	�n�3M�z꺸�۶u�ʬ�W]��G��_;�tǈT�`TȄp��y���dy�Tʕ*eO���F�jw�S+���O�xߧ?)���5޽��Xq��!�f��7�q�B������WbM�ɽ�P�s*n�>���C�+��3����	��2_�o'��#�4�����Lo¢�S{>k�}����K�
�@�0s�'8G8/h%X����G�j��>�>��j��ܪ�-C�*
%B�_��wP��p��*e,?������B&D"d~����s�^�n�?�g���(�(εS��)v��Γ8��u�\������52�l2�����S5	��V�T+�z�N{��ܝ����D�
��\O~�uP�*2!�E�?l�%B�(>Q���P߽�!��}�/��̥��oI�^.��ݢP/��*e�+������dB&D�%L�s���vjf�iS+�jer��}�XqJ�w�}z�wz{�ʄ�T+�9���C�ȄxsϧW�	wvܥ�{Èjq
�m뾍N�:B�qʅr�TPn��h�ĠK��S�~�X�I�1@���^��C�jµ
��|�S;�L�D��r���z�!";��ߖ�Q����Ǣ}"�V���s��s�Nz��l&���X㩥�$.�n��ȍ�Ѣ�{���5�;�]w���O��s�|���eB&D-�T�o�tod3�-�T+q¡[Ͼ����8T*{,=~>�ޯ��k��u�^~��89P�W*2'���F�؝!\/��ʬ��vj�]�DȄ|��u��"3�{��}��OOyס9��Ϊ�D"dOؕ2�<����L��*er�L�G���]a�,2�(C*p�?��}�����p�������p�Vo��v\��Y��z¡�q
���z5;C�*dB9Aʅ}��tq�!P��
��\;�{��_��qP�՞������oR_r ��5\0�%'���td�Y���騼q��oL��N(��/�\W����yZ�ל=��U-�$���9���>!
�F�S-���|�����S#G*eB<������8%L�s�;;��Ȳ�[^Mґ}b���M����V�����s���u3P���Sm��F��a�
���<������T��B�~�{�nN��o��u߿�!\�T**w��53P�����$٫�w�C���{�����2�2��A��u����vw�W�������q*eK�n��f�jv%L�Q�����<����2!9�ʅ��uߝT8�>P%f{�����|Z�CP�=��%�4Kۮ�Ѥh�0Շ���+&6��uE���~��wm�]��?!��?m뾍N�:B�D"dB>������!�T�T*T+��uߝ�8��j��l<{�'���C�ge��y��S;:�S#\���W�y������Q���_��ͮ���3S�\=�^y�s����jeC��_j��82������¸��O���(��*�
�~�ÈTȄL�G8���:�q2!"	����ӯ����މ�LJ��A�I��l���v�L�G��tc�52!-�\<�{���eB&D�Tʝ�����Ϸ����j|%L�V�W+^~�~�!͆T%�T-ɇ��Ϊx8T+n����7Z�$��'1
���z57}�P|�|���&D#��
���ΰ�
�1*
�
�O��;�qÃP��T�a�߼���׽���:��?͏Ͽ��?>��2��/��v{�j�Z\W���z��_��g=�7?W��;Џ_T���-u�z��M�;S{�^:s�5��/���\/�i��!A��}�'�ʟ�vu��iIn�#���giĮu�z�s&W.52�B�*[��C:B����~�gO�W�B��Ϻ�8�NT*dB9S���:�8�1ʅr�P�Q*}��:5��
��sޱ<���;������l��Ms��D�ؽ��tiޡB`H�P�E3��35.�m�v���ڇ?��W~����S8L�`W���ּ8�[�TʄL��yѩ���L�wᳯ��߼��띍y���8�L�Nd2�i0�~�ε<*��}�_�%��r�u�!��>�z����HW(�B�w�;�7_�v�?�-~����ǲ��Ę�$(B�D�W����P�À�*dB&R��yѩ��P*dk�2�~��j���׿IU�g���&/�Q�Ӕ������ʜ�}��ε�+��P�a�?[���C:B�P�p�W�^��3߷��6{�v�L�D��B�A<�;�C�p�W+�
���~�S5�����7wl�V��|B8q�W�>��߷���|������ë����L���(�2�Ϸ~�S5��������;C��ӿ�~�������!6P�a��=�P��
�m�=��MֳV;���Tݿ{ѩ�!��9P�W*��w�9bLK0��Y��bbR%��(>Q�oi��B�D"e,>�����
��L���������&T���޷�2��/�����嶭�*��uR��4�F���۶�����nܹT�r} �'5Hw�rg��Ã&%b[�Le������Y.O����譀��e7��\P	��'�K�SA>�{v�^B�r��l�m�Y	ێ�vx�n�\zk����tmrk�"�r���ӮqZz�ۤ��f�mb��n�����6q�rs�F ^D��	z��9��:��qp
�����v���]�g��&��|kx�a��g��痶��D��ic���6M.�HJwjK���Ҽ��{9��5�ۻ\���n�l�˹��n۶4h��o&C��Q�;.Ϯ��9�.x{;��vk~����֔��;���3��	\:����C����T"dOm�΍�!�!l2�[�
�o�����
�]u�}��~C�t���]!�9��
��T*T���:5��
�O>�Ñ�d��v7{�8������y��52�%�9�����������|���D�_D"dO�*eO���F�jv�2�Z�\�_y�]a�9�P��	���>�[������κC��
�ns�gW�Y7M�I������K�ﾎ����W*ˎT+��>룘�����o�|~�y��~��8��P��L�a~�y��f�#�9S+G+��>�8�J�R����ղnm]��&T#���?uӓ�dy�M�}�q�Z�P��'/?tu��
�����u��"8�B�R�����9n�����%���3���T(�/W�:C�N���z���$Վ����z����q�2�2�p�w��C�����������dL�?	S*N�~�t��D��mL�Q�=��Èr�*�ʅ����u�y�
�y���G��s�'��n�۔�%؎�5HKʻ�}v6wg��{4�ٶ��'OI����?����=Yű��5�*]�}��f��ʅr�T+��}�G8�B�P�T�W
_������dB8K��=o?Y��L�9y�GI�@���T��+��~�8�J�R��<y]t��cd���3����k�L�_ŋ�>���%��p��]��k$y�^k�Sʐ�ඟtg��EҦ� �V��7��h��8y����$�����;g�ם�3F=~�r2�g��<N���F�j�P��
�o�{�}��"pB�R�P�Q/����8����>�(�&�[�Z.���L_}z�S5��?{��ݲMڻ��p�P����c�*e,
�l
�=��:��9�ʄL�DȖ��>��ݷϹ�}zjf���2�#�k�~����2!8ʅ�����8�*�=}��K�̦�{ÈjdO�뮍N���_7�9|<���T+�ʅwϺ�������W
_{���C�jµ
�r��yѩ��^z����}��w��S"2:�|�u�N%L�rs��4�nm]��&T�W�9�+������yѽ�ΐ����?���v����O�	A)�گ����B�D#�K���*ˎT**}��:5�:B�|o���﯇����n�	;;6����gc'Z�㮶�;Y�7z�d�۔VB6;0�������֤�I&���G��~�u�s!S"2�\'��κx9���*eJ%L�����I��%�}���=_�vVvw1}���}�Xv��JC*���߾u�L�G�]��nSkY��C��B���ލN��
�1ʅs~���{���z��ʇ���}u�hD8�
�ĨW��yޡ�Ȅp��*dO��Γԧ�@��������r����߾�.��Xz�	S*S�9��uڲ݋f�f�q9�\:����C����P��T��|���!nC*2!2?~�r_hGu1ѻ���7�
%{�������9�Lԃ���x#�\�s��J�����E�W���[|L-��\�5���f-=��������ޖ/c���築ݞ`������'/��Ω�9�F�����;�d)���8t�T�N�� Y/�p�7��i�����Z����;����Nŕ�K�v�Ǡ�i��d��t�+��}�0�ୱ+��-���}�ޅ��.����G j��^@�zWPZ�d�-x���Zǵ�5�^Dyf��uI��=���ݮ����X��}����o�+ș�e3�nr�)/b�9��xv�^��=�I7-f8׻{o�ٴ�IӜE�iA鷧z�������z�o����{G�4�>���zU����Bw,*�v��+ۿ��kF�q5x�VZѓ7U�7��h����q�i�SZ�M�n��G�c^�e��|�K�̏I�o\����x,��5y\3rx�H��iV�S�y�F-��OpriÌ�z@;�_d�S(��| �w�����ɛ����}�^+������m�z6����q��qr=�9
ų;���B��,'�F�y"�xz��=͐�#�Ρ��=:@����)}G@?uŽ1*³��꯼GF�.����V���e��pcɕ��,��X�ؽw���-f˦���L���Sީ�z�j.�s�<r��}M�(-2��w1^���?��N�,j���������or�緳�>��=��X�Yw J$��q����]���]�������8��&E8�q["+����"*���
�,kZ6dV�U��2�I����1#m�!\E��QW$���,$��"�
����E.J���$�%�r̲հ#Y����
��
��"Il�*W�(����E�Y+�Q-��3"(GE�$�G+k�\L+$�A�J�"1l��&B2�Y$��r(��$d�q�#e�j��`���(��Ii\��DUQH�nI$�!-�EVŘ��Ă���Y��$��8���Kh��pd�R�X��qj�D�c1�d"Ԙ��
8�#�A�E�ĬQ�#�Ȉ�����&�Q �(��U�-dr����X�E��&I��QTq�3����D�B�R�P�\O���:�8��qʅB�O��tj�t�p����8�������+ J߲e(\�V{����s��B&~�*e��~��ε��+\��(�2����F�jv�2�q���5�}�Xq>{���o�!7!�f߼��C�*����_�d�l�mw�8��*}���5;�
��W+�
��Ϻ��9�*�2�9]'��}�/)�ߺ���+!
�Z�L����ѩ��L�x9S+\�<��É�J�S������yכ��<?����G-�O+��S�:�׌+�\��w���W2vn����_,��Ww��ʟ	\?o���P�29���a�?[��C:B�eB�*�<���ÈD��	@�w�\s_��@��O�R�K�qʅr�P�Q*{��:5�:B�_�O�4�v�i$�{�ÃP�����P���ǒ�}K�0[���l~̝|�ek�2�J�R�n��f�jw�S+����5���8�,2�#�gkH�7�L^V[L�}�9{Fg���$+n����E��h�{�P�pB���ލN���Qʅr�T+�߾룎q
����}ϟ>~��Wz����{�P��ơ\(�*dO��΍L��L��������8��T�y��l�h�6+����'�o���s��r~��z�����|���ʅ,2���}�C:B�P�����{�xq�P%�%P}��6X��ou�w�wAaiz{%s�t�]�N�-����b���	)|������}S�����g'�ۑ��"�<���w��5I��/<�u����}y�T8�Õ
���|�P�N������l����P�1�W}��]!S.X2�\=���y�q2��~�}�3�ȄL�~����L�"ds�jer�_~�޺Èp�ʄ�ʅ�����ε<*甓]�=�Q����M�Nx�<u�÷1�X����ۉN6ǻ&��������`�=M�~Èj|�O���F�j2!�r�_�y�]s�T*T**¬�i�X�𗏗��'}���}
<���tjggP*dk�2�=��ô�%L�s���W��mM����ʜį˝��>�X��� _@�kS^���;��~Ko�7�gH[�V�T+O}���ÈD��B�B�\?_�y֡ۜr�A�#��#�žy�^�Ț�R/���P�:B�_קӛ��c4�k���ơ_��z�8�������}����8�P��*Tʝu����[�u���w�53S�T���P��>�������	��~���uP�dB<.����"�l�3gxjNT�o��jO����y��z7������t��B�G*���z����Q*
�
�~��wP�dB8pj2�}��:53Ύ��g�|����x�G�*ek���?u�B&D�~���ٮіlWogI�N	\:��{�s��ʄL�Dȟ[��3�"�*T�����|�JSuu_+��B�S"ˉ�οy�C�pr�\�T**}��:5Ӥ+���~�9_���kv\P~��b��{��l���@��g��<����/�V��+6��;�%�L ��Ng��OV趶z{��b�IO��z:�'&H	x5q�,�瓟/g�P�,7R�^�sӤl`�Wv�Ž��獸��vU�R`�Q�t<77u׵!�X+����M���8�(5�:-�-����[�A��s����ckPn�7�:�Y�]r����Gl���y��yʻ�o`zre�s/=[x���k<��<<Ę�����]S/Q�/�p�����v��ٺÏm;��3�Y�ն:5��Y��tZG�t�u���
+Ü.S��V�-i�_�1G���>x�L�L��\=�y�x�+G*eB&D����f�jw�S+�κ?w߿u��s��>dr�~V%j<��/G�T-�{�_���Ȅyϟz��͛�e7]�!��>���5?!\��>yn�y<�>�,"������J�P%P�T+��οy�C�ơ\(�*e��o�tjf�#ە2�����y�z��W�����˅�
�
�tG����a�w{8�S�\=�|���eB&D.XeO���F��ΐ�P��\nWt~s[�^ˬ��X���P%��#�O|���T8��W.9P�\J���΍C�:B�}��76��d��]�x�Z��(6���O_*�[���%b������+�o9�C���r�T�S*yo�tjf�iS*2!~��ô?x����r�p�ЖP�a��{�U<*�����t�m��5ӂ:����t�r�P�Qʅw��*���@��o7��)���\$İP�p��u��8��j2!)a�߼���B&G�*ek����8�ĩ�97�O9�����xWXI�wn�Jq���8�M��&/��B����1�\6y����rZy�mWo�I�'ؕï���W9�+��P��=��:7���*2!��3�/
Д	@���_���K@�9����P�dB9�ʅB�SͿyѩ��p�?~��.���K��p��+�������*e�*g�?��v_���������W-�)᭖=�����������WF�+����S>1N���j�׵>��H�Ү���o���V�����žＺ�v��_��>������fT"dJ%L�s���vjf�bT���\�^~��Ès,2�"���������͘�~>P%+���8��̦���58�Ov��F�b!\��
����������P�P��u��&�������C�����X}��:53��TȄL��?{�]a��%L�N_~�rI��a5w{8�D�|�_d������ei��_�}����a�=��:53P����P��������*(�B�~�y�B���^���]ߟ��o�$Ͽ@�	@�=��΍C��
��w�76��d��]�"�����!S"2�-��fG�/����O�/��]�����Tʔ�w��53S�*er�2�F���u��XeBXeBه���U<
�}������<������iM]N��/<�q�w`5���y�>9��g��9������˺Q�ɴ�_��<O�
�m�ލN��
�r�\�T+��룃�B�R�P�P���~�"���Y켞~�v��,/��}&vu�F�S+\��|����pJ�S�9��&���خގ�;N%p���U�#�jeC���t���g��}�MmE~#�Q��D	��������T*dB9S��~���B�AʅC��y���o�txDtt��t�p�y�Ǆ��k��.��qÃP����ô"g2����������dx�L�q*eOgZ����M�`F���/eZ���%�/egY=n�X�R���������󿷜�<ʘ�^A2���J���,ř9ߟ��|�{��S�z��3S�*er�S+�k����XqP�P�2a��y�C�*��_g���7ve7]� �hJ��T����u���	Y�|}P�W*���룃�B�R�S"�����wP��p�B�R��~���<|o�y�f�<�#ӕ2�r����u��S*^_>�rI��a5w{8�S�W{��:�q�er�2�K�?G�4���%�B����}�^3��P���:�Љ�
�JT+����:�v�*2!�T�_���3P�A���!����z��!���S	"P8��)�ӻ<��Ҡ!����uk���m���������lt����!>j��{�A�x�L��S-�\<�y�x�+G*eK��
??�JE�!@���g��t�����u�B&D'2P��{�_��ǃ�B�/�?Zl�;I5�C��
����'b!S"�i�]y�ju���H���eo��%P�P%R�\<�~�C�5
���'��::L�:�S#G*eY��w��%�����u���S*S�9�r:��b�{:L�q+�[�=�\����jeB&D�_|��gHZC*�
���y�N~��=�����a�"z�B�*ʞ�P��W(9P�\J����!�t�p������Xn�d�֡ۇ�G߲e+��~������7��&/�%�}�`W��s�x9���*eJ%L�=�y��f�iS*29F����u��}�U�>���_��R��0���ҒAl����ݭ�ۉ�q�;eV<�es�O���t�}���i����w� 7��ٯ=���ΐ�d2�nL:�w��C�1¡[ϟ�^�컻3K����ȓ��]'���Qʅr�T+��>ӎq!�O�������ĨW
��yޡ�5
�q�T����&w�@���Tʄy����2$�޽������M�j��6>��b�(a����+��,z�qA{u4��a���\�ۚ0VO}�͵�nֳWw��ʟ	\>���s����jeB�R~����pΐ�!�
�¡[��}�C��
�O:�w��[��믎����'[�}֡�9��
�r�P��/��&jü�����l�Ѥ�{�Ø�+�9���q2�y(�n~�:��T��
�.>W�,��&V�S*Q*eI��Ύ�5���ן��p��2�.C*��A���?�]���X�A��z�C!?G��Y�xj`��y�W3�̘�p���nv�"Ď_k��Ǟ�������C����P��,/��::L�"d{�������8�N&T���9٫n�-��&q8%p�~�k�����?w��B&D>��?_�tu��
��*��}��8��
�B�A�!c��,JϷ��?��J(����@�ȄC��/��z:L�#�߹��]k*��.��v��P�����&Dy(�J�Gf�,����ٓ��uI���L�5*eKw~����NҦW(52�Z������2!9�ʅ����bVY�(;��ە=d�ń���.KUj�:}����9J�����M?|�8����>RI2郗�;���B��o^\ͭ��pz��f����*&�F�a�ð�E��0ۣBVQ�̆.c��s旎q�1������+uP�u���f�bŬ���R=��V�T�sn��]p ݐƸ�]&w��{Vuq\Z�rz1��HhC��q�p' �k����g;����E�������g���:�6[F@�%���k���rrq�Dp�Şݵ��+k6���G�]!��v"��¤ړm��\H�T���_7���!b�F�Ll�,h11/'sȮ�8;;csz�&����/�v]ݙ�������/��}'ht�r�T+�r�_y�]a�%B�D#���~�C�jþ�������qS.X_o9��f�#ە2����Ϻ�'�T����l�7k$����T�Ww�|�\��ʄL�^���܇�f˂���zcJ���D�!�
�¡[��>�8�NT*Q
�r�����js�T+�r�P��z�~&k���:�s���B8}7��t��Ѧ�z����+�=��AǈT�`T�`W/߼�^9���*eJ%L�����ߞ;�����5<�T"dr���}�8�2�*�ʅ����:�8�p�V�>��]i��m,׼5&D�~���������]�]}|����TȄy��tq�!P�T*dB8}~��Z�n�p�B�P��_���3��U;��Ԥ_xď�_A�=��g�b"dO�u��n�[u�-��3���u�s޵�<L�PjeB�R}}����!7=6�����	Q������!�T*T*�	���ε9�ʅr�
�����GHw��}S��/�&E*��D�Chd�$�gs�L�b2���>�;����M�# HQږ��|���%n�ۿjp��W|��t!S.X2�����:ט�+G*eJ�2����GI���S+��/���Γ5���߹����,2�"�?o���P�dB<�~���wvf�M�!�dI�뮎�5��*ϻ~�{���߷���<��כ&��u�?U�� ��N���3�swj�=8��ǡp�7�g�c>|�:��{1)?��2	׾�>s�TȄB�P�����P�ÍB�Q�T�a~�y��ggP*dk�/�ޡy�t~����M����K����q���l�l�I5w{8�S������:�9�+���
R~�y��pΐ��@��	x��ڿ+�W�~�����o?�/��T*T*�'���:�8�*�9P��'��::L�#�����Ҳ�V��"dB>u�:�<6���=�{���T������+�/��Z�s����2��T����gI���T���\�ן������/'>�fq	�2�l����:�8�p�V���o���	��^��8�B����GI؇HW(9P�Qʅ{��ts�M��s���ژ�	h�J�7�򘕟+ J"2���&w�@����/;����|(�,��ʏ�gTg�r���0�kWm����n���8.�c��z�ung5Ym�n��|��V�a~:L�>�u���Z�&W.52�l2����GI��L�G�
�o?}�}��"q�s����K/��Qs�p��_��L�G9�T**_��::L�#�ks8-7�G�x�tĬ�Z J��g�"g��W���~כ�7�qd�����A~����"Uin/�B�Ϟ%q��M@�-��,N݆�NU@���$�'{yj>����>�?Yy(��������ۥ<�\N�l�=z�D�d@<n�Z���ۓ�����M����{�8���� � ��~�wp}f��`�A�M&�K^����p(�7��J�NU GvuZ�H���w{�͸6ˌ��u���d����-�\@uo�ŀ;��CY��ޮ�n�\l�9������ǻ�����-�����#P��:6��/8nۭz�d�0����u�u��{3cn�w�7�&�̂s �������w`�A��;�
�O&v����d��L@ng;�#�G�ᱥ2�L�Jz��E�WI�G��Mx�Mx�r� ���j�I\�c� uq��)�|�{{Y^{��¨m�&G"�sW;|�,>�[��q ����n����.�No� 3s]� ��{�q��ɨ���'�\݇O~2}~�ϔ��W�ao�Ұ>�w��� q��C]��*C�~V_��~7���w���7����;�x$6{ �j�YHž!���.G4�������o�p
ޱ|XI��D[�oTy���ė}{|����|�e!4��-{� /�UN�;�/ٓ����wV��>�c���N�*R����������&���m�j2sQ��k��\���h�e�&w2��م�_���$L�JZ!�|�� f��X@$��sA^늪���[y�i�Z�%p��w n��.d�����v���^.S+.�jfn�+6�w���D����  ��S����x�,'�n �=��KSL��}z�\K��)$�/_����{)X��v�D�����¨n&A�e����3һ޽͘����Ҹ 2s�'	??~���a���z'�0 |����Zɨi9mJj\K�a�ӯ�| g��-�±L?j���xeXWw�����i���" �������+�!-w��v�mNW֚�Vk�S���eLK|��T��G�?u�7^Z;!�y��_(Y�B�L�9d;���z8�g!�:��K�<\$�W���5�A�/������}tt������%����W�h�0��]���W�kV'��`�(�BC��e�s�����+��[f�� (���o����@�㯏�OmC3<g!3I����מ2'9��J~
)Z$�y��Җ��e<��|s��L8���]��s(�%�����Wy�����w�p�;-IS&T�]ګ韦��g�c\{|�_�J�}���<�퓟���w-0�
���`]��%���7��}��l;�J.=ܗ]~��ι��u�Yu'�˗����cu>#|��G�G���K'_wb�aܰ=��|��Յd���<Z��9���
�k��燮2�1�����s	�+ۅto��6���ۑ�?=Q�P��k����.=���8q���C�d�ґ���=a����_;SX�������g�{}�<��ƅ�f�{|G�x��g�r�u!"��h�FΚ{0���i�W����m�՛���k�ō峂���o-S�`�}���9����	�x��)��w��-�S��c�j�jžـ'�a����x��HcI-�yp����t�9xK�����W/y��-�b�lv�oe��T��҃�mx��M��7����%P�1�~w&�	d>��xC�7�8$n<y���U1z\+8�����z�[��l�|��eR[�+��s�n��w�D�]���"O|���|%c�2G*Aa"��A)�� ��R��m��qB��j
,W��� ⊤��+1�B�#�E�bE��lAF�G,"���$ �qB&[hT"��qEq#0F2!�Q�,�H�P�,�0�h[��UTr�W\��$��1��Ѩ\�H,T�lal,X�����AV2�X�QUR$�R*
�F A�%��E�,�.!$�D,�8IEB0Y�!E96EQB"�L�l��l���)AȲ!���+�TY��X�T� ���H��U-�� ȑ�F���#R
�3 �����T�V1&B��	�Ub�JXƳ
�H�kl�s�]�?�.�<�;�{�v3���5�N�N4'v����N��Pr����g����i`���g7u�M%��R�V3�`Ë���jc��K`�
EÀ9�������mS�F�6U.�%�Oa<���s��w7c��,df��n::Ҡ�K̺�]������9ؙ�{]��g#S3��h"qz�r�:l��v.4�����a;'u�vގ�+���ӹ�h�A������u&�X`Gs�M��;:kb�,m<m�۴&�#i�c���m�����eۋ�v�K��<ۭ�J�l��{��ٱ��me뫈Ύ�4�]��x����o<�ާ3��5�N�����M�C��5�=z��3�u�m�{R�՗⶚�$�;-�"<�۫v��yx<�6�8_i�.J9�WF#\��ݻr;4�8���o�;��n0��ՁN���]ٻ&�%Ն�CQ�4�"R��-����v��Ci`�^^yH�cgZ��vs���k�g\n��s4��J�P���9=�kpj�q��)�#گ�s�{=��aÒ�%'b<V#�������㛮pgss6��U\�us�Ғ;H��,��Z����Mn�=wG[n���)tl���@Z8�v�V��]Ѵƞ-��OI���m�a�N�z���mp�W[��;���n\G��	���{I�������rq�5i����Y�r��h�kf�T��㇩�wNx�1O ]&�s�A�u��=�1�{vr����3�n�Ys�&,���8���\q��I�eC���#u==�K��uu��U<$o)[�Ǻ+��/+v6��������� �tv5��(��n�	��G��ۜ<���x\��Q���wmO	����chS��ۮĜ�"�B�6�w�eX/n�FCڵ��q�ƭ� �9̮��m<C�Ј�ۍ\����h�`ܝ;�7�vpI�^<��|7�|0�~F�:]t��j^]��]����n8������i�3�ry��qۑ���4�-�|Y��g���M�v�[g��9N2vۀ6u�Ӌ�^�U���(�� �n�z�79��LV���
<�^��Kk��u�v�Lޫ�X/4�kX��ɑc��}uW��Ě�#��egbm����X�p�c9�a�b]�k�Hvq:����GF�ݷl[ݕ{5۫����Ҙ��F��t.]dP�3wn��<�����Њ:�\]��v�9m�����^u�j2�m�_ߟ����������Ϭ ^7C�" �wU���W�n����'�1�;�  �q�0�*�H�ID��D;W�U� ��O�jsB�p���d��5~����o:�D�5������OzG#l�s(h�n�U �y�X N�SC�|ѯ.n'��l���M�������Q�l�)�@��Ҟ�v��n�=p��Q ��ڵ`����O���wM*�� <:t�37��h�����	랸�H���wCO-�9��Hw�1* ��ۿ�I��̟����f ש��5�7m�p�Ms��:���ݲN��S=��kaۍv�ِ�y�4�i�Ը�o��iԀ��۹" �^�c��]���O�=2sN�G�A���rZ���P17E�[����W�*.{w�%��z�E����3ט{�-����O�3�6��t�i��n�j&�d�π�5��چ�_h^WVj�s�ɤv-���~��MοD��������:�G�F�����"�1̒�i6�t����r@$����*y��Ӟ���&�@�f���H�>���wpv�����CrH�ӯ}�U���;�p%������3}�� ��w���޾}��� :r�4NK���7��t��k���u$���׶�+�7=�W��ye�7��+��D��z�f�y�:�)e��#aBd9��t�8ph�;[�'O�`��
�ɜξ��{���$�����;qr�w����>즫�Ϻhʲ5)���z�D@�c��#kє�I���K�v�:鴪��n<��Vר������H���w  wcu�"��i{"�[���ޑ��Na@�ݗ���"� �^�m*� $w*%���-U)'��ג�h� u�I�s��޾׍�xm�TĽޥ�Q8�ս��jJs3�O����o���G����n{�A���ϝ��)p,�c��H���� [Yp�2J&6�v� 2�����|�;��V%��s��b@fe5@��޼��̣��I�Ĥ^��*E>��4�drRS��  {N�y{;�_<Z
}��� }���/�����{}J3V��Ei��l$?�#�(�%��J;��V�n�#YW���0pr�,<�?>���uͮ��]����[�n��>/5��D�B�}ź�j��� zq����,M���e�����Y쇾��sq�w�-�Ǒ |��j����g�"	?���^�F�c~�����[NF�ĺit�|	잢�_{�7/�����y=��$���g�䵽r�Ne9�t\m�ނ���u�Y<���  7�;E����ǰͫ?�����ny�F�}����wG[D�Bgt��u�������xS���22�칥��j�hf�Ӷ�ba��� �;m*��.�f`�p�!ڰʹ�,����&;�`����d�˦� ޝ�� A��w]�O��=�FU�ܷ0�R�W6q�gn�q����Šl^*iinkn%5U���+r6�y�$����9�.g8kiP�����wad�ױ}�]L:x�@�O]Ğ�����p�875��qa�\�����/5����D��}bW� {��� �:4ӻ�a'�彐�nap7���	�]� -�c��Oݵr�#�\�������H���:J���m4�n�j\K�a�4�kqN^�2.)#������ @��Iߕ�`h���Ko���$�s븐��M̦�9�A�.�q��$�����#%X�v�ʀ7��e�$|n{��vM3Obs������MOmr��K'�e��@2^���OU�{��=�M���̊}XUex�S+u
mֿ�u`<�`���Njm|������~KOgm�p�-�Ā�C����&�:���nL�
���.bv����ݘ�t�2�$(<n��3��u�mzҼ+�c<k���V�����[v9z^����	��5l�5uy|ͷgoi�e�������N.6�qS1��<%
A89�fOd��g+*�C�;)�ga*���;>79�5lUۑ��rn;֛&x�uA�:F�����V�n�p�	[���:�.�՘ N[]`����O���z�fbe8�?/��s�$ �]��	9���R )sw��⥇��[D$�Yu�$�=��F ����K��!�8�����3��PU�NO�� ��{����N1�W���*%�و��y�qbѸN���_��a ���SҋS��^_q�|g�j� �d�f�d���2F��w��n˳}����[ ]7`	zgrf��>/�=m���!���}�RNj|�ޞ�@[��h[�^��SPĈ�O\\�wm
s���<�\�l݁ |t��LD�~��yD�9�k^���D�n���n"wp�I!�	2��e��o[���m`�u�n��n=�����_��L&��q�[�v ��rk� D~����3<�3�#��E'�d�I�������i�$ʑ�
��2�z��>Y����ƞ���o��o�b�O_>6yK��xD^�����ݜ���%�m�=?��t"��0��>)H��׻�u��`y)q��2$�K�H$���/���8L����s�Κw�0�h�Q����r��ݎvvj@����������{�u}��׶{� ���� �rz�$=��7�7��ړ�eNn��i=�����fS���"3�����דo��y�V�[���䰙�s@v�M���`C$n�'z}E�m��gBܲ�^s��� �$�|���>��������%E}x���	�8��>q�#���BE)�1e[����;�%�Z���������pچ�����*\���F�G�������b�^��;[���j��P���HY�36�s	�D�Vl�T�P���C��.j�H��{2� =5�7`���I��W�t���9$�R6�C��UOe� ��7`�y��Y�jV����/;�
����R~Tѝ�f�]��߇��nY�1d�j����c[��f�;��7��NM]fY��5wO��).�{���$D���&� �4�I*�2mI��$��L?_�U6��Oy�ͣ�'	9�u�w t�9�6���]Ub�I+=�9b�y���l�-��sjG�9a ��R�}}���>}�� ��d��t�9K}��vm�q�]�JJ'f�vM��˹�ݓ
ӹ�_7[ћ������w�^��*g۟���&�C$�J�&���%�nM+ �{*R[V��ĉ�>���N��" ��d��{�M5#��pڗmq[�͖!߿wxy�1��� ��x ���� �s����B�{�۲f�$�Ж�3��W  ���p�I�������� ��N�� �s��\�n�L�`��K]>�x~h~�x�`�BNa(Ω�  r)���@8X��3���H����|����uzy²���G��ȷw��U��nt���������� p^��x{�B�Xױ�ğ���o	9���	�ڇ2n�s�� K�{�.��¿xeV�̫\LH�g�q �ğ�Y�w8�����Nr�PSj[hjU5��i|�ۑ��89%�[A�O\V]���d���ٝ���%�3-���f��$���U ��ާa8��Y�m�ӝ�w� |�n���ɸ%�M��Hݤ-�Ϯ��ޔ��1�6}` .�6� ���qB '˼��Ǹ��gMl{��Ԏm�j]�v�����t�^w�Ź��r�wM{3�� @�7@�>-f��E���2��*fR�v��o$�{y7>s˺������� ������̩���t���$�7{0�?<�jT�*F�>v��]�	a]�v)�J拙�<;�>� ��4�K���~� ]��O_m�M
�3][}6�{ӚO���t����x/b�
�n�ls�V+ۅS�{�Lu\'���s��f����ݽ�W���߱���J���^]��nU�m6�ػJ/v:m���sm�ы6�0�\���<))fy�X�W�L���˽���>Ü vy�r]�/v����g����l��1l�v�u��[mЁ
k63]+���n3s���.ݒ1	���[q�bw��$�n�!��/U�痭ݜ����݁ۅݻ�ln��-�h�ݡײ�VR�L�Dri.��j��jM��;k��z����
��+s���_U���r�$�';�<�9%��FO��n� <���� Wc��evNL����Q�;����U A�;n�(>y���l�ɗ3w �Ұɢv�����!)OѨ���	$G�n�%������#���*�7���̚�Z��d��B޺x .��v @cѺ��m[W  y{z�@Wc��#or���-��.��s���N���.� ������ �+1��{�g\%��횽�p�I>�|K��H��h�V�^��[�+�.����\�ٜ�6�)�L�c��pe�;� ��si\�̽�j���Bm6�y��q=\���5ɧ�W�6+Мe�8��ϯ����H�G�RZ�g}t|	a{�v{���+��������.�@a}�V�EM�M̿��3w � tV^��/Q|͵g_�������O�Iu{�g=Q�c�����k�4~�
Cү���-b�}����t߃hz/#��L���S2}qӼcJ�_t] l���� @w���D��ڜ�B�rfq=lI��:7�	jM�uw�'��H��Ҩ�u���ڭ߸:�ߢ &�&����Gfd���'L�wa+}��c�{kw�X{�i_� {�MW����,��^�O�O�E����}���9n\2]���m�D�珂����1�	9�G�7��$�{[IP�޶�N̊�8�en���50���֋��ӎA����vys���459t6�A#��)l�&a5K��zv�7a /{[�"�޷a��k6;K�n]\݂@o���!k�ܐL�#m;V��]�%6�$wg�gb� �ST	�~*�v
�ɤ��xQV�Mˆ��3w5� -޸�,����u
�O:S���.ON����}�隮U..�и��t��ukn<���Q���ޜ��NsoE���Aw{3�m��%<2i�[X����U[�l���P����sx9�}l���S�YfI{^{d;�y>G'���a�����~�qﷄV9�h[M0��h/���d2�����^�9��"���V�o�2n+�hh��qr��$�6yL�u�9�=���y���$eA�G��!7:�]���H�H�4ջ>6<e��E%�r[~�~Y��a.�g�RX�:����$��/;B׉_e��c;��ty���*�珇��Ɍ�g>w���O��xn��V4���~��ލ�pȬ� I	
1��z��ir�ʷ7?�-�[�"�"���faS�9��3�"
��x�`�,�5���FOH2��c~Ʌ�hR��O��g��A�D����^�r�m�{� ��x���rp����^�)���?N{�VS�'v�D�̺ߟ���2�93���T�ȼ�}�{��xЭ!��Ov����|i�r�;�k*l������p@]��xl��Vb������4z~ߤ�=�N�T>��9���z�y���o�i��<(F>5������g9{�O��ݺNH
7�}��}~����tu?�J-�����@Sn�;;�;�=B��^ʼۀ��nT����Y1Z���Ok�nMm.sK�y�Ο-�7���	E���,�NLa8iOVoEl�|���t���b.ŋƗ��[p�o]�F{R@�?`�� �����""�Œ`�H�*���+�D�"-��$�qH�(���㕮c�-��Z�+6�d�RF
$#2ł�b��3-�I&5*�H���4�iJA�J ��E�2��9YT�21�\�ģ�����[�E,�HD�AV+[!"���`�X,�m%\� �!-ʤ�����X�H,�$pl��kiEZ�X���X�AbAD��$b(�I �X��R�+#	$��H�b��H��E�Dr"�
ɄX�BI�0$$Lb�!H�X1�d�$���	mZHb��`��dc"�c	$a!"�����.H�
���0�L�W�!$XLa�2E�d���IA$q*Fɉ �92E	20��E���E%�E��o9|U_����� ���qyd�68&\9��v}�T�{�T .�m$� �ݶ�&�&ɞ/k�{ai� �n��ܶ��M'-��J�˺ /ro�\�=ݿ^w���� ��i*�˳n�D�ɻ����Ωw�M9���n��=>uM�X9�웍K^�e�ǵЮǮ�����g{9Ș�9n\'.�-�� )<|p�I����'���S��~�7��[�ww�t�Vڙ�MC%ڿ���M�az�;�\u9\����>�� �>��d݀9��خOݵۧfU�{ +�,d)���mXj����'	����2'�L�gt���W�[k �Y�m+���M%g�QV�Mˆ����n���L�L�V�β� �z��  "2orn�Zv9����s�1	����	'����yO�7w`<q�M؍�o����|���{�u�=v���c�r���ݞ���g/p�����m\e�q)��Cp���	�훋�.=�j�_CV>U�� 9?m;�>�y�w� >�5 ����ۃG�u�YpĐ�r��gd�T�YWs��͹������;war87&�u�����a�(p�e�w�+�.�$��ɸ�� �� /��y�V^����q�MO���o�ND�')����.���yey y��wm�D�5`����9p���8�Ѽ�{�;"��&a5�jΝ�M�a ��s��ß�u;G?։�P&��d�O����{|C�$B��?&��IJn_�=W���w��,.=�U@
�ޫ��N�/Ue;�o�G�D�^M�f�������9���s� ���������'���RMVD�d�1K��K��~�̈]��^�*'oe����wf>��HD��7ۉgtF?Df��+9,����{5k����K�ޙQ�lf��K��4N��oLD3�e0"Tеj"�����]��E.��U���.Lm��n�/\n�Mِ�Zf�Y���u�ս��:1�m��;c�s�닫���)&�d�������y�Y���@npTV^1�΂t�)�aB*(���'`�Ó���ƣm��u�Cs�Cn{-���̑]iW.ݻt�{��t�;r'aᇩ.C�[GObU�%�1����gx��7����4��Ri&݂�7��/F;v��W�zzx79�FL��u�2b���9��wM�bIq�r�@��\�$����s�}G}�l݁ |z}�h�3-'-B�&&[���=�l� �yT��, �uJ� ��޻b ,\犽��ȷ�L����-����m���R�C���<vݰ ䷜��L9���Y��{�|��r�J��;��aމ�<�i5�jö�߽�2A�RI��s@���M� A���fqZ�iM�&_9�>��L�[�}6�6��Ű Y}��s������髩U |�n��� e�;�ش��6wG����vv�͡<�nH۹�{9���q��1ӶͶ�y���痾�&�Ї&tw\���{��| ,��V#�~�3���%@|{�u��2�e�Cpᴤ���&�]'�!����|u��=�W���}Ĵ����^�z~?{ �W����H=���ܲŸ��Ņq����Y/�0x��l�����}�Оz��H���8 _c�����>����n�.]9�"73-!�$D�D�v��{"����ŀ��0��N]��+>{�u[D}�ҽ����$N%�˹x-z�'?yk��bՄ���[o@$�������s���ԛ�&_�|���?�L_�d�ssF$�����D�8H���	�p��j�fs���+��ɻ��h���S�uT���=�Q��Ü��k�-��gd�ʗ9.Iy��$�͛�i!w���zk%����>�F]o@8M/�<d� ���� ���VM��^L��w�t�d��(��W?&�Ї%\{\������{�;1�:������MX ��s@��].ۮJc8�X�츽���r�6��7pL�lҸ��r�@��=��][�Y�8<_�������>;��Z,��y�\����=Υ�~��ajuπ���:�!y>���#����o9���@�̛����c�s1X��B!�C���'zs�\U� |8��8@
���X@$G�2�P Ay��F�w�u+���ۻ}㩤��m�r�W�� 3�=D���]J�u�X-��V d�9�D��up4��ϣ��Mk������:xV�ܺ�C�ㅌru��v�K�u$��Y�$�'�~}��5ؚj[^.���wa @x�sP������%���Ad��nS߷E�}u��8b�ut� �h&be���a�|�����$�����5|�,H���U� |9��� +���3���ĨUN�x�9�|�.SB���s� ��{{��`]�Y���힐���I\����u`}�U�>c�p�L����Ю��e����m��> 3�Ε� }��mM��s��U���o΄�(2�C?��r�0��y�3S�8��Rj��)�A�D��A�����l����[3��,yٗˮ;������5 E��W
e���wpݎ�� �}����w^��q����Q��U ��u`���up\ux���V|�.9zD��|�å��
�uq�	[d�×� �dлsi+�������.j�o��}7�~@ ��5����wa�����>��:}�RU���Ҹ�J�����2�Xs�wbY�8�9�vu��"37��W D��w�f���kR����s�|����f&[�>�W�|�, ��t� P��쭉���㜭�H������g{�������.SB�s���v.5��P٣��y݉ |{���   ��9s��^��k�w`G��Ks�K��dͤuk�� |{\�@El*e�L�Z��h�#=}V�  ��;I+6}�jQ�~z/[/,�������b�Rzʪ��;ý妖|���;�G}3���˝�9����#=q{�~�^���)N鐷�AR�*&w^�\�^�n��[��p'Ds�x=QۭvN0�ʮv���aW`ݮķ^�n�UH<�pηV���4r���y���x��tfm��	��=�v]c���5��3ٹ�t6k��s�q�]�������14 �+�m���H�j짶��B�}\�d��]�7hC�6���ee���s�s�)r����;���v'Z	6��J0�z�/�vܻS�����M�7l�tٸ���J����ip{�{��?�]�t)�@C��-������Ĉ��w������U�z�#�^��N�o�_�� ���@o�ڇ�8��7.�Ηnk� #��E��]}�}` o��W >�)$�Rս���\mV^��"3Ҳf��!��v�^ۿ�  Y�m*���c�>';,��;��}�g{� o����H�h������pw�ݞ/we.w� ��f����sj� W�Ϊ9��\\xY u�w�."�P�.SB��n� � =���,��g&4��(+{�� {[��s��.�3���,7q��\�H�ɗs)�mK�G�{wo]����3ju��	��n�_����>���&L�|Y��Ē[�n� >��J��:�w.�в���ۮ �6�fG��IsO�1�ςw��X�}�=��OP��t�U+��M抶t{Bkr�MVSk=i��������%S^��E�Q��ݜ���nnS1Y��H��O#^6�s��I��K�� �u5@�^o6�	�X[V��B��]�ߦ�a'=!ژ�%�˹�v�@$@g��+ =�S�ji˝|�" =�n� ^w;�;ґ�K`Cj2�Xvյ������~՗�}� �7P	$F��ZJ� ��v�ֺ�P���Q� {��T�ԋ����&����u޻��Y}����UU�.�mP$��w ���t�� ��٪�48����<�3�{�^���nX�.m֜v��t����ߧo�өa�!��{�����w$����/ﮪ��6gO@OL�D n{�S^�*$����*��MP�6��Ҹ��Ε�����(��
v
3-�6��b�����w[Ȱ�>#�q�(H�������{e�W��e�X}��� �?k�ߗb��wc�É�(^L�K5�5#���.I��w>Z����� 2��j�z5����~nk�9�zn��K�/���٤ ���">+��z#�)�A�7���uz���g����rԠFe󓣺6�k�:�ח7T�F��B��ru״#"�x��M��朡2z�7 k!0U�$�Mn�nh�����y��2"!{МF��[U@!en9
��~�w4�b�՗� wm�C�^c�Z��TCnX�䥏9�,�t)��r������r�
���(���eK}���Gz�t�c��i�����r�}z� �,��ӫ�;.��kq����vb�*""���h���Jrf���B�r�B���)Yݼ���K�'������,�|_]���|��b&{/���"΢��ޅE9��\Z�#�pb(OJ�r9��8�����*�w3nBg)����~�6��s�k�( �����^��[���յ_��P G]�Y��H���_{|c�?f�t�f�)I�����k��
i�lk�]����ʆ�&�	�B7��8hS.:�(�r��
�{f��{�Ez����:k��-��('�ORq�/zPAK'���^ߖ���� Y���VwmP�Ǡ�ó7 ��r�>�Ǜ����'<� ����T.1�ꪸ�4ʊT8�S�.� 7��}�U�u9�dJpڑ��n���Tz�}�w}򊾖� ̽ʯ�#���#�ѻ�(e��;�A�U��D7�?��ѓ�9��V�ȟ_{#V��ch���u��@�]�N����w�,/�ϻ�&�\���S0?]���Ŝ�	U�U�Ý��Q=�hz�m�@��
��@�rYL>��w[��1Z�Ȝ[+7�M3cl��8A[��o���O?b��{��o!�[� ��>Ğ�d�_2w��p��k7��Vj��f�o�����$
5��0޷Ĕ^+GCMԆ�&f�?�͘/H�'/�Z�bo��9�~���y^���U�It�(��ݚ��v���7��v�5�w��~��r��7tu��wQ�w�ߘ���a�pTy�p%7��{����T�ʁ��43�.<��}�ۣnymag�0��=k[𝝯k�U�`{퇝Y�P<�虁��ۤ,{�S%fy[z�Թ�,Z��1��y�v�|�Cg����2ך�gf�ծW��Ot��n3!V�7�*<�zм}[�ik=�{=��=~�>���VE�0�z�-\a���b]ܦw��:A=W�s�I'�OßTkOT?������^�-��^6aɾˁ�:a�~"}�;sn{4�tz�&Uc��*�]�����g�\��,��)��=N�;Q;Sq:C���ӱ�r������ӗ�<J�q�|79���ݚ�w�ڧ+�_+�E��#���o���wH�N���>�����4N��Y���Ģ�K���c{�7�\G�r�z���=�A��V�{��z����K)���A9蔜^���ֽ�7��{<o�������{���Y�y1K���qx�]}�<0k���8�� Ȋ��8̐fI��\d�R
��ȮH��*0cY�+EX�c �� H��DU�G�c�"�\dURAc	��b"d�&Ac1$Q�"��J��$Da̂�$��b�ɐ&H3$���B"�0a �1��1dȌ�	$Q�a!1�#�b�"�,�+a$UdFHF#YT�`F�B ��Adq$��H�c�q� ��Y0aV$�2d�"����G�pI�EH��$�Ec�!��dc"�(�d��l1�X�\�b��H�`��HFH\�HH��8����\��$�$V1E�)"�!&B0�H��qYEqU�L-�e�ZB1�e�$aTŐ���p�Y"�� �B##dl�,dW	+ �F
� ɓUc1�Fc&Eq�QL"�RfD���"*��$ȋ��L�!�H�����H$�	&2$�29E2Fd�"��fB�L�(�	d�3&&.(����L���U�W����n�����k[��/�-����E=��d�ف!�u�;f���X��:�疫r�l�Mu����aD����+��n����[��3�SG)�ֻUH�ۉێ<Y��Of��]�r�l�Ν����կno��k���!]��z�h@v��c���&5���u�勝��u3le�t]-�J̈́�H3��N:��B ���N����on����sG'0�7a�썻l��]۝����4���������=q�mN��%ܪPu���H�;�MU�"�T��=t��&��;��-e�&�n[u�nގ&�2�k:t��&�䣣��qm�nk�3v��M���|���j�vǯ��nU��덀�֣V�m�9,2�)��[p]�0n7��:6�،�5��['uۅ�,����-�1a�ui�ٸ�Ue!�]�\\!ԗTِ�;V-�I0�ꬭ��؋�u�ugi�0q������V��:���ú$�]��wa��v�7&�K�X��-l����Dq�N�g�W��9�F�.�v���v�s��=��m��;�.G�c`y�`p�U����}��H���ce�;�.ܧFR��{j�j�<�����6���{��������*{\s�i�۹��=uʣ�<Z6�ܨ�v�76]�[��m���t��8۷9l��ծ�pn͚ú��/��Y����ݵ����9�n^�|�]����w�9������cm�m��v�cn��Xw]DN�GN=f��M��-v���\�.[��6�헜x��ۉ;z�ë;v����x��D�mu�[��9m�֋�����<�	��uη.��떺�͐��ph�o�*�q�Cq�7Y6��[�b�㫊@7��c����;��0Mƽ;�ܼ�vm�9��38#a8�I�f�)�˓2�oi4c��7!�r8ne����cv��n�Gk�s���n�^N���)��7�u�`��H0�=�u�y�+7
�L�s�[U�^�.�C�=�ѳ��;%v�@� ܤ����t�҆��Nރ���[��c�#�J8s����v��
xpm��;���,Y�[+uda
:�K2�,��<�waUCt��9�<s�V� Ȝ� XV�0��eJ����:�K�L ���h�;r;�v(o�c��V��xx������vv�P
�i�8���+���nt�0����P÷X90�����Yb��a]u�n6�������cNnj���$GT4>:�r� ���e���]����3��ك �=[��`>�n?	�x�jN�/�������͇Ѡ�_nU!��jQrO��{'`��&@�"�Bp()d�VQ�!ev9	�[�ռ��Tk���_.@��*�}�����(�$�drFON'��Qx�Mú]�ԕ ��s� +z'�� ⳡKB�wT�]9�~P4�l~�U#��� �ۘq��[q5l�ؐY�WT mv5 Wt-|����r��έ�<���ل��m��s�4���(6�nY0�vWI �0)r��-��-�%?�i��ٵG��;�����M��9��W�OgUP����? Jw�~�G��m���ꆠ��ng.*��W��19�]s%��f,���z�I�>'`���f%�F�����Y?Iz�U���K�r�h����c�����B2{�^�3�v��p���g�����z�!������\�nt?����#��}]��\!9�P/��[����i�V�{}8��Ƶ���|����r��.�6�m��կ��^�� ��L��
����|*���M���e�u���]D�;c�
{/��/z���_�{UTD�?#�M݋nd�ۙ�I냮]��7��OhOS�ѱ�[���l��KR6�NpWt�|�Kݲ�|���꤇J�̭ɧ��k��N��q�ۇ)��M�+3��I�8G*���A���N��W�r�q�y��c6��}�h*�_7�jhm�":a4Fv{j�JD��`�FiP>S�����]�Ϸ"��[$�[�Ɔ�u@�w/���uY_����"S�W�{͓�ʷ)�1p���\p .��{/�Ul#ױG����f������|*�@o��
�~�|��ՠjlB5"�)Ay�SY@!d�9�Mj���H9i� �������Sѹy��k��&�{{6�[�ϳv�&��Q�L�7��Ʃ���0�V�o-��tg-d0��rג�$�_��qj!!t�5n��s�ݠ���H�������Ki�65S$m4M�"�]B_.+.2jc��3]@}�w�HB:{�5W����8U��]J\y�N���gb� �w�k��'�2�gb �����c�W�^7�jhm����ۡ�z+��A�N��>/z=<��{�L�{Sv'���Fi��ܯB��/���i���ܙ�"�ҤN�Qsמ=;�b�9J՘M��y��_�3�\����w��9����[��V��x���\����69��ꮯ�o����c��	����lϣ�������zRN�r�W���7N;P&/gh��ZڼY�!�c�!("^���C�?L�rg|����6��!_sM*{�[�#�s�kc�� �ެrr��%��n<��y��k�`{r+ܩɳ�wB�"�����b=�|�{�Lc�vO �\���|�����U${kZ�v��^����}��\�#6���{��.���0�(M��Y���s�sUy<��
r���� [��@�z�ڻR�D_��V��j�n��P�Cn���`,콪�U���f���nA۰�|O�?s��=���Yq���a����x�����z5g���|�Mf7��{�Wl�?��R�<�on�	�����U�-����3J�<��"J��X����F Xn�.}ud.n}�./]�8�j�.�/��c�N_+]^øs��:�q�S9�l[�z;����G�nݫ!�=dkQǝ�K����c��dz��wZ��\���9�rs����˛I#n#ul؈��\��%�n���Ouy��������v��R3m٫q۷�k��:wcV���;U����z�a��q�{�ezǮs�}n�R�2�;�A��^fBB��&I?~�|������O�o�� �6��M�j�+���yt�$^t(�.��>�!���3��i������{y��폚'j�RYݛލΧ���K��Z�47.g�0���A�u�*�]�]��&lc���OU���xۏ�3�z'�j�f�Y�$����z�*��8��a��cض=�]�A4���!�??!68C����l�"ֻ�9�wۜ�_KO� �����t�Z�1Ȳ�9�}���+�( R08���U$P�0���,����z����v4��,����~~ӕ.j�_�����Y�B��=��f�[�D�����S�
�~j=h!���r�F������\-�:��D��s��ܗ����fg�~������-+��9K2G������pɁ�G�}7.��*vaV_���Cd8~*����ݪ��_c���w������sp�֫��C=�n�V�B>�?©�y����w���@�k����}�N�J��ܹ��¾Z�j��S��ޮ7tR������R�����׾��Ѱ�[}�k[�m��\�,�	�En��v�؜ߎ� I�ܪ�.�̉ GgC�6o;��>�̶�oЅ�?>�]�]�{x��Ғ�c�uU�3Aн��v�;����#��T~^�&��ɱ���{��>8{�(>s��т?f��{o�����̉E�+���!�p�ۚH�0��=����b�m�_ʐw��O��6�{��A�$���!^ұ� MJ]�s�{�Єc;����=~|8Q4:�(����$�ۛ��ͤje{�Q�<2[�b>�sS}W��Y�'��ɥ����z��O@݇t7��.����~����`C��0~��nbS=���`(i7��vi;ޜ[ɣ�4������'=9Ք�g���;�^P�А]d��lԩ�˙��bЏ��Ϊs5�]k�Y�A>�Ȕ�#���N�u*�u�]�����'ǭ��[�e�����.����vV�w#4Of�ѓS���"�����Ơn&e���f�$���b	�Κ����V��U�6"H͍�|_d'Ԯ�J�17^M�%#әԨE��!��0@WcO���J�����j�n���]��t��!���^���>@�yB�g:��U�_�_�G���D5=�s={ٶ�a��@	oM�P�}��wG~�편�;iT,���H���x��Gێ�v����p�4wF����5����j���'cu��O����M�(��}w��[��"�p{�B��8>��7S�X>Ȕ��6�����z&>�[L+����dJ=���y�)C��:s�3��Y��d�nWxk0�S��c���iۮG"n&��ܵ�˙�9NtÄ�W쭯�B�Ưa�
w�h�ߊ����Ҏ��nZ�\L�A�Ev�I�sp�S���.�� 5�t�:{�b݉^+}V�ظ�V�N�Ģ���lp���@$.��(�K�y�v���F, ǵ�I �{���x�5uG>���Şs���SX�"�+�Q��\�9@��ǢWT���Evm*U�_��G��D5?#uːB��i��P��dB�ʪ@=�H#�{ss���ߺ���\�7<�]N��L�4_��:��q���M�ya���p�]��m�W5%�����l�����o&�m�a N:J��32��W�ݻ:��ױq`�5�l�wB���1�c�t :7���Z+��,�V��;\[[���q���S�uͶW�a:گ\�8.ys�m�;=\���6z���j��m��cA��t1�Q�q4�+���V���a �ʘ���n�nI����]l�U�7�v�ҵ�fz[E��'ہV� @G=;U�\"k��p�_V��`�!�0S=�:d��z�����z�Y��5
�<�y�w_RN��}�ԗ�"2bc�N=׽N��I(]]�+`��Lhn\��aP��8�S��"<On�y�G���1P�ݼ�B�_���ot��Ϫ��M�5����/9߽�� Ww9@D�L�.�����;ә ���!I�zW���zs:Q��%߾���>({q'��ޕ")��bY��ӈ����s�R�V����!�p�۪_�NR>ח�]�Z���/ٕ��r <��1}u�{�B�Ьq��'8�~���K��ʸ� ���<��;V�sá�V�8�����.;�zϭ�H��� %�l�}�L�mw��$y�PLb��G��g�n�)�G��'�̷���i��3p΃��5n�|M���4L�w2l��.{jf���QY�m?{WY�u�)�Ǫsť3���۪��:�0> [�ҧ�<���uo��K�݋H�-�_����|y��s�r [���8����5^��%���o=�q	GS2�%�2����+�Ho#��͝�(\����U K}=��g���wf|�m��Xu)C�PBlq'��f��w"R,��/����@�̩�=��H;����x�c��w�������a%���R۞���{;� sgl�;�-��h+��YrNw����z5u�vӔ\����}=�?#k�Ͻ5��d��p#�����w�H�^�["CLy�{���k[��y�K(����mh���Ho���̧]��z��;z�W�!L�"I���vvee%@#	�@����>�ף%�l����fӚ��\��k�jבw���SܰBA�������{ͥ�]B��F��E3����7�e�x�p���X�%s.-�/F�kO��lC��]sܡE���zߧf���:{����>���>��.{��n��|���t����c��إ���W�U��r{�т��s�/YS�|�a�)�Ï)�ճ��/.
��%w�vƣDWץ�3sH��@�o��]�
�k�/�M؊i��/�H�Ln�;�Ʒ$݉}z�n>�/(�������59ޤ�nO)WՖ��7��}�1���f��LÝ�S|�xL������d�*����߁*�^�W�����:��w{-���yt5��y��g5��u����/{��5O��_l�M5Vk�v�JQq�d̞i�>�W���"���w׫�����5�7S�m^s��J�]o�w8�Y��UnL��d�{}�u�ǜ&�?n���*����Ǿ��C���|}�j�e��J��`��R��΁zr;�B�����`c���Mr�z�f���;�	�7~mT�Z�F�qsk�罚�,�7Z�d*�}��L�t��G��/K��L�3��{˃���z�|j��\0��Xq&g�/���?E�cQ]�w��
<��;�W���~�([�ؓ�i�x��㚹<w�KB�U�,�kl�ڵ��^�K&��,�������:#�G![��>%񼆿k����_�m~��G�Dޟ4<N�sD�#n�dE�ac`��`�O��!\QQ�DP��*�$�*����,��8.G",qrf"#G�X��r"0\q1B0E�8�HŌ$���સ�J��FG1#UQ�q\V0X�!"*D$dT�2`�E��c�6�,�qa1�X�X\\V�V,�$d���cU!5ɃdEF[qUqJ�1�I!$EA��H�TUH��2d�"HBH�20�I �d�"EQ`�1"��&"��d`���$�,�2,L"�"*�($I&(82@��Qc�!�U�a ��.F$a��"�f��	!"V�B��1$e�Ȣ�H�DE�.A!&(1��$�$#$�#��H��2H�F9 +&HL��
���2�)1� ��Q�B ��B"�E��b�EQ"H�E\QcW!0���ȒBF$0XC#DA����"�Bb����qQ�&ABD��2cm�Q��"
䐉!1��H��$"0rFHF8EcIL�c"F0H�*�#"���1� �>V�2��{!r��0ls?!��c�s�]��iM9E�u{IP��{"@>+����|D���ĭ�Jl�d1�)�'Y[�I|���K�d��5>��_�1�6	���>��rY��a�I���J>jС�`�hݷ����Ж;l�=q��=mn�^g���pf-C�#Л!�o*GƑ�� A{�*Nθ�-]Z���L������fD���cl�&�p�۪DwS�
ta�Uߙ�n�[���dvB�H��s��N?L��q�W��mj�1� �?�����w�=o�� ���NR�FwR���( ��hy���(�G�?.��e�j1���V �ܸ`���8 ���g�����r!�I9h{W?K� ��64���LV<ݠ�a��^}{��L����/O}�sn�ݯ�L5�6_1��g�g3E���3�]�z�T���aK�믒J!y���F�M�蚟���eD�s���}{5�+��t\�ڋ�����a �gC��3ؘ냡7��yX�q�,�6�1�6�����?5�9s2��9�wMBI+��P�Qo�j��oO�Fl��U��ٗ(AW��@]CI�Ĥ�m9�+�n�Ƥ�s����vm/VS��
�֤S�ڤ���5���6����2� ]U�[g�7p�����@	���@v/b�R���Y}�Q��׵H�^�[=��G�\K�����V!OL��$���F�c�Uxf��;��˟��}�<B�B��EQ��)Q�>��r[�J�G����k�S��,���B��s�<9�3	���M	���h�c�G9��N����X�kE���O]�� SaB~}��e��Df龸��QӜ^J�Q3t��2<i9O21�?IH��SD	�r9�N��UԌ���59�Ne�y�ۭ�Y�������u6�7]�3شq[s�jϰu���m;���9:�H���na�q�C�t��[;�x�ona;O�[��컬��9�ö��mU��v5�����"�j��{b�k�q�m�;m6�X�N�O�: ��2��<g�&99l��O����5�GvV����8ܮ�pml[�;JLn�<�W\۝�;oc�mY�s�;f�2��`��]6�L������I�Gm=�SnC�\�������X�,\�@J�n���*���f1��s2�A7p��u	BǦV�[vVԽkA|;}T�:;�,��=SȘ�u�}rJA��=�Ny��|	�q�@��+|V�O�C�^*@�d��W���!SZ��=	��n���x��kq9�����c�s�
�y�͜7�>����U|	V���=��G�$�t� ��rX�q������iR=�"
��(/�s�L��N"�>~P��<��Y�&�;�XL[n�bĽE�n:z�;�϶:����F*���Bc�r�
��R��E�c�7ΫL�����1���Kq��(q�2�����;�*����4B���1��J���Vi�Ys<ta@b+^��$��Z3o"��^��Ft�P��y�=���vҽ��d[n��6E~��wY�*>���"�yȁ_�ꌇ���lls�ю}��#̈m{��I�u� Ews�����c� A��� �y������7
B`p�[ڻ��_�/ݲB��<��!ofʟ�)�ezv��\�����ge����8g��p����N~	�r�Z����2��� >%��@��}�����y���{��i�@�Ab+h�Z�khSSHܓ.�K��ųk�7gk�y8�=v��>���͞��?6r3�9���~�V�eP{n#��0"���
�y�^�� ��|�o�lz^��;��%=������֤El�W�Ϻ3{!���x.In<6�B�=?�\��^�e}@̕p�{.��/ݓ��ε���=%
e>��ns�R��W�=щ~߇�U/�?E_fm�y��*Rʗw�;cY���U�| m�9>+g����s�dje�&�T���]r�}���:����E�fU �{B���t��e�F"w��e)p/B�N$�V�}@!On9E,��mҷYy_ s�*~��T�;�不��t�qqw&p�{9��*��,��Ża�X�=q۳�^�τ};bz��:^A#R�=���`�7��y��B��ܯ� '{�K|���e�Lb*.�� ��ɠ��E��?��͒��NA��ꉭ��c�չU�����"���>�9߭���������B0���g+� S}�A2��w}:N��W|�_V�P��=����-��N!B�Y/���>�/�-���	���� ���r Vo:�~�܉~ȯ[n&n�H��F��`���{U$���ϛ\����>�Lw9/tw�U�}�����5^�����'�}��ٯ��d�݃���23�R�u�4�O9��#�'�{��I���H[����Q۝����.�zs*����Rf�V�f�Y������gL�{ɼ<SE�f��#�B�L��I̖���y�lc5o1)M�g�N��շχ�V�mIb���{k��=���+7�I�D�Q�z��m(U�wT���j�dC=�ڙCu)��_%u��T�&�>��.��(�;�����"�s�s�7{{~��Q��!C��y�~=�n~�>/9����Bʝ��t��V��x��;����px���!��EQ��K�֏X:�|�QݎO���Jj������S{�T���u��Q-��N!B���u� E��U�D�3j��*#� >"�� Ggk� >��ꯐ�;/��*c�'��l�k����<_��m_f����w��թf>�jʞ�6�.lo������15���d򆩎`�����d�Ӿn��uu��;T�=X���x��c�"c���P��;n9��dP�ۈ�Ɓg�x��gMn��cS���!:ɣ;x<`��l�mgo!n��\V���ּ�>|��qu�Lw[�N9.%�[��ڦrY�/v6���Nc�n,S8�g�¦��xX	�7P9��t��ཛ����^�v��h6설�I��(��	��!7Q��LJt�H�k[m�=l���xmh�]�����RJ�G�x�H��\�A;���ws�H
˾�3�,q�Y:����jP}�P%R��!^z<4����T�y��vggu8,�n���*A��ꯁ=�{޾�Q{��N뗺C�����|G_9��{T!z<έ��srހ��D$
�/��@�j�8��4�6.ȧ�&7�m����MS������=�S�Y�i��W}X�"sp<B�C�����ڥHB��rux�c*�%
��T��׵_Oc��{��μ����7<���Ll=��n0�Pl��DK�OZӻ6�ݫkA��~���5�i�(P��eu9 ���٥�$Oc�r�9U�;z���^���A�וp�ۣZ�"S�sݢ�]|�����{����ǎ�hg���{��ۍ����̻Uk<��Z���ʗc�en]D)�շ!��8��Q�W�~���ȯ'�o����A�#�����q~��U�6�c���q�l��H@ן�!4���ܣ�N㟁���_U�G�%�߁V^Ut�9W/d8�����|�����t��vmuť	ef:H#3y����<��k��@�Z���P�l^l��۔����y>՗�ˋgR=;�*�=�P�����.��tާi71s�s�$ �s)�%�?/j9�j`�8N4���v��m4��Eۇ��|�}��vޅC@���u^�P�
�q� A��*~4#��y���Ҡ���jw��;t,��K-G���`V����C���|#�q� Ff��FJ��������=�5��%9naMB{�`$V�9�ʸܹ���B�WqWD���Լ�ٞ�/כ�xY
ׅ�'x^��ș��|3~�:�إ�k���0�J��b��f�����+�����p GNc���37��U(�R?�O�����&n�.}N~���ޕ(G�Y}[��츒�J�#����Z�C�kÇJ:��6���F�66�@�gd@���(��~�Ue�W�ok۹\�V��t-�-�^M��3�2��Ev=��±a�wc\��l�V��<�I;k ����kb���N����6�\�|Y}T��<#s<ɿn�:�\�gf��N� �#��&�-�ٜH��舫��0�ms�*��S��U�ԭK��Ξ���-ꙷ�F��܉��^q哲Պ�/���[c"�����a�^w9�
����>��@�G�E!��uf�aڷĀ�r� @�����l�:W53�H�u�]MWgNj8�pd=M�P+w�i2�Q5����s���sn�����+���N��3ё�S[�Z�s�_�X��l�{�@��ƍi��4�M?Z=�{4����Ҏ�lvTy9��An��*@���?�����<�:l��/#Q�-`컛&|�n��t\��Y����G��<h�|__�~2��:Qs��Ge�� -�ƣ�L{��Q�~".��(m�R�^Y-�i�����nPq���-�蘛����Ҥ	]�RZݚ�zo��3�)x���"��juH۽��
��2�7�yϧ:�G�ـ�n]�R]��%��Sm	���䥷�t{�~Uݔ��r�HQY���.��3:8Ȏy�(}�����Ǖ�^�P�5n�	����(B/v:}ʥ��V<����3(�:�7�Uy�/�O���3?����f�30�#�ffff�3̸�a�	C��({�J*��BP�P�9T%3?��033��032`fa����fa����f���fa����f���fa����f��@fa���3%��e5�O�} >kŘ ?�s2}p"!�\                     �                � �z��PH 
R� 
����@PQ �
(P  �*@� U D( ��� PQ P�                                    �         (�^�.N���9�[nn��.n�Ɔˀ�-�c��kK��X���vPʜ���� ꝲ�c�)8κ�P� Q�  Ώ��a9eA֬� nDQ��L���u\U���*�����n ��CrhT�GM˩�j��7�r@�AI�           z{
q�seN1�� �+�U'\�{�Oe�붫a��+m�qn�^���v����15@���$H��p   7��@� `  L�!��(rh"�M �  ;�
��P3aUA��� (��   p        � Ū d=��݀��� 4,�@,� �ت�` @A�m (  �   `���k��t�  C* �m
(�� �� Ů�l�G�\��wt��)V�- �           "���-K�QJ�҄�iT���BZ�)T�7 �J*���(\�
.f�70R��{��P)W�p ;P�����V����O 4�J    ��J�s4�B� U%BW���9���S�:@*� wP�� �l;�T��s2�jj��Q'��(@        �
�f���sn��Tr;�mY��]� �:-����P��GfR�nڦ&���h�� nQ!��6�'�
*���@uOy�N	rb�emp ��m���mn[��\��,�l� 8trnn�a[[���Z.`�1���� 5<�Ғ����S�%%T�@h2d0��zD�  Ob���I@ h5Oz��*UM4�&C	4�S� ji�h]���f=H��4�[B1#���P$�	&�O5����$���BC��IO�$ I?���$d D�ɪ���I�̫.��&��d@�&����`*��Qwv���ϷfO�i=����k=�u-՛Gǈ��JR���5�R0�����o4w5�흀�Sy�&�,o���έ�Ru㓁�N=��톌�7�o`�����kMƄ��,�/&8g��8�z�k��ϞQ�^gwG�7w���8Klp��x�5L.���$#��m����9؁�Kr��y�+�=�fZ,��F��u��oڣJ����%���Nŗp�\��(&�0Aa�t�j8�K�Н�#(Kɲn�q^q9�i=	dM�w6�\�'^6[$�6=�.]�u&&�ln���ηE�v�y��S��ٌL*6��k��5�m(��p楙��E6�Z:L�DsxÖmw�g`�K���:���4rwxHu��s$�*^�yBr�7,GC!�}΍BQ ����	r	�.L�!`��6���K���ɒ�3��ڳ�����V������<y ��e�����fr\ㅔ������g��J{k���~q�j2�ت�ЌN��f�=��蹼��n��YK��ɽ1��s4�NN�]:�.�r)�_��{��y�޽�0�14aB�-�'3	������j����o!����0�I�$5��*�}�u=τ�;5ѓa�Ѫ8w)�ZbSQ=�w���}/e{p^�N��&Û���L�a�]���΄���x���s�1�C�ˇj�%�;�����.��	��F���{���k���9B[.��ۇR�[cwI�X׈�#���c�W�\C�����<�}ۚo��M	��ǔc����B8{W3@kFiwan��d�)m_%�L�pv���!@��ǎҧa�teI0�t܀wm%q���w���X%I��t#yaxg �:%�о��*�d{���àɳ���B��P�X��ԛ��V&1\Zv6�� ��׷���FPށ�z�[��Y�-���'��6�:mM���y�y+O���{L/RMC�/k��Bwf[�-o.?�,9!�K�Gt;����jw7cfq�&�|����>����U#"�2lG�+Y$�|~=��M��2���E������'�߽��k=�z�4��'B�U��O���b����0�4.���˺	�j�5<�)�;T�ɱ���@=#w�Pw�k:��˵����Po+���� Ĕ�6Ė�F��y]����`j��w����}�(�y�`o>d�D���	NovX>��N[�6	�f�G�y�9�US�ȺrC7�V��x�6�dL&�x�wwjk7�}���Ɯ�.���c
�I�`qkr�����Q�������2�𾯦;����Ap�n���tt�ǎS��<����4��u w���E��{H�^^р\G9�؝Y�Ȧ��Թbނ�#��B^hlY�	��b/>:���F�[Jhq={ov�20�$����.�����.�{�i�:�J�*fc/��c�_n��؋=`a�&�9��X�fO,�xU;�+C��2*�Wvٺ�td
�$c(�;�*)��0�3zb�;A�ݛ��qK��ߨ��v�!�a�Wn�N�`�A9�S94�]e�Wn7�lԲ!���)#���WC=ё'����ʓ7R���-iZs���8�$�f�S�u���k��>��9s�l70����v���~ݒY��MɹaG^ȷ��8p/��x<%���[w�6��p I8Re�HV>��N�n���e�6�5P4[r
0Q1nN3�7 ��y��
3v��Iα֬��!��4�%nki9i�s>�Lx�۫�Ǎ������[$�N�%�5l&]��{�jۘA��:�˦��)$����΃��ء�w	6��a2W�-rR�a�U�;a$���}�u�%ͧ7�S�r�]v\��A��e����G Z�9�]͡t�@�ưbO�<\g�3���C�/�$�Ɣur�K r�#�Un�B#P�\�  ͦa�oEza8�v!�N-{�VN�dH���}�v�2Y��l.,�5VJF�Vh��ۏ������J�
�[!�Ll��ҍ�]s�1t�d�R��!̌�I�e0�R�oP��b���B��-!��w>���M�v���E��z(��E�U��|[�\Yf,*����*P[Ӥ��{x�aٛǦ�\KOd�Ӝ��}�Xd��v�-���}�ãܭ7����sQ�J	�O�bq=;l��t}4s�;��� U�>1q�}.��zQ�����r�F�r��V�8��q.��[-���ڰ�-kS*�gj9��90��һ�����y��ۿR7O-�#�38;ѳ�d��c�i��R�a��@3"�vB:����`�t�y���iO�N@
�sGb���gE.��Y���?�q�?w��yG����,�Li�c�q{���	ɉ�ڔC6��`i%��sb��S��s��Η�dy�� �r�Y���vh���k�����2�+�q��ص��1/u�p�z$֒ƫ�nht�\q�:�d/��X�V� c�v郑졋�,���i�{̭�d�[z�z�2Z��sP�b���ܛI���e,�b�����7�:cq4y"��%_>=�x��ع�˱��s|�Fۦ��8ZY-���κ�ˎL�����$����m���
N�C,�-�%Mc o^�>fѝ�k���+q8��J�m��*>�t��������*= ۺ�u�����@���N��ѝݗnHK�����Tqo7�gr�Ow��n�c)r�u�7��46^fō�����8��	gy��q���V��t�,��jB�ݕ��,��Ng=;r��ܔ}V�m��J����d�[f-�j1E�$wUK����mL'�S��wW�hm)�1.��sTm7��h�Ǧr���ۑ�}�k�}wM�t´|<��R��˴������7/aOPb��:+���݁�\Dq�m���]����%�r�iѷ�� ��cE�����p�r-͙n�
�Y�,+�ɨQu�4s$�C�zgO�}����rc�]���8��j���F�7�:2`�-���y��v�5�9/݆D��Ra��gS�z�e�Վ���eN��Cv`�lnp4m�l{�v�1hf$N��5���,�eͿr�Ƿ��=��c���l��;y.�Ʈ��i�f���gb�b,�t=r���./�rMP��N�����K��pi���Ȝ��v3Joiٖ�F��z5"Zt��ݲq�m�uv[��ł+�V
�yv�3��mr5N�-ٝèJP��7V�}���Y^��1f�f�z���-��.�՝������6$��C�s���޻�{s�����-5��nI�<�[d�{�#�tǰ)�T`��}eWU�n໛u�X.i��f-�wd�a�W�4=�n��{�%ܢ<a�)�MFa}��,�W|Bԙ\��{n�ĕ{�˦հ��w]�cݏA��` �/w_��t�yM�l�y0Pc?"c���z�aIs�v*��f^��q��Cv65�q�-x��Ԧ����F����%�]�E�~�yϦ��\rh�I���Szb�����.r������{�ۅ��kvL�@
��ΊP������+wF]����fjĞҊ;�Z�X �Ϸz
��9J�è��æ��[z�\{VOK0r5n����t���ժ*�=��B4������f��]�u��ۉ��/!��Y��Y/v��[]�'J.�V\��>��m��,�Mmu�<!�1��}�FA�Dfتg�bG�v��T���jP��0
=�Oh�9�:1�y��y����yd���L�Y��q��Vy¡=Jy�a:��{a"�)	{�`l ��v>��;V�S�r��{ݥW���ͷ.��Z�aq������������a[X�����[�oY8����q��]��5wv�U����1�{6�r=�����D)��lWL(�}�;��i�+�X�^Uц!S�`e�[~�Л��-�M��-(�:��c��M�"��=�%Ǻ4�J�6��Of�j��x��8h���ܝ�*QM��ntL�R��Sk�n��qӒ��E�5ˁ,�nF��)C�L|��ƭ�o�&�3��p��֮���lR�#܁��Ӄx���٦lSOG9n�]�M�z�݄pL
ň���_�|��dk��J�<��}csk1�~�L\�Ѽ�x�w�/�[��a�C��ܫ����u�v"C�\���yD!Z�N7��rm��m���� ��n��(�f�E��0o�\�&����*��<0c�a� �N�e�׳�ѴL
<y��n�{�9q��.Ԯ��[�Ս��YَY�jRA�L���j&j�l��vvS:䏃��&ܠ�&�r�n 'mܦS/fQ٥A��Cx��鉈�!�+O�bp.�jÜ�Nk���7�i����� 2��菈8���t�0P�}eQ��'n.�z�)�����L�Wp��{��8�×x�U'�p]&�h&� X|l1=Ĵr�ɝz�䙓�[�sFj�;Ж�b���|��Ӯ2�#YGnnu݋=���(�۶
�b]/X�W���cuκ��=Iq��X���P����K�3s^��J�����������$�ΘD��Jؒ`@��v(��8��ƣ���[���E���݈� yT�%]n�Iv�4>39ZD�(T&Ұ�v#�ct>Xu��$�F�uilN�=�wy6�Ru����Чj E���� T�hi7�^d����v�S�r���]9��L�E�M����t���l����WdX���|�8�[l���7���q4��M<�_
&=�
�^��#N�{����۩����*�/I��4�Ǹ
�ج~�D��9 �7:����,_W����$��cS(8���`�lU4�'��z��s�U��1��q�m�D�G���X��̻�c��#�/::����hհ`w���ˎ$��^��c��䋁G�`s���u�T۹�F�I䖹f��Z�
�a%N�+���H������%�]�q�-�(��%0r]ɦ�d:2UgRgg.*���Ō�k���Du�ֻr�"]�Zӂ�j��c�s����;���G��=�@�3l���3�����ń=�+m�N�uv�:���(t���M�g��Nv���`8'>Q�KH�8��ӹbm�G�u.ֶeKF����t_?c��/ds����&��4�CF��&io�F�S���o<�KW�nU��y��7�T{\	1k��e'5=Yq'hc��Hq��Ӎv�ۇ�N	�[���l�e6�<��9�:Z�ak�flPv-���7�B��\J�����G(aԭ7w[��A�0V	�9�/�]�y�����qq���G$�8&1/qŽ[𻓖�
�b����
q�)'Z1�p��&�u.�[9*�O����ͪ�;�����x�0u�������μ���%�u�f�ĉ��/w_q�.$2��=�R�K�pW����s���t��x���u(v���OC�ώҕ�Gwck�ۍ���`�� ;vǶ4����Rڢӗe�8�5��;�G^�e�;�в��;l8���Mԙ:_])��wm�3�ex r���AG��d�f��>�1��k��?6�}}���]�&�E�a�)�z�Q�|���)�=:䆄�Z�Q����&1��>���F%nlQA�5^��5�e��ڌ��.qW�n�M�����2ܦ8�j�9u�ˮs��}�qC�;��nvY8� (=FgN�O
�Z�曫h*�P��G�]�td�Χ��Y��<��q�֖��)x��O�n���x���2ghTB�8�Q�%��u;����8���H�y^e+7v�s�u,߂���*�����踩��S�V˅Gai����AօJ!�4^&J�f�#�b6�՛ۖ�2�pէIO���@p�
^rB�N�NUKVlިrq����.P�U�O=�>�;D%m�p�7��̻zM�5� �`�N����
eWe��˶� ��.b�i���M��u�u.��^��- r����v)�0��{�΋&��ZJ�R���2�7��yAG`Cyh��bÑM�sy���{5b���Sl��P/g8
)eX�c'����N�H���<���p᭜CK����:f�Ǽ[��O-ˣ1cm���C5��p�8�I�T�.��\���^E:<����S*��7nZwB�آ�v�Gulν��]a�p��_Y����q)�}f,���/&��	Q�3]t�4�uN=��+�٧Y�l}�7o:���N���M<Y�b}0f�I�ػ��fY���	�4�
G�z�c��c�+�q朹�;��7�g\�52ν�lS~��Ya�Xc�iG��$L�3���5��=��U��ٽRŽȃ���3v�iXɑ��F[옸�P>� ���[Q\M��w&�0�m���tv����-`Ӫ��� ��Ѣi��D�(�Zz��/>WH�iY�4N�J�p�(���N�]݉ccM�5��7��/f���J���c|ޓ&����C��׶��syc����,ڱ�om��j�f��ʲ��ǽ�F�������Iz� � �, ��H,��(V@�������ABI+! J2$XH(��P��BB� T�$�,	$X@��XABH		Y!�, ��VHX@H ��,!I $� �B+B�a
d�!!*I�"�,��,��T!�T��T(A@��+$"°�
�$���*"��a 

�B  �a �BH$(I�I"�H��H@XH�(@XA@V B�
@$RB�	Y! (I�� � �$T�`H�B����HB, VI+�� BBO�HB!!�P$�"�^���ə�ȉcHuD�v�u���������6�u �0��8�^�+^��޾:���y�6��éJ�����I����I��)�j�<��K���9e^s��m�lחy��X[w̞c�i��S���؅'PCj��y��P�Dj!��[�0��'vf�І-��q.XgO{ǣ4�;O�6�N�4�qo+���f���ggDGR�,��=���c�=7[�p�d�/2=�R�>�nsu���q{�?ʤ�p���s��1����дD�܊{j���n�ŗ�u�|�ی�cU,ll2��6�9"T*�F�F��F�4�`;��˕��W����ls��[b�D�Ȼ���7|�=���������%�|6�-�h	�}��	�ѫ�Q~��OG�)�,{��2��:c��������]����۝|�|�~Ź��/�{��G�4��MݰЩ��D!)�sS�tǾ�p�~ɉ����A@7wM�6��M?�����ˉ{f�5�R�Tsc��#�,Q�.۷��d��yzf���/vz�6
���z���M��F�oNc'<�n�x�Y�~ӧ�.�W�����N��If�,9�,V]�t5�(��<��K�omh�`����>��}������q���nQ���(=��;�k�/�� ��yhz�1�s����1�|��'��T�Ϻ#�݋�X�UL3;�N{�Y�y�k�o�]�KԺ�L>葿o�i�I1���l*��w�A�ݞ�����od}<���77���^\��#���rrZ�ǎcb��>Ѳ)e�[D��x"۹�w�z�����SW�K���0�/���斟C�q^�S',c[��Ɲ��O���-���Ǣ�|�@�%k{L!�K�ؖ�ބ�v��_b���x�&j�����a�]���i���j36��In�	J��N�ɫlhcI��˜�EQ��c;���͝�]9�����)<��s�xNS�pKۢӻ�9�:�~��#�v�NK�qa��63c8Ok,��/'-�~�X����l bg�����z������J�s<��=�n�|Ԃ]��w�l���0�}��2�Ӝ���Ϯ��n��=�oO>��t��ꝇ�=Y�n5��i���>>��|������|Ȁ#ub",Y�>7��o��\��Z�:F��lٸ��o��>谈�u��8=sOI�B���=��)��7�e+��W�ĥ��n�on?xj�O���!��p��wB�v��q2Ι��z$=y_`\y{��W�|�ɷ$%0/g{^�d�����M�QbMVN�%8j���&�J�2���v3��{oZ�^��Mh�����~^p=�w�jۇۏWF�u�x��KŘ��é�P�]�^i�IȔ����}���9A����E��ًw�w/���Ň��	�3���#�:�U�ڕ,�y~![�Ǌ�ɫȺ�l���޷μ������R�|��ɍ��0���斦������kZ�v\⇏�P����>��f{[�=}�w�����iWxr�0���<g�ǃ��� ���B�����<tD��}��%�L8�xm��o$��|�g��·��B�A|��z3����]��E�~���uCr�%�٪��<}N���+�	�}��������h/s�.���Օ�3�������V�Ǐ���y��϶<�}I�{��I=ۉv�!<֔Va�;�d h�`�7�t���p�����Qo�бn򴵗�_�ڱD����	�Ǯ��
���YBRlǤ��a�*ǧ��0{���+�^˷�8j>w�[�ts˔hu��w�S�p�i��֯���O��/n�g�Q���h�z��=�uv�]!f���I�2�e����t.���cjb5�I��\�_�*gy����ǯ�~x�9V��ֻ��U!��[3�#h�w�m����q!}�,C�y��<���\�Jn�A�Ϸy_[�[p���Bk�x{��5I��q��Ķ��-�3��s�a��[!26ٍ][��'^\�^���؍<���鴬�S�T�n��뇡����fK�	rY�x�t��Eڎ��v�]�{V�r�o���Za�U������従���ם�k~E��v�'J(�NOyĆ�d<ٺ4�{s��5J�B����=�������ݝ3޾� Z��e��!���r�%��s�y���ra��2byO��z�Q�K(���Ul�k���P�O�7��{��7 ������5A�]Y�T���M�:6.�f�R�l2^&hY�5�Mb++f�j��Ş�F���~�m0�H�ۑb�@�|t���Ct�"�\��˵�܍v���D����4{W����UC�O0�G�u,� u:cs!�!2i�9*'�ރ�I���D���i��>�'I�\�c��T ��"���8xt+ؠ��5nn��ڽ���ۇɧ�BaaY�ʇ"�u@l+ʁ`��u��p�2�K�W��q�nv/z�W����}�k�}vbI.Iw�o����v��o�mZ�u�º[��o���w���
��_i !t�k�xy&��	�;�34�3�'[�bf!��{��1����K�>��m�˄"E��U�rT�d�g�d�^w����3+t����6:��C"�6vѪ�Ca��j�4�nUP�N3G���@��M�g��>�y������
;�������=�˴�\ν��SLrk�B��{��q���P]��P�L����r�6�>/^�h�<�����p�ۃodK}�������lh�Vt�㤧'\�͉�X�t)u��*��7�y���|h�wfo����l��7�G��Vy�`tJ�Ky`Y����H�;ϲ���4�Պ����d$��I�47t]$��R*q���:�1E����2�IvM�0��:�F��\�#c��#�x�X��wm9��|���b��sF�^���N�ڋ���EK�l��s�;M<�꠾gپ]wf�av������Y�%��->��|7�gq�\��F�p��5�Pݰ�ᚵ��El]��դbE�;���2{�Qk��Z����e>�7����x{5vh��;Ǫ�5��F@�y��\S��0�TݣN�,��y�>ݜax��h%N��~9<� �پƟ-ۧQ^�A�:��P���p�x�+���2h�!���x����y��>�H�`��l]��dg[��!��9�{�y���'ol	��{���k~=l��%+�n�z�W��U,)�� ��փ���7z�;���#|$ ge�G�v�ڽ���|�=�'�U�
/��Ӟ��K}�-ulf����_�؟��G�U����I���sK�~�P�go��N��%�Ԟ�ܮB��˱U��yE�C�������gm���k��n�;�OI`�٢����p>w�O��7�s��`��7��ΐLX��n<�k�}rwc')��1u��`�^w�io�@����No�'���z�zX�I���O���X��'��ȅw5�f������B�tD��/�"�Vn����{���t�1��1��˯쾈�շ�c���{�@Ň����=���3e�v�װ:��Јg��A�v� ���u���L(��zy8�e��c�yz?(�r��n��w�/������F�nm�i/|��$�̊W�r�X��Y;���"Xp���n���{��=]�6��Y��ᝳ�@�CK�y2;d��_��%a�8�a�5���Kۋ.P�;�[���N�%
n���:�8����n��Yr��o]�%�O��}L�,�M���-��k�[�/5�"�n��3G���k{�P�{���Pu�ed{o"�/sr���(�n��J�oݳ�=!u߻��;V*v�#�&��x�n���x�{8M��Or�cG�_м�^�l�m�Y�����c�DQ�
�>��pbí�r÷FdA��w%�ج��^K~ҫޞ0<��G��w�-,��(����ؕ�.��|�Ǔ�D��� ��:JF��k����a;��Vi���%�~�n�{V���&Q��85�j-�R]�o0C�(�k��l�Ҍ'h��b�ݬr���
���Gu�Ӭ��T���pW����T%#ў�#���4/QK+��g-�����b��W���{Ϣ�i2y�|�*B��u�7D�e�g���>{��S��{�������������<�N9��;�ރW/n���t.^�������y*�vn����%��еLU�tرWK]a��~�=�:�Gy����p.��S��&��%o��gyv��mO�I���2�LL�ٺ���.�ǖ��)~K����D�Y6
�`��Oޔ��Nn�����yݯw�.S'��Z ���zࣗ�y�F�w�_��f�u�]��o��?x'ݡ�J�ǯ,}yl4��HǼ���/H��V���>c�:T��)؀J�,��qǛ�����LL[��3�lx�"��^{pl����Vvჭ�v)����۝�U��fso�{��y(�8�j��Wi�P�>��o����Da˄O �.���![/�[�fN;"x@�yan��EK�Q�J����v\8^�Z���g��B1!�}N����:)�EC��G2���P����(�H�;�/��3ˎ�7;j�v0v��ƾ͸�{��wؤ���������:�i8�Fog���(]�j�W
�t���ɻ��a
o��ua�{M����x��(�ڽ�%���wp���������#,�k�͜/���lv��/X/�ܞ��\�H�2�� `eFO��	�x|�t��+䁴��'���\��@���x�O{��Wvn�:�&�u�2�9ٽ����u^��P�������*�-����9�\h���@��x�#}�8x�$��C{�W�Oz������<"���2#�f�f���e]�W�p`�קk+��2^�Y�ˉ޸g-ɩ����Ǝ���[2�aT�j���,�h���Yj�׻6�x�U8-�d��2p#q�O�4�ϩ���^y�"^�{�f������|3��z1�N�,�9��y�z��2�Ж�t�y-i��;,�XZ������:�U3�n��)��K�N��_��&���nn���Us��ٳBo�6��3�G����Eث���fs7���������2��c���H��x�֠7���T����:���(<�a�Ι]�GE[���芙�]!K�l��}����zA�{�d"@MNv�q7|M;u�Da�s�j�mD�h��څ;�'���L�=�:<=.�LX�su�l�OWro��41�}��iU��S�⡈�&�R�c;�R�����'f���wU��7��G�+9��.��o�U{w6���Y}����O�ڷ���ly���H4��5���彺ы�;q�T���sۡP�Q�����p��|h^�f�9فwZ0��8<vFbQ�Onh�z�dy�͆��`�W��2�� �C�xi���n���>�f�7�V�Y7���g%�y��m"8��;�4U�RL�Mۊ~n���u���+���P���E���{�j����xc�n���n�������Ao�h�W��ۈC��\�B���D�]M�������:K��%�C&�����|�~�&׷V8)�vP5[+"P���L�kn!j{��7�A�W9Ү(y4�)����Mu����U��8HY���^���X���э�(O��D]^"n�e3F�m ΄��S
��y�.ǹ�l��NWX=%��n��7�IO�#��u��ջ|���K�5�/��/���� 铡�->����7�z�����$��=�8�����x����b�('	:���D��QU���v1b���G�ކ��w�L��5�����OU��7x<F��>O�8����R��h;���үg���7,*x�ռB;�^���{���~]�>hc�y��б���Z�6j����3J�~��h?�l���FU.�n�,����s��i�5���۾v�Oʍdn�=��80�:)��r3;L;���#瀓,�k�������U$�1豊�*�*�zy�t�gd��_��8�9v�K��}�u��sR���e�-Y/��4�ǎ�_Z���1��Q_����\5��s�j�[�3�;��gI{�cZ�0���H8jY��[��:{/�i�l1A��s����m��~��އ��\2�������^tмy��x��J7��I�G�o��٫����g+x;��A���}W��u&kaP����
�b�q�ֲ]��rn�B�l�q���7olat�������<"�N���A��l�=u�"]�7��,}���;ݞ> Ǻ���<G�����*�(^��oG�P��7GVc5j�fn���y^}�ۥ\Z^=����]��(�óJu�F�Q�|=Wy���8�e1�_�G�C�ث��#1�Ѳ�iY"!eN�/HuM�"�����.�{4=�_P�ܟ��n�]3�B)*��i�#��)vn;!2+�u�Ώ��d����n�2��/���t{����GܪO���+��k������K���rE&�o��L��?��q�9�~Wy��>}ޗ��V����Y����b$�<Z�.��A�KT��vD[��-Ǩ+�sB7ZԨzY��|VUnw-��LE��uB�����D�^��1yx��^��˒�'��>�ܧ���O��Բl�d�
�Ƚ*�%�o��=��ڧ��y�}�C�ܳ�sG����uE��L�{��/ݸP�Y瞏)sq���ڞ ��]"�����Xy8�t�ԭU�ҩ�mc�R�EEb��<���=�}���{��|ݯ6D�z�s���W�κq��:��r�nx���t�0�p�A[�]��ʶ�n5���]wdT�,h��5���K��bym/�9�p��]q8��n;v�p�u�$���q�]�����F�f��-�=�c=q�ѭ�wk��׏oWi;g�C��;�u��j}���YZ���Ct!���r��ɹ�{;yא�s��=S��l�t��ݲc��9��<`�oj0��Wn^��=n{	���Q;�ɺ��Gf۶x-�g�}s8ln�0Ϸ�c��K��ql��n�����G:{ěӌC8�K`���kgi���v���ዸ�6���M.}<�s�M�o[�wMcc��VLsݳ���ً9^3�^v{G�\����y]n�{k�dF�=�ne磚vKvٷ�8��u�D֓��T��];�N.8�U�b�U�\�ǅM�Or��cG]�C���3�u����&8ɶ���f��.�Q��;�`fLv.���'[��c��me�jw�c��n�'d�}�v4&�:4��r�ܚ�nhP�mc�]'q̆�M���n���gzά�8�V:�λHs�;rkc���q���<�3��un��X�1�3��N#�ؼZ�6-��D�66M�[Ϸk���W%��ӷA�.���]�nݫ����;n-����]���+�l�pӹ뷷pg�t'�B�^7,x;
u\���U����wqϜ��)۞�l6vv<u���݇��VYq� G1��b���
�ai�=t���>U6�v�a�q8��E�ZN6q(B�c����]���;agFqVۇ���1��ݺV�a���;=D���k�v�=�u�m�ʂ�A��=���Τ�e�u�rUgE2G:`�G;�v�3:q�8ܵƅ���tMr]Z3ܷLu��i����\���Nm�든Ì��ł�ȡ�v�)��nrI�vr1��7g�z�ۆ�+�dڝ�یt`n��[9�l����Fn�d��K�k��㤝���lX*���;FK����w�&�3���dWi�<�W;���Y�0�Pr7	�uW�FH�t¹��d%w&[\t;�ڛ\k�[C�iK���i#��ۅ����r��2[85s��u���9�\q��Ρ��� ��<zqnk�1�d3&z*{`8®d*mt�������������7d�v��wQX-�õ�L�a�{q���$Ӻ=�nK��]Oh7\lɻ[��)�}+��:�\6{n{v�z����C�ۄ��lF�<�c�ɭ,:0��[��^9�y1ۮ���P������ܐq��gs�nظ�˶�Z㋃q�qۢ��36���7spvG�,8��+���GK�l���������n�p[��<�ݱz����7m���뮤z��v������m��x�@[���/D�ݺ��v�Y��:��<=��y�]����HSc��<�V�瓮�m�CΣ�M�>;{K̮3���;t����F8�v'�ΑY�7]�5�]�<���[�8}��ཷ[��r�Ź��ւ�<��d݊2�Ń�2-<9��V�[�t�9%K[]���W��7=������:���\�¬v���R��6�kی84�LUŲ��ޝ��9c�9:��zs��޹�'kn��J�m��Cϓ���,�֓�ݭ�`ևv���x
Ӹ�LK>��67n��)ٺf�ݛ{nG�sĚ���㵵�m���|��[�]%ێP;��<\l󶻐vvչ���m��^���vЖ�N��բ8J��Oh1
q�.���n[���0���y$K�Z��љ8/Y��=u�V�ڹ���8����V[b�0�g���p�ln0�[�m�Gk�f�{kh�yۀ1�9Ngkyջ=9�n��5a�[Lq��ڝ�h�����1�䎝����6�utQ�Lv�rv6r�:j�n�!Lc��)n��m��k���!�����5���
qt�p&�G��Ocv�n�v�C����E��{���vy�y��^	���{\9�sl`��+�=Z�}fݏ#sv��1Ȧ�`��9��d(:�nڋN\�<�n�]ڕ�1�9��C��p�N�pc�0��ۮ�R�'��'����:�:v���ͻ��d�K�K��u��=n�F�n��4u��hh��k���I���Z��U�+cn۬[q�Dܴ�؞cͷ ��fM�-��8�r�sg�n�w'v�����h|=�ζ�g����-n�v�D�������x�#�Ws�HhNi8�-�m���U�Vm�Rx�w>����9�z�f;n;3��������x^�i��z�%x���dA�R��q��d��q��5���;S��:+��s۳�.���hӻ9��i\��j��ۣ9��Ƕz��5�t�Wع�ma ��m.����u�ڣ��OR�́nK��מ
{�9e.v��v۩'�q�p��˧tQ�ݑwn���Wc���(��bɹ�;Uؼ�9{m��x��΢7�M���&N�ȝ�o;O��y.t�xL�����`����)�S!��p�\;�-�S�����,�v�:���{N88��m�6���]sf��_Q��l����\6��A�C3�s�hɴu��A=�u���#�����ðI�d�6��U�ŵ�q��m��Er�G �� �r��t���9��o<g�|�`�	�oG�������ѵ3��tE�+����jx׎�/b�fG ���.�4v�>,�K��c�=��w5�}ۋ��8��wh6n,�<�0��ZP�=<��WY[��8L^�q[��b��<��qGW�C��ފM�vSq�p��Џ%�U�0.�6�n*ۇ�/�\���C��{&r����v3n\f�Żl�r/t���Z����P�����3A�to$q{v��s�u�y#{H����)�qg�=�9s���O
�t�GLp[{�iڎٔ�e�[Tr�l��p�a���-<v�췣Z�s��y�g���;a27.����e�+�^�������m����M��=u��d	{S=]��ApnŶ���<R�ti<6��H��W�X�����N#"p�q�+\!�����Ybkj�c.k�r�#������S4�U�Y�Y�q���rd������pQk���_<�v3�Ϸk��C�kϨ�rY���=p��m�e�V]9箅݋Q�s{Z��Uڒ���Ԯ��m�ʰ�ShN�\�۶\3��G�z��u�f$6�� ���.�[�Q�]\pw5ӳ�=��l])�Av�ݶ3��];f|Bu�I�˻FL��v�n�5o\�kȅh뮌�8G����706]���1=v��}�{v6�خ*�u-��U�Xۡ淮*	�����I�ͼuBcs��[R\i�u�|*F���c�xɴ"����s�vti��Y����n�:�ǩ��׫n��%&ݧiVw<�`�뱽�ɭ��^�����ů;	s�yM�mq-p]�y��r��<mF2@=�m�����8z�����%V��m�Wj6n����G�c:����"��6�����6X-3��<�Ytf��L��/��y�X4 �;G(�u�n{���|��7DY7��\��׳�&��T��Y�^Gl��8�7m��P<�El㞻h�n�Ȣp/l�kPx��7V�; -tV�@�q���ƴ<�D�Hs�cl]q�}�m����0�p�C���¡ۀ1���O;3s�c9�M�]�r�v2��B�Z�n�g�؝�F�۴7m=�H�6\�;	�kn�N�3�.=ۭzv�l����G�^۵kۮ�q�m�7\����**�1��-��{N{8��S< =q�g�ڞ�]�^�����s�i�7[K��˱��9�� ��y�cn���Eu�F�Q�m;�vhH7^e�NZ���౸�J�7vWi�[C�r�p���8:G����`��"Rs��#�o�n@=;���]�s,O'v۶�ɝ����ݸ��m�F�����*C�]e�a�&y���]1k�OY���D3;vp''�vFh�v۰�#]�q�v#�x��v�Ϸ�nk�U�ȭ��8�f�1�l��ۉ�����Cў.�az�']���ֱ��� �.���>Ǘp�׳#ؙ���f�kg�e�v�O���n���j�k�vT�pշ�����C���ݼ����t�ڭ��m�CA�h��F���97�v5�n�NZqg��&�#m�7i�H�N�jl��{*���{Lk����n%DދjʚN��s:zϻH�&=����wbۭh=ۓ��жݐ;�j��n�V���s�;���g��pn��Wb��r	�E���������8�.�<geM\��N7��#��ڻ�pp�Z�s�ݣ]��^��b�^ݰ����x�>�,����5�;�L��#�]�=>��uڶ[�+��g���ݶ�[�F��Cpn+����)�������;$�\�7^nݡk��>��C٧��iص9E��#a�<�lI����o<��za�@e�f����t�-ۂ#t�j\�xḇ8#�۞�!!�EՐ�mY�l���
i�[����ź��n���@㫻U���
�n�Ӷ뮹��۸���U���װ�\����.�V���a�� 6�c����v[�wn��l+m�GG)t公\ {b��{^u�y���7�Շ��"�&��W	nw.�]k��,6÷-�\F�
FϞ}gt�/m�[uz���'�we�Fݹ��u�.��v'�v{&-�n�u��FKJ q\wEp1[�уX�7n��v펴�F�q̆�'vn�x9���.�I�qh�kj�bۋ�==[:y����+m;�lN���nz�[�Vx�:��\f��[l-VrZێ��m��͙�8j2ݧk�.ڪ�Y���z讧��um��mSz�b��s�η<X=���E�ۛ�Z�v�ٯ#�8����g��m(�J"�+PZ��Ne"�cZ��F���e�Q�,4ܢхJ�Դ��ˉ����p�J����r�5�����K�Ze*GT��0�q�0jk.E����R�4����Ds0�V҅���r�e����j]Z3
k1�c\�F���UQˍf
�Q��C2��mC-�ť2�1Ձ��QEҍcn52"�V��QY�M4�U�̚sYEr�+1
�+P��ڊ�L�`�b�q�4B���ҥ�Uˎ���)��Օ1�-2�0SH������-l�J��(�j�*,X���DF�J���6�[h������-3)������K\jZfJ�n�Y����c1
*"0�Uh��,Z0t�J�t�W�Q�(��mU��։�jʒ�Im�V�m��b�����,�KE����m�����ب��J��X�1�$�h��5�ӱ�敹Su�q�%m�(���{n����� �=�8�k���}w׾����Ǧ��N���s���S��	��61Ň�6�����a0�ֵ�q���s�<r�SY��{v�;M)�������X��7���O8B.{�������3�Ě+եݳq�áT�득�s�<7e\�Oq�s�K��[[Y���פq%�;w;�ol�y�QЙލ�M��Sk�c��3��q-`y��q�3�-�g[��e&���ϧ�c�8;:Ŏ�ݷ<�c��N�޻g�R����kl��X��n�Y��kKn;5��㛎���;h+WO�y�ܡm�D�d��I��ge��z3�|�n�ly�y�9뭲JƷg^k��G:��z�'N�;���&��-���� o%������קw,�v�cH��8<6����-�=��Wp��-����v���nD�2a��7�s9�-Q�=�:�۝�:�ͬu�^��!1b���IΧ1X�%��Y�O�>��ؾ��8�vˍ=dz8���K���0�_+�Yک�������ٍ�d�GE��A�y����� ��"iyx.GlW����m�;u���9u=��ۮ�gm�8�њ�j3հ�[b�.b�ɸ�x��n����t�%7������D�]���gX�pq�vp�q�D�8֞�C������4��GU�����m�q�q\�,'����ͷ:y�l)�א�3��vr�q��qȡpt���˪|k�ݫ[Ӣ�@�
�7X�<��j��lh=���|�UN�x��-��'��۶l������nͻ�Ǜm�ѫw�\���rn�8������۱u� �m�rC۲s�`�ԫ�F���;�L��#�{u%���S��s�;t�z\��4��(&�n;�_[f.��'mm!֍�]:.�������%��6ĉ��t�n�kn6u�>9xΌ��S�q�շ>�p&�WBN:��UY�i멬�f�6�G��}^���}q�}q��@���G<
;rl��vr#���l8ܯ��QGr�2c��*&�����n9���r=�lc��s�˄�rq����9s�M�y�xy�8^<wnQxN{m�9�xC��`s�cs�wg�^r��s��6�p)��8��vܸv�6������\��siC`˔0�y�;g���v78T;d]Á�^�o�����=Y5�������� >�;��� �shv�U7���F�������k��a�6��d'�i5��l�L�{�߄�3��u���ϰ ��nS` 0�k��'��1��=lbBd�`LD��cAY歀|����3��:���(��}� V�?��,=��!�c
�SDI*Fά�dhεu9��D��vZ�D�5��I�$�^�d��rL�]����s~�z�ag�T��LE��{�C�{��U���;Մ�%���<�h ��ۦ ��vf��nc,�td�1HD�}B���Y9M�T{�Mب{n½/�^������|�;��L�Y4��zl�Y����K�w�	����VJ�qO8�I�[�&�w�-�S�C>/ߧX)?�k�:1����̫��&yT��1�F&R��\9�F��ȭ�;˜�Rأ���B��)��Y9#N��pg��;9���U�3¯v2f^�Ϫ'ΦU�e�0"���i �z�z�b)*���-�s7S��GF�d�E5�Q5.�ј۰���s���۹��if��	$��:�I�׻ً�;�6T��%SiY���}ۂ�9���&k���I$����$�	k�[#v/��m0���lP����*b�����~׿`�F�cV�c�G�l8��]���t��4�/}��� ��vS��=ȸ�T5�k=�l� PL�8��1�^�=h�M`9�&l�-<�[nc-��urv�$�=�Hߪ����LC�^�� /��x� D	��l=����P��6�.��9h {�nfǖ��ꉚ�%D�l�Yյh�@�>��F+�N�W��7�  z�)��	q'Wj��Lz}7��qܴ���&��"�6��3 "#kq�DqKG�O�)VGdnU���*���Nȩݕ9�/L8�}]�r	��U)���\�ɮC�)����׎ݑ~���;��ɴ=3&�=��?W| 	���X@�=]��%�w� �'�e5>�����ۉ�C|��[�� �=]�lû]b��	�#~]�?��t�I����J�S0Sh��{�k� ���WH��n�
?W�%}os0�#�r� @aݮ���߆�ߍ�X$�M�l4Ji�0q��J=&SM��a�7l�M�i\2�}����p�f*`������� ��ʶ��si�qc�k���1�;=�b��G��6X%��������i$ЇQop�`���V�|�We8��#�n��*����;L�ν��Hyh��l���3Q12����ݱ �cwm�` I�Tb�yq^~������>aݮ�w�AU3EE+�����PD{]��3\�m��D�)��Ʌ&ְ}����ӹG4����^~��=\�&���pp�I�������峷�w��cþ��v4�����ݕ�} l5)(~$�^�2��t ����3��o� W{����OGdW='Xw�� i���������+5lK���Jp��d�CA���y��%E����ʹ!�&ՃcT��8����o�������SS(���Y�+qGv۰A%=�ل�n�\<A��]VM�Ey-=����&&�*`��Og�3 ���.�g^�1;ޫA$���ܒM�����	)��-w5#����k'�Ϫ����LC����Ȁ+��x� ��U���]�s;.��� M�t��"�}�0山3�ST����P�y]��Z�����n(I^	��*ŀ+{��F �նwl�k�Q��������UUUL�RcF�?f` 6��o#���7�T�� Z<�M� ��vb���}M2:=��T�?H�월~�צz%���#��[��-^��f:}��Rv�2�m�#=�.��nك��heͩ�����X�M��g������ca��  Y��|ں�����oVا��}�O��x��9cs�u77�����'�ܦ͟dѸ(��ȸ:�R&ӽ��qT�y;��=��8�m�$�ްO�X���:�\����[8��j�#�!�nn�1d��ďVtiS�nH�ќV�]�&�8N��:.��������c�z�v@�� �{'D6�Q�}��;njՒ��.��:5��=��i��[�[vT�lm�����ywVг?7�ρ�g���Tz��������`|����Aڝ����m)�~�ܺ��{��~��	40�ᄏ>鰓�������s��� W���� S�l��v��vz��s[R�+@�W[D̩���%h��ng� m>v�>�QXr�\@S��nԾ��'����ݒNx=O����Dg�E@WԦ!��{����1D��p����� z��aO���ѽ�Gfb�.���GGav4�)�
a"]�6@��{f���F�/;��|�2# A��O�@��''�֗�X�C��F�E���ɇ���{jعw(���p�v����h�M����|pU�MULRӑ�o٘ mf�` }���`t󢰎~ų���{����W�8~�"T��ET�h���Vl�"a1!f�!>R��d`�G&������{��N�f�D��{�ܶ��������fb�w���\SW�#]�� l�t� dom�A���'��w��e)��M�zg���sJ��Ddom�T���G���}{���:k�-&A�ok��WK�T("&�P�
緱�ST�W�$�#ޛ`����Dy���y�
	�(u�Ĝ:��S�N2|���/�!�\osv ����,��]o�S�����M��t�k���sŇ���\=H~D�3 `�ac`4�W0�k�9�f��a{;oj2��CV�:y�fV������������b/�3�_�� ��� D}��ėEf�mq��]�X�+:����Â�$33E��U�gR���ѪWLn�}n��l�h����)7�f�|?~�����Bx�\�$��U.��6��	F>�<��A�ʵH����,L�s�Ӯ����S�3��bh�/%ȥ;�ڍV.�B�ʉ�Z�n�=숭K�"a
��b���s�br�b&\� �ݝ�-@�>�e��y�CXXh|K����������ת�"���@�@/=��b ��t���EEz��i��tr�_��4�������>1�zܤ�I�}�SǴ{�[Es�=��r� ��n8	?|y>��>�?п�%���2����T�f���W�2�le�t8Ɠ���0۷i�0�MQ��;颢J���{�ӹ�"=ߥ�I O�(�;�H��뫼�	 [ט1 �3�!Ɉ�L��e�TρtT�?#���]�״���1 ��� ]e�//xچ_f�9ˆ�R�33E&�]�Y��+6m��1�V�fmX�u�� E����DA�=5�-����%M}AUN��6�v[��r�[�cŀ�f�������sS-O��b�r�N�����^w��Lu���,㧁�:����y	�K�{q��A��Ъ���{-�22v�tp�v=d�T�<��s��|�����ȸ@�W^�	'�f��1}�4���_^[�i�n��� �Kd�vܰ�Gw�;��1+��뜆�:�ۡ����˳�N�*�	0�RQ3����aML�@��gnf)��� l��`�~�U����|��oԃ�I<���+<�'("�b	�򦻮���ѹga�'�^vM�v� @%�[�� 7��DE�Em]ߗ^󷸒�Ř��%L�*	��V����A&u��a"fԝ��gk(Vp��y�H �ܛ�h��� �������i�����u�����g~��Vxz� ��:q�a��Q"����11���7uxI)k��H1�tJ(����3N���۰�����u��������ٶ� �΢�"����6���ϱ�*�4!�o��G���1�j�;=��צ�1��{+{�����Ã&4|�~Ѵ�`��;��x$%]H��>� �(`8��4
 Ol���v=.�(`��}�@�[b�nzݻb�N�J�s���F��k�nw7W�R[��,�[YN��n��v��\M���|gZ�e:�<���ݺ��O��8[`������m��of��9z�v�v}��9���1F�k���@�ݸX���\�v�m�rtW�o��6�7c��ga�3�76ܷ�^C���ã�Z�qSnv��2'ۉ�n�T��z�n�w9M8�0�F6���i�5?�����X�cy+H��ʘ dw�݀}�sq*�/��9�l�l�� t{�t��Wk(��L!@J�Gf�f"fJ����O���@�	q��L"_{ݘ��9Ƭ��ێr�(��N1$"TS�M�<��X �_���`|A�)��7���̝ ��t������V����L�������&�lcp>�ȽSז��(�;�WI$���^a9�	��F�>�I�؊@Y��0�9j��L�T��+#k�� 8�ƕ7<�}��z!���̈́��AWn�Y$�	��E�Ӝ�w����{?��q��kur�!�壗Hp;n�#�H�v��˵n!�Q]��������C<ނ��2]�Dp_{����]��;���$�빰�&��^Q<qz&JD��)�ir�ۛ$v�����\;�9�Fb�j�FF���i�13@�R��S���c������c���=�[��ns�ݴ�;<<����%�&�6F��u'�A*׮�H�=�b�IN��������<�x!T2�"��R�����f,�+��q ]׼��;W��WTF�^o�1a�vK`e�� S1
}"I�S}s$p]M���-(�n�` 5�-�@�7��殱{��E|���a]O��*�PTE�fssd��{��Zq�q��v'�����{��yOd]�J;�K��{[��p?����ɏ���h6^Z��+d��Ӝ����w�d&c�´�������ٵ�ڤ���wz���> 8�Ʃ� #7��	Ƴ.��c|��;;3 �MnK�������?�-���Y&��������@���<XDDl�䶀@Fok� Y�8q�Pu�;ُؗ����(% �Si�ҳ��q ,��l @�OU��D�uß��1G����Oׇn/� ���9�Vn�1}���۸:��֎�d�^�cp2�%�~z�a��n"�Ԛ'o�|O��쨾C*Ѭ�n=�3�˯�� ����T�D�]ό��2�;��;s���z�2���9+�o��f�.�Dg�x .i�rޒIpѡ^C��	1S�U��=���j�>U?Skm^Ҡ��o5��:m�SoM=��l�=T�w5_�UV�vw��<z���d��|ԕw�g������qZ�q3�V���.Sw޾�~��3������7{�l��~�G�~Z��R�d����n:Q�N��V�o����Z�Z:w5���U�6�/Kl�UR�;ʵ�QQ�oۛ|`V;N�uL����wwrnoF6X���)�iؚp+w�g#h��\7�x���������69�"~N�e�Ww̮�F�_�1��6A#3��_��[?�w��_��\����~�@�NH�>p�פrXx�~�x�B���ň���5N���+gp�Ψ}t���{lȸ�ON3Z��YFZ�ն�*��d��=K��ݘ_o�l����	#=&{��ڱxoF4.���Ӕ{'|��ߟ�\��f���6Li��v���<!pyP���P��ԟ��;�b��"�X�0z�Mj���n=��٫����g�r�zk��ڦ�vA�Jf�+*��S�T�Df�ɉaV�k�x������8���g��:���e�T��k������Tn���H=گrr�πHU��/h>���p5��%�UQF+Z5*"[E*[V��6���\kUTh��[*mj�uLTĶ�h�h�U+m�E-���s�:nfW+PUs.5*"(��X)PKU���cQLj+��mX���a1Uq�Q���J�G��1q(�)hօ�ŭB�h�iQUDX�mE��ŭƬF�$���ETb������QDm�*���eAX��YiZ�Q�%���-Z��m��m(�1�cQs3 ��ۍs,�EUm�Z�ҋmA�,cl�aUG-]R��B���(֣Dr��kUX�DKj�eAP`�(��2���fZ*��XX���QjS��6*�KkEZʂ�E�`�+F�h���3Y��cZV���,Z����Kd� �Z"B��+KJ�*"�ҍ
֌��X���khQ�T���j��U-��Ƃ��R��-m��QF5-Z�T+4�+ְ�i[
�T�ik������K@�[�q��+��d���(�P['�ݖ^��9�� e>*q�I���7�U۽���dXզ4W��Y�D
b�d��TCb��m0@ �w��O(��D;+=6� �{{]�> ���3
˹�MןR�ʮy������^=���
�'a�/�]�Tm�s��O9�N���e�j:��|������ٵ����=�m��-��� ��٘;����N�4R�ȱh��<��XIwGLI�a���g���u�H��\a�	�k~T�o�n�� _{ݘ��9����w�O۷���]�,X�̖�sv6�A}�sŀ n�T����bo3g0Ѿ�v� H���g�K�>[��S�1�|]�?Ws�NO�O���m�� /����>�]��(�b̼���В�'S��tiĹ�j�ӽ�:H��v��u�Ww�fDМ��]]G;m��Ξ������g�@�۫�K�T��1 ��YN�ݖ�-Oe�ϗ]"����������H���  2���mE�S�[8܇��#�y6��ڷn.�#���:9ŧ�]1�����W'i����L�L*U�
���` _�z��H$��d݄�k��z#���뺴�J���{he�Q��1&e)%���ڶ ���1�=S��U�w� %[��	ė���EKdn�r�V���`-��QQ5EPS��ً  ҷT�Aw��[2���n��;������_a �얘OuI>DJ%W�R��m��j��Lc�� f�9��@�7��v�ټ��ǅn�u��H�o�.RS�p�n2IO�\ x��� -�m���k�k�g��πW�ۘI'�u��	 �;�	:[�m:�ʌ-U�'�U�^FZ�4S�Y��T׹Jx39�B��%1�[���O�^�C{�f��w�z�Ol�G�b��8R�4��K[��<�.�ʆ(|��C�K
g�sTgu�m�O%���g�r;�1��&u�f�^�[	Ӟ�n�/=�l��h���GT^�*���\i�ǔ�oN�kr�ɱ�����۞�*���<�8簪�[��OFF�n����l�������<Xڗ��M�=�J�۵�n5��ɱ�tv7m��������.9י@�9��::ի#���"v*�{p���%�6$
��>�n�=f�������+�߿���� f
�`���٘�H����&� }�k��y��e�����ϰ��MnKL�nQ�*j�T�!�k�wh���';n#��W�vI䚞Ȣo��uVK���>k/n�k�Hyw�Q��P1&a)&�5�ZZI$1�V�Da>qѻ�q5��� AչM2 {ݮ��yz"j�5EPRcH��좦o)�T1�F�|Ҷ|��k�H�f�d��z)�%��M�^�x��R%W�R�5�w�*~�<X�j�e{��Y~��O�� ����`|������R��1E4�:����������`v�&��%mWMPc�39g�������SK�98�$N5ήQ)$^�fbQ�����8��tk��>��?���7nZ�+��be(��$@*�.���ļ�݀�f����F�`pdX�U�G�1HgF\�b\K�Yw����}Ｄ��e��j]=�{���8�v'T[@�0��^�4^bjwm�����ޫ$����$�Au��Y8��ttD����FxyU�(��R���|w7@��<�����ڊ9���͜%�-��A6�����w���P0&b�L$o:��]P�2	��kv�	 �=�f` z�*��7Ei�����P�Ky�d��b�jӬ�$�#���;&ܧ�|I\�tS�����|��l��^Mk���^pN�N�P�AFB���L	�H�����{;��Qq�=���	Z�h8��E������p��*����s�g=� �We[���辱�_K�, �=��K
U��L2IO�zfa#����ZjC�v��y�A�}���We\CA�/u1��o�w�s^t@��4x�:_����]��A�U^�ԯ,q�]Q�)��VP<gf7z�u9ޫu�&�jo-K8��X��*D�S�uǜL��qqY�s	u�ש�z�S�+��f��"#�^, H �vU�F�yT�2�LJ$����u�D�w&sF��2�9�� �V�[�";u���Ӯ��b��?{m��}�������5�C�m[ �ݷ����4�V��s��m�3�	��6@�÷]4�Ɯc/��Ǉf��O
 ���m�vV�m��i��;n٭�<��n�M��⢸57�ߟ7�j��URJӾ=z�����j��t����f�*�sDF���̕��=�<+�k\��m�i?���^s;�tߵ��_���N!�û\ߒ'����2���p��vYbD���IL�&Tڰ��͚$�=�LRA"y���w�5.��[�  z�*�	a��I�&Ed�0`ȀU�]9���,������)��� >�ݺa~�d��͸B���M�Oq�U�n�ƂS��v ���j٨�h�<k4���mw�j�{ߨ�=�Τ�uxն�ژ���oe=��,��\�"37]�8��I*��8E�q�̞�$���ｋ5��xGj���Sk� �w]0_�ٟa7X��@��u��8k-V cd�q�����F�''m۞��wI:�Of�+~���៖�&��*"� ���� :7v�"����A�������ù��̃��t�	��3�	���[h��.�d�I>��v���~Ƚ���t�u���%L/�ۉ˝��+D
�$�K��w� ��ݯ0 A���^�D\uQ�~��;������Ł*�����*�TQLaY�'�lSmƢ��"~�f[��[}��� ��1R��bg�;��A�U**d��J���� _c����(�-W<�w� ���L >6��1," =7�-�Os�y�3�������ڦ��}�(�{f;��RD���37�m��zC�۽�;G��Vw��ղ�a�EKR�MT"���{��������������$u���l螕�gk�{<j���lܶǎ�ҹ{v�^5N]�Ӻ:�[[��`�d�q�n{�ts��A"�ۏ��[���7n9K�:����{c�b���sV�pn)˅=����.soj-s�vպ�r�X�]��b/=�z7M�G��ӥ�e���{O�v�ng����qMƌq��a {<�of�D�̠k%���kV��slb��kKE\7m��g��w\f����i�6۲�S12�߹}�I@���(H�w�T{�݂ =}�� ���d����]��8y�N��I.��3|��!f ������=�����}\},����X|�.����@�얙 +�i�P����o�W�?^�>��
E���D���`|���:g� ���mgލ�y�,�ݸ�"#�s�a+�yd,hc�Ǚ��Y����{b$��x�,  ^�ܖ����u��^�^��ʞ��	�����J�p��*�TQL�j�����⩻�~��f ��M�4�8ݹ�k��tTFB�� ��P"f`)���.�v��@^.���=rvz1i�,�q������?�&b
�[9�,��&��(�	!��E8��]����b$��Wd_�|�T"jh*U*��_�����,�q�8H��S����ǣb�f���m�D{5ҳ"��6j����b��f��ND��B�)b�/\V��;=�`���NZx��R[�f�*�{�x�̼�ļ��_d�@$~��1�����7�3p��Wg7�K˃:Lh���3��&�u��b�mP �T��ˣԽ�|�8 �{��"#8ݹa��Q5CH��Y���m*�Nݸ��$�0��Q6|��i%�|���[�����7�-���>�R�W�StγQ �>׉`���{�}�dr':��$K��E�"Om���&�s�����~|�{��䱧۷]�u�M���9g�WH뵥^�Oa���>7[�-;�ҳZ�| {N�j��]�ۙ�Ø���N/����d�vܴ*��TS$�*P7��}��>���ۻ�{�8� �Ӻ�@|w�n8�A
+^�Z̻�Z"s�q�;G�P(��*eR�����m* >s�n3�N�|�O׆<�~��Gz��I�ˉ3�k��ӏ+3�u���ݑ����VB4��+�����\غ�ӭ��I%���~@o��r�@��s0텑�HQ*�d���{��2Ύ!��]��Ҡ��=��@y%�]���p���-�N�yqh>�ڝ�����*�ILi���X ����x��<P<:o�4�;ϵ���w�)�'/29��oA�r$���c�͕��p�hӸ�s����n�sȑ�uEp8�s/����ax�6��=�Ȅ��Wm�vq"W��v��J���֩���t��ē���m+?t,Z �0�^�<U��%p��r�����	/��I�[��I�b�����gsy<�
+�A12LR���}�� N���Z	�=�&z�Q��ա"W�o�1a=u�\4o���D��S*�D7������7�wL�ٓ~��ۺA:�^` n�F�D��qK��M�gr�Z������)W$��������t�"���н��&�@�Mê��i��ғ|��w�3�C�5�yK����$#���߾���/ާW<
���� �_�w�8O�������I�� X�{3 F�n��|��k~*���v_�\�=���&0c(�vܲ5���v�Nv8��we=�Bf^l�WW������o��*�IV~���1`|��.!��ud��l,�5��u�e��$v��l�tW��*iT*�t�6�)�O��r������ 6�|[�,�m�h ym�|z�VO�Ｐ%g8�E)ET"�têsK�a��h ;q�+jKso^|�u�̈��m\?�W*�⠘��&)R��:�{>�C�}뜮�wj4 �/�K .�m�i�{;r$�m⌹{Ѡ$W��6	=W�%� H�l�}4�D���o0����bˍ�h�՚6����d�H��;�^Ջ�K���hm�sJM�aϤ��?a7��@�����T��:)�:��[}�����"�Ve���sH@��2ӥ����$��35z]8T��wIeUF�g)4\�Wg+,��� ^��م%{�lY���
��AQ�Ӄ��`]3��9Ŷ ��{n�N/���]�Ҕ����Bӟ����=3���s���[��L/Og�q�����8{�N���n�_+tl��������&����R�}��M37�rFƺ{u���ȧ+��`�(����g/a�W˶�'{5B��po"dQF˷���f�^��P�P���n��՝�.v�C8�2��k�Z�듙�X�rXn��B��v{�:��xY�QSdV��Z��%�N�A,H��uu�n\6��©�r�^� 7����r,��=�� �wt�L1w��r�綩�ݺ���>����y����gV�ν��<}�\jN�6�����O|%�]޻�Y�jkY�m�n�Z.)x��[b'�ux�N�p�bV^E�c��6��M����^�ǽ8��k�Z�:�z�W��٠q���Ͻ5��ll彧��"���v�Dd<�+ReN�0��c/}I�ډ6��� g��p���6
��l���9����H_v>9>��������u��+<����w�{J:t����>���Z}�1cN��5u�0J*yL�K�����Æ.�iy�����y̱U
V�-Ff��*�70C{i�eץ�F%@׆]�oC��ynsv�B�MZ�����T�Me���^�SK��[�~�6~���0�')R�5�TB�V�[T�Q-
e�ŶUX(�����PL��X�TD�V�����Z��S2�
̪h�օ-E�%�ڬMR�[�"�IQڣ4J�m���`���U5h��"�Ԩ,*�&� �U��Uj���F"1m!]%Db�-EXVTQ�H�b�m��+ұGT+����2�Qb�e�Zň�0�E+�miX�b�j�-j"�,)�F ����-�AM0��VԴ��E��eu�)A�Y�S,���T-�A����UQ�Dc�WL
�T���*�j�-�DF"�ѭYm��V2[+*����(�Qk%Q����ȰRV�ѕB��,-���b�[TAF�
�Z����Z���+QTQU�*��dR]Rb(cU���-��mb�21�3-G����J��Ձ��j,T�TR1�3,2ũ�e,�Ţ�jc�6��O�'��N�l��zm��h�'ٹ�u�n;6�t;�:�.d�7]���L�W�xŌ{FӔ�[`�NÚ�޷%�q��`�9M��r��F9�ԯe����㮟nn99t�K�۰�v�d9�76hpr�
*�̝���M���۝������vqֽ��x�j��m�ݷ;P ���Z�e{m��p�@��=U@�[;��eP6z䭈��ۆ��v��7cX=vy<hp츢�T%�(��Z�.u��aǍ��Vn7U�y��u�;D]�nR��v؍��G= ��{sõ�t3��!'�#�|㰔Lsι!��ݵ���5�!�3�v�'[�r�[kr�n;���ݱ�]�
�0s+�+�@��qĜg<i�m��x��ԋ��m���tٮ�A��0��v܏��g�ک����X��OB=fA��N�����$�읙�^*Ŷ�뭃��t����D�^ۋU���u���c���d��\�=�];�r��[\�g�:�[��F�7iȉ��n�t3�`ݞ��&:1j��V����[��c1�Nݺ�V-v7µ/nӞ-u�ڳ�n�u����3��껗�s׈��NO'�+��l\8�t/`�Yi�G^�n+^8��㊎7:�'�>��Xv�τ�v{l�b�9c=۷6�pkaU��燞��nq�y�}=�w=p�۷G7/m����THZ/	y��Z�1��;F[����WnݻI96vՍ��Cܓ>���v�%�2u�[th��a��㱏\ݥ�s�����]�h��y�ۮu����s6x�Ei'=�e}Om�eW�(�Vݸ-�����ѻ�u��<gz�AW"F�!D<��dRT����6��z�dӓvuۆ�\>:�}��밍����oXNsٳI���d�蹎�G�tp�ַh$�D�9;��N���v���K�u��@=sT�`.s�^�Bp���v�)�ѧ�� �l>u�˺4Σ���ܧJ^�utN��6Z�J�k�
���M9��@ fl�e�pK�n`�!���A7�;�4�ôxy�G]�g��;�	�8 ��֗��\=V�l>��~�뺱�-����gur=tش�a�=�����l�:P��7�ks��v{O�gI�۴O	[� ����,	��:�ڶgxg�������h� D�%2s�l�̚ӭ�X����k�[GW��pbݪ��'��:�.%30q�ZթF����{	��r;��AWnp�]sŔ�'C��>$�u������|L�`L�L��W��b,�Ou�i ���y���3",e���6!9��Q��[��ޭ�5�%UI)�ݹ�s�&��l�k���K���ȴH$޹�~H��s�f"N0���	՝�*����7�e�ˊ 4x�6����M�@���[��" [�Ş�y�� ���i�Gy��XJ�q`�R�hE�T�ד��`����S����`g>���u�pJ����4��H����|Ik7G���i<�[�V 6紶���HU�n��׺�F|�}�هJ��=9������i���x�x���cl������l����OK���[Omj���%������pά�!�{i�;_kİ 4�ٶ���gFNR�ڜn�4�|�s0����U3R������;֋��&������=�M�7yL��x���5�޺���Oɾ����ӹF��2<C���on�}}�f�J���{�dd�'��(>�y��$�W�(��WX�d��*�s��/g9rM}IURJc:�ٙ��A��������J�3��Y7��gf�b�=7�-�����P�TM*�5.�F�Kn�7��zw���<X  �o�\C@}���ff*Q��N�
,gofg����"���E:������[˝A��5�2�g�-�ƒ��y�� �ײ�Ν�/�,Mt��[j�ɳ��W5�.3h�+����`�8ݸ��].��l�WDȘPLDV�����f!A� ��}]٘ ���> >Ν�1��#��6w���y� y�4�#|fJ��fLMߕ�M79uΛ�ѕYݚ�, �{M� YӺ�!����O9�$:9`"2�30�H�;���:�ubRH����A��./O_���o!�}���t���w_W�2��w�yCf�Y�xL���$5��v��w�{t��Ɣ^�ߘGǟ��>�xo?$��$�%�{��o=����u�ouz�T��T�U$�GV�~b!��a:� �Eֶ��|Ӷ��I%�or��'s�`8�:PIx�dP����P�J�R\��p�t~�~�&�k�bƳ�$�M�	�7Q~Iy$u�����-�<�p���
l�%E�y�]�&�u��s�rn�7k���f����/g�!��Ԣ������l����@��}���s��@�g�6@�4ݹaEC�52���"�(-����`ݨ���':ǣ.��[ H;Nۖ�#9���{Ls���U�n5�d��"�Ҩ��ù�0���/�� ^٣kgٻqYs�=<�� >Ξ�, ��s0=:b���DR���P����7�e�=;�}�� fm� ����3zy���[�6��-oR�<��17�ګ'�l�Ў�YH�oU�m�>n>�y�\�(�}ڲB�/w5K��{тz$"��i�.I� ��2Of\�V��\�Q>�13	d0�o��H�OLr���m�'�u��D�I,�o,�N���j&� U+������gY,�Q���A���ўݦ�� n}���QW����ղ,�����������j=C��� A�}��|��e�
�rs+/�^�`|�{����P"�R��QW^A�^�L@���"|c�y@ {�u� �O=�� o�U9�V�z� ���SS*jI�)R�����`ļ�-u��m-�I�\�:2㻞 >3��g�D@�O=����PDD�"LH�h�.ꣷ�p�L�{�	jH�7���`|�#�{6�q�sK����9�'�,$��7�,��X�T�$L�Ԩo��mS>��7m�G�lr�Ɍ�S���  GN�����7�:����λ��
)B	�jK�-F�vK���/5�ۙwY6�afuM�U��)���P���˶
_7t��ƥ�\ّm	�kY�2�#� ��ZL�˸������=���烶���c۶�����E�u�<n�Y6��-�u�YvГ�l{%�W� ��=Cd�ڇ�}\�g[�E}�UpiLu�L[��i4U��T�pM�]ǝ�;��p��b��nN�����*�Չ�q�[ �`��[�ۋ��[]����y��[�s��*�g]l�q9�m5�m��sv�G��n�GV�8�����k7��N��ݓ]m��v݂����l(q�^*UMo����������V����f}��I�n��^I��Z]��[��G1��Ow�3I$�ۊ6 h��$�D�"&.K3uRI���w��v]�䗒���h"�n��~�K#��ڻQ��or��S�Qb�UJjQE:a�^ʹ�#�ݶҰ@ʲ{Hά�u��� =:�n!��n� ME⪘
aD#"AW~W��)]ov���h�O'ݳd������Ig[y�w��w�;�<;	?��HI�쵦�,�'�	0����`���`���T��S�^������4��Q �给�{�v`�7��'N�CD -�X���C�k��6c��ŧrv옷c;�[74���ڄ����[Z*�jT_=ͪb���ۨa,给�;�r�gR�$�2svZd /�u�Di��S30�Rau=��bI:Ƕ\�U����3N����I1���Y���3@��=	�y�a>O=�x7�m�GVe��U�3vmN�������N�~Tπx���3���������WY�)�U5E�Ꭱ%H2 ��t΋�ڰ������u}�eս=������Ib�w$�av�yg�N���\s0�U�����9�d��
�ݺ��s��������;��b/|DDR��ΘP����$�)R���[�V���Ա���as�2O��/Θ���F {��l����~�4�CV��+6[۩�� ������ؓ���6�Jh)�����Mչ����㻝C@ �}�>� ����6Վ42�.��S{s~I�]��`Ć��Y��M&�I����(~&%="rFeE�^��n���I$;���I;�X��W�]���ݼ�zc��ߒY�0�)���Ed3��m��I'�S��1(/���l�^�s�T-g\�eDG�ts�a��Ot�*��,�O<�q��3��C���=�{ۓF�:�>�s�y{n�r�m9?x  ����O�I$��}��1 ����4�)^Y�"���R�SR�x��d����Ƨ ���b �i�q�n�W�S��ʿzPG>{x1!+�ɑ ʛ�z�^���	i�ub�_t��\��[U�0�p���÷]?��+�o�ާ����\������]�b�$�&�m2]�v9�q���囎:]w����E����>���>@|�z_���dv���/���;�n����'H.sz���OA7� ���!���шH�s��EV�#Y�r��� οK �t�"/p�2M�P����{���SLLD�6���m�����vj���V)��]�{0��?K��Gn�0�Ꝋ&�D�T���+�ٛ���b�(=�� 0�����rc��/���_7��4�}<�?{���P�[ڥO��0�'Ԗ<�ꀍ펍��]�R.iT��;o��s`�d�� �u����y����L=;���4a�MG~�$� ?�{��O��Co��˸�0�� .�۶�#��szcw�<������mb	��D3�H��\�륶���`�d�jۊ�9���M������ߎL��T���`w���VA'ݴ�·����^�{�D�E�s�&��
S
 )Q뗵d�;�bc)]�}�3^t����:	��~��7^-N�J�7"��H���0L�"M���~ �_Wm�� �Ύ���{��$���v	$�{~��V`SLLD�4Ev��©��q�ʩ�#/�hX 㧷`�Aά���#�(�Ov�ݒ9��D�*&d��V���u�_��W�ǵ0J��b� ��m$�ɢ�吅V

�:����h������R��Y�W�RK4O����Y����ocy`�ӹ�K�m�E9�o+�^\+*(�����7;��]��\̷*��5�"���]v3���۵On�-����jSmհ�wx&�z��u�g vc�;oF�yX�ۘ��֪ݹv'�:���U��n7nf�.W'c��yy�ll�
��4ܼ��º|�}G����C��X����ܓv��ݫ7�I��Ū��ݜ�����;&�8�/5���n�����뵭��o1������D���H+Q��'�N�Ig/=��j�û�]'OM�vS�e��GLWc���m�|�z�D�Te��H=��Œ9ՓF���j�l(��n�W:	�<�Z�\ �1&`̃**�y.h\"�!Guu�۴���:�h���f��j��O 0E)`�
aD"A������YB�"�hw����;�^q�{v��ά��zJ�A ���b��~�j*޺V~�ۀ�������d�$󛷛j�2�]vb�v~�����iI�=�I�n�ŵdN7n�y��{vH��ɠO�9���v��5�d��o������o͞�S���wf�p���'c�n#�w
{9V	b^m��������N�����:��X$s��Q$��6��V�FA�}��<�&��ht�@�"D�n�8?����_�v�NT��7m�| v�1=��'ת){V>�_V�њb�'�����.��� K(l������k�%��z�X��j�����*��Y$��ɠAg�ݓ�������*��Q| �f�2��9.����ud�@*��t���ɬ��ǉ�dQ>'���$BVQ0����(�1@���;h��{�Y����A>�����۾�T 0� q���0�x���?��7~���/���8�ŕv�g��;č[�	�9���'ă�Mس�x�N`?���<,��$�5��lKk��<u�������rm�'C��9yٶB�_>~�:r��&"`4{j(|u��X��M՛�w�5���k��5"�O�[w`�>퀼�C)��0/��2D�]�Y���
$��y���>$�nłe`{y�b��eOx����>�"D�"&"��.�m7~��|x�֯IWΏJ�V�U,�fk<��X�������)>^N�n0�;��$���t(�����O�Qn{��]�i�\���n�==����zc	�u�O)�q�7cB����G	���ҍ����DjNt]�Ӑګg�O�t�o�9{;�q�,y�ڴ�*2��G��z��Υ5�O�xL�ܕt�ש�=���~����F;t`�ӷ.n�;Zêr'���Ptjp�XE�d�e Q��2'�1I�le�}{�y��6�Ks�We��n�N������	�^��1�:⾶�s�*9���c�i�sbp��o��'r�/p��&�9� �,p����^.��=*��q<��w*���yz�VqX﯐�o�K[�ۚ{%]�����%y{��t�B�x�Dw�>���
�a�ĻtzM�γ���N��>&�۝rl(y{u_w�K�>�o#�޲�B��J�9S��M�f�݆Q����{�ވ�^ūQ��;^d8;����qL�y��Iu�>_<��O>�ڻ4UV7㡜s�U�M�?ݳM~O<' d�C���We쮧}v�����N� ?���#�us��jO��7��Ҡ4���yߨ\��b�UP�Լ��u_.�^�Rk����{��棯;�<��6� pe�]���[��k4�)�-���A��c��a�����~`�;���ݺJ�x���x��h���7����w"��1������ؖ�m^�Dl]1�K��<��Ml�U�� �	�E?\���e��f�c3W2�U���jW-�XT�YG��ʩ�X�[R����e�i�S����nek�*�X�*�L�PU�F1EQ�أmQ���Um

��#�Q`�Z�X�E�ц
B֎S-Z(�*j�.Z,bE�ne�J�D\j��*�Ȫ,�f#iQk+�D�&2k(���"�%�DGIcR�6�MVVk

�Ƞ�%X�1V1b����*V*�����R6� �Y*4�Q�LZ�����X�QT�,P�2�
ȣr�QUb�CEDEE@X����-��D11�t�e��j%�X�mZ�b�EH��7W�T��ȢŕP�уl��QjQ�Yh�*Db�d��T5(-E��UV6��j�����b��lT�h�P�`�E�Yl���,D��5���U"�,QmFTi�cFɦ����C
(��eVڈ�(,)h�(�kXUB8���\e-E��PX��aDDDWL�*��R۔�UE1�¿ x'R>'����I>?m7b�Q}�fh�Q/�s����A�ڈ}mۅ	D/ms�X9Փ����ŻD�޻�Jb��f" J2P=r��i��Κ�B�t�K}�v	$�\��8z�(X#[��?�E{���x�.i��H��pt�eH{I����>�\u8�D�??v���g}���I�/�����]Y�Һ��m�����\���0a)�LJ��t=�BI��8®E�O>̶���8��(��� �vc ������fL@��{v�.���AP.D]�7��m�~�]Y	YiG�'<CKs�Y&�R�w���v�	$��ȢI���r ��w�f�@��� �/t�
���C{	Q�[��을��ޥVr��kD���X!J_Xs]���eU��߀��q&�;lY
/�(�B�1*B�g�K�'ă��u`�[�t����݂I��h�}����;��Ot�Ђ�B)/�	�a��Ć���=r�:7Oob�m���a����j��9������|q��\�b�'�k��_om?e\�3zV�o���|Iͬ�$<`ٌ�J!)���u�� ��GE�wѷϬ7k$P��y݂N�(�5Y���ݦض���$Ĩ���SD�����$��1t2���Y`�O�}Y4I=���s�;d��2b�ݔ�	)��� �Fu9�I�۱`��z���2�Ǵ�\�+m ��D� ����wv,�ۏlY+N�٧�[�3�f�&�yՓ�A�ǖ/zO
#�*z�_�#F�k��x��} �2��|�{��[ɷ�;w�K`�X���g��6B�q�]�ܡXFڇF����FlW� ww燐?69
��1Oc�v|���q��;>N0/1���v�N�ݲ��e�m..P漮ԙ/�]����xGzܕ.�9śc�m���NN� D�&��q��#�<��ug�2x6��l����p9su�.G[���q�4n)�$p�u<�q)�n�t�mD�+����@�^9��K���I��b8{r�:�F���;st4�ӰQ�V�qa���#M�;C۵�K�GnWu��;�rn�V�Z]\M�����u�$)Q_�̗B�'�_s�~ ��˰F�ԛ��N}^ǯn�4�,
�TDIJ��^زh�d'iyL
U8(�M�=�$�{q�:5�*��GH���,���g�.x����;.�>;��|��m�U{R�I:���H=����3af�ĩ�
�G^����ӓH�s����㽝�d���Y8ʈ�B�H��۰O>q ̑�dL@�1ݷvA�:ʬ[��O����'����;k&�R�Ճ�T�'�iB�)F�FfHcu��E���b��7>���D4���כ�H��?C��wH�"D�9�v,���,�I ��Mjm�NbJ�5}X	#;�/�@S��?���L�h�z�<_�����)=+>�����fN�4K� 7q(��'Qc��NcC*�)�Cw�v���✆��wO���ۿ�� #f�W��@<�2�Ēs�ɠD�(��w<�H2mhT�2�"JPPo�l&���\*�Ηn_wg���W�9.�o�Q�,�j!-�P3 �J�&F���yݕ��'��7JA>;Y}V	�'*�I$k�ۑ:Ȝ�12�7ջ~�=�,(�H&%L�T��4H9��Y��,���T��[t	���d�A��{�v9=C���|*-?�D3��<	_/Ξ����]�y{q�Z�Ǥ�Jn0�C`��_�>(pfH�Qf 0���Y���I�m����w9����w�:�h�*�rUQ�L)���zۄݹ����WN�y�g��|so&�/�w��/}6���C��Պ^�L3�L(�����|H=�νd,��/�,��P��ED#�����Վ����<�{��f�{d9W[[������-u��X��i%n�#;\� ���{�� DD�� ���@��?zL��:pcH�Ax��=�y��<ؽ�8}U�B��o;�	�����칽~�nԊނ�bI#D������,�_ve�| ^�z�	5Ss@�o�w~���ٔ�,��X���ǂ��U�e'�u��/�9=M��͋ɲpG����2�[N�BN�a@��A1*f�+�P�@9�άH'��.�F�vlIȫ�-Ӛ�c�H~���7�Ra��������&Mu!ݻ,���VH$יv9Z͝@�[=S�;R�H�
Sd�2 �����g�$י~�H*wT����)�NgI1�V	'ǵ�_��<0�&��R&]�K���7�ηv	#;�� ��}�@ �JۉC�ys�|�=�.yJ�[�E�f��~cV�zMlΫQ�������uf�O��z�vˊo����LLf)yY��wLFRڧ91��|O���`�{58�-�/߇��ސ` ���U=}�:���>'ٵ�b�%�̡`�s�&�S����k^F�ȩJR�S1j5F�7n[�2;\m��
rEv�I��TĤ��+�h�`H�b��� I%�f]��Nu�׏V<c�kj3k��'w��x�1 �O��e������w�n�8��rJz���)�I�o2����ɠIS:�Mϵ����~:��`1&J�&bY��v�H{yB�>=6�}U{�������H9ד@���0"D"S]6��P�����`���vI� ��M�v�vٓ*4��g���u)��&bT��dvK�$�w:�c/k(@�on�$�ɠI=ͻ���n`��6%ߗ�-��{n�Oz��3ϝ�]�[d����1,�akl�aϧ5��A��IK;���xs�ٺ�LX��~����s���*\]����{��~����o�p�<\#��ö��k3�{x����r�N�y�y۷r=����tQ�-=����p��Q��۝���(3��l�[q�<��U��k6�t�`���`�ݎ�vqr���zr��o���l���p�ۛ1XNBǀ1J�9T{4�os3p��p�ʋ�:���R��7cv���=����÷5��]��հQ�V�H�9�=��rݔ"���kuu$�{Vaݤ㍂�T+������|���JW�쫝�ωo^U	�m݃	��U�*��=O�`��y4	J��R0$I1
�z;���><*�,vNYk�K��;�d�@9��(��Y>6��.��S7;]�G8Yb �Q>10fR�)�PA �n��ќ֦:��(t�$�&� �m���>�Q���B��1��uJ/u��ѫ�����]P$�kw`Ok̙�E�V4X!�9l(ZH��A
b3f�زOḵj�ٍ�Џ�����/����יb�.[����T)��'g��/n롸�)#r8��u&�5N5��*�]0
�����LL32�L�~ۍ� �>�W�I=�2����/)U���v�
 ��۱`�%�D�&!L��@���M���,�6����s$�a�:5'4�~WeCF0r��i�iLI�l�\��^!�g�m5�@��/�Ց��Ʋ-�7wq������J\�՗�pP�� {�&�A$�����X�n��*М��-O�#k�%#L������'��ݙB��J>n�g�F��@�m݀A��y�,�6X�0�O�L��=�W,ͦ^��-�ڲA$��̿_�u�b�e�'z�A�}�`��сmSx�́~�� �0xt����(�S=~� ���,�}�v	>�בGf+��_�n����v�m����ٞθ��>���٤���%�SLWc��~|�����w�~\��� ���,Y���"���w{:A������޶de�~ƃ��eH9.�$�w��v���`�@�ٗ`��]y�cw������4��$�1
d% �;n�ŒN���$'��zv^Z�n����ɝs
�֒o6��f�uF�U�j�]�)V�=���Έ���VF�jI-C�;�VT� Y><Q{3�����w�c�H;�fX��"��F��&Q�Ub;��t��C�/�[A}[`Y�@�O W�#��cv�`���	;[W�X�`��3)W�u@I#�[�=v%�aEO�άw`�F*܊#��VycJ#~B0�'�W,uq]��N.�;r���õ�[��q���V	��M��������mSx������H ����I'ľmݑ��#R�7�E>�!�x�`��nEx�%���@����P�w`l��91�jnj�#vEI|ۻ�����3y���yw�Wg��v4M[.A�+�`e�����,��}�mlDۦ	�f�"�'�ͻ�O��V�d��m�-�~���%o!�J�6{2���svk��E�M T�i���(T�� S9��މ*�`Ў'Qm�U��J�&��q���RS.�2�ܩ�>S��q`^�+ݦ3?{�����{��p5�b�)J�e�[�﷮�I%�f]�d�SQK��P$v�;�O�=�2��)�
�1��&4���$^��@��%���A���"j1�ۂ��;�T����B0O�L��=� ���� k̡���P'�Y	\�W�"�b�i��aI��L�[�3\�p�������f:�I$��;�A�2��;6��1p�.����	@��b)ͻ�'ă��.�'��=�.�fƒH�mز|ḳ��LJ2�T�f�K6���]R��@19�d�	��.�H�]yoz-l�R�+���T�THH&�/������8~�_�g*�~��3.r�3^�#u�]�p��Q~��K���V6V�-�Ә�K�5o^�U"����,f���v	<ܞ'6����v�Z4os�+���Q��Y��A�2�"�Ԋ�kj^��FN��i�DaO=Y�ʃ�JVf�,r���u���mL�E<O^���K�;��,�ɺ��s;��*7f��������E�Ś,�1��2��7�Q�QB&�����<[��e�w|1��>�g�<�GB���NI�=;7bF�	�rGw�y�{Ϧ-��v�q랧�57�P�{�[ǌ(����{
��קOkD�x�=����������b�{�N�֞�(�Ĺ��=�F�����C#�R��y!��̑QP�A8��A{���um	�K�q����	ܵӓ_�]T�q���G��c�x�R���d�U�˗����C\7*�R{���)���.w�g]�wNX2�5�2�j��B��X%�'S�7b�$�SJ�E�kc�2��=Ч��|2;��r�Ə`��w��=�
�����-^��v� ��e��Z���ܫ��Z�-���=����A^<�L�wh����#9�9��zM9#!�Ŋ�	$"#���&`�X+���v�`�/y=�}��reM���{�#�T���3�%I٤c�.ɦ�j,���39�*�[�Nr�ԙf�r^�ǜ�Zb��i�y@t+r��SZ��Ȓmy{����f��n{ֶ/�I�6Ǘ�H��)�fX*^➽�"	�I�`��������W��Ȏo�R� /��_k�h�|��6An�o������o7g��"�	���X~M�Ⱥ���DAb2�AE�X�ұQ��E��Rah�(�UPƶ�`��(�
�Q��Z�"()mU�"#��U�Ŗ�V�X�1�D-�Ƣ�VJ"� ��V��Q
���QkGWI&5
�B�dY��jl� ��`�� ��I��b��T�����Y��"iK�F�UUEp�UX�F*��Pm�YR�̪�UUL�tª�-UQ�,TDj�TT�rŹTZʋmF,U�T�*�j�[��Fj�ePX����te�	#����c��V�Z$T`����Eb�T�naD��c���QQL���EIWWW"6��+�F�,-��j���r�J��5�1V���*���Q+E4�X�Z8�Jj�CN�
���1G(֕EV�`�����[eE���V(�-�ZJ:�a���&�&Z]R�5lDR�I,\��J��UA�UeB�1�+b�,U"�*�X"ƶ�������Z[bռ�k'�0�uڥ�v��v��m��og�v����.뾋����p���5ƺ� �v�tS��!U�j��,nn0K7%���r��Ӷ����ճ�u6s�5ܐ��d�9�خ{e�ns��L�o:�T�v��m��U��˞�k��[��W<e���ltts���Pۣ���T;z$v�f[���=\�l�aި;���9wFv������m9iح���=\�]�zne����+�)܃��S�j�w61=^�Kûlb�^���XIM&�]�<5����#˹��������W�m�v+��ώho=�r�ƪD��x��4�M����������xh�ͦ.6��5�6�N����<=�E:��uͳS�ڨ��c��sK��S�]#7,� (����.���jU��]�Z�t�� ��ً\�h��2OZ7n��:�0��w�1��������kl[��.�e��.��ص�7��Wg۱�ݗ�,�Ξ���M_W��\��m�oV�ivz�xM��7O[�|l=�g p�8��3Ǌ+q��vB��oeCDwbx�=�����=���$b�y��u�j�<�s��Y��Ԧ7F���n��%x�ƀ��s3\��;��kCk-�x5���`���Su�jc���9�q����Ϯ�]�緮���M��Wm�;���ѝ������lpv�䓝�xu�-A�i�-9��a�qu[j���=�n��V���M���c����;s���Nۮnչ��&�گ^�0��,������͹,jx��<u���oV�����{e.!,���k�x�i���+Ρ6�A��j���;��7\���6�;�Mo]vE�7r]��;lM�8�<7Q<V�?�8�>�O���.-dO^^�2��r��#;�Gg�6��j7�ݰ,.�U(�tp���g>�`ɻkj���bv�od��y��M;mp�y�	���V��v�}[K���6���V;g1�^���ݹL�3
6��-f*:�����-���w{��^���隣ß{����Y)pLt��ָώ�����j|;&�w[ƺ�hN�אvy���@���0�xu�l�E��q�l��܊����̱G��tێ�Uv�X�v��gcdڸA�9��V����؋�����Ƭu�Y�x��ƨ����l=�
��M��p��a��9x�ڮ�'�㮷Ov��2�<Ym\E�h�VnU{A�������\�\f�c���rA^��[J�J�g���~!%0dJ1
������K�̫�z�(�m��}��rFT�X�0^�l�^&�D,	��A�w0h�۬РI'v�ԷZO���U�H�בD���zGAP���$�=) ȉ���c�	go+�@$�wR󑋎� ���]�N.��E`��a@B&��W�mݢ��@ݾZ�xӺ��8��Q$�ͻh]�}U{�ě�N�`�	�DLJ&fblq�p4�w:�\j	}U7�Ċ���'��V�EH�sn�v/p������`÷5�z�S˛��燲��.�n��cT�o<Y�fܽ�_�����=xj������ݟt��I �����ܳ;���<{��}�LOJ�����
�	-%B�w��,�j���������%YY#��=r�Ng	��C';|Pא�Eɡa�T2�7b(;nb��*�NF�M�ùL�Ε,}��x�u�_����$>�[��$�Y�Z�t([z��%� (
'Ц�BK��O�[u~$�`N��j̕]{�CA#^E_kwd���tB���.���oMҙ�]$�|tͺ�Ay�ݐ@=�2r�I3�� �]��Z�P� )�讪��Gḵs���Mg]-�eE8�	�g7v	 ��yb�yۍ`J�@D�	�bk�5m{e��a���
u��ζ@��:�H�@�K�����!L�P�Q�$�s�:=����w^[�]�&�(�3���#*P�F��*���ز`��#��I �����Hv��	S�M��]=5]�e��0ELR�I��s���Gѽ�h���w=���������u�%��޹�&�R���o��=�h���sow f��α8����{��}��D� ]V��#j�(J�� .>w}�F��~���U�6X���%0f�h�ձ7���䇣����ʲ@ ��̻�'Č]yi� ��7��[�wd�����$0" ]��wV	�go(M��6�%פ����$���_�O�.���������$N��$��x��M��I�kѝ��� n}���Ea��x��ȤG���߿�0� )��9�wd�w{2�A�ב@�:�{�)��;G{y�Q��n�9Q�8�mI���ی����`��$	��.�H'^Ex�ͺ{��z�H3C*PRT10���w�H�בD��lv�gY}Q��A�on]��]yM�rJ0�B`ȕ
ۜ��>监�"6a��n!�>.��'؝�Q;y���]=�����s2&�f�)
����m�#����V���[j��Fb��,���\�s��rNه��I��{���}�A����V
��Sa*��T$6�d�\�{�B�α~'�S��� ��������/$����P�WŐH/��m7��n:�W��٫�;�u��wsڡ���ϛ�rI`�x�wW�|Y����A�gs� ��S:mC��;��,H��"� �����B�#0����� ��i���]��č]y���s�$�p�]}6�+ޯ�z�f�F4����I ��s���?r��N�q����@�}��ذnFQ���&baD�t��/��鞚�EP$���O� ����{]�][��N�0����e�$JB`ȕ
Xy]�,���o�މ`�Tl H��QD�����Xv�����������e�Ԃ5͵N����H폮���.xd/]�Ā����Ve�&!N>d���=��SX�s�.�Nm��Ȝ�v�n���=��zO�^�H�6�EF.�8T���zM���t6�ٺ�q�˻&��m�)f��z���s����R������[[YκJ��%�խ�m'&�{q�����-���K�6�.��q��z\�[wm�u��oV���<O�$�z�\f8۰��y��G�5Rc8�<����uZ�#�&جvȤ�uխN;�������˰h��:�գE�N�Nw�Z�xSa�Sj�[fӞ��v�W5msO%���%��(
�!)�0��h�	9�VH ��킪ܬ��W�ys�<�^'u��;�z���3D����6O7�9^�R�.'`�Ӓ	�n�v,x�޼�`�����%�p�>+��I�>Fa-��I=�yv|H/�=�=��uD8���p��K'�����2�m���+%-��A^�Ȑs&�Y��yvI8��)U�^�3�;2��H5#��RT�b"����'O^Tه�Qݛ��;q�v�n�'Ğ}yv��ב@�fC�w$ ��L�i2�@�d��}�3N��L�cG�"q�S��R	2��2Pzt�P���� ��yvA'^E�O�U5�Mc��nłNk��9�Y* �3$%0f�ڡ$��^��[�����֊rKS������1zo���{yC�n#�wOC��0���GT�ݼ�(̨�YY2�_����{_A_^X���Ȣ|g��'I�:*�����4DǊ�0@� �c�A%���'��h�v�p�Q{��H�ח~8��(�1$z"B"aW�^]�GV��dH;}�vI����$�kv�4��tP�I���FA�B32���7`�R�}��ՕU�W*ك �{wd��k Q���f�.�]��Ș������ k�}+����˵d�\;��x���沱.��;���R�T�D@1�nqг��(	 �{�����ٺ[�n��O�S�j�λ�#['�D�Pn����|ocaAζb���� �ru�@����;�73�]�T�?Y��b
&d����/j+�������bq]�*��eWL
f��lD@NnMlLD�n�2�CTǦ򃱺ӛk^�FD��U=�,�ivF����T涯�;���Z��%���W}�ط�W1�L,.yO�^ñ-�
=�BA'7w�|Gm<�TMD��NVaB�k�x
�ȜD�D�D®�˰;e۴�-DFC�i;��>��q@�m�w~'���O/�3S�,`�9�$�{0�us����+v�煬^{�	�u�l͝�U3&Q31�wGA��̨*f�Y�u�$�o�_�v�ʳW��O�54��(F�s�T��)JPJ�1P�l��9�fޡ��f���=n��On�Ϧ������ب��l��,��6��S$��.ω;R,�d�;[ѻ�4�su`�|{i���c��(�Fa*�m��� ���вI�d� ?��=���RR����t���A�ϲY<��ާ��K�p.����8�Bz>n-4t�$��s�e4�%Z��r��_�������������	y�vN���D�(�!D畢Ϗ��U!;0���]}v	�u�~�I9ՓD��5�2b��Ε2;8��M����]"�\�.��ϫ:�[Y9��g�BL���۲� x��4}Y ���O.�$�Y"�J�Um/+�n�Om<�=(t�ʂ�`ߜ��P�ܹӐ(P��|�2A8��Nud׉񭿿8��o��5����-#�n�{j�#z���|jR��]���I#��̘_�^�w�M4��2�I����<��n���<I�Ƿ�$���"�/��o��U���M[���R��$CD��T=�Gă�۫�w���± �����������u�y�%|�����ۮ�X�*p�UV�Fr��vV[�,R�!v�M��"w��[.��tt����T)	�Lh�	dK���̋�Y�/q�l}� <��'��I��	R�J��`5�7Feeۮfj��ۈ�2�o��Q��ɺ�n�6����V�������&m��#y��Y[Gm��]��=�bvp�YF�ŻC�xh�n.� r8�1��j/e��|���� �n��s��1�^8F���:�3��I�]a�N�<�}vY�1̑v�^М��m<����"}��ځ��0�c�գ}C���Ӟ$ڕ�C\];9ownX��׭�tay��l+�mT�ߟ��|��J���
 W�c^��� ����A!��vș��Yz$f�L����X ���h�ys�=(�aWK˻������=zşG^��'ǻ[�$��hg�&�_A�B12`��5��tQ� �>ud�3{�sj�N����A{S@�ݭ݂|jC�D�PLJ��Q�kw]�[�H"�.���s�wd���V��w7OU��p�A��$y���^��)DA����~$}W���5CA�@4�&�$v�v,{������s�j��7��s�:ב�^'������գ���v�gnzP�*�=��������4v��!��(�^����Gu[�$ǉZ�B����og��>��w`��)���0fB�`�:�K���E>8�TE�{n�5W��7+v�[�Nj5$TؠT5�t��	'����b���49�9紡ߪ#��a3��K������� ýϨ�I߻�b�G�W�`���x�:�J���`�e���D�D­��w�@$�����'ǯwgcҎ8Qn���H��wd���W�g���!�0��7�����k�1|�Vfu}�n�Ēr�e�P�fg��jp�A&P��B
(��u�'�s�E �ƈ�ݰd]�6	���|IΫ��.y��x?D�=��'
),A��! AG�힭k�3�`t;\��؂��Ѯ֍�.���>1�R�D�#sz����}VA�Ⱦ����g��/wO�߶zAyL�3��HR��T��� ��ɓ75��*���k��[�w`��r/��O�q�Y����=�#wJcD�)L���1ζ�8ܡ@����z���Ϻ"N�5z%l*�yE�L��>q��x��P\F�dQ^����\�><W��\�������f�!���G��������z�:s���;�G����؞�5�M����:a')��>�n/y�8����:%Cag��|Fo=�Nni��ow=���xW?o�2Ư��&0������Mol���.�<�2���T��<�-��W��X��μ/���/��עu��ވ75o&�s�No�}u��m��s�uɓٺ���p򡵣;j���v�{7�0�������~H��B;;�D��քY�$�����	�������qj���O��5�&�GTQYX��K+���l^>CЮ��?[2���m�t�k�=�����f����X�M��~����5� �N���}s��e�Ow�}�S/'w+�����8�)E��n^�|#ez�μѯS���l	�����p]��grk�q�=ô����º���Ģ�[�����l�����G�	����;�4��ǀ�z�=�C9�ᆷE��Ƙ�>��!� Xv��_�`���<�o��l	�ٚ��wM�7D�9�ۼ�O[%6{Ь��=����Sf��JZ��E�zjj�noi�H��w��;z��z�O��CfK���z�'r6��;�x����ٽ㷠'5z��w)������pհ=�W<]y��-T�F:}�v좟?z�'��K����h�@����n����OC"����ؽ�i�'�����6y�	y��]m׋�V'�i\aC(V*Ŋ�"��T��]P���UA��QV�bTZ�8ʭ�F!���
�"2ڊ"��TF1S\�īIE[j��1*��2��#*娬1�X��]\0Q]Z� ��X���YmQb���1����G-UV"�V

[,Pm((�PUQ����1R#+X* �Q��TmR��YTm*&3I�2���Pb*��
�)D[lX��2�h�Q�L�����e���cQ�ATQE���Dc+%�X�6����,���-�Eej��V"-�e@��UU@F)Z�A���JKeAA[C��0F*��e�)ZȌU��֡l��PP��l��Z��"���(��6"�,[i��`�U��* �(�eb��R�En�b��P�U��Ub�Qm�D��b�m�V�b�ilR�A���[dQQ���1eJ"�DF*�-~�O5����U����NG�4I{$�3�=!0��/.ƭͭ�s=d�������r;&�=��fh�G�RM]�5�#��U�&p���)L�w�:)У�3�:���hё9w`	9�D���n�n��ǰ�f3O��!ע�ϗ�ݶ�u�"��yݺN9Ǟ긳�c�Y(�&����be(���z�]� �6W��;���w�r���7n�������-3�L�RBE��� ���%�ҟgzω$�ɠO���nŃ{��U�e�:��t�R��"
"�-V�H=���A1�N�J��1�{Ēr�Ov�vN���D�)L���1��n�g7���UY~$�}"�>��Y>��T>��ȟnݮ.1���BP�R�a�Cb$bh�䕛P6��uoݳs�/)㈤���AG�)���ZE�gf�걦�pkl�d�Ͻ��>9ϵ�_ޚ+ڎL�5�g�����>�yv*���N�j��	��߉� �S��d�+��C+�Љ�
����jڭ�z���[�lz�9��᝱��W\��Kf1�_��>��T�S�Dw�:�I �SʰD�,�Mm*Aփ[�4E�B�eU�$@�EO�P=ӛb#��ۊ��QyB"���E�vI>=����J흃H�|^����?Zg�d�����vI#ź�>$�l�Ԥ�u�"�����$�S���ػE)%J$�EJ>���V�ɂ[8����#��ՒI>ͮ˰���F���Wѱ �S�v/wOA�(JSd(�aV�h�	!�m
�3����od�z��ŒmvP�O�]t��P�%��b�T*���c�9��!q}���܂�2�a"��99u��ݏ\�����㼴���O�˴��.��WN�9a}��E�M�("&d�$Նؼa��+Yl��:����(6�1���o�-��ۆ�'�<]�]�� ׭��sk�9�;v��[h�Sc[��=��%wrՎ�PxyȚe����w-�
m.�����+c�ݠ�Y{n�]q�]��㮨�q��H�텹Z�1�����k��-d�k�N.:2��i�/m��Nw��>����9W�(3�DFٰ]�,�Vx$���:h����V�mΎ�x��z���ʤG���>vȃ����_����N�<�de�M�Í���s�Y��b��=&}�2/�mm�-��p���m�@$�u�b� ��MH��W��\�5���$H�EO�Q�9�d�6몉 �¾3Օ�gd�˽�O�'6�/�$��M}�U�R�>��)DA���Y�ͩ%�R�	�9ՂIf����n¦q�Y����W}vCqv2J�IR��k�Tc�Q� ����ET��E�@$Mo;�I'grh�{���q��#6�d�TI9��Z���6׋mQ�'��q�]�=n�\�d]�a�J��=��)L����wd|C�ʢ>}�ؑM�j#.7e�����9/&�I�Q�D""%L*�yw~$�;�{�����"Fݨ˛�"�ۉ��8C�E����Bf��x�gy��a�v��O+�G����+vw.��X=�`��0�_�������I'��&� ����2�F~]?M�E�^�2�y��I�ed=��$��΅�X�V�%�����bߘ9/&��#�[�"��PA�$D���y�kɁq;Yem�Y}u$�O�m݂A>=�yAuc�kEx�	���ɮR���ĩJ"؇��g����r�no����d��"�>'���vA=�ywBFYbG�����w̆;���d�'N�a�,��'��F^ܯ۱�u]�e�{N�B__?~|��bv�e(�9��N�7B���˿E���K��ՙ�ݒ�K��W��3D
��� �ػS\t=W�I'ݯ���;]��I��8���w��`���DDHFL���>��,Y$�ɓ��}T+���=H�HӢ���r-�3��N"�����L:�/���_�	�F��ؤ:��99�kn����h���W�#��}�$~�yvG��&}*$PdXf\�mi���u F��аI�ו`�F.����{Y��z����ۻ�9B�H���(�[�ڲN���:ވ�W{W��
��d��ח`�1u�Qv�vG�CGB	)���%b<�� �,�ɫ��X����3:�5 �)�������� �������$�^U�qu�P=��pS:�m�|��K�/k������N�|v���*Kݡ�I&�v� �Fw^]��p��Q ����0;�/p�yFĤ�dD@���h�3��$��trv��)�-�v[����łN.�h�>�E#�#C~�����:��g�`� i�m�$x��o Q#�[���H�7I��*0k����8�R�VT9��W*�,����f�V�zr��(m�r�&�����)��=�˳�|;Q�ɤ�rj��߇��E�{�dp�B`Ȼ<i�	$��ϝ_�Ѧ�	8K�f`m���j�e�E@'����:~9�O˽2~$��G�#41����yЮIܽ���z��+F�V���u��߿��[��㷔��>:{2� ���n��q��(�8(�g+��'̊rl���31)DA���L&�Ev���}M�����D�ݭݒ
�<a�����m�n^� �#ph������_�0��H������ǝ���[y����|�Z��H#2%H���c��om:���I�{t$���n�� ���Y��f���%������""Q`Ӟ˻����+����;���}�6����H$n�ؑ�,��>�"�q�J�tW
\�4�v�����Ĳ*պqu-R�uU���YT,�wڟ�7W�_��f�� %�,��5��{�����׻~wB1\�#g��T��\���zݹ�vs��<)��獳Þ=�q��gJ<���]�o'3��[=sl�0HBn1����w h�r�V�L�;��v:��󇀸:R�n�ے�:v4m���3Ŏ������=��l\hβs���'�l�Ů�����-���q�[lq��8�d�bw\>;s����1��y��wRn�.s�
��.x�2����Nz;��޶�m�7Tk�[����tvf�+���U�����|���I�!�Y�U ��� �7yw�Ѥ�m(w2a�	�ۻ$
Bt� �&J�" u9ݲ\�9YuPb"�I�NH$|�݂A���%�-����Fu�+*F�Q>�3�Db;;��$�yb���uI�r�	^C �5�vO�<�����7�E�dF��^�<w7��}�*.��ں�|H��וd�� �=o�۷Ӄ���zL;��r`��b$%��w~�H�̩3�����1��B� ��˰@'f@���F����>��h���k�Ɓ�r�-�N�՝fx�nnx�$�i��{װ�!�21�5YU����*� �]��ٹ�]�~��w~$���X�8E�f��"�2�4�R��ǑG9�YمC���'rҋ%�ݠ��8�{�j]���(c����q7�pQ�Qkz�_WǼ��We��[���2*�������w_x�	�%���� �1}�&a&��ξkj�'Ԅ�A�$Lʈ�E�Vز	OfT��onǕ�������w����2(�P�Jg�fbR��w����i�<I���,��Zy�@�kw��S����NE=�x��HQ�(�DI�ܓ�A�m՝Y݁�1h��n�v�ē�s"�>'ϵ���˷Q��g!�������ݮM�;P�� ��WNv���[��r��r�؞-�7����?��"�p=���:��I<w2(��[����(T��9�m�kޙ>��Y�ϰp�F$�� �;��G�G�Dl��p��-������ĝB��,aXP�>����AI�
G�#�}�0��|��'����w��ͬ�M�V���:����� ��a�2%H�L]:����{͇�AH[@��~�g�`V�*g�k��3Z�������V���U�U{N��T-=7��j�1d���B������C�w� �i���ڝ;���{�x��vU��~�y���*eO3�߷$8$�Q��=�gXv0�9M�򣤑3*"W��>��������_�^��4��VJ2��w�vr3l�e@�T
���xu�ѩ!KO�翶'뿦sj�?\tp�<�ED�W���H��:�&L��C#����#�����Ͽl�I�=/|<翛��?$�}��CI'�(������AH,�S�y�퓢uӾs�/�kO����޿�������F�g0����F����X�G�8n%{O`*u�����v����������~nHp��������v����0*S�y����@���_>��y�+4�7ﻆ����RT�����>�.��QFbB�����
���;��H,�߯���nq�|�͞3��@��}�:�X
#� �����1����큝���m�0*?o���\����s`T��y���@����2T��{�gD�B�+
0�3�~N~��þ�����a�
��T�<��}��N��X��YS�y�퓩��><ִ���F�0:��z����7��A�[���v��`T����{��u: T� #�B߷k�Cy�
+�W}J��m�O�|7��@X���`�܊'	�aT^p@�j����w��!��x�K��Ok6��&�N�������?�J��k��~�Ԃç0��ʎ�F�W.�i�#
�w�y��ID+<�|���hX>��gw�|EQ�"���J�����gjAH[O<����Qo۵�Dx��ۙ��
���ϟ�rnv�^^��7=N�C��lR;^-ɰE{�\�2a ����K �d���̣3_���|����T���gRu��#���~ݿ
>�#��]/7�>��_RT�?s�βted�*AO|���N������r�im�n����P�^���|���R'�NI~��i�ʴ`V�K��w� �AN�
�"߷k�$y3��"�[��}���0�aXY��>��i-��E�ra�¦���vC�(�d��|��g�d���?{�g~��_��yy��R
AHyi�w���i �B�����o-�~	�35SNp
�I���ݝL���~}v~��O�4̃%e*k�s݁�:$�(°���rH(��#��Ϻ�z�tڍ!��{�H��R����tN�_��<<ִ���G�:����G�i
Z�{��/�D��뇶x� �>��: Y
vD
ʗ�;�p�82T(��}���>|�>����,���љB3&v0��歗�N�E��!�k�U���gǙ�G��܋x%+��3Ol;������sZ�	�s_3�����	�63�(Oaž{괫�$��m
��56�IO\Z<)N��7
�`Ȩ�["��肽w���"aje��ڸ=�,�f�`<��[ޝ�8�����O�3�"�ozNˁz}��ۢ�W�F1֊\�5��%�=`&��z w�n[ʚ���w�d=XtuzY�|�{�����9�&�&�m��t�<"r�����L��;�n��+7����e�����K��oۻ�l�]�=�z����E�k��W�t{/,N��|�e粼h䛺�����H�^w����O8�WO��ߖ��c�ڶW�������ݛ�'��&�<��f�D�ۓ�+N�F���n���լ�����*���2��]�i��u9|;��oj�J�Yt��Y7�K���B׊q滨��I��CH��Jp�FNo������;L�)�c���/��U[G����N�]:=n�����,z��ʋ~8㎈d���Vww
7�m��(����Rz�v��o�K��A.@_tK}��/&�.���Jz�k�1%�x�=[Zj�25+]N~�x`���Q;�z�0���>N`����ۻev����h�ޞ�t~�6Fs�����~]=^gFV��Q�(�-��<�����޻�m�P�&΋�&!�q t-΁Zƣry�Ea���X��$�.�]�0ւ���'l:�&f�q�.v��I�p.�ՠ�2�PP���b�����TTA�
DE�1��m�Kj�%�X+EE�0`���T��1�EH��"(�U�,bT�VT�QX�#�e��5���RcYmY���*��Vi���G-�%Ku���`������UDV�,�b�"��Ma��E�̵X�KKUb�A�Z*1�
��*�RڰU�PE%j��&��r���ATV�0�R�Ɏ���h��Z�DV"�J�UX���Pb*i��,��b�eEȢ1b�EL���AV���5(��6��(�6��+�7i������`���Օm�Pĩ�r��������bR��dUUf�*�1A�B�QH�[�X��E��ֶ�M�n�HT4�Z���jX-,E��lƎ��Tm������\���m,��m����}���F���V�O����u\��؛8z��8�l�c��]]�m�]���s�6u^��7�Su�{Gk�xyݍ�g�E�=�q�������c��=�FA�2��*�4o���q��]teѢ�cQz��ܮ7@'[<�S�o)�P˽D�
�Iܞ��Gf5���c����qg\�y�y!��v6�bE�h�y��ͭ]���q�.�wd�n�N�p���K��{��=��ny���ʆ����q���E����y̽��I�I��]�	�z�r�<]F�.�d���h�;f����̀'2��3���{zS�}^�Gָ���6�&Gۋ�]��eݒ�������/#ȣ�>��)���>zu�fzv�q:�Cѹ�/;�o�����ċ��)�e��G/�i,�z6,r&�s�u�z�v�nClwWQ���j�ێ%��v��\��θ��h��x%-�C��IS�׶3��9����[�����=�{I��ޭ�4n'�Q�}k��7<��V�n�m���7e����xK�މ�k�-��G!u{];
�w0i��
��ѱt��V��|s�ks���Yv�c,9䬫�r��4�n���0q�,��%��b����Onܹ+qn��Yzv[�OVy� �v���Ij�pI��q՗�9�vD #K�p/A��n�L��o[#��p�.�gc.�]��O'nے�-�WG�ן�lk'}[g��N�u�s��=�����E��>i�Z���muΚ]���e6K��.��&͘Ǭ�qã�X�v]n��s�]OU���7�Ӄ!�;es��ɴ�ni�㗄z���,��7n�h������4����t�:����=�A�M�.-�������u;m���]��h��R�8m��=�S.�<u�<Ѹ�'X��z��p���7I�e+�qN$[�,�zYs����q;/;3C��:��pxp��F�s,�ϧjpq���guq8�]u�s��q���it�k��Z"?��yowѹU�.6k��N��Km9{6ݸnq!øs��;G�sێ8|+�v�[���G������NQ�uW�~߮�����v�}�㭰�pun��\�5�k�46����,���j�y�a�]��/n�kC����Y�p��:�]��� K���Uۋlf�fH�v1u�l�g&�N�۔�8w�g��s۰���붅�`{V.RuO3��`Nq�[m�0�:�y�'n�����:�zyd�t�e����7i4k5r��$���͇�!Ԕ�����m �pJ���{��0:5�U�W�ºs��#������c���q|�v�(�E�u����#2e%0�S�5�����YFJ���~��_�I�������� �����ra�%�T�O���vu����߫������D����@�=9a%L���t�5��w�Ãą����}����E �>?(���r+��`O�( VT�y���p*A@�|��a��|��(q$$�$)	@�8ã
�����k���k����N�+%X>��6����@��~�g	�	��h95��]�̌�������ۆ�0*R����ʙ�Zi�S�O�����u��VQ���sݠ���"q��Z=x�nf���*J�Ib}��{���������#���0��j�bV��Dn�OD�f��E��[���x���^W����݌�ԘRw�e�P�2�~fJ�$D)>�|߼�6�R-Ͻ�ݜ�R�
�H_u���$}�����, I��1�H(q%B�~�߽�Ԃü�8r��֜�e�9$���͇���W޿���_��"�X�%��btN��� ��g�g�Km����C�s[�z���y���+J�ԇ�.����Ft��������j�+��"�~���vq�Ѭ
ԅ������;H6���ϼ�n�t9�k��O��D*����3�fD���0���߾��u�Q���s��:��T��aX}ϫ�7����������i ��
�����ݝd�+%eH)������:��PJ )�R����_S�>����M鿾u��C���-��<�Ă�^�*y����8�*T
ʟ���p����571T�����"<���[��Xy��?f�۬�t[������?}݇P�J!Ro����'��������;��������������R
B�Ow�߶{H6R���;�i ���%E0ty����#ND&2K|�	�e�v��W+�^:r�q�Ͷ��͘wOOn��P�����ؾ�3Z�Ӟ�S�I���ݝN�VPd��%O7���u'P�*AaO����I�|����?B�4G���{���VJ2�VT����d�@��y_�5�7ZS2���Z���9��� ^Hx�U��WF�, �����|h��O��߸R
Agb~Ϲ��I	*wo[�f[{���C��6|���aNg�5�5�p�CI>�{���:��
�YXy~�vpf�
 �@!��Jh�65!S�(*���t��>���g �&s2�N�:�W�7�w�Q�N��۞�`��{��=2�?&=���`����W˺�]���gH�y������R���~�� �B������o,޼�~2�R��))�`#��P�"7���U� s>++%N��}�ԝBĕ�aX>���a�¤�T���vq���^�*0����'ް�]��7gl+�k5[tۧ�`q�}�6$-��	 >o����т+��U��.7�u�
�����N�H,�_}�w����D�
��{�:ì+�{��7�}6�l)[�*0�A鈘A0v�s�<a��w.�[5ڞ1�sjܸ獦1~|_�Im�h�-��z��My���;�J!Y++�9ݜg(ʐP=��}�dx�%@�o�"%���}� �1m!Z���{�m�����*f�i�6@�\��8����Vk>�6?v�>��y'�}���IԂ���/�{�Cl8¤�%߽�ݝd�eG�>�,�O����c�~#{�6�|ִ�iLˣ�R��͇�������}��t�+Fh��������_ݗ�����@��@��+�d�X��P��}�gXtV9���@ɓ*&!@���g����oMc�>|�:��
�Xr��ۆ�
"T
~��}��Z��R
}�}��5�����J~�XmM��h�XNw�/lC.��+!�Bc]�kv�V�Y!�y�wf&*��Jw!�
1�x�����2���˘��94��=?��#�����p����w����u�]h�n��@Ͽ�}���e+,d��=��΂N������y��+#
����na�%�,O�{�:�ѕ���VT����a 8u����~�衉"���B�Ѹ�d��{Anq��W��q�+��y��v�B�l�EB�))I�#�>o��ą���<��vs��k�`Rݝ� �<	}�Q%��>˭ #�!W��6�2T(��D;�{��:0�)����4��f���9��¦����u��VO�:7�Ͼ>�������=g+*A@����`u�
Ԃ�{�P1��Eګ���O�L�����c��k�/�r�kV�s�T��y����Q������:��X����>���MFgN�������ID��~�gY:��FT��{���u:�C��-�Z�u�3.�`u�y�6?
?nb[�>[��H��$ ����^�
�O>�}�N�T�������;�t�Z1�����A%B�w~�ΰ�
×�����5sY��4Ã
���<�u��������}�Y�Z�aQ����������:5�F�,����݁����h����nx0*d�?~�����	��G�Z���5p�n�d��8��7�L���G�cquާW���8�q�-9E[�Q7v���k-�0��ɋ�������߳��i���f���]Ie�^�d�VS�i��M�q��`8�ñ��Wq�6���z��W1���0��mW[�ۮ���۟s� ZL��L���ËU�q�b����{>�t�Z���<cn���b�l�;v;pU<���纗�C����<n:�\wb{V��ۊ��$���]"��۹ #�6��j� nW��M�ksѴf^����`]"ι�µ��γ\nU��>;f�F�76����p�+������^5[��'�M}��l�t*Aed����Τ�AH,)}����q�I�=�k�����>�6�i�����'FT��S�;���5�����cn�t����]f��Iu�q"��ә�-����S�{����J VT�����l�2T*J��7�s>�:�_�8�0|�@v��lϒQ&
P/�u�Mwϻ��ID+%e`�����g+*J�����z��������?`V�,���}��;�A�!Z!}����FJ_u��S5�M9� }7�B�UG����i��>�>L�9��ݝI�(���
����a�¤�%O���vu���wY�Y=�����|��c�r��֛�)�tl�ư}���6�R-Ͼ���x"�s�|�GQ����C���:�� �}��6��
$����,�`>�5| n�r��i�l)�;@뛝C�G�.��'9��ȋ�c˂���R�U���{��{Z]j��u��4��?k���u��VJ2�|���6�P8%@��y�:�������k׸�SY���8��h���wp���R�ߟ��]jWZ�[�xS�5�����@G�����B��g�+vI'�K��j�a�=^���H����ac��}Au��J���OVV�E)�:�w.���
�bɑ��'c�%w�����S��l�uT�����;�m �z������}�|���;���)�H�:�F�1B�*`%&�>��>�- �}����)
сZ��ߵ�b����߷�'� ��{��g*%B�}������~���|֋iu�U�C�3Ͽsa�}볩��)=����y�m��*�_~��xu �:5!mS�п[��Bc�hx"�
~�
x��ou�7�kV�s�T������:�*Ae��>ߞ��ԝC��k�׏����ϻ�����/�<�!��*J�Iby�{����������m`#G����$�~��Q2g��c�w=f�v�gC+��\��LZ�c�m�eNf�32�qlB�bB�$DL|���z�8<HR��=��vs��� $/���� DO��9U�@|�E����l��P�%@���gu�aNg����s5��i�T�]�͇D:��Y?{�{�-��w�`�>�g�d���@���{��;�R
}���!�PC���@ܝ��^�7{�m�.����ni+�i-ռ�Ԛ���l�v VVJ��S���흂N�RV�`�<���i﮽�sy����g��DaZ�m��_l8��3=Q����n�.����Y�a�c0�,�����]k��F(\y�ض��6p㳏n����濡Ԃ��
����}�βu� �Q�?��߶N�u�x~�ֵ�ȕ(%&�>�Q������Egv<H~-!K@����g;HV��Z����� Y� ����>|�C�3퓩�{�ΰ�aXP���e�ZGZ5[p�:ã
���;��RQ
�FV�����2g����ޛ��j%@��~��;�R��������A��h!�wP��G�{��6O�F�<�I����7�^3m�s�u'�+�G�U��bK5����߿����s@iπ����vu �td������ĝBĕ �������aR~��{�}>��ӟ��x�������Y(��YS�<������kw�s�]ZS3X����=�<�q�B�H2N��}���=���w�< �A;��w� �w�4��y�<������q ���kw�.�t�f��ra�§�����;+%ea�>��%e@�T ��5?}7󻹨?��| ���$)i��{�`w��aHV��u�����Q$)S$B���`#��?�a��Q���x�>�"�~��=�
���+��u��aRT*�{�,�݂����'�%@1BQ7>PH�Q97Ӟ5��������ST}=��X�]�;���2E����/�ިs�������2�VT��}�`q�oӼ�ֵ����R�����!e�� ?7�B�<�y��bf��H��=z��M{�{�:�@��%��wp�82T($�Q���vu�XV�=ʍ�^��G�ED�@T
h�D)A%�p§����;��.��ڳbx����ߟ�����ڭ���8��Mw�{���K+%e`��;��8�YP,J�}��}�Ԃ|�T��vl�H}[�@�<
�	����;�m �%�^#jf�Y��18������t@����>~{˞o^'��'���}͟��Bĕ ����w��*J�ID��}�gY:��c+=�G�9������2�6���@8��WE֔��;8��X>�nHp���>��vs��H-=��8��ï|�
~
ʗ����iD�߽�ݜaхa�ٻҗZ���ᛆ�
}����͜Ӎ����t�*O�B�X���߾�6��T�S�������Dx>�;h ����c믭��+���᷌
��߯Ź�����V�'Rk߼�gS��+(2T����3�{_�^4��"��>|�=�y�m�#
��RX����vu����>G�@����@ 
�U�g�NR�v����R^�y��E9��.*޹ǘ��RNT���m�JKQ�!�՟���.0=���7K��kw
V�������?�:hY��j���9V�x�����q���;s�u\�k��s������s�I��mѥ�v4��N��#Wuu�S�p's�{��N�]Vv%7Hs�;H����M�{\����P�'��E9�#��k�s�q�m���m�h-���]�\W��I��l�i�h�P�Rs�`�;ro)�8u7���ۓ�Mƃ=�FВuf��gskU���Cm��G�x��w<�
�َQ�r����y	�Y�)��d�����|��@Y������{��}�Δ�k�`T_}�� �0#��s����Q
���6�2T��C�y�:�X}߯�u���Z[\70��Mwϻ�8�Y;uӟ�����[��m��y�����P)�=��H)!�O�￶{H)�ߙ��@��u�E� �K��5B��j�N$�}��:�*Ae��>�����IԂ+w��u�~ӿ��yÙ���m��*J!RX'�y�:��VJ2�X2��s��'S�k��s�]ZS3X���X>�l/���k8����;�~�g:R��Z��O��߸R
A`����6Ϲ���[��?$:����vu�XV9��xau��.ip�CI=�]�a�IA
�YX>w����2\p���o~���(�~�����A�
5!KO��߶gi ���wp��N^���~������������v�sʼ�E�%��;�z��x0U�+e�ѱe�����󅎑�����My�϶u ����2T��}�gRu
$�,aX?��w��
��qӞ��9}����bN�ss͝d�*Ad��C���R�b� �
d���Dx�k~�M�༐�ދ�s��>�W�f��n��o^}�y��5��3]�e�l�f�q/�S�u����D���"$�0�ƞ�w��/�
��оC���AJ{�?�p�P*X�Yb_����G���"<	6t����a�j�����aO߾��kQ�ִ��rH)���l$�
�c+��ݜ�J2�T��v}��e�����҈�$x5߿�i
���wp�AN_u�~�DLR(T4��K�v;Ng+_�����>d��9�vu'P�J°�-�����F%�('�y�:�皷��_n�?i��"7�(d�qv9残�)��xu�ְ}�<�q�Bʇ�H �ﺅ��F�*��r�p�()ϼ���u: T��K�~��q��,C��ݝaхas����>��e��)^RՑ��Wn;]
1��6�ݻqoG]��㮞Y&�=�_������,������*}��{��RQ
�YX>w���8�YP(�Ͼ��xu�Ѭ���������$}��b�P���wp��������35��榮��N��߾�gS���Vy����8�����ܩ�}���Z�6|��T���/�����q�ID*J�}���'c+� |���M��Uo��ߨ{|F���p\.����X��ﹰ�<H[H(~��vq ��
�%ߢ?�ӿ����WuBb��qt����78���n�zH;<�𜏟�v���$�c�~�Q�AOyS̝��e���/��z	V��--kў>˴ �]װ-8������tWq�K)�t�}�tN~�ޞ�î/j>c�'Q�a~��U���=j=�ܫܡq���ᾓz�<����ν����H�d�o�܊�u�������θ�>�Kj:5b^�h����Qwq��z���k�������(�p��oTL��M�Ľ��Q*��O�� G�%��=�N�<~mf��/�X��]�{<�c���s��Q���=�/�ݨ�/{ذ��AjSfQ�h�:�����!��;�R�Ҍu��ǘ������kA)lғ��=���yjhnuQ���M���z����T[�R`��zIz�L�@ŗR����zD�PۣTwE�E�z��S�	�
���;封Cb�xt97�:�\�W9^��@)r/�9�q��|Q=��Ӻ��ܗ�;^޴��Fh�x-�ż8]儞����c�$\~����q��������?f�S�`Ƙ�_������f.ME�	�ˋ�;��1�(�k-c�C,fӄܻ�r50�J�G������(=���m�w�DL���0OVj;ä�h��!��&�{��2�9���*�]�v��f)h���%<��n���!;��]�ju�B�&n��k`��s ���{Ρ�;x�.�"�S��o�g4j�+���A�0�:�7�!�gY0Np��Qg���>S�l�3W�N�Yh��y�bn��x�|�(��)��1U浆�����m��Q�
��E�ZEc��k(�" -�h�V\���k�U��Ey��L����c32�ce�BT��"
0Z��;�P��PUA�QeC0n[�ծ��J(i*"j��c�6�G,�Kv��#���1Xi��T`(�m�n��PQʵ[D.�*��lb�TQs.
�[�G3]%"�AmSL1X�R�+cs0ݨ�PE�K��B�������T5cJ�RҪ�("�F �AA- �J�Keb����k�&9���TsWc�R�QV
�Pu��N�a\jJ�b�T(��!F�UE��PUƫ-(��ADm�i�(+�)L�M7Hڪ�SH*%��U�ɂ�0յ�luh*��3-��4���*J�-(�0�feȻ��"����Dbȿs������(�YR��;�m��%B��}�����>���<���ִ��9��y�6�k��}῾�ǳ]�6���e`����8�YP,J�g����`v5�F�,���{�`Z���?w߮��ސu)
�/�����
�����\mr�.���1�}�l�~+(2VX�S����/>�����_n�'���,�}����q�IP�(�{����'c+%�+%eO�翶N�P>���M\?�p�3��6PE�_��)=��뵋v |=v�y�'��L��ƻM1����~�~E�v�k�0>k�s��iKH[@��~�g���,��{��u ������W�~g�_}߻���d�X��D;�����:0�(^j�8at�W.hp�C��ծ�G�����{�w^_W7M�m����g�8�HʁbT<��}��cX5 ��s���i����u=�Y���y���(�>�X�5sXi����v�&����:�@����d����Τ�%aXV�g�oy���f����ID*J�}����Ad�ʐS�����'+��sEn�� �w߷���{���7��AH}h�>�gсR
{�=��8�@�beK��wp�=�{~�Y�����P7",��\"�5�º����
"��Ly�e�^�ٺ+���[^\�y6�1�*�δZ3�hŷj�0�Ќ8���ݻ��E�F&%g{�@��@�{�gu�a��o��.7Z����8�S9���x�RQ
�YX>����8��2ub�o�#���>�| �<	S������i �B����6�`Tl�ÕD]}3��%*&d�� ��I�櫥��<�\>�v�m�s��<�Wn�e]$���|�nٖ�)�ꚿ�k��g�Yc%ed�����Τ�V�ag��ݿ	>������;vl1J~�\�մq��ed�� ��9�퓱:�a�w~�|�h�й�ǇX�a��<�pv��
�������w /�e��x"�|*0*_�s�����T���������RT5�լ���<?h��g>�gXu�ae�ǆN�\�3��T����a�:�R/~��Fm ��@d���;Vv}6V�1|0�(����������i��lC�w��H)�i��s55r���_~��O������s���x2VQ����蒰��a|���CL80Dyx���#�}�0�ع��q�yq��H,�eM�����������\.h��°8����ᤂ�P>��l���*�_>�����|G�!
�̰�
�@���w�C
IP�{��]>|��[�!��}9���DZʉ���<��etV*��qx.�����ކb�9�H��!X����4�:���G�{gt.1ŠLe��?�ݥ��ۍ��٤礊p�b����tہ
��0q�{Q;.��zڄ+u�pZ���NX]�v6�g\��λiQo9��^���7[�.�M�Q�i��u��O�X:_��a�sռ'��s��0�%�y��ݕ݆��t�wg������w>���B�]���#]u�s��g��y�2�2�9y�R&0)֖�=���uj�W�g^G��ט;-m����wU�[Sf{�I��l��J�z�:`�!L�)�8�~�9���u��VJ����4l���$ �;��c��|��W�Ð��I>�>�`xv�RP�;桎����&"0��(J�d{���F ����9��}�9y�w��ݟ�N�aX_s�n�l*J�IS﷝>�#�/#�foԵnbTؾK}$)����� R��d(�LD���Z��h6�ZB���͜짂( ��"7ھ�*5d<݉]��R
Ag�~���c6�P���}��|���+y�q�ӭW3CL�1�>���~߼|�k/AH)���h�f�(ʁ`��{�8�X�G�	��� }}�u)u����G\�A�sC~��dI��J������'�ed��%O}�߶tI�<�zɭ�ly�H
#�H�����Gm�ƛwO�;e����r� D���R�Fu��.�\�7YZNSe�q�J4g0��v�'0���$�
%���9�nsڰ$�u�w�U�9E��j���ݏ4�j�*� )6�_���E;�"V���G���Y�٘�H��4�ٵ!�GnW6D�t�{s�dd�J�T���_R]AB���h�����H$��ݱ~#�vP�u˷�F����yX��]z	QABDJ�{e�݂@$�S�	�6!ɻ�u�/7�	�۰I�e����&�,xhI��-��b���S���וd�@$wS˰	$��B��qk�\�Ug>i�ϦȔTU3J%���߬�O���y�ߩ�;$��޻�1�e�>'�/�L^Ek]�5����k��rfCh�uVޕ�n��4�lD٘�'U�4%4���$����G~�_������]�,�I/�A��N"��]ꑄOv]� ���]�3��d�D��@�Ι�-�
�.�ψ�˲A'/�HT����]�ڵ/gπ��j@
M�{�b�$;�@$�-��g=�M��4-�-W(�a��հft�h�������Θ;��r2]ᮛ��h�i�]�=d}�3=kL^�@�홡!�_M��C3nܹ�s9�I'��.�$��g���(��3������ߓ��\��~>.�H �{��f"yX03$��]�A�B?!ɼ	�hI���^1�|s��Y�7o�F�\9�����$�}H�=�
��Fd��`�U�	�)�I�Ctz���7l\g��r����%uQ-�c�;y�� �3(�H(B�s'�Y$���$���j��1V^MW�=���jv�����O�!]�����̓;�kb�V$����#��ՂA��ѧ�H�S8N�d��h�zђD�RMX��A'�^ՐA�ѐ{o2��cvw|Hu���#{}�����"$�� )7�̚��`�
Y�*ωtd� ��{B�$�}�'�'��J�]�2I5{E����S�V+4���'	hK$����;�w�5����$���s&c�B��[�-��R�4-�>�q�F�M8^��DBF
��%�]U�${���j�r(R�UM�D��q�ڲ	n�)t�������x�:�#Ȇ�ΐ�j��F�h�����vqL~~�q��{6�g>!�L�A��`�Cw}V�t2���D�K�ǃ�{�f�W�1b�!'��Tt�ݒ�޾��d��|�j�H����/��]E
��w0)��陙�J���#v!�v,���]�`�t۽���F���H$}o�n� �w}w���ђD�RMG8� �gjo�n_uY$��v���'د����DNʼ�$w_;�Nf�щ"aD�E)l�h$�{"-���s[k0d�F�/{:���ۻ��|��<�޺���۟�;��Z���Cel�7�p^ȩT���"X�RI�Ƙ�ۛɪf��.�T�3����ݾ|L����w׶��~s�z\.p�`띧���G���n}������Z����8*�ܳӚ[s'#vu�cc�{5��C��]�;;�&��ѲY�X#���Rںb<����pv�q��v֓�s������"v�L>v�q7O�F�V.�w4]�-��Ն�:xy��5���nW��vxuq�s��魠9H��mϘ1�$�ղ<��n�тd;�듮:�ܼf��v�{u�Z���1���M�?��{�ʆqs�'Oͦ�v������۽����i�V�z���>$��d�+�l�I��7e��=�Os6I��R�����$�yvI b�R	1�L��0�{�r�`US,a�x#��2�'�|H+��+�M��< �w��z�_)�4�O��o )��"߯���[1���/��u�e'ح� ��f�xwUs�bN�ӱ|L�J@Pg�I�h�$�{5�Y�oU��/o�F��1���u�'U�$���n�X�MO��D�І��������M��2G3�wm��@��5���L�ɉ��N9$I���JE|��v,����`�K�v�g��y�9s� Þm5
#��(Y�{�RR"�B�S�'�|&}s`^?����Ǐ �u�l�f�ش��;A��Q��gݲ�;h�f�*IWM݇�b]��V�����=�o�hW�����o�ݏ��
`^��aT)V��H$5mH$��vO�E;�}2���s�gnJb6f�(�7~,��>;�ՒI���F�k5Nt� �W�O��^��*I��P���sT�uh�����RA��ۿH<ﳪD�{�Ś� �7Tb":A*'���ok�d���u��Q�֛7HI��ڰO��}�/�m'Yw$N�c���Uѩ��(ݐ�%�����뱳e5�#�)��f�k�)@�
�I<h�L^k�	�w�w�ǨM.)Fx�R�|{s&���P& `PS��V'�a��sE��A�on�O��}�,zh�z��m`#6��D$DLd�T:m��$�8�{�m�.\ⲯ���gҲ��o�P�Y^� uW��dc�VVdK7`��#��z��fR�W�>�#q!�"�,�J��Ll�Ŭۨ�H-��f �_e4ò�&訉���c�اn���&�~�w{�a|�9�S`$ꙸ��� �����?\����&i@��ug�VπA��U�,z��"������ A�M&@��.ڊ	Mo/��t��WBv�(����7]Ϟ�<n�zx쓮��t�^:ɀ*��OH�����m� ��K
��}?fR~$Dk�` gz��L��lU��˩�ծXZ��3I��4o�Eo�a (3�Q�>ۿ��2-��峒k3�7� G>�m >3�u`�C���yu�!�9��cؐ9�x��H��m?sv�o�Wa�D;�7\�1꘷7�$��ɢm%㝵5�:�?DBDD�FL+�����-T����Ѹ�� ����,���/���ʩ޾�/4SD�t�:���ERop�{�vv��m��/��.���\@�}�/���2�{��ަ���c�	"}⅞��9 {��Le�LM�QJ50����Z 3�u���כ=Gn��I�nj�^I y�My%��m��^�&����G;*�UP|M}UT���YB���ƕ�W�B�����!k<2�ߟ���L�&"ABv/{�h$��hR%%��ݓf�O23U�����D�{���՝3D� ��S(��'�ۙ���7��q8����ey��
;�u` �w7�ሓ.��`.�_���쌘HR�5�TC	��� ����������FL����g�Gv������$�#ʐ�	�$�HH��yM�S��Xπ����4��ۙ� �잱1b���g�/d�HE<�&�n� ��
�B*$r�6�٘��@m�U����c�o�7uD�IWky��P	 ��d߭W�5!��2ć�N̑Y(%ɬN�w���8v�9Oʯq�����.���\�t,C0�\̸Of��{pߧ�m����ͼ`N�a2�˞�Փ�O�S��~-����Ǜ�uo���zt�g�+9753AUg��o�0+�Hzﶃ_'u�Ǜ%�a�D4���lmH��ʹ��UdDm�i�Dob�-+�]<�r*[K�8�T�|X܏U��X�K���}��ۨl��D�h�Ư"aдV#P�h�]�w���������&���Y��q-�W7u�}4�9R�J�l,��跤�.+ ؊ʔݙ��X�,O6l���'�T��ɪuq.��W&�1H��lF��[�w��y몌����]f/�3��tg�}��x9ov�� �b��d��L`��ȋ4�I�@�!5X!�]ػ�3�#!v��·XO^��ׂf{��.�i]`����hQ'{��W3��{��z���#�%�^�ˈ���c��X�@�6�n�46{M���$[�|���t��)u�����F32۬[F��ce3q�:p*�{����F�%�7�ܫ��Q�uc��Z4�䝻/-6�����Lr�}�q{��3�ґMу�t�[���\@�����*j���
XpQW|}�-�7D�ȨwӀܾ�jo[��C����S�P�gs�������o����c���w��è�ny
��8�G$i�2�4h.��^��[��\͛�I�k̸bf�$�5�D��,�9��QL��vxu,�y��0{�������{V�q�{�܃��}�w�=Iy/K�J��I�mAV�qr�Eb�T`[E�(��Y-�Y�a�CR�Y��j#Y��-��Q?%`�ZT�TFc,k1��V�jTb����%\��PW2�ƍkJԩ�X(�h�R��k.)��#[�̑AU�1�X�b��J�`�V�Q"�֨�S&R�J�8�*!ܥ���;�ݶs�&���[&����E��k+���Ҩf �ț6���m��y;.��to%Ó���x87v܅�;�=۶��a6�9�CX��[
�i��\���xd-(�:AmT��Q��m�J�[��5�m�1[vᔪ;L�.Ts\��m���]�#�ݺAM[Z-wq�ʣ+DJ]\1�\խ�*�n��Z���ج��T�f�\2�����naQM�t�&Z�hk�q�xq�om�we��߽+�DQ���8�[��q�v�W1wanˎ�2v��1͝�׎�pb{����V;`�ù{��2�����$��!竅�:�������৭;9u��������5�;�\�M�;�q>�P]���7�^.E�c��-\�m�n�8��뷮�n�Ag��ꜞ}]���uٷeh۶aʂ�\�\��۠2�u��v�Wn�Tlg������8ۭn.���Q��М�=.xx�t�f)V�v�;qף.���e��G3÷�����;Sq����:��Ccu��us= ���эv�eznn�H5e���i۶UQf�3±���%I��͋mc�ln�=����Sm�A����@���X���Ai˳�H��L�z�77:��|�W&��7>��`���;p���^E��5Ky�$�.�v6�8�xy�5;��9�\6�w�jԧ0����ې��]K��w\��'��:������{-/Zћc������0Bn�% �WN�#�L�i݄چ�kgZ��.x�77�.FոT��[�x셓�]��t�b�����G5j�}]���j�ۡnwg�7)�� <틪��cnrk���vr�m���GSkd.緫.8�<��0WRԷ����7ns�v�f�Q7n���`������R�CO;$�����5z�uX�u�mQ
ǆ�v!������F�.�yg�V�)�5�qp�g�|��nw[��x��\u�ݻ6$�<Nb��� ��s�o<p�zl�[�'i�[���`��kJ���AGZ�.��&���0㪣���FI:��+���Fx�jw�s&�rK��z���s��bK��k�2�}�R��U�u�հZh/j�'�u��z�ku�p�6^1ڇ���nL2�s^�]c�u��<�L�oc�َ^=���]�){V��FۍZ����9�,ᩎ�j����qkggX�B��9����;��童�fH�*-[<ݥ��B�ٮ�ۮny8�z{��Mn�;�J�\r�A�3��&�������{�W&z�{\�Y�Z�h���}v^AԮÄգ���D�2u��F�Mڔ�v�k�b*�;���.����N�='8��K�lEen6�ɲa۱7N�].�TCn�u<��ȸa�(�*�0+av�0��7888��pӞ�<<����in�ۛu�bt�Z���V�K�u��(��ؔ�tu��vv�r����B��X�im26�����,�aM?�:�&d"��ۯ0���o��ѱUQ
/���� ���Js(%UO�$yޙ��9߫�uj�^���~a�y���_e6@���+p��x�K�i\A� �2D�"['sw3 "#o��l@|��w9Z�wVz��P������즘#ކ,���M}����;s���ng;{9�� �ܦ�Fo;��W�fɀ���3�Y���Q�H %C?sj؀@�wm�l��:�=�K���a8'k�n�A$ok����)��1lW�Ģ��)S����꺘ݑ7`��۝e�S�h䲮�?�s
"����U�����OS�d��>wV�K�FI~��U(����W���l�鉪*"iB&�,s�a*���6��k�л���	��=ْ/��tX,�7�hX�S����n�ƿ?�{8��e�ݴ믭��{�'�tw;����$��t�I�"���@ f��iB��#�������~��@kkO�$z�Mg�|��w GT��ʬ=���|� 7�S�2�Q��퀲j�J� �2D�j;��TuoՔ� 2I*ꦸ$J��n�I*�o���W�'�������C$�B$&���I3��o|�����$vc��#�ul ]�۷���x���Tߧ����
$�)J�
T}SB�(�v+x���=1�q���P����鿿�}�� �d�{\*�A ���i$J��f%"�����-���� G����{��J) �H��o��~%m���|�A1�Fw:������}��ń�wx��7�O�2�&訉���c�7p������n��>�����W$^t�D䅐�(�l�{�K�j6��MTB�4��>�k���	��]�<������1�����뽺� >Qݺ퀂/���d\��f��b$&��E�o0w���_D؀�<v�" /=��� ��sLQ��'�Y쬺�$�I�0&%L©�Kd�{s����~��yж���f;h 
�n�,  ���le��3��\g ��@DQ$�l�>�6��d����|�/W;f2�KH\���%������"�TC�'�s�a^�ן`  �z_d����{qNv�i��˷z�� +��3 ��O�UQ ����L�I��/)݅ �Rg�}� ��u��H�v�&��RNttA��wOkH���
) �H��s���N ��z� 3S���=������ń�ϲ�a��9L�T�4�S�����v����{�<�
��<XD �)��I���ޤ�G-Y᛾˅$���a��)3��,3�S�LS��#�p��v�_=��sck���+��˕L�����N`�� 5��BO���""���7Vt?��\�"3]��� 9�Sd�gv�����۩x�㠁L��:����ƣs2x�E�s���K�<M�CTVjJ&"�Á(�Tɓ"4��ݒ{�F�ʶ�@Fwk�J��u^�� _e?�${�ŕ�"�TCb}��]ZVz��s��ߖ D	�)�>3�]�O�γ-���A=���Fq�T�&���m?sj�w]Q$��t;�Z��*��-���%䗑�r�̃�gv��q��Ȑ�**d��b�{o�u��S�%�t$�;�����,�۶ݻ����^�n�&��2}�-0}�K��&�"ja�^6� Wv��5��E��Kf�˃a!��U������1Y�dw�ex�᮲˿9Mtc��辝�/�����D�e�q�Csv��7"�7"�3P����5��L���[sI���>��'v�]�~��Yֻl��R�\sk�����^�^��n�&x��Q��\q�e���ѱ:�ѓ&���ŭ`C�+ӐzK͹w����gi�a 6��n���磧�'n�ڜ*����Ѵ��n��V��t��+��`ݻ������9qM��K�I���)��㨻cq��!��]�r��8۶��#v��<�,p�����ݭzCq:έY5���d��M'SY��GBy��'��]�"l���N��jjt�~�~��m=Je�
��A�f�L ���`��s3�~W;���;�z}y-&A���v��̇ al0�%!_�w���i=�o]�ʣ{�SD-�۶ݻ��#|a�F���?W����v�8ʉ(B&d�$ݡ}�tm$�|��$�8��fW�r�/�!{{n� 
���Xx��*Q5�%C=�
�K2oj� �v� u�nf ��O��Gݡ&1TNW+��H�wV�����)@0�P�_���@8O��[�]LGD�����w�1�nf >>�3a��x�u����A51U�Je�[n�9�F2D��]{<upf3U��wgWkSE�{�E�3Q��ӾB���<�u��|y�Si�������f��^c���ۯ0#)�EJ�$&d&��=9�*ɒ��ʔ�ܜ}p����ү]/�>W�v��/]�����𭛨�� �һ����H�ˮ�G����`_�N��#��w=�W�v�g,R#��dӾL���2"#_e4�If�a�.c�u$�UBQ��&!L�z�ێ1�F�ƾ� z��=L����wZ ���XD@�y�U�F�E��D̐d�����+Mw>Ǚi/�3��`@���q=�u������~��{s٘މ�L�R ��?sj��n�VwY:�������f$_e?����ۦl�(ۂ�~@yd?�?�8i�p�����G�nm����r��&��ۃ	���߿�?{�ܙ*�fb���E{}������A��]0�~m���1��fa u�S��Ϣ�H��b�!Sh��m��<�я����}|1/$J��ݠ��v�i ���_���o}�E^�L��$��
�Z��U�?�{{m�� 5w9Xv;#k�������k�9�c�������
�O_zg����m�ˋ���P4�S1[�+c����)�x�R��IL�j���^ =}����k���ȫp*�QTT��q��^��S���@|w��G_;�H�]��U��h�S]�$�ܮ���'@����؟w;��H/������V߼�\G�:�)�� C�wV��F�y�bo(�Si������co̝�q��=l�q��+�D���;;��vÞn�3�tT����|���-u�o��}�ۈ.��D��ۙ�,��3Gy@��%��7�E$����#�8�6�A�ux�u��n:o��'�Ete��l�"��v���v�, ITig�Fk!Of�ZWƸB1$ML1��& ��^` 5W��Uh�u�aַ�N�De˴�I��D_{���7�Dʪ"I)@��AY���:x���< *��� /7�-�I$��կ1�}�|ټ��u���3��j}�o?{v5 ���t�9R���L�zw����9<���>���
�R+�:���_��+�˶�2*�
�AU$�-�{7s>X ��5;>zb����*D��鼺�$�:���a@ ��S�����]2g����n�=j��歭N�c-���n
6\򖶋i�z��Ad���}�o��ÃV�m��{��`�#ϻ^, ����z76;��y�:ї�퀀G>��X���򚙚�@����մs�`dM��S��;�|}��  A���H�	u��z�����jCwY(�&e��a�P�~�m'	 {}^�@ģ��=8��ٗ�9��b��_e5��z�WS14�Ss�]Uc�ܜ��4 ?[�` ={�m  H����[��*��
U�xI�w���.�S�R&$��-ug��@����d]��U�h�2�73 �_e6A�,�۶�ڄ�r�J���76W=��٨=��w/%ը�x� ��_��{�MKRފ��e�ʔ]4l�Pӗ!�b��k�5*�g���k�o����˘o�sU`l{\g	N��n��1�M�ln�6���[u���]�b�gv�'�Ɔ෷M��S�W:��dN�<q뱥�nާ�gcgq6�q��u��g��x���Db��ͱ�Ź�V�:g'U�J��9.�ooc�v�5�/&�3��ɮ��q�u�$��܆�X�q@[m�����^�< �v�q۶蓧k�����"C�^�9K�v�Y��Z�d�*���uq���p���L�m�x�x��Ϟ����I��Rb���)��0���_yFgvg�	 �+{�π@}��o�E�Uz�p��w�7٘@��i�����I�[�6��̒�ⳋ���������|f���0F-QּMnb�G���򚙪T�%C{9��?�o���g=�3ҷ/���%y)}�v�Ix��&�v�(�&fff�W�e�=�)��׫�$�V���"��m �E��sTK�Ɇ��?\P7si�Z�)��M(ET�|.�m�D ��kq1�2��V�mh��:��������ݹ�W�:�_�����k�Ϧ�u]��ٚ㍖7n{sZ�7UrNw�n��M�e�=6�����������#��V �Y��i��y��K��F�:�C���Y(�o%�A�
;��ldU�1�ML
F�'��3EFw"w�N��î�qS�)��1�9����Ӷ���4{<�WM��/fNi�v��i�9T:)�nD�������=8���S�FÆ�M��A�gw�� �������8j<du���@�JW�!����q�s�a~�טD7`�U�ݫ��4�	 }�D�IWo<��[�:"bfU)T6�ϵ�&�]FyB��]��D���f�AmObj�&�"7wjo(����l���"f&fdɕq`']������9o�,X<������Usw�}���@�=u�4�z�*�/�w}Vz��ك�
���@ݺ:w{8�q�OG=�N]�����o��������v������ɀD_{u����&�n��2&�Y81��ZD�*m���.�&"!7�^��O���a<�揖�Z���x� ��v�f| �e?��b�Vi�v�<��Z
`�ĩPP����{����[ ����|�:����;=J&S֔�+��F$.#/���j�x7���rFj��WpS�v��y�h�5��,��`�2��C�%����fi5�c{�ٺžq�oia�5N�e����j1aN�DRaf�Y�6�Q�R�9�Y�t���{��$5*��q���˓�V{ox����������|$�B�~�d������<�(�a�w�Xm��Fc��t]��o,���}�vF��'x��:�r�o����FkG8�/���� ����D�=6�vr2"��U���[�SaU�K����ݨa���-�U���oq�٫����C|��]��J>�hF�ā���"�����`��e�y����|�vrryѽn����f�[�ylh���O�p��Q[-�3E46g	�q��e��cѾy�׸�Y�M���)��^.An��̺u�N�v�ep`{�������ȶ��;�2��3���
��Q��I�c��"��ƕf���gi�X��(���C5��LҤ�K}2�M���܍��r�w��^�[���M���bq�F9�\�o�ޭ���el��=u����շnl�wBښ.������l�J�bwH���];�\&m��������c�ؖ睯k�]*6�۽�ҋ����x��p���VJh]H�\���h\8w]��1i=�w�O�'-���z]�F��v]���ի��#�8"��v��Y����x\[=Ĭ�/��3IQ���i��Gh�}��0�ĒJ'1�Wmm���+\�6���L�[m�Ur˂���T�V�ITs*e3)��2�m�q&*�\J�aR���rڈ�U��mt�F1Z�J�j�EmZ5�X�E�)X�)T�a��Z�f&%E�h�jK��mR�R�a���э����v�� ����Os�܇;����0�Vꕶ�̶E��P���[�b�X[j�J��-n��!�jcQk��4R�I��fe����Y�J�*��9����e)EJ�Z�j�:�Ʈ�KH�t�X��r��f�j"*�,V��RQ+Ŷ�`ඍCN֚Q4�˥be%�\feL̮G-U�ˍeF�r�eTDQ
��?_$����1Eoe?���I�|�$�H2M��_mTJ;:E��`�w<�@ ���mB�λD�����OX�O���1 �� 왉�U0A*�s�i }�m���C���X	��f`�V�S�����S�',���$�$�-2�u+r�D��獻/c�Q���<�ؒ#��=$����|�	�h���#���,��"�q�D����*e�$h���ń �ܦ�sW�Eu3JU#�/Lw�����������/{)� ���o� �*���T�[�j��~�i"�xq �vl$�':{����O=�ٚDCכ�� {r�̃�#�2�%E��ϝ�:��%���$�/�ߪ�C�#��ui���y���j�dbQ��f���ܝ�!
P�Y��p���,nU8\��yՑBp��5�D!�FӚʊ�fΊ{�U�9ے����,�t����I�<��f}��}J���l"�ݭ�-O:�+*H��YW� #_uՄ�^S��3\��M��JzP1���K3���gg,��n� �՚�m�z^��9���eK�� �32f
*|��뺴�!޺�D����y��{wb�ڟ�٫��L
5�;`(��(	(&*j�d���fg��ݬ�E,��gj�| /?u����v�X@����N�׀��^�ת��
�R�$���h����N����X g}��w���ms���G_zl$�$����
�����`� ��#ӛB��z:����k�}A"F�]X |�=���  �� ��y��`}���<�r������H�'s�3ؐH���].^��&�<'A�t� V{���� o��,�p�q��352�XV2ɷ�]D�Ǿ~�3�:�L�j��/^�����o2�5���f��z��=Ss�Π��C��}o}�o�?���v��ɦw\zg�F5μ��)ln�7�t��n���8㥧p��Q�>����\e��c؅HNNy�b=l':��m��;�6��E�8˸��5r�W��/\���G�6�z��16�ܼ۷c����a��qsǵ��	�Ch�&sn<�{�Òهv]O\��g&{���n��7�i1��򦑆�A�s�Ů����ֺ����wHg����qr��ۍ&d^v���1��`�urv�/������yL�v��������W���b@񯲜E��S��P�������ŀn��m��BD��f�KZo���*Z�ij��]�� Vw{3	 �_e4�_�����y�mWS���g����b��&A���f8�9�;`'��q�W��z�7�Y��� ��lC��A�Q&"I13
�
��]FӒ�.��w��`Dsܫ ����}=��1�	,$�����S�+Q%0P���ZG�6��$[}Tpi�WF}��>H������ʸ��P��퇽�2C^��NmӠ�8�X�-���J�\K�O��/B9v�^y�xk`�����~|?�=�ym*
��Q�ݖI�$]vM~Ix�޺1{;�,����f, �r�a��$��K��L9���BI�9���=��zx���C[��ǳ�7�/�p�m��ͱ=mÜK{[�f�t,�s}Ξ�#�@C�[�^�8w�w�� � #��V���� N�m֞�|�bAs,��13"b ݤoz��O}������Z�ٙ��� �A��M�y�w��D%�MTE�z�ٞ"�"��e�A��ؐ ��󸆂+��g��c7�'Y� �眆�{
��I����>�nBIW{��a�3S.�t��yM� ��]XI���ܳ5�fs�0.	e-[َ�F�ܶ/[��j�ʜW^"l�qV�0麚��%�+G"�J�fAJn	7������� 
�w��L�3�Ӿ���}l<�ܤ �I��4l:`�xʁH�=���v�f�iuD�h뽦 .����+�ۘ��D�"����]��%q��x�ه'{�Ѵ���w�ĒA)����H5L���jN��\��>vf���{o���������\��0N������r��8��iK#��%��-jctt�����Oy%㹮��I%=��1$�dF���TJ�%C`�s��ު]�-��g{��@ :�w3 F��O�8���{پtF���m�o��I@���"S^�ff 8�Ʃ�V�U~�Tq�?^;h����@�}�q&�턬�g����-�vL@ۣ��nv���c�I�^L1��s���=�ruv��}|?�w��n�O��n�0����ט-�����`TH��{�<z��&�K癉D�\)T2
SpO(��З;uDu��חq�+�s3�> پ�l�$�?Y�b��/?ӴC��oD�2;�X �㿬p����G����^� ��v�, �l�d�ŮI�L�O�"n³��كr��}u$�wg<XD -���	�v��Um�b4�j!���"o)�[ �O^eF�dX����h��'(QÑ�3d7�����poqu七у]6S��o��L/g`l�˧O�Iͽ�ēP���x��!0��?I��ϴ��\_�<�;���e��� �M�K�RXs�M�!5YU�FA��	͔S6��F�n��r����G�l7��õ���s�0��!#޶
P�!3�0�^�g� >/q�L@�v�a�7w�lߔ(��sx�� t�䴘%��H��%0mC��O��	��E�W=�� ]7�-�FG��M �c#�b�M{��>�Md��j	�)S+=6� �o��� ٗݵ�]:�sw��7�-2�{���E�*c�QR
F�:�ݑ��!���;����1A���?�@$s��.W[�3�{}�G����G-rN}TJ���f�>�$���병=��sh�Sy7� N���`|�~�f`�B�Z�	bp?0�����o|��ͳu8�Ћ��ǰi�MXo��۷/o��eU����w����Gmi��P$�ϟ�l���ƹ75ۓ����WY��[�q�\ �mu\M���q`wƮ�e
Mɍ�]�|��h�m�\��ї�c�� ��<�㧍��cy3���k��M�e��y�=rt��mk���A�$��6�ͱ��ո��ty��\tcۮ8�7Cq�wZ�:�N�ѩ����H�]k����F^`����F��÷g�ʘ�-ˌ��b�]k��GZ����N�{rk�cO=t�(�a�n^p\�^���'�Z,�-�27����9�e�'������|�sl����iX| ��ّ�ުk%Ov56(�ɸ��Xw��@%ݱ%�� �Lh�������ND54鮅�d��8��x�k�� ��vf ȕ�7l��x����vC���l��"�jncb[��_��0 Aq�i�z�?:�0F{�� ~�f,��9\�5��)�8���W�-�$�s�$�$=���`I�q=�]�5o�Y��I��u$�U�U�>� ������f`F���9�����j���Θ�}ً�vK��omi��13��0�OL�l�8���v�z�Q�Y��H۷E9��������?=C�����w�C <���@�k�]�	{/D�[�r����9}�vq0�A�
l��	`�	����p��g
$��W<г6b��vꄠg�j���ۇv��jV�v��G�޳cr�s*�2�T��OK����k۲?c�W|a���̿E�G�q���D����F��/�@��
'/'�6����t�#{V�������Lh���ŀ�[��b .^/[�,���V| ?{s?�̄���JM�&����E#�A�{�0 ���lwz��&�5=q�_FM$AMs���cb��MYxAp�<�vl?a$�ޫ��̬��t��:�I�=��3�"RWe6A�{�4���N{^���?~�ʻ��1���d띻KP�8z���g�Y �^�F.8�����?�y�v�����~�ۙ��"6�V�{��wt�/}���f����}��a@V�4��Ng�T��7aQo�M�!b먨2����n"=�V�7� ���D1r�8!�V'ư�����;%D�*����������� >A�2�aF�Q�T�屍���n��g+�p��6�D�އ�`����=B�h��
R910��"���*�V��pY{g˾S�j�_`�]�.p���q� 0�s��
;�j���5PI�u׸u��^V�Q̜H�[�U��^Ž�� _{ݑ$e��k��t�L9;�$�15�T�K����ڲ""���#'��S�ˈh��M����rM�$v�e�����˩u�\�tIL�Ʈ V�>X�n�T1��Rq's��۬g�Z�ZU��US}��A%4R �9N�b���Ղ�_{ݙ�#�]Ч��^��3=��" Zoy�����T����{=٘A�p{�Q���S��<��7lAi���_{ݙ�� +zä����V����i�W����LCe��7`��{�|�i���Aؙ����v�gt$����K�%]�ك�ڃ�TL���XH�u�I�/�u�[������o���T���N��wV�n���D^�z��G����� fC��za;�(���7;�=�nǢ�&��o
@55�0Nd�tx$�m]̈́�m�1&bɄdZ.z��$<�r������yn�e7Y�i/R�w7�4�����ʸz��}1\3*UE�,zeG���Z����"���ZM�j�#�b�:���Ȣ�O��kW�<-�f�H�������߃��n�����n�c���q����HX�ea�	w�f�HG�S��х�J13ܮ���RI$�޻�_A�z�)��6��OZ=:�WV�1��STQ3*G/��` ���@�;�o=�Z�Ӭt�����z\� N�dѰ�Rb3�*
S�Mڢ��t�q�yk�Nn��X |�GV�6�}��]*��g<� ��٘�T(&&&T6�V�����j��ԫ����mW� ���� �mY�����$�	'��IO��$�	'��IKH@��B���IO�@�$����$�hB���$�	'� IO�!$ I=�$ I,	!I���$�rB���$��BH@��B��`IO�$ I;H@���d�Md�,<u�~�Ad����v@�����|�                          ` �)@      
�(�P  �� �  �  Pg=$�����)%DH���P�%���%�"�T��T
!'�C�*�B�J
�|���v��u]�9���!��Qs�7n�]�tӧB��sǥW���z�W�pB�����ǽ��vN��Q�!m��M֧,�c�����Ooz�=�-� {���{������r�� $� >�bT*!E�/z7�}t^a�u͊t�����{���}��k��=�;�=�]*{ϥ>�l���G�[�@  g��=��o�-[>��-�z^����w�����{hS�ޔ����y��s�����:2� C�*�<�R��I)R�TJx�4t�hs���O/�c����ݝrj��{���z���=c�  �}�o�@}��Jz��U���=Wc]�]�݁w�K�R�=���e݊nڣ�� 
}鶴��R�QTJD�W��!못����<������Ew�e���z���`z�p��{�y��PA�=ѐ��h��{�C�.��` �w���͇  c�G� �� @=٠;`v�� �QA��z EERR��U� a�٠ A�t �q�<���7`��]�V�C��*��U����yP  n ��|]b_'����A�6܊�5�����p��Wmv�=��:�V6�d>      ��T�BCL��F�� i��T�JU(       ��U&5)$	�0C 0a	��d�@�?�#4`	���4d0 j~�I�R�# �4��h�1$"RL��di�Iꞧ��OS��d𧚓���?��W�_oڄ}ε��fF�����BbG�U"��!$!��1Di	 �HHB(A���e !�����������6���t!��@�$	B ��A�q BB��4�� ��B�#��3'n�BM3�~߻��鴁!F��.d����
�@��՟��*_l�܏����QB!�$~#������fg����-^N�6��
	��oc����W9�����2�|��T!TC�G�\���bj=�0��� Gd�yvsAȎn*��BѹÝRh�g]�P׵�{�+�V��t�����8��.�v�坒��܄���5q��<$p��eq�d+��X@/IaUjW��7Sh��{�w�8֑�eF<3�Z��w�����Avi&����vwg�=��Η0Q�Jۓ�F�Ha<��ϟ,z��t��ܮ"Guz�N�2�Kx�&jmM�y��u+�-h�t��CWA���ɽ��F�YgR��hLq��n�<�I��7��-��A�x��.��8+o�vv��;�$��#��W�p;��8�3�t��Bj7L�us;&)�\�ur3����!���چtP"��P��"-�;�S��[��Q����4=>}�hw"j;ó�.�`��q�G|���)(;�p�R��i�w;���v�]���s[���9�����kZ�͛mm���8
�Tc)��J`�0:�������B�&��jxL�<%��E��k|J����ש/p,�}�Ͽ,�{b�g�,,��1S7fG����S+�U���wQ����`��{�od�X�u�f��j������,=�y�}���3;��ɓ7��V��9�%��,�d8���lk�̛y���n&@'$#)�2�F��M�%��z�q(d\���ƒޫ����J��c���n��*}�9c9L�9�k�>uZ4�����s]|��N�0����c��4�kZU7�KIّ�^�Ӑ�)��"�{q��MDŦv���im0iˀg1"�c[ٸ7%,JA}Gv���U0�l$G{h�)
��WF	]ص�ǔ�i�@k��b�ʶ�+��z�4����5#m�d�Q[�b8���˰�?�f�3�u fA�A�\5a�o'ӧhW9��"��pp'�B�յ7�u����J��\�u��j�������jP���~�9٬�ZJ���N=,[Wk�ҍɒue���s�a�lb��0�ޓ�t�H�ma�&���KkX��w��u�t��"�=�@x����≷z��-�[��F�=>���b�?tL�UO�IK+xU���A0=�Y̡y��B����$or��n-��8�v%C �ۑ���*����`<z�m+�i%^�ٔ�y�r�}R�2DBN�
�T')������=s �#Un#�r �XQ|"\�jup��voK�RӨ]1���5�&�wn���IL�4Ui��O��l���#`�!Nk�4���k6�n�h��띸�҇"5���.N�{W�X�jC�fe��f���E�8!�$Щ{�I�#��3�������KHAts���,e6Ӎ-=f��Ŗw�h�7.�+���3@X�h�׸Iٸ���S��w�7��t�t'�*��'c�0�8����_gC�vO��,��%���<��/l7	�"C��&\��ź��a 6>r��V�uÍh�N���:�)�ݛ�H�%Aj���B�-�Cn
8IȜ����ҳݐɼ���v�yJ5����I�6	�˺7F� �ۢكPūS�N�sV�)��<d�3p�)l���=��a��9t��0���[���ۚg5�4�����k$X� t�
5��y��E���6��xy �7y����4ع��W�����5Ʋ	Y:����1:iG��NpÝ5�j���z�m�=hj{�nKv�NM�'Ew���d�˫�K�eI�\qQ�����E�g�w���]!��$���
�vS�y�VT{Cn�˽�!�h����QN?p���?��w��ˮv�jZ�NƩ�������!öu/Y����Q;�nV�.e4ՙݝ�w蚊�7JU�)9m���^��RÖ�{�j� �m'�1e�!oE ���e~;ۆ�c��36�;Jt�f�19������I�7v�������C���_��?%Gn�{��<9�����~�sz��!�_�]y0���q`Ň�Dw�4���Dk7y��?>�{�b�"�{p&�hJ��TFɐ氉}�7�!��-�j`�Zrݐ�'�����.�Kw'��k��(�酭�`v��/,����+�d��:��y��c��`@Ά�!�9�fW�`ݠ&Ƕ�`ɳ�n+,Ur1�y����.�5�*u�{�Q�]��N��R���Wamw��1��qO[�o����ڞt7^�Ϭ��Y�v�0=7�L�m֬����ӌճ�v�O%��l��X�b#5*�uÚ���|���c���*��כ�����x��K�Z�L�\D0���z�+T'n�=a�]�t���<��R�B�}*�z�(it������7�X:�q�e��9♩\� v����#+�ԧb�W\ոM���XnѨ��[��R;����f�hU�t�hq֚t� �u�ᘰ�;��˧M�g+��b��^:�8Au�:�w�I�z��k�p�'$�1�͗ ��ۮ��6&�ض��1���cp�� F�*��%Q�a�28dų�����B7��n�N�:2~�C=�;4@2C�
0����GZ�V�����QgZWܸv.�JtW�ݛ��XWo9Ow �2AN�d9)��W���;�>���Q[���.���ؤ��w�K;G��g�<u]-v��R�k`����oi+��L�lZ��N��/L�k���7;j�_3�.K��ݒf�]�^�b�LZ8���
Be�.躨�4m�*�'6��S�՛�[�����Q�yW��h�٪q�ʈ����unYyT��=@�e���s����N��34��Ӵ;�w5	v���78P�a��gY�I���u9ڋԱ	
���<ʓ��;8��苟nicN���m�f���b�j�An�,#��7�J7��2�y;gn��8����Lw6�h�U���6_ᴯ>���h*,�NԿ<S�`{7(�Yle�����%ObX�c
��β���T��fq�8��s`	���M���RE���'C���7��7yr'�#�0n��ؗ����@{�Y`�S���,�|��opE�˻��'�[�!��H�3I0C���$^�����۬.�('�I�s�u��*n�*��U��<�eiDA�[r��x�~�h�y�-�2��*`���
7j�=���is;��a��/[��Y���g<_��Nv��B����*��ڞ�.W������6�����廛c:M]�i��~���q�A�F׼�X���o�='��ќ�AZ�n���wp�w�n�v@��Z)ݽ�����7���]ǹ�컹&�������i��q���p�7�^���f�VKw����)��ߣ2;�^�X�޺0�%T(����%˯9�鸱�39�F	K�w����Ќ�A�2@�^�"I&1���i�Q��M�;:!�\ZXTr���,�:o5�!�:T���qѻ��&�r���=80�8�:�5 q�2���a⌖�ǆ�9U��<���^grv��'�e�QLO�*a��s�%������06��@����p,�(nǚ�#f�ӡ&m1M9ð8�d�]q�쪡��{n�;���c['>�z�!� 9q��2`o:�D4�GV��6n�����hԯ���r��c��KX:���:jÄ�ؒ�\�M��Y���+Xa�6����H$�Y���9���ł�v��OO�],Ko^�[I+��a�8���3�\x��w-���)��ͧ��FЃ1��-��;rPּ�ݔ](�m�s���o+�kv����� ���pW9lӜ�27�L:�9:�ڃBk�4(M�V5#�5��(�X�����v�
��\ݨ�׉���}Pը(3s��ۃ��Qږ�����-l]�nk��U��I�ڷ�ໄ��rr��f��{/~}�`Wv<�\�rŻ�Sa���4�L R״j5V�`�dѣ�t���8*'"������Cq*\���۱n��/�՛�+s��u^6�ݔ�ޭ��8�Zrw��䱩�?à��,�.�NNr��xx����2\�w��V��7�����;6��rٻ�
��:Z��ۇsw������* oyjS���:�܌m���&Z���nrK$�V������p×YZ����3�`�K��tށ��5�z<�E����B�7����k�uQ�:����P�����p:�O\\�2��Bп\��DRq����L;�a�H�x#����ɬ�Ʈ�yː�� � 	~����trֱ�:�u�z�"Ί{pu���_�2���4K���n���l�ފ		���ژ�~�kpw�G���B�]�,Uҥ�I\2f��ޝrn�JcIp,1:�E�0�]
MGoI��2q�?6�+�����w\�9c�O����O�Y�7�f�����gn���^��"�����v�n@�B�1�gvl1RA܀̓��ygo���j���֔&NWF�N�5�3v��4�ΐ�E�r�k���<oXo���ŷ]C���f�7��ivH�wdl���Rۑa��3���.��B�hsn5������m�EZL�,��U�ש� ��S��>�����1,͘����U;��J��C��nYOxG����F���?�QY�15K�a�|���u����)�-|����M���6hHlI��6$$�$6��BI���� `�h#�bIhHmI	�!�Ch�ĒQ�B�$��@�6	#hCb�	"1	F$�!
0&�!�Q�Cb4	F$$���А6��I� �h�BI����@ؒ`	&���؁�� l@��@hH#I� ���$"1 bI��BH�B@�6�M�lH�BI ��6�6$�@!F$"4�&В��bBG���ϡ�|w�*���g�&;��!$!�C3���!!,�@���q��E�IB?A���c/C��O�� ���k��j-yt����nMm�V�Ү��Zr8��^ף�z?z=^���ۀ����LW����2��pj�=��vx�n
c����J�8��̏z�>�n�v��y���78f��Qν�J�T������w��?��L����Ng0�>�`SӗRa^�w�A�پnz�6-䟐y/���� �>���_������ٽj�{"�H��I+�N"�n�;t62k�#�U�}�Sۙ���o�6M1��o���o�����o'�O�/oO��uǱ��e��U�"�(q�z&��.�Gw��� F�ި�����w�}OoW�a��vs�}�۞E�}ܜ��c6�����ϭ���mȯ�f���7��XKw�
qb����w�Fƍ��ېǇ�8|Γ���.�ǆ������D�Km��<��淠���ͣ��pC=�;��3pvx,z�s;���v\�G7!+�ʸ=j�S^f��{^��%ؑh����&e��x�Gk�g/p���L��Rz��L��=��tf�$�޻�;�����p�uh�\ļ���<���f]Â��dN�`MH��nkޫU;y�Pʷ��m�+! /,8H�;�!�Ù���G�k�����T�OL��F��E����zo�{��S�zr�D��[2a�4{IY����s���Þ$u=���0�^1�7C͘��3ܽ�h)L�$zN����xy'��Ү���nC��a�n�W��O'��dY��﹪�%���"#c��9��}��h�ΐ�Ͱ����J:w�_��	=�����zOw�"_a}��}����ۓA\�{�՜���`�덉�@H*��J{�y-�'ywrl��6FP�5ѣ��i$��
hv��̚Q]C/���A�Gh�9p)r�JS�77�@�w��M*����^����v���l�X�y��ؚ�qȗv��˗/"�F=/��L�W��"�'/�uY��b2{p����r��o��沇�Q/��;�<��c�o;N���ʽ�e>}��һ/�e��ygEѫ�o���n5P��ǈ��Ni����(��_vu�吇8�v����S�����IT�Ct�%zb�U�ʳ��%��Ջ�^q��1���r��^���o����=<f�W���t~�Hi�?fj��1\���"�����}UJ~��������4N�a�������4�r�*p^8�NU�a6r�N����y�{���l;��k�����Vz�G©�Bը���>�'7�k#��vL;��o���ՠ��\���׬� �3��T��y�)�;	o=���#�ޞ�:�݇�%�},����2��8�6.��8f��t�7O��1mo�����Ƭ��|��e��k{�'��#{��Y챗�V!&�Z{p�ѵg-��B}���}[a��6)���&�r�D�{��m*�׋}�oy�f��sK��)� &z{�\0�5�n�'�B˾.q���!��̦����1�ɏ[$��4z��<Ɵ��Z�R9��M-��{Oy��	^�{��(λs��o����cl���{/��'{ݙ��;(T��d����ؒ������;�sV��*��ǩn�2�k�xF2��M�}�^��z�'7;�v��,j��G���lD<�K�zLYy����5x��99��-]v�`���O!�L|�������g��x���	�JR�~�2z��
˞ػ�Y2�病�dj�7�3sپ��B���,���.��y��
�FOc�Y=A \AA��Ė��O;���2���ѝ���@�ݫ�I�h��xg��� Ӂ�7�7��#���ti�w���7%��
}��!ݏ�`�O�]Ç��g�|�&@�վ�}�,�_qVN�]U���mN/Ρw��ɽ��%�Hv�Ixlk�{�/�w�A�����6;���<�(b��ނ臲�s���=�8�1^�%E&���g~1�=�\㒻�'���R��u����<P�����q��]�-�g��G�yƦ�D1�cg�4���ɸ���~��F=�?e��h�
x��n����w��<Օ����ك��}���Sk݌���]�μdX,���:1�ݔF]M�M��J������}ԋw�Cӷ5��\@`���6p]���-�{ۅ�:�cw�x?K��{��A�������>��9@k�FC����������.��@<�蠏���|;o�4��O��12(|�p8rh������x"���;�Nɛ��z���0P(�PuDd��;��i��63n��a⏯��9{�w:<���y�q��o�h�7�-�p�U���|pk׬�o�!��Z�t
��ZG��(���/߆�������3^"����h nk���=��w�G�'	=Y�σ�/t�ac>�=zU���|��$�ە�鈬T�w�۞Z	��/����hG���^�l5��p��gd9���l��s�8q�6!��yc�aG�L�G��ny��~;�:�*�1E�YF��t_-��{����'��y�������������8d�̜��O��Fz+ݺ&�`�f��T$�yF�D��n�B-5b;��IW=^8���	�P��LҼ�՛{��u��d�e~Q�fuE;���/4f�7o\������ޕ���=tZ��ǲ��H0g^Ӂ��u�>9��ȟ�M^��:���^7�ⴌw�_E��0_��.!���x�&�cw��^s�<�wA==*�����QSr��-h����9���Do��׼�9�3�˃ߗ��s�=��]>�����bb����Mz{e���p�'7
Is�S�Ċ�D�,3m3�v����G'4}���K���g<���\�Vk$l�^�]�=a��&]��(;�W��M q�9ZUs�N�j�l7��R.��U�x���Q�3�<�8�DK�+���cH�|��O�ǰ��Vj�����=�q��.�Ҳ���w!Oi�=s�n���\ �]��r�{���o��q�;��-�Ew��8�y��[��O/�_o�4���Q^�����8ލ0�x�O�E�i�`['�O��w����]΍F=�;7�=Q�)�w@u�B��|1�Ǘ�\�����a�{x�ڈ<��$���v�����#�)������9�ö���K��r���v�p{Gu��g�zf�.-���go�9�1�?���t�p9�D?�����7�,� �!05��~����T�Z$��L����<��L�/7��f�A��䠪�h`�;D��Յ��K�x���|��ZS��ư}�Ӂ�g�N�;��x����j���E�gd�n]Kܻ��J1�9[Ȱo��5�qD%W(��w-y(�ڨ��q�^�=�zqY��o��vu{�>/�������`��d/�Wf���V�����+Y�y�#\#m޻��^P{�d��^.��=��\��s�!�x�A��<�г��p�\���g�Y������%�u��\'zy�0j��u5�7iK���S]���f�|�sEg�"��y�����/OI�'NĻ�˵"��3�w������ �׻8<<9�oAe�=��}8�pK�P�E��BkHfں�y��sw�YÇ�iL���l�<FU���Hsь{�8�]/�VoY��w-�"����P���o�?a7R�w�˻ѯ.�$՞���};5�=ާ<�V���=}�\����p!�;C-3��7�6��\���ߢw<�N�@���&akC�{�/u�D^���ϽڵШot��B6�^(�o�u����9_2(��G��^پ��w_<Y�����mŭڑf!�'�ԍ���&�8�@:�xf�����L*�e|���!���?n=��W��{<� �{Ԁ��m��J�L��W�'ow��]��|3^oN�U/U@qzzOe{vc��h�D������2 �t��v�����]Ǌ,ᯗo��G���]��h�|㥏v��ܗ����Q<��~�t[��9���:-އ��P�<��j/������;7CI��}�_^��wx]{v�-n�+u)r��'.w��iQ�MįP{�����,ʢ�j��}�,�=�4����(������%N��A>V�:�t����Ť��\M<����wݖ�2�0Ż�я_dy���S;u
��X��3�e�['�{�0�����n�}ةL��W�����*�-����p��'�;�ev�ұ�^��f����r>+�VЇ�e���6�vt�a������T�5����W���I��[��	�8w���;�X��G6������d-/_22��&;�Z��g�<}���6Wi�ͻ���콜|��R&?p�_5����-x��%Y[�/v??f��|9]�����vda��J���;��=\����>��x�V��Nw�0`���{��=�9\e�:F�j�=�{:��sw��8������V�Տ�~������}X�s���=�}�����a�ӛ '5�p��P���ҫ��œٺ{���v�f�l"4r�����:�x�c/�U�߀�z toD[�}�g�ܷN/-��|D�ͼ^��GDK�ɷ�y�n�@�t��5t�,�Jл�)~$�����/�z63��y�	G��'}0�Oc0��iu<��\܅�δ�o�)n�W���(1�!���p�y3�<E�@�9�N����[��K��(63h�k�$ �������d�'����NQ�4��ot���ҥƂ4�\�tmU�(�X�ޜ�����rӻ��qu�7���+�?���X�z����}��㤌����g�vt��{����z�������=1��+-�^ok	�q��ͮ�#�\�I��������w��wP��a�	��Z�?�|�	B1�M�D�H�vh ���@k�
T�j���*�,���#j��9��aʳ%cZ��-�v��R��nV;Rh�WH�f�6��l5�Z�*ܪmn��v�8tW��\��Y�c5%M������B�A�T��KV��0j���rѳ*S+��
8p,���mlVbR�:�FWUu���*M����h�iq����l%�rd
�!�̐��"Fi[��H�B�,�̘����K������JXqܖGWKYp�� ��+6�P���ѧ	��f����c]���T+,b�#�Z[EQ��M�j턘cwCkM���CYld�&C' �p��.X��xoXC�e��#q�e�6�
\�"l:g�k��6Cee�a��05��l��p�0�Un�R��b�;W&�60B��3e�����ڶ[��(YL���ȼ����X�s����ڛ[���J�C$9vn���8��Ĭ`�7k%R]Z�4&�T����s�،[,�0ծ4-��u��`.�54�j��=�F;K� ,�c��%���s5IY�v��U�a����Y��S�K�����0�D��v���V5T-��AQ�C թJ!�<��@e�cfٖ����ґs��d�1
�LYvl��צ���V�\K�ZS�ā�lf��;i��CT �l%�+����]��ZV[��0��A�k4f4�ch��B�&� �4�]���U&��CQ�-���uDØ�ƅ.6#�{�d�)k�u��j@���`Jͬm7a2f�l ���Ml�j�������k�	�����i�V���2��m��n�B��A�V�m	`�[k��R+�mwk\�b70ui�a�s]��`��(Z�keN,�:��-�jL���q5��Bg`�s.[lSZQ�卵P֠7 �ы�f�ek�䭔��c5����2$5��(ٹ�����K�GA�M��˒\ŋ��Pv1LCi���d+foQfy!�Sp��[0L\��:85+y��c`�	X���t�Qս���ij�*���޴̮���/)%����\]���HĮp�u��M�ꁥH+�3���1�̲�.�g9�:C7L^�7q�EBj��tn��q
��RӴnsj\K P]�36ȵ�mt���������Ս�t�A������]H�"V�mc�0Ѯ[n2��1IeVaM��b6�n�
Д��\�X4�6Hk�jn&tX����Z­^1ru��\��ZU	e�fw�smyu�	��]�ɶ�s���(�[z�7]�a`6i���x�ݶU��([��n֗����ɴA.�f�heᴅ���5�ip0Ym`!�Z[W2�t �%�J�k�[1r��ٍ�Գ�#q��h���V��d�H�m�Rd��4hyU�[�^ID�fR`]n���)�al�iYL�eV*��1f��Z��b�u�Pf��"�ښ��3DK��Ba�݌�	��"઄֐H�:$mt� ���$�%���ĎSJ6�l3�	�����ѫ26sk����a�KA,#J`ula�t���Z-4��&8Ĺ�X�V5����3�]X$p
���#͉��T��Eă�����s[(v���c^�6�v�{T+2�b�ЦВ� j83Ki�u�X)��
�C\����B-Ÿ���X,"�]��L���MhЮ�tK�e�+�,��v^����M3ec��ث��[a�#i4�V�H�M���fÄ0M��*%"�[�Ď�i,	�����+m͍D��fK�ԙc��J�LѤ!zf3,�]��K+B6��e��s�\�K�Fj�Ś��B�[�.�1+C7#�gb�T3��$t�ѭ������T�nv e����h�����f�k�i+pDm�Fe2[vR���,t�$\[��7�Ќ�E�k�,X[�@���h�"ud��9���0��!a����Ye�TK1X�	���=����],ƭ(��Ŵ�Ԑ�Mp�۳*�a�6T[�]e�����;#�̷,&n��k#b�+6�41�cL�,b�e�)-�k/^ԂZf�)�< R�L\<ʠk��m�K�h��L\cm��T���5�2�]Np��2+]V6�Ev��\���Q��J1�,I�k	q���r��2�]6��а{X&��֒��i�HY��Q#�e!)�ڮōƌ3
����aL���k�� �3��n�.%J��кږ3�ktx�b�-�ʹѫ�
@�خ]ueЭXٚ�T��-�
��ո-�D��lŲ�p�k�� �/���R����]-D�u�P�ř`�	q1�]@�T��xū2ˋ."k2L[1�4�H�P�c�F4�N�%u!l�.v�6��p��[�	]փ.��u�B1��C���:��&X.b�iEMwhu��2�ٲl@�r�t���-ŕm�̬��m%l�l\�3MƝ�;h6�W%*�t���d�6��$I�Z�\��9���t5�-�!ap�"��mR�����E��4�T�]G�2Mc �C9�q���22�]c�eK"J�M6tp��[����-)�εа��e�V�`c��9bL��%
£R�E�KK��w��u!���&ijɮba�;t�ˠ�(�2�Ÿ��Ɣ�SP^�F�Z[6bY	.�c-�j�i�@q5���i1������ųb�����*�4%ᱹl��(�eAhm)(`����.��61؋Z�Bf�W�KoPʐ�0ਸ��Sq�]#�:�de�k]���a�`kYvշC]�h	lGPJ&&���o1A#h2��Z�͖э�6�ڎ����1�CB������]�R+�=�m�f���J�� l\G(�	���[t[�uI�B��72�4��	m��H��i��5�8���9�oh��ʖ�U.�Sq���j�0�nia��5��ud�ܡ�m��Y@ta��v@���F��J���h��S��]Z2��,w]��9ҫc��L�uPl����53aa(ܹv5\�4��e�JV pI��Pδ��kJ���2�/R���J�d�6��nb�W9�Jl���UGe�h���8KnB�B�H�)��1��M`b�q�L�M��M�nQ�j

���Z�cc�\��V�<��l̬�L�q�ܵUʭV�Ѫ-;cj�k5Q%�����mn�E��J�Մ�l5�8r5�0�"�:�u�.B�E�T�p�79�:�����S�W*�UʹUr�v�ur����`�.��-�$"��W�K�3��s�+X�svUU`ZA�� ]Y\e�*���.4�tri�Gb����p!���A�F8��f�۱��.qb`�N��p�3B�.���k���k�0�-+r���\W8B�;b#1,j��Y\Gm2�:��ŷs.@�MAVS<x�n�g�a3e�K�����cNB�I�s��TD��<��H��ѵI�4��K6՘B1�Ŷ���g%m��.k�Eδ4��r� G��4F6�14É���(�KzK/�������I1���@5�&6��'� ����K��Iu�!$	N�aH�qi��	C^�� !ķ�ޤ�8 8G[b	�P�&�B8"�� t �8�Iz�Ԝ$	Ia�� �R��Nl�5� C�JZR�-7&&� �p�[L,K� 8'�I@ ��@����\-�AA@�qG��
Y�@�	(C�z�JJ^8):��Mz]i�JS�q!�HpC�� ����B[, �
H�i���6�6��ltŴ�F�[���ߟ%����R�V�h�a�5&�R͠�r쩳�af��c4���ņ못Fj�X��"�44��ԥ�ن�:��v�Y��Zj�_�z�_Q��kn�a!�t���#)�,l�Q�e��e�%�2��k-4�B.I�s�au�i�oT�R��qs*�n�;f�X[�fa⸲�<Ř��5ev��.r$Ç��/d�K6��@m�)�ΐYW<��#v��1�Qr`��؁�qAP2jͭ$f6�vv� %�:噓(��[FY�6`�5��A��&��хf�$�kk��jm1�+kmH�Fw]�h����/���ڃ��J:�L	�Fa�D���+]������i-�[�nE�o=�Ҭh�̰Y����e��R]�S�[xDxK	�.�^��u�B+b�\�Z6:.
[�/Rճ�T8֖�jc2�ѹ#��)F�K��s�`:#����h^�m��&p�a,�A]-���V�����)�;&Ľ���pc�f&�\���30.�k�J�H�6ȬŔ.k(�z���H�[�=#��efD��ZT�a�P����v�K�Q��q�4Me�j;Zm`dKi����ڛ6$n�,vf̹�̬,�B��.�i-X�WZW2���T+Yj��B����nU�[K�M��J죰�{QB�eT��i|-����%�C-,��R[�����2Y��KP-U��B[i)�ѱiT,U�V�m!)-(����ť�h��-�j�`� UVPaVD�aF�� ���2)���YH�`�F��@#��"0�kE��k^D��JD`�%�D��*ؐbH"�����?O�	D�&��gf�O� H$�[Tx؟����kۉ'Gh�3��O��V�$t�1�����D��u�	iUM�[���H�*�d����P$�mQ'�4�4�u��9۪#��38��"���.3������H=�ʈ!���~S5V����@_�7@R��A%��&��w�q$�C������E���ɯ���hV\%@�\��d5r飩���ȃ��W�� ��Bfe/�{c�i��$����v���p,K�����䔡&��ͪ�<_�2�3G���O�s�tN���x���3��������!�'o��=���h�π��Js�c~����oj�N{�z�קN�
񺥑��J����I�yU��jjB�I�m
'w{w�[�\�#����{Ց��.�s-�{��(���{��|��@S8$�"���^�	 �q%EVk���/��i{Z�A�ݸzU*$��� f\�lav�nsƅ���
�R���f&q�՚��[۪$��$�T)mc��=��H1w�D�y���� �N864�˛X	$w;�$�$��o��3�R�P���5Q$^@�M�y'y93x{S�jF.G�g�V�۾�^���ݺ��E�z\}��V�r��7�^�չK_�|�
#�I;��3j�K�{���>��h8}6��ߚ�[�K&b���HM�W��*�ɘ1)M�*�9��_^^(]�{v!� Hu��R���s��J))����}����5��U���6�;l��zO(�Z]w�V���ͫ=ϣJ�v�?=���ؒS5b���D���q��ڀ��UDM�I �[��C�[a��5}~'�ڐg<���C�a#�S�'�P6&�����.-�d�q$�w�׫6���T�HMYn�0m佪8lp#6$�HڷT;���.� n�ܢW���oM3g�x�'���E���g�#���-�{ں�r�s}�F�]�K�j�c�};�,��S����]G1�WP���.�A$��P�w�*=;{'���a�Jk�4	�Sc�T0��WGF�Vm�mQU_��#0bR�eTO�!ݵDsx��O�;����q�Oy�/� ��W�}Һb���w��ۥ�]�(ð��w�ycuAW����=�e؃�~b���� �;_�˾}ڈ}�)$�^-��ۚ񗪉&��
7D�ښِC�J�,Dv���݂��́x�Yy���eQ$��UH�a�H�3���yY�����~��i:��jBw��}PK�ot��^V,Q�6j�h�S6W-%��6��bm���W@.6��4�U-]�	�Ki�6�]3�j��1������s��U�-i�X�v�۰��d�%�i��Ճ1����l	�A�t6�kLJ�͆�f鶺�i�4�hh��)U\�p¹�0�K5X皙��l4v��4���
JIJZ�����0)`��TH��
$�Cp6�#5����:��x�9�P'��=Dc�S1n =ن�D�-Z���D��O�1�5�b��A��3�@1"���>>�O�+�.9ȵ�
��>۪>n$��.��L$J��9+C�ξ[���Ȓ/��_	� �(Q!�ڣ��A��3)Qn$��bY+�GWv��Ǵ(,�$o[�/U�T��u���I ̰r��
l\�Mu��6�n��:�U|��o�0�}𾽡Dp�	'���*mh�ηPqJ�]�-} {�}dQ�u߳���E��on�uIH�4cjk��b
���K��"p�qg�R��<+ޞo'r
/�bR�P����$�vРn��˨m��l4L����G���$L�X"�dDKs�C:D�Inڮ��T��j�/{��^�f9�d�!˽j�>|���b�h�8�&�鸘���W`��B���\Z����5���Ȁ]�v�{r����u5���JR���Xq��-Fl�,�QRJ%;ΐa�	�����$��w����&�gA���]��n�&JBn�;ڠ5��x/gA����ۺ� �[�Ր�-{ЦE�R���؀�wB�"�+v�!`��D�4z"�����WM=�#��h�B�v.Kk���7�Qzx�إ�2�"Hd�|�������0�2"R�Eǻ���	/j���r�z�~���Z�m^]���T��j�ox�,�닪����$>}TI��B��ȥ�s:�@�	�2T�*bAA;��-���*R[3���Q*���DĠV0V�UH-� �ɐ�EeD���hQ#q�P$^MȈ�n$�����@��������Z���>'3n�]�'�]��%W�(���cH��Xn�E r��F�q�%Q�0��T	$t2'4wI�2&�!�[�����{d�]�Dv0�$��w�����{k����=~��AH��}Vl�vo_�Sqb�u,�����'M`&��F����*���x��D��T�V�nm��z�p6��`��9�f��f�/|s����Ln��)�=�-���+o4��i�YU�פڦ�ZK�jÆ�' -�t1K��L���]uP$r�V�Z��1(V
���!R�E��u�y�>���c2�W]Fk�6�̛��Bfe*�d>̪hj�i�� ��̐A�n�p����������j�'�t�$��U�I��M�8��A1D����(�:�n��|;����S���v@@o{�����ߵ�c���I�$�J�5J�[�������-)��W�p��;V ^4N��n���x���֡��ň���
�lI���öbx��5MF(T�:P�+٭v��`��Y�W8e�s�tش��e-�!v�4�U,K2;:Z��5�"�A1L拍��]�֣ظ#)-si�G1���չL���˙Y��9.U��WFݵu]`WF��c����h���2L�JRW�p��JSTQ��J�j��{j<�v��2����}W͞���i���^����پ�4��_���|�パ���j��bd�J]�{�P-�Uz�l3da ו^#��Q7�r"3�L̥N����p�}u@�y�Uz���w��������bIVw�@�8dOv�5�׷vւI�H}>���ݩ$�ڪ�)T��bgLۮck8�%B:��T���.L���H��tA>7���=�]W��'�kP�[�'�<bB)M����^��ȑ+	Rc4��ػ�܏cù���I�=�0L^/ח{;Zf�=��^��TI.�6�\R�*��M��Ji���K�݀x�D���]j�����Vx�#o/#��R*Ļa4��,�@�ۯQ��2O�޷=��<�]W�a��"o���/_��bZTc�$�����d�5۪�J%x��G_�[�BH�IE:� D�TɆ,
nK3��ל(퍽=%��`���޽�Qa�$�O���1z�ݞ��>q�A n��jLH��Mﲽ^Qe�R��	.�I��3���VZ�v��tHPe%]QFI$������	>���v�D��#��X�¦U��R7}��2��7�rJ����|7�v�|�h�e������kQ7�\Ȗ�#��}�u���~��=�(n���o@����[0?/Is�84�x���1���2�
7�s¬�����6�j�g�x��W;:�m���S��b����"�o&7���x�ǄO�W��I=�5�������=�/^�Y��W�i:�N�����|��IGT����z�}����7�i�X��X�041)M)KE�� 4r��0LD]ۋ����������3�ѱw������ދ�1�u^V4I���e�ϧj����R{��z��V��->�8���g�H�����g8=����9� �8�WI��`\9.���w	��w�VQ�#�q���k�l�M�a�=��G��Y�2�'<�Nv�,�mY<r����h����_l�.쫦Kԫ�L�������~����ܻ�_�'��Ѭ��oe��d���|��]��b�&���3�яc�x���_;��5��Q���bU}����g��8��?����6i�:ά�b�m��>��
O�mj	|�&61��A�!%��@	Ŵ�e:�
X��:C�B� 'JRH�H�@�8%&:Q�bjH��c#	L����[%�@Z�a q �޼��А!��,8![,ŝ C�������@ �8 pB'�����%-��!	 Md�-��q �N�ȅ�X�h�J	3�B]i�������+e�i17��!	)ԓ^�� ��� @�[N� t�)��� HV� ��!ou�w D�H�:kF�wbIN�;Mw0�S�v%1I^ׯ� �X;���P��ҍ��)�r+b�yz�o���A�?3���dS!Cq5d���@�g�>"�$���}~b��Yc}�|G���s3(�+�uD���u��Z�	Q&A$�{�Q-����LE����<���f��h,����&�W3v�KRj�m\�_�o���'$��ϟ�������ܻ�[�x�jW��	�%�ڣznBH��sk�������]f�D�[��O:���Z��5�I��N����wB�$����vO��3����
-�B�)+�QFu^]mE��MX$���Q�$)&y�����mΝ$����b[����_@���,x�sϹ���swB�[+)6d���Y�~*��.�����_m
!ΩrQ���ٞ��|~?�ל9'F*�����@�	Ͼ�.�^d���}�8I�%NRl��k�Rm��mrvJ�n�I)K������@�2�6��=�D�q&�e�ov���u@�ɋ1�"fT�n'�e<�P���R��@���Q�I�_�gk�]l��i,�c#���j�;�@�2�OE�R���4�Ax�	-ĝ�w�� )S@��C��U��V;� �;�A$���f�Ur�羽mw.�I��n*d�����ۿ�᳂�[ʯQ�I��_!]��c��낮�U��H�ddwW�}1G���������~����R�%��X���,�L�#�C��d%�TP6�W+�7u������D3�Mf]���u���[s(�D6��61C;�t�3<gY*l���K,\Te��Z��(0�6��y�C3i�"�6L���6�I���a*��Y�uc�U+���̹��[�ٗ.TJ����:ʑC-��W,�m���0c�2�U�����7�Kt��׿�� G8�A>$7n�s!���1;�T	����ח�����V�o�#����};��X ���}�J�&c2��7�������K7\	���*�\�[��ؐH'��[�*�dn0Q�MYo6�Z�X���\q���� _;C:�+I.�K�oJ�!P6��x�o�c��D��mW��T�{���MÚ�2�@H2��B���MQ�934���U�����>�pPe%��IN��6�ȼ��c��lp8��]����B��j�{�UYP_�a���+~Rk� W���5:���.���������,�E��sE�3G#�tF������|��G?���Kǯ���"�%n'᾽�[ۡ^��lon>ފ�U��y�B�,?i	G��%G��~z� wuТA����;w9��b��{pdn$�(���mQ�3"I���j����˰u�|�̫�;��S�*�D��7Z���QƆ��@�Pj��UUJ��;��q:%5��j�#x�Q�q ��Wsb�w����P3/���UUx���.�;��2��)�o��D��PQ��s�"nT�(�ʢ}�$NJ�YsE5�n�M��q���供E,��}5o�w-˗d]�'��ʏ����K���������t>$w��A/����"dĠfĻt�Q�w�x[Z��A�9��szz�� �߮�.�5��)�6����z��c����<z0]�n�l�I�o�y���"vXr�X���RGZ��Gl�s
��ћ9��.ua$�vw ��O2�6�p�I$��uEVy�;AZ��<x�'�A�4�H�eE}��)����r�p��N ��|�w�i���[/��o�H���*(�$���	~�s'SZIg�����V/M��Ji���^�}�b�$�̂I'��Ux�n��4����������!��r缞wx�zx�0�����,݃�R��w��Ԉ\&�l�~��q^��������!��T��{Ҕ;öH�� �n�_;TV�'�1��V� �l����ͩh��]	`J����?|�g�y�&bG>�}B�$�����UVF�0�ᷞ�3˿N�"���=��Ո�ߐ)�q�~$]��$��u@�V�z�,D$.$bD#*8�����
 ���GhU�Y	*�P �6�����ffa��m;.���]P$�ۻ@�4���.��{�]�6�ʔD✄�=@���%@M:[v�3&Q�;FGs}�R���9��H���x ��Ҹ��C�E�u��/޾z��*'�Y?/�/�Bkc�(D�#�M	ae�33v��ɖ���$�SJ�Ue��`�l.��f�L��.!�����H�1#"5�hB�F�^��,�ks����J�J��"Fl-6��������6��,60\�i���ڋ�v�fh�騡�ٕ\�J��ѤpT�i�ݠʢp�3��v�h�\5��V��>���cf��nu
$���,��Q�{���:ɻ���{.��k��oM:!�A�9=�I$v��@�t3$����TLv�[L_s�d2�݂�j�AÄO�'.�c��u3�V�'9�Qt3 ��1�J"AFTQwّ�7n�]�����D�FF�$���OF����g����38���J�Dh!;uR���Fؑ*�݈KH�}��s��;�@��6G��+]��X��*1�M+lKe)JIJYo�4��$35�B�,�O�v���u��xs��D�a]�% ��R����Y�z����_#�.�c� Q5���1�x��"��Ex�u`�6Y���ol�Q�۟ĸdI���p$D�K-6�h�؋��
1x� ��Q&1��6�]�'2	!�j��l�L�6<CFoWXlɒ��*��u8�g��9F͑Y���AE(���P$�۪��F�U�\d����M������Р���ë��i�;[f]WP�1�BR�k�]����l�W�߿����V�m�
��v��ܫ3ʔK\  -��"D�]�QF��u�%�4B���!�@��ff������O���DL��ݕ����
 �!�G������"�+r��V !|'V�5g����3����nBX]��6xɪ(R7�����'���B�??�
��&b)�8+D�m���5P���T.�W�"6t�[ڠ(�{�g�Tʃw��5
8p��/���2O��U{:��3>9S�ż��:A�ث�]G8��6g��4�3n���Jc5U~|�/���[>z���z��Q� �d"m��*�rׯ3n��n�J	%H�~$�zD��f�ڲA"ۺOC>�B�T4���ZJIqN:�k��ƐWw�kN�J��,{u�Y�ݨ��2���S�JeV����6� ��m\u^�\Y��p�c�R#�{�����ڙ{1�Li&�KTM#8IȮ5ե�[u}�G�v���13쪓Gg����1��g:���{uD�\q�A��_uݽ���i�$�B_z��EJ�]�p���Ĭ��3f�+s�����M�OS��}����  ��͵�vP��:�����̂}���Q ��P�e
��R�H>p̐Kv�8�S��N{A����EU^,vD W�o�L/4�|wwVMq>%ƙ$x����s"�RLH��]�\nM��$�'�	��T	/���o�i�%|nx�5�T3$�U�j"&L�b짎�{�EUl
��͙$uΨ���|*�WIh�?��b�1;�L}�V�'�[U���<�a���[�q^���~O����܉��z���Uo���t��ݣf�[�poX�wé�g�A;�_s|�h��
�`oG�@�<W���A�.��a/���b�Z�4��V���Y��x��ڷF�;}�����ۺ[�ɢZえ�L�c��D�Jγ	4T=��W��:wF)�]�3�oql�ڄ�.�ȥ����C�����
6\�[���m<'#�,�o{gk��j��3�3�M��gr�YG<}��Ř�����h]���/=p�w{��O�'���J���ϯ�k^P��đ�� QNn���PGOzCu]V��ë�#���<0*�#�tEl�IԶlla�H�X���@��o��I��	��৿>�p���aY�7�,>�}4#.�Ӷ�>��0Ցڸ{���/xw���"y���ν�:�O!���0j�3N#y�w4��f6<p{��2��R���e��o!����j�7r�aٶ��������ݎdۅY�L�JsU/��ǴCu�E�i����	>�&��S�"� v�Hpu%��I%��&:b4�ԓ�;�)�)I1I��c��8� r�p�֒S�& JBp$��&$C�pKl�f�tNu�ى�3eK��Zp�/$JS���S�8'@����ӂuS�,!Ԇ�H�pJLt��8&:À�t �I�݀�	�):@��c��1�%$�D�N���8X^��[:Ѕ)���Y:gZ��\=YA����Jc�b��u8�x�SEI��iK��1�I
b�F&5� ���ʮ�,�˲����s�h��5
�6	i`왭ٚaF���^т�4��*���IKtz���&Eu�@���SjX�2�YXڡ�:lj�c Za�[p[6���®�X���-�������<����%1t�UM�(�8z�Bq�
MN��K���Z�2�DJ�+�Eɨ�jޡqd��3�	��ZX!+5s��l&���բ����٨hW'�M��K�cK�3�Vl!LZ�j.��B����<�Rʺh�*[��;:�ˤ��(�mٮ� �%�:�׶��M6e]v�<�Kf+f����q`�P[j&2�\���e��kZP&eR�	���\*�l\�ԣM��u˦����l1vv�c�������t�L��3Z����!]u���k
��$Д[u���	�I5]A��-�kj2�� `5��hafqt�u���M��P��Z�i���RR�,�Q���T�n&�m�LncV[�k��H�1�V��2��j4Gd�4Ҭ�֕�K�������FܑKn6Q��4.ȕZ�[Y�(�l-�8���R Jb�pd؄h�kb�X�{:`e�,^��]�4�бN��k��5��a��Y�����@@��Y2�MH1��F8�f�`�Z	��;"u��r��J�V�GG39�eP6[r��։���V�`�M\�6�Qm*���Ʋ�@2e�&�H2��iv�F6���i\F��(�SM)YeW�����ŀ;ip�� �)5�Z�]0����mb�+P@ҳU��-�t��Q!q+�jP�X �k�Q��RjM�V� L0���J�s�]�i��)V�d]��S!����F��.�6�0ћgMF3[T�Ĺ]O̵��3z�m��2�h4{D��2 u�]j��;{�o���	tP��8�$�}U�D��TC����� }�m�/�+�sJZC���x��9|�!� �*�%�j�D�Q��t�9�FM�����@"�ڢL�s�lI��T	mڢci�S1("����Yy���(�uv�'�{�P$�����nD�/P���H�*`ĉ�'�(��93�u��a�u^$���Q �d]����6���.�lbm���m@��R%�q�r�����۱��o�6 ��c��;� �h�e#s�J�ﲕ�]�;E)��)�rv��<�}d�l]�ӎe�V?2���oP�_#�0gtE�6I9^d䬾]b�߾bW���6�=�a���jf�k��ꌬ�UiУ�4N"���췻v ���R�}3���~�w-Z8���:QQ(�J(��m�OM�H�	 �ğs�C،z 2��X�LĤBJ�(�|H)۪�������p �wj�v�f8����!L�ec�2�hX%� nڦX�\���y~�Z]4���'�.�I'�����$��HH.�A=�spff%e<j�݄�M��aI;�$������T��p�T����Exq$O�Q"=ⷶ�v.�tQ����=��y:����>5>)���~R����s3�<�*���D�m�����Yy�k�t��g{o�yӯ�$��$w�*��'BbeA���hݍ�Ө��	:�hQ-�^�ʇ�7e�`'��w����:6�#�ګY������#v��:�N�Kǅ�w���u'�w���5QNi�&.n�mȸ�U�����<[�b+��2� +so� �}�T�hVS���E(�%��Q�1eJPbdP-\�x�5�����ou�Sm"|z1y:�$Sۛ�31(�)�$[h M�r�HN(���+7vPr�eK��d�ٺ�>+-B�x�	�W���qכ���^�*r�"�&v��-�ltI����ɫlN��Q{+��l{����'g�����ٗ�1��7�Ƣ��ʃB��Q>��1��B{4�[ܪ�H	-ă����3b�?֊�=H����i����M�K�ʹ|��_��ՠ�î�Q6Q$7
���N����'�$	ݶ҉�^I+�U����"�M�'��iI�A���p��o['�S��SS��0�� wW���{a�p���A[�<������~*�Mܡ��{)"Ip$�m�EU�{b�j��� �zT��H��>w��z�K����T�B��p$[n�Vr��;j�X��ێ����B�~�:�������|�|��3����υ]����wSv U<�j��Ӫ�i�\5�J؛kK����
۠�[Qáe���
(�5ZL�%p��[kcΔ)m6B�l��^q�ې�\�*�H"���-�V�f��T�-&�vZ6V͚��0E+b���꺘Z��Z�&��6Y��kj�\���U�,�hl�UH&�iK�V��,fڹ�\�Z��>�}�$Q�L���G3@���ڴS��:�.`֢��7��T���FPr& ҩ���$7$=m
7f^=�/��������W`�@�6�K5�zW)�SZ	$�Ē|�
1��EUSQZ6���{��Wh��[ʠ	%�����sZ���"q��Q�&A��c �=�~ϸ��n����^�����mR>�W�E\�kN8�A��v�p^R�R�ì�#m*���[��REL���=�p�s֬H	�C��G&Sk�x.�>��W�شb�Je����kQ��P��9w��X����8-����8���k����z<��i����FK���c�s?x{��[A:۪�|���1O4�-���:�)D�����^y�������,qD��z�
=�P�_4�bPE%v��}Ҩ���S�|us�@��Ƒ$�k���X���M�%UBB+F�U"n$����e���V�M�H���Y��7�_���R�.� �d��tM��+	��q�p�wǯ�����o�W����m*n�����~�rۻ��}T��wREL��G��3��R���`�ڡ��{��N^VX��ӌb2&&T�t�.�H ��>n�/&F���ثFu���2M�4�~�Y��sW��T�g��^ً���Y�I�Y��r�m��Ҟ���)�(��N�a˦��b�t�A��$���7]9O�rēv�&��3�	+�X$�n�HN���Ӳ7(�N��w�vE�J����R�|IᏃ�nVź$r���jh�,ȈRJR�|YI)����]$!�I �n��nө+��� �~ɌrGI�·�V�~󩾃��^��A�~ݺ����������N���3!A���_� ��Å�^�����3\@/}��Ï
�*ٶ��Do�7ˁ$dĂI$[ݡG��#k�S:p��d���z9��:�wg��|�Kw�ϓ�H�닽��K]�ښ*�\ƈ_{���>������Q*Q&&(�_ez� �f�f�s�*}�k5�x�i��MAYH��|����9�2���Ml^lYAhM7`�\���<�SU���`]�T�m��w3|m��T���;M�:�4�Ow~�1�ӥUS�H�.�1��+���6�|o}�]��D7	xD@�HI��Eĝ�;�V��}`9#�ڰ���1��g��6��3ϟ���+� Y~r���w	yK�$T���{�f�/�����7u���6�gu�m��{�]��{����u�ұ����� �����O�\��k���o|�`�~�	�ma��=4�Ͼ���r��<�0����goz�]�bڷ��su�2�|_������/��C��;֣��r�*:���ۛ��L��:9�����.8/=Rh0lRh&��jVmX 6ʓ�5a�&�r�A��p8�n(UeR�E�Թқ'&ț��؁�̶�0��\�4��1eP��te���fU��iY�e��f��U��)��]ak��5�U�B��j�[\�qtG �UW���� ��O��2C��E㹤�$�}��'/�����/��ΒI|V�$��?n�Z�n�6f�O�߇H_��� ~: ����Fdud=ؗ۾��8*f&Fcw�����0i�o��}w{y�����m�ߵ�7���C�:M�	���RD�S�$��n%z ��t��^ϸRI�wp���If����� �n��癮��G-�6�m7����i���,s2����?���8j���ŋ%�6��q	�,�MM{a	UNWp��rS.����
�`f:����7	^��M�)�$�$�CzP̭Z *)�����'���ω6?��R�Ϸ(�#��O;J�Y���>$�w�}N�[�5[���#�����f�Y�Iw�<��#rgr�$�I7�{93 �X���W�>�N_�>�:�,��!2��K�}$$�'s�g޾��{�����m�]r��m��nf6�Z�UQ�2L�\>��;��N9��I$����BI$�����z��w�N�Cm�&�;�����!$��/�,]�$}�*""�u`\��n�;Nu��
��Sנ�\�W�hZ.�,�r�KŔ�����>}���F�_[�ߟa�$��p�����wd�E� ���F%μ�%���G	��&��S�6�y������S{�-_}�O��&{�?2�f�* =���BI�F�,��{>F��xoVkx&I���(��U{��b{ހ�4j9� �(�U�Lߞ�(_m�u��fO��՛'��\���t�L���;|R����n rng�<����3�����>�}�7z�}�3�Oz^�p=�W�����m�F�\�O�\���=�\Ӭ�N� ����l�Q"�
m
�����q�ᇰ�Ŝ��Fj��T�u�G�����pï)����7�������/Z�e����Kw۵�Tw���I���7��׎<`�i�����װ��Ũ�;��wf.(~^F���y�}��	8����n�}�fK�ߖ���{Y=��b3��=^��;�z��{�@}��Y�p����w�~]8�����m�D���K8-ѧ���o���m��*7�-ejB���T��<R�9=�������Es�T���ؚЇZ?_$��R_Ĉ;x��yG���M����{(<�뢘������0\�Rֳ޾��_1ޞ�Үx&/{�����o�ѕ�璉����#�L��)�\OB�Jޏ>>g��4v��O:�y\�����]���ꨴ� 9�& ��6KdP8�	8�P@���H��� $!�)ؤ$8;�HF��〒'LM�l�R�L,�	��pw@������!J7��1)'$��/[ҝ�&1:����u�����e ޜ��ڄ�;�LN�$Ie�� Im,�H�F1��	d:��#�9$�BKia��@�IzM
v8%'u%� @�J@�Im��N�R�&1F���$���F�3���G�����x?��u,��&!�o8�ړ/�u�'	_I 8I�o��'	�z���{��$�g�B;x�;�t��\;�I$�>��̧Yg�}d�H��$����>�H=��UEH�Cqӡj5�H\��؅���ݟ�`H��N_���́0���8I��n�v�����.����>��"�NjK4��S	��@O�<�k쐖�i�]Rm����1�������ݝ^�j&�]�7��*m��fc�S Y�q���~�q�o�tOf��t���5�O�^v7�1��@�sH���B ��۸;u��151Enk���{��&�b�#���/<�zq�{fI���F��f�����D|=�{���m��o�u��#�UK���g��$���x?D8�����+I �7������Ih���� �wB�JZ`Ǜ�а�m�h�8���X�)$�$�6Re#"؈��* ��PL��vJa��(Qgu�l$"	�OqCr�� (��NHL}2@<�?�;�S�i=�T�M���nf06��Wz�x�X�\ʍRrL��ߜ�{��� 8N�i�9��W���X���(�I���Bn^��,%-"8O��/?gf�=��$��� N>��	8}�؂�D�I?|P�x��9�
�~'�O��;�L�0�s+3m�����b��DCp�A�(���Sc1�b�Ѵ��c\$�o�]������ӏ"��r7*3��)�5W��^��Q�4��I;���_k���ƌ�fJ[Z`4�U�3j��vS=mu����%�wk�Wb��\V� �渥#�;�б�a3��!Թ)�TU�X��7K�e�6����\��혴��i2��H��6p�������Y���;BV2�T*��WTZbP#�sRSa�^��*��t���uZ�_���.�ge���m���Xf�f>6�7\
w���[ڴ�ۮS0O���VӋ�1)���,�dq�v��ogo�'č�t(��H>ښ�o&ݙT9)6�[�K��P�;t��'����۾u�[�.�T���n�TL��UcB��%�j�(��-��'�/�Й*
�a��B镳��mr����ڤo��~gy��A�)���첛��G��ZM�K3�R��cOJ�����ݚ�yH�r7�:�]�u�T	$�����2���H�c2�����,�Ίy5��o<װ�cӏ�8w��8���:�%��{^�[�S\<���OҲ���������Ϋ��D��$�K������m��/�T�aM��=>)���rIif�CȒAܦUL��-��Z�7�I#i��or�s4��xاVz�Tj��fp�}Tp8{{��H�)���aIn�^{�z�'xK��H���JKc���uv3/m���:�V��������n�F�Iws�Ψ�ft�,�,�$��e�0Υvy��	P!Yva��<pA{�|�&�͈������Xb7�I	Q����7|�Q"7я�:j����WoC�Bf��P��[L`ހ�G�k�wÈ�z_��8�{A����5�?o:�}ｌ����ww%��E����
�'fב�u�'��3e�pM�v�#cR��Fe�F��Z4U���V��v��o�Є�莗�;f/s²��չ�	������f�;u���U��<��Х"I�+ޔ���݀�A��;��;�)�o�Uvs0faIL��/�s��r>���D���ݏ��ܓu���8�P169�-"�>��7"W;^�x�$t3 �͂��)I	P�*p@�cP�IpȒ9��=OL��̻�7f��G�w/�)����#Ӕ���ܺ��{��C㻍Q��|�:v��s<�4��D<�7��M���2�ID)�h���C(s��y�`�׵D�X��7�Tj�|�mg�4'O���#]�SI����͆���&AH(JRQ*�v��Fe��,��-ݪG���/�[�۰@}�u6���݂��H��Qk��h����� M��{���u��AL�RUq$�K�@"GO[������H$�nW��ө@@��n𓱘s�&	��=��@������n�#�����R���U�@ݿ���no��r�c�]�x�Ψ$��ܚ�(�?iT;���w�]�Mʷ��r�M���Ʉ;6`���QS�6�s�����I:�B�}<�eP�Gkj�n�R�Q�3Z��*��f1�#�����2�B�4ё�]~��jK���k�40[Q1A`Z�	T-�W$k��`CV�툅lNѳ@xl�l�2�mm%�홖�)u �&r��2�, ک*��A�d�e�����]]]����6@r�XRTÖ�L͆k2�s�4K-�U���>���r�����>}��>��}�1��Lw��[H�iTD#2�@�K��vC�����lB ��fjD�Р
��m���ɍ'�/*nH��؝s���$�^�B���eƒB�Kۭ�Wg0�SeL���d����
$�����	����c�%_������q0�h�iR����q�������p�۔��*
�C����z�]kY��f�)JK����
RBTT��|��̠}&��2*��)�U�����`w���F��uL�r`u�ھ/�ބ�5�["?Fy��:?�?��ˉ=.����:k8�>?j��N�O�z}A��B�HB11��7�v�6��Oy���b|�>���XۢJM��u��U�=����@��jR�\y�H�]����qZ�Bx�fUC�C��;k�h%�U
�#(J�3*fq�4�#�����C=���zN�����>���z|qc�vi@�8�ɱk�n��2̀uE�U�ߐ��T��j7{��@�� #��\�Rn�BI�Ԁ8o���'SS�UIӲ�%"�s�+2���A&�zK�!�MX��u�$^
�Q���W>=M ��C%:y�� 6�ݮ��w�ѽ�]�Q�:��;}�:�i[���[y�T�]�3��I$���;����a�q�3�&���jce�.�����B���yޮ�A�u�_.��n���������$}Yav	 �����Hm� ˻*�b�H1�-��n�uH�*l�5-./VF���nV���/ϳ;;V{�|�m�D��u@���=K8�|Fe�}׀�8�PLM�o5W�&��	�3� i ��@�5�>갓��D&�JR�(�lj�B�Mo@�Ƕ��,�v$'5��s�S(�JaMY��O��s���^j	�n�O��]�+Q8�E[����?Q���1�
�~D��q۹]mGa�Q|*c�z��*�g�x ��>)�\'��B�H�z�(��C�$����V�ZI-� ��Gj���7�;��3z^�Վ�D���,�;:[hX6Z�m\�_ϧ��r������"	�-�����vu�76� ��u@�]l,2�JJbUx� ��*w�WeW��n�HGo:n=U�:(j�/%�4�)A169�mE�z|a��be�^7U��p'3D&�JR�(����}�暾�+�tI$��>|���n�U.7��wuN
��[.'HQ@3�}u�=� �CnhNyM(��U�&�ˊN��þ�?��kr�k��!2ۦ��z�n�r�>�c������sotˈ�܇0�����S<�9_j�W�{m{�j�y�#�V��/E���L��[�w�c��wcagf;�������|��r�ņ�ʖ[����/ɂ���Tq�3���_�ʯs���(�,Mx�K�+�G����D+�-��mL�|�<)KUR�8N�x� ���eæη�Υ0%����=tҺ=^E�dU��J`�[��Ị�_��9����ΛX�_U�@Vt��ߊ���u�.��Eoy�Dl~��6w���Ɯ�Ú�.����~��g\���fyD�Þ8�v����Owެo{��9٠�Q��Z�^SGj+n�ޣ�j�8�9)ʊ�g��	_�E��w�����&1LJ�;��,�㐄(��Y��iH[)%EÚk�������{��M;壷�_
�^Q�U����L��������A�q�~�i�;f�$�^���%�8��L�ξ�:&{�O`Cоˍ�I�c2�G?9X�s�M���`�_Q!�ט�J0����UA����"�!*F�&JL�:�Ru1ؐ)$��M��pB�n�Q11��� �i�JeDF�	PQ�����9$�"pu0���RIu�:�1�*b��)�����b$��^�$	���Ρҝ1�����I�Ĥ�111�)$N�t�a9;II�v8:I�d�b��)1� ĝ�&����b������@�BR@��md��@�qe��-�JI�� R����ɢwS��@�� n I����a��s6�m����̘1	��L.�4!-x���m(��3]1��%���r����PT���7d�Թ�kk77��:�e�!Z�P֜�fIa�x�e��.�R삜�WU����v�W����u�]a-�`�X���cuVͲZ���mI���E�1@U����zòֺ��F��m�����gg�W��2ؕ1U�h�fc�f��}knq��ͅjrlnк�H[Fl6�ݗ8	F�F��,x��W��2&�&M[	��P�-K���B��P�YU�M���e�%�4�u[jbZ[T�/���L�T��ModJղ,D��jgU�L�X�57ҥ�dc�p�T&%����[���������h]��ĩ�NHAى�	����4"MH�KH;8��FK�Y���k-��ܚ��M!�fD�U� @HĊ��bPa���vq[�Mwf��l�����6mH�6���J:�9Jq63h�K�esc6��+�!�� �b��]WF1�D��lE�6%�֚���st��gKp�H:�j-ŨVٓXYM��k\f+�C�2�P����x�&���|������	p��Rk3�ݖ^1����j����3I��T����1��6U�:3qQ��ʰf`��V2��+�]V9q`���nUUF9�l�W�G(��[�aa��:F�i��ɳW%֌&\��j�t�nDq�W�$��^�H�m�.6�T��!��6�[�k�B7�uה�&f�d��%Ɇ*���b5ҋ�{Vj)sin�s*8{s���p,�����ʚ[t�fr�Xl2�h�h@�<ѩ��3��U���v���p��h�e�%VYY��6L3c�w	�\-���¡LV��k��V�iS�R�.�U��~�/��k]T�1��힉�ȒA'��:Y�S�-��7�$�QꈴB�3699�J��o�	n$�y��늾I�+���Tʄ�%P=�$N����JcK{��"H �if`1�J	��-漎�Q�W\H$�V4/�X�<䳁� ��h̥(�Nׂ$]�W���R�9��!LH$�V9��TeEJܹ�"���)A�� ���MK(#�Y���	�fRRIJKX�eD$�)�n�H'���$����ҫ���9_����b�F`Y���L};n>�3L�JCg�1X����y���	��� ��b|��{��2�Q�췉��k��X��|��7� �d��� ���}TI�W���\�nd/�b�
�՞��>$��������^f��q�$szB'��{���2�i+X��;~k߯1��� %����B��LN�F�1�^D^i1�HH�������ݮ��	�/��x�Kp2�w77a�Bў����!,p[X�ve�ٷ.�srK�(JW�J&R�aCm�|H7m�	�p2�é�TGXSix�>��MD��6*��I`��+K����ۛ�A>���{�V�[�=�yZ�S	�)ה#�	�QoC��瑈\.�C��jǲ^>��Z���x����`w����M�3{��G1`��x]g{���A ��J]&�
��i��0�y�GU�!oR�A�H �}����j���sz�^XTJR�BTu���)��X;_d��N2	�}T>=�$���`��W]�wk�?��Qۨ7	Rm�5�#���l����r�)�&4��"q���da$�2Z���d�^ݫ@f�wʶ��N�!@�V�B���݁s�O�"I$�iGU�0o4b����P��T�$�9^$�qC��r�q������B�H�
4�oe��$���H$��D6���3}�夾�;!�� mҞD���i�ު���6Sݛ/M�}������Ks0�Y�%��I �6<\�����&��R����������%��-ĂH�����u@�����C^�jC
�zM.���3���ɜ����]�:�U~x{�<Z����&��D���a���O�$�Ĉ��c���a��*�<���$�"������t.�)̘2�-�
�Q@�h"�n�}��d�qd�⛟f����U5RJ݃wP>:U���i*B�������<������I�H*&<��
$��$�
�j�"H�m�$8�dk6�?��\�s5�]/*�9XO�
��@3��)��z�/9�\.I�6�5cʘ곐����/��xaf��l�f�Y�B�X�meuC�X%"�."�Tu�h�1����R���:�Vir��l�٘C]k]E�]�$�0@��YX����C=L��%�֦m^�fm�6&\]��Ƙt!��u���v�"���+k����E��*��Bl������޶���B�M/0��I)����?"�ρ��D7�Q$7
�佦�#����	#7Q�90qQ1�p$�p��ܹ�A#��P$�,"9P���%��e� �.jа�<[�TO�̉�d4�����������A�#�xJ��P���؋��Y�^;��A>#\H$�����\U�N���M)JW`��H$Nk�Óu�4� Iē�A��]ї{��o�7�}��LkX�p6.t�]3��XL)�����.����%VT�igU�q'ǛH�;{a�]���UI΁!
�&o���i���5�u���`�ٴ|����7(f��}�G:UW
�]�.jX&f7v�񋹏�=�{e�晴�"I-�>��Mm3Q�b���3�:q�U|��@E�UO}Nz��8!k� �#}��]΍���S���[�t����O�"I�j^$|�.��UB�d�3x'*$BIB�.��&�����`�̓�|[���ϝP1�� �������-�Da�+�B\�M*	tf�aDU��挃��F�~$]>M�TH1���؞��E��N���#	BS,�7|�ײ�����,���P����b��ȾT��.L_�3v]9^'Ǟ:O�� 0�y���π�F�ˍ{�v�@�tl��o  �#�`�Yƌ�\�#�2�K"�f]M�}���<)Q��3zB%���,mD�F
��,��Eet@�"_*��wn� ס�9�iX��G}�uJ$D�n�ip�1���u��5u+�w��sƋz�9o;��@H�2R�P���jW-KGbi������oJ��P���(�W�Q�&6���Cs>b�z����DJ*m"����9�vB-�B��̑*&m��l�W7�]�1*Q�f�hQ�,��4�1�;���$�}�@�:Mt�����6��^��V5�#�ݪ*B��(�pV�Uy��=�+��T�����|�Q�m��'���%f,�&:-�ʙ��w������ĭ� �p�����%]�_]�6/�{Y�1{�w�7�(@`�{��Twll�$*��q4T�,6��lT�ڒ�+�.dZ�__~���\�.�>���ÆA�9fDzi��7���L�I(Q�;Hv�{;�o� ��2H!��@�����"V
�0��"bQSwQdI �izr&�nōn�FGH:�E�wH̢��&��[ܩ��2A;w+Ău��p��1@�&&�M"	-�Py �qA.� I|�zu�;����WU�4َw]�5��p��%&rB��s��	��+b����⦌j��{�j �����6҆V�ꋡ�2��X��e�-���4�c���R#e�&)�K��㑚Zͦ��]* ��l嚸��:���љc��B'ςq�Z�Xy�(+M��5ҋT,��]R��Z�\8���r<�����Bhs]��5˥\G;-
�,�u�u�6�]h��
=A�yܷ[�D���&!/��}[kȓ��Q��'�M�|��{���~�*"Zn�3�5�2F@$��H���"k:z�8���50;��*$�IDƔ���EZع��s&��D��T	�r&e7~5q�`ZW@�|g���Ϯ����5�w���^�v�Q�*T@�f��D7we�{�L�AC��	-�W�=BF�e��\��)���ܚ��Mŉ�B�����%L)IJ\;\�`�&&�-�Ȑ�:�	��A���wn����o]Q66�I�Ba!�0��nk#n�t�֬�gB��Z�T�,��Ԍ���eC��x!;��d���؛�B3�ۮ��  ��~$��~U�o�R\��7gj�_'�i�TC�-�$�ȒH�V���Ǫ��$�3CRT�IL(ڈ�ͫV7TO�`I �uz�Y�;hWpZ&�D�)]��p���O:̘77n�ߟ">ݛkf}H�A������N��Q��k�q-f��)p�L*��7}Q�U)��%}۱ ��A��ײ(�H6�@�R5�b�(LM�t����އv��nD�kk��"�*��˅'<a	��� S��$���>A�=���������=���F��g�d[�v5���(v;��~^v�益�,u�8@:=�zL{;��܋���vJG��J>�s��}�L��G�<�S7��cڙ	O2����9�5g���n�����vވv����3��!��.�N�9)ڴa��5�a�ߋí���� ��2:�C�;�tY�X9h�3ܔy�魐����loK��ow~��w�ꧽ�_�z��N��.���Uq��<g���-�M��ܱ�� q&�z�������4���fy��xN�}|��2z�^{
�ov#�icr��i��n��z�z{#5�^\�=&�7�uq���m��ǟv]��ro=}���Ĺ�����'��^����sy�:zs��˩p�=ɩ���ã]Y���5����#]��w;ɕ���7|�q���0��{��o��Z.C2i��ǝ&�ѳ��nwٶ��Ʈ�m1e����/\;�e�+oy���,�S�p~�!��v������z�'��Q�����Xz߯�;�.���څ�˔΋��20�{�S�#Phl:j��7�襊2Fʒ�����l�8	B�u�LL` ru8�%%��J[KqLw:�Ґ"7��fи'4!�
Y6��9)�1�iҐ!l��Y",-����ɒj@����d!;�(WR6���t	�$Ĥ�	1;�N�P�H�$C�;�t��҉ɉ8�{�:�o[�$�ix�V�7���� ��A"�� "v;��6��LLu$�ob@���YN�� Yosa{��6F�l��0$��RpN����e0*U��}�g�ɷϔ(g�]�ƍqD�LXn�^���y�b�K���(�m�Ú�m�9�ML	���%J�J"b�[iA�n�%��	YI�'[K�9���}�93(��3!B0�5�-�B�WHׁa�͵�$�%�v��2�V��� ��� �H����@Ԃ�	[�]%�B�*eDz%���_E�8#  I.�^$�6�ĖZӊ���h���$!15~9](x��4L�"��D�Bƛ�7�&����v+	4�|���^����z''�V��
1x�L���ʳm:�Z����j�������o=��ۃڬ�8H�O/|�cɕ�]���'�r7W͗�j�IÆA���4Kv����Ip�7��r}��G6
�"���1�a��c��
ծ�.�V�Y���*%(��V�v�P$����ϰ^���Z64t^�A;��D�����4Uf[�B����_WG����w}w�l3�[��*o,+v�fJ�Q�ma �d�(Esv��T ��d���c�T������=��} �� ^}"Iy�s���ý��i�'<bD�\x� �v���M�ף��^�H:�L�J����X1�/��=�*=���&d�����!,�S�kj��~�t���yn�I�i�RZ��M2�� ���m	e�̫$ȸ�!����t�M�KI��QQ&�Q�����M���[�+�������KE�F��..���X�e�d�f[KY���v���thhh�W,��ǚ���R��2�sM�V�)�������](Cb:]D.�WF�f�1)(K�0�$J�7o>�ÄI�9^1!�r��7oI��$��ChjҴiK�h�fR� �y� �����H�ޭ�a�͎�,MH��	W
�2O��ioj�U\�q߬���N�^E�wQ3%L��^)7<&|pC$�A}�H{۷��گ?� �k���!16�@�x���i(�/{h�@�f|Amϐo�W�ʷ�q����d��`4�.��^�A�5U�d�s��U_s��󋦫��~�I4�H;��^oN`rǑϷV�4�$�nUp�z�H2����B��ӳ�p�oY�҆��"�d]r��Y<!F��q_q+�ۀn���]��i[�jL��̵��2}�#/E��^�ںޫ�MM�� u�ʒ�D��f�]r7mЯt�3�q]��dC͐�N6�zS�r&���,�Cj����H4�UPp�o��TI��r�M�r)D���<O����
;�x�.�Q ����q����f�����M��4>D� SXM��c	hv(�2����LN3��"H<� ��A�7F�z�Qj����Q X�jNxĉ���0�ݝ��Z���D��fA&U��;�R�/,�S���n�변�� ���܆�[�P�k;w����3�5�V�7�Ϳ/g�H��y?�ٹ��p�P�2��b`����A���D���A#7K�	(�L�N���a�<�e
��2	�#[bTl��|��P-��6�uN���������v'�H���zN7v�YY��~D��vB	�̺7h��.��A�u����M279uϩ���*d��g��Ԁig�O6�1��2���Y�%*�����=M!j���&r�
$��>����-�i��t�8i�'<bD�T6I�i{�7��c"��޲I�$m#X0^��1v[��}+='�I��"_7[T5����8٢�WT�y;��^��y�:�f���^���͵Q�yw�^��2e�ݲ��߱�D���qA"���+�Q տ���t͢8@B�ب7wn�~�X��>�Xj�D؋��ڳ3ff�L���q�Є�P�Ѣ�H$\�%��x�in�w'���@����x+��(|sv�]Vn���(��@}�� ��ĥ���| {}�&h�0�� �_!G;]���� f\�5�*�Bs�&e�)��+��Ix�c�@�퇻��u�$Ӵ�1��1vy�G3!�H�iAm�D�}�̃M��Ll�B8a���E�vm�wVl�K��LF��#������,윔*���&�<�zK~ٙ�ϰ��_{��+�q2��ktv�z��YR��3f<[F\ܹ�뺘)�vыv�V�c�$v��'U�c�v�Й
Ci.XM��3J�V%�gK��Hl�eaI�vv�B��%ήb�V�27l�e�-�$65�ډ�����k�9�ΫSK��l����E9�T��A�q)P��cWll�I}�.>%(�)��"I��\2.8�"K�!Ekڢ�C��&R���!@��rj�Bs@�y�P%�>�W]9���Z��:��W�W�Z�Ƒ,��Ta�\Am��I�C"R�@���b�����������Z�פ}�umQ|�������w��J�YC�Ae;'�*ɾ�TI!�I��<�j��Z�ci���*)HNS�jJ�[�fSB�W�;"ժ��yT��y�ТIÆA��I�N��{B���Nn��JQ�SEݠ��Z*���Ѧ���(U�nn�N��K}���P�[�E��,�MLŘj��:杖EG���u��ΐ�E��zZ�7;P��Q*�\Y�	'���D���+^��k�Z�X`�� ��͠�'ED��M�u�K�/,�,�+�o��&���! *�kSX����-����Fʛ��6}X�^z����޵��#Q;�9M�p��7MŖ�i+�$w-��n~ϧ�f��2����;V� �3y���N^F$���k�
Dʓ6�� �ȞLFW�m������$�gs����p�Fv�$��SEݤH�mQ�6�Ɔd� �9]<����C��v��B�6k�������V��%{��g�$W>ެ������ �W�w��Q|��H�J%U=���I>�6�"O���x�Yetn<�C�bI�tT(RaD
3[�D�d�Q;Щ��ʬ�Iڐ$7w���#��7�mgE��K��Sգ.�[���B1Jq��Z�* ��U��埲�"�S|��� �4(����W۹�:�'�7��{..�)*�kӕ��A����ՋM�G��u��˞\��Y��O��^�2�"H���ˢ�q�����@�Y�s��A#)��.�&7�G�W�8�$�y�3�_t6�Q��ͻ�g%X��4�������oy{�}��{��JӋ���<��$
̺���D�Q*��̒IO��O퓗x��� ��vU{ػ���CQ7�ʔFʊj���ԅ�3k�n�&�
�%�ޖ��aDzZd�x�$���m쮝��wo�<uE��1PG/8V죞MmF+Vւq�@ ���6v21U;_-ߥ�7��v���ǎ�p��@����y�vO]�����2H'�[����B������o�ܳ	�vA���H$;�#u���s��a���"������H���~x΂6�γ48dO� ��'���WU{k+l��]Z옏/�_q[�p@h�M����쌼�|��T&^_`V;h�LR"6�J���B+˘�_-k�-��'���,���i�{�"s`ɘ�=ϰ���<pz��m�>l���"�\���?.����l���:�7�*��<(�������f�y<�(�g���S��{ۮ�X���U���"+Þ�����l�ݲ�ƻ��s��9���R<���O{���2��IHY}�/x/uD�#s��}��à)�\�yɩn"�=�}�f�,Kn�wkOw���^���7�TҥG��$�b���n?D'��;q����s�66�p]�_��y��k�����(m�_c[��+�a�#�{���,�`�\kz��v>��E�����N��J��'��8y{�}�qt��矽�}���n�-��E���?.���/�[Zw�p9�`�|
;�� ��O7Q������w	����w�y�:�_^�����#и�&dWlVDbР���~�b�7����F���<p��w��"`
>g�Yn��+��f�,��Q��6�6�ȇ	Ko@�l��)I�Bb�Y�����B��H�e��'LN��	:���6A�� !-�5��N)l�S��[:T��$mKa{��K{�C�e���(u��,,�v��v����5�RR@�I@Ʒ��ZY��y�[�:��Rsy����-��aM���5$DF�N�--$� ��N .�Ð�I�)%��8�t�� 8L$%�`�c�L�1�ע[e�^u1Ғ\Yt��8���08F	�\%�
��m�Pc�U׵��Ck5�e X�l�DXS.\�kM�.��yƖ�Xc�a��僴̡��[/�,u&��/[C.���S�H��+JE�09֜�۞�Z��ȗX�]�1p%��!κe3f�h���K�W0*�lMa(�K���l؆�ܗKp���	N�rR$��GMƨ8� zQ�F�[���ke$���)4;B�d�5�0�vR�&Ef��-��5h���ͫ�l�ۈ��#1�X��%��Ĭs.u��`��q�*�[׌�In�uy��l�.��KllX& ��a,��u�%��k�#�5f͛%��2S��k���ʪ	�[�XSc)�r QBڤ`v �#j6���\��_� ���G�X�R�i��KX.asa0�Rj�m@4*��% ���h.�T� òk0I� �.a�7�f�e�.0�ʚ��F��^Zv��D�E�i���I�H��\�Ц&�e���AX��J�5l%2�Z�4�vK���%�3@#Z�E��l��U���<<'���%�kWW0,6İ�.�"m�s���0ݐ&lpJuZk:��]��֎�Y����Y�fԑS@aU#n7��Z۵��8�1]p�rl�ui	�@e4�eM�� ��An�����[r�KWlʺ��٣�.�Wenv�=\�nAX֌ֹ,�e2�q�Zʚh��Z@34��f�6�t6��-��?�woL��V	Ʒ)4Ut��D�-�6�CT֤�'7�q�	q�#���"lSrڨTL����-,΅v����Җ"j:�M�M)�c[�%F\jS�`���B�2�T�:������k��J�:ь��uH�7jꬱ�+�S9f��5e٩l�9b�*��ku�bD �-�y�ګ�A��|�<�7�T6n?��	6���n�"*�RY�I.ܱ<�(HQ������p�/;�E	�Ĉ!�:�	)Tq뭊��sD9=�DPD�M`+5 |]�B�9(��{z�7�A ���'u�@�Td�fL�T����@���G��]�N��,�A��%�!%36:�h�H8p�����6��փ~�I��.�Әt��Ť���'І�6�(�6%�Q�̫�;$��Z��=��"�@���L"��P$�̃�[��%�t)�s��3*%Z�H3wR;�n��UJ2�!ҡVf��yq<���q�D'21�����R��QQ��.(�:lƱ���y$9ǭ�a�s��lo�Άj���Q�Ư"��T(HQ���|Im�+j{��Kf�.����hn�R��DR �M_�n��[�hD���N7Ż��O���@f�֯;s�D��T� �K�����qه15D��$�F�g�[=�ߤ!nJr����"A6(�Y��Q�yMz�k���XR������$�@�	��N�m]z����y"�$L�U6Y�5­��+	8��Cm AޠÉ�ǻq������	)�ʷ�W�P�\�C�{�8��I%X|�>z_�"A�Q�ṃ�D(�7#��r����-�GUqꭝ���7�$�z�8��QM����Y��T(HQ��m]3f�9� ��<&��wsYp\�xdT'��%"A�4���@ܵ;﫞�۹�q���	v���h/���[��5�m��`@�DBfe�@�.V�khEn��e2�S
I+\s�"&&R��2\�I�����$�Km"+��
%1e��E����i�����u^!���7����i=H���U"���B�w!�I �4�}��
|��$LʉV��ڈ�x�M A����\�	�q�~EX$�)���Ώ9��6�z��΋��u����F;^�}x&�oLF�1�{G���ω���ʨP�0�;n�D���$�-Vd���Z4W4���@��5��y(T��׫[�(^4 8wV�a��m��ñE]���Ro�w�����z�B�!�
Z�!��Q[r&@��ݻGPu�#M�%W���8{<T��g� �>��܉k�3������6pF$�v]�TÍ �H7��E�x�>�{^��I#;	�Fa$
S^.��uO������#}@��柝�%�:�[u8�BeD�U���-��	'r�svr!n��ju߉�-�.P���X�(Dl�n<o�*�ʒ �0�i:;_>�}H��/���\�S��b�������t�߹R|�^B
��R�s��[Fz�x�����n]���Q�ڀX���[���g%,	�b	X:�f�o+�X��c+QҲ�n��rԭ����m �mB���-���f��)˫�m �y�)��3.�Z�]12�eM��ꬱ�*l�욵�F�֤�-l���p�m^�sv���3l�#W*����?v���������s�H$49_]}:пBܯP͑$�w�(Cs��PKϞ��ʫ�b	�;	�$b�b��O����0"&&R��V�v]v�ܕ�*� ��$��"�d�(��E�x�.���HӦI$�z�v�V��wn�ܡ`��m�8��I��.�@$�Ɩ���NYH9M I۪&�����,��!M�M�HXꣵ��9�aDU��翻}Ѧv~y��pAkH|���v!�2Q&H&���r�V���~v01��{�4��_r��@x��C�����&L��l�॔/�u����x{��4~ �o9"��+�^H�Wk�:H�8nܐb&��>v��R3�u7�Y�i{[j�22�D��T��h�Q�cAx�x�k�Cr:$Q���pgyD�b,;y�Q���.�2����>%��	��߼f)}��f�PԪ�e"�
�F3[P,f����b�T��'�3	 R�uL"I�ƅCs��qSB� A>���6��HS0��\�#�牻�J��S��3�InD�AW�3y�����)�����u<�	�	��5ӂ���v+7NA�8t�v�5���,G7x,���<ALm��q ���zo�ov�����/��4����#:޸�l9�w߽+��̬���)�jv�76�#j�P ����ۓQ�U,v����Z�#���䒪�ؠ����#�/D�n��@���|I����7�>�-��>C�jnn��b�+��s,��GdZ�_����D�b9��=�G�^@�A[CG%=4��@��Ǆ���H�:���5�BIShĐAm�	qQ���gq��N����JB�
!]��BnQ%��oYu�H����nV�.�JD��
2�˱]x�0k� ���Km�qk���P�%�q��=;+�[̺_:y�T:�j~����G�5¬�<�}2�R5C}fq�9c4TD�� {�Y~㦠Z�"n��!x�:�t��[;t	H ���ͺ�]����\��O��_u�u���I�u�;�X�����xCϞ[K��=��ڴ$3����wp5w�+�pgyL�b*��{B��28���&c	��)�Ć۪���3rj�p�����R
SG��$�OW�]�W���"@.�Km��8�!%
!U��BT	�$nB-�TI'�e;�+��ܪ-T��J��5|'s�V-�
7�gtb��Ƒ^�РInE�,i#��@t9Otˇ��#9E.{��]pf���>[��f'�҃��^��+N��?Wx�&��T:�eH*$b����3��!��6W3Mj�Mih�Vn�Y,6Dy���\��כ�l�e�гf�i�[0�b)j�I6wF\\	��[p�@�S������ݦj\�n\iusSCȑT�t���2��.ɝjds+D�s��^�Z�Zl]���T�(8N(ka*�:�U|�x~����_����$�n�ķ�g\�h/q I�kڡ@�l$��[�0{��E�=��߻%pD	��B�<�H.�Z�����;/~ԳA2����Zq ;_�r���� ۿ]��#�t=*�"�_W�*�%u
�UQ$�_D�A�E���U�In�
�[r�Q
��ĒH)�����hȻ&��Q�p$�m���0����-m�v�$s%qbe)�f�6���6�V��<�玪L����$��ܢ�9�g5f��ڢI\	Zl�YS �M�oB'�Q�b5��>ڲ4沈a�&'O�5�0�!��j|u�|�_G�Vn	�rMU��.�5�U�%�rt8���}�$��$��� M[���[��	�#�2L��J�q��wh"��� ��	"� m�`7� )��Eh-��a�č��tz|K�H���1}��-��n@��%�I�����@�V�Q��]�w��� ����[Tl�����l���FB�����jm�ⅥK�@�Rb�\�RR����%0��n�|AsAI��Q�����04�	���a"ff=�Q2�|�8A����Q}�N`f��QeL�6%��"Cx�Q����O�n�ȴ�訥�0�ʕ�xn���y<r>���#�z?`G�~�LG�r��Ͻ4�����U�����S��<t�3{F1�D�:��?1h �=��)yi�`�='�C��7K�<��ί�%�Jv^W{}{O�O征f��w�W3�E�@��=sV�f�̸cƓ��6��ǹj$� �ov�dote��P���bGh�X96�@]��y�l��M�_n�'I�r5�X�W�g_u��M�;�}�����x�k�^;��7��T����ɞ�<c�>L?{�d"Ov��_zعpa3�tF��;�������)�����o����.��.���}�3D��͎�}�*6)���S�߾�cz7NI��ٻk���]8w�GQ��#n�`��;��&�`������w��� �����-�sv����UyUv��R���<�8;�l[�� u��y��|߆��_uX����V�=������ȯ.��꼭���=��9��<ӊ;��\�	�Υ�ݫ���O���2�s��=�%�|V:���֐ �k��=�s+��-����n�@D4�+)saK!z[-��o� �#aN�t��x�/[l�;�	il��H����uz�N��l�B�-S�z��Y-P��Y!b�u�0�B�������%�	ŀsKP6sD���IF�.��t'�Le$M���SAP�5MTJ1-��% j���K�70�Lt!s�-��{C�mzu�5��D�t�$HY�t��pIց)G���%U�����0�y/`��3��ݬ�`�)�q�)N䒒ka]�$�:^z3^��]�Z��У���	P��$�%�HB[HN!Ԕ8��K	B6�vպ`���@���.u�? ?���F`�fe ��I��ב$涨s�;Su~p�7��6��]��ݯQ�y���jD��9��;���p��W�t_!3A�ڥ!J[��H�*�ܛhۅ�R����R
R�U��[u@7�@�^O�r8�y�9˙�
eLZn�A&�	=�ed��	>�{B���IU�+Ovuj���Jd��%�Ԭ^�x�.�B�؛�y:	4�P�9Ă��j�L�5`��E�DF�QK��I;�$�_=��z�8���K����Tu�V8! �8
���1v���ug\MP�uZ11wRH��i���yQ2��T�wi;�Ȅ�k7��c�,��#��k����\�����'"��l;b�{nJ&�g����(��IBZ���D�b-��گY� �N�H�"���N�P$60���4�% �!����֓s��)�
:0�� �h/ldE��.����H(�0Uuő$��K܅]jwy���G �ە�e4��33��y]wxT݊,�	�M	��[6�Eh�\3$�:M\)�b&��Q ��rU��Ps�H��}���@}�wi�0}V�Y�}�:C>�Z���;K�{��
��Sر�ϗ�0��d�� q�_��3d�}�M��d����!H�fm�%K���`C��Ql5��ITj�Bk5V6��9�+e����Ke��R�
mbZ,˅*c\4�v7'[��"�q �R%����2Iv��F��oc�j��.6�(Y��Z��9�30M�]�V�p��ZD.2�m��6�lh���be�V���d��y�.�|�~Hwn�w�U�N��D�N�Y �逢B1e��"z�m��QŐ�H'i�y��ө[�W�+D�`�3B�R�;Wʉ7��� ���5\�����j�*���
˫R&%Lth�D�h�n�r����o{*��6������ �FUm�9򒶥U7$j�v��t�c��+E�?���g e�`F�4�Pf���2�,Q��A��Ch�y�'�ݷ�λ��b:`���8S�֮T�,%�v(�����}�Ò���y0�ƹ�,�Q5;�n̵�!� ��Bw�M��L�{�]gLF$1~���!��a��v���7������T���e�=ꦭ��_���NOmΎ$~Gn�ð_�V��B@�Imm�IO_�؉ŵ�ň&c��:�E�c}ݞCX��6���xFX�ő�iFN���m+�a���6{>����A�����l�bG}��q�lD$@���mq����W�޳�����x��bQ�߷h��(�6h��S�-w�'j�K��QlCg��XW�[�f9z��Q�m�fцFF!�Mz頱Ƃ1C��
�/��W6!���½��2�6d��s���]GyM�j��J5Q��1��̱e��_;1r��v&Ѷ��1�w�XF(�4��Ҷ�J5��gޱe�h*��ѳu�z��3,�"͎�����641iQ��W�����9�mC��Ƌ��h��Izz�ݍdLȽ�{ e�Lַ�L�n��5L���FX��)�4���m��u.SrV�-#1�z�#���i=w��z��gx��C`i24�ˍ��G�!���s6!������]��3Y|ܪŎUK�fZ^�Tj�J1�l�w�2Ŗ�4A�A�����c�&�NTn}#gBY{ ���.�i;�t˯|���J��U��}qO�\�k���q9�/M�ⶣJ5��gޱe�h&�ro�]¦t�6�{{��{�|f����X��vD�Q�A��6{=큆e���9�nц��Lg��S1F�՚�Ch�k��VIwC��-�,#=�n�#��Q��߷fF���:>Q�`hz�q�lCb1�������G{۴e�l�c�;u���f��i�[��9V-˶�a!�(Z��}~����M$�Z��k�J5�a(�gݳ,Ya�Dh����#,Ya������U�bJƣ�׻�Y��p��J��mS��n�#�$������A隌C|h#�7�{ e�lCk)���h��F�0�:1��f��k�0�&��<�\�䬣LCe�\�0��Q�Q���`e��c�Jf�s��;8�G�Hc:݁����G��h�2�����16��0�DY�����]�}7���Ҍ ���e�,#h�Dh���e�b�Ҍ�z�K�sY~�Y��?��=a�ύx	� aG6���7K���͏5[�Mְ�B6?y�_`�����5b:2B��~��}�� df�X�����77�.�SbG}��0�p�Ch57Q�Aw��v��3l���`a�`F!�k�գ2���vz�E�Dh���L͕[���ic�$����Q��c�GLi�Gmr��{�/��e]�L0��{6e��(�h���2�X��F�v�q��Ƃ�qgq��^�`a�o-q=��іd`FN��U�nQV� i�ij�Q�m[J0ֹ��hT���`a�mh��;�#,CbK#;^��6!�9�ݏ�4�{z�y�h6]oWWW$�xlCh�wv�1$$A����6!�3�ǷX�\�n�}�4�0#�5�jцLQ�LQ�h�z��/��.�$��LCe�^��'��7[�[K�F���3h� ��6�j�q�m��BC�׬X�5���c۴e�l�95UX��Լ����Mu��(�Q��w`a�ŗ�]�2,����Z0ű�b�#J&Oz��cQ�l���Fe��s\�=��s��n[ϷrŖwn�T!���O�;B5��Z�2�s�ۤ{�>�#�v��=L��z�t&()*2�]S!�E��.�$�D�v��z�۰Gh��:Ĥ�"6�4�v)a)��r�ЈA�"=��4���&�e���@"�ڗKr2�5h��Á��(��A�Uqen�S:�d]��.��j���9�30K�vY�*:V������st�Qم͹�e��]23(ʄ�%�w%@����O�=��X� ��=n��A�0#9�z���}�9[�f��q,5{~�,21F�0�D���-�4C��;U�]���b=���l2ҍF��Ǚ�xYh�����Xdb@��!���{^�3�!��G����~7���mb;�>�M�.��f���j��մ�ُk���6��w��b�ib��1F�Mz��cQ�Q�F{���#2�C�ߵuud�[A��F3��J{��sV�R�Ch�T�7md`Fc]݁�e���=�jц���Y�����Fb� �/LCh�~�oSWD$��LZa���e��Ch���2��c�����|6��#@���!��$1�����Z�{ڴe�����F:�?ݝ����wq0��[`��X��������v��gW�'�~���LCb�9�ṉe�LQ�m�h�ػ]yۮ���q�~��!����23��,4�Nq�ꭕY�A�=�r�#�؆%������z÷�3^C�{�t)��6�}�~^�c~y�:-ocS���������R���6A�3�� e�L�6�=�jіLQ�I�0ֆs<zw�{ӌChɎx���*�yE���u`a���J55�j̵�d`FF�XΙ�ۮ�\�A����k�V`��AL=�jі!�==�MSr�����S]�w�{:KmdQ�b��1�21e�m4F�sٴa�,#F��Ki{��׫+LC`pdf��h7n����$��؆�x��8<��Ch;�NƂ<e�8߽��6r���fFj4�F���0�)�0��zSE�F���ceb���3!��U\�0[68�[c�Ժ����}���	+�����y`a���J5=�f̵�L���N���m�y�W�Y[B׷�@�.���jj�P�J�is�J��7�c8�6/3��l�XF(�#D﹜#,Cb��4�������Q�k�����N2��Xh;g'v�uv�����Ǝ�����$$A��v�G�0 ��>��������4����U��Fz"9�>�M���ʳ��]��=��\���1u��,�׀�<��F�j3��a�(�&(�4N�����&�����*%~�G���gD�a�z�V�iD�h���2�Xd`FF�)�]4�Ab;�z��k�;�j������0�u�FX�̭��֩����@�4�SY�j�Q�Ҍ#f;�Y��,'K��I�	�a�4OoY�2ő�b�#J2k�M+�(5��{^�e�h&�����ўq��R��)]�,sk�u��0��f*��jIJW���T�0~'�|
��6G��6���LCb-�=�{ e�m`�B��J�%���{>�e�l2�A�w�LCh�5���	+�����a�iA���OxQ�������##�Ov頷�����s6!���޸��{^գ�Cg�٧U����0�>r��mu�D��wve�,#bF��e��_;����-�#L#@��!��c#=�zŖe��Nq�Iv��IƏ{��w^���|b:��~�v�G�1�߹`a�L�6�wڴa�7^λ+�ߚ��0�R�,*�%��nd@�ܩ�`��]��>W��}TxǕ�l��ۋU�a���@񊦋#DY·꧒�r�(�XFc�݆S��j1�[����X�g}�������24s�M�4�"Ho�偆!��������H���x��Nv��l�ĵ)�)�b�ĩ���CQ��:Gm����_���/�L���?N���c�ҍF�b;�ẕe��DM�.���2�6'������e��Nb��cQ����{ޱe�h9o���VIQ�q���2��6#�z3̙@�꧶�8��0#&=�`�#5�j�}�FXe�0�Q�q��7�"�����F��j=I��	+(����~���,CbG}�Y�������g;�|������lCb=����!���{�Z2̰#5�n��X�T�����Mh��.Vtc�JڃJ0�g;�Y��,#h�����b��U4���y���m.�df/ݱdfZ	̛�۪�V��!�w�݇X� �H��uNƂ=��kAl�d=�o e�`F�J5o�ݣ,2�����bGR�s��0����?���{��2�����;���>��z�1���!?ovj�J�����?;��=����S
ҷ
�T#s{����r(��b��g���
��ۧ�����N$���W��9�ܕ��1=|�ͻ�y��z��#�F��	;��^,��=q`=��?����;�[�;bF�g����������!��Q2�bZ
�T���U
6B�ҳ+�/��#1ՙ�Q�y�
'���i�C��I{oT���r�}�!�?3�/��a�v�y��=����s0e�4<Ʈ���6����+DN�8�՗�(���0��S�Mg��,���j��I=Ցr�y��o�q��?_y�����̯"�1~�Zoض���w���-�z�v��}�g�����aL;E���W����=�R�9]�q�$3O���W����X^�&����㷎�����{�mdf��{<ފ	�W�\�9��x\�B;�7|mxM��s}�r�ݻ�M��?Y���.%��1y�t�I3g�Y},�4��ޚ��0R̋z��|4�;�W�����8�hm�@��l$��R@�d�D�'JK	�;�cy��������ŠYm��Jpt�II		�Ԅ)%$�I5�	d�iذ��$����I� ���$�N�u8���N��  pԘ���@1��N���!І8'Y��Rè��H)Ɓ�1���F(�m�����%&1&I�8! �)H�N�m�@��8@  @�B@(ƴ%v���Mi��$!�� �P�:v( '@N�	�[@ HB 	B�%%% �D@� v�(C�x	)� �!q!BMhp!q�8��Ҁ w� 'BB�	pBv;�k� $��!�B O��|��E�H�<�鴨:l�9el3��h��#�H�kbmm��4�;sj�d�)6�-�:�
Md@\�2��n�##[kÝLM��K��	��mZƹ�@�+d�j��Y`jܠ��qe�J�5B��k�X��)��F��J:,f��&n�.�fI���X4-���9څF��)���GCLm�b.�\1�ѕ]���]�j�f�WYJ���&5Ŕ����JA�[a����*f�n6����cH�������Krv#F9����kj�n�����qq6��`�\�y�Xڍ��br�3RR�b�����j�e���Z�n�f0s���Z�8�[�-�b�84��A����b#��K�8�j�k��0Lj����Q��4-Ԗ3YklF�BVܵ#W4�f����#����8%�Yn�jp����
���It�e^�]R�W�JM��	�a6��)k�&cL�L��
�����ݫZ�,p��؅[�*��Lm�rRb�q�`�ea�[�*1Ђ�ia\%�=l�Kh+X���G�)@\�]1�����:�]��;:`X̓FIU��S �5�ōs����XכEТ��va1��0�Ü�f:،/�3G&&�-+	�̄�]�U��Umʬ�Y\�Qc���V�*勭t�$a��em�.�.	X�n��-��jݮ��2`b	[���j�eo+wV�E���3])�s�2Vܭ��It&�l9�ַ��X��`��gmm��"�ֈ�÷А˴��2����1^���5�É^A�J�A
]�VC!�Ks��5CΉ6q���m��֘s,b�\�rƽ��fL��X0H�2��Ј�,�V���:j�cj-W/�v>U>�˗~F���wa��,CbF���0��#24{�M��jw�߻��w�E�g]�������0���FX�Ξ�fi�E[��piMf��lCa��9ν�kV��9Y͛b����=�o�ز0�漢VF�j0/���ɞ���p�'/6.��A5o���t�T�m\h�5��,D�D$@��!�Mb'3s�;��n��8�6�ҍA��h��F�0��w�M��zsUn^�-#=�z�������譆X��6�ox��Yb&F�On�m�1�Ͻ`Q�of6!�{�ݣ����+շuv9U/ a�|�S[�j(�6g�ݙb�s���6&�6�g���,�#F�d�*�V5Pj0 ��羱e3-�o���=UT����!j�1�fJ2��3]4�Y+v�W?�����n�{?������-b�D[�v4Ƃ20#;����2��z���y�[h�ޭb1F���LCh���~��S.U�b��s۰����i^��S7�P�?^)�Jcҧ�3�+;���9�q�T��=aQ/
��y����ϝf���冊�7g���6!�}�h-Ƃ8�BC���1�o�v�{��{������$}���I3"QV ���SZiF�Ҍ#g��Y��,#h����Z��z�2���b�҃&�TҶ�J5���}`a��-�r����-�m��û�{��s;�Cb@���!���l�7�`�#5J5�{v���so�jة���@����h����U�$�#,ZFwz偆!���h���2�X�8g��+u�,Ch}T�qƂ1��7`a�o-q0���FY���\�B_��߲����6��&v��%[��&�׶W!Z�U�ϟ���$���g���*���bٞ�vdb��4s�ݣYa�Nٞ^}Sa��FLz��mF��ٮ�,�-7����WR��:h4�G��Xe刄�+�n�@�ʧ��1�`Fg]���d`F!��{v���a(�z�v��4��5M�#�t?Q�t�uxF��3>��20��Q�ѭ�ve�� ����_����2�kK����;�2���gr�������wQZX��E�	����v�U!�3�F�'�!�w����G��h�2���z�7)ջ�f�SY�jo}�1̾��M�4���k���6��a��#��U4�Cw�w|���3��a�mFdg7�X�̴�K{���É`�+�z���������v�����Ɛm�l�u��`F!�{�ݣCa��0�D���,h��z�;�����*z�%Ҷ�6���If��nZ���;�������U�$�#l^Fwz큆!��F����-e�lCh}T�6����>;ͱ$5�j��`���F�s۴a�lɬ�+n]�R�� a�iN���lCay�Q��Xf}��a�(�6�{|��!�e�i@d���V5Q���7����e�^=b�̴�;�����M�h���,D$$@���cAh##3���}Y�y�g]lCbG9�Z0�6�@�ꦋM�o��ͺc���Cf9�X^s��W���A�!���h�u�2�X����z�SAn1���}`j���H�D��>�E��Q�����U1���	G],�������[��{���
w�l�ܜ��(�� ���4^��F��Þz�9U��h1T�6!��1FwZ��b�����3�e���3�fц!���N���mF�j0##=��ő�h+��k���٧���.�b�kz����3�y��5�c*5r�����/�ݦL2|���@}�����Q��ۈ��'1p$��;�F�TH�Ue�4����s��!�O� �[B�t��i����vtuT��U-�����X!uϠ�P�_R���N8�Ou�^�7D�P��U��<*��#�+�k��Wn�I�w[����%�H%�$R2AR��@��uJ/�"�:�S�qğ:���n������+!Qs[z��z+�J_�L<����t��\�v�~���߇G���>%�s+��l8 ��k���0sZ��qi.��(ݖ��e�X��cB�vlWK6sf@h��i��Z�iih��l0r��qmZYw,�NNu�=��4�qS$!-� ڸ��������`�밵�١ֶ3_���n�*�����)US!*�Y����d���v�&�	��v��P�mEj�O>}<�d�W�p��]���ʾ�~��mlw�@���ضk��S�A��W�� ���ў7�0C�$M�eQ�T	+�����g.\rf�"V���9ߝy��H����C�u@�Cn�S��JB"fR��0�M�����Т׶�E�٨��˽[絼+P��B
T9�mH��vs:�Z����m���p�WW�U� NҪ�P騥H�Qη�Y�ɩRm0X�U���!�$�*BηD��hQ'�I���*��/��=�Txk�rfJ�VTzz�[�[X_k�؇Q3!��S���w9�Mt�ԣrʪ�;j4�.�S2�r�$�	-Ă/!*/Ƚk��DZQ12``Sʠ9ĒEM��Y�|0�m�$��I+���Q"!]���U�w��P$�Ϊ�$�z��-�BIN�����¥!3)р�A�x�]6O��j��q �|]6���9���6��ve��"٢��ժYkH�tt�3V������`��o^1@^D�I>'��	{�-ӭWd�+��w����B j՛�J�O�5�v�Y>!��.�B���*M�>�p�Q�V�6q��>׀iiVZ�].ii,άW3ԥh�1�'&8!Y�7��� ��r�j�����٫v"aY:�0Iy �n���"'��1�OB�ב��*�'����@�os]�?�/w�h"8��0�+J�ve��	�U��w	�>$��I��ܡ@F�{\�����y��fc��	(%��&mq\���֙J%f�2�fe&w�I ��B��yT[�Q�}y�b�mD Q3Zy�(GtՍ�z4�|H}�T>|�V���\��
�!7y� �ǔAG/��*����_kB�:�Ux��]�S ĥ7`�E�.sHwmQ �m�Q ��NE龥�U�"�zTt����r�wb�;2g&��p����~���(7�۷��V��}�
�HJ��$��p�{R	{��@[ܪ �p�5�v|x��[8���X�Ոn#�e�T�l�e
�e��������)
�r����[ܪ ��I��n�L�극Tn�dF% �̤�$ƃ/�w�U	-đ������j�f����;Q�(%���ܴpY� 8WXW�NAuk콠A�(Q�A��\���
T�5���V��S�$�{"H �n1+�y�o����JnǍTI$�V�{x)�%�Un3��ۡK�4��ؾ_1��F�f����L��4¨A�u_]���;"�÷���m��o#���l�Ɔ)#�Hn���IiY��6rv"���-�-��1m�n�Y���!Q�
�d��u�LM3mj�amul�F�Ɗ�X�k3��lM�uGB�B�Y�yt�mv���`�4Z�d�k��2�:���l�Q�uGA�Ŏ̳E�J��*
�sʹ��LZ��9i-h˖��h|�IQH�UUS;�D税A�*�����|��ͻ?O;6~R�R����� �qqfd$*�~��Q��JtŅ�/�P$��H<�Up��q����|zߢs��U-�����V)�g��߾]w\���b���������gp-D�@%��K�U֮T�H,H�p~�j�U*Y{�v몪�J6���E�I���'���ߟ��uT>7B**����ԷGizb�9���\�����HD�	�ĝ됁#{���}53��itV  ��xǷ�XUЊ@����w9��j�,6�E�-Th�v(�ꌙ�7���r�o^�6p���|h�(��$dCEn�P �uTI�҆l�ԌQ �n�\\�P��ݗOU�j�La��[�	9Oj�Cn�U����1)Qn"Cz�tH#��Q��W�s���*��x���FΝ��eD��o5Q$^@���s*�\���O8����y���l�Xh�׮қR���9�M36@�GTZ�_>y/�%6�TU���3�w`��{d�M�q�}�x���SQ�V�6P��z���m�!��Cp$Ƚ5�{�����Uk!�D�ɑEV�Cq$�p|8f����V ���q�L;υ���ĥ5S�����3�B��"��)D�'���O�Ϋ���֟�u��۫-�o�����
�{�~������z/���o__2�H�~��9�����ۍ��%b�8�og�~}��+x�C��^�߽ӈ�:�$Q9�<�����M�Q�`�;.\��x� e5��i�����V> :�M�2o�������3���=��-ʼ|�.m��6xo������r�D��o�	n�y����?���C%U�ǆ`>5{��K'��00
|9�<��������4�@Э�������{�j��1	���H����7����v�8Ｍ�/���Ik��0^��T�=2u�L�6������T�{}1�f��������|[���c?���D�qy#�q��*w�{u�C�p����l}�N#�������מ�G;��9�O�ft4���^~�f�K�ɛ���;Z!=�*���}@��)Yˋ���9�7Û��q��VC�-k/�O������)> s�|&q`i �����)x�$�!NBbX q��B����@ BoS�/ '���-�H�!��� 8  LP$ � �pBR�t!Ҕ ��K�BC���R�d���ZwR�� kנ��Ԑ��B��KK�m�I�������-���ٸ:@�� ����  ト�:b�@ -��������LuR�@��RX@��$����628F�I1��BS�oXMBÎ��l%,%���ZK!R�R���p�HBRZXI�JB�m��'b�p H���[x�p)`ZZ�[-��B
[Ɛݭ_���ڱ~k���a�QT���t����9`}Z�]TI$� �o-r(Ϧ�ӵ�&�r`�
�����$�w�S��u"=n��ĂD�oomZ�nD�����ۑG29C���G��a4�L�H:JݮV�o~6���'W~���� ��*��W�bNfl[x��=�!�((��HN�;����/u/q͉$�o+����wzg���f�fҀbR��]�y��Kǵ�n���|��� {ٷg��������Eϲ�_u�Hx�����q�쎷�n"im��ֿf�Qz�Z�{'W�������n��B}���Ʒo Z}3��@Nf�Q�ffƫkI�ڗCr본��U�"\	���O7u@��k'-b{&'�D��vj���8����T���Pur�����M�`����$�M�z�o;�=�����M3�H$|�&vL`�!69�o���NEt{)�Ux����n1��U�]�� �QJ���a>7��$��v�v'o#<H$���ŷuD�뙴�DJJ��Ct
�ۈ��SyDA!���An'
��N��I
��=.��L̙�qP ��H��Aͫ۴!n�]�����y�a�+��jd%�z�DM@Wܶ���{�nv��d��Y;�<��1o��n�����ؿ��R�\���Z�+7��"�R��KK� p	p�ݡ�����7laIt���di�5�U�SC��V��
֎�e�ftH�L�ؘ�n͘�S0��iw)r��F��[tҥJ��
G�Վ��ҭԙ̳E�J��0�(�o��l�0��B�J�ò�PBY�b��~�y>��d�85^/�<��O8�U�]��q���6`�
���� �P�)>��1�̠OgZG8�NV��O=\�rg�	������� �/�n�3B���c�Cq$�� �QJ��櫙162w�;OUH9����m�]R�T�'ʠN=��JD��%�.�Ь��5>�ۥ� ۉ$�M�@"eҫ�'o��]�v2f6�P�mtݩ�nʶ��_=��M��v7g�Hn��n�*��P��T%�ż&H���% ��6�3��4���I���a�<}�kUc��o&��'��j��^��g��l��j���\�3�ؓ�M�D̶�3F�un�aڌ��32��H �ו@^Y����ȒA���;�W���&���n����,�	y�Q$�<�.ֽ�gLI"��9��I�Z�}���~����T�{� ���S�	��QJ�y�t����f`���]0o9ѭ�i
�m��a����2ҁ)-��H$wʼCo���+�W_�%��	7�����A+���5�́9o��A$t�|�2��Hm�Q ��3b�^[�M��q�T����3�uo�sq�q��O����
*:���anmO�;��\�7��#BB_��|;�zo���Uz�������@�u;"'&fe �w��d��|����J� s>�݂���]�f���]z��������������2��l%�^�TA�*�%���^c�X�2��8@�A��L��-#`4q]f�B��r����?Dm	�*o�v�`#;���n�3�d=��n�j�oqQ<��m(	%vU�}������Z{��9�j͊�e�}�Ǯ�y�B38���>�۔O��$�ʕ��NWU�M���$p
�&T�D�wL1U�'�κ �qǤ�7=��:��V"+�*��w;�RS��xu�[��f�>�#�7�����:d�L�>Ws��>���<�,*��I-���  ��Q�����}�g� >�m_��>3ya�m��:�����Ƌ[�Ȁ��c��R�\���>cx0�e��I��$Ws�0k7a��#)��3c	�!ȨP �R6���1n�r�3��P �$�J|צ����n&�F"RWf�$�MSj�P����].�uA`O�	�U��L�"\�VU�ؽ�G�P�8p��ڰ�o�}�au�@�	TxU�L����Kwh�KǵQiQ��U+��D�GSʠA#[ڣ���!frylmPǙǏn�ب��HV���Q�;���{rnu [�c�z�a��y�y�Z�F��J�I�8��=R��X婨 g3hB�)��f�S1���u���c��9d�d��D�;Z�i(��6ۢb��s`��WmL���0,�0m�h`� k̺&(b�-h�L]Υ���Y���RT�4p�h��:�ݛj�I��4PK����dR���FjS��)�[�� 0�QX��Аw5�US��݉��)$��=����[�B��w�b`H$�>�G�cvL�H�Bl:x�]�wU���8|A�����6 ���K��	x�0��t�
T�����B�`[qZ���I��B�m�P$7�h�)+	G��e�X�ymUx�=�� �9�q�c���{�v����D�@�'&��Vp�p��,]�Hǎ������A]���^#|�J�ˉ�K!*�NJ��T1���)
gQ�����>x~ݴ�ύ��P%�ڠA%����s�E�m�೿}v�eO�s��$�Vn�E]�Y=p9���3�"��"�B)	zd=}�<��#ꯛ��甞�E��2X}=�fzI2��~�@���]�V77Bb2]�v�ġD&���(�f8���Ҳ^�����߮�[����L�*T��xU��ͨ"��@�Cp$���9��'�N������ݸ�	DD��MTI$W[N/5{ �Mx���	/"A��Qf�6�Q��"0��5�7���S*��]N�%E"�UT����O*M�9>��bo@�A\�f�7/,7�T}�O���q3"P3b�=�VH!=��/���$���G�Н�i�Q>ՊA��3)Q}@>���A� ���~K%�!�{߬�>��,�g{H0��s���������{�I.n�e��9*@Bj�v��/����$@Ov���;������Q��J���w���
v�.ha���NS��-�TM���.�j�3��1�
�H��[i)���0���gU&e%)'a�𙈉I[*�
�yD��X�����x� �_վ_��JŌ�k�Aq�]�-�#^u{[ž'��܆�i�1��K�;�W�G������S�<�(��ռ��[2�)I%R�s]��xR�.Ѓ�߮��o�g�t�d����#��h)�y(�~:}j��r����9�����.��.����&.����c��9�u�7`��Q�'\�^0�*�$�{�b֧oo�qO|�@~Q�Ȧ�F�f�L�vsff�5@�GT�	$�9񈘀�K����m�U	n=�WG��eP ��@��t؉��fp�j"��y��Tt3	��7~�؄{\@��o�_�$ݯ�8I��qE�V�
�q��]'5�����ZO�k�(�yĒ�ݛ�����^[����Ps� ��Т$<� �M�`an�
\��!32�}H$ּZ���e�]�c�(m�����>��?��g��lm�����@��"�?�$!��r.$	B<�#���5���
QU�Z��������,�6,d����2L��V]cEc	�䨆HB������m�"�M^T( �`"S��|�S$!��&�Z������>X���A�>�A������Ȱ`>�R�5VE��h?��v@�B�|mB!�7����A��iXk�!!G�Pw���_��K�� LKI/���#���I $!��6���g���">`�#�܂��?�����q���X_p|����>�� HB�����?���hc�����HF�P�e~�P����u ��̆
hD������X��g����4�>??��fT�?�b� HB͟V��1ʔa��}�c>���@B6���.'m���04Ҕ�O뒄}%��س��H�|%���m�����/�,}g�_�/����a����ꋈ�}A��}k�#̴�������D�?��~�z��?���MD���#�Q&�P@�)#'ރ�>����d���g��B��"DZH?��'��~~�Ծ���K	�/Ҿ�����+�%���A�3�-3�$!���&�����	�_����6mal(c?�h}�A�$�	CL����!�����<��?����_�(%�䙳 G��K��� $!��0m�*T?�a����M�BB���h�}g�K��»Ԙf��P�� ���Yʋ��b��qh`�j�z��� ��!T���~ӨG֑��;�O���BL>k��B_jh�������w�|��t�?�P��(~�>����~�0���G��~��������U�#����#a��2�}�⾘��G�I!���I/����6���!/���Oj����������:���� �������YcZI5Hg��ac)��?�1c�~i/�������#�_���������������/��d@��#_�#��_���j�?M�F�~Z3�_/�#��1����>͘i(�B?_���	!G�A1/�1PD`#��~_�������$!����44dV����,�a<�%��cU�i���$6���x3��~>/}����H�
�kZ�