BZh91AY&SY���t��߀`q����� ����bC^�    �>T��CZ	*�
��z�R�)k6�V�mj�Me�Z��֭5B�b+TkfSZ�i��k���4�[l�U��4���KYl�B�@6�X�"���E�6Z�5�hɵ���i�,�6iVլ��2�̊E
��6�j�֖�Lڔk��(3J=���M�eb�lj�Z� ���l���XkX�֫R�j�Ҷ���֑5�Z��T��Yƥ6Y��-(�ڌm�Ŷ�Z�h+R�Z�Z�i�cJ.   ���t��̺��M����D��c�NՅ����3Z�@v��{޽�P�v)��R�f��e7�Wu¶����Ǡm�y�<��j�͵[`��KZ6| t  8����t������).�.7�-ҥ62������Nڮ���*PT����z@��07���UIJ󓎖���T�^�=*Wb���j����Խ�Y�f�j��;[fR����g�  ��AU�R��ܪT��Jg_n����ҩ�WsL��jR޻��J�J���.Uݽ�I���UJ�J����W�ӧOZ�^y��J���K��"����T��-&֍W֮��j�S]� ���_Z��]���T�)nG�^˦���L�]� ��=��*J�С����)�����j�!*���zJT����Wާ�>��},o�����^ڒ�|�MhҨ�[��U-�π �{�f��C-�w�j}�Tw����U_g��N��ཥR��u7tЩ)���*��{2oS�iB��;sܮ{�*��m7{�^xJT�{���*k*��ힽV6֭5���S[)2ʟ  ���JJ�_m��{�t��{އi^�ev�eޚ�ԭ�v���z��ҷ�J�n��Mg��������RU��y�Zn��ow��R�ޝ�v<��t<�.����d���)�S
�_  n�U|낕]Ǐ<�R��n�ܩJ�큸�Ǒ�*�s�m�u�H�{.��U%#z=s{+�P�3����������Ίi�<q@z��I��Vm4֥&Z��T�|   ��}*�z����kV�Ҧ��h���C�K ק�����8�[ײ(4q�WT�n��S�:4u���v�٭6�4mj�4��b�   ׾��ZWWU��]��w�:��yy�Ӻ��Uֹ�;�Wlp�t{��x���{�� Yޞ=P=�5f��k
��)�f��   �����I�n=5�uڏx�<WuW@j�� ���Zѡ�.{gzP���w��^�n��^����ht>   t ( �*R�i�	�`�	� ��ъRT�       �{%*��i�	�F  L "�� ��� h 4�  ����i�@� �4����Rh4�2	�O)�f�zC!�'����o��~/�>�3�'����9M�!׏w9M��^������־�O��O�� *ﯞ%TW�
 ��� U�� ��<	����O��?�������� ����x� *��~��g��rC�EW�����{��?� x�2�a�`�d�������e=aXC�@�=dXC� ��=`Y>���z������=eXC� ���� z���!�+�eY�@������W� ����=e}e~��� z������ z��������Ք=dY��=`Y� ����=`Y�����������
/рD�0�DO�(�2�|dQ=d=`U=`Q=`=d>�('�*'��'���*���'�*� ���'� '��'�(�ـD��P��D��eU������D��P�������2������=`A=d=e=e=dQ=`=a=`A>쪇�*��"��C����D�T�S�E�U����"��*�zʢz�z¨z��z�(z�"z�z��vA� 0�>������	� 	�*��"�� �a��D� XS�(�������?Y� ��=`Y����� z�x��+� z��'��ѐ>�݀>�ݕ���>��e~��z��C� ��=e}`<e��=e}`YC� ��>���
zȹ��O_�@��4��������z�#S��j��u@MhjJ��.��ǆ���׷��-��Tw:6NB�m�5<����kd
ZXnQkm��RY�Z��݊U�+Q��E�⳸��ճRSm��o��n�k]�)kQ�a�C]��jЩ`�ām��B�=���a�"�Xԧ�nk#b:�֫�'e�ɮ �3`�h�B �5u�Rk5�����:��Ӣ�2k��Y-�ZV�ZkJt�ڂШ��څo.�%K@�*ee#p应�'�Q�&;��x �YtUФ�WZ���:���aJ���1�+��.�E����pe�K�;B�D6��x/P[�pݱ.\@b��L��˒!z�6)}����S���b��˫я-V�óat��6��7��'%����VC3[Z*A�l����J ब�j�L5?:�(�7�V�nq]n���Y�t�0���-�R���M�0V��'�)��J�f�On���Cմ`���8��M�� �!�%"�8b��b�����Ѡ��0h�ҡX�Fm��R�Q�/���[{�Q�"Ax�+�)SY�tӻ���&U�f��k�#Z�1�Qց����j�͡�f&F���f֍�y��*��U��CW]��-���Rwh��q��k��X� ���u2wY���&�wO#P�����?+��'V�`�`X�vL�䷑D1�˗V"�'lZ�i���*{W	¬`�e�q�:6%�0��p�����K����L�Q��A�aѷDCX����2�kB}M�\��ҡn�V=�g56�6P�/oA���0<ժ]�u��t�l(��3%YC2��/`,Pu��e�n�0J��:��2若*X�!2KqJ@�f�(Ƴl����]�Y�����ȍ�%n<�r8�1еJ���k��Y�J>��T��S� R��J�@�N�d�10tҼ;�b���xFH褅�w�Ed�����QD[��jCh��$��}c�Eck)R��G%��d�j�h>��B����-���eԭ��ܽ��6��a� ���,'`ee�Љ�h�{�-�!�K?��Jl�(�T��6ڱN�`MUe��Xl b�T�E��]�yp�z&[��3YRm��#A���Ǥ�Y���6�r��U�􌷛�GvP�	���cj��q��FV���;�w��Zj��\�C�9H��:�n�H�ɘ����b�`)�3^�43f�ІM!sd�I���"q��^���@������-M�p��T��\�f��I[��{�
�H`�h�5wne��,�7�$�Y7��a��l��k�K�� �9��%�j�c0�ǒ	�*�Z�jT����n�u��&c͔�6f��EL�aض��m�8JG[*T��u#Z%�̡Xv��WD̛���K�t��Z�ly�bK��u�W�TI�J`B���A\�କ�u�G/f��#����:Dn,�WYC1���嘕f�E�yt�R;H�n��U��c�^�������^��n�Á�吂���p��I�X�p,�w���&kK�BT���÷i�ţ5�p[���91�C(�Y�(۫���������xVn�ӓ&��p]-�H4f��q�J��i:�-	��:�^n�f�����VPZ��)�!��M^[�x��[*i��^J�+��lkp-�*�֡l��'Ew��O�e�ԡKr�2 P�Q1F�9/D�c+2S�݅ ̡,��L��c �q2,*,!�q���7��f�mG�emmn�!	���B��f!�P���Ѐ�	�@*cwD�qa��x !�2����HI���wt��y�J�LRydm㊯[w�f�R�T6�e(]F�ʚ�� z]cdҳb@�.:i�4b���Z5��mB*�WBQҬ(�Vf"N�I-Q����=9Gnn��ach��jn�`{,l2c�)����*�Z�HB���Ar�)����|�HU͊8( N �m��˭Y������u�j":�	�M�]i,0d×n�ּI^�Ɇ���l�ĭ�3H��|̊�塧D��lX�jZ�+"��Դ0Fa�� eґ^(��e];��hE�f
҆<�T�B���x��2j�+r��kF�eK
X87J#/t)���ˇK�4K3I%�J&�I3\���L憓7���;!�m���P[�G�9B�HB�M��g(`�7h�Ln��w^�[������)M�r�f�@t2��g_�w���]�5�-���O �<A�V�Aܲۡ� �E�+.��Ԋ��<�vSDH��F6B�Š��=�܂*�ߦf팖/��[���To�봯���n�:"⥸^∀n�[�N��aF��[�G��=cj�ةIy�Q�aצ�&]�E�ZcOi&]ۑn���/4�t��\��w���V¸8 ���|��Ud݌F^
qj�2��3QU���<�2�r"��(�e���d��G�-����"� 5z��1��6�P����{���Yn��U��N�Y�G��@������
����-+ G^S8kE���,X�#6�ˢ덻u�M�M�1�IR!�Z�|\Ư�5��;�4.�#�e��R�m+�<��Mvj	��:��w
و�+q�������f�˧��˧59@p  �i)^�E��3�g��֛-��@����1��hX�nQb���Ͳ)���8�QX�� ���E��.�<��[`'�/ {5��������˛��FͺL/�7�	��Y
�������d��Z�f�b�m=K
�YN-�x�^��e^�h�O��7v��J	�`D$�F�� 3W�[�Zka��&�p��{M����M����u���4
T�J�#�,*0T�"���Յxd׶)�@���扙��o+S���Q��Y����S�#�7M���+)a���:��F����j��U�+!ɇ��3�F�^����U�����&���@�%.�2%�ilx��ḽ���oS,^�u.�,M�@�������uⒷVcyp�+�TR�-wXv���M���m��k#1,5��`n�r�%��%N�B�ѫ�DۇVhŨk��)�;���v�ʄ)��T��7h��m3�Tb���sE��6հ)+w��;��X
Jh�����U��7r�r�젎��X6�1�`2�ͥ�t'=y�Š$4T{i����t�qJ�6r�v����#aC6�j�w	�&�;��A0캽˺U/v�z�L�	��hl��n�SFܐ��Ú3m����ʲwVH������e�I�'�by�d4��3\�qSxH��n�Gl��M�\V��37`�`���Lu1Z����
�n�קv��r�ʚ����]:0Q&��\����3u�y.l�+uY��m��ڍ h��W�V��!��p���悪C׵r����_.C2I+�v[!<���s�--�[tT|��`��j���-�t�.�茌�❺�u�̩�2��M��+k4Ry��M�f��Lͤf�z�p+��בbv�F�l��*�DzQ��AE�%W�3M+1[�}�H�*B��l�2fL��������B��T.�H���&�`��U�;�ݭ��4]aZИ�'�\c6P�cqowr=)�J�,��
�[*�,6(�<�uq Z��qiI$ީ�D�@TU/$7Dhh6�2ޜ)b��n"C�w`f��*����&ZH�׈6��F���Kf��F�L�E�'Y�0KqL�wU215T�[��7݋��J�8͌�{xSͺ\� K[�FL�Y1�l��1�6L���(���������eh0��ڬq1Xh3B�ei�٪FTA-�1[�.��+4\3���Þ��X�Ҷ��G��x���O��I��z]�u�6�V���F§jfK�=�eV0��1fF�ս�D�2nS�R�h;ZJ��q��"�b&(�����im�UG4��f�fP.տ��«Iժ����؃�'�1R&R\Ub�#Y�61�3q�\��ؒԒ�7��;�Q�.�{S:��n�4����p�37d�X�8"����-�-0%G���v��.�k��;Y���E �ל,��5z?AQ��ei9�+ׄ��Z��Ӫd:ܴ�o@ݕ�j�G^�s��qj+58
i��ڷ�=��R��U��Zwg�t��n�8�+�dT>��^m�Rzr=@7V�\�I�wc�!�F�7�IG�/3&] i^լ*�I�L�]��݇j$*<ݟbͺn;��O�f�<�;Vr�{�6ö��V������Yy���{�ͧ���˺}th8-^��Q�n�wy{1"�b����$v�ڐ�un�Ei/��d�uckt�J[rV�P1]AKT�X������=Z3Rx
�_e��.�_��4l�a�R�Q�{Ru{�N��q!��Cu�^<U�4�P�iѭd���*� �#sY��[��Y�oj�i���X*aOa��u)�f�����C����0�
Y2e�ܗ�(�Gw�7�kFi�i�m��ٳ�X��zdT�@�/��wfY@�����s~�,l��A� ��7]�@��v1�`SVa�p�ٰ�PH`�4�`�-���U,@ͪ���U(7J��YF�43�tw�4r��sh�wWi���Z��5�fi���V�>o ���M��Ŗ-� J�Z�rXE!�����]�L�͛C*�����N�x��f^�����l�wL!���6#�$�#e���HJ��^��V�J4�:�q�[�oF	 �5lMȨ�7�5J�MKcdǂ�xu�lB;ۙ�l����e���yE�i+B�6�V�;�2�������$��7"t�e��f�n���8�)�Oػ��y��E�V��k@X)ۣ[(�]���6�h�!d8��m��Q&'p�ωܥ#n�G�L<�@�&UƓ�n#a���r(���9�˷]]�ms���t��*0wn�כf��Hh�VdT�m��J"�rMۂ�T5�u�^�`�2�3PQ`�>'�k�Je�%�G���k��%4�$VP�f�߄������1��p`�:4na�S��RZl���`�*!+qV��o2L�v�n�c�&�,�;�"�osp[Ϡ�W+!ê�e��U��R��70٥�4
�F�a��cر`�nbA���-]�G@�F�o��3�G@� �lЬ�4ʴ���6�PZ�y�1VR�lCV�i�A�3
tk �jIK͵�\�:�Y�u�W��CZ���Ȗ*V�TŘpQ%K�u�D	A+�T��f�8!��t�L��5e&jT��nޜae�d �sԲ�n��%#�����4�����s�lo<���uZ�yu�m��V���B��3a����ؚ��A9k0�O�
4�.�]J�=V���|9Tͥ$��ʖ�Cc��f�l�mZ1f�GPGEc����4	��̼�G��߱(��^���5Чy4j�!?�Xu��[Y��kܐRI.֔�Qۣ��h�5h�bصP�Z]�q_��0?d�H
�0J�4R�O����jL#�y�)�Rڈ�b{�ɦ2�	G���4L9���$�e`���i")����ܩ���ff:�-��-1�ayDʓ%dc2��W�=8S���J��J(d��QH���[+La��Ln�m�Vkr�W�k�ct�lt&��`�$(aű^��m�Ǹ�g1=�3-�oOي�E2M=s%�մ�GVj��Q�Nؤ��ޢuf�O��O ���(� �t��U�&��˴6�	)&婂f���bUʈ��E�X�F	�lBP�3�N�@��i5��zB�qRU����v�if��,����:L�=ZE��)
6�;����5���Y�_k9�o��-��+SX�/零�S(,�v�m�ã)nр�(���]k ;vPۖ��F2��kXA�2%|(3�:������B����+qcq��f�7M���P*�+L���`���^�Ŕ0�R:T`� na�we�)�[b`�☣.�:�T�p�³�Uؕ��cf�C�o�G&F7"BZ�0���f@EDC�f����-ܙ��%�WY��4�k�N�M��j[��v� �t��=����M���Y�����L����5�SF݇b���Unǡ!�m6�'*%������<���6��2�T4&� ܖ��6�L	��c���TU���VD��)Xwt�JR�Y&���2$�uv�f���U� ���%��eX5���9MKO�F	��4)�&$eҲc{���QI��:�D�+5
�7�Q���%m��r��t�$b�nL�m�N��i��skxJ�9%���"m��y+0K��2俲R[!�%i9T��ye���K�'0Ho,dZm;#1�R<��	`vu����wu#՘�o#C*h�6������e�PLD��c�o �\������T��V�Ǵ&�r�*�V*�[��h˩�����L��0�!���r�a=�@"�Zm��l�s!-E�����Y��cJ��W)�>�i�-� 5-�(��Xy�c�h�5Ef�PZ�P���ɶe��{L��M�V��341>�sK��*�͘��x��oYFf�,ْ�Ѷ�Gw�3d�s���O
�5��ݝ�@�yg������W�y�t�yUû�ә5�uM��'y�_9G�k�1`e� ��V�T�ONFֆ���8������D���� Z�V���J�<+"º�K���tDn���Z��j�s*
�d�)ٚg�mWt�b`s'n�B�P�qGf6�	�)�8兙Gb����EՕ;��o9�G:&�̀xGK6�ՕO�T�]6�"Ά�Λh�X\H�t̵�Q�"��StۂN�����l��[Wr5/rYF�+���GD\ԁ7��y�y{�9׿T��}}��?v��� &mh�����y�u��N��lr2�1�7	����Ǧb�VNY����;�Ӵl�mn����N���E�w�R���,/KŔ����we�%�'éSͽ�]��̣ 6�w�^�N`�����~ޫ�)*��7�RA���r������Ƚ�ڙz�@����3W�~���l�@v�W��Ǎ1�;W*^.�[V�%b���R�f-�$�̈*^v���8wq������F���9�b�T�{��U:p�;��m���t{q���Z�1���Q���P��1�#aF��v��oi��9��և�ìǅ���.�f�ݞ�i��P���aV���-��eN���J]�5ߙƞi�� v��1��A�\��`$��P�1����̀���u�Uy��¨Zsdڹ:�	��UG�Τ����[0���3�Z�*��T��jZ"����p���Q�;KEku�"�ʁ�v÷��Wo`��ö��5*.|��\q�fa4�̱K~h�����=j���u�;�eϹ���7��R��LX;:*s&�a�syu�L'�>��s�%��e�h�}p��fA�x������`��Y�C6M�-��>�,�s��\SNX�a�u��.�u֪HJOn�FfP9XLV:TM@�r4�v�ބ��s�1�ۖ��ѭ�Ig9%j5��UR��󋲴�t�
�����g+˷7EQ}Ըl���/�M0�l#�XSH��������ˮ/n�m?/E=�ق]��cv)���;/��hY�������֡��
δ���\�WnM8���,i��%�\��6q�yaE���gYE���h[v�-[xɺ�u�w4[gD7�s�)b5j*g)�Yg��^�z�շ�a��µ�vlLo@��b�oH����hWJ�l[v�<QU*c�\�%�y͓����/G7 ��NF>���I��������}�BZ�u�DIQ�r��T�eQ�J��U 4Qg�څ�3�9t�W]�(݉@��n�Zr�����ٯfR�9�����ё�N w�anh�1Q�ؓ�ϼk��z� �L�Τ[�E�eC�,q䕹Wx�� u�_B�]L;��uD��0o�S mv��H���꽙7\w.Vf��w��&QN��� �*�l�aR��5�7�v& fp�6�ABm����a���6�^ۙ[:u�9��0�b��y��]J���nM�ͨ�frU������!�a��I��a�wrr�g69|�Y/@1� r�0�j۠�r#DJR+`��Q�):T���K�X�]ܭ�nV����!&�}�x���*n�J�r���·��J݁�q����Ц�`����t�ޚ���t� �$ǝ��ǵo2h˫����j�[��k-�۫��.��[{wq�+�=8��9�p{�wN��ɗ*7,b�� �QV�ޮG��/�l%R�$M
���T�����$&b4Dښ�i�_S�{�7vn��)q������*�O������+���u:w/7��T��������ݭ��C��}��3z���sP��:�k'fw϶�\��a��I(��5d��d��6�q�ٻ��H㑹�.����9�u�Qy)+yv�nTc�-������㖂+��3�4"]�Y:}�F:��M!��*�]w&�76��mX}yg�Pq�s�x�%���jݮ�ܹ��ɇ0����:�m,S�L{x!/�1����s�!vz�yԤ�-���i	�sO�5b�U��u�E�3Wb�%���̲�/z���`N/��O�����St_)w���Z��`0mpԖ�5��sF%�Wi��7z$狒�kVV�l�uWmY��Ա"��!��
:�AԚ�Ծ��]�}n�*خ o;��1$$�n���^m���5�2�
ɜ�mlذ,�J^rJW(�Bη��Ќ��)f�Yd��\�7����K\9m˳x�B���F�x�޾��( b}'v,����c�	#���51�v2RW+�w�4��2[[ӸvWk��H]���&g_t�X��L�[�b*d�9�f]�7�6�.�8�\�#�:̦�zb�p��)o����}ʓ�d��V6�r繃�<\vof�S+�T����ƐE��d�c�g:{�ۈݶ��m��5�P�#ż�-LU�ܛ��F������|�B4}��R�L���E�����@r�L�5��w��9RqfY�7e^���bڃ]`Q��C��� w���T��^�SGE��ū�0s�r����7���,.��K�y,���8��E���ڷj-ɸ�E��ٗWu����d}]�ڱi!Fd�P��C���T^қ������k$����#�m]쫛������N�a_o-�w�J�\d�7��ոSo)��U��A�o�WX�J���"F;k#QRʝY��6�+WwI�)F~��]����i�A�w���$����\��.f�K�Y��������]�����Q9p�7e���n3M^M�[��v��G2�<�[�#�6kt�Y�q�tn����9�Lo�LT]�p��;tG�i.����&���OYri������y7�Wm��)�[�Lg�J�+c�k/��<����%��髝��#��5umN��?YO���;c�SZѕ��6�Za�gk���wV�o#ǽ���s	/Mc�Z)��p�Yv��:�@^d�-.��+���ٮ����f�J�}����	��2H�[�˓vHX�m^˽B�`fK�}n��>�s�� ��ܦ���;�utr�s��X���7f�����D�^�3)S���_e�����I�4a�c0V����(-�ʲ���/�<x"2�M���o;vtZw���r�"ō�KǓ��yʀ�P��O.2f1���%�*\�0����J!h��O�N��"�8���Yx�v]X�X���Q%D�s��z��W���F@P!�Ȼ9wgTX���������S��X�D=�uc(���j�ht��t�Jt��Z��2���w)m���EtH��b�֛B����M��ఔ�k6ԋ��i�+zcRj�ެ�`q�p����]���F��V֪Y�;7vo���F���$;I�Z�^o�n����G쓽n�[�-R�ڬҤ��#o���g���E�9-�4bq�tn�$a,��LjAjG��!�\��X�ݷ���jJ�ʙ���@�����˺6�u>�_�Þ��&O�X�Z������7��x.Ti�6�J.��s
R�fVe lV���Ͱ�㾱-o���v�,��zZ%�:Z���} �n��Ȉ���̋�pn#�@.Kn�5A����0��Qqy�)N�ڝ��<ônA+P��a<}+�J@T�%���x!b�T��}�x���q�]l�٨J��&/î"& ��$5�G��<��V�$�{Vk(�ʂ�-%ϑ]u�����(�7�֨8�Jg\�Q����T�h�8|�\"��n�߱���0�[:���X��h�\��3Nma6tr���*�8r�Wz#-�C,��(J#`R�r(�,UҬ�Q��]�s�PY��;�xL;��3P׳����q��q�<�aia���U�@"�L�x�7R�(�+4-���RT{����v����C�Á�,��*ѫ��a�w�&c�*�[���6���pt{��!>� ̉.�m�ƙk-�4�N=�+SJm(dC�o�����uCNun����wWK���}2�^jhv��d��4}��Բ�W97b��#m�Lp��*�V�	ќ��%F:�.�	);��
<��z�k\�nb��Jl�&� �� �D)XY����Z�#�3>7X��e�B,��|lr|ă_
.}�Ή�6��3i7V�en9����yg�w�I]m��ߜU.���-���t���S��A�(Ev4��p��a�$��vP�uӦ�ͼ�ʲ�o��c����>�y��Q�<��ϱ�>�7]O%/��!��FJ�(2���ӆX}��-k���}��uY�vk�\4��;8m>�KQxr1+ �n���nCY|7���,Y.�� �se:�����n���f�Q*���@���Cw��
�J$vr��[p�rf�N�}a�:�$�
�L�n�$ZQ��] �{���+z�� 1�.��R;�������cV�rڗ����3r�2�*9��ʚ[�.���ǂ�,:� V�r�7���� �A��J�#���v�1+�;��t�G�	t����D,���N6a�^�4=� �o[�0e��v�n�t$;�.����`�f]��I�Z0�]ؓӯ�7�"�t��|d�R�qv��[66Vd�yt�GK����
����ͬ�bGu`���}Q�XѢ�ث�fn�|4��"!��,�ͳ:���g�I!l(8b���4m7�띸,Z9��~��h�Xٽ���v�m�ۃ)�&o�t-�)���o��4S/�ɘ�g}�5�3#�9��sEu�go[.�_��ci��pV8pS�+j,�&V��7���euN���Τ��M͠ZO Ka�#�li�hΗ��vXE��6^dK�{W��{wآG��SПpSu��Br��.i�[φ^(ig4%�٭���n���Lc3�Y��\�n�[�'}��{������+�BfG����We���]"�ݜe����X��PH�ls��������6u�Y�^��O�&Ï��m�f(�n��J��ф;D6=<ۂU�ޒ�V�}g�3u��nY��ZZC�ʕ�-<�6gwP��:��8����z�H���h�%��3CN�� �[�룖?$�Ǟc�JQ%%�s�#+et]Ͼj}��5$��c���.9n�u��0;G��ɔ��|����b[^�&�Sko�)d)Xd�"q����,�d�$��-��w�\,-��7�CK�{>�ŌW��bY�r.���-�Lvc�ړ �}]��,J�S�ꘆ��r��M�8�&�Ap���WK�0m��{���Yv���4mt�o�F䒔���R�EK���o0�*���s�*ax�Ϫ�5�p���wx�<�J�Q���n"��K�P'ΏW4�p�;Wb��ckH�H7r�,����G/���<�m*yIX�d��}3@;���i�6���2gP�V�����fT��Zʶ0S��9ʹd:�0��P��YQY�{;#�k��0��^�uQmH�gIwY%%t��(*�1��A-V���jl�hopw�ŻI�'T����.r������;SYk�C7mī��8���V�Or]rf�Ѯ�<x<�;�`�w�a�gV����L������t��&�/ �j���p��wVH�q�5 ��u����Gr�:�MuǷ$P
��sHK�/q�{��$d�Tx1�[,V��%��"[�99��b�B��a�^-vc���A�;-Z�S��E���Y��;N��*C�{�jKھ⅐�-wS]�����W\��VF/�br�o��6�\K�<8��վ���U�5�8�BV����'a����m�?�Ytԥ���?>���KoKS�����l�һs�M�eYH��M�n� x�_f�6�p,���Y��:�2�#�d�W�Vf8���3:_V�y���{�F�ș�8�o������?�75[�H���T˰��h[+UA��x�'"}��p�CX�"t�����x�)uq{z��Z<���v���͉����+�=ɤ�I�XX׼9gu�J�9���+k�����u����6�"��N��^����I�w	��kg9
{��`�W�)B���y]@j�H��yNh�G��&F�v�M�Gơ��F�>��iN�6����+��&t��+餫zh����+rv3v��L↟١v_��zWN�S�KNgϞK3��p�vwGy^f��%��KTt�va�����3�����;N=z��b�N9�]hW�Sw5���jFxpO7pML��WY��n6`���"V�j�m���m�F�b]Z��3��e��\G�,����(��Xv���ƶN�Σslu�&!��@�B��4	}�t�+(_n�XR�ۑ]1����J_i��G5�(b�g �.��xԈ����� rU��x;�e������<z]8���R�Ef��0�j��Vd�5�A@d46;4`|i�Wh�)Ц������ � fl
j�t�s6�b��=�V�aU�c�.�n�@�\�4zk��E�3�	pW̳����j�@��ii������[�j^1N�]q�tȬcN�L�-�����{�҄1#��B���Tܬ��ݼTF����;w��6�#[f����e��^�1:��)Ԇ�����}��`�.�����o��>l��6�6�R�dv*�.�-��-�ci�;��w��G�r䣧B�e��}VMq�n����]хl�k�zC�l�+���:�R,q�f+�iZ�|D+��!����S6��c��w;���;-�Vcd�,Tw�՘51W6��#��W���|;��!��'��rxCɁZ��S`����GS^�YS����^J��fչ4V�f��Y�m+�K��
�K;x6V�ʜ��7l���{�(����ƫve
�6��8���u#���3V�W�8Y��c
�n�t�0Ԯ��E3�Q���'$�+'ZQA��u�%qi]M��rI$Mɂu#q��x��N!�ӵmIX%bu��u�����M��LmgM��Pe�$���kR���H�Ԃ$�L���� GmG�y���2�:�Ud�,
D#vn����A$��'AQ��mNn�#k�ƀ�(�-�E(�ƈ�`��蒱;�2�]��!x2��."�Q_���%�N�e�e *�q�K���Y) �,;]��
�B&+E���N�5��!!	P�#���R*(������ A�������)���z�{����O����}�P️��~1��7��ʺ��U3$�<x�bZXz��/F��'6�+`�ِ��q5��vI{:CvWCNt��h�
�;�����ה8ه��q��L��l�j�4��G�s�����j�{+"V�lյ�+{Ze���+\�8g.5��ԋyon+C������)PH"ǲ[�̬Hu��Ւ�o]���&�$������*p`�%�g))V*߳RFh�p�͜F��RT��a͋�k!5�Zx)虭(7�*���l�E�\�f�:N;�``U�u7�a�Ύ�kw�3[�2��7����˓�\$ǥ]�[n��[V�P$F�慃�����B(^�;�%u�]NMm;�b����LOdڥ�Z}�wD�\jfu���d�0����Ȧe>��9jk��`��Yw��B� q�E��+�b�+�m|�f�rGJ��!��Օ}U8٥+���s�\�I'Qܾw�e��\��!���
dΕɀ�ֵ�33\oy�����R���1cQ+���;�V5���y�.��ǫ���j)0���qS��U�Y�NVV
�H�C7*�Pb^E���A��V��]C�j#bҫy�fk����j�����0��[�L�K��E/���Y�}���c�pf9	GL��\˔�h`ĳj��c
ݗH��i�wN���;�L�� ��)  ���>�k@F�ҟ^]ʐ�X�u�A���,�_�y3�83��<�P-���p`��z�0�Ù%�X5�n�y�ˌZ2YP`\mǰKnjCd��Ge+�:oE�J��T�q�"�����R����Z�ڵT��䚃�k�u����y����v���huvz�5S&[~2�m���Eձ�Ƶ��4��m+���a���7cZW1uu��v��ڙ\r��u5.�uިZ.�` 5��g�R�2�F�hEG7���tN�vcE�v�7T��6p��kDf�Ry�xu4o��@�V�Z��*��{�}.�$<90n�u��|/.�=���=��&��8�,�j�����3E�4�Δ�c�mf����U��C�"�CD��S�
�,ç6�����X�)�r�*��C�+��&�z�:���u0�S�hYv�gq�n��1H�[���C~5�*l�/���EɪV�}̊�'&��F�� ��gyE����I�F��$�� "�w�p�ۄe�	Ρ��|Ďc��禃��#��#z�f��λkVk�����Ūns�ϧ+�@�X�����G�᷀8�e�2����0�7p����sh5l*��䴗�X�I,�ҫn�I{�7h&F�	ԶL���&��*+���˱ ]V��:ė��S8��(�� q�&2;��\3�I]d�|�ct��HU�d�DN�^3d�3/��ަr8�%�Z�Q9}-\Ȥ�jt;[Z)>m�>�E%j�(to�;	�� ��{X��R�V�����2�^"�R�� 0y��q�q��͚���
���Tk���yf�T�k�����yQ��%-�
`S/�즄v�|�^���¢.M�4,j�/8*�>%f])�s�nV��EM��Td�������&ƤF_F'
1\g ����\���mA����WU�U ��>�p��ݚ�#%V�<0��a���֞�e�J�<�/;�b���%��J���αt�\U8ۆtT.+Z:\�辷%���c�Y�^�6t�N�R�����SL�	c�9����.��뷍��1`O-�"�n�NG5��t�j�ݩtt�-��F3nm���J�;)�X�g�/A��K	�ܨ�Rna�{y�m��� ��fM[*HK��Un����"�t`&Q�v�U���c���>+v���'D�ӽcH�q�0�Z��b9�u �A� ���[hV���*�����x�5y�:�aaD��u`|�g���_\|��\�ܺ��
	�#��˻f��i�ͩ'��@�g=8���ղK�#�r���k��J'8蝪��9/k%^�%k�;rȆm��1f�͛�}�&�Q�dJ���c���Pm\�ζ��v[�m�ړ�|�i��*4���<�U���@�9�Y�>�U��]C�e�[�98�gIX˛�J�ͫ�Y���_k��qK�
�l���P��*aF��Y����Z�uvS)"��֎!�K�������-a����Kz�h}|��@�,"��=��eEk���Ý��cǼ��k�߸pm�[����]�9�o�9Ǒ.V�� ���gnL�H���v_&���T��'2��293邀-�{+e@�go�i畵/vY��	Ѯ��&h��r�|%�ʯ9�5�'%�H���2в�?̎��q���(��$�g>BލXz�U��+2DM�2�/Y4:�t��B>TZU1lH�2Z�b��\-L��w�yEdt�M�������n�jf`N��7�œ+�os�S�k�{f��������ʽ��;r�rw����͙�IQD,�(�w.�w���D���n��ba���d$R7�ew��g!R������5��t��tNtd՜����w5�:vس��&�����9���T��<��V	��+�'`�:n�II�II[.�Kz��*���C�)�"3����&�ĝ�T�E���2�܉�\�:����3G]��ꈡA����1�Z]s�|��`ߕu���%;u�.�0�X!���,=�kCm���ܺT�"V��zQz�D�,�.�S������Mjx���;IA,�z��ܢz��W�T���WYye;�Z�9G������� i�,^!�H:����VEJT���
 �P\�p�J ��m�.��ِ���s����w"k.���ky�4Ccy�v���P��1�Ij�R�{��=�{:��3k���} �
DI�)r�M��b�^]��\累��]@<̎��m�G��Z����#�ݲu��#R��k���Z�[k*<��ݍ�*���CE,�� [H�<�j��ɜ]Y�t<{�S�`C�+��t1�dY�#�&o,Z���jL�N����M�\�|hYs�i�O6�v"��+%��{7xUA �fZ����F�j侨F��HIsh�6Q�3�Jܬ�-�
�8���.4���<������ʘ
��vmA�۩��_T�IY�vɳ,q��� �W!�+��#�3%a�/pT����N�����ؘA�������h
`H�	�5ۙW� ���W�u}}e�Ub[�ꫩڈ�XXI}#���XڱY�/��[g�NJwl�L$���w�����t-��v�u�1�m�x�I�rHF^Q_+�ך���L ���YY���i����#M�it���Mw����}N��Ň՛�Q}BNyPU� �¾�7fWN�m��\���AQ
����9�i�i��SI�{��ˤ�\(Cs���5l��El�F�����={)ƺLβv�j��T�z�^���,�I��ܢ�$̲FԚ��(VA�H��XNm��ʼ�5�)U]#Tw�T)��KŝjT�]��ȼT��U��Qh-��N��!��,�Ab��pU��%�xkwZ���6��R�'��`�`+��8=�c��x��NJIX͟<y�9E�y�q]tq׆9�c�z�Ɏ������ĕ��T9c��]��ۏ.�����:�e�=��$�q�,���*W}WWE	[P��9�z;4��@n��v��sc_Wp���]
�\c�zd��s����-^��ڼSu��S�5�D�kͦ�}�8�ӕ��<]��|G[d[6�ssܳ2���u[�\];���T����F|˘�/��Vy���fi�!�ڨ�i֡�\��3��d:1H��ʹ����G(���6x5�I�
�|�U���=�����sc���\<ú����A�ǪN�9�n���\��:��3�	��7kI�+����{�>{��ʗ��7W�:G�Z�zX'�S�x����ޭu1e��+����uxlѸc�������u��vV̒N�E.�t$_�m�0��Wj�\��ۼ�|R�-;�ӧ+���	˵Р_	Zn��(�i��gU�Ɛ-��I��ٚ�7ާ�Y�3�Ωi$M�<ط��v�m��h��7���(�T���ÖS�+-cD��}6{CHc�۱f�4���4�ާV�K&��V��D5�@�+���5_Wճ��+)�{�J)�����tu�vX���H�^A!�k�$UoI�'����uPi�K]bc��eY˕f.���i��k�T<N_:Eؘn ���E�6�㝼6+��M�>)�B������N�wX� ��A��V��)�g^��;,���w�m���^:î�:�K�Y8�*�5��Q�M����pʸ{f'Rh��1���`=p-hJ��-�W:���>�ppu{5�B-VU�PcG�w�!�I�պ^"֖����Tpq���i�.rF�nj]��
K�l����5U���s&�k��&��y��Vȵ� #դ�u�����P[�	; ��^������t!p̺wh�04U��j%��0��*ȧ]i��o43�A��\����a��o�T'�j^���W��4��a��6��8�F7@[�]���}��9uT&�θ��q�@��[>W���Au��q}�őY��Ã:�C�0�R��̛�u@ـ����x{������<4�����lKi�Ufu� m�,ڞt�=:�(A֩e�C9d; 5�2Ҁ��c\��T¨�}tg*Өv�MU8`Y�KZw	���#2�@)P�����"[��H�5�r���#9_��݄�u��2���w�$���%Y��4j "b��K�&S5�E=v+5�3f\���ZƵ ͱ��p/8�<����َ�r���\	umGy;VVJ�!N���S/,E��fA�T4�t�k�t� =�L�,�N��b�gC<�����lk_���d.��R��q�:�!�i���S��ɯtq���TG	����4k�X`��R�Z�蠦�eK��&j��}3�尷�v�k,a�Щ�Zy���w���k�0�1�Z�J��m���˲�t��d��zrKu�I:l��6��(��W� �����E��A��J�1Q�����y)U��Kc(�F�+��kݣv�f3 ��?a���(�r,L<�Ջs�Vw4�����p5z3C3AH��u�[��VWe�y�0P���Ѻw�����#m���J����f����oP픞 ,�R�<�8Om��@�� H@-����v)й����1����}v�v��b��w5Q�/㵇7J:�muv[**��:�J�Y����&��؍K�V�+%�A�@��ܝR�p�y{K�^�'��n���.{'�hu�T�)V���U�:;6^�N�J��������e���"�7���#:4%.�A�G�-�z_mt{|�n��{a���Ntt�7�47�`���(�M������ՐAO+%t|��M�'�B��$��r�-q[�J�՘��Ή��ԾU�+��ʁ�Vdӡ��îێ��`d�Ƈ8`���:�5��t�pl.-��O�'S�K�lxt9���FSCb���z8�Z�b�ͫm�V��a��C�v���T��7E�t�o`�Y�) ��ʷNք|;u쥆:lL�צI�qVh�8��F_����n.X�������Ic�i��Rzy]�����j��K���t��]�x���5M4~;zV����,iN��(�KE+�ه�w���q���m=B�bq6���� �pީ�����6k�'��.�o�5��5r�g]�+w�I>Ѯ��瘸���5#6�U�Wn%{qν�ܛS7+8-u�D@\Cna�(m.��0'���ցQ[�ʧ�+�Oo+�8}��B�.{=J1A�HJ3/�m���(R��!�Z%ԃ����gZ�l�c(�'��|���Dw1(cJ'��ȹ�4viX&`#��S[@@Ә�S����і��0 �G&T��h%������Չ�'�p�g��7���r���uf�Cp��Z�/��0j������C\�����'9�B,?�)�K��З/�mT����%n�)S��iK��WCn�v��X�#�iۭ&��";�%bKC&ʢ�[��j�S��5�i�iᬰ����b��w, o6��WD�}VJ���c�jt[qn��B#"�Wn�]�m3�w#�Jw����f�Ӱ^\�{ʭ|ى<�(i�9 %��]�0�����o����r��Hc.��l	Y!�l˔���U֢��Í�Qq9qY2u*��%���.���)�S���
ӭn���M|�cَiח������W0�B��5�*��~/�auڭ���̎ׁ�|,+�MPX ���x	{�� j�j��H+1Էt�ʛ���T]�*��X{\+�cV��$�{8Y�yQm�Ԍ�[u�[Vwc뿉�ǵ��S�A)]��7��+�:�ϴb��v�8-�r!��$�mq=�O�G��ħ.'n>��@���k&HT�❋nd"#`s�Dww�c[5	�V2�[�ʼy)�X�!���������f�ԕ�/�^[�Af��Bd7���sS���e�"��'A��oE�`�(ޣnN�,�;B���l
wP�Z.��m`�1�]��3%r��%�
�tI�*��_k3w8ր%:F?��4f���i��us��:P�Q�b��\uo_J�3%AvP;�J}3^өa(b��1`6UΫ
�<�Y1tJ�w�f��0WG#i�)q�{���`�躻QѦ�q�JŘ;���[:P���]^h��U�/{�h���e3�,\��L&���:�)�	üG�|��_����� 
��O����O��������?�������o��~?������߻����i_��l{~�(4�Ĥ!,����!��������������E,�a`�yR�D�]��Ix���)�Y �\^�!@��/)����C�iN蜦��S{�뫢F�2���3b��gWnf�BKH�8�\�l<.��u2�ܗ��m5�r��Ъ�T��/Ft�[���@
�o��Zt�^��˭�x��ED#�v�B7'M��g�C�,�j_`���Tum���e&r�]0݀k���3rt��ض��rg�uG�DE���Uh�C1��r��U�bo6@�f)]#+����ݔ�w�SRăY�-*yOEi��җ��A[q�@�������Y�����d�e�j���&��%\����κ{�:�\��9�޴
IǩwN{��umʗ{��g+or��(�B��Xy�>�VT�������#�n	J��._�Q+��v�՚�]��Y0bˌ��-3�n�SDq7�&��{��j���cY�H�m vȾh����.�$ud޷�{�l��Փ��yX X�QGb��༾�.8{�%�:w�nbOK�:U��q���z9��/(��x*U*t��,/�9�t��\x�,J�b�\F�]P���!WV2��9�:�q��2�#�_2$y���q���d��+��,��Ch�b6���^Kê9���]ovՓF�S�t`�!X�ut��ѤU��|Έ�gv5Cۣ�Fg�ݞ��;�wb�m�Ί�xب*��Ӣ2�*jz;��h��G�h�gk'wv�T�<�(*ւ*���EM��*�o;�����m�"M�DM]�1WF�**7���,GZ*4n��5L���������h`��b��#��-�g���DkETS�雱��כS%�A>v<�UQFӳ�lDDEMEvėcv1�;)����QP�m�*1�N�A��ƻ����E1mN"*���f#�Gh��wtUDV�SUTI��؜U5D�Pn�ɺ��V��v�6��uUǘ�b��E^l]b��;�WZ���v�5'Gˣ�U�m�Z�cy�1�MPA�,m��b���ۣ��(�)�Żj����0S�4���y|�7`�WZݹ�Q5�"����A�ږ)���6�w��"�ۧ�K�m:|��E[b&���lDQQ&ڼ��w�����ww����O\v]���ۻ�OU���Ƣ(v�3E]j����^ �B}c��Ad�V�.�UE.G�s��)�ܲ�"�Fh�X�Ds�WF�:��{��	���+ܭ�?�ًZ�t�$�O�>�Ȋ	3�M�29ӈ���\~��T|-����S���j���"�v1����h��N�s��{�������z k���������R�&};���S��J�粻&|�{�z������y��&W��5.3�{|)w�^a#W��^�5]+�R�i��g�����{�R��ʭ�|;y'���+}������%s9܇��:���_��ma�O��N����X�O�G����^��q��Q�ڎ����Ԇ{�L9m|pfE�uT��n�ܦ'���I�Ld�����B�5���0N�AY��ȶ�]���F�%��L�R�I�O)�����{K{^6�;�|�� ��3��Γ�a�D;�mLd�����'t����b滌�4w�P;W#dߨ�=Ә�Չ��߽�{����U�>�J�C �ST1Y��� ��2$ma+.�_ �Vp��sZ���=�ԋ/e��O{�F����*�����/ݽ����P�G�UY�䫣.́Ĵ�	��������ċ���[6R�uw�Z�5ԾjY�v���h��zB]}��]N����"��(���%p�9%��?`T�^���D��km��9L��Y�~�H�k>���1Frhw�!�y<���B����62n�9%�m5"t�ں
�A�rj�j�/������R1n��(��9�ۋ2�Nޭ��{�+�~�Rg�6��قC%�g���53G�<��8;�[�{�m�g�ޥ;��;��>3Ƥ,�'/OOS�������N�
��2dd��K�y�z�[���t�����=5{2�>�쒵{�go��N�F�������w/���oU	^�_��q8��:��{d�K�N��}��>�&Jà�����Ȍ�7�����I8(��oe���^}~��#�=F�M�'z���,�x�O%���Mچ��5Y=k�m����;n�&����r�ʻ��ϟ�S�z��j��,T�ۗZk��o�B5�@Z� X�o�]Э۾��ؽ�yd��pj:�/��vա��F�fMʽ"n��ƻ�L�}�v6�@�L��;n��+�V\�@�������`�6u)��Vvvc.��0��19C�^\�дVR ԀT]8���#9X���=��ۧ~��n���.۞�<����+{�����6ظ�n�㓬o����3�67�=�����?c�f�&�s�کg�ϫ�'خ��Ϯ��v��FZ�X��p��/|ۡ�	ŏ�:L�|=��)��c�
>���Z���7���^_�u�ς�3C� �ļ��G���vV�kӃ��C��]�<�z�����}O��u�S����tJ��f�tY�I(m���k|���y��zk�D7���C����ךE ����t��fۜ�w�)Fx}��o�y����돮d�pո-K>��������7�0O�����I�eO{�����s�˛.fԩ��p�^ZR��}������ ?x�����\�j�i�^y�Zd �޵[�TJNٵ�%8��,h؇��El"�P�Ŋ��-W=�j������g���\����p����=�X�ϣE�|EЃeM�],�,3�z=�T+z�QZkE�*V�SFj�V�����PXpf԰ �mS�����ܧ��X�T��dc[֊���q�"ό5�^���]�]%,�̀�V$�Zt��'e�K�YfU����vKر�ӗYy�;P���z�F�z����c��*�	��{~�}����E����	s����	'�Ɓ79@�L��;��5}�sOůW�C��߲��Ǥ�w�z�j�^�5�ؙ�]'������s����<�n�;����=���f��k���"�na}�k�s96I�6k��O{>���|Q���>���;6g4�p�k�Ad_��Okt6P�����]p�#����Ǳ��F�g��t�|8�7������Q4٤��m�4�����
e�#S��{�'��Wq����y���W�_���Ҫ�����x�'f�K�F�N��F�����Z���[�����N	��y$[kؚs�]Lk��{�{�my1��o����5�}l����*����=��3� ���y�8O�$�v�Ɂ����oI�1��<c�y��_%Έ��[	ݼ��Nmo���|���T���`� �Hv+��7�C��pW3�ժWݜz�#��S�L���|��T��/l=��*���&��jd��o�����uŎ�V5O��ne��X�.�l�1
����Cb�acR����l���:� � _�U���iz���S�0e\�����z���>e	���8�y՜]�Y��Fr�<������߇�=��X�qK/�({�ܿ����[���L�J�`�pߩ��)9�j�g�ՎYw8��"�y������uԒ���Ә���/��k8Ѝ2�@�l2������V�6�x�1�_�$�_s�5=�^�7��^S��۷t@����##��8�S͕��z��4uW��ܱ�ux���b����l�0+V�'�Ժ':�I%��K~�K*��!������9C�A�̝���S'���J#��f�r����_��X5�޹)���4�h����xb�Ys�w�E�iU'2`���zB~T�*:m����A�c���`���5p8�w�@n��2wo���={��q>ꘫ��]�^f����O��^�T�j\Z]���b����{�z�6{��<RY.fʾe��a��cu	�hf0�j훲���E�]��=9y�$�ek�ꎒt�F�(��{dQ���4'�M�ܠ�p������ĩC�ʞ^.��D��l�O5�O:�(C�%iʇ_���hH�x����<A�ÇvI7� ������8�g�W�<ih1M�Q���w�<��6w������ON�6k�C?Gw��DL�����z%�&p:��W���ۉ��w�_E�a�܇��ߗW�g��-����w�����%��U����?nb�x��������>�#�~Ss��������ٿ/��eNY���r���~'��ƚ�n�཯�83���ץ#�b�)1_�KG<q�Ѕ��
U�B�k+���Ʈ��߈��mrK�5Q�#����ǫ�(;��X(�g	Gr�Ń稾�A����á��oY��-F�4���\�s��g��P�H�T>�w���Lg��}B@~3u<�(�]�S7~�y�5���q
�Gy�-�V��A���x�v1�G���u[oL�����ެ���K�E�\��$mT�Nح���@��Φ �`Ne���������v�~��i	̣a(x:N��&']�s�Ww�]�A�pN�v��0��ڔ[͹6�[����������f<K���U�Gy1�4s1򉻃;wv>�D3o�	}}�E�{�P�U�W��,c6�zc�#��^�r���W�/l�V��-ڥ�ם�7�}A��{�'BY���^�n������Q���/I�(��{{v���W��C{U��e�Me�z_���%Wm�73�F��n�r�M㳚����<[�����2���X45�m�p�\
�f��OV�5�2s/�t�f��m&�Q���{"U���*���5�3�JyU��KX���zxߗ���xﻰ)]���L�՘
�_�)���������;��n�:��9�n�p�F�e�ц����ͺ�0�hM@�_��ά����S7il����/D�����k܇� U?b����yC�}uKB���}���Oyh��y�6�c�y��c��=W��Ͳ�ϸ�s9�g�l������J�3�����;~�@�ӱL����ߊ�1>ȱ��I0�_Z�܃�Z���S��o\����!^M�Z���u�Xx_Mu$+�n����JY,堌��skhs�K3A}�S{�t�@�4��+�\���2U�j����ك���$��zQ�{.��K��(��~��~ʝ�]�*F��ݛ�0�}{tq�A�!�Ɉ��àAM��V�`2��B�d��C3nD��J͝Z�>��uj�sk��c�ܞ�rj�Q��0fCcs��x���󕣻�I�|�h;˩�z <����ѕ�_Vj������ځ3=�ao���9�ƈP����{��eG|/4[8��O[�W�>�`|t\�t�޴�Ny�J'�<w�{�i�w����ǹ�⟗���c�DM��Lߙ����_�'�/���A�K�z�L�|��C�z<��w�ny{]{#� ����a�j|���4��&�c]�ӷ�o�������(�K|懒mA�������������I!z�B'���Vr��8�s�p�_��;@6��sWWV�]1���Ƣ��~���r��y!�}�~��;��Jl��c�-Wܦԅ��GqIA�|5
���xW?{t����Up*��� ��G�I�do�IY 9c���5��ww�S~�wM20�ny�_"4*9�5�Z�A���:����/WR���s���/zƍ����įx�C�M:9g�Sit4 ����r�:�w'2'Y�>�7�ON��u�e~Yґz�{z�� ��7��=Yч������;@��7ϰq��Fkٲ���"];釺�ݏgM>��=�=�r\�꡼K�Ú���s��6����:ʒ���Z�'�+�^�?t�N'֜�$�U�8��Ӟ*�������#��~�ߴ /O��F�>���R�N��>���Ri��e_�o��N=�yI��Dw'����ף9�O������"�n^_yU�@fc�\�h�C3�{����VUO/+�W��s�>���禁�dr��u���@=���w"��X�j��zV��X�W8J�v�5��������m�
���
X3uzz��Õ��߈ח���yV͜�����!�׸��-Tx�j�w�ڭί�L��ԍ�N|v����Un��W'ǐRُ���^MevEQP���h���`gPKK'6�]�ܾ�Km"�(�A��Tx�kaw�r�>͢�/3�c��d�wg*͕x䲎S���N9�<*}���80�9���\3%�����,Π����3P����pr�i$���:����Y�b�b��N�(y	�"�4�oL���O��s�y�z����}1ܑ�n���on��7�5Wݖg���](n�M�n���f{ң���m��>���I�,8��Ě�cU6.��Jm����R�z[��Tr��tpa�֥�Oz����7�|�������������xONs���G
oރuK=��矶�}�͚��@�IޓvBʼ�%�2wI����� �:�D+�>{��{s���^n'1�^z���h]�̕�y��=�Z �#ú��:�|����*�=\�L�8�<	̾~��4A��W��o���.n蝯W��e�`�筏3[gq��o��`�~��*���3�DE����N�f�9��r�z����0a�u��J�*���w�����Y�,q~�eD��Brǽ�~�7�����x����_������y�|�opѲF��WC
��b7^�&�Ĝ��]��]����֤w2�k�wrGmm"�^������}���e!|A䭭��uV�9���VݹC���)M%�u���ºfs�w7���XU:��>��Z��s��:�:iZ�N����D��!Wk5��J���;l�}Ҏ�_&�Ŕ �&˘�ѓ��à�"���]�7B��v�]�-S��_�u��c��7E�;����y0�t���r
��� ��˹۝|9.����c+FN���+��4�^��#Z�uk���/�G�;[�1�ׯ�����B��UI\e&�K�������C���5�9����vv��U�k�ʺ�M2
���c!�i��yi�@73)(֌J�gv�U�"��_u�If]�V���˾ۓZ�'F�Ah�.�+��v)�Z�l ؋�X��WI�S�n�:�b�V���NwR��fc�:u��2���u�[���g��VSݛ��n�-���hز'j�˧e������Y�����нuqΥ�f�Y=�����ʾ�<�Su��6�3��m�m��r�z7PO�ʈ0ӣ<Ɖ���:6��].��L��8l^�] =�Q-���|�k+�>��=�c*�*]���!�4r����tk�c?'��s5vM�S���mP�Ԩ�fL@f�5�8_\SN��X�Frį��\ҵ��D��A���������%uB���ˡ��7R��Wc�`ؐ76�xU����a�Ta�𽺱EZu�ΦU��ţL�J4�$�6��G�O�Qwֲ`����k+�/�ձ��3��Pus:�ԻQS����p7�j]�o +7/`j��Uf^d�U�1^��>���y�ro^'˕�_`����:*%$#���9�f�2'
�T�S��k0U�?��=��T~�V��r���g��tU�i�1[au������W�NhŹ%�fw(��K	�9��u����qV�[��֝u9�ɯ:�g�p%�J���RAfT;Z��1�����]n�%�[���>pLR�W�RU�8Eg�8�J��Mǥ�����y�p7Oi���8�J��V���MC&�I�ʴ�-�fj��_ʋT����iK�͡�i p�a6nQ��q8CS���=�OჀ��p;�#�T�wr�ǋH��̕j�=���ΥQæ��v�:��8�1,�j���:%�=f�KgP�{n~��0�HFl�Ћ9S��rm�Tf` a�3�B�q�%�'a��pK���U���8��H�k�邵�õc�$#r@���Baz/�4�J����R^��R���Bh*�ek���(]8��b�A�{���`[�]|,A�ut?\��������ۚЫ=--���3k��tX�!�^����uwn���%�I�$mc�L�gH	ƶ��)dq9�je�Y�wс˭e�{{܃q�r�4t���堦�}u(�4��Z˗h�����`��Uw���+���l�(�A� �����T�?>c����[b"���"m�|�1��/�;�,_#q�S[h���^mqf���td5��1��ULSy������cl;{��A������Ty��iǅ�+�;��5��:�8���w���yk�ƚ
#��o��tb����5T�S�G���A�(���n�5[���QWc��ѣ�u^x��w�h���Q��e:e�!.~;�Ruݷ���y��g�v����&<���
l�k����i7c��V�C��#��Ρ��n/�݈f�͎��mv��e-Qmm�m�mYM��D�͍�j*팝�;�d��DX��ص�i�WZ��tuG�xo-Ŷݞ5�u�]'\mc`�X-b��y��v�"��[V�=���'TE��Qi뢪�&N�Glv�MMv1v�F��Z"m����m��Y�1AEžmV�2�v�QDE�$Z�DѪ�Em�N�(""*K������N�-j�g��O���*(�������;A��6�h���4WN�J
.���93ECE�&���m�N������d��_?�L��eme���/T��N�b�d�y�c�J"Q:ܬעc0Lۭ��̟B�c�ܭ	���}\�vk����嘾�t�������F'r��`u/���R��"3�~��ڊֶ։w���������?�ϲ�ӿ��B�8��m���@���J�N�f��0�v���/��K],<c/)�&/�Y���E���oa�5O�.`U��/����[������xk���=�A̢g-�]޾�T�ء+�	�Ѥ�il�울�aՉM{��'��w��h���Ӊ�����]yB���i��O�c"�g����x?�����p�wQ�]�j���J��;�dJ8�E5Z�u�M^���+�.���37�l������w�7#(Du;�������[�k5���ڨ(uS�[�<�Z�5E'6�E6�h�jeG*���/ �zf���ɻݛUq�6;:�K-w-ö!��v(�����aJ��ӓ�U�Sl5��	��y�ge��άۚ����rg��D,/�lc���y(����s�÷�q�	��ڲ�.���w���B���s�I������0���Hsbc���Lx��dns��nk����!���T�k`�Q;W�˒ρ��6��訢fA��u6�ln�pH��m���gT��P说��pT�T�@w@:F^�t�Y�OM�I��[NO��<�K��S	j��Y������lԳ��P�Zؒ9L�똬�VM��	�[�q�UH�vuc�u�ŗ(�*�}b7��9[��n���l��v�`U��[�b�嚽�|N2��I��m�u�ǧ귊�+a�C�~�q`�%�p<y��gJO��"�*-k!j�LZ֐25̸CK)m�w6��w?�t�
R����s��[�{�����֌1��J�me �D-aG��Ij|�ީ���z3-u>2��P݋/�x��&�8��E�$����� �Q�֠�LD U���N4?"�;[���n���R :��hqͿ�#��9�����-޼L���6�͗�"��F�o.�Z#�{yٱ�P����L�Z�e�L�zE�.�i7��� ����6���ۅ��_oa�|C��m�ZL�qd�ЪzZ�p���C�v����q�M$�B$�-Hg4��~u�qٲ�n��8�e���b��9�F7���vOiq1��L�/�����\g�s�TɋWվ�C�2�Zt$r�,h.��yFm����G�u�w���	 kV��\bofb�^�I�1�e�Vb��+o�ş1��vd�m,��?�G���Ȥ[��T��Wzę̗�(ӌ�7��<��**�m�["����Y�rJ���[�p�R�^��c�<��>���1{WI�C.ٹf(�;�Ԓ���p㝮a�sr�j����c����v��t��}1�E���ά�WG�Q ��N��k���ןɹɌ[���98��ɖ9�����Uf��wWR"��K�=�d*jx�l�+����qG�i>���h:�(8~m'���03��o���<BO�G��R�{�9fbj/.���)�d*ɗ�_n^��+���o��e��CG����w�:ד4�3/^=e���@ǟ�qU�Vn�ԙ�v�XjT�E�q�P��*-�hǅ�ɛ*�=i�k|������A�D߭0�P�Ӑ�2��9��R��zsC����>��ߟ�C�����v�>_���̼F5K'���N"=�����sy���l;�9�}�PR���g�.D!�rjwp��B���UV5�k�0�Ly������ �|U ���ިOAdw8�	Ia>Z�/�8/���u�c��1n��ēq�/�$��$oV��dl��%u�o$�*
���m��R�'�b��^zK��%�@�A�p�L�_�9��
�3�%���`93����)��l(���j;ϳ�X
}j*��}'`29Z��ԉ��vǃ��jbyQ/��{W���\Y�&26g\$�������R��� %[1/�uf��P���T�oT�
������`���b=C�ϸޠ��C�g�F�p��2��Y�u�I���F��-�{��¹`>�CvWo:�����+`[:;���0�/fsGm��9v�������L7Nn�Y�Sw���2D������8g�[�P3��s#=��(��~2˔��kl3z�ָf�^
�۪��cm]��Qы��c�8�d[�mܕ�͠��a#���g<匕�γ�����kH�����$��{���B7���A�ʓ'j�ܱ�M��e���,u�bi�P3� b#����d���9w<�9�3�uA�ooԥж���`:��U�k`�!4H�!2���c�ƭ/�������GWf[��z��T#D�2NsADc��7�S=��+�	9�Ǖ��k��5i=R�WW���R��}�6&@��^b��W��T�(2Q�F$s��U���n�
���;Z��OM6i���h�k[� �K�jb��y9�Do5S��K��$��v�2瞂̊�x��f#��6�����"��z�4Kۘ��&�Jn⦛x�j=t��Ƭ8�e!����b�]?'˞�0{�Q�ρ��z�Ɨ��?��ڇ�JJ{��sX�ܔ+z�?Ra�S��12��[}�[R������\�A~j�����Xϯ�;{���*3��ͺ�k��b ��d��|a��������GE��{	�0K������gY,�O���A;��#S�qk�h�ʓ�X\Mչ�n����+[0%t�,w^x t���7_G^��%Z�>�[C��oک�cA�j��c2��G]p݈We7n;2�>�i�YF�rݩ�6�����K�^��_�&�$�aa�]htM�;3q��-���VXl��:��6;�u�)M����ʙ�;�24�Z��p��-'Z�m�cl�3O���f8Ny��O��:sm"5����k���v�X;UFH�Uh	��}/R?�|�z/���G5`�ad��@6ݪ<U�s��;��>U���,{])RP|ޥϺ`{)�km�3jO�a�-8	���blr���z�^�0��7��E�S���9$Wc��n�N�,������qF�c4�Gћ�,-ׄ��(��ۺ-���ծsh�Eνc>�'D�,x=���Y�D�}ɩ������9��4���Ƀ��u]��d���*KZWN�Q�M�.�	=	��8��s^^USov��T��G��M�]5��\����I�K/j�����c�3� �j�,eԶa����9P�V׆%4=�Z�|e�-��<�k�a.�؛�׻��6���$׮�ˌ!�Y��֔��\�7j��q1�f��H���n��b�h�j�	x�Jױ�`U��M�7� ܍�37�l�����
Jh�∯��߮��OD�RJVS[Q�7��;�AP��s�CV*Y�*��)�	Ė/�����*@��^��æ���V�vse�Ҫo����y�=�ǥ0�qn��;�n^f���H.W��ʔ�ր���!>2�L��q�[{K�]n󨔭B�{Vjr�k	W����S�J)�����|�/�GTtIǿwE|����l	lԦ����{�yt�4��L��<�u�fK��;#��E�%F_9�����\��\[�T��%���B���g�7�F�qi�!��h�;:�˯q�e�g�?q-���p����E��'P��<�UU��"X6����ݻV�ض\2ge@��F��f�6<�l�.%1����u��[K>�!d�s�ӱuY6��+x�]�s*3^�ꑳ�a� l� �e�f(�nY� ��=�§C
!E���1)
bv�.SJ�E����[?��d�Ԥ�6�~\�C�6jv���hj-=	_w]V�/��.,�AW�c7��ɻ|-�:���9��PW�6�>3"v	+EcV��GH��s�Y�U�2��iO�<hu���N7F�5�p�=�k5H-���ێ�!vu�����D���.��.���[~�Ρ����f�����E�M��kK���lk�W!��)]!֨�+�	���k[�m8�8\w�S�G\��8�״��m�Ú���"^�y5�Μ �f�gb�vvJL��#�ˮ�C8�a6����5����'�Ƚ�B��}�VPz�w�Cu�3�*{�]݀(�3L�ӛV빃X2�i��8Js*��G�=�O!-��A�^k��3돵����eAڜ�V���w�Wne(u<q�> {·z+0�-�2��w����o�Uy+������t�?��i�nO`V�u�rc��s2�J��/�p�u��=�ϸP����i��&��b��;��mQ"u�=�^���Qj����,��uR�p2Ff�C�?R�T n�9� �צI��Rb�d2����V��]�߶ZK�΋d��z��gCY�!	��M-|�A�<�J):�%�+m�ت"��k���Δk8�}�~N��4i���+�3��m�❬���d��neω�>���Y������\�vݧݩ}��R��˱�#� ��_Ij,w�u��b�b��%��%Rm~�_z�f�V�s�*'}1<;�M��P.Fmź�i9�aP�����A��f���tS�_V��8}Hh����tL��'�Z���u�1��"��Ꝡb�R�3Qpq�P�A1��^ݞ�����������l뢓�y�޴���LS��Ru���r=��H@nc�K�[E(�f��9����:��W,\�{��N�O�y���P�dÉ�U�,&�#�x����(�z��U��W8]�o�E�Y5==����F�fR�ghG�G\6�h�P��V2Q>�XY�nec�kj�����z:.�K4���TZ��^�yz��yoG�{�_Zw�3�
S����;�G����W�7L�&�LO4�Ы7��ۻ�b���hm&���a�ˁ[O��[|7���x�˞7�dd��s7��L���ڦ`�W�tGfqѺ
��Af�'����,��&��Y�ffnV��l6�r�ڈ7n
�	o-m穘���QL��:�z�N�~Jz2���y��-j�V���h��ULZ�t[G(��+m�%���Cfr ���c鿶\�O��~;�W��$�/%c8�4�b��c
����s�z�26�.��X���d<V�j7eHobh�"�����΍00�4�U��A�'yߎ�b˲����m�5ÿ�x��G)=Ռ�j�[���S��mq fS�⭷R�#Y��-2;�H9<�[�{���#p�p�w:*�^)�^`B�s����#��⿭`��1�F����0�!��-"r���=6(�톒w!�-��a��#��do *x)ƶ�&�Bb0���D��D9z���y����F�,��_��ƣ5_��o��ʈy�*.��'>4d2
����3�Ncs�6O���p��b{�νM�I)�}}�0"���ĪK�@	U'��dd���La���Zn��ƃ|��	x�%�nºl%�j�/B�R�	u�ђ:�V�E1V:w(:VG(�����/Ss�=�R�@U�_u�;r
�,��\�����I6��c^tB�����p�U�0N���xh(R6�vV9�k%��N�nM�x�ß�}U�W��{�\񧬙�C~JaAt�e��S"����2,�^�g#Na�`e��B�ojA���.lD]�lK��i���"8��?D�L,-WI��4�>�=��=8�/^���~D5ukC�KQx��ݹL�Dv��tݹ4z����2��򧋧�6�[~n�P	Q׶~���1eV��1�خV�2<S{�Z���Y�s�*��7���J�O~u�#�ɝ6�|�*����eͮ���c ;p�]��gI�haa�V��vf�y>�so뮍2g�}�-����I]=S��]��$tT �&�@s���f���,1��Uy���+"�F��߾�|1��[��נ�zx�!�X���j�3��Z��ц�f kC��]���d1녗��M.i�OE�g�km�N�c�l��&C�zLפw��u��I�I��^�����Y���M��8����͎w�����1b�9;׊�+$��/`�Xha7�j�؈S���f�r�14ƛ}���o4R&�.�#W��NH��MF�q@�D�M}Y~��&5n_�-�.S#~�V
]�8㡜�
}J����*^�ѥ�-h\K�6 v��{�y���+H��Z��W0G5�x���b�e�ޔ&+T�UX\�[v�;�)Y���m<쾉����ɷ2��!u-��fH�$��$O��������x^P�cܭDed*��S0ԠZt���y��O&-�yS�Q�zKi�kS��dNH^g��~y^~j߉��Yg�y)�q�0���5JY0�=�S*Wj�<7�#��$n�O���6�Rhjd�/q�my@�,��
��ɾ�D=wy�ݣڡ*�����N ����:mWb]�Rf��tj�tO[ǳ���ǏXΨ�s�Qff�� �5;ݾ�wC�n�y�E�\7Һ�o*!S�]d�뵴�x8����>����-���
r��o�4���jF&atӇkL���,<�Z�׌��6�*�0�u��U"��ZrpV����ݓ�)M"b�z���V�u�%��d�nǲ�>�Kz�X����n�[|����2�E��vE�"Ȓ-e���2q���e���E�,YC�ye�jފ�EЇ��1�uj�u�ђ��L������b鴃�B��Ss������1���\-��XjI�XFWn6<������6®+�5��M��,�ъ�=��&���)m{Sy��8D*�b�7b؂�+ �������=~�G�����}>���x��G�=Zw��o�W��^�"�4A�D��2�n�kD������\�4jH2���"X�VP��Fq�e+,��2؜����g\Y'V����r&4������q�;M�|Q����s��m�ivvk��V�-���x�T%+�J�gU��:���(���C�P�% ��ˣ�9���#\J-���A)f�"�X�@���W�v��C&��p=eu�z����cr�Q�\S^�m'c�P�Wu�7	��)/4ʒ����]4[�X:c1׺MX/�Тo�l�5f��b<ŷ���������Vܒ�@f��okz�B]w�$�G�Ľ(����C�X%b}+�hט��y�;x�.t(:�4N�GSLn��:�\�ə��b��Ɍ
��̇�A+aMs= ��y����8���ؽ�K��'��}$Z7
3��I����ՖHE�+"�Ct�J��Z���B\J=� ���Zꓽ�:���s�Ζ��j^ɛ�
�/%��5W���\[���-�t��Kh����ˍ����
�֖CFؤ�n�(�=��S��Ǝ��p����`�y�M'{�$�F�VL�YE������o�5���6L��*K/z�eq�Xy)��_F�Ҵ�]g��Mf���;AEI�g�5���n\s�[�K��i��L��)��%��}&�r��CsEMe��[�wy��t'/L9�+V��BRYc�5���Ӫ�ӬXʘ�
�ū��rk�93^��w�$�F7���x��k("�b;�A=u\�p[�V-�Oy(蕖.��vK,�Ҏv�������JA��ݡHh�4�"b�Jw��Y���<)	�Xe��/6�Ĝ���UR�C������X#DU��t{6�(u_h%�b�S�Ww٨��Rj�AmAvlQ�%�;|��m�v^�Ya��k�H%�A��An�Nԛ�����ͮ�G
�u�)��
��Z��buq�뫙Vb}����dV��Ǜ_g�=���CU��Zct�އ���q/-���Äʀe(�}K��s�.�fLS�9�|�]����ӥb���BWl��G�f�)P�.�ӧ��EIvK�I|����y�w	9ҵ���LKYw����TP����A��S���1\�c���njB���oC������	f��wTU�˽d�D����
K�x���>}s��-���:�E��);p�%�V�L�����U�C(��4��/D-� �]_�a�bHQq���X���;}������6*^
�ԣ,b���--r}�;3 �X���a:����Ҿ�8ӻR�����N�$�;�5׫���Li<j�lJ���={ќ�{WY�r'�t���`��i�Z�2�l9x[�l	.)�]�f����	�)vw
���-���p�l�Gmguo�!i3��U�k�ps�& ]9�IB��p�8lB��O2M晪Ӗ4��Л]Ǎ���{n�CF�ծ�M����(�]�}Я�I��H<��}8� �[�$��RAT�B�)�_�I��� b�*+�l��uUAQQ�E�����mRE?n�EUQ&�55�e����mZ�Dli����(4�����(���TE%ֶ��us��6b""*���Z��y�DU�QF�"Jd�$��E�6��h��gF�ƶtE�K�QTGwlTth"�����`���#`�5�c��TTU���������������j{<��OZ�l�4U�jB�1I֦"���A|�TQ�b٪���͚��cF*��F

"z1T�%4EUUAd�ڢ-�i5����$�i����#���w��$�f&"�T�E����fڂ���kQPQ���ӣ����l��-6�6�5m���glD�Wgv4IY�X�
����Z��Q5ڳM $P�~�ɬ3�7�^1��5*�H��uȇq�ڑ�h^��ĨWp�;Z#���1I}�y����ku�-�4�n�R_l�a����,]Y��*������t0�������{��S�udW<Ew��r��4�3��J
�`F�#C�5�[��6���ҭ�C�(Ź��Z���X�dvۗ�8�H�ơk�>��[!{��pZ�v�Qo����p�4M$S�H�m/�]Kb�z���`ᐷb̌���R�R�n\�;Ga����1Y�F'J�i�\�jqO���z=NMq�q���a�s�qTE���A@'��t���g�W)��-�1:W��=����4���v'N��f�FӞśj�#�ԀIMCV�����mGij%���VsK.�X��gd`!x�-ٗȢK�g�K�c,�[{�5�5G�Ġʞ�9(7_�l��p� j����j�2k��qDD�[�Wu���g����P�	�����W�A���6��\��F��6ws��\�[�XD�3��eU�̸�Fp*5@���XΔj�Ji����d�cq�S��Xq�pϽ���U�i����Cm
�q�.�*�.EZG��i#ײZ��6�B(%�ڭb�&�x	&�������ѻ�PͲ�dSL��2�P 5G�.���{YϮ��L�ʥnl�}6�R�]EZ����v���6!��:=o�pd���U���7FA[�9�I�9�f� ���>ER.��^!��Ko��{E�T��vn�c��O�Y:�9�W��ه_�}� �vv����������W��n�ͯW�P.s�-�R��(G�y�(�r�n4�ȪM��cU�ng��U�e<	�������)ՆQL��(�����$�S�3
����eǱ`��C)ͤ�w�1��o:<������a�q�LS��M׹�v@��A���>J��M,*�ZIͷ湱ՙe3�����x;;�<����.���f�sH�dp��i9VTE��4�;�9�n,�^�O؊�;�f��L��_��L�6*=�����J���|�[�=����i��TK��3G:D���#w<��.�A�&�
�	oQ��f;\߶��?Aoe�%`�P"�j2���O%�,�z�1;��T�=7��L>D1��[Tj ����P6�CTt_J����ry҂�]Ғ����=V����y�'��ʎ�­F�>�d:;z�26�˓���X�g5����<��[�E��Y��59`�r�#�M�:�����Fk
%��8�֗,�1��Z�����,Z����ɽ����n�\��=�'2-�gAN��zd���`��H9��~�ڱ����:�m)�JQM��|���ת��7I�7�^J��8���3N����ǡr)c���̧��Y��Wz[��tM�t��g�9�'���o�/�F�Ε+iٮ��cG�aS�
j�ac�-����I��()�h�e�kP�Ȇh�
�)�qO�Ք��g29O����_}�>�u|�y[5�~X�&3�k!�`Σe�Ԝ˷s&U��e _��qp������Cu�Sٷ��I; ��SE�F����9Y�J�����#�$��]�A�Z <](�`�!�8��E��]�M�۪	��ʘ}�i^��]a���A��v`A�)�a�-�'#�3�	��3�;݌��lx��8�\/��X��M�,]��.��3@Gx��d�^y�M�-fNzr4݀�J�9������=����wA��m�-]c

rr�#ci��9�$c�K��6%��q����\���u��H���N�ZU)���/�K<�����ϻ�Yό�S=�i�\��c�9��q7[�fi�Ë	�.��.ʞ.��2�ݪh_X{~P�5����nT��-�p*��Q>A��Q�����Lzg:�րۼ���W*�DA�η�`{%m9�H\����5bI����ֆ�v�;7멖��%��dl5���bq	��^��2\�7�u�{�����:7���0�Y`��O��PX���¹Ѩ���'�����Z�u�GL�Ou)�lpՂ��_r���f�v�s����EFK�R���m;�.\gg$JZ��F��*2�;�ކ���Jx�P�M5��[��d�F�֨���
��+����,�ܴN;�m�t�U�u��ƿ��0���Y��������QO���GuG��k5��2��bvae�k�����zN)O3N��f�)18#����>�r��!_�^?5c�2�?|����b��[�9]�W����R٦��؍�v��s����,w6��`Rlt�Ǩt�&F71s]���3E�T솄��@gd��[�w=|xT(�C��	����m6
�k�M�]�E�6��ba����5�;��N"V�]���c�u�R���Z����C|Po弙���?�؟�T�u��06�I�1]|JǮE���`�{8��{!0S��0�eq��ЪzFbR�����@Xe���~s[=p3�;�p'�ݵ�a�(���0��R�̞�W4�`.چ(��d��)�eT�-��xòfpu�nFF��J`ay��H�ރZ���A�P�[�Ϸz�NW�^�Es�&.%s3]2�¡Jt4&h~����Gt���ơ��5�G�H5�����|�����Ȧ��y�7pc�kLˡ�iZ|�,u�:��G�o+ք���#v)��l"��~�%Tu����_]����L��gҿ�tY�.��`��ϕ�5M`��}��=���A�w٦�'_T��"���S���/�C!En�ҧЅ���k@^��G,�C[M �v�vђU[�gox�=N��XWO��6�v��nn�ҙ(p���t�{����:��7��v��#;�)X)��*�/����������@<�V���#X��qڔ��@*���/��O���%��Y.�hQ��T�O�z�N�f�9�޺��4	zP���1�؝�͡�4bc��)�i�zˀ���t��v�vH�Rժ�Y�2�r���ݳp;I1VE��ƱY��^]�tJb�\�i�k˸F\�^Dn�~��:��)�=����KǷ�%�(lc�m��`㜎g�R�D�������oR�\��z�t�`_Hc�g��V�i�g�cm����G�pi��r���|�J�S���c-�8:�t�Z��Q�#���ri��`KJ�:Ź��-;k�gjŸ3l�Lt:�֠[D,�4�*�"���p����m��PGvm�P�8�-K��F*!W?A����Зײ/u�
��V'I�j����4���z���|�Uf�s�������V0�3K
�I�*Z�p�u.�FA�wK��0/�N{������:K墶�㮓��@vq&7�͌U%l������\ͭ҃���6�m�_G0�q��ˢ��W3�j���6�a�복�����yFc6�=����l�hV��cW�w(U�v+>�wK�J{���x��dN�ȥ�*�r���Nv<��+*��)�݊'�|�u�sjk�\�����=#��[�GL�ė^�t݃nt���/{��@   �̆�6J��p+���-��}��UCr81����FD�W��Oǰe�T�bg�Ą�33�~޶jb�����zXS�솯K�����S��:��W=�3��xad�����zʜ�z�ݒ���t�<�*��SCj^a�҇���;Yŉ�ɡ��W9�]@��N���eE޲m�n=�B�y�4�X��b�i��*O��Kя]�����E�.3$�-��[8����<L���O�[b��U��6��ke�������qJ��n7�j������c!��JC4�o%���N��S.~�_r���J��9\:��'/=��׊�y��~l�*�~w�2�\C�R����~�4�W�ż���˳�y����(B�?%�u�2�\��q��_�ϗ��d��sU�O��W'���C��	�u�kH�dK�0jO��<&��ϗ���ߓ��kLKk:�Z�򠝷��۟t��B�qT���ިO��s*�s�jn�)����je�/%%���\���A�qL�ÀV_�E�3�fYˮ?��4���Y�u��S��$�D��/E��$�ɇ�[0������or�x�mv���v+<ju �Ik�8���8}Q�L"���q���/�e����`�yP��$�:�V<Ƹ���9C���7�S|����b�D.�ƯL�hb�#8���Ňl��� {�G���3����fVN!�I��Y�u�UM��Ѫ�s\&�,�	ͷႳ9٫P��[*�)�)�a���s[j
�Zks��7V�5�fί,J<�����ޫgmx����p�t%eJ�WM��uf:�ii9��z_F��ed�S	Ҡf��_z#�kL�����J��u�u���.n�7+fH��@5䈐���N"�->ֱ�&)�o��*�Z��Ƈ�$��>����4�#�
���{�7�"�+Pw��j�fs�i��ky�����Tr���ծX��r'g5m+�4�+��������L�q�0�>;#\SyA���P��!��M?tɳ��g���z^ O\҉�+Bƅ�smt+u�	�bʈX]*3��u��`C ��a�٫X��VNM�6�mg��<8��d��_��Yfy���\Q��D����ĪK�BUI�Pd���"?����%�m)�h�/#������J�e��t�mWX¼TfL
x�	Ȩ�֑sMO�j�*��xV[�P�4�(���	g?b�-g��G�wLq��蓓Ͳ��U�s	��T�}�����S*z�cP66�]��ޙM���k|�	[K{����3݁݋���p�l�{�����)��؎�_Ń\�$��֤e�%9ݸ?���V�.ܖ{�Y�n9
�(뜱��t豔�q�
u��u��F�l��\��W���}U\�n\��#/���� ��Y���F�`Zl�=Hq`'4�y�mC�4����)?7@�nI�st$m����l:֥�{5ɀ�<���8
���-:����s�'#���7S�\��3L����6ږl��R_�k����a��W4�'5L�aa��U���N�_덍y���?�E��(��'ȇ�T��.S*�d(�c���1��Y�F�x酂�Y��l�/¹���n���l:<�U����n|�uͅOK��_DY�0��޹[dt,�:M�=!�Y5�E-`�������{BB��x�Ս��4.^<�6�����^�U)��qqRFW)k!�aN9�{�6��}ʁ���b�E�x�xh��&�z�N5�b�C&'��f�X���-��w)����q���Н�D���o6�/+�T9,f7��]#;����N���J�ܧ���pIYp�pT�b����y��ȧ��y진�\�zC4m�i��
�i�d��Z�/��FîO��8�ҚAa+���g�No��� �a~є�R?1�B���[��Vz���Q�$���s�F�=��]�+K���x��T�۷�y*��x�q]T4p�{faJ^u'kl!����rE�m"���,��y�ȋ�C+Vj�s:[��d?P�{!������]�F�y9Z���[�f�foD� �9��y*6>��i�����\���])�A�R˜��7��瘙�8�?�V~���N�wJ���Ui�Z���2b7��M�K*�J�ƭ�a1�.��}��f�,�iX�\
����s_�l�$g��l7Cc>ҜƎ]���G-�܁',`+.K��ժف]x�%a�n��l�L Xy愤��#v.�����B��U-x��A�b��u��g�cYW�q�R�]4j������9+йz(�D.����<�H|%��B(�P$,I�;��̓E1Ef"��Ts�m?q���Z�bMІ��/���3�|�74@��3�����muGnoL�1��Vy��o�q���$��Q��:/Ӻ����`qY]u�۷ib�tB*�����f�HH�fx��R���6�������v���M)�jIȭ�m���QO7w5s��91�)l!��y1l\_}��B8Ȫ��V�v�X����V��Y�f�Ѵ�;p���lژ�pЍ*p�D���ܴ�Z�)G'�́�u����ti(�ز:�Ҫ���z��'{5�i��v�!{E�-wӫ���mu+A��[���S�fMm�����l�[����G��.^!*A����鞛|��o$i<�k� lWI�����A�?X<T<�P��\wïN8��]��r�f�c̋w��˔v^0NW���o� +2�3{QU�=���{Մ�g�&����K�\�c�Rئ���Λ~�M�Xzs�j����J�K������j�1:W��M��V�������0��u�+~U��mI%^�ة���Yw�q�lUBl1�qd�g�.���]��S��~��b�5�Gy��橊�L�@���(O�q4�J�h�)��yeэ�|Ǆ��:g~�#�ٟ��%O���(�7�7=l$Ϻȷ
��)���+y����At�;���ꤵ������C� �hDz�12*�E���*:���G��J����'�h��j�7c	�
'��FF�ƜU«��τ�d�2|�Grj4���,gJ#��y=T=��2n4pw^�-؊�5uSث'oZ��u��l�͹p;��	���b R�� ����{E�~�?X����_?���(��^I?���7Y�no���be'8��q��s�e��#�F�ò�{�O�ol�+Y\�X��'u��A��@]�Xf����!'V��	O����t��E�����\��������_��~��}g���e��Ĥ<�(�YW�i�Ǐ$��qi�+4�y���o����c���K2�������&�n�^��������

 �dR�r�YAݘp�	\��#�l��1LWv��!{���L���*̘��9��ʴk��ՏfGWl�K�]G�"׻$��2��e��ye	(�;@�B�r���V�X	:˃�`�k�����ޚ�J��5W����'�Q��d�4T;�.�b}����Ӌ2��\�F�tUC����+?]F/IyX�S�<�F�{����$R�,#�_�s垺��2��e�h���1�C�G܏B�#N����i�kÙq��t.e({9B���帅_:�9�ĳ];1\�囁��L��QNm�ǔ���xz�pk��ZYJ(�*����W<�Y+�:���.�˯��e٨��Y�3�����O/�>�+-�p���ft�jó��Ƙ��~��u 3lɝ�f��[<����~���_f�2�Dv3�&��5X�FJ��T�
̹oM�k��|�&�0�@D�Vm�pע�m�TPa�+����;�X�:P���I�H�38IN){�^�+�`LI��%ʎЈ�pJ�`vQ̣��	-8�����5{���>�aٗ��݌2��2�ʍ
ms�|���לec�
y.<�����n��SB	��7�-�l�e^�WuϤ�r�N�)\����f�sK�(d�)�6n��ׄ��\��R�pN�ԙ)E�pV��ϴ1Mr����fD��(�� ��z5�U2��w��G���s�����Ǘ�u\��]@;�҆�;���ɶx��I}�u���b��Z��D��v�tm8�a�ZMV�Sw��#+{��N�Ņ��o�v�U��"�	�IC�f�t�B�Hrtndٛ��s����|�e3�ᙐjw��ӃN>d1�)SF���r�!k��-h��u��u��Q_�K��M�Ʒ��4cr�n��(�%��b�m����E�BJ���#���g��e�BM�mq���9R�1>�U���c.��̩���J{��vM�r���y�2�-:��;6��9��Xظ�z7�h��-��G1��a���/n��!��5��*�Q Y�Pԧq7&�T�v�H7��	I���Ӭ*�{u���n�G:���z�	vZ4/&�1ٗ�eA*����(�y��Ǹ���f]yS�=������2=n�v��˂}%�wF�d�3p�<�8E��!�W�e�OВ�8�fB����y'�ڠK�N�������Y9K��}6#aYُܹ치q��XFLm��	X�#YC&D.Z�tݣ]��WKRW�/�N���"����1�����z��x�Y�"�Y/��W*&;����=/�E���R�.d����I���nI��fy��TU�
���A�x�ubkX��3��y�ئ<6h�F����QSTTL�3D�Q;h���h�4V��TI�AUUGlk5u��u��Eݹ��"���3�EDTv�tf&��u�*�j�����UUR݊�STU�NΤ�ӒJb����]:���D�U�)�5]��h�5Q�c���j��T�L�I�4[h-&�m�*�*�lLT��Ѣ���]�Ԛ5%kU4�Ay�/'��4Q4�y�vj��3֘��f�f;&�ƣU,JEQMN�:���'X-b�-��TPW�j)(K�C�������4Um����ԏ�M�r��w��׺9^�����V�m�F�^������8�f֜�xDf�����`lg[�YsL�wy�rbv��C~x�{��E#ћu{[�C�Zz����|������}׆�a1Oa�Jc�:'���c�����ܓ�4��s�,���K���K�S�������N"���BF�>.�n;z�,4Pn];�����B��C�X`�H&�$�VrV��wn宽}|kJm4r�N���fg]��uΘ�^���B�}�g�a��h�o,��a��	e����|�Ӟ�N�ُb{U�k��e��s�bH�c�Y�u*���o�ΣQ5���Ma��g����9g,U�j���Z��7��Mh�j2�_
���V�tv0&�?�FH����v�һ��:z�Brs��.���'�b��6��ԃ	ҳϬ(�U&�-�֎L"a��˥��^;p��V+�3z�`�5��w�}�"Ѵ*�����G����t��}\��pPn�EE��r���~�\掟Oԓ�b�SG
�Bj,�^>7H���45� ��6��u��M(�x0�Gj8�Bf����C��͊F�}|��SC�-d~�������C�8Oi�����k�|�*�S�u$R���;��n����o0q��Y"`�0���a�Zh{}B��>��w���%�a�Ί� Uz˝�Emv�X����m�auOzT�����7e@Fcݦ����N��Usj�r`Be��Ge�SLw����{��0����&�UT���
�%���A7Z��N��E�YD����@K���K\�J����񑓪vw{�/X�m�k��j�2�d���=qG��jD�K�+�Iv"j�cJ�^4�Vѵ����e����4z��UXWt�e�⪙+��m��m���YX��Ȓ����Z���k���O4�pK���5N�N⋶�kq��|V����0��Sw`*��E�F�ߡ��jƛ����WU���N��/%�K�l�kT���C &���{�"��1J�{˘�.�6�GUv��,�r�e��T�7��+?0�)����$���}��b6��D��fr�o,����lM��7��/a'�������
$w=Qm�@�;<>��!�k�^��a1m�aG�fD��V�L�vC��SZ�J�[Je�YaE͇+��ӝf�`{�6�[�껔eN��|Z�-w�>�1P�t�^<5�4S��,�;N{�V��v;�ީ�.�.�!�!�8��t�yN�O�M��Ώ*��r��qe��y�t7gی�,��f�Ԑ�s2�t�Ⱦ�4�i�5�v61�s��D���(-ۗ Tj^b��9}�lXE{I�F���|�Q��W{�Mw�@�43Ά��
@�5�D �^;�Qɽ#�P]�g*R��.��U�����0ɲ�X�ޫ5ukw��IM��s�EC|�C��ajpp�9ܦ�A���<AY�MSM�d�!�;'_^���>���њ6#i��)ߋ+?Z���blb� 2��sV��ik��H�XYé^��<%�M�J)F�VV�v����6���W��҉�������O� t+y�����ub�vt������%}����˦�9�Y��C����(טnQ��VIAо(g����8�{ywMv�Ӓ�/׋S��2�1�S6�,q�٪�P�l�.�K�����v�.Q�P��y0{N0���ÃZ��1c������ޙ���`ln��ZvOh�3c���c�Ȇ�տkӜ���x���5~�W�B37���ַ�eW�m[	�L��`vډZ���&�J%�e�9T�iekZ��û���dO:��,y�1�@��)2�츨�6BFh	�}4�9Нc��)?9py���Ԟ���-V�B�LU�2=�Z��x����JK��p)���� ,�E���}<���+�r��8!��W���Qe����&�kI7 s���l2��zX��KL1��X�V�®w��;�'gc�d�1E'��UO����e�*�CH��2k���`���[���m����Ҫ_��ع���]͊�A7�ߞ9�C���V�Y[�(�Z�kx������#9;���s� =�%F-�B��ā03�s�g��!{��4f �vr�1��h�©[VS�����Z�9�v��q���=�9]���� u�l6�W_@mo���/�|fX���X�=ˢ�Lkm�X6&$��Yn_�����g��	~g�l�+*8R��K�tn�O<��"���d��˔_���}=u���)��}��U<4��T�����J	�F9��`�7����΋Ч�y:hY�����	��5|g�pA��Rtz������ O�� �{�Ѝ�	I-�Me�����iaw���W�9��L��+��~LR���/��|$��9��H�j�d`j �o$M1W�
�>�u��v)�]�g+!�SM�
�s�-^�	܊�}�\�IN�o���d6�uK%{a06�˘"���ũ<�[��W���9�j�C�����b��y�I]�iԳY��f�ܣ؝+�L=���#(��졑�b�7����橠��&�:..�4�ͤڏv��\oL"�9�;+�x�.����y�w�^�X�&�����>�x*[� t��7p������#����������{��~���(=���I~���w�P/*:�E�SJ>�����]?�6��F1��Sʘ5�:���%�
����L���*X��{���y*�R(�]�`W ����'#7F��F8Gj�;8���`�L͏e^X9�3��[�OHjM�{JHw���˻�O�m��a���p��D����"_��� �ɼ��V�E]G?����>o{�f�����6�r�r��n���m��j!��z]�c���3Q��[+�����2a=fԻwj��r^"N`�v�խkd
�c�cR~��(^߂U�>�v��a U�=�`$���K�c�Pɨ�6Ч������󎱛I�ne@4Z�12����͑�"mD���놵� ��Q2�#�s.Y婎��p|�4��!����~ ���(�\��O�}H卿I�ɂ25؍z��ʳ;r㮅/��7h��u��(����0U���G�Ԧ)�:�L�D�u�=�j�3U"f{[�8��k�^X.���R��e|9�㚬R|O�|�&Ek�!�фNrD#��v2���Y8����S	;L�P�h�HQ-��g}���wi��oc{+6DјP���q	=U�C�8���	�����|HT���C��.�@�E�p�,0+�-��x�;����+�?=eF�F��cm(t���<���rs5�#���=.l�-����������["!��r�nw`G:�5Fm�H�*=p*�N���ln�Z�֣*=�U�}��lGb��+W��P�Z�a[3%�P��N��u5F&��U%}��+���AW-�H��ܩw-ޭ<8,���7M�\����E	T�8�I�h]����-�$2�J7�m�S`xg��MZ�5�ۙFl�[��]�ު�*�wȓB�6@`�$w�_����x@����x :F�U3�d�V������A��d8����ʹE���=���[�I47�8�>���]7IIM	(�ӉJZYG{��Ű�l�p����C�>�h���w5�x�>�^��	�#ǟ��f|a��fL�Y�ó�H/��[Uc�e�U��x )�ʣ�������l!��8gQ��<�>��u�%i�ޜ��L�·b'����i�+yIT�y��N-du�v�"��}�b�� 5M�u�C&�-HM�⮅c��yX��E�Ny�̚(��-%��wl�U�O-]�v����!x�K�ʖ��{�2��OC'ӊi?X[8�Ԫ�V�*!�[㾧w��FeU��#I�A�����.�@d���9XWt�e�
�d\�\M���u�6��!�e�˳\J5֏MU<��2��ܡt�mf8�j��������� 6tv���q��~9�Ff�Ȣ]�I��i��λf�1��+;ϯL�Ơ�;x�Iv�tl��/�ËNip�flv��)	lO&2"���Y����9�/�cLsrP���~a�S�a7�yY�mf	g:G��.s�D��n�%-e�r�qv�ߴS����a��*"M�6�ح8�T��_y>��$R�ɣ�<C5�^s+���q}]uu71��,�74n95dyi�L�n���c[G\���fA�9g�p�CLr��(7.Ш�U�����it-{Q����� ��w��p�ƺ��q�0�ĦI���=��O��	B	T�#B>�����}�G�N��J�^���A.� �hf)�.5bI�i�+�G��XB[w�)�q8^��s{���r�9u2ܽ�SSQĪZ��
~nY�`��j�m�to0�[-�VP�J�)3."��&��?Y�2�|#,hz������ǲ���:�����Y�3L�;�����1J��Z��)���(�S��m���V)G?F�m��-{�>�g�=#b��'63�)���՘!4?{��Yq�����y���`T�^�;c�G��PL�n����|]�(�-u�[W��+�(O���6�j���i#Y^LM1����u�Z��¢���gmD:�P���l2�ģ���5���iU�ך2&a�F'JˤƟ�N&/���^^9-��Г����{4|��_~�\
��s���^=����"Od&�r�P�� �=�q������&Z���5�"x9^��ס5�q6�d%5�a�Ą�3'���6_�mC	�� �ƶ�7ڇGD���&��jY���18uĪ`��b�H�U�
Z�� ɨ^Ĳm����j�e3�I��	.P����JFT�#t����MQ��P�f��F1sS�#�dK2��&��ݹ�y��<wR�"�2p4��q�<cS�g=��ͅ����kD���M�1fhu�)GS`[W؅!�#k*��rQ�;� ~ �)JR	�}�| ����@� Z3��u=��Q�s�^��g1H�t�ˏ� 3d$�A@M�4�\�q�wE'\�f�BS�/d��S�'�S�jsX9�ƉP{����*�B��hJLy������W>y�����ي�zp��.��ԪZ�Qi��5P��-V0�k�'ge��e�z!o��yT�NQB��y�7'"�������oj7����6�g
�K�X��X�u$�}M�
��A�]s�����5ɲ�Fm�\�pu��q)��tb��^��R�j:��gܺ3���#�uH�}pRY�M�����̡j���������t݊=�O�6@���Tt	20�n�4�����Kǔo'��[�,~��_�fJy=ٮZ�̛���F�Kh���6�j���v���eFl��w���
5�:ݦ�6ǒ"���on��U=O�����m(+�+��1&��+�i�"��j��g��pHD9�̑�W�{2�V�����V�C�UZ��04,�᠑4�*�"�W>�Rב!�v��!��v�/V/$�"��\O�\u�������[?y�yP��|r�BW�k�J8�����5Й��n�j��ީ��s�Cϲ���΍`�Om�QS?+�F`�N��5r���&�s��U�TF���|�J	��yn2nΣMq=�|����n�w<�����NE�f`�*jӽ��up�Z1�I�Z�ݵY�VuZRe�F����|[�}U����e��"�*�( '�� �x���n�Â7���Lς��<���/5�,ңR�dd25������.�c����呜nq�DpX��i�56񗆓ڧ������f� o6�j;KQ.3z���t{S�FH��ӰrJ~IOo�p�Г��K�W�U!&&Xc�U��M���S���t�n�Ӗ�G�r2�4�N�MHr��y]�7��Y���������}Q�q)Z�Ua�*���l�����ԅz�pl�^J+�x܉�ְ��Q�:��pTj�6���ͼ�����g�t��u����R��/���=�QI�,�y�y����EM2=�I�얣	�UE�֭�������`�=4P���\_N�3����*�n.U�V�Z�)_Sxm��5�Xt�(\ዱh��&TӾ��쵖K6 �r_�=�$��2��J/nfRtE2��{�J7c`7 �I"�|$�VgN�P�ƾ�іaK�G��P�1QnUYz�(�����sU-��]z�A5S*zs��E��1ݯ��ıJ�)��y�i�C�j�z������̙q� {ύ�Ҽ�ɦ�.��讦y�vE�\��;D���p����Ԯ�YU<>�Z�tL�ؖ�W"�wd=�ϺN�N|!���<�C�۶��m�m��
l#pi*�K�x�;)�f��j�t�ov@kkw��t>��N�i�`�����dj�����:�pW��}__�%�BHД4�(BI@���@$�� x�@�ͽ��꨺y��#�w>���|#[(*�EPHQ-��g+Xiݷ����;�-�Φ˶��n�RE!�R�oO'����-),u�uj1o���˚�>���/t圹���ʽ�w��]�1��CA�&�z��V5(1pB�择UM�\b��v�^k�D�:z����.�p�D^��)#����@���c#:t�Z�h@�nkz�\ϯ@I�-^sB]�y6��5h�޲��l�ٱ���Z�L��3kW&'�bB��.�,ǖ0�'ژN��aD��h��Olz��L���֗,�-��Y��+�4y��Pg��W��z�F*�5?<Qm�5+�gm�v(���!�M-�"wH.3^r����@fso�M�?�WsS���2�e��ѓ�לKA�x5+�qj��쒎cD����]YFt���l&s@�(2�eV�J~����V���b[�4�#'��c`�!4?�yzz&R�;)8����8�	Q&L����=�}��Up�9<�/��!�U���̚�j�S�ްܥ��Fi��ol��ػ�.e׀w�G�����z�^�W�����g�������M�.���1��c�m3�\���Y�-Kʼ��Β���-�b���=�߆����+��'�e�e<�����������"�9�b����L���vr[�5���V�g��Q�#̺�����;/�r��ڲC:Fp�Oj�:��9'qPe��ڋ��9�h�m�8r��:ur6ܳ��Y���Vpc�wF��X	�V̧:Z��&�ݖ���Y�$�@�1X���j_s]�Vڵ8��"ޥ�)Nm�C4�k��p��mڮ�G�)<�~	QÂ#FY}Sf3yPv�죱Ö�Muܕh�+9Z�;�.�L⬬�cr�e�[�9�$nk%c�Ա[Esa�̊��5�C��_ĩ��tqM�h�r�ƕ]��gNEgp:�f;�4%L�*V)eE7 ����3Gݚv������Q"�|���E�&�*2�^��t<�'<9v�$7���G��y�ѝ��sk!n���a�f�%3.��w�}�	���]o��y��&��(�˷]7��, u����4���J�x����:�n��W�5�j�w-x/)*+�y)pb��ӓ�+��a�捧��;W+�D`)nʱ�d���j�]���5�&�If�t�A\���:�.i��s2�o4Fug���[�����B��(�ER�j.�$��@�ٝB�wRa��̓9�� Wb8n�q�aS�<�q��jȓ�o17��ۺ"�Y���Q���qPR�v˩u��hѺ�*/�oK!��͚� ��ol�BC�9W�[��r9֓Gl�7\v_Kr���si��=��;�]�@[�TR���f݇QeQ	�vh	Jt�!���ʻ � ��� Q�x]U��T{[�)A�
���֘�4���q�hj����w�ٗݽ���d.+ΌX@_o2/,
E�A��	�Y)a��R�T�yk�.-��)���(�z�n�]ا�5&ѹՎ
�\� *U�ڽ���{+G6� �4@	8��]Ir�ƪÐ�Ӱ\F��w��{�a�����A�$�S������Lh�;)v���M�=�̔څ�*�J��g�
�س�&k�ݎ๵�p��_n�sWk�[�q�YԦl-ɝ�+f�VEd+��ћR��Q�7�d��A1�e������g9X�K�$�sRɫ�b]q�>n��Zs�$r��$�A�t�n�rQ�g� ZrP�E��ovN�E�w����6,%Rz��{s26��v�\5ww�'w��g�VF��U��Y�@o��Py҅U�[S֚�5���T:�n��v�Z�Me����|�\R�0(1{��3�#�[ھy([+%��:�j�>i=��7Q2�h�M-�j�DQc��1?����Ǹ�"4%N[4:���ݝ]z�Gd�T����C) ���]K����3��J���G����0s�fU�C4��$<�q�3x*�'S2��{V�v�䏠�*N/j�9���-[\���n���m1��VU.3���E�!��Į�6s�ٙ�J��r-ϳ/�KN��LIQ_�,& DS�J�� e4�d$
@ �$I�lR"���;&5�(ѷ�=m]�RPAq�k:*�&�4Um���Dl�*�����DSEQh�)�*��b��b
�4c�h�"���0E�L;�p[h�����`���QEy��QEII��U�I�֗QIDTLZ2�E4EULAlb�4�-ѬF��IS���DvƱcF��=.�T�CT�I1�������i�)��b-��H�`�:��M�X1E�C5�sEm�bh�0�<ښ)/3��Ӷ@Qk:ѬZ̳V�*�l�SED���j
�5TV�EV���`լL4[&�*��'A�����	� �Z"
Z�C����ߜ��#��r�ˣ�Wbs�{)= 	2��eLUǺkG���jX�ǳ5��L�D��+D���z�|����}�����W��I
h�� �"�a�j����V�I=5����t���_A(2_̯
���������a���L�m8UL������#�G��c�����u���H�@�e���{,�S���ؠR�Xd����Pq�|�r�%�n`��:�K��iV���mx�Um=fN?g��km=�p����m�F�>�L8��\�5�6�G%�:a���M��5O�ܤ��ެ7��~��|��X�X�2
ok�7+5=��D�(�q��'��0�I�om_c�n�|��15��\e��sI��d�a�� 'mpx�����ʷn�"���P�DAnV*e�N*-m`J��d��aζ�Zsìâ�0&�))��1P��i|���hဗ�J�\���vi�7���g��}x��-�^����9��1b�%ř��ŌaS��b�5�%���Xn���Z��*͓��ʨ���Qs��M	�S,���]�d���]�ݹ.Ya���f&�ͤ;n�^����H�,��`S�n��ס]|�F�dE�x����I|Y�!ų#Y &&���R��F�{є@J۸�"��wg|�.��آ�ٶ��.GJ�)=�B@1�+֓C`���(���gL1��ٸ%�u�M�+x��;M�j�rl�EL;���^˜�>�B�&�8>�U2��Ŷ�0i�	e���@�9��6��y�]@2# ^*�cS���	$��"� `�
X*ZJ�J����T��3]h;|8i���[(n�y�Q����|N��	1�N&g8pL0L0!�r1i.��hV��A��M?������:/�{c���E�S����1BWǟ%�S�3�2�c��{�?P���a�h��&~󀯘�tR��vd�ͯ��[)vT0�ou�s�z�h�Sbo�1�fm.���ʩ:�q0S�3�8��T����D�p<_�'��-*�@��ryNr�b���Kk��t���Qm�7�L�ؤ[>��&B�Z�ZZ��a���ƬM�����.O_��y�K���g>ے���l�m�U���[['L�H^��Д��dn�v��"��bi��7+�n����5Z�	��q}&V�OI�j��_@�X�Z�99.u�t�AM>Q�a��2v���oH�Y�k#&]:f�z���{�����)�%E��O��U��@�
�[Ol�u���O�|��8�1S�����<_�u�Vr�jnQu��{�E�ƶ�n�Q|!pł�Ki��5d,}��U���
y�1]J�t��W�B��W8�+_]mCq~X;������3j9����ͳ'n���^�>z����W��Z,��v��u7�4G���CP�]W+�>�7�vR0��y���@�h.kT��ݑ��֓5���������5o6��m�/�Ϣ�a�%'4^��eoJ���p� S�ř9�����������������((�����9}�ߟ|�.�0���;�f��#����έ������EP�*���ո���嵻���R�����.��棬��>mbTH��P+yi�:Z�_����OU�4�#r0����/:5��PˠQi�p�t�3�v�mP5p�	LU�E�s���\�%�Xs$T���5�5��c���〵��6�Yx�K5����Ơv-T1:W����X�����U'9>�ڍ���Lf�Gz�!=o���%r1[�%�̃C�]5 b)�T@S��%�*[;�w:��'����m�M��V>��aR��u{��r�i?�Ki0�b�nE�<�Jt��T����QȮ�'�j=m�z�|ъ�qX���B����{[�BU�~x�m��,�Me^Cr�75t�5/"[+L�;��_N���W�zL~5���E�Ȍ�g3�Ʀ`ޝ���=��2�Oʯ��E��"WK�'�dx����c:Q�:�N�!ߛz��V�J[n��n������9�-z����gr�킫5ž��a�v#T��>��NV_�$XVl:-���m�nQ�������z��&c|��	���&�T/�]��� �w���7	O}AjS&�ܱ�3����f�}	;3@y;6,ԻR>�Ӥ�g�'-s�[ÏL��E5���H���G�{�%!�j��������o � ����8X�F2-�I�H�LЭV�k��E���O��.+U��ᗒ7�ɗ�}�[���R�=q}r��A�J�p/�6:C4�)E���N��S.~J=���j�!6G̺�]��	z��Gޮ�G�5�?\#|�Qk�� 􅘨�*ڴ�8����^&�1N�0�*�I�*��Neڶ��g�=��H@nl,���RR3Q�˔�x���Ԫ}L֧���b��s�R5�/��.�K�U�s�FK#��v�[(*�ERB�og#�X_�a1<�_2�浪^0��m�z��IX�|�OBٮֺUړ����2��D�	��+&�n�6��)�u	eX����]	�%���c==E�\N����m�,d���h��i-�5s^pN#~�n��т8\k���m!�i��%��.�l�[�4���{4�k�V�ϰ�fܥʦ�GdU#�<��f�iF�koR&�-����T:<���G W=�X�h��xY�*ҧ��dw���&{���"��q�WdEPŗb:jZ}�e�cz������}�6���T� G���_Ct	�
�=��$��B����T�捍�����̓"����"�\�.{�RTc�~-V��k�vz�x����{l��,������H�u[ޫ��V5t�I��	O��-�P dt�ն�rۼ�8�\2�����㚂�9�(u�g�,0%ٝ��  � '���v��t��U���46"�,g��`�9M��?Oԓ�/
t�{�R�W�E*׌n�	�W.x�d=)J7m[�C��(2�"�'MÇ�WP�}��v%�C-�'���{ƶ�Y�8y��a�}���.��{�-��D�ja�lx��/_^H�ŕ��N��m��-��dw*ȶ�Y�!��{� ���׋P�Sm]�Y?a�e������,Y���m�GMG=Ӝi��+Y�{V�eҙD�1�d���5<!�5�H��E��5LX��	13�i�h�]�5x��p혢|s����M��0�ˣQ�aǱ@l����	��SףkT�V��K��\�c��p�tNJ�|`�5<�`��[u�2u�(��|	ŵ9f��m�F�>��aŖθ�3�(*��.%��E�)s�Q���"i'�INC���ת9�����bT��Wk��I/���h5��t䨌Jg��%<�e����#��ۀ�7z3��ͺ�y0�U��6���TyPFYr�2���0W�D��K��i��QkkR��`�lB�J5��g��iZ�Ɗ��\���O���z��RQC1�߬�.QZa�)h�t�q[�]��۴�L<h�^X+.hd�N��W<f�kޮ��^�w�F���� 6E�������\��4��9�t^s�s�U׮*��:]�vM=�?ɫa�G�v�2���:�k���{�Ev�W~��*��7���J	{�2��#,hz�����Rc����L=cVC�oTEPY�q�)���Gma�fNk۵C���@������G�1޹TnOD1d)�2ړ�*j1�6��K:�C����hr����cͦ�cή��Wj�]Օ'.���i��vpmA�FF6�|�@��b<���@,C�ّ��ĩ�K��|+��Bd�޵������Eى�ow�[.�P����X*)8tf����P�a`�BV�,�ۿ=���{T�bs���:��B��[�U�*�aT ١v�yf;v��=�e7d�����-�w�x�!�4��OBj=�B�m�aQ>��,�R�͏�\�g]Y`�ΘhИ�g^�D�Ȭ͇q*Pp�I�ﰕ�+���VO�Ӹ��Wx<yq�3���b�x¤�v,�:q�:�^�3��nwj,ğz����o��I�n<3D�]y@M�A�E�����ka��AU�f*���y�:�u8M�8�E6Ws�)���m�U�=1�O���
K�W��#�� ���nX��@�rή%�� }1Pؗ�e���L�Nc7��B��?`���&_�P}�V1Ե590�tS'�HO:�tڋZޗ�1|h�Q��,2]�K,]�L�mض�؜�Ƶ�̳�ҥ������<.�%�	[��Cv;mwn�~���` ������XI�a�����ÙTu�zO�@�B���g�#�o�|�lb����~ɥ�����!�����{���UG�����E�ލ3�f��QI�J�yͥ�:���F�s�{g������t�pi�8'~B�:Ԡ�8[�$3�0�'E��l7j��׶׮�u��CA�Kr0N�n��fR1�י�O[�M����͛��st�N����~/ɖk!6�"(�Vܬ�0LU�F����Cd��0)�$m٬����P>.�0��6��a�y,t]L�J:����������l�.�)�`#�l����F�8�b�pm���.�D1k�t��e�P�	�3�l��[,z]t���1��1.�M޳�6+ƪu�`h�"�D���;Ą�� �D��/*��,U�kg>���TyX-A�ͱ��JY��V�>��-��Tbt�m�"0X�Ll�ə�c����im����s ���-���b� ͌TjO���/��~*��%���i�j���%��W1hZp?�ũ��G��s�J��Gr��qgT&mx�A�!*�hբ������� � �7�ł�
��0K�n�=������r����+Ԇ����4�9b�� ���7����m�՜W��Ī+}5Z6/ߚ& 6��^J�:�
�W�5�P ʚEd�2�r�gr�H��{|r�=�kn<ӳ&U�;5�F������������������U:�Y�]t���7k�ͪ&u��fE�AO���-��/�֬�v'bv�6�O(������a�n�ݬ����?��Ǔd���ʘ��S>g�������*��u(5�`�^]�t�1�e/V���W"s|�k
j�s�:��d�N
�^�qE����n��͌�˵n��IF�_'��c�179��Z�+�9g\Ȭ��5������jI��ݛS��&+���I�>ݚ/E�hB��%�z,Ƨ�h��)>�[���z�k2��l�_o�ʞ)wv;ڬ��j�8�}�8��m���m���{9R��0����s�P����9=
��w�ׅ�Avn�9Ma�Ç3�,��c'�{��/��<�*�k���X�)��q}O�7S;����w}���ǧ�sE�̄K�0���7�L8���R|Z̝�Y�oe0���a;��� �T8�J�kL\�O7��Q���&����|��Z+?k�~�싆����3r�2;�����y�Tx�aV/K�R�{f���q��a�k\���@�[����&��������Vڬ傈̷E)��Vѕ�����"��(�w��Ă-�ϰ��j
�6F���=Z���d��ثH=�o��h����|��c͋qcr�뾧�[�xc²�A�x�S�]"���V�P��A2*\��t�f���J�Ic�� z+}�F�6*�faW�U�cց�-�����3|��S0g�����=E�C��cR�dsE�iN*�Z���[S��>�
/*d�;����c���L&S�� �i�Y��K�㱑ц�ő�����m���ݫ�<e��,��zl�Bh~�u�#�+�=�I�k[V����=Ies�>�q��X"Q+�5����E�kx����Nc����F3�kR��֒�#��|�yg�PJ���;=�b���7�i-'���iZ�f�j7K���D�W'�d�m��ǒ��iky�&�Ή�^L�=K�igTv�)��_gwj��/c�C�*7���vE2�Y�L9�vF��53�4�~��}--g��w��Sd��vb"f�bS-���"SMzԄ�@��X��X�"+���b�Fљճ��n԰�Th���d�T�����CǸ��y�3��S���.�-�onOc%�E[�;u]���w��3��-3�7iٔKmrUI��.!��ڀC`��GD��	�ES,j!�skS²�W6��QM�F��s���[*9�m:7`;3�)h-����d���E�E;�t��aV�[��#�*�y�۽�|;3�]��#�mT��:�w��!8Pҳ�a� ��z#���zw�)�%�s�8��xublGqR�w7��b�j��dB�l]Å*ǳ�N�w�]vꘕ��r�[�	��t{�S>�s��Ӳ���UU'w;�6��.�����充��1:�t���;uO�f~��J�^���>���n�nRz��+x���Yx��(���E�?%����yO������c��a��Ў ���������vZT�їz�}�AlG�3�q9Џ��[�4_��*�=��]
$w={T[sP/��S=;o�+�.�4��/|�ם6��ӽ�uM��RZ���W6��uE%ܶ0)��8��cZjE�Z��^�:v�8����?]Ay�cWx�_�e�^��}�O'���f���5NS>7����Z�"�����F���^��,��̀��v�'Ub��������ֺM����uz�@��9�x+�,g��"4�O��f-3�Z���H2��㚵UzR�T��������n�}	��B*��F�iԣ7 X��׍P�@,_��$k!14��ic�b�v47%u�O��]�I/����S�5�����叹�>���- ����&g�П���tS�.{b;c�����\��O�o�|�u�����0��^�"���7�tFZ��N��=��w����z�^�W���<���o@�oЂV��,5��}Z�Ȉ�󹯲�;+��YDj�VvvYȶ=HГ��ʈ��
0�ͱH���*����{��*����e����3�U��	 �GK��l��q_W%q��坎�ߐ9���i�j�Km�Ƥ�AS�\��C�;��Ҙv�]fU�h�̮�T}YΗ��N�T�R�@��s�"�6�{w�	��yѺ[�D���cIOs�m3A"�!�VgU��tNc�-�H�6E7V�Lշ�s�'K�W7L�Öz��gb�f�
¤Tf$6!a	���U�T#�Ӕ��o�R��
��zΥ�Z���l{�Ϭ� =��uoYx+���:U�sK9�����T�w�"B����%�x��Aи��������ɶfTѰu���+����@܏6������
�F�N��V�hd,ņ�fgc׋� R��F��)ct��6��������&�"��(��o,JH$��>r�i���c���]��m���:�_���3-�Y��
O��OC�0�1�:*V�gp�1Be>�z��5}xWo��^����b�-ZΚ���7���7,Cc-S�^�ʊ��#�嘦��%M���Ѣ��e���ӯW�v�9�6��/AF�_{��A�-{��qĪ�D��j��0�]�R��\uf�ʾYG��}5�Q�EqJޡ���<t^p��^rlP�e7a�����=����PںV7�j�]Q���"M��p��=�杀���5���VWm�b �Kz�An
���98t��.�i��4I��$�Q)��CZ�sr�n�����Vn�`*'�@틨�L��0��?e�-��W�o�ǝ�9��ނ6�)�l���I������;�[�o�bK,u��W�yL�8kz>�}uv��"P�
�Q�Vq��3vv���~,�`� �qֈwiޫW`n�&�L���mTO��F�4�e8[��ުݥ˝Y�*so�W��5-���eY�ٖ;/,���S���DM��7rIoc�)kb�R�}��+���n!�N>5�2M���Vs�/k���F��j��Qֵ����hY\���ll���߻k�p�\��u��(�H�6����������:5�<���˨z�ra4���+62�.��|D�WK��/35�����q�ej��RҐ������[)P�������޽�o�������z=��HQ.]��RJ̀�]K��mc��&�h�C�{�ګ�T��c�u�o�.	�h��;��q���ZM�ٗ�g�X�^����{[�2�5�H欥zzr5x6��v�P�tp��.%�yHi[�B��!�����Y�3�w�d.\�{T��i������Ah�6	s�����(;��F���N�bv9�Qͣ�Y����IRm]�UU�f�>�����h����أQCF�N���"�"Jb����MQTUU^Z*�*���ڼ�D�H��Ѥ�b��M�E��E-1S��ش&��`��
~Z�A��4TIZ�C�C��h4��ѣ]7,��S�=:)�(
b6��&��Jo0�@�+Al�L�G���E[.*Z�)�"��.�1%1O\^Zk˧�)h�jR��rl�J�*�|ƨ���{h�ց��%��͎�˻���\�	IE,ESQDS3�o6j��"����ɪ!�u�JK͏1�I���[8
*��Ӧ*�e)#�5u-h�ԑ���*�(:M�K�||I����>G��Q�L���� �[$gq&��M݊��ֲ�Z,��YGzA��Cr����^��p�K��J��Ԍ���4��T�{��)�`�J���<H*S2yW��J���RwOlcb��g��������S��*��yĪ`�%�f��07}F%sح���N��/�7�;\�3�plds�ӛƯz�L�n`�	����g�Re�ˊ�͐��C�e��xy����k0�3����n�=]'��)9�Ȧ�5�U�f�?���-���Д�m*ڲ�*����)�l��J�	i�Gz[_�=����B/�E��j�}B�cj<v�����=�V����I�E���nv�~�Iop�ud	m&og2��M;��)�='�~*�/B��)X�]CM���X�hbnXE�f�9��The�[�&���.ӷ����jua�{t�Ѻ���v'Tou����Z��,��ʲ�4[1Ht��m���m�4;�s��޶7�� �Jqӻ�0��{��O]g��ΕZ�����.l4�˼g�e����C8���tb�<�)�1��۰�0E"����y�=,��_(|;IA^��ǧtKxXl+Q�ވ��~?�h�y�Q��Ne%ӻ��W�J:B]S�UbZH�E^_2)�t�S��E`��;r�ij�5�'�~� �[@~��,�+�I6�� �ج֩�!�޼{z��nY�GT<�+��{�2�����Ӧ�%v���ע�˩�ku7�b��(�^3P~j>	��)���N7/�z��
���{5��Qx����Yp��顪f&y���.X��Y<���=��5'6�ax�w�3�\k�j`2��r�/�E�n��I�d��&SA�-�y8��&��۸^V�9#SN���[�Fh؅�4�����Om��xu/�{���(�+�	�{L��3����'9O�/c
�xc�J�U�]U�1��X�7=$��t�G2a��yeэ�|�CE�	̋�NJOB^��5]�%:�^i�̛k�\�5m=�#N4��t<���(A����?��%���z#��/֨{�P��Uog2��!O��	<nNֺ�wCL�	ގ���!������,�[hְ���� ���4>�r����q��}�gS}���Z���?z[u?����c?g����Z���anP����8��d�~ʾ��N^`�љymK���{��潒�`:�(8��$�V)�r�#Mu�t:O�)'�N.�|�e�����i���&�'(�|�+{'%�ԭ!���uJ<�An�)Ƃ�+\G���(��ٔ�0�����5]����e�ʛS*�X�3���M-ÎChH-�8�$=)�|Z�$��/�@�4'�꾮ѩ�u�����t����.�.�T���[�/S�*M
���*�5kL;��+�%��fM�Í0\$o���1���n,�ך��)�
�tOD�B9/���Wٓ�Y�W��֬���w�cYX�?�ُ�rU�ޱ�r��d}���8>8���#���g�;����^���2�ٍ�;�Fw#������΃����'��+W�G4;��A8;?2���x�?�w�O9<�����렒y]����,ڮai-ݥ��l��1��L��Xk9uDޘ�|]���|�4j�}e3>߶��Fq�U�%]*���������-),$-ki֡���3<����݃�_����������hp�Й�\��.���<N��-���l-1��f9 '��lz�)nbԷQ��`m�
��6g(xd���Yf/z�A1�o��r܅{v�jc��S��¡s�=W�������?���%��u�_���=*�P>��g�emF�����!Z�P	̌§��	a����eܘ�[l޶��H����)��m�\�q��o�9�c�F-���'b��r��J)�X�4��?v��#��I�c�3�s�"K���(웪��Ã�V�S�9wWhȥ�mo.���z�;"�x'�C�C�ڇ�n�V}jͰ�ӽ�&��a^��^������ֱ٬ga�l�+c2��@�+���1,��RL9�~��T烻"���8��4l�\x�(�E�&�rt�÷��Ht�i�YصE�
iMO@�Q�ېl��Wt�7)�U}	^�>~ ]����Ey�DSMK�u]75��hRm%t+�cH�J,�K`f�O��fz�C���JL�u��d2
��ƛ�r1�$���k���-2� �g5�G^W+e�1'�òjDȫ��u Z��7B�V�^
�e�|�������c>�}JVue��9��[6�sm�⪘�85��*�o4㰏M2�hJ�^ˣL��t�V�����$�߲�e������,胡�N��:`��m�U[uZ�:���P�,��%�qdl�'0͟ �q���}�/(�𴇐;�"��b��飕�兽}ϴ��~a�Q�2-�c#���C��`��s9o�{�*� E_ߏ�,)�NC��E�oH�&(A*y;'�}���q��_4�=61c��
+ `,ºj����[R�:�\C%��!����Qkk:�KPYaBN���Q��孪)�%�u�*��X�nc���	�*��R�p�l����t�����$�s_+��T��10�smU�O[��?�v�""�gtr��0��f�B��A�N�タe�1`]��U�F�{%*T���}�C��d5�Է�������E��}
B[�իjv�4�`��o8mϖҙ2��V�Q!�q����󔱚o�q<�8�ݿf�u����&ጫW1n���䧽���8���kPV�њ��LĄͳ�����i�*�����˜	��q��@}�S^�������p�M�ZD2��{w=���B���!٣�x�ߌ#��C7�*��#����E�W�g{�mJ^��y)A
u��?͜͵�P�ç7e�k]^yeYS�R�8�z�5�2�B7�n�`��Mn�(o<�
��rq����r�w��E�GW:Xy$�A�L`>�i򇆣�M�15Qo׻,�T �|��ly��I�2�\`�}˱��I*҃���F���� ��:,>@��E��5뫉�^�%5���'����@��ݸ0�UP������>��7_�IU��<�f=�Tg���k��WA��g��H���Ǻ���9O��Lx�oTA��z1~�{d�����:������h���CO���~�����vۡM��j��]������N��7�4�w��Y�V��@����`��L��囹F	��i;m�l=�^�H�]�8��K�*R��J��a(����B��V0�&����J�qCdCT�M�����͛�H]��>lc��Ka-7��.gt�1���zO�eTy�v�=O�\vӕ���EO;ً_�^ʂ�!{!������]|x��G��m��*� Ǐ���<��K����)mf�{5��	ٻK+T<��e�'0��s2�L�m�:�Żm.RpN�^a������:�"�c�p	�զĥ�k�+F��&ݴ�OtV������ݽEu��¾���;�	����@G��3�)ւB���+^���9N�7(�|���M��c6/GVe�Q�Ja6�7@�������:�2��������>uҩƗ�gOܚ�b�F�1�s�����%s�<�,�7��:Uj�F�=a8]|!�V��"(�s�O{�aR��Tw����ITB��]�b�i�f�7'�,���r��G_�c��DC�,U\?v�vS_|U��؛{F�i�}e�pOEc�y����3�ƮoipOc�q�jkPe�/X�����v;�\�`�竷�</J�H�S�f�ߖ|�j7�v~��=�3���!wW�pN�5��VV@g�[�M!ʖJ��iw�,�ӊ-;�)ɣ�y��+�Z����өo^��:{���eN�}���V�oԠ^9��O�Y�<���
��|�s��A{�T��.G*��ێ��V��g��m�e�D��*I�wL1O��ˣ���̞ө�O���!�0�v�J�s��Z��ճ�(%�P�f82����`����}�nE��Ú(wG�99J�L�LZ�����Beۆ&�wy��m����^�e-��0s��F�J����q'w��{�O����l-0dW"�������23�r�S4�u�I�e'@ \.���K����@�5�C3eK�93u�u�@b�?���N�/'����̥����@��a>�d��l �^�E'ԮD�Z��V~����F�ߴ6AQ2�mxɛ���3�a�|WZ�\��co'�����AQ[���X����H�s�hK�U�^o5_�MT���K����#� ���KQs�PoB�{i����dk;��oW�U��v�=ӧ���Vĳ�� D�z!�öj�;�\=�� �{ΩC�u�Cv�;������[R�I��ʵ��2�c��
�t�9b��&s&7�5��(L�W"o��'�����f�jL��gB��n�y�t�Ox�PjS��Ƿ��No7J��֒N��&j9�&��S���ݷ+���Buд�E�H��4e�f�sT�G^9�,�����U$(���[0�h��Vy�7�iyBJU�a��!��"dގt.V�BzY�2�RX-j�ףWF��Rޞk�XC��!#�TA,��;����4힢��	]C-)�8��t�zd�keƓU~��dNf�M�撹G�s����9��\�Sa��sǴ���)[�x�~j�mt.9�U��yiM�gJ��Fk�����F,��tNv�+��ٹ�V���:�F���-��ic�\�2V�bSU�z̖9r���`���)��lp*Y�ǰ�Ւ�{�Kɋ���]��}-܁��G�h�F���B%��Vv��h}�/�&���[�v���� 5?�*�}x�?	��S#ҹP��G�T���2�VC����m	�<�gm=�h,�=���8�++�!S�n��w���,�^����ȉ����u�sb�u��iM9c1�
��\9��qU���w��Ce KH�)M�i�4О�a�tg7��;å���Tke^q��p%�)��]�̗ H���'���v���ud8y���YP�fcnD��X�{{���w�C({R���f�w��aUM�~�"SMZ��k�]
�z��=�L�`�ȉ&͈����L��%��5�*.��/��a��*`so��x���z�O��	�Ȑ?V���ֿ[<��D�)�*S��g�vjDȮ�fN%RW�U'J�wQ��8�g���2xm�{��7��gfV�N�RÌG7bU2.WD��1Do*�a�CZTZ�]�aǱbhY����R���i�Xm'dJ'��rН0��Jn�*���I��9�^��	[=���A��߬����A�"�����d3������iW'��f����s�+-��1^����6i�A[MO������ȧ����]���v�{�^ҫ�%�A&�����yrk�T.�i�70s�TWy�=j��)��w\<�)3Zg ����q2l�:������d�1�X��?;�yJJ� �)i������8�_g��3�7���̽���������1��N"|J�On`�E<��N��vi�fyt�����V�c�,9]hs�K3s���L��ܥe����jN1�Rs���'l�g�z�F;-ô��)CQ�AL:�n��"����r�R��q�醃f��\{��U'q���Ef�}�9�7��\9��q�Fב`v�tv5��f[��۵18�Ti�h"SGC!&���\�Շu�
T�N�?:�������r�O̿�w��=n�����һ�B%��̘�I�(�Md7j��p2;^���HZ�p&�7e޽Ǩh�/9�<���i$gG�WK�Q���N���00�s�������#Ѧ]
�h��ݸмڄ@�(a�t���{��jq�]p�/�ʇ15�d�Ó����������riRve��&�!���E���
��W�LD-�t��v�U�����u�7��4�!���;�(}�aR�WsǱ�wB}Jʙ���O[��V�O��{&�l3��b0
�fq��H�#�XFS2��5{�dTʹ�wu�c�frKɶN�k爈ܗ{��-��D��]��Ǜ{֫%���ʚ/�oXю���]�������1F��M)�$]�9oe�ίl�4�󾜺NN�ΰ`ϣ�KU�u�m���9��΢wF;�V�K��|�J��u����~�nzg�~�>����l�Ab��%u�0C&�j%�m��ݷ`Y:�M����j���‗�~��'#;�*�0��7�_V;�/�=}�:��N=��):��o)��6��J�>`Q�����zu�U�:Lu^d�6��V���������3v���y�x?)EŹ�K_3�wc���"��3������k����u��oQ����px��71�q-�����gj䤳�qzO�ݺ��X��,�1f$��[N�S��e`Iʆ@��b�Z��<\\�t_�Y��泄h�jr]�ĥչ�of�v9Lc��]� �TwmH�v�o��'��Ӧ�P��fȹ�����ۅ��!��m�S���ҧ��-��#&����%�(la$kKh*?U.�˼f}�G��p�2�weW����=�6J�w�Ra�cr��E�=����vmc�j%��b؛2:y��w�X�4핥M+0�jiO����q��-8�K�cY��$�Z���j1�i�>k����E]3�Jn�Kq���&X��������[Hz��_H�Kn�fM0�f��!w�/_������}?����{�������	-�����1hLUxעYB� Voa��ͤ�u�v��h��n;��6\B��Rh��"ku��V1ugvX�푨�,��G0�
R���e�NJ������:�S�Jy7����WGU�U��V�la8C�X-r��\��::om,��F�+o��8��G�tgNA\�ks�E!���:�-�cp��4H���dM��n�Bp�79����ٿܺ���l1g-����T�-}J�^�N�\f������K���-�Uc�2��I������z�᫵��nя�+X�ﭠ�T*�Cu()ÖV��9����
���� �+q�{��ί�b���r�m33�Y��٧R���Iϴ�u��7��9�4k���"��&^>$ 3i�ܾ��S�V��{���y♞}~
�y�sl��h��%�h���F�\g&��,X.*��f�[ޝW���d�Wt"9��LC/�F���L�ĎW�� ��8��NKS����T�'S2�wRwf\��RrtN��>��j+BH8^ܾܻ,�K�Vۧeӱ�:o.1�Ӭ߶5N��5c�1��ܠݪ�aSME�sk>��pvugl��<�imYޠ&�U�p���u-r�N�/W�c�s�xY�.�/�,}�o��N�կprH�0���NE'VS�{�l��b�'bAtY�]���[�I�6�|��&f��1�k�0ˠ���%���9��:����(���\�}R��-�w�9 �(�MQ/t�ǔ��-0h�*�wjЉu�)�[ʒ�>b�d��x�L}
'��.��U�u-a���x����2��nݘp&m�J��GM�r���Xy9[�+�v�f��vr��>gP<�%�PH�m�;#x�s�9X��Qk6�=�|�FP�-]K�74��a��[���;*X�2(��S,��#@�"eU�;Iuyf�qb�`��ݭ��[�,*�����`�P=Ʈ�lSJe�f���{����_>���+vj�_�M��x�{�jli>]N�v���^����@�d"��ӣ��"�k�Et�̖���TVJ�S[�[w���ǹ��-{��$4Z�1�ٗ}�q�3Vv���_7�w9t8����$e;�۔�f#6�;5�Wm<�y�
Tc����W7�,-r�p;PedT��t%�+sP}sG"�ue�B]Պ	�R�L�-*-��}���-���|�y��/Z�wo��Y|���ud�nvdyܤ���ehI�Y)*���x	�C�#�"T�gig��)��zi�dT��=5��`3�Vʾ�e1c_Z#YXK�1ۛ,b���j�g.S�e���\
{Ĺ�8�U���&|p�Y����k�[���1�ƻu����&��fn���d����8�c؆���Y���q+�s��_��&./z,�G�8�6��q���iQs�s0ʁS�"�����JݺRi���"�$�EBh4
d�R��y��_1�f�i��� ��0�Q1Hn�WcQ�݄�M���fh-�'MW��+�)Ѫ�i-�U-%�m�AEPtѪ��αy'E�Z��G�]�����C����4�j�:덩SJō��<�y�QQ4��kS���s���4P��>`�W�h5��Ԕul=��@QUM)u��QAvtV���Bm`|��z1��[�O#/Zz��y']6�^Z��O�i�%�ڪ���_-Z��w�O�yi*��
Ӣ���:kE/@uA�8��"&��]�?]�Ɋؼ�f������'�2SI�R�kIX���M TPQ1�:�N���v�F�(�7mL�v���1U'A���:�i)�!mI�uf �w��W΁u�뽂�8{�W'ho�m�c{�V�c�f�O��烮�.����2��(u�_N�99Q��P!3}x`��������=R���Yd�~�i�0E�[N&����6wu~��xN�;�/\a�L���3�5y2{9��_ג�c���ad�l��:�zM��S�MX�P��s̡��
�r�`X��,�����*#ݭ�ځ�Z�~��;C��W/�~M��7�W?|W=�JB�ŕ|����k#vz;YT��@��d������C(y[2��-��n璄\���Vn����"{��ļ����?T��Fu���G[ȳSl+L-z�J��yՕ����5[�ʮ�N�DR����/��Vs��-f����XΔr�WU賔ɸ��\s��}Wî�M�(Z���5����oQ�Vԡ�7�4��Ai>a}%�í���X\�M�4-�cL��Jc5���N&L��s�`��Օg�V�zDځ8ޚB�nn�WI�JV�S��e��kkP��9����;e�׫���� ���))�M#�6��d�3ߙ��.=�<��YR-gT9�z�˪�nu{�Q��/!��xl��fo)�����G�s� ������
��ݧ{�X<�ߨV�]i`��"c9vk�t���Ԏ�w:��j�V��%(e��Y���`�ܟ�+R���}�a�����a��ɣ�=dU��늇Cuc�/����BJn���wn�g*�*-|���{�ݍ��'���`��#�I����v�\#W*Ӛ3�=���H�Rn\q�ۗU׷͕Ձ�� ���_t�.F�CW���>4s�'�Ta�.,Ҟa�,���0��e�Z);�0E�gR���5����Z��.�!����#J�.6��Bz#��%��Mom���=��W�x�6�j����U�����г��_�1L�t��q:�n%&26���oAz��^�]�[�5������-[�er�D��L�Y���n!�+�)ɧ�Lh�\�v�7z����6�Y���&�r��%dTtZ�L.хZ�>��f�!�@�ާ���X4��A�Y�TD��ŬdhY�mH$�501�50�* f�c�����,�1��[޶�p��|P5���:��&��e�$Y�]!��_5Y6���t^����;���.(w4g9�,d�uT�����f�:��X~}�@�J��WX� xi�i�F2�jY�o`���R��ԉ�]Y,���ܪ>:��Y{�d���H��g4�>jn��S/;��Z���p�{:�WJwhu�s�N���v�|��7����<��j�	r�ÿ����b;�DoRi#J��G���U�wj ^��e����k�v�ӝI��_���������(���P���R�W�\��јr.��`�%�೭�\�\�Ѱ6�%���rƹ�wxڎ�g(�����(lt:�^�S�O���'�S�w5Xǎ����c��6Igf������9�o'՛�R&��.�.�MR%�`iS�Ay{�fb-Q�k8�2��\.T�a~��/�U1Ns˦ۭT�*3&xM2�hJ�{.�ge����qLUUl�f�gi����r�2 �4��"��	�t�)�۽�R�cc:N���n��P{MsIl{Y���ޅ�h�Y��]�T�	��@M�Z���\w�ҮO�b��cTsu%+�ZH�|{�suY]�a�)(vt8[��XNAM�IZ�.a���%���Nޞ�b�Q*�;'0XF��G-���k3b�>L���AD�¡w(8tGol,8+m�M�8fn7�S-��KSaԪZcwF6�ؤ�Y�95�M�*[���s�������:7�xP�{����aq�]2Ƌ��Lz��Kl����u�aS �O��Z,��;T�5Vc٦]��Aî�,��p���z�7up#`eW<�f)j]\-"����0�S�/u��T���l<{6��A��ŭ��17w6狹��6�8EÛ�̻�|0>1��82���Z�G�����gu�8���aC[^5jN���=VT:c���
�5ѕ�«�@Y{��K��8������Iֺ�ڸ����ׁ�7,�R��L���tDd�[E�=���x�#�f
�X����/�C>d��F/hl�ԛ�39��f�6 �d�%φu�����.S��|bi-��x�|G/�&&�,,a��G�[�u�l{.���wJgt�Л�����r�7S�ga�(�Þa�@��Yt��3Ɍʂ�%���{�r����j��d�A(A|�ӱ&C��s��XkV���/v��l:��q�&�*a%�Kv�u�xMn؜!�9A[�Yk���=�����*�m&���/�ˆ!�sK3>(Jx:������3��ƕ�>����:��^�����ЮX��<_�3��n{�3ت����Lp��j�%7.c|#�|�ҏTU�TB�vU�Z�=q�):��򟏑��aEc�Qm��{�C�QJ�1:u��Zv�MY�u&�Ѹ��Xes�9�W���ֻ�s�T/�m��XCci��m��ޣ��=��zu�����Q�/�Q�n!���|(�gti�-a��!���['�)���\�q���e���Tz���\��;�2�&jC`:n�փ���ǋ��tWa�M=/M(}
�܎x��W+��e�Ɯv�q���bJ�VE���!f'�nY�{b+y���Ƥ�:��R4�6h`��[�J��dM���#�����Ϋ�J�x�Z�+����k�u`:���G��QVB:aڱB�
������w�f�pH��=�7���]�^�x�Z�����eXQ���!ݳ��lWa7N�d�{q�j�#E9t�m��Q9M��1��#C�?���j�2e�N��n]��+�Sy�QgJ�[D�V	�3�j�f�ȑ9�]ټ�صΟV�zO#���*��-�hOK6}\���l}*�*[��?�}5}�6[�f!���0�P�uq���%�c^��;�|��Jk���*�|���v��-SRj�.`Z�D-䉠w�0s������R9�Tf�`/n�3��L��k1��k�Q��p��r��.�JԀ��,�qG�.;іD#gcs�v>��Q��=���z����Xx�{�Ѡ{��ֳAnQ�ҽ���8F��ȉU�*&)�>�����!V+�1ϗ��Ia��-�8�3'����f�WP�<�����X�ө�-�nm'��UFs�V{z�s�K�8��w�L6�A�=M�۵Ú����8�,���eKq��Ϻ�P�ؕ���}׸�]"��LʅO�1L/�����Zέ���^K(Q�vő!���8�ƾ��*o)1\̻��d X
4���gJ#[y'�q����Nb�ִW4r�=��r�67��M�x!��N@�ŗ��nK_�o��x�
�$^E�k��Rf]I�L� �gj�R�R����:�i��D&�2��ٚ�����-��n�4�d"�g�[F�V�ۣ�F,\:!y�rBr���� TE��剚�֜�SEv\�9�`�8���_�H@�I������LWt�E�L��x�z��6�هU��M����ε�nZ�NZ��5D�#-�Kq��{N� E&ؗ�θ�P)ZB�,V�Q�Z9d
a�؂�"�u���;���W�ϳC2�&R{fRt�-}������R._^��1a�N�f���͑9���#��UfnJ'��@m�-�7K�z�L$R����U�\z&��+:~hwmSEo�1�Z�+6�YL�&9�Q����p'�{Ċ~�F\Y�<Ò2Y�0�C�z�INu�:�w�`V����Hs0�L�b�P�2�ب�@��b�	V:W����M�����u�i��17�*Cƹ;����7�g�	)�$�W3���,쮲ްN��{�`x�ںy��V���#:rWEB(拯I�mj�E��W������f�B�!��9]�N��Y���.Kt>u����]8��.(q�ktg����>1Ba�����F��`��������d�.[&�o�͞.���q�[,c�+#ژN����Cz#��b˪���lz�ƽ�=��89$۾���G���K��d�{�,��|��v���3��%n�0����44��m��l�r�X𰥍��l]_v|��p=Z�hK�{z�I±�[��Z��*��Z�� MM6�tu=��[��-�l�z17��m_�ū��߷W����V���hS*����,��h5�.(w4s��r�y�ndvM�~z׍USEX찒nX�&3��j�TF�t���*�e������i,a�th{�+���������ܪ��I���t�:-��p �Z���p�a��;�Ⱦ�f|2�?���V�۷<E:Ҋ��_ 'ZEV����^���I��5�H��)��[��+��X�L��}�X�~:P���!��.����*��f-���o���o���I� ԧ����WFR�%�y��]��ϯ���,�UL���M���"7���D�.�&�����+q��H�&�@��Pg���vv�
ZU�7���,gդk!3�l��փw�&L+�J�S�Z'b�z��f8#��Y�����8``r�"�&�/�I����"��iQO��R~mO͸����M+��eUҶޛ�X['�##�7�ٛ���meS9��M���xEUrzu�\��u��M�H[�������v'�kI��$-����t�C�7W�)�m��F�>�4Ʒ�����{��i��i�m.�<���0�3V�\T�������ٍ&z �تw�Y�ַ��I���k+���᮰ ��Al^Ʒ��ʽ�8Z�7�>�z���sjܷ�t��]r��6Pds.�:d)�K���±�i��l]���0�y���@1�CR��tl>�~��56�����f8C�jbظ�	���;�ًr]�_C.�PH�]��z��Q<cdqjb�A{�]S;�f�Mq����͝�����_�}El� Od���Z;�Y;����3;#��2;�bdv�u�+�=m��+�@k�����ك���nGL������%��e���{�9�����L���Z~1�s�3
�c�3�6׹��8�=���Ӻ�+֦x���Y�Kb?� �ݣރ`&��3��n���zw�Wp�$��lf�芮6њJy+}y#wM�M�:���ς��|�/�3�2Ҧ6�f�7mqg���@!D��HJ��n:Y�GܮyU	���c�}�Ú��MW�;C^����.kk�܌{��EaUW�X��)6�zM�&������f�۬��-���jQkL��7^��[�d�U���`��y��ju���eo�%��0��%+�����`�&�o�p��Bv���+�)V)�v^���W��&�s�a�/fg�w�����-�VN��ku+A�f���s�ْ�yR�@����v-���_U�xk	ֈ���+�<��c�3�3�y���T�]����f]��./d�Jc���4�8����W8vi��J(�9^*�tQ/a�L��Ȭ��պ�A�R[���ܪg�)������ݒ�����{c��T���f��kv�F�v��o(A8�����e�e�ޑp��&*�M���ܥ��!�y��Gzۗ.�ѻ%�y�dN~�@�~O�^��ѿ�z��E�L��?uB_��RN���K/ہ�`g��L�<�j�]DU��m�����D�{j���V��Q�Y�u�z|���CGU�xwlb�]�`�ۇ�m=�j����J�w��:,�g�uk��D�
-�w�,�V���/0OPy�3|�6�s?��������O2�,�T�C���Ş�7��3ފc�8����6:��dI��71�ï�D���vT�Nf)Q,�1zmZ�.[�������m#�:��m46%����X}��5��"Wv����y橫������2Ho~�C����j�����΋���E�)&����N7�-���-��t�(��G��Q�u@��nK��pΪz�0y�q�GΘ�O��������5�Oa3Ur6ץ�=_I�%�����;�����׌������ fd��-�
CQj���u>�ڧ���U!b{:ڏ
��u3kH��/{7�DM��v�0��g�Ȍ�ȯ�E��}�}3�AVl���TN,�3ͼ�aj�5bz��kJ[^�A@���'k�����)�3sp�ށk�S�2�Ϛ��K��HE[�[�+��R���D��׳z����ܲnr|7��j���[q�̄�H�"7�֜F��FTCa���9�.��}�$�E`���[���=xƅװ��!mTSWS���v������{�o4`�㉨i&X�&��+v�]4�/u�X�'�d3�.�e��_M�1�j�nz�;�K��p; \��@�䨚E_�ӊO����ڨ\��j$R2�gL^���{t9Ua���s�������ۣ�M�\�T�qE��j�1�����rS>K�3���c�}�W�om�a�ƨ0%(�5�����������W�����=^���x����^������h�Q2#��{\���n�5��B�8�:Js!�Q�-	�EbVw"EY-2�"�9�U�z5vXuY�Goh2���ﻐ�����-!�CP�Uɚ���췖�jo�a[Kt�M4V4���=�	ǫ�(.��̻���-�z�*F�9�L�3�t�.����c���d�4���-�:��
�0S��c
1�{��K7c�����W����#�^��	�a�pfryiu�o]��+���(Mr�f�/-#���R���KEk�Q�]���l�@�ځ4sp)0*S`�\*��sS�2�#L�2�Pz�q�R�zZKr\S���[��vѣV��4Pe�|�|޾k5�b�V���(�I��4�ɰ�/f��Z�r��W�P&�ϼ+\�=���r����.BO&��8��J2�U������L�I9����8������ˮ�	���V(�4�YҲ�u5O�=�ر^V��v�P�0�X�6IM��-u���v*ζ��@���u!�#
����W�<�@��;\�55����Z*�Ԗ�(1��zN��_s8$�5��|:	XØb��5g�r��Tݲ���X6�q�귩4�tΐY���7y\1_�(�Z�pZ���,.ۻ��,��*�6��E�6^m2g٫O������q�]*Dྩ(��%j2&b��� eNh�\v�c�Yk���q
fZ��p�L�P�n%A�'c&�F����ܤ�4\Y�A��(��(�O�w�:r!��� ���rLt� �Fn�m+xl��#/�+F�kyx@���5c�D*�sm��5�Vҝ|.A�N��&��qP��s+#V��o�x��{6���c@��&�7ɝךJ��+kb�K�t�y�r����WKu:��T�I*zV�s�&(.�ݽ\����aK�Z����L���Cm�疑�rZ�(wQ���5�DB�d��wz�w��O��z3I��f��/�k�7���.�M!��r�i%���9qL�g+@�;�G-����As�t��0�F��)m�;eJs��,˴0Q�$9�Jͮ0�h�S�����e75��L�f�%��j�uFĨd���UX�f�Zu��kT�:�%�K�m��p� ��6�`�����ptꂵf����PW�l�V%�V����r�I��g��0M��!�a�ĺ������	JZ�XR'nLX7QV������e���]�踯H�&T�x�ثK��QM��pA���}��4��Rlr�\�P&ɴF�ɎՀ_q�S��$ň�ל����qt��ʲ^v���<!Ut�*Wl"]b�r�����<o���4�̇A�;hG���wLI=\n�f��AְR���3�'#<ǲ�u,��;���dS���u��R�M��Փ�Y��n,ڷ;�Zn�2�^�vzM���a�-;��!��q8��[n�YW��h̜�oX�6r�v�/�a�'�'n'%G�w|�Mɛl����*���v��bB$���*���UDUL��d��Lɶ
ъ�CF�5�(-���b��cAMD᎚x����ъ�AN��::���N��Z�AM�sI�y�J;X�N �:֓ki�6�%�h
�&������"(4ETt���&6���h(�G�CF"TS۸5N�(�kK��ki4tn�1.�v��V�j��U�J(��yݻ��Z-�-�0kKAy�tQV2h
�-&�E�6�M�:'_'��*[8;��lF�4'GOZ)i�=[U��]���ƪ�$Ck��ۧ���l��t3=`��GDí:
{u��l�tWE���m��km����cV����sˮ���ڝ�O'^Ty�M�]�Wa�G%��JN�X���6�Zf
1��1`ӧM���8��#�<ڣlmlh�4��t^d�+N#K�V�4U[[Jm��A���$h 
5��;��Rݕ�쁝{��G9Ҿ���m�����=`���ί%��x-�0��M��Cfќ��,l���U}�\�l��R�}U��<u�����7��,��#Q�[q��
��aIV17
Ȱ�|ܣ8f��u�M���e��pc��5��Xj끷�Y*�Ƹ�<�"���l(;M���I�j�j��'mm|N8�7��-����3ae���,�۳9H�����:ݍE��t��T���S��s�s�ɖi(ehL��VNT^D'��A��Zf�׋G=�'���-ŴV�~�5\��9�ncU0����*{q(I>�Xݺj`תc��7W}̜���bAH)�N)�r�1Kt�e�hx.�l��]���<�k���R�i���M�Olٴ��E�f�Qq��;dDO#��N�i�|�@��/wʥ��>_�A�=\k/G�{@bNnG�Rv�Z��W�����l�]��Ep��T��c����Bڿ���-�{�=V���r�Б���Kg$�"afH�~����R��S���$���M��m��W��Z��;��������b�vG�<�q���tl\�|6ͅ��q��T�ݽk���c����"�����(��M��<&0tl�:�ޏ�2RN�	Y��ѳˋ�X�$!��R�\\o��^7��;�bN���^u�z:eu��vr��������=k�$�G���	g��K���A*Z��٥Y�1"�`�;y���ѐX�m�
�g��������ٔo̸�6�Ә�k�	�޹n��}���Q��'z� qf e�5T>{�죹�#I��y�L�q�2�-���ENz^�i/T�oj��a���ʷǮQ�K�3��	<�n��K__[�h}'LHүI��Z��.���w6F�C��q@naֱx����5V�j^�1�U]�e��A�� q��-M�����7�	��3���1s�}{���>Ǐ��wb�'�h�>��6���7��E_(�5�˽�(+v���yўh�`����Ų��z��i{0̊�k���X�M<�Y��ݞp�]���:��1�;z/dK�?m�P�p�Y=���/ö/�h*�����:�lL���|�!(���_x�.���>5� ��r�@����Ի]-:�(�/@02�ZX�TϞ}ԁ.n�E�S��I��=R�m0��Я�˾Fb۾T�!�ɿ��2�vѤ�z��N��ˍ��
�����c4T����sy#VJ$fJȓg`^�mPn��չ1��h��ڳ��j��y	��Nu�z^ԕ�)�������]K%+v�ʝv��hx��Y�.|T�x�t�)�����P��k?��'���O���P}�I����2xջ�KY�>zזb��+fm�ȥ/�M=\�&.r�ҫ�	ޏTL{Y^�@��m�r�+*�ۊ���W�8�S�&���~��,��W��+�z�􌎕��d�3��i����Ύ�X���ߺ}��|)���{���㪚�)�WK:�G8LAt�������y�R��m��x�;���?��2$UZ�)��Y��?�^���1H����ߴ�#��1H��n�������Q>3�y��#Ll�4�T�R�8����><��#������R�|��
6Ŵ[dܲ����o�?���1��f��2:����f�R��x��P���w�d^
vDl4d�\Wu��!�Z�uLaN�Ϸ���XV�{��rα�щ��|�·O��V������jv�����{eX���^1���p��kݧ�6VWU�4��*i̦�̦����@c����ֺ�q��Z�eԐd��\����yw2�f�s�.�'G2���ԖJ#w�_fu��e��(���ܒ���L�2�n �6�����ɟ);Ƴ�]uaDF6�s�yԙ��/��'�g��s#���`�� 6(p������ٔ���x�e�蜘�=���1$���c�0$����	Q�����*V�oN�k�J�Z�C�4�G� b�noF9�+F�)Bz�pյ�M�E�;kq(����u}��91�E�i�����e�L�>��-�6�fN	i���k�>���^)M����ܗ���ȍ����t�,֑���x(c 1KF�^K���Խ����h;v����7p*����@�p�5�th����P���̧����#��Y�[��u���0�fA���:_s���gZ���Ksh)��v�@�e��6�9M�,������#�<ul���n*2o��0gL�	K����Us��$=[�f?�f��lN j��e��E�F���u`vc�q��R�B�v��rrKh��]�N;s�mAW/�>\��d�c��l^��ޛ=2�&T��������;���k���S{��5kU��M��Ov�T��Y[6�e�i��J���RJ3��/t��V<�~UfΛ�l�������M �y�%^FN�WM#�B�O�*�}P�M>���h���ӧn69�YU��Au��/>y���"���Ź����0��ֵ�`u�rx��Cc�l����޷V:����;Ե$N��6�������̬��L�/E%Nd�3ݽ~��wK��m$�[����o\Q����&���Sc�ob������xf�|��h�(m�I�a�gMј:��3g�I.Ӷ����7��;O��״qa�<]֨���n��[��Fz2g�K�d��*���H�Z���5��=��\i="%�-���q4��	�׀�z�`�}�g�݇�Qm�� �S�P�:��+��T}�NeJ���h�g<B�hNB�X�����H������a���{�Y�R�I��W}g4�BWh�x�V/���&�I��7z Te�S
�N[U�;�f6c�n�k����EK�@q���s2Tfr2���}h�·R�w�^��>e4��e� Ry{���g�F��q1o4J�s�T-k�[r����֚��93�]�9ż�T�;���oPah&;���j��t�78/t˰S}O���6�z��c���S���2l��d�)��i۬���"��حG$%rkڭ�֩��Qk�nU =ɼޤ�^n�C�kz��чkz�<�;#���S�Pr��j�oMDWRP/ݔȱ�B5��P첅��ZS��8^�)<yҾ	IT�p��ժ*q�Ju=wp*u�u�ض��g]U���5��:�3���pԸs�\tvd�E�Gr`A2t�3vڻ�R��O��,��Š>�+T^o3H䌆姁$�C�::dT�dWa~�3�����R�+�+%80i��w���Dpا1��݊�d�Ɋ����Xq��{I��c�k�2@%_Q�g�e�D>������Fv�t2�η��l�L����KM �a�j�ul�t56l�����!*�'"Fv�2���ly�'Gr��nw���7�z�'ܧg�S@�m���n�?W�7����VFF��xa����V_���yo���؊oC!�E�����o-���J���l�<t��2��R��5�7�r����or�`j�5�i+���m�boi̜� Z�S��}�8�k9m%3�V{@�{P��'Q�!h�����m]=�̺�`�C�U�Q�� �p5�O?�}��������?zj�0�W�i�NϜ�yöP�Qx6��* >o��[��#�a��U�3o4���Q�J1�\�U,�;Yg�6�{qI���ە�)�����go`ý�h�ʎ};wY�݊�2q���ܤ�x�E�Ս��/|�!(��rt�5�l|$��1�����CADY��C�Ql�\���͖P%H���7�Z-E�Í���;��%T��20���(II�e:^�n�dwh;����/*�p�ݓ>��WBc���a7>��yB��B�*�
�֝�-Q�w�ϔcv��Ɔwr
c�=���h�%���*�Զ��޺��yD-%lZ�?z���H�Ͻ9�>ǏU��t�S�ӣ��u>�LO5�[�2����y��I��k(���wj|هҦ�A`W�g�x]���.��˹�.I˰Y��rf"t���V��^���ԼO"���7���-c{�nc9�8��Ֆ� ���1���HO�˻4F�bz���jI�v(&�<���!u�\R&ذ����u����!��r���5z��6Y�+�;D7h����z�Oq4ܑVJݿr��sF%m���KO.���y�#��{d��J���[G��ޕ��IIE�o+ߧ<.�p=��9��z���8n��"����UWa14k<��S�����S�.�V�wy�R��'�c��᧔�<�Q�O>�i��VR�u ���QkL1�
w�x�F��gf��2z=^���|�?j=��tq���g�ȁyoY���Gt����<V�����|;�`!H��5��ɜ����۬��/U"M^�
�I���ݝ��9��~���1 ��"��%S��>d�Q`�#��T���{t�S��������56�AG�{�c溷FN�j�ɾ��Zf���y��7`��Py�f� �����r�Sb3W�B��ؓ��{���~�QV�o�����{�^}XN�(r��yN?��fr������R2ڤeM�7׮uaR��<�!�sE��FL��	g6�!5�V};c�<�,�5�$��+���'�x��	�F��w~��;�2(��O/3�]��5�9�Z�-Uz_p���^�}:����\[��HvƧ-s��"�^�`���Wyp�c����A%�τ)�.47U6Wg?&���MN��<�%���D�&������jy��G���Ã&��T��).�b��*�%WTr�^2�w�Y>����ls�F�[��Ot�͞�s��).Y8�U�+{�Vě���>^��Œ�n�x�c���.���E��VSrG�J��;��o*	̗���5	�[Zv��[��]K_Gv�i��fw��	���;X�w�A�-����f��C�Ҩ唈֐w�]N#V�d{Q�z8t�]�KXAA3�M�וy��^S�Q �R��hf���=��x�����ң2�'y���wq=�''��svI���,�&%kSmq�v��n-���bic%�i�[(�T��ro��v.K�0ezJ7��*��d��r&���`h�X�8I�L©X�9�p�k0�j�FB-�~�v���5�2���2X��BʋPfP[ҳ�hֵ������s�7%ie�$%5���έ�V=�I��Y�c�Bj6ޕ)O�IW������e�}i%���	�þ@�;�ԁL[XK����0��5�md��;&�$6�`��l�cL����ӻ�5�0eG^VP;�cc�h�j� @�R,Z=��7u���� ����iҫuP�6�[�W��N9-�|�h��p�QSb�=ٍ���@�[M+�����E��kM-��,2���Z�c^��[���
����"!]�1��~-�n���9�9e�81Y{eچ�u��s�d&=\��o���Ub;�1�li�A=2+��I)m�����;�5{�nT*��3B���x��2��xǴ��t��9C�"���6�x�W{mL
�,�.h�cu57w1Xr4�$��������5ɽy ��KO+:B�hgx���YE�v�ð缀����Inp[�_R��tVU.�8��F����o�L��-uVy�wA~�X���e��{�����?�������z�^?�����>���uN;1�[䭗�:gA1��Tz*�`��^���^��=S�[�-ӈ�ۻ�5ʸ�k�x�79u��b �N�̭�XI����m�:Ygy�c(S�+������#���������sP�D�v���YNT�����̊�����'H�E���j���ۨ���Xsic�k���g\t��1\�d=��\�cqM���eG��d�8u�*n>w�u��)p��B�80�t/p��l�Ixr/�&gur�Q�gF�|饽�w��lQ[��8^|�B*���'R8U�,�Lu�:���﹒)���)���m]Iu(��\7+7�FZ��9:,{3`ˏ�Ʋ��E�x4�䭵�-L�XT�Y�q���,Ѳ	8�B򼃵�ͷJ�*.;�i5[[��7�K4'��N�suc+j^�s%��h\��h[�7�gD�	ZHbyU�s��>U' �<�J�����Ho]J�l\Z���i�'&�{���]�e�Dɹ�2=��J�y��gI�`�ki-�P9}@��+s~���]Ef�"2�cT�6h��a�84F�a�u�A��F]C ˂�� �o� �V7�V�u<�r�ֶ���7�R[q6]̫�޳+r�Q�M���:��"q��P�N�Jh{�d%���5e��r�rW�sH�<�jq��-٥��1R��9w��Ť*��o1-�h������VE :4VaCi�����|&[*��Ͷ��m�{a�l���3H���m\�$^|d�5uv����"M������2�9���pNڅyt*������l$����3N�'�u�Ȗ��@��s��K/hb�+:-�q�����Ik#��
�Ҷ.��(��X���!�"�+��܃'��*'�&�Ku��-�������]#r��ʶ�:�e���Wj�
<��K�cy��!2,��7K2�X:���y�N���W]�Z�:�(�Ӯ�X����g���:��%8�f�c�P���x�5�v\R��Cy�t6vL�߬8�,�m_XX"���/:ķM
�%^�*����D�t�X7�^lr�������\�[���v\&��+kkn�j������F��w9Z^ޅ���J�e���Gi���Y��8�5�.����@��Xp�Z@�9I��{$�IF��au��us��㙂�u"�-�k���v࿉ٸB�a�+�MuDќ.��3*���[��2��o��ޛ�pgD�ax�t}B�=��c�;��M���'���R���L�r��P�	%�ٜ�.�YNb"Ÿ�A��Y>�dHx�]�S@��n�Z���_e��,
\��Mٚ��hPviu�G�,0h/�`�(���8+�v �˫��c�;W6*pwI��n�-J�Kj�f2���e[F0"�!��}�m��-vG\0���Vq��X�r���bv�0^P9��l�Ӻ����λw�ۨ���/:�x�ǞV��~��gQ|�n㘚:+���i�mlk�ښ����&#�ڴ��F�Kb5P˪�Ƅ��#AA��Mhh)���)�ӻ��)h4�m[kZ��ct�h�5y���Ԛ
��y��n�|�h�#��
�m��f�;k�uA��U��Y��xbƦ�h������@Q��j��^kNي��F	{b#�ȚN�l�v8��A��kTV�lV�
�li"�h4�m���Vq��).�1A��M�ƚ����ٰ���
(�II��E���ȱ��bѣl8�آ���ƪ�|��E�km[m�5�i�b���EE�3��ų�1j(1�!���(���m�y�tmX�����u�gεb1i6���h4�N�^y�͓Vڪ(��63li2E�)��U�AVə������)�Yٵj����M;n���h<ڈ���6��CT1[:.��~�C�>��g��
�{F?�(�Yݫ.�jV��Z�"\tT�K|P�ܽ!fex)�&��������L�\̮߬��d�Cj5'4I&�Z���,����?�c;��|{�%���Ĕ���o�l��[D�Ĩ֍Pj�(,��ȫ�d���i*^��,��{�0�\u��va�}��cc��y�{Z���S"�ɚ�/�����	w,O�C��׉�u�ѹFy��r.[�s�4dՓ�s�Q4�lΟ;�����C�5֞���-LGWN�u����p��`�jI��2.Tli�n����W*�y�d�4��C|������FY�!/.��O��v���p@Xs0�u���ɤL�/�s�ac׳���V6:C�	�:�~En�;��(ؤvպ��6��s�6W���%�G�Uv�]6ƹ�joĻ����"�(�[�k):��gue�d��Z
 �<�'�[�w�����V<\i.�>˞W��z	����oqD�M���:GY
$#�jj���Q�]~���
����$���my�=��m�����6���3zo9�eq���I�y�^^�Gc'�]��Ĩ�t��ַQW�LBK��w7J�{�1��q�-��ӂw=��_J��j4�v��7`	X�T��u���7َSǳ�9�ͼ����3����u@�5:�O����,��j��f�j�����]�������&]0�r��7F�ꔫ�����ܑh�i�;Z/�7�H�otGO��r�9V�3-яV�i�BB+������v�N��}97� ��Gsfo&~�Oi�f�h���L�n��j��eh�T{"9F]�K��WƟ��xG�o��E)Xl��슏5e7E�'QT]A|ʦ�N�n�0Dp�7l�mrͅ���ήS܌�:��:�����q٘�r����[?�"xȸݴ�;	��$�q�е �sh�M�{���h�A9�z&I������g�L:���V��u�Uuc1v��oO.��Uv�O�}�G��6�{z�Џv,�ۧ�Y��NtI/5k,k�h{Ӥ������V�uz6n4�|}�c��ƇG�F`���>+��ނ)�2$ݳ�Ew��z+fM�S�+�͂�G�|�=H�B���5^	.�+�X�@��,ٿc�=P$T��_l�ҭ�����9�Y��!KN�Z�������	�v7�U�հ7��V*����Ǵ��F+��:�$��km�T��G�{b��>��|}���{e�Z$�7���{N�3Do�q�'��9O��W��v�ol^na��(���#x�qm���aѓ#�T*P�ZJ�ȧO.�6D��5yRnKU�ޫ6�n�m����[H%!�j�%B"]��^������vG<BK���?�[8�{�3�L��Ԛ�V_ެ�[�ι�	�̚�S����t+����Uh|4�1=>���V�y�+���xDݍ�	�ޘ�6��c�t��j�ˀ��j��<�z�t�,#O�j���e�EmZ��e�WT�e ^2釻�V��RРS���xk�;U�@�q����poB9dߒ��׽���U�"���ɧ^�~���ګ��~z���-y.� Gv��{����&�1�h��rK����oyC���M���c%���a���#4p="��h��H��'��绅=87��o�=�bq��P��iW,����ܼ�͏0� kV��N�}HEk�Ty�Aj�)�Gg��y	�s�b� �04󻔣�:�^�f=?v�<�K3m]�[��f=��ztw�������t|'b�aC6gWYca�{v��hM�����O�V���;0��g�����qS"���f�VVe$��V�1��o�Q�z����-�>[�q�4�E�K%��۰�Q$��Vk��WyS���\�
�W������E �`��RΪ�}�.�J�qՔ�ʹ_�(���{����Zޓ�?U����N��i����P6O�v�:rہ��18d>�\���p�nv��,^ӛSY�r�ӫ`~�=���#Kb�yٓU7p����ͮz�{!�@n[�Zf3�7оH��oa]�\�;���w�<;����n�.���P��<O���$��,�?A�ۏ�������i܂V�R$g��i�0�%��[���jos� 3�������I���[��j�z��B�▕Qx5[^*��*i̊���v��8*~3�ף��!��t��K�F1��
��/	[D���ȜOo����$N����3�:*F��m_=���T�t�},!���Y�1�	�1��ӂ��lF�]�'}Z��.^�3���5S�v���2��t�GN�eG[�Γt[��D�ީe)A���C���F����}1��.��e��F�k6�u���VI���1q����r
iA��8�M�V�]�>	���:g[�U��l�
�2�=�V���uk�l��c�]�+�d�"��`��e^�۽t�Ȑ����0��P8���p�؈�9�&��Զڤ�FM��L���U�U�5���̙g�s��#�f�,�u?�_0��Hc:��m)������e�����ew$�j�8���-���w<yީ]\�D�:�����k��%�a0�J�@2�49�$�}@�����UN�q�N1سٯ$f�B �lm��6�0�)���Z��e����~���<���_�0��ޥ�)������\��c:���g��h��z��L	7uu7���U��$�A�=��G�&�1Fc��J�ӠKwr���9�\^�0��ק쉉������H���k��t���B�vw{}_�c�_���
��?K���<j��:%V"��i�ym�����j_��0�|' �(�n�}������K/��/	�N�շT�4�}`�c�3����YX̕�)��oc���H�D�/���9�\oc5v�ՓRh�-VX���q%��w��6\f�:��,ȶ5�� W�7N;Oo(�:|�Y-���5���S�	6z��e�G�T��zt�j��V*ƺ$�X�l���^�o�&;�u�h�S�����4�(�<��%n�3�v
�2S�L�����:\���o}�ף	�s")_	�;p�%
�
�W����wi���c�ܴg��dV�\�с��W�*_WW�V�i3��>���>􌀱���Wƛ�ӻ��>&�������--�1��׏�l~�5�۩_FV���P��܋���Z�\�V�*�l�:s���7{�c|F�8��J����;��͎��ɾH:)�^�{���Qqklr�n�x���b�����[�&j�n��"�h U�	ǥ�.W�2�l�+��Fxwvo��5Ŷ��r�k{�"kMs��m���w�q%���{�_�������+"�S�������O+�g��S��|i��C�v��%�XMl#1��Q԰�AN��:��3SWO4�f�:��´���:7�?^��k�NXV���,1��q��4:m���8�ylsE��elo�\m�y��90�b�U[2��ʱ�L.3q�=��v�2_�)PK4�^�ڽ��M���n�}r>I���nmBޘ���=�zk<���YC	�mz��/7}���^��gGoVm�7C,�0	���8؍��|�\�̞�����jI��ueyg>�)��s�ݐ`�a����T��z��x=�`��d�,Ma���:bN4��c�e"NZZ��^���p��P�V�{�-����^�O�؄M7s�����*m�n1���r���唘���^�����83 ����益��ȴ�f'�kTL�N����7�n�渭�0*W�M���Ny&�/|\��J��6�Z���;�z**D�qS��n�Ɵ��ߜ�*k�rf: LN����\"��{�g���>$�(��MM�Ê�;Ǻ[`4�7i�>e<��Y�V�����p�q1vr��#�P�C��B�T�5K8vs��t�b�V~{��O�����z'��å�Lma���\��/6��L��ǜ�λ����C�IܲK�S+^�p��j�Q���z_1����T�p��&^��GL4���V���1��+^���i:���J��岏^2�l˂�ɯR][5B�xwGT�??s�A�֦�9��)hB����UD4_`�r�4ͬ��×��{{�W��|�a.sM�H��j2wl(��0�^��U�8����^���h��틫�{�*�@�w����T[.`���U��Uz&h���N�=j��hm�f��&^�\hl(6\Z��"�Xl=�2�wzU���uPX�Gc�T��j�x���!��ݏ�n-7��m]�C�m�k�ZWa%��wiw�EkCm��s`��kQ������i��p)�ܪ1�ё���,�ܫi������$�=vS8f�V�T�ޮ��:�u! �H��ʱ>��[�rX�B:�`�z�<�����1��;��96�LSm���ؾ�Y�݇�Qc��W7zW~���9m�I�_�F+�o�G\���W�u�K}��맾PEG�!Gܻ����)��thqciRU��I���_.��+:��畝�D�ǔ�yL�ޢ��|�V"}��OiBbZ�(��diN��Պ�71#�f>������$�n�@�o
ns2�ɨqn���ٷ�6#:r��u�B�1eM����{����q�����6���=�c���V띶��p�ɡ	\��6����ב3�3z�77��4=1#�r�)E���v�i�S���4rH�kN)��Б�a]]��{h(�K�{�Y�xR�K���ި��gQ���۳z�K�u&��U�в�܂�Pr���]~+6��.ӫ��ʥ���!�߆ؙ,��>�`�CЕọ�<�|
��fm��S���'rc'�i!ݏ���`�-R=���[���a���"!���7�_I���3�W��*�9�;*o{��jCT�)��,�W�Sft��5����2o#��{#����6ͪ� �|䭿�r�]�B�:��ȮW�yw����S��s�<�0�eW�3'���z�Ȱ�0<����a�Zl���(*�*T���z,�fepJ�3�<|�C���,!��0]�jƙ5�2VDa�o�t���Sy��f#�;�|2Ne�:�v���36��S-u�>�m�Sn��Y�\��#�,�e0f��_N�R�ݒةh��'���}����>��3 6���%�֌+gk˶�[FpoP~su�Q��)��|$;j]1�L�li��U�n&�B���sKedf&ZRwvm�zk�O�S�@wj�ٗQ��k�݇&�f:�K�ǭ3NoLE���[d��4��o�<˹���Ϯ�ɜ�1����F����Y��iG�\�H�Z��R�:0����9�ZFM��g����܎dg,m�&����H/N�l6)�����'3�VY�X�v��n3���u�/9�ZJ"��,��XgB힔WR/7*̆O��ٹ6̅ix��*�����)_H§�v�|�)E���z������Ș��jy�(�<���A�L���t��D����p{vF햑��x�g3{d��	q�@e�@�M�^��~+�z����W������z�^�W�����������x��xl�e����: ��͌��˔�@�t����t�ŝ2Txh7yu���<�����o{jW�HJM�H�ө�K�@�������{������?<�o\#�%M
D̔�g\[�r�]�h[=�%�����ϳ('�\����mmG�s3��X�[��H#{r��ŭ5�I�Vح�{��ue��n�����I�՝D��XcMde���2�LE�wEm�2ky{�C�B��W�'�i�Y�6V��XkN��A$X}����\�L�3�ɺ{n�=xM�'2���8�Q>v+.�TB��ii"�����}�ҩ�o'��8=r5s��j]�sDS�{n�ei�쪶}vb �Z��VL���7y�O�������a�z�V���@���8-U���z�ܴҋs���c�cnH�t|�5ݝ�"�S.Y7.Rӵ��X��犅I��`v�s�&�M���TZ@�z��?�+� ։C1��`X��Eg��.�<���͜U��0tVS�Ӷd�!\ �ŉ���{��� J���2����0)ۣ�R���/k��#Vb��e����kk�n���y�$]��Zn��̈́6gK˥ѳ��Fm�i9�2��][N<a���6�%�J1�+I�
�W]�?�u��s�	T�*��8#S//��D�#e��0�X+���*�l:�����4�,.�D%n��� a� �y�휟K�Q�R1\;r�b�-�MZ̜mm]��Y �7y��Wrә9R�k�ʅ����@o��/��Ӛ�hƛږ�1�#1�I�kskX��&R��9W��Lf�_Z��0�J�#h`��N/��z�8>�(���e���+�u����8b��u�ФO�5��k��fF��=���ɔ`����Wj�⥾"k����kK�MV� q:FSɘ�:�A�9u/5=�9O&'�f�,ôu�R�\Ϲ^S���R�嗗{l���9�aC�q�륆#3tQ�����0�_P�g,ܩ]�j����w�,��Ź�bFg<�`��ve�u��f���K���^�����є��ΗD�����|iP_�iݞ��cs)L�/՞�F�k�#F�Ml�L���wWYȆbV����b��^pw͓�����B�0����>᭲�C&V�]3t��>5ӷpw49Rɡ�,U�-�x��SxDqd���D�����x)&��N-�/����K�Q�D��7E�����K)�\�¹��J���j�:��ǎ�M�]OP����T�}�e�\������*��}���+�@�ܣ>I
q�ܮ�)�b�T��#�u�"V���;|4M����+b�3:�od:ѭz�ﻳE����F�=�E[�܃3��5�w�C{�j�q����8��B���!ؾ� uh�go�����|JrW3�i�f<�2��v�06m:*��B��i:���{r��9p�ئ^)�wvx�%"$ �H ���v����U�^wt�����A��8�]���4��je�7v�F��L�cIt�"��"���l���cV��Ma�:�=&�m1��QE�TF�����=bN��ϑ^v�8���:�+��熻u[��r��٭h�SF�%UQ��ъ��Ӫ
���UlQ����61V��m-QV�A�u��cUZ�m6-���m�����-�[b��F�[X(�V�v�ڈ�����b��l��b��Q�i4�5T��G��u��gin�K$ڵm�F'8ѬE5ZmlZ�E���j-d��b"��z��֨�tc�Mj�IThmF��lkZ�3�2�S,Zum����"+N/.��my��i�y���\c3UT��S�i�6tMӦ.�l��8�ƷϘ�-��6�*��LQ���Χ���[Ry8���,R^Z��݂(�m��C�K8/wt��L�~udKH��w��c舷�x���x�]���xo[���q��wtvT��X)5����jS�LcF��v5��������o�zh��ӳ���⭖σ�Mr ��P�nn�o�yON=�')�AtoK���M��~A�dդ�Xϗa�������V���G�d7����+k��l�n��+�*:�cF�v�xsQ7UN������@����#�}�*o��ۙ˝q+�u�oKn&��S�����U<��`znC,N˯иȸ���U^�&$
4�cjm��*{�S��K�_O|���&|f|X�[����6��U�^�L�]=VCD���]V�l�q���	�{����=x�PF���/���Ţ�� �Ȩ� =>��d򵝑��5=����6��.:�?�i<lr�5�a[dz�r�]���-�I�8�c#�<��G,�ђ�>|A}�w�O˞��>���"�d@��#;��8�E�H6���w����&�y��g���9�����.��y[�X�W���N��T_!��V�:rն�d�7<kFe$�2p�4j�q�5�L1]��?N�V�洹��y�t�
��N� .U���gJ�F�G�+��֠�d��Vb������P��{M�Z&v�\}E�y�V���7ʆ]��-�
A!NS�M�^�f�޳�ր}���/ө�O�6�YW��\��ys!��UQH���zpD�i6=�ܝ��9E��v�T�a�˜����R#��}x�3���v|����x=X۔w��׏\U=XmUX���:[c�T9u^�W/�K�2�ů�^�ö}�O+���"�T��/$WTe�ݧP�n�[J�ً�ͫ����[�3,��Zm�2�$��Hqoǋ��n��I<�$�xX���U-q���"���%�u�K�>�*��^�z�$8���1����cu�Iܾ^���K�Y1�t���[���u��F�4�ieYy|[�����iHn�X|r���/�)knH�Xv#�KPCO���3�����'������FL�C��.G�[�P�B�d�ώ��AӹS�s�}w��-�[��7��=3��y����t��[�Q��]ױ�n���v^"ܔ:�ԛ;smb��f*����l7;�8��4_�f����쪔�:�UC� óǷֵ� ��t�F-*:S˻^�E���H�{F�L6�-Q]�Z���� ��]�~��_�.��E(�+�3�wVYF֖���/C�N>*{��u2j���@���C�j��M����z/9TwR��z�$��G&��/~�!��N��8r��>�c*�{ad�j�M�h����/3q��i����M<1H~����q�ĶٱY��_���^��%�נ�=��~1��]��b9_�Ou���Py �_O��"�,3�Gz�H�ͻ{]��nC�0U�3Ғo�»q��"C{68�t�|cw�ML信<D��G�^f:�n��y�3�v�W�����-q��i��e���*)��ߢ3V2w����s/��������XĦv�Q ��*��jƁj�Ƭh�~��1�{�����Լ���Z��#"L�t��	PMq��v7uaw],��75�^��i=���������I�K��8�t����~C�-�\w�T����n��y[lR�IU���+�jc��X��K_n���fĹs7�t��L'3h���4�Phr��g/2�Z�p����u:�t���5���������_k)�v��R�F����׵m���q�\�5�\�wȃ7&b8�d~�箹?ʽ�q�g�PF��8l��!�\��*I
�yU��H���9�RJ�s9�Z���w�7R�d�`�M,Bc�1�#��)�!M@u��2đˏ2qY]Ғ��E������	�>Rπ�"�f=��QiՋ�E��J���/Er�Yǟ/<J�<�uW'�ʷ၁��pf���#_�_����mL��qN�%ܲ��2��v̝�7��ײ��y3{v|�����#Q����޻���r@ �Ǻzݳt��U8�OH�2KSG�{6�)��|�7��cN��oo,3�Vm��ϙu9D
��6�39<l?I���[�]�������2��}��l��h����}�ɤ�q̑��ƱФx��i��uJ�tgƚ9`�s7-G�ƛ%���Ր8�f����8�e�؟.�b��A�P(Jw�]Q�l�u+��5���m�t��ȝ��^�.���J'�[XxAB���eӱS@-	�%�Ŕc�a^�X�?fJ���k���o���%Ԭ��VI�:����[B̉�m�9\�oVd��-@�o��[а�4ָݣ�$�V�|�dttG{W������;Gh��y�,W
�Y���v�W
�{n���E���{$nC�@jU>s�j�л��J�Y�)|i��wb�}�OO���@0�T��n���zYΎ��/d��yBN�Dǳ���M�|��=d��y�����%em�k�"��28�p��i��e��5)���7�9��e�7?Q��v�ӊ����W���e�(�/�,�e��(�-�s�7/���v�6��>�h0�ZG���O�[\�"|u��5��"�6�&Ujk�]�Z풂͐�� n���((Y�V��՛�8^�����b�{$�5���e���� vb�u�W,�[���-^T��Ȁ�I���f'-��W��˦�d]��="}�Z�J�	����=�׌m���t^\eD���x�:б�Ӌ�	FB �Z�yK{[0y���se�9,D�oם�SyY �v�<�M����8�:�I}����L#*[���N�/@���!M��d�M�[��$��]�����ќ W�,U�ȣc�Y1Po��diu�}�:P
룛��	a���n��f��1^ *<)�Lȇ@���pٔ�p�Q;��g�o:�{�B�?���g�PF�{$��ګ���l�FJ����򲳟f���M�?`�;��Ob���%$�{�X<ض\y�Q�I)�j�Mf�e�Gi�hϘ�bcH�]K#�����7qNԝͫ�ї�׻��}->�aW=��wVi�UY�L;K΍]V���L�:�q`��.�|b�x�5�#PBڨ[��=�\:8s�L�:Z�f����\Φ�>,��R"k��7g���*�|~����4��>�s^����%u;g�S�CY��SA�Ӣ�%,K���r|f���﫷�%v��N#�8���U�V������:U�#�
~���1y�2�6L\tm�K�4�֡���J��岾�����k)�,�Ύ�}|qM[��[&�}������#��J\V�X������j��h͇3T7Ok9��R�yp�903�i[�.�%Nq`ox��3T�CE�V���&���V~��}ٯ�o-1GY��To3I\��i��N��zav���٣��Ӛ�Aӗ����Z�:
Ѡ����9�-u�z���%��^f#�׆�l[v����J�2Q��w븫o��a�ɂ�E��^��0���Kx�6���a[Gb�f"wJ�Nm7q>���\(a��\���bz8�-M[����On�E�"d�^��+�߷g��E�����W��=��Q!UpT|ι�q��|�� ngt�qԗrI�NK��Dy�D2ޞD�J!q�oL�9���~�C�i�(��#e'SOݹ���Z[g��cHh�����ě�;|ϑcA)��eH�%�c�wj�h%�s�m:�=um���ti�3uv�wd(�@n����J�nt��+���@�����Ro�}�k ��k�&O���&�6��T�g +2,_F��;��}J[*�1�,�d1�"�X�ˑ����5�}>�`E�a�E�'���f�h-7��onm_SंI��y�_�GsX�T�F�q���>d3���wz:�����UB#��"��/r�/^	��RE���A,ݖ�Rn�T�7:��'0�C��`FF(��x�9�-�K\v�_l����/��~B���+�8ehP�[�e[PwJ����O�J̱ˏ�4��rܥ�)��F��͢��݄�A�3Kеo.���Ik1�߾�]:�*�b}x���Hl��i�S)��a���魱�ρCV6�x��sk��?N��!A(悮r��l�fD�Fe.הn��ٓ-y��JX�w�I�/�.4����]w �Ԡ�>���9M��1����9w~�����J� m��c�.����P����m?�+r �vc�l5��� 8��rrI�T
̉��*�]�G%�|7�3?P��Y2��r��b�Ά�&���iR�R��������5`|L�fG,��B:�r��6)R<��y��i�h��q��h�S��IgP��S�:���)P)�2U��ɛ�Ҝ�����Lk�I�w9C�,.kZz� �%^�:rZ�j�����6�'Y��j&aʑ���j���)�y.�Rw!�,긫��x�6�wK�5ƅ��˳R��w�ב�b��!g+�j��ƫ�V���DU:���dj�����O%E�Y���'�i*�Ft�*��&H(9-�_��8�v��{��R�t  k��cxjVm�YMdr���p��b�5�����;Ĺ��()㺽���7(-�E5�⣙��ˉ��w�zwv3m=|�j������3Ś��o>�b�g슜jb��Z̔1�nֵ�����p��Ⱥ:�VHu����q��{�ᅻ.�F
�KLM֣�Z`WI��#e�a�&;�n﷬���=��Kt�26>��a���s Sn]e�BML|��P�Ѥ�ni����-�
�>/N�������gc��h�J=��}��gm^4A�}����w�Oƀ��32^sIX2oQ'Q��ݮ��M�
�u���?��H��q�L/n�]Y�����!L�f���^Z+�~�� �#6�#L��_���6c����������˟g}���,�AV�^��r���S�w�˱����9�ʹ<uT)mWo.�*��e�.�@��N��^�}Fx�8�i+ʠU�
�[>c�UCa�Z4�[�Q�������z��d���Ǎ���+;�d��a�g)n�Y^O}ܱ������	����m�E�XJ<(_Ƈ��p�9�#KK}�r�H�V��_YA�ypF@/���x�2����6��3,7�I<�>��8]72��\�ĝ>J�^c����%׵�Fle��*<���Zu��}�SvxAN��tza���g��䊿1��io^k[]B�m��s�ĝ�8�rDQ:��3�:["�n���ӷ�GBq^d�2�g��9w�#�*jF���y�8������e<��иȸ�iT��p� 73#�͎ݝ8�cFltf;��СcKd��g�a�o:�+X��<��$����'����=T�+p��:*�=}Y�\�
�j����K���O�u�a�����w�
�q�9�;�,�s�S�Ɯ�׏�hP��<&渚����CeC_C���E*#�t&l�Kf����8�"��>�tg���c:�����TB�=֌��6�7׳�Fc�iBR��Ӄ1:�7e{����U�Cj���k=�YR"o��`��͗#�74��L;h]�����]-���$�X�k<�lim�:}\b*��W����?������ w�*�(��~��/�Q� ����A��O���Q����!�`2�0,02���L2��ʳ!�!
!���	�YAĊ@@  ��x0��|�Up� �"-��U\;" a� !�U� �@ � �[� C" C C  C C C(�C* C(�C(@�"ȨȈʀȀ� �  �*�   C
����2�2��� ʪ�" C @ª�  C*�� � ��"��ʰ���0,2�0�2,�°ʰ2,2�0,2�0,0� C�*��ʰȰ�0,2�2,2�2�0,2��O����>��x ��H ���`޿��O���߬?q��o�}��0G������?(H~��?QC�������������@_���w�O�E��ʀ�@����� }�����%����b� *���������sD;����O��a��>�����~��k�AXU
  �P hUZ ( � � "P � ! !Ud! P �d A� $UVQ� $H  d�!]  P� ;�X?��<~��DEE�F� h@���c�G��/��?XP~����~�c���-���� *�����A��}���������� �s�$~������>�@W��H$�?�j}`PW�T �C����������
 ���a��z( ��	?/�L���	��`���߫�x~������ *��?{�����O���� ����������C������~�������$�����p ��C�G��J� ��������D>'�~i���?��~_��ϰ���}_�@W�}h>����?�<�}`��C��e��~��?����_�" ��%��ՃӄD_�����?�� �~����d�Mg��?\x�f�A@��̟\�o�y"QUD���DD(�UJRTTRRJQ(�$QI*I
IBPR*���* �JT��J�PJ^�*���P�C�D�¡�$D�jO�PD�T�*���
PU@AR"*%��N�$kER�TJT˾��A�
J��D*A�PJ�))
"E*��*�I R��JPBPIJ!(T$	/�dK͐���}�   Ğ��ڻran]t�.��Wj�*�7S.����j��n�.�ڧZ�wG��[ںճMң9wZ�45�rKt�\']�m�C��`�T�N��A�PJBU	J*%H���  i�B� H�
z�=44(P��N�
$(z.
(t5���X�ݻ�GV������]�+�7vj��Z���s���k]�]������˖ڕ3��i	**U�(�E$�   �����H:�\�m�m���rr+�wn��2�m�e����l�[m:�J�R�uwUmY+��)N����u��b��Ut�e�nWWWF��4�r�cJ���J��P�m�  ���[Ww8�]�5�֍u�Y�u��U�,��m�۶�Z�st�S:���ڪ���λd��uuʋ���#�;������R+k��]h��T�H�PQ%U$P<  ��<ն�����ڵOJ����Z�f�s��Rv��&�Nt��Z��cq��]`ֵ����Z����guZ�$��]j�B�$�Q_  ;ն�UR�t�F�Mul��T�i�%*;���� v�S�]���;��n�7h���㢝v���p�l���*P��l��J��]� ;��k�v�惋�tt�U��ٍU�N�kk,N,�%N�a�j�������Z �u,  ܎  R�HD Dm���D�  8� FyE��tΌ @�,@�i� J #S  ��@tu8l 0��NjUH�PE*�dA�  p  ��E�����@ и�� Z, �Uڦ  j�4)�KuN  t8r�  u)!TUTB�H�*��   wZ Nq�  Q�V  �0�˳t���t  WX:� ��. ���� �  x���R�  E=�	)*S���T�C�@m@ �JTH  5<�j�� �	4�i6UH� ��z��y�
9Opm��C[m�������,�3�n��m<�ӎf��ɿ�BH�{����$�$�$���d$�	'�HIO�BH�2HBI	�ￗ?������Ӵ�6�^�A�e�&~&b8��ˍ$��yR�BHf4:�v4����T��h���1R"�V[�5L{�`��qXɂ�4T��
�vM�#D���dnV��6�8U`��9w��	R��e��,�\�pu�����c�G���1f��a`���H��#SI�Ĕa��jb���Y���(\O��qY��2�ǩ�z�ޱ��;��ɯ�V��^�3U\�a�N���d]Ҁ�%�b���v�f1�Ea�N5����M��Q/��GB�����J<��R̫@��h-:��@1uZ����0`�{p^�<
��RP�JԠ����ĕ��@J��I�;D��w�����S��;�(���Ӧu�h,ɖ�w���nAAX�Z���B�=H
i�{����2<%B�T�f�B�3FU��E���`-���;bM�,�W��T�%K6�����4]�-�`�X�y��vU�o�kr��z
-��L⢠���M� �IX�^��Mf�C�ّ�%�W�P�t�A��w�5�Vl���j�Q'5��&D���ǑU�J��Z5) ��Z6Xq�'a��i�w���/n�6�VP�圧X�K���W�*hcVV��h���Ԫ��Yj�="��7u�Z�
JkJ������[v+5����ЅG����c7
�;���5�T����7t��P롵gM]$݊n�j�w)���I*hT�.�6�{P ʚ�7[��m�M�a,�b�iVő��
��j�wc(�PQ潑�w��9����ʸ��8�S�N��8���/���iǲ�ī�mj@�3�j���B����.�E�DF�ȨѵF�ڗ���Ҥo~D�8݋F*�*\T�����Y��d-Me�N�96� u�y4(��ت"�6�Z��Fnf}S�rdnս�.�jeR�NP�d��f�l8�d��B
HK̭Q��.�3S.�Xi��ӏ`̸��O[)�v���m�V��1�A���4+cH\��1ϥ���9xL(]$�f'��-hyL-O�.�B�NvLݖ��gM\�PT�*��fQ	X��:�N��F5I�mZ(r����Ⱥ�]D�p����XY�۩�àˊ���+G�2����n�5M��n��2��e`9J�&�E���EB��+ ӉP1��z�а3a5u�˥2�e�4.�boS��X�ubdI��6VUۙf�ⷭ�Z�0.L�F��"wW�5��Ȋm�Ǫ�ꎠՋ�R����t�(iƦ=n��!@�bAua^1�qT�(c��i�La�^^}��&�Z�@kEۦbE�ֻ���W��-�*3L\ڵ�aķ,0�d�W(���`)	7x��Z4��	V]3:o2�&dߦ���,��Q���A��M�R��,��d)��LY�HL�OS2���)�9�dE �S�E��p�E`$�fa�E\6�*�`D�!6�CWl�BH]ӭ�M�Q�ww��])W�z�<��I2�-���U���`Z�K��i��-�;hIn�#a�*a�3D�D�L��bs캀�͂�Y"�U�Yo����/63&�"�F��&��r�Ci�Y��{a�G~�ݗv�\o!Z+hRѐ��W,���҅a���f=�d����J83(�S�F�^�@9U(<GVk2޸*�*�iYxIb�Rw�o�J;ueȅ����ً:�Yf�r�&c�4E���E
Y����d�֜hj1��Q�1q	���MRZ�I�Q�u�Xf�d�Vgol*�je�2�٥yS"�3!?=�u��%&wA�C�ˢ�L{z�KA�ٶ鷚��	.�?fз�R���]�6���y �1����Jm���LC)����D+��8��LLZ)�-��Ȕ��P���Dѣ�nE�I5fA	�r2�O�c)�)���ӎ��Qw��KSP���V�m�CQ�r�5s�^D�<Gj�l��x��7IҖ�.�MۨЇ���-����M	�ʑXq�.�Ӵ�3D���ܬ�JL��� �.��a�0��CDu�!g��l�ױ�������*hiKlͅ]�n��.:ט�7�1զ���B�m�x���h�EWt�ŀM�t�U����Y��+m^u�8���Ã^^���;L�(�3���S�El���X��7#D܎e�Î�j���Z�J�R�}��e�V���F�]�p55M"�4�Ê^�&�� m��q��Z���[׃iKt4�3 (i4@4(�xPz7p�Jl���w��*��8] ���æ��5��0���B��W���Q��zi���w�+w`8ra�Q��֛H�2�(�VF"C�ue$���z�
���#n�j5f����Y����t|��D�/��YIaBT-X9���������bݼw>�Q	n漡A�̣
�܅M��ܬ��Y,� �\Ә��J62ƁsM]��9��Z�P�&�4i`��*�j�nӶ�[AUʭ'rɦ��(3DP�	��f�VֵT�m{��1������ff��u�Ӥ,-;HjVHf���
q%�k�X�*�A�+�V�9%��W�䄪��-�{
L�́M;D�u1�Z����kG��[�PNl���D/Zs^�eM�[�Y�(�v�+���H4T�v�%Ǣ|�mhY��j�6.�;�
�Ǵ�D�@�rb?=h��XSvYX�5"A{DQ+��H�/sfŦ����;�/5&�\t1e�{q?��b�Y;�5�����WG.2��J�N�*�����)�U7�^�5���)�-|���Rcч~�V�h�9�0��T�A^�n�� ��^����V�E�� Wr��^<nB�
��J��ұh��T7��R+h]<
fZHjؐ�cj�6D��E]b����{yh��I��T�JS�i�gP���U�/�iӨ��G-7��-]��.j	�k(�����f����(�:��) 5y�:�9d<f�ɎWf�VE6	Z���F�X�6�4��A��!�d2��$�n�����l=� �Ыhؕ�M�1C(�hV�$�#d�v�gٻ��Z�on-MRL]�eB,
�/�Y����Ӡ��o^����7f"�of����r��<#E��ғr�u��WN�<B�.��Pmn��9����:�+�($am] �R�b� G�	�e�à�_Ś��vI�cZJ�	�b�4)u����x�҇�\�>:���������ݠ�%��͑������6-��,����A��ج�p$R�a���mlǤjMbL�'�.�Rk6<@�ͻ-���%�٬���3�/TD⩒d����.UC��VU�g�*�L*h�LpP��XU�[�A,�p毭��Gq�w�zٺ˻�3jXN�G��C%���{i�N���јi�D0�mj��5�Q���N���a������)��c$�I�ƥ���uJ��YF�R<�p[
�{������Wd)��k�F�T��H�N��G`ҭ���ZJ)1Y2���(^ˬX$�Z{YYYr�̧�j���OiZ���n�dN-D�ޠH6��U<o���XȺ�6�MA�O2�j�(��Den8�nѴ�1�XQ�b�d6�V��H�H\JlV�`2���w[.eV֪�7��zB,:�������ÅJ���m�����fN�hRK��WG1�Wt���a)�n^,3��e����q��$��{�(b^�e:��I�N�2��.f�H&v��e���6�`[0C���y���c4�wM��^[@�wW.���$��O(][��m��N�=9�n��p�� ���k[q�ɁZ���R뛫ǘ)e��\��KYD��2����8���L�4�ޗAKfPMe4�L�*��!�rĥٚ�K�9R\���nSu�����[kUe��p�lã
z�ź�=2�XgN�&��0�-)�P���n@�j!��y`����r�T ]��9N�m��Y���ghޫ��Vv@�Q�pQ�9"�m��ܩ��[�!�%��me*�;L���y��)�ƒR��9�>�.�7����2</�*
[l�X�1�I,Q�6�n֪PdpIZ+@7��HC5�ˈ���n׫$�[��k0[2�qZ�U�˕h�ҭokY�͆ލ[I-:~T2�w�k�B���p�������ͫ���Km!�S!]AB�(LI��&�V0�f���h����L��b��Z�bSD���6'n[)[�/[Ur��I�ؙ�X�p��Lr�$������W�R�l�t��Шf'S�+7WʲP�#)`2=-��.	+ov�Ld� Ư�xQ*چ��r�<�SkL.J)���/s\چ�7u`���I�t��Lf�Wa���/��![���U��Ṣ�h�ÛO�X��/1RY�uR�*�Y�1�y�-�Q��F�W�=2�
B�E�!�2�Mz0���%e���-+L�[:c3&f�I0�H5����ȕ��1ҩ�Il�����i�%+�>�R/��f���.��M����;�lp��e�׳ w�#y-�KLލI�L1Y�-��
�F�u{���.� ;�3��u.�G�T�,�4G6�i��cs)�Z��`� �2f���Kr-
Φq�Dl�u��36l�QGY�#U��3fH��pj���޳����ee� �mXm�qH��PZA%lA�Q�����6Y͚�)kPԓ��4�W�V�Z*e���t�b˭3D���i����ũ2ͪ���`���3i�� �R݇A��ݱDѠ�n�n9�i:t�W1�ǔzt��;%�D�y�m�����ma˃Ka��^(�԰&e�����_�jam�z֒�ҍ����B��`�(=�v���۶�>�WU��q�7��9{R�,�Z����bV��O7�b�VZ�f���n�xn�S&n��q�l�k{�!EjĶ�r&m��874�ͼ�2��0,�-�>Q'dP�wE]��6X4��e�#f�F��Rl��;&^�Xj]ԭ�,�uٺL�U�^��a���Q���`��Sf'u%�{rbv�&��/�A��)%R�ѣr��GV<�U�A;A�crޖ�efT��n�:2�1k5����H�n���P��l �,QF��ԑ�����������U��X-M�����0d"V[�O	�n�e�F�R캒�5�[s0��i�D^��9���7 ��MϤ�$Z��WWJ�i|�/��H%ȶ��5����1+{H tԬׂ�4TU�u&�1(N��[u�K��R�ٗ%��q:�qm�;b�%��B֩h���V2�6�U�`��I�w	P��j��[b��<�B�����P{�v�b����*��d�I�Sd�.=���Z+v]�X٧&�4b�J�X���m捋�1e�l�4��I�*i�ji��<`�2��+rA��Q�I�l�=�U��4� e5�&���y�˳�6�h����2����j5wGwr$�P�m�p4U_�+���e�rQ�y�1�R��t{�b��	�N�z��Sv*mk����1&�#�Zu�Gi��ۣ�wfнv�$D��J�L���'Y�j�
VlC��JrZ'wq��M����/6����BPM˻��\��C�L�L����t)eeY�%�VQ�6	�$v�T\��i�n'�YH�J�y�.��Ze*��7�+~���&�t�F��'w�D[�O	i�c1�fn-zX�Oo↥譊њ/!bnn�y4ЏQ0d�-��h�.�P�M&�d��Z.�
�W���JQę�-<�Al��2&�L�V�͡�Mw �#
M��t6];'[��@.V$t���)�tFD���L(�˥�H�[�����
�y%���*ȡ%�dJaٰ��q�ҫD�c��H�A�Bղš������fD�+!��1m	�n�"��Ub=�ba���n���쵖�$`���	 V5u���_^�)lT�I��c��`e�Y�Ѓ�8fIV�ɸ^8�D��&hm�W�F���&[�՘�ǧ���	�/
�!� �4e����U�gZC+uG��d ˅[r�Am�b"0]Ũ�[�"�P蔁�tc���ӆ^4Py��4B�HςZf���]Y�֨�IE���naD-7��]�;ki��,'����a�����xQ��*-ں�g��.���j��'qԋ%j�WwkVe� M��]�[V�4���f�@��+D1�/`�aZtk�M_̊!P[���i5'K��IF��ut5a�����.&��"��SF5���co@@c��/�#1l�sA����or҄Gc��p F��6ʰK7M��.�m�k�\�l�7����W�I�d�IV�bP�᳖F��]�b:�7L�h�t���Cf'x�j��i�{�5��j+d���b�SX�/o�R��EnU�Ga��J�N�D+R�ͅ�m�ҡ3
������,��բ�j�"����#�Y�tl�w�P��s2X1:�i�v#u��V���Lb�+0�w���A*X�EnS���6�4e��3/�)%�LH.♱ԗYB��݊ړY�\5�����(��*Ɗ6II��u/ -�V�cj)��f�Wp��B�٠p�$��ǀ[�9�骛Kr�,�d� �� �3@ݳm�Ԭm�)�Fa1e�&2f��WdM���V�]�F&r���ʎ��Zݕ�m�����0���DHTZM=Q���6�DM�j��$m�n�'�\^��o�`yj�*7/ajm�N8�:3#��B�'v�ժx�P��[����w�X��� ��,�s��Bع�hl�c�w���gCP#l|��dt�*̶��#7]x5e�g}�I���������-3+\�<W�B��@;�}bm3�8��p�Sf���c�[��KD����+5�q���bɛ�VXu���_5��F6Fu�0eY�W�K�/�*�$��g���}�u�g:��;|��*&���
/f=�8��RUi����OEn�-#]a������s;5���aGK(��/��aN��^�-*!�i[�H̷�\�7u�UN|�r������ʚ���\�_'�W�U�%�O^U�X�z�E�[v�_E�*�+t���ݵ*.��s*�[�����d�cy�����7��v��뤬K@�7�Mf�65v�W���P,F����-^vQ���^�+�� �	��B�(�|gso��{��X3�\7o�
�ų͜xbt��ۃ����z��]FWB��*�Z�T(N2�h%3��J�#�1�X8�n���٫G]J��tb
�	��8��sfR��Q3A��GA�ەaɿ=ݧ켣������ŉ�3w]�\j���L�촑��	�
�R��"�_ ���WMH�gr��=F�%EN��Q�`��kN�R��Kr��:�L�;�}!�wj���ݢuu^�+4;o2�]�n�n_r �����0V�Ѯ�rX̧W}B�����3X�f��{��Zyn�N@�Dq쩃.��rӍs�*ӛx�[�2��oN��#o�ٔ�,a���jԴ.�ڮ;'�S��hj��!x�@�_VCr�v�z�f@�@Zu�W1�o��2��P�Ko.�[�wbW��Y���\�D�.��M5n���S(��&�7L+��:�H��{1��cۧ�gNW%�2�Ҳֽ��	��թ��2��=60TܫӖl�1K;�i--Пn^�V�t	�MA7y�	''���T�,�{'hCFI2�1�&V>�v��-���K-ĝ,�|�4�R��Q�Apw.�^4_rX�F�����2f�g�{��˰�����a��m�c�fd9�M�1�k1N��ىP�K�F���Ղ�imv�v�h�Hh>��oK,�*C�_gr�7�4��Z��/E	V�ә���-��bt�L��Zս�P.�a���Y���عW[�6 /��'/�/�N�
n���=�\\���I�|��7Y���g�q\MhZ�̚z#]C���-}l�޽�{U����u,#���5�pw�oH���[�
5�Y��$H��N��刲��;!"��3�!�NA�p�$���8�>���w{��#家5�&��{k���#�����/��Y� 9���X��l=��s�@mr��d��bƌ��(�T���ߎv}ۦ�v���OF�R-(U�H��<5ko�:�:h_}Y�WŇ֍�C��b�4<8R��7�}��{Q�mƔ.�3`��I:��M��*�%F��"�̶���'�kY�r5{&�4�:��a��kG-�-=�X���e=#p=ˌ�t�A�S��-����oE!:��n�F署N�&�.��ڢ99��e𥹽M�˱u;�ثH=�C�k%��Tf�-Us�@9�+>�Q�&P��@��.���wX��>H庮P[�%-�eoFD�����K�֌͢s����6l�h6�� �����|�ڵ&CO3~��T��Jln�:�e]'=1��[E���LЬ�$�4@n�pͣ�[a5@�U�������祧��%��b�MP�0�z�y��|���u_p�G*�p��pmt�H*�y��H��8�H���L�P�Fa�.�O-ϱ|o�T��WZ� n�U����΋�'Ptlu�^R�rй��뮬�wL�6	���+�o�K��,"mP�RJ�SEء�TR ��f=Ł�]���.פ�Z*��&�ZR.���g�>viM�Zd)ְ�V0�P���

/��Gr�|�lXY/P��eӪ�U�]5W �B��ĝ3�:Vk�<�93�G�	q�u
ٽb�kz:Q�.u�ۃ:;E#�*�.�����p���[ܐ;��|93a�8Y�Y�XY��Rޫ�l����`���jkR��^'v�YY:J'��Ň�tj�ia�|(�G�3�̑T�F�'�ǫ+��>�F`k�Q���w*�����P��x'Y��la<7!���i� jv25���f=zb�G_t�8�p�	d4xk�Z9���Dݣ�\��[���P��{q�'[��-놺��!�i��@zYdQ�n�m	��r��X���+$sY/*�WV�tᲧv�Ґ�t�L�Z*n�K:k'"�������ۜ;o^]љ���zD�BkY5T�̃1���WmobԝåZV+����%dI���3�:^r��)�%2�S}@;���k��r������U�J��h�S��-n����L�"'��Q�y3�;�j�R�;���B��S,M@�,�V'v�ɡ�j^�4�^�{��
B�Ï-�u���I[4�4͛��̓�z��nLd�e�BLE��]�;��YC�	wڍ8���F�,��q]_ru3IŇ�NU�_Nޫ���F�.^LGZR�B/��gY�u��E�sh� ��+͌l�Ҽ|=��!C��
iv�[,���fLuH�
�S�V���q��Ń)* E���y�vz�X9��&_�/;�m-�ӭ��L����P�y}�l<S��AM�-���WB�ڧ9ސ_҉�x�k��N�C��5�	y��tf�o:7�:��It7:�u]"7�U�Э�h��1:�os��O���;q����h(�|�8L�����s�=wn��6e6*�Y��p<�ؔz�(����q�Y����	���%С7�K�dpV��@�L�`Zӛ��6�¹�2һ�����m��\�)2E��Wj�@�$�QX]���T��%,(7nl�NVӖL�3v�2��uђ���Ȋ�L��:3�����FE��e+�u:T�ϛu7���C(�˧m�`tq�o�l���8���b����!�˺O mf����[/�]�͑�Rخ˵�s3aܱꏝ�a���������8:g"��#<bd.b��Or@o.�9WSr%њV��}c]����iڪ��}3LâLo��Y�	���
g�`�$RP.i��F[���w�gGى��r�}�i]�](��-G��w�h��c��n�+���C�*��v�/��Q�Ԏ=wH*���Xb�@���QԆ��L�X7��f��Z�V�igv6�^2�ܙ}Np̨�֢w���
��9v]i��۽х\���p�K,V�rK]'-;��
��͂c��m�"+v��(�oe��
2%�rR��,e�;��[�V��m�W2�]C8>su�OO����Q}��o�K<=uq�}�g,s1X�e�]f^蹸��u���;Wv*�*[L�Hݗ�ģ]�k3��s��Y�S�ָ�� yݾAs�78�!�x���+ H�}{�zo�eЦK*ղ�F�&wAB�6o�^[��	��U�0��[�r�7i��u�Wxd���w�v$�!p�9Aǰ�W<�ÝKT��[9���Ī�oHP�k��%b͠L�9�y�_p�RyFge����2�_;ʇ��h�Z0o�_n�Lm!J>f�ֳ����c)]��;X��9-6&����������ծ�h�5�-�6������ʵ�M8r��jZ��Soo������]۳����^�l��qe��)�b$[�!77tT̶&���Ѣ��&d�����}��
��꼾C8��yT�mo^I�I�Th���s3�w����7��o��_9�]�S��fR2[Ec�s���J��P�s�G��KU�:\�*��b<�
�L-�7oc6��g��n�^h*�>���̹��'ĭ|��sb�ޝb����}9�{ñ=&����ڻ���k�o1�;i�NT�Y�AW�q�XL��H1n�v�Y"\�K�ac����m@1��@5�Cz�p,$%L��Wv�+hꁶ��<{T,�wr�9�A�,Q��@i9<H$�� B�m뛃/*�m�� �}Ժ�zU�T�&�k�*guZ�6�.Yݽ�v��s����]
���v�%u�<�9>�X��Z��ʟa[�ᶴ�S1
��&�EQwnA�Lp�;�摸� ��H}٠j�E.j\-�Imq����S��c,'�W<Kvϯ���/��1�ȴ��F��Aق�}��܀�s�����g���k�4��K,�5\✢��r�Hr�7����)�J*�:#]&:	�#���6-S�o&{o��Qd��%^�m��u'�X)j*,�y�J�ҮEr̍�!���JɣY�fq�X��E�Ef����
�P�B�����ObiۧrM��pt+��z��P�����i�	�Fޒ�*��:T鋪�N�/3O3R84��7,cn��.����'ܐ邺0�gP�RE��i� }� �y�o��t��}r�18��C-e����/{�6��
`C�X:K»�Ί����!"����0��ܷK���Վ�M�7Ϩ��7f������<�×Q�3Ց�&�Ӎrk���Y�����|�|����v�T�P�1�L��2�RHƊ\�E{y\����9�&�r�M���Ck�j���:������ά;(R, �i�#MnE��sag*�]��(_R�5p��|T\S%v���q�� ��N��Q��[��4�]@](;����h�6��)wQ���z��W0����\"L�0�q�7����{J�Y991S�NeL���2��I(X̛7�>Y/)�u������ޠ�o<v��_	�At��%U0����K3Qbf �^QA�Z�̕�V`�����At��Rn8�ai�u��ˋ����,�)�ٛAf�Dw̻�Q�3�c����1Њ��X����`����%#�\Ԏv%(����M�C��\��ZTU��,Z��!��z$j*rp���:���|��Q�l��df��[s'fur'y!��]Oo����#��Ҽ�-&h����M��7*�p�lw1o_�T"C��U����E�5ӆ�G5��YsUTՂ*R	k�_.��4뭝���t*sU�:���_[��\���bw�����3�#�5mXq�.��1Ê��V_s GYUoѵ��)r�\B�¸����Үu�;��R�^*𤧕f���*���٪ovAM��Y&:snq�������:Ni���l+k"6M����M�����5�3�2�:�U*�,=���_=����#|Qws����K�ׇr��i�?=��Ff��F��I��͂t��iEu�oh�r�X��ÐS��б9��*v$���}�N�������w�`s�m'q[хyø�`d��<e��-�+��
��ưH��壮���i	v��\ʘyR���=��V�(Hʩ���i�'=�
�8�+�����e%�ڀ��p4�"�����C�y9t��[��xBX�[A�)5�vf�V��J�ِTsU�}��hU@H�h�ʰ�%��^]��!z��WmȺ�y]�o3 $7J]��\'IdKKN �p��2���,���.��˛fg����	:S��ص���iٛ�n�L�D%3�k*����7d��>��uL��m�/Fd�4k�F�Y߇d����%�ZS��M�;M��V��7�I�T�1J=��fc�q ��j\��~�*�þ}6W-WV�s.�Ji]��q=�7���I�\nl��o^�Y;��K��T쒵�+@v�I�~v\���u�̰ւ6 2�:F�N=�c��Sn6�(hvq��~C�8���<��xlVjQoUK� VJy�\��n
�gKԖɰ`:.�aL�B��ABt�

ɔ����0����ӧ��J5�F��kioK��������G�}a_.���<��ſ^�|�U�H/xæګ��F$TܕYϲ#R�j��ƚ'-H-��m�]�h��RwK���֊�/�`�e�.�c�X�̧��:�V�m��en�j+����ҝu�V�i�yyt�2��fκ���J�Ŕ�
�=�sB�M ���z�no\N���%Z�]<N�tT5.�k1���g�Ā��jgN�t4��% 8�,��W�8��1%d�Of������X�g��+�׊���V;���n�X�`$�����c�n�#o����+�%f=Ԥ]F�U�v#��}a)x/�t�^kٕ��$��]���a/L|^�En��+يЭ�����K���W���>/:�ft�[��ŝ\�iurn��L�=m���T��ӡ�,�U�J�q�[o��kt/�<K%��b�����N��Ŏ����J�L�ZZ7��)h�}����TN,���A��Q��76��'�bbxF���EZ.mt�m�ɇ����Y:S�r�흈iЙ���7b�֨��ެJ�/J1��t˚²[���4r9�C�2c�-`Hݝ�0��u�}�jd��X�{oZ��_���"�Rp8"���d\��
�����ƽO�7�P��ȍ�
��ɾS]ue޼ů��}�_v��K�Be ��p���Æ�dY���N��>�g��Z��6�h[x�8�-xޣ�3�\o�,g�G��r������ТaB�E��n�Y�����6�Rڮ��[�˵�e�Y9.���}�(Xk���+�okA��7�y�h�E'_^5]��	����\oT��h��c��P�Vf������.����q`һ�p��#7�شF�v�����<���+e�y�]EܲvѾ��Z���]ѭ��Y<:�}7{�&;և�Q���𷝪����;���N)UέC��F;6�:ڝ�*�����!���Y�Ѝ���})��M�dBN��m��T�{����٢=5{,���Y;H��ৃ������Rƺpٝ�gcS:��oR��i	���5#{!yեY�	Dڥk1.]�k���� ����]
E�w#��9n��nw+�����=�ٺ�"�por���=��  �@�$����IO����ù�h꧉����}�ʠ9��:�O+:R�:u�[F�)v��1�I�yE��U�hbc�0���q�5��,f�����E�۲�=4�\|�x�_�Br�ĳ��0�J'�ՎB/]p�1��ej�׏��W�5��}ó� ]�z�n�oSt-j}�Y�R��d��#�%��i����
Z�� mq������"�_\����oƮ
&�5�{ƅ*:�<y�(Zz���M��<Bv�b��kr���W�w)�{����)|�Ui,�Vtې}ks���wOM�Y\�ט�꡺�����Ry7�%�d�qMՔH���!���jv
����j�3\�v�U��>:�!�s�F#x��o���V��LnQ[%4����W�ݩR��GGS�uwX�T���X)�mQU ۹
"�� �.̾��Õ���[;����w�����.ə�ݐz��g�:���{ݴYG��s`;kc��b�r�k��@��O��۱���U[t0�6uX�A����R�v9QY��H�^u�����/��A��0e6��Z-�o3��S�sz�$d��6�rAYM��h�[��ٚ��yۤ�[�����JN1�Z�����6������ ԣ�:l�J��3����S`ot[
j�n��wR^{�r�<�q�{FJS\�EX���i��0�*v�!�p#z��5v3\ZJ��� �w�Rs����N����N;Xb���F�� V����1���ҳ���8qr<�go15da���ԕ���f��Į�8)I1�`�{C��`]�VPc(�ی���eB��l�n�V�"�j��ډ��v/0���n���9��x�Du]gtܨ��n����2S��d�}'l��93��I������Ѣsc�n��0�@)Q|�_*x"pţ��'�sp#��y�~��,����.`�q�s5d��� ���1���j��]J
���Y��B�ZR��O\�5XW�޻*�J�٬��M�6��u������ͷ(Ű`��T�t{d��[s�Ķ朊e�*��Z/��l�!���G��/A<��я�ɖ^�jK������sT��:��\�s!�9`YlA	�q��A�.Y���U����}��V:�W��M؂Z�z8Z�|ɭN.bոjR�;��G9�εg�ԭ�.�LLr���V���Wu5Z�uT__At;膪�.^䩥��7�}P,�y8��7>`X|�l�R�/��E� � ۣm��ea`�g�׹hc׶2b�Rn����'Y����vܵ�X��¦o�ۮ�3#1u49�,�o����Õ/������j���J&��H�:�;����CC��
�(Fn�˱�GV(�IJ1�NGv��7#���yC8�}ϟ����a2;��u�\�Z}wUC�l5����n��(�r�޻��h�WS"a}}VVV�f�rޥHF��W���Fv]\�%"q��X�o�Od�rzWgFR�m�9A�Y�����:���j�7Mo��\��>|�	�9��d��6�qf�\�xݍ{�=<��we��2F4g7���.-�-��Y��Q3.��[�}��{�G-,)X�[���(K֥{����C��V1S*�th�k�5l�HY�o�m����3[�ʘ��WA����t%Ch�[u��w[�̙m���7�'������#2հ����ٜXR�L!�+X/T�]��F���C(`��� 8Le�n�|�t#��0�ḫ�s�Go��FC������,���MY^̥Y5U�.����3��>���k��u�5�N��rU��3숒��x�n�ծ�2=�*��c��#��wWזB��.�1X���0�]Ț��3/���]�Ig> S�w��v'�D%s�!s&�-ը�����g6J��.�݀������_ZVwt�wo�m�o�˶����h�،�L9�oY�svf� }ˊn$S�ᝒ����J�7�����fˮ��J+z����F.5����]r�NY�j ���:�f`��s9xC��J�+��3��K.���ؒ�Ow9��xrݮ]����Y��32�%`��@x�4����F�c��b�&�wv �$���u��^�J
� ���;�*]�����$C�N��J�B���w6�51	��M�����nV�-�k3{qJᶪS�&�)v�v��rc��)�Y*��3-*Y)���a�X��V��4r"�YE�T�ӱג�475�{qo�u���V)�Cǜ�S�N;n�K�q VU��X�Wu"�Sy��}4A�ʺ��<�DT{]��<wڨ����X|�����WYܸ��hW�+��D��U������Pه�^�s�Eg��p\�|k;ղc�Э^oI]/�F@"��[=���b��9!�f�����k���3.nHP��l����Pb�9pJҀ]�puz��W;Ϋh�,��p�v+C�R�:��p�㺯;luo6n��L��8��S:m��wu��V���
�n
/��wT.�i�		�܏6K�ö�\�}د��t��Y�u`�n��T�+���/CpM�΂\\�
�����;źpv&��\,���b�!+�ұ� ���ۇ1���^�)�Ym��rR�\61�M!��p��-Y�s�Pʠ[i�\΂�n�W]/�ѽ3�%A@��{s��Y�6%Ŷ�X�tX/�	d�� w\��<b�������U[��$-�M�8����0��{�
[]z�єT�a5xG<� ���N�AWb>4l���e���(M��:��I���%��hp�6�[)��42um�pХ�-�X�l�&��}�#��w&rv�W��Ν0���ʳ�ebQdhm�	�T�ݟ[��������=���v.V��p	l��u)��n�r�XĶ'C:��dCj��.�!\��*��p'�"�ϲ�fN�pωRt���c��m��`,��m`-�)NWD�|�k�2�9��S�j�w?���YE�Jv�D7S7k��\�7p�
�Dwvo�R�MǜΓP�t��Vi�s��[�q�_p�}��)Tf�n6�*Z^��Z�lE;y�~��A��MH��h�	1u6{���T�]�-Vsy����sp�0��UZ�Z[���������gSXU���U���-�Wnԥ�p��Dq�܋���/��P5��2��Ռ�Qog�� �/N��I���O�wq7���-��r-���}.eąX�QoE9>,³^���Gf����tS�u��PFQ�G(�\�f:�J��du��}�ݻ�Y/B�ͪw�vJlJօk�c�6������N�_Ý�x5�SZJȬ&����D͌�_guXǡ�Qr<�a��s��V��U�MP���z�UԵ�Ӧ�!ٕ�Ԧ��g ���fe,����!�3s�����ދ2���K��J�7�Q��
��×>ֱLSs#�sb���U�ҁ6G:0Q��.�jݓ%x#Pl8)^�Vkb�e&ܛ8��j����W���d�}�W �n)�Ҳ�Ŵ���݋L4�wϳ���bdQ
=.���i�:�ɕ�ͥ�(R��Ѧa��K�H'
�5'U�9tӥٓ�Ƶo�6���V-vs���yB6�b`ouC�=Ϻ�����Y@�x93.ܥ�o*� j{�����o,�9	Y|���A���D"�(�T�V^9H��g:pm�듯Le�X%Ҙ�Ad
�}`՗���f�ԝ+�t+fm�K���;��������JZ�3�Q�� ;x�:��.z�@/�<2���.� �<���S�����PB��[������+l�nh� �����H*��,��Ր��q�/��W��y�x|��Y�� �CsYzw�N��RCW�Oc��@Y�/S:�N�����
/�i\Ļ*^-Cjk�b0\j�h|���6����bI�fSZ��֌ٸ#Z�G4坻��ݭ�4��!(�X(Ӱ�!mTa�u*:�֠T��5�\1̝f��_9oN�Y.U�$�)^lu��I�A�+/Z�ۋ��o3�:���Ԥu�{P<��fDe���r�MZ$�z�/��(����*C���[γ�r��`�L�j�ȐI��T���V�*-C8�`+ͮ��Xdr�\�����(V)v�V��!zQ����i��-#�r���:A��2� �9�oN�ZE%G^gurL^_&۫����N9*�&*K��R�͸R���9m\��j<��;�Pq�a6��ykB;YH@n�?�,ʘ~�B��b���YW+)f�N�]��gMμv;��
D���dq�L�B|2[�X�-q�[Zt`=�U�b�Z��uv��t������g*kA:�AX�>��׃��v�k��[�Y�ًk�G����ֆ�
΍l�9b�|$��j��jYת����w��lF���l����FL�Zv�uv�+v���vL���m�M+�V�[�g�_K�5�۾�_X��:���WW^�m�ᖖ�^��a�ǝ�&��*ZZMK�$c����y�-W\�y]t�q�i\K��(�Y퍔zop]�I�v%Aw�ۭ�-\�fM/��;���-1|����F�ݾ�}�t5��9el&����(����̚;���������wy�39Օ�����<�B�Y��b�Gq{,�����cz�67�R[��OV��W��q�����1Q���n��}�,53k�C;��#��.��i�j�'>�M��U�	JT���W2���w��ĎboL��'耝аY̚zeQB���OL��ހ��D7�b��M%/Q���,В��ݮa]l�|�~LU���׈�QޭY�&,+pSp�5T��[�B�y���sh�; ��X*�K��raȉ�^p3���}E�����Z˺�[ 73P��^�[�%b�*JSMkqGEӎ���O8�V�d�z�\��ƕޚz�٨Vu"�j:�]]�m�����u���p��v���a�*5�ڸ���4w!	1me��.�V[�h����l��:�*+��ˑ�CyXV���ή&ξ(������7�����-"Ϟ�>��S��cF!��Z-�G���̵�	ܳ�Τ���l����Q"Ȼa+[��̍�ݰ1s%N���.��Nj�(�N��T����3yZ��K��۝�#��E8C{��36؎,54͎�6��<�:��xk��euJU��rr�T]Ʒ{h��!���|�t�v9�$��S��%�v�jKB].���Z��*�H`uu��V8Y��,��/CS�[ٻ'G\�W���n	0m��m�/D�7�^Ŵ���ΝL��t*ڀIHW�'|2ɮD{g+o]���]Y����6Zm1#�wTH���z��a�x��
t��C�f��ws'" ����:�u4��hb �QQ�l9b`�2k鶱5���<�XqQi�n�,�L��Wtۮ�A��Kc����%��ѡs&^����
���7��W|�e�W�e��о��ӿ��;f�M�r`��Ǖ��ͳ�.M8�����'[_F��-6�+3a�j´�ה����V<YzI��-��f%��U�����͝/q�Zo-�֟.��8n���ۮ��z�ց`�͏����;�Y`�AWQq������u�7�73Qi
�֩���6�,��v�Ef=��7[Cm��k�-�&q��:��	�B�T�]N��K�GI��D�j�_��+�:Ki�M��ڽĬ��M��EӬy��"R����%K��w���'�P�'a3��^o
�yP֏���Q�벉�X[�v���Ls�̓�K�K����+r���g��3s�N��{C*ڒ�s��t�y��H��|��ȕ��vC��%���Of�t�$}��Q����_n%��׶мq�L�1r��kq<�y��Ki���s5�Qr�e�]���8}w���s��J�+0AHK�\���#c�������WI�,��b,�q��,�ԆX���Wl@k�q�l2)́`约)z*�m��tʾ}�Y�z����d���r����ri�|w��u�O���v����_� �s]�b����Wl�A]'^#�^�2�*]���[��'cz̊�*jR�����4GJ���l+��# ;֩wTu�P�Og+�]��޾�ol�W '*��D�[.�Z�(����M)��>犦����C������ŵ3t�1̤�����#���I�E;6���ƥ����rt:�zU��RtҵQ��7�,T�9FXҊF�",իv�8+R������ٱg���
��5�\h��ov�L<r�L'�a9�Er�x�49(f���q4h�ݍHv�WT{F!4���u�t{i�6�\ЬTZyY�[���4�׽����v��N��w.��Ί�[�1`�G�f�r�k�3��&����=YY�MǕ��2�Dn���3)��ӛG�ʇ��=Wb�RUێʛ�h7 �F���I�pk���X:uI\�r��f�[�L�!�)�GȐ������yS�M�y�g�e����3;��_}�k�h�Í.���׽Q�
s�clZI��ZK��F��[$�i���;JX��kokT�yPC8uI��'Gz��ǫn�����f!	K�k�yw��5��c䮛BYi�޴(�̼��̡L+���.U�m�2*�*T�5s'r���RJ�����X����w���y:k����I���;{��'H�l�U3�.e)(�8����K��8��ͻyҥz��ŗ�����{F!M ��q��O��c�]���\D�����������[�┈�u飕��ͶS7��XP%ԋRZOn��V�U����P�W�ȇA�b �i�����4M���:�KȆ�Y]����Q}3�i9[�����w��"n�;"�Y��}��x{� Ú���)W���v�I�3a�!F�T��p��0<�f]It<6[k�kD�#5�V�=۷����'hgJ��WgG�\�:�<ʎ��v[�B;�Wwӵ3���L2�<(;K��vJ�+)��o�UNw ru�Ȧ�eVH.��sOp�Xv�׵���m��wTɯ�����]d�@#��d���J0zpz��%;��|���ە��@읗�rN,z�*ٝ0�#y�Ar|�"�YYK��Î.����a�u'.=*���0S��ڋ���x4�ڬ�f�ūb.HGngM�TJ�N1j���/E�7F{ʔ��Q}�p�h9/]��d���Υ�����a}$��� ��l]�؊+��w5��F�kZ8�!�������.�Ksya��gM�[]B?�ӡ��mj<xqꕆ�X��*Cb��ݔ�9�mE �b� /Q}h��.}sB�*U��ÃOgZ�Z�+�=�w\�O��^[��\��y���
0��q+v�^͵
�g}r�j��)7�7��2�=����m����3I���q���9�P�g+e���*J�����}4��:�$����ǖ�emM�×f�� 5��e|����ِ�oؼ�>gs�>v�ح=���tdRS2�$4��V^��Z��Y8{�X�g�Oi����/O��a	s��Jܽ�㝃�fP(�6��g8�\xQ-+����Y&-.RV�]՗9<��`@ ��>�ı,PAe�Y5�J�kEFڋm**�h�-�����(�UB�����J�Q�)R��A`��(����,��d�S�����X�AE�E��ZXTF
,bZT�Ԙ����( ZETA,1��ň �-����$EE��$Pr�X1G(J�2�LJ�T-U�����kQ@EEU�S�c-Db2T���kE�*���*J�UB�UUPbCQU�Y\J+*�T�Ubȫ*!��e32V&R��PT[T�Y-�ZE����1������edTamQT���dD%j5�ն�����F�b[VЩ�PPX�i,��X��̄+R��b *�\-�Ũ��V(���Kk*�H#QEb��-lI�e��%`��[���Q�H���(�1(�
Z�A���"��V)"�X,��ır�Y�1��rIZԬ��C�U�TK[,b�E�nd��lX��(�
d�m�Q��EXV)b���2�\��p�T�u��gt-�J�p�[�Q�hVY��<X�L�M�ӯo1��BI�ǉ��K�XY��v&�q��u�<H��b�S���$���M�=Z!]m�ʗN����:���٣�Ez:~Zkqg�ͻ�,��0
�\7Y_p�R���爺��|̮�Xq���{���;ӵH.�v�|����%�wU�=I%�4�/�d8k�o�u��V�aK�t|�&�媎���wO/�e.�2�~� �&�,�v�S�T�ځ;Jav�!\qd].˴&��u�N^ky�
ӝjp07�\1��hi�).h��!������6�ڸ�<T6ݱ�:/�泓4lūh��e�;��5��~nt�F�}��a�H@���d���T�{����>`wi�7g:���Cb��<�� W_:���c����̱����ލ�˸������p+�A�e|�8g�/8������m`��e��o9�P$<�S�A��O��K�lǿ6=�g�Y�0A	���xp9�L���V��ث�c�˄�{N�S�Ĝp�M�k(^PN �{�-����Є����㳲y��/���9�vL��<2�uS�=�6l�Gn3T���.���L�(S���f\�f��qX}����h]������m,nk��6��@������l����pn�@�\�>�����m�s��( �f��Ns��[����Q�׳ ��R���sY��Q��V��JjE�}�R��y��iY�ƭ�^n���z��#+�#�H ���Yӈxx*c1����CJE,}~�DO9����V1�-2M�n��l-�鄖�'H�wk����{�}X�T{k�9(HZ�XHiu^젶Ge�	��v�ײ�n@B!l7�w1��Ddj�(L���7`�c(�$f�hTA[O�����)4�&��s5&D]Vgv�6�c�id��{������<Q��X"8�����->^���v
汅V/�q��=�W�ӫ�T�#~�I�^4.�'T�n�R)�'T���\*��Ds�5�~�GUr�c�w����t���7.%!���qP9�<Z#�ˠT��&�Z�BrDL��;��R�m]Fm�ܤ�Qc��R\0���a��U�f�pz��I�$<�; �QFC�cl�B�v��y�
��o��Xp�R��:����U�_�倧�+�uxxJ��6�NCr$�/���d@ܼ��e��b}�x'3�3�k�?/M��F�����@
�e)d�sq�CGi�	�eE;�W~��.��)/�v�Tr\�ft��(�d�7�s�]�7d�o�{��2S�� V�ou=�w��C��a{�܈�1��e�@�7R���ք��ƻ�S6�VG�ze���n�I�V���WP��S!.�,R�Lܰ;q����Sdڕ�p�K�+�l�O����珅��+�ԥs��4��j�|{(m=L(v� �؍���ڵ����Vʵ���R��}����C=�yf�	Y����o5&8�原q�����v�uݪr�C�ty�����ʝ�oٗ���]7�,uD�fVA�t��L�䶷Vz�/޾�L���|*
�.�(F�iXb��s����HQ��lBÎʢ��cOTl�=W�-�^��L�S�.�yPרXCM˄�܅�]-��zuL1U�Q�,��*�e�'�)��2���bۗ��]pC�<��|���3����ܾ%T�Z���&�5���Ws�eY�V���+�'�
�T)�ڝ�T�qɜ=���MOb�VF��8%��J@@#��	���]pQ���~�
�>�QbR��S�y�I���5�q8-ҩ	�D�`����9�H*���j�l.<ˋt��)9oۜ�"-0/a�&��t&F�Srms�Dj�Rx��a��"�J0�&�P�9�od����8*V��\���z�	Q��q����r�jU�b&6G��qo/o������Λ
dc,�bPX=j�I�>�8�b�+�S�J�5�0@�y��} .ׅ�kԓ�uy��t����^w|w�b\+p�d�s�w��ک؝K´�����7�wP�X<]�B7�Z���K�<� ���f�3�`�����$Q��umc�&:(4� �O��7}7j�U�Rn���E�ۖ=Y�A�;]4>�rOaB��cBTe�FD!Pڠ6������B�����]X�u�|0 �'���0�9eI֪�m�U�����ߧ$}~߸ejֆY~��j�G����Z�8k�za��!���8��x~ԩ9���_W<H����͞����.J��)9Y��*�,��A�S��^M�0�W���Ǚ��7�&׹�}Y�g)Uo_�ۮu�H:���_���^s��*��'ډ�S�>|�CEiY!e��7m�F ��Vxи��@7��u���� �v��'�F�7�ò#�ܣ,\�IG)B�z�&!
#& =Caq������pY�H���K��[��釒�t)�R��.Ӽ�l�����h^1��>ȯ�R�1�˧ݕC�����,�F̘!�v��j)6�.�Lc�Hh�u�hd�"�W ���3�S<��
p��8;�V�M�R{Hʙ.�+}�u*��w�1�㷝���h7:Sd�����,kv)X��*_]�Y���<k���i��]< ��K`8ܩԇ!W�����E�;{B���.�mq/u�s�U�Z��]ȑݢ�k!��\�e�w#$)�oR;P'k�PImێp����d3��5�'j#�H��d�)�0�.
�s�]z��|�����. �arj�7�w!~�:u��f��
�;�E#��K%f��v۞�1�����\_��� ��.�S	ꯧ�g5i�7����z��Bꀁ�lsn��c:�~�r^r��_@�YY^�
��Yi�����uH��M�7Xh�s�s��G��)��eg��� �,��j��x�S0 Ol��̭R8�|�5���n���㔍C̭;�؃�H�fI6�u�Fk��	�XQ�9W��n�N���\c�u/�C#i=+R�ݑk �o�*T�	mP�u^��I@��`(da�<vj��"�ڈ�I���t���X0��婺�hfy,w��I|}��$<ٌTʠ��b� ��0���JI<%6x�sr�MK��Q�8`�{��x��f���zzv�m�ŵJf�=�C~���_\�K��[QIof�F�
q*��Y�,\���}�<L�`W8F�<� ןN{S�3BU)+�b�2�*�U�9��3:.O/�x�`�~c����K��G��ߢ�<[��M�pP��3i1:2��щ�;�q�GKW����&�e`�<�C���Y]�Ky>[��ROb��D�<9�U��f)�7;�w��'7ki��e&$˶��|�z�d�d7�ѥ���ew@Jb�!d��\6��=��ߍ��+��+�g"s�e��[������
��G&�Y����q:ި��;�t�i�*x�'�8��uW�|����ҋ�x�\�_���Y����N3_�Ka���8�Xs�ŭq���s��A0a.:VV�]�Q~5Ʃfp�Y���s�_H���+K�n�Z,<*l�9�j8\3H�
��Z%j��1N�*nAM��w3�;�Y%�JBəy���-!�Wi��O��z�v��2��:SV6�c�\��ż��h�ZQ|Mp�/�w�e���<����곸��K n��1w��^9��	&�;l��Z�%e,u\�{)4��^��@뎥�.������"�%:�-�CP,�SשL�%��Xz�� �)]`��j������]����[��c���B ]��9��)C�1�{�F�~u�v:I�"a
vI(!h�J�Ð9�`�r�a�]��{�y�<��d3@'��]PN�FQt��B�ڮ���9�G�� e�v���5���Wζ��+�[ғug�V�^�]b�{97��{Y)2���p�$�{(
�i�{��*�v��������2�ݬG9�.>T�nN���\;$֡l��.P=}H��e. Ս������]�k�#:�ɩS��Nk0IK��떚%r�zp��,8+�l�Szܭ�Տ�1�����}:�*��c�j�+���;��6��lgM���%����U�C�a�,�"/l������܋9K�B��&;e�Ԗ:��)�BL5s�Ю�#Y��X��btV�������;q����N8¢jG`nܲ��y#ڏ��î�흱:�A�.�'���y%�ͩyq��.�fzq�rz?����y8 ž^'4����J�݊��޺��O��+R�b�=�M�[�O�xO��引�׺,S����i4	w��R��^�KN�ݿy������Y�b"��\����Q;]2�X�om�ɾǙ���:�'�ΙTKku`�3�}^���5zH�Y����+y.R�6��L=�H��X��"ۋ����Fȓ�j/Po������kP��z���sH0�\,;�N���`ᅂ2��F^�ƚUhq��v%�:���f�[�
n��I�����}c�T�oռRv-�U"4�=C�2j�ȏq^�:�Zֻ.0�LO<��rr8��CbDV��ͣ[Y���<˩<)L��}|a��ru��1�׌ڗ�3>������+{��3,�'���Xj��mu�f���Ws뉛А����_Nÿz�E��V�ˡ�Gr�'}ѪX9�����E���9M��f>����7�����B}�4V} ���s��<���.�(�}�0�²A�cf��t�q{??�t��@��E���F�U �ق���]P��/)nU�b�3r2Y�]�F�s͞j�7Bk�u��p0�4�i^<�L�(��Lpژ�沞�����j�[���"z�p�����/~�O(v8.=1��̅��A	7�2��.;z�xob��1�b��{1#c2:P�Q��Ni����"LX�c;%z4����\�Ī�}w�݃�g@�a�象�>ǁ��^���Z��t/ø�^�,��#c�l>��w�	vX�l!V(WpGM2xeʢ�֯.h��iB���8[�m����I؈t�/�X��o$x��-`^��@YG��L!�2��qa����쫫S���를���W3���Ҹl�(��`i����vs�&0Pc��.SQ�<m�k���|*�˃�*��r����v�d;U����uP}}Bk�V �vH�m��8��<Ӎ]vu��,��y��ЁT�,��^A��f�q�ɴҹ�9:<2�`{3q�D�{:e���ԭ�g���Zww2u�'ԁ�}��C��%�z��{h��]�^1:�f�����d������8,m�u�:
�jꨝ��ү
��S���i��z��;[{�<��|!
Ie�kَ����C�3UBFL@mH;+����N��W��:�N���cF@�b��6Y���=�~�9��7�Ь��KK�xw)I�Fu�,1ȥU	�/��O��g��ۼ��X�r�5�����*���[B�rl�N8�+��OHdQ�]��ov��H��#����X���F���7�P�sNx3����+��h�Oц�u���>��PS�.u�S�@ÃQ�UHVxi��u܅�X�֯�{4�zC�Ƃ��ZΜ%�gQ��0�֖�?W��T�]��},�x<��HL�4�N��{�� M��G�r��m�p�1�Tt!����@}"���X]�	v�tv8���k�D��i[�2i+�LD��'�5����q�=`;��|��92�Ѥ���Dئ���9*��3�^�#��;�5�A��)ht,�r刯?�l�?�IAq�N�FQ��(�(3�*=��Z.c��c�����8�7�u�|եs!k���]H.q���%LN<py'��*6pW@+y���)Ir��4׷[kr�l}��(�"��ݗ|��\��]��M�Fq������u=�B��e�����[DiRK�g+o>#�fIm��tEM�HQ�M�������{y �J�:��c��ָI�H�{�ڵ~}�I��g�QHǟC%h,F���WoackjrO$�5�r)�{�j̿���f�t���ϫ\�H6c7�A�W1j�t�v�������+i���t[��Z6�����!֜�Y�'��8��E�&=�N�/�$aT�*�LK{K����T'E����޷o̅�}T�X�J�p��xT-��:I�8�B9�65�Ӈd:yy��սT=��p�����/Ԣ��Af�;g���Pخs�!�#��_g[���tɕDk��+�ڳz��Z�x\+���ߞ�u�t�0e~�9�q.q!�����?���t���1��s̗�M͇��c&E�:z��.�{�05���^��O%7�*����V+����+�ۮ�o9�cJc���V��m�e#�&4TB5�2�T{����C�z�"�ڝ�WK:ФSڤ���+������F[8!�N��^��>?��.�[�j�V��oW�s�σ����+�whL� Υ Rֻ;e���o����W��l�Mf�fl��{z�3V�O��.��J�ʸ�`,oڭ���5�^R��4n��P�<�#nY�
�M��[�{�lu�+E����u�q@���gL����q���8����y7����CHa�7j�t�� ��,=�����o�p��$�Ly�Z��	v�1�����63��v�#/w��BnIf�v'��k��yTل5%	�d��Uj�՛Z��Ю\x�;�kzp�R�Ǥ�h���/_8�5�r3i��oz��u�������ϸ,�u�4��L���f�h�CN�	h��
]6���:��[	N���`ӫ�w-v>sP�>,B��R����l[i��m�M�ͩ�5�+��5y���2��w�:�������.��܇C�n��b��6�43K�#��8Ů���¯+Xy:�$fk�]ˡ��	����u�x{�Nj����.��CP�#u��2�,�ts��o�T�H�k�4i����m,��@ȓ)o��a���ξ;jsj|^�����O�Ӄ�6���w(�<�dyM�n���P)ܛ��hn��PfM���ZC6M�c:�U�D!��I�ռ�N�fؖ��
�7��6�9C����[�D�É���S\1Dh�:Di�;Neu�q�st�V��/*���M����l�H��4�b1�߀�L��)n�@��w�9�����Yۙ0�N�1�1���T6"�L�ß�i��.(���1�B;b)FWqT�����ѳ�9�Ӈ��@����k���'d��:�	v��VJ!,�[C�����9�����5�ý�-ӫrJ:+�z��u�Suˠ�3N��)5�}�rb�v��Kꋵܔ6vj�%L�kp��jx����*0���8��R��W��76��M���k�`���&�zWw�ٴ�m��B���7�������;�A�\8��o�{t���������L-��Z�������m�;���c��7��r�LZ�������j��B��3,��o{b���t�ٖ^�7-TV�i��Fk�nR�a%!B���x��(�Ch"���v�E��Soy�@3����)awA�
f���n�zo=ŕgsdo�r�`�v'χ���}l�swZ�RI��j�Y���]ak�)a�Ϫj_f霮���HƆJ�+,sD�y��ϖh�H�]��\��w�����}l�����6�\��uۖ9���8�i\)��8����v���Y2�J�75�R�(�操���N:�t,�=gۺ�R��3`[&����]���C5:��Z��U�����&{Kj�f����[Pf�r����S	�֑3k�x(��&�!3˲�K���r�5�W�]�#��]�U�(�Գ(��Z��¸�&�r�r�;a�zQ��1�=��Ѷ�)qcF��׏l|ڨ�8���.�(�����
�nSI�b��M��	��'^f��{���{9o7�Y��%�rQ��&4@�I��KD6n����3�#Z�;9Y0ҝ{9�mH��կ�}F����� V
Ŋ��F*�UZʂ�Qd�%�)EU[h���Qd�2T& VH�#�,dd��AX��h��+,TA`�Pn\SUE�2VEc`�L�+PDRQX1F��EX,�B")��XT���Ys2 �+*���"�d�-�QX*� ,�
�@m�X�m��j�����V*�H*1dZ�A\i�2�`�����,�(��P���aD�X�R�TeHU`()�YUE2�iA@U���6�V*Q�E����H- �2��*�R-�*��RJ���X�A�
%Ys((��ȡ����U��(�b�"
����,�ȌQU���*��H� ��2�LIV2�T�VE�*��U�Pb�����eTH����"嵅E�X(((
�kP�(�H�*�)(uB�k�h��\�7�w�%�T_;������BJ���Q�f,-�Gd5Ĉ���A��7б��A���Z�U:]pԳU�w��P�%Z�����(�|,���������AT�["$��bMP��C��ߔ�0�1 �e>gP�8��b��a4�|§P�������s���IS>�#�x�>�;>��BW)�m��_�n�i����9lRm
Ͳ^����d��];H,�{a�P�1R~J���N&>��>a��ex����i�?eg�1ɧũ#��G�>E��}�u/�|�#���3�y�=��x�x�C䃪��<Ag��M�u�O~B�?$��si>B��U|�w�<I�Vs5�W��|�C��4�į̕b�Rq�*|©��h������8}�w-Hߺ��b���ﻮ�C�6�O��1�s��c8�����;hx�U��i�4��V��w^{@�bt�O��~O++8����C6v�VT����e�Ax�2g��5v����}߮�3O��{����.t8��d�8�,S��qX��~CO�>C��d�C�+��k'�LH,�����Ӷi ��u�����l5̓N���ܼރ�cL>���� A��#1։���E�ݼ[B���u0$���$A@�<	�?'Ol�Y�J��y�`q%&�1:�Cԗ-C�l1'�Y99�4;�`bIw��x½v�Y��$�T?3'{�t+I��:�x~�f�g�t�oG�s����Ϝ�c%q�^Ͼ�P�����6j��>f!�75�Ă�:�M�!�z�$��b;���$�
����E'�+�����
��T��d񇎹d�4�=9Yr�n#j�1��_�� B4}<d�4�����&3�`,���!���&;a��C�>q'��5�8���aߨx�U�n�����Rz�xèb�C���hJ�YS�������P�'O�������}'��>C��|�<Vq%��g{�i����?$��Ns2J�m�����&2m�d�Rq
���Ǻ� i$���l<�M�|��hk��v�0=�;�v~�J9���j�\|�> �=�����쁧�P�����m�a���/�+=g�b~C�=�siP��N���� �!���*��J����iI_S�L�N!�m%�S٫&$�
Υ�{]�K���c�{ JY77�X��b��/F0F�|G�=9�fr�0U��e`�Q�w٘��G'��.[N��
՘�]�V7��e@T������,�/'�Md&$�'Y�ڔ�.n�-'5m�[�#�Q��R�S2���cs{2�7wk"0�Mo��5��A��SZ�q㤂�k��:ɴ�c1Y��C
M��:�0�
�{�<C�u1>I�c�y�@����o����m �nO�d��!�-_�*>~I"�Z��F*i�W��'F�9^!Vve/�:J��J�L`~`(i���9�$��N0޽�O�����i��7i�O�O��C�8����\�a�'�����#��֐�S7�:=�ߦ��>��PĂ�YĝB���/>Lgɤ�4�Ԭ��<�O��1�Cs�!ė�s��H/�=9�h�hu& i/�a��k=d���(b|��`�|>����Shn�����ޑ ����̝>��|=���x���y&�M$~x������?C����UH/����4ϘbbIY�:�r�׆�d���.��h���A�x��3�l�{��>�G������g�Ȧ��J�O�=��6��P����h��u
����'���8���2���HL�3�J�3�C

q8������q�Ɍ:�0�>�gG}]b�l�V�pG�>��A~�P� ��}��Y�8�C:��Ag�f��)�6�N����M���7��<L@�8�Zc
¼��ӌRT%x��a�Y�J��;��������y_���۝�k���>�$����z�w��ځ�a��a��m ��3)��>�`|���>B�ý�4�OS����@Ĭ���O��t��HT>I}�����tҋהn~��x�,�l�#���Cbg��H�u����2èi>d��n��T�B�����x�Y�'ƻ�<d�i���39��L�']3HbJ�����{����o/���s��J�����}.�}�"�}���>��ϙ��3z�CĂ��xn�r�ă��0ҳI+=�܇�:��'��[$�P��a|�*O��9N�k��3��q'��:��G������g���.�����i��C�v_�Ғ�R��%M0��q��I�8�Ɍ?&�v�$q��|����Ă�nì��Hc'��Az�!�>�hJ��|捸��N�Y�{���}�ǜ%�7Tfbhi�|-V�����3:�V-c�R;�%i���ʈ��ߡ�:�Gy���T��3/;���}ةy���Չz�ߐ��wfb�U���9G�$�岁8�o׽r����hp�[uj�=�s �X3lRQo.h�N!�~�U T��}��+
��'�5�|1��J�,��+%C��
����1Xy�1'�������������=M$q�]$���Ϭ�g��G���_��	�N��n�_F���Y� �0�N�����R��c1�x����k�*AV~I{�4O� �G��T�IR~N�"��Y����T��n>�̀���<��G�DE��3ն��PNf:�`c�M�M0:r�:�~���4�~�4�CG����m �I��!�8�3���wD4�ϐ�y��$C��CI�m@����CR_ >!8�#�X������S'��{վɴ�!P�����-`):�7tβ_/�w�:ɫ@���=�	�q��C�s�kF�'P�����$��La�
��hC�La�w�u>M�x��Ǒ��o6,Gf���A�y[_/�ϼ�IYP�8�3����J��_��X(J�i��i<}dĝB�=��W��_rqaXW�Xo�;����>�}�=d���W����vɧ�I�
p=${HW�r���q��ݺrduO�;
�*>�>,�|5���>LH)봕Ĝ�a�VM�I��՚H<�u3���� q+<=�x�<I�P���
��y���'�bA}���<:��l�&3�޿]�ϴvV�f�N(���=��A>|���ﾀx��T��f�������Rbx�`T>�~�i����d�՘�2^Rq�l�� �&�~z��*�|�C�?oF�8Ρ��������`��5D{�T��^ucѢ!��*��a�8��bM��O�V|������C�J�{��M��s��1<V���04��u~@�!�%ea���P1�d�SS�q�I���#�e|:����:ws^?Q�,�a��C=��l
�!������>M�u=��4��b�ִ*���~O�g���8 �Gw��&�:�'��I�̘���Led����$�#����[:��)��m��3s��|'�|����|�~d���ۉ8��b����1���O���CL�}�:�'��߻����O�C�ـ*��V��<H/7{� ���� d%n�;�����e^�ت���gn���Fr�K<�:7]�ju/mn�Z�47]��Zb��I.�(�l�~Áp6KYyx�'��z�n'��|b��;x�Ny�۳c�KwC:̺��Uꇮ�^���{��䲜|su=t��Ѥ=˾��S���kc�>ȳ�z�I����Y�:P��O�)���L���1��'H�u�۳�a<I�*q�Ý��OU���/m~d�c�Nv�I��L�4�b>���>��<�g���f>��&b�������^ʐU�G��O�3I�v�.!�|�3�cĂϙ��n�'�1 ��0?0��=C�,���b���~�����;�<N2bO��v�$ז�;����u�u���#�G_:`�$��}�	���� a�������Ԃ�d��0:�+>d��aRq?&0�>՚k��?&y7��*i ��P��C�x�0���'YP���gه��
������r�	ۋY���~`�Q Q���2�׬���gt�aU���r�'�T��÷��%M��*9C��*,�h��B�d�<2�X
N!S�t�'�HT>|��$��Ld��~�����^��:~u8���G���@Gß�CJ��+;�*�]���0�m��a���4x�YY׉1��}�6��
�w��3)1I������L��=ˤ�E��S�|d�8�O��{Di�k�l�H[�~����xp�#�Ɛ>K�C�?~�A�J�ɚ��P1��%퇓��_Y�AVM������1 �w�<���1���چ�i�3s���1P�%�
�V>ChaS����'E�/�T��ߗ� 3���p�@�T8����}���k�O����������ԝ4�*�Wh�����v�(��H���TYzP��p�)��NH������M`�MOH�$�@�{(<��/�J��bV�Y�#�>����R�t��r����:z��V&g�x3��D���8��R�گq�[�;-�~c~�'
���k"�is��Q��~TE��uv�����4�ҥI�c4��Bb�U9��,V������qqf��r9o@Dac�x����6B��5��B89�}�yK�䋸�L��4�C�]�PhY�^s嚺�Tt���݃A�F]1���o�:�xʭ��q��g1��t�cA��s��#\q�+=mi���A˦��nլ�g>'U��^�-�G �{�5[.h�I��A�mw,�gܧP��-��b,n2�ۉ^�/���u21��T�97����R������G4�����}�g\�Z���t҅$K#Y@�ϟF��%ݭ���ע�y`A�����B ��k��rn>+��Z>���7�&�ۭ�����P>�D�=�&z�Q�K|Lpwx�T,��!&���u��-6��� �"���]���
�:sp��m��q�˳Ĥw]�4'e���r�
9��S�,w5"�tj|���n��&�J'�尳�t�ai�X���MK�̃�m���\����C�\���������rrVP`7t���Z�C�W9V���^N��s��aQ�?<�v@C�z��pj�{��.����ϛ[��]�)+�Գn�@����S�o��;�w���9�Ȳ�3������j4<Z����4R�{\��ǒ��Ks�o'tT��0|�IF��X��N�ٴL���!�r'�QI��`��ڼ��\��|�\�{�*��	�{�zZ����W�A�H3���:��{R�h������,�.Q��Δ&kY�h�~5)�srQ���v�]l��j����.��:2~�١	����J��p)�TH#�0$�����Βv�bx��瑴��ٜo#��rNϺ:�G��jtDv��FH�T/��KV��Ľ���JO��5To`c��� 8��J&�na6����i��w ,=�٧D�3�k���Z���C
f��}���1\�혍F㊁���g�c[�)װϛ��'ÏaZ�Q�eC�+�<��I.��3�sDv��o�1�y
�s�o:eS�mn���R�+���O��A�t��݁B�h.͂!i8huZ��0œ��Em���ŉ�T��ږ�g��|t��+�B� ���dT�.D�G}O\oԨK��L[�w5;œxa_,����E�%�1�ɞ�� >����Ҹk۫FNrh�]���$9�z;�R��u��>�[�xX9�耞�MX��攻�3g)�t	��ˆ2����0�\�<{��T���-�bB̒�󚈥:�mԊ[�ǜn�n	ʅ�fݫ���H\	l��0PEi4��u�%�X"�a+F�+��cVVi�=�L`P��w�Zn�(n�.��u0-^f�9��eY�T���D���:��Y���V�]��s�W�����j�l�5�[�2�OJ�Y��DV�:r&�i>'��ȷN���� 7����MNP}�ol�"�uy}1�*M]� �վ%E�q<�?S���=9�l�^%Q]3��e��])g����:Hv*ۖ��w�*s�.���PC.cR~���	��t����;p����눡 Ն�}uևb+��;Fm)<I5?fܲ�z{dA�/���6���6;��]�g:8�W�he0��������Qc��:%�;u�-����]Y�^O�xh�\6-VNͨ�������ёRK����a* ��-@�9EIַ׏k�'��x �*X�9;�ϻ���HYO2Fr��2����^��a���-�gk3� ~�]e�W��\�9�|���>�6�y�z���iL��C�9��.K9��>9Y��ʵZ�C�����A��f�����Ԧ��V�9L�*�m��8�����ܜ�c���*�J��a�ȩ��k@�g9�
P`b&�O�27PfeE."��"ko��ֺ��9xa��s�c����Tt�ӑ�̈́�����n���q�F�ƕw���J�������#R'�U���x����G�3�Gn���;�^�s��ɾ��$��7S*Y��d�m����{;l�P[�1����mv�LL���9䪽Ȥ�|�����ʥ�[,����z!P�XrRm!Y���ښ�x�i徜�ȫ�y��Ԙhn�1�]B:aF^t}����7R��75�����r���9@uO��=S�o ��IA)���κ�d�Etiԙ�co����t�MW�vm�f6\��¬�B�U���5�Ee҆������eD^�V�!�b�N��+T�y�|�6sO�n��(E|�[��H� B}i��mz�[5����Ѽ�}N�\��册Z�#�
JxR�IP㡵B׬Ľ�Ë�.�2؎UY��]*{�qh'�jy���3䵭�~�3U},�ΟF��j�^���w*�6�0c��[�o�F��� FTt!�/U��\�T�B%av�.�.�v8��=+nX�щE���^Oy#��]�w^�~���[̂*˘b.	\v�@Zm��-������[��Ք�B��jb�[X�B�b�����4[�E�\h�����=n ��v�(���vf�oor"�*.�i��IqjuG!�)	�\�ȴ�������{q$��ᮌ�D20��͈i�ZǺ�G��<�V�]7�qxb]�B�\[n��@k�y	�����Pw^6Ր��N�n�F�������H�%^y�=
�`�%�c���6��+�|���U󾙴��9�e��mmW
Lw��k�.�M���^0�L��QetԺ�s���!8�d�֮����d��x�ͼ�`�ds|GR�\�t[���{��w��꯾��L�NFxA@e�6�mp�TlX��)�/�i@v۸a�ڄ"�:�4J뱱FT+���S�x��S���(�=y5�������}I��@ًWȐ�.x����x,M�%Q�6�'.�Z�����z��uls�9A�נȾ�6kl�b�B�O�L���j��<�� N�$�b�M��g�O_rtf���zPD���{����/����S�t�K��R���}'��~���-��.:�\T[�Ѳ�l`8Ճ`]xo:z�=���>�Z�8;�ն2!	q�v
��Ldg*�V�Ī��N�Sۅy�\a��8�d��3�Ts��j�8v�ଖ5���&^�8K5�J$[��`Lcp�i�7�f�ku�CT>Vl��1Pn��;f�P�Q���������Dm��"��T�\�S.T�!�R�Rֻ/ݽpD��a�C[��N��iRDz��a��	ر��(���;�֧���%��Dl u�R�����\��*��l�"Cn�{Q�C�yR�� E�9����G(22@@w)��C�Y̍�y�5M�~�$�ړ2�@��,�2��oP�����H�v��u�s~+v�Ru��ᔛ]�>��JP5�h�2���iwˮfbhn�Wi�[\�b��֞���;T����ô����o����B9���ӭ�֪k)+Tp�U
����  ��1r-����;>���B8��K��+ly��9��u�Z�<4VQ��ҭ_l����*���:��L��s��|��`gy3_R}LYsh�9�����4�`�!T����e�!����N�-A^����k��趰j�Z9JB�s����מ��*T���l�mnU�9:Iq�,��t�h�I��n�s��t8X#p���UrX�B��6�Q=��Q��Hozl���hZ�d_o�FA��b=�%,y�vk�Z�ag��� X�I�j�Tӕ�U��4�*�h|��t��(�bA
��_�<��9:�3�����Պ��\�wjX���B���j�EҖM�9�8�W3zdRR
��N�P�lz.8��ݻ�����j������K�gC+u�J��z��a��V����h���+��[�ٜ��������=H��'g�NyV��c��?�q;`�Je�Ϭ��M⿭v�܍�Kَ�瘳=��)j
���������T�s8��շ\OTPW�Z?6��Ώ��x�d�3qt�)-���̇UM,f�Ʈv�UǎsS)��� ���7��]6��"��$8_v6/fs�nИ{z��D`�*�!-�F���Kr��������#�,�7D��ȌD��b]����|i[<�j��x�~8�l9ro�Tδ��)����J�.�^M�hD�Y{.�x���e�=�ڋe(&�l��K},Xt�Q*��V����e�H\�Ŏ{ji{':�z1w8ʸh�,R�=f%׷�]i���	z��X��9�&YIj�We˩�{��#C���h���K:�VԤ5�~����MB;c�tvA�w������n���\�GXJ�ō�M���!�,��n���X�w�~���x�WX���t��b��׫-��Wc/.���Fwm:��v�a�T�]m����[%�����)�o���
%�ԧ��H�caE3�=/�ц��̤Y�9w��:6�/, z�9�l`�+�*ӓ�Q�Ov\-'��w�^;-�Z�G����8�{y���raWn탍���Yx���n_u19NU;DJ�4�v�TҴ�oG>�wǶt�ζ!�;��K�#8˖��
�}�p�O9BNx���˝���`����}�Vtٮ���g-\5�iϗ@nT�kd�ly���,�k�\�=����h34���s����G$م�����v��C]"��������:7���=�R[�P�;YS�q�ţ9������;��o��
�o�k�&�]�a3-T ]�����9|���+T�!\ �Vvy �qܹ�a��V��Ѵ�����V\1:{B�:4�n�pr���)[h�~W�N��D`c+i��u��Ku��̫���r�k���L�s@;�ǲ]KF�WZ�ta(ʂ�x;H��͗���&*䍶��vtvF��/:��}GE�)��+���G7-�/xF�u]�-���-G�8k��e�w���g�YN|��,� \3�E�eMǠW3�U�+x�����z�K*�|s�N6Sj�iѧʱe�8X�:k�d,�x<+0n6�|�G���PN��Z��%�&[Y�(�n�Z�m�E�4q�P�A[Y���؇'ؓ�*�t���@V�=]�`����~��Y��N.wo4l�Tz%���f�K��hw3J�������oȤIv*R�q�k�P���ӹ�>�!�uLX�qQ��՝r�Wsu�pH�y+Rfw:����j�2æ7z��+[w8X�npޛ��*4B:/1��As�nՆ�,P�~6.�\^n,�%cY�N��K�ф����j�ʎ>���[\ y0�fod���i�pH�U�I�����Dr����(�����r�es��t5�����d
����S)�޹�3/��Գ�k�MrqF�@G�ڛKNWh�f��������C��J9�@X�I�#��!��M�^\���T�[�M�{D���k*o.��:o�?ky�υR�Fѵ�X�QT�H��Ƃ�T+XT�Le���Kib��E"ʅA@R,P�T1���ejR�6�"E�������X�T�@�)2�b�##�����B��j���V�+PX�Q���V[l�Z$�ED
��SEQH�����cR-d��AE�(��`���-��QQE�+"�Q\eA�����F,U�UT�1QaP��n9Q�*��5*J�"֠*��`��(,Qb+�V	j¸�Q���ęeEAET`�e�,��� ��������Ld1�DE"����*Q�
*�ԩ�(�,�amc
�XK�DP��*��TDUT�1�**�QE��ID��Q�AEP�"(��A�@EH��콓ٴB�؋�x�ݒ�����ﮕZ�N^���R/����o��u�Z����w�;��'w������s���ө56���X�U�4��ؿL�11��T-�#��s�tK��L�`�!�V��pN���<�<U�|0r�Za�,eB��a0꬜�4�&�<�}�.��;���g����}zL�`BS�>����v2�����k�47SI�(������!ǹ�[�"�' �y��%ʊu��v���R-���pn�\\��Ԇ{��(7�?����w6��^ec��O�0e�1�ѭ
q�UW��<nD��íRp0�4�k���.�.+:7lvX�8����)�:O���R�s�l!O@f�'k۫��s�;^q��rT\�!��<�S�t�}���'���Uw��R}er:LG�z|��E�i>�H_Y����+�q�(�-	����M�8���a7%�_�
%�.A>�>ft��z��T�ڹ�^�q��\C�����}����5B��o,v��f������nꌜ4A(s0�	K�]yEj����R�M��Z�y����P�W�;���kU�wL��2��~�,���Pv\�U��e�2����{3'\�C��Yܹ6�b�<�����:f�E�;[v<2��)�#L�7����ZY&��c'�S* �7u���:%]u��:c'q�خk��L]�9��J��Δf��Ԃ��ZJ�k8j��ڂv��=�Y�2��g8n^����.�������< ����kٜ���N�;[{댜���½@fܺ9��-K�_d���f���y�;ܻ����c$�A�0[V�.[z�!�R�W��W�?\�:7]�H�hkVb]���\4���c"�hi&�X��=�@�Qꉵƅ��/9�{�����@L:3���t�ړ��ky��tå�ò�Ar��V����2@���\l
��N2g�+T�:As*�k$�v$�!Lguv�\�9n?�����Yz6�������<���PQT��"��G�Y���s9�4�=�:[�q܆ߥ�8h�ι6:�H���V�Q�#��w�[��O��d�C^(P<k�^뇈�l�i��q�P�sN���R�ŏS�{j�z��lovY#I�Nd\�~a�f���+����Xbw��hg��u����'6	��7
�l���#��k'ai��=�&6T�-kmZ��},��^�	�զ�I1���&�=<6i�1rۑ*yt?w�ҭ�U��5�(���*U�q�4���W��B��c����ծ���k�
�0V��$�2;�{C޷m��QV�wN���L�C�cJ�o`w��Z��R�.��s�����*�yI;:���"�k�m�#��/w��+�։��el/��\�g,�����z���7���q����A�k�"櫙���c@
�+7�� {�wv]��݅�=:����4E�P+h
��k ��\��pJ㤀��[�d7�9N-�c^C�j�1F�������f���VrH��I;��4����	�X
=�4�.7�_2�NQ��k#�W"�֓���L:�DU���î�`v��u�T���q;�B��X޳�Us[��o��D:�\��T^��\3�"}���X�רr�<b"��8̫��"(=Ol9�cu���B�&��;��\=(���QXb���(��/6��_FH���rxȮ�'#.k���E���Ѕ:�x�`�h,��G��>6b��A!�\�4�m��ZwX��W�R�·���}L@��
���#������_X���[���9�yL��Q��t[��ɐ?Vtc�����5zq��]o��j��߶��9�h<?h����F�ї{������,��)��}e��U�Ѕ�s�����]t�x��n�0�F���T��v��+�wo�t�M�U -*��2�1p�a3sά<%�j��kM�P,ϵN!wL^��fw6*t�GQ�9; ၬu��NLJ1"/�]`�;�U��6�[!V	,��{�N�
n��2˝uwz�S2���`9G�O�#;�9�q	
�`ku9�Ӎ�U�bx���{!��4_���B�-J��:���U�f�4T�+�b;=����<<���ۇv�u�P�����,@W?��	��#-h�N��F��^u➪4_�����!
�-"��w �wSRu;w�ȼ��R 3e6���ф��,��E'�xͱ�֨�m��sS�xNv�+��1�Cōkt�3am��P>�P�{�ge	], GV�b��4u�ɢ�q+z:?�vC�H��+�,���]Rl�.(�.|��Q;K��rn6�.]X�u�\�y.E���;�|�&���K��g�x�� �ѐ���Q'�����qѸXJ��
޽�W��;9Ȁ[;� Vw�5�iT0��3RnH��p_>��x&�x�}Q��]ei�)]EN�\�dm/W*jߎ���)
��qP)��Ց5sO8\_/3u�T��&Oݱ�v$F��D��\�=I���5&+�҃�J�K�'���\�Po���k&��8��b�_��|iuC�Y!qÓ�Qs�aa��c\�2���L�4�9-��6( ��-��]%�M�r$���g���8GjŐ:�<�t�z1-�'��q�g��-�MLW뻝,ct�y��a��'Z����a�z1@�㰹-��i�<$շ�t�޴�O�s-�L�{���N������C����(�8fu��s�;b'�+7��'Vnl7�p�3�_�mr�s���	�����DG�}��r�>�����rx�(yL�@�"czU��
��v��Į6,k&�����S~!�3¶��8Ý����+؀��gC(n�iQ�z��a����לYj�k���p�1��YH[�Dr.vpRX��氼'\�N����_e�lS;�Y�,拽s0�M=)��Qs�s?1[��%7�*��8?�%}�t�="z����-��4k[3Z5�q��k��_n�t��b�󹆽��`��R\����kF���+xw��f��՟tV��5|l�YC��̡�9ĭ0��e�ף��0��sN������w="��6NB2�º<O���
z�~���yA��'#�z؎9����!����R�����<1�'}|N��D���˔��������܅���~�)�ql����\e*�p�THT��匰�_f���{`[^�G���G����mUy��_kR4�ִ'��M���"x�,6x㵍�{ �)a1b `�4��T�S�3D����<nw�qۇJ��XZ�ZS�}d�[������Z�^i�귱}pg]�h���u'z�g�th�G@�ͮ�Ɨg�G�ߏ��7L�؊Ĵ�.g#
�˹
Y�p�����n7�n'���ݨK}�4V��݂�%�����N��&���{�9ι�gC���m�z��o7�{pa���{����4�N�ې���|d���)�O��7H����T^&�S�t���������k
�,_T��}���a�/� Y[�5*��n+Ѕ���gJ�^Ӓ�u�k,���GX�PZ�a'V�M�r;�U`5�D?m�5��K5���A/4�TY���`��)qˠ��2U�j�x����;o�w����������6�ove��"�4>�}3
�e7��!�z＆�k��uQ��G=�h�|�p�c�ҭc�>���J^����'5Ȣv�Ɔ���|�����ia�O�y��i�j�-�~+&�u\�Xp��BT-�b+�ֳ������!�yL$��W���q���1.�4�vZ<+�k�����-*�b����<��u�}y���4r-���{#m�.0�y��;o��!B��r�Q�*�CY��WŰ^�X&vN�8�ɧwQ)R���U�3�͈�\���S\��s��y���+ְl�Ajt����U�6�����eA*��
��HH���p��M_����)���1�M�p�=m
���9
J��i�D�ɖ(��U�E�ݣ���u�6epfe�I��`�];�^�P�e���r�-��`�U�'�Y��m��_�.t�MZ���{��xW>�ĝ����so��v�rF��	��N�iV�P.f�.�W�������g�NsLUl����Ț[˨.2V����Yl���7N2�O�n�0L�ڭv�]ad�]��Y��&�+�E��q\R�J*��-$wB�'���-c�ZM��cn�F�c��z�R�-���0�H�?)S�h�g���*��ȇ���(~Ǟ�S��&�Ԇ�ݝ�C�����alaƠ�`t�BD.�!�o[n�B��\�=V����06�ɧ��7����i[A��z�n�m��J㄀��
-�nݽ-q6^�S��o�iK6��1��E���<�j�nIK�Y'��]�5�<�;����Ѭӹ���+�e�䣵Ӳv4�.�F0jRDeD.w6nTG9�O�JIL�]ߢ��`[��ڛfԓ��+�`uA�忼�+�N�p�������[@���ՈD�29���G��3��Z)F�g*p�����������R���p 7��0IS���N,�<u
N�׼r�*WO�c��ޟ��Cg�#KAeu�#�uҰB\��
C�=�sV�Q|A���r��tݨ�ݾ
��'/��)y��"8�[a`����Z�	���Cr��Ny|�����E�Yo����.m7^7�{�6�ۥ�o[� GE��-��0F����\�.����Hu(���2�dϧi��U�i���RV`���y^kt�A�u)�V�ͨ��'s������ۅ\^n\��~���Wl5��W�g�:���J�0�������rھmgW��{O-)��
Wv{����p�R��8˭����?1�mQ!h�Ip��5Z�2��Y�`���&G1�U�"��ECZ��t7�=V�w��6'�{K�r	�a���`��ε�O��������edFu���q�	uAf��4���pܦR.�`�A]���hI'�]�<�L{u;*�I�H�L��.4�:�`��y�O�Y�}�xs�x��o�Y�Ǿ��q�j��ҧ� �؄i!������Ȇ�*��:R�07;NJr���Aot�����dڀ���6��W���� A��fL�Oo!��Yh��֝1���2���wCL�wU����e����\P� ���ܰhA����;W5j�3{OA<��)���O��7λ�|}��� )S�d:↮FYGo��upp����8Y����!�4rB��!�Z�+��VQ�S���@��|�#.�������-{hP�3�WS���k+1��� ����Y��r�.�}K�<I�3i'/|�dẖ�;��,���fJl�]p�S����]��n�pG
K���0j�Fk��g�h�V�񊰆W�����2�6+nu�iG𼀎)
j�RȚh��?*��;��\�5��zyZ�x<��}~�@c��f�7�V��ׅ}p��R�IG�CK�"4ڈ�.E���18X#p���������ċ n����ZF��;� �\�׏T�����و������ٮ�j��!#�;P/C��y�D�P��C�2�,��ޅc��5�y�%W�����pȗi�T��Y�S}mMp��H�;�[n}�bÌ=�^N :��kl��tl�xP����l����q^4�{��<�IA!�.�7W9Aи}Q@bڑ��7a�K�k����vE�B�g�(�S<y�����.��b�C�|<�蝞��zd��B��>��tʠ�y�ԯ��&^�s�$*Yu��1�ƯI�tQYS<D5���[g���Җ�c���)��8;e�wOp<Rf����t�����Ob��}tkB�^ө�� �� :��j_uH�&�٪o�C`�MN����dt�6k��n!A�g:&t��O!|:Lx��6���/i6����b����:�P]J鬖���98�p�>#Ko�U���QhQ�&��AXKo%�ҕ����GT�T�����e��v���AL�;2չZ��N�T�V����L�nU�����V�u�6�u-�mT�WTO��_U}_Uvc��i������{��|�E��v����'j�����O*C4B��
=ЈҲ����s��Q�71	}sڞX�)����wU���V�Yu=:!�@B���=�7��ػ��{Hh$��?@L��@�t=@q�S��y�k�4#'Z�'Үr�iB�a���aۤyb�;���m̹D�!�$@��~��ib�=�/������2mH�K�+�/����� ��^^UZ��(���Γt�q���u��O�ҽ�vz���U��3���3d��n�]5ҽF@׮�����F�ÀO��K�|v��d��5i\u�q���7�]7%��9�]hh�J�1p��B�mP���� hI�J��%�2�1\d���闖����)�0S�U�P��Y��s%�8}a5U
�m919	j��L���8�����]?���g��F�G<�z}k)�%���zj�l~���)ֹ,��ek؍k$DF=�.�ى���f���Ն8h���V����C8�qX�������ӹ�53�boLI��i�M���;P��,�r�\4�Z�W8�`+G��#o�<Ύ�΂�1k��l�6n ��|��:W�� �R�IWo'���MEb�R�cRt�g��7Y�.����Őp�Z(P �%���-	'���톆�����ޫ��Ց�s�[���SY%k��3��Z�b�(٧]���]ܮ�<{U��g�0����a�!�
Ja+��݋�Z��}]M���j����K�܆e�.���#���iE/�i
����J�bKcOJu����]N�r�Yc�a9yd"�ٛ�R�X�kVĤ�02�@�L���;}3Q׆�t��U�D ���YiwΙ�24�={v��	a|�g�>Dm>"���P:�;�7kF-�������LK�S6]l��]G
�M.�W�����d���[�2���#"f�
�^�'Ml����%�[om����Ps2���Ôw`�aI�8pci7O��H��sa��f� �QBx�l��Z�И6�&�6��A�]�Gj���u١l�����5 �������ɳi�CS7i^,5�l�%	��DG8Pk0r̻v� 2_r�1�|��=Mҗ�ut�W�9�2W;9B�xQ�f�<�\Iho+��ZmXn�剥�|e<��#+&���jP��ݓ�v�C���I���c��5FᲝ0�6/lC��+:8��5x���N[g%sѣ���5ĺ�-�yx^��s�X�8s��<Um`���0�=��9�=�;��0��b�&�+�z�
�|��^<ۛ���英��}Mؙ۠���;ث]ܚ������ �����x�B%@�}Q������=\ܧy�ѽ`�Xg�j�y�oJg��&fh�͗w����������(�û��F�gYWGd^}]Ӌ`ur�cǜP�Q%e7��,G�q����k/*�I��ٻ�����}�.\�5vR4P�qV�h){5+�ߐ'i�H��uhUk�����]_R̰��n���k.��ֻj��K�"�@&��j�YL`v[)Sӹ�hB���kZ��f�%q��3dA���ɻu��ۮ9F���(6�e��M8����7��nn�m�s��j���ܹ�A�\�,F�����c�e[��F��O �"�E���ܱ{����r����%f�@�H���/k��q�C.+Ne(�0���ڭ�(�YS�wV�w*ãJ��.���3k��D�q`ݰ;^kҬw`gq����d��U�z�2ug�i�0v#��Vv�gA͘�9���9��'w�ChW)�oY�\�����rڂ�sB����F��s�e&$����l&�k-�L�YCP��h�{U�sB��ż�vh�V���3v�;:�LZ��.�R+��ev����˹���Z	H���Dx"<�*ʐ����#"��I�1�E�Y1A`�1F���R(�RT+%H�A�b����j[B�����2�E�A�k�*��PX��"�\Ɋ"�,Q��(+`����P��APT�A�,��# �(��eE�D�U��AB�H�h,F6�E!jZ�Jȵ0Y((**�E�`(�d�(-IF %��X,����f%Uk�� ��������[J�$E �H��,�)R�+"1a������I\H�TX����� ��խV1���IڃQX
(�k-�X�DdU��b��F,PQ-*U*���p��EEcl��1L�d�V,DQYR*�]~|w�sW߮���Uh䜛���ŋ��XW	�\D@�j�8��6�Fg\m��t�ʡZ�&�nm����H|hˋ���ꯪ�r�X׽��D�
������i��v��G�{b�D��k�(_/�I&��<)[��Td�aNU̱���n["��N7s�5�R�*��r�B����5���� �{�����x��1yC�8��3�J˔.��Wj��F�sގ��X�޲�m�%���墥{�j�����VjT��˘N �����p��M_���x��6�ؘe�鬮6��/6j��A��;r�2T'��$��	M�G���PdO�o.���Z�o=��ܜ��b��W����,M��y�Lֹw3j�W����?R�|zpTm����A�Rу���5�Rx������pRV�5���
v��W��"��P�^.���h-�(/ttl�	k[h��t3�)Vhr�=����4�z�3����-4���oabt.(�ꎄ6��bkϣ�i|�YZ=��X��gh�ް��q�X�=K�f�i��u���t,�)�ȟ%ڶ�	�S�BR�z�1�P��#(j���L1�|j�I��\�i�	�$e.4I���=N �"Nu�JLK�S����΢�udQ&����#�6BV}}���	%	gFt��s�3�8h�l�˭b����bT�n�%��c�5�f�WIGKMv�B�
wf�Q�X�+�Yn�pV�00�֦�X���[�wo�X�}�ޘ�&Z���U��Q�h�m5�=#�w����x{�����Ff��F/���r��#������X�����bV��[A8�WVn
�Gs�&#r1��H�BR���`�꼯��f2�(��ŷU^�p ���6���G�{;��i��n��m�0h�6�=�J����Ԭ�}��x����r��f'C}�g(a~���Fs��@��7M�,CY[kD!��.G�'��1k0�Ҕ��R��5�J��+@�{Ԁ�p+�#\�x�A���{u�2/�M��ٌ`�Cܷ~7v>ְ���ȽW��I�)�h�t6`�2�y*�/�2����Pn���I�kJ�.�+�
��f�c���:��65���8j�](�Cx�\�]o:z��wz�`�p�N�Y��9����g���EA=����rS|��w	F�	��I��,,5�r�H�-�$����Q[=ؕes���roPƅ5��1�b$;��`	��
�ƞP��C����C�Η���6�fZ��]j��Y���U�u�;Hq^�%�@f�@�	���ΛNJ+w�9�i���R�̘.>шa��E�@����<x��o
ޜ5��_Y�]�k<�@�����y*3�}�g)N�ú���u/]��oc��ϸM��n`��q㛑�mvuKjB*9�Ե��N��6kz�I1]��-Ư2�#�����_K�g���D\�a��{�߶�ڽL�mˠ�-j=���<�{��=F)hJR��E�c���J�V�d�w�Rˎ*S���"b���d'$o�C4Y��c6�,�y��,l�붌D�}sB��xp���||�&�����kT㮴���$@����͎sj��k5�(r�|����Ύ��R�s		����rf����,��\�}pt�M������UI:���3���1�]8G��m�E�[X5q���b���e�T���n��
��	O�L���P�^��{�Z1��[����X�`��,a�����iO<5���7k�r�����CN�����v�T>{ĕ�N��~��0���$�>��L�u�h�I�**$�ݎ,�}3���' 7"L}f}�,S���X���L�w�%W1ϽEe+�C�ד�^�`M�\4⩧>�0��@�}�=��^T��V^�$N<��W�6P?�f��(m���@[YɃy��@ؽ9�������V�N�G�7��Ye��sRc�`�ͨ���7�b�x��u�׏���:��K,xo������:+U���W�<{+u�ۉ+��tf%�1Kz�KWe�Sf�QF.�7*���UNW�B[���42�m�% �u�mw��x@��Y��eDП�ŐβE�k��u��1��Y�q�9��3S�t�B[�\PבyF���%�31r�M�����>�n�1PQ�c��ʦ��U��į���G�����՗�\,я\�=�n/0�KՙN^�1[�T5갆�!�ؙ�&Vj$�Rj�����t�Rg��buL��J��xO�.h^�b;���&Κ�3BD�+�ߛ�����
�:��vo:���۶�+� :'�Pv99m���F:'�uY�E#�)�E;"bd��p����sa����Ldz<u�*j;S���IO�	�E�!#�.+�3U�7}��E:[gY��%��G$K��T0C�(�mUz�y�x�	��:�jƔ�{@2����Eu�_ꝁi~D^�u�́8֌4k\zJ|���>[f�����f ��읪ߣ�׾x/Ե�G�\��PhmL��9C�L�]˪*}�Y1���E�W��^��53ʲ��V9^\d�3�暴�K�Q.K�O�>ft��z�L�U;Ph��)�ޣ}�t[���vM:9��;�����K	�����J�v %]bq�'K��a��"to������C|��s:����I·>D`��u���|^qX�XDm6M�Yَm��7�5ԫ��cz8#��y�9:�}�1��V#�5�!�|&��տ�U}�UC� �\�oZ�j�_�GE�l��,�D3��Q/��<�0h��)j�j�0�v��=�9�����E��B��\�P�\kz�Y��ѥ��`�r���+9�u'�e�}�2��?�)��꟝�J���<?jR޺���P�3��_I�`�_s]��9\]�H��L�N��Ͼ��Ն<4[�[�r�4�P+�߰�u��f�K���g�Ⱥ�a�E�#5V�)���T����E����.�G�{b�g�ե^�NSȶ��]Uy7V��@��롫L� $z�s�gh7��l�K��.�w*�!DeD�&T @y*n�(�O@�tΣy3>��VvP�ޞ��z�i�u,���Y����LU�]�n��0�ά����բ����O��nHd����T9����,�'Ί1�����ݨɩ��MP�av,wС_���a���F	L���EZ�R1"��}P�.�9~Ct�N&�B�]�u�ޡD=���]D5�D�0A��Er�F.�Jxh�"�-�p��/2�"�i��ڒ���]�W�*����1�����e[���X�z�N���'z-����&�S�(m��
�pք�fL
��uǗ�;���kR/yS��,f�!}�^��f#�z�S^u
��r"���2�@;��V�V6u��ts{0���٪k�2�?=��x�ͳs�f��9���Z��=�E.#���q�]�B�$g���L1}��Һ�:a��,��������Zi��]��W4|#�\6����@�eeOm�)���|�x�њjd<���O!�_���,;�:Ii�}4E�i[@7XOU����P�i�Y7G��q"�V΋��x���;)�蘤�h��3;�BZ�7�>MUѸ��u u7�ȇ����چ�Ft�2u;S�Aa7s��p��@�؜��`H��\�l�6����d,7	$�;y���p�u���M�r[�20ɐ�^O�o)���4��t��{���:x�7{6�֪�J����1���T;��xD�����Z=��\=>5vy�a�"�Pv��q�aj���1��%�6���;CH�еHysF[�V�k1��K[�k�ߘ�zamA ��7؋���0��.I'��p�{u�2��rѯs?e�cm}��k!�<v@Ь0�vܖ�-��T>�����̈́ �}�&�x��e����v�~c~�a&�
�]u�Ϳ3�ƫ	�!a-ZM��nӳY�n�(<� ��r�$���kc��  x�j�\���<�x̮wz�Ӕ���������0�G�������ނ�n�ۺ�:�A��\,�b�w��u�V�12��j#�ꐜM@s��������μ,�	��0���h��U3���O������o���#/�Ξ��8��>x��G��S<��Ӹ%*�.�P}���}���w*�0+�������Y-m%1��U���n*�i��Y�t�Y1���9p�WmNw���f�"��G\�/����-�`
۳�9,�z��or#^���~M�4w$1�8f�$�v,��T뮫�W�x���:˾p�sޚ�m+�\v��8�n���+��l%q��k6"��U�=�as��
k3w��M���ޠ�U�S.P
�u��O)�h)˖�u��f�l���.̿�'_&�����7���W���n*���t�'c���t����N���V�W����%�H�|���l�L�\�gcANZaf��d&4q[��j-�]�#=�V�s��C�]�9���ބ�F���)t-pUÅ \CLvٰiu^b���b�f�m
�r@�g)�f��,S�P0�5�Odۘq��#��5�e��9�Z���܈`��U�+�v�|��yN��JN۱�|`�:2�.Ą��9B�ރ�Χ&i��-��ƶ�ܫ�ȍ`خ߀���l[�m�f`4UVo��C��@o`��k)�V�����4rs7&���|)�+[�V�.{�A���M�5%p��e����ekbTU�z,Z�Ns��.�P�v�|P){�mQ}Y�A�+�=Wq��S�4�G9����|� ��ѻ�'\m̪��d_rs;����˂En7n�kn���3���/ՙ5{ �vL����Oa��ךΩ�?k2��^7�J�[s�RS7���n�[��>=t;�����Z�E�M�=�n�l�n�g@<�8��'*�Ym�۔ޣ]s��{`�����ˋrv�0u��v�T^*����{����4����ж72�m�v��P�3]]�E���&�9''=ˣl�9���Wъ:�|{�V�vW����CW�G]�ә��ɣZ�v��j�\��TZ疴t��4S��@�
b��:����6�`d�����G'G�87����|N��/�{Sy/7��C�Ԣ������4M���<�b�����-M���]���Yz�4��U�4�ʚ/��y'+�L��ܓE=�QӗН�+%'���J�g�Y�D_J`�]lvi��'���xA\؎���+�Zj5J�b�	et���.˸�O^���������<�w�k�Gr���u��+p�ӱH��.�1�b�Z��>̝��$M��8+.W��;��������5|݈�l�� �ڋb��^��.�U����&�[-�]�ZR{>ԝ��4Rt��>gL���v�!U��<���DM�uE�3�<r���T_2�7��yuK��C��{"�̇��T-B�f��d���K髷>o$gaQ���U=�6�9��#yإ-��Y�7q�<�쉪q�ܰ5zq����Nb��r�9���;̹H�>���]\��Q���d7f�Y˔��+�*/f�\�u�����WY&B���Kt��Sޔ�x�t3�^視m�KKj�C_g������Mp*�6�'{����`�^�r��ٗm������f��\�&��m��]n-��e������+��Ĺ��m�^WN�=�xl�o%[z+7o
�r�77�H�x� k�u���Z���Jor��y�d�Ʈ��ś���1���rf'�2o
����C��J\d�<�0����\�m���\���Z��D�g�,�NJ��WVd�VuQά�䵮qDk}G��<;͡�YW��9Є&�J���v5��D`^�niou|����������P���WrZ����J>��$�h��b��pn=���g5Թ1�|�ZVU��:�K���x�(`�c���#�)�v�8�t������l�q.i�����Z��O�D��=-J�7��6��bQ�2b�%����Z�}V)$���c��o"\^�)e������9���<��o�с�Dv䀆��I|8&b�n���q�Yc^e�n�O�+�=�E֝�ݎ�N�Rq�^a�6����K/�9��V�1{Z.^��'�qVRL�&��P�+���$�nr���*U�9��9 ?��G��ϯLS�8��w-�J�R�kn�аMqO�v��#m��P����h���[x��£ۜ�Ñq��"l���Q������V˾�|��M�Dt77�wJ;�YI��]���#;c��-�{��V�%�~or���.�k��!;��ǥ+e5B���v�le�����J�f�GJW�4j����={w#�W�r�A˔��8U�{��Gf�<�Fc�>�P��9I��X�0�(u�JV�w_ڈ��EuFx!j�#pw�����w.n���P:�4��u��3�5�ȶJ��\c��3:.ԕ�գ�86/�\��ǵ��r���|7N�ѺY<�e��-�v9������cm
��xbo3	�:����bB臭��mr���Y+5l�/�&U��:���G�5�!>|�8�qV���L�1��z��<�Z�RZz{<F��&�ڃ]��L��ƻ7����A��W��	�A3W[[���8�g>T+-p�Y�H���1}�-��Y9�7��en2�liy:��>��2�7u%����0ʅԫ�om�!��\wDZw+h1�p��v*�e��W�m���e
�@�\��ζ�v�Suc�����.�J:x4lw�t�ā���71��ԑ`���ÍM��`>�v����N��7��_��.�k}U;J�i�-/������+v8���tA��wA�n��*���ܩWC'z��!�f� ��v\'�1b��6P�������q��6��}�6�R�k��&��Bj���*g9>�(YK�W�sw+P�cB=lw,�����U�����/SV>�@
�<(�;�6��T�b��>mhu��)���m�c3�f@۵|'-5�nt��N�u�/��wMυ��렄�7)���p4z�h^e�Z̉���]�\��7a� ����w��}Z�iJ�|�C+Iŷ�������e9��swr�N�aGt��r�h�tY�;�l��ڬ�K���uⱵf�R뺤�:�m�#�Բ�*r�,��S���\���U:�'���?Iw:� ��� ���+�z�7ź_���P.�/4�����܁��n���R����y�V8�F�6p�)�����ا�%�Kި-.��f����A��Q
{��/B=`�ף12;ja����\
�oKr�O3���}�&d�.vZ�ݎ*�I��;Y���+3F�SU��1)c*!|��7��;k-��V^k��kGgC&��8����6����S��ste���WFg��FćM2I���(6�j��T�d��b4��N�����s����D�T�GX��t� 4��}t����)�Ke�p��NCY��0�퇆bp�o!)�}D-�=\��j��f�-��u�jjn��+\$��Hn�\/�N�k7/����i:<�U�Y*qWq���wqns��[����k%�����]��Rܾ*qX�ujg���ȬG\��<�Vk�J����X����)�FR��s���kb�����PA ��*��h�iaDQDKJ6�J�(�P��\j�T�AE�lm"ԁY�2
R�# FLITdY�PD�E`�VEb �+\J��(�Z�P��()�E�X*��)("E��QT�X��`����X�U�B����R��X���b��Qd���T�
���TQF+"2ڤ*
J�(,����EG.eA�(�F*"��+"�Z���(��ee`(,,"��X��dQL�ZH�E�,X)�TS%���/\{f�W��Z�NQǋy����zo.|+��0��Fn��Sc�p�Θ���!0��jr�B��d����A�O���U}����Yr�嗪H.Uy�VC^Y����htV�̥�V"�zY�˕O�^�ݽ��x*��8 ����{�g���yZ��j�Aq[����ua����而�=�����[��.�������ϥ�s{��3�R�m#�h�e�k��.C�}Y�q{hǺ��k��~o�θ]N�{�y�dkӶ���;5|��N��3imm�y�my�>���j3��~���6�/y���`�⏣I�Qۺ��gu�A��
����j�&��c��X�@����=(��0w���^���ܷ����V�X1Ȏњ�E�]ie�;"��"6��X������wk�_���B����OE7��<: N����)���'/Ss{�G7ܐ�ř��Q��\��br���;ТB��H�4�TG�s������颟u��pW�1ܩ�e-��\�����i�����j��׵����Q;Ҥ?`�D���Z��;J�#ӊ��6��=�R��I�-a��k�w��(���P���*/�0�q+/���`Mk������p�oL���x�e��E����e5h'��x{�n�*N�,��7���U�݅ٗ��N���y�/4)�J/�4�6�r��z����c���hWzk����̸ⲹ3�%�{�SP�0V(����3��v��	��n�SZp.۟<���b	r��v���sSu���W����]{[3!�nB�`��<�ڴ�%OM)v��LÞ�{[�U9y�4N6=��u	Qu�*�����*�EnC��fH=_�ro~���ܦ���vV��M�WR�cc�����`P���l�������}�H�[^��߂�O>ұj�1��g�oV�9Gf�Z�Ѿ1��t�`�߃]��;r�&׳,[��흜��u1C������8���k�<��gS;�{��D�Hk�=������m��=�E|�:�ս�E�S!�z�N��6�{�ק
r_�dK��.o�M�nP�oDpBq���g�5bvn1��L ]�j({P�y�0���	�����ȥS�)��N��X7�y�Ok��8k�����}*,V#��ptJ���ԾU}[t���ᫀh��ћ�zugmK͘ �����/F���s�J �\��p�A��3ap�Z��������r��5�5��g �]E����)�������z`���%���n-�����g��ʆ�D�cU�\�|֖��y�7���E��.��Dd��c�p_3Cu`��־������m����ŭ!T�X'������;����B�����\��U�x�v�O�K=�����H��\g��uS�I��d�S4��W���BY�?��.�?)�P��c�@7iW��˝n<�98g�;�Qn��)F+�h�y\%k���p�j�7s!^`�ಭmc
����w�3p]�T7bU˞WmZ�H�=ͦz3��bw
��iiMFkݸ���u�ӸC�)d8��/xh��[���ܥ�j��3�-i�X�k䤾�mT6��U,�17PŻae���Ep�w-��r�K�<�U;�:�v�9�P���Ę	dX��+�򷒣�j^���m��8�u����Λ����PC��w)<�V/[1ƞW.��j�/:�90��r�o�M�M�Tg.㖖�������N����uE�Iso��F��IsW<�dS�]���Jw����`�ޱ��� O�n���u�%�|�����/���r�{M}z��h��-K�N*F]\�Y7���5�6�VD��޳��=�򾩨��qdi�F�R��Ɯ��cs�<�u��g�y��36�ra��q�9��>�tvv���[����{Z
�8�x�}���ݺ٠��}���圑TwV��sV7�X�^�?1��\�fyQ��8ᠦ������U�罛�}@5��FǸ��%Z���W*e�[wT�Q���%iu�qϝio/9��O�0UObؼ�59���*����mx�y#�ã��e&*�*�T:���~��{w������e�c�4ݎ���Jb��D���2+�\D���O��{S����F~���i�pgp�*�k�M����un�V/%�����I��������3zO�4�)�/{��Z�AB�S�!v��q��x|��p�e�Gvu=�ѦH�Y���k7�SćL�LH���mQ��@���to��i��h%�z����z�.��]W^9x8��Z~+u��xw��hv�Yنэhp���u�X�8KV�L;x�������y���!K;3RyƶR��8�}�U\i���V���ҹ�.����im�ZV�A[P��T���N�P{��n9�p�~�4��6%nMF'�|VW�3��S��=�"ad�{fK��x&k�Y�S�N7l�-��9��s+|�U��8���qz�3@�n�]��ʕ�n��8�d�����$=�*玲����Qg��[1x�r���&����=�;�ᳵ���tV�i0xlm�Ra�ƽ��r}���;3�⣥:���C!���eӫ��7*
�b�W�)3e�W�?v"���X����՟E��5�},׹��C3~\���S��]��Oy�m��|	P��9Gi��J1j7�^�B�Wۜ�]�6�,C��װVS*&X���NէG&5����J٦7�%VZk6����#R��Ȭ�S�R���w�MZ�v{z2I\6�EkY��N�mw��K�xeGe��ߕL=J"����@%2[Ү��xr��f��+�[�P÷�t�V���V��k���Ք����kOn��/��Xk�\���h#}��3���*��w�v"3�Pu�����9rY���k]����|��#3x�������g��a쯼�����ݺ�m�ڰ���c���� ݍ6�=��E�g-��}8��K��[���)|2V����7{F��,��%Qәu4oZ�����Z;�=<�K\v�43��C��ݳ�!��Udaռ��E'���zdr�λ�H-�6��o4+�q��FH
�.t����I�1ۧ\@����U��]�ٗ9:�4��ۘ�R7k]�W�{�g�^K�=����d�:=�]�e�摫�$nr2]ٖ���^���v[ct��Ǎѯ�L�T6Ct:�Ӌ��Od�S=Ӷ���{�OlgmV����l�O)T�	e|��L�6���p��%�;.�4���no�^hV�*�y�q'��r�N��7���V�R�q6WVt'�Z59U3�mg�v����i��ϵug�o��%p�|6[���s�LQ�1���]O��](�:t̹�E#Rmߝ��0�	WW�\��*W��»���{�T�^S
�>������H�q*]+�S��F�j)����7C6��Ek9.����-�$ �M��	�fS���$Z��Gs�]�}R�+�����z��뜳�6�虜v�����|�h�Z�y�O�T;�Q��p$�iv�Etu�V/��:m��3_T�r�����=��Lk�{_z���>�n������K��6��fo��� ���⾂�9�4��׽i�;ϩ�+��u&+_�y_f��Zo.)��ڽ��mD]��nD��HuԵ�*�H�Z�lz3����VuR�����i��y�LF��zT&�ë�����A`�l�>����h^�� Nn����z�ٰ�_��n�n㢫8賱 �n��4��O-�7�2 �#���2+_]�'����ㅻ�Le��:��̰�.tvۍ�=��Ƹ��TZ�	L��\�K�b�w�)w�ĉ�u�cĺ%�nw�:���|�]��N\��f�Jk�����w�.ɛ���*�n������t]a��o�S�#��D�C\	��`�5[Q�ۏVZ`��J�ɗs�����ܤ\1�0n�6�5@�gn(��Q�-D��m�����Vn����d�	�Ԛ�,�:���fi��1�f�9&�*�آSh��5�Şǣ���ĸ�g�y��X�p�7��]�(V��G����}��{=<�xr̰��k;����m���t3V�<4��Sa�xR��֡k��v�}�,�^�u8��@�]�<����$���V�N��5�� <z�ۿP䶨le3�3��ٰ��B[r�[P�`�F1����r���HL�p��������:��x�cV�5��r�n0pq�1s7s�6Vv����|�OϮ�u
Ͽ4��YG߭���}��K��چE���"��T�T=�J�[��8Š�D��܍g,��
��^������+����c�S��㍯�S䣳�7��f.!�������B���t�rtZ�ס̬J�u9�q���S��l�v�e�{�h{�iٶ)^�ɷ�5�>����
��,e}-_Jȳ�[ˆ)N���k�|g&���w�|����K��� v�jT֪,�]�φ��Cv��HS3dr�8�����n�]b�`��������dY�~��<�[~�{���m��:�����asv���8�ތ��5�:�Ԗ�S�{�j����ZH��%4�E��<���&Q�K�D09�ϝj'����;%,���!��UUO�����Ҏn�Z֦��\��� �k�PbRb��o-�������<wQ[���m�?�.�}�擱�R�-�.a.tAʺΚ�ά����	0��k�M+�q���l\�����P#��Ҙ�d��5B�oR\�w�M]�k^��k��sB�	O��L+����3���[AW���Eq��!k�^���qɴ�ۈ/��|:ἅ�rs��;v�Y&
��QC��,3�r��f���E_=�Ӄ��ɪ�j��cs�n��7�����y�_g��=�F�Үf�\��Rs�p+E�ҡ�^�5_&��E:1�k����z{O�4u�g۠C#��y��U���}T�t��#hc�t����-���cK�7�u���YU/[�W�l]�*+���u�3����ʘ����k��^����-�L�'�5ȇbM���������1䪸yp��9�m�A�PR s�we��<�g�X��ٸ[Y��eG�ɻaɹ�
��o���a뇝 ı;�L�Ú�o,"�uu�Zơ�Qje��/����`v�v�w^6�"=�3�u>��US��5��{���8w��
]K�E�E7�;���֚��$E6��X�y9�����ߣ��x�9�i���y��[T_u�#Ͷ��=��:j�7����l�~�vA����o�M|����z��عߊ=/�&�۽�uGq{C�%6{���x�d>�[��V����8���ur�0�o��'�1�U�����[|�l:y#�v�i�v��c�!Õ��,]��T�б	V�ɥ�/�>u��^({�	�څ�ݍiB�l.c�7�����o��asܖZ����������%�mJ��*u<�WtgR�*v5�; �n}����ð:��a��{�p�-�cɸ6�d�S<Н�-�B��ၝD>���'bc��]�c���:2�k�B�����u�Nc;\v�ݎ�N�uGF�]�G;�xGe��﫣q���7�:�T����´h�G�AwsY�����܌G��.�(6XH�m�@��9�_`��wM�{EomI��]�� w4���mvv��]F]^9��ǐf�tT�[�]Yy�r2`�S���c�ս��r���Kn�|�������[�ĦF�nX��Mv�,�n�4E(�e������G�B�] �y+ �d�=�,���>�z�fkt�ޘ��e4*�������殨z������\�:�6`y;���VnR�J���|�/��;��3m^���`Mܛ�0$�7���1(��t��GzQ=��=�.��Uoy�"R��Z'tUw<}x�i��srpc��Ӱ�[��!I���m�}�J�{�����П���I݅D�;������b��#�YY�3_:A}Og&E��P�.���]��6;X�UY�b�j�iC��r�Dq��l�pÍ���MHA[�x,p�̒W��%RY5}c��-샚¬�8; �N ��n
:�sK�R�gn^P|_NO�]ױ\��o��]ΤA�^�FA];z�m`�6�-�λ7uF:�(M�uu��<�&�!�]�N�p�\4�Bve#!���X�θ�x6��:�;6�pO����VV�P*��_U65lf����뎫�Z���P���{�_ҷmF��/$��	�����r��F�� O��uc���|���M���q"��V���|�Ǹ�
g]�A}:�5�d�(x�	�
��x�}g�m]��ɍ�O�K��ڭ�Y��WZKq)�%N�ݐ1hl%��g�.��F�f�Ϙޭ�xM���ʠG0E��/^���>9���!�`E�n!P̩�4��^��I�M�}ח�i�ʂ�u���%K�Yy��N�9R�2 Cp���hٙ��̋
a���v�'���4���:n7�ZȹIj�d�~6�
�]m�w���$d�����R�����Ԋ�K,����\�8�%���dN�Ϫ��t|(TC�fhuɝ��Ӄ�7"ST����ޣ�$���Oq�����%�j���h�&�O*�*e'���v��Y��&���]�VQ�5�P��7��2(k�G&VV�(b�;�w8�v�T*�n��m�e�t8�*�P��5[I�#�O=|��i��	�����^]��I��`�2�76���j$ګy���x��;ug�H�:}-34�|j������H�W�!2�-�G��w݄��3�u�s����*6bۻx���f]Z|���
&	9]�ެ���ʌ�vEB!��K/F-��7)��<P7[���] Mq	���ʙ�Ux{��RW�6�-J'+{)��.�3A��itm�l�����iga�Y�T�T�%�$�\�
��'�ct(3��9i[ֶh�lva��)�g�4�c+n9PnTO�en��aX�[��&������z�v5�qt�^)+���ǳ9[*:�n�w}D�<��鵯���{!�Nr�PjWs�~f����`�Y++*
�iUq�P��\aQb�*������R�P�SJ�*1U�Q�%T��"�b�
`�̶EQb�*��"�ZfJ��Ȳ,TX�V��`� \�-�QE�(���T1 ����c"�i-�� ������QQYUAT��`�EcT���aU�&+�R*����DJ�R(,Q��q��)�T�QX�IY[KAJȰR����
�@ƦZE�EH�*�*�`)E
��B�Q�A*����DQY���c**ȰX�ƤRV�F-��r�iE���*A�����v�/g:�`Z7ƶZ�2�;é8�a飝K�]�ݘ���mՔ6��:�ۡ� ���@�Ў�?}}��3Οh����SI[��=�q���֓�V�O�����r�2�Lڮ���^�Yisۈ	eBTo�2އ�ds=$��v���蚱�1\1qA{�Eѽ�^|�O1��X�������i��O%��lrY�U�*sv�g4�'d�S��x*�H���-�l'����Q:*@�u�N�p���Bk���k_���z+]���
��ch���-PEt˓�M�d&��bN��X|�>�����i_o����i���|I�G�=������sմ,Wgbܝ�z�w�{�����V�Khq�'���i�|o��v�����U}O�F�����P�=ܭ������I�4q����Jz�7�a��EC�K:��w��s�vks���[�gf��#ϭ�d�#_j��xoR�2��X�c��Օ�H�t�g���8�o�m�� �hF��!ЭI_tT��.�[c��ݎ-��l�g���\�H���h��qv��
t�e��b�FIa=��p��]Sw�,
����WCS�����>�V���-J9��1ҙ�5t�o�i�����|����ր{�n3��]r�_��S5}\w#ۙ�f�y�Tǲ�2�?�Y�/J�橩�I�*ZX�R��k+m�M9iM���ݨ�n�u��9H�J�̄�TE�ykGr蚵l#�5Yܕ���k��ı�S�\Ӎ�푻�{O���Y�v�^PJYG%8���;Q�{��	8��,��#��ߌs�/띥�[�����Vu�uC]pϲ�{.�u�Rt6CtcÎ{%��!��~R[��zvF}T4����_d�'�c�.U7��M>��w����*7Fxcx�VZc��.а�주��4�����y�v�o��}G�ʎ�O�y ��K��uj���x��ϫ��֍�ڢ�o�y�vj�Jas��6n�%/����\��7�wT�g#ϥWì]G��.YG��E��M-ۘ���e��s��S�N����x.w*�yY�z�V'�o�b6��"j��6�>"���C��jD|��9X=n����᮳�C������i���̮�.�a�P�����66�֢(��T�E8�!8ID��^�U��]�!�.zx��S��%��u���v%ٕ�R��V'R	�I/�����d��cUq]�Qi��#�hw�����q���i=nۂ�<��aq��F��[�����ǲRv��-!���iK��~qs�#ݛڽ����B��Պ�:�Zد�7��Kv���׳S��^�'�m����{�f�����{��o�ㆃp���^S�Q[���O}����Z�Y��Խ_x�
�2�H7��V?+�-���rj��!(�(:�ѝ��C�ӤU��ٳ�\#���L��:�V$�_$.���g)�Sq�L�,sѳ�)�y���_�Ko7V��5��no��*���ޯ��v>���cy>U�n딕a���.��W�5�&�Ƹ�X����ەp!%mG�w���j'iХJ�#�6�u�s���<Jh��i��nb�v���N�
\}�F<�}t��^�Up2��ٝ�M>������vv�`t�.	��W��{(:�|o>g&K?G�
畾�U��o˼ك��x9�}�3�!�8\%��S�L�b���~�q$����]�Ը�� A�sY&.�~p��zőM�;�\k�{z���\�Z���Q�cȝ����{xk���¾�I=�v�5�:�ĝn����X��k�'�^S���W�3�e������,��+g�A}�y�s|��r�L��܉��;�l���ȝC;���r�M��*\)�}v�]W���g��[�X���Ե�~�J�+�̄�`�W)�V.��Evs��nd�6���sZX�/'+���(����L��Sڙ���mUƌ٧�?Q���X�ު	-���V-�Լ_S�-�_ys�D��)뭑��7��^E���w>Շ+lfQV��\�s���U�3��-��u�ܠ��:76����豧��Iе��qm6�'��7���� ���&n��� RoS��oy-�z�5��s�������	���έ~�|9zj������yi����.�w�9u���O��;*�z��pttkݾz�h�T��ܦ�����n�Qu����\cs+��H���.�a5�gVʟna�� 0&f
�S2��[�|n�ۛG`ԗO<q78���巂��͙u���<�lBο��rÝ�W�G��+.njwf�T���vc�N�Yz%�E<E\�
��u}Y�x$�+��]i�@չ�Z�,�]�m�f�]îw��b�f�ֆ���47dB^:��\�_дt�$�Bi'��8��*c�����j��af��C��t�؀u�P��ñ�؟.{�<�yZ;^�+��Qǟ�R�G8q�C�tk�Sԇg��r����
ɾ��,��c_H�.rNpI�TG��H�bt�#��p���wb�랸��L�\��t�j��܎����_[��[�Oe����v�K�r竹�A8���f�v@V���̧�CX]���l�U��YaQX����*,��^gZӱ���S���d-mAچ����Ν�LXחW³>rd�]�G����j5�3��+���� n�c�v2��������z�h�-�-��h.4�m��5� u�r�X�o*��f�����>Q����s/7�Zڨm-}�tq^��g�}�b�F�B%MAP�yܝ;��f
��� ��7���oc�7�_�A�(��S�?9G��kE�]<e�r�Rtl�r`w�ު}�n�q�L!���%C�K�
��ɥ���g&�r�</�J�A�ú^ۥ�r�3�h���pТ�vg�/Dٍ����D$��l*�L�����j!�/睸�'ղ�ս�Ҿ�j�{zƍ�J\F7s�,+��%�;:�n96*'��Kv�ŷ�����V�;����qk�.Q=C��1K��o�+��T�5}�}��z�u���<J��8'���=���=C�r�Mf�\oHp���[�lne9�'a���=�\�es��f�o�콵
cc^}*D�¾�k.1GM'��[ҵ^4 U_]�E���
s��ʝN���А��
���ˑޙ9*&?o=y��s�ѳO�M)2�!�Ϻ��Վ/i�1P�*�%����n�A��[�免�Wѽt󛧉M��֎�Lb�C"��˴�{c�5}�C��ۘ��W<��2�,�M���ք�l��8�5���bL�X��Z���8����c��+:,ߗy�W;�Y�;C�4�vܾĮ.D����A	kPo������"&P䗒7����;gf_J	�X���n/stt�jx��QR��y}aP+�3R1og0Ͱ�/4Wu	Z{0:}�N�)*R_Nx9�ۜr�t��noU�����}����*K��-;�c�?;Eek[�l\o�`�����UxV| �Ok4�$_��������귦~ŎisԕK��ʷ-��7�f�T�����%.m�PV��Qy����$L�f��
y~�hZ֘޷��&B���Ɉn�X�Q���Z�8c�'ԧ�T��{��*��/t���jy��s��E�u�ޚ�n�>����ǁ�g$�z�'_�S��9�-�n(ݏ�{^J;��z�K�z�!�mv�i�N+���3V�:�QnE+r𾡑γ!sb�����G������l�F8�N�H7Y��yT���o��e�wy�l��	�s5�:�K�H^���Z�s]����Wq*.u���-���Ү��.%�nF]���������c�[kl	o�Np����ã�#���w���_$]K�����7w�%.Z�.��n�Y�i���R�-����7���L�S6śPel�t,EB����0�f��d��g)V�ou����j����WT�
�5��c�9����[�J���,������{ꐿ�k��w�b����D�.����7�	��d�LZ����r�k��^�س+d�;r��U}#f=�c{���bow;���rikakcs�\d�ހ������iEf�[ �ӻ29����O��u|�pW�8ŐE��"l���Z��q�BdC�Ӵ#�(�9�V���2�rv���Ywv)2�@Ӕ5��� ��-�xn�xQ]��SV��b{��e���a�;��uu���Y�ܩ�j��\st+b^�E�y�q��{1q{#�o|�ﻅiW3�د�q���O��*]@T��;��K���E���)�]�����&����E���9��u�Hy�d���9�u�fl� J��~;��v�!p�s�W}>qr�T	�3e�s�t1���a��Cn�gL���C�Z�ʂ�:����r�c��Q1�I�OT�1c��Y
t�Vލj�p�(�����Cih��?g8�O���]����՗��<��/+ғ��n�qX�,1=j���S���Ț�S2�����>�|��M짛�e�%ˉ����|�-�GmQtN�%j+�V�񺲧�L������V$N�����̝��>��/��r�Ţt���.��/5�������N<��Ǥ�D���!ۅ6��7����\7��vm���A��fj �T�m�y�-��벱ؐ�>-�gV׃��uk����}���N��xZ�m>�v��*��V��-Ն��o�Y.k�)�4(�f��B�.����k.weBkk����ֽt/iJ��������h(S/�6& loT�;�R�h���ic��5&i���d]*��=�[�����zr�w`t�؏{Tk��cë4��s�����C(l��=������q�n�����wD�@���Ah�ځT����։���yì��8�b&��	��â�s�o�{�b������5-���L��ڳoq3p^B��U3¢
X�����g96�ev'�
��t�K�Ƿ�����3Tڇ�\8RsQ�C)�,XVx���&�j�t|�ʆ��ެ��C�� G4�^Ƽ�o8�4�
�5oҎWjv=r�-���F��=�w�z<��Zgzj<�]����:� ]�,w7�sw�F��+fTc�Aŵ���r���<E���`N�^@���GJA�p�d��3a��oP�c^��8�6�+g"C,m�+v��u^c���q`3�n'p��-m��E�<���y4��{ֶ�?xz�ô<օ=�.�+�i���]RcjdT����F=81N����-�bVYc��j�j���m��1VD[�W���b�Ud�{t��'��noY5�q�����S'E0�9�v�������vN^�y�������S��f��#���ğ�&�^�3|ս���m�E��0i���p'ݷ=^���,�]S����Sb�9�{���4�����4�x��zf2B��z�c�퍩�5�՜N�+��T��-e�i�����͹.�U"���z�窜�5P�9���X��&��)�kKy�)nt\����ne��m.���|�k���4-�
f�u*%.s܊ꛘ�{]���j�=V�����\`ro�����.r� v�u;���q=�_���Gq�AE��9�:Bλ�ɵ>4�������@�cJ^�٬��3��ީ�Θ��Gz�zVG����X��&�d�.�Y�]������ʁd�z��kM�6z+D��K�;�wn��B�q�Ba�Y�wu�r��{.�����-m9�fP����AR���\�"����\-�c�k �R��"�9^��ز�̳�V��h���%��0����Mq�.=ݩX&���dR���/J��'d�����۬P���YC����ɗ��[Ä�I@�.�r�y\lE]BM}i*̗[!�Vgr�Y�� +�qB�&�`�A�����-�֏df�)<尝�O(�r���U2��+��ȣv�0h�m�5��+mb���s���cU��es�y[���h�i.XM�Q�C�P�d��󩓁�^�ڭN�c�e��(q�VƘj�0shvQ�VN���ot���u����[���6�;ωut^����p豣�;�F�n�Of��(F5�5�;�!��ލ�Mn�DZ�5��
\�G�l�E�Y�^:��P(�i��
3&�0%�+9�����q��6�Ԭ���j���9�zm�;��c��LK�T+��b�l/�b����Q�r��gm�VM:7{�{>Z(:x���{ǲ����`��n�I��Ê���"vJT�ŲL�oy��g��m'��뫕BT,e	�롩�
�ʳx���V|(����d��J���U�մ����Xz��i�71\J��'�6N�e�\�8�UՄ���c�1�j���@��;�d�,>o�OV��>�튀�	�,�O*����qΉ\�J�P��ɕj�La��P�WZ��:�+�1�g)-;�����ÊƸ�@1�QC[O.>+y3��7v�,e�Zo���w�رEcm (��q�?c��kGf�Q���%k"j���=g�
�V-#S�5�w䠼q�N�k%�2W9Z'.[�ݖ�d�mg�T�U�Hj���W'���|k��{��i�u�	�)Z��x�캻ǭ������ܤ�5#��1�vd��ʁ�׍����N�"Ѻ5+:LH�N���:n��s��/5Q�u&����m�9��a���:�0��ݖ@ ����'ͥ��S�鼑F,4��]m <�u����nϳ�,��X������V�8�el�w��z��ʛv�q��م�����IS�&Qϧ^$&�{2�[��G7gBJt����Db��[7u;�����Ri�2�������g7���:U!Yz.]]ε�DعojfM���ٛtL}G�0ZZ��H���efց#��SuW���5 P�V���M,pv�DȫLx���A�(d�9v�rE��S�(����ƷF��.��\�
�<o���m�S��N��yy[�2�q���b�qϚ\z���muZ��-�b�ЮC!8�R�PK0���)���ݓf�i�NP���љ�J���h�H'��	�d���5%H�SiD��"�HW󌈚j���RŊ:����*�dY(�UATU1*�q	V1H��IQ�TQb$AB��d��]8��D`*(�"1A�L@���(���`"����-�QDt����1X�e� ���b�ڤX,D�̺q&������U
���b%J�,QZʥ���V�Y!��:J���Zə@�1���,J�L�Ch(a���Lh����cR�`"i+��uL�����L\��FШ���"��PFLj*�ZkTj�"֡��M:a#ē�ID73�s;�ᵺz��5��u�B���9̾�ͺ����&�++�ӂa�HLr\��+7&(�'�� ����m��;V`���+�sߡpsI%6_sq�(�1N�L�]�0�\^Zp�2{:�Y׈-b�]�O.󓧉M��֎��*�v&�������uu��^E[^T�r�z/3cӅCκ/n����C��S�o���[�#�R�sZ�.�L�z��PWe|i�E�evMF'�YP���¶�Q2V؛�Ê���e��
��%&8UE�7��R���K��zy��@m�{��meJB��khi��1�ިk˅�gπ���[��Υ�9~�iEģ��^�p�k'��ei�p�mݽD8�z2[�Q�+>��ˈ-eA�n�nMv������5Ӭv�Ƚx�
�p�{�gi�c#�覟����PxB��������5P�6���Q��)F�w&*�T6���մvÙ��xs"�;�b�[�Un���N�hC���i[7»s�����/y�jWK�~ݛ�n}�a���'&/�I\��ھ��PK���C)V�x�5��r�r1�5���@�T-w}�I�V'��X���f��7�4�!Sn�[߯o{�4��](�ł�{���#��s��k�WB���Ӿ(e�۝Z�m��m�V8!-���1~~Bi7&�{Y��3{H]��Y5q�B��O*\����v8��[���N�oFA�+��J�:ՎJ�P����M�:�Z���Kyx���v���)���u	�?nu<P]�>TK)�3��em��w����[��l��9��:�GCUu9���}�ggs+X���E[��I���Z�ү�y4���W�2����8�KW����ɮ�p!l�nc��#�]�\��&���q�wC/4$k�����O^+=��Bo�����+��9�W���fG'�	��)���!��sV%�|����:��o!U�
�� �6-��%nM���I���,ĺL��FT?Vk[^o�=�n�W��Λ�Me[Qx;0�:���������--sK��Tr�3U	�}eK�
���vY]�;6#˪n3,���"���y��O1�y�ȼ��c!��p��ʻ�]�.�&5�{1B���v������{z�/n"�'47y�h�O7���-=�R� ����*�ɻ��M=��<<�ۋt�3��}�����M"��x�WE6/��`3��T�Ԟ_6��CR闃)@�e�醱w�/"x�k�9-����r�0f�D��7����4;~�4�W�!i�0�n혞�;m\�9r���.'ϥ�i^}N����eԡ[�SDS����\Y���+�񯖋���S
vb�E<���u,Hy�1���w	��w�R^��k�f��C�p��؞Ts�5��R�$^_���M��w�y<^Bn~v���^�9v��T\w�]Z\���iP�;2�,�-�es��������ʷ�[��gq�Wxg�n��Ҧ/cY\�l*ݟF#3\�,���_oK{��۷	�o�U��P�FJ%�[��&��ϰ8�lc� ��3�����=�m$�`\���0�rg�2:�tS}-�;Kg�nǍ���k�zx��rZ��!�����|a�k%�(��t���^g9������٩���d��W����_������cWz�D����O��V��ߗ#��`ִ��X��Y�k4NM=�����9�M[yݒn�;{�+�]b�wu"��H�r�:���^`�\������5��%�5�n�J�eO1�c�=9u�噫[JyU���)	�w9,Ώs݉	�t�:�vӣQѦ�vц�+�OV@������=��bVu�8��w>�w<�]�Z���Pr�;|%�^��<}�m3����|4���Po<�{��U#�G�a�-��������qu	튷Gn2��`��1������P����}{��Oe�R�	~�G"��:7(��k��:!�:�eϖ�j�}V�;
�	�e���'�-����;Y�7�e��gϨ��;UvTWmlUͺ̫���I3Y��I՞[�9Gf�Z��^mw+[R��~AqZ���3byu_%��>��Ju=�w��}w�5����{P�Vg�l�\C��x���c��Ugd�T���l'���-ڈo1�;�JF����tM��-I���y+vK�jʾ�����;u�U�j�J���V�EU���X�f3:�*��*>�! �9x����6�ʅk�tD��\B��0�@��@�{�tŭR[�!5�}�*�F�w��\���o6ˬ�빳��oJ�����lx�gx��muͶ�������Ʀ��_f�#���J*��t{Y���8���|w)y��jKy��	F��>�rWer�r����V�U���!�:�,tk�{�oQ�[����#OA��/�ɤ��C��u<s��?2�=��^��z�Hˈ�ۀ��64�"���-��,j�]yT������.��\'��n;�4�Rv�_��ה��Tx 78iE<�3O��M\��U���ru�-r�o8'	tQv"Rr�܊�UΚ}=1Ɏ��A�N�#�� r�f�y�W��t]iu۽X����2�kΣ*:x�tS�[�Q��v|(�s<��T:�b�K{W��8��`ް��t <%i�Z�+r�)ᘵ�w+�FKHwc3��T�X�*qʌ�6|ڇ�T�
�^���e�����W��D���m�,�]3��Z5�mo�Zk(��f��w0oN�/�G�E�
]�КG�Pt�W���3:4�e��M���w��%M�B�W�Y���t�����I��v�h��v�v�ߓ�O��<�';�[��-�p��hw �d���.w�;��+�<�u�R3{�=In�	�3���U:���OFM���V]}�Y�O�_T�3��]�;z��xo"3���Q�-��ή�g�g��]v^���B��'eOUn�n��a]��\��{4��������m�2�l�yt���?J/ۄ�7yt=oG�퓢f��8���.�������XU��w��a��;�d��)o��7�1/�s>��[��^�k΁ry���WV�q7u����q�-��>܇�9�e����B_K#�b��}=^^�=׭5$U/!k���5��Q��aN�����7�s?u	�?+"�-���[��x��Q��&����>�^�|Z���f6����r�]�Q��І<|Yݩz������2 zg���m���{����̟�QN�a��W����9Y`!��p�,ղ} �@݁�f��uB�`un��S�Aʲ��1�����Uҭ*��Й��}���]e_z�.�Gs��iL�W�V�+�_�=�䊨�&����u��]I�.�%��`�9W����-�ٛ�E���#Bj�O]\ݱ�;'wqdc;I��6D�{B�*������[��:��F��CR�ܳ.x.Qn�	�*{�ٱ9���V��	us��A5hl8�`��\�����5���݉�\�{r�s����.װ+�y����i��cL��raTv�`M&8Qۘ�=�Z�c{�y	�,��8ؔ��nv�,�Z�v����pv�� J�;�`5�gB�Kx���ڱ�']]�Z�8���*u�Bo���yOe�6�C��[��w)2ـeQ�
��]��w"�3��e���zc�W{�ކ�\n��֝Y��wq.�o��~<���b�\�J�<�Qnu2��9R;^�n�#����N�9��q�Œ� ����q���7�紗�e��M�{$�L�<.�A�Uyγ��^���vͯ9n��U�b�o�7ٙ��8f�K�$�����6�U�ʬ�M����{��&���R.]]���xZ3 �6��z��G�]u���\��J�P`h���'_<�Mu�rHy�.��,Pw-�E%�N�Op�ݫ=�p����N*y�����nw^Ҥ�gh�KBԻ�:�����9\ۭ�=n������-��E�0�fp�"��4sL�[F����9_!� D���%�gP�ޞ�=觗T�0�Z�>q-�t��=3ֳM�@�[P�ӻxv�!ҟT���_�ȩ�|M�L���ǯ���>>���AL9���g[{c����g���n~���g�}q��U���q5�J���J�}���E�u�gn��mw���'�D���/!^	ly_����pVT��r�4�b�4+�H\ah�y�^���@{�=��F�E�늿���9����o�tW�����-�` ���gQԟC&���6��w�+��yO�_�n��'�k� �s�G#����n�[�r���-�O�с�%���eu��Ǣ}�&i��ч��;�����5�Uzae/L����
��ˇrvs����pV�ٽ�X}�Q>�����.���11Ӓk�S����������C�r=�z��[���Wz����@g�vA�� |qM�>����=='�J��ǅ�vk�_���g�e3�~��O
&�x�9Z��ǋ�H��\�=��y@U܇^���iz�F/��s�W;�W52�fgfNx��
	�iWU���W��]��W���S�v� ���T;~��R��m4�M�5�x�J)�e0�d��=ˇ��a�:�Bt��X��L5� ������cgm���{�A@n��8���cXZ�]��|�er�Z�Ŭ��3x��J1_Ho�ǒ�lg��t�;��~���_�
�}�(��2��q;,e���v<=�_�M�>��>����t��<��wS�,wL�gO����8����+���m�(66\��|#��#��yzxW�o�֗y,P��r3�j�_˞xl�:=���ى�=�<b�x��1�Qz�����g�&�tς�ɭ>3�7���}鑽�u�-�q���p�#}ܭc���PȞ�3�Ϣ�����ق{�ğa=3����'Y򭻄�K��?S�Δ�驝1f�«Q��q�[�:���8l{6���ӱ%�鹨@Mw�*,�*���f��C2���tG�=�SIw�}/���o��c����d�,�9f }7PI_���jI���ǳ|�ۇ=ʠx�}�����x�wO�}:*=���g�eK/"�Pz@]�e��/}�Y)�w�z��7���܈}D*�ֲ^��3���v<F�[�^�t|��[�Ie�'sǗd{4ߦ&���5�>fʞ�̍Tǯ�트�W#�eqR�H���i�ʿz7�r�fe��������Ⱦd`�Q�����|Ȗ){��AVv�;:�4]�(P���wK���!�����N���0b��n���8�t�;۝�t]2����W�N%#�s�����H��k/h�%R*��K�����$^U٧G2vlR>�2��Z��u�qK��;C���&��LO�O��p����(z�N����(��qf*T�¨{4��Y����Zj��S�}2���f�	��}[GC���
��|u��9q7��y��k�\E�P��:���@{���{�(��?QD�L�-���c�3jE��Nϫ������S��u��5G�eqj�Ǣ���{�#�s۸�Dx�i6�
�cx�M��{tԹ���y_�V�0W�?|�xTicL�|�|='���^�.b��'MG��pй�;��/L֏߷j*���y5R3��F����D� �2{K����}>�/i�ܯ����#�Mc�U�lZ�=����|Q�BBwM��;q;Qv}��Mi�� o���i�������#����ˣ�{�qN���#7n�P��5�Na�?���aY��ڌ�L���_:�׃��S��q��{¼�sȟB�Lwk����Hh����	��C�|�Ϊ�J�V�~J�섢|���lQJ��W|���d{޷�#�>�]�ˍԫo��QW��X�rW�ߪ��֔���� ��e-b�������7����k@��[�ݐ���Q�g��	&�ʵj-���?��.n����73Tma�I�Uk�y��Gs:�g>���/0S�.T1���Eʰ5��/���d㽕'�=L� ������d�(����p֞�F9]d=�Έ�P�"�����1؛@ro�����x��R�7��ᯯ���V�F���O����A=��}y�93]j�bs���keAq��܁�r�����Sĳq�t.�u��cqm����!���&�,����-�ho ���,�k*[wc���Խ���uj��K ��S�S�H����^A%���.t�%Y�PY�����K����'�gkV;��@ ;�J���#�vf�Z���z*Y�UaT5kUE�����NV�[O�����b21�}�k�o탇�UvL��[��(t��UϠ�M�$�]GJ��4�%�E��km���X�e��hE���SiD��ܷ;���΄�����K+!��%�wVT]�2����*�}�yE��z��V� Ok6�7�Z*:���.��Y���3�lne� �+V�����6��S$�3U��]#�+��7�N�vkP�A���-�T����Xo]	;�h�U-r�ThMY���I],s��w��,���6���Τnh, 6��C�^W`��o�$�I�]�� NN�إ׺�R� ��Sܳ��PX��lp[@[��BP@�킷/�ʡ��m���e�*5'][�p��εw^ ��������u�q�}��ڔ��! �+,��(;r<凄S���(�L��~[���V�׉�M��x�R�|NF����x�tP+OV�3��m�']6��0؏���{�扒�oc�W�����y�d�q� tC
� @��o;i���*��J4��Mh)]Z=��yu�
y��3��_�sT�˝�<���,��etN�,�N�1���v�f^c��v��N�*��nk�m!��^{	�Z��P�j�%�Y���bI �C�ލ��tM�P8/c�Үَ�ړ0��N-Z4cŧt���U��梪n�$�k���.ʾ=d��L�UΣ9k�v6�ş
��XK�f�U����5��#ظѻQj-ՋՊ�1ҝB��x+��#�	��Ȳ"&���=�]�%��G/
��FXƔ�]�F��B���g�ǉ%�av�=�|z�a�P�QK�]�w3���ȶg>��wJ��9j�&4����I�u�%)��.@[�o����]�4^���z&�Oa�]M�9�}M��o/����q�`��O~�y�Q#\�+�HVb�ҹ9�-�V�g��燅� `;֫0�6�E�aUw���_[���R�w��##��Kl6�Y ��B��?ȼ�{�R~:��E�Z�Z�|��6Tۭ��Y��>�S�v���3��$��r���������X*��qȄ'�"B$�,=�t�,lәU�E��5�(�`��kB���S���H,X�a�r�"�Q�őS(��X�(�̹l�լ��ȡ�f0��B�b:B��
��fB��j��EĨSVb�B��U�*�,�1EATQf��k%�Y�r�B�Y��X�`b�DeD�P�Z�*9�kCl��֊��h��!�DAV)��,X����X
)X��%E�t�&9�Ĺ�)�[Tժ1��)r�1*6R�R��Ŋ(�%m��ŕ�-)b*�XU���T��IZ�DY�Q"*��
���Q�P�*TY�ql��`�R�(��VZc�B֪6����*Z��,jZn���Q;���p��sw{�jPo�}m"-v��+Bũ�󝏜�v��`jA�
B�U���3��S�l�����I/{�N���
�#?��e9���,���Ǵz]���x�w��o縮.Ig���ȱ̩�׆g����wR��[視	��{���������h{!�1y�U�}���U���Z��|31���Sf,�`>�X�ߧy��#���#�l�n0�,��GT,^�,c�/}̚����}[�ܜ�=J3�_���8d�n-�!�*Lq^����G7���_���
��L�3��J�{�W}���`�F���Q~�"�z��,5=s /�1O��v	h���mU�^t�r�A������K޸��jߎ��
��z��{,�_C�<ML��n&
���D\��3�}�i�H�ݘ��y��e��rϴ����u�����c�K�w��I�s���p��oMدV��+��`y����#��鑯gá)c[�"�������?8�C�䤪��鰣F�0�>KS���}%�뉺������9�t�C�n�x_��z��=�Bzn��p�ٛ�D{j���3�7�QQ@J ���=����N�����c6�>����_��Z}��)�!�@�k̩��l��Yf-x�tw��1h���VE�}FB����^ק?r����Y��+	�(�=�*)��|9ڵ; ܨ䕻�Ӕ�a�.0������2�k[	���X�5�N�Q(.x2�ų�;�F*B&��oj	��|�E����F~��iY�_��s�Y���c�����R{�oK��OA����7�v{�xR���h�:d��E��:}��CW�V���t���:Ǟ�V�\�G��v�kO��?V�9��d��7�|������7��{��z�q���Ҝ���i�u��^V��I�(��\\yfC�o�x��5���ɝ���!9_uz�jg��_�����gQ�{���ܣ^��q]�ื���7�K����z�	���&u�r+n�g�PkL���q��qS�П���ڻ�eo	��]{��al��|T̰2*y�S-�HS��S7/�®+KC�AF\�h�W?b̏.=�z�8�CÊ��!���w��bb��M��x�����zT�ݝ9=���{�H9h�}�v�������3ⲥ� 7=�<su�E�@�b|vf.�Y��}_��8iy%�>7�Tm��$o�O�q�v�tU��z2=2���sq0X|0�)ػ�Y~�u*�� �A��s =�3U?��qW��}9ģ��H����Y��D����͜+�?��Up�z�Ax�ݻ��\�&v�9�������w�;�GϨ�Q஺���W�O�]��%�}͂o�}E!jʘ÷�u)��:!B'˚���9*wCy\�u�l�ӫE7Ɛ���i�O������ۍ�» ��JV�Z���e���mj���&���3^�gFJӸ�7	?_�>�S0��zd�N ߟL�0Ԏ��k��z��� }�fפ�7%����G�'���U�o\�wg�Sp�\����h�]-�bB��^Q��Ճs6��߇d�6�vA߅ I�8ja��a�~���K�긆�Çy9v=�]��Np���[CO��ͻ�G�@Jn�xw��,��IG.e���ͅ�y�P�g�t���_a��Lf�m��Kv=ZL��j>~̿�Q�+�ƾ�{.��Q�}�(��2��q;,dV��W��ʶ�{����|��X�5U��6et�q`J��G�z�����n=�Wq�Tp�#�wN�I��m���}��kR���֌�ɭ>���:��Ov��;�+�Z���Wq��_Jx��y����~��z}m�0ǖ	�$z�]UᕓZX����t���c�9���u�}��X�i�������mv���F/0JF�'�a��+�/&u�gja1���{��ۘ�&������&����\w����u����2�a�Ia)����1]�y)��z�+��:2(j��x�=٫�Nܦk/�fY�)�^�]�&ظ׀���bHd�L&���Ԕ~nH��Λ����2�϶�`��W�t����ΑaT�m������|t���c�"��-����=19M�;J�Œ����!�ܴ�����hE���E�V���r�^�G�����)�����vD_����u�ج�TY� J�3�w��$g?o�,ر0|�U�S�S�����[>�4
)����6s}!��o��U��0��e�epg�ű��>�np�ߞ`߉��Mԙ�N�Td�y��}D*�j�M�	��1���tf_��?'~G>u�!H����su�E/�\D�ǽV���V.W�?�|G�Zq.��{%<�xJ�~�0:u��Ω�Y#Wu�辦n�z�&��LO����"	kga<���â�{4�[�OM���w$p�v���Y���=�B� �~��D>[B ���(X�������a����P��s��Fi�~��gǢ�@{�����E[�M��-�3a���!rw�<��ԜC��O{$�|}Fڗ�۳Q�z��{΀�9/.���I;s��I�Zu�<�j���Y}���>Ѿ��Bþ3Ѳ��4�X�י���T}1q�:��{�w�g*p�}�9+^�H��Ω}�t�~�+��>���������Zn5��f�m�Q�����:�K�8�����,g�T�/2�3{��t�2��30����h�/w��:(��bFɫS�4؛iZA+þ���ߦ=W^^�k�C�'-���4���>,��o3v��Ċ�O-k|,�ލپ���l������1���X�Y�)T��eC\��d��W^o�^��̆(�?^F`���ǵ�V��֘����o�;m�_.���#��v�^�b�n:��W{���v����r�4^�Mh�X't���uT<5[P�3��nu���l�V9T7��L�p��G�F/���n=���y�Q綇�����̒��L���B�Wp�$7DVݑv��W�Vҹ�J��|s�Uq	���>�T�Zｗ����_r����X`�"���U3��=��~2�>`y��XOz|�㊽V=�����{�����qsJ�5��eA�|a�f{�j�6z9�>�����&���7��f��H��?c�J�3�Њ£=�h���ѣ/�7��rʞqU��aZ������F�l�o�¼^�C�!S�_
�t�X�����O�zb��N��j<��g�������T`/J���}���~��z����B��+צ��T���i� 1��g���3@�9w 6j-M
���a~���]��df�Uߏ�7���Y�P���y����Z���{Հ��e�_<�t���,.7��c�Y/Ԧ��g��?��U�=x���!f��yt%Ē��nS�ca�:��-*�5��tɽf�\��՜�P�`��ۍ{({/n����>�z�{�o"�,����gM�zsn�u9�,�WS��3�6��:ܬ��ĵ�Io;��Z�,���PU
ו�pN��S+�y�wA����Oƣ�ʫ�A�V��'� 5TI�s�Q~"Y�#�9q�铛�͜�r�q�Sc}�D:�Zdk;㼌�7�vj6ӯM�_�·����^��w���c��dҬ�{ǥI�{J'p�$�51�[���>&�\�3P���c�'�;���>�3~���j&ub�Q��j}��ׁ���h7���z~ǵߖ4+ғ����X�.�'؝\e&G�I��r���/����]����_zO�����d�+�f ���o=u�}�<�ȹy�=�v}��ڭ߉��x�+��G�:�_���N���3��vX�u>��8r�\�Y�6�qh��ў�t�ޟ���>z�~&����{��y⸫�m�Y$n��n	�9��\�{ܲ�=3�}�Mi��d��b�]�:�V7��{���7K��n㮖`��+Ʈ��Nyw�]�l���%���7=����T_�>ڔ�;��L��F{μ�/�]�56�W��WV�\^�GU���w���F��5|�����G��6r��C�C��>a�̜�T�?<�/v^�Mȸ�[Ʋ%�+e�V(�4c<�Z�U� �8��Rj�J��Q���G,��
�����T� �S���	�<�6s��ۍ������t;QUkw$֭������ds�j\��ɭ�G�Q`�r��t�1�i�i-�䞊G*�gY�K}c�{�>=����t�Wq���h��q5LSt������`@
*�1�(�|�O�t���x�Tg�|;�7����xQRYN ܁�7;^�1����y�rmy))�>�<��!��F��q%��+ސ�3�����n�_��^�� ��v֣���E��FUWz�1��YT* �^9����~/�o��ȉ�&�W���H����Y�u���]�;��>��4�:3�E��x��=�dS=�x�8��6�����W錃��Ku��ed������r���='���#�u�2�LM5[GY���X�ڼ���!�i��̭����w9�	�A�� ���������}FV�y��5^�V-Q��*f=�͍��X�y��L\?Un=�@yg�^]���G�%ؙc��3ax�n�9��F�H�����Uy�����|�}���/��/�ws��w	~˸���p�zJ8K��2�������n;H�w�����ٽ)��y�����c�s(��i��g\UǞ�Ҿ���o�"��}1]շî�v�H��}�2��6S�5�W��i��Yt�MÙ���+vA����=��q��}�T�O|��}lZ�W\ڽٟCvc�{��{�l�}�7��k�tI0�� �+U��LBU�Λh�s����[\���)�fJ݁_;2e�LO�ѝ���"
m+��[�4��9N�&�M����x�;��Ӌ0���'���~��f��g��V��9���I灼�E�k޿"r��*�U(�z쭇Y���ў���1,�n$�>YT�a�,nL��:[^��}^�"f<������ozg�m%HZ}�=���綇dw������,��~5��ɝg��V��s�#=Ҩ����r�(�Y��r���'^g��y|�و1��(,El`���P7�ߨ?����䏇�{;H��~>�9�J�;�#��q�����wų�����ͪ`+�g[�%Q��/�`�����d�D�=������fRћ]��>١��~W��l���Q�h�i=�c��,��υU�����]Y��s����w���T�q,y�}$%m_	��m�ϻЫ���H�G*� n�'ي]m��~���qpKV�~G�4x[�	\���y��S��bT��(as�x�-�����'ޭ���E�"���$j�n�C,�(�)�����11O��s�Z;��Tǌǉ>#n�F7쪵���:=�_�A�R{Հ5�̂)�zm�-�K�>������O�7��Dɛ8�2S�z�������[��	V�'u+���mv^KBF6��y�=�B��V��pm+�eVR��+��u��WJX�&|�M
�gS�;)�3�rÓjHޗg�{0X�%u�gr���І]�+�e���UM�����)���@{�� ��`�+�~����|����)�B|�X�u=dn�>�(e�C���RkOiTn��۳Q�z��{΀�9��=�Q&��|K�RF����d��4��Y���G�rü���'Q���3+��n��^˹sD���w�pI�un�\ׄϧO��H�9[;q;^��vN�Ӭ�k)��9_�<3ι�/`~���F�:#��~�ݶ�r���:�0k�3X�����z�'��~˷���`^��"��W��Q���/�����}�ò=����|kB�w�x|�*���ه~��q�36��>��5��.X�N�G\{}~&���v��
��mw���Qۏ�X��qEo��9b}s�ѱ�� ��g�8|*#��������#�>�]���7������u�����5b�l�`7�]�y���=a�P��=q�+��>�~8���VD>���x�����K�q
�\j�S����W⻆n����)|jz@�qU�(����%�ڙ�^�����:27Ы��P�����vE*���[�%,+-��a��g�J+�V$n]���(����6�={S��H���1uMw�B�D��7K�*̻��! #=�]=���o/!��l3�/�@��3g;h�hC�%c]����x(��]�J���B���v��T6�P��o� ��X��UZ�����q.�A���z��D��;���Q�؄�5�׽$���%��{�Oy�C��q���~���=�n=����U*1_�Xp�����Xؤ��n�D�,���i��_�#�{�H��0W�Ԁ��B�G��-��tI��T5CF�5��s�֞O��t�3ݢc�4��Ė��J��i�Ӏ��D;�u�v&X|]X�f���k�[;������]/N����t�zm?��~W~8}8Ϥ�r�{,�Km��1�ڙ؟KN��/�OA��;st�\F:#����"�\�`]LsTj3�϶�.9��)I~cچ���NKz^׬o���oJ%a!�]7P���[��d�t��\�2���sR|Һ�"�{����ow�/=�(���'Bzo�=��(�+�	XnK�;P���a�O����3¹�e��h��f��uN���S� {�c��O�K�Ы�ۘ,d<���'N��ǵ�
�6��~�Q�������?÷�]�^�>g�zn>ο )m��9���̣��pt����x'Y'N���1gzܿ�~����c�����=Pv��u�׸u�����)�
���O�o%N�Z�}7b=�ٕj��m�9�%]��MZ8{x�Dh��}�0�D=�$�L\:Wn���vP�HͳD�̘��G�{�t綉��Z"��$0F��<��ƭ��c��ӝ!x{]�HY�.ޢBDt��[bE��!c�kzΫG ��C��7Ul�^�S�%Q�A�f]�ڬ�\�b�h�/2BI]x���e�5�<��iٱԞ��:���WwW��XƧ���u9-m1;@��y��zӓT��:�l/��poU�܄��`#����A�ޣ�1a�`ҁnfU�롭F��Z,��Y�%�ikbC-v�
�N����Y��T�5�����~H�_��v��i��-��x��o:�<��u�`�ET��Ȋ����@\TE��_\rd�.ȁ�[��85S�z�9�*�|��c�6�
dc��{jњ�G����m��X�L�6IԌ�}W]V�i�=��諕�K�:nn`���R��@hVI�_�*�g>%|��2�N*�]]��<���]��%�#�S�+:����U��"iPʒX��koA��>�ZX���:����U$(ݎ���wd�6�/1�f�1S%51�3#��_k������X�<����9b�W�n����e�Zඌ	^M��qeB]ְr��rK�"�c�bW2�E���+wF��cA�cڸ�mE[���uIA9���u�`ZhLv�8�y
���u�N�Z�J��o���z4M��OuUݛA�N�@>#D@h�-��sx�on�/���7���f���s�����#���i]o	N���U�	��
���7���G�dvS�'8�5z����}��-��[I��,�ňd�.����6��ƭ=mfڸ��� תї�]�լ�}sh�9�GnV�[Nk[�ڕ{73��bݷm,j;%P�V5���ܕǸp���2�#��\˻Y���풯.�'�"�W�Q�Т�q�u�XDQ�7O.D_7�M�-�ܳ$-gJw�l W8I����Q�ʡbԸ�l�XiPF�4rVI{���.�n���V�!ۊ����9xhfc�zGR�IU�뜆���G2>s�^�Ba5�³�6Yr��S�N8*PYF�
�֨���V�g7V7&N�[,)CwLƟwj���<za9�V�v����z쀪�uv)�)�25M�ͥ�
"�e�Y��
�s%_j��!eRV[Օ-!�]��Zu��Dt�pp��ï/vl4��hmݦx���b��t�8j`h�.��Bh��=����ܝg�Rm6�*^U���J����mr"��B�@;���o$��sy�Qp�l�{vI9�	dɆ����Z��X��m_a��>���ku����ޝ���^oO���l�Z*բ��()U""ʨ��%�YZխ[R���Z*q*\̪l-h�*",��)b��E��Z+�Z5&c�0�Uj6X�b".f��*+�`��V"�Ĺ�".VQ�"
��D���cr�*�DTj���r�Q�2C�%U�D����q̅���aQ\��*��h�r���r�6������eZ��D��Ym�8�\i*-\��&%b��ARڋ��D��j�#*��F�iTK�EeE(�h�+"6�A�)�m�ѴiX��*Ԭ`�+*1X��T�eE���լ��Q�c�cX������E2�bE�ʢ#2Ҷ��aX�n`UEVcAFҫmQ�Q`ڱA�E̡�,H�˖�e�Z,AkP��6��X��1U��Z��*�b0�Ō"��"�
�(�Ī'�n���������=��L;�n�Iܝ	����5�$�p���-�<6Z\�'���Ca(�xg۝BΘ��/{x8�&��W%y�G9ڇ�%�����|�îz�M��s)t{�MTm��۞7�(�z�{�3���Ǉ�-X�����Ux*ɭ>���L\렜��hgB~�q�x�gt��1|��*�xt�\g�Y��o��r�F%#O��E�x�q3�ӊ�.�Ϲ������3~�_�}�F[�/��c����;�O�u�:TI�*n��1S����oj������̐�Ks&���qc�9��ǳޯq�ut�Yu��:�8��Cܢu*q�w�]�#S�ھ��s^��ۇ����~~W���;�,-�P�~�������'�ne��u��쭮|�]\Lr}�z@ݔ�_��}pQ���q7/֑��GY�A���[��>����En������`^T�3���As�r�j��{[���5��`��Q�zC/�.':��<}3'sRS2���ܟ#��(��s�:0�V�Ȁ����lq���ǯ����݋�
�g[(}�xFœ��
|�~��P��exEH{q�C=�}9*��ú��8��|j�uA +�����{���1�.�i�tU�4y��4�A^a����^�;�7�k���[�o�7�%֛��b�Mw�4���=V�b�z�̩�����K^�Ҷu[���
7Roi���3��N�a���c�;�5c	.�i��
�1�y�WY/�gDӘ��u3@�,b
[�5cپ�uw����Cщ����|�yN�&��|=�A��� I�9�u�2�L+�WI�~���:����y���Щ�tg�y��y�A�P���QbJ9s,vٛ�=Sr�혬�z�v'�ܥ_����x>&{r��)�ׇ}�U/��yT5�nd{E�a���Q�nteX}~��J���H�
���3�C��������p+���dzu�M�ޑ��ݝqUg�����/
.�Fr��xq;��>�4��^�d֕y>����M��,�\���G���&��V�#h;2����&���؇���2 �\��~C�-�ZC������P��~����Hw���ͳ�+�g}����^G��^�ք㽷(���%#q%�=UC�WL^L�>���؇�nw���u�3k�k�_��n�����:�=����Yhm��(+��*jK��j�y%U5�z��+ўΤϺf��^�x���+gs҇JU�̲����������mr�hّ�z)��7��w�c�O��؏������qȍ��7�_���1Os�H%���a8$�3^���)�+�\���|;�Rw���^p�zA�hu ��ۺWR�� �m���+�`E<쎱_
+r���s�)�}]�f���q��	��s�(-WD_M�ƨ)��Pud�a.���5�\��J�0���O�.�.���
.Z&�X�;��܇y���~���uj/Y����`�z:��b��>N��χK�Ř-�`�{J�A+�a�Q����1e�)���>���^��i�,r�eO��F��fA%�B�h��Lw���/g�D�Wf�+k&C瀠"�,x�O>�������:�7�(q���]��PDǃ��qT"YB ��k�_�j;�uu�9��z\7ش����vDQ�-��~U~9΀�g�� ��,Y�� �/�-���˱^�;�kIn�!��{��_[��Q��}Fҗ�۳Q���V��P���Tz�<}�I5�or�z��u����n&兛8=�;�5��fk��Ǯ���/U1q�U<kc�蜏R��-�!���Mw�|�T���/NDI�;s����2wO�2tV�.Y,�����<gy�y���9��{�g��mX�t�1���nKgnv���{��l֝d���AP�����Ϻ�`��Xܑ�{�M�y��,�(_��֋X#1P��}��v�2�d�?�t�WXq��Q�b"��9�{���\��8���Ƿ�8��5�twճ�CS;��� {�]6�w�wl��%����ԆGs����B���P-Ժ}�4�}e���;qtF� ;��L����.ս��D��7�ү�c��~�^��_lG������{6���(m̱��{.w��������W�]U��z��_��\d��N��'���O�Wz�7O/c��G��'5꼣/�nf�4X=��S��~ɔ��"]?�^���޷�c��+�G������x�g5�q�P�Z���EחYEi �p��e�⧗��J���R=k޴=�ϙ��C=�ug��Z�bp��25�.帾M}C��=s�K�Pz@�3�8Kea^/q���i��#�$]������W�q�"�t���xSEq�=�_�<0���<75�n��Tb��,.bT>Yu$�j��L�_�ߧ?C��T<����H�{�H��ED_�܇���4󞸙�>��8N	����_F���^C��< w�g|G�m���>�^*���������P�ғ����p��:��m�v�.����!�(+�f������_��ȅ*����P��U�q��珤䬠�tҩ���&�<����e�d���ݟ��Ǒۉ����Q�.V��|{�6����bs驃@Y^��*�&���yI����t�k��9v�Al�UA��Kpf9���/N�|m�:�{vu|,8��U�ֲ�v4j	���uF�K���&���Hq�:f3����b�}�K�8�9|����wuG��\Ɔ��e�k��-S��N��x��+�/d�>�d#�����ζ�����ӡ�wD�ωXzO�뛨j�K���{\�3K��tN�~ɞ��w����H�u=�Pw�#\ߞՏd�A@gd�;q;P�q��a�f׸�l"(mw��J��՜��Ľ}�l_{���!z����yQQ�eؠ��po�ޓ�.&Z:va�fF_z��Gz�y�vgY9{|��jS8}W�Nu0|���دO{�*�߶��]���vj�`a����kM��mZS�
ϥΌ�ڏvO��Ɩ�n9χ.�x��G�}넍�⸨��ns���cT�ã��UE���b�/�a�/rg}0{�	r��M�O��n#���R-].:�O�߲��z���Q��x�,�)̓�,���b�ɝ~��ۤO;��W�ǌ���#"k����`X����˥q�G����uj�s��񅑱2�I�*n��?T�>&�0�\e�������P�y���ǝ�#������_�Hw�WlU�N�ې�@�;�a���u�n�j�,Wj��d�a:9�}pQ����|ϩ���ǲ7��z�^eK/�����Ɣo�'H��P��'5V�*��bP�ŝ��W��跴R��0W�k!�F�ɛ�.�e�����t�����:�=b=��w�0u���YXա�����v�ח�w+�ls/l��������OZvk(sq��o�b�]�Y���lv;�ܟH�h�[��ɛ2=��7�KGۑ�
6Ҩ��������y�@����{,W��t]�9�
�U*�� ,�����}j�T>G2ai�R�_��n���Z�ȃ��%~G4�:�ɋ���p�W����ydWeR���>G�鉅�D�9�wԸ��,eB~����=꺮j�oy����x�m�L�O�@~U]פ�nKgo麇�>&6���q�|;�xD�1'��yd�g�T뵸�N�N���_�:�ȉs�zǮ�"�<�)s>Gn&�^V�l���<n�ag��C<�k��}�/��ެa�B|)z��y�����x(����J9L�۠���긫b�����j�{�������9mB�ͯq�/��ʇ�]x53(�}Pt��˸�D�p��ìEJ]���7�7I�ư[�.�q��X��b(Zd�{�`�>�ew�2��|�q���fk{�ɪ�W�v�Ŀ���g�ѥ���~�`����7�t�9s����B�����5{+���V'����r�Zk�dAG��`���"��������;�u���}p��K�u�������vخ�[��Ͷ�yw�L���P��ަ�^�� ]u':\�Pl�gv`�Dt��+�⦺�7շF�w��v����kWQ�c���s�Q��=V�rWoU�(�,�����v�(Q�A��=�C�۵;�i�P��H���zw�9���;��(��0JF��𞸊�~5��^�>��ٝ	�s~��o�Jf5��F3����^G��^n��ѐ���[�C����\���AB��C��ø�������㎼�=����;���q~���*bனg�;#��&;)�ʸu�o��5�8Stx	������)�q���;��x�o�x�o��jd��I.�0�`%Б��p�D�U� y���+�]
��o�<���!U�|&�?[f<}���=���#3/�瞘�^�[#�[�y��W���`�x���.�%x�9����]x7��a��u]s��9q���t]>�}^�c#ޔ\�I»��\^�sp�4w���^��D��O��M����/h���������Y�u!�z�<2'ʯ�z���z��dO+�h���\���з���FW�w!8�r2��<T����&=��~6�G���Ϗ� z� ~�De�QdȰMf�=�w�|�0�\��6�f���h�V�d��^�Q���n�F��=�:ȗuQ�䀚��dTf��;:F���Y��n�I�,v�����,���JT�Y�m�F�>Q�Y�E����`��*�"��u��Q�_u�:ӽ�)AG%ѸBdcg>�w�a+� �[T��t��*vv=��r�ar�#�{���=�e�����^mhw��3_wSfo����̏d$�ϦI�c���}U�;ܺE�ϛ븫��᯿2���s�k������Zn5��f��=k"w�"n���EtMtj�F��'\���C�}�ʱW�m�1w���9�N�<��f�i��T�Q�i�y�'٘�x�r�`_���H���d�μ8�W
c�:��$zݴ�z�"��r�)�Y�z�f�w���z�j�޿~�����×�Z3����%޳|��'HL{�k�U�;�Ǩ3�裃��Wq�ɝ��>	��S��ϓ�_��x���G��loY8{E1�o��i����� �����( z��L_z��d�s�����U��>���>��*o���Z�=R3����mvu�ЅW;A���i����Ó˼D���L	���7�H6vNw�޴=�ב���>w1�]S�{�o�N}	��#�o����w�>����a8Z�;�B�Ke�x����G��������s΍�����}��lg��Ƿ�w�~���)�bX[�L����"U]E��K�Jy��J�#�:{k����Z�蛼�&#��J�ѯ���t�wHe1��0���{vx���7�v��vѫ��
Us:�R�YB�gR��|f�w�(��/�r��H�Z�ݍ��-;��K���v4w���";PiN�2�kD'��Q]x��ΥR��Dȼ��"]����_�"��{i�������^����8�\b�K� ]u�c7�j���G�VnM�}gIc2�T?�׮&�}ּr=9\
��@g��35/��*];����t��>U�}���LE�"��9���8�^��'�^S>+�Ϥ��	�\g�0���z�0WD�_J%�1�v�鎿��C��ZdTk���E����a�<����hZ���We���S����p���9.tz��Q�>%i#��M�5q��^���A�R^���)����'��N!�ᾍurX������y�=5��ǡܐF�+�%���^��0��u��>f����^v�4}ܰf�m +�V�����9�DuD{�v(_��kE�zO�����R瓷�ǘ�^�9��>�u�ڭ7�i~=9��m߉���Q�;���^��/�8�Ҿ�#�e;���ɞ��e��g&8=��͔<�r�p�q��n�����J�jw��
�1\���
�`�z+ڶ��Y#p��p�CۓZ^����A9Ϻ�V7>O��o}�+��J�/���L�}�(W<�S�[�q�3"tB�X���]f����t��oS�p�ϻ/sYy�P�!˒XT%�#��B���7���v�=����eN��1���Vp�X@�8C�@ �[��jW�!�(�ٶ��T��1��Vw`�Z�7��6�n�w>�|{��G������Z���R%���d�F������_�*x���hG��M:�B�v+�'^g�G���Ͻ��7
�\nG��>0�be�O�SuL	��|MN�+���_��nW�L�,�+��gޚ�>��^���W�^n��c �.����<z�&}'̏2Mv~�WO��1�L��x�}PQW��#�z}�흤;��	~�_�A�G՛�L�����~͇������M�M �(-c}pQ�����D�ZG>��#���'@Ǐ�l}�'���o��+���RU�{7L���6�����/ƽ�\U���Q{^�����~�q��idߩϠ��+#���t��[<`�����&��Ҵ�|���@�s!��ٙ���}�}�=�ߦ3��霟N@W�e����(��-����^&&)��3��=�7Ig۱ޜ��~�j�;<��࿟��mO�b�qzt_��x�~�'ȭ��|�;�&�h�i�F�2�y	���'^�ZV�V��p���^�E���t��c� �Ey�(�����]�X�F�uP:h���Ϥ[Lt�^RpRW��N�h���UocGR�/)��̓�S�B��fZ���w�A�F�:[}��p�ojP�S�}���-ZЙ:�]��{,`�05��
	��I����T\t��En���u`+�a��Ҙ�����W�Z<�����q�)7O��F�}0�Z��SR�90Q��Gٛ{8F��x*�*�QT,d�ZM�v���qU������{��%�f�r��]nSӥo>M4{�Y��ܘӥK�����o�P3!�qHj��W7\V���Z��-���nc͆�;�R\�w�������좳>@R��.�=}�T�[=��賻�0;�:w��X��3'	��aX�X��d˲�c�!7���:E����^�{�{pfF�Ue=S�Ԗ��0��9H��}Ū!�N�wn��47V��H'\@�´�X�s�wR��bK����XB�.'t�H�����%����Ny�}5Qa��{��(&3���u0�'.�Y0�Kb�4�xk�<5a��� �<7�;�[=8Tu�����)��`��$���5��@RH�nU���}�`+�p�Vp:�#`�o�^�9}���r�3WN9���/�j�;�OO�,��0��ۚi��u��<�J�*dE�F'pz�͵�wE�$-�Ǖ��V}�=vE�wX�<�d��{m�(-©/�WZ�+���P���%̠]c��]w\��Sv�=/z!]!P鸓=��Զ(V�["ӏiTwMhՔ�\�N�4V<gl�Ee�͎Q��ۗ�����[!L�Ϛ�NJ�TH̽��Z�X��I����LU�Ro�$�%G���)eɘ��������b��mF'm����X�-���b������}z�XZ��.aV�3:�-
��v�y�s����᱐�������'T|��Mϯ��b.�'�Κ�4{B̬���sn�jD�V����Hsx�� (�D�zy�X�Y���Uaa/:�:C�������,�Fj���cFH�wQB���oO۴pb�n��NJ����[�}��fj�j���Z��&�&]q�S�N�j9ث�%I���ٽ3�T�^��%�W��ɹ%`���ثqw{r�T7�8g8����v3.��i8���tke4-J�.���PÍ�ۺx�uԬ�u��Z�[�so���3�N�w�v,/o��J=T���B���e��{�ў�IN2]���5`oa.r�J�Wo7)f��T\#%��E^�x��9V 71���Un<F�uJ�y�+�}	F�������߸��jW�VUꍊ������)L���R�]l�]�{v˹�;!O.��@��&�L�ޕ�wT���7]}��Q^&2�j�	w.�Z�f {�J�,!��j�[��m�����a�޼#mt�Z�\:0:ۦV�����HЩe�();������O�E��M�j���}���R�,�X�j	��wH�X��wp*�Z��IY䑄��T�ڴP� �@� |���A��֠�++JZVT�������)-�1*
̥c�(1clX�
��F�"�V�UV�S�r�[[+PX�-��,�1R�B�UmY*�� �"�"V�ĵh�m(���0Q��֪�YX�Ke-��,b U��UUZ�\j"��m1�Qlj,�����F	�&S2��VQ
$D�ʊ�,R�("���*�(����-��1dQF$��U���UPP��1c#Y*�����,���m��m-�X��*�B�V�1Ɔ6[� 6�+PUkdTE\[F"��-KB�
�V(Qm��m-T+
Z)m�U��`�-Z"�X��*(�Um���TQ�J���ְ��)TVTUEZш"*��W)�Z�
��1k+kJ�-��%���(�+D**�j1���X��FD[LLˉ�2�AQEb�(��Aeb��P+��T���E�@V0�V�H C��j�y�5��wwv����y�{5�0V���P�!}�f�pAyҺ��7��먣�:��,��K�9QKn�\v^)<�~#k�A�	��څq�K�q3ۗ�����ߡ�������|��̋��}���co;ޭ5J0G��oIӗ3��챗��r�t1�ﳥ�P����~�ew�{�OVV�8ux%R���\U��7����ᒖ?�Zxz}k�xg��3�z�6��ߺ*�\O޾�����A�{��(~��};���dAF�^6!��=e����g|E{�o���[�]�ꯙ��;��������W��ۮ~����F.3�nK�z��!-V��d�V�ꑐ��6�|�y�J븗���b�->��:�=^���m�BPW"zv;)����b$�#n/ugC������ )*�oђ�v���:��q�{No���z�4'X���(�����f��}Ҷ�X�}������2)��7��w�:�Q��~y��M��}!��u��;f0h��%g��ж�e�Mx� 6F�5/��t*����X�;�>��\'6�����&<���֩�;ė�Ǘ����F�F����Aߏ�?Jf��mm���!.�u���x�آ5�g�{�Xclm�j�+�=�Rh���s���"t�U�9�}�8��F��i�����ǘNnB�c,��:ga�P�lg>�[IV�Y��ŇxD�er�`�E��]�,J�c1�st��]��9,+���[���o�N�4�,�7[sa��m\w!�t��ͤ��z�{S�
�n�,o�RqC�[����#��>Y^���䆼�;�#g�P���圽���}㻟^~�΅>U~8}��Y�^���pF��M�Ih��k�ɏ�o5�9�Ͼ�	���V����F��oƸ[��ώ��Zf��B��cc�M粣=+̍�lex�>�cv��c�6��E��Mf���9�5٨|�F���q�Y>[��h�e�K:��,L�F���5���^��\o�af�ћ^��3+K7���<4�
��&=�u���X��'�vc�su<o|�2=r������"O���v�?_�;��tNg�2-<<jc���H���3}�y{=��㎘*;�8�{��U�m�1q��Hh���Cˌ�qc�|�=|]�G��ʧ�������}q�~��?I���9�\:���B��3�V	�7%�򭉇*��V��ys�ڒ�A��&�1WY:�}��f;!���O��=�=\�֖w~�<u`"E����eI�c�g����=7G�Tb��_�3����3��9z��{��+�=��<�8���X�~��CH�
p]WEO��ȡ��F-\��;3=k]?\�=��!�h@����!1�7-V��o.�J�WܮbZ[�<5��m�L��C�L��i7X� ��$��TMN�J5�X̊�]�x���]si�<f��;���*��TR�a�E�*��زf�]c���j|Vl�*�3������7޸w�Iφ��/����Xx�]���S�A}C`z��.s&�5��q�-���JU5�,���%���2�ȩ��7(6^���|�i#aM�yV}CR������*�9��>��Q�W2�kq.�A����gĶPΟ]�Ŭ�E/��C'�n�g�C{ͼ������=�Li�Oi����e�#� �5��PK��_�]t�Ryuy컕�ǟ�Ǻ��_�̇�<���~�����o������[��^���Ŗ]߃ƌ��z�_���D�F���Du<8KGw *��o���(�S���xc޽ 7�s�0������7�<����vI(,;0X�Z�'�s�v��(���~5?+���z�Vu���㑄���b}�zI�;��e�j-ϊ�L4pԱ��!��Zdk���E����a��{��1v%�5g�^���d�?z���2ǫ��d�gļ${�50�fއd�t�i�Ӷ��l�J��n�O/w`{����U��^��/�yО��ڱ�(�+�	Xn$�:va{k<F񛧳ym�����$��r�!�����u�R�h3u�m��H̕�j��N�%l���ò��j_,��;����}��W%EG��U���� |���]e逼u�Hᾥ�%&�<�L�.e��-�֎P=�[o�_n�A�k�Ee^�[x�+��j�1l�j�J+�5���S�׾�`	J�~�:��'"<��W���b���8+�'N_�Fv��O�C�M(��^wF�>Xo�*��n3��כU��O�zo:�m:�=�̣�wMG�:�TKѳ�ܔ(D�q=t���쓧o��:|/r��a��,��u:����+�9�s��SWW�WH=C����Մ~��yQU�k��,;5��bfu�y5��d��`된��U�凢}�Sݛ��D�HW������;��{��;;�r���R%����1s�,^L��ϼ�G���h�T�Me�ίX�K��y�����9�;�x����^��w����G��R����^�Ɠ���4�
V�'Ћg��۸~f|����z�gѾ�\{ޟsU�aw��:�>>�����={�(h�MF	����L�O�
5���}M����x%Ӄ�^�6=tn;�#�sº^Fm�Ԛ���MA<�ό���H�v�>��T[J�n_�#��g������t�=��I�ƅ~W�C����)�(��,���2��]���W���������oʼF���Lm	�o�����EV�P�ʩ����1D����j��x��ީy�J��#LF�6p�����Nv
��;Y�2v�|�B��M2X�jT�X���݊6u)�^�'s*�a"����YH%g��+����)V�t�冷{�h���(��ޡ�ٷZ$;�r�+�'�j�@��	q�,6���bt{s�.�Nz�|<e�>Ѿ�>��T����zb��+ޙ>6�{2<�IDܖ��õ�V���!�s�����U�)�;�=>�9c��6ẹ8/��W�<�{eD��=c�d��(}�Tn�~���<��V�ne^���w�R�
�1�I��>��j�4sד~�T||��/.ǆ���~�غ%�<���<w�2�����ܘ���N���]B��{��uR��+����{�=�
�3���(���j_�a��x\���yԶ�����R�z����lz�z������}��o2�V��'��t�ouF�{gM��{M��P۝�2�&��>�u��J���\�ɍ/(��>��`���mk<G�]����qV�l��`��C���Led֖@�k��`/1N�w�[X�oya�����R5����ǽ��C�=�=�r��_��/	�V�j��5��X�6�D�B�g}��ۨ^�������o��ϸ�exs��0?a�n2�UP#�E�ˬ���aA�Q$�;G�p�5P9�΋�ֺ�|����|p�M�������s:��T��k!�ѧv��پ��o�[���b�j��[���;�� �����MY ��}OlL���9���J�R���w;,����B�<�JW��;	f�>�}xj���~���\sN�ڠ�V�����}���m=������zx���\n��\Uo�W���V�	Tg@�7E�Mׁܔ˸�V
)�Ty��l�{2+&�&��5�� 6���e,�M�3�y��:c�VT���Q�W^�\�M�KgrQ	ˑ���뮩7�=�y!��O����0��_��^���ŗ'�@H����v�@�Yl	q��OF��]GwA��>�/ܩ�\G��q>�E�{i9�5�{2y.j�T��������ٶ'7�1�2c�;�zF�흁��?RE��*����{�Z�+�'�u��z �5V<�`y4Ug�Uy����1�&&�մn4�ǻ�z[�ʯ� �������b9����]S���棙2<G��G���P[����m�/ղj#K��)t�+�Bck����\�K�X|��sw�`vD���{�i6ϋ����F���l�}�N��l�&M.�<x��B�z�����l����c��s)����ƪ���[WS�����ӑ'���ׇ�����'Ei���M������Y�}��E�w{���ӵc��D�ϻ��:V�݉�ˣ��'��m㼶��s͵���J���w|*u�t��gE�6����:�ϧX��Y��Z�3q�d��*N�W4/�;\jo)=�zk��N�4�����ϣ����=����!��ʱW�m�1���Ih��;P��<.��/g�]�Lr|�<���75��7��������Hϟ��'"<�_�Z.5��=�.�VL+W�ݾ��ڬ�de���P�;J�����_Ro~�{�]�:C���0¼�?E�e���������GO��gT���󾒝��O��eGS������q��o��>]_�3�|���i~U�� �M�e���pZA+�e�_�L	��\;��N|1����U��b�=�t�j�IӔ:���Q�,>NS)����ڨۆ��+H����S��n2Pl�F�nb��2�=��OGN���^��
�h<���z��}�O�۫�ǫ �,�_�%Ѩ; r��Qw
��TQ�}���vW]5>�p�ql�rY
���H��;c;�+�f��ڈ���g���!�u��gzNz�紩�!y��0�Y�Z>����U�Ǎ��[/�9@��=`h��֮E�}fI�.���{��C�-ӣ*}
 ݝ�� y��S@>�Y�Z;����U��Z��NW��h�~����v�+������9��Ն�#��y����`|��#���0�s\�����sT+L�7��"������R�X�=fZ�|�L�}ENN��e�v�NP�i��O�6_C U:�Q��(�)�w�3F�F�#+]����Χ]n�Sy��|���~��:�oϑ����>T|?:��O�p���
�3�>��)�r���9��ԧ#-�C���q� *���$���ĳpf;q7LvzH}+L�g|wn�P��#��
�����g����u鹋~t<�%ΏXwD����#���CW��]��q�{ᾬ޵�ynߐ�>�ޮ��=P�\����dg��A)ȏ{���TA@J�I|w�����=��(���Ӿ��C���׸�s�j���J�~�%���DuG��b�����LX��b+��_����o���ٍ�q�rzmx��i�/Ǧ��[ \.�~'>��Y�y�O�{�=n0F���T^^+��`�����:t�-���2��\g�Y���O}�|9w�Ĵ�{+��YU4z�.���L���넍���7���F鿥��Hz�kK�ɝ���렜�ގ}�Uwo�Uޡ�N]�r=���bΣQ�{^G��F���,�=2���,s���e5����꼿x����)]p�Oz�<��ϙџ{μ�l_��nb����_lL�Q|����������GZ@��|T��q%[{��;�w�XZ�	��-v�v{/[q����+Vx�9�H��T�b��mZ�PE �7�)�M��8����<\�x���Vc����E;B�hVc��C:]��c�{��7�Ey�8�`��V�+�Y��Z�tyJ��K��}����,�ݞ��d��3�(z:_�FF�E4V�z�:�Re�:�I���c=^�R����K{Ô���1�)z�7���>}pQ�~�d3�l��%����w�vcA4�>^�.Rɞ�
��U���'�,%��	�$�nx�O�����S�/֑�U���ǲ���*�m��'E�u���Iv������.|�d�ә���ur�F���������^D��+�Jv�r�8�sޑ��{,��.�'�KG�^߭Y�x�+н�One�N<7���*9�P�'����ʯL\*^�>6�{2���OD����u��^w@��.26�>�2c�:7��=�Km���m���y��J��8�z�*<�)�1܃�`E���yW���F+�+t��='�K��j�8_�ٯ�y]�9� y\�ǆc�:\����ݸ�fz)2<G��t�̡�pf��ݨw�m{���n\?Or�<�e�?i��n^Exж��wEk]0=���GG\�>���p���b�l:7;/K��7����~���o�ǿ?T*9ϋ�P��1`���YRp~�^����Xr"�g��C���\��vc�oo�ɠu�u�!oQ=�������Y��h�}xa[����IEu�KY���q_.�[Λ9Wg���&�������t3C"�sF<�.�А;�z���?o=���N�uDך����=��҆��1�U�a�5S���'����gM%�]]�9>ӡ��VN3��ޮ�q������N鿤�>Y�S{����-��2����y���s)����Ϲ�,v|���G���;Nto����G����)YOj�M3ѻ�v���H-�H�3��ׅ��;�숭���ov����>�܏e1�
����"�����ܻ�k�:s���敚>�~��!�f��O�޸xP]��p�\�Ty��{No����k���c'ҳ�+Wt�s����՝|2��ǳ� J�3�w��)��;)�x��Fտ,�{9��ؒ�O�Uk���ω�wNDqziջ�ϏeJ>�@l�A��׮�-q�Ǚ�'��U#~���d*o:7�w��7�����U���F��:�C��(3��7R����޳P��V3ԫ��qó�磧��{�W)��a�%�HÃ;��#�.j;~�}}��˩�t]�nw���a14���%#�
a���GAg9K�5���s�z�sZ+��$��BH��BH����!$�$�	'�!$I?�	 BI�$$�	'�!$I?���!$��@����IO�BH�p��!$�$�	&�@����$�؄�!$��$�	'�!$I?�	 BI��IOHIO�1AY&SY��^z #P߀RY��=�ݐ?���`�?z�T�T�


�T�"���p�$�)J��URs�u(*�E*U�
���0s���
HPBAP��M�8���j��-� h�Wl��hmCG�ma�M[f��66�ji
p�rțml���knj�m�'s�����h�5���N������(v�ѻu�R���sr�3Z5���ed���u�E5��Z5%U ��(+��d��'l�փPi�p��[EKlIM��PT
���DJ��m����,�    �44��I�4h  hO$�)P�!���dh�@s �	������`���`E?�$#&h�h�hɣC@1�`&F F&&	�bi��Q% �i4��'�d��123MM�'�����o��k��_F��'�ag� $�撠LB��K��C$ 	,��_����������g�F0&@ 	��O�� ��	p@�E!� $�W�_�������W��|8  I�'5e^jW����H}�۽�*QB/1�]��?�tӂ���gV��^�7��Ka�
RͦC&��L&�����NCa�l[;[xΧ�kt[�0V��6Mcz,�!�[�[�v+E\�iB�ۖ�H%bG�5JpR�4��F��y���yjX�$�M�Lm�Y{7mʆ�
D�3v��r���ܕh��˭5��5�(��C3u�t�M8l��j�طB�uR��+$�e��J���-=��^�&����1RTL�.LN��j�srD�Z����l`!����($�p�7{{�Tj�.�{�#�Yw��c+N��y�j�dkŵ2��&:�*D[�����G[��YV��"ۻ�,�e6V�n����\Jё
Н����˘ �ֻ���:��t+�D5�T�m:2>�F��CI;���yP�E��lJ���m��.�%=-�In�*�'�X�v%eg�9Y��WIC�L9d)�2����Ǔ]�'m�4��[���yqm�[��ޤ�h�1Fq�-\È�b�@P ���X�e��ޔ�^Q@V�@����f��)����oT��h7kE
0Yk+Cu4Jm �s4���L�bV�&r��l�>��ci��fZ���Ӻ�"]iԕ+�F�N�N��6��6m�Xʎ��100^�ou^3&�P#5���t�Vj� c�s~L ѻ�Z���d�M7�`я�J^��p吪^)7C�u�m�Ok.
�w`�Vf�#�1�j�]n�эh���D� �A%��H�xYq��t�%
W
��R���t��#�z��`��M�5Zn8&r�⥗�v�[�հ�ض�Ie�Z�O�C8-I���U	����a�$b4Pǰ�T.CN�X�d�`Ub�Yv�GZu�@[���T�
U3[��$�&��fő�3E�36a|/&$*}tL(c]�kl��JB��
�1���PZ�̣��mS��CN�T*�ۭ��S���L�(����N^����V�l��z���gj��M��:"�����%�w�(�#7xI*T�%^��p���u���J��slVևx��5m�¼���5!��UР�*�V��a���ᶲ���"���Y�i*�@*k�K%��À���ةeV��3`�S�U�;+#�ڄ|��d�;�5��-F�S��f��Yr C�V�M���js2� �*s��Enl�;,Ht�[ �;N��g,el L����&ǛF�bZ�Mz4T9�*|u0"�/NR1�����Ȗ:d��5��t�[l��:ƭ[0i�/����Ka�m����W�V*I�suU�RҀ��s,M�ڋx���îP��(���f}����X�̡��)((f�Q$�ټ�2I�L�e�YYb���M��!�2���  Sn�Xۚ��V��������݂
ؓ���Pނi�ȵ������v��ҷB�g+%�r�<��5�j�"`J�[Jb�b�r���H�r̊V�`i���J%. �W����iQ�b��� �H��2���~X�RK�#*�,��	��l�]�e��me�Z#Ba��зL��Flܼ���Y�&�^��������8�%���#����,����g϶�y?p�J�T�Ѫ�K��l�!u��H�֊`��!CT�\9��e��m����Yu�1�k��-�s�滗O+�Ӥ��n�O��#�2�]ا{��]B}�K�a��}GC� �>�1�ζ���.�K���9�,�|�����xS�5�v�(Y��n�z�U�p�\��答�p����S�+����S�5
$c�K ����|�o�@E��Ю�RY��ͫ���n��!4��֝�)�g\r�,��J��Ц�S�]�;5�A�">ҳ�"�j��ʳr"�w�u�t��>)�݄Q�6v�1�g|��j���C ���9@���m�̷9YR0,��,1^�����Tmu�����J�Mw)�9m��F4�/���I�� �y�}���J���Ίv0�a(�\S��Jf���ڜ�3��FbV-�Je3[�nt46&ta�>�#i�v�gU�l�SL.�c(�m�i��v.���4�v� d��"gZ���`������Ѣ�����}���x燷ew#�ݱmE����7ro���+������7ڴ��0�NS��I7�:t]�C��V�co{3���Lc��Wl�mL��v{�DB'\�/7f��2N�ǈ� :�������1&��gy
`�O<���6�9�y�+��!G��'�(^���3��<�^�	�]������jrv������B�M��;���Z$Mֲ�s�觱X��jpxss���)��b�`���%�V%C�r��GnХݮ�ó3L���S-<p�ER7e��z�5�(AًekF��Te�k�1�:�b4MK�u,��#@y]���&3�ծ�HȖ�7�9��o{��)�J��7SX+��R:�.)R�G��C�>$�TxF�B��f�*^�bi�����Rљ�V�����u{!7C���T/y5ۣ�b�~�J9qq�E��Od�f���@��
�}��o��8���3����l�5�V%Έh�\���Xy�\Q��y���DWkCz���W�lLTy�)��K�R�R�s/3j��Fr:�:��N[��Q�3uJbvQ:Ӝ��X$�fi�՝�@����ׁ��X�_\%��x+�DR����[�Wk���V�q��l�/���j��oIغ[�M�V6Wd'������쾔%�]%�<M�}E���v���3��(g���ʻ]���m[Y|�[���]Y�XOJ9�[N8�Iwm
���`Zk8Qv�RB]N��4b���Y�/gh���R԰�Ȭ�B�j�I �[x:��"�=���d2�M��B�3V���Us;o��P<��ZF�G���o�Ѿ�9��1�N�c�oP\���0Ծtr���0��9�%�_ݜ���i�Z��N�y���g,�Y�$���7�Qi�sLSz�����$��})��I;���So�6�9'wT��������|S�x�:��5�}�uc��X"6�TH35e��Z�*ᦶȇ�S�7��Y}YV�Y=&�W�v΃W���O>�ޡڤ�c-N��Տ{R��_n��I_u�u���f�*�'+��p��IX�]"i;�{�r�rJUX3�kf���>�y���綮�%~� $��%��� $	=kw�yː 	>��h���������G�3p^��wr����#t삤��;��nqo�&�{����h ��������<���]|d���b��^��.W["m;��w6�S<9Z�����7at~��9J��UwB���N��#9<��8%�P�Z�8���';G��e�U�[u�ƽŦX"�n�ѩ)�-�p5;���n��*�]\��(�&D�DI�I�}j����!ov��k�9�%�Åc��ii��{�ٌtS��mV��H��ɤ2�f!jP�A��ˑ��4���w����9�lqڲ�k����,�ך$�S._�|]V+U�����{\:w�ac�Տ�㭻��\��l�lX�[x�t���{�=vG���TTWvT��=\:��
ky6Yȅ������;D�=H�;JƑ���
��r"dB�6�#��a�	�j,˫�}J�xNА�gOϱ�4�4�trb3<d��.WܵB��S{�^GD^B���_%�����Fܬy�ku��/N��|�Q&7C�Ȫ[ЭY�[]��'.�e�Md<��󵮀��_V�=�IY��M�:+3�N�M�B�+���7�!�+0�Մ�y���Ս;e�·A��ë�e�<*n�AMȫe15�7�|�HU��A\:ČHh��:��喅Z���l�"f�`$9'K>-�J��̣N��VO�|�r3V-7��� ����>�ܮ}�H��ц�� TF(�Я���q۳�������`��S#��Tyw���{����mN���;PІ�P�L�pRT,R˗*��)}˥C�cÈ�=�s#�9-��z�
b��X�g8�饌�{�,5wG;7!\�]��6`ӊ���8�E����|#�+wR��UYm�b}sR�[�T�#q�aC��؄E+B���Z@�v�[���[��L���M���q9�ٖQ�QY9�8̃��k�6��*V �&%�[��o6�ih�hD���V�7k ��k[����֣ôS����Jf�${�Uԁnގ[�xӮ0Z��)���빜i���\(�W��kR[�KP�7���5=s��7��a��,��۝�wq�V��]���.�(�u�tV�-��9�Yܠ�(�3
�Yo�,�.�*�@u�Č���	�k��v2�f�xɻeI������RT�Eq���+(}��3���l�g^J��j�h��G��m�(�e�i
�a����r�t��ٱ.B6�Y<�Z��4ȤrӠ�Z��z�S���7���	#�����i:��*k��2ry���QWkO<<+��uV���co�oG����.�©�'��9` ������5�U�7��n�˦nY��[�ӌ�c޹ĒX�h"����yOP 9B�U�c�^dL^�;��>�N��f�b�s*�Ӻ/K�<D3�N���uf�M�-P�6{k:ⰺƾH�$�;øi\v����z��i��#���IҐ��X��_^�(GlQ����f�C��쇮�&YC��+�˛��r.�Md|��o��  �� ���
�cH��'u�B�ʭǩ?}Y��I�,���\��UÞR01�ek������/<ܗ�=x�D�bWP�����D���єݚ._R�$o+2ܠU+-��}"�6q�P���[Ů��#_i�.>/�b�/,'���mŠ��ֺ̥�:���kvys���9K5���;�n0�_l�C���Tv�-�����{��Z��ih��R��--Kb�D��:�E9�9�wgn��\�k�,��M0j�1F�R�r��l�JUL�V�U
�[��0��7Tȭ�[B���,�qwkK��K��e%��b�uEEb�Y�alU�E�B���"hD;v��1:�?g�}�z��BP�ұ�
)�U�?�O.�ʈ�n=98��zd5���-�3^!��t�VX��s����x���:v�w_t���\Ua��ܾϘ�������iz(Y;H���8GW^�x���Y�ۏ>�{k�~�8p�$���2�J7�6�"�Q*����l2?ʱ�������*��J�������:�]�^�X^P�>�'x�e�~`����0a�4�O����q:[I�����Bg�����yOMHXi>?Y��R�l_.B���:��piщ�Q�c���W;�5��)��Z�*�;��8;��r��v���&K�G����*ql�b9�칺-�2݌�)Yڶ�s����G6��o�j�X�Y��Z�a���0u��g��9��v��^����Y��>�%VB��f!���=���CV��X�
'�wj�ׅ�H�!�=�b�*�+MehaU��8ĽvM��Hv�F��%w_q�D�<9���J���<���M��L����\ޞ��KW�ꃇl�NE�r:���;~�{D^Z�u�\���a��]Ԟɽ����E�S�ǟ�]�sk ӷ~K��y��ʒٖ�,01�q(���>��7�w����`y��K^��)
�ζF�\*��kcI�_wHL����d;�t�|Ӝ��mj^��{EM�������.-��Ϟ�7� �t��Ǎ2|<�38H�M���2���3)��g�_��d�	P�l�o�����OZWyt�#���5�]���z���>�y^�r�/p,�\͈^W�B������}�C���[GU�kw�9�9�J�p���k�Si���Q�,o&�tkh$�TaP���ѽ�ȃ�Ϳx�r�1����Eokf��)Y(xfx��^�7ִ7���O�<��G��o��+uz�r�;,�OtҰx>��г媽YC���+s{������a��ܫ>�����W�����ϴ@�C>���@���82q��k��Ǖ�X�_{���,�]�Ay/ Pi�n�СţN��LF�W���������~���[g~�mΝcx{��Cw*��"�{���lꕇ��]�@X�v��1���X�5R:b�6��g�|�7.���WX&���0V-�<� |��лt��X�ll3
��J����|Pv��V��Y�hAZ5z��-w5^�^�~ĩ1޽�W[Ǫ���	'�'Iǋ�;��V�޸��[��l�iQ@_r�O6<�B��Ұ���z�ng//1�ޕ�iG۴��x�i;��@�ס��cs���^t�"Żܵ��u���ITd�4��q�C�Z{ʼשhܹQ���\�����[��o��3��R��81�Uʆ��V�,6y)��Є���s�5\F�vj)�o-�,���b[�#l_

怕���wʺ�f������"��j';�b�1��?fX|���r�zfIg���M7g�c�;}/�p�Z7�yg�����t�y&�S7 vm�Fڽ	�{n��'�-�^Ǐo�$D��"�e�Snj���`��+v�mf9��O0*4������܀e�p�8`�L�(c%G�x$�%AAd1HXv���8�-�����)�	^�e� �q[t�/v�Z4�WR]�y�Yb��A	T�ˉ�
�dR��1�p�r�ȍ�gd;���N�������WR��ln�	��Kb�Kka�����j�(����(����(,-Y(�
`����(�"���%UP�H-P��]Km�WB���)j�UHZK������F�S�Uw,B�EX*�A���EJ(�XԦ�R�U
�kB8Jb��*���uC(R�
VRR)-[����"�U[.&�� 8p[������d�Ҵ����9λ��ZC������_���)ԃ�3�*g)��/�_o|�O�/q$�)��k?-j����f*+�P�ѯ�����]�x�G�r�,G0����/p����i�T5�ag���7{A���T�^�!����[�TU��x�Lɟ�9�p,E�	��w��]���y]Q�at}��^43
=\w�O�o<�\V�]�m�+ڴ!�~~��ښ^;7������79A��I���-�-�p��;;"3=�Ci<=��'��7��e�AGT�|��/��v,<�b�������w#O��R�cM������^�e��'�Q���C�(D�����Ta}�í�=�Fj�N����m���=^�<�R�ۄd���W2n�z��/�^��K�V����MaC=��s���s��1�r�5z���k�^�z���\��7��݈�|��*r��^:c�1m�b���[7�4Q�;��T�+�e���f့a�`�im���@�2��^z�l!L��a�����{Rd�
`M!��c[��g{$"�ꉦ�=$�l� d��H�󗼄�@�Z�-'L��2+0�fv`�0�0����"�}��˃��Ʒ�#C�;yo�-��ѧ�=����դ���� [!I�	2�B39P� y͛k\��<I��d!H��l��&Y6���=�6Hq����ц�$:�C,�C�JI�����'Y�!�8�<C���$:�L�"e S$H���!�M�Y!�e��2�!�	!���	I
d�h�u��YHԐ��XN$�B8�$�I�Hu&X�s�̒,0��!�OL���i�r�$��z�3��q��d0�-$�dRCl!���c����x�Cx�6��I��["���$��H���fP��!�I�!�!�M!�Hei�I�&�'��x�zߘ�g�]d��u#0v�d�/�v���F�&����)w�s�@
Bq�M��2Cۺ��{=Q�!�M��,&1�bE���$�NUI0��!�Bm i���7f{�	�x��G/E;��WJx�͔�k�J�c�i�⫇ں��]Oz;�M����MCf�8J��ݪ��X�]�����a�r�	���o����K�h~8�=�m�S�8_V�r�N�A
��� &���5*���x�mι���#���=��a��e%/E͜ZW�~1�کn�Y�и������Wv2(�BIb�A��v=d\	I>�mΎ���#���j�j���X0k��_	���&Sh5�D�EI]Yo�-��L1��n3<�ϳ�Q6��2�kJ�W�Z+��eY���pp��s<�p�f�^4SβL��Su��P�6����QU���|�p�D��,�W�vR�­.�Gj3�����V�X�-]飸�{b��5	��C	V��0'�����~V�x+_�~�W�¦8�R��w*J{�O��|�o����9�W]���sef9����cЏ�6�o=X���ECŪ^>�.��n�Mu��nU�	�#�vg��E�aO�vʉVf ^�lp�!Se�}v��_�);���W����q��܊!����)���y�_�74w�����)DgN��[K~���E��^d�Fw>gV+%��F�&y_���βM�d�Dd�/'`�>"�5�h^d�q�kD=����ʇǠ���9��2-L\4n�\��Jj7eGt󳈬ҭ���$�>�������Ŝ�`{��ZW�w�5��hй���#�%\�땗ă�جX�a�My�d;�7���������|XRx�]������R���#Q�bGݶ��Y���Kp>��r"���м��}�/��w��ʝ9������ն0Pd+��W3%e��+��IP��J���w���'Vkh���b���n���Ƞ�Z�<��b����B#YK�5B:
�e�E଴��1����O.�@���Q��3J�7ET���VkյN�����4�)�V�6b�xUy���S��r�Tj��Lch���iL���TL7r��J�(JQAe!J*�*�qx�MSJ�KT�4,"+TU�GQU���PP�  (�×�찕?�3���l��ǵ���0g����@���՛�ףsdN�$����Ua��yoc.`+g�zo9Y�u� �u�l\i���ko}=N����L����jrڍP���3�����LgmP߈����By?{5n��k4�V�@�;���u�J�7n
�������ߞX�6�����a��+ȳ��0��8���ۋ�_-��c�pyҿ=�[`p����v�oz��Rb��V��-t�z�t���:����ަ����.)�C�1LȖw-��B��K'��`���Ϡ������G��;�����������T�����~�^������\����@��$�觫��R�F�^�����2�1�s�^���
|�_�!Sʦ��V`/1W
kv5c���ZP�©/�8������~4���3 �7O����]o������.��S��{iA�*� ����T��;T6������;�{NR���3���Ǘv9~��T���4�Xid2"+ٚ�^��X4T��H9����`�ݝ��3#���ݏ�"|��z��w�jtx�cz3��}��k�:��ׁ��&W	���7{�wy�����N���o��dz�A�Ֆ��_��Z�В	�3v"6�V�X����S����bvSX�]������fO �v���m)3v����cc)�<�I4U�Y��A�r����<��p��x�1�̱ *��3�==�s����U�j��^�T�B3�]Y����Rц�jSh�*��T]�]���۽ڸ��k�h�Ce�˴�f`Ƌ�s�?��R�dg?:�Y���d�ZF!Lr�ߋGoP��r�uW���d���eT)O��86����E�����P�2{�i�s�y齈�b�۬�z5륖��o��������� =_���T�L/z�%�i{KE���؂��z������0D��u���G��S�ܱg#SJ줝k`��W6����Э�e`9�@.f�y�Uٓ���ø���r�O"WJW��}�4���f�V�l�o���=�z:�p'�����s���1��{U0���Q�g���5������/e�����;����ҩ\\�R.	��^��ב��z=��*�D3@�ڄ�[��Jٹ�6F��^�jˡ"s�RC_�P)iM徽�FP���8���5������dl)m���c���OZ9��n\�ɞ#�Y���DV+G`�ͩwTж
\�����Km����\VdLޤolD���9��W*{���+��b2���S�1��g������*2�e���˒G��鏥M��s�A�,ǙL�6�5ױ�o�������`�u�s��3\^8��D��x #xB�m��e`�� L[�����Ds3˲�嫫���X0��  z�����
�.=Pk4&��*ھ�'-jMe>�+ލ
f��v}q_�.CiL⢾uzȺ��������n��x������B)��p�mˢE]��fP)��B��
+A��J.��8��jVIeVՉ%'Yw�t�]L�LŊ��>�b�ቱ}N
骪(e4�)�vܪ�P�2���M6�ꩤ�����b��)��hhhj�(���Pj���.��M4�����R�P"")��M�۪��?{ɴ���;Ju>�3�ҩ��M�z��GnNd*Rߍ���f+/�Jp�QOuw��^�VP�9�L[y9�q��L�QMT�+Y�����葫d�6�A��y.����񾶪G�yo��T��R��A����TU9�V����Kp)��M�Ҋj#�  bH�c�p��ovh\��%#N�)Z�x�ͬ��5������P�'�.������$�3�Ht#�p�n\�4=����N���_�Vv/\�$P;�B.1 rs-��3�/�c�0�}]^1E�Ufe���1��1��=o��#��F���9Y��
��7�	]p��<�y��=��r��]�G���^ӧ'���s���D���7��$H���>�x��J���o��%茻G�HYf�W��2ci�J�R��3����^�<��3i��"2~\�ŕ��8�K�Y����ة��N'�6�����^��X-�{˔񲡽b��K^om�H򣡝^*��=�~�/qd��)^�[����25*��5c�fkh^*�����&�����ff&Na�&:k�<�=Ɔ���P���븺��G��N.�R<m��|��W��3��Î�R���C�^�����:��}��������uq�[g
t#�� ���:\�A�u�&�,y,���Sx.�"������ϣ�-���f�d��I�7)>��f&}��U:�ʍV�G��2>�#5e^X��L�u�
HWy�,{��ATkƩT�r�h�nKlx
W��s�(�����v��ۻ�.��k_ =�7��^ړ| ��l�S��PG��g�mȽͅ;� ��0���=�R�~PU�y�Gi 0U���)�x��;�h��8��x_�T�u��K�T�a���3��T�5�<��8�-��:ӎqO���,�����*	v���f���Jaˣ��/��Kߕ^n�5��@���_�;J�٨�5�痜�k�y}��|K�%��Tݾ�z$kF�s$��Z�"V��7{��1�R�yv�ojp# '��Sk��흲�8�`Ce4w]����0��g���e��a��f�y�w�a�vs���P���Öx�<L�C.1�s=��ąUNs�m[(�<�<��8�2�S�%�N��}�|�����a��j��!e�_+�Ѥ�Ka�:��<������V�u2��}V���Ǡ�1����X/=ٜ�c��ٍG"&�T�59����N�^ 0��A<�u=b���Pi�^�><*�VjlJ}3m��z�f�wF�YlO;�
C�n4����E���P�F�S[>��k׭��Ɋ����Za�C���ݝ����K�5F����ZNԭ�N���,�5�w�"�YWEo˞<M�i�t�2W�}�o��Sʕx�a^ܱ���PG�>5��'����WoNKܠ��߂�H��t���D0f������ I�TyG���v�f�ǃ�ڊ�`� �^F����ڦ����B�ͧ��L���8�M��{��1�6�Y�s1��k�q����p��Dx�8���5-�2���Tm��Ï*q-{�g)��7Tu--)�����v��'T���T��e��5}[�pz��=���
k
�mC�O}px�D�.�aO�+)�_�_W������:K���ص��pe�&��Ģ�+������9[����q��yg�p��;A��l�d�j����7.�7ғ��R[h��qT)Y�ҟJVs��ñq�%�3��n���U��Gn4���vđ�ع���܍�wW��1p	J�%5����Š���&�^�<`[{(E
��qKۍ��76�<�8�7|/���
�WLs��E����R�w`��\�@LWƅ����l}�˒�忸�y�NW
�"�(�K,-�Ĩ��g\
�������u�S��4d�A�����<�];��Y#"k�WbA|�ڝ�v�,�",E�
5T�^�*��(Q�VU�QF��QTR��TV��PE+E����U���Ji���"ň���)��T��� �(�ճ)^��˕�F/Z�љ���|J�?8.\+����S��4G�b�aۨ2�T���F���V�a��O
31����G%&���r��U�;k��̜>m۫�anՕ"��5��M'�1��'D�4�C͗�Y{��U�F:JE�e��C��s8�7˲���S�M������eX��!���>�v\M�$9YkI��nn]�	�a����mb2�|�(a©!�^;Y��=y��L������b����5P��qöi�z��ڳ��0�����&���r��4W�־��G�7�gz:�0�m:��x���汣�i�Un�ڜapz�>�N�:�t��/TC	�wY�y�#&W�i��u��w����(m��e6��Y�]�mV�TGğ��_�V�����Y�G/瞕zȑkNpק�ڛκ�.��l�30��ǝ���8.ӏVN]z��6Í��3M�����M�n�'��0ì��(ˇI���;�۴X,�1���6�M��M��µEGx䩑)�i�t�e�ט�2�0�<����Kg�$�|���rv������2�3������eow�^;�"7Sl2���NF[4�Ǘ��77T����Z`ަ{1-s�սD�ݮ쭬^�U���]�=;Q�л��7� �ת<�|t�v�9yLn�B�X���ݹ�w<����80�5�s�Y��Dӷ��Ц�FU�j���r�o��7\d�Z[Ǻ���)�q�jg^Y��9��:���$�x��I�\Ֆ#�
�;�h�M%�6�3X��Lav�ק������~:�l�D۹�K��!Ʈ�{����tt�d�C��3�r�/3 I8��n0%�K����8�����9���ORi
Km:����.�3Hi�5�-��.����޳hzCi���������5��Fe2'h�4q�e�������U1A�4>�
�8��k<t��h�m�dj�]��ݙ�|O:�;"݅������T���_n��놹Rq��k88�R/Y�P��x� ����ju3�[��<1��^֮��5��}g:�U�a!w;��fj%��)���i1�3t^}c/9xܜt�0�3ŏ1�a�]ه����fjm�;�`�x�&���`�[;�2f�b�٫<3�v�e��aI|���-/��a��L�̦�N�i��͏.���c�"��!C��Ķ�.5�U����=8,�Q��A8.����n�U���xQR��0U��/d�k�C�%�M��V�d�k�v�J��R�gu�ו�g(ύM&\4��}>k]@�R��i�����x�4�e'�t����_lDe��NC�ɑ�Ĝ$k�N!M$�-��V��g{:��8�P�F���u����-7��(�q��4�9�.u4��k56��i�&:��L���N�a:�[�b���(�FR�l�{�[����2�k��y!����1[���Ш��P��j� 	����cò8of�������Bݙ���)1��8�b�|댛��㝹��;�N��VcT�8��v�FS��WnP�H��i�p"����j�yT������Ztg^��o	0�(�g.��9�ec�������L�T0���9��SZ�L)+�{�֦�3���a�U������8�\zVj�W(��B@<�;�R�t,;}]����Lk�}Z߫nq-�*z�;�	��.�z�N��!�zL8N�r�ti1�w�'���f9��v����/�SĦ�r��Bٔ�Ѵ[g[p�1W�VZ�􆪌����Al�ܹ����m���Ѷ5R�Y{]ƆguPV(�T��a�N�ƹ��0âc�%�Wv��]_?8�[��ᦡ���zud�<oI�¶�=ğn>�W�^�;����;� ����',{`y�Bsn}QY�wR,��-���i6��[���Z��Ψ�L�\7�L�Ę~��u��Uu��!�i������x�Ѿ�S)�L!~T�1�ٶ�"������n�\N��g.�`���[���y���5gY��ŇY��e��N<��Ѻ��ܙaO�2>af��X>B�q�>5N����(^>�|�}��+-x��n�����a�K�;9h�a��-
k��.*���v�ͣw�HSn�[�\��ũ)Zt�}��>Ő�o9�!��e`ei.v��i��uscn0hޥe���/���1�L��Ԁ�h��6�gJ�w�YX���u+�*�¦*ˢ�Y�S8I54��c��=T�ր1��*>�WQЇO��+��f�Y[ͭ��]D
�1i����EY���C���"p�wwu��n�\v�I
,ؽ�x(i�ޫ!��� ���ӧĭP*� ;j�!��6����g(*q6ؾ6w��#�X��b�g����d�w���9�,�̦Tw����P�%Np���u�>�4{������e�TaS��R��� �
�YUJTX5D*��S\�wH�j��"��X�S)@��I��!I*��U�-,r��KdR
RSa
f*��<޹�u�<��E���
�mn�� ,��;��❄��:�ox�M�r��y����u�o|��F�;FSM��0�Zk�f^&7�4˺+TΦ_4���¦�S.ަ�hۦa��ˤ)�s�:��l�sU��Ja����dx�6a���r���_lλ���0���
-4�/�ۯ2V�Ve�����9�i��VF]d~���7j�ehk'%8P�fb-�5MC��v���>\p���n0+���E�v�[�H1o���v��.9�S�00&��O\#�c�S�mv�砋�����Y��*��p#��B�vV�lpf�c�pL4���b�)��gN������gP�����)�[�(�0&o��'����2�L��q���UP����5�h�T���+/�b�[���o��6� �\����i��Zyρ�0a����+)�W}%�꣄6��U�R�Ù���xz͊����gÖ`8Z�Ź%3��f�`��ם��\Yb�U8D:C2���Q��-ߢ�s�Yʶ.����/`���&��gTHO�Lkŉ��pm�ǀ;1�q�n��*^�$z<�_�1���!dC���������ݿ
ֽ�Eהb�[C��]��5��ڢ͡k�/qu=��/�^92�ٿqƬ��	LSTG�k��гv���ǌ�^��v�oJY&)�[N���*�|oQ/�+�|�}�^�s'e0w.�JI�o~��~���E�b�Y�����}*�v���)��/=ᾄ�tȆ���{9T����/���ZW�K͊�S�ƚ�=j�������+h�e��!�0{z`���������^ �=]��g{"��k�c�sg�;���ٯw�'+j�3�A2;Ҏ�{+�SEz�v���:u��ed�����(�|k��秱�o���l�j0��AzׄΝ��b`��z�T�JԤ�����. 0�]�U�^"i�e)�7�[��7�/�K���aՎ�մ��97G����~�ޫ�z��{<Z�Ֆ�z߱N>��b�+nG�S�,�������Og"Jޥ����c_-��������=�b�ïC��]�/<�SߢT���fSǬ��J��̧!Eq_5ץ����(�T���'����7YG>{��ɼc2�))W��ד�����ε�{� R�rF�{J5
gx��x�
��w5|+�R���2@�仑ks�	�К/#nW������@F�ca��ᅅB��j��°Bm����n-��T��j��yUb�6��׭�g���]<�D�TsE/xAy}vZ�!�Op&��Ry9����Y�<�m�*��3��_��,Itۣh�S��-�6P��ha(��]BG�υd��aGm^���\՚�j���8�-�E^�=]Vs��/{�����K9���R��k1+�������ݓ:w�y'솆��^^|)�?�Y��Hz�����SR��j��[�Bݔ��-������=Ŭ�m`�`F��b���G�Υ�d���5|ҵ�,���l.��O����M��E��Ё�5Sw+Wt<���|��Ȳ(�e��N���=�w8M��PR�sn�Fi����2�59r��L9�6stf��Wխ#��"�dո�	�KL�L]��
�ʲc)����1�iѦ�Ѭ'�1�ĀN�#Ei�ef���dJ��$���-�6��y���^1t@��Ԗ�B��r��Lys,J�%B�`�N6	�%����wIm�/3�Ab��l֩�SՕ�P��A���	N[*�	)�����SwV�,���),C	i�a�,�*[��d������-*Ub��^.�H�LRa�-�v�.��j���hUTSKX�m���1R�1��k�39jU��g{�8q�L+Z�;��NC�c�5�f&kcܖ�L�nl�mlzɞ��F���{ٴ|����p�o
`N��`��q�6l�;n��[h�1uʍ�5/ݣ��]]�����Ҽ���+6�J����oÓ��en��S���0 j�s��4v�/R��;�f�ًux���v�����ܶ�1+�&4�β��ϙ5���yWXZ�:t�q�Š�*���Z��y�6��V�{inE[�ު�E�q�#����'} ��qY��Ww�In?��w�F���z�)u+��[:��?vx9���cޕs��u����(��z�]���������ި�^�X���ۻ7��lh��J^:��@il��Bp��Qf;E��!:�3�{:�K�N>��.�w��N��>�=����Òf=,�~w|xՇB2U_���U_���=O����l~)�&Q��t��1\�QR�����{p����svQݩ�c�p^�7.��`��{<�����ˡ�(�6[E\�d)>���������6���H��������nhcֿ*-�v:g�Ik�<�G����u�g���-�)��׶�������sB��z�Nw��rn�����շ�W�D�5L3�l�9��}�c�to�k[��s�eP��bZ��]��EK�$�ԼI���!�g�q�����ztzV3~˿j)sv3�/���I=�K�7�3S�,�xtJ�Z���-�o/�]�rڵ�����B��IoT���Y��ʗƖ r��42�K�Bf�Õ�#��8���D�G:_u��t���dO,�&�y��\��ρyb��K�gǠ�oE���^�>:���F�,^^|VE���>��w��T�������ѣ�W���՘_v��+޿xCf��q�q���e��ܝ���9�;#�rX]R��[K� %ꛢ��*iʹ.3lϕ��LΓ"$�� �^|��2b�l��p��9�꾂b�+ �z�/ls�U��P.���D=��X �Aj�ٗ��`�L��e�xz��왻 �KƑ�l5��k�;��rk��'�߫r��p�Yj�n�h]e��[:7a����T���ץ>E�E��&�+ܩx�C�z��A����?c�'�h]7�>� ւ,�0���^��.�<BV�6��nS7�����Pw]����d��ڄK���ǵ-��<�]�է���V��s��`�W�u�z�CuA^��C��{2P�V��/gf��u�6�����Ũ��$���6�<O��%�%����!�$�#8�8���<|F��f�
����q6�]��w�����(K�-\���6�Ò�hC�b���A�1"�U��t�Z�V��θΥw�ĵl@�5��������"��d�9y��x[��uy�Gr)HQ$l�+�)W]�\l��k��K�j�d_��c�
���o���>��,fY�+Xy��a]��g䰐�a8�By�2�D��e�����d^R���mK���V]�0�J���&$\�X�@�t�P"�h�,�2�`�@b]%Af�����L���K<N�E���h�$��Z@�wWtFe=�H`_��Wrb̦������0�k.���gc[/�Ɛ(j��R-r�T�JyKM]�KT7E��M�kPh�*��e�YX��즩�����J�F��-�t�]]��آ*�0��lb
�B��P��*Z�4�h�b�DV�V��qBҫU��E+*��}`�5fv�իd��(��Q��{��`��SQ��d��e�HN��eQt���v�d�+<���"���j�1�v�u-����tlo۫Ô��\k�(v陓�ǯ�B-�r[��/�������䧪=�����#ٺ��Aܖ�]�N�݀FxmX�����9�^q�!�
#ȋ��Ą�w�`f�Tv֫�:�3��oݼ�R�N�f�����9���]�'��v�3��2�6�؝=��Н��=�2X�_:|�b�Y�O�Mэ��lg�k-l���3w��n�x"�(���aͭ�[�s�dakG��[7��!\D��n�Y͑���㣐��l
�6����xp�fwtP�i�;��!�;3�v�r����_
xY���gM�=s!FG������%�ղN�9u�݀B;mʙ̆�H<lv����e�ξ\k�K�Ж�d������T��r��¼�h�b�-�&S������7����ю�۵��Xn26�i-^9�ok�7��h�m��XΟC�<+M�m���ez�B��O¤B�l�sF�2��9�ћ���{�S}�>=o�m���ҴC��D��䬏
~���OE%��"�<��{�����٫ n�4z�sݚ�Btt����m)3L��C}Q���t!s}ˠ��ܣ��z@��,M����|UI��+�V�P趒�jc����w&A#��(��3R�w7�wP?%�/�:�v�����꘻�D�5�`��[�_f^��X�k��wX���8�5���#~�W�-@A�t箻o2�qH��.5%���/۩Y�,�xߺ��nBŪ�$9]��C��q��JN�ɽ����o�ͯ@N�N����j�j�ȴ�ط�j١gN���Wq��'�s7����5_#�_6&�}�����!��s�k�C^FcZ�{j�u�T2�=g4P��拖=�<b��x�B�f��:�o�-���k��-O�Ro"q�83kX��;�l����7m�w����ʼ��W� �Z����Ӥ7Y۾�P�����y���mL��4cک�S[�-�Z��E?V�\�͉X�o��O��M��v�F�ӮY�*�9�1w=�E��u�g���������6������(U�����#�9�UAѱ*Ż��P���j3�B�s�+/f��֧���v��ǥv�{�����Y�:><�E�����U�SpkN(��eRw@�Yy�1�OT봬v�b	څ��B����%�X�V�wk�T{<0��n�~��R-���U���>y�H:�Y�����>ߓ6����V�+˳d�?6�3��B�32�O?jbj{no����Uya�<P�`���X�P#� �b���w�������^Sַq���	�GO�xN;��"W;@"�2�1`��\�7{�ӌ����4��ת�7����|/4�(�+z2MRC(XB�%r��m�$	�k��;Y����BXx
"�XN��vm]Ӱ;��6���5�^���^=Q8���ۻ�V율�f�M��X��[����g)+8!�c*�IP�iIi�WyP,R'faQ��P� ��� aBm�],q��.�ːW��T�R�ʹb�	�蛹9���GT00����[^^9�y,�ee�믅PPQ�P���ŗT��j5L���QbRJX��U��Iww(VRP�Ei��D[J*U"SQ��Z��)3���E����aIJ�e�E�EU5)���P*�f����E��*��N(��,�F,+����<�x�;��Fl�V���j�n2�-��ыkKɷ�u.��t�~�T0^"����M3#����yR�o.�Z=喠��ʊ�o��J���9���K�N�x��%�e�UL���Y�s�r��i~��ÂW�\; ^WIӪ�]�l˪�������YIӔL»o�0�i|�²>��n4�&�`�`K�n*�9��������X���0���2̑�X^�U���}�I�rSaW�e��`�*P���<��� ���{Q�nv�`qv^;EoQܔ�lj��_��υ��b)�}��/Sh؇�u���Ka�yǹ���ב����E��"W���.{��YE7�t�I&����=U4Fj���q�c��FZ>x���-H�sW�ej&"/�{�Wt����bb�`�A�\�.ʛΥ`�;:��' ����w����׹�Ef!ஷG.R�59�ne>���d~�� �٦_���Z�} /v��
ge�<��<���՚�̍|ϺY��Oh����F]jyz�Wݏ���ϰ�@���0 ��h}�ê^�nG]�@�H6!��z#fz���g�vy��qdQ�C<ڱ�,����~K��u_�66$��+�ǌ Me�̊^-Q�hw�5��NB6��[s/4����,u��4�]bQ��<:�F�Wp��G!�N|���]�t�*�.��Э����"��ËZe��=�,K�xf�{����jDX�]B�>�J�te�ٲ�n+�B�Z����d�[��{���7�ߕ,�u�xmZ��;FX���t�o��	ߧ�T��ȞU�,�.'/�B�p��ѰeA\Fo�%�9uz[9J� ����[9���X����tv�˓�4��p��2�ǔU��n��Vbۮ�^�&�h�x�q鮲XZ��]�S���V��/f����P@�}�Ҟ�fl���K^��̜+6wRθ���>ݞ��6
��iQ;渫-5�ՙ9(�<��/I=����������u��Y�A�s(̣ zEB�cG�'���)��q��/P|���[��ꔉn2r������x���|rz?{W���~�@��I8 ^��c��5�~�_��'�~6&�Wz�A�.l�`y20��e��W�,�	j���P�Gl��ݓ����wd�(�]��w�2� }���q�� A�͙�g��Wqp�6��������a�k
�ռ)qa۔��IN�; �v^zE �u�v9b�]v�><�Oj��/;hf�l�H����؂H+��л�F/A�z���I[/�U�ܕdc�`Hzr��YB�+�.$��Å�;�����]kO,УE���mǑ¥�_f�=�;VЍh�[��](���:�Z�kys[Y:�7�&N�*�]a=]@��e ���j���;̔l�QLٚ��i�rx�QC��+��!���g͈�N5a�}s�\���x�\����d8A��l�p�k9&4*�[���r�a�剝΂�mv��8*�n2�c��ȉ%�1�`���P�7k ��>�,���hWQz�R��!�8C1�V���w�;q�Xh|b��2�2�I�.U�ZTE�P;���ptro���\Բ�*Uǆ��K��d��:��]�}�i��a�vJ�.s ��qN7�c�L�
<�[�9_\�p���Ww�YaQ��2���(�AW(R
��T�U*�cUBҴ""�R��)B�X��V��H&%��-.!N%��[J��R�b�Xa�+7.�e�D�JmX��@
 $�4E2Ss����+_w��Y}֛�̕�w�t*�ҨP��xN��(z�u�Ɉ��l_]zMiob0�ZѴ�������eaͭ����ǶUꞸ����쵓���֮b˫ٯ%�R�ʶ^5Ұ���K<��Xy\��:�5{����H��>�*g��X(���7,�Vr_�x��E?Z���擹��*�\*}�x�k�]!o ��u��
�G��H�d�}���=�}{=�6��݃ϒ0��Y�ѯ?V_�*<������b��Ч�hz-�<)u��n����w��4������W�ʞ�C��6��TT�{�{3�Q�q�~�Lu��ͦwL��Jby�kW�����Os7<2����_�Ċ��e�gf����<�\�e�W�A��?<\9+�LW�EX�|6���~<W��l�{�Z�5�.ws #;Xv��8��{�َr³'��M#k�KҐ��-|�In�ߧ5gxWe߲�>�e��֦x&q+*ɣʅC������_�nN�fs��a[@U�{���@�Ӻ�{��͌+�1ت#��Uɺd�����wvgo�J�˲h�gg��d��kc�n?tYB��P�G|!��E�S(�uP|Y�f�úD�!�a��7)x�~m]Խ��.m���S<m"��3fz�.6�>ͺL�3&�d��`)`Ͳ|o	�~S_I}6��=A�r�-\W���گl�y�M�ڍ�/-Q�D����j]C.�t����sF.Rk��ɾܨ�	<}]������;�DPĳT��ֵ�^�����&J�i%YPo�N�C8p�{cwl��G&C-;#����}��,��39����tK��QS7xӃ=��v������y:�l^V���F�G�--^Fߔ=�R`��ɹ�����N���]���LV��8�G���T`��5f�J����/�7�q�˯���^8�����/la��/���bK� pi�}���8�������GM�L�cb]��0��������h�u	��[��i� .��'��=�/�g��>N��W1
7ʼ���o�`�f��ߢ�C1�}w�K�������q��G�ЬSɠer����pR�����;��#�\��[�e�BqPӛYN�]�Ð=��c���]�*��@�3���𲯧n����s2��Mk��gy�����8Q�N��+|/R}��I���XqF�^-�[tf���)	�g���n��契���+�����{fN��Oyo wn�_��&.lvv]#��e��{J.M<�|��i�]Qm�Al��f��֗�;�b��M�N�^G�j���ma�OxNa����ؼv�b�K�p E���/������?�?��� ���~�Ҫ��0�� [G��  ~_�*t  ����.��*�+J�{8Q�?���:1�|����wf6Y�2G1���=��c��Oc1�m�d3*J���/�T�I$'�$_ky_���������������g?,�)x��C�p@q�i��g�fr$p-��   �����>}�c����@l�\  I���D '���aRY�����ʃ��'��'��%��͇��ϼ����� h��  N@?:��>�����I��,!��X���(���z`����I_�W�z����'އ����8�q��j&��bO��  H�/�c�^���#� LOŰ�0@�r�!��+^��%]���&��f�A��z?  Od�4�_#_|>?�c�?��b���`=�ԇ����I?���}�����?�����ʏg�� &~�Sʍ���n�������K4b��Ov�s�(
�	����������X���L�������d����?#�M���  I�P�|�/��?��=��939b���j�Ϫ�� @	3�p '��8��������Y1����6d(!��?i���$���U��叾��G	�w$ �ɒ��bI�>A��1��_�A��IPO��3�\j��l*�ݙɎXPq� 'e���>���'�  G����A�O��ɇ�w������{ �'��?��'�����b��O���\�O��}ޖ�����|/��}�����  }�>���/�
���?���P %I�d5�ǒ���!��z?�>��{�� �{C��~CY��h��G�������o�_?jL�D���������_����nw�����ې O��>FC�`o��~���j��P���o�'О��7�j�<2$����'��=� $���~dO|	�9��3�7�����'�O����4�h>������R�������ɨ{DP�H'�(�������rE8P�'٤