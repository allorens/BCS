BZh91AY&SY9�~^~ߔpyg����߰����  aP~X �I)     @ �    @UEJ
��@ �HP     %@��@  ��J�T4YRFE�%kl��N��@π �Ԑ��
�  �����U���M=��v����C�힁�;c�ˮ�\��<��;5��  �9�A�:��<�:  4�5�D����8 {c�A� �h    �	���G �kA펝N��H�+�fQ<��;�)s��xs�ƻ��  .����Kݸ�9�A���rq�=���{��z�g�����we8�ָ� \��g\ 9��]�j�s��ؕh�����{
�nX��N�����/�x�2��4 / F���uѓ��bȭ��=Ͷr�{������/]������ˣ���  3� ����u;Wn���;�D{ǵݑVq��l��wk�!�׳�n�WN �n.���{�{����r�r7u�^���t�S����ҹ�˛�c���  
��`D=��s����3v9Y�����:=n�v7f���z:v�֋��l�{Ǽ �;k��]�ͧSs�=�\�wM��W�\�֪v��zOY̽k�#�����           *                ��A��*R���`L�0M4�di���DI*��# �h0M0 	��'�T�)  h      �H"j�$0�	�`� 0CL�&JDɈ&L�4���mM'��F�2z�������i��*�0 LL � F�A�m���$�	��	�lq:���-�b���Y�cؠ��^( "<� *��b*"��YP�z{�������\!��ȩ>P�$�� ��`E-`y!_�J��MW���pa���&AUUU��) 0�[:>޳��i:��������?�t�����M"#�"5V�����B'�'
viĹ<d�b"#�����8���,DN""`��DD���D؛6Z""&�ҁW�h��b%�"Y�6v�&"P��$1:"&��DY�""Z$f�P����"`���D��w:"t��A0Â;��"r�"'DYbX��N��#�<"#����5�ob"xy<Q�:'��"tF�J�DL�pDL:s�"a�Ȉ��dG"""r�"">��$�K'���Kg��D��#H�>�"#���n��M�t��'DN�D����&��h�"��G^�t��Fީ4��&"$) ��"Z.��F�H��O#n"#q�QMDR-��8�����"ND�:b"&��"A�#�x��|�;b	�b��"Ԉ�F޴�GѤi�[��Z8�F�N�>|�8����(L���Ĝ"#H�\DG���Fքok*"-6�Giȋu��""y,�f��""t���R`�DL�"&	���� �^�"":��N"%��<�M�8"'8lDN3��tuؖ&�v"&��DKg�R�""'9�V�<�
��a�� ��"UDDM�=�"&""A<ΗE�DJ�O	�"WA=�<a�'%D��""&��Dؖ��b4L ��D�	O	,�����c�DDO$-�d�O"%"""s�X�X�����6:���76"p���"&�h�"74�0�J:"&��"t��X�͈��M�LDD�6�`��:�B"R$D�%<&���8"<�DL�M������Ȉ�"N���D��""&�	�2""sL�"'�D�DD�<X�����0��b"p��8p����#����"#���'`�&	�7bQ�_�l�MNUHsE70w6a��sT<�M��_�6K���#�ӣ�B,���DD� ""9 ���˔""X�'�e���j!b"}�����"&�pDK6>�B"lr"&ą<P��'O	�Ʌ���O�#�8"%�� ""9���&���,j"X���'��9� ꄽ�E�,��#q<'��#s���&�6tFJ(舉�OO!Y��DJȈ��;r�JDK6"#q��_��d�DѰ�!'��ݙٱ0}!�p�Ȉ��K���N�(K��6�-������g
(�YDɂ`���᳼0Y��MBnA%��*�`��i����0���'K��DG��2��",�C��q��0��z�	bVDٜ�"y<�i�ʹ�x����F��mţ��Du��GQ�-��Z4J�g�<8p�����{ ���t��ؐ�8';:&	^�x���G��:I6t��""%�a��pF�d�#Q0������A�"#��=� �Ȉ�͔"58A��P����Nb%	�!��'DrtDM��(yg
Ȉ�>����ڇ�0�	4����J� �7p�����bpIQň���"'��p�C6"m<P�����
8��`��DM���DL0�DDM���:���B:���m"9uh�1��c�1�����m����DDzM�<P�67��"<���l��AȈ��DG��K����DK�DJ6:�0D�OzP�t��DDD�"7<2tDK�DL82"""�""9��"#؉�Iu�E�Yb#��"'I��@�""l���b"P����Ȟ<x��D�d�^��lD���"%T舉��D��"""w�(K%�DDO1(L�D��K:'j"x�;�!l�,D��'�dd0DNr%9�ӧ;:c �DN2 �Y�nA�Jd<aB\�K��8&B�����pD�bQ�N	���0��D�Se�^͉�&O,M�Oe"x�lJ8P�G�ř�x�����b$M�����,D�""#����9�e\�"'�DLc������xD��qbnM���K�WbM�2�iÛ����䴣�3ǰN��r�����<N����8�~&�bM�M�&B�Ôsbu(�$0�(�Ht����
�6=��f��D�A�P�qɃ�
�M�0�npOT��X�9��7Ȟ�㇋:t�8"sfP"&i<'��	iÆ͉��e��R׮!�Q���J�h�pr&'`�<&naE�%��&� �ؐK8͖a��	�>���䇁*�Qe�'x&�',�8Q��DD}�`���H'L� �����͏�Q�7Se���p؜vġ�:X�g�0��"#ؔ"X�(HB�""t{��G�	�&2���'w��pL<%�t�7�t�;"'�<:�K,K�2L�:A2M""&��"&�b"lM�DA|�D�!��""l�K&DDL��lD���0M��ț(Dt���"pْ"%��0�����:P��bpM��i:"#�N�+�M�"'�<�Y��H�#��:�T��qDm<��B%y ���7��	�b{e���	6""{b	bX�R"&��ZAK8:��D�g�:'D���������<�bX�gJ�&:":DN��,K�A,DD�A�Z""'И""&�"%��n"#n�u<���q�6��"X����:"x��P��c��j>�H�#֢#���d,��bY�:����77�un�z�ն�>E"6�ZGl�HDSqM7��+��z��q�Du�#�筴�mZ�=BQ�!�a�}:V�ӂ{f�Q�QƎ���}6�w�|��u�b&�wPެI�����<rӉvp9��,啢�^���LÉ��Ƹ��<ۍ.6���m�mF��8$N"lN�ؗ��noI�Ŧ,FDD�;,t����� �DD��"x�B�&FM76e-8<�`�a�f��:t¬؉f�'D�D��I�:pHY|��|��Ω��D{��&ıd0Dji:&Ӧ	�l��al�`ɮ#�G�6:f0���؈�D��D�����D�f͛8�+ӥ9�؝0t��D�7�t��p���%	�rp�w6&��c����,�{��`�a���<>�6^�$����Of����_�>�v�W�5��Qrj��w%)=7��&��kك��gaE��p���A3�g�gN����>yb����W.Os|�����qy��9ޕ]��:V5�n�#0�k�}��s��C���3�k�ۓ���>�OG�:��d����O�͆����#��t�'9;v��4�� ��{���s���~>����{۔�ɾ�<�������{X3�g%������=���e�$�Rs��*m�쥒�.��h���F����y|x��>=���ϰ�����'	�_=�-Y\�n���ؼ� ���|ۑ`w�^�����٩�~sή�ٿt~���߯m=��5��f߻�w+�8�jˉ�ӥ�u���~��͛���.f�U��9�m����Љ|��ާ��g���Ӷ>�����������h?;$F@��������9�Ϲ��C9��rY�ݷ�ٗ�����O3n����_�~��y�f�����MϬ>�L�q�=�f�M����s��}.����w��껞�ON����d��FT��Sڻ���y\�s3����ﹻ�_[�����Y����{O�����K$�%�ެn\�~���d�g||<�F��������g�����Sɸ<DҼNI�K����b�lƋ�g^�)Sn���P���ّ;������'���k�����/��7z��K�*�7Ǔ}�;�s۫�e�˴�I����o��w�rC�w�}�ǞB�g�;��5E���Fh��XI"t����}2�f�3��Nϑ�&�3�]3*�\Tƭ-'vv�a�&�����C��gV]�ﭻ�j^������f��OzQ�5k�py3�g�����f�f��qo����]�lx�={���r��;���m�9�YϾ������Gܗ/'��no����ޞ<�����~0��L�>�g�q�~.{O{a� �����2����Y�f|J�)9+��O�o��{��:}}�ی�=�[=�nM�u=2'�v�Sl熵^���9R�t��U�O]�7��px����6D���U�o{;:W;��}�P�s��|�Bow0����竾�T�\�No��ˮ&�g�5~|�g��3"�zM�2�J��4̒L�|�{|pK��3vU�笚L�Eͧg�>{ڽ��37�t3S:�K�&���,�0���{JL��$�{�Bz*��zN͗%h��ߞWyww7�2�s�;��3w�Fo��ߦ	'��%>�����|t�� t�wػ��~�ᛲ���Ov�?}!��|EZ�}������^y��p�z+��"�Ѿn{(�q��s6�϶[��{�_��N�G�Hf}ߣ���=��%�=���]�k���~˯�[/�����溇��-ɧ���{�:����v�oݳ�o�Ӈ�Ϧ۽,��gg�v�M��x]S-)^����9�����2{=����r���	��=�z|r|�� e�}�i��C;̞��nnn�9�v��;�{Ē�74Wl����ꢴNP��;r�|�s:��>�ڝT�'�6J�����	t��[ ���_�4�ҭ2R�0s��;|%O���w����9=:e�=�Ʊ��b>�rw���U�҉S�g���ߞ�4�x�6�%�f|��ӝó(���g}߰0]�{�]�1�s�f����*�N9�.�ߦs�ߦf~#V��w�b�K�O���f�t�۽�3�3^��}��w�;���f�g=m���Q�r/f�Ny�y�xy�=g;g��KrM���Xwp��=���	
q��L�ә�XQ�0�B|q��X	��{�,��M:���Nv�Z��'���K���ﻝ7~��;��鯘m��rn�Ё1x�D�__�v��f'��Ff{�����eojy�G���}����9ȷ��=�t˔7�|x��9��r�M�L��v*.��3�O���c8�������{�\ʻSRgƒ��c��c��w�����<�?"�x凍��ͲI҅�����s��7{;0��}٘���hY;��V>��>���{/p~̟��)��3>i��:�ʭ%���>���0��/����ͬ�;d˓⛐����*�a6)@�Y��ɞٽ�ǒ|nl\��Ʌ1{~�f�g���(�债���� ��}�=p$��v�%����S���7����zl�����h���Z�Q�<*��!���2|dN��ǋh��,�lݲf"t�e{����Q���JN����L�	�o�5��vߍ�'�Ǧ�!���?�׳��d�x�d��g���a��܆.������>����g�2m�]"���O���8S�:z�f�:i�Lp"y3몿������!�Ɵgӫ����=�:%��k���w����)��]�O�E�k���g��xy73�藌��e����fy:��;��I�Ûgggq]��i���=��m>Q�f��\����o�{>!�����=;��'&�[9����Ese��Ι��rOn�|��~�|U���+�\���&|ǳ����ӥ�w���.��sL��͈��=�^�7��_�t�yy^{���;�����|�/۳W����}�/���{�֞8fG�)�:\�����7��?�s�tsd/ �)F��L��I����w'�7_6�3>�јN�2�掏�v�ǆ�3cZ��9�G�Ůw����@�����j'��������g�w1`�7�?_g���2ϋ�-GӺ���!�V֫��/l��y]���[Ν�=�����Zd�_e{;�&YCϲҝ������>���ϧҬ��_?�=+>vwd
gK�}~�Vl����L���=}>����~��{.H}C�۷�u��{W��z�o��'~��|3@�w3rO{73����~��޽�azUfl̍�Nf�U��Խ>�7�q�zz�BK=���5S������+�|x$�Nd���ƺ�0$�:z��W׳���t�������x��.6�� ��x�դ
e�b����ܧ_ѩ����.E����N�M�]�];}c<x�|[������s��!�ַ7��ۼv�{�.�>���y����(�~ɤ���3;!��xȞ��N�A�v`��$�;�Ґ�d���\�όY�����̔��:�u���{ع��6����n5�gǳ�]>��ҡ�y�.d᝘Y#����l����t3$��jV���7��>�;d�?�.X�;�٘1؝xg���9�����~J�YY��/�/{����gf�H�.W�ɮ[3����x�rQ�t�-��~���_���N�OO~����G�K��.��?d;��d���`�6��,�O33G,�=��5��8���E����}x�;EWh��
�N�<Q�z3N=�zΧ�]۟5��k����٫���H�����2�'}7v���di����?����/�^�������g^H�?�o~�m�]�!��Jg���Ϗ�gޑ��Qכ�"��$��]c&���-����{v���29��x����$����9��e�m�}!��=���w�_��	���r]��h���s�	�F.�{���wӳӻ��Ɗu�S?g;����Ϥ�]�����|兞w������~�����t�;��&I���=��7�DK���Ǿ��s����r|q=��|w������K��}����ϵ^N�>�����zu�<~���0�����2�fl/g���7�]�s���Hͽ֥������;ݜݭj��U��Xw}uף����[����e�+6��vQˇl~�:����|�}��m9�m��wy�}����f��:���3�k��;S]#�Z�ٸ-��Wx/�b� �٘7Z�d�+��|�v,���o�rS;������_�s&va�?dW^���w����;�bpϧs���%����{ࣞ�X�9rc�{{�ك߻��|.�t�E1�l������]���S�?�3���y�$�F.�~���ڤ�{���T�ǷM�x����s�Mo_���<�*�����cY��̓;%����U�c���n�,c/���rN���3]�\�\�8n��e]�#/r�s������������Rǔ%��,��V�!!�ܛ��
�}B��H�ȋD�G��g�8��F��W$��-]�ۃ)�p��\mnݭE��.�N�n��N���/�^��cdr9C. 1 �	tu��@�.�7ݾ��Sǽݿ~����y;���r70:NE��#2,TqZ6��e��Y�[��:���n[S���	�Y���g�JV�4�8�(�p��,j�4�QHA#Q�l�=��e�mv��X��ԁ�˳z�����v��[�Yz���d� ��n/�k��R��DQR��$8��c���gps�c��pkzp@�K�qƨ�)�ӸǺմ�E�f�w<`9��Q1ӇeŶzB9�:���Du�6��f� �q�Z{
��� ��$C�s���}��Re���CJd���$��*�U7?g3���ʮ�p5�Z�3�d�{��VE脓�����^��UN�&p��v����gYs�P1�l�9o(�`sn�:��`ߑ�z��{�k�S\ZHz�=,���ݶ��Љ�gx��ۚ��6ފ���0��+B�9t�H7]�,�Z�����7Bc"y�E��6s��]q�i<\����Ɠ��JJ.�E�C�֩�@�Ud	Ŀ�j���T���Ҽj�p�q�Цn��1�m̯�z��:�v��:i�V���qQ�y��v��wu=����}zW�޸7�8��.��۶�8)N3ݳ�n7g�Z��؊ָ�u�kQÌ����GEȧ$��`1@+�\�]X4���]��P"fIXY/�S��6L��Վ1�qڏM�먣lK����bq�8a+-|�\PKe�U#��Q\�����b��x��n�3)��w!�n�����m���}�����2� 7�hƘ�����B\ד,�F�jQ6��B�B���U G8�!%H��m�UV�Պ1��J�۬��� ��#�{�9�Dt�L�kM0��A����4���18�,jژ	Tc��+PI�:�$u��B2�T��P�!T��T\eU��d��-Ul�s.]jb���z9#�꣯=>8��tq!I����焢S�o�� �pm�ƚ�pb������f|Q���\d���1!P����L������u��������mM����v��֮$���y��O��XGPr������Go%c
F�k�ʵg�����;n����on�Q��9m��)U��9�ģ������MR��0����l�1���BU�k��A|X�:ekd*p/`�V=���7��w�����ysE1��s%CiE�X!ġʜP�����$�|**~��g�YߢմS(�D�QJ�N2�����e���������V�K�Mv��M4׳$ֿq��@�S���I�m�~|M�L�B"@dA�A�VDGqZH�0�
I"* ��o�^��������\U]�⴪�V*��EUUEUUEUUEUUEUW�UU|�U^�*���ڭ��dUb���UUQUU�=���W]�ڪ�b���UW�J��kA&� 5� n��Ȍ��7DUiR0	d@$$UkJ*+$�d�0

�z�/��}�⪪���ZU]�⫊�եUz�*��F�W����V�U괪�V*��U_1Uv���n�\Uv�j��W\��|�U^�*��qU�j��Ҫ�X��p��&��5�I�� B"��D���b@ԁ� �W�}�o�|��i⴪�QUU�Uz����Uڮ*��mU^+j��m���\UqUڭ��*��j��Uz���եU^���͢������*��iU�Wj��h���6�IYbR�� *�,(�=ed"������X�"�%IFT*1�U�2�UADTX&0��q��#�5��Dbz��6l�� (��>?߇��g�X����C��8%Nc##"�)����#h��Q���-DqǨG���q�>|��">DF��DZ">DG�"4����Gu�DG΢��E�!���=D|��-|��ԄiHDR"8��"4����"#�DF�i����m�"4�"#ׯQ�֎�����DihґE�F��z��B"��z��ۈ�Z"8�8�u�DDGQũ�q�|�"�DF�Dq�R"="6���"ޭ��q��z�<�E#H��Du���Kױ��i.���]��Z^��Kax�`��Zu&��b�C�Dc+����@�UO�b/>�޶9n��]�g}�|�J����A�vߢ��?nq���@'Ea��YuZ5,US�N	�����5��G'ď��}:��pq�8V�����).4x�1]x}ع�Ku�A�;����{lz��6Վ[OC�H��k`�2fw[r%���pqg�[�d�n����=���y]���R�=X�lv'v�%�݅�%�:la��M�x�砗�N]�����<:�9D���jV�9d�"��[SB�i��1�j�q�*+����v����g�˝��c�ܮ!TX��� A/'D��!oYeq]�E6۪#^.%1����]�Zu���[OiBL<�kt�</��F۝�bIۮ^3�8�=�����c[m�3�)��<��v��GN����\��:����������v*�|a6َp��u����/"9N�`������v��d���1ǞV�[���e��S	��KY��c��9�2��.<'2��=�bi�Og�ݶ'V2������x���� yˆ�x7O���+;n;<��38�{vW,�[�ݻt�v˄l��aYƙۭ���շ�U�1pG<�ofu�?W����:�����k[��!\�(�GD�����>�fSQٽ��zz���5p�r�������:�c���(ve.;SU�Y	H�	业s���\�ݬ��|}|��\��q92 �`�+���1E�P�ro�Wj����! �Q����Y���<d��tu��BGk�1;v���Sq��=v5e���r�y�ɒ�Ef�%ש8m��c��&��쭻\�:7qX�"���8{Thp܎P�����sí�� ���`�f��'~z���y�D��۲p�U�'���	���c�;�����Bu�a�0(���P���/�����6�{Zri��͎������`�n�w ��\�x���̹�l��aH�:��f��|�n<mm�a{38�y�u����얌�u�e��g���WwS���sj���5{Fn��7=��e���ԣv�3�{1��\[[��r��v�	E1�����\���Ç�k���.��Z��l�<��y��n��z�v���lܽ��ڹ�����wB�ݭ�U���L�nz�t�T��q	�b���g��s���z��Ŧ�v�����9�m9��8밅5�(�װ�����j^�<�u;o��4ݍmu�s|���2\�ʺk��/I��l��[�u������Yre�]�ƍk@��oX�����w[��x��y�ٙ�̬�$�w��n������fgs+2I$��}���<<8������1�R:�>Du�Q�f�0���˞�?M�i֍5�du8�D�ܢEq��5Ŷ�Vtä�G`�n/6M�y��T#�hLn!@M��b�P��F۞B̈́{g��m�^Sh��g9̨H!�������9�nw*���r��|.���_��g��9�Q�L�bMr��[d,<��V4�+i�q;v�<�u9��M�we�Q�?/�����ݢ�Z�5�GJ��S�nܖ2v.x��'F­�f�]ӏv8�q�QF�"��4�,geX\�ހs�4���v!��E�v��6��I�]k1\�m���U3���7w��w;w��rz���~ᾤ7,�L�14h�)��`�S�g:h��6L5���?�����ԝ�{\>>09�r�p�a삤��u+m�5(��aᇃ3Vt��q��K�̻���B����E���N4'���ƣ������ ��e,F2�˘�kb:Xi�}�VF�`�m1�F: `��u�C��ț�{�Tn6�5��b母�����껭��շ�O��b#q�E#���GQE>R�z�٭*��eޭ,���9���'e��r��.���9�}��;�K�O[�4�������l+ɿˊ��G;ޱ6͌n�y�:���"t�$?0�C~w��>SK��q�p*���������Yn~�w�.y��{�nS��8M�3H�NMI��`_6�6h�S�B%<<"'�:pDA<xN�:z'M�0�E��d�2��UCR�ٹd������2J�Q1Y��1&�P�T���}T�B��xny)����J�/��p�V�~/����a�����)C�w�yff&�e��>r&�Ю��=�u#���*���BQ
!o��'<pD޵z��앇�J8��ՆOL�B��~�ö8P�F�=(~�xd<8P�'L,����ԛ#~Z������<=TUښq�6���"!u":���)��TQT-�<�� Kʨ�\^�Mm�fj�U�ÇC�Á���J0h������Ge��,m��ɠ�3�w�s�t�ӆ����||�Op���f�g=MU����ӆ�G�f�Y=)gby�=��̸�[p�]�hKA���*�Ԁ��p�gN�=���x�*˰�Y��O��)�CC�aUD���R��L�{箭�}:����q����DG��m�M*��}ER�̎V�R�J��;n:eB��,O���Ǖ�J���3n��G�k�l���1�(X�Gܻ�Dc�X�ꑆ�9Eh�,��e�K�=/ NC"P��6���ם���P!E�Y�f�2���֛�E�֏�kEw �W���1OO�y���t��8��HL,y�"�dc��]^��n�j�z���nRV��.L�WWT�z>�6l�S�Pb��U;6I�ၞ;�*%���\��P�C���9.�=�́���n�N_���O)=��,�a����v$�$?͌��xt'����b�3��̩�<��'�`s��!����,�
>3�Iw�
�NR:��%U��M���/˻�S����r��3kM�4&�E�i���������&�6rӇM="8��D#���GQG�f�0Ѳ��=f$�H,ImY�8����<�ӓ�������k���-��~?�<)Ҕ6=���O���;6R�18�'��:p�l0?2SGM�.�~h��y(�=��b&i|��8ّ�|AZG��rW/hs�d��]Ra�W	��>;g����"`rk�:���h]q�ɰܢ!刧�9�|���\�c[����SҚm�\q�"")�Q��xD�(!�,��D�7��u�*���)����4Od���u�+!�� Rx=�ᐣ'�:l�[k��4Vl�����o�T����	'�@�T-������T�� �>�9kS5�ƺ��&�Rb���	p���Bx�8~2M��������^�\�~6lJ&_-�C�����<���
����j�>b��i��Z�ߝ�z�|��8��DE:�>DuDqf�0�{�ٕڪ�u��5)����32�3SV@��{�,��7�a���p�{�Um��̫���(��'Ayl�a�1Yv����q�ɔ�P����SS\ц�:ә.����x\'��[J�Ar`�Z��N+�����?NƛG'�	�x6?7����P�B�p����g����(�j~<ٲ�����(�2��IϤJÎ����æ�QG�U/�ck���<�[G�q��DGV�>Duu󭬧�Zi�=k����*m�W���v�鋟��f�Dm��:��RX���Li��	4Է�h�X��f�V�4�S�m�[t�HC����$"�" lm�K� K���6A�h��׽��<��O[
�<��şG'�]�zF�3�&V'ﾗ|	�{�|e��Sr�;Ղ��Iq�v���ۣ]�K;��<0x8hѠ��y������o��	�T���UU瘏_/h�t�h��o��}�i���=4nxl�E�_���'Y���x�����'L��36t��8sT�u�
���Th��Fx!�0�ҙ�����J~=��%ej�V�Q3��V��! ��'�m�n�_/��Z���L�L��ƺt�6{0��k,?;��>��ߛ|�GX�8��"#�u":�:���S׭4����J5*\�@�,ဟx��:�dM��K���I=
p蔝\F���Nl��]�{��[��@���%U[כc�y��zڟZ��>�@�n9UɆ��;=66Ʌ��	ú,p��_լ�rQyrd�\n"��06�>۷�i�����W&�vS�F�f&�'9�ۘ�y)�7.z.e���Q���&�L�$�����&�?o�9�ION��!��N��B���i�:�4�b�Q���^2��[�b��]b���_=cTţ�/l^1}b�b�kl/�X���/_U�W��yu�1�+�-�^1q��b����k�XƸ�1x���/x���^1x�T�H���Ԫ����/H�!�X�c�^1x�=f��������1���c�U�4�V��/l^����Vؾ+��U�꽪���^)�1�b�b�Q���X�Z�/J�c�k�W�/�m{mx�4�+�/JҰ�ivˬ]���Zi��1x�ŽQj��y����_+�M"��t�����/�^ظ���/u�5�_�ձT�E�Lk��^1x��_��m#�".*"���������5��#|�1v��[1x����U�u^��6�Q^b�i��m�tW��LR�Q_�o��׏��b���XT�zgA��N��ĭ|�"`�B�p`��]S�-)�QޗL�}rx�U�\,�bn�}̙�X�g3҅8BzD��u�-�,�$obӼ���MY{�[�Sw�P�ZV	� ݊�����1l�Z��*Օ����l���m��Y��*&1�����
4a���ZҺ������qB��$s;�e����|�޷}�����5z�}����.�k�ϻ�~��*��{��ܮr����}Ͼ��U}�����9f�r}��wﾯ�U��߾��k�xm�c�q��DGV�>Duu��M��m��׊�LӘ[KiA�dJ1r`�Ł蓑c:$�Փ�R��/��e��L�i���:�Ad����Z�6$���2I�a
	�:������1n���4Q�YH�7'D�8pلؑNM{���ن�C�	:��kr����	!%L�:~��$42lB������&�Vr.ω��s9���05l{oQ��f��km���"�4'�SF`1J���D����`PB�f�B~8&��z'���"�FD&I�zXĆ����<�`v��Z&�����ʲf~����� �>��:|���)A�?p{��n�����J�6j�FM�F� ��^��[Q�l� �'A�Y(�x&�B��2���82Obm��d��eR�+�������q���u�\u��4���M�z�~x�y�Gc�[E@����'����I���H��߼�����]7.p�66��8����bCiFI�����Z({�'�8�L,MB���O�m;{M9�[Xș9
P�����6�����k����zޫ����¯��!�����A�� ��!�@�``�2��w����Mh�DC�ݶ���,@0M��6�)��zP8&@�<l��[ ��s>.8 ~9,�D���OUXҔ����(�Sˡ�O�`�(���� x2xx��8l���	"tHz0�=(gڹ���,�C�
%?	聰d�F&�HlI�0�'�R0�?D����a̚�!?j�g�鐝0J@��a0I���%%z������M	��d�ů�-��i����:�q����GȎ���u��YKm�޽X�;��8�*�������$���-7Z`*�U8KQ��a$�1��lxك�D6l�fb�+���1�TZC���8"I2ǐN�)n�(��LM���5:����9�.�.�a�/���>� 0�7*��s϶�S'A֕��5� �		/���}�ȏ�>�=�{y?�;��۽��5����;�rDm��Nhdy3.'�B�J�*�k/�㸥s������կ�:�����Sˠ���OD�'�	R1��ГbM�0?I��,Ě�,ꆕ����~�ыX�^��( l"l@�!���,{a����nM�C	�!��m��O8P��X����P���˺i4拭`�O�O�B�0`�����n�2M����B2)�����9)8	��y?}�����=ҋ��:	=aA�H2~����C�&�𥁿V��>v06!�'u��0���J$(�CA�Q��l��#&аBCF'�	B��07�d'���p�!�''
Mp��`�#!��J�$����ꍲ��Z�G
4V�MW�i��L�]�� ~B�;�u5=C�IN��&�� |��(����C�"�$����ߜ([t� b�뭽q�~c�8�Dun��GQ�_:��iJ[m6��ooO�m]T��@�!���Ȉd��~5,�2G<�K����Q5$` |���a��7��<�C�2l��pI�d�8h_>n{�����vCtJ��[	�Nlh0�zLlK>ID�@� 11~~}c��NQ=�a8 ��l,�0���X���c!�{ؑ4R�(���G���32�ћ��������x�UA�i�*��Q'���@Ѐ�>5�z0:@�Ѳ�8$6��g��Un~э�p��|l�	��N8�b`��O��x!��!��p��O�=�rD$�qi���ዩ�#b�ӑ��4���4�n����q�"#�u":�:���iJ[m�hѳ��H���È���a�� t��td0(�f����H�s�O�)��n��aN Y��"hBı���B��I`l�62o��f`�Ї�1?�Ǳ�a�O�F*���!�����䭰�h(��!F�ДC��X�(�Ě$,�����
@��#`&��b{ů�{s]�~0�tjo����O"^�J�_�W�)�xڃ��@Q���:P��d�)����c�;I�t`� 鹿wh���q&����l�)�@�m��]�{}ֵk�?�9�Z�ǝ)��2��#Kex���:��PQ�405���\	I������E��»��@�m���"OD���}m��Bm��U�H��)�R+����?6��1�q��Du֑�#���ζ�JQM�0�FœKE𕈬QQQY=���qTL��D?��$,P��ߟ�J�Z�|�߰~<��tK���d6I4X ��14'��	�8$��Ò�;�R��5<)�"��*yРzs7�9kV3�u�IU����������2����vHz3�"������IK���C�)����ft2��&�4|S&���h���X���Ț@�`�û3�]y��W5����=��&���8!�I��a�X��p�$���jI�o�����G��C����4�L�e�e,bCF�Oc'=[ �(r��m2@�D�����h"N�$���O�:Rm�a�I20��a�dؒ{�h����?1��b":�H��|��/�!Mb�TX�x�$�;Z�Q4���O���� ��u�U�ʮ
l�7��lԉ�V�dsY�?\��Q�T��H��X�G�<m��"X����;V�l��X녏9�	���[l���lQ�>�E��F������a��L�s��+ȱ�76k껜"��:c"�)��̌���F�׮lu��;>Y�}/ٲ�~����0M�b &嫏�D�d/��1���&@�X`$I	���
� q(���Da5��f���'�4 �N0�`Q�a�CB`�B0Г�604y)����W��W��oIJy 3g6JzxV��DD���4�"|2"C�(2�-��(�<g�۾f�������}%80�z$<� ���h`D)���D	'6��n	��w?�?F�V��2#8P�0���n&,�<C�HkeFO�^z��ns�T�	�x�ō�~RD&�r�[ί���C�DD�����"X�0��G�00~HpM���CC%�Om�&��	�??<=>q����#�GQ�m��l٣F��i���X�!�M�5&��da�	���M�2O����o?��u\Y���z �?F����A'y�z[nI��d�!�~�����~<�K�ȷ�A���0A �zP���"!�P�d��dd=7 "�=��jd�10驰J��{��I�_s�FO"~�,hB"p���Ӆ��:��>���n��\�ԫ,��tEV2������fY�X��d:{(d�@�z'���h��8 ���C8�d8	��O:����>�~}҅�a4�J {V��6$�MF ����L<z5>4|2pA9=�`��KR+�|�Ƒ����\q�����_":������KSm�z�˺�IeChU�O�E �l�� 	z9!������F��(2O|\2M�M<����'�tH~�!(2M�}PB`�/ki��x$�â��0S$�D1���Q\	:�!�d=:&��}�%�e�v0�&Gfǁ95E�L�16�NBF�I3�ߖ'���u�\sV���&��sP�a�&�U���2r��!�)`�ԭр���2vp��$�����>5'��a����Ѵ�C#!D>�ip�z06$�6XN��L'�8%7�nnᅆP<�0C�W�˘#�n��pNQE����2CQ5��?���G��뭴�����u��G]G��F�|�lh���޽m������g���z(�� �����(�{��nό,5 ~I �HlF"#؇��80NICc!�D` ����/�sWM]fb M�7jw����/-C���������ke<<��NO�>�gD>=(x	��S�=5/|(jD{�@�"�Ͷ�5"�=L:��;�_Ə�,8{B�M�#���8��F�a�>[տ�:S�l�������m��a?H�~� &�9�������'da<��.�<�0gbz&`%1:%)��&���f�ߍ�� ld�ݭ�N�ON�D�e7(��J|R`��z�����F5���1lE��c�^-�c��/��_�|���i�5Lq�V��X�V+�c\W�^-�����k�WU�W����.1���^1x��b���+c�t���/�/�1x�b��z�+�H���1�b���~]�v�5�]�x�uxS�Tz�Ue���Skαx�V+��_Ub��ұT�U1x�|ƱX�q+�X�W�V1�V1x��k��/�׫���/u�/�b�[�����폚��k�/JiXV�Lz�4�V)�KҰ���z���qx�4�+[J������~_�Z�+��墽W��+�c\U�cJb�YU�[_+�b���ӭ5�W�W�~W�1�������c�qX�5��l[��l_�[��Ɜ�+�b�V��꺮����R��|��ֱKb�[m�b�X�꘨�5���iT�.���g��س*o���Ǌc�젟�%Н������zg��N8���i![���=t�69$��8�vnon�n7�Y\̳}Oy�'1����Wv�p�1�s%�L�Z��5��x�S{�t}�e���!&Fdf�̃��55�����;��Y_����<�={��8���A�����hk1�X19�~3]����n��5��J
�g]���)	���ovK�z�wY{�&ʨ�S���V����ǫ:��޾��[H���#]����oV�a�巽�������o@�X�ܸ�l�7���h�q����l]���%5w��~��V4�B�&�<̄l�Lw;�t���xfvPB���j#��r��e^���{ga�&����H"��c��rfC�n=�H�r��3,�B��E������-i�W���i6��Uך\wٳ��{!�\����O��qF-8��1�]-W4��ں�{�zOguW��i��d0�X�jp_�R�O�H�{�:x����Cr���z��5��A�R�kU8���6�5Ʊ�pN&�6h��i뵔��;<�z&X����\܎5�7#��t[ձ<���bVk�Ϯ�]��(�ΰ]!ߍ�۩�֋�1�جZq5S�UC�V�
��+MF�$F�\�Z9`���27\��%�[�Z�;n�,��O���cF-��nnon9X����W�����du�������p�J�o��}���}��>�{��s������w3=�������}������ff�33$��g�}�_1�\cu�1�Q�#���|�lh���޽m�uj�WW��&ފ1�9J��7Ng4qc��h�^���]����=�
1*���~��O�2a���>�%��]�:��4�V3@�D�#q�r+]�����/+�Y7lf�sٸ�nڴ�/]�oc��;NL�Gs�$ͺ�vݍ���� l����$�z������l0Rm�p�1�1T݃�!�{L/6�'��<u�9qNvl��Sرڎ5�/o������[v8mkG�z������1��G5��/�6�-�j�~@�!!p�Z���ڝ{��v�2P_!����y\�3�v�*�N��ض��@�l�9^�ƞ�.��s4��{��K�j0>B,���B��Jh��LA	�1(�b	~>\���w:"$���0B�<�X�S�5Q z0�h{Q
&A���ܸ�ό��?j"&c	�d($Ԁ1"�G�oZ���S0��80Г�2j"&D��rۖ��6!�N����Y=d�I�N	��c,C�;G�"1�@�d[�)�K(��
!D�0(2Q�C�T�ɱ'FbPI���?��6�'j�/'����nZ�3Z٘�M��"��~��F&zX4	87��"!�
!ұxTrL�>��)��6���뮱�G]GȎ�|�lh���޶ۨ�s����*�E��xh�0>)Ʉѫ'�{�{��g�}����w�\�֦��a�΍&��A��O*�`|!��3�'����{�A����M�O�6���6&�Oٖ�<�Jh�404t����Hh@(�|�|��q)�C�ҞA��L�h26O�$���&����J�nbo+�K�n�KCMK\Ac���NG�'w������煹)���SBPI�� ���|~���f��Wj�<��kR'�Ӣl�hh�
`����(û)N�0��A"A6t�\7>>_�}��ߥyM�z㍺���u�1�u�|��!�ζƊ[km�f�3iU��\��QA�	�?<������|�m>W����?=6Q�C�	�pd�$�D��%0}�S�4x�4脠�S�5���Q;�ic �ϩ���07�%�bi۫eY��EP��"�e��أ��֥�a臂hK8?��a����W%�5���u��zQE=_�nUW�θ�"�ҥTOa������%�C���ě�B��r���AD��7o�.9����"2{J�PC�{��0Ҥ�7Oߢ��8!�Cf҇�E�ȝ!�l���ףX%r��:~:p���뮱�c���#��_:�)f�lѳg�5�E"���!L(�����C�},;>)�=�j�S|����Ȕ���0����4��t'���]M�i�h9 �R�_M�:R�\Ң�xv�(�Sa�7��:aK:��ϧ���}5*��'J
���ֶ��n?y6^�`��[~�8z_��3�:{R���� {��ˇ5���.�VUQy2�!d���zL8p�5~g�~Cҋ���#^y����vSz�˽xM�67��x�s�����S�?1�����"1�#��\<l���(ن�Ůަz�Mee�K+��p.)�="�贶��5,NI4Ń�f�S1�Te�����W$�.HمP� v��jҗ��͍�Y��x��;'B��Z�m7i\`wZ�=����!'���W��7��6�R�;tu1�ᙙ���Q�B�G��3�weZ�ThX9S8���ݞ���7�^�{5\�_N�	32_�aI�N������Bvx}��h�X���k�M>>1���s�}���:s!f|<�����-��S�&�&|u���B������*C��h�O߿3Y����A��g��!H���?��V罛c�U�E?4~E?U�^z���Fyj|���)ּTY,����W����gaL���6M�\���1���ap�\��S��O'�|��!��t����\9�i�32�k-���\�U~F��#�κ�1��|�u��[cE-�޽m���I�Y���M$8(�A,Нz��7UU���v���4���v�t��y������{�m�Ν[S���ժ�����~Y�/.]�[_��(�X�d=�	�������p�h����k�������YA/����Д�M�+Q)$�Y�α�@ͮ����y%�������4P@��~�{5��Ԛ�bX���|�&�����J�ptx�Z����Ww'ŔYÇ�}'x��~c��8����F>cD:����Km��[s���U<���^Z��kN�c�>ݷ�%*��_:YF��0�x~c�W��-�i�4QG���U�J�d��o�~g��Ϟ�~kB_�5��]uNY88�VYV��5���L�\ˢ�͚�v{=<8Y�U|zQ�<1��}��X��]+�~�r3_�+�������-߇Oߗ᲍�S�i�>o���_ϛ(�<��*��|��W�}y�w�8QG}m�Θ�Z�њ50���a�A72d�r��m��zמw�-�θ�?8㮿1�Dc�1�C��m��͚6o���YZ�o�!����>�������W����'O���
:w�t�[�4X@ϻ<�v��6ώ.��w'`Sg��b�Ѻ��a���Y�ldN�Ǝoͯ���N�5���;����>DѽsSa�òPC�|�<W�:�Ce�y^uս8w�皹uz�:��G�e*�Ux������l�:'��Ι=�~>�N�y~o�&���e�il�Wγ�F�-��8��q�c�F1�:�:ۭ����o[j�骾׾ݞ�y�^�1�:���qq�+�Iwj����q�~��d�*���ƻ�S�"�{mDw@-���H�z�ی�m<-�/F�#99e�ƣ�@�pHK���Q����rM-������, �!ɑ@�j�����������YT�ݢ%����޵���]�VR��/
xY��ٳ�&��M�>%9��g�ЌˡZ�O:&8&k���(���+>�����\0��V`|lѯ���l��┶��}9,,��2���e,��<a�E�T��nʆ�S=U�N��� ��@ц���k��n�&�'5:3�֚4|rL�p��a���~�aϷ���	��'b����Lʪ|k�ɮ���ϝi<�4ۥ��ީ�f����y]���諣��8���\q��1�u����lh�����Jq+4$���`ʺ࢑f[���i��|���޿U�!�JmJ1̻�������0 C𙪫���0�`��#�0��5<<�WAND�0CG�PM�E���-�a����4	HI)�?|'g&�$(�5|�(�����̅n�(�j�-Q�D�J BD��ˊ���r�6���>i�<���:����:�������=�2|iT���'��?~�)����jq�}��ߤ���>�|�N�R����ǭq�����ű��/�X�X���^+�q�bыڴ��1x�����+^+ǫ�.ؼ[��k�:���/�.��^1xڗ�^1x���c��k�m|cMc�/�bⱊ��ⱋ�-ڭ�ڪ���#H��׌^1xٍ~~~�~m��/������YU��X��b�b���˪c��.��R��S�V+��c�uX�V"�\S�b��c�cX���ǯZ�^��^1x���5��/c\b�W��k�˶/�+J�W�4�b��b���ũ�k�[�<�EqX�4�⭵�N���/�V������Tj������~T|��k�R�X��z��b�X�+�Zu�]_U���~~~{k^+*��c���ixV+^+�����1|S��z�Q�b���8��S�aT��b��[M5�c��W���_T�����'Ŝɻ����w���@H�ds$2�0�L���.��	g!E�L�C[(��y�I�Hq��(f,����!6�h�?c���7��j>yl���'�T]>�v{���bk�����/+,T��<N�g�J���.	�Y��� }�1��os~�9Y_w���w���߭_�|�����7�s��>��U�W>����Ͼ����qd�$�3���O��8�":�F1��c�u�u�[cE��޶��6(�A;��v���E=��сޜ^�z�sr|<��g�����5�o��´�:x���e��/�2��0��P���+i����L,N�)�>O�/��N}ݫs���5��V��V�#�Y#n�+��+X2��E����MO<�85��	�
l���o�M����7��oF�D��x-��I�|B�X���t�j�C��������r�S^�E|�8�����)JZy��m�jm^�Mo��w�KLʍ�h؈�Vc�5ʯ��t�}�4���q��κ��1��:�bm���km���*e�G[PDDO�/���ߵ�˃��f�0��L8h�"n@�����Jz�k|�ߞʥ[�:�)]���w���3��S���C$��C-��cj�Tg7��+ϒ�1�JR��Ŵ�<���wM)Lq�DDM��٩�xSb""ǿ��q���|{?��DO0�J�x����2��>��N)DD�����7�V�)MuX��ֱ_��w*�돿3ɶԥ?yg}�ŭ�ʹ�1X�8�q���1��1�"1�^��-m�������}�S�ո;,�US&,q5��-��c��U�I�&��ܹtaX���,ݎ}w2<,;H��+J�(�q��o��T��6)�\ld��Ր<�b�m�nv|�h��h���GcEj��	B���b�y�\X��?���6����B��m�K+�Yc��P���"�	1�8��1M'[��޼��1�.&�!e�Z�����ܽf��Q�aBae��'yz��~pឞ��ԛ4l��t`����*���՛П�Յ�����C��ㅈ��|co�+]�8&=ۇl�Z��Gޝ6"&@��S���>7?4p�fbϹm�8R
M��B�h��{��Vv|y=(!��qR�k�S��0��τ����	��kLb��@%c����[�������9�;����>0 }�������U�֪m���T�c�>m���u�1�#�F0��[cE��޶�Ɣ+[U*�(����
O��#?I�����	 �Mu��֫׾��#oT�(��V�~ϛi����{{�e�����f�䛯YU���0 Y
7<��Eg���?? �<5,	ϕX��=���r+kCi¹c��]��܊s�LU��Y��t�����O��l��?up<����~z��11^Z�<�N+�G�!�w�������ҵZهB�������]u���1�"1�^��X�ٳ�?v�V�t�4��|PA1�M+��Y}�?e��+V�mE9^����\�����@�Y!�\��J�=��֝W�Ϫ�|��n߿Um^SJH�=<�r8@@R����G)x�c��F�$����D(���r��v?�<6!INx~�b�k��[�Bt�D8xd��i�b��?2���<�|$�u�׺��>4_[Q�_�x�[�>�J�������2��NB�s��<���y���/Ϙ�8���1��1��Q��m��~s�=��<����r���X�th�F���`��"��i���DC~~�2��ݶ�f�]��F%�=�1�kV�u�6l�D��=<0H�Q8����ϛ��i0O�?a�����&�+��txnjaOM�ꌆ���z�!�����0������,)��}�coˡf�7��M���&|gus�~?��*6�<��|ژ���0��1�~~~u�_��#�b1�#�^�KBk(����F��C@G%��U14��r��6���\Cݯs�fff<BlcykVy���؇7#��;~E����9l���kHb�~Q����-sy�\�z�������?� HBX�ͭO�o����?Q���3��V�f��w�Ӳ^�<���K���NI��,tWL��;�����N�r�o|���<NM�s��O�z�7����S�Q������6�z��E4��j��j�m�zdW�͸@O�{d�-�N�t6Ok�L l�'�.O�&co7���5��~��MC���}��F��V����j�.���[nyk��Q�����6��xj"D�R��R�IDTrj'���O����nu�ɬZyrvsvw�����w�m;˅��lG�}W�R�:x!��W���x���Q��Z�d��x�ߏǎ=q�??:��c�1�F1�z�Q��m��o�;�����ﯭ��M�7�O/)[��>7g��;6s�e3=8S�'���S?�b�����_�2:ZYE�L�Ӿ�$t(���
""��W��x{�仺ʪ�ÂQ�� o��<�OҞa�Ѕ��iw��̮9K�9b��Ƀی���e"!(��Չ5�w�W���yTB�Jq��!�)u��Tw�g��)�畴��tvn~�l0Cu����~���S�im[u�q|��u�X�#c�cc�z�-Km��f��݊("��<5�F=��}Wu}�Hl�a�D�ޒ\�c��ׁD;7�����֮�?	�qJ)�����j�1��(����Ӂ�'$���� S�/�-.�0�{�*�'�u�Y�� YZ��\i�>g*�SW��R�Z�)^�1��<��˫�6��%��Ӽ���B7�hΐ���N!���t'=!�k��6�Ex�[�����c������b#�cc�z�KR͛0����?FL��u.����~�("JrS0,p�w�ѣ�g��R�;���Y��� �y��3V�5���d���M��+�3�6��򑴚-h�CS���5{U	})M�I>;>�p=��t؆�|T���^��Ν���f=�r���ʪ������!��E����,�N����Z�:�s�M	B��,ȋ�Ӈ�'O�QI�_�~|�~~~l?}�6c�4�ȤGȈ�GQz�����DG�B8��z�D|�"�DK�&:t�Â""aDD�DDD���艅�����DN�'�'�:b""=DZ"6���H��8�"8�>uhY�""6�Du#H�����DE�M-"4�Q�޽z�DZք"-h�6������ulb�a�b�F�R8��GϘa�m�)�DDq�S�=q��!�1DZ����#�iƑh�>m�y�R�H�=F�D��{�T��/�*��fHO�u}���OZӃ��2�B���%�ĺ������3&s�Lί��Ն�k�（��ϝ�گ�����X�{�umy���*ŷL�co5��o3.�d�����X��P������B���z�nܒ��p��z�j�s�9_L�I�	����Y*w�vo$���r�W��#��v�-/�ĝ����Na���_�7��W��֧��E�}[����!ikn��nf-��y��uZ�M/GoćD�
�8q�H��.go�v���\[���~ۊ��ӿWg�h��ܶ��|:��bPm��d4ύ��I3R�XF��Qـ���IB�nY>�V�^`�g�UΨjr���
HY��@�wr����d�W�۲�UK��?���usa��G�U�����������~�z���s�e��ֈ���l]1L�v��)-�1%�<�h�z�{Gc�x�Em#:a�h� ��Qf����a}Fm�����~���k;�k���kѺ�[0Y�tt4��d�%e�9C�*�mme�r�g(�u�k�n,Q�ܝ��87V/�ú�ֵ�ł=���N�9ݳ��Aݱ�ɫ�n?M�\�J��;B�[ͼs�܏K�5����${:���2�"(20#��p�y��_y*9��=��_|���9��}����|�W�+<�9�>��U]��s�>>|��:�c���#�&,�l�f���*�N�f^u��.6���ݹث�n7V��ܞK�)���t��o<;g=�3㵃s�MZ�s�����<b���8Mƨ�[�ǎ2r��x�lF��%����y6*vn9j�v�\���H���姲)��w�h�M�n<�"q��G �ד�!{�\]=g{v��ӷ�*\�t�F.tة�]������ü�d1G�Mc�5��q��u[���+���ݧ��Z�j$�T�>�	K)�l���-��ߛm��r����h�������o��}���dph�P���L]�9��nW������i�oo��o�V�����4���������My�Z�T1ׯ����ׯQn+�ijy�?^�D̢�}��6a�{
lΎ���p�ߧ��\:l�4�%��N�4$b9���8`�Fp�����������ߏ���{%�NI�=B�۬�ED,����l�{5<5a,V�Hݒ%�J�@9�$���t� ���T��b���Q<.�g�9��'����inQL)i�\�*�TՐ����� �����u�1��DF#�=G��Z��km��眬�=�U*�Qc��4qX~'���!�%�)�rIzu��ϴl���bwS5�u��<Y���2��n�]5o�F�?~�P������p�	�>�V,��_���&��0?G����UMKo����#�jFQB��^�$�����,�]'j�g{�H"c)_����^k�iJ'�?|�o�~Z���8�-�uKO��T�J-Lͫ�2�{;�e�K���6pzpOƎ����#����cc�6�0�)�e6R.\Т�!��2jx�U��֥�o�yJ/�G���M�:lІz�ba�|����NL�'�9>�/�{���鼹��H�T�L��B�y�ma+�Os�[�U�n�t-��+ʿ/�~E�H]z�<���)��]�{sWz������r���4d�Ȍc8h�L/~�s)�rM�K�D=3)}=�9$�I>~J���%B����(�_W��>sͶ���S���κ�]c�1c�6�_4�)�e63�$Ό��ex(��uKW���*�JŸ��ΛQ��f��
!þ�߄��M\n�kC�
���#`ϖ�2�ܒ�>����Ç�6a=إ������)���ݠ����A8S��A�|74"!�p���K2g�l��g������4}�c���F B���Ky���g
}�ˋ�Ɇ��ᩣ��(���xc�^}��(�kZ���ө��mH�#��]c����c��1�mm��m���}�מ�U�j���ɐ$�hpv\�cve��]i��z��c���P1 y����j>:�cEu䢑KS�2�����[LRX�[�ש���S��Ì���3n;l�r��-��nUTcm�J(�%n�fb�	KdƷ�go����E�����Ws�������E�@ -�<�|E�d܁,�X_e��죏0�쫭���k�<l�h��YL)���B�Ó����R�h^Ώ��O""!��5x��Z15��10��
Q���[����R�̓�����gL��]��?L7����
!������K�������}8Q86�MC'M���b���A�����etd�l�pU�:�cVA�T��`.����ч�a�b��$�A}�9j�� �DT�V( ,"�	4kg`wگ�\.��	��p��?8��u���c��1�m�0�)�e5��m"�7B��6Sf	�CA>)���-,Ѩ�u���g%:aD<��Oơ���>8~W��M=*�u�-��iwW�[b��)G8�h�����>,��D=�۫���&��u���,���//�r�	��^�7^�!�a�=�<' MS�jΐ޾�9ùے�:C�Ő-)��4S�&��a����8S��T����m1�:�]c�1Dc�6�KZ�mo��eW��u�EC�p��=�S������J=_K��gB��0����'u��ag��˺���ɒ��wPuE��~«����Y�K��^ܽ'�X�k��wQ^7m�6pG]?�6x�ѐɭa���o�w����?��m�Ye'U"L�|O�Ha@��%�X;%B/�8=2l�5���-:Q�
|�=�=.a|��قq��]�)���5�ߗUM1�����q���u�:�"1�cDc�6�KZ�6R�`���%�����Ø9�U����a��)D=������Z�%��ǐ�?ؚ�e�Dy7��t.%t!��h�n�T��WL(����x��|�k3L�D:hA%��Y�G�h�#�$������ɚ�I��?ԭs�ԧ�nT�x�/�0�~���9ed���T��I�x�_*WO8B=Ja��a:t�rJ!�7F�OQ���Q��1��#�O�����e�QF͔s�n拔�ܙAŢ�����T�ѷ���E��f�̩�D�hq�·�lB��M� ������4\
,QUE��k5K�&37q۷n�����k,[��.8�܉�O��B�D�Uco���bu�gn#H��i�[�h�m�8�oG7�&�m�Fn�26�4:�mr)Ә��~ HBV�&������K�W����8f���{���(K�";����W=�o�ns�΁�H�)�`���Ǐ�e��w��.����s�ܹU�i�����>׏t�@�5/_��<J�O	���
����OZkΆ�Q�����=C�F`z0�hG=..?�˱��QkWGC���hَ���PlDD5<WzC�?}m�����~�R���*���~��ܪ�������Э��ƔU�Р�@j�L�d�l��v�L�	��o�̹���6�O�%uh&2�)�����O��|��q��X�b#�b"1�mm��m��v�d+R"W&Ւ
,J�(�5u��R���,���"��qГT���EC����۳�8pДD7�G?am+�کR�^�x�X|M����8�ԾM�|����}yT����j)�Uǫ���4pۻm�膁�qQx�=����2��w�n��e^Δه�ƍ�~0��ڜ�z��]&��x��vn���v���j���y�����k7�B ����?I=�Ua�}'�F@��P��%̇�^~M�тB3ɇ���~N?0�<��+e\i�>?8��Ȉ�h��GȈ�">DF��"#�")�"#��a���K:t�ӇDD[Z"#h��">DE4��D|��H����8��un����""#h��M����#�"#���!B"��-DR4��">u��i��""""""#�#m���kZ��G�[z��=b؎��iht�شF��Q�":��M��X�)�1�cn�qŸ��c�1�E�#h�ȋq�Z4�6��y�Z#�i�D�Q����.]�h/�[��&��&���_�7�u����I��l�8�kl�^�R�7^��wVo�fڞ�ߚ�A��v{����KB���ś��|�d��7g[䞜ncDi�S9�ͻ����r,y��J��w�U�{�#3��J����RQ�t�۹ZlӐ�o2Ǔ���q�Y~�"]i��
��U��`���!)"��}y��f�'�-͚�yC;b]y��ھ���_�g2_2���fz�s�7�߽�˵}y�s�}�֪���k�s�����U^/�����9�p��1�\q����b1���0��f�6l��<��
("�%�/�l��Ç�;�m>4Q'K;�5��DC�Bt�,��J֟�Y����4���7�V�׌�V�6"	w� �4O܎6ݖW�r+H6ڴr����5NX�V� �
�-�,���b߶�R���k*�mGim�žz�L��QJ�wΝ�U�>�w�[�qO����QЌ]��l�0a�ܵV��&�D �L4��'��ޭ��8�X�b#�b"1�mm��m���}^A@%gY$�ָ(��k�-�����^��Dό�Y���ȉ��Rϯ鲈f���)J�'����4�N2IkM30hK0L����p�C�!Ą���6����xaD6%9��[qt%=_4"�0�0�a��M{�b�C Ld�gg�?�k�r}wVY�#�tu�pؓ[,�ҽ'
��6l��e�k�9��ǧ��P�p�_��=?M��<8n�("�[�oǧD@�y(����gȎ-�#q�1��F1�1��cF�ik[m�s�m�ߋ�7Y��n��e������Ks�c��m���vӭ\d���z��c�����$]�����9�f�����>^5����$!(�������}a���׈�;s�ݎ�Y�a'\���pr�82A�����3"��8Ɏ���X�@1��TXT��}���m�b��~�l�ޯ�30�J�:~6a�Jp�~�R����6iE8����U�9*�D���h�S&���?�XkY�����6���ᔘ" �֛r�{߿8Hڢ}Z��	�	_؛�Bj���UB��� H}N�*�G��2Z�bi�/^�R��������G���w��I��}��}���z�m��q�c��c�c�6���ֶ�[�}G��;KT1�E'�vD�sҲ�;5:�:x!I9=�g߿w�\q݊>>0�؆��h�a��٣�8�x�5��Ӟq�[[�s�^���?S�N}�*Wb'C8dDC�_�k_�_���Ī=V�dv5�\Jn�\`q �߷؟��1�����4S�Қ\(��|~�~Q��,<���\�-�s3��8!�î���М6@�J�m�U���ee]ݕs�ÂM~�N:�ȶ:�:�����:�1��16�ֵ��غ_�U~�!���\Tj�	K� �nl��*���6!�P��/�6'�83A0��7�J��E�f��S4}��g�&1�����}=����u�4J����&���
2��s���7ӆ����؆��'N6�����ƭ����W�g�u��8��U|c���8�?S�wkm�󯵇5�(:C��&VoW��P��~������j�8Xa��Y)�p�H���~G_���:�1��0��e)Jl�����آ��T�}�G�y��UJ��l��}�4
J�`��0����@�8U"+6P���6}���k�B�Ÿ2�n��0���+��[ vQWS|�&�]�ij��DZ���Yj�.��`rwsc����M��=�����6S��/�ܢ��Ķ��E��N�}���Ut�H?�E�rV������Pxߎ�m�{�������M������m�/��?U_�#m���c�8���F1�1�c�|�kZ��ov7�������h�# r��g�D�-X�d`c��
eH+j���̲՟��--��peLv��H��4�l�3�)���ח&_b^�����tW���)��8�.���o�r�$RA)�ȿ-����X���l����O=��k8+''��ˆ��wdBɷ �L��6�UY�����~pn�/J�y`v<7����ɚ�G��<��a7�ч�~���\�V���/�>�Cf��(`�Hg݌�w�/_��a��o_js�0��W�
p����|h�z�0��߰0��|p��]�0�wl��4�CBRh�ɢ�'��DЎ���k�bi�H���*��j�pX�',�T;f,Z�U�N�!��S��>MD�5�>Მ��������|'��?1q�"#�X�1�c�e)Jl����X"o��k��;'�!�ֹ ����?]��XaO�򇿦J�/��=><&����:xl��ך=[�e������UсD��y:^���Þ>���{G�DD؝��A<����(�H������&�Ί�xv{g�c���U��<8S��f��FҪp�0N�-��-�t��<,�+ϼ�yʫ���G����m��~~~u���:�1�c��e)Jl٢���lngQ`�v�?�C9��C�?zz��~���Cbl����g�T���|�����=���CGB�~2CK�S�a�AжJ��&�3v�5۲̩K����x~�Ò�3��?y�W��!~�B*�Ն����']q�:iӽV���ϼ��=#��xDO��[�h_9,/��(�)׶���̿Dٓ�~4~��߄�xtt5_s0�~��Æ�w[:Y��0�F#�8�Db#��1�cӆ͔�)�f���p-�E1���:��Q`�?M�\�0����g��.���<?�ٳ��ib�im_�1���L2���Щ�+IZȤ�zީsA�RP�Ü��RR>`U]�KQl�O�Z�M�G�j��������<��0�]|[��/��}�.p���I�c��Y�IӇ��&��,æ쥲�S�᳆�~7)��l���E��~���ߎa��,x=yʈ��ܛ<)D�Jd�"��_���R�i�ϔz߃�Ҽ�W��q��b1��6�Dz�Dqh��"�DF����">i��G�""#�T��8㥈����0D�8""u$R"!�DDD|���V�#�4������E�Dm�ǭ�Ԅ!H��#��=F�h�"#N!���F��kz�DZք")����R=q�1�V�Lm�cG^�B#��4���i�:�\q델��c�""":DR)E>Dq��ӈ|��H��L<"%�t���p��پy�ݨ�c��ȞG~|�p�nJQbs(�L��(�p�A��7k2Bǯ��w�`�fгq�i���I3� �96Mj�����2Ɍ2p�ʭ�ȮFU�ȧqnذ�ڪm��[�2A�tέ�`<�����T�8�(���#��	�opqIqV��3?^�ƅ��7Ǟ�75��k��M��Ƭ�y1�!��^Q�>�##�N�+���X���/f{%y9�� -� �m�]l庫3��"7�a���3d؍����s#S|�Ǔ�y��S���.n:f)�t�G.��bw�Y��&B]@[-������"h=[Ɂ�̘�*,0�*�+��꒘���+��v�aX?m�������ٗ��2b�N�V!j�M����۾��t� �q��@8y�m�3��9�p8�k:�^�a2q�;��ծ�5��{���9�XQXJ@����:�F����*��|���qr8��9�7]	ۡ�HI\k<�X�k�����~ ���;�.���w����a�ե�#�[Vd��N�A�c=�	u��4k�G>{.y���vp�}s.�/5wy�F^\/3/2��R���>Ux���>���������*�}�|}��}�~��Y''{�g�߻m�1�1�b"1�u�c�16�ֵ������ې�!nW�MF㣇�m���Z�w��0`�c%��]��a����ۗ�8<)Лk�΋���S�v��"��n5)�if���v�˪8����pl� NL�>�p�v�϶�F)�R�&H絳3����%����%8.VK�F���n��$��kq��N4�vl���-ƪŹ�-v�Uw	�<Kt)r�M��^��"`�q�nv�v�ѷ=���8�Í��.����nѤ�q��I�(rZ��;O=t[O[�ƃ�[x�*�:�v���� �`��H�i�����o'݈�B���WѾ��
w�uܚ�|�.��1�T��f��N�����y�l���r!��Mj��EQg���іSs�i�Z�V��p�"n~�WF��`�
t�v��us��p�;�4�;0�ԧ�k��;=�pr"qym5��ꩿ�$�pUU�O�����6xY)�L����f�鸘h)�ޮO�3�(�6oO�csT��AT��D#�|��|@���U'�;�8vI��{R�@��S�(���K��᫖��|jvk�ki���#�qq��Db#��1�b>m��km���<U��I��.a�1bh��UC��E�S��QѨ���ᇟ�߲�zl?D�))HH~�6hב�E"�~=��ϲ�ѩ�OӮ~m:= �蟦	�BR�|S�p���һ��M�0��[o�Jd��}�|�kz}'� C�����x�/�ԢXfd^�:�6����b=><�|�7�;�ó��&��O�����{w���Lp�S�׮�~�Ĥ��͞����.q�	�q�|�^uo_��ׯ�θ�b#��1�|�խkm�O�nBBM��'�	�����5�/�ڧ�h��SaL���鳇�:,��ac��f0�56|l�rK�i�����
D�Z��i��N��F��SC��DD0�,T�:Lm^�r�U�<tOi�̈́ CP���x�]f���|��:㎽--do�<4j~>�b�=��4hMMa�%=g�K�퓇�k��_������6�^�����m��=u��~G�#��c�|�խkm�ɦ��SJ(�Mhp᨞z��wƛ�i�O=,���]�|㏼�ގ		{?�J@���B�����q?��	�5�C%X���.���j�w-��*J��sS���CD�x����U!+��T>?@�����A�/�Μ,2PK��᳟��G�ژ8!N�L�zf���&�>Q�?eoO�ms�\��(���0,�%?qDx�:zjznhA=?$F�<����0aD����z�θ��u��:�1�?/��U4�Mb��;��ř���^~	�63�n.r��?.,��\.e��0Yf+Tqb��e<k,��u����-��;�8�ہL�\�������G�oe�\1�=^���ã��D8���Y~��Xشlo����wZ���Γ&|�����l��m>ޅ�5�\A�n�#}��W^�c{3$_Vw}:��C<w�+w�s��	Ϥ���y:]��K��bv}ެ�ɝ=��1.[�Р��\)��Ҕ��L��Q;��33a�5,�|��6����q�W��=�OV���<�h�����AΜ5g�ᄖ`����U.x��娷��z��>��z�]�@��%���V�l@6�+�~6k���A=�D����N��h����=cq�#�먌u�b1�16�kZ�m���J����^qX!��X?��M���|��ݚ4n%4h)�O[���<0���(ち�~|[om��<�F+Ͻ֑ي���O��?��5)�f�R!�]�E�}�p�,�9�)��=s�;���i��z��j�F�����[#T+��W9#t���b�̍���?���>}ÑDB	G��
%z}�%��'u�����_�,Æ�~�a���XC'�.���̒gN��p���@Cg��8a�u�G]Dc�c�q����Z��l�Zg��UUQM��W��~�����Ԛmx��l'Jx~?���	���T�60=�rL?n�}G�,\���ٳ
	����E���!�`�}�6� ��g%O��_"�B82ɮ�fk�I\-����bQ��旿��3Aw�M������C���ϧrt�R�)�Fl���4xl��Ssf	��m��+�#:�'�S
j��?x��]S�-���1��[c�8����Q�c�c��ӆ��)�bHmE��iUM�����K���tXlG�'�9�G?�J/�Y�.��	�ln��e^Q�̖AfdQo?����r��↋�BE�Cن��x8b"'�/�(�HY����qi��p���?&���),>��wQ��j˰��:W�e�d8}�Ě���Kֵ�����o��x�+��<�|��Z��F��g���5������ύ=~m��D|�����#����*�i��b��XgOc���F��Yy���s�[�]
#���ݳɋ0�7�a��{p�M������n�.�����-nݔ��غ�Y�����պ���*9%�ˈ�k$��~�BʟbwL�Ϳ�����1��|�����f��3:����Q�:�~ى�ۿnb�[�)Y�&�)�)��y�坛���u0��a��Q^/�n�6���Ⱦ�J�V����A<S��M��7���E6YA=Z6��UdQ��*i+��quu	�ڕTƜ�� ;@��<��)q�����
y�&mp�3a��x~�8|e��S30�L��tኝ5�Z=�<}G��^�.T.�&e֪J�tp��b��Ǘ0ƾrb��1��z��UܟQ���p�0��ѬL������8|'�O?:t�N#��8�1��>ch�֖��ܩ�Ĩ�L�fZ�'x��vQ8za������#�>Ҹy��FG�����J�a��fU̼R{^0������}_�T>鉱�J�}��6Mtܓ5����̅Uo�5�O���?|�:[�KZ�ִ��pnV(;A^Y!\	��#=�U~��$z��96h�\3g��'�� ��xj"f�����95��t�Â�u[��]>|m�|c��>Du�8��DGQH�"#JDDi#�G��-p��G][h����G��؈����DDDK<(�u�G]uN��)�Dqh��z��8�뎢8�h�!DR"">D"=m����|��F��"""""""#�m��z�DZև�Dih�KDDi�֑���B�8�=c�[a�GG�B#�DG�Q�u�zێ1�|�1�=c�1�E"-�|�G^��F�G�|�h��G��QDF���f_Ebh�z�Ӥ�A��5ګ���t�6H�;Xg[��Q�L���u����;ؘ���P$�`�k�&��o�����4s������2L�v;�~��OfAw	dH_d�����G=��5�=�y;�^ww99����}+�7#���g�ʯ_{�s{����?O��U��{��o{����U�rw��}���m��b6�8��:�#�c�c�6��ik[m��UA=��i��ѯʞ�[#=7�[^:��껫�W|s�X���y�uXp�	���!���	��	��/3��BQoV�N�ʥj񖢢��6ܒZ���h��rE���EN3"�=�\�s�*��Q[�zr���@���t氽^���0�!�q�� M�M����>�����xB��U������8}5�%{�ҢΩM6�GGq��u�1�F1�F޴����}@"G)J�F�eH��8��oC������Q�<
Y�:�&�!^U��M}�����c;�7Bd�=s�qҘz�u���f��V�������Z��UP@���O�����!.�[1�0e+���ST���U��QY�P�c �4~�y�;/�A<�������0�R������_O-�w��A��	��N&Mt4:0&���69���S����S�4�9M��y��y�_��8��ߜq��|����1�F1�6��ik5�9�s�@m�(7\� D�c$�ZV�~Y�� <�f9��:��#�U.VE2z�C#��\���۶k{N�۟KrX�Q���\B���@�����6���7����z}�.�F���ISV���|k:���u��qD�����~�g{�~kL.μ�&�$�"�7̳2To"�5�!z�Ț��?ӭhnG���6y5N�j�&p�QZ��ʫ��g�x���Ptx3�~������t�D�y/�6[��˔��|���zz�>b�U����{o��ٱ=�����z�<\F��~�[s%M��RU��bb}Jl醃e�����79:s��a�ן��z�U#�_�c���8�|����?1��6�ѷ�-km�^x�P����J²T-�* T犨&MO|kCF͟���l��B�	��奵��K��4;?a�'��jt6l.�:�h��c&�0�͘	��2�|ƥ���SG�y袧
��D|�?���$���4S
h�A�����Sv|ɉ�TD�n&�e�
.]5sG�wwn��nr|t��𳧆�:oVf�~ߏ�?SV]՗~ԟhqn����}���8l�4�m8o�=|�믜F8�8㈍���8�c�m��oZZ��oUV�n�d���������a�xy���߮��:�?�'�M��O�:y�'%��Γ.M�0��:=��d���hÚ�Q���v��Cfj��Q,�u� (ϖ����Ǩ^�C��V��h����k����X�Ӄ�q��5��v�9����!5Ԣ���9R�~�[���,A?	�����q�ו_��N#K���VߋR>i���Ϝq�#h먎#�c~6zlх)M�/稳j�	��2�����y��t�{�~?7��:m�ߟ��_ٽ��_9'�&��\l�h�h�gڞ��������Q'4x�I����Ð�`NY�����+Xc)�~a@��Z%�	�F}���j�9�~��-_�}��e��<<h��陼�@C<�D�Ej��D�����'Np���������q��:�#��b1�_�/�*�i��b�?1��*]MF�7�a�u��ݹ��`��Q�i�������5ت�t�����G����K�g<'�H�ݞ�k����m�Q����!H�wv���g�Ȼ�Χ�w�q�O5U=����\�U����}f޶=���22�����;t�~�O�Ww0����/���ڥ����Yu��N�����$�I�N���|'&J~���g)�8j��W��áz.}RT�"^�s[x�<_�|P�`���\>��#��6އ
jl��xsS_����tf���*�檡����~!�r�~?�l�}+��!�y��m����Z;,vg��αƓRܥDGӓ��_���'�3��د]JV4��{�|��8��8�#h먎"#�i��oZZ�ٲ��CJ�	���d�����@��O���ky�8&���h�aᱻ,r�~��r�p�s2Y�Jө(�ؖfI��d>dF��.h�}�'�M�iV���!�%S��u���>�L���Q�.naw�7�!Ɗ�2�c����un�FK�i_8�|�m^z�h����~S������/^W�\�ag�>00�>�]U_�J��ک�i��[���X���8��6����":�b��6����f�p���sS=�$��O	r���+��Uy���׊��X���6��'x?`ht��x}��E�;)��Ԅ�`��~g�զ�u�E��1�ɺ��������';����K���_��i!����C�hC�ǿ�.e�6�:>3f��D�l�D�M�;2U���ٮK?Oř�kW��^�Wܓt��z��Q>�|�|SO�|����8��u�Du��6��ik[m���u�[�U�=[����؃:,����'`��D��p?AB���n��.T��*�\��]]�͔x���.J��a��#T��wQ��fڣz�z���Qa��L�=[��7+r��}ɩ�H�zx�޹B$
�i l0���td�{�R�����N��h��ϡ�Ä!?�6�d�pgB��
5⼎��4�u|���#�GiDD">DB#��B"#H���8����h��㏔���qH�GQxDDDH""""xE��#��H���O����DZ"-�h�":㨎6��B��DD|���Ǩ�"#�[��z�M"":�DDG�Q��iH�-hB"-ih�Dz�E�R#Kp�c������Dqh�HDz���Dz�]u����1��ű�X����)�bا�c�8�>u��4�>SoV�!H�=DmH"t���ǎ����	se��U���&Dau謶�r+#ؚ�b�����:-�W����L�WEwٹW�˯y�h+�`��y��b1�G��q��6�j	�Ri!��'z>f�LOSk��.��Ūn�=�	ͥ��Y$̿,��Z#��3���h�������'޵(�d�bd!_L�W� ,k�ws�wfM�깛��?�h���O��f(nY��"ژ�F�"J�8�Z@W6+5����IH��KjB|��o��E���V/<"+���s�{���/W�N^�~��e�o��~'Y�"-o-������߽�-͔�5�J�cY��9��2�7��N�D�\�n+߽�Ӣ��^�2vj��n�a�p�cmW]�Y���� G�k�F�dJ�6�����kD�,�����^nc��Za��9k�BH(���D'�s+b�Vȕ� �ؚ+K-b�P��n�٦���i�D�6�@�pd�]t�dˋ�L׀T�� � ��j��b'��Sv:sL7�\n�M��l}�����������/߳�5|���y�q�R����̽�M�NN7�;�j�CӺ�1ć[�m&[�c�}=r�b3�e���d׺�g��ng�5��kVZN6�v48���\''�av.s�zs�,�f�/+?f!Ab�
WkU�imMї]ǻQ��
��b�vb�� �LAb_fcȘ�2���H���!���������4�߭�`:�`3��D�MG�m���Q�hY��� �Y��̣���g���W�������UU}�{���{���U_{�����c�]q�b=G]DqF1Lmz�ֶ�b]�_w~����k�6x��3��n.ŧm>9���g���!���X�l�}v; ��N�G��Lq`��r3�h�vmM#����y�nۉ�[;��<����ۺ�s��^���Ap��R�%��vF36XST�̶���{mkrf�=�E�<�ӎR�۝Y���v�vlm�M���v�� Q������B��e8��gl�V��%JKwVpy���0�]/7&�8ݞx3�2���o����ն�)a�u�&5[~� ��}ӿ��k�H8�,�qͺ�,�sٞ�kmB!���Ϳ��ck%>�H�b1�1c��j��gf��nkΟnV�uٽ�d�:�kV�����kT���?ɩ�7ʮ>S���>c6���4*�6��m�2���y�.xy(��:j:&�ɳ���[k?O&���6V�����e�p��2]Q
�_kg���!�k��]Ey�j�sR��9!l�WZ-U�^\���&���国���(�'�>y��UUR�R�m�ޣ#q����8����6��ikSf�^���Ԇ���Uݔ�S���p6s��)��L,�����-S����&�����<�\?]Hx�R�/W{B���,����٣�æ�9��k���������ͺ8�&�����͇<o���^%�s��'x�[co;�)'�^�6Q4	�O�J\�ًs1z�'���	�����IG4f��I�Ćc��������ϝb8�"=G]DqF1Lmjz��z��ʥ�9�T���>���pU~<>�����/p��sG!I�B�v���Ra�S�>՚��\�����ׄ){��a����mE����YUqH�QM*rrpĨ�Q4���s~)���Ζ��<��g�{���ٱ>�gߎ�fĠ�����.�c��y�|�6o���V��V8�:��h�8㈏Q�QDGQ��~6Q4R�55ك����1�������ת�E1��ޘQص�Қz����j�� ��t����-pKd�����zPUG.f,�/~���<>cޮÇN���t1��lS�^mן?y���Z8�ϫ������bpN�`h��zjj�1�̬�9�$���TCbp�x�_���H�X�����4��;aQ�c��Q8p�G�\=)���Mޣq��8��u�Dt���D0��0�����U��3.��7����s�|o�o�M������L��w̼emF���2��E�C8`�Yq0k\�,��9ɸ3�JgC��\�S���ns�uY�8My�s�&w;%�z�>
�� HR��6��Œ<���T����]���zv_YFo&U��/�}&��/?V�{����7�]\�yޙ7tg_yo��c�wѢ�lm��l?�~�GƦ���/����1���gR��M���<�Bq�M���=�OO^W�e̦�F�/
$�c�F���d�>���g&箵R��q�C�&��8H�GM�S���w۫�cvt��áO�xjl���G��l�Y6�%���>`iHLHVAji*BcLr��e�n�������K�j�\A�1(��I����|ʖefeɮ:{Xp��:t��:�#���1�ckSխ�;.�.猶ｒHĕ��/a���l��rx�U�]U�g��3�Fh�v��g��\?ŸZ�M��<_ҵ�%�|B��I�w��̭�o]<:s
8^���7�˒nf���yw�ێ]�×�k���i�r�r��m^�56�����?X�����Ҍ��Ohқ7�>ƍ2�Á�%�4j����� �럿jB�˩w���	�(!񇍜:~q�"4����G�)��F�SF�I�!���F��,aP�T	Y%�*���O��'O��I�sG5����IZ��ѳ��[��N�0��/��`��Gs��G�c���9���>�˭_u������<�[����lQ���n�(ޓ�/S�Uf�zO�g�UF��2�_�{��۝V��/��-��Q칌�OgA;�Ы���͘�!7���낌?@E�<B�ᦍ�U~zR�-���8�:����8��:�>DDu�Ŷ�=Z�<�N$<d9�TQ6p�?��ɖ�2�;;�>!��h���0���k�	���1YZ|��� FZ���͛�:���)���<��C���䙣��:	��OK)��A��u�f�)��=;:�`t��2���&�e��s���� �(�=��v��>4��d�:	�o]\,N�)m>����u0����'��Ki��n��>q��iu""��⍐�Q�=5,��T��q�8�Q���"ey0Bn�-�4ʱ\%n�Q!\�1"�F��MnI2��"T�F��Df�6� �q�<�$��!�A:PVH��Etn>� �����;�+��ow}��ox��cS�y�\�UYVL��C�b�X��,dnҹP�ɦ��
O��{��-g�)�B�����16ޭ[�
�nd��O��K�:}��;<HtJ(ku(�sZ�΅#)a��̞�:=��|���ٹJj!N yӇ��tNC|�0�_��eO��ִ#�ʯ2~�{E0��rL���%M������Y�~�+Y�诸�9��*�>�n�{�ǥ���	#��rb�&!��H�T}���fA�xH�lۻ��+�k��~������Z����zVed�$=�bQ��ߜ|�\|��E����DGQ��[jSխ��y�%V��ߚ����I$x����Q��͘�,�\�YR��ΐ��tه���[08oU��ߤ�8ᨓ�0��l�Z�*
�4�.�ܪ��յ:��s��1ohE��j���"ą�|�q������vv��:Du��9���{�>�觅p��ѠD��2�Ja����l���vE�2E����@��TX���S����y���O{$�T?8x�v{����e�g�����g\~q��GQH��!h��DDE�)DZDu�D|��8����#�Dq�[����z����H������DDm��㮢""#�:�-Du�E�"���q����Q�Z��E"#��"#H���D|���޽GȎ�m�h����6�m")�!H�#M-�|�4�uH���B#�X����1ZB#H����E��]u�|����4�#�Dq�)�R#1ű�����q��[�#�DR4�QDGP����o�W���8��9��6%����8�u�~E<�Cq��;N�ߓ����#���Ӕ�T����ߟf�c}CO�M53t�խ6e�]Z��v�1CD���[�y��|�uxw���9&���6��w���s[���N�9�|�0]�bͲ����7��kJ�eOt��h�4�㴩�5�f�>�y���Z�9s���Qߧ~��y��Ԝ��v����7@���WnenMԪ��>����=�ޟ?*���}�������U_{����}��|*�����[��m���u�|�h���F1M�OT���yW�UU��u�I0�>'L9��j4T��|��?:,,9:��xt�x'0����4y�]�쭸q�тj��B���"�"�8~?�ɇ/N��o7�nN�C��a��T��J���Zc<��z��c�+g�:S�ߥ��?M�&������C�u�~H�(�Uu!���Yf��q=W����~G�8���Z<xN��?�a,ÏL����Gr������aÆ�����U�Qb�����L�Z��7r�W]�m��C�E���J������µ���+�=����J>�#G����4O�5�OݒH��~:zl�j�G�sשw�J6p��Y�� {�x|If�JՉd�\��t����|o�m��'�<u����Zk������/|�o\(��,9�e�@Nk�<���8��8���Z:�>DDDF1M�M��O]���[IV{O9e�,���ƫ�*H����q3�+�+el�\	�+S�	B�(�h�U�)��9EEv�n�'!>��c\P�{w[��V���V�-ں��^���n�'�d�n������o�7T��SM��� $O�zU������0�bo�S��L��g	��{�٘Mda�b�N��M1�g�g��f��e�=�)�}ܸ��w�:�tV6T�]�$0��;�$N�N��+�{�f�B�������Y�^���͛S�|�-�kMk~��+�|�f1U��ѷK�n��֋k�N�����v�� Yf�J%+�z{���)���[����Ƹg��7OJ��""e����G\8ձ�-q����]��zv'�ql���ϭsz�4]
��<�V6�׮6�1�8�Z:�>DDDF1M�M��OQ߯;nQ�I@+v>D'�>\� 	U��,�Cf���6:y���$OΊ/���A����,'�Qg��mY��8N3�U�V�IgHo��a��5:`���:z�8~?|{�Qz6d��d���!s�~��J�n�$�7�s,�L:k:��Qj�����;/R�T9$���?Xs�f�`a�O�ɿ���V?�B������0s�y�1�Kq�:�"8���G]GȈ���)�)�=i��ԙʦ�M���37��l���\̕���� 7�����}��]9��4!}���b�f'є�ԡ�X~����>0O����%]�P�ǿ=��0>u�;n1�#oۛ��N�񸝆���x&�xl���l�(�@Ú�%�s�����h�w���x��ּ}�J�DI�J8fp���No�M�(���4f���o[����'��[�Oƈ��-�����|�h���6�6�L4h�4�?3l̠T�� !�UB�0󩊕���s���<�6S��&�.�æ�w�/u������M2r,���r�m9e��U^]�ɟo�.��w�jW���˲��	�~���r�950�>;�����{\2��
�|p���c�P��K?M�+ȟ&��=E��C���c��M&�ڇu���5	p�ˁ>�M��X�\�����+���� c���H<8r����m��]G|�h���"'��8B0��3u�t�Ire�d�����R�@�����Zۭ}���?}򯡻@0o��4�ҟo��]뮝Ć�f�֒�vp����ˑ�6���{flGl�n�w� �G_�綐9���ڬ��g3��;�_'��^�����ݾ��]x;���jDd�e���*���j�UDK��Ǜ��3����h��J��erdɼ�O���WM	�u�d�j�cd��=)�d��kj��iJ7�8O5?D��۩�bߴZ�����t{�6�k�����_-�����|��=[*R��͞�����4����`jl�ǇK�z�w���)�ɩ��GN�aL�#�ï�ӎ���]����<j{f�<u�.rbշI�}�L;.
j~4'!��k�j�iW�>����?6�o�G|�QH���DF1O��ޭ��Xɫ�I�	��/D8x��[�=0�C����f�׎j���0�����M�2z��DCA��3�M�j_�ٳS4<�R��{�n����KXh�ݓ�M��.��J>7����'I��y~8>5qGI����� �5�k���'ǈ@��;�W!z��ޚ�e�Q����
d0�BhϡRS~���{GZ4��kXO*�kO�#m�8�:㏑�R:�8"xDD���CfY�9	�;D
�
��Ъ ��ԁ��IEY��e��*�V(
J�֔�Z�[QDR�1��j�Kem����(�)F�C9�T7)M�0:hיB��;)�Xxd짾�U�d���D��ӡ���*�8y8h?qi�B�=E��j�V��]k�R��ۖʼ{�࿽�ꫛ�E�"a���F�/M0��}<0�Y}]�~a$	⠬ئ���u><�S��8h���!���L�n~����hߴ��ζ��+��Zq�~u�q��΢��Q�#���`�6h�5<w�Ȫ��L*�W���Ϊ����sr�؞{�3�fA�մ���C�g�����뙊8����*(7[���AurK.�GO8C�>,<�,��0ٚ��R��G�a����8NxrN���P�M����D��o^:V����؝<2�J~��6p��.b�6n}�!�h�ϰ�ч�ܥ��c6s�*���:�N1jR}Tm�=<���G����$HD�t�I	$����P����/��c��'�5{֥I�
"� �����坪�al
���D�D$6XC �$A� � Ȃ1� � ���
��AH�dA`�" ��$A"H�2 �	d�`�DAA`� Ȃ�"	H�"	`2DADA"	A�A�2 �dA`�DdD` �0A"2 ��2" �A `� �H�"	`�D2FDADA�@A��  �H�A��D � �� � �AA� �" �A ��22D`� � �A�� �$A$AD�D�(22 $A`�DA�� �DA` � �A#$` ��D �2 �
�DA� � ��0A#$H�" �DA"H��D2 �D2F  �1"d� �A$A"A��0A Ȃ$A��"2F �AdAH�H� ȂDA��22 �$A$AH�A"  Ȃ ȂDA�2��!�A�0A"A� �"DA�H�A� �� ��2 �� ���A�A"� �DA� �" �#" �#"$F"�dDA"0D`�" "�Ȉ"Ȉ"ȉda"Ȉ"Ȉ#""$a��D��"0+Y`�"�D�$aFDAFDH�H�AdD��A�dD��"D`�dD�"�"D`�#"0D#�D�Ȉ"�FDF �A@F� �2"�0FDA�"�#AF�FDA"0D��dDa�d"$F�"�2#"0D"0DdD��""�FDH��## D`�#D`�0�FDb�c `�� �#F"""#�22DDF" �A0��H�#FDH��"DH���"$" ��
��D��"D`���AF �#" ���FDA"$F$F�aȌ� ���#" �H#���"#"$aH�H��$D��"!" �"�D��0D���"�1�D`��H�"#"F�d� �AFFH$b$DFDA�`�H����2"2F�A �F���b �A� b"D� b""0DF"DD`�0�FȈ�#`�#A"#b �1F ��#(�A�ȃD`���"1FD#@a�"�H��D������Db ��DD��DF""�0�DdD�" ���2""�F��2"0��� �`�#"" �1FȈ��0DFFD`�#"" �dd""DdDF� �DA$#!��R�"��R"1H��!!��(�
1
Pb�Q�D)�U"�U�@)�Pb�T�1D�AFHA`A�AT�@XA�@(�@  2H��� @I ���d��%�hc "���Đd@� F$�Ȁ�Y@D�I ��@b �$� 1� �1A$$D�H�#�A#"�"F	��"�2�($`����Hȑ ��A���D"F	$bDH�A�DH���"$bDB0HDH����H�!!#��`��	�@H�"	� ��"FD�$R$H�"!�B$1"$@H�"	B"�"F	0H�A��Hȑ ��"D�"�L@�	���H�FD�$`��A"	#"D0H�F	"D ȑ0H�"$dH� � ȑ��H�"$H� �2! $dH�#�$D��$`�"FD���"D���H�A���H�H�"D���DB�Ĉ�2$D��!0H�FDH�FFD�!0H�"D��$dH�"	
�D �FD�H�$A"	 ���H�#"D$H�"D��$H�$A"D� � ��$dH�H��"	H�FD��#"D�$bD��$H�FD�A"D�$ ��"	Hȑ ���"D��H�FD ���H�F	H�"D�2$dH� ��	H�" �DA"@dA"	dA �H��LAH Ȃ �"$A��H ȂD  �  �$H�" �� �A$DAA� �"� �A""	`$A`�D$d �A""2DA� �D �"�$AdAA���"2 �A`�b ��PY" Ȃ$A�� ��@A"�0d �0AD� �d���Ab �H�(P`� ��$ �(FDd�AD� 0@c$���� �$b� ��d��b�b��BKDA��D� �FH0A�A��AD� � Ȃ �H��b �1�� �AA ��`� Ȁ�"A��b �d������c$A`�$A� �D�F�!d@` �1A"A���" �A"	c  � �A`�D �$A �0A"�" ��$A��2 ��" ��A� �AA"H� � �A �A� �DA"A�A�	`� �` �$DAD`�+�3�oT��u]M�9�R�^PL������H�!�.�Q����m>8����?g��2��[��@�Z�1���-�ƿ����9����!hk�K���)�ݦ���I�~���<M�j뻆|�����O���,���D��+9~ԡ�
"�矊��e�x��~t↥P  ���$DP<���h�=�kT����ǈ��K��V%4����������g?[�!�m�:�|Er�����:!$�J�j�G��D����:�P�ŅX�ɂ�~(�Oja�hF�Ӎ��y�w'/|/��r�nKB�Rd{�C�<kyF �+Mu*��DR�U�P(
"�
)"9�lE�Q@�U�VE��(P(4fS%+F�}Gm�����.�X�:��� � $�B�E� �EI �	 � @	 � %w�Pq�`�%���/����#������d��������]��C����������Q8�
J�ǵ|���.'�o��:\H�b�K���gqLDy���������KP�>�@�|�8�������'���= (��� 3%��Y~���Jtd`d{��`ǒ *('�@�o|����4�Z���r��Evɉ���B`�R��w��*  \ܴ�F��
�l�%C8
��Q��y�j�p7A�xca��%|R��z%/���:X��b���nJ�1���#��"�D��q$&χ��R��o���vz˄� 3�7;A;9-Q���W�z�y�ȟV����դ���(�GG�1���H)�P����yv	�YE@�EtT�X^��DP/}��߁��#-���Mg�9E�Kh��m�n(�0T�=�Fŀ�-		%��[�z�Ӫ��A���>��q��J�w��-����g�//DP"z���:^X�JD����v��ځ�ʎ�������1�"< HS�ʔ�LϿИ�k�6�� �1N��@��p ��������u2U  �
%������sR����ݔ.O��Nr��*�)��������H�
5���