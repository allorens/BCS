BZh91AY&SY���X߀`q���"� ����bG�}          =���
�-��(�F�@ ���Y(��3`ƌIDA�J45m�d CMm���������ʢ��Qf�[5�m,Z��M�ul*ƣR�f�m�,��-`�aQE���֔��j�h�ZJ��[m�-FhM&MlU$��ٶ��ƙ�V�UmC��P ��B�S#\nɲk4J��v�ٵ���8��P�Ym��k�յ��U��5aZ��m�a�ڤ�l�m�F�ka	Yi�mljVm�V���Y�I��   �����6�]�:i�Y��T(�ei'vve��1�*�ij�Sc[���S�:�܅*��ֻm��C�q�ؖef�$���x   ��A*(f��R��\ ("mv :6���(�v��u�AC�m�=��
����J�hR��{�=oj�Z�oyT��=�ֲT�F�h�j4�   s��zP���{��G���:^��P����^�S� ����=t頷g�|����<�AU{i��N��t=���ٷ��@{��G��z@���&a��Zf��l"U�  "y�^�1���})�>��mү;�^������=zP}L���B�������` �󞂪���W��(zf��ӷ��M4P�=�OL*��α5���Vd�
����Xx  �;Ά�@��G��*��E�_x��m��wm���V��y��Ԫ{ۥ*V����oC����t)J�6����A���۩Q����à��@��ڛD`���Ee��&� ����@
���
�ɽ�B���],�� .;�vU(��p�{h;�^����AJ���t���kZj*�tp����s#)��35��S6kX��A�  7������0 �A��@p�U@k� Gjwtݍfs�颅��(����v��86  Cvl�ն�I"�Y)[&7�  �Z��֔P;Us��� �;\���wt�� -G8 � ɴ ��9қ5�ժ�Pj՘R�U`�   �[� S�` h`(wc�T��n�\  wt�� �s� �� ���� Q� 
�ζ�+Q�Y��EKm�  ��;5 j\�V��&�	�J�W ���]� ;;m�Z�8+���(V�O�   R  ��� ʔ�F` �a0 "��b���#LCM �C&@"�����HM     ��@��J &���M0T@ߪ�O4�oP�(􇤇�1��M&d��E*4�F�    _��o.�7x�N�v<��:�x�k;�\jņ�q����.1��n��W�o�w9EQW�EO�D_��
�a�'���>���DW���c�>{�
�p>����{�|�pn���2s'0�����̜�̼�̜���s'2s'2s'0s'0�1�L<��<��<��<��<�30�s'2s'2s'2s��ə9��9��9���fy��y��9����d�N9��9��9��9��y��a�a�e�^a�3<Øy��9��9��9�nd�Nd�Na�Nd�Nd�&a�a�Na�Na�y�0s0s'2s0�'2g����y��9��9��&�a�e�Nd�Nd�i��9�a�d�d�N`�9��9��9����L��s�0�2s'0s'2s9�a�<�̜��<��<�'0�0�'0�2sf`�<��<��<�̜�͙9�2s'0s/0�0�L�0�0�2s'2s'4�̜�̜�̜�̜Û�3�0�e2��9���0����ȯ0 s 2��'0̠�*<�/2�̀�<ȏ2�0�̈� <�2���"<�2���*��/0+� �*���0��� �ʧ0�0�0���*��0̪s<�12�̪s*���2�̀�<�2)�
s,�09�Ne0�̪s"<§2�̠�(s
̂s(<§0�(�<ȇ2���"��2�� �<ʧ2̊s<ʧ0�̠�"�ȹ�9��0� � <�2#̠� <�0s
� �ȯ0��*s*<�2��(��2�̀�(<�0�̀�(��2��<�0�̪s(��0�̈���'23*���2)̀����(�(<�&e9�Lȧ2� �"<�0�̈�<��e9��2̪�"<�̈��2!0s
��y�S2*s"'2�aC�Ü���/0�s<ʏ2̃2�̠�̪�"��/2�0���(��/2̈���/0��S�@3 2�s0 s '2(f^dD̂�/0��
<ʯ2#�L	̪s
<¯0�s
���2̠�s ��/2̈�2s/2s�<Ùy��y��Y�`9��y��y���9��y��y��a�Ne�y���y��y��9��y�<�̼�̼��2�12�/2�'2�'2�$��̼�̼�̼��<��2s/0�̼�s̜�����<�̼��<�̜�̼��p�&a�Ne�Na�Na�Na�Ni��9��a��y��e�&y��9��y��y��3<˘y��y��9��`�e��N`9��3�fd9��d9�眳!�2���̼�̼��12s'0�A������=z�������e�6����jNU�͋�`��E��3�7E�]��ݷ.G{��fB����ƙ��*�RU�5������aB��j�燁Z�t7���j�j�A��o��)�Ҳ!��(M36Õ�樖J��ӏ&j�ĵkPb(��w{pnVVl�+�$x�(E7~���&:��Uf��B��-hQ0n���hr����$!�-�C ���uGAk�o��[�F.b�^�z�3[�Z2N����[	�7�9Z쿝�8��#ͬ���(\wu��0� f��׈'�[�#0�øV:�x2�Fµ�Q�QK�U�-�=���ڥ�,�N�J��ҽ+V�<�aVX��ِ�;P�%faR	�5D!9kS�ǡ P�cR�C��WY6�ck`f����3v2V�[J�@c��M�ѕz?�sۼ�(����8)�mf�(@��nn�M5|ys���<.�?��a���f����ή��or�TK�Ǌ9n���D4^ Tl��:�j��˃���j�yahUy�1>V��/�f��Ձ���	�X�hK7i�).˷ҩ+S*H����f�i�ȍ��̐dw�Yz�S+r�B��W����-UК� �At�mU�21�����O*t��8b��ls �
[�R�-0���U��k`|Vٽw�kY`2ڕ�f�)1X�Q�xR��B��Gn���4�9l�`sr5T����0ͼq�1�����H+^AKsq�5vڲ附�g[�cJ�ݸ֋lĎ�6��t(Z���%d�&���WBMgG���`Ԩ��[7[��f��y
���6�/�V,��߂Y1�i��3FR��puf�;�3]:!4��X�#]ʨ�� �\*/��4-2�7E���әϞ)%�)`�a�h�mQ%�y�b�on���o����-%x!�1ndoF
t�H�5�
0�n�[��(�#uA,f�W�ֵ@��O�}�3B�b,�ÑӬW,�����n����ۇk6h�G$�i�*��YM�Uxw#�s��`B��zp�8�!���fU�[w��jY����V����K�)I\v���
Yu����k�V"��3�m)�(nՠ��_چ���$m�b00�L]���V�["2j�6n,/4'�u�����U����6����F���J[PIX�T>�qe"n��Yo0�X�*�Jf��wԩ�wt�2�A�E�h�6��)f�e9+ub�AV[ʹ����.��T�7CҚ�m	��5y�N�X@�Z,��T�E�L���^���ʹ"$[���إ7yG#ۆ�؋�;�+J��l*�6�ت-:�*�g��V�:6A�*0��2�%���S��˗�i֍���X�A��̡�"�El�Cf`*e�,l�/�!ә��C�=�3)DG�/3k�%�K9DD��L��h��YwR��ff](��C݂��L9p�C��C#X/u�$k6Pb��j�-엪3N��H��^�#;�k��v�z�3l����WC���7�X//�s%(S������6�Vm�4 ��G�N�6^bɍ��m�	d��`���>���dK�%;%̘q��gtR&�!�2�m�^#5�ᝇ9X������p^�d"B�Ӡ�mJz�؁�H:i���z1�H^�woHL��y�mLm��N�ūb5n��!"O)ӊ��{VLdm2@}����e�h!��gm�G���m�&���P�Fe̦mk��ҥse���2]L��ܩ�(M7	V��c�n:���ȷc�5���#�a�Ö�;@�yYGj!ٓL�{2�<���ݍڗ5i�o6�a�d�HјQ�#pMZ5����ki&i�˫���3Å=ۗM�m%.�B\�h.�=h^k%�IqR4ü7 ��`0Pw"1�i,�λ����f��3h���9��-Z���V�h)�G��J�4�=����NoZ�����7����a�A٘�Q���́�F�Z�.�62��e)�5=��Y�!���h�2��63u�k B��N@�]�U�hc0Qŀn	W�q�Q5��O]'�'�7�h�̮#�G&�z�^�􉈊 +���J�����ݐ}.���KqfJ+�1fv\�
ǇV��)�/*�ǨO������;[v��fh��tI$�扷.wS4Sz� �2�f|�o4��d�=�x�{sR�sw)$�M���[ ����.�/u�[Y�a���7%@�Hss	W�o2n���Ѳ�ZTmc��"��ĵ1��g��F�
��l�J(&��lZb�IKܺ$EFP�����7y�q򎕒f�zQ�JcR
�hvI?��{�1-֞�!X6�kI�b�w�-<�[n �۽
����M�YU��F�T�e&�Pt�V�&,�������NYG ?<�c�cM�Q��$ˉ������b�^fM�iUb���q^�+7ຝ�A4�a
�h:F�f�h̫��vU��rˢ"�j�n�=L����5�y��S4�{bZ�����Y1F�"�QnYzv�
ɷ�0K��Q�n��;�ê�6�%2M�p嶅��G���Z�˽��܌������@~x�'e�m���];L�$#�Pxj�]Э���]Mw����f�
-�J�W-���6,���଀�d�Mݔt�c�$@�X���d^�&�Tn�р�XXF�?B�42�J��Ɋ��5t���Q`p�`����XgG2icc����-ҵ3I"i��Ro��ƣէnD��"��k!��ۗdk���t��[Sf��"Q)qD��?U�u��2�0R�z�w���˙se���;��hUA�*2�ŹlfQ�-ok%�)#R�Mqj�5���wI�L�0ƌS.�X��J�d���Ԫ*L��NE�b�^cЌ���Nq��lT��ǘ��� �t+y��KZ�����/b�lZ�7�i�6x���s�x�-��K�3����>�8n��m��	$3DdL� �ڻ��om�+7e䵪�P|�(�[c�Y�
)�D˒

�m����&f�����P��C��S�.��=�ؽi[�Z�P�a���/!�E������#��"�Ѵ�Xs�ae�	���RV���h�!�YN[��4'�+Jk̅���7�崬7-�1Ӗf��Ů��̠{J�1�Y�"ݭ�e庉���­��Q��{)U��͍��C�c��0��5��]' p�?���H���淍���6���bcZ�b׵x-��N*�2Uֲ�Ǔ\#Vqd.�K�>Ii�U�2Y�-��!x��X7+]�D�>����H����rH��aTݼwL�1���a��N��d�U;��
	jR�V�Z���7��+˾<��篒	�X�+]��P�#Vjܓ���n��u�@���Ӹi�/�TeQ�X��F;V9h۪����B�ETv:�r��)&i�hpj�?,�@�Z�^j��;�*n�"a��2�C�]nU�-v��5�c$�51��lS�����bF%�l�2LЙ���`�8�J1�*�i�ķkTwrڄ�a�&,�2�U
9����R�#�7�"�)I72ј���Cye���M�T�x亽��r�jK!K�NED8��6�%�;��7MŮ�H3V�nd8)�o�k�ma�wm�w��x�#��XOqA[B-���wb��H��-�م�͙�G�*�P���nɬy�cҘCÁ=I�ˡ�	��rKV`����]k"x���s�(Y�,�!�f���h6�G5��R��0�D%ݼ�X0�T��tX������k#3h�t*nU�����[Ɂ�)Hh��r��а3z�X�YChFt��y��	s�p���.LhZ7�0M[�i��E�7i�Z7>�1d�Ln�Z�S�����ե�v-���O�[� r�Uʰ��̢�Q��X1�%�n�/�`M�"��eC���L�d�kC�x.ɷxm�����$jV�Rl+C��Z����j<F�q&���2�ۤ�).jҨ&<��0�Z����m��e���wu��J��xȨ�Ye�E�� {�,��8�KU5�ӷ��n]�j�~�6�.`��&�ث����Y��Feڤ,(h�.�Q�˭�n�Ȱ	�]�[2����U+(\S^���ȭ䢥���r|Ξs�urd��{������Է���B2�Vc5F�Q�mRܷV��ؤ�6�H���K�B�eە��p⥉]b��@Ze�إԭӆ:8��/vMܘ.�
�	��+EP�7NJ�6�whP.�m���B`��J:���Y�e+[�]$�AM�SX�k3�jf�ܩG,<�z+L0v��60��Qv4�X8+��j�ʣ�0ʦ�te��ѸD�"}�I.�5�v�M;e'я+�R*1�MmGJXD<%ڨ�EawE�P��L�n�Ķ�7��5q�&S!m�ǽ��7E����T����u���Jp��he��Bb�0D���im���[�R�ҁ�b����"ŷؗ��(�:á��*��<u�,W�40��f⼹��SwN�`*5f��p��<�ř�\eaT�T�kjn�w�	��9�ޝ���#�0���gdH����'���!���6��vqMj$�>ɖ�����͒��FX�jBN^��ڛ4-�{&�j�-��­�X!"����0K�kÓІc�)EW�����oBU�e��%�&U#l�kE'��Y�hG"���ʺ9n&�2A�ˉukn�T��.m����^����_�̈��^A$n�wY�uE�M!�k�@qdj������� ��x���hP.�x�]�F�2��D��֎7{lme8\1p��#jVf�fc�+2���.��ȱ�[�/a�0��T`�*�L'e���X���^�x�ŗ�Y��ØP�����DZۏ~�2�M�&��˅�Ynl�KU�C�����1����{@��E:r�ܩY�i���ESV\5A���z&�VٽS�xDʰ�Y��ѧ�6Uɚ���wY��-6
F0a�Q���:�,�$���ywt�m�N����V���K6BnۗG]�Ly�c�M�n��YD��h�q�{6�kܼ{�(�E#��AT[w%@�T/^@T ���	���;/	�uw����!"�F��v$��.��cw�S�	�,���1�y�҈�ݎlx�[sk;��7��kk{;�V��V�zR�2��D�6M���rƭ���dn:X�aI6�{�QGS�3%Y�M��u��u<��[�	(��U�HG�����m:ʂ�B�R��gH��`�P�w��5���I�t�U�Pν(���W�>�O�lkkC����ܬ�9uC�����jʵ���]D���Ư*^�5*�pT�������D��j�[S4H0�g~e(�v!��@����ly*ɬ�-��Ne&h����t�+M*�m�tU�n�in]|jnT���G]Uo�R}i>�mX6�n���ѠEÏ�z�Zʓ��%�a�kytk2%���Cq�$0vJ��6�PY�'j[Q��ёaT�^�1��kg1��]�Ow��s�P�-|��wZ��ti��?n2c)`sR�Wc�Sd�KϵV]�C�0�ɶ�A,:�E�U��w��oٵ(��r�XfmI5A�X�
���7 ��Ml u��j��%37[��E�n��r�ԖZ
V��5r�!x��VI,Si�j��sRXÐ��Qq�c��L̓7pͽ����'"b�qoY���GT��ۭ��2�B����*�,aKv��3o[�z�8%'*l.�`ݼ8Vw�k!�w�E�h�Ÿ�jZ�.�[XR� ��Xٺ�R�ڍ#40h��*��d���S&FN���J�
���z2X.�McE�8���1ϪnдƩ��6�ɻ�:!�8�fs�AT������J��O�Dڹ�|�E�6��ku�d�֠�l��l���kZ�L���	���$�"���m��Ynۗ�!��ecUl�
���x�6�^�6<YuN�Ec6��
i�3c���yfm魻�1,�Wklm7��xi��5�S[J���d@�˻&�YSdZ� ��\܏M��t�~̢��q�[/Kw�01z+�̻�'�1�Y/ dGq%�6�#�e���_����!�-�5�z��F�r��DB�̞7�;9R��OnR��E��y��R�o��D��i̦F�'�|�E�W����ü��6�=�7���i��n����%�}�{XrY�S� W�`O/q�(d�+.pw,�NwI��}�`��]u�����K;1K�/���9\h�Я���1N����sL�H��Xư�-��6�F��8yn�zi,�岭�˷Y�.����i$��?=�6b��ˠ���](�ienM�qt��ahJd��Z�i
���s��s%��R�T*����M���GU�!�g������s��9) � #��^��I̖��ʛ��P��pی�Ѯ�۵�s6H�]�`�S$:x��)�8CR=�!Tv��̦EE���E�������#*"0%��=y�xh�T%���ul�fu�7Eܭ����f�`�TA�-��n�����R.=!n�]!�nV���4ʹV�cm�n2�Ӄq,�a��/GP 4���s:3tV�d��އddҬ2V+�
R�e�ۖ�GS��)��7��h�V3�n<�B.���]f���NfV����m�fk�X��Ui)P����ۜM�ĳx�64dw˹����j��á�sg�/N"������yj*�ܙH��Q�0G��L��\nM!stg�M*��~Ys.ؼ�B[tR+�Z��^k`һN��Z.����������KT��o"�Nǈ�3{�=慞(�b�X�������ʘX��+X�hn8H|f�{�\e!�1��ɹPzY�p�;.l����d�H����<|e�՝}��xQ���Y�Yc�!��!Pu��A:J����5��[�-��VCO;��Ճ�{�8}��-�`?��/�'�f�FE�↛�sމ��2d��M�m]�ic���[vO�o�R�լ�OZ�f���6��K{(�Quɕ̄-�\�l����u�8�th�̙+��
X��R`�C���N�2�"��c��U��w��(������=�)jna����o!m�l�4x`l\���p��ԍ�7s�ɴ(�'U�Hd׬jt�^���f�:��k��ٕP�{]�Y KH5��BM��[I����s�R����
�;=Zۥ�Cd��ip<���sU����̥sfqh*�|�8��pt�Ӻ��]a�7R��ݺ5:��(jd�h�f�A^gRڝ�e�$�9X�WaӸo�q켘�4i��XK�vs}6_RW�v9Q���}ce\|	�w>��n���c=�t��r���G�	k�I
z܂�n�]l4�<Eas������\y���l��U]y�D�1z�/Uwb����5+��'S���kQ�w�&�lUƅ�4��ZA\���Um�T�Xu�/4��c69�Qcy�z���n��澁��t���bc��ׁ:%�Ӭ��V���FR�e[3X�����:�5$�ٯ�Sw�M�7�Ed�[Yy�Kgnj@V�&��*�CE������6���V7�����c���:��s��n^C��.�[ʀ����S�cꕁU���}�^�:z�-�#�y��F�'��&��2>�КWu�{ �u�X�Z �0�T�o�!���D���9�
��}�n;����!�i�f����ͫ���9VpFa�u���yn3��ϗ#��M䕷g��Jg!��U�n��PG+V_^jm�:[�-)�6]��M�p�g){�_l�b��v�
���'X��7)���M��gD-�p����Â�%%/���2�d�c)�8Hl�Ų1�hU��n.w��_�R��$�}�;�N�����'cza2�j6�����8(��qu�o��lU�Ay�:Ru���n���!��z;�eˢd�Gc�gwT���{��F)jY�ϵw@/bƫ~8���`42րD�	���B���0���hSh!��.�vg���-�&�����kR�2�vsF�!G�T��7�)R{`���ne���a�vu�$�U1�$���z9"��Z��<V�Z��V�2�}�xk��E�`�g�wGwWw�G`�Z�����vh�aX|/vΥ���y�G�'^y���n����N�`�z�Z�5f\`��@^C{S�}�*�4������ҙ��;�>�Vݭ���Үx&N����a>n'���F��6��;��ySg4T�Ht&�Ү^ŧq�ΌzNJ���81�(��vDGF�9vze�q��hYQ�k�����%:X�:�@]��K�fL���Z�v/��e���C��5�rR�����Zefm�$���;�Iz=Pu������6������Y�J��2���f�r�,^r�c�A����
!�	+X������˧�H�8#�y��w[�k[�Z�,X���1��wfh���ϭ��<��w�#w0̖]0���K��]�/gb襡�Y������Q�=�~�[Z��>堽�vq��}sx�\Ku��E�o��`�MP}eX��mY�d���>���Ų*���	�./q%9�� "�sCIl�Σ�«�%9�:�#�X���^���̷.�n\n�a{�[���`@JH9ӶĈ��oN;���f�fVcq�̏3�#)���7NF8�N��Ԓ��ڵP�#�1&���{�Z�W���	<ː��+;9X[Ӧ���¯]��^��4n����=�ec���L�IW��\V����q�Th�g7V�Q��I��y���(�3!u�����3�7�C��s�.{ܶ�{~B,�-�@aTO���^�y}��֡�IrS^8ėV�iڣu���|�@-��.��
��3�l�n�R΢s^�H(Ra�-ؓ�����a�Ў�b�<ՠ��f�+��Z(��D�N�S��:�����n�_)��밾l�:�jr��
�Ɋa�&�p�y�x��F8��l�I�=V�F�a�yn�kI�ݢ�q�vW3���E6Y]t�J4����ő�-Xz��f� &Hz�2�VU�f5S%�β�"��˒[�}�A�7pF������_ic��Y��۝A�O��"�CZ���T��1l�E`z�r^�<㧺��K�@�wC�����+A�@��
�����x�
p
�S��/w
{bH��ZDꓴ\z�������X��v*��Tr�s] �U�2a�F*.����]��b�]k�t���ntO]���wd�Nt͘�{�G)�V��7jN��ى��[l���ڱ!p+�q6!FcZ�m�k/'\�H�dC8����ՊdM7��ܺx��w�4�98�Й4��*ٕ���/Xt4R�
JR��s(�ך��LZ�ln�f�s�#�E>5Օ|,�7X��C�>�X\|N�W7����	�b䣴��>�,�kc:ᢶ��[��(��-.��P\7O�V.�bݴ&K�5���w�S�ڸ�^�8?�G�]V���p�Kx���v���E_�M�mʜ��9?�]�_�m�W20-�۽������Ր�ڵRؠ��ͨ��~w���n>O����c�O+�s���ܲ�{Y5spy],�J������z�{T�4��Ś�+�2��'��;P��_��]p�#�s$�8'N6m�{ܛ즸"��T�A�\�2��ݛ�6��R�'��|`u�]�M��P��.�4�O�>�]����GW�,�K��l�-�Pu��(.��J���K��EI�Ao\5ǯ5f�ʔ�F�h3�d����T��sJ�!f�М�
�.c�ڼ����v)�6ۖx`w����<�D9I��WB1nj\�x���\�f�S�4b�y@��'=�E��9�N�3C�h�tAWbZy���Y�3@w%�7T�c�h�z�V���7F��{���!%f)AHI���s��B��hq	�т�!���vd����_)sD�q[o���[�/_7���Z�t����ǋ�tɒ��<@�0���l]�m���n��;���;��z�z��'�<u{�d��`95T+���jי�#�ּ@.��skX�E�Һ����^3W�$:ژ���������v��g[��\���6�u�YH�[�4�f���Kҭ�WkxLG{�Tz�}�z�_	2��2r,�q�-Gr_Vir���sap�ğ%�^��(6��7M��fI}�q$���/.]3��Z�㩽i�mhT��zg��yg�W^w	��ٺ����q
��-:ف�MbuԁD{�{i����݅Y$��t��W�)f��II������dYa�[2�������/c;}}Rr��7�o5�9�8j
�:��:����k��U*=�K�1ϔ����)�Y��b��f�2Ꮮ'��N=��K�%��[<f����T|X��N�9]��s(e,�VB��u$�:����ۮtm�0	�m<�r�[�w��.����8���9�>�4��\ϹP�02�/�i;®Wv!��:tv.�;Bv+!X9��t�~V����Y�o���k2	niH�̇C��rt��+jm�u/_l=�Bi�l����[��!̎9�N�u��ҕ�l�1��#� ��_F��Ws��i�#c�oR��w�
5kxlq�ΧqC�)�c������\л�1�u ��.sV	�w]I���"�b�{]*�M���Q�[�E4�Hz���(���0�u�C��a[��Q[�3j���?q�굝,��Ʋ6ia�l���1�9t���L��\�Egfã��M.����]�l�)�P�=�g].'H1X0��'Ne^�,F闙O_ljH�(E0zi�ݔ���^��s��+E�qP�=�[��p{q}��G�c���A��:���:�.�Z��mm@""�H�)Bh����Xq�G
6J�2��Ӳ����59"��;$�1>0q�Z7U|4}\"��ym�\��&�&etk7VZ1�}�x'��SS`M��y��k��V�djU�X�����1blX��,o�m�5�u�A�ê��'�B*��'r�U$4��S�Sj�� ����_s�I���k��m��G�;�Z���fJs ��hCr�Q�<����7�Ӣꔂ�"q��S4f
�
�i^���l�/>"gq`�]ϊ�1E�&fʰNeD-r)�M����7��W�&v����g\٤�"v��Þ��ÊA��i�K���۬�>�:��-��ĺ�2��t��y�͸�->��̭�P:�,��PG��-nX�����e��7�rC6����]`S]�6vf��#��S���CZZ(�^����T�}&��$�F��d��^��5l&���Y�	���&1��V��m�9�=�PA_*O��Y%N�[�7���.yA��qk��P�F#�uů>�>y�ۿ�X��|�%�F&AOB�Sgn��0�@�#z�`�������!���p62��k9V�.��XbjS!�瘳%�m�Y��Wo��7��씲r�tJvE�;g�Z�M�k1�?Y%"-��aζ�h�Ta�R�4�V�;k���0�X��`��-�uא\��*f�3y�Y���/�_\֋l���r�r��~V����-�����t
��ɋܨM71���*�E�ھI&�e���m�s;���k��ޗv�D�ì�.
#e*�@R�2�dT�Kx�m�z�ֵ]���+@�$孬���,�s+Tޑ�ƺ=��K���4S�(�'$��b���0���Ѣˣ����[��a~{�n�W�ֱfc��=��g��KI=���;ui.�Κ�d,7r=�g2ݫ�t!�[��N�YN�T����"EWyv�J,p����r�� L��3{T��\`���$xu#ۮu��s�Q^
ݽ�)�T�X���2:ǌX�$Q�x�[ǫgm���$Y����usT;�NG��Ց`�ڱ�9����^�ԙٍHk�#�׃��G;�D����:ÍFT�K��l�yZx�����/��M�;���w�u�af��q��	-���өY��m�
luŢ����JSh����9-`�t�+c)����`S�oS5c��zk^X�Y����j�G�� W ��^^��E�\:3�M�界ٛ���l��#Bh�x��y�Eɺa[��9o�3�XOQ߽"z:���VNq+P�v�G%��jr�uS�pK�"��z�T���*���6ۤ��Ux�y���/ Z{-���0���@c{8��Uن��@g��u��V�y5�
�0Y�x�������V��x�×�p�[�Sw��s>���f�u�W��@��k_^M�r.�S�����aQ���3D��Қ����MO���V�Ҿ�yˮ(/��K�s����U�3N���w���Z8�v8����B���o��3�[\�p�9X&�d@��j�X�;R�>������T�ZPu�Z۾-�8��qt�"���V�WA]�,��|R���U0/��!Р �,��a�d-t%�68V�3��)F!;J^u��ow�;��oC�'v�Lr^(�<��a_m�߻�Zॻ���������K��rlF>���<��X~C31���Cm�������b��+,�h��f����*zk��^]9��{aEJ�������YZm�#
9�>�J�+��-���5F���{Co7���%;�:Nip��mw�EG-�|�d��S�>GP�v��"�ʊi�G�����ʲ�J:27��^��
�Rq祗R��� ��u@x��_k�@�/��m��Y������D�iV���,ݭ��Ӆ�wfk��=]����q��>͎�ƲƸk�[�1��BsN�%�ۈ:�{v��0�����U�,�%M>]A�gVe[U&�&�8�Φ�Kh��^Yݼ{�-[�ls��n�br]��a����m�ə��	x�˼$<l��*�R踃�(�%��V�C����n��\ʩ&>ʍ!87$�'l�;�8������JW,u'��oa���o_���I�$�>{5;���t��c�0�n�{��a��"U/Lu7)g$�IK�:���>r��Y�ΎPђ��r��d�)Bm꼝�{B�I^v�ٻݽէ�*@�3� N �rB�*3�@�qST5�Q<��4A�Ԅ$QrpH	&R��c m�5 ���NN:%�&�.�YJl �FF����]J�[g$Ug��}*�t)2@��i1i	E���[�HbC�*�Ze ������h&�J�>�1� ���S�h�[��Av$T� �E������#Re��Ԋ�m]]B:�2��Ѳ�<ӭ�)T
R��U�f�m�v�*"�	�FXs�a_��B��7�a�@��b2�l��"��T�$a ��Ǡ�(
�""��!j0��4ap`���#aj�nOާr�6�o�I��:���WI[�~_~i��A;-&	�	��d_�$e$���uRQ�|H_�D���-�M�@ƋL��*L�&#*�!2YM��
ؤ'̣ʹD�wm�(��8I�A���&�T� ԁ�.��Q�$G��Ge�h�AKTUE#$��("K8r��U�#E��jM�S�bU�0�؉Ch�DH^l3�?�~�>i����Ӷw��DAG���=�Q
�0g�oW��"
?���ۼ5������᱿����3α�����8#����4�Sȵi{yN����WP9!چ�9�R�$��l�Z/���A�|;�j�����%r���>`�`��a��"l��<u�'s���ou�:�e�V_eU��3c�q�X3U�\�vm����n�L���vh�&�����&�-@ǘt	��H[�b�q�b������Yt�����}���4mv�w�yTNie^��,��(+�cm��:�:��Ŝ.����z��Z)9�i�w>�O{en�z���lw'6%�Fh:�ˌpj��.��ܬ������8'�#K����2P�om��)�;9շ�gYO�f�F�Vk��nR�B|�Z�N��6�*����̌@�s_n���t,��u�����ƚid��F��$��(䕬����k��*-6����0ڍ��'�椲����t,՝�e�\�u�¥�Ne��ͥ(Vp���d�6�rH-��0^��ڙv;/f�����^
����
_[hQyJt���$��fF,��ea.�T#yլ�R��p��x��kz�E"%tr�-�jP���
�bж����Yި�Іq��-,J���;'d`�AЧ�8u6��V�w�ﻡ��v�S.��g�����������8ff�噝������ٙ�����Y�3333:a�����3�g���ٙ�ݙ����333=33�fffza�����3Ӗgffxffw�333338fffxffwfg,��ӧ�N�:vt���,�����3�sɽ�s��5�����[�{j�V�2��b'��ˬ�7*2�)�ӷy�g+���tm�z�2 ��q�޻ǳ�	���� �MXpy�ȷ�]:p�W��$�	��2;wLVD�[n�po/�d�F
�ޫ���E5�͓Mvi&���l��#�ͥ�c��>�¥՝�E�ɳ�vZ�D~���a�:�Fa��{2��Ӣ�J�_��/5+�''bںt*"��z��9u�7-Ƿ7�J��Jq�RV�0T��[P�΂�rݠ>�N�'�tQOT�tj��b�n�{vV�P�C*Z;�Hv5��9b���z(X�=�����Vؖ��t�f&�ü�=X�}�P�̻��2�Û\gFJw�H}�ف��=��Z��b:��>ݎR��t�|������]�0��]��UR[��Zv�#t��l�+�\�F�5��;M�AԖdj�[����S�V�8.��GcY�^�|��3�R�U���Gf��\�@�z�a�R:+��j��:� kGO�����ͮKm^p�wXֳ�A
��K�4���3�B�"��b�	������ĭ�G�t0gP�k.ց֦���I�*�:���k2^��~��R»���.6��&k{�0쓤-AZk�bOɤ͎�*V�[��>ߛ�9fffg�g���Θffffzfr��������33�33<33�fffza�ffzfr������噙��Y�ٙ��ᙙݙ�ٙ���fffg�g#33�333��Y���3�,����:vt�ӧL���噙��>�O����}>߇˕g&�>JM��]�2�1�jv���;Ю�M�@�c^7�ڝ]��qHov���1'ea��ާ����ؾ�yܒz{$tT���s-��:���R�
��mJ�M�X,�U	�5�u�[۫��g$�F�A���Kf\.�2g�N!X'T��e��<��E���f˟q�Y��5"h�	�mʼ�}\�^�*�ڻ��;V�u��"J� ��#&8���ĥ\���x�oM7F��1�يH�˼��Q��*3c*v��M��uv��}mmJ��^��llP�4�\�QV,W�o#�2�{��KXG��c)5X��"�ɹUXl9�jJ^Y�\x�s���}�a�kdB�ve��_���h�ɦ�}��6��R��]�-�W���o,����a��*�;3fʲs�^VT�p(Z�f���j��V�^�����ǁ�n��4N)����:����Q���Puk����-��(-��*QˍQ����2�Ո����3lb��s����B2����=�O,�`�K� R���V��h:�<�|�x�Rə(+ݤ�]��Ǘ��/V.�����3�+��:1�Z���[ �M�ʚA�t�D��W�6�U-S��Uu�۷��`m��C��߷���>�_����}>���ٙ�ݙ����333=0����Ι�333<�3�333�33�3�g,���L�����0������33333�p����,����Y���鐙���Y�ٙ��333���Ν:t:t�Ӧffa�ٙ��w��|��e��l�u<ժ�����
i[�X^��z�^����^]��AԌ���Q��}R�UW";��)�����D:�Z�71�X���+$����LS)?�VE���*6�0�M]wW�9�7r:W�����_v�Ŕހ#��t�x�̃�wi[�@����)�ځ�Q��ݧ/euw 'ݭ�Bծ��IN�<$��J���{q��ci3y�&��c*([��rWU��4�]�`�bݑ؜�bwN�R�R�%�^ӑp�>�b���f�)���ݮĵ �XZ������g���sU�.��W�
v��-YР��RĀH�����q�	�k�7��[����9��ї�BuȬdeX�Z�u�j�VggeKR�;�����νAـ�U���]�����'��7�V�oD=��e)K��=8��\�$�k4̬'��]�\���NPd�C�q$#wWS�x������[�
yd��P��Y7U�s�=�'V����K�9�c���W�+V��B@�g�)���@u�Fa�f�F;e�"3n&��0�̨�Pa�f7Y���<���V��Np֘������8��,1:�:CS	n?�u*lf�;$��9 �?, ]wsz���E�B%Y*�eP�B[����M2��]�	�Kd0k��tG�0H�f]X傊�y�=����)S!O��GL��x(�+V��n$�<��z�L����]��OyԜN���h��̼w*:�G��ٶ�u���P`����+d�2�Δ��8t�h�U�e�W��=K���H󴎻x�K�i���=7��.KJ���P�a������B�k�$8U�r<V�3�}O�^A -aΝf��b�ڊ+`��n��zN�����RڐI�wr�z��A�1����t+��emTl������m>eS�7Z�_p�?a�~��ȧ2f͊��4�|1���d�`9���r}��v�� c15��||9W^<���{t����Xve-�n�=�:�j��۹�4]
�c�\�5HpF�o9Va�U��_07��UHJ��p(��8f��kHYU(��o��R��}�b��[+5լ/;(���}�,ۭPQ)�\��،�#���%}�B�EW��"�xy�-Qb���i�m���n�!k��h�,s�)tc*�aWHTxWʓh�3M=X��S��/�2��������F[f�i�'�Zv�e�vc�9�0)�VnT[PK�*����ֽhV���j��=)��}#���U9&;�hf�9��j�m_�}�P�f�C���tL�A��1W&�yq���Rg���@��Fk����FRb�q!@M��;���
{%�[g�f��)�{�ݘ�r�}���d��E*|)7{2���8I ��2�v��r�:&��x�*�\�ߪ��&�+T�d�2u�g	ޫ�4���(�$\��J�Sk	q�F��V�	����Z��U{�=��PY-]�u�h�T�@�H0sx9�f�N;�0��8|к�O˷��t]8�L2P��`ن���f}o;�N7����D�gng�[ރ3yU�j6)η��;%%�˺M7�J_}3f��}*�K��	��!1T{u*AW�|F%څ1��� %V݁j�$����a^)�CX�[�+C����e!Xپ:6�|v�,)l���|��[���:��šE>�OO*m�X�0�Ðc���m�}KF�����ҏb�)��8����]����.rQ�e2�_�v͖ �w{ff��Dh\�-uԪ���<DT�Ɖ5�� ��'�̓��ǿQU)��𼇄ܝ�c�o�kl%x��'��u}�J�v���
3�P�Y�R,�M��чx���̫5¯����Q�io�C��+;J8�\9�9�������o�dZыF�O腲�^@�h�F݌�Z^�JKx(�3`Ӷ�m���](�͟8�f�>w�M�]_]f�sz.(��,��hw��v$�غ��Mic�N���٩�xj��wbs�&ݼxn��q�6��r�I�_ӻ�z8�F��z�G-��+��J�[9�5"'*䅆�Ud�{"���拹�>z�ES%�D�u`1�[�L���	vJ�h*E#r��,Zy�*o33��MP���=�+R��
ם��H�SZ�ڬ��{�*���uZO2��q�r�rgA�R�wwG��kD�3��z4GG�f����S����=�������!m���sD�u�D���f��;)*�b�հ���n�����6x�U�34�56�o�_J"�im�(�0J)����o���RP;ގ�QR��B֬q�Vd�ǇQ��e$�R�;ni����K�E@�ST;H�Iٓ�j/��lLl����Z/��U�,`Ӷ��\���Q<͟��7X�^��!<�2I(���i�6�����$[�S\6U3ǉ�}Ō:U8PN�}�Q-}�w����XN�Fu
�
�33+�v��
)�m$#{6���3LXz0^�[��4��5�F��H��f�t�}������N �Nu�M'�<�z��p����[L� �v�t��32��a�o-�.�<��V����\ �F ����E_h!�yX��xH��ݴrF��T3G(vL���L�w����4A8�K���n���mG���O�.k��d�
��XR�lЦjw�Y�E�u���j����ǚщf!��=בnV���6�k��5��ڼ q�޴�G��Ô]�E���e�.�i�h���6�ۭ�i&�k���S����\�4J�%��ɋM ���x�2#!�&+ODѢ��T̡y�NO	��]��QU���]���B~��RS���E�ƹ��Z���z��G�㻽�,��LO!_U_bL]=l;"���y��6�D�F�p�|�oܰ�t��]I#TD3/�Y5W�Nn���c��� �:U5���eت�s�ˆ���fb}7�PWm�N�%Ʌ)* �9}�(w.*�eT���q=
",�0у^��]rb�`lմ�Jx��˔�yf���B�l�}��qL�Xq�PN����;!ڑ\�5���y۰��F#�Ō��[���f.��!���ڋi���K3p��z,6k/�J�
X|t�͸0|FՆ3P;�++�����ɖ~ŕ7Ǧr����9YeZ��eX�^s]�ʸ�5�Y���_c��=Ӹ�MM|���)V\"��t�]vԜ*uNP��.�%oYc.�P�"a�a#��:�
�M �*E\����54�-9�w�7���j��8�D;Ƕ�\�oE���5�vb��D���0�y�����Ȋ��=Fcc3����2o`����
��=nd��t�_H��fIw�AL<�����i�uI�P�A�.�t�Bkv�C�3�r��v^=nu���*�0��q��#����N���ǭڭ]q��U��J�ݎ�mh[�����)�oV�w���\���fk��N6	�W�B��#��!��z�3�P�C�3V>9;�*��V�;R_@é��uڬaV�woN����Y����){NeL�,J�Ov�l^n�:!����:�Տ*�_WD1�N5��5vn��9,��!�b'�[Q�2کD�[�D�����lVQ�Mt���ܷ���%��}�j���Ry�XX��l��΁��8z�.��V0�e�ǘn�ϱ��n�^�KP�aNQ�_'CU��%�1[(�3��,��"�t�^-/> ���X88*�T˘�A��
������n��YXU��P��j���OgS�T��V�e�).Ђ�-uc&*�EW'\�y\-%r�S+_r�r���W��[�ŏY�G1�F�;L��t']npDZ�x��[�F�Ǌ���-���D�� �h|�iݧD¬���&���m:�!��iQ�ϸd�j��e֍���D�%��=�v�+��ҦFܰO)�մ����⺴�U�n�Q<�kƫ$�[�Ȓ�����os�ͅ��t�	�G�(���\�s����k`mb8Kɦ��m��땘���t�hոumk���k�3�J�$�m�N�n�|�h��Nm��НJfo}�q'��9�ְ)Ռd��	�i�ԯe")�!� ��͛9=�24�-��h�����g�����z�aB�N�,HI�r��z�����%̂��E�[	��Ž6�H�u��ng<�n�u֕�9�@x��ދ�J�'NL h�ٜ��U�B�'�K����*c���s+ndvTBJFJ�u#��s���2�����0؎N5;.ٌ���TUa���	P�dF��V�j/��d���k�(�����m��Ŝ�B2U{��Y=��\ߦ�>�B�6)��-�^mb[�� �OX[�� �T@�=��h�iL͋�wӝ�A>�۫�h��lN�fe�9��Z�e�x��Қ�B�)��D�ʔ^�Pe��#U&&�>׉O�C�Ct������m�E�= �r��	�՜�����-���Z���+�ߎ*��S[ƳfD���e=i8ܡ�v�>O��:o���MK&��̄E�\B�G+rݗ.�,],��˛��W-w�HWV3���5�����)�;�=Pͮ�5���-ݜ��M�@�cr���2��!��[B��du�'���
�O[}5>'C���ש�|H7�3ɶn9��kkn1�8�{��~�Q U�ǿo�������W���Ɍc۾��/n��7�v�)$T?�Q�D�@�&&E�,� D�	T�0�
e6"h���)4#5O��W�ʲ��{,@
]�CĆ�T�ffV��sk��<���;E�����ՕY2�7x:#��P�Y8�t��Eĵ-�W�	�	ւ9>�vu
�czf���qª��b-�.�c�ǹ��v��*k0ӣb��kK(�Z������/:΃�bD�����a�7�+&�����$oe
�&�Da��{(m��p�J�٨1մ�e��_Cj�R�Æ�cw_uv۝f5��qU��n;�`��o4��Ns�v�yl���>JV=7�JJ���ʪl�	�0���Xz"}:��\�ei?^�-'���ԳϸQ�J[�^ЈT��J��Ar��4v���l���� ���5���m���H�ɮ����R޺�kepL�]�aЖ^f�q*EENع��=���zl�ܝ���*��%���y�;܋,e�Q���ɠ������ٓC�d�f�'�iC�Y���9	���� 50Ӭ��d�����)��$����d��3k�)vM雝V�����.�,"����滠�-Ψ��6z��{ܞ���]0����:���n�𾛙V�x�Ӥ�h+�ր=�}�6>��r��a9(uGA�;(a\pRj������XlB�"0JH�m��m���#b4B�(�l��!
!J��Q�щ�0���m�Q��rB#A���U$?�􉸄hJl8J"��*�R���F��?S`8�mlSڰh�AMPS�&�LlK��y��~>���������:����U��T]�P4ղ�Xv�N��@��>?��������?���
��au��)�A�n�d��45�c���i(<y�9���}>������?���3����$� }��բ�5���]��4fu��������!�{[n�4�Gs����vo-1MBm��!��=Y%��c�^� ���@�iJ/0�.���<ǐ�L��B�m�V�즍nե�#��5w{��M	�6ѭ4�y�/E�:���:�Jt#��R����ZE�7�i*��1њ�U����������IV�y�4|� <��ձ�cn�ۻA��~^���6���8�.������M�^^E:�q�.��ݻ��P�]v����y�y۝�d�g]�<��'Z7;G6�:	֘������Z=Ovo[�w�q�3�1�F��ƍuF�\Mz��d��gI��t�y̺�=N��%���v�����Ty��z<#��������{��]M#C�0��;Wn��T(����I��xO���|ڻE�cSU��`��4�ǥ�<�bϑA2�����iם�m���`M���y园Օ��n�[�RNg���_�iK��S���� p�.T�i�Ԩ$�QBB� >�}�B
����� �h���H���׫����&�c�|o��2�Gf-�l���֎�3� ".`	���z�vA~�9�`Q4M�aJ����ߙ�Rm`�u���wwW��f�O	�
ͧ^�6��f�|Ǹ��ޙ�w�?�ǣ�v͊�{rԓ���|w'X��4�&��5��[���','z�j�Tq`��Y}�m�jH;w>ͦ�e^4̆����.�|D���;��)u.d��nv%��o=^�y��Օ^�5��Za�]�kۓ�=��"%f�G�b��O����&�Ӆ��Tڷ����Q��ޭ��7;Ո��3�l���S�2y�޽k���?�a��x �<����;(U
��jb��[��tzh�O[N��:4�-�����m�r��߄���
��	k�*��uv)v�{�[�L�}S��$X�tV���x�����ᥚ=��1Q\�n��5�f_e+V�&m�e����l��L�Aׅ}PI����=����:'�.�zS��U�s0VNe�ޗu�]r�M�P�{�i{5��T�VMu&
y����Աv���>�xhx�P,�w������51g������j^3����`y�*��ޮ�/>�j����4������׺g�]U�rK�#��.J���9�)u-���T9 �9�`�p���/:/�,d?��.}��zh(�������,��ߩ���s}��إ`��'(K�=�������㞼�u�`�q���OiѾ�m�4�0�",c*�b�룚$=A�ٗ�e^=��xU����OR��܁>��Z�#�!�l�8��_p�=�4
M�.�k�ö�`\52����7��g�.ٚ}�^�z��$��ޫ��i�s��zrt��y�b��t���n��M���,�~��r�ȱݻy�2n������=ׄ��샛}7ƪl�a�������K���Kކ��zn��r���X޳�-{��k=�h�;7��Y�[�Zl�0b�Oze�����ac({^�-bjx��Ԝ8w {u�����$�s�<��Vf�q�������g����O|�w����a����̙(R.�w]����n�/Gv'���2���.`�o^��/+׻��k#�eP�y�;�8~��˔�4dO�TY��5������*���R�y����M�����]�Hr�o%���YH�=]7u����0+u�V�yǍӔ%���z�'�e�`��{L/�=Y'{�C������n�s]2����'/_�6��u����ߧ7ݙF������J��{zR[�wz��u�pб.㇯d�C��v���#�#���?�]�H�%{�>��[+sك��t�+}���B?vԝ�賭LRe	�>D}�&z�$�{�U����=��{*�
r������3%K���;�w�,�f��$��]O|8ʱ\����w��%50�	S:���}��k\�wY�P~��XVT�t�OMW����2o{}Q����w�7!��{��ZZ;��/��G2�8�N�Ҹ�_>���h�����z��GC�e�I7跻�r��6�(V��T���.op����u7�Zo��=�pb7� :�zu�W]�2��!��� ��d#�H�y��+�NK�(W��=^l2��ktbܶF�n�Fc��7�s�ķ��<ǭ��_��3$z�&����R������A����Q�'����׷ݼ>򙈠�?t�E�pXolֆ���$���92r���.�p4sx��öX�Q=|j3dk���t��'ol�Lٷ�[��!��e�7tA��z��,Qʟc�ϵ���@�����}���Һ��{��W��Z-W����/X�宦��E�#oӡ�'�-O,)���;�d����z-���6��{.�+��ջ�E���������R6z�߹��m��}㞑��_�V��7E���e}�%u��'A���of�A��M�N��L�zI�#:�V��}�d-m%��ўf��t�Y�[h���j�������RU=�^C�5TUyf��ׂ_{����5^�U�.����n��v�]s���g��&U�e�at�����q�^�8mי����s\�X�fn����h�^�Տ]`x$<6��up�{��EgB�W2d��#(�e��0Z��f�З������n��8�}�/)�lV�R�84���t��n����x:'}Y)�	�k�&c��u��$H��H��5.������LkY'��N��0!�02�>l-�@zZ�٧�ʿ��������r#=�BHN��Y�N��z������J?�2'�rB�ײ5��/]mX��O�W���i���n���������K��o5����{)�V\^�t�C&�A��ݧ�[6��Ԫ�mIk��Gy��|.Y���yދ�J����=v���ռ
=r�7�Vf�SA8b �� ��|U��z�ۏ}g6�f��ɉ�%懪���>8x��]�Yko9�q��t��Y���ࠠ3�ܖ)�9J�<R$ּg�;����T����Od��_�ųT�X�<q��gf�������U�enUw�o�ny���'~�~<N(ʹ��O�7��)n�)z�x����ƭ此Ϟ�����N�����j&�2��ufO
��z�d�c��k$�A��8S�L^����<!��̧�t1��}�sT�@��	Vi�6�S����q��Ea��]|I.��A˶OZ�뫕d׏�����8dv]8�1<�Ӻ�#[ָ�:�lꎥh�Х���O�H����g����{�Z��n	�T�s�9�z���U�>���,��A��g�t�w�:����cu\�^�D���$�����l �t{Eq��Y�a��q�7'l��N׾�y2�{M�%	=�4į�!��������:�=�I�6_C���2�q��Ɯ	������*��ϭ��|�̱�����j&{.E�=C|��OV76o���+�[�1��z|��N
^�`���Y��#�x��n�뽯-�6䃛s�z� t�}���8�L�_Z�N�w�u��Vҵ��ް�Q���Z��ҧ$�H��^̇h�Ȏ�k�1��ɪ�2�q�jr�v��~�HQx|�^�f�fu��z�ϼ�O��f�c��{��X�u��^�����{���܆��}]n����p^��J꟪_�� ��n�:�@����f\9�z��,�V���������D�H��%�7����2�vض=���!]�j��C$��յ�-?Kj�
9b��ukT� �E�+m5���ⴧE��m�=��^�_Zo�$�$�Aɳ�v]��ԩ�c|�f4ʩN��R�_i�5}���,�m���I�W���Sdpm�+=��`;T�l��t;�Eg{>�+�NtR����Ϲb5�i��Yd���5v���;�J�h*Wr���#���=��B���#�V6ֽY���#2x���f���v�'^���N�x�r`�u�^�-��b�� ��P�V(�{�~�ԍ�=�^S��䞯v%&��E�?z��~�̫�8�u�d^S3�A���+�n�a;#_���{�T�y����&��z�Ю���:=�W-f[v�p����X��=��^�%����=��3�Gi����D��_|�m�]�ݪ����Uj��>oV���w��V)�y���<ǅ
�n�IP[�_�%�,ƶ{l. ����z�����ogϑ�኷�9��ñm��;C\3��;ךEƎ��*L=��#ޜ�ɝ�ʓ�?���S�k�U����Q�Z�[W�NG����G���Y�+"�S*i�}gQ�8���)��;j52�]�59��ϡp�K�z�5˳�����B�e]gip��lYŜy���Uqg��P:�e@Er�ou����q��Y��Gq�:j���﫜�X����dܺ�.�T��EJ&�#�6��ˠ�g�Lpx9x����8+���3��h�a�<�|�I��������0����{/��ԣJ��
�[�?|=��)��X:��p�~ﺙ��W8c��ۉ�93/<�	t���
��^��Ǧ�W�X�  '��Ş���ݒ���V�Z�� ^t+�����u3�n���\����`���9�����oo�{�kI����ϕ]�4'0ٺ�'.NP��{N?�NK<l��x��yg��.8�K~#����ޗYL'�r{�Ӑs@����1��T���{��.���De�j�$����(ߔA���k�?yo
�y~K#��}��܎rZ��9���ʮ�vQ��YH��}���buޝ�:E瓓m=v�U�}p��3))���+d�1y�=�q�۶H=XY³;dڏh��mȥ�.�A���V�Uz\r���L��`�F��u��%{O�juw�zʡ��ݙ eb��)�H�ePH�Y�ٗ�w`l7:�jHa*C7Z�U.��:[pd��Aq���piaLY��wC���2�o(a��.�
��K�b�9u`�
��Pef}��Lt��`}����yO����?��E�ρS*���휎Z7M�=���s"�{}W�z�s�M��`P�p�� P��t���r[r���᧼�6T7��R�����{=�����!�|�O�����a�}�#���Q�S��2]S�~tTԧ��o��1U�1{�ܷ��뙞��c}�D_@q�Ĵy��q���ް�9�s�ޤ���!ou+ۥ����k>3~t��G�굳*��ή�Ⱥ�u�6EC��w��ƚ�롽c�\
��UX^�(����2��,�Z����ǧ��|Avqם�x^o
M���x]9[w���斦��=[U�Ti�/�t.�7l	��	xGO��L�;^;�I���d�xܨ���z�	}��A��6��*DU��c���쬰��s�����v1*�;NRfEZO)������ܼ��W�{�%���S�f�2bDY��Z.��/^Yqf)���NG}x�n$�[��޲wv�jA�Z�Pc��޽:8Ě��δe��ڔv>���I���y>/;�����N}ʞ�&���ǲ�Ws����5A��-����W=d�:��I�Ŷ�d�T��\�� U��wkLһw}rpMh������:�}�.��u;o+�9s�fV�&��ٸ��3N��Ԇ���ݔ	�G��^��%��1&����u ����;�9�Ʋ|o���I��50��:�8F���;X��a��"�%���l��t�� Tr��9Uy{�ߥ���eN��,r�M6�˷:���9�/շ�y�������rx�T����i�r�3��e��B�
ρ�ৈzLN���L��r!�^�]��#�~�������Ĵ���m�2���C8��]�g���뿕:��~�r�"#~��I�U�ph��)5�j�O|pK�t�gݞX�i���Ǚ>��w9~!�n�{\UL��\����+�~�yWG���}����yü}���՗P�2�j���Cq��_c1��u�a`x�^��yOij� /(Jr��B��X�e�Z0�͙��ܲ�K��NF����g�Q]�����崡锤}�Dާ�V޺��:3���wЊU����V�7�[Zw��8�݉�7B�Ä����u6#�,�]����nH��9(����ޝ�Un(˗A_i��%�!��g�h�v?s��,�ÞH�ӯ^�,R���nR�,���rѪ��NE\ɪ�6��m��if�����MH)�7�>UY��-+[��%��M��U�br�N�/8F�o*n���A��1�Ŵ�Va�쬷p�B�摒�9�K7m<��P\�ӭ'}J`!Z��mbQ�{i�K�A,�I!�;���7@�P��]ޥ��-���aŁ+	:^�a�5��q��!�Hc�M�Mb7��Tr�-#NI^�r��2��"�V���9/k$�9fC����d��B��Ƶ��b�> �������h�$���5����i´��ur�fT'>pٕ�$�Qh��M�4Z-���FXP:vS��NƧR����4�G��-}�4��N�̶.����ދ�X��SԄga6�!��΄���Q9�m=B�����pSMn�����].8���rD���,$�WC�WӁ�][�n^�0G�.*_/����'4~!*���טwш;�2ì1դH-��#��'D�!zҾ��.R���^��PШ��5�9HU�ɠX
JÛmT3�<Xl�oɺ��C��E���F@��}3z7Չ��7sn��;�L��J�X�>�}�"w��`;�Z����]V���#�/�g`8��+d�gON��Su��[�lo�V�&<���|��������u�2!W�H��6��}�O*���Ϡ&.WNT�޾Y�Ě�j[wIv��[���9��j���fp4�u��r�Mt��!r��t�s�й˝G���u3,���wXFe�ź�p;���ɺ\�Y�ˎ���>��Q�,;�M�2ݶ�=����$z�:U��_R���j�뺢^o���<�L���}��W]���h�[��&�9VyQ�����̋k8�k����z�3&ͽhu)�8.�y���O�	g_9l�B�-��N��4�J�6��K2�x�x�)]�ܦ+��MJ�3'r������ͬ�&�|c��������7�Ҿ��Q��)c��X��X�9��9-v��)�ȋN��U�2�yq�v��"v�k k�V�ssX��p�H5y��Y�#x%̻EM�qbC���z-\q�L�C!�Yc�P�˘'Dvx�[�ד��N�-w<ʒGM�֋P�����I�*��+��ѵlG�5�m��gV�kU�l�kF$�AAwU��vl�\�s��?O������?���3��~�{/S�wv��b*Ӫ;���U���/��t��EjM�w`��1����~��O�����_�י���پ�uIݓ���E8�:Ӣ�T�:+]��Qb;�U�Z
KXO�>9��~��O�������\�ןߔ��fJ(45m�&�1i�PU�.K��ъ'TPU�l���.�q~1�v΃F%�kN���o$��lh���6�P���H^�F�"�~�::R󸠵�֨
(b��lݨ
��zlb��v�M:4Z���m����Ӌ�v�������QE����@t�:������(�ζ��bx�Ί�U&�m�N����t:+T�ւ���4�PPkN���(;��G�y&�kU�ش�lm�5)���DII��v�M,C�thzqƈ�&���nW�f����9�4{�k8L�ͥI���Ɯ�K�fs�.̰��o��R������3n?�����0<+s��� z��]s�~�3�9�F6��� ��OH�b��ރC	�g@!���d�c���ߛEk3}|w����,2mN5K�o����lo�(;t��7@-��D���=A�t��St!��y8`�/�o^l����	{���X�xj�5���L�Ž�������;F��)A��f��)���������K,/��}���_S_	���h��ߓ����G{��� >O\�
嘎��ޮ���`��������,N����" ��i�?*J�*�f<�ʑmꌊau08�.�t��$G	���#���]��\X����������:i�v���U��lcy��٘~�L X�b�6g��Y�֗\�Z�β쇇�nKtW��9�m��S��ּ��0%��eV���)�}`��ۨ8��^�[ ��8�;�to;d��w-��,�nonk;4�4���t�qq����)�>�]^�&�kh&�%�8�1�z���D���m���{���!킕��ob�O��/��mĦy�.�sJ�Ϧ��mۛ��r�Utr!Π=4fG/*��#>�1w��??B�˄_�ā�Zl�}]����&<�\e7�%�X�gB��ж����״NĳF#�B䤆��vw*��?/S�T��tdK�@�5��mD�:�4��}��=6�Aߏ��	 ��o�->>�{V���O���M糥�n��ՐM��I>��.�����xŞU����bj�53�gH��mF�(y����`����]�}�;?�v���~������z��iO��)�ܺ^[ɸ�"y�=y���x;��� �X���^����{b5�:y��ǀpm��`1�/�"��*�E��e4��S�.E��5ӒKE�^�s�!���-�����oU��`��gz}r����v {o8����?LO����{�br��k���f�nE��?<1��M��zo&Dv��d���="��Ǆ�Y{=iV��@	�3���`���3]yѕ���� 5��!�]�>t�<�ո��}�5�>����޽�9�2�͗���\�M�'w��z|G��B {r���i�Ͼ,���Z��ޯ�Bp��fH�a�l�x���9���$Ms��ڣ�: h����XW*�[�	�~�>?@��� q����h�D��xϊtd.h̽�	��pw!�]��/�k;�S�gg�L�y�W�<ڡ����d]	�)�UC������S����\�é� 9�4�0Vd�c/a:�l�2%�����.o�V��薮?.������B`�0�,�y�Y.A��ǪFK�;y��l*�8l7��?c�}>d�mx>�������Ĕ��Ԑ�t�$~�A�	m˴d.$�cf��Ss9.���n(D!��}bbXY=8p�����X�!�E�D�Յ�3@T?DK��?S��eV���i��8;^s�^(%��d=�E^]-���f`�ⱄ5� ���Q;l�zd�Qb��В��BL"r�$����D���`y����	f�"��f�ӣ�����!�\K!g��lqyɍ`:�"KkX�L���Ȥ��$S{4%;�-Ofh�it���_�d�T\Cx/.�Mz]v�a���lj�:O�"ܳ)�`}z���ɟss3�O���ȮZ�c@�f�s�<ˋ�H�W���p}{w������ * �v!�^�	��`3G���P,Ϛ�\�a�.`ڕ�y������x�M�`:{���w{�!�k��T��Q~`2ރ�4�e�K���X��L{6_ ��U۪�i  <:��d���5%���L�9�k�Ob�X~|Y�=�g�P8W��M�转-���XoOi���v�}�p$�{�*�8��S�FK �9oN{�jv��������h��2��]
�wu�/ C�{�!�~U��4ػ�5�ǆ朧OK#���,%�̵�=�n��;*轝��[F���
����<(<M	c�i������T�������T2���c�g�^�,��ف��-%J�ow>��"���ƃ�Y��<+>��@ �9�	#���/����� ��R�ZC�pbz6ܯZuڧG6x� & �ű���H�-NlK�\3i}�f��##cǼ�)�?0�3c%+����#~G��9��������V�����坻��4!'oF��j$%ٳ�������9��+�Y.�y[J&�>���i��GR~���=��5�Xik�z�˼N���b��n�M{���w
x���[%=V�c-�}�{�Z������l��O�y�����e���Qb�\@�p2�ڤjr��T�f�o;o��gק_�{i�%N��MJSh�[h�Ҏ�!׼�a��IٽL2�چ�&�mk�Cm"|,O�Sl|L�L���:{�8��:��N�3�;�z�[% �-��l���1錌��Ee{}I�4��``:�O���ڜM��=r����DNGvL,{�!�
�v �%�70�{�OB_Ú�����m0�-��顼K�ě�6�3��3�'��i����x�| �e�~�ڀj��	Y���|��^���p��Q>a�z�b2��v��]t�sc?6�물S�%���η�x��UyfS��(c��	���T��|���~�U��"Y�a��K�/7�T$����@����<d� w�\�1E������OW�^C�����]��|� [2�;�g��̵<��k��O�'�~�CħL,�M݉U�Ќ[����C�W��[Kz_���*������KƝOe���� \÷��Xи�-}�p&��o7{�qz1�XG4m�k�~�;�s���3ڲ5��+��q�����\�]���xdޑJ9@fh�a�^\U��9�[`��n?�����v��3�m���&��v�V]aYze�Fg%:����Z/<R�S�N�k��m��\�P;{b���+q�Voe!@`��܉�x6�6�J�5o�ҽ<�3'q�q�W�/oo��'���rE�6
���:�����η��������>?  $���1��������/�����u�z^9�>j��&�b�XO��
i�����:��&�M�;����������`xz0��(k��>Lh$�
��n/R�Κ�p9�F��[6U��#�
����c�;�iX�y���?��<L�M�q>�wj�6�LG��y�=�#����>�wk�9��ɲ��ݚlX[�����:��j8��CwVH���7,�X�ٙ�����yBa$���Z�7�/I`�a�={*1�X`>wO|0h��������_���t�6:&�Y\�Y5�}p�0�9���v{�,�� c3d�̿@�sᣜ���o4�6\[�3S��.��t���t<��i�&r|U�2� ?o�3������9r=�hj<e�|���b���DF�к{�7އE�"{�L�Kf�o�T�%z�R*ȳ_;}�]\\����}Ù=���r޵L��ɪ�ٹO	)�mz�Jj<�~�L'�şD�������*ET���u0� ��M�L�L)�A�b�Ã�zV>k�ŊȖ��	mSm���R��xi΀��"���'���n�~��?�K�N5�x4��:�<�
Sr��\��l����m�K��>���I[i)�(���̌;�.��;k�~�_������a�ʄ�H��w��jͣ<��%a������7{���+��̪st���f�7zy#o��o��|ua�p쬐��=����~�)�O8M�i���f�7��#Ep}�R)���ǻ�S��x﮳MCȌ��F��%�׳_�ˣ�AR�6��]�}� �q]�k犄��8��mnU�֍H�_��G������g2'��z�7�n1e9���x�Y�c|@�O�ᑾ.�NL�h�~�ֱ1���)�
k��+���cw����☜�������~�i�]s��!��[�&��v�Pv�S҉*��Z�[������?�dP�l�VX�!���k�>^�:�A��_~��W+��o8#�۱��<����X�v��K�0K��;,�m�#:�1�jƊl�ю�;@w�̟T(�}�Ǉ���,:"�\.�cO|�ŕ�"�i�a�Ѭ��9ͯ]�����gO��Y(�6?d�_oOJ����u���}e.1C��i�#v
{�a3"����&�ZA1l��+XD�Һ��0�1f`�3�;�-�{,<и�3����Y���_	��2���@���o�Q��?<����B�/�>��O~�0i?�0��|���-�g��O�z���5���~�Z�A5�]�#��s�\���������d�$af��V��Lqc�%�=���ƍ�D�T]�2�f���A1�ߊ�А����WF���&�]�N�)=��`�-�;�Tñ�x�7�$�p3v���:scm�ٙ�F�MΥ�EIq]�����V��z��v-k��W�^O��0a�@��#�|	�|	��&e���^�皩�����@��Q;�R��^���0G߃�d�g͆l��ܟO�I�*e���h1�|3}���>^���w���⮃�9���D�μ��v�a9{ ��ygïwz��,Ҧ\s%p+����t]���"Z�T���!�q��r#�5X�M14�X �e��ޙ��5תּm(;��E�L�cW��[�Z�P��j�^qm~��x|��8fy���{KoC��\C�͒>s���9O�0;Y�Sn�m����q6��j�q ��q7W"+Q3��$�)���kC	��{��??����y	���'��W1��<����yC�M{�M/Wb�^={��nr�F��0���1�1��4Y�<�.ý�~s�?uŭ����>7x]QL��S�Vj�ͻ�s�\�N�m@mBe�r�2.�if��A��=�������k���!�gu��)��y�������gz�P��s�;;��4��;s�wRֈ<��8��c�z�]#`��sj��J2Ys>�@Z��/F����֊ͯ�i���M\�kW��,�N�����a��0�	�K9�azk�H�e�F�s3匬#!�~Z�uA���a�3;��w�OT��x�)��4��M۟ @l\4Y���	v>f��g�C�TY� �32��7yr�&9W�F��m�C����x|@���D�a�,�Ry�����;��ῇ���#X�bך!��mG�Z6�~S����K��b��,� ��LeV�!�6*�zχ�=�}�ύ%���_�u1���^Yw����x�Z8ξF��ֶ�ў�j�Y��r)���x����C<�+��O~AC����}���m�5D�4�݄�J��S��c.|� !��g����R��VG>T��ȍ(�"Dlaz�X�!A��i;&�*�-��AKI�z [ey���l����9�!m&�tnS;�dKD:���pA�<�P�]=�kA����7SC�c�ʱA��"CNLj}k~�Im�"F	[7�p�	�gNaߞ������읊u����C��b5��L��Q�:��eg����J��> .i�p�����<lEdc�_��#���ݯ��Eυ����>�Ȇ5ME7H*e��p��@�	�S�̩xb��k�J;x�����/���"p��?4��3SQ=�E�����q~{�%Oh�j���{6
��޽���/jh��kXw��̡Z3v�VI�Ʈ��S&�+��`L)/ͪ�SUn��CF��|��x��F�Zؗ�r� ~��3+����_��!��p���ܙϫ5�hj��Q�5���b���k�͉���J�L��WG1�ƙ���t����}j���v���a̚��˶o��b��#������ǐ&T�"P�z��Or�QHe���{zd�ҦYk��6vǲY�y�6+�ƽn�!�7��Sti<�N�vM5��ke��v�r�5n@[й����S�N��Z�E5z�f�&�x��}�2u����xB�k�vЄ&���p��܀l=��Qq@��/ze�6�[<��e)8��I��ů2����|=�U�/�8ޭ/���>���0��`4���g��Uۧ}k:6�b�2^��/ə���{G�a�f�.������qkX>�^Y\ ��_���7>��
�j���qNkl�k*Y����s���>?������5O� f�0��o�z�i�[z,9��,<�c����D�)eiIm�����9^v�c[8��P�<��BꋙG(z�x��t��+K�ۋ4�oj[e�It!@��#��oH���_@���\o�8~L4N~�{��M�(}�w7��떰P�c�#E/�l��-�1���4��2�J�V'N�-J� �9��S����mC��l�B�-@K�TW��f�5���~�������ݷ�6�ݡb�X�!�Z���awT	z&���,���Z����_A;e
=���o.]�&c�|�u�
[h�LͦM��|��~�sz�0�RRbAlQ�=�_j�$�Ԙ5h'K�7L����zw�S���ʟnk]�������W�������da���d�
���_ϝ���?�����_����>^��iii��9�e�K�+�;����)�����^Hz��G՚�,ua�3du���M��X�f�!�:����c��騿oM^l⌾�🰜
-����?�����Q+��y{#k���͏�ᨍYN����s�3ǪZ��VԺb`��κ�I�ONA��AT�❷�A�p7ɕ�������[8����ć|�]��W��:�a���vl`� ���P�-7;���<��hLZ=8���o4���7�n��;L-2�@��$��m����-l(��ʍ�z#-p,J�0�]�r~�����~yg3ڦ��܆���dN�_f���I\�{�=O��"��>���h�^�f��	W5���dkȄ2�A۹����c���~��W�Z�Ô0�]mހ�d/���T@~���>3���o���L�����Pv����x��g��z��ߐ�b�CRmQO��e{�u0��%��'<�v��h<��ZC����3�&��~��:�= -h�(�w�{x���߱+��D�y�?/�w��D=P߳����+�bc �����)ї>]�-�F�nըd��c�"Mk���jR�5R�.�Y��@Q��5���rgtgz��-�J'j��Ѩ��<�CA�\s��r��w��h.�\��w9`��5�lQ骷���W+���'����w𓺹D�^�ݍ����Ѣ���m�t5G�tԷy�D�zG�G	q�>wFN��ns'�ڶo^���f*,�9� Q���v����rc�Mgi�y�/g|3Gu�愇R�Qh��*����:�N�������PCB��5s��P��0�� `�2��̛w�-�]\Ǜ���|���f�S��ٽ�E㹲�w�-`lA�fK:O(�F�7����=���&4*�i��ᔦ�v�'j:BU�sw��t7��|ய��k��0�����!V;�xvI����Jݗ����`o�+�g�{j�f�t��ȞVD�sTY�X�{����%��̦Ιd:�f�_x�Ri�.m`}��T7�s���L��7��������m��j��x�<��>��D:�cV�	V�Mжʳ��8��$zPu��9E3oq��l��̫0���9�%n��;��倳�	��5a�-�ֽ�2��ux���n�ܾPVr²p��%l�q�j�`��H�a����Z�^�Wm�l���[/'Y�ѳG�w��mw�5�H��m)�k�^\����N���
�_]1E����ϫ�*��ܮĒ���򜾩#�V����g;*�������B�9�	�f�%�̿m��7H�{��$��H7,�5x���SR���ϗ)/n�?��d`c%��K�5���Y��������{��U��e��6�۵ujM(���VP�g(�0I9��i]�VZ��Xou8g�R�����{�j���sF*<\	Q·+ �:���Ui#�n�s�D��ž�@�:�w�NW�kof��Ov��%�ê��9��x\���r�ԣ�mC��Tܻ�zQ��'���ԛ���m֪�*���{:�)X��X:��'��u�*[���eZ۱�Y���qQ�<�
"�s�{��0K�D@�;߭�ET��! �����P����-p��d��?4J�ᩍ ����)f>�vY��Ȓ�q���-�z����`�ͼі�`�� �)��/Ah^[[�Q�/n�]d�v�٬n�ѮN]s�����"qmn�]r�쌮8�M�OY9`��]K~L�ʾL<ZO!��Q��Ǽs'-�w̵4.��|7�͸�oE��ռ��t�;�zD��v�ĥ{N!�c��BAW9�0�{M�+��V������0��V���:4f�	��I)A�_	;+\���[Dpr�v�w߱��^Gu�e!�[���MB��ݽ��F�b�N�pL��L>����I5���MYը�k�����3���0��KnnP�A��䵚3��T���ޜ���<�N'��o�U!��|u<ۏ*P1Y[�&Լ�T&�0��;h�DQ	�����%$�&80�)	���jP��i�2#!Hщ�l�$"u%S�,S�T+/�Fm�����$n�J�ґ0Am��D/�ӯ}x@�I #�[N�4Q�Z}A�N��?/˼�Q��t��+��?	=uX���g<��y��}>�O�����~����ʝ���|����ODQ��Hv2h�Ѧ�4�z��;t��������O������}������s9�O�E$ӧ@|��]�QT6��t��m)��Gh�J}}><��y��o����������>�*4:vɭ�$�=[t�����J�͚��i%���-������xG�M�T[��OE[Yz5�=<Wd-�q�m��-��В�:GKA�t[b��pb�k�`�u��vtww=/N;�38�N�g��a)��ɧZu�����f�v�R{�t���F���v�]e�b�1�53ZJ11�γ^�����4bZJhh&�^[��D_�wl��wi*��F�:���:4tuC�EZ+�(�<��iǗs���1:���[F�&�h.��V՝PUV#TkT�k�1����F5���9��IJB���HP˱W��kUī��M��<�:����i����[�Y2��sg(�Ʈ�1�S��OL'��(FI$(T�Y�9F�;�v/<ݽn��z�;���#���C � �}����_���ޙ�0f�"����~����[��}��Z��7˦0���*1���x�?GDO���+���I�3�Vo
�%�5�hg��K��1�>F��4�v
�I���:Df�U�[2�.�WXN����v�f]K=�	�6���;�v-�f�\d:���8�kc����6�����3�
"j��4Ȱ��B���X���'�SS�z}2d��~��Sp�m֣ذڊ\�٦ 3V�;���O����L"�]��04�rZ���\�[��o���X��'�HX��w�����'WV��u��y��:�9��ͯ�=3bWA���;�6�v1�=�Bf����1��w-�B^��jp��v�Y	�=#҃u���U��"+��;��|r�뵌7R����Ⱦ��W�rEP���/�U�{a![�̂K�Δ�r�x5V0����iJ�݂�e������wBR�ɯSG�Vn~��Q-I�w>op�<&��wG;sߎ�'�,�����<F(�m�k�Mo(9�!�3-
�S�AA�֠#���W��x��<�k�^�Iq�w�<ޡ���W��J_k�,�Џ6m���OFW&u�ll����;:��p�/��S���{7����6�f�S�t��0e��;-�z�Y���ӹ>���c⤧u|˶����q�T�-���7a�8�ͻކ�M��&b���}�}����UB��a�~B�!L�)@���aD���ն��S�����Ae�j.>��
3�n|s���׼�c�okLv=��C�V��E�h3%�T=F���ǫ�f�s�Q��f�m�SyC�]TT=�ɖE��a��uY�}�>�����q���a0���7�)��*-֡c�ꗎhi�\�[���j��;�D�&�J��m�0�1�<b�3#���}��x`Vd�/���1E��p�o%"r3���7���Y�wBK46Ae���:Su��lF�V���}����E�������Fw_8��:�%���4��`�B<=�SƵ�����^{�P��E�y=�P��3�N'�JK�n�p�,�2�<�z�����r�c�ᷙƵ�!�	�����>tڋ��w������������r�hǠj�H&ĻuO0����7<�R&ivr���L��èS�izk�$1�����a�c X�*�Y0w��_������/d��g���xy=*6�i�܄!97��#���lq6�љ�Y����$X�$�X��zJm��}�RNN+S�W�r��5�\U��E=���B���zJ3���}�p+j�V�=��J��gT�(pf���ǭ���Ao!� �p���FM8�Ꝿmڱ�s6�q��1Ԋ%ڴ��'�\+������˵/ge��;y�Ds,�L�P�s����B�����׻�{��m�O�+�WAJ�� ����~�?�������?6�0�����q [��\
h}́E�>L!5�HLܭ,����U���ߤ,�?�FE{��do�WT6��b�Qz��*��ڈa���� ���.K]Yٙ�k��a
�={'���0G��/���I�,�07��Xw�\��?n��/���Ku�8��ϻ�״����g�Y_�=�i��]��Yݗ��vd^|�v��A>G4X;����_RPQ�o�x�t�G�3�1:2��<�: �Ħ[��4��0�ﲰ��t��X���W��6F����8���X��E��"t��nx.�0�t�Vڲ1�I�n�i86���U���FS>4	=.�D�76կHf�}�|�@r���8�I�۸*)�l���{����M�;b���@O�Gw��E}>Xtr:~N�?�Ϗ�z�⧓��\��Qא9�d��'CJ��AD��A�����,�\�&!?C
�46�KM��eݜ��C=\��՝����1IG[�yL炘���	�И�X�;����r���Y��T��=��]��4S��V0�iS�e�&��i���-gT-+V�`��D��=���k����˯x��k��端�����΀��h�kq*I��ԜOt<wB{U�sz���HQv���}�M.uJ������~? CQ�
�R�JC0/xW'�	�g��}f��##({��/?c�����Q7�J��Fv��˱�l��vp��u/�S�="Y�3���p��L϶��}pu_�W34�Ĝg�u����i��g��9����hb�xl�}�'矖>�������d��t>3E��x����Q�g�o����m���]Q�����w2��7L��n�[Wf�>{F�Q�p��  �޸m��A���v��P�������������DC����1M��36���.�_�b�2�-�Y�O~�^U�"w�į��lQ�;}�Bj=Y�6#X��	Eۧ���1[^�zs�����^��k���nW��x��1� �a��FEґX��n�	r����c�rԽ04���ܦڅ� Ũ�K&�Eu�s��>Y6�:�DOir�$����na����-��K�k���9�Z�\��oBe�alR}��E6P*s��&z�NJuqYfq�d�+gdC�� ���tl���5X�>���˵O�ؼ��d�e�Pi�������*��e\eLNGVė�Wg[v�Ӧ�{Ϳ ���%ܫ�p�6eD��D�uy�yي�ү;3Y�/5p=Ge@�E�Ă�ҳ�*ʱ�#V���/�α[��^�M����3�R��}��������6�%s����EӥEV���Ꭽ.F��&�s=}7���&��Q!4�UT�[F��<���~TхԬd@; �� ����nCg���&r����%X�ԕ�c�FS�N0�$��}>^C�{��)� 
�{�@S��m+��P���÷ҝ���<���1��t�m1P%�����DL"��K_��>�ώ�ڃ�I]�\T�5֌��HJ�3�DȐ3�{�%�zc[+���5���3?�H�g\�8'2���CMk�p�0ӦV�KH���˒Ɋ0Y�o4 ���9��٘��AJ:�;1�_�Լ�I�����H��<�j�y�잁�g�<\O6�fka���sH8;U� yz�R�Zbʊ��4y�C(��q��gz-=GT���I����{ �;l.3Ւ���7$���X����õ��� +�K�ᕿ`��3��;O��I^�pu�U�[���	e��b�a�k�r�̕�|���^a�����Ax��5�(R��tSz�D��n���f��~b���mg�wCT� ����-�=s˾�x�6��2��aeǣ�G���2xG�Mx�󊚘f􌄜H=]���3����E;��v�y�W=;�!�$�~#�w��#���{����ı,p2b��^W6��޲�FD$�5	٭E:��f�5s��FF������ N/�[[��ķl���ꥧ�Q�k0v��(��ƅf�Bɲ���}�~8��=j���q��D��*�P>H��H���z�������o7���z�@ƿf@�P�b�(t]��"Z�T��3n⻳wE�=�вDg x�Eb>>���"+��:������7 �_�$��>��7�2����h%�+5��7&'�f\��'��Da��쉯�M�b�Jc�w�yjNSแӠ<&��t�]��A��f8v�(��]O�rO�RS���k�چ��|�m���l��&���	��؍S�m�]��nc$�{Kn��2�]S���yo-�x����
�r�Ķdd��id�s��x�h��y�we+n�5
�P��n�lL��^Yc�Q�5�*��׊.џ��x2;ƍ\�S3�h~`�.���xbۯc�����9M�>�7T�_<�R�lj�m��c����m��;؝	ּ�X���*\Am�ݯ"�Sȵ,$U��q��Y�Z���/�a�]���9�h��zR����C�f	��#\I��/�*=�hЪ�������Ɋ1	=�*���ާ�ȏ����<5�H�U���N��D��
C�%��{1��K�)����>�Uc�`Sv��T�-��+���!�y�r�m�gmW18(�/e�|��#3R�d��˺��43��t��r]Օ<�s�b�4)����%7�W�o����m��c��']��a��4k@����W�|�7������{�_��
���z��B�_~���;~�?�?��w���pm���&���b�˖`���5�]�~����� a�6��O�`�L�v���k%��(��Y��:{К�ư.ML�&Ļutm/>��>���xȽTD�zμ�@�NÔ��4�0B������\H���,��`[4�b�QkrY�F�3�i]
RjZk�bi��Fti�M�""���?%�x��jɵ]�L^�ˏ����BB��4�R�v!����F���G��=��&tZ�-���q_�y�sr�nAcAA�AY��^ ��ɽ��`�2{��i�Qbi?��@5ϊ�(xX^�%u�Ǿ�^�<w���8�$ �y��ֽf(RIAKA����(V+�i�=M�|�+0%f�w��ĵHP8�5���� 
��#`�1x�~�l���� �[a*���+2��-�(���o�d6KM��V���o��o>L�>MI@M�#������p��s߱E6W����J3b�<��.��m�T�wj�jP@#�Q7k�u��^��Ӫ=?D�L
�S���%X�^Y(;�?Խ����K����!YP��hձ���k,�}��<i2�R�*�k�Y|<�Y���.T�2�c��h.�Cݜ+9��#� ~>*�E��垍H��q�Js:�![��u��ԺN�J��*�9jݒ��6��QJ��Z�6�oE�j}u�ۑ^oW)͏��@ хJa�4�A�G,x{���a���Y�S��RЭ�\�������DD�'㸇�_0�s��w����b)>�mַQ0�[a:8d����D�jIOc�Zĝ�i3��=>2*!?4[��3��S��])tR�=lAg��T�Uo��r�^����x���u8�Ŷ�.�^���s�R�XH��ڦ!���V��q�gճ��8n�BY�2i`�)�#���Ƭ>z��������l/�۲��3��7
�z�YI��}��/�>X��g��U�^�q|�(��=��[�����&��I����بK���*�r��W����'���ڨ���>U�,�t�,��Ȕ�v'�h.��^ ��u��^�ؽ�Clcj}�/D�U�dvn=�a�;]F�U������of]���;`7^ =S�TW��6������b��k��c9����{�ڵ	$3|�b߮*O�Q�8g!Yə����%4'���? ��ܜ��N�y��?�Ve;gC�P�)��X���t� �:º$T=�-�?qfV�W�H�כ3F�H^m�Z��h��T���,��H�b���(t�VH�RSF�^�5U�l]��**�=�|(�I���C�6��F�c�G{�}���k��y�[���`J	w[�X���8u��hyN�3y��q��;�z�b��q���(�J>�eJT	� ]�ו����`S� a�S@R�J@���{޿|���u��;@��REO�_�#?��|���<#	�A1-t5e;	żD�zw���ӭ[nz����'�{٨j��Mt&s��J�y1j��$�tӞ��M�VХ�n�Ȧ��,�4¯�uk�*2�>A���ZrR�b �/����95���:e��b��J���gm�2�3y٪L���3%�0��,6˷��9E5�]1�p-��Ϟ��F�%��&��	�"
�L���\O,#�5��y���s>4�����?]*{�����\\�!�����tĺu�H�e+d)q;��Q�R�7��k@Tn�2�]i=�0���p��\��-gnN���#m�s�J��}ކ�vB�H�oT�:�^<�E���r���l8mxw���Y#�^Գr�.�WZ����x�P^������1H�}w��Qi��b�o��A�})��� c�z�9xߙ5�i_�z�y�=>�%�����" ��ʢ�_��R�{����
}J�����z�޹���k�X���O���Dc0NC9�� -b�rQC^��4Ȝ����`���	w!�*~Ǆ�����]�u���i6fK��J�
�QT,���@�ɚ�J�w���I�w�X��U��,�Y^֫�L��/�=2������}R�вۛ�է[�Vu(�+Y}|Z����֭{}�sn�%1��tw��WD�f>����W�ꯟ L2"CFJJ��)RbC+��#=F�X�����.���|��L�]�Cڑ"��A���dkM��:��3�M؉�37K��״��$m�R�/��\��;�|�:����;��G��fdN�Q]�O�"��k`�L�Ғ�A�47�����oeKW��)�=s˾�7��Ll�8�-��X޷]�z�y���x̣�m�$�������#�,̕Oy��;���j�Zc�vü�|�����Oy!Ӟ|�n)�=��e�*ే�#6�P!�T[���H��:�3�z9L¶�0@�=�TG�T��j�W���E=0��J��c9���&N�Վ�1
-��suU��{w�x���U�(�nD�M�f�+�/��P�����>0��,�z��<'�~sE�w���5ⶮu�t�s�ܑ�
�..�{m�V=����������b�Җ�����~}�$fZLY����Ju�*|��Z��YW#��z��F��[P|�T�\�U]�l�QZ0JL�]��2h�x����f+^�#���S-s�*}����&o&65,�	����{���oѼ7(4�#Re�n)�5 �L�n�[��/f6��K��郍$u̢��nйV0'AT��+]u݇*	z�1�;�ޗK:l�/�����O�j�1,���Q�׎����k�/^w40dy�n9����ٵ�\�6h��F�va&.J��Y���Ye�F��8�17B�۷g���]�;d��F:Ĺ�"f�m��.9n�������0��U�������2�f̃��[Ot�l�e�K��M2r�Lu�P��9Gw}��,N��X_aW��7�v�]�s2��S.Xb&�m�VLt��Ot��E:��x,������5�/:*��N�Ѩ���\r���l��'�r�WV".��l5��(��y'�R�ib-]���g^v��7}�lz�e�_�{�%��,!7|�k�7A�<�O.�:�ZR^��!P�`�"��/d��Y]�yq�f^�;��0���?�7`4Ix]]�D�f�Y��!�����1V����2�߹5�]�u��1�sCT����iL�8�#hb_,D�]��6����0�RZ�Yh@��d$uY�8��FZW���8K�lۣ�m7X��B����P9��w>嬆�����x�����u ��ԦЀ��b�vX�G�NG�Y�rPV��	��U�n��(-gD*�<�c��>��yۜUjZ�Йu��oZ	(a���p�"1e+��U)�G���?jק:�(Bۻz�5jߞW���;�i��L�v��z�<�ۦ+���f�RP�d��͌/i��e�QGr���4�hż�WuÈ�L�'�I��f<m#g3��i��,Qt�	X��L.����0�L�@�Ysz�U�^�l��N.v�pg<��2��uݏ���/�).���������e)6����N��c��:W���;0�=���K�jB#�[g:����Cy�(B9�P��PW���K�����u�lpdB��:��`,�:�X�.�H��WtwJ��6�ѝZ�Z�'����拒��6�����eq�9��3����՛��ikm���N��[��B��]H��>����r�ݼeҠ���j(��-]c��X�8��Z��Cե��i�+{�H��[����g��v��"��ةm�\%��Z�ek����C8]�lu ��y���~i�y��sI]g*y:�w���%�NV	Pc�}4;Ԗd����/]f�9G$��Ÿ,"���ې u��ek�2��`��]�A�2�C��VԨI-�Fml����gq��n��*b��;1�w9�1 �d��ݒ����!	H����w����̓M���z����2D�w�\̬�4g0v�~u{瞧�޽���֚���i��햝V;r������F t�O�<��y��?������G����9��!��Q�����u�%�H�4v��Oc[Q�C�@t�!KI�_ny���|~�������~�����s�>���j%�k[z눋|ƃ�""�ډ�F����Ӊ���'�������|_O����}?G����g��}&���tS%1��m�0�A���hi4����\R`>G>F������t�5��U�4����k1����6���Y������Tl��[`��l-{�qPDh��\I�-��ꚭ.ֈւv�i(h6˦'Z8���F�%m�ₗ���4j����cM[kG����%�(+Z-�`�)���"���@�m�&4>����x�d��y��>Wt�%;{L�#��۱m���*�	�ղ���c�xݶ�a
4A�6~Ic�� ��D��
��p��)hEF�������]�ϧ������[�^��G�n�(�rѝ�Ei�á�qr�	�3ͥB��W�F>NZ�����{�����:�REq�����S�a�*��peG0���Ǐ�m��|'�b����Rb��f���������N(�q=���"�s`����K��}.-%���S�5s�oHx a���]G'�3�R��6o �p����i���a�K�ok�ㆤZ�]O�q�pCs�@��r�n����C4{���4�[nl��l�CԵJ
i�L(c�|�N(oAk�3����$lK�P��]ٵա�m��G��i\�{@π��~���HS��}��`�Ő2��q�4�����4	Ϣ��������ƶ�ȥL�}�ǳ��R�����)������2>���-�D
��ݡ�]U������En��ƵD��n�X�9*ME��a�w>�7 ��"8P8�鮹��3,B��ˎ6�T���p�7�FEj$g�ح��� k?_���_�-�i���Y�����#��+&�-;Ɓ�Y�k&���[�Fw�r!�ĨEb9s�}�iB��{:}�Ю/vsx�u2�M�`
`~5��3[m*2��,�w��J�c��=�VW�z�MH��Ǽ���:�u�2��C�6
=5�<u�9����nw��x�Q08D:���*)@ ���߯ÿ�X���	���h&�p"��,34���u�񤙱�"��]�e̡������ޮ�����S��::i�v)d��94�R��?���V�/D�{���ή�����B�G�Of���xQ �_�jgi/K ��<���{�ES.{��Eec
	E�@l��7Sqq������9��X��&�h��B�ȟe��3+4�O/�U)�J�l޼�b�;�s��P�LS\����kƶZ�&v����M��#T�q�c��R��xM�;��w�um�*��9�Z������TB���eO�z�����9
�)O7�M�(�ڐ����ƭ#+)AwRO~Q�K��������F���\,��=gv�nE�x��ɱ8I)�]Қ��'P��u�* Bƙ[�6^�����q�>p
�+9 e����N_�E��Q��� �x��������߈������d7񢃱<W�8������A�|�d�r[<��ؗ�«ym}����YOz�����U���� ��(q�H�z/Ҹ�¼Hި%"��cf�q��[JM�_V{7��Z2��t�m�۴s�y`t�Z�Ʊ�µ@1�W�mO�*���y�tM�嫟>�*w>;�tYjތEc܂�k��ޙ�yd���i�ɿ՛���!�l;����@�-�7��"ޛ���ťҘ�߮�w���y����U�3�ZIp¢R�D}��}�T�������D����o����{� wf����|&HQ��⑳����z��q{��x���jYYcx��]�<�u�ꀢ/᭣��',�"� �y�\"�1ٰ�O�y��DLR�퇹�7u�f�1t�4�M�!7X�X�{��!K������ZbL�*�3��6w�3��>?������^���$F��A��3b
����t���f�/j8�7Խ���\�X��e��K�߼���`k׳�Nʽk�3k�F&޷�Yu��� H>�r��^����P��B6̪ǘ�,��z���陦B`�O�ŁT�c�:E��yd؎L��f�qaF=�iy4��ʍ�jT���Y��a��<�!�8�>���:ӑ=�V:})���qI�n�7]�� 3$o���k��1�wE�Ѭf�|����LA-p.y�g�r�_�ݐ��u�wew'�U��[�K�o4/.�q�����z�Ǩ5��*}!B����,@�ݓ������2�fI '���F,�R|��U�fef�n�S�`�>��4#8A��>;����o%}�t.��¥#S�9o����9oS8�b���%���.�1-�R�r�G�͊5�u�S ?e6�:�^�=Ӱ_wJ��i�5kr�R���m�4�1ZgYwK�v�<�[u��o�m��\a;� �T$W��Ȋ�@N���.���47�<2jއl�2'z����%�{9���	^Xv�p��D���;�+k.v�+Dw9�࿶+�,!1�$I�+	i�s�v�k]ķG���_kY�=Y�'F@|��r]��<��g,n/��	�	mk�Ej�az"��kB{;���AL��� �V�_��Ca��>�D#�,�o�C�`�^�G�R�c�qw_oQ���}ż��܄tr�uS�G^���'��|� �9�><#B�"��~��%�+i�3*w4�Gu6�X�4+5Iǰ_�d��.)�	:_����UʈhV#�z�t}��K��vu�p`�୲ݚ|_�l��m��.K�0k\���1l��s˾�x�aP��Fք��|!zrS	��M�\��Oώ���{�����,�>�jSt��Ļ�p���F����r���iO���`��C��6;�#����x�k��K]n�=�����&�R����qƀ�������RW��Ⱥ��D?���j��_�+Qo��Y[�y���o�iH��e!��E�;�%�\�W �����;�<�"�u�k*H9ڳ�}i��oI܈:�^1�Zm�ytM�G�Ӕ�d7��-d:��!U�$ƹH�a�-T�����c���K�uε��c:��[[��	�8"���P02�:V� ���w����篿���~g�V_�Y�����kb\���+���<t
� ���jV�i�D���V��_[��K��-��
��`b�dO�>��s��ݘ��f׳N�ð�v�ݩ+E��d�ߚ=������$锟m�h�i��UB�������B��@�p���E__,��Yk�P�nT�C�]^�4z��C��e�0�����.}��!Y�*���U�����D���z�?p}�i�z�>��$N�Ely�_Cz��ML��4�o	�Է�b�6��<۱W�1L���v�;�������!Phs?�j1㼨S�FE��^��㊭�mm�a՟zj-#�p�]�n�Ja�嵰���f�Q���#o��t��}H��g�7~�.o�����F���e8^G������!��*Kw��5�5�?9����4y�iz��jx���By��O^���k[")��<�i~ڎ[�*$CX��r�	����ў�8�v*u��no�OS�A�C >�4.i�L_K��~N7��`&�\ӏf�����Ļ*����W��箽9:��$�QC˗�ZæQ9f��v�?s�qVL|��Sx9�Ɣ��� )f-�;���i�*!�
�.p�#��;��u(���Nᛛ �kHuκ��ܫw��(�;����F�ju�[]�9+��S�����R
�FC!*a �@M")7�=�o���\�=Է�c#��%۟M�A< �ՙD��
85|"����+~J�,�b�C�d [D��aa50`�h���_�c���7�����_�W؎ �,b3ła���7r����G���ϕ-$� �><=�ޔ�Gʳ�&����>�?�y
���;������k���"�j�=��ޮ�!ι�D��Sn��#t�'z�M��Ͳ�S=���K�jLݙ���B�t�T�LzoDsBFBm^��ؽ{�֑��!����xi�=��"�m68�%r�QkO���z�8 �(R�����c���P�ͼ'���{k���kv�E�6���6kܰ�KU�tO.��C�{� �Z��1����3*���U/[�{y����YX�ã�e�`�c��sbS�oT:��ˡ��l@���[�1�4z�H�5A��]0��Sw7:9E��09Q4.+�wBv�mK�t�b��qm/��1�dx�Ȅ�~���}��J�n��"����9S�"�ֺI�q�`6���|_ ��0(��xn}j�mzgbCd�~uT��c��L:�����Oya�͍���nj�	ۈ�:�̈́L�&㌓�e�Q�g)�D�Vew�;ㆱ�ݮL}�=8��b�:S�|ĵV��熒�v�J᷎���*oog�q�b�j�Uh����ǡ��!�v��Z�6G��b�`������V���th�n<���ǟ�E� �2��P��zߗ��W%����B"�a˛߁j4 �<���9��R;�(����#`�\*]�|��x\��y�Ψ������3���1Bԉ8+��<�3�'QIAn;�7���FV�f͐�46��l
��M^O�|�(��z��顡��3����l��ޝgG'�Ӏ�����5���T�c/o4ˮ�hL��7;hA�qz�\r��� W�'�W��~0���.a�El���)D�f��3A����)q���&'ǟ��~c ��?*ń��Ghn�����Tt���3���9
~�^�z�o}��u��~t
#RG8�m���;:��h���c�ek��w�Վ�5v[wp���Gv���B�&�4$�W��~����K���U�L����t�'Z� �G:�ʆ�_p8�_����E����,XFm&������	�_X;��|n��݃v���tQ��++�)6�����
�Gxa��y8��B:������L��� 5YN�|�^��w�k��E�i�y����%ݩ�6�E�F��`�a���M%����~O�L��B[>�m4a�C�Rm`��W��t{��Z�[�q��ݥ|e��Ǚ�SC�hX�pbhU���`:�¥�J�*�wc�օf�ěo��.��t�r�W!���zc��S��l�h.e-�Z�T��:�dKL��SWW^息\QqF~�_��2����2�	�7��ox{��6	S��S0�}�S���9��J��낾�����,W��k7�2��m�����&s��d���0%��~L��@i��F`�`.^��C:6i�"ۃR��8�6/9ړ<�/����bv��lp���Z�mⶅ�x,�a�^�s�W���>5@�!*K`�����ϖ�!��O�h��S)6��Te�چ�k�� ]�>�Y��Y�`�{��3��y��4���ù������z_C&8��rۓJ��o�@�oT�����]�_�ݒ��C��s�D�?��Nm-���z26��K��Y"y� 1�B�9瞝����L��,�9�gh������~�]����ֿ*��HH �i�K��kA/<"?�yP�y{�I��7Τ��EG��WUߠ�~b�^����^�O���zq���/�B)m�N�v"!'-~��PǤ��x�i����m���.ط��.����:Y���L[9z�K�-�-�~N�F,���}��tL>l*��K�������D3>��.��.��*�`�|�<%˷�vK3��n���i��s�*�Gi��0R�v/�r���:ǝ����߶�r�K�l�Z^wC�mno��8�+��[E��P��sN��3� ���Z�oeK,CX�܎�[���`6G"�e��*x��nR�
���G�q����_}ҏ�`a�He�%(�*�R�P�������������(U�D9}>����xＫ'���E����Bz��b��*���l�/z�~Y���]����Bj�r��钆[�p��6?��BG,5ƍ�[���}A�/.{�&z�(�Q�̉ي��`��~�J��9f�H����.E��/�6�����3s5��1��[��;�����㚈��"��7�w��S�K
	B�����r��aK�s�>���lPH^(��6�,�YcUk
e���z_��=������-Rh� қ*�du���G!��SV�<�����U�#��1
���;p�ԏ�w�����f�
�����U9~�Ȏ��j$�z1���ҩ6�^EfЫuu�0#s����ޘ\J�^9����fZ�$]��=q̡��6Y��z<���G��;�c�W��]݌���cS��Rړq�H�B��,*]�����M��%�1�c��&C��=�R[��V�9vN*���#$��ۛ�J�I���=/�$=Ek�w K�m�	��q佣���]�?߽yu��{�GW��ɂ[�n�����O}�c�S*8k^��C������ۙ�nS��]j:|�{�c�>�������t���#��>\��(�u�_!8���J!P�O�Ɇ��7����Q�V���.�m�#��}�U1�U���Hl���A����_>o�O�~�=0�˺S#���	���_]�����cu	���[ɺ^��M�����|\GوLyJ�qcz5=%�2ʒ�V�N�$�oɍł��'m-�Oߪ�0�(��.�[�8Ó�T*zj�2���)P�1�q� =I45�	q8�4�`����?o� ���w��]���E�F�k�4��1�>G'��$�X�<�ӱ����f���cF�#Q�3u�sH��+�矕��AaY���@��W_χsH�����>�ֽ����u{�~��ii$��w�x�`o�g��OL�&?x���.�31�夿׶��C���Ӓq���
'��l/�@UlߤkT	3������0�}O<�Ӆ~��++$�Nw_l���3W=�C�f��xA{�I������'��_��f29>*}7Th�ܪ����5����ћ^��B�\u�A1�v�k���a����ܡ6 ��W�Uǯ�C�͡�ߞ�Ef7�1�8������X��K7�;)��=�L�ۊ���
��w�[���y�K�@e�ZQ����X�Fb�Pą����1��i*|#\s	S�����oK{�+ܨ��斀�D�V:*g0�������v����A�R�§�[�jN���jEG�57��3.�p�M�<F��]�GN7�9���:�ӳdJ�O������s���ra:�'heZ�\ۢE�vm)��}�l��S��JWB������K�f4�:Ώe�/�R�rm�,��*�G���G7�5E&Em��ge+ƢƮ4�(�=
�[�j������f��R���]b ���Һ�{���l� z{_g	B��'b�AH�K��d��D\��n�<�Bŭ�S�F1C�E�tpnIw���|���d'��i��v����T�3E����j1��p����Ɋ�otRQ͠�7�m�ظ��Y���D���h\�N�7L������J!M�hg^V�k[���IFU\\o�H#�+�z��Dr��mR�
��9���Sw�܆���SjGԏs�W�Jۤ>ƴڹ�^�V��]��-�M�%����B��G)�].J��M�#�d�ra��z�\���P+κD�alet�5G/�on=�.s�)�h�� �M�\��F��[rK�u�S�M�Ώd��	Y��^�Wd���ǻ�c��X��]����e�6��"0�=֏�z��X�|L �tOӕ�?a�gD�W�H]��u��`-$�����P�P
�2�5X�
�*d��؄d�0�.�c�)hV6/gTұ�J�����`7k^��u������{�/��&�)����uպ9���ӈ��Y�Iz�g_f�g^u�o)���&��.j�o��]կV�"����D�/��na�
uac��*�k��׭�9Y�ll$��p=|EvY��"����$�T�$-�|��L�9��#��SV:�\�2b��k�����w)�W_cn�����-tlT���4��1�6�Vswz��:fK�̸�Cm�|�d5�C+w&6�^�Z�7��3�Ыͱ\����b�ӄ���-ћ�}�<$n�!��Ptr��ɷ7E�Hc�$�u�k�iQv��k���ЭW��q�@J_v�x�kn@gu�s�^Q���"�q�uMp"f;�
�:�4ft).��rƬZ+7%��)����F�s]�'��l�JŸٮ����VRޫFv�t)T绂I:g�ZyT�䣀md��%�m���h�h��ZWJ�ܧOYsR�@�V��+�~��_��2���Of�"jg�'��.�d��z��}@f�M����ֻe
B]m*�ř����ѥ�w�L$j��đ
���M��!�[�fPW�_Niܸ����pj:�ͬ�,�x�s��<Uȋ��3`����I��J�Z�Y��E�R;�Xh���EKTH@��Eӂ��e�"A0K���D�J��?R& kA�"r$�Q��r>����S��S'TE���}uJSM��M&�.A����yy��-�C�h���ڛX�Q�]��΍6�-�lb����|y���|~�������G����g��_f��k���ׇ�T5�֘(�[:�_�y������}?��������~���~gmcZ�E|�j5A%$DIZ(�[qE��C�,�}O>?������>�o���?_��s?�DD|�U��E5��Aj�V-�lV�Z�a��&"g�2|�U{Ϊ����6��睝D�5N�#�u��'F�������i��v�A��M�h�͍]燍�:�7E��Z4h��u����mۊ ���n�q�w�{�e'UX�Z��y��y���sn�߇0Et�,vM1l�n۫(����6�v=[N��n8�J�່�Q���4��]�Z��.�T�Tj��Qyh��h.�(#�~��R^�^��]Ë{�`�

)Q�*u�<zN��7�ۼ�݅v͂�8��(��fciN�df�v��Yb�H�wuO����W�ffwn�|��1")`�
�y��^w��;�?�/�`r�&4"� �������������I�I�w��Dn�X��G����^}��r�7�S$T�-r1_��'[F�y͒�^��=8��baS�/"��o��CGT_6<}�����~�`f�P�1F�����綅�3�sMP)����cg/#V�G&�<f�)�������
�H|>O�0_t��e�� DI��\�ε��x>�Nż�ۓ�g+��@v���}�i~:��kނ����2g��RF�N�LcyU�6 ���������F}����D�w� s�3�~��*|y�z��i;��G'`�Ds�S-~���~馯����{Ϗ{^F��$8�WUy����f�Z�h��������H�
z��審�4Sso��i�b�J`3�5�q��O���?##1=ύ�F�خ��hg!�ؾO�; �:������B���*v���'��>�ǔX�F\�4K������w�!��\jh]P` |�_Q����V��|�j �e��t��}&2���|e�<7#b�_���O�{�mz�1d����nb��<�v�텝�-;@vV���p��S5�y3�Ud$�8��K�s�$ӎ,�����^��nH[�q,����R��uҬ�S֥:Z]\�y��ŞbV�ҽ�����Pb�#����mD,�[V��wӲ��^nh�Q���A�۽�d������de��m��s��'��0Ô!��*�xxM�N?B<-3oz�
+����4s��H�@�6�PsR����[<��� =W����=_<���y�i�}�SXk��a^M#2���T���vxŰƟm!��n�={���ʃ?c\s��SƤܞ�SLlz���oL�>qXe��%�3s�xk�R�2:�)�Pr�=��^M��?*J�W�Yk}W���э���qP�z3^�,�kVh��^2Ѭ׹��k���hUv�I� ��5K끥�^�>�wNM-�~�hX���������72mF��X�Α�/�0υ6�1�-�h�\;.����T��ЗH�6m��c�6�J�[2�7�W!_��-�T�3*{_AP��B򼲭��r��z �z����
�g�b爂�"b �V �G���K�r�5lk��b �Y����R�nf�m�nE��v��gC���=]�)�0A\����u���s뾈��J����r��S���}�$n���;�p�����g �����݁�>�]�xZ�.�7��	��03���<�;.S'��FIu��-��8�_1��`y7/j^���y����X����w�ch�y����K������A��3��^}ɂk�����j�!���[�<�}O��1.^��ŭ���]�ׂ�iL�jF�6�ucʛay���uf�\F�NN<�Ӳ`K/[�g{���1�!�8�08D�x\�f�_�0~`>0���o��������Dΰ�
:޽/?:/~��0&�s]�V����rʮ�1��\ӎ���]��rC�5K���ql��%��W�/��+��s��zN���A�adɪ��i���pݸ�/�I��(�Ơ��FT�+��/�,�K	��V�H���i��y�<��N���U����G��a��/�(o9��Lss\`sB_����6Af;?��{lN�����,���)��𯟙���?|���&ϼ���l�}�/e��UIjbڽR�ʳ'�J�
�|s�O��Q��ϲ�=hR���'��?*��ȵݒ�<.z����_��GgG;�2�)�|oP���8�ZW�#������lw����nX�ت��45q��^j��TV)5���$�w�#W��#�F��=��/�> 4�/5����h>�-j3�ޙ��З�Ǟ�B`6����U�)�-%�<� x�;u��\�0����:�kUKK���r��WVh�;j�-�p�eD�[^�e�G"�O��;Ck�/V���}�a���n�?~�X���tk��a���e��F;pm��mL�83��rM��i�c<�M���o	���x�\5X*��z\��j��є�j��Er�u�r<�X��wv�hF�j���t�AR�U�\u�͵�Qěf�s�Ѳ_UW�K�d0����iA�'�W�d�9L�K�nf��ӌ����'ze'ң�x�j����y"7=Äe�,:�Y�g��E�3CϛĶr_��g�lNu�bg�߇�k�>��j酫���+�=�n�����~�u�ΌjQ�/�$��Pܥ�5}���oJa;�%���Ojp�VZ�&Z�7����,�T�qP�9�F��ס�񐨇Z� oS8����Դ�ߗ���S�^�X{ ��,,�%�"�'��g�5�jM�0��^�Q�_��M3u�:�ǼTSb�0�T*�Z��
\�������{n	Aa>Z� kP�fޑ�ƆWITi��T�Q�w�{���y�S1������9�x���^:.8�3Ԃv��=�X�����P��Qp�����{w{����20���u�M��_�%��🾤O�\�k\����^0s�m�#�jfi|<v)����(ٯ"��сj��G��l�_������u��V�&O<����u[��u�A�=��iEW��[�2t�OM�|i�� +c�v�C���7߄��Vײ���dh��ʏ6V`;��5Nq3:�5P:v[.�Cmv��tӈm>�e��:a�M�G���W�2��ʉV#vv�+���7:=W�RK��\�s��;>�בν:��59���M��s;y���U�ܘznF�B6~@���������u������+���>$|>ŋo�w��Y�5�4�C�)׶��&�		o5�JV0p��g��䖯hl�Ï���E� 3�?z�����ZeA;�uN��O�e!���5*ӏ�a�t�"�ڦ���"��W�a��ĶB��}���:�8g�>@[B�ݿ�ے,G.�B\kT���O��A�q)�����/{(V.�b�Mϣ��Ҩ�r�F��X�Ӛb˲-�KT�����)��z��׎F��n �s{���Dz�1,
���(F��Ւ���ꢏ謁@�����6Mh��*e{�4�`�Z��3����N���k�����M5a�X�D�jAvV0��k�/�~.�TA���qp/�["w�x\��3y_2��ܾ�=�LJ=Mͷ�3M�M��D��g�����as�O����c9���J���[Û��q?n^M<m��;�#x��W��h*9����~k�;q=a�x��%�ݓ��mg�]Q�u��KM��_���ǆSy:���|M�eT�Q�K��[�;<h~\��;��ÌT��@���?�w����U�hO�I��5�dW���5p�D��v3�W�K�L����㿸ۿzhѝ`�T�(�^t\���f3jtf���1Wq`e��M��p�RuX��h��f��P6�ZUKƩ�������J|��s�`M�׬ML�ѫ�H��a',�u��k+w&���1�}��-v�����e!��E>@�)�ﯚ��m��1����!�~/�&�.}O�B4Ǽ�8�]Cl^0�gU����O������ޅ{�����D�A���d���xnl5趤�#.C��~OyR�S�i�[�P�n��"}��Y"/�}}�
\j�2���?�@�{�G��$�'���e��{��C����)Sz749��g�>mje����w�c���4T����C=�P����+���w3���ۻ������^N̠�^_�d�5�xL5�Jl�c0���;b��Y�֊/���쀎[���c�V�i&1�X>-p��B.�f�3	�%zj>����~���JTJ�_��������
A�����11O�0�!Ќ��ﲰ	�ڄ~�j�@�2��2��aəf�T�ZQn�l'�?ȏo���{��)��5�,\�(����ʮ�{���y��8n�<��Yt�[4�r��r*�/���j�Qݧ4��`/���|Wy�j��,$���PPE-��a�e��j��6����Z�yts{#XE'��S�E��:�׎�u��$õ�N*�{��T�X���+/�g��Rw]QN��8ܓ&�n�E1�b������pr���.l�X�s��A�jG�#��*;b֎�O�]�|yT��g3u�r�Kv�HrW�9���{U�ٛO-�Ԝ���b7A�A�9��u�e������W��y������9���{x��HՁ��0��s���T���{Л���ٶ���z��^�Ğ�U���o�������^�\6m�y��_o�̅�lJ5�l@�bØ���
��#����P)����kj�urK�
h����y�nh��M]��Z�v�J�8^<�E�ҧ�D����k.Çʧ[ѽ�/��#���A̹��.��d��oE��]��P�6�i�E]z�x����Wك<�g8���<����p�kԂ8���yTS�ߕ��zdVX˳QM	�U	�w��I���Z�W���^��}u�G�����zx;>>o~�L�Y���o�9"���;j�D�"-u�]>�PI�����u��ދ��PC@ Lz����4��p���|p���@��r�/W�Ciz�ے7��os_�s^a��.��(��n��ӇV��b�=�vt�]{(Ac#!���G�uNG������q ���$��Κ�gy�-��Kr��l��Er��K6�R�g�s�	������x8w(�[D*ȻƟ�x;��e�7���:�����|��u�[#X�iѧk{k�2���ɫNaՆ�wT���&�J��:�_Rc�]�$��4�#23/�Sk�����3�m�O��}2[�%N�E2^��aX��%�(���ʻ�N�����a��k1,�qܷ�Ϫ���7�0��M���ҊNג3���_})����E���
�@�~��"�B�]��l9�h�PEѷ�r3W\������-�I�Y�q�!�MÉ0�c��TST=����ܖ�J,*�\4��.7�P�vg��^Y�G4��������c�V�F��Pu&β���g��9�jky�+���@�[�v�҆�|.��F� Z���&� 8��`�Zss�����y�š��d^$w��ޗ�p3Y劕o�������C�q%�4T��Z���~j)>���u��x��2����#d�?^f~no��~�w��4�uK�m�D�6r˫$�\3VZ��c�=1L��� E�*�E5�Q��/��8y^�G.�S���m���m喽	~��{�:i�pM�L&�B��������mD���שMҟ>��ģ-��?$����?g��я�C���m�n=�e9��5��C���mo��ه#%�/>�a׊q�������cw�)���,�y:�_
��V��7��]��.(�:y�댱�K�1��,3�)��x=��g�
���ȅ�]� $d�SN7�^i��;�� �7�˒�{��z=��S�p�H���L���Efo船M*�pK�e�A	E�y,��x����c�H�|�toCNwY;�z����å��]2��V-��WUv&�1Lᑧ�,̾Dw0m�d�֙qƌ*D�E�ʄ9��^�3�7��<��< ��Υ�ף��R�"NuO���*��EH��|����f�d�EzH��Dж��^�6΢������������)��@��� aM!__�,�ϟ��ӈ��Z����w�yˎ��$�����]�PC�B#�}+�TI��z��
D|�������~�*�^�ٿԏyB������1�]�}�b��$��}�!~�R�SO�_b�?z�7��{�N�{�xF��|Yrl���E;�)Ec�79h�7�(`�{߫�*�e{�(�-I�aq���#X΂�8�Z���Tl]�v��L��� �\D���m�EC�v�a�['w�x�~B�^�YQk�I��CMR��������x�0�ͤ܉�Ս�DC����\�R�,_����/ĕ�*>�ɉ!��;�;+�СM5�,^�Dߝ:S��g�����9�*I��r���T!�b�xy�cw2s0�߶?}�ey�[�~�O�oL�M����sS�Ń�+��n����h�c�yk�7E�OW2񢓻^d@L���5P�!�o�u��;�3.��'�;�xӧ:-s�V��Ý��֪G�nb�I����Og�{��y��mnp�L$\<62�1�G��}�NR�t��dT�m�Ӑ��*�,x�j#%N3,$p��Z��X.<���"��Ч�-��r�����W��|<y�/���tP�s�P�Wo�Q;	�q�Mǔ�d��m���l���,��%O���o&���
1�����h4F�L���y�t8�Q���"��YQʹ��U�z0���WQ~��,�	�7��̮u(/�9d�T��������ȍ*t���Z^��_$�,�zŴ'N�l�&��t39�b� y���2�&"#�[�~�y}�fD���ms^8Z���n[
T�7��:���c.<�E�L템hj���ر��~U��_��ZS���~9�Е���#�5�y�-ם�%��pND;_�z�����V*O1�1��c��<�Vu���-45���=���0~���}��\ ���K�}�Q�vǀ�a0�>FE�
'�ae��(�h��~�w�;Z��T��Ql1�]�����G�����ȥ .�� �zך6a��l�i�9W�������q��c3c{�̚�5{;��f�@-�"A�͗f?4;�h�̲m7E̫���Hz��c��#u�*��j�����O��۳8p��k��i[Hw rVf���vWM<����m[�)��`n#��w�C��r�mi�$���Oh��{c+z�fj���q:]n�m/�چ� ����ھ����ǜRt9J���T%�Ǘ����8�k�Ҧu�	�xnԛ0���b>H���1A+��X���-�6f۸n󞻩T�����A�旘�W��^�"TkAUĤ�v�PJA����2�y,�x"h�����v�kb��9����8���/�cIL�B0�M|�teL|�t�쫾T���=�هq�s��޹"x^�)bۭ���b�S���ݲ�v�MO���B����Z�ʶKyXA�@��p�����M����Rv� >vF�ݘ�S���u�Ĺ��S���Y��ش9��)��z�K
��i�K����;��o�9(.�dr��q��}W�	�F#T:��RX�%�.K�rۡ:ޭʝ�d� �}."S؍�ѡi��.e
B�=���gzM�cj'���ӭ�Z�5v� ����jIر�sәwr��Gp�㫋9C;�>�h��V�s�!�;e�ѵ����uj�Z�w+�.Kz����ڍˮ�����*��
�yu�Q���%X�3#M��T`�/��y���y�w��R4`k�j+�7x[�ڦ�#bн��<�t�[onWNY�B�QCP�\栜��7���,U��"N�%�-nw�)z��GW-�^aW�������Ь���� R���Z|-���,�w6��q�+�"V����@�.u�nj��̧S1�(eIĳj�?�*�R���
ʸ���ɤfiD;cG�DMu6c�K#�f�&����NZ��7`�����3�U��el'Mݶ�֜���je��Q%����z�p��]lɚ
} �ݑ�Yˋ��"��7�go�u��Ш+)��Y�i�E���L/q..��g93{���ΧJ`ӑ��ݟG�g*�V��%R�,�M"U����̹�vElx�C2C����������?"��jS8*n���ɭ�5��������vcw����dQ�GsM�8�	�	�ܖ-�6h5��_Z5��2��mL�#��^>Ew9�Mp�K��6��7^h���i|�]������8��ɲ�uuѨE��s�XJ��V�=��G��F�����(�̲{U���Y�dZos�Q,�����5d�4�}�z�`��M�#�T��Y�t6�A67vܲ]�]�T��/.^D�S�6�K��s�CBv��Z�j%���	+��6:S��Y��Ť�o.�������i�9D�6��Kg���|�^;=��9��h�\�3�s�_*�sb�9wT��vu�i��3B�'��g^��DǦL�⹓����kڕ���3����Z���(K�)?��i��m��+��ƧF#X�����Ӡ��_y���O����}�����f~�ߨm��	�}��:���/�=������v��L}|y������}>��������g�����owE�c̞��;[Q�v:j��#��m4h-lLE]����l�}9���~�_O����}�ߣ����~��OӬ.�<Wi(���(��������U���;fU�חm��c�;Íy�*.�'l]� �Ed�<��U�j���5�=Ƌ��F�ō�h1�����6������C]�FM���)|�1b6����5U4��m1D�#n��b.�vrM��6��m"~ ��(Ē�1�ͮ��4�խ�b������5��5Z�k;��\�∢+n�����UC5��0L]���U�n����rn1D�ΰ�������F���z2�)өO�6*U����j��e��;��jv#�9dqQS�[��?��`���`<���\����|wA�����1t��<][_;i�Z�z�gC��f/���[���z���{�\�g�ߏ��i�ʒ�暲y�_;��Ҧ�fOBr�HN��3���'mߑ~���uhjc�
��el�mx��T�s
�xj �+�!J�����tPK�x���~�$Ա�uctn��HƝ�L��yO�+i��u�k;?��]�����c���OOF���� �M�ʔ���꬜ad��\<)��
��~X�=K͛�j�����p4Fǟ˷H���k'6+6P����0Y~�X��/�����h��U���9�1i�_�P�+7Cn��9*`�v�Otk�����^���p1�J�ǩr���5�t�M_7�
�T.se��LK�0J;�q]n��g)�J�R]����I���m��A�w߶	���7z�ix�/sYT7��.����{�x�������x�m,	/<"��ϡ���?5��nA��~�u��ۊ�m;JJK�fu�9͏o�|g��C��OĜ[��$���~?�[i�O��.�߯*�-��>��&�Ћ(�D�U�,����CuJ%v+��ӓf����11o���V��7��@�٠O�B��@�{ʅ�4�vq1u�-ų �%��m7e�{���i�Į�m �T����Ӹ��f^A܂�.%�/��c�ݝ���a����
�F.%jB�؂�_�w�,��.2��j:B�^oE׼�>.��PШ�21��������ȊG����D���=W>�"�i}9B��ܗ��(��?<�y'��d��UBG��K�������'3.�x���`�W����R��[&�_��ݸ��/^&h�p���8�1F�t����E���ח},�Y�E{^�E00½S�S���qU�:�K���h���H�{��8��Y��n1�w����zm׫7��^p5���5���w�+�(л�zPv�}k;6��M4��0:N�޵�K���D1Ɂs�m�#�\80�tD{!��T".<�,[wuw�1^�ަk[N��Cb}��tK��[�jK(Vj�:h���PwA��QX��X���$�s�ΝM4����(G���݌���n{^Sn:c��b����o6׉U��3۲�:+#Yp=[fX�=e��{)�{� PO���{vz�tBO����b���������Z�3�uH��xxw�cU�ֱ!Fk����|׏�!�Y������rz�Q
��;��	��~���1^7�nw+�ݭ��lϞ�י-�(�&U�>���}y�tn��� +��2!W�٤i��*��,�Qc��hC*�]1}�-�;���]1���M��e��L����fյ�:�e̅@����{''����w�ojc��"� �D6��k���<{�<��?����mL��Yr�[�,�;=���}��{����c�GZ�����j��/j��r����!����j���{Q�+�kX����Bm�ؔp���� V�;�t	xM�0o>��|u
��م��H��!�+$M�qqC����Jd礼� �::k���5�$4���tW~��M��:��1d�^��O���ϓ�bT*�����k�~�Q��/�I`������ͽ�9��>MU����9�0C����y�)=	��z��@>G7�T2�=Q�^8ހ� ��v.F��vE�2�u��9��zB_�³��F����
|�N7���1�E>����WNu�GY}�������>��t�(���>�#c�2|aP�MڣJ�snn9�-9���L{�ܺ�]�*�-~oܳ��^��t�%�a��Kߛ*#Q�Π 냅³���{e:g� ��㽏l��{������'���Sl
��:4�����3�Y��yf�d_�p�z`D����Uȶ���fţ7QBEχt۸tj]����36\�N�|wnh����zg�zYP9��1��ߦ0����W�nj=���XU���=k��D��@Z2[̡]�ZI;�(�>�Ί��*E��P&�o:g
��u�y��j�e�Z���m_�:���\��K��b�Ni̽�)sތյ����͡��y���=;.�bx.g����Ϧ5��h�QL����ך������h�+�kH�[N#�G�����ϣ�y��%G��e��Iޖs��!�]�CM��J�Vת���eڠd���C=�i�5UqS��c�*oR�,��w+~�Ǧ�殕�Bf��w�/�+� ����Z��Ԫ�f��խ|�UL����'$���:�f�����-}���
����w�1m5��h��q4sИR�M�s�gf�n�����[d<�03��8�7gBؽ���%��y�S0X�b�U�-QFCΙ<��{�O�S�G�)X��	P/��;�v-v�x�ȫ������Уp��V�z˾=�kz�<7!��
��6tЊ�|��ڈ�[`čǤ�ڽ�Soi�߮\q�c��2.�n|Ԇ�9q^no"o_�e��O�
k]�}:����E.����2�_&�"PI4�U��Hx~g�;"D(��/<�h�����j>�s�������q�t�j]���ių�i�ӍŪ�����@Ƈސ��r!'�_E�*�b��6�z�v�cc~�(v��Yғ�;�2;���^Tu08��yV��
;3_U��M@jY�@�2�`�j��Un���2�hj��.�;�~�gQiN�HG-��n�Θ2�衒�r�7Ox]���4��[��V��X�330 �|I��m~�<�?D�ڻ`=�U{�a��� ��<��~��c��8,��ёW'O�s�4�����S�HѮ,`{���u�5��~��J�H��(IoE[M?����{�I��)��e�ؙ�\5ٵO���YCm�m�H�bR�.+�j];��n�Q��-s��/"��V�fO>)�=���72#3��=� �x�?�[>�w�zPۉ���\ق8EDG��*�Qb嬝�&'#hB��V�j=R*)����+��ٖ/R�
�ֆ~={�1Q9�*�����m�;.�F��٩\�,��5e��
'�c1��MA�S�Z��UcƩk��ZS^��;���xd̷ؕi[B��l�4�pˢ^���f�q ٬��Us��k�v�l��7��{�D��oBe�kb����Sex7�vT�8�we�������0�����g����nc	H�r'c;�+5I��*v�Õ	�����.���a�C��K�k��*n����sX��3�k��]��\s4_H�;ϡ)�^�t�4`���Ҩs0Hn{�E���O�����_�kE�7���K�@O,h�Wu�Ve�ݧW15wD;ĳ7��w���4��+C�>z��u�lZMN�g���/�r�H�fU�P�
|2��sx{�xgi�L�������$I�\--�n�jI{Fb`D����-n�I�����W���y��{���0����z8o�T��;O}��1�	0��c�C	��]�\t�^�7�W9�y��`�
o{�]uW�K��0��0�xq9b�8�x����$u��3�߷"�ɋ�·����r�ёQ���{[����c'����}�Sg>;��<F7���|�]�*��Ax��Y*vGtO�L��@f��c#[�9��3� �=?�hv���5�C�BD�"%j-!yd�⢽�I�����S�6X3��׆�>P5Z�L[��l0���/Q�G ��F-��qf�y�v�͑>��o����̠���;O[Ѭ2�6��`���c
�N��,yZ��Y�K`L�N��x�@�B���m$+׃g�>�*4��\�#����=5����]k6���ћ�l��ĂzY8������Me�xө�ex�٧c��a3s�(E�N����LӺ��>gQ"[��̇�)���n-�(;��2�lXS�)&��[��9��q�kT�ϵMÉ�1hdy�&�pQ�$�ކT�n��������E]O�t��=�7���K(��{��W�/&�ӌ&�&z�j�mM���˩�8�X3{�Y`l#L���a
��ʁk�����g:�@���硋�"J{ջ-q�F:�]S�L�Ǜw�n��T0t�M��i:�m��0�A=k���/#w\^o1���C<���3gT�&a��}��/����V��C�Gx�&�2�e�aMAnK�����B/&^,�U�5�د3�O�6EWB/��n�	������xrc�3���~Rgk����~ww��ܢP�㳰s�^q�4'�kTַ4�d�ޙ)�(��W��;&,�$��i�4[ o�\}��ӝg�︢k|�ҧ�̺��hb��ӊ=JnH�$���6�7��;�MNK�}@��j���Y7~������<�����C=Q��b����b[�V+��hCkt��F���_<b�|��)7.��#���x��8�}��M�[�>������ݽdG�i�A<��eH�f8��~�\�
2[y�a����]�c5F����ݸ[UF:��g�+��'�^�E�_ՂѡZ�������(�q�T�HZ�:�U��;�3}w=�u_Z�Ml�ɬ�lhei��^�*1��K�)�d�{%Y�m&L\W� Tgo8������ݰ�D7�}t5 �����׶9q��}B���\�x*�98f�����<C캺ݑ2!+mM��j�W����m�́�!��J�v�\�u���f:c�<N8��The���]J6�ӲK5S�d'))O_2��R�xz�\��I�sx@���&^�B'a���)��!qM���]���C��3{ى�E"�ٌh���M	v���^a�e�xR$F��d����F6���w;z��E����+������OBz3O�AU�� (���w���B#�8���8\mA9XyS'�V��=_�׼� ��+�3'�q������"Ą��4�����s
���xl6��+��R�wE��8�|`W���F0[���1����`ƅq2��ZAA�E2}���7y�;�M�{�3^ƌ����@Rn[��~�� �Jh�d&��9^��X���;��\�#����i�ɂɂ�R�Xv`q�s�h
���Ιb�V�="^�L=G�[׃p3�*n�z^�:��'2��y[��w���4g֙����x߶̞�V�fEs�шM�_5[x���\j�s���(��aA(��/!��;�jEЈ	�le���!�r.mƵ(j�ܗH��S��9�:aIT���U[m,�m�L�>5�!��Rۚ%�n�3|ˋO7//:X�a�*��=(\�}�gy�� ��ɵ��)9>�k�"���Dy/;t�7Vן�7�;�1�=3p���C|ع�G�������W�/>���Ï�k/%���j;�:�H�6�w�)��ފ�N�1��X��u�֗�[�dn��<�U]̾���8ȍ����v	��˰�|<zk-�Ơ����w���F^F�K%��-�)<Ui{��q,�l�����o�6v�p��jՃ��y�?��x � �j�'�Fߎ�ԇg�=_
'���^�xM\'�����+I_�v}9o��uk��] [�(~��	������(t����a�z�Vin�\Ժ9��e�;\��t���'"��o�9�v?yP��l�.�5�;B㰟��mط������ڼ�0/>�w�3�,�eAr����є�ؾ��2�����^����cM�%��|��"}�S��>2�26[X�������x?L��@����G��Cn�7kU>��
53 ;@��-B\q1�͒w+Ϻo=cG8-�pH�>H�;ߛ��(�g��:9�:O.�wZ(����Z�`:v{ד�/��;��J�~�0�z.Y���sk��2���Y�Mۥˉ;�	���ӷ��MG��Xm���Ebh��nE�Fum�����yt�6�bZ�YN�Q�x��{���k�2�&І����\���8B�sJD �H�D�#0������½��۬���<��	������*[##�R�wF��߆W_NyI����	�e�^`��N��JWt�_3%k㌉8]�z�++IǗ%-]����Վt��ӗʘ�u#=��3����<�r�`7��~o�Tz���PYɰ"�O���d+&��\21>��,nEn=t�X��8i^Ɂr�+�GW<,z�˟�E'�����J��3�_��2��^�z��Y��}7��`i3]�޿����R����$D�=���E�j�Y�6�)F0���7�U?��*P���>�S/�G`�Y����lu�ۜ��ǣ0�%��{a5O��a��\s4�؈����v���9y)��o�e�ȷ�v������x�ԅ2K��ߺ�������a{Ҏ�)�76��&�D˴�R�j�}(�D\�tf똈[O�����X�l���,���;����ZC��a���]7�f�}TF=�@�F�Lq���C+JI{ʂɨ��b��g�i�)�����fO�*o9VU�{�3�Owg�w���
t�eH����B�u�=ِ��_�b-��i��m- ����d����ٙzy��Ո2g�|j��EE{�����)�q��,��3��ų��I�R�&��W���E|��L�G�^� a�ߨ\y�Cu�,ȝ�z�0Xf�`^k4n����$X��ܔ`�UfN���a�����S"�;E:Fũ�ɯw�rÚ5"�3.������ ��v���}�d���&��s�]�U�J�6�Z����Z�Ci`���B����ؤF���#&��)Y	�s�q����)`r�G�:�M�[�q����� �����*)�iC�3�+6".%��j��R��Ǖ�R�6ze�U|�h��T�a�6��L�k�N駮<���.C�b�e�Է9�*C�[��X�>+C<�������`��{��*/I�y�$UI����ϐͼ\�z�C1��WF.mb�۲�'ӵh���k;�wV7:���H��a���f ��O�R��*'� �����19p�ě����6�WO�c�d��|Gpǜ�W9|v��8��u/"�7���G�7ON�c����R:|,�����F�a��P���N�U�O$�:��e��v-V\r�sU8��̣Z��S[ɷf��]Z���1ۇ�lh@�b����Z�T��v��fA���1`�AF�t�)t'p�ר���l�y7�*v��U�|I٤A�p�����]Y�n����HN�}c���T�&�xS��u�1սyY�d�O@���xf��:���*H�7��-s�c��]"�h�Ю%��`kN�Gi�hbn�Yp�T��$e���G-˹n�C���g���q���d��(I��W�Z_ۧd���9�n�0���!q�m��3Ga�:�K�Rmu���(��HB8A�]!��m!t9�fu�Z�nH�Y��\b�4�l�;&	}�M�\�ʵ��;�cs��::ы�5mV��ಮ�IC���8�Z	:)��}	�{���!��v���������.1whN鲻_fi���Lm�e�h9��P������F�����`�n1������U;�
_Y䶪��3�Wj�c�&g1l�f�B(�f����W=㬨�U�f�j���4�y
��*[��
����)�8�Eؑ (0{aW�!����ܼ�ȥu� �)�Nb'���7aF<j�h��gXl`LKiTcz���n\�Փx�B4����򇼞u�{����O���ziI�d[&䊖��.P��.�ӽ7et��tcVȺ
6�2������f+�jsg��u[���9����idZ1k�]e����z�r;RR)e�.ww U�VV��
���'ay��r���KEڷ,m���(��N:%��*S�:�ЖvNB +��v�V��/-��}NS���sǖ4dN2Wu����\���+Eٽ�VG!�᥂��]��q�6p�I��	,h�y���*���ڒ��7f
͋1Vȭj��U��̥Eu%�N�pռ�/������9��eC�o�-l;D����o�R�c�ҩ&�bs��&�!��Ha@n+dh�(;��!����h4I���o
�c�1�أTu�Ճ��Td2�Q�2���	!
�˪uq�!ǔ���uB� ���AAV��cWX�4U��v+6��RG��5���i?���}>������}?����~?Y��ϥE(TW�d��cu��U�1LA$��uzآcͪ�8����}|�z=>�O������|G�������I-�i�6ߛ��)�m��޼M���N�""
�+�"�ǖ�lV~��>>����������?_�����b5{=��n�lmmG�_cDEQQᴛ���N���Wcyi�*���F�t�.������um�*#��c��b��DZ�c�5ET_�q���QU�5WX���'�g��U�v)�`�:3t�Mv�Q��ձ�K���DG�%5���A�����EAz�m�Uu���5���)":+C�v��Qln��w�L�V�Am�7�MPw��8�M������Z$�(�[3E�s���؈�.����b�{��n���AU�h"�Fi�+�q����%��y�|�'���e"�	IAXn�h8Zr����b� �*mu�{�d����Z��vv�����ٴz�r�1�%:�M*�lk�}�����8Ƙ�J&�-��`��$D�%/���q���,�������[��j����֗�E����C�Sp�m�-<��tַ6Z�7Ce��s,���wT��9�gOC�]�Px[���G�`q��+��X��{����j�2���Y�Y�됋f�%t��u�mQ>��yfD�@?��d��L��!�NfU��Je�2
�cڗld�s�ܸȖ�^��w�8t��eKٓ;��(Y=��f��=��v@��p/���HN��܆R�ri$M�j5�Q?G�yaҭL���ΟmyGA��1L�������bZ�b��^݁�ΚZ}�	�>��R~:���Ҙ�%e�荎3Hg���a"��@�?m+6�/���d��-�2�Х2�E���f�ξ��y�t��;1ӯ/?�Lh�
g~P;&Z�I�0h��׸�ٞf�ܪ£=vjgo�MsA�ux&�ʇ�:=�p�ڬ��s��O��ɀZ��k�v@b��K�Ck�*d��y�U���)����f`ҵ�OK6$ޅn65LC�3]���9��D���Py�vm_-Q��d=f�)V�-�7�8��W(/4ܰ��a���|��N*ͼ�u���"��+V���ա�h�pP2�t�I}B��P�4ݞ������c�=R{XJ���E��/M���ӛ]��f.5���N�{�Ew����<�1��)�1����s)���ы�aA=6���v�;O�˩��΢.4��f�K�\D;���*=�,��8����ג��� �,�j��.7w��]�,�C��c�wl��ީ��yC0f��^�9Ok�s�%�B�vfob,����l�7�*r���W.r��
��f�wE���{z\7��f�H*�.�&.%حfU��.�p��H-�y�A�y��5-�.5�vQ��
���$aQY�v�K`� ��s��m��W��ĎTe����e�#̋��y�~��x�vm^g�o����>Ρ�<����sN�nӵ�B4�A�OB��h���p�׏���	�S�9_߅}nI6j��C}}��K�"P�c3\6��Z[� ɭΜ�~�H�fHs�Ц��Ȏ�UГ����+q��y镻7V3W��!o��Vm�_?��e��{��nU/sR>���:��v�b٨�A������ʻ�8����-j��>�G8WS -ń��^�Z�F٘9Q^�K���)ʨ�c �2�J�]9�duc�x���XҀ����p��/�,��A9�E��]P�>�oh��'�m���r<��~��G���z�h)n��=ץ��j��v:q�򨨫I���eDٍ�w�o��������©bY�7��C?��A�{�	���м8m���g��*��קyw3��U-�)^н���x�:��;鷗����U�n�1�)u�5�K�\�P�j�퐒�������|(T��8����Zӄ���l�c��z����Gl��V��l�ɨ>y���-.M��	��ܬ���݀���O��xLt��E�����A0���j�H��Y��+֝¶��ٺ����b#R����oY��d�9�Uq����m�c=i��Ū;א��y�1I��Y��gr�Un��<-�lԚ� +2��=�s�~�1F�<	��}���}fz�8���q.�ؗ��O�,鋳!c��l�'��q�t����z̹]��¨ThR6�WiɫPQ�ރp��n�-��ɱ�e$�^��1U�l�ؠ6���R�ɝk4�3Xh��UZ>Cº��N�>a��_R¦�Qޡ�)n@�[r�l���\���~�+3خq6�N���lN���(��G��ɘ��?��Q�p���?8�����Ϙ2E>�<-���9m�$�|Z����⟱�(g6�:gCQ�lL�Mi�
����{\�{�����L���{���v+�(o������+���i��E����<ߢ��T���ފ��nM��!�ʺ�8�h����ڟf���o��|�O�q���3�A��[��^n�o�}�wP�H�Ŝ�ARnVQ99Ic�db�M瑊�H�f�鴃�/n�k�tw	�||����&��nsry-96�W��&J�P�6� Ӷ�ι2Ս\Y?�Uϟzpp ��b�x%�R�r���������8�עj"�\�Ff�k������n�hi�RpI�w���휼̴{c�����)�w�م{���;�����k3�Yő{��_���''��p�����Hׇܹ��	�:X :�f���;x�ʸjAo���}�����ִ�,]29W��0�r_�3M) S��<M�n`��:�;mE�6C�����PJ�u$a(����5�^�=���E�Mf�^�������2^��>�k�`*�^\1ʮT6��Z��n�/U����(PԵ�24З��xɽ�c]r`�C�cDl��ȶ`���HW�z�* ��6ܠB�G�G��z`3�����M�L���x"#{!x���r����n7ox��i���S�*�9�bv�F'3�\7ӫ�#���Q;"�C�®��r�6@�f���Gg���N���O�C�c�E���U�+��bѦ�8�d��nL�XQ[��s5Q���Hm�ˆ,�p�;���P(WDR.6���g�kM3��&���8�T띱5��0��&�j�W�n\���n�ဦZ��<x�#��*��K)�S>�Y�l��\�wm�����:���^��6����!�9���V����"K0��X����>�c�G�m�s*�fG�4MH~��B���%^c��J���{*Kq�ƫ��%u��g=-Q檆¥�ԂTW8�S e�z���b��?���+y��@:?<ΌoF�^�������ԝE!�޹Y��� �&�e^˽�&J�t��q�9�>ug�y��T�����L���G�[7��z!.��mSJO��i��j{I�Aq:�hW�m���Y=+$�}{���1���x	�:w^.eWuB�ϦuГG�Cߟ�R��{i��Ē�f���� ��k�̹����Tm��]U�\U��l|nX�m��l��ݾ�b2� ���ʴ�ͱ�j�[�j�}��q)oz��+U"Ҹ cx�%����pf�C{��ѧT�V����/J=��S��է\�v����.�,�s;Ϻl�M��s�)�U�`4[�24���Z��	F�wH�S�7YѶ�f:|�nnfQ�����X�m�FW���l�D��8����Z�&Ɖ�Q���P�߈V�J�������~�O{�P��7ޟ7�o��W�I=M
{�9����'t��z�����8|݃�ħ�2��)/��F�D^�����#7�G.{�.�?&�i������1M~W��_[�;����<�]�O;���l�;���2�,m��K���6���Q�|H��n�b�[�^ftƆd:/���T���lmwd�EY'&�ϳ�h�^Ԡ*~�}��_b��
ul�?n=��]#�2CD9`�۷k�o���mS�;m��Ĳy�.����>�J������N�o)�kWvD�t<�u^_��v(�o|rū����G�9M$�(��СY���D)�]j�톖��/��^/v�;���nA1^E�"����Z�}��7�}���T3������)��
s�����T���'������B���ݻ�Ne����hwcY�y���>|�nU>{�����pR�����a��_�����(Md�����ɵ��ݪ�g�b^�=<�n9D��^Ž�jL�:kO���;Җߒ��j����^5�����pk��iUq ��/��g�(���+Wzw���48��͚�5í����d[��C�)��@;"�@��K���s�C�U���Qu�{�e�ឍ AN��=mF �Z�^�� C�����"��+�y�������������3���{<3���~ޡ=:��9��y~��vfάM�.�b���Mm[Z���L%{J�4P"����ê�%R��ZI)R�'�7� �8e#F� �	��I�/�`��m���cu���ֵo7�<m�JK�3Y�5��]�{�{3a.!R37��	1�lN�9�a�M���!��nQ㭻��E�H����4T�M�/>���>�\c�k9많ک���x���5���Y�'s�T޽���nT�^Wآ��'Ea�"9�é�6՘5srwϫsͶ���}z�/�3�(N�s������o�|5_��!��͇�2������/���;�+T��b7���������\c�Q�~��#�U�z���sϵ�0��7K�^9�]�үӞ�g�>S_<E��y~Yyѹ��.����t�rx��'8t��J^�d���y��<d5�:�iO;7IٝN�������s�V|	U��E�Nzn�+d������N��AN���·���y�3�JtǪo�;��>�����Ī;
ɕ���V�D�����g�a����<ϓ j��Z��U}�i�9�UaWs�ߠӦ���WK��EsK�ݨ��t�v�7�N�]
.�^���o.]�Lf���9��jw-�[��{�N��b�Zu��&w���Q�q�j\�����N����k$��9��`��%]us�BC��/�,��z��L�GQ&�LA!�@5-?�|�������E�R��_�t�O��GC�Մ]e�~�K]�Y"(����R����9�3}��7����;�!�
�>!m�5�+5�^M����/+g�a@��Î�j�z�֮Xp½t%-t:=����סa�tL��i�ù��9��ٮ�����s���g;.m�3�37-[��hF<a
�����t�#����-
�ey�9ü��hg���hd�����,����9zbWT���2���(���4�[��!�`�D���#e�v�{����a�c�Oᖓ�T����շC{M՞��+.�4L�܍��0��]�� #�!y���p5�Q�\�}�F����)��Y��`��xf���.��Q!��y�;$��ίHJ=B=Ps�A���xUkNΒF�;��m����/�����;���V@%s������#�io�QO�5��Ӂ�A4���h���r�l4�yjg%םm<0����h=��r�)��.a�5-�mo&���]������^��~.�J�<�G)�9';
��-�|�3~���`Iw�So�����'"�f�����noL��U! �{���,�ȍ�G�v�7��3|8�	H�{i���	�3�_4y���V"k��z�`'9�U+��2h�_W!���7�ٳ�;��nUŭ[�,ԋ�����-������>�5�:bbnJY>��p��|j�&�-�tӂ.N]����i܍�B���?MH
<T��e�<�
Fwv%��[Ǉ�Mn3��U�}TGq�w�u/L.}����!�a��S��X%n�����y��Y�q઺Q�z�3�y�,e������ndu�.���C0f�(S@�ݬ�`�+7�82�z�^�\ML��vF�6��O9֎Y!)��KG����G�ՙx�w�Z�]�+�߯i]�GNۉ����
#DS>s?���foP;ި�-T���j⻊��c-�#�%3��^3+���8N���<��>ǝ����ή2(�+>�6��0y�/�*\��*�7��̢�=�G+)!�Q"���B1[�-�S>]`.�
�=��rr*��1P��G@�6���עt��g+k�2��)�5�/F�hB8��`�b�f��D���=�^�eR�Wѱ�Hݪ��ı]*l�TWee>�fE��XӬCw3���E.:�DP��ͻ����VC5Ŵ�%u�9Im�W�����j1�OvѼMY	� ,^�,e�St%q���;.IYR=�F�=Iİ0U՝pW%|Miݤ���+����د5Y�MDd��ܠ����f��%	��m+���n�r�'*�,��x��329W���	jT���Q��[�9�S��0�c�½F��l_��U�����?s�c)Q`��ngzݶѕ�޾������ᕆ�w}I�A�wm�=-�h.�ip����ʻs� JV�:M9�6�;X���[ ��o2����Ov��R����9n���A'z(�SM�R��Y���m1�d<��c�+���6%F�d��jJ�B�uj��ju\�*9���2�GinH벉鴷��d�ugV�<f�ӑU�7)B�����[���b�<af�8ғ9��.�IZ3;�j�6v\5�W��ZX�QY&_g.�tl��8���&�7{{$0��e�,_c��u���<3'*%#�W)o���S�c�p�:���tS$H~�(?K������n^�9�bzŻ6�S��ٲC�>*����Ha��.ۨ�B�^��e�(Tߥ�r�^Ȟ����kf�,<ϕg]�ѐo/g "�r�y�U��}�`��#nݪޖ��VjKNut��E��1:�o]�+9��_R1}%m�	���n�`N�Ib|r����C9���O��`J�t�1��C�QH鬫B��HW,����̍J�tu>�D��bh�#z*�a�Z�P��6�|�+P�@7�L�/����+���Wgp�gM�h�\7��_!2W%�P�z�HP<��69Ļ+.�{�q)[�cz�\�fd ՋZ>�$�w�dN*SU3-��X9S�f��gb��tݥ�#�1��WQ���sR�P9�n=�!l�2����^�x�*w\��Un\[�[���ؐ�n;h�YY����v]�swr�%���	��rY�=��4�u��Ҭ!'oy���ƍ��_l��^�����vӸ]�U��7w)�Hɚvv��s^���j.<c2j��{��y����6.��K�eeE��hB9���$���y2�oƋi��\��^�W	\&�y)}�C�4���Mk�]\e���M��f96=������4m�˵��I���m�D,�3��^K��V��zޛ�sne6�K�����:5f�e��H�o86��)	|Y�V�H�O7�J����of�;x����� ��Fg f�6L
(�Q�������tsvՐ�QGͫZ��E�l4U]�c�ŬW����Y������������G����}���1��KQ� ��LZ�N�f;m�11�&���3QѶ�W���>?_���������~�Y��־}�(�X1�Lpq�S;��Y:
ԕj�W8���ݞ����>>����������~?Y�ߵ�V�*�SZ�}�UQEt`���� �i;&(�ݎ�]Wh�g��7����j�m�QZ��m]��E�u�uGT�l:ִk������11QE1SF�A�эb$�gzٶ�󸚪
���I5IOOO]��VƵ���:h��L[�]X���׮��57�h��mѻGk���Ѯ���j3�c~OO^lQ��JGs�mhڂ�:�E������6���E�իGZ���[`Š�Pe��SE4OZ,kh�,E�۸�f�a��ԅ]i
���:-��[�"8��mi���yw��Pz��k��#��ړ��+[�:�5�N�j&-�G���4�Q
��RM�>弸.�������Gb�nv�1����ř��+���7p�#B����mF����s��_��:j������|3`>�o42�>��1	�� �cC+��wS��I¼c)cLs}>&-�����`7�ؒ�	��᫅z9��V;z����b-���`1�[�w����.Hm���ϜhE�S]�Vڷ�����r�f����ٜ�k��Ô�hW�u��,���#i~��E:R�0A��q+
��KA���7
omy�d�
�x>���^ ���=�g{�&;�|g���0u/T�,�|wg.[}|�h���A|��nqJE���_S6d�	��>x��^�LwT�� '�0�N7]M<kfr���#��ή�9:���[��џ=����-q+�)8�TB�9����`ۤ�� �º��+2in5�E���0j�f���P��x.Ӽq�A/$�ng��ʐa?�
��w+��U���Ň�_�����@���飱��D�.���`���Nk��Co����v<f�|ʒ	F���Or��J��z]���u�c���xآ�U����M�D��-��7m=���L�-4�%xn�k�ҧ#{&S�*�Ay��}�!����$�E���:Zs����GCr[�j�Ud�����z��NNs��t.��T�/�`L���
�;�/�Iu1}�iV�Ud�R�{��w����jmJ�ꈛ �L}6�����������scл��Ɖ���i�S�;,>Ya�(�=�:�Y`��l}0֙L>�8��{����+;���7����E�_���^Y���� %Ʃ>Rs��[|��]��vk��=�E�D�R��q����n1��^��Ū�>����� F�yN�j�*O�= ؇��϶.�e~Y�?t�ec�l����m�Y�"r��{J���rg���2�cR�(��hfTY��M�I���t^�ptKa�ˆ�0nf5�#�T0a����f��g��p�[Z�J���Y��V#z�0��}���Ǜ-�BL���<�C� �4�Ç��-�/(Brur���޺,�Y��{��Bת9�o�񂝀H{�S���xo���6ߝ���y��g/p�8��r��Q`��]ږ�H	�<'�#����*�٫D뮀I�=���b�\�6�����y�]d�jl��_���+�c
!RD��%!A��n�~�hL��d�l��d��]=p~��&Y_P���h5>|�UP�BO��nv_k5J���u_�E��C	s��m+�����Z%�����R$gi�=3��p��W^�詿BJ�<n�%��~K�P�P(7wt����c?~�ۀ1�m�DL.9j�Gl,�j[>7$ՕX�40��C@M�Z�n*����q��m�,��ߜ��pT�M�u����X��=Qs��n�z��=5�*�V/o��^;>o�VPt/o��
���r��r��h���v���R���V��5�Q>�[\F��Ao��ڥ�#���ȱ�Ջg�H#I8�\5� f���K	�ܟ$n@r����Yi�*�'���g~`��Y�Z8ho[p��} ����g�}�p�1[�l�Ь�n��QPk<+s94lli�x��DrS���2�����ta~�R.�j�[j#�z�?�6U��j�{��u��$�P���O"
�������('ܯ��$��t�1ZU��d����5���)M�5�޵���5�u��M�^��3����X�S��5� ���=�c��.S-v�vow9L�YhWﾪ�5ݎx�3�������>2I��J��c0��oi�η�޵�|{��W��o�:'�}O� �{T^cg���^�]>�Fqh�"%��x�h��w�[Ӥ^nu���><�T��TXc���4&=���	#�$NC�D�l%��$ϔ �l��F��ܭ�;7�h}p���Tڨ�TF_L9-¹��	��^�bj���N#4o
pC�`<���US-���Mz��S�Q��j���,2�ꇽ�4�����Q�\�iQX5c5SL�׎9��gZ����=��-C/"��-������/j���1|�J[�0��ma���7n��^~K������Վt��w����6��J�k]*~�X�;��iߊ����x��+�Gj������۩��@k��n5��!���B�����wiF�QW��pk�=�"od��a��ޭ�O�*�|��_�o�ɰw�Lz2����Iev���6�;Ͳ�K�����$�5a���s�6U����ӥ�F^�;��wF͢�Mt�p���R[xr��S��7��*������]Iu,�[�/׹��ݳ���C�WH#�|av.cKC����6i�׎44�;+eY��)��ы�f��Z�q[,�j3� w㰁=x�h�O���^Vb��"mw��ĻI�=�|hx�]e���Y������yHa�z�=>�Qi@��+WO)��s�w��#��l��w��T�m�p��3>�e��h���j��}���U�~S I9[bh�(3����L����0�XtƇn-cL�{T�&QO��L!F��S�F���)$�P&:.�D?��q���ffe��z�[���3<89����Y�j�c؉�d���>��k $��2�����d;�͢��:(���:/��;�az�40cj�,�[m���}>��9Q4�A���^�����ሽ�M6S*���EǠ�X��Ǽ'd����@�cG�W/���uޜu<|=�9�a��5w9+"g�^���L�zLf_t��S�wS�T����A���� 5K� ��Df��U╙%��;��D#�QųU���xӄ���B�lŸ��y�a.��x�Bvr����:�=׭L]E>�Ak\�١�JKuZ5ﷷ���Pj_D������������i����{���Ǧ@�G�NZ�/}���F������B��;<�MjƏT�-���f*��j�ƕO!CӺ�v̝B�J�hP��He�߾��E�A�WD�Ү��=�� khj�]
3�F�<a��"޷������7'r8׺ҡ.����ڠ�㄂l��i+�:����S^5�Fi�vo��E^�5�H׎J�*�k{
���a]�3��{�^N�Osjٗ�"�����K�P�`���a�,�Y�}��k�(��E�rG)������'3����q5�Ih�����Z�6晘3^�W;��I��L��51פU�=��4_[�(teH����}�,��������B==���a�z�[��&*�N�j+��H��@�&g3��%�;-je9�j���Ē�������-{�`%Q��c7�^�<�B�͊��>V���<Pn��S{�f\�iv�Q�za�Y��mpn����;B��ڙ�f�(e�>�V���Yh���YDP����w�V�t���76Uȥ[�)�m����י�����C�c9�L5�t��z�'�v�<%�ݙ���8-+$��
�_"�`��m
��
���e��3Z�ݿ� ~���!�G�MT�����f�dŖoFr��v\���F8Ҳ_5�(��jn��ּ}~�yLa.�ً���7�o�B����Tg+'[��`����^�?g��/;+�\�`�a̅�}�.�.i3�goS?���ͩu>�}-N#�uLg��//���x�Y� و���={�ݴF$9�I��E��H�
�lЍ2�|@L53�c[i8KiУWW���ñ�H����(r��&*q[)F��t��d��n{��Z��<�����ˎ+=u��A�fJĮ/
ȝ�WU���<�����N<�-4�AL�}O}蚆>=!� ���5=�i�9�ދ�����0ש׼84n�`��nM��n]P��V�A�4�u?�2��mm	�8n%ޠ�j�&���֒N�x�\�t���ږ�Ě䅮�{�^	��c?h�-z�+�ͥ����u���[Y7Tf�T3�Xk�Ռ}َJ�N(vl�����L.�ȧd�i����޵��c*��#��Yٍ��Y�k�1ٮE� ņR��)��H�*�Ǹv�$��Î�'ʣ7����9W�(��ԑ{����7�2�ls۾�syQ%��o����_��X�//h��������8�

�`^o��-힂�6��#��^<�9YoZ𚬛��j�ѯKD�x>��s�O�EL�oH뤌.��ӊBn�]�Yˇ����X��`�n�P�_��S���a�ū(_k) ��k�|�:��l�jx�MJ{�͂K�>΋���)��J�k5��c��Y��;�$�l1�	����a�����Xb�8]��I0��tu��p�`\�l#M�!���0q�ٰ}���h�cA�G0`I�/���;��ڹ"b+Ό����o1�3�y��7���!�����C6���d��\_s��SeVz�y��3��EJ�� �2�ɪ����K�t���=o*�䧋�5dy�t���v6�T�/>\�O���L���#v�c�[�8M�O��M�b��ݑ���Z�++mMݽ�'�V��jn@��ED1��/(�[�h'e�{.PhD���t��˂������R����1g(8����-�������"�R4nk���sy�@zrsI�%��ץ�x����YM5����Ě��{�Cu�d���x���ڇ8jr�qVwΖ��UG����c�Enuql�7��W|��$K�iyڳ�q�;+�]��)�5�׬�zk#�sr:��Q�Y�3n�W�����ّ���)^�Y*��W��\ձ�d�7K�4�G�3���%�\��L�0����oD�������W�K� K *��&׶z�me�d�]l�����y��{�ûE���->�z������%�C,ƨ���H�5��Y�bz��9�P�&5h^�0*�:o�:��T:�$0�s7���ON}{����Q��!38�a���n���ţ!A�Y?x��Y������kouڽ�AkN�Q���9��*�vm�Qw�g+��%�7��ל�-����D�q� ���	�������047/2g��ÙFX�>���:ොcȞ74r�i��+��X9�+�G]�~�up�63�"~��ͧ��?A�+E#Ec^>�{mW��$"Dɤ�!�)�a��x��P�#�7,e$�Y�]��^[���Y=4�gVO�j��� �E�
G1P8��ʀ�r�/���q�u��2���-����4Ԥ���cO�Z0q�L��jj�>�k�e6�_���R��v�SLm��ڦ�k�T�n��gj��]���</%m�붡��@��s͜ܧ��1M��CMXpORi��}��嫺D"�\�u8��|A<1��^婃|�zm	�{ˈ�mq�Y�#M���>x��!1\�;�5��Q9u]L�%vU�!"�h��i+'4v\T�e����$O����Kx�I}���F���-��G����X��@܅z-��b�f�oX(b�l�y�[�U�=[5uŕ�VK��:�gzR�ҩu�WL
�n,�;F���v.�a��5-�4�w, �������䒥����#!L�5�6�nN�Nq���'����Or9\��@n&�E�/��w�^��rR�G&b9?n�v��m�0LX�G�^����Ņh�J⁈ڷ���!�DMw�]P���׻V�0�K4���#w@$A�b�o6\ai��� è�9�nk57a�EVj�V'\�4��(,�u:䓵��ةΙӻ��1s�v{9�xc��6�N�6&Vq�T�:�f�I�`��>֑����sZ���|�N�ۄE+��WV�F���dEA��\�;�1;kewVL�Ľ��G���>� x�����"&�P<j�1J�^E6�E�b`�w%)�Tɥ2w����%>��`e�R��T�v�w8ƨ�ri�Q��.H�Q�Ժ�XΘ�sQ=p�`d4���bksM"�sR�qW�S��$K][�A����a2���]��X�.L�+\cC.)o�Xrު�6�u���9�l"-!A�8�n�6Sy�$4x�r[���6"�Mh��.���Q��Is�ZW�A#���ˮ�ײє�)��Fw�ԗb��9L\u�#oh�Z��M��
��"��;���:嗣PIc��Y���x�]�ڗ�ʽS�b��Mv�Ǖ���!��Y�$[��Xq�w�^�u0���ۚ��:)�����9��#e�s�5+�o������'D�d�I1D��+�Ͷ]���v���|��o�I���bgA�+]��o���ݮaOU�"q�<��n�Ǹ����\d��Ǥ��m��`#�؝q#X!���
@��Q�#����j�=1�?Bz�
jV�͏>ʈ+OT�v���!��5�/��@Kz6�ý�2�}n�$�4"K����d;aV-�zN�1k9(N�
�Ѡ㹎��7��.7�X�	���[��f�y|c��j���a�Z���y�Ib��i�C�Ԕ�Mq��tB9�ߍ�ʣ-��p�&�Y}`kY��-m�XW=�3-�Z��3��8�F�6�B3�IN�U�����c��T���[�(S�24w!�Sk;�������.���c�̨`�X��LVԱA�M���k�p�̼���t�t+J�{Y#;yxjwt�$��ԈĂ��������J��üb�{i�=�-R}4{�x������c��h��z,�ں����N6qt<��%԰����\�g_i���[0���Փ2v�z�ZQrW�w=������'������]I�(�M��Ĥ:�U�W��S�n\l�Fn�ĥҷ�Y�4���i<��U��\"�]�vM�Ys!�5+��t��k#`��e�Ntĭ73f���e�VԶMpO:WgYs������!y�����J�L��t�9)�^�ը��T$�Bݽ��y��,���*�u=5dǜ۹X�������!�q�	zV�rfV_7Td}Zՙ{37��n����zE7.3��qF)뎇*�uV��L�ZVܪ�$[+�A�C�(B!Pe��2"�*I�[D���d�T$��!Dd�MJu�/��	�&�Ш�uL0�A7�`���	��d�b$SJ�(�����{��V��M��u�-�GF"�݃lU>Ƽ�(�lz��yݵ=ӈ�~&z��ꪯ���>y��?_o����g���6���`����n�k�:&��塨�ƘZ���֬d�S��q[lh{��������������?G����>�Z��}��lwu[c�O/<����b����u�og�u�M���9�;cF���k_������������������f~��Z��_���cl�k5�6�T�G�݃EE�ֶ���Z��)�:�m�CAT��:l`�U�A�W߻�υ�ԝ���b���.�ۢ(�Vn�Κ;n�Wm�s]}<�]6��뢲c��&�IHu���7|�]�kE[b"���آj�*$���-Q4MUM]���7w\I�ml�{N�Q�4W1h����V�cww�7������zɱh��:N�����wgX�:��F�w�U�EV��F�sF����Z��۵����i�E3Xڛv�5llo]�]���d��"|0!��Y��U,jqXa��4�\H��'ֻ�z[-��N���=�\ @�0�=u��6�T�'3%�@��rN�p"�H��6�Q��_��@��6�k�`����Q��[�j�����sѼ�K�z��r��*�˛*�_�KI�I�����Uv�,9��`2���=�h��*�ޛ1dNtN��b'sf�'TWr�
)	��v_E�j�rmgf����ɚ׌'��t��ǟ:g�Uϫq�����O�X�q�ڶ����r	��>�.�KCn��I˛��$6#s��{�x�F!��.��_���&PA�G{0���K���赖�sm��y3���`���`�Yò�ϟk�@e~�l2��2���^*���i���w7��,&�uT2��(Yg�A��r�V����������BW}�0�;;k�M�wox3d����[�b��C���Y�c��>��y��mG�F.�k9�;,fc�5��_l��HWu�Q���^VrI�*e!f��GC��Ui�!�V��S_��n��^G�2r��d����Տw���a�^�ƻ�Hl�]�]�4,�w�P��]�rQ���3Y��v:I���@�.�_by�C��ʷ*ӹbZ��r�c��-o)7CS��2��~ �KM�sJ{2���NuJ^ԡ��,���oL�4R��˜��&f,�x��w�k��tL�r�[�ʸwy$5�)�Տ��I�{�}\q�v��*����
ם�u%���t��3�6�ҋ'��6b��J�[{��gÕ�t�9W �-F��2EnlB��л$��.��6�Dl�H�9��Za����j����z��<y�ل��9�O���m��/ѭ��U?*��+�l_��	r�s���7�{��s�I�V�����}�����C�a���!�tW�F{#`RS"��J��&���]�cT<uA�St����hD�;��7�7�P������"�L����c�Ms��R-��Yy&W�=�c}��8m��G�T>��7*�=��Y?���6�t�߾K�^�%гG�hk��]�`T� d�0;s-��3O��tE-%����s+�ߎH:��e�Ok%���e�j�ƀj��,��&[TY�_��W)��[�HUW�� P-�d��\J���V��s�j�el���_�v����Ns���T̷���'ҊZŎ��W\�|�w������ךч���e���9Fww�3fC�8a�d0f�OZK�t���V���Ӭ�8~�03��t
��9^��gi�!ʓM��hPܩ����/.�CTu���Ů�^'���`ɡ#/{q��	P�u���q���}r��ۉM�>�C�S�]t.�� Yg�%�2�<�;L��F8X?L�Kؼh�:P����,Au�v��CZc���i{51�gRU��S�Y)�7u�z&x]��D�I뛡�Sb��E���l3�^|9��PK�9Ƚ�c-���F:�E����'l+^�V�𫺡gM�.��q�y�E�z[*�b3��] �-�pǞ��3a,�)q�J��fL�ןU���i��ol)u�}���.{f�� W&V�;^����W[�(�����48�k2r�cUgts=.�z� ��jxKv�p=6�Q-�Hޣ���׻��=�D��<�@�_�Y� y�Ź��!���eA�;�T���s�K�O�;���0>۟jW�{y�L	/��Q���]�V«�䯮a�N(=��][����`�-�;;�ٮ:�_}S�E����U�H�ߣ���vi�tK����̣��f=��������_H��N�KJF�wO�V�k*��B���d�]����@6�����1���d]�fg����t�c$V�}�|�U���[��}��7�DU_N���"
��qY^'���NgtC7i�u�~��=��� �t&�^����5Z�@W�M�1�k�hoi���=�=A�]��q��݂����Py�Ty��)�u��}ٿ���{���].E�Juˍ"�p$�X���>g����� �1{Rdfy�7��WiD񃧶1�SA�.�m�4 x;�ϔz��넃�֚�2�Nu3�i����B�x��� r�G���2_������m׷H��*�qn��,-�C�Ct�\�Df\��eD�ee��Kh�/e(�H�+k����V3o�>��7@�n���չ���'��p�EY��%tdDsl63{�ذ����7� e���3�yۼo������b���S:�Z�-2���!"��c���I��%Xv-3�e�V&yL��x&M�+��9���cu����3(\ۉ�Wڪ�f�n���Ӷ�X�) �T���14�p�4`&�L����[��t�i�ݦ`���ti�7j�e5�A�W@��ֲϪ��?,�m��,N����Bx��Y^K�\�}��#_���Kl����iz����^�g�m�cFf%.W����P�j�9-��F#�N�rE�#�����
ꕸ^�n��Փ��/z&��M��8,�U���~���L�M˺�J��Y��sɵet�k�,�
u���;٦`�s�8S$f�m�|��켞
N4�N)�`K�_˗'�:�D��睆Фɚh��p�s�$n��ΐz����٭��tWr��)���ٮ
[�3&�)6����bx����~����8��W��^��Lx����6�U�0�j�j�v�_�]�;@v��z� u��0)8�:.T�Hl�uݷ��u����.�V���ܼt-�,�]�v����n�z�z|۔7��=
8v����μ�1���9�v}΍�1g�9V)5�'��w}'K��w`�
��LrO�N���d�.��NTԛ��\\5��k�p��>Z0fu��>? M
�\BsOa�-�7��6�������z|ޥ�V��2VG:\獍��yx�w�ކ�>�)�I�:���dl6q�3*�Es�H�T��w��}�$@��A�����F�N�*R�YN�K�Hx����ؤ����*��0��E���i��]��K���#��Y/���I$���n�T��C�z���x�~>jV�s"njO�+3����(�T�e�0�FlG*z��KU�M�i��j�S�)�%R.��B�Uyjۜ�r������ѵ�p�Ϸ-��]!��1��+�z���Y�)��=�MU0���m#h�F�����dg|�(�*�X�[-�/��|��w����^KGxCONi��*�j��2tA��W�.���n��V��;.��Xq,B��KT^]�%��e�ky���u��c+6�[WVtJ|��|{j��j��jQ�x6L��t՛��W��E@��Q�r�_��=��7#X 7���-^�Ի˃;j�����{�v5���A�n��~��=�E�5Y��t�7'
v�E7�@D?.���޵fNс�t�X���HhZ5�wMA����8��_d�E�t3�e�5�U3�n-��$�]~Y��;�9}q�A$�{�$1.�&�͜���}=6�d]��zm�%Ev{���zg���clf��DIo�_
�@�l 7^����3=b�W�+��#�6v�K8�[��;�R���AƜ��6���؍�&�T:��q�fr���|8����͆4�n��!��6(�険E3NEޛ3�-�Y�0q���肵fsi��'��r�� �n�|�OmG5���a���Xp���"������͡��;��7UC�K��n�;d����j���6�M�Qzv�w6�$�0U6_vb�>m��X-4��am_���lZxD�Ά����vY�**�Uuл��<�/I�{�wB�f��d��f*�$I¦�|�i�s��T�ɐU;�Uty�r�(�&"��N6p;�^G`tH�9>&���qU{;��m�z�D�"�T��帆�S�\p�8�Ri��;��U�����nV��(dw��|¹VZ���r�VZ�Ozc4�m�\wMK�DR/��
�f���C1�Y������"7�=��x[�Z\��i�������6�U;�ڽ��n~����M=�/y]�|�i.��z!��߲�{=�/}��H�E�,)�5P{fa�#J��Mܖ�پT9�5ҼR�mUR���^f?x�ѿq|��, Fp�W&��@��˨��6�1wKtb�2�oÉ�.�z�u;Qn%r|�͖��� �F�T��؛�#��{`�
%���oQ�qh$&�܁�y��u�Ӎљ�|M��֜��`��i��u�#V�d�#�U���qJ��E���:��q�`��J��ͭ:��̖a!�t�aܣ8+s��j�ة$fp�"�2����X(¶���%�>%��{��{f�w�}�q���c��"9�V"��hC�,�ټjo4�{�P�D���{��5�ܒHz���(���턥B%�O|�/*��R�S�q<f�{t��2,��6l���#���Vf�/��o��o)���N��fk���y���J־�WR���ڷ�W�b�ƛ��������\�{2�y��ϣ���;|
�� w9'yBR@Q� -�@���gtU�RtS�_;�I&��\��������Ա�
�sHՏq����J���ٜ�q�Zj^��w��X���M��'�d��!�����gk��$�5X�=�v�n�K�,/ee�6���*��*c�${M�\����P�i4�i�S��[5�~����Ԟ�l����j��\3;����+ȡ�8��,W�S)�l,�m|k2�3s���D,���p��QKL�b�7,����mƳqN�WI<����:k+�u� "hr��.�oP2ºKĳ����.�D"�T��㖘h�r7�)��QlU_�P+��C�-���x�k�%�ڷ[t����'n�o[d�1�8f�?%�p	����='���f�3�=�٭�U;���%g�ZaY*�$5"��
�7�+V{�&��U&.X�A��F�߽Z��NU�٧�t��9}�ZL�=<(���Mؙ����p�:7�nm�8�9��9+�\	Y�9��U�L���ץuuz��h�n�'|��T;	h0Y�zoJ�y�j[P��RٹF��yzH%�ـe�Ա1^�\��:�ͳѴ'h�mN��.w(�l-飈۽B����I5�)k�\E�k$:.v�\ޮW���T(� 6���M���mAI%�e�P��^�V���A�7�����s��C�y�	|N�=1�J!���'\
�9`¶�E�]<S˳��]�ݧY��� Ï6�:�`�5(�k0|؍���Q�����{}���� �f]ωj��u�g���_�n*C{pg*�w��*�7uUC!���J�>ONGu��{0��P�D����Un�Y��Y�B5<���6��l�#�\��f��C(�8j�5>�k.�h�̷��]��jzׂ�g2=��1���_���VdYs;�,8�L7�9qeH���m��s�#i���UM�ģC+x,������0�ۼ�ѭ�M#x�L6V�"�Ul{9����(o�����s���2���8��z_�N��Z�V�e��S#-]5~�*]%R.��W��^�ˎ�k�Q���a��{��xÀ��/`\4/��Ar�\|�n�E�F�1b�t�纷?;q��m�	��Xp,���K�ؕˤ���w9�:��qT��2]�{	�#ܒ�M�&�/㶭�e�ֻ-����_I,�yׇ�7@��[������{���n6JVs��t�yF�C�@46,hs��>�%���Wp-�4]��vi�>Ѫk��{o>lf�8�.�:/c�3q-QV���yF����5��%B��U��謔����������a�(��}>�3i�����L5�cXr�s����{�[u�{p��k[����5��w��A�P�K�p3`M��&L��X���сWe�r;�)�U�L=���h�c�1\�T��5N��'"lˣ�M��bNR��U-�yb[�(�,��A��q?n4w��5�įBʔ�ob����9�8F�9��ۇ(�cBq���R��n�4��K`�����ә�7j%�z��s����prd�yTmY)�INv^�Ɓ"�Jk��]�VXo.��zW�;��L���;��.�����f�%�4��C(��V���[́��9^\�ƻ��'P���w;\�ijYb�q��,�
��gGXκ�7��oSB��Q���otK�٥����5�J͂j���.�Z��29s�h��Dp��t`W�����96��Qr��绉\N����Y��+[�P�������m�]����{���y*�7ٻ�V�*Jᡜ�\3Z+��*!R=.�<��������B����t���uy���N����^L�N�Z�_M��G��{ܬ�A�=Y&&;�[���I��Q_,�V��b̮#��5�Z�8��P��׳��Z���i�	(��`eN��L�
�s��]��ANa�s������3����}|*>x���V��%&�rr�(3(��<��h(Vg>f���Ōḇ����w�<ر�n��f�ɂ�#r�ʻ�%i�<ª	��JJL2���3�B�B�^��0�#HN���ٹo+ja�Ue���6�M_:ל��913J�3�E�]�Ǖͦ�dov����Q�`V~�<U�X��G���q���qA�6�Jέ{�D
K���\��I�+��rj�<�z��/K�+7���,��^pF�	
���X���tP�L�6f {�����b���0
���e7Y#l�^`�Ɗ��c	l�ߌLm��.�I<�]�M�~�)M�[4��[=o��ܱ h4l�O�	%���ٻ9��yw��쭈�v3`[���=\�X��-M���\U�)Q�qŊݻה���f��9wؠ��A2�$�0��7G�BO[��b���2�-:�=����U7{m�IoU�a2딸_�cq���,��ԕ��|�H$4�I$EF-�Q��Qأ7Z�'l�:H�h��9�����������?����>G�kgE�ۋ�n4�]4Ѻ�{���ݪ�+����T�y�DQ��||}�_���������s?���}4����c�E<U���̝)���sT��SqcG���|}9�|}?_O��������~�����:�6��F����<�U��ѡ4��[j�Z*;X������k��M�8��Ѯ��%�mEU-%�Am����jh�;mT=G]p��� +�]����u�C��U�ɭ������Ե�T���u�6zkl���i֪�v;�N�A����[P�jΓkV�c]��k���;:����`�Ji�ڣm�M.��Ti)#S��[mh�h�6�60h�Tm������S�Z(�j���'כ��v�&�u����׫v4m�Z�tn??Z�+}�S�=r+��4дl��2����;�Q@�\�rr�]������K�Y��Y�T]L�wW	EuG��2s��xc|'��>��O�6�{p�{T�To�V?z��%ݝ�Ł�ʥс\���X�ݫrxm�넆.�gJ�Y���n}Kl#����b[e��(���]}k��G7& �pU��,�s��yY�VB���t��G>_(g�ïx��m�KS�-s�Ղ�Ws_��k���(��܃��r�ӗm���iI��+�|�{��0ϡ�H�����iM:n��x{��,4�G�xge�S��rB�@�g��׌�\h�F����l3��lކ�n4�s���n5�K�@8|������p���v�|�RnQۯ���U��/��+Øn���V�؜y3���6�A�襔�uԿc��]�f��R��B+\�Jv1��i���i7A�ݢ�-��Vۛx��|֛�z@��B���k� ��U�~��WQI�qL[Kg=7��ە�������/Y0+ؽx�pW�:E��Հjm;�WG�:��jE���qv�g@ʹQw6e,�]I�{�ȉ�������xm��7u�M�+fĝ��u<H����7I�rE޴���
��ٴ`�2��)lW��	�7��D�,��}#q��("b6�6q;�����������Kj�:��ߢ��ǹ���X��7 [Om�m�ű��e���fGnX�9E�k%8��6&[~e�>{��'����x�׌�{0���Itށ�<���@����mU���I�����wV�'�,�j�m�ޖCi���E�Ĺ�����[f�WuOgV�:���O�k���f� �`(a~n��)n�#n;Y+��.W��]V�^Y;��Z�&���3q����r��k|ՌV��Ǽ�6�o[�-0���sf�[A�'o�������TNYQ�q�����Ɏ��� �-�K
�<�Z3���.sv��\���{8��P�sc81A��>d�ս�E�.n��]���cY�ܽܗ]J�Q݊w��c5����ȪW{-��8�f���J�gw:n��w��`�g�
�=���BӃ7凨On:z�xu�x�������p��V5pguA枊� ,բ7,�l��G@{ �(k��m��_a&�Lf���N��M�۝8D��M&F㢭Rށ�4���h^�w;�MR��t�N��^&Z�Y*�?&
BA��������~{��u�R�Z!�3���k�F�2(�(�wV����I�G�ȹ~�5dw�֨�����|����å1 =�a*��{�m1R+�=�� hB�Z��3�����K���^}i�Qc��^��M�RO[^���i"h��b�N�������@���l�VhWR����p���/O���>�%X�`��k-�`2.���U{I�%��V
��tD�l�����H��4�GChk�v�讱��r��=][����pɞ��vӹ�B(f��T����ag��:��-�g���oC���yΑjEPҁBy�+k��-��C��0�-�޾++j��0>���%�w>m�L�{��z�=���]ޕԝQ�^�5�s���Qc�L���Q���J�.[>x���j��\��ο�=�[��R�n�B����2p�m��m+����5��-g��{r\U��{�����,����������f�nL�:�]1�4���f]��%8�mhҺ�k�X8 �җor�.L9���.�$��p�[�åH�~��,ޝ�y�d]mRô2�ڐ��Ƚ�{Z�a��MK����)k�՜ke�Ъ���A�oP%�
�4���VJ��n��X��wjV�YW���M�F�IkW�]�θ��KA\}�+�Ic���}�Ԉѯ9tn�Bx�~1���0���\�I�x��J��g4甘�����+.ƺ�"u���r!ઘ���/^��;|�ܬ��<E.�W��Mff�n�g�
l,��-�9�1�L� ��=�g�4�wh�sr��7�<�d3iq�Sk�t� !��4	!�l��-���\�|8��3����6^�ݹG�W��K���b*$�U����1���lB��-��ׄ�%��}$ř�� �d9�ާyga��ށ��L����=�XU��G�t���G݊����g��hY� ��4���{
��׽��0�Ug�����T4�o�1��	Sy��ʎ�1跫��ăJ�`/?\��'���2�i�l�N��������E)gZ$�H�$!������6`�����]E�+���<iӫ��H�Y��˘ӫ�X��N=m��ޅ��WK}�������8E��y_O��w�+v��=7l�yB)y���*�fL[�DH��1O���;	��#1��R��w�&�h
�Qɾ�1��0�֖hHMn�N�w���#���l��wS���[�MF���	+���%�ɘ�vv�+�w����BY�k�rω���p�7D��O��H&/J(���踪��n
!D�F��E
�������}�s�ʬ�s*�X�Y���K\T�7���^woT a�!�����S�	e���x仂A.:�?�����ۭ�=� ��)��W��B� '�K��"�=p����"Z�]�UՕ���֘ q���ܸ���.�f�+�v�#w�}���f���+h��2���F��NC�O[&��d�gH�и���	o������C��Pr��a��l3����.�!Z@���̯�G�s~FyGv�ኝ�{��v��+q@�.зx�2X�WG;�q�O���3Ws��u�>[s4���$����U�=�x��T�`�µW)�w�������-V����Ί2����L�XSS�;�m�����o����	D{=�g{����1�E�G����d���>-m���|C�(��nJhgX#�r�;+;���RJ
T:Q�U����a��3ц���q�:&�hZ	���]V2����F_�����at\�"�b�m7�gv��^�L�1���Y=��U|��dt�<���ZwW�}|����m=�tm��w)h\kb}{�&s�>�9 9R�^�7�]	�����B�~u��ϋ�����q�۵����b��#4���Fȡs�X��LdrnR4ZkKbk���[aa7������Ȃ#���T�Ռ�������!��ݘ���J5��/��D��w���	&Tbۑ����M��Ê�[�Cf�W�t[)f��Zo6��J����N�j�YGh��Y���ͺ���q}^��|d>�Cg��fW�4���h�8��[�6��\qM��t��^��=wޥ���!R�"�^������O����ܮ��;��-b��:���p��A��9�[p$�@JQ/RQHv�3m]�4h9����2SmI]�=��V���д�^����S�!&.}���gr�^��Ԛ캾E��dҲ��aW�ͿM�?M�_`-�<˴Vt�ճ���c�[��m�uűy�2�
Z@�5�TƬ�*�E�$���l�7� ���T=?��,����D���H��ͭ���.�N�x�kJ��-���+�]�:�����?�U�N�V�_4>���� ��$��]�����X+�J�I7w{l�5�3�:�6Q�	�XB�=�w����}�r욥�$�)=���Fָ>��!����Y���kmwpq�ŝ0��"7dD7��;դ�ܛi�g#T�{���'��p��!�ť�0]��9�y)wf/U�vE�5&��do��uZ֙�Q[5u}�ݜl�~x&\fHc5��H�I���/�����S��C;K� ��������4���v�݁�B�ޘ��BjZ^��&^��p+�n�I�sN��'xP�i4�_���چ|�`��q��..���6���Վ���p�[m��$�j�Sx�zo>�ZH�y2�͐_�/�s����
�}f���j���pwaQ��/���ˮ"��2+;_5��j�8&�FmӤ�^�L�[z�[B�[_q�c�a�fuNN)g��R��9����UW�{t����Q�wV\U6ZJCX����qn�e�ïl^��DG�����	�&geJf�d��!?qY��r��e�y����/p����?U)�k3�R��L\��} 'U;�7%�ɞ�Mn&��y3��x�?{�c{��+�e��WݷIJ�~�%�,:�k(h@��Y{uW�{�z��7>�v�+Ǒxʤ6Aj�r[9¶Շ����I��Ђ*�}�n;:��_�]�\r�>οg� �tH&�|��S���N��R��v���4�8PE4�}$���o_��9�^���쀑�1͞]�'.'VSҖ~�[��­Ac��2E@�[���^@�訉�3��}j(���>�qW�J�V�
}��|�l��u�^l�>���w��iC�����=a(�v!���:�"#v��1�Ė�:lR|v]q�<��D|MW?g�kY��޺"{{��ނ�ʺ��zu(��l:KU{a���<���G]9@G�]��ܔs�:�X��bj�r��W	��fߏ*܉Ѭ���N~L}C��W���~]�΍�v���AS���+�,D^)5��˻f<8�v̬�(u�C�q5I<�ΐ�PWVx����^הH�f=xC��+)�A�qj�w�!� y�����9r����%�޳o������Y}��&�����4׻ـ0>��Lm�dE^dĦ��ڻ�{]?!GT ��-`ϯ06�O\��&P�;ߊ�Ѭ���T��������s��0�X;ڻ;cr�u��Q"|+�;�C<=n�Ƿ�U��^�U�F�Ŷ�A��V�L�{�-��^�߸���/z �g�&QC7���O����7F�bWV��&a�:Z����g�jT���n�Ul#���ĵ�Q)�˦Y��;H|�9�.D1�7m��l�;=O��{p�L�=I��嫸P���r���<׹>��:P9+����8���]�Q�~��|��i�4�]^Gav�\��v:�ږ�7'<o
���2����l�|��T[D����b��#?SON�3��.�gI`ɨ�e"s]x
�nsu��:q���h��
Uf��uZ�I\�iM9%CZ�xI~�Rz�"��A�7����(_!3A0��:/��
�wv
����:��Ѹ�*�ĕ���A��X2�ڤ!oP0���lP�q�Y�]D���	���';�B y���ɖc�>^^e�÷�Q�悲=�ܺ��f�t2�1�'�zw���K����9o��؂�`9M��
��W(:���<XlnIX���߱�F ���H���AF�dx�S���a	����PSA?��ee)�=�ؽӾ�����-
��f�`��&}zb (�ٚ�V��M��x��=6�ɽz;X�5yu��4e����(��Ds�����:�����0���f)���]��=�Vy�L�Mӗ�����띾�5���n��;�Cl�q��I%^���Ƨ5���3��.�t��~�Ⱥ�'����z���;_��_8�%b��R�j�G�ck���ؗ�sƭz
>�ƽ=�(/�}�����/�H���0c���� 9ƽvٖ^�t��\��$d�w
�M�ca�����հm�<�����~^kᜣ� U��@D~N�y�2�~ @��8�9��>�7��Q�$! 0�2�2)C(0��@�ʤ! 0�2)!"���C*�42�!"3¤� {��"�l����DLʁe���"��Q�!�B��{@!	D�|��(!  B�! �B!"�B(�� ��H���J ��J ��H����!(�B(!"�B�!(�B�!
 B�! �@��J���B ��@ �Hs
��@!$PBPXB!@�$B�HBD!	D�%��HB!	P���HBD!��IP���$B$!� R�A!@� �HB!�P�(B!	T�!D!	���Hhhea�H�!�`G����s�'8����+�(�"p ���A�S���~� ���?f�������=�>x���o����k������Q U�����*�(����� �������@�����D������_��3�w�	�P}?�=�?A5����=xɌg�ʨ�J$�	�H@$�$A �0�0�	��$$�H@�@B$
$�@J��H�$�
B!+
�$�J))(�0!+��@�))�
B�� @$B)+*��K(�$J@$�H���A ��@B� �(ă2�-�#H4�4�!J��?�I@Q��B�(D(RҨL�� �"@$@A"H��$�	!�A"
�����c��X�����'�����
P!� c��������ü1����iצ{�P]��!����;��ݺ�e��˃��M�[ܨ�*��Ԟ�S�d�
(��� �����~a� ����=� TW��'������c��!��A��	�;a�;��n��;��^_�Q U���g7`��OߧA�h@a?O`|C��
 ��`���DW���(n�v^��'`1��>܇�v�@�=I��^�]i�@�_X���~����� 
��Q���⪢������?��2����e5���ߐd�� ?�s2}p#�<�RAS��J*�R�)k%%��ld����6ք�%Zl�BJ[dBJT� �b�[4U
�*�%6�(�J�����M����4��͖�d���HE6*�L���ڬV�*�ZʱE�(�3![ki��mMh�ٷv�[f��	��EJ��FSZ����2#B6�-��J9(���K)(IUi�X�Ŕ*Q�
�ͅ���2��DU��[5��жJ�m�bԍ�Il��k*M*�Y��FV�6ա��̶�Vj��  'u���Wvn��m�ۍ�٣�ۭ6�yw��v���E���ᶭ�m�t^���i�����ܪ�v��k�Mv�;���W��i^�eT�������u]�(��H�H+^�P��6�IY�|  ���P�B�
Hy�O�ECB�
$H���D��v4(P����y���ݙ]j���:�z�M�5�O=�ӅӮ�[�m��n�k��v�Os���NwN��r�u5��z.�v�uW+�����Զ2i���{h;-Z��*�o� �^}kFk������ιmۭ��{^��
��nw\�k��]�4�s�[��v҆��j뽗/Nݹ����*�--8���[m������/t�]v��{��B�֮�緤mZhe��k�v�-i���/� ׾���Z^��J�ꪠ5ν\zV�UT�j� Ӧ�ڻѕUt�un�z��㷳CG�6��C��]OE�U+��֢x��F���*�m��M%ZUZ�  �=��	�gm���e���z�̭mr��w9��(����\ ;ۻ,�uW����:�݋%P��i���U� <���mmf�e6��i��l���  ��J�K�P��G��� �f;������yuz�Ue�4ׯW^��Um����z�l1���Gl�1ʪ��VY�bY�Ֆ��kl͍5��  � �}\N�=� �[N�C@��`��� �N4�tP�4�u��iB�iX@�׷�� v ��7��jdm�5[f�5�|  � �����h` M ���h Ǘ� ���  ���� (M���=�-U� ���p  -�-F��VRj��ڲ�ck|  ׀ ���� ��-<�@=�x�  ���  un tц� �e-� �� �D�X zQ�-l�,��l	l�2ү� ��>;�4 wO\ (�Ӏ  �:�: ��  ��ㆁC�ث(��������N ���. �S�	�T�A�� Oh�JJT� h �?S4�T�?ToT h�JR�  S����F#CJD��T� �j~�_��>?����;I�=����;�~�ׇ���"�j�#U�v{���?� �|>/�s�������UE?��x"+���� ����?����������A����A�x�џK���So�+!�B­�"�26��.�Ζ�pYaLn��k�cF�J�3�Hډඡ8,�B�8����)]G�m���`F����vo��l���f���.�M,Zh7���Ԑ�:-F(�nRt)0����Cbe;�9�Đ"�e�i��Ui�+I�)0帱
K@ʹ�6�*�@�cB��}3R�H�͖5+ddY�ɚi��n��P�3) ���#)�7Sc[Z@�Mbܻ�Z��2bؾc)+��A�C�4�!D܈8I��Gd�ne8�������*J�B�Ɏ��,c(�*�Yx�$�Y4�P2]�6�mm��']��e+�QJ �.����k�JS����9��	���˷�*U"Ɗ�:Х�
p��ը\�[$�,���W4	B����.��7+1R	��Dq�>ލ��
)��k�0t�o1��:V\V[���"Wb\��T��̄��B��di����f5��l���n�ѫ��Ѿ�wgMH?�0��X��ʌ�p�v�U�v���TD+r��J�L拙i�N�.5���#y�Ԭ�z�ڍ��,ؖ�ˆ�����VZX��T���+iՂ��z$(-v�f�l��U��x"�x�ܕb�ec�!��ƥ�J�����{��l�/2]a�TR���eI�Ѱj�:�m��\SKJ����6*$)����(���T�ȱڻj1x�o5%y�����)���Q�(6!MֶP����.�i��c�4��M)�z�Q��0�ޫ�DFT�oC-Vm��q7X5m�뢁J�2�Ac#�v�5�f��$��*nkL�QS��SŷZ�oi��4�a}�9qX��/m<�� �1��Ɩ��X�%2�V�=ٔ�?��1������WY>��.�Ggk$�V�K���d1wt����+YrQ6�^�Uuu�i��Z]�H���Cp�J��t�Z��;ך�MǮ��d��Y�K^�
����[1�k���n�����V�7L�B���k��Յ6�j��.Cn��^%�uҔ�M��
b�������.�K���ŭS�q��@�u��Ux�FT����%����H�Nཫ�K�E�-e��`Q����f�A{.,;�֤'.
�z���܎*����u�SL�M
eL���0㼗L0&3-L+T��bZ�
����Z����Sh�5�pj�L`��`�;3Aa��gIy�ut��ϦT��Y�1a�8C��@Ų�p��7l'��v�0K8H��� Э�i"M����A�V�駌R�^��pE�CP�e舅[��Q����9.�&�jk �M�([�*�����Q�l֚�T��U�A9Q7)E�Z�+11Vf��vui�r���Jk5�hD���	����M'�	�f�$dh��E@T���+P<�-��^0�b�ظ#cV�j�ֹb��yY�&Ձ��8��H$]�Km���[eDf�X�å��ƛg/�V�������
tf`�ۈ�-��g�N�ʗAAy��¬�qj� �GV¤�f���
����6��5a�؋�&1J�P
��WB7�!�H,��U �л�H�
V�P��F��͇JX
P6�e��U�QJ����j@:Lt�����Q3�n�`��å�n��%�դ-lV�����'H4��G��x$|��F��*u�����[U67Z@ەyc��%��
Öt��i�j�[@Lqe�
��kAf*n���� 4/iY�f�ًIu,1�`�)�����t�Y���2lu�JX��M�͘��Zk!�-�YN���8�P��׌k�Ȑ�#E��f�A-Cn]@�vAZ�$S'�Ec���[�j�U�V���K =Ǧ��H�l�`���Ş�A8w�r}�8A�T P����Q��J��Nm5(貚� !9@��WZ�17n]�d�,� �e�B�w{BE�B��tj�З#�cV�UX��0-�+wv�� ��,5yJ
��$���ڧE���+q�۱��YE��p03:�O,�M3�,ة����Gb.���ݖ+4vιY�	V!p�L:�.�,�w1^u���������G�v��e��/\kwL� �b�^������������W�]���Ս�U%��=�-wV������a�b�*njv�C�)�u���[���x �)�Qy�i���+Op�IU�)��C,L�m��"^8(���T��n��r
6E۴mڰ�Y�qr�Å�B����b����:n�M�wX�䉁���TGM#�f(���ʕ2����Xh0l����]m�&8���JL֭F�������U2�c*�M+)��k�+����"q�m�Цv<w�c�ȵp	��O��,7G(^�b�*^|�6\�C1�! %��^� �%1�*�L�D)���	�]�~V7lc��)-ܠw*��	� �y�N����U-	�����2avp|��w%-_��5�b���K���f��)�cF�m�H�`����-ڵV�o[�Fը3
�x�ܫ4�Ky�K;���g&=�1jU���n�k��sl',����ʚ�[�oBsckk�VP��� `:o�e����EVCb��2I�'
G���c[˵�!MP"��f��ĕ{�җ��R�%�ˬ� ��
(`��Ԉ�,��J��a�	{�����zj^}���'D��ê�ћWb��4�ʁQ(�2d4�T�V��H�G-�W/�˻Ôf�s"@��˶�ƽVq�ALͷ5VQf�7A��^�[�nѡ�X���M!���7�������o\7Pu�rI�իv�m8���XC^��7��,D�ƃ#HFH.8.zU7����	p����q%�-BBr%���tu(�yGv�!�)=�й6T���ŋ7f�h�%aӵ�*'6�Jr���8�E0j��V���,��i�����#��ѧ�q��#,��N�d1fPsA�N��ؕ��́ �hX[ó��H=�®�d�R��:p�\`�Ji*��M`:kLI��e�F9n�4v�H\I�C(7�h
r���5	5���;�8N���<Y������>�F\޸:{Q�D#h ɘ=V@�,�!��lݪ)Vᕹc[����X@M[���"m�t��'ѻTr0�;��Q$�Nj�t�8!Vu��2��T�&f���"���3v��A
�E��Me��Jfvf��������e���2X�6�U���`qPɦ�A�� ��"�3#ɰ�I�t��hhzi����t)���ֹ�$�H� �zp�P*U��T,`ҷ�76��p0�����U>G[_�[�Bu��
�%yZC�h�N��9M��%3�Ϳch���&�<w4�05F��L���+�PWM}�[�4
 �C,6�,827r�\ª�$BC9HѦչ�P�e�U<�RAVd
̀J*�5�� ��B+J���I�b�٭�[,�Dn�r�f5a�D1�s7j",衹%���PR��m\��
��N��7�41��̆�Ѷ!�Ak�;���3y�2pE ���t4�b�6���l�8�Xl6�8�C�X�u�qr���E\"؛�����d�⦕d�m+v�ʘ찛T��%{M��jI�5*�"����]fE| z6�2ɹg4A�Y�4L�0���7h��rTp7�Sq�<z-�q��q�ah���[�[hbQ�@�(�r�ȷl�����6Ƚ�R:.��xfK�L=���\�U)�gq�E���]�
f�U��  v�Sq溶Ec¥:�m�v�:�wI�Ѱ�-��KB�D�$!��.���B�RK$���X�mZ�
�&�'�R���QMT���\��DP�4Zp�b�����C6[�#Ԙ{�#m�KwAe�o'�l8�	+X�iT7G[�F�骚�6KAmu�����*y���Ӕ𽱸�,˙E;.��T��ce�ó[�/�eb�|8��x/�z�of�����HK��&�����"�ʤ�Z�]������v�|u--Y�M]@�����s��@u��iN��GSSR6M�,*�-39l{7`VD_-���Q0h�!�5��tF��0p��QL�ߧ/P��F\��5��%f�Щ����(�[y&l*އ��A���!��	�����F�\�x�ys&�m퇍�u,U��U��4� ��J�N�Ur3���F�.؋.%��-��Ĕȋ�0wUAJ��+q�M(��y@f�TH�q��jөD諶�i��haֲ������4�\[����`��#R8�CU�ѻD��Yuz滧�+�)��k�cB�u����,�]�5�.���jD-��߅�3r)�V�=ON�*`��H�D��Z���l�]F��O.Mu��R�lYa;1�ؙ��St֐�o7.^;�
CjcVY!C5��N����i�e	*J�V�qCM���+:�p7��6���&��S�ej`m)��8ݱ���4�`�����$�du�+~3�,��:�A�gvV0�$����X�C�����v���k�Sƪ�RgM�6�K*h��LeV��Z?�̥Y�+���,�e�bSt:L�,Jl�mR�Ѭ�-�����+ǵ1R@�J��Q�X�z��pP׋m��m� �&��Š��"=V�9VZ����Z�Vq��΁�1L��z�nRf-�/%J?'RV�N�KwB�$z	¯��;U�6��V�]ǀM��t�ɜ�A���hT�J�.�(3䣛��+ũ�^RKe�v�Q���[�o㯭-���n�T
���G��V!#I���X��V�"��\2�AQa{�n�q��"Ҧ�D��:���%$wB�}���::m���MԉFĎVgҞ�Ѵ�V
�r��+4�h�%nj�;�:EӨs-�� ���w��^�񠒘�(4TZ������F��-�O��j��C��WW���P\�;5�·���X�:6eViI����(�ބ��t^�w������5�S�pc��ŀ�X�ʝ,���Ḙp��Ż�Ս4��qV�+
E=D�X�ڋo7l	�N���0���� Êw9�nl^8V�� ����e�a��`8�A�R���i��ٱ|4M��Y6nn��Ȭ1�H��tU^���ǌ�Y���u�Y�.3v�v�)�6@�"�B�צ��Z�!�e!$��mY�-*ņr�Ty"�YV��s
їk0'kski%&1��Ʀ�B�����`ʻ�4�o�Sb�.���^/�!@�`��x���m�6`sr�Yq�e��<� ����˚�ϥ�4�ճwl��I��YrшE�(�)�6��ͦ�l���J�F�s�w�3_�T1����l�#+]��Pہ\�W�j=��^Bٗ�7&��fZd�FM�2�#cPLe�L54M�l`�2i�B�����%z���?c���`E�n��Y��Y2ROO[ R�֍f�	�iN�d��^�c��L����G,lia�L�RFҶl�$Z2���5�л�F�tS��r�����q<�o*_��zr�-������#V�5A@�V�l!����"&ޔR8���u�n���:GcMj%���elѷ(�ʼ!�h�M�+Ԯ,M����,��^j@t4�0��X�%TGj�qJ�ߋ�h�f
��E��j��/&n^�.�[FZ��+.�Ϡ�K%��!kI�De-����;n�X��N��~ѿ%>a�4�6�^��I�5���@u�a����ǡ���b�3,kU�JSlAZ�����&��f|(��4l��a�E	�7)ފ�Ԏ�:4P����&�CU'a��X ^}�����Y+#�m�cE!r�V껦���t�Sֲ�D�LUՌ��%.�ۆ�x1������dJ2	-�ϋEuz���[�Lb ���*Sj���z]��(^G�J�ʃ��&�J�
���5�kE+�'�f+� Q��qQ^r�۱�xQ��.�����h��°ɼ:��j-ajr���t��X\�D�/1��|G��k���S�������6Rͻy���	�/5"d|��##XM+o�f���1P�*G�鐶ء&��ۧ�����:Tll�m�iF��j�&��\ЪC�^Օ6ZB��i�5�CF�wl[ր���)��Sq�����V/�[�V৩��wX�ZY)]KU�a;O)�
��J�^̔ ��h4з�ޭu�Q�q�h�թ�,{�Ŀ�FS�e�0:��@Vi��cDhs��r���1��3����D>�!�-&��RFnhB\�2	 �	��#�E��R�N٢��Y���h��.�PPb��r�ֺv�	 w��
��\qis5)��n���8��7{[)���0ET��-6�]`"���*X�PF�������a֙U�A��H\F�

c�܆i�s+7vU�h��b�q�n����t��wV��F������H�hk��,33^���C6 ��PD�"�o0m^D��5ⶭ��HU�ٲ���d�+:��ݕ��L��F�Nm9);X.n���|��t�ޠ�<h�ܡ��]�v7T�.0�[M�Efe�!j��i�P��m�Π�T�V���M��r��{���T跭̔�= ���=}yt�T��Rk;R�e��@^ei�8��w��!dNV�Чi71��R�&:�o V��n�;��	g"��=�LX)�F�t��Kʶ������*��%i6���q݇b�ܻ��fi�m4UJ��*��u)�؋0��[��Y��ș�0;t�-R����[U�
�I!-���C�a�v�\8ڷZ�7��=�4��+�a��nƶ�������aI�h=��o_�}`_=[�c�+��_b�U/u�5�u����z��)�e�<P��H��+����ӛ4t�gUṺ����Jt��M�Ԁ�[���sǝ�ຘsb�;db�gQ���ƉB�׺�cn�9�e��~��,p��7Y˔<�Y�}k�)��VՈF�x �mP�x�7�;Mӈ�Z�3�&�l�LsR�f9�S�/u��y���w7��i&�-��\�*���;��m���.�\(�i�	���l�����G��(�P P,a*3�@kc.�Ԋ"��x_+[X{�
�Z��ܮ�X ��ndn��P��Y/0Ձt�q�e������l��{�ÛyHO��(��u�����*=��#� �]�Kn�6�ө��5Q�w�u��p<�o�"��E�>���l���nnF�5b%���ڜ����e
�A]��[��*�tW�a��dH�ȫv��u�
ȼk�I�'��"�6���	��3��Z��hfغ�Y��fBr��]��F�w�ߎm�)ԕ����aj嵢�_w5�
}�;b/�����Ex�A�k��3�7W��,�z��١�3u�Sii�:����E��֏m.��٣t��4�����x��ޒ��Z�pP%]rK*	V.(�x<���^oUц<Uk3����	��G{��&�4o<��	�\�M�wD�xY�n�x��S��	k|�X�Ux*���F�Ĺ�=�V����"9i�k�f������؂��ӑ�����hy��U���f	M *4�J�w.�<YZ,�_ZCn
����̷��4j>�'<2�4�R�����-�����k$�ꏈY"׫�ɑͳݏsc��8<���@(v#��H�������ǆ�����hb>��n)5)�^f�9&n+�,�w+�֜�����д��c��j��\3�</X`�%�4�����^\�$ce�9x�$N�fc�8�}Iـ�;`���EϗY��;+i�	|�2�5����-*��z`:�׹N��vgo1k�������n�D73/�i�pͅ������ÃC՟w�ٺ�z���f�u�],����gn	{����-���0ʗj��	v��f6���!�r-^u����h'���Zl����G}�̵R�(+J�z�ea�6���e:�0C��W��gܰA"��cQW{�ݺuF��<������Y2��[���E��:.�֩�;X=m�\0���욼w8�M�ӡQ�����b�}ȉ���Sǵ;	,x�u�mS��h��te��ـh����g�^u~Q�+�	�Iʺ4Ty��y�����Y<���*Se��=��<=ܕ;D��,H���c<���٨��`*���Re��85:���+Yb\�3N��L�;ʲ��߽^ڻ5Ҷ4�}+4&�
����2��S��*XU�-���ʾƪcA1vEh����+��J���m��JM^V*���1b-��Ԡ���ߝ`ӷQWG'}>�� {�$;�1s�b)c/;���M��
C1��&=��O6_^���h�0�Ef�S�����U(%���"�&.^(�\�ی����\���kfn$�i�ĉ��m��p]�4�������+`x���-aU�$ì�`ɷ�G�T��f�=R�=�7�ӽ�S޶fxQ�(�A��eP�l,�'u�{�.����|�e.��1���H:V�ʮ(񿔄�2�R�(	 ���PU���׬�cZ��������9�����|3��7�ď�t�e�Mz�C޳A���q�(b$y�{{n͠�~̶�ݗ�{{ׯexb��.T�u�ں�{���ͨc<)6@�w:�%�.P8�fe�E-Z�7�\��{wm��1<=�K�O�Yc�H�B�˞Z|��DT6'G��	�)�,�{�
;}y�y�j��	g<�l�n�^���!��Đ�C�K#��D�p��#o��y����'c?ڼR�o�Bmx��4���N
Σ,�xl�u��<��dnfdE|5�׎��8��(Q�>�g���3�����=�W�VE�^D���.���Ǯ�!� ���̊wP����:w�*�j2���X6�3'4��-	�òJ�j�^���/@�2�m{�硹��JI���Ion�/�(�/����+3Od�=��gf��q�ۘ���-L��\O�x����n�l�T�;��G��>�U�M1��9d��x�W�Jy��y	g�%�f�7y»ݝ��}�D	^�u����WC�ZEr��r6;��k��2i�@Vj!�%���)����KzƬ*���	^���B�t'o��i�W���*QSG�3��G!ڪ���{r�H⡏��#��t�)H3꽻:V�T�e$ի�V���S�7V_J���HeZI|b��=��rگ���rB�dB`�[��Y��u��YtD�)ёm��UoI�=�5ٸ����;�aԡNm#���b��6Z���b�|��ݴ��h�7��(�z�h#±���j���r�{c{��I�fQY1n�ig*�ps!�T��'�y�z�kp�߰�%ր������qH�����yX��(�ת��xm0���I��y�U��m��C��oXV��	���5E�	�:{{�^h�H&a�\�Ge�bOy�W#G�*��>�U�J1�E�E�|����e16sJ�!����Vr��/�B�-P��v	�2G���2����N�� ��\��Z��T`wNJ/�]�Xt<�Aw��5�}����18��Ɨ9�;3Һ�ђ���Y�[p�X8��������WeSg��LE�f�#ZEȞޘ8���ZAnu��e��Z�C��ua�[eR!�a����Ō��r�e�Y)��iu��[;��g 0�\����V:5:{������;ݰ�4�V]]�V+��9����2]�Z�bl-j�����uN��$y���փ�����qI3���Xm5�2�|�y0=�dXm��v_F�v���f�cO��a���;Gwg�~����lZ?X{�^�n�^���&C�j@s۽O�4�E�	|��Jam	�����Yb�kE�4t�ć1�b�۳D����"�	��6�5�fNbT:��O6�]�"&V�껇����z�-��p�Z��o�|�J�ʰ�c'Ƥ{��Z��B��-��N	���p�N�3��K�YrU%c�����K����a��y]���0Po�W�H��/����/!�f��l�� =�pT��J؃��KsP��5�u�t�Ɇ���t@k�M)���������t{r�Z6�>9�b���E����Ϩ����He��������FE�3�:�Gz�E詏5��q㦥t�(f�eYT�յ��"W]�N����.j�N�3E]pmk�9;�XK�Y� ���-$-�꾖-L���F��R�ӌ
��j�L]��$Uϝt7wR���[�X��:n-0nmuԢ�N%�z�����Ln��r�����)��i�O,��q`��ϝ�>�%c�+��ȉ��	t5Ү7;F��:���������bO��dH�eC�r�Ӣ�a�`^驻�L�:�����o��qJ�Z�P0��έ&�o}�ed"v�����fɝ.8��};VL@9��)f�,����,�vQ�)e��@���M7��m��D���ܭv��aG��j/fw�:_[�v��w9�>�(j��&���S���طe�9ty��pɛ��s�ڡ�Lv�K��D��@��� ]�\�X��7���D:�\ޘ��i�-/��g�k��%[Ji�e��7,k������ĵ�������r�񽴼��{c��x�
�2m|-�}pEm���,��r��h��9��#��J8��:�XU=��(���{t�l�Wo=�ˬȧ$\�����I�k(X��j5��#�u�/��X^?,�{:s�(�����oZ�{���t�p^j��GBrgxm�@59:��
&T�4p�=�J�3�w�!��MM���`�qau���R�*�%s@(�X�-J�!A٢�M�O�#m�P�We��^����ه��j.�f�{Ҡ��ߖRWw>��3�>���:�!rL�f����M]>�� L�X���'��7�K�]�}�R��@o
α�Eצ���Fk���;L�6���P��R0�ؑ�q�[s3Bv�uD�x�l��wv$/��S�e!��r�Z(�I;���aS�l�M�'���]|����=�7z6���-X���戞jC2Գ��%i5�9ei�˶9�Y�1խ�I��3�u�B/j}��)Q�`���@�7��F��y�<%s�v�e��傁��kwB]т�����3j�sC7���oi�[�I�c�ʭ6Ɨ��`|�.�Ĺff��<E�4�u!`h�4{H�ʋ�寸���mh�w�Cs�{��m�99H�YWu��e 1`GEǋPIL��^%;�Zr��8�.y|�N k��	;��}��Y�C!�8s$yؚ62�}�N�Y��dK.K(:�iAV
�ya�� �
�̗!,,X���K�f�!z���C��5��K5�O.O)؋b���v�o�J,�,v�@��v-�=�PSY<7t�8���bT=��w���u�������n���M�E=�yDҺL���I%�FW@�*�����w`X��8N��|��,4���sY�ds�>iY�Ş�[�����c*ݽ��(�om�u �9�f�[43nc�7�s��{{w|���V_;¨e�_D�i:f��wQ.��JV������}�1�is4G%���[��k�t'%�B�T�V�Od�KƺM�� ������'�ُy�2D�5ӻ����|nq�b�G9�M3G-Z�y�n�줚�Ov���q��"wIn�م>�
X���
�Y;���2�f�kx�f��+����f#�-\4Q�y=�M�&�.�"::�|�V�p��yXn�l.�)�ٛr��g�,��S�&x�͢�C0� wf)f����{�5d-�mom��89()��;�\P���}֙��0��{����lU�u/P�� Z�Lq;��m���VGKݬ�M[�掹��.�vt���bYl�]�;gIy^v�\�����c���3�	�NQp�cN�
��=3�N��~/7�zH��ڭ��fm^��"ǫp=�#�/8n�ၼ�4�ʱH��Xۙ�N�������(r���q�,8�"��8dX��FWA����u�͞/O�4>��0a�k6[����lv�������X�2��3z��+�B�BJÐ��+���3�"٭��V��n�� L�NM+iw^�c�է��_�S�e�*��;×]��ԖVf��zմ9`T&��ܷ^���|��v���*��sc�8�wv;�ڵ�c�3m��r�3�Z�-Y۽=m���sU�4�̥�ܼjty��޸���a���M�"���ٓ��=�Á�L��9�uR��$���4��v1����Ԏ�vȸ�֗e�g�V�Q�G ���aH������s܋fOXݝ}����g�&|�w(
K��í��c��كZ]fTE��W��˘��]�T�����ziA>�yk��k�����b(t&��ë|]�Z�\�X2c;9)/.U�6��Jgx���$(�Fe����]��	�d�y���am[&\ȰMɋ���:ViD��I��wyg���ZD�w��
��]�?�z�M�����`q�λJ��x�ǀ�4_<�;x\1\^`���[�
F�=y���j;�a8�d�A�d-*�^<��	��J�u��-/����i���B���{���Y���Y�A^T�o,7,]эb @���A����Ϯ�Lz������t�Ǘ�Hm���הV�5�E���et�鋻���.o��-͏[��:�3�ô�����iP	�Ԙ��>�VQ����V��Q=�7�
��K��];�!��֮���b[��Ǻ��h!�2,O�o��՘�X��ǳ �-���ۭ���'Vފa��r_ĺ�7(,��-���ww�Ǳ���������^�b�}3��@�=��Zw�Np�C�}�;���\F����0)��5W�ѯI�hj�:�Z��*$Ŵk��1�;Ԗw*x�qx������ʉ��ܭ���Ԍfw�u5r8~�n;K-r{3Ȇ>�۱y|k�L^!�bc4�̒c��H�����<�x�r�ꆶ�#/c���@�:xF��a�Ae�Ch֬]�J�`�̼ ޔ2�-�g[��(����c@�'�	$�5m���e���j��F:����8A����O���}a�;;BF��g5�3�"M��C��,�b!Ԏ���×:Ү�u�3C8��\É�Q��M�oj���OY��J�N�����p�\���f]�Ȫ2�΀,t��Qᬎ`����L��4�u�6h(s��7gv[��Dߕ�M�TY��}����\�H��)�]���}(X������Z��Rt��1k3%��Æ���î2�ei�;�7��o7�J��GV.�\�Q�&P���d*��1�³B�q]bx�m �
�wZ�2����-�i����e�iמ�E�Y3pw�^c����<������"Ϧ_s�.�n��-��?�����j+���gqщ�/n�|��	�φ.X�Y�T�)Mp�`�t��f���<]��&8H�b��ԟV���D��/�^��C��#���?`���.���\g��A}�<"�s���{�W�0ɇu�Q��[8�0Z ����3ɸ���;Z��ް� (Y�h�
����Zy��y6��3H ��1fLՈ��E�y!���DǼ�{B�s��~c����Wϟ��������� DG���A��g��O�JIj�lu0TR\�Aa� d����6I���{��Q=�!��e8Y��S��Rp�����}�0xp^��"�g=񀼤wgJE�`ܫ}s��7�Iu�۶C��Q��]GV^�z��4��9Y�T���"�D�/0�չȭ����ᔮ[w2��j���zS0&s�ϜG���mXI���TB�4i�]mՐ2���Ŝ(T����Xn,=|8Z��_wpgf2z�W/a([�E���B3.�oڝ��g!���W����j TbW*P��Z�PX�J���&To11t4��ֶc3U�Rs{@4�]s\b�6as
.�����\˻/	�D�6=�9�#�Y��3-e�x�.c�w]
�éA3�ў��;��25�م�uy,ήq��`No`oN�e&q���yd��z�l)A��bF�Z �C#nb�n���������{�� x%���W]��j�b����W�������S+A�}�����{��Hu�JP!6�l�cc�p\�y��Z���������oU���/$	��΅-�k�A`3�5f�Y�no�*�]�Z�h����|�E�NW�+	�
��KtpJ�u��4�ʇ���3�{&h�煁sD��[wLX����r�,��٧�EI}'�"}��bP�P�{�����F�t����Z;q�/We{�a��^���݆w�V���7ORw��=Wi��7��jV֬,  ���C��UL��C3��4�����I>���٩R��1�J�w�fU:V9!j�㗧w+n�k/f���e�W��oc Y5�;&6>�%ڨ�̠NM<(J�Ʊ9��gh m0vg-��
�Z����;/�i��E�A���s�K|۷H��Q��6�o-u!I�=�[���|4
�on�	���9����R�.��6m�����m��J��|��]�dm\xج86�@��jj��+P:�s��ն\
Y,�D]�t��ʾ��j*Jɹ��=�r3�<Qk��#�Y��Q��V>�v�:yZ*�"o7�ܨ��e>U��)*7tP��t��F?��V��1�)d��n���j��(����X�.��DMO�:yz�'4����Ɛut*cF��k��lk�lE��\ʊvf��F�E�8��(nn�u��T�]!�q�w�ܭw�B�o09GF���Q���K<���/ZK�X'ef�Z�?sa�[.�d# �x���<�m-:(nQ�OW���z���`lI�uQjN�`����Z�f�A���z�.�,�]�l�ͼ����.��dC$�Z;��{�M������"';%�yDĒ���f��{�_V�|�%On�k/N����iýE�FU��:�Ɂ�G+(3��d�Qw`f�f��'T�\�r�{�E��L	���}ʖm��Zg;��e]5�6�8��Һ�H�T*̲a
e朽m��L�ÞGU8������K��3��B�k�(Ҭ�V(��B;�,r���h�W{��w�gXzZ�GM�q�|�$�IY\�.!����K���4�C�j=,>�6��u*�q�W��p,W�P��o�*�C��� E﵇҇�6~��Ø
yi��3ٶ�t{�Dr�+���l�6'(+D�c�樬�K7,5�:�������	c{��ܯ=��b��yM�Q�P��f-��j���'�B�Xf�c�׷b�a���K��wƘ�m�f`��S�
���ͩ'��!�tiaY,` G}�0*��0m4�����������W�;�1p�^ٲ�#�i:O�QR�����p�2�8P@^m^]��7o6�hU�b�{�y���q�}է�t���*�R�Qkw�2���L�4�"�M<�I
�F��U�iJ����'N.�3��_uI��KN�qTl��o΅=u�=��� �]�}�_]�)����!�\S��]��OP�r����b�V���^�҃�j˜��t`Yw ����/]sR�XV��
�G��sPL:`�nwZ�Pb]}u�vP�Ւi���x�"���4y��q4]�Uc*�32*�� �X�j�7����+(`��q�˴�O���Iq�x�z��Bk݉�l*<�\�V�0ʽ;O"��..�X7����WV�.��2��������o:���#[���{V
�i�*���:Seu�/^	3N,���ͮ80-�t��=���ς�*p�}���M©����P�e.�\7t�����}R���a�a-�TUY���Ka伢'-��S��X�/+@P.6z��2�|�޶��t���4�P:fk�OOwN�y̐N�W�v^�����#���m��j��N��9Jt�e��q��e�����tg�a�e�:d��/����'�S�J��W�պ:pݥ�����~C^�u0�s/��^bq���p>o9������4�ge��^�B�
���q��Թ�s�ݡ�u�5S7!��U�ot/��	3v_&Q��;wvt�
��(1��[�;��	�V�.�Ah����Ev���4j��#������8R{8v�z�-tǖd;�~͜H�X
�������ŋ��r���(�����w7}R����w�;�����͘��"~�PX�0���g7��N�3"�x8������d�P��<;Ω`+�p|���ev_�X�
S7Wm�a/�^ڶ�튷����]�BZ:x��c��hb}�l�����j\�!���ӽ⊅W���"���Aм�79�ͤ�vq�~oM�E-'�ii*>Ò�px5|��v,B��].](��v�)�u�Y�m��Є��1N��`�[64��˨�.��7��(��iԧ�f��5#�
�e��бzb���B��w;gˋz����2�iS�b�N��Hfplo�6W�Wy�[���e/B�A�$���̤���_{d�
ɀ�w�4�Q��N��Ve-�=�e��:&T���|�b�)>ұ�Al�c�VY��n�Г�3��XZD�/�LI6��`WU�m�R
����e��59d�WS��Q�,L�maK�dV`��9�zF/�_J�@2_a�.�sP;K��k���^�����q�c��U�(Fi6�:�G����
�!G������er�V��eh�s+�䛬Mb�a#�� wh�ۣs9��Dtт�謝��5I��d���]��e@5Q�4	�ᓛN��V�uC;8+���L5����`\�k�x],U��-�(������X[e����s"�@�T�i��"����ɡ�Ϣ�vh5[�����k�P \\́��̀[�s�r�(��%*9[r[�+��`�94��T�Y�0��'�Hբ)R�kqpv^0�*cV7{h����b=a]�U��w���p�q�/Iۗ5�S�WmY��X�E̸lH�g:��(-Ku�XF `���̣+�����{�?��C�]�v���p�c;��7����d��:���xh�sATz��b�����!��5ȩǇQ�ĭ�lc=a�u,���b�n��N���]�u9�Ď�θ4��s/I.2�\�M�<�j���s.^P�.]^�����s��.�����tca��|�_̫�s�q��է;KM|�|q�����R����F�6��4
�Y]�O��"
�%#�ͦ�}���d\��!�O0? ������ym0�>$^:X���쬮ozvҖ`\����	{]�9]q�o�����,�n?��_s������y��uǝ�n"�Mb6V�7���;9��Ƒ�j�5���*��Ww�+�]��^M�g�3D�S�̭�w ��.�J�<�s����ip�6����L�uwZs�%�5��X� g.um�������ki�]�h�{o-���u7W�=Z�l��(ḉq���U��\�B7���R�jG�m�������P[.�е�}�r���t���4f��䃶ۡ�z�N��X�4�TjZn�ꇲF;7$��,�
,��գ\��6�gE��W�.	wm��^����A3H���gV��k��`���Dwe�dX�K�nW8�ὢ��gd|j<g�r�w���\`�wE��aK���ˬQ/Z��戽O���U�'��UZ]����mŸ�[�LEN4�����*������TvKƍ4��m즸m,�@��1J.��[�rm��U�v��ObD�H��M9@aIg.�#U �'��l:������3x*͔ATQ��Uaۥ1�rQ�r�9�R��f=W���{����)��r�؍��<��6�q'�7p6V�_�`�9���||ofW�}(��[�[���w����M�3�0�����]��Zy��:5��F����sz1��f��'ҍڳ�@y�pug��cG�z_��bBޣ������=�����%�9c��F����u�4���s��Fg����}�bDz���Z7H�yv9�%[�"5�߷���a���s̰���C�;$��Mľr��dd
y��H�Dٗžu�%���#��%�����+�X!$0��8�3�����V/5��; (r��g�#��{�����X�%Bh��Ӱu0u����L���)׀�I�2���0n�z�+�C2/�~= �>�)���~`L��xH�(�9�/�Eѳ������a���B1����<���}��,����ҫ�k���=�x��k2�y!M�ֆyǔ
�_4�ĳ�*5�Υ�c�4��/u�a��<]�'�Kf�K"7������rP�vԬ^�5�2,Ժ����i3w��%5j�d^��ܵF�h������S�$B_j+�sK�4��@i�)�t����Mj�&(��=˦EnЗ,6��mY����m��F���X��&�۸+N��+j؋���{��S{��lwӝ�#�<�E^�S��w:&�s1�qQ��x��`^}fh�;�I&$6nj��E����2Q�Ke�Ul#5��Li�Et��PZ�޺�+u˒�q9��~�=H���;"�j��&�Ot���{���jI�egV��E�v��.r[������.*.�i��b�سx�;`��c�Q�i]r�߯�p8�Xi�d�+�8,�Ʈ��W�w=B
=^�9���evy�E�o,�.��|���i7*�g��J���ͳ:�H��o��V����:p#�-��$�6	ޚ��tFuʁ��z0Y�X*	zS���cY�Q�`��Rs�cT�{�Z�8펍����%�Z���L�]�>v�\�1$��J��&j�A�7ǊG�g�d{뺞��5]�͝5���c�W�9��+��&��4�]w��3�.���Fl�Dx&�#֮���$�]W0�Z1;��-b�h5�;���{Ύ�Xc`���8�H�̌���<<�59�g#CHC4VFy��b<ȓh���F�0a��P'��\;m31w(���8("K���=`�I�����k2#s��`�ͿPsےwvﻵ�^�"~��Y)�S�k��R�xdO�\c�]H��TZ� n����~d�P��[��Ǐ��:	�x��S�w,R��ҫ���IgA���+��P.pOl��/��W׭�`�AR,��B�[9�.�wea* �%��w1b�ҫ��W�%gYQ'B�
���W�wi��n;<7ͧ��z������3;|='����ot���Lt*��F�^����c��8o�^H�o8��`��ڛY5jI�n%��5�V ��e*v�]`15R��c�C9�=Ω.�v�1Z&>��
��²t��nFc���21�Q���^'��Y�j��8��V�l[�$5���L
M
�]�;m̝m��Ŭ�N��f�UXo�ͦ�-7�X[Xmai��\�y�<0�^{ȟp��ů�nj�Q<������p�6ů�k�������:ܿ�î�SkFX���cr�gur�z��-��XŚ�����Ԗ` ȯR��.���;RȽ��m8��'���I��7{^3�ǹ��|1sF��a;#|��jt�=�)�"��d�O���ze���:h�|���<��Q��9��L�Y�o7c�\�q�S�hS�W'�T�^��t/oc/��a���$Dג�n��S)֖,�5|*�e�c
�gs����p\�mbM�$H.�����vn������;XB�9��� �ymeȌEZ.���(k��ȟZ�*�-\��o}ς\��57��mG��1�gWgj;3�ppZʄ_Yb��m ��m/��V�Y��#�dly0D��O�Z7=.��wm�����+�G�e�]Hc}��x��7hF����s���ĩ �ڱ�l� {w�c�����x���"Ʀ@vj�G�&�v�{�C��&�(����x�.���4p����ٍ���ɰ
�;:P�����x�5�g	|�ی)���h�\�"��!{{��w��ю��m	a�n��$ }{��6F́^\�,a�T��O���f�8�E���&n��^��=���,���,cW�%��H���i��,s�b(-�]�a 2^!Xi9�� ���f�9)��\����t�Lh���o�Om�Q���W����;��-]d�U��#�x%�B�<�3�r�g�����F�ɔ�sX%\�3��o��V��:�t�u}w��,��wӌ�C*��i=� J*�RO�Nh�W��sC��\Q��w�LedSDi��YGE$��ʭ ����'��Y��x�zP �`XU٭��ưW-·m����{����L��X���t�;��JF���A��Z7;]��o�w��M(���1r�X����Ct݃� �����>�!ɇ娲P��=�{�l�9��.˅�-	´��'��c��:x���a*v<���XS�y�˛���h0���G!d������w����ܧ6���7���Ԭ0��n�+�
k�a]I�i�\YÔ����Dz�Y��衂�}$�d�)n	���� ��n��h��d��vc]I�m����xF����nrۈ����V++c�����z�/Qm�;���K��JP��6����3�B���3h-/WTcl�d߻���̛�=�s�j�C����+�n��Cn�%]sQ�/�r�t6ú�$,ev���c[�@|K�{N�Y8\(����ㄭP�:���`���Y�MB�t�)�d��47O9�R��q�;�!ՁnGKr��hH��	���);Ə{������ϖ����+{g["�FŎ�<E+��r�Db̻/�5�_��g���AT�aNxR3iE��/
�h;V��c���tX�X�d-�q]P�]����l�W6���i�uLtR��ۗ�i�cT�0V�ͪ�v���Q���mq�[<��G��o)-o/�,ݍ�^,w��6�1}�N<��O�3E���\.YA�8O3�$�n�v���a��v��x��m�t�_2|1o��D�)\���F6eW*�v�3�͇�jѬ�s��ut� |�?aM����htQ�\�!EDp�����;e�B�F�Ԏ�uMj�Zt%i�Ӣ�
i4i]Zֶ�%+N�C@sj�h�J�PP�<�Iɢ���"���䦞C�4��� 5���l�Ї'���[�A�䍵A��hM&��QAAIBV6Z4	�j�F��<�֐�<��Ֆ��DIl�B���liu�`h8C�ѥA���K�5�a��)���4Q
\�5TRii�7,%�4�\�5�F��H�h���;�4�Lr+$l�P⦪ah4r� ]���6�[�)���I�5G#A���`W!�'+`đPR���PQIX���A�O6�lPsQ�.`t�#���.���!I�U�.��l`h�$sh9�1}�3X����u0>
���*xy'A���1��嗘'13�5[���"s���N]����W1ѧ{/��N�ד�,*Q;�g�+�Xh���G����*˭{�V}ָ0w���(4��ѝ@�f']��)Y�G8��u�� ��6�������>���0O�@�����$�qy�@�G��#�'K�%@4rU`�G ]9*�������[���_�Z�,�ҟO�yO;�ז��U,���hJ��5
�Qiދw&��k0B�rZ00��1�S%��}�5�����s��b�U�\
��b(�C��`�F��\W'�]5>� ��~�l��-�:�-��׺���Lz���aY_ +αp�|b,�}�#�vag�_�/��VtwF�|i��,:ґ�F��]Q��W�7��<�C���hxT�@ei�<q�s�A�:gc^CS�;2N��J6�o��pk=�ؘ�u��\O�DR�߈p4PAZ�����3��h��53�y��*�zF���81�jL�r�
'q�T�J�V��5���� �+���v�k.z�� j{;ø?���pzjv�<s��0�����ז*�����ǰǍh�MA�dB�Ε�X���>�掜�Vy��Gh�t�&�#�N(��Č�f@�K��Tz��n�֮:�̠�H��#tyZ.p�,b��@k��a(s��;}���Z�:��%���(�������5*#�������P��ʗn�].���ٞ�����~�Fv3�a����\���Gc��]K�u��N�i�:��j��dY�<3 ̋���&���@�u��k=������#87�C�����֏9�i]����s(Bک�);[:&A����
8#��Ңa�0��NyW��pдp��8�U���8���_
]S図6��=�
���"��{�,Wa�4�f��W��6Oj�^�􄷇�\�)� "��ʐ�
H�ޡ��EZ��Ƃ_X�ª��V�bmG;=��e�������Շ��K����6�M�o*`�J��#p�撅0*�["ov&�3t9F|v����aT%L�������*������}��*�9R٬;\�kI�{6s����m!���E��dҳ���< �<��j�1�g�z2�P�	�(�[�)��񮛾r��)��)�R�m�n�x6��κ&�u���8�V�����n�*��F�VZ��.�u�MJ�^c�T����yKz̿k��-U�V{��| UDo����^��'�l��x�r��=₻�C�߲�
�Q�f{K��Jk�)��A�s�l u�o{�q/]����s^3�R�>|�������V��!��}�lfZ�Y�r_����T��ޭz�u�O�9�C�IL<m>�yP42R��h��KuM*g��9`r��M��58w�[���`��R� e�����~ͮ塊4=�e �YuKY�~Y�8X�^�Vo%�瓫kK�⽔���@h�;Y
�B~{y)ϼ�V�De�+V�G�����V�:\�G*�n�� �*��##���7��+O��c<[�_y�Q҄X���++,E�n��!WEv>����yҍKw �/�ɗ�dl�T=�l��Ĵs"��Q$����ϋ�AGbcE��&YY����c�f�<T���(� S0�����R�ŏC��ܿ�WZ�b+33eP��>A�-��u�+}I��瀪�>ڎ����Eʾ�>�}�l*.VŸ�׽�VYY�ϰ����H�|�`���Yv��`3�O�0R:E����u�_�u�����;�D{�����!{�c�>��Eo���=:!+��!����Bpx��g��u�=&:oƧ� �[ݲ�^�d��0�m�,G�hE���R@+v�q
10`�-��%����'&k>�y�jFZ���d�e^{N�:3��Vt��R�W�5��w� �a�ܶ�[��u4ʏxs�B��������9Q]�,}��&��z�E�.�5�Nv�;T�����e�u;�g��z*M8������P�_Z$U]��C�{��z�u�B*�7���-3)�[M�ě�:r���vW�%T�FdU�Qz��v��2�ي�BZ���]	Sp#@s�sSP쥽2���/g�]��o)�J]��V�]�m�O�uN��lsJ;�dC�j�{��s�~��*u�u���X��}�!w�ׂ
���W�
ok�'��>�X(��Wx�H�-P�m�r�g��g����+J�۪�[F�|��CȤ��1�f,V8~Ď�t�x�WwAaѸ{�sePU 5�p>sZ�!4�q�.�λ�՟q$�C�4[V�\��"�(��f��y�䀘=�nx�j�(҈�
�����O7iN;Z�f�^��v���Da)�UM4�v�������8lY5�8�;��{8���ki�tv7�`�/����������l��΂�����XMs65�Q+�-/
�X�Q���ԃ�چ�u��I4c����ۿ=�<����G�z����R0o(��ig�t���_�.�u�o���Ն=���}2�sr�=�di���n�⍕m
��0J���l�
�:�=��M!�m��oΤ�eU)�м��֥�2ҳ���gk���и/�`g���MC�˹ʚ��(�b�1c�5r:�o����iv�v�FA��$�G\�ItxN5��w>���V����K 6M%e�=3e�s�㨲�ǅ����:��-W�-}��_@�M��]1�r<P�S�4ܔu}� BU �2D<�	����Uh��m�>�����^�&tl.�O��B��t���P9n�F��RS�D��C���cN*fѭ��*�Ol�3Ӄc:��*�� �Y�LȘַ0
YJ�rF�7�5D�j3�u�&)YX��D��Q�Xa=����nD<'jb�������(�sWSB.��U>�x*!��_C�Y z�OI��fa���\+��q�3x�6f��%�ȅ�t��/`�<΋ mk�e��<d1��?!n��9�<����f��zWO7���iZ��M�ٿ��7�:���� .�~G���+x[�����7��X��eR���J��橃&����ʄ3�*|[���<�fƈlԹh��b[|�}��c��˗��	�~�f����j"�㯃�/pN���5q�쮑�DQ�b�*Mn��|4:%��P��8��tX�8j1��PtR n�~}�Ͻ�>Aw�����-�!��G >f	�ZY4OzQ�u/c�o��
�P "'2�9�c���-�<�T��[�2:v�y��m�8�W/+;/��A�֢�lsEP�r��E�]�Lފ��m^��5����� ;�yV����Fyp�/�Ѵ�һ����3{�h�~�F6@�;-��ߍ�W]s�!� N�hxT�@e^�㮳e7�+��΢%��n�0^[�8�z�h|2�^x0�C�ʾ��P������@p��m,z�;��*�x�uz+ڜ�W����ň�:Ό	�Qӹh
�l v۰L���Z\~���+���O��Y�e�
[LkW�x'���	��C�c�5�Uo�x�� ������01=Z)�2��X�4�[,\/UC����xݞ��}�?��kE\�u>��{�y͊�ڱ���w`v����U�@[��^����ܒ�h��}=��lж��qϷ�w�x�}�Z��?f�T�$1�����Ƈy0�n�B�V�nTN����E"`��}6�h�������߰�)
�ؖ�<D�;�4��^F���&�W�����S��n��l�+��!�ԑ(�.��Rb�0cG������a���6�+J�<z�F)C���&�ɿ[FÇ3j|��y�g�씝O: -Ti�T��Nܐ^��n}Bz��ay�ɋ��܏�.�AH�+�%<�t$o��������6��d#�ws�}ےk��2M�º�ڻ.�j^f���Ff慗/p^�H1�VuA�L��p|�t^�X�չ۲a�='f`��y_Qv�WaJo2��&PQ�rb:�e�-|^R��u
����t�����4���J
��f/�����u�3�-�%��`�GySm]������>@��Սqp�X�8+<<��p��!�O��
t��
��0_�)h�+�5�@S��Z�N�󿚐�KU�/9`)���n��2Yƒ�
����m	p��T[�z+��B���K�ԯNU����PA�79: �,��Ux�3l��_�5��HN����"�9#Dx�dYߧ%�����K��"��u�����^lP�hEv��~��Z��|����l��������Z�9�s�E�%�X�>�ņ�W%�b�Ï)'�?+�����@��c}�y�%ѺlL��b�,�%�]�M��m~�eK��s��ft>ّ1���~mKӎ�.i��ol����N�H�:ɽ�Ij�1�'Q�9�WS�puQ.��'�°Æ占%d{|��|]��"s]��x��3�Di�}�2�R�ۋ�@�&�/��[���l,�2�ҝ=�8\ҭ]�r�n���R�I��q�wQW���^P���vx�=�ra���u��9�	,l�,o��!�-��;�&�yggj�&m��Ds�i��� }*jޡX��I�ΗZ)���ɣl��cP��)�s�m(̼��s3xNƓ�KͬTQ��	��!���!�8k���V�}�Ī؟�hw'�@|�Ӏ����x��_��Z����s��f���2շ:���������*���Gx����5�c)����uH��؜�h6}�Qw�P��)���c<�N�}�Q�[v�F� ���E��W��@6jWE( =]2��?�"��yP����:�s8�i<��MOȀ6fm�w[{伳���U%���ԧ��|�3.�����]�s�ꏹ�r�� �D��l�gW�r�:ꈻҰRot�ҷ^���*~V�+�%���fN�n�2��u&�Y���'d�]P�7��F���j�+�7����׿1J�e��}XhicnE�]DG71J�wA���L0�ܩ�<�
���!��p�L!���&e��d;[}E�.67	ʽ�,˔b�_�:�����Mk��˪�!��Zyz����J��W-n-���#�)�+��n��`[T��u�k��X�
i㮉��#mb��>�DN�#0�݋���h�)�.� q�%��;:3c�/]��q��9Vtj\I�&u�n�>�;���;̉Gg���[��������E-��HE%������_�WXْt�V]���(���C��O���wZX���.�X��<�DUQ;4�yV�먍Y�P�4�(��r�d8�=�i��M�4��B�E�S�80W���Z �+	���C������>�/x�w����/��)j��,R�9c�S�(��Ϲ^ˋ�n�{|��ؽ��q�ʧ΀Ux�E]w��0�m�|�]���5FG6m�b�}�huJ�͗s�V�w��B�y̍/z��e0F�A��Y��+���r�+�P6g��Nm��mPF��S����й���ݍ�u��}`���_�?���Ac�N�1�Z/��`�NX�p=.J`�;#%|^�ƀAӏ+^)<���
�$���O��5���V/������y��*��GM�&��EɜK��=����x[��R1�Ȧf[�jpzD����<<��{��
��|�idt��\_]�����Q�X�5��(8y����7��g��ڬo�k��\��7x1�5$�]=��tZ]/���d�� 5�z����e�+��29�<Ga��e�V,ڔv�8��� � fAk2��N��2pέ�hnU��]'��އI��9�xn^�:���7}���o=Lµ4��أ��Hl�ν{/�z�à�u��;�q�9c�v!�6_,��3Q9�^�������6Gל�w��<�cf�"�����pg��jY����K���oTHX@���d��j@hܹb+�h e��;vc�AQ|��|�a�=z�$vs�U>)_y�m��u������ߕ50�mEO��u^�"�h�6�e�h�����s�m�'3,����W9
�t�j�ڈ�q�p]P��u ��)>�B�u���p}ñ�s�1v��?AU����,+.��:��*:-LA/m���o��X��ssO��h%'�z�����/t�.B�O�/�L�Z�C(h��ׅ)����e��uٿH����P��\�h����Dg��_T%�Q�^x0�C�ϭ����uP�6U��7��V^Z`�/t���V��a���_��`��D���%�݀�zWo��}��\�`�fN��{�װ��p]�|ܦPϩ�xV��u���9��N,���&�ឮ�$�<M\����pz�̯j�~����V�/	�1��w�Z)�$�X��O��~>��SlÈ�|�Z����o�;�|)S�O;�}/�{  ��䝰��5f�P[�[�>�J�v2�eZ�,±�fa��������|��t3��9�o��)��dr�,Ԯ"��au��h�/z���{�y՝�(�-�]��"�բ#��U�Dؚ��[JL�$�r�sªw��8u";�.�>�2�*��Ȓ��ݜ}7�q-�T}�f��KZ|#�I��;Pu�:�K認c�ٽ��( λ�N��*-Mh� ��-�@XT�3u��(��b�}�E���t�5M	S%�XW�t�ݒ}/V���%�9��
L��)`�}��F[:�hh����]��s�%���X5��"L,-��:*S��Z#Wd������0\�@��v�XjVSb�Dwkm��2�0��s�41�c���^��q��V��I��/��8����-.�[�	��N�҇]I�^Y5��/Vk���v������-����q;c;�P�oZw�e�D�����sr�(L�y[������@��3��n�H��U/��We��%���{(�#ݜ �l�����A�ռ�:�Z�]3�ТN-�N���%]r�0�&��*��� \seE�nfm�]����\����\-�5�]@��:u��P�[6�Jݯ�,D��~g	�xőnc�瓃�w�ѐ��ΧC�^4t���L��NUb��B�1�ص�� �E�mو�#v��b�΁NVfr�7�$�i���paM�%�N�[��������D���]�.{p����gFc�g�o���f�wvL~�ѕPt�8��t��v���3�T*�h9�͍�0��b� �ٔp�#�51q�sr
꾦re^q9�7N��W
h�&�����74�0�!.�#�"h�E�v�t�}�ʵG��d�ev��u.���%یt�`���fZUyi[4��#C) �����j�m�!�{0��51F͡�{L�����w���S�#{Vd(wv=XI��.·n�Dv6��b�{�N��=�
Y1[���U�H)ȶnL�����(�j3/���Q�֭��![��{������S��5�.�)�Q�LG��StH�3 �e�^Ӛ�����Jp^,���Ժ�����W��1��o�����ܚ����C��Y%����9�gW�>��nr�"�x�/x�v�W�Y�vea���H�=�t�G4�q�r�w��On�;R5����Z��"y���RXrN��JLy����\����4(-n#]h�ITMV̥f�/��d�FF�R��x�����K�[�J7BK�+TIIc�t��V#�<r��W�vU����~����h0�X��(�p]E--#k���zV9P8�(���E�>u(�UiWZ�qq�S:�Q�z��SHR�bbή.H���	�Q�b���ĢK����7�av.��7���;k@WP:����w<�(�q����xü*w[f�9���X��"�����oɇ��wz�M�-�Җ�D#��+˕P�%�Qih�.���(�����伅���]ss��:4R-��JꆓBQ����N�O%�����t:�됅:
)l�s��rP����n�N��N��ӡ4[#�%#Jng*�*i9 r\���&��t8�����C@i�%+F��9*)4i�Tæ��Д�-�%)�)S�-r�� ѡ@:#��<���(j��F�AHкMS�N�H41!�4��M!�4�xIɢ�K\�MrM�'"�����ht:t��(�:F�E'#IȡJ
(
 �et�Ӧ����h4�h����������ѻK.�ű�\LXVo�p�Q�I4jX�Dt��k���N��9V��ѩe^���`"Y�$���7�둩{����#�O��9�]y�������,C��yo0r�������x���Z����;� 4?���&�`����w	y���7u?a�F���|�����"4�1�H��/|o�h����g��"<��r����h���.�󾼐�z�Oa����_!)�?���iu@tHW�?G����r�CN�A�u'��9�9>A���|~� >�����h�fu詏\�̫H��w	`���O���]��C��C���|��캮����z�I��:�5�YA��|��c���8�����c욤)8��A��_G�<>�W�烝��Q���ˊ}$G�<�^�z�O�~ܟ�~���U'~��u�i�<���� ��N_����˧O����C�%/�sʞC�����(4:�>����ܽ@y)�疖�>�ُK4���}�����H��>i��ܩ�? ��A��=�y����~���!)�N��~��<�����HD>ߧ���/W�
�{��4i����w>�pr<������G�j}��	ty��"��D!F>A�%A�?��O�:���ï�Լ���w�A����|�^��޿to����w��:{����J}�/#K����A�HW�������u�����z�h�7�Zɧ>���H� ���_;����A�u���g�}��`��GG{�>G�9	^_�r
}���>���u�4r���	I���r�C�?��ǹ;��C�k��ھ���G/ܓ���} D!"$`���z�B^�}���{�
{��\��_$�׼��~���u��p�����O`�%S�����h~A�$�A�u߻�ѥӣ�y��:��K�o]]�6��ň�D} Dw[��� ���u��`�Q�^�w >F�<��׫O�t�2r4�nT���P�5�_������!��I��#��>�<~���>���H���-�չ�&m]�� } G�0}#���"
�w����>@h���<�?'�9e���w	T������>BWp|}����?a����A�u�?��������wݣ�Yy�i����r����B�8b���[S#]fJ]��u�u-T��_�=	��ڝ��3����1���	�� 3��z7|E�nx�k�UN�-X��u�)�����hU3�^1��[5KD�^7���<WsX�9�A/%���~Igў����r�o���v��3��Í��ö�������G�0���<7| ��#�L�e�iuO�켄�d���G��I�@y���=�G�~�/�ΐ���������{�����A��$>���@1��1H��G�^����w���n����G��u�y�������w������~nBy��������y/����O�y/����ϜS�?K�ι>����̋���]4�b̟oxOP�G�J���ţ�A����|��rGQ��=�|�.�����y	G2{=A�:N�n�� ���O￸|��y�o����O��{}���=���zŤ���k~�U��.~`{�	�}������0�����׸�����K��zu��!�~��Z�����c�~��ϙ=�����/�}�P����x{��W�>y�џB�۸��9�>��]��� 1i=��::��:�d��;����~�����`���_:^���G���I���g�p�|�F�U�̇!+���?G��d�$������$�~ʲ.x�gӢ��V��F��D} |�F�=�� ������? �<���}�/�h)�y>��C���{�%�	OQ���'q�����I�מd9i��}����N��=K��;����\ǍU��-��H����>��@��7��/��A�\�����w	O�|z��C�C�}�PcC�=�\��9��~q;��4�|�粒��B_}�i�!�|��p���|�㹮�Ve;q[���",G�"�G}g赃����p�)}��K��2����=�-�5�?�p�>_�4��׼��_��J��p�.�/'�~=�� >B��G���e��ʇ�8�����W1�P��A�?|D����9g׬�BRGGy��<���]��>��OP�����u���}�NBPw�޸^�4>A��<����>����zX��|G����s�*jEy�=�������{���"��+���<���?I�O޻���~�I�?���w	O�}���|��J:�'�������M{=A�@x ��AP�F	}b>�>����f��ecNV��+�V��t���fl�B���&�QN��3�!�{�`MB*�q�������c�R��81`;f����������V��5�����f�t[J���ԥ�;F�uq��X̭6g����9��	�� 	��vG��^�����F��t`�9o�N�A���_�ʓ{������5�䆃�?�G�����S������`���<��C�>�ן>W>��y���J��@>�!i�>��=1��?oa��}��uO�wg��=��?�k��|��I����~{�9��?$�xw	G��_��*>b �\a��<>�"!�°�[V4X�Gf�}W���>��b��̏�}�g����B ��^Op��>yë�>ǰrF��ΐ��z� �_~pBU��:N�>A����u̜���;���h?C��]�~o�O�_,<,��S��D} D`��1�����=�7S�]������K��}�����<�%Ѥ�矺>T%P�s��?���O�k����#�x�����|��V��U!__P���;����6k��<�V��􏈈�"$}�E)���t�_nI@y��u|����Iʽ����>AԚMy���pu��>�߷w�t��q�?}�� }��>�h�:~�<��цk|W�:�9�}��}
s��� tx}���\{������:�>A���N�_���|:�P�����Rr�i�9''��<���NK�� ��:���#�"�CJ��{��}�d�0���u��Ͼ{y���b�����C�x�Q�^���wR?�k�~qtu}��~����������=˼���!*���:��{=�W�>0r�}��pDFI�Dp#�>�>��ٵ��~�~������;��=��d�� �?>�����r�����=��u�]��/p�>y��r;�
�=���t�����A�:t�_n��?%ф(��P>� ����:sy췝��lw^�/�?G��O�b䆃�G#߿8�?c�%>EO ���tj���}��s�=��:��
z{�罯�#C������^@v���S��~���~�>�>��������/Nr;��χ��>C�������CN�������윫��C���'_�'������9	z�ӡ���h����4�����J�/��@��  �Mf��=x��Q'�k���e�+��UE�����w&�ad.���[a�%���Y�w��k#�ڱ�P�:kT�V8�8����1��es����p��ĺ�GY�%����ϱ����F ��Gk����u����j��2�L��[���_s���i�=����9���:��;�P����uy���?���s/�P�>��`��D����Z��(\s�*q̑�9e�f��Ij�f��M��ņ���<6�	}�w����A�������߄{�5R����/`���m	c������P�#.��_LN�.���F�7�1�g��M��p�È�mת��;D]���| ��t�\}p�H Gͪ+��y��U5�;�2Y��6�>�e�Hy��&<ϣ��_$�ٶ� �.��#@�\��A�b<"�.X��b��~�����~���2���^Rx?�z	��9P�=����9�d�_�:�l���뵒xf;�2��;�a�Kf3��E}�>;|ݞ�����,]�L$c������>I�U�HiDQ��S�`V�A��< ����^Y��-O�w�<:�(bra�zX�R�"ݥ��	U.��1y=)c���Z�y�� :�S Ap�o��1���(iP�ui*�C�1�z�5���b�5�߷�ha��k�&e������^Z�p��hM�3%_��E��87�Fb��5�����?fz�iR��d������;3���ǹuq�t�)��t�nhp��\bT��!�3vV��	6�ʧ�����o.�}o��y�K�k�[��	�告��
��X|��,<��4P�3i�gv��ne^�|C+�;d�0���K��r����}!֪�6lL�w��WBR�沸���c��,��ª���$2�*�X$���r�Zi���oLe�'PYۇ���5���κv��=}ʧV����`*j��Q{O	ih����<+�l_�$΀��ڴ���S##6�A�O��k��r�s>�.`v�Sv�j� ���J�� �[��Q�5
}<���Sҥ��FS��B]y���^{ ��Srv�\mK��6+G�U��`��8㛗������;�}wܥ��81�|����붫
k��穇G��������L��p$��������_�0٢�N����@F!��R%FؓgM�T�h�hm�]�P#qR;�?����^�j��/i�M"��06w� 盢�U�s��a���:�Ӟgn-��F!!�#B��F7^�P��Ӷ$���l3�eI�� ����BHi��INY뜙ut:;eC̘����t!���2�=�d�aHsO��1����9��G�Y�^�74��W,|̗-㐋���8�;l�0+@w�p�ǩ��.�p�/m�oLe=�`�|�zܞpvw+o�Kt���鄬���78�[A��َ�<��v���.��
9�o=v�
\��̣0�ѥ���kgeX������a��+�[���ċ��y9�����
�+�6��jB��^ÇWG���](seG�n��n�;qd1_)�_S��K��%,u�e_�����x�%�F>,U��;]��.���2mK�UAD>�xݔw�{�8i��l�k�ʫy+n�����ML�m�������©xk�m)��n/b������w�5�;�y]��õ���[��\ʴu�S���vצj ��)�[��E���oxt�P~���@(�\�{}�]��KӘ���k->�m��V��W3��L�+�n�g��ٰ�yC!MK w���wO������|~��x/����>n ���*��%�}����.2,�$����Q=G�u/����+�M.���g���sU]�}(����'y�K��,<7<�]�ˊs�8��Xl�ێ��t_���Q�u&^9�Hc�~��R:{]� ۟�O�.*e����R��m�����XI�G���8���V���6`N�҇����$���ӆ{Z��>�{�����%���i��k\�;�1O58s��;�۬Y���{訫i}C�&�\�zG`��0�� �8���ŕ���ɭ=�N��\n����vWVw�Տ�l/['���)��э=.Ɨ��O ��o�ݶ�5ƻr	ͳ~��`�w��=�>]�݅4OVl�u1�c�y*!l��g�"���Q�][wW��g��0�*w\L�%���*�l#�`7@#�\���nA��fb,k��_Z��M/�c�_/���pS}x��t܉�#�2.L>�h�-��qxc6Ϩy�K���2�~÷�]����?*~V��<+���c�(�<���sxe:��~�9A�(E
�Z��)�f�rt��Ա����=�g��+K�eٖM�vUԭ�
�`�.lv�{��d�C���<G*l�6&F�=|��^�1`ڋ��ZG��;��:�3��e��sUc�	���Mk��u(�x��ʜ7d�2�@��Gc�%�=�'��U���Y�P�xB�:�taDw�f`����ItT�e�:��a��3Z�iM��C�#|J E�*�D��C/���{8 ��}>�Ў]�`�D�kk���9Ql�⍺�d\~�Y>5jUп����J�e_���Hp��}3%����>��n���/����wZ^�W{mId񢳝��\�"�O}�[�E=�wA��n/>��QV��&�97����J�w1�M�v�� b�+xlN�ܳ0O1���C�;E��{��j7r��Cj��f�P¹�������6��0�s������t���s�|��8�O�y�\ � l6߼B*m;������)񚅒ʻ���{8�&ko��h��l�����}9=�*Ю��5~^���L�߽֕�Uﻩ{��.����]#�8ݔ�@&�e�;V��+�젨�I�o��kM���%2E��L
��ьn��|§iH�0i􍁑��a��Эɛ����r�^_����lz�R�G�m$5�%�'gD�3҃~ο%!�0C}fU,�L��x�r�����3��!?W�R�WJB���y�����~��lu��x:�/���R(g�[8�����
��H_[̂"��F|܆�I�rhT�k� W��yzu�>c�!u��+�z���Eh����/)�6P��y`MD,w Q���?!yn�o|���b���m�q(��fb�!^T>�s�6� R�q ����(�+�7�!�zᜉ9G-�GGvW������57ҡ�Y�R!��к����C�nfX7�DY��x�S�g&Pɴ$p;"����\�w}�V0Q�-�׻-��Gǻ:�]�M��&
��'��P���!;u��vsn^���Wq�������퍧�n�IH1����5������Ƌ���x��в��k`�Y�[�4KìZu�Lh\����O\8�~���=�y���B(����j|qp�����c����p�W�}���g��5nٹR���D�]���/�,�~^fAK��@���kqmu��y��V�\	�BLZ������%�uʠx`I�$4Mi�`s�nz��ٽ��}6L���Y�K�?���<����W|7�Ui2�*"�&�DX��\��;�|��j���+��"�&e�Υ����}[6m:�M�^�+��5�w[f���,DÍ�^9��8=�S��6����p�يՈ;Z�R�s��%�����칵��f1���8}�|~���Ӕg�j��L��^
r�Qa�R���t���Wp��K��`*���T\�(a:)�W��)��}��~:g�]��j0��.OV�{��/���~�}\���m�	���z�Ǟ.���	��|0�lnX!�8m��+6�$z���`hS��g妾%@YqU!��;��5HT�%��yܛ��fL�#����|�J/��#DJdT'Neu�C�}����=�@jA�M�n\;��aG����5�{T�����`t�ί{sC���B���9�B�YJ��o��թ<�U�@�{q� R��3xNr����i�3�o#���w��ǰQX���t����4�S5�wD��!}ʹp�yV2��k��pI��o�1�
�lu=�����.�~�_�wf�}����D�6k��x����Rr]�gB�*��0e�7N/n�juw_Zz����[;�03��^�����a�H�'��� �eF:�1p���ݹ��x�ly�jlC��#F���xs`Jٸ7��=t:g�ͫ�!�(C�,�7U��s���{���c�t��j�\Q׮[����]<a����C�\��+�tq�^.5Ɲ�!ɯk��C��ٔ���m[���]��5�9O��ͬ��\����&\v\cΔpyʡ��Tt���B���#�~ǢN���m��=�@�/=�J�}���~:b��Wî��UD��?qC&ԨĮÁoi	�p�a�P����O�z�7�9�j+k�E߷ �W)����o�9�}�u^7��׋���j�([6ώ7hchо��eLv�[*���U�]���kX�bǩ�NϥU���g��N�*��z�R���+o�~��b����	�ݖ׵�!�t؋��yX�SQ��qd�ҳfG������6>����m�L�Or�z��!�Gc0��8����[��2wX3sCWw<w]�8�:�Ž-U��Ƭu�0�b<�Y����\�[l�y���;���+���Q�t�ge���L&�u��O���������q��Y��^��%9�dʙ����ջ�\� *݃�=��[)�Kd���E���!ܨ�K���q���fZ:���-��܌�Gr�NǓ�n<�M�v��OW��3xF�m��("6sK�`x�2��Yz
���e�5�ƤrQX��Ўڕ�W�ۂ�WAT7]/y��Rӳp������!�mg��������\��5+&��<���d�[x��+t��c�!b���dc�YX&$	�M�vN�-X�θfZ�,�2C�}���]Ų�r�A���Y��әs*nniU�V;ܣ�U��s^#غ}ī�P����pg%�n�U�p*"�^�.pz�zH�I�ZO5q�H��)��;ηG^�!��n&��v��Ԭ`K� �=�+;P+��)�֩�ºcGU�I�S�y�S)^��`�Z�$y�����$ZWI^`:��hכ�gdތx�.v�S,D����jxJ�eu�k�!Tj�I�R�$sz��`h�ԝ5�f���mA��]���i��t��(x3f�*ʀ�U�P}CUۚ����x�����T���$��7+E��P���w�{��=�c�gAY�RH�e9����"J��g%טرFM�*On��yh�=moMw��#O�K(�g��',���+J�-���mR\һ���� 0S��v%ԣ"���u����VZ���z��o@wz������h��erò����v�f�Oq�(��O�e���s�ؕ��������z�O;�r3�{����c�Ik�J�g07� 軩�vǆ�I�	�۸�XT�-�䭜2l�N�M��"�I�8Sn(3����8c�
�@B���:�j��d�*�=�t��]}HS�f��(��+����v�.�։8^�s�K��0��(�}ҥ>�i�5N<9M8�W ��d�NU�k����N��~
������n�&�Ե*!�t�8I�mC5t��<{۝���s�m�?Cm��^9��icͨ�7I9ĤGrEPȻf%�ǖ.F�k�oY����l�n�dp�Z��"��a3ٜ;u�����}�QJ��.;2����,�����0[S����G$
,Nx���]��k3�Br�
�c������6�|�L�.���&��
D`��j��P�5..�]��k qh�Xo5����5�I��0S�)�{�P�G���#w���
q�C}�I�t�N�����!p�a��,��F=��!���^�:�gm۲�ҝ�s�n!*�y�^=�x�Ξs-av�}��g�`
�Yj��
�<D������Y�8�U�W:!-�W�G�բ�u�y4���A�y+AZCE�1@r����ӣ�5�4��1ˆ�N�@�(�M-	�F�К
��(
y�#l%��M�-c:��̇!���D4�"e)*���%�D��N��Im�4j*�)��K��hh��b9���� [t�9��
)9:��U�ٶJ
�j4����kl4i�IV��4�5�b��M[:ss���Qr
tM!Z�m�;dt�Q���N1�B��!�1�9'%i���s�4��*���(�4QZ�Q�h��EVֹ���9r>sW��9$���=�݊���-u��{T�v�p\ �}�Γ����pt�]�(#֍��t�X�w��>U0W�UT��>K��T6��y�*��Ο���p|jq�)�k<xJ����R���J���{�w��1F��]��jّ�*��3�ƈ��C���Z��S�~�)��:��6�ďy���H�а�\a49��1tS����;uশ8��r~K@�S�~��4��=�xO"�����}�u�����IS����"8nlgζ��/*$+�"
����v�s��K�g��\'2S���T\�9�i��&�ʮ�e����e>˨�l�z����OM�3�Θ�9��U*��4tu�{O�xXv�5�������ʥrV<y^_�[��B)�lV䅪�>��6�/A� yP���R��^&��t��^×�<-���+����؞�����poy�b��D.L���@5�����=��9���d�������c�y��7-Vn����Ǧu�cf(S���K���0 a7Q��o���/Aw��+�oG�;]Z1S�|�z��t3�8k�Z�v��00L7T��G*l��&˞��֏@᭺)5���Y�J�Rsݰf�ču9)Z܉ǒ'69p�n:��+���}K�XDl��]���x).��ޔ\�w�ykG���ø,-�n��ݶ.�#Z[�VYۀU�&�{���3W��&p�� V5���*�(j�=9e�}_}UG�ƘU�r���j�4����xLU
�|kώm����'���o����@�+HRX�vp�����I4ǆбn�[�r���ó*��x��*�n�_����!��ڊ����2]N����B��k�V�#0��
���HU�Ɛʾ@.?=��4�뻩v��hM�h�^����nieh�������䘱S~̮�nh� /K�w\��-ً�K{�S�Y\o\�E��N�n�Y��{���1�W6�=
NU�O����5g�ӝ�����bC괴g�֞g�*{9��9C�pc
�Zc��P��	U
k@�5O&�aB�0�_��/.��Q=�+`ąƼ�P�J���a 'N�ǎ4ە&�	_5
ݮ[֐��kr�-�~��q�Vxm0:�o1�^U�r�`��u��l���y�O���K=3X���p"`n�C]%�;f�<��O�p�S��W�Lb8V�� ]��t����U?7Q�~5N����K4��P�ה�3O�pzAH���}�'��
wu5��s�/�Q�F#�lPf�Q��Ahr�;��,��h�1��q��=�)�(���d�'�k)��fz&�JH��nM*��}Y�vη� B��v��q�M�8�v�bW;j�d�Ӽ0h��Q:#�B�����H�v�3/�蕲�xm��� Umd_�1�KS�I�.hT�}�lP�f��f_�s�)Q#5�&4DǛ��{V�AyLAQ&19���i(a�3�T|�A�k�8߼��ʐ[a`B�+/>焉�K�m�M~���� �'�̾��K�ǖ{�d�\9�X�;[ ���ܷ�8��Y�,�b�����^�RVr�����������ԸG�8�rp���N��YG��<��ǅ?��N� �g��/|ê��_��5��:.�Ju�魦]y��WHj"n4}�j�\C�< �����E����"=P������b�D���3g�TC�?e���5Y��6@<,�}��u�i�$�c�6)n�+\k���@ g���qeF9�n�7]_M���5��lL_h�HWS���1\�{�wt�(�������2���'#��7-;���0W��G�׽D!�����W+5e���kf����f��U������ʮ�g<�'=�t:,�j�xC���\�u{k�����oRƱ$���b�]�a<*��z��7��܄R���m_7c5jDDsdn�������;���{�3� ����H�f0�93�G���T����W��〽>��}����r���*��ȷ|"�yhōJ�C������?&x��Q��*���Q% ���^��U�0���� ��=�2��D`��uoU�n���Pe�t���LS��N��7`/�� *z�ܝ�.��X�}[����o�XGx
>��O�����r��ݼ�0�`�"�+�!�)R&���y�"1ї}w��,���FN�8��b�L��U� W�ۜ��F>��t�1۵�?H6w�������.e��޿(��	U�[}S���^ƃ��"{��഼�����78�ж)>8u`�>�Y�M_�Z�aG��-^���Aj�	�}|k�����V��*p�k®y\6�����OlJ��I����n��^fx�ОU��k;�����q��z�3��j�d�u�uc�^�p�ϰ�^jd�������G���R6��<IXf0��|��"S����7�?��vk����r�V�H�Oo|�N]��ե�!�ɰǜ�d3ZM�{͏	�(_ν�2R�rR�]d�=��.�N�X;w��o�i�Ի��tv�6��qGM������瓡6���.V�X�l�L��D.��mhg}k/���A�*S}++��J4jk-��l���ԯj�&�'|�ܹ��sr�4�����]u^%��)�y�_NVR�� �iB�<+?�����n�kg��$~E�鿾�ր(R,W�U���qFp�	�GBɞ��]D���_9�wT�	���131n9dk���i_Vt��z�® ��8�[�f͋��`tjBz����m�Jr�/%�±�R>�����U�Y�a���[�s��t*NWN���2��ص����{��2O��u��>�*�^�Q@v}M�k�U��@\c������M�1�ۘη�!�1�3�����JDѡ��d����\q�ǔn �x�ϭ*��\5��-=�T.�#�)W=&��q���>���6�fh��T;��J����R�`?>�%2�d���n����%�w�Ϭ.�@�����qA�����R�D�J�ΩD)Z\����p&�;y�v^��b{g�ry����_�$�)�j`85���j�d�b�=�('9G}S�S�����,7{�pf��#}As����i�'����tT��.�_a�iY����f�/���ʕp8:�SzK�^_ǖ٩�]�4zןO*����Ny�0�sI�˞T�f
82�D
���L�m,��W�;�.��~jۛ�f��+=k0��׍
*�*Y�Eo�GNu�X�|Ck��c���[�6B�����j�!�q��vԂ��H�������m�_�F�V� ��zT�Jdmi2u��3��=� m�Upm�R�U�U\�뒓���k��_[>&���aߺ��o�9OQ����0gp����z�(E�n�M�!��"��N��o��9_&��n���o	�S�YE��+�R�񋹟2}�|�
Ջ���,E
�5@=�5C��8@i�F�=�ga��uө����rj���@ք��U7�6��͎�ݪ9Us����uN�����c&�)ГƦ�����g��x[�^��j�ic׆�����*�I�5�Q�5�@ƝJ7�~7KeΪ"��%�}���WS�$Ň@ч%�ϣ%�Vp(n����gӤ�{���\��&;�/VSo{�ϕ��2~T�^3f���Fa���e*�!Vx]�S�}1��� wA^��X^-��q�=}op�����n����qyU�ؕt/��c*���:3�O:ڮ�Rb^UFƿ���yL1�X��~��KY:����}[u�����y�Q�Q�'n*�}@A3�.�U^^�P�p7I�.��AW�8wZB�}��/�j�kHѽ�˔$��A������%X{[i瀹���`�w��9z��V��.�"ܙ/͋vL������Ӟ�z�'��)f-SQۧ���v�����y�w��6��1慏k3)+��]zXZ�e��t�*!������U_}���V��_x^��f�T��&{|��!�.����҅ӡ	����Ǫ:�
���T��.8_�� �!�\�ԏ(����c���#�O�\�b�f��];�É�(ό0����|��.�8�P�4���z�*��u1��̡J��s5Ga����OX���P�'��U��&��A;�r��.�қ�i��Ё�j9�/�r��X�s��a���F�y��O$�u��0�5K��>喐��WK��ʁ)�;��1�1���☤�V�AYLA��G 
�<����!G�j��aSX��w%$Dm�1����u�W�6K�ftL��j $���{ =.%��-���G���R�x�E���|+x\��d^«%��F���\#���T�ďj��w��)��vC؆�(�CQ��>�Bφ᫳�+�<���|�ǡ�f���˹-�܌q�#@`�U�W�V�"�^�õH���+u���< ���
5���~[o�i�9(JMf�A��eNi�Y8�^-?A7/,Kw��⺮�&�x�H
�4֓]�̩�(},�Pj�t��j{kB�x��P�L)^Ӛ���Q��K�{h�������� �-W��YU����+{em�6)�w��jf!
M���Pax����?C�� c�*s.l��lR Tf�� =@�y���z˱�����rU,@�����<�H�����4L�Q���D
�w`ʌs׾o��\p�o�ؾ�����V*�7�o���ė�{�w>uc5�`k0�-vɸ�0��"%�Ӂʎ��ɗ�2��x��,"��KWNiz�+% ��zW�֖�5��3�p���ei���4R�N���D�{�|�<yDi�f��gc��
1&��Hq{O	���ҫ9�ΰ��&'̄��)E�܎���3��k���6*�Y�R�<u��7`3\ ��o�;Ơ.�s���]���:�-5j*
��b����0��ڸc�W����C�P����J��P�͔r;b��uQ�u�&;��]�,t(�NɝlR���6/��$���+�
i���B��/�%��5�X���O�}�|�\�+�=�^`p�F��P�E{=PC)�����o���Y:��0X�����J�#��/O�p���&��/j�s6����@i>�P�B�IP�,(I��2�0��VrJȍ�oWo=84��D�#��I=��D@4>ԡ����hKLz��c�s0).��f�D�X/���Q��-����;ϓ��{���Z��܍�ށ::{p��?}���{�q��Nj�eY���6""����Ա������K���W�hT�����]��I�J�f��m�1w�w��/)@��`/t~g���h��t����c��D�Lz�:�N�)B`,gڳ�	�p�LkR���0;���7��U��p���A"�����i�d��u�����&�X0��:�Q��\� ]�?n߬װ��ks�p3�k���K�A=9�ז��Z���}R�s�c� ٦X�J����6�a��"�|�T�*��5�P�cd�/{:b*���ZX��R�k�uG���k~Bq�?\��&t;�L��qnl���i�NJ�x�{�
����iϕ�"<#���������Q�:<�@�Z�p.��1�z��b�ǲ�m�n�4Z�+���7�1�3��v�7�n�1��J�ʴ����!�b�Z��#�T��T7����]�=ޗM�676vT��HJU`��&�Ǆ������!<�=�s�{�<�әYY��<j�lg��l�����
����UƱ��0�J�j����1իx��1��[S6������gĜXxm73pY�ӵ1h	N�"М+lS%
�#�/���ހ��0��gޏ�����5�����T�B�YR3-�^�i��J|���5.�]�n��3���ԩRT�&l�v��B\�rԎ�d������%��j�������÷�⃖�A��˨�z:��,s�:U��)��*�:��GL�D9�U�=1Z�1����ig�ağ�`�X6S+2al�=~����G���T���,QT�j�yW��Z�Gf�����uQ��D39�\���i�As��20�
v�Jn����o��çQ��Yf�N�q��"�;�e�|`���t��RlB��:�I0���8��
��r��>����A�X� �݊�1U���@�4~��^&�b�.���fPp�mB ��7H���ƥr)����IU�����h�Ҩ�U���3�ߴ�ҷ]���9h�}7`�q��(뺖�<|,n��f�
a�����c<l SN�Hɺp{���*�H�$kE����Xie2�`���R���=j�n�n�xT9�3FJ�2n
�T��]����T�~Z�7	�2[��ZǊV�����A6�=���CN��W����$�p]D)6g���e�������U��]Y�{ˮ��ORqT��,K�o�c+�,\&U�c�;y��V����ǂ]$Q��n�&�LW�YƇ�/������:�]���e�ȖAXP�1����a�Fm��w\�Ӧ�_N�x��[1Kmv�9�+'f-y�۱4S���l�vs"w$��i��.�7X�5��z9��覾��Q�h'2c43�K����F�S�O�5K������+h��nm$�/�r���G�{ɋ;��h��(T���ـ��<�|�=��e;S��4�kOr���3z���҃K{_4�%��ݪYo�gW^|p�*�{,QW�R�z��@��A�y�`ʼ�&`�3���l��y���;]��i�}����Ӻ=�I}*���%��(Z2	o��"������}(�'jk�l�PX��q�@؏1��wh3H4l����Ţ�}mR-��ܱ��\�g-	'^�f��U�ۭ]p���9g,-����EY�vy{T�B;�G�m�`�V]pz�$�tQkB��
W7�����(A�&G{��//�����/Y���i�r�*ǎ�6���X���ǯI�]�-hj�s�,Y��� b��įz)�h:f��cd�ۀ�v����U6A&�����C7�T�;�1��W>�r��|���t�W5h�N���f�2��L��Vp�oyS�u���˯�\�)m��o��gH����`�]>�/Y��1��=$]®o<yy [+9!���UȜ5�S��S�����v��U�ĞOfŃ�fő ���m����3Tvn���e�R�7�&��*�
u�S��NDڽ�'�A������h�x�8���%��M���͓!ڼ�x��:�I�٢����۠����ֻ;�Fi�eX���bX/{z�5-FB!Ȏ��AW�/%`���[jT@*����Q�s�	x�+-��P�Q.�dT�꘦_Y[�5���Ȋ����-3s3�[*�h|RK4���v�]�x�wq���5m�,:&޿iѕ)�����뙊>�S��YZ<�)��:�ԪB���xM�0��p���Yw�Uڲ2���j�od<�v�-�!�7�[��m�V	1DN�K��@�u��rTl֩��9´� ��}+t����ҽ�\�]�J�7 ����w�����Z'�):A="�85��5}�E���ʶ7����ז�:zE�M�1	j�n����1����:ǚ	��2e�k�m�I��ck����UO���IK1M3{>;���;�WB�y�L��k=�ɻsTg;a�m@�v���\�,��q]#q���H2X����ލ�����7Bm��%L�����Coy��� qi�����Kc�/Q� c��K
3FY�ƽsu���^�c���cv���)M>�pA����\��o���o������8��U%�i4Ri�F���)��i���К�H��m�P�u��
��4�B�B�ִ��1:60Rm��kU��颎C�I�yrĥPhR�-m�������]���F�]R�Ri-b��V�"t�-4�[m�Ѥ��咀�CM�hq- �Q���TE��4�:+E&ч���
J�h4TF�l�%%KȤ4i9'9�m����Mk$��Ӷ(t�Bh��ci�ִQ�lV�("Zv�ˁ�E5N�M�Z�m��-c[m�p�M��"'Z���h����fH�� x�~'�n����x�NxG��9�o�y�W���m�8�oG��H���v�|����z�NxK�R��x��lO~��� x���)49�����Еj6�bȼ���1Q�H��Ĺ/e*�D��W�L:�����v=�4�6���W���]��Q�q��θk܌��y��Fұ�
7Q�WRJ>N����%Tm�]0��u�q��^>���(��c���� �Ř;�.ԉ��%̉dHᗙ�(w���ɘ.reAr|U߬GO�y�rK��s'��hV�'8��3&T�}ϒ[J"���3UF��U-�P����p��{�Ӗ 뗢��S̓�2���\Q�~wp��;�MD-�]�ܤ+�Z9�з�ĖҾO��^��9Zh����F�Z�p�:�6ʸ�����OȐ6~%�X�p���D����������:Ko�,�6�)���� ��9�\�q��znbX���Ji��9�Cu��_�7~R��'��d�XL�	�K$={;:F>�ʋ9����A���G=�����|f�C����zR�<����o7�B�ӻ)ȥL�+y���VE�3���'D�hD{��m�/w��^U�h�e��3��w�%���%g���"Ⱥb#�ɜhi)�Bw�G��6zغ�d[�'�i�U�NȴS��"��1���'r�;��iI/�p�㉅1�y�uy�&�x��Q�(�}�G�G�~a4��()��P>Z}s>؆//3���)8o�wzn��nħ�.��z��iV�5ak*�Ԥ�f�Lo���O����.�S�}�5P�Ǆ�����0荒�ԑ:ѭu6�}���{њ�j�\W�~v1u��22���7kock�G��v������ضw�3�V���Aqߏ�m�
;�NOv�wĩ�ڹc��j�%c�y���o��׹[dz��������Z��$��#�2���ƾc/�'>�o���U��:�m�'�.9i]�4#+��k�5i�̋��Ld��
=/l"�Xƙ�y������]jd���\Y���<�`�`�_5~��~�e���~m5�&�;!'�9j�^���ޞ�^����I)�V+��[*�yޖ�:	T�fA8�Vm�X���=��5�$7�o��\ ��û�M�Hu��R�lTр�1���v�Y��H�;�ƚ���P<�aݞ��~�{/�%��+1�A��t��Q]��e�iśC,�H�����F��n�*��D�09DP��۽�b̊�[s�zx����Q�*g��Ι �qv	HK��Q��s
�m�s��J ����-W�ټ�ί��֍$�v�������=&�>��!�
��{j�^��%�Di�)���~H��F�}��)�����g[�i9r�%Y�6�[t�����і�N���D#�����V���]q��}���:ٸv�4���ewKsԨ=0M�@YH�+�,=̰�cu뿋�w�6�
�Ǒ�0V�+��j,,�F�
٫T�X5��{W���gf����V9���,��'���-�1�t6�C�F	/�ɯG{��O�����wئYK����}^���\+ �2�|}*��,�� ��Ke����\%\O�+� ������c,��ҩ,ǃ�C��y�׊rnو9~�{���#��Wk;<|=���6��6�����!zm��c�+��ڴ�w���-�9{��ba����o����챕���[�c��m{
<}��>ޔ�H�ۯ9ϗ���ˏ/~�wJ%��Q��5��HI�+[�6����� �r^w[� ����xxq���k�Z�݁�fK�h���y���}9)�:�|uvhۉ�@�[���jʆ�M;r� Z�$e��쎭�   Vn�Q�i��9��+a�{m�^�곎Q��B��<�c�~-�^+���D�ռ�[ �n\�Jq^��l�`%ך����_������mQ��#������۫:����,z�\��Ugq��qp�j�)�X$W5��E���ߝ${�~/���3*G,�Cɼ���~�d�J+���~��ubY��r��[.;Wp!�8,���G�"J'�}��˭�7�3��U��n
�6�UidWƂ�e�S������,�M����Q���w�)��W\m�ֳ������`��z#b�В�d"������)�����Rw�YwӬ�����Tq�j��Vأ���;�8�rU�կZ9�h�[�aoWs�c��\)�_H_�|iy͆��?�-@D�����hN���7�eҮ,A���٦����K1ш�w���n&h&dD�-F�3.�ǹ^�J�MBM�æ��&K,h�i��4���o1:ݙ6S"����=����#g qq�����ʜV�P�&[ЯF1����o�}fN��f(�E��k'mf�-�A�3�� U�ɟ����
�mǧ��.�3�\֊�IE����뙱!� t��r�+�������¤��G̃�L׷�U��hr�rqv14�.p��?6�,;9���9o�ԣ�ܖ&ڱ��4�jؚ�q�\�����kՑg��6���Z3�\������������M�(M�*�4+O1�����v�]�~�r̃��l���=QZ�T|�~+�>t��5%��a��k����cZ�l��^N�z���9Gi���pĊ�C�ۨ�YP'�[gi���r|�5��䒟t2�77��}w�̰�5����zVG�'�1���+Qo�]����]�g`�Q)��Du���X��x�n����m�|C/��#��ܴt6kʉ��d�	���q���q�T�����e۔W�c���m'|�t#�a��D>f��7J[A6w�U{��>��+�(.����%�ک����>3\������|���_��҃R�����ꏸ�<��\�k���A��'�n�#9�� ��u_;��Xz:���+3��2+Pv��βO��ݛx��t��na��u\�����+��`�c.��f�n� n�vd�)u�1qV2� � �(j1ơ�w��P=�5(�-���0Bك�K9�x�k7��^٠kM",�a�e�t,c�jBnV@g�rzk�B��laRd�z�䳹5�m-LC����\���Cރ��W�{R�~.2N$������>!2�h��[�!�܅�%��ڹ��sbV����ӎ"�E��oyx]�h�dù�	wL=�����!eq�W�]��0��n�f_^w�p�aC���&�M���Ŷ3uX��^ձ5�N��㐦�D��*a����
sð��m�v!dE�/�����ߊ]�Q^z��E����Pn�^Ôu�C/^xr�a����_����3~�l������,���K��n�]��H�l_�������{�l�W�1݂X��5Q�X�}�xz.�y=�)�^�k]�	��5�1����ok�d�f��ڮ�ng�`/)fM��i9%��D�@3y�^{������z�9*�AKqn'>�o\{�՛7!�vИ�R�� �Wy0���
�3A���r"�u����oa��b��޳�A37�i�.&���(��ِ�,ՙ4>�e3O�g�h�ze������v+��|�}x��9xMtW}=�,����N�@�&y�s޽�=�x����QOMY�ez��x��5��N3H��5��8��VT�G7��u������4�Y�ܦ�
�\��JĬJf�WV��E���9�k��@�ξ�=�'����h�Z��*<a��0�xg�!s4P�Ó��,�zl��bޫ2��5݃X��JY����'z��EU����;r�o?Of��7��@_r���[����*�)�:[�S�2NRV�Z�D�@I_��,����jwܹW7�w��q��g�ɋ��q1���+]*�f�Kܳ|(Ċ\�3����6%��B�Hl�r�?%�{���ո�P�[�²�_8F�>��oԻ͚��q�Y51z�ՠ��|�QM�o! �yVa�
 �tc&�赛��W�}:ě�yq^����"��6�����n���A�-q��vQ'�끼c� m��m9�<��מsB����/�5Ӄ����5�g����3��^׼Un%F��j|H�>�Wd{g�L{VA��=�xyYҮM��.�=���=��6�h	8,��4��z}VF�:�:��I�i��&��^K1�`�S���^97a����Eh�Y�#�|gE[�1a�[z�M�Bl�j�c�'�jRʋ����8cF��ҕ����-����?��m|����,�:���^�]�+d��p�k���y�n����zc�9���D/m.��Ǔ�F���f��v[
j�����h�zz��.o%}Ƈ��k<p��k�Jƹ��yڏN�4����J{�3�������6
W�
���q��"V�����F��r>,�X��)�Œ��J�V r�cb���OE/[6���]Zubh�C��Y�o�3`u"p�W_��N-t(��P��j�f�q������/�b�&�=�F���I���(���~��xo��j�ϯ���;�,7Kw1�C�'}һ:�;f��P5���C|U�s3�[(^���J%�^������\�a�$ �_bSqV��w`w��=�̧��FC1{��Z;]���w����0M�g��R[�nڜ���]���W�UW,B;�~�(/�F�j�!/�RjK9���Ζ;�34��~��{&���K�0e�ys�eY�!������6��5yݙ=9o�a��dS�P�3m�y
�嘚LF����ɦ"�F�^q���s�P��ݺ�(qp�pkA�vB�tcD�]�s�;�U7�k�l�s��m�"уB��z���k�ܮLO�P���;G"\�̬��3SY�<ף�q�@�oFh-){h�\�f����Y�:�4X��� M�vDHM��d'��'��D������~�(���W~�CP�m��c"�Y8N�����Ru�U�Ao��[��E�>}�V%�}�{�	X�M���m'�=����0OZ�������6r{�$TP�Y�(��yX=�pP-D�UU=��]��bc�m��G����X{9�n��y�Rv:*���T.%Ӱ�x.<�q�ፘ�;��]}Z�Q�)侅-	N^�7�Z�9,���M�zYEj�%�u�mݪ���4V�Y}����EG9s�q���q೸uƠ:��LsTlx����1���kӅ��yT*�ia�Ah}+	]�>j� =�yQ�FЪq}�7ד����Ҷ�-�ip�o>6[~|�J�;5owGndc����:���/���U��^r�b9=�M"�=2{:qL��;��ʬ����	�
W(��V&���R�m'ˑ�����
���nz�s�,�j�`GB׬;"[`T�JB�j��YyPz�3�eǄ��Z�M繃ݬg�q��	�Lo]���j{{��a����Z
��ʆN#�oͽ
��e9G>N��τ5?ԋ�nE`�3�/AԬ���E)�U�D��U�?�j����{�q=
�=�)PRw!�TfA��Djz{l�o��)-�r4��}���^%�M+j19�D���:2�����JM�cyH�P�����������B��p�'ŊGN��(w�8�r�����mg��|&���<�<Ϙ�\�e.���]��=��d��sgY�6X��N�����\��/���.������h4�f�3�K�OeOt���{����6wyB2�C]���2�n*.K�i�L}�P�b�iQ|i���V����|��S���M|y���!./,��՗eh��Y����
�v�5x�-��ӥc��F�y-���bꜭ��޳m+�1� ͛K�n3*3M��$]�����ްۻ@dW�r��v�o�$�t���Z�x�W՛�]�S���zg�Z��qGm���+�d'r��l����w`�X7��к�m'|��rз�[����KهTedR�'���æ+�;���B =%�+��Ev��M[Ҹ.������R7{9`�J�$�]���,T���+n�V*�uy`��3ͅ�l}��S���gIHX����+Kkpl1q�i�T�ǃ���w���~�=c\��}b0e����G��O��cݝE>é�G5A��G;��5����]Ճ�0����Py� �R�ݱ�9��N�u�q�)*�]�F��Wq�`ki�$f��Z�;����;)n\̲էOrL�<�N}���[�nQ4{@r��Ż%�4ngP[�=�Fh�}�1�a!݀eL�|�]]%���sl�4t�]a����>��氻�����J�p�9��疃�`U��u_z�w7�<NpC��dB\�E���rC�sԪU2��21��^;�ej�r�Ϭ^:�$u.�Z�
 m^�����d-s2a������dSd�/��>A�Rݣ���~�d{�z���h�m�L���b��9w��/�om;Fp�xh�1[��3�9�`�Մ�)mm<+q��G�o�1����� E�~\ث+[���ɧ1M�0��`\��8mW��x����)�d��ĥ�@Q�x�e��BT\bb�Lݾ4��mp�|7Q��Q�l�Tၴ�f�莑���Q2'H�g9\�t�0�Wc�^R����J�ڳ/��dlI��)���v��|���҇B�X=�;���BPG.m]6�r��������A���_��XĽYC&iwRO��/l�o��#[Z��rM{V�Ν���q ���_=����(z�gHmb�dǘe{3����,ŝ�V�f�r���U����}v�L��ʝ�k����֋��Y;k�X/q��.���D�����?5\7�M�7*���$�r�,��`�٬�&�v�}�!�1�K��<1�E��\��Y`��2�ؘ�.�6��-��C�j�F2��h᧫{Zx�.wH����Ww{�=�.-�ڸ���Is�Q梴�:�!S�0u��<3j�:��p�qrQվ�k��V����Qs��r䆇�}���(si��	}��nç/qj\�T�R�=��xrn	���_���1[f��D����Z̐i�o�����伽M�Ga7�z�ᾰ�g�p�h銷9���8vY<��yQ�K/s$x7�Y'��*6�=˸ϸ�hXն������������y�!��kC[f�J�-��*��-4��r(���Ulb��#Ti�D�VƁ����V�d��g�m��&R�g�V��A�%�%�*���,Z�KD@U�����"�:i�!�E%���\�F�ZMjb���-�LDB�Mi�Y1�F��	��-�܃HPsb*�ZX�""�����F���*���cF��j�qE�5���85c5�[QSU;`��N-�R��M�QSEE[hŪ���1��`����ESkM:UZŶ��LhsEEb �P �  ���ױ%�j�*�)`��x�[�YYo�НG0Ӓd�Q�8T*Y�Yt�Si��v�򒮡�4�j�r�u(�ڴ��|/�}_}_�w��/�A���i	��8��f މl��R⼢X���9f^���eOCfSy��W\K��ig�T1~|����Ղ�u�@����پ�h���,yK���mɤGh����lsfаK�3̩6=Հ<ݰ����Q�̉��˹#<+#z�V��c7zƸ�3}��Z��h���^Gz/O\����w,�8�����G:YYZ�5��U����q~ƙ��gU���~�'w\���׾�W7�J��U�`��'U��VT�)�`Ќ(�MV��tz1nfqD��[t��`Oe�|)B���V$WB�C+l�q[���Q���*�nN�8����'��v6�M\�]`6ߔ��`�[0�G.�x�[5��g���W�T�����}��;JX#`�B�9
�g.'��6:�8��NT����5�\����J}�ݩcdFS�yh��6s_(�)�V�q������ ��a׏�1�h�Z;��[;<���fʹ.�Y�χX|>�����.�f{��a����Q��G�D6k�^�}$�Wp��/���n:�]\��x����%�3����E��P�:�:�<��UW�3�}��;�C1��*M�����t:�\�Εk��9{Ц���6U�QC�Y��"~>�s�4���Ю�:'˟���H��OO^yl>gVx�Ӑٽ�_�h6��Z�"��G�mn8�r������܆�J�˛�76�4Wl���u$4�*z!؂؞�%����=��7GwZ��9�����a�԰�V9m{�ð9T;	��J�x�&( �6uv��Xt�oM��;w��ܺ'�'?%v��K���S��ⵎ�d����>��sq>��V'�����O/iX�S�r,�iN0C*L[��=�=],b�����f�w�:�Y��+�U<��v!�0�j��G!��5E
�AP,����]��i;y�����*������K�v_n�)�#v��F��qW��P��{}o�����v��K<%���N/���t���	����s8d��J�������Ю�C�=�7I}Gc�U�t���pq*T�n�0�����il����8����n���
��8W�\�Qhvop�Mn�D�Ei��X(��]"�ٱ���6��3��YJ������Xw��J#��_/�����5q�7��d�x	�p������ֵ�J�����!�F��_>��uߗ��4�q�%�J/,]	�Œ��
���M��n��3z��[d�uC�uӝYBK�Av
�I�e$�7�|�q������|оmxw�k����+���8��*	.�ق�OBF4bksQ���4���D��}d4�n2b�5a۔i
�۩�\"z���+��k�Y����?i��x��):s�ș�G��vC��Y&%k�bV�\̽/m�oV�TkK��s���,p[��{�B�9GFEr�n�����vJf��q��/�Ϫ��vy\\6�3R�����
f���(Kͣ�Z��U�SOf��ˬr��e�� ����:�����p&��?p��%�hl��<��}��,c��,��:: �3��n'D�Ԕ�g��P�=]KJ�2V��@�T_����$>����-g\*�Q7�ý�����N�?u���s��vj��e�[3�28V�T8�>t�&�i����v�?�\,����5�)4�k1k55>��/�/\�'�����;V+c�xv�-�z(�|���s��_�1�^NTF.qC;���^�Fv�ur�����u�g.V5�̈́�vوkhz��������[�:���U쫖RZ�*E[�ٴ/ĭf5�7�rf��[<�f�z�����ٗ��VwP����:�����׬c�xw� ��վM�(��^�Z݅�71;�Φ�`B�����ڻ��-fvƺ9C��N��
�ҵ�g]���j˴��U�+�+8��ث}�J���`�|Ռ��%��Q�Os��i��@�*{~���M0�we�h����V&������gܹ���NY��+Gu.I>���P{�6�����g!vj
� ��r�)%�����.�'��եz�ه�Ln�����=Ꮧy3�ˠ��2�_Ԏ�u)\����h��g�r"Q��/Ћ�D�r�L��~П�˔TBr�\a��耑���� ��d��>��4u��-�$_���M!1���f��
�*�5˩�3N�Vϼl�}��/�o֝�����;��4
aG�@���iT��2���ʹ8ǻ3���˹��@����.��W��Nia��^r�7�O�0��&J�����?����_y�p�<�j�Q���B;�>�XTKz�4\��n٬�6��˓��urU*C���b}K�r��(��6���|��&j�e���k�����ʲ���ٗ���_��e.^f��9�ڡ{���;+rRqe���/�A��B�i剄z=��6�]��b�b}T}^^��]��7=Qm���/;��O�q����;C���I������ǒq�f�0���C|i;�PŇ�z�������u���rⷤIg�<�N�yVӕX��f�h��lri^0��7۵i����UԬ4���P�^�yn���l�̝V�����1�3�+V�`#���f	w��>�9��[.�}��2�}s���:����BlbW���S��FVm���[����+rS��X�s�o���,ںվ���.qZ�稰��=HЗ]��^�R@a��&����dv�!fv�_/p�8��Hf�[�e�ɘUe��۩*��C~�c7��f^۞�$��
r��L>�3���z�u4�Ӂ]K��f�1R��]CK���(��W�UɆ|ö�z$�r��+�.3ݟ'���(�V%9V$WL:ޤ�F����ܫVs��o_�W>V��Oq�>�m��*��A�]���Ԡ��j�]O3.����Ѱ��e�^�M֢E�F$.�ݚ�u�n���M@����ލK�ݾE�ES�I��!3���F��Ҭ&M�;�>��}Nѝ��4�.���UfCzM솯�-�Q���`�w3ڝ�Vst���TeC���Օ�1�l��㍏�&����j��Vأ)s��3��B���jdd\)�G��\J�Uj4y�[��"���oz�|�i��v����<.�O�V;�!�U��m��g��*�a\�����8h>*�;pP/�&����ԣ�bC�su�=3��!�J��ߒso����uǼ��[�<���kaFv<�{��	���b��.q큛���z�.����K1�*�)���8
�wv�FGo�/7�7L�$�+��~y�.]�0fxC��[i��A'Q.��{�K�~R_�Xp��V���U������G����:.]|us�Uƥ۶s^�崨�`�b�[����?+��wE��2�M�ַ9��x+����r�j{���D������\t�q@��a�-��诘�ݾ�	�&"�$L������^�]�(z�Z�TqC�U.��}IR�0�b���{���Em�|����go�j����k�eCY�(������`+�M�Pw��e�� �ʁ8�'(�j,ao/�mhu���y�*-`���8�f�Q�FΥ�yWS"�?)ޱ��Ε֋{�3��6Y�o`��*z�%��ˑ5�=M�q���2�V+S�(��r�L��ȦN�ӡj󎨚*�4L��	Ŷ�k�O;��Al蔂���m#|�X�OH~�~mve8<m ��'�Ҝ4�}��W�J�P�I�����Me��f��M��L��:����Vo��x��	>����C�v�U �b�Ԗp"�!kq=���O���R��(!�J�s-��0��"�).^ՄQ�Oл}�{}H1P�͌���2�Muuz�j��q��еc4M���$�cn9�f@o����]��`vC�kΎ����c"@L�Ks^����%��B7<p������%�(\����0S�d,�Ke>¸f���,����T��鮡�h�wj����"�FS��v���3����ǹ��]�={j\�5���VxF=pk��)˽����zX��5�����l��h3�U��OGt�������_e�~w���qn� �ߌ�����Ŏj<�kvʸLL�{��3d@�Yc]uq�t\ J,9�L��U��o�}6�]�xb�aw���5�bϨkzrp$�Zr52�ly�P}P��l�|���s���e^c��'+6�k�O�T���sjU�kՎ�N�F46bڣ_'�*�k~��.:|��(z���x?I��Y��Z=��fв^���8j��cK���c4���;�Q�S
�y=Vwx��F=��]�yk]P���U�R��z	�9��-]��\L���bN�v
Y���>��
�t��[��M}�Mzi֡�1�0��/o/Û��3z⒛0z�_5�%^K/��J{=��u��6M� �bP���ǒ�x%:�+&h�̈��k]�o��C�b�Իgў�pQ�ѯ�*��]X0X�c����S+V��y�B�O�2�YZɗkҸ_xC9Y���C}�*vR��En�	YQ�̚j����U};+}�=����k��	.�o��>�R�U��2�K=����]Cc(;8�󾊕��2¢� !����5i�3��=�+��� ��Hv�u2��.���j��5�����m,�0{����n��8�f�H��i�Sښ�ǥq[�Ĝ�ݝF�{Э�9ޅ�aM;S~	ҧv]<Dk��w��潗Y���~�~}�3�]H;��'^=�®o!�A�ބ�n���e�����Z��W�)T%�h��}���O_�{��)tcd����e�a�r�$;�CB]�mm�p�^�ŏ!T�U@�kڪY���+tKisҰ;Sb��&��l�N-�f�c����r�agu�]Ɏwži��Ӊ�{�~녗-��竔EqZbl\)=�����F�a��]ڄ�m��*�-���_����vkk%j��}N�p8rG@]���M����ׁ��Y�A����*��f����J`-v3wY���EQ�l/�M�!��et0a�@Uh�����x�i�u+m�9o�}n��U��O�r��:Jպ�%j�Nck�qN�x~����� y��p*����y͢�o˼������Ճ��3�+	��1�������A���>��|�xt@��P\HS|��z��a�(���=��&H�ҹ�7����dƼ����f� ��[dy+�8��}D/oԺ�m1�-j3H�����/R�;+�3no��>6Ko���w!%'#��E�W��(ll��U}v�=6���9Q�O9��o��aV�	�6�R�eOU����x)ͪ�Ծ��$rg�.��C�����,(t,����^����AV�f���&��[�\(���U�Q����J�{��5Iv�l����h;�����7;�:p�ً����58J�d�lsU��d���U+�|Y�4ٿ%v�y/r3ҡ3��jd_rފ�+ � jW�n���+q�9�\BcʞY�r�5��F���%y凹����Í��پ;�r��OIx�*h�)�O�EvK�.��*5�AN����Ie&�-�)&���Q�M�{McnJ.5�����ګ+��+�&�>^��'�$�������U��6#������m3kە�^��9}���{��x��������/���a�3@g1�ΐ�B�@r�=N���,e�3WA�OF�"ԏ��^�^��(C�e	���s�f5]ƐjΜ[H���%�um`ٟ]\�GS��K.R]��,��_
5�0
��5Z�����8;�c%\�[�+)���1��
׎�.ٞ,��p�9W �������#�s��{����[Zc�쭪&��؃�CK�+룃װYzX!�j>�t٢�4^֨`כA��ҡj��h{&Q��x���~a��[��F�+�2�,u����4�ة�Jm�Uj��\`��x�,�Y:���n_C�N�E������ά��1��Z�b�f�q�ɠp��gt雬	8�D�m��K��'�1�1ύ�n������7{+H�Ģ�-��L�G�vcѫ���p���Qg&F��&yn�X�(s}��Ŭ��q�����o����PVx
8�
iܭ��kܧ;n�4f#7FH�Z������{�t�3Bc�U����ݥ�ּ��B�c��J꼉��V�M���y�U��s����Im�CI[�"�[ʹ��̙ԛ�̚=w���9��1���R̙��&pw$�xu>��
ťB��a�� !�l�V�e
�#��UG泓��ӵa��{z/5=htq��v��F���/WȖTs鲬������ɚ�rs�Q��qZt�v����e��{r�N._1�_3Z'É�|H�ѝ8���MD�J�sK}/�ئ��m��&��ؘ�ֶĵ�f6�`�op���T����X"h#ulN"��Ef��+pl�5��(��˕��ä{s�t6�[�V�,�L��l��͛4��G/'�Ldþ��Z[1V�ɻ+���|�"�����K-���;V+2�K����ɎI��k F�7���4p[�yY���H"b�%�bȢ�O�u��ٶ]�l��mR���k�<;�_p5��%�cɸI�P/J�����T�Z�S�y�#k�.UZ�����C(��7�

p�fV^��ز�[�1б8�:H�Vw%˱���ir��[���X&v^o�,�x-rcl��D{����O-�]l.�Nf��.���\�e0���k��,�:���v�YW��>��r�D���w3M��xlsJ�R��t�sO�����Q|֜�b��y��Ҳ�k���o��xeM�,�x�hm�$�Ul�U��Y#����8sa�������U��[۟k�����hɁ�0���G��έ?9:Z�X�B�?��+��Wt�v�q���rR��������˖EY��6��J̪-Z㺣{&�`�Jh����cm�*+N�4D�$�EUSEDU������IU���gEF�f"������h4�ƋPb��P�PTZ4m�)����(�A��(т��$*&�Jb)"���[X�A5M1l��
b(-M�5EF�i!�m5�V�ִ�f���(63,�LQ2�킪cZ
*i����"f6��[�[E1�h��T��TD��h2�6qQ43QA�m�kj�0AU����T����sQ�DAi��$�[E�s5DQ����j����?� �H����5�����7/��3]xyw;�!��Sз�ڳ��'um'\3��L �;]Y���-�[BF��F͙���� �oN8A�ʊ������"ӗ$OdU���Grmn8�����$S�^I�]۬C��p��;ysʰ;pQx��M3�w7)�7��"�^˓�F��=�]s�n�ʡ���kfq�Rf2]3(�ۇ�;X6�W���m���׵:K1��Pŀ�O1}\qM��|��=�9��#w��Qh\v��q@��s~�,�{��4��nM��	����M��紕�j�P��
3�K���n�����	1;�Tu
g��v�g�E�5���[[�b������>��j��#��,v��R��ǖ�E�^��G�I�{�3�o%}��nf�C��Kak�Us��N��Y�r��i��iҫ|}�rb���A���6q�[�{}�1"Kؔ�X��$��Y�_J{�|\���t�Lp3/�י��^�|�%���/%.�kv��;� �V��
d��k(�u؝�@xV�zяgd�Tf%���D}�Ŗ.��F��GYV��#��'���#~��ƅC�*�9�%������wέY���s'*�2bKtL�]Q�v����
�nmR�/��h��+�`�i!B�K6���bWs�b��{�bM�v�\���no���WE�,l��9Av
��HŌMn{Q���c��.�-�e�Z�i�`�Z�ջK s�P�H�[0pId�ց���2��څ�f{��T��E�ߗ3a�ބ�kB2�ԙV�l@Ka&s_N���U�5��R���Hտ$j���R
�r�W�5j����ʍۋ�w�.��)�V�f?1"�mj{�;��[W7�v��58^$�]z�[I�ebau�JhC�OE�-�}�6m\��O��9}O�zo�V�Y{V�F:zo�n5Ɛ{�q?�A,r��=��{��3���.�7�z��&[5K\�{ʫ\7tv�m��e:���k���?_�ߑG̬I�̖�м��f?�&vc�������kʓc^ܧ����`폂�FEzv��5���Z���I*�|����-lw���&�t�*���c�H�:�#�٨��Ǘ���M��Sd��r,/��@��,�ڰ�d���4��	�����5�v��Fm�渽g{���4���ɺUZqiB���t�V-�]�E�U�ݜΊ[p�)^^�]f(���Q�E�׷l�7�J�Ʊ��1"͡d�f4;\p'�u;9S��'k��F��#�q����,We��c^���K��8��թ�a���++έ����/������K(a�~��c*ɥ�[��2�ld1Ufb�9i�`��f��k5�U ��8+�[�U��%�Q�z59�MSX��.��E��UgQ�\C�J� �h`�"�l�F�&��Y9:K�;õ��ԍ���Gc�m�
���As��!m��d=ĩ��[�T񎤆�:��з��ist�X��x 㥔�wA�<U���w.8R����Q�VR�����_r�L�2��gzݩ�Bg��%��v���������S�����aЙ�Kʹ�����!LNU�W��$�:��Ƞ����2ׅ�+���gâ���.Z)U�1o��M�h�E�-�
ZY��yN�&��m��%��������g,���ZZ�J�X@)�6e��}��j������r�1�7� қeL���$K=��yǹ�ס�������޽"򶔲r�#(.*�;��].����B�ͩY	�b�s��J��a�V�ŏ�m��3b�o�P��?�斖S��+m�L3��;�M89�m��N-��DK���蚩yoMM��W�.1�3�|n�r�m�:\�p�!��z%�ׂ�T��V����g�K�6�J�?;���N7�T1cV��Ղ�v��/4�v과=�t�~�n�ؖ�|;G��V%�SÐ�fп���!,2:�����ҧ~�'?W~AmtV��u�qӊi�7kc���3�'"�)�w$L;G!��
��G���=�V����8��o�'��<�A곌�NL;�m����S�i��{�����	J݃�bo��e��o P��O:��{�q�q��ϔ�:[���G�lrv[�|�O0$�S(�P{���z(h��	V`!������E�zS��}�<��U������J3��W�Q�V���*��8�;V�^ϧ�c{��9ɒ���A�7y�̗�k�yۙ��R������R�۫AVF�N�#�+��7�<J�'�����4.�#b���U$�	�7��[~[��w��5�����cFh�5���4g��Q��d��NYY������,U��j'�_M�i�3��n8;���ʞY2eƧ8�Mg��4Hj�u�$5��*R1c{�Q��V���gfU�Y�m�UY�[��I�q��:f�:t��!/�*f琎�j}/���)�
��w��]�VOm�Ҝ=0��5P�&��Ƞ�3�E�� �3���MwZ"6��J��+ܙx%�x�Nqփc�e>^4��;rQ}w�Z�x1����R��~Kv�y�d<���XI��l��x"�dIo"�9�HYj:���0��(�_03u^>��׮�s���|���9�*�����Dh���Nr��jUף�k~FA�R�����S}���]�Uq��b�0��_
�ɝ{&p�V�p(�������˴�[K���>�쪌�O�[T�ժ�۾Fs�����k���]�Ǫ-������ɯc�[*v�qL��Ek�%wm�,�L�낽,���MqB'�x����s9��
��4�Zg+=XQ%��NkN���EU���/{��|����Ú���l�kr�����t������M4�����*�	�����/�I�_�9ة�v�=�5�+e��1*��0U��o������_�}$����r�4��'.���vz��Ijt��5�<ќ����}����V�%c��a�p�:�:�Vei{����η����]+�o�v�� ����8��D![�wQ��x�7�J`KħX�+��+�J,����y󞐐^������"���VN �!�6)Z�g��B���m#ϔ��:��f��p��Rz�I[�������=�= �,���IOg,Y5��(��i�
z�wi[��8�6��J�:p��\ rقCȇ���f�ʙ��|�mtۚ}}<S&����q�0��j��4R���in`P���z��^-���$p�n�П{�/�r�����&��"����/����4q����E���z�?D��Ow�g���]q�a��������l�b�~��=t�9I���雋{��O��$BO�w�������mMPT�nz��k{�y�?mH�ur��{rnC¾
4��j��f�sW�M٨�h�;W����\�C��l%����ٰ��*:��`׻EWy���a<��i���4Y(�e/T�\w���:3�<���� x�#�	�UI[�㖺����ͩ;����S�n'歕6i��ʋ�W��1`6r����a{��>**�=��L7�N������|���?_�ݕ��6���yl�U���D���ǝ��MD��{Ƶ�:���yS_=0�ʂ�g����"�}��XQ)���>m�+�>o�l�K�1�����|����Q�:$v�7y�|:�S������7W�|�Ğ�����Sj��k���Egh<��[]9���vܳ�p
Y���>�]5���ߙ���7�A��#���[��s9���`*�le�VIW�˺L�{)w
%l�Jfw�h�;m��9+��>�g%�+���!�cyYZM���:����jj��GWC�mi�I��]�*pA�ybf��eu�9:�T���=�sp/w���pl����d�H�X��7��Y��0>6mk��u��=�;�iXja)-��6X�zu�y��B�ҧ�xg���t�bȸ����,���b�Ij㷿���Չ��|��fC�?fv�9���{�Ik�˾7m�;nu��0����ct}|����^���m,�D���徃X�d+��U�,��t�IH�p�WR�3{���ׯ�XT����}j��4K���m)Y�*����cd%p9l��\�#��{����t��XQ��.�v�.;c&5�f���bu��C�z�fXO2d�����YqE�u�1h�@�Rf�0����t,��w�W���؀^��{�T�"7�Rf*������'A��X��A�+/�:�=F��{�N��Ny�+�+er���Xs�m_yHuڃ�fߠ,�f މ1��o����;�jZY�z˒����5o{�D��'��y֮j7����Ļ�6��0n��RŒ_�D�@�ט�f�ߵ>��'�͡~%�
\=.��
|=���^B!9���ܭ��iUAq!G����|�~�����)&kُj��EV�s�����λK��G�3p�:��z�P^�g�C�>�q['h�x��ܚs�|tl��.,�]k�Թ�;��SfZ�'C>exk)U�M@cO��P9�`�N�yu(��;&+�g8�W���o�C^�2����V�J��m�>�P��3Wi��˃��Ã��q�>���~*�������]��F��w^���-��Lt�^K+I�l��6��o�W���9�|)/{!��I�[��-M��)u�Ejh�(���}I�q��g�Y�Ud��ϫ,2<�9<����J:�`�HU��f�^��̢sˡ�@��rY�Z���Bdb2J�rэ�� ��NP��b/�^��I#6V����d1fm�.tZ��|���=�u�/p�U#VTI0�.f�i�T;p��osME<�&y��;�q8�~{�)b�@�j�r�0�������zp2�4Dn:GSN�B�%��Kk'9�s��+f&�9a-�spe��ꇌ�]A��嵺�vY\n��硠�*��]���}7n8�upr��y�i�].��g������TCZ]��B;��f�Zi�;w՜�3�W��8��y�A��C������l��ˮ����Kk�n��1�e���of$��`BD%�ٺ�rQ��vn�+�x�+u�;8tN�It���e�rň;(ֹR��s�e����!A�B�� �I=�Y��ꥲgp:�o�9�@�{��֭uyϬq�W�8��+���Ɍ�p�ᓋzXho"������S=�sȣΊ��|�b�ew�Z���J��s�R����S��k�97l��Kv�.;���o˼��t1���gor��al��'�ֱ��[g����s<�<�.:qB&ӑ1]�{�o�u��G�'�m�
�Ǐ�[&��V�c����-CMT�1D|�E�q����Lͼ�w�j����p�����b���r�5n�O!�	�+lI~�c�ށ�݌�W���[ȷ��5��FfM�gk�,[�z�U�r�*�Hf��JĬ*f�W5c$�(��_�S�q2b#,�L��B'N�XA�c°GB�X�����p�HU��m#n���F��ڽw�fx��������cx�%�.P��W���WTj_�����������"����̼	�N6����{ik8,QT+�|M�q�!��>R�Wfu��QW�ims�Fw�y���*�-t�%�[�-���U ٹJ���E�^͍μ��X��Z�.��;�������l2�5���Bg'�9UY0R��v51�v�u�Ƅ��TGE�iow\[����I�R���+8�)O������.�	�-�hf2M[�7��p.��(�Y�sj��j�h�,
2f�u�84c���GRVxG{2�I-��Pa�4R�Ǳv;�Vq�)�jS.b�::�ʇ2����\t�f�����uf�yy'�e֑��i󴊴3y�j�>�!�_B�����'��=9���Cn�a��[ ��Y\D+xҫ�41¬*LzL���-�dX~��7�_�S换E��@������­Q�J�ٝ�Zh-��![�bӾ�G`�Jw<ܯk�=�^B��}�M���k��F�E�v
_)��7Ȼ��i�D[�Ww��K���~�]��x�4���x�tWr�ǲ�6�)�:ʊn%Z�Y�/AT@|*:'>w�v4� U�x��
�ӑ����y!@�G�5r�2}r|~�c�y(Γ����Z�^���_�\g��d�O"l���X-���9f片�|}(^�Z�7J�ذ�.+M�EE�u+��4p�Η�����`��k��OD�,��>�"����͌^��{�^��i�l+�֎i�z���!މ�*n����m��P��۠��p��I5�6�K�bMe��|�Bb$b�v��u�B�j�r'N����f��)�Ki�m��e�i������5��J�z�������\�m�9�{��u��`�-yړy�.�N�#g>@@��M��}�[�*pg����_fA�#����vʏn%�6��ˑ����b���)�`u��B�WS�We�PB6^(b�;�.�i��{�p���-�N��z� �z����7�1����7s�-*��_� ��wN��y:���n��Y�ϯ���Up;S5G����l
��J�tu3� #O���h���ê�}Z`���:Wkehj�l��ht��3Y�7���REN��Ɏ�d�F�-v]7s���3{`�GG`Kr����t��(�t�>�O]OM�}2�=��gG<�O4�y�4�9���֕%Z��H&�X��(�zx_%WE�T]l\����<�G� �W݇���,����Ξ�)���2b�%���w�o+BO͞O�*�;�^Ѹn��h_P�i��̝+�C�Ys��f�O.f��$��%���kh^� 3.D��%о=��VW���;��
������]���s7�Y]�6��t��J�Q�x�q|����o=�^=��ǘ8�u���:k8����+�����N�֏T�!�[8���;X<}ܗJ����v�.\�i�q�#���l��h��ų)�:���ĝ�Z��:���X����h&*"�h"" �Hj"h��`�TA��%%���VƵ�&�b��U:5�(��4SEDM6�MEF��SETDA�i��"�������0PE0��C-lU8���������e��("��
#X)�*�)���щh)i	�gRTKQUV�;b (��f(��"(
Jh�����f�"����(u�:J�H��t�

&��(i�h"+Z��-e�j���&M&"&��:�(+N��!���j����gE4��C�PRQ4ӣA5�E5j������h�+Z(�)�6ֵMU4T�T�T�htQCAL��SQli��c%U<��î�Y���Kz���|w8��Ώ��w1��7���{z�|�n�MM���R��y��U'?p�n���J[̞����~M'�� Fзic��K� ���m���o�OYz�pލ̷�k'����d��O��ܚ��To�2{z�#�� ӕ#�5u�n�QK�o���'G��&��h%<TL�Y+#ݺ[iv+��q�@�#�$=�q4�kS��8�|6���;��z��G�H<�����X4�E���V�n���g[&���ysU���wO�P^��Um�k �hlg�[*l��Y����������E��W�l-v��|�yݻ��C~Pq�m�#f��	e�{���o�B=��rQKFQ�T���ħ�5�	��N0�� y�Ny�����1�a�g$Vމ�'^a�y8}�k�C}�а^1a����u��7y�N�	���u<q��0���!EC�p��竨�c�i��x�fLΊ�/m֥�o��k/�^AshN��� �3P�pM�X��x!�Co��ó�:�o���7i��nR�d/�K�w��.Of�g�+5����!��w1�J�k5���}�2^��pΘ�¨�.%	��j�wa�D߫b�[X�
[�`�'7c|��~~Br7��M��L�_��}S��7;�	�޼�^q��2���o��w��GsTR�X��`��
ԈYo5qe���g��S�m2]�!U��aq|)_��h]e��3q6b2����3�$���o+����a�����nS��G(�#�)ټ�����:=��>�ͤ38�H��&[ U��.�,%��xp��팍蕧s�u�:�J�dr[#�}��1�����L�R��2B���Z=��j�פ���Wuz�\�]5���ӹ�nY�o�h�\C�{~���29M� 7�d��Q-z>+ޘt��s�]>۝��S��Ǡ�R�u� ��ʧDZ�<X�0xcRFS���@/��mjN<;�U��-�6=�B�Z����i���wrx&zJ�]��z�2�I�ύK}$w��ү`�����rbs�2T_B�ds��;��V.�\nb��S�D��l�\�J��s�_��{'��g�q'�3� h�����I���B��ud�U�Њ8���\Su����Q�K{2}E֭��Dh�5:�ަRէnWDk1P���������^�*r[����0M���-�j��g��R�3b�=[���a�k����O��[��Q��A�@���=� ��xn�h	�++�r:��� �0�}�k̭lW��v�ޝj=L �up����.O�{�\�k�'���e�#��!|��9q.�Oeu����w�����m�EX�ʨ�qP����wN5�ΤGD7v�"��R;A���Eb��'��d��Y�^,t�/{±\���o��ŝP'�^v<��;^�H�s�qW�����o���߆;O���q�~A��q��=��鎏)�p��{�����\{OY���Ǒ�����s�ٹn�
u��+��w�"��{=J��v��t��&}��&R=�2G��<3��#���F�b��y��_HS�I���#���%������*z� ������ɖf���ƪ}�7x��X�tny/Q��|&<tR潬nWP�=�Tm���c�p��1�2��*Ԯ.��T4j/�P��]$|��د�t�u=;L������7@xTs��eK/��<K�2��h.2Z=��CGr������Amzh�Fh��ʈv�5P.� f�Q��M�1̼���k��l���$Mz����p��5Js,5\���7���.�˽�N��w�NY�X�땢�1Y������0U��|zh�؃[R墐�X�+חן|�!<�T�9��+e�7mM�2�
���R�[+tyN�G�>����ݟ�u#������7
g�S 3�{,C�k�.���^^"==����	����v��ζ���J+��t��ԇs.�	p�f���T;9�ϻ�Z;�*9�Nx�{l�*�C�'�_Ldt�>���Z���E���d���i΢}/ε~�~9Q]7Q޼�LM%^�q�<7r<i�\yU����7�}C�s�S�8�W��#�=��W�Uh�}M��'��e�17�r�[��*�a�K����=_��%f��uG��������{��ව��r���J>������&���ӡ�3��|q<����TH�\4�,�˟jW����J#�҇�����9Sf��$���� �n},ft�{>�Or�=���o��.�t0)Ҹ\�׸��o:(�ݾ��[�\��#���=�����K�g���eo���&�c�҄��t�tޞ����mw�P>����S����1p�ƷN.�YG����Ε
�eyz����2�&�x\dϑ��H{$v{6��X���t�{�+G�1E��y��#�>���E$�����e�d���&η8�3;��[K���=���	X��|ש�t��=wI⳷x/
kD�$��~�X��/�����5��)�;v�<���U�౩a&��q=Lggb�ٺ��m�|�-zV�N�ͥp��'���q��+�Թ���V~���[��k�WL\dϙ����}�!�k�����︯nc��uO�㗜�b�q�\����c!�(m��Hܩ����X[���o&X\s^T8�OJ�}C!�D�սBwU�G���^����ëV�|VT���;sL�"�����',ה�0�̮�{�[AY�J�}*�OC#���W#�^�W��x	����Ȋ�<S�����v��½����x��׵���l�r
�9�'���C�s�Pp|%�f�P���y�^��f�/G`��U#�-ß+�x�J��;j�qc�;H��#���q T�E@�Rzl��{e����1;���a���D�=���%��Ac���Kڶs��x���z�@������,�P�ǐ��D���3p/�B�ȉ��}�bi�z�ǋ㻐&�\+��#�w7_3D�mt����D|�V 9��] ��3a���Q���ڦ<����Y�[�M�z���=�{�*:��6o���C�������uļ�u�i�����x=��}��В�g}��^���m�;.�5ȡ�l��_MW��n����K�m���k���,m�[�3In�<UϺN���5cH�����	�i�Eǜ�=d2��ŧ�o.�>�>ᅉ4>���CE\/����|8�~]��E}�j���q�3��35~�����2zcc���Mǻ��w���e�?��}pm����0���N"{;���X�X�t�3^����G�u���ʛ�w�������^�0.܎��yQ�WH��JJ@���;#O�'�.2�K��=���o��\����n�q�5��sWϔo��(r~�����FY�UP�v�����Nxs��y�uG`<�"�,�9��>C�w8������Υ鮆�|��ћ�4��z�:zpaS!����d�O}��&vt��F�
���
C<��z�|�O���P��џr�G�N�����v��W���k�AL�P'���ݛ鎏L��Ϸ���.�Ǹ�;��O#:�q�k�,��YQ-�f�P>��u�U�����<��{3G��s�"��Y�/�ɔ:�����-���t�wu6}c�
Mː[�8�]5���::�����:=���R2��\@�R��ϽL*��ף�Gs�.=�;�r=����������5w���3^�s������ʊ�����L����԰�����CU[���uԑ?|�����<�'�y���F{�@1���Å<z\�Fޭ�ŒA+����3�1��=�.���R�Q��3v�:�w�BOJ&WWV��΋}P���8v���R��gQv�w�-�n�o%�S��lB����Zk"���r
,Uw�pO��_wf��|�=c7��G+#¯��E�uq�y29� '��M
/k��-{��bz/��ӟ]�>�;���,�t.�w�[:
_w_��ȧ�N��]G����)���衝Un���Rj�i�'���
�{2��s���u��}���I�UD4w>����]�����I��O�NT�/߫�1���ϙ܀xeFj��ڞۘP��J��f�
]��]������4�.�"�2;�b�l����K?\���o}�f�ǣ]���:f�MpZ}Eq��Q5�{���Mqty�;���);0�b2��==�Ӡ�z�*���N����gA�>Ӓ;|sTȐ�N���N�D��mrzmq��X,z�woI�4?R+y��by��;��"29S����[߰����;k���X�.U�����Fk�[����3�u�sy5���~X�2V.�*��X��9��T{y����H���c�n��7x}?Vo��G��?�~�'����H]7�Gz���n#:���Gd�M�v;�ϣ���q��[7>��g����m��( ��nmG6o�J�Y��e�{�����sՑ����b�{S=e������1P)�-c]� ƪ��o�r���u6��Nc�J�����(Q��eu��[Br�w��f_�8�&O�HO�f�%�g�	t���*.�r��y�q��۾���7���M��g�>g	�_���k����\�����őٴ��dLf��Hv�[�<�О6b�3�.�"�s�Z�� _����6�/����'���9v�_s�XZ�[Xq��{�t:�A/\nwEu�s,�5b��+�R����EE���	��"��;~9��T���0��޴4_�]\.
��e���,�أ#t���-�<��=˷2stO�֡F�p��yuG)t�O�����D�_S����L(x�G|r4�u��r˶{'���Ӧ�P��\
�\�_D���G����ڇp�o��tϴ�s�O����^e���ȼ��j��i������޸��*�3[+��A�^>ȀX�K���W��NS��@V���M��er�<s#��N�yfc� vЖ���Y�&&)����%��Ud���k��t;�z�(��oس�]�d��8^��#� V��6�%�퉺��^�yղk���l�����NJs��zFb���|Q�m����{�9� �	GO�6;�=�y��8e������� ~讅��9�eA�
��nh��(�uʥ7.��z 6��7)Q��Gx��y��7��#j�n��(ܛ�&.��5�Eb'����1\ԇ��(�.���}x��sT=�}L�f��uFfȾ�Ǟ��Dg�G�L9Q���$q+��M,�%�p�V�z*�˺c�o���t�t�uS���!%= ,'����h��x�r���I�l�=���O3����@M�y��׸����Q��\U�>�ϊvp��V.��`z]�1���czǴ�gD��t�t�`g�������}ݖ���Q5��:c�b�ߤ.���n��Ѷz��f����[�O�*���Vy������xP�Wi�_V��������:���*��9֞�7�3�������Ȟ�x��Q�k�3�p�	��k]]�aň^����
�ySH�YH+�y�h�g��D�_:�ɘ�2+z��)�ɖ�㘼x��W��3��u��'gi��W��e��q
�_�+*Y��)ۚ`=���4���L!�#��8�ܿw����Aq�ن��H��d��9�/M�g_S�Yy2g�����b�����*�d<�;^χqxX�������1�soQ�#�u���r����C<�����ՠ���#���A����Hu/�Å���
�kC�U�P�����v�u����okL�K��!s�-���%�8��J�TF�_���vV��P�:�`��ѹ/6�z;w^��f�7�G��������TU>tq�͌�\+�%��V�5���{1m���Q@p+@!���gJ��$c���×Q�Х��z覐���;VU�����#ٸ0t?\U"bi�w�A-z�
wO�m^ISO�v'�E>~y��1�����	\1]\n�*���}2�S�������0��lP�N�������=�H������� ����`T<κ�W�p1��=D:��I�B���=�/:�ޣ^���EQ�r��0�!uz��������}@S��.��G>����c�*�[�y�y>~�ޠ��	�K35�õ]�?F����&|{�pr3G�����u���{[~������,7�O��"d������;�����oަµ����N��#e뛏wm�>N�*��j�@z�n�	�'�}-�tG�#zX��c���-�����~˷�����V��%޾n�ɻ��*�8.ǟ�������B�o�xZ~5�rH��P��}��yնo�@��#�k�Å��<:%轞�p�g��{Y�k����:C�Vw�S���~|0�g�g֖~J*�+��������\�������]0�L��}]�D{��{辸����w���TW�DSfl V�U�/�uE{�1�j�9vXYe̾<�:r������GP���ٌ}�L��ڋ�Y�0����fޢ`@b=�R�B�^�n��8�����V���lV��{��ybey��:����SX�Y��Q����o-{�Û4θl�2�k�q�ه�1��*�����ȝ<����aE����7w	�΍������Vc4ɶ'�ؾ�[�)�h#+1�j�p�m�]�t���C��k3z�R��
�ԥ0�����x�]3�^n�$�ea�mcչ�]������t�Z]m[�M��	��a{�Jv�./]m�b*��{��^��r�:�	�vY]��39�Z���-�����+��p�Va*6'Hw_�e�b��拘�=��1ְ����Z�@޻�Y֨��y�ZKgj W5�ig�R�vݲ����ݠ�Ȕ>�Gn��Է�Q�yԀ�B�e�q��}7�)����L��nf�<ك3lR�Q��&��*��s���{��弌�D*�]�I��YK:��!��6�1rI�.��$�wq����Qw�6�7��w*��FXDE�T�q�-�9'm@*�gfd!�n<ym�U��������=�5���9��/i�.�w+*wR�Ο4�;e�WT����Z��/�m"����ms�Hi��$>��x��&\ݾ���l:�ӥz�7@m1{)mZ`m�yE�A�����,�`�*����l�8J�XU�Ɇ�'��z�m�;�1!`��Suw��;|R�Vm��S\�����_{٦�&qy=�6=�"���Vz	��iJ4� ���3���(�;O�@��Y�!�r\$�L�[۽�RU�]�0d�`��~,s|�C��2�;��	�+7%���� �ûSq9#�ٛO6�$
S�UҒ�>(�i]�Z�Q��¸��o�vxFi��:�A�L��Aŗ[���������x-�;���0��iѽ�y��7����#J�*Ws�b�0%�M.\�C�����R;���E/:g��Yb���㼪:\M��fW�.w*+ksSB��>k0A`��t�.̣w3�=e��>: �%���.�,h���\�lJ>�K
☭g-���on�G��.��`�zl�_��[�U��ܥ��_|��j�;�,�h�z���Wt�B�u��[SaU��M,�/X7�^-����`�	uyR͜_^�L�[A�b��b��B��L킵�F���u��;�_U����l��$R6�5����26P*�˶{l5v%u\��U��W"-������<��R%�j�/�J�ey������v;N_f�[����u���a�y���plz�GZ�)_}3hs��1<Rk�(k]j���B����SUv��3s�T�;�8U���jإ���S,b�LU��@�z:Goe4���DZ첷Pz��xU�M�|¨z<�8-�z�n���|��pna��1#=bEyx����z��mq{(֗뿿���w��\NER�IT�US�QDKT������LIE0LQ`�Jf�"h"��5N�18�QS�CDQUQTUQQPTƓS�4�QCj*)6ɣVƌcT��*
���
���b��C���
��)�(�*�)����-.+�PP�(gAl��TQP�QF�5UD�:�S0Q8����)����i��Z�����h��� �6sQAA6�T��STPU�j��)��f
��"6C���]��D�A&�5I΂�m@�AN�,D@�-��$�Ʈ`֐(M#IE%%�%-rDF�A@�tӣEI��G��g��p̪8�v����0M�R=��5cr+6z����@Dp�GX2C}}�2.�7%2� 8:+����1,�v#�uʇ�J/���^�Jb�g�Nk��K����|R=}#J��W��TYW�`Z*k�]�ʫ����9׫��k�*�	��"�y.#&P��Ah��z:�NGt���W�u�@֛T}b�W`�+՚7WӦ/��{��s�Q2��Ԯ.�=L*��^����:϶[�W��<��9a��ŭ���w��dX�!���D��T�*WR�G�G���,y�ɋCq�z����������_Gm��__[��\nG��spH	�n�Т��A-xy�|��$�ѐ�=]�f�.T�wN��#���ѝ�@y.H��<X��IQ\�WU��=�ꞎ��s�|
G�9��Lv�r��tϙ�9����z�����S��jL���
O�Χ�i�ʤv{Q��n��/�G�ޮ��ڬ\;���s�{��rE@�= :�u�"�9;��������Ab��?&]���s�ck�SQ���.#]�|�M�u����ٙ�NC�P�%��<��@J�K�GN�vle{�z{�~ޝ},�__	�,] ߿_�E�ةm&��5�rj��wi��C]hmPԶ��JWKOmҚ�_.�bN�����-]vK6�RV�x����%��qpASڻPm�Bd��{&n��^�-x��u�njc)����哭��v�e1Bx��%5w�wI.���t�����H�C�rt���}P��nW���Xw���AM�{����eb���{]@ͷ`\oO�����N�����v��$��OP�|X�FW����*�ZKc��3��P�.�7�
����ע;�7��v�;ߨ��ӓ��k@M�=����l��As���ɟt��HNt��evp9���4-���p�9z�".��������]G���?@7����U�`M���q3�o&y��!Tx�3�#��#���|�@�d���^�;י�J�Ss�u�j��+{L۩�\��:����n2e��O4�<;:����>C�͚���}�*P�AX]���*��}5i��Ԯ.�0Ѭ�9A���+��� �ܯc�XS�̪�q���<;�����,���-��L�;g ����7�':����U��B=f��s}RwzB���0�RF�����g��'ò��y̹=xd��-�W���{�v锻L�[[�9����sǸ�ݨw���GL�IGI�ｗ"��9 8K���S����&ޝ��6�%ڹV�ӳ�$�{���>�Y���J��p��p��	A���u��nc`ӥ�jR=yONS2���X��s �黚��#͌�c
�EG&��&cږ�b�s{��1*��8��vX�,�p�YT@�v���i�ٳ�W�G�xw��D�9�|2J��|�_-]lq�u3��/�o���4���m�/ї�ot{َW���{lF�\}su����5>����%��Ud�m�_��z�֘9��v;֎�}�x%=��:�G. N�i�U��D�C�O���έ�_x����}zZ�Y]�3���+�'�w5w(��%_Τ>,�PIGO�|gx�{����]C��옘�`�G�u��D��k=ٗ�#]Q�/���=�8;Yʛ7��g�����q~�]��S��:pǻ��&�ǺFr�W����Kb-_dsfs�iW#��늸�G>���3~
{����rk<7����l�����������o�,Tby�WgN��;�����`�*�Aus�nΒ��c4c�9x�ӓ�0�eSY5���dϸ��1�ڡ���`	�^�3��uW�
ܥ��{�"��[�c}�֙��xKf�z_�YU��]1q�>g	����m�ޝ�;��S]Y.��ҷe#���]����Ǵ)�é���MF[��L�����<�wJ���S�:o���8�skq٦�ʒ�7�gnk����e�Y�̮�#�S:+&����#���~��7ٵ(s�vg���^I\��-���G���o�W\:��Y��`��8��t���9iޕ�MƳ��J�A㔬�o,��ʡq�!���	)w�J�J㻝��4��*K>q�`[�(0�r�w�Wjt�{��WB�w����������A�q�����"��>�Q�/M�Y��>S�Yy����׾O�Y�ʎ�,������ˢ�F,
(4y�XU����l��.=w���C��6_�C�\�g������A����UHU2��9������;u[���E�Y3�U�{y���%�>>��̉���3�ق���&2)�w�ק��,r;���`;>z���sM��<��,<VR�.��;�Q�����T�ș���{^�x�;�rO�gwcsu�=��i,�=�L\Cٮ7���ovX�@�ʫ��}p1��Q��R�� ��{=ڐǲy���n4��b���4{���y�V�g�}�+��dM���^�s��GwFs_�r����[�Kמ``�=��[����8�3}�^��Ѯ�Mѡ%1%����]y���4��S��N�g�팟
���ϥ��u��ݐ29S��P֍�C�~���K��Lf��J��	�f�����)��t��e ���mp�Or�V�u�O6���W�ەF���}w����DvkB�!�i��{_c�7��t9|y�U��as�௥��l<ϯo�!\�R��{o��]�+���7�^~���b� ��ӊ'�.2�K�8}� {�i�7��*㇟�BT]�k���G�U�h�:�<�������5�rzF,�����P�3�l��1�f��y����ggH�]����ug�|��W��ћ�4�u˓�����[r�oڳpFj�\-H}�s�Zٲ�zz<T�q2ǚ��*=�O�*�Ң;��F�(�����jkj�ѧH�3��+���s�Q�Z�7	]1���q��4�=�c�_���y�X�=�z�|���mNzs֢�.�J��(�N��}U`LT�e���L���|&����:W��mr7c}�)n|��͵��F���U;U����N��T���l�V�qu�a(���8\.�ltq����{��׬za�7���w�0��y�����P��TJ�X@h���CO�k2��^O�Vp�[Ӟuj�˾�����v�/#�ﳲF}��G_�dr��@o�(��/k��Μ�q��1�]w�w\��p�\{va뭾�;'AJ;��y�dSʧD\.�ŋ?Z��������{��%����u{PU��p��(-vt��wn<֑y�o;�~K��S�\���S�l�cI�M�;�?��Ï�6D�G�/KF��/R�bF�n�D[-֨#�ڔ�ޛ���xgm��m:�܂=]�=�/@ry�(�PZ��k�u->h�7�����R/V�S�r����da���0�=���Q��]��L�=%���q�
}td����;�\c����C���56=ю����xȨ�O����ڬT6�Los��r\�^�¶0gL�x�S�T�>�e,��weIVznZ:nc��^�w�O�Q�>o��l)�X�t:������EL:=)f{J�o��{V7��`#b	XOG�;Q޸���;��Wi�ޝk���ج����maB�=�̭ڮC��E�ӓ��T$R�4��܄�9s���>�xo;jzg����PL\���R�3=�nT�[�`t'9�v��{2�7�5�wv�Ez&pg�ϥ����l�o�� ���x����_'[gÀΝ�O@�Df��:�;]��s�q]�GN�~�������DL��%׷:T�u���R���댙�t����3���_q��qZ}��k���4ڈ��T�'���n.�(�C��:�D�W�YU`Y�,{&|��d�"�fB��g��ι�ܟq>�0��(�J�
-�OG�ǗeO��L�:�e�́�S��Q})��&X_��!럹t?�9X���)�7�E� �I�AI���x[�(�pĝ���P�YӄN���[�M��V�<F��g.�39���uT��%��|˷lU����A:�#~����2Wsd�t	T�p͑q�{�����R����~к1�Φ�1Ƒ�55Χvv�E���Ә��z�3=�s�+N�wX�PcJ��7>��7�XL���n��R����wZ�hE<�ʤ�5>�X�(��m�(e"�~�w�������d�,��-��t��b�FZ�G�^���$+���\�.����r��gިh�׻P�u�q��S9�𯯭܋��]E猀�@���Y��=���}�����Tȓ��/ �dz_��\<�J�����o�����\��V*c�Y�{j5MI]}��3�H�;��0P~��dO��x�d���X��.�;"z���}Ӕ�g�A��܊��&}V}��+����6̹ z	�w"n���+���j�F��ӹ ���xK��yx_z.�ޓ>��حzF_/�t'e���w T.Λ`��r;���^�yղ|�V��kӚwޭ٣1���e,�l3�(Z�>��΀��{�C�P�J>���C�`������}9Pj�o�Ŏ�7�����vQ�y5�L�Cy��5;��j�=�GuV�jM@�6z@�'$J~�F�w����t3�v����7��vMƖھ������<��o�qO����T�譵�+��~q�U՝�A4�=L�rX��\�>�z�Z�k`B�Q����f�i��k{����E�ˁ|���Ȼ�e���F�z6������2�:�<�v/��Y�U� kS�W����b��)x����6�{���1��Y��>����Α��[ɷOH�+HL�&<�ڙ�Ǵ�$�.��%,~*������y���y�����`��g1��׮�g�Mz۝x<n�Y^f�=�0�2����b�g�|��jGz�m�5�U����A����Ip[w��iO�����<��0JG�'��+���5�+�/��8OǊ�Q|�k������"EtC:��}����8o`�6��ص$Xnv&�@���5����{�����Κ��jW�y��yP�4����\R�e�B�Z�0��gs���9���Uy�����^��n;�@bU��O��d4}ޘN5�F�Tx�}��K��
�,���Ϧ��vdUo�K�SJ�N���=���Y�T��U�TE��g��{>~o�����v�����;Y^�� &T[j~EL3�M��Ǥ�C�pth��H����	��6<6��Uy���t&b|�V/ݱ�=�O��#��]���5
��F��a���{�����%��G���/y��;�ҽӧ���g���gu�q�̉n���T�ș���S��h�u9y�^� %2C9�;���\��_�7Qr*��O�'� zJ����]Mڈ��p2��a�J� �9q�ͩ|��a{aS���s{b��|�>��z���w3��[���}����;�������.���y8���+T\;?:>Pcl�۽��g)�#��ܢ� +�e�P�.�G��4��\(�x���9�g�q�cx��>��;���i�T&�_Y���ҾuU�����IU�\��W���}U�����-��������'��zX��|}�2��k˹��t�wU1��3�Dxْ��:��{WON���I�r\��;_��'�=d�W����f�L	�+��ݐ6az`� d��w1Q� �:q�jr|�hOF��|a��ߧ�#�T<�����zk�́��L	���zj���f��ʶ�;}T@�oր�U���]p�Q���/��5�rzF,��xj2�P�h��f͡��z��V���W�uG���T�=x����:�;^�����yhh���.�E�ϧ���NQc2�ɭ{��֮�{�:�#q��.7�,zᮾ���K�����*�<����+<�k�3�:���m�����)���k�h>��:��;	Nb���i:�W���q|^���%^�����aNQ�jbk���z�N(4��	G����'Q<��(u�W��po�GV���z崏�����y�ͧ�����\�0���:�{0�y�\���4�摄VV!������V̜�$9�CDwv�iY�m��Mf��qN}	
�ʽ�WҺ���7`5���5��!Q\!�9��q���{�2��;3��u����,�PT���vn:] �*�eD�d
�ԮsY���W������{�=!�ʶ�D��w�@���c㛎����Ĩ�U!
�WRÐKG�Bgg�wh�*{\�ƭ�w��-S��w��v�����.#��ø��n	_����ͱ47���&�b�L���� 4s8Ls+va릳��B��� =���e���<*f�����6�X��q�.�DV�����gЗ
�|�����zN:� ���\r�V��"��3n���{$vU��M�_��GT\��>��؏+���b��X�:RY�f0E�s��b�P�s���7@R��D�zQ���+�/��s�f�Lu}���7њ_N�{(�*�IH�ԍ���n��|dgh~����7=<���Gz�+�0�=]��ޝn����4oi������HV^[	̖Gz_����b���}ˍN�d�3�T<7�v�2���м$K�3�z�*�b�?QA�������	u{���LJ=��C��Ƽ9�>؞�3�~�غ�#߯���2��+V��!��`F���gO-�F�]�}�8%7�/x�u�YF�	��{�	�9�Gǜ%��6��n�4=�[�MI]h�r��5���+���=\+�Љ^E��0��B�dYl_]$9�fv!��,N�j���Î���Z?]��R�(t�HW`DEvm������v=��xL/Oi�+�����T�U5OE��8�e��K�nLⷎ�z��BG-�G�y�N�[.����s�C0�Ë���Ir�̢�*�w`�:�a�F��h�"��m�U�At�Ny�*:{���JT
{�?,�u�E�O���+�J���_4m���B��Hu��|H�9ʢ��q�&q+1��4��N؀�ܴw'��x��� ���e]_W*|%b�Q�t[��rh׼qL����4�w���k]*�i���{;@,kzqq�ip�`7HmY���'wo���̺!D�����woMڬ��m��׷�Z������-�H;���	����b��
-�+�w�\�5_R�ǚ�Q��a��j��=z,�h�j�������XZ\ 2ϗP�eM��n&�>(vnP���B'o\ZN�F�\r˜F��<=�$����z`�݂ȭ|��˵Ը����­�	��\�����,��7�0��v����:w��D����9G�ѻ�h�ˬ�o����k��n+���G���s]@I��V�Z(�}��7/�)����	{�nB��Lc��yh��a-�V���S��Q��b���:�u�YSҵᇥ�Ж�{2��WK��=�z��F�$��0�_��Pr
�����ܙq�n��@&�"����1�]6���dcy�+h=�����6hf�X�JA��t޺8,`/�W�Ǹ�՘��e�#ɧ�M�\�j�U#��s4'�t�{�����'���TeЃ��/B1їY�U�`�S.o.��$'�3��;n�n�^���&��㙔Q�mX�m�|�75�B�V�LkK�v�_}���_fr��e3���`�N�<%��t5%1q5�RQ�����fGOH�0���;S˕��C^�֎���6I�n}�$"���N��#��H�i�^�c]x�G��J��2�)�n�R�z#Kv1-�yÉ��XN���8f,��^�t{���s��<��璋[�Q�|�7v}Ɍ<�L���Gz�U�����=�Y����0#b�bP�ta�z��2�Wʘ�(����V���lIDԻr���S����e���:��9����J3[y]3��ksA�L���0Ќj�4���2�Ҍ��UX%��`P�D����#)D�F�J_:je��y��p^3R�n�>�R�ʳW5�g���1�]�c'U��	z�7tK���+�~�~�:������+�� j���IC0R�AJV�4iMD%W�T�JrGH�͒��M4��A�i����9�W6c	DIKM!C��)]6�:])�4QCE4��3i�%6�l$JRU RU\ƚ(CmA��CSM<�QM4�-h�Q\�U-:4��%%4��KECC\�O9����r�f
b5H�()�Z"h��G.A���)*�@mcX���(b����!����H���s����SM1D���l)AM�(im�U%#Z9�[S��41RU��(Q�@�HU� 9&�����Ak%<�E͡(f��a�4�U4P�E	�9�﮾o���7}���p��d+���,�|pt�b�Yhq�����q8n�5a���w��s�n,�k4��jV����L���3�F׮:�%+��Ǡ{�ƞ���`R�w�*�T$Zj�n;^�\�%}���5�Ad�V�+��=�����Up��~ɟt���Nn#L���]��S���}�����a�j�ff1�W9Y��F���^�Ǽp��y8���	��,_�3�o&y��!W��<7�l6gy�S�6m_��Cܮ��x�#}��7��1�;�.�Ϥ�.n�@��D
��L�L��H�"�!Qٙz+��&t�����D�����:�A���.�s��\ۙ`=Ț��4� �Ws��ܮ�6�rݗY�ʮ�j�]�'I��x-��<+���aU�L�|nk�XҽdE�x���7b�k�hJU��7�����'x��0ѯza�u֑|J:ˏtO�_[�����y�P�Q���זf|�9�*����$t����2#�����=������%��q�Wd*�@����L)���� RQ-�0t?_�H��;�� ��@b�	u��ԯ�;���__r=rzz�������÷��_y]p
�{"m�� z	h驇���bi��Y��n���������;�6ΐC�w�k���~�U�T�'Ԧ������$��!L���jliK��ڥ}�O���x��]v��I}��B�BM��H�YF���`�c/z頮o˵�
RN���7&Y����8��3wsx]��lW��z{��DG8�޾�RB@��k+��,��f�g~d���{�q�Kv9Ϥ�\U��:m�U��D�C��W�a�ul�A� ��Y����85�9��������b��Tx�C�@rfdg�Ϩ
]Q�����=��Ƌ�0T�{պ�j̞���V�=�ϦCy��"5�"�i��}�w���,��{�3ҩs�>�p���9�U��vxe�c�d��7��l�ėoW\v|��.#��t�Go�qT�����ё��R�O�Nx�v��^��%R��r�������Ν���'p�_O�|���Ւ�����E�M��U��|c�OƷND�>YLeFMx�q�>�q� y�mH�g,;�K*��:�5슿x�tq�� �ݦ����u��oz���
l���Ĭ���X��h�����θM���Ϳ�ߔ�����=З_x���\���P��Qϻ�PV��9�u8�1`{jI��E��~��WQ~���H�L����kj]�������v�/�J�\�,��_�G�Ve��B�Νg���Rw��K�M����;��#�C�<wOi~=7�ƿz-�~�ͬ�j�k*JL�GJ�su�&�h3ox�<k�����O-^&F�:�K+eC&}�m~��ُz%�v#K��v�Z%�U�H�*�GJ�V0t|���=�b�ʌZ��V�u����iv��������{�r��Ζ����w�fPn�N;.���]�`�=H�ч�����2#���U#*]0*.X�{ń�ٷ���l��{Fޣ�Ǟ\
��N��iS�崠�sk*7�ʓ��	h���R}2��8\�9���gC���^�W��^a�:�K�i����#���fD���9�Yby����Ok�s�Z>�{4��8# �`���(Z����ЇDKUro槁]ư�P@��*|�79) =��?^5/�ey�R�2�l�?��-~�����³�F����㇝ې]`\>��g]p��-��@s��u�]���"�!��F�Z�I�����U��q�vN��P�Ùc�O�;nz��uq�OF���R5�&�T��M�3��W���3��3*<X�Y�\����M�*�U��z�AƲ�����.�6{�,�+��?��N����'�=��p�<��3Q�`L%}����?�~�̭^��rs�t�nT�wz�U�*8b����`^�=�"���I�_����X�S�̭�u֦2Sΐ6��Ͻ|G*�ێܾ.=�5�k�kt�OH��Uf���Q��S����T���\c �u�Jǡ;}�F�fX��Ӂ���<�|3��b��E�w\�_&�)bw�8V�|�A�~�R��2��1-��o��泶��r�=�KJ�V&����v�3��nL�\�m�,�{���������T8{>��b��.�V�Q<�л6�q�Ǯz��R�jNL��8��]�`����*���&}�q��&ofX�]]�}���uFx��;ё�/QEg�=&��W����j ��ף��Fl }�X��\u�L�1q�<�u�}�;�>�8�+N_Oq���[~��sX�ONcI����z�*�`[9��U�MN�*�b�&P��ʸ;�->�9|7��؜��TVHy���:����W��eK1�q.��:] �"�FTL�@�WY,mk�J<.���OE�-�+u#�xw;��)��>����Y�p�#�Csq��$ WJ�M��!P��a�N�����;(�ЪT]n��#��@��dx_S��7"<ds��@O�9c����㜋O�z�@W;g��>�|&�0�m�=��VB�� w�py�S�=b�2�M��{d��m�lq��9I�|}����#f_��3�j��9���s�^�[����P�3~��S���}�D��!i�R�tgQW+�Eyϸ�|Z�\;��71��q�UuTb�2(��#��-� K|C'��y�ve�O����*Mb_4������n�v���2�����Y�s.��]v���ܜւ��Y���jsż�yg�L������To)N(uֱP�:�e�X��fk*d�����[yRlޓ��>�x�Ȯ�{�'����;®�,����<��Yj
�����������S�9
�2��*�M�!b��?-lx���0?c�_�6����r�W��%�K	�ڄ��<�kǰ?QW %a���Grv��y^�g����Uy���;#����3ʸ>��c#]Q�;e���uP�P�!|��8zB9��Cõyȟa��x�WX6�=��^7����F� &-{����F>�+��g�~��gFfå���t\̣���W����=��^W�6�y\�x����=��D,u�v��7J��;ъ����x��qj����қ�r�HZ\��+j��FMx�ɟtǙ	��#�mvp7�ţ�&��gf=��VT�y�خ�=���(���l�W�YU`M��c	�6Oin6d-�o��\+�5��b���x���6w��\��U�*xƾتf�N2�*�	���@�)����<�ye_z�\<ް�k�	���2:#����:�ت7�����#�Y:{5T]�W���y���"�d"��x��=Y�h��ިv���C�=�s��#»���W2�C�[���먝͋� ��+��`�{�iAN�@zp'&ͭ��8U%��#�����ʱ�2�ՙ������8�H�h<<m�k��+^OXԋl�΋��CL+X�b
J��Ti1�{mT�L��'����������=�:���śͤ�;9�����XR_D�l�h��=Pѫݨw��>=:�g��pLC���J����yڼ�������&�L��D㞈��1�i�,7��Ƣ/v����T��Q�˄*q:����%�J�yD��9�7�"��) _��O2  ��H��;�� ��`,e|�Z���:�����Đ���ILw�u�]3�����}Vd�q�[:jaﲸ�����Q���xn�e�V^��W�;cR�ݵd𿵺�9�t9NC��:��������Y���X�����{�,*!���b�3��}gT��ei�Ͷ4\*£]Q�k���U��>���Iҽ��l6s!��N	�>��ȝ��Fi�[�y�zn4�&k�T>5�_�Tx���bt�L��g*l�U�/WE�&�q�aW����:��0xL�H~�y֍/���X��a�ٛ�0+5vGo��q�΋3��۶(�m`��ū�V���|nu2V����2,~*����_��>�!����2�҃j�<9�������@��Q��)�uN��b�����1p�ƷNOH��LeFMx�y3�7r��˚71�<���)��A��X �D,:{�IK�{��M��|��,�.Vkn� xf���v�x���+�E��[5�*� ����I��ƸJ��V��.�<5�����*���UY9Os�j��I�%�Z{0*����گ�"Qf���5�W��Uv�����lZ�i��t���H{ݕ:a�	H����YU��]1:=��u>iU��Ǫx���z6e���Ԏmu��}�\����+�Whxw`�5=��m��nGʩ7�X�^C�-sЀ�^ۅa��	aq�ৰ�v�◣��)c~������;B�b38}��_�ʔ�����l���Q�&�\
����zh4g{j3�\C��;�>{=���v�F�� e� ���Sxt�{Es���9�*@~کR�W,r=��aU�x;o�����6�-���ީ8���<7��}'ƣ��뇑�+���|%�f
�R+����q̏O>������ћ^V�e\�ik'�o}T���(�}�>)��$u˚���������/p���'5� �,��
����.�(u}Ӻx9٦t�W�#���]ď[�7�E4w>��=ݗ]��H�^~�s%���R�Wrţ�+���>���|3���=@N�*@_we����)�^]C=V�r�F߅���O���m1���ck����~��6n;�ȹ���7q������<�e27���P�'�V-�(�����o,*��~�%yˣ�8Z��W@@k�밯oy4xV�Z�3����"��bK�Dr��gT��wĺ�К�Z�� ��r�[V��/s{����pn����?9�%�;��,g����'�f�,x�׋Z�2�U=1x��^)���h��L㓱����^p��6�����*�����	�֢�����z�~���G��qF�u��xN�[�)��Ut!�s�,��r�*o�w���>�ό\rw��	�=�%����y�G;ו���|�Q�y7��W���) ��8� ��x�;���r�};w�Gvz�6���,��UC�:�ǎ�
�44���w}R�=�Нm�q;~ڑ�����X�;f��q�-��H?d�}/a!�s�q���|�ҧ�y��?{�~ч�g������괳�@L�ٖ<���*7����]Fq���<�y3���˲|��2����c�W%�E�hp+~��&���L�1d�.�fC_iu�9�/�Dyj{qT-����UAD�eװo���"��yV+�dB~���������UXS����E�%�*��@G���_tt�ཝ������[��Oi�}Q�%e�0�%t�9�/&[ W֥qtB5*<�w����=�:�����蕧r=����:���P�nv	��R���C���E�Or�����o��ĶI�`�,m
#�ޫ�Żs}x ���'*�Yx7=@�!���</�]���k�f]�=J��rW�����{.tg3$�a��dS��^�C&��;���A�[��x6��cr�G]M~ eM�d�QH䮳�#n�c\�r���m���~K��ߎ�<.>uԑ������__�t�wdr�s9�Ccp���B�E�;8nz)M
��Ä��ba��T;�[}�vN��w_�:�UWxFĪ�.�c��=^��fyQtQB�_5DLS���@/��@v}	.7�����Iup ӻ[ޞ�h/p��`T[~�$\)��R��3�����"���v�V.Oޑ;0�"�ݓ����G�0���"zr1R.��*�D��;��ו�q��d�yρ��w:�`�����=b��Y</yYy��]4C� �}�	XO�[Q��6��:���}���;�y%A<����83Q�`	�J���uG���rw�dH�.�Hr齞�����0{r���XeSƖ{�0�n�B���W�������[�.���ԭ�G>�̩��Dm�	�J=���)��k�ܷ
�Y���Y+\WP�ٟa@3^.yH���n�t�ŏq�{������7n+�?Y�ݒF����;2�8ɯy3��'7�Gz�~���2��O�G�`+ ~�aM��iN<�>D@MD1�!������^�e3y`=��R�(f�>�w�©;99C7u�
�}BZ��ǤTjǖ�Ȓ�|���}|[w��e˫�b���K��*x������A�)Ĥ2�<L�3���J����\�cQW�h�O�y>�q���o\�)�|Kg"%��
Ϫ�	�����w��]8�����m�^ѥ쎤���	�)��s��;+�ګW}�xƨ튦m��.r*�	��D
̿`���h����݁x,μ8J}��q���3��=�s��m��A����lwEu�s,��W�kJdp��*�7�/��@Ĥ�R��dG�7�چ�t�Ϗ�\7}�P&!���6�Q�>r�=U�j�u��oxҮr��5Sѳ,��FFԁ���qꆍ��=�]i}%�G�'�}E7}�fZ���V����Ǌkz@��[%\x���:Ϯ*dIs�{ax�}�|j�j¦���u}��pG};)O�����C7��RG��S�����D�~[���v���u�Ӵ-O�ĉ۽�z�f�����}1��)��uO�+�޸��5�@�BZ;�u��eq11MW������5�Ȫ�̽ήbv2�B��5w�4ǽ�D���k���������:����i�sU�VNT?Y�j��ywb^��{+��ʌ>�*Rj<W����	Q�=��΀����,䀗D�}���l~E���pG+�{{��Or�5�*+����:�#V��Ɔ�s��RI��W�Qk��P�n��h�V�:��&���d�S����x�v�3����7hl�p���<�P-��S��Wq���* t�5�mr��t��M��ph��9h��KSW?�RH�$�w����]Y��\�m�V�|D�{6�/�����~�z*��A��i\[gTkη{�)oq@X聥2�ҺNa��<!b���ͧ���˫	6P���V��m{���l�gg��⾞yR�kY��"+ǷJ^�:Vq5w�_h�.��T��8Ec6�BE\+�p¨\�u| %�cek�ʇ�"	2��\�]���^^ŝ���i���ֺ]�q��c-od匔��{�(Ԩ�!띟-�Wr�L�x˾^��W��*��u9��`R�-�q�p�W)��ZI^�`��kŘx���M٪��nd�	����"����`V[����J"�ar���Y�w	��r�r�71��'+s��%l�T��:�K���C�j(k�U�.���UhS����_>��	(�^��h�fu��[T�Cm[c�{�?@��ہZGU;%�X�`��E�qF�8�nn��3s�;ժYQp�	�|B]�L�b��[�����-�:�������$�e�(MY�dP��s�����v)8�r�McD�J���;*Іf�ƴ�1& Z��{�S��y���T��3tv/���zm9�.oד�J�1[��U}�!ǣN4�W�{�/�Ǧ*<Hn��S�<��YYfiE��;�O1������7�����s*0f�\a��<	�%�3��/����]�ų��
clec�g.}��Z��
�J�6Z���qާ#�jQ<�L;�N�V}�O8G��4����Ӯ�S٫F*W;� �AG+�~>�l
�G��;�-[�����S��}�F�1���A���������m�/B������G�C�g�	%� �[�6���(�F�dձ�Ӏ�b�ꖄ�W%"L����GZp ���:9/6	/Q[N��1:$����+s��T4޿�k���K�z�!J�o�<Fx܆|"�岨�'�j�^��9ί7A�Ǚ��7Q�2FU���m3D՗n��m�]��s{w�S.	7\�CݙA�a��h������Ց��pL�qH�[2�{x����5,iT��Q���wf��Eо�j9�� �5S q�%��z1�����)�c�9�po��]��氁8�"�rz{����nдk�u�~�{Rٴ$Zݨ���"��sҬdȞ�Wu'����}k���q���v���p��s���v��1�co�zpH���V1ՎF
Eٲy��Kb9uc��B�������4����ܪq�-Y�Սv�z���7H�!���.���!�G_qy�[����oq��;2Y��я���6 �e`ި�p8������Y��(�{c��۫�ܛֱ��A��){�<��ӧ���F��6�=K�~ �H��ď{���M�JJJѡ�lP�PSI��s�i�(b9�q(�h��������)9b
j��:
B�.d���4�P�M�\�#X�j�:����c�HS�
����٦���1)E��G0�&�T �71MkMR�R�%U4QI��V���!���;i����46��f��Mib%4����4��Q4E[/'�-	ȣT4���:qh4
��N�ljCl6�+ Қ�(�RD֐�ZJ]�д�%1��.��;`\A��\��э��N�h�u��*R�j����
9�փF!�ؠ�5�t!����cd��AUF�IN�' ��ZM���h}HI>1�{�K����fr���ʵ�J�)�HO�,eEZ�L���}W ��3���{oG��ps{囊A��*�]�Ky���/���_��W���ok�Oz��=�~���_��'Tx����o�]讆-�X߽Qݤ'�-�}�J>ɜ�q>����\�l�1ޙ�,	�W���{�~�hAո{��]Y�ԋ6v����⻰^�+�tN�~��'���X{~�_��+<�~Z<u��L��!�=�岗f��c�Y���)-��v���w��Rڦ2�kŋ�ɟq�щ��v�ףwq(Q�W!�9�R��W�
���O{��m�we����b�~���Jت�Ò*����T[�u���r�]l�?�:�3�?Bhu]]�{�s;�ΰ�v[3��6�����d�1M�SP��z�f�z���@�:��a�����s	���x�l�)z;/��[G��F��.k�͎//<2{��t;�sL��G �n�U�'/>��h��Q+]$^��x�*��X3F��M.�����AM�2��].�Nd��t����9�K
�|����#k՛N�zq�UUn]���f:��p��}n��q��,x�l�:���Y�r������3���s5�^�
kͻ�Rݧ�!+�Q��DI(��(=��	�/��i�>�����-fR㴉
%�v�U�fuY;>{"�K9c��W�"au�{`|���,�ɃcOT�ú��v�U�6kG�m�1ü�a]�奉N�}�Qt����f���.Pu."��� ��L��e7�#�z�&�x�B��ߌ�T����B�~�{�Vi׾cΒ�����'�W�wO��ճ�_��Y���{2$U��p.U�f=�F�<����`n��z&&�W�ߋ㻐&\'���ޞv/����د\�� P�/b����i#U���cw����Q�}'�/Ǩ�xuP�n5��7�s�9��T$1}
M�yjyB��aw���G<�%��NNOg���p����3Q��j��~���gG�vG����;1ɸ����^��Y���<<¬����,��l�l~?,w�������Elw/��Z����܎�w㶺vo��7����;�OHG�>�yq]��N��`�׮LhW�fE����{�G��ݲ��֪���_�p{�u���5�p�ƷI�,��{��T��d�:Q^���
�����6�ϸ��v�p��˰.��]>�����Hz=����:�b�3ԝ�9Ǝt�xx��_b��y3�2�ٖ=p�_x�_�����}�����r7Ƅ	��1�]{�t�O�U~S���'j��=�
�0���`X��k��՗���x��]�b����$�tNr��a.����1�0�ev��8���px�2y��тI:���ܒ{���B�$���ن��Ȩ;"�t������`�Õ�3kq7=c��+>�Q��5���*�	��y2����<�s\�z5�x���S5��M�z9E.eB�⏰���R7)Tz�z嗑�@S7-�r"�����E�E�ɔ;0����-�\u���n�:;B����ӟwOi�W��eK1����K��UHʉ��Z���ޜ`{pq��UmYU�Hu_��pϻ�1g��w�>�=}]p��3b
��%�~��v��k���7֡l�9��',�A;ǳ=P�D]n���Twm ^v���C��w�(�hK=�5Oc<7B�Y<�|Hޛ��4*�xp����a�ԕCP�_Q�t� �/5�FD��%g���� ^z��퐏
�_%DM9�d@/��p���K�G[�w�<9��t8>Wz�L'"ף��rN�H˽`T[��"�QϦ�^u����^~��� �+�ٺ�r���-�����90��N�e��}9`[��.���iF�z3�����%���ybw20̎3�:*��.}��*���d�t:���vnMv|��*9+	���gj;���jd��*��F������:;�ưd�E���
�����Y��vY�1n��8�.k�r�vKڻ��i��^5RL���aY�ev��	r��v�Sx�� R|���]ݳ���pN�o!���/7G���q6	�Lb�J~z��3��9�g��1�V9k����J�0W�dg�΃>� J��?�]Q�.9+tVwU	Д+�\jt��ۗ&1�N�/�{h�D��Ý�	}����{L?Z�`Z]^�3�1(�o�t'��������z�٢�v�QGK�/���\ez�^O+���o�����@J�Y��,��ˌ�#鼡��U���g�l�:�y��ר��t��_�<��o�Zx}*��ʥg��7������MSKƄ��JU���-�Ei�Gd�M�c��YE�>%�^N�����w�O��V��ػ���]�w/u#��#c�+��y�gewuj���C�j�B휓������9ۮn�߯�}S{�F�?y_�j w�R73�v}���`��=�s��m���2
��7#��\��#]��f�{߻�-�}`/tMF@�r2��Ʌ��z��"�#��\�֏����(��ӑ:a��^�*cg��:��7�L�;g(���[��fL=.�j��H�>��evFa��vE+�Nx%���sk*GCuN���p`�}$������<_{��=�yu�Qߝ2Ot���)�(��Ư�́G�%wD��=�a�H+�-�ᛌ�,}Z܈�z��G�����G:�̾=���b���W}r� P]Qg��c��q��������y��K���!lw���\ź�#��E�Uu���/U5��8�e>����^�\�=�y���D�S��ᇥx�����A�P�c�����4�G[����9]�9S���D�[�$ �s�u�\LM�d��9}�q5��.[�G�����	ᕪ��-��㇝S�:��8���:m�5\��zK�=LX�=mud��Dt%Ы�1��d��=N#k��ZXm�n�x�r�;�!�P�8��~�zN��>����KȾے��G9Ӵ����o=ꇞ���/I���C�_7�|25�#�X��G��*np����OF4w�.�9Sf㐒� ,'�8D^Ui��c�gC׋;��{�f��C��CQ���G7E��*=wz����'|nz%\O������W<+���G�Zp�B�M�b���<�z�@����Ӡ�N����"
?w�6@?!t�����ǯe�}�"���x��y���jC��� *<������h��9j��S�)��=>�+w�w���$��g�]A�t^��+�.2g�o&X]�R�k��s���vW:�C�;�)OH���ǩ]az=R@��F]y��7�C���IJY2���3;Z1����%t�_A�Y�b��,v�*���4w��,��RPT`"M��b _�^ǳge��鑦�2dj�q�>��oUƋ�<�%)N�n������GLa��C�n���r\^<%O��J{��&��:��)���aq�O�{N��#����o��S�9�+:{�e�^�H���
脪�� Kft�h��7p*��/"=47����H��ۯ_󗿿	�}��829�ǰ���S�Yy���پ�@=ʩQ.�r�#�,'G��yP��b�0^^$�]6ĭ��^V���]�vC�rx^LKF��a�������a����e�U�N��^�r���D)c���;��o3�i9�$y���ȑ_<�7�e|`��������N��]]�0+�{���ƾ�:�N���f�ݗ���Dq��;�)�P:u)��O �t�{��u~S�Ծ���&&)�z����q݃ϵp��U�ȃ΀��� 
�iG-�{��w�k��d''w[�W�����U��%^2=Q}^�^/Ǩ��*�_Y�F�k�#w>�ի�>�=����w��MOK�5<5���N���3Q�~&O�(ƌ^.����E��U8wl��[Uл�����>;�^�Q�}�K/��?��N����_�� �d��2�]���M��~ڙ����\07�SI� �,�z,�bN"*��|��CÝ���b����ˡS��G]ŭ�.31mL���!���z�o.p��} ׷��AM��{g��:�j�xOo5ҹ��n��!���.Qu�+�ו�.#in疩%%�����'���a�ꀣ�����z�M��ό_.&��-���㣞�ߝO��z���eg�~�_���׏����\Ū�@����gܫ�o�/��w�x_˼kt���}���M][n��7ez��gV��1�mH���5�	y�q�]Hmrv����P5U�鉮5���Y�1d�80��E2�1]ü��M��	�%��5��9�|^��gV�H�����F�/���,1�.�R���jV
Ϫ�ި~ɔ�0��*5�OpF.��b��=��T�i��2����Ax�=pҹev�ʖ���U�1S����E�s��e�t���(�8W���V�a`-�:�O3�*_\u%��8�G���$Z�}6�z��m�k���:!�=Y�aT_W������@����Vt�?������Y�]7��y��UH�*�9�{3�T,����wJ�z��v�B�ElEDy!�Qh�T��{e�J����y>�SB�/k��Ĵ}��-ڇp�o���{ՠ�)-�E�I�^��Zj�}�aq����hȆ�\*uf6@�"݉��u8[оi�/q��A�N���v��Fw����p�F���=���1��>�:8�	�"i0RG�>wY3f/>�VL�r�uI_w[R=��_\��Ѯp�M�17��+����4+M�z75$,��9�Y&U�N�/��STDӝ�����	xR�5��LѮ��xG�������d��d暓Д�����y]$\C�!��7Lz�΢:��^2<ϸ�l��:���4�<�v����Q������#�S��p�P_.����e|��m����l?����s��p����
���P3Q�A�'��[���t5NGt���5d<���科��\�^�mS�MN^�ͬ�+��g�c{=ON��gb=L)__�uG���rv����H]g:�7��q|�W~T�^���u9Ð��-�� W���UI�~c߄���B������!r��r�����z} '��M��P���>8cCړ=��#Q����d��lgR�x�=ӣ�g�3]��t�<ƭ���W���tnr�~�v�k�H�yq�5�2 ?{�E��z�r���1�s�1��uZǳ��u{]c֭q�Hb�}��z}q�����ޅ�Q��d�M�\Uhs�X�?s�q�W�=���ػ���2��F̅C�����\�����mի�g�޳�lL����.a'}+�%�0e�����x��ǰ�D��W�
[刧�z���q�>�� ���aѩmL�/�j��Sh����`ji��J�ҶQ�{7l�s��C5�)���%g��Z��m��n�z���;�R)�n�8y���7�]�c�Jf����_^��q�,.ͧ���}~�Oi��c�.�b���C��!�Y��K߸���R���L��X	��d	�}@TZ���z��__z��.�9�O��<��n�S7g+h��.��|����TYv='��t��r"��-��-�G�5�P��ZG3b���.���w�qF�ﻸV������zKQ�@h���L�.{O`,/Ͻ/��H��>����q;��}��g���� ��%}'��w��U��$��ق��Ҳ'�s�|�WH��Ļ���;���]����+Z�c��ʮ�����9�T��.'��8Q}�}�e(�����K��G"�Y�g�g�S#��������q�U̸����t9N:���\P�:m�53���ux�FI9���?V-�����x������U����*2Ǿ֮�G9�3!��yӚ�;��4U0;�I��H-ȃ8�{&�z�M�zL�z��̾���ѕ��	�t��J��.gBp�U^�#�6o愔r�z�^7�c/����+f��|vM�`l}͂��.*����YcM���9n�F�Z�GY�	�ǵ�Z���S��x�.�	�\�0	��]�� KfR���"�+パ��g{
�2�#�l2v�"���NxMp1;Ͱv��-TpYT�Ϯ�����m}�F(���Wb��TǓG�q����׮e���Mxpϧ��G��'��\��s�N����z"}LfL�+<'g+ȱ~K��=�k3'�\���]�*SΝ�wJ�X�*�}gL\.��������Y���5��������C�ϑ��t���6��*�=�+F��f!�s�a?xSe�l�}qBR�������o���m�ږ,�G�&x'���ad%��9S�}���ne��Xނ�e��/Vv�b9���]7�8��j0	���������~{v���Nm=���6������V� �g�����2�~���Su.y9y���ۇmt�ޢ�ݤO���w����i~5V�F�QG������$^˦E��zcazct{=�w�������*A��lÎARg;d��_[�u�t����lك���Bq�1��5���/m�6�+�x�J��;���=�L��ޙ�����7#�O��.���;&;�|�D���)8��bb���@H�A��Xj�����`�u�o�;���@����_������\ ����DW��_� ""����"+��DW� ��� ""� ""�� ""�� ����DW�@_� DE�"+�`���"+���e5��K:0��!�?���}����
��EJ�DTT�*J�H����dB�J%+fD��[P�\�J�)�)"IT
�R	<�r� ..�V�f%��f[R�mKa�]#
���� ג�ٱ*b��iZ��ݒ�KM�҅��v��̪����u� u�;�)���2
���HCE����nƇ j�#J� m�$v�(�Z�J��u��mb�l+V���խ����(�j�D��i�e�ƵY$��P�5�bd3ilcmU�d��;WZi�l�MbM���d�Y���
�n��m��kM!�SkkCw��   L�2�(��2`�@�S�	)R�` L 	��  $M	�F�z&M�A�M�O��J4 0 ��A�d�0	����L&i��S� IR�f�d�  A��&s�ʺzo����;uug��V������a�	��%�2���s���?U	IV���o�W��~Y�ަ�%J��D-F�~��H��C(��HʐH���ϕ���~�n��� �,�b�_��R�SJ�OOm��^�B�����?�t�o��g16A�;�y�N���7XE�����n&��n9Z(^��M�2$K0TB����b�mk,YT�YT���2�h�ٹ��ͧ@�A�ļ�.��[s$�\����-�11T����X�8,({zq��M9�i������F� ��j�!5nf�

�1�g^Y	Z�0�E��f�� �Uc-�y�4��;���N+�Lg6��AGX� �>&�L��荭ڲֶ�+:UX�%��SsP�#xK�yR��������0�ua3�_7ͨ�Ƶ��(�P�N�j�u58����jefJ�kP%��Xh|��J�whD^iD�"��,<�l�N�����C+)�ܰim
2��`��e��)��5I�X��(U�*X�"{Hi�y&�<���	�AQ�Lb`t�hTjڥH�V���R̩p�Qķ>g0�,��RW�vA@xcIR�m	���	et���܅;���,��b�T1\q� R�K�gP��@�+ZU��7���!���%`͔�[�:�afU��l8HǠ��2�F���0E�D���"��E���iԂǂi `)��92�h:Ͳ���Z�Xn��I�L�Ź�q:��f�v^��r��fa�.�Y/c�r9w�EMz�� �(aIX���P�I�u34�b n����a80�&U��lV½�h����>�̶�ک5�g�3l�H�ʸ�5:���c�j�7��5CZ��uo!��ٗCr��Ȇ��DӢ�Y�TA��6ˇ(��J�hr�{�5f�AL��N��8Uw�Z��/=pc�BB�g ��]����-Z��6�jYwS�w�o�F�T��$�m�b� �x	��#-l�t,+�AJ'�âG�F%zd�ui�"v�z��Fc.t�$;ݙt>4P.-�k�7[YSw]AC4A��;�!�s/#�ܑ��� ��o.��)co/&����5��k:�DŻ�0-ծ`z2E�)t�^e�`.�:�D��*�
���p\����Z�$ح�kn�;��m^)���nn��u��LX�.,�
�C^�e`8(˨�M^���]+ӛF韀!'2���Ab;�����zh	j]��RYFƘ��wSF�M`7;2�}�Z���T�v���vsT/���
͚# ̰��5P��peM4!�.f�VVC�N�Wq�7�$8�
����j��*�3���U�k�����R�K$�bd����'�Ga��[h���k"MU7Vq�8�����U�)�l$,���ҌsHGU���ݴr��)b���,d�5--�������)�:��T5���j�*�,[i��{�cюu<q�Z����Û����ݽx���-��T���gȍ�C��vS �F?�J�+jm�ʫ̺Eh���h�q�����u zզ�\!��Q��-kq�����'��:Xŧ1�.�ɄDNb�B�X�q7
�j���a�,'���YT�i��dƅ�DۛB�&UɄ
����dR"��X�zc5kˢtZ�YB�0�9���`Ķ�H62L]�v�cr�q��
��JSC���hfJU���0�O㱃o��������1�$j�+y��,iv�ŲF1+�A�2��/�e,خ�M�mIHff�9XӢ(�ce�:�U�B���27n�8Y&*�АkуlKIڻ�47�G$�+ST*��ˈ�ۀ�٤�zte;�m�!�[��e2�҅�yz��^+X�WE�ѻ�JRx2�1j��cd�N�$�Y�E����I���tٴ�:���kv}��KE�,�m&��jAM�R���%"%�OE݌�-|6��^��Ž'k�٪�rj�jJY��^�T���ݽv�W�_�_��F�2��;F7��	Q�b�و�X�T N &��+��3,Qm�c��xR/�P D�ϱ���w#�ې�z(0��Q�(�/y��㨳4u�_Q����	���3�K�J�gI�c��Q��-,K�8�	�_Q|
�_u*a�f荀��ge��6�����,�s�'jI7���%i��Lt^@�[��黭m��\m��?�y��y�RQ�3U�=�v
�Z�k2�+�6�x����Z9>�mYE�C��^w!�����<V&(YNj�&��������<���`��t��w�8/{'U�(-Ŗ8I*o^ (����1[Ӛ�����6���gE��7�B�Y:u�=&V�Es�n��Bޓ:	��f����B����{h�����ʛ|9�D<����sb����0sl.S:T[��{�Mv\6�̡4ԭ��w�WoaZ�"�C���Tv���� �2
k��;��!�F�w�E��;l�ˬ�J�Tb�^$Ҙ7N�ى�``�f��=*l԰��F���]�|��]�yS�ˋ�u����
9vY�P�;�N�`NV0�<EwÕ�����z&���N1b��Ů\�DgN��3�C��n�N'(
��}j�o��`��_s�Am*����q_wB�!�dqX��=Z������}�|�RI.��s�ç��jFҸ��z3:�|���9����![�;\�Z;�?\BC�H�z[�z'J9����T�[���D�Ԭ��,�n���'��Zm�cZW�&;'m�n�3�����w!����r��e��N�V�
�W+�;���[hї�[��ri�Q���4�n�;`K9��b�����Y\�tn��:��K�
��Sղ�RWױH ��O���%���,	�j�7�6ֺf����)��!�A�͠�t&L�T��me�{;u �����R�t{%k�b�Ƨ,{.J`��`̮D
�wzmu�%�Gp`�r4-WׄZ�X�!r����j]W�\��y�G'ۄ�*8�x��W*�&�W3}w.,�y��|�u��1�2_o1��ɠ�4/�Z�=u�P�Q�Y��:(�]<;Zzhz�i���vY��p��w���v���<���P�Q�4aD����9]��Ѕ�����f��]��N��[�Ҭ�븫��kh(���]��
�}2�f��*�qw�TZJ���۷M���85�c�.ńR�F��-�+-�e__TncA�_s�vrZ
�ծ���o4P;��p�Ċ��aJ����7�3���.������[94>�0��7tJkmq+
Lr��Y�;,L[i�y�I��B�`�آ_NNn���/���1���T]��(
(n-�"��o������]�{@Z9JW k5jv�����5֥	��O�^������RI�m5c
Q���e-�rS�ķ�ү�&:��õd�@";�.#7���T >��|u��K��ԝeb�H�5ht��,��H]]q��wVSdҩtU7�{�b��Q-���֯�W.�\���}Y�L�J�ѝduL�ӛ�l��U�48od�.���Sy.��燘�u�)qX��J���6Ѓ�gJ�n���XZ�S�v��P��iU��ΛZ�	��5��D��-a�>��G'M|�l����R�����o���~9G�D�7(q�vA�wWw'z�Y'}i%
eX�o�N���V\ŤT�E1_v��[����/�N*�b�J�Q�ެ�P��i1M_N��u�U&k��U�<Yz�����]�/�t���"1�J]LY�d�����V�2���70Ż´�[��c_%�/e���)'�V�)�gQ5"p����#�/9QS�Q��M����X�������w:�����/���+��M�[w8{��dS^/�D���Lh�ir"��T�7���mn����3�[�+0�3�[ȣ�����mY+B�{q�3_,T�t)Du	�����;��t�5�0�]����i;Y%���!��P��5��9���sB�f�ACmp�c��V]�v�S����<5$G���s���fF��е�!�;�)mH��������Чs�e9�僨���'S�W��J�B��Gb�m��0�G���*q]�3�:<z·Mm«a�����mj��-�Z��掋��<�	�yx_]fD��L�GyW�$��WU���Ñ%v,u���F��ٹ�s�!�Ն�f�M�87f: ���h:v[��i�@ݩ=ܫi����U�+E��X%s���/ �L���	WR^�JR����@�%B�8��Ƶ���k^����-"M�E](�5�)��m��=�A�&����k(�]v�_:��sD�1S캕��[p����%�q��Q�om���s�l1:^����)T��+�ô�ۖ4=,��}��kG[�0	y���{��k���ꨂV_}ww�IT�Je�����,�o�ΐ�ZJ���8��j/	��ak>v��~1\ZÑ�)ݼG���[��7�ԗu��,�����Z6
U����f���{�WV�]�P���5��3�f�b�}���v#;.�I�d�n�{WTv�
�W:����~�>�_G�tdL��u����`�e�rZ�������+�t���hl�g�Z(s����6Bu��Ҡ�+�c����{bR��ro����Ψ�aY���Ž��ZĶy#I�♪��U ��/�u���0����wX�b�N�O'9Zy��4�������c%��5�ڰ"��f��7��k�s�cY��Y�O���oX��nf������S���.��rZ��]��]�}�nUHF�W�D1�e�18/��LX*�!�b}sn�9���D���3(�T�zM"k��T�
^g<b�-�Tn�T.�c�^ ��������G�Sw�D��Qb���b*��Zm������6�ژۄ�X԰�rժ�**���l��nm���^��u�j<��Mh���ru9�N�7�أ;�d��X��$`�&������9�����l����kY���Pz9Ȏqk!���:�!���ͬ�wC�(�S�4;�t@I��˜��m�]i��aZS[�R]��|9IB���B-��ŷOY��^�I؁����V~o!��oq�X�u����yc��i��n'֏̾�)ֳ�p�ǭ��vv�w/]lL��r%c�NK�8]�X*���JV��U�f�>�AnP�>�+*Mf/�=.���J�d�k�GY��<�( �}�/0P�0	�j�h�!c�U���J�a�N�*;��OcH�v1ۘyk|,��uڥ�D%�gm(Nms!�!�5��}%���c)�u�3+i��Hy�;n��C���ocxً�:(V�O6��������	�Bܾ�v�������	�P�-�fX�˾5nK���;{#��F�0(%�][��ˣ���׏[9D���ȱ��oK��w����թ��5�5uL�QC�[`�j��6�s)�Sd�|�������gJ�A��Ӑ �+H������<'y�Ի�<=w\WuHj*K�'$�L��j�"t�7��5k��פ�笼�w��b��ʺ��h�΂�
�9%�3.g�q
�!������DT�"�Q��ja�6�ذo��End���l�ڤ���p�!��OU�.f�שwT�]G�GLѠ3"��]�{ܨǘko�pi�e�[M�V�N�3;���wYACh)�ٝ�5�Y�ģ����N�_ٌӥLZ�i	r��d������j����  �B�z�T]P���ߢ4�������'��G�~�d[� ��4^JҾ��vn���̔�T4c<�$m�-�I��o��[��V^c��UBT�5�v�[���[�5닔C�ݽ�jP�)������?lKY�q�n�4���'8N���eR����Z���Ts����(��Ul�}��A'�.mn�����er]}�r�EX 2���1��N�Uz�]N����w�2цE�N���7&F��r�;7�����R�:�e�e�Iw��Q-��e�[�������m˺���0�L���%���bF�G%��&\����$$�ɍ�P�E�nYp��9-lk�r�e��R�S0��.��0�#$�\���˦�c�$�&]��T��eʒ7y�,n�!r�fB[̳"Z\��0�*H�nB�Fլ�9d��[bܹdV�H�r�P�ET�����_��{��S+�c����k�
�����j����
g@��ɜ���]�/Û��]��sOZ����:go�r�M<�v6km�A����)u{VV�$@��q��0i�<�}�͎*��g�k���'�������6^n�r��FhNwv��}���u���6�w:�Q4�;��Z&3c}��Iqu�K���wW�w\�3Qf�7�4Eȴ�>fY��go�Y����ս/酞~@��>i��{U�'�X�Q#0d��wlt[�xIF���g�4�������a�=sE=�%��N�৘�0!1Pv�OG]K����w�йs��SʝD�6�]�g�����b�CS��(�N�]g^�zxԙFۄ6�=3�2p�v�F0fMܸ���OW�ח��V�1�\[�C4��,��U�tEN�ْ�-�1R!��^CO�0�xU��]}' �f'YVL(&��FNXM�=�'�t+�ZnH�}Gj��D�OrՉ� N�o�VV���م�<z) ��$V�w��!��ΧIH�I����z\SQ���u�wE	�]�������v5���}�'/;������Օ�Q��)��m�ҁ�˔
����mR����3`)t!�s�Ƒu�td���$�;���d)�j�09@�/�Iu79RY���w���I$LW��{��dX��9�@�X'����𤧍���w����ǽm�<��uX�R�\�f����]�w3E��Z�ֱ��j�T�û3���>{�NO�A��~5u䳏��b�{)�:>�Ey�����)mk�ݜ��ܠ��e�w(àr��	�i|�*T7d��\�a"�+;�#sD�-Jg��E�f�U�.:E.��>@S�}�7��=��V.C������M�년cN�z��uwޅ�&+�����(��՚;����m�Am�����w��]֠ڙ��k�������ݙ�wntΦ�;}[(s!S��G�Tv�B������/8����G�Kk`{I�TK��U�^�YstxX���_Y<$���8(�ׅ�rn6V�-�B���oz����uʯ��Ǩ<�T�f��=p�b�k�h+��F5�V�$���h�[�ڵ�vh�&z{��Z�L���]S3���N��"�zK9�DA^�f�X��O{�9�1��N�f�
{->�H��(���خ�B�>Re�ۗ�jܢ�uF��u�ع��evRpV��z�`%�P- ����۸�Z�Wѝ�a����\&5D�ם��<]�\�g�B����U�����N�#GjK�Q���������lx�je���y��Ja{&ĤT��-p��U4����TY�}Mg,�b�xN���Iv���4Q��^�z����L�@��v��_��EK��ڙ]ܘۊ����W�'Ќ��4���+�ot���=�|;evj���Y8/I����]��6��q���`��̵@�m��ۊ���@[]�C*����������L���W��qkEe5�Ym���sb�-������A�82�uM��f��ڜ[�gr��Er��#�B��l��Z0[WTkO�}DJ�Akq�v[<�c�*%���&�RU�>�_���j7&y{t�0C.�7��0 pڹw����L1�J�!i�%S�@F(��wX�3>j"K�R�Ŕ�٢Ky1�PXQ9�ɣq��p�lő�yJU�J�ػ��(I .O�	8u!���+OS��D|kC�V�8�er��X�e�@�j�R���LH�2���-ݳ/ ��1���*#�|�r��d�Lr�	.U�,`҈�(^e�ˬe�ZZ[w�$j*\�-�eܔ���`D����&$$�Z#)���%�d��%��Ks�BI%*�%�̗0Ɍ�)�F��*Z�H#-��rH���-���n(�p˩��Kę�0��Ѣ�O߿0�M��ުs���l!��g'�wJ[/DM�W����ޥS���>�M�R��*���FW�~anϯ��w�?��zQ��귛E�,�$p�Q[�y4�Y.��v6.N5(��]R2�\`�R�A˸��\:q�N�nRbG���C^Ҭ���\�X�߉C�aA���W]�==Gr��z�,�؞ַ^���GL*��徒��t�c'�%i�z�VꜴ��l��|�$\��֭�ݔ��-[!��u���i����y�E4�֗b	��E�~�� r.�W�&��{b^\N<p��b@)�k�����!!.<���q�K�%	ޠD��Z�Kz;5�̘ �U��m��q3[��uo\�����0] �SK�,g��������h,_f4���^]Ȁ�Ϗ(ت�Oy�)a�����H�T'��/��Y���f��]A�+E<?���p��F����R��z���ƕ��>�}1�GR�4Tj�}(�L�p�~�?5UX��
�A^��U�T~Jƀƪ�4h�mV��U��_!GZ�J�h�檉�Em 7��4�~�˾��n�+B�j����@0J���m�Uj��op�;���U���2�*�1I&ʌ�t�jC:"�*�J�@�ߌ��ޙ;��Tm
�����b�6P�$¢l��	��U �9>�6�A�q�������q����WR�� �A߫�ފ�Z�U	�Eu���W��Pq��Q���GZ%U|�N�z����Dj�#AU��*��z u�������5U�g7r{���U[TQ<�Q�%�R�ƨ�P~h�/]�����^���C�X�C�7�s �M\���o���ʛK���t`Gk�/�z=��߄ǽu�*�E�Z�6�u�Km�gH[V\����Q�
-(�j��*�
�B��UV����js9��m(4�Ԡ�cA�+�A�!���Z5TX�j��T9
� �o}��UƩM�G��UkmW�+mQ�
�V5U֪��@�E���?�y������u�AhQƠך��F҃ʪ��*��EZQJ�9﷩�k6u���Q��\h<5Fҍ'檪%VjUQ�
6ֿo�s?9/y�(�h���J)�Ti��UW��[�G�<��{6U|�m��ڔ�V%Ui�R���UW�6�G�m���__5UGw�E@��U�� -�� y��g�W+MW���{���V�/���_�F����ǆ%|2��s�.����US�^�_
�\���r"�]�����~���O��nA�ۺ���$b?�<.?x��9,�� hv���'�r��*'K�ŷ���v�$��z�r�U�X�O����N��*c}qWg�}���v�'y�0��gI�#SV8s��u��gF(8\�)7J =��7.�R�PInћ��3]B�r�����z��������q��iR�O�b�������w�ȍ��������j��9b�"���Y1�	�p�
����\t�x��A�l��"b���s�4_IKWޞ�w[8Eg����9�W��V��F�%).�_/P�(8����j�=i�[�U-�;������������>�1���� g=dJja�K&kvud�GT,gm��j˶;��MV�+_��*��E]3�=�Y%sT����C�me�����9Q3�ʵ��=;�>�
�"����k���r]dNu� �2]]X
��];tc����e��'� ���?����#yo��'ur��z=��6cBwo�3n�ת�W�9��g�^��f�ͼ�'�{�<�� �՗Q
~+���f������7)V���fm�L"�}<�j"s�O�#{q���:.t���,��.e��d���U���x{�r&�^��P9�PZ��zc�ԭI�VWU{�����Cik�3�!��73�Vu}��re�L���й�;��8[/;�C*����}n�/�j!}3$@kV@�W8�'�Qu��̵�5��Ȑ2ĝ�coU����y�����u9U�T�Hc��w�7]�g�>���儻��D~́jH6q�w�;U�Z� Mm\�L�qek��Zp����٪ٵ+��@��*�c���̦J�J��]34'ٌWJ�78����t쫌�Qi�ܓE���y;P9}�y��	���z�x���쵯��Rh��.	������L��gK9��#DX�$�-���7S��7�;w&N/%��iW8R��f��v����52�g�+E$���M��:u���A�Ŕ����H"q�ti*m9��0����Y�#b�0���q�6�
�u�Ôi~��D l��Ɇ��Yk%���,ɗ�YicN<W�ژ/䚧ę��V��L��I��40�11,i�P�IQ9r�V���K
�(/9�s.��ֳ�^��}��k�iF�'����0QJ�ə\UA�l����d��.*�����w�Cu��T�������r4�he˃����d��B�QU�q1,�$$#%J%�x^9�EQ�.T�H��.�H$�ܫ���s�R*��h-F�wr��6�ԤbKb���.'��o_���ٟ���.����<�j�����F���{Wߟ�kw~��RK֭��W|#�w4��2���ތ�Tՠt�ׇ��G~��qY�����:��z�)�́Xi_ і*�x��F�7�y�ljh��9�b�z�6��풸y
��ڜe!���X��q�`���և��]��:w����Dkj-��J��^���U�b���M=�1M#7t5H��}k '-.�-=���N]i��x���Y#B�|���^[�f�Nf��#�1���ap̥g<kʵ���evEv4��x������Ĝ��5p�*���R��7)d�<�wT!����b�ڶe`���[��{��|���\,U���ۿ���ц{�tVe�ᬵq�z��2���'��ӛ�w"S��S��^]�>E$<�w���z�y�%�P㎻�W��mg���=~��u�ʬ]g��ݞs��J��(m�YR�A)aȟBNʍ
M(���3'/������y7�@y�c��:�w��D��3R�}��.�NE��Lj�:���P/ٙu�0r���6�����L�z���U2�)��A�V�WW����S�t�N�W�Z�)��ғ�<E���^Ҍ�g�J�!Xw6���⢏�gSO��5y�;^	T�h������g}G�����TI�E�74�{�T�.�95����CI��~���{�/�*O�J�۷�G)%u��e�ґ&��o�®�&�l�+��,��z�g��ҿ	�y�5���9��;���b�zc�� 5��m`Ϋݠ����{��F'��{��n�hG:J�B�����&�k�
�Do�j�T��QU&&c=<�FY��ն.h�V�MMό���G��eou���בC�#��#�y����)�H�P�D�t��wNom9�]5��-��ڲ�/�^�<��AZI�ts�J����΢f�}2n���F�kz��F��U�0����+�B������"<�:�Ei��\hH�j���{5��uح���o�dbYvy�F� [O{"ꢧw,T��B�f�P&N����-fXx`k��H��f�c�M��!����[d��V�7��_2�k)�Z����8y���\ǖ�a��Np1���u(�B������=�>���{�aJ��wig�=�G�j�<��FS1�B��;����a�-N�~nz�k��>.�{�{M�Ø®��s���Ɵ�`��:���Y�/Ș�q'u�>n�B{�vA�r��k,�A�f�٘U"��)ç5n�u����������++^Xݭ�Nk�UG=ߺ������~ۆ��}0���/l��2^3�sBuֱx�a�wp�e�-�	��"���+R2]_J��OD�����1ߴ�1R�IJ�!�;�iٸ�y�1�6��u��:�珜�N`.��xx��m�=��6�LC(1�Qa=��r��v(�YiD�p�I}��y�y�e�%�(l.Dn���+���V�yW���ꜞ����`�5�\ۖ�?O��f��ɫkw'vN}d�L�]���F���\���I��o�}�������G
�O󿞖"��&.��wf����
��:��.��&T�F��sDTU���s8*����vM�ܦ9�#�rg(���\s'�y��h��$/l�룼r��|��������G���]Id�	#�鳑max+���=�#t������1�sE�L���e�9ҹ�g(�7K�b[��	�nb:�Ư6�dgb>��|����`U����f�s�� 
YZ���թp������;k��O)��k���(,�4�Js�I'��i�h6idf��G�cØ��v^�2Ţ�)�m����U�"F��
�һ��WP
`�X�r�"���.���)�$&�j$�6r��cm˱��wWXbL��$�m�,�E0fժ�8���ʟ}���B$Qn��(�$��rљdU��e����IX���PiB�J���,���r�]D�Є��,�%��M%HE���X���w(D�.֔-a��!@��:w���Uewq��p�+�b_��"#ɦ��u_4.'���6�gq���'M=Z�g��p�7=Q�����5�j4[��6E�����c�Cݔ{.�K��J��?!��ϝrV�ly�|��D~�зڕ�TL�P���r�5D`B����Xc�i}�'�o�t�yƭ1�ɧ����};���ð�YG԰lH[�x{��+w*Pv:��}W��i�X98�R� kl�����(��������y�X5��>圞��7�E�s�O�����{S�d�����5��_��ݳ�ާZ�K�V�=ih�muǉ��߳w�>^�5d6�>ChL�X�2���w�N��\�0�����+j������V�Ƶ�}�]{��ı;��;�/p�3{���U�����4��y���_&*K���Wɋ�;�y{�O"���`א���\5�A��Pșݜ�5ݤRć��G����6֓��՟:K�9��m�F�X*��%%�}�{�MT��>�~G%�� �Rv^{��{�_�Nӭ7-��u�o>7[ܯ���&�wS���[��ٛ�}�M�yƖ#ۼk9+�C�}�y�\O8ҞE=��}�o&����Y��-<��ƴ�5��v���gɷrv�nW}8�fO[�y�nY�j�~|����cKI�&�kdۓ���D�[z�5�R��9��ˮ�p���}�HZ�!.��䓩���1R�M�������,�=L;�uV�hj�zA�m?&ǯ���^k�X����Y�7	�w�6M���n�����Q��כg��zM'�|j-m:����8�ޝ�|w^�_��qjT�/��])N<O��ݟ''��h�H�v#"}S;>sr&2��aeF�f'Si�-�P���c��f���}x����b?Cw4��$=���}�3�b��D���������x�.���1�=��~�₃�{�ȟ�g�Ӵ�?���+I�f���.���o�YcV����]�{j�q:֑Mk�m�X��i��~Ѥ1����6��19��ϓ3�����D�%�\6�Ój���z�[1nA;���{Ϧg�9���o����4[�B�ws�l֠[��LHy�ɋ��V۵I��S���c���J�����M����M;�2��V
��@b.��>�A����a�߇
l�_]���FBzrچ����G�ƱkF�FwLTq]�Z%G�<~
������5���k߹u�{������rm�\C�b�R�#c$������bm"D�m|���i�s��`���>t��*y4�`����ƽ��y�X5��7���4��E�1�u6�i�f�߳��wc��R�n�Z_��k9g[����>߶��O=ih��vV?'_a�o�v{�����t����@R�����*���|~ct�LI՗6{#�5�u�Sɳ�_9��vl��9:Oy~C����%O���u�ܲ��q7 bsP�kv_��U��߲������u��&*ga�޳�+e��]�}�6��'�`�q#�n���_|�5|�0��5�bLh�C��H��b��D��8}PW�1��hI�9��ڹ'�J��V�7�;��q�3�Aa���b����4hL5��}j�����f,��/�ǆ���T�QQX������0+S��/
6j�Б��b�D�&w�/�N��ty�8,r{�TU}������k�<tҖ��d3�9��3�&��)i�ϛh���][��a��P4ktzpR��*�>���.�:T�T�d�f�3s�@�u�-u �0t�ׯW��z�vi+hM��az�]M�ϋ�r���؂��N�^�r�Sd���P7�Z�J4�����s~p�N�;H��]��Ny�s�Ǜkɷ�ݗ�m��8�꽑�3AB�F�G:6��A�����5�y�^������|� Uk�g��*��x��'5ƾ�,�q�!�9���}���|��gҶ$z�7+�m��+��7�'>�V�h�O����=��MC�%��'vM$cW���~�M=LI���M��}
y�ܱ���t�Z��{�m�����Ӎ�'aE7~�o����Ͻ���j��_�o�{�Mgu�/��-���&�g��z��|�|կ!�8�1*ݦ����s�8N�ح�.�qN2���6��%�z#og��M����D=k���+�ߧ������1K��\��p9��������.�74��~�:��v�u�7so�s�V������O8�T��ɦ��i|���=������85湸w���H�ط}'T!^*�����������{�p�B��L~MSn�}�oڮf����ɷ��N&&��J:�*{�J}��t��ۖ}��W9v[�_��<*q��"��*�xz`&C�{m���3@F5I���(f�+�W��O��j.<{�ī����'le,�;�E`�OwB��)t�/�2k;=#i������	�.p��{Tn��,�;���tz�O-��γLjҝpV�9U�ڵ4��H��5�y�k�@�ɶ��6N�����H�In^�ɰ��JjȖЦ�����+�EWb�U��7�ȱ�S����;���(h�Mu�:�q
Q�]�1G%3�C�H�7H�=�0�2���u�3v�9o���N۾V뻲c�ɫ����s�&o!OV��q:�]��Ӛ�[�(q����m���ej�/�JK�a.A����S����Y�|�n���]�/��u�Gb��X��4[�ƻ+t 8�6em.��]>���'
��|�j�[�us��<s��|_ ��_H]�U���e�|��M[p!$Ys,�0Z��Ƣ��Ց��r�!2Z9��Y�"(�p���:��L��0t�qm��k�]1˅����	h���ݑr@TiK�ńP4��A�s���}�;c;7��LU�����m�z�	��G�"LNTZ�nyײ_o�j�iO!mN�\ߥ�_l�ǎ�=�w�i�r��q�'އ}=�c��X��5w�κcN�g�Vv����|Xw1,��__�X�/MK��[�]����~���:'��&����W:���/�q<�c�b`׬��������l��sX"֛b/�5_�����<��1�J4�M?$�u7����+�if���+�tD���P ��;[�Z�N���}+����U��Ҳᦍ_�Zm�r�Z�Mju�ɦ�;p�*n[�G��y���Jަ	�iz��Y�������޾��i���m-zK~L�y�}���C;�k�^3R�"{5'��k��4����-M&�j��Y�w1�׷?15��ԯ��=Y��J�V<M��6+I��/�����<�5[N��<�:���������ij�(#T��
7
�X��=���ig��:6].�v׭4��Ԇ�i�Q�s~��@}�h�_�!����4[ְL>s���ƿzu<�E����l����!�t��Wȵi;;�Y��!���~��@����W�Ι\7T�6�55�.�<O9�}�ljƴ׵+n��&�m�d�o٠�tM�4}��ƲJ���ɿpǧ!7vcn$��h��id���i���]�K5�c���=���5Ƣm�^����k���P+c�y��Ĩ����86U��U��9)a4�+�wBSAV��ߢ=��y�~h���LT;�i��d�o�D���nWZS�mD}1��I���D�!��4��%î����z��t�O<&쭦"��_�_N��HJ��]�UX4`��4���׎x��{��?ru5�n�<&�H[���O�n��^��/����M����`� �@����*��/�9��,t���y�j=y���f�I�1^0�G��?3�J�:�s�뫮�����p\m��vP�[w޾�����;�l��?g��i5�ZD��|��[־���;�Ț��i�'�&��:d��s�0�ߡ^c[ԣ�w�X�w�{�/Zu뮹�B�cBzm��>�>�vQƬ�J8����g�׽ަ�V���2��iKB��#5�{�������>�/�YܛH��ƞ��4�>O�?'9r����Z~����푮������[O���{p�k��Y먕i��s-> �4�=�2�ߜC�gHk3�K�(��|��Iޡ�{	���]N�������}�����i�[^LT�C.mØq�����#���o�kI�oS�2w�nm>wp��M�cX���a�j�H,L䴬O%���Ǘ��V�xפ1�>˩�mAW���:�i��4c���oZ���|�����ە���I}��+7�����lx���[K�2[�7w��Y�+}���붾N<ԥ"oӛ��캐�{��C;�SO����y�������)V�=���õ�1Ʀ�5�b+�:�a���I�"����_T�\�}w����Ϝ�nϿ^�������o�qT�ϟ������1��܍=���.�2��;���;��rR��w����D��f&�N'�u���[�V�ӝ~�l����g��b��5��u�}ϟ>C�Cn���+G�����SI�������lw���x�������i6����{�S[�����}���1�1�	��}�_;m/��Ǉ~/is}|s'���V���P��R��8�Ӌ�q��ᷩ}�=nǾ�"��LEL�3^�#��毒ͧK�8��z��Cn�~��wv���M'jԬWc�m�w�4U�����݆�lk���<���kN��<�q�a��s[׹]{�\q���ǯ]����y����Î�^�Z�����wC5����x�>&�p��(�s��v'_�'�}�mǞ����u��q;�>��7���5V��WGiw��AִͩtF�U�u��)�ciTb�{���]�G��{ﺟ�^���~�Y�Y�I�Y����o��!��?&*q4����k���Mm�]z:nz|b|�ݘ<�<�t$=L󲴅�\�ڗ�^�jșr�i�'�$Kw�w�wJ<5כM:{������JƢc�>K|��M�g�t\���P��"5�����߽j��ƛ��[�h=}��zQ�LLH1�Z|��Nw�l���ō��1X +=鱻^�y2�ep���l���n�yӧb��1�b܎�Q�K��}�4�ϣM�����s&;��adf3<�Wjŷ	"��sӺ[;��	r���ڔ���&Au��.�k���|i[2�W9�i��YK�K1���NsqM�2Da�p��rY;�
"�af1k/�I�JyxH�n���o2�Q�V��~�����͍�c.m]�p�FWe�`R��d�n�4u�X�31"��8dw�K��]��@���w>��r������1��k�z�$�e ���
�-/V�Ț{�fndB��FV�f��ހ�l���9��ct�9[�i�P}C�����;EX!�K�\�A�^�6l��ڋ�M������:.S���
m��	;;=��n���x���EU�!�ΛU��ɥ���333��]���M#b�z!4��]Cp���,��%�φ��RK5��1�o�ut�
m�����FL��%W��З��F�Lb�A;tQ�9T��Ϋ|_bx3�+�f,v��\w]�9-�Me�AI;f���G�v��ż�'\��lս5�J�}ת�|Q��������յ�&J4���R�<�{�3_��^h������U��[-!���8���R���r-,�M��m�j ZD��jF؊b[n#uvZ �#VյD��-Am�m�R"bhU��u^}�6��!ԫ��V�Ck�/�=�|����=���s�[\y��ݙb!���sC��J��|U�JrUx�2.��)�^!ٗ���9ޭ�i>=�yzI���"����绩˺�¸��{�@+��&�K���^S���oT�1��j/e@��0����!��RÓ��8+x��R���{ܦzN��{�E%����0|M�J��NK�*�s�x%��ܤO���K��6�V����z��Mm����+֎��T0!���(�]WD+1���rot�0am�2�C���F��|�uլd��:W�Ү#Q-MR���I�4TH�sR���׎2�2h��n��]�R��ڔ�����ܱ}_f�7�~C}��O�:+n�1�|��k���s�2�Y���&[�%״����nα�N���dySO�úl�A��8�X
�RU�E�Rx�4�j�,��H�h
ňF��*��C7!mMGB�y�V������Z���x�ʪ
O|�7��8��y�g����Pk���;&o�"�"�����b�(��v�4��t��p�ɉ`��v[���Xm']����걆�Oa3���� 3�I��87A�/�,�Gn���ж�btV�	�{7K*I�]����]'!ei�1ӏs�d���w��������{F����0~{'����z�͎�=l�8U���e�ׇ=#�T�͕[��2$ I{�����􎧁g�a��(x�3Wp앨�5�M�>.^���Æ�d=�V����UNo[/���P��=��S�j(k���$��]Ӯ���с��_y�����+�;�����������ϩ>��׊�V
�0��<�~���̞l?`�K����Ħ{@��"fy�F��FP�7�ځ���y�b���xبjyۑ���4Ұ�*��\e߄��)/Y���Z<��x��i�\,$�{��9�q��!_X��n']'#g&v^QA�R�j����9�����]*��U`&;]��SO�S>E2:U�;���4�3zCc�YWέ�������/��.�L����u\�Zٿu_��LZ2q�3#(��9Kǀ^�(n���p��#yENC:[�����1�c�V0"�F�D��!��&�8s�}�����;��V�+j뱲�?��r������;���+R�A�z����x�-؃q�m�����[���ݘg�d�S��|UEgy{P8��+$9�{st���y�F=��1y��ۯ"	��L�LKF��Y�uvc�Q�{nr��.���nu���{���U-�;�����D4��R)|Lg'��p�r9@3����w�1�A:����X��:�t�{@�r�0��{F�n�޶.�,�GН�vmងs��Y����*�T|�Eځw�f�h��)����|e%B����w�m˺\���#SS��������cWs��*=����Dy�8�2��]�aW�]u�l�E��b�d�=w� 6������ػ��l��wޣb���{n��Q��RU�}�H^]�a��1�h�(m�P��!���w�u�f�y��o�3
������6m�������/-�4�ʥ�EE�Y�zYXM�Le� �^E��������"cݢG-�ۋ��O]'}G�G0˲�5�ur���9Ky���m�c���h%��{�
pN�X��YC��&K�t/w&
Y-�y�~���Tx��::��Y/�t����-��t)���S�»� ���2���B`w@n��o3-��y��(AFl�UЕ|�E0Py��vV��.�^<g��>5��	f�BE0�v����ᴙB���j�(���M�e�s� u2[6YL.�)��E�T�2�%���eT�vhˠ��ѻ8n������GB��a�bc�Kt�ed�n�ؒp4>�M�I����#y�N��������JVu�,Yǅc�`�u��J��h� �:�I�c�� �TbEc8���Z$r�Y-�BҖ��-(��!��m-�jd�֖Hܖ��E1���jTdX�H�!1rJEEjX�U��J�����!w�e9%(�Pc�A���еH���^7�w5,R�+wWӌ#�h��"����Fj��+?��Dy�����;�nt���;l�\�\\n,U9S\��a埌0ߓh�k�jI�{Q^\���'f���w�d�`s�"x�˃��N Z� x��teJ��F�6<�V�\j�e�G��|i�Җ,=�/����r�X�@#�iE�`�c��U�s��n��6��>�~r#K$�(�y���	z��ne9o;xfn2��F��k�{��9M�����Î��ȧa+j�N�4r�+/0�9i�]�<���Y�\�;�Of���A�q����Iz�_4Oe/tО7\��>��8Ot?��~�\G>��:+�\l�w-�=���{�5�#��,���OzG�X���|h�S�.!=�����iKw�U�
o�-�aO7;�n��υ5)n�5�P�n��h�f���<�j|.ꣴ��N����V�ؗ9�qlF�L���K̎��_wN���u:�?7�؇*G}�K0��r��H����T�$�;��wg�؋���ކ��}�wh���~��50"~<2I�F<{���1����}�)���Or�%Em;�50�Y��� %R��5 zY�*��y<&�n���	��m����>-
Q@��<��om	�ґ�͑���ré'3j7^����z�����xGbOeI��q�9Y��w�R��>����}�c8O(F�}���Z�^Zn�{��%�dҏ�K����*�\9�+lZ���C���Z�# ĻU�m�J�WZ�9� !��Qf�Np��3�Ԩ�r`�E���6�F��]�}ǟ��mm_;q��~����U۩.�{x��k�M�ԑ1d�m<�CH+;�b�Ssc�>�Z����{�p�������i��:��Q�{m9ЌW4����������~�Sw޲xQ���X6�5V�P����zJXYlhUܯ�W�E&��c`�lW.GW���襘7^�ՐI��:�W3T꘺��<�J�]�m��SH�;�����^�'
���Rf���	������5蠵[����P��Dc#��8����������S�f6�6lqz�����Q���db�yqRwW�q�Un*�7'^�}0��C��P��{Hq3Z׵���3���NA�����7X���r��4ۭ���{� ��j"���5<O��,��}h�
�r��lZV^�cƯ�zG�J��U�#�I��3�(���%�AS�{�⧯v!ݔ��oTp�^���E3�����P�a��#�?�j��P�U���1s�L�٪wt�]٭z�y��/GJ���㞻"M+^����ƾ���V)�*��A,��\��3���j�eǝ�w�yI)�x�֒Ini3�9�6��A�aohӯ��{k�lh��̄��Y�j5� +�{*�h�=��cTN7��[�e�#��멆�-�Tz¬�H��o��Y�V'���#]c,1��t�vc�b�[��ڄ��Q>5��[[)����v^�A�*��y<=��ӿ�s�>��}��s���clj�W����X�I'_��� g���7ö�c~U��K�"8��2�g;tsQ����ދ�6V�20��]�����,�b�qi�w;`��0�V>��hJ�}۸%�׍'��a_*�8�w�^iqܖ�48�4�:�[X�!;����n���)��ze %v�m�Ͷ��˧�� �)����{���o��z�[����.��{BȦV�̩ĊҦCqV���*��IJF,��V�*�������9w������Mb���,��D$��<H�P¬�kf�\�p*�+��i�L��
�Mc��1uf��j�� ']^;���yxmIF�[���L�LIZ����K�'�Dۡ�:x�c���|嚾Y����E�,f]]1X�ԨrEqS���0��<��e�����4��KiIm�K��Ʊ��-���W.˸��S$,��������"-c.,a"%�qm���ı��̊Z!��Y&LLʻ[��Q�R�#�e�%9��o��A!&6Ц0k#��6��7����̗J�����R幄���L���+):T�w�6o
Q3\��j�3�k.j�Ʌ�3yd�h��;ة��źCC�=�������T�Rm�(�nF|����[\�o�Ufϴ+Bw��O|�w'�BvE�S��񏬤��H��c�ɪpeTl��^�i�yU�NЬ��֨$���5�v;V�����l$�P�Nl�ĺ(�1A�{jo`�5��\���a�AO�X{D(�1�N�;�� ��f��W�ڼ�Xn��ok�6(3[|�Z9|0�^V�R�[�7,�S��t1s�w7�
^��a5J;�qqn�X�('R#��i����ͮh���b��Y5��Yܹe��;ouh�Fz�ݴ�r�#s��Tfb�1s}8�~Cl�T(�ʼ"�0z�w�i���p��r6�C5C^|�b�ʡ[�/�t��q��G��K-����=ƙT�풮U.Q� j�=�;u5tK��͋3Z1��%WM�%�9o���EZID�W��;\�I+��EF�`%�X���K=[�����l���AQ�g���ao����i�) A��ۧ��#g���X�I�\W�����Ű�Ďb���H^]z$�K6D�jt�?CIt�_JH��X�:w�Vc��n\S:�.��u�޾"H��ˈ�F��G$~��k����z���d�^5 ��j��#��)��Qyj��m����hk9:w5+�4)��Ф�ҍxw�LncP!���V���+̼��i��5P.�[ۨW��ߗFf=�2H����;{A�|�#�e�+���'�
Z^��7�3�WI�LL{��u�u��x`�����X�m#���,1ѭ�QmO(S��(�w�Q��q��@X|}hZ�:�;�ޝsUK5a�.����a}z�D�0���B��Cب��॰�͌w@��xf�R����VV�.�!�����x�4 �e��bXio���սpC8a<_v�EZ�s�)��tG+�ʾ��`�c���.ƍ���-X�m��{��MP�5xa+��7ٕ�.G	�q��G-e���DJ��d�� ����x���=���^�:�����ll`�Z>���Ӟ�i�W�k'̠��
=^�1�k4��j���0Nٞ gj�r��W�N���0���S�,�!��*ஜ:�qe�<��6(k�qB�mɂ���Z�A�vD�E�n�{����3���ܸ���s�xP�r�P��|{�uoTT�<L��t����Q�W�F*��K�ɝc8lWn��-����1�ȴ�k�� ���X�gk�[]�pu��0�ɂ�l'�K���1��eq��((!�tR�������3�=+�*�^]�@_3��}{*�I���C�w%~����x�X:	+������^[���Ԗ^�sU�Px��Բ���՘O�o�E��3b��f��є�aG�7��J�!PyV.��\����s��v�Og:�IҀߙD�є�.������y\�g�w�j;�y��5��m��pC6㮣{�7ԛ�(��q�ΧpPz�ga�����(R)�§K����VQ��3���:�@��}��e��<�eh㘉��� �/>�i=��3�����q��`��奓B3�i�����p��� ��]�EC)C(�j�Ňd��x�FS�p��F�ot/䎲f�
$���]&����R�ש�x&���B�=jBvŻ�4��Y<��{n�|RglJ�5ݜx�܄�|��t:��z�8�����[p�~�J�i��hj�S�j��P�bρV�Q1)/*ګS��d���]ȈT�Ģ
m�]���VHD7�P��L�S%�9���`���,k9�v�fU��x�׌T�(��%���@ǗH	�ec�:NG��` ��R��gm+B��B����: M0����TD[��7wZk1�[�̐�b���T��V�u��m1�IWu$�.-�cu��%�XLm\2[L%�%Km��Z\��		RK��1e�ayr�,j�L���!x9��Ƣ8�$�����$,rL��d�d����]�1[`Ȳ1�\�p����F]���Y-�l�YR
�Z-̻���  D�2DT��|��'Do�ƶ��:��o)ܟ����x_O.���7�\^��!�K�m'{ױ��0P��7|_����^�1�]Z��QEU�X�Kx���Ҳh:>�N�NFq������=��HW�AZ!M���;�.�_`Q};Q��Ձ�b�T�R��op�I@�v�7]n�c[��^R�grS��Mm�]g�)�q�Vp��o�:@�Ȧx�\����x��uw��=�|�ZC�~��x�4�Ew}�Eny=�힎	�il�����]�ɮ�1[���A�Hj��,xc����E��,�yZ�a�m=���ř�2u_�����}0�FŬ	���2q���h�g�k�,�qC����yt�D+-Ems�(oR�����,�=W�^��cauf{�Y|�ώ��0�3��Q��0�b���b�{*�Z㷗榓=�x盼��k�����v�����s�����R�ھh������m5��ˠGjb�1kV0��kȺ�+�h�ǘ�y�'nV{N�>��ƨ��Y	I�hm��"�=5���Mn�������.ir=�N��	.f��#|VJ� S����c�,��r��b���bu�ݘQ�-�[�9E�m�/�>�8!8�_շƲTv��fqֺ):w;�y�+Ǿ��+=5]�Bz�}p�I�l��^�d.AW�F���J^�4#�wg� ٪cFd=�K!�v��-����x�W��c�(q��*���M�[R#���yh��;�Rg(v�Wq�P���Bǥ)�rfM^+:��ݻJ9�qr3dX�j�-��@ﯰ\�Ilu#kU��Ҋ�8�C�.k,��%x<�:�{W�Zrz�3.���6�,����1[y��rP�G��̡����n�CY�񊡚��V�"�����8�,�/G_j�yGY�i�n�CZR��4�+�aݮf��:�o�(v�{J�������f۞�^9��d/{ ̒T^��e��ϑ�������+�����kt?]��01�ي;dүtv"sԮx��8K�DA��~�$�6�s;�F���n������ �۔z��{euEI�B�S���v�������1䒹G���Y�����clc��'�H�n�)�dJ�uc�AW2Bf}uB���cgRQvWN&��t��L(c��Y�_e.���ɸty��ݡ<5�*�x�!�Op�x��m>\]c�:=���ad�~ɲ��S;\�F��P��H[J#3���C�ţ:��k=;�s-YP����O�����1v
?��Q�����U}۪�t!����ף���A���+N��p�"{e�C{+�uӪ��^vu_9y��a���q�x���]��l�p��OT�c\�N�*�j�Ʊ5.�/e>�����IUZbR�H�(;5��w.J\r�͓#�s� X�����S��ɀ�,qx&��?l��wf�[�d����Z�^k@]<Bu�G�Z٤tY��+��������{�ٝ�4�T�z��CzeK�����h�CΟ��ݲ.���;otٵˊ�:���4c�1S׼j�t讇ʷ�=R��M#��e.��"��	;eP0��sh����WuXWomݭt7݋Q�ŪO�J���GB���X���i�r�(XYM'��ub����UAq�Uѩ����Q�ݒtV�&�g�ٝX��u�T�qԹ8҆T��:'��uP��U�0�G��V��ٯ���5L%l�@\~���Թ+��6ܗ*�Tu��̎�hV��OL�z.������O�(�LNػeY
G��[�u�/__gKrWm��9���ݝn��ƽO�2_��J��'�-�e�Mmt
�X��v�J�긺��˂�(I�^�D3f�a]+ڋ#룴��>:�cɔ9� &gd��H����#�VY[�HR#�q��ar2�n5�-�r�&Ym̕�s2�o*^Qy��\UQ�5e�1���	%�Z��.Zɍ��e���*\F�4Ą��Ke���n�2d�2B��m�B27hK�.2Ii-!4�Z0�on�Z�Xԑ�-Ō�e�-��M�E$��@�m ��l�˘L��X�r��-Ed�EF�1�/,�"�H+D*\��,*d��m A���w+�|�d֛Ꙝٝ�v���k<���;e���xzm;��7`��2%ŉ�W+�����J����*m+�<O�s^�]��TK�8�onL��n��ڑ��+;�x����C��	4Uay��������c���F���6����'�X;�]���5��'N��|L�rϺ/hu��,�7�t�3���� E��=(S����^P�9��P�n�Π�so�ߖ�{�yռ�Y��'�����ܖ
7�9�Y�U/�"�*�����I���s����(�b�&iR��>����ұ(������k�?I}Y���;���҅.\����+�W�^�� ��ݬF�l���+0��oA�����E���. 6zx��Ҙ���-V����+�'76�=���rWē��~x�.*0EtY=�P�7�V|V��<�����]&��.��i.Y����d�5UFW"��k��`g#h�#i5�㳁�kg���Ć[������+V�C};aV��
�؃�S0�~���}�;}n���Q��M�Y�Ge�'8Gu�
/��u���R�:=,�������3l^�Uzl8U�gu.	v�	]�ʽ��w�\�����V�����xR��R-�5;���*�.M�4�L�T�iQ'���w�W�I}��)��m�����aF˲�t<�3%�쫝�*ۘ���ъ��啡س�04���z�Z�擁gwNB��,cwnЃ��ܟ_����T�Q�|���O������ff�]���}h��|�/�)4��y��C��1�ܶ�P#�Va	f��u;Ё-�]c��\,�5��b��pys�3�T�����O[�e;�����ԩ��\�J�M���|��t꽃��{�d��(��e�fT�]|���`���P���o{���x��P�>�{��\�-��W��W�"����3ZS��s(�eE>ū��t1�Lt��ņE�@�_��b�N�����P�mȚ'��ko�.��A�9 �f`��{��*��˳,	۽I�]�rмRCH��pEF�8�Rѯ'C=x�K�ͱ�	.:�ո�3�]��{{�8Q|{O����D���]g-�Яw��zm�U�T	]�5׈A]��E�*t��2*�,��
���h������U;4V$�u�ij��+��\�ê����=}(i^���p�i�����k�{�ū3���N�)4�x/�[���gɞ�y����+����IS��ͽENur�g���o���nU���:�߯Y� fb��:Lw-�)p�1�^��'�^.s�_��S�w[���N4�/x�ۯn�_�b��Ȓ�Rݽ(��okH�$kylǻM'��yl�����k�>J��_,i���[B/��m�J:���HM��iz�I�hＳ��r0����O��?���1S���UV��qkA�;�X"������+>���{V��l���۵,�:���&6g�u� �����,���Y���΍�y�n��7�&f%���轂 =JJ��iZ��nZ��ߔm9K�?z��/a�.��T�������7?v�߿Uj4�ZJ��݌M1��MpD�>f��uvJ����" ?B�4H���q*��]����/�c�������>�Y�n����_�����;�;<��_1�o��OmJ�M�K�Z��c�]Fs�Y��ZӢ�Z�޶/I-�e�kz/�*c��.>�Uo˾�9L�~�'��f�Z�[(�]�ѓ�|Ԭ@d�]dd��YUUHׄ��c}��-{�~�hrb7�>Y6�`��2gKsg�f992�=o��E��u�����Q�ko�$��y�ؖy�>7�<����ʖ� 1薛-*�q=ѿ>��������Y�ӆ|my�KM	��_{>�D�Ub8Ɂ����Q��}��g���{���xD	֢�j��ԕS��n�j�15]T�qf���S�ɾA 1*���ϰ��Y{�;��ZN7L�+e�9�����{Y��� 33p�UR�'�/.����&��HH
T�Y0�I99��L���ٲ+;ڭKE=u��"��;<J����^�a���>�HD�s����֓�s���ݣ�)�wp�>��r}�[8��c���'�����ZW��J.�.�:����Q�b�D_��sC/��X"��8�Ƹ�UyE������5EzB -'�~�Z�߿�>�|v������q%��V����i/{<,�JQy/]���I�$��۬�}�Z����U�����k�qc�o�Do[���N|⯾ݙ3�Jx�YN��#d�B��4��ܵ0d�Ƕ0�Ѵ�RD@�y�:!9W����M9��H���쎈�3-ٝ]VL�1+9i5*�������*��S�N�m�4��]��BB��ND